BZh91AY&SY�����߀@q����� ����bB/�          Ξ�
kETU*P	U�P����IR"2ֲ�����ai��I@D"�0��M�J�ԩkU��hl44	{�9 ��*�F�Z$��6��ң3mKU�cf�f+`�llƲ�f��km�%KZ��[lY���ج�m+l�H�bӭ��m�Ne��a��l��*����� �v��d�aG ���`Q�l��l�	m��ƩUkk�Ŷ�Z�m�cKZ�kY��[jԓl�[� �S-��M6@ �JP� �G��
�� 먺��Vt鮝�����;k�۷n`2���kHiU@F��8�qh���v%ޞy5��Y�#QV��Y>yJ� �w�u��z�y�4 ={v��4��z���=)��^oyV� �����g�<��A]���,��< �*����US�Z�E	�+M�[1���J� ���
�G��tC��ǇJ�l�wAT 9��}��
*�!��  qâB���Ǐ@��җt�w�( =��< z7�*x��FQ���e'�T� ��|�UUK����AU����΀��7x���iOA����z
kJ=���=�j���������F�7 
zje>� �����I �Zik�dkc-�mDm&l�KV��P���J��tnWwA@�.�U@�n����(/Ms׽PD �6�U픠��*P�<ݞ�Wa�F9��E*G<^��*�om7;T�[U��5���a>�UP> ����=��PGU���@[�{�B��I�{�� ��t{��]�� ]F��ݮ�m���:�]	��F�ٚ�I�+i6���r| ��q�(�\ �;'� ;�Ƕ�:�Gs� z� �^�٠�̸W@����@�E͍�U�����d���e|@{�ۨN��g�v��@z��� s�q� .S���p(��� ��p �ٳ*���m�-Z����ʼ�y> t��Op z����N  wk� 6�k� 1��
8��Et�z�@i����ݬZ�fmj�+,m��ɒJ[歹 �Ӣ�{� �<�x��c�h:��������
�ۺ�� :m�ʭ n�r��`��  	R���� ��2�*��Ԁ�bT��*Q���b`a���)*T �     �O��%JT�LC��`���J	�R�� 0   &$��ҒI��i=56�S���	��MO����C����ˈ��%��i�}�״[�=�v���G7��7�.1�y�ʾo� U�DX
�"��@U���Ƞ�*�`���O�?2����TX��$���^�6S�E���~�����`��%�m�l[a[�Ŷ�m�l[b[# ��-�l`[�Ķ��LbSؖĶ%�-�lc`[ؖĶ%�-�l`�
alKbi�lKb[ؖĶ�b[L`[ؖĶ�-�l�1�lK`[ؖĶ�-�l�m�l`��Ķ%�-�li�Ķ&����%�-�lK`[�lcؖŶ�m�lKb[��ؖ��%�-�lKb[��b[LK`��6��clJt�[�Ķ%�-�lb[�hc�6���-�lK`[�F6��%�-�lKb[ؖ�0��-�l`[�Ķ�-�`��Ķ%�-�lKb[1�1-�lK`[���:alZb� � [ؖ�0��-�l`[�6���-��lJ`[ؖ��6Ķ�-�le0-�ltĶ�-�lKb[ؖ��F%�-�lKb[����-�����2ؖ���-�li��-���-�lm�l`[2�Ķ�-��-�lm�l`[)��-��%�-�l`[���%�0-�[
b)L@m��T�"��Jb��T� :b	lPm����*��� S�"6�Lm���U�*��V� �)�6�F؈銥�T�
��F؀�b#lD4�m��1�"6�R� �K`lUm���@�"[K`�l-���� 6�R� � `)l1� ��F� �Kb)l-���T�(����lm��A�
6�ت[`#lD�A�
��؊[Kb�l@m���Q�+ [`lQm��Q���F���m���A�*��آ[Kb	lQ-�%��
���F
��"[Kb�l-����
��؀�b�� �` [ ��`#lQm��(�Zb�[�(�`l�T-��� �`)��`l@m��� �!lA`#�*6�V�*� b#l�Q���U�
6�F� � `�lPm�F
�F؊[`l@m���A�
���ؠ�b�lPm���E� 6�ة �b�lTm����
6�Fؠ��� �`#l blb�lA� ��-��6�Fت[ `#lt�� 4�F� �b�l m���A�*���!��[b�lB��m���-�4��%�-�l`F�K`[ؖ��%�-�l`[4��1-�lb[ؖ���h-�L�%�-��%��%�-�lK`[b[2ؖ���-�l`[ؖ���Ħ�-�l`�ؖ�L-�L`�ؖ���-�lKa[�6��-�-�lKb[�S����Ķ%�-�lJe�-��%�-�lb[ؖ�Lm�Lb[�Ķ%�-�ldb[`��6���-�l�m�l`[ؖĶ�m�m4Ķ�������-�-�n�`S����-�lKb[-�`��6��%�-�lK`[#���%�-��m��-��)�Ķ���%�-�lK`[ؖ�����%�m�lK`[ؖ��&�l
`�ؖ��%�-�lalcؖ����IS�g���O��-�nT�H�|��(P7�Ĕf�4��d�̽jܩH,���R�i��Sj�洫����V�]�.�gX�Ib�۪~��kï �7���<��[�T+̕��\�C�������d��t�R�SxݗyV쥲�����Tj��:��.���������	�x�U]�ʖ��Y��ɉ�5��˷���4�j�!K2]U�۶CZj�jO-�nִdB�����j�9��n�	^(��iٯQ%`�Ѯ�U���j7@���sN�we-���Ӳow�M̻�D���4����5�Vj�-�09M�CXJ]^�ey�9�a�~�b���ٻ��c�̱�<�BK���i�0Yy4%��r�H��7��Y�q���>ډ�㥧S�ʚ��^�ɭߦ�s�l:ww�e�	w�&���w2��$��V�coK��)�/ѝ	�)���Zð�n;ܠl�A��Z[��^	�+h���ԈK�ѸK�����e�wp䲜�����6�d��E�n\�4��Ne�̹�H<2��r��{i%V]L�[W5��Ӭ���Md�Yn�VRȥ���.���U�6�md5��K֪˽y�ƺq�k�����jQ8������FP�F�̽$◫�d�͒ۼ�z)ъf�q�Յ���e��]�uB�nb)�O��*+"r�5��MT774�!���$��y��w���I&�ui7����ZkzJ�EZ��2^�3&إm����J����T����j!�KmN��Ne6��B̗�f�
T�K�,���-%W�`9�Tm��F�չ��P�0��VC�uHn�wr��ZT�RJA�Ö�7�!dSoLYF3�Se՜h<�(o����4�[�)�F}x�-�EǶ.V��h�\��A�Qĝ��iɎ�l�6T�&h��MRV��{=��㳲��+e�y�qU�Wz�tܙ���z.�{nc1�Me˫k�.�3J�Of��{�B�2m�TP��X�wX�˙��QL8�:��)aڗ�z�T��E��1t��증C��b<��t�b*[a�t.�f;�W�� ۷.IL�4��w��*�F�N�E1ښ�X�	��t�q��U���L���YJ��tB�7wW7�:�=����S�S{BH�j�/�+Lr]�=��f�Y��kJ�X��f	�aPj	pdd�� ��3TQՓA�];�ܛ��ņ�q)x�����E$eb��b��,
2���E�[*Y�D7GjZ�N�U����rkx�kK���Ï�Dh:�K��o[n�)�x-g������x����T:���7���2Am�T��[�ɲ�(��[����9˭b"��zVah���]_]#��J��,ĩ��+�+Z�4��h�$]�ܘرA��0�{ ��kSu��o*2����dm��4��Km#$�.�݌f��0(T?�iz�F�EY�����e,LXûL�μycÛ���z(M�L�:�Q��v��V�ou�%�xe«e�=�a,[����©�W�����N8���+#ROmJg廗���x퍩zմ)aZ��ja�Hb�i���-��DkL4�#��7`�i�k.V���ZY�X��n�GcV&�d���Q�Oo%i�(�vZ�ۻB@�fc'wJ�1���c+v�BR�!^=l<�����
�6]��a�X\HR�a�Q�.�.�M��v�=�岞���Q&��"�1j��l�B�v�&~�a+�%6���{��%ni՘c0��E*�0:Om]L�2J�V�RU�dE^x�5V�ޱ��q�$Ej�6�Tp`ƚy�U#"�f�-�ڿY�%�;N�����C$)�e��bщ=�9V^�Xvhsm+B�еYXp�l=çF7i�&t`*�4�̧V�F�2����Ά�'[�`Ĕ�N��׌*IB��X�є�J!�cX4�̦�V���A'm�a��`�V[k�6p �
�[RJ�d�y�e�-��A���V����S�+#���b�t������!d�Õ(���V�zb���D�3^�����rӧ����>:���;��7*�����i�eP�����f9�q�$��i�ڡ���(��h7�U�ۦt�*R�̭9.��U��޺pՑu$Q�����aqZ����2�"��J,Z�1��mc1*Uo#1^@�g�܄=�����
W���!�pL.�i�N�VJK3j��m�jjۼ�#�BƭM�dk�[��n��D����H�5��8%M�+�*�{��ԑ��
��w��ƴ��M7i~{Ǻ�Az�+qf�����[��i�YQ�3,�zV��	�$e�S	
�T�הQ�[4e�5��AT��]`�E�oV��k,�*�l��ö3ie�2��K&pJ$�cq���0��n6�:�̗�E�xw�����e�!��S"��5{
�q�"�ZZY���)���cb���MF�k��R&ۊ��ע�c�ej{�*�1ů^C���yV��yt�k"ih�	v�T��%Y/uVe�/wG����öLѸc�l�%P~�sn�ӣcRv�Yc%��D+���vVXa�����ɗ�-�AK+5�9,ؒ�C�]nT��os�*��{�@��X:�\�&C�7�7#9�[���o멏$�)H��Č���Q�w$�UN���Hս�7I���%�oxmɱ�9N�0�7�%�5b�B��ɮ/Q�TwH֎�[����N�]�ff&l;��Uh(����i�٣k]���eZ�VF�sPc7J����ɠ�Z*��M�&�ҍ�t6���y��a��ہ����)b�V��Y�<�¥֙��g�(�O_g�WX�5u��ݕ���{b���w��*ڋ\�d2C��z�T[��܃i�r�j���u��s!�t��cMG{*^�
��Tf)v�[jj ��ie7x)T�YeĮ�I;x�'{�a��M��w.m���Ze7��D�l�F�cfh�-%P�Fʲr�:5�q;4��g�f]�U�	��el�.:ISb�VV\۬H�xӽݩpҵ����f���v�^�N�BÅAy��̬�Yg'��S<���.�nX9���/j=uʆ�����h��9AC�������y��w]�I��MoSԮ1��%e�C��9�܏we�Ğ;���ت�M����m[��l7,��S��v���F�ZS��\wQ���(�2�e*!G2��1��[#h�X�1C�+'v�^�:oj]�;�$-��Y,+r�nb�kZ��7
���gZ����Mj�dFM���
.�Ijk-�L�.��0�/*�3Cm*[Vᵛ�Sn�f�z���r���gC`��7#�!HB쩗�OK*�t˵Z-��ak��F��5�ɪF�ޠu��/a��]�d�mm��kf��U!-LdWc��]s�a��v������6Zm�j�{�`۔��&�f"߲���j�&(�U���t�v���J��ąi�l��U��n[�ڌ֘�(P%̢)]�G�"3w,���N^�8�$(���͑��X!�f�� (�9���hm��S\i?��|f���R`�$˛(ndW-0F
�P塦F�<	�w���i^0�i�,Ǖ���bJ��˳��z.� �d�X����sR5-M�(鼬�{���ǻb�l�pc4^��ǌڄ�f���WPY��9*Mt����0Ͷ�Q6�Ƣ5+oU�ʓ��{H�췩$,���\E�z	���Axq$����le!��Xfc�U�R�]e���4��6i��ܥ�ر�C㶱h� ���9��-*Ь���f�x��B]�Nm^KʥX���Q^�=Cwd��6m�&�+Rd�w6���+I����E�J�n�x&KWM��Z���6���F���!��T�;�r���gC�n��
���v�M��d���RT�K�yw���ǐ��8�/N�{Y�MVX"Ѡ�-jd�u�����B�XT�TTQ+m��^(:��ܘ��/#��R�]A���:v�V�y�	��*�*����ӷ��{��9#��Q���X3e�X�t�*�;�îb�kU�u�u�S�� �Ȓ���G�\�V�k.δ	&\��Ej8퇒l;6c��)]SlS�� ��ei��0�fkR�sfL���K�� ۫d9���U�#`k) �u�" �U������v�;z�R�୸T�ʹ�VӐF��Ɩ�ù��ג*�eY+Ǘ�7F�5=B��Y���"�Z�a;�8�Լȍ�|�Lj�5a��V�-���L��y�jLymٖ�f�N�F���"�%��1,�����5ސ�l���Ɂ�Ru�㔦b��da�D[��X�F��#2��J[�����)�䦅cu�6�ZҚ������V���Df��B������̬w��Z��+M�A�1�dRݱ���J�6�tid̷�(���a+c2�͸I9���t��1�$��]w��{�gd&�x5I)�4м��eb�)V�V�5.d�&�eSѕ���e��^Ńh��"T.��uZ��´J�M���ݱ*J�ԩN�
1b�f��4R[�)]�o^ʶ.`ل���!I!I��(����݉7n�Wc��`زQ�	f,�w��ю�����W�'�ֵ1���X01���a��]�X�)B�<�eK�\�ʡ��ŲC��Y#�o�Jى�a��Y�#�٥y��ַRƊl�]H�,�{G+$t�*(Kt0��k?�72KM]�*bz�1�Wt0�E�C]ݘ��x��<Y�Fm͵Qʸ.���a��1f2�%6�ݭ����r���k��Ķ�n�zK�8fVn;0�+V�`xi��mQ�!���Y�s�SZC�Y�6��UO	ɶ�21��{�)��ǖ�:xѦ`����B� �k�ծ���m�+�,ǿ�4�EԢ�VT�[ù��� z58�k,n��[��/q�2��m봶��Z�ͽ,�%]��37lXR�1r1�v�^c&�Ŗ �;�L^���K�X&��Rӻ��viH^1R6��9�Pd�����+(c��6f���Bbcm��J�{72�-z���3Ve�"b�qb�j�V9\+-�ޥ[��s6�F-����VF���!����6X�9i\�N,���'f�㛷/$������"&�f,7�y�5X	������Ya�@��@��atÉ+!ٺ��	�MQz���2΋֭�5�j�z�Z���;�J�i��N�[H�Q	V�ԛ��l5�b�nX���)�ni���X��6j�wx^LQ��R�9vD;��۹�}i�͒U^��X�&��<�Q<��U/#��0����ͩ�ê�Kl�6;2��!����'�]5,�Ão]��@�\q�%G~ؔg1��4��vg`����m���̦��&U���Mm.�-<�r�n*�Y�wq�,�1L�����`-���̖�D��e�A���iܻ�
��ލ:*����n�J˲IDe�Xè
��^iC.��gb�3��t{ҚKHS\�k�]��u]wbH�.�ܫ}��#R�#*a �ACDbB��ʨ]`���7m�R�C�+�(�4D*	��ɔ�x+c�5yL^ʬw�Bm�-��Y�lu��	ֶ�㘮aQRj�̌h�#:Ne�,�rU6�ѓ`��ۻ:0d-�{�9J�8V��N�yTV���m�ZX;�ޖJ�w��Ul���N�Q�K×zpR��3�6�IЕe�!֍n46KUG9�V��a>��%�����tǎe����Ú��m���M̪a&�"�b�:���sx]@y�mKT����~����l�����2���Sf��wP��{g1խ#4�[�-��v�O1^��wj���OP�-V1��x�>Z+v\~�S�*�ͬ;f��KӉ"��f]�UJv���7�r�Ĩ^�hP[-T\ȱE��Z�5,��Jv���[*LI�Xq����u��2�\�{�I
8e;{�b�Q%IX��f��#!�zN����]�h뻩JȂd Rd!E(�I-�Ou	s0�ōm���9L�^wNTf�礝l�9=o3�y�r�������J��#R$��"̸�*4�"Т�Ⱥ-�(bukyS�6ZD���fd����g(M�Y��n�FF��T��z˲܂��܀���ũlH�C*�<�Ò�#���&�Ê�����2�`\Wb|�9Wq��֡���-k�u6��Gw��㹜V��+s-C��9��M��Sg�h.>{R�n�����I֓��V�2�OTIg#˱bW�\oc�Gp��"ә���cW�s�hn�P��(@��ڔ��-vڸ)˧h��y�BM:B�W$�5iWir1Q�j�X�����5M,'i$�}UIZiY�b\��f��A�I+䁻]i�@�N�b�F�.�jґLK�J|�.ԢQ0v҈��3s���������e]n��j�x*e�V�J$�4�̪�r�^��\��j�T�P��ř��=X��"����5�b;I\K�KN~�V�-#UӤ�X>I�X�w���rS\J2b�ۊt���cK�'[3RO/z�������6Mٵԫ2j��z�D*� ̢
�ش�/j��Q�N�5�jT����U)jR5�eś;cJJ-n'b�J#j�4�N�r���4���y5$A#H6�9j�i�qU��z�8��b�G�#m;Fײo���JK���]�|�+.7����92��|�u�&�jjT�4�IPj�r�.Qoef�%ZX���ݪ�yZOkn��r�E��G�bCb�S�����w'�$�e�j�[��MR�P��i�֖�Uh/S'�M.f�*UWz�Ԧ���ڬP���*-Du��v��Z�\�X�]R�;l�����jr1v)��f���U�1u	q.��D��i�6"ky�}uI2(�A�M�Hڭ�L�x�ѥ�u#��D,�cU8�6��0V����e0u��J�;#6�J��L�=Rb����郵�}�-p��#y�s���wY-�Z5VZ�hTɑ;�u;�֐��MbTlIؖ��<G��G翺?淳�����J^�����G������m�R��j�5:N퓳j�JXo`�En4�,���Z{�\p+��������R:r+�낕C���4�X�9l���w�uCB<�1Θd-8�6�n]a�i,E)��l�F\ȯ�Gd��^Q�<�mƇv�(u8�����9�
B�
ӳ�˾��q�Y,v�#�����Z)T��ȶ����ܬh��To���᩹���'⠵},�d��C;_tֈ���)�hl��=����@�NfJ�3�t����s���%��>�w��ʬ9ð�;	W�uv^cYrc�t�E��-1�(v2�Z�-Z^2�L�x���Ȁ�d�=���cs*V�N[b����8����+x�]��ǥNӕ|���1��x�������APOiH�lM:{���޶z���{�WJ̱���;a�Ӥ�jxy�vP"8��,�xN�|S=}�ccVTz���J������/jL:Ɇ���q��h֜K�!I��z�`��vIZfY�	��=��0������eS/eӕK[o3.���jWH�Zo�q.��e�f��yݓ��n�0A�\�k7������16���� ���h��6�c��rLs/0�P�ӻ��LNx��õ�;.ꥑ�uסه��ޒm�y�ۭ�	��3�]��2��CKH�UݜyK!J�Ռ�U�5�zD��{ڶ�lW��.�K	��ݸUc{�u
8�x�j���%��u�*���۴�ns�_,�RA�Uݛbyr���;�yz���R�n�T[a��q�6�E:�����{M�P蒻�j3u�-�1���)kՄR6D��;A\�r�8Z�5rC0Z�m�j��ox����h�Ia��be"��˪��Rr�N7�
ƙ�]�b�Ipbi�r�{��Q7w}s�K5{�IG^�l��7���ҋ���[0����"w�SvL3F�әn�w:iэ�Y|#U��a-ʥ�dD}�3پ����{rm3�nuj��u���Q�+��\;�J�)ԸB��6���>�3f�����K79+�/��4�=���B���{�j��ҽ}�Aǡ��FMp�+UI�*��)�Z�f�;�ۮt5�)�"p��^��\Z|�z_>O{c���U��:r��'J�x�9,�պ��qF�;�2�p_-�D��7�5�u���֝����h]F�x�u�p,�R[�
�ŝ�8����ۨT�P�c��M�W��"�9�w�t''M�ͱ��2�U�(��0�ް����
!�s���V�L*�M����C�8�kҫ�""�[�&��^:i�dK�y@�``��]��)S����&^R`��ö�ɧwnk/2�>�f���ڝjd�L	t3���Wʙ�r�]%˱�s�rq�Eq4w<AK��+l�f�He��$�l2o�c1�ƱK�WR�W�]m]�xkgc���}�����v��"<Hο�0F�L+z�x��������7hkK8�vLܒ��Z+��*�ؐʃ�BM�W�ܡ�:c�սV���7g��?���}8�kHg�q���D*��ol[�%��u��G��V��L��~H�{�goA:h�/�l�}ϖB�=(�uN@��wW��k�Y*�	AFK�䥒�Ǌ��4�s��wn�˅�Qr�ґOLG��wuT�%�d]AŦ�V�JZdI���T�[ڭ��c�j�x�L9:���縒���\&S�5f_0�?!݆���������n��wRU��ʩ;vǺ�_Q�+tr�X~�6��Z�\VY(b9��\w1{����z򊓬֮�{n���vPaqCe��r:!�o���H��M#gH(Lr<�}D�::TB-(g8at)��3����ׯ{�U�t����^f�\BR����J����0��,�GU֞�o`����]�1�`��ܕԘ�J�YٔwM�Q�j�;ux�i3�k�)�X��<���V�=�w����D��ut�ܲlԗ��a>U*nb!h����od�!l���=���Swv��8ݨ�1��ͿҒZ�Vn�{��V�QuU�:�NP����n�y�-i��61����r��
��u��ʣ#3_T&��[{%dj	:�V��f��cV���yd*#hg5g5��B�s��D�0��Uq&�}+��ݒ�.�UJ��i
�˭&��R{_���Ӭ��ٹ}�>�U+k|�t�Yl�&���A�����b]ì�xГ~]I�p�|�j��>ceP]���(�3IƮE΅�;3�nQ.��Dj	�.T4n��sz58)�; ̻�=����q˗x��^"2L}�﷗�]x����7AiP�.��L�ƋbA&W�n�[��32�g�/�-@��^V(�+z^p��
�ƪ�#�BҸ�]^��1'�ۡa6JW{�F�H[��Auc0^|mQ �u�i���#�*���(e�󛯎�TB��Xf	i���j�u��vTޣ:�=����eq"9|�/4�C#�m�k��BpR¹}sKt��T��9���ζ��+G;M-����H�:-őzR+w9L\�&��ލ��Wl���Ǻ��AL��������b*�-+�̝B���r�;��y+N�F��
�;j-G��F�FX�6�kO��4�T�:�<4�h�u�+8�`yυ�&üz[{�b�֊ѹ,�2�F�e,nΈq-�jZ뙥��c��T���ܐ��3���/h���3i�X5��-��	Go[O/��=�-VXн���Y*�}j��P��!ƅP��i��Lv���u�bۘL&��b�V*rQ�om��ռ�-��̎���X��<�R�U�Ұ�����ě��L���`���4�i�N�eJ���)�/4��1cvLBU���ͷ��]Ѓ���P�µ�T�t�}GRA`cG8��d�o��Kr�d/z�U�8ek�pM{%\�w�*9wFђ�l�R��:�*�Sj��]B���se��n�͊b��"]6f��n�{�w5:492�5��W������p�Ĩ�'�lf�H-YnpvLW��D����1�t��j���}�Z��L)FƹG���dC4�Vv��vI�|���ɘ"0���Իc���T�\�5wV��JVG�(�s]6�\���*\��}t���n��7�7�N*\yH���+M��N������mMҶ�ξ����nG6��<�˙��uS}�,�8���m��:k����Nt��^���z%J���MB펵Ty^[��l]d�׊f����,�e.l�Vu�n�h�$d��Į��	�s�M�A� 5�u2_8z��ʫ�z����r�'s��e\��?�M��X�a����X�δk���Ue���T��K,��CJ�r�����w��	�Gr�	�w�J�)����gg6ը��I&�º�ۤb8/�����8��uϺˏ��zsC�sS޻T�hj¶>�.:f'5�Z��֪��%*�}G�\ܠ��r�[X�w	�����2�Ҩ�E�˻����=�z���V�R�U�O!]w�$%NBT���n�%�anl���pOd7[���9��A����\u�Ne�����ByB�!�/�6^���Ð�MM�0:Ldl!jν����)S�G��9��N]��\�\/�.�B�gY��iL=G���n��絋�:��,w�ރ�.^vT5��ݾ�|:.F�m�2���L'7�Y���5�u�3	�������[h��y2�^�����X��
	�Jh�E���|���K;�]H�;x�j�c���R����w؍�gp�����gb��O%�zL�I݃�v�'dg*#5�e�k��-��S�ٚ:�7�b��'U䓸`W+��[|���ܡL�Q�g�w�{�f�Z�9֦�)q�78��-+fN�_P��c��%�A)�v��#<㧗�\�b��m����Y�����ИkA%��r�f��ї!���3.>då��Oe[��#��.�T-�-���V_�@x�B-]�%li�K��]�ڂe��;mQ�%lӇ,��4o~�$��Ѳ�yW��譶9du��U��9��vPd�=ƶ��b�-ఴ#����<�QhEr����Ae_Oq������k�ږCM�#�wZ��54yu��.�[�M��Y@"m����,)<��KgXλ2`[{8uV.ME�D�0����}xV�َ��̠�ݢ\�(���,�G��`�
��1�vr�u�yF�C����K�!�9��SewKL�ג�s�����ֆ�wk-��b����s���%�U������9;�[Ƴ�ݴeͬ�"�[��n�����u)3�����iV�gJ����e�ᥝ>�o�n"�lmM��;}�$7u�r8K��PRJ`��E�-�\gY�J�RR2�]�3�ܹ���T]�a�RZn�,̛��cX3�M�V�ʴ��E�j�6vv�Vۙk�C-�����o^t��ĝ�UN��2XZ8��y8i,7x4]��������ܲ�w�б�^��z��r����6�G���g3�wT\���*�a�sV+�����7�'�=�3�z��:.+��W�M�k��q̭�n�q1kA>'����̾6�VfvEf��	VV^���HF���l];UD�;���3J�tQX���6:���%�,�Eu]PiP���w1q��q��*����E㵛��4�V�����/p�/%c�܅I��{9GmZ�w��qLK�\�+���9to��a��G=�����:D���u���ڄuaU�ȕ�7GI/eSy��ٚ�;�"o㯷uP��[��"WL��~�i*�R�OE�yX�[3����l��Xf����Go{�qҧ�Tp����[�azݜ�]3Q���O�pT��B�d鈼@�_`֭��o����N�Д��Y�uS	�-�t2���vF�9GCm�ş���G:�Wl��(�qN
���<5�H/�\o���>�̫����ܖ�Q׬eYJ�k�Y��I��([]�Ygv��U��A�S���U��s],�;��B�JH]�}����F��L$n)��SY���+�ζ�Mt^��d{�]Z:���l�E-�;DBn�v��������,̰�B���{{&;��M�z̲ ��}�u��5����v�R�]������t�7ֶ�斻na�\�kl �ٹ0�ܷ����K
t]�Q�U�Wf�
�-L�;�:��f�]���+Y��N�w1m�r��1��e�Zs�)�qf���J�R(�Үp�/�8gP�Vgm�;Ѧ�����竷im������gigV���neDͬ]bӕύ9ݰ���Bi�aP�d��m���;�ѣ�&�M�Dd2mk;�9Y9_|[9V�
�~���d.���Sv�Q�-��[b�9�`��c�o�of���Eo[�o����<+�4˕�iR3��MVo#6N8D.�~�M�u�CN�Ȩƾ�ngq�D8�,Zj��[�#��J
6��ň�k�m��vr��[��咎l��j��Gu��\惘,�t��{2g�i;R3#�(m��:��j.�6kj� ����/W.ܲ��y�)�ʕcC�+�ݰ���!��3\���޴��'f�
�|��]��D�b��ثO7��"�RK���+o{��
+{tou���f6�̺07��$�բ-�m�˭ǏpU�/t�����&2���(1uu�r�d���R��先��áY�K������a3�����LZ8f��m>�X�6�K��Ǹ�37a֪�}��}�zqUX�f��CɄ\��SYү���n��L�&&oV��]�P����]��]f�"-��i�*�"��6�by�Ie�ꂖ�)S�e��2dfĲ��y����;�ٻ�ju�S�'n�/��t�.ssS�v���X"�e��ݛ��Z:C��{�u�0³�t�
r�Y|%�g�a�������R��20U��U)>����ݷ�d훗yIfÆ*��6r6��S��]2`1��%A�K�{\ ��bZ�u���y�M6��op��B�+�$��[X����S���y9$�Ȥ�I�]2�	����Us��^�H�ybK�k/}�k�@��%^"����Y`a��R������1D�� da��k�5�e�7���ƍ�u.��g��6:��rj &+�mV�,�{1Q�}Q�����|t2R*~D�\G��x@��v�(���,l�V����0\^��m�W4MV�Y�^$r`�
�UKS^��WW�y'�P*"y+�ѭ�]��V�yu{�7�(xY�v|:���>�eoA�<ו��A�ˢ�z7�
���U=�5Q�n�U�S�ʠ��DCiU�(�Je��>�[Kn��	�t��>D 	��)7a�+��]���#���ڡ��!X�d����KsX�k�[d ���`a SH���D�A�Z�����&�6r4�_�I�r�d.����%,e�k��N-U��.9�b�2ܸ67��u��Ӻ��H��\n���nȠ+��uV����#���B�����A�"�M/�Q#�%Z�;��Z�D7�הD�����h�(�ϟ�������>""�?�����>|�'��}����$����/��V�e�B �ݳM�>�8�q^L�A�tu�t�Th��`�cC�8���qs4*�-&�^mv�x�g4�0����g�k�(�j��9�f�rY/�+8-y���%%����H1$t6��p�ڨ�2���T"�-�+�Bw\GƢ�c�e޺�q�ep�j�S�|���z��A�
���[�\����8�j�tR�q�mnL����F$p��J�ékyMWs�ڕ	ϲKmR�Z�3`u��I�j,�Ă�L��~GK�w*E>�z�~�,�&Ibm�K
�������/��ΐ!�ܱ�N�5��_;����nZ�F��v���HA�X3Hb��u}}����G#ol��
g ��ʾ��B�ũ�y��<`ԯo�ܒݺ�=DO׫c�r�ہ�&;4����ܣ)�p3���H�xr乊�����DI�a�Bd�3 W��=]��k��8:���z��Q�N��yʩm�{z�4��Zռ��5�Ƨڭ��jS^T�o%J=�@�7��0��+F[��p�����|��Z|�Cq�ܶMEW�l����4qS1�Z�u�|�T���51���ȦF��VqYÝXk���|x8��q�x�q�q�x�q��t��q�q�|q�m�q��q�|q�q�q۷n�_]>��8��8��q�\qƜq�q�N�q�\q�n8ӎ8�>8�6�8�n8�>8�8ێ8㏎8�N8�8�c�8�8��c�8��n����)��7���#�8l�u���hn�ܐQ�H�8;2��i�櫢�!�^Wr��h�˻ԏ�h���!�f<����Fw��,�v^�=�/:,|�� b֧uŪ�n�-�=��v��թ�L[ש�������x�W]�w:VE����Ω�~獑f�s�G��5�K�P<���9|s>{`�h�n�J�j�@�}
y%1�|w���!U֎nX��/\$^�Z�z�35�-�0<��di�?SFEWݹ�A�T]S"l��-�7\�C�A¢�nE��ኹQ�xh3�ۨޑ�L������jr&��Y7{%��B�x��n��wU�m�-�~��z�r��`�ǌ�j[0��S���_j�(�iu\AA���\ڎ7Xҍ�D	���9���j�˭9����ʢMo,��v`'C}Ϡ�ƛ/���:��t�m)����5v�AXS��x��L��u.+UX��F��zi�n��s���*��r��i�0^�I4:�/j}EL�*��v�UA��YP�+i��� w�p��m����m����أs��[އ����T&s��M�<;��[w��b�~�T����!e�,�����#��
��~l������
�=��hZ��p���|9&�[��|��O8q��ǎݼi�q�v�q�q�x��8�8�8�8��q�q�q�n>���q�q۷nݻv���q��q�q��q�q�q�q��i�q�v��8�8��q�c�8�iǎ8�>�㎜q�q��q�q�q��y����w��c��=�Y`�)FUd@���· ���wCFfѰ�制1�F�u�t���'� ���
�Rhѳ�n���h�;��Vn�g8�ёF�Bc��M���'k��y�L�Ve�����QT������ť�������nO]�d-���A��T���Ҕ^�8ս�+D���ʋª>�Kw�ى���Rv[��l�\q�N�wU�B�K\N���ѷw"��"ݺ������L����K-rV��u�*ץ�*���u���;J�Wgb����jMn3��rX���֩�n��C�D҄g\��J=74�V�jۓ�wI޺���}gn��%�Q�Z�Wp�{ͼh*B����:��f�tK��Z#����ۺm�UV�0i|��Ўcw���K��i��GU����BZk�z��U�e��d͖����I�ZFӐ�ͭ��ظu����Y;T3�[���0ˆ��7j��º�|z^���f�!sa�jx�J.F��8`�vH���N�,�-2�v�F��v�@��5n��Ǳ�s+�_\��B���U#S�����o[P[�ͪ���}w����{}Ϯ�v��q�q��qӎ8�>��8�8��q�8�8�q�q�q��q�q۷c�nݻq���N8�8��q�q�q��t�8�n8�>8�q�q�88�8�8ノ8�8�c�8�8��q�q��qӎ8㏹{�����ٗ7���ܻ�Z\����2�ᯠw�K1���r	��=j����SvQ�̓��ݲx�ɔ{�^�LޚR�Չ�3�������x-��f�S3y����t-�7�K.e���u�u���k1�j���w��eZL���H�c���Q��X��Y[O.�Y�ۇH�zP'VT�����b�"�m����}�1֤h�:5��|E\y.�C�����Ҋ�*�6�Z�ޤ���H/�aٗ��yɎ���@�B�Tk|�23�m*��e�cne�L��o�!kJ}}:�!��k����#Ul�{��:F���-��ۆ��	jv᧲�s8�uZ,mg�&l�2�&XɅ0+���yU�E�w�%M�J�u8��Oc�ǌ���y��j��ٓ��nWIż�H
�޽�zZJ��+���ТSCZ�^�����ꗑ��g��Y��l�����G3��ͤ� �m*���_*��7�2#en�q"��z�Cb�����٨T�IWwkS��XK	���ףP_Tf��q�ks��b�Q[�j�ОֱXäI"O�d�%>��Ț/��@
�7k�2��ƚ/Pr�岨�j��H�*�K	.���Y�|����gP����3P�HR�6�c�W�W�����.޳�y}�kԧa�;�=�+9�'����w��G!7�o"=�o�#���u��Ü���S�i�n�Zi�q�]��q�|q�m�q��q�|q�t�8㏮8�N8�8�c�8�8�۷lv�۷qǎ8�8�8��8�8���8�>�㎜q�8�8��1�q�q�1�q�qノ8�8�88�8�8ㇻ���{����lX�W��H��m��@Uj�K;}&�ʝ�FF6]J
Q�0�hz]�I�AfɻWN�cB�m��b����j����vh����FP}�s��C��x��@}y8ܣ�mV��ڍ-bh.��j�V��Me��Ͼ]�RX��e귃Q����Ӹa#o�hm%��Ss����?��ile��ګ���;�Vu����MA��5
�J��4F�}�L��.�ìś��2'�b��uwK^������xi�5+R�ؕ��� �B�6�i5����N؎���B{�i�Z�p�3.��xx�x��Z�Q�غB�'aA8��o,���n���wOu����7\�%�Κ  i��ί��,FQ#Bqv��f��(��Fʗ9���tz`��Yn��5�'��Bޘ`�8��=�}��{WVnAlٽ��y�N�POIo�z�n��7����� �1�d�U����o|B�#�]�M�u���^�,�YZ���u�0��[t髚�j��b�]ܶ�7bZ�f���7zK��>n��u�#�}�jXr���i�ku�ԍhQ�	�t���:�Y��hd]`�9�/�[�S�u��W	���.�4�����ID���Ѧ�lR��E�YY�z�IK11T�6��,����mY��!��Y����#3]Qj��I�έT�'u���Z!{Q�M*G�Y��
 ��:����`2N*<�n�9�{��5VNCJ5��(�̎��/b��r���`뷘O>�^n7ܛmZ+u9�VH8~�s�P���Y�W�W��芦��4�x�yj�w�����r]j��w}X���%�vJ�ӯYA�|ipÖ
 _��ôUF�Q׫�])�.�����T�]�M�u�Ζ�������R��n�:ǹȻT2:vj�Ù��(��X��V���d�N���F셣4gs�y�r��l����X$��$��3�#sT��p�f�Z	�B�U�4��:�Un�	X��WE�nt�E��t�L�c�w�5���3I׮e��o�y����[}�,�)gjww���2����>,n]݅���"V.�(�.�D��6�ǔi�
4�)����UTd�����n*��M֝Mh�b������n� r�-U�ɭ@�e�T�!�6g.���^l7���T����X��-�YJ��Ńһ��;u��
��*�����]�n��&ӽ�*�ٷ��9U�y�E�%�5x�C䀼�T�܌�%���Vv���Y�l������ǻl��l\U^L��<�[��1s��ŧ��3������k�`��WWE`�]����Z�mY��wJ-����e�6�D���-��Vx�ˉqqC&<Ԡ�᷇>�������*�6��Cp�s���_��h,U&�(A���6%
ݻa��C�Dl��Jm1�V�ƞw�yM����\Q��G}p��ͼ�;6���Н�O�+&�I־�5y-�����v�Ѹ*�Y�'ڍ�'��.�l\���+�f3A�R�k�����1>t��d�Һ,Ԋ5��k�yx%c����<|������Ee`v3��c�\jӊ۶(�q���c�:V/�-���M.��5�D9
��VX�v�S���ft;UMU[�ͧr>_=�zwc�ykT�bw��)�#ڻr���+3Uv�֞�2@k�滥w�_�+�75MI�ǽ���so�h^S:"��>��i�x�gw����Y/����������$3-��	���ڬͭI�RV2izq��qv�B�6���-���3�N	u�c�dL�oS�$�N���7Y�I�\U�L �j�덚���	��VOe��Y
3aaz�3S_U��P^%��d�N�-��R%�ϯo���s�r��s��@�����]���8�{yLf�"#�-$=;��v��%��qf��?2��,ڗ�X������8���)N	s�n}�z������Au+�i�}x��g{�=��Z�h�>*J��KfS��UGe>��*%E�,z�l��W��U���]C�ޜ�|[(��k�UgI�y�ݚ����Ӊ�kWdU��0o'�_�'^���٢E�OS�LO2L��Kv�ݙ��V��U�ע�vl�n�	nt݇e񳕚�tKʧ�;���|�w
%3�����Z�Q��d�Cs�*����h�\�C���j�$_0`.;�vM�C��F���n;���kfӲ�9Ϯ�Wy��ݯ2�L��2���ft�e�+�)�C�&��8^QZ�N���D�偪\�e�P��ƥj�%��ec����UNH��A�+:-��Vd�}�6��;*`7gB�Q�r�N;��2�M���f_]��uVtM�[���A���3E �������Wc�4��ja򚺒]���FK.�(����wx����EuZ��okI��{��aȪ�<�9W�&�C�U�ZP��F�Qj3�:���^��Eʮ�1#������l�p�X�!��Z͸E̖V��3j�qo%��ӆ��M��%�#|3�����]�2*�il�"�>�����ʙu�VS+5�v�eJ�s�����5�T��T{1LxGD�
��h!���%R�*�\��i�حk���_1��°��Uc�V�[9Uzv���Qf��'�eJ�m��y(s�v�k�E8�f>���1M��˩+�7�z�X*�b��-�U4H�^Wr��r����2=Q��쩭��S�p&��ʃy��.���E��yw-<۪X��2p{[>���`��lP�ԩfN��U���.,�X�S7}h���4o�oa�t�˴�A�ʝ��+�k�^ԴqFm�ݼ(�s��ĳ���x�A�I^Ib�%y�{Ім��1�c&��!%�'�f3��ui7N�쁄.آ�]+�-a䶲��>�q+���&]�hʹ��)X�}��>R�9b�W���5��F+lm7|���roLU�+܊���:�t���늚7����o{/aWnYo$�{��eЃ��7���٢�jdZB���^��7�x�$%E�M�]��y՚fѕ�i����m[#<����Ӻ�G��*;�YV��w����I�q�s��հB��y}&1ζ��&=�+M�of��|���0�V��u�&E�hk!q�<�]�`��yX�\Ba�:±�vUTcm�;Gp`CvQ��u��1fM�e_,U�B4�V�\�s�$�+0����IP[ (��lM�����ri��>+��Y�])z�c�i��;��(p��"ں�Mq��V���.���M���U�b�핃F���ݼ��.��'��]�~t�?�G�j�G:�T*�uj��l�R�;�v�;�t&��0�yLs�1���X��l)��]�GP�N��N^$��jmQ���Y�r��J���/�^��ץH3lՠ�$�J�z�ѪS%HĲ�"�7E�̑;n޸8u݊_;j��W>}7�u�33����c����KEf�Sk:R��9d}V>ͫׄ�J1�o2��d�T4=��GaZ��ئ��J� �Rf�٪*�+vw�Jn;i�d��Wʝ��qn�]Ʊ�qq�t�-g���DUf�e[�[��\tm�h�P�L:U+�3�:�Z+zJ���D����f[Ն�e����7bS#�\Y+��b��2����(�q�Q'�Z%��̣}P�<[dsrأZ����d���gj����soEa��id&U-M�PSɽ�)�mYy�5���kx��0Rҍe��y�3��Жђ����4�e�+��J�YϺu���Ty�*v��psE.�Ec�*�����۹Wvw�U��l����P���ʎ�d8�.jb�#]h�ò5�h_o��04y\�Je�����{e��q2U���[ܵh�Zq:ܲ�6��?��M�fQ\
6;Y�zm�D��e<O��"hh�sYǰ�����{>ݳ��ʤ�'��]S����ŒM��|�w��W��?C�� 
�{!����������j��#��$���?�~s�g�yeh� ¢'�`��/͗�&�M��C�Ʃ�42�H�m��L��:B:NJ�J�i
��衒��E��(& 1ȍDBj1"PBS��8Z��QƩQ�1�q���J"��nJ�BR��h�$�2)[B�Q��")!$XN��# �����&���1�e��"�&)K�`�r��FC0��d�8�F9�3I�SD��
��z_�{�w�(-��r^ʽ[�B���A�[�q���U���'�Z��O/�Zv��U5��}$C�t���L�|ܩ�d�qY��N�"L`��v�z>�HbŚ�Y}Q�y2n_fK5Ҷ�F.,!��<��fs�1ͳ|�s��,��}��5����/���q�B��姷1:�K��3Nۜ�*]��N9j.4Wrt�e�W`�,�"�5���+��wG:�f^.6�mզ���Ś^!3�r�֤�ųu�:�q���Pɽ�o���3u֠�]:�t�Y �HYR�q���٭�׽�guƽ�f6������TM�&�Y�:2�^7̪����J<ޱg�:�F����e��b�u��Z�-����Ʊ����7y��t�I�TN=�\p�j���չ��M�u$���|z������j��wJŇ�2�}�7���)or�D�=X2�P'gx��Gy�.nL���2��M�88d��a�8����w���Χ6�g47/��}��*���\�'�-��I�y9���L#�
�\q^tc{����'��L��L�ս]l9B��ڴ�F^��9m������f�u�h�5f�E�����
*6�I#
a��M�"���!2�*	#$`�)Q��h�X1@�D�NC'�B�B8 -��� R�a��*�0XHF�d�?�YU4)�.@�!�d� r\."A�$�R"�p�	E�L�(���qB (9"����Tb����aBb��*�`��&��0��8� ��"A@�h��L�g�DZ�d�aU?&�o����F�q��4Q*2
��D��IE2aL��L[s�D@\i���iU�1�	H��6&#_����(�ڤ�rB�!��	i���i"$�
 ��0�F���!��SP�#p&
#`��%�$��	0�AE%!�B(�N4�m ��Y�H���	��a��-�R&����vC)4�5$�(�wh�fB��[�}﷎ݻv�۷n8�$!$��^�wu/]�O+ˮ5	}�E2��p��I)E�iD��q��nݻv�۷�1��	$@�I��L *)�s�Q0R�UMQ
��j�O^�z�۷nݻv��[�oU�CF�]=�1&�\�C������Wn�sw'W]ԝõ�s���wk�ҹÝ�gup�d��$a�5*���ǯ^�v�۷nݽz8@!Х*T�J! F��˻�\Lm��ݹ].\����/�nwvۛ-W1�T]
��K�[nk��.sx�]��r��,Uwv�n%�q�ꡡ�.m���s��%Wwp仳��۶�ܸ�uڻ��n�gx�n�˸�s��vN��]���]]uȺ�rN�q��:�<�3��ˎݹt]�]Νvjy�)�<�:\<^O��9]���u�
e��1!t톙��x�Ñ�&PO&��Ρ%h���qH"O;�
�ۓ2cB� $�#	�#&��
L���a1$Gn�oL%"���u lH��ՠ�Q�OB@�CkQ(?Ɉ[��n1��M2$N8"��Fw�ٮ&�yˋZ�*�9NÂ�:n-�q@�*�����M���b�2l��#a��^�p�5n����<[UU����oYf �$8� ��#L����B�Ap6hQ8$@��&!��l�eS	���La�K4I�b�����=�y����}{�6<Z�n��i��H��%[��y�Ǔ���yn�\S�hl��p��O
ky��{F���h�rLC���{ق��^�N��g�ۆ���ʙ �^c�Ϟg�}����n-�nk�����.vn��u_��.@�u�{�k�j�O��׼@L{g+�{<�����z���u+�t��COX�~T!����3���*Ț��/o?S�3���̿{���4g�"<l�
�h��������|��6D
d�Ŵg:x֗�\u�z��.;��i��v��������	�g��!vzg�ݘz��`혦����/�s��� ���g�=¨�������yP�(2Jn��ݜ��z��ϙ�7I8�Lt��s�٪��_��2�J߂���Jov�߰&K���r�"�-b�X�;�{���Q����[v�t��E��1��4#�L�w�����s�F���j�w�ޜ�����mk$��2�MP=f'W�318顱uqZJUfv�*�<�:ݩ�MVWyȔd<�*���|�ޓ@�]�*l�y�uB�>B�upz���`�������h�u��GD�q�g�}��F�Ǫqoؘcp�V������[�{��U��\Y��:��=����~O�J2	�KȆ��Y�n��"�5��4*D���̓i�O����_a	<�����JK7�+�!��@ �e�o9�c8��U���&^��|�6g�[H��/s]G4螘�.�4ߵ�����8���"#ƏH�<����9�=�۵զ�BB�{�[�%TM��V
��Ӯ^c�9�Ż���<��橈��x�&s�Ir�L�rg�˒c�k?Zf�|H�}\п�����5��U�:&v����(��we��;���z{io>���M����bƼU��噖�\�P�7���l�$�9oq֞�;��{V���Ά���̾�_]�+��mG��'Pߍܒ�CF�Y$�70��v5(��qUWq�ʦ4��s;��G���[q)o~Y>�#�<YxN������˔紏kg|z1�[A]�x����+9�7�V�zxKZ�c�d%d���hg7zǥ(����-1��e�W*�6���"��8�� f��gQ�a�ǎ;DFO�)��ݧ����~�����yg��|�\Gq�N�;��lO7w���]1�����"�=�@�e�� �%�}�}u6�y�%)�s�U��s�Mu��ç������_�mw���'�X���]��Ql���r��ݲ������Ⴊ��.f
��[jG���hDR_��ǵ��#�ϙN��*���ݮ����}�O�S�)t<�O��"�W|����>Ʊ����nzߞ�(�~K~Cx��~e{ڞ.�۾�0v�����8\
�{�d���N������?xg��;|�,����8�׻���{�_�=��8f�vng�߶Bo�E�ƽʽ��B�xy.#�j��F��@�����Uv`]yi��Z�sE8�/e�Herl�wh�X�8�;ι��Ǎ��l��Z���%E��p��5k&��tr�yT]m��A�j�]�g���:Z���}ȚB���9��Cn�-E�ja�kE��Jɓ�g���+E` d=w�d����?vB'���P��o��{O�2O��n�X/���t����s�����j�{��&2;ð
�ͫz>˱�	�?W���қq=�0�S*�V<�_G��ɸ��ݦ��Ğx�e`ܧ����M�~�ޭ��>�<S���:I�<Hמ�N�!��n����1Vm�@��z~��^.��g�<�ETW�\�򪪌����Jej��P?D�k�"����g<�W��"4�^�_�q�;���]�wxsֶzC�vm�Ǜ���9��9q�r�Q��]��_�����k��|����)6��_h����^���>sS���y������o�%���OI��ydE3O�ޕ�����,]�(��G>���|�{>��X��9��J���3��#���O����M�Yfh�qT�h�c�p�mNxS*�r;˕��θ�!l��ʁ,Nh���Ws�����Ƨ�d������u��%`�iȊ��V�v������T̈UYT$�:N���NX�;��v8��{,r���v#�$����!*W�����'sm��;��e'szoл�{'�C�˲3x��ŒI�`/�`�������?�4�N����y�`�\�_{��z��t����,z�C�_���.A�m!O������.�N�UV���} �^t���7�\�E~�r��N�I�k�l���xG����kk�$0xzA�=��Le
�����T�Z��x��=�C�>��J��k��|��j��T���(��QKrQF����4r~� ~�X}�o>���0~����������wC�Eߑ1U�K�W� ��E�צ��,t����\�=�x�.٧X�.��Ɩ3��@sWhmL���)/�ox[�w��P�'�Z��n`��{��$N�M���jw�9&|�[-T�(8��G��>:g��3<�{g����y�gKʦ�xo�?O2����7�#��:=��Z�mN�2�o<zknJ�'�sO�6��_	���B1�qm�v6���8���^]��ث�+�z[�7��h�Jȳ�H�fGU����E�V7R��>�R��oK*d��N��.Nۓ:�U����AҤ����}Ō�Zc^t��^^b�_o��o�/J~�j�v�����03���径!S���]��f�5�K��/�m�s�O�;(�߇]���O
���)$T^��#Ȏ��߬7����z���!�q�{���������k�`���d	~f@�/�	c�z�z,v�f�G�k�uU�u�����7��N�i������$?V,|>�U�����z���7b~͕�g��n���)q	�-�`��]p��u>��cm��?O������O��H�v���qF�=�N��<�P�$��j����c�ۏZ2Z�=g�zR�Y���^GLĢ��`�$�e;69��>O�I/*�6��?l|2�o���}������b���v:c�n9��ֻ�a���,F����<�]�XxO�W�H0��"z*�#L=��b0e���"��C|݃�n��;b��:���ݢ]�U��)т�y�ƨ�X+�� �fʢ�ßwI՞ }�:��]Ҵ9���׎���zZ��&���F)D�������RTJ�k��DI//f�iV�ym5# 2������̪��[�ܸ����pίM����L�1Mj͜=�Ϲ1Ʈ0��8��D�AɊ��g���9�W��^�<I�zO�5��~��Oo��z{v�g���{eX:���{/=@�t�wL��!�l������:=��I�h8'�"=�WT�}��K׾���{�@3hF��_�����[���/�^F�:A�r�2��Q�oG�������O|� ~�#c�0F��c&��i��h�<�kEE۟zu����sw�J�5���_{+��O����Fc�����-�>��k�e{�^�߳A�㜍p�@�|�bz]�3�J~�i�w�u�h��]���ݜ)�}���T^Z��G�@E�ȧ��+2�U�����|E{��n���`��]��6%�\�t��O�����/ʽ�u�m���f��fo�o�5��+]X2��F��x/�r�^b+�٨�JB;1]P����̷o�֕dCz�щg'�m�Ȫq�ҳU�����%�r
5�etзpvR���K:1���{;r ��"z3w�G�>�\�5��q���>����>V���-�v�ߗ�:�W�}<Jt|r�!v<5����ｴ{�Y�0�� ������f�>�3Mk�.X^�����\߰X�U����ӏ&wY*����~��x�Ҳב~���';�[��G��zH��~v�!{{]j7n�Y��d��ܘ��;���4=�����tz���n�h�^@��.t~9�ü�y]�7V&�w��œ�3��j'�(�&m{�XS#�+9�3�ǒhOa������l\I��Y�E�;���5�
��z�h� �q/{����%�U0���~����q��9������P��륊��{`�uv����\6�/13K�|yG}�ז��gl�����x+�f;F""�|V�q�y�;�2�]]�O^C��$g� ��Z�K�7EZV�"銺V���0a���ϒ��L��a��ܩɩ�1�-���to#K�*͗������K���&䕝��f����F�9*�����<�V���}w��Aϛ�#ojb�a0�^�{���Px��ZŏZ�u�wI�6�]r�$��:�ky����Ȓw�[�=$󗞺�g#�}�D���I������s�����y�M��|���>���� ڰ���|����Y�����?_cm��7������[���I��)���m6��GϦ�$_���09A�:g����wڟ��5|�q�꣤����'����3+��!?�y���`�+����}�l�zk9+�DoZ�z�{�쬞J��j�8o��j;���!�/=���]׼k���E�^^9ތ���v���w�Zw��>_j����]e���a����|�C�K�ro���4��,n�Y]!������n���U�b�r���W��{[ٞ"�
.��u1�}��9&!z��N��t^{��/nq��-���vt9�)��tv���s ��̯h7�OQ���t����|�gث�}\S�Z�K�\�;w*�b�g��KTc��\J��N�2���.��"�Wƥ�����	|7ӱ�Ƞemo�׶i˩O'��5vG5��2o)̮����W-���(��U�ae�6�]�����勒c�Z��,��FuL�uWcެ��r�E���[y�ڸʳٹrg���ȫ�ӱ�o�G��p�z�N���L6h���A�$��)�^����u���ߖ�u�����;�=�5�V���?zx��4߹P�7��?q�ᦴK����Ic��Xf{_����~�}��1PV(��z�;'��γ/��I=�f�ˋ�j�C�^��<No��HW����ɴ�f��(���.׻OV��}�a������ך����G�9�N��y[Me�2�9�v�p�Yg4�a�9��p@a�7t��=����g�c[6x�i#���2kc<���az�n<�~�wk�y���l-��H'����*g�ʞ��w�Za�c����@`�}PVܾ���r�od�D��%�x��g�bm�K´�@�н�<���C�����͝��C�5�ß*��u��sTh~�e~ջ��6U(ȍ��t�ۗy�y�UPƹ�e�|�;�q�Z�鐻��%���{����}$23�g�UDU��zxDs&�qU�,�!���.ݹ>��Hν9�2jųZ�u�%VB9H�{C!������ͳ5P�{�^����tOpojD�3[�n�#� w�a����/a>�eO"�:k�oM�]�.ȣ!u0K��ˬ��R>׼�M����	��ؖOIK'��qި&�S39�����Fv��˻�ej�|A{����|��x�����v���͌Ã5�ĥ�a8�\i��Ti���c��x�+��65M��q��廅5����9Y*�۾���LÒ�v��jwRn�95��p<;:����*���+.��^A�ƮMC]��؈=���	.2Ǿe�����Iږ�SdF�9�\m�:��TVco���3��tb��k��h�70��$����/�6bΓ��._;�f��⛬@n᪳"GS�n�T9�r��ۅ~;H�=|�bT�A*�}՚s^��	�bfƾ�m<r�~��-�U�!z�j�]ɼ�] ���ݜ��f:��� ��3���uu-Q��r�0�R��V�I6�E���Y�d��CQg85Zʾ��oxd�uW���)R��s;4s���L��F�j�L�(qו��8���dn�*�mb
K��)v,�.�h��o��L7�s]����=�^�׹�8K8oq=e�Ywu��O3��I/�va�=��΢�j��-G��`re�`�c�&�P�7��*����|�l����#�Ӷ*�t��[�4)˘#�v̚R��f�nv4�n�ۂꌅ*�w�	5<��eٷm���o'&����ż,�P���P$.�[��qs��X�)Up��a�j��V�ʳN�ַ�6���A$���=�TI�7V�&˺��`�M���.U�fڐ���Z��{�N��*����ZS}�r��Y�;�w�Dǝ	��l��#���s��h3O���k{xջy�ɨ.�LaP�mY��r��m�U>4P��
�Z�[��̼c�����1�"���V�nKn��ڳ�i�Z{VM���X}[8�,q�qC�5'^�O�[�B�^�We�MK{YJ�{ܵݪpm<��%)�uШ�\���*g�%RJ�f�.�/�b|->��7[u��$�Nq��GS�8�s5��d�f^q���o213:M�x2�ΡW��_7^۴}��9V�][��a�����)Lڊ���ɭ*%%
慪V~Ews&е�9�d
§����U�v�Cr�\a�oSz"2�-�j���V�,b��nv!���u�;[��FM��w��y~&D���0B1��W�7I"�p�#$$��<�H�M���<q۷nݸ��ǎ=�c	I$�j�!$"ĞNБ�H�|�c)�B$���o\q�nݻv�۷����2Hd9BBHI	4J�()H���z���nݻv�۷zǫ�Iں�A2|�R�R�e1d(�II�޽z��ǎݻv��ף�@ªt�d$��	&�!Dd�}׵w��+��/vT��n��A�ݠ�ꮷ� '7Q�h��ݞ��"�#I�����3
(�����R���ܣi��	��H���/k�(јA��|.�"$@2/��a(��������w���Rj�#z�Z�f^�s{F���1�>0��tė�;�����kh��`�d�o<��3[�s]x�1�`x�J�s+����Q<`�����8��f�E�$8:	5��p�lz�=�p.�D����1Rfz�����u���pa���n��U����Tϰ����ǯ�07Qa(��/���8�ȶ�m��&&{b�B��}��Ͼu� !>
Y_1������/ml<�ǣ�i��J�Wb�ņM���y���n!�B@ vl��5b����R@1a~X��y��KzB{`M\�ƨ���[��vVR��؝����b|���s�4�k`#)׉3���-馞Ŷ�<�AG��xav"� �AlB+�E��Y��[���\	d.#qG�X��Q����* Uo����� �>W�Rp|���.E�6;Dv�uO��/K��X`���n> ���~�(�*����2����p0s�������
¹D��/�Y�u=��1�2�^ ��M�_�s2�HL��w�Bb�y�57�G0�����-�w8�S-;�CGw9 �0m�?=�� �#�7�L ><��S��W?�Fo��;��8I�No|�|9�_�s
����;�����������i�io',�<{�+)��t�^<���E��S�ry}�m�^���;��I�_V۸�M��uޒŪO��W*R�\n��fr�uh����*��3ns���b1��{�w<�(������=U^�^4*��rW161�X��:��Ò��Z�`�z��r��M���L��U�c����9.�~_���q#Č|�9yʮn|=��X
�W��I�K߲#����[�J�, �,�~n4&|'hB�T
m����3<���ͭ���� n?���'���	6��7��݌�υzQ�
��`p|ןC�8��as�Z7f�nn^��Q%�C/;��ff�l�͐Xbc�,\�[�wAɳ��)�S��,�8D���b���
{�~��Խ�(4���s�.����FI�	�:���5����x�T X��q3��k�\L��è�@�3������`�^�c�2Y��_G���s�p4�NÌ;x#wl-���;�-�����𺷶�vD����2���y>K�fyB��<��hM�k�/�l�5�t �$0=b�j/�e��x86|��	�! [xC�["�ަ�X��|i�gH٧����t�^ o8����M��QY$5g���i���H��ϋӼ,:N�y���0�Z�5��D�,��2 �wُ}�����q��2�o8�>Q�nB	�,�,�ԑ�`������sCo��� �b[ʲ(�ի��Ug�
������W��,�|})�$���޿�����R����-��/&o�E�~X�f��>��j-3�j�P���O��ۑ�%�(��z;�!�Ⱦ�L��V�h�Ukگ6�z��*�]��	'm��53��<x������2K�2^�*��B�{�I���Aͺ�ϳ��{H���J��t��+��L5����)��[��ϭZ6��x�������{�*N2t�/�I��Y�)ϼ=ꅑD���9o$����ѯFy�Å:lk��ߢS�)W��2��Q�"Pނq
��@xk��Y�hO�������@�{�:oP������	�I���&-�3e�ٶ�yo���}~^���z[�>	�,�D0����̤�
/���Z~�1�Ay���U�.�g^�t��Jk��4�x��7s�1LS��s�-+y�ii�$Z��_ˁ��~��zv1vɃvv�^mt�{���e���+���� ��* ,kˍCxJxw��`V�?� >;�xf|B3�l� V^�$��zXSat%���X�5�V6���*i����f�V��z�csH/N�G8`�1k/<�-]=yT��٢������9a��t8�T��SlipI��������Q��'ju��b2l��Ъ�gs!���Tx0}�gC}f��А��h�˹��Mz�����m���COs��M%Sjm����e�{�:^���;Gg�h<%�r�����f�0�ȚM���q����m�߫��k)����%=�F�A��xo<ӫ�v�Y���t0!�sW���1����?5>VB?�����G\�������j+.�m�����U��.j��uH���o������/[�/n��]��/u�����i'�Ks+��b]݅
�[�v@{��}����E��=�����]���EXu9�5�K3�q�vJ��c1��s^v��Ө9$>]�lM�ߘ��Q�a� ��� ��x���k�L�H��H{.:;h@��R^��< �|�%z-ޚ���Nd.xj��M�d�8$�y��_�L\?��C^��u�K�>!�9����;|������q7"U��
�z�"m��!ܮ��^c��8��ئ�8��k?P���v; J xc�C�ygo C�h���	��)����K6|���)����3*��^�B��Z����`�*�l6����Μ��E��5j�3 ,��H?@0��@��l=�
���<��9�tG�74	�Fi�/�B��i�6 ����������V�+��i8��}�#�/��$�Ӂ�Vm?t��=r^&C<w�ǔʣ����	n/z�
cID:��g_����U1�+ׄ������g�给������O7��/-���f .��)�3��<�#���o�:fo�zk�.�/W]tFF>���=�ݼ����	���Y��+�ކgk���X��Zʂ���%ߚ�	l�~�N�WR��P@x������C����p#���6����<��⏩������PWC���)^��lL+�u�R�~���IVB�U�mv9A+}Hl��eJ4ER�yE���<�q��^�7c��݅�؟V�\��ӸK���Q}f�xJ�^�j�p�s��ȥΑ��)�A�ݽX�)ot�}5�av6�9y����\+^o�s����1���s�g�gftS���O,���k9����\�Y�c蹦@ϲA��@q���P�^eѨ�쵼�5=m�ի� y��u[~��66&B�@� �K��U���D�u����������TZ���ht;�xa0*���|o Lx�� 2�ۤG��0h����FƎ�V>�H@��jKYp)5��6ܗ�ƕtId<?"b�G� k��Ob���Bō��z�E���ʺ���¸�~��9��55�A&���5�p�4�z&=̼���.2��l�_U��u�rC�q����-ǤlEC���>��B��L� [k �PX	�z��7���O����'v�#u�A��	M{�e�Lt�_k���xi�痢��
`!����p0!�-���n���硎�yr�>`,�$2��hM � D*�4?pDx{u�2܏,p�Xt�|`-���S�Xk�y,2G�>O��$yS^ZF�.m���G/v��`7r40�Ȕ���xz����ʭ�?��� 8CK��"�Ǣ
�U�V��ޮ��x[��#��#���H;�Y�I�(YH���
9������^@V-I��?�������Y��n�ͤ��Umk#�:�ɍ��H��C��	���m�����U�G�UnJ/^C�ۙ۝�3�ˮ7nܦ�mƸ*��`�._E�r=={��Ѱ�sg>2�v�I��s����u���q>y�[���{��u��1���A����s;��Z��DkH���i�B�N�x�;�u�<%�$i5��;"��z_��>t�#�*q\E��,�����d
`&;$;�����`�/�΃���� u˺b�<�Sx�M<���_`��<�ze\�;�����{�X4e�sΞ�Q
=^oL!��^���7�K�(��r�(u�-?7����Ow��Bv��� �-��y���w��ҷ#<=)��d𻆡���xe�S�,��&བྷ�!�K�re0�������xxsv<7�de@Tq����Āji1��!��o��+�����X"uѫfݙwh�Riun�����/=8ԣy���t���R�)��=;���8!��y�2a�q ^�U�gU���D$�r��_K�+����mz}��g���/�㊟��*�jO�n�l����n�V#|]5z��vO��� ^�O�ŀ�8��k�K�9k��r
e�5�C�ֽʭך=D 9�;�/���!� �	��pLزc篬Э��Iz�72~f#��e�yY�e���W���#<�u���ζ;����o�?|��7��/ҧA�tw_#ԏ��T�+<2��u���ǅ:��g(NL�������B^$�xa�l��-*��£k�8/G��f��J����K�UJ�ex��y��u[�%��V��35m\���^�-��:�3�IKuG���Y�M?�3�Cޭ� �vt�3z7漲�Z�����~�)��i�B���՜y~�sY]�[�m������q�M�WX���v�3�E~}r��/��A&a�ִ��6�kd3`."P�aS2Ƚ��#Ӻ�a!��SL�j��38v� jeu�+r}$1kKd�JCM��*���hOT�� X0Xt���l���fb���zJ 
h��
�k=	>5�B	�d	c@�Z�@�[��n�3r�؟3�X�(l�U3<��q
a�/��^�]uyLP�|�U>Og&��7S�_��,2&�UE��綳�:�C��^��5a��}\�\��tm�~g��sx��v&{g�p����.!7sߟ�S� �]�Q�3�D���� ����^�6���Gt[{d=�80���!��k?�<�ޑ#�U& �W���0v3u[��,*m( 7\?���<�O\I�O�}>��Q@̵DX�c�M�`k�]Q�����t�6�Xe�Բ7���p��N�}�G�/����������ʂ@�a=4B2b"�R2G2��F���a����3����NY��U��a�-~ro��{�[q�o		��Gd>;0�f�:�7n:AeG+)��({�ػ�cn�/%�J��}<\]�*�
�y�ʝa��*J��|Y�%��)Y�p�V�;f��b�1L5D1�U�[�����m�-d�[�f�w�y�~�M���Y�����vU|���1�Yr��X�����WD/�\G/x�|5��[{�FA4�z����,�Ncχ����_����i���aE�_~w;��N�> r7�_��僦��Le6dR������{ �%�ң��9��q�ޚf���{��}8ŭܠ�0q�<��lsH���;2��`��Un�1�[=��p£�F���ډ^�q|��Ks�^�9�
��<���|`]��[�<y�S�;5��mJ��ۭ:�I@x�Ű^��OEC�cׇtD���l��k˿yqZϡ�=�Λ�Z���3{��=4����;�������C�I1�+�&*&{�J�o���6{J��S��{CE�^��^�/V��omq��m�r_�W!
�_��\e:j鋇|���N����&�"��<����Ã"���h��K����ly@���!�9C�6��f�GKT���ʟ�o����F�U��E1�~6`����W�Y���>��	���	���>^Xrc5�Ƽ/��V$���a�ųS�1�4l|>�S_�Y� !O�h���L�T�<�����@{7�G��y45�M��N��#�Z���L��~��R�!�O��V1�"��i�{���핚�&�'x�{�䨙��U�s�����q�g]�H�M5�U���76��i6�C���w�B'1��9	���gÝ7*��5���ݘ��6	8;b�SwO:��!���ǩ_]\��gw��7��j��{���̒��s��7u����)����F�hI�d	���o���+W��35�����@�3��3��TS#I�>���{���Z�	Lc�s�7Lj�K�-�(KSe�~��H7Н�ڀs6��r�E��LkP��-N����.�iȑ�u��!�>�C�*=Ds(p�r�D�am������C����⠱�.�-\Ol�ٖ��Q�K =�g8|�P`��΃�\<'T&}<��3O%B��c=�Q,a�E�B�� Rۢ�6����w1|;�,��*I�0���G?��sL��S"Y�s�o}X&|+�dGK$�y�y�/yTS�z�Z썚��@����D���D��j���'��|������oLUɡ�ϩ�G�����v��G�m����Lx?�U�r��5��r�^����O��z�3]d"�����Л���V��,h;ǞƼ���á�f�>�∊��wJ��G3�x�
C�q �Yϒ��rf_U����%��I7>/�����l�G���`��bP�sJ�Y�| C@B�زO��o�skו�|Ճ�@��H"[X�Vʴ���7X��g���|^�x��}���ԧ��E� ���:�/�s{�o9L]6���/y/wc�Rd����Ԇ���� ����j��L�f�Ғ$�Ǘ6$#��ܼ�*m.w+�ި.m��e:��ͅ�ۦ���{|�+�}�'��'�MM4�M4M4 �|����=���?g(��o��W����
b��!@��na����zhR�ޞ�zk�j5��1�I�/!�fN0-C��Y���c�:���T=��a�y��L����/Kk�p�.�{�י����H�������,�OE���馞�\?����K�T��6S>N��wG8@zXauJM��^��2�=�9H�F8V.�{�w��e|��$������x���[�v�o�.:X*�O��~�N�<��f���y��$J�M���"��:�n��!V'@{9���8�f
F5D����Tk"�y�oJ������Q�h����]�6��@�=|�yáQ���{^q<y�t���E���6��^�?�;�r!���gDKt��a���)fc����~�p���.�c�$}��A~�s�;�����*��s7�^�v��W��7lc�-���~��D�y4��(�>�;������u�x�~��R����"�|�*E79��ޔ�P�Ӽ�g����7�:��Ha �ം /����U�L0e����SS�C���&gm��6��g�7�$u+��������D��uu[�nY���[�B�mں3���I\�q�/ޒ��Q��:��6��z{7�s �YT^ؖ�HFa����vh�T]kIV�������kOG��8�j�)%{Pec�m�鷭�hT��ۣ�O��^V5�뼆�v��r�i��m�wF�j�ww埱]��r��$U׭�-\5�����e�
�82����9���|��[򻛖o�f[����zb/���z�*Ԧ�('����b�L�;��e�vH�Ҝ����
�[J�,t�;#��嵞�z���VV>�D�t�sp�CQG���0�ڹ��4��L�����2m�웛�Ks,��j���c<q�(�7��Nme"�C�А��AZ��)��RĄ5�\ֵP��-q����bu��iQʩ�����o��*'�=�4�G+���9øM��Yw��+/S�lK��WV��-�8\4��;����w�-��GKrKZ�6�՜ݤLN���j��Z�i��A����fŋm�-L<]�XWX��#y�"J�V`��{]�I`�#�Y�u,{�f������'�Z�M�lf��uH:����kE��x#��.�Ǽl���.ՓG�^b4���b�
��nX[�W h���wp��y+nM�qJ邴�+�L�8�.���D6��n� (���BB��U ��&���{�B�A��mZL�Y��x�-ɍ>�՗�w�u�B��5�|���W���������8v�S��Cj�t�9��Q�8S��G/�+�Ȍ�]e5d]b�Ө����³�i`C�e�k�5}��a�ҕ�25��D�e��CM(����=^���W��/�n'U��+Zje�������-����}��5�ݪRt/o0!onE0�H�u_f��
x-^�fW#��L��L
�V�W��7b��-�-����k_e®^m��RJU���7��.Ak��oA.c�h��m�}����5��3jf��9b��trt-���V���3yօ�Ү:�u�Z�v�t_.�,ݑ��p�X"�!'.���x��`v���Þ��[US�T/�m	����*��m����"Z�D�ʬ�uNk��΍���8z9ڧ�����#��U�>\��A�Ӗs�.��{m.b��G((mtb���&�ǲ�Rj�4M�����G��fv}��l���.*I�܏b�[�
t�|����ݖ.��W��A@����&�rvN��̲���u�.��+�soL�s�,�G�j�,����J�|z姉C�e���lY{�(b�����<��6���f��<wrn�Ǡ��I�����T)�K����}���:�ٺ�2EEQB�@�1�1�"#Mـ�T�*D���t[M)%�X�����ں������������yٱ!���Q��ut���x���Ǯ<x��nݸ�q�$��X�c�4�_}�JBf��o��z����ߍǏ<v������$@�$�h���FB24㏎8��Ǐ<x�����޺�F�i,��v�z�3H��) ٤�|m�q�׏<x��G���Ih�T�1E�F�� A$�uҹt���iSQ2�zs��+%�M`�( Ğu�4Q�b61�R	����b4E�$�Q�cjH�[��s\��b4h�w�`�F$�h���\�U���Eb�.]}v�4QD	�DX� o��޻�������ǯ��W�K�M����)�N5o��{W���>UҧQ}�����k�-3����.�Q��o;'[Yu����ze��9�.�!�uv���$� ��f MM]�E6�H�N��,R�@*!�Ҥɀ�.]�E֥�YuwZ�^�:�v�)4�BH,���@H*SM*�*2"����5�z�������f�ww�
؄L��ZClY
ZCe�Q8A���?,�B.��_�WǞ�V2� q��P�~�b�O��ЇmXm���i�&R��tFW����������Y��{l��Xb��כ���`ǚ��3��Gn��c5�_	��Ϗ,|��C�*P~ "�`�/�u�>?}�U��4�g�sW�+g2��~��L�8_���r��l�"^#3Č�4*7���=5�7�㔈:�x�z��h�HB'h���Љ�b���PZm�<0y��#ȉ�`��Fvg�TkqMl�Ƽ�Lԯr1M}�)Ŏ�A�W�d�{)�lؖ��ΞG=;׬�s���SS)�+��k�XR]r^�T\W�O��ƞt��%�kY�z:�\=_�c��r�&
����K�pP	��Ƽ��Mm�~��K �z;\�+U
Fd��Qz1�I�m��"�j��i�i�O�짡��`y����v0�$cXȄ��~~�N���斅��7��k�@ͤ-d����m�����Hp-�$���e5�ozO��ʲ�]7�<���ٺ����Ø�T��a�/TBޫy;���7=+��q�����Pn	n��v1�[e$�ٓX��,x-Υ�"�g��dYwXn����4���}8wCH>�Un.�ܝׇ�d����};h@)��E ��	Zi�FDDX�RA@u����'~]w{��[>��h�W�W�d�#�϶o��-���cL:O� D���h�k3h�fI��Ox�7/Q&�Ӆ�z�߸�2�9?��}����\� u;d;0|�ؐ�|�6Z,�������K�u�3Gfg8���`��u��^�PX��Q~qAO����}z4��vz����n�1����Rf|{���?��g8�8��&k���Ҭ������{<�F�a����󿫾Ծ�+��Ѕ�4�O�X�aV`J�3��ҵ�r^�_	�[��Af��(`���Ԟ��z �3��=�|̄=�@|O"�/e]�zT;l�X݋|��j��f��K4��@nZ]z�+�Y�G7�ncz<�^r5�׸E0i����FO�]���Fd@���k]��13u��P�.0����x�c\ŕ�/]%��p_��-����x���v��]����-��M<�,���@!��0�tE���<7c�i&pΪ[�	�[���/h��%��A���ݽ5��N��nA/A,��yO�7O�����/'Ȇz y��m�3wA�]cN��k0��"��Kus��!�}}�宧re(Ԉ��ZMZT�C����k���VX�Ȍ	��{��U�rO���#"�uT�C�Ub��b"���ɸ�#�w��&S�z�s/{�ek~��Y��P>�iA)���hQ)��R,@dREdE	�yߝϕY����k.�5+��)����{��4�\�h\�[V�����kj�8��NǍ�p�b�+��r{b����ŴXPZD8�yOl�d�w�_�߀��o�%qݎ�;rІ�/dO*]�8�P0�~���!��;���y�F�4��<u^��R��AibK�e7�j
J�w�ɼz��cBz��1^�C�-�Y��֤�#+��-k�<j`��au��#כ2���b�є!M�Hʫ����s�sBl��W���s,�;�
d!�6���_Io;Hފ.��T�t��cڜ���-UԦ�]^�Uw)�.����4s�;����r#�k�6��T;)C��񞇧�6��PX�l$��7�ּ7E=�bX���!����x���ig��������Z��#���͋�1��\��a���u�R����+ߏ�{�����_���X+��?+G?0��g�� �OܽTu,h;͛��
����_���Wlz����_�xs��x/E:�&�#�P/��/��߉9؎$3vBLui�k����\�b���Z�04���p;+�q�V��ۯ�{���}��i;��7Z�y�(h�S&'&)�9�MVD˭�+nk�O7.��Q3�Ѯ̓��)F��N�����:�$L����J�)�/ƚZi���E�i$IBDCU�2�w��y���z�\�l�^�gӯ����j9P(��	Z9�x|�����,�w�n
mݹ��3s�8f�+'�����l��#�������Ű]�C��|Z�&sP��3n�3� �3v�F��
����e�d��m�h���8��i^��k�3������o�e�8��yj��O��_|Q���`�S�2~���ovK���R�+h��l:�����5&�4%�..�7��X}?"~!�����z9�����n�&��ٳ��΂R���x��P|ش��λ�S�Xqmâ�"���Fb���;������>�"U�҃&X��~�V,/Lf�[ռs�`����lQ5��y�yT�h,a(D�#�Z�l؂�W�D�=�����T�U(�|j�t�ג&]$�����R�x��dF�k��1���l�!�>��K�DIu`�ƒ4�ٖ:qc������t�0mx�,Q��]�^i��5�ЮD�rH��u�s���J�r�b����c��;��2VMt��b��Ne+��Zn�6u�6�c�����?h�X��PtJ����Ϫ�<���׉t���=a��Õ���J��ȟ�������Y�;gER�^�� ��n��9�̨����vT��=Y�#���*������zy�e)��8��_a�W��� �� �i�P)��@��	��m���Դ����[P�=�ɿ�P)��T�6����!��YE������s���jΔF���;��cD[AG�"mLpm�{鶢���2���ի�S�DJ����oW7C�^�뤚7-瑴vk<���p�h�'ָr9�̵�e1�z/��V��-��4*�����	�=Λ�xTwy�����`�;�}�#�;*Jٳ
�;�dJs@L	n�F�&���)�Z���*=��Fk�B� A�Vf���r���������|�dꞥ��}jE*~�a��Yc��Uz�O�G�f �X�A�{�)�*��k�'mB��>��D�_��>2/B"|r������u�.�Gx��_%M�]������u�|n����+9���@3����ֲ�?}_���}~��ͧ�Q�j��'hӚ�
u�ŧxˑ&\�Y]��`.6����-i̦{��͙�76{;�b 0��=fК͒^�TB&a������6�kd3>e��}�*fYw�fk�Fr���㩸晫��HY��q�/�Zҹ ��
2�%�{�[:~iw*/���)}N��z^�H�4�m�uz,�w<fR�U�H�ON��.��]+��m�X��\�-P"�`���3f%Y�,E��3�O�$H5:~c��lmyz�Iޤ}{��U���fa�e�n��+C$�+�=���ʳl����*f*�͞nf����>��m�D)��V�h
i�Dd@ $I9���V5���O,>��v����:[走)�Z5����]X9�b!s�جN�~e�ހ	p̼�@ɱ�&9�'�M{�����4��l4�S5$�I���3�>�*�,)��[t�C�S>�0��^Pdd:��q����=�E7s��!&7�]�h��n����y�	�%�:�m��E�.�od��L����˲9�6b|wވy�o�n�n��;w�y����dY�b����\��=]A ��N�o$nG�=�!�~s�W3ΫX۫���ˇCF��dI��f~��Y�x�yl����ٮv`���z�=����X��2*Z����@��2OYP��@���I�U��xj����-`�,w��桄��&��Mn��'n���	��w6L@��Qt��A�h�}�QaV�y��*�����p��U;Y��b��T����|n�^�ɋu�*F�����.4���OZ�tZ5��s�^1������NF��ڝn^{�:Dy���_Y�D���q{�V6��ŗ���~�@�r��R�w�(}^l��b�޹�ۋq��|��4�@������ۋLp��f�	_�'>�J���N�/k4m���J&lڷ���*�h�L�6�<6�=�گ���RC5��zf�ɞ��s[ǪB"��M(�4Њ�M�	"(SM ��(� 	��s�;�~jW�g<�<"#u
���s�8�����4���^�9���灠�x��0���|�e
�
����q�vL׮���EѢމ/\a��"����E[G8�r�<��A@�WAl�g^_���}����N^"�;>� f-��-���E��Cb���k�<7K+����J\ԡ��g��W8��6��z������\�չ�a,��F|g��B�/H>�e�[񮔒8G��8յ�� !N��?!�>�y��X�>�4yi�cݰC*ll�,�7xS\Rds�e�Kײ���͛`��{&*ll_�����q��^�d��>��(��S"�n�7�T���и��żo�It��
<�c_�������>vg�B�[cޫ��:����"�����2����D��OD�V
��5%P�ȫ}jgO-N�$8��l!(�\��T�r�̱ޔ�<�f/�E{�6�@%�/Ҝ�QLk�L]z��1o�v�Ù�1�+R�E!��J�G0,�C#�_Iw�y.�r�\�oD�FAƝ�i*�,����j�[��'kΘ�7���xu,"I�4F��F/���4�C�nZ�9|�ҵ����Bo%�H���
v�M�����S�{gSZ�ͣ[��s�$����e�W׸�NV����\u̸}�������~ֳ��>�CQ�i�)��E��IJi�$�AII[�>o4.C��c|�k�w��C���!6И	��< ��&�L�=q�O�+K3�7���\V;��i��y��R����Z�[?��!|p��韚~_5�w-�]�K��Qab�w<!���s�~F��Dst ��X�ߞ��v�xG7����:�t=	�lS]�J��E�+�5����r�Q�»��~�)>Kج�j eΰ�a��3�p }���9��C.�6�j��t�����ǞEdSkꑭ��:^��~.�S��%WS�|Eִ��xo�Hw,��C�~.�T���l�_D�[܋�L�=_�V�Y��ln1��c�Z<sGi�K^��FT�L��qƃL�<7�����K��I�/��ˆPi�}V�w`�HptCJf��,wr\_:�Z�Z�<�5�c�?�g�k���A��Yk�߲|⮍xL���	�����k�ٳ�/ݭ�,w �&zH�i���y薠�)��>!a[�����OL�i�s�ֽ��}�gU5M����Ɗ�`Z���Y���|�д
�
�DM��	i�X�<_��ܷ5��orAG�L��.��ձډ��xz.��,��5������Z:���N�=b����ݾ�4�fe���e��h���gD��K�B6�v���7���D���Ӻ�d;�a�=��w�Y����]S���=W�Gl�TYv�b��:����� ��ii���iPi������$��ϛ��|�o����v_��;����w�-�׌�����f�k^" 3��מ}��0��s�����S/f#T5 �%=x$gXW����{Ǭx/V�͵=�P�b������-	X"Xq����V*�>���EӤ���m�R�I��څ��tv:qN*�P�����ѐ�=>.x���L&YB���LBb^�f�wX
�M�x܇u�f�ce��f3(�eîN�2�fH8�ކ�������KP��L?T��p�^�;ך����E}�~�Lj9/���f�j�$�l!�"�.�a�K��y����͌a(�y�Bm������ݍ��%MVv.������n���-?,�y����n��M��`9��҆8p\
g��r9�K/�326����G$��.އ�g�_�Ù\�B̄������ �;�׻������<yc�l]0Rr&z_sp�V]r����E���B:���ڿH.�x�إ>�S#+b���-��Ԡ��ª��f��n���^!��pu���킟%���	M��0k�+}��Ǥ��5�)xA--$.cv8�q|Oo��B7��z\2H�ki��t^�}�j�FH���u�p��/�[3��f�U��mQ�W�d*؋η�^���B?͝�Vg:�i�,�����ֺw�sэ�BP�B���KZ��W�g's'�#�7*��ez����T��)��1lZ+q'cR-ذ�lW��:��k^��\��[�7�����~�%!M)QIH�H�M4*� �Y P�^�C��-�B��^�1n�LZ���v}#��![��`&J�O�c�3WB�nR�?���sݹhU�\����<a�@8;�n��l�;"]���o���:�ZI��)��zeSg?s�jL�CvIr� ��	�i/�i�m��s8j٠Ǆ�n*���oJW��3���0A�9�{�.=3Q>�P�8���Œ�!��"�i�8�t����{e�GriN��sȇ�zaQp;������3���ģ8���������w�}�(�Z}*:j�w�~�y���.,��4X�>Tl��Ӟ�,s{��˹*��Y�)&���Z�n�+Z��!�|��a��
Rk�.asȼ�p�Yk~�q7�ͨ�z7ϐ�*�s]�5αj��I�'�%�7���8;��?|�� k��W]2a�ʎ���cm|�1���t�����f�Hd�hK�
�|��>��./m
���T��z ��=
��L/2�	��)���nZ��O��t�<��Y����򨜭�j���6su
��\�T�?���-�n���:���ک��u�pJӶ-��B��HgmLv�q��؋/sB���"�h3B���2
���et�56�&IO�-���2x�����cc�<�JEB���%��
�`���/��Czk&��tZ�J�ܬ���uT�K����$�!����T��*�=7�N����Aǝ|J˥��� �h_
M���W��KDL�t�l��v��4�1��J�p�����{\�j���ح�w���Ӭy����u�3#:w�B���+��P���1�_J�R��ڝF����NX��%䡒2���vc�o�0¼5;Gr<�T']U���M�6�15{m���_�uD2�]����T��ꉙ�ϧ�Ɗ%:���j�m0��5+J���5��oI��N��1�x���R��ͺ����Sؖv�C����aȚV�܂�)�殩��|1Lz�Օ�LAK�a�Vd�ᗻ��X"�lۢ�A�5�+S��4U�2�LR�N�#�C�y�952�Q�&��"Vk�m=�Gg�1l��K�ñZ����Isuo�"#�KH��WA9�A����s;�ָ�UA��XI����렵�ơ���s7�t��۩����ib&��:�;y���̳��|,V�{5����-IJ꼙Z�7n���}I�+W�5)ٜ��t�֢f����+��N��a��:1X�`�>�l�`i\4�2���P �Z!O��2l��N���Ӣ����{�A�o���?�k�?������I��2�8��������+��>�y��K�)R�-�]�'a��΋,��j�b�[ׄ.g��w�a��*�Q���]i`�ά����Q�s�s(�ך���K���0l�v�g�iW{7�*2�]�}������E�E�
Cz	[�ĳ;�3q*#z���ϟ=$f���^��[�;ֽ��|��5�:��0"���N�#qo�A�d����v�f��vX��Ȼ�mL�},<�:a�#Mtٗ�+�~�3��:<�Bk���(�Uu��0��޷�3+�����e9����Y�do����t��x6��n@���P�ˡ��s�yu�y�9���d���4;����ڇ+(pt������_$�p:͜0�2���b^��9ӥ�GV�g�}3v��[)�c��L]�W���M�y��Luy��e���7�Q�_ ue���.Ʃ�?��Tͣt =���oV&�ոTӗ���V�f��L����������2����z��A���YLT���kLp�R��1c�M0�c}b�mRu6�f���Ff�-��x��n�r�Bu}8*�	�(�Od�P���6�s���&O�xDp��=�N=�*#Rp��"��y���+w5�(̕U�S����>�#��1���Ƒ#�,i��$�ȝ�Q$#덽q�<x��Ǐ^�c#$��2#�Z��`'.�l���dI�Ԓ8��q�׏<x���{��z�0�z�0��(�Fآ�	1`���lq�x��Ǐ<x����p�0�26�(э�z����#ޛW#V4�����N>8�ǎ޼x��Ǐ^�N��D��X��nQ�bKE��sAb#lAQ�67*��W�4hЁ�'ź捂w\�!�̮mFKEI�,�!�aF��Q��1E�:X��|�Ta+F�9����`,k�\�+�WMcO��+�*(��U�J��ci�� �h4QF��(�cF��II����r�����7+ȋ�)���uef�k�&*��[���N��9h�q�z�:�FN<�6ɯu�?=�K0��v���{�W��I�4��J�DX�@�DBET�Tb�Q�5�w��ϯ�e��E�ii/a�=K���2'���xU_I熯Y�E���0òZ�g{��
ޔ���fgP�c����c��w�2u=K�u]]�a�a��.Ǹ�,*�O1�N#emz�?���"t��������%�`ǥ��@������������7�N�d�R��v�gҩ�7K,�Z]gA/mr���y�j%��������,xk� ao�W�蟪����pǹ�"3=��o�+��0�%}�S,��p=n��,�49���,ZC9�<�����io�Ձ�*�`�o��X�^ИfE�vk�վ���LIza۱P�0����ŕ�3]#�^:�������)��lh���Cs�B{ap��`�d$*�E��;�w��>�A���Y�eO)�R�n�b�@/結�ă������@O�;�f�a�_yC��:7 �܇,�jf���m9���?kz��,�Ju���o�Vhdv35B����8�軝�%��@�йH��#3��ý��Ѓ޾R�fP4L�p��dP��j�_�H��c��A�V~��?�U>t��7t��{K����i�ͱ�+��+{�5�p]
u�Z��l�
Ùd���Ђ��Ʒ�����x�N��/��@�����ֵf�ܕ/T$�+e����
)��腒rW�g9=�j�5���� ��*+$�Cv�n�mM���ݻmsj��EE$I�}���{=�>�ל�v�cAa�I�*;@�վoV��)YG�$y�����p��pk\�Nr+q��5��
>3�['�y��0F���P���`������W���������^����m�������Ƈ�W �3��(����=�TU���#I�xLt�q����J+u�Oy�5����y�/D�!�1��B����E�S�\�1z�~�բ�Ӗ�ltX���i��w��i����e�0l��F���q���C�"��XDF��C��9�)�a2�9��~d���}�P9�!����S��O����/ק��Qٰ���wY��{��lw܆%ʶ�F���x���9��;�dB=Æ3�k�X�ş��i]�|�Y1��x1��S"[���gr��`�%�^�(jdf�0�`0b9�6M	h;,��j�fq��`�C���Wm�����o����5P����kH��A���\�����WO�x�����h~��r���{C-�+e���Ӽ�7+z�f²�(��ڻ�ڀ+��	���v�r��s�fc<a�A�����Pp�$�5(��!��
/��}�J�x�c*���YW{��'['��V3��2]�O�Af�n�
n�se ����]��o\�rj��=9�yUʒkU����M�CPF4��#M*@�Ʋ~���K,N��\ڒ�ޜ�Q�]|�6�Xen��L�� h�M���
/^�S��u3��UM��K�%����C(����R�7s%���@��A}�<��e~va���Om�����hՀ�߉6��vL����z7�;�nI�3K��4�3���8wk�hV�l�R=7��*�-3(S����H������{F�׮���E�����}�����|ݎ�.*q�j�r��͜O�L�:E;Ň���u� �_Fφ=��ru�5;�:��A��t[3r��?�!)�� ɏ�D�(�0��{�%�=b�K�P�v\H9wٷ�ѩ
L��Q�eP"X\��@Y�q�lA��I��4��*k��8xU�y]�>�X˕��b¾R�%��Bx�9�W��Ra��0H��t��L����Y������/u�ч;�sR��[={K��v<k����y�1��F���ܜ��x�gy#N}��<7L��P���q��޺�-���Q��������#��q^A@�{EI���ʬ�
�9�f������Qx�s���i�YC��1�O��敼�6��0�w@~{�1J6 �=��۪�|�.��:��ֶ���v�o.��oQ��ue_��kA��&�ŗ��S��[���4-�m~(��]�rXz@��h����M���3�O��})yΊ�fb�*�)�2J���¦:�2�+s^��\��Ue���]{2���Ѹ�B~�J�������i �� �"��H�$ ������M�|������C.zv%��ꡗy��6�`Q��Á@����$�~q�5QD{�TK9-�|w3}�����F��P�M_P�C���͘����~���b�=^W07[^�y&)Uڍ�c��������`�a��j �5 h������>�ӈ��?Z�=>��,�!�P�c�Z����?���8H/�`�xWŖ/�c懲Qѓ�of�<㜍O��$�x������T°����W��<�$�OC���<B��	���jgyw�z��#S���b^�������a��}��������{�E�!p[���3˶�����q�a�&�7`f�)�=��{����K���H���Z��w���ߺC5]Sv�$�K/ڨ"���߃b���hObn=�ZB.(nG-^K��`6�~ɦW��t<��,u.��mg/�3�	f��;�S�.4.m�.��P��n@�=/�ۻ׳q�X�/��ak:�V�}uꗇ���h�a�����Y񖰼oA�����|S���EL��{�e]���Q^g:ٜ��k�}e׽e>��'��c�X,���P�wRxt�W���*΅ː��R!�T��y����J�N�a���0R�t2�Q��K�&�dt�^���,I���pK��L���݉�������՛�Wjm7n��۶��2*������95�N��st[��{�l� @aLv�ۻ�/���}`0fs�L$}��ŝ���������j-�#K�<\R��)���.���Ǧ��8މm:N6+�ߧ��&���X��m6L�ҩ2����ZEk�ރ�_�|��WjDc}|�d)�sG:���e����^��!�˨k�6��{b�Y�x�ع�i؞sqfNIx��QVke�7��������!����kBrsׄ�n�fD��z�xW�7�b��/eA�9�B��,l�]�]ӭc��d|94��_�x�#����(6<w�@K��#�_O|{g`͎ð*d׀����3��k��,{mn�=Cؚ!:�p8�C֎���/F�˷�]��j������M��|��~����p���ڬ}���Vn|��lzx���w0B���dsL��l�f{-k�k������0N�u����xu�n�Ǿ0'+�z�=�x�*z~\D�a|M����k���7cv�ΰ��ޙr��a��зf{��L/z$�{�;v={�/4��)��:y᪅��i��uL�P֬��Տ�+�*r������&*����s6Vk���vP�Np�.��ؓ7n�*�#
��6kޅC+&^Al��v�7I_s}XYW}�ҩ��B�ZL�>~���յ��s�m9�UG���v��"�v똛�m͵"�"� H���\޹w��3��xü�����D�}��yOl+����3qM�#��8!�f���\�{���o��L����-��P&Ae�ۤ�%�ޚژ���-^�h%���֙�0�z��ҵ�x�=\w�0m�O|4}���@K瞽0|�.����k�/H��B�4^���H��&�!jb^in�Ym�~���[/��ʬ��8��^͛o	��P�E0>��"����h>V>���b�7�wie�n�������g�&K�K��m
�;���L�+3�_(jzl��TɾJ���҄4x���I�Ȏl��P��LW��B�2o����Y������[�t.aLFz0�C��8����Y�@͙E�{�%�}O-���]E��g8Y�S�Vkq�O62�p���~��" \�����a�t}o�|�r�]��vw����NM5 ٥�j��������-A�6�{jY�7�ڐQ�D �И�������%&�UV����{���t�=c� � �⠱��a��'�<v��4z}�t��#�[L0x.�Kk�M/����4��[��_U�o����,�GF=y3�v��Q`�-`u���6�_���r����T
*��9�x���I`��2�X<�Sƒ}����\6&*�e`��72�ȁ=��f����!�؁-��xʗZ[[�T$a��3n���_3�J�F�x}�� }��`����usv�k��ѯ�}�~F��.����u���Q�I#w�E��ͽ��.�:�^uE7=0E��v��T��z�X��ù譐��K����5�Ha�3����#�����Y�f�~S�Й�f��L;�,~A/r�)@52���'�6~��/���w�����p`�S�0�\�óe�ҊcB5P�g�����u�sg�L�2�v�[[�x��k����m8f�fr]C�b£ՈK��Ǘ����U��ln}���>��^�9&�wrtg8ː�bʃ���2��1�{�'�,��V$�fU]�B�끱��<��֛��������@��z�-�bQ��p���B3����6�(�Ox���g���}T[+�grTx�}ZS ������J�˰ygz�:L�(S��¼>g�Oʼ��}���>X�zd�=���T}�H�{ǜ�x�z$2�����Sy��f��Ƕu#�S�W^�m"7����4�#�l�p��[`j�Qp)��K��."Q�A��$������������[>�Uv��}�ʶ���]}G8��� D_� '5�����N(b�d^�SL�WZT��/��E�U����v��lO�C�ܹ�� �r�D�u�C7��Y�����l��M�.J�j��[�ve�l��Ax�_����h��y�?�ʐ�K����uԆ��b���K��`���:�%��^��Mb����*[-��=���3.��������SEH�MH��RIB#		/��;U�'�9���C�ְ��er����A�d����t#��YC�8��1�.��E�E��6��4O����dS*Ml�p:ޡ��y� ���JD�~�@Ⱥ�	�U�b�a�r�v�o8-�^�f_Bb�sȢ��Ú���#��
=���6��{.�+jj�95�5B�څ��yL�M�&0��1i����O�y�m�a#���D��3R���۞O/��E���h!��먦�Q%������ǡ��	�9O�����#���h��C�@��w[AM�Y�#�7̵�C9nS�:ꁦ�n��վ^�*鼘^uzx�j}����CҺ[w�����Lk<
�!;��.� B7�ٓ����F��<�k�Ѭ��m�$�|�p�M�z˶�Wv�}��^-(uc�_�� �+h�����Bs;c"�%�>Y��T�j�Ʒ8Gi�t���4¸��3�4{A��-^�V)��8>@��.R���>����3"+��2ۨt�犲��G<oh��<gy�<�`k�겺l'�A�ִR��)�ư:jn[�0��ݬ��}2�n�<GH� D�5��Y��{�Ar�gf��/9T[mfG�It��A��l�k��8_�볦5�g�"ju�j�������&ͮ+�#:��<�V����L����!gV����W���vv�[�FI��ƫ��׿����k�o�cdÈzk5�����z�wQ��� �'
e�ΘG>��y��0��>��K�GoriA�-�	��$��<�O藖�n�(��9�Wk�`3�>���*e�r�A�Z�Z�\��y���qSl
z��zaP�=@\�.t������s���Uh\Р�!MJ�T�k��&�8�y�Y�;����8��y�;s�Ol�� ��	�*'��f`��<D3?<D4^�	��*�*�Yam`��5��y��x�[РȺ	=k&�o\���>U���W������Ys�<_���]x%��؟e[
ڋhUӐ�i趘b�f�Xh4qW#����*���5Ӗ!��H��&�"��y�K�
��_;5ظ��C��}t��of���\�v#�k����(�ؘ�q�6���f:��ӣ�c*#�d�HM�m0V׶C6z��1p�`�����6�3�>Yz�ܪ/����(%_O���ܙ�m�%l8ׁߓ���2�^���hϩ��b�v5h��㱱�{����ꄙ}\W��+1��Q�[,ܝ��F�h;��U�.���Z�3RwF>���ӽ��R�Q}�ǻ�"����i��9Zp�E�!ܿZ�鬫(��dlz�{$��s*G�eQ2�v��٢&������$�m3�2�@���eS�5t{!�N]�+&�����ߗv�v�ɻ8�����P��y���������a{�̲�R�"~�Z�ޞ Ħ�AC�a�Z�^����Y���R����_GVRZ������`�%�J�a �N�{w�������Q^��^����KpVwٟ3��[�o�LE<x�d��k���8��/h�6;������Nq��yٴ�@c��E���\�lu��A�M-��Ncq�6!^�	��L�y�L |��홮�M�ޚ/f�۱��^,z6*z�~�X#*��fs�ug���t4 B��!�=�y{dVK0�z�y��W�%��* ��,l�2�ӓ��???:�{*+έƂ���)Ӎ���	oHA�W~��~�2R,��u�Q�b�~T�w�ٮ�Os���LݐEx�5�K�����E_�B����%���d.��	���V�@���������psj�v����n�j�K�}g��X�/|rz�������Q�,׋L�0C]�:n5���BS]��PL�N�£�(Q�z���̥e�S��O�~qoڕ��_��1ıw��6���m�"u��7��(t�Jo�
�Z#&��������Ց2�rs��۲��VF3R���bgf:r
���u�.
����rY�Hvs�Ë��\;x��AN'	�� k�TV+,�YRPuP:�е�s�����.�F
�\W;=ݏ9�Է)�b��N�ӻ�@~�W���%'_�i
P~��Y6�^>����3q]�!SP��8��Ѳ�N��09]c0N�٭�D��b�9��s�e�١�+{:�F>˗H��<�Sׄ���e�6��X��+E��X�e�9]����r�e�k��j�r���_\M���B�fÚ
��.u&�2X���!�x�'(�Y�+	��9T͘�+F�Y6�<P����Ym|Ai;��b�!��}�>���`n7]T�y����ͫ���ay�5�t�؇�Vo�,G�e����?WG��YXMإ���v��1G|yoc}qS�3h�Z�k��)a�6��PP38H�m�kB\P}��)�L��
ﷁr��6�Nf7���dα;�����-�G��R�:��\⽩؈�{�\�`̳씠U*���M�]�.�!6�g�WkA�}�{I@��Y�J���c��m{���f���՛���WZXZ�)gn䕓���*a�U�}x:eJ!�Vx�RĲ�<�}�hº��=���,��od�ՏcRNcn��4m�b��WF�z�:��{s�Nfl�8>uL�ׇ�8o�И�Ro�R�u�U6�87l�N�����I�nm�1�ʉ�l]o&>=�A�)�NA�hR������՚�X����rS��)]�^S�:]�7��x���B
CH"ˬ���W��D����`�坃*�=7~���7�Vv7�L1��[���|#*k�{R�ZT���m��K�P�cF+Vu���5PF�
�nrN�9��9�ϫh���֮�4sKX�j�.evnI�b)K���T��TM:V�+����0��&��T�3�u&4��i�I�L�d���f�.Yh�!��q���Mj��_%tz:��릂Ǌ��Z�(;F[V��p�5�IW[cnv�R��7*�<�����M%�1P5Q������[�s ��vVK메��5�:Hou,ǵ)��YI�5O���2�.�KCZsC����u�.��]8�gb[5`�Fi�eWd��Mɯ�X�0֒�����K��k�;N+jW_p��f�b����e�[w�w.薆X;+Pze|�t�R�`vZ]�	���m#d�_��8N�=����2�ڡ�SK�T�)������w(���: �w;��jQ�1����kw.1�[6�0��f���ɴ�vPAq
�ݾC����2��iu��A���>9[Wg���3�a��٧���鶚/�it��{q��K��*1���W��ƕ����!s��}Nm`sh%B�G��^d�֒�J�`�*�(��I=�����2�V�O��P�J-�f�&�3�/²�R\�P-�� �wy#@d���ϭ�4Ai(�Im���		DdY��ݻq����Ǐ<z��� B	#��O]�4Z�FѰZI�	��ێ8�Ǐ^<x��ǯ^��/H� y
B� �bѪ���Ʈm;��Q��q�Ǐ^<x��ǯ^�� �?�+%�1V*�4t�n8�=x��Ǐ�z�2��*-%��X���DRT�-]+�\���%bѹnQQ�66�oSmr��F�6
�5��ű%cV+�Z������5;�¢*�Am�V�d�5ʋlO����ݪ劊�F���Z1����%cEEIE#��6�V@$	�M���&5�^]��i�����bQ�������p0���>�ފ�@�Z�V��K[�[o����s�D��sz>Ȍ�'������Y�)<�=�������ʺp�D�b���q!0[��`�
�T�� D,��,�If�.7`�LT�	NE��`���(�c���/_��IILcU!$#��<�H?�;Fn~_�d�]ے�w�K��	�Xr@鷗��vj�$�x�_��%�_���I�ǘ��>�3^eA����5T���ke۬����d��/�~�1afGkH�<���#���t~��Qt��f���^���^�zs'ր�yZ�1�a��7�r��S	W�(>�ap��쾖k��]�i�r��Iz��F/xٝ����������i��!~���s!}�����JpR5x�n���&�
��Px��d��Sz��Z�c
����4��~�=#Xv&�i��+*S��=��`V������q��cv��wZ�,�K�>R��+����*n,G �"g�1%\]���0��#B�Th���Œr�~��б��^��=��>�؎1�	���%`~��3SqmjA��ɀ�� �����?5�<��Y-�n�����dBa��m�[9��uU��\���иB����C�vy�k��,ֵY*��u�l��5�)��.y�K���k�vE3Q�Vs�wi������$@-�$�4��-ĳ{b*�"Y��d��'���O**��p���0��_(<*���E߲�Ͻ�����F/{oi%�\�l�䧺�~r�E{rg�tL���j�{9UN������Ӝ�k6w�.-9*st�����U�X{BN��br�֚x�N�29���=�{9�V��2s�+�~0#�H���ځq}�g�)�o��.®�i�v
yA��|��x��߬y�&g�J&���yl��i�4a����K ��\ߦ=	饨-*h?��!�Qx�G$=7��lc<�(��k�ʤ�cu�32�!Á��8:2"-�2b�݉�m#̸�Mg�LC�q,^�Q�a�F��W�z_no��Ԑ�������r*$�j��ÄE��J�2B��m�lA��,��q��*��]�,N������U{�f�F[�W��4d=��z$�����O0��$T^;rݡ�Z����1
$�$�<�dD�	7�S������uC���j�����~��^��.�}�1�፲b����FmH.�� ���D��9��b���Cp6-� z�V쉐�RWx7q\����L�7��Z��sb9̿���<�G4�v%�͝����^f�پ��Bݚ�a����ׇ!M{S��ؽ^�N�}�ـ���*;���1ŋ��{.r����I|E�o��}�t�0s�!�'��:�Cc��0������a=
 ����"��ڹI�*���Z췲�?�������������n�g��tg��wY�1��uD-��g�}2�m����c���yn���Tǳ5��^���5Va�[k*�켝Y�Mt9%���ޣ:�U[���w�~����o0������V"y2�^��(����ҏ�)�(g�?|r���U
�2b����������7c)ex����~4߈��@x�/�GsY	?ɰ8?�D~�K�_<�������L��e�w�f V\�pl�M0�-����f��n[ƂL��M�~(��?�{p^��O�rƮۃX�_�	�*�]�=}j�{y�*�4x��6}�T sCU��`�|��ť�.��9X=��h�x��kX/̢akס��YuYq�*�M��KǊ�>A�ș��ކk	�l���V�[*�m'�f�b��k�#�p�!{p�{�N2.NG�j)���ۑ��RY$7>>;;�R"dNN����A�ħ��1��{=^��lS�0ƅ��j�U C�>�wi�|j��ŶrOevm�v�P�{
�^��X�.�4���wQ0潰���yO��Y��<+�\w*�?`.��1J���n���Z��ɞ�7�;ʀX�R�TaLv��=C�*i����3	-�Pda���ؤ�]��&�5(.���F64�D������K0�L�Rzk��a���y[�������U��7��τ��F��W=�Ut�½W�s�y{��mҲ:��[�K�o=K~��p{fЊeϑ�v���1�e����}>C���c�V]7�wP`��֞s�sZ���W\y�K�D��B&2�"3�#��b�f���g�wd�~���0#�9�5���;>{MM��]p�i�k ��؆l�4����O<�Qx��y�p9��u�+e
��A���� rc=y�~�S��Èu}M�{َO��9\�/�K�UKK��b-6x�M��_��sP��iQ`|{wO�s̻{��~�,Ȟ�_R�fˁ�F�)��٠��"'����ٶ�װ��&���L�~M&	�k �����@Pm2m�g��d��Dt��ђ�5����t��%�7�i���G1�J�������N�(x,:!MA!���om�Cc�y��H�`P��P$�u)8�zV߇��TQl�H9�����s�`0�<�s8�c���4��0�W��J����xC��S���R^�q��ײ�N8���1b��Ϳ$�h�ëA�5F67�f_�[	�4O�o�=b8�^�)u�PNa���]E{=��~�@�<���~:G�π�,�ZZU����^��+!Eg�hO�HUn���w/����.uuNژ�ҳ��V)����Hؚ~�J�c����I�w��>�3)C����@'���C�L��z�vC�U��'q.�ChZ7��4,�
�3����Xx��]�1D�B2�q_������W�C�����y�N|�΄�R�=�����7]k�p�����iܼ�oh�G6�*��o<7���엑T=���V�	[񂑁�7|g�wƃ>\ټ}�5.!�iA��K7N�� ���g�xx�{�ӷ��\��$!^D׍����Pj�?��3���|�.�W����r��twmU!�ց�P����2& ��~��������tas���3=�!��v��z<r+���З^j/m��d�w����"�d��y�>���=[�[�DB��mui�GQ��i���Ce��v*��J1�Ȏl��D��J�8MaR�����w7\�\��f���x���iE���/��,������,��]?7x�W�r�ɳ��W=��g��%�����J�QaO�\��s	�\?��cX�}a7HW�]�#���(�'s<���-5'����):�7z���XOc��p��� ���͞DKmL��4�K�<�_��.���Fs���}JO���z����)xb�t~l	Ĵ��->2�k(�b�7H\>�GTlM�<'�Z5�4^�B���f �Q�fJ���q�Z_��dg�����QqWO�̣�S{�0e]�e�K�?�p矨LKbl3�ݜ�"N����k �y\W_0ǪA�wf'§�o��V��V�C��~7����F�.��t�]�xP"�=���i�М0�1�0\Q�&}H�o�[r�uù�Fޡ��=;7*	�i{�-�v+�����I�?��"�׷�6G��.�Ҝ�����|+����o0�m.�1Oa�
��8m�B�(��/�4Nb�΀3�Uw�ȭ�m���'b�$;]��,�V.�f�W !��yP(��Mh���ο��DS���M����D���T���<Ar���߉�P���_�hp�:�E~x�_�V�� �������<�Z��f��wf�F�Cb�Um�Ķk���@���� |�Z��P�T1���0��[�.8A�~���UMj:	���K�w�b�8������}�<��A	�>��Zfb�9Oo�]������i��p� �\_:����x��Z�w�� �Y�*��j�e�ٴ�A#��]v�F��=�(�?O�i����b�yG�3�!��@F���M^Y&2����Ԧo�n
�0������o�l��x���_��>�>��ө{IbP��Ǟ5��x#a��E�d!�f��+J6��=����{�����\\:au�4N�u#�;��>��F\F6��z$��)�K[JSS>�솸�^�@0-�)o5�J"�GU��-.��'K�W�K>�;,�ͥUjWXJ4��Lw���M�k�{q�]��4��`���+�2���s�]2U�=ʮyh:�=搶Y䯡�Rۑ�nL��5�c�N`��^����[�r:�1	u-�j�6P�c����.o�]�˔N��	�a�rL�Fob���Q�^K���*�Ժ,�c�hq�l.Qb]��s��':�಼��Al�1����	�L;e�s(z㞜O�S�-#;�iؖ29wJL�U]c �6���z����!�G@q��^9�Z�H�������vLe��Gr��D�sr��_�w;�ߗ|�o�F��(�Ƈ����.��)��|�g@Y���oJN#gs�ycF����<ͬ�mO�'��� ��+��H�䙋�����̊UKTSF���HY���}�뱬�
B�6_q����s~��k��o�A�����t�R���X~�g��j����u3w����V�'e�i�q�<���s_��r��w�� p��ԧ�On2}5�����A���s���W����8ė����8ð��6�Vk1~�jq&��ؚ�~l!�BC�h!Bi0Sע}�\��j�Uv�/`���&&Y�l6��ǽ1��{Xyͺ��bvԢ�m�o�[�D�FgA������)�*)��5� k�����Λ�k9������"�QsJ��1
Ok�r[}A�0�ɳ�숧�����f��3�,����bLW�|O��Q��ARK�_������;���4�����A��W���U]b�C���ܼΑC�wn��t�v�nnEO��s|��9����b����|*�p+�?Xw�2��4�@�Ξz��a}�F�B!���Ea�7M{y����=��U�Du��}�;b�	�d	c@�@iU�ք�q�^�`�+��X���勦M��c�u��$Ew�J5��<�W��ƀZ�R���i��c_T\<�{g� ������p�^�S)�ڏg�������P�r �P��~��㼰
f�žE0���wխ+��Ʀ��]�:o���^� p7��<�1�Ԧ;� �V9�T�p�Zg1mV,}�(X�]n6�������1���<&�y�ʄ�T4���~/,�������od[�m��ͽy�c8��A��E�����;�A+�p��2��K��*o�kW�|7аq��j�p!�*0��K�N��-�C�;��nC�˸�2m���y�L(���ڜ-�%\ᾬ�
�ە�.�⨳y�Z��3cԫX/�������i��?�|@d���y>U,ͬ�V`J��p[���]@?O'�5�es��%�Ts_����v=���#Qz7TFF��M1tM�=�����<ËxavG��׌:�z�9wҸ�uY��殂����b��t�WLjMn�\e��i��|��鴘�J<d7�HY�w���{l���Ŗ%��2�L�V���]�S�ìS{�7čs&Mi܅��U{2J�T�^�X�`F1���!�^:~.ؿ�|߷;:j���M]���Q�]��}������埨FO�}gԘ\0v�dp;n�ށG�v`&�w8ċlf��+��Y�\�T�g�=�\��p�yk�FO�#dg�������E��sɁ�h�)5wy����v�u�ʾ@��"[�Ξ@חxб爌E_,"�����q���e�_y��I�m��߽ݗ�7��~�َ�\L�H<"ۙ���g@�y����n�Ȫ�������ʗ�>ךG��2����������4���MC�.Z�� a^�!'�^q�����1o��*Vc�q5"�����~���Sy���������P�E>���/R~�Z/��c�܎[0J<��9��C�ǔ��������zdB�^���hP��ȉ�	�QD���+4��jgM~5����bA��O�l��h��Z��K�J`��{"YA�=_+��=�q�;q�\c����߿;���++�
V��,/��� g�9P�2!�6e+n�MK�B%lб�ǯ4۬ؿ[����(ϠW��`�{\8��膷�L2}�i��"41]T���~l6��B�'x/����5�����0�f�ۛ����9]�����oP���].��oNÖ�	��)^�G�%�xlH'>�	�X�أ��-�qyw����6�Nٓ���ѐk	)ݏ�"�����,�>\��$�=�ՙ�9���䒟�c1��{���20¾�ܡ��Y��9L"�x�U�=���c��S�nxw�A;y��	��v�u�ub�$�*/�s:r'��8�.+9I�<�������F�#��I�4x��'��T}n�:̃�;U���{���O�%����t%亡0XsH��qqw�Q����U�I�H�-N�脄*)?M��2-���}N5�(�:�����dK)�}�a�J׿�E��q)l<C���m��-o�1tc �`�
�f�Oο5��M$�Ԯt}��7G&��U��<Q��M��_��g����W���e��L|�(��_�G��&��"[�~d�������BB@���ݥW�W��[��D����a�SE�O��w�Ņht�<tY�!����4٧?�w��b~��v~�j��4��%��jv��3�_���nڼL���Nf�>�싓�ߤ�\��������*r���z�r�	�n�a #R����o"��X/X�Ҟ{ʹ�Oo۲������{����f��P�,�_�=��~������P�W��`Z�G(;�H��~�.D�R���y/6&��2ߖޱ�(��i7���9V�h&�n���u��s�[�)efb.���ի=غ�z�v�m�kv���b�ƆvD���誓ZFg)^�}Q���.��R��v.���9�9��HOhY����BS����f�����r��z�Ht��ͽǽT�ɲ��2^��z���:�:����Őا3!"v�}��Et[\��K�,B��=2�&R*����VF�Ւ��8�2�T�L��n���zk�%˪�k4b+)�Zgm6Ѽ����W�t��FB\9�s�u��f��%�b����h��a�*�v�O�����F��_�r
�����%k�s��W|��P�!_vQ��	V5-�o�ݛ�n���p��1�8�o*��l�/]�A�oC����]��.��rǯ���!�kFTo������3U�6f3@��i�Ϋ�79;(�u5-����$�y�5h�dm��{�'QL9����R��D�V�˔�7�6uI峖�B�bK�{WZ^7��^	mm�#}kGYѪҲ2�՘0�#N��֞��`���s�9�T�|�ӓ�RX(M)���)�:[f�C��CX���H��};����~�j��3�;%,=r���wps���/b�8���pa/��[�G�Vz��׳t�1�sq���7!q3}C^�[{C�}{�J�]'A��<�h.O+}G+2���u�^����i=C���G�7�>�Ӓ�u��q�C�[]3�
�+�ެ;����|R�$�[n�ⲄT�x�C5�"3Q�r�E�.�6E��3���m�t��i��s;���N*�8:����u�J��}�Ү� /,����T[Q��3�c�^(��R�Xz�I�=�Ѻܶ�4����-,FI/j�;�ag@�ef��G<Rʧ3���/9�T�lr!6�*�ۼ��U��CZN��_�\�t��^��]�ܪ^�%c�F��f��Ls�;d�=y���"�os컹H�ڧ���0��*�t��6AAuHK8S��C�v�|�.�әݶ&f���N��j��,p�*�3Z�#-Jt�s��34��r��4f�w��Ӄt%�0�V.��9˃d�"ڜ� �wQ��/k������%�Z�#�m��x������CʼDYZ{A�{V�'�V:��R�x/(2���[f8i���I^Le��x��A'@2�����߫E��������b<��'����[Ou��P6W�f�t^v��J"w��\{k>H9WBB�7l'gV�m���M�%��E�wj�t�R	Q��,��k�3١��Ἐ�s{E�-a�jG*_��@$��Z��j�kE[�W*-(�!#PJ��G��v��<v�Ǐ<z��=�I�5$RA�	2mx�
KbѤ���s���8��<z��Ǐ�z�	"H!�Ѷ4jEE�[4@�[m�q�Ǐ^<x��ׯ@�F�ƋcZ-_��z�n8�<z��Ǐ�zX mbأl^�6�����o���kr�Z��b4�F�5�[cm�fܢ�/�QYI�m5&Ŵ��׍kɰQ��IX�|9h�^�r�F��⹍ZMQ���,m%�+c&���U�ة�H��$�=�.�U�������%)�t}��N�ʥ�����+.H0̈́m����7׽��`�7ֲ��^��z�sh��o7��{��i+*J����Z_���|dS�[U�0��".�U(��2V2|�pJk�zPd�u���v��Krf�7���B�zo�a�l�4�žzݙ�L�]��b u�Z�i�Xg��^Zn��oWp�"[S�J@�V*J6���l�����y��B`�g-Lt�r��&�4��J�瞈,��DIuc�����jn7$Od\:��� �65M�{��aFg���5b
Cwz�KxOd!3z�$��O�*��"�].9��Yz|�?.w�|�UZ���I'ã��"9�zaٸ�kT�Hq��K$�Z�>Pq������7>�N���AzSf��`�(�4[7�=��Za��Y���W틮�j���U5�����L��Bf\�fxWc�6��v�\��	���׶v; o�sߣ�	�P���`Kl�7j����'t����Z�Ok�͍/(R�*�z� �|ZD�@o(>_yP�NE;sF�?6ena��nMe!E�9��>1�����/�{��1�]Cl���p��~��So�����cɸ��$�<�Lc\\,.uXfYs���o�f����d8�jS�t�6�0�;G�,O8X�f{�^�_`����@~5V��==j�&�AZ.q��@WU0�Ԭ��}R�[z�w%j6-�SqMۥ[�=�=��s�}&�1��QO�ϟs�}
[*-�4�1}��,6GX��>F�_��P: v�� �K���1�h- k�<c�\s�jwB�V3�m����F�Hlx��Cy��?5������=z8ʇ��wX�fu�Ta��Ѓ?\l8���vr/^?�.�D���Tx ф%;/]�]:~���Z�]z�V<Ul��x��g�F0���h/sq隊enK�~X��i�f�z�)��K`l��`��ٹ:�C���*�Η�a�_|�Wj��i/�W����K�MU��x��5+g��g>5��q<ߕ@�;�E^��q�1P��� `\��IqT�u�0u��gF�~:L������h��Խ���}h"b���c~��+UE�5�8�K���|g:������'������T��p�T�|�M��~�N���BN+Db�c	��Ы��޶��{����oD��M��͞�`ނP�������1�x��y\��^u.R��j8����\�+�P�ْ�Tk;$��#��X�Yvd�V�r|������EgL�xk�8]ޢ����j޽gq`I��k���6G9PsŌ�oW���c�6�O����CW{s�ޭ%��{v��z�F��bi,ȝ[�Ǫ�Ǹ\J\���T��J�z�,|Ws�`�Q�8�S��5��sv�%�U}��˲D��؋�r//7���� ����i�
��J�[���;�����ꃫi��e����T$�s�;k��ؘ�}���W"A����-���2�t�6dO�9h�Jg�f�s�
ͽE���y��$�T ֣N�~M �f~�(��B��l|w�1ߧń�K���rxS��p52K��8�,*�3�sSJ���=������w�4��Uz͋J�콋�|���a7��~jWL$k��̀y��
mr���"Ts	ji�:�;k��9�B�3}��;�	'����j���w>^�e�.K�}ʇ[����-��j����w�wE-+�1�Se�m�ͬ�2/A�ϺC3���0yk�FO�VI�����+��G3Y�7���ˌʣ�w�s����������q��
g��,�E��;!5E,���6mhc������=�Z��j�d`�I�c��^)Ẳ3�`L��� �9
�*��1�(f��r/����Z|~d^�\?�E
�D{�D�zd�1	)�vGS�����y���:#X[�7113zՔ�t
y�L�=ˈUZ��"�q�1�g(u2q���4y��Ӎ{��|�)�PQe�V���+5��3W�[��gf��e��!���ݻ��7�O��]Te�^��}�v#��W��ܴ�{��^�}G�������[��������;5m[���du�}�^�UV��Fjv�=;�=ߗ^y�=7�շ�g<�I��#�?T�f��r�VyCD��������q2�!E�U���	��j ���=!2���'�Ghe�`�֚�����ΧF��n:��xi�������CiW��`�~�.�zqh|ٽ�i��s�n�j�uy�0�C&<�Ņ߄l�={����/FDz$Pq�	�T�I�^{�^�/�^9���+e���b�����c�1v�!���Qz��lhk�)s�B��*P@1�.7�cZ�Nt �A����ِ�#s���%�7�����x�C5cb��l^p`�^}p���nxw��:=����ֻ/��mʀ(,iـ[�=��juYJ_(�}b��ނ�WI��s������=.�%�Q�~T\�����'^�Oߧ߈^:`z�? :a�Z��#��i���x��K so�y�FZ�#7g��;ϖ#�)a�����>�Y7� ���q�5��A/r��v:k�62-!��v��6�1>���<9��]�h����8ňQ���U��lkt[�`81C�a�r��ӯ^I���;'��;t�`38��/��_����G�{������g�^�v%eѐĔ�ejG`͹�֖����Z����\�z�%��*M����Ou���?�^!Ct�R��.���~��?pb�9�b��ndj�v���<�j�G^W�5�q��p�Mo+1���]�n�ȶ{����x�Q'����f`.����W�3he�u;������(m�ޯϴ8x�C�4p�͹��D?�{;�/�飨n-���c��1Y��i�6��E��jA}��lEC�dK=�*�ˎ͋��3l�!�{BM��i�:b�m�\{]u	݂�������ߗ_b���_���wU�����Y��g�HS�$N4~C;�k_�~|���B(�8�7Ú/e�F����.�5`l�y�{�K$�{�_J��9ެ+�z
S�-�	�ȋ��j�cW>p�_�i��pcL5Y�"2�p�`)��Iz ��\��F3^���ջ7���"X\��+ -���
z�SB���l�Cy7��ȍ�/S��SL��N��sS=���A��ˋ�.����X�E����%[	�xwL@/�%�P%�i5��ۑ����Ϻ�+�-YX��˃�#�����k�0ɿ2�!��[�`ԩ'�_�1`��F�'���ay�,���D,gq��>�0@pQ����1��n�Z��ۙO�o��'Ł<�f��q~zsG��'2E��!�`�\1_K������4�=pcS�A����E�]^�Y�ࢯ"	�к;���|D����p�X�u�S�,�ArU]tf�����R�O���Ȧ�͋`H��+3_����39���BG�i�i��h��eO����j��|T�	=�Z-��ZD9#���^93�A:�}��~��'��9Yc��߷5�0��]���u���|w������t�+���6�_�T��H'/��MY�d�ݽ~�~���h�M�L���E�x��Ⅾ�/6)O� *del[��1�0}a ���xv.��t�V�zqw3G���P'�Υ0��-3s�ǣ��g�=+�W�����<�V8X�;�{�Obv��ޖf
Z�~b������"�y8��~�a����ƹ�����y��=4p�0��[�����>-��h0.��ج|~��﹆7�:{�GJ�/�脫����GⲲf^Q[�*jM��}���Z���B6)i���ʿ5F���c�X�&�f[ļsLַs�K��4��c'1	6b��Z˯�x@WHf`P&|D[ql�ߦ��>�������9l��9�����!�V����
�"�i�8�t����؇�p)�Tw��j�������L�Zm������4�p(ֳ��u�ì*r^k 38A@����O����}��6��\�(�j̦ì<¹��D6�ʥ�ZFv�]D��
�x�����)�aB�X�y�;6��}�v`��ɲ���B�2�zn�];�p+<���U;_V�*B���]���fY�V2��������*�wO�y��o7�����єL)�kW0������gX�V̹��ާ})�.���=�@���V�?���Y��c֯��r��JS<�����0�/P씛j����y��d")L���66s͖*8��c��P[FD�Sw;s�tF�APS)8�@��P�ӹ��d��v�B�[B�<±�4X�t�؆R��m��eRc^`�Y*�DS�7u�Z�;�m:q����dA�����b?�]B1���vV6�CW;Q�yc�����Ik���j����&<f}����򴁴�T_�/��*|{6�O�����kmQb|���4g9
(_RaUfW<5z��OeAc^�i�Jxw����6:m���/�q�ł'*�sj����K�sBzA������,�t��J������ӽ;��:�C��hƆ�51YFL����&X0.[�`c)�"�?O	�u-|*���Ts	;S~�u�����;;�kD�3�=/� 0|�gC��������様O����U�f�Ž�X���G'������(O��磍���n�r��cÚ\�s���zo�:aS&�7���<۳\z��`d�\���v��&}\83%�<n�N�4#�s8%Y�eeӤ��Ə:���h��k+��{-n�q�<;�OZ�eK�o�y�!��N"�ɘԛ�c;�)�ѽ=t�>u�����{2�wh��H���F�������|�vps�����Y���C����ү�1�畆��ȧN��5�o��x9e���`(jfL�4I�p��X��?��:4{�G����htt����	_@�E�$�S�d��L�庯TZ�F6z�*�k�n?'*����4���V��X\�yg�s��q��C���6?ie
�H�u�=~
0"��a����Ɓ�|��8�㇯fͿ�h���s�DE�iw����r�b���@��
����yO����wP��g��.�.V/]f[���B�9��ucA��A{�^=z����v�4+��H/mL���S�)F4��'3�5�o�?/�;�پ�H���ϛ�Ǖ�S�:J�w7��L�����[@N��8I����h7B���<��}P������w\��,S�y`x{�W�S�����i���3'q�������h��~Q~LUd���;���9T��9�P��:�u�j�mx��Y��Yږh��#��K�Ϣm	��2%���T8�|ń��{���5�N%2��0�Ʉ1���ФQ����}�!0H�s8ݰL�����P�]�qwZ�d�f�[[��ۼ�g=�t��	Wcs����*�N�C�j':9���j�-�ɂl�3��f��+-�uN��V�fgmA���d�`��|c�1��_�ᛙ�~�UU�MaO��^�#Y�ӫDsi�F�߸�0�j��^;��$�mg���T���J��T��tۼ{����Xt���k�&w�~�O�]ޟr�7�̝�Fͮ���(�8¡z�x����>�
���]�3���&9��s������ߗ�Jc;�-:�����nә����O>0{j~`(������H��;w2|=����wO4�V.g�U����~x*�l>�Ϣ�ύ+Z߳��x�Xh��K�x�qn��15�d���4���xleݒ/����a�O�C�$�1mq�؋���S˗�Hƚ�6��gD@�����`�xi��p/�W]"w׵�,+���LL8���ǡ9]xى��izh��@���pCP�`5��0�~ym��W��2�i;Y�دS3�[c;4�kkӲgM�ᢾ��RLXB˰���o�����'��ԡ9��h��{5�Ds���o#C6�Ί2ϜW�FSս[�z����Xp�H{��f������yS�Du�Spbo���l��a䬙>����W�����G�f�~M*��V��]�m�zQ�u7>쏾��z
�>�Q�PpS��1�Z�rv�0̭%@�'gN
٪��{y��XƪΔ�2����<�םT��+U�����q{���������SL�oQ�`�zy��N<2OE8�v)UЪ
6�����i�����eA���;Vm��A���}�08MBא���{�DIt�)Ķ�����!��=Z���M�-���]V#Ih0�?�}��/�����p?AOH�~ܜПoR���LW1�}J��7Vs�N�&����De���<���kB#��Bm���p �j��{~d^���fתNM�� �5vjѴ^F�zi����@h���i�#�;<x�>\x˷V�ЬƜ|�覊x�XE�&w7���^��P���r�>X�cɤ�YD?�c_r����xL��\C/�����7L��;Cw!ءkZ��O�
1T��3��f�i��/La���h���*߾�vj,�o�������|pDJz)�����gX/�V��8����,�`��[QѴI�k�A�(둹��q�_����<�5�G$.��[8���u]^�)Vq]G8�y����\lA�s��|�I���Շ!Ӂk���2w\��X�[:�P�u�z����Cv���x�s�@^��X��V���q;��ӱ�2�e�c�v�D��k7�Hs@�>큸雳Y}[�Ӌ/g8�f�\ܶv�4��r��:���
�@�4vn�R�?4OX�R���^e��n�&�������=d"�Y�}�sd�ܭL+F�Ll�d��7/(:b�;&�\Sul`����s��G5꺇�"���uU���MQ����=��z	,�T�.�"�3z�%"�jGr��u'w^Hmp��q��J�tqj�`�A�zJ����1��cx��۫�oU����[���ۘ��R
t5v�*х��r�h��>�ks��k��#�މ�����WtHK^q��v��_.�ٽ,�.�t�x��EGx�����v��&��		U��0�V����ϭTsmPc5HK�be.A�s�7��Yri̊�w*3jF�юe��Q��I�B�x��i%���k/��Z���Hwq�w�^��˿���޻}N��6�w�2ow�G��q�W*�,�na�wҸ�e�<Ħ���N��L�yiښ���g�@�]J��p]�]�X�8��;]�\͙X�VQ�՗�ti��F�,y�M�5Ybyh.������Cb��ڭ��gs��'�,���(��d�殠B�r��rzd�����x1����sAٵpYH:���hňbm ��H[�շ�m9���b��r=\t�L�V^B:��SŖ�f�K��H.�r]�� nM�漾Y�("kN��ք�-م�7C�e95:7A���w�U����뭑�3,b�M�����K���-�k5F���
|�Lӷw���H#C�7C�`{ejA�lҵ�.�[�6�'�l��׵��,�qe澁��	��c6Q|�Cܢ�6���v^M�UA�J6�)����Q!�m�]N���Y�r�[}PN�`�sqÏ�*HoAyV�fq"��5�����ml��J �}-�$�{�]��rk;�M�t�ͱQ*c~{���F?��*1�6����˷��j�CJ_dR��߳a�/�-#mr��e�f��5�E�gP.Ļ�Wd.H�*��p�}/t<Ě��魒+/eG��Y�*R7�O/�/���C����[	�������2��ݮ�ώ��,�H+n���&a�Q	�G��Hfdo�G�MVj�{�s��
��""�wmJ�B�f�3j��Q�m��j���*!�i���CYϖܳ)7!X����K�M7xn`���>W}��E���.���~��%����}7l��rRvKU}��5�^�YJ5{dMݑ�[o	�3o��1��;SS��W�ok{���m6�������1ɉdQ<��p����ЊNO��AU�ta�D�,�B��W�/��VƠ�� �IA�QY	�6��뷏<v�<x��ׯF���[AE�cZ����m��<x��׏<z�轌� �m�sb����"+�[��T�H�����q�<x��Ǐ=z��!Q��XC�.(��\�jĨ���F�6�8��Ǐ^<x��ש `�HH� Hkb.m�7�ݍ��r�\ۛ\�5o}ޚ��ҹX��Z�`ѭ�e�V���žg�Z�>[\�X��{�*�Z4m��I�Ɗ�s���j�[\�+��F�(TY+RO95P�j�Z4^��.�_����G'�1�JD\h��(�*7?�F):���vJ�b��v�W�Sل��g�Ҩ�������Yk: o�B:t��Ɖ��*����w�W"%�I�@g�1C&"��	%H�	$P(!	�
�����A� �"��%9�32$�e��ԓW��\��u�c�򲰩��d�^l+v�ww'��l]΅'9�Q��8s�4m���)�ea����}�y�n��ų[ƚ|ƭ,ڎL��ix=�}w�w<[k��拸
2��f�mz*��]���rڔ�"���٘�Hng�rU����+%j�]@𠔇�ǧ��QOkd���J{z��dy�+�/PY���D���j*%��0O)Gt�$P��i�Mχ�����ƏG�H3�E���5�OyY��\7��L:��l]ee�
u�������;L�Y��P�t��4J��<z��,����*��E�-e[Mґ�y�vFH�+�!Eo��E�j:7�����0e6�b��1�H�L���R�/8B�r+}F9gA��t�V�b�}�\o���Wl�65џb��;=!����Л��p|Rqf*��gh�gp��6z�U�<��%@��y��g�`��ڞiD��Md�V��)ͥu��v�ݜ��}�"�l4��u��W�B�����z�7��󝽧�2�Vny=��XR��+0t�2���/z�����Z��@�6���!"�M��5�Ǚ�}�ڵ�<�%���H��x��������]�QݶpW|��r�t�$o.Uk��Jݕ{�a2;��cG=���ڛS7���2�䮣�H�)�,=�+�u}b}˔������Z6�����K!���tV@`����8��T	�R/O�_���xoW�ї�Fwpd5%�[7�v% �c4G����}~
�Vq�`ЖMTF����5۔�̔Su`����/��v�E�xU�+�P��`[�ݧs�x���
��я����	/�����Qu��yq�����S��oTɽ�Qx���ޔ���P�[���zbv�*��ܚoiOE<EN���_�W��D���0�rk��'����q�oe>wri����Ϻ�$���¦=Q{��o�ߩns���)g2ё�r��ݹ�t��"���7j�%�ճ���KXrc��")gL�Ҙ,MC-��c�g�{.��]�Ov�-`���a���b��"^�e�y�;!�[K{
z�S����"�����r����Ot����s�s�Ź��i�M��)�]�9�k���{�SQ}��1o��W[�f���QW};�@}���o0�v9�C��7�+���9)R�>L�5`m��^6H9 Ba��!#�#����v�3I���fv����K9K�<P�#���4ө���k�e4��*qG=�u��Azrh��r�R�f����H[y�j�ӵ�{��W� =���+�ˣ]�_V���\
o+���잁/����j�F�s?��Һ�5(a���wJc��gI��ȥ����v6G�܎�ƛ��/^tq�C����o?�ޑ�b�����2� ��df a�e�[��%�b�V��G��s�8�ն e�t6+Ƭ�����M����%]9?؜���.كP��k/��DZ��Qݓ3��ά��T	{ ���_矾�l괽�hnV���'C9"k�~�?"R�Jt���c.\��M�K�������ѡb���$n�$� �<�E���3=#�峆���0w�����d`�pɴ�����u��]�ƶ��d�#n�b���Z�`?��� �T�K����ƭ��nW�y`&�y�iN�ശ�9k��I�a���}g�軰Lޘ���<��9\�ק�ck�������w]s^|.Ƈ!@t�F
a�-y*����a�g�8=�&�R�˘��O�_�a��yu��9􅾏=�5�0f���]�}�1a�����hG��݁����4�Z��卛+�(,��o���,"��RI���/�˼̜�W�P���^��e\t���=y��jXC;�b"���N�Q���O�ݎ��,�v_���Ze"�.
zNM^�t�C@�`m�ij�˷�e7�7�6���H�B=Ga?�~K�TQ(��w�m⛗*���Gqx�����Wu���L��?�^�w^4ɔ��^{8�ӡ�tlK�f�9���\��>l�ۮ
���}���6^r�.����l�>v>�*�o��q>=��\��b?��_	p�F�[F���tl��VU�ny~�'/���{յ��W$�����C�ƨz������9�f���U%{�Ș�3�r��O:񳻾l1D=6p�WZ9/v�Օ	��̣cO�{�a�>9��^�.�$G��LBr�����ݳ�s��hΐ��7}�)�yH�ٹ�ݻSh�D�䥣҃.[}�̢yX7��*�	��;��zrFZ})����~�������U��?7:�I��ou]V�[�ܙ��"��d+���W����'��w�
R^�3�y��';�LL�#��[�|���)��=��>Y��]T���@�*+��}{�G���~�n�Ä�u��"���Q�Ԇ���5�Go❵󖼬����������j����uZ�R�s�Nt{��2��Ne��̓ٍ*m��T�7F_�פ f8G����4M{v��-�lrm6�1gw.2�� �s�-�]�tX/Q��G���9�-�\�jW#Op��Y�^�λu#��X7r����ԣn�V��_�S�-�\f����W��i=P*%�V���P��mN�k�ሒ5a��e7�;��5���/b�;��T����&9Ovx�O�ю����Y8�p��{l��x�7���#�X��\%]�.���y�����J7�'/����ܭWpR��7�hi*<��Q����J�ĞL��oiY+ƞ��ر��3ݦ^�b�B��o��LGBܔ�{��y+���Nd��]&���c�7B(^��d���Ӻ��K�f��͛{���Ԑ���1�c/��Oy�]�)�_5����2w-��d����ezQ]�u-N�׍�}�,�1�k,s�����-���v�)>m�.oّ��[�o[ũ�{Wq����S�zӱż��\u��b��g�0�(Ґ�gg�x3�
f�nm��6'��+a'�߶��Ӟ�>wض�(�gc>Pݍ�FV�ί,����XXe@uݴ"9Lo���4�o.U�]�!n�f�a1~�q&5}]�m0q�L0��J3�E�3��'�ڳ�t��,��V��`��,&xw�Ɋo:�p$��
�������G�F�y�&
���%^��[2e�P<3���_+ؾ;��L� �!������6�u���9t˻3�7��Kp�n"�nSwI�-��}}�_�F�e��3F���I�[fЍ���۵Ы'H���t��O"A;n�ߤ�$V�9�,����/%�ぺ_�	;L�FRb9i��L�T��U���g����߶�v�<�-�η��ߦfT�qW-ֺ�\��X�|�x����,#SkXg��4���2�;$2����*[���N�wy(��5юtz��䫾�c]���W����y��p�ܮ��5�5���J����f��2��=�U�w��&��c��ڑ����+#�]����C�ɨ~�L�F�p�t`����&�C�}�
���ә�n밋K�+Jm��
Z��Vs�U��n[�)͓^2p���Ӛ���&�&�DV��"�dc��x�@���^�>��z\��)()�;7����C0�	���L���g�}bqZ�D�<�;Dqq^�k��T�[� |�A�snD)�e��Ŀ�r#�����{�GE7���fnj`�e��q��7�F��57
^���vH�-��3؞=\u�z}[����P#������m�-ݏ�4��<�mG�)�mz}�*;�"��7a���l+����}@��q��͚s��z�����0ހ����y�_fyeQ��%olWk�X�й��t^�+��X���{5��R�[P��������熺f�'�˒
�t��^*�KW��y�5�������N�LJv�^b��Ũ�
�G/�_3���#����a�ȃ7�n�P2�+q�2��������su�Q��c�1�{���7�f�{���o�"ME	\}Q���{�s���ԁL:���b�=F.�jR<�&��:\�|9CyN���b��c9�h�tȳ�k?[��Oc����]��Mg�w��Ύ�W�=�r���8�� ݄Q���˺�z�s�|Z��Ty!������^m@������7�Ē`-���n1����/�1/TS�_�!���%��_9=N>��qY�U���}��?�#�#Rg�3�"<�^j�CͿ���d �5R4#�����w��q�]!��;k�e�ŜB����(�f��t�6Y�}.q#�2_%yk~�-�`yob�ϲ{>(o���S�q�ǱP�./��D�iȈ�}�gUp6)J�Ѽ�Z[�1����9&p�IJ���NV�+�
�m#��˯{�W�Y����b0�O��#�+�5�<�J��4QUV[�V�����ɮ��9FԜ�N�i�@�s�^�(.����UU.��Z��H1EʽM[���aR�m=SBkj,�R��7�'V��r1��W"w��(��]cw(�n1���Fq˕X0���::���
6������������[�;�l.��;8�}[��	��Ψ�IêXN����{'o��F�å��H�ꑹ�x����:���Gn�:6�9���쥸������+b7ˢ�9�8��Kn�ݼ�YPx4���^֥i�f�u���g(fy������ߤ��n���7��Sg��H��Ċ���]� �8�kY��P�8r�!D-]Mw�U|v$}�c^?��s�v���ޏ%@B�1R��ˍ������)��U�\�Zwx��q`O!t�X}ӵ��Ք8��t�d�neo!����9�]���
���ރ;R�@��1�Գ�v{h"}���J�,;�h����B���o��������Al
C_��\q[���������튆��ui�_{l�%�P��,5烂���C:ޝ
��U��Sw����3{za�w���N��z�G�s��Q���9��Bۻ�iS�
m4��Y��D�K�o+�w��e�uvܥ3C�w����'����K���E�HRW�X����! �z|�GW��B��"�`H��iUtz����eN���2��0J�q�_p1�\Gp)�!��y���Wj��}�Lo��T�t������;2��q����
�՞����AVD��VB���N�=�l��㿾5�_WX�h��T��1U���iW&z��i��a��[�,�(�O��������x<���*<�Щ~�m4O?��Y��h��N�3͖C�c[
�V��y��p�.�n��	@Y�CiI=�O>���i���-�x���L��T�Kg�ΰvdH�����!@��H2�Xcl�򃝼ELfu�ڈJ��)>l��UA��l�v<�[�v���e'�~頛�]�މ�+�4��]+|����E���������4d[Ԭ,��oA� ��gm�|y�m�IP+�p�$������mw�n y���i����j���h�Uo.T-w�J�Sr�6�*�j�w7c��g���7���B;�5�T��I� ١К�+�ہ�������n����jǞ�6˽�ԣM{n��Ǣ�:�FZЬ�@�����ɔkF<O]��C�8����{|{�:8d��-��}2���.�����F^ٖ��P�{��m��(�<VVkT�#�r;�҅]Ӿ�n��rb��N��$�{�S.��<�ۈAL���v���W)��
OX
���i��Y��Ћ����}�S3�(t7��8�v+�^�8�aj+�kZi=�(�'M��6�.W���#�Vv�┺��8!Y	��k��jշ}��%�G�wi���m5ψ�x��'���l;5�E����ԏ��5���k`#f��b���C:�h{Ctb&�fn���6����7*�����&�m����MDݨ.5�/�R�����wn�g`Q�v&�3�N"m9�B)l[Ink�.�*���}�e_ãz�mq,���f�j�<�n仏�+�1��J����E�x�������P�Fo����.!�1��w���*��v˼�ҰIh�!	2%���]>yKt+*�n�u>��/*���MYc��<6�Kq�v�5��u�mͪ���FR���Ʋ�:��,�W�ۊ�i��j�2r�XM����4&��x�(���l��c;~P�c�CWhȁ�6��E+�y��:>�ʑ��d��K'��3��Q�5m����ڵ�g��U7�ɧr��r	f�戽�#�dJm��ź��@�U����Dޘ���;u��嫢�՛�Dkˢ+^�>���t�e��}�5DuoH�b�ΝȅAȐ��i���}��H%[�fFz?^3b�2��Z{xy�*��6��<��h:*.����ݚ���Y�e��+뗗�5Sc���\�qv>���a�dM�C&$k8oU�3����F�n*�ض:�[&v�ɡ�Ժ!]�=:�7�{w�ȳ*W+l�]vi	�,�]��=Ҧu;�������e�=��9��_QI�w^r�G�d��!�dr�`,�m�U�Rǡ>bΛ�zu꼘R�I�� ��wO�bf��le��3��.8�.��a��^n�G�aV�<r�9d:f��ns������i{��K�;�ݖ�e�X�OS,����X��3�j0�e:Co�/^�Kx�G]2��p}��Ώ��WG7~S/����B�T��4�}1�#�r�N����Yg�:[�[t�\E�ג��C-���0�6��o,U�5�����îJk���,%�U���c*K��
�گ
̰r�B�|FZ�1��t��^��y%�Ue��b)!ܬÔz�]u�8A�-�� v��F1ϫ��:Iٛ�u����])�M���_��@�^U�I�ڶ�Y5�߷�߳��2@<"H��`J�>BB�H3�j�:|m�ǯ^<x�Ǐ<z���CPE�Dd�(��i��q�x���o^<x��Ց�v���E�*2��PJ;H:i���q�Ǐ=x��ׯRA{E*$��$��@��O^�|q�<x��׏=z�Y�N"��B!;I�����l��P�&�B�U%��h�V��W͛}�kƨھj�Z����o-}���n%DdZ��*��T)�Kx���sm�r�-n[F��AY�H@�����ֻ�˼Y�뻦6�nk�9t���t�MI=�N�v�r׈k�����+�n1b{�39�ߓ�9w<����ͽc�1�]�׽S�_�֬^�%��}6b��Y�>�G�*�'��͎�h��1#�vm�������>���p�c��>��}������UM�m+��'Iv�x���'��oI�-���`��9�m�0+#��q�qg���k8����(EY���"��3O�$^�Q�y~�ӱ-W�9�i�p��%��n0N�^�EY����gcl�{�p'�X�Őں���(�|��QO�k����W�k��ζ�� �֠����~1��41i�K�'�����O�}OC}��kS�iY��R&x����h���kJ��UyI�j��T�gE���{$-���,)!�x�X�����c�k�[�G]zGA
w�*�E*RUS�\�2�>��rUu��[UPv���`��1�z ��|�U{�%����Z��
S2ma=W��[�ظ�M�ʰ�*�ɰ�I��ଇ9�X�%�oA�t�f<��;�7�}UD����֎*c���>gmI��=�^�6�;������";f�.�q{���l�2Wp��y�fviFF��֋�\�y��{]	�||@>>>9���H��1��fP �W��<��T�K�9�^�E��/��^[ܔV���ڟ��C��,����{�=q>����j7�]0��a�"��v��с�o8�m������!st� 0�b6��?o��9]5�i�1U��,�ow��0��;���L㱟ʽ�����	���EVf9�����>y�T;�yp�0�Љ����r�=�s��;uء;M����(����bE:qչl"]��5�����<�@�S��s�����%Hk�? �
5����vv���^��p���iģ���o:)^5L4�.ש=[�����R���ZV.�mtN�2	`ޫ�o�9�$����r����%��\��E\�7�{}ުgU;���i��`�=�=����l*���<�d����c�<Bv�E���Av���֙���xضc��m�[&��DF��fV����Rbڲ�M��M�12��O*�\�Fj��޿]I�/�G�y�t���]rAY�"M!>�1�듪�Wau&G,�#��-UV�׊�8�=��8�e.��h��W��)uo]�h�ӤS�=������粲"��f�ev��We�._xR��������;d�hEiͥ7L�l�Մy�*f�����v�L5�l)u�dY�W��g�\�O�b=wەndXLҧv➭���V������� �E[��ޯgw��y%(��O�H�ڷy�F*v�,us��]�s����@��L#�"�@N�W���ʉo*=�2]�3�,��o~����'����p�Y<���K&����U�pR+iL�8��K�u�V(]�ՋV�c�SF������f<�AEǠ���4S�x�UJXKj���n�u��r�tW�.&�[ϓ㒧����kt1�#zlom���-J�)QhTd={<�Er�+�Wc�.��\z�m�����.j�c����6`f3��r@��9,>��z�x7��Ww(�JNN�S�������8�bE���hZކ���eH}^�ź���:�C�sl���b6�nuT�8�n'9�KJf�	�ㇵ���;2}]ֱ�@Q�����v{���V1z��ŝΑ;b����0�F۹�]ȣJ��$o�����oL�yU�����R�%���:��|��qL�U_o͗�{�y��xK��я�1�c��<3&���zCr����wvd�������b�l�o*����V�
���X5�u^�ټ>�1�F�89�f�
�Aī�0㇟Xf1	;���*���P��*�G��ş��c��e�� b'5�	h��;f�a�����{ę�����׭�t�(���x��E�����F�}c�gV�E�]k����Vw!sSF��v��#U���P> �+%b�Uk�dHǇ۴+m��e����©��v��<�Ea}Vbz��g��]����~��U�y����Q&�"�)���_��X�ߠ*F}y�^�j�Tx�x��m~��������m$�s6�g4/f��Gj��xLA�/�zVw�UR��vKV�Te۲&�uݳ�I%&8�=ҝ�u=� H����KS:�V��	�3�Kn��ϔ�����ts��|�dBN9�i��\���@��e����{v��Qܺ�y��nYd^Ż�����>dQuuq��b��{��쪣���M���Zl�����!��Y"��dv�\�s����t:q"N����o�dcУ�\��9�t�b�-s�l��d3��[�o0�����W�x��������&wI7,.~�"�:}Z�+g�i�������)�3��j�����_:����'���8=Ǹ�S�ϣo+u��;�EH��:�k^y��8t"��N	0�g1�l�.n@t��D$��v��߸`u8W��1K�;"޺�a�1�oR�()m���o��؎����%��LE�g��KJ�S�d���̳3����b;m�(0�M�xfi#�|�P�(׃��1s����5�Ǆ��.�Z�;w��f��]�}YYD@=)��*�������_�D�s��cO�[*	�S�oh�d<Uhװc��ǳ��RBROEL�2˶�w{�r��am3��Bͽ%>��뫫=���j�f���1�Z�s�|��m,oaW�^Ίt:�C������?@�>��oJ~wk�N��jjtEB�m��}�yo(�זf�Ͷ-7���ic�Z˧�Rm�oOO�;�������'��6�!�\S���N��'O������/5
�Q3�Q�V6���r��"�yb��h���Wh��e��젽��������_o¸A7�*��wi���q.v#ρz��ҭ"+�2�M�ض�u�����X�"�qXk��J�HΫ��S?U��M������גU�\\�7�}]ŢB���:����@�t%\JT���>U϶�@�m���Uo��QJ�c{Aкl���g�P���	�Ub�<x��]k�U�<D����{��������_��A�j+�Fl�V9R*�<����.ԃ�h�ּ��e��x��`[{��h������1l�A�O��:���6ߥ���v��ٱ��!|��+������]�q�`L7�^��=t�%¥��iƨ��Z�=��g���h�<�/w��M��{<�z-��v�
;Sӵ<��<Ӿ��B7�%�U����\�-����v��ӹH�9��2"�f���eH�]�s��㳼{Aُt��l	E=�6���]Ս���(�h>;�a����7���pҶP��:��_:���6�Zy抺�$�Dzg%=6ٕ|�ݢ$Y�@e[�r�ɧ_-g��C��e��NN�4�wo9����R�3F�أ�]�}[�or��rn8��+���=�hIY�sK,��ZIQA:��~���������x����&W�3y��A�����s�̓scٳ���@?1�-��݋�'�V�X��?N�m���Ջ6:HT͑9q��[XLe�h#�Y�ʀ:#�][����C�K;v�L���:=:�?	em���Kg�e	xW??�*���m�^��Q��;K�vݡX�4D��YG+{ՑCA
�U"�a�+T��?� ����=7k��q�#m#��Q��fҹezs35��{sz��N8dU�\��q�g����\D�a<�yl���v|��ɧ<���i�͗�;���}����8��[�ޡ�$�	O�%�j��s��.o,��O��i[�����T��E��&G��9c7e�bL�:;����ŷ����t�K�L�P2B�.�$ns�1U0�W5IbѣI���>��h���:��@�#-�mlBݎ}詴Cv�����w:ʹz�V�w��o[oTj�G�ԖV=FXQӭvx��gq�=�	�j�ޯ��׌6S[ઃ&�����{�
�H�7P��S8;����ݙ%r�\G���XzÕ�k&<�ǎޅ4��8����T��׬CI��3n���7w�/7����y�y����^��ekV��L�%�<s]���Y+��<���4�#Q�W�\Ƕ�ċD���g��8yM.��Y����c�v�k�������5(����*p����P]��#1P�_ߺo�u[�M-�$�Q>�<6�dr���f5���<�7@����&�F�z�ƫ��w+���@q�Z�a���kV�����چ��gAڕ&�_�w������(�֤}�Í
Oi��^�,�m�ߌ�<�����3���&jh���E�2���Q�8���1�1����kr�,����06�#�,�{:�y��#mK����޵���=7�c����x;�{q���K����׿b��4��y���+Gw8*ȟ�Ed��x����5;���ms���^�P�?z\yu���R+3\g���k䩧'�~�_�Q��}׷�S����>�7�\w<��Vt��mn�Z	8�����3�[go��P�wU���숒ZU�6�
�7����ӱ�������1���b�ֲݲ^i��<;y�{b+ݽ�~��� ���_a��c���D3V����{��ֱ>�N���l��_q��t��9G�t7ǒ.�{��ʴ���xL뙁2'�H��7��=|�lǦrc+���o�oA�ZM��U��8���Ԏ�u ϳ&��I]At��.�X���:*����9���:���J\k�/e���Kmx�B��8��VƂ���G�X5�R���h�dV�El�W5������������w��I�7̀�m���5�-\	�Ί1�h�����J���&H���'e���7���g>��mv�k�+}���\�p&M}7�.�`s����1���:Y���+�%�a�/��Ϧ�z���U����Hھټ��=J��%����=:��\v6=c��|�9�,z\b��Gm��=!��-�{��	��P�o�6�Ӛ^���M086��ij:����մf�����kTЯ��������L��6Q����A�����W;�����M��erJ�M����2� <���7��x���SŢӸ�x����c�Ʒ�����39sl�њͪ����){vy���erF�J��+M21�ǝ1�c�1�{��}��xk�Ek;�;d���#�G�.;v�rx�<=C�v�W·A�d4f�Y̬��+�3m]g�C�28�$���8���oi���*���5�o0�o/��� f��y*���q��;elOT�_�v�a�s�fH"��M׶�{��ݷ�c��K:7h��Dlzkէ��dub&�9����i9���z�|�Ǳ�fџ\ә��/G�S�&�����WX�mv[m͚��j�rIa��{'��\��\+oc��7�0�o�wQa�ހ��J��5s3-	�w�=K c����K��I>V��Ǻ���PD�P1����}ã�z��Y~;��������8)෕�z��ʦ�r�5wdMM՗����1��g�u��Ty�c�+��c�<|�����ӂ�%S������`f��v��d�O��O�Vϯ��k�:���E#Lɭ��y����e�U����5���v(��3gY)��"{�O&���t���u!h�qt�`��4�צs�K�'�Aɜ�ԙU�=����'�-����1�tF<k����|�N��UA.�6����4��*�Gr�f��W�J����Un�<1Y;�Q��>I^�u3�ʈT��s+֚�F�=��Ǥ�e�i�ܴŴ�e���2�8�7q=����γ����ۖbI���U)J�u-ԙ�<�p��Ѳ4��y��b��R��U�;xU�Ѳ��[W[#�J�9�%\9n���B�RkCpZ|m�M�+��ڝx����ˏSC2L�tʵ��m����J���z�΃��\.�NtQ��ǚ�'��3Q��'�/V�mC]q���������ɷv5ؖ��X�D����+���I9�eI�qg6cS���=˿�k�G����ǫkAɹUCB�'iW%e,�oBoN�Bb�T����.��a���2����W�`H��Y���6�^W8����KM���C��3�9�M��JE�Uոc����m��J�_@��H���\�?4椮�G3z��#���މ�K�3�9D�:�)��Vw��[�1���+�����^�޼:�|��U��,V�r���1�3zk�s�¢�!��eA��5_I�0�yy7m;]�]�hք����&B�� B��q͠C���s�6 ��hA��l��1U�C7�\��_+�Qa��e�qDh�7�U֓�^���A^�D�6q����<�h�v�v8n�k�P�֜]����{�
��i�e�5���L�I^Գo	Ű��Ws��i����Л·�N�і&ݱ�	|[7�rt�v�s�.�h��ׇ/y�}�򊅬�3�k��\vK�!���S=k������lE�{\
ӈ��H��3�rO��²i��Y�Q���j̒v"'j8��܁���Gtt^�4㗎>�j�櫺q�����msy�w:�F�
�zܵ�Q}��ͭ�d�
Q��C<_��\�I;b�h��V�L^8�N\��=�yI+r����z�+3C�jcP��3�V���$]J�_:�B�q�m���ƙY�cw�{(�ML�rls��n�����۷V��8cԖ!�[��[���wW|��Vd�M79��uR�IǶ!�ec�T�
�
Zgl�aI$'݄gr�yY�!�Nтȓ_]d��=܄��[�bE�����g0�,לj!�p{S5]�Ǽ%ιc3pJ:���iG��鋎ܬ7���p��T�A�� ��.��l4Ă��uJ٤�s.�����*��j��=tu��M�Lb����Ƶl9�xfD�ɱ����)[�hR����2��vE��JK�D�.�D������)q�Q��~_� ��<�n,"���F;|x��ݻv��;v�z����{B�r��$��ӧ�_q۷nݽv�ǯ^��)� H����`Q ��^�>��۷n޻v��ׯ`��*2$�%J�U5**ʠ�Di�׮>��۷nݽv��׬��FID%J
&��k��[��nm���u���m�����R�ג�nssj,w+���z��R�P�S��p*5�"��]7+�\��_-\آ5�Qm�\�n��c\ب���Q�r�T�GQ��I����U�\ך�J���fQEE���!�e�
	G*3�O԰g�Wy���Ns�j�R����i����A٩�c{����[��w�;���c�k�۷f�]���K�'%Ȍ`�eB��/�8$I"�%4�(b	�TA���M&\@�R�:NBH�a�D��jH�H�UeU��� 7Sw��S�.�gҦh+�^}ݲ�4�՚y1�x�k��<r�U��eq~��:�M��d?��
��/����feq��W���qE�s��4��G������vq���5F.�r�R�0&�ߴ����*��҉��F^��+p1������nob��7�G�0.�eإ']w�y�mq�k�A�yy�5t��'�=0�s �})�h,�qe�Ş�7E��b;^~��4s{r9G	0�\*c�EMd����wro����g����#o
��`�`ǻ�������i�	C��Ԯ�F�y�?�Ͷ��~~�}�'���ȸ�-r1�N�7l;��x�5�jG* �>VQ��~�d��߇�#��γ�����~�Ե��QEy���o�M��K��gl�<m���Ҝ��B��hD�}ՂjƮ�aB;!��A���^�r��R�O�^=y�;��L���{+j�m�ܻ��tw_ep�]]��#����j��2w�:��_J�{�v�n�̵�o�)�7�q���ܷLC��Xvu�uZ"�Ǌ�Z؟W)g���E�R.ķ}�&��y�R]33�T��%%����3*?�1�I�;��3���|0�"�+�����������JTl]��Ӛ����]�c[�4F�~��\�50�
�G#��k.Y�{ͳ��7	&�l��T�%�����[:�4� �:\��9�}������5�X�&���b�}�[��38�s�lv N��p�f=�r��� ��[G>�2�� YpL��4a�����X���6�Z~����}���d	�uf�X��Eh*D�l홭Z��@����x.�	�#Z�E��򧎰��k�^���-�n�+�����R��^�U="�N��?% R����*x�L��Wf��/5�<��g��1I�$zve�R��h�>8��"p�X׵�ƚ{�3б�w짟m��o�*`y�Q��ȥq�%�YV�&o-����tZ�U�f�=�L{��:���z���ؗ�QR��z�����R��8����%ێV�T9?>�/�����u��F���Ez��v�k$^�w���M�;42���W�+�ۙ؎�;�oȺaض{9:���\�����/7�UyY��J�n�m�L�5��y5�0ɜ�g9�U���1�c��w|�_��:������o�c��;ͦx����jn��CB�����{k��w��L�����r��'t���G��{j�-νQ4*��Ts���o.N�j%΂�=�盉��v��>*�+��N%���[A��Σo�Ū�8�V� �=��
����@麿B�szAq"Zm�4,�z5�q:/Z6�lk��CukN�Sê�΂����f��Q��Q�U��q�˝��ni�G��3ʪ�p6�i�i�Π��ג��S�Ԯ&Η�ܸ��[�h=�:��xJ�JA�5Ot�寠�3 ���S��=e<=�mNr����|�pĊ�f�.�x�)g<�H��>�Ct����ڡ��}�L�ኅ��Aq;`=����
ky�V�*��\o^���6�]~sX]��͚�;���!�;K��zB�]%������yz4�V�>�~�����U����^J�<���v��<��L����ǣ����԰�u��[�vw07�[i=EwV���@��hy��Ji=�P�����J4�.NYl��Y��˺�W)�;V�7��'S�r�:U�;l��.;<�y��o7���Z������U���Wz_��ۼ��o;���Wi��P��o^��Y߯w��Q@D���i�:Y������p��+�GZ�fKȥ$�+ޚ�7��w��y*�+�I�^����u��`�#y^X����)��������m���,[��=�b�{c����w��m�m����GVbޡ΅�,�x���y�8h�����{�ɋ��7f����\�C?�_3�7h��������"Dͅ��X\�r�s�L6EG���ƽ���Q���Z���޷�X�7׋�m&n9�7��Βy����Eܑ>'SM���>8���w�3u��X�So;�
���;;$
�W���}<z��Nճ����!'��:�T�l
�׎�}�egY�^ۈ��R��ʠ��N՟\���vlJz����5i��qw�����f��ٔ��c�l���W[^N�U�3td*�ec�F�"��x���G]�;�muQ�в��d�b��Ŏ�b�h�pǮ���ɳ-�oXGk�]Jţ��3�:e,�%�Ө�J�4u�>c���EY��h�{��������?����[�����+����O12�_��޽��͙����3�X�)S�ޅd@���r;�C��%*򒪟*��zU�­��\��ܒ��y,cY��=Y0�w� oG�J���V�[t�{q]h��O3ta;�� �O���G$�ar�+�v�d�F�é�M�{tj�`�s..�8������M����^���@}gы��pK��n�o�/1gr�Θ͈�N���:����j3[c�]��~�B��C�ʬ�~���v}�l�U��
Y�<u{�,��c��\^6u�5����Y���9�) ��G�M�݃x�����N@���[}����fD_�5���D��7���>����jv��ƣ���T����w7�X=����i�-�"�f�+��b�<�߹�eLFrV�ת��ƭ"���3��C���,�)3f�Z��l�������f'��'������
蜳ϰ���߳��2Y	\}�=��V�Ϟ]��eV��!;���"�l�2�$��:ү ����ٷוvfn�T}]�A	\MeIZ����
�ӪjL���Lr���
��'�w�
7;Sx�}�����������@ԗ�ѯBz�`9�D-�r�qº�I����oq��F�wL�nꚓ�ŹO�r(��/ג�;=�t,��z�����󺀅
Eg�9V�
GF�8���R.�n6Pƈ���U;�{��c�!w2ϧĸ��*'�R�q�\��e3���I4��s�}A�TX�-���U�����&2���-�^3Z�~��������}�5}��E��c�ۘ�&�Y� ����d��6�5�^lL�={�D<��D����Q�N�K�6�P~	5�͚�����q��6�r��G���]�KtU�3�uw�.�v�Y���Gn�RJ碅��p��<���w\f�qu��}��_'�Uz�st�7��V�f����]�z��`Go��M��v�Ng��]��WoPG^qA(�>�Zx)�6b�Gw�r��L�XFl�*��=8�,t�%����:�<W;�rM��뵺SP<�����fX�[H�e�ss6�pf_oq�U��ʫƃ��)��].c��zm�ܖ�rA��hr<��=j��[��9�A��c�3�o��;��o^kZ֠4GH�G���}}�0=tL��N'1�q�U����1��$�tދ�2pD��o,��m���r�6��Z����r��&1Rӓ��sl�̿kq��Uc�r}�c������t;�37j.؇uÁ��zA���ѺY�����^ �Β;$q���:C��?�s8D��f�σ)��5ݜ�h;�pg�3=���"�@`ǣH��.S�z�y��'��ʴ�3��� {{B�Y�4I*���,h��hDi.L-�P9��(a3�5�[�TT�z"�x"�y�Ѩ��N��np5�+�c鶧�&ԭ���t6�u�O�
�7�,�1���	C�]�W��	��WW��;?
mb��`�;�~'	��Ł���=H�N�`Mň1�~]�Oͭ��]��{�"�I��G��G)���W�z�/�rsI��E5/U6t�%twK��)��u[����7�\�ɪL�G'�&Q��.˴.y^�7P�>��Y{Ʋ������:���oH�?	������ؕЬ
��(�r�-���b�x��X�Ң��1�����V����u�5�̧��1�9�S�eq�鰄���G��ĔR�"8�˅@v��fvϪ/\*V�h���_'oh�B���W^��fbR��!���nlLtg��_M��:��ӻ�p���!�� ~K��歎Y�W];��*��X(��b����Ѿ�����x.�к=D��F��=���Vg[r���O����<�+��@�GLB(%�>��r�'��%9�չ�������ŀn~��s��Y^�p��j�6�A\ecc�tN3�=�Ӥ�`�թ^U��Ք8�1�*9� �h��7�9���`i��4ՓVϫ;T	k�@�2�{��Ǧc�1x7�p���k�A�J���}�%��4Q�Ƃ���<y��b�Nk��d5��tW��U�f���3���Mŵ�A�u����8@�0'�&��9��B���$<n�"�)�i�o ���89�g]LU��Æ�˶�v&:���v�d�u7�)�㛹4�H��}X���4�ު�X���K��!8Sŷ�g5%Y��15v7̪����G�p�S���pq�7W�p��ݍG�fb����;y�}��9�m�o��8�/F��{~1�c��Nw�̣}��g�rf��:ԓn��x��B�58,7��Mi�T�8(�c�IN�����*"C�O��Y�Q7����;u4�Q痯l_�,wA	\�{�A�:�9��t�V��l�7��N�+��A�F̎=m"���ní�΅/C1=)�7s�:�q���a]��!II���~�K�0�~�f��?z����	DR���Sr�dE,�NA;Е9N
V���C�����Ch�cmU1�&��\o,u o���(��<��s��6Gk�;�홮�t�������B����P�G�TW&C;��{�ŉno+q^Β����gݵ���R
CpY1����x�%�v��Z�1}�[���=o{;]zGzK3�މ���}�޺x+fy�wu?6�Ca�6����D�>{��#Uͥ>�o*y�O>�}�B-t�g�cQ���Z�a9�Ի{�3��P��F�$�Ź@[�[^D�Q�GX�d6�cVh�r�gv�FU��"��}�����N�	�Y\+(�uL�P�����V��g,��Qq�nvR"���T��}��ޮ�K�B.�Jf�B��٠���������5f���>���8=����3���[E��R�G�N��ݯ"�e�37����ŨW�($����6Vz�N:��ś��t*��<Jd#���pރ���"��v13��r��.�7�{�GUb"����M�h��S6���{s X�mmo3�Z�ቢ��V#=��؈-.��/�թ�Z�`��Q�H��ĳ��OA�������]�,��д��+^���e��^�����v��A�qY&����d��u��6�t�FX�y϶\lf43����A�j��S �Z���"dq�J6ג���M<l���i�n�m
����d+F}���<����,�%�2.���Ճ@u�t\s�7��r����/�8*���b���cP�/WY]��a���Q��&:0�^�u4���`a9����@���Դ��A��A=�h6&p��ݳmS���Rb,�!���\!��]���p̕����L�:�o3kS�����K�V
\�9�1 �}��8_�;U�j"x��{�k���`�#K7J��`�݄�v���vqv��6jd��p���w#��׽�r�@μ�����㱬+]����N����b�e��i��<[.����k{�VwR�Au%U��0ꙷ��f]��Ҭ���*�E�ݚ�k���aw���c�;d�<�Ue)���HAe��O4V�q��ÙMKy��q��Ѵ�/�m��Q[�)�}�1]�ɍ]���ŝ3T��br`]�^���]�Y�gk{
h$Cbv܆�a\�v�Uf��u�;��7lX�|􇉉SkU��&=���ꧩ3=;
\���p�/ �Dr��$���{��j�U�G+J�*�v5_=���Y4�əԬN�������2|���.�}�l\S��/3�N�͔��Գ Y>�I��wx���=͘���i���i��.��f�>bY���T���T��wVI�-�ޥw�b�B=/�ŹANΓ��e�]�O����]���K|Q}�x�����ȸ�̓m������[���H��� ދr�w=b������g�V�Q�v�梮�S�q\]u��/�jo�qT��;Մf��)����W`�X4mt�+%�}m�Ŝi��݇��}^�,[�����υ	g��YfReɦͷO:�$�cl�U���ڪzZD.C��4��G��~0�"A��buz#,O.�7��6z�C\hU����]gq���+|�s���>Q*A�*�$ĭ�4�/���G�8�7�y�'�̮�ϻfe�ҚN�O��WR�O��j����ĥ��m�vkc�K.d��əFMg�y0�a�s#�v+���
�ǆu��q�6GS�)����0�՗5H9�K!Q�w�	��w����jk��#K��Yf@�8��N ���V��q)�|�r�z�N�vp��n+o*७C��VZiC��|4j���9�y��0Q�'O7q�-r���G���敒["�u���Mۛ�Ƌ�Tnur��s��'�-������u,��VT���В�]�%%T����pe�e��.�1�3�ف
�9�m��`$* �.{�ct�I��yd�4��uɻ9�峟�jv򳝕��w��%��}�����g$�s�Ö�첯q��tT5�dLݻ���3�ŗ;���;c�̮���m�j���)���9��"r��wfxGf�A��&��a��ÙS0��oB�Sp5��7%�:rݖf����K����3�#�y��7F����7t���]�9>�	�X��]��T4+W��r7*N\PT�p���p/��U]U*J�3��x�f�e�ɍ��w��f:2 hWE�Cκ�TJ��:���JkS�{�xd��9O��Ɍe�)fK�F4��A#�5����5��-Ζ"��D$a|m�^;v�۷o�o^�}ƽ��Dh��qҌUUP
�Sׯ^���۷nݽv������i9�lw]�����D�Q���$�:z���ݻv���o^�zHIڡ*A��*��)F���4�wK�9Td�)�ׯ\v�۷nݻz���쑉 ��`��]�^8� �r��kƞwK���m�"4w]S
�9Ўv71v�.�H��q�×
�xב�z�1����77Ll.�ۗwn�̹�܃D����g�l'�q��I�� ��`�ח�a�-ۘK�D�;��t �4���\�Q2J(����s�E}�I�J"� �Ai;�e%�g���%`Z��FU�����a��y�(dkz�c6L�6�j+��fsF'�bc����c�3��>r�]��!��7[����|<T�
J�ϵ�.�i�W���ڢ�*��o\�f��P�&��8^7�%|�6�I:��:f<��C^��/\��<-'�q��ui��
��4��~O�k��J��uQ�Y��,��-��z�S̞��ݵ�t���V�L�z�{W��K8��k|�$T$~��ۧ�t�� �R#'t>�Ӽ�@ƾa%��^ѝۯmGT��i����2ǿz�p���B�z�IiO�=.�f�*^���{���8�������~�St즭-m
�Zsk���R��kl7m*��~���� 鎐�C?�sE�k7S+(?����WP����9?����ִ�o �H��pOl�B�xַ���V��-����#�P���VmuYqWF'u�"_=�hDڷ�q�Vݚ�#ki|s�igG�L[f�˹�ҫ�au;߹�gt�\��tM���o�΅s�Z�'&���޼�w��H�,�\OM�k(�S����'2�WY]���t��e-��9���d]a��T��Z���'v��c���}��d��VF?!V:��H�U�M+'hnp<Zz�&ʹ����ݙ}�􈽓<�́��`�XI��ޏh��b�ndv��c��(�t��@l݋�Er��'OTTK���+�b7L<L��e��9������H����ԭQ��z��C��*����Mm��iFm1��e���B�ź=�Η���T�N�J���B�mV���j����z��\�|%�d����]c\����&<������MN��ױS�uk8h�>��>�k��-�����dx�!V�C��Is�Wf�Wۙ��7�5L�m@����i@��s�e�F6vѿ]�k�A���g���!��^�9�ea��8y���xC?�Z�6���ż�Q�,��y{^5J������룕Cx�U����+�:�B��!ߙ̣�h��ŵ��dNӸ�S
�2k��ԛ+k5I�׋,����{NF���xI�e��=�v��=l-��g%�� ���	��P'z�)v���0+ڜ\�c�-N�T�ܾ�Sf���2�+��SI�W&����w�c�S6f+<���Kq(.�rsW���]��)�<�O�1�cy��]j��M�͗��M�ĂU%̷t�3����T����ՕǺ��W������p���4ql�p�L�S��+�+��%�v9Zb�ol�3Z���մ��٫�Wh9���xo����|�]y��	�7���6�S�SQG�`�U�EE^;�u����+u;�
tY�����*Ѡ2<�Wn�Jٷi�Y��wb��㺈�V\�h~��t �l=$�Q�4�&�3m��k�2�YlP�7YxF����@���ܟ������+D���+qS�;�/��L��z��*����f��=M��n%��]T�r�DX۴3q��z��z��dϯs���╆�pYR��f�w��qU��'7k2���w��&k ;��%-�~k"�<�Y^/�Z���	W�6�֯X4]����e;H9����M]�`��]=;ѪQ:,��̵n宆�4�A���b��6�g�[�n���0�]�2���t��0{P{�������+�$�e�O3�����tC�y����7E�ǫ�4N«�j:F��2^�k���l��<���;�v��N��"�݉�����1��^��3ɝ�|ןG���{� �<���N�\�����&|8n2��Q��w��N���B֎B�l���ɶR
[��jB[��;L>��A���̀0�9*�ǫ��G]�w ��#��|�U��ޅ�kx�C�g�'�����>��m�5\Qy���8�ɵ�7L;�#��*����^t{a��\�:�0�Y0���7��(���@Ȍ�\�z�ܞx�%�5����2|�Ba�.�@ˮ�cc|��>�س�b�6�]�SV���Q ���we뮀��~��|>�lϠ+�H��x75=�%[��ձ�z{r�[��ŷ/�������Pl;ǈ�����<�ᖗj���q��ݨh�k��N��F��m�3�Oz��-���.f�#Dd�Oc�5��Z��zV/P��W*'��#�x�e�=����O����&��{���ާ��qi�eEh7��z�;� �Y�]Y����sk�i��[쓔Y%���N���2(��1������s.Cse�]�2���͢椚7s��p�����r�R��Z*\��H�4��jo���Oiڪ���0#��Κ�|ϓ�{�+Thִ\�K7@�j��O��R��B�6�F��6!�g#���"��S\�qA\Z���\B�<���mt�J�#���l�ɧ�gv^H��S�^gz�D]��{F�βzpou~��e���WW�R�)铕z��z���������9�kϷ~۟���d�&�����ط^(�tQ��RUA����N��wB���gmcr��{�6'������)_:��'W���c��=�v5v��Η��\����ȭP�اQ���Yܢ�\�n�f�x��<�2jo}�4V�`h�#��-���^�{��ga�##dm����\���J�k�ί5U�}R�e��������*�3m���Fl0]u�b1O�|k����uq��1j��Z�w&��A�
�5���^��o0(ߣo,úO���-�!��=��nm�SJU��7v�U��ʗ��qf����d420��k��.k�"���X�n�uJ�W���~��"q_^�"�x��sub_o�g��iխ�lVx�fb�u&�{�&��7�]T�h/>>>>>>����A����˫�VW�����e�!��;ຶsiJx!��c��r��+ܽG�1�$����������Z�hrM����	3tg��u�h)���5����z��	���m��:c��ͤ�=�~#�l���^J��rY����ӦC��f�(��g*��#^��[�F�$C�5gV�;��_��ÜJ�u��Y��Y������1���H��N�3*�$1�=[V�g@���h!��dT뇺Y�	4�s���1���ՙ�95v絹#�ʫK�������=�G�M��~!A]z����ڛ��x�^��Sz1���.�@�*=W�t���hA�}L��Dˈ[����Z@c���z}h=w�$c�&��%%��T�K�'���1���{�9l����_O���{�d���om�����+xk��4��U
�������LIݬt��R:#҅���n��\�vi��>�(����[|�X���N.���(ú�΍HW�T������E�.b:�db�{w��:J�&����T�����^wttq��sw����c�C0����X�F.�UfS�����������>料}�q�]�
��wq��U$	t�)+r��R�Ha���MUr��c��,c��7�W sEl��mp�EE���H'9q���+ҟ�Dc�����]E�bn��B�����j���h=�e�%���j-2��n�_e��$>����u����:�E�"��ms{�w��;�U�l�؀K�{q���{�҇�Q�^5y��5�2S������)���;J���J�:�����|�`�̭���H��>���T�i�]m��S;6���%z���3w�e��u)���Yb[Yg�4�!�B-�� %�z�R��D��Q��wa� ���������uS��g���£ё�4#*4k����0��yź�����$en]�	/&���\{��t/��K�Sv݌��]5�t�Pn���n�(���6�vͲ�zo	U���{��TsR������j���܆om<5Ch��p�N��g{��-f���UR��<C��1��ʎ�sUn�3<���!q��j���;�Ml����+V���k�5�IoT�76��<�w���T����y��o7�ٞ��F��������;|�����i��Y������ܼS����Q�8���c��A�O Փ^��aWi"B��nf�����v�G{�>�6�P�����
����9���I����{f٪�훏;��T�W*��*��3MP9�7^�9�d�ܥ��L�Y}�0o#�nE�a&;G*�k�]\��:-��֝���T�]���iZћ<U�EW<�+vz���l45T������.�9����籋�� ����m�������үڻ����=07[u�?q��%�����)!�n�EDr���u����d�(�{�+�)�ٺH�{чp�O���|�����վ�����3�ݛ�I[�6{ck*.�FfW��;���)g�F��<(z�F{��
݋�2,�[x�|��k�8o[o�� ���̫̭�C��f�4!8�zO^/G�f�pY���#t?5\��.�1�R����[����m���������$μ�B�u�������G��e�x���s�n�c��.�n;�H��٧�j�:�����Y�q{��|�zh~�^cs��"3ݰLl��֯o���r�Qp�v���8�*_��䙷�S�~�gy��8�������M�?33��ǂ��{c
��G��3�X����H��|3ڴ
x����.�z�����/�0�#��F^i*�Sљ�-��������Ya{��S峩���4������0ᰇW�=T���˅���T�.�d�{�yڂ��hm�o�fnz���,₠�y��Q�.J�ioaVo_m��n��@���wv*=q��\Ά�
�ty��
�7U�ص�맯u����/f��B1���Y6�M^@�Nh�2�!�C��~�p��J�<��9;^m�IV#%%T�Q���:ދ�y��iB345�σg��׿W�����eS�?����.pU�&�����/�s�6�m����mˎ�l�Mc��g���@�ܗz-gK�U�T�s*��["c�@s�^�&��2��T���ok�A�E�y�D�#[���|�sv,�C��)UrrG3�wQ��99El�5_;c5u�w;��՝o܃t�+n;p��16��z��q��|ɨ�{Wr��=�H9Q��ݿ	���0��2 �@������f�k�`al�5�ȳ�M�>&m�f�W�咷��C<�mi��u�" ���evAk�x��6F�5#�ԝ�O&C�ߵpf�}�X�Y��|W23�;vӠ�Ur}���6���3�/����-�m��"(����A��!������Ⱦ��"��2&G��5M��+�Y����zz_τ�ﮋ��ٯ�_�q_9��$�c<^����	~z�u��Y�k��Kb�k�ݫ�i�6����!�7� �	K�a�z��������.��STG5�B��,��_����]r9�̌!
,�l^&.�����ܴ�������a�+�)V�dI�������h�g(���<���~����r��p" �_�A���?���("�2�*�G�ڀߔ@$BF[i�͵++iY�JͶ��m1�m�em++iV[i�ɛZVUeem+-YYV�,�i�J�ƥ�+5��fLe��1�����������Y��I��X�UeeU2̖mi�KmfS6��m1�e[2b�m��K5YdɕTͳ&L��1���ԙ�ic)��m��m�Ŗ�ml�c6�X�kY�So���dԪ����S�Z�jmifY�ef�̱��Y,��Q��ͳR�,�j�ͫ�-�R����MT����T֌���m�v,el����YVVj�f�+5ee�VVʳU,Y�,Y[+-ef�cSVVV��Yb�l���cR�����YY���YY[+*��l���ͬ�5ee��������C `1FckѰ|�(�1D�
�P0DUj��Z�Y[U+-�T  @`���H�T���J�کY��+-j�f�T��j�e�T�Q ִ�Q ��Pf��Vm�R��U+-j �� �A�کY����j�f��Vj�J�mT���JͭT�
�@`"�րt�@`)�$(��@b���(��@b�T�B�"2���ZVmiY��em)��*�kZЉ����+-���J�m+6���Ҳ�+6��v�1���em5m��+iYm�f֕��VU�em��
��
=�� �,b��(
��������_po������?����G�����f���z5�*��������_��@3��������
���q��=(���@�@b�O��	�P��؇�@���?P����t�
���6����NX�~���(��`���͵3kJ[R�ZKm)��miMZKZ5��֍�6jҖ�6ԥm4��KZ5��miR��J�����"�Q �P�T�@#H)� *�5M�-eZU��Ֆ�"ER �	HE#H,A"� $Q"���Zm5��ͭ*�m&֕�֚�SJٶ����MY����Sk)k-+X����j���k)���Z��ڍ[mcj�F�*) ����P��B!�kI�h��͵���dHED�!�~A	C����S����kU���TU���}����������
����B�������*�~�?�������0O�z���g�����a�������_�~Hb~�a�r* 
��A U�(xA��j  �����^�@|O�������G�a4������>ã��l4�j�������>�W���@=����?#�O�����C���?���@}�C�����_�����D,$O�zs�M������~g����s�����I{?��߸ߵ��3��UU~���{ન�S�l�'����)�?�1AY&SY}�_@��ـpP��3'� b8����6��-j��M�7u��֦�M5Z�l5kCUF�&��ح��i�m�f�[mP�+Si�M�gGdMm�q�F��:Ź���Ff0�̺�wvݫ��s���6ݫrTl��ݱni�iZ��7rͳ��M�sv�wb��륇sZ��ik�ή�L��9�mٶ�g-���K�ۥ-un�n�;n�����%٫����V���c��e;m�u�䭹nr�t�K[65ձs�fڹַe�K�����Z]�]�nW:�ܬ�Kc�v�V��һ�m�;;�tՊ��9m��NN�7n�5ۻ�;�3��]n��cj�x  om�JA�]���m:��[ݡ�y�\������eP�/v{{Tmj�����y��M��<��W^�@9+W�k�=�u���� W��v�:��[�C��ӭ���.L+��l��wm3���ce�   ����P�B�
(n����
(P����� �P�B��ﯞz����m�w�� u^n�ݫ���l�;�n����T��wE����:]nݝ�^������w�h5�;�]��N�sw�v֧uwm������  x��������]]�wv�W��v�5������כnӥ:�k�����4�N���ph���;n{Phӯr�{��[ݪz��sj�Z)���8V�\܅��s���v���� �(�h���n�P��y�]��eO{{�ֶ���^�Z���G�[e�ւ[=nP�u�]��S� w{7z�֝��o8z�v�v���{�{�2�ڥw].ٖM.� 9��A�+|�\�kV�ikˍ:+����Ǡ:=�=��F�w����U{���Mb祸�GGv�{��m��]�� $��.�����kf�wk3.�tu���}�o�]
:����oF�)�7`k{޻[glt��Z�כ�z�E�r ������խ�p�{wz������;wl�sm�u�[v�vm��5��  �|�  �=��  ���  ޙ�  {ޭ΀ ��< @w��  �ۼ  YF
@	�V�ov0��v���u���ݶ�v7_ />  ���  ;n  wk� 4ۼx  ������o@ ��ۀ ��{�
 r` 
ݼ�v��wM�m��U��v��׽� ]�� ��S�@ {׷���;�p ==���A� f�n �{��{�  �s�� y�@.��  ��ZZ2�-��V�n���nr>  �|�@ 6qp:>���t����{�  x �]�� ���{� �w��  �p  ��  �S�)J�A� �{#R�   O`��*   "��Д�$h 4d6�1R�M2 �B�4��@ j~_����W�s����ua���Y3���-/2p�Σ��t~�=w�G�fw��F���"+�^u׹��TDE|D S�U_�TDE��"+"  �ק��?�?�a ��P����p���^	�p��f��H�R��=`dئ��tҢ�c�-�,�):iK�Viֹ�4���em塳6J��j��C%�&C�a�LDڧu�SdJڛ)6�i���$�
F�ݢ�&n�*:$4���zUFn�t�<��IP��3E��-��x�;����31��cw�8`�	nȝ�EAOL��C�6*��J�eТZ��-�e2E��x� R���ӳ�:��&�G%�K51�SH-�0�
��sT��n�]Kƥ����y�Z'd�lfC���F�����@U�kF�L�&�����]٘��u6t����)��;AY�Vdt��[�	�J��]Hb��T;D��,�C{�\݊C+f���-T��Т�m�j�7S���N�`%�$;��,o���|h�W+Bš\��)�9'-�-���<r���P��M�Hsi��ɲ��n��:c�֍�krT�f?��N�3�4���d�tm���P�D�D��|��r�wov�h�4�R�h�4��cX@���ǯD"œ�S�u��S��6XTE;�v�QdH�u����&��=�6Ԗ�"	Mdgf,͌���V�@�Və�#e:�Oj�b���k>�cU�06�3v��f�"�d� ��+s�G�SH�tM�1[�2*k-���V�)/] .�Mh�C]�*;{E����,YH�rV�
�Çj^4ckF�*�����7� ��LTڠq�<׶��(��	N����Y�'ҊPfl�H9O5�Z�Vt�����U*4���W��۸-�cU�E֢cTf$+Lgc܂3��vu4z�ON�mh��Ő7´mo@�&��Y!ԃ\vf^��*�M����՛T��e+6�{W� 9N�+
H�2�7�4�����W���!
�ք�k�U�%s8���]���+��5-��\��Ի���`�d42�ꁜi�śd�X�҈*�-d�E�f��$�f�7�$�҅Be�VpM����F���	���d��RL.� @�INM1��t�>̽���r�db
V�N^:�k(�����=ț��m�a=F�Tśzw��D�	3�V���U�l�����H�0��db�ۮ��k�A�b0��3dô̋M%��`u4#n��T@os�7�H�CI*�_P5�7j;�Az�2i���Q3�]�nF�E��P�>-Q��
�jm��N�,;�f��h�t;7B�J̐�n���ۡ�*�o�^�Z���we�_m�B�x\M��U�Bk`T�Re���b����emd,c��(i�A��4����\K��U��ѡ�V�4�k�6��㶁cq��Qav��w�q�t@h��]��f��I��eJ����
�I�:>���w#AEܸ/k劎w�[c$�4ެ�,B4+��K��8 �����J��9�hV�vq޼TN��&�nնwq�vOrm�
����>�kn=3�: �Cd܀��rb�����!A�.�6�E�����)�Z�܆H�<)`fx��R&@Әc`���,kz��cV�����Z�鍔~����]2�SQ�%����Ŧ�v�͂�)�teHո�v�r���+�Re^K�Ze�V��.<n�����l�߱����(��v% ]��j�k���`PYri��[�Z�C�[%��-�u�!6�&��:�*���t��-�  �E�LB����V���Vq���!YeU����7/la��Y�j�*XY��QzcdM��Eޤ�Q�됼T��a[����a�ll���ݺN�-��4�Gh��YVb���"�Z㽥"̱�wLu��h��RYt�`��.�܎#��d�X�:�RB`�wǷm��w���j�?��:���DlS�G@b�taH�Ѧ�A���1� MF|ց��퉦�H�A�j�‒T�a��l)�tf�;x�'Eث��s.�fm��̗���
W����nAZ�eaE(�˷e"Y�,�yB�A�n�H�	;J���c8����"���r-r�07$�Q�����H�75�>N�g4M�A�6JPm�Y�#��^�ڻ�\�r�v��ԨX��.�Utӕ
J�s]�[�å�T��:�F�*ZͻsS��p�ވ�׎�P�V�6D��U�L�����I��c/nSZ-��݂&ˋ�ڈ�Fc�t�b�M�*��e�ӕd�Θ��1	@#�fB&��u(�%S�e�Jؚ݁��n�	4��,`JR`����:H���71��=J�bKyze��b��9�-Z��b��)��������*#J�0�t&�mS�V��t�����v��/tRlAD�C��=�I?c�O0��u{%G��Rkw��ş*d�ئfQ�-����l��ZrV�b�<C�W�c��K{GEl�:J��*�۪;�x�фᕅ)�r2Bְ��4K�Wux1˙���	�n�5[���C�k�30͂�Fʻ�*bG*x^S��̶&AZ�JNI���n-7J�Y �%�܂�7P�ZQ$��Z�Nj��5R��1G
�����~�eR�L,�%�!�T���ю����"���F�ڮ�2��	�)�����QX],m5�1�EɁ��f[�}ݒ$\���d\n�A���tNQ���,�IP�ۚк5�jQё��^Kݎ��o�M@Kɕ��Hb�n�uJA�܉�n& W��MVK�V-M��e,PS���{���&Y�@�3h��o1�j����̼b�3qԤ�&N���Mxq6(	�-%BR6c�s�Y/m�$!�`R�	���)�e&|(*�6�^i�c.�.���&�i�X�f�y)��T�P�_b"[�/ UiR�sF\��Rw)���R�yx��T;7ztn�*V$��Kt΂chd��kGƋ��EjE֊��>�L�c7$ӗrHe��!��Ƶ-��62�㦪����Cq=���T�lL���I%$"aG�{w��Ȯ��X��j�:��b��D�3,���[H����w,ȩf�pcy@n��T��=�ւ*�X�{MP���g�7�6�pԢ�Y��ͽBd�Q&�Ŏ)�S-���i���z��4U�3L��]:U��W�$d�!`a'/`k,3��VY��/t�n8f���N@�ZB`2�t4�f��v�	�/�$�uh��fRt�k�,(���)��	?,���L����Ρ����#[״Ҁ���,����MQl���F������2�Z��� �+����b����������'�m:�e�0'V�ld�����^���+^к�ci�aƫ>,���m$�c	 $ȩ�V�Woq
k^^Qyw�Zy���s �e&�$'�U���r�wK-/�K��c�.��)��M��V�/wբJx��cL�p}�)�l�5����y(;څi�`��S�T�qD��Rs$"���SB��õ��4�ū2�BS4[�L�ܕ5��8^���EY�n�2��yW�1�4�m��h�V��C�m�ئ�&GR�H��͊�
���J[n�H 72�HJ�!ufA�"-�zY�݃�]��t�F�eʛ�"�1�8UڧX�+v�ct;YLT ��t[�@��Q*��뽋%m��3�����76"ݥ���5=�]�B-�`��H�cG�dddg$���D��m�px�m<giʵt[Z4��s51h�u�+���d�(��ħDQ Օe���BD�iY�Q��t�ջ.��̀d���&�r�ZZMH."���5�OE��e��R@U��C�1�^���#������V� ��&+��rjh*�
�aK&�̦U��w�Yڶ&��6�E9��M7�"sFD��`DU�42�j�hk��l�V[����
C�=H��=b�l�7"�k D�-���j�Y&RW�)^�n���%$vS��۠Ln,۷1&h������5�)mf�4�,��:&�����<���0`��ٺt��}��Vje�Kk]p=���I �w�������fܥ�ZRC���`V�RG"���@F�v�+1V@R4U,Y�V�ݹ0��;��w2�����~D���@�:27VE�eY���)���n��Z5m�i\4��)��*����E��Wgp��F��3��){�6������b�N�Q��X���mƂ�Zһfm��l�7c6�-���7$��Aԧ�n��ՉnJ�+)��� (T��nC�3��V���AC��»�� RIkY5 �#bz�J��!&�ME�H��,�`	w�L:=ѯ*���Xu�Wkk+V4�b�M :��` ��5A��lY�Gz�2��o��!�� ;����pS+4�c[�lPn&� ��ʭ!e��z����%]���Jӡ��-%�єDЎ�f�1d�䣲т�A��!MUn땲�l�S��{&k,�D�T�����I�.���53!�읫�N����*r��%݈m8�ݺ�B��-f�ʱ�"r�Rc+avq���(�H��양�Ěh��f�ʗ`�r�^�A��<��:�:0Ԁ�@���p�{�}�G�N��Kq^(�ܺx4��D�[�&�V��P������y!.�)9��A>��K�ڻSM[թ�A�
��s&���in�E^��-��0ȓTQ��r�
h��pLr䬼(��Z�^�(�[�5�M	�9bL�r�U_�����*2Z�5Fݰ���a7��洲����;z9��4��B�$($h�x�,H뺸"_fE1ن��+Eh �PK2^ټ��a	�r��Pu�k,`gL��hմ%[�e^�Y�I^�S"L�5�P���:L�����V��b�"[Q�z�]ү]�+J^[t>U�Q%eH�1)�(V3
z4˽x���j�H�Z4b�,C2`����o� ��U�N�����@ñ�V@��i��� ^l��b`n�[���b�Y��R�[�a;Ő	)	"�W�V�&��h�ïo$���Y�E<a���lfQ*Ɗ�Ŗo)[X�i�Z�3T�%��7�X�z\Ȗ(���ˊ%�g̱ ���eh�Ɔ-�+x�[�����N�ݹz�z��@����yJ��[�U%�f���rj�Y�&X�+Sq]�Vv+�I7M�I"0���A�iܘ��ٱD]#��[�U�jC"�Ғa`�2��iƚ������P���R�wopR�8T��4�Sц�Jڢ�\Ճ-��	c!��<Z+.@��l8�֭-2M��\d���6F�ʺ!)a\z���9��.�/`�����Ÿ����L��l��R�ЭW��L ,2L�UL�qp�c�Z7m�F�^/[u��4���>z�ڽ�;��RR�����GU��3c��ڻ�y��C/T+��Jyԇi:�I&�ʹ*=YSU=�����Uj2�˄��-`(ҷ{�q��bb�3[f
� ӊ��:M��y�ᵚ%�m�A��1��&fํ֨�=��X��'d�S�GY�2(��H�\uE�$P��mL�1+ɸ̹t����(ۭn���pJ�l:�2a�:����#���$U��@�Ћq�goi������U���Yj���aTɏl�7��.���hT�-�U\ Q�s2��DD)t1]F�&�"��86ë�&Tx�-XD�nm����4�]���H�xݡs!Fc�g4�	��X,*V`�z-�"P�����Sid�>E4��*Z���"����QL�oq�ۺ1��+ɺ.�	o(-���6������򒺆��2^e�.4�ʵj�cM���5%e��M�����4���Ǎlx 6�t�.�9���Q�Z쪹{ �h:Yt��Y��g��,���]29�l�Pcǹ���l��5�ʱb��S.�lP��lX�͵f^T��e���]��".Tmލ�r�2�=�����@i�V4���w��BR���j�o�ui�eRzs�p[Ѧ b����VsD�4�..��3��f�Ƽ�	��W!��eH)ZoV��T�X�ʄE�ɚ�j���A|��D���eҍ�5�3h�G1��Z1M��+QS`�f�rP��ܧ(�$І��:��n��Zim���c0���!p`̭1�P���pmf����]���M-c�;����q�7%<Z�[7��s692��LǳQ{��(�.@d�h'�h�ul���ghҎGw��cW׊�M��qX�1 �e[̽;�2�E�2e:6>�!Q*j�̵��ѓi2��ijp'�jY���Q"tl�]�yi�jhk6c�ި�owJX,B*��PVv�H=h�2�٢1fǌ�ù�^]��[��[�L���[��](հ�ї�����ܵ��4s\� �FT�lQ�VJz^ޖ��լ�Q'1�A�k�lВ�z��Yg2�M���q$)�5�2���t	`J{{x+]��Ce��z���`Zv�h�e���v��
F��E�v��(���ӧ YtV�f�ژNPD��f��d�!C;�NW�8,@j]�����N�صSi�)Q�j0E�6D�������}���Y"��tI�e�LY��/"Dt�\=d�)e��#E�B4��*�9��urX�VPX6]^ҵ�M�z��d���S9�kQ(U��g+F����4اs:��-�%�hh��Xh���bj��:�S�>C6�@���������T�+�1'I�3!���2���nd4&���ƬZ#���jN���3i%l6dR�t
��tr�*o퀐{��)+d��+	#�6�Q֘SW�p��B��Da6ȱkhO���J��we�[��e��o0�7u�
�ӉlsM�m����A[�y�]��۷�s����Z���Vd���*3�Uj�Wd����;)�;�mu�o��l!|���vv��i��J�E�!g�n�_S�܋�w����Öx��ǅD7;��ʓ��-Vx�:�&�0�&�#n�Hv�z\�k�[�Rq��+�eѫc6�m�</>FZ���g=��A�`;�B�U�.�9�^*U�0@��ʝ[C
w�Q�d�8!�(�Z�t�Ũ��s�i�{!������ښ��܀t��9D1�d�0cz�)�^w9�ɝcB���n��Ȗ+oR�7�����ܻ��P��ץ�\uwV�����R�	Jδ#A����]�G=L����p���'�F�<r3�{Ŧ���<�<�ԗ�k}>��3Kmc�w}C�o�Ã)�y+�O��ט.��ݸ�pY�҂P�'61�cʷӝL1��f�3-
��In���A��K,b�(=�t!b���f!�m�^����;7A*J�i�}�hJ�B�p���{R��4)��N<~�\1ُ�=�d�T����i�T7o-��,%G����rr*�]f�a:g���ۚ�u��Vih/�5usI��7X��f�Y'�_&��ub�NPv����M�\˛�m��W�����}�W)�w^���xq3��;T�l�-n�r/'�:��<%I��l����޴V��c�hE�$�l���ա{u��W%��2LP8��=.�����v+��O���*��:�z��2��մ���,�bR��+-��l�C���]�Ɓ��mcl��\/���ra�J'c���α~@���
y7�i#u~c���v�����3
��9ٵ�ά�z4�:i|z�P�ՠ*i7�$�Y*��� �*�Lه�>Vw�{sVL"<Oe���A�S��df��#;Wb�-h
j׷!���R�R^�L�.�Y�j���E�7*a8��+i�V[�Mؽ�1��S�'��y�i��E�w�s&�v�G̷��e�l��8hÉ��OA;�W��ds��&�1��9n�z���TԡY&�x�Q)�w��V�b��a���;�y��D�n:����0S�)�L���[�����-�4��p�[TĽ�h��V�*�Y{��
�4dﲅo]���}^O�T;��)��	z:�q�}��ܩ���>\Z�m�c�v)t����)��'Z�;-V�O�i��\�,ȥ��ɍ15�;�^�=T���&�આ�E}�)Jڕ.՜.�@U�Aл�z�h�mPv&8�U�kz�XS{�lT��1WyJ�koT��B�n�/����MӬ�':2�lޱ�jU7m�+����H?lV�(�����D+�i���YX1*k8$�7y���2.�lL��Wq��؏�uڀ�Z�����NKh�7��@�w&M�-ggQ��nZ�+���3�L_W>����oyhn��2�C����ɱ�0�����+PLoj-�Y�`�{�)>mS�� :��Ҷq�\�oV���4�Ou�����0�5v�!��ْ�����Ƿ-B�C�C8*W��V��H\p�-Qrƃ�d�g�F�Ǒ[(IJ�mL��7��e�����,�t���ӫyK�䓷W�T�;s�줊�ֹøn��x���a9 R��Isa�RVh� ҃����9�j����}����
@�>���t9��<�8bC&3� jN�!E>s{��B(hӤd�H���F+^�j���Iô�h>R*ǚ
n�I�G�V���f��8M5*𖸚tJǵi/�-�ӹ�Q�={{��~��1�5����<U��=s&�a�0��q�ˤ�e��� "O(��l��<370a)m�_v:Ǌ=8i�h���x�؀Q�"ee�KF���f��t,�)�V��,�i��˗fiS�%v�S�l6�Ҩ�1^�뼛j�iq�]��A5����eÔ�Q�g����^;֚s.G]��W94T�ڷ���g�%�$�<ك;�La�YN���ZT��Q��*Br��˓�G3]S/�=x̍�BCO���|�n��[�o̜.h��I���dy�����|�ҹM�[B�^c\����i�Si	ȅ{}��H�q��;��Us8{[ǻd5u��]H�&e o5�]gi:�JJ�Mc�A���k�82�)���gg8a
������ԅ��E�����Kܽ���d��x gu]���L���W�=���� ��G��i��e+椣Yg�vqv�y6�DX}���a�)��x*��q"��P;��^��z��k��ƥe�U����.hհ`w���g��ȟM:�K�o,޻`m$#�"4�iv��W|���}�e��X�;r��cѩ7���ܽ���F����`x八c� �� t�'!�C������M��jl��=4��?kX*�ɴ�յ[6@�
1c��ݾ�=��,�ۦ��z��|�z�$M��)4���	���Z��h'�Ǜ*J�A.S4<��][j�fZ7���V�V��]p�d���+�WM[t�2GXEv�/��	k��gSD�gm:8��իS�}�
�6ùS�QO�����-ʁu
���gH�3��S.�)��`�C7�n �|)�"'%u�ݛ��+T�A��lQ�YJ2�b�EmJ9�(��Z���hKL�D��母�7N⽱m�Q�a�L ]���w�ܿ���ΰ�\ӑ	e��'hs+�EM��WN�'�n�$���Q���BT�������ׅ�
�G�:���������o�,���%�t�w�Z�qMY�*�2��թnCޝ��t���_���zKʇh��c����fX�����cw���2Iz����P	�pYw�4�X�۽v2�s7B]�-#��tB��2�P#w��J���yDoE�es�-�]�#'M��h����%�ZT?!y���5Xȷ�msT��I)fNŻ�s�� �ջץ����cZ�^��N�@[�tv�ՙ�y�Vʾեë.}�f��%M��<�E�L�:����$ٯ��8R�R�۸OZ%�;9��N���V��rsy�l��J������ٱA�R�����Nu��9�ڕ�,zP�-i\,�C=���#�0͙nM��3�Μ��
"Y�X��������]:O��12v4^�+T)Ͷr˶��|(;-5������M�f���ԁB4���:q\/C�:S�� L]!�����-�ť:�jyK:(��Y��2�:����m�(V�v�TE_nBAB������:�^"(�u��[�L;��B����l�.b޶����&�K���܈\j\�v�h���J�'Դ��������]h���WBSV��Q�lf_3�p��m���5OB\C��$��ڗ���M���g.T�J���S!�W2<��[ǖw2˨���V�O<�g�@[��B���F¢�ot̎WR�I�t��B�����gb�[�1(G���ǑA���_fQ38��S!�\�*�9K�pe�|*P�t���ի+y��̼êr5l����ڂ�Mbsu5�%z����I��!髗�v���˖�_;�Д���F� ɴ���T�Meq���cM�(Z��i�5z飛@.�M������V:g}�`2�b�̭�*P���EC��Lڐǲj�X;	����r��g�ɋuAI
�Ӄ8��ZY���o%:��b7����\�[E�3=u
�N�yq��j1I-�A���[�æ�C ��FmF�d!��-N���7i����G&�.�-�D��O7�\�a�|��i�&k�ڭ^�ժ���P �w�s!�J,�*uD�QG����Jz���8�Ũh�(B�Ò���Ǟ��8���؀]e�lr���Ze��h��C�bq�1Q\�H�͜}��s6̍>���r+Z��h���-��:�Z	��T➈��c�k>GqP�KMw���5K�a��*@�'���t�Ut}Y�nmDzR|aז�P�L3G�Xe:��U3o��R�2��Q��Wbf���K7��C|��mmpLpzŸ+b%[۴��>}��tu�]͋6m���u�4h���:�o�j����i��UFO���o=cr�kw+`���%��NwP��I �[.�:t��N��3�X��S Y��`�}��;P-�D�l�f�.3R���0��uj�V��9�n�>ݵ�W�� oC�8_9�w:��\{ݵ�E���۩r��48Gt����-i��$�О�S��� �\�̷J�uqV�њ���97`�|�l�-,���X4�tL'I��s��;Ǧ:q>���ɖ��Ruu}b��`a�s�͕��@{���sr\a�9�(���HM66sT6��c�%W%]����6���vm��D)��R&�b���_�JR�Y��se\�,^w��fQ��m�2�����7���0�s�w�~�Ԁ��[N�i@4Ѡ�d�$�xk��*j��>��$�Xh�6n�#җQo8�"�V�F���1nMb�M4(�CR[��b��Q��u:�'OC�H�pA�7R%nP��r���[�ۨohc./���Ix�JH��T�J���Xn2�Ǹ�g0��Y�E����B-�DgT�[T+��l(�^S�V+	M�Z���z*�[��٫۟ �I�X�igz�:��i��٠�luv��:���H��Ts(���+9n��;���5DE6�<N�-G�7GT��	�K��v�,./izdʴ����f�g1"xd�["�:AA� ��Ҭ����"���T��vz��ְD��7z�س�1M�ܒIXɧ�`���X<,>��DQ��n�������\\p%n�:vKD}i��u�)<!P�e�k�׻\~�K|���й����4��Kl�/�ۄU���t�u,��j	u��|��Z�WA@�ŝt_:�Z_Mo����GV�U�Q2U�@�VFw�J�U��-J���[2�m��³j��=���dX)u��9��O&��Z�l��x�Z˻�W�u�CsS�t��	�K���Q�2�u�1u��引]L�ea�bY��s4�Ì��B��8}�H�J�f�����u���:���Y[��uoh̕`A�RK��8U�����!�ף�y*0��g74[���tv�^躵$�w�'o,
����d�P��K����9C]m����L���c_c���+_io��
�1$p�%�ǵ �G�Z��ɉ;ʐ���^^BH��u����m`q��:K�f�h��ٺ�'q��Uty�(�Rڽ4�����g!�-�)�j%>�"1�=��b�+ad�����[���ZVA��H@���U�^֦�s�j��42���}���� Y�'WNWC�fҸ�wds[�7�q��ǚ1\�=6�'9Y��`�H#/�������-�T���%:��-E�ϩ}�`�p�wr^6��.mӣ8Lh�DC���+�N4�w_S�/�m;Ur�ud橽�b9&l�󲞋����Gr���­#�6�#�-�V=� %�j5���ۦ�|�NB���j��n�k��YV�\In<��;�Ye$��_t�ʛ5R�����gN�p/�c�b�Qи�&'��v9vѧO��� ���H����&ӒXmpmRI����+T�v��;�)l<�U�Q:-�y�Xm@��d��F��-�+��丮�Վh9WV��P�u�0�a$���ᄥ�����Wa-1�[�'vݢb����MDMof�ܻ�H�����GL���Օf���#�t7�s�P��*ӝq=�Nf-Z��l;/Xk��d줎�jN�9'>�m�zDsf[�~���CP�ɻR�5аT�KA�/�_�u��e���$�Z)��17�441��OP\mtH N- �M;����<Y�:����󈥲���k�Wz�S���s;q��,wc���-స�$>��C�~�V�c�R�-�e�������Y(u(�.j�Kw�"��g�Xu�K3�2&�n�8ӛ�	XՎ:+:���wr9Mr�H�b�ά���-��R�&ݍ��sx�1Y�B]Lp�s��W48k$�+y���c��4#q���k.�:
��\mJ�:�������3���.Q*�*��;��5ǹW�7��3c�6�%n�$C��z���^��É�u��q���R��&�юX��W�RVK�Ȑ%6VTT�d"�L�t!+q{/@�rhM��߲U(�d1p���7l���V&P��D��k�Js^R�����M��;�|�����ӥ&�;���]����-�2�j*{�bT�DS�{�����d�)��)"@�j���wf�E4�c��W X`i�<Œ��hh��p�β��Aڂ�bN�ֶ�O>x�����c�\K��V��r�3�n�iV7h'�Kb�n\b��.6���?kuP����y�@��D.�u�v_eq	���2�ֆ;��Z	t3�F��7۶n�p�������}��=�Nj�����X�ǫN>	���!�j�,�w�/���J&`�
�+vgR�W���ͱN��,ڭ��`uxk"jՇ����қ�l,R}�v��N��|��$tz	ieDܛX�-+>W���\m1F��+-5�+#���[��l53�M��e�c�Ļ+td\Zr����)��T(�vv<�}�A��(Gt�Rw�f�1���2�\�}�H��e���h[|����w}:-��<��u`�����q��P����9R�Lf�	���k�� �Vܥh�8�g��ZZƛ4���9�4)��G�A��797��3]m<}K��FpM�`Yx�m��UA[�]�*Xs�@M�2K��F6�L�#"��oI���L�f�� �N+��H��Vh�*1fXr:��F��.�3�8^��Ĥ�6����UUUU�?��"+�9���:��u������7�[ױ�.�uy�����/��ɸ��d��y�f����w	;[��Mo��R��/]�=ɻ�N���t��í$v���C�ٷY@El
\��:�q�e*"����1��u+E��v߀rR��v6j3��Ӽ#�o=;�I�yD�<]`�^��+�U�J���kZ�5�ĉV�cY��Ǧ�m������7Be��2��)r�m�T�[�6�7#�2S��FX�Ю�`X�,b6��"�z�1`*��mw6�����m���xu�1:��z��T�`L�1r������gq[J2�ƚ��x:�8*�Fa�Kzݲ�ɓ�2�$v�k��۝Z'+:=�3�
ə�̆[JѰ�7�Y6\:�,&���؆ʎ�L7ʳ��ǔ����;���`.�\nc.�]`G{t;�tVj6�9Iq]�f,W�dI���m��n�2�t��Z뻪�=_��S�p,��m[�uF�pL�gtV�p���l�1�.�.��B��́՛��ADT�v�xw7:ֆ2�ބ�=�0�T���
-�ʃT�L%սA�����ur�vJ�e�,r!�i�<z_f�n0�a�4�/�R�Z�}�{]�Įw�u���01٣!��t/OV�`�]VvۡW�L���u�J����L��5v���M�ҳ]��m�PFw�w`�s��UsE٬̸xR�Y�i��T���U��2LZ"]�WTWp�5U�]v�k~u'<�5].�q]�/��E�u.����CQ3�̭}�`��]�S�1�Nڤk����|�G��Q�@�ۚ*+}]O3u�c�%^]N	��T�]�F��=�>,�nWu7E�c��ß*��&�\����i^�Sѭ,N��2kP���عY���Dj�}b�u�=z�e�9n�i�5��lL�<�g�.����,�qNb�����`U��mev�R�.�E��h�M�>b�k��n�_LzT-p�w{@U��6j�;�:��ԣN� *;�k��5aPRCQE9<a���VpS�8��{;.^��H��c֝��!q2Ro.�k���2]�:�ge�`�.=��x'f�:��v��s��5l��\�M«�s�[�Y]�����e�fiMj�,I|L:N��������{��S��h.��Mp��*Y?ih�I��9R��1\Q��\>��:�*�o_9�eq�+���Ǻ��^�*��$@����K��T����b��]��JZ
�Δ���&撽6%����A�T�ŗ��c|I\�W�3��e
Ѵ��.��U��,�^م�Ұ��|�%Y���Tf�}�u���!;�J��7z[�������N4��i�.�*U��އt��)��\���P1�=�x!��-��z\�m��|�i�P�<˗H�w^��ȭI6�_h��7*VE�F�jn��؎��7zQ�����Jl�ވ�w�%LV
*�4;x",taʏ���^���z+a9���b���W�3�ΰ`�i���!e<�S��hڐ�++��u�Ȍ�Z���2�6��guIZ)�(tۥZ��&��x+�(�Qú�M�Ś;K���v��|�/���D���Ӣ�>ʐ�Շ^k�1���V�ce�ʜ�{�IҌ��ͦ4e0܉��Jw!�E7�T6����U¢
QI0�ڶ�����:��ڗ����Au|��r�����i�;����#.Q|3!��b����ϓB�9i�X�.d�P�J�ʶuhђ]]A�U��,$@*N߷�v���aV3�β�u��3Ph��D��j�Ieh�נ-�p;NРl3L-z�*�r�����'�!o{`׹MÒ��n�:��E�
��4t��e�ή��ʽmՈ.����}��m�!�l��-��<�ޭ&�v��I�6���Kٍ�Uͷ 7�=�'o������!��kT����%!X�_D=�d�өFr�Ů��@�W���Q�a�W+[�l�VF�qV�m�;�#k�sZ�+�n㬲���Q:d�cnj��aw�R�r��Z^]<��wSQ�u�*,�'�v�AT]r��'�Qꕴ��E�֙�Y V����ƴ(�Lw,�u�ÛOD�:떥8M�!7���W��׶m�Zk�m�5�����U���o�@�Ӥ�a��X�%yY1:�Ş|M�ҥt_s̈́c9�{y���J�}عC�o5�(W<x���Ɣkgf��PHe.���F�T:H5errk�&�lc��|wl!}K �sWf
�j�P�����Z����V��Zrj8�
fGyB�����|{w�][b��E�A�`��V��"w#'���"�hl�F��:LtCB�gh2��b$��jI�-�Hn=|HX��|�Ѷ��=7�R�$3zueuԝ�z��oJf��u01������&�<%+�L��'�L݈h��Nͳ}����+�j�S��n�3{�������P= �
��{C58j.�n�F���s<n�`���(�h_`�����1���u�nP�^
��^����uu� �Hw`���ڛww����kn;*@���j�c]��	�����>O�����z�A�XegL��fСV�{��PT9�IY�}Y�x�N�,����O����o�hhL5���vkrd�-JV·������Q�ךԡ�o��(���.]Ps�t�J�Qt�\[H��SH�A��@aӁ��W�q�.�M,��x�_)�I�<皲i��J�� 50:K`95FnG}/�r�0�Nbj��$�O1���sR��	Џ��c4��m��XQ-}��#f�-�9�+k57��G(�*}j��֮��"��f�,����90K�:�6U����#��G�nTւ&���s7�]�MD*5�sj��*Պ��Ǒ��	vh^Q�u �ui�Lͼ�v𐓗m�wr�u{���yz����z�W0����s.ŕ,�V;��F�x
�B���*ņ&��0��J��i^-�v��DMU�������J}c*�RZ^��L��G]L�x�Q�������p����U-�#}wƷ(��h���u�0�7d�Hx���]=<��m*9B��O/G��wF��5��z�H5��New3��PU{�eĮl�X���ݙ (i�f�Y��\��B�����Y�
<�ڮ�����n4˕��'J qu���}��Z���j�ۅ�h�G/wzt���O�z5��&�J�����(�#��qu�ԀSc�P�D�	�bC���Y���f.���P��d��`�E��Wb�r�Q��a:�u���le�j���Z���FE]Y����4K�9/f]��5�)�@b����w6q������z��̀k����魔;ffN�^��	B�����Q��s�s���δ5��mk�	¾�:��]�e�z;^�5��xc�XٵX"}:�v>�1�k�tK���n�� Zʴ��ҫ��%2R�U�GM=+.���\�wb���(k!ض��M�p�o�"S�T��c��ɓ1�Ƶ4�*���Z���k�N�]#��Rۛȴ��O6]8% �=���S�)!.�z���ۣ�gp��d&pF����7:ۼB���A����*d�# s.�.��kE��w1P0�ŀb��¶���y��nӧ	�V�f�ȃ�}���vp�ϴv
�;n�4���%��l��%�ڕ���5�He���P�n�!�U��]ɦ���۲�ɮ�pj�}�b��W:8�w���4\�m��kP����iް�jz�7vV��bh|JW�ގ���Ue����^�)N2㶡�,@ϻ�8;L&eR�6㗸��a�ns�!�ֹ��\���-��m[����V��U�y`�B���y3i孹s�A�����Bu8Z��V]�4�P�yP�p9Xg�{Fu�[m6����y�Q�ks\����w;�$����d�N� #�o�[c��k�R�kG|��}Y��単�ƕ	���]"�
�e;�]��iCtP
yV.�^bAf����+m�9>U�Y����Nqu(j��q�aM�o�.9j� >��.6q�w�o,�sp:Kp
o/c�v��1 ����R���T����5����� vۧ j�Y�hJ)̫�L��+��_p*��t.8B+;����ୁJ��SzIm��_��ܥ�I{�E��Z"��U�u�u�b��RWS�����H�Y㭸K�"h=�w}d �,%R��n,/DbN9r�I���`�-��O[�����ê�Wŧa�Sxp-D��7*�P�9ٻg���iq�MP���6
	·�wLܤ[8���l�o�ivU�iq�-lj��X�F�t�F3�����홗��9�L�6�V��]B�3��t��D��S��U��@F�)��1�W����k�ʶ�������cZ�iΛ���mt��̙�E=a�6n�,��Dh����id���hf�Ҙ���hǙ�������'��m^Ά1d���z����7���G-��);�-^�9��n����ޜ����먎Q��xV<Kq�Ju��wۍ�C���0�=ox��L�/���f�7)��u���B�9��9X��-�4�35���X;4�d�K"���YԶ�9���PZ�]�����&��r�2�I;�V�����ֹ��"��f����Su�2�1�/o�m3��E'^EQ*����/)dv�y>w3R��2�=Ѱ\�B7$z�q�9�FR�HK;J�F	QW��uvlf�i¶����'
˘�(g\f��k�*�qi$#s	�Gm�9�h%q�;_RfQɗf�2Wcr�YӠTM�T����V�t�(������q��|l�.�5�'5��d�˺e�;0-;�Z��zp�NF֊�`-� ��ˇ���s�7����I���P�۠�M�՘�@�K�㮠�t�������43���u���z$2*�Lr\']������RS�|HDt�;=� �Z�f�� ���sE���ES4��yBx����Sy9�7�����ˮ��8��Ko�B/,u��
��g0�0���@���b*V�t���L
��4*mn��K�G�=�.z*X��4����zv�X���og��u(kȺ��]���8L'����T]��M�跻$�E���Tl�I�Re��fK����4x�I�������A�u:���-���g��!|�n'��t��_Uݰ4��,�e�y�2HN�[�� ��v��(ndݠƬ��KI��{w���X2j���Vf��ѫ��Ɩ��iv:��)�Ʒ9�k��yJ�u/�-юܫ�I�y��Yz���N�B�4�S�����/����{LJ
5��X���X0�r57��n��|����֞�k���%����)�J�4t�6��*��ޫ������p������(\W����+�f��V�WTv�h����N_s�q
�.��=H������q��Ap�F�]ݿ��,K@*`��]�Xݱ}�d��{a���%[���n��\��pw;��ȶ� .�n�/Hx�Y˺N�f��	�Ry�g +��C
�-z�Q�/$�s%��0�:�^���+^1��19�p,[���][]W�	.v�Bw!r����,r�2�� !�Fe�i��}�>}�syڵ�6�NX�Z�=3�����\�lF���vH�-	Iot���4�n�Y�'hz�#��V�c�N�]�f��aiוj���WB��-�]�j�*q��pԱ,Õ����$��Rss�����P�5$��cj-� �Y�D�u:���+V��{c�\EE��7u��洝��=v���X�&�H�e�Ϫm�/QK.��v[*�6�8&CP�ŗM�;Z�ڲim�����F�.���fu���Il��{V��lڹ�KN�J^��ۇ`��®���tt�{��#�MD��tVR���[4�]��������a���|3�Q�CAǏ2��_rr�u�0���T�H"M�=n�T��>�Y'���lab�RQ�SM���������Z끻�-q�Φ)��V^�PNdv�H[�+]b��9&��IZ1^ �֬G���7x�q�]�v,�b���nay��0 FV�R��P �Ћoi@��K�]�SnW�ʀԕ�"�	cv����G:��t;:�c�;ǡ2��O�"���?6t�t�ؚ���XUi"[�aT����N������cE�I{2�o[�^t��=��}�jrԷf�苝R̳��N�^��1I���7��}=yh�"�����t]M�Ė����z����ʸSQ-[�C�Nd�,�{v�2	�BPi�E�Ӵ�o.@���]�ucYWQU��)�U���r�9DD�{)��b�T̰ͫ�wg�~ֻ	��ڹV��<R��p�wg��Y}�f����z0��!��{�:]V0�jLmb�ۊ��ނ��t�RT#�F�B�X����!V��dj5N�zw�;�r�M㾀�����S��%t)�i:��n�Z��-Z+�]Me�ͻ�� Zl6�%;f���7�mo�6lgJ�j ʭP���y�khٵY�� ݻY�t}zCDu�4�c�'Q�.��˩,n��w�t]
�w��N��SS�tN�Y�v�s�j=��� ���;FX�@֛�˔�������H��9���K]Cf�(X-�ޜ���,���'|y�V��H�0r��%��bVQ|yJI��cVR�p4l��<WR�b�z]'t��2�톐`.7x^r���(Җ)k�r��OC.��Y]�{����wx��H���hH6�D,<6�DF���q7YX{+8:A4�:�w��W��C�I�W��SR�WE�zty	��tՕK��^��#�F0M&oy��[:��~������{�>�]�=�|-x_�Sg��f�t϶�˻��,����!]��r�}M��+��_��l�f��;���0��&͖Tɐ����T�u5p7@1찞�����+nd��'>�z7e�����*6��K���mH\�m�iؼa�^|~TL��=+��3/�"�e2!�n�Sk�ݷEդ��#���Ӳ�%�"Vn��hю��*��΋qG����O��J����GJ�/,B���Ai�&��N���̰U�cZ�+byӊ�n�0Mie��f�RV{��lvC�ѐR�+[�hK�&�of�LUb��ʾ.LиGR��q*�HFb��q�Uٷ5��Nֵ	؞A���Λ��f�w��!�S�M�x�*���T�T4�k�y��w-�%��>������A�Su o���!�t�� �5������C�� K9}f����"�$`Wi?���b��9qƮ�*�yIY ru�Mm_v��̍���n�O7�@VՉ����4n�_�c���������_uG����3YQ<Vj��+Ă]���Gn��x�ɢ�E*�W�o���v�8�.����C�Ru�T38�R���3�3C��e>�&��ź����ػ�=�]K�F��;��W%�LŴs�/cv�jǡ�N^R�!
�)���;����+�tHͽ��M��g��\<8!L��B���%�[T���������(���Z���,����bc,J��"�j*����h&`��&h��"(�����h��&
���h�h���"��*(*h����*k,()�"j)j`���"*a��j���*�����("��`�*�)���b�B���
��i��Ț"����&�*#033
��0ɪ2�"�j�3&"0̦�*�*	���(j��������p���
�0,q����2�,�������11j���$�(����j�"j����!���X�j*""*b*��(("���*���)���!�����`���(��"`�**�f��������j�2L�*���"�)���h��B��
h)���ff��(
"��$��fj)�h
J���^����U�����+�&�hU�m���2t�1>	6��u+`��|�9kGvw$�ޱh�`C���3�8��V5SP�Śr�;�^R�oP-}~�uZZ�;�4hn(��+�kn�sQ��R*,�@������:�e^�V&%��4�#�@��,��{[����ޘ�1�bv[�bMAKt��������� ���@�����DI���k�؋�k�	uMv��%��7���4wff�9Mi�:���;���L=1���官��Q"~Nbģz�!��6�vl�"g;��mtԬ�R~q.Y9q��MgvB��}$�Y|e���c�ƠP�v��3�G����L]��`����*��9�Ea`M�_�M<��c�N��7�+�Yy]YkM��k�����.,�=��B���ƾ� >��� E@�@��\�ּ�!N܂�lOJ9X�;��p�-!c�7��%�C��$�#�YZ�h״��4M��:� d<�Gv�}�"�>T�h��%p��t��'G��s�j��' ��u�M!��c��V$�Y�S���WF��hˋjޜJK/ND��jဍ��l�n�TN �j�a�k9;̘����ۍ�U�B�Zr��b�����mh
~����_�
��q=9��}Îz���Q���1r�_^�كh5IP��5���q2���:hY�D��ٳzU���闥9Ǵ��oH��p�t�q��E�V�#f�3��B�w1$Ţ��}4�0[Z�#�Iү����RuC��9E��Yeg�U�ɗ���_5��@� 87:�j���P����B���q7]��?9.f��ɬ��7U%i%K��	D�TA1��{j Cbj�g'���Lu<����US��~����?Uy�JvPCC�@~��$a��g��*����N�{�����w�y)��gj�S4��քB(�;���t���_���?t״�7���9a�!�Jw��i�)��U))L�-�Z�
�����Vt�,F�4X�R�y���F>�_�l��4��ڙ��ɋ�?2j>N\	ۆ���Tp�Q��j���al����z�A[}��pTS�f.4��r��7���}��S�]g��`u���5���=鎑̼\��%G���aɎ�+��A���+�j�������tX~z|��#���P::^�}��r��^B����ncD�d��L ����S0��>~�X�I�u�G�S��v9�'�u�`&��ԧ�s�6}���V�B�^��3f�@;[�[?��ʛ�8]u�Y�ní�Y��d�X]e.��[��VI:o3��&������#�n�+M��}
�\�U���f�����o�[ӘDk��a.!gJ=xu�����w�{�K���d��^x�V��t�B�u���*���P����Ǜ���n.Q9V�����p_VC�k}3¦_�u���<gD������u�R�`�٫+�VQ�k{yeb��Th����07��ˢ�L�v������>Y�0\J@��t̩�{����sDPs;Z/�i�,��ᮘ���t�3��M\>�*��N@\vջ����1��Y&{��=��\'�Ox�f��X�pЖ�_�d���8*�Ķ{�ge?�f?�7����"
�e*��ݚd�Ng��?}�fCN���q�{�$Fک*�]�qx.�.;f �2�n���D ����*��'��UyQ���f�d�2�Y��C[֢wmq)���s����F� %���h~u�"_r(�Ts�n��7���r5�]ms1���<OJ� u�9⇒T��R#��;z��n�8l�P�r�p�D��+
�]�D;S¤�BI�g"��hLT'"���-6hR�npȥ¨\�,��l|5��������f'R'��c�L"�����H�6�=�ˬ�4�@��N�쾭ǡ軶D�X�9�b���;{��tTA�iNJh[�Rr��QL��{'��Z��%o2�S3�n^�1t��w�ۛqBi�X��{�}'}ޱ�G�U-�=��!����.9+�!L�Br��@��/Y�nY�1XS�{�ӽz�z���Gi���Yǌ�>g�{/v�o9�]k��U)�8�#n�[�w\�%4"�(ʑ�'�Pzx��)�xP�c!����rMP�=랐�'��|4����b��1\������D�_�����Q���t��'�z�����+��=ܠ�C�{p�L� ),k6�W�kk�f�p�N��2����R��"�MO[͛ݽJ2T��C�(��쎗\��N�+~5f7m��+_���]mԞ�oN��#kͷ}S��=�+��LSZ�����φu��[<�,�yC���A��?'�s}@Hg�~���1�,P<~�(�|.�^�mH�mPAg�[���-=�mFZ���AU��8�?g�<5����{`��`>0�"��o�c��r~��l��� t�N�ש���)���zV����|���U� r�8�L5g�d��"x��{.l�,�������=�b�`W o(iluhq��GK�51T�[7�Ӧ����P��}��[^����ukxgg���j�-VR����7]}"�es�&��\z�W\ld�ԋ�P`������PJܡ�5����qq�RU���wai�@�vݑ���:$EB�8��n��r�V�-r=�y��}�������և���~�����h�x�'U2�*�$x>�w[��I�ð-����Z vdДc��Xꎝ*I�c�����M6��sn��}�1�=2�9��[�Z�!�� A�:�����d��;z�B�G���m�� 9`s�[FB��˹H���Û�}X>���F㌒�:�*=�t�z�QW]�=_w��;����q�盝�~���G��^`SC.�0'��P��ƾ��a�unHv �T�N�졽�����HU�k�ޜ��&�b F�uC.5�ٛZ0��B/��8 Bj����/D2G�J���ht�4N�����zai��⹙^��Lt�x�����tk�W$��)���N,��{�C�1����x�	��)UX>�Iֳ��i�[��L^������<d�`�_^�5Wi����𪹬7�)`���|�i������H^�J���*��*=ל�����ސ]��6Df�ʚ%*�ْ��(����q`\���w�u�዁�y)�[»y���b��w��ww�	�1%ց�&��	�#�����o�-##�Yyk��˂�݂dƄ[8�T�h�c�En�G��D	�kuJh8���LвVl��#�ƾ� >���P1'yW75��pEF��|���]N'�Z�gު��{�� ��	���]|ǥ[�z"~��YP�]����U����R9��p8F���LÕ,g}+/���WQ���O�X}P��Gg�\3�!���*��P�"&����v�zr��ӑD1���b੶^��D� �:�M���Q&�9�����1u3V��E,5���jN�y<>�N��w�(�X�z��Y�d�˲�<T�p�������Q��E���B���7]���]��֭���M2��R���&�O3ъ}L]_ʄ��JT|L`j-�ۀ�I�C!��3˥�����T��C�Yi.;����S�}���.���w��*��%C�Z��f�-A�N|Ҽ4�M������n�+ :��E�ݰmUc��Witq|��?t״�=�G�|��%�f����t�a�B~'�))L�7�}(y�j����Ǟ�mxS���U8�^P��(^v����[��oϨ��<n ޣu�Ap�¤%�t�-
$i��U3�����k�Գ�y� �eZ֏����Ϧ�w����*d+��i�#�@�t4���{��:w8�ꉉ�Y��޹|f	Wq���Wf9��cD�BCKK���+ij�g�8�\d�5ח����Ȗ��������8@�?ԱwTNS8�:=��U�૆:5���|��_�xGF3a��}���(y0��u�i�C�v��/c2gQ�f4ǳ�*�U�s��|a�2�b�.���(�)K�#t��gu.b�M'8\ܗG���y��h۟i�35�!�_*,ԵDo��F��1��إpV�={��F*�iUah���p�n8�c����E�Y\/�ы��\d�
�U�����B����-E	4�J��u�D�s@u�� LFk�D?!�
X��n�
ƫh�ȼ��(�.	ЂEE���X���g*S�@b�L1�1�
�@���r�X�_��)�,���Jw�nWK;J�O9�܎q Ȏ2��Os��Y4!\@�L}oC�1��|��}�V#�n�7j,)��齕8ڋ��48g	.����S0�'�=�b�/�R����b�{%�׋�d;^Q	��5�_R�,1�E�i��6�NX�VhHnχ� ��u�#��Fd4�c~�.ΫX�u��e�)��*��
a*�W�e<.�Ά�͸�&�8��Ɣ'^N������5L��b˕�#��Y{|�HV㬴v��KR�ʤ{X��M�0�M���r���iob����6a��9���j���t�MݽA針.��Kq=�a�����Q�`�4�n��@ ���BCV}k'��������b��� ���G����]��t��3�9v�m�u^�b��H�Z=��(���]k]Qf�߼ן�^��f�˞��2�;��h㙎��\�%16��3"�7Hi$v��]�~��ݑs[�i����( ��aL�v��O
��vYS�\:�b��0�O+�)'e��26U����h�~�ك�1c"T�5pa��1�UH�	��k��Q5�6l�]�Z,��o�'3������YGn���~��B�
��| bݮY�{t�ʝ�G�/;dq\�a��<���SB+�eH�ē��6���+������Ҽ�'���fn�������z�xA'���_�j�������%�\�:���XD�{��z^�n��RJ�-�7�p�:��2Kˮ�_c�S�߮AYo�GD�˷SeP��6:1�~�vNNC���Y:>��Y��S��ߍY���8�F��<Dˊڋ$[�ǑZ6�YY�&:�f�1���K�|K�cec������B��s���mo�����Q�@����:��I�xz̨�noECY.�D�U�v���u��0ic���dCL�{;EA��M-]����ͺ��pUiS�IW�k���-��D�@uԝ+.����V�
���
��g]_B��X��r�N�����3����.�[��%�T��0p�q���_D[j�>��|1{�-����,���H�����Ĭ��Q�G�<|��أ)%�G�\����(*-g6f��{����rQ���@=6��ȗ���l��T���L�!����V��B��|�K��T{��n(z��S.9��n��wV�Ȁ����� 2_��rf+��k���[7P�@��1��C�t��3�J�˥��F?6��In�x����p�[=�_@9�?����0�_���:>T��e�,�c&����}�XeD}I��]�R^�Q����n�"=��@V�E�K"���dpCY���eN%��U:��U�9qy��3�!t�����qk�:�@��CZ�{^3uLׄN���=/�������[�G�WC�ǹQqa�*��Ƚ���	�uJ���0�}][�B���=�0}�b)|�P˫βo�f|�ҒBƝ�~���K6��}ﳶ���v�K^��cPn����eD���[[o�|팇��k�(:Z����Q`���k/���d�/.��CI�{fT�mZ��S��w��hM�۔W�O�:l{2�+�m��]͢:�����o��۬(��&����Pˍt6f� Gg�*�~�A}�|gG��{����^����zy�/o/�ޘzc��T>�b��F�xӳ��x�6a5�$K�X%*�&���k�����|U9��C"UV�'Z�>�g�:�0�Iy%�Ϩx?>ywy�|�3�4����n��p�>^8xW�z��~�J�7�f;��ʾ�w�j.l��#沐�Ժ��8Jۃ?XDu�'�R�X�`��"օmN���m�����y�R�X�i\���pѸ��Սm�싞$0.A���_0n�[�7v��~5m��U\�w7b��
�`����Lź��]����"��v gي�=3Rʕ��~۫i��Q9^�2�׈�^�1,�-v��RYzph�6�5p��6ϥX��EtF�x��P���~��<�1$�#����R�-�v��jN���ש�1h����"b�J��ʇKp��C�����c�ʱR���g�M@B7�֊�_��6��n��}_; ��� ac]zZks��}wj�^E�'j�O|kB�&�R[�@U�A���Ĝ���k�p|�op�R�x�`���L��%�f��K������gn�R�����O�ǡ�{N�́%��po)1y��4�K� �(���HEu�d���1ns���Ԉ���v�8�!:���b$'�ˇU�ǖ��K��RV�5<��a�s��Y�h���u���M������t�(Di%~U���\覆�;}S&���I��P��ǖ�wE+r�t���kb���VrZ}K��,5R��\��P,��k3-P���U��$��u43ъ��E7竵"#'��C���P��	C�����[] c��,0��j�8�s�ޭ�Z�7lr��:�:�'ө�T�5b���x�{}��k7�q�G-��Z���C���Xt�׸��TP�ᇀm;���#N�S��6�7n�ZX�X�D�{��.�kX�ji�J �*NpW��Zu�䬒^m�@�d
�9"��4��&���s5�T��\\��s�mHGh��d��|���L_n$`}z6vG&{[�%��B��9e5��E,}�/��j&V)�P$�߳D*�����6��bȭ�Ž���l4�ld�'n�ntj��l�ٻ�{�:�h���|���l�6ݝuC;i>KW1�`L����T�p�
GFP
��{Υj2��Z1���sbݫ�Q��}u���E+"��	WA�K�%��ś��+���k6�wD*C)�f�d=�2⼧�mA�&J�Ŕ�q����("J�L]8Z���u����㎈y�8���E�"��s����`;���k�X�bm��˺����JM-����nʘ�Z�>ةs�#o:��G�7$�Y�	SvJ=Y�#��"�܉��jd�6d��x��R>�ŝJY�D�G��tS4��לhU�sv�7�O���F7���X��,i�k�X�46Y���u!���:�,�	�xl�)V�N�����W�A�W�$�u�:���Η��n��!�qtA�%�9��^:�0��W9e>e��$U���g��T��a��vޑ�&K�u��|�UFh�B�;Z������^�F�i��f�*H�)T�:C�������)�-���V9 �X�
J��J��-�i�Zw�f���&��`�ߞӈ�7l���Ç]�������;e�m���p�)��}[��L�Jvw y�b���q���GAx��,o-]����Gq�����t�]�<�V&�$"���vεy6,��VH�軄:�vZ��A;�,8��)�<i����d�7>f*T[����x̤{�T\�H�؈���ʝ��#�z�cp�+O���]zrS�H�ҍ��4�uQ�w��u0��w�c+�Ny1��v�<�!��*�#Wj��D�I��!e&ֶ�t |�$^��*ᛆ�h��^�4�%�������]/�#�����E�TEDL�IEPTUQ��)�`���&(�*�����"�J�"�� ���J)��&`�i��h)j�
�����������j���(����ih��*��%ij����)����*�&b���H�*���J��Jj�")b
Z����bh��������&"����H�"&��%���&��b�����R��j�����	����'#**(���������������(����bj���R�)J(�������
��������h�Z��%�*��$&����*

�����(�"Z)��$h

)��&��������&�
��$�������(��h��*���*
*f����MP 
�U ��˝L�nE/vN����{%^������*bj�	���R�*s�z#o"�-`c#_v�4D&�f:.s�9_>TЏ������=��rr5��ZN���%Q︚�G�jA��NOװs0�FK���b�# ���?K�`��P�0�_|�t����>������"!�����m���b�g<��D1^���C�sNC�~�Q��y�Bu>K��u���?BS�w��3x�r2��TY=�Ւ����9��n=���>����{&��|�P�_xG�\*�����53K9�T����#蹁�7��F�Կ}�����sX��>�PFO��.��C�;9�����L�A�s�=G�~��	vX�\�y���$�HRe��7��XZ��R�g�e����R����",}""��5|}�j|����{�6�BU'O9�èwHs��`��V���ؼ�ɒdyr���� ���zj��rw����ϳ�}���gr���}y�
�&�
w�uҧ�_g���}��_������:���y?]C���ػ�C�:}�����Jy'��GRu;�BWkKE#Pj~9��bӓ������:�������u�PGF�>�宷�퉬���ܽ }�x{�.��O��u?��F���Or�~:��7~���A� ˹|5��������t�^��Jy϶�f.Z����h7P����\7�]5gw&6���=W˂��G��!	�w��:���sS�Ԛ��|f�p�O�tfj�'�5	s��p��캃�09?��c�������\��[܅ ���[��ט&N�~6���Äw�sv��&�т��!B�ѹ�\�w���'�7R���{����?`����A��ѸJy��Ӭ>�����xw��C��5��j5{f��d�&;6bti�ފ�NK��ح$�}��# ��:��\�2�9�4C���}���?����}�'s��\�����u�/S�����:�pgy��!��?�OZ�s�u	O��X}I������K�t���{����
�@� ��j���ش��tf���FK��~����.�2��k�J���v�z��K�O}��'���<��S��;��v��5QӬ]Cʨ�*��W���m'��Q�x���0ֳ�,Ο�z��n���Y��N,�b�0�M�a�����A�i��,�o�f��w�]	����'VKm=�r�p�U��bwT��`gn��qJs�A�z>Q�yC.Vʖ6[�zv���4,��ѝݪ�����no:2�Q�IPݐJ��t�����G�>��f�?}�E8J�}.�/c'�_�����}?sA�K1=�7���MG����!��}&����c�J����.��Ht��o�n>�Q(����oy��[���{�>��~���&K���S�;�fc��m������Hr/a��R��~�א\����<����	@��h������紒���
����<��g�9����A�C�2�pu���j��c�#$�6�}{.�9�a�wrC$��n��9�}/㟹���.@u�ε��rK��󟠈��c���+��f��+��w7�ϼ��5�|���jG�as��=ھ9�s�w	O���h<����5E����n������!�# ��?N��Խ����S��������19ۈ?J����;�v����O%�>�������j|��a���K�k��&��2�oI�g0L��\�A�X����v�S��b���fb��A���P�`�?p����H�#�D���u��{ǵ��ۄ���MG�sC�u	A����~��~`d5�r]~~���:������^�7>G�bo�!�s�n7.�s˯p�]ơ���X����>��Nϗ{~����v��Y���>�!��?���>�?g�1O�{:�����#P��G9����9�����}�!���������j�}����2L�}���}.�:�����P�P� ��5pU��f)�#;c8r�˽����9������{� 5�%�rw._���3�_ө����y?Z����vk��=�߻�:�ơ+�Ò}I��55��pPy]�Zz��?|O�4;��ZN�ns�K��_���!�FG��w;��b�O���p��Nc�0{�P�[��%���=���n>����2J��r���:����{�m{���d��K����?g�����ݝn�]s�����\�\�^fj����1.�7	fǼ�~��F��{'fgq�Jy��oG���BQӼ>�w�?A�;:��02�<��0����\�ﭽ˸FO�w�9�:�Z�Vu�f����~�����6�;ka�Y��K�Q٦~kg�W���$^�q/pMSt�<A�N��,���{�H��[l\�/�Uu5̼��2�E���.o/��횁����К�̭�2�%;�ʼ��4Wk�f�P�����8a�=������뙒?�6FK���߷�����;��v�����.T����reI�����j5�u���L���u� �:���gX����<�K�ʓ�pg^f}�}�\�������˱J�h�>�f>�"=�\>�ђ~��i���.�;�>��W؆vy�����=���Or�<��d��������3X��Uִ��}��".$ƈ��A1�R�!3ևK^����}�4�}�>�!>���x}�����0T�Pk}���;�����[���r@dg������]Gg>��BUG<��x?A�s�����s���n5/�S�Z�]���k��>������=�^�;�������HP�=����k�	�a�K����7o�:������:߱��@{���}�P�a�δ�]�#�5�5֞�P�}��T�ߗ�V���!_P�	�:��s���������}�>"�ЄD��O���k��:5��FOrQ���u�e��]o2B�7� �d���f~�nz�#�}�g��p��u�7���5'�eO篴;���jO3þvy���L�&kf��~������B=�ԁ�>�BQ�3�~��r{���5Rd��cB\��f��p����rn>��Rv��#pd9\��n��r�zg�m~����?��o\��e�+��_�L>��jF��":�h����Q�{�_#|ΪB�����I���2yY�ݒjy��c��MF���e�J������5	s����yr@vu������������|ߝ�xq���UJ=�7="D} ��:����5��7�>�U>I��7�����^�y��z��e�����HP���h7~�Q�b���K�����u�S치3^�BU���Z��<��z���P����D��=5_v���MG�~�c�w	OQ��Q�=Ơ<9����'�k�y���`d5�u��m{��d����A�x�]@s��3>���I.��5��N��^��L�ݯ. c�-� �3�,B�=��<t�𽗇�����Q;n�١Br6���j�pD�mg�����j�>+��#����b��i!ѭcH/��jԙV�n뀻--m+rZe>W����v��x���r��jQ?]sc%����:�.׎d�_m�{���-�+Q�"v� n�vuu�Ї(e��F�:M����	?���K�;=�[�]�)�V�]4Z�l����١(���W�:>T��e�,�c&�,�^�����M��{��I�"����1 A�:����_d���޲�G��9C��}�\��Z�{3���U"���鏑�ts�2K����v��F<"up��Uܗ��{�"�Ʃ������Vܪ��"�9`iyM(��uJ�~|h��w�un����	���v�q�W�5G��	ݺ���w�#S�����uC5�ɚ:�f5�
�7s[�'W���{�<�cX�5{y^����N��}T�,ډ�Ńè��)P=VT<����,�RvG`V�p����SO���..|�W	K���Nq���y.̨5��%f�3j$���cz��p�3gDv��.(dU�a�X#c
o��"㩧�6�������F�����Z���|�sq۪_G�z�g�Lp`�إ >�L�]�ة��s3`�c��a�U��;�#WΫ����-���o������
����x"O�kي#6���ڱ��p�fwn(��������y���=L�,v�I�ߊz2;c-j�-m=-�9Q6�eq$���]ݘŗۏ�U+K(��}\#:�eڴ��Q�4 P{B�a%Qoi	8h�I��e�ٰ��ɚ[�yN��T�B2���k���uc��<;"8��`����lÕ,g}+/��E�[D; 0���
,�H���N
/�nE�#8��fщFk�ޜjK/N@�jj���2���(�ޢe�;[��y��2t	��_ژ���f��j��R��K��p�eD�ӧ9�V��+�܎���,�A�� B T�}5�@(D���E�K��m�DFP�ʵ��%��9;KI{�q<nR��!9��" 5P$�J��&05�ݷ !��C�<vlŖ�n��(yݎ+�W�i3�,���ռ��"B� \h��~)�Q������A�S�o��<�7��S�Pz��넪5��^Z"ы~N킦m��-<v~��v2{Wh�r1�IW�;WI���8�ѽ/Mw!_%�!#̙.!�@s�6�O�9�맇�	`�'u�C"�ut[½B	yt?].�����u�ΪL?��̚��������yr�l��*�����@����B*쿂�<�t0:}8�\F�2�Q����O�3S�[Ь;�ف=~=]���7���⏓��S e�!����^\��ohr�*���zu�S�Fr�h�\�z���m)��
�n��7j-N�&#rsu��CK��qwL��+l,�*Iʖ�(Z�:�;��b���Lv�7�:wA�Ң�sYع�}Ujz��{��������`}��� k��V$���8@d\<3%��z%��{7��o��aH�.9R�9M�7�k��.FgN����T=���fZ�7�ib�V������l��( �����`qA�}3��n�W�-���,B�p�K�s��[�;��9�t/�^9�<��ӉU�T� 'y�22%W�m�b3[�C���ǂZ�DG��ïOo�Q�����ubg�\T�S��cxb�ҁeѴ�2�*�:
�΀���S�F,���邗d�=_�h\	ա#�R���B��L}qC�3�ge
;N�H@i�)R���z�=��k���t�̬U�</�pi-�]:`c�b�LvU��R3o�$%�k��a�Σ���-'��}��l ��p\��'�os�j��tM���w�0�U8�w.�>;�'@j7� �sA	Nf\�  ��>�`�P'gaS�	t��s��munu��1Ȭݯ��Is:!��M������JbIB������&E��IOwBF�gVS-�fQfDکj��KB�(��L�,�o���̏���΍�(�z���q,�	 a ��N���ϝ-�GJ��ѭǪ�+�1E�v5	o���0R�u�so�'v��\�9���6��J�T�*��2������7~'=|�����a���)�2��4U	u�Y1���2T�.�w��W�ȴ�	���פ�׹�}�bCS$>��b��0����a���z�Aq�1��vYϠ��ֺ�RY����vn�l>E�����@�tw�R~���b��R�����?�n�{�7�5D��kͦ��ޓ;Np�O�3�w���ڬ�EV��F�l�mc�T|s�!��!�E�mu�z��8�zg9���p��ջ��>�+�N�i_/��s�������6;�
r^�o��F�ٳC٪����hڿp~��z�U�I�Ž�b��X�O*$g�t�k+oM:���������9^�3����zbD�ۅ��5ȁ�X�o��ճl�3hE��[��̙��oM��K�:_kJق�~CڰpT��}��3�;L�5f7E;�]:M,�6]@uTr�ע���⼃��˱�At�TD�������
[<��[���V�zt2p��e��j�׽ѭ;f��G�Ҫ�����7O��&��Q���o���\4n๸�]�Ni�[�沟3J��#pD�ϖ�$����-л�y��<)m�{��t��lP�B-���.�'^W��j����[J*2���B�m���'�t�#�mFΗr�Pi��B/!6�y���L�*`��U}B*	�����Y�cڄ�=�g�����epY ��`hg�_�T�
��r�)�E��b�_�mAH�Y5w��i��M���/+�Ѧp�) r���d�ѱ�m�F�z5>U����� ��ߖ-��Q�;	L0��k�#�۲2�գ��`"��y+���/ԍ�M]����D	p!i��u��tه ���ٌ��N��.��\�z�p5��8���4��f��0-��)�2�ӣ�_BN�A���x�gGP��������@}T��Q�͛F`ψd����#�ĸ��}��B0�VWj��q��)y��D�#��钡��DX�1�D)�tn#�������][F��d�0�Fγ[i-.��F�{�-�����健�2/`��c�C���~|j͇�{F�m��@mȸ�-�kp{�' �T�[�W�o�é�LZ F%2-롳7q�#��ӿ)
~�KW�xv)�����:Z��M{	�zy�ں�x����_L�\�6�A�*#�&�z�`���L���/a�TL,��05�t�bͱ���^YP��8Z{0�顁��0�� j�9�t���{gyV$}.h��}�"�ń�U�:�y��ls�Q��B��1�$�z(h�d�����8��i���%A��f:���8y�sI��Alr=O���;gB���DG�vk��X�K���4}���?�֍T"��槏Η(L�����pڕU��Iֳ�7{����e,�l���m?���o�B ���W5��KTa@O������h�G��'+���Go��UQ��|�}�y���ֺ�Ѐ���h3S��x]�3 ̳����H�J�rf�$@{ι��r�l��v�u}��}�d0�c>��t��d�&����ޅj'��1���S8��A;�;��\C�LnD���d�[�X/xz�\)h5�c�א>�}NR�/j�L�Q'�2�ec��q(�/�ڄ���Sl�iTrqGn�QΛ�ފ��<[� �'@�x�RSLs;�_MB��pֻH�5'J��:ܧ[�D�ڽ��_���]GzG���*3�O�� <�kAB;�Rڈ6Doa�}�;������Ľ������?bs����JTA1��0�N�x�-�+�HZ�C�ݠ�O31�	�mցp�E_�D�+� ��Q#
��z�:ߩT+�|�wA�������*���ؼ��k����@�/.���&Vz-ׅA72����D�㕡-=��0xue<^�8���b�ѩ,�(]M�VV������oV�1���!�O�GG��J9W1�n[�ni��K��XE�oͭ6�������D��5��-��]�?11٢��%Pɦ�p/>�0B@d'v���U���u��c�tF��x'�(����|"�u)��iZk���.�	Jdɸm��C� �|�u��(�t�4]j홳�ˆ�^���N�`�����]�����˅�rwrb��̚N\	ܸ=�Χ����^����n�PS�tk�G�FY�9ѯC��x��3c��l�h��<i���Z�n�y%ؿUFk����K��Ơ�^� ������
�H״��G��r����a�nH�]�
o�ob�W��������S�-:{�ͦ��	0�b�QfZ�0=�}���K:�n�PR۲y�0c�c~�U(1�����Y\/�ыG	���1��0����Ԁ{���Q�)Uq���p7�@	��\��U�jX����B���<.�rҎ(��[���u���&�x�D������b������F�9L��j�ۆ�.������Z�Z�@�����aؖ��ԵY���&_)ȅ�B�t���:c��ҝK��ʽ�:D1�w]���q���f��{y&�|���:�l`���{n r�ʮ��
�-S��]TR^�9%i]C���)a���>�[�+���7��n��k��K��Qѵ�f״9������.���5�>Դ���٪I<�*�=�F��֓6x�5�46pV�uԭvMu�����9b��R����j�Ԍ��g%H�4Wyr�ܽ%���e&�or�p��IC!S{"w��([�nԾ�A���P'1�h	��&[DEl�,�3��U�� ��l�ȝ�DX��Z�[�ɬ@�\�5{W+krƕ��� u�l�}B��4�S�i+ PW�\�eG�'��7j�̳�s5]�R�+s90�#-��.�н�����еK�֝�k��lXM;؀��K����;���3Huس����4��2 ߵg-��}��:����h�}���b���+U�sn[�K2�h�3-����h)L���J���X�0��WƳDү�s�c�\�S.J�m�d)O���M�.��ζ�Z�*U:p��Nvv�ڴ���o((������|����w9eqw�ㇾ����N�3+�R h��*t��R�*`����3h0���-���w
�֕�h/�з, �|������W˷Fz�޺���G�XyMA�$  }nݬYJ�jC��]������yA��8��kk7J|.U�x����fQ��SR�v���mv�Z�]�nh/�Rt��-��~L2���}t��ŏ��=�+;�r5�7[��=r�˾�	1�X絒^�N D2�k�nam�	�M&%r�|����Y�%����*n�K�QQ�!�/*� Kʔ"��f5��l}�F m�^���M��gKj�pV�[B(�{k��r���b�nL���WG��ܵs"oTGW>��O��Qs���t����p5J�9l8k�C�/���yX4��L���(�T���;:Drp�0�N�l��Y����AzMp����}{�PO*�0L�8�Of�ٽw���Ǉn�.��E��KX�p;�N�y��S�έ���}�E��i�2��!�c�b�9�����O(
�Fn���
�+��}�[y5��(�bH����e>tř
]fV��t����>��;�SNj���p�5����K{s��l{b��7�g��Ѡ�9�$��������<���y#����щml�[a�����<]4��wѲP2��[� ̭�{��uf�ׇ:�
-���ބ�cqoZ��Q�����[u�o�kD�䨞颠��Ԍ�h�=����!u��5��m��n��ʋ��V�mj�+n�Z�*ÏsI
7jf ܤ6���j�߯���ΖjY"�Շ��.�Ýwp��\A񨞛*M=�a޹1��z��+қ�N��;�w�.�|�t�YB�
�C�f$������"i"hiO,��*��
��F���������$	��" �"(�iZ������("
�*�ij���)�ZB����fi)J�"Zbj�!&H���(Z *���
���B��I�����i(&���)hJ��J
��(�������Z���(���)h(J�Z(JV��(Zi��J&��"%�JJZ)i2@2*��b�)JF���JX��*�����"F��(J�

R���"�����ZR�R�b�)&"�!�J*�b�?u������{�wx�*bճ�e����]�n�E�S�R5�/��|�P(�r�66��5lA�X�Kem�J�Vtݹ�%.g�ު�W��b���M�4��Q���Q���+�x�̬�<.�U��$�o�t遁�!st�e�B�"/���	G9�|����$����l
��P\�V��˴�pg^s�����Z�8�On*�;�ܾ9����9�1�N'U.P 6�,��7�h��rv���l���E�|you�p��G>s:!��v��H�SB'�x\P�a�T�eE���Wl��d�o"��,f���4T�[G!��b��Jϙ� �V�3®&7�:�S��u�=�i��UD�$��6�WҦ�P�1Q�3]�D+���)Wwy�>\��+[`%7�}R*��]{��!�G�o�K�`�k���<5pa������u��F������C��Y!��s)� h�(�q���=@���w�.s�!�Hmi�i��z�nI�88W(\jub.��Ø��e�"6>�R"���z����ݨSV�8�N
^�{������[~A���^� ;;�N��.�1]��f�옑h�5� �
��6G�n�w�I�7��\&�I�}~��z��1�����֎���ۂ�"V��tx�!y2�gY�)-�@KZ{s�Ue��ΚFB�T;a�#�e�1ӥ�K�=h3`���oS�hdcbty��L�w>���A,˷�Mu"��WB}�e��]Ga.Х������� �u��1�}�����*����i�?M��Y�T�"}%�fӪ�VͲ�0_���L��m�S�,�]~�Ј#'DuC��i[0.#ڷ ��z>z��Ɔ*v�YyՓG���C�
��^�W�r��ث������?&)�C�؉�l��tn�S��K�Eӳ`��&����Ǒ�S�s�3�)��<sE]���Ň���3�7�e�G>Zͼ�P��mMΨwyBŰӼ���Pz���|��N.�X�T Ϩe{�*,v]my����po�f��˲1�/?�r~�Χ㏤��Hxz!�R���z��H��{Y�L�aTq��U�/^V��H���Q�-��X����R0�Ҿ� GW�ݑ���FFA���n�����GA����P+�c�����u��Ν�c �z[1�<���R��Z��O���8���ͼ
�[k��+UP�baq��xk՗�'�\��I�i���+ww��Oa��,��������\*�tn#�HJ��`�6�a�������E�f���
Y6�EBenibc��{j�S����ݟ��-O��B��vv/�[�W��%Yj�u�۬����pw�՗	Ig�ɻ�+�4\1	��L�5���z��*--x3�{��sD�����wf_*�)(�M�X�M������fC���Q�jNK�����[��2v��?⪾����HvͪI����?ql�_6�p�Z�",	N���G�%�S+�@�.��oWp�x�:��Ɲ�Or_���7��&X_#42��0&9�9*���F�]Vjۻm@�Д��8����i<�*AV+fsc*o09�p�����!��+�ۯnIw� +G��w�����#���Q5���
u9�s9����r��Tt��2�lh�4����	��xmCF�����.����\%.n���Ԍ�'�R+��|�r�.!��yo���L_�o�`��0����
���t��*0�zk��Ztu�����CN-8t���5ϓ����<��]#�p��g��:#��F��V�^����OT���
��"o:��S��h܈ko�ƶ�r� ab�´�x��Es��C��ct��f��0�8��`���1q�1�]p\rLJ����Q��Kg5�V	+�X����M!��>���Fik����������3!����u��D�i�G�]r5�֍�ہ��%u�u#�B�+;N9��eEh�{�iI���n���5Nedz��Y�ܻv�a��=$���L�Pҫ���F4m�1��B��Un����J��݅ݲ�q�c���'�ֺ����}}��}�p7k��u��N�F�JH!�!�A`��U��|o�������Z�#�{q�ס�0��rC����8R��IT1E�gaA�A�c�a &�>�Ͼ��u���F�7m��Z�u��#h����=]��T��N`�P���|$R�* ���Cp�6]L����ٽ��傺:�;�8$� ���3ф�6�@sn�!� Z@�j��:j�ژ�2��tތ�2��?pvh�IL2[S��ֆ�F,	��`��u?k�Tj�62���x������\T�;F�J������H_%)�&�t6&��ɹ�Pؔ�������u1o���O����-��T{�Zp��㮛�l�u<~��V�+��V����ә�Ԟ:�ޭ���B�?��E]�A΍z>SƯ��l!N�F)i�
n>yZ��n�"�L!:�D��y�Xq�$�|2~�0¸��Ƃ-{V]�PZ6i[٦� �����e�ҧ�q����ǋ��i[���1�5�*���]�aT�y�~[\*��K�����m.��{ʺ��z�ގ�n!ϥ�*鲻qv ������X�/�<��d��;M�w˦7�]ר��6X�_T��dQ��Ʉu�F�l� J�v��
����e]��v5�)����ٮ��r<�Ib���ZI�UU_UW������~o�K���Lp �.�2UT0/��r����E��b��v�����+�\f�_40'��T;���tb��u@(������R�f�P��Zu
*�+��#�}���,gG���d����_L\R�8T�c�አWJ�F�9L�7+lnU)f�*��(�[��q�K�����+��-z.�^�R�&)\t��ݲ�$^w̝�9�Lv��p�
�F#l��<IUg@�_�u�L��n���۾oh��OSs�P}R��HKF/�Y�c��������D��Ux$7u��J�����[ڭ;I�ܲ�~b�SWj��n_N@�/�P��̹�@=T�#���q�S[�VT
�r�U�&�����t�ȇ3�8�k����SB$[��-�} ���L��VK$#��V�3 Ɔh0��h�3!���)�"��e;i�Y�붪�o(���=���,^��Z�ۡ��\��W-�\'��ȹ�0pW.S���=����[ga54��:�)�������{kZ~���kf�e��&�mn�~��#=yg�)�	ǅi�msf����հ��-=F��*�ҙ�U�Ĭ$���si;��7q+n���Rd�qCgm�+��4Q����Qz���Q�j:N~���[���}����.�m=�:�Ԫ�n����� =�~f�/�}c�{K>�1]sn�vދ�ǳy�����s�ꌯ����l���������
~��*`g<�'�\���N���|d��l~���t��T�ˮ��z�`�us��yU��Z�3V�()�lȎqs"C�$�@6�{[�j�[�ll��|oa:��7c`����� ;:��!��,V��vh���������Yh_����zAsվ�Z4alOS�ḣ̝7���on}�5ȁ�X�m:��/w��FZ�w���O�m�໶χ�:ɳs�%x��+f��!�X8�ǣꎗ\��:�:\+˸:���vulg%&&+��]�6�n��z��1֢)�(�{`d�}y���e�yo��� o�:r�Y���A��1M�gD�����>�]m�^hܮ�]Y׷ИG)�:��dn�d>e��dC���*���F�G�=F~��NE��q�3o���1Rq�PH����c�����K1���z^���"^��4ܔ;b��]���ȸ��T'��PeF�,W{���ԛ��{Q���]�9����ћҼ�"e�6�1��4s�������Nf��@�r�����.'���*q]�2*��P�$i�����b�:t^�o-SҔ�ܧC;r�v��ۣM���'^Ԡ�E���菾���3�t�������H(}!��Q�)�k*+���n�aq�� G[tEĉ6X���J��H�K6�@�"AUD�!*�Ps<"���9��;l�@9���tf�7YByʏ��u�sF�k���$�����6=�Ja���q���v�����{Њ98���E.�88Rݖrɨm��Nm�U��tx��wL��&�^JH'UT\����Q�N5;#�����^,yDE�0�1�D)�to�2K�g���]����8���6�M�]5E�c&�����+�假ӊbY�CAV�ב���2޾`�,�-/uy�v�����ǰm1J�sb�;�9� ���@���e�a읰�X�x�6���%xm��٠ϯ_�΢]`�+IÃ�Q{yoxc�8�d�9`ty�m浽���t�s�P�q��@��׆��Pu�5<~k�&8z�Ҟ�]z@X�q��M�B�}���c��V���;��pÍ7�p�0`0��!�Bl��,�$	MT�}z�
	��x'��S+�!��R��AY|[k�q�L�,X��/C�N�z�D��ΠҖ�j�#1���B��Z��qu�x�A��*���K9>�)�ot�c[��·� �#o��:�̍��>���W���^�����ݪN>�,v��GKN�(uQ��D'^lk����D�4ph�m�
��|�%{uj�Ec�ڵ�';z!<]t�ݍ� ��c Lo*���1n���k+�kn�Q�OѴ��U�BĢ�mB�b�H9?8��|#�s+fX]]P0B	�w��J�܉Y|�7.���P�W���f�5�`$㤰��u�M!����:�J3_-v��5%�� h�4jG��"+�I��	t�t8�*43�h�i�(�%$0N�?|:x�ZSS1�ڵ_J(1a��v+�Pݥ=���ή���9:U�O�9�!�i�,���� i��P��I-��Pg�������<�:g�:��#l��n��z�'O@�S�'0Y��D�H$�@d��h��=��W}z��,�U�"y�&9�-����9��~c����/�u�"�Ȑ�F����m����)����U	F���݃�٢�ZU�M����P	ݰmԅ��ΆL�U}���L��!�Y�gN|�#P����T�JS&M��g��w<:��j.��ݛ����|j�Z��������oh�	�9��h�'P |����%��ۦ$c���ё+�79?������|C�rK_P�՜��:��]�+�Gz��Ն1!#0�����ɯ��?���,\c}�Wr}�W�}U���w����7w�q����a�N�>�B��v���7Uݽ�Ȫ=�*ݛ
u�
nB��'�Fz���ۖ�݁���5|"��
��F��5uXxA�sz�Vn��n껵�8ۓA�.��N�"�L!;m�V��u�"�N�@���f[�L>;�b����y�G!ʄ�}8q�u_GA�J�9hȉ�o'����P �]��	�J�O�vF��y�i����Ɗ��=q c����*�-��{\"��p�Ǖ�cY�C� ���8ѱ�I��ܖ���LC(.u������ip�`�f�.K[3�T��}t�d�}�M�O
��×G���b��0�gB��}1(��Y��9�z�3�� ͔<��N���e4Q�;W����I�,�=Dexk�P���>m{yJ蘮�U9QA�-�9�
r��x|��3>s����삫Q��nA$�3�O��*��+�b�%����WW�q/�s����<�h5��=��r����8/�L�r�4a����صXT��)�#�����HV`��u�ﳑWvaRV�I�S�&��j���O�j�S+OK�t[�.mf�ᆯ�U_{'.�(��S��҉G��&+o;�Y8�SB|�bsl+,=|&��B�iet�F�x�Sr�0%D�������8*.��ޭ��@�U'r�i9Eww���N/z�P�8�x�3s�Ej��Vۋǧ��g�(���g�uZ�����|���ݺYW{�E"zs��d!oy��'���2P�?]5��y�١TB\��/�fV�k����V�����I�s��Ϡ�����~*�Dr�z9|���v��8��������q$9��Z	�F�s�?U�?imQ�#�J���2x�Ӯ��dfsu�9�����獵'����c�io���X�k���S�S����泫�9�N����˫{�vӄ_�)N�7;\�>����x������Ms�gm}6����~��W��D$�]��s߽�3'�?Ȉ\%���=�n[�n���Ř�1���Ť�Sכ2G_s����vI{3R#��4�R�÷eAW0*�l��=^�K�T],��=�=�B���򙿅eۧ@V#P�B�u7�Rtܦ�bI" �v��)rц=PG��K%k*0�n#�t�7�{�oO����)h�3YdY�q�ċ\k@ ԾÇ�A8�B�Vmeح֦�.�O]��+e&�:��w�M�eT�'��4��W�J��/b�6;U�E� J&�w�e(O]�|U����%��ɒ���0e���C_g#Ա��O
U��yo��O��@KW��&���iK���ȊW�v],��f������OB�I�:�O��7�a���,�]�mt芣C#ζ%�^u;ЮY����ԢR]�s�F>��]�r����R5��6�"�U܉�Գ�yݵ�r�f�L�5�q�7�A�\n�6'	�X�WqN*q{���[�AgN�8�<�o�%����w֩Q��\���T2�T0�#�WSʴf�"á��w�]j,in�*���ۭ����.�j������+�#�\�D�Lԗ��Ktҽ�z�6�Pm�E�%���*p47�z��ބ�ۤ*�f�ŀȤ�� #�B�	����� u1+������:{�^X�t�N��0�"��FJ�փ�o�w3���c��@���ޝP���m��J�Zޟ	dR�M�u��S��9n��YOb��t�HN��B:�/)"�]��L�h� �xy��8���m^�&dّu) M�]���f�����=0s��]�qo5�^���(ķ*ś۴1`��n�ؒ)h��A�ƋX�9���ric[ЌB��|KnMyC��H�t���k�k7E�B�*j=jS:�N�.:,��ݵ�w�j�W�T�`X.fܨr�}���tx@f�13�ɖ;���]F�*�%�u��6�:@�к����3((*��ۊq;�yͳq0~߸g��U��r��(0m�+y�V9�q�INj��)I��h^�QS�yS�aƆT�)����wq��4n� �w�U�J�J�뵚7`�e�)<���`�vxV(�0��Ϯ@)�O�YQM���jG�����б�9]���)s�6�a7x���4�fܭ���u��bS��u�;���Hzd��hx��F��k2�����jp��7e7 ���C����	� '&PK��{������j^9��>�h�]��N�f\5��Ig8�&��+2p��b�W�Q˦qyW:�����9R9yn޸�s�L*�����=(SJ{�+��W��(��R/����<�e(i���2��l�C�s�{Q��� ��!�{�ԸY3v
V����7�k#��a��!V��
�o(��C��Ri��ݥ��o������"u���>(��;�%=��3;C�t,G��qɋ�Du�wv��S��]�n%�)',W�#�W�Ꞿ�=j,���+�Ӛ<���{�J��W�!�(λ`���o��X�}�{�]v��Ì��rn�!���Y���x��+Y��N����N@�
���( " )j���
Ji

j�
�(()����
J����� (B���L�2R�����!h����F�!������h��J�i��JQ�J��(B�\�$(F����iF��h"h���)
*�"�2"Q�f) �Z)B����(*�V��2F��\��JZJL��))i �+,�C (
2J "%rC%2��"�J)��ɤL�����b	�)0�hj�!���J����'# 
j��׾{�����i9���zwe5�䱕j1Y�� ���Ej�+X�ē��j�|��l�y]�s�6�޵yЅ���5^�Uz��9vM֤�E���)I�:�������늱�E\W犅ɺ=WN<��]k^*��L7P�?�nr�j�s�������8.��yq%m�wѴ�.���n77\*R�ӑ���V5���������	�mZ�Gv���ݐ�f&V�J�;�9�'�I�j�Ȏ�n��kn���mӽ'hg	%��I��˅�_bg`��Dr}]r��+��ֻ)�����U�k.�ק��\��-2f���k�B3BQ07�M���]�i]t�<��˱�K��չT�^��,gj!��T�����6�X"�j"^![N��]�V��k�[i���q����Nm�%�}�.��\����H��ӝt�'�7=+nfZ����.e���ƴ*2�*ۚ��6ES�y�<i.���J������%;�W���J��s�7�����B uW[\7l�0�G@:B�;D�ʱ�q���w
>�xM�zJd���GJs�ɗѝ��<�[r��Ko��rʫ�X�g�W1��jWQ�O_����{���ڹ}�n�<]��9PZHZR�ꐍ�<�I�l��p:�ck��*_s���]��q\	��������ARd]��t��^)���-��Fio9ŉ�5�j����b�\߽Ó��WuB�hnP��BNk�5�G��8�y��p��U ��D�ܹ��7����Os��&y��C�j��_��(jFqH�;'ZX����J�$���|�~k>^�V�+K>��ʎ�C��9g7�u�8W4(wυt�p�Ų�����3��fnm�}�Nլt>�<�v�9t��q=9_K��u@�˛�v�9�Ư�5��,`���λ�;Cg�����эe�YݘY����_-��4���'i�����=V`��ѵ�]#~��w$g�%ܷY}8\��N޵����K��t	z��{����ڔ�o�X�"xZp���*۱�U.��Y'�ڵ�5��Y[�eϋ7�&��T��[ϱ�ί����:n�Ӂ�B����0�ϦH"�qw�7�X�ۗif�l��k�ͺ�]�)����r0=1Z!~t_fe��N�ɬ ��A!0��R���X,ޭ�Ni)�[u��PgEfQ�{$�e�d��L�4���)�L;��q;]Z5�F�1��؍�1G�P���益NT��Oۆv}���O�ѷۍ��x�ӪSQ�r]B����'����#�ɥ�k����b}p�f�I4��o#��6�*!͵ĞO\�:�Î���*:�_/n�S�K۸OoP�3P����
���cչF��Lk����G_e�������ڒ��DK욌Y?n���I0{FB�o��Rxz�e5�6�T��ky���_^;�Q�C9��O�x9��r�O&]Tޥ��G;�	�;P��z^Ѫ~���s����Xyy�-�h��ξki5��+_:�j����5)N�k�����k�'O2Si�IHxsm/�A<}�YJB�o�By��w���%�_���������ad�1]��uB�ثN&�*_�����󲧜\��{S~��?/��Xy���%ob(��ʈ*��_K���C�Q�1D����7_z�՝����U��g��>ڂ� e�D������κ4�Y%f� ���w�Ѭ�$�gD�z����na6��or5����N��^c�v�w[+f���<q,��qŬؓ^q!Q|�w'n�bN�%���d^�6�h���=�];[�=9.����Q�'��#�T2Z��(���/c�Ķz�*�uAW�H�]Z>����iN>d�,w��ݢ5�i'�랅]���<o�_O�8}X� ���O:KV����M��q�w���_��=��On
�V7
]wΨ:~�+�E�!VN�c<\�%N90��v�ƶ;쩨ipɨpT���vu�����uo_l8��3]IY[M�|�w\B8�S�޶�9�6%cyupy��rl�'��_ZpcOÔHS�W]L������l���r�_�&���o�Qv����N�#����a�p����5�ϻ��5���3��.�m��Hle��*�ۚ�2清�jJ�����-�0n���X�KY�u�^��7��$ø�\k�p�Lts�5_U�49��Մ7�x�u?5��q/���E?n�.JM'��k�
n�5�����ꀻU5�^^�s�`@<�P�]�y���:�P3Q�]n�nP��m��rW&�Z͠�[��x{�~yY��$�s�<�]�[H��H��_`b�\kUL"�jo1�T����ܲ�;n�wV��6	E�'�+ۮ]�4�n�R��2�]�'H�<7pŝ�Bq��T��ꪯ��2�^��1w�k*�����-9�����yJv�ڎq���`�̛W�z*�����]`s��_M���9�VV�闗��oK������[OsG����τu]�"�~�Urr,�G\_N�_��i;նx9]r�u�ⳏe��#��B�ҋ��������}�~��GJ��躄5���9q)�u[J�UҒ��->�W���}�l��V;���U|f���+�1��'�\�`���#�q=�79�4պ���W��=<i]-��P*�
	n�ׯ{�7�#���g3���oCv󖸇I��|�njxɝ22.h}�f��V���"���	�u�����C����-����b*zrKǣ�-���U��9j��y��CU��j�M)]�c[�v%��L���L����_S&M�u�}<�xRrVUZ<�\Qy���G��3��Z>每	K�K�Tn��!�����EB��?P��ތ��2^��p*Q�K����r�oh]�Ug�md-�)	��.N�x�IƐ�������=9���6��ܻ�oKu�q��YE����j	��I�
u�iܙb5�sSB�p�5&��}U�a�
�6�N��|�'������|�ҙ*���4���J׊���7$q�Q����c�`�����I�l��g�m�S�sJe�}�.��DӅ�6�t]��Y��U��6�k5Oݼ}�.f�m�p�c�n%;as0�d�Tu�(��/�p2�y%+��f�Itʵ�Mƴ2��ر7�39���]N�;��1�Zߎ>�^Ŏq_d���[q��2r)4�S���:��r�z�*J�S�ozg֗g��B�9�}YV���$dLSê�$T$��J9�=�=x�[�*�\ʈ/�f*���+F`�SǤ�.���O�7����$�+5�k��W7�,�U�|'�g��]I���f\��juq-X��\�yP�z����]�&��܌�Y�tX�]X�y��-3�{��T�+�axA�]P1�TQ���N��u۶�+�2.d���7�Fu�˼=��V���VCL\��J�j�ɪ=��/d�|�`�f����2XZK��UnV�],�����E�'�G�L��y�k�3��r���.u�Z\T�9c���Y�æ��[}����FE��G��	_)+�s]�=� ُ��Q��Qʾ[-_�\J��M��ŷ5��SnSgz:��G?�A�-5�|]����|�$�T��p�T�n�OK{��<픢xn�pX�4��n��U�Cb�p�ү��9�qy!_�v��k�ҥ���\%�v>�o�T'Mޜ�ܦ ���ǖ�W���ckÛ��D��Ü�������ې�hx�k�S_'%�/�y��8���P���.�Y�,�	�p�hI>�淐�m�l9�0�LR�Z�yپ*�Y��I����T���F���ҷ2�	�f��3ɾ�7��+�]{�y��)��Rk;�Ź]����Jf���>���~o���0�1Fn�ȶg��������������_V��x�y����K���S�z43��,R���z�2kjTm8g�7j�=N�z�O�;\�������[,9�P���$��.�H���B__�b�tec�͵,�'� ���XC�ޟc�Q��Qo��I�s�:����Qwk�T���:1���z�� v������[��p�����=��:�٧L��|�"�I}�2 ����ޛԒ�_UP5�=��Z���aQ>gJۈ�ᗒ�6��W4��o�Cۍ��-ﻈ~��Ź�V��x��}����o��\cܤ�'&�<��w��3x9;�v�.���j&�+��:�v>h�p������=.�M�L�u�c��}�������l9���G�ꔺ����N�f3z\;��9��2������*ƶz��us �!�D�]_M;�[�+�3Za�YZ���R)���}n���U�Bke�p@�{���/>�`U�u�7�γ8���@��zˇ��i�AY��nP�66�7�Ő�(���W�5��."M��-��k&����k^��8�Btދ	�3]�;L��U��*Q!�B��i�����q��q�m��6�v\�$"�Ky�K�\7%w܄f�J'���[?vn�ZI�֯ru�ڝj�ɧ/�H&عqK���Rh�+�N/�����#Z5�5u]p����#S�-�0P�J��*2N����{z�D��/&�NO^���[.�\ba���KD!�ux�&���������v��M�c��Q��y��)�G��#tJN50uh�v����NW;!��:��Q��^�'|� �^\�!��b�fj��'�¸W�7��Uq>*�_j��~������s�6$����f�B�z��F��o��I�2�]�Y�qQ<��q}_����	$���T�Ox�i�r�d�j��I�N�Mƻ����qq1��ʉ9/�T���#;ֵg�ZXb��|�b��=�~�N�yJv۝�=�챬�9s6�}�~n�>��6�jNϨ�E��ro�E��^ZN9�we,�U�j�y^I��Z���S��*9[9/ʃb6p��ܠ~�u��E�`i� ��-����wg�w���މ��.EC�{zQf*���OR��d൓�j���G�^��;϶_(��KO��W�m�cY=�V;���U�֫�F%W��p����0���c�&�)���>���Zz��њm���\VY5n*{et(܇i+m�ȡ�ɨ������o�>]��^u��2ڄZ-O�b�;`��~0���S����G���S�%��M;:��a����%�+c5�>�rub��4tPj�	ux6����RX�y�F���&��_}J�5�������T��=֔��oCwo��I�U�*z;5��,��r���Z�:`��T��K�p�L�g7p�5��=���F���N֭p�x�gq=����շyUHk�C7T��Fk�{$:����{3������Lc�J��ܦ Ɵ�Q07�M�[p6���].v3��y�)�g�LV�op8x�ӪsP�J������#��<'���-�<�k[v��VL��f��ID2�;�q����}m�|�\����Yn�����N9�D�Ը��j3���\������n5�7��/)B�&��*�٩k7��ɟUp���8{���[���&}�ޱ�&�]5�0lR�'�h��]��y�뺕7Ƿ��L�{����#Q��8b�qb��@Ɛ��{�uɮ�/�A��r����P��Ĝפk�����}v8�����j5�y�Ĵ�:a;f�K9�i��7�R�Iʘ9��z�L�=(ۃ]�x��N[|F�;�K�y�DL�o�dWV�`B�2�ٸ�J!Ke��AD�^q��k��Wz��:��,�:��#մ6ƭ���=LtA	�չ@511zsi[�̛8��"�����_e%�mf۠�������+mۇeЦ&Q�{-MR�f�����p��Zҭ��]��Wm�Dޜ��]�k[�m+u.�
;�72;x>��� )Y�we1Y-r��IB;p4D���:}�܍�^l�M�/{y�{q����EtoL$iL��e��@ܶ��[-���E:マ4�+Qnp|95@<F�߰�6�7���~̭uw�F�Q1�f�7F��5Pl*n�K��N�e���:di����>=F^뢞���{\r�Z�
,�*��f���I�����Z��d����p&�Q��w�s�f�/&� �8�V���W�N�����k��1�2	ۄ��QNJ[%��f:�Mw&)]:]�dj�[w�J�C�d+�$/���!�����ۣ8/qw�Z����E�����\ժsއ�԰�_2"Vw\��l5��6�_.8,�oBN�nՔ6:���(>;y.�7]ql�ܘW�/9�P�J.��P��2f,�-��L�$)e�ĉ��42�I�6�!d�I�E�{m]�J�mmcۮ��Y�;�֋�_���H�RR���T۩g�uu�LU�Y[S+6Nu�ٖ��}�1-K�����l�Y7�Zp�VN�q]S�r�/i+7�-
��@E�-Z��
�=4�`�\bKu]Y���.Y� ��
�\8{�Ө����(�ވ�kN��e
���#V�[�IކI�8ܵ! ������_H�X�)%s]Bu��(���G|��%���g'tav���0�.kqu�"��3J��ެ-j�b�Yr� |뮢��WY��� w�wVC+sW)��r�R�6�#��k�U2���Fi�����u��Phuƻ����U������44��l_={�ҕ����7��}*SJ9�-~	��'r&\�f������>�i�7�:a!�q�/:��8Vi���M��mh���IΓ���h�=����oL��J],�W��Q��ӫ�8�B�v�ݧ���޺ջ�ev�yv!��Ĕl���۩�N�)�YEk��Շ�o��j�Ę'5N$�� ����U;#�f�';B��������s�t*h��y($��<z�Q%�Y��!�	���Qq�W��r=�خ�ADI��{��DU�}Bn����s�sI�x[�ڳ�
{M����]˩eC���,�Y���Mn��B�����X�ɼkt��S�/�9��l���bz�[Њ�����l�-
�ֽ"N�٭���v�_��ii
��
*��(
B$"ZZB��
B�����2i��i(J��)�"�i
��
B��%)b��( ��"ZF�hhiJX��%��$hZih�����(i
�($h)F��J ���J!)D��
JiP�iR�J��i)�ij�(B�
JZ�@�)i�bR (Zi�)D�(J��.�uuwUUW~��|��	��x�3F�lJZ��Ž��J�v#w���f�qQ�r�T����[��a���;���{Sݦ��5(�U}�:���=���-����v�\�3��YW����}03D���G�k(_ո%�,Q��ȧ��j�ҴZO]����.�\څ�2��|�`hJ�b9��ꇽ�C�8��z��ˇ�8��q	�u�<�����ڴe�8,d޴D�(|��[=r
ڗ=Q��@�P1D�˛�I�u۠B�f�eV�w3�y%��@���Q��Il�iq0�$�LHC�u��R �"܂��C��D�bk&�wn���8����W*[J�m�ݺ�qU���՜5Z������m�eR�ب�`4�r&б�)��Yv��-h�f���QҞ[Z�c�Q�e'M�i��ܶ�9oz�a9y���p�%[7 U�1۽�f�R��}��7�+��|ꔦO�[QWɪ[��0��o�"�eg������Ъi\C9����
���.Gt��[�"|�ŏ,اuh�@b?W Ϝ��[G��ճ��P�F%�Yͨ�d����'����{���婨;��C���}.Yב���	���+��]8o=�َ��4䒔u��>s;S}��{�{}LiV3��]/�m753�@�؄ʊv�YyS��~��tA7��ԓ�x?}�P�1�o��V�\���
�.f�7���Ѱa���e!2�u�]ctT8��_maP��G��3=|I�̶�i�9��Qǔ���5	��p���=N����^���l����ʛ�D�
�˻�ܛk��ٹY�i4���M�y^������pծt���s�=OބSvz�����X�{&+*�����N�x��x��8_�혩{�\{��[�0�ob�M��x3ܺ�q�+E���=>:���H����&C��;&m/(a^��ZYA鸻�'�5�>����J���`�e�w[�&Ý�t�5��^N�A#=k�s_��:]^�:�	�Fw�S%ձ&��ھmJ(��8+��*y���^�f�fܗ�V���z�=m,��^��u;:й7L7��7�}p�\}_&�]��_O���%�EL�ܭ�N�g;r�YN�H��=�Ś�(|�c��W�3d������ j�X��}�4�����Tl:�*p��<Ě��Wв���֖�-U�K�V�T����c2<��{�B�q�n+m�۶����ԭ�����V��GI#��d�|�&��]+�L�;�r����ކ���{M��_.�WˀP�]q����SFi�(y�Nq��N���Jym��x�M�E�b�+����Q��[�����W>��dIY����Wr���{�8�6h�R�9�T9��5�%���������WC�l��^2�7�xݑ��E˾��V]R���	3�ꜢJΐ��F�>���/��k��Ȼx��[�m��g��>�c�ڶ_�+���N��r^N���1���<2��z�iF�Ӻ=�K��z����#�Q����,���(�o��M��)V���<fI�/|"Yr�Mb��oy*5�3Q	��p�F���s�e�Y��Y�[KAN^��R�/����t?R���,u;���Bb�zS�n�xrs3��y�m_�P������o��9�>��F��l=� n(��ێ����FVuB���AQ	��GJ��O���7��ԍYP���pp;`����-#��0.,��w:���+�mM#^N�]�j��/l�Ԏ�7�-�S4�掜m��B�-fI��!���#��Y�K��|gnZX�rk��˥O/ަmǘ�t��Us��/>�����P�^�k9W8���(������\��z��V�|;M_���:eѦ�(U1I�7;
���-KO�^�_c[=uc���t#�WT�tCr��o$��n%�������'�&�>�i�uς�ߡ����k@��e��{�¹�3����v~�DI�.9,+���7��>r�,˹�;��*ﻜ�I��Wp6(.D%�_%D�vsv�5�� J��**G����;S\}od��	K�S`�;�����Y7b\��P7�i֓Y�J�x������le:�� <.�ܤ��QCy���+�u�꼃5|q�ׂv\s{�SJٽz���xί����$r�~�7Y�ee�\m��o�=֣���ڗ����|�J���lkob��6�˛��+udeFuF��o[����|u�]�Hc���l���i�.��44��Χ��B�{Ϣ@�F�y��ׯ�F�-Vͮ��:s��}�Nui�Z�fՈ� [��ݙmS0���\�o�8�Fh�"�ܡG���m�ג�b 8�8_�Y����v����O�����x�4Wz'}�r�j|��]�7,'�/��+5L-�����+��f�.3V�P���G�_bɍ׊�IT�ZL;Eڢy\1��ZH(��X��GtdJ��K큶�e�nm^��6�)P5@ ؽ]�G��.�[ԡ�x��Cs��0ָ���1TQ�C��}�����gf��/�"bP�Pl��JlY1�L�L!��}Ƅ�mW5&_�5�I�촧����8A�{���-��I�}/{^]����fF_o���rB�W�P\��z�W��t���s>^�[;��9K����DsΖ�a�G�N�e��Z�ݔ�nW�\�:�<T=��o-j\;O�Z�2�uܵ9JqYծ����c�v�����A�5��Ԧr-�qغx�|��}n��UY1ݵ�U�������s�"��g'Wr3�-��h��A�̼v�Ò�fMc�²]ɣ��ߞٚ?7����<���8Ki�C<�1�@�u���G��}�����Ni#���c(.�*�A�~Ѕ�$ZΑ������ە�]'Ϯ�b��jo�Ҭ�D|.��Uh{�\�X*�����˚�m<\�C�M=F���T�'`��s��Dآ�F�f�eӈ�x�JS�kZ�|3���N��Ӂ�B����]�g�wzv�[]�-������{4�w\B8�[��T�:�t5���2��od�c�ﮐ�r��;�of���B�(Yb����7����	�?����E����«	�M�����iG�[}�U�ϻ��ڜsG/S��RF�U$5��:Ѹ�Nإ6��W�h-s��&�ņ �E,�y��q��c��R�`�6�]�q:��c���O���z% �o���jG�Wv�h�y�iΣV�3I�:Ѽ�\\Lk��1i�]d�q�������ox������:s��=��jR��nv��y7��h�|�e��v��w)��Z^#���.��j�<��{}u�^Z�7��U=��z�`p�J& ��:;(�Z軷t�㌌G���dc��&�s��/���5�T�-+in�� ���Q�{�������Xq8�~:6Kيu%�b<�[�BS�S��S������Q[�em���B9
�,.w	�c�(͒
,�t�V�EieP����B_c�����'\o$-]�;J��P���=^����2���{���l9�G�a��ϩuM��u���7����P7!�IE�W-�O6��Q�l���
�b!���0�� ��y�X�$�1I����{nm���s낯�!5������-evo{�^�������-;W)X��ކ��yͧ��Y���D��ʍ�;����U��5:�5���IԖ�$�;V�k�R�\4ס�6�n⎐��y��$�7"3��O���Q��vɟx�=&��z4��<��Gw�j�)'�LF���+�3��>5<�
B���W��D�'B��돁��}���O|�&������$�����F��J�q�����f>�V���i�����K������x¶n%;sJe�}�.���뫯Lp'oO��+טu��!|��U�����\��n���/�(�֥���R��2 �x��N�fҜX �R��hx�gJ����^�r���Ȇ��w�i��Xk�E��f�m��z�֥nk��Y3fp�Σ�*G��;]O���X�@���:Q�S&a�*��WB}Fy��9~u:`ϻ���\k�p�Lts�8��5��"��[�8r[̿�,�W���Tk�N��k�j�MD��P�>����7#k���j��b���H:zg�Ш�?�|��p��y;����u��m'�\���e{��~�BNt������������iTz]6�\8�n9(���ޏ{r�޶s������̞�ʹ73#v-:�ͺ䁸�X�t�8��)��6�:{xvԹf����a���:dB�p��F#.zV(�\8�p���>u{��uF5��C�z�hT�hn=
9�� 믧��zV}cLv$��O����WܔjH��\��Wo�����؞��v��lr������l��<[ƟN�3[Ypr;Z����A�]p7
��t�v|�JU%�TNvsq)�1��Ӗ��:�9XKi�}�A���o�3�#{���%q������.�U*��`���Դ�܌�fE'�A���zŌ�]� {<�^ۜ�_�9:�$�a-al|:�FZevD7R}J�F�	gg.�ـ��k2��!nԠ���v�C��S�w�(�Q��R+�i��;��+/��TB��د�p�*��ιp��(���qE�Jם<��T���x����le|꒸�_r�`%�ڨ؞ި�����t��zr��58X���L��J�nZ���*�^+�$v��E�Z�]�/��qlvdԦ��>��	&��e�w��ب�6�Ѷcw�A̞g�L�n�=K%�!�| F�RV��'1��W.f�����^�%��R�/f%;/�e�����_��}����
���S���>�$�O�:XNgZ�of��e���zћ�q�<�ʱO� m��e[�N�+�w��{�{Yu��R=Yܱ���5��5ř�p:E���b�y�k�+�kdŅb%�y-�(N7�e_^����Z{.z�̷VV�{�f3yrr{���t	��0��+sϷ�ҴZO]����kܬw���cFv��y�^������
���4�L ��e�T������X<�3]M[ojbU�d�K/��A��復�<%���Z��;:��j��}ft7"���}�WJ�:.W%�óc����c�6���F���!IYn��m?|<�_{WŘ;׹U:�Sޗ�T>�����E]�'4�ۍ3�ar�w!�S{�.��`U@;Ş*Ÿ�1D�����J%O�r��h��:��\�[Ϳ��Q�l��\LA]?@:��/��Qʖ�J����������w��#��8sw�}n�����[�*xӰ`>U'����6q[��5��p�#6���Dv���Wn?�OmM�p6ʯ� ���p��a]tě�\���
�_Im*W(�nֻ�|/a:oE�'�>����(�����!k�+>�q����it�@[��w�R��}��������%�yfq/7[��L�O8��T�X[١jM+�g5�a��
����GB��գ���j��+���L��>��C��[W�1;�a��[7�$��9�Z�܋�|�W����N�F��z��Z侹q�̗���q��, �ݳOu���	�F{��$���H����a[92�g�������2􍣕dcw{�A�A\'I��m���Q�i��v�`&�W��(�ː鈗�w.mp��W���,�kf�ͺB��0�
�ݐj�p#if9�(V�XK��/���W�*Uضp�/x�d�T@��b���٠*��{�J4+�L�t\���i5e�r]
*�������K��or�'섇nj�b��ج�����x��\5-ⳡ��U��)P��vR�r�/� *�R}jE��e�V��&����7S��Y�I��uj�GI���-���p���XXt�ŷ��4aW�u�nf](U�u-n-��<tvZplysw4�G��Ywț傟v�j��h�w����>����Q�Bmu\���h�wi�&d�����r��eԱQ��Z�,���mIS���(8GN�+�'cwp��>玣x2J�W2�}Mg��cU�%3d��qC.�e�-W"�x��,����R���h��˛E�"���M�3�kI���m"1�קEs�"	ݝ���"�V.A���d�����>�Bn�*�'M�����s2��l��F��U0w�;�=���q�v�;�^j�2Iw�r�k�9j
T�5�Hǵ|ѥԴ��]2�E�Nu�.���l1ǣ��l�[YQ^��\�.�4Kfq�
��5L��Gk%�/��#iF�^���k{�f�G�����S*D�k�s��of��ʼ",t{�����,�6ی�K��m֚��D�Ya=У��9z/�_�5
��{Df�S�@�c�<��>�u�$KT�o'2����6�i��e��k���w���Mu%Ѯ�}w.rɓ��mm[��Z�54^:�oeɰ&�ҏ
��6p�Rʏ�r�<���W����B^������|���3�T=K�+���K�w���R��n�(�8/M�k�Ql�<i�s�9ܽ�R|o�;��LR����tTX��ǧ��1tH���J�n�)!�b���t��m�6�j�-s���N��C%���E�k5�������w;g]��dW'=��̽7At��`�%̽�A[�����G����u���#	��uL��"Ŵ6��;�w�`[�c#4N�xTp=4X��Fzխwdo:�:�[����R��ͺi����v54��tD&@��N���И��hf^��oe�w��9ϒ�#�˺�s]Ax�i�:���NƆ�W�a�s~u3[�{��e4o�$�v�����{���y4];Op�:�eФ�� �Q��\S�6�B���KY�@�,_j�2�M�YB�W�/U��rf76�2�et�GɑG4��%WR <�Rnt���H�o����*�9 n�s�#���:1�&ۂ	4��V��E��^�f2��]'ͮ��iRb�U��G���@,ؖ-c��O�}����5�۽Pu�@5�RV��
�����y����3ΐ=��)�iZF��h
 ����T�ZhB���h���Z)�hB��(@��D(Z)�R���hR�j��)D�B��iJ�iB�)�(ZB�B�(A�hhPR�
d�R�K@!�H�U�UU�W�]MM��,1�����j�m���V��Ŭ�I�]�d��αNBe���w���{��V�R8��$Z/@h�K��Lڀ��W"&=�9��R}SQ	&|ۍv��Ƹ��v�_FS�w��yR���b�;�ӹ`|ϧd�m[��F�-8f�pv���qq:�uS��}��r����U�yTbXyy�>ED��i�N�xuz.9�	�ʵF2cL�eM�R{�s��VpP��BNt�����f'�u��X5'�B{�n
���/=�f�ޭg��d�L���T9קJ,ʉ�:�v>{��v-3��3�y�A}^�9�w�9U<�R������;M�0������=���c���e�J')�Q,'��\�n<�o5��V;���S���~���5�u��P�O?�a������c�����s낯�X\��g٢*�7 k���e��WW��i�����j�\5�����z�i한�Q��X쌝�/qT��x���C�RR���5J�aJym���p�v�tv?
� =�����,5)��@6A���Gn�f��$mY������2];�����q��Y�+��f�B�|[4t!f�*ok��SuY���!�qn�ǝ&؜�
*�\���%�x�Ʌ��f�;q��3�j�N3�f�C��*R�?��i�}<�1(�*�J͖�T��Jgn9=[�b�633q+�[�K���:�1��:�)��ڑ�0�����[���X�������)�Z�s�m[9�1�5�v�S�����P�L�������K��õ�k}�՗3�c���歗�öC7�������_M3S9m��@2������ܒ��F'=�Dr�4�a�2�\+�N*U��^n�dWH+�k���B��ne�)��bɎ׎㒣Qi�5	��k�2l����ou�x����hԛcUZ�UW/��G���t*'پ0 �׌�C��pɽz�ѥ�m)�Jv�9�/���m	9ҿF�	7ѥ��Ǟt#�o)���r����z�$���}��[9~`fTt��F�@\=��v;/Gt!�w�QQ\��?���o�_�3�x����<��u��K6���������b���HSn���")����8R��2�4��*e�E�2��R���ڱf��J2,���/TLkV���{*�2-Nˋc���Y@�E�B6�]���ٌ�'��Q�l[6��]Ҧ��=W�*��"�)l�S5�VT��
J���n����b	ڪz��
�|��KO�^�w��'k���"u��;'�����P�pr�-��=R�u}�}cO݉72�����s0v�Y/�mVgqR��֗u�p]`���G%�.����;#n�H�D�F��&������P�����AP����	��]�W�m@:�X�5
6�֪�=B�S��9�i�-���+~_r������n�v��a��N��Tn��q
�M)}�	k]�>�ؽ�T�;/~_r�1��-N� �#��3�%F-J�n�No��1�]�m+f��B}���9N��|�J[;.�c�JU��1~����d.߻4*��W��b�{o9*$b�4*�h�׼�f���9���P��\�JܜOb;x*�\�o�rΫz3�����[�ܽWd��ջ|8�)ZG����4p���\���th!Z�_k=3<�+p�kY�`�I���S��z�v�%�C��)Z�n�����aZ܅�Y����E�n�s�*����&�g>'��*��5&v��=[Zo_4z�K���+;\��|��l۪\wfT��f	,�'��r�4�q ��շ6byg&���P�q�/�m�_&�]�7_k��������[�g�%�yx����R�cbv��x���X��V�s���ᚈx��cz�}\
��щ�tϔp*k��hҎ��A�������ś����ީ�1����ue_��fN���yhV��Md�10��+-ͭ/�87OU����'��Kޙ�ez#k=�.Ƶ�������{�V���:(w�oT������N>}4M$M�^e+�o�3�x�O�5��1-��yU�;Ş*�q� g"ꯖ�.�j�G��g�i[x��Q�l����]�aC��}Y)����#~L�	X�M��a�����M>�t���_T-�u�t����b��,�b�j��k�L�;w.V�oC�F8{I���۱�R�휧\�5��ކ+��u{�µ��w�k]��uE���6�o;'���S^�v�^7�}�q�d�y�[�<�a�U�'�k���TD����z�ɳ+V�۷��[��Es��= �"�T4�K�E��b�:���@�������o����B/s)�Ҭ=�:�/��,��j��\�V���� �=��f*1��\֞h�os�osvU{���.uϦ��c��ҕ�p�>܆�E*%�pX��^��)�:����K���R#HJ&Ʈَ�
�I�s,�G���+T��ʚ\�;,8��E|���)�������}�r�4���DF�fr���ͅl�� �j��56i7�æB7��Jm�G�6n
�;��\��pF^M�g����f_�2~���ꚈI0jq�
�����K��ue\A'���x�r�窆�Q�B�C��|�|�}��]�P�^�3ԩ��J0\��me�{��'�W�3}/0�y��+&�F����8g<��y�P	����G�ݏ�⵹7N{�@d�}C1}�D���e֫��Z�I����~s���z��v�:����W7�.®��TM�c����!�:GS�0�S�u�I�������'6yL�p㮗%�v3G�P���	���4����LA���(%2-�eފ5)�\�#���@̫�{�տ^��ϲ
oaf�0>�Q�ʀY�5�uͲ�Q���_$�ԣ��I��������^�)�{ނf�x����]��y���q�Ϙ$�F�y��1��tc��y�gB��7����ݴ;D�_���v�t�}��eW�U���b��E���O�s�*��mig�?,ǆj�y�vLdwdD�䨥�nކ�C��������M[����W(=ؓ
����򯤤Gs�V�j����]^#]���3�Td[й����9P�7zp*��!�_�idIY_<������<��O�/`���7�'S��Z����З���O��m�8�{AZ�Y���E�{�9 ���>~���i[9�d3�)�v��9�S%Tt��WO�D�q��R=�ׇ�w�I5_��y[/��LTg�ۚ�2�'a<�B+3m�^��Ѩv�]���T�{���9��oQ˨�I�l��ad6sr����z"ق�����x�]Rf�T2ޚ��ޅT�ks��{�T���x�)�j��J$;��,$�i��P�;뫡2����.�$x�1v��*�9�5���G�Un҇�f�Cl��3��-������J��0�7J����m� ��բ8!��$U���,q��](�j4Ϋݚ�ʅ�E��oVj�a�mD�1���U���{��o;G������u�
��8�iS�,����6�Ï+��E��S��7;\�S�:E�����m�X/2PDtm,i�Z1J�α�)��8����nW�l�ǘ���L@�TgOWR���)�x���<�y�Kc+��?M����Qq=i�Ŗ��s�,���8ׇ����u���(�YEצ/A�\8�p��^���sb��] �f*�ӵ��)^n�qV7j
���Y�����(��I���.��q"b�k%�T��}��u�i�����`U_T��P�R���P^t�)Pu��C�ۥ#F�p�}p�=�*�\i����t��!�)TD��4�o �^��W��jQ�K�)���Z�<眶������N4�K5���R���u���-�B�˷&��w(���Z�c�V�ʈu��W�=������Ҋf�5�2O�� ��P����Ь�:�H�ꎠ��;G�|�O&�Q[u�9*Y�Y�m,�6������a ��E_G	£$�.�:�� ޽S���m��V;��.Wc�����:�
>�F��mto�ؘ���-�z�����
Ѷ��^�a��LE)���%m$e�|��[;��.��Щ&��/��g�#R�(��!�oT��7w{�G)�� �L��|�p�Gx�r�'O�>:�	�o+���s4��5F��q1	�
m�}�>����[�S��g!�(왗�N�n�Ҋ٬qܪm&&�]�3u�z��?v�������4���"��w���|��'��Ѧ�f��cڥޯ����^�Oՠ�~���ޔꄬOy� �,�z�|[C��S؎rp��.�Oo�\��n����M#Jуy�ON�[�}C�ե᱿�+YK�Uny�Ї��O]�����><�_D���qg;)��c�r/�����Y���UT�{oG��	[Ȝ;���x���W#�����;f�"�6�Ͱ�Q�G��>��Fe]��pN6�$��JWݔi�Ζ
n���(�r1i�h�� jj�u���+W�JR������QaU�[9:��+�/NEd��E�X��.��x�Ӏ�hM����-rttK��c��Ԃ_;�I��66�Yβ���Q�Hk�Ϋ��ӧx�w����OR�36�%�#����(�O/O�K�B��)lڻŗ��F�q����N�M>�t��WԷ�U�\L�ӕO`wr��7�!��ׯ�h��2�TT�-o.���ڄ��Sm��U���������s��U���	mg�{�µ�_)O.ֻ���6�@skX���$܎��a>����!(�Ϧ9��=Ǥ��Dfu1R��W�}��완Fn&9Iա�iޙS���K�ڀ�HXՅ�١.C��"��Ec3��֢{W4q5,l6�)͹���U�H]P#O�>����d�db�V�
�n;m�}�9/�LuB\�o�A�
���Snk��p`i��8<Ua�vq=s�/|��5�,��]3�	&Cn5�Q��.'�����&vث�U��t���e$�\�k2�,�œ�V�yѫNM�͆��$��==�وe�[f���mu�Y�{�N�O��%��Nv��R^�뾜�m��z�\h���wpͤ�xq�S�ڔW6P����7e��}Bcun�����or��Ӎi���� ֳ�P��8®��L)]��L����!|��Y���-	�$[�R��~�ت�O���Y�B�Un�c����.��gvզ��s��S��dݾ$[ꓲ�����N�ga�Ƥ��A�Mw�JV7�S}.z��T'y9v���<Us��w��8�f
�������V�N:g�YO_g����<�us��fP7�З+6��ܫZow5C�2�vTb���'y�+�ڧ�p�*z���X�&ө޽�r���r�ݩ/�C�/�b��E��m>�uϮ
�����u�ry���7ً����j�w�#�]�d�'�.�;ޫ�'�;��#�*�Ȩm�.�}�D��}�goB��H�}��Y��f�D�Fc�L*�te�u2���x��;��������_�n�W����7�q���m��߇�%�9 '5x	��@��l�Q���߲9��wG�9T=\���������9��\_���=�#}SL��?U	�pB,�:�u">��~.3��Q�c�~�c�b��M{R�ԏTw�̶���+�2�@�[qz�D6�=N��jә�A�t��ޫdy�}.��=[����t39��U��|�o8���;v2T���.��-�r�Wx.�7]�ܳ���N��{g���a�-���� i��[���G��V.�v�2��x�̠q�+�v�
�G�rЭ42���ݶ�L���WW]���s��ܓBu�w��5��Y����$.�*i*oL�u�&��݉ޛ��2n�Gs_
�x:_In:�Q��{)�Ꝥ�'WR�SGz^�ىX�&��`�7x-�!�e�1��Q]er6ҶfQYN�rD;���������Y	�/]�: �5���Q�t�����Uf�N	��*�4t�E��^m��`dZ=�����A�*��v���jm�>�Ń��YO��ʓJɳ���p�XF 4�b�m�����m�f��{��b%2h�t��-��Ņ	k��������ܩ�u�锌:�̝��3p(�֘��e�0ё^�O���;F��pg"�v�e�wA��V��$��Wk4�^ʓ\=�],'@�!G-��ld�a�$1Ιo"�V�����A�&\�E�U5�"u�2�Lr�Bƀ�� ���j���.m�M�u�"*୲����Z��^�*FԶ,7*l;a\2�6��{j��{j#P�r�#����]��S|��4�N3d4�|5^0����mJ]�U��N���sOvã,�H;$s���K%` I&����؊K��dq��!�'��4/��V�V`�(���KFaޅ�z���F27Y�M�9�Ҝ�t=���:�g �f������,niTJt!�Y,��7�xW:��;��ȅsu�Qe��R���&֙���4ӮӲp�<��d���ajP)�Zu��9��֟�$�+8��pt�!�����c�GE�Mh��rX�֍Ӭ��]5��y�g0n0����M��lL�=��F	0}+{z6m�f��ZGk�+��oBY����@CE��{���ҏ���������##�F!�k�t⺬N�W��VdG2u��޽� R#�zܙ��Z�-8#��G�S ���c
���y�� ���N�Մ��]��t9*/PVgrL��h�X�7�v�E���GXqb�CL�� w]��R�Q%�r�ɻ�U�2v�gP��؉�Q�v��(l�8䡻-��pY;�X�	�b���2�Hak�����H�O���M�Е�ܲ�J��h}$�isF� t��ճ�΅:ٸ�s�^��^�����+�KV/\F��(LSY�gƏDo ��W�l �'�mc�<�-�5���B��З!֦V�r��լ�.!9M��)4L����d3O\�ɛ�@�7������5o�vq�w�;.�eg^:\��$�e6��Zu}�K��1xőO�.�H�f����0�n�L`D�ֈ.�l=���l�}�xi
Sr���B����9�d�	J�.J��B咴�I@�9�PB� Rd!�d�J��NJRѐP�!B���dH��BR(� P�R4&Y-Pي�"(�D&H(dW�_U�_1Eژ��W;w�Ňxe_����5-w&5�J��{�#�\�9,��̝]թ�)F�̵.��]ٸ [�Z$i���ش�7�v��_�=���^��g�z��Ǧ{I�{�����YRHh{c=�M��z3����}:����V�Ж|�p,*[�C���1����N���x�d
����L(�Y�V̼�]^���v7o�{��̑�qz�TD��ѿ���W,z�\��-5w"�u�}�3�;�r`�N�9����NNNXIj����.��FCF�eA};�h����zj{o�!7W&s�ߏ�j����sI������9��躁��XfU�a�;8�w�z}�8�>�`o�6b�*���[�3&��Ui���@zM��b�=���6f�<����t>��61{��������V�<�<�4N�3�5��I��:�R�ȏuW�/߫p�߿NxΜ�ޒvv����]�q��{	UBO�5�����v��,����1��1U'�3����#7�^�ǻ2���]�ޞ0�u����9z�d�zǲ�J�B�kM�z@򸍦�H�������y��q[W��F���I���M�]��.�g>���pf�3���H����MP�X5��������V6�7���'�n;����!{+��Y{@��+�F��@1�/�������=�4�M�Ô�vt��!Ud�s@����,�㎐՘Z��S�c�x�F�ڇ&�L�^4i�
���Ӕ�[�'�Η�
�I�Vga�p.2��4�B�u��q�D��buH!ޗ���ϮBȹD�jKF�2���2�>�a�ax�f
��nH���V}�9(�w��K���엖��3��r�%W�<��rKs�[��W����|� �#���dК�V�r#�O������W������D�q	��8�c�3����=��˳�h�^��p>�o��S>nq���;�����):U����ۏ]�0�{j|t����Ū{�$�Οl07�d�u�*��5����xd���Ͻ9����K����p��w>�W�1[�Fs�S����W�SR���@�	�)�Q���>�T-�!���;c=>�O���T־9W���	�e��9@�!���W ���9��J�%�d�~���7E�ڸڇ�P�
�3���p�?�W���9>����/ z� �d3XC�_��uY꘸S'�l�ة}Z*�_���v�&Z����/�[o�*>�>���?;�7���6�������"����A��Q�ǳ�2ɃJ�j��V�÷�Ttz+xU�l�5��ˏr�V�Z��7��	�������f�x�V	�9;��$f����������n��3��2,XPg�-jX&6%�����ƴ�ø�q�y[5Tq�cA�é���Na��{�;fՀ�Ĥ0��q9y3r-�QsfL�����W);W`i9V��^�U��V��KF�XQ1�t�O��d��{Ezt���P��U�9O���s�G�kƖF��U\y���T��ۉIGۥ~::/��vYlW�?��T�A��`	��[����{�%l_���S�65�����3���\kͺ�����yL=�ʭ7E��q����"�t��w���Vy��G}���C_O���Y������QYs���2���>�Gb���J�^6fhQ��{�䤎�/�ޠ9zW���P��W���y�1q�u�Pȵ$�Q2¯����uI�/�x;���)�El���G�k���@��Y~/���[��6���i�jH)
#�Mz��۹��}�  V$��芩KӐ�h:�}��ё�=LnG���\C��7�aoW{����S��e,s��x�'�x	�|��rٸ����x�E/Ճ�ϫ̭�g�	���ב�V�>��P���:}��,�|n�3`�@TA�^*��0���u�\:k���z��k��f�{9nM/&s�	�M���#�=wlU�UO�� y�A#�n`@z|�	����H�r[���r���Ʒs����u�]�MDMֺ�����ȅ�-Ȼw��pE�Ei+]����J��$�ܝ�4f��E���w�ά;�H��i���s,_E�$H���A테f�p�]�s�Q���������,mJ΁@V��0q,�e����
0wm�R�8�}���������������@��Vxә�,lB�-M�H҅:R"Z�T����*;�3r�v��=�Q�� �D-�Q�m_�����O�|}9�}��O՞$\:��S$5
/Ңl��w��O�>��D��4."��M\l�=ޒ}UF^�'���y����P� �k�i誕����:o��ƒ��.cz��b�-���j�e�]Ua����C�/��N��_{���)iQ{f�9n;�Qs��UD�}p'tú�n�����X��{yld%U�%�(c���$�Y�[�e���סuXuӉ����ܡ�TI���;�r|�QzN��/�̝�������(Ux����u�sʫ}���o�[Gr�:v�&^���I�>�,� j�7�K}.
^�%|Ϡ-��C���K�w��~ێY
��}�}�<1�;q2�:^�w�Q���ϳ[X=���#=�J���#�o�>W�]��^��%�g���{#޽f.>�>�Gz��*ڪ�7N<�zɺ�� ���H�9�4<���*���z�����^xwՖ�<m�Z����0�x��tY��{������U�sЈ���w��7�������{�M�p�Y!F��׳�馳��D�;Dd�ki�pnU�)%���Ħ��z�#3��m�d}y҅ͽ�	�z��vmX__�h�5v�K����S�vQ2��]'��xW�g}eU|f5U1u2��>	�<�<�����p�x���F�x�㵛F�������k�qȗ��χmK7�K: �}F[7S(/x��#=~��9�b���"��ϡ9+����}�dg|�w�����-�s�x	��l�7p\w�ʪu�u�mĭ�%a��m�9�$W�g|W��F������i�U	����@�o������RiY��{7��N|+|j�p�:��c=;��v=3�M��z�z��w�B��T��xb�8���ލ�++��J����q^���	f�.�}E�N���5 �簽�������W��Mm��#�Q��_W��Qkf��=K��Ŧ��[n�O��A��}{~��G<�����E��q�%P1<�Q�d�":�2_V�Ϩ��ڇ�w��f?t����-��I#��>�:��^O�����F\
���2�����};�C��.��Ǭd�θ�u�6��nI���������9��P��b�����6f�ʈ(�|r|����q2�H�t'Ѯ��<�S��a�KS�ѵ�-Z���z��[4�M��AN�03E�M�z�w��Æ@�A �;���v���Q;�+�C�a�Y��Rf�էx<_6뙻p&䔺���s���g')��j��fk�Zv�]�6�����Ծ7"onND`ze���Z��X�}S�N�����T5&}�~�^>�
�������~��?�I����W_����ӣ:N�����E�����&eb���2Ry �V���[�}���ۗ��˕wiE���,�<t����,���3�Yܶ�] F���@�u^~�����p���Ӈ
���k%k}t�}p����Fz�ϦQا 5q��x,����~3��[�4���E�]5�tǖG���Y�пy��Y(��Ih����z����
��J���ګ�q������a|O���=�9��ׇdK�A�8K�(UD�Sӽ�zcoݷ&wG?�yG�_�d��r��vgƹ��|��z}�������վ>�:%�p@NR�pU�F�s;�'�c9c@xl�k�{�1u2���x�E9t�o�m�^{�o�v�9��
�3���ʽ�}4}������� \��5��Է���'�v�G�:�;a���#�-�)����H
U�}����f�<����+��d>>΁0�D-�!��o��?}��Ԩ����{(U�E���� ��{�c�������s�ێ�vǇ2��n٬}okn��X]
c�.�
ȵ�p�{;7n�Y�q�2�|j�9��C��[)�L.`C��:�������=��,\��M�m�������V�'V������r����>$��G9d�y�Ώp߫���g�*��W�m%�pH�O��Q|v�j����'u�5/K������'���|�� ;��`�~��g�b����`����7�lyT�v�ls�T�yѪ,fjʏ$���b��d�?z��dC5C/�CH������B���~�A܁���+���ﾩ�:.+�^��ߗ^\<�9z�f�EzM�g�z�롽�f�9ki�`�Y�Q5w�¹��%�1}�Z�O��s������j�1�ʽ����#�5�J\;=�3��ΗW�˛�Gq�y�Xr�N홏*�N�9>��S�vXc/�ld�w����W���D��עiN^^w!����(vj��	�m�� 5�g�}��Ui���a@L�PO�_��앛k�i���Ӧ��u^��?m ��п�κ��d��/A��W^�G����z����w���Td2�{ᾠ*9z���b�p�VEy\ody�1~s������&XL5��F+���3�ezGI;����}5��w�=�Ϗ��?K�Y���{��8{G`^W�i\�/�`������K`w��$��By�.��S�1�Raq��H�lh�n�&C͖b���7N��r��Y��i��Լ���d�R�-=:�=��[������u��
bn�����E#=���5uj�[օ������N��Q-2ه~ ό�>\��U>NrMW��g�����7=�|z�~w�W��3�#bcf�]t
�����f��(�"�.��
D��>���������F}���V��{M{�b`����'�x�}������;G���D���p[�*J�U�a��)w�{#<�ދ���^-n��/!�;OǶ=�C�����u��ث~��M� �-�
�������#���k�W=��=��Tu�1�o��Ͻ3�}�}ՠ�ެ�=U�5q���p�KSpH����%�����΅z�|tnȭ�1�m_��"|Y���`k�g��Q��9�6�M���������%z mX�r�h\E9Zj�^��;�D;�����~�&����|�FA�D�����U�T�� y����\�W��-m�ȧ>�W,mB�r�T���=3�{����
5��D��T]	��p����%�Zo�js�2U��}bwL;��[��>쎦4U��Y�z�1����]����\<�]�ͺ5qڱ����ֽ��3<��� ��7wj�W����'OUC�c����ؔ���u�y������^�6:�]]\������u�b�e��w�բ\�Z�FR
R{+��s9D>67gd�����!uƙz��[��cuB���F�2"�wQw���\���P׋x,���<B�[��!Pb�鴣������2!�W��n���υr��f�뜣��Aӷ/A��{��^1S�G���ެ���}��5zQ�x�t(Z��C���K�w���劳�c�mO{'N�_Yۙ�.��e��xz�xL��Ԫ:'��>P�p+��x�ȗ�~+}yq����1��1K�x3�IF$+ۛ��hY;��~x�$��rQ�G�w W�Y��W�/Ǡ��Tg���T��^�C���^�.��-��^9�YD�Pf<�|eS2����O]|;޼�P�z(�G�x�"4{��RC�{�Ǹ�K�A�d�<�$�3b�C�2ْP^!ç8�L��n��ܔS���ެ�3�����q��=��ڪF�?]�{>�:K������Hn�E+΋��^���]�e��]Y���^8��qW��s�3�+��HҮ3޲6��V�[�P�pB.(Y1WY"��_���;�m�����P8�,V|��-���z�1��޿3�zg���{����`-���ET���+\��>�RG�ā� ����9���R޲�j��O��>��.'x�S�L����|i�՝�@�� Lru��";Q�Ov���e�Ns6����������}G�)5����;�Uy�3�]���L�9�O���S�[���$v���6�:{j��V�e5����	M�e����	*�����B����
aNL���ʿߺc���S�)�<��=f*_W��Qkf�e�.TC���$D���u/�2+mo�U�w[���O{����q�W��w�^��	>G�]A};�C��ɇ�r�3�J�g��j+&��yMI���@zo���}Ƚ�F\
^P�ÿhc�5�f����?~aL	u:|�|�m/<5g̭7�uy;�:� zK��t�vG�t:�^��7q�DF5�+U�9}������|}��+���T�'Mƕ�W��M{LdC~�^9�
Y���7�~�9�:M�����B��y���I���S��~�,mFp]>_�ˬ^��u�ʩ<��K���C�׏.6,N�����O��<����ُ��nY�gIݸ3��X��&����-���h*��@�N��!�u���Ҁ�ݕ�쾾��]`�9�{H\o�]#�g	J���_�q^�FY��MP�^�>������V���w���'魋�1垻C�t�{ϮBȹD�j$�AS"��O.�L��L�,���F�`M�D/Ux,�>�a����T7�����엖�ϸΒ��IU����������ZZ��\=�yu��@E[;�PF���>���-m8�e�ۂDU�%����̦�Xxk���'����X���8�b�����
��o�Q��fv���]v>Y1��[�,֩M��w�����"#o��{���VI��W]�I6F{�SV���7��@�qi��*ٕņ��yP�ٻg�aV�ir\�f�n4����G�
+��ʂ�U%��M=���׹}N�;=�p]�Q�IՓ'B٧�equ=�c�RR����l��(V��뻳ҍ�A DE�r�	�oiUś�V-:ਫ਼=vt�i�>$ʸf� ��Pj�T��uM��v���6�f��B&��U垊�
��iYt���2��Зm[q��Gp��p%�cj�s�LΘ�[��rB����Ƃ(�kJ�e(h�T.�uI�=���|@����M����U��ae���mԨ����B��D���n�.��9�U#�i�b����Ĭ�6�������F�jt1c3vJ|B��
�;G=�1��kq��`��-|�����\��Kw��(��0)�ܙm�$�yg����QӸ�U�Q�V8ǻ&��t�u\v�n����J���c��tS.Ʋ�\��i�Mi.�)��مKǍO���O�י�j�ｩOSˊ�C�n�N�w��*ݜk����:Wv;1��̭�mc7\����.���Gu����Hօ]�ZU��v#\��lkR�M�tk���3�l��"3:2f!�G�a����U�,�yo��qNq��)��Rϐڇ;r���1�ȣ
��ʷ'�$P2CC�Q9��X��j6��c��{b6J����N�ܙv
�H27�'�X��7�X]�5�rP����|m�v�٭[���:)eI��ʉ��-�Z���8�A/����*U�G[�n=�W �G�T��WWVox,fhP����}�Z��ˌe[qo]E�6X���9c�ۧ	]Yu͎ 5���Y�t�õ�L�������T�r�+Ѩ�0P�-��� ��L�k��f�6�s����E�o�f ��m��|��MVX����H:����)d�Qo��Vju�J��m�%��`5*��s��|�}��F����C���ݨj��o,��:a�t��1��,���;�`�� |�z��feay��o }ƕ��6����Zp�MT�t8q�;v���V��9;#�&GM#�5f�X��J�6v�۱A�A�%N��"��-��N��E�����}+�e�O7��E&��a�8�HZ�\+U�c�z'aף�S�q�|���	R��#W�9��$�!�Nl̘:�7�uҨ�pYg�R�c�-�jn4\YϦƊ�"�@r�B	�,\��)�f�#�C�Kj<�a�s�]�o&��b�|5�&��M���.]�)TDқ�%cn����[sApi:2;�j����<��n�y�%PW�JR	�咆@�%#AJ+��ERJ��4�&T�1&@R��DIHҔ�(P��R	�
Xb�d�@�R�Jd��`�Ӓ�@�@�b��P- !4�IH�9	@�QFY
Y�d��EH	�dICI��!�ׇ�~]��q��+GV=w��=(S�a�Ev|g5��7M�t�,���<}�F*�2���o�~\���[�ÍL!(S���c&ëWv���3�1qS�~9�i�|��}���/Ig}�p�zs���ӢY�S��i���ST��.U�A�`�>nb�S���h�.�������Rt��z����S(Mz�Ɖ�]���/m^gh���	���zW��|K}|<2'�v�zs�Ï>�:,]�
�#7��zv[�}����7
��:��n!�	+��d>>�0�|���7٬���uھ��J��=آ�/ ��J����7�z��g�*��W�m%�pH�%�z��|v������}�h��F�����W�7���� ;��`���o�U���S'�Gr�T���9M�~��6��x��+�T�ѽ/MGrۏg�ۻ�q�_����|�����B���)b�<g��H�XdZ�C��0��DT�:.�ׅ\F��_B�ˇ��w�3_��&�����]q��V2�bj����li�>JA*�1����}�E�S�'o��C��x�U���~��"x��8�����ewD�{98^xiy���m��a��wnǕD	�0�'�z��;����4���}~��YB=��7`���x3�������+���;���	F�CJf��f�tT�;`��;�[}\���]ǂ\}C�T����lY����E.�]H;�^�,��\٫�(�6Vփ}�}��7�+��9�5�+a�Q�9=�n�1)�Ղ�,仯�<�S]��<����Z���J^�}�tק<���N���^�6�k8Nf��xk��P�+*��Q~%*�
�q��{��	�ܠ�����"��K�d:�ju�i�����~��:|���:��~�t�x�9���N��QP=�pv}\�����;���Y^W�}�_��IC-I%/l�V�e^��76=j�@�=#�&xu�ϔ��)�o��^�@{�QP�/�z�G�Au���M/D����{P��
�{��5����<��b��T��O����A�����#�z��t��^qn�����Vwr��ޅ�ƿA��adq�,�̢K�3�L|
D�>���S(/;w��:~�z����m�>��:���|�GJ�t��q��dq�>6Ȁ�|f:��
=+�V	���>g��o�B�����O8Ξ�W�����ב�~�8����m��ث���}6��@Cs������=ՙۻ�յ�j���ׄ��*=7�l�w��t��A���z��<j��T�-T������yYo�u_�]x�@ݭqR�tn�j�w�6��m�|������f�
�~��#�����o�+7}��(hB���x�%���/�_��qM�"�\=�R{�K����c���EǕ��a�&�J�{��&_;���6OX��=�X��rF;����9��԰sh�1�α��s\��t�ts�ro�诵Ҙ-5���$o�I��������2G����f��zV���^����CmUQ�ר���>�޻��������c9n���@��^���5��D���>�>�ZX����Z��~�76�<a׼��B��)��xtϗKzἊ�qލ��%\�}bwL9���/O�:���o>k}[cTNU�o/o(̚�N���ޡ�W���z�q�hu�n��*$�@8<��ڇ9>G����2��G�����G�����/��3/I�N��}U^������ul���X���ۙ�C�kz}b��mW��J7}V�\{$�x�q)׼V���r���w��E�9RwEA�~�&wGr���e�X��^��7�����Wܽk�D�[�^���F3Dצ9蚎5q����1����ƅ��c(���S>F✆U�١�5�P��_�7i�C��<�:����D/V���6�w�Ϯ�s�(���y�*���e#qU>	�ˠ�U��zG�o�:�6�@Yޱ�bW��{��u��Ǹ���P;jYa_|f:�*�Q��r�ԽW�x��K�thJ�9�<�|���4�WJ�9�E��w�!+�`��ʛ]+��w۔G�9��Tjݛ��Q%��#M�m��x��	}����1D�,0*�Ws+(n�����g3��LT�ur�'������gd����HZ�P�.��Щߴ真9���*#ڪF��߇���.��9�<�����q�ڣq*;|�lہ�s��>+��eE)U�\9��\w�~��^{�F�z�٫��>6��z�>�����^�R�<4� _�k���
���-���׭����;��n=�\OO�E�����1��xN��n37ˍz����<�H542"�����K6�o�m_��+><��������em���ˉ�D#Q��Q[��F�L�������F�(��W,z�+!��e�^��>��q��u�q=��=�W�y��;�TXї�^���FI�5�Gڳ���ኝK'e��o��G>�g)����;�)��ԟc��~�����\w�.}Նe_��|l��}���U�Z�t*pnҟPKy�Eg�x<={yq�^�������LWg�t9zFL��Q���]x8����=���e��cn��N�Ҽj���⩯i���E/�UxR����GG���U]]ߦ���%U��՟w���%p97'E)�;���Y��c%Ry �Vx����Uu���' 則{�F`�V��o����BU�Z �%mķT1����u+�ZEc��֩�n�� ݚ/:Ia��z[;�$vi�S+K�5��2�n%���T�kt!緪=#iD�Y��J��	�v���9�"3E����R`�k?{��a�eO�t�ۈ3(O�bpΝ�r�������#��ԍ$.J&�۾	v��:e'=��������H�% a��=P�+�H� 5��rvxf{}�ީ�|�Ϥ`�n@�s��z�Lyg��<K�A��PTx��}%�FUC��Q�nϤ�n=;ۮ�R>��7��3��z}g�{���w��K���엖��3�����{�]ӎ���;���i�[�>@z�C��^���x�2�-U�>�������gT-�e�o�+`N��n��18m�5���~@����J��Ē���:�V��1���v<��[˶|�4G�Z5��F��T8�Aު�c����� t�-�(��)�w-���ȟy���\��D����v�ʥ�c=�.%�'��Q-�Գh�A����7E����i��w��2t)�Q��\�hb�����������>���o��Wq�dUê�T�#$�l��~���G#=P^x�#��^x�R�e�C��\�G�5~�~����z� �dC5�?]xuY꘿���]��!)1��?Q�Q��^*1�@�)s܎�x�;����������l]�l�����s�{�r�ܸ3yM޵H?*J�����f2��3e�����y4�a���X�R�,r��C+x��om�:V�x%M�z�K�k��\�ug|E��7��畽��A���x���h��^����p�uTTc��d�?z��g���H�=8<�o��c�NF�,k^AS�|ntu����Zt\W��+Kë�.r�����I��@����\�e�
�TU3w����p�}	��6o��L5:DT�N��s�������ʽ���/L ��6*�7����Wxb�|��4��w��~ͺ�� ��3UwL;��i^8�~ {��S6�2�9��o���8Uy��T����ӞSCܧ���o���8c�k�/��U��`)u?�F��ˤ����T,ud�,�^VE��/�:�ju�i�/m�{�]Ed\�(m��Õ�}��9�����g��UZdz��;>��\��rt�}[~�~++��{<���s���_����p���5��L�"g�T	��R��Br�Mx����>>���~+��=۞����[9lD����i��g�{Ҹ�9������T�Bd�9�Aվ�xhȏ!�c_�o]��=ワ���8��/�������q�,�2�,�����n*e쇏4P��X�+�ѐ����y�čT*u��S.��M�Yn���K�y�S(��5�j�X�|֭�lKY"%�{���}ic\�[�xX%��낚�"�7��S-czVN{ݺ8q�ѕ0��B�Ͳ3�[��Z# \�7�0S�Y�K�e^1������o�N��Z����'ԼW��<��� t������h��2 'Fc�In���J�U�6+�Nh\n��;��OEz:ϗ��n���;^G��&���z�ا��� 4�$i�Yx+�/����س�?U��Ղa�*=m��9��>�؃���^�~���uU%��kMy�F�U���ev�*}H#UxT�q���[�a�j�&ߧȟ�~'�M����6��|����!��Q�L��c��DK��u�ZkKÿwz�w��1q�Y��f�tM���;B��5[�E�o��Ȥ�a�����<����koFS�i�,f��_dT/?9wv�G�^J�]���;��{�����'y{"���&�w�̕b�\	�0�[��>�����.�]��.���ή��U^��C�o�V=]/�F���P̏*$�D���Aݨn�~�t�����v����N��<�}�}l)�zOBu�r<��+�7ݚ�r�l)�t�v��"��Mi��G�������ӱ|�F���|�=�g�@�N����B��5%�;g��g����b��]v�.�w"��T`Oo��h2��`e�l�Bv��3�/�wu��*b��ܞ�F����~g��nmU�S!Ů艧�J;"�@��m�TN]\�Jv��ǥj@\�n˒����ܧ��>�@�ͽ�\a�m���\ǃ:�ݧ�~X���~�0c�}r�����YdyODi`*���Wܽk�DK��׎�T��3�o/=CfqFoC�}����|�����c* ���S>F�)�eF�]]�]������FO�'wV��{�+���Y����m�~}u�A �Ǒ�2������T�'��U=v=�l�_nʛ:�]��������|'�;�=�=�c�s�{H<��R��2�.��@�>U^dy�;;�j��H��k�>����9=�n��NG��9��P�~�R6���=�gIv� ��qX�{`W����Z��<;�D��(�9�v��E��+K�{��Y~��kV���VC�O�ۖv��r�E�_�@�	�
��
�_��\:��c=;��w�<�޸��m�����l��}r�D���ޚUR*:d�u�dfAGY�t�f�
�V��-j�ީ5.�|�/{Wu��K���+��������ר��d��OY��}Gh��W,y���X��%��>#F��m׉�@���C7�]@��Q�FI�7�먨�պv}�)�z|��{�z���N���q�W�ƐWuv�3�l��m6"�u�'k@��ݶ����|	���q!`�rխ�Y��>��-�Jv0�@��]C��ef�"QOL}�.��~��� N�nB��iX�'Q@��%kmޤ�<:�N�S;�tj�ꅦ������q������C2-��.B�a�V��K	n�g�D���݁Y��[OC����n(�O��xz�����V��@zM�n���z�u����n2T:u�=cs/'��d}σ��l��䡒^����/o��>��)x�{��)Gw�_�ѕ޺��ʼH�w��<��8����?���·qS�t\E)�N�`lV{�ȕI�<�-�z]�vz��Gr'9�G��<�毴ǶDtmx`��Vp��
�ꗍ��x��JU�9F_�4]�g_r����M�����+�67OG�������9��% a��=P�+�H˳���;«۝��")T�p�B���z��5�~�<�T��/��?>�.Q%�-C�z�q���m������eq�>��m�S8���#�'�۟o�=�9�^���ygIv1kQ�y7/}[)W�g�3�O���]L�1u>��Cɦj��i�)>/�G�O�\{U��ףM���?TU�";��W�ftmA:3�B(�71$���x�E\:v�������Py^ZߞЛ��7�dN��u��^Y]��#�G��3ջ���g��K����恤�i��}l1}XK����-vAe��H�	իQ��3��Ye>}�)+EA�VF���i�H�rƵ�r��n`�Ս��Q�S�6ip�I���Y�-��
��/���ڻ�a������[ Q�^SYP�����g8^;�lOWh�򱕋�y�;��z{I^�\O��߮*�u5,�ȈT	�^���Q|}��]#,��5w�o��(��t�vG��sĿxΏoޮ��~ȫuU�FIh�#�ͥ����������ު>���;WQ���*�j�&���Hg�=^ w��_����T����Dw@��F�}�����A�S�V����Ѹ���w���Cn���_��?z��d3T2�c��O}3���L�x"=��9�@���Zt]=�
���.��y�/]�~����d[�ğ���uo�(����䮆�*:f����� d�Q���T�N��s��������
�rG�*���]���~�Bn���{��ido�+���=�T�l����A�^x���g�����xLΣ��U%C���=��m�gʫ���>�O��{���Z7וC7�:N���xG�à�s������Y�+v�wZ������K�� �MY�ԼF|�9�~���{m�:�+.p�6��ڒ��x�lṽwt��Cq������j1���X��r�`��M��Ϯ��n��(5���M�FE���C��crK���qm�E�����:X[ί�LO��'�j��f賯��Yg���5|E�E8��!,���]Y\ꃾr�⇌R�����{b`P�\��[cX02;�C{���wJEn��#I��8��:�]�ac4{�-��6oo�)���ލS6u�Ĵ!�=�78#���sB͇�6��E�I$�y�j���{{&��Y<�I��n^4��Ŋj�Z��Q�$��Yw�S͢iz��ZXn�^�ks�R�v�G;�d5;���9���6��tP����YZV���8��Q:ժcF���&>��C���5�����n
��rk�=�a���y�t�%��ظ�H��%�)�ґ�<�_Y٤GSY�Jn�d9P�l�]��2���k|)�%�D����V
F��Yi�+��Rޟp�an8,a+��>)�p����R}��rx���g��&1Y�4R�z$��JX��5�m�5$�&pd L%���07�7�TI�n�q|ۺu��S�1�w2���Bz���[&�+2����ƿ�śC��E�H�ׇ�yϩ�q�EHJWԥ#j�rv�7|�=�q�Z�d�@8�� r7nr�v�M��]/R�**k��i=��¯^à�B)X�,�L��s�]�J�d�
/��0�kkt+H�*R�6u����S��H��nYlhX����
k��H����۝+�N6�_JBb�b"���'�[[L
ABl�c�Z�x�>��ޢn3���,|����YgMZ�B�cVnZL���g��-da��Ż�,�Hs��R�q9ʙJ��!U������e�)���Y�b��0�:S��.��M����(�,�l�9��S�T��#3+���P��nݰ�3���oU̸/`2刚B�w�x#�"Í�9a��d�k��W��&>��pWYN��i�ٌJ-V���9J��1\2~���0�%V�3E��%r�1�Rͽ��kn`嚖�d��ۗ�*[��^��[���K �~�z*q�yn�r�th6\����Yahz��A�e#���|_af��J�ܩ��`J��W#;��'�nmE�i5��+'F�j��Zc\s��i.ҹ{Y��W* �F�L˾z?b����#�w!!�5�l�k�A������+����G��҉�Ey'�z�� �aU5���q��֓n�N�܊��ή6�݁l��Q�+[OO�[}��,n�4��6|Ժ�Е�������˶<�
搲�5h-�Ԡ� ň��Z�_	3\�p[��r��O�Lv�������S��+�s��Z��}qM����|y4�
����4���t�����7�ʚ��m�
ηQø/�hP �HYߦ�~���֥D� �9�����"���f�fY%&I�b-4�!�䴅SE!@d�@VJa$�AK�8Q
RU@�d!��PP�EQ#BSHPSK��&BeY��Pd999$DLKMITSTP9a5@fbE54PAE%�feMUT5fd�BQM!1EIM994�BTLAAQVf14QM��EUSS��E$FFEe�41AIQ��%-35IQ�ADFF6a�T��LE���Q)E�U  �I�>
�Kw�d��%��&��p#v�^�:��1�ٵ�\z�����8������彽vAC�!���]A;VEab���C�i&�UH��T#pv}X�@rr�}N/��dW���y�1����P6��9��ڏ׈���9�KG����1,���׋�ި��>>���K�X��N�®&f'�Tv���]�F�A��W��QjH*���b���H\UO��fC����	S��G���-��LN����t|y��{TY�Ȏ;E�e]A�D�>���L��Hvz�Er(�ms�Q�>b����F|�W�[�GJ�J?_�=�$��C"tf:��+����#>��4�{�exug��ׄ�񨇾늷Mb��~�O��ꑷ�b����q� 9��OA�Fh�&�ѓ�_O{<4���e��τǸ�����r=3�}�=������.=U�5�(���Sa�9��OW��U'�7� t���
���̀_�-�P�W�7��O�|}9�}�uoOʵ��D�I�ͯſ�w�.��^�)�<�U��xП��l�5��!�Cj�ue]a1��\Զ����gx��B�p9c5�@��QY�<��=�+�koFE9����c\��˯]�NF�)h ��a�a�7_��k����u�rz'�ڰ�;� N��܋�O��f�6���犛ݷI�W)��.V9ً�t��'�N�z{N�T�7��D�bk����IZ�)P`�:OK�4���³8����%�:���d���	;�+ �ǒo'���Əswr1�G�S��	�^ȭ7ލ��{,�ٯk���
��fR�~#٫����d���޿GR�Y��!��/-��_�CƮ=�c�ӏ�C��.��I'8<��m���{L�aEw�o���ur7^�������aL��S�g�U^پ��p���u���xw��V���&sa�_�9�������eV�	��}�����wrex�_�Y�C��r�=�+�'&fR���r{g�NmK	Û2�A<�I��S��7���]@���^06�Ӿd޼�~���ήgg}|S������1q�}r�Y�R�,dŌ���#q�2� l��.b�L�e�T��ZU��@�l��z��Ͻt��|]b0����E�ITf<�T��L�j���K�>��ڹ�u��g_����C�q��VG�O�w=�G���c�r^�;&Yc�,�0f��;��cWE^�N����G�S>��x��;�����=���=��=��m�]�{8Β���5��e�@�i�[=�U0��$��`\Kf⌢���=�p��E��+J�~��g�De<+����M�.Z��۰q>k���}���m>��LV|AN�I��f9�c���cw���I'�#=���R����[6a�~{��}�Г�Z��sK��s�Yh ���d�2L.�_Q�YC�U�eh0U�7#��9M��d��]s+��
�dQӛ��B^Ti��,����:~�
���
��\:��c�:�ϼ"�3����B{����>�W\OZ��h\C��f�T��; �4%���?�>Ͳ=�gS�~��:�F��yS$޷��ǡO�e�������Q�*��n��F��\	�0_O���i깟Wx��� nz���r����*���>χ��w��n0
��ˁK�~�p���l��W�åB��N病����Ľz}G|v�j���o�!7W&�����?_�����}�ˁKՆev��V�����@�Y�=A3�ʶah:��~�A�3�z���w�����=�LWg�t;mnmrߪ��]ң����Pw~3^��QP[����'�6*^���Ҽj���⩯i���E/Ov5(Y�t�nzP������
^���?)��2��"qa?ðb��j3����'/b�ݐǪc��t��>��(HV�Kw�9��׏-�+�1q�ݹ�Γ�pfA�,lVMi���S{.�D��}�9���F?_.:��@�U��[��>������r,�)Y�xj�C�e ���'lB����잘�do\�ޣ���,ԛ��(r��o���O71�2���_.kobӃ�2�7�,�x�T���Ḍ|k))�[O%�T�ܦ �n'���F��,�s��=��YNNسn�Ι�Ү�5�����2��Mn��"I���76�w���O��]l~>����{�^�c��iW\[T;�r�(���������������Lo�ϑ���/}T�������O��>�\{�s�[�ȉyh;{$�ĵ�t��b����JG'�3�L���s�O�3��i���;����O���'�`���.
����8Q�\k���VG�Y�p@L�)@�>nb�e?N<u���C��LV�7~�<�']w-�����N�c���US0��h���	�\|d
�Ҽ��1ҡ�3�nvߧ�gO�Cҽ�c=9����R�o����TVé�f�����~+��v�2 �K�7/�?Z��^�4�&��aߝ��G�ԉ�G���7ޮ�u�?ғ�K�/�p}����\�|vǵW��9G�E��l����T;�5~�~���� ;��`�~�d�ƹW���Zl<�o0���!ô!�ʣҴU�R�v�Ɨ�����<�m���_����s�}ْ���/d�۳��'/�9)G�J�z���V:pz�i�t��*�^��ח���Ǻs&}�[�'*�gr&ͨ;��*�y�"B�/k���֛�^QZyr�{�����1x"	��4{�5>�J����R�[PX�_i��|L��ߋ��l���Suݥ�Q��gC'6�����-��A݆Qkwfl����Bn�n��7�gt�����������l��%pɆ�ևu>Ӣ��:N���G�����G��Yܮ�j�q�^�Ǜ���#�.=�^4�}q\w�~OqS��k�PlW�,� ��V~*|�9�޾�AJ9[�sʼ ��]ld*�|7^^���=�}�t7�;�fo@�U�LLU����~5���EmW�+�k�	�VE�J�/���Z����п�|먪�0��ꓺ�9�!�A�V�O�s���*����H~��6v}X�@Trt�}[�Ⲽ�7�1?Vp���p�F�\n�<�����c�jI*�e�_	��g�bY	�>��x;������{ѵހ��N�ٿz�D/V����.����4�}jH*�3�H>E��T���s�<����]����9�ܠvy�xo�O���q���<c�������<�� x�q�%�)����W���Z1zEg�y��B�S������+b<��W�'M�_�=�q�>7�	�����"���s9P�J�o�{�s���L.5}��A|�k����!��}23�T�?�������DU��W�T��jQ-Vi�K�ʣCN�O�f��rs��<��=�l6\Y�OJ�����Xb���mm��(��}Od9S���M隰��ɓ}6��nXu۵�8��m�qh���.(B�7M�c,5#�o��NrpV-T�ة�&��N�uJ2٘o
�n��}weO�F9�+��D	��o	��7�l�w��w����^�m뉿X��w�l�c��/|�ף�U%���O��G�(R���F�~<��C�m_�����f�x!���ŘqX��ot����{��IV2E����2CW��K��>+ll�5�wz�s��].�������]~.:�Όz;���7�>��ϙ�Ȯ� /\���1�P'��D���)ϴ�ugT���P��SS�[�飓�7]U�uR=�?P���?O�����w�j}��2U��}bwL<t]}��D�
�\��N��>������yld%U�q��x��jǫ�!�hu���P��N�f(����po+ؘ}���UGNKG����7_�E����e�)χ3�����T?Fpߌ��cfBZRV{����9��5N�u�Zax�{�0�����ix��/��+���w�m{=��ܡ$Wn6��E�U��9�:=��:t�/"�EO�踊r<���|5�
�I;�/�"�d��5"�;�F�;~+cח��^��}r�Y�R�ρ�,\Tϑ�C<��{?R�nz.��1���IճQ�����'�e~�j8rN�����ܓ�u=/+;m���4��5)o'���
��ɭ!������#���,��J<ƫ�|,�:���F,,�*2qz���@������T��l��-ٞ�H%��̦:�p����A�m��B��2Ẁ=|}~��?�=�������׍I\f<�A�L:�y}��7}���s�fN~�]���G�O�w#�D{�=�c�r^�mK7�K��4,��^���V�@��g�d��CǷn��NG��9���7�U#m����{��d��;��}U�5W��v>%{��;�_I�'��P* z[2
/�B�m�[�i�3�+���#Jɫ9[��`��H����
�ޅulեT'������:Cu?J��������0�^Xf&�����]�n�sh����ߪ'{�w�A�̳��Hj�
�N{�p�۴��G�cL�H�t{���C���w�~g��ώzg|K���������ר�)���`��Q�J�R.�O�||�8�޻��p?B�dx\&��[n�O���o�3q�S�e��^���d�"eQ-ō����u�+��Ǣ%un��+&�exrSRm9ϡ��`sC/�p;NY���x���ͯ4��e��zF���7G�}�8�5{yp���k��7�b�hz���x���3�]�պ�j&H���f��A�Ej�-����IJ�
6��U�7f��
���x��L1u{e	��n�R��ێ] 8�Z:TKZO6�@�Ì���etˊ�d���FG�VP�m\���q�`^�}��nΪi�\v��0�׷���c��|�)F+6��)��ÿCt6f� �G'�F����6K�p��W�^�\<�M{Lyz���\�^�{܋6�z�)5��Et�ޏ޾�~�9�Zs�������P���(踥?�ۍ��w��G���6�f�q.��==.��/׾9�^<���Lo�Ӿ8Ne�^�/�|-���5��{oZ�n�W�]x~�x���U�쁎��ҷ�X;�D{�H\o�]#B�K����z�<�N�['�~�U�|@��T<@�@Tbt�魏e1��<5K�A��P^O�&,�2�����d��}eTz��FG�&zU0�z���O�����9�^�����P{*N����pw��6��$��x	T;��e����RgM3O�{
�)>/�n��꺀�5��.�=��_�d[���:6���A�~
P5 �����S��s������Rx*��y�R�y�,z>^�~G|��Y�T��ݳ�$��td���J��}8#�9��zx��Ղ_
��޾g�����_�l{Ը�����~���93,� >P$�Fz��vɼ*g`��=1�9��wK�����T������CpR��j��G$�ϟp�2뫞���`������4���Gz�q��ԧ-���'P�ӭ�C =֝�dJ*��86�8�)N��Ϟ���ؔݎ�5��7�ʼ/Α�4$�n��Wx;;�纏裬�r�U{��팈���>�'��Z���p��>}^�q�����7o�����GČ3�z��G�&����Ba���>��� }���{�p{0z�b�ʾ�b��u=k�
����t�jnM��tVԿ�izj;��!*�n1��2J}�
?_�;�b�ױ����X��i	�S�G�F���e��/֝a���c�7<�c�~E$\ޅ�w7�=�W��O�N��t6��l�GzA*0�Z6�9>ӃiΓ��o"��b�����r[�S�;�/]����^��_�/N{��ido�+���m��� n٘�9��l��.͔}�ޔe�z6�?e��2S���z_�SCܧ���=yT1��wk������4G,K����:���Zn��*�� ���+ԼF|�5�~���{m}鞅�z6��9l����؏z��4�*8�Ο�҇Pcc�ъ@��I��0���R��NQ��=�Ww������z�u2�ET�
	��|�.)�f��x��N��B�\mP[���Y4�q�땨RtD��w�}
��Av]ۺ��n������E��/�eY��J��㲦ˬ�*Wo[�X��ͼb�X�S����bf̃q֊,�s$�2�n�X]HÎ���4{z:�؁��u^���"�=�V�j�(��'/�dz�=�Mq��\i��$Pf:�bJ�&O��v���d/3]�}��kczۡv�1ahr�z=�|zߝǻ>.�C�9EG�*����~��|�)�v_�ԡV�����W��C�?^��9�=�{��������Q�v��D@嫍o�}1^��<[�����uGg�n(����TWD:k�;^G���Q��ޢ7�T�N���Q��� �;�\�r�5>������6S>��0��Bިw߭�����t��A��{Ӗ���{W����n&��B���WURP��I����:G���Z|3`ⷄ����o��	u��白ۊ���<F�d�����<b��z�!���b�\�����f�%x�}�Q�b��֯�����^���ͿY�O�w���~�d���7#Pz��XNx�o�y^���f�):���#�����Drwr1�G�T?O��ꉳ�w�jB�Y���>���|.����xF%�]����n����P�ۗ������P��ՏWO�do/mȽ�䏉�~?�q2�R���wN�Q��3�4�z_A�[�nwW�GN�W�V�A�UŎ����l���_l;�ʺ�������Z���@np�{V[��2�"E��;v�K���!(��R��iO��xx�Xվ Ժǆ(�1�����Bu�O�\̎	����w-Z��L��૙sse�����1�T��+����IQ�6����کã�38��lD^�j��ҋCO��ߔ��J��d�_L�MX��H�.޷'�˹���7�x�]x�"�R�7,4"�-�q���S�gN��eA���C��%�1"�'=��O��:�47�&1��ʜ�Ӻۏ`^t�M\v���vҹ[��J���T�^�׷D,&�̭g{e�O�����'o3:�P ����������Э.�⎋I4�C�:����[��](��������:�e輔�jФ��%  e��g����4t������� ���l�+`�����x��p�i���e�x�GuVb�ڽ*�۷�7��j"%8e�9IY}Y�ᦴ��6�嵦��f�_E�}��4�Bu<�L����\�gp��o�&đfL�t��y�{�A艍�!1Q�Ǚ���[o�no�Bf	�$�u���&�����}E���q���{3,�4�����,���w�q���.���[nm�Y����7Re��&]+HiQV�K�h������A�n��'p�(;3[[��v�6��RZ&L'#kh�����1ʖhK8h5�c�5��}�B%j�u��60\���凸1Iк&V�H�������Wf�h��#X:7�M�Vl�y�(��u1wX[����5�'Q{��֑�m%m���n:�ʾ˼B��L�I���ʡ#CM'�&�E�]Dm<<4*��R]G}9K�
�12 ܜsA��h7`\߳u�b�;����e��8@Z�2C|��n��/�w>0��ۡBަ2um	�ҭ���$Zrn�m֭�z����Yr��fQ⩡����.��_L�t�"MEyB��7����,�ed�դ�E!�t��+���E����!�ehc)���R����Ɓ�:bwK�X�F�X�a���L%xz�u8H%�d������}GC:=6��+������v)%�`o%9[�*ˎ��:onS�Юۺ�&-�rQz:����2է���7-�&��ҵ�y��j�2�2W�������[ �"�IYm�x;�3N���VI� �5��2ڤv+����٤�简�6֥"5�r��ټ�_5eXg�Sz��@�Aғc[i���99��X-Ţ�v��B���6��L��=�0�o��1����Z`��
�ۭ�ҬP��kMq8��F5ҌDfi��`:F̛ǜ*k�|�IԞu�f�Qڵ[]��a`�6��ɸ�Ͷ�X�ž˝I�uEׂ��
�@�"�0�\�����
������������1r���2��r#,�jb
�b����)����� ����  ����,�fff*�(�����3,�c1�*&��,�*�**X�""�)�Y�������������0�2�""( �30�*�����

�"��"h��*J�����jh	��	 ��*������i(����
j)�����3)�&"��b�)�����&
�*�J(��J����"(�!������d�������b��j����!����b!��j2ʠ�il�b"*(�	(�d�"i���������r���&��*�� (|*��ܳ�q�k����(�ݠ˩���W$��E˰n�B�e4t�OkUxs~=�k!{+pi����A����6���S�V��3�o��r���A��NJ;&�a^5�ֆB��iL�w���U�]~�����ڊ͘����s��=G��T!��Ҩ�`�iC�:���g���ʦ� =��d>O���q�݃��I�G�1��q�6�����	a�+�0*�zx)>��b��)�,~�_M�U��I�s�;>=9�;��@\�#K��{�^\wd{ע*=�nxв{��P�O�]�t��ӫ}�ZВ��Yp̅��o� ����O�/�8�]!��#Ϯ��$�0���m�_/V�)���݋S{幾���7|���A��U����uG��޶<�y(8ܙf�N(�"�����*N��a'�l �ǲ��n*g�x�Ƀ0�_�r<���do�q�����0/��	�y�\��ݞ��Β�H9�<#<R;Fx���ۊ�Nж�|Wt"�L#T��xTq�wqs������WV���:'���@�n`?��`�5�o����語���|����w|я9�~��=��ި��]ߍ�UR���A�/jci�o�K�<�b����d��sOb�f7⍛I^�M��^�Y���m�F���e�f��]̲�b��N�|�{lQ��;!��s���uJk���1�4��9�*����F����x-�{7=���|���ݖ5�,�^z�|���G���N	�$9�*
L�һV	�O���넝�1���㞙�~�F�����93�;�!��?�
�w��@�9�}%�.�Q���\l����Ȋ�]�۟���;���Q�p){/�d�������0��Kg�n��}��r[9W�T=5��curo�zn��q�(y1����癯�����{�|2V���n�J���gg�>�[��>�᥷��������'w>��}�z|T�q�]�%.�b_�+��Hɚ߹���Z��e�_���H� ��w��5^E��q�Aܥ��hEy�J'�{2�w�T~�����]��Ŗ����Ł�7�p.?��\��n5q���y�}M"}�g=�c�*�p.��?Mx�����ݺ��pfT	�*�ns�U]�Mx�u�C�Ϩ��m01:@�U���|Ψ~����A}�}t�}p�~g�'�b}�ꎎA�i�ڏJ�Gb����ڏc]Q�����=�ǖz�ۏ<�7�Tn��@�>�6��T�}AQ�N�Ih��u&}�B�ȭ��Q��XJ)�P�H]�߹	���V�~u����-�b����2���R�{Z�9w�"�mt�U�$���*<R���T���c�7/Ƽ�[�|a�G�'�BmM=Ԥ9Xd�WY�$��Ph�^��w��2����]t�0�lTr:.rw�[jG<7�g�2vJ*�W��v��(�>Џ]!��:KeJ�~UIF2&}\�,�F�z���p�f�9E\{��OS�=�ĳ�������F���0x
P5 ����a=�~&�I���خ΍��?�POGt���W��C{�|}���s����0����n	��c��[ ,y'�=3���J�u�Y뻚�(z���@mRߩ�n{I���\O�]�M/MK6��ױ{�]z͜�%o�����`�[QPK�o>�d0ߕ!�L���ztx��Nޫ�EOs~0'�7^V��g��Dͯ5KW��3$���H�'ާF�㷳Ɩ�w�����Hg���G=29�g�2hw��9����o�]����\���?���*��LT��v4�5�w��ڻ��L�½���9OO���W5�D���@r��2��,�Uߜ�)��u�P?��`�}�����Q�,	w���TfM8�G7v"���%���}�]�7��U@ه�6�;��i�9T�j�q^���劓��ꓜt:ʫ{�T�#"5����f���z�:��A��o�+�f}��6�����+b�J�ƙ��źT��k��ώ0���{pQ�}����dڱ�=&�J�|r��lΙ���s�n�
�^�",�ԓ�����|x�z�O�Y%�!_�z��3J�R�Z��գz�7���q�3/_}s)Dۦ�#���]��﫫���s���xle����T������d{�{&���6�m�������H{������c�j�:���L�� �^WzW�_:�j_�xtW�7�T_f㽙�V��9s����8Js/�q^�\q���uTG/R�9�����|C�>\��EY^�=~������|먡�B*�e�Qg���򘸧!��|Ww/2Hub�G������,�F�rϨ������{�
��qҸ�9�����|�T�|1�`H���}j�o�5���O�Y4=k��`�O�{d����q�ϋ��\�u$��<�I���w2�ؗW�,�g��s��Tχ��x(s��ўs�{#�u~�Bt�?_�=�$�[�|"|/�EH�[������@�����>��ч��=늸t�!�v��?Lg����P�u������̊�)n�Aoz�z���� #$�!)�p6W�� L>5z��C~��}���fuuT�I�ȫ��Q��\�p>���m��uU%��RZ��@��zxMT�>��B�Q�s��5��xxܾ�GNe޽p����Ӣ��,�<Q{��v������4�:�r ��rݜ�\�b�]���Z�޻*���שH�A�l�@S����M���-�lC���Gs�$g�%�M{�k�����ؓ�3p\ᨾ��j+��{�}�Y����ư
~��s��7
d��U��s�4$u��/@���ҭ���]$�=ü䆟UQ�6�d\{���j2)��+��QB<���9	.i�MUT��y�,�ī�=�l�M\l�Oj�r�܋����~�����05{,�W����=�__��7'П��4������yqwz��C�P��ՏWO�diF���(��';�ݷ>���="��:$��p$F����𤾸'�a^5�ւ��a���x�W�x��:����f�@�^�O�q;�yc��q�A`�����D��~��=�놦�6,���s��; �w�� �x��n��>����~=��ڞ�N�����������NG�䥻H�uHʍu`,����P��~����3zߊ�^\wg�z"�<��'��� �Qk�Ǟ���<��K�p���Et�\�X7� -~�	^�?��<�����~}t.�zpy�:=YdF��ڍS��P��x��RS>F蠽p��0�w�x3�p�x�D{�=��1�*^��P쮳�S?L�5$��e���c��n4�V)2�)v�5(��Z�`�]�U�@]^	�nrυvPK�j7��^&e��e�h�(�+cT�[�\4��Wx�d�Z��Wf�hM��ҋ8���ӟk��a,����ݰ�* ��W�q���K����A�������,a'����}FR7S>�L����G��9��P��'ђ��a���������yv�8Β� '='�����Ϩ�㐳�qW��=���{dz�$�9��y����F�q��F�z��~8'��[���7P w�	�i&|n��"EL5|i�y�)�Ы��c=;�����~��'�=w~4.UK7��	�/t���omF��e��������TT~Y�G�w��}���zg|M��Tl
����\:��S$5����z7����	�{�ܛ����W���*"7�z�[n�O���o�7C�\����jA��s�.^�>�w��+�}%��^T==��c�uto�s����}{FE�aH�'wb���Nc��n2�T%Y%\A�;8�W�t�z|;K�Ko.r��4 �������S�Ms��K������Cfn��P�91�������xm�K�t�i^+=�V�wG]�߻uw������<ߢ���g¹G���5��]��ŗ�%�9�X7�pa�������K�4ȭ�[����,�4h�	�����rB'Afip��&��@wZ-t�v�u p��<��6�S���ު�gtT^��h.��>�0s�0�`���ݰ��n�6�9"�13j�V�ǈaY�׈=Դ��;�%�R�~`?�}���S�S�J�p-�^��?Mx���_i���Pb�݀ו���a*N�]#�y�������t|<�|���E���@�U�y�ln�������^3X0�$�={��*�.[�&�+5]FϦx�9���
5������=�Ǘ���=Y]p���](*=a�*UbA9K|����]QD�{�-��:�>�tTEtσ_�E=����q�.�Ny('/����}�W�t�kU�]	+�x	�U�e)��Jg�M3W�de�,:���w(�V}��>�|uG��=��x�4��[RAu�~
P5 ���͇���c�TxvR��8��W��|�բ�S��޶�ǔ�*��+���w��|y�:3�\w~���&���f�y��ڞ���[��B��ա�9�Z��.&����x߮��?�v��JU^�1����t��^���(��{"��[�C��9=���ф��ՠz8TgJ�OE��42���35k��}ꪗ<$�#Ď3ޥF�;�&����~�~���,#U�#�V~�]/�R�f�H.� �O�U:��ϓw
��-f�ь�xWq	��FK�PǚΜ�S�w��NVӻ&�.��s��P��ZQ��(b�oJ�Ƹ��!�<�F�JXw��J&o�e�b�ɀIz��6�R��Q\GJ\Ts�h�w#��`�"����'�Ь����y����S%�hd��
���;F��5��P����מ�Ǹ���;y�=Ïy��[&O��@w��� �H�2��N�c�}.V��Z*�}Bx*������ʷ�7�l�����ˏ7�0���%���y��*8@�J߆�>�Z��ڏb��ðgm�]��,:=]+ǳ���n�1�ʽ���=3~ٶk�޸�6��u�#�I;+�|�1��o��x.�F����h�zt��c¾���cS�"�/NyMR���V�p�M�=�'��ܧ՘�[����'t�8V�;�ʭ2�Y, ���~ꗈs>�{v����=�?,��0�������kh�C�'F���L,��V���y��*�ڱ�&a���ef��Dz"]B��w�����󮢆^IE��	��|�%��Ԍ�UL�:��ٜ�ڭ�^>�7��@[�QO��Vz�ǻ"�F�~�Ƽi
Ð2��L�6��M��F�n�ſF��[^c�U;���M<�޿�����Q���q������h�l�KF���@-�z���w��ð�h� Lwg�o��Gڛ���:�m�"�N�g7\�lU�v�G2-T��E(�'	R�WuNre���M����˾=΍�HIr讀
���8aڙQ�а2Vn�0��t������zj��[��v�;�x��a-�i�M�p���7���;S(/;w��:~����3��>=q�'M�_�=j��h�9�YGg*�u�f����@�T��?����q3M���\Uæ��;^G�!���r�< Q��᮪y~�(]^!{�whW)���d ���G-�
/�V	��ouCN�m��C��	|$9�es�yu^h�}�h7��o�kƶUIaI-H l/O
���g���︊���/��{����s�����O�����<k ���<d[��QD��D�.{ƀ�^��>�V������tig˕����߬��@�11pߨa�{+�o�S1�Pa���F�֯Wg�LzV��ȧ>�W>_.���ϓwr1�G�S���C7���F���Wj�)��{k�<�͖��/��θ�aϧp��n��屜�V�C�P�l�u�^��5���L{�n�0��9(ʑ^�D�@��6wj�Y^�!�8p/{}lb��i�}���n��^����M��ULR�}٢߶���)�:vϑ�����Օ\n��:o�.}��� ���f�fj%���	8v7ԟ �HSvN6���!�����c*�9�L#�u�P��R4nMyKu^�$��Ja����xݡh���^�/WR{�+�����%��Qr��M8(�I홎�N�Y��!�6���hu�[�s`j�j��N���v�l �ݸ�r�ٞ���~��ȇ���׾7��wjxd=��n&X���NQ�=�N�Y����^��PP�X�>���|�������Vǯ.;�޽F/|������pe��~��]������g�NE)�3�<W�X5�P��g�l_����]!��1�Ϯ��GnA��
�4gz�d�>2��IH�Ez@M�Ha����Ͻ�}��c�+�Ǒڸ��,�Z+`;����l?@�Գh�J�1�$�P��2�}.|8�&�Z��9R|穘���/UT����N=���g�7�/o��gIv� ���x	�%Pcų ��[Ƿ8"�ut�ur���yT����N��w�r4��=�#n=ul���p��]DL������҅tL`�[Z�T�x������������ϝz�1��޿q�~��߷����n��� �HH��^L�#��s�n��{:懾���]z���~����Y��9�z=�\t�g�*��ׅ}�Ȣ�j����ܻS�o�<����ѿ��٫�f�����'DSn�����TX����>�W��_�_�TDEqQ�_ꨈ��ʢ"+�*""�������"+�ʈ���TDEx����"+ب���EDDW�TDE��"+�U_�Q�j����DDW��PVI��Z�c V7��@���y�d���GF>K�zP(�H$�$A@P� � PI@���uJ��
�T���$�*E$�B@ � ��c�@($P(�J*��P ����J)!@J
�:�N g.�5���B-�@��2$�*�H(�1@L�K`h+�vPJ�Q�*K�@  �(
Y�  	���
��J:e)e!*l�Q �RD�LiKmV�Q2Q�T@T��խ�MT����� �٬���r�i��6a@M�kST�3�.fʩ�M��[*ؔR*Up  ���Pʹ���k�k��R�-)�M���l�jYj��m�v�M���L��(ZdD\ b��cEh�bL�j�5X�e���Ś�3���9�mB͒�,f��
)P��9-ݎe�S[cTQD�թV�مV�fIH���,�&V�hV�	4��Z#F�d4���$��ʔ�ZZȳb�[b��2Y��"���e��T.��ڴ�F�SBF�Q�kl�e(�խiD"���*@
� 44ʕ%i�&	���i��L"�������   �I@&D��yF!�i��G�h�hO$"��	R��'�C@@�&MLL`��I��M&M�ڞHy@  ���n�μx�|1ÎY�c�+�cmu"g���t�����RY"I$GdBDIr0�)�U�q�1H�:�~�*~1���
�!�և��
�$<H��:�!!I�b$H��
��2�p�e����`S��~=���I�	4�i|�r�3�iFt=����M��?�?_a��,/r�~�?�*�+	n����؝��0�0�S8(�a0ȸ��7{���.f��W�w[����Lr�=�lY�^؀�ĥ��E+4�1j�{�uV�i�E/�۫U��i��	�����qᢶ���p;�vF-:B�hk��5��A��А�w�Y�w�	V%��gN�&c�M�k�e�[� �U��]�)˥�a�j�opd�n�+KjԧXe�B��i�cD@�+r��؊Y.�y�m2>X
��B��j���Ig3wJ��Fu�n� ���pl�Dc��7��LaW���ot�z�3A/t[B޺w�NS7n?��ښ��b�hM�#��86��ܕ6,�k-m�]]���ū	"˃s)����X�������eD,d4���N� ��U�:COE4z�.�:�Y�V���Rvj\��K��üB�&��A�+ijI�kځ��jܶ�b��eaW�!Y6�Rw�3�J�D��7E�E/jk��Uҫm�5�O.[yq%<F�����0u�����Ix����&� ��VVb�Yߙ�̡8D�2�i����]�
���A��ʹ_Ҙ���1���ڼ^�G�ӗuk��r2~Kv��ğԲ:6���n�Ԋ5�]�L�=f�o:�m� x��e�yMd��C���յ&��n6m�^��A�W@���4�NU�`)#1�M�w��]����R�����E�D%Qխ�Y����4�7�q�ցoAև�� MlJ�v�@0��JQ`��#3r�حڠ�K����m1u[�}�� �E鷍k�= ��h"t����9�k�Q$Α��q���X/6��^���f�on�
���{��,#�S.��R�T���{%[D��vZ�m�U�v��,�t�a����ù����lF���Xu��f��G�1���e��`˨�#��,��-|(&B�OVb��s�w4n��X�)�"����q�=�M]&o�L�$�p�	��e�KM��bι�C��Ҷa����Z-V7�"�h�Œ��h����clHn���ܘ�e�8D�2�lEO^��^]űHq7�Ň��b;��0QO.�7�] ����crP-i����fE���
��4��B���t��jJ�P�7)"��L��A��
8�dh��F�l��U�$Ry�Y�ًN�6��%M��@�{o2��Q�(k�G#��l��,�|����)i�4Yn��׫i�M_c�I����Y�f��ek��3a&�L��-e*�0j��%�u�&j�V�,��N^c���(�������5y�aD��͆]+KUl��7-�SoA[E�r�����j�>j��َ�U�E�w��dh�n�'�śF^c `�b�)WsDu꧕���*��,��̍�ǵ0���Bӗ4�Յ�e�Tml���������Ѽ#K���N�*.��fRe��C�K�U���l�c{�u%tqA`�0������a76��5`��d�F}-B� س>c�h�u��qݖ6��R�N���(n�S2���ڃ�&���̉"��b��j��I�,^��X�xf_[WO�m�]A�'�L�A�<��5�e�T��Y�4�/e;0�%�s6;rQ֌W.��gw�R����U�K�"��wzڃK�ì�+��l�0�3m�o (�ٚ��^hyS(KHHJ�A�vY�V��#0���(�vڀ��ʈ��kk�V�	��TV�^���ܫ�#�C*�� G���M^^>�b���k̬A��d�5-�2�2\:^���K9�f�Y���hcQ;u0f�-2 �)=��nj/u�en�6c�v���,Y�;{L2ސ�D�n`���s�L���g.(j&��Će]�Jb��$ю��ݚ���ZtJ��$S������n��[{�*��V��������M,�D�
&��ڬ��u�
��T�����u-�OcШ���Pm�D�J6(-��rKJ�M�۽ŏ"�V�96|�jTt�
��;��scXg��K�ҷ�)Y@�v�2	��p8�Ae���ؐ�e��iS����oF����BN�c��f�F:w��a��Y
�̆+n����b�w����S)�ikI\њd�բk�C@廧�u1e�[��)Y��:��z".���l�՝.ͭ���'�;9CkqQ�R��2�v+cm�ɍ�J�����kU��®�u-�VW�R�kk+�����`ۚ��D7m�2A��ޛ�*i.��U�c)���A����IC&:с�L�;yt����U�J��u���&mF��IG3lP0)���� �8���`�S7v��m��k�k!t�hړ~Ê��e�%aڣJb�vu��u�uz�����r�=i�$ևd]kV��ge����润T����n��.pV9,&����0�ospd�n�7��S����^����ㆅp����h5zѬ�F�S��C��ƈm�Ů��w$�O.l�NZX�H
i�
6
n,4�5Y{�i�nLD�G]p����LFأhʽ�r�(,,ձ�*�ް[2�����3cW��B�'
��дF��-�͛Y�7]���/�4J	��)^���o.Q�vЅN�5� �wf���Хw��W����^`�yw��qrI�ܗ��iه]^Cr�"�
+I擶�9�6�}�j�}�Bu�{���Ҝ�k��yB��c�ˤ��t�`ֺu�Y给cN��|I��L-�v���՗ɑ��V\�ZN��)G[��Cc���N�::�Z�ص�i��/H�yi]�>@W.2V*�{��n(��ڷ�iU����7�����b��r�dV�[C�н�+�.�����`��2��,U?�S�°H��z��t�&^[gt:٭X�7Q�ϯT�[�Q��R�}�a�m�ڶ 2�c�fo�J݁��BM�k!wX��B�ӎf*�(��%M�W����2Ht�e�Z0�2�ځoʲj�h��v���`�p)[�V�-�T�8iғ9,E��)��i^ ��/e�LX�i��9D���j��u���+Oc%�J\��1K0���	�E���U���9����i����
��s�o<��#8��K�� e얩$"�/"�D��(���kK��W`Y����{N�&	z]��%�S��������ܫW4��V]��s ��݌pe
յ%Ё=[�7!�(�����nk�@���-ћ6;WqF�Y�$��٘skh�އ�Q�ٕ5[���I�ތ�\�����W�7��?����J���
&v�&9�M�#1?��?7��z�n�G�~y�����(q�&�o	�F�=�j
����)���ِ�Ļ>���`Ӥ�8vofȤ�;��ݲ�`\��R�]ud[�T��f<�F�w	�wZ	��xZ��y$�
H+"Zڥ�z�������!��2zʺ�MR�{>q\��X<���T��PT�m6���Or{�]^5�49�krl����° v�XD9.o;���m;�GQ�
�`�%>�u�1��~��wrr�ڬ�Ƨ)YR:�EIe�t�4�0~T+�Vh���^�f[�eMH͝T��#;hXu;�v����}��d�8�C>SVL7��ָ�)�5��t��)D
5q%���+Wl�3.�"\��pA���1W\(B.T�t����/sA;��{UBU:f�9I�/��/���镩��W�	��P�s �4�����D�wZ�b����1�g,Z�b=l����b�,�9� �
eR�l�n+T��ۨ^R\UE+�"���0��M�\*�+:�6!Wd��?D�WP��j������:Z�yr���tĭ	wH�[�F�E���&�L�s����`:�'L]��t�N��3��T�t���:0ED�Qn�TBgY0���©i 1��6��N�7H����i��LR�W7�9��+�6������p��m�B��j�*�*z+�!SN����²�*��̉'�.��y.�M|z�k{��.��A��;����ywc`��lb��:,	k{�}6l�l�
��a�*�d}��5�sLFl���� �|<;��4N�ѽ�ڐg��Ks�	�+w��u�9���l;��osX�Wj��n����6CuvU�]�6�-�^ꕕ֭�@�(P��vn��"k�汦��v����P~rcZ+���̞��v�s5���	���CU+0i��5z�Y��T��˔f��V�g�'���˻("���N�s>U����ؗ���΂w���T��^{���};g�Y��3������bZ�T��TsX�V���E�Y}z�9�`G�i_R�A漳���Ý����d;�5�+�ݤ�/L�|\�%̥/A��Ŝ�hI/O1V�m��y��t�|�����<*�r�fg8nj�̓\��.�M�S�����W���[����IqBfZS��ٹ6��pCʃ���3]�F$��������:���y>�9ɩ�Kfн��"�M�[m#;LU�G�G�4��	�tX�gC��O3u�%Y}�yS1��.�Ղ+V���u��-������jR�Ng�gnj	��8�C	+e�ԭ�*�]Ao�wmJ��A�����iF��,��)�L��nZ�!��6*!1`���}�S5�F>s���c�&��-���:T���`JDd��\5��hUݼ=�(0|������B�e��1���{���!�}\z�T�:r�8:$::#پh!�:9Hb�ήS|;%��/Zۂ��z%�Pi��9����/�XLސ�e@��¢����kͼ�Σ�˳wR�N��oZ���f��:���5��)���V�g��l]���8�cw�!���u-���0�m��0��Z�L@�Reew}�rK���|�4u�x�\q�w���t��ZVrV�q%������w�:��ն͝�fF���Nd�}6.�k(8�Qw�뿢��&��s(����z;�v�yum��6���8��Jl�bɫ��6�N����/o�h�ѤT����2�<߬8���i-c�LG5��ֺ���*Ӎ5��:��.'����_E�/e�[+����&�	�0ao��ڽ�xV�tΓl�� �[{�b��g%l8�ʽq��pbݢ�!9��v&��L��g� ղ��JKk��gqf��Syt��di���Kш���kK8E]�rd.8�����L�%B�8	AJ�4bw!ʺ�Om�2]�V�-g;Ƥ�����}�|�8y+��Ucie.�tW�lt�+k�$L̵�H�=��
�����O�Fg���V�ů. n3�%=��ܖ�)���p6����;i�,fNN*#�Of_q�U���j���iJ������N�3A�otf��<'��TZ2��i<�;��f��7ui������z��o�SkC��OV�1�EV�wh
��)Z{��U�I�42��-t�����\W5��z�CsMY�w֊Ûձ�˓=��	�?N��ʍ�Uե�7L��s���\fV�G+;&	94�r�uY���MlӀ�{��k�Sn�P�z�#CW��=���&��>郟+��_s�WiJ(ICx�	�����A�Aa�f�I=;�ћ&\J=Y{Mu&f�ZYQ�(d�*R�2�:�s3��(k�v*�#w��ӷ&���r�������ɷ�rkJ9�p�"ue��[zc�sY���(��3�p�y91W�i��u�-cY)2򳳰Vn��58u(2�XhjX���Ld��z��z�.��D�ǘ�����9���W&��V���Y|�>V���^�H\��o�3��,c���!»�G`]t�8(��!�V�kiq���wkv�P�9s�n;=���ڎL�74�{�Ҹ�n)of��p��d'�]e��@��N�9 �#r_jrI�I$�I$�I$�M��7S��a����"RwaΝ:�K�1��-*ŵ��b���2�ސ��[�!����⡗MG��B�]$�f�l��
D�v�����4
|]�[�F�sew'�p�ݣd��p[���:wi����n '6����6����Q�ۻ�A
�+)
�{x�w��  ZV!L0�Us�Q�h��#X:�Q�p���^�D�z�P�$]wFԇh�N�u�GU�cP{��Op��M�2HT�|*U��Y�v���2�n��6+ "�T2�j�4��ٷLE�l���6*b����j��tU��)�!JB�$�������B���6�B��Ňs�G5|��p�f��V�_ ��b��B\�u��	�c
W�-�]ܪ�P�s��}F���jY6�=|P����J5��3�ت�kN+����P�
�[J��l����CEʬB��yw�,�ؾgE�CA���-X7��r���W$��E�`� ��:R�*���B�ٮ	�Xh�Z�]�V^8׌�|��^��ncJ�\ڽ?�٪(ov�U1¯�����D$���) C��KG�8`��
��tBh���%�D3|ڕvy5�W�4(���:tt�}���I]� �l:܎�b@
�KZ��`ѭ*�ފ𪶛]X�W�V:4�������i�ݲ�v�ݞڕ�V��8_N(�$I�-7I�5i�UVg�!�I BO�8Ο{yҭ�����Ɍ`�������Z�[��3z�V]!O,>x
X&N�.��c��������"�`�t�`��,v��8;Mtp4-U�<x�1��ť=�]N˻�z���Ww6�!\��Ǚi:^-3\$ 42�m��\�����߇Qm��)������)�6�c��JA�u8����6�j@˼�p�Z�@��M�UE��;GR����a��fFZ���vN��n�����L��*�m�"]�]w��sK���lx�qu;�ʌ��Q�dRh�4��-
�&wb�(�n^w`9x�+�:+zֈ0b��VB�2L1��T�8wn���F�K�m���SZBh�AbᲭ���s��@���T�S�U�Uۘ��J����,�4j�P�}d�k�ͻ�4(�tϡq���|~��hA�	z��$Q�r��B��)�R&twY��B�@�t3
p���t+�<u��*	H]�m�J���h�C�ӽBm7DP�f^[q�1˼�|Q�Y��c�K��h��0U��[��YM۽��Z��]չ�2[�9D�\�/���i�P�;��G0��݂X�����Hn#N�S��%P���\Y�9�U�y�2NpJ�(:�Kty�#ĕ�8lN��5�g?�]�����]|`S/�E71Û�8]�:hp-�l�k�p�&Mv�#��A7A��G��f.�*^��:�]���ù8L3��
���+�\f�Y��*��I�桑:��ċ��Tz2]�- ��}h�m�=���u�U�Ô4����KcF�2]��<�˧kM�y �%U��u���ȫ�l24�c�w��k(
g]c��G��(*ȮeP��q���Y������(�k,���[ghFyӵKoWS�f_T�i������ĸ^V,ͪ�,t�w2��ҢF��Q+���Y��u�j��Ma,J�M*�d�b����hR��.Y�i6�P!�KUV���n?��ʭ�_^=0��P�:3NQ�k��K���(s����Q�%1KV�x�Wu�%���ܸAg�r�����[�[�-��CAP֟��$��D��
���@[G1G�}��B�J�t;�[}/b�kfr�y���t��$F�!��Mwݕ�"֚�ҳ6�Wn!�l0�Ғuv
*�0a9`��>}��q����� orBq����Z�s#{�f��	�	*���)NTm�f�L)n]�s��A��o9��F�^\��ج��*���̤퉼FK��M�E�l5�XBٽS����2���lZܹ�����='S���C�W�Hݜb���)s>x���Vt���b����	�T>W�bt�un�����qSɶ���7�<Nv��u���Y1�uҤ�tWeC%�"�ЉЙ�p�f�D6�e�f���hR�)��[�-khTN
�ѩ7r��.�^t��P�v��,��F3m3��L�T�hL�2���c�İ�V�@�Xj�e s*?�&����Ac(�й��4�%�]i�л�N�^�4�l�F�J�����7M��A�k�U���GN�xR�C�p�j�]Û��avʁ�\j��3�+P@��xM
LI�
#�wAN��dB��+t�{�q�.�j� cgJۛگP��#8U�j;)���\�ϡ�F��@0�1wr��O��j�b�T�F2DxL��bVrBHQ�C�W���]Z�Wn�שU˹X�\�#� �%��T�c:ӧK�����\+"ŊP��Q2R3k:��Omb��@�0ՓRV��ӗXme�u*n��@���:��K-Ҵ�8W�v@�B����R���.k�]�>�{������'X(�F��vkY�;oD�Cr#�a؋<U�w��+]*So��]2�bb���ܳu���������c#f�mT�%,(�������U������JN���s�xc<�+�͙�(�!9�.�+��:�]�1X��ȅ",�],�
���/�H]�s{���U�}�h��Xd�苃��Mp'B�v���nE��tӡ�\5}q��t�Pm��Jmgװ�`��wή���m�s�����[!`n�s~CS�«It[n��`���+�h��k	���Zp]�A�ڥ��m˳��캴y��Jh�#ifS��+�+�N&o���&a�E,���*���+2%��Y�g]�nQl���@{M�e�c��%iQgk�
��slԴ�(r��]Ҽ8x�YW�:eʻAV���lד,܊��X�H��0�
k���uu��_R%Y����1j�^¬W*��$���M��H�h]�m;fPba�X#�4S_/����ӈb���f[���
��<t ���N������8=s�s�<ߚ�}�
U�s�MQӢ��N+��ξ`�;������^`�\��:�1�|r�P��ʅ�	R��4�ĩoYpG֌ϭ=��Ў�|���n���c�-����y����ݒJQ� XWmKvg�n���ʅab��ąb���)���g�κ�כ*@;g�+X���LJF�ѬLL���p�0r��>�*C)� �Ҧm�Z�����i��;iPާu ���5��u�5]O��9��V�SUAc0ݳp���ҭRW�j�smf�g[��CI㭛X�N�v労.Q�k\���<�a�3L�`#x���X�z ��7M+��jY(U��bI\7�:��̅9���Z-Z���؝u³uMp��	<�#q:�f�+n�@V���W�	_]���EZ��� &�<+�
Uh�4���}*v�f��r�T�m|4S	�61%܁�g���`�q�nP�k���숋��֍����Ie���ASq���On:Q:xU�Q�,?��U!7���Yr�'Q�e�x��SwD7�T�J{�앨W;4��XU5�/mk���W�j�MF#�0Ȕs;.T���B��7j�"���'V�p��Ix��h]YV�u!�W�$�giQ�eZ�w
����*�>�L�䂗Z
�V�C!����W�u�P��o�4q\�[��蕶h��
��`��b�0��)#T~ّcΖ��j�R�,�����b�q*<��F��9��T�y�e�RБ��|�����Z��(�'[���MJ
�Iv��wx��.T�0P.��\fs2�=C8�BE�秺��z����Q#t�FbTB�������忈�foS�X��_����TT�@)B�#�%�<6|�` &����V�l'2u�?��+���e��Nm`��2Q������}�UW�|�XE����i$����:z�}���7��~3�{gjY`؝���v��7�Y���;x�����c" Vf#[�ѥ��(���ጎ@�o&W7��+�7[�TO���,s���w6+�,HV�,�I�u��37;c��`:xt���9v�J�ꀡ�nN<�m��Ws��&j��Iu�
��JY�܋�q�ޭ�W]�� �Wyk@�����(uv�-jm=��{ݔ��ⰾ�ΊE�i��S����̓M��.փ�N���������Q����'gc�47E��(��7#������IvM�zd$4��r�w���0H^�����E�wRU�;��{�෧KD�$};�r�ić�O�s��=�+<!׬�E`�*(�"�Fb��UQDV#rY���D`�,X"�	�(��
�b�UV�Ab
̉QDAETAX�����,�YE"ŉ����TU���X���Ū�QD1l�QX(VTEa�ńc0¤R
�
,�H��d�o�3�]}�����c�p& -��u�V�=Fl'��zf��b_S���.��������Ǖ���$���������B5	�D��+�x =�A��Jh�0��t��*��1a�d��9��ǚүj����&5u����1P�R�;�����2�S����qf:�K`��ͽ
ÑJ��܊,���}��Lӫ����_�=��9������ePX���Cƪ�Y�=��2��u�WK�
�D4��=J Y�~�e���\a��7����4U��~���l[�b����C�QA��M�LY���Pw@dM��ֲ��͗��x�Q�r������ؔS}7�|��A{���ФφW�n���ܤI��uؚإ��Eݢ�f5��g�0G���ۺ�OY��ƽX�-˞�b�6�TN1/o�&��C�q{іx�f����n����r�ȹ}��G��G����εQ���<z��Û%y(&�{�h��l���vs}��mJ�^��6����W�E��N�n獵**~��ϋ��a�G��H7#��i���u	��`w`�DpK�f��牒-F��`������>�7WJ�_QS�X���2��GIc�^��M}<�Ҧ�>)�g{Q�������a�(6m�v��Q����{P4x��*c:7"����c.��YHb��z�)�X�K";j�J/���13�U�`�g��獜�6s�q��m���M���e��?,����N�T��)��z����}[|�&u3ָ�h����o̽�5[��d�'iw	ĎFs$.��xVA�^�^��%B<^TN06�W�v�ٗ'L=�����I�@Ie\��^���O�D�&@�V�
�IRV���^y�^��|�s�TFq�����[Q%�q�u�zz��07m�q�TU�wW[����՟����N��{B�������9�¨J���g�S����1��O�$�&m�,f�Ϣ�I���+z;�gs9@���Wv�;�����8q�MN���h�#����Ɔ�Pگ�du�k�8�g�voQ��s���j����*��qg�=�}�4�S���6q�xRx��Ob[��XA���B�5�A����90�Y�
�%�fR�$اU�m�ѻ�r�6�r��s+)�Ӛ�!kY�%bG�߸3���Ur.+X�~���\��j>�hF0�1�������{���*E�ˋ�����(��[��{��u��=��b�Fy$���=��)�m-;���<��:�F��ڞ���Ne�����~/.(��tM9%��|<�]F.xazx�8|��rAު�W��j7�Cs�k�Qe[�..`�*����r�d/ռ&os�	����/�.Fz�l�Wq���b+�����]�\R�/glYBKس�� �̔i�+�L����fi����~LQ��b�����Z�_Q�A��|rX�)����CG�k��njk�v#:�5qe��O�׵�~KK�i����}u仰���i�eSy�A�@w/aU��{�^u����]�,7���>�k��H�����=�M>0���r�ӶΪig��<<	ucTx�����J�����u.�l���(^�-��5<缍>�g,����qE�N�Ǫ�;?M�G!X�ݳev�,��%Gἷ�l��-�H���,����^��.�i�w���T���(ѓ������0ז�0�q�xd���=8�j�Ҫ��q�&�m�顕�	�H��ni���ߧ��������:�2�}{��*~�I�<�n�;�*2o];�QZg����4��?3�ZЌ&���*�"�Z���c���&���;C����c8���ɭM=�t�9;��b�x���Ui���#��i��j�Z)ST�\e^2���q����ߘfn��4F�W�{}�D�6D(T��g�zH�'�R�9�9u�m��s�e�[���E5޵j��:����Tk]\f�l75��˽~�Y�"�$t����5��:�izfPx�ť�N��!����]o��ͳP�e�A��Po�V�Ο�Q[k�M�Ȳ:4���y���i�W���<ڭ\�-��{�Y���]����ҡ��z�� N�ͺA^W�Ώ,H�4:�Թ��&<�{؝kU7�W�')�u2�t����mk۰f[盵=w���:@�E&�Fo����;�,<ځmD�j\u��u��Ֆ�k����w��l"�uF�Z^늵��WKx�FvGMs�w���rە��9vU1 �)��{�T}JX��}ŋT�ԛ�Š�	����\|�?m�mx.��ϗQ��z߆T�ֵVi��Yh�7Z}ǣ��$�ls;��>q�x
�?dQ�_�+z^Y�ϙ-�^�F/���c���C<7���<3���8szr{6�U��6d��.}u�o����]�H)�if�:����kx��,�������hW�0[>���)��/�'y�di{Cm���͐�M��0Dێ�-cYkA6����=7�P������ɖ�^h�r*���$�X��ުÞuu�L�j_I�ˊĻ#��� ����f�MVb� ,��c����rn{:�W����x&��YH���h�Tc���[j�q�u�^l�����|�t�����zq��Y�/6���L;Gc[�Ϝ����nw4i�ͱN��.h{���i��k����[�h����m
\�(T`i>]�L�6���〱za��3xS9���7c�{�A�F\~^��b����&�\41�}Z��hU�~:�u���d��w�j.X�12c3z���U����*�'��.�N�u\V[���F����ݱ1�8���]\�/����w����PY�������F:��e.�Y<wbO�N��Ѭ|�{�����\���v��rs�w�Zq�}[F�J�\��*�Y�HgF���0nZF�x^�x�h��.��p[ݻF�9bs�p|i�[BA�א`�ʣ*���PX0�i��hR����d��5oZ�y�ݪ���#�]_Y�H���D-��U�3y��R�kx�񂉛s�[7g����� �@o.�:�9Z��,��r�(�kq�E�M���1偹S1��#�	������(=��Tf?��;h}jv;�	���ӽם�+5kZ2bcF�cw^��� �xX �����!oD|h�W��2��᠚�:��'�V)��61c�uy�
W�em��� ��VaJr�u�.`�Y���Ç��}�bN�YW� ��c��L3�h���V��; u�9��y΃M�s�f�:Ba�������1X
Yu�lkX���ִ�3=n�ڭJ����_cy[R�f�Q!�����0��ݺ'�(�\�a�v*Z�vs0���7�q&H�FέᄉC�N�q�ݱ��'9a6A��jۻ}yc�s�4�xٚ�*��Ӥ����̃f�8x�����}>������,&-�P�""�%B�`���q`T� ,��"H(
E�a���TPQE-�"�0�*ER� �"�4���(V`)	����*��b�#T�1��`# �(("fO�e��@�	��U}1#��*�lă���OZo��I�U�F��s�����SS5��ṛ�U�{��m��z�8�|���!1m��wG��>Q�mW�����_6���۔JE�"�]o2׽Q�3����[�Tih,*���M��-s�ko	�Hixyq�]�q�2,��U��Ｉ�}�.QQ�{��q8�J[5tWo|�CI�x�c���Os6����W��8��Q�]�/_a��y8������
O�L\O��cKu3��ݡ�0K��*LO�nuޒ���@nG`����@��'V#���sjV�S�h��I�Xi���Kˡ���~�o^��@�f����'g��o;�,��=clB^ȍ߽��zNj������	n*.'5���T�2c�L��mg\��O�}&�0i����=X�*w�R5i�=��7}�a��	�]�U�%���&�Ù��z�/~�l3d�u?r�9?>К����y��x<�."�|��W#�7��:M?gg�"���q{�v��-4iR�/��m{$悏�q���7h�Ve�Y��6B���+.>�9�9�a��Z��%�;�'{cc0E�E������\��K�sP���՟H��K���hz5=:]��v�ud�BN�:��rj�-����΁;ʅ*���ga��
u)Rcǒ9��`LWn��\j��:Q�੭���H�8�$ZG�����1z`������x:�N�1÷	�ƹ3gT1�}��u���IA;Eu@�םi���n�\8�k��֍:̀~���}'^��~����P�����@>�	Ć�u0�a$�^2M��g4�Ӗ`,l�Y;�w���q�,�����Z?df�9Cq)j�)�Z����E��[�����c���֥H2�K�$�5���Cﾬ�i�g�C��M$�x�:ɔ!�t��� Y0�!�4���/i0�6���}�}���HC�M z�����h4���$����'�:�5�1$0�Cl��dI4��;�漯��{�d�0�=�$0�l�2Z2m	���P�4��'S��a'��P�C�L�|�]�������I�Re���!�c��|�a���CԘH�8�zϐ�@�'S	'��8s|������C�I�9��&�
�Hi)�
@�=IP���2O�i$8���'P;�s�����|�2gP�C��b�����N$�Hq������@�!ԕ	�P=a�w�����@�$��0�<`��C�� �'i�I���$�'X$�&��`u1���N��w��|�zv��VT0n�
x�d:���C���d��0�1��Y'�Y8�M$�[�;מ��0�	��Ձ�e	�@��'Y%L��!���N�8�u���@ެ�d�^gϜ��}��&�i!�d�f5I'Y�'Rhݐ�!�>RO��!�����0��&�d�'����L���{�p��w�GM�L�j̳7->�a�{�^���}i{M���6��:N���λdȣTel����4�bcޏ��=}��q8�Ba�H�Y<C�C����c�2L�:��!�s�{��<}׺����<I�Y6��RO�'�O�d�eO�!yC�C���>}�yQ3S�f�&�-,�Qc�C�0�M�z�q�u&$�@4���I�u��Y����wN~Ͼo[כ޸L������@�0��6��	��Ԟ g�M�M��N��L���d�C�ϟ]k��Ͼ������`e'�:�}��'zϙ[��C� z��!���N0 ����|��vP�!�@�=œ��8�� `��'P��'e �&�L{&=��"!ϼ.�>����iHs�_��Hz3�:�i�4��I4����L -�u�̴8ɶC'������8�XBu�q�;�s�}�o|�N�{�ϸ!�I�@�I��:���8̰�'��L0Ra1�9������L��e��:���O��$�����q&RCl�M�aB�1��PǷ�52��
c�cҒz���0*I�!�:�P� w���q�I�M��l�g���;.�G�}'�k� ����0�e�p�Bm ���IY���X���yA�\��~��Z͊�MW��<�(BU���1�w�C�η��HC�$�O�?Y=d���C�:�u�� �OX=�!�P3�<<�0�}rw�]����0��	8̳��2��!����a��Hx�RHu���&�H):�Y� ����ϳ�1�=��}d��Ԑ�L3(N2C䁙큖|�x��,6����S�!����y��^��s�s��d�$Y<��!��:��L�'�����Nr�a��I�>a�N���^���{���L�C��a�I�t����I+&�C���I>M�Hm���m�H�H|�r���������|߲P�,��<O�!��Ru��M�|���,�����g&Ҧ,��q�w��q�>��$>@�vM!�&uBm'�q�Hj���'�Hd�O9@:���,q��g�}7��߻���ŀ,��&P�@��!�fP�I��0��>@�	�����lRx��.��\{�w_{�C��`|�m� |�a�	6��&RP�ힲN0�q�3��2ɓ|ޜ}�c<߽����C(u�`OP�!�@�+x�6`,{d:��3��'d�����������y���>.�����W�zm�4���
-���;�/`�z'[�Tͦ1Jt�[�R�p�6�B�Y�����E�z����˄DG2g�2N�ؤ��'�x�I�J�r��@�!��u��<}�;�����Ha��IĞ���I�	�=d���!�I�6�O�I�w�"&^�w�dekQ�T��:_1'+Kz�>��v�bfX�(���ڱk�������ǭ�w7�zLN��D��/V�@�}�U�0���vv�\z�	�T,W�tfL�/��R~�b�}Ey�R���"���uZ^3�\��Z;]̩�����g��O�qUe�x=0z���G_`P���	��0@���
�T�%_+��
%/yS���S~{����OV���Ved���\��1W��9K�V8���=�i"���������I��p�-Zz���W�m�/�������}�Z}ǣ��oV��D�>{�Z��������bD�;6{4���_唹;�Gú�^��1�E�E2�v����9�M��3;Q��	��q�-�c@g����{C�k���{U��9=�JSfg�⍾�h:#8W�R���0_��/9�wje���6+�2��o/_d�]�j��'�s�n[#��u�w�櫱Z���)��n�x>�H��'�檗��u�;��,����E?t�`�(�sv?J�m���2=*V9ڦD����������g��ϩ1ಭ�渱��uun+Ky��b�p"�h�ty-+��8�^��FL^��Z�6���{��:좯��H�(��;v�=0�+�|�j߾�$:���پ\��j/�4�o�7(��hz4�v����9k�-mѓ�']��#i�:�Z��kQ�@xLt�5zbd�m���U��C��:A�a{��ԭ�`d��6�6�Է��^BoL/zT�_F�t�7��b�/���o\�c0e������{8C���0�
�C�-�x`�q�pZ -J8/�U_U|s6F�&wf���}_�u��>3�J�ˍ�C9kj1�u���!�C���u�7q��A�7�r�v&���Y=���y�y<��K:��g���Jf�
^�Z1!��c����d
���l��b��P{�ֹ�㈝�;1��F��2�5�*OQ�ޥG�r��<O��:�h�e墈%h+���,yhڨ���Z%|y�YѽpF�s���mOտD������$���>���R��T҂ң��k7���Z/3vSv�؈�}WHE�V�Gxu���v�ht8���Џ�fb�d��.�-ދ��r�q,�%�&8�r�E)Њ2��VV�ٻ:�A����Uj]�}���ܥot|c�)WG���肰/_1כ]��I#Qt��X�)6�s1�f �JD��/%+�yϫqr\m�:d�֏L���C�8o����*:i�,#�.�P#@ߦΌWi���N�+n���6]�"����ʺ��(�vJx^�I;P!�E�h�[S���ƀ��g<=6�}�t�fb���X�ZU;���-���b��*�!�n30,f�X�t2d�tg�t9�+��c���>�T*f�zs�ko�����w��S�)bEˇ$vɽ����V��$'����V{���R����H^�dW] *u\ި�U\x�=i|�k��Y�G���j�f�,�bn����m��K[ ,���R^R�7�׻X2�q����D��k�ۛ�3�ܳQ*��#��2�/j�mԟk�:��b�Cjm�2^����]�l9�?���͵Z#�ov�&徛�����s.��ͮw�j��\IKmP�t|��Y,��\��:)#�5�Ƭd�}��۱c��i6�O��nV���#�!t��*��t �I;R�K��g�P�wf˖�Ű���W���I�2
M4a.�AfH�,U�,�d�(,U�X֕"����R5*+ T�+��(T�m�ѰYX*��$+&c	PDűb��P���\
,�j��Vb��BTY+U�AUdRa�I��J�2)
���V-(�a!YZ""� �m
b����DEX�Řa��:f��j��1��o|X{�p{�R��H蒯��w�{��X'W����W0@��L�
>����w���O>�a�J��������B���Ev�c����qaK׋69c��%�f^�z:��%���Qשx���k}&�\y�o��k��S	V�8|���m\Ybb�{���q��m֗�`��[��w-�n˂D%�8Q��#��^-N����p�a��؞ ��������
�s4�xy�Ҍ�4�a��CF��wh`��`ÛȲ���TD��A1;�j��0�tx^9I�l@ݵ��3�.W��C=(���|��^�{�芫��X��>ο}[�a�}ǋ�����oSTc���M��ky���7���G:�����t'�)�;�V�]��2GEPL������;�������^{f�`�#V�,B�Qy�w�@ؿ8�5�S>�b6�i�Ǌ{r/vߖr�d��ܥ�����9R��չѷ�i)�u����f�L�q�z�<y���b���@���j��;4�΋���|T���APw^R��F�p�J���>wp��aD���fP����vj����|�TZMCo�H̜�0�Y���_}U�`��8O����G\�g����g���^s�w�0ȝi�6�8ڷ��b��۱00�@W�����]D���QTN��o9K)WK�o�"�ze�қO���kSX�[E����{3�b�k �9{�: &=����P[�U��Γ��]N[{�EV�!VQ��W\���t��-���P� �6��M8��u=[Z\aldᨡp�?$R�����cKQn�*�=�ћׄ�G-�2�0�{'tr�������^c�x"�}�JI�3���zl<�v9��W9_Ϫ���O	��,?�9=&�̯�N{�:��H�]_t^��6��b9��+u���M��8��Ҕ�X�]��SC`p�<ޥ����H�[g�o��{ז��k`�w<^�F�u,=��9��i(U�2X�IKkq�.�O��F�؃�-_6�B���7q'����<Mf`�^r���85,���R~X{=�7Qۺ34Z�o-���qϺ�/UU�W���0�mhݽ�pd)[��Z�w�/m�w���oPZ�q�M�w�!̨!�U�.���CtN;t�-�?~������fj%/����j2cg Ř���	���k3y \,��:{l���4y�M��hiĘed5�5V�����}����yQz��V-b��x��m���jD
Աv��3:�[�/ǃ C�)���dJ��]9c{M�옶��A��}��2�S�a��V=�W�E\g/@܎�	ĳ���W��ށp���pp�5�}�!�8�1�1��2+j^�̐���ML5e#nT�t~�WQwy���%���Ը g�?v�	�g0*������|wo�Z�F���t�������������]�P�Y��yUi��=cL,�{��
�B|#8
0H�;��GV@yu��"��;;�;�_s�����>��Lm���;�<��W��Dm(��K�����<,���#tk,�H�[������㚲���ء���]�N;���ǹ�j+�g�=-i$/��v�����D��v|S��@���>�u��|�oP�����+��͔�Y���ŭ����ӂaV�����w��͡�;��r�֋���:]Ӕ��v��E%oRE��������_^otl�L�3�l��5���1��Gs;�q�>1�`�9�j�پ�0������>�wvG�������ǟF��t��>~�>���7H���m9�[eny���7���Gs�$�4�z�N���R|�:�&+�f�s�l5a����jZszxEN�'w�h��g�����v;�� ��N+���H�r7�dY��w��H�[��*h��u�>��V�0�o�u%�qv�'G��VS��f��"�n��r[�������-�΍M����7�89A�+�g%�z=�'
k~W:"��
ޙ8��*���(����oj�a���9	���5����F�ӻ�<�,����y�B"�H�YxT	ܞ�y�oY�M�i�y�Q��h����m��僫S���6��,��D5Q�Y�$�i��{Nf��OP�K7`o^����c��m�;�w4��ޥ�X<TK�7������,�d��v��i<FY�	&;�ki��u���B��v�b���j���9r�쐬/�B
�M4��m �oκis��F�/��H5�[�m�s}��UU4���;�Y������>��Q�q+;����^3jy���Gv��eç<�ɉ���1�-���cn�����}s9�������#/x�w��f�=�׸A��`��7����ώ ޘ�î���5i�5��eQS�6��֙�X��!�7��f���x,ξbq�.0��;]�9��comhOx����1&������n�
�V�<Om !��Zߵ�^�)<,��V�5�I���b4��xxx�ﶻ�v��;��8��I}Aų�;%������ŦQ��u�oG�6��Ș��3�i��#ճ:���ǳU(u���cI�>k��j 2�>}�n�GJ�FT��mE�DGeGN���,h�~�5�~�s�Y�ZyS�DW���WNՃ����f�e��`�LS�@��ފ��qCl�������R��Q��s���6b:�ꡱO���G�i��Jjt��^�3��U����c�bdC"׎NŎ*�b��e
�<1����/��ӳDd6+D�Щ׎�֓<f$tm����mA	33�0�á�>�����[Xt_��B瞏�`Fx��\8h5_�>�%�r����V�}�^k�uA]�M\9N�g�cV�q�3��%*!��Hys�3�O���V�J�uE���ȍ�_ob9S{H�Km6Ҥ���I������V0o��>���hÓ��5g)�x&Ҋ�wgӮs,�\�"��O p,An2�n�wj���ZP�nm�Ҿ.&�!NGw�2P�-�3
<�%�����9+���Ai��Via�2t��o�
oB1;��s{-{,n��ɹw-$��3O:mĮ��j�EK��"�ڵz�r#n]�'/_��bv���{�V�A1�R���2�A�2��ښ�uͻb?��EJlɜ�W�p��]9��t{���TA�SY�S&��~ͬ��ײ��N����Js�X�%v%���h���zf9�L���lf+g�m�@ی�빆�fh?2�v��)�\1b];GU��:�[��v�I���9]�T�j8�7�������y2T	���y_02]���"\{*č�-ogN	�9�R�ٻ��x�Ö�����v�I��I��r`=N�uHFI�qU�v�x����a%sN�s-=�Ƅ����5�b��kX.���ϵ�� S ᇪv��ј1.��k�m�U����HۑIY�f�[�f]ܾ�'mL�<�w��q���*G�$r�p�x��Zg�Q�ǃm����r�x���m��~��P@}�
) J� �d��
8�Ap��%A�@RR��V�Ɇ0���VUH-q������j�
�-�J�,(&b�W�-b°���d+ �J¶�Z�Im-��J��Z�q� �m�
�P�a��qV�T
��Vi`eV�DC�Ţ¸q�)�Pk�-��%E��*,,�Q�P�Ɩ�
�(���2�mV�"�X��-m��*V
�K*��֕��m�  P�'�����a�ƭ�vNR���列2fjqk�r��"��W�����_�M?+5�-�!������ ��9�L�[}Rf5�VӜ�R{KuJ�]8*x���[�xS���/�>�7գ.�^�(��Un�H�7*�"�Ɛu�}���4�K�9����>��K���ßO�����2+�s�ؚo��30����C��Ft�d:�d���WH����"Y]��H^�����|�o)AX�QB�zj��B�q<��*q"��Up�2�֍[�l׆���}�4ֺ`T�D�}Vo�P�\�A��R���5��Qm�+�W7�B���I�^U7��6�gX=e�N�W��<�f�u�;]Dc�kEK��u�H�s��mb�6��Wk��=c�<�8�d��̬��%���d�p�����+��:x�?<js=�^���-Mv�O9��)!�B��4%��ަ���Eۢ>"� M���t:�k8O�`ʞT��V�Ǯ�W�3��ef>�c�h�5��S;u�`�]t��.���y�3y"iںB��8)s^��,Z�
c_���s�5�C�Ӄ�EX�N4Eg�eMȖ�2_��d���3������(��lR&� ��YO{.����HM5v���*nV^�+ 7=�@k��è*�L6M9ʗ�`xj��bi�h_-��0h�Caq��m<4}�Å2*�ىjK�_��G��-^`�����-Ѿ��v�;�̜�ZOok��.�nn����ڊ�+k1�2�Q��)������)*�����g���]��>��2���c�{�%���a�]��0G�
�j~T�xs��i���$��g*�
���J���>s��Q�b��g1�*T�=�f�K���UAj����hy�q�����)^�P���R��C�v5Hxh�4Q�`L�&���s�o���p"�\�7[U�Rl_��
Y��MΨC���8�T~#I���Dׇ�1���+�>��\4T��*�G�|<P��W����]*��G5�y�,n���]+�R�_s����|������Y&;��(Y�:r�b��?�tŊ�h�*�⥴�o,�Ѹ9f�ހ�60^�\ ��&V�uuol�H%\�T�6�Y���E��H���=�㸃���oCs��W�}=s۰t�f��`�W��p[ȅX~�v�+�E���Y��*�?c5�q��8 ?Y�K��\q��,��;ݹDxR8\4�~V8X��*�NT�t�^ɺ��~�n�x>7[r��)���<����;rƴU1�������ׂ��`�<G�4�:�τ�^�|Ί�4U��R����"����¶L��X��<*
C��3X=�_h��}��Ng�'�A��tz�4X�����4ɡ/s1��iA�M�^5^�����>'F�>�^��r�^*R,b�A���15b�I��[ �Y^����wP��^⤋�x�8���c��n��6�<z-u��X��_V1�yH��B�x
� ���d�]����{�����G�W���|�1PU���F�������͟dN�vQ�t���6�r�z���맮�BM�򎨕��d�������*���]���$��gi3�{U �ОZ>�u�
�h�j�Չ�ox9��>$��Uof�C��*�5+��ЭѭKV�7�+���V�QV�X�Ƞ��G��������������T�5��_5b2�t>f͞��\��Ҧ�)�����=���*��8�/��\M�u�>��׾8�#��	5^��F���,"s�`�N���8��*W�Rӡ��[��d�L��e�I�l���(eM�[3���誵�8 u,/GN#�h��!a��t�t�gE����Fy9�ﾯ��i�@�=��!�
�HO���g*OUR�5�ױ���s� B��Bɪu��������w٬��Ovبs+.a�Ŋ��ʐ��i���<��C�w7��Mg��|)
�Wf��W��/*���ps��@c��&�FS�t��Q��*n;��A�`Ы��=�w'a���N���(t�*�=�{ML�mz�vֶ���q{_s5:��tW	5W���f���	�O@1�{�4רp��o5M�
�$��R`˕1�Řw5w�T�H=0�l�D��01�O��pװ�>>��K�y�ج��<<(i�PU���ƫ<pK(O=�ե\�u��X�}Q>|z�T]̮է�c������wђ�ׅ��:��w��&�Rn.��rގ��r���>��}�|���o�=�T�½���LF�L:�>5c������F�����ø��¹���;�s���4Q�O�T�-*_NU�p`�9��,�s�a�a�P����1[C����xx�-��
w{%n���� �_j�� b���sB��6U��;J隊|:nj}�Fa�FHuT�ܙdgq=s��x":jrK�s|/���LYXoJ'Y���3�#��G]Q�V>��]�4+�L��7EN� <�^1�q#�tV����m�h�}W�4�aV�)�,س�N`'^���@��:���mq��T2*wap��a�f�T�"νcOI��ƙ��8��eZ+4���ﾪ5��R"�f��?����>'����C�(���Q �>���s�o��*��)���ç)�uW��h[7��;L�pb��P��_!�iLd�Z�7��%��(���*�Ճ�v*�eTfA0��xF��I���\��M6!
P�
�k��pxk��D,5nbd��t�҉�9;#���b��&flh�Ƭ
�j�t�{ْ��`�LV�f��*����i����&m�?q~ӣB�Ռ�4<h��0T���޼nF���B����w�F^X�t}���b8�;@�:9��}Jzt��J�2zcdp��s|���� "�E�}��Q��a��B�Zd�����+��"��R*��R�1Eyy�LoD!�$Bl���;Ѽ�����T�*Y�~b���{�h�x���R�n�e������þ�=yZ�����U0"��}��λ�B�Ph��7u�j�P�]�w��AGM�;����Z+Dv/��HV��~U��z�+��V���کf���X���B���;�[@Z�Nƪ�D����5ҧǔ٦2f�9l��gl�3ơ����R�E���g0�P�}ཱུ������1�GI�5P
��3���J����J]jç�G�J�����[�G}��A��b��R�^�`���nW��0W�|A�^�Fυٯ��x��}CĀ��+$�*B��e�(�:V�2�r�A�\�Ԣe�W(���0��)�@�	��u���*������]����оd*�1�1�`d��0!`rn�^o{��:��5^��/�5�4�ة,P��m�=�c�@rvnvS#کN=/Ms���Ha3��{׿W�r�,R��fe
�>�:��WPy[���~Ⓙ]0x�j4FP�®��_j�����F��"��C^�麻�^�ļ�;�T*���h��Y��E�˺�;#j9%�����\�!Ձ����c�̔��5o����3X)U�"�D�x��f��ٸ[^&T��ʕ#£�0�O*�@�Ƽ>;n_�Y7B�5�~C�xQ� {ML��r��$n�'��,�!�Ő̼�ɞx�[�x��/Ɩ�Z���ҷ������p���g���!Y7v�F�u �靈���٭�o`F�e���j r���EWn!n�c�N���Ff9�w��j�h��d��ڋvv�"-٦�ŗ,�6�wƴ�X*J�U�Ѻ�AwvMJ�,?M�᫚�zҥ)wa��U ������O��Dw>��=�f����ÒLY�ɮ��fԙ�庸k#݋ra��+�?�c�ŝz>�v���R�tT�du3]Xu�3��]b�)T6.�La*9f�9o&dI������48�Lwf*:��.])@�����3��R�T��.�y�Q|��྾�
K8Iʄ2+�Yh�i�4�E<�Qeqݔh��?:4�߆��Of�:V���Ã{���Sg5*��(pw�]Xr��I(z%v�o*�ޑ:͗�Y«h��"`��Z��}��+�Q�O9�w+�fr1#s��һ:�*��_C{�˘��В��נC�1N�ɒ�n��[\�t�h���<Y����]��|Vp}w�GPo`2�S%2#��M+0Hv�,U�;�8��������Z%m-4�Kn��EE1���-��K�09��>\E\�fK����ݦ��u�IR�1uHy�r9"h�f��\���wwV�s��Do%l��7�x�Nf��CM����s/��<����8P�����+B�I�����H�1��Ŵ�*�
�B�[iUm�`�KR��V[QZ�����������,[J��D�kAbVW�3j��X�+(�dE֖Ш�EQ�E�ԣm��DAX"֨ʕR1�%J�J�V��U�1EDEU
���m���PF#`�k�J-�+b�DJ��Dk
�����"����QX0jX¡KJ��+Uū"���,X�,8�X�T�T*0cb��Q�
�b��QbԕV҈��Z�

�5(�
��B�AJ��%b1hT��F�X(6�(�Z*TDJ�X�0R����)mU��j(��*���@����$F��b�[TUH�UR�h�R1U�j�����
�1F,T�lQ���h�kIi,�Q#H�Tm*EZ �Q"(���g�=�珘�p��q���,��LA�ێ(����%��n;���՘�7�g[���)���8B�-FYVS8sOj����;9.a�7I�
W���ƍCX=j򁶺���lV���*Ch��gµ+��oۋ�w4�S�]!ґ
�k��ك>S0]�/z���KW=;"K��53~V=�S�ϸ�v�mכ��x�%e��U�y���u�i�*����P����n�V+�ı\�xh�(}0�J���pX�9,sCVƻ*`�9��4��yQ�"�MTs�������+�>��"���� ;њ��L�R��~��W�E���Z"�P�2���J�?�K�Ŀ,�W���˭��J:�\��w�-��rs��˭�Ӥ�WYN8Gv�.,,��륉k��L �y&Ա=�gt<�s�l��r��DBom���:VW�X�驂���AL*��Xs���lP���=�b��w���V�{_�2������=Z,�h���x�4G����~�׻�� ��*�Ң�1�+�K��;�R?�Юt��
v��U��Vo��z�}�Z��G�9�)�����YZ@�*�����xc&���\�����c�h���^*���x�*�IAy������pxP5^T�O� �\>��6'g����°�Nu1�4��H��
�5�k��\7��3�Om�ׅ��X>>�b5�4� ����gҏ���F�M_�Z-9���@��B���r�I5��o��t�qyL�)8�5��p���V�k���}�g>���4W�-`�?!�<3�Vma�t��&�����Jlҗ"}&�f'�v�������\n��[b�f��!�����ϵ�Y��=Ql��Z�hFeXꆼ��4:�U#4���i?Q�+f�_z]EZ�i��+>�L.�Z�*��4���%�{�'"?X��p�:�C�o����c:9�^�@Q�>c�&
�LWa_P/����H�VS��:6�\B�zl�wN�����en��xq�{�%�u�Wp�
�`��Z�x���ɩ��ǌgY�]O�;12��S��%�ř�r����Ho�y��}�)2�
v�pV�|��������P��z���g�S�AS���ȵ<Qnm�F-�Jt+\eJM�'~����y��t��:��s?&�:M�k�C��|�}v�����gB�T�y��԰�۽�[�+t��M,��Y�83�T�U��jC��*USʯ�-�Mw=������@AX�k��xk,zm.�������tL"��S1�s�*��n�e
L�7�e��~��I	�QJ�Q�:�\���ى���i�j{�#�s�>��u����+ִ=5���[]~�fvgw�TT��BY*�p/��
�dê��KI7&}r������G(!Z(�4�j����vp|�m�u�����fŋW���fY���W�Ͼ��J�YWG<�_�\5��D�+B�c;[�^/b���e�݆76�9K���Ӯ���	�J��5��_`�?�վ4�OU*��6*
��T����1�\m����T}7>��b���f�U�b���Ż�oo�YU�5�~T<8xU�#Z��p{ʐ�]��ֶ�|�\LWT^qu�%��5>3� ���ܻ�dΰ6����U�ex�)�N�F��2�p�T�AaWo�+/�D� z���B���F�˩�q�4Ɗ�c�<+Q�חC2������p�T�8P��p���*I���w�H�( ������Vuw?��шߺ�cY�y�!���T�m�ܭT�񩇇>Ph~5+f>��[�`/r���볢�ݝ���L:���;����l�8X�쨳S��[���m�\�)	��g\�ʫ\ҌO��U��3�X(ߥLE��p��f�l�קV�j��AZ t+�V��x:��� �U��R���e��tw
�5*��n(
��\���ؾ8�&_f��6�M�t�xQ�jpWF���Ջ�o�R�(݁7�J�Q��ю�2򌳃կ.#�<+d�=0'�z�q�Ei�K�X ��sX�+��f�-X�9+z�ݏ��5aUxן��<1��~0��R�z�__�",Qp|Ez��?���a5�<9�����G�ss�]q
�R�u/�`Vr������ޤ�ͷ�Z�����h�:q�� S������X2�8�R�q-(������O�Na пQ���r��,��r�tx-�۔�{tS��M�ӨQ�v�$w^����=��N�?U�'�����]jݩB^1S+��p}�X�U�mX}��n��2��b��@�K� X������ݕ�z��m���١70d����R�0�+��@�5|�R���E�tl �+V�o��Mp�4�� ��ރ�鹸Ŋ�lA\)�j�����+�o��l��n���]C�B#93ҤJ������-xVv���^��4V��ч<k��V5��񲂠G���5�=��K��ȫ�Z��8kW/5R��z~�V4�ω�������Er�}�0xVY�;k5�=+�7�Kvwy�UQ�c�d��g��ٹkC�C=�[�6�l�mE�I~+E�N��پ�f-�[s������M�Ya��F��0�� (���N�^٣�|K*If��cr-��8��ڥ�t�&�X� W�+p�P!rN��&$e��g!�)�m	s<թ��έ��d�Xه��ȋĚ�i�E�]*�3D}�5uY�嘀B
�}�H�&�"'�uw��.�A. ��r����rz�oֽ����0:g�5���eX�
��t��^Z����\���Tg���M<�}����ӯ�@Ʀ�����~T���Z5!��,��i���H��~ }�x�a�C�C^U�ӝ�s�2���f2�"mp��Q0d*�1�=��.�NwO�8&ł
�� �U^�V�CY� ��i��N��7�*FGע3��O���Ýk���((kf�łwb���Mvգ�0k��%�Ż��Z��(�Y��p;�.&b>�{{9�}9&Q�a�Z����}��y�kTC'�߳��)�"�R�f��U����Iǝt��d|�V��� �Q�}�����)nl�i�n*���ܰX"�@�^�-�T|wi�iW�Y�l�^Tm�ʅ�G��:��F�n'f�'e�!}�E���.�ʭo)�<�����n�3M�R���c�q'��ͣت�R��@�\|)5��J��#��Y�i�o"b��+�a w*g���i�MW&�-��\ mq�]o��8�^�R��F-�2ց���^� т���V3�W���>�s�Z ڔ���*o�t�N�/���S��;UE���ܕ'�ě6.���7!���~�l��Xm�nTђOE�_�@{���0���Ꞡ��=1���xT���QN�a�{n-p�\�w-Ta��(!�q<GUOeɫ�x�^k�f�ܾ�Z� ��S7ܥ��,�T�S�p�_�0���R�n�Nn�ײ��
$S��Vm�QB�dC�"'�hF�#8B�L�� �eܱ���&�E�>�:-��um%�t��E�����^������^Ջ__��j��=�S����TS*���[�Gڴ0E�¾�^kױ���]Hz��/������W��Dlg�����s���ˡ�v�g���0)*��TE;lWK���^����|L1_)���|o��T�Q�*{�,�^�7�����H3%�k��r�%��B��)��np��L<w��GlZ��R�]�>�֋��j�E��2R���:VP�뜘!��n:靡*�Q�{6��h�5�sY����-o�a����
�xou�V2XW0��k��(a���@Ѻ�`TM)����\��X��L�ho-�2�%l,��p���b�O������#n�a�.�&q��pަ��2�&��n[]cˏ}�����d�)�5%j���CM���`,�ʋ�k�n1D1�ۓu;�)��3R�2�Gzu�ʀL�8��l�Ӯټx$f^����t�K4rc�-�q��AL��L�qM���4�n���U�Na�HQ�L>�|2����*;�^b(�h��Ё��ή-ӯt��]��ն3 ƹ"Lj}n��8:�jpSo�q���k�d����e;=<ޜ�����e�1f����L�7/�W,%J�����\����ފB�Pa���{%u�1>Z�}HtṜ�_�;9���_=��gc�_:/�,�V�lf�zKI�7\�r�[:�G���^s���Wʌrec0tן���G��_b9�׸���6���GL��>�F�SÈ�v�q&�M�䉢M�4W��1�*��㨭�$�׃�C$����fL�`�c��$����QH�.�l$�n�r��H��i���"�eEE�֏[b�F
E��bDQ���Db �b����X����1�QcR��QAH�+iD@D`���D�b�j���IR�(,ZZAb�jVT*�$m+��ň�E�h���ʢ�XK�"�mBڢ��*[h�����Ŷ��E��������ؕ��l�QV[DQ�Z�Z�*�X��e�n1(��*� �EDE&P���ض�j�_������O|�|ݯך��+���|p;������$t�rK�����2~�u]+��R͚��_3��>p������p��!�F��,|�i��F�ax��e^�p7��M�^�k�*�T���%����{���14���^���v�)eU��J��Q�Ֆ#~ɒ��c��aI��uB�G*�4������ɋ��~>+ōZ��^ +��N�*cJon��3�^�`ɚ�0l��� W�%�����5fӶ��P|@Ϯ�b���3^ƚ��6�Go>�h��u��׍�#LT��>�ǀ,^�r�6��SƼ*q����AЪUf���[��	j_+�[j.�1\��.��4���9f0ǵ=��/�k�J�9�-F�؈���T�9OZ�=�ކ^̅sm������%uF:!P��},��v�;����D�߅*x���b�����C̺�Dh���L��!����V�����3���Hz�0����,�^�G�}(z����{+ P�x&tJ (�w��զ���*Q*^8�	0R�DV�D�����{�e�N�t�ѡ׊o�p���\i�����3�^�80
���)V���f��f *����^���U�g������SJaʕ�GJ�=�*:
1b�%�s9���F�xhl�����|eU���I���>�~aЃ�!��4�g��k�|&����x�}�*���F����J�/|��A_�Ұd�� ̠�?�ri�e�s�;��G:�+��jS��Yz���33��2���P7[�Q�gh���B�zN-c�Rea�h�@5����EZ�7{%�����r��kP��U�q�t֊�B��X����j�����p��� ᪕���𬷢�#D��Q�u~A���w�o�g�~!�b��������٤�oҘ�����yR)	dH��8/z>�'Oe�ۥ����
���Κ��P�E�]i��������Qע yT4����7'�^�'l�u�:��h�]ӟ$j��j��_=T��T�a�V*ǅ$�F�4��: tqhuj,|N��Gc4����{�O>�*�-��2PӉh����V4JpT��첝d�����/�Wg��T���n�|S��k3]Y�Q����}�UUa%)gG�
��P�2�O�T�Q��K+^�K�{�T����P�Y2���Z>U���.�-���R��!2z/+�؍`�P�g����u��5ՠx�W�?1�n��cº *;~���x n��ܷu�-��d����\��\��}����P׼tk�/����CO
vh���>���X��< !7O���Vk}��V��r�<^��J+��o�E�݈��~5��[��i��Y:��־a�5�*6D*r=>�[U��'�c!����Q�B�X�}�B����[C�ܫ=�(�A^���U���.}���&���ֽm�Z�䢙�l�V��+���,��J�eʗ$J�s7=�UUW�kܾ�c��|��|?�^�f�p��@�!�tѮ�2�1�bfwk���w U�Vu����h�)��|+O��ks2$�
������_GU�#c<�ВT9�o=���4UڭhP�]�CU��#l׃��Cn,9���������]KwIl�z���9#�O{��R�+/wL}`X��4�ax��n��g�%Ȼs�P�L��:���#���E��%��'��z�w�o�;�ٵ~�4jf���F��Dl�3�)��"����E)�棕yuH�����saϞ���,��Oj�*�xTT�-���8_&-W��5�V V��IQ�r�(�.�`��w�_H��t��fQ��(��Ih2���������Vx��udÜJ@͚.��A��b:I���l���*�L�*�&�3vD>DW���e�5�;��W[7��f�˺��;�\^���tʖ��'*��F^,!�c6([:q'5p�T|ՊZh��i���ƫ_@D�hee/�7�lX�f�7����
����5��ֻc"\����Q�2F^	�&O�+W�u���g�NkWr�]H)Z��nͻ7� ][�P;DK��fp���������i����h���+«p��V��(�!N����Wj��2����o�wB��|����b�,C�1$^F5�/q�u��-߽�\_?����Ӄho�xܙ�X��9�J�/��C�!H�Z�諭��{͋�dz����wN
|T
�.D�gܫ��'na�<� �
|b\ƺR���`z�μ��uz��M9g�]yN7��Y�}׹��񧌻C=۝y��Iq5RˡLT�1��Uۺ�]4�0Ϣ�J��n�ܺ�y.q�����W�Ѧ
_��f/�m_�/��&?P��to�!��no[lv�����B����´V��H�����֫�^�,�2��W�b�Ɛ��w2�t��k��P�&��7떸+�����C��s�o		e9]9}��^�_xQȺ��h�����9uco^���9���C���b���f��7R�N^��U���C�����̗��=*؋�f�K��k�B�44�����ѓ��]>��2�X�&&�1��ݧA���Y�ňUV
��x+U�ԅ��_{���b�us�@F�-�s�G0 zQ���o�˿M�k�lב����`p�"��Mc��j4R�s�[����� ��2�zEr��6��	�R<*;����䚇�)���VQ�Kʗ�|�g�C�BmSMkM�;>�� z�;>����(�9�=�Dmyt���ؕ+#���a�HA��B��P�=�wq��I6)���xR��4��_h��l}B���|X�º5��Y�A�¼:�(uj�Z���k2�NΧf�j�YUw�<H���&�T�N#e����ՙ��YN�bNˌZ���ы��	5�IʲI��NeI�y:�V~,��p?����9ח��L�^َg �6�4���Ί��X6`X�n�:�=�xM���@�Ս�3���EO��A��d�(Յ�ªae��N�o��f���Tp�PTp�iд�DX�5���ɇ�t�f�¥1ƣg�7�����e���*ǀO�U�*�
�Jγ���G����L���3^&��\xs�F���U��le"��}�fR'y@��ؘ�Qp����u�|��ۃ�D�/f!�Q�\lp�t*�5�x�>Z,�
��[-�o9��-;��!��Z*ŀ,|�a�T�����Bm��@�F=�Ryn���ۋ�wI���c��ֿh�3����ީFJ�˙ ���\��G���ḣZ���Α�;X��+l]ר�=f���87&S���u�G��ξz�����4����p�F*�j��Vw1���H��	�Qs�e�E)P���͋�-q�ߵǸ��:h�4η��i�s�]�5�w�����%^���Sӷ^n��ԛ��W&b�pr��TNTmGKURf6tW�ߝ�b�-Y��g�|f�� ᢭=�T�3LT������	[�=��j��b�]tջ?x��Ռ�zÖ_�:�h�]��5b�T�Y�������8w۲��+�s�I�S���w���Lj;�z5&%/Nu���I]�IV���ym��>��EF3! ����#Cf^�cy���DL�&�l��X啬*��h��e;���V�L��X�V�lWt�>u�֧n(��c�mf󆴙͂�	Z�5f7t�#Z�آf*$,��C�!���o/���M�ܤ��l�*%Te�8�3#�m�ᔚ�����6��T�/+���}�XgY故��;��m��p�I#�8E���b��%A���jŞG;t"����e�]�w}����)�Z'�F����b>��N]4��V���)Z��Щ�-ݴ��f��w���������I��&�<w
��o[H�O<SI�&'O�:�[��^ȗp�x�ϵe�lX9�@�:������s��)�u�����G��<,W��ڮWO��quk� �S�Jq�9&ڕ��Mk�:�$�S���n��s�������ϣ��{-�c�*�Oy�ԫ�q����j�{{:��<]9v0�$��8n��Ǎ3�et�B����*q���(����Mf��X�W�n�'o�}���̀�P�SM
�qYBM*�Lɼ�t�j׌.yc	d� ٹ��G�g�1���;h�)���`�#=g]����e�ڍ7$�'��q�{M�"9}�>5�}��r7g_wwnws$� ٦���ЦH�d4�N����ٴL��a6n�!��4�xɌr�BiU+ETW�SQ��V�-,DX�AdVa�V�)�J��T-e�FҶ���J�"�Ek;�CU���,R6��H�Z�`,�,��f�a���R*��"$U&R�D`"�"�E�Qb�,R<n񽝺���z[�ړ��gB�E���W(r�*$�����AH~}�R�}b�Mӌ�0xR�*�Z͛�R��!�ܾ�p�8>@�W�@�o��'�zE�~!���w[��5���)W�qފN��̣gh����[�4h�(`��.��AzG^m�@^���UāN���]�f*|��`����Q;ɖ-�����ǫ¢f���&�Õ+H�NQvDzo	K˲�*�����:t&~8h{�E@Eu��ݞɚ�A�)VG *���b���KꉕUZ�Mo�5t9��g�L%�V����e����>2�y7�v�9f��|�\r�㩺�&V�Ow��(��e���oVW�қ�*��z��2D&�B�ݩ�4�bݫ$y��g�5\�L78�%3�X����#��E	}t�h�pQ�WI��!��Lt�N�6�U��4.�EИ9Fw*��TC�ճ:Q�g�{	.�A"�Ѩ���#eK��e���������왂>w�5 Q&#�}1S�S� �k�pV���r���[0!p�����¿`�j�â����K��iL�-5W��{�
�}m�l�ϭvԕT��ɨ�C^5�Lv�7}�[��C����X �]>k����x��Lݭ���X�Vf���Mo,�k��okp]�b���Ǎ�8�`)���Df���-���a�AqL��S���S��Z��^�J����ch+-�J�d,�����f�8[��v�OyQ�v�b�k��gg"�q���>z�����9���rk�s-�6��t{�6�Ps�;g:�?0ŭ3x�E��,m�����&�sj�b�lT1�
����>���
V�q�1��"&6�d������׌x�	u��#66�耣��%�ml�n��5K(�O�3`;y^�CU���u>�O�5=w�M��`�q���>ͯ[��+`n���.ڼ���� ���T6;n@��w2m����6�-��3�fċyTV�+�˜�Y����I��� ��K��/:�Ϩ ��~s}����D��GܵOO�~c������xq-�N���s/����P���F���]�r���}<o���^�<�Kt�˽��s���f�u�q�c�}:p�xj U����o�����f�:/q=(��|�=���Yܣs|-3y72��d'�j�����5��GF��=!���������V��]f'ܫe��m��B�v�Ъ"Ȯw]��˽4��[��v�v���zfVJ5%���s�6r�&)/�fo`�jk~pR�u���=km��R�����t�h��;;j���<��F�4�u8����	����qf����:7'eOh(u�b���@�1մք^��!�k�L��Ѭ$Mg+�Dcs3P�t�˃������շǊa�@�!^q����`��y��Ń1��e>�W����R	��ᚌ�w�'VQy��0Bu7�oѣ��Y碩�w���K�i^l�Wְ�wl�u�B�(T�|�@�8�"�
�]����buղ�,�o-�v��͵`[��u��C	eH��l"�Rjlf��w�b�C29��o��&��ڬ(�Y�v	�W1��(���	#x����s���!:�fb.9~��q��6�mf̨Y�q����e�k�̑�I�~�C�����P�ʀ���m��ZB�݇�5�m;כșw4o`g(m�V�>�͉�q9�q9�bj��y�p:�1���L�qя�u ��h���o ��b��TBJ��*sv��Z_�%	�p8��yE-��I�����K�zC6���z�N�rU�[F���m�-���:m���w)Y�v�u��sP1ul��+�I��z�GH��4[^aq�35cIn���vC�����|�ØyJ��r6Yoӕ`���nV^���'%���豏vIɲ�en���1����̘�γ�ү]�X.7le���zl-�&�a2�3|v�T�E,[�w��s��cp����l�LQ㳀 �6{!��|R�2�>>�j^��)�����8�a��c�}�K=^:}R�#冽�gm�ᝎ��a�nV˴!iEr�`��ݧ���rӕ�I���� f�i�����VY�w�61gkH�f�a���C����x7�S���p51ü�a���C�%��;�-S���^�w�O��� �#�e�MoG~o�\�H������l����k����.�;�y{WxA\�W�ϚLx�ȁ�>��iy��t�_�L��l
�$�1�^���2���=��bh���{)O I��ݐy�4M�� ���K~�~��]��j�׼
4�kb��	|�(Ж,�sD�A^N�Wtn��£�*�+�73jLR���<Jt���
�h�U�ݾ�S4-ã�y5U���n5LȘq�¹�� zduC�<=�(C{�=�Qo��g��eqS[1����׌wom����1Q�Dh�A��qVl��ʁ9;܍���{%zri�_m,�TZ1�3����M�/����#��g;V��i�4�;<�.,
�sv2+��`��љ�&z����pފ^V��@�#���|�Έ��>�һWZ7�z��I����.ܑ2��IE{�GIr�F�I{Ϥ�-M�8�</��-����+����{D��6�g+V=4\V�����#���5�ݻ�u���8ler��7v����]�3JQvv%���9���O�4Y�C�����i,�|�E�򏼃-
强��X���Q��
5�슞���F�4�\"�����0{x&+���S
��glg`[�|>��͍9E��VaV�z�6��z$C�'f�Sݯ�w��7g�֬`m��ڴi_����F��+����*�[�;/=�Rf�1�\�Z�iO ��j,��(t��V�K{1h]S�t���m�2l6�����n�ya��VLT%�P)��.QKBw��[Ӯ��J{8�u�����
	(+XT�d1&ui������5�p���4�S�kKW��y�j��q@�n�wBVWSuVkR����pvn�	�`��9��oo)5�9����wղs�@��_۱�����w]�-�t�u��u��Noge�y,�|�V9���Wf5K��w�-Ť��)��=xN��i�N�+rh��ʙ�g��eJo�N]�I��fU��L*�ۊ��,`��������8쿥��á�a�Z,��[�K�h�@�q�{+
�z�� ��*����urE�돪�#���ѭ<���4a���>*���2��G�;��ͬn�0	YEj)9�%iWu���k��?9�>΅qظt�۴�ܹ��m�3M�D	$"K�1� �.��K��(���7����.qc}� ��yC`�"Q���[���Oz]edŖ�z�ò������N����ʭV��WJ/1��������f`6��$
��	ܓ��o�5����ͬ�CmT�'Mp���㵰��wv���R��6���H�6[6w8�]r7L���t�1����Y�BԾ��K��h����9.��Ӣ��F��a��4�d&2zo��5���T���db!*[E4�aqp�C,�R��H�eb�R!Y!R��%�$�*HZ6������
��!�k����;u.fC�/2d��i�3��ќ�Ө����յ.��~:}/^SE��+�w8�$�'=�����
���p9���������\_\�Y���j����JTm�q��`�o	�<�5����G��\�}��{���I�����[h���ُr��я�N��ǥ����P�����'�mA��sw�Ĺm7+���w�z�;Y�;��_;�n�������f�<�������{J�K�U��P�g����9�6r[Wv��m[�|�#{X����l5ȵզz-i8�K���ԗ��5S�]�+O�2�vI{��6-�pB�i�o�&bL��d�л�sB(�l{�)�=P'�fR+в<w��{n:�>�`v$F�M����˞�'��ZѦ�M^=�Z�F�׷o!�P�����6▬�q����zMgo>/i�9�k<f��q^�y��׼�gr�h�����S�b��NA��n4��c]O� *��=�uJ��1n�-&�Ef�6j���̨��;u8JU��x�C����oZ����j��e�ĩ��rF�f��֔YڽAI:�4��~9������VF(��F/|�&Yڳn�X�$�CC��ۿ\���"xxV�/��[�w^?J�ͧ��d"���W;h��69�}̮.,V��q�8��=�ymS�q8M;{���ݓ�y�Mp��D�/��!u��T��r�f,��$�q�x��U�27�k�j�CvٴՊ���O��/�.<��Q���W{H���.Ehlv�F����8��
�sd��B=6j6�IS^�wy��Hӣ�}�/�є��U���F�g�g>�џz�e��Y�ً%hv5���{��O��5�W�;��ף�p�h��:>�-B(�G�sUm��ft��H�;F����!��M������}�m	���s���{��{o���Dgy��o���	gqov>���r�ϫ��c�����ڣ[�љ;xY���\�����F%��ޗ;q&������b�PęW�U�����E�7{���|/�;x��y��a�~�*5�V��̈M�(p<�;�9B#h���oD�g�C��j�u9��Y{C���om�HkŤm�0��O2E���^���7\�M������07��)%��c]��}��],�v(��s��>/�S)���FD�%�2{�a�f��ȾX�{��N�
���K��{���Ԛ�kG���C���fn&�z*��<J,��3r�$xG�}��y�
�Λ������B=�u�W���:�+0�1��f�g���ٶ�$�-��Ķ�u+:�&�ī�Gq�y�-�)��S[#��&����Ƀ�H��Q�CU��.�Z��)���%���Y�<�4����n;��i��7F'&n���c���ۓ�y����B��^��ٚ�6�F:$��jbOk'7w�b�Y��Zg�\�X�w������賛T�VaF�%"��(ߐp(�^�Xi��G�=9��8�x+���U�x2�\AM�X��!��=�o}���!�nj0+���	[|��5�ߏ�*q�{v����L�@M�#��v��錮�t:�,�c>�e�1�5��=�e$�2�u�ȫ3����Y=��@͝>�z�5W��r���gX�A�rW+f�ɧ�:|�.�i��ƣy�J��Hsv��K�I��A��[�iI�v�o4�k��gH��2g�-���O4�eZ�A�u������l^�q��$�;���FD�|2���xv��ʋ��鮚n�ɪ}ę^��}q��[�'|k������t\V�T���+���>�+<�1N*��ޱ[����tf�wD�R-�ؐu]0ح�� m0:anEO���s9:�6�>5�#��=��d+\��5��OJ4�S��iU�.�TFo�.	�)g���Ld���Wh!x�`�ʴ������mu��'r��=ó|�r���
�䳻��
6q8Fv'�ѹ�y=X��P͝���u�A�n����v�n=x5�Z�oHױV �� ;���0�([W֓�!Ӣ�f�뮲W����1��V�7w]�a²�����E�5�<GK�ߘPZ0]����2�\��arX�d=�^3B��zd�����4|��Q�6LR4�M�s�Q�i,�1�yV�"�r�>�DgF+�h^���zr.���%Cn�EK�yz�f=��;��,rp�4����~f����»��\�W��\�p�[:rk;gV*U�z)�Kb��5�ww�ez;0F�ٸ�Lt�Y�gr��..�-�3�rUM6E���i�{ ��҂#kbk���~/�@i譺�`��u��:[�G�V^��0I��\��W��:�r	��`�y��x�ǎX�!d�7��;���5C��e��J=�VJ���`�#�/��0GX}L��>ao�U3��p�OT��������5s�,����u4+c�����ϻ�>�e�����{�����xCF�������F�nA�e���D��t�s��$qP�s��6w�o���B㗥<�eQ6���������\:1�y��!5���*:|�y�,=}�j�7��p�Vs�7��[�/���ގ:�V7L[;�s�"ߌ5��ʑ�B�Msi���f��k.�&�%1����m
�}��;b�6r����;��Q��e�ݙ�5��|r܆��|&2�\��z�Z��k�Ҟ�thU���؅�P��Ȩ�':��C���@��2`�ɛ�˾U�j�ΛD��p%(輈c+^��9�������@7x�E�8���M,ܫ�#��*w�7�r�w�6�	|z�b�����Bk�Z�{�y�#�(d�E�:�؃��Ω�:�)��t�wa���+1\��ژh`bd֍rFv-5}(.t��	H������j������ '`��"�W�u|�H���,z�I6�|?n���_
2������,��H�X�*��;	/9�)��u9K3y�X�ki_'�\&+[�ѷZ�HQ��^�u�5P�y�Q�8�z�)�ݰ�3(��.��{Zl��w�lm�KC��qL��ʬ�Ӣ�:�	(���>\Y}�]{}����謰xӕe_]<��&�8�+�7��Y��C1�Ѥ�w�QՖ&!ˡZ-�pP������0����k#6$V��4��ĩ8�zC�`G/mp�[�tbj�Uӗ�+1
�T5վ#��$�Qe���U�Y�����YV�z��s���v7#�5���Q�VU*� �vsuH:��5w.���Æ�b1D�:��vs�׋�u>��b�'wu��I�ӹ�|�޷B���Ve`T*ƥU*�h��QU\U*j�X�Bԫ�0"ņ�
�b����a�H��m�*��REQ��"�P������8Ͼ�9�-��4XaIx�y�/e;%b"�I]tV���̎%pG��fk:�%1�����8���k���9�{�2��A�O{���ߌx�y���3ڌ\���U���k7M0�������O�Mѩ<~�]X�Nz�{�v��\����cӌ�Z���:-�ʲ�`��s��w@�0j������7�u{f��^{Z% ���j�ǜ�u�cC��>d�:3�U��T���4�4�-�Fi�w�Cp!/>�ivL�m)k�\���I~F�����k���N����Q�
����
�ӷ_��~��Z�����	�f�Ө�x{T�4g��<��ڗX�Z}����'˻�uSуn����l9/N��'Y���M�|{������6��:�P��-�L�3�qBu{<�*��f����b�K6��^�	�į�֑�2�Y[���[E�����I�{�ĝm�g{WZ�W\|g�%wJU<X����T5��W=��~%v���+B��#��U{��X��xh[�Z�2m?�Rɗcrh�A�5�B/_l|_�1.ػ�c��'�?�Y0�& h]���-�Q��oD�ϙ�'�h��y���.�O�kf���fӞWkM~ͺ{�u�]0N-fy�νz*(���!�?8�r ��'�qs}��2���ܞ��(ͥ��(OY�0r�Lm�|��y[�e��I�ș)*۞�穎�Z\v���~I��;ئt	���j⻸��=L��B�x�g�xx�I[��N�(��R��TT�+����NU�X���>5�멪#ny��YGT"��Z��Bi�3mgt�yw�[2(�p�5g7�7��q۠�;�6���Ot,��b1�v�]�C�;�AYE�w�)[���FM;U!�i�����wG�Չ���ϱpxE'�Dٿ�\��:�8)^��Q�.�}N;�Ͳ���CձM��]��9����϶ܻ�7/Wu�h�t��V��`.�E@<{+��CyV���k�;�����|�v� ���\iz��̧_bSʹ⬯poI�6>���^�������1ʖ1Lc��b(�K�uԡn�g�D�����R�Zřm��9[9�;1:��T6ܓ:�M��:���S�Ti"cj�"/�}����Ǌ�ՇK��W�.���fm�>�u<�w-����ڨg���M��v���7Rl���_�l��t���⾘�|���MI����7�ECT�f�&5w�p�c����^j>��^�>E�׹@��\@�=�4�����WJ�%����Wh��a�^�<|J��E�ϼd/5��1f�Ө6�5�^l��A����a��V����LZ��ט&k�ӛP(S'ԡ�:U۔��V�ٹ%v�I�2J����(iƑ�-|��S���O$Sw��Յx���W}G��`��W}�=YA�9��j�����;PpE��W�8�`�&�{L�$��iuy��n�.ɞ+����������q��Ϧ�i�&4]%�3+C�i�^�6jz3E�cDo�*�WP\���d;��i�z�������鮄��i�%������Q�f�J�B��5��B
*p����6��ۻ������GPa*�9ܶ��t���.t$�nv%�O���9Vr��[��!�JL��D��]{���u�3��xf��s}��y"4^:��㓽ˈ�Z]��'�����i������-�:&��̙^H��&��y�yױ'M�����E��Α�YΎ���b⢒�^K���4�^�Q=~����nq�QwX�Z+�9��n\���؀<6�b�����3�%ws`���T�����S����LK�p���6J���+ڝ�rT^a���`L7[��G_z0�NUٌ��:�n@f1�%��P�(����t<�s�+�;��H9�[1�r.��Y�N��L����OE赮D\ܶ�9��<��\���уU�	@�#^v��11l�c�̍8���w2�̇`[g�tWwS��� �E��,Ek�v�ɩ�����M��.��i�W�Foo4wѵc+\��ǻ����o�\C���cK;���O	��d�b�{�І�d�o4<r����!.|���\l>���+����ܫ7��}l��U2Z�,��hmΚ�\���,k�[�Vu����(&e=�;�y$�A��TF)��;o�����S��{���右���;d��@��#3�]ә�CV����|[jcDOj4t�p^��ӵzӮ-a���S�����a&�X|�%Yca�/L�ZG\�ͽH�yחgh��v\��n7�y5�=��:X��fn�=v�w���� �r{�np[�h(�G��3�~�u%�
��7�xOv���zv�J�ʭ��,GU�/|��^6�T_+&D��"����X�O}��c���T�ܖ�����3/Z����2W�9H�����/$)zV�"l��t^��!�:	�H_H��,Ӧ���M����W����4`g,����{�O��x#4�)Dw�|�e��i�v�����OvQuXr/&�[��٨Pu�w�V���Aʃ�\�d����nT�OQ�B�W.]�.��к\�o���e�9Ng�U�X�N��Y�M�sǼ�n��Z�1�1-�s%>x�z|�	P�H��Xw���u=k�f���Fn��p�Wt⽙�Z��NSK[7� �]�6����}u��p֑��vm�]�9��,[4+.���EZ��Y}R��p��D���(��`�9��0���A0���.�4�5����tV����M��(VM5z�t�;���K��M�J�r<{*A�RCo�h���O2���6�7�Wp����g�����\9�����V`
��X#��b8v:�]|��A�*�܎�ۥ�e�+`mMn:삮��M��V֑�e5���$�ن�yuٛ�\��&�,�-��%��=x��0T�J�nBgN�	��o$5�"Z��=��1.x�u�O.��w��E� �w�ic�E�]���I�s�1�Vcw��ׅL���f�l�g�7�����{�Em;���F��Z��v2��9e%5K�9��SN�l��ˠ��VLY��e�}�Myh=�%Y��Ź�n��a���`�3rsf�k���7B�x{�+��J��v�г�ݓ]AN�Q ��	ތ�(�yJe�Xr�m�[�s�L�%������`om>,�G�	cZ��n�.��
<�.պ��H�;����Ur�-Cd�խ��v)���g,f;�R�elg#Y����U(�Wt�/��<��n��8O@�`H��69*:`nح����+Fv��7��5�<�>�H���nK����T���KR��kZŒ�++EEF
�B����X�1n,�()EUZ��`TX,FҨ����"��,F�V+AX"�X �0TG�*UQTQE��"�TF*""a�[lX(��DQ��s���>�ם[��˘t�f�B�
�19R�J1_<33J.5�9!���q�]��m��E�L}��
���Y��^�q�;U�9@h�`ž}9�JE���d����86�}�@�{%(]�4x�}z�4�v�zb�\���C^��[����Y�Z!c��u�|����}���9����)�uz��B�;����8�3�n���噢u�����i��1��Z�c��/P~�\��m]�m���Sܐ,
��C+^̡.ȥ��GK�n��}���E�{�q�-��-1��{�Vݩ\�S[-<�Y{XɎY�A���9._�0:ɜuϒ��+�	�~�u���F�{���{h�%��oUyi����u5Dn��yaq^MWJ�C*y�x���d�Q}*�a��V�0'X����L��S�c��������V���}��WOL���Z��bnw�1�ʫ;����{�ż�"�����k��pp3���א���=6U��i�b�J�o�Tz�.�����$��+\ܮ9�_Oy(����zaJ1����X�^�8Ƅ�{r+ƖV��1��8�Om����C�溜|T��ڿ.�i����-^uA�Kg���;�܋��g�z�����sJ��B8�L���U���=ͦr��tB��Z@���)�n�=]�G@����!�M�T�f���E��EǸ��:��ɥj��l�V�zfU;Ʋ�����|I]�w�j{�o �{����1%��2�rO:�G���{�;��4jx�:��bxkycτ�×��ڂ�U���k�k
/�]ӷ�&��d�R�/4	]����xڼ����GT�Z��`2�������w=�G+�7n�̼��l����udIߓe�;졉�6�.m���>�{�AS�视�`��,�{�����ÔࢨW�b��,���i\W��<��o{�9я���l^�O�K6ӽ����"W������e^���H!�`Ģ�1C;��m1����㽏U�q5��b��fv�M��q4V'���/,!�� ��9=K��s��᫝����pn���`��U������n��)���Z�C3ZeVK�)n�\���il����������wK{!Z��Etg��;�L�|8T�P���j�ǚɻ�k����Z!vN�<!�r�{�rԮ�-�szȃ*#����z�$���L�3�5�[�WQ�b�kq�K����㸊�4���Q���d�%N)ѯ{������Sf�x.��0�Xz0�Ů�u���6�T�Ǟ�>�=oFذ�1�Ҋu���D����t�Y5��@�D]�2)BW,P\�5^�|mj�qױ���B�O7.����d�j'�SqO�i�id;[oIŭ�T�/
��4�oM�0����8ޤƙ8�M0�eʐ�J�n,ZZ�|Few���M�L[�j`�qo�f8Ui��߹$�j���n�zq�ܮ��C�ZĎ���8�sVU���f�����3�7��]��G���iVo��2��{�֎m�C�t�<wP˧��ϑv�Ԓ�7� ���7�5�)݋Yf��%�@�#����Z�6���6j��K�y�	��N��c![��Bmg,徠��Ɏ:h��륯�&��N�v@zv����e���UaSz�L�W�)����Z�NK�)HG�ֶl2�U�d_s�Q�f��e9/u椗�ݚ�0i�0-��r�k7����"��ͷ�Pxy�L����,�}Հ��z;Ϊ��<�z����Z]���h���1˵����[W|��յ����8u`s��3���\�7��x��L@�hڼ>MKAߕ��+�*�X�4�+bA��[պ�3��u1[xo�\"��OwW�M#�v�S�+r��ː�����Kp�NiQ�����H[.���z�c�mm֫M���{��ju���P��80���� ��&*C��\�p�\7F�B�
Ge>���@�����e��X��R�)���a�PR�E@��I�ež�ߝ]v��`�'�j�ڮ��v$���a���:1�S#����+aFױUﱍ���h�,~^�7�5�ng`����Tc���#z�nv�\Wdڲ�^��(}󎊦�(�y>�;��&�3=������i��Y�g/s�	��M��1n���z�t^���O��h�+�.|�n^�w�MNY��g%��7[��e4J�>۽m�M�G��4b9�[�{�R���_Ji��#�V�ҥR�f�a"����W%r@N��V��|�⦳�R��M��!��K�3͙�F��>�:�{�� �-!Q�<Γg���&�S��5��L�d6���+
��y<{�;���e���ߜ�څ(J���d���
���'���vr+�"��7��pv�����R����ķ�{P�����̷V��vg��=�Ą��c�Fm�M��G�q���_:��
�z�=������i�d�hP"5�@U���;6biN�)޽�+���w���|�����-�(9ժE�mv&�n_s%j�ہ5J�ly�B�<�Wk��5	���2���w|�k3��,h��Ž:=�Z٣Y���S���S�W�P���gڅ�ڽ�Dd�Ռ��m�`�)p4��ʳє/^��޸�|��*�GE]�ѳ�E��:���"4�Q�.ŵ��sK�ڌp5�b���g(�ϯ7�g|ϔ1���Os䰿tc޾�
	G�� �[.�����x!��X��iZ��_���B$�Y��	!x�"ɤI�Y�������2
��7`Xe�������$�F}�:�d$�BHH���BB@*B���c|٢o�D�a`ꅁ��6���C���C��J�k jB�~��!����!'�/�v���e��寃��}�a�t?��&&���?ND1?HD1����Y��7����)5;��ɿ���Q��9��D�'�F�s���ݲi��II3ؒB$�
�1�?(u�UE���u��â6,u��,��G���˚?����N����IVv��HD���e��;JJR��d\���E�C��O�D��S_�8z����S�
E��E�ܾRJ1���GTs���g�;�|�5.�a'��(@�����ؓ�k�ܚL?���L�$I�~�Ēt�Hh�-.���f���\ǣ�6��u����脐�6ɔ��*����#�7��6s��#��R���M)����p�dc�:����l^ã�{?˾�����f�IRĒ&<��TԼ8R6�rG��Cw��}��e�˦�ZE����[�ǣ.��Ub��ğ��@�K�t�x�Oi���I�p�(�~�2QG��l�44��Ox���8�E�-imD��(��<$�I�>���'A���'�6-!�����?$��
hc$mbHɶ�dd:�Bz&��D?�p��.�HBX2xY<&�I�~�Ԟ���ܾ�a�V�� 8;!=�D�$�Գ��I�����xd��/�s!�sD$�	=�<��7{ZG\��$"J��'rOܤ�����JO��؟y��{b>)�p��nM�#���&�J��Ԣ���'�Y�j�Q�Z%�#�F#Da��	!v:M��7��^(��AϿ�F��@�%���e�V�w�>���&�Y��=z�r6M�]����#<���R�OWK0T�%��6�|<C�~��23t��G���U����x�4���øې�%��GZ2�9F}}qW6۷,U��YMƓn�n�U�Q�f|r�Q�=i�Gv��TI!�'�������;���3���B$�'c�7�&I���;{l��+"�4J�9��xz/|YH�R�Q���:klD׾g?���)���/�