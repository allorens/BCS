BZh91AY&SY�o;�_�py����������  `�;�S��      �(�  T��b�@�� � U(I��I*V0       �   �{��_y޻9�Ǜ){�w+v�zl��7t�v=�C�}������v���֨�fmvv�{����܍:�ʟ5��t�b�\������N��`]�gs]:��g�����լ�W��_:�uo�^������֝�#��s�oov7�)�{�Ʒ-���ù�����,�j�x;�VjzS�����=w�9vݻ��u��	��;۽��z�Xt7��p�@M�|���q֫۸���)z�w��p7lͼ�I�z�>��ף�[ӭ�w��׮���6�� � ��p>:�1���[���s�u���7�V�sݸ} �׹e��v�wm�x��pn�{��n����pr�    �  B��  �S�*J�Pd  ��4d 0�А�T�0F Fb` �i���%6�&EJ�	�F����a �0�J<�U# L  � 	� �$@�T�di��T��OB=C<$�@TI)U!�Q� �0�1	�CL���?$�����1��$	-B�	�m�j�HHI%T/r�%'�}���|G����,��?�D�G���|�D>������8*�g���J�ç���u킬��"I$E�T���u�̶��� $v�:FBp1UUUB�@�Iq#���y>���o��u�V*�/���+Nܰ��.RU	��ך��`�cP܏1���L�Ǆ�EF�tIx�#`mƓr*�3��U{=�4A@�����X�PJ�L��be��m�[�?0O�$=$X� ��C2[,�&w��C�C�7]��9d��bë=�I���b���Z�v�	�..	��0��� �d�+`��n�"ɂh�aH�I�T��2F��,A
Y�3����TcE[������A~zI�hQ/% ��K9��M�zm��p�Ī��Y$��4]���$伒�	���i9���J�%0*�K����i:�S��d�4AҖXR�.�vq�S�K���15�ţ&I�/A�Ea�3Tj�QZ!�Q&]�ٴ�Zp+&K
I�V�^�/il��d�Eb1h�FZ*�h�.˲M2i���ueM�U�$ac�M��&R�K����BCG%�m���l��P%NĐ���֕l�2�ٻ)vS��J�K%�YKL,)QvU�/
d�d�)���5H�K����)�ʶj�Y�ݕve�O�*���(�%�D�E�����%�Z����HL��
Z]����U3���#7�"�d��Jlղ���R8H�vv�+x�=K^���-JZ"(J�:�����!�C�40�"M"Z)�x[:�g\��$�E4i��h�G����U��')&�X�i,i,h�'\��$�AVK�MQ��A<��I�K�3J�ˬembS�q#tcI�zI�6K��	��.�"���B�&�B7cd\,��!� N��Tj��RSN
t\�N��i&�x�o��)i����i[6�[�U�8&J�h�$Ś�v^ZN˹*�4�{6҉���J�%D��-QKME�I�YM��K'H:R�d�vS��Jd�d�t�5��Td�5��J�dS>�p��vn�tS�;e6m2��VU�IYJJXV��i�6DI�V#��e����vI�M4�d�V��*p�YB�Cd�Y��ZnɌK"�2wI-��M$RJѻEX$=-���*��e�vn��)�ׅQ%��,��V��.�2Kd�SGI�f�(�!�Jl�2���Va7ee+0�f��8L��p�2����s�Kd���ԜJNN0���nJ�oT���	�FE�EC$�14�zSg7J�;���vw1+x�=H#�JzN�-��vݽ8��g������N)�i�O"��u�e�KZKZ)�M��ਣ�R�	4Y-��7	k(����4�4S��Rn��dܗ���R�J�i�������Gr�%,K.l�t�Rh4\��0!���њ.�b$��CҘ�IV"�:��QR���oMq�a�jq��F��3��P�B�&���X�Lk���A�X�YR@�>0ԚeD���ȏ&�L���p�%��YZ3EBY��$d� �I����Aդ�
�!&�^a��#}���*�t�:)�v��J�)�r��,j60ƼKd�Dd�,U$��V.�'TT��&��?���0F���MȖIb��Q�!L[��4�4S�v�vU6��)�N�K:�z�5�a0�z�أݬ<)�m*�V�Ɩc*��s̒Ʋ2N��0��'xT���$�+�Y��'�&��e��)��$;J�W��ĕ�S�%���M
K�M�*��a�J�+�2��d�*J��%�b��V7a+tS���)�z��)�Ԕ9&�ѡW	;��5I5Ey�?�A�I8 �IbJ���0M?1��k��k���h�q+�)@�b�!����D�� C>,�]%�b[JF��1��١�	��,=9��!�\�2K��pN�K�&*�R
!�,�,�`�O��d����D�`�^b���&0�l����L���9��Q!�0.�.�0 �I,�_����N�m�A��AC��#Y3�'��.�wf�u�H�D�Ԛ���#C#}���*�t��.
b���[�:1�Z/q+xS�+zS�*�UR�FAPT�TW���`i>�pAL��6�d�`����4�4S��T�LE�1^��Ri�������L�Ġ=:$6dk80[9l�$������/҉1-��L4�Y�ء(!2� @��^=[�z=)�l�l�ك��S��N�d�`��'Y4�����9��4�r8/p��{Fc��	��t���d�0h<�^H0D��X�`�M�b���	i`�$��X�L1�5����BDXM��,dP,e0X�4h�cn��@b�Ʊؐ��A��C�@����1n����"�U	4,R&�b���s���
��;�F}�$�ѱ��a�/Km-ӡ��^�G���1���)�+ۅ�|}�9�*��k;`O�-7*'��2���φB\��𥄗����7s�٫η,�Y����\�W��yq�u�u�ӊ������!����)>>�@�;	�&_o����<n8?���Z����_~��Ǝ�x)y[L���|���gM'�v��¸Y
hFZ2L���W���xqU\�HD*���J���Cy��UOV�1�&K�r�0����p��Sz1���;~�(�"�goO����νm�0�%�֥+ɋ��h��F�Ww]�� ��W�Fx霙��D���T��l�14��Պ�F)�Ǒ&�w\��b�@���,��*�t�j��аK3x�ܨ��)c��2%n��,\�"O��n{"��lTb1q��fx]��/"˚�ȼH���oew�l�`��r���ݺ��VJ�D��3"ΕrmU�8��-�de��x��ud��#"TE�E����,r�3���ͻgM/T�ѧ{D�$�Sf�v�ex�T��3PB���]�1E��*L��(�����u�u�fNBt�6#M^H�nCQ���HwQ���8��Ğ5�>zo�Iý	#�uY^l51j׳.�n����/;J�'[)\�R������3X�\��is���������%�Yѷ#j�GYEiD�ȉʟ�yb|��+����i��_��9���rDR��o��۝S��^\t�c�J�lN8Q�T���=4c.T;���Y��g"+��5�(��0����*b8�ʶAQ*�^��Q�!�݊R�XD�Vb��ɨ�В0�L���*��N
T�QYv���k�($DzQ�*���E:�N2
Ș����m�����Mͻ��dM�F�H<�t&=�#]�(٨���j��U�C�kQ�u�����\��0`�E½W1>��yT�
TB1���Tm�|}�	e�M7J�FH�\��'#��af��ʋ����z�׵T'�!%����l�Ƶ3]8�!CI����؍��g`(��J��d�Wo(�Vl\E�]i�F,�=+0\�
�w)��3��ό��}�/y�>M��,��s�k�9U*�&�%��;#'��0�B�tro�uY�}n�%>�8�M����-���V�<���K$U(��T!�v����7�S	Hp�B���*����NDR[s��mE]����HN&f�u��9^zt� �����qr�S�h]�:²kaȲ���U�꒖�ˈ��8KC�s��J6��%�e�8^LdDLi#e��"�Ynr�Cu�.ɨ��N��M��)A�dD�ˈ�3�2�O��̎���NVc�'���#H&`�I��J�\�{�KB�];�b�'�fd��F�-��~4ݜ��G�&ӊ|�p�#��.�I�16��+v���[�h�'Hy4Tag�m%;�,��n��YW<B_��^:dm��tb�	���rTa��Pz"y����*RIYI��$��iRDBw��{������Q�6sw�y�zz�kI;1�2Q0.��q8v�EvS.2%(��,��Qp�#gi����*m�+��zL�(v��!��A�صQy��f˂w���j1�PYsXnԃ�(���d-h('~v�_(�
C⨒�:{2�6�RFD�6wٙ�u")�#QGLמvj�"��5)J��$R��!-N�۠�4��� ���h�å�;�=�����x�9B0!�9=,�8=�UDǬ���͐��Q6:�����EUBjug���Q�������E��U���&OLf/��4���\±��q�Y��pԒT�(��Ed�䍇X�MMI�;.���Ϣ�C��dQ����ϧAݒGd��������s�|j�,��C�&���
�^�=~={?�>�}yC�>�9|R��j���y�Yy�Օo�dG��$�e��k�0˚.��[�(\�;Ѳ�
e��,�h�Beˊ5(on9a8�ޮx���Ǿ��?��Ӧ�S_9]n�J�u��^���WQ�d���ѭ��b�E�I2��Y7L��'J���w�d��qx4��w��,Hcvײ�f����:uD',e�-�W]���w��s��{�g���^F�J�	F���2��QܸH�Q����n�XK{t�V��7rE��o#�������p����o�_C�7K��T�M�8���:�l�Eu��\����IBP�A�7G\��i��7PzBY�&�3P�1z^٫$�T����Y3RM	r���b0�i�Q2��%����L[\ެiȤ�q�]aE�l����8G��b�mKd����B{y.��"�(Y����!���ю�x�Ѐ�����Ѱ�.8�Rb�*t�}���ݐ=���e;�k�N��QF#c7�	��{0⻻���x�fcH�?Z��H�(�]����s���^�������q2�7�}�o{[�
��L����Sgq�Q1�"iL\dѩ����lD��4"���c*h;ʦ��&�v�p�[����f�!=�u\�K���e����Nk�{��H��GF���(AGJ��'ʷ�$��r�x��-�w{%Ti���w�s����EmV�ni)[�An��T���A��l+T�E$Jtv\^����n�$�ߏ�-9����:zeS�;`d�'2�f�]ʙջK&��A����W�79����c�C�����?9vJ/������ć�e>T���r|�GēPH1~�D,��|_��}g�%Y TZ�����䩬�X��S2 ����+y:p�R͏(F %D�$A��~�L��ƊR�S�*rAS2�I�Ufr�i:�?���3D��VED�]�r�$������1�T(�ʁ	�)�!Q�ƛ��5eqtΙ.��[y7���9&�_�{y�U�&Y$���%�ڊRIl��~3�p&:h���Tu�"����n屨����󻚧p���d�^n���Sc��Eݳ\�Q���lP�V�EP+���ճ4�ӦE�%c�r�څ-S7"�ϳ�=���J��z�G�>�V���Lm���^
�y�cu���j"��ͷO��UH�D��pp�s��8��`��l�w�{�[�6���H۶
��B�ki�:I,nG"$(���8��m}�wM��^֎�5ċ na�r�`H�$!�?��rM�����ž��6)ͼ_'���L�������(��~U1n��Ǜ\o\��*�"!�*�cc63<��@W��kM ��q�*'pb+��"�����\�*��>ݢ#M4��A�v%�T�%Z���X�Lu���
=FY �ƌ"��ɢΔ�Z��#�n��rq�FuL��X�j����ȇ\���m�����yK�
��ʢ챶4T���k|�m���B����9AH�׵�j�B���F6�N(4�{]oZ��M�Mt�jliݨ��L��ڪu619+�;2Ni�ƴ��3cP�B�h�u`QLƫ���Pq�{�\啹1PC��,�ȥo��.9$j����5�A�-VPO��_cA6�y�`��� ���>ƾd�?g��PG��d�Ϟ�G���h��?���C�y����!���������~J����}�����m�i�m�m�m�m�M���6�m���n�n[m�m�m�m���۶�m��x����m�޲�m�m�m6�v�N���m�޺���0x 0��� a� <��m�a��m�-��x��M����6ܶۖ�t�I6�6�m�m�m���ܶۦ�m��0�m�m�l�m��m�����n�ƶ۶�m��ڪ���x{�����xyxy�SM�m��m�a��m�m���m��m��嶒m����m�i��vۆ�n�n[nm�a��vۀ�p�m��鷮�m�{�;�����۷UUT��a${��{���wEOwwSm6�o-��z�m��l6�m�e��o	�[m��m��l6�m�e��vۆ�n�n[-��m��n[m�e��m��m����������K���c��G���x���U;m�m�m�M��ݶ[m����m��m��z�fm����l7�6�m��m���[m�m�m��m��m�M�-��m�a����;���z�t�sm���V����6�6�m�m�m�-���۶�m��6[m����r�n�nm�m��m�e��m���x�m�m�����oM���6[m����m��~y�y�<�s�y�֒��"3�PO��>����@��O�_�������������L?���?���Nճf�V�6鶛v�n�|�lz��6l�j���O�+m�m�m�v��m�m��V͛6��lcm�m�M�m���m��6�Ǎ:m��>z�o�i�o�|��]���m�1�f͛Wn�v�Ǐ]���V͛6l�j�i��m���!��t���'������P��cǖ"Pq�d���F6�x�YTv�줣j5eQ�4����M���m��A�&M�H�l���Ft[�A��nF�,	N�B�UYZn���5NmZcB���u��;kjtRRٵ�0bqh�7a*4��ks�Q��l���R�(����j5H<�HRd�u0N���Eknب�[U�@��\a�fA7r�MWɵTjc���	h��+��X�[M�v�r���3wIS�㖌�
ZY",���T�d��ad�5[�9	DH��7���ƦP
�Z�n���h֥啨봯%��Il݈Nl���]#�(�BkB�J�C�W�4�X)�mN_fj�E��*Va*jFXڵ��*T%l�*��-�Ph��`���N)hZ.\����$��`�6W"��º!Q�A���-�`��kyc�{�b�[��jWۥ��!*�h�8Ƌme�L�dd��!�9,`�:㠮��NF���l7��(�V:�
(*(i��
�(&�"jؤ�6�i��!.h��kQc���Ҫ�U�Q�&%A����CU�T�D����+HOr�+����B���B�Ӆ������f�]cٿy�q�c�}��Tw���s�c7��]UQg{;��8�1�}��D'{˻��g�w�����˻�.��oq+UI�����8��ӝ압�h:(()�<_--_�w3���b�Y��cЏ~�V�8�����jkc�Kd�:tNf�oS��M�H�n:2X�i0w���Յ\�8�е�p�,��49#�jq�.J��[m6�L,Z)ƙx
D7"�R�K$۲��r�[�b(�/,n���(wM~��	����IL�%�|v�tbj���e۔�a �[�&�%8�#j*GWm���E-�rԊ�?��q���O���q��0���DNcF��Z؉�L�U5�y��xЊ#��1}0�,,paɣ�B`p�L�1Iͱ��C�U�eL�x�>�g�ME4/�}�Ÿb�/��k&<HV]��2��'d�Y;<a�>UW4�1����0��h�Q����H��>���R�\Ġ-S�a�����$R6؜�0S��֕fŇ�l��iE��a���*'�`���#΁�����'��u�)�1�Ut��1��`�����X��VE�*躆�$�^bR�-���A����R
��	ș[P!y�Y��⥨����j�Y���s-|����f�*�6�$�!e�4-�`Z[N�:!�Ĳ�Hdk���M�8p�;&�����<"Am=sd�+ڹhs\�%�o[B�'ʞ区�����Yp���BcW�&G.a�Z��-Q8��P���9�	d*v��&��r&�@�	�-�I��7.�˹�rD�
��Q����є!��b�eQ�7�1�39�h�54��0�t�2�3�Ӕ��7��$��w�lH��+�E�zO	���5��a�>UW�Zc����_n�gZ,z�%H4xp�D�N8�:���Zq-,��5�B��m4�.Sa��
��fe��Ńn&�9�5��\K���<#���0�ӭ�X�籨��OXa�UU�֘�:��Eӽ������K��̆!�s_��ۤѤźN奾�BHJM�Q��)��b�%�jZR[UF�f4�(<s�ٓ��N�m-6[z��i>��#nGѩ=6�l��4��,��y��iϒ�7�Ť�y��z��yxOmV���M��1ਐ~KAi�e7�Dѐ9�_�!�[��q,Ŧ"w���O+x�C{g�mnvz����3Rn���b|���5�O~H\^QEQ|<"3p+F�v�i��n�T����L�YvD�t��D�4d�m�z6l6�?�I{���1H;!�((�2���G�Z��D�i�����6Ek@Pj���Iq~��������jyˌ�Rh�M[2q��bc��ʢ�����o��l���Q�֙�}a�����+j5S|s����C{4�q$NcQ�ึ��Q�w�+���A}����� ۝u,�H�L�p�e�Yg��������O�Q���%���;x�n���o2��dԐ�H��v�� 陷��ʢ�s�RI� ��j�.ns�A�S�סyA��х�,���M��+E>m=lh�4q�2��N��TO
3�ಊ=
Y�!����x4�b>	|4��{WǬ��8�^/q�b�������p�/���b�~?U�DG�'
#�8?>|?/�>á>���N��������G�Ί>i�9T��tz���l�|r�/�-��|l��$4XX�+�"��%p,��%�=:==��d�r&���I�:<TO�|7�x96_���;mnOW%<`�|����xǇã�L'�x~|�>	���}��E�]@���\�_�����5���P6��U��4��mHö,�qS5�פ�v>�I5���5��~��ӌ�5p(E�Ne�.#�4a��R"���[���I�s���x�JL��>�Q5P+ox��G��zD�����]E��xZ�W�U39�{�*|{�wuT����%O�w.���� {�wuT����wtwUT��G�������s�NN[���ռ+�4�M4�w��1W.1\EQE�,�9Q���Z�V4�ʞ�{6�i �E1�Ih�B'��lV"-��(�^r���P�$�LcN4��d���K��w&q���R�8�?�� �sٹ�s8��.n��Y��	1�%�1��C(ď�s�v�ϴ�H�G�l�b�du;�bj�Q�<���x���F��(�dB9H�`��%���!���Q0��4V����4�M4����OY4ŦOȢ�(��I�%�4�U`D��L�eP���kZ�\O"��_y@jҮ�G*Z���j�b��J&uy���p�>�ˡ���A�Sq���9��D��G�=H��H���Kԕ�a��G^��2�0�<��FZSJO\O2h���]]��Cԉ���6��k#v���oԡ�c��i��,�Ԩ�(�!T0���4U���C���Ye�7�r�̳�ő��Q���ȄY,oż{iƚm�����U���ӏs�"�j�
�n݉�dnE�P@�	)k5�[m�q��*�-�A6����Jj�N����)�������ip� ��e-Ô�ȥ:�BC� �����&���,�)m&�E��g�N����)$3C&E�j~WS@�V�pfg֖�n����)X��aB4��(��) �' �i�=OR�Ӱ�0��]'�E1g�a�	��dQ��	��5$z��L��$ ��F��#�e6��D�{��`a&��cCY4zp��,�#�3�7$������"�(��`�� �n2��D�*z�.��!h��醀�GfH�Zv6A�,m"[jRa"f%�i�#���Y�oڏlr,xX�F*=�1d#�ذ���@������\�����L*�{�>E�=?tQ{2�g�%	�%�Ox�`���"xn꩒�qĉPv�6G�i^�(@5ju`��Ǖ�9;�S���LV���i��iپ[��f"�=ft��QEX�~ή���'v���a�h����D�b���y�19��b�V�9	�+����U�ǋ�Sq4���]'�[���	�a�`
�-���z�u��a���ba�'�\�ڮh:�5���#����a��=1�m4�(�#P��1�ʪ%����RzBM&�´�R�����u��lvZ�R ‹ᜊ2�ȝ%{�p6��:��u�M��=�c�����h�S\�i�D�[�9Fc��!0�+�84���_���
��4]��ʒ|���O<����x�9��a�bx	���Ye�)7�v[헽������]s�9L�U�[�ZUl�*��gMS^��Έյ;F��1�M�q���f4ؓY�,�S�"55��Z(�Ͱ�4�Q��$�W0��)�9X 5����g��%�� kXǮI� wnR�i���5�������=t�H�1L%�o1�Vx��i����i��'�&H�z����|�Gk_ms[��W	[c	+��+rrx�@�3��Q��s��0h�$,Np��,�A�\�]$}�V�9��s���+�b'P�v�O]6�6�aٛ�I��9L�30�֣GnR�׮0Q�����<)-��2�,t٘�nVG��(����w��ԕ��i-�z�������Ne���5�UN��˪8%L�S��1�;�?~�tF�Z��Q{����0�`/I�&��H,I����?\��]�˘�~8��A+����ݚJ���FJ��b�+�_�������D�Q,#��Xt�2�wo0�t>���6�¥���L5o��0&�K0᫠����8co�cva����s�j.�b�"�L��/���>q7�I,J1�����&,%�2}A�̸{�
��}����*�G�g��=Kp#���!��h�Pf3.g&@׼t�+,)qRp�D���v^5{���j���	iFn���Sn�0{o�6�.���3��|tu/�ӗn�Y���'�M���E�Q�Ux��>Yƙśt�k��x��Y��x�4�+kū��/�lb�(��Q��Q�g�?
'�G�ī��OX�V~t����8��3�x�|'GG��fϋ�~~�"?
?�O�U��u����o�\��o��)�o�\88(-��G	���ڊX83��t�:c�3����\/��c��p�M�
��	�8@H�Q��|(�|S�<>�Bz|Ybz�	�L7��_#^�ш�vۊI��ۦ��~�-���Y��t��tT��Q܊�+�bj�����5Ɖl�Q�N������YU"?8��=;�ʵ�ۄ=l�dm�C/���IK=
b�eDZP+
�_���6��m#��cғi��9�t%|*�c��3����rPф7����k�M�j��%��ɲ7Mkn�л&�],㵭}&�6�\69;:m���^��H޻p��ǫy�-�-�':ⴷSSW�#�⮵�)�M��7;�gJqm�p���ù���	7��w7�|��\ژ�e�N���H��v�B�mniȅ(��`�zG�~㍞lQ�1
r�a���+��3e��D9 ��T1��`�m���8ժ�k�߹��{��I�pN�Q�]lB�z�sGL*�D���P��k���6�E��sVq��/ښ��&�vv�$d�qm�����Y�ڪ����+������=��=�w3ß"��wGv]�W|�~=��ݗwUß"����컻�ܒ`�Á%�OB�ODD�'��)Y�hC
��eamdP�rQ��T��A�F�huEb�xPN#j�kT����!RR4�C��'
6��$m��ݎ6��N�d��
�d�mu\��R��tM<Hu�ӊ�����D�楊�Zj�͍U#q�:9j��+rœe2����e�>�TYx�ћ���9w!���b`���kZ�Ӧlgq0iY����e��g�I6��cp\�;���_9-�m�殹���%	��O~'8�9�?{+!�5����uV&b�q3����3�8�����`�Ra���"z{!�v�4t�,���,����a��_����Q]��r`L���9��f|�&գ�JښL�L���iW�(��a�@�Pk޴�9c �VH�Z{������2�N[�	��J&��]�\����︸K����S]�Q�
GҀ�=JN8�,�7!�i�.F����yV}���H�VV�՞"i�V���ƞ��1�N�\�2��q�7&C�SSH�n��6a�&�h˸y��^#���i㶀�i�JOR�<wY�]Ũ(8y�Y.�ow�MO*v�'m1琄=&��ju��M�LOr��Z�!
Zi2��[b$py%�]�Q�Ƨ���اͫ
�La����,�Hnrv>���HQ���6��ls�
Hs�Y�fjw��a��3��g�Rc��TT�ʺ�hl������\fRx��SX.[Jh�$�m�}4�`s�I&�'SG�N�� `}��pn29R��q�/���RS�NUUJ5�I\<�N��0�S�y�M{!7Fl���O�����N��$��Tu8/����|���Sk�|��:�Q�e�c,�75�un����b�i�=[��B7"�cEu�8�;TN��U�֘�f袨QVߒūb5�	��	k&�`"FЙZ$�ph�fYr��,�;Z]��(�l�TYX�0[�7Ϫ�	��N�g�/�:��q<M�4�oP�[DM����N�mOs��N%dx������2��P�R��2���-Q%��Y�E(5$���1\^p��Th�f0쾜� ��}X��g�}��ϓ����O	A0X���d!��:�Cpa8�K53��3�MD�<�w������m�Y�B�|L���'c�Xk	���G p�6����@SC�&DM��ǔs*^Li�ci��~�d��:��mZ�R�)pUP��`'����Y]SI�=k	f�:S�N�0�,��&�:���Q�{I� �,�ψC��s�2�n4	��L4 a�z��S-z���797
���:s�J��
a8�$<Nm�o�<M��`Op�j˪j��h�>��е^@�>����٫�GC��d�dl�>Z��r-����p,w�܆��,����]�֞E4ڰ�4�8i�W��<"�"r$��7t$��	I�Ϝ��Tl̐�i�N�"Z[�S����0�E��PPa�J��W���ƪ��$v��Zz���Ԥ�d��gѷM���Ro2HǩI��r2��m���Bt���D���Q�J	m�=����}��c����J´��ӊ����7�	�s��"_޳�o6���M@�)l�c�'kҍ�(H��k�d���em�aeen�a�1A2ppA��
&�%Ac�	�h�crƫx��-�v�+�P��>�M�$���2��@�f�.��	�N�˧���ڒH��`F�m�!iI��I�&݁Q4���ʭ����~��$�q�\�@�5u�r��}GMՁ�����n8����D(�RyC;�,��=��}��1nZ�����P��J	D�t0lD�yl�.l�Y���C(E*��Í$<r���������8~�W��`X3�{kR�T&�j�&_8y�/���qWX�/��m�vT{�'BC����.��sR_��%�M7�d��>�2�v�sR���Ӽ��;,�&����>z
'DG����E~1W��1��8����x��Ǭq\_��g����m2�����g�
>��>�D���S���)x'�d~��x�|Wq�q[^/�X�]9�����M�'�	���?	����������3�zt}'I���m���`\5pap,�0xhX9G��q����V�/¸^ó����xx�^c��Ȟ0S�[�2�
�x^/g�����_��K���.v��������Jm�(D��ϓ{�Y�;�k��4�w�� n�tO}ʶnwW"F�{Ui0LA��4!�<ظ���8"�a�Z`NҖ�ZaV��*��F���ȽW�0�=tr�d/aԙ2Y5�0v�2G릧0��.�|�;�wt�Ϝ�g������wrI���˻����&{��z���w$��wt�e���Ii���˻�ܒ��b��N*�Ӣ<�:��Σ�����1����a���!���U8c��!��p���cxŻZ%��r�,i���J'q��%����9w�2Y�9kP�=UHp�� �m&��Rm2��;L<2��ۓ]$��0�L���%��c�����b�ګOU_4���D��&��4���M��O(�@;g!kq�JR�"�0'���qN��5iD�I���qO#��G��fq�	��aH�i0����ZR�l80�x��&CI��v�`ZNa0��0�0X�������'L���9L�ˊ�S%��3>nj8���_f���^M������:r��!?���d� FM��p���c�925+Q����Z�%R>��p��b��7f��	���Qj�j��Fc�*ӎL��g�FZ^�3T7�,%5�"rx��� ,�N�0�N��Y�FL���`g+I��ɂ�=�wp���}.�*���U�Ov�p����/�]��?S"כPQɌ��\��%'����ͩ��xL=2�]�Fে�+
�i��>Ux�AU0	�����i�,daӹ�*4����d;�����ŸִkMӬ\������I7\� W��h�S�*�Z4Wh��k�9M�{m�߿6�h)Kcd�%b ~i���V1F*��8�Z��8x��H�5��K+Ř<�W�O�G�E4ڨ%�0pD���k�V��e���i��q��>m�<<��$�]�*��L��N6��m0��9.�E�6ԍغ�J�����=�tl�<�C0��Qb2l����-<�-8�G�yz�Jdi�@x&�nTN�2����'�8�`!��aX�<+O^�˧y&��]2�L����=��i��ӑ����j�TV�o�k�S��2m4�ҙH�`G��I�(be�)O�,x`a5�a-���$��"k&����WFm���f9��a2�Q��YG�F���h���aX�:Ui�W��������I�ע���m�TNWy��8p���$m�=���
��KX�d�wJ֨-(UY�P�q�l^X��U�2��bvDUe��M�9di��0���W9��"���HUQR��V8��a+~�n�C%�<�$:��O�=H��yr�M��lhӚy1$D���% [��p�0�G���4\��&��+\�V�\b�jp�且�Ó�}�S0�3C����M�0pD��Y�++*+�rfb��K+b8Oi<J�]���櫉ӛ|�K�Yz�<r��<�@G)�i㴠=}{��RBN����tn��D�рew!�X�AZ�Q�%J�!�8}�G���x�9�����#i�a�o3FL���_�k���NͶ�+�i��\w��� ��e����a�`Q�$��k�
���E���f�5;��!�(�z�33-���WǕڀ]q�1��s�N[6�\$��رR5By=L�2JJL����	e%��`�D�l�K`�H)�>�K��0��')��1��%\pͦ>�L�ꭅ��!��0��"'N�I���Q�u_����X��GUW��$a�=��Z�u���t�)v6�wJyb�n@�X�b�m�w5%��~�#�����E6ysy�i�i�ͩ�B���CK�*�K��*���S:�##'km����uLr:��&���8���N�pHC�Bt�,G�tQ>]���OU<R��gC���|S�+��	㲾)�8z����җ��O
>���E��j�tD�pS��>���:_�������|S�p�c��D|(�+�G«�8�/n�iǙy���qx��o/�Ӣ{'Y�����>	��������p}^������z<;]�����r>�[G����)�%8:8_���8�.�'����am�O�����x�WO̕q�[~!�`�8�B���~��6(�@F1��<���y�������&Fp��j�J�
V�vW���^H�%�����v	��(KT� �؆j#�{�8��0��yÖXڷx7���9 ���.��^��z��Q�j�"ซ$SՇ�I�X٩�6a^B���-la�
�j.��1�SB�'&�Z��mՊ ������E`��L�wfl��U�ی�6����������Ǡ� �-
rÂ݃����j��qI�;x���c�ո�weBG�)tεu�	��l����E�@���% E^�k"�=!�gEꢱdTa�K���H5��&�N���=���7tzy���ɭ1D����|�R��,�؊�Z۲B5T�-���8��Д� v9e���V5ʚ]�9�S�9���ҵ[�+Ih�u0�C�9j��]����7&����X�#(�S8+4zI���(�Zdh��kE�D&�D`�TɑR��wӓ�-�d�q9bI�W?\0�'7D}{U�wz>q�t�wwUe��������˻�Ǒ����U�w|;�#��������wGwwuUe���<�8p! D���������չ�P�0ʌlnYnL����ER��h9p��*�,i�\����m��v�7�)k,��
���b�G#m���2F�T�E3���;��R6Ւ�emJ�< ���a�1�P6�G	�7�F�*�WԱl�mժڔcm�,����C�6�����0c�s �y%a��M�6T������U��9D�I4n���X�.����C^�h�/�yw���e��$�}cБ�9<���{?$$��%
6%�|0l�)����V��G_���!�:OCS#�aP6��U|}&a3/a���m��Z��%�a�(���&�튇 �Tu����(٘e��;���r��?vCõ5j��E�Ȫy�5SO�w���c�G<p4x�&kJqý�KplѸ�((�
0�	���uUǭ~�B�]�h�,\�� f%��y�S��o����vӻ�C�f��sR\��ҥh�pb߆ٿ�I;>9=ӌw���b[�c�:�_l��Sp�#����L��K���^5c����*���T�|�"t�5/���Ӣ�(�
x�R������< L�7
���fS��>{/��:ɰi��M�
r~�G��c����/��ɧ\$f[4�&�S�򒲝�e0m0��^�޶��ǝNsO\8������2<((H`'����r��r��2F�b�Pb�[�;�6~�h����u��i=�sJ�h���M�"���T�N*�J�N5���H	��[|�W/)��M2嵸�I��I!2��G�"6����n�r�İ�C`a�|���)M�{D�뤐�$���&��'�nI!I���]s���4J�<*����upY�\�c�p�[H1�^f�i�A�>9�h����mU����8���s`}G�UxFf�5�d�F��V�J�de�l�:���r$�)�n	5��o��Z �M'�&�G,{��M���}��g�߳��%4���IQ��M��a㤷��	�����Z�p�!�n��)��(��A4hDON�$����6�%���]�lᖶæ�ϱ0`�ն��-1˾C�C� x��3Ͷ��.�ZEX��i�Iyy�>=%}G\16�E�Jx�7�h0߁i��D��m8�6�����YvYE����V��w�2���Q�:�M=z���ᢔ���;چ�53L�E�4�:@�tn��8�`i�1.���dy3r��h{v3��U��s�0Ɠ/��a�l�q��V��G�^�����ݘ7��Zh��d;��y�G�����a����|��B"l֟����t⚳0���f�u��mr9��Zv��
)���2Z��vK5���Q�6���Q@j(�j���ԸՐ��I9���򖶕 �H64 ��ʠ�	\�SB�SIU�Qp�p�;�.Ƕ�[�Cӝ��zbH��#�0a�8��C(a�����rbP�CM@�>�(g��-0������EڿWh�r��!�;�_XԨ�f�l0p�J'� ��А�a)[��93R�1�g7u�D��=KL8��$���Lz`��[݅zH�S�v3	�X�@�`;��z�����f�ì
M�Zq09�HC���߸�FTy>ɸ�B���G""tDL�?���D�U|">=c�������K�v�_\a��)���|8����*>|">�����U�(�W�i�M?+�����]�1���8OG�t�N�cOW��xQ࣑G�<'��������\p`..2dh���<0.�80�.�	���0j6E���|8aiOE/���x<,���|px|��l�|8O�'�"c����j�q�\m�W��~]!�Y�d�8��>%3�u{��������� f1���(d��$U@ĕ�1vDCY%��h쒶�u����V�Fיּ��i:N�n:�%co,j���;ub*"=��T�:�^T^:��X�ٝZ��ը���>3���I��dv[�����wwuUe���'����˻��O=���U�wø�{����.�q=������.�w�"�q�1\Uc���?����s	�HL8���4���M�$'8�O.Im) s�R�SӉ��"e���a2H%$����)��]N��9��C�I`b\�	�20�,/o�wq�݆�#�Պ�nX�ӓ���;6�b�Uc�WM�9m57+�.e�eZ�/3���g��v��sR����EB��"�~�q�.1ro��&'3�|���0:�� ?d��f{�$OK�OQ���B�hz��O���-�m�x6�Gf�F��O'p��L1�����וg�>�&a�H `E\q�,MX�bi�_���(e��4<��o^(�Ч�m��Lwkq5I"`��*�E�]���2�U6��I+��>V�-��G2̨�H�eUA�?Un0���V?���w@�}�c�XY�wy%w�s��B�M9���!9O��3���R�O e9�[}M/�'��X0�Z��[������f�0�+�V6������f��M&�����h}J�M�q�o�������1e��A3;�-�>	$�������b☴��=�NJ������`�F�&S���f{<���o�^�N�0�+��6l4~N3x��+�(a$�{$���L�C�$v��(7���?Oy~4;06P�ѭ�c�8܈i�B�f�?���Po�:�wd$��G(q6��ӄǃE����\�h֟����*����0��&�9&�)]��V;Ux���}x���
s�m���'���T�4]ԕ�7u�r��Y��}�ä���˄���M�<��iÄ�Z�Ϩ�y���[l���a���+08NSi���`��(Q�)�f���k\�7ܜc����~�6��D��1<���Ib�=-��wNN���9g$�wWM޵��3Ϊ����ڠ�������T!S�x�+0ի^D��M�(��$�(ѭ�#c�2R��Q�ʚ��F�J
'&9r/��)٭J�M��8�G�9�T���9u������a�f%�5)��Ѯ���4�̧�ll�����'�ʳT0/��ǘ�]�cjd�.D�KsN~ݪ�� ��ر��߯+s�FO��OLR�W�V?*�������qS)���v���������X"�����XS��=��M���=C�L����!�D��s�/�/�_ ݕ�E �#"��[���I�p�*%>�7�/�u�uJ~���Ut�}�`��V��'C��C���[n]�8��v�y��
l0����&q䊪��O+T%�'jQ�=즙\Q�� ��7r	!�T�K,=NN�����2x>QD���Զ����1X)e����k��Q�k���q���D蟄JlD٭:��N��pެ<���^��)����Hy��5��q��n�1��u�H���uT'S[L8Kr�2v.���0q����D��Ơvb��f�a�eOhvM��a`{򪎧'p��-�b����Å۾̆�}`�<<Q����hS��Q�ρ<*�
��W��֚ⴽ/�یq}q�	�:x�D��h��D|(�Q����FpQ8?��W�D�R���á�~���xOOtN����=U
z��(�U�C�xpx�8o�p�_��Q�18I��`�p.��pи!��hp�8&�F�-.3���x�1�*�Z��/��G�zpN�c�l�z8OK��.�EW�����qs��/����Waq
(����p1������v�n�ݵXq\f��l��/D�n��{�j8�Ђ�KEP�o+��Cg+j��K�񻫕2G�*�w��ro;z�6k���S{��V� v>;�B;yŲFC�_{��Z���������t8[&5%rU�y]q�Jj��ܹ��q8q��1%%+�`0߯�%d]M��u���F�M�E*��BtM�i�"cn��]��~إh���B��؂jn\���N�[݇wA}t�Em���J-s�y�ǐ[�5]{��B5�v�s�����k�qf#h�5v�19;��>oϦ�o�A�B]VYZ�9d�ݗ�jH`���'`_�+�;�T�� ���R?�@��
�53�t�v[jR�-��]r���Q"n
��:����(�"b+VJ����Ѓ�[R�ei��z8&�U*��.'0�7��%&�Li?K4Z���Y��y�f��1���'�țGj|����vﹻ��9���=���UYwø�����UU�|;��=��33u�;�����39Yø����κ�;�����qU�*��)�NȠ���H�J֭�ۼڗ�NI�I"�l��+�����+լ�ҵK,����[���M?nAOmV��$��m(�*
ѡ�����[��X�S$M����[PN.���2ڐ������\]����]��Vd޹��'l��wu�
�Ej��w���j�`��{�sա����A�;sA
���,0ٶ���ܸ:��[$�5�"D yёEu>���a���ߺ�K[-������`�� ��X$xN�����u�S�7�p��lC��ѕϹ^a�V�T�������HD�t��S���'��B�>��y<,nh�%��Z�B��T܉�8P�I$�§���BL�zk���s7��EKcb"�E*��V�5&�Y���؂`N��Љ����|��U^�r*���K��q�i�]���ͪ<������bznzh5��5`��#[+��T0ȣ���em�f1FpޔQ�vf?j�UT{�7�/!4c�(b���BIl�ӂY�!�o�>�禍�U�%���enyc��JV�ګ*�u?X*��B�p�}Y���Ex!�F�z�2�5d<9ۖ�Uܪ����堘��YF�}�Y�K����('!�u�s�"�*��
��bl��l��35�`�U)�Yz��PH���o-�����(�h�4'DD��}�C�ָ��յ��~{�{���/k׼���a�د{�:{�o��'(���#�8���]B5�wK�jl$Y)�ջ���vZ�,ȮכaQa���9DRD!JR;*_�1{��K^-�N�{��c��zh(�VsUR���!�F	y����nN�����M�ј;�eUȁ�>>��9�Z֥����d�)��l�2 ��N�8?biӻa\1�\Nbv�0�>Mb��c�2����R�9�I��P`�|!�)�`�9�[��jXb��`��=o�:�2r���u����C��Ii�֫&�%���7�t�Rg)c��+jvǬc9��rj�f���iĤIfm!�r�7�&$����v�d������lkeOh���=���ii7GJ}�G.�亲��m(�Zm{u�Y]�'�Y�UUR�E����3�����m�|���?�Y�K��&�4S�)O�V�v�E��ufT��&g��e^H��М�\���%�H2��m���;$��IFݺbiɣ�-=��"-aC�f��SPK�J�G����Z�O�4r�}豑\5Ph��Їy���}4iU��}f$4���"xz3<�����O$��j(Y�mٛ�3��F���(�8�n�X�M	�Nꉻf��"��N�6Hd�<z�䖄d\uKe�[�� ㎪e�1ۓ^�Z������eCqDG�ƪa ��X����_˘{�;2��X�9��>$�5�w��h��9ii�z�l:q�0j�/>�_�T��d��6(�RQA�c-�Y�y8n��U�؉����~)J~1Q���Y�}U�=�|$$�t��d&L��FS(n�O�9UUR�a5�8z���:�e2��Y�v7��jʦT!�Lv\�M����C��W6�~?Cʟ�Z̥2|�rd�w1�s��s�M�S��nl�ÇW�q�t�o6�m���m�V͛6l��������q�n�qێ=�v����i^�l��M�m�6ۦ޼m�������i�N�m���m�;m�o�6��N�v�m6�lٳf����Oz��o]��M嵳n��cň0��b�$'U��sq�̌�_HO�=;�_]rPdn@���'p{�K�w��{h���ڍ#!Z@)��2�R���ƤCkY]�V�vc�q!3!��ԔT����e��oK7�ߠ���w�xk^���.��uy����G����v�O$I@d�\����;���wwL����g�wwL����dp��陙���L���陙���L��wwL����d{�p �8��8��n:��~�c3�?G��Ȟ	ĉ'����I�ʢt���&1&�~m��n�]��C�4��ͧS�&#��=L&�����Z~���g�t���-B�gHjh��L�uۺ�|�9���=�c�� ���)J|'�R{��0��.m�o���%�Hi��WR�dN��5�f��.��,���]�}H�t�O�&? p������7{��Z-jna(��Ze:c�$��N�0�L���u�z�cz����=Ox�R2 ��!`����3˾231�r�	[׿�&�F�ݯ����L��n��V��Q]Rٺ�����j����v&�9!�K����]�'��Le�,�P4X��M�h�Sx�����i��0��!�E���dOo]���Ӎp��i��m4�3�%j��U���4��Q"t�s0�o�g�����6���0�=�ϫ��0VӸ;M'���x$gSI�6B>R����~c��7H��:�*7_l����h��'R�'��)�XRq/��T��2�|�{�)��i��A�&���1�5��b�(��s&UUp��9�Z�O�f|M0���e4�8:�=L��H��!��g�c��g��E�I�6��Y��UEUi)8�e=�i�f�����G ��:d5��kJ�iU�N�U2�ZCY���f���v>)�kH�umY����Y���E]��=�|pɓ�a��2Є=!hM��Z!A�L>ې�~	aa����w����rf�s�i𖅶'$pr&��EU�M���m�[�zر�T�5r�ΧS��]�-�p���Ô�2{��&R'Ӱ�4w믏��HdDOC�!��������W�5����M$��4n�ֶ vɪ�aj��vSwy.����J��s����IPN.n�tR)�W��',�yWdZ�tU5%h��f�$���� ��;�z�T5P��c��A4���Em=?B��3�ҍZY�ɋ=��ʨ�s�6���&b�L'���I$#�D�=S̒G���'��ֹ�[c�XեsD�$'�V�]b���cȓ��]�<���20(��('�D�M��<~6�oW�+�	TN�@��c��D�����Ucn����m�ɛ�Ǒ�u;�$`i�c2C%��-<8i�j��ҟ�Ҍv��,RED��Vb}����N��%m̔Γp�?FG���Z~�NM�Gʮ��US�hDO}w����#��WYҾ�/NS���l�f����Χo�9N�S&f�8����UV���Ca�~�S�N�#?A0��a�H�ǩ�\I��$���s;���S�\$��Gd!
4B���$=�	�Ŋ�S�K�_��6�f)�sн���idd,+�V2�5ʏ)�-���#=�Z�k�kf�G�јI�mY��E�!���\k	�'�v�L'��Μ�����%f�zMu��H�2>��W��;4��4�f�q�=8��M8�\m�����[6lٶ������ǏU�t��n8��|��m���6Si�ն�m�M�m�oX���6ǎ�t��z�獾m�o�|�׍����m�ٳfͫ�m;m�׭�t��olٷjٳm�cm�ۇ��n.��NV�)��X6a���\����eE�J�\k�
*M�b���!W�nN��U"�$��L��V�*R�o�P�[�����h�ƾ�j���!���)��ŭ�+������-=��?M�k����qk�{U�pO���0�n4��V�������c��d`M5Y�� �[�CL�N6��T/^ڻ�nÓ#\��0�ټn�p�2Q��޶�gok}��+���{���v{|qU碃�|�ȵ�m��ج��/*��ݜ�)�����V�.�K1˪�������棏\�n���+�[��2=oML�;^���.�#O\�n
��#��Ͳ9����5`"�+q<��btvFơ��m��ԕ�I2.Dŵr>�>�i���bɲ�6���v�]��(ӎQS*�ڈ5D֍u��r�
�m�"r����N�4��yy��`�ʑ����ϵ38|�L���陙���L���陙���Lp��陙���Lp��陙���Lp��{9�s�x����(S�"x��Q=?��gS3��$=޳,ݨ�X�f�\�Br��zYZ�ԥ�]��0h#n�ۋ�ǏT5T	�^Rn�o�횸�h��N��G�P*��Z(Gv
cV-zM�hUUGimM�5ye(�!*�'|�%�e��]��)mL.=�!�J=�%i#������!C)W�Ӕ�J��e�Yu�+��NK�0�Ԇ9�ܧSg��&��N�
�K/�ҵ-,��j�'kh�G��!4�2�7�*5�N=O\��������6�1�Ҡ�i: �L3)��9L�3n	�z�!�n3,a�{�in� �qa��F�&R:}M���N&�s�n\l�._����3LL�wv�w��1x�!=4�5��@��#��vh���;UWl|�1���O��c0�<��}�K�a�0�9s,��SʯG�p�Զ��sZ�t��mCc6�5$m��&f�;��~L�(W̄��4g�����L���$�2�[��)��bx{|� �A>!z'D�%���&�A�&�R��~#��]�{9�(��h�{�$������&,�#P��	�&Iƻ�|����	�/�^����=�:}�]�?*70�X�!��b�~�zکro�p�w�<��OBb"zDזz[l��F�k�SUo8�E8nג(��:�9"�i��EF��������ɹ&��hU��7i�����cSI�[�˂�������O��j�Z�TUv���lq��c��0�˵.�3�U�!,�+6&j�"��i�-Ot�1'%JM;O��0{��%�,��n(�9B��z��!�4�DFќ��(��ys��MǒҪP��D�-��/8��n�Ü���n.�yx[y52kp��U^��
(�WҌ\j%��m�i�m���Q��]��]]�Ww:P�1g���^�]UJ+	i�l���^��%�R���Y�*gX�qp3�7��z�ħ�!���#E'������Dݞ�M�3�I��B�0"'�l�)��~�kd�a�%���3�d��e<0���Ӑ�xʵkQnw���"���<�͸��BH�j?�Ƹ#��O/�E���.>VR�8�O�H��:��1�%�_#��ƧF���c�Uz'DD�����*�	��Q��TU"C����NV�T'�x]������ڲ��fM&S��	�l�I�"5�(�Q��3sQ�;1&u�i׷�*T*��By�w�#8�O`Z`r��::�`����"�nj�ꨭ?�|S�ɕ[0nbHY�{�KA6BМ�$ť�"Oe�H�K��Rl2�}���B������j�YY�Q��px�$�!�4�F��G1D*�D%����1ZH����(��R�\��&��Q0�nm9z�e;7�`!����K�bߐxf��b�i���0�1��e��F�B�ҷ�4�a�n`�A��>��|�����6ZzH}%��-������B�0"�X��1��)9r�e���<j<L��r�$=���S��Y��HN�=q�������a���M����z]�Ql{Z� ��$��9����i_ǻ��.I�}
~�&��YP�D*Ky��:����ռv�c0�����*�6~4ٳf�V�m�[]�m�m����Vح�6m����������\^;���z㏛z����lڶ��i��6��6z�o�c�m:m��6����o�|��޼|�m6�li��6lڻvӶ�<z�j�lV͛6l�ն�m��p���w�Џ�y�W���]M�M��?Γ��%+krD{��ؽ���`HA}'8���I�٭j|�/yv{~QouM�ő��ھ{o���gx�O��؎���鵵�M�}W��B�Q�105z�[��+��*+6�#�d��r�1�bhH�S,��v�ffs?O���G�Oq���G�Oq���G�Oq���G�Oq���K�tp�1�Uq�1�q�~�ԉ�0�g!���le��_�i��}�̨_kV�����[���`c_/�"�L�*��H����2�=h�vCǕZx����bb���+.�_w�7����Ѷc�U|ǌc}f�ޮ�Y�[&��s�ɷ�����'��Ҵpcj\vHs8:��{EIUrѤ����}��9UUU�h���0��^�$�:���dy�*`��)��}M���
Ȑ���DO�h��"��A�����!D�r(�Sic�NV������nX���t��K@��T��MA�TMT��n���\�9j�I
�D�<�v���4FI�N1�ӱ��p��C��L�=2�щ�(����t����ԺUL���8�qN��8M	i(ˤ��5��%1w#k����m�Z��t%[v�6�Y�2V1\�v�ZG.C�Ȟ�<���p�1�UvǬc4�~z��Ym����M'���o����桂S��s6k*���"���"�׾��x�H�O�d������n�V3�;8�2�F�W' h�dW�7�����ݎNO�Cs�-�>Gg&���ړ��c�Uq��c'ꎵ��}9C[���Yh�Syc�s�SPs�<n����KD���c�N�6m�#
,���ǫ��<Jq�i窰T��� �B��~�FV�y*�C-��R�NUV��y��K�����I�Ud�V�NEcqw���%�ԃ�@�0�_��n��J{�;�f�Ҏ�����MϱZ����5��݇�P��U=>��2j8�㊎�!�	������{Yj��j����@E��H�S;�U�Owd�&P�5���iv<rm�o$J��`�dp���q�E�Y-i��AEKa[�����#2IHs�=--�VU����/,���y?  �)�l��~�Q�+�X����^\+y�+��x�˴��}M�uC�2���/�(b����"�*曼S���&�ۃ#B3ۋ�/����ヨ�<�VWR|t�iUN��1�HI���u�ο�8r�W'`�8!�K;�Dȓ��˄���i{L%�i��T�QM��K�j�U�NMUT�J\�6��U�ƿQ��e��9tj�Qt<%L=8�q�FgXyMPt�"I0�L���d6(P�D�M�;���,�g���p�vp���l�N��)��s=����ӈ��C���ى�vΗ|ITN)�Zj��R,2ق!��12YkwrW=���.�T=�Mp��a�8D����rl)�+��<����=q{v�ML)�1�Q4S�)LQ�	��0���P�;������~�]�G_1{.#q/� ��C����9:~����ݢ'M��i�&[M8<��/H�	�˜)�x�]J�1�*��fR�ߟ�����$HD��$�I$����E�?s���?��� I�G��l�B vf�J �A!����xKa���BVU�(��R(}Q�R��a)!H��	H	H,U �,`�,���
��
J"���(�B�(�H�E	E�Qd�EIT�EDQHjT�,���(�aIX�E$�T�E�X�E�EEH�ʑ���%���,QeQh�E���-(�X��,QR�Z5�#QE�X��b�E�T��,�ʑ��E�-(��(��Y��j(��T�R�(�Qb�*FJ,Q��,Qh�EJ,QekY��Uū��twHԢ�,Qe(U(X�ʑ���,Qe(���-(�b�d��*Qb�(��(�E�b��E�X��,��QR�YI,Qe*YR�(��(�E���Qb�(�(�E�YE�,RK(�EJ,Qe(���*RK(�E�TQb�YE,RJ�YE�*Qb�QE�,�,QR�(�E�X��*Qb�,.b#"�QeQb�(�E�T��$��YE�YE�,��QR�u���,Qe(��QE�TRK(�E�X��,��,��,��(��E��YE�QI,Qb�(��YLH0`ă#1 ă��T��EK*X��Qe(�EX��(��)%�,��*(�EE(�E�X��Qb�(�E�YE�X��(ғ)%�X��(��,Qb�(����EJ,��(�E�X�b���YR��B"�F$H���"��-,R��E,Q-,�ZZ-,��YK(�(�-,R�,Qe-$��J�X���K%,R�QK�R�,�Y(�)E*�)b�JX���)d�TR�E��)b�K�J�1HdR�K�R�,��K%,R�D�K�R�,��K%R��d��K�R�,��J�U�--,R���)d��-)T�K�R�J%�Y)b�)d��Y)ib�J%��R�,R�K%,R�*)b�d��U,R�K�K%*R�D�K%,R�K�Qd��D�R�,��K%,R��)T�IJX��Y)b�J))b��ib�JX�R�)E��%R�)d�%X�d�"�V*�V*�QK%X�%H����"#"0FDȬU��Ub��b��b�2#dFD@FD`���dI#"0D`����2$�`�"DQF�`��,RʲEB�1"R,D�TIH�$�P��IP�&�а��E�$TaIH�
EAH�"�d%"�)R*eBaH�E�%"�)H�
E�"ĤQ�B�a$z�N�����=�|�zД&�C���)�1TP# Q��P #�Oi+�����9��s.�W��'���)�XY������y������1�^����Hb�2�,������(��C�~�g�k4�U�?|??��a����_���S����|��ӧ�EU�����������?�A�$?x���:��`��'�!LB���b|G�L������C����)�����������Bxh��D?�?���$�	����ߖ@�V����>�-�7C�[�M��dJJO����4�5�k[�p>�}���W��Z�1���?���>�ފ` )�SU����	B*5j
��� ������!kL�¹���?�~��ë����I���ER�UZ*��P�(�$�-PQY����������5�~�A�����)ڥ?b;��?�~�����_�\����QUD��ZtK_����:����C���{��g��M��J������p}��!�2?��?�|BS����u����O�l���?���'�~�	�/���C��W��O�y����#�W�?8 �)�}��UD�?�,W�?N��QW`}�C�|�F��4�����*(\�|�$'�$�����+ H�����x����bY���RQ�Jh_��4'.�G������k��'"�O��  )C ����������hk�"����q�?���>��)�������:?�x|��R}C`��'�u? �	�������3���"~~R��H�h�>Bu0����)�S�)���b���&��L��}�?����>��|O�������i]$����~��� CI	��-�����-"�ߗ��? ��||Ȗ~}&������2"�����}C����!T�D�� ~C�6�E�X�C�7��6�=�H��![сȥ�t��'>?���O�@���S�`C�����-���pPP�|�P;���j]v�6R}�ߐ���+�!����;�M�������)�4cx�