BZh91AY&SY(n"��_�`q���"� ����b3�                                             *�  ,�_lP)� � ��   �`� 3a@@ؠ  ,   � P �   �      ���PDQAT)>�"@� TH�	JMh� �ءR��!T)% H �P($	� �*�PQ���6h(P��@�4�t��"����`F ��.t(�c���=u-4� Ҟ�:г��o#u����P�
���   �"��!J�徟}oR�)J�;�U{��eR%�s��4}eK^��J���`��2P#���������
=;B�   
<   �PP� ���k�H ��zr�C�` s�T����z x�p=��@K��X <����
/>��C>`��x   �   -����zO�� �x�$� ws�{�{�}����z��c��@R>���J>���ﲇ��G@K��(   3�4  )�� 6i
�"���| -�Ϙ�����`/G������> ;��|�w�נ{�Ͼ��` �{�B�p�)�'���   �  ���x�;�П}��R c���=�=����|����H^ =�>��`����8�  ( �  T`� ���Q��C�ly��`x�{ �{�Ϡ�< x H�� �>`��z�}�}������y 2tp ( ������a�ؽ� ^��R $<��:P 4=� 8y�Z� ww @����� �   z�   7���*�EU�$!U$���d���#u�����z!��Cu�[���  ;�E ��   `s���`��+ ��3�9u�9�g"
�t�: b@w` f��     �O *Q      ���J   b  O�*�S�L�!� &#CCOd�U)       %=CRJ� @  � � ����L�dѤ����&��hf��'���>����p}5���<������w>޼�G�����{x��WG�����$$��QT��E�������WgP����g������#��E�.����J%_;\�?�*�U��}�����j'v�?T~��~٥��Fe2����*8ĜdN2��D�E8ԧ�����q�WUƪ�b.2��8®2��Tvqң�	Ɗq���S�P�Ȝe22�v��P�(q�8�<5)�P�*8ʮ2������a\d����(�+�\e�eƎ0�G�2q�q��\a�ˍ\e�j���j�.�\j�W�ˌ8�Ɯj��j�N5q����Ʈ2�Wq��8�Ƽ��\a٫�\h�'8Í\h�G��M8�Ʈ5q�8�٫�8Κ�Ì8�Ʈ5q�ٓ�a�;5Ǝ4q���彚�æaƎ5q�-8�Ǝ�\a�aƮ4q��j�3.5q�q�8��N0�Wq��8Ì���e嫌�Ì�ˌ�ˌ�ˆh�Gq��8Ì8��h�W�Í�q�f�0�2q���h�=�q���2q��8��N58�Ƨ�8��S�\d�G8��d�GN:�4q���d�f�4q�8�Ǝ5q��8��Y�2wd�'�ÍN5\j�L�q�q��Ì8ˍ\eƮ0�<4�G�˻2�.5q�q���ӌ̸ˌ8Í\a�.4q��˦q��8Ì8Ì=�q�q��݇8�Ǝ4xh�0�4q��q��8�ݕ�'�j��8�Ʈ0�G��4q��a����N58�ݣ�\a�h�Oq��8�ݣ��d�Ǝ2q�8Ì�û2�2�Wq��{1Ʈ��Íh�58��W�it��.2��q��q��aƏ\h�Gq�q�����:j�Wq�q��Ì8����\h�'q��=�8Ì8��g�\aƎ5]ڸ�Ǝ5q��8�,8��Gf��eq��wj�K�N1q���0�;:�4�ʸ���f��ʏRxb���q�hN4��D��Ht�Ơ�UN1��R�j�ْ8�.2���fQƪ8�N1S���ydN1')�"�%wj�0W�ƒ��Qᢗ�A�)ƥ8ʧ��$�R�h��
q��b�I��)q��0�*�UO(�J8Ԯ4'^+��ƪ8ʎ��Rq�8d�%Ʃyb��8ĝ��I���ߟ�w׏o{�����k$�2*�[��[��aC���1�jgo�{�P�|��h�7l��j!�~ �oU�ȥ-�N�)���G���������XZJ�t��hɳ��w������mOv��z�X�^�hV�]�I��Ѯi�*��1��i�D��XO��v���f�!�i�q����V�k������XsT����Vt���7w�P�y�2S�����Ԙ$��{zF�r��Y��G�K4�{�5ʀ��X��ֺ��-Ky�c4�c�z�I�qI*\@Y�B�y�b,���2��2��m��!iӨ46���g1/nA����"����A��ʩPh׈���+^��t	k�Ю<q����89�}��ͮ�m���[J��"�!!����>�<0i��8���L�z�����%�N���Y�sg�%z���� �\�:�qɓp� :Vt��B�v1:רb
b{� ����`�ݕ}ҭ'��)&� R��<�un�]�(ԊB74���g��}a��n�W��y��Ķ�n�\Y�l*�ޛ�o^�κ�U�&�C��5C��Y�!��4�V�Vk�ֶ�Å�����v0�d�2#t�x���~��]�L����
�u�ﵪ��Ç��>��p��on�'9Y�f˪�*:�v>:�H$���`\v��
�Gx�۶B~�nYԨLwx����sh�.o-��{v�z�.���9����0�=�u��4�.!Iqz���f���dҧ=48qu���S�o1���cw�{�Qz��]�?��NGǬ���x��S�r��)���Z#c��6Mffǔ�уZ��iZBX��ĳsn�ͽ4�O ��;-X8ov�yl�Ɂ�vr��L�����Zx��oVe��c���*@mNmX�������;l�s�L����2r�ʵ͝����tΖaе��P�o2D��K���@��bB�{�,p[ ť�'+ܖ�)��S�njw��n�����	`<�!C��l�{K���v;�	�����݊��4�X�	y|/3����3b�gE�b{r��sZ8�������&v���w4�8hs�y�n�W�'��B�����i�����ێ���cͦk+]���B�sID\����l��oB���H��twZ :�F���O-�^Zn�Gk�.+UL�y����+JH@j̛��`���U�ܰї|��H����3��͔�x��BynW� ��hͼ�N�y�ɠ��[.�X!M���'�pV�Ӽ� ��MahZ�d�	�b�_���<x� 	.q�i�j@s��a`|���@\k+�;�ץaԣ��{�Ψ!�9�r�+�@���Z�����[�vr�r��[��V���v��L�=
or���5|�f����	`�d�V|{�����JL�ݺ��F���v�౭sbz.��61+�٢h�!�t�tX&)!�0���[��j��;��P��gN8h��O@6��2���U۔�z��p�:�K����6eE�e��7B��6��x�<gN ��bŊl_B�?��=V4�[7F��ǵ�;��6�F���ughv3�G1�Q�P���Q[ڱ�����ѳy�Wv"�V;�97~|w���z�B�Tv�L9��a�y����gV�6r���9ǥ��s���=��{Us<�Rtd�5�v�l�ד`���h�rE�%�'�ݷc���O�Og�����<�QMH�0���ݬNy��v��ݽ�j�zl=ǲgoq���S$jCR� M����AX�, �c����V�c^��2�4e95�C����WsC�Z�0Q���N�Μ;��Ι'-���#m�w6��.^%Ŷf݌!��۷UH��c�M�ˢ9ˆ1a�!���#4G���Q�q%>�ܔ��l��]�v��ч5�$��ۛ]���ň�>k�厨;YU8�9c��N"�GZ�`MOd��y$����w<Ea�K�w�߭ �^3/-�$�x�$����Ը�*���t�4�Z[��th��5�v��!75�dW�y�D3��wY�U�]%h��n�x���-�ڣl�MX"�2K�3t��[� ��s�E�v
8^�� ݟ^u�p�0�=S�a��W4�8鋎:�p�vI����8��x!z�̽�#�:PLh�gg|�`��/���<E�p�Ғr/@��������3gI��y9��`��,b�Z�^�t��ˠ��2�]��^�b��T�*��f����\I�:�9����)e���[2�+�PL��Wgg^������y#��z�B��ᐫ� ��%�H�-Γi���S��vQ�L1��n{��)^�7���:��V1���>��.����X�D��sosj������,�9��n�@5T�)���QОK�c`>u7ss�����xt��xV�Gw�WB'h��cG�D�x�@��q悻#��[�!��)��pf�\I̺YY`"�/j�U{�X��
f�:�8�1Z,�D����]*蕘�b>o7b��3�"3Dګor���JA��n�b����8���N�Nƛ��Yg���t6Pl�Lλ�Y2ϑ=��zٽ=W^s�[j�8�)lw����s��}i�*k8nj�s��z� �c��5��1�׀=�L���[+��{_�ϸ��껮���9[i�<Gv���kE�$���0�y�X/LwC&�qɯszmgf�n‚�8�RQÙI���t�2�7�-1�>����oWۏ_���x�[���s���6@],�ƻ�Kòi�Y1v�f}��y-;�ko9�6RM��F8wR6��U�w��0����V�C��]uKr�f���Z{�W�� �_cۮ���a�n�K�뎼Ռ��F�;x��wl<8���Q��shUC28JT�}隅T8���*���zT�R��]�� �l��`Ɩ�$QCJ^�����he�c��r�����Zɋ.������΃s���ͮ ,Z�EYۋ&�{�|Ȁ����4��U�G�z��hzn�5�E�(h�Q0M�ό��t0���;��,+g-�ۑ�7����b�
⸗�^��=� ��`�S�52���bxya��S��'��jbI�=Dp�d*� ]/�;� Tf#�3��
J�CY����w�]�4V[|K�E;7G'[/�k_:��v��|������=��k����j��� Y��i�M���)�*��
��t�� �S��j��=H|��u�]���U2���t
V�EU��Er�v3�Z�s^�9��>U�77��aҜ���tذLn��n��!���q������+	̹:�mт���ȫR��~��}:J���ػF��ƴ]�
Bp�r�]Wk����G ���ja�{���a6:ʳLs��Ѽ �{[��17`5k�pǄ�z`���J#5f�{:��	������*�w-;{�ȗ#yak(f���o0Jʃ�8�_9�z�2U�넔
k�V��{�ONE�&�ݩs[� �h�[�1=΍\��:i\��]ۼ��WQݜ��7�'f��ձHs��.���6��c-t|��d�s���{]S[���qV�{����86���hÉ����G�JZH��v���9;rn&�@���9 ��a9d	�#���������[x�0D��ݠJ�*F�3a�v��H���q�ﮬ��I��N�Ki��$���A�״�ѣ��ٹ�r��:}���º��G�;f�vt�~��A�i@�z�6]��w@dҷDX�v�uO���\�m��ԯp��=ɇ"���4�q���u��x�3{�3���^Sq��A���8���J9�Y�L.]���V;�Q�z�,W	9�DÄ5gX��Wd����;)�
&|^��=������ڳ�e�uB��X*���7�9WY������-�4^��
�۳i�.<���wZ:�@�-]ao�9v����e��;�v%�c�d�uX�IӀ�F7�!bdL�GB�i�>������rL��w���8�W�re�>7��*q��]C�2I�q�E���@I���xs��d˵7��5�>�,�ɸ�!�n�XIW���QY܌xrP�YO~����Y��N��D[׆���۩���!s��\�X˵��&fr \�M� Wl#ou�Q�j� �ܾ�lM����'12�S^v��{:	�f=�S�kf��^���e߭�ô[6�ɧ��f��*$G&�s�׻��LK-��Q}q�i3����q��I�v���ׯ,ԭ.�0Z�m4�g>�7%ٹs��d�ܝ8-��~]���`w�l�Ox>�b�ޠR�ע���c^P͇f �1������N���`�AK:g����gh���Zp�B��3�_�F���ʞ��A�\���V���W%�8�6r�ג@j�5!�Q�X�Vؙ�_�$���E)ݢ�Z�HLLic��)��2��k�3smi�tcb��?�rβ��KqL��vU\Uo�nܧ8���"��ޒ&�r��{
6�+��q��9�b8�f��U��*b�<9�`���m@<sV�5ͽs�e9qp]�ñ��j�$�J.���LI��O�q�Hb����F�L�.�Ct.x�f���n��_�����@��w�v���a�*��W�u���RVE�1ƦN�������=,Jݛ:��8�F]��7�A|&�\n��)V�`0���`���^��2¡�É��=.^Q�J]���y���{����B27"�F�i���;�K�j<�BC��E��>�V�[��wZb��i�h����Y	�n�l�׽��7p��H2|#�)��&l7�N�^	e��.��ۈ�<iZ���:c)ݽ�0�y9���|��~�fk���>SI�7Y3%6U�%uH��
]�&(�J�D">���^�e��*`Ź�p�Q>��4A�%N��>���YOpsa�w[����|�r]����I�,�r��Lz����Z�*��7G \=1AJo��'o�MLQ�Y=�w�f.;nD�C��$�������r`P�8�����|5����eCr�3�����ۻǔ���}�ٗ`�T�Żq\�hE�������Z�X��h���d���{t������՚"!ßO���ם��:��[d�����z���ظ�@�lf�u������/M5�0l#z`!�Qc�Q��kN��<^�w��f��G�X��4v�cm9�������Fq���q"���*z#~]��4ŧ7�{��g^��H���H�E����sC�[��,�H�N�&	���s:n,MI&tg$�7�P:��#y��-�Ov�>��s&�Q4
�6F���Z7� ^l�����Iru�N�g-T뀘��&6FKR�C�!�q�cyBI�]N��d�4��
-=�攃W�@�=˳f��Rr���V�/d�T�n^N����Ъ'R��vmq����K�����VޏY��	S���;��Ҹp�$�FI�zs�sw&�Ó�<ZF˫�ݻ���Y���] ˎ:��ɛOQ��˃��Q�ݴ�53�F1�d��]8�݃��Y;�ԅL�B0@Kk���Z����P�t3G%8�á�f��%y�Q��<����!����y��'B�i�9��ӝW��U��|��]�3e˜�ќѿmX	�k��s:�s���p�#zn�#���&56�{A0q���	�Xy0v�&�
T�[V/�����g�ǻd9�c�1f��+rnm������`��;�&\�z1�9�ѣyˠ:�mhq��툜�#���:y�8>�7�ǀz�$f�<j��������\E�1���o���ԣCyh3/IR��4�y</�I���h{3w/M86�!��WOU��u,�'>�Oaܷ��G��ڛu�~��W�{�*A��N��S���nP�7�[��G^�Q[rIL�5�/DeߵsG5�����;�-l�Q�){�B�YV����}���?�wT�<���1�s�2�4�	���:VA98�Ƿ�p.��v: ��l��D��1�"p�zΡ�ķ��\O{3w!�+���5�Tt�Z����)ćI�N�YQxP��I��Ϭ�x��x�{/2&Ό�v�x�a'���o���'J��oE�JB	��忼�ܽ����=0˚u-R���Nt���Cuw.ua������}3����`Àg�,�wvc��zK��أ��^BzgF�7n(����]`o��Q��Vnh��^���y3� ������d� �D�m�3���{%[�GȶͲ�ܕ���R���0p��F?S������ճ�&�{<�6V��,�G������x5Ǉ��9�j�]�m�T�1&�'B�e4�"��ԷPԑ�{�88�VUr�7j)�&b3j�Ö�^��9�a1K܈�0Ĳ��/&�#�:�np���3 Ǉh����Arg�ՉS6�b���mi|�)8�&��2\����oXԝ�!��.��G�Ϻl��%�.����xn=���G�ݲ�� ���9��>�ض��+Q���W�x�鯣����a�9H{�l����A����ſg��ˤ�5�lK�i�N_yr�|��f��f����Oq?��?'��H��{����<��|�;v�>�(�+e�Wב֥��M��.�WY�U�Pl$u�-��(���I6D�U֫j'ZHڐu��[IM�K���+eT�U�%����e["��[EmWZ@�*M�&�ڡ��T�UIM�M�6��JlؕlKj$�F�eu�Z�:�)���HR��Vº�N�Jl�]j�M�)�Kj���*F�l:ҫ�$�P�)�!���N��N��[M�M�Җմ�	�lCiTu�֒[Ql���mI:�`V�6C�� {�����3\�%���"?+���b�q���zC�['��5��X���S�$��>���
;�8S�^-���sQm�M�zuc�1��>w2d~m��zg���_ٯW
p�%�fd�M�9�;��+,����ń�V��L"/ϴ��_mI�M�d�mJ2�#�<K�Q����cM�B�U�X=4�p�����i�X@Y	ǚ挓�F!Q�sX��O���p������Q_Ww�bq'IK�3�6`S2���ߞ����Ztu_�q�)(����$,#����^#�	����Ho�IB0�7�7���Xi������8R��Hhɂ�ǉ�ꘫ��%8��G�!��H�"an4ujp�Nz'v��QXV�21�s�ʶ��r1��<��qLŐ`�R�t|�����1�m�e�,dgr��WX>B|�I^\{+%(�t}��t�X�/J�q07o=��IB����;(�7���ǅ���D�_������?����z��}?7~�g�������{s��\w��Sa���v�� ��q�Vn�=���u�juh��Gޞ�k���Ι�����y��r�x;6#�w�\n�e��s3n;��yL�}�h�=�<�O,�*��s���%�^	i�6١����n�2)���{m���w�_2=�g;oз���'.��w����������=�b8f�l�vu|<�]��{���	��hBNzy���:=��C��������8��4��z�F��Z��A��o���@���˒���<�h0�^��N�;�r�d�y1|��Y9`��n�f�<�'d�qBj�47/�ܺ��z��z�҄8�w�v��W:�O�'�^g5L:��1T�eM��0�X�$+,Q�QMB��N�������Q� g��"��/{�?��BX��Y~�ҫ>[�Y˽���;�[6��=�1�%5�
��x������s�(��.h�C������4\t��H��ܒ{����t����X���A�A/��V6f��w�Y���3|�����wb�v=��{uT��s�m3���O��z�;csG_^9��7~�G;.,���n�H+z/Y�ظg7<�toO�,k����ni0k9�5U�ތq�������o���47�	'�x���sH�<�v��w��Vp��w�������H��!�sL2f[3g�8��`��:|C�N��ӧON�=:t�ҝ:t�ӧ�N�!ӧN�:t���:t�!ӧA��g�gz��y�wf��N�z���@���з�f��3�/�u;7F
{��ڹe>/6���zy��#�\�m{�hc.�=-8/��=�*s�x�#����({�9��Ŝ�����h�O�؃{���o�Q����J���|k�"k~��5�"����FS�t ��<^w9o6���\�����3<JA�,���(3���w�٥E�\!Oo�t�W`o6�nI�0/��p�8z�N=���}����R���7}�8[͚x"zj"���ٻ���~�s{���5��}�*����'a[��5%�ӯ�z�Y�vR�9r�`����Q�!R���������=n����^4cg~����CL�Ν�2����p]I��E޼>/j�ݞ�������^v��_bS�ED�}X>�G�G�.�E�4g�8�໯��f��0q�����>�]ӦLK�S��>7�8�>��"���7ψ>L ��٬���i� 0�C�%[vP��v��<�%٫�{|�w�ؼ�3F����ۅ��dD��XzdK\�#��x-��y�������> vWY��6��rKͳ1���h/n�
�������C~�L����c�ފ.[��q4�s}�`�;sl܇����$ rN�m=c�n�[��^����l���ОG��wH�{��.�8s�	��.���9��&�e��
(P��0`��0`a�0H�� açN�:t�ҝ:t�ӧ�N�!Ҕ���yi�s"�f��D�(���O{Y>Y�trO�ޞ���'��1Q���t6����
,�s�)�%��J����GeX����a\T�8ax�qP7��3����g�������A���T��e��(��O/xp 2e�n������X���y����w'���s`a�ׅ�U�\�l�Jv�0�j�����*������8���}��������P�&(]��=3ڏ��������hV�	��U՝�l�|Ax�����˙N��6T�:�)� �w�lW7hPQ��$I�yUJ���*�b������᠄;�Z�`�纽�:Y`$��Zs�ޡs;����ܼ;|c��>�O�E5�Y܇����-��4d��mܷD�K��j^���F���o��l�*0�}۰���W��͹ؙ�O>��ݾߊ��a�`�����|�m/݃�������y�	�[H��sk��]h��Į(���*�{qadkw���#hhk�ͼ��"_� �Ǡff�����r.?W��ߎT�����pK���/����t�8���,rmJY��-ۄ]�ի�ϰӾ��wr��$����_�����Ӛ�����y2����|۠x��<���5h�n#�Ш�Fv��vC��ޖ��h;VS�s���6z���v���Ê}��/������e�˞�:iӧN�8t�ӧN�:t��N�:t�ӇN�:iӧN�8C�N�8t�ӡ�0`��
��]�S�l�D�a�zH����(<�W�*�p��}7c0�:{��]�f�s�x�q��>���<��s���F�lӢ�j�W�e}�|=ӹמ�3��w��Z�SQ��l0+�;N��-����f��o�Bg���e���L��gkH/#W_
��޻	wqj;�fb�~JՁ3pd~��{�W=�s�d��Vݘtr��h��ݯf]O�}揵_>���O;�7���^On������ƾ����^��̻��J���n{n�}��F������˱�gڮ�y������z�ʫ��x�廆p��Ѻ�պ{�\�W�����{Q��lz{Ǘ��]vOI�W{�ǽݳǠ�E��~<�N�}���6��[a�7�����l~���o�T�Rޭ�bP��g1\R�j�U���e�b7!���^Jc��c�C�4��L��V���b���%�;o�����ը�.�R~
{�"< Mσy�K�y��=^��zK���L>��[�s�@���ڣ����=�ί�dUq�Fy��&����ľ;�."4�͛��w���S����(���̠}�u��4C����s��>L���_��x�[p�
F}�}��(�{������=�]�������Ow���X�J�{�w�f��q����4�5�N��J:\�{���s����ON�:t�çN�4�ӧN�:xt�ҝ:t�ӧN��:C�N�:t�ӧN�t`���8���2�&p�4̃|8�o�XF�G����UN�1�}ږySr����y�Y�w�<{3���3�2�3\�^Q�}�c��1M��V
�䌇-��aE��y�w|Up�p~�8�Җ���ܬ}��(�\�nM�c�;���ˈ1u�o���Qݵr�}!d�#�?{��+x�W1���2$=�������?m�3{��'��D��;��߯z��{����^�6{+؝��_��R�O{=�3��ٓ�.!�a�b�S������~{���Y�Y'��+F����@����h��.�`���!�1��~�O�0E3.0��j����sɦ`��J�&�|���=���V��l�j�����7��)�ol.� �š[�g9�s4��-~��@�7�x���Or���C����BH����s{{-�G\�?	w�a^p�*�^������m3'��,@˽&nH��;�w+no�~���N��F���%��L1`���s$�:/���%޳�7���7y�u�z�v�}U�bk�үob�I��g)�Lp/p�w�v��>/)i���1f{_z���?L�S��F���^EOn/(�*���I)�
^���b^��͚r'�ٿs�k6c����0x@�q��yuk���3k�XǓr矙�]��@�{�@>$��~���ע�flA�0@���0`���!ӧN�:t��Ӥ:t�ӧN�:|tN�:t�ӧ�N�)ӧN��M4�N�����`�V��o�K�fX͈]M��ĀϺ}���^�Ҥ�.��1Z95�^ݞU�^?>^k�]Lf��r=g}�֞
_U�:=����ߗ=���|�j��2���¡w�l�dק�ѣ��xC}�pPЮT�Ǿ��q�8;���!,��K�M������s>���!�H&f˾��[s��or�g�"���#bi{���FSd�,�'=��v��s�}�I٠:1?o9F����ng�� �n.!���c/t3�V>�Y�Y^��l5�ܳP�yo�eW�q3=�ۂ0e�������NМ�zL�7�M��3iA�x��ýK��O<CڲQ.sey��U�,��<!a�.ytÐl@<�Hom�Rnk�<�=~{�)��@�7&��d�l�=J1JV�����F�T�5���0g�ھ^�g�w�f�ӡn�� �uOn�P��G|��YD��5�(���p}����?'��w�`N������k�U�^|s��6��CY��{�����]yV�����k�/���g�yk�|q?�n^c��|��/�=��^�A�K��u��~�zzp�k��G�8�zOgj8��;��n��Է{;g�N\��ᙡ&׺y��i�_;��ž��R���y��W������1V��%9Nj��8�O`�g9@�����0`���0`��0X�F:t�ӧN��:t�ӧN�::t��0`C0a��0`�u#*����ca�h��y�l}����������U�<<5�pؗN�|;4�8�f�aq�X{�����j���d��%�9��`�>l���<.{QAe}�S�2��<��xx�#�WZ�L������,��f��@3�?��e�6�3s�[���]:kf�p̧���)%�z��<e��@O��-����7w��׼fW�c!�qӾ��,[嚼Ob�A1�QJ�����d7�U���On`��#����wؖ� ��L�+ދ,��^���CNo�G(\${.M���=�a1.����|�5����V
�XD<l��G2E��\��t^Χ&��)��!�WC���4�}�΃Nhp�3��5����<d�ww.�'��@V���܂�$��#���H׹���/����NZ���y�o^=����}�{h�d��h�z4ۡq�|I4C�jP[9~������Ɣ7�K�a�2�ǳ��.JS�h]�����i�o*��;�#�'H���wۈ���Y�� ����ݸ���|�O��׽����YO oY�QP���xd{�([a�	|j�3H|罦s.%��� �\8�����+6��SO�u�_��;��!��aF����Kzκ�p�����P�~��t�B7��%zIp�~~v,���hŨ��뜎3����J��'��*��/����&�'����4�.����;3ۙ�q®�Y!��,@�"�0`��0`0t�ӧN�:t:t�ӧN�:t�t�ӧN�:t���ӧJR��t�ӧy���#�Tvr��a��Ȕ��b,�{��^l��Ą/}��^��j�����ö&bXs�9�ܷ�����5=����j<=N��g������,�W�hø���{<|��g^��mʈy�=��U2�+��>я [s��uϳ��_�+}�Y���^]��gT+]_^��W�s��Ɗ��E��4{�}�7���x_v�jշ����S�ꖺ<Gz�@�<+^��I۾|3}����q��!c��L[�G�{��$*7,�b���+W�9�i���=�)Ɏ�ϋ�n�X2_7�z؎�;�I�C"T�F��r���wU�t�({��䳱{�%�!��S�deۺ-/�,�o�����7�f`�����s�����	��!���)b{���nv������*�瀞�I�#͎�a4Lr�zʽ�TX}/����zO�s��=���?/o�fLQ�ȱ��vn	�9셉���6Q�.y�f��'v#�K��=��8��곧;Ü\b/�{˴u�r�⻮1�����4A�g���4uH���e�C�i�F��ᛨx>�Rז�	�Z���xA�j�qN��!�$}�*m��G3!����������3�P�k�[���I�{����;��9�s	��<�{9��5�v{�X�x����^������O�Xv����:3ٙt������<��_WǷE��}���;Z�1>�׹���}��B�g��㏦�.Ǔ��g����L{�7�}�6|P��'+y�|n\y�3ٝ�0`��00`��0`��:t�ӧ�N�ӧN�:t����ӧJR��t�ӧ��aa϶���w���i�"Yw1������q�9>Xs�k���n������e�k���{�r��7ֽ��>g}���2��xߔ����#L;ٽ{�z(5�q�3 ޑ5�(�v{)��^ܗ��b��������!�-6o�s;��ن��׸"�h!�e�E�2۰����wl�[H=�w�NRspv�3N}�A��y�5���yrasiG�`92��|�-��+��Y�j;�~ż2QE[����8	�1�ռc�� ���=�f�����˯���4->~�/y���b���q���]u�Kq���x�y�������KkEi�'��|�i�f�x���+�b	/b���ϧQOrܾ���-�x�!zmy.��׋�p���O�.�"��{�f!;�E���C[ߙ�u�L0���|�o��pYڑ��1��)1珀��� O}W<[&nqx.��_qq����)�aB2џY	�^@dZ. }�^�`���Z�^@��?5�\��X�V���N�v�PA�JU�׽��=������g�N���y��w��]����ř��4q���]�;�g��8������xkğ4vhg��������s�g�Ovl��_i}>}�,�l��%���ˤ��(I�¨V+@'
RŚ����l��E���5U�3��7v��J͑����y�ktӾE�T����M$	:��n��9g�������=�����!��V�I��bdIfq�t�R�cN���lp{���+���C���^���S�}'�a��S\�����n��\�#6%����g�*�"���E��,w��}��H��w�
�ǅ�f
|�N�t��۞�{�����������o���RT��ox* }�W��F�������w�o����d�N�F!�)<s�Գ{��ɷۄg�����M�2&���H3�	�o.�S���{{G��F{W��:���<,ԟ/f��p�^׿ �����\^5���f�	��_>뺼�+���[�ݛ|��6��ٸ�"4������J�>��i�
�q~��6��W���=�e;�L�Q%B|��+���&��4{^\��ۛ�p�����a���X�2{������O3��"��vo��R"�^ex,�o-]� [��x�;{y�lC�ݙ��8}�����~,p�����-E ��ҵ�"1�jQ$y+)^����G�٦=	�@�\�M�6���d��s{�9��އ�^�N��{o�>�.�8�nu�&\W�{7ޣ�.�)=�ˊ�	}����%|�=�/y#�=�z�t���e������@#�W�_,�͛�I!�-`/WN�������䉃��_{�>��n܂��w�
^f�x^ۧv����c���W�?_����O���ꊿ�:��H�����JP�6�G0�	��GDv]�5��f0��zэ�"qT�k%��*ԛ�݆-�z���=����x��X�ʤNe7>��W*�ϵe�M�+͈�Mŋ���i6�e�a�p�Z�<��!q�Ujŵ���b�8�q4k�E��B�u����6�y��[u��<RZ-R�̥[��vGT�ֳb�z�'	&ú)-�ax�X��<�s�MuRl>{S�]%Q֋�k�7O�g�)�#nq��U�Ŷ�c�n2y��v�*�&�d�H�&9ZJa-�ͩ� ��	8�I7gm��]5�8�u	��hEɶb��k.�˃��2�8�m"C;]���6�	j4I��6#���Y����:B��a4�1l=����<��^�����G[ǵ�q���=n��<�vL�z^��|�ˏK��n��Σn{��6ݕ���0n�ۣ5�W5�nx�K���.�w ����! �̤*F2�h[��e�&���8zi.݋��$�q�M���-��a]�y�z��ݝ���O�m.{U�M�ø1ښ���S���6�:���CP��ya�[�YS�Y�護7[�n�4��1�tH��y�N�����l� ��=��v<lOk�vl�+�W<ųس��7ռt'Ex���#vWb]6%yI�*�l�,s�+���7�mcNڲ�7�4
ш�R("]UyeS�p>�/
�֜��u�Ǟ`�Ʋ����]��.��Yz6���v{����w	"���զ뜝�S�p��*��ԥG�;�s�V���q��'"=���G��6ܓ4���x�� Zh�e�C7#ʷ"�6�e�4aR��5���	+EkRd(�[9�
�e�@�q�yHՎ6�����F�����qal��Xw6:�����Hp[�J�f����98�������-�YkA�����3�sM�tDە�Z�"�囍Wc�lm�����'C�u�N��:��k\\u��4�ׂ9w����j3�^`�d,��Z��)�9�8�:ŜQ-�
\�2��!��.�[�I�I[`�N�8uϳ�n7n7�z���Z�ۅ.7�M�e1�[\BD���볧�7�]��Ɡ��ݓ����k�۵�)��2[<K��I����ci@�Y�`K�§0�%`Yv1d��hݝi$�����o�k��6�����88X��E4ݮ���C-��[�}��ۼ�CL��]��t.
:܄ñ��s�=ێ�S��,�Ds����Y�P�H�nbx�C�g��{n���4r�1�t�N-�G{EsۀMI�,=ru�a�u��p��\�t��8v�`��Q�J�o���v:y�0v�-9xn^,�t�׍"1�Ie�LC]�)IR��Y�<,O<�x��Còh��)Bb��݄�Hh�����J"SL@��Y)�X��Ri��j����B�聎�զޒ2x��ym�m".^�崶�oL�5�A�s6�m1V�:Y�9��SWY�B�Sl�@�P�r�JLF�aX����4�dN:� ���b�[h���B�(&��Տ.%��4ɠkL$bls-4��.5��d�A1������h�MQ5��k���(�x�y���ަuY7sv��m����OS�֌�����t';RP�	�z�X�����v�q�������6�]1.̇LY��W���.�� ͋n���4/���r�v0;�YN�]�Yv�iE9MX�È,��]ͦB�p@(f���]K��I����LƄ%,ړ*K�\�0ͼ�R�8a��Ms0�
wT����h����3�2<����$9����{z�����k�"n�Y�,ѵtR�غxv�,\v���M�k �L�	-l��:Mx��7����Pٺܴ�&��r��qS�L�yv�4tc��eѴ�	�s��Y�=vG���o&fm��V�Ѐcj��n:��N-n�q>tulA�y1�X
�Ս�ZH{v�
7�{#�����9q��=[�3���g�R�H+�sj�:,*Q�T��!���FNV{wŜ\`������ �U�n;q`룯j�s��C�iznp.�n����4(db���{�Rhg[Y�{[4p�.�����z��okZ���R2��f%2]V�6��p��]�M���t�/'>Ss0���c�FR���"d
$:�����{��y��=q؇n��h����0�	��9�t����8C�ʧB=S��d� )�5��;V.�v�	�6�8������f��`�y:�>�W�v��]�ۥ�[p�Wz;Y������P+����=Om�
�q�X���7=��)�B��F1`d.��y�4�mʰ�OB��#����<���9�vS'V�Ua{���u�^`��a�섑2�n��e=R\�/lt���v8��I;M�Őx���]�(uڣ��\9�u�vw�awj�ۜ7��}��A��n��Hׅ1��<n�W��f��m�=�Xض��1�M��ٷ����ɤ�EtRU+c7#k&�EmB^3e���F�M/.�`���6&M@�ΎҴ�G��=5��9轇�Čk�=�ω�4yjN��rۋ=V�Pֶ�Qɤ�s3[v��5g�k��헺��M�q�����8$wgG���i�\l�s�,����)��Z}�8�i�p���]���a-��hE�-��u�,K����/N�u�)�,=>|��X)6 �]�H:$]u��;cM�!FtV�(.1�ݎ��M����C諆��dA�̕���af���7�ۍ�75�V��5d�m���n^4����&�<s��qX�c)@����.И�[.��:��3r�� �cE[���<e����,��mGQtYm.S#p�!�0�˴��(:aH�V���)��(�t���
Va�%%u&�YC�sĬ�юP��Q��1��%)�<�:��_b�nTz���m���n��F��f�Z��(��������K�R��tr9�'`N8��m��`mU�l
�[N�blAG�89c�2��۸���J)Wb��Q�&4s!& m63m�{Z8��#��j'�6�.�ws�i�F�{9x��M��K�Q��9����&6�u��
�h�l���PT1Y�*[	KK/#F���M����ڰ�5���99L�PV�݊��>�N7<i�-�`�@JM��3ai���6u��ؚ�S�cISW&���Iq\i��ۯ0j.�������q�Ҁ��h[�pP��PJ`�멬/B`n�2@t����K��!���v�9�Nl�`�f�:�>��'����7m�n��Mwd�͝��)]0<rGc��{m�+�ts.�%��Gl���z��7`��wn��Z��\�v�+c��d&5[�NW�89��vgnx�̓v���WmN�����. ���ek+�B;k�U�m#\\l5�h��eb�X�ؐ�5t)C��c���L=�<��E���'nBgF�OnH��7�-=�Mʷ��)֌�,��q0%%�����À]�!�hi�$f]v����ڬ�W^`ݦ3&�k8yY�Ҩn�D^�Q�B�l��Xj/V�yd�N��L]�*ع�t��kmf�ձh_iН��oyh��Q#�mL�nŦP�s���i��.�ճ�/n����6u�Z�5�Ԝ��7'J�6ͮ�\6g��x��4M;FL��G�	g��q�.Ӳ��k�9�f:R�����ԇ,�%^�
���ۋŒ�]a��x_v��Yƫ���q��y�����g5�E6x�Ƿ���X�*���zc�;��9s��8�P2{����Ϫ��ӬZ�v1ҕf�9���@��2XXC����]�|ٽ��Íb�V�s�=�t�n��:�<v5��bXy��rSp�	ö�ʛ��=
��a���i��D-\�N��d�����&�[n@��]R�+ �0�#KeV�H�mΧ���.��(p(�]%��9�V��tv�C�2D]��u�$]qO���<,s��'Ө�b5ch�'cb�[v�X:�.m<fu,%�J�5�Z [��AAՔ��,5�\�ѵr���*�ӳe��v��J㗏b�Pf�K��Ѽf��s�v��L������T��$�W=olq��+U������:�������vxz�T��f�i��A�s�Hݓq[q>Gt�)����Nݢ1j[f��h۰&�/uۋ�-���"�g;�9d{e��]��U�g�8�i��-����r���a�C��j7i rWX�%h��*&0p%͊&��4͚�֌
Z:Y�9n���3L��a7��-Iq���5�Ɲ.G���ݏQl�:a���l�!�ldS��&�v�d��=�wGq;�U�N��	jq,��j�`�[��=��5sL�r�uvR����X8��Yv�m�M�kMky^1M[d�8&�i�v�B��u��1��J3{v�ĭ=�,Ax��U�6�q�lmз\b�����������(���Li2c�������a������+�v�6�Tө$�kss9[]�Aj�S:���-�3��ҽ�L����-:fvqa��[���j��e�QlEΎ�֮����� @4u��)��D�����e6�m`ah/�����aq�ό��LG���t�@�@7`.��_>ur;���s����6����.Sy�����6�x '5����*�8G	��a�U�,���+�-�I�W�
⢪�>m���B�æ����$	������ �" �e�H��%I����Rb""��
��$vE���`��!M8xox�W���I���8���H�T_l���M�K6ZL�"(��(��b*�s6�u�D�4�����e��3.K	�Ec�<ٹ10E�B<���NX|Z����������#$�HLԶ|$)Ç��sd�I9-&���

�#��'��R9"��j�Q�+ XL�c蔦����<�AO.�#ِQ!B���*�a�"Slq�n%��LX�d��u�`��e�d��}4��<=9�G?B5=�kl�^<)P����\�걖@2)�2ܙc&0��j�H����L�B�d"��`�²�Df%Hc�����l!0ą�0�4���x����+1H���<Haq�B�Y'L�DVL��\��r5�W&W&e%KP���V@� �T�H��ܰ@}a����x���q�IR�,����0DK-$��Ӈ�OL<W�g�ȤE��D�ԁY1� ���q�c���r�dA#�m��,���8�@���6�G*I Er��	0qTfLF#-#(6P-�ZD�q���� XZJ�)�#�"�BC�ka�; �cV[3�"�993F%R8J��Eq��9�﻽�}���!=xXz.�KuE�T�JH.£3[v��j�9k�th��R�y�R&��y�U����;�իv���K��Y���n::guvۦ��6��u�5m�#Bl��h�<$��r�-�v�"9z�!;T���`1%.s����Fm¦X�[)�њ�
174*$KM�b�\�ƺ�A��r��<v�������
"9�](�&���Y[sQ�i�Л<��DP�v؆�u��p�Q�(�J�l�%b���h��'<e�5�u�ث�pg���qɭ6�K&��ڧ�p9g�k5�G������eH^�1
�\����hq}Z�M��^s��5��S'v0xƌ,Mm�ݬ�̷P\���&�	����y�D��`��q��{i�!��;�����G3N�����Xlj��+c1z�漛c�u8�h%�\$��l�D���C�j�1�Xw[��<ýe�Ɓm������{�-�<Sx.&�+-�a�-3�Xk`Hfx��U��p�A��1���<�qڧ��h�{\lt�m�F���٫tOOn�x'�r���@:���dَ-�b�lQ�(W*���<r;X.L�h���Ç�nj�YɊ��!�X�⬏��N� C�[E�������ۚR�^�#�1f��s�A��[��j�Ї6 �s�5kn�[Q[�K���p�8����+v$�v��j�P+��Qy�ݸ�����K�۫!��}�UݪS�U]a	���`�Nj�wI�7�l	s�Fiw:�:�4tOBH-mν�A��.ף��rs�+؅��� �@Z��4�6*Oo%�.'�v��R�v���x-ø�;�{XΛ��ՠx���n9�ݹ�q"����v�l��1y'�.D��>s�z�kn����5[f�,��6��\���j�Z�t�Mf,�C�����3�,��Ţ�AVFA�iT��6FE�H�U-��V����H����Ki���"��c�I,�"BŖ������N �mT��`R
Z��Yl����j�mE�U,!RT����m^ �U�8ѷ��%Z(�-,Y< �[m^l�r�9�2��Ds�X�EmlYYZĥ,eR�Qk K�w����5��K>�VHrE�c��A>X�\��fL�4e���8rI1q��,N��AI���[1�5�K�E�P��z0 �f" %�C[f�$��T<-��R6\Y�R�K��M!M���{��È�</�߼ʩ˭�V�c.��
F�h(�؏-V���18�&L�k�L9ѷޢ���LH:Ѱ#	)�K58���z�ۆb��SۏC��n���wA�VPh�z��l,�b
L�55��T�5�b<	%Km� ��p���Dj�u1�'u��9��Ѭ0stR�J�`I]ecfјx2�M�!�f�ͱ���w�ĺ�Ү�c�� ���� ����޻nDD�(358�~U���
�c6�a��?�ح�p�qW�UL�v��ABb�*ƶqX�7V<(l�ǘ�f(�J�«�e�+�ˢ8�k=����6�ڷ!��(��c��"�zw�v����
[q@�@m��8�kі�qE���H%;9`��o�Jɀ�	nc6��*1�ڴ�U�
�X���`��(�]����ƞLxMr��^�A�2چ7����F�rA&j6̼������ z�S0��c
)��_ʰ�	5���!cf���#����㰰lwf Z�S�h)/ �}tM8��ܸ�m�:��,r]��87toA�07D������PEܻ��AjS��k1��Y�@�x�4�gdk^�m�kj�Z'79����Y�$_Ļ��)�ق�|˷k���u�A�
�����؀A�B
���
v�P�J�i�-u!wHNa�y���o"�~��{��q�jg���D�^O��{}�Wye#ٴ����3�����1��A����Y/�6�͝)¶%:ǉ�.��bo6�&�,K4j�A/r H"66=�6��)���A�[;���յ��j�^Y��A/PH��YB�Z��֪�a�Ԩ�������M\YA�d� ���hURV,�a
3#�`�,D2� �C[n�.u�^_�K�	���^R��E7���v�X���<��ORE�[�6:�ȀO>���kqP�-,4�E\c� �m��X$-r�\N{�����7&"4C���Eܻ��-Q4���
�)	f��N|O�E��,�
|h/)�c���D�Ь�t��D��w��b	
��*�Ҍxշ��TT�� �n��+V�2-1�c�L]�z�1��μd�.v���y�
	yS]��$�ek��E��(�ANw�����^���K��i�w
h2)��[͚vx p�{wg�����u�z�x�<6K����t}d�h�=B �z�tÖ�@.��	�_�䫘Aq��wX8.�(��m6��Y�	ə�� 2���ZZ���~�<�_�	A�
3Bg���R�o����M(6e�kR�.�Ͷ�6 �%���)�Jp�g�w�#j"��5H$�5�嗍y�Q9�d�sb�@�pSc3�}��ƞR09E�:,'^�?���Z������_fm��E���#���N�6/l6�֜|����"��wt��-�	5z���T�2E�H&����v�[w`A>$mk���ۅ�rI�2gvQl�-4'p����������:/���`b��������1�3�a��mp�v�b(L=���5n �H���H�فgHHRfv}g5LtP#_���[�y��e���qx�v{�v��H�} ��ƹIzLE�8}�}�}s��j���qĲ����'�(���6]4W6]\K�����IZ5փ6�۲r����qɂ\����jh�4&5�Xƶ:�n�X��O�u�چ33�ݖ��Ų��x�('���o1�Xyt�{z:���j"OH>�p���ֳ<��g�ڍ�qm4!/5�q%r�.Ҁ�+Kh! �c2��5�iv1�T:�Sn�qYW��v����ac�;�{H��ˋ�Gk��B��ӻi�,E^b�8�h+�����t유��
�he����X%�����S8��o.�V�� PH��hO�%� �X����vg��������v�^�$�r�Ó�u6�́ ��ȳF&j(<��z�	��p:f�0f#"�8 ����O�
x�����Va�Af`�A9V�wvb	A�l�,A��������_���C������3*b!���`q�ZLƴ-F[e��n�C�	/�Y�N�K�$��{i+��|O����L]�z$�<�u�oK��s�,���pvU��^"����/K��y9SRH�ג��Co?}��l%;���q��@�n��O���א���v�F��H$�Us A0�c`d�Π\l�x�
�u���'7
���1��M��>7�g���Ps7V�w������xym{�v®��:����U�?l���Iz�#u�������H��$��	!]V{[7��L嗾+�!<8���_�?��& ���`/yz���gPH÷.�p0�UL@$���q�#@�t���1h֖z6�����L�I/x�}v���ҐSTEe���ݲ����'	���4��m�"O�o-��4F�ˈ�&B�O�6�E��]���p�.��v>��|�cv�R��j�J����`Xla��lB�?��
���3�3Wp`Y�%�K<�n:$�l1�H;��`B�]��ݭs�����u�{<;i娳jmf���	!9��|j�i���1�'k\^L?�\y-�������X�f�&u"�ZlA>;��L I���*O�y~�y���L���w`qI��uY37�� s7��4e���Q;K�q��db��PZ��Y*�D>Ê��k������}�M�O<��������:����#|�آ�`��m�Ɋ�����1R����,!@$؜�	�%�:1����c�3)d��4�eT^�8p||I�وƆl���`�i1�ݿ���و����ɽr0���W1�GٱG���%��I�8랛�� ����ޝA�Aܳ��@-�����	'7j �:�ϵwW$��\`" $e������%�������ꐀU�V��	�n�Â1 ��9$3�����D����nwdc�m9+U� �ዸ2��G�� +n"&гn��ֽE|�$���� ���Л�t� t��	�G���>]�񴒻sX�Ry�e�s;R��M���_]��5��l����R�/-��g��}ٴsۓp���YR�6D�YV��Y��;cTLV#�K_��r�z�X����u��l�7ޟ��"[s���Y۪� xM����%���2pC�D�|]k�ڐt���;�3P�����a
6��lg�E�.�����{-/���T�0ؗ[4`�O��q�%dƳ����lЛB��Gfu���[���1f�ia�	�x� ��}0p=ԍ##f�$/3�^3OP ������l�f�?/������rX��|	�و$��}0I���}8��M�B�-,�l֐�'D�,�#6/�|Cn6B���5*/oB�T��l��d ��b
O�w<׮�>����Կ�vtA$�{>��qI��K�S��}��E��;1r�gP+%��2�7����Qg3<�QRۭWm��$@���7��˧计��~�Lf�ty�FC�P��'�sn�0��!f�'�������5.�� �p���s93��f,"%3x0���r�ra����~=�{��hA��6L�e6R^k�
q�<�m���S��ԑ�r֌nժ{n�����F8����=O��bݖ�g����l������=r�Y�y��k��9�^Ѓnu=B��_k=�7X�뎭���xq���ƮK[�ݱ�^\����(<Zf��U�]�څ�N,dmU�[Z����;k�u�.5m�3�x��n��0M�NǞZ�L�7`z�7;��79�M5sȲv���0�.�5��d4%����WĬƞ��w*�v�.^g��LaY�wM��a��_���v��@3���M4�l[��6����|�2������Z��$^5��1��]�zl��jn�vgɿ{{�_��M�C30j]�l+w�zw���6��`�H�k�Hػjp�p�g���׼��QOt!��kk�-D,}p�l�Í$^��rsw�<!��fԻ��/h\��|}����o���cz�` n�'���i�qF���f��6���OQ����s����y(�'j�������p�ʫԝ���PL��j���Y�J^$��8��r���2�)	����E�Y�,8�u��F��N�lP]�dn��Sq�ɻ��Й��$4���d}of��~~���OCS~��o�ɡ���{�VK%2��37�<��r�=���8$wv`@ �3��O��h�h(Q:3'vE��c�'�$kjc�A �N�B�S�T�<O��ոpH$����g�?$1��8������û9~�g��+o)����4�����'��zd�%��]ߗ{p=Ռ
��d$�A�!��%H�ױ�N�M�V�^f����I>;U1^/��`�hB����߫w\9aQ�GM�M׎yy�J�]�PC%u�{i�GV��b`��ʑW�Ӹ_<��ҷt��(=��4����s���F�C�ug_ Wn	�و"�a�ٌ�`����u��|G� ^��{��;@ڗ�	]���'Wh�3���̘&��~�8V2���`��ylA �x�{����k��:"�R��Oy�q�<{�N�Z���Nk�G��n�/t|�<�o�v�qi�^�x�?��.���m�>�����B�ѳJ�-�w=�iRf����뽔C!�ݤ<=w6����=/�g[W<�w�y�I�R8ox���%1��};�Op���ڢ�&��w<=�E-A�{B�gވ���^�n�۞XƸQCs�P�y˲�����Hg���e]�ތ�f�N)�����|]�(wv2r�}�s�޸��a� ��	r���E�f�bV:�Y-�������c;�g��O'��.��nu��;x�v�욇�#����R]�L�e�ꟻ`��񬁾HǾ}�Wpn&R�kre��݉:��	m�Ӻ����Fif�oc��<npn����4�牦���>�L��� 2��x=����mny�y����8�rOz)_y���:���Ib�����}�Γ|��8gh�Q�wt��V(�DV�R�F�c�q���Ù��~Uo9�S�?,�s�;ܼv�����}�_M��������OOctzxM��W�p�O`��9	�޹Ӹe���w�r<:9q&nK����0��V�:���}���ӓ�óz�W�����Of���}hs��{��=��Y����X��sܫC�y��,��e��]Z��bD�F��2oJӡm �S�[ v����hѺ�ל�h}�<�<Wz�=�x�3�/���A5������ �Z{�KC	��V%���ߧ0�;^��=��b�g_Y�_(k����q�x�&T�ND�3pc s2F �XK���K.a-GQ
����'"ʤ�W��7rcw͸�?.��T�#��@�M4����o�5��G|�h�Y��er�&�a5����bA��sf����dזf�-���H���c�RLD����r��Sɵa	>)<>&�䙒(Y"�G8�3+L�
ƭK�4��ɭ�FH��a�[����h���q�G*LI9�SÇ�'=���dR"�m�tV#�ǉ�UǑrY�5��y'��*����_ml�$F	���d���M�U��#�j��X�LPUDN��%��Qّ�
a���\��"l�v��#�"m#�"%�������G�e��"�X=���TEr�rʅʖ�$"��8�(�T��m�d�w��<��s�!N:]Â���&."!��[�L�Ym�d���H(��.0��v�9��9UEd����q_m�T蔦���$qWR`�(�!�䌇�l"Ă�e��qr"E��b(���6HA�pU���'�ۻ?�:~>4�"r3��1�DD�H5��� ��h�"2r��S��b�E�v#����AF0]�nKaT�0D<���TEPU\�E�OR8���Q�Z���q�$�d���qON����a�10�L84��}��s�r�ej����G������Y������<(��p��1�k}����N~@�Ls"{��nxg�A̎28n{���#�(A��Q�￼�̿�.���˦;`
 
>G�"}O�a�(����!b�;��b����G�6߹���S=6��Ha��۫�-7��������g�G0�2�w�x���q8s��|�1̈ÄD￹���|H�:"�����/�Ģ�8� -� �l�̛O�v�����iL�8���v)?�p�g��#��#/��'<s"̘�p��鿹����"<_D�|,�C��fJv���z�-!;T�z�xx�xD܉��D�8?�)?$Ҳ���y������8A!���E�O_|��'���|�x�(�\L������xdL�� Lp�~(����R���1�=\�L���!���D��_ϟ7����f���b��������0\�L?��uy��`��\O��@�Ғ�`��\xY|>^ rv��ዘ({�dC=�����28%�� �.\��G���!�-���K���D#����?����L#�9��?�۪D�ja1�a!���<=M����z���iKº����%-r�Wu��q��\���	ă����NŒ��{OT:)s^_-�slL��ɛAD���G�>�>'����<ዘ)���g�M���[}0�8�ߞ{x׆jl�j�>9���W�8g������fz9�y����\������CLC��y�q��}��T�<'�^�Pu�\� �U�N�����uq^����tq�bBv���}�cV�a�7���?|�9��1�$�d�>���0L" |#{�Ǆ'�#�
WU�� c�'=��p��<C�T(�����ÂdpLdۻ$�C�x�=@�":���O��x�5D5��^�F�DzA�DX>�+�LH�L>�7���V&��u8�+��(x1��5��}�+xb�z T��}8GΕ&ֲ��L/���s��bALEO����������1�b<���%�{��-SY�χ��̎~���.Þ9\�Ow��C��0����>�����f�����Qc�]�r�֊�?b�c�C������n�4�Á��#�������z8ɈȜ���pā�O�խ�擾����DG���È|������T����l�ǦD�G��/��#�1῿�s���G�%��t���F��G�>3���`��������&�L#�����$H�";gR���w�1r�UץO߯{���?ݓ�y���M&��ޱ�~%J���~�',��6xN�A!��ޛ߮�GW�r^[~���X�x��IIt��ud�s��_��v�d�B��fu�`�o^�5��s�ݗ�`��A����M�A&ۀY=n� �l�(�$�9�X�\��2*zX�5>��n1у��Τv�oX�gl6�m�E�(6��xuњ|�(�Дr�lf�!��D��î{�n���x���[p�[rW��ƽn=pa�g]�N��xڝ���~g�]u�L�����0��	p)k`&:x�G���Ki�U��kˮ.�<�9�Of9j�9>���޶�?îer�D#��߯�����x���2<H��G�L��(�#�_W3�GR<���s<����VN��1r霹g�#>]qQ���oxTt*��iO����@�VWZ�>>>;y��Sjmy����ǟbO���>� m��{��sNO���#��EO;�N�0p�g��#��"�u $���p !7���3����
	\	�{�y�;V��T����1��Hu���	��P>�b����0<I�8!���,|�Sm������Ó�iL�x�} �yL}�9"p"}��f�s#�#�7���y�&x8D��4J9���5s��q�M����8� H>G��Ք��=�-��!�9vb�h�
�G��#�J>���	���L��U��������2���D���08�sț���)����5
&w�O��|6�[��HC���>D��.6#�u�pM�16�]�q��a�XB�6�e�� ]�����s�M��6�����§�OLÎg��s�}���1s�D<Ĩg��wTØQ����I���"Wr�='����̌L��~�)��D�����>?]��m����������bp��^^���č�
,[t��Y�ƤY����0e^9ˏoO,��諰9��U������Y�oG�k�x���|�WvK|�3h�����?l���L��_\+�<���xb��p�̃��'ޏ  |��m=m4��rrftO	z<�����벛����c��}�a��HQ��~�����	��T�����{w������e>2�6{��\�7��ϟcͫ�u��3����ÂdB���;����K��w��>�$O.���;���<,���z�>y1���g�)��z�@@k�&߽�Ã�0��<��+�5�[ؼN����&��E�\��<?T����?}\��%>�8�o۫�u����F��w�z�$S]"��(���y{r+ǅ��Yu�Z���||y�6Z�` 1˩{�D���r�f�h'x�������.�Ev�k����AGeX���
e�6�)�Ό��|�;�Ś��=s�~����0�f���߷W��x�F��^|>ƃ�����S߼���� 9�0������L�����n}�a&ͷ�0P���`|$�Ȁ���әL���G�^^c�+��!�?���S10�s�y!��W��^�%��ʴ�>��y�*z8'~\�礗f�[}0�>�>>���\�p��ˉ�B�~��{M$��ov/��K�dÜ��1�9T���vlKÐ'&�ˮ���N'ٵDL߽��{p����}G1~7o�ꈙr^""����S�`x���ݡ>|I�Pw��%*��W��xz�1LC�`��5��cU���5��$H �K�����Hv?J�I�^�}�g�)GD-�}	�q��uU��b�^g�"�]m�!��	d,�"R3�%��=y�^]�#k�[��A`���ݓ攘�_<~�z���~I=�O��m�3kF�$�^ɴ�l��c�x5�3!�. �CoI���Kﭚ�2L&8'��I%x�2ޛ	2KÔ�O�R��:O6�D�hQ�x�&H�R�Hw�Z�`��UD=�F	X��n���f"�\4o���zI$�_�I2�C�2�&��r�,�uy��=����s�l6������>_�4lc0�Έ2��C��krؚ�0�}�%]�&	&A�ޘ>3��EO0��S:w,Y�n������&YeG���	dSԩ!�H�ɂe$���Y,��2 (u~��g�&{Ү�<���+�X�4{G=�ͻ�g4Ū�\ζ���^��γ�1se����TYd�W�^�V��1� s�I,��3)<�d�b�X;�u2��t�})yHf��Ø���זn3i�������K�!��)%���!�;��D�vo3`�	��.�dC�5��8U�%-��vB�ݵ�cw/(���MϿ~��̹�v	y�K�^��Pȑ��2(;	ywD�0��UR��2��-�q�1� �_���k�}�ϰ���:�A 5��u��2�/����z�����NLD��2���2��:!itJ9��CTl����˃���vE��!�2��'�\D$Ipo8�{6��'ӡ0dX�gL�I��G�Y`�ؗ����:я�(�~XuZ���F�d�H�Q�!$�J�`D,������
�(k���?pd=z�I��g���l ��m�0�C�]|�}���Y�E�`�O��%�DH7�!H-�2��{L�#f�͜E�]��5�p�h�A����?E�l��������h۾רl�vj�� ��	�"�_2sE��b[���
��rc_ٙ�,���V��\֣KD.��m^�'�����d��]m�?��|���b�Xj��^'����UA��&�1vd-pA�ț<$�#�d��sM��x˥,��L�1��b6�E�P��b��X2�5�i;Oe����s]\��3VGfm�\YZ 4�a*��ʬq,�j��A�Z�*���5\���֮����S�q+��̕	���59a�	���ͦ�-M)� ˁ�=��'�%n�s�u��P��C��3���gD��o&$$�^�k�h��O��'�Ivt�$%�U��b�^g�"���%��Ӹ���J�e^�ؠ���If�&K{^L�(�O<9Bf�:�E>fCZJ�5��!�2L**�;�H��H/,�y94/%y�g�ZDI۽����@���	�y$��,��Yye��f�"�}8���u+��mXZ�w���A/t[���\8;�}س%�^3�މ~l�����!��h$^�Ò �_I�e��@����>��*:t���K�[9J�)cl��j�w�Kˇ��	!m}�f�l��h�iIUv߰׮sO#`�p�Rٶ�[���q�HѪy��5�<qw�e�4v��m���y�6�pYy �^Yz�*W�3y�#����N�c�۝��[\92��̸�"R��`dvE�3��.�ע�>ګcT�j����ޭ�̯H�`0 k���9��Mpv�_i�oj9��4�Zce03���ͬS��DH�&hf`�Mђ�TZ�B��� Mm8�H$�Y}fBK��P���T^	S#�����p�}3��gA�^g�"��ש��!��N7D�I%�@lق���JFx�	 �ױ&�4�k_�KHIr���`r3$�EziF�
PP��'c��!'�z���d��'eH�k�y�V��y���2A?tY�+�a�c��f�"���e7J2�Evl�6�U�h���ra��)�2C&ߥI����X�v��6'�Nm!�4��d�e��8�;�i��s庴��r3&Π�YK��\
������ߜ�	8u��lS��Nf�&�m�Hd��Hw�t����
�PA�y)اB���,��>�(��cg�BO��Fg.�4��.���@w�Y��x���)���$��*BT��t��������,�N�F�!bxp(�.�9g����T`d�H%y� K��%��a�����t]� �=��b������z�ŭӸ��Or�������k��:a�Ir��=O��9Ij?��_{'\E׆�޴����+nl� %��1�v8�"YH�Ҝ�gA�^g��%��z��y�y[��ڧ�8:�&̺��=!�($�vBD���$�n��9���+|h$�9�T���i*Y�X�ٙ&�:G��f'���N������I���I
�z� �B*��@,PIywdQ�\-Ō��������)7a��ԛ(�M.F:Ȏ��N��t/8S���p��۝j�w�~���U��q؞��N	��̹��	$�K�"O����+#'��b�zv8F���In�]���3��# p�ٓ��RUq&W�����;G2ba�-K�$/2@	$��P��B��|D�U�����|���>�Iy� ����úf�Tۘ����bL��]4V����Ӱ	%��4�S�=����|	��O%6M��eds\�vW55���KĽc��H%5�	����%8H9���ژ�z�އI��k�*�d1ɖ��3��ջ����h~���$Hf�K��ߪ�S�Z�]��1%i�c������a2})��t��b2	w�rH8iS!neV�仺Ky�a7y���B��}�y'����Pv���33��d�j@K�$��Ę&RO��&BN2pu�{��P]�:�:�*F� H���M�=�u�VS���N��ƕ�\ޠ}�c���*3ν�:��S�tH%y�3�)$^��>2�YX_��><�zq6���O�/�"�c�I�^[�e�y�7����W�2�Id�
mL�/۴��a �(n�I�H���g� ���f+K�!593�W�`G]$�`D&0��ZK����$�1�~��HN�Z���U���d��ȓ�QI&��X���Aс�;�t�B�=8�z�A�m����Uz��I$�a�B�@$���I"|Q)m��IC\����� ��m%����
-������_��ۄ�%ysf��1��exʕ�ߵze"W��bL�4�/nt!��3�� N�"����s�0�E�^2^�X�g��aI���󏏢�<�f'��O�<�p��ϴڻ��mX;�">gs�ݺ�X��e��	��*�����8f���D_��d�n�o���=�yvLC�P�6����<7�1`���A��(a��[�3��s^/x1N�{F=��; g� �%>^�^w�zo��m��g�or��uΏ���}�ں�s�p�)P�P����G,^+�{�<��4/nR(��s�q�6Fĭ��=��h��ݑ]S��n������q|�����z�=�o���U�=>~{�O���Ɵh�ޔ%����(�uû�ܹ�q���ؿV|���,�ڼ}7���wn�Kp:�t/^�� �� �n�~�&�֡�n��O�hy�!-[&Q��V�U�4	1�}�.����Bs\�z[Õߝ6ٸ�(����+6<nģ�qXI~�}��Q�K���T�FU>1kɼ��vJ�jG|��<b�w���C��]3��פ��U��}#ޯ�f�g��(#�pH���'�qΎc��yu>S�՞���a�ɝKv����h\��+�w����`���k���������z�3�k;��+�胐"$�H�K��o��q��Z���^�f�ď`O�Onkz���Pq������I�AE1]��n�g���=��;�U\�}�D�����.��Ƚ�8.r���p��oM��g.�����R%#�QdL�d1��.��ϴ(�K�'���|����G�e�(@�)�yL����
d��3!��H�W����?��Iiǭ��3��R�Fʬ}�8qJr�l��[$���ϳ�^3��
�(����%�I,̠�#�X*Kh��5	���1I#���l��	
p��� �8��z�-������"�B�5%��Zl&ȺH�Ka6�E! EB��H��dsfC��^�
iӦ��S��ߋ/�v�*+6Wd\ԮeH����MI�,�DBI�����*E$�1qē"��^��8t��Q�?BUgU%��L�
+;M]fAq$�����%$��$AϒY���J��$�Ȋ(�DS�)�����̣+�L���8#�Er�@��D�&���qϦB�d,��E��O��؊l�$��Q���(V�bOR�����@�Z=�d u&b�!72���Y��$�����K��\�\�[��$P��f8��*�lFv��&r�L�DŐ ��(��)'�U������ɉ6��4(�d��6�NH"*�<��Q�L*Wf+��NB�kq�$H�T��")��H�G�||COO�sUGz�)�^��Wd[1Ȋb��Sd��]�I�fG���"�8�Y$�8�qA+$�R&����pr�qJ8�[:��7�[N3b�`w�ɤ�nC��7=�Ƌr��@�v՗�u�ƟP��%p��N�<�������SYic�i��J+�ֹl��B�֭v=s�#�<\�-��]�\`N�G;v}��U-���ۖ�w%˸�#�x�%��m���pJR���Gt�ݽh��:[�-���۳L�s:��xZ��y��8���2F�ÅW�����.�eά5���ww]==�f�kcC�C��OV��;�w����K��"�F2MJU�E��ˍ-҆v��.
�'L����݊�m��!�؂\�����GL�]M�u��|[�c���� ��Ŏלs��sջk��LhB�Dc�4C6+n�<��-��q\���=��Z1�d�ۺN�)����]�='SVƻ`��+K�!�G#�t\���^:�Ǖ�+���-�ax��g�#�8��s�b�7.�5�$%��˲E��	z�ܜf�s��6�	�Ku��������8��ϣ����k&�\��Qd޳�lvF�d;m�v6�y���*�یV[m�\��z�;J�2�=O�:�ֺ�3N��1�`��%�K� m�p�{vtV��9���N��/1O��63gq��^�'
Tv�����:-��0�WM�U�bQ�n8���m���j�eDL�:��Z�>��e�5=�_G7)����۶�+�u��Mc�\O�Ap��)����Y8N�]M���7A��V����vZ��w.��n��V�nr��by��({v� -�6a���f�hbY�3�&�P�l��m�VK�!��<=�պL�m/7lv<&b�[A����M[,I��IL��U��dѤ0[/,pGM��c5��v��GB��Ըpa �b�AF$턥l���j��뒵ʝ�og�ƫ��gb�lX77<��3<�=v�asT��o��P��g���EF2��P�H�@<<,���7uɶ^�*�`f�u[��b��[���\V�a[���h������Zj�g9�e\(up�q�V7��$.�0VP�8�j�jm5��97���ٓ��ۍ�S&���u����i۸��cs�ڸ�[�<Be��Zݢ��}m6���ґ��X*��5[���N,�Zn�we6펞?:9�򛵠ڝ�j�0LQx�`XsE�-!F.������e���p�����-a���;��m�78�;�����ʖ�RO��伒@$���0L�����ɇ7ls��>2O۱&@IB�36�QvfL�l���	���i�ݵ�LH���H�Q��&��!���b�J��C����`�r�A��n�6"�,����Zd��J��;��&��LX���vzڗ���fב&|���p�
V֓��.�LꚒ~jށ�ѬC�چ�9�O��I���I1��I��b���_���wLI���p���;�iK��@�^D��R�ӷg217�=�>J����Z�{��K˹����"!�`�yG]~���h:`r�(- �f���j�j��.<���n .�Y~}��;�.�s��k���;��'��n!��fU�����h��6f�v�ѝd$���^�0*!�ٲuػ:��=��.���I&�ۼ�e7*���>Ě��_(�:愞۠�k7����/��F�
�?!R�_�u{��yil�]����7ܢ����l&��{�"e� ��X��{,f�
�����j	���6�N�p����[ę5��d�HE�2g4�Ol�f��l��$��ʚ��Wo�\Ů���\qPfd�����*Y���J@��K(�A��wwbfi\O<�;��?t%�Y5�`���V���x�'�F�>�O�}QVс�CS��ӄ���	�XoZLA�1tgV�~j�$�	p`��!'�[���!f�u��^A$S�)T:S�2w�q�7uU�_����ix��p�`6�\;w&���qɽ�FXV3��z)�"�$Yı���ݖ�\���B^I��vCJ�����)@z�o�Y�Cl������"�	%�1�e _������'R[z�.�7�%���I82��`���K�^�J�A&��)$��,�1�V�y��ԏ�28�|�����m�K������I���L��O{��nC��Y$�ڼL�o[�o�o1���x���q��h�s���_I8�V�u��'/��w"�Z���h���K�+��%�n�2A��jY0�"陙�yPS�*�����g涤�I�j$���$��L��I.������t��FW�
EȐg_��I-����g�K���<�!>-��M2<ͺr�^�ۉ�e�X�t���$�D ���ҒH���4Л{�c��ĳ&�	��C�F5��p���K�mt�
��ͬ���-�RL��0v�L�1t�w]�#�|���A&՛��$����/(��%��c��W�30~l�i�Hq�Υ�]×�X�]W}	a�2n^��,1Y���fH@�c���&��:���+{����;;)x���I��X�M�fe$����H$|w���B�Q�J�֋�m쑎���$�Avd◳I��Z��3���ϙ��f�"&"�62�!wq�u�����aw�+�8fd��@�.%�$��GH�������w�P��tn��=���!U��������^����Ǻ1e��WʧnyusA�«��$��}�	�)k� ~<A>׉9�����*� ����L;ȗb���V�@�Gě�r'�D�]WpK~��J��2��%x-�%o^�ӿM�~����K���md�k�e�؈сkծb!D�L�gV*�{��c��V���w���e$�[��"RD!�;e$m����P�`zzf$����^~�	3h�_��I;��z�];q>PKZ�aV�NPg��\��Hu�>dJMӲ��E$�+�QX���� ��
qc2g,�;�V�!u㈄��I_O@��^I��p�ڄB�f�),0,sa�B+�%�;"e,1�Ib̝���'U�9�2Td��	 ��8�	.�2Uu2�BI$y���T:�oOMF�/��}���+]�3�`�g�&6:3�RI!���&RWїy�kgu$6�zI ��$A$�:����gZ�f�5D�s�{yn�W��p�F�ˡ�h�vZA�"��z�SF���n��v�էk������v���{h�q�`�@ב�F�1��f�ԛ���pG1�LG�G<7��Yn��%e��2p�t���{X��.��,uh����v�u�o)͵m��G>��T̀��3VI�Y�7"��(��#P5n��GW&�E���0��!�ݹI�o5SV5�Q0�6��m�,E�m��K���k�š1�^��ׇCa��&�����ύvΖ9���{I­4�V6gb��Wb��.��<�t�-ϗ��j7=��Z�l̬j���$9�����7��a����Ծ�S��
1'r"/��D�����X���i������U��&W���k����gtj�'7�>�I&��b��ͣ��P���I��4�� �;�����Q�w:;�&�eQL�1t�wib[�`E��t��H��A(ֱR:�$��rD�E����əq���,���'t�U�p'�I���� �D�0�$@o&A$6[:X�K�V���z�p�"f� H�����ɋ�;:E�R�[r�#!-�qc��ɦ�j�aj�N��М32U�-!$��w8�A�Rf�����C�왚���j���-E�d�%���z�(ڈݎon ⒝t�@G���⇹��a��ꞁ�����>&{�?�vہ���N�2&QI,v얕� :��2a��'��[X[}! ��뜇�qQg���Y9tE�J�-�9|�4���0��|���7|sNg@UN��|px�c5FλdY�������-ݣX0G~tw׎vvst�;�ze��L�5�9�������9�|�$�����e�$�U�@���q�"ݹ��a��\��\�1T��~���zo-���4렀D����8l�t˶lI�����ײ���N��G��/��$3�K���X��˃��27�ZX)�ULK�Di�/"�>A%��]#*�kLX�G�%��~�jIr`h�F�d��:83���	/%偯����ٮky�W��-Y,M�fI��8����7ü3��&<���%CG-H��eu�e����M��MF�`a��5�6�p5�����(ݜ���<���|I
��	$��ղ&B]{JgZ��ђ��2�ɷ`9�)wt���=��.��J�N�;�L�t]D�D[%��+�}#���I�%!���=pˊh��'�u��fc��S���cb�Q�&p2�Y�"|�	6ɬ�z��:����ٷ�,�w�Q���\]s�h�Â�:�Xk���xp�|��ڷ�g���v9���0�O8s��������ۗ�}9�?�g��b9�9�iY��,�fQ�Ƿ���^�uԗ�Gݝ!O�N���[�-�;���坑���-�V�/)���W�� �\��B^Ic3vWHBd2BCy�m��u{0f���O�;$�fBDM*L�_��E3��[rc��,�e�ͱ,���؍�ںa�̒ʈ $���͞�"QA�3~~�>G}u^����ߞI��D�p�l�Q)mi�ڷq��n(�0����l�fi�8h��������l���j�D{C0d�Ms�"D30Idk��	�~]y'sv����B$��9r�1�}�8�-KI�����<Ia]��X���c��$%gOH!$(1���lZ�a�' ��Ud�	9a�$��_th�	�npZ8�]�Å�|��e$�X���A/LTA��� ���$��vmH�aW�/d�D�!x����f:��p���
s�5��A�W�~��%J�D�љ�)/����mk�O�3^_���z�yw5� ���4�:M����=�O��������}�H���.�k-Zez,C��&^q�k����}߳�λ�cz#�A�Vb���#0Y��y�|3�z���R
A�8cXwE�3�vF.�|��gʾ��K͚�):�Υ�8"���d��K��&R^H�e��"�澘�㧯?_{�hB��ⴳE"�a0In�N��/�׵�f�sd�)4���~��Ry#1G7"[3�Iɉ��x���H��@�	-#*�Q/��"��j�"Q���t�ę�Hh��<5wt��ػ]W"Y���-xS��cktXi>)*�ǃ)$�_8���5=�E�{\��zKг)���d.���	M�8�^$�`����I��i�0[5׳BD��<	/$���!6�8��Å�y�����n��ה��ue��H$���L���In��$���iՈ�y��ԪLT[�,�O\I�N(0�L�j>.v@�R���I$�|��&���ne�L���%!�&�\G�PL�� 6�>����5�9ֳ�Dė�q�,��/ż�(ٚ�yt�O��/;~�4�p���.�u�r�c�"
i	'��P�*�57!M�����}��������oܓ���̈����􇦤�+5d��LL�0133=9��6�͒V��3���t�	:ɲ�7[l����8��/N�U��mҔ]�v�������e7`3���CX\Օˡ1hMv�&4YkqJ�Xe�T�13�2��N�CƤ����]vn6t2�ئ1=vN�:�Ӯ^�q�N�^v^b=5kqrqV�7U�ǒn�6��2�]jCI��ҜvR��:���D����c�;=\�]�񧳈��ts�nt]�=���zC�]�m-â����f��d�����y���'ۚ�%�]�:�BP�u��ϋ*!�j��f�L��GoD$�a�x���2
k�a��]�_��1n�ݿ�vw�,$J �P��!�[�Z�W�	{���m��ᱬ�FBH����394*�M��D���zCJ	 ��ʘ�toc��"AI#w��I��D�(|L�A��p�1����y��izނ�3-$˧H�J���	$��tO��i'5L�Q=pl�-�3�v���G�j��W?�X�4��9I����oTq��{&x�&�z�"|�^\��B�5iN,�賳�t��-0�n4�al�v�jlA�,5��X���Ͻ�`s�Y$��c���>9�9-(-�y�z$�TdN����ϑ-�qVԝÉ�
�����ú)�9wdj�}1A"㙶9%<M����x�l���Hs�3E����������B�带j[w��<7��q'`�r�4���߷~o��Y�zT�e��Qf�f��FiVb'�^�������nx�2&���&������+E�7�#a"/&,t�giS��A
�	k�<HI$L�E���z�H$}��j�L���<d��PCF"��ٜ�ze�6a�K=B��I ���&}��~d`$��R�ئd����yꦠA7^$���T% �#���g.�:Lj�[
�%��D�k���Z�fݱ�:�Gz�$���ګ�$��n��H^I$���[�� *_
�#�C3}�5Z �-��<b��;��{��Ld덞)�<��-0Y�~O���m���{}���/D�ᙖB݆2A//wd�m�kث^2u�0��O<j�Tż��!%�DJ��1,QNҥOl�$����W5M��D!c�In�햔�32���pa"�����4AK���s�JU��a�$Ŝ��5ꠞ�T˯ �	v눌���Y�{����VN)H��u��I��9��{���a�w��s}�)��;y������w۞;�e�q������������	�<4�?{C Qr_��K~ԇ�]66�9����;{4{YK��F�Ks��=��=�s�e�r-�!�<� }A�����������l�4�:�.��{�X���s}��ʳ�y�<	�s�NG�(v��㚖����}���3��S���R��&xɈ�:�y��zI�]��/�$ڃot�y\H�<�x` �����E�
��^���A�!��ʱl��+�o��c{N�W���m�'F+��<Y�gc�{9H��[���g6p~쮏�]� �=��pW'yw�F��y�Ǿ�k���OM�&����S;='s;yTӽ�HV2'Y3`�|���V�Bp##�;`]}3�\�;��v>��2�;<��x;�jԊ[՟���}�ugd�]7[n���ؕp��T�=��g�:�����jF�����g(�D.� N�|��/����;5o#=��|Dѹ���k<[2�z�<3�g�E�ޣS�X{8�ԝ~,6�i�.�K���;��]}p�Ho���X�{=��~,����į!�n׽u�{�
������qW&,x;֭Xc�\x����[��o{&9��Wb��5n��N�,�0�x�.yb���k�?@����b��Mrf{o�E�6'b����6]4O�>r(�����s����>�<c����hO�U�39&g�m3������X9��p�^�PKHd}�C��#^+;�E��}��૲8�dOK
�Vy3"
��M�Lu
��������\$%�O����!$\R2!H�MJ4TQE
��	&FH{"��������
i���y9"��p|y)Dq�"�'�ATEl&
8$q�\�LE�J�!r��:i��.�8#���#��{2�6��	Q�+�qq�UI�DD�Q;!��/��Jzp�n��H
0��Ȩ��g�~J�|��3Ă.��&8�EX98�UNBaD�H�>)����.((�����೛KEB"�\�`SfV�5&#d�6c2(��k$ ���>,܏YfLDE���.�_�,�Lu"G� ���b���TdGQ~>!N>44u�$D^�r�v�.!�wK���'%V<.�O��\�/fC�֣��l�!,ȯ�t�9�
V�p��Od�	�U1qV$}`�'��T���*���y�䀖f�U�m�TR�)��*Y0�A7v��$�<n3Fe�t�9߷S=����$f(�C2�0Lж��0��>�}?�ĐH������$H��^�T���:,��%�%�Ս���9�̟��%bėޟVNp�T=wP�2A$���x�q�F�O$f�6A�k�SRI�Ŕ����vg&ştˉ����%��R��y�k��2�+BA�p��Ғ	 �r�L�l���W�y��9�Ǒ��m������F�- `��J�͎.��[�c���G�W�m���hq-�r�äǎ�����$W��.f�Hs�ʙ�LI3�܇:���MK#2K���9����û����UIu7T�����̪��]
�łDЮ�p/Hj� 2n��S(���8��z��/xġA�	�"�)��y�L$'{�)+r�>�f�d�bm�$�K���91��ِ&x3�,��	A0�#wp�?�{���l���(32�D��+f�I2C����޷%#|�G#Y��L�A>[�s�-Ͷ��}0��&�%����f�G��xY�'7}�;�C���{�Z�9ݏ�-�#ᢙ�fA���C5T�I�	�wzv�o?/���`lєŏ�0tY��_����|e��_:ϡ��5�!=ϱe֓�c�D�I.��(S��CoKO��nMΗ�J_�_�C��^}��cch� ��"en��Ƿ(��mj%���]��ޒ��{��S���qВGǮ:'�|�H$�ۺX���8N�N��o)���t+��d�jxie`�r�ä��\*�:402Gll���t��ْ�� �X�t�	��+]�$�BTe��ns�8��d%��)��Yû���ϒM�th3�,N��t�A-��v��U0 Z>'Μ��	&澖�����p��$���T���B^��H%���W�A����R	%ݐ	�����P��<ٶ~�O�2&|������vF�ֲ%�d2^I%ۮ"���hy{g�Y��LUH�^I&�ǃ>I����C������"�Y �ld�-�6E�n(�Z�5]���
��I�
���k�k�EN�Fe�S���ECS�`�وa ��$�d�9�����ڒ��?Ø#�&e6Uf(�0L�� a�w��f�Xn���e���l��.g(�V��.�2g�c���C��-���{��n
c������٭O`y(��0��H�]GG��XYt�J�����\Js�@���p)��5��+��6.q���޻8��X�\��+Ҳoj�nѰm�v�L��N
K���k�Ȩ�[
��DA\K]a�G!vճKm$�Pū��<j]�� [`�uGq<�{N�j���ɵ�B��
�0۟���LC|E���|^�c��)/$�w^	&@I{{ ��ګ[�zF�0�l���E�ns�����
��S�B�˪�@�����"�Ñ7}���PL�&�׃)pI�>@�B����rd�s�/ϗ
�YH!��p왂�
6��BI"k����I$�w�~ǰ]l�]֐l�	&��)��@q ���bg	�ܕ�z�K�z#���d�*���/&�ׂg�$���BI$�t�.�֌�%e�d�\�eyh%���وI;B�)΀�	WFD�g��n�.�3��	�v���^[�� �C�lS����۟�u1�3Xu�)�8H�x�GqA �v_Y{PGYƗM1��X*hU�~��C���vF{�D�̤�In�'Ę�tt���^Jcٙ���lI��"����҆.�X�m������?������N�[D%3qX^b^gr��2D����g;3c%�ȗ/Oq���qn*�-�6��j���^ti�֞м�17��:��*ǃ�$	.�������}�A0���|�]Csۑ�?� ��%��3I3Bf�"�&�3��y�$ɒL�g�^�&RAs��&QAy[�֗��g�p٦BI�^%�w)±f�\_�$�\��"@^K�I���ww��@f'�7l�`d�"���"R��*4-F�)�wɍR��Ȩ���U���u��sʰ��E�wnXFB���� �A*�3繗�P=��|���䰃I��j�k����i��&�p�I����$3�>1�
���ʵ�D-�k];���J�Q:��Cd50I%:�$#V-��n�ֺHuT&<�����"}(��ݑ>2��v�v	8~φzK��a��v5X��3Ҏ)e�Z�`n,������]��2(�<�;x�v�bi�z�I*�ȓ$��n�'��O�Ȭؘ��n�6��!�6rD�C;,���3p�����V�2�JUn�e���?J��N�&	%�7=$4t3/?oD�ey_�����&SO�l츈H�2���:t(ܨ�C�kb�b$�Hpfy�-�P#L�*�oυc�M
���T��m�=1jV�P����4o'!Fث7����;NYu=$a�[�����+;����Ug D��<߲�X6E�e�҇�OM(̔�#1Fa�3*3=������]:�{|���<�^(k3?G�&BHV�%�w,�S�89�,�w9=j�^3�]{q@�  Ǘ�}���8w/�z{��g�tFڃa$��O�z��`��p��D��v�e$�0K7�9o�sӃr�益y��$��o7�{bL���� @�'��_oϝo>W��w
�]�SVS�;vQ����GPY��r��i�I�qm������i���^w���l|ex$���3�	��T�9�BUm5R�g�L	bKx?nę	'1ҙ�8b��
�jU���,�1�S��E�)$n�x$O�'�@����;e�[S��������3`���x�>�1قH%� 0�3 ��Znj�t;G��5�$�j���'�偘��$�i�Hc�o0wd,�z['_�"��J�Ě�$$��.�p���	/.��7��Jw�ͽO\��]
<����U[�.��`Tڂ$I�T�gТ�)�Ln4�e^�Y��dxƦ��Cx~�����(�1u~8�}�}C��̓�
�C4Fa�3�P�$w�z�^|�����|/�%#��%��2T*��j�I�>~"A�~א��s��r���%��K�r������=dJٰi�8lTE3�I�N����e&v���-��伻ˣ7nŨ�̉�A�.��1oD�<N�S���*�sF�<�I�3f��^^]�bR��[�ҧ�Ff�绉2X��>8s>kӔ�çm�_7�������H�,�n��g����fjfd���@I{C7�N>��/&u'����X�����`fa���t�8grv�D��l��It[��JH�Ue�sc�ݣq��Iyvd�+	���.��0f�1&��f�ӥUA\O<��Iz���&�1�
C#��q$A@$�ط�Ϝ33��In]wg^*Wb]�ČM8c?���lbX�h�����G���/��4��\����Цd#bBD��y�^4��Iy�z$�I��%a֔��C�&�m�K��ޘZ���c,������[��7�;�X/{�٥{P�_o���I��eO.���
/���ޝ:�]�ww�7]�����ĶS2�h�Y�c�f"�������M�$��wd�p�˰5��]�+sϬ<���������gqB[�9��a*�v!p��:�(k��s;sS�ȸ�l�m��{5��<fǑ�y�wl�F�,3�ƙ!�K��u�y��vm��]�.��Y�!N�(��e�vU:j�6g^k44��%�q�y�ln�`춺�8���֫t rX�N�l�,�0�U��f}�d�*�:�z�=m�mt��x��u���M��gr3���%�:f]�����! ��S�*P	 �lމ2��ܷ��m~�+}2}��D)��.v�<a� ���Pi��7�*�Iy/c�E�X]����a��p�d��C�#L�H$���I$��qp�mȸJ��.���w����lzA�%�9��Iy(�~��8e�y�hI$��/�H��J�z$�3!�YZ��3��J1��d�d�m#nrh$�yۉ2����n�x2��,����0M��2<��$JYy�6�0v�.vɊy�C{�=Xh�"=F�Y���0�W�;����30ёB�y"P[�˽�i�FKs�;�8�	A��eeڶ[��$��t���U���V��I�k��Ⱥd����Z�����������H2�^I&�׈̗f]��ȏ�υ-�+�y��d�	ln�	/g`	��2�U�P�Bk������B[7�A��F���͆͊����/!��wݏoz�^̸��M����{��I�^�;˯������a��À9�Y���@�R̪� �2�[x�	$��^�������"�ygP	<�;l_� �P2INK������;M��3^s��JJ.����]z"גK�u��>I��B!M�sn\N����5=�Ջc5�aÉ��>��" :@���@�	$�[��է�ن�.�귙R�V!��n��w!iR�vI'��"O�L�'��:r�޷,�w���	XO�Ă�	hU=�"�|�ng���Tǃ;�:g؅��{�m�Xݝ�f1��8i�k�XCiu6�0O��轂�0v�+�bۜ�M���zĳ.dY��@��eo��'6dN�������ǎ��}N�\$���~�ř�:~e�I��gS����!�I$��@H���&QIT<n�̪;�%�X��K�a#a�:fR'�MD�Q)&��d��m��F�[�)if4��tB�O��sDe��|.츲u衏���>��(|W�ӟ6%��wH=e�x�d�
Qo9��P���L�B|=�����4�j�Vj�j��x�uR��H+΁Iy�}�$JBF,@�%9t�t�T�\���3�x9P���m�q t��[;�&B�^K]_C},�/u,3%p"	�lӗ��	�w�VL��`2JKgD�U��Z��c6\1��'��pvo^����̗���&B��W��6��6G8>w6��t�
v�b6l�XNܡ��gz���.1�В��^Y��b�,t]�r���̒Kg6$>).u}#����!�����X��GD�$X$::�3�����Ʊ�N���,�L�5���1�����͇�H�	!q{#������[U�JD VM�W �T�8�B�G=i3�,�ػ(i�]�Q&RK�k��c�I%QN�x�ïΨf���S�"�:˲<���:JXӦeLP��B{qG&��#�5d�N�xs�̴��H�s��e\1�*h�dd�ҧ����{���۹T}�K�l�Oa��{n�A���S�;L�UP�v��I}����{U	��4���
����*̪�S1Vd��3 � ؙ�)[�T����@�%�::f�]r��Pu�A,�q��3�+��/�N��L�宻a�ʃ8h�9Õ�����uN��
u��7J1� ֔�RŋI�	���)��]���8�j�O�y{�K]�6m��H���``�	d-ؗH$�H{��D�^�,�Z�7��hɑ>�|M�톐�8K�b���3��ۅ5���1� �7{!�]�vVTƙ%/%�v���J��@��#ׯ��'P`�4*���]{���Qff0|�_�?���8���p8�UF�D2t�lM�)	tslz�oK81��8b����M��׷;�7Os	7�/ �AJ;`>�ƕ6K=gL�X	.0��;�L�@��7I��x�nX��oFF�l Z7g�'{&= ���p��� 3qV��l����^\li{����Q^��ZuXi&Ցa�zm� :j�zn�(Ns�z��ϧz�_�8���lQ�k`6zF^���R�*�@Bj�ȸ@�j�����v*�D�5��:d-}o{!%�7��;��2���K�w�ov
����F�B��m��<�7==�g���}�Yy�������sM���D�5^Ҙ��+x�ծ6l��A�j
��7���`ߋ
|$��]�ea��G���.��,��w�1=s�vz�q�M����l�Y/{6E��j0��H~�O�ѫ{�=�NY�j܇x��^�ϭ�1�JV�{ß�J��]�y�}���w��nzJVM~���Ǟ=�;��u�䰐���X<L�`��[��(z�4�)c�ߗ�1�8�?N�'�����yɏ���|lp��՜����d��w1㻺{s���q[�f�f�A#��cZYz-'!tٻ�����5�wY��w�{9��Q���ym�Μ��^����j�����|���z�h`�<�oz��=�.�����z,�s���)�L����O@����9��W%u�>��+�Ѝ �}/�O��'��V{�c�c[�M��}�ڷ�oOy ��у��p7�XW�GN,��IaN��YO������P����������9����X[}n����_�{�qt3��v�������N,��̴��~�ݘ��K�,W��o�ծ�@�:���9���6y�w��R�i}���v��/��=��³d�^��9�ύ��36��6�;JEA����\PƚᎳ��L�͢�m�Ca~���T��Q�Z�$o��Q}(���E�6AAW��s9�Yf�-15���|�8�,�3����isl��LE1<H��*&YW�W#���$�� ɐsX���zS�����$�2�0�����.F�+���$s�bF5lPQo�R~x��$������o��b��!r1Y%b䰸�}	�`�b��DT�dٜH���'�8p�� ��A����2,����ܴ���9����K�ɩ�D�S�M8zNf�bq�`�j|吞3$fD�Q\ʇ�QqÒ�y h�)��N��N�.ͳ`���G\�1��
(���#�*!�)�d2�B����X����'�c��*Y�SY��OI���BR�<H��k�ClE$:iç8�$xHQŒ��EŊ&2"*�"���,HV�)��� ɬA	�8AKyz��#�;�-$8�bEq�,���8RM|c�y��ږ��u�v�n����a�{h������Bq-�c�۳kn�c6��`&7Wr��-%Żsn��y�)\񸡍�̏b�U����p]��g�躧��׍�7�s�<ttr�cM��������ch�9�G��B��0i�e��u�:�����+wlkd;'[$uƛ�"l�<�eƉ�֮���vh3��o������nnF�Yې��|��鑤�����g9���*@rB�ێ��q�k���nc�ja�Xng0���d�[c��[�!�\v���	,�� Χ�-`�:�c1��=����8��a��b�4gs�#5�������� ��qT]���]�[:΄3n:��������y�g�{\�!ᣯ:��Ύ�j������nB��N��v+Bj��Es8��l�n�{#�7��9���Q����4l=؞�Hu�Hsm�;��M���2�89���BH]!�7wa�����<�'��$�c�vq+�\Y�۪��k�^[r\��:�0dT���y.�:��j�8��&M�M`:��"LjY3��M�WE� �����ol�,\���ps� {�m��0�KN<n��mv$��d]�R�6]�h���9�l֚��xp��dc��6pZ��m�����������i���fܷ̑hL�)fu�50G\ֱ%h�8.l��t]���^�	i-(�G�`���j�x��TWY������qK��á�\yg��Iw��F����\ҁv��9�c�K	�
��Gg�O�==�hŝ���.�-�ƚ',In�vl��t�cu0�z[��;��d��v��n۪me�*���1�y.l�X7<�Fíw]����nw��v2Xa��y��ّl���#���B�,nu �(�A��)�k�6V����'PE$��ݮx.i����ݫ��f�<^�덑�j[���Q!hR�s���P��Ilun�}H=2�a�Y�3K1��s�L�iǞ��$�m�F϶m�:�t릌��h��ɋ�/�3y�	��E0\
�[��L��5��"b�����b��57e|.�� �Fގ"�י�n��u�x6���qqm&����I���9.�q6}7�&�iל�������p[��X�祭O��׎AWOnF6������l����Д/]��y,jwb��n��r9��	��5/R�(��X����1`�Bh����V6�=����˻~�OZ������Qs �X+�x�I��� ����*	P�k��E��� �@Z7�x�y˴��,�b��Gs�#_��u�F���"C/ ,$J�">���q����7{n�s����2,&��S9]�]�n�A �^8�O��G�c���f����';*�l�ǣ��;;"��O�S���\�[�-QZ%��]|7p#��Bn�Y����nQ �NG�׺�!l���ػ)��r�Eۏ�>3jv*xH��~D�>�Iȼ���-�}2Zm��3�K���0!�� �dHK�Og��s����!�^8y幘���n殩u��Ko����;�fc��`[W� �/]\<x��B�Ι>��޹)�ӆ�uZ�Ijy�#��&#��ZIv�9M�3�wY<�6�ͺiP��iL�)=��%�cb�Z��[3�^*��N�E�;B�I?x��8��{�aQk���ow�۷�vg�|�P�A��5T�D̨�UfT��{��ǧ�f{��|�
�}��g�5�|�ѻ��n;�F�ێ��)���՘��H-}�! �=�O���C�ބ�77�($#�ތ���	���&ck/�_[�*�ɱ&�K�
=�� ������$�7:Q�?+f획�}oy�e�v:vvE�҉��mL��@�ٰ�h��㓞bj��0�A/}{2d �=}/0o9�\^)BޱRue�L�.�k,�)�c �nQ/�B�X���Sf �}���N�k(ͮO�����oi�>8��$����r�f_q�j���u��K�B��&F�$��R�� ¼��	f�H�U}��#n��$�6`O� ��LB���)�&]-�{�����e��]0gt�5SumL��N�D�oj��(n�WƮF5�'��r�������ɗ|�5���]��91zmK'J��g��]=ٺ*Pk�#��+�㿵w�}5�2��#���f�f��E�K4�i'<��xz�:�|{����m�νw���vN	v�Λ���wP���t챾�U�����>#BZ�oT@�$ʞ���'�$�O�C=B�oj�%���"���];�����F@'��@��m��;Zx�����UW]�|z�\A>�;̄yGX7������-��SKmA)t����q��pݻXlDŸ��D����qwϟ��wLd��K��WL�	/;�d ����h*�.�K�ƆU���s$`J���!n΁N˲���rsF���Sq�ʨ�	n��-�%�S����l��궈��~d��K+��0�6����ހ �/��Iȭc�/B�'���MwK� ��炛0�VK����&B$?WL��5-A>��UǠ�	==o E��b��j�-�V�:g�Q9f��0�S���%��L��N绂�g�k�/z��{cˏ^�Lh��z���k��pf�3� ˃��}��|Vd��f��)�����@���2���Y�t�v�L���)��pٻ�9�d\SB��$.멝	5��N�D��:j������	.��MăM�*9�(}^9yn�1�&%���YsfWZ�X3�;kӃy˒K���x�FDi t��8>%�{fIz�.�B�e5,��C*{���������vt��1�zd�C��C�L�Ne��@��~��Sx�m[�zov�&v�Y*}�O�>���k6���;�ew�"ل �6#lH$��F���gf�	T�4A��H�>\OiH�K`wI����U9�O8��Z&�p|\'�ͩ�$����z#��`��<&3<Se����8wg	�CemI�|H���c2�B�ĺ.��1�4��X��=/�ֵ����W��M��옉VQk��Y�gMq2:�:f#!�,8VO_=�m� ���<��xj�����{ҏog8K�6�܂.��I����� c2��iY��3V`��y�vѓt�M)&�4]M�2:�a�C�c5M�r�cY��/o~���x�g ntO��r�Ň�谬�#�X-�K��h��Xl�5����z�F.x���do 7�FT"�,wM�S����k�ز�X�ōnw�d}�Ak�â��l3]m�A�Vʎ�0�a�;K��,.[�� c;�L�릶��;B���y��!-M�v�g��7�m%k=��t���,�6�a��_}��Y�t�v�^����IW��< �~���� �Q�l,������̼�$0�c�$�r��6������-���&t9 �O�v�'Ǳ�< Erջ�,jq�`%��,Swb�;�Bߣ�}〣��	�A_�z���C&���J�؀H$���fHA[�rS�r�ii���z/�<����vT\I  �ks�`����.ѻ�2����;2O$@�KXp�|I�{�=0�-�chF� Hw빀d�[�"D�O�s�;��w�v��g>�"sXm�Mƻ,v2�K�*�,A�/MG1���І�R��ԟ>��`r�˳���m�d�W��	���mκ�ױ9K*�����h?fXvpΛ���5P0{� s�@]F3�as�<�����7V�b��/i� �l��R�N�u�������K�N�=v��!��^�S�)y�2��y�"��<e��u�u���zb�f���b����b�A���������㮛|z��ǀI?*�a ��E<Wuųd\���H�[���vNC)�gz^o*�L�u��������C�y�� @'Ou4\u�-û��]�vo�1��M[�t�L�	Q*�b	!�o��(��`h��f�H�=2}���V�\��û4�MFC�KngD�4'�Ù��;�v��$-���$�j��<H-�}u���������:E>ٻ�̣��n�̊�Ý:�aZ��[�Hnn1�5���ݳ����L���Ukǉ���I+:�dn�J�w�����?o8���%^[A#DT﵃�,��3�PsS� ��1}���܎�?uw`���U��I-�}2X%���_5(�R�r�w���&/���r�v���=u�A�^�b$�A��D��H馗�v�-:�1��:��,��4�X꺷=��{�8楣^Y��`�b�ܴN�|:�K�L0�%M�����z`�S4Y�f+2�� �x{=�~��'�M/�g��u�]�,��gvcF�M4��,Nn� �����a��4���E���3�:E�q3���nLC�3]�5�D�xh��:d7:��וy��!l�/iًN��"����Ü�ڰb��wi�{,�4���3��{�;Ѻ8wf�&_p-���NPL7:�VbE��U�M2�!"_�vd��C�$��	�Aٛ�A�a�����8 ���|���6g��)eD�8"���Q��X6K0�':����`��;:g�-�=2	��+Ι�꾽���v���n�� v�`\�om�]S�Y�r�v��� ��1��Q���yR�`�$T]�$��ӳ������T�
���1M�~~�:�g�_�Q���}�fw������y��e���p����'H~�o$�����3�p�sBf�0f�e��{y������2%n9wD��C��]��* �A����79Ӳt�U�]���1 �� �g�	�������8!�˂]܄��^fZ��À�b�k
G�3�-t��Ʈ�-:�0���`��ӂ����ީ�I�. F��h��-����x5�&g��|{rc�XV좭��8p��EAX��p��Ƀ��}�0�UƒH9y/ ��g� �Rj�뎴��ӳ�8���0Ik�"E��D��Q��#�3і�x6��c����y0#�D�]P�O�5�,����p�K�:;vC^;�sOn�C�}"	2������ޕB����������8=�[�t\����j��=I/y��0�kWY�2���Dx�v���u���g�L�c	�we��*�b6_uK��F���)��YqzM}���=�b�N��]Kw��.\�6n��Ԛ������'����v/4��̩0���_{��@�̙��235ҡ�w�}�ū�������z�"��!w7���gk����L���dF*�u�WΙ
F�9v��f�Gk�G��by��v�v�=��5��t݋�l�Bl s�g2U�����AdL�w"��a�f��x�U析��% ��%3�j�M�Ms��A�hu4'oE��u�.�!j:II`��f��j�����?$�xƭ�ַ�#g^m�vq�âǪ�X�)�V偅����������\����@'�1N(�$�>���7}���!@�^�� �sj�F
â�8fr�1/X��h	��̯��v��U=�'ǹN���P�왟�_�S�'����������Lҹ�iŝ�3�M�3��y���ٖC��R����:d$h�aj�9)�B�L�^'�̚:X�l�O�r��P)�ِH$��˱��ge��
1۴�n��CoL��ˋ��� �{�ϘFN�zY�-�-z"�rd�X%���5��6��X~�֠���d���!��W@u!��� �-.�5�)
D��ܮ�,��P���/������w�� 1��݉'�	gL@5�-)�X�o]4b�|c�:$���]����0�pOY�`i�_�{��e�l�U�E��sMvwo{h��A����246(c�F<�n�!�Ļږh�E�]��E�c���Ŗp�	�E:�OLVdf&af&j0�� �� �-��B�ޙ2D��Tz<� gSA��p�ђ�Y�"�39wE��}؍$n����=�K3TK�'Ľ^d�$����+v�w$�N໳L�|kV�q��@�1wQ W3x���������Ś���W9����>������)8&D����p^F�2�Om����=cXsgX1[u	:��ف �C����S���<�Z|���.�PK��Z�nk�6��!۶/k2n�6��Y�S]�)�'~�����]�3�~��S�$�o6b��Й�y���q5�S��������J˷,�o;t�>"6z�:�y��&#�t�dƝ'ĭ�$�u���/۔��kU��}�H��;�K�o:t�%����<`�ُA*� 6��P��1���'r��2K��B�o�������C���Ԁ(�����=��<�O1)����Z�ZA��^�3{��4��������'�H���?&���G��ws�c��������nT�=�5z��rN����h�y~���6�ՠ�"�g��vuzI�}�j�eW�w{<�:�u�$�C��>�j�A����;5�tj�ޠ����}��.�e�]�
A���xf��������[��s}�m�8��ӧ�i�u��f{�|f.��#������]�/����.p;�M�o�S�������Qe�r�����1�m�}����e������9y���m^~��v{�7�e�{�`�eM�����d� ���{[��ۄ���([�6��N�;9��y�zt��6�x�� LO�{^k��uz�����㗟����vY-����6C��7.L�q��VvY�`�g�z͢��[���ټׁ�����X��y`���p�;ܖ��o
��w#�W����=��*��5q�$�U�����bOG��\dk�q$;������֙F�5����n�ٯp�P�s$ǖ���s����&����{�wz�#�}� 缳��}��pЇ��y�����|m�������Lz�G�-om����\ͻ�{��闸�q��퐾����yOu������8zW�����<&�Ĳ�T(x{�W�(��\[t>�\sL��'P��);���q�TB}������J�d���}L^�+�3��2A�9���/��HgK�컧J����n�xi4�H�ǂ�3����r���������a�_ز�
G��ŨE=v�pD�!"�Y����EqDEPTB�� ���<4���(��/���n#�$�=�y!XG7n����>�&���i����������,���9���\K�S��~$\\\\�M�	��o<j����-)c`�d�i"~�NN%�(�0ATԈ�#�l�6� (�\�#iJ|p����C4��I�,��%,�l�8�"���Gd�f�,�����@PP�R���4H|i����}�� ����D��̒W�$ݔ8�""��!N=9�dW*�`�ơl�dpD"���
�W>p�qѼ��/j.�i�����q�m�n���.%��dٚ�R$Dq��Q��-�rI���)�����8�^CZ� ���4E��5�����I"'a��� �\�Q{�Sl0d�>X�rɊآ��«d���Q�#����H�L_A��fVjY��0f,>��� �w�}�A�و�y������fr���Q��҂<�gĂ��e��$ ���*�?q6�:�/bb���V������5@��ȃ����b|zZm��Zny���	���2<H�&/��Ă|�]�>-\/,#�����%��\K�"lnؖc�D]�	Kk���2�Л-����Z��=?�d��VmW�~�;�.
w���J���B�4X���_3�<	
�Q���3�p��}���B����Z������	y�x$��~ʐl%y�vs�-��ר@���n�����U`��<�KgnD�O��T�@M�2�ިi��P1W�$���!t]�.��Ӑ��F�����6{iG�̘Ex�^tI��[�t�L􉨦舭s:�tE�1������h�dק�iN��^�{�=N�4�'{m{�ga�wO����%��e���g����#�ė]wz/X�&j�Sj̛L�ʹ3)��zϗ��������ي`�
�g��Au���>�l���NgE��M�י����E��d'�������8��h���l�ݖ]t���ɮH��ݡ#�c�6ˣ8�E�[|�ߡ���霮�6��	%�7`O�$wz^=f�¢^���֗�C�{vD�8�R���t��У�9S'Y&�7M�z	`
[ד��w�pd������K�
��ҙ�$��<����H<s�"�tI��V�ۺ�I��b|A�����yn�����D�񽫳�N�����?VƒH�[�d���3ح�H��*�ӗ�!N側�m5�6�'����"*vo`[3Fc��?
�����>$���.�y��������4��n����7{�g�6Ӣ�\͛֌���fN����>�����sP��ݳ���7����M���28[oD�X�����g�q`�	z/L���F`�&`Ø���y�m�a�c����ܴ\��on�˼U]'u[p�S�Щ��[e�f.b�3a�q��dݰ�,Ck�8U��+�ئĬ�BU�<�c�^�Up��v��a�G�61�ulu��I!:3U���H^�ֶ7XL���m����d�i���r�)��V�tu�؉[��Xs�hɬ�C�i0l
�g���Q�����`gm��q�>�6��ϓQj���n��q������G�3�w`Ƀ��������]𓐵��]��(�<=�c�1�>$����R-�᜗g�ʯ�9j/��9��)��wa�5�	З��� [y@$R��Yl<��tf��X���2�d�10(:�kq/+yA''R����,M�D����	�`����=����sw��mnn�A~���V�!$A�zfwp]"J��� ?^ۤ�o',]��B���F鷸U�=r��9c�	�؀$	
ڹ@$���2=[�,Ȥ�bAْN�;�����뷧���qc[c��ח[gs6J�C���/R��~��d����̫�u�z/����
���4�Dt��EH����O��=����Ÿgp����y2O�u_ig��>�������u~�T�R�.�dŞ�owp�~�__7�w��� �w�o���s�fV�Ff[m�A���}�əY��٭f�b�;�||^	x�c���}�}2[Mu�i�;]`�0g�_į7��S��=�;�]��n���93�Q�W^o�$�PRjgڎ�.4l�ŭػ:LL��蝽���25�f���u�����[\((�Qq�X@���&A ���V�5�"g���`�",YI���}�n:o�I$��.�h0�VS�Ł��H���	���E�cm��`������'	1.�]�nnyA�n#Nڙ��ι7/?��:-�o\Hg~�?y����.��`�,�׉�&]�}i�ᛲ=�B{y춣&B���Da5;x�����י]�R�bm�S;r��ε'��F�χ�$��i�2��$�h�6	�<.Æv�30y��ْ$��� �n���(�::Lͦ�m�K�c�Aw�9�;}<��6���J�}��5�^ނ����B���7��N�}����,t��K��(��d�>34f�ՙ3,�0ֈ#�v�~?>���d|g�+rf��&p�죩,�����֭��"�y �6�w��v�A>'��U���,����3��GT�#�I\�&��Γ"�D�z$�n>ۇ��f©m�g��F
��>Dh!t����:�8a��v�`XO��d2�fS�e!���t�&��]�h����è���s�(�h�^M�p'Ĝ�ȊJ��7'�����6�E���$�㻹B���8%�鋵P&5�Q���;�*����|I>�술����?B7\��&/XQݝ"E�n[|�����י@�����6B$�����x���~cCuS�ȃ�� @ �i?(u��A�v�30|*ڻjh\8��kC4���N�6> �;�ӣ���m	�1���?�
,�3������R��7���ȗ�s)���qh������|��l1��Z�j���=�1ܽ&K�&�{��}=��?��G1�LEDpG0G���?߸q���r6�t�;we3�md@5�W�9�t�[;�5�2�-�K�D@$a��  �v�(��Q�O��W[#1I`0��令Fg��
ݖ�z:#�t��4�y�E����r-~��[G�g,����؀Aچ��%���BB�.d�'�Z��t��q'�p�`}��W{wI3���Y]Y2	7�����_,#a���%xu���$���~� �2 �}�H �>�y��)�.��L]�]\�l�KNnD�	<�+�\�Ό��||	�� H����g��,�1wu�P�7Vu!�8s����$�����>$�1ޜ��Jf=9��`�r�	ؖÑ̍�ٙ ��q���9�c�cVp&�Lx�MN�̂	�܏F�,�Ғ���#��OS}�"�B�Ow17:H�Ƣ�(c�����z��K�;ozC�D�Fsۦ�Z����^�f~�]�e��Q�FK:�=6Řf3L�3L�6Yl���:�2WJ�r�R�K5�q=�L��z5q��m����ú����l��6��ᰵ��㫁���u����֚�5�u`�Q���͹���u�;ͭ���!^.W�3g��Ӷ��g��T*f��XC-8��`s.�e	�f(]mCt0mP�9�v	2��n6|�Dd�u���풉��v�E�QD��Q������E�^Ʊ�=�\��Yu�c�Mt�rMlh��-��[/����s�N�gv]�m־
� �����O^�Av�ט�m��}�Ú_�I9;}"��,�R��##雈���d���i�w֨�|O�{�d�I�ۈ��Ͷz���g��|	��38,�}�}U�A{p�"%�m�Ң�6K8��� �΁$��$���)���,�`�S�����r���>�k�!"A��x�=�p4�lB��X٠�Fm��"sHN��w^u&@Q�(=��#�(9ς�:�-��!ٽr$�w��@�Y��d�Pz+{*��I�dͮ�筍�]��t ��]������� ���5jڡVs��	ؖÑ��ɑ$�͸����WM&�u�e����w��u2O���눑]��lr��;��h|k���d�����U,�94َ�QQ�i��oww�2i'�y<]1S������w�!>t�R���<���*՞绵����՚3,��,������y0/Ă}ٷ	 ��	`�b���1������͟�%p��Y� �Y�dp`�鞀!�&z[` Yv
{)�b���H$�m��:��` [��Z.2pX;���G_Os�j�Ŏz�i3��;�L8�m��$B/�%��8s�_���\{˧)���d�D�9Ј'��;bK������J���/!�� ��tE�D�G��5;#�#�f�MfK4݃R�Z=rW3;�!v��0����9|Qwf,]�+x��D3b�A!�w�J��f1�W��=�X(�Z��@�Xo��	�1N��w�y3�~�ڎ,ugNkb��j$9C�A$���$�nfaB�Z;\�Esl�D+6QM]�'��O����P۝�.$X�lz�ߧ����3`(��yJ�9�bj����lw����S�Qf�-��u�F�M���^^X��������NŲk��3����q1�GpG�p���s��!�����DA>���!L��	��圦F����y]]7<���)�K��@�	��ۅ���k��#�\up7�qIæNYz��=2 �}�^��Z� �ݒ��~��|F��E#I���R&Xy��V{Y�n3��h�+D��R��u�H/�c׆�t�P�[���n9�31�|�7���ݏf�ݑ�ʡ�BF#n�� ����>n�p!��ƙ��'��b�w��fP�Ψ#ĂX>�mPAC���� ��^��=��H*���dS�A�]��Ԃ4)���-"�tm��·��Ap^D?f��ƻj�`���!&���'���s����T��� ��\H$8HC�DG�$��cu�������E�=_�m=\&�"�V9i���t�yUw"ٵ҆�0ua�n
T置W{}��`9�a�<bz�wϟy�q�}9�>z����`�1�ADLGA�������?xx|w��w.�22'Ǧq��'c�5��C���o��s ��^�@!!��"L��]��������R�A.sJm�LmCA(���CB��(�`�1R�;l���]qGbw����6�fvI;��5>�{���H�q��%�m��oX�ewl� �ߪ}3Q*71ç�;��:�"v9��\u�Ǟ.'oZ�c> �ݘ��I�����<�1a���Ok>�!�E�n��kB��΃�U�c��@'�FG���=�n[FK=	�3z�O�o�x���z�p��dS�A�E��L��%e�|����I'�M��}�*�br�i,����4�$�>��SXN�'��̞uwA�[�;���γ=i�bc�b>Ў(� ���'@{�86��;�xO��a|�n.����ݯϸ�h��;�^]à�������i�{��'(�Zc� S�.N{���%����������{��ri��[��ׅ��{vxe�/4�K��Ý�a!2�4� p���6�w%~����}�U�!���ۺ=�������|��o��(2H����y�I/]�1l���i�Y���%�}w<�!%�sݚ?d�p�Q��R��I��I=#�C��}�+;�Q��=�Q��~
���}N�TEs���[ц��ls�˧7����r���;_P����;�~��`�&]=�{V=d��p�>'�yo�.A�9�JV �toop*����}u�7�?}p���L�Wf�o!Jk@���y{�l{2dպ�C����}z��$�����u�_x��n1{GfjN~�`��-8"����U��+�^eYla�*�z�R�L\�ݷD�7�N�{� ���c�hf�>!1��Y��;̜�Q�u��;�u{N���mYʦ���=~h�:�¤�ۼx�����;��(Y��4�Ww�=�y���?[�ђ�����[`{=�.�m�oqz�!7��5�rs�u�v�����d��_:�N�S����aBon>h�]�x.��e�go��$�V_h����I��uzq�w��j����m�i�5M+ݐ^�g{:I����L�3��0tz7�n�M\���=�`�|;�H����-'��v��~�}&����C��p0������%��q���v>�А���7��� �I������]x�#
�㦽/X��3h�OUl�@��#+
���M��cv�Qq��1��vGarE$�MI�U�>9��9�B߆�T�]G<����]�jl�w�S��^H�5,��X�̉P+��4JS��+����8�g���,�l�ɶ*�E�]�H�J�[	1!ON��SX%E�ɑ�W*K*�V(Ff�D�$�f�����<8xo+�E���G6�R�4��v��"��q2%��vE����N���7xB2m*XLX'�&se>����l�'�g�C�QN$wb-�d˟�8|xn�9B�;4A�M����R�ݼ��%��q�+\�?%i�[?yH�4�ǧ8o4�*�+�H��-jbોS5"5���F$$��$)�t�9tw.�["�Hk��m���E`��ь���x��r~���*[i)��Ke����m�Q���8l\� ��Y���_��Sh:j-�\ʌt�ٙ�E���l�����-�%K@65�l*�4L�6x�d�����E,Xݻ4\�z�u�vMYt�6"�G],\q6�k�v!8cLxsp@�9�_�;�UEA�o)�����\=��`���.���:;�"�:Y��Q*�v��8l�oP�����6̈�Gs��lю�vY^�2�q�	���d�N���+��JMg�#U��u5��!.��Gt�[��84i���,C� ;��A��tq�p1�lN�Dp����<S���x��y�6���m�����6����9�%���w;.�-!�	
��P��liJ���[�۴�sb��Fm3��9���F� 1]�Q�i�����<����]�#�:,�/kCs����m�E��'h��tqy���q�9ƙd�0���vmlm�\q�Wa�^}u\<�t����kmnc�㎉���ѥ/m��4�oo��G\xn��9�W1gq��=d'�d�:�Ǯ;gì�:6ܖc�;��Y�܏��g\I��p�;;m'l����:����/q�OL�����Iu��ϟ<R�Iv#Y��q`q��`�;2�%�R�l;���j���׫k.��rQ�v��)��듢/X�l�Dv�\�9<���p��`ZKx��W��厯7a���d'�c�3�s��p�k�@f��,� /N��ޭk�U���4�;���X���+�;�U�d�:�#���L���]�gBB�`���,���R<g\��T�uНA�\��m����w%��[�;��u-��6�۷b��V��`9�YoZ-��!�āɉ�u^�"Z�.��\�$���8	yJa^kr��Ŷ���aj<C5��49�M��M؍v�ǲ�E���j�q�N�����|����k\�e��r�;`[�Y��a���M�{��v�m��M瓞1���G1Gq�Gt�O<.��,�Klۻ��F9(�ϧn5r�`%;�ݲ�);����7�g���]úӂ7U�����X�j����}���y�v�cHb���jhJ�"m��hV�B��瘎�}��K���рsAe�2kF��v��h��SF���&�LY�m44%#�ֻ[`b���ˊG�GB-s���p�O:��V�pŖU���������qa�B$66�n��ḹR�onz<xy@mv���p��vd����)��3��,���ٜ�F�
�N��Q�� �p���0֏K�i1َ �֎P	V"�ɝ�fvI;��wML��3��y�&q�6lHH�mfā� H�c{:���s���Ū�_6l �]A����b�P�O���*�:$8KĂ�.�1C_u�ǏZ��I �a+�"K4�9L�*$�ݾ����_! �y�J �lci5h������+���
�E�3��}�$������pJ��oF H�k� ��rd����"c�!]-��ǈqX��V$�n��LhMrB��Y���\�f��{���!�4Gk＿���e��؟�@'{j ܶFG\�ٜ�W�$�#.�Ran�ؔ���霈 ���(j��0tT�t
f�E���57��2�v��L��m����r�CQɯ��yc;
v7���ie����F���g�� �b8b8b8*&#����ɼ�TQ����q���=G���V�!����iR:sŝ�&t��ą�="@��&�xl%�g!?NM/4nt ���(;��Y`�EQ�Q�sS��ó��o��%`�F����$G[E����[�r#:'�K��:L.Q&3�E�˵wN�����3}2I>=�O��ޟ�v�+i��u(l_VZQ �F盧;���ұv�қj�)��b�f�"�}�����d]�0~�UnL��@�w6�H�	R5G(6!��Y��s�!S9�@� �m��j	f�S"�2gs�ܮ�5����U������cp� ���� H�i����!�td�뽿F��I0���Fh���f"mG@�|v{1jc�{=�9�������a?A�u�N��~a4������9��w}��%0I�.#�`��1�<��O^N}��>٧�?��&"� �#�"����<?�ٓ���'9��'���x�pɝ$��y��T<3��l�g�Qw;�$o3|N��C�LuwC�Z��჆�#���ڞ�Z]؆p�C�u#�۴o��8��>&�Wd(������`���Dx��zۤtM�CY�<煽��R�(gK�ц\��Z��l�7j�2{{G�8u/H`�/',���{��&��*8�mG��y�������huM�U79��݈�Θ� �J�A�Ļ&`�"�zdM��ϙ�q������N$�}Uf��e�h�"��;����t�w$��)�N3��-��`�c�:$�3�E:ڏ'ɠ�;��`��۾�����&�39A#B��8&��Kh8�u�Q�	����^D��AwL��C�)� 0��Q<��Z�0��l�k�ap��3@�"p'
�L�E�ΰ��#^T�8���|���󛳾��>[�?�8��9���њ�Vh�F��x���^v���Wx�p��v~G�麡D�r��FF���i�S��$l�ё(��� ����e���+��{>? �Q08u�&�Ve*0��]]4�0Yb�������Y>Gn&���OФ�	��}��R&owb@'Ğ���ZM�K�ܗ����=}��	���ϻ2	gr���B͢~�#�Ĭ������/6�q�<�i �n�g�H�|y���t�k��4�u���&�U��%�3�����A�ہo�ڪ�C�2ٝA�p�!��O;�����W�T0n\!nFmfD�}�� �l?B6Y�V#"_,���<"&g($a���9;P�Z\�H!�-uxHx����Twd� �Hm���ܤ�ɓ��S�%��6��;E�<1��6�ج�+���V�BjiU��=X�{�#s���O��r�ʍ���}7�g���=��N�?B�$�bo�������7�r,���uh��\WA�G��u���L��%�,�1�tsH������M1Y��v��Y㤍z��m��;&`ѹ���g[���]��λ���Vu���壡ՠ�n�	�v��裦;p�!^۲�nZa�8}Wg��ڳ�n7u7ns��I��Guw�w>.1����ݐ&|m�S=������ZY�7n9�np�h�u��8������n�zz���/R���aG���~϶`���?|>��$ov��|I#:��I��q�3�gT� ����4G]c'f�7����T5�X
T][h�~���A&�i�D��~0E)�b�&tu�^f��p��p�S ݘ�����@��懨�9T���`���&z��+����%�&/7�qE�ĝw�Q��'���	��c�D�Z��RڳK���&6'ω�ɭ�9�۸I�p�Ϧ@-��`A���4���7A���q{!
��`�	�uoL�;w�QW=��ց�n;����6�l׮lz�6*��\�^{��;B�h\��23N�'`�xp73q �m-[� ����A�H���q���}�%���g��3�a�;��23��1���?�����"����Ç���'1q��h����w�I��t<)�q�E��t���8v� c���߿=��l��kf3M�+Z5��A �i��I�($���|I���OR�:�vm�~��vf	�o;V*�=m= 1";��I$��s��~�l�PK��XѨ`�=���B:�1�p\���UF:9\�h8j�t�A7ͷ����ދ �[�mo�7NН�'I �J�� $p�kE'D0vI���ə��읁
D��p�Y��� �Ǐ$%���$�;'ba;����HM�$��{:�A��tx�k�{ZT^�/bX��@� �]�i�tɓ�v���&w=�6��"�6$�'�ӱ=r���k��R����=�S$��1�E�:z��	�"�k�ע�P���PH>���BQ$���JP{�j�Z�6�G<We�L��fy�g�ْ|H7�1� �!p��ۙ	�==L(궇�vYV�ǳۋz�Z�ҳ#,
��I��"G0�ﴇ���]˃S�6�F�v|��}i���LqQ1QQApm���s�Hy{���
���و h���vf	�o;U@��ϭ��T����{�f��O�H$�옂	Ύ|Og53��	@��#:�dO��`\,�`��Fx@$^FD-�*4��<�ē�|o�bI͞x����9#�|����?vԷ\MB��]n@����ٞ�H��]�<Sm��seD6Yz������fA/�u�3@�=�P �H	m?<������՗�q��j�	�-���H�.�1{�A���"��"q��n��H���XV��R?&1����yg�E�$x�A3��K����*���ú�S�$�Ɵ�2���!�u�9��yx<,�Ȝ���D�s� �[�k։|;�{`������K��N<Ue�fp��3<�]�%�ʜf�Q�L؁ ���@A@7ѯ�����]S�m�$C��G�Z����`�y,e��J�y5f�����7f܇p�%`ț�,�_n�Շ��`ɕ;1X��A��{�	��a�\�*:����������5�����͙��mfj���?�?}:���8M�`�}��`� g>�� �e�4��:�'��v�@�r��A���bΧ��1���p	C�y��f��6�K42���=z���g��w^4:�1�ʿvn�.�pK2v��e�b���<�H�}2��P��n6�c]p 5��z����_��b�7]�2E�5�Сv&�Ɍ��I4�-��"	�}3�MR DփO�m�
����׀�p�,�	�;�@��Z��Q��F��N�:��O���M,�h@Nlt���'V���L袕
����S])���b��I'�]�>�@$�#�W��us@��fp��3=�y�gfI��}�K�h��曶�I1W�2x �6Ή$�ev�gu��$�SL�4Ǿˬ��ݖKwd���93ny?oa�릫�_�w�հ��X�yI�q�:����nv�� ,� �prٓ��y�'6�� ��=lM>��]�c���W=0�K�ˇFf��Q��f\c^��#��/fhݑ:�4���Tۦ*�4,�<�^W[��#��1�2˒��p��<����u�^=�^#FmX�6�mx�b��5��#�&��cm�8�=5�=#nU$�{&����{ ��uaq��'��a�U=��L��K���'O8l��b��a�raO�wml���qy��6���_�w�+��������ށ&={�I �l�C��]KI��}��預H��ِ�W8.rK2v���b	�}����4SP6
�	̝�$�x�t��<3��Ow�k���p<��e۲H��9d��^j[3 �|{6`A�ِt�Cf.1ډ �y� 	����]��2tX8L���Fj�#������8@'kw$O� �[�&�Z�y��T��!�h�0.���TLP=$��V	˄R�gjnp�t=ʀ-��m54���B޺fL�׸� W�%haޖ�y`��h3x* ��)̓:rY����� �f0�a��v4��	NY�ES!�Ō��݃B,�]�æg�X�s>'��ͨ�I��.<P���1�v���O9�@'��eG��T�3b���Ӊ���`&�i<݆�2Yt��ܛ��⭩�©9��0m��Q>Y#���6��U��C};��������3���Ex��*�R��Vڔ�Ŝ��>>��!/��y�	}�� H��Zy�_(:��o�0*����s���w$�'g#:v	$N������w��g�3q�$x�t�pK��)ْ/�Y1s3�]X+3��tDl���Hh� z	$�˧��PA5v�v聅��h��K�����&�;��Cu[� �ΌVޓ';Q}��#+�#Ēr�^ ��ޙ327Cjɒ+�+ł`C� 8`�I`��X�\\V�������4�0].փ����6��;D%���� @$ut�D�w@:�dk���VХ�<T��sr\`j�v�;Q5�;�}��Ϟ�����>�4��*,�fLd�Ğݗ�|O�"{zP�"����>P��z��ݙ��M�`��Sт=��&E����yk�"��a���.�[g*}ػ?����3��gz#|�B�{ӭ��m[�jvh<���߄��{������G��v�����AᗒX_��g��`~9u!û¯W�˥��<��/\��6{����!i�����/>����3�;����||	?�j暼!���#�ϼo��	��"h:Q��=�=��f����=J�����Վ�9y��3�{;/�g8%�����z����N�����?�X7Н)E~�W�-��{<���n�Ɋ�{ٗx������Wf��Q�|�<Pg|K�O��B=7Xt*n2\�Vl���d�;$}�	܁�kυ�<ٚ{l�&�b�X���l�SȥtoU�չ�{D��5ب��{��iK:�ذuy�`�7}ܹ�w<���*�k��aT�����q���X�i���RY�����������w���]���xZ>������u���XqՃ�:zbV�04k���o�ڡ>���e(p�D���B$��<E^�=;|ApC�����vx/g�����f�<��3j����R4�S����ܾ��F��.�;���Ü��^r�'I��вq͗zk�z	�\ ]�k����;�Vd�cZ���h�1��]ޞ�װQ��eÒ�]�����??�tKW����~�+,��~r��[�Y�E��"d�zp<�9�/-<|�z�5�^����=oe���+�/N�N^�4&z���a�N�ʧ��\ㆹS��\�N�k��Nv���>�~x�j�8pg�7��bu0� n�y��^G�G� c|���ʮRo9>y�������7F�v(ȐG�$Fk�f����U����H8��
2ZV���Hi��M2���.
Y%�Gf���TvA�B[*7��ۈ ���-ą�s�G������6�A(��K賋��c���u��dl6b0�ql̋����4��QԈ�2����E9mF,RlȉdQ"��r��r1STF�qHB�p��J�a�.>r�#�>�<�ѵ���RRtB�s�@��Au��P�A*[�$b��Jp��⛜EǑ��e,!l�"��-�W%���"N&���rAf����#�Ou��)�������@��8����>��`�!P��A�v��5l�	�JCM8zly��ԞN��Ŋ����H�A�K2�YX��<6���L ���H�X/�!O����{b�|��rH��[0�J�g.V�����ԥ��u��+~�I��_!UX�0�*>]��u�j�l���`������a�f]"(�.G� ��x�@MN��E�K�t�"'{�S��3��.��CwEgcm3�uv
9z����$��ː��<Hi�q`�W�S���̛N�Hv,�6���(.�ȉ�ʦJ�+�n{�	eQ��3}2H#{.!�:��,��.):o�y�.�a���mB6l�u���I�+c�㲜��E����g�t�#������L^f��;�q��kcfp6�b�A��Ȑ���
�8w�*2z�"`�Q��h5��f9�H�R��gƅ�	K��@ ����Z#kc��W�JW������+��h�{n �K�n2֧�Ǎ"��z��m�����pv���鷛IcI#��6\:Z;+^�"Un�����H$pG��	�ñ͚akaf�N�LӬ5dL�){:˸��H�{F2_9Q�'#��oz�j=n��vYN����d��|s��b����Ls�pA> I&�dm�t��T�����L�4@/�LD������������������s��$U��/<��߹��r.��K��f�	vm=I����Mtت)�9h�1f�"���|��.��س��ݺ� �A�ځ$|O�lsAф�[d3s*���Nd��"�[+��$X���3�3��jʆ%���a,}�;6�o�h$�ܨ�H��S�ДT鳝�Fk4J��ܶL���b
�t�`��Q��$o6�l��NK�w�CQ<�1>�h� 3|J.���&O��!���8����MwpA$�֌H@���}�C''�� ���wfg,ɐtL�ԣa�'ǧ7bNX-��N2�[�ӕ�uC�ĳ]D�@�� �:v�d�⍧'uOI�e���wi���8ܫ�9z�\����\�n�d��I#�Q�kY�i��6�b�u��T�@���g��D��aa�r��cN^_���3��LC}y�<������/e�\��n(*���l�g���M������d77�<�Z';mѺέ܎w�ur΋\]s�ֽ`�Y�c�����6���V��(sYv{ˣ�iv��#(��c5��qn�>��~���e-��%�t8�h���Ж;&pl&�(Yi���^,���!�=�c�n�h�lI[��4K���<��=.&��j���9�nٶz�c��y���5��<=m����ۏ�����d��8�;W����}��y�e�<��$�����b��f'�sT�	��= �}5f<H}&��I�%س���ڙ!6Z��N�-�/`�!/f��H==�a"�m�%<*s��M~|��C��b�fq#��M�d%U��$�J��Xr�,��|`��H���Hi'`{l̝��b
�`�NP޸=	J��f�}�I*!� ���8 &�wN̒<	�Ʉr7�XMO���ǉ�%wvvN'"g��3�D+��0X������"��	=y3�A>{f"ŷI;��)��2�D"���;;�3vpdv�Ϝmn(�q�l܏F�~N��N~'<L��	3Y����Y��v��e�A��'k��A`P'{b ���
r#�ICO;����"A<&.�ӦE�b�3�Qz�}������a�Ͱ�S>\�م��g��e��=�CrroΠ{���F�ֿ���w�Y��X�]�^��Z�i��j6���q呓�0H!�0��A	`:�����E�ٳT6�]�\��nC�eقE���m�3�@��E��EL��,//m��
9:�^6G�t��3��U]�2	wl�zD���ᘸb��U�j�ʬw����,@H��LO�t�Lʼ"O��{x����|v���m��M�p5���`[�;u�;$�?����c���s�H�d��J��n�aAQ53�H�Ɂ �A��x2&⚟|њb{8TL�hAK�`�,ּm��*%���"fmF.���xh��]aP��}���"���ӱb���#f|A�ُF�H:z�H&1]��&j0"A�ځ�v��&f`�D�6��7�j^hf����ĂI$od�H6���]O4�u9�Y��e���X�"�M�_�Ӡ�[�DL���s��^�S����
u����W
�a��W��ه�T���SJ��TyL��e���c��	�����p5{�Mon�ەz�#���I$�O�U�~�~�"D����|	�Dӄ��v.�dE���quKr{`���<x�~� $�2v�g����{wd@G�g�=�=�C;�b�d���+f��՛��mcm��k��8�m��gnDx�|i�dD�I�V�H�GT���W���Ƚ�.�voR�d���n<k��<�j�`��d�Y8g�\8��H羁����&�u��OYm"���r�4�A>�����3xRr��;22�GL�.��.�j�N>O�=��$�z�@���|o%��fmn��o�x���;'r����u2׮�s۱ cGfk���v�m���� ����aL]qw%����gz��N�s�*�K���ѳ	��ft�wtϘ���o<��X@�EA�&��p���y�*8�3j�+ڪ*[^�9�k�.���|.�Ճ��Ѥ��7��&KCDږ�8��\�G�h�x��l��/�	�vH�����q�g	�v.��؝ȹ�H$`]�0"�-�?Eǈ��q�����I.�T�28x�rgZhÑZW�R����bɠ<�R0���1�jmm�5n�h�q�M���b긱�t�sj{&�bA��#p!�W�jߞ *{zgĆ�_��ɜ�p�	Wd�������I�H�X"��<bv�d|GwL{�d�����G�k���N]û�vA���t̄�&���HF1��2��� �EVt�$�ݳ�6��æLΘ;L�F�v�F�t��v�(h��{���<�X3T$A+	x1�٘H;|]�g$��3�
��d%�M���:�n�x��̙2� ��Dx�;���:k�����wt��)�"Z4�Ḏ���8�L�w����8N�d<=�\mTb~��_i��"0r؃��[���eW$���#"J7��ŕQ�w���f����;^��p9��/^�K��v<�5ś�FCDL��͛��������i2庶*3�	�`�f#..ghM.-ڐn�l��Oa�Q��CnF.ݻm��V4�g�Y{T��j۶�v5��ېyi�f�
6лp�u��x�I[st�cI�]V����ĝ���4Vv�mu\n�%lAˉ[L��.jL��;G0��y�L@�kx��0�5؟���y��0���}����$�N��A�,�nx7��j�d4(#F�Wٳ$�z�`Dnᐙ�3�2p�$=wL	�)�w:�&|M����O� ��<HThc�r�97]6g�&�8%P�vb�$����H�e����wj�����̗`c�@�O8�pk����\3�t�=PQQ�N/�=S'�Y��n�@�
/��$���[�V��#Y�wl�H-Q��gd��&gL���;>�%�{2=�c�!��U����'ӗ1$����#��$��S��y�@�/?�?�&�[n�uܬ�,��ۍ�G����C`�MR妣w}���f�&��ݓ�>K��''"$;}3��`�O�B���@�I�x$n�8���&	ػ,�OQ6����S<�uD��ZC�2CAV)�A�f��sE���fn����M�g��}?���;���j�N��������nx����;3� �d2��d��Ȕ9��3DCKngc��L^ڐ��3�2q2;w0A>7;}H$|�͋D���Uf�ME�-���"g�Q���I��r�	Y6
×Z��wgy�5��ǌ����d�|{�N�*�ovWa��D��Ǐs�Q�)���A�U�_��	Dn�"�ݕ�xm�c�l$�9�ꚽ�$�{�lL��k>F��g�8�b����f`��;mÇ��󎻍�N�O�5�QX�Զݾ����ݝq#3��뗾��uotH$�]��@������{����G�9����fLŊ@���^���Րx��VE���A &{:g��@��!�v6Ӏ��q���*���3����m̓^$m�i�]�e��e�^�����/���a��en��"W���t�+G̿DO
|X��<���x.#v��ASCM�ۉp�K�'�/�|x
�XF�	�3�A�'��6й�(��'h�@����	�9߭�ѱ���^M�W#�Y8z�`�ó�Z��S A$����l1G�����W�s��.�x$�s���[W�n����������!�S��.o8�Ln1�u��]��D�j�l����v'﷚�39fv.���2	'����O�x��<�p�W6��,ws�q}2$${Pp���wN��gt��l��A���������I �	툏����a �4��c�F������t�aL�رH:gi��LAѐ�"�v�hm��O�	$����A6�9��@n�*q��3���N�n���D����A&��:���T���r=�숹x���i#�����
��;�Q\����4�[�5x�GL�o�X� zn�)�h4Z_mUX��P$�C��ly@�O�A+�����M�tM��I��� X3������I;�2GO1qU���$@Kڲm�x��؉6���WtF�j�����g�M���4F�Hk�kI�L��&,tcrl�uS3���8r�ْx�Hf��Çg�P<v�"�$}�9��ӷ�&��%���P$.�ـI�q����!��3�t�<ʍQ�#ė~{���.j�����+���Y:�I>��_H�^�B�G���u`�*sY�:N�Ӈz�ƣ�@�Wl���ڬ�"(G+� �V�4pCU_D�E�9U�S:v!������n[Ζv����fv<���VdI��Cy�,��L����'=�!�S�Θ2NΘ�������ǳb �*��nP��&�h�չ	'�{f��� ����GX8�֦y�����B���׫���C|�z��{��Ej<	���Ļ�.;�î1�L���9�1�(��=Ңn�C�[�ѧ�����;���8A�I6�������Ld�Gܞ�̺��NP o�P�uwu<��� ��o?���}�_�==�P���M�y;f����q-���^��o{\^��>+�����1-U��;��A�׎y����]��=���Y��λ=����rF��G:~�Y�M�/��(�]���S �^U��n�e�_�7�S�!�x��GR�ux+G�
Z������B�����v�X��ZL�A�=�T#�xa��&�l�Vov��z����6��
yM)h�9굟�F9��k��܁�P��hd�!w���.����<<}B�5=F� �wy�% |�w=��z�����n�GIs��g��	�7��߯�oM޷w�\��q��gw|Ǫ�r��jTq6Y�U�'ϸ��m4����5ë��-�_�;�Ɯ�^Nxߠ��
�}�_�s�f�h>;��N{;ٶ\�I]��v;R]�%�[�gR/z��!1��^����Nd��	�5�����yx�~��q���c��釼�g���|]��/��;i����fL3	����r/���xxm��u��<z=���;���8f�n��׷= 6&������T�kuxU�\z����'��<���{��=a���3�I�l����B5�T�KY;�!���fO�d>�˓R�*�����[o���B��4���r���מw<����域�6�7��QN��*�8�0L�5��X���Z�:)�=U�#�a���q�ab/ogqw���3Ji3����]���|z�B�F۴f��y5C�K �/$�Y	��ɓmQ�QJ�p�b��)�����q?���1~��*m��̋f`ȸ(���噩UUPkŰ�!
iӥ��qk��EDd̊⌖A�^�RH�D�@A���������a�c��b96A<ks�!N=8qW�"��.��8��	�ea�"��R�!����8�|$)����H���B	"��wV�Œն��$ )�"��(I�=!
i��w�`��$�%����H9"E"L�2�.8�A�-er���}�S��ÇƜ�BHǗ	Y���8�qkW#�DrM�2�UURH��E�x��+�cd�Hi���N+�2a1V9	Ƽ��\������e[H�d�T�㰶Bd`���	����OJB�<=9��$�prKn!�P��VJ�(��"F}wsK$*W�L��$l��H�`�!b╥d��϶(�X���*��,b�1�MbY%b̎BH�**,�0��
�!Z"��Z4V�����+Sݥ��9�f��&c��2�;�ˇ�ؐ�GWm�oj�Z9�v��p�qr��d�-�\\7Ok,���41�|t�ŋ�)��V���a�f�°��i5�t��Jm�5�.i&��V�۱���S�y<ںC��cڅ۝�����J'���`��[�]���u�:d��t�ƞ8{\`):s��4M�������<1�n��.I�[��n��zk�n����No0sqŧT����������#K�BS�ָ���n8�{�ؗ��̓���� d����<�:�%��5���=E��yF:u��	:�lK��0��ݹ\Y��f�=j���ϳ��:ؒ;\��%�c�0��b���kj[1���!�zi��0zĦ�D�т�x��\�ЂS���|��s�nnm\�)��8S�	�tyc��am�H�)3�F�]�6e6�0!��4s�zճ�7t�VM�����5�]/�,o3ՅB5�:��8�[�0��F�@[eKxR�e�����e�S`�lV�bk��7 (�sM��U�A3�h�q���ѷ�%"D�,���S	M��-c��ș�Gm��Mt$X�l�&U��aި;\ꮉz�ǌ���Nu��
��/&t��mrv��b�4���M�]�7<vz�m��;L�r%���қCq��D�X����Ysp��s�rK̄���s���u����K�sBm.�C1�%fBG��g���k��Qf�祍;v�)�M.���u'-ӄ�kA����s&8��u�[�	�W`�2;a�=�հ�y���5�`�<��"#f�t���X��4i���2�	Z](	�n	^mѸ��f㲌j�l�9�$�[&%��|f�dsI�ɻX��ncPN�n#�6��˺�#k��L�V�������:R��L۫�m5��s�u�W�uH�ζٳ���!ĢbE֬�f��]nsU�! s�!j���&q��
�m�V�u���#���J3W��jLMYI���z��[v�t���z8ܹ��8�S̭)�Q��4#5��6r،����l5p��s@�v������G��]���x����HP�'�V�u�C��� �M6�l��)�]PO5ki��n�ۮ&�w	v2�ǫF�P���WT-��!�Ͳ�4E�N���;3�D�g��-��Y�$��F��~�=.���[0�a��k�r%����g"�Ä�j�XZ�xٓ��U���.yd���޽�H5�1 ��R�޽�iU�J@$(��!��3�t�:<�j*�$헏le�ݥ�h�f��� �/VU�ω�{�b�;��'N���z�����Ѧ��bN�OD����3���wn�ԛH{(�@<S��=�)��"1�������87��L"�4�����'�=3�lĀo��@$��{0xv*���m����%2l�ݘ��v����,�x˲0�]�5���{\��-N�Z��Wc�����=�;��H �츂Fܿ�ꫤ��rcZ�{*�� ���k����);����qv���=�j�1	��i����ʨ��/:�ކ^YӖ�,��������^A�6���n7����wT;Yv��+��8�FmI�Aڕ\U't$�+����q�8|I v��}��r�� ��z3x�J���Ȱp�3�(�/pI��� pw<�tV\�hZ�Х�3@$wLH�~Ps�x��!��2p��z�L�r���&�1��K���C�*H$'[%z��N��?;��A����;Y:N�˻�� �����U�fU�K��	��A$��Z�@�u���'I�����})�F]tҹ)]k3$t k�W�d��4� �i�x��P�3�[��<��4j]Wo��ۘI��@r
=Q���-�l�]	\�q �A�ւ{�M����vt�f3:�A"B5Զ�Б/���5�;=I���� �mOt�>1]��ߧ	�c-�8O�������0g*�(��9#s'`O��]�y��!:-d5N��2@ͯF���)\�����:}��:���-3G��N��`�og� A9Qh�(��{�e�����4尀N�OL�����^��Ä��j���OUuq,�k�	(�l9 �j�H�{��\�i6I�h'C�v����N��6�\�!�wd̵LL�ݘx@g�M=�H۹ِ�wdDtt��3Gc2Pb���|��*�cG[i���x��b�!���6utxW�O�\`��w"j��.��:wt��G��{�	;�;I'�����p��s1�§��c�$���쌀n*��t�"�ް뗀TUC)Ue��䎡��� ��snzdd!��p��T#ǧ��b�/�����/�l��I�����	�r Vj[���v;1�L;�� ����x%N��`�"|h�ˉa`VU;��$�>LI$�v�糙<_dZ3�IJ�^K�eQ���a�T�IL��ϑVQ�@c��T�XI)�᫴��>��[���H��uo�}p�O��ߗ(yTX��R��<X6Tp� ��O��_<C�g��b��c�#�m��=L�H;����2���a�����ל�{m������@k+m�J���.`���V��bl��i����-Ɣ4�&�֍�� �}��,�����'`�a��#:jD�E�dA#�����ݝ�0g�v\��>��A��㘼����H����Ė;}L��+�QXO�Ѳ	�ZPgp�E�3�Iw�yx�X��@2H����n�-����${;A>e���	�U�mb'wLH�s�9A��mTGI�Y�$�e�I2�>4I�=-��b�4Dn{"#�%�^������bY��cWmӂ�OD���Ҏ��냤ٕ8$\��@��$+�:dy�Zq6s�h4i�TDfk��3�Ќ���.�û��6Z�M�+wUiol�����U��S(vn���웸�\b�[{0v��/d�$0�%��pn��>9n�A�7IK>ܸ�t>��/<k��M�n
�鷋�Z����q��)�%��w�N�s�k��A�p�.6,�<��ѱ6�^��u� %��̈́5`!i��na�����3�KՑ��-�A�[y�mqQ#�;�u[4ۙ�x��Jd��,l��I)$jh��[J֮���6��9�v��V��n��G]0t�V��NvND`�@5���Ȥ�uʠ]n��ˬ��e�iG:�q ]�/�_|a�d\8A����Ȍ�$�Ʒ`9��힙]4�~m�Â�؁>e�m�ŖK�'%܇����I:��D��b4%�f�1��O���ْ@xS�z�����ǳ��H��ibz��rFgNĂ	��5.��������wy� �k�rS@53\�gp�E�3��"�D��۪�wޓ�� �u��&� �v�c��&	��4w���H��U2kb'wLg_r�%�܋�����-�XP�.����0Dξ� �A�n\b�i��0RI^ä�r���ܖ2ڕ�Uܮ�rF�)-��1,6�3T���ᨺvwp�q�p��9 �la�؟A��\A�1MI�C�{���O��vd�R. ��H�DlAc��n0�T�i���(���0���_�N�9���e�?w{�- �q�ؙ��p�ve���]��R��^7|UYg�Su�-c�F���	/I$8,��O��="@$���Mwm?Bt�qS5��.�Id�仐�#�dO�/����@2���5<
��@�U�tPБ<�q�4#fֹf	�:v`΅P,�k��Y~��\?r�(CN�а}�D��#_"u�&D3_9��|pH[�S!�R-� ���t��@�t�c׌#����SV��D1`u�P���� �w�<Yu�G���6Y��Ǌ*ٔ�n#C��D���ȂF���ഘ��^�ո|���gvX
�;L���8;��s$�A��qbB/��� tq��OZjphݸ�	;.:o�����0,�`��lM����Xs7��$��܉$���>`�s-�S��}�j�� ��_N.<R. ��X��\7D�Էa�5�ϼ�KHh�+�!������������[b.gj������2T��v�uw�Y�go���U�%�i�}�ow��j�;�<<���o����4�e��Ĥ仐��/�\��xNi&v�=�E�>($r�zr���2x/u���Ae�����L]˳x�N���y�1 @U�T�o���!�|||#�^	Ц���PF�gl�:�����_d{��(kZ̉*�p�h��f�1ԙ�֐�Ki����]�������;3�q�Ɉ �[dy�:`O��zd����Z�`�6ݡ�ѡ�� Ck^(&�m����I�˚���$�UYu�����>�j�`���"��NC�:��Y�.Uv�����f�HN]��3�(U�\ǃoc:$��5K6X�mGQ�ؐq�1��}v����i���EÄ9i�;꜈��d�x��l8e@�Iӝ2��w�:��A��8=����n�����|�����ˠz?��������~8;ɟ�Z�7nFW�c�c=����#U(�Wi��������K��H��K0tAN�܇�mz���a��u�<R��;��	9��8$<H+� �h<ɇr�~�p>z�Q��)Z�b*������ѹlp9�ּ�e�����J7k�;�［ﯗ�iݎ�H �vD	0�WY���<���>�� �]� �b�o��Q('fv�B{��m�!��x��p�s�6d�@=ݑ�Αݽ�����O9�h�(wX*�n�I�ܹ����L�I�܈#�$3k���CS��l�'B��Q�@��yon����!9gwp�8���t�/Z��r����I6'{v0O�$ ���.e��v�Jv�e
L��. ��H�v#b�-Z�w��|>��>�~ɐH4�|q ��~"�l:x8ټ��/��X����B��~;��@����c���t��fx��|��?9ޟ�r^�N�:��mK]�]݂�H):���5�`j�ٴ滑k�f�r�4�˹bv�ܼ�D��,Zf�8��#��Ý�E�kv��k�՜�ȥ�k���]��L;���)���"Y��R�\lsF�$��QƼ(�g����s������:�j����ɮ,;��)�n!s�h0A��T�b���S�J��x+,�m�)�%�*Ķ.�us��"���u烙�����۵�J���c��0)�-l2�1�P]���3�w�)ػ��w��*�d$	5� �	�v?�ǌ��1L2:dI����R.]˳{E�[�̚��2y�,��ӕ��dH'���~0H='*yz���Z��ݞ:.�� ��D�읦��ف�ݍ����K�[��5�}W�����`HK��V�g�L����d�K&�W�D�� �� �Kg>�_��j#��0ts��+���pn�E���ð,≮����|Ήom�V{����4i��q��%�zd�8tOt�$	� ��Ȃ�<����n�����G]��f�8��D���}�, �]�k��BE��!x�O��vd�1�O[FN�=oq �C^=��(7*�%;<I�k�A	���͈�g
mY��|��\�/�j���p�-����7�p0��|�l�M(/�,L0��s�/N�=�x���LXIan7��c=��4��B�y����H_dFsc����w��b(�w.��L�6Ǒ&�NtD�XT�Kh����k���>%ĝޙ ��rH�t�A�v�;d�6��9DnU-���I�=GH�Ov��"�騰�����<Ot�&�$�;�3ckvN�� k6�D��hN��d��9��^U9�2���x�6OU�Hj��o�hĳe�M),��&�ہ*ۭn��G	�i�&fg~��Ȼ3��v�wz��`G�36�C��������d��#y��	^�oP�����8"���
��gf����y]�cg��	>'�/�A@��AeU����?DY0u`��Q)ٓ��3�Ț_u��*ͩ��vL�*�4�1H�{0v�e��>�r�\��Ƕ�����)�x{޹j�.m+���pJ���R��� `��P��ЀD�{���}������=�o��1����<wY-�{���TĻ���?���SQӾ6�*a�"��'n���ۉ�&!�P���������o���k>뮨�h�꾜�ǯ�c��{m���6�M�io�����+�T�jz��[��9h��у۔!L�	��nѳ��"Tn1�t��M)�wA�.����C���6n�SF�A��y�]0��y��c<xNҕÍ��l�\��ؠ�Wq3����e^��%��{����;��(v�5M̾>b&�3,�t�-e�'Ab��	qy>ů<"���s� ���^�j����8�bF�~�W/�&����D_����:��rq�~=w}�A^��E��X�[�7ٯҗ���:]y�^[�A ='�&{]^�%ȡ����j<���l�o���zW�z�o�m��}퇞�|��.=�c��a�M9�Φ{��q���i՗����ۺ��\/�A*���[���7}��ol\�n��%�G48� ���P�̼�ǪV�B쌇�=�U�S8������||1<^�/bze�*ͳo��"V�S=<�ug�ڼ�Kq��D��Vl��Owm^�M��򪌿c���~�����Wt'��7{���?xh����rJ'a~�6H��~>�<��d%{lh~�y���Ds�}�=����2�z�\�ݜ65oql�>^������BL�W�^1�LM!*ȑ\�)�ّZѣ�U��)���y��8���/3H0qD��_�i�)�̌V�c$�T��Ń�ZŮF5��/HCM<:p8"i&*�BZw6�QQ�¦Ř��H�2L`�����ڸ�7>x||oS�"g-1k-**�r��D��pr�9Y���M�hTd|hJ�/e�Ӈ�K��+���eb�20�)!>��5��d���GaER0fH+&,$
��>���p��o6ȓ��*)�B��w��TdqNʕg���m�>��n� �"m �ԘI�X�s𐦞��E�h���\Q$f0H9��g}����|�_6se�����,�q�O�&"�=xxt�p^21�	��*��%�+�-�?C[��HȈ��qq�̊��S��ٍQQ
��B�:o^I����X�&��gy^�Q\S�xk�H;	��*���H�?�E��z�p��j<�DQDqjT���dX2<��u��b�d���H(ɐDT��� (�&8��e2���_��5��2
�}���H�js�AЈgwN�8bfA�MO���,��	uS�>$fK<x�A��yD]�U�Ñ{�zZ�I��U��d��������@�AQ�!EV��3ۼ#��>$fK����o��Y}~?F;�p7\nX+k�kl\ge�5uՍ�,�ڞ�d���H��e�|�)�=�.�g�<�F�d�$��I���./.�7L]��-�6fv��f�RvL��;��,h�Wmh�1��/��'��3Qd�z�b��$o��<��we��e��G��r0"����b-�@#n: ��a�hbdwY�zņ�r�"�3g�A!L��%'b�y��=��\=�g�B�~Ȃ�9o� Dv�Keԧ؈��r;o��F���|��6�H���w�SZ�R�ѥ0�C���Mv�e �·���Zц-���ʱ8��`x
�׀� E'�!��;�`��Ȃ�OllH9s�h뇂j9��^�;��KM��9ѭ��~7���f�M�9�78�Cgr\mP��O��.|�╼ae��L�N����*L����3{:"A$^���B7�&|Z���İ��p [�o ��JM�33��&�6�`6�Z2�!��q�lsǉ��N^�W�%@97Sɺ⯴��2��vZt���9p��ٓ�0�|b�$��տs<��1����j�X8&{�06�C�X8A����L��GHk�*�Q� �Օ�&���I'������&0yT�G�$��K�Iؿ��g��:D�A��DC�h+�4ԓ���$���>$�u��3����eG`�
�ӗ�Ć`�OV�Ynl���z��;=�b6����J_?=�C`T���M��}�S����1�3�R��#�)��)S3q���0�h{ԓ���G��63ȯP����91m\˹�cM��f��k Xֆ��k�v9�k�7������>��GlG3a�:����fbc2�]�ԘK��<�s[u�X��V1����i�c�WSb[��`�u�4+m��ptŇ�, r�ΰt�6��&�n��F�V6�����Dy�1�e"EF�bKy���	vSq�m�7���C� a��4��vt�'�V|���Q��<H$�츀]��v�LJ���&�@A��y�ȟ\5k� �;K	��q���^�s`�Y\�p0>��̙ ���C�ռ��]�O,$`ܰU$�39N«6s&A͸�H5]����n6w��WcȒN�\>���Ӧ�;��.�n��l��+Kv��$���I��@lm�X_^S0������ʐHT�<`�1!�X=���}�C�A����6��j��F�����ګ��"�nvV��*�p�P�R���h��N"5�-��u>hu�s����Pg,��Z��ä
t_��9��k�wCÄ�o!��h��8E�d�Ow\A;�M�C;:t��ڛ�1we*�9�~�-�
�/[0�)���*�n�u	�\ZP;���}���{�A����>Bt�Zޤm��3גb�jr�;�5�RR��d��f�p��}[��cw($���y��6l �uox�X`]$�j�gz}
	�أăw�ݺ��9�n�ϻ�� �@�w('�$��*�l��'awwՓ��'��־[� �zb���\�,�g�8x�JyG(8��홝�4���-#3ĕ]Q� d𶐁g.�3�F�u@A �v�H:*go3U�#�qq � �-v����oL�W�R�:���d� ��c������mn
gJqΈp5����y��C��W��8�.����{�³A�����u�R%�_�h����쪓LXb����������6B��K�
t_�b��I��zZ��k{�̘�V�f휠�O�;:dJ��Xc�#2r�b�0CD1�d�D3��A=P-J����������ECҪ
f�*q�7%#��F�e<�@Q�ZI��X���ȹ�6=ޒQ�>J��� n�?-y ����<��J���\3#�(��Ccȴ�mڄ�������0.�r���WD��Ŋ4w8=@�-&	9S�	 ��Қ�$g�#a�/8H�~0>��T��3�N��@F�d�A�ف���;;3t0��`|n�rD�{�_0mƛ����.�;I����r火1v��(mm�n����1]��c�s� �P�WYϟ�C�%��m0�﷿�?:�8Km�bA �N�LG�=�N�� i�l:d$n�zd����\�"�8dK�
4�q�<g���q�uO��(u�m��"<W�X&d1`��0̌�m����0�����p��'�I'7�A+R�nQ�.��܍ӄ�H����AI]��M���'Q�;:t��n~��</�Q�`~���S�	�}�x$�O�i������j����S49U�SW��76��]^X��룎��z���s�����Ϯ{��>>G7P�s���Aw��c	���M���<:�8�[��2H6����t���F�\0L5sd��7s��[?O{	�yɐI ��ǣ�5k�ꇗ7���w�bM��)�JY���`���:�f����a�Mu��6rTCo}�)�ێ+�.ù�r�ĀI�ʈ>$�կ� 0�oL�WA�w�3��"|h��x6H ��w��L��.����U��mv�E�m.�F�'͍ؠ�A���"�3�[; �C͵i��łpȗj%t>@�H�_@b ��WT.�Gp�پ�A&�*!�^�!SokM�	���P(�5�TFNu�8˯����<@"S�5� �ۮ��[�/�zZ�Z&.� �|M��v.�'����>&�k`d�{���Q��������!�^�m�D��3Ί"�9=D��*B���9<�ݨq�V4-���%��{���h�3`0T�Vo/s��X�w������X�������o��������n<�
��:�d7P:��&�:��Z��2Ljܮ�8��b^��גj�ۻn�̛\��Ud%�����`�0q�(d-�ۗF�ї�L�����p��ږ�[�f�*���g����x�1a�7��{E��Ae;����-�]bٰ ���uv,�k��X G;dwnF1�Q�N׷�מ��;��FnWT�z��J(�$�H� 5F��C'j�����kk[S"���b#��N��ߕ و\���Lz$�ca�	�`�n��k�δ�(�dP]4C�tH>[܅$��u��c!��ذ���ܪ�%���!T�`A��'��	$w]t��F��І�����<���b-��-��jz\X���c��ٟI�ג�o��wt$�_<B���Xb�8dK��=s*��&{��	'�U�2	v�31Ω� �uof	��)X;�A"��ީi���(,�Zȇm7cX]|���!�#e��7��<�b4�*]"���'��\6����m�CvA�p��pd���x��%�sc��5{�=���,rma��W���>4W������o(;efC���\��>$OnDx��#8[���	�P5�1�<����Cs�N&��n��2 ��1;�����w�Pxp�m�{Ud�-/f��ǡ�=�R\�����A�;;/�YpH����x�V��LDCm.���
�u�ȃ���L�9�I�9�f�㠗�
9L��d��۴��A'�* ��Bkm�@}iS�A"��#ē����:O�BA���3���u<w3n��h&��A�~H!U�@$�˷�����:��"����d�ui��őp�K�
AsƼ�܀�YhC���P|@窀����q v�G�i�������]J|E�~��ن�sq\<,!���1�0�-�[�f]5�e���{�y/v̒.����{�Ąu���dr�̿\���m�. |k�� �4Y:���g�:8Ccd��W��Gi3���z���̨�	wC�mm�2a~}�}��)�LAr\��";���Ư��$�X�z�_���v�<�1d����D>x�>���4���eQf�������j �A�M�}�v�����+��i�����᜽
Thp�;[�6q�m��;�ѩwX+U3.�ӄ(U�r��۳��B_����h���A!�f�ϑ'�{�q�;eW�O<�'X% ����ύ����s�Rx���S��	{c�#B@�Z ��n�d��^��y�L,��KəQ�<�h�˯kq��=msU��q�멐������P4R]��������6@rI��x/����z�s��	eY� 6A��6�����3�� �%�z^�G*����I�,�1������m�$���nӾ�B��{� F8�!����E�{��p%����3,L:���.sN���c���ވ �~�LBb��i���R�L��x�(��z�qBP���Mm�7�g��V:+��l��\���C�)d0���k̡C�8ͺ�%��[��t^�d}l׈�VЪ��Z�A�xHB�v���I��3�����v���ި�i9������9�p�q���/���#^� I��~�J:�c�V�s����@ɴmZyĈF;+آ��nJ�ϋ]���]���"��_<����Q]����,J2�fk��	�D.�ȸ6i7sA ���H��Z�F1b���P<� �Е�y℈7;b	:sT�FH�>�����j$`n�7���U�]�D�ΨA>4�s��ik4�9}-`/M��K���%0�.�Ar��3�G��7^��� �IDÈ��O�	-�f��z]�e�@.)��#�U��Aw(�n`��P�H0���E����S֏ H����5�~-u��ߧw�z?o�����~�O�E���_����>�(V�������vM��ll٘5B���j��5UCR0j��R��`�#��+�w��:D`Č[��Q2��0j��B0j��I���2#�e�b����5�+0bF��;vjC��MR�#��2��+EX2��EXl;t�tUۨ��
�ٱ��V�f�f�R��jU��͖��a��VJ���U��&R�v�.���Vf[*�ų)X�l�U�͍�͚*��͖��ccfƊ�e�k4��Y�f�Y��3��W]Y��[6j���J&%Q���;��} ��I["ֿo��?���{O����������\�����Ο��_��7ݿ׷g�u�����w��_���TQ*�?��������J���*%_���y}R��~�?���꾋���U�_���K��ƾ/?���/���������}{��e%%fE��j���i�V�VY*֔�e+YJ�kT��+i�@V�#iB6�6-��*�)Y�+5J�R��Xҕ�%c
��V�J�i�Z�Ve+XU��cEZ4��T�YJ�IZe+K�e+Q��J��V���Z�`�VF�X�J�i+ej��¬���e+Q���R��Jڥb�+e�Xe+S)Ze+R��I]*�T��w����w�}�a��J�)�)�߱�Ou���[\�>��y_����~��Q*��ë�����v�]�����͞_#���QD��^��_y��_'��j�J�(�U�/��=��W��W�(�qe��~Bg��Æ\I��s�6O��?��9�7)�f�Q*�g����}eJ����K���o���~C�>W�Z�c�u��%_o��D��o�޻[E�~��طW�_���������?+����W��ͮ_CK�/s��~���=/u�QD���]�W�Q*�o�>����K����
�2��.� )b� ���9�>�#�.                  ��h        � @   �^  ��� 4h@R����JCZ

P @��$ �  � �� RR� 4 |                                     EJ(   @  )Jw@�T�3j��f�` a�2@;�@���4` `f1QL�T�� �: )F]���S P̀���jT�����U({/ �%C!�϶�B�A��U^f���^0^`:�
��"E�         �*�T+ �*�73�J绑OҊO���W�Ԩ(u�� ��(�%*��aм�:}u�3TQK�i�d	
�p 8h 3 \��P�U)@N ����� � `!�U�
g��K� s� ��v�d4^�s�\@Q �           u�+f��u��U8���2�Ҫ�^� g�.fs���u5��Ì�*N� ��/cs��`����ѐ�J��   9�y�ꕵj��*� A��v���&�kj��=^��7l+�{�zқ��*V�-�T��˥Y�,�j��DJ��Q^   �        ��+m������D��ͤ+��y��N ����r�N!��2��jv���IN� �jPr7&l˘g	M���  9W��N���"�� ���Ә�͒q�s�tMYst��u� ��T���P��Z��u��3�n���P  ^  �         =�����H�b\Z.']5f��:�,� �l�=�9�m��X"$�0�W�㴡K�� �);$����x���;t r 4` @���@ɡ@�T� k   d��`F ��CAJT� ��JJ� 4ha"Fh�j  ��U&eJ��   j���T�A�F�i"jz)J���`NO�������� Tkϩ��cE<vι�$ I=�3���$ I4 �H@��H@��B�"BE�~x�#���_��'OQZw��l�[0-������Y�*�;;�5�>q��T�MyЌ��l�VN�T�k��B����,�pjbb�s[*�����~�A�bg;{��Z��`����� �u��7w^ռ�t�jbrGD�������o� �Ws���,�ܠ�7��
��p��f�}����:���-CR(`�m�ˏ���	9��i�k=Э W����9�B¥��J�3�=��3`	�.�q�ul��\Ԯ"��w�	lXQ�:3�q!\QY��D�q������Z�����E�BO!���/
Fjk�y椬N�K��@�_̮��kݒ�`�3^^)d��[iW�b�OQ�LӵK�wA9�X0��+#�^Jd%���{�!4�lYk�/4&�u���h�!�;*�pY[�KzG6(��p+�k�k�3�ΐ+�P3v>)j� 6J���B����4I�D��wW<���@�V�q��q�ʖ�͠$�on�a�_Zv�W��,��N�yJ�i�k��!)Z��T<\�(�mcr��Ē���A��q�D�u.) k�j�	�q� �v��,�z�q]�7�p-
�誳�- ���gL�Ҕ6�n��(�u���$�Z�5��}���3or�T�̚-\��3�Fz����ነ9���5��-Uj2��# �%���O������y�i��m`��V��NTtLK|��g�s�ӫ�u�}����4����nezzd���vN�ⵞ��Y��G���Y����oJ<�|����J�n[k�K���
@��;�Xͬrg��2i�3L��P�������.h�8e[�t�h��9��κ2�����sAǔ��l<0v�`Ft�:u6���Q.���u�W[��Mv53ka��K��o��c�׫��Hte�vA�lRG�QSv���۳j�Q�K�B�ո���gyv$8�Že������@�;�r5�+x�ï�D�]��u���q�J�{�	X��u��5����N���j%g.ط��z{�F��s�o ��;wR�yn�^]��ksx��\� 2���)h\ɫ7�h}�P)�#�E"4Z�EF����\�>Nb�{���\��x�ݝ�z�)�<�6n�u'FV��0p��_�����4n��I�(��hW��S�^��md���sQ�]��I�"��	��G��[��ň��,՗��!o���7���8��G�`��K�HvZ�	e�^ � Dû�C�0�	���S%!e٢m�M��_ћ�;X��H*t9�Ώ#��o]����R׸-7�'֜Yv=�m^���QυbW F�ν;�]3v�a'�n�P�zn�a3o=>�A(X9F�lڈy�����f���dZ�on����r	�����K����±5�Jq�Y�4��`}Ǝ٪��M��w��ͬ:�X.���cJf��Ɉ&h��;Ǜ^l9�i�����c���FPq�E��фם���L�t���\�ICu��\Qש����ʓ�f�7��i3�IHO����t˫��g���2�)wF<nη�,��Wb]��J�k�!�xjѹ����E���դ.�D�,���c���4��o)�J{�A{���.x�/��y�^Z �t�#���d׹QÅ�GB�t�㐜�˞'������6�xk��|����Gt��m�1 `�wd	����C���$�����^�vG��z�hYz^��[�N��y��ݝ��B8�Nք�P��)l[P@l��ڬ�(3��q�D%9�ڕ췛��S�x;yΜ�{V�0��t|p�a+�r̛��5���h˫_b�#{S�zt�z�;Nާww3f��6����҂֢v���o|#���dv�tM}��J%+�h� w��%R�v�D�%��P,oR˘�Qػ�,ook:��'�~/��Y�J�o�����!˛R�UJ�������$�Z�8o �8�oQ�3wuA������c���έ�=�(���P��C�K����gm8/]�I��:����׸�o�c�Y�9L[����Kp����.S��J�.]�gl�Ӣӓ��L�w���WGDӃdktӣ�ۑ#�hD�Z����iI�dӌ��C��yu�ꡫ������ ��A6r/p;������5&p����+�]A_=�	X7�/��w����]��U�-�!9T*����v�6�.��B4���mPJ�w ��I��Ϋ����u�X�$<���=݈Y������CN�ћ�cť��D����B�N؆�jUvf�y�7��yd�ɕ���v���V�>^;����r0�Q����ۋ/Qr·Nu[J蛫�!��F_��k֨�49]8.5��R�2����\��|8]��˜���K�� ��k@Q�h$���ʜ���S��	P$-H.o=y%Vĸ�竨KtYr\�(u(Y��E�~���0�itB�����b͎P�]��Ƕ>gf�_a�)凶G�O�+�H�����w7��\�~�u±��)X�:���g8c�B�#�o%���9�ڹ�6��UEWac��ŏ7xf�1�O;'v;��(ZF�CtV�,u�Lڨy���U�h�c�oUE)��ҧl<�u�
�n��!��g�n4�E�&�7����	�Y5��Z�{��1X37]�t+��� ��\�ݖX����I�fۄ�ƭ��Kz5��D�v"�F/�H�j�(�V�we�>���E�{����yYp��m��t���{8�3�z:P�/�Փ���� ��:;�F��4��:7pN��m՝� vkS�N��c9q��Q���Łr3;���%�������Bw��W���D"N�zÂ��呜�j�gE�}��[0wo{�(>ʝ�y=��Q�V��d��5�^p�otgd˷�n���b��!�;MX$Yw��ٸu�	�83y��>']���;���������ʌ���ֺ���,\t;2��qzVq��e��4�sKD��<�[��4��r��;U
%{7Z�_�����m}�v*vsO�6��{9]D�坒-�g�Uܸ�;.��L�L��̷C�Ѯ\ �5�)��5���K���Bv�IN�Gp��&��k�(�_R��B�MW��.�8�TojFt]s��wT�S���@P�7�zmut����0v�&�6(�Nw;��mPb2����nm'�AO4a].qpۊ��x�h�;Q�^�`OU=�a�&�VY�a�� M���Tv<L�)���SS��"�����W�V��Q\qa-Q�:g,8'.�,�a4
�`��[��oO	0�K���I�c%Ih`��l��g���pb9B�����6�׼���}J�s���/f�WM��n�8����c�KF���Z�É�^G������t�������3�>�,鴮��{M�iY��� H#y0��o6�^�*�6owoHTQ����N�to�;���9bX!�Y�γ�:��܅�4󻶞ֆC���5��ލ\�EZ~&e�n�$2n�)��t�����J�����q�)�]Ǆ;�N�h��*�N�:'�>]ת�F˧��𭕲!�|f�Pc��ƞ�����@��@���>\q�o�?N�l~O��7zU�wKĢ��P{uS�f��G9��Vw+0�`�E}��7$̙�n�����S��u�M��1�M��wc��Dt홝I��Z�a�����f'v�n$��a0��c�\�5����x.���y>��=;@7��,gVΝ�����ozƻ�~��'O4Ǽa��ݜO�~�[�S$�:WoPl�d[b�8vĠ+y`���`����*g^����{�kb�r�L�s��w1�z7q�0�&��TA��i���(�u\�o=�yy�4ftt�46��{��M*;�Gf��N��������܇W#��Z���>?�T`g�&mp�4�ܙ�7�x��ӵw}��f�D�<����!J,ق�t��8![���O��Æ��t�������Ϝ�u�����l���vN��!*Lp���Nq�[y&��u�Y:� ���@.�y
O�m�j���Q1�Z�}���t��u#�$�.��D&+e)� �A�K�Dsi�s�,j�ɺ���#�Ezlmc�3�=���^�&�����E63c�nۏ �x�lGg�)2�V�X5%��!���B3�hݝ�F�L�^Qy]�;���2l��Ǳ�����<u�mQ��-቞X��X�w�Q���]!�t���x�3^rRя�Nɨ�	��FoK���fW�b<��7�8v��.��9H�����f���{�&���*F�e2Ir縳��Ðj��c�nи��=�*�����#&��l��6�ޣ�M�������Wve���t�xUe���r��t{���{�;z<�By�nQ�Q/��Z�h�EC�|l�m;��8b�܂�Dl�gp#6l<.�9ʡ��h���nv4�uY�� A��c�����Y�&���]�^
U|f-ђh����ױw���3�1�hG3l�A�2+3�A��zw�3f8����� ��hGY�K��W[�.q��m�T�T�[3�h�F�k�s���:��غ��6�uu�Zj���ؾ�r��VnwZ�
�pmMc�f��`Õ�Osͱ�PI�W�^;�%;J��I�&�3l�k���83��mh����"��×�)ժ�w�W`��\d�m�Z5J7۱��|g����{� Xr�vh��|@�3y�*�6�@Mr�D���Rol��kDr�e%�"j�댶5m�j�p�����4�O��Q�m���ym������5�:p�8�������A�S��%Sغ����>%�=';�(��������ר���8����jۦ�N��[~�h����(���M�Z+8�v�v���y��L�קpU�Kt�Ȧ��r����;��v�r�{���R�*'RN�h	�;���`S7]ov�˹�Y�bR؍����N�D��%��PP2�'��t�3�컻s�����N�%=�����݉c�,�pQ�&s�Mw�tA^
j
�^�ɷ7#�zusB�W|�7���[����vf�[�t�7ս�A �jd�i�=SNR�ib����Z�r2��Ε���w|Q��sc�L���O��@C��	pyq� YTY��c��!��;ti�.��[Ԃ_I�P�,�Ʋ'�~��T�e�-���Ҟ�q�Sk�'	�}Jd
KsVn�-�Yr{Fm�:�I�qh`���ݛ�K\�W;7��G��C(�7'֞#v�MV�nU���b�����۴��ҹ�u�M�*H��@E�D�;FE�m���g�Bf��f2��
{�Լ�#9}�����>��#�-#�7v���B������^*�Y�f�ȣK ���jk��2�޹���`꣜˳�����1T��/)*t�p�w�G�iY�`��h�4�v\���3Q��5ohf�[�r��V6�w�쭜j����3y݌��L��������#Wq�07c�5
�����^ǥ�B�gQ�*0c2#@v���s[�9��c|��.��5������ѽwK��.0�oU����3>���i9h8M%-�WF0;�LT��*[��
�[.)4-Ü��9�LLmDGv޺l{�_G2���#���60I�b���k7o1�\|����[h��j����s7�R�-����(�u|y7��2Cxm�fo^M� �n���v��1�M�ܽ]�ɝ'~�q�r�ގ�%��BR�@v�_pӶv����:B�^���ڻ$�臩�n�@j�{!+w��.�Mr�܋��5^+T��U��pS�n�>͓[��;85���q����St`�f������k�=NEvٮ��t����|�8��Ü�X�GQ[U,� �V��Mr�f��M�{r/�w�v-��Y�W^�	�NN]i�%�,�����/cC���<F�̃ٱ��c�U��u�*��(695�8�_��Ծ����l[���FsjMvZ���&1�u�0j����⺀ۼ�2�yo]�&�����Ɂ��"`�h۪ȇ$@p@��˓(*7�:��=��i x0&�ok(X��Nv=V>X+ ̯�yӶt�9nI*�c�^�?a�S.�Z�Z9�ūv��;�r'�A�����s{����%�֨|k=x㍒���q��m����{[׊���c��.��r�\ZVǔ@��ݶ��q�
Jݜ�A3X��;�����5��2��2���{�*[ KC�&�G�oaVi�eK��࣐�Z�gt�{V�8)}{b�7pLppQջ�u[�d�{7��3�O�:�p�-��:f]����摅�5����L�p3��o9F�Y\ӽ�9^F�	�gEŶޥ�4M�1;����#w���,y7��K.-�Q���^���;V�J
���I��vgh�wqһB}�݄�K��i�f1�����IA�6���x P�W�+1�tѐ�1vAu9b٪�*�!4*�P�0�uo�l�u��<����=��$��E$�����B�BBB,@ ( � `, T�Ha	R@+a XRH@Y 
"�+"��R
�)$��VBE�E�J��!$� ��E� �I ,�E!$R@�� J�BB�
� T�%BB(HE!B(@!�X, �H)$X"�BV�d��d��!$(I!!!�!E�	P$�IE��!
�V �$$X@�d�I�!"��	 �!@a ���Ed�"���HJ�%BJ����@�! �H �AH�@ XX��J�B�I ��D��RBB��מϳ�E�e��9��ŷ��s+tj򰌭2,Ц��f��Τ��3r�_�h���=s����/E�42�M�*��\f��� �oN����7},���0��h?��O{C���p����M�yd~�W��>�D�����'�����Ӽ�����ʧ�垯�D��ޱ�q�i�IQ
��PT�N�y�ֽ�0^�L�ɝcbE6o7r7C�K#Զ"��)f�A��ascpc�����T��{P��ݚ*��{vo{�&�_���b�Qw��xM��ʯ+p�ظ3���9� %�7�9��B�{��(o��Nۻ�Y��������=���\��W�N$�EV��܈����F#F��4��ۧĖz�d��Hd�Q��	&#�j����h�j���:o�'�wi���ji���M�}�$ֺc�Zx_�Ҳo�~;�:����o������q�𷧐���V�&���K����5�-�1G�d9�ҥ�vz�p~����}�6��v�.z�L�=HI;�nlO�������ؗh�g?Q��
��q,݉�H^�����'�ۛ�i��0�d��eLߙN6�)���O��۷S�=��]'���&����!�{ǖ�M��l,Q�BÈ�8�އ�g��{���SD­u{�zf��df-̜ܵ�kr�԰�ӻ�N�N�����zG=Ni�/ޚ����zl�?�ﳲh�|�ƚ���8��,�b} +���y{�s��{~;�H��7�n�䜫�y{<�OS���{���Nj�fV��2+�<<�\�Oݨ�_%Q$��j�ۅ��}��碄{6�G]�}�#�>;����<��c��ճo��Ӱ&,�Axx5+Ó��+��훴��x�������^�����n-�/�SEL.�3xm�ٞ>۫f��㋆�7��f���d"kD=��7�9��S��>F٥�ʂ�WUti�ׂ�nO52�<�B���\3GK�_yi�Y��5�*�o�q��X��L�A�����f��{�%-6 qQ��=�j�;
�x��g������Ob�v�uX�ŋ��>W�;do�s�e�R�>��>W{�p���xU��cQ�mAvY��6-9��]o=���Oxxn�����9ЖF6yE����_��/�(���8{�'Y�֋�Md��E�:*�lP����>y/p�g!<G�6������P��ԓ��&���Z���(�=�ݍ{�7���3�Ƹ�>n��_C��_Y������@Mz��+w���{�s�z
|�F8:�6���֡#+f7t�m������p�e^�.�������t��Wu�{n�H=��导����Iwp�Q��r�5�Cۺ%����M�G���X(͈���'�w��e�z����y���y�2ʨ��6�ٲ!�ў#�f���v9��Xg�G�p�;�.�޺�UMgrF��~��vwhpny����1[��"�݊��n��57�$=ء/gY�j3i�����4���p�:%���{*W�+��l�.���7N���p�W�1\E���w{��.��V��t�����)g|���s����(nwC<d�.��H/���7��#2��qgk�}�J��l�T!5��������<��@�4���3�${���Z�z�ӫ�7��L�zF��)�l@z�N�צg�����M�V�5����nw���7�d���}�;������@��묏g��A�٧f�l��kF�i\��-�.���B��z-���F���aݱ�3�;Õ^O=h<11:�L$��ﺝ�hT�����㈮�Y��C��u^H@lW�[l 5��{�
=@k���W۲�Vku*���CbZ�I�l�����\"�ڶ&
)h�X�ȣ�i�fq���xrj+�x	��]�x�e����x�E��f2I7������n�]���ku�U��Ѓ&�2��á�o�
��Z�94w�����'\fPѦ��0cci0���Mn����aᣠ�|�^����{�!|��O�l��|4��MO��z{m��1��-CƯ+޼������=�\��Q�Z�ÿy=f{¿4Y�� ���}�/&o��E��$c�j���q�v��}$W��'e����!͡.�g���M�.;P�z�!	I�t�eR��3�W���ı	V�f�?��]:M6���'2�U�4G=���� >+�'*��.�C/�t>�L�mk{v�blFY��CM����Q���3%Lm�O@kӏo���!�Heg=q�b�p�׫w�>Y���~Y����A�$����?Y�g)O�[�9�\ vd��ԗW�z_n)��e�2iY{��ף�ټ���*�@���Z$^����v}Խ�zW��/�p���t7���͈F�d�!ha�E��{m�H���R�mj�5����n���ą0��;M��%8��2����S��n���7�E��Z� �w{�O�\')����߲���{�R�*9�z
�	��ּ�;�ڢoWz�`��Ojǐ�����<�|ޙ9�-Z2Fኙ^�q�¼�UѕN��4�͉L�7�6����BV��6F��L�'v\�UF��B��;f�@}��Y\��>7ٿ��^l~d�i��~շvr�G��O}����?){ HC�f����>���V|�qx�%�����=g�uɺn�����mec���-�n\�۩sTv���'kr�g��@�o`_ ����|�*�
Om��xl]���K����o��Y���o�)9�.[�S2N�)�/C���9t�v�l�
�ǵ�u��ׂe<�h+�{��h�0e3���L����w*����+�u�?Y�On�:ó{��ˊ��"��vv��^\Ϧ��pSo�>`n�4�i���|��l#�!�]f�'oc�%~�6���5�w==�o��>�M�_sr]ȓ�U���Y�+���a�����:��,^t��C]n_��#/n�.�%�\9�6	�ݹ.װ������:u�����B�Ѿ��z� z5�kħ�\	��>>��,k��5��9�|$&v������U�H�N=�K�+�Ut���ռ��5��3}J<��@�F��S����>x{�p�p[F�͟D<-ݚ=�m�����A������w��X���r��_���L�pwvA��/^}���e o���ݗr{���-Ȝo�,�Ȼ�S�����u���(W�|�{I�zĳڽ�,�~~���]�ղ�$W��Kn����Ѕ>����vii�6�垷�&���B���ɜ�ٷ^)��<.Ƒ�#��u��|�.y���V����g[�-m�u
q��}�%��p]��v-<�Y��X^�W�9��.�[�2��Y8͗�=�����<N�����5��H�j���çd!�Oz���k���z�|'S_a���==��k���V����$�n���:y�=6�C��=u��;���v=�6l�H�^y��.��CR�^O�'��7�h$��g0��y���w��᯹�y��_ޖ�=y<��w������y�!���G��k�����GQ~~9�Xjw����gȈ�^��D���s��=��G'@�-�LT�[�P,騇��ܙ�m�;��{��(峐��(u�izo
rtM�~�/��_���������㌚|;��<�5�N��u�Z�W�ι�����վ�q�*���ww���F���lo{�>qf�Z=�L��ۅ�Z�,��n��i�Y<�&�]��������0�2��mhĈ��c��>�`��
����9�C�q[ �<�hR���g�}��� _�Wj�<�w�u�Q6��4�U�;����s#N+������o	���4e�>�v���öG[�|���9ǙK��K_����xz�컅�2��[V,]9�Y>Y$�.c�,����%b��2g�x�����o�LK8��<�y��=#z��qD��6��F��"e���<�td��!����;��[6e6%�̻S=�X^;°�ٳ��js����۪��&�m蓮0Q�A�Ū��F��Etg��{J�i�?z�q�}�A{�Ga�r#���Eb'[� �Ə�����j��l�^��<��z{�,ͺ���E���.W�(DA�T�Z���Z���ᄫ��`��//S7rι��*�Z�!{��Z�!Ы���&s�Z��"���È�0�u�^>~��Y�vg?4Ӌ��1�������1��;��*���_!�iʛ
?]������Ef���]u�}������l+�)�>�#�wov�����/�ĝ��C�H��FV�v��Dw����C�.�yM�eCgi��|CEz87;B�wY��ܷd���+��Ik�`���z��bZ���_iH�Y�b��H�R��>!w���J��͔0�����9�w_�ѐVD�:}�q�R����^7櫚Ma^ֱnU��K� @N�|�����E�GAE��>^B�։�ݛ{�[$�f�^�E�MD�,=c}��yFe����幼b~n?x�8��A����n"�~҂�T�/І/U��-M>�ܴ���q<���K���Z���W�f��#<us~�^!h�e\O^��:�������r`<���::x���V����_K����t��(�7�I�y�����QG��< �&k��{�2E�>�7IH�z������Gצt>gm¢�;��/v�λ�`�U�����g��zm���-z�����E�ݓ��k����W��+�5)3�q馯?3�����o��s|A����b��Љ�9��ot�(f�a���XA�o��O\��;(��@���icc�:5;�!=?2,�,�[�{����ᳳA®��Ol}1o>&���kd������pk�&�޻��A�8)��5��Jf�<Ta9�8���	V�?n'ఔrg��\�A2<n�N��]���Ɯ�	��u�[)$M7޷Q����:�kV�6�sV�Ka��R���ΑFj¥�z���ީ��^���;����p�-�Ùּ�!�;�����^��>�7|n�>VwL�O.�:�gr:��.>psz��lô���e ����{^���Z���ڻ�v���w���f��}y53^��F��}�nm�7ξ�4�ើje�o�w�'��,�>�+ޅ�h�٦�r�����ؖ70kq��B�x�7�b˦���3�R����^�����螥��U��'����oz���K!�)q>g�Ü����V1����2�:���[��-<D���^�@�9����z�7�MW�>�gUnMN�eF�#jRS����{��,U�]'6ݳ3[�V'.�ƫʆ��f���FS��L"��(N�'q\�&.蚠��)�͡�FN�.�p����iLY���z�oO`}�(@�L���%�w�|�K{/���^�d�~xg5Q�^['y��\�wދ��v�6k��.[$1�s}�^��-��?��xH,���(�}^篾ӊo����\ݝWz֡�+��rg^��ҊG�Y�F(�����$��p@���G6� 1���^3xE��:��/xZ˻�w�Ҩ��Z��ۃH���V��sƌ�A_��<��C}�&?�5�7����_xA�a��c�͢ｴ�.����w�{�A�b�bɾ��O�{k�U]������t�i�7F0��_��A��4joНD�E�-��7�TxW���C�"�5q�K�E�9��.
�ۜ���n��Ƚ̇�X��P�S��`=��)�٤����Q�ў�^�����7{�jO����V�͗ %f���}gC�8.������¦O	R�mܞ��<:y��,��C�`͵0gDN�����5RU�zgPv*���x���of[9����=��?2�X�Ԡ���'Z�+x���l1a�F��.�w��3�Ćj%�6{m�d��}�4�:��~�y��}T��v���4g��	���{YE�k��90m�ӝE<��QS�z+�n���Y�[��O�!���Zt�h�^��^��%�4���M�lr�P���]D:������ې�U+��t�}1��|߼���XH�%D{ę�2eۧ�R�7t��l�,Wn��7ki^%�P�c|���י�� <�����3�(��$�g�1;�s�+�7H^�|�b���SG��+s(j2^���v�]0w�%�ذ�lZ��]��Ξ��ΜWj~ل{����*2�c�[���G�xn7x�8�/{l\C��n�n����s�x�����=��y�z{�
����
_gx��y����r���R��32o��ڇ��Bdy���F��N8<�������{�l>���[�(�˄xy���R(龕�/���6�7&�}���ٰ��c3�-�Ӎ�!꺩͂�D:x�U�M�5��-�:d����/Fޒ^����9.�k���������#��W�k����7'�Ia�~�������N�aXG�^����|�p�H;:���������s��O;��Χ���Cv�˽�6z��eSQ�vTt7�ޜ�~y=��z価�G�6�`��+�����؄���w{=�_\��z@z?��y۾��*���>щxU�@sa޺9TK���(���Jי�J7
d�����:L���m�^ASz��zIv$���wbWO5�Oa�����n;H8+��>�|9�����+�� �O<�];��N����9K?5eS/�\�~��ɑV|N��}�V^ԍ�W66�=�ᧃ�4q�0��r�����F)�\�����-�7�vi��?O�����]��ׂ��j��N���|��{��[`x#L�E��/`�O�Eꮯ<�{��o�s����INI7���������AS�u���Nl�nuu;�آ�+�p�q&�x��獞+��^Ws� cg�[�.�{�(�n��œ0�FN��^�����=�j�i�q˞�^���F���e%�˔�nkoDWg\a��{V�!�V{9�mF��1�Tn��us�B��n��c=[�� ��'�^��0�g�ܮG����3b�&�۬c�ҕ�*��v�w5#�Ɍ=s�i�x�oT�s�mq�wmtg���uݭ��k��m�`�S�-��u�OtۛNS��[�C�l�۞{>W�۰l�h{�z�zq�Cb�n�N k�¯�9��$0��<�p�Ļ$[/gzS;�V��e�tS9�Ϧ�R�<�<Ƕ��LW=
FÛV�(�9�]�m�f6��֥;�]�H�@&8�s�)��LnƗ��<N.V�Xs�c����ryi�|�����ͭ=�H,%����d�v���1���=m�ñ������7m��;g����gr�9�d�Lc���۱���["ܗ.�xm��@=��.a��ݛ�c�tm��o.�mfo7n�nx����uC۷��޻�쉯�x�E�6�N��<��ު�P��m8�I�]�1�D�]Ƹ��1�3�\���8����qٗ��	�����n�Y�s;nO�v��n;{R�v�L�u�=u�H�\�Yp��U�g1��z�t�����ۙ;��lx����x�M۰kpkvy�`{cvݤ`q��Z���4<�:M����v.����w�!jp^�ˬ��瞺5�f�]8zEb�Y]WN#XM��UOk�։D�5���n�ݲ�@����3�5VRpSZ�h�݇��M�铸닫�t��˧���1s9���Z���G1� F��r�3��gmE��kqvr�n���s���D�fW�+�5�MU�tn�s�lwn2q�;g�-n��-��΂�}����m�h���NV&�ܝ���iN��9#nn�; ���9�@��s��ǬK�=���������V���\��k���C��������K˻l���N2�X箖;q	��
�q�H=E��c�������Q^�G,n���������wX�n�N��Sv4��ノN�ee���0E[{d�B��������v�'r�կ^s��v�qӈ�;�F�헐.'e�7�y�;��[���y�\���[����5�f�ڝm[�֙;L�ڈ=�v�qk8:�6�����n�uլ�>�	��9��Ú�)d�녽�q�%�ָv�\�Z�!n��2fiy�cm��vd㮝�Ѓ�.-׫vn�ᕹ���za8t�vsv�:'�+u�;D���u�pC�]��׶�א�8,k��xz�e:8���N�ؙlq�%���q���ێ�oi�.����766�U�Qٻ��{VR���
����pz�V��Q�(읰��npP�����Y��]j��K�e��qf�l�ݖ=����R������^��lǰ2.D�>+������6�ݨ�\�7�����0j�0�FN۞1Ս͸��M�>�ܱ�;�d�n�uv֍ŭaJ2d3�5؃`zSl��w���1�"�ۗ\�C��nۓ���n����8���棊��c^�ώ��s�ͥ����=��5nolsr���ls���tI���q=�{W�f��n��G��K��$�ݮY���2�W���v�2l秫��pmƽ�v�|u�lkBE� �UFpz�/1Ӂ�\]S�z���w�xA��v�گK���	��Ɯsv�g��À���BR7<��mqz͙���I��+�]<Fˌ�d{wln��mi��:�+���x�i6{;tn;GF�:�gg&�� O��[�mj�r�!����Y,6Ŏ87iz���$�'=A�wn��ym�cn׀�C[r;uqBG�ڦ�cv�����zm̜��4�>w+���[��&'W=�<����b:��m4��l\����*��Ϯ=�t9�q�:z��g��u�]�=��=�v�����Y�ܳv�Ԧ������x� �.�����Լ��]�u��9�\c��=���s�<Kc]�vx��x��"x�I]�����gY�Z�g��6�pqm��/=m�xzM���ۦ�9�n\��1v��H���]��[T��`��%�\y��5d9x�=u����;�]�{w;v�&u"�:˽bX2���'[�.MJ6��[�9�6���v�L<c<���V�M���]�Ӷ���;\����`��v�]7m��l&�ٻ ^3ڮxSW q�=�����{�[`K�s�������wV�5רv=c��&��l)!\���	�n�;v��{��[v��D�[iI�En;s���׬�Ӻ��X�ݪ�ݺ�&��v��Sۮ�5�q�@7d��D�r��m���M���b��Η��_<q�=�l9���K=��%|��L�b(���yWuˮ�;sv��{6�k��;v�6iyjw�xu>oA��ͯ\UX�I�;�k���=n�9�����Gf1�^'��[��˳ڰ�����nö��r��ۂ�С�b9���W\���F\4�y8��n8�uՃ�t@Vw#��
C�Kڇ
]��dɝF��۱n��ۮ�ݷ-�g���2b�n66����z��p��d7m�':�9�V���9�]�j��6z�/WlF�7�<��WX�P�<�rs�Q L��*���v��9��X��b���;vP��$u��6��v�rv�=ha��WX�rl��{>��r�mm�t��T����ۤ�+��1�`D9����$xy*7�]vU�<�[�;��:�B�WD{}g]�muنܴ�Ϟ����ڼ��9c��Ս��;s۱�p��Ϸek��v�k�����G7`w���)�ЄIG�b��m��qV{l�<�@vN��[�݅��
䑭�� �)��	����(�*��s��u�5�M����@�iz|2��{,GN��ʔǮUy=u�=�n͖�u������d�6�c� �ٴtk�ګ&_�a� /m9�m�����nvR�1!�ė;�h�ON��r׋nם��q��[�=� �5I3XmX�c��g�ہ�Lx)�r�����f����.G���Q�c�d9�%s��S�cf�<oh6v���
ٹ/6�یyе��m�}�j�cX�2�]ڎ�C>_��8�uҷ.��<n;���w\K�v7�2��r�a�k;������a���^��Z�;xg1�ơ��z.9B]����ҽ3���m��یe�W��]�	��Cu�W<�b��\K�P���x�����8C��..8��Yޭ�8�:G���p	�9�nW<`�1h�Gl�S��l;nOm�1�ݦ����`�f�Ѯ���Ŕ;b�'n=u�rg�8wnK��5���.N��x�睟tt���9^���v��P�s�]��5�%��qn�P����e680�!t�x[g�W#v�����:�Iݴ�XC]�؃3����J��F��؅	-��xkq�E�y.c�u�b�lX1ی==ӛ�.�cs�e{Y��l^9�+���6�GS6:�׷�N��갬���6_��W\�o�qP��z��E����_F�c�S�qv���	c��^�����<�=K�/n�'=n�q�<�4�u��mƔ����\�ctuJ띹RW��M��
A˵2m�:��H�]���pvz�kp�g��,��2��q�;;����:�c��	�l��n�8������l1���F���[q��m�Y�Z޶Y��e.�]u�nϭ��zy,�q�N;W�:w�bvn��ˬ��n3��n��n�<2�2ݳoln�8N�}�GIή�Ǯ���;�6��Sq���涻/��*Z�c��\�y��nw\��9���Z�p��n'�g8�\�[$�ۮ�oO:�Oc�K��� Khx�,��)m̓ �\$LV6�e��t�h�ٶ+�����sɵbȧd�V�:��;)��y;w@��kvn�239��۹��nc����^�sY���'\r�F�	��j���x�ʗ
�n%�1��0����fܻp�7��t�LW78���g+�p��s=�����]�M�Hn��m�3����c�!cUg���VusҾn{3����������m��3��r��#v�����*�a�V͜m����y"�����A�c���g3�}�B%0`��ٲkMr�y��\Ʈ���gP݃gh�z$yu���{4�FN|��v�Zw::8^�y�n��!
1͓���.%u��#�l)�.yن ф��z�OtY]vg�w-8��v�� ������9�N�y�paLy��k�A���s��v ������5#����m�ԕ����nn��$�&z��`�nL��:���{c&����{�ݸ��;�ېrb��q;{zk�8�
c�J7nQnt��Qk�t�u[;@..mwf����yAhsU��&�s��;H�Q�9�O�����=��rPY�\�n4i�T��W��i���n��� �(��7[:܂�:�vyM��\/k6J�n�%,݂8#dx;&�nū�X�wklA�z��kb�,��ݳ��Gf����j��D��"��y��k�q�ȼ^�ON��N5����1��W[s��r��h��������=U�6��]���uc���^��iS��O��۸�j�Q�7/b�c���v�'<Ymlic>:�j̽Qۤ�::�tg���^�5���V�u�;#ӽ�`��I7z�d\\ݮ��X����R�v��'5����9;=�'������{]dk���m�Y{�;�q6��0Ν�K�z�������������*�kŵ6�èRY���׵W�m���m����\s(���.5R9h���3�i�Q�i�j��\C)d����V�JZ��l�
%�֠m� �;�|�w��1�ϱ�3��+iK�2�
)�2�YTFܴ�H"�R�sj�EA��V�U��-*U���W�R����Z�s,J�+�F\����b��r1DiKm��墩KD��-�����ZS+s+��Q���J��2dT�vE7pvw�˽�b*+iQnR�YU�\j��2�Zf*-+�m��w&P�D�o�v������+�30q��"�5�Q�Q˗��Zֵ���lVʪ�pɘ6��L��F�(�����n<;���۞<dc+��1e�b�J�X�+�VێѵE�ˍq����[kYQL��eR�Ls*-�PEAS.5��nZ�8��.E0f*�E�U̷
�732�I�(֥���\\[DB�\�+��6I$��z��V�M[��{7Edx�l���<U��i��ۍ�&@����W<��������Ճ��잚��;�����U�[pb8�y�%ؼ�l��Ӎ�d��k��>���x�8�v�B#w��k��Vyz��9�=u��8����֎���f
��n���#�^���-.m�vw;n��y�ٺ�vͷmE�ۍq�l�g��ލ��2b�9���[5�`7�v`���h��v듶zUq���	b��v��휙��kSm�8��9⍃�[='����v����ŏ[=�;��.^�uu��PԢF��J���n�v�HlQ����ٱͮ���\g�#�7M�gu�RO=��P��������!�z��vi!]m�����϶������8�m�t�y�8�=��)��a{hܻ��.�9Ņ56]�h�;E]h�n.�ɍ&�79��nކt�h��]n�x��ۺ;Ry��-�t���b.A!�%�0y����r��F{��U��u�;J{c�ۜ�D�.y�v�	qpu�����;=�6du�E��p;�ל��]�F�ĎCm]t",���s�<vٗlӥJn�T٦f�㫅��n��g���CΧ�kN�V:���d뭬��!�ڵ��v�y9�-�k�������kX�[�X3��m��g�Є�%�9\��9����7['9X�{i��<Ҿ�ܷf��:q�ǭ��;WA>��ĳy�s�v�pwn�^�pq�<1ϋ��&�m֕{Wh2Ѹ9zۜ��u�.�Ƕݹ���=���OP����E��%e�+�t��s��x:����m�;6�Ep�o-�1n��ϧ8�2����{�������i ��s�U�i�7Wg�c�ڮ�����v�����IC�{U�c����J���0g&�c����8�'W�r>�r��sp��R|����Ec��{v�U��="Yոg�V��>;O'Q�mue�����n���N���o
dQ_+��9��y�!�ro۟eC�*nw≠.[.[�D�\�6W*��>���ܛ��g�@��;>�� n�q��nLryp��"�e�\-����0��8�c�ݜ�}�r��3�r������=�0�����{�f٩����7p�)r�p�rm�lc.w 'n��q�N�ll�68C��7;."&'�~R$�"}0��3*�3}.�� ��-���Wl<��]���Ċ��a���0�A�"b!*��T$�����.����_WH���$����P/�`�q�0�9@��鉔�HR!B����I�;��\Py�zj�%�Wfs~$�<�(����$�D�#Us�ՕB��'�"�(2A#;�@���s�6wV�s�������q(�fD�RȅL/.��q�ut��YC"��0{�6�'����t$M��l�Ս�b�����g&!D@�"#�cS�h�b�s��G��Wmd\�=�]��;k�s��&�w�Ͽ��D�& �		w���~$�:|H�����.ׄ���7Z	$<�(m��"�!H�L�4�y�J�/�UÕ4�a���#��&^�6*������o6�iR"��z�;�&�쓻GgcQ���ɻ��[�_C''�$_o�Pجۦۮ$�qs��z���#������/����ĉx�E-?VГ�|��|Iǰ�%Ll�ԧ�0��j�Q���d�z��L��B`-쾶�F��Zy��o��8��wRI$]�s���{nE�4$=�R#1\ȟD�I$��z�e�S=���
k Q ]�s~$@���ˮ<�p�����w���5ure.j�ah�an����<]�.�{m<��e�-�V� ����o�mk�������n��|O�m�?2	����;������3�Y�:�	����"J�"`�RQ��Ve�`�	ᕻ�
G^�7��H�^�k~*�y�O���Dd�S�����wd� ĉ"$L�1<���m����/]��A��&g���-�OP-L���I�5:ӝ���/��ͺ�5خ3��k9���3gnw1o�����n��!F7�H��ڷ�������A�����F�0�(Fd�%^�=��4u�{f�Vk(��9͒|H���>���1㼮�3�by�.'���Y�&Tġ""���]m��9t&��Ɍ�ʓ������$V^���z�"/�3ԓ�1��A��0�MT<�#��g���N�X��[��\Y���Z���d�ߪ��?�d�6S��� /K�~����24S��m����D����|?&����y�Q�\$w�OĂN��D��R��[;�ƳƂac�e��� ��Ę��]j��ݎ�����d�N��ru�fL�&P���s��.W@�GI>*1�2	#���q����DB��ú:�]{��,��<F��=���li�R��Vk��UN��"qR�m��ۂot�����k<�}~C��X�7�9�"�'��f��[;�_�>k�� ��*a@P"$D�0$�މ �y��b�nĕ����"o��	6gn�q��`��ٻ�Wru�p��܄�@�F=��ѡ��nɞ�b�#wa�`CbyC6M�o?����&�L�! �~n����ٸ�`�7�7t�Ğ�w�����ǌ�Г�W�1&}3(�L�^:�d#����wwus��A>�9qDy��&Q¸�����+���h�t�"ARȅL9w@I$���`��&h>[�1]d��l�]	1�sdҩZ�%"L	J�Uyw�`���R�^mJ�~$;WRA��y�v����)�d�d�x��zO���"T�"&L�6k;9��|v�m2;3�d�^.�(	�٭��{͚g�J�^�v/��2˧ݍ�����Y��������.�P�>��-�Kz�;�������qo��i~�wÉ>C�B�Q�����7��`��I��^B{g���Y�j`�x��c���N:�۝��o^�ˮ�t��=4-�\�V�G�n� ��j1U��t��1�:Ί1��a����n�<Ύϫ�Iv�x�ܽ<Y<�5[<����Cl�dB�IǴG'c��g/-�9�5��m�t��ƍAҰv�@P��on�脻le0	��&�^�zslӺ�Nn�N֚���H�֘��4�����X㳵��s��I�[_�����.x]EJ3h�]H ���d�.����:��%N��骺	 [���>��8ĉ��L	F%���l��\z2˩�D���|O��9��{�?��f��]3o��� ������Dcl�@M������'�-�P`�a�]ۏG���el:���$��o��4mGzD���	��ͮ��l0p5��O�����z��`�H:g������1TK��=�yA�U+T�Q>"R�"Un]�~ �ٞ���;df��7Z�����d�6�kd3�R�ڣp;�`S9�g`��N�����K�m�;b�l`�!��5��r�[���c�C�H>��Nq��$�����5ۛA���i�H:��(2"�d'J+��	��ɔoY��(%J3h�mIv�FH����r�{bص��ܳ}b+��]��j�=�I$/l��#�U�Y�f�d���Rk&�10{��o�*�J���F��M섬dN�k$��}��A>:z���=[c.7���z��H���`J1-���l�I㕔$��2u�S��\n�US�Aw�����*L*�31L�%$�;��/ݦ��o����'"�>�^��0��c�2s�d�M�zDLȄ�<^]	 ��y���gwVq7�;_ ks��$��ʐI�e�6
����.��`���Dq����\�f�qv�3�=�e����zx&���\��?~?K��D�"D����H"�NEI���Z���j���߰�w��0
+��z?Y-I1(�ߍn�0�;�vj�]��*��#�NEs/y��/��S�}��@��( �%B3�GkhO�/��|Fgg@��R�|1Ej������tY�J��wE�ȁ0o2���W�V�(󭎬1���uΜ�j�qyё{Р�US}=V�I��y�f�[ʂ0��wq�$�=9^�A#2���8ĈS"�M8�|�s��I��qD�y{��$���h�#qF�\2�Ysj�$�U�bb��J&&I�z��'.�i�#L��ǆ	j��'���$w}��g�VJC��f��g�o	Ӥ�����"��tf�p]q�bK��[��\jr����wϟ����x���!W�K�$ng6H���g�z���� ������ ��Q�0b'�BR$J�o�	$�x��G�ܐH'�3Xd��sd���"�5�a�'�a��qZ2�IfICf������}�� �C�W0�a���p,���͒	�y͂D�x�(J� �A�zt�.Z�����V�S���L�p�a�&�
�o�Ts77N�P�qS���1�w�Hز��ߔ�f	8�%���%rYK����x�*�\��z���wұA=��*��i��1"Ȁ��Rߦw��I'��P��i�Q��N�%�o�m�6 
�
��/���B���R#�<�0�nىvۜ���Z-��+g��qv�o������u5��t�"`�(��'�t�l����I$b��ֻ���ꪫ$����#\����"`@��<r��nD�2��1����A#�lN��j��ǿs[��q���&����/3C��$�l�eI ��ޑJ�T`Փ�5��$�{͒	��=�'�s��*T�be��[��2���w���D�S����<�r(�@���|�%C��u�H9�a@�T	&!�4g���v�����Y'I��]��A'��P�A=���8o����Z���������˱K��>~�&vwn�zw�W�����v����h���~X���M��0��u�{�O"Z��ЃÉ#��!���b�v�c8��M;�Z͎�uۧ�u����p!`,	��q�74��/j3�qQ�-F�㡣�Ṋ�g�u��V���̵)Ҡt�N.�s��-�K������q�'%�hRi$u�M��*t��H��l)�4O!�6�q-m�=�)�p�8����r1�/���7�:l�ݙj�j��95\;s�{g���C\�P�f��7U�4��]�vMt���p���V�WK�i _���fL)�	P���7Ym��I�9� �w79�Qc	��]X	$���5�ƄD��Q32��V=����*�c�r�w+I'ĎS�I�����eQp��e�WLeԠU痐�`Bl�˺��Iy��̂L<��fv��A �3�BA�'ۛ��"cb`��D�R$J�w|��m�Rmо�@�uT$�A���&��:�7�˹�|t�:��:�30Q2�Wohd��"����u�:Qɨ�|z�:�'�Oy��)wF�u��[pu(�p<	�<-�V�ly�Ʊ�ŀ�7=�9wY�ܳ���=m��ϟ�r<�=l���3yBA;���$�u{̓zB(LU�b���@�O��9��x��Ʌ2 !*�'k��As\�Ws�M#7,kNً�?(}�zS�룒�2�U�����[N�P00��(t�R���W�����.���,�������9���&�s�> ��g6I"����$�.5�1��3�$(��1���hO��� e��H!� �s1����>�i��u{��$�@��/!��ߏ�ӑ�+1�Ɠ�w�����oĂN����w�)?����1{���j&�xX(���X���	6g�����N�[�B$6���y��|I�=�%�(q�g-�O�:�U�}�;v^��.+t�W:�(#c���q%Ç ,,����Ch��޹��j�i�Aا�(�;+8���ff�	����&B�f%@�b��h�mzI���O���Q��|�$��[� �p�d
 �Y3�L�{�ٺH�kt̘Q&2�K��u��@<g2��N�L�ٵpY]S'	�����E	f�X�@��<���Q�������=���JF��j��	=���v˞;�=��=���f���V�W�̀��DS|;��ъ��^�D�sj>	c�
��뮬�L٣���>S�r����Z��ӣ���F���63M���\�4�7��:^3���>�6�}�%�J2���J74�s�B61K����U6/�N���v�bhغ�7j7Ɯ���L8V�C4�jكú������������/G�C��2WZ��/f����-Xvv��;f�cL1�+�X��B�?;���پ|a��>�l��}����ў%��6Q0us%�+F��'_�C��tV��eȪ�,�����ޣt��O+�a�����c�܎]NՋ�g�i�޺=h�]��F�P�{��"�����p2�3ڍln9�(�;�*�� U�bNՃ�IgcE�б��"��@�]ʯ���$��
Ͻ�:�0"�O#2�{��E���w3u�!�|�[��{�O�S��÷��n-����m��mS�U u�.��$�����d�g�{���Z�UvF���{��N���KW�H������ $�3u{S|c]���=��>�.�F�tS�P��s)4�Ht%{�c�Ʀ�2������}A��u�>������l�0pr�<��=�z����幩��07����xt��򺗺�0�6�*N��C�c���Z�ng�-�����5����fZ���<�«�0��$uAP)"�%,�������`��L\�1lSr���B�h��֪\nS��V��eYe���-jԩ�UP���1Eq�2�e)m�֙aKp��KF"�\e�&f`��B�\s�f�ff8�1��kKUJ�[K\LQ��ڹ����fV��eǗ�v�]�C��v��Z	[-�3
6�
�X,ʉ�*9n.Je�V�2�8c\�-�s)R��l[E*��*.+E���W0��,�����8�
*2��֖���J��-ʵ�4�0�kZ���Z�.b�s.	�e�(��
`���2�kFF6U�4��IELl�*9-��66ڗ-��h�����R��X�ᒢ*�ѭ�m�eZ��mE����ۀ;�8�U� �s�"��R��KR�ԢULLf)�QfK\��[��R�K�v���]��v�;{ov�J��p�+ZR�e���m*����*��mK,��--�c�Җ8��A*�������g9�y�|H8g��$J�P�&���̚;��mf\-�����~$�{"�>���]�o`tT������l�P*���@�0!6��� ��Χ�n�����6H$�{*A ���bU�z���C��Ds��M�N���ku�]�s{��R��$�;����<z������1qa�+�n�A ٝʒH$��l�Z�+�+��������>�ۯ���@\&i�{���Eg-�_l�pLf�$A�;�Df�s~$�D�NS��N���P$�*bhэد㽹�2O�d�j�,����Gp�	:gr��͓Oq�0�I�L����u�������! l�:I���lM޾dU��;�
������n�ݝ!�̌t����|nX۴#�cTTt����ހ6�K�qK��Ş3m^�^�wH�;��s� ��-��$���`�:m�2��2�mI;j"�&-Wt
'ö�[$�w��Փ=.m��k���c���q���{<�nzq���{[�n:��<S�2�Q
"*��|��p<vr�y�����`�呻��.k�H}y��I���&B"$T3.��fP�ݝ���[:I��~$�����H��͂,D�2CP.M�ԑ�5����L&[��H��� �Y����^ı��#A���7כOēw����M��_��Qi�����:3��͒Lum�`�|�>��]��a�e'��5ַLI�L0f�;n��I�*l�Pyw��uسԲ��QX��$�o���'<�<[Fs�@�ۯ��I���7�cGV}�z��(HS��ν�IX�A��v��W�{*;*]ã7s))�v�uq�˗a�_����]� ���C���ɯ< ��
��n1L��n���ҥ�Ň
d�ρ�\j=��6s��cN�
Tt�v�H�X�m3�8�ⱽss06-l��[,Ӯ���s`ʛ�������β��;�'kk�M�9�/���O�*�ٌ�����1u��Ů�������2k�s���j�9�vz��.V��Y���h��{uN���i��;�����Ȥ� ���]�,��a�]�n��(�u�r���x��qjNXoQ�����߿�C�ݰ�2L���?�M��N^=�|F.ys.�ҎF,��o���}Cj)�D� @���^��c�r�>�S.�ĂE�_6H$����p��Yu7/�ǂM~��	"������ �d�� ��]66Ek�٤����2I8y�	=o���� ��Xp����_��g8&���2�s��{7s�{m�J}�H���$@[\ ��P$�
bh��ڒF�液��:�N湆I�+��9���!�3��u�MĤT��
bȸ��]k ���A]�5�]՛����:��v�}��|�L"��4~nY��f�q���.�sf��Y՜W�*2���� �l�ʓ
����d��f$�ޛo̔ok�N���X^$':'��*�e{t$c��iD`���d5"3��Q$#�)6�>|�P5�朊R��^�E[9��\O�$r�ȢNv�S#.�(S��5�E�}l�D���H�0!P�Z��H���$<1]�a��o*A�ns�QfeJ&"�*�<�}�|7!2#	 ��ʟ۹�0o2������'��C� CdR����� ��Xf���s>$�e�2�������j'b�>'�3[�$��/��=�B�# /�&�������*�GX;\��s���]ŗN��^y�;GnMv�m�u��wj�w��ϼ��=lfg��st'ݻ��`��e�2�)�EU$Cp�&=WR��gS$V��1&H�QR%�=]l3�E���Q;5f�\�	35�O�2��A�C	�E��'Щ,O�H��
bM�6�>����Ϩ;�	yW��F�:�Q�Qi�Y���
�xT�M���f3�h��9��F>4ϓs�W*'�Y�)/`!�9��ڃ2�p8����4~�w[����*T
�	����p�8�Yc%B�������pIX_|�[��]kO�υ�����(�o�(d���	#��1
þ��vpg
�S����@���F�(׷���v'{����d?�|��.�|*�v���SK�Z�t71sFk���;϶x�R:2W���vx�C[w���^����Aa�Z���!�T�������' >Dx�����Q ��E�0��߿�._��N"킱=�����!�5�Q�.9m��۞�Z���|���%S�J������,7��{��<`X5 �{�{��JB�B��[;�~�4�.�����:��m�	�y��Ì��YFJ�����gh�����4���m ��k����y3�PӅ6��gۇ����Q*��}�Ă��X�����R!��ճ���:9�b2��Ο �1w$B(�������Ă�R����=d�T,#��*�9:_}��Q������_��>,aRT�����$N2����ܞ	�
k<����i5����xT��ߵ�l��EOd��<H��hx*R��_����O
�YS��߫�ϣn�7S�GP~��U���T"m�`[Iȃ�Vo��/o��0�U�n�c
���!WM��h$�R�\��˙�{�k�/��~;���I�%B����~�ĂÇ���zb�ц���8À¿^{�p4��*J!Xw����<d�_�gqQ��}��޲ d" _Uw1d`�D��{����7H6R���ۇ�?U�n��7���i&�@0a"%=�v����m�R�P�rܳbzK<����+��6.����j�c�h�}�s��g�e*A_�wg��B��Q%a��w���aXk�����4������8�Y82�Q�����O6����]kZ��k30u�Ă��y��c�jB�~��>����V�Ik�~O��� Q�D~���4� ���߻���q���<�f���$�z�7�2<��b3����a���g����~�<a��!R{�}���2VT
	P5��������`��@�<	�m�p4�|�-��߻��ǌ
������2"
*d�dX#��<�dv�p�#o-�c=+(�_�}�g��Bĕ
$�/~��y0�¤�?s��gc5��~���"/> ��O��>F���y�H������kY����P<��_~����F�)h�{��9H_{�ӳ��s�G������>�'�H,;��p񜌕�d�Q��~��8����ݮ���UU����ŮQ�Y�1���u/T=כ��q��W5w������A:��'v�=ǳT]f�ϧ9Z���T����3x�=���|�Ɩ8"Sp�,���Ǣ�۰X�s�U��ݬ䶺ݑ�6�]��WLB�'F7�F�n��n�� ��YϨn��;��X�p�V]ش�����;l���u���Ʒ݆ٗg��`]���x{z�]�.��ȅ�qٱ\��6�n����۶b+d�E68�a��g����OTt=f��2g�כ�\����{�͞�&���_��6��؝[��7mv+=lu��0Vڮ�h�n��W"5�-GZ~��߳�+�4��C��
�y�퇃��
þ��n2q��P,?s��È�X�租�y����{��Z������n�m!iaϾ�ۂ̓�S֙�JD(�1"%�!��w�P�,��=��Σ[���B��T����~�a� ��~�{��$����w�7��k��xګ���� ^���
ff
S1�G���s�Ƥ,������R �������Ϲ�>m���`i: T��'���w3�%H(����Ă�e��a���f���~�77��ڼ7��m'�T�B��߿{��8�YP*T�?{�8� �����UDKs�w����$x�����g�#\sx�����5��O}�,�����W��;���h_����m|���%Cĕ�>��;�8Ã
*���<I�+%Y++����Ohkzy�����nx���Z�6�������ivۄN���ݣ֫��{S���%
7>�����~wݼ[�3Z�_�蕇����x��H[@��{��
B��Ϲ� i<*g�|���[��x��g�s�É�d�T;���g�J���V�ύWFi�3�p�y>�O��@Dy[o��I��n�ub����P^뭉�^l@:CZnam�6��\�����Gb.y�{���s����X�^ڎ�׃�~�#NvI.��|�9k���� 0Ͼ�ݟ�8�YP,J�O{�� pJ�R��s������8���D��9�L􊊾J;g��'���K@��x�}��pϿ�o��N VVJ�+�����hPIP��#�]O�`�o�|�Ȉx3�g�0�(��{�vq'��� ������&�,������Y���Z��ׇ8%a}�}@H��1Zk�W��0Q	 Mg�<�HZR����w�O*P@�;߾�p�޵�c���6�*��~��8���3�x��&a����!�F��~�<a���X{߽�g�NEg���񏔍��	��X� �� �(���;�������}��Ï#���G�Ov�����\3L���OYnT����џ5�nxT��%����c��9]}���in�e�Z~���&������e+(�_o���6�T(����}��!��+|����f��g�w��$�&���l�N!Y+*A{|����U���ӭfkY��@�����䅎؆�=�w��ɻ�`��$�JB�B��_��wp4�R<���>��"<	���:Ig��o�?$�����tf�3<�pW��l<a���Xw��휌�%PD �l�6#��GE9g_'��-9=C^ˇ��r�ç�<n��F��+I���C���Nz����{�<�#�c�R�=s����N�[����q�<���湖������������F�(�������������< ��ė�`�R(�0e�@����������xx����%w~��FM�D�
$�)�{�|�r0�%O߻߶q'��w��5���~�,�FVJ�~[{^�Q +��!(������&X���߽�p�Ƥ(Z}�vx�����t���|)��?$?
�YS��w$q��D?~�~��x���5U���!@�
!+��r�Ӷ����'=g�3�p��]
�S[Pn=m�u��te�.:����a�
���wI<�(�a�{��3��eH(O߷~b��G�|�1�~t�Z����Q�u�w�t�e!ia�w�Ï#�5���6�F�m֟ q8�z���8�YcJ��s2�i�c�Q�̖Җ�T�����{���+
 ~����Ĝ�����i��u����9�j�/�W��Q )�_'�I����L<��a��� �w�{��9)i(�j3��=�&��+���x	#�'�~ﻇ�J�2T,C����C�+��_��Fi�3p��_e���_H�~�#Ȁ��'�o��Ă�D�?~���q �8�_^׀����ͩ�ό3h�ј]ҼNk�1�+�?�m�׷f�AvM�w�%���+��\һ�Yqh�>��Q��ݏӝ�ם7��Nͬ;}��&��{�H���HV�����Ǒ�Zo4��њ.9�X��<w������R(�_�����d��y�����to����%a��}���0�(¤�������8!Y++%e}�s����w��v�%O~����7*8B^H��A�K_'nU9�3�gJo�;��<Ӹ��kf�/��ػ_߿��25�mֵ�����}���<`V������ �)
с[�}��I�O>����{��}�q�+(�P;�����8$�.�u�hˊ\u5sY�4����~�<m%�9�i��_�����~��p���P/��߼8�ȕ�cX���wp4�|�/��f�YAL�5��xi� ��8r[�F���O�8�o_}�g�������^�<d�IP�J�y���7Ͼ���a�aXR0�*~��~�Ĝ�VJ��Y^߹����@�_?�!2��J�H����2��|�Y��%�=��`~jA@��}��9H[)
с[�w���ȁR�
�'{�~�8��^n����|��c4�P�׼��!�%a���q�к4f�37q�~�����ID*J�a�{߶pg0�����=<���@�J�f����q�XjA}�s�����HV��p����/��|v��n:Xɜy4�|��XX�Ŏ�gS�3���{�ِo�w�ճ��� �Y%�<�2���C;���j��T�4�������2{�������-h��L���[�ݗb ������.���Qφ�� i�{�q�5�^�&��W>p��o��{�o��j�ӵrKd�\��5j9��T>~�m<���]�ݺ/�ه�#I9R�:��*u����� 6B�s�8j�:q���U!,�������;ä����P�-��1���z���,��������]	kݽ�`��=�q����=���s����#�w�ٽ��+�fՃ�Dfڪ�u#.LU�GzT�n��=R�!�m���icm:Wz��
!�ɽ�������l�'��o�}��z��]{c?<V���U���xٓ�ъ������&̷F?���NN�ބ����,�������~Γ$8W���U�+�R磆VW`�X�sw8�v�8 ���N�ÌA
���DKfJ$� m�ҿv��bf'�ݻ������ۨW�b�'Y����!�[��C4gޝ�9O:����
c�)�6�o�n؍���+j�+5
�2R�����5��6#���Dp�����GݍF�5�YW�N��O7Le�iuC*١e�W��c��e���?�~׽��� Ҋ3��5P*�C\�����wNMv�{ٳvpq��l���9_U�ű��on��3��{;
^���B�=ȡ{��!:b�o�+Lv*+/��K�#�;��݇}� Vf�g1�S����	0���J�����>JP��_���w����ɺ6�m��j҉Kb��̳+iT�R��ik��)X�JU�F�F��2����)X�2�Z5+[��#��s&J���KZ���QjX�m�L�Z�+*-��i�qQ2�J�Pq�Ŷ[-�D�s������#�`�y���|�c��v��=�a�aFT��+EX-��feZZ�����\��ڊ�h��r�����ȶ���0�2��V�<� ��!���yM�wn6������{yx{q·����W
UR�����*Pq31�Z��D�k�250�*�1J65hڪ���ƈ�n��;l<a7q�x����cU-��Q�ˎY�-(��T�Ɔ+kR��W���Km��*�Z�3&��2�*���K�r��T��h�5l˙1.6�d�YZ�1�V�Eb\��nS��]��6݇+���=���JR�QR��,R�-���QW����¦E�UDH����Y�[Tq���U�3w�pv�n���Ӛ�ў����r��vc�mn^#����Y.;p�G�&=a����,@����'c��R*ٶ9c��p���64�[lS����;n"�U�������-^����9�v�ź^��`ȓ�^'�����c^���<�ӳ�[��c!��e�����)�˶�6F��q�v���1�.-�l���ۙ�����3s��������aеûN�(�;[���"�$ݶμ	�;�U�,����[�=gn�F<���ŷ8vݜV
�����na�j��vԙ|�ku�G��w.D�ǝ�Wn���%��q��e���l�<��v�g4.u���:�㐵᜼���:�m>��Iˬ�ζ���e���`H��v��t����w��fJG��:z^/vۢ��`�;ծiy�o;X�.��h�ۤ���B��Hm��6�v6z�-����"m����`�2 '9�77-۷nn:���"uI+��v^l�{q�푸z���d��W����1�D����#Ǜ{=�aԧ`@]m5Ɲ���Y�r�Zv#nٯX����ՙ��^M�N<D�ۉ����]]�H,E��۳��S[����r��۶�[uǢ�`%xP��2�s���r7\ԋ�2rtg�ݤm���f'��ɥ��td"mv���V�[�k�ڏ	��{A���v'%���Z\�-��	��[cv�N��-��oW4Oad��^jt
��ù+ׇ�4��5\�8/[&{W����5i���؍��1��Kӻ<��g/Q[�]\ev��xŵ�i9��}
ѐ�v㤥�gckv��$�w(�ۇ��m�>���.�a�WnSmyd��� �-Ůθ��r��ܗn�1��wV���f��ͽkku�6z�s�&�zr�c�[��;�l���Rj7Oef�\�������t���q�x!V��s�n�.�t.CC/��:�O&ma���R�bݣ5u����w{���������3�����m�,�&�\�g�ɹsb��Мl`�ȹ�ܼ�x�k�1�uf�6�y������{e�wm.��;��*�v�F�:^X�Z��y��[�Xx9z�:�З���yq���8�e��li����ۇ
u���x�x�pv��B3�{e8�����gm[��V���z{Us��kr�_Y���.;�͟Xiw ,U��-�j��l�@���\U��7���]�Ų�^]u�[r���?�}�X�K�e�:� T�������q�����%_yݞ2m
$��w����w����_*����]�n�$�B�VT��~�wH~߿��֝V�k0��8��JÞ���0(G��R��o]�3�t���(�>�y� i ��߾�<g�%H��{��U��*�+�wC�<����_sFW*fjj��i ��k݇��
Aa�~�8�$
�����3��K���f���@B> Q�������y�A���ý��nx0+�^���H�"S&�"��O�e#s^�?�X��R5+���g�&Щ*Aa{�~~|,�"<	 fn�A�����޾gׯ���ɰe|�����M�SX󏢔�]9�]_ ��=�6��
5!e�w�{��9H]y�_o�;�������$�����w3������37~��G���<���ձ{h�����SF-��&�]kM"��㦀W,��f{s����}����/���ow��W��l<a��!RX�a�{��9�J2�T�~�����	Xק�_�{��_�H._>��H?R�w�}�p����34�.�Ne�:�O"N���q8 VQ������]5���������3�����,�(�s���H����ݣs����UOn4UK�՚��bq�`I�_f������Z�S�ɝ����s}�B}'�����ɴ*J�X_�}��+T�?~����$	���{�{���Mi�����u�o�� C6��(�2������dd#�}�}��<H)-��}��)
р���A��EEF���G�#��h"���8�2VVJ�C������pIXX~bv�@PH��J���'��iO�@r�1��s����5�)>�T�
�{�>�<d�eH(~���|8�ȕ�F��������3��8R�����7<���~��4hշZ|���M�߿l�p@��� ����<6�y���q�����$�3Ϲ���aXQ�IS��{��$��d�+%_�wrx�@��f1_�� w���O
�&4egݫ�[!�[�`�ŢF��͕x����~���m�f��֮����V��?l8<`V�-�w���������������� DC�S"4ws�Y: ��������T��C��{��$�����к�油�C�����ta��
��o�nm�7��E��p|>s�^��x���{����q�Xk��w�w��G��5�$MFB8����|�+� ����B�
L��� ����� �d����w�vx2m�
���	���Vw�YB�ٍ�fj��������_���6B�~�ٟ�|������JsEpw�ym�M�ݿ{�b˝]�U���=c�� �����GLCh�Ibw�￶q'*Ad�����u#!��s��$�JfBX�<	�}}@$��g���37��x<1 U���HT��_��ui<+,N�߽�8��~���~���3]��nO�g���.L�vCbMg��ld�'�nv��z���1wR����~��P.y����"V�(��������|���w$᯾�4��{�^����~1<���y��lv�ֱ�:�{#ӹ`���nL]+;&i�x�������[]n������O;������YFJ�2W���<<B�*%aw߽�H,��os�������>�I�>�wgq
�FVJ��wRy�7�x�)L�ӭi��PGç���l�G�<��F��Q�^{�6y��-�+F{���O
�@�������g��:y���b�T�{=�/���dx����&'�d���g��+�~�x�ĕ
�Xw����3��P(���<����Y�y���ӈ�*A`Q�w�ځ甃iAxf��^l�W�$���J�(A���@Sě�}����������:�2VQ��{�h�<B�J�IX}����x|/��| <���#ӝ�믫~���������n�!bxM0�tE��͊w0^���s5��k���'��R�I���"�<�1[Z�xHܬ.�\�Wy&w�]��#\�/�.CJW���nOh{��p��.�YJkÉ��s�퇣����<����
<��h\:��_p�G�"�W[�C *Q������8�YFJ�C�߽���,�#�[l�%v��c �3&V��R�rۆ�s�盅��Y�<w^M{t�^�>��v�?�����.jk2��i��+��߶FIP�(�a�}����N�J�g���@B>����v�5��8�`��}��
A����{��ǃ�ޝ��*bf��H~ȰG���BȲ G����������7a��w�O.�(i���IP�+
{����8�Xr*J������ #� |�����k����?O�?wr|&�.���b�5t�Zu|+��~�q��R���~��%!l�*Ay�|���7��k[�I��Q;����Ă�FJ�������q%as�>��:�M�7Y\�!��幔NdG�6ME/�|8�2#���￷82�Q*y�߼8�Ĭ
��]����~.�~�~m�;)l=�|��ǃ�t����[��c��]�S�'|��vq8 T���_�wg�JXg;þ��7��1CD������%�~��8�Y82�Q�8��$ ���^����4V7wZ�.��&'��E��L��%;��1N^�(\��rP��+#@����HK��J��%�*����.��Cb#�;����s�禗33Z-2WFZ�ִ� 9.�4�v���m=P]��s7S�탠7k�U8K�]�Y�6K�.ٱ�JUͽh�ѹ�B�u�9<��<YǶP�lY3`#�q�9��v�L��G'K�t�c��9[��D�^�⑺�v��؋�˰�g��'h�D[[g��;�y{�=Q�8���s�7W*��Sˋ�ƏrF:�C��/��W1F�b^:8��;V݌�s�ė[.9�wb���R[�����{�-vPq�����Xs���Ï5 �w���g��-�+X��o��I��S�Ǐ��]��2�~��ۇ
A@��}���%ap�����u�!��ۯ�߀�=����q��u�]�3���:��d��*����8%H)�k� �Hx���5��:G�KF�/�y�u���߿�O���їYnh��&��߶q8�YY*A}��vxɴ*J�V��~���߼5�s��XT�������g'T�������6�K��}�L�Ӭѫ�x������nM�}<�Ϟٽ���#����;x[HV�+f��4� ���߾�p�>����ϓ�vJ�P�>����8	+�w�sN��u��W3�q �^󛁤��*�}���2}�y��o�<�6���{��sÈ�Xk�������A�!m������0+��'�{�5m��ڶᙊ��Vڈ�tP�I4�:�niN��O��^��pp<��~���Ţc��}���>������H,�������&Щ*%a��}���0�9��w�o���Ԟ'����H,�ed�+�߽ܞ&�)�w�\֪R沔� q+v}�x3�,G���9�c��UC��ZaY��.;�ơU�/^uH��]�<�bZ+�n[ֺ�k��k�"�tP1 �Fn	��^��������$�!��~�g��!RX�ٿ��$��������,�}`y2>]�몧�f��}�M~��Ρ�Jp׮q����u�!�0�]���i ���{�x��ʐ${�����s��$x�,���k�=��-��߾�p��l�^�cu���Q!� 	���22��\���kV�u���%{}�g��hQ%B�+���wq�aF%�����gs~}�y�Ɍ��^�o�����?q�-3WN�Zo��X{������Z���w�����!|�zw����!������|���@�P+,N~���g(j�033�IL,b���o/���[����}?�����s�rv��zz����ƢQ�U�7�N�7Jcr\h�߿���Zz��L�|x�^�y͇�6�� ������N2�Q*߿{��8���~>?w_o���uH.�y�p?��K���y˧�t].����ֵwOw��P�<	��y,ƣr�#�����7{:2m
��bJ��߻��C�8°�*J��~��H,�VM������;=r���'�������aZ\�R���V������jB�~�ݞp��Q���T_р}_E����fŤ~[�۠!M:���|�������aKǧ �����������£Y}ַۨ1��q�@��^^x�l�`T�a���p�d�
!����q$�)��^���%�K�Z�a���*��	p�/czW�Gxa�#��k�9���d���@����|8��+��c_�wp5�}���������D.{��Ũ�"_���HT���&h��&��߶q8�YY+(�_o|씚R�
�W/��`�
��9��)�,80�*{���l�ND+%ed���k�dQ LW,�6]�Q#P` �lR�܅���x�(����ݻscj��dc+u���׽;ߪ-1֋���(D�=�~�q��!K@��{��8��![+�#���$�@���v벡��}��ɝ�~�8�2VVJ�C��{��$Of�bH����~G�<�]x	"v!R{���|k��a��y��Y�KP(��߻�|8�R�_����t�JB��߻�߿C���z��Ȣ�B�
bdI��O� ݻ��� &VJ��^߹ݞ&Щ*%a�}�3)�{�}���<H,8¤����l�NVKY++������u�磓L �1dd#�}��@NK��3�``Ԃ����ݞr����[�w�|����Y����w3������kj�|/S�I=�CsF��?.�'<��+���{���*盛g�X�瞳�&�O,mLZ}_~�L]��~� �i�̕~{��!Ȓ���g����d��tk^CL<W/�{���"#�����}g���O�Bu��=��9�>��A`q�
��������ý��w<�y�߯�����r�������GV7m�z:���[�ʭ��:�%X��=#����������$�o�����_��������������6�R
w�}��A`�^~�����k����O�y϶q'*Ad�+����Oh�gؐ%zfDD�L d#�����π�
#����ݵ���t��;���!Z���}��@�x�R�VX�����g*AC����흷�o�~��=V��[��Ӭr��3�q����<m%B������8�YP(�|����c�3�t��V�+^��wp<�)e�������EDQ��0!)�ffS���^��,�>���N���p�`�Dxj��x2m
$�Q%ag�{�C��#
����߶q%������]�Ad������[�ryh?yמ�:kL�f�$�}����R�����w���w���G��G�#���WW�� ���߻�����������ő�O���i>��!����LU׍8��S��a�w� ���y���αUHi��:�8�>�~��NSѩ8��\W)\�'2�+%�қۃjhy_�����|L�$�ڏv�����\�Y໫��_���������^��躅ݠ��ښA׋��.qs	�s<u�'k��t@�cB�)���� c�ti�d��6����ccv�g99��N8�GsNDfX�ucs�n�3򩽍q�i@L���T��u8�<��q�\ḍ]� 5�9�ו|c�c���m���N�N�:{F���)��\ql;V����]$��g2���k�G�1��k5�3Uhht��>m2\Ժ5��H-��y��IP�*��}����NFT������8	X�wo��]�S��遍}�o���A�!l��ouxY� ����B�LDL��,�k���g����폴����ߤ�Z��iD�
������0�aR
��߶x����VMy����7����>�p4��.����ɬ�֌�R���~0,jB��{���$��]s˿���׺���@�~@�D
�'�{��������
!�{߶q ���_s����˗V��C�8+���7��������*N%�=���g�JʁR�S�߼8�ĩ�Z�����wޛ�?w�����B��ÿ~��Ï˧����kF[���<}�~����
�2T�����<��B��}�/=?��%ak�}�8Ã

���{�8��
�FVJ2�Y�׼�E�U���nɦ�H(���b{;�:�n�i'o=sܱ�Mb��\��A������~S5kLu�)~:��V����8<`V�(Z~��󔅥 �>Y������9UM���8Ͷ� �ٻL��0-$(�)1E�@I�;�5L�%�e	�������Ul�������o���h��s~^�8�9��εJ���֠�G֍MF�Y6
F_%�)������σ$��gkg�o� �o�������g�ɜ��
LHQ1"[��~$��+�|	�1��w*x��fn��$Y�ȯ�@�1鈉��u�v�>�Rl�w�A�m_dP$�w���o1+��c�H6��H�ǉB�*�(�6t�آA������꭭P'�P���`�8�eO��mv�w�����_4m�I,�KM��hI�\U��7�uڜOgTl��ٶ��2���?~�ϷO%L�0�a.���A�{�$�K��a��Ӛ�^�a���+�F�����f` ��}�4���팮����$j�"�H%����"��.ڞ��؍0-��)1@���I$�ݧ�O��=��ڿj��~�k�ǭ�u+؂
�vۺڡ�Q�/7^��]�s�a�;����L�����4yջ��i���>.�i7�e;N��V�����prk�H3o�
�ƍ�������g�O����}���Pg�]�a�O{��H X��6&J�,��N�F�j�e����P�Y%�{���^Ѿ���ro�y�=��~�Ӑt�?y����7yA�=�Ǻ���DC7 ���.��ꆗ�9�Nhu���㼆�WJ�4{լFn��sfAsEiD��
��6Yܪdyy�Ir�m�{��ۤ�A�O�WU�Ë�OP��6T�&��6;w��s��ų~�GoOy����Gv�{ݬ���}ޏǪ��-��zo2�t璻�C���f�D)�	eO���̩۴�P�_�Wy�o�V���f��-^��LM�%�`8,���o����n�D�ieR��}F�r8sK�������.|�}�?.a�~C+a�<=+�K�'aM�j�Y˱c_�(;5P[��N�ɼzEhn����H���f�:=<g�}�VX���{�
���$]��r��,q���#b�I!;�Ár���-F�����ǜ��Jg�˚�˝pWP&�f��z/N;��q]��ddyb��Ӏ,pg.��꟝�G'��=�7|��U��Z��V�LR�$�jdB�����!�I��3��7|4t'�>�;��'�F��|hWg��w�����Ǔ���q^\��y���`Zam�����eD黖5:3�����Q0�NeJ�n�V��� ҙ��?q����-�ؔ���ʭ)V�m�Qk)P\��T�Z�Ÿ�be�h�G2S00�j���j�V2ѡ���kVe̸���jRTQ��%��c��Z���1kh�a��=���@���q�m�w�c��=�Ǖ|)�Lv�ȹCiG2�i[mh�R�[���1�ƹRᘦ��3+�ĩ��W-E�R�T�ܥ����-J�m�l�˕0�2�R�Z�krְ\��mj�i�q�8x�!�G.ۄS���--�T�J��X�Z�4E��J��YB��m���U�d܏d�r�ێ��2��nQ�p��h�)T-�-2�b���rc���c���kQq�R�eZ,TkE��j�JZ���y8Ì탗�!ېwm�qjQj*5i\�b�j�����Lj���	j�DE(�j�jʅ[V5��Q�������e�J�-VԵFۗŠ�Ym����Z��[mk,-�+(�iK�(5mUdZ%J[Z��Ŭ��Y�.JER-cA��F�lckډ�r��HBMk�߹�(����H$�ﵲD�莃�B�Q%�-�m�ә����ݪ������$�^v�����5�;q4o&��,��J�Z��J��+�;�	^gS;�78$ˋ̚$��P$�okd����gA�a9�wYx*!���B�[���9ڶ�=d�y�]k�V@7Z+1��J͸�~���Q��0�(�"����$�Nnv�|O����c�I�9e	qcJ�^�I����!D
�
�2 ��(l�s~��o\Ìn��;s	�w���A>׹͒IyW���9�H��\H�H�L�&*�����ͦH$����lU�qD�33��N��Pb،0�(�D���r��K��:\��ܥ�I ��m0H$mfsd��6��艩�u|:-�a���c3�k'�U�Vv�v���ñy:�}�7{��0/`�k����KtjA�l*�ӈ���ax�M���	�u�#�Ĩ��T)�߫�|t��^���qaiD���a��ͯ0l��}S��$f�x]VWO`$j�.K7e�Hf�,t�k��7\��d���י�����1�12$w�ݻa�Vf��l��H���~��\�X`���l��=��
�0�:k.��J+&ywv�U�����z�5�|l��|Z���T�"�'�"N̙�)�L!�9Հ�p��H$���v����3Ă}��͒E�}Rz��bR(L�Bl��v�].Q�s5�̿�޺���� A����3>��Ă�4o;u�\rbJ'�"f(r�(x�w�u�V�����[� ���ԃ�}���\^!��7��O�z�ۼ�z�5�c��ɗ������.T�˿��`�P
�.`�"�꾦vmΛ�Fo:_k@��A�T��������.]Ƴū�°6�����f��dvm������ۜ���p�p��t���*6�ˋn��mō=sr��v6��d�V��΄�<�u�nv#��ӽh��.J���;vu��c��a�r=�xx�dח�O<rnG������R��zf��6��u��iv�&�=sۗ��.����Y���م��*�X7���q�muͬ�>@�G\v����q`�Q�=n<�GK���]y�����Z�3�|}}�_�6S!4����a�op |<*�A"�{[�ܙ�����&r��e�ă��b��\.0��
fD�y�a�0t	�G��DD�VH'^�����9=)s{�U��5�l��H�Ę�T	�L��t$��r����nGu��6v�=�$���#���ZO�D��"D��L!Cf��^�ᅓ�摆���;ݻLr�9����44�h��I#k*R(L�BoŽ�~��f�uteE!<w�(<Onn��I�����N�ޭ��о 3�B�!���nyH�h����oW�=��F�Aٻ_�����9�O�D�p(˺�I����$�ens`�YԚB:ߌ��H �nv�`*�t��LB�-������ثJ�.sv�s;U_3q�s��(�x����o���b��|2?=�n����=��4vf��rغu
}�=��gG��O����I����>8&M�B7R4��zO��V.<�Ǧ̉�uS�A'k3���	"榄��+���` �n���͂GGVb(S
!�t����lg�{�	.��H�f��^hp��?��>���cd �x�h瓿��I�W�P'p��*�'�	���l���{��j[e	_����,)|��Y�4�e���q;���3d:[ke�:�X8�3��ĉó�*R(L�@��-�s� �f��M����;PW9�s^�3�$�������� Q>�1EΩ ���	v´Rw��$�ՙ�?����Q�j*��V�[z#�̨�bb�l-��� �3yRI�ͫ��\�DҐ�w�҉s�{�k
�5]��|)�k�YJ�GY;�h�d�t�ݣyS�zgw���g:����ׇ�FU�yۨ���r�����<�k2�Ď��6&���$�´\�A�L)�(���^ b��Y׾$�n�$I�7�@�{7��w��o�m��`*ۼ����I%��ΜwBA7���ˍ��������?0l��H's{i��/�l�5a����UU�ۢ0mmp���C�u��R�jH=������ A)��-�����SH���4���7�@�}ٽ�����Y��]s`�l��zzE���0�2A�Bk{�|E����'�>�)��h$�F)�� �O�w���tT��.�o��$N� �%%�3��ԐI���� �\tG^�u^q p��zA'w{[�>w�c�̨�bb�mF�9\�<�$�x�h�u'����٭��F7�ș��+Q�7{��hW�s��w)��
��S/hƓ�I���\H{(�G�7��y ��S�KsA���Zwo�l+�yޗ��Ͽ�f}	_
�������K���Q2$Qߪ���5���؞����y�v8Z�q^$���lO����e��S�4����{��L{����[�+�zz��hǨQx)s��u�[��2\X���7��,��F��t��	 y��3�O����e	b�D>h-=�}�5�	����"J2���&��O�eF
k:�.�3[D���l�1���ܗmq��]�ʊ�.����&fI04�y�M��L�|�c��_t�۝L��a�Ò ��}2&b�S��+���:}V럃$}z�$�FWf^�����gfMyx�_c`�;�1�&b%B�JD������ �y��56�A;�\�$�����W��:��jmm:���C��*�hD��W-��qX��������ܱq�Z��x��j�1�J�tG��x~u�s�k̹�f`�?�޼��(����ͣ�3�~Xq��n9�]�.���Ct�]�v�-Π�j�c�ۗV�뮄�C%��nA6|�u�b���Ox㳎g�a�T�8u�A�������]�5<��8z����ݫ�7+��H�.�v�����nm֞N:N�T����S͊��(���`6�C����:��U諶][n�1�\�7=�*�Џ��9ˏ]s��9�qƜ��T8�"ծ݀NKnKխ��q�8�9:��Y��&\u�޷�G2���a��}�8��.���c�!�ݓ�nˊ���#v�i����2��B1	Kdv��⧟V͚��]���{n��I �}�@����ا~��}g�)0s͔q��	�6n��I�(
 ��K�gVܺ�Y���w�?F>ɮ�u�(L$̒`6i���vgbP'�x�YwOĂA'�d��۹�vi̇bؤu�s`���"��dL�x�;�+�ۚ�w9�&��fV�N�x�}�+�v�s`����� n0KM����������q�v�ɞ\���3d��ps�:ɯ������ʑ/�Y�m��יTI�ns~;t*:ԉه\�*�	#�eQ(.�>1�*&��[�9�jڮ7m��F-�Pu4mgUn�]-,䤰�gX��d���ɾ���^��Ӹq���`�8���ɧWsjR�}L�ܚ���K�H���߶|*��;�[X����~(�<n�8\۬��8f$�Q �L�4��u� ���~`�C���o7�`�H�{>�u�s`��$��*��!D�+j�Qƭ��N�>���D�G�79�I9����uR�sU,>uB�����$̒`15���=�Bs6.hڃ�$�nM"�s� ���l��yvp��<td�5��|�d����\�[OK�Q��Wk�A�2	��[�<Q�񇍿�q�n�2I#k�����Y�"�ȠM�f�K�&&�))H����l��^Ӻb���	9��߉$mwcd[\"�`]y�:����C�'b|b�J(�S�$mv�2��.;r�X���]�N4:���ӊ���3�g0g�;6L��- ��࢕��*�T���w�R���y���������3�	n9�����~��$m}��3�+&"L������k��V���;���� ������Au�u^Ne{.�&/�$���Ga��9����p �n��c�s�s��xϯ$.�q�A�"\�Î���B�Pa ��Q��%�:M�A}'�d.�y�q]���ㅶk�v�p7����䊒D��LY���H7[�L�|E�t���S��jz���lVrD�$�H�"fh������'+7�YF�����I���	�E�uz�1׸Y}�}����o{"�	�Z������6�(Q����dp�XI#��6	�u�� ܄�O�B(��B}�4�>����2�nOO1���t>$�ɢ�{���w�՗� ���i7r����j��x����y��4��6�=6i�Q������[Y= �cǓ��Y�N�tK���=����k���L�����W����=T�R�'�4�3I��'Ă.�$W�����+#�hҳ�?LlH�ac`& 	�I�Mk��I�h��s��p��;��{z��1��'���C��|�$���h}ם�fT�d<�����l�Aok�dn�y"��&d��i�s�$��Q�2*���N�'���h	����H<�R�on \�}]�b�Xg$@jHĉ2&f�B��I=��L���r��<b�wI�oq��@.���}Q4M)T���pb�d�C�u��	��]�m$����vb�Gf8���eN�Uu!e؈���>Vb���U4*M�o;˴�> %�s)�6��p6iP9��ʧ�I��f7�R�k�I�ח1��Bٹ�"����q�����Ty�a�)ױ�PJ�pn@��{�>s��x��M�ǈ����H�C�6z�z��5l۾��8mv�Ugg�;���VΔHǷU�н2nA=���Y����K/{��J!,[v�ӹ� S���^	+�^霻�ux.�;}�ٛw��Q���G͢	1��4�;l�z0'\N�U�d�l��[�[:pN��O���a�P�x*����4���{iz;B;*R�'f精��p����P�:�|u'O������8>=��Z���~>jzM�q��S��h<�H]��7�^������sy�~p�^ʤ��A�3�w�k�fM�ڏ.zD��Q)��{���Cpj{���D��5���$Ӊ�6�MZլA�q��>L�:HoYJ�Xy-^M[�i÷.ag��o�ڰq�$�Y����[Wo���z��=_+W"pp����t��Inl��	����*��MU�Ēf,>4ɑ��uҚ�eW�i	a�<����/im'H{��3�b���+��9�==��}��f��s9��G�r��|_����r�Oo��~�9� ��o�d�x/q���|5��r�8,^�M<m{�|J���6Y���\�Wz��{���"�;!}�ܽ�/ۢ���#�=�g���#;�n��ˏ�+�*��n�VT.����^�Ϸ+��%>h
�|�Y����9�^,�O�Z0�2q	y=~,�P��6G���}}=URuR�M^���t)��ahǉT`O?^~y�.��y�svcR��+4+j�Rҵj"6�Vڨ�V��[*��ڣQ���-��KV�ōU�Q[ZԪ%��e��j�ղ���b�Q�m��Z�Td���f[A��*QkYR,Ym$��*�U�*(�E(�Kj
�4Ae�V����M5D��*���Q�	V����ؖرr�	A�(+R�VQ
���Z��U�����R�m�iihPm�0���Z�VѲ�T��QQ��e���n��"��ZҶ�2��TV�Ҩ��J�,U��**�+��
�*��iR�XZ[,���ѥm��+����R6�DZ�UƬb�lhҲ�5mTU���*�B�U����W%m���e5LŢ*����mQ����mhZUiE�L���m�F�ieF�+-�((�TQ�+P�mV6��Rˣ.QP��R$e�V�ƭU��*V�TQ��
ҵE�m�KVҋZ[jT��V����Em���E�F�Rڵ�*�Z�-�i�ST��DT[V¶#�Ԫ�kV����+���{�uf8�{g�l��1�x9����⮞^.w6;�H{p��*m�7&�4ⵎ�s�8@�^.�{4���덷;��4Q�	��ڝ�]�L�=�E[���up�A���ݍ�P��s����\{>��m���2���;��{\�^�v������V+%�`=v0G+�n ��=�1�`W��rq+�9N�u@�3\2����]���\��hj,ͮ����i�������v�n���ڃ��j��<u;�����9v���=��؛oN<���<�ێj- �n���r]�űX��W��k�N�'h�I�cd�u&/�V��N]猼Eљ��;n6���H�pq�	�lx(�q��ڏUN�&���s��;&�O��\p·d�l�+9u�Y멫ے7����'j5�\ӎ�\/\�ߗ�_���G�z�e��S���=�Pua������n�Re���Tvz��%�e֧byu��n���uv�[]э��2���ܽ`���۰g���n��,��;u��N����m�3�Q��%qԻ���k�j��r�q�f�7����[�-e\� ���Оy��d�ժ�ʆ<�=6��,��v{��6 ���+R8���+��ȠrX��J�{�k�N[G]n��gq�ti4dw�c��;�Ul�8p���b��O���y.�X�qnݤ���~\��c�����i��ۣ����rМ.���=:[���$v�ݯDx�K���k�;���뎮=�����Vcg����ۓ`�}v7n+fu�����j��s�v:}�ylh2=���q�Jj�5;%�JmΒ6�-s��l򻣓\*h9�\�s��N�)>�t���LnL��uغ9Sq�9�z�w2�ԫό����ۊ�
cv�ٴ�%��۞gX����W+�7m�踠օ�c[�[�ݎp��
�>�t[�����7Z�a-���W�B��h��:;�:^!�<���g������a�ٺPݴ����F�na�e5�| I.]&e��1�hp�j�E�S�r�[��2�yC�w<��P���b�q�@�g��˧lll^�#
�2�G��ۅ����Oq��<Nِ�X�����9�ݴOF�c
��bO��ƺ;�v��������߉vE��]���T��s1X���7W�xR�]p�A�F�ay�Ϯ�q����G<����m�"��KF�N��њ��6�]]�cn� ����Nۖ���3bv��r^^��sul񮋵�b7UC��~�;��%EDJ�iM/e�M� ���j�$�Kڻ1�5jZ ��9�m�]��w`*��D�D����jG���D�ȧ��8�L6�I+��&��Z{1�$�j,ي5�r������ֈ)($I�$�p���uݤ^Kfy�A�6�j�{QN�u��� 3{���o�iQ7*n	�"j�R���>����Sw� 9�k� �s�� V��Y�/��r"#��컈�}�e�MP�UK���Lb Z�pU��;���3$��wv �3J���z�Kj���>�����w��U.�9����{,9�ָv�`qY5�ZדoK@''���$��8��Ӹ�Nb����PH[��a.:�"m�LK#�� 	'���ȏ~4X`ax�x����o����<F��������켬��r��>��q|$�t�q5\L �d��t��u=�V&�!�I�=q��\��EiY�[�a���$�KM���Ȁ%�de'��IYw�b�&.��NL���n���Oͭ$+�#��Jh���w} �A�����8��:yY� vN6�� \;�ׂ��ل�)3$���3;��b7b�A(wOВ ��t� ���mV�]e{c�������6�����7�5P�U?4�o� ;������[�zN��X��w������wa��˨�J�?l�3�<8i��%��`����}�n�킭��M�S��[[Z��֎7��x��b0V�z��7��ԑ�y�`���q�o�bq�;�:ܐ|��Qg�r��hL2+ [���ZA('�֓;9Mk��}S��  �x���wh�����~^��Ni���/oM�F�?���� �?�(��!@�	k�љo싱�5NEx=����NًG�|�u�L�6�]5JW��<�_*%w�oyɹ��F�{&6~������*��%�\^�x��~��w`/��<QQ"���j�Zױn�����;{/� �v�t`@}{��w�gl�u߱�^+܋Y���%ud��L��L7��bȀ3�s�I^��������"@0��Q 3�������?�����<>W��n�}�F݁�7cpѺMͻ]k�N5��G;btd;^�G7k������7���ϡ1���|���+ �������9��Q��[��+��=�@UB	U-�ޞo� g��[�ͽO����v Fv�x��X������l��U}@*��)6���.���G��D��)3��q�Na&�{���@�W{?yC�4S80�i�O9����]��Ѿ�[RA+���&����D0���������_)�=l�z�;�3N%�>��wytjdo@f��34�6����S�p�e��tHL]�Lb!r��*дxh�TIݬ�����
`�������Y�%�y�w䐙1EuED�j�&�p�9��iH �#�����S�T�}.K� ����� ����H,=x�-�A�}S�S�����L�����ܓҜ�R6m�㚺�Ax˷N�.�khT�"�j�*)R�[=��v�� �LB^I��u�k�QŚj�F�1]����8ܓ����2_R+�iG=i���,��$naۘ��	����K� ���I�g��3ǎ�K�}��^��(���	T6��O2	iq���$���9`�(�]]�^턀>3vu������o�z�U}AS��S�ھ��NIȞ�Jh��S�N@��/D?�Y��wK�^���6ⱴ׳�r�κ�hP�U3Q4��n4� ����ۺ=���B�G�{U�w*��H���u���w���J�,�&�؊[Z&�Ju�S���s�X�dp�	g��m�����˹��QA�i@���KdP�nmXf�X��:����w��yL����@��n����`��P9�8m�<���չx�<sf���nM�nY�\n9�bv���1���<��jCeՃ2��]v�ݣ�u�lޖ'�ݮS���.��J�%n��n{�!����p�:��r6��m=����.��w
����e�l�Olr0<�igcv����Ƹ��l=��Ǳ�ͬm���@�:M������T z��c�<���r�m�Gcq����y�9�Z:Gu��3�WX�5i�t�`�\���ҺH�"&T��G�WF7	$N��a$��fw]���F�L���9�D��o��V��@J���J%9h{��j�>td��T��� ��מ���n�S,��lL�tO�r�H}9J� �ԉ~aQ�[�@���� �OwL���i�؈�q�Qw��AV�U��I?�X��^;����럳m�߀z߄��n�����z&TS:�㯩���,J�1蘑L�̻V�t���F�,�׾�u���!��n�]� g������֖��
�$p���G��T����uۥl�ۮ=k*s1�g�C=nJ��ݻl���~�4(E*���^���_��n�;V�gN���Kc=��^������	!ۻ�dؙ0��"`��S	���nR	
2xoCꃱ�w�w�/�;������'���*���-Y{魉�+p�Tf��}�����'i�&�w�w"�rS���ʭγ'~$�庬�S߷����>��Q�姱���=��06�H)@&L	&F��=���w��u_)�C�z�L/��X�@}���w�����7$U
�/�G�TǤ���� ��wi �(oF�ZG죹u�����]<�����ڒ��k�T6���9$���SC�V�0dӳ�$;1�ݠ����o� d>�׌SaW�n���q����QN9d���km�8zC�����V�a�r�v}x�Rx������:�iG�������s.ՀDtn�^ !�z�,���SN���� dv�x6l�&�
�
���h:5�O������Ss����";5�C�� /�]�s�eu޲���������$�>�ߩN�a�	$�r7b�mw./2�d˷�wXڷh,7/������5�B��u��5ʰx�ָC4�C��kn/([͌U6�w�/���{n��|  ؿ��� ���mxJ�eD�L�L�{{�h�����<f���D��c�� +�޻Z�a{/T��8�m����TŁ$U
)K��=�'� w���ڡt�ݧǸ� ��[��##7��>+�޹>$7]c?Qb?���� �	$ٗp����v�������������H�����%" ��"�QwUԒI-8�$���޻%C�[�ɓ��v��)a獊Hd[G��fd)���ٗ~��\X�gvI饸�w\)�^����W��v <�����x5)޹��P��&p���$��ӗ�my"swy߭/$L�{=Ur���u�|�Y�L�/;y��S%3�d�3&aD��k^��tk�:�_Dh*���� wo]�Z��롳�M�br����s�B��1��S=^]��^MS��K���?�����0[Ы��#Tx5{&���g���1;y[-���,���� y���"3{���Gτ��d��`4��׿[6K�a��t��s8�n�QfwR@�u�i/��o]�~H��ڒU���@]����_��|r���B�^9��/�9��륓c��k:��ΝD�����}��&	��~~w��b���������L6�}�M�p+��~�����Eo*�Fd�>��*�A�m�I!Ha��=]�b���� GF���F^��v:�D�ΰ��E�;$�3&yT�o�חv ��s|� N�r6w�n�3���y��q�:77�Ɩ���
T��	�������#w@ ���Շ�}�f��`!]�>���W]�8̄���d؉0A�D̙��ƫ[��I���9�{i�7���� tnkx�+��4����cZ���o{M�����R��z9�B*�
��_"sH��Qr5�*ō�Y�U0�wk!6��*thT�Te�pl5Y�� n�� ���9W�`ԭ�a�=�n��;ri���t2q�n�U�pk�^�z: ��ڣ�pu\<�f�;N�˓�99������aӼ��v����L�r-����v�ol�]�nެ<�;&�����\p�V�Ц����Wj�˶���c)mc������l�c�r㪊�uu�k���[�ݶ���ط<,ci�k/7�=W\r�8���.ǘ���6���k0�]���튀�93FgnɈ������JE*"�UD������w��� �ͧI�w�L���N���W�v�@#cs[�x*�*l �AUA���x����	V9����Y 8��M  ��l���79�[����n��H�JT��2�l��m� ��` ٺ�9��n��G 275�R$����m!�m�A��
<�$6������=�)G	�u�$�D��o ���뾬�Y�M0���.�T&Λ��*�"�%6�m�؀A�����l���tĲ]Ց����[w��E�7��J�s}�oh�v�.�үk,a��΅�mZ��WN�w�gR�j�[���?$��e�U�Hcl4SZ?a�w(`|.��  ���@��󈾜�f�1,���(��JE?E�$-?'��v-$�m������bBXV۸9e����{������"�p:�ͳ�>�od����M݃�wxT��ʽ��=k����{����ܶ����� fw�n"�GM:�e<:�;ܠS��6D����R����l�������e�3�4��b�����[w��@���븋����D��U2�o�O��;��n�o}U8| )�uD�$�gw]�H�ܷh�ι���N��q���Cb���1"yLHmuu�ش�H%ڷj	��UՓ��GN_��"����� �7\ñj��{Ңe�yבWs���/;��V�O��iף����/agq$�B�U���1(&�1��̀ ����� .��r�OL��w�6�ڔ+�m���n�u�������fR�����5�@�]�v�j��
��m$J{{��"Oݦ)�f�}�.^��WnpiB{��B<LϥcC�޷���H������:L�%��cfc�B�Bp �,{�E���O��O���\�㎢��f����c�d�X[A���g��5Ou2
��y>������}�R0%�����$����k�ߴ(��/��y׾Ґ^�����+��ˈ���7��3z�Q�$���	���Nڳ����v����>c|���|��rh���
Ƿ�:|���\F�3ܰ���yY��?dz�ֵnk�;�%�w�ܝ0�݊%�c���s}�w6#<���s79؏���g*�f�7�eF��z�^�t���n]gX;�n�W����	Þ˩� 9 �z�=�B�vc����!pL]Td��a�H�P��ف9�zwffV썉���=Cݩ�7ZnnC�i
�>н�9�Xz|����!��`��� M�畧����h�O-��uk����ɞï�xq)��G�aP�[����17
!�wlUPݓ����ok+q�W����@�2�x��^�d��hǧ)����=sL��o��<��۔�[�y�8��
U�2j�Ȋ�d*z����[�=wL�,]�/�s��\qjP��2)Ѧ޽#`��ٝ��e�0��I��Y�����eH�ذv�Y Ω4����vg�ח�ہ�ݹ�"�mq���	A���$�4&�:E£����Bs�3�^�n�z��T���\���z����}[�3��U��o�P��ġ��=r�'���7y���SC�Bׇ��bFc��3�o,�{�ܗ�b!p)e��U�Wu��|�� ��L���
��m��(��Q�R�Kj�Z�i+E�Z�ԩm+Kim�QUZ�Q)JB�l�-Zh�l�*�@QV6��ҋm(��U��aQ�ծZT�����%bֶ�Ub��լ��[F���VҫBʭ[,R���-,J�%�1�m�UX��EffTR����1E���H���
ҭJ��X�h�mm(Te��j���J�m��UEF�E�-ҕ��U�j5���Q�cm�G��"���Lj�2�J����F*ԫm�U��eQATV)[h�bT-��U3.E1��cADUs1����Y[EV"e�EV���*ڶ��[KK*(��*�\�X"Eb3.Z�6���K�E]aqDQKD�X֭j��M[,[J)YQ�5(�m�4�PZؔ��������"*b�+��K��QJ�iE�QQ��ԥ�Z�F���-���DX�Z	j�K(�bXk4�+��Kh��کT�Z0Ƥq��eaV�4J�ij�Ӭ�2���\M&Zi[VY�	%��?~��m(~���v�߂r2���QAJ_�'��y����oOP �3]�I"t��K	F>�3��;���$���w �x��U2J��S*�Ɏ�7� �C�c�轪�Zr����$��v�ߒ 275�,}�l��ۜ�&&��pX��`�J�k�3k���1�e���cqɮ+� ��SxX�9<?b��o
XO'�>�2�X �ꆐ	 �c�E����*Χ�;˳���,c�[^�:Z��I���@o�������Aޤ&��g62�� nk��>��aA-�
lp�f����:$L�(D*����o�� �>�������mn���7P��ۭ��,}�� `OhR�S�Z5�y����8ȺA�T_?5� �����q�0��3�n��m6p�Ɠ�&K��^|w,ڬ���.:��3]Jx�l�Mv���Dᝒ�Ex:����ԁӳ���,s�*��������_$l�m:Kч�"PU(��?0Oߵ�$���yڵ��D��w���5���H�y�����wh6)˩Uwo��(&��W��z5+�y���c��Z�h���֊x7GZ8�\���D�D	�& J}���$�#�cM����v�<߽�*�i��ۮ�Z�`]���@U)�Q4�H�u�L�?h-�٪�I�H��tK	fv�v {�����}��f��M
&*(��S`�}�6| ^��qa{N�2}R����M�TF-{�i2���lH��P�"&T�XZg[W���3�3���M� wo]�� �=�T磆���U�稓a4�/�Uf���蚑T�p�׽w�� 2;w�x�}��:=;]�%�����݀2;u�ܶ;6j�Rqy�٪�G�f�Fn:W����u^N�ю߬���������w�H]h���i��z�__ߘJ�:{4�[�61�pF�zw��g�}��~'�8i%O�Ѥ^:w�<�u۶k'��Rv0�CjMV�-�l�N,����z��W鬛�2e�/\yԯ ���ļV��vq�����H�v�D:��s�m�܆��嘋<�0�"Y�ݞmt��q˓7"uc�I/n��s�X仍�ϱ�r]��8�[����؋c�<�Ls�����w+�H-n�3�B��y��vxKOg���m�uv�G��cD�7F:]ۥs�2�d���tU�v�(&�*)���clH����Ν�/�W��QSe܊o��@��w��3j�6����Dʡ�O�� ]����5F��k�� >��n����u� A���t��ճ����UnrL�\Ơ*iT҅SI�w�2�X �t��T"'o8u���1�K7���$�,ʃ�b�E��0��M�ݼ�7��vNw�R@��nҲ" Y��倐V�t�y�J0�ӌ��˻�U)�P�aL�AU.:�m���������t7
�}H��.�"g���!_~��J����
 �)aE|�	ԶЇ^��G<�t-��@f�]���''�m�]n�ۮ��߿>�J�R*�m޾�@q��I}��I���j{99
��u��v@|n���	�ʛ"PMDTR���t��e������qe��@�L���\�5�^�ݼE	Yy�{���۷u�{7����y��$<�۞.���((�!�[Ƒ��%���x�}�xM��sq���7�� ·�d	���B������V����3U�T6O�1���U�I%ō����$�̞d�I��mQ 
�c�E��j��M(U2(��ۗg/}�p�R');�%��6�K���Q�n��E;	/��nR赗&&`Dzd�fa��ݼ~l����wd�9;��^�z,- �k�tKIfwu�=��xs���I/�)QS�GGcq��Lf�n�u��]�,��;h���ͮ�ع��{��97-&��o�|��ҐH�����A,��l�l���dB�趉i/!ϱ�f�# ����6��� V�i�Rzg�\��b� �ʢIy��vM��1;���龈u��{c�l@J	T�(�����Ā��v�;��k����Cg{	�T}w<�[��3�wk�V}=M���<Or*��"��iZ���p�{���Á�
��%{{�9<��t���W���$�!w��� >���w�~�"�LL�@SS+z*�%.c�gq�bD�����B@}}��q���ַ�ȏL�#���a$��7D�N�̙�LH�
w�.�����ɥ�yM���P{�E���������9]Q>����]��Uُ��\�7�QљZ�5ۂz.��kmk5<�:�:I�;�z�o�߇߶i��DDUO�޼m����Ȁ�:��<�֭�Lق��o�A�vou݁���3�I4k��k�E�R�����b ��3�Y�)9�|c'/�%ɳ�}��ɐ1|�E�\��:Ie�m1�E��,*���4���A$e��Hz�*l@�%D�!�H9�uf�/�j�4b�MD >��wa�	�N�`| �ݎ�b��g;MZ�����٨�ԠD[B��N��%׏���p)��'wj��ځF�凳�}���uR�mZ8TeQ0�3�Y,�uz�L�Q��<��]�����%����2 �L������6�"IY��{�={UC4����� ����D�����cmB����(=`�J*p�)è�7�G�ٓ�N���=^Î���u㱛�ݶ�Yzl� *�*j"*izm��A���j@��/���t�-d�_�o;[� _N��6c�19R�~��
�[@�3`mm_F��F��i�7�}Z�	����I����(Y읗].�NbƳ� ��MR��uՠna e�}� �2�bv6��@ ���o��W΋ ̞ȔH��`��{}ֲ�6�{���A,�sD��G��Iw��w�s�r�y��馒�1�pP�2A��� ��%���w;�OM�?(���?Q�2����z� y��v��B:2�����7�3��ZG��+X��5G�u��K9#�]O��Ë�n7ۛ�p��!jy��ij������ٟ-0�:@�[G.nfH�DVw>q��c<~l�����ڴ��js�u=�^���K�-���1�K�N�1�6�$�0�{r�Q�J���J�l�8aM�����YE�L.jR��$�n͞.����Og�Z�d�nյ`&�h�W;�,�4<F�W Y[q�`�q8zdѹ���p]��vc��7	�p�c�#�����[�,z����� u�����F�.����<s���C��/#�5ĺ;=v�v��S]���)LU�T?�x��4���䗯7��V�{xU�|�炛ۦ� ����X�5UQSQSI���x��$��Nkr��N��M0�-��y��^wsv -�F{�W�U�^]�i'3���m �l`����_�>n�7� ��H�qR�sb �C&�4IW��wa%`>�&0�&�$p�9맗T�YDA|� ���π@^wuݠ6��u��>Y�DG5ն��=�(� ��Q�,��������^h.�9O*Z�q2�
+�ߘ���w� #o:�	���K���j��$��	b�Y�6�Ev���͈I&�.ۍUt��bx�=����|~&3ʕ��}�u��;;�݂ ����wf��ȟ!3\�D���n�Hc�[5�	��T�]^ĀA�p�f��X:t�w��\h�R��t���(�h���׳E�W�o��;�����=��N;����>���o�p�@o���w� ���M�+�ӪG��M��r{���l1���	4�7ݙwa�Du�ך  ��<]�wӴ�=鷹���^wu݀�73���>P���M�x Mwa9�(৩@Mژ�_� ��v  ;3��B��ۍ3}	�T���ҁ(<�&0��(CF�m ����o��[Nv�3.�����뻻H�;3����B籰����#uuRӆD"nI13'��y��3�u�������n��K[s�.͛�ve" 
3���m�	$�3��� ��~ �7�s���{?9$$�?[���UȂ$�`��Hs�TM�{�n���i$�Cs6�a%�\�:%�I�8ރS]ϲ�3]�-zϓ)���gA^�� .�v�w �7�T������q����È��.���u��9O����g���p}�'	�\Llb�38��n�h�����آ.F�r��'��3}�O�I ���m	 +���`]��DAT����i6��f[O�/�a��ѽ@ �n��DDu�������ʺl�~��Z�aݵ�Yjzh���iB����i6 �7;�ٵ5^��{Ҟ�h'��p��]n6� Y��w�{�p~����~��ߣ��kH<h��ݺ������b�����R�q�Og�vn�=r��~w�����<n˩@z9�-� �Y[�6 37��YUm�@��+#��"��=��'ve" �2J*E��m߭$�航�)n�w�A  Q������n�#=71��3���#���*��H��n���97|�����n䣯�B�ݘ��!uf{��3�������
`�����)�~�wD_�|.R ��A����3'��ۻ�M[�2~�����-��
{�s�z�{A�tbv�媩��3��i�+lnLhn�
��"6�� �ښ�M�pqT]��B���`e��DEM ��	�پw�j� �;��X���P�]�9`(��?D?���7�����r_r�fvO����Q��쪻�n��f㪗L�k�����E���Έ��^:/�'Χ����]��7nw;V d�9hE4�Ю��PBڪ�l%ݝ͓t*�3(�LD�Rd�JI]��ë�X�6�v��h ���� �a��!����4oc��>�~	�V��`< �e���m߭$�Y�:��I.2(rL��_� �o]���3�J���6\R" ���LM �r6q�����O�$~�wa�D��寀 W]�q9�nA'b�����[�̄$��!T���7����6��ۂ7�oion�`f����+������Ȥ�讦���Ytb�TK�ʌ���;�W�٭�yco^{D0�ևu�L`+"���obҼ{��wvD<�T���q[_��S��}����z�V���d7�| ���Gk�<��x���y{ciq 
Uᬏ_{7��z�*Di�-�=���FZHX����4�U��ku������[o*�r;S�03R�0�f�m3��8�@Φ�mM�7Bq�W��smM"�R�����,8!#�"5��R~�oMІM�C�-��3۪��`���u�\�6Dߓ��ܹ��(`��g�wW���{�t��6+)E���9�!G]��2!Ί��E�OQ�S9�0�*E��7���b;σ�ᯧ��x�G�$�O�ɢ�%�l3�N搬���1%���1P��b��O��	�ݞ\��/�sх����R�L� o˼gz�2;\�~W�wC¶��
�Pӻ���d@Ȉ�{Aٸ{Lk^2�{���t�ɮJ�a�|�w��r�ݿlv�����=y����m�A,uU�^��TE�p����ٴ&W�����u�}�/]H���2W�_���T;�·%�
��<�s��*srp�BDEZz+	�Z��k��!��`�_"\Nl�5�{|V�.�5�Ś.��lT^7˘fKyL<S#q�>�nls7Cz��W_������z2�������K�_t��G��^ɺ'?}��m���JVȅ�� �b��ƪ�Mc�0.�b�[������k�':�Cx=}N;�waF�%����Z	KUbZQx�(]%1-4�5( �c�*%M&*�J��VԨ���m-��"��k,m�0��N8���D���%h",�jWWTDKi[mb�X���4YEr�mTh�EKJ�Z��Z�Q\�h�U�����i�-�5�B��M5Q*5�ʥm�m�1:h��64m�k-��eAZ�j��Ԩ�* �iGTTY��[*R��Qm��Kj�����*4eb�l\��Ҋ��e�iKh�ی1���
��eb"�V�UЕEkP���E�ŭբ�J�kH�en�Uq*�u�	�6T�J�J���TU���bԩZ�D��FUcl��fQ��ڰ�n&e��U
V�A�D�$�ZP���2UE���PF���E��-�ʃ-�1E�0kU�EE-Z"�mQ��E0�J�.j��Mk0�QPE*�ZV��k�-J�U���m�`�ak,e�V��M$��ĬE(�kEQR,UQ\�qm���-e��j���+*YmE�,uLUb1*(�o;���%\�feq�#ӣ'0��vv]����֋�j�� �j9j��k����������'<�q���[���ώ�r�[v�kK����!��m����]� O6ђ���)�V6�'��ы����&���V��q�vݶM�j�����MrY8��i�}�U��:۶^��wZ�=����2�vwa��t�,�@��l��zwX�s��k���=���,p�c��y�k�]�0㱍�n�w�v?��g񞂹�8\���s��{!q�q����f��5���jV��s�!�E8��8ɓnn޶���]�ێd� ��m��uv�	K<n�7ۙ9Pg�l�Q<�/�2�����A�ď�9:vOӬ�F�nlX��A�@��̮yݬh�%��:+\=� �p]���V�N��j6�N�^�ߏ�ߝ�k:���[������l^���&x��K8zS��q8�8�(Xs�sl�<ɎϹ��íb��mi�޸��۵��~~[v���v��pi��ۊT�=s��A�l���X�C��]�n�n���B9w�yǜv5��7������wG䡸�纯��/N�ݬ��n:��:7a��κ�{������=��w⽠y!�	c�Y	�.��A�Pc�;�;ݣq�o	��Y�ŇrI�cNr�7g� ���O6N|��vN�w+��Y�K�\lt�&=n�m�N\tl[n���z�rƹ۬Зr]��k���N�s�Ž.-���ʽL��m�nݬ�m��u�8�n'!l���;��n�Y��ZeK={
a�㓍�ct�[�g��zO'm�2v��r�֮�6�y��;<7[�=i�.�lo=x�u��h씾%�E��lѽ��{v���wk����Y|MWP=n��v�w��a��1#]�ڌ<���n�sg*�"��v�y�:�iL�v���Bs�eM�uǶ�q�ګy�u��.�._	��x��&�y���OWT���ζl���݁���=���spt���nΗR]Gm���v�������0L�^t��w���������[��nqlk �7�.��ڜ��n�,�WCӰd��q���a8+͜�64��I�\�۹�w��8�c�݊1����λpq�iw�[cu��qt�lۨ)K��'A�St2����[��tU{7v%)`�vٶ(^3[��3ezc`5������5�H4a�����ݩ�CɊv<�nX�v6mN���=4�.����W.3.�v	�,M\����2O	E�S���.[������@.��w����nOV3]�iśLJ^ȵb	�(A���M�$7/�'��#Xpz��M�w�����@�u��S��4)��ѡ�nz��$ T3�`���Q �7K���+��� �ׯ5��Vϰ�� ��9�D
�͂Q4wfPF�d��2��θ�k:��4����@ "�1���gw]���Z������7�?E<�)'�,�~H9�~my"w7�߭Nd��y;��\F�Oc������� ��n�=�C���Jg=&~=���,%���B�y���i��s��e���]Z ��G�Ͽ~+�����U*��%ߺ����m��;��!ꐚ�[�z��k/�T@B����$3�<<%RO7����p�"�389�5 qf
�PF��P.p���d�Ԅ�&�&���O�KlA�ݓ�{���/����6Ő��m�`R��9���Lw�|k3�k�>3{���_�Q��dx����l�̇*��LRT��v^4���w��f�v��t}��t�Vg� �37��P���$�D�K���o.꼆��w�0󻛿�H�̎dH����U�
J2�C*�~i�&�ERQ
i8�s�z�	fOy�,�t��ȼ���3[�%vwuݤJf\sb���箝T�\�Q�|���`�����bmƭwt\3�q�<�'.+d+^�H�<֏�����x˿��v�6 �{��`�2����XD"[�rd�����nn��B����3b����� �a�D��Ҫ�L�?&��]��wh ��RDD���f�_eL�1L���{J*iID��H���݂�w;� �@�/�G��b�*��,�黭�WKM�grI�ݠT��E�u�=�D�����,�t����T�K��^�2�K�^����{^z���L׽�"�{����6�͹�9P�SD
jS`�o>�z�&��y�_� �{���>w=ᄐI!��U�9St�,�%�����Ҷe
�Q3DDG<�܀ �;w{~{Y*v�8hݎ����sͩ H)���7�z*6&\t��E�R''��-����<�-�[d��J����7c��I"II���t���D�"F�5w���� ˹�5 �&��^1~�fa�=Ű�'�9wN7XS2��Q$#�!�������:r�ͤ==�ӝ�ՀDwZȈ��7��d�2��N����3�uHU5P��T�Ml�I [Y�6F�x����̼��@ l]󨆐��~�]���bB@��d6u]ن#;����&���x GWc�Cn�u�8���_��X�B�I&N�R=���ŕ��W�}L�e�6�j��}��ɨԪgS�'�ő�]%��S|f~Kv	��z�q�m�黙�
E4@��8��w�Db��wa=N/w۹�dr@*;��CWW�i�|]��wh����Ͽ[�Jmwv\�Y�WM5��u�Z���D8��,iz]�;Z8�
o$=��s�߿>���F��GC��� e��lA}ٽ�vY �ۘ���++@�IHmֺ,��C,C#�p��ߧ TOW��uK�q��Tp��{��	vou݀��B홒WU�!�
I
 D�`U4/�� Aݽ�Հ����Y��e�$�Y;\$���$�;S�%B&��S*��c}�ruX�\�wr2���z�l ��> �w�>9ۧ5H�.��hvv��"�yJ�����M�oz�����:��1��99~~�˴�P���� ��{��$�n��=�`C��RX���{�_;;ݜWk��{��T��4Mau̓j"����7ԬV0d�V��V(4K�q�S��ctm`UXH��4�i�~o��acdMj�K�8퍽F'��n�Of��Qn�M��6��v���G9	K��:3nVQ��U�c~_���<�&�p&�6��wWg[�v�t�s�����X��%oQ,�g�s��	�IF�9�h��
ٖ\G����4��l��[��97s�z�q�9Y�<�k�u7,���run9�t��W�@Iӧ��[:����]v�wW��~w�\���u��tV�y�u���3���Y����m�|���ޞ�b5+߁m�4��	n�;� ���L(�<�ѵ�O�����d���ؗ�K��J1�)�\^6�)5��p7g��$^���I�.7|ؤI�v�1>ފ�.����2�)I	$D��=��v� �2.��x>@ "'-f\��f�S�I��$�<{2��$�!]D*�eM"%?4	纫��Deh�:� ]��v |�m� Ww�=����d{�/����vnj
�ME
�D�jW6)�Hm�?7�)3T�+�77��"�FF�6�A���m���9�&|)ΜX {
�E6@a���fW�.u��\�l���ΥN�v�����������BH� ȑG"�}h�ӷ��%�@��?0��N����P�;Ϯ���oC�U�'*�MDԦ�m�?�Kp/lSU8��-���q�Nr�S^#@�ݚh��A�l��X,��!3.\��-{�z���ݭ蝛����-.��y���U:]^>V �^:h���l�*e�>������P�qP*DD��t{-�0>�|� ���0��z��3�.q�o� tu�/ ��Lz�f*�J�2aV����pj1�D�^J�^��	/$�v�K���]�|��@J��<��n���E�"a(1!O���������,�շs5������O� ��m�vn�݇�Cq�S�������|�N݌��p2�|��X�ۍ��]�v5m=���'�vz�����;_�����Xm/T�"��� m�4؀H���v�����{<��v��Ww�l��E"�)J%E*M�����|��+������$ 
2�޻����iiS��ɞ�;wn��5�Q���$��M�oq� �7w��}�$z���	X�u��-.�u�$��&k�Z��8�]�8��}sU�"����;���I�~n;�m˾�FyH7�?L�O������"��|� @vn�ݤS���R"*� C:=���Fz���k�	��� �	n��݁�x��+�W��;jL$Dnm6����PT))I���z�ZI��)Һ£���u����~` �����:?K��xc���$���(`�ZC��3΋������i�Ǯ�u<�\Q<I�\y���|��}����ĭ� O��� 7{yڰ ::����U��vq
o��d{��v�W��栨D�P�f�[*;�߀;�*7����^�����4 FF��^  ���םm�2��ELR�J�T�D�;��ȃ����5��k")Ϲ���ڽ�g� �o]�{���8���@�H&����雲��G��Du;�iX��-6���X�=QY��������lmjM�rY��VW�	��ش|������r���#j�d��b8�+M�����e��N]l�|[�ݤ��q"*!EM(����[t��I!������o]L��m�]�a$���b�I�yL��f�M�)�2f")d�>M9�2P��6�C4{f#ڧ��Hv�Һ�ޞ�7���Ϭ8K[���k�ۻD����Ia$�9׎���}U��o^���	 ��׭���(V��P�"}]0�[i%[S573qR���Qvs�w`� Xm�@$,����ok��S�~�+�{�����J�I�&"L6��sb�$����	30��8U<�N��Ԁ@z�� Bμ�`���Q$T�*D��I�Os�u"ʜ�(`Ү�H�3��$�H_^U�J�w��Ol���Ѱ��K�A�ۤ���GLT�SJq���6 >�7wyݏ�s����Adr�$���a�J���GP��{���=��#5R�����W�OM���^1_aa���7��5�d)�dݚ��]��1�Ɔvᇄ��(��D��ژ��9G�U"L�2���5͒v�=h�7��e�,wc��;���ը�������\�"�,�
Tu�������^^Z�`λxc�r9�m�6&ßc��)��]���9wI�ƗNz�.8�l�{=��b�:��qՌ;��1�3��ɲ،g��݊{d�ۡה�p\EK��p~q�t붡��\H��������\Z�l�E[�h�+ ������U��ȱ�&;�u��e�T\4v��$`���R	3J���u�&,���� _n�݄�g�esmƎn�H$��z��;��i� �xD�XZ�z���Zr��qȗe����	$Fu��@{��v�C�޼�>�z�3�z�ँޠ���Q>�.���[b 3{yݑ�:�"�̭U�o�zk��,���כ�w`,��uPI
$�&����&-,/{���$5��Ā��޻�##s_g�{��U��-��|>:�I1J�*)Rm���Z�����Q�W�j�m��}��}��v F���[s��a�	%
b�ĩ�P���������SC\h�g�&\��΄�мt_����~�pR)�.y�6F��;� �t�C��ڗVE\�F�{[^ A�����Ut����DC���e�����}9�h��T���m"�
�݂�������Y�����!������b޺9(L�̫�����t`��k��ܻ�]�9����B��Aܽ�H�3wz��K�;yN�A.�ʕ��I.���D�]Q*dT�LDRp���iX �c�<� �.y��cݥoWFow7a$��{��p9Iɍ�����'�V�g�?��$���wh�ӷ�-"M���s���dl$w�v<��i�**�L�O�\sn��c/�o���.>�(���ۻ� �/�W�IY���d�{ ��R(�aRc4g5�yu�A�Fn�[7�GpɌs.f�9+���ĕ�{<D�IJ�*)R|nz��Z��/}0�.:���w�ܥ[ۗv�i��TmM�=1ST�4EJ�A��~�ڤ�~m:��}d@ݝ�1�^7H�5�9������d�	��	
�R �Z�O[�'�a�$���o��Οߝ��@m�g��k�;�罌�zWp,o�wM�H\�u�O��Ł���WD��%�WQ�ȳ��q���W��p������z5���9�G�^n��T��w���6lٻ"ϡV����������\�y��Ԍi�a�}��d�������p~륁�ò����3p0�o���kpr���I�'��@{N���gKðD�JCÙZ=}��5�S=u���8�w�!��� ^�fw9��/�T�⍫��޹��{K�O��u͓�'A=v��sa�u���o�!��n�T9��U�T�Q�ݡ�⇚�K�;=�Bʯ�.�z�pMo{��Fh�e�N�7��N��>���8�+f���FϦ2���lc[vb{hvm���1�璕�1�v�;�*G3�,����|��X4��ӻ�Lr?=�=�/�9�=.z�xv�#aR0O/LX�u�@�S�v{�7��� ǙOHCmH�F��*@�2���0h�k[J�v6��H&	QcvV�CBz�0^�۞�����ٌY�z���<�S~�f/ovy�����q\�z�|s�[9S���P��$��à
�&�Prӆ#
u�2y#�pvQ�ۇx�k*���}������Ɣ�qаa���5�K���yMݨ?6�JU�l�w����>��+��z:�S��7��cԷFx^ĩ"�����'{IV�"iv��]��]Gz{�F�L]��{qu[�nk�x��Q>��C<}�ʖ?\sM������w�a���iQc��ݬL�FԊ�uq�bUm�Q��U�օ2�h�e����JԔQ*V�T�"**�b�h�*�t����Ѵ��
V�m+ՖeD���X�KF�KZ**[,F�-�VV��`4�im��j�F(��Qb��Dh����V$��mŅh��mYA�m*Z����]&�Ķ�E�jU�bR��G320X����+Kj��R�"�]R��P�Ԣk)���-��R�Vڵ�7.6�Y�����fV���%�����R�3e-R�m�fk,L�*�1�K�,]Z�Ŕ��3"��is3+5�)-�cV5�ж�\�kQT��R��Kn\`���T�CZ֍.+(�+QT�[-2�*#K�������N9��n-�T���KB�����\��D�YFڹT�Lp2�R��)Qr��%J�j\mu��뿼���P��Y��$�e�7�H�s*B�C-=����}���VTI�'|��Y� X�0 W��v�!;�l������A�
�+�I��1#�Bfw_�����`Z�"೮�ez$S
m >���- 2c��ם�whf��yV���R�`�ТJB"$Kd�š�{q�7'V�3@��sbݺ�����D��U5J_$U��T �y������]� ���CϭĬ��x�o� @$d>��y}A%R�J�T��������d�ԩ�R/�f� 4��t�D��w` ���&�S����\7e��s�q���g�{���? ���X \�m���7�k:��C�o� �7���
U:\�)J*TH�Y:f���
��u�<�$�\i�������q�����ǔ��~O�M�"�w���혟ny�w�Y��<�.}�6{qz��nU3}����b�/�<[��t�۞���`{�/g^n�#�/)4�t���&`AF}$�25���� �f��kvn���9��|���{�� �6;7���E�xn�^�_�o�������awF����wc�g���!u�\g7�;�6�ϟ?��k�-''���q~��| v�sqi ���]Ѻ���-��7H��w���뉓B�2D�Ȇ���u��ڃ{T�7�? >�����Gf��@Mm�j��*�a���״Q%*D��I�O6�� >����� v�.�V�t�=���9���6K�f�,l͙�"��(&�)6�b��֒jʭ�w�z4 �o]�`�,;5�@|..���l2̊�NoW6JP.!1 �:��i��uJ1W]��0����"�H���Q\]�K�d){F]z��B����ܺ\�Zc̓�u1f�4�+� Q�)����rPU�5�z�k$m�M3��J����{}������@	c����K��u��u�Qr�$�z�/��#�˞f�GX�K@����m���ױՄ,����5�nۙ���u�=u�|�dl#� v��3��ݹ�ym&�^ݮ�,��:�sn:�_A��e6�"����.H��^yܤrp��5�n�/g�Sųٝ�[cdf�u�v�޺�����ݑAr�vl�+\�6m�Xw�^��h��X���l������]'����K��u��Ӷ��v�n����Q�I0�&�޾�Ii�ڒ�I\]�����p��A��-on���>2?_wi8̨�"�-b]����_�N�a���7o�PI{Wf�i����~�ITr��:���t�u�Ixs�ؙ3$($�̈l*=ͿRA$��*I~K^��,k�ǹ�$Ja����D.�k���:IS34���&ͮww�S�t���[�k��-�ZW����R�.e,���9�K��18E)*`&�
M���4��o;J�� ,�e�&�V�,$�:_e?R�/3y�
�7�ik���d�iH�u3*���X����[�D�b+q��mEu��h����y�`�3
DG���H$�d>�S� ������/���Q7��$�\^ct���&`AI(J,���uݢhp��V�s
;5����<���+ǈ��jѴ>��"(��:�\�nر]��w$�P��u��)xtW����| G���y�w`-�TunS���^
7��_T�J�Q/���o�@��7��E���\��^K	���ؤRI�w]�y[U6,x�m��:?{�g�䒳��!��G>i�@�� ���ܬ�~�zۢ u�h}sĔL�)�iCh��]ڰ��y��\f��O����}㭺 O�z�"��rs�s*0���2<�� 
UH�.wi��#&I1��R�3��j��������_�R��j`����^z� ���%b��,y,���s&s�O��i�%���͓lM��0D�L���YkKz� q�=����mD��h ]��݀�H���Q .r��sQ����)7��)F����[��l�Iy-=�RIa.��i������W�k��qY1h�%J��~��pa��m7'�n*D����,��4C�"IJ�)�_?)�֞�����g���T��K��$�����v ���ׁQkf."��*�T�_���Yީ���!�TE�޼�j��适6g�՚Ez�Y)�]�@'����o��j���J���y�;�k�^K��a���2v�D�]�w`$�K��H����ߩN���vbԉ1��ߨ��G���ր�#��ծ�z���}:�{�CD�}/�JO
E$�oﰩ�N�ln��| h�?�=�*�[�M���ۻ #w]C�*�&x�RR�&�
M�F�?����J����2�����| qۮ�@ l>�׈�f���5�ח~I
}B%Q*,������ $�� )��)�f����߈ F��u�;��Q"&�"�q�����sW�;�סּ�Q�t����R�H$����j/E�#d-=B�Wb]�W��򮈸31O42���OJ��/�l���}I���4��f�LƜ�7B��(�qZ�N��I:,�ٚN:�� �x�»X'[�7nw7�*�̺p9H��n�@�ci� 33z�������a�����  ���DrX��oC�H��n��n9�/6��#�^t�~~�|>N��%T�ET�Ǣ����1�������%��d���{.LᓛUԊ !k�o�w<IRLҘ��)S���V�7�^��:Us���x G>�L$�K3w��&�`��;#-��n.��ٛ1��R!R��H�w������vD�2"fb:��j+�� 	_c2 >����vyL�TAUJeZ�޹��[/�e��Iy!��S>��޻� 2;uůL���&xn+��H���t����$�Q0���kn����I-=�RiTI�\�ɬI[X�!��W��w`$�ۭ��d�*6������(ن��h1:X�#���7$�Z'�{I����4�g����5wu�v�E��Bbm������a���{|�;a�쮋]1�aj]�luњ����.	�Rtbc�{;v�v�|mv�Z��gv�=m���l��ۍ�(�>8��m=�i���5C˧//]�6g�<c����#����t��+v��<mc�<�{fn{�9M�ո��;n/W���4���5箖w]<�s�P�6^3�n������B@�JWmV�5�䷧	Av9�U�`��Շ������7sDAt�&Ô��k��4���e �a7�,+�������gv�`��;u���K����߲�'���ݶ�@�ݽwh2�VL���"L�*���G��ob��ɸ�֟��gn�ݠ2;s��DSGm�����o���cf��S2%��y�شI:wr���I-�ե��Y���0�u�|go]�X���P�ٛ1��R!2L��K��,���]oTox|F�d@O1ڰ� 0��M  H�}����\�4Y1�/����VPQIS33&Be�6��%�,/��%�͚׳�[A����dn�!���6)�98�ě+9�ᖨ@Vd!���{{�B��];j�=���۪-�����z���]5�{�U5 MHE"�9�m���6;s�xD	`�0fO�f�yww(�o���$$�O��{�K�T �`�M&g����ڗlv�X��������r<Q��d�Ft�s�C�+I"��-o�7��������^j��0n�}8����I��bU�.��ng9~�o��Di��� ������}3���b��1������"fA�D���u�� A���� t�Δ��wgobI#Ƿ)�$�/��$��;�"(FD���.ط�]�1��Iu��$%j{�I%���Z�t'�ͷI��pL%! fI��KN�0� ���Y�'N���v�{[�@$d>��@�;{��3;bj�&W;;����F��V"۴����uٶ��Y}�3U��!bGi�ФD��L�Zm�t C�?	 �Y��wa������^��I�ƶ��� �	#J9[���:g2z�v)C�W��D�i�9$���o�K�v�(\��q����`�&}&fA�4����D����ݢW����vθ�ci��*�n�]*9ѩ�dE	��x%3ū7y�[ޫ|�M�am�9�Q�v��uf�����P���Z�y�����ӽ�x$��x�(7{�� ��7(�$"�EEi&w���phf��voBK�i��� ��O����! �^��B��:#a!��ۨc{1�
�(�	"�89�x��@ �Ϳ?u�Q�����*<�� �;����ο?޺���2�C�;��S�����u�9��N�i]<�Mk&����0(�ǻ�UHM(�|��3��H7{�݇�|���ʽ�".�6<��|ٻ�w`)��)M!&`@�OyX=Iy'�b=[Q�Vq���"�w���@$tg[���}�f�'?r��Ak�4�sŶ�$�h���ao^uشI:s��� �6UN���2�����$�ݺ��I�:���`�&}&fI�:~I���6A��7���6�1݀3m�H"\[���a��z�b(\�e���PHȵ�\�u�I^�V�{����V�J{n�8=�,��j�]�n��o��r�m׌~�OM�HI�s��KlC@��y�� l[Ɵ��Ν�n� ���������"��7��SVd�|�~~]����v���T6x涒�i��m�q��I�8�.Z�Y+���K�߿y�GVGjT��n��F�m��� V[�O����Z��kY�wh ��o��W��H��N#a�����m��p���-��@q���� ��}�@t/џ��ޘJ����`�L��#�����I,7}R�A*�g65�WV� �##w^ H"��y���ª� �h����������a^Kğ������ ��:�`f�u�=��ޚ���\k��HN��6L	"bA�:a'�߄ fosq)��Ɉ�Oo"�.Ou�-$�;�D���v�]ߒ�z�~ێ�Z�7��3�y6�k��CI`���3d�f{�'h�u&�c��"���=\1�h�,�P�u`��Fc/����J���g]�X�<hR�{�j�A�w�K�x�1K�^�{�^�j���.;�,y7wo+�����L�װ�@�A�&����	2,X�c���啫��󃉉,���=;�vy����B
�F�NL��ۜpgiվ��G��N�����xCp��ߒ/un��o�ƶ7��������O�{�X�t��Ȳ�B͗�m��݋�
�ѓ(�"�V��=���_
�@N��S��A��t�S�[�J��s���\�q>�ء�s�i��>,�;�TDܾ��={�F�=����TEuʯ��sv�ɪ-���CǾ|0N�ݾC�g��9�gi���^T��Tn�W*n�p�����`UOs�¹}GQ2'�Y7:��I��5
��8��M��l	�s�y����S�q�r���0�+*��r<� �d�ˌc~=�N�w!ȀX�Z7�{}��ob��qC-{����˂���9!-���Z3S"�cW@ͭ���&ڃ�3F��G�==�Jm�>F
�o����cS��V|����Sq�}�Ĵ���t)����V���jɥU�H#�*�7>+���^y!��+.I����[�}./a��R���á�,t��׬���w�L^T7æ*�q�Za���CÏ���{*�r���/ݑ��i��ro�#샼D����^�x��g&�7C������j'D��� ����~�R�Ģ�mc-��9�V�ɊV֨�
�fR���ҋq�L��Q)��֮R�V,a��`�WV�1�Lʢ��W0X"�ֺE��Z�*�i���uJ�t�@ՙ���P��l�s1L[j�jʈ�Tb(�le��YD�a�٪S-�*��n\���b��2�Ct��J[,�DEWM�F�t�
�e0�l����LL��
��q�\���i�E(V�e-�� �V���Tq�q�Z��EZ�b�P�kB��T��44Ekh�-m�mZ[X1Ėҳ�EE�DQK�-�mU[L�ܦ7G+J(QYR��,�Qʶ
�uL�Ԫ�*(�-WMm֋����Tf6TQ�X�e��5+*�C�X��Aq2�Yf��у�����,Պ\aq,P���U1*53,Km*6\p�ccm����0���q1�+��T1*,ƣ�UB�fZ9j�-m��ն嘶Z+¸�Oޟ;�ݠ�y��h-d��H1�yWl\���8��*c�u�9����>ID�0g烯=vLU��t��am���`�M��/FpI�Ē�ѬY���)����խM+G,<qis9�qvxqh؞m��&^{q�:;S�"睻nk��Aj�Lz�tSt�\��l;dw6��U8�7I�`�����5�Ű���C�6�!�(3M׵��u[j��[k�u�7>�#�۟L�\�=h7/\��n9�;r�iy�qע��<nu�Q.��vݚ�%�n��m��m�Pl�Me6;^��vA��/=p�sZ�q������Tq �|��͕;s<��&�Q����q[�����t�ܚcay69��]�O\����\q�2evۣ�:�*v��o4s����:܋�z:.]��Y�-�=���t�v�0���յ�kq�W8���kO;92����rOOcZ�F��9���^�ǭ����t��k�����0`��E�凌��̯[���Gv�ݷ'�n��<n�8�gj-��QN�Å��b�<׎ts�{����`�o^�A�n�9�Ɏ��r�������{cap��v&�}ۂ��(#'-�*v�M�v��]�<�*vW���۷Et�qnK���:�urn˺�t�;��bY�����m%�h��%mnõw���4F�q�����m�A;rc^Z��hwY�k<���[M�u�\ն ���JGn��zu�����([��m�(u��u�i���r�u�K�6v���{)v��:u�������u��h��[��9����3tf<ԗ��8☔�e�nn�M=�qE�^;6Վ;v��ap�-�N���ڱ����=���fƎ����kmrK�T���iP絵�lg;胳�J۵גJ��]����n�Ie�N�X��s������m��w��;u�7	6N��c�]��֙��l�+f�V��1:{��1��۶p]��s�<��8�r��<.�	���M���7R'��v���$r,�6�`���b��pWd�k�wlu��9��{b���rd�#��b�OC�܇8�=N���k�ܶ��:���ݮ�ב�����x�E�*�8�W��x�Ժ�K]��]��E�r���nTAz7bգ�/`Tڳ�Η����3c��s��{6�j����v�sg�l=�+.쩬��m�{`��r�B�Z궇t�=8N��{ZU4/\���5ͮWV��f���Jx7=�w@Y5΄4v�����?��"��r^6���-w��  ���J���+�gOOWR+�n��G��#�ETI0E*m�������R��4��N�V
I$@�tKI���!'�}���x�&�K�I����S��)H��)6�1�$ n��`��uw^)�o�̬H >;��a@$�fo]�J���0dD�32�z��}9k����8 �s��w7��$��۴Jl��ۻ��)-ߛ
*���!A3U%1�{�w�� 6;w�x}��m�_q�j��~`$]��wi��n��`�v��<M��2����rz�����X�ռ���f�r�����b7�z*I��{h�$LH*IY\�sz�bvo;� 6;w��*�v�]��͌eyVZB��~��ks7�� 6�l‣�d�
"i��߅"On�A�U�-��ۺx�Py{�j�)F�$�BӗF�T�
.�b�,�����k��9�jP9ې{��Ѵ��}=�G����g��6 ���� #c�|�A��fi�6Siz��#���

P��o�6��Ց�ѻ��`H���+2I����u���N���"PX{u�
H\͘ʠ)H��)6�v�z-U��޼Y⻖O�~�"+����q��� -}��5N���'0�L�m�I
��dĩ(ș�!���Ԓs�}���h���(��f�]�(�v�6���ۮI%�k�m&\]��m�����$�R��6J���;;J�]gv��7
k������{u-��*j�Q35SR�$e��݂ 4��1I$��_c��A.�&r��۽�[��8wv��8� I
�US�A�k��/��l��]ϟ+  KM�t� ���d#m�{����S.�- �ҭ�%�UA1	�=�YH��l��%�\�Gz/�ȉ�~~ճx%����(���� ~�$��ى1������;�\���!��I�..}�r�?6#��ͧ�����X{u�E��j��x��!L�$R�4N���>�=&=�t�z*��"I^8�4��Y��wR���0$�$����z���ف$��D�RHn�?�H%��͗�ȭ`������- \���|������:4�����������jݽb�ț���=vմ���8���͵��������������f,k�]��t[�׃��X�l���v�-�x�����p��q�?R���m4I���߽&BI��������#�~��A`�4 ��wi9ڈ�=�k
��)O�E�DĂ� ��������Ղ��G�8��ufV�.c��fw]��T�!��A)#�G�۹��%�Ĝ'Gm�����w` ���w�n������o���4���msI�.��m&Ĭ��'X��9����{�m�v��Ѫ�VSջ���BiN什�7�- �;�z_�D��L�	el�yh����1J��ܼ��C��>�O�ngsv�##�}Q{i�A��hwp�x^�P �Ԉ
"#�W�m���i�KlM��y��4�FJ�P��|��<��2�d���6:�� n�s�dDA�n���T��w�9�lq^��@�w]�@/tK����*����[o[`w�������Q�]9n����޻��H!gn�� Q�=}���3%�ۨ���~M_&�?�X�a�ˏ��ޓ! B�����B�3eߍ�Xw����%�3�]�vbD�1 �%U`	3=�^cw#ku"cw�߭�H�`���{��v�0�@%}�n��]Cj2 D�%�!2+���y$����@�
�i$wF�����	���m2�2c~3��>�'É��bιmwO��;�p�-%�� �"�}����ܪ]�ݻ�ЛuMCc!l��Ah^M��n��8��PkU`�/޻<�J7<NԬ�v}�+u�λ>�Y�ɩ��5]��M^M�N:yM1��N�� �46p�,IǮ����s�J�sm:����FƉ�{lN㎺���{k�ٯnֻ<��,���g�Ώc�[^qZ�ƭ��׮��H��O�����c�K���5v��j��vie{�ω���E�u��]���l��h1\<��Ż"�j3�]��9wI��$�mh�2l�ٞ���au����s;n����!�߈�L�)����T�mŁ�-��?�  ��:auQ6��7^���˻ -���{5d��PT�2���aѷ�����Ef�������%��;َ�H���*Iid��C�w�>Ե��|I��F�`���@.�6�?C ���S�8�Muqu�=�q��cl�##�<ׁ)��MT��Pb&L���޳�����RtJ�B{�ވ����u÷w��((�ܳ*Ը�"/�)���tA�2}1 �%U4�o���|��;{yݗ�9^�L��րJ*�ߚ@ dm㨆���	�u擜�\��84䣙�J\u����Xj��`&x4]��Z�'vvK������$�k���?�����fG�	�6� >��i� �3wy��Ϻ���,]�[dD����R�T�D̒IJ�w�����g�>�s�l�}{��,C��K��-Tm�5�*��`T
�3GUiM�����L�?���s�f>͆��k7/��[���r����S@ ��z����{��Qջ�drv�W�c�Q�YyD񬺒u-��w�i �Iq��U�cs��8S�_g� >.6�}��q�X��Ǎ4�:/�s���2��O�ߺ�9 ���DA�n�]� 6��Q[ϙ�.q��,��1�HEE�L������2S����:�#:������xO�'��{��CA���� !f޶2j:��ۛ�-�� G��$���L:�u��i�g��&l�[�ݗ<gv�sY��<����}�<&O�$$��	3u�K� �oo;���>�����O��odp������fn�ݠG�&"b
��&dlO�Ͱ���bۙ��}������w��",Y��� 3 `�|]ɻN;��x�;�SQ2I%*�D�<��@�w)�4JI���#�L���k�r�=9f��!j��ٺ�#QS��"+lZT֛���ډ�e\^�y�\�;2��$뻊�\zm���� ۻ�v�f�6�*�\��TĊ�)z#��sL�^�E�MF)����Շ�|Ƿq�,$�Xz��#N���ޣ�\t$�շ�v��Ʋ�(H���U����`���i�Z�F�{o4�@/u���D��m� >2;1�ya잿.����wۮ��������q5Dպ/=ƺ�]��ȍt��E�1�<�f���\_~}i�ܪUB.y#��n� ��|� �_c� �6b��w#[�ݾ��� Yۭ���)�UQ�T����s�4�9�vi���o�����on�4�H�%�u�zT^�4i�ǾIW�qD�JBI�m� |���O��,�쾝�S��`�s͑��o�	Ԧ$��aH����.ͣ��~���.�@����|�#��*XI$����$��G��鼇[��Y9AT%5��e�λ�=B�������~qE>��~�O�#����<�om�Hj����yr��9WiC���F��P��$��E�r]�ځ�e!*�2t�� �J�{��h�uZ
'�m��H���lR$�;w���Y��c���;\�Z����n������ۧ���؟M��r��qq�7~������]2�~h�~�w� �"�~>|ow]��0�W��v�ˍV�H�t��Iu1�30
fbj�C����w��7�)��c׿�b�������4 v�sq��
#�x)QѾ�'�$%$��q�֟� v�s�� �\������V$ FE���x��������u!(��2L��Í�s{�۲�l0��3�~� Y��w`$:/��{�ꎡs6��K��n�%.x�S ̘�J�GU�]�`��{~kË!��u����.1ߩ��{��@���myH�5��u�bpm��kDi���<��җ-;lh��O�kP�7$����d&��TQ�fɍ�OH�{�K�.#j�U�o1�ؖ��0��
*�U"U�Eà���u�u��dwd����ې��을�.� ��c�1�=Pݪ�4��<*�b�+e��0qn��v9��۞x�X'L��3c��Br���퍣T:�r:�ϔm���u�1��l9n7]<k����#�cA���gG!�N֬�t��5m�*C��N:�G��xA��Yq�ܻ\����ժ����
i�q�բpv9s���Pq�{t�y�$�n��b�;Z�7�l�-qھ~�$�3�S&E���ԓ�^��-  ��n���[Xn���l.�k�	���v�QKGrD�*���?��^6"r����b�Vjo��+�ٽwi$�\o��I���KWM#�t�*�����	�B��9w��+���N�H�����D2[�}�rOy$3�z���'���J���X�>Q ��g#Ue�H�bp� {ٚ�Y ��n� #"�9%֞~q�����5!"�i33-�7�� �y1�F�軜x�l$��˻	/$p޺t�Hᾚ�������L���*bNq��뫵��X�"�q]=�1��'� �����]�堋�ɔ��,$�{d�BI�΄�	j�7`�^�����ܶ�=sX��$�3�S&E��bʪ�@siqi�������Q%�j>� �E��e�w���~��͜�U�gjh!Ӈ:;E�
�t�z�*F��eʊ��)<��H�A��E{}TH�=�|��6�nޞ�7=�$��i���/'��N�A��LUN�vY �F�u^>���Q�3)D#
bfTn_=QϮ��ϴ��ڢ	;��D��w� Z��H0c�:pw�'�$$$*WӠ��}�̐q���I߉�\P$��� ��K�{�k�`��lί�
	m���*܃��.Z�y�Z��j���^!�\�Q���ę ��tA�"HQh�:�H:�(Q$��y̓j��W�{\��ə�	!��t0j��Fd�&$S�߉�����w�U�V���U}���oĀVH|�3t�3�����6��LʅS&E}uD����0�L�1�a�r���[��'b��[���2����yy�w���>�L^�s/���<q5�GQ��Cj�n(fN{�P�ll��pC/���Ȉn��~�U�����W#�5#�`����e�[��;ޕ�w���h����~7�6�P�����^a�K]j�2�X��7,�V�&)�ME���srzN7�iul��wqТ�=n�{�;S�o��6�lN푑8�@^=�'���${��ծ}�@�B�Oy��wc��|˪��q~��Fw�����/w^�W��:�<�(�8b����/������$� zN���S=�O�a��&�蟼��o�����5V�����[ɽ0�<��3g�����q�su5�?WGwsQ��4�)T�9,�p2Ȳڧ.���w$*�{6�F����Kڸ�r��콑v��|:�o
�!�Y�)�Ǿ|}�s|��/J����sb>���7{c��~�CES=�����y���1�,�H��ɜ�{:<��o��׹���m���̢E�5�1|@�m1��$���-��8}}�!\�-��WtuG���4���q��#_Lђ;׽�z��)]$h��#��=y엷 I��7M_��mJ�a�F���:���j��F��[��)n2ғWAn�G���]>F.�\��m�S3�XKm��1gU���=�q�j�ƾ�Ym@���s���2�I�Ҟsg4�,/�=�>*�V��o�Z�Z��I�ÈLx�?�JY@J-t�=��L~%֨��I1�
�TU���I��LD��80O�ij��5Ypf#i��qZ�+r�P�lZ�*�8�f�ZEK�`�m�ZSLm�-��1-��52̷��W-R�b��TB��ʃ���feQQfd��SD���JT�e�
�b�Ĵ��*���Z2��Yh���9����m�v˸ݰx�<yN�#ٖ���e*�GeG-�6�����C۷�q�'����`�(�(�� ��AJ�eJ����L�f.d�Z�bE�F0P����#q�e���#L���Z[QƫQ˂.\m
,J���ƆaG.9mE�R��h���cs�;�Oc��0	ܫȻ����%�4���9��,�.2㌹Gm-��EA�a�S1�m�+S[i������T�Q�r���)��c1�.J�n%k�������Tˍ�1�C�Z�R�D(P������:�wo9�Fn?���i���~�y��[sYr��
Gu�6H$/�
�<�
h2�������m���Zma.׵��l�u:��*�u���$tf�	yy͂@$/�	��"�3��ʨF
��h�m�������vz���:�8��[g(�K����zkL���E��w�wf�Aݾ�`�	:_8�A�}��컺��=/����pA!��BE%�E����|ud�Q�Ro���}}̓�7Χ��LR����>�CF���fJ�bC=<�	���В	����J�'�L<�~'�w��$�F�uQ��Lʈ�H�ms��a��3�3Ug���MO��U���f]��F���y�5sQ/���nE�zzEк���8:��I4�i�;�j��N����t��pL�`�5�^I�1�B�����͒.���$)bT��mfP�	��}^�Qw�����ܚ�l.�*�6����o.��U�^��D0_A�V����vv��'�ٍ�N�`1��v����s�M�E�v�Lʈ����{x�>$.�j�$�}�GF�ܶ����p��$�6�
>V3ɉ������<"��cg^k��Q�X	�N\�� �{�@�[Q�aE�,\=٬н3F
�D�0�"����$���Q$��<�b]�H���������T̙!A1!���﫧����+��H{=T	8憎'�v���'�țu����������A�T""D� ��РA{}��4�eW\�L�9����r(�e��|wo���w�(g! ��Ea�7$�6s�}ηw$�<�z�g�����˥*�gb�v�X�U&v�q���Ä(}�UK!_68,+ӸG!�3"`��$%!v|�I8䞴�:������&֕����۹űc��ċt�!����a�ŋ�����*��U�\�Z���rp��
���t�s��{-��g���n,o6S��	ݖ�r�+��x�Ok]ø�m�+*Dn��lCpzݑ��Z[��ne�.�dΔܶ�t=v5.y���Ōg�nׅ�`v+�c�Y�f����Kv3S7�s˧cm��ٺ�aK�"s=l��-Z���r���
�2fJ�f%H*�:�*�'.����}����ٙ[�!��H�����숙3JbfU���oĀoy��w!vV���_U}�}���l��ȑ�St{Y�&&O��HHM�O:h�{oz��ބym�1�4	$v�UA=����0�+���i��r�Y�f�f�u�k~$�1�Uc�5kn��_MM�ClX�2&DJ2Hoa�~Q�*9E�b(�@�n����a��1�P;e����A�������Д©i�Mm�[��zŨ-�'��QZ��sOl�����*a@�"G�n��/v�$A�=4u�)�\��έP��B���u��`�mQ]fL�Rĩ?t���׸�8�<4d�����QD���;��{U�n��!�������OCt�?p��m�w���ޜr,��/%п_��nv:}@���m0O��9�|bF���{_��%bM�q����޽ـ�'uP|H.b�Vgo6	����A#U
=�畉��"Qf�s=Sv
�I��u�H6������b����$��l�FQ⤙��ڿQ��y^�6�yu���߉����H$5�O�>��;{Nb���
!\%)@��=����,���ӧP׮�n�Gm[�gr1���~���¦DL&B�jj� �5�U	'�o����s��fM_6A����9PtAe���<߅�#��W2�_�vn��i$����hK��H��#�^S���GM�d̕"TLH)�F���'.��|k���#���]�F�MN�.���8���t���L��F�W2+��d�Yuest������������iEH����QKKГ���H�����"#�"d�@S0�޽|��E�7����4H'6� Oon�f#m�k���� ��UDn��V&O��DHM�y�(��|�*ٶe������M�]�P�;{u�\ޓ8�@��@��	aN��!�<��8�nk'�v��sn�F�[]��<��XΌ�`%3 �(��)�'Ƕ�I n��f��yS��C�W�	uC4��bD�!L��<�'����D�o]Q�$���N�n���s_Boh�6!�� �5D�S
�(�I�n� �G>ux"rrۑ�������ݦ	ڐ�	1!H�
~�yN������@��{i�I#_7W�w ��D٭����c�f�����e�1��S���th�o�y�[:�w^��k��[�h95������=�;�3n��9��໹�ҿ�l2 D4��w7�u�@$�}uQ�D�+=bH�	���^���� �F����q��K��;=���xn�^��6���M� lf�WLvˎ2Q�v.�L�PA�}�yp�>R$#!h�wޣ�N�v�cĂ@:��E�=��܈�����wݭ�|��PA`�Eg:�|US�������$Fwv�����Q{s�w��jVw_�t/��&$I0�lts��	� �yuG���37��a���{w:��$�}uD���3`A��>���LI��fI's���u����8�7{� ��l�	�����S�MfG��㾡VN�T7�� H�׍�	sˑD�}�^5W�q%S���!�p=W>���u��܂�Q��W�����}�3�jL�/`aƙ�UAY�7��g�����糾��N�묉"P���x#�WS��Cm�p��=�����7Fr���ٞ;wl���h䵍��v�m�(pnu;��݊7N:5�mm���y��=���Yo��]�N�n��cpl8<�c��:��;��g��/F��D��nͮ�!���+�E���x{#��mlo����n4#d{�ݿ88�~v�n���ٱ�C�v6{s�B]����{=�7v����Ƭ/�Ch�#\�J���]�\ԛ�\���ߟV�m��/%�s�a��-��@&�uW�P��MY��O�[~���T}��z�̟)��5��D� o<�%�*�;i�	"���'��oz���w���SQ���d�q��AR�DEx��t(�u���|t�;�5�ED^f��������oS��o�F$L$�Ildu��[1����r	w:�$ϻ���j����Eh��3o��B#�0�@�"E}V�&73�V�{s�|][r3W�@�[���}[�Pw*w��\s��X��=T��u�f;V�8+�o:v.��W�)�D���1"��bD����W6�MN;�l�|cs:����Nr�D�B��gS�Qj&L�d��*UX�'ƻcF�3�7��;k�Vu葑u��t�}��x�Y7xz�^-��=:��MNu��W:����!�{}ȴ��)S7w�j�
 �	���~b33���}Yd���7��~ۣ��3'�D�H-�Y}͒LogS$���B�v1����k���I���O�39�|�ƋPA	HS��X�򧕘�,�l|H&73� ���*��X��\����ct�>x�鉔�D�ID��:��컯V�M��jޜ�R2'	u�~$#{5��N���N��3[.�"�_PS�x�"6�csM�(��d�;�e{ZplW��\��0B/3P��L(DL��}V�$��u0Ij븣�b�ġ\7=��$���b�����0f"bAU��y^�+jss�wE�����ۼl�H���$���٢*K���׵ĊQK�d�&R��P�ך� �g��H�ɭU�K�]��u6�jݢ���f2C�Da�ٝ��5^�0�?S��A>�k��m+%����r��f���{:���S�[:���e�uo8�9�͒I��u'��0�O���X���..槍�h���OĒ	��qD�E��f7+��6.;�L��q@�����F�k� �u�ks�ʜ������>$=w��v��/O����ɠ̒���5P���*��I�v%������r�>½	P�Һp_�����4�(�_s�m�i˺�	&�o6V�v;��W�2}6�$�g��	>9�=�1"$��=m�+Ec�]=��d�I��(�M��oă����ek����(�fD��S
l�o+�Hǹ��;"��eۍnʌ�	�u�o;��|)E+��	��d%X�s����H/�%��$�{��	Y���՛�;����xz$�9��t~;n�"q�v�ÿsV�n���ȥp}���G,�������U��z�p�z�&]]�\F͡'�(�
D��O��٬��'k����N��^�'n(�H�}�?��͂�Aڱ;Q&q��v���2=sq^\&c�3��>��=��7\k��9��a9���u����>�����C�o�yU$�u��2A>Y��<���'��v0ٙ�H�y�7:w�L�2Q����m�NK�{<�H��8I'Ď}�߉$Nfs��]�'cFq��A��Jfa$"&I�9�a�L�gS�I\!^�H1�v,����l	��߉Ȕ_	3"DL)�1ƫ3*;��łA���̐}[��?��<b�UN�Up�vad��� .��1*)lH�$̨"BT+^s~$����;�n �eWD�Km�����owro�$�	/��$$ ��I	O���$�HH@�����$�`$�	'�䄄	'��	O�$ I?�$$ I:��$�`$�	'�BB��	O$���$�P$�	'��$ I?�	!I��IO�H@��HH@�rHH@��(+$�k%;�9�ڣ��B
 ���[����E����  @�                           
        ]��x  {�(@銨
�*"�(���RE
�
��
(����@��U �)A"��"�($�UR���   E((  �
  �R�     �  � (P        � t \�� (@ @��Ҟm\Z���:�f���i!��d��p .�R��u�iNms$I�����U+p -�nv:�7,t�HD��S覊P<i}5 *�+�ո 'R�L��MR��Nڜ�%E3a�i��r�)i��R�Z�'-R謮Z��F(��J��7�� |       ��Z�*1�����͝5&���b�#�x �S6�<�*W��=�rW�!Oyܽa�y� {�zr�m�� �x�4��URU*���= ��� ��րP�� }� �����Jx���l��������h�� >�@s}a�h� ���o3�B������@P
;� �C�j�   ��(s|�С�0uv�4QsB��`{�)����>�굣������Gy�;ؗN�ҧ��<=�����;��*U"	I|   ��z|��'���WZc�> �,�����ͽQ� tWOz޵MG� �r���ّ�3�����{��֥UU	-�  �@ 

   �{�T9�K�hy��ng^�G�`� ���8�f��`r+s]Us��p ;Q��c����R��IO�  }���JP�UV b�k8�7XP��I\�+�� ��˳CWwS�;��Ss�����(JJg�  ��  *�   ��;4��9Tu[���}4S�����!T�j���������'\F��è
��x   -*��J�J�����8 ��-����h9�ִH�hu��ͧmI5�� �J�e��kZ�ݖ54��%�kn�Al� |�  5<�Ғ�C@    *�	%*��L� �@Aت�bE(422�����@JJ�M0#	�0	O%)�TD�      I����!���MM��mOI�����̿������?���O��{�h(�f��ǑPz�5���$�}�b?�B@!$���i(&$$��� BI�,��	 ��������������?�����X	"����I ����	?c&RBO����[���������?��m��m6�]��mv۶ڭ��(��m�[m��j���m�m��m��m��m�l�[m��m��E��M��m�m��i����n[m��m��m��E��m�m��E��-�ڭ˶�m�m��m��� �BN!$� !8��� q ! �	'	8�N!HN!$�H@8��$$!8��	8��$�@8�� @�!�Ha � @�@�$ q�@�q�!�$28���H�8�Ya$8�C�0�$�BHq ����`Hq��$2H@!ĒI0 q���L�qC� N$�0�� q���@� e�0$� a$!��$Iq���2�$� q$��N0�q� � d �!&�@�I%! �!�8�@�!�	28�l�8�BS		�'@$�! a��d�8���P q��ā! �	' q !	��ĒJd �N2@8��� 8�I� a �	�	!S' 8��ĒC�����	� , 2����$�9�wwu�l��m��v�U��m�۶ڭ��n�m��{�-?�~[�;�߮��Eu�J#�I���߬m�q=\�Fw~M�ѷz����#�ǼN^��EV'��h�^�o�g�i���0F���;f܀�׶���eC9��*r�{*74+ȤD�s�j�k1͏���.���ɨ���^��,��M��9V3E��c�ƍ64!(���<�kc�5˜-�eU��<�vs��^��\��&�[�7ʰE�NX���W{��z�Ɏ敆^�}3�1�=�}��N>ǈL��Ǝ��ƴT,G�g�{ }:�N�xH3w9IH�#����z3{���5����غ�q�奼�k��f�	�4��Ҧ�.����:������9���:R����f�����R�2���sig+O@��Δ�\�9=g#E0�* ��.t���n��ƍ�ii�i������O*n4�n1�͸��d�Ⱂ�2��(6�Τ�9�aeu'��ޠ�{9!�k���9�h쫗EP�m��d&�jr��gfG�G�U�����Y0f�z�iy�v�#���h}m�5�f�q�g@t��ƒ��{�;��!N�%ɜF�v���I��<��l�:�;wΏ�a�q�1�|&���4�i�=5vD+Ύ.�ܦsl���oIo�w]ųj�w���j�-ۑi8ޖ��{���;���mSzn�v�ŹD�-��ӈ�Z.��M��᝹OW�p��_5=�3�^k7v�LO^�$��(��,�m�]e,a̻9�ȼ��8�������#{
,��xa4���J�ywnt� �^���!�i��c<-�
�7�O��~������Ӵ������f��{���'��W�z��%�+/���1ǨI��ou�I^���Wk�cS���t�d{���:q�� �����H�Oi�L ����t�1W��L�����v�y�"D����]x;��.p��.�	�qE�L�%�����Ǹ`����Y>��pU�:6�z�&EQ����ڍ��-'f�J�;yt���aS�L��v׻��e��f�"�:tx luKAˢ)h�W �V뫎nGΈ.�-9'=����D2���P@.���8�Y��ҧj�D=��W�%�9�� #�����M�N`а��oi�8-�qJήG�+�`��t���nMFdչ�P�ց�C\r�����lU(��iSNIe(՚h,�n.��i.�q��$��y�cAgcc��@���T�Ŀ�axF '<�-;��:gdj����S��E�t�SŐ�״Q���V�e<�v���	��/�t�#�w�
q���6tZ@}}T�w~�Zj�|�2��Zo^{�og]����ɿ��ۯ��;�����q���>q���X�[p6	�4#�nQ)��u���4�{�v��^t�-��ɄI0�h8�S�׵Y�ՃX��ڝ���'*ì�m�s��lw Z���9�����^;���+k�m�ᅼH�;t��wRj�>����bn5q5���,�CHH%:�\ʮ�OYPN���K�kCt>y����ͷ8�t[��Ø����Qɮ�A�7����Ζ~9��p\[L[��!K���҃���.�9B�Ɓա�̼��ҮL)r�d��{��LźC��X��ޤ�>��g<�q��ӌ�G��!���T%[�˛ߥK6���lK�:����]�^.�zq0�SV k��k�7A�ro	zC7:Cn����L��;p�.��{�x�r�mu��S,h):�"�&61�лx�'�M'v�jX���6����\���ᝬ!o�f�<��v����ݠN�@�؉��S�ƀ���@֫��p�&q7y�����؄�]�'vU�ʱws�V�5ۋa�0��rd�۽����ur�.�m�g�꼷����!���y��Ǌ���w#n�l[�a��eo�T�VtK��5��/v������Y$;��ͻ���+b�j��d�DD'�M��9�ۉ� SZ�Т�.-��������6��ߗ��F`�6�)�mtV��L�k��0.9�z\IÃ�k���5�2�gtz-6lZw�O���y�9�Xz��Q8Ꜻ�Ţw+�7j���q��gp�� �(I���q�԰:B�o^'��g�]�m�g?ǌ&L�݈�7���Û�&q;����yWW2eeA�x(�c�$f���ًFu�t�w�ut�\ڣnǬ���T��Q*9o#^��re	��1rB��F�9��.��Ī8��\���r�ч)ꜫ�:�?�Տ�q���M�g着vW��.�c�d��e3�⪪�o9�Wn̹3Lv��6�f6�t����ښ�v�*���g����ɳ�*�FJwu�S��	�-ܫ�f-�O\hU��ꛬ��=�U�n�k����{w5ȈL˰�\�ޙ�H9�NS.KSGGv���v��t�K*�ڡ�c������Q�(Ra��~g�-dx �����0�A�d�]���/�D�=��'Y���n�m�����	�aep���a��dK�H���f�to,�l+5�<n=��W]9�����s��/�f��m\-AT����k��אj
��es��Ð^� ���˯b��u8��e�t�X��\yW���:�<�O_({�kV%e�(��tDڅ�՞[a	�k7�a��lڛ|e{F7���P��u��h@v�5�9����W5��p�;��Ex+�4w��p��t�2:�G#�GY�3��=[�����3�qU���mՊǻ�ϻ�TJ��}�Q�.�`�g�����8i�hy ��#{����=v�Np0]�:b{�2M��άQ ��EnopjoO�����V��8��m3AX��mڍ';�p�,�b���t�SnǱ�u��J�1����w����8�;��~�����*+cn��w�i��קr =���-)� ���_����n���Gno@d�i'�C�0;E]�v둻c�PGMî1�׊���N���!��|lhG��{�w{Q�r`�̝[�K��x�b�.�2w�BQ�{�k�]1ۨ�p�1�זi�5�T5�Ck����FC�ݛP�ic5�w�⮘��Y�[�"�����>q��*I�k�ӱ��s�؎̮ۂ����Y�:*��㻫�����h��-d	�.�#ڷ�"��<Ҙ���V�Gp�qyOa��-l>�T�C������0i�~�W������;�S�g!�y�9V�&f����'H	C8��ܙ�-�1�d�ܻ5�Lk:)͂��wk�7#����*0eI�$ά]�m�ܷa�S��v������N��Wc�!y�B�U�(�q�. ��e��7�á����n��s��!��C�We��wy��83c�7����I���[0ܡ,�o;Pq1�f��͎()�4)���cl-�h�ˏQ z#@�í5u�
CDx�]���C,���Ȧ7���,��NBG7�{����P�[t:�r�a��zAҏ=X�Z�����.%�	g�"�c�wV� ���*���F��3z<����%t�wr	��f��&��\�,[t��,,<雈��R#�:��z;�oI,�񆃤,s��s�K�,��L��y�'�N��w�xc:=<�\�h��*�b��h�� ��'eE8��A &+�+!Ip�L�
�t�Y�k�Lぜ� g]6�+V</sr�sL��v�2�Yaq�j9�s�Q�8N��������z�vv�y�3E�ێ2�f��Ë���CՇ#�N�ݽfK�뽠&�����n�i�[M�K�ے1�zzůf���%�'�`
�c��9��`�GcVJ�	�\&IV>cZ�0�զnJ��.�9gcY�4�b�)sb�@`ͼP�b�x�ܴ��_%D�)j�m빨��.�]��cR˲ �&�#9�(��Օ������m�2(�Q��U����R��#�cQ����,��ƙ/s.�Ҋ0n[Ob=ݭs����b�4�M]��nܘ�G���nС�a}��6H*�fj�志*�ە�Tv+����Č-n����g;������Wp/HK�Ϡ���F�V쳣��ͦnH�q,�s����bfn�;��w�ë�{j�1�B�x]i�4����oh�N�4�$A�R�W
�C�.�	B�;� mJ��9�I�S_�p��N�\�)�V�������H�T���:s�nS�;]��3݌n�=2�	�u�-�|�7u� �DDs�&�d-P��}SɅ�ַ�-�m٦Lhd�=�l�;����3ٖ��B+�1.���v�d7�Zկ ڴnɛ�s�5�	���6��]ۓF�n��x=<+y6��L��Gc}���.��ѡ�Nz�ܻ����3 �-�7�������ش��c����t `�-�*K�<�-ˣJ���%�*�~\E�ިT��$SZ�5���l���4qr���΍��^^z9��ˎ���+k�=X*�aY���G7��Q��%C�+�ӆR�������n�:u�H��c�$6��@X9$�/=�����\q��5�=��I�v�cܽ�A���\so�e.T��,,�&��ruc:��~�gaɫ��bN9&P6Z;4di��S���=$�nK�g�f*�n����oS0�k���>Ņ=�vvSm���ͭ<����#�dz�n�����ҽ��%�4_{q�0E�����̻���ѻ8cڨ}1<�����\n�N���#���*�@_D�~ �GR�}�	��m]���=Ud۠Q#�yM�]��=I�F��%�Pt��^K�R��BdG:�E�9(�aH�̙�{��l�}�C�6^��²�`��ur�#7�XNk�9w;A?�K� @)�d�a����[7���{D��݋��FN��`��F68�;�(�sy�	&�����4����ig'$8�d�
�'w	�E�&q���.����b�UD`�3XY�x@�1e|�^=���p0w;��U>j�8ᤅ�,�:���6�^���@��Z��YF~w:k����i"6��V�P3vi^/�.D�Zxi�ĸ^m(fƝ���;^�ooszyا\I�,L��:!a-Z?r�4�����篊�,���Ryn�l�&K�N'ss���{��0�vu�{p��I��wUQ�Ş𫛮�1�t�1�ǁ�۲�.�v�o�N+
W�ѽ�:(9K8Hh���Uj�C�4jt+�7o$���v�ثpTp 
��E�Kۆ���8m�UK&ni�qNs()2�1��ż���$]��"�a0k{^�7;�)Oʮd�5\��Bh� ���u�g�T�#��n�ē���D����%�3D�v�m��,1׃-͚�Q+e-`�T	�y��UP��7DTݚVu�d�N��I!�G�\�R D�x�ʌ_�wpcP�t�Y4�W%@�"�ܘ��3Vxd�/p���SO��Yw��@�z�|��U�^�ᙻr��/��u�cJ��çT�ʗC���C:��G1�yu.��f��":MY���O:���8�ޘc�y�w���h\��&��n�ݘ{�n����Gr�r�8�O��g���U1��C���w������7Fqɵ��\��X�Om �́�d���T'8�n^3��P�X��_�=_�J�YʶZ��2�- +tq˺Vk�ܸ��&^�ݭf�"�vu��F1�G������Ca�離��m��,;�nsz�L��Rr�s�����u���q~��r�itǻ�c(�������qB ^F��[]���.Rsw�L���pv��z��w# �û:���W-uED��p<t���"eΎ�ڃq�#A�?��=��n fM��é`f��ޙshnv��
v��9��5Lo�*�R^;T��3��^ 6>��x�A�:;�tp�F�"%ȷuÊ�3��ؔ-�\}	I�������ߵ�^�=�z�89�<��j?���]$��ְm�����N�Й��:�Yǹ��6d���-���xl��I���;C9:��|��.ۜt�q�L�2)��rb�ｧ<3A����y�mS�:T�X�<+�!�7��8���x���������n���8�Vno�"İ0��.}&��D��n�=5�FhhNޚJ�&,<*������B����è�r��n45b�-}�o�D�on��n�
�3����$�8C!3y�S�w(ݚ���]�2X�n���%]yϘ飬���x.�]X�
)�|��=`�9���;z��wh �q���Jn��R-�Vm�WO�^'����{�L[���Ni�46�P}ӵ�%��u�"8l�Gq����1�$f�c��N��#���>�k�ݓ7v����L��n<�n�q�I�}^M{o�$�J� W&-�����;L"���̋�C8��F5pn��n
�r���� �=�������)(l���`q����-6W�&o�9���	�U_I�<�ת5,�!�X�F��g9L�nv��1D��"�О�p�rX��Z�h��Λl�в�(�3�=����"Rc	�j��'�҉�vH���y\�/��h���q�����5��9���@�w�F�FFI#s��'&���d�j\�7r�Wd�rs2W0��j3f4�j��)*n9���ܽ[Pl�dD噽��Y�S���7?OϤ|�o�����I?Q�H�H		�	$�H�) 	�A@�P��Y$� Y$���B�� � �XE��!
HI�d"�B�H*@��II �I P, !L��(I$P�$!)���$�))  �I�,���R���
@�Y�)������B�	)$�� � ��H�E!)$!�E��	@�B��
d�Ad	�����S$)�!I$���"�!�@�2)�I R@�(�BE�B
)H�E��X ,E���	) Ad�L��@��R�E$��`� ��,�$��]������9	 $$g��Y�H�� �! ��������h����Q_�_�A#�1G0E���O�N^�'�A��F����f�j�œ��H��D�]��]����E�ϸ��������W�i	�H���'�Kki��ɦ�ٸ��rSp	�0*�{�ch������\�+������B0s�ir��y�{_�x����T˻3e�~�S�O*8��04e�Ȝ���9�Ա�M�>�b�n�d������r�Z��Zdg�Q��̾��XW+8��ő���ۯn�eՓ���o�^"{U����:M��Κ��6�ƕ8��;�v�g���N���{ۤ_�DO��E^~�f��m� ��m��OW��������,Q�|�}�n�H��nOw�ax��21��<-�N�&ng���݋V6�6�~j��*s|��6z�]/r�'�ۯ۽�ٶc${E˯�@���{�x�c3m����e]CQ�,b��Q����w{.�+%	�38{6�%�c�<4� vy�wwu=�i.]E����\6{�G�\��77]b��N��}b�_�ݏӲ����W6���:�]~ ���)gr����q���Vzo{F�������q��Z,���ҡ���o9�K��E�Hݮ2Vl ܺK��ܹ�M�+�2�J��`�;&�'���m�C-������J|�4���6d�ƃ�v��3qcP���"�0��m�m�����۶�m��6�l��V�[�`���P/#;w����~��r7�m�Ӫ@��3��Y�Ul6��1M*bw[���q,_��ɖ龶i���~�kaJ�30�[o-D<�J��m#+�(��̽�z�7��;'�r	3�^)��ӽ`���'d{6_,�x�����Y�5����r���xܤn��'��#ƛ��vK�b!��n����:s��v�-Z���{���{SG�'����'=F��;��I���բ���S��{6B�TC;���Zw�����b[��������{�ya�Zj�����9�����a��E��4�M�vl�W;�}�g���c�=d}���h�]x���HX��7�� p���6?m��[�;��dd�v��}b�43�5��y��NE/{4ڎ�c�Yf�dN7 ӭ�ڹ�s�m���K)���¸�6u�u�=�d>����9K7�jDU#"��u15�d�'��˾�ʇo�"��0�1�on��8��.�U��d�׎t��
��F�G�o��	_�p@ץM��=>�G�u��Z)&»ٵ�9��ĩ�y�U3]'=A�Q���y�I&]�7Y��}���<Y��wH5�~�&�Z筮Å�T9᧡} <�j�hrh�Ka���4�7UϘ�+m�`���r;�N���Wd��.����n�"��4��ͶW�"ۃ8,��C��m6�onm�n�t�M��ݶ�m����WJ��E܈]ߌ���ӗ6�!��V�w��Gh>^F�H��M��hPg����X��^��[�*��E�>݇��垘�$
qTSڣWRݧ���BV��M�~�Z���Oc&�� ��q����Ǿ�ܳ)���C�z܃�Os�S�n�cO�lCZ7m��'bQ�"НIf�#��Q���>�xj��5th~~���8]c�y	w��Ƌ��Ӗ���7.ou�Θ��9���%������
�������iKޡsE�6�q̓)8Y�Y�Ye�sb�ٸG+)�����@)�*��Ƽ�n���/!�)����M����/���yA4�B��(O_=���V6�'�w�	��Ǫ^M�!7�!�@����{��������m����Oߎ�`S���w��ڼ��dD'a��Ř�g2qȦ�6u�s|�>������4o����l@HL�e����
e8���6�ג�y��W7"���삡/�lpY�k��W�Z��p�ݚߖ�ʷ.���LMR���7�F�u��؋��GQV��ե��]ɪ�׷����wW1�M�*a~��M빋��,9ot=����ܷܗ=2�����km��N_�f&!ر6u�ć��gwk˻7��k��{�Ůj��k�M�Z}�zI�O���:{�u�l�w�pme�3�-���6�t�r�m�m�m��t�m���d�kN��c8fKV�{0��웜Ft9���#�@�^e�v���縷܊fWt���1^SOG�ӭ׷�܀Lԅ)z=]qI�_%@��[��O��ŬP&�3�R���=�T�;�����1r�Ī �wB���\��6�Mӥ6^�-y77��61&*��g�=B���of�L�������2�44,�;�)�N�d]�"�VȂ�ŭ=aT��`[�d&v�5x�L�L��.��n?x�,o|ʭ��7v� NP�.����sF�W����{��d=�j�9�97����-���������7L�<Y+H]�]H��{u�C�ת���y6��D��ۜw�%a9DՒ�߽��.�����ݱf�q1T�h/�r�n���<�ۜ������Q�w�)��Q�~\��[�jb�0ֵM�X�{Zk�Ir؁��
WaO=��s%�.���,E��e��\m^L2��C�V�i6��դ�,��3����{6ב�z���P��f�0�2b��U��ڷLK�X�]S9x�cݽ��ʄ=g�'����%��5ڃ�ˣJS8K0`�9��؊H.�T.�;˴�Z+CL��v�wS�(�Ë ��L��� 7r΍��e�F1>�������6ܶ�n�p�m����n�ni�y{���٢�i��&+�o_�ܦ�2+#SV�����up�j�lCx���_�$8q�.�z@s����QH��U)Z��Jt�~�!9V`|<�#�6�c'ٮ�G�6on.>�bפ�'����$���:��(K=�p����-����|��h�wn)�{���g�C���5��3����z��4�㔝�s2�//��*�A�:D��`���EfJ�=��tK�rzP�/àe��lM\l��.ȄS�i��X�EN�5�>���3�j�`7hu�؜������滌��a:�:U�=夎d/Vn�}p�y��g��k�xБ8b�eY�2hSؓ�U�gT�;/8l��#m=�^��C��j�;���l�}x�;���ָ�b^'9g�W�,no.|�C�<��k��9���xd�;���=���k���g���7ע���}��2��Ti�kdeh�^��q(�d��A�����i8����1���n30�UXN��#u�u�@㳧���rN�.�7l�t*������A3��aԕ��=���w�L�O�����m�E�嚦�M���{}���Da�Y~R������r( �q�se:��}4�'w��>�D_���*�?s	��])���k�_�=���aӞ���]�޽�u+p'����v`)���P���dcm���m����m����n�m�i��7���?	n�f��pOۼ�\�{ox�÷��~���n��a�|�h�Ȗ۰�,v�z{�%�a��a�������}}no871�qdl酻P���3�"umb�A��9*6������8+s�Oh��kɏ����۰������ �'r��`���W~�8v�As��I�#�L[�o���&��w�v�ې{A��DT�i�s{7��HU�{}��)�&}��Z��b.�N*´���g���q���(���2�dr0V�J����V�~�~z9�<L]��7���1�{p����k��w���\|}��������i��9��t��V�=�;_��q�F���ѭ�K����� ��] �)�%���p�_薫U�|;;nn˞��͏���7BUe��n�����}���td^��/V���ny�ՑmY�=q���މ�7�Ocx�ãVQᚵ���ǒ�ytxE�廋/�O��6�d�� >v��n�hD��"�����/�-C���*��޾-��g�g���]���5Ne��DP�!a�^DX�l��w*���ۆ���Sʵ����X��1`PTG����[��[��<��/L8������%�f:�������-t�zn�=�r,�٧|��b�>�]`�M8}������/e��hۻos��W�ӕRF�����ٱp�ܲ��-��׋u��z�m��l6�m��m��6��[ݜQ2^nF	�׳j�7DlQ��8JY=�M��.'ۅ�'c�s�.�g��G�f{N�ŜA�*^[eW����LN��n�3�8��R��]ݚ���L{�z�6hˍTQ�40t�E�o��<��})��SX��7���r~O���2�����X��٪y�ܝ�px9����;��^yL^��vl�b����n����u�'�@��Xh��B#{ln�u�,e]�/E=�po-��=�MѦv�dpF�)x���/Os� �
������Y���N-��xi�J�r����������=��l\5���b�{%������{���������]{#�8�g�K{s�l��z$Z5�TD:�Ge�:cM���td\Yx6�խM.]���w�^m]�=ty������F��a��f��tͷaΰ��+�ӳ4s�U[sˮ��.RqK��	����!>]h��/���U^�����H���J�8��{�4��Բ(����GVL$4V[$9XdBb�ݱ�l�qA�x˛���Q�ӘN�I��NC����u{:��2�[3ʿН"{�u�
_�����·}	�Q�r+�^���3��Y���5PT\�unR�������6v���HI����h��=�j��Ѝ��=�«(��Ң�.��(ˇ-��of͞���7횽W���m��m��m��m��m��m��m��{��]X��Fئ^�)��F�T�A���s}8�ڞ�鸵2O�nYhXW�*/���e�18�y�w�*_�����Z��{�H��6 Ԥz���a7��x0����P'�ʎ{/w���u�pC9oC�p-����9p�o���pI�tX�z�:�s���{UL`Z �\�}�
���WÞ�}%���J���i�aܩ`��n�z�����{�{̼Zyq��ܐ���=vnx�O����C7hʈMð�{�D��73��x��z�L�dZ�3F�'⛋�;��[��觖<�������a������<Ҳ�{��� '�y��FRp�>Ko��y9Q"��^��}���{8o���{�P�n�bt���C�
��M~<"]���x$�0n�cr�ȭ�4Ý����©��VA���[����=�.:�k<�/|T4]>�X�%�x��}�df�ǣ6i��V���֚S��"���|��뷧�?5����ں����rxa�۴��=ݞxى���K�_K�,3�#*˧��[���ȸ�!zwp\�M��y����;D��ɇwC�����S��@<�Ɖ�.�+-��\���d8t��������#��4vT��c�֞·�z�N�gd���h��X'������9wD0�T1T��懭��l6�m��M����m�޶�a�����%o����Vn��s��cd�@p�EΛ��R�i�e�R�������AX�k���.j��'6u1}:��zc^��v�������������Q7�શ�<�vuӦ�c��jg����D����t�N<ܓ���L�^9��钶מ��}�Un�5�3�=bۼ�<e�����s)2x��*���»m3Of�'Q����qз+$fԼR3.�_�Ҷ�yG��lAwgj�A/�p�_�y���u��È�h�d�?p!S2w�w��'i�/�zL�!n�D��,����<����:�f�1N�//o��$����������ۉk]�N�;���q�{������=�g^ޒ����T�+�^����w
������V���yg*=��j���s���۱{�E���<��w��YV��֏D=����t)����{�.*ƃ_�n�s�[������"0��"���,dAw��`�9-��Y���$��j4<k;����3�Ҫ�AC5NN��9�����0Iڳ+V0QB�F���j�=B��?8�*j.rc!-	�^z=��W�Ѽo�{�{rF�� �����3ȧ��P��L�:j^��h5`�a��2��3{�m��N�l���6�
��*��JF�$�sW�z��nҷa�
�״!���O%{y�9[*����}|��zf��C�0����O�o���ǔ�����U�H�o��������&�����28y8�1r�rvUy4���q5gi�0k�j��\l���ڽH�1)���}��8y>Y����_{�ȍSn�nix������F��ږ�jz�)2�
��HZ;B�=��ܻ3�����>W�QL>�s:4РȦk��~>΋no
绗�
?QϦ�:T��E���OR���FO+�5+��-f�֔�P{��#��G��%0�r����Qu[ި3r��f^Y�V�	
�X��ti�NuĝF1��E�ANO"MV�E�$���>Si׋ʊ�PF���
�x��x�3�v k�V\���Y�n�m=�wB���^����/�)��l$�"Ru��f�7$Lu�ع;�;Iދ���o��x	}G��O3�Z]1�>�j?>Z�A7�s{fُ�2��*�?[��O��������n[���y���ՎL~.E���!��MF�Z�2�#f�ɏ9��J�[�w]���q��<��1n���W��t^+���d�A��5��ͶR��q��g
��"�.,O5��z�����޻�8�Sb�`�̳����"�2��ܔ�����x��m��.Ҏ����i��޷���qr�=��^
{՛�Ռ�g7 �zN֐DZ)�9q�'�;�o��M�y���w��RB	"��w�1��X����_��ah��)�F�Ć�;gu���;n<,���-�d�xȝO*n٭ ��0;^��vF�D���ך�u����t�������y�v�5��O\��=z�uݮܙ�Zz*!�c�On�Ѹ
uy��=<�>{:�͞E/Nn��y�oF��=@�檍n"nΦ�;T
;u4�ٸV����<x\��Yrt�gl��ڥ�Ħ�,�f�W�0�ɮ����ݝ�:���������ϝ���ˍ:�������C��w[1:z���N�o#�s�v�ꊹ%2��d'cv�[�����s��ٶ���7 ��1n��u�klgQ�Fl*��(�(�R����\�DN÷���<chb$gl�����;Yr��n`ݎ����6��Wp�Y#��'m��E��(b=#�d�'+����c��Trle�6_@Z�y��;s�����/X[�ms��m��5֣m�k���Zq�V�gb;���/bu<�un�)r���]�kY�9湮��㞘\v��Ѹ{�ۭ�p�Wu�����z�K��7f��=��]���n��r=Hu�`�<1�c��[��u�GA5��ۮ�ೋvv�����Vw\mU�2�j���ӵ�&|^�7�Wo
�6+q���we/��	�=:�n�v���6��� y6��Cd�v��p��O{.-x��z�o:Rc޻q��*�v�&٣ƅ藃pk�;��;�ǚ��F��vk�O�p�:	�n�^w;ES����.nL�ۂ[^��]���&paS��hk{�6�����Exu�Q禖���B��Hus��hZ�c.$�"8�����&�u�m����Ƃ��[Z�X���S'Y͑{:��m�uG]U�Н���Ƹz��Ξ{&Ri��j2݋��x�ܚN�/[֮s��]6�km�vfųXy��&4F֟m#֤���;]n��6��FD���Nyn^p{\v�q
��v��務.;r��9�u�z�.޴ps����]���x���nӛ���|���s��h)��h��ʻmuu�Ե<ڎ^6w]��<���͹ܵ��s�m�e;K�{=�$��v
����GnR�=�:^�/n6{��5��k���$\�����g�=���r�s�pL\W���t�%u���5��Ț�*s����,.�ݳ�=v6��\�GL9ƎH��ݝq�n�m��W����8N����ն�9�Ys��wStU۱q����n�Sܼ4n�,:�ϕ�׀���a_8s��5�>�Ϻ��f�rx�B��Zj���r��+hXθ7kT�k��N��вy�m�p��m��
lu�������C�8w\n۝�y�]Ť�ͺwJy�B\��6'Ga����tYFE�8��p���v����
4�Զ<*����޺���ۗ��n�v�Hk�|e�qB���Q�z�׆�8�۞�j���z�ĕ�W8�<�g�����\n{2��(⭹y��k�9͛�N�շg�Yv��c�KۜV�\��Bt�eګ���ۄ��κ�/�����Kp�=u���&6�e���=n3�rcݮ���p��6z^]Wfm����e���u�n,�;^��]����y�]��ݮ޸z�r�]�h�v.��8�k�F޷��9�v��s�ny%ϡ:�.n�%R�]��z�e�O��9݇y�v�n8�n�]��]��a�F��P#�Ǣe�
Ŗ&������1�+oE>���5^!/H�c�k�:̓�vH�Ɂ�c����= 6��3m;���v˜S�x���xy:�We�b�u�pu��j�zn6�s�n� �ruƶwR�W3�nq��C�ٵoVa�+����E^�v^8:�*wT�-�i۳�я-��v��'c�\�r��dTÇq�����0z���6ѫn�wV/&:�� <]gُa{Vz�H����j_Yy_g�1l֓��<�Wb��ЏA�WW����7]���h�vӆyxz�k���I��LVp����'��ɲ�vfʯK�{m�����3�k�H����؈v덕}Oc���sF1�s��6z��t�3�Ku.��{0�[�s�G0x�9�A�O<i69���U��t=ٌ��'���oe���n�b+(s��D��m�2��n]n9*Nd�!��]��#n��uθ,�{F���c��;��'�K��.�:�{ű�Z|�l�%D�=^�n��=vy�v}���=ф�*�ς���6wu�=��Q� $�/\]�&j�)�y�ӵA w&�+�c��>:�<���Cq�q�歮�v��v�\�a[�J8��1kcN/g׵Ƨ�<�%�V�W�� �>�uvg�����M��F���W��Lۚ�З���g�v��L�u�씜�y����뎺x,��k@u�y�vwg��֬3��٪σͬ������8Ն��%�q�k�qqb5� �۬^��A�]�����I�[q����:�,��=��/>����^�.�;���{����v|�i,d�mcQ�y7��$���^���	�[�۳��R�kOd�ݹ���n���v 8��d�b5�7�������Gp���΢{v �۠�v��i8^�����J�fW����).�	�P����:����vjS�n%޷V�d��s %|������ù4��'(r���.�K�q���m����۞���-<w8N{�Y�Gn����^p�E����su���On�g*�����]f�N`���2�. ����s����w�t���k�!�㕳s�nƑmnr1m�ɸ�z����mp��]�a-���Zcz}�H�z���[cˆ�.��N���I\�\��N��B�ʯ�n����6�kf��y�㓖ѻ��mg������m7Yo[غ�N����Ä��s��Gg�cn{oL�+���m�on����_:��E�%�C�M��/j�V�V�����s�xz�7�Y�]�<3�\���Yݝb1��(tq�����vE;\�[].1��q��lnb�wNC��9����v�g���eɳ�(�m��qk��f�sȲs��!�-��a]m�Q!�vv�޽Pn��H��r���p�ˬm���n^2����T�Պywm����=��N�j��y�I�w�c�N�ǉh��2k�܉�nf�v.]�QN����k�,�G��{FK]����y�rV&���<�wY����l���f�Ё�%;7PU��v�g��n.�Nq�ݩr��$���<�\8���d���=���^˨yc���ev�Nn��ɝ�6����^L%cy�1��Gng�
�3<z]��Sp/rj�v-�c�:����[a��]wO����n��n��64�;�F�=q��5�˻;���Z�Z��g��z}H���0�/;�Q���,��݄�p<]lv�nZ�i�;'��dS���Ů�/g�m��:c��s'`77W�����^΋:���P����ku{mOPu�9�:ְBn��l�t���L	a���'�\�t!�pmƴp�v�<�Z���0� ��ֵظ���ti��m*V�n͹��������J�}[y�D�-y����/�ϭ�;o	��eq�<�p�k���3Qi�5�G<�صt���V�b�۵<��{ {<D��Ջi��ә�ڏv{ް�ʵ{g�y1kS�z��wL��_VkN�K���`�p�uΝ�c���RY�N��\�Ų�=�Żf6�[[K��p��Ή'�;��|�wV���x����q��N�Ҝ<���%��n�^W,%��`R�����źH�M�v�n@|��]�U�Ѻ���u����v�s��:�9��[Ӷ�DcN�ܘ��8)7=�ݶ@*���9�ۭ��uA\;u�XW��ƲU�후�^qn�7TpS�ʉ��m��]uϩE�\="��r�����;k��q���N�-��/Wn.��<���#�n[��1ڋ^{Y;c�m�D4;�O2�@�J���3�.���Nv�[W�Zo9�n�h*]" 6ְ�_n���8Ktm�z鲦�Z�q�x�/O\s(ێ�6f��LvQ��v�����زe���X%����&݅�n�1�k"[��¼�n&k�D=���[���=�n1�Х�c�(�z彶��.s�k�q�y���p�eg5��<�r�pgf�ݎt���u����6��y�m��$�aG�U�a��6+�8nN�ckJm3ʔ�[Om��7=K5�2mfn2��������kD9��"q��NCa�mpsv�q4�;.��{]����'.��I����� &��v��6GFK��m2�&�q��6������)�.�K�nz�z�`]�Gtp�����hv��9��k�K.��؄ۍzۮ��&���<s�t].KE�T��=��8^(�ݝ4+���]��뎽��q�\Qv�WE\�q�TݧO[�m8饽.�c��;s����:e9�^s���Z�b���.�%��WM�����֫���ث·��tGn��z�v�Xc�Y87k����N���u��㔺Ɩ�v�q�#ֹй��^.�']7����ֆ�q`����'�c� Nɮ�x+�ێ)��+��k;ޮ�qmd�s���f7PY�;W�[��岷G���Cim�<H�v�n�V����vR�%(j��j*����5�rjg��j�B#��bЖ;puq��}�[x�j;=�J�P��Nzy����v:x�n-�(U���v���Ԗ�9��uƎ�A�Nf�cK9ӈ��f�F�n��G]�2����4/���{tۇv�7:��6��Im��r��v�]ŷ%lv$�oI��^�p[�v[��p�l��UkK7��HĦ��b�O��:Ū�i�yVF�YYS�)�$�Rd�x�K��E�W��{�~�?�.DQ�L��By��3�9/�Y�E��O#$��Ă�/p��M��}�{�y�fAE�T�"�TR{���k�yU?��U�DT�_�K��y�{;~��~��J$�TR�̛�I	h�	gs��HI^U�hKGa�|k�﷽O'�yz�������K���
;~��xхzb��*:��	'��3!�yU�~��������5=�&��$��B�UW:9~o3�Sǜ�C�Cģu��L��:+u�&��Ĉ:��cU"�d�{{�WB�����󞞮f�&z�̞<���y�SH�O)�ln,ܦ�F��XL���}��~��g4_����#�2B���ﷅ�~עj���x�|����u�f٣"�{Ft�F��iKESƠ�`��*//�$��P�=ϒ�1�Q�������i�����g=Є��www��ۯ�O��*��	(�c�f-K��p�
�ĺ���&��"u.�b�޺9��'��<ؽ�:%(�)���)ŝ�Ӡ��	^ٹɳ���1���<;��GZy޽��X�BT������j��v�ku����y���vݸ���L��Q�xu�%���K��96�G]9	.�	{t͕�ۇxs�)9ݎc��C�x��</�D�H��+��}��i,*{o&e/s�nh54��e8:�b�A���?���$��ñwl��7<�b�Hs<[d�e�����u��ӭ���nq��a��nݝT��v%�]7�8��򋳊�{q烠��[n�.�1�s��Y�ȥ�{ylg�.�Nm��V⃮��nk=8�64p]��϶�t%���o�>K>ǞN���^�V����P��;�n�<�l�6�.vvR Z�ŵ�X����3��v ��9��5�N�a�����|�]=�De5��ӂ|���x)�Y�I�]]�9l�%ۇW�:{[���n��]w��vσ�Ѷ<'�κ�ɗ���q��3��pPf,��c�
Q�N���&0�7��/j�'c����ۄr�����5�>#�ٰs�OU&����5�Vv�Fws�ǔ�C�3����Ź����A�W�r�[��ݎb�hw�ωb)�;����7�n�8�̺���k�"Q���X7ZɑJ��鷄|kӽ��숩����x������vs[���o����t���c�{:�kr�	lu��ԋ��瘹��v�Z�q��[8n:��,K ;�3vL�n�S� �g�]=q�h�o)����'q��qM�[ga��b���=�^�O��V���I�궝�i���ꮝ���r�v�x���ܖ��vv��j������_I��S��gO%Ո�nb/���"�i���Q���h�����9ɹ�9�_jq��Y�s����{���m������yӵ.%Ӳ-��Y1����m���͜�.g�6�͇�#mSN��3S�du�i�u�ƵN�ɩs/D����j�3�Z�'W21�mU�gr����f�ۨ�:G,B��ٵ�F̘è�v��6e��Ѭ��[��'(�vh�2�3i6�w.���D�Ӑ���N��`�fUQ0Io���o`����� �����v����[���E$�ا�v��ȧ2`B�>Q$��[�T���!����O{�F"
�H8�س	�hM�⴨��)F����ؗ�����jԎ�C[����� ���/G�8Q5���"�ˉ�׸��H$�*�.�H={�W(�0۞V��
�,�����,���G򷼒)[{ooi*	#�(I��K�{2M��N���s����q��Z��?z�r��V�H]���F����D4ttt���H�.�K� o��גA$yݹ��qUU�z*V��U��ۏ��x�#!��l���ܝ��]��]�Q�'s�9��;�����]�u�A����Cw�(�H<r*�+�<�wx�]��*�mT������WQ����r�h�nZ�<�&UwW{�x$��\T9��8��+�����{��s�3�ŀF�-{��/�S�轼wQ��L=E�<n�I}�k��]
����=�_�k�6Na$��M$M'��x"�R�I�\�U��Ƃ�5�Z�
�	Zz����  	^w;��I���]�w��V$J=���  ������E���뎫e����Z	�s�̑�j�W�6E
I$���f$�H'S�Of'�g�ܚ;����8 �7�Ha#J8v{��I�7~��΍�a�=�4q0!�癈���u՛ĭ���Tl	���|��٧P�d�m`��cjp�\/�sb|<���Q�T�Ed�ߘ��Q�ԕZf�SۡT�H�z��ZP�!�u����l���M�;UBh�Ku����5<
0��dH�V�-��'
���.���"�$�	!���bIDD8�qv�H�9�����.�G�uݞ�~�0	˩`;�N��b�����$�z��I$�1Ҷpb8���sݛ;����[��:���=����-�>3��o7�@��?OƗ�קm�[|���^s��'8� ~;3oU�QYXڵ:��D�D�����Ԑ]�(�]y�HPT�� ݡ��42�{/����泯�@I��}M��shNGb�4j���J���{���V��Z++Mkx=�vg@��U~�^����GDHk[�����9#�X$�-�� ��rkn�[�Q\���6�/7GnuΒ���I�c=�9�������� �q[%VB^�m���!Y��;�5�wp�<_zb� E�<O	�{����7�F+����%.���j���T�DD����̡B�	{�9Jv�s7��;ֺ�	 ��5��R�w�+�ܒ�w��)��Z�{vs�3Μ��a'&���t` \ߪ�@�%=�O�ow��eUi-%��o���PIΡ4^�s��'iIl�|�����M+Ν��I�7�&ג �Α4�(���"b�-΅m)��sU��^��m�Y��zl~3�嫟f�G%R�*�h�E����U���G�����{�M!s=	 �*�/֗���8�2f�� ��t+tG�o;w��"!�+�Ŵ�'r.�K�d�hM �K�s����WI�ʄ�Aوu��n-�{m���T[qt�N�����y6�v��%��,��\\^��h��5� �{WI8�A�$�ks��bS��=S~�]S�7����X�4�o<�fi8 wؑE(RUՀ���,�[�{e�0յ*3=� ��UrݴE���c��ݦ����|����a�p;�RRU2�l!(U$H�sw��	<!�D��]qd�H<�A$8�;Ǳ~����8:��5��7�t���m�߻�X%W��H�RI$����y$-^�v^ʫv:v+��'/dM
���	�XN�Ғ�[�[�ۙI$��>�R� Hf��^1�Bk�$���x1�q���=���dwE��$j��@�gU<���I��-�Փ�v���a;�z9:�ș�rz����c�;u����F�\�W{��ާW4<�AN���5xq�7���w�{W;ip��x�t��Kx�X�����.�v6/]��q`T��׈{c6�6���ӷ=I�-[�ltݏg��ml�u��F��0��s\����\�^��Ӟb욎��ϭ�H��F�Ip\������	';�+{f�r�;V�ݣ�;	��3u6c���G&�\�e�z؞nՇ��љ�<ի+#�nW���@���YLV/X�;Gc��݌:����׭�%��}�)U�w�{��������W�����(��j�s�V]u	�nH��]������U��YZkZ@�g\�J���s6[�C���B�ۻ'Alv8�Z+�*���{L��X���gm�I�kR�Y�	�s��� ��sd��WU5�i��*�0N�KƷ�w{Kc ;=�̽(U���d(��eF��K�=��o�XI_u���"Pq���"FgH�w)��jV<�N�b�{ז�y�oU�PuUt6��А/��u�Κ��1ݛ�i,���N$���Ɂ	"ߞ&M�t��W��3qj�AA�iq�Qm�ޓk��zޝ=����9�y��e����":bBQ�S3�ڼ�΄c��v$�H�牓�^	m3s��g���l`;���h1���8�Tv����X���;m��&����a�fk�˲ɐL��ݼ��d�h�"�@4� 56�L������8�I�v�Qr]��[�ǣ�K ��}�|�$��g�&�D�U���D�$7�/^$�&E"LL�*"�=��ZH���(RIQfu��6F�K���X�?$�@;�]h`{�T��y�l����W/�A]�9Ԅ���v*גI"�hM�H.��9b+�hT�j��Q<��4*��,������W���2�ۼ�'1�;R2l���y7i$�x�M$J]��3س�����Ⱦ�m=�!F��ˠ������Lr%[��=z�k�Ўu�H������PuUvy����"Gc�T��<������3y�z�f��˫�Y�'��*�;�#}vT���NN��&����#폱Ä�pOs�� ��K�t�^~\�T��,��j�_�DH�0�Q>5hV�
��&���b%�鑹$��'���m���p�3�,��o&��|M��QK^�bA-��~|�Q�Q~y����_y���
����])y_X�!;B�9�x$/6D�D��ߘ؋�M�.}12�( �$�[���1�R^I���^�����u�\�I8O��_M��jƖt� x/��?ğȺ 7{�J(��m$p$u�ߪ�[�,�qW����H�I����1B�	y.�ٿ_Lå��N������D����f�أ�Um�4{x���Hu�\�yc�-���%�p��ЊV��׻�M�
��I&�wgH$��͛���f>:zZ�;C�"w��=o!g�P[��|$!�FD���!]=ʲM�+}5�a��H��%{5���H�仳f����6̮�$ë�Z%��)O�L��m���LԖ�>��p�$�xcڻֶS�K_��:%�J�z��{%%�6or#��20L)��!D���!�u�G:����	Vm��ĒK�^lݪ���mP�}�z�za�F�N�Y3Z&�DW�D+u4Oq�
��Ӱ��l^����Rd����]����]��E�o�&�}�Rr{2˙�D�JA�9��8I�N^�:��g8�]v����W��vfy"RZ�f��&�ݚ��_�gI���c��D�N�%j�F�4�Sɾ'����x\�s�5f���T����J���s����e��&J��+����#� �:�f���=�Bi(��w/f﯎R�긚z���)�{|�Z\=�t"��-u��Z��ϩlDeqH�]e���o��$�	/.�ٻ	�nP��D��fS�O��0��g�[�/UBsuUti��������$,�S}ق�:����I"{�˭��n��3׬���Tw��X\�3��V�q]��q~I$k_M_�%{BI��	���^�n�d*�蒒�nh����0L)��ED��x!��*��7��ө�%�/U@�Ҿ���H��^H�o;�Y�ݳ5��%B��ٰ��̊fPۻ�]�bL�ʩ���_m�뤙�8�w>��z.����m�S���v�ʔ�+*�����,����M�M��ۯ�x��O(u!�"��g�-�ؖ^���g�����^�Hn�&�vgk��B��qٷf巐6���9��#��4.��:��Zs;��<�j���x�u���"���x�]��۝��3;�{9����vn���%l<=%U�0cn��&�9Þ�k���{��K�����F��lrFRg@*F1�����>ӡy⨁�uFu������l%�9��"��.]Ѣk�<O7 j�7N�����²QIk�w�Y�b�r��$���y��m
�:H����<�ֹ�h�����<@<�P��� 5S�� ă�f���wV��@�9A$�]���Ey mLZB��^M�H��($�L�77�"�
�"R\�wd�H�t���
�Ps���IQ��M؈^Nw�M��<$ cЌ�h�0�46(50'q�Gx$���`RA%䗻9���Iy$\�eԵm�h�^c����}�G����5�k���ZkHזּ���}\r��lk��Ȓj���D���y��RI.w�E�s]��&�X�Z��qM]�׫���BsQNJ�R%�I�en�+duEm,�]�Z갸���Hoe
�"\Df�;�b%$��{7iY�݄9y['�(I4�[��`Īh�ACBb�� ���}��ZHn�'
٘h��hic�{����������f��z�Aۣ��6��BBdYM�mMU:0b�}�ag��V��ۯﲻ���Y�U�x$�Hkm�g�A$���߭�vo��Ow%ʹ9�ߤ���]f��5_v`ĆDBE�w�PH���B4(D��n4N��A^syd�Io^���LDɓR�n����ͺ"�I$�}��4�I��I��~x��n8�蚫�G���bX�/l9%DB2$M�H�n_��D�Α����A��;Ry�'BKr��`Iy%������ݪ^K����MzU4јG=Z���0�$��d[]�;3������.њn��u��E~w���n���I-4��gZ�� ��sY� ���(����#(.���'H%��o֖��n	*}("�|p�]!�I.���g�9���$�Z�f� �H�u	��q7>�at�~�^������ԡG��H��ud�D�D�I�(x ?�D�s��~��E��.0��:����M�3����s#i|0�$/���i��h�n���l	�Og�Gg����x�x\~�
+��f�%��.��-i�k]�/wf�"�a��V<v?Wg��C7�({�hSz쳬bc~�1{lS�Ὕ���Kh�+�i#�����oFn��٩��	.X�`��N�l��+�5Q.�� �Q8gbڇY�R��Ա1�Z�9q�\	�m�:1)O���c �8���:����{�xi��]������5k����y��`�矎�O>�Uۻ�ӁXz�N���~>��;|���Z&
WnZ�=�Ol��gO{�Q�Ļ$��Ӓ7���n�#HdʧS6�Bv3%��r���p��E�W!�k����qze<�,��,�A���=옭� �!�X�:�w��MO�Z���Lؼ55:��ޘv��5��z��㞖r�!<����G]}��SsA;��y<-�~4a���h��W��zf��:��|8�Ӻ�^{�8ļ�Ӱ�Y�gQSY����.���ə�$Ғe�R]�~t�g����<��qe��ك"�/'�d�K^�7�5����I�nz��ٍ]=���4�&t������s�n__�qe�� Ӛ�c��N�^�վ�}.�Wl��~p*[,)�h�S�*�J�uq�f �uv-�b�:INpY�{YB�x\���%���yr�:��K}S���ͻʝ1l��׷ٻɂio�`Q�7dM�l_�z/"�r܆J�'���<��g�H���:�O=[��Η��z��}�o����3�W�L���
/b�����c"��^a�����I�)VEB�fO2�<����￿���ݞ��W�ǟ�#>1 ��9�闔R�D��b�.��!�ngMi�ҏmD�alA**�DP��Ǆ>o^��d�bbyyF.M�{���K`�fqc0��{��"��ӭ�K!���G��*��8{5t�g���=g�B(a�{�k)ߵ˓����x������mm��
1vZSQ��](�ޡ�=�	�<.gbʁ'2�/n����\���CY�E�������D�0�I�h�����z1H���`�(����ȼ����r<�,�ڗ�^�-/��Wn��奶5� F!���6�i�*A�����ag���EOmɔYjW�W�Qa垑�)�8ad�
5\�{��@��RG��D͊{6�<���%L�\��a�d�j�y�=S�G�{Ǳ9�2oK���N	�P��j�<����&C��~a�t�y�Etmd���{Q��&WQ=-x�s8�I&>�G�f�X"� =�D��! �Y ��(�$ę*��w��_] �+'�D�gMpI$KΑ4iL�����~{Gm���\��㧗�U�k�>��=�+ԂI���x1Cf�(�?tQٷ�D@R��I$��P�h$��v�w1yk6u9�i��V��DV�*�ŪsX��V�q���U�n�͊ƣx��ƭiQk%��>��0����f�s�w]��j ؽ���� �Lv���]���J����B��U�E��k��Gq$����Z֟�!�X�~��h�v"�g�&��^_>����P!�9��gϺxZ���n*}("�|~��BM$No|�%ꈁ�3���3Fp�����9�I�.��5䗒K���n�HL�F�����P��Y'�ٝ�v��&]��HU\���%��}�fI$O�n�8i�G~\7v���j6k�-��.2XOEߞ@���P�[pڻeY¥����XTTT-Fb÷����(ꊽƫۗrH7tm� x���{�r���m�uD9]f��k��ك�_DA|���@����wH��"��w���[���s�Z/�:��}�g�����IKp��|��UU�5�Q���)�y��]J��+%�<���!G-�y�B��*�_DM��x1/$J_}�7a �st����h��	�>��$�����ĆY?Ib���Ut6��A�|�w�O+/lC�D��o$}WB�!���0$�D�w&��ϟ$ț�s|���n�x���k���O�����9�p}��h �N�I����{�ku�t%��_{����K�	�{u��^�(����p����:�O%0���ߵt���.h0�>n��	$�;P�Cgm������3Ϸ�����LzD;�&��g��H���(}q�oe�	@K:�ۼI$�p�b���	ϤI8�>����S�|�˞q��S��d|#Jn���w��݂j��\\��=��UPڪ�m��lg�P>z��]�=���y��Rwv>w=�!#�j�L��+f�Dq!�������[�݋Ag��7E��O�9��mx�v�78�㜵�F3�����6�F�܏n���;�k%�R��6�m�qsk]�5-��^!x(�������N�e�Y��<���u��kT>{]\O
u�ݩkv��/p] m3�ݹ���h�dŴ�.�k����
]�A��Ƚ5d[����=��\�\�TA\�j��ٻFםs�I�n/R*v�^3��5�A%U�%��l�X�����}�E�����y��-��ü�t#�LD���&�����ϫ�
��G�v�Kg�ɭ}"P�}�Z7]���wUmd2#�L��.3�]�ć��K����H���&�p"-�s���~�׸�.c��G���h�֮���X���9@&~g쭋??���Y5o:3D$I����c���U�Dg�-twKL��{36��w�K3�(}j��I�~�^�H���w�򊩂������'+�m-Y�8y�����H_g�YK  {9�م�tT|��mUVM�H���'��BU#�����R�S�V�SPI|&����{��uϑ@*b�#i���k���k����\۶���v��.���J)HL5��7﷭���i$�|�ݹ�b�y������͋�ġ��J�i���(�u�7F}?����w��;'�vMp���LNm��S0K-�8�%a�n�L�LQ���L��]�<��C�z=�G ��yqҩ�[f�	�
�����	�I w:��I8�G���q%�ڮd��c�?FNE?C>�vѺ�g����G	�w��{�HuE�Kr���coR��t��W8��w�oN�m�|ؤr�D��JN�>�,UV�a�i���$��K;��N�;�kDY��Rs�e\�rs�\��6Z�.!-��Q�}��ļ�	�ѿ8��=HT[��y/�-�lM�K�ﻞf"��[��ˬ�P�i��~}����7�&�dfi���vXy�Ga�Sv6��=X�#.-�%�;��z�����\�i,߾��H$�Hl_��D)�D'����`��B($��/��yf�A�BJ�"T(��>���Ӊ+�E�4�;-F�r6R	 �}��3BD�'���f=$Υ��:�%�Eʍ�<��R
9h��`Z����ޤS�<s��.��/���o��l'4n�vT�07n���P�=����N��D��y�g3뛾��_�M3w��N\�׻�%.����_~��^��8�m�~�|=]5| �y�.Q�"9����RE��zl�+�s�>	h$�B�`_<�����'W����\���|�c�1ٿrkH ���7b6��d/��/����I(�o3ؐ��O���RB��]�=�u+�  ���F�}��Y����V��K��7�� ��glX�I{�C�F{��wO۟P�~�u]��5��Շ8㮒ڷ�]L���ym��^�7�Z�K����k������浯bI/%�;n~�>�I!��_|��eܷ	�ݙ����^_F�������H��D�����ꑲ�=uy	b��c�<'�}�D�K��|[�ҍ�+Wy-+��ܨ��*P�P��U�����3�bg{Vh �"����g��}θI�~���Ā_�T�;$���B8ʄ ��'B�����n��tFB�I���u�@���L� >���&%{/l���sV�-��y�����)VĂuC�v�lH����N�b��YS��9��;�1P�ۚ��N-�d����g����ۚK@��]^v��ҽ]#N�>z���	}������ʬ�{v:2f�EߒI/����q����r�FQ�1�b���Wu�fq^fR�q�����A,�t������2P�Ee��-=�/���a*�<([�sg�r(zFB0ȏw_�wtB�������
c^ŋ�D�'� �(P�~�qzL��@���kpb&$۝�ݩY�\�W��N�E�(!��ܳ�Fi�F<֖���S6�,�23n�Q>7~_t(uA0�s��{�H��mm�����$N�r"��/����6-���&P�P��f��_��5C]�1(k�������<�I{�����H.����7#UQ����)t�@s\���8㶴{y�7�}���6$�,�����W�b>.dE%	t���{��	$��رiȁQ�͘}@ߑ��D��|��~;����x���aD�
{9��;���A�Wz�Ob]"�g�^���}���{Ogmf?$��r�Tj؈��\4X浱mS|�-���c�z����pc�{P�V�ݞ苅���^�/H����\6�â;J�l����*���s�\�ݼs<9����<a�:��淝��YݺS��b�t:9&��:�W���{B����iׅ9���n��ݲTp��ص֋ũ:��= =p�꭮f�Y�N|;��4=]����q��A�Y��=vD&����wkSl���n�m���e��Q��J��^��//����g��m
�A'�����h��^q�8�H���g���F��(}6$���w��N�?j/���a*�>�RS�n,���*w����ፑ�����y��I'����^H�յ��3/훾�!�/�CQ!F!-6���Z���>>�v��o�럾�=�b"�G�����b)$�}�}7/���a	A%�q�ܰ����}i�9�S��$�]w��n���DGGձfR��݈k�}�?�v\lU��Y�s0b�=�f���>u�JBa��6}���6�ʲ�E���^��͸�X��U	������K��ٱ~��"D%�uB($�|��6��!�E�!���J���'�#[�=��.��n66��97�[�aT�7Ku��tq�Z��y��u�?9 ���w��\�C���L��6і�8��oB�<�q}�q�ŋBN���
I���Pjl-�NŉI.���_�T�ɪ�{[�?nn�95m.7�	��X�%�5�ۼW}~��f���NQ���(~<Ϟ��c d�=xs�R؎Sb�w9�
L���[�@c��95���ǽ�6���������c�]@aA��	D�gܒ����Ќȡ��*�(��t��)��6'���D�1��q��*:b�:�[Q�)Qq	og�����n�=}��<�9��7$Փ�vs(�5� \��J�Zw+�E-�����]�v(���n�	p���ee@�5�}�o3.s�M�'��֑��9�e�1�����͓�7>�j��5r�1U�b��k&"�G���JT�<5�P#��5z@R3ӊ����}s�QɁs���ЎI�N��+ �	 >o����ZvVx�A�Ww}w��.};�����tq�e��w��� ���r�����C|����s�p�]��%{Mz;��1Y�Krr~��g�:�q��V���˚=W$��Ϲ�H.���2������d�X_�����W�l�W��=2w�c������O����VI�/e�A��#�T\Y��N�M�n���ݛ�H$��A�������z
BpYu�G$�%F��L�Sw[��gg70rE|n���0���{{� v}�G�M;ϟC���-�K*@$�T��8D�>���w��ٙ|�� %�����v��u� >��Q�E#9���8���0�ϻ٭
����k��w���k+F��)TI��\j���8J����F�:�v����3��{��t��.~8�����rB{��Z{@�Kc�ߧ	�wFG��#f��{e����19�����}r��9�jQɃ���9���%�f��|�~.dpS<����}��������I���W�grL�M�\���8�v�f��s߷���@���gIb�o�>웑������� t�_{�!8��Ҁ[�$�Sl��l�o/*�|�@���;�I"Pq��]�$G~���lv��Z�{�$�j"��ƶ��wMW��\!(��9��Ěѷ�{ϣ�5���Z�F��,�Tw<�D����@x��{�$	�$��i=o� r?����l&�~��Ih�f��tc�DX��ܭd��h��b��w3�BI����$��m	���*��F�[Erf��]��؈�k@���<��mXWx1��;[4݁��buM��۾��9�jIi�};�s��o�>>�5t ��W�~����j����ų��ܹ�(i	��~6��P�q�J���H]�YY�ۀ��'���ȩ-�xb_DG7i$�;�КI'��vUv�&�r��|6ݓ��q$D��3<���w6J�\[�Ʌ�s	o��J?��3�KN��b%�澺o`*s��] ����A���\����7��m���|�|�K块6�H$��hK��H/���t`�QG���τ��(rg��zïǟ�
ݒ�k������	$�}���e=C^L��L}R���	$���	����du��tq~G� ��ߦ����"�
"��d��A��j����V4f��N��i�{÷�]:��^��>����Y�M�o`�M����ʃ�3�v���_q��J�l��6�UZփ#D;��D�O�=}^���8syQ���|��;�`��Ү60����?������:_�����e��k����c��Ȇ�:�1X�S�up�&޷��4g��3p���7�#mTÁ1��be�м7�����[d�-�[�3���;&o3�-�_�ǋ+�~gI��rBEt>f��!B��q�WO3y@���0�KA�Z.�k�=Dq�Â�}�j�t�E����s:��'�<+F��gf�xZ"���	���d+{��{xv<��r�u�9m���J��^~4��ਫ����yɧz��0�a�徃�"�>ŔeV.���Ѹ�a�qI�cb35U��$[���7�9ۂ���ox��7W���{����{Nj��=����������-�bv��%��v�[h��<���r���(��7�����F]�$�[�s	��ڌ�f�,5e�|"�'d-گ�1Ӑ���1�8��C�{\�nN횆$��p}�Ք�+����ǻ�o���Lҙ���CJ[U�\USY�Ej{1��H~y����޵��D\��Mo.����Ѐ�Oc����"��U��.���@%�ޕM�� �g�l��F �^�]��r�Z|�wCkX�\sI��TT��{��nМ�q�X����e��=;y��w<�J�>8�Ns�ąZ#��Ȭf��%��е��n6�'���sdu�W(5��O���n����{���+�F�+Ċ����Y	���T�"U�%װ��{��}Vj"a�*
�;�d�3t���������U�Nόz�{!
ɣ
e�Turhɂ�<��&Uy�mP�<���Օ��L�������̟�!���d��B����uG+�vdַ2_�y�:�+���<����>C	ٷ����I?�Ey����:I���9���W�3���vø�ް��=��͢NY�����{�<���&����'�zG�NUB�WT��^�=+[*��0/v��'�����~�>�DP^QEv���6�藽�vL�(
/
*"PM7C���������<�� ��
B)AN��]�@^�����d�^QyN��(B�n:�W
�4���Z��<��tk��j{��3��}��x�U$?�~���?����/(� �8�^��ͻ�#ںҮN�&S7�����g�^�<Q���'�Z�A�^TW��&�pe��%;�m��s�w�ma�?>ns�~�j�xqe�QiKE1d����}<�=n-g�]lv�q[����죨�s�k>��8�d.���n�ݸ� �<h{n���v��
ۢ�u�Y����i�т��3v�6�۠�;��k�z�K�2xw�_O�za��S]��َ��3�&g�=��\`0;m9�v����]<��۬�y��v�Nvy��̆n9^�K]����.g&�7�Ř�������;9������n�c!\%��QK�u��; �gs;�����Z�����Wd�-�+�#���:4���N9�m���E��f���9�r��l7;n�-�3���8[��ͫ=�#���9�Kة����= ���.��q�\D�ю'�� ��|�4w&�Y�b��Ɣq��rv�I�]C�kX���.UݔSGl��:n8����0:��Ir���]�+S�Ս�ە���ᶷ���M�ݴ��SqJ����.��*v%����5m�*v,�6��UF��4M�[�7c=b���r�v�\�����Z�͇v��Ƨ���]�cv���G'/L]��Hݜx��ɞ�a�,�^a��Y���e�ӑ�	�
uX��K��O[�v93r��b;=j:2��;۔�]�QC�W��&.�f�8{o�ls�^ �km��-�'���WS�O9Nak�ǆ��n�c��۲{zA��^ɹ�{l��ùv��ӆ����G�r�/؃�t�����+Z�qㅹ%xL���m�[c�\8����.#ظ�;���t�rol�w�6]�����y�����W;I<3sjm{$]d�v�����:s��oav ��ӎd��{e={Og9x�z�&���#l�q���.��/i�4�غ�&w\^0 l����ӫ���#�k�1%޽�1��s��s=X���9c{�l�9:��]��M���b��;z�H��b���c��a*&�����#f��q���;x�g�����y]��αx����,&Md֛֣�4�}�'��m���� u�u9.;t˞��<���K���]Kٲr��:�����8�펭��͛b�G�5���jzv6.݈�<�]q����#���>\�R��N<��tsùlm��㵎�h�zy{Uڵ�q��f���'.��M��r랏a�����J�9�\v�]Z�]��a�(n^{uͧ��Q�D6��3�Y� �36�m��m�Z�s[��]�J{zm�ֻMqXn����K`IS��f�g� .��eg�"!%�wf	}�Xc��uz;EpYW}4�|L@~��W %����E��I2�Z�o�3K�a�Ld3A����GwЁ�>w�W) LO�����m�;7�7+��
m��)J!^�"d"�ύZ/�,X���L��;�Kb	���nX�ϡ�Iw��Bh%��_}_<�F�]8�q$D��*�]�g_��8�*y�g�N��VVO���s�{{� ��6|��W:;��~�)/�t$����Q?I�e	�FM�����1 ���C�|�}�h�'VКKzfR��vn�K����w��zER�����mwgŵ�����ׄӸM�K+� �$j�2�ITVJ�����AUd����~���ʯ `1����sr���^�ւOh�nr�ve˼��`�O���ok`o=k������A�;�MC�V��{�Z�y� �˛��.-M�J��qͼ������sOZR���'&�yUXm���_]���~���ѯ/���g��0`��?X�R)���m	?-��?O��K�����y���߶�s�aK�S�^���W$�-�rKM>��Z�>�n`>�w���ϔ}���?Fnd�$�I+{ۘ3�D�_z���Ԡ-z:�C�zо��� ��]KR� B����Ѩ��]Ӹ���A!�䏩N^������^VY7�M�fH�Q5iG2D�QB��ߢ�$Hײ*����W�"�%���Ù������h���d:GA;{G���ż�UH��R�SeY�ջE�B�|�Mv��\n��]�Uc��{���En'��ƹ��z{ =���
h,��D���U�g��qS�O9���v|H�^�փ�/Ek��i�"���w�0�wV�W^7�mm�ļ�+\�+��!$~n��I@�R�v���6���r�}�<�%�IS��-�w4"I9��V�����C���ٻ�X��j��t���m��;��/gјwtfnҪ��W0����{'6J��9e�J���T�������ď"�AH,�����
�
��~�;�ֆ ��̫��^CrO"�Ii�r;�Y�I�^�]�I4�"�>Ԉ\��I �7��l}�����N!|XU�΋�fkz�jL?��:����d"����K|1����si�T�76.�^K�8n�RI$���lȈ���ȁ���*zy�����I0�u�.����M;]�ɻ;8vW�el��m���N�+V���?���6�H�{"��!/'�}���`�f�~n���LKȻF҆��_DB\�� |QK����[I����-�&�-l�zo�D$����I��<�D�V��*{^lj�����e�(D�,���<��%C  ߹��{>��lC<D�o��Qk�	5;B)$�Y��}���}�����YS�Іw��ҳy���^| ,�U�������Z����ݸjl�	��m�7T��s,S��͟EJ�tV���A��/�f�W����_��(���ܥ��~�qn,�+M3y#�7tn�.V�������� '��dH$@�_W�UG��Ɍ�H������'�v�䖙�'5��{=��繥u{��pn(��ҳ㗠*n�E$~+&7���'-|�/֍�׎^�Sv�����`��:��rhnG�.3��{sV������ˋeEy���v�j�v���o��� �}��k`ӷ�roA��v}�l}bJ��A%�}��w�׶:}3锢<�k�lM�����Va��j!	 �����"O)x#�d�U�L��~�&|�IT�
�� �FQ[���N��Y��"�ݱW�/�"~��;B��Ey,�fR����'E��E�ҵG>��%VYm{��yQwN�]�n` �w��x�$����9�J�� ��M|�c*>����[�Ϣ���D�	*{��� ���ed���}�l�@-g���� ��_G���+�#�m	��Tq���,G��Z�5��)�{�	��ve���ʳձ�F)�^$���s*�cN�W�/���h^�ӏ������O"�{^N�nV�@�p�Z7����51��?��,�����H,d�^CJЦ����,%�wKۥ�-�����ыF��ޭ&y�N�q֎܇b����`ؑ͸3�+��SO
Wv�hͭ���@�$��[L�q�s�+[�೸�Ǟ$��uѮ=t;�O��^<��v��2�X�o�G5x���G�M�O#�����6�黭����n��n�n�pmu��*M���U�8s���٨��5���U���bF��ɶ�MK���V���y-���7�Ղ��eo������`䖝�7{��{2W��kxwQ ���;C�>~��1��B��70b$��;v,z����$�(�*D3>6C���/�/����G���{�{��M|�Q"��Ț	$��vr�n�����0�y�ϥbP�σ���΍�[��+?H� <1�IB���$�K��ذ-�7�B� a�x�c�l��WX3�������e� Al9�+��V�$��r�Pbs߳0�����>��(}���iyS/�E�1J����v�����d A��wg�S���pd�x}�.�H��	��Htw?�wغ��H�͐a$@W5��Н[M�Y#���#pA�R�"�ŷ��+%�Zs�(�YS��7�kBK��k�}����&o���y�
�M�L��Z||�S��Ɩ�Ј�ҰrK+���fY�=&6 l�o>���D�F��6
��}��V�rg�o��-^t��xC�Db4��G�*�`�W·��~Ẻ�ct��;�� ��$Y )$(Y�k>��k� �g�GM�I//��v`�@��}=�{y3�߳7�VP��5!n����"	�u�%�R�l`����2��Ӝ�A(]�"�H(��y���/8���1(I�kA�_{_o'}�J�H��="��BP����GBq�8�����5���w*e~�א`;[�V�r�ϳ�o{>���w�oS�V&^����ʪ�RN"�:���킒	8ߜ]�N�d_y]|��K
���N�2)Ik��g����[w-�s��J+ ���[���~���)��jM�F�GzW�qϻ/=�D���}�v���f�9��Q�؂h$���<�S���J12���m`J���Ϟ�qXOAi�|�ʾ�����j�����w��[�Y��ѽ��`�ñ��l���+$��p����{[����u�M���g"H'���D�6l஘�v�!SW:��*Iv(��Ȁ�4�Z��ѧ6,�Ｙ�nU�y���o��m��y�7��H�$P��`E$�Y� ���UQY�����s��h���rkE(	�u���:8��W3v��@�=ľ̍L��[��y� �?,�`�<�j�Њ1�?Q���IQv�F,��ܸf%	0-iM}߶�� }�YT�P扢.|d|�Ok�o{@�GN���	���ߘwu"e����M2��hd0�N���n�.Eפ�ۍ�m�7�[�aT�7K}�yC�n�[���3�������'��$�Z��^I��M���^w��b@���/TY��Y!
�e���S~��d�K'���w�o�׶ !5�c��\�5�P�H���;�O�9�M���\�&&RS}z��.m$�_�h$�M}�;	�����S���I8�رkR05s�*>��|T
؁�-6��ִl��p��Zº 	/5�_&�?s��u��� ʼGr����[{I�n	X1͹�+/&��
�˻������6	�ja��{�W�\��|k�]��~�a���H�I�E���E$"��IcO�UL^��֮�L�Ŋ9	Z{�8��Vo�F<�����@�VDB�O+R^]�d݀�	|^Ȃi'>��m���jcD�nm��}���D��u�8�CN�J)1\���v���H}�p�$(�%V2�s���3R��	��X`�[�Sq�	/����K�a��:�	fk�����˺�RH�+�/�0�ϣ$��]vXK)�D�F%�����%xr�B($J����g��&k_�O�K�6����I;��7t�X�-�WI��Y���{���I /�����D�d�����MЊ�I$���l6��v�UK@����~��~��i��ws3� �u�e*dJ�;�kh�l�7���W��)��E���φ��	�ԍ�~S�m FO}f;��V.�.tx*4d�HP��JO��,����������2������j������S�3�.o����}����3f/o�ο�s�]Ơ���������|Q7���â!9_n�í�Ѫ�F��	!����H�ABH�Y 
BE�3U��?��/!�.�m��bҽ8����N���-ګrs&6v�����c�۩�\3��{��3�(9�p���m���W0𫓺E�pC� )�6��rmOd�X����r'^�^ν������¶2��<2����d���x��GOl�ݘ�;��ӑ.���6]��=Zy��e�vc����r�2Eslְ�.��ԙ�[�3L��Kш��[85�,m�'xx�[c�5`�v�����ϟ�!�%������ңa&���ތI$���MXJK?K�����l}aPH �;�w����Gf�i�6�x�{^��}�V�d�|N^U}}Ue��	$����癋� ����f�B����،���Wv��2�/�ȓg�S~U�o3�	$�wm���,�;�M����N}s�|���k��b)$��M��3��DBP�׼��=���ne�پ ��}��`$�����	�Y,���2����	o��zOz���E-ʞϸ���l�?�R��?3V<���6�(]~g5��G�=����� _{�Z�'����ԓ�5���o�>��v7S�V��=�9��$������M��Œ�LN��w����~k�$���]w{��>�?��5�6����O��`���>J�OO�1>#�'�飜��� p�Kd�*[%����>�a�i�[X���="$�hx���ߦ��>��#�!{�}7}r�(�o�uU2�l���_��^�h=΄��i@x(:�p�4%�=��n����.�Ɉ!)����0���$�E��`����� ��P� E��Y!�XHE$��0��������:�2S)0��iw�뚆Y����l�e�ӟ��,�5[-hZ�c?b?k����&��w=d�)�o��GŲ�,�O��i_o�d6��.��d�*[v���-��	l�ؖ�h޲r����{7��w��<�m����KL8��>�a�i�����L9��sZu����^x]�pZ^1+P�2�I���gl��j�z�/���W�3���B�hZW���n3L�%2�\Ke��_��0�Q�ZmG�%3ｿ��6��<���k�7�9��K�T�%�������.���#TZ��!
�Yi��cMq57��)���wR[,������go�e�㜣T�=��y4�S-���y���m7�d�S.'/��b�!��B�)�����w�g�9����������X�<�-��y7�&��k<�5�j�7��׭k���a����?�η\����xm����y��3l�ta�&T������L�[)��H�}�}��m8�n�����`�c���Y��{���]����,��Ke6$�ZOW��E�M0�ZY�Y�v�FX�����l�����vΈq�ˈ[-Y��u�o�l�W���7�g�-���[-��_�kB�$��-2�#�a����}���9R�*�[%��U�3���6)�﹘e�M�F��֛rt�p�ű�k�q�p�zȦ��[,.��Yu%�����6����Kal�����8�j�f���/+ԍ8�G����;��gOL�m*��f,���Z��ëe�0�ёOw��>�\\�2{�1�ڷF�Wr��%�v��ä0e˰�����s�*����o�|w_w�����D�w�J���:���0Mg�����*��w��/�N!|��9���'yc�yLcm齗���ݳ�{�ɒl�y�� ����NL���@KyU�ky���;<������{W����{|9�o��}�����"��fr.��+��x���$���O��F4���E$B�gpe���s�f&�;��\�q��ŉ���s���r��%��o��~�r�:�J���*���y����-����2퇻T��h޺֚�0�zbΘ�ks2in�cP�:��^�{I�0Ϥo۾�u-9B3v{X�B��3b��q��3R˒aBݵ*{z˨m���͢/d�nA��ݖŢg��{��{V )y��.�Eȶ� �뛝f1�nx螌�.o<�������0� $�Y��&��T�Ū��c>q���;��<Y�����;N`EK;���N�q��%a�p���쵲�<pgo�����d���˭S2�ٻ����\���q29���cm�qkʪP�f
a��E��U�=#�Z
��,�~� �_��}3rV��+2�ѓմ��7�S����מ��۸݈{�ty�)�!�2�Qp���v�v����s�|Vw�E%�}=��0k3m����u�b�uפ���v�S�(
����0U5_	Ъ��4��x��缐�g��mTx��[��?���\�?��*>��y�t�l��L�� ��p��Z���<�=����{����#萟�Ȣ<:!�_�iW�!9{��wH�����J��=�s��{����UW*�S���L�**����?c�?-"��RS��g{�L��V�b+
��Zo.��rfG{oQ!(ffL!�%����?�����_ʯ2J�6���5B:�O<������*�Jp�~���׻����u"*�ɦ��לT����*���ε��Rg!�*�\cF-0"n۽�SmziFH�Qќ�ԛ��mk��4���:�������]=��������/_ht#���g$9r����q�̘лX��yzzI	J�&L�ʢ�d�릒��'�Pv�96��2\���/1���!'�! �$P ) 
� �@����y���0�[%��]}��Y�42�h�v��~}�ϳ�M��p�g�Gu/>��#�B���R�c�|�l}��Q��S'�R�b���,�%:�-��JV���\d�)����Ke�E���I�]n�o��λ��ѝs�0�w[-:�޷��0�#e����t�m�ixĭÌ�pIi���g�ױ����S%2��q�Cho������ru��ķ)��9|��,�Ml���-�ˣ�w�g���Kd�*[%�2���w0�4񁫻���3�8�w�霙R"���jk�Ѫ`X-\:��^��WW���p��e���>$�*�e��xƞ�潜��Ι-�u%���KN��}�o�e�[-,al�����2�&��fy�g����2;��|f�?}��Y�
e2S)�i߻����[8_�1�5X����lm������,��ԶO�-�/�#Ǿ�ݯ���9{Tyz�}&m�a�%�Zs����&�L�)��I_o��2ϷR[)��f��]���l9~�r,�n0�Z^5�_U���X���8g�
m>���v�!�[,B�hX�e�w��a�i��l.%��c���ٽp��e'�l���-�ˣ���g����l�eKd��Z_y��v�d���j�}uKwx��d�m�}�dS��u���̚g.�`�߷����'��Ke���a�LK���P�6�[-��L���wYe�d߱{��y���c탭g��:���熴��
}��fvi�)<��uq�D�[p��7��j�!�c)�E���UZq}��mi�C̄"�XE$$X��RH �g	��!�-�����x���[5��?\a�Mܽ6�m�ҽ�ϲtͲ]ԶK.��{��#��@����g�9�{:���L�<Kd���w�k��e2Rpd�]�~���2��9Ra���l���}��0�al�{��׌��o-ϱ�1Vvm��ݫ9�ܳ�s�\k]�����:J�$nv�UGl�X������uF��>���^1I�s]��6�g��ZhZW����Y��-�Â[-�+��E�d�Rq}�\ot��zD!�=���h�yG�[%�	i}���2�6�i��^{�]�B��oO�\q�S~�SkO/�\z�Y�����k�/ �sY���l�Je2S)9}���2ͲS)��[-�+��E)0��a��L3����>��&o��xɶSc~���S1�����-��IW�k0�4�I�1S��a�g�ȳ��%�[il����Gї��{>��N��|8d�\m��wE�s0�4�L�i-��!��u�fQ���ZoH�(�L�[�(��[xQ���s<x�Z��޽��gY�-��L��}�d��3hX�e���[���hY�F�i-�[%ˣ�{��J�w�����[�HST�Kn%�1���a�m�!��s��R�O��n�7HN��wzȦ��[.�Ke�RZo�}�v�I�[�{���&o��O3�鋸a���>��3i���e�l�Zz��dY�42�h[-����#�����a�>LQ�����K��U\�{�`:L`�D1{9lk!�ڀ����`t��� �'�L"�rsQ�a+�� =�cNɲjhI: �Z�D��0�{Г�$"�(�"�B,r�r�q�������j�׼f�۞x��@xvݝuNgk�N�ݟ]l�x�p����:�$��3˝�8랒8q�8�$;bY��l�i�I�1�gv�9�M����ۏ�|}7e����6R�ݳ�]=�'Ak^ݰ����t{g%v�8z륮7\�u$��<=�ۗ/�hޛ�\]p\�V�u!�'ݶX�</c8�i�aî.�˳Q�07%G�kI�w�W��轝�5��,��emٷhݮCi��6�ݪ����󇿬�Z_?��2~�l����l�l��m��l1]�r:*e��Kd�ĶKK=���\e��-�"�8���>�!�0�L޵��Ẓ�M�>L31~�,�hal��מJv���#�m�M�����x�!�[,Bд3����9����n��ͧo[�O��me���l,���hY�Je'�ۆa�ˣ{��{���!�I���}9�u�!ok�	x�_<(�9ڻ��	*�-�|xƚ�1[�,�%3R�Ke�RZ{����l��Ke���K�3�������9�3�w{��L"�2S)�B�l����ȳ��CL�Z2���ĜN2�_{�Sj�k*z[x�ciǈ՞���|��ϻ[�{�iL�]Kd����{9a��%�[bZ��������l��d�\�;�{�-�g�.�&YO��lz����,�%!I�����bƮ��-�d��=��l�!�[,B�l��O���a�i�kF���osL�%2�|z��hP�%2�)�ɢ���}�x���Kd�
��l��q�wD�����M[���[眵?i}��UcVB���)eWN�H�mk�C�^+��TU&1KˉeR��k̓~����`�2i<�Ww��i�%�S%&��}��q��%���e���=�C�%2��`��낞Yކ�hO���E�CL�Zl��N}���pN2�\�͕gͮ0⨻��gr6�O�~�Cc�m�T>�������ӫƉ=��v%�q�����;"�i��3ܪ�KzqY�n�\�Η�ӡ+/��������o�^�7ىVj���(I�t�Є��R�	"���d (��0�o��
�@��-��L��߿?>�8�d���-�tw���6͛�-��%����=�4��l�t9���a4��i}�5�t����1Ì�pai�k��6�d�S%2�����6��-��L�־����^���0��p�$��m�&1G}���2rp�l�e�[);�sӴ�%���>�$p���]��k�N<*o��m<y�^��~�$�j�k��3�p`S ��}� �h@���M���-�V��h?||�\ (�Hϳ6��h	�[��>�tS��/�����l�Ƿ�L8t�2l.��Yu-����A'�G,<Y���N���0��#�",[��\d�pm����-�]s��6�2S)ؒ�m�r��dP�%2����W�}߽>[��ۈ�r��d�\h�m��n��\u�5�^�6��aeo�{��称�~{�|�I�k����2�)����i�{�6ͳh[-��L�9~�,�&�e��\{cb�M�)��to����Nr��Uʖ�m�-;Ϲ�m�M�Z^��-S�o᢮�7HN������f)�.��p��k��}\�����ߒq��Il����i�}�CL�a��[W���0�F[-��-{cY湭	�{u���sY޳�D�-��y���k��)w4a�I��i���ݳl�u-�˨�{���!I�<�i��i���s�7���+��"���4��Q�6"؊������UH#"�5��{�o�|6�f��C�c��p��-���� 
E���$Y
B� �o��@|���X}[��a�j R���7���"�X{8�t�K�i��r����3�����k�?{����M�ihu-��;�0�&�I���>�,I8����z!�� MG�5�=��������xP�}�*���;~�$d����2��/��YЁI�JOw�}�bM�����8����-��)��wz�j0��;e����r,�e2P�d�����}�lf�(��v��熯�Ǳ����`�q>�`��f����e��j��	�F
��Y-�׎|�V;\,������oy9HQTB�W�}��R��Hm��Ͼ���M�R?w%��Ľ�L�n�ff�RZ��7�w9aL*�jg�Qf,j���m�'��o i&ĤY;}�Z�W}ܝ�JH	H���E!��4�/$;����H�%q�j㷲���.���	=�r�N��Cwx��6�k�}��)��C%$����0��>|:���]>��ۛ��~��P�$�O���"��S%�Zq��->���I����hl���^-DG��>
>���Y���06�a�`�)@}��9J!I����s�}�M�RAa�߷�a��v���mQ���i���d�r�<��?ݹ�n���[ms�h�I�b@�Bγ�j3����*�u��#2njbh���)LV��~�̀ ���X@����C�%!B����I��0����])�^L^#�m��Rg��^�n!���JL>��y��L��|�s�y���@�AL}P0b�{?}�7� Ԣ���y�
75�qrY��Z�?o�eP��+n(Tb��};&��Q�Soa�!��ś��!���u_]�����qn*��ǀ���g"�R<�I���lI�(IL)%0�r���a���������⹿x2��dR���Q�����@���V�L[x!L�4,�]�@Y�<K���^y�լ���y����[l
h`RW��{@m6 RWj�ӷ�o0��R�����c$�cce����||:S{���V�I-�x�mzg<�\im%S%2�v��fd�)�BR��y�~��,��|,����
o���stR��;|��:`RT�r�g(�����` ���+�_��T�ٍ�� �
aL�&��� i���Õ���a�����ZKO���"�÷�}������ZAd�I�{��@٭cCG�F*�
��а44�ڿw!��awR(�>y�}���=�j��T��j��Y�J�y����)
��u�[5)
IHP����|,�#�xp��_?���LU�	��Wb�s��"Ig�s�~��F���g��u���۽�|{�{p,:yl�+��%˺3S�9=��]��kl,�QH�~�I"�X$ ���p(pq�ޯ���U�%s�z=�91k9���^ƪ-m�璤�ڮ�m�����y;i{��)�ܻ��㗳��7I�.�:ñ�V��Ξg�ϮM�緺9[S���5)�H�Y����L;u؁���li6g�pf���5qC���X��on;-�j������hN�I���/ۤ.G�v]@Y�vӞ�î.��<�qΉ�Hc��˞+�6:gNO1�NX��vyY�f�`x���
���[�{�A���
�p�ǚ� ���u���JB��۾�0�M���G���B�X�y�.1�ɜ��9ԇ*�g��@��%6$)�=�gYI�!�E��:5#�:�K��ZKZǾօ: S ��xs�o�m�S�ȧ/�s'Xe�$�	)�O����[)%D)%D�}�dY4�d��d��(|�̋���{� S����1"1����_׽䖐�Q
*�����uD) ���k�u�f���s�o>��`�IB2�����-�@�(R����"�C
aZ��o�]�07wx�B�
z���u�>���|I�)��Sn�̚�JS��=�{��CL>��iG��}�/^������X�?Q
ig�an�%�����o,qw���I�kzȦ�)�
e0�Zo��쁤3�u�w�?{Z�}'�:0�|���-����������Zd�)��L��O��}�n&�5�~���o;�ż���Ԫ�P������q+�L;��*v��m'��N+�����y���aZ�~S%0�o��-!�B��7ϻ����S0���o�h⍈��y��;��7�ԙI��֡l�������9�wYaL(�s���8Ä����aI����6��(H��cm�ڎ?GD��T(��q��
3��$�g��^o�����r�u���f���MM=�s,Ƕ�������Y/5��^[��⻗n�|ɿ� y$�I��X (H
B��@�fwׯd��J��
�(;��օ���� �����f�R�S��S�����^�γ�RxHhB�<
G,wxq�0�5�}��j RAeRZ{���8�hRJaC
aw�֯\�h������~��
N�I(�}�dY4�d��H)��-�M�+�<6}���o̓�� �>�fP#zr�y�NH�U�{��tB��)S}߽�6�@��
e'7�k0�s�r��͝�nL$o��E�Xg%�_.�q�����Ì)=����m%!L-�0���ɦa;��E �T���hXi �|˺;�{ف���!I�>�>�p��K�
5��w�\�Ө��I�L��N�<��@n�uQ�"�e�n�抴s:���-}��Ŏ.��|�I�kzȧ�Y�JN}�o&��(P��S
aG7�kD�.�igo�ϸ�9�i&��7�dY4�`��HR{�ײM�l�oZ�F�m1wXV�^� ��o��- �=�s�+�1����g#ꐦ�40)+��~�H)��sx��KH(hIH53�}���ko"Ì)��x6>Gp�q�6�i)5��y�m%!L��a��ɡ�d�RA`}���y����B�&?���l�A/��z�#U��`�hdd�nV�&�Y_!j��F{_���sb/�h����skMQ��ѻ�w[-�k~����$Y	�HE��Bd���=��$����@�Aܩ
a���H)�vs^N�t�-�*��`a7ﳑK��{�s<l��HTd�����Hm%0�Q����-��%$��$����,����S�|o�L:��d��L�\�I����'�~��r�[[���\c��Rӭa��bs+�(N�5�J����%2)F1���6�IԴ�@�R^��f�2R)
�{��,43)���������,�E3�++u%$��`Mu���.�U�� w==�c
�X.t����ߟc�����������<�{�IpB�(e0���ɨ�2S)�BRO���B�,��>�.�TD�}o�9Ǒ��{� 4����B��=�wy��
k��k���X��4�i=�oYU ��d�w�m7w�2��s���$�W��u�ZAI�)��s�d�)�S%a�Ny��{H�� Y w���_2b#
��а4�j��CC��U�����GU!MA�M
L}���;�{�π�x@�N��}��y��q���%!Bﻬ�
a[��cbuq����0�`�|���^�������P)�,���y4�$q)�% #[��(�Q	!��� ��{gkM8����g$�ǎ����F�xgn���0��o'�.ȁ��7���_���g�N��Ar�b�sS8��38�v�w_�	��AB`H��� �`Hf� Q�Q
i��{0�Q�IA�=���]7��8�M��7��)�) ��{ϲlI�r�����l�I�)�ox�5a���
IPN���E�L��i��GWϨdٯ9��S1�8�b6�6�ësv<y$vtr�棒�t<s�K��]�T�ۥ�ӳ��r�[[�y�/����ND(��w������
J��s����Ż�vb���u/��3f�JM��-��s�a�aL9�s?]��񁻻��Ì)7�k�>G�D{����������CA�
% {��r)�
H)J���b |B�<��^�*�����}���
J�r��`q�8��:i�'}��"�@�aL��I����lI��£
a����{Ʊ~޻�-��R�>����&�I ���{�&������/wxV�/B�m�1�P5�M��_,��G�� +*��Au�m�I~���&�%z����y���sZ�`����O!i)
Cz�0i��
aG3�-���1R�:��m�&��}��IB�L�n���f>�����.;��
�����&�`SI
*�{�w l�j�SQo�amh��K ��{oޯ��^��n1��{�CW[�{��{|��)k�<1��߽�F��J� 7˥���7�1�2L�[{��+=S1l�u;����z����q>��{7/uǛ��t�gDM��Rl�d:܊مlf���+Λ�"��i6A��6 ryl�f�.���}����%��n�E�<��!M�h8�L�b��brTh!Ӭ�u�qW���;VH6�m�T�o�Yӳ���[U�!M��e[�$�=���%'�T��O�/n�����<�oZ�Ǹ|@�S���I>r�i��n���瞡vArE��m�+�������4T��sl�v��x�4x]�>�{9y�F��٭&��z�PټB�[�Ƈl����&����Y���y�u�"���_�i��.K���_/\���V5�|�>��8>��5vy�	d�8��Q�|��9�N�z�v	ٷ�����7���"@�}��f����+�u��\�<�MpD��s�㛡��gv�/�vL�`Vz�|�S]ĸ�����^���_{���n;U��.�yo��秃�6�MFV��Y�f��.);.��B�2���i�N�;^M1��c>-��l�שZ0������r@�ޢ��^����옷��4>$m0�����^~(ܱC3���=���tB��(*\m�m�,��z˅����g�^���a��nu��=���]�F�1�5V�V7�d��/H���E���)�ɛ��T��n6ҝ-f
�D�F�]����ïn��Y�YUbY�0��)�=���sJ�"�*Fpj�ę�m����#�D˦�%>�g��)*�AL��aM��<C'�����C�=3�:��3R�M������<~?Y3м�T��I^ʄ�i��^�s�R��������߻��$=?�n�ўɩfB�	�$��WeE9�ȣy~����|����h�LMD��a�܎yeN\���Qmv~�����|�=<I$W$�4"�Ĭ���F�"e�ٶaTrXXn$'����M�_�=��e�'��Ѣ얕fz{=�ex�Kb��}����R��&�a��$��&E9ѲlC�{���'�K8��￿}���s_����L&MN ��B�!5�&yd�b��F�T��F������ڡb�d�QI�	:e|;JI2���a�k��!�Э��n���W�~Z�j���qa�u��\k�v�v�=����^R�����d���.Ύ�b^j"��/m�r\[���啌�[��N���6�s<�66\m���`����xMex��_c3Q�o�z�~![1�5����]���7V�:���u�;��>��%zQ�����Tq�[��헛�n:#6���ᬝ��"�q'`qed�q+�W6��w)���쉛q��;W�1v�����.��ȳ���Z��(���!���J�4��uI�sMeT�u�8��x04���;g"C��Ԝ�.�^˝��<=&EP�������;2�Hn�1]��[���r
۳���Ϗ3��D'UƠ�V���z�Wj��m+6YXn}�6�%[���b�7ᬀxM>�,h�"׵h���l�x{t��>�����ͮs���u��L�&�c3����	l2b�cOn�_I�TX�|[ã�u��<Lp��q؄1Q�]np�7<���<h�6��3ølOX�7Y�ݷ;!r'Yn$��q����{f0e��u�m�f�={�֫]���q��.�;ĩ�`�(]�c��F�7aN܇�$�\�7Zq�I��ݜ�ȱ�����l�s����7/���Ev9\����Y�7<�d{��m�X�ʝ'�g���v��n7�����Ia6��cl�Zwd]��a;n��9�Q�FvU.+gs�2]Z��j�{H.�K��E��V �H�\�Z�� g�����Q�񃬒����p����B1죅�sU����p�-�ޤ	�s�x�n�\����Ht�i� a6ov8(X�ы��q�)ۊ˿�-8ʻb䍹wm'm��]���n� dc�s�n��9�.}��WC����2Nz��Iax;]��Kۜ��pqn&(n�5oY�ZN�y�;�x&�;m�Ok02�Vx渳�Vֹ�I�g�=�ɋ��.�ޑ�d���5:Z�����k��vsÈt�+x�
�չ��ojZ�k0sɷ<��b�P�� E�"�E�A@�x�^8�������ox�j�Ůs���ΊѸpIYє�h�Su��NLGI�fӣ �M�iI����QV�����u�N랞���I����i�y�y���9w�玡�9�S׶��q��zAʲ���ϰ��p�WK�ؓHHn �����\��!n���#���{����`����]��k*9E����b�e�5n9U,����v��n��\��.�J����;!�i���s�F"��o����������]�ǀ�o_`�Ag��L�eN���@��) ��sx��a�����Z�u���M	���Ja�[%2�(���������Gk���.�]��84�|E� ̑��C�%�,p�����g��Bam�)9���I[�-)�Bsx��f������X��ڰ>#��>|���581X��W!l8�k��n!���2Te0���ɦa����BR�-��1��X�3�l�&YI!ʣ�{�d��Q
�����`R{9_��1V����@#<G���Eo{���o^����al�JN��}�pI��£
a^�>ޡl<m
IB{��2p�1�z�ϯy=���N�S%FRwײM�m�w��k	x���5�Z�a�_���p���0,.��=����k�8�pj�F%s�ߴ�b%�۾�0��L��D��{��0�����o�o7gѭD���*�eR�(#�	�y�mp�{�e��Z�ĭ��j�Kt�����k��1R�>�Xxe"��u�CbI@�0R,>��y4�2P�H(���,4��S���6��r�
g��2�
A{����:`RT���<�}���U��0�Y�0e:��l�JdM�7�£�wU�����;2�fxu�L�P��|�7��H6� FDN\,&��<�w������b�p �k-ۭ⹗7�~��9t~�@ R ��
X@#'S��w��$�AH,(���z�weB�P� sߟ`�&�I���Ͻ�}����b���:Vw��}~b������L.���r���T��pgEILR
��Dn�حk_n���"�� �0�"	�V�������-
�{�4�Xj�+�?U�q����j�C
Oco!��_5�R|S%��{��	IH}�pe����HUQ���������}��c���;�0�`Rs9__0`�0��^+ iﳬN�f�\d�Td����y6$�����c$�0�j���i0��� {���he0X(2��{��ci���������}5��bp�5��w��.3s�+usx�z�}�6���v�m75[���Ѯ�����%|)��<�0�C�Q
*�h<��2�]0)�%����H)�;�}w�__i��@Xn��fH"�)
C��pi ��}�,N�1��q�4�Ͱ������IHS&\��"�w~���q�y" @�{�w&�M$�J��{�����<��`�㱏�+�o�_�k��%�&��Y�_U*���I*ךƯޫI��@�L�JOw��M��$�|�����zjh������^�AM^���-�Y�)
�ڔ-E�le�r&�E���MÅő� ��)����靈
��f�˸��:�=��!R�h� C�	"�Ad`� �dd W5��l?�)*'ߟ�����~��0�C)/��w isK�}~aS������oyKZY��E�﷭�o�HnU��s���At!��`RQ�}���؁L9���esZ���מ��II<��>��aL('��>��%n�9%9���������R�L���y4̠}��Ok-��Qֵ��'f��N	h1���H,�$*U�~�@��D�Ї/~�p�zO	y���{�5�#�u��	��ϳ[��u���ESf޹�<��C��΂������0]�\b��6�}���I�I�[-��L��Ǿ�M�6�	)IL,����0�L)#_?}x��>LY��M�׹�d�e2P�N�������$�M�V5�ik͸���8ĭ�cL9_:�<,$<+;a�u��:"X������`SQ�IG{���M�RP�L����0�2R���]g|���=^���Q���buqx��u��
M}�}��I@�2Te0���>�<	 " �����>Ϥ�ٝ�F7���X`Ti!UG>�����
Ai^������^z�o����E��\��,������:���g̔�����dؓhP��V���5RAI]����6�^�{��Q�LU���`�w9.���D���]�j(h��$�������#x0LL\�y�A��@�Zγ��B1����w��BO�$X �d�� �I �2~�|���?���:�q��_W��q���1�F��0����ӖaLY.����2�]�.��o�� [�%{=��>JND
e	�緘a�d����{�I0�<.M/����;�4�8�mLR�i�d���k���n��+��&h���d���Ue$�K����x\`���^���x޻�؆�R�L�V��M�A@��
>结L4�ߦq߬��߫�Cꣾ޽�4�wD)��ׯk0æ'>֗��f/�6�"O{[���2�W��G�����f��=2���z, 	'�mE|��b˪5�۴bfIp ʈ� ����]�(��"�;AK��[��AyY�7��}���jR}�t�b|��Tnu;������`���͆t̺�AHf��$A}�H�\yMG*v("��3��,���#�KIK3���e6��wV,l���x �'Q8��-UdQ$�n��>/����tcPlP˩���TD\e{r48<�O���{Ox�c�����[�̿���.�kX��7u����c������_u���5eR�����H��X �E,�L[�]��/L�m��C�{�t��Y�����q���|��+��_ Zyݬz#�6<�#l�E���ۈ�L�D��C�������IL;��)�[��.�^�'c�*���}����k�Բ/��x�M��Q5�:�'s�+�=�v��T��
��sbD5�����/]�h=r��k�t
������{HNey�{/�p��v.<ӹ�E�{]�s�Ջ�K�nD�����+��^��K}�ߏ������mzM�9�b�{���2G=�:�,f��[��+ĂC��<��>	 �����W���'��d,7gz��I�j��w=�`��y����;_�I�[3I\�ڱa��ն���	7���[��aHP/y��1i?І��Z�M�����O6��b�I ��
:z�]B��T������&R��}�����2���_����Z�����F:4 �ɘ��7f�S��v�/�7��z\���	9���I���qF���ữ�m�yR��Bc�ݸ����uN�6�n����k�E�͔s��0�N���;�7F�	n���讷�`C�yɀ
z�(����Z���T�����>(��p10D���9�(�\	Ӎ`Y6$P�qXE�q�0QPdk��vxl75y�(7���5�N���5N{d���<Xvn<s�"�.�e�ǀ��� 
B, �a"�E$w=��~�C����$�츠H���8��N�&hGfI�(�D�@��$�=�RI7Z���ur�\����D����$��.�q�$D	&L��`�������_c��4H���A$��pi"�gmtɫ9	�O $}�ه�Q ��D)��=[���٠qըz��U��"n�]����Hy�T���t+��9>�����e�}�kd�QJx�펛����6���If�0��%�,*���l����o�������u� ������{;j�̥�51Y5zg�A#V��C��	&�D��r�Q&���S�W�>��ʁE�l�2�8e�ܲ�+j���'WGI���XB]t'�V��R(3H�Y9�O��\:9��%re�H��ޡ��L�K�(���kM7P0�ZZ&q˓WSm+�.��&cKLAuU	�"0���@?� �E�(�	�]�c��츠I?������������힊m��'���8~��$�ݡ@o==xm�ʐ�A-e�P'(Hqd(����w���-��/s��r���ِ�*ڊ�$�;���H��wy�k�Ϲ,���ƙ�56��B�q<=�Zݴ���O<�u�"i�L,;��ږ��~�__���1Wxĺ�O�O5��1A����#�>��B����\�6(bD��B�Ӣ�xJ�����v�a���j�W��c2;ĂG?���Oo�lXK�q���joz�ދ�r/h�݊�9c��Y�g}��h�����Ch����i�h w=�$s{w��éZ�b`�1wJ5�7c��|�Nu�ǒO5Ւ	 ������]w8nD�� �֒���Nߠ�5y�5"9��~�pRXtl�g����$��p��QD�`b��{7���u�f���jr����}�Ad���H,���/5�d���R��d���DJB�?Uo�,��w���y��
�и���z�X$�]w��ۗ�\��
Çl����@u�5�{#���[����=��k[��]�CU~~���\A�D�̇��=�I�<�Y$����U-8���_U�����\zb&g���9��hzq"91���9�\l���VO����b3�7�.Ӿ�=|0A&ĨRA��i�;��E�������5᷹a�1݀�H/u�A���5�
�ś��@KRZ�����zJ �n������v�
��ˎ�2Rkr�?K2�o��I�0�F"bM�5�Hf :��fmFl~���g�L�e?Y�>H���TVۛ����� lGg�#��SR���s�ߒ�0�q>К���3��> ��gs7������۹�s���o�����W�;�_�� ,�, Y"�
B,"�$ɬ	�X��3r��h��xԽ�ɜgm�S]�v�6qd��y���J�rv�l���\r:]Ã=��fӣn�93��u�mۖ���k]�[��G7b�A����Bz�A��<aǶ�s^����u/�������l��ε.N.����=��9�<�:�E\f�v�N痛�ݗ]���<������D�j�����sغ1�7�����u��4=s\��g����@^�WL��������j���!j���,��RI$<�1��X��̪�r�mۻ�	�� nP��0�Pd�337�^�L���Y�	U�駀Y��r�$GgUP#qR��}�F�%���}������|>�� A7��@�bEm�V�;��F���>6�7r(<�f�$��^�X�bP3�Vi�7[�zeV�����D�����{7j� ���j�Eު�倬�u-Sw�F)8�QPb`�31U� ��/��
����m��y�wA���x�Av�'��\��q�֟QT�Y!jj��aٻ����j�m2��mتUڂUB���q�~� �3s�F��H'^������)���+Ā�v��MX2$@���@�˻A�P������;���V�y��]\.�;�)�{��y%���H]	}�)�e��>+�9/�����h��WU"-fM��瓽淾��� ,�Y�"��(��w�����̫����45������ x��/m3y���BJs $}�nȤ�zu�c�ԩw����D�A|�߬���K�D̩""H"�������+Ɨ��lׁ �@���vH����!�}�O׌�gەD��@1Ĩ�|n�>�Qa�;^��&;DF�1��8K��y��вC��ȳ}�/z��Ӝ�[��Q6씃�=֮v&5�	Ѭ�絓��P���c7�p��7����"
�A%�=�6 :�� ���d�{F[T�`��r�'{{b��)ʂ�ELĚӨ:B�2�-����s�_�u�Q�\��I:���]5b��D���JR�\�زH4�fX��ǖ�x ��gGO}5l0T�l,7�E+��1�v�2z�~�
�Gk~�ږ�R�5��bv�sc��[��.
-��e��d��1��%z`e�N[36EG�^ⱅ�ވ���y����xw���O7�~GA����� 8�D;/*:]�qmFG��m�N��H�ې`�W�4ҋ�'N�{rK%lc�J�Y��^�2�TC��DP������H.���ӱ#"g�p�N"��,��f��:��^�m]V{K����窝1a9�Ͳ��mF��@I����쟵ۑ�܄����2�WgF��]B0C��R3�e���eg!�w���y���w�X�q��"���)�H�"h?;�C!���)���Ðe�5��}{t�x���fN�6�FF��k�Y�_{�!����(��2�.��/t���y�a����0�Ή��+�
�3jB�VJ�H݅T7(6��A�]�(F�����[N̓[�7ټNzT��wb<�Sx�q�f��"H#�=�A����?w�T��&����|��v%xd�6�xm����_���rS4��w�UOT}5~�޺Ъ���s�.��6�"c��on.N:1�$l2�5���Kmݹ*�&�M�ԸJ$[y��B4�F5�EŜCc�'}���r#F<8�ԑ�T9y9�f9���d�˨��n�޵� ,̬	d���ŪcX�����U�lŗ��֒�����oww�{|I�}ޔnh�<�Z�����,��Zb�z�x/A������зF+�w>�~[+�����b��)y�C5љT�)�}�b=\eyx}Na$^�Zz��/���"{�T�<"St��)	B��e���l=(�"�vzU�ۊ�Eo���||/0��ewS�_���$PP���H�a��)����'��Ao����~I.r$4)��!LɜaeW]��W"�]rU�И�3(�{���qU-ǜ����t�=IvV�*U�t�U� �)UtOH��<�W����<��S*5~�NEz�����Q8Q	��9�yy�Pe�Zkiy��j�}���!��<��=3��,�9�,���\��i�A��k+�[����"�?4��<�J��@�ĕ$�
�׫�ʇȥڑyj�~�߇�'� QCV�!�]X�D��%�J��֍�pG2O(�I]p/
�\�O����=!�ȱ��%\�3�V[m����-4R~ m�(E)H
P"�����b����5���p���[ǲ�luR����_{Z����6��J�ܫ$wqD�gmU���z�[�?
����d kӉ#�6$�,z�>>7�f�f�Ɍ���9�W�0�5o"��v��!:�c��;]v�$��`c���䵓��l�r�榹aK�2Z�Uc��\�Ny�ڋ��<�&kj��

�xV�мj�݌���]'�ACV�[�,���<y�b��z,'C*�(?��+��~߶��
�%W�2��c�/鞨�8V�ELěe˯I�{�^��l7Vp�R�κ��ǭu�`���ڢ}4!h,ȑ�	J�e]���c�L�Lث+����v���y�q�[8�d԰K�gݵ����gG{�aV�q��F��<a�&�^W��������-;�]^�}x~�k���dX
 ������
j�}��w�hk��1�0�]�zF�����F���q�O9�j�I|wf�A�����k{TŮ���>�n��x�*q�]�y@��\�鄺�Cuϛ��	�t'ei�]����m�֥�5%i�'����A�{4O�=ݎ�Π�F,�]�y�P���@w^�Eu`�@1���
|s���z;�����O�$v=���A��}�,]k�ݽ������k.V�g��aHWlV�N����o�ZM�g�G���j�I;��@�H=ݎ�f��]�V��HLd��*�C�k #����H�;�]v	�>ʎ�p+#�`霒���/#�P�~*�b�(.f^�H����Av�=;���� ��|�аHQԨ�����Iq,_C�(kPb��?v��r��**�n ׹�1��a��|oxG�M9��9��ף�ؼ;��=�����}=O�E���#�C�����PE�7�)��dy�������h�g��͕���z�k>nI�5�c��v
��`w�cg��0&����1��n^;{z��̰�k�÷�Ѹ�0�ɲ�S��]���{�����ɑ�+�Z���ȞN�W3#玎�����ص�Eĸx.����x�6��Ms��tæ�mu���8盦��'�?:, �P�v�qWo3l��Prȍ�q�f刧�n�Ӭ˴���
�ŭ�n��'X��s3����|?#�H��D����wT	�>uvAK�z*:2�GuK^���� �y��Y�������"$�0K\�����-�;5!��8��Y$�GR�I��w۳��#�I[d��3!O�ٮ�t,�[U����g����I=�������=�g�w\=��ح��z�
 �CW���̻D 6��P6�_�>���,���m9�sٹ�l���RQ3&�)��F����uf\aS��"�������E��T����Ӌ{s�ԫ=���jz؁�X����]'vr��mG]��g����f%�����+~�;����v�t�O�D�d ~g��Qt{�7�{�e�g�unX�@'�j��ț%A�b`�337`mu�A�o&�mmJG���u�(�&u�y�k	w����ݘ��2�-Vn�z8�{����D.�YLH-L)Sx6�M��P�?
E �� ) ���Ms]�~���~�+��~٠I����xGV[ݽܫ!��:U��b�K�"m�k��b;�٠A7:s��"Et�Q��ج�o�f�n�B�T̅>5f�W[{����Z��jqP$��hP$|޼|Aص�y�&�e��5�++rƭ������O��b��g�\�uUA?7�D��7`Z��u���l.x�*H&bd��JN��<��
�Uy��V�r�7��Ÿ��b^�����g�T�	m{��{�i���\�PD7���]�/�]0��=�u[j9o������VLg���+#��o�ʩ2 mI��Q\qB�TA۵^'ăϛ�X�{�߳�}��fVG���� IM��wF�G���|݋ ���:"yE�tp���R��A[��_,�âN��ڼY(ߍ���gr(�h[�$��k��yw���+]�w�����Ed�`)C:�y_�揮�����?�kv,�D�D*`�A㴻Z���Nws�MAq� U��v	�>ˎ�Kn�ʞ�Gvz��zR���B�3!O�`��߬���C����R��b+��~���w%x��Z�՛r�Z�Vo�������Ն��b�*�ңI2�nѻ8I�n8�az�tz�zF��__��V՝Q�}�"�j��$�|�ω'*:�DnA��k�(W�;���e\���52L�fN`+VeA5f�v��ޑ��6	$75��	9Q֫�U��)���g�*� `���&��)J�\�ݒ}��;U�EdK�P
鞆�A�'n�`�QҨ�	#O�@�\;��y�p]����6jE�A�̻�>'*:����ξ��kc#�p��۝�U�a�̧q{Dm!�2`Db��8&ؕ�-�7��ImK��V��=��C���D���F�30���1�9Ţ�Ќ~��DQdAdQB�Q��ﳨg7��*`�A����B=���n���؟����$�ȩJ�:��������vBe�S�18�D0�Mʣ������;If��{<�5y�
���e�}�B��-��|��w�Ҳ	�Ś2����i��F�����	�˶>��Vj(���l��0�ۺ��ݜ���> ���"�^ŝU��}��Ռ����ϻe�O9���mt�U�]J^M��	&�vk�bۡ|�_�C�ڻk)7�7�r�ʆ�2�UT����溲�M���'�D��6k�|y�T���r�	����T�F'| $���q� �%�vjzo|�5�Fb�F�Κ$�6�|^wm۞�v��}�!_`8Z�Ρ]
M]k�=[���xR��W�A����L�W��rz}��{�^�X��jM�E[�5��qw����gn���ڶ���"�R)���d<i�]8�J�Z:�ɴr���p�l���͐2�m���v�´r�+�w���9�-���S�-9����8�BU=��[�&4,��A�FE���0r�F;"�[;�ɀ�M���{jp�;qnN�6l]vų�g�����_bGiGe�C7]s���v���s�@d�WZ�P��u�s���Ԇz�#�����`Nғ�jwv��w5>,�;S��!�mɤ��ֶ�ry�I�t{r<3l�`l�G7j[�����rY�m����/�������2�A����؝ۧ1"o��PǛTO��$����
|n�Gs�.R��(۰�w+��"	�#{P$���b���3X̙$��=6ό̒dI�0�f*�]P���^����J�F(gC*���#�mQ>�{Ѷ,�W�\a��`%2l��~��)��P�'j\��~��I$}��v�?�Cjn�Er��~���`�m�	Z,AD��������W� yq��^ ���߉� ��0g�
�p�$��,��絜�n&��fQ[%v�u�����C�U�̗\Ń[�ب�m��.�K���~�A���&I332�:@7��vA>'/����F�M�
� �om_�b� 4�
""H"�n�6��F���vt ��͜y�_^0n?z�n�+��-���ro�{|�{��窍��`�}%����Av�_d3x�p�B�?�f~2(X��ߚ��/?=�h�w�����+���l�uM���S2�������E��L���N� 	}�d��,�P�Ҿ�V�bD-)&�_y�����<����L��C�	᝵�c�D�En�=��"fy�3~�3)�`%2lqx�=٣ݖ�j�kY;��vH$;s��$C�ڣ3�v3-���6ٵ���(�,UH*��u��n�fڮv�2���F�R�2�f�~�7�ߖ���X���˱d:�eI ������Fg�Qwn��!��M>��F	s�@I+s/�xƨ=^^1���D�2�h�$��� ���7Z�V�A34N6�Q�IZx�������\��\�M����z�Z��18�'6S�ێ�˾֜a�����:ش��S�r�MM/l�[d���?/Y�Ӎ��^�^[��Й��lӫ����� �@$�I}��r��>��X$3:�A:�������d)��񬟸�
/ge�A[Ѵ���T	��{Rq��0q���^D��o��`d퇾(�bD-)-�g��}��'k)���{��W��7��D�=��ގo��o�5q�*+hK���ep���b��{mz��v�'g�i����d����߇����	D̛�f'h��@�F&���{���,��hN�R�A{�"��T&H�fJ��'7�Y��h���"��]�	#�ov׬y�u��+���5��/�r��D$`1$���{�߳*�`G����� �mY]��n�q�a���� �x������`\������s��afdq�ޚ$J^$W]�㖻Afk/�AƽyQ3���i��u��M;]��`ĺ��(^͛5���=��E���~�0��8�ч������5T����f>�~�W��b�(*(�Qt��Q>qB /��L���o�d�]����͙5���Q�=)��:%�H�������-BU��a���$�Ĵ�l�����5��<�vp�S�����\�=Q7����&D�S31¢����|w{�$�r�Q����[^蝪� �&!�v"e����&d�	D̝��`�vnX���I$oؔ��&���0|�X����o�݌����#$��+.e�>$o���	&cgbbzc��H 'w�&O��1�23I0����sr�㯉��$���$��� P=����Qѕ'��x��yvLf� �kcRV���}̫�o~�j��I�HR��qf��A ���@�<f^;��Jm�_�j��=��ʖZ�'q����n=*��1��f�.�$���7��#=�wTf��cI6���ӆ��,\'"�#����G�x���9~��°�@�*\d�lV\�!%�Cm�k�i��& �c�	����}Ӫ�
v������͞\�;��������Y�i���q���ZU@�	�no�^�'~��N��u�Y�-X�9�._@HʿHN�������0�q��sM��G-��Ή���1�������W��R��^�{�a�Z��Uνtc��Q1B�9�>��{Ưg�
�{�𰐒��x������lP��{۽�Ox�#ͭ�m�<ovh
+�]ح�Υ�ê�naȃ�Kc(�@������s]%X:W���l����`Ǵ"��������W�L��m�0P�� K���~�gy=�h}��{��;�p镚�6~��Nѝ^Fn�z!촞&�w��wpX�T�n��o�Hb�8���g����ުG#�eh���ۅ��V��^1�b���ױ����+[��\��Ĺm�qT�q��v^�?4�z���ד��5��W��}�X7Cr�äNX�<�>��V��g�1��Xv"�cˑ81E{��ܣB����J/H���Ɇ�&���p-@����k��@>^|�R��Jj���%f���E;���*���8��E�3;�nY��yM��P�:!�����	�� kWK^&iü��V��Zʊ�7bs(�#��k����{ol{����SA8K�������mvp�\.�Ʀ�\mѫ���o����~>�!W�-p��:y	�zIEv[2":�V�έ��{�Z��s<����!r�=.IxUA�r�VxƤ���v=���}��߾�S��T�o�^\�9����j�S�^��BE����Ч/_F+��ۙ$�L�h����$��z���������l*�s=�R5Ң���:��d�f��g�S��Udo������E��Ē뗵�1G"�"��TP�4v\�U�����'��b^�T�aዩ���\)T �I5���7L���0�v������2�u��S!~�0�-TG<�#��K�ڕAuH�(���	0��PRA ����j��\��-5Η�`�Mj|Kc��Z�3-�ۣB��:Ñ�(1����u���c�l!�0�2Z�ۧx�^ ov+;-���]��]pUM��7X^M˻s-��)���Zs���(�F|�=�`�F�J�+��s���]�����ֻ��jnŹBNO7��t�¡;S ���V�c8]�.;i��f&�2:�׻$[� ��f�Uw��j:�qv��\�!���<Z�Z92�Aӻ���8� �K�/U�Wq렻E�5����ld��ٻr/b�#���v��N�>�g)���];m@���:l�9-��.�x�&;qf��c r+I�綰���[N����Tԇl���n�����*j����nO8�v�sΜt�O��Cy�ا�M�'��.�-r�|����Ƒ3F�+�>vv�����8N�!���<��ˮ���9gq�����7g��y۸�˹�v�	c��bc^��v����-6c ��v+�%���,��x3�\���nK�c5|y���έG��{�j��QKwo�ƌ�1Y��5;(Sl`����>�f�gM�Nz�C�`����55�m�>�F��2����k����^]V�;Dp�9#���[l��3/3�����1��!�#z�����ԯ�}a�Mnn��wP������2���v�ۭX��m���/n]Z���d`8���f�\����+�m@k��)e]�1��q��۾po����OU��Ft]՗n���ӭ��us�m����xs]J�zn�p��֢�\�]�U��/>l��s��Wl���h^��k7Y�r�8�z,&.peN
L�nܧj���c�:7��ۮݡ5�a��m������8��)��:�;����RT��v����ŀJչ69'�,OgW�S���W+�ƹJWun�\�h�b��t�:��Ӷ�����=j�Ìbґ-v��0��;�2T�V�d�(j���j�Z��uvFn��c�T�����NWhUo���v�v���|�l�m�W � �6 S�η:݇s1w=�g1����K��^S��8qűm�qt)�Z���
�$�ب��8�����\=6��.mn+�۞R��F6�;GY���l�Mz��;Mͷ+{k���^\��v-�(����n\����D���*��T�t�̶X�G���)�9��n�B`�ҭiڝ�[h��T�ɞ׮�X�NN�=�6t�]�X<����	�ۚ$�x���Uc�����~���.?a'��vł��=�$�A�͚ �fQ:E���L��|g]��9�$���{���v�g�VgwqS�&��\����X����~�]�}1d�:r�M���4�Wku��m&>�yJ��x~��s�'����4t�gV0���"� ��Tg=�]���������U_�m��ʒ	� oc�4�'����Q�T#on�ؐ	j������B�������A Z/yؾ��Ͱ�z&V%]�A/%��@�GfuQ$�{�+/�%W#�FV7���9�Yc[d����#;��ٺ���=sn�ʨi�l��mv�s��H}��IZk���S��sD��y�:�VL��l�\	�́���Ӈ�-K5~���/p��F�f�6f��݂0S�[.�u8t�v��\�O;��hDh�%X���9��f���7fA�21�A������L��PQU�]wW�.���hM���;�`�D�TM:H?����H[.L�*T�13�Z�$E.���g.`8�J�����}���6��O�oyݐf���a:� �����$L O���i\>w~$u_dC�pgMJ��E+�^G�P��&�2%H2���~�K7�S|���}�4A���v,t�dQ�K��5����P�Ez`�bI�N��O@	r�R��mFp�1�e[����,j��������$O�����[���@I���w���b�EF�Dli����D�ۡ`�TD$�bB""H?ƾoө?��|����k�@���:o�(��܍�+_E𹉱�B`�L���+���dK7�RA>��g:��q����p��X���mw�yx�b�h�?���k6K���@�Τx�ڄ�'{��h���!i��SP�%3�VM���n0���Ă����߿~wpP:o�@�g��T�n����=b~�0
OzA�~�}q^$�y��dҊ����x�9Bv��}���ܠ̃ ����
=���^���Z����K&q�(�´r�nώ��r��r���U5�hZ�=�V��e!�;TC�Ę���s�>�L����ۓ�O'��T$������C�*T�R���r�_������/���^�|ns2�(|��z�+yj]yB��7RN}�[��d���2M�Y�s��CW�i��6
}Zk.��ڰb�wmU<0Z]� ��ܼ��{�b�m虭�z7/��7H�o"�O�y�T	c���12"|s<i�p����1׫���(_��ۯH>�9����\�=�rɘ���
��T,�܁��6�#Vt�Y���;��ȾXy��>�~Uw���ç��;#����{zv�z{ W�	A��{Q��	�~�)��&վ7&A�� ���Ŋ��TI ���ﺯR8o���o#l"K{�^�m�m����5��|��3����n�ҤV6��z�y�R�kq7j�]ذ�PWk�EKy��s�9[�����̩ ��6hH'��m��m3Qr)H��b�';Q>W%p%J�*A���<��(��rM��L�"s���VomA�p�=��<�VvuE�S��
#
��������E��dK;���A\�^�Q~'�:��O�=�g9��؃	!�}"H>�8��fa��ר�@�\��t�r����7��kl:��w&�x\u�P'�'!$��ȉ��y߬�K7�s�9$ƍ�Q�>:��*Z�7���SI,{m�o8ȉ��~�
�j޾�^�R���������ڜ�k�P$�mu��W|����A����HY=�oE��=����C<����߀'đ��oդ��mO\8}]'T�U��8Ɏ��77�Gmox6�gpn�J�ty{9��ű��ص�f����o8 y�GVu��6�<�H\Q���5��n	�y�+���drc�BX �G؞p�Ή���5��7n9.ɓ�!q��9�b|؝ع��Ǯ;F;+cv)����'T�9W���ul�z��9�VNΑ�i�/n��FZM������(�;��Y�α�N5g�8���]����io��?���,n�m���m����ŐO����3�b�/�d��VU��ݷ멱�sPbI�R���(�eN���޵rf&�9۱�ga͓��_m���Kگ�(Cӂ�D��d�ܡOZ�*�N�_&��%�u����D�I����Qw$�#��X>$5}qD��z!C�dG�L�߹�P����Fb6(��D���Y$7��'#;�j���T��:�:�vo=�4�D̎ ��#���S�϶�$s3��L�%�"lvꩩ�#z������1d����U^A�+�4�Q2.{0c�wn��ٸ6������,ӣy.�ϣW�3�q���`�`��1>;��n�X��"y@I�3���t"��G]�J?m\� �����hXՠ%�$�D��3 ���yg��#���F���֞���HzuW��Ӿ��>7���xkjICW��smN�����PY�t��=���h��v���o�Ng��(�~﹭�hS�{Xʋ�o�9\�vJ޻�����d�����e
>$�6h�|a��JlM�*ޚo���������:���Ib)bՆR��}vTL��d� ��꾴	$��������^˜�gu�#<H79S��bI�(��絕@�[���:�s���:iNk�^�H�|݋���{���w{�܌X[dp�E����Gn�3��v㫻s�0�(6Jơ��ʈ���A�+��$�N�9������}�c�?�m�����MQCtꉤ"l�	Z&"TO�a���le���jM�ǳ�	!�mMA ��v,c*YY9S��2��A�fb`�����Zꏻu����&���b� q���'r��ٹf�1�vnna�=����� ��7��p-h���z�u$�ݦ��*������:�Һ�/��?Ց��jO�	#���Ϫla\��g�D��&��/ΕD�ZC��^$	u�N�뇵�:����u�-�#��'�KK����ϣɃ�=!zF����s�l�s�^�����F���s��Zgsw��V7�,���tr�G5�wn,��Di�"[F���ĝ�Yy�%���_��甆fA�(��ݵ���|I�����!�ي�F����m�1aW[����~�uqB#�LD�E�k�zDza�w���'�$kt�fx�KYjI �"+LK���}�*8����Q ՑO��� �{qD*"�M[в6�<	����|t�j,�{���,nYl�Fy���S���e���ļ�dvX��[��|�t�������H��S��z��M��t=t]J�^{��"�}�l��dLvc���^ƥ��Þ;�O�<�TT��9��d�59�*��xM|�WWԨi]�$�:�?~O�� �דٕ���>��X�ح�W�&�uQ��������������xxg����<;�f�9V���r��#&��aX\YB�-����mT�YS��=F�ݐI�O&��M��ųKh��B�v�/�.7��oX�Iչ�@���D(�(��5%'|��9�}�X��[O�='��WfB4o��� �ܭU��,��q�YY\�����$�I`#[�&�f9�Z^%f�U�U���{ox?/2+֑+���*,�JLL̨��V�d� Tz��
0]��H's:�X@�o�ޕ�s����v`^:o�(��+D�3 D��Ex*�^�{[v-J�U1P��6H��Q>/sf�y"V�8����8kj���Dcs۾�۰�:������y+8t\�tЭ�u�X$�#mU�n�t�́�e��[��4�u�a��U흞�M��@��T{3fLR�a ���t�Z���$��Z���"�\�%ۂ�-�:�6�f�M�[u��Y,�Sr�편�+��sn�k���l�t�r)G;n��=m��x2�nYc�{<�ݳL'=��N�*����;3��Nյ��Q���C���&�K��
K�lr��>�n��^�&��\����2t�|�[	��<�ZDNΐ�����Pl�{	g�PU�TP7UQ������͹zn�Ж��/�=w8�j�V[������ �]&�}���k��.Si�O��;�T
[�<��p(��ڠJ�uNEevJYS��wY�Zl���w���p�����;�A:�m���z�FE�D]��L��H���YU�|E��VInylmoE5���A#^:�>��?W��� ��7P��|,����2����� �=��I��w�CL�l�{�\_{F��1:
:\"fb'���O;��Ago#s��'<훶�S��)�A{/o֌���ճeu�|3���}�"�Q��E�N7�m���)��s��69��	�G.(�*�������S�U&&b8TvUI���/�o^H��7�`���Sj�$�|�ő60��bBI(���D[��c���p�Ⲯ���r�^��:n�4���I`Y�2%�������0��Iu퓑���3W��9UNv�+o ~ b�������wm��	;��׈���2zx�`��s݈9]��-An��`D���� 0g�J�<c���G�Ǜ�I ޾۾(��ɠ�sb"T������W\҃�ӳ��NZ9��wn�$�ɻZ���rv/�]H�S�$�݋""*�R�$Ɉ��z(��y�45@;��
'f�)��>'���� ����!�ꩾ�+nv�iB(�Z��v�����4<W8�s���#�[��x��ʬd��P.�]E�K���gw�֚M��PI'ݙ�D�(dIp��#������*`8��
ŃV�9�Rݏg��H�=�.{ܠ��[��ω� �y>���DE+2&��'�������LL��S17��w��w���Gl ��>������j�_dOBΝw�6t��J<��@.-UQc��3�φ��P�~�{q@�4|��i�TU�Oy���w��'F�q9�U����g��׃W���L̓΋n-�J=I��{x����x�QV�i�U>���A�*YK�R�a�k���	��"=�<�zzt�S��F9�����vҬ[6��xX]�DZ0��Z)���]�Y��e�-Aͤ��!�B���pjk/�s܍�P�p���ܦ�� �y6fR|���"Þ�g��SOT�ħ�������+Y����,�_��Y۲z��z�o��-��=���e�Ivځ���{|��G}y��Wntl˥��GE�|fT,W]2�N)�E��䙬.i�j+5K���]10w?x��ñ�XW(�gn��:b`�t��Ҥ=Z�
D+�6N<2+!���}�/Y|������g5���W��Q�s�z���5�c�s:�#֋�A�œ%�<��r��R/���,V`;̥���.)�f��C�CQ��2�=��f��)�gsq"���hf�V���*,����Ww�ɭ��E'���#)�b&:��!Ul4q�4-�=�95��Wo��6�4O�@2�^7��v	T��PTʋ�7L���m@w�vo!a���n���*6�2���U�[�E
�PV[�#1��zn>�6a��]�C�t���ޥ�ʍn�xTc�1{q�٬�������l0UF�mm����SF^@��//�r�*"����J�v�I�z��}��_8ܪ�����ޤܢ�vLV���50U��USw�Gv~����/�jZG������<�9�O��$׶���Y0��;��y�}[�׻ĨLW�Fz�Z�����E=T�L{K�5�2#	 ������B���eK�zV�eH�N[�V�树�1��I�n��Re������
/��$��DRHfh%Q垑I��G�#<{J��t������c�I��B"L<��$�Ct�u
0�"(*�*�ʪ��G�o߽�C���M11�3(�<��(�S"�"/Ұ�]��C3Уմ:������yaF�cd%E�d������E^AVL�3#]]������y^T��3"���gD�Z�鈴U#"%5R�C�}�w�H?��h	���P$m���T��*t4�����P��:V����^O�箬O��������a���5�(��B@��S@�]�Y�.D�!3��u�@��F�߮]�Ö|d�$�nh�/s��$������	�eZW��sʂ�E��vnAC�l�ѩB��{zun��i���]V��5�0
��L�� �X拓M�9�I}{}����c�����<;V�����O�٧<��U[��+�;�_��A�/�I���;�[>�ơ�$H11!A����Q���I�olX&q	���10�L���8�{=��
~��8�"I%-R2{6�Yɗ�|1N����J�s@�5cs�`��d��*�;�yc$;B:�v^���f %�q}�OL��^�ә�d�6_o9 ���l�f���piT�9�.�U~��}����:���*LLLLH2������{���A�;��p�"�w:�7�|7��~%�d��}1�VS��V�L�	�oc�N�>.�Ij`��;�s�⻲�,j�Li*f���dȐ�����:����b�D㽙4]i(7"�*]�E"!�� ���j �t1A}n��E�A�!C�S�3@�I��u~$�_fHg�� �(�fQL%���L�D��Ny݃��P|D���lY��]sgD��lX �ٓ@��1�A�R�2���9��t���	�����ޟ8?^�Dվ����NgF�h�b.�ř�bւ�(�JZ�g�c ���X�y�~�Z�� �UWA ��4I"����:w.��L!�� ��<����o�O��v����8ȡr3�Mr4�x����]��r��@��E����H��ӌ�}3�m�T��u?�E�7SQP��{^�kg��nz1mE�62U��ءv�	���MP����e܂���9�jwn���s��`;:y�e�i�.���p:�²����{^:N]��^�a�r6���Ɯ=G��&V�Mv=qz�&l-�x�<��c�9��kNq�����&�����}��9�[��Am^��wV��pٖ[k�|N���*�f���i���j�&FSB�<�6�>"�d�������O'�'�hI[����E��,���z�޵�?���/��r���xξڠu����Y���b�|u�Mj�W��
D�L��oeP"�B
]8ܜ��V	�)�O���U��)ܻ���&t�V�y� �"$~TRV��k��2���s{�����	;�\�z��$���f��}�^'�SX���hS3>;�4�F䠅��Ă�V�ٟA��B�'��kj.8n0�i�#����U����&&$�;]8H ��������e�ِ�N]��	z� ����3�s��j�w�M�C�����2�9#Vک��MڞGz��Q���/yj���R�{X�����w��Uq@��&� ��u~3�ui�ׯ:�Ӥ�6���u�q&TDLLLH2L�&��8l0ϧ�������Z9�PG�Λ��,Z��I鲬&����s��ŷ���޸pb}֬a.�\8s�F҇[�q&a��g#2�)��{�c\w0� m�'�O���X'�S������s~�ͻDGL"B&g.:�m��1��!%�*�e+O�f#>��ij�U�H������
 �"$���Q���*���$n/��<������@�]�H#Tt^�I�MuQ=3M�13>:'�{��Hw�@Ti�ҳ�4n몁���$��[�&Pۗ�{��׽���i������;I+�Zy���P��㶰�AB����El�Ys���1�I��*{��P�7u���veX=O����3�@����J���AL�E%3L�d�"/W�"lօǌ_�5�E�A$�o;��}sT�ile]��e�?+���]$�[eT���v�k��Y�ZM���1���J�cF^`\���Y��Q�%�F͘�I���p6glS��S�9ѕx�]�N�8���R�!�m"!H&n�nnǘ�(ج�����Đ���U�7�w_n�7���jv�UP���\��Ծ���x�?��d�`}1< �ﺟi�gs�"r���� DAbP���6��^t�S4�1T���FN�]�n�P����
�u��2���j�f+��5W, i�����Oo�<����]��ϣW���%��/�у^ǭ-����s>�Z$��ר��r����[F�d�A����@.�� {
7��LLIRv�p
���Q�mꩪ��_\�$��P�vb����_fg�}9��)3$��boǮ�>.�٢|}5jr��4���~��< ����2Ozj��Ԗ�E=׵*��3@ufUH7ٴ(�������֏�f+�퐷�i��{�����V�;ԀkX��'��3:S06kl0.�&L�"�V6��n���y~�]���V[Q�*D�L͕E����Q��G�;��O>D>ڪ%7�఺������ˀZs&y�g�k:��ݟA\z��v#�d�=C�el��/:�b����5浞�9i�s1ȯH���Bj`m�1��[5Rt�׉'wQ���J��T�L����u;AO��sE��#��U�@ �{
��=�~'l*��h�s�/�^���ۖVZ{w�������֛E��ܷ�=t�g����W����,a[�	 IKT�0����[F����GI�#�{w�
��ɾ*�loFN�c��!츪�<*�+��
&&f&J&��;�8����ݧ1�e�����ۿ��4_H��ԅL���^u�3D٨Y�-ʈ:sic�У��)7�h�"S}�{k����Ϟ\\�_v��#{�q��9˘�j�%�l�m�$�[��^-;���<�]le�'Nt�h�;c�ƆU-0����ln�<��i�a�����c��#��n�\x�p�н���d�s�
7X�ѡi�.�\l��#����5�Сz����&#�%r�Z�k���m%�F�����^x��f宅�ķ��y��a�a�+���i�V�iwh�䶜]��Q=�ԝU�����Ez9ȋө�^��_.:bNݎ�����io�__J��a�P13/��U@$�{W� v����8ܧ63�����j!*�b`DI=��&tr�Q���7�Z@���m��'o�k�PK[Uq�EH3ոH��@�x��b$���]������d�����3�QRk�@#��ۻ+��[;-S�1�(ĐbT�6C�Q}F�g,rXt27���'n����X���k���̻Sa�܂�2JJf&Ť�#I=���_bS�r��h�U�~ �g]`����֎��ٹ���+�9b:XR�u�����8��r5���{I�f�i�R�zY"�ۮ��mr9e���=NkY��5�jR�H�ΪsU��:V�Ei`���A>^�Q"��t@p��3��V��R[^�f�~��H�Y%�]ojL��.�+�]6v��k�o�`�RS躻0�mUCIɔ	�"g-��I�fm<0�g+����9�	�o:E M!է�z��{\־�1j���IZ"����~�Ff}4����tFթ|�3�`���@�}�U@�5�r� ���� րk��@Б��uB����T �[��7Q�A]�����D��O ������#P���U���=d ;[���#�,��h�ߨ�A;ٵD�}�`�8}�}�{!,4N��RKR��t=�� �{u>�;�1v��i�bI�L�ҫa/����D�RS17�ws���l׉$���ߏy%w��Y�o�֮]�zT�W��A�""&Aq�v,��#{`��Q$���h���݃�2�3�4��-7<[��֍9�sJX��;θ& ��0~g��ቦ���&�˹�5^C����hՀG�A����x?3�q��ER���`tU��>��b�{�>ٳ*��5v��e�ea˄�og�>�9�Io{nτ̉*��10"$�,��gTA���I�7mX ��əǂ)t8��t����\Iӱ:L�D�k0�U:��{�Y!N�����!|ߡ ~�>���:}SڃO�� �3��ϳX��cm��y�v�"3�#����C�h����ѨU%Q[/u�z�9Zr���������g�}�G]�oC��Iz��T) E��bȪ��>B L������#wk�<w��yʽ�$%,�����y��`����3��R����n���f�bff%h�w~�O���P�Hgk�o�i[I��w`�N�d�I�Mp!J�p$����Gܹ�>6��� *��`O_rb7��go����oǽ���;�J��@�N�?T�LM�*Y��/�Y���#b���3=
1�g2b�;/6)��k�U�β�ڌ>�ᚯ�I�O7:L���Z�D���hṽ��7d���n�	 v�&���C\�s�9��n�=g(�!QJmQJ����t=�p�덒�Ug�+!��r�-ӆ�}oϱ��LDD�ox��;ϥy��z��>��<�eŚ�p�Ń�A�ܚ"m�L@�bH1*J�o���sS ��I��_|��/y�x���G�6b%՝߮����|�Ɲ�!D)E3�	�PA }�(�VX�������$j�ȯr@�i��3ޫ5h%$� ���d�u׾�{zٷ�8��I ���P6G'��|s��^.�+�VS����'m�䮝$m�x���kM��r�*��@�m�x���o�^ ���y)�EJR�pn�7*��L���q�������ވ�s�?�,��+��q�=���\<�9n�)�U�
>
p��=5;�H����	��n�p�N����Őfr�n��ջ�p�r� �{c�^Wv��԰>�{v#Lᩄ�Q3FĹ��F�҅g�4�5�D�v��̃Ҧ�Fj��'�>Bf���˃dN�h�2�黳�][�n��Y��=v,�*�n<(�l@��-���M;��F�U���^Scsd�2�M�v��<Eny���L"�ul�=��Qu᜿v�*>��� ���w�����[�y�kס�QjWn��w��v�٧Ζ�0w���3�YG�ʈl��R�=Qu���*`MLUf���i▲Z�ѵ�Eb�\�!m�x0w�q��RC��態���"p�Z��o��"2�������w��4o$SuZ�	�9�B���6�R��x��'9;��y�yN�w]ў���{�۰G�Y��>XY�\5�󹥌��F�S�~���f[��I0�5�,��)D~������&�{�}��V�y�Ob��{o`j1(jfJ�llT(M���6rJt.Ħ"�ln���j5�����:�{\��3�[�J��|ud��l;�a�Q��wZ�y��un5#qxgnb��-��b�܃u�p���{�Zǹ�=٨�ۻ��'W�5v�(hXr6�u~YoJw��7�'��ߦ7���63��дS��V�N�ރ�N>���_\�ovF^���!Qǭ��]�oV��
(v���e%�^����n��b�coi�v#��]u�>[h�����H���hloL���"�I<��2l�3�![k\j�nG�Ʒ���ޡB��i�dA�jG�f�V�UTV�M�Aq-Q���YUt3�p�e'�e^�x^_�`����&�D�|����$"�Ho�{�oRCKS4�*}�3t+�
��#�0(��b ����FK�!>���<���(���Ve�X̷A���="��򧞸u����～�$�K��F�$������+R�x��˩�JSTB��߾�yTO}Y)��l����Q+��e��nA�Ѵ�LU�"�B�7�QuM�o}�ޡ��A��6�Af���0* ���hEQ�7\�/�/���}3I#(���R��*��ʋr4��7t Ќ�T�\�R��BRsʢȢ��DL�-ʱH�K����9b��G0��n�P��<&�xYݜcp��>�T�K���ݱ���<��=���u�F\�dS�|1x��6'i*�뗵����V��\��!��v��chŻc��7)�j\z�m{+�׹�Sr�����]�m�7�ՎP��8و�g���즻OF�d'�鱴�K�݌jvm�K� oP�y;D�����Q	d�j�nT\�.ٚ��W-�N�u�&;�Ʒ:��d��F��繷I�2; C����ʶTѻ�Ίe�콳���Z`v�������c�R)h�&N}��Y+�w9��78"�������=I<tόy�^���pa{
�jL\NnzK-���G<�2vL�۩���j�<� w(��#��	Ĩ�ƚȸ�=���=Ds�q�$sΛ˸���]��Ɏ��{iӸ�Ϲ�X�n���<l�Oj�����q";3���+�m.�qթ���Vx�e�\i�&�D���sc���';k�zSb8��0,�=��c��n�_n;]�����g�qݮ-�۰��]��[K#t1�:��d����]��q�����[����tv!�M<��FpGuý�糳Dݢ0�w�w���<���=�cd8w0�z��F�ıͩR<���5�Ϻ�K�{R,��K���"���m��/	�\��V[�axn�ۮ��r��q���vҦ�74�g�].�ݛ�糲q��d+��Cv���qX��`�:��!�R��ka�Ơ�v�ֺ�a�[:sr[��r���;;Ƨ2�S���&�Ԝ��">����ہ��شF��ibN�N�`:,��s��.�n���b۟)���V8�t{G�c��k���(�*/1��.tޚ[hE��#�h�\�nv=��<:���m����V��t�v��Fݳ��r����
'WG�;5��1��m�.\���8�)�2nܽq�3�s��鶙J��i���ql��8u�zčy��٠�Mur�k��1�OK�)�-�[u���Ľ��^L�q�77k�y���-�]�v�]����;���C�vUEh����+���Eq�z�;�7v����c�E ���Vi�Jûk��B�������m�uј�����������'VG&���ѐ�mjń�x���Uv�45�X5�x�-��ɱ2X�ڜqю���'h!�kómEܥ[V�셰��L6���=��[uOd��i���[l��Z>�b�v)+~6kz��F[�	��U�RjNA5���g�����~dC���%`��*��b���a][3P�~��/�7]� 	���@����X&/զ.⻶a��g9��F$���;s���;�E�.�]��JV�8Ԕ*�� ���b�iO�J&!"�bs
/0��|�#�� ���@vv;�CU��՘b;�����7�~[��ƭ��j ��+&A� Y�ʓ԰�����&1�P$y�;�I�U��Ơ����͹�������g��vm�<�̼mu�-C���������7�_ikV�:�s��z)e@����}�r�&��@'�����\�{��8�����^��ő�f����AɈA���$�}\�FD��~��́Q7��h����7�-�����K�r/n����1.�:�'��X�Wю�E̍\�Tj���X���#s�ᛇ�#�O����(vkٙjw��L�P�{3����T+��&""H6'����If�"�TH��N��kQ{,|I�ol�}�%���(9Zq����CUu�=^���哱�mnnX ��vG��u-$�A�/u��w/���44��
�FS17e�B}��hޟh�$D��$���4�f�W����\����(�w�ѩj�I,uLqu��㵞�yLNb8�1h�j_U���%o����2,'PE" ���ɀx_W�`������M#�߰MfU+�������6�{�Sff�}=�^$��a^X��4j(D_f�z�$���&� ���}�8�y��_M�/W��$2n�O��9�$����@$��M	�f�K�?��}_��>��T,�������ժs$���3V�����cu�P��жf�MCx\�&s���J�[Bb{����Ț�u5�����D��U���t��"�.�$���q��}��]�Y^� �0O���TA$��Uk��ű�ۛ�ݸҬ�ӫ8ɝx�����+B�:�T	� �s���ا�u�@��h�����~����׬z��~w�\�z�Ge�n�ܮ��v�MȽm�6���8y�ζM:��V���t�D�G �]a�Z�k���I^�U��̎|��ujq�>H<}U����LJ*$D�}��g������آ	���*;z�_��!injy��ӓĀ��[!LHH��q�;�y���HJk��i�[w6	$.�۲Hǽ�q��%(q	RA�a�f�+�I�ޚ�$m�]����tvҬ�!z�'�z��!ڣR�$$d֘��0��	��-"��l�G�����Y��
x�9S�Y�q��q�E��I�ݚ$��y@����_���b�$���K���*�{=�(�1�B�����;ۓ@�7�y�R@�,D�R�E��(7����s^	-ŵ�=g��.�Og�n�g�{����`̥=Nv���u�m��$��rh�o���֦�oQ$����B��{�H�IKS����:��g)3z�=��ɢ@$4�t��~'�܊͆e�$��>��
EdI3*&&F)^���zר)��w�������/�/���� �s�yb�'ܞ�Q"�RA�Ą���}/(�L	��x� ��ɀg��w�ߕ�i� ��}�8	���v]�J���RA,����/e�9y�8FC��B�>����	>kw"����ŕh0�r�D��zs�� �}7�^gK����+��x�bTo��H��+^؃s�ϛ��f�hoI{����k:E^��p���pp�$��u�u��v�;�*X��rg��Fގ����k�\V�i��v��ڝ���sȫ�5�v��<��xo9�Fպ�;q6ci-r)���st>��q/���r�f�:�n���ۨ��n�3�v��LX���G.�pt;���v��N��.�/INB�>���Qy��Ȇ�"�R���|���z�b��Dvz�ۙ���j+4�⠣�����-�d�j���������K���ٶ�=���L���,�ߑ�qO)$�=����ii���*H$՝T����+�h,�wv	�ې+�0��e)�+'�� ��=�mu1�$��1g���;�����gMx�
���jc�}�\�Ϊ���
eIL��xه���S٠H$�=8Q�5Wu�x:��~"�׿U�Վ�x���AZ ���nRMW� �u$�C��(v�\�_U�=$���zn0�$��aZ��	$�r�o���t�F��UJZ���٬2F}o���y�]���u��
DL�RIl����-<<��I���c�絞��l�I��۩��/;�rFyѨV�8���V���v�Nv�U�h\voNR�ȠAOj�HSa3b""H7`��v,�л��Q'�����7��YIw���>��xkz��Y�>5��[��ϣ�s̚�%��6�J�?�r�V�
�v��'j2�n�݊�	���H%��I';{n�}�9�s|��ok�I�u�
�HFe)��8O��ol ��8(�7�����Z�+khu�"v7�Őv�ڣ�
d$H��{fƈ>�p�<.㛿d``ݵ� ߉��w`��D]�jD��A#�����<�l#��V� ?|�������v����B��O�{�߬y[ȠV�N��\�����i\ʘo3t���F8�p�C3��ny|�tAc�:����D�K�t�4Z�Ӷ��e��m&�׷�ņ�坰D��D�d�̵^�ͪ ���{�Zh�F`�F�Zk8k�>�k�׶4v:5q�`�����$����|I�y"���A�E��.�ċɦp �� �Y�Y� ���:/N���^ɋ��e��C�r谝��N�;�a�S���~dݱ�2I�x���z��p��H��d�n�X�s�&��4�O�7�w�z�D�$Â9=!���l�*�P��5����~$��vMH�Ψ�j�73!�0�F�ú�H�c_���؟�șL��S�3�#��Е�����B���ϯ:�����Mx�76��zkZ�v���~ġ�����뜫������k�����a�4�b�Y,"��ͭ�u��u6���s�Y>��I"	y]T��̗{�R7A��w~%���9uI �
d����>��F�����e�-.�٠RD^gP�����z���D �J9J"�l߈w�^A&�:k��aK�����ʋ7s\����{>�ۛB�Qa�
������O�J�<'�nn��R[�AV{�C�9��]�y{Sծ+v>��)��i���&�Q���Z��f�+����:�ֱ0��X��ӄ6����6�Ѱ�:޼������~1�&�)�2zB3)M���l���mu����>73����Ms��
��{���yV�{t޻j��\�V�e��m���᭻ss�ӈܐD+$N�o!��Ul��iy�z�bL�*eN�s+�A �fȠ	����Һ���r�t�ӥ4I>��TO�U���5`Z ����2h�q��W�*s�A$�Ϊ �	<���3�u�>���U_Nrn�C���L���YT	'��{jaX=�����]�m�қ��^�'w�/��������� ��	�F�H"���ƅH3�bh�2��Y@���łI�.�cZ
�1$9Ƀ���}w�~%G�J�"H7`Ӟv,�w�B��D��� �n��:�t�вN�d��xN�ї3�t�9]u��pm�p�ܳ�k(f^�[Gco�Uct�^�}�N�>�r�V����D�n;a��f�j>5�n.��[\	p� k;u�=9�EH;���k@����9��a��!���h{	�a���]�р��F���A{zst*���;yqi�'���ϲZ<��텃X�fN�?��Z����Bj'�v+�}�ۓ� ��c������r�7:*�i��g��p�P9ۓ.-č�=uIhNNp����;A����犵�5DO��!PK��d�)v9�����na}u��g��K�;
��+e�<���u8�c�/�;�z`;��s>���]���wT��TH����`������I�bL��2kƨ�������yS��I=�����d�$�T�����MՇ�r�$D��e[���;z�5q�O��Md� �{��'��vMWTR��XW�N���Դ|I��q��f@I�;��+ļ��I�H�����LKǖ@ʚ�AH��$B���E��:2�>��]*���v^`�Ix�EC�}a{�#V#�Ur!L�PdF]�Iqn�� H�-����5E�d:�"�b���~��+�J9��n�i�9�+	�w��+��j2n�e)ύq�����{�2�p
��:�lv�s��^w�=�%3�^�ECQS�T��w"�GH���8�\��>��l�r���4!郣8Ծ���k�ꝗ�����FFC;{�VK�Ʒ]��z�/���9�刑A$�1�`�I�7��C����40�9(D��*$�ա(W�$��\�r� %�;��nmYV0��x�#�dM�����l�����[*zbIȼ<�m>�ִ(Ԑ�B�ȡH����>�{ ���R^n> ��~y�Y�xԕ���~�}��|�a��}��S̀���#l�7�BI'��w��nX�돚�j4} 6�J����Q;��������]��!� h�ڵ��$��L��5������e�<����i���ss*�� J�;�$�ISڮ�[��vA�;���]	��A%���$�l���L�A��q�qi+|wEd�n3!�I$�nofbK�/'Sڨ�	(�ݡ���~x�:����@�1�}���y���ZI%~��f��qE�OX����{�,)+7ڕrU�œ���8wx��L*oo|��ǾY�����)}�2��1�c�;���<^^��v�;�mj��J���L/o���&(��C���
0�>h��"��nh�Og2��*�V��}��g��������#�v���{W{H�����b��G��V�S��Έ`�ٙ�\�6�m
�[y	fU��&Q����y��z���ј�ʼ㵮���#v(�e=�CJ8H�ĵ{[uC��fD��QQ����r�܏� ��R>B67�B�������<sL�®'ǵkone�ԮG��O.�nL`��"7�8�wF-���:[ZO��=�wf�_�@�>����H��{�O$/?(�85:�.���s�z*�)]і���gmԱ,ֳ�ҙ�˷'le%��i��ɧ�T��Dk�o�-�L5v���ݰ�������VXx��lD���0�|��LZ�Î��R�E��Lg��y,��٨M�������o-��U�ux�q|��^�����Ѭ��/l#$�&��ӗx&��P;�	���cN��:h�r��P��9�G������^,:%ZuE��pS ��ވ����)g��6��n̹��uC�]�����<��L��,|=@�z������St��x���xx��摧;6d|w�\�^Թ��Ɇ%�1N�h[Q�}��{Wo����ڻX�F����~�޾ c(�h�f.�����5������TK�2K�Kn�09Pk"�N�f�ģ�HI�'Ʋ�4�D�_�s�%W��J�y��E$~��M�[m��?R)��T�����-J�0Ƴ	P�*��Wl�H�y�!�E9�����<����ތ�B�<�>v��yiA�>L>I���<����Q{I2l�/V4i_[{�{�T<�T7<�T
<�6�^W=�@�*I2�1S3~�"�k�^A�)�*��o~��<~s�ī�Q��b������6��L��2Z�jS�D��/<��2����{{���y���Q*�C�'OI	2/��4�L�\�fixg��FAU��M[�z�D�����B	<�!(��ʽLg����'�O�xEMJ
*�����
�����!�zj釉T���W����G�7��A{� k���{zV�9T�*yA������lB<.�U�ʧ5D��C2��I�Ԣ�=ś��zU�Fr*"�*�UrE7+^���a��&jEQ�2!c�H�K��}
Iu��Q��C��5�AG?�����v���K��ȏI�yט�I :��]�%䗎�P�k0kbv�$zj����h�ѐ`�"��� �s�I9��ǌ���_r~|��$�����A$��Wh������x�V�(����MC4��r��k��j�N�$��\C��;&���mûHk�Lj�g{��q�ö��{浽��Gj�I���@%���%"�]v�{[��p˶֌�7U�+O�|�u
���U牚�4�n]ݞI%���/�%���^I%6赿<��t�wul.jcfT�������s=�aM a �dU"RZj�'wc�JJ�v��+��=���� 0��eV���'�R��P1�1w�^Aܼٞ>X�ڙ'	���$����^I${3��E�eVD���}RJ�*�ӓ���k᱾�ﻵ}�RpdH������j������'�,����:zJ�C U�4{�$�N��3�>� sR+�
�9��T���Lt滲��;���\��D���'�s*��0��=���Ρ9v��Tm����IJ71 ��Ɇ)P��n�S7k�d�91h�[!I/6�vxq�Tn���
^<�a($!��"a(y�ل�#�7i�oB������BHJ�v&�HUVނr��e���ֵ�l k�5�kz]�6�eɝk�] `>��W(0���}` G~����_���r��C��8pB&	�) ��3��R^I%y�׃	/$�>k,b�]1����:���H��=�e��V8%B� ������c�.��Iqۺ$�'�vNy#�{b�7 ԃs�����4P⸖�AR��v�V�fbI$���&��{�&�Z��� ��}��$v'�.���~w��ͦt��i�j���};��F9���n'�@�@Ҷe��w��u���8�8�w%4�$@7�X�*F���%���� �����^ֹw"u�n}Za'�hu���.]���[O���,J���s�nT͞68�gf�f[����Mn�]'k�8r`�ۊ����E�6�;n���N�x4x��W9�6�;�oC;;��Ў���l$N�ǯ,W8�>���k8�a�Z�^�=�3�wnl�ks���n��a�5G�ݲ�=�[��Վy�P�����#��3��h��m��]X�:.�*�mŽh���t��ֺ�闝�^��R��%sZ�ཞeg {��=�$�A����Gb%m�u�v�`6�	�%'��3��H�2H�"DZ	�e��'�,�o�~��b�Y1��������>�ܚЙ�]������ �⿰���	�}��V/�jF��\�`�榀7s�[����Aw[y��I�{U���%`�H�䤂+�A���= ���=�$�Wf^��m�7��=�w{2t�C�[갓���T� �x7��P��B~q��ZI���&\Nd�6'&N�z�>{��8�I:�j�@��IkZ]�^�.O{Q>-"Y
�w(�[+�E�e������;���7H�=���Q�?_{o���6�DVWr��գe�K�:�XU�HP�J��ϨE:0y�N�����sUڞ45���-%RW5��.��edo��Ӕ��D�ʃ{��d���R�����v[�0u܎����Ӳ�u��M����� %vgi�D�eڻ�K�}� j��S��jf�w}��釪�� ���I ��Y��ah�5����{���(
��������Љ��U�� &�X����;�x��zk{R^I-�z�Z)'|� ���{w�_�Ԍ��׼DÅAU^�D���"gH�J�!.�}�C��(�H�5j�/D�*�"Dh�%$s}BM$M�>��(:{�l˽��	!y7��$�D@s�M�	}��}�1X����6%F�g�B�3���z��ۗ�ڈ��]2A�����<vK�ț�]^��Ikr˿q�G���!+Mo��g=��r!�*�%�1�{��{�wz1����)!��&�B�%dt�2��=�}>��!C~����~�t؀`���M�K�9哉m7�
0�g5Ӻ�wX��b���+��GuU{@O<n��H�:��dGT��U�׼ǁ�iy�Xݽ�-kh��JEc쉥e=�;�v*(�e�m�6+f���I/Ρ$גAvc쳗���L�H�$E�JثZ�ɾ�{},�Oծ�O�r(��'	 �K{�@�I>k�3(��巡�O�}k����j�3�12aqUw�ĂI'Q�b-�=�uոE$��H�	//з���q�T}�ū��mP���~8"LJ!D�0gBGK��uU�d����bz�w�XC^���~���"8O���C/hI��&�;��8���WiXV�Y�v�"{�\xDݾ��%�tQH�Na
$�3<���Io���7V���8�E�N�ϻ_<��	 �)�Nb���Έ����9ق�X��WGI�!1%e`W/{3$Ë����J��M�Ҿ��؎	���y۰W�AtelX��q���LA�K��vG��ym�n^��CI�
}yy���e :d]���A����uW9MX`\��tx�y_?����T?fDc4���G�D53CI�1��=�x�6���c���#w��	����=��f]�<k���K��]dȔ�UL��s����w곓=ݡ�&����H^}���I$�迶,Z$�Ϥ\��y�h��ȼ�|��m������Ƹ�9���z�V�c�3�16}�n�}st�7�����i|b&S�,ڼ�8'�����D�w=�rFz��/�S;D�緽����ŋHL�lB$�&|��E���
H$f��̘�9�����MLH��زl�:��<'�w�c�w�\��9�^���,c3 �!+Me�3��M���H�A%��5�P��6��;��H��׹5�	��~ʹԓ���a�yZ1V֫��Ξ땑�6z$���=��I7���H.��)V����x��Ok�/O����)i,�gB��VR�`�E��{[٪�qy�<����%��I$�y�	�$��]��f#SE���,�'�Ƌ*��%��12C��c�u��{�+���ի,�H��~'�oW{�����rȤ�ö#Z�רM�9�"#uC`-jgM�\]��N��I�"h��S��i�k�C�۫1���.�����m����gWt#�o؝���9^����v��,��n7�es��.Ny{;���.�Y�%pv��۰�c6mqv�rV���{�cqe�i��%�m�6M�v�XB͐M/i�ڶ�I�r�4e�t�1^�c23O�v�!��Kۄ͵c�jՕ�T�K���w�)�v��:W�b�b*n׍u��:6��GZ�6ezj����>�6�UU��s[�А6�ߪ�2 "?���=��OM�:�\Q)&.��V���X��9-5�{�����.�t��.ʹ�J�H�u	�	$��0b)%Ox�i�pu�oTQ�3�)?ۇ+O-s=��܊w� !=l�g�ݢy���k}=r$�Iy�wzvF2��9	Zk<A��vzCݤE�.:��"�$�	,�o3%�{Q�N��1	 i�	'H�%'��(��*髜��ĂH]Cۋ��DO-�4�6ˡ5�E���0dIvkܚ����ϟT{)�8ӓu2����R�ܱ�k�ŷ-m�-�A>�C���S���\%ԭ������*���(o-�^��C��w�����N+�.�M���Sʨ�5�H,��g�$+<�Y(B!@�"iX	B��
���wb���Ë6�X�ֱ���Qd[W�HGb���y��1�h������4���{7z�燲���]^s�0�U��4���I�!7\��$�	�vE�Ey)V��h1w�\��Jj���"$J3�2��:���D�]�V�	M	���{��D�I%���b)$�Wdkn5���r��weN�9U>���O�x1J+�.�^I�x�%ߗ�ND�����DX�/G�RF!D�EX��W� �%$9IA��S��ne/����|��jE�^�ֆ �����s��KkdEY=�F�T�0�$;����'�y\Q���5l�w\ލ%�s�ߟ����L�P����+����JI�y`$^�~x�4}�����~w�� �Qɟnih�m���Y-��g��4�RI7yw�;�!��ļ�+�+�.�� Hڡ5�V�M�b�]Ӹ�bC;�Oe�D2*��4�3�0��Y�$�Jϯ���Y��o ���V��[�N�_�@y�k,�K`�Y]U�+:���߂}���������F����ʱ.�>	/$��SآI�s9�d���h߷5b!~�p�����:��z�D�DB�&גI s6�גA%���Ahs+�D
�'ƿ�0ŷ�[�f�b�V����{*��0���*�70g�_Z��+q�X! w]	���I7��tU��I�e�ktv��
<���etU�MJ��ŉT�z)涮'��Z2RUc%]������	Zk��b����I$76ERI C���bO�e#
��GvN��I�o�$��ps#��%�*���y�q����72r�%WQXA$gP�I�����@	��E���[�}��CG\#�Y���Љ��#~�2p����{��� �hx���H$/:D�M��bC�:{-�UU��^h̷>�<@ �s�h�W���0��BAD}{�ׅ�0�[/�P��F���t��tR�fh�x>�*a�H�4v�����A�4�۾������+=��ڄ����8�~o���*� 1n�:�TwKMi���O�I>?N�-�8}�}9,ӓ���PRF3�n���k�ŋV�gu֞�.�qhhS����iFZ�u�!��۫t�՝��HZKq��cDuEm,�����ew�7�Vu
��D�>��D����~JV>���x-��@��K��ލ��J&&T��K_\�<_\Fe��do\BD��ݹ�A y;qb�A+���b��M�xRLP�%e��l,��D��nm$��ˢ����-+K���n�$�_VC܈���^J�(�Љ�g�Y���~�=��������f=;�Mh@�~�2�W|�S�&Ԏ\I���٘�=y�N�BP$H���%*�w=X�IޑT�p��s�)������f��g���F ��� {�?���o���D$O���BO��$ ���Ĩ�u������ 2�% � ���$@I �J$� @a�	"H��� !   � I  � �	 �	$�  I  �� @ � �  	 D@P D@P@P@DAQ ���$��n��/(��$��� I"��_�����?�:>�h�ߴ��5���$O�9����/�W�@$$�?$D��A��`?�p���a���g���?_���	 �����������͙���������������������+��* HI��?�Y�$?��BBXf��J�������@		?V�J'�~����	��S��u�o�����?�?�����?h	&�I_������ �Q�x�������4?�O��ş�	 ���+��~����~�e�	 �~�$O���n ��AޖD����d�	"2d���`+��l�j��Z��K'�c�6d�F �I�~���~��	 ����nO������������??���
����?����!_岿����BI�'�O���?G�O��?�� �T��?����w�Y��Q�?Ǝ�:j������n!B��������~�῾@!$���e~��0������D�_�������ʏ���d��O�@$$���?���g����$�!�FI �3��?�d��������?y��~ə���
�2�� �@ ��������>���� C�Ӱ=��D�� �
�9�L�����a0CLM0�'�a$ �    *~�@��   �  ��H�=M&��M  5 9�L�����a0CLM0
� ��h4SO
e3Si=M�!�zzSk�Q�Y�$j�KH0�F�"��{Y�ct�+��o�?h�1��a#�q��*�U�0!QiPؑ��A��.TL"���0�2�v��k~�w��a�ŕ�����BI$�I$�I$�I=`�tCkf�l+܎�v2�(*]������t��@�CI���r��;��K�Z]�n��-WH�v�y�!-_��ar]l9��i��,E�Du�b��Z�`�:t��72�3�����5-=���V�Um�$%��h���$$k��ɡ�Nk��kU3fk$��I$�I& H� 
��QW

AA��N�Ab��d�]%2�M�5�_���w��m6�4�����[&g;z�YnI#X������f-]р���0B���m'��vy�f���=/�ݽ�9��L�U��s,������b��!�Z²�iY������H	F�=�5�Ŭ52����xy�fT/1���Q�WP%�vH��\-�Q)�VIiz¬
�΀�^QDz�@q���zƲƨ�H����" Ĩ��W+V�F��s`������2�ɥֶѭٳ,�!>#�x����23�ƛM�6!8wzy�v���������e�Kݒ���^B
��>b���Mu�ڤ����V�`��)6�n��D�$H�4&�_��n��1�8��J#���\�v�
¬�Vt�eo���ז����)���Y겔�)1��1c��^Q�\���U�#��(2CU	3����]hvj6�c,ok�|I��d��jz$��}�g�*Ma9��U!TY.v'G�Xw�t��~��<	u?m�2�����\g��fq49I'_�G�?�����,�r�*P�'}H���D�&|���J���%��0�E�����v��C�u� uO�����t�]�]o�jr<�,�.�֖0�>�w��6"�CL@l��!�QF&�i��k�����.��CM���[��11T���)P���i�L��t&S�H��ڢ�����G9�F�o���}���YO8��S��|����m�,#�(V��9ބ�O�?bvuH�ϿH`����.yf��vK{:�3�8��O�c�vݐ�7��G�����3�q!��A�IE]�ǂQG����MsY��Ox��s%����QR�q�x'�"��/uD�KJ�#�\`���4�I���łh�CКZI��v6�hh{�JQK�7w�	��Iw�t�p+X���iA1�V(��D�^FYK�)/E���3�j�*��U�4��e������Ly�w%��C�P(�vjI�R]�:�w���t�'�&��?#GA.ˑ�S%~n�1D��wM}^G�Ig�7Ƕ��/��ޛ#��n$h��%Q��ND8'�=�Y�=G��w�����M$M��=ٓFrgFAI���R��Ƚp��<#�	�ɨ��ȴ]���Zȡ]`��N���ИE�F�4h�`in��*N����6P��؆0ʆ:�:t."��Odq�N��tp�}IQ<��h��8m�&['^�4��K�&CY���d��ȴ�2��P��GdUJQRG\P����[��?�w$S�	<�Ѡ