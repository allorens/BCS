BZh91AY&SY�9��_�`qc���b� ����b�    `                                       |��a�(           @� �  �  (    T   
     3ϥ*���P��*"(R� �R�%T��J!%D�U@J��D� R�$J�I
%TP���(�(��$�   mDB
�T��UX�3ς�1([��@��:�6(#�Tq��XH��B����
��	� ,�뀠  Q����-��}>�  w0��yB��Ц�r(�tP ��� �uEH`:zo0�M�������� p $ | z
�)A%"�QIR� (> ��� {��W�o0.�=�׻ʥUp 3�W���=�"�w� zK�x"���yz ��xR  � ����A�t�I�`4
�=QRs�������`���{� :2 z���(���su����s`�{ <�70�`   �>�hi (� �U$�U_f!"�:N�� <�S�������W��$� ُ/@�p� MGf�p ���c�@�>AA݁��  �}�E}
ʏ�p���y�P� �@�@\��� ��s� m� v�,��{��P��   W���� �����@ *�!�}&�M�[��9�Aް q�{=�q���`����9�<�P�p�@`��  ���  � =� 7PJ����C�lX	� � `�� d@4d�P  �  }DQ
�)D
�
��� �9����R� ��w`��#��[�X' ��� ��   ����`�AN���� ;���F�M d�f��      jz��*   �  S���%T�2 ��  ��T��J� h     �d�&%)#      &RR�G��� ���Ѩ���M���MSCG�Ѵ�OD��?�>����j�W"�:������gY緎��� *�q���
�U S���*�� _�d��O�~=*�  ���U_�*��l	S�`EW���~o��݀~�� � 0�,#�*��G��S�ReOG��; ��m�vʛd]���Sl��U�aCla���al"m��6�&�C� �:`X^YM2m�6��6���a���l2;d��`��l� � m���Wl!�P�"m�6��6���m��l!�Wl��m�6�`�l�� �0�l��Wl��l��0ev�exav�d���Cl��l�� m��+�+�� m�6�a�L�l#�@�P�P��C��2(v�"v�(m�A�"��Sl���� �0��	�P�(	� l*��E��eD6�(m�@�#�"�C ���*aQ6ʪm�� ��t��TCl��� NA��aU6m��,(&�UM�(;e vʈ�:dvʬʪ�`Ev��ev���yd6���  m�U�
�t�&�@d 	�6ȁ�Q�
m��@��6�;el��m�{a\��l�,.�Sl��Q� d]����|d\������Ɨ0z燖��arW�uP��)D�E�C/����wc��z�wd\��)�v�t r4.�zd\�f�su��ޥ$�BB�.8�E�%}ŷ!�V�����6���:�]�/�a��>�m���źE[������xA�#ہ壵NC���w���8��(������0��ܴi9���fL3%��y�+r�a�Ͱ�[��ue��i�gv񁯮>Ś�(;�����ri7�\{�Տ�͠��3��R7;��:�N�mɜ�ڊ��s �A��ڞWn.�:�0<" GwuX0C�}.������O�>-��Q�����;Қ�q������2�Ҽ�YA�N;�(ɹ�b9D'�9�v�=79��0V�S�Oa ����Q��:�{��^t��l!-��Ot�"��; ��p�&�H�
35bƷ"��shm;�-ۭq�]��`e���r���o6V�I���e�Þ^���M;�W��Ғ�L`���Ǉ�&�q�$pyn�9ر������:\��*o�)�ݝ"�]+��Je��^u��V����ǵ���Fc�:4Q"��s���¬m�/�8��[}s�����%^�,�2�K�K��~`��3n���Fڶ��o	_\�;���hf����ň��.�(.��2
���֒k9++��bC;-b��Tvi��_n����;WGͳ;K\����%�S�d�Z��Li��
8���sy����a��5�O7;�Z��2,z7^�H�Ҟ�sn�+�j�&�Ki4�d�y�D� �z��Cu���Q8��`�Vk`Ƕf��i����n���tc�s�GQBC��WL�d��.�L`
��nK(��r��-���[n���vM���X	�1� ۷NR�l� %ٳs�<8��X�Ft�ÛF3��rw���z��}�&��R��n�Ƿ�A�lի.ϷT��'��SI�]t����X�³pL���sV�dչ;��jN�K�i������p�~�Xǈ��V�,k�9�������V�=S/25���
�<��}銸-�;���C��ʳi����u�d&��[5=��Ʌ��m�)�mK����'wPg���O*ѕ��p��Uw
LAlKf�+O7sa�ڥs��Èy�U�Зͭth��wļ������`r��]�vꪙ��K`���1���r[��,�q�����J-\��p�&i�ft���wZ�E1$9�u-#�C� ��
���H�B�+f�s�N@m�x�ݹvXM���;U��!DM���f�xI�ȼVVlա���������D���dr�;s�.��r�a�Z�1ur���i�,�5�淖<���+*é��ᗦ�u�rӭ&��Q;��܍��%����˵+�$dI�b�D�ƕ�>��o��!s�)���6�Oc�����{\�bR��� �Ґ$J՜CA�ie�.ͽ**8⭅���/+bve�$]�T����#/r��܆mi��Bθv\�$���N�|�Mv��|���3v��L]��c�ٴ�k]�`�����W,�zc��l ��e�n��n��.��`ط�k��$�i����
�������V,�����z��wC��V���}�F��G�]CP��gv<����]òU��{d�e.�{� �.˹bw�$��**�
�0Ԡ��b�#ur����iK[;�S�^7H����uW��p�2�!z��H��]���˯��s�R�<g�Cw��^i�I���8��Vj�N/mG`Mod/��Ħ�i�5F�3� .'j\UnI܆�L�۫��L����[{���ylzV
̠�?s���LԪ�Pxv��C�M��Y������F#	�E��B�ޓ�ע��f�w:yv[:���,�ʏWr�-�(����p�������ޔ��)����8�\�R4��-��-��/4:n����������f��$�`99b��ܘ���&�,�Ж�,r��LQ��C����2�v�wVq�{)/���Е���T�b��/t��m���/y���v�n�%�m�ǹԌ[�޵�bL�Л�	� �0=-ogDs6-�Z��T�noa�ɸ^���C<�W5��5װ&�ߎ���)���]��u�^̱�:��	��*�p>�L���ab"7QC'$�cW".�n�<)̜���f�9+�5��q�d��Z�^wV��9g8�,���#��dw��y��,X���=��+�pXrQ�����ut$i����$�:�^�}�5��9���"v>v蜳u*�e g~圥s��9!��|I<9w�t��g�vݬ5�JHr�|��#{%i�O8����.w/�i(�Vtkj,!,�+��j�t��ѥ	K�e�>5מQ�75��j7��"����%�NmF�V���l������z�zW��K�p�:������&t�(�C�
�^d�*B
{R�aW*~E�8�~�P���×ol"Y���B[�#2���{w��8u�5�g�j�
y1�}�l}Գxv+�(+$撣r��+�^��f=3Eǁlc:�vm�HK���ƥ'&�yӂ�B߸�jP>Iݲ����Aڞ��xw��_׮�,�D]���3B}ݰ}�T�{�zn���w�vK��C	{�������7D����b=���R���wP$��e�ц��|�����B]��3fͅO���ڱ��VY�_#�V��͙�Nۂ��`W��^:lxm�$��+��=�ʇjސ��KU�Le�}\VP���<@��8�5���3;+�v�2,�`�8�1��gn�7�K�'gS߈5i��kwQ����v��e�����M\�������sn��K�n0�-�����sG����v�v����W7g)!���9dGX�
��gC��<�b�w8b�w)����U��wVs}�P�X�B@	��>J��w�U�mgh�z���5e��k�`�������26���3F&!��Af��C��i�9y�=�����3��κ@]�Q�c��gKs�NCܱ]�Vf�WO��5����tB:lH.��!,r�i4�mB[{�+�+:�:���o�c�>"q�e�un�]�n�~���1e��<��9�7iV�V*������}��e��F>�7R����35]�(/$�^����7��,�6��V�N>1���j��;J�dKv�,v�Aq�p�hKU�vn���c8�ݰv���K3R���g�ْ�:r!=CB�������S�B(�8�͑v%�7��~Wy��/E��-o�&5����
;��g?2<&�0/b� �J��[�j�[Im�IL�p�˕�S��бq&��yǴ<���.AM,^*�����+�J�np�s^��JۙU�B{�ۊI�{��6�����sIFu�L>7'���#幠в�����0�`�����ƃ<K�+&�4�S�gn���$��S�3����(-����Έ�q��[��v��.���svu�*��Y{ ���%"����F[�͖\&�����pnz���3�r13��X7���l��Nǆ���n6-�I����K���XiUGn6�k7.𜨸c�;L駨Uq��L��9��DEpn�f���ȱr�eboNv�w��r䇉+:,������p��z2���,-<W믂����p����`*�J�5.��m��{��Ѧ\�~ZzXqc�c��*H��6���w��9��Y�.�Mz	.k����ް��Z��h<h�sX��.T���n�Ӛ�wP��
 {�i���b�4n�'%Δ��:k�U	���6�{t��29&"c!Wv��D�^��}N�LU��45���T�]�٢�ލ��iA,a	Q��M0vJF�n��c�7�q[oF-lc��L�JsVN�;e8�g(�@���xv>�/3
v(E�y�(�R��)�|�݊���x,]б.�Z1�ʜ��Q�ҕ8�v�yoK�w�`|��w���su�{��A�R��h�͚�C�XIg=��u�=���R�C��2��!NH�r=j�I�����*�>�e���V���9⹶���{+a.��L%XAql�c#{r��r���GF#��0�����-o$�����S)#_`��nB�[�AC!�7��m�lk���7���trx��93����Z#�-�v�����1-��v:�JP*k*�3�.L�ܭ��&ǡ���ӑ���!V�8���]�.�*�ɮ��i�wj�9�sзsf��ղ��6��n����n΋&����9^�(�lx�u$$�RH��	n�לߴ���ed�v�T�%��ܙ��+��-��Oi��$�a	1�8wú�Q�^�8Uh�u��Z��0;+�zy������rߞ��'�����Ų����H�W��B�wL`���}��-�'�X��9�dvrq=�����Nݖ�{9�r�}UC�}��-�D���:
z�Sv�b�N��_�γ@Z�2�3�q;���]��z+�{�\9�vr�t�Swr���-lQ�����Xs��V�/�j�z��zZ�7g3�JI+�ݒ�[��\��yx�ܚU�m�������Hgv�x���\�3q8�\%Ѳ%�N)���&-�a�ؗ!�j�wD�o.���g|�n�ȴ����@���1����O��Z��D	(��V߶�0�T�r��\Z9��n>,�l��\�D�w��؃H�)�pQ2G�c�i��/-=�r��Gx��0f����+��k��|�:�ͯ��ԋt���.�n�C�~��:1����l��s�!V��6'D ���r[��T�M�kn���uG��gm�a�;w8;�!�pI�ND՚U�̷w$�t�c]�;f�cE�hɷFU��f��)jOjAC��yU8���Y��5�T��,��M �0��=ݛ��1�VU{X�C������[KAz�1��.}��{��b��)<�;����^B0�lv�ټ��neszd�no'�"�z��VA:�����XT�(WRv�
*��˂B��)���1Q�Ĳa��U�~�w'n�$74N���!5y�mo�F� F><���w\B\���cŪ�ǚ�[d(k7Oګ[�6]�XsX��W�_����`��g_n�o~�gG��js$i�ߘ+���v�rl�7���!gu�J3q-�H+��v��;��MS9�׀�^�N�Z��õ���(C��frץ���h3�f�G ����km�Ť,��m��'&^]=+a,h����[��'K7C�wU�l��c�y���Vpxw{g^��W{u��p���4����"*�gnp<
1U,O�t޺)s&����ە��{�֦�9�k�d�j��ljZ���
��-*�4����'u�Z>fS�8A�� *�1����{�
3R�t��<�w\�6��-%ĝ�^Y�4���Üq$hd��ar�ڪƷ����k��4o8���/U���&�x��m 7��623��Y�;A�V��!�f��3��т͉�L�n�xI����M鏶S��pݯX,�v�s��L�n�~�ӄ���&�ܜ2� ϵb��d&�aL��׸�%ǵ.�.n�Jp�͆�1v�IF�.�N$�]>����/�(M&�&�ad�W ��`O���7e�w����cx5�Ý�x��c����[T��)�5���o�9fuY��[���-^�y��E9��h��JW���+����K�:�}n�~�p<F�۸����cֱZE��j���S�HY��7�	v�	0��֐���Y���Wf\�$��AA�P<�4ٹ*�z��u��v6Yw�Y�K�йv<��фe���jXp,��:���i*c��8J�����4rh}Ci�����͝{)�z�۳���9�E�y��ؚbFh�P��leM�L�ܣ2TL}�M��Y�z�kz�$�ɜ��nK&.7m�.S8i&s�;Ov�0˄���p{|�V���I��b�<U%i�K˞ɐn��І��1p�E���Z��c�r�Ō��xMɶ�%^�����<"r�&�]s��&W�\gM�)�Hk՛��q�f�}��x�u��[����K_Xe��vSr�B�:ͻpc�9���K/I����ȑj�^���2��{m�7���}��)��J�e)��o#Z�����`����Β�ô�h`a��o0EN�Z���䑙J�#Xl��.���%��A�;�،���yL�r���S������C�6�z�EPV!5>s�8۽Nq��G������¤FM�5�D$!��;w`��6kVţm�Z����Gr�:/q�^�6��Ȃ���ׄJ�nq@��{^����U���_Xr]�xЕ�i�7��-��ڰX;��YOa#�^�Ji��y�v���)	�,�{��|.�1�]�˹�j�ob�E��SFo���mY�6'��Z;
g_�Rg��3q/�aD�
������p4��o!�`�o�<|��wo�Dih8�����5Bi�h�d�i;���,���l�Z#H�4���}��pBB?���(�'$2��ۯy��OS�}�C��ǧ}�߰~��;����М#{�&��[/��*u��3[�e�w&%��#Y�o`�L$��x�+��vn��т����ߵ�G���zs�������/�~-�
�Q.�x��C�>�i��'撙��>����'ۤ������Ǒ$�ˤ���y�w�#5���~!��,ǿ='!l�
E�P)F�AhZ �i�E����ZB���D�Pi�F�(ZPZJD �)iUB� �EE�U�
TV�Q�h
�(U(U�T)�)@�(i�F�Z@JB�J
�
JUR�(EJ�hU)��� (1�0�e ��M��0.0� �H*�"P%��ҭ�% �(����4Ѐ�"R�P���B�ҨЀ4 @�ҪP
P � )�a@�q��L.0��x�3�x�f�Q��uI��&.��>Z�/s�8�0u70:�]�Y��Naq!���wqy)�0P�Fd8�a;���<����8����;�8��;�
u R��!���C��G�q�MZ��_�����P ��}?{�t)���r�QE�����o�������S����K�w�z�ミ:���s՗��+�����?{���G�ݓ�/E÷�5� .:;�q\����y��zg;������|��=��[�e>��B�|�}�Ȯ��v��!���[;%d��c�B6$2(N�3f,�3!Ĉ3�Q�=���L����Z|"�SB��xC������菎>~�VX�g�ӏ���xoփ����x��,	`{,!g�W��D��"��؆�k
nԘ�xo
�8ζN@ƽ�nr�{�}�(a͘;ޜ�J%�p<���ܹ��DFUE2�d�K>Y��jɛ���0-��'z�!�r7�~��r��dK�S���ۅaR���0�v�l�GL 
��|}�{!���:�rt��8<%�vs�)��Tn��u��9�ˀ�{}��|�ݽ����jN��h=�#=�So��&�^�{������fJ�i犚��o������Kn�<ٓ}����
���耹�����٢{=4�b�w��j�/ɠ4�����M�[O���D���w���-���p�E�9��	��o����S��Ė��Q+ˑ���X��Y��Z�ۥj��݇&�"��%|����	y��0�
k��mڪ��xﺫ@��î��}���ި���ޅ�fƻ}�C�*�����N��_o{Z��Η��������tb���:+qH	�g��OM�Gwy�|�ݮ��lT��c���k)K����gAg�ύ��������]�z|ǽ��I�sUG�G%}���_,�i��N�~�Ҟ�jx��p�#�y��ع�j��[���F,��f��y�a�~�_�����Cd������2g�}ٻ�;�O����$F1o��Ş(�>�98���8oz瑋����zq��7�.��Nf�zB=���>!w<�9>�o�ȭ��ۧwɮ���]�^�7�f�7�.�� �S٬{ğ�<SӞ��8����N��8��������s��\&{*�n6��o٬�U��oh;���y�wLz�q���ד�E]^wy�gf��~�}�w���E�a�<��왡�R�ww5��`�r�;�^O�Jܞ� O<Bp���	�mh;�ބb��m����_?�o�?B�=]�o�F;�B�kk��|�§����\Lq8���zf�;��7S�ŷ珽y�O�s�G��ԾO�w�G�KNr�OrÙ{�Tޝk�Y梁��T�n��Y]�{��e��bn0�����9{�&ʤ�v�Tq?�����G<�=�ns�g�nyn��V������ӹye� �R���'�pF5S����7)�������w��->0̇�vz+�򲏴���� �˽��tC��R��P�z��_�D�u�^<{����s�wލO,���rj���!_���d�㫸f�"��{X�n>����3s�7t?y�&�}�Q�2ķ�$K��$g�NLջ�#�qu֧��rt>����O0y*'��App0��.�Bs�K�7��cË��Ǯ�>��t�*Z,�����6�]�9���iU�k��� 	��]��}��j[����M[��ŏٯp�:�f��}2x�^c{)�tl�vz�h��{ogs�ai�p�+���kK<��7;���C�<��^��n�שܙ5��O������`X��u���n"s��-���׭پ]�݇�.�͢�X�s����%�\^8�\���S�5:PB7;{:�=<�77W�2��r^G�o����5F��z�=�l�}�Y�u�#<�Xh�P�n]�%�}�N�M�G�޸&Bx#�g�c�,���I�d��b�>H�`�yM�s(��>�w�~��ޣ��4�a��:���7���#y�f�Rox7�����vb��i�<W�;ˢ�x/[v�t�x{��<u(�Z�=	�=++G��%e���	��jȎu�y�Zl#ڭWk�,���������fi��ݞ]6r�7����ޞ�^ѩ,��1݋��/�>^3��"�%���A��y�I!���SfC�s����p�v_C�t4���I��ar"9���Ƕ�D�:�>Wڼu��M�9��~�Ԗ����漲7���[�[�]����z�������7$����K��`w�jl����l��`��Ӊ�����gY���Ǜ(�~y�\��:���9�^�����9��V�{}��/���3_�[�ba�>��C1��k$)�����v^��آ��)�3�A�ݍ>�;uꌴM}(���/w�{�C��E��{۞f��4&��Ӎ�zq��yՇ�㜸�ʢt���1���-<�nykxo?b��Շ<���YQ����������Z�����;s�}����% �F[�|=�m���y�wf�vi~L91�;���5�=�Κ��frݚ<v�[qՔd�͹��^�;����(��o�l���e�7�G۰�AoX"������ުz�9C,�.�at�f�0�A�<�d���h�b2�W}�m��ܝw�sL��k��=P��gI��v֙v��g�ò ����[��a~�{�M��D�WLS�6��}�x��o�x:k�<������<=��A�w6�WUL\(�γ��|r��Ğ�1��9�����kO5S�H<�	>X���KbF2#1��6�l>�R�L�f,��F,d�y�3,rٹ�;^�/����S�7�7Z/����["�'���4ٔg�b����ۺf�o��L�<s}�������asζ��.�'_)���^��U4|T�NGws����?q�/���m r����N�����s����=G����X��7�v9�Cpƭ�o�p�V�����_#�4����=�����^����Ku,��J���U0���{=��'�M� c��&�Ϊ��{B!x�!�\:X�27�|tu�����g.�w� \�\��%
^ܹ޳<�p�q��{X}wf=љ�lH��hʥ��c����������H�g�Ι�6)��"]������t{D��3��g�o{�]�H#��=F�����f��Pz�v��Zq���;��N�1�ǿy6ǀm��G�%��Tg��bT1��MZ���rrT�%�ϡU��;�BC@\��q���r���d�<L�-Ľ_�����" ����{���3�-�jdu�3޸u3�g�������y����o�WG��1@�S۱��O���s�<��oq5�μܘ�mX޵� ��n�8&��y�ė9v�]��#�Z��m�����xp����}Ɲ�^A��/���/�Mˈ;�U��޾��|��,^�?g����;^�pN[�b����?\ң��Fʹ&���f�y���E~-�g��x�c��M�<6��޽�vNn�wbn9�~�}���Dƾ����Q����h�ޞ����z-�טȳ�|j#�ض+���e~e%l�4h�M��N^� ��K ŧ���iH�����I,q�5�����mo�pC#�U`P,^���:C���A���^8[��Mӄ��ca��g������wa�=�D�g0q{���:��0)_E�����N�pϼ�8�z'���C�)�w��������#��0����ݖ��W<U+�O=���>j|w׎C�K(�qDH���@�r�`�3�Y7��6�{&�֭�/�yvk/w�҅��b��Aʙ�Of��o$��p��WU��f��c}����˂�������v �y{fv���To�l��W̟P�ۧ:�=�W7B�z{v��Vj�p:���-|����nr���j���9s�;�j܏���=��{��=��Ro�(Lo������{�0��a>�μ>��Ow F,zA����Z� ^�}dIrv���S��>��}�t.�@E�Tx_���==�L�,���ka�^΁v�&>Ȕ��D��o����J�Q�{��>��m��ޔ/"FQ�L�VԽ�������3���"~A_z�S9}�j��t.n���;������~�f���������XsD�=����sW���p'�<�l	����Ҙ��&{txܾF� �a�(wm���Cѓ�Y\r_�{;�������0ޔ�Z��o��7��g��Q�t[����]�3�^нlL�1!��<�C%B��ʊ
9'��8
��=����3�v�U1i3�#�[�,�=����6�3�g�ׯm���>�=�oK�izؗy�Oqg��]���R|�DY��4!� 6�d�\J>eǋ�)ޞ�����w)�yw)�;���6��z��[����v�1��l�ԮOlM6��wo����'^�q(2��O{�x����6�ˀDn�R�t_Hsσ��s�����q�ͻ��W���1fi���\>��Q�r;�ޅ��j�	�F�x�yѬcP3.�+��9������P�o�6eWˌtzQN���)���L�Ww�RY�ɪU� !xqX�֍ڽnN;�}��bnv��[���i+o���"�N^�®��;�<�6<4���ǋ�w�0���,.��"�>����=���wٝ1�^9>n���=����}�!w��6�o������I�	�<)�귆�z��U�{�.�x.��Pva���ت~���La��x��{��e�����m��!�g�=|���5�=�|߻��{�	,�<(�ņ�D�x�<�gw�9{��������`Ļ{�E�zq>��{������/X��d��t2����v^�>�{A�Y�<���u{R�N1"��o����o=��j�ξ�jɌ��������a���<CAv���=f�s��{��h�p��/��z_,��	_sz����[5w�r]�9c���N�#���ko|-�|��HsH�c�/��Q��=�k��sqg���c�0U�z�� g�Ti,nx�O^ཏ��{۾^�CK85���O)�q����;����o{�:W՜�W�ޒ�j�F+��qf����ˬ��[���<���_3A=�p�ϧ�C�����P�}�	*��Yޛ2�he��LgH����h�z=����v�S��2�{�>'�����
ĸ�7��lI0}�n����xP�
L�(�DeTɄc[���)��,S�F@��83C��`O��V-FN2�B��a�ëئ�e���̭/�G�p��x�7�a�_[w��1{�z�f@���>>��	���Wo��6���ϧNսd3��?g�ҥ�Z�lÂ���!���Ð��M3g%�^��9
r<����?5�콇���F���q[��Y��'�r��!Ī�Dnwx�"���g�+���۾���n�g�������r�MQN����
n{��>�tM�O��,�g�<}{<wA }�,�>��y]��N��"��ܫ�}�����	�V�s#�٣���O��tL�`�ðO���;�/{�4?˨m$�o�5���X�6I��m<�ӻ�dh}�5-z�tQ�
x_�Ѹ�����ݹ�����ۏ�ʻ����H,o]��2���:;��=!W�W�Z̞�
�t���T�;t�e���-
��}�/�S�BH��;���s\��e�@�{kS
�g�4+���|}w�?c�|P,�I�����;힋�x�v�z�Z�D�zS�pu�;�}��x���;�����VyY�{�o?)CK�}�[7x禍�/}��Ġ��e�����^�'A�:�jLx��<�9��h0=��7�oz�r�#�ȀY���m�G&#=�g���N��q9�J�Y�GS�z
�#ğz+�wpS�d��U´���������]���:�v�����(^��}�gKU#D��5�a�7�b�*�Q�,Ec�y%�5�	=��?G���ދn/!0�o����"2���W�z�S4��#|���T��z��{Wq.yL�E񎫩k�����l��5��T^ߎ�2�~��¨}�lGǻ/�z��$�ͽ�F�S}�㳀��7���9r�����R����#����bWfݛ}�q� {�|����Sit_]ۊ�����zM�����#�~J���5|���^����J+�Mdn=J/o��#�,~�*x��{ҙWq�|��ͩ���/�F}�+:nѧ���<�@�F�?S�{�mb�em����x/z�.�9Z��2A1o���od��#���bۇ7(2��o�N�jǏ#PǼ�^9�-��XR��W����������}۫��L<��1�O�	�c��4��n��qOza]��'��G��D��W�/o�̆̍>�c<8-�3z�ª�S�e������<x�ڲ.T�5{�<��,�q`���/y�l�`�$R���(�����������]�jg=3�Bo���f�����3+?z�5���
gW�	��&M\�&*����>S����xA�\R{���;�.�?l�tc1/:�]=[�4{ ~ý��:)_=~*�k�nP�36�v��^�{�6)�=Sw��L��7�t��I��W�K���tN�$ܗӲ����w�A�^�aa�r�q,���BJd�23 �'Vu��fq�Y��HQ�y�O��w�٥�1�'�8�2��=�mOU�^�1�i�xz�{n��Z�B�n##�{۾�تT��E��^Y��W��`������s�{;��ޞɹ!�u�{��I-獫W���L�N\C=�y��x<�{�\����^�-yË����K�;h�x�(H��n6�sԿE����qr&��y�z;�ix��l�Nb9Cd�q�1qG- E�g���|��v{w˧�����A���^�����$���O���Q훗���J�u�o�w�;���l����v�$k�>à���wic}��gyl`x+�h`/35�ݻx�ۤaw�{7L��n��3){�c��Ac���˾�Gvm�ͼ;�Vk�^Ӽ�7q�:����_��j �Ч���������~K�P��p��3?7��߫�xxxxx~�������0}�O��q�x\L\f�V�i6nJ1`9f�#]Q�(Z�kX�@LVjA�||=x_^,l�!Cym��R��:]|�q��Qt��f�.�^H����L+ku*��M�a�%�,,��Չ4e�.�jj�QY���0����u�M���̮�G�#�! ̝u�,����2�v������E�J$B6k�+`�х�U+Mk��.�f6e�2[��rFf�nJ��2��5�MR���%Z�^u,f�tK�������+���Y�[iq��Kڀ툐���-�6�̤d��f#qo�-'[hԋm��3f����1�f��`��uҚ���GUڣ11ƆLP
�i����׭mz�Y���k��;H��VJ5�\����F��0ٍ�Kvt&�HB�.Ƌ0�4����X̺�7^�Ͱ!��Gs�l�e.B�S�ҍ��	fV��.em.3s��/Ya��Gh:`�ٶf��uK�a0��I����v���pka��W���TшFm���U."�jьu��l����.mq��{G%Y5�A���Vd����M�[�#���.i�)�%��-�&��/XM�[Z��Y�E�i��ۆ�5p5��taV1��;r�H��	`���lA�;B���h2���!�Mtvt6&5��l,�l��j:���iZ����KƷ4J�V�&։c�k��L�1k��c�\��h�YWL^Qf�2��gF�v�KX��np�B����Z����a�t��k�cEj��TH\6������IkH�b�b*�
�vx�Q�)��Zql��\��5�;�j��-6TիJf���p�v��ٕ �n��#�i̥|H��0`��5�j֬�kV,�@3E���0L2�-�l%�n��!�V0#!�:�b�Ff��q�L�UYXf�F�o+孩���l6*V�RӪЊAIq���L[��tBV^������F���A��c8��%�M(ֺkU.x�,��`̼(���`Le�;���`B�ǂ4N��l(�e�TF�J�m���h��8Y�� CdQѬLme��"v��cT�B�B��R�W]Smsv���ivaa]jv�-�5�B�duv��M�v�R��w)�2Lbi��l���z:#G.6�f��@�`6�+��PlŔ�ʹ��h��K/# ѾxO7�*&�e�k͢@� �MԈ+p0��8�6D5#y�q,
��H�˜�*��]2�3d�i���8�M.�\�Sh�3h�hK-몪��Z�.���%��&��JI^d!�G0�ڻ�a�B������ZC�70e�F��YR�o(���+Nq�Z�ɶٮ���6��cp�U#q�ͅ�Ma\�
n����QpG&�u�f�+3�����tqU"Tn%���m7$�F�+bKq�6��䆏3���l��A�h-ɱ*au(�&����FP�&q�1����	�q��D��Ԍ�by�m<�465�XǊ�4�1h�,u��d�t^����2vs�	n�0��X�WK�� �	�� ,-�\��α�R��)2q�Z�l�F�"�gXď)��4����l�l�W�avM���74P�sL��nŉ��m��
v5�����05�@� 2%��W`c�7.��ٰ�ŵ
0��v�0`�����Ë�B�:��#�"����nP��M`�+B�n6c	k*�h�-���(�驦�0Ŗ�3���
��1�A�6(�;\Ǟ���0��&���k�ی04��\�gK�����4�H�+��!��wٲ�E�l�Y��[��T"b�c4��͊Ys-m��1B:mn�Y��b[�j�nx�8��c)
�@6����ؤ��6`rĳ1���gL�ibk1�B�0PfҲ�f����k�kٷsn
�A�G]N�a�Z�.�2^��]�L�I���J[���3a�e+i�P&�X�4!�N.�V��ez�Ŷ^�i�La��3E��j��=����!ͩA^���y�V�lf5�:Ԛ%�&�-����::U���l(���[��R=F�Hjх�6K�#iƬ+e��8m���.���$��GhY`��K��X�LX8����.qx冻%�A�y!b�
J��riF�̒fpu,�@r�щ2:͗�[(� �]�`#ፑF���%ԘYk{Kf4�M�h��.f����
�.���ƽX �JQ��gXI��y����n)�ٮ���3��%z�8�F�W�Ɖ�p��(��RYB�1pm��#�]�5:c ծ�[�4���ն각l5��\K�k�tҺ���u�1r�j��m�4L�Ix�RK�c�EҸ�4Ҕ�6�:�E��6��Ƌ���
�UJM�E��at&�evəsfѱ@��[�j7���y����[-�	�aiB�y�2TЃjEG8%vk\����6e�:͵�-с)�]JL�e��i2��v�s��1�)M\��*�佊�k��[.��]u2;&�j^�%JSb���la�֑%�2d��٨��̰nBh�i\��rcZ��KiHAP��h%�m��@�����+�v&|�#�K%��a[�L�,�FW\�3%�:�+�ff�Ս�̻MNy�s��̂BmnvڌÑfm��PR�35W���$n�7\���`d%vk5�(hl-l91��7�A58%g��:$ա��&&�I���3��i��(�v	M�pf\�( K%�V)���l+t2j4V2Ӵ���
��MF亃t�-��Bb�hK����kN׳,3��$��0D&Dt(���5ړm*�7,�76iw)[.�Zd�]��7@�"���K�nkvрB�YQJ�ƻ.]1+*�cJ(�K�g5ԍ�ҖR�f�9�yX�KY�&����r�2�ɬ��Mv�JK�M6����!�n�Il(Q�J�'3��w!B5.4,��+--�����E%���YhB8�fv3JӪ�SBh�3�kH��3����fZ�E�k��+���H�V۞v[Vclʖ
 c�)Xd�j�]]I��e&��,���=0g�Qi<���pm�V����tnH�X7u�yJU�%Q� K28qb�3�E*�m3m��2�#e���b��:�L�:����Xi�)î�4�]n+u�	��eJ�]���!�u���Y�����lո��0�Y�ZJ��6ZZ��1K]3�GV�)G �Zg�GQfٷv�C,бb%C����i5P֤�t-16����r��8҉j�M��ͮ#Y�ܯn���D,,JM���\�5B�֤��t���[���f���`��[hB��]�m�f�gU�@��sl[��r����ֻX��H�W�K��c��Ldn��-%�TH YfK��e�q��D����1�SǱ��)�sH��� <k�(�/\&�#(���٭���Bn�kX�eK�-	��3I@u��s��'���+����l2X�6�-WZJ��Z�av%�[��Ci��U����әM�1"#u�l�h"ꨨ�.�i�JK�E9GvVMٛ-Ж�pM �&��%�K8 #fm�����%n%��Ԣ���t.n�"��5���)af�ilͥ ���� �6雐��E�AB!e����e�ѳ1C'*j���m����Qm�5u�+Lx>B�y<��Qk0;+MI�Xr�iB�j72[414��r0�Tj���1w1�3��f6 �u4�]��r����qv(m�cMo
�������^Ĵ|�J��Ҁ󭣴p�V"m�]��#���,����4\FƯRЦ"7]�a�aN(�,�(�5�QY���n5����H�emK��	e�\ �34͠ա\J(K�f�5Q�.�3+���V��ٮ��E�4L�j�a��^�ԥA���8����JM��l!
c;m	+�.S9�kk׳�ʞy��Jyt��=i0o.4�Y�]AWI�m��Z�P����֮�$�W,�̅!`J��mnp��vQ�5�56,԰r��h ���M)���.��X�$^�2m��Z� �FP�Sd�^�p�Q�bV7 C�p�14�0X&���1��]����mV��^uե��!R��Y�T���n�`�K� �^�c���0k�e��ٞ�5���(��d+�®���F���)m�e�
�!��R�ykG���||�Vxifv�1*��k��4&.��bjM��eL$1�!x�FJ�{S�VR�\^��x.5�X��*`�u�\����Y��3-���x[k�H�e�1�z�H�^�tХj]�͝����6�s�R����Jk�a��Yw5�#�%�#*K.4��\f˂Y��)32�2l���n,�R#M�+]F���`GWWhj9JT6m��u��&�#�ŕ�-�j�X����i��ha�������[�[0�5�Z����M����).e&�2�����)�5t�� �׆]��ir�0Ԫ��h�,jى�\��Ã3UI�pe-�����<ks0��\�*������&����k0��4�b7FIDn���s�1.��`a�Y[1M������X٦&�L<�Ѷ&�q���֐�Cd4�f�Ҁg/.� b��u�tZ�с2�eԄɦS�cZŶ��h�As�v��+�h�.��M-fm5�ԠdF�]�[���T�_7�2�-�b$лbtwVR$-,	���tH)؉6�a���s��2�,f�a�&S8�6�L[B<���-������b[�������%��ε�� ��l���1���Ҧ��6�������љ�6�����$������]uS&��˘�W<����%����q���%�&���4��)�����Q�._<����L��Z`� ��1y��B.�k0�[J��Q��m�c�����+�\VE�Ѧ��ɍ�bڰ��0,�vI��lʉ�Q��U�4M5���r��@/�7l��i���lfK]^�}�u��B�YfR^�X�GG���.�uK���%Y�X-�n��Ж_4S%m��!�*�k�hb��f�ĥL%�"L�bgf�7��}hE�2�+uj�bL�U'�eˑ^E�ˑr)�K�"�YG"5(�QnH����u���+�Q:,�9H)IQ�7tO�\��IB�G$�! s"�"���A��Ba	!ʢ'W"���*����TU�D�vF����"�UEG�T��OE�ez;�n�BI�Ü��s�*�H(�j�L�9�֝���vr9EȢ�ŤAʢ=�XY���&J�"��T�TrT�e(�w2���u�� 󘰢�e�6�ʮGN��E�aQE�E�(*�I���29du�*�*(�D�!ՔUD��i*�Tp(���$�NTr#���Ü�� �<�����gj&ʙDQ3�F�t�3�����s/M
3
����<��$�.��X�ȎR��Gs�E��tȧS�5
(��΂��l }���W��x�ޞ|���3��`Z�nVRͥ�L4��	n0�3�b^�M�c������6�sWf2�p�"�	�jAc/]�^�[)bmal���Z��̈g9]V3�ּ2���b*ݝȸZ�c	[Dd�B�h���́�u!j��l��Z��^�����J�K��H�X�H�����T��΋*C��<<�z��Ŗb�0�UI+e0��4"�\�+"���� �D�-(�k�!��\Vm��'f�1���k.b�f�FX�ͨD�e�L�90&cvu1�a�A�m)!]�CSiD�z�F��J7G�\+n,�K�Z<��A��e�::�
�.M��XKc6 {J�&���b��C:VE5l���0G��4܅��&�M���,�{CE@��5l�eH�Y-���1��f��a�c-�JdK��(D�t�jZ��Yt�s�GD��K��Me�2�Ж��ՕbT�@�qU��p6���[������5!q2�i�2�̼@�kb��v �e��K-L����e�k[t0��3&�M5и�f�MLe�l�e�D!������� Um�w;%қWMy��c-Ύ���$ul���B`�i�Z�Q[m�kb�B̩t�
h�@֏i���WG)
�T�4�tc2ݪaجe+M4J�t��C6�3��ʗ�4��	Mٺ0/g1B2��Q1]��՚jJ�3�鑱�� �.+��,��u5�pɀ���.f�����e�����V\f;��j�Fͪ^�v6�����@CLn�M-�D��l��64��鈺�V�`6�ƛ�eb@Lu�1�k���b�%�V�1�v.��p�HkT.[pD��4JK���� �2�Sh�8�t%�H[�Y��bPQ	vv��R���K���6�`�%x�i�.#i�kV8k]��b���UD�Y�&�K(�sM��h�Ѹ�@���c�<�_�k���ܥq4Ux��J4���3���gt�uܵ��9�RE�K�襷ݑ8�s�+�����!\��1��̰����y�� QcK+X�a(�RZ�Ue�[�S����x��@���	�TO*�+E/ws�1�p��9���<R����,���lJ�X�cN�bHu-k^JX�icm�ly�b��R��ܿ#?�[����Y�ųQ�jf3������gr�jU3�3��[�����~�"�Bڜ����Wv�,��d�?�d����9$ߤ��C��_ďri���Q���i�dP���UA�ۗ�e�Ҙm��I4��ʭ2�5�G�F�
��&	0I0�k�Rd;�{�����f];>�6�8I�k����/dQh����3D�U�୽����Mc���Q׹�ʶf�U���[�An1�٧3mR���$�b�Tֶ�X���"*(^�]4���m���d����ñ���C�W��"�^�"ak�r\4�bj�u�5�V��A����K��o�*��{q�o��+���L�]!�i��l��S��^���`o$�y&���=�ڏ�~x#b��hy����yEi��^{���D�{�=;�݀�:[�ػ�]ΰ�:g��R�Ûq�Pe+<�Bh&W����U���&k^�f����Vbb�=W���Jc=U�
����E�?r�������H�;T/��^9�мi��m�����u��������I>P˻���ֺXr�3��k��.n`[���0�N`����j��>1�7o��C4�sW���M��5�I���,9��l���)i����l�y�8aGmaW�ivM��1�Q#4�&����14u���~{�>0�ħ�&9-Y�,����&w����v��Ƨ��Y�/��5g�z�Y�q���u5i�����ۻWY3�P��g�M��t��ښ�i����c�Y��L�w#ω�c�{Y�p �2��G;��^�z!0vZ}�:���H���0��w���Y#��*�?R�C{��\���ksu��B���z�|�eLN>(T37J��7��������+n��o��N����x��L#rj2#n���;��L車���-�F��+l'�}w>��l9�h��0���u��7�.�F����	0J �˻ܝ}ƨf�C�gw�i���7M���L�7h�+6��I�j�-a�e]#=9y�L=X�$�I��ֽ���*��L�4���[�]�Fzq��|��;����z���P�B�e�=f����2k&b6�;�;w�L�7���*u��M�L�H;P)k�V�'%O��N�A�ҬV�!�V�el��`˸g�{S�wI��	K'Q���Uz.Il^�i�$���ƽT7E�]�&tY�,,�ra�hg�z0Q����ч/$���p�f��۱�H`�j�����"2r��Ӝ�Yjk)c��C�{k��ٺ[����;/Y��������$�$�$�>>��۴�-L�Zt�`��93����I?��iM-���2�{�[~��0�X0X���F,j÷&3t�ˬ"��H,�ZM"�A0����Y�L� �qt2e]�F���w,��f�Uݦͻ��2��m�$�&7cT�ئ�9���S>���'ֽT0m�]�m�����/R��P����$�I�K�0X"/&e�mӽ��x�[}8�-d����p��:��Y-�Z��%r1�Z��ܬ�i3�a
�;���^�*�[��q��I'�sD�$��O5�%7���9��ۚW�e�ދ���`�A�H�V�������������(w��s��x��\�7=�t�3��8�7�r�Z�Jt���A�?ݓG��K��cҜ�@f`O��=���^�]��,͂b7jRL���6���R�j9�	�ݱUqBl��i���3+ɀFD���!��9��D5��^s��L����Tm�b�u�ֶllaKMluk�m ��n!lQ���:\&��)�H��2e-q0HŲ�ց-���ݴ���lnG\(b\#̹�eu��&���ˡ��(�ZGW�(�Q�&��ƃSm��Ɉ�	J�S��'��8�K��5�2V6�cE�m�5�Y�i�`"���p%�	�̭���^�s��U�$�nEd��ۧ}n�̶�
��L/���c�]��y$�3&�KRlUMk #6�rFD�٬��K]&}����Iz#�7����_gS!�,�A�퇬�6"�i�ZU��]e�=6�.��5��8��V�̆��w��6�>��H���۪6�k�6��mq�)����r��_}yN�y)�P�$��69���V)�tm�[��s*��լ=w��%�9Q7�&�&o�?>���k��L4�����i����ΗU��Q��҅�YM"��}�#�}<~��?IO��0/sNwuV�u�������7R���^ǒO�~��z��mQ:"�e�3�S)/{
2^dK2{��:Vm�u�^ [��!�/m�w��'�_\��m��&�tP����$�o�݌�V!
{�\�_b��6!r��Ƿ�g�z/b�e�m�����o�kx$�:z�anѹdQh�=�Ja�nd�%������A�P5�lmm���9�l�+[��_�0	$�Ef�TS��J`j�Ny鲭�I��ӝ�Xص��Twޛ�
Y*��g�����eZ�&�LU$�n�9��(��kl�m̼f�[<6��;�N7��I?���{�7��T���y��m��`��Xm�uX����cɶ��qn11��J%���kī��y}��I&�v+-̃yu��\H3j_!��l��z��LN<�
wlɀ��Kn�z���ӝ��k��ƪ;7nkG����7��K�U�55BqV��I�d�{K;j�~�K��=�g��ӟ�|��}�wE'o:@Nr�}v	�k�XZ8�?~��ٚcC�༖��*!�!E]��N21d̼&Ł����h����$�I���|S�	�|���)7�O�2&�,[y�oﶛ׌ρ��٧fv�q186!��`0I8�M�Y# g ;0*�ܭ������j�M��	 ֖\�d�K⿟B ����F��n�mT�u�j�V�I����^"�00�l��NڲC��w���Y-kX�ۼz�K��wo�p�u�J��@I�.��ibAJ�K�ڞ�)�)������ݣYY����a}Onh���ŭe1W-u�2�!��L<�$��K2u\�KczU�q.TⰆ���j�n�f�	'	7�I��eĐj"�����ɗ�kZ�Z��L6�@��V�ݩs���U4r_���������n��	3r`S�����Os��o{7�nt+�ћ>G����Y:��K,��M�g�1���h��e'��zvZd32E�����ڑN���|�HP���Vmc��X_F����2J��<�|Y������I�Y�Yn�m](��)�d#E�#���B]ft6b��l{q�Nc4�3s�Y��+$�bq��o��lNo$�*J�j1t���ʬ���e�m^Q/�q��o$�ڂ�9w<��2~�2p�o�fu9!�D퐳a����t*}��u�8Y\�/�i���$�'�S��DiiGT���p�ɧ1��׺��B�U�X�D���03	�L�I�o �p��������5q�73�9m{p^Y/�ۉ)�Iǐ˻��T�5���=���UgV�GW��_j��5�v�w���������§m�E�hma0�[oE�_A�j42��"��{�80g�� q���L�`�u��H���6��M�Č��WFړf�(����kcF��.S��he�v؏kklf%����)TsU��E�!.nl5��qd�L:���y��Ʋ��qY��L]�Yz�[[نj�s�W6�9 �-vQ�ԺԖ��f�5�&���I�i����UIcu�k�i�m6�f�ؔ�P"%+v���� ծs�S\��uډA$_~������=����Բ�c,Ƌ	E�R�4[��Wb%Z��t;C �5���ؘ$���6]U��8Z�V՗�Rۻ�ko;O�iŦ�M�I��"�1�
�5�C�6�iG�Xɧ1�zPm�Yf@�})h�jRv\�>�������"��R����M��5�Z�Uۍ6�!^��*k\yeگE������;jږ-�<89#)��'#aеY[����a}�la�����mJ}����	��C��܇[�v�8�����'0�Ƣv�e�GE]��[�0	(���{e����O�x߾P���:�J@�������i�L�j���i�ru �Jx���܏��Φ~���NH�3*rg#(,Z���.�-���O�o[��!&	7�' ����D;5���S�k=�H�ᇲf�_޾��K���iy�1?oqv{<O"���Y�o��ߥ͒�ǅy��vQ��Yn.Fˡj�V��K��u��)2X^�=���HJ����)0J_�*׸|=VVC���V5��Y�w<U��7�Nb���<�V�u^���&�ʕ9�b�^�)f�3̬�A�O��+Y$��$���S2v�[myn��.��2CZU��5�B�u��!gߴ��~��[�g�9��
16��[,��'=���K�2eX�h�����SL�i^�o������9���Z�e�}.���Kb��
kwD��X^0I8o$�$ۦJl��C)��ލڬ��1Ym�
Y���-�7� rb5���|g����LL�Z]�8~�v�����������{v��嬇Q�vq��AU��R����)~�#����������0;��c��c^k�xS������*ｨ�7��=+�!���Z���SG�Jzc��7�h����QSޱ��#���9�,~���=�vA��h�js�)�fx'�7O��C�a�x�r��C���G��7��ۚ�Ph��t��.�6�T"%���ɡt)X3��d4r���N��ӗ֭.��{�y����ɚ��%�=�A��tXH�!e-M�/�*�1���bi��d�M��7���w4�{��-���嬢𫇴�?a{��{��{�����W�{�@�Q��d������N,�<j4�p��j�Mzb;���{��{�g��gm��Ij�	�Ձ��y�Ⱦ˲���,��Ye��E�����N}���3z�la%w�t�tt�o��H��l��g���/��y<oޛD��9����Os�^7/Rϳ�︾Ju�W�;\�d�VY���#���v��=ek6��Tf�O���c�u�������zܝ-���t�VFy�靼霹{9q�({ 巩�<���G}�sf���A��:E�x,�'�NTz��1�qx!�\g}먙����W��%��9���n�?]#qm���2;"�z��uCo�Be�w��}����Θ��&b:qhOL����ػ��sܣcz=뜲g�l3fi�T���^g_q��7%��P�L���8�>8���Fn+�ܖJ`|�lb�m/ٲv;�Gۦz{���n�,���^>l���0�Q����֢v�1͂�SH�0�l����9r̪��QW(̙UC�(�QW��\��"(�q��ݤr*��J�"��U��I�)Ցl�*�*Ԣ�%6G*����D�*�E$��e�H+����Ujz4+�r�=U{���kd�8p��Z�ӓ��rM��$�L�$ᣙzf�
��i%��D�ݑ�Kbq+*�u���pE�j�y�<M�s�ӑtL
*B ����BÂllb5���yX��r*�h:�RGwڋ�ǊS����ɸ�jO\%��!	22^��h�H�Ra�,N|�җY^�$!�w:�{t"*/u�QN�=����e��kI�8v�f�V\鎁
T�x�S���6¬ΩY�N/q+NE�]d���@��&�m� 6㨕U�
�"��Z�Zn�.Eϛ;�D��E��3�9g�H���$�,I"u�/w"��&ǧ��a^eBBATp�(�K�����(�A}J��I>w9K��Ӓ��ͅ�*B�81U���Y5k��F��ܐ֖-�>�}�#�탐Eۇwn �ʭ�"ޢQ|W8�
 ͸r����4� �ts�Yf��q�*���$\X�����$�&�y<EE�Nb�-�QG������+C���[��^���2Y�CC�t�r�-��]���[� S%Uqѳ��!��>���䫻ApX�ZF�� �[jR��`�l��9��CDC�4��'m �WS�#�붐_�]�ϫK؅�]�hZX� b��c�Ω-�i������Anwp f��q�r_a���;��G�5�ci���^��+m��A7��Ao?�����t&�'�F�~w0�/�����`��#1��Ne��	�Ջ2��r�K��vb�v��� � �|��w<n��n�{69�Z��;��|*��{Ϯ��p��]��Y�����|���/��������YR�ཊ�&T�On�w6e��*w��ͯE��+�{���z������2�4�h9��8tnF��Q^�ԈL�5�VK�5l��E���v�]�0["��rj�i���uv;J��kS6�A���r�y�R`�V,�C?�Ll��1�i����<akm�"�֌rܹhX� ��S&���3q�Կ��>�eވ���q �v���	��ͭR�����}�3GG�N�V�8�r͗�$@�p���~ ]��A����%��w;��r	�ox�؈]��*X�n�0r��n��aմ6�d�y�]Ñ�@@�J�턑wn=v޺76U�K{c�DB��[��5ɘV�A�9�gwo"��>�:�Y�,�<��n�8\�6uK��ŊW�C48�w9��K�ld$�ٌ�I�ݼn���jn���hd,�C����Fb��E�=V�`3�[�� �b{�'L>��o9L��F*��q9v�Y�q511�<c\!�FN`�z����֝�:1��W��u�y����{����'��M+�����h�H��b�OB�"��� �-��a1T{&�P�U�� ;9��[
�������M���v�-�����y^mF��̳
`��;t�$.�k��(i�iY�Z��P��m"i���GK�I�
�ر��CF��W��l��:�`ΠL9�J�[�+��]5/Z��E��
%�9�J)v.qlf2d��gl�]j���D����a�m��)�͑�x�%�ꐻ���%a��if�Y�>̰���q0pA�k�]�G����=c��kxE��������ڲ;����`�v�po�A7v�a���c
!gp~�݀R�U0�EۇZ�#uL.�%�W�C4p	�`�"������*��â���ީ�������_�v~ű�cG}�Y�1
X�n ����#�탐Eہwn9�S:���C�T��3�3�gC���y�q"��ռ"��\���3ѓrr��
��D6��|���Z~��@��Nyd�މ�����ɅyR���S�ıJ�H�w�[ �/�޻��xݿ�L#K\��vb�7.�s!6��6�`k4�.�ui.F�EJ�r����S{A���;����g ���rlC�j��R���q�j�Ҝ�� ��`����["퀻�	�`���϶,�������H%���i�vU��Fl�c��
�����M������^E��Eʘ�X�4e,!�ɦv\v܍z��������)\G�����i;G_�Ӽ"��\����< F�y�m�q��e�u�`�Ԭz�řmZs�2Փ�:��x�oY��1���^�+��;���w�7���"������s�=Ŗ╓��ވul7�(�.dm;�9X��Y�3,Z7J��l�5U����+X9َwn ݷ��nws��3^Y�t�������w��fS��Krf�A�W� ���v�]ۮ�˖��}w�?g��h@�^�m)P%V\�F�A1�J�%������Ҏ�.���o$�������`��p ���������3S�U�.R��C;��۪l��4F$�_��9�#���J�`��a�Q�_^l>�\� j��NCm�y�[�3+]�a��
��z���~k�w�c#�?��:�� �pA�p.�.�z�|�����V�0En�S��ǝa+�v9y?[s�M<�`�R��ysL������{�֝r󭑌VZT%#�A�λI�.V@�|��|}�<�Un�==�­,ɛ���x#y��휂ݼv�<C��V�L����n#�c��o�㪥tf����g)^w�߇�{99dşdY�x,�̯G�[�81l�n���.���lƑ��Lc��|��]/ -��6�������W0}� ��r�q5���9�[���8	�����H�)	V��b��ʀfj�W�U�G�\q�-X��%ߣ�l�u���wpx����y:����u�����xs�zN=)�@�s�p v��� �ܒ�4P�s8 �����Y���u��9J󇡟� ���A�Â.��f�;��]�X=sO����X]���-�r	�����4k�z�0S�v^d^�\7���}���A�ۇ�w0�imge�VE�<��+޵u"��bqS���V�<
�f�}7�>��&�ݎRm��j��9�T�Sf\q�i�sfR1��푒�E��� ��ޑ���N�V\{�f�<�'��{�n.�w���n�z��<=�'�R���D��Wzo��x�l��v�7u�W�j��� .p�T_\w'K�ݜ��އw{��E�Ǡz��s#�w��Z|�#f�m�I��Z78�:e/m*��u��%F������(��dݏn<�ݳ�A����%��;{�5v�n"���o2��
y��ܶ|�+�8 ݸ^"��Q탑X��tc�TPj��dv�z<o�'U<mOEj��`��`;�7�o8l�{9�$a��W�rh��� ׳2D�����פ2��n��5�m���U�އ~��c����À|-\����ݳ�!�p�c2nW��: �8�V��]�Ǻ����{"�)��+�s���%��l�B����v� ���p ]�w��8����t��7+�9�b�B�x+���|3z��`.���ww������8ܾ��t��݊�8$��k��_/U�?������n�5��S�)�;�绦��~ZN�� �>�<1��OB|���E�l�bva�����x ;�wt���<����mr�\�B��E���g ��2�8�`r��P2��b��.,n�TX\bԃV83XshleX̐���X�W٥.��1��*�\�v�,�[�*A��e8ש.;=�l\�����`��R:��#�(n �[e��YbR���0.ev �i�]lB��O<�!4�C���ܔ��cbZ:\%�kX�]���x4�2����9��I��ZY����1��sV���b����c]fs�i�%B�i���sF�G����>���A��8��n�nmT��k*��.�Vgz���u�׋[���ܸr7�="����|n�Ǳ�w�^�i��,[�����:��E�S]ރ-��.`�΁ ݰ��a|��Vh�d[2:"Xp"���=���]�pEݿ�����elR-�O��J�x+��n�u���|��j�c-+T_����8r��o�S>]�p2��c5���,�Vgy�����C�=�.��I͝p�8�ַ��=o.t�c,E�}���x^������-�Pm�	j^НQ���x���n>\���=�<n�9^,-�S�\��S
�O�"�p�m���#��@ǈgP�%�a��]+��\��� PJʤ#��??%�������^���Eݸ�]�o5��5ۥj��pW;7x��������a�o��� ��������;dK�߯�똩~gݛ��ii��օ�rC8���˳Y5�v�l=��������R^ ��v6E�µ��3N8�n�.d3�)�^^d�>w�x�Y�z�����AJPP:�[^8}����d���g
�;ţ�z�8 �?��E�ӄU�LƖ�~�i_��8pԳ�-+���S�=�E4%�2���̋�L��yn ��<{`A�`� ݸr-\&�(��.��S�ÂNwDx���M����8+]��9c�7vnAͽ<p/�.n��c���cA� �0p>��n�p���-�ּt�=��K{1���g3C�����1�8"��G�ۏ\�Kc�=ϋ��c?"G�tM]kR�ք�1Ƃ�`UЦ%����%�v�w���G�,���]e�5����wo�Rq۽��x�+��{�611<��K �\` #��v��v��e���ͼ���=�]���"����̈́8n�E?3G-d��
�f�\�A��}v��鈾�U��`��x"��a����=f�x�����׎��ب�@b�xɚ�گ�+uoN���ŉ�������%��{$�c� �v�x�U7fLf_FR����޳)����xS]mzԳ��\�}��@'���Wn=fȠn�Ƚ�,����U�u���x�5��i �������v�f5�$��A������t�S�bjߴIG�|�Â.�Ϩ���V,m�
;��� o�=�}aO�˙.�c\���2���q�붒���~g߻w��_ G�Í���mBaIu�c7[.�l�[Sf�����f� �o'�k���0u��f˂�ۇ�Ա�Z���3����C�����6Ҳob����Z9Ð����p�@1�Nf?�KnS�0G4��v�y��׍�(u�wu�+Ģ��$�0 �`���q�6_dK�}�v�#��y2a�Ƽ����ݙ;�X���w+X����S��d��m���+���q���붒	����>�9�Zw+CmZ.�V�pA�Q�6h�.���>�ó����^U���t�p@�՘�m��&1�/����ҳ;ٷ�^��Q�i~p?�9-���n�2��'kh�m�]ɫ�Q$a���xN܏������4�Mپy�,�Ϝ�Op��"�B'>d��~�#�sq�sv�A񻷏fϮھWw�B�4��P�b8b��[�^%z$�7�0r�@�f����Q��}kv~�9����h-�3�@�e��2Zkj[G!��Lge�l� ��x�D��.び��v�r.�[Y�R����JK��vn##P��n]{�� Sa�l���-��Î�jB;n�_{�
w��ٰA���K���Y�ʾ�~�i���E�Η��n]��t�;,���o �md9�gݼIM��{!�6�1]k�)�S7���X.� HM�v�Ȼ���S\���<xީ/z�B��q�Ti>��pIvc2�f�+^���6�Ӡ䑅c9�^�.��}v�� ��� ݰȐ���Vv���K��l��m�ժ�3�u}��G��8 ��w=v޷����<On�ݼ:yyyy}����ї�`�5�y;e���ŋ�CSfz*��vOz�rs>�t,"�y��=w���.����� ���
��ݠN�vG��|C�.b~�&H<bz������} T���P	ô����]А�3Jf^}ػǋ��w���7��B���-���v�`����>s������B�Bj]���/U��	�o=�eG���Kt�������Z�=�>��L��l�+�«�&&�m뚹(W���^�]�G��&D�}覯^~�]5�A�rnSn,��mri�`���}|H>�A�������d~[��s��o��>�j0���ר��� _?K:M�<J5��^�Y��Hs�	Ȼ�[���/w�\���!�L�k`����1w�I<]ۭ#v�3�J�zR�K8M6e����捦�\�CV�x<�M^�;t��������n����k�l ���K�31g�xU��{s�ow��]8щg�'��t�Dc>mB]� �l�hh����a���9��9��Z��R֗�����ܨj;vyj�}�0��禳�t���壷$O���i̓8Db��M�J�:cGd�2J~~~'���>E�5{��B���;Ʈ{�p���x�>|<	�"���XVZG�z1�򦸎�O����{���:����X}*��F�Vg�yp�q��&Ş:��?f�l���C6�@ Q��y��ގl�H�GP�s�ӯ��͓"�:G�=[Y�ٍ[����g�q�"sECp껱f�G	f�{����ǧ��c'��1Նs��S13'�!F���$��w.DE�ҡ\��}�]�UU�V�D*p�y�'#�J�k�㣄Y猋�Gy!y�ZJ��k��7����K�"�">"Ey,�iu>��y;��E"�H���^�e���)��(�}G	��TAÜ�R���;����۞W*�޻��wo<��""a�)Q{��:��z�@!��Y<:P	Ƹ���%AN�V�8M̼wj�.E9�r�J(*��Yʏ)�]|�ddYPUpºq�����r��I�_P�ՔFZ��UJ�E;t�&�`�!�Rc�	� �)�=.����;�".���q�-B"u���	� S=J�c���h$�y�,���B���GH�'��=�wr�_u���]̢��!2��EZ��^xuB9�!G�眾sD���^NG9����F�[�E�$��t%�͞WP��*�F�[�^ke�ާ��s�_��}�ڄ��"�B���Q�F��9e�K5�Qf��si��U��U+�&�1�"V�(5�BZ�0�Ɲ���W8l���3,���\���6*�aY.JjQ�bc2Y�u Ŗ��/4�tarF�U���u SE�&�*�6)�_���5�c4l��ٰ�&Fl�4݆�aq\�Yh9֌MkM�FVf+��K5%���`�tͲ��p�l#�6WZW\M�Te�YTT�1�����	��q�9�qr�ql�:�@v��Mk3c1T
�Zd�,��� Ix�f�\渁jBh�k[,�Ÿ*�4")��Y,6�B:����&�ݎ��u������Ȱ���E�ܗDlƉ���-t�,!�n�ln�fi��Mұnd�d�P5���6�f�qn3�[R����*�Xݬ�(�3K�4��Yt��4�f%�**�J8�h`��L�Q3��A-��h4��q��LjA�˪�ؼ�ݢ�i���f�KJ��ee�	E��f4.�k���JSK1�O�xR�\��M��f�)4)�I���R����5)�c(Ъ�viKk k!n�c�����]s��;M�	J�IVPs5�n���Q�M�
��`Fy���ΙJ�����vQ7��B�$�b���;���]������D�[�\�d��lhA��E��q3+]��7@`ڠ�x���nڊ0���Bd�����!�e���R���	f�HQ˂�ӛ�[*��B�	CU/@%�b�]��ͳ�7��9�p��5;k�wQ��Q1XW$���������
�2�
�BR�#�:�,�&�Ī�F�h�v�-]{jh�6JQ�u�cp�1+fkkhF�dhM�LB㮚U���E��И��ғ.��E�J�@�6�ј�fb�a���^SM-K��2ڍ��m�V(G;@ڋv�]�A��Rkfl�3a�)�%_<�%<�QM�X�ZkTj�9D��.�L���V���pC��L�7l�-3�6f�0-͹k��\��*�. �}8���B^�8��Ι]�Y��� �����I�?	;��H����4���qe�E��l��Z�#@Gp�R/:���P1eĦu�� ��$b˩���)�@�slt)H҈]w�,MC��Mח]3c��B]L �`CJ���4�ɦ����^�����)`1��pR�cL'i�Y�`�sLP�t2�Ɠ�n5Վ�+R��+h��YIG��.�yb�dl`[�ԻZ���K��ޣ��d&V ]���/�u?e��P��[�.��TZ��K����4��%dņ��]/�|����>�Ow�n�� ��x�P���{��x�/���Fh����s.X"��=v7n���v��o[��D�e�=��,5q�o?=Q��ϑ�%ٌ����Z��o8�g��9�����9��\-i�/X8 �/#�l�V$>2��nZf�V'�W�\]���� w9_8pE�Ǆz퀻i��ӯ٩��2v���� �?��ݬ�f<u	\n7yp�W�b�Bn>�`���n�d��}I�Y�`����.��v��E��OՎ�[{���u�[l�G�f3^�7x�
�xg7�v�swoUTi�����u�h.�9�#%mL�� ��E��9K��k.M��^,��F��1�*��%9��ӻN��j�b�������mX��aDe����o���x �m���c5�zqUV"2����3>w���&n"����B;r&�&MKl6�@�O�&e�=���j�i����^�f�Z����^u�>w���=kO�=� �(��ЂRЈu��z���^��6�]o�.�x�/��_0pA}�=,�d��c����aW� z�8�p�]�����{��{���Z�{�).�f�vn �
�xv����]����bj�D�5'Aj�@;�n�8m楇5�j������C��w?�7�R_/�C��y��]��퀻����s�?�?E��+�.�<eַF+Ǖ7|o�\�� ��ý�d�����߿hC&rs0�unbu�8[���%�M�f�KZ�- �X
$&�O��E�F�S��?S�;��]�z=v�}uF�q|�).�f�vn ��8�.9�����A��H �.�����v���U=�5ݾ�a����u���jڳ��]_z!����E��v�AÈ��g��T���k�[z��8 ��z���a����t�\&�D8(�cM�Qhhw'������t�r�^���c
�UfZ��Q)<Nl�Si��g��Z�n3���jo8�1^�E=�� < �eˈ����ƪ�	��	�`� ��G��Q�Â.�e_31�F��Yl[�x���uF�s�pT��k�f�J�xW�jY^jdj_GT;���t�i��W� ����&�⃿T ��[9�8o5N��⮯��8�����������~�XK~ѹ1�l�Y��6sJ,�Q,ʈf�ZUņ��F)k���q�c$H�g&�A7z�n8m����RM�w3���fKTpN�{��c�a<����\q�qlz�ہwtz탂/�5�Y܎y~���;_�ʉU���IZ�vow�տ�v�l�Q{d��)dt�m��ɜ���]��`]��ɶ<bz���wƩz+��D?@>;�|��E��x����ݳ��Н���*Tm���pA7v����ky�%�8'nz�� ,��l�gA��S�"��b;-�R�P\�?G�v��찬�}�����
x��e~�c>"�Uס���.���*��dw�"% �(������_^�e/��v} @&m��Eۇ"ՠi�|��T��ip��D����I.�͜���w�U�A���ݳ�7v����w�mS�>���[��� ��R��l&�
�]��X��j��@V���޽��6~����߲6_~�>?XwZ�m�`����5k�v���Ɇx����A��w�G�S��ݴ��n����k�d4lOo��r5��6�jg۝��U�-Q�;w��X��3Oy�yZj�fDc{� ���A�p�"����7o�/��o�	������}
���s�q��Gkv�A7v��av�GwU�Dړ�� ���p g@��u���
�����;��li��(�����	�v�A76��Ao��h�5"\��w>�ɢ��]�)d����oX8 �]<nۼ`���ae;�m�e@��Љ�'��L��L%�4�k�� xю�d����ս��-*&%�;J6]zAj��a�ӭ��3[��c����U܈� @��]z�!�͸˦%�+vIa,�a����H��8IX9�sb���GM�붦��)k��v�-�)3�U�����kt#�1%�`�#�5sl��c�M�ۍ�K)�cZ�Ѩ�%�y�u�4(K���6�)	kQ�+�yp�h�e��,`��Z�Uů1��<�C14�+�s��Z�FcZ]J;�mt��e�X&��a7Z��)�����6��r_�P�ƌ��.�b"�գ���ÀT�k0�7�`�<!�A�m�� �0z���]��>����Lp\��$�;7���F��:.{:�_l�I�&��l� �v��ꚭݦ:x7j�7\)��{�>�
��v�0WW�/ ��pA���p��h9۹�7;�'�L��V�����r����,ؔ�Ǯ�w�|���K�
f�A7�F�� ݰpA�z��_PЗ�\�W�s�#�ǣ�m�򂷽1�n���vn�i����X�coM����y3�M_<_�g��휒����R�&t���~��s���E����G�7XA9Ñwq�ovz�s]�m�e����&���-"Xn�܂�+vi���j��i*X�m���i4`�����Ne��ڟ�pN�{��,���-�0�.:�!y��#�z��ۇ����`��{b�w[MXy9U�osmn��b���Q|K[�˻���.��-�ի`T5�yTl�OF��tx0��N8��O{}N�'�R�<�ɅPMB�/��TӗTn�"Tl}�_d Э"+@�P��q �J=�o?��������s���&�<Gk��n�X�(ݛ����5����0ofd{1�3+ӽ�9<�=P�hw����1#۬�8wQ�.��k��;�.�(�-P�]�w�N�����R�3����Ia���w�w�z��<P!��A�U'�`��#1�����@ ݰn��W�q�jhI'��5���s��ªo�vn ����A�����gwo�kC]w:�Zh�+Cd����c�ܭr�J�e��U2������\Ói�t�A� �l탏O��w8Wc5�V_
���#�nA�k�ޠڡ����Z��.���A ��ǈ7Z�������ɼ��c��L_��k�X/\�V�7�����6�sjzA����9tǳ8 �v�U�G����Ox8`��rSi��aB�ېm��S���b��>d9n]�xL��w��
�x�z�:<�@kƻ���瑟�����ϴp4 4����.�)�S (=S=g�t>�R��fe?ޏ0m��v� ����0�o���N��uT{1�}v���m�ց[|+��<?@'5��&��YZ�`�S�6�C�n�������!�M����)N3�ּ{�%9~��;5}t�\	�Lf�Z��Gt�6l��"��$xv�4�&Ig㲭p{l�a��!c.�m���&�+3U�U\��к��E?�/��!�UY�>�N_�����k!�*���i�ªY�vogH'4T�vu����3�Mݼ.���C
9#M6�-��������[cu�V�
���� �qS/�T��|=�6z_��o{��N�x�.���v�A7v�{3f`X�y��l�|��1�y6�<7xJ�����k���p�"��LG��f�L�g�͠#�m�VoctB�/K,�;7��O �n�y�y!�x�͍���'��u��i�(�|���U��>d{U�L<�� �y�ݥ|S�~���W�b���"]ވ杔�gԮ�]êjY��>���<	ZJEU(hG���}�����s�m��`��뻁�e
OH�XU�
������W7�x~5�{�E��x����=�Z�ܼo'��}Op1�n3k6�][@f^�Dt-�wV�ڥ�HK����_S�'�W�!���!�����gwo)��c�S[�t���pp�h2�j��#/�G�X��>�p�]��탂/Mgs�Fk�~�GNG��˟���Uvݳ�WzYg9ٸ�
��y��b�koo#�βX��ѯ�֯M� ����l(n�t�i�ysֲ����Y�����\�y����`��_8pEݿ�����x!�/�{(@��/���W���1v�:*Y��4��z飁��+X��ǡ�{�cEZ7�q��l�m_Zs�`�b������۳꼾�|�[6p%���]��%Zx��pn�����ɻ0}�z��ʩb��EPy�>�n���U^��U��9��hOc���9D�{Ŏ�9'� '�/����8p�7��#�4*�>�m2�]����	B%" P�KgwN��?�g�6[�}�D��f ��Gm�R2�q����*�k��[Ĥ#�j倬p��M�2���P��A��Xٴ2D�ب�v�PʃIX�i�][IZruX�j��d�Y�j�^V惖��L��f%�pݮ�(�1p��4BR�Z��QH��)0��Э�mL)��`tA�c�v�㳛�#�4�2���į:Zbf�۰���1%��ߞ������ᘚSk��%�$���l�	�����Z��U�Żc>�C�}��|���2{�]����?lV���!wab�o���d/oQ����؆A�ި������9����!�1��\U��g>�o@�2����z飄3{���l��tuCh������8�0<��`��E���v�u3:���93"���ڲ��
T���sv��x]��F�c6���x�[�����p��V��`.�,VM�����O8;lݲ1��{Q>�9�g�v�7o�7l�sm���#����Aݷ�0�R��
j����8;0�ÐE�@�� ݸ̺����_>o��{�䇞�a���lu�9�l����Y�ڕ�j�*���j�3��gר|�������=n�]����Wc�����Yvٮ��Ql7:��qR� U?��r	����Q�� ۻm.�`;�a{\���;���0�zsh��ss՞��{�tõtގ���-�Y�]nZ7ޅ?y�Eٲ�c'�^'MW��{�=� 	�B��:�e��<���~��}�{��VM���k �8r.��]1������g ��x ���v���ݼ@�nu�-l��6�:�����l����V�r�G��Q����7��v���vGs+Ĭ]�����;Epv��l�f�x�O o�2����j/X��gy��U��J�+`.�X�+�n�3��f��T�`�?��|�:ɾ���sX8 �������zQ�}�jy����~ҥ���;\djiaE):���U�1��9Q��lmJas���տ}'�-����{�9���n��lѤ�����m����.��V�֔�%�A���v����ݸ���6Mk�a;.�%�A�<|���
�n�Q\�.�5ٽ��?�w?��ֺ�.��N�Tn���=��������|i�.�1w�N�����C��=��/O����o����k�"�e�,�:��|d��cr�t�²���!��;�nE���=6̇:5v��x9&=�!�A4�͔���>ۨ��,Av?r�R
��7/��w��f��Wz���7�^�h^;�O=��ڮ���v�pL�g�.e![��8���=_��&<]��򛝷BI/)B��7=����J�4u�����*� H����e�K���[��:���稌��<{��O��n,����������.$����)Yy���f`�|̧��P7ϱ�:B����*{�<W�N%�hⱊ�Ƒ�b��X�i��e]�S�V"�H`�v�w]��z۷�D�A����_g�]��Ow��ݹA*�uY�[���+o�B�A�{�*\���SD7�=F{�O��vJ7<rix�����&J�rS����u���$��#��ݞT�i �o{���s}�f�+��{����z���v^����8�ȼj��k:>}�w�F3�]L�@���m͢|qg���{�{a��z�5[��9�}��=s�	��]���PV�D�|�vs>��`����%A�bgo'�S�blwō"{����k�`�;�9�S���s�^�]v�wI�>�{պ{�i���>>�Ծ�R�����wy�an���i��?`�h��a���˛O�l�����qn.�������b��I����{��v�����e�ѹs��T�Y5�uL���*��ԟi��Dayż�r�+6Z��xf�����c{�(ڱ|7�h���x�5�� 3/�,�8[� �Ls�T_��2Ī������2�$ ��E	�Y�vb+їsÁC��\�ܜ���]�!z["8G�/$��$�y\�܂�f�G%G0�D����
�"�w�'N�����iE�Rn~�r��<�Q.y'u�"��D�=nBs��I�9Eb���C�҅/�ӞO����Y�Rm{��K��K�9�K��q��
aL��#2"�D:[����.� �/<�;���J���' "q�x����좮K�s��^�s���*���&g�����ٝΟ8!�7v�2=����2y2�y��������m���Ȝ[)�;�;r*�E�H�_)ܓt ��h_=�S��*|��|��/1սH�9��Xw�<���� �9��oS<��lNS޸p����J�K,V6���N��'����DihV�ךם�{�����<�^��k�"���<���<@�p.�HK�eV���U�%_!|~Y�ڟ��䵶By�=e�;7x�k��}��1��.�����"���&x��p��9���g�*s�??���f��n��m���5�x�o8�?�L�JL��(.�!�e@�}sɳt�f�!�1�cՖ���nMg��ˮ�g�R�\;mT+K4��B`��18r� ��8��W� u�M��cš��Y���QY}��-y���˭a�Z�2���2Ŝ���&�z7@{oi�g̓K��x�'z�pvn ��pA�$�`8�;���h���L�޳��w�$��d��S-�e�F���}'9Z	F���e��f�	��#y�I���8!&�t��������Ӷ��A�p����]��l���?�X9 j���s;1��s�{~�F���sf'0x��	̓�����Rɮf�B����j��cJ4gZov�δ�g���E��9޲w�,��9�z�"�Qi�2�ã^�{n����"�˟��Oʞ>a%�r�a�g�������'�ٸ;7Nkx�ĲL �L6kU��M�����0� -��4�&���˻g��T�/0��ʶݜ��J)\��o����<�=��	�`�98�y�mm͎mě�=,G5ٸ�y��;��!���H&�܃�b�Dv��P�1fJg���i��s8���9�H��R�=�;w�۬���y��m6�D5�;��y�T�>9��&^ ��	��]e�`f��1Q�\#(Na����}��� ���$8�`�b������{t��Cz��� ?�o=�]X;��pg��g37 AS8.����r�9�g �L��m�7l�]�pRa������bld���y�H��R�=�;s��!s9�N�7�M�O1}��FCAraձ��Ν�8�"�l�M�I�P�v�KᬷM�3r�w����`꽸Wi������
dI��0�"�<��n`�i���,���=ʫ@��a���x�"8�8�^m�X�Ɍ���.؆5�	��E�SZ����gTm�˻�Il��XP�z�J׮4W7Iqc�U�f��*�C ꮁv�2�ƌ��b�Y��I�rq�H�G`��2lh�:3r��YsS���+�\:�"D�J�[�ط�.Q��Vԛ��n�4�f�B9�	�u[L��ۮ��4k4Hk�]flIB[e��'ϓ�	�.ƫW�����u��!e!e�.�`��U�2�>{o��
�pA�M �Rm�4����2��m��Ǟ�^�$Thi�<�x�����$X�H��9}w�N����F˿���[s`��M��V���A*�����I����A��x���L�_3��Os ���R`�!&صpn+����j���ȫੲ;Hv���sX?�+�9	8w�O��I��b����(�h:��=�kH ���d�C��4̡=�ہf�	�`�wtT"2L�"����'�\[C�n�8 ��J���9ð����̭��VvZn�,�f��L���r�9�j��o �����/~�8�A'��	H�Nl�Iq]���K&m٦�@��4n*5�I���-������I���[^]�S�W���!ۜd�\d���X8��9;����
L&�
��}�5�3������x����^!ݝ
��cd���m2���B|�3�N���Ǫn!��[����fF���;.�֍���G],����>x�Kě�;�轨���{ޗQ����s��iq��h�B��m��q�pE�)0ؓ��-z6z�w�u�,q�rV�Æε�1�d�=k/w�Y[1��啀��9��Jo?s��L��
L����oxB���wzj�V���`��2ns�P3s����N~ �8pﭷ^�An�k6��f�p�m	��M,��60�row��P ��pA����Lj�wsi�lSi$�q�'�c�cLJ���,��� ����	$�ZL�@���c��;3�vG��l(-�6�bj3+�٠�։��ÓZ,KW�T��v0pA�@�.�?��q��r�5�MSaf�7㌾�U7
Ӻ��B���pA)3��9���#uo�6e��l,��ö�]�.�|��������`�%s���!*L�וN��]���f{�2E�eͭc$CkX]u���� �l�=/�"f;j)�X�)��n=�H��3��=�����I?C���C�6��ۄ����O3��dưC�}��Ǚ�}�	�hh���ߎ���*���<7� �������&A�]��.�l�zCa]Y3��;���"ݼ�?�ZZ��־	��,�f�A�g[�n�y]P��c������|E�r��I��.Y�-[J`l���O�Ư��#��f�`;9Ð���BO��Ƶ������S���;�h�!��K����tѺ!�¹%-��bƑ��S�#/���}�7Ok8 �e����%&��k�d��$[��,��3s�O��S0�[�6�	8��7l�����To�6[ϸ��蝋�|UXY��� �ͻ��?�MՕ&��9`��ފ`:���&�
N�dr�Q!�WO�W3�\H*�ʲ7Hv���A�p�!'�8)3����7���\��o��8 �Rg�
��z�y�H�Y���A+�ǫ0�у�����Vz�0�3��T�]_^�D�k��e���7n�l#9,ni��SZ�,��Kdȵ�ebZ1���a����(��R�ōw�>���� �Y:.����y��ֺpL&�
N�$rI�����f&TN�C�����NFq�)��,�f�&m�w��
L��2rb�
�"�C7[�.�3�Ն�dң��5��.a�]��T��������#c`�l��0E��I���`�7��5tJ-{�Y�;0<�n��d�aD�I�?�O�&JM�kX��gC4�G>���`*���l�l�M$g��fn���A\?�L7n<7]�i.�1������v�� ��9	8��g3QB몓lν&���&��9���Ӎ��<�&p%&rg��^1�n&-郂'�&$�Hk���]�_yVGmy�C�`/�b_����j�XpX�_��|0	
��$_/��_r�䇗�2�bV�V�T�FvΆf�	V��;o�����Z�0���v.��q)�(ܟ�q A�Ѹ��Q˽z����U�,R�͛4a��S��RT��j��te^�i�"KI�fw�+� �m�q��}޾�nE���g�<�R\�c%��l�t+��.��� encm-%����7h0�
.ΰ�b-n��m"�iI�����Z�.�5kE{V:�蘎I��]lv��8\�,5��%Q�Z�kV��LCM��r2�f��YEfݵ���3ѫ2�U�1��Vi�B�H�bV�15�]R�[a	ilFk�I�lc�\,���|����+-��5m3s�T �t{-m&�kK1�Jm��3bR������@���8��p���8$����T�74`�����g37{�k.d3ߘ�7�<��-��䵬e�kgZ�X�]���ѱ@�0�öe]�u�"��K#���P��s�v�#���F��彠޳��sY����z<n��&���)dz9��ͪ��9R�i�<n����ۇ)0Rq�]�w'��5vs�/n;
u�r.�?�o8�&֌ؙ=X��f�Iq����n���;�-l��m @&���|w�����[p����4��gu�Yk�%��C�8>7�|3�?�I�����SQ��4q��M��z��:�f�)�S��rِ�5mT,1]�\��+�L��!�� �/}���_W�?V�����*��G�3{={<�rT>�;ɖ�u��=8;]��$<w�gc����)��6i4L��]S�h�������ߵk�' �k�|�YIu��T�gDޗwf�C:S��b�D8X�y���=��hZD�(JB�+����B����-��������5���A3������0i�֏`@�ט,h׬Eۇ&I�!�9bz�H����]J�*�f�F��8�FsfI��/���k������U��+w ���U-����Tι������v��G,��K ��y�v�Uۇ�dķbw����YޯE���v��,wbt�f�7F3���rR?�MU�1n_�b�Tu��C�w�\0f0�SmjX��Z%�a(��WGV\�ژf\�=Ͻ~N�`� �p�&��������yE�݄R�� ��ʷ��5�3�k0��a�Æa ?�I��&JM�c����9,��o��p �m�+e�6yI�\��f��;n��<cJ��)
lX6F��H���kY3��YB����
��K�pf*�����2�cS:�͑�M=}����oh7;݋u�Z������/��(���1v�����r{Op-@ĉIBo����8}؝=�Y����K9y�����부E�9Ӭ̻ornp��v�9�8~}���W(idv�_�^0I_W.��pB���������mn�����)4�J��B��>�	��j��Bi�j�c��zpc�`��x�}��kX/;o}����MAݝ�������pt`��k�aC&5-��bdV�f���-�;>�C�O�r{Ѐ�`�X�BR&<�zM.M�:�̲��f������e�g�����g��	3��R`�m���])�����`��z��W69�Y������� �8pJDN,�ܗꧦ0;�M�5��|s��A	?��&&x��9+iɩj��Bi֣��p>�o�ێ����8^ �q�/C�p�#R�v뀵�!'��\��,u�]̺��wp2X��� �m���1���}���pыg�,��E<t'��VtS�B�]7~����0�ٔ���~7vn�P���+n�֟vH�*����W/����	Ă@� x�#B4�'�����g��1�c1L���)0����^�q���r��%��cn�]����>�p��$��_>�O��������{o�Q��g+�;KE&�(gk��	���l��]/f�Ōx��}B����W�L��#��Rg �������z�α4��,޵UՑUڳ�~��{�9��!'$���&��>l��3�^7���->U,�֜u�s.�9�����~Y���_		�v�\�a��/�rI��	�q�oe.��ˉ15��/Ai|Xݤ;pp|s9��J|����Rg ��Qp�Fu6�k_���r�8�T�l�Db�4��,�`��}�2w��ޘ艭�O[ �Ð���?����:�3�x�l���F�Y������i��]w2�s���A1��w7���-k��ۇ�힞���:yyy�o�0m���hI��*�5�ّf�7�X�8ʏ��[�NL�jO�'��c��Z7� {5��i���z���%U弋v�I�<go��W��էXT�wP�a���<$��k�=��g��>S���1>ay*��-�<��g�=����O{�xIzѷ��&�ݠtZ�o�Q���w���LQz�]�o��2{Ow,��5ݏ������}��>(:Vwg��;=�7������-����;�k��gx�1���v-J�z%�g����#ȡw	��7t@��N�T_����v'�ŵv�Nr��=������G])��W�J��?��w��{�n�^~�x鎣�x�f͞�&ٸ������.{��\���h�3�<(<��nA��f���_��i�c��DN_������Vs>�αO��C�9��5�xv�����n��wʭ�!z�x;N��FW��dT4z=#δˋW�6��od��V�Ɗ�m��m[]�*�'�a�����o�G����y��s{��\#�Œ{��ub���5�ٶ�H�k�8�W	^9���d3_"�ܾX�G��|2�=�<��U\�U�3��=�#VU�_,��ͻ����gu�z���;}�\�ڔ�H��~�--��a�o���Oo�x���:�:�Y����6�ymه��â�r۶x�z8�D:��W�<钡�+���oed��-����6�^��}}ڄ9(7�������]��	��|o���0sh�>���ǻ9m�8���;����p}�0�"~����ތ��T�����ה)�Ht&��¹`z�#�t��q�kp�6������t�I*h��w��/{��>�Қ/����'��ۺS=
����|�Y$��<=�=�^��-�R�o��iv��r+����<y����{��č�SB,>������tr��:@}N9$*!/��Uy���+�E�/���=���y�*�>c��r�rnw�^|��=D��vz������9����y	�E7��t(NU�)�N	m�%�t-��J&��,��9ݓz�<��TEQ�eDξ�!g�����z�ʧE�<�P�V��r/D��iȇ?�V�в�RhY�U{>�ŅG��̴z��d�޺m,{�p���}ם�݉TUv��I	��
N}�$��˅ܛ��(�]N�.�{�P�^��	����	�6��N>O_?-�ͦ��:�oD�G��w�
���@J������5�k��59���Lָh٪(��Yk�(E3�Ү���+�IpB.U�u:�l7Cv�͘;M�+�����-ٮ���e��7�.�y�-0Pҝ�Ԕ����Z\:if@v�&�GD9�m�F3l�M��k�RK��̮�R�c.6q�Ƃٚ�lk��Q���-����,ɪ͈��&��ܺԦ��E�&�(�5U�3��]��Ѧ6,4.��X�IM������+asC&2�ʋB�Y��7:=v�`Mb�z����12�YI��e�b�tp���:�SFґ� sq��(�	�!M����J�ʄ,%qi��4+Va�ش�\m��\A�ݵ�&��e��6��f�f���)\D�jb�j�j]��2�iV��2�5D����LaKn���������:�ݫ�l�� [���B1��JSe֋�&���&�H����T(����ڑ�m)B��i�V�r�{gU����h�D�^�b˭�Uce�Ku��*JB.���N�F���@�mIY��7�2�4�WB�����cD2\�A"b�.䩩mMc��b�����b��n,���X,&�A�����K�����%����aZ@YkmCmW;K�b�xA.N�	���������^�^F���h:�Pj�.��R��Kutڂֶ�ⵠ���4
��P7R�h9����!�6�2a�&�1a-ń`�형�n�V�ɼs5��jnr]	
�U�6mFҐe�vB�RĚ��Φ̎�i��� ��9;�X����5�Ye���ж9WV�eк��i^L6]�(�,ݯ1���+jr�ҤWS�D8B<�v#m33�n�	�P�q=e�i��"�f����sā]�6�Wi0kl!�t��k2�Íl�u�HRQ�JTK�����+��69h��ڰ+f�:%����H�K��cAc��h�8�&�^T,�||���k�f�T��D�޺W���A)���s�lؾ"���N�h��X���}P��-���ځ���U�����o!eVYA1k���2�Su�Vb�F]�l�e��2[Y���v2s3�a&�f`Ĵju%��"`0ܩl�"�I�ۺ��&�J�Ds.�ö��=Ublbn�R�5!f#P SD����k��b2�6��lѻ��:.u0�ZfZ�[��ظ���5��4n��塀�B�&�����fɞ�5�"W�����gF�ni]1���f4Ȁ��G"\�5��ZѰfU�Y|���_W��><�?�>���L
N9�37y[ކi|Xۤ;7��r�|����l
b:%���p/%�R9I�$�;MW��E��b���o8=��ʙ:ڇ|\i:�<7	�`� ��r|RasS��2m]�%��뜙�Z�I��H�k&cZía��x�n�4��])���n\˩�fn ��s����Rg ����orؓ��%�0�����'�]�������b��!۟�8BrZ�ë�S��������������:�BC��N���9��5��M���޳�']G�f�*X8 ޸p
L��n�&�}7Vv������\\�6n�1T1P�p����JR�]y)�2�g1������^��\������	;���x�˹����]Ns3q�=5t��mo-d�p�1���sٍ �n�8 ��L�}�w9�
�.��p�n�'�2oA�}M���:����'s`^��M�t��b����zk�,V�-�� K�̺w2��p#Ā#C�)24�3�d��� ݸq��>��[��g9xݤ;pp@7l}|��IRw�M%��_����p���)8	4���^���+v�����z�<9�܂�e, ���&!'�.�8��Ʒm�na ����HS��M�U���pr�˙u9^�v�	�g�xD��A��'�������Ma0pBL�&�].-ĉ�+X����Q��31�H/�7l�	$���$�}[����2�^��+�1!ʇխ\.\3���[ل��	��r�Z:,G7ۺ��L�n�}���/�Rg>�&}ԩ�m3Mo:O=G�3w�P�o��>y=M�;�^"8�&[]��F��$kYrE�`�G��ʵ���S�<�o=s��uK�kN�칗S���A9,����pRi�k����eۃ����c��fְu���Mpsu?;�	��!\�T36j�^� \|��͋���b�`�`hY�1���_���T���H���;�E�Pk�������w���l׿s4�)L� L�ERRSCǝ������동�f[v�_�lE�$��BNM ����u��F*����?��p|�8��iԟ������\�pD(l���	�m��}Z��	8pJL�'KsC-�w�5?�k��f����5����3��q�&��㯛��;k�w����]�3���8v.�j��ؠISVNVt��I��۳0��ϓ�-��8���O�L���!'6�7z���3-�Hv��z��d,m`��58p����d�r�9�&��K���!Vfz���3)"�i�'J�[��fn ��pO��o$� 6W�lf�^�p6�H+X9'	8��P�͗Z؍�J�%S=S�sOs���A�w }��pRg �����M �<���3a�c?���`o+�;�Z��Fe���U��[�i�&�,�b�T�U���{�\��+���į��"3R�ۓuw��-Iڻ�\=���+�Z$�I҉̲�e<ő)�+Z��>$��9��8Es���W��|��h�������x���fS/�zpQ�gUiQ:WȷI��� �z��R`���$:��f��=�`hP��q����b�jY�S4���*a�BY��E�����	�R��u�rp��'����dvWUT�Z���fn(�̘��j����0y|�̥�W�X~��`��C�Yd�y����m����p�;x��:H̶�!ۜU�r/X8!)<f��4�{��~;�����'�Rg ����/1�q�Ԣ�j!��[$�fn� ��A�p��?�$$��BM��׽��v>�8"����?�\Ү��骞X�\�37��mg"uy4�^m�X=���pBL� ����I��<R`˲�ZaV��3ݮ�wo;��C���n��w���z��I������=!���CD4��3�"o�Qnm�᪏x?�SU�i"ʑ��K.d��k�p\�O�1e���s�bzȸJ����-�}�G[Ws8:�xw���V�{OuU%%SS�������u��8rWL֐��K��t�l��<谥y2�ash�vS[5��"�6m���YtXgl���{�-�che�ض�k��1*ha2ޭ׈뵻1$�m(�4��b�[	��غ�5D�B��D�C�q��b,1a�X�\������@�1f5f��&e�]�&�%`�rlL����ie ۣ�l�`!6�3
P��0S�M6B@��|������3Y���Ѭ.A]��:kAu��w+��+��a;��w�;��Є�8)3��Rg<�O�����I����ѕW�Q�x�	:\89����!'����mð�����)�뮙��5�k3w�>1���o7��&m�F,L�:Z���� ��I��	 �⇧T����%⩺ꬪ�$]�o��i0rZ�Q�S��SzN�k���Dky�X�<|�?�q"���iG9~����d�q^`�!�������*�FL��R�������p�%v�ֶD��J�TTV��k!��l�蚞X��s���&9��5���@&��]�y�����xO4'���n���^��ң�v��s5lZ�h4�iB��fU�Y"}�u�=��q|X^8r�.A'�ڳ�u���p�i��7:�Ai�]+l��A���B����ȇo2M �
L�"&��8�/�m��(�Y.���f�<+h)�a��e���s��#���'K/�Ị�"ъf9.R������{�'�>�%%ì�=��8�Dx�߼pqΤ��j��S��<9����AZ��L,wqצ.��E�����f�@9lv�%/����y˓���ݩn�{��YF�sY�����7��Rg�?�I��j�us�эԑo�`0�X�� ���l彣��X�-�H.ÁV��K����tP!�P"m���o8)7���'��*`!Ρ'u�
��L��rAn����N������I��
N'�$�mlf����x,��
��˪���qYSKj��f�E�
m��s��\�x��FN{��7`˧6O7�,y���E�ʕ��M�S�(��s3q��yD���95��T�s�����I�$��y�3�Z�yzs�������Vv�J(v&q�C��[ ��Â���*�lx��̹��;�E�8r�YrZ�3�au���5���V��Ҩ&�bI�M�:&��]���N_�j"߼@7�Vo� C�������5��x�w˸6י��K�ȫ�Cv��9��	 G�oW��~�i�C7�x37�����Z��LBN@���wI� cO
x��� x�R����I��JVl���YF�s����F�wK�,����g���zAI��AIÂ�	N���O�X�w�yzK{G%;���%��[/�9	3x�	?�d���@�4X���fj����J�`h(Hl�vZ�`7#���iwk�r��f�-� ��w����r�8 �i3�rI���K�sC���Lnҕt\C2ժ�q�W�Nn,Y��,	,#Eȑ���]��NJ�.�?����r�dv@���5s����	�9�@��v.���-��y��z%�8�'�	0pR`���pP�[�\D����5:�������U�p7���?�o=y�7�C�Y�gi��3�_!!_B��zt(l�K�X��<��A���@7���n���������`tI�e���(>塇�]��O|!�=��Ḹ�*����j�q�e��z�{ǤƑGwپ>����zl`��`��׼����y�#ZɒAI��]�`vL���Z�j�ϣ�uGVI���f�=,� ���?� �v��y��}��Z?0K@0�T��X�)���b�	��g$���H��u�c�O��g����W?��I'�}�Ǔ�ԛv�k�o@+���q�y�j\8"����?�y�g���Fms�~���<��
�x�T��L4�u�~��������^�l�������'!�e�p��$��:MhJ��U*����Y&�s���}��;��&pA)7�ib���ܦ�?�&� ��kn��N�^�XѺA�pJ�D{��7c�e�*����p?��8	4�M&r
O�)7E^Q��g5��n�i��x������㩃���Y0p)8�w[��?/��Y����uv���?_5����W�t�K�W�`1���^��d�N,2[n���}���⏵᪝��}U�����@��[KT!�DA0��=e�eE��Xk��L����c5���#\[�n!,9����n��F�B��p��͓�Yq�]��R,�i�&�Ձ�U.)�Y����c��1�#�gV�Pmت�j�%l���vF��I��)CcTwZ�W�P���l�sy`�1�<׏>��w��K�6�4`�'Y���+	�csCMH��7p�u�L\E#�p�(������)��JF�'ԃ��6��L8��F ��Ŧql0J��ݙ3������
���8$�����U��":��$��s3p!#�����uDTm��4u8���c,kX�D��,vyߢ��0v��Ek=������Τ_IX��E7l�8r)cl��YS~QO�9l�j��!'^i�g �ŷq��ӗ�Pl\��Ľ\��c�����������L��� ��8�%��ۚ���avGKx8$�p�7�t���'�:�M�Ώ;�@=-�d'���z�����r	�g!&�9	0q�k���Oc��Hj��x�}6�Ž�n�Sr�[Oi��7l������<��T�cnw�������V�gjل��cB�EGkZrRRnZ�)Yv�E��aZ0/�P������.!�_7a&q�`�ݳ���N�1/Y-��f�����x:��V��=����?�`��6�3S�
"��ڋ�*5ܲ���[���_�}������{�=�0Z!�퇕��K��S�s}���#�O��6|���V�g"Med	Ƶ����|>R?�|�d���r�Q�$ڜ�f�=L�Gs��I�4�����;p��ox��?�7��I��>I����{�Gi?�jU��WC �i� �y�탑e�ɫ��	
���3e��:>��\yɻw �&q�S2�iz�m��<7@:�9B4m�v��۔貭�����p�0r�p�!-d�c=U+���ܽ�M��ܱ���f`6[�=��)7��&��������-�\�0Ì!��H��AI���A�ݛ����6T0Z҅Q�3����H�.a�-�p��I�BN3/s��u��*�wH5����9��s{S�����9I���9WϮl�=l:������Ay�F�[nL�G?K��7
��<�o�3[�!#標:w\������'!� ��r.�9	0	0�������;{|p������������V�֫V.�,(f��z�~	
!]����W�}%��}79��2��E������%���ǜ�c|�}a�[��}^\u1㸳ܽ��j{Q�.<a�Rg��sݜ��O�Ś�'� w<�4z�k���S�c��Lj���=�Z������,N1@S���)v�����{R�ĸA]�w�E�fr�0{yE�3����_{{P��]<���yw�����q'�;r/s�h��[yv�O
�g�*��� ���z�A�W�f,�	Z-�h{Wu!Q�ѣ!���y���(�Y��;Ӣ]nn�l�9V���9$���p������Wn5�e*�#��wa�W�XL�߆�z}�\���/�8!���2�={��c��^�8\�\Y�;�c���p7��9"������e"�[��k�~$�\%o<r�����vG#���ou��w��+����V���Q���p���>e<�ĭy<�]�r���=�4����w�Rt-���I��\��xvG��<�9>�y�d��Aކ(����ɩx�r[�WUt�*"s,ACa�����9,[8�W�=���[���b�}���ۓdŽ��u��m��Қ�C���]����γz���G3�_`'�k9���� 3V@��L���S��{�?n;��>i�q�b�ߪ������T���9t�h�t�Qz���/*{�w7#�!�(��ϲu�^���只�^�������Y������p�wpV˲�@����}���Zo���{[�n��O��y�-8bbf]s[�YR�g��\���y޷g���$�SD���|G� �_'�"]�8��B+u�'s�e��L@�5���ܖ�t�����D��1*��ZGx�ϒs���r)̮ku A��5v�@���0���=� ��2��f�q�{��ot�
p8D�5X&��$������ĥ% UX�RJ���[�ed��g���<͖-�^|KM��!Hb��{\,��.�9巏^NK�w��#ŉJ��+�9�G�\��#�%̼�sn�s�r4S����X��7wDC�q�!)P,W��MF�,N-�������s���]���w2��zN�֔���8�p�kƴ��V^��Bޥ����! �Y�y,*""vU������ݮٵm׈� ��1�:��*����z��Bª���	)m��z&�:{s���*)�L$/��Ϲ�$��=�x]u�v����X�*�fo�����w���I��Rg��P�������KN��l0�/\֒`��2�[�WZ����i�q
�ȑyK`f����xK&��w������v� ݷ�v�I����|�cz�1��i��)�I��l���6���oX3��d�k�k&�y��a��@�^Ի�yaiem��4p�K@�@�&м�B�r��lCD*5�;���g���_� ����D8�̸F��N�,dʳ���hoQ���#�6u�M�?�X��	I��v�&C�VՈ�h�6+�/��p�:2WZ����w�s�
6\���BT�� f@���M�9�`+HE�&�v��Û|���i�4ET5��pb�K� ��w�(������8���/�7l��r�mÑ��&D?�z�:�v��;*�fn ����+x�=�M���������q|b]5�[�� m��Wbi�(ͤԱ��C�ǻ��ޗf�o{���Xvk��3G(����X��-���Zݳ����{@��=�z�H��x�ӃV3�����8r�%�T
Z�����p�5��K�Ofs�k����c�!'�7�?�Ϟ����f��F"km�Ae����-+%*2�n`�3�(hF覱��.�ف}}}B�<�8`����$+�>�|���D]�ˏGs�pb�=�
^�6�Sd;>�p�[
.!'E&�(��.}��"��F���a���S�Ք�9������[��fS�h���oӭ~#�oF�	0��.AI�fɐ�ǧ�5�ym�ir�d�g;�s�Q�����$�!����Zh ���g��k��E5��;�L���N�b)�;�������:�K�h�J�+E�:\����BN��Q�
!Ix�x�3�e��E�[Mb����k��f�	�g �5��&r	I��tϥ2-��Lq4#2�`&��+W�n�3s�����r�G��l�!Y�V(Ќ��T���zc/�r2���wϴ�.�@��;i�4Kʖ�clݠP�f����t:�錆�T�k���-���f�`��WF�2�u���"���^a�,����M�l3XLainƕ��J����ґ�s���fU��n�X"D�����5�[3ju	B���9���HB�[\6X�����t�B�s*����1�t^�!�k��˄�i[����"�ĩ��CJ���{���X
`�����b.�re3$pѫ�lg�ٯg��>M߳���	s ��x���';�n��\����Wy��Gq��Nx�)8r+Ι$ޒ�8uԸ�h|��@9L�׍�a�������vm[��#mÂ�<�49p��v��у�Ñ)܂N�\���!&�Ȉ|�|n���S�-d�|��7Y��w�A=,����4�)3��Y���kr��Vto3�XA��>n�&����˙���w�ppAFˏ�-xS�gg��M��c"�&��L�"�.II���;jڗ��m�oz��V���Ց�������A�"��
N+*8t�!��}�f�X�	����.��(�ckeԪ��Y��\̓E�6��]#���g�\�G��V�rw�L�x�Um��Lc���f�}�t�%��]���l!��� ���Q��&� ��qG�NK��&���׻O�@�d�»��vX(�|�#�4��oc ���������xym�B6b�eT�ws�YX�/���E�F	�Y�����V�$�����gdݟ��M˙����2��g�����E��o�ލk!���A=�� �Dw��퀹d��޵��Rs�r,sC�SCVE��ň�v�9mÂ�.A	8q�a��T�liR�t9�邈9��7K��dC��U���Dc���f�A���F�SA��+��e^�
�r	�o"����'QG�kʈ�yi!���)�=�)�s[��\<ɇfϖ��BO���0b�-?��t�y�?��@��e�@&.�]�F��s����Jg����hB�ao��{�����;O�?1	
_"B�}�땥_=��������0�2xlQ0�m��x����(� ��?�	;�E��E��7i�g�0N��M�8��WqktC`���wpA=l����1����6#3�- �]�z�� $�E ��m�w��ӳ�}�GљWƯh�;L����V뵙���Lǻ�M{���<�i2C���l;��վ�l�p{f�ݩ����ѯO�u3;oL��V���x���
�>��v����|�.A\9	;��ȇ&r3��-/[m�ۍd85lM>��p�qM-]�[��0 ��4ɷ�X���ŝ:\��BO��.A'Iɭc�v���sխd8���z�]g37�����&r)3�����I���9���pq0i�H���`�ܺ�"֚S��ηEE�\%s�����<���߿����E8	8q��F��Tu�k9|��y��D��H�3�� "���Fۇ�	�Ro9I��g���R��k`��g �Zѝ�uD�to9m[�`N�9 ���LK���[.�L8)���x��)8r?�O��j�:�Ims�e�8{ݳ���9��A�g �?��8 ��9	3��ӓ`���S>��`�$��n]�]4�e��̻���g$��������;j{�Ǭ�{���;�K� ��q��~����Uۺ���&��w��o{������P:-0�k�J
��U����{��Cp�|n?��ݯ�7l���?�)?���*ca��$�3�_v��tLVl������>!&�$���bl1���7Qe����8lsI��	n�1� ���o-����qf[��CMi�2�ϒ% `S�&9����	?�;U\;�ݾhw�u�[��+y�b�3�f�s�6R�bi�7�i ��9#s/�A�,�>6�8���2��u.SO�^�/�˃�n�8�Â�J˗|U��;�*�.����ԙȪ`(��4�Y2�5G'�}0C=P1]�0?f-��N���`��
88��K=OV�8h�Z��Fc��dC�b�Ƿo���M�kw� �7�-V��)F�rELo�;��"m��Xìk��c3kX˫U�KfM��
����Q��SS�^�3�ɇf˜�az�Ȼw� �;	�D��{�c��ou�v)f�7ݪ�����F"���5���@�sBT&��!�f6��4aʴ^#k^q�-{��f+[ͫj���M*%�� �	��Z9�KD\a�b��hM�AQ�]h%���%�-Pv����*����]3Z���2�0Pi�1&1+)k��C��%�[5]1u��:B���ԗ6�c?�>b�s^`&�ɨ�Q/l��̎V�z�",�6jl%,�ʶ�t�j�g9��B����Ũ�z�׍�*���q�]�R�Q�Z��i��+����&�3MB��'��-�����,��.�����L�r�f�:]��
®��~)��}���aRg>I�Gfر�@������Ż�:	�l�a5sw�#�6��p�pII��N�		3��k�h���Q�D'���o+P�w{��|y��[q�0r�%<Yd�/ϝk�������
�E&I���v���*^+_�òG�]��NY{l��.	m�\��	;���`�&pj�eL�e�dS?)��m�;�G�y�)g�ͻ�]Gc�w�����"pδ��S&��������n��p��6\z#rD�8�n!j��C��j�nm��e�M�;7	�g �q�d�ϡ2���`������#u)�iփ�l��X����.S	�G]uNc� �8x��K�z���Ek�\����to{��nz��fw�s�7���ι�]?\��j\9�?�L�pRg�9 0Ǚ��M���g� Z�U:ç^<z�8P��*��zߜ2vj����$8g��\��\��R��;��!�"�BF%���1��q��u3�܅�/t*m���w��G&�(��jhS��:V.\�Ȯwǎ� ���	7�2 ���Hr/���÷2��g ��{aہ췴�Rg�?��,�0�Z����9��>t��F����$��v]�멋��tٝ�\�}ծ.s!ߚ��	�&�<�m ��r�����/-�c<k[qufF����,G;n0�97��$���᭽��~�����Y2�ք45����Ya�QC6�Wî,u
��h\ɿ'�>���:�ى����z|"�z�C�6��3�f󝛼C(����l{yoi��s���af�7ly��E�(�-7R\��<p�r��˫l��7M��e�	���0��˓;6�M����i!��`�`�g!C����{٦�����J�H����.��y3��=e�]�݃�UE��ܾy{� u�����9~��ը��7�u��ư�ӹ���{�a�n�l�`�N~O~WL�-���f�-������(��$�����>[�ȶ�X�}I������Ֆ�����frM�K7N�8#�z���ҘCóܐN&���7�G�0D�ȣ�SX;}����&/��[��np�k��2��� ��Ú�B��A���K&���*$2�mF�#4�7E˳��n�#�e� �d��V�-�{�~� Գ�A�|�$�8��B�KE��k�Y�1n`�1��YN�/
�'l��IÂw�(��!k�(b��;��l!�w+B64�a�|�������a��n�0�����^����Ě������X�l����O�:���-E��s�^�M¬n��̸?��~`��w�	��M�z�ⷔ�t��<W�����}��.��8wK7,G�A�g�h�����L�*+�_ȶu���z ��
���t�7%/���f*��탴��z�n�+�p0{ߏE�Ւ#}��F��%jՖ#Zɖ4�^Sup��g!���!�R;��dK,��� ����5���7��&ŽT�ζ�:����P��ͨ���:�`�1&�gA��Mk�)P�X�8�,��{��Q�����S�����N/���z&�Wz���̻��Zo'P���?��#-��[�Rj��f���m�M��r�����9m��NlI�'������0�IE�l�=[��A�p|GT�&Ο:N���(����3Q�e�hr�7�-YVm�{��8 �u�q�-?!iC(����[�z�� ࣅ� ���d����ʭ����2��.C]�C���V�{m����mDv�B6C��Uf��ծ�ѥ��V��2��Z���9n`c͸���K� ���kY8[n��9p�������������{|�vVu)�����Pm��d�٘�5���姳d�X=}�:�������o%�`�V���{���NM\��7�3� f��#i�9�5C��^����6�]% ������<�E��׼򧋲�C}�,ܛ�s�/(�`0;N)Z���������n{�8��{t�g��t�+��z��&-^��>�l�Y������5�����٭n��J�I9�Q���^Z��,��~���o�YQY끋���?j~kV�j`���w=x����J�2^�y��騟7������Ǘ{Ц{"`���S�q9����c�/��{F�z�v�Ӱ$;�aL3^\��'#�>ؽ��Y��;�=��e��8F���,;�]'�����p���d�^ ���|Ͼ��z��y�y�Qa�i�����ۺ����yw�w���B{�{RKzh��,]����>�)�W��[��S=���rm�[㻏�}�<]�6{U���s�/y�T�Dp����I�7�{��nn�oj�uOiy*|��@,�����ͽ��C�õ�<�������${->k2��^��P����*�k�'�p�~�z��@�� ���~{��K�ޫ��}������g��ݞ�I������i[FL(��?z���w˔��:g"�����ݛƟq��qxg�z��Ǿ��y_+6��%f��et�|}��<{A<�mMO������gc�:	r;��?#��o<��.�g���n%Q.��Ȑ�xS% ��I�`�D�ް-�M�5�5�Q��>3��q�t�z|0h#`f�&�Vj6*����lȌ������
���xkA�Ժ�P.�:�V��1�!拂��u�%r���JM͖T��FYZ�Xc��Y��FT��w��}2�KȨ�����(�Mz���N�tS眧�y't.���+����q�7WD(\�F��I�w�C�9p�Z;���y;�e��+�E�^��Gsq�ێVe :�Lu��1^����e��,�w�W̏�#�ݜ��ATQvR��vVqe�j$�)BR0ú�%T�"	k3�8�KIs�-��+R�J�3	t�)"���غ��ۏ{�e\�H�!�<��E2)�T&r�|�T^q���u�B�fm���yլ�����D*j�tp��ϨPPE�UQ����e�(��=KB�� ������	� �$���܋$AMJ���r����YUY���idU&��ARQ��M-%�B*�X_�����Xf��)̡�f,�f��u
�&2ոJ�f[d*ff�te�l��9��͇���3hS7L��R\h-U���	���$4�M���#�Xh5��apXƵ [��f�*MVgb�WLf����h
�<�ǭ�`��h�1څ�Uc-իl#�X0L�����u�h����b�k@\��b�3�;;
�+*陱u�6�.���p���JMISZ����ۂ�K2v���k ۆK���qj��n��X�Â(�h�R�;.Ƅh��Fb[�B�6m1SR���n�ʨ��X9��ƗX�e*[i1[6� ��d�85؆�`�u����t�ʥ��#��+K�l��l)����6e�z�b�imIfQS(��6X�ű_��{�M���(@1��Yi�nF�l��M �MvX���u��Ff�ɒ54��b�Vg`���n,�b��2�jX��@�%ƅ5�ى	����h�yU��V���Enlv8�P�b�(ݞ�����Iee��2a�t��Y��MP5G�5,v#@Ô�غʹةca� -f$�e��ST����s�X��
��]je(�&�k�C�e��e� .�X���"�c�uŤ�̕�usRT���]���pb�4ѥ"ؚ�ǵ"LS]ZfPu�(SF������1��ڛ�X��+���R�k���Qq�VX0L��D�-���L�v!w�!@5�,��ɸ�6�w;[[��#G�Z�(3CV8cHbW������[p#q�DD	nҸ��4�$@%"] ��0[����hˁ*�Ա��Mt!�%�.�E�1m{bٜ�c]+��l*�F��t��& \2͢�*�M�JMU�X�θ�\�5h{Mee��%fn!�,Ck�U�m��2�����.f%B.2�y�����E5t1��1����39���Sl��8!��Ge�p��6lV�+M�Z`���X��]�.J�f6M+Wj9i8��դ�é\��ֈ��2�F
�e�zŤr�S:�ƒ���. �Wm���6��$3.�e"����*
kn����va�7lb��,Ң��ó�!�t��5�E&�=u4#�����B���J�k�n�#XҎe��ڳ� Ѯ27L��2�c��^t�$41]�em�ԁ;R$y�m���k-��^��͍�J�W��]���n9�U�)芐�1���E�v�u��2��P&�]�tk-��p�B�S����q���GU2
͵�#���[���Y	��2as���������/���E���R�!2!��Z�'�%� �ζo>���hT�Y�Di�7��E8	I���y���e�kh�r��[V��3r�v��̹����B[X��y�(����w�y�3�Nsy�dC����*����^g�XJ�-s��FlzpIo��ֲe-Z����vǠ5�L���j;��5���A\���o"�����݉<�f�̬�f�A�;l�=M��;�,���o9�g����I��`�y�6��o�r�C�����Y;}�7]i����2�4_��)"��|ǍU��e�`MzI�u����T�̮%�5�]���cf�[D��2Q�������l�����^�;y�L㶴�2�lOq�]G���ۄ��16�S�=k�u��k�u���k9���=�/1�{�f�0&"b�<NS�d�����hOy�{��ٻ�w�=�y��gy賮�o$�������9�v2��-��-��\���}�V��Q��+�ζn"��8 ������󶧮&��Q���28-aͮ�d�kKZ��5�oģX�gU�WB���j���e�pJ�A�p�$�$�p�d�<Ds�Zf`^���?�[y�L�gWfXM���t�!��'q���l�T6�|Νz�9
����I��
N�%4YL�Otӣ�����k5qآܹ:ٸ�㩟���q^d���)55��]��⃜ y�|M��Xƭ����U-[�s�[��Cf���My�]1�~�a�^����_�g�=�&�]����Ɏ휻�K/|ɅC�(}\9���z��T���L���%�aͭa��ɷ�zw��r�A��g���̰�5�-��C7�o��\?�L/q���c���堩�.9��������R����H����YM-�,���&���5o���4�;u��&G�1X�"1Y�Y�HE����aT)��|��d�қ���1���oE�j�/;�cԕ�c,A笹mkgZíc��z�{��W���>0�Fc7l��&W�1{ӗsB�e�w��0r7n��L6�z`�tG]g,�ysÍkE�q�5ju�czҽʛ��g�v�ZH��m�-Л��1<wo綳�'㵓?�B��u��꽪0�8��r�B�ͲY�P��fS���.Y��y5h(�pA�poJdC�U��E�r�/:ٸu��[:խPª�"Hs��>)4��UL����8���#�+ ?���휝�̹Bme��pQG��!,�v��^�����2޹�X��c1�Q���d'Z����[?ct�\H��Ovga7-�	�`��QE� ��BR��5��7������Ïȍ�W\u�V�b�m���;l��"����Cu<�7p��5�5�_}3А߱鷄T�Ŵ��92�Z!��P�f���^��DM�b�A��Q�r�������v����8"�I��
N�����3J����w��r'zs2"�Y}�L�<�e�7�I���ȅ���!����w��=���$��r�V����2�Pj��5a��Q���i4u-�.�=z�����|,�Ow�7����ZU�&�S���M�p`���j�cTn�0�^,=���$0�TK�"����v��V�ꆃ�F�����Z��,�\���l�A:��#���&����EƇ�@h�j[э� �BN����8Xm��J_�w�N�fc����L;ƭ����8!'�����Rg"f���'n��n�!c����Rgg5��7�\+�7f�A�`���8j�v`���,p��
o$�|AIÂ�Ut3���r�����������\0<,�-��u7�g?���
M�.5�#?D��u��6�Me��;�=p�o��=��!=��Y`����Ե��P���Ύ��;e�3��r�2���f��x�3`�@��G2F�F*[b����Dң�k̺�R6�X�ФA`4���+��ݑ��(r±4��S,it&��WLm����K-�]���,Is�
B�!�X@ζ�5�mdk&)��E��!K��fe�13x��骚�+ɀ�1I��,�+�!o��qS#nJ۸�������4 7M��Kq�A�F֑�Tc1u\eH�����}���iOz!z���X�e�,�Yu3,s3�&3�uJ\����'o�Yǲ"�X2���6��9q�gZɓ3���c��2M+��Wy�6�g,�91e�������E뿒o8�5�@ �v�C3����c����pA;�㧹���!'\:⟄3�È=n���5(�>y�'.��(���Zɒ5�9ֲ����\�Tt�)���͕X0<,�f��L����9I����E?� �?n��zWwݩ�x��x�r
Nf�ڷ�ޜ9�F��y����'K���6�4�Q�z�߇����,cq�8��AkY����&p��Vŭe5Eg�D_[+<�!']�⣄>�a��s�pQE�
��H����rŜ���8��`���6���;��pmU8pE�2:��֐�O�y|������� �x��BN���{\�l6�7Up�𳭛ݷ]�m3_�#���S8 �� �$��9 v��$�KS�T'�wA�p"9��2�tO����e�/G0��̓�>u��ۙ�Ӊ����R� ��y�_
f���� ��y����1���;\8�6��7�ffQ�k�����A�p�!%zⳓ(�!�GS�w.�0��\�׬d�}�$]��7}��@)5�u4>��ZHu���L.�:�����c��Ô�8 ��9	;�����|�/I���p�#u��$�q�U��nz�Vu�q�S9���쭋�eY����s��I�%&�Bw��ז��'����&ލ�y����i�8 �>�p�$���z��V;N�￞���>v��.ޛ\�j�Lcc��lj�tnW	u]���j�cmk9}z�����p.��o?�M�)3��gXNJe���!�����ZÛYV�0�A��p�:�9��!&i0����Kh/۸�p���S��+�e��`yY��� ������$̟�a͌C9���)8pR`� ��G�G�:Ê�ݯFq�D���i�-15UY��hKp���������Hlv�Z�"���k���ꧼ����B]��g_���Oy>������6G��2{����iZ�4w�Z��"�����y�O�<�m ��/}/o�k9��GSz=�Y� ,�dg!zbq�~淘p,��o8;���9z��l���^�e���g$Z�.��1�d�1��bס��ᔮ��l�=r8Vu�q�g �?�����QfTm�97�2�WK"���D�����ܙܱ2�յƫ�,v���3�U�e����dֲd��"D�?�vl�}�켱j�w�883EB��~*�i�L#�,`�U���&pA&�{�k,fp�E����3�`�?��u�l�J4��t�U��ӡ��X�ƈw+Mh�~2�8�5��E�u]]��dlC�G�p�"�����:Nx���"#tp`K6Rwδ�t6=b8Vm�=W[�b<Ǩ�kX��c���`���V�^y�-��	 ��.BL7���{.�ڪ����Q���'4Ap�r���YSQn9^@5��^��y�_�J�����.�o�I���=�62b��V3������8��Ҳ�=dx�X2k~��X|w�N��Iֱ�#X�fI�S5w7y5��U�l�]r:��,|���E��(����D�ޠH�[o�{ ͐�311�Z5��EفUk��]��*�r�%���'��GK�n�$���"�ۼ�A��J|+6ٸ��\ɺ�LK�ѭ�> �a[?� ��E8o$�ț�kRݘ!��O����
���Onsy�^[ҵ�w���_0r�b�2�(P�H��շ��ǈ &D9�$�>0�E�U�x�|�"y�eKl�}��3>�,G���b{��6�Y"5���)��#[)uj�$6Ėjl�f�V�v��|������l6�&Vu�p �:�E�2t�;���x��x��\��	I��'
L'v�A{��Q��Q�9��췞�e�+�!߃�ⵃ��!'��3f�ء��ޓ�YTf���5Jy�B�4�#�9·S�[V�jR����-���w��N�}�ǆ�&z:��֥��K��"f��a��0q/���q��=�¸�Ќ�5��RJ���;:]�Ci�,l-�`-�4`�2���A�-U��a��v-���H�Ecn�5���`�a5�-�S�6��@咙���B�ٺ:�,J�6ݳr�`�҅�Q�Ҷ�^z�3p��M�׉v��	#7a�tJ��X�o6�6��E���u�t��1GV�B]o0$�v&��l�LX��mOϟ>Y�ueî��M.���)M���aK�אŲ�Q��V�-���!y�4���7l�i3��s�ƶK6ݿ#�����->�B���#�Ô�8 �Jw�]��U�r7#��n�tX")��f��W_!�ܥN	��l�����&]�������GS9 �Ƀ�R$�|BL9��6'�;B�'���Ee��]�����Z��A��I��}�|1뽀Cw�t�h·���~BC�c5��Z����#��>�`��^���l��z����`����J|6=v�������gg9����k�$���nJ���L����3���&z�x0)غ�ϱ=�������OvhuE��b���샤P1+�V����f1��B�#����}��>^��F�=c��)0pAIƶr�.�����h�~��4��7�����&�l5;��D82M�)7��Ixs{6xT;�Q-,�������M7�/cX2^���W�l���g��.(��4��n�R՞��t�����u��o�Hx���&s]�����r1\ � ���A�{�f�N�������ȩoa� ��y'I���L���:��t��ݽE��%+�gS7	�g �qI��
L�!�#��Z�^C ��
(� ��;vjWN۽��-_Ky�7�:\���/�}1ɝKՇ�����)3�|Rg!Fz]���z5�q���r��Jj����h���0�An`M�����3�$9��w�uLGg�ќ�!�0�6̱l͢�H�)Z$v�ҡ��S�e �O~O<�4���`��<oA
]��!Ū����g�%�f���ݡS�����{R�Aȇ9l��3�0%���	\��=G��@84l�U�9յu��S��w{1��?��E�!)�[��b�Xl�@�����w������6��O�.�t��������z=^�p���TF��C�˸��z��hL{��s}5��.��8�l _U��O���Y���I4	9�}����7��)�t�8���,���C��{v�#[M���]����q�j����<|����By�]�.�
�p��Gc�Ǐ��s���܃��!y����H���pc�u�@o[��W�`;�=�{,��Z�X���`�Ȝ����l���^ʹ��网���.k����׎{vȼ�u��ҽt:��'�<,,���<rQ���S��$�
�߽�N~{:_sXO��G.�A���$���0��w��k��*{�/>�1L���c`Ft�	��z�y��<ż���d0��c����`�_.J:n�NRN�w�R�:^S��5u�Bg��g�c�p�͑y�!��ȴ�&D=HWw����U~����y��<���=�*�J�_M��k�����OFuT�j;�,�rA�pGש�3u�'OK2�sf�n���Q;��g{�3�h��ya��{���>I�ϰ �;�]&i�fku��$����1�v��ј�Aج��S^�nj?Wv�ӽ����9J�%������\�NB��q'x��C�Wqĵ-�ٳ��ވ�w�xvOX����܍L>���� ��w�1N�q�~R��盛��'�A���+w�ű�X���gl�|��K7V$�ފ5�sXR{}MG=��wjd�2=��CQ A��Ӌ�u)�8	g��s��&�iiW�Ov��v������˶w��4{p!��QǷ���ڰ��o? �x�o�MO�)4�S����$IPf�$��G�����O�?v�gO�����:z�88�5+��ª�U���i�$�(��$�MJ.�L*��T�uj�!(�r+@�!(�;���TQ��\�դ�h�؁ʢ�J��i�uB����tYEҧ!�VMք���U3�DU�:�aka.r.��(�w0ҭ�Ȋ����*�G(���u2�����I99!n�BQEB�\�Cn�R�x�\�(�D����:�Y�!�"��w
�U^��d�r���ZZ�F[R4�j����wD�2")�*'Z:� �sU̢K���U�W<¨�*�0Q�#��eW��'���r�"#��¢�Qu:"�5�Q3��Te�0�
.P�-4�.�� ��V+EL��EҪ��s%5B(VFEr(��#Q���}�_��d�(���xZ ����`����/�
N�$�%D�&Ϝ*p.��?�dC�V-�Ӯ+�%�f����A��g�3��E��>�n݌�"��)0Rp�jH�cf �`��_gm�?oDb�k��"��O��Âw�	�<�����������R���r�6��Dŷ��kêL�r��L�z�)�`G/�߶��!��{}߄9&r	I��9Z�o��F��J���3u'��V�6����0�>�p���IÐ���E�D�5�,k�4:���8C�Z���b�X&+:��m3��C��wN1|���v����� ��� ��9E����!:ݍ����S���W�v�H��8>8t��A�󀔿�y:"
L��L�	p�^�Ap���g�3��k�s��o��\ �0�3-`��.-�yԆ�i�ݴ
1c�aX훳�ߧ�����������Et E�➨8�c�aa���D��������󑎡�G�>p���0����g�.��*����z=-$8׻���o�%�b����'i�u��&���C�n��Sv'�O�߳��=��a"�����P�kt1�l��G5�s(��"G9a4R9���w����}��_H���w�F|AI���u�S�GE��V�H��	�c$�lE�������$��)3��0�S�����8�3�N&qs����wd�6%�Ab8��`ࢍ�t�5ko�#%�|�ceː@I���?�DvB��v3��,�rm�%b"������kqRg ��yD���ot�����Ec�
2'!��������+��!��8t�"6�2��&b� ���)��M> ���A	�Rk����@f�*,X.�꺮�C�l��Q+���0pA�QpAI�ݯy��H�ol���,��'�*&r���W��y��V�C�p��KTwMR0���p@��j]����]��%�b�>�{l�����Wѵ��P�mt
3YR�Q���cI��H�M�q��R���4H�b;4��6�	h ����&f�p��[��:��.�  ��j��E�<R�6�^B�yj�4)�U䦚ce4��uc�n%z�^*XR�Y���i�Kf�02�\��Kq����J:
�j���l�nYw6�����`B;��񶦰���}��P'��n��D��8�%,VXmGvh�La�]@�B�*ud���{����>���wBN�&D>*����m�Ջ����8�����JZ�sY�&�)3��T0%&�lHn|ld,��� ����t���֯]t��	ӥ�_8r�u�e߈c�$�3�N[8!��[�R`nP$�ۊQz���#�-�eS���]y�,N��%�VX������&�y�*;��6q��p3�?�dC�K{4���ہ��8 �s0��<,+�+ǎ��+�����í`�kY2�]�R��CpKK��Զ�y�^[�t���8'N�_8	K��Ds�ټm�=Nfm���E�遥�Vѫ6�Ʒ�D�k�Rҍ�]�c ���� ��Y�p́췸��M�I�\���m�*�W-�`��wz��*�`"�(�pA	8�ydL�ӏ��f䕗~�if���4�����츴<
� cf���1d���y<���~��n���T������%�Ģx��'j�������x�q��K�4�k���э���Ѳl�<�)������l�J�B�v�|�h�vT��fkUfD-W�q=-<=��็�a䓄�ܲV����4�����
m�:n���ё���2�%?7
���جM�ح�3m���o��]ۋ��S2�{�PUQ����um���}Yb�2��u���I�S��k�W#U�v&1d�xùw�aؖ �ٮ]+�m�#�9G�J�
��`��!6o��g�?z"�$�v�\��:!r����i����^w��F���I=����i��0!@�𫨞��bn����uhx���eTR~n����T��v����IoVc��$�$��P��6к!�qn�y���Vm璩����x+��Nu�W��l������"T���A�S������&"����3,��n2��m0�w?�og��O��:^�Ig�F8�iT��0��L����Z��娞�~�θxP[��'42�jof넘�y$�\�#�K���QV��cS摕QI��Ս�Ԕ���;�_�g��p{ ʀÏƓ"[/��2�\7�^س
L3��fCA, ����� f~�z}"x՛�l�=�^S6�;kѭ��Vy��'�7��Q���4�_TE&Ȏ�u����m��W�Et���u��Jy�zv��2Y�b���d��&��m�}yv��o/�T��xFT�'��X�N�I�L��hk��%�Ɏ���k�$��{4��T�Y-yL�5w�9��@��uⱽG��E�k�--=���>"tV���3��3��р��2�����8n���X�L�dݚ��rɜ)��~m�a�l�Po$���m�a��` Af�M\�5[���OL��q��G�K�����|��gp���%6�_�:u��e�XfR�J��nK�l�\������}�|��OϿY���(o��N��Gs��x���z�[��y��p�$�$�y�N�M�j0"v�ni	S|l5�3ux�f��&{�Gc=�{�C���$�-�.]�kt0�l�X�*Vs媞���N����M䓤Å_ssd.b���~�ד:�1�g��I��XÏv�Q�bU�ؠ+Iw��ރ��{f�\s���ͫ�"��7��^S6��m����(y��`�M;@�7B�/�͓�SH�.A
�@�0���O(�ɾ�Uic�i��|��������x{� l����>⚓���M�F@s�2�`LKH6��np�X(-�[4
1teffJk2�0���c���H��k����"F�i�$SUա.t7��1��`�tc`5΃��F��n�.+6a#�CV�\Z��퓋-i(L�Y������[j7J̳��B�䡦�
�u�r��I�M4t ]n�N�3�t��QWq�-�v� �Т3��5J=��O�����a&բu.�M�,HuT�\�)�i���Z���j�-t����y��`�q�>>�L;����V��c�L\QcT�<6Za���z�lx$�o��p.ܩ�Ê�)"�lJg�3ɮ^h�������V7�RT�8,a�i���aY��I���<wT���CiX��j�XJ�9`�S6�j`3��`�Jwp�J����z!�-��S���_UL�����em�N�@7���M� ����(��nS��Z��ki�7���[sw��	'	,u���Sk&��ic��Dv�1��v�:�)5�]��V��Q�X���iU�@�~������=�����hҰ�b��̢�f�se4����O{Ҕ��I�'�I�{"t�O�z$��QBr%�^5ȣt7SY2�2��	G]ټ_w�j�4�Wv��p٭�gu��M5�^��#�
L#UcQc�a���yrfE��pky��ja�]�d�ꨞ�V�\�64��Qz]���s	I��xR۬�:�Rkv��SL��;��*ۛ�/�$�����t�h�ˈ	����>����O�ŗ�M�7f��̢����ko=`��uο<����$�I��$��`Q7�������;V��W�Q=ծ0I�[�s˄Uc<��*��XK4F�Ƙ61��cD6�ոfQ�0��5�.bC�]l3Yeh �H�`=�޴��5��.f���v��nn{v�={qn�X�t��2I���m�t���M�[o����m�����s$����;�%��a̸%�I�I�>J|��}E�-�Wz�A
���x��Pp�E
2	�x���YV"��y���%;��g�á�ʹ�lٻ���q������Êw�,�z��=��<��l9�e�+����������*N�����b�V^���Pl�ٮA�f���w��nn�k�v΍eS�B7_�lo$��@��:�!���]����]w���������[|6�����L�����Q4H<�33�x!���-P`-�˫-n%^�l��6��Xs5�F�_'��or~}Y>{�$�'�մ�{���W�Q=��8#�t�Mu��o$����p��fL��&�erA�b���w��nn�^�~��He��Gs�f�����Q��d)������X��ۭmm�Y�3 ��m����o$�$��[�=k�NP�Wk�'���w,�1_J���ծ���Π�X�坠�48U�p"�9�,����!�N挨�}wLfӚ�#8�@񼰋6e�F�(y��y�w��V,V2�F���X�=���I�j�	�Cl��P�R�y-V�g;[շ7	��`�p��l�:���%��1o�n�)5b��SU����ir�Z�&�#Zl�%�ݺD�@�h��o0I�I�N���md�՘#2hxSm���,+�z���C���m�ݽf��Qo�:�`�k����{���̻����N��$����A�>�{��o�S��r���8TB|�-V��mV����I?�@({��6e��D��o���_>�k.v��9�[v�k���L�hQ���ެ�]�]��w��<��0���&r.��r�Ym8����:��Z��ֶ#�N�Ӗv������������=�gܛj��	����e�[��ۭ��t�)=��s��{_���0Y�ˋy�jmM��o�v4�����;�v�훞MlI��ǖ{��{t��X{/M.< 0��b'�h��3��:�J��ި�߇���u��OS<O����<���=Ӿ�e#�#��1�����W9!{S^I��R	=ĝӄ��� [�m�%5��͹5�U����{:�BJ��.سe����U��w�|����v���8{>�0�Hozm���'�;�V./��B�G��=ðF��-ڲ�fnSb>�:������E+��h����X�2'��M�80_/?:��͞��RH�_X1;~���G��=h��y�	�E�%����ʲ�����K�z矱���Xۋݽ���GK������4fvs)��w���y�f�z{'��E)���C���sٻ�ᷰ+���	��L��o6:Z緻�����M]@z����![�WU���9˽��wˆ��}����0}A�����<�H�3����{��bݯ*�#��s���;��	�>��3�����X;C`�{.��s��#�����_m�s-zr6��D2�ʏ4�}���m�+�9��x��p�7��N�,�c����={�&��=����S��5��H3����\њ����y�R�=q{f��]V�`cC��z�87p�bbWO)� {_�s���vW��}5���ɑ��nz�{V�[&��w��`//k�Z�kn{��d�L>1��A�.��o�FϿZ>�q/2)����8ed�Ȥ�Q(��fPArβ���9�$��ʮQt�.]>q	��5�Ȣ�"��+��eY���j�H̥B���a\���&�Q�	�����G��L���q@�Ut�;�\�Њ��K
�*���(��F��(�B��q�V�E�+�������d H�WuVT9�"���W9ˑ䊔됊9�U:!s3�V��9]�ʮ�PR���w/<�.Ws#�*�9�AU��Ur�Z����]�B":�sС(�C͖N^��R)�)0rĢi�E:��xeTy�*�it��\#�:�/0�Ny�B";�QA$f"r�Ur�w/
�B����Q^��dEʡ'&^����K�P�^�L�9Qe�Y�:Fr��@	�Ԗ�	�;~��~z?t\�Y�l�n�+jݣ�ece�,GO�u2MI|���1��6�
$K])Sl+ͬ�-`���Hmh�4n�F��2!0J6�4.
k	���֗8d,Av�0J2��oZ�� �c&�cjHһGp��6A��Yaf�!k%.17h��+i2k�j���MJ���͜��p�q�Ȗ�U n^-�W�b�[�s���Qm!]�t�eXK��.e)4d%Ō�����gj���F\���ΘAѪj�C5��v��6��Yܱ��ƳJ�\b�)��q�JV�,�`��c�ĵ�mâ�T
Ԛ ���nV].vY��E-X[�f��0��4�veR�UG�h�����i
�bY�٘���\���PtF�k���� �mr��:�-f�C,m�J@�[Qƴ�0%�mT��μg���`֑�6�@�MeRT��X L6��h��F,27�`��klqL�y53v[rl�׫i`�Z��3B�K76�&�d�Qm�+�t��lE0�4�,��]6amX��l�P�Ζ�32���#5�� �F��Q-cl�:�0� [ZͲ�YK6���R,�ʷp�[GRR] �\gCTX'�KR��+̍���+]�9Ś2�A��t�MB+�x�@\���R�)*�-��RnCY��`ˇ
�a�i�Z��5� T�8������uiIXJ��\�u��:�s.��f�d��qY�қX6+\7f���E3{ŉas�\ebaa�[n\]�yŘ���;&vBP��v%�C�K.�����Y�]-`K��T���mj�ֵ�2;:���k���3�F>Vg\��7'%��6�5��A��95���3E%	�L��@c�+Vf�0::�����	�Û�WR��%��&�V�[����!R�s�[7f��C: P��2�Q�Xk�Xq]�6��J ��-���s�3K�ba�Q���m�.L��]�jj���
�ζ-���6��#kl��Vi���X�	-���;�%��u�g<摖5�K��]6\�̃�ɭ:2õġŘj��&���hq�P��!�4�����)�����d��fL����5eIJ9���\��&6�SmX�]��E�f���b@oSK2[�t�rb���$��k˜��ճkbWAsVfݣE5��BL�GM��h����!VZa���m�B��V�lEԻ�MfR��:|����S��-q�\͕](\%eȖX2�!���a�!��`�E?�*oW۞��]���NU����c�nn�-g���ˣ��U�gk�$���c:=�`E�{J{�����멧0Nd�{-����]��ޞ�����M^���$�$��]��y��2ďcNj�Ym5�n��_7�o����ƭ���r-i4�8��m�l�5f�í~�ۛ��x1���;^G�3 I?��FG	sb�x��l����0edܶܔ��]ƨ�[�:|�6�� �g.ׂ�6,,��n�n\
k��7M��K�[������g�\��R¹��$��yVv�w�Se��u�������ck*�	&�S��!�T�]�?�ѯ	ㄱ�ݽ��y��-ų���f�}���/�G���r�ߕ�Ƒ���z���֒3��㸡�2NK;�j�j�R�e����ov@��j
�M�쨌�m��m�c ��*��u�[��l.[׺�&	$�XnIU���үa�����_F��HI�I��Pl��)�J�`3m�nכ��Ӽ���泭߽�|�r�/w���6r$�x$�ֶ�\�ݻj���>NsH�t�[q�d�nnSĔ�#�/y����e!�� �-��|v�LN�Fi�F��1��* )�+�����h�o����
�{�(I8��g��q��Y�D�&tZ��
��M��⒥#Ԯ��L�7i��{�f�u�o,�{y��w�t�_$Do?Ej��������`N�%C�m��֡���qH�ayH�MB����jc������f�>]
x��H�xm^���_{��{ˎ�P��w�(ؗ��p�$MH�9uo��2nۛ��>�I��P;��­7���V{e�� ���|ֵ�q�X2�K��z�E�e�'�w@�o$���$�W[u�T�&I�bw��6���j�ˬky��w��z��k���想٭[����K,��hb xp��c���שGv��65aW�	���C@`Z� ��KH�OXm��p�x$�#��
��u�����ޏ�?L#53{"y��:]�v����`����d{'U�e���9Y%�n5�:Z�O?@ڜ�7\�}=�7��y %�N�w��{��{��^e�5�Vu����V@�v�I8I�����I�>뀵����]VUe՞n���<Ȍi��i��&�)��oz�b����l��z�Ǹ��{����ӡv�x�� �ylN^�����/A�l�/y�v�F=-]�Loy$�$�%����0�g3 -N//w
�uՙg+$���Y��%>J���CkF�>���{�f� ��Li��YF(A���m-t,L�#n�M0@�)6O��{������2E��7b9��.1��g[�Xs0w�98I��I;���G��yCG3GR���:�6��,�H͐���uY�˫<�#�Ja����Fn�D���o��Y�	���G�y$�z#	1�8���sVe����7.�{��}v�{I7^�6��@�|ɯ�9�n����OU�n��i�=����*2Ekos����]��������cT!��ii��B���]Y��Vy��Sv2Iҁ�ѹ�E�=�Z����Wi��ҿ��O0g�q,_����t��F�tiy:dqaV5�D�C-�~[G<`��Uo��1�& Iō�Sp6�Ev�mؓ-Ŵm2��A��M5a�ݐ*֣ۭ�chat��]f��1��ܠ�7���R<��V��0ҭtr$��Sd�[���rq3�`��Qc� #��l$R�A���f�J���u�*��R�b��͍�8�wgd�jY�rĳ�͉Y��:!A��)TX��)k���q@�a���������G������݅HۮJE2�uf�U��mI�K3�kms!pF`�;��&U�f[��1���I�N;m_�����V"���'١�h��˯P	��'I�^��S��`�������M��7ݗ�곭߀���`��r��u�Sm���~L���t����5��C�[���l���U�vy�Jov2I��&�E�y�p�3�í�I��nwf��e����2�y��1���gk ��IJI(�K��M��ۥ>7�Y쪳��߇�1�rPOr�t�vɅm�]�'�}��qG`�2)L�4�)p��$҄c�B�W���\��$To���w8I�I�GD�5?r۳U�h�q����tt׳��ڒI�I8a��5�����n&�#�."�*Mȇ�[e)q��U��y��Ձ����Dr��2Q���g�"������T� ��ۼV5-P�'b1M�h�޵�(�J��(�]��7���	S�ۊ��n`m&>����y&	'	�,�rA�<��:q��*η~8�9y�)��p��9��4�2֟˥�'��0�Zi���j��G����>g;��4N�5\Lw`�s^E�I?�I�|]8��:���]�\���U�}�/�)H�w�(\�_���?-���&��x�,h&�&��-![v��v�kԢ��؇��C���'±�I8�[N,͛8��v[�>%�B	Ua�C���'I�����˱�9؟1�ۍ#���tu%�5�ty��S{���g�`.������I@����ʼ�3\�U����+{sR��S4w�U�6�Z'��LG�����?Ҷ��g.xw�<c�eu���r��+����eɭN��U�}�}����2��q���FMXMYo�MՎ�Μ|vK�[7����̝s(N��n<�yC �t�3"X���#1��J��Ԗ�V]���M��$�	4ٳ�4��Epp%�H�=T��A�)��&��lۄ4�.����i��������'�.���k�����_[.A�fb��}/��d���O��!����^S���l�X�k���d�.�p8�9���H5Kzc��J�@�y��$^2I�`��w�S#9mE\�%S�s^n~���IO�IG�v��gR&�����,e��z�����k�+���_F��\2��ܽ���-k_��O���w�7(7S�=����=ޮ��I��ۼ>�fn�S>��~/��J	y�����F>EԲ��^͜���Z�۝ut3��wp.��	.���2��@�fSl+8w6t�2]�e��:�9�oy$��ȡ�K�o<��S���{.���̤2��w$#�h���)4KfZ�+�< � #�W;N{����絞�٭ꤞ#r��5ƅœ#6�U;��$�$��Ϫ�n��h5��wsB�}�R��VY}���t�M��YL�15c=��ِ)7�o$�����]l�rslV���Fחe�g�3������hcJ�`k 6#.e�X�&�:�MoT��ny�J`���^�<��jݗ����%.L��6�h�A>ץ���}}�s�O)V�VY}>>�o_k���p��������އa�I�Ʋ
{�$Ȳȅ!��>�f�[ؚk��S�C7ۯ]�������{�fj���bK�fˢj�	>��������ծi�����]4n�,V&�t�%�p�3Vm��U�&śM``��#�M1E�Du�7@�PՔ��K,��FӁGSMM-P@�X�]S�]��n<�B�,f�%�[Hu�K��Fմ���!��itl�j+Ι���JХ�snː�*�D�hMV1�����R ܭ��mc�-nu�l�#5�%#fL��c[��}���fH0"�h]*.�͐)���0m�,)0,�f�vx���D�p����awn�au|z�8�a]yh�����7U.Dv_���.���y&�in{x������<�Ԧ��iDF�۞i�xR`:��Y�q�NIg����3z��/t��La>T�L^��p���s��jo���U�Ye�ۍᝮ`�:Iƈ{ױ3���ɧq�ͽ��f8��=��0��H���)^o]�ku�Rm�'��o�$���"����6h���ٛQ�v盽)���R��vp��>[=������JX�!h�V�,j��^j�7�~���?�2LI�^���5HZ�] �e�ca� ���`�޻���۶�8���"�~��������s՜��p.�7���\�>�����ᇍ��Q,��0��7{lƳ ��m��_s�M��k���vd�kċw��\z�-wա�����Փ"�y$�$�qk�6"9��;�˔�f�Dn+s��Jn�	*�2Mo �uE����@�k�I8ݷ�k�M)�c/,�{��Z�e��w�?hY$�I(�I.��k�)�X%|��mّ�׉���������U��f\p$���5�!(������:�Ԡ�3\�-Wg�ֆ�l�x��Ӟ�o.�I�)8��6���Q���7��!�:)��;�Rog��z����{����$�m0�ʼ��Z��Β���_��7�ҥ�w�Pr��mu�k$Ƶ�k���n����������÷O����W���� ^��.(�ҷW?v]����g���9��� ��e����y��UW;wjٓxxd;�'�� 5^�<v�׋X���^�`���\|��&ѩw���u{��-�O��=��-pͣn�r�h���p���˼oQ8�Z8ŗ�5�o��vZ}�^o��W�f9��+H�=��}�B��'}=�fRFM	�\�àf��a���������E���v������^h��������Dw
y4��Y��f鉥��od�/>�L���b��F&�m�ێ_���C�7��M�:����ب�bx{�3rY���������b.���Xl��]zx���*�����=�_���I�c����d��=���+1'�f��|uO.yO<��*���6�Ƨj�]�>]���n������|�GIݔ�h�za]�K(�����KR��'!��Ք�T�7dDU�#�j�WoM�W��h�9)cF;�NC�����~�c��F? i~�C@�����t�q�~�_#��২�|�Q�:{���Sܞx��gn���G�pm��⫑�m �=��pĻQk���{�ڐp��՞��l�l9{��qЂ��-[Y'�]������\;��;���ݫ4�N����ܞ�k��S�3i�~6O��u郛-;�<�iX	�a=T��49w|=ݜ�)��E�v����p�v�𹪠�_M<Mp��� ]��R�_��9hH����Y��C�]��<b�@_3���ׯx6�x��S������.Tr����H��ա�#R*""9¹J�L�UG#�F�Nc�ʝ@�\�(��\(��L���AUUu*�r��BM��P�jZ4't�"��^J+�):ʼ��Fg.�T�E&�w�UȦ�E����Nd+���15C%D��NHjĨ��P�UQs�(�JTiD�I���%=q�e�G"�� ���V�G8�QȠ�ṪqY
����R�]
��4�
�TE�	Pd;���D���i�YY ����1eDU螡R���9��]� ����y��2�j�:�Q��^V��+��-֑Q^u�mdQ�I��!Tz�u+�'
)��ʽbsA�9U��I�U*;��s�n�&Dr#�#�r+�*�25"u"(�(�)srp��X�],���r��E9�r=0D���ՑD����`�z�퍹��ىᷮ��$�g��>6c�y&i
5�����&�ZRԺ&�7/�p��\��t�Y+��57�o$��+���-���w=nn`\��Ε���/�n6���a^>MpL����Q�ևｋ<�$��H5��0��E"���ka�ǵ�ԁv����<(��@�8��a�}��g~�7�0��v����!sf*/�]l�{w^��}4��oz��$�$Ӟ�UX'rL��ͬai�"����&�7/�w���l���__�7$�?O�3�
�p/��v���8������K=l���eB�9y%�e���)&��,�.g�u)O�L1��_���|\�����i�{���j���H��j�n�O�����P��d;�VV��;�qNz��i?��� ���}2�EK��d<L�3Cs�V�od�<�:o�p��t�\�4�E��)��l�\���n^9��&ۀ���%o��|�o��L��~�SΣ�`vH��\	A�9t�XL�fleV�1�,����Ͼ�����$�{o(��P��^I~�E�M�8�7����$�&�|�5-&q��λ�x�kn4���6u�.|�E�j��J�B��i�WK@]n:�±������]�j8qk�h&�f�n/����Ո���<��tXu�I��$õmƞ5,#��\U��?�7�0�I�]�x���
����e��U���z�p�G�p���hm}��=V�3�M�k���/�2��j׾d�$��qr[�أ��v�zzK�MFD�4�<:��'�B�1�1�R�\L;���͊b�{A�b^^�e6a�a���շ�ړz+߉��E�)`��ڍШGKT���Vˮ�Y�R4*	��P˱�&Ѭ75����:��V��Me�X��Z-��5�iX�-��n����f]�Uж�ۭ��b+�ֳK]DW0lM`�`i���i!����t���"VfW�
q��3]��Hخ����e�MD���R�l�X�m�4��PF\G4y���c4�Y�4�؛*![�}���t�c[Al��I�2�c�F;29�j�n̒�6�`Z�%����M�c�&��*��n��X�ܼs�ޕԨTd'�4���l����n��v:�r��]���[˹�{o��0���/$��-�����퓌͍{q^zg���L�t���\�$�=6��U��de3����/�&�I%"���
n�U}�)��BM�\�7I��ܼs���NU���W3��s�"�$��i�������UWz�I��v�y%�,`7��d���c����V��dxS',`�l�]�F�J�Y���2�l�^R��Z�Pٙ����=_��IO�am��y�`�����w�쀵V����W-���'�]�� ��6ɫ�=4���iV'6h[����.��`���e�m�UGֆ��-^6��塊(����ef�'eE�K�G�d�,�������Uͳt���m��<�&�s$����\K��dk+q��#�'�]L}T�P�n�o`�*�1�$ʽ����k�
���\?tܶ�\O��OM칿a�n�y�`���k�vᵯ����<�3 �8�O����%f�����;,�¦5&ٺI��m��<�&�	�:I_g8f��xߓ׭ �-��:k���m�1�%�m��-�6z�C32�7)0hr1���Ѧf��W{.\f�U�Un�[�"E��=䙯p�az�)ʿ�p6Xy&I?�I�͸�����^wu�kcF2잀�%_G5�p���o%`�%K.��Zw\ 1�&	'	7��暆�[6��*�H)S��'h_X��>'�
���k�}�t�|{���(�y��/���I�%����M"tN<N�4e�1Ǉ�L0��1�A���n�{�[2��7M��d���7��ܳQzw�yM�%Y�x+q��]�c��=���y*j��ĭ�i�
��o$�$�$��n��ƶ�;
h��s��~�y.��q|�0Iou��_5�y��8�Sg�K�D�Ywd�e��+�c�Ĵf�ÐHfv��K����%>I��V�����`���<�#d��m��=�� �PN�ٗ�׈;;��Z�սמ��yw�����q���|���|9Nٖ�c�S�`��0�R���'h6	My���{k\_2M䓃䝐�F��l�~���M��f.RuĶ��<�=6������M<:po�x,:�X���:<�Ӌu�Ơ�=��W��ν��/�����\�	G����֗�?��7n{-�v�x�ġRp�%�r�[N3�n߯m�E��z�3��a��^��)@����~ϐ}х��D�#kACH�%��K��l)t�a�0�]��9q$g<�x
�	'I����'�6IF����@"\F�n.㉆�K=wwy�B�kn��V[xn��jul��N��x�+�2�%f�1<�b��du׫WcݰI�Z�����; �L�z�[$Z�OWtn7���`IO	+��5��ۺ��v�ҫc'�6QF��v��8D=,�x�m��{Ӹ�v��ݼ�&F�c�C{%fLܤ�mW�y�Joe�Iҁ����.n<�s�ꘅt"7�Q��{/��͹����&̵n9�������o��<�U����\��?��
�P�׊�4\��m ��P���E���u�]�X�(	�˭���ŷ��јq�Y�ٮ��c�D�m��lTf��ݦ����@Zڛ�:�+P�������MR�bVP�-fE��+��=b�Bl��ך�V�ͅ��b90�Rka3���� #R66���[�z��u 6j��鵨
m&��IAM+���v�H��i��uHM�Y��h����d�b�nJ�o�����k�A��݈�-�Ҳ�NL�m,���Zu�#C0`��� f��~߇�$�	'���0�tP���\�4Q|�l�Sټ�L�po��Z�fNH3��Mr�V7���b3�>"�bn�v�l�|�,��H����'�o�L�t��d����u��M'Vj�s��/fm���	(`Cƾu<��x���$����0�tPK1:�3�q��M��-������&�Y�&��49�s
[(��h�lO�ݳ��I+��﯆O.QN��" ����-YcN�mX�=Zū�YpG
 Rݦ�fB_=C����{��_�m�^����M*�گ�w�/�1�?D��4g�cWs�$�$����鬾����8޴m+��^v=�����;�,cͻt�30��%&�`Z5��L�Uꬱ0�֠c���C�iK5�f&��fjT�Ih���W���E��չ�q��!��W"F[ݲI$����W�u���QZ؟���g]�|�$ʓ���S�����v�	�[/�¼S7��wnn��umW�y�ұ����T;=�����J<�p� �+hR�R��M���ݓ�M�չ��Ὦ����|�z1�'�������e�*����c.���;an��[̼5��\j\�@.�"��][{���p�kF-�Μ0�sb~�v덜�j= _G�]���&J1�tGK�un�zn��ݷ�Y�*jUumW�y���l�l�1���H�G8�^�q���v�y�D{.��\C�ܼ���c�?"K����|��įj���`���0�6�z�r���(�c&`K� +���g�h�e�nk���k��Nc��������I�'�i���zm��1|� �hű����2��wn:�»��g�m����lݸK���Tt��3�ؚ�˚uYE�U�n���$��Oe�������9Q��8�6�h�e�󭌷U�,�b#01��e&����]���ϯ��}����F��*N-j�zے'��Ǜ��;e�6ݱ�1�#t�a]o��&	'�JV�}AJ;��!q�f;f�;�e����s����nIY)���W���z=��Rt�����#���r;&�VS3b�{n~�����k�$�)��L5M���5�|�'ŷf��$O%9�70��iW�
#?�L��+$��˥*{����"�q���{�+�r��U��=��&�O�B���?9����P#o�����vT�kp�`jJ@I�I-�fKz%�5V��:K����u�1�ۀ����0�L�wM���ֺ��p`
� ��� +c�1�fCD�e�[�\F����۱�@�FXaȿ\�t���%2+>�2��-���7(d5�9�@6���s}s�&I8���,'I��/���k.��ۙ<�aɸ/�n6��K{��9�O��x�f&I8	^p�UL�a�<R�y��T�Q�X���u̓$�/?�p��C��x�����յ�y&��V&��UG1m��<��5�LD�J|�^9wpݿ�d��&�����mw[��xۓ%=�Ű�7$�	~���������X�?D@W�
(��׷�/�� ?t�("c�r2t9��8��<Õ��aeedaaa`�a��a�f�Fa !� !� !�@!�P!�!�!�!��( 8���ea��X`�"+�0���
��VTXaQa�E�@VTX`a��DVXc�U�V X`Ea��Q��TXXaa�E�DX`Qa�E�DXax��TE�TXaa�E�TDXea�E�K�a�E�QVFFeI�a�s��9A����Q�T�A��Q�E��FFFRFFF�u��AΠ�����	��TUR*��1������׿������~?�����C�����ȿ���1�.����?� *���_���Ҩ ���� U��X��� ~�����|�֠ *���>?S�<9Hq����4������1���+c�� �@
P )	Q%	�	� %AXTY�E�ETYaQa!`!`!Q`�E���X�E�DY�E�YX	DYXHDXTXBD�E�$``Qd%f�E�ɀE��0X���?21E�A�
Zo��?����~A���� ����h��C��}~���à�B~��������N�� U�>h~��m��5 �
� W�C����" ���}G=� *���L��G!k!��~����{��� p ���C���  ��%�ۯ>��>g�8��|C�@���?`hp� *���� 
� =�N��)>���`�`4�Ӏ�'����`m;�$�ǐ@W�ꚓZ>���8�2���<�� D_������ �+��߽��/�>�>����e5���P;�� ?�s2}p!O��                                 @   �(=�(                    @            P  �QUR��*UR� �TBT�T�HEQ	EJH��EJQ"D�*UT�UH!�P(�R�   �!*Q�*��	A �[���{��(��(��R��PEg{/y� m{�
Wv:�� �U,�� n��  �  ����t��� : )��zD砠�
��B�((){���XG� �m��{(P�I
��(�`{�&��i�:u�-Pu@  �  O�PR���*�%@�QA)\ 3`��^a݀6:�޼@-�%G���q�۠Y�@�-�B��F{9HUw�@     ����G=��
�ꪩ�ɷ{�P�O@�5�`zQ��sА���ж'Gl6�z�zP24�ް�R�   | �*��JPT��($���O}�u!Uϰt<�(
���*Jw�Q���M�f9�����)GN{��HU�@� Ӗ�   ���E� }7���r���4��ɢ�nΊ:�ܥV������(   ��_S�RR)!%I$���JU��9��S;: d4v�(�����;!\� r�4+9B'p)� "    �} ��x � �(`��� �@#� f�' G&�@d �q��   �   	ꢨ���"�@� m��
�gBT���L��gJ�QUޞ�<� �{�J�0ݩ*�ΝiVԫ��L�֣�Ξ�h   |   &�'J�!�҇PN�5y�J�2*S{:����#�%
�;�9���{��
��3����н� ��Ɗ�Bb 44S���)J��  ��R�D����46J�$�F�di�M��RT�ʚh	� �Q)�R��z�&��>�_��Z���W��]�hI'����g2�'(ۏ�r��bm�H	&j���h	'���	 ���P$O�@!$B@�������?���?����z���媔i��ª�^[��6��yG�T2�c��Ue�.�!�ʕ33u�5O��]�UDQ[B;ʼ�`F]S(��r�/4l{�;B��cnPJ�R�X��oh�V���>�����cS6PT��'�T���(KE����e���ދ�f�Zb�U����aR8Z���#1H ҉5�E#n�LE�)ki����nA�$��ٷ�0�8�Z	�zt^Lm�iى[�)cS~P�Nցe*��6�h�9.�l̤jS��YLPٙ�����m�ż�f���rV]\��a`�T2KB��Ģ��ǚ�0�Ul�(�ly��c�yGj���uGhK���A�f�a��@��������N㢲�e�F�,ڬ�x-��j}0m���8�b ���ɰ�ۥF�	��j��Ӫ�F*ztV��V�e�0Ф��4�^�{�t�X2�Q�����ҝr�6�ӻ��[VI��y��ә��;��]�[�u7$��홦�K��P"��Q}��rU�Z�Qn:�.�;�jnv��m�S�a1MU�d���I�AQ�Ut�� ț��y�U2��h��D��R��6�Y�AeV
w,Z��Ӵ�扮����Э)(���N��P�ɗ���27Z�F8�T��h�퍳� {�J�r��I�ևY2�۔�b��ٮ�]b��f��N�JQ�^\E�76V�B��]�X��F�W2��'bD�/%�6�g��<7��3"�b�m4,-ψ�I
�ɐ'X�UN��Tki	�@��n��s]��f��v���6J'#��ZZ��bK$�z��;ݖ�vU��+��U�G6��%G>կ)zu�׊�M��B$�b��cl�`�̪̀ʚ�t�{z�����:zF6q,{���rq��J�����hb����k-j��wE�F��Y�1^�(n�X�����X2�V�.��ڳWwVlZ���Z�H�F�7u`L�i���M�Z!�ڛ%�D^։���U�y��r�(���]ay�5&n�XN�'��X��Cj�`�L52e�x��P�U�K8��^X,Ș,�gj�/]ѭt�������0^�)Qɬ�s,�h�̬f�H�.9����Z`�Q�X�ueY��H�Z۳{V.}/YY	.�d�p�X�ʅ�P��Å��e�^nJeX�U+�FVc ܴ]+{L��� ٰ%��f՘U:#YqdM,���Z�5�v��X���hau�mJ�Y"�n땕�9F�5�[��j�Pd���,��ӃhK��z)!�V���w��[.��bi�n
J����c�Z��������򅶤�YOA�Ӹ��P�)�&`h���lQ��\�Ph�S.��^�d1{�(�6B��֢����$s	�0��[PnY�U-w��Ѣ63!�&[���N�Ĕ��0c��Nc��%W⪽��[,0j����K*{�fI��f�Q���̈��uk
a�z�[i���K��0�ǚ��Go^\v�N'���$�l6�CN�s#�W6��vP��ŨoZ^����Zt�������v�,u�U5X��,�(iӛ��&V�#W���p�AfV;�D��I�V�ՓMV�U&)z�5#���v)0�C�f�kr��X����D�[B��͵��jH�p����A�J��PP�*L�̸̚ⱌRZ�S��t6�2�a6rR����+n1Q:%h'm�1^\8�����f��]m���VU�����+,�*�b�+owt���'b�f�D��� ו���W�dx�$#�M�#zlՍJ��1��[ˡA��A[�uu�]Z�^����U=-���(ά̴`��� /�ӹsnW�7u�"��q[L8cj���9Z��LԥM��J�Sb�Q�x��qJ��j����bU*nC[j^��-^��:�2_ʄ�a`�*	�YB���ba:�P�#uق�U:ԫ&���=�
;T��t�
�{C/nn,�5�M��`Y�BZ�w7wM1*&A8��ɅPCm�6��b�j����H-�ƴP�U�4̃�ݣ�ee�����͂YP봬KY���N�Yǘc�7��Wn��cN��)i6�V�?T���)`TlH�͠c�l#���՘*�Y,���C1�lvUR���w�wq�4�{��x�%���^Q8�t%^���-P���d��&8�9{�Rr�!խ��-Ŷ&mY�b �6�@Ś([�ɓ�9Ck	�m=�Xt�̨ƩMfï$_Ie-Wz.��v*�jI�	ٖ�u��'aX+���BwVۚ2���hc���,֊F��mC��Xȷ$��z��L3t�b�)�w�c�������Y�%eA]�ob�E8�ͪ��1R��]X�ٗ��H�lPʙ���^孭�PV�or;'é;Ui}��j��hԋ)��Y.m���5���Ԫ�:�"]�n�-���2�{u�[i�
X�3fhƝ�b���*�V��]�zaZ�c�3�f]����#��f<�Aӌc��Kf��cS�ۡy.�y�g,�������3Rt��uV������w���2�<Ud2�Gv�M��z�-�kx&*-�hT{�ͽ�h�ujHƌ�e�x���EGjW0Jª�����/Cݩ�ګ�ET,�������l��Q�DQ�T��+72�m;��S��9i
��U�B�ϯ^M�f䭼E)�1,�slaT�E���R�x-��Q�bͥ��/r�]=�2�.�mһ�#���o�Wr�Ut��{/,R��AzqZB��u�Ң/os7T�$!��VQz�nMƞ~Ǥ=��I�ỡ�$qr���'(���K���/d��x��(Yh��:���3NbSj�\P*[���Ճckl����-�(mVc�urCkj&�n��)�e'��9Bhr��h����K�w�/+t�ɘ�YD�۴����"Z���tX�0�e��^��Xs_hp��&dZr�R�,����Kyy�,R�.j��h�6]���(hA��ZXԗ�l�Y&�/R;5���,��2���O#��M-se���V��@杻�/fh9�e$meC�`����wH�ต�)�͹��`m���kh�Ͳ�e������Җ3>6�lټ��N$�]LrB��Y	��Ʈ�f*�`���AJ�ϔ�Uu"�hi ���tE-;�EͶ-�w�l����4RbH�m�h�Z��)^ຣT3�����T�^	Nf�&6��{��aosrSZBc'ل]�ܥN��cw��֡G���)`�7*�-�f��$G�����;�����vs-&^�j�͟c��k���W���yCp���x�������(kv�sn�ʫ8$�3��aH�"�SV�&�w`�%����Iq`x��؛ 8-y1n'5eAXm�on���	�Y�}5�oژd�u��w	U�T��vi-?,ݭ����.�mT��H�Q�*�Z�mW��an�8E����gR	f��yPV�^F֚ה0�n𕗔vд{wT�t�y�eQ�4:�J5E�f��V��E=�a���,94h&V&��K5Ѻ�����u4u]7��cG2梴�d�v+�[F���mP'lێ�@�!��FQ�uN�/Q�r�ws�.�Tj�����Yy�DKҝ�z��2�z�dڼWKV함a�r�qJ��vkS[���wN�WٹJ��wQ`1����\;��d�V�S!`N#���NڥF��Rn�ٔ��9d�T����Tݳ�˿�fl���vۣ��J��G
hk��e�MB��ElH���7w0�4��trn��3]��3c&b�S ��Zn���5V�r���h�ĕ�ٱ�Y��4��2෮1����]ŗ6�B���^�R���0���0ʛF��^���4�T����דU��[��Q�����b�3&��Z�$�՝��Q��l��[d�iL�&�*��v�Yt�Bj�H�Gf�kSEb��7UD��2��ܺʥ1l��M�q२���\;Om^+�׻ZXH\�F�j�Beq7m[�M��B���4����K(���e �=�4i�.�fV1H�����sdq�)�3���T��ZȂ��nK�9K�F-P��!�)*R+6SV~��\Sv���KN8�`+j���̌�5�UjV-%�$�Yx�]*K~$�fU3�-u�n*�-gߓ͙JI�4�Xqm�Y�A�ӏt\�{��h�ugX����a��8�ݥqQ4�5iH��j4�Ne[�:�z�I+�N�Kxn��8qQk��
.VS�an� �f������N	�Csv�Ȧ|j�L
��ۼ��XTb���0�u�:�5�w]�caմ��S�9��fA�ǓFY�ɸ�[;��b�{�Tz����u��t��C�uw�{6���ю�N�7.fUʺ͎��.�i��<W��������̚��5VĻo`o/,�.Qt^�[N�*3��5�g0Wص���"��%E�:r��Z��޺���#��~4ӣr��jl{��������+��I�l_ҫr�ƽ��a���6���Zl˚�p�4�Cr��fӲV�+c��n��v��h�1�TsmL˦��x��v�Z��᬴oU���u�*�a˪E�����+~�������hWt$7���YP�WT�Y�R�I��6[Ǹ30�J���I-�mK���m��(�V���=d2"Jk�Sf[���J�Ձfv�R��t���Tq��/D�I롌f�x���b�)m�Rڟ��cUT6�#8[O��	^nU}�bM�{$���kj�sc5��&4Y�ի�w�j�z��R�f�3J���]�ڲ�k��3͒'4kIw*�/k�����x)6���F�u�ቦ�[��X�б�ܺ���U�)�r�D�w}�r��G]V�+,��[y�NK?f�l��I8�Th��γ&�h�j�u�;X�j�G�҂�8�����i�h�^�#������A��X�9w/�nVS7J�l��[�ڻ�+�Wb�b@�Iյ�Y7y��i����X˰��iR�Zش�ǸЧ�U���/��X����rʪ�GQ�$̎��+R�mn72U��(��R�.�lL+���,9b�U���#V*��Ԃ3�k.��a��y'��j���a`�-� �+XҎPlmvՐL�x��r�榴j4r��@�i[n����9y^H^�J���0\�Z���s>CM�Q��5l��%vR�����&���XH��j�(�fЗ�o^4���c�����"]���ȶM;��6�v6+@֣Xi>6��o>��ZNi޴��
���YH�H�f�m⩖�L�n�7�R�b�ef��j*v*�	[Y3��ä�b����S�j�5.�G!�� �z3�.�Zi77h��y�H^�s.�eVR�d۵ko��������j��4��R�K+o�v�R��V�جͤ�j��"􂪆�����n;�b	�&����k���6�Ub�q�R�SL����`Ow&��̕B�R��uL\ʋj�f�G�I]�J�9+���U���t��;�F��ܽ�Zaf���TS�Qմ�Ta�!�F���]���.� ��캫yz3^�8���j��v���rӢ�����ݲ6�����']D��SN������4l�ӡ�"�:���4⫏r����H�J��ڼSF�I��C���UUVyK`E+v���Ԉgب��Ef*!�y�}����������B��j���[S/M��AKu� V�kU*�R��nXwN��xA��RE�X�ӂ�H�a���a����,�p�t�WA�T���ľ��ћ��mh�n��`̥uW�:�譬�Xq��ڽ���]�)5���;.\���h�5=Y�/l��W��1&��CM��+d]Z���׻Z
q��ɳmM�Y��K3B4�ktVCc+-:��Y��e�9pd�g�����j����z71,��"K76��wff�gB�u�������C.��;��"˫�\�ڼ�d�.��7�P��ŵ�ܓ+#��X�7MQ0p�̀k�+4��-mR��[�����=�̽-�m��V!G�v�ͅ�ե{�qi��1Mi�5�&�Bn���[f��j������+i��U���0�}@�a-��nm�P��+>9iÖ+p���T9d֪�E�'n���۴�ܺ-ݜ�\ ̱�h�i��T!�JX�[�c!�T��E�p��8��wj�Jv����P*̷�N�5ZC3,ޔl^���˖,�ű��tȯ!�{��i���Kz4ʹ�
ŵ����'̥�~_��)��`�%��*��mYxF)��R��5�Cr�F2���Pڌ�Z�V�դZU��vx�H����䫗���3u��$�d�9,�=C`u@��;���ѵ�E>wb$l�sq��M�ȍj.�%i�{$�]L*��re�e��̚��W��|ޕ��_ѽ�*<�f��Z�vD�'7k�uxˁU�.�hv�U��#ռ��4k�&�٨�QCn��͛2CY�Y�LV����Kw.㎪Xf�ʛ��x�5T��4�ו�ڨ�P��m�F��Ub;n�b�צ�T�st������-a��VMA6��f���u��[3,D�8�7F�ZLR�Mn͔~�!��bV6��CYn�kF�W%Q�s���5�1���+wv�����ck,�(������[���t6T����Pj�m�1l�F���X��i�5�#�̬B�:�ج��j�^Tr��Ղ���г'��çr��7!�[���[yAQa���^ڍQ����j�W�+6)YT��AʂItڱJKܿ�b��1T͑=�5nS�e�NKA�;Jf��f�6K��tt-��gf�;ҐR���[�6�iJ�HJ��pڂػp4��B^#�aJ8��G[S��ʕtv��ݸ��Y`�۷�[��	\�ʼ����	X�J�"ƫN���P�v"b�q{�5��S]�3�%���s+n�9�Y�0�7�Ꝍ�6��]Yc�*��K�T�ԗF�IT���+�b�K"5m�j�`�;Iފ
�����Ul��s�_�����`BE H��HE	�@! ,�H��$�X��A` �,�I!I 
BH�H�BE� �AaE! (�XIE �H(��$��BE	 P$���(BB)$��I"�	 ,!"�	�㺮���*諪+��"�$���,�"�$X���B,a �$R YB,�AH,���H(��H)X�H���EAd�A`H,��㫨�:�㪎�*$���PX,�$X( 
B(XRHE��
 )!����X@XI"�@��P�H@� E�y��	%W�WD�����YwV"(E{�,wt��H�ЪV����Z:P�f�.#ҵڶk��+��7~*����V�M��]һ���*��K,��n�BݖsuLN����ƪ]����7/xdu
j��l��6��ʅ�M�U�sZX��B���A<%��rp���=3Y��]��d�ډ9�5���\����׊f�³�3��UVj�ss���p�1ދ,$5��6��&f#�d�0����^�mZ̸���48yHPs�<70^�ᕸ.��������X��/VE:+�<�<*���{6�7n��ݮmmZ���j� �>�mmf�M��¬���f��r2gl[�h��c%٨��6�-?1��j;[Ւ�h`n��G;%�HT/l<5��Hh9b��ŝ�6�x�a�\q�wz3*�$Z���]W�u^T�l��M`�אᕊ��&5U�S[Mҭ��y�Rb�(Z�E��#��4Ƒ�H��9:��'z��+��t���-�h�_�$&�Q�Gc��M�	�Yei˄�8 ����X�tt��s�̖��+z-j��Օ��!Y�z)�t����T읽���(�`�u�����쇷�NVa�}R��]jnC��U�5MWs��İ��@��i�:�Nt���3��+c�a�yz]����֎��������,��D�v;G�fG��ox��e9[�/���oZ���M����S8��-��4��hΒp���dǐ]�U{�0Qow
�N\�&η����4�q̷}:�Y̲�vA}�N־��s��g-�+EI$�`�R,�<�O4��͆K5��6�٭�V~��x��6��y�*ƥ��;�
*Y:&̢���']���'u��.Fm��ݡy�N��@�T�vt��&U^
��4b��]�����O0�.����;(e�6^I��(j������(�Rl�3����:vu<r�]e��惒���s�)v����ua�-8�T���~�ۣX:c��х�qŷ�v�e7L����qn-Æ�,�so.4:_9����E⻶���ukt*��b��R���h)U�L_,��)[��:��r݇�ͩի+1VF�WZ�t�ճ�����'cܙ�3^|��ڰ�s�ԩ!�w�`!_<V��H�q�oVi�@�ڝ0��U>�$YF-�e�XX+l��
f+��N�V+3������o�U�{��y2���kU˾������F+)M�.�U�5�}��ڣN�@�}��������������[�j��>���4&���`�qg+k]
��#�t���^v!F�叞K
�*g_j՚��f�-䴍�ǴP�	��d�{a�oٛT�m�Z�7��.���/��8)��]��Wf�}���I�y�7[҉��b�Գ+���w�;~��v����R΄�oǂ��� ��UW��	�'Y��S����@�t?���jky�RżW��:��6���"�e��Sku��4v�cs-n�J���=��pZ�pd��m��X�Kn�XqWwb����VT ��ح��B�T��{k�^�Ӽ��i���]�@�{%��.P�kI�r��ܸ�m�������.�쳝k�-Ve^Mw]�kb����[��msC4��Ǌ۴��:כ+/`Y{��g���4�Z5f���;=1i4qj�w��ei��}HK��R�Y.���ЧP��b]���b�+:�^��F.�[6�7n*���s��K�a���7�l�39�G5ݺ���M,WMw���� t��LG^�J�b��zfgQ��^�ɧ�ۤ���k����K؎>4�h�B�;0�-�Ųj��ٙ1]T0ܕ�J�vڕ�M��T/8j�6������:β��h��%�`[ ڗ��Y{�R�7�Rû��
��ӷ`<������k(e�=7i�J��Ѣ��T�ռê�u�]�:V�hk�k%:�fu����s�Ugm����P��ż�M�qӨ�ŵ.�a݉�n�:�A���i]WM���'�2�r�!�]Ӳ��m'p��Kli�ʮ��q��TQ���*�G�8Ղ�oQ���f>�¿��}j�B]Y*���ze�ު�|�7X��*�=��U1T1d�	s�b<��Ao�oas^�em���m�]{Γ
٣URkloq�P��X`\6��E]f*���P���K���ܽov�onb̠`���5VL7�wki��tfa:��.&��C�o:�g�z�8�'�f��J�ʏ;�D;S4�+��j>h�%A�tr�̲�% +C�2Kf�h˲(�S:�;+V�m�2�d5���k�ѹK9�A��ϧ2����N朡Z���{���3.-K��jңͺ3D9ש���n�E��tN�}�V�f�kE�x'e<cK�p����j�t�6v�5�b���ݘ~��ӳ:��]X4�GRU��ṄFШȷ�V�b�qཱ�Uy���oU��+�&n��V�����qS5�WH�P4���Eu�vҡ̻�zl�r�qf��j�d�4�����;��s����f�fm����X����N����E��� ۟GY��WK���̀����rź|i��k��2�����9\G97���J��er�W�uq�p=�Fp�����(D���-[n�O}ISOg#Em\&_G�r������ob���/i�]�6��`��â���|C��O�<{{���Φk{���Z�
V*�Y9���9��T/E������ƴhr�xm�W(������͏:�Vuǯ]���\���[��4ڗ����� �]��J�����i�߶����Eq].��n�˅���^������eVo7�s���ХX���tyһ�+q��i���j�+���+>`�c�G^���+6Ӽ�dX$���
�^h۱YKD��}
3v�5��0Uݜs�e��Q������5)<5ؚlR���+򾼕 d�r䫭���$"�X��ׇ4SUݶ�/��M�<B�|��ZFn,��n`��� H�[Y�#t]�ÛYc+n�y�bE��Id��C1�G]E�fԵ�0��L�.�t���E�2�.��(��W\��:E��\�
�G�o1Q��t�NR1��������rj�.t�U�bvL���y۰\�ARZ�H��U
��5�]`P{��C��u�{���[��Ckz;��kԩ
����К��pfn�A���B���j�������]��gT�����8q�#/1R]�w����%֐K�;���D��w�*�[tv��b���A�G`벮�JM�u�QZ�ӛ]��5m����⺜ENe�_������0�eмhC2��{c���_'��u�Hh0��;��{�8�h�7�����t�hn��b��o3���ٽ��vZ�R��ۺ�uU��ӭ�W�[Xu��q\�y����[����I���h�^7��iSG�/t��֮��V��bfsJ�lS�s���mU�0n�������ګ�W�'��p��ƪ�0�L��^n&�e��<�u�Ҫ�z�L�S�N��2�ݭ*��.op�օ��v��y���\Os�ݫヰ�*����씺�]�K+�f�IP�'��?�i�W3�=�#w)�	+V�ns��|�
;ٚ�������,[�Ҭ��/w�ИM]A������ۆ��m�������xJ����"��\^sƵ�tR,��\^Xy��F�g���ڟUo�S�P���1�|v�-2mu��`���g�W�	;��v^��6[�`{v����қ|�9���Y�U�c�T����A�Oλ<�ݶ�g�K�ј�ڳ���6{q/6�}�R�t�+������{V��Τ�v�7�!Du�q�ؙ��r�l�;��Nxzs/{i�t-N��ܱ4�U�����+�K+��ۣ)B��b��uš�%qA�o&�kP���*�v���n�N��˙X��ۻ��0u���^��C��V�Ci�)f���X�� �\��I6���5�����޸*�Y��Hnt������ؕ��NԱ���#�L������Y�ن�ֆ�����x+Vu�*�E���l���]C.=�A�\GN�W�4�nNK�qΪ�MQ׷z�VV'[���£I��2�X!���,�.Н$�Rل���[o�3�}�a7D�|���ȷ8�A�D�ÕF����ꢍ�pP���m��{����	5ϏH�J�ۗNS{�"2E��4E���$���u�	(�l��
ªTQl�N�v���h�=Y���K`�4��S8(R�1��\�b���r�<魺�����꽈�z� �����mb��t�Lڦ�#{u�vY�ŭS䉭�s�zq�eY�mR�UD���U�y���;{n{��ɜ���a�7oU�d-E���+�^�Iܝ��H��a=�FN�u#r���w�ظ�ƪ�A��e����[���o]����X��w�����(�)���°�T]��2��d�[�2��v�({ooe�����Og<X2��~.��;��p�TҮ,ܪX�ޫu��ݏH��������zrޘ	����ݭ�,-�f�_��;v��A^ik(�Xi�h��$�I�&[}��ӂ�+r��kٮM{�}�Q�8���ټ�U��u��K.;��`ڵ[�αi����V�G)r�<΍V]�>6��U|�>SgnM�T��c=�/Y\y�����-���+��� �f�&�Z�٫�t��n��|N�0��9����7N��{+��h$țܺq��2�F匒P[W��B3w&��A��ŵ��t���l�.��ԧW�V33nH���]`��W׿i�`�׵�T|+VH�uV��Yq���8_mX\	�+x+��S��ŕc1�ϵ��AG�����a\�����/YM]|,����f���̊����K�4�5��Y��-h���L���
��-�/���j��۴5mLx��ײP�XH,m�1Cn]�]n���mK;gG�{�=�&�v��:F�Β8Us�b^�;t(�nb��un'�7��ս��;;u��ubۂ�c������S������.�"� �X�ʟc�P9�d�kS�]��>�;n�ꗮ��Ҫ\�v�Ud�W+,$㷽VVf��[է$�\��1��{[�]Gt�[;�	�4�nxS�����O�R�66��ڡS����s�K�޸ay�F�.þu���7���d���P���G�7"�sw��ʽ�7�.8��ulzڪ�q�T��ku�&�t7���cfRO���44����;ũ�Y���n]�9IU7�d��w��T�<oNYJ����.����ګm��(wrI�f���JD���W�ol�5��2iǗ�2�US�Ըu�P����-�b��u��*�ܨ7/�+������[�O��綕�<X��P�ù���I6!�Ҿ;�.ﳏ+�ٳC��t�;[!mXw���e�'-ݢ8����	�%j<b�J���T::�xi��F�m`������,�XSp��[++�Cz��ӗ�1������x+F�Čw��<����fI��ݫ�G�6$.�KLe��X,vL�󞪻Æ�D�.�]�w�}t&SK�b�
B=ܚ7����2��w��٪g,lK�ު{��W|��om/Va��B���f�i��v`��]uu4s�x�}Wg����Z7v�٨��}�Sz�qQk��Ϲ�����:t7�"�hmb�D2D�X{��.�ï��jƳ}��{�T=���͈�xeܮ3;3K��vj'%#ni���m}]Dn�ڰ��,��B�f��L�n�xtH2_m.�-Uu!��gc�����`��g�p#	����1��`�YB�]��s��1ɴ�6���I�5����h勪ގ������s(MY��t�ɸ]
c5���Щ�N��ֳ��{�k�׮e)�6m] ��uuW�L��Ds'�/9�y�1n��];����k,du>�%dM�N�W�5|.!&�~��J��*=YՊ��;�H�}g��Y�r�R}f���˺�������b�2���}ٲ���=�pc� _VStܺq7h�|���v��Kw49K��TN"4�77����\�
:�����9h�30U�z&Kc�����K̮82������#�sQ���};�����K���l��9D@�s���7ٽ�t�_ڽ�-�2���k$��h���X���hk����M�:�^o\��M9�]nZ������+u��H�Ȼ��{[c�"\_8Hژ��������ժ�֜9�1�6pmU�;LǕ�2Y�<-��k��v+{�v�J<nS��]E>�]L�|�je��Ō�
��e�Vz�/J�Q�'��s'Н��V����)N��������s�wV�1T����i��0]��qu�+!#�|�;8�헡�㶦�thk$�7vs4u�2q�Po��}u�tUf��t�:6ފ�%����U�Z�F��w�K$�b7]�}��mX4_�6m�j��G�cG}�i��w���TmP}uݔ�DD8�q�5�&J�����ʈ���*[�U�qj��$��U�R�ב�6��c1+�<$��-`]M�u5i��/�ۍ�����PZ�!��l*�kq]��xv�%��
��a���w[�৙��_���O��k�Z���۠���6Ү�s�;q��n���a	tr�Yf�>!���-j�,v
S�j��v��/�v0�C�,��Oj�q�A�rdt�L�j5y�C����W����;(+t��Z���i�����鹎�ڻ=�^o]NŶ�TdP^r��s�Jh9�۸+mU����a}u�v����wX��7����\p^L�P�S#ϲn�mj�3U�{R����Rэ��T���GE��:C���W���rg]�蠮��ô5î֖A��{�gY�Q�2���F�D\�{u���٫6��1���CT�٪�3�w��]��3���D�,�����,¶R7��f_S��z3BS[��ʕm=|r��T�]�SPG+��RS:|Mjb�ze�k]��w#�ڭ/��u[:1�幂�	�N�F�a)+v���\��!N2���)3W�5���Îm��^���%�O�����@I$���߬�cٖ�.���u��F����tl¸�X�,!�MbM����#l�h��6j�frF7@��ñf��&ZF�0�j�"C4j�S4��+�i�M1V�mֆl4$"Pگdp�Q4%I�ٻRa���ׯl�c	�oLV�Zl"P�m5i�K\R����SQZhSg�]��)	l��N�G!��v�����Qص��pR�v�Ljd�k�^�u"��6m�[� �8��U����Wq�p	K�`n��Y��%܃���P��*=+�L׈����f��WbjD�QU�����`P�庎l[�x� _Y�_z�6�\�i�a�VQ���Ֆ��\2�8�]c26�!�i�Z��M��I�4�]6�daU�%�%�DB��׮����Z���{d(�̬ژ�mb�UR6��Єԗ�+1��s��i��-+M��k�K�MB��7d��U,n�e	��6��*�[)��4 A Y���P�k�3uLl�-XP���5��2�4����YR�Y��XX�&����و٬J,�E���@m�Mu���k�X�ˬmj�v��
��+��,��1�LL�+X\d��m��nR���s���mp:۠�V;��h�d��(�f��Q�u�^��f��E�H.���Qٙ����a &k�Á�J��h��&(��H�K�CX�4ث+��*V:��T���j���:ƕf ���ML�I��iB9�m���,�F��
�r�Mf���f�^\�8�$j�0
�qe�G�ZQ-,
�`kI��mVdH×Gnt6f����0-��I�K�]��e�om�k�tt����fu]v�I�ttl���
V;��鯮��&5P��K/S����+P�F���:4
�1�1.h�tU�p�]Mkf֒J��er��qm\Һ٢yP�WYF�ۚ8�zԶ^c��MjJ���/��%!�ڭ��G����j���ޱJ�Y���"в�$���W���lΔ�D�,���[�"��)4J5���hLc��mb�dK*��A�)e6�s(�4���插�#i�u*"­@2F��]L�貅2�/;4��DW`ջ��r�ֱ�J�#���*6�LU��i��4���G�*�M-SmD���ƾ�x��h���,�6���!��!te�K��1��h�K]I�7G;6�Bj����m�Q�t�@�6A�ל��]Y��5i����Ѡ���s5�eMS�a�)�e%�\�"���4A��0٭�jT*�j9��h��֔D\����5v+
�99����
f$�G�@��rM�a��ͫ��sv�3�F��R���sa^n/�۳���(%�6�a��5�b8#�2��k�h�F�02�ΘͰ!��� H�Lܪ`�IaGM��K]�3bٞ�mR"^#ҥՓ4��
j`�)�a�A�lٖ!��:B�ʩ/����ݘ\���ͯ�Z�!��k�)1H�W<��a;V��4��L�P�KJ�K��L��]e��u�J]sɐ�Lu�9�b�`k2\j&8�QVř��\�6���k��n	�o-�Ʉ��m��"K��]cc�)���P�p��Ƴ^�[e FM�b��mV�:�u0�r-�c#X2��Q�i�+����6�Ł3�s�;D�aS1Yq.#��D��e��pK�1���;dW@[�,]�S�M]T�L�k�h���	��l�.ń�v�++�}�����-�F�0qy��3:��pJś�A1f&kj�u.XK�ф��]���Qxi��8Zj��6�8�v�RfS���3b@p^�ذ�$�/Xm�L4���L�M/&�9�cJ1��)-�Vͣǜ�t�e��&Ј[-�P��,i4��jz�)�kuz��-jD�4� :�.v6�,!Q���*]��..*7<,�sLEJ�l�6:��nu3
�X��fn,P�l7c"B2���B���+��uVp�b��-��N��[����q����e5.WW�YY��j�ǌauex0�
��Y���ڍ�e�CR!��75��� ���\2��{!����ljmf�-R�K5��P��iu��GZ�nQ��v�s�eB�f�]�M5&���5mF�m-��6@WhZ6Z4��a�6�t[[f[b��R�Է�)�L��8��n�f�#]��, �`�7ȶ�R®�*A��T�]�RcY��Z����M2T`N�Яk+c	@�yH�ZYRiJMd��]Tfƌ�UD�,��q3\�ؘq�N���$&d�4]vjkXJ�R���Ѝ�"5���w4�Vh�5�U�1�(�l��GF���6��pWlLhi��f(m.�oP��˲���G;@֍��� ��Y�i��hg9ћ�2�^!-�'Xk�Y{l��m�^��6ڹ�̃�-��f5�٪�Jʦc[��̮:�Ir	���h����n����":`,�ڌ2���.5��vF&��uJ�m+�1t6#M#6%��,1�6�0.Z��r�ڣ�K���./Z�
��Yfp݋�͵���,+)k+6����*]\�,!c��1y�b!�.B��Qr21;`Im������Y���A�j9amҹ&��L���@�3�̅��Tq*��W:]/�L����	j6,f.4�	��,�f�����:�0,�V��-v&���:�P�5]2l���.� ��fUv2�J4&�`�ice�[\�� �f��Iv�*�+��K�JKu�&�tX$6������%�e�@�B�ik	�6#�X0�d�L��lmSm.�6V��f�5��m��(�M�͸;%Me�4e3Ld,\�Z�j�q�KkJ�S�[��`��`�ݒ�X���tb&C7��u�E$���.�8;d�E��mX(��4��WD��[cc	��샪�j�jg��8�q�c�6�=e<zkx��L���ݘ�Cl���=H�d������-�]��b�\��RkŎ��e�bٳce���+r�b;[,�0M[�W6j*��XX�b��R��w�l��gp<cXɭ��9u�)f� \�LbT1n�e��{0�#-�d���5�3��G�a!,-K�f�khB(±&yb��)��K]f ����T�MZ1�
V1� JC[�t �B�+���cj椬���ka�%�(;$�F���L���C�J���X���Nu�FC�]J諊6\M�Sb�K��0-�43��ޔ���]nm��[��K���ڄ	V�cn��%�m���`qp�U�fl�s��x0+Xe��n�)[��hkT�)tP`WgTwT3��Y��) &3Fh�d�M����T��f��uB0�N5bK��fr��`ٴ6��ɑ`k+��f��B4fՔ��R�W��.�6��[�A��+�SP�m+�	t�ґh�L7g#M��20v�v�p�������.t4r\n4�W�-�:���Ŏ�J9�����.�m�V����Ȑ����Q���-��)0���:��Ԑ-f2[Etv�: m4P�Y�芵�B�337�t��-S�0o���) �i@�yu�%mR���:c�L�0�f�LBkٵ��/I`-���,�c��R�f�R+�-��y�*h˚�M-�+TѳB2��%6��ta����Ψ�XZ�ە�͂0��l����6�R�kP�[cJTGF�a���8�)^�sf��Օ4�� �D�pJ�q/@��Z�+��kVٖ�ӆ���,Y���0wY�s��ʁsWFX�k�� Zm������JF��v���Z���[c%�X �f��mX�r�I�4MJ](�r��p2�R�]6Ö�1�F���p��h�TM��M.��^�V��1���
V�6�孕�4�ݸXKְ���&ڶ�E�1���t��͕�]v�rB1��\�K�!��MSP���n�[��R����ײ��.�lA+Wr��qS�'aV;]�eɀ�:=XMĮ�X�i�I��5��F�YW�c�Ee��ˣ.I�mv�X��Rh������3F�sr]���a��ѓfSG�\�]j0��.���e�&*ͩn���9ե� 	����-����K�m�Q�
�&�f5Ι01ͬ{SX,���+��a��C.�e.�u�Ԃeh\M.�<`�H�]m-n����e�v����v ZKbc�RX�rZʳA�U�5��f�c4����V��5�q�
Z�v�mHBmnP�U/1[�!1
¸�0Y�
�Ke)u̲��hZ[Ƥe���Tt*���7P��ፎ��Bh%%�U_,�n���CXZ�f�c����{��q�e�%�أ
�c�	7�XS,]����]Vn�q�9b:����t����-����Ĭ�Yf��8��Z�t�s�j9��R��T���c��XU&��\8"�2�����p��Ԁ��
�fڭ&�Lۖ:SJ�N�N��V��2��8�f��0�n��cmÙQ8�eöf��Q���9�+��4"ٶ*d�M�n�cq[6K64R.�kb���e�k�6ŕ�K�45�*��K�,�Q�K(�Kz�c2�d�3̰ID��׋,�q�\�Mdт]2���a4�M��t��]��b�4�uGR�s�t "j+t4��6�Д�K��G:T��h�2�R�g]Q�f��ݦ[3r��k6�l�1++���ۖ5����f)JM��bV�[^���h8��5a���;a�G6�HD�+����M�,u�
�ĶԲ��Xj�&��CWu���j��Z�Z��$%"]�fK�l���B�M���[tե@R�8ٖ���ō��]VT�)m��+mD��-�e�$\]*˘�i(lh� \���5u��R����<�K��F$�R[v�a�ݡ6t� ƛe��lᅚ��Y�X�6�hZF���6�ͪ�b�L"D�paԷV5b�S7Fb�Ѣ����V;GR��9�-���i�nf�Z�+]�o1ͭ�]�1ٺ�yÍ�l;U�J��	�([�|�f�̦ku{S�-�`�o�����mA�'�g@PFQ�c�����n�����8��Gvwd{۫�:C.�!�"ˬ��D�#<���F��'#nmm���;��GTvٵ��1�\m��8����:˲�#�ʌ�ru$SlN��=��n�����C���&nN�ޯ"󳸳+H�mv�e�l�5��Ȭ���8��Qe�ڛY�X^XtDvg9�i�gu��Q�t��8K���;�����,���++���]�G�Sk0����8�󲢛e6�ӽ�Vu��n���8�,�����m���y�YkwvT�{n�Σ�/;�;����y�m��f��(�{W�{l.��wiAyok��8l֫"��gi�i�gNs�彬���!��8:�N���:OI$�{�"�ڊ:isC3͂������s���b���+�&Cl��^x���CL�(��mںc%Zs0�=dnг#�0m�fiZM�0n�T�@#L�q�� 6Cj�.P�0#.�U��5�D�ͺ�P�l��A�[)X�ol�J�e�tU�U-Ś�;m 0B`�V2�V�v�Yf�l(�sR`�׭�L����.6�m���)Jt�����R���YZ��iX���*�m��̴�΍���qDD�m�&ƗR���]x��v�.W�(H�X�`z�G	�fȄI�S�󫢑f�f��۶�УV$Տ#+3�
�aRً�J��(m����u���j&�m�.��nlf1�l#C��l�j�ÌW݋x���P͠MLۉtCnًG��G�fp�ʭ�5�:�u�ե./�8Z���ˁ,r����(Shj�׍G���j��wX�5�&�M	H�,9)
�p6ј���e4U�*�':Y��&-ee�u��]�Klƙt�$��IQ���R0�KX�#�]����E��n��X7]1�5��yuTɥLZ7C\m�L����jԖ�b���탩�����6��6�hD]���j8���31�`�D`� ]6ҖG����*KՉljnƭ �
mv.����U���r��L@SYV7j�ۄ���cdu�f�Q�r��Z�p4JFkK�Y�۲e�P`T�4�B�������\X�$�V[��[���L�mFk0��:j&�u�%�f����cbVd�K�b����7i�f��l�{���[u��W�.�ڢ����u%Z��x��+]h�-`L���Z�lcys�)LYJ�c�RB���Qi�Y�8�Uƌ�e�Xb\�ζYtl+���a�o�FU�#c�an��F`��R�F�ڨĢ((��*�p�.n�M��ZQ�Gb���m��@�mf�ڴZ�B3&���Z�a�V�ˊ��rZ0kv]]2���f�zI$�m���&)��֬$BV6<Ԃ��Ж��h�V�m�
@Z������VEDy�YP��U��N��X-��l���u%m�cml��<�@i@���aAX�eeJ�[+Y�[#�Ƌ*�^)Q��+XIJż�K�B���E��me�H'Z����K�6�)�:U�&v�4�[��1{@�h��%�Y�L���=�f ~|���n���/��<]�I(1���e�r��5��{<.m22PG�r��"�"t�!�M^��S���{�yH��R��v�l�2{僀��>� �:�����[�0�?f��u Am~m���2o`�Vb*��l�ؔ��t����ޠ�n��D7_]�mT�뛕I@`�j� ^���<�K���Kl�(c���@_c�B�^�{�O�I|G��H	������9��.�Eh�l�W^��Y���0*�w`/�=L�t�-�y�-�.�
���lغ+1�f!�m\�����H�g�&���2��L���})�(G���{(�8��Y`�}�w��/̌�;%xWVN]X35�x�#��E�~o��E��|�}��f��-]���ie�|�Dab�L�[��'����>;��A�K2gg^`�v]�t��;���V�˘Y���/Wb��򙔉V���l��isA\/����n*�a�����!���v��e׎��� ���� ��(��"�/�%�eп+�u6\����	���p�'ޠ���������P�
�+M끆�F�#���.�ۻ�}l{p�#��F���W�V��/����A0��m Kt��I�
��UD@��P���xk}q^P�gި��GJ���ht=\���S;���q���#��:A��еSA���2�eٔ�`� &c��R.�|>�zϿF�>}c/�c��m����������k�Au?k�k�����C��n�?7A����*Pe���ă�4�?[A}���[�����#͎�^�=Ԁ#z��;,�%Gn���@��Fec�� ����n���^�����o��+��fj�Ux��y��e�X��n��Җ��c���c�<nv�d�N��S���~�{��W�Z�ݵ{2����Q��Zǘi��yWi�f�/��~�?6�������O!=C	��6�@�A�H~!�Co7%]͞��^�?z���x�9�ʺd�����H�/�-��?7��tό����=���C/Ќ����D��D��۩��WI@�^	�	��X�[-�e̸lq]T��k^�H��J����M]ފ����}�GyE�9V��C+��^��}v��f}���u��s�����Ќ��,fz�q�9e��Z)�T����0�3m�1 �B �ͅ^�{aL���}���1�}�PDy�_��rW��{x�	�/����� Cu�n�ϛAz�b&i�UO=q�cwQ83'p�l?di] F��n����Y�E�U[�B� �{h#:�M���z��]��W3>���u"({�a�{~����CS��rYV��B~G���&j���;T��t�)����ϲ\�v�V�c����RhhxX��w�������A�Hn��-� �����ˤ3�r+��qk=���1���ޠ��΂-���CE����C�[Hp�hJ��uwWvh_к63�=m�����
�5u�1��b9ʭ(3^���)�������h!Ѻ3_�N���"��^#� �S�ڄt������/�m @-�@��g���P��R#}AR�o�z��OV���3� A���vc"U��E��҂� �C�@���H�Cu*��^z�OK��;��q�;�� ��>�~�A�"m���3���&ckA|~z��p4�9��_�s��vJ���W˳3s��,ɃW�~�y��Oz�Nr˜���Qd-��^U���}���Aj�g;�C���z��ϳ|�u G:�~m��p\�T\��b��g'+�y�r���'�t���1�N���8}�R�u�4CC�v*��9ޣ^���M�P�k��knR5V���肯Ҝ�����V��Fʰ*�5WgM��kJl���4�GQ��F��l�f+c1YWZ�+�X��Ք��9�+��1�ib[��t�E�E),�a[�naH�K2ŷ.!+bX�l�2ն��Ͱ�k�(�n�k,ey�Be��t�I�^�rBk�BK$ұ&��U��պ7��Lj�r�46ک��s[`�*�1�݇gV�6cT����5�?'��������[j�cM����[���#Yb@l�,��S1Y�-M�����K�$��n�������;�E��0@1�}�e��`�J)DNrˌ�,��U��7�_v�=^�?31��/�4nks�k7��#H$n��"�{����YO-<�1����=� ��"�"���W-����;���]���>��@�:�sA�K���*�'}|�1�ۭ?�Yd{ڴ`������g��Y�����^��~鋫��(/����n���@���k��+���O!��;�j�{ӿ��Oz����*�"s��]��o_?|�K�e���GD :���Q���"�RĥԴ7$qŚ��Vo��}~Y�q� [�?6�ĸ{���]�[�gپ�(�q:ݮ�Ax�g������!�@�{=U�v�p����}�ßl���y�ƽ�@SU�j���%]VsR�J�Mgy{���x�Z-����k\�ʍ8ޯ^���"��{㒐5��=��W.j��`�c���P@�y�@���a��x{�kf ����:���k��/�hEw^{�,$��Kg|���������A��z�b�H��|�!��5%A�����Aҗ�AJ��uz���3�� ~u/��F؄]�կ���PE�DCt����ָ�͌[~�Ӹ={oW�j��`�c��P@�y�E�D�Cr�k>��YIU^�R@�c4ƊM�4�m�r��.���1��BR���gkD�l·�?y�~��>|c{߶={ݠ�n�./D�n-��F���ԋ�ReP�"���.R �� Ci|��x�H"f.>n���ۜ�4�u��3��	�H�t?6�P�|^n�?Vb��k�Ct-� ��k��e���8k�r}|�U���Rĺ�k([��&�<��9���Ⴚv"l�|�`&L9�F�ӻ�(��A+��Nu@�L��)�8 �x�󯛬!���h|�/�]�o�A���h/�ۨ�A}�w^7���FCLe�{�	�"(K�e�~����H��!����~n��=io�<�C� ����振j�Ԫ~9�V��/�"�~��Ŵ/}���l�=�.�0��*�زݡ�l�!/
�q,e4�]��)p[q��j��\AzR �A� A!�C��1����\��8 �����]�=�Hn� �~���"m~m�t�#�.�<�0�P?^%�h 4E���U�U�!�2�<�=�@��-�Ϳ��K�<�ۢ��Qb/9Eǜ���͵��6f���d�<�moa�n�/�R ������_��0�9R�3k� �_7Y����1�w�=e�~@���C(�gz���E;�{՝��/(A��|:����5�R�A�F�{r���3��;ݺ��� ���}Z2R)���
���u����~mźD�G���4�~����M���[Ks��\#���z��"�"	���ϯ|��}����>������Z(� 9�h�6�bd��D4��SbdWC���e���=�YvP_���fU�L�����i�n�/��Or�e�T�?���_��H|A!�@���0l�^�m|�r�݌c����� < �� ~�_7IS(z�G:���c����_wS��� ~m��������m>�_����g.�A{ԁkA|t���������jt0AΠ�<���}��=�<�<�{�g۞@�gR��Tz���O��?gW�>A|[�$7H�� [�琶�N�[��|B�Q��s�S��͡b��}ޠ�'�[�A��cqV����Z��<�5����n�u���śf[&+����j��K=�/Օz*���}��C���8(r(^�N��{�vn㯓���稲О�SX�#��^�d�ݝF$�F$×u.���Ѵ��� ���-�q]lڡ1�Lf�75E��l�iV��(��k�lit�Y���g��j!(GW��nvjiKԈ��6;].�Wl�4Nhڙ:�)V9�B]�S��CQٰ�҂ڐĥZ��!�X0F��UV�M���e3l�-��D���ef��KK��X�͍���'���aS2�P��=����n+����f\�6�M2�-��V(׾�����������~m/���go_v~�W��{�y^������&gۙ��5��H�Ct������C��7w·�����,�gzV{��왪��Ϸ<ө�_�x���iןu���$s��m�n����ͱ����d���o�͠�g� ��y�E�@���7�EU':����j��#��Ŵ#;��q��3�i�~� �����
�s s)Hn��6���@�[��-�J���蟉����ֽq{z��d�W��}���3�|A���}�6��c�`�D���T�����F�*�
TƔlһ��qAIlP�!�/��d�Vj�l�[���!=�~�t��n�����n���A��u�^R� Lp� ܠ�t��G��@�[��	���P��;�q�?���5��um�8��9��hoUWa�����e�x���������g�����)�]�X�i�����풚:�?N����n*v�Bm�;�h ��R�@�YL��f�)7�@�w�"	n�-� ����g�o�7��H�;5^����'��#z�����H���q�׫$M�C������]���}�G=����{6��x�� ~�ޢ�*�g�� A�G��@�u�����x9:�x��ߕ���l�����ֹ�{��{���[�?�Vu��D�׽���l�H�B&��*7lܹ��4��r��nm�)Yo#a*��:7t{�[��DgPE�@�����^�$~��W��}~��y�	�CF��!����/�m|�a�Ct�!�����v�Au:尾6���7G�o��ݞ͠�%�~�A��z���ћ8{hC�b@��_m|��-���д��I�ܾ|q5UX�U{.�{m����V��w9^nL�9]�֧J�a��d�Fa���)]z\Ϣ���3J�(��7�DU�(�ڲ]%e���d采�T���O��"8�ut܆�_s������N��Z�9��sX���27H����-ւ��ˮ���U�
h.�rw;��3$�k����J�W��}e�8j��b��3�t�y��K�sk��(�bB3�ݭ��̮�������ox��ۺ�Ǜ%YHM�뙙��}ɠ��.�����y�x7�=�Uf'�7�w�ȶ�X<�*lZ�^c�غ�F����&Iӵެ�:��a=�|��UUȃݩ�MU���J����7t�j��-pQ���kWp�me%ܮ�U;������$�km����';�\n>;��Gk�W٬=�˭�3^�Xi��b����oO��z��a<�e��V�R�ʩI��ou]�n���>L�sz^u��eP� 2����w2�*����v�|�&�z�7�.�t�޺9�ή����}�l꺃�Q]v��F�W��=���R�7����o%��ִe���q�����\v���s�a}Ԋ�g�je�bx���,�ή���ꗀ�0_U
�A�T�J�W�G�m٭5�Ү���¬�j���	7%oZ/C�/\���5���zV;�l:ѮH�<컳����S#Ydf���\���M���g�s;a���5�W[��:��4�jT�[w�34�Cj��9�f��6*��J'����/�~?s��ufEvGEVؔ���-�6�m����3��<���{������֎�<��w9m�,�"���;$�6�m���m�����S۹���:�,�:��M�Onħ��Am��3��uOk�mVڶ�{�wzQ��gQ�T�gfgKj�8�ʌ���,�{W��^E�[�Χ�ێ�����mնH��ygY�^^s�q�T�m<ʃ˷�YA�Q��m͛t��ADFu��Q�mk2첛t�H^6�"���:B3NN�N��H��I��qDsn��ˬ8�GGDqE�v���y�ۄ���D�iݶ��μ�O0����(�8������H��*��fu!^Y�ww)�Q�y��gbEr[=����
J�x���Y|.wZ��� �A��@�R
������Xh�\4�XhaH�ZM!I �e����XfPl$�����t�����wD) �W�P- ��)�~�ZAH(i�4�Xh�����~���}��w��ߡԂ���i ��B�	@i�|u��^�G����	}���� ��B���H�Zi�)��2�ZII�Lˆ�
A@̢�p�mv�l�����_ �G�c��^���8R���I �{�- ��Z+٨�SH�2�i �?3 I~��7�"��[w�0��7��\�j��g$2l96��c�655��M���KՕsW���
ެ>a�����ܨ[&�) �Vv�$�H+�p5� ��fT4�]{9��:����_��־�����Y��j���ik�hr$��ݸi ��;�-&�) �S)s.�j%$���
B��3(���!I�ׯ����f���
j S��i�� I6��'�"��tt��gK�S^��:�W7a�$�þ�ZAH(9�4�R
A\ˁ������?_�R����`Rz�M�YC%/ݸ��%$f\4�XhaH�ZMRAd�R�\]����p��(�*}��i��@���H,7��$�@w�- �Q
H-B���i4�L3*���P�C2�$�) �e��i ������x�C�7ʅ�y��P3(����4�W��MQ �C2>G��ܼɷ�U�=Ց����i e@�� RAe��}p- ���᧗�y콉�hr-��|s�aMqm�`���V�u&ggmT2Yo�滮ѵ(u�_gV��S���zo�ۻ�s��Aa�aH�E��B�%)�*�j%$�t�RU�E���]�I4�L3*�	�~3��CWR����m��Me)��� �G�}��n> +�X��*��9@���u�pޱb}�#-�&J��A+4f2�Ixu�f`D �1�i*�����ݙ�(�zMd��=��BΖ�2S�TCBJH,(��H)2�H)�q��T@���ߏׯsst~>>�ü�ZAHk5ﾢ�Uo��E���^w.�
i�gj�FJH(�ZAa��$2�ZAH,3*ɶRA@���U׫?}����Ă�R����
A��eCI�=���;���+�s�������->@���_}P-D��XVe�I����E��c;}�p1 �X�wʁh����AH(�- ���TH)�eBك%$(C2�$����*�o�޵//1�:U���&r>
O���B�
A@��Y����I̨�RT3*H.����-4�I��������]��l�k�W�~y���II�2�i�������B�%2�ʁh��|n��o�n�Ǐ
Aa��}$�J�;��R
Asj�}3������W�q �D
a�uf�JH(R��$�) ��a����)�eB�4�H(�f�
AH.e@篮�{�]}��<AH9PתH/�9]=��[wmV� ����2S���%$s.H,40��-&��Y*2�ʁh��u�Lo5]���@����^���(�GX�/�7I)�-$v+T�+�w3ͬ�w�6��sၮEn��_��'ɂP�r��m�)uvf� M��� ;)STö�K[�7-��e܂���6m�Fe8�Gh��6mfq��F�]��lxe���H�9��	�M-۪�k��sXT��4��3Kt5����*��JE�4�Ժ�a��0��B����co��0/�uؚ�F��Ҕ.GV�.h�V�2��F�t4	[�20u���M-A�Mfɬ\�3?~>����F�).�lF1�#u&�kc]iVfd����K%FR�Lm���N���zZAH
�9�- ��껚�i4�L3*�2RAB�3(�A~�3�i����_��4��&q��$AI���i�i�ߪ��ۨ['�RA@������Is�F���h�fT4�]0)2�H)�)s.��RAa��w|3���Y�é���̢�i
H,��_z� Hv;��]uÇG���8�$�����QiR�RAj��@�����2�l���U��/{�&$,C_��Aa��$��44�RP�0�jɦRA@��4�Xi �e���RJ�eCI�C��|%9}U,R��j�� ]@Dp�I��K�����
̸i ��aH�ZM!I��)s.�hJH,3(5$��֯��+tZA�D) �W}��SB0�����P3(��õ�3�}������w[�?>��
��i ��j��) �f�����NH,4�W�\MQ ��T- ��-6�I�2R�\CI) ��2�G������ ̀���{q�|������:�Y:�]�����u�����7����� ��(>t�RT~��
AH+ܸ�Rʅ�) �B�i �ｭӿe���l�ת�a�	��^P52 �֡��]oZ�+��-c6e��U��סIw�i'P�eB�5I��f�CIs.�C�H��G���Vog�?^�Y�|��stZ|�I�羣�������uv�ZAH,0�.H,4>��I�) �S)s.�j%$�H)@fQi ���Ͼ�F�P���M���wǢ�&Ι�L���I>j�na�4:66�8�ݙ��ҷ`�^�����Yԝ���U���B5�3;�3�+�5Z��D?|#�H�@��B٦JH(R�4�Xh���OV��ϜW�O|4��%���$|	 ����R
�z�$��
�\��u�8AH8T3�$L
@�h��@���d��n����XT̸i ��
@̢�i
H'������u.5;�Tc��f�B+�����㧅 ��*�R@w�- �RAj�5�
Aa�P�m��
�eH,40����a���]�_3����t1�=P�Le$
3�i �4�A^��kTAH5PfG�H�6�"����)w��s}��*����(d���hi%$���������}��0���I�
H,�K�\@�JH,3(4:H)2�H:(�$���H)�
a�P�Wu�Vk��d�H(y�	#�O�ue���s�d{�'�G��\H)>��ި[&�I�=f�
AH+�p6�
A�P̏���&ە�+]�`��W�Ht�F[�kX�`�SF":�V)�dJ�e�GB��+5[�Q@���H)�d�����%$g�$�)2�I�) �̸����\������描� ��P}$���/�����^����D) �=p- ��)�r�l�2RAB�̣I �̰�a������H)]w;>~}o�O$�
�.�D�R>��>�fy-���+EM7�߀d[���
H,�������Fe�I��Re�7�.��f�k~���^$K���.�i) ����R�ݢ��!I��5�
h@��f�) �B�i O�!Qrxv��j5���E��1��j<��}�&nޣ������u��[g#峵F���V8`�j�fr����tVּȰ�1	�/�7���|>o*�]j��jN{֏|4��%����%!L=ꅲj2�
�4�Xi �e�֨��h�fT4�]
@̢�B$o�����߲N�߮��JH,*s높
A@��i �m����4f��;�Z����<�����I!U@}�- �Q
H/�{��\�w_��տ@��� S�B�
AC@�r�$��W2�c$�!L3*ɡ��P(̳I�������}���7����$|��z>G��얖�Up��SO���@����()~��Z�) �̨ZAa���E�Ѕ$Je.e����L{gSu{uU���lb�mK��PZԖ��kHǭ1is7 ,�X�a�<���>�I������@w(���!I���@���)�eB١��
2�H,=_s/߾��s����C�{��ᆒ
M_�gݮޏ��0�T-��) �~��H) ��p- ��C2����`Re�@���W2�ZII�r{{�{�s��}����e�HRAd�R�.�k9ιߊ����9�
Aa��ZAH}*���ZA����fj�� Sʅ����U�������7�4�P��4�Xi�$��40�AIB��[&�I�,�A`hH+�p55D�Uʆ��]����w��߳������Z&4T��_| 
���q1d|.��v��V�����L�sc��l:�����Ø�TT?�h@��"5����:op�1���?�ez��D���.�f<�f�ߺB�SYh�qoX�_.7��4�Ԃ��<*;!��R7��?� ��p�T�9��r�9ʴyh#w@]Q��R<�l���:ߵ���@���[��t�-��-��^j�J.������]s t2H��nu�tmS4��E
FФE��R�q�!��������Yr��9�-��W�5jf�ժ���N�9�q9ʜ���y�,�a�`�r�xp����6�K��ú�����@�_�w47;س�9��eg�C�"h t� ���Mn��2L�A�����F�Uc��n� [��k��&g��Z��� ��u|�ho�����L�Ҝܯ	�/�����dޞ
Z6�|A{Ԁ!��-�D[��uK������F�u�,p�kS�6��f}ꊇ�-�����Ŵ-lw~�Tm⫬�ay7�u�����֖w��zs�9�_>���n��;ৼ��pnWQ��ڧa�W~�n|j���H�m�������>��O���.F Db��X�R�.I�ЖB��+i��͔9���q	Nt���Y��+Q,��vb\�\Ɏ*�T�V��6�AF5J��fHD)��º*�Gn4ғK-�l���Nx[i,��G#���ކ`ؤ�S5�^C]t��u��Z֚�ؠ`һ:0Ű�\v�B�aq�cȶ�9���v4 ��4au���(Z�)نvM\:�'����^#Yu�D���ka����:��	l;����Ǝ&f��>��Ye�>��� �t�$7K���+7��=��7h\(m��MT �g�{�v�?]��?���f^7������p��W2�S�+�z�n�n��vp+�_�����6�%��[��-��-�k�7y'�zo�o3kj}� ��ޠ��������@�溔��-�7�������-�Ct��7��[��F�U�^�@��/h9ܿ ��_�] ;�����H��m���.�7i�J�߶m-���\��N<�|�|�A�|A!���x��k������_�Bѐ��4s�-dɭV�S:�[�M�����hScV���=}�[��(;+��!��g>̩����^iڟE��U�r�z���|A�A|~~��h"�"!�G�;���\	q�U���;!�Λ�^�������뱦���U˅�nUa\��mξ�����,s����}[�0�3A̪�֣)�^�����|=V��k�ߝ�_�y���0*��6���b��F˚"����>�/�!�?6��6�����g�1� |�gd.<��G�_&�E�D�|Ct378���=��X+(x������o>̊������mO���� F?w�j�������A� ?�/�-����#�3Vg3QD�];��W�{̳�<�|���?s��u�m������χ�>���!�3�̦L�*.-��C��W\h沬�u��`�J3^���2����{�2��|��#λ�<<=L�Ǖ��wf{�i�*��_g��;ԁ�/�m ~7p�Af�ϡ���G΢�h!�Z�2+�{�_cѵ>�� Ar�#z��RU�//?�âԁ�)~m[��7V9na[�q�SB�.���=lop�:�oQL>�VeuFn���\��]�4w_fS�.Y���Л~in�:�Y���&D)W魍� ��R�M�ǫ]�����,c����yʴ�(��r������{ �J>����}wі�v��s;arex�G�H��ْ������R�7�q9�,c�Qq�*q�Kj�X~��RT7Փ�&�{��_l��}�%����o�������]F�=�������16�0=u).ap]1F�4�em¢SA5�R�,b�j�ټ�_� Oz�C�昷H!�A�aΫ���t6ǀݯ�}1^̾���@�}�� ��G��@��7�E+Uf�_�L�(!X��1�e�Kˣ����ʭ�bB�!�@�_k���u�u�ChD��g�����w�#�d��}S�|�"4���_�|[��\G��W[��`����A7K瑍��Y�n�T��Bp#�=��C�.��&�o�����`���~�6��Vp̆�9`�,�YT�����T޺�9�Ӯ����P9��$��3�}�danT��wE^㣥�~���Zt}$���G۫�gh ~m�t� ����U��`H��q�l1�|�������A!� 5h [�����*W}]^?Q�D P����)c���%*��1�5�17ki)��U��=ޠN���_7XCt8������M�k>�ЄT��a/@��(7���i|�u�!�C�!�{�o��U}�@�y}~��J�=�@�V��z� ��A�|k]����@�t�!�����T��P���>�^�'�w#�.W�w���u��Ct����C{�{+��'v�>�"mվ���]7CS�@�)�%f�����F{�K���o9WNr�9Cu�h<7�/b eV��oz���<��x9�X��E�}��W�"s�2j�U�f�~$�V賻"�w1�V͎r-�`��r��i2e�;bm�L�A}t�$�[.�����1\�|s����!��u���
�&lf�;7�R3��2g����uA*�SMQ@��R���D�Դs����;��\���񥹗��\���ԍ��z���m��W:�|f9ҍ��G&ou�ŒB�nRe+;�=�],��0U�J��&��7���9Qә2f]Gdwh���1�����
�GŲ*��y��������L �gA51ve)w�N��-�&]���ܣ[�����Z�U]�7x�:�2t%{�z�r�[*��[��!�W�*�T[K���s*��ՆƑ�������c9�ݭK�3�9�YGm�{�aul���r�Z]պ����<KJ[ל���wN�L�LܫH��Ԟ�yҪt�3�rq�Jr��cW�)uu(�oP˦��W�V��w��nW�:�#6��,��3F�S�.=;w�5����
2���E�\x��77�m�y��_me�]�uԩ�4����1Yv���Q;��wo.�]k'��LZ�t-���y��"Т�o=�Zl�v�2z�ôt��e�j�:f^t&pݷ�N��ew�_^^�=��N�7��{��C�U]�,��\��9�	\�|����Z���X�]��N+��4��+
=��v�z&操�M�36
̾o+����i�]��{�G9V^Zɘ^���_m*jCz^��I��m]�PV>��[�j�8�X}��J=u�k��'*�v���Ng:��/F��̻Yͪ#b��	�(�������f��}/��R����l�*J�~�k��muvۻ.�%����/7y��RNq���"��B���8:�(�+�;��ʼ�N�.=�uޝ$%Y�]�\�]��wǙErOkίo{����
��:̬�˻+�9+��ݖwG���.�';���������󳢊r⼴��(8���u�'QDtsێ������ӹ;��L�9�:���Β(�����,�(;�{]gvvVq�%$��n��/:8��yn��̨����t]tvg]��8;���wIWPVwY�t]E-�ȸ��8���N�
�����H��^yt�pQy�E�TuGvێ�볎�8���<��J�;���~?3����L�썆�R�U�@���N�vs[�&7\\�8��[���Q��e�lvn�:��Mښ%�����q�+b��'�]O)Ҩ3Vݠʢ���.5e����\=�і��@�v*MQ�(L1��6c�����E���ִ��3I�Ų�Ch�6�"�s,R��&!4��I�Fca���2Z��Ի8��S.�Xl�-��\L�&`CV���e[z�0i�pF�,D&�Yi�e���Vdt�][6�ePƅp���6��֒±���3�9�C������G���7�֖Q�]����v����1�WC\��gKjLA(Q)(��6��ƕ�%�Q�M�ʰ�uCDm�oVݶvʸ����2�%()�T�u�0�6�!t��9��G$ZE�����ш5F0����3��h��Z���4���U�j�ĥ5�հ�SM���.c�Yp��i�M6X3a��5��c¦���L�1��,�F��a�l��a�-o+���Bgl���u�lH�貍�F36ۤl�Y��
���o7��k{4Q���M\֬�Z3!��,�8��p�++ea�u����c#Ef��m�tm2�J�����NC]&i����͌F�5p�Xi���-3�M(�Yib*����]H�]L�v(B�uår��Yc��z�]&���<� 4���a��X14ۖ��TIk� C"�2$4锼�!dɴ]���!�3m����v�Jb9��h&�&��bfQ�OP���.l̫�0�@����4+h[+qiD�aYN���G4�i�,�mK��\�W++�G�cUԳ*���y�ݥ0](Sb²��\�s%�`
�Иyqr��Z5�8��f�p�����]�[p���%CS�p�[�c6f��p��#66�[[���� ��ScLX��Z�7+�]mv�P�V�i^m��Yj�D��*Y�
ښAY�]fՎ�uB��lѩk���+��X�]�`��W뤒wH1�m4=�b0�Q��Wu+�q��]���`��������^��F� �m���iWd� �irlČ��2�Ʀ�@M��l��G�ఄ���WG`�!�dĬ_{�Ob���l(SaP3	��ˈ	Smti��HݬXX,6�..���cl�"��ZP�2ʤPxˊm	�mcJ�*lư�6"G*�zل"遡��+�����2���t2�V3KY�GTΘ�F\���^^RXf����a��:r��/_>��� ~m/�͠�����c��qt�r�����[F�{���n�N�1� 7H��[���ۄ�uW�+��^����{��tE>��\�<�G��v����=C�R��Gz�A�n���n�֯W�)�^;:aM�3�l@���_7X!�?6�]fn嵵����2 ����h/�!���x�k�hɕ�� E����e��.����)���n�@�A�9�nf�������=��"�5�	r�o ����C�;�y�\��C��Yf�&a�T��R�\�n�-5�J���lFQ�ssWA��>~>Y}c/�c,���~c��<�� {��l�3ݯ���T���_{՟Ch ~m��_?Z�˗Z=�W��;��s�x�YW���2��az���=_oAMs���w�.�y���9z��V��,d<U�WI�uZ��gwѾ~�qެ����I 7��~���@�Oc�s>Qo2���}�=�AZ�[���N��b�)|Gj�����"hk>]��i���9����%O�� ~.R����!�ź���{ؙ܇�9�ic*��@��	��1�<1oO3���=�_OPBW����u��g�]wtX�uq���q����H���۫�-�vH`7Uxw����ؓ}2� �� Aւ9W�9��^�k3�y��uъ�`�c���k[��(�KR��a�s\�tXD[m��K����b���z�t�-���z<��{�Wu��gՔ(d��@�n�;� ~q/�h"� A7H���:����/�$w�|3ь��zy�/�>� oƜ�2#[Wq��I�C.���,.{�i�Q`�r�!�Y�+���~�a�4�*b��*�/2
a]oAtEY�b�̭s��B'&�:�^9�eq���"��ff\�E�U�a��^�]c���yֺ��^�w��s�D���ɕ��Gz� �A|[�A ����l�*�:��A��W���m+}sz��ʺ�w�e�H���~�Ҽ0Y�Z|_�GM@#v� �SY�fX�A�}�-���̋x8�@�=A����B�k�s!������1W��Ҫ*蚫��,eM��+W�uΡ�:�Xgb��r���D+k�s��W>�3����Yr��r����-y�ё׀"�o��yQ�����A�#�H�Ch An�"� �W�NryC 7��}Az��w7���X��>�h��~���sC�0�[GbR����@��R�_���z�>����ʰ���~��̄�pk����C��H[A ~m/���U�������w ��r_�AU��ü��GFG^ �Gz�-}�U]�Z*��xИi�I(��\&����5*�nf�,�ڲ^���lH��Y׵yjl2gfQ#�����W_�����A��ʵ˕�[�2�K���t��ʖ&}S��b<���T�(���M�8 G�"b�G[��wQ�����}���Dh/��k���N�|�yvf�2�R�e0̃�w7b�+�]4 ˶35F\��YV39��7������B}�i��"�7Hd����Є�p|�B��ֱ+p�^��A|zR�G����DL4%���Ue��>���
��0|:;��*���@�R��t��T���|�W������+��x�� ��/�t�!���)^չLk�;��N<���>�z�{V"o�X�r���Yq�*Ļ�������Ԉ?_�_"!�C$�p���=O ������#�ދ'���t�JDy~n���m��OL�]���qx���q�g|O��gCRJ� �Gz�Z���Hn�����Q�F���r:��	[k�z�V�=�:�M�R��Z��*]�VSԆ��ِaCH�e�����ݲ,_o�U:�~�sY�?HHI6W���[���ڪ֪��6Tj�	3����u�6��x�3u��is6��	0�h�nbR�4���lDe1���uiI��)p��\lEU-�5ՁM�v�"ڰ^ٚ�i�Z�c[r�m�*�Xìee(��f�tEi�0�.�8�6oQ�Q��ŵ4�E��ؔ��9��`��nf�Sd昧�sq�t��c��H7l����tj�X��u�_~�^���.S�04�����m��[QX��2�v��7kB�-�8�t�2ߞ��'\}w ݯ�o��Y�B��ϢuɆU��y�B���C�ޯ�͠�t��f{��������K�	�!���p9�'�0p| �P@���H���}�<�K��ՠ������"m~n�M�}�ây7^�}H�"oe� �}.e�5$�|A#�H���@�����p��;^���B���_S��.�Eӧ8��	�6s�[���f<��%��g�4�3�"�"	� ��h [�*��������E*A�f{�oI�EL�/��/��("�/�l����}|��˯������������^1H3[]5&q�PN���Jr6{hf�JU����Bsԁ���|�h!V߽e���_CRJ�g5�Kڽ���OcBu}�l_7XA!�D7A�
���8�d�_v��9�y�o�r+)s���g��uP�z[�ڶ��V`��:�n��-��}^�^�f]�Z���z��o5u!wu�8����@�����s��>p���g>�Ё �� �my<s�5f�'��$�HA�mn���ql�a�<ǲ�w��w$��*`�� L�A;("� A�������쒰>�ޯ��|6b���m�����~�2��W��� F�����Cr��� @����-�_���u���	�E�qf��B�s^�o_�$1d�>����F������
���A3o<������2��XݘL�	H��fk`�]vb��R3i�e�}'�e�|�s��������\�<��wU��{������YA<�"�|�h ~m/��BX�Qo+����_�*������~w2��W� �ޯ�ւ��azm�_�m�v$	�AAn�-�@�ǅU�/eX��.RS���U����%��9{�]9��Y�.������r�$5��Ђhj�B�ķ�qX�3��}�nL�Y[NsQG���}� �l���@/�h [��?_oz%;���Hޯ�VHn�)2x�=�U�+�{����t����~ʣ���#yK���C��i[��͠����{���g��
�k��#�|���5#�~#�H�t-�Cu�s���|I+�ё	�2��3F�,�CҗGj欪Hk��a2�9,�T�/
� A�P_A��-������k)Ӝ�Q��3�G�:k[r���̞�E�~|���@� @n� �]����u�"�Y�r>���Պ����3����c��gU0��s�R ���_C�*ٞ��<�er;'.��H��;Ԉ#Z�H�m P1ع�EY{B�&�;+���'v����GN3�� Ou}]Z^��Լ5���h��#��)��C,�<�6#�*	\:	[�9��f�v���wjF)�0��.�\)���Q(e�R�ei�>����?g �?���D�!�-�fy���9Q�7#@�N�xf��[�,I��~@���	ޠ�t� ����?���i���6��P�-�G�XJ�7]�maKT�k�c[����gZ������=�K۫Gܲ�s�.<����֫?qN���׈͵��U�2t�b37e�ʱ9ʱ9˖#�Qb+��6��z�r������P@s��غz�8�q�Vx	��4��E��/Ǭz����:/�� �G�|�A|[� ��=��t8���Ʀ���ujԠ�u �P@�H���7�2]ͫ/z�m_y֐{G�D��<�{C��U�N1Y���77����ϗ��6R6�@����"�T�ܭ�+����v��gOY�k'�g� �R ��@�����e�e��^��_]i��pu�����vs�� !�T���>F����[�^cڂ�,��Y��v��q+\U��^�,B�hw�$����ղť����j�ZR��������4lnu�`�vmY�r�kprmP��Mv�+Q�e6-o9�eeɬ	�&��7���ԍk5�]t-b�攗�a��EpZô�����m�0դ8ض��@��B�d���±��m
hqr�V�E�r�q1n�JE��X)�;6��@���Մ/AlJ�j�r�r�EE�뮊4�A����U��_������x2ݩYb�k�U)Xf�h��αMe(�h�mP�cׯ�Y��{��-� �CuqI<�����R�;hK$+���S�P�A9���D�@��@�� FVp�Z|vh��`��_/4M��5k=�:�8WG^;�����ηޞ��k��i�	�n��D�AW�r�heu��o��|^�d����g՞@��D�~m|�-����G�,�r����|�` 7Hg\�˶���2*([��h�q�59���
v� ����%�@���۳�/w��ڈ*��;��{|��o�H����_F��u�t�:��kA��6�}��,��1��cM@F�,h�K�2bkf) �b�.�N�Uz;���9E�ǽ��r�D6���mL�0���}Y�*���Ც��\=_�K�A� A ���dn�b��{r*a���ȓG6���(�2�*bS����
^�e�ɛ�����n���W�D3�Q�AյC'���k>ێ3�{�3#��٭�dTxZ�9�Ӏ�7p�k���0lп���������-�A��"G�ާq���o�ؗ�*G^ �Gz�Z�H�7_7�j�ו�Ҕ/��u}�X> ����9[t�6�q�G�q��k���U����0�4�#�n����h [���K����K�Fz������0n��u�/�`#��t���9n֑����q3m-���&#�Un�V6��E�bfJrC�yP*�_UZ�[���/����7_7A�ܯ^�S;[u#&��̍"Z���.���U}���/�|A7HAt�Y'B`�!����@���v�ח��n�d�>����K�@��^�.էۼ� �R ��_7C>-��n�}Y��w�{'G�H�����{���-��	�T�U��Z�,6�E&J��m<�'�z��`���U�����a_L{N�Q.��8��ˮ�v�:��׉2�˳Ά/�x׫����U]n�#�ˏ����:���3wGrw[j^�uk��񪕱qz97�w(̒�9
��뚨����j���Y�u�<�2U5���l��!^ܐWw���.���\[z�ş+k��P'E�$qZXK�sf�w&T�꾫i���͝Q�ʺ�����t��o�%1�K�.�Q�r��������ɳ�����k����zm�I��a\ۯ�:ِfV��9�D�(I:��w#l�S��T�_	׊m������Zy�r��T�1�^֫���b�Qu�f��Q�R�\�\���v��;F��g�b��']_Z�rIc�B�k�z��07��}��ԂY	lɛHȺ}"��gun�3�;C����c�n�}U�L�]�f�bS�tĘ����uZ�N���؁�\��˻�m��Rʸ��Y�,R�ޮ�Ey��[�4�4Aun>J��r��Q�/����b����7�=�w�I�x:Ѹ��B:��ɇ��^��Ӕ�R�)��%���u���I¾�y��7Xx�ޮז���y�u�X�U���.����4$�8���--Ӷ뫎@��E�gC�A�|T�fQ���˙]���ƻ4��N�����r�k,��r|��fZ���i�^�Wp��u�u��ʘ7�R�nL�.��{���T¶���]r�u�>�rf�qf�I���ٶ���sl�K3+��lf��ս��ߟ�����P���N�⋸��y]��Ywgf�6�/mGw6��.��#�8���;;�q/3����2��H-��;��.(N�/mw9ܒn�㊈��J;�D��);���qQp�vY�tT�Yl�ie�[h�F�VS�=��㓮(��쮰��Y�g�trW�ŉqu=���4�)�[�Ivۉ��wm�έ�gy�gew�ΰ�����"+˶�W�]e�嶣���<�;�������u�$�XZq1L�� w���K�$%9����#fӏ6�o^�pD�%�Z	�vU��è�#,�3�%!I-���`����ާ0߳[�7g�:���뀈 Ӏ���� ݠ����)#���q0+�F��������q��-��C|�G+���Bvc����jw���Ns741̢� �A$^�űS~����;���f_������}[_I���~��BIay���O����Q�X�p�۔�[��+�-Y�u�Z�	���������6h��~?Y>|?}��2R �D���_t<<绲���M�nz>�מ'C�A�PG��dIA�A�+ �)������}��5z<��_���L�eG+��Gz���d��~����������������+ �J ��{5ׯ�j���],�{�~@����J�%�X����#ҳG��T'��_f�ذg�|A"J��������k��~>���K��}�S�)\Ӣ�N��k���n^e�ʬڻ��:��R�'εq�*������j�����3�!`T}qRZ~���|&�.ڒ'�#�d��D�@�Y�+l������A���J�S�}���Q����"�b̔� �$�����G��7�"@cؔpiYAR��v�q��R�3V:i���!���V�j�E�[��1�(-�T��،̹:[�X�{�j�d��S�F�~�VH��}������K��$IH&���O(��@}K�}��)��'���0	���z��1�h�3-;���,��:�j�/�ܾ��A�A|d�]�����N�n�b���a�YyA!�/�5y"A��% D��_��;u��Z;�����t_l���2nS��]U���}O�{����-�ԂsZ?lA|zu���HH��"H���sW_��r���@�U��
xzI�婌m�X?z����+��(�a�&�4�A���������o-�s!�y�=/a���d!�SZ���~�&�LH8F)� ��cEd����UJ��[�L���}�*��F�l��-	�ԤR����V���� @�a�SIi���R����;+��6a��#M��\�t(��FF�e���QEҴ���拶\+e�8�v��1��00j��r��ډ�������u�.�	Y�[+,J�m̯b(��K-��P���͵�ɭ���K/�fŤm���0;�T�L%e"˰���4+Z��c�c�++�������M��)RR��v�q<Sǜ�aЁ�����X3�MkZ(�����;��c���N}e�2��$�atx{�]p�-�|�)��+�-��0�Ylv,) A"J@�%� �A׻����گ=�۠�:�}o�@�9����x�Y�8�����yX ���$�~�q�>�9:�>��Z?�?I/�+H?%$�`�o�3�=���z��<'��`�z������"�I�����^�5�n=T��k����'����vK��%�����{����u�Ǘ��t4���^�H���/��4�_I�yٻ@�ɢǚ��z^�{��m�g^��c�פ�Ql̻�fh�uS4�Q�Ⱥ�7���2I��T�F�˚D;f�bL��h� �lJZɦtSZ��������!���+AJ_Z������ש���N�!�<6�d����v�����ܬD� ~� ~2E� (�])�*�j��2���l$����҅Y�x.�s51u�̴2��]+ڕ�F�����R�ZNǰj��.۩�������}.R�>���8�����E��GF���KN��^ w��b����\��i�c�#] D�B�~�J�H�D�sa1(�^��q`�p��/��-�C��"�}$B̔�������^�k�A68������ w�Hn���0�v��yKA�.���b�fd*���۪�=@�"@�$VA�~��i���=U��t�j�Y�t1q���\,���� �W�$)	V��lp���m�"�Uq4�X�b�5�c��V�Vʬ�\4��k�Yq P,fn�U�۽��ޠ� �� d��"Dy�ٳ�Rq���:��_�W�3U�e�3;e�ff�G2�C2�/�M>ø#t���!��|�!�z������r��l�m}�C���}A$D*�x�wS8��	��� LqY	@�"�$�=.�y4��}�w���gk�m�M�g��Y�r��:ȶ�q�YH�AI��3N�<s����A+�(3a��y��߁�
Hܞ|>U��w�d�o���Jl���Gz�\����r�K4M�ݬ���WýB��2 ���veη^td��5� �y}�t��Wtt{�`?^ �#����$�I,Y��U��e0��D�_e�Ǡ��.z�{�pgw�}�-�Qq���9�Y�rmQݭ�Uh��D$l�t��Ժj����J�Rg�A�ԍ�v�ãH&�t=�2�=�q��+���ń�8�[��)M��~��]]�/�=b갃�}�,�ԁ�+�"� �M����~��.�g��A��w�����xUѓ�|א �y}� ~��������|�Ù��CA�HHr�I,_�J_H����c�NN�����5��6Χdwh#�J��dA�A��ܟ��u��^����|~�X���v��cۗ=+#~ �7a|E?���NF�cr^ܠV�aڭ�[Z�~KMiS�UELE:��W�s��%S[ �uo����`�]�#��\���>��s��DO�S37��,F9�32�{���zWN4ƨ��:Mf��*`�2��� A���b��%����^[O~>g��40�+l]�`ԲѸ����0-ki��hGN�Z���E]z����\�˙�6����OA3�u=3r��m��}����}-P�~�A�/�D �"��Y5]yG�{^U9�(������ۑkl?i��+::=�M��^rř*��[�<�+���Dv���� �(#$VA�H��,���7=�Ǽ��&N=�?=�VA�L�|D����Y�u^�(Bnr�o�5�3n~n(�̄t^���nUzb�|�vAvxl1�	!����z�;�W�@�"@�"��/��Og�rS���v/�-c���"����*l��Gz�d�fJD���|sIx��\e�uy��o�5��oUN4o�6�9g����:X���xU-����3&;�m�K�=�ZT��V�Y������q�V�U���Mq�Ar��P�4LJ��K3`��[@n5)M�(Ǝر&s�7liUgZ�X�V��c�He�a����э�-�e@Rh�1ƴf�9���&,�0�Lm�l�le��U�mV4t`ZWLQ1�,mvL�aM�-ƅ�L�b٬
�;�V��V��W�e�%y  4�B�uĠʰ!��v*�3��k���V;L�pٝ���������Fh$Ÿ���ar��j�Q�)X�6�CF&���Rș�(�)	���H'n E�s1H ���:˭�9�%VL|{�~����=���޻s������q���Q̫��̫O���K�T5����;�r�	�=S�7.���o�}�A}A$C7f.]����8�G�o��� ~��K���5ױ�xR�e�%����m�ey;��f�eX�fU�fH��6*=荶�l�TwqIH�g���N~������'��df<�n����D�����$�A�X����dW�+�_�T�Dxh"�!�	<'��OK��F�徰A���$V2!t��mr%a�*�*6(!V�J�ҿ��	��/��a�b"j��&�nY�ڣ�V��g��/�ڲ�����hs㿽�%������3����w�-?9^"z!�̫��V&fkB�Qb�񶪪�a���ۯ{e���r�%�KF֠�K>��˕O����V�͹�7+F>�u�dݝ���i��}��pv=ko�|>��P8�Z�A�/��M��o:bP�9׳w�ď}�Ќ�Y`���޷y��]��n!t�=H���ř)"J�o��q�%�3�/8��jz]�5�-��z�@����X"J�A	���ͬ�no�0A�Z������,\���ֲUƻ��̍ �7c�YFf��u�v�s�t�X�OeL���̢ٙE�$RQ��:�X��-Ac�K�t��Vh�������{�Џ;e�fYs3,7��>�Y}�|@�6���I�����]�����k�J#i-�θCY�{�󥗬��������K��܋|_���E{n�}�|,B+���e{�h �΂>�V2 �� �H�#�ۙV��V�=��z������s���>\��)�^ w��%�2RW=�^m�x`$c������� �( �X&l��cH�w�3`̣�M��R��n�[�x�E�Nb*l;iײ�dC�i�]�|�YG��Շ}�q|.��޶����Vf@�G���|5x?�o6�P��p���	{�H6�G�_I����I��VR�T��J�A{��z�����o�����W���ݷ�w�/��6�Ǽo(a}�9~� A�/�D?IYV2M��y�n}v,v�g}��t������$w�~�,X2R��%{��\�KN�S�IW��E:��b��lb\	�������]f�ي���v:�� :Oz������OfT�ޭ�,d��hW�5�g�Yk�� ��!)H�� �&�z����� �G���ų{��"UY1����� ��2D�0|]N�|\�����?�Y����$�5w�U}���[p0���Y����7+�ޥ�\�`�HAR����	�ԟ����}A�~9��{��"��Ϗ��X���V������+&��f��.�N͹I=Ѻ��e���MA�����	����[��;�]�p�k�":�mѕtr��;��}�Ԕ3�%^���U\�t_� 5�32�{�Y�s*�S2�#������?O>"Т.�\c'�u�Zl���X ��_PFH��"�{�����/���ˆ��11�;m42Q^s1�ٕl�� ���LWn���Q2X�����/�>:Q=_	+�K��7�{����G NJ��}��ʏ����?k�u""JDI.���5ʩ�Mw��]�����H H��ħ�mм3�}[��{��?��
:�G��?G�N�D��@�F�_~�,_�J_$����g�2{oû���^���5�-C���/�%�}$Z2 ��$8��9J��Z���B���/��H��lӹ֌�C�>��24Ac��6�Բ{�޸*p��Ԉ�/���d���fj����G�����=�v�����4��Ё7T�m��ى}$C~�1b����К[�o�ٺ��q�Q�jIZ�Ǹ���f̃��caj�:�a�J���g���D�n����f���ق�����^[$��ù����ON�;>ǽ�X$=Υ�����:]P�v�k������9���N�p��������r�:*���܅#*���Pu,��8�s]Q�37&�X6�,��ktv�@�Q�×�O��*�R����M�5Up"/�w���w��N����,������ǀ�vy��T�"��`��m��bi�.�R�b�\��fL�l�y�X�-#AŜF�p���Z��p��.̳��PptO�u6�+P�y�5�Wfg*}D�{1�/y2΁����̹����#Cr���&qhZ����J���@�K���}�a�����ky�xJ��+w��V���Z���z�kB�w�%� >*��4r�^Ͳ)�ܭ�����%e!A���iu+$��+�*�KkL�=�ɳ���ܦ�U��)뭽�;>����e�}�t0U�T��[ �tJ�r�]û{[\��W�]RX:U��T��X���a�˂��a����-Ҳ.MX�}Y�T�.OQ���GgRܝVse}4Ǎiܼ���M��U)��O���T4YΪ���f ����,<	��e�k��%"c5�S��vWU��/JBn.��K�N�5��<;��<�f���v)��"�T�*)�E���30=}�n�:�ov�]�����UV(�Wx#̶2��H�wU�j�UC���R�C�����3��;4�4^0鍊�v���:֍xu��e2�P��W0�U����Ӈd)M5T,���)�JΊ������3��3Yqy��gY��gYqQŶ˿.��:-*;��!*��VM����޻<��ӽ�����e����⣻;:�[l��:8�lQq���m�����n��8��R<�&�YVwiVFw�Au���=$��^��էqW����ә�eݝ��@��^:H7���oJD����{]�U�ZgYtEae���y��:�ӻ�gg/��Gt��Ɨ{ۊ�*.ɶu���1(.���_k��
�����|���+涍���Zy��Ygn�̣;������(B%��Y�����15Ir�Y\��j�a�e���a��[��Y�,�`L��1v&���1V�8�ĸ���ٴԤ.�əd�R��E�l�`��R�f�!Q��.�:������2�hJ�[�n)M&��Yb��Q����\��S#Mq͵W�Mu���v�f��Tk�[�ۦJ颗�˥2�$.F���,�լ���bQ�U�(b�0�5��)jH:\�0�1��ͤ\�iY�M��)�0Ԅ�hƯi� �f��t�IX,����قU���/Q��[б��e���WQ֜�J�躴242�n	�̱,)-V:W%�-�@�Ã5�ԕ�1B�wYy\�D��bUM*��v��GY���^�-�0ʄ�n�.Ph�4u�tS�r���Ҭ���K��.�WUj�
R-�Mc*5�m.�$I�e�*6�X����Մ�nv�)Q.�B�,j\]!H�1n��Q�ehYFJZ���.e�_�Y}���D���K�a�֥��v�RZ�T��ל͆��n���<���Y���5�j)�hfW1!4��s����ae1KQ&1��jf�2ݴYx�Hb�z�4Ks����"�"J/e�F���X�+������ux�kMt6��p^�M�J��!��K����!�L���rl1��S�7h�+�h�e�+���d�.������,
��6��أ�˝@�L:�v��]ZJeٚ��`ƶ�f �L��M����2ѵA�cV�+,�[���p�[1Y���av�l:����vYZ��а�tJf�Z�慣�x��"������f���Q:���1�HhC(ɀ4#F��S(6�fb$\��.��
`�Vg&ݥBK�JX�ˍi�p�	���A̤�J�8���ZE��#�s��(T�eeufoP�JXl�E�����sK2��cq4CE�H�y.F����u�e:R�e��dm�f-��:֪�cXYZc3L� ����IGZK�V
\��9�uHB6�d�'	eqc�)^��^P��V�+s�6Q�Z�WSU3�L����]uv �V]���5�Z[h��j�lnŸ*��+��+,nZ�m���Eu�i�"p[��CF"k��km�Q�&%@pLړb��Iaȉ7V�Y�̵�u	��k��nTc5�3b���i�摫Lj�T(��a�X)o-Nr�f�s���_�fIra��1SM����r
�k`50`T�t�b�E�Ƴf�h?�d��e����hd�AIH{xc�{�/Hi6
���պ����s�~ ���jH f ��D�E`������F�y�?f����bǣ��x����{9+�:�A�d�+�#����*����.�3�"J�H���ZL��m��޴:�H��Âu�մ<g�������H��d���7��Mm�0�3�"N�|�#2t�^�8���+�[�,ޠ�t���t'��U�Aq��J���#���y箺F��W��K��;���ߥs�S��${Ԁ �����߈���P�˥�|���;Tl2
��mn.�cV�STn��f��#�:��oK���0��嘇� d��H���OC��ݕ���j��w���)-2Ȃ��2K�� �% ���_���5�xH/>���f��(F��H���A����b�Z��E�
��v�z��v�*J`�v��k�%���>}�tq���v�LU�緓[���W�R����Tf�񼹵}�{�ᙈ��d@�"_Ij�z�糑���^�NJ��G�K��IZA��)$�~�C����П�( g���"
�o	���+�g�Ԡh9��<DH���~t����I[�% "II]^9Sn�%��mX������]��j���/#�"��}�O;�4�="�K��D�j�"�#2�Q�xy��jB�CF�L
���!\b;2��SF֊�L��b���}�X32�Ǚ�5�3����7�\��
rW�M�޳�Z{�[������X�\���9H�%�`�(/��6����s���~��D��3�9���ÂL�|��y}o�G�1X�B�;�:���Z ґI,Y��@�+'�/he�/����Sj�K���º�Ĝ��Dp%h��F�؋�r�+�6�Ǌ�����N�Q#���rN�����l����Jc�)Y��  �}�'������]��B��v��f^�����{�x�s�j��VA�6� �=_ �H��~p�e�;��M1����@���O=�=��|q� ���_�	�� �(/���� ���{���7�%O>>�C0I��g� �yX �� ~�/��Ŀ��U�3ׄ�|-*��ժ�����^���f	s� �X���`�L�dMu���^�)�\��2W�%gp�'���|Jl��V�X�"���;8�mv<�����?H��( d��S��)ׁ� �~�G�q
-�=~,N�;LE�F�!� A�,X2W�_�ݹ��}��x�J��P��ҾP�$VD���W;���,5��v˜���G�	�� �/�G�+�$����?gj�h���,�����i�)|3�c��/�M�uo��~=������z�F�M�ũ_�;7I�P�v�݂�(F-{����G&Ӕ�R���CR;Av�v�5yn�x�]}b[�g&��J��fʔ�.�d�?| �������~��"�"�A���H���d�r������O�{�����bi���� �ޯ��b����$��ɫ��V(o�<�k���f�Z
]�%��8m�t���1Hl� �4����ߦ���FK-��2E`��+���*w@��o}Y�n�#��V�ۉ�F4�y/��ř)��+�;~����6��>�S�"ug��'����JzM�{}`�ޠ� ���,�YM�V�����A�j�|�+��(/��%��
��]5gn�-v:A��w��ҹ����V#33F�ʴ`�+�&ؕ�;Ou�(m|�ZA!�n�T�@��7���	����1D2��C�y?�w�Ӽ��%"�� �$�`�]���ߨa�}���oמ�����;�X'�A�J"���۞�L'�(��u��N��a��V�q�r���.��RW%9����C]�#6b���	J�ˡn��[������)�:������|�5� �"��(ZN+X�%��G1������!��daȐ)�/g۠r��cJ�f���i5���.�����U,m�P��bViK�j0�4�NK�S#�scXrduR�M�.�l��IR�Q]l3#cm- �K�)^�F��Ԅ�fal�7(u�;1�u\X`+�x�H$�u�l�B-��*F�V#�b�%�YavUd���i���lk�.�j{�����l��;*a�M[-H]1\E�t]`��,i�B��[��k�Y+T}���L�̲�33F���Ow�8z��-�x�B���^�nt�76��_R��D��K��2P���.��c���}�Y܂�A�Y��/se?�������@�����4�ǫ>��hs�,�V�fh�9�h�e0�z>o`Z��.4]�5��*B��9p��VA��Ψ�ol]�Z[O�-#v���Ҿ�!���샐�b�
r�H$n� �VDJ�mK��n��|Fd�( A�"��=Z]��
�1����f{�^���(x�VA|���H�\�ڽL���R�f�R�0��a��SV���+T�
\a�hԌt�FWK�v(����[���U�'{�4�T�3*�f�V����_���l�V��_��ǔ�2P6�A;�}�D�/��P_"��h���j7�`��1�'O�z[��w2uCh�zV�ٻ��2KDΡS�x����S��"�1^[��U�Y��ǽ�k7�۫��}$!]�}{�.3�{F�����'X���b/*7�!�|��D���Gk�� �q��\��&J�H��$Cm5A�]���u�ҏ|�������@�;e�̻���2����cM�t1$��eH����űa�^��4U�3���m�㉚�!�q��_h�A������H���$
u\h�������o����P���� �;Ծrř) A��*�-���8;��İ ��v;\D0��X륺��g[M�8F�j���Z:�]U޴���41稸������� �v:ewt��`�}�/!��E��z�~=�\g�����Lʛ��SG�������q��h5p��!��/]�w��O	��W��A�P҂2E^�R�2��)����G���yX �"�I�|d�+�t���<�!Pn��ؚu���B��ޣ'�rekw/�vȼ�w�]���40�t��L�-ٝ��j��3\�s��T)�eC!�}��}��a�`�y�����R �rř)H���o�<*cܽ���T!쯷�i�@^���&�F��
v���	y�H�q�!�y]����c7�.s�f��W��R�fH�s!��`���#v{썆��w��vp_���_��A�A"�A�U|��|���|޾�ci��FZc��*���Ǖ�PNͺ�m���	�k��ɄVk�>��_?{o��_	0/�������7<}C;��
yQ�kq�wpL� �2�D���fG�"H��%��Uy�����4����L��WM�^.�Ϩ��7�}���V/��G�ɭ?>�?��{�,z� ��ř)|A�%?p{K�3��a�:OѰ�����6'�~�Z>�@9��#$VD��Cr���O�\�� �_�A|d�/ӟ3�����O8�h#v>�Z�(F=�y�*f�ȟ�;�5���D4�`�y�ֱ��㻄V��qXT:;R`�;����cWuRZ�����}9�/M�}W�RgZZ
�fK��u�t?��I~�����q��bff�L�2W�E3K/��?�$ҧ~����^�%��s�^_t�/�G���,_�/�����<�l]�T+Í�*�YvQ�f[.e��p��XK.��"#|�ߒ'ת �=b�2R �%/�=ڮ�r~�oQb�_���ë�ޝ�ݠ��/�~_\� ~�	�+U�otWK�Џ��_��M�nˌڍ��j�����#v>A�b����`���qv=cYH��/�� �+�"�~����޾����b��
2��9�/|������ ��%��IIZg���T�0�"�q��%i%cܪ�?/E��X��r�L�Z1ݚ�<{��G��G�?���A�/���H���#�f�{Ѫ���̱}<��E��-��M����"r������aQqS���+�-��+sS3ugrl&��bĶw�q���c�t�nǺ�SC��!��m����oXw]�ʨv0�N��<2�2��g  �;����~S�0f�[��J��H�[e�����&���k%�.��p�/�s����־Q�v�[`������=i�Z���/Q&��W�&k�5�W��xi�MR���#er�!s	�Xݘ��ٹ����j�Hh�
�R���g�;�	����L�`6Tneb4Y�IZ-��[kTWe͛J��F[RcfU���[��uq���?|�?���L�FV�Skv�N4�Y����c�pʶ�L�.7aK�X �@/���2EdA��sw:���b�������	�&	$��}\��^~�#1�<��2����D:z����4'�h�)�������I����V�I�D$�爛�����u�|��NO8�����q	($BH�h�����6�����k�Ww:���:y
�]�}�{��~�%I� $�Ѷ=x߻�m�W��z��j���� ����}$@He׾]b.�ī���K�M���/ZʃYi�5�l�:l� 3�A5t0��[����V+j��C����}$A�l��WxM���{���Af_��2�V������I�/����Vebv���~��q��V��i^�)z]�7��l\�=�7dS7�=���XgeK[˅·��ģ�3[Q���ۅؒ����#޻T?�}I~�_}ޠm~�S��^�1{��/�I2�f�+<��_>�BJ�I��Z���w*�?
��mSE�w����!��	$���VnrN���:E$Nv�8��anr�7[��UD'끋cm����3�(}C�&T�5-�~�S��Ⱥa��)���r��}��>�`�I��l���I��o�|u�:\n
�B��jP�����9�%[]�)X4E�EZ�J�V��gE)+�$C4W����ʋF�O��~��5'o>��ݯ����Ib�]�s�W>΋�: �l�����{�o��w���I�^7�Z��Y�K�5}�BI$�$���Y=�S!�;\��ÛĐ����d���a����sv�������
��Gf�E �U,�n�HvZ��s�z��j+�y�]�]\ʅT�_tݡ�i�*��B��Z,U�͊¹j�K�`�A�"����(��v�k�}uGE��ffL��>I��sK�6���>��-�]/�3c��%*��%6�r�I�����U�u(Y|2[h\�uSkm�L̎έ�"���{Jrk5��]�꒨��S2�:���_>�*�n���:�G��,UQ�<Z�̿]�A�[�n�e�M���fѾ{�]ݚ�`��Ҫ�l.#\�ux��Շ��Z9��5iB��L�,���Xl*��2�����l�[�GX�к�F\�2�(()V�DC.� wbÍ�+n�slؾK�>z^m�]�
�4���u���:ʇx��9{�	(�$�i�.�ٚ9�]�+7�F*��̕��@�&%�����[(挏p@���iלhY���a�J3�i1o��zI�λ��f.�2��T��uy��|
uN;���Q����U�[T�dҲ���������,�����Q�y}P]��V�{�*��{�:�<�=f�
w���	���j����Ļk��g%����S�݋�I��^f���2-�9�2W�{1�eu+UGx�RJy�C.
��ٽ����b�/J������7j<��ui<��sEΛ�j�9.iwOճ��m>��n���k�(�z�K	�m�4��ͭU�b���u�L�+ZJ��o-�Ѓ�	�)�V�y�̓�[3�X�R�n��~mgFg���7����m)-���i-Lf�7D*��M��;���$�ǭ�Oj��[���gq|��mYYo�n����1����|=�Vf]�xW�y����6�O��	�Yw�ٟ<J��#,�
R�e�u�F��]@ˠ�XI�]�&8:bb�!ɉ-� �h��ޢt�I)IH[ؗ�����$�,�RɶI���_m|�h���q�%����󬳼��M����/�EF���ŶD帓�)�g$��I%9$��R"F��@�wov��|����{gYv%��(���B�kF�Jk�� �d�?����ړ%{��E�-\�ý��$_I�iT0���>����I��;�+��i��Y���`�h�d�w�T�|$��(I/rX�k���蟓� +�ruK����� $�I@IR�j�n�2"br�.�m�)1�E�H�Y��X�!�uF+�(٨A����$R�3�l����@���o�Wt�S��ڎj�(�<}S+��Y�Γ �!%|$��x��{/;v���3E�����ZT�Y�����)!����n�_��nl�LI�/�G��$���{�Y:���o�{�AȤ�$RM�+{�����U��G���I�[缤�Sܱ���;�_;gA��Y)\Sَ����v��RUq�V�-JJ���PW��r̝3����%3T���e�ͮ����OҫN���AE5U}����e���3#�"H��	Y��Ha��Þ�'��]*zWz{{�	"�I۶�3��b���҅5����]�����&��]�!Yq��
�L����eL(������ըvFf!���c`��c�߁��K�������vI�E��|$��V�#E���ކx��s�J4��yt�Sܱ�����T�2���o��7�W�g��	"W�I=���;�O&3�ttd��J�����z��)"JD�^ߢ��w��7(>� I����9�U���=� 3��|G���Ƕ���H�P�I":�{_J�lKa���t�Tܱ����_(I��w(C^㕞����v�#b9��Z�k=N�﷠̻�I�뱵���k��طhv%E�4��%/Y[X���~L~|;��B���.�6�\�KՃK�"�.,��7W0�A��׬lԡS66����7*���Äep5���������a6�/[ &�E8�f.�WG1��V%�l��LY	�J�R,:�Nof�:��K cem�Z@��ym˥v��q�1 ��-��v���a�l��X�8����!Z��s���7du�es�tVct����h�������Ycf�U���z�,c,�Z�E7T�R�$��?]R�`���us�	�I3F����������z%ԫŸ�>��Z�J�/��s��Ut��xhM��z��:WVd�r>��� �c��#:�ȅ�WL�3bW�E$@I���6�����ut~��cj9O�{�_$�$�IS�]y\�.��_OW�Iٺn�����ixq�s���w+��=��tC��$_	"�I!�J�ʠ;9V���=^��*�|~����IRE_xL{��T�W`�бR��.�$��r�mcwX0f
�]
B�meaK����}W�t�@��n�ή�Փ,mG)���y^�J���H��L�]��2�r�~���4fy�T]GI�F'�k�	N�eR�=l��q��G풷�y빙y���Z���\�R��Y��/ݤa�׽�}��f�mG��z��mg"������}=_����͜�'׫Z�NBJD$���6�E������\�	o�{���!%��	"N��o�}o���*�ѳ����Y34�r������
B{s9}��g�H��I���R���������o���u��M32�#��'������* �(�sa�t#�b��ڵJ���U�����v�k�Є&`ɋWBeХ�.%�e����}=RE$3���x�nGWB[�ܞ�����=�\��+�$�D����,c"�z�z����Ѿ����Y34��~���r��^V��_�%��٪u|;ܾ�/��$��hYߝr����-�����9w4�Q�Cl�}(�+��5t�1�~�7+$&:�
����r�q��.���X<�˪���(Y�F�}���7:�Y��i���9߾���RE$�����i�Au�W�3ю�e��^ˉ�xMށ�P>�k��v/h�nV>��{��!�����$�Փ��*Q�P���������Y/6�q߇����L�H��ۿz:�"�Ҡ���a4*�t3
�.n�h`[���V]��A�%A��I�c��l����f�Vu���wSH�x:��xU���7�BJE��f8�Z��N�6u ��ݶ������-���y|$�I�ԑѣdSW�E$_I��B��ʦ1��d�Q8����I3�$��|V=��JE���s���pk<o��ћ:N�l=(��W�U��gU���bS<_vt[F�<%c��m1�'����W����;5m�%v��n�s;U�4:7\�ެ0N7!�,�p��־���f/��$�?:a���=���ַJt�[��y �_IBHg��fZ%U��W�l6�� �2����;$�q�C)U�sSk�4�U���G����H����uݓ}o^�E�?���z�`��P�W�yI���+n��������^�Q�N3F��`���z3cg/��X`�r^���l�6I2H��E�nn�޵n��{S�]��{���E%|$�I.�N�KD��Wϻ~���[O�[�Ӛ��dއ��kbvܚa��{k����{���$�H����}Waq�1z�����p��{W]�=_l��Ho.�),��f��t^�nU
�_JT7.�����W��ga͠�}Î�sCdb:���I��z^�M��mf>�V������| ��E$��`�.u(u%ٳ7Mc��TT�,ָٙlV[)Hh����&�8�貯��	��C/d.D��P�t�%�]�I��ġ�UQ�e&���ѥGC�U��lWG��i�`4���.������=IL],L�M�`��ɐ`@�^�_<��H� nN&(�'1�옋���-�n�U�I]�4�P�XR#�-X)��m�� Q�߿�������S�P�V����{�<�mcu��1a0�P���]5�8�|*�}�fb��u�[�m���m�<���O{�G��;�}$�>�![
���eW�����J��o>]�����SJ�kF����8VBcw>�Kᾯ����	(Io=e�[s*W���`oh�xOP��MI%o�X�{�G�G�q��ᙛ�e�+i�L7��F�C���G���g������y	"�JI"0��f»�n"o7u?:�I�9S�Z��I2I��^�&���)�?Z_U*���.����uCBR��1Dͮ:��L\�^ڿ��~ސ���IBH�V�W�w���0=�9ʝ �}����%�Nߤ�$BH��t~���[V���a���C��Ws���0�;��+HJ�Rݜ��.�ȉ��ս,r�`�r�<z��Ы���}���CS�����ךyPn�=�ffd�[��<}�;���MK���"�H9�r��9{=����s7���r��	"P~��96��f|7��	"�[Y[��Bo�ѡ��8�)#����ymb�ޡ$_I�T�����X�kV6'p������h��{�	$�$��7���w�zl��3��:,]K3	Kn�(���`̭�LZ�HhA�6�k��|��$��(U�􋳷�:��yw7}���5�m�n�l��H������>>�J>Y[�#�xz���N��	�g)&�2��k�e)=�^�褒`C�}s�'�N�4Q�׃���ZG6��ɢ9G�nwm���	��OB����,������(��Dg�o5݂�-�:�/f��={�f�T�qwmw��v	�=5-<�9}���}������]{z
k�u}��О�$����?:����NV�����R*\|}^ŀ[��JE��D5�L�^��E6����՝�`�tg{���>RE�^+p�7��zOa�5Uf�7v��I\/mlTn)�Wqv�ie��tY�f��J�S���A$^Y�{�]g�v�t�1ѳ�[��^W~�tF�W�E$@H��7�m�������E���ܜ�������rHNo��Ƹ���u�_I$���u�>��r�+�&v�=�%ugu�&��z��� $�"�ڸ:���U��S�?s���Ū��lL{tԴ���ٺ��孹2����p�4�:Z���<p��bU'V.*��Y��J�n�d�����z���PCo��t���8�\�p��j�5��{
���{}�3�"���/��]z^^]��.��s~�ݹ���������I�HGi<�����,g媦��\d(Uf�@qnV���5���]��#V�$lS�;}��%}���ݕ{�i�,`�z�|�Q2����ݬȒ/����1�H�s��:���V�W>���m_W=���I&[�Y�޷�>d<�7ӽ�}$@I�{�{4��Y���K�m��{k&��{���>�Iۏ��d�����;��ݎ���;ˇ�;�z��k=��c/��BI&	"�IRM��c��ٙ�t�����wj�u/F{��$BJI�|k9�u]��:�`b�v(oLi���v��Y��
��^�����-3;a�F�R׍۱bĎ<%��}y�wO��\�Jl6^Zv��3ԣ�e<|���]X<�O�����(N'�4��W�/��V�!p�*�'6v�匳Z�"�SZ�����Q6+��]#VQDme�����l�2��[G���ܘ9�����9e�rf�&e�Ў�T��4`��Tr��6������^�N�Z�RL�U�����]����hч&�2r���U9�[#�l��QΗ��@�Ppǖ�,�5u�sw�v����[�w`Ǉ�s6�7Eu<�>�k9�[c+/.�6��e.y���ӴV��U�}�fv�̸��:��|��[p5�Z{j�O���;O�ܡ����,;hh1gfUw��㐓����qv������ki��8cT�<6�4�s��q����cڿ��q{��̓��W��C����A�Uͬ9ϱowf��7H����D��fa����u�y��f|�c;/7M���(��9l��,]�NAs��SIk��Y�e���q�B/ܷT�v���TifYݾ��n�NYs3�gb�Tv�YSU�Y�z�����MaWD�{cmc��N��i΍
��ro��ə��M�Ӭ�xiU��[:�E��8;�V(Ke�baR%��J���Mc�yW}�{w�^깐*�β��G��R��C�m�~�e�Л�Y��Xy��;��+��t�vP��������)N,(N!>k���H��R[C��:�@�D�Y.���-�R4���5�/T�׶Օ�F�#zZ�q����Xn�4)-��5�XXSh@�k�ŲLH�lm����{��PB�+z�#&z����bt۱�VEo�z�/��/-�nQ|�=�u��΋0���ݧw�{u�x�Үl��X�d]���RF���g�|��Χ�y�V\G�Qy�]�Xq�x�m޽��mhqu����f<����|�-�U�-�̬+[,	�idl����gGW�Z�>|�8^j��ͷ¼�{d����+��]��8 Mv��)���F���y�&гY��R�,�ם)���[`wf�� �΀��C[*uK=w�Q{;axܦ��h��l
�`e�aQ��*��
8�����Tc[��&�`Y .m��GR��!��ͤ�e���-l%1,cJ��a�D��m�v5m�1,���ډ3�ѱ���UyѷR�L.�/R�ٲE!��[�l�\Jl�`�5Z�J�iM�����2�Xsj��K��C-4���-J5O�r����ČI�Ѱcc����e�j��#U�I\�acX�D���p��1`���!���gv�lbS,[B�W]) D#�S�l�nmVG��{"�ڳXԫt�\�sE�ڵ#Dv+��*�+rs-�)1s�l��Y��L���).��h�k0��K�[5��fUToTq*Y�F��U�19��R"��K����6����%����8MtrR�#���g4�M����5v���X�5̓�`��&����W+2��\��X%���GY��SSb�ܚ�F��+s��JC0D��Ŵ4uR�#�lҔ�v��e�x���]KymQv��vrcE�\��=k�qm�+�3Z�9j��r��K�V��u�Q�����V��i��dΣyj�Yec4P4�2��Mv%*3Es[4Z��W���4�����5��	�а���lkK#ՎIl�L��[e�4��e�.�r���:�IZ����	rͬ.�w]��]�{E6Ύ*+����n��r[�j�6*�4����v#x�1i��,`S:5���k��f�������
���jJ�y�Z:��q5��aD,��qX[��h�bU����+

��WD.e�D�z�����-��&t�)��ԥ�6CR�L9��D
���GVJ���k�4e�!���R�t8�%E�(FnVCM��m�V��2!n�`ƥ#]�7�µ�����u���,%�RLh��B����]�섵;U�*m�%[YH4�S@ج�E���i��1�h�&�+0c2�m���&��릦쭬���a�����lh5�����b�1f:�8xFP`�C�MT2��;f9�$�)����#
@bZ��l� �mjQn!�H�ռ��2M�v��kBd!`�����LA�qQ�S�mΩ�9��z��u��ֶ�J@!��U���D��Aؼ6��c����5+6	l��Ís���P[��C	�pYH�bbŦ|L�L����
�5p�mj��]�1�����a�-P��5e�K̯Tu5�Q�j9�f=��}im��#�v���ih�R.4%�Bg*ـ���g"���������脑}!�q���J��ݭ�{=�vHC�����|��I$τ����94�#<o�[�|��Ez���wM4�U�}:�����u'�j��o��	*H��&�9~����0���|��~�yI���I��By��Y�ؾ��2�jwmzC�Nӛ�{�A6/$%��sWH��$��$���ieo<����/�;˸��'�ӫ�9I$�
��a���ߟ���ǋrq2� hE�3����&O6i��4�fT9H�K���Hĩ�� �#���Uۙ����Mz���~���c��9T���A���$�"P����fe�D����E��]I�^��
"i��)^M�%:��}i�J�2��vHs\���.�����2��y�wr�0� O,��5y�~��	�x�S��k�-9����ʒ/#��$
o��=�M�I_	#�2�>��-)sV�sn���c�={�3�D�$B�7�9X��!��yf�q�Xݨf]������g����s>��t�hP�!$46���e�:�y����8&�ꖤ�}�y|�	"�^_�|S���������[�Fͺ�bU�*���l`���$�j�Pҭ�Y����6m_�$��2~�����"�5f����Y�LF?�B3jc��>�F�N_I$Ϥ�Rշ�\��r����e�	cv��wPr��Vf!��^cWr}��z7��$RD$}�%^��F����+뗼f�6�\ɊPg����������"{{V0�nrS����w��nf�X�٫�6��ir���<�{�9�����������ˇ�S�����rI�I���Ge�W�7vcz2E��"�<�O[���`Z5��ԙ�n��W�мw��ٝ��_I�/��$g<�X�+���i�=Rχ���]�F?� $�I@I3Ng |iݽ��￴�:�6����#�-�5��Yk2F]�[+������VQ�`M����/�����/÷���.n��T����V:�/�$�H����V�n�y�-��e�Vx?{�����`Z5�N���$�{Z�@� n��m�3��z�
�%�����ymg���޵�4G����LI#k���G];Z���jo�&�fO{��ڋ�1y�b��פ�Y~%���a��e�Gp�&��2��S�W/�7���+)+鴸�4��V�uc{��m|r�߂�_|�RW�E$RV�}\ޒ�|����u:���&�_��A�I4}'��T]�4a^eTW�顗uk�0�6e�����Zh��v�-q5u�A�7vhҫ�繯��I�I=M�s��3E9^b�ހ��1
nZԣ��W�D$��0��6�Oeɜ�s_t�Y1���ݙ0N�2{��y|�$����J{�3���KBz���������o����p��}�QZ5������D�$B���D&�i��lt�I�o��(z)��.��ւ5	Q��197 ^ӑ|$�JI�\�=��z	A�W=��[���ɂv���{�C�*H�O���]z��ޚ(�g���&�x��YF�*j�����HrjѪ�nm2�����Ug�FP�{^�[�2{m�z;���~z��ۉ_�9r�j�1���L�лi����ְ���fS:�8Bj+�B�K�ם�f僳��v���bM������ML�9�İ�Љk�%`�2ز�K��Xۄ�5�-n�+����W�G\���`�J�-�R&��+u�#���1����4���E��
Z�t%�X���[)6u�MQ�Ƌ�;`V�,�l�@�-�25�s���ϕD�B�)i�(��e��0�#u�Ebma�L�;&�Фh�"�C���ϟ^���%}$�^�T|<9�Eh�N�(���o�܃}&	"I�S#$�������E�&���Y^�ε�47�	"������ɋ�i+V��J�&��0i���l������^��b��;���y|�}$@IM��w�*e����H�W����^7q�U�������{^��h�6�=�"D$�$�7�D���圵H�{�u�᡿zy|$�`M�O�/�׮��=�F��XoQ�Ûku�C��ƀFmc�*R�X��K0�mv�V�__O�{�w߿�	(
������=&	�d�|v�V�����h�o�����I$Ϥ���x�/\����,���=3ɽh�����\we�aY�N��fN�L�v��z�0�]sa��\���p�N�!O�]U",�N�>�f���l�ʇ���DB�Y��^431��y;�[1�gT}y�z�J�)"��I�����v��ה�:�^���[�C~��	"W�D$����������d�߀����������2`�fM���d�~k᳔��I�yn�ݬ�J*����v��!��۸�R+7�qs�� ��:=���^F|5P�J��h)6���ޤ��O���l3S���،5q5c�����W!{3٘�����O˶a�S�]���������}@I�}%}l'bڣYx>��C��w-���R�}fM�����POX3&�+ �ޗ�|�@I$Ϥ� ,�{��+4�IZl�|�Ooks���Ψ렑��{C�u�8`\q�+����ò��gR�$Ȑ��0�R깘�Ȭ��3����Ϊ���u9	$�u .���s
�}��'��E��3;=~����}ފ��Xi����-�{>�$BJ�H�e����ܾ>���[���JD������JE��{L��+��Vn�*����p9���m�'�l��MŽ�afd"������߿&	"�����~њ�xg��{�V����_
�����8��$�Iﾭy�
�5�sٹ4'��ԧ� wD�}$��{��9�ްK��]��I$��u?U�X��g��r{6�Io�ܞ�y}%}$@I�8�ܵ���8t.���_t�$�5����΍嘅>9��)�;��n�_����lG}yW���B��X�Q7|3n��t�e�=�F���V,����w��'��*��K3G�,�I.K^����$@I�T�R��WU�ޮ�TV����)۞����;�9���n.�|�O>~����P��� �K�Ys�[b6h�`���b$m�)-�A��'W[�j��}�~=�����Jzouv_z��9}2��o`u��r}V��t�I@I�%(���׫�����,������Fj���|;�9	 !T^�7ʫ_��{�	$�$�d̏n/[SGM��z��\0G��|�JD�}X�3Na�[%�ӑ	(R��[���D,�y��f���y������a��H�~�JD$��7#Aʚ�-�~�{�;���ﻨ|�$R	7}�tn���$�V˛��B;m�!���P]V�l�mض"(�(9>����J"�i�QE�Æ���uYB��	k]7�-�h*V*�QWܛX95��&5ؽ[�J���
�y��o.��ٱ��J��U�7j]v�6��K��.rV�6�b�[�֒�K���X2�g����e��*�\Зu�+��8�����,�IX�f�����u����34�͙zfX����6�`qJ�1���	a-��/Ynfe#(�]�pՆS.
;k1��9�B�a(�G
�s�}�����h���éf���]*�MqYF�2�q2�㶉k�x��[H���v��٘�1m];g�kkc���?K5������73�ͯ��_I�E��S�N���v��u
^��;/�3
�:e\��y+�%S�t�Zoծ!��~�	"���f��X6�L��z�?u����3���n�� ;��'!$RT�۞<]_G~�u���H�7��gL��x�LP�߷mK�W���k�y��k3���I��:�]�G7ў�\��)�}�$�����`�ILi��?N9l��%mh�@>��hѮ� A�,4ԗM��`.�� ��pi���%J��*
�u�G�#�0	"����q����b����N�g����w/�����"L��W��e��FL��0^��ҽ��D����W�h��Wmk�,��T��9>�M3�.�l�>X��;�r�g�<�k[Xz��uGyw���/=��g+�C���O}���>�9u�ߴ���n���u ;���	"�߼��ʣ�������T�����{�$�$�IuA̍]��^��S�I��y�����T���;�n��Y��⽟nj��$@I���ގ�^Ox��A�W����3˳��>\��{|�}��}~�~��ޟ>G���O��v�df��Il��yɣ"J�ѸD��L44{P�����Sk����|$������J����u�xf&>�r{�5�<�D=Ѥ�}���"�IIV
��ոxv�oϢW������T���:����oV{؍���I�=��*H��I����So�]�䔚4sY�]�Z$�[A�iܩ/�2�i�*0��5����GU<�MbW}W�̻���d�t�VVf�To>=1�CMC$"�BU+�[N�K�*�! �:����k/g��]�i\bm��X\4Mʺ����ɡYG�oP:�}�,����~�,ݐ޹�-��ܕ�*�oi�*�]L�9�a�U�!y�,XP�E�sw�&�0��b��ӢC2�V
]r��J��Gj��r�]&��R�-7����aU豎�SNW^Y".���q��5�5�M�x��L���9æ�cy��Kv�ו_jz��ڗ���z�gmUe�߸�;s1<�6[Тֈ���=g�Yܡ�E� <VT���9��o�WK���;��Y��\9�yJ�ܫ�uV���`�����le]������J��r���sn(�Z���1�܆K��Sw/�}�Gh؃��R�}�~#)�.�1�^��H�I�oRλe��w�g蒛X����N�2:�J��ͻ�M�Ie�~�t0�ʨp1�䓉�X�>.��\����UG���'n��V����5*�ݳ�LU@��Gb$����i}�NR2X]R9Cf��צ�2^V�zrN��	r��"������*Si.��5�V�|�ڕ}�ܥT��ga�̗.Վ�%�Z�q}���-�7�>%N���9sl@�$�Y}�h�n�i�d�ȁxs�w��x)�N�]-7w"P:8�*�_�G++��+�,���K;o/B�Ōi2��5n��_��g����a?*(q
P�,�����f���γH���n��}��=�"���_z���Yd5$m�'LS����m�9�|�8�{{�D�$P�K��<�ô��6ܑN6���b����G!��v��|�u�I=�9'$%�n����,�/kp��^^9�Y�ye�m�.�ԛ۽à����Zv��0�N(�o��u��<��'�^��-,�F����Y��2D8�^ץ�u��g���Ol��h��o��u�g���<��;m�J��<{n�hW��>��:N�e�n���X��{���bA���Y�H����K,��(u��!v:)R7���hvKu1l�@�XYj� �&�/m`	I�Jq5t-��E���J���n��Z�jK-�$���S���C����$;��[cgXJ��I�E[�}�)�pN�_$��@>��E$_a��l1����4>OqIF_���}�S�����_`���ޚ�G�����!%	"D$�s0_	���}7s9V�z��ޣ2xRb�xN�')"q���y
�.���РMV�o��Cv���f���me�ن.Ś��0�A���{|��Ir.v���]���k�0�W
�5r�2z�������I �1X��{��n���	���u���'3{���'(I=����8�܊/0#��H��$��;�ʺr��Q~�(̝E1hgx|;��'/��I$�ĉy��v_fP��$C��|s�W��}���y��Ð��y��K	�+�m���hm,���P=	�'q)��p��.�Ń�l���֘�qKღ��kIx�.�:�	�OB���W�dBH��$�H5�����|=�T�^������W��&f��5ƻ��T�ۺީ�]VT��k������U-�G�&B�ؖ ������yq{ܾ���%��
noB�z�1hl��֞n��^���1�sP�y%9�D����1�:���{.7�+��k������w��"��=�XL{�^m����M�I��K{;l94;�s��W��w��7���P��}%Ig6v�֧PE�Y��u��VOQ�-�ʂ��;n�G8�$�I���� �=������J�~����~�ht�JI��z�S�����y�5N��o�(�'/ElEٿ_/L{���^�x8G�(<ؒ�/TB��^
�_gk�lD�ܐ"���}��b}�m��B|++un��f�,4s�����1P�`�Sk�������l@)`��Sa�ޡC=D������]�m	��ZjcYJ��B؎�FT��Q�5�ܕJ)�qm�7$s	k]��tqo0V��଻ki�D*�C(�e��˵��r��h��i��u([�(k�a��b$к�a�\e��
�c5rEq�1�7e�+�a�e|��_�ߺ�95�K��5�e�-¤Y�6ց�\e���(�������|�t�_I��Y5��]�e��޳rx� ��W��V�ݠ'r�I&}$_m��P���==sM���P�������\�8š��������q�6�m}]�K�p��/����	 ��N�}�o����볃�y�="���E��|n��.N��g!�wc݈y���˚��]���`޳rww�+՜�r��3Ⱦ�	+�$@I�+֝��}�)9��k�̞G�6{��BN@I�l���7�̻�nՂ���n�nA��G\:\�],�i^ �d,f�l�K0�5F�X������z��H��͇���Y���~ڬ�
���æɟ	"�/�׆%��2ޕ]��=7�y.���{�Y���ӱ�:���3k�o_�Q9�e�ۺy;��[T�W��u��L=l*Bo�O��|=J5������y�еls9"���5��w)#�m��<!�Q����8��H�P��-�n �ۑ���}pg����3��o��ej>������� ��Cng�A�RC���5�!���U�����	m��q����=�˖,py�}��H�������&�I^���$��A�rn���mȐCnI9%�j�>?*BU[|����H�'}�}��R� [k�����[J�<od#0 ��"~�i�I�轭�p
h�.6f��A�����҃Ze#��=��	�В��$���mș��'���u���.���Cp8�����;ؠAܹ뿧�_6�	m���N�����ߖyq���W�G���.X��s��|��G6��[���:�{Qo�y��(�wL�l|�nD�ۑ?C�rV���(�P�Y�p��D�Q���
���W�̢)��7s�ڋ����O��U�DM�n�;��Ft�ջpbF�&�u��@��eӴ�8l\�r{���w) �k�ڣ�mO�6�jkm�O������B��k��nD�VqmK�]������{�pt�T���&(��'�܂-���S��E��{�N����kU�ʼ<<�a�Ŏ��=|����H-� ��U�Ŕ==��b`(~���Vٻf4��p�"����&��I����[rLJ�Q&N���A:�m�۱?���f��c���������]�FҍLٱ����nV~�A��H%����@��E'8���z�F{���_u􅵜�&r�es������ �_B ��Cn7�w�T��瑑�*���}F��Ch"�R ���S9�Ւ�f���p<6�X���|_ '����6П�m̂���>��J>��4����hz)�t�N:���NN���o)���w����k"�}QR%Υf�k0���}���7{�\is���36��`�N�����rP�����Vs�nf�����z�P`�*��������a��~� ���!�%���m���<�ǌm(bݠ��_t??^�E��b+�^��_Cݑ ���Ŵ)��lF�4��gLF�	Kao�n�Y� V�:84L�mا:m���D�
�4��~[�#?Gʹmm���=����X����Ϸ,��qܾn>�܉6�A����ǆ}>����{"~:�_R��V���brE9=���K�RAm|�W}��i���.1���+��@�u�Cm	-��ș�3סG�����{�i����{��� F� �_7�m���%�qI�n�E�@6Ս��֣�農̱C��}��;�+K��;�b�� ���$ۙ��D�nD��{5%�w����=��(.ɻ�/N�S�)��]���n-�$�m7����
���O����xE�;ShҺ�A�p+z�O�u4ľ�s����t�p�*�Y��y����:�0��IT)c`ͭ�F὚�T��Y��)`EYz�R[!f���--K*����#�VP�v��G��1ma[v�Q�#Q�8�tB%J�+�s)2�au�B-�j.M���E���m�$$^b�va\0Фh�-L�[�ͺ�&ڨ� iv��hV��c+{XGQ�RӴ��;R�"L�"[�6�Ȩ��a��0�*��T����?O٭��. Q��a� Զ	(�.�����w1z�XX��XQ
%½�/��	!��%��6�H�z���^���0��+�V�g�{�����9�s"��$[����m� �ڒ7n�{������z��{fxx�4ƺ��qD{��1CE� ����������̋&ǆ�H�bA�������Й��³ڑ�j�:Q��2�ly�8�9=�����A��-�?Am� ��!>��^u�1^��'�k�%� A܉�^��U���r��U�)�}v�gn?��ف���]"~{ڐA�������R�FW�BA��#5�樏=�ܦ(p���s��#9Ȑ[�-��bQ�TP?r!DAE&cƋۋ�h-�X�l6ԤԸ�)q*�W��5~E��A5Ё� 6�~nR���'�'�����n�q4�Q�8��A�@��$�_7K����1�۷�yf��#W���t�nN��c���t��4�k����u$s�saw]��f�Ε���2'���>θ2�ۯ�|s#干���Uz�:ܯK
�E>	}��ȐCo��~���U[�c��_P;�I�����m��M�W� �]l�Q��z-�b���! y�[�A��r2��L}tˍ ����@��hz��2��ab��W	��?9�ϝFфƃ�j~ �Ƥ���6�In;&�w�ȯ1*}"~�������s�^L*��p/�������·�������Q
T��0�D��sWE05Ŗ0�lM��\�LM��LB`fC齺A����~�_6�	m��ݶ�y��1C�� ����N�5�X��x�-� �,	4 A��=cd���n�9_��+r@��h/�Oن^���a�Oǽ���o)��A�sGO����tT��h�RGR@�o�	܉-��7!w���T�#>��9v".n���U ��c��t"#��z�^�l\��j�U�ṣ|ҍߪY�XqMǦRL47N��_>�l��Z��[���^nz�y��&p����D�d݉���_�S�!���!��}����� �m����iG���nS8^����!$W=�5dY�G�n}����$6�H%�D܉!�1�lq�w��\��I��]�#z��"��ej�~�� �_6�Km[�����?B	��e�j��*��iH�����m�)��L(��jQ"4E���В-�p�m�"}{�߫׹q|=*��#�u�ҋ����;F�BA�"~?6�m��ڐFG]���/�JA��S����t�
r���s�'���7"Kq7�م�'���f���� ��݉���W{½��"�����h�چ�~=����{yH �_6���!��p܆���ː� ۹�9Ё�܉���o���7|=*��${a3�4����~�i8���S����,��Z�0;��NN�w�Uݕ�;lU;�f�V�(�^��)E[p.8��	�o;4�
�ں�����|{lO��8ڟ�%����_��P�=R3�~1��=�x��n���)�p@�o�#��%��|ۑ���g�����[�@���	l^&V�c��p�5d)��4I���72ڰjUm���?~o�?.!'�l�!�����fQ�����"�������<��f`����r�A-�$6��W��Db�����G��$*��o��ї|=/p��Ƕ�ȐCo�)x���5�uh guO��z�[A�R%��uNz;�}��+S2�u��9}}�H �r$� �X���;��d�H�g�{ڀ���@���ՙOVҝ��4��V� ��REq�z�n⧧����R?�S���m�$���+LV�Hn�B�m/==2$&������/��^����/�^�۱?����M�x��;8�l_wy�#.��k��[�����tw�`uV0�v�9�L�zދ��$�:�j�Tzơ�������Ț��f�ְ�ڧV���#�vn[[7��ׯ����X��j��0>*�Y�.E�A�>�{���׋0:�F��7ee;Y!J����
}׊����ch��V���m۫Ǆ����|/�m]nQ}uY��Y
��N�.�T\6�v��V�k+�1t;�u&j����%���mww-�ǪV�� �:k�v�l.�-�eM�v�9V�緷��C��n�*�T�]حY���\I�黬�[���Oqp�}�o���o/���Φч�]ίs����z�mJ3�ޮ#g}]���
�hd�*l��J�A�WY-�᥵�j��Z�Av��-*�ju�&�,`YS��;w������bz������4E�]]���UR#���v����/�e�f�jԖ7r����w�ZSrV¶�����TtgOzVm,�{Χ-y���C��������N�$vgV|d�,�cv�`�'��C'g��]q���/sC���5��3l:.���C,��gp\jĮ��=+%5]�Q���.gv����֨�r晼��K[�B�S7�_	kR�t	V��{�VpS䈷+�
s�M���ؕ����lU��{F�SZ}F��$�]���)(p*�f�w+����x���-�\Z�H����O��ڭ�g���ȸ]r���*��m5���Í�WrVK�T��V����Sh*�F�T�g	�~7����ﱫ�	��m���\���D���%.�Z���u��#���<J*�VB�Dm�Ą�������ΜH�2�lַ`ٯz��hm�ζ�m֬�I<�μ��{Konܗ���b��f�;vd^^t���!<��ћ�Iv�[3kkG�I9"#��Z��ml�fl���8{6X�'�;�&�$��3�{��H�ٜ�r��s����G qDD�D��$I86��jܔ�E��R�����w�e�m�v�@@��JYn�sm�W�ͷ%`f۳̤3$t��nC�km��r�:��Lk�=�z"��9m�۳���n+[��Z�����lq��AqF�mn���ּ��km�Y3�2�Q�te�oo{eM�ȷ��j[KkH�d��9-��m��ۭ9I�Qs����]��qJ�1��!#�jӜ9�H�6ӳ#��"8����'�&t�����kZ�e�qA�[���\s)kWYJ-Hrڐ��v�Fh6�v{$tJ�[�-��B�(�L������.�Ή
�i�\�ة�s�ZmBY���كcr���v{����x��+[�Iht�.�	��#��kK��bj`��t5�i�ȽN�B[�)\�P�z�ݰ�f�e�nV��b�`J<ڈ؋2XfS�K��qlm��S�eɰ��̲���X�0v�*h1v����ȴ
J�W��K2�4նA�n��3D%	G�k�5r�A�(q���ݢk,!�0hB��O�ٮ-퍌�a�Mt �Ա�3�f��L˓MR�˞U+M2�CZB[C.�)qe�	L5��t�'ib3B�4��ʚ	uM3Q�������h��4�1���ҫe]����T�4X���S	5`Lm��Z�3`YSd�m������3�1�Dٮ:m-m�FT�١
٠�4(������v��% V�f,ҰG�1������M.n%IJe��v�2	J��uq�A�4 �Ҝ��M��+[5"�Ҷ+�h�*q-�x��5.]Z椺j�݃L����z"*TZ�Ձ-��u¶�3��:X��"lgBY���
�j��dť3K/9[Hjd���lƠ�i\��l6;f9d f���0ҳb��Q�^�5�g:l*@g�-�)r���u)YlU�Kpk��K5S0�6��5u��w
��%�����w�=|���[�����q�@����`��䴬�v�LIpZ�5������$3
��1�� ��:��+j�*�!��Z�ք{ԔV���k��y%���*[�z����Y`����.e�Ԫi�a)�A���e��֚�.�G5/bcMz���qec�l�D�f�F䘭�L��4l4�`��R���Se��bIZl�c[X�A�"��
��[�Qp�K��k`Gc��{Z3u�1�-��Ճ��31YH����ЛP�v�3Ƶ�K�:m�f�:.J:�J��]���⌥�d��ME�qf�����y]V\�(�k�1��yc�#.�k+��X,��n��a����P��E\�;6jk��	��M�9�[C�K�jv[
up��Xk����P`��kl,�) B�nu*�����u:]���lb���v
�sfl���KLb&���m�њ)7��C�������F�XA�D����rm"�1�o��ҟ��,�H��0V��S�<P����lƌ��c��.��-6��f����6��=z���|[jH%��w+c�ѷ���#C���	��]��ݍ6��͑ ��A�Cm	�_3v �b��{�z���~{
���^ٝ�a�?����_r�A��k���X��pH5R���P��-�[�Cmg����uǬ����˗^�e�ϡ���/�{�n����ԑc���҆i�����=�#��������4�Lh��j�E��! �U��eg�����+��rn�[����I�ݻ;���H!�y���ӽ&*��V5�K�_Kh [jA��M�5�,�U.e�����Ҝ�Waع��*�&�+2�Qkl`����J:2x/��	�vD��/�-���Nr�{��ϡ�Z-o�V��̜�s�g���dH#;�O�6���ԐKmH!�u��O��E�>��Js�V�Wmn�.c�]��_u,�O-KV^+�N�'�V����+�5c���;���"�Q��f���B*�]S$���s�/���Ho�Ɍ|Mnp��-�_w@D{��d17+�}]Ro�A�ɐ~=Ѐ ���fd�?�b}@�����:����f��0���8�	�� sّ�9��3A��G�B�!�^�A�iȟ�p�̀��=���^�1����[�H ���9ױ�2#n����:���/�@�B �"�A�d�c'�r�ƚM_��B}o��γu��� OtA��s#���ϯ��}����/~l�\�S��f�Mn�Y�*�6�&����e�����eM�6���$>�aFj��'�3_U޾�ٟwz#^~<�;�-��V�ò�9�\F��r� �$V�/���!�y�$z�~��Ѽ,�� ��&��g��{�/Ŋ�����6�#3�n�B��^oУ��	�jH̀�̄A��b"/_:�Sf�'���Pg_���d�n66��&l���{,�W}`���|9n���.�el��Q˒#˩�3(���u����,�
�4K��i�;4cÅ�_o@Dܑ �B ȂI,Xܿ��+�,U貸f �!�ȟ��A]�v��>��Ca{<y�p?gj�ѻOY�tby�z�O_)��ā2PI,Y���z#�`��U��	�/��V��ќ.�X�p��	}�٨̩���-3�;�u�E���z�aJ�`n,4�V�,ҩP��4��^&�l�Lͥma�^�����_Oõ}���f)���%�j��U��<8[��Y�{��>��}�}�d�b�=+�� D���)?W	��D�_HƂ��݌�=]�����q�g�+�dA+۟�C�2���{{|A��̄A�B{�-��&�z���~�=\.7��}/�j3(�L�.9�q9����~�����z�s1O���8]�Kr���xp��;�(o`�sw�E^{���x���
c꼲0��GyN�mm�J$�hd'M��F�G�y�3tx�.~������L���U��Ps
����.a\Ɉ�c���8t�>�$�`�+�(aOxm�x��Ѩ'�xwK�������p�\Fdd ~�į��:/�򉂠A& ��	����+�T���e6Z�jEp�YS�d��WC臈o� 9}"Nd/�?f!4��w>ќ.�z�\o!d�|�ӫ1>����#_���@�H�d�ȭFQ���N
��6ڑ���S�4�n�xĎ��"���d5��*��"��A����DK���O\�;��� �|��9}E6#����';T��A�Ds1H#1 �
>��^����@��?nE~�AS�t��9����W[������O���Gws��F�+�d��"D2W#�þş����~S�_�O)�+��0��� ��JD"�&��B����񓶒�P�u�ٷ�I���������f�n�~�6�f��.����>z}�;ަ�>���k����%��X��tʰQ����ρꬵc0KZ�aZZCeasm���2��؅C��s*��&���e9\̙���;S��M�2*�Q��h��Ed$��4�*�+4�[r�с�Xb� ��ZًbX!�C;;B��R�oX���dD5��ƥ�.�
š��wk�4���D��,qfe�;:9����nVa& $���\b#N"b�#�3��ݞ���n"�6��߄������BUښե�3��q��674�qbUe�(]��!��}���_N{��>|����`���^�M����8���tN�����_3�z���z��e��-0�2����{�q)O�����.�zk��FW�Uh���A��D����#޽I�po|��@��ܷ��D2R���u�&~���㪽���N1��� ~�����J�d@I4g=���^ƂZ�ܑ?3C7,n���)���w�)"{:���[���#��)#1|�2 �d���Dwgm���W���A}z��n�VEp�Pǫ���A�:�@�̟��Fb~�tN��#9n�JKm�K��O3��d�j�\�J���Y.��1i��V����ֽʯ#_�ޑ?�e�2���r��mw�vn��)�S贕dM�@�=腃Ґ"JI����V�`���gb�v�}�m�nh�{�;��BJ���aV�n���fn��#�h�7:X��]ͻz���UL^�_��ڂΡ��c���^�x�8�	����#%*��EZ�`�}�� A�A$�I̅��4qn�i�S��ɚ���5��C���	�:�Dfd�ِ̄A�왎���sk�~�A��|s1H�81�򝛥�|R���@_9?YC2���[�o&t��-wՑ@���̻%}%��&ct�~_����(p����Gu������p毻��̄٘���0�t/q��t��"�B�1p�4�,��mCW�MFcXؒ�,#.�+��?�G�}$o��s!�A]w�^u]mW�{8^�H޻�.^r�'WL��l�?��̏	��$.+�_�f���"5mH�81��N���>)�{�".���T�<'���h��`�g�|A�A FfH��bs�^�s���3*�	*7��Ө��r�Z���4�8��{��#�������c�����3���tf�b���b���<���q����/ #%/���dH����k�:�HX|W�X ���?�� � ���.zi�c�%{8Z�	݄��:��1բ�#�$	���d�A2E`@�d��y��ߢ���NMp�K�~��d�8^r�@���f�eM�Y�v�����3�4�4ԩ1�f�ts{4�Zh놊�!N�p�������6�V��.�h"32D�sY\y��OM�&�z�p"|8�<��ę�4��~���e9��Nu[����|u�"�VΧ+�u�J�h��$�����bfe=����ed��Yc��q;�+ �_)	�.���μ��]=�4�L����|A��$H9����"Ibŷ�۸-Un��:U��A���b���׽�<��<5��� ��v�"�Q�;�кΚ�8���R�Û�wkqa�,���B�3��YÜ㇪�h��"�Db��3��ޣ��Oٷ0�̸�ywÁ}~5�I� ~2P@D���d����害ՉT?$n���^���%�p���H'v�����]�dBU���eY���ԏ)]��ke�6
�ƚAL�E�	b�M��F]	��SQ�ܢB���z��C��2<'3�����m�.�%!�����f�5�y��A=�����pG2�37��e\K7���������4�n��~�A{69�tO+�OMx�8�	�� �/ِc��ֺ٪����8�}���Ad�,%|� _{&�&�/��J���J��:�|��`��e���ML�.9�/�W{������ s1H�x18��l��2e�'���8S��;���^��c����354.eL��=�o/z4�w�����Ϝw=�W�^5�Ց��}�ʙ��#���	�v���կ���?M~��oF\}X��������Q���5����j�����v�:9)�v�oz4����!Z�r�>���[������r�Z]uNW&�$M#V�&��ai{Ee�Yn�d�2K�l��%!m�N6Ҍ�Yb�F�J�]29�ͦ��cDX�F�LͲm,4Wm7l8Όc6Ma��DWEl��(k[mz�\����]���d�a*⌵]�{Fm�-��6�u\F���t��ժɣh[��2YY�M,x�KL��[�qi�{��g�n��8v�t�1Y�iy;�>�>��[I�)-Ֆi�3���.;L,jܺe���L�GW�T�A]����d�����$�@���w��J���aCU���k5D�V��x�m�� a̅��b���^����2Ɵt A=���/'����&P�y�����_fGB��N͊��69�^� �{~�A FfL�D�-W�ש�����W��f?i�
������H7�#�#��A�%WQΙ��յ?=��������ˮ|"$���._O۰�"�S6x���}�cA�_c���AH��"+�o߷��٬{��V����w�k��(p��'� �ܟ�"�� |>�4u�����^`� �E�YV1,�lYzխj���bEZ҄Z�P�����K�ԯ�����m�]�xv��XKl���1��<5��?�n�?�"�H�H���~S�W�G��m���m������RJ:��wƘ�7����Jg���)��N���F����(�C���T�Z��#wsIC�[⁞����侮�U��b����s��^� �A|FI)��7�ۗ���}�J_��_��_IXAH��~ݽ�f߬��f7��5vx̣����9�ѧ2��Ybff����z�o����h G>��Ȃ���owi�_Y��=��\q�;������R����7��?�/���J�$���{5ضϮ.�}H��z��}E��m�p�q8���p/aF�#3$O�f!^ʳ��M~�A�r ��2a	!H0� ���{�U0���uW�n&ʘ\��U�mf����gߔ�o�G2�R�^��{o�����[ydc�V�6�-��pX����DK2W�K?�{r�Jj<��/�6���ow3�ͳa�O�}q�s�H ��̆��o=�1Iǵh��>�D�Qne#33S2�#�g�>����G��Z���WPG��M=o7�\�Rڀ�d⣦���0�Dhu�^Za��u�\hZ��h�����7���*���؎Ua��q/�vwR��
�c�ٮ�0�1]��`�gu�Y�r��C9Gsk�q/�4�'*�b��{�� �;��v�B�ҭ^Ån[�w5O��)�7��BܘS�4�x �ݷ��W4^r�fe�P��ۃw�rD��w�̈#���`�]_Ƃީ�ð7�=�ʰ�H�VS�R��W������g�Q�r۵���|�#�w`i����WT��������ɂ�Պ����������݇�����b)������B���S�P÷��"���n��ys ���eR�P5)X��S;-�
��}�s �����D��m,�]ip����]9b�5nV�˼�|c��n�#����o�)�ϷGr9n�9�<8��􍩦��.އ>ߔג��>��>���Vi����/�b���r�����hd9���ܼ��#7{:뷩νu�N^K�|��2F�W'R�SmE\�]�lW�U(����
-C�ԝIJSX�^��XAYx���i"�O.Jڮ��ꥸR(��X�e	{�q�J����������Z��:V�	]���%<ݧ�N\�zA���ʭ�y��2��O�VV[����66^Q����Jx���1�s���*<��왺]p��_Z��+tn<ɶ�v<�*�U�⦶��LV��vS6��b������]E��5�N4���`�H�ْ-�i����Vv�fWm׻w�ot�@kv�;����\�o�������{IK��ƧX�bU�|�h�aR�߯����k&��+2��m�mkk3�6�!�I6�{N���yd��Y�I	JN6�	�N�/o{���H�`��Fmf����Q��htP ��"!�Ӝ�G\�!��' ��L��Eoz�j)D[V��l'3m��S����kb��!˼����.ΎO<�p�Qݦ���I�+��:���VtgVYYĖbHN۬���#���w%�bYiL�VHkK:���������GE��V�E6���3����T;i�[�9Y�ru��۰:BmfTgf�/{�^�u�v&�l�yd$q��fՕ琧p%wTEǭ�6�q[��h�%Egn�]�d�]a�e-j�y����mgm��lq�j:���mj���ۮ;:-�$��fA��\)�����~��_!܂"Iw�}%g���z=N���?�3�����3��7�>��\a!�3�'���+��}��Vg�}���X�r�D��d�A�$z=��3˾�h/���oolg���q��w�8�s�I��dxNf.Y^��6"�>��`�`EL�D 1�aK�c2"�{E`ͦ+#�`Lb���bu2���}] !���dQ����c�W��[��8\��
L���;�9�UD�O{���e�ʱ��qտg����[����p��[�b����@��E�H�dt��J�k�sSC�)@��ϳZ�U���,L���fe��{�J�r����Q9gs=�σ��Gz��r�A~_IX&H����4�4x�yA|CƄ���f ����c��g�Zk#8\�/a Gy��k�:/I^Σ]��.���v�ț�����XΕKz��\0��h�l��ۊ��lU���M�����䨇4�p!��~ހ�̄A9�����2)�#�7�b[: T�,���Q=]�#�%!��@�{�"��̏�وE��ʕ�2��z��I`F)�S`s2�i�̱t�1��hF��ݳ������*m	>4� A�#3&~?f ��lk��s:σ��G{#�QםB/��m��Hu�}����e��R㙗���b9�X����%����#գ\"j
z���V��6��_�����f;�q÷����/U�E���3,�2��bu�Wm�ܒ�9�ћ��ड�� �@_~���̏��@fe}#\�p>�����#�]��st�5������ɨ�dp ����<��r����0� �kV�2PD��,+=b�o���N5s��!��1�ם�E����6���"H��"zV��#h��E*��72_��(�3�kOS<�{?LF��M��=���J��]�!����hc}J���6�ڭ�,�5F�%����]fi`q��^�mS�ZYX��!(��KK�[m����v��F�SWK��ʂ7aΌ�u�n����W
�veI����,��M�;��)gQKH�`k�a��݉��3��P�,��R�T#f*��/jB]e`��	HU�3Y�����Re�:�*%�&-��]��svL���-�3��sqp1n����-1�ϣ����,�[���vek��֠��iF���6Ȅup���("�.�A����Gj�2=��b�=O$�3�òx�(p��*���Q��@�o$OǺ����̙��?V9�U��	z�g�3P[ouh}�Y��
���;�ǻT���C��;��κЏ^+#ޯ�P��X����!^e{�E,�*ǽ�5W��ΣQo&/��� ���;�.	��5�,s*�_|m{��H#ւ�����Ľ��e�޲�vbB39���Lﾋ����_�@�?r�%�&J�H�"H>��֛���1��Lf�VN�UX�dp ��S����J@��^�x{�ؒ!M3A`$Ԗ�!`]�z�%��Z�Q�Qq�,�K#�-�Yv�!�Z� A��H9���Ayn������y1|%�H[�o~�G��"�7H"7�`_�D2W���}V$V{��K����':m��a���j�q+��մ6��z���[zS[}��=��r�*`�r��rS��κ���p3�f��&X��z��2P�� Ot?m�9����3o�!���*��X�~2R"JI��q������Q��U��*�w�8�����J@�$W�/�y���_�wB7q	����&8�����7nM藜$�l/�HVZD[k�N�=�����d��H��#%;�s��Jw�&p{�\<�)(h��Ǻ��$�@�������Y��+����L�
&l�lQ�72�5�%H�7V&�[r�K���GE�r	�����f/�1�Ǝ��g�����{#��[~��9��H � �7о �s1}�Hd�Tj+��G��i�˹��������v��	y�	��@fe���2R�uo���QD�o) � �d A�^kW������3k7"yQ~s�1k��^d��Km���"vN���������H���G��c:V得��E:������'}���=�q2����0�ʒ���}�~����M���.����..�A� F��?�9���/�Y{�CUcg#� ���H�g��}�4"�_�Q� �r�D�/��� �$�fJ����Wy=���R
�y���8xU�F�K��A\"m��?f@���������(]��C�4W�U�d-2d���!�ۍ2�Ɋ!r鶉P�ߔ}�ߩI�2 ��3nї���z��3�e����Oh�>�����e�"�D�ł��!E�ϽW��T�Y��"����� ����>�˞$5V:r>�w�H ���9����Q{>���niH#5 N� �2D�s!�g��k�'6#ҩP���'�ǅ]4o���$=_.��o���+>#��_F��n��S �H u� ���@���~;��s��#�g Ot�f�Q0�7��P�_���lr����;[z�nl����������*��tޥ׮˶�]�7��d_[
+"��9~����[�XtXs5��y�X���H�f`ҝ�{'���`gf^���Ud��`�dp��� �z���B ��[�������F�'�H��X	���d���2�E�Z8���%��\Q�R�Zmu����>�E�u�9��́���/zc��®���/:Fg��Я]�Z��{xg =辒�2R?I���I�s
�}��v���-��fX�6�Y^24^w����6�	9�o�n�foKX���Oj��Dfd��1'�����s��UY!�f�w�8�����̏����e![TcL�٬��y?f��yhי�8��п+��C��/���nc3M��*����[s?܂9�� ��_Oو#��Ӝ�ó�[.��7n7_��#E�����$�D�"���ށ�����W0��r���ދ3�+Aҝ6t��ʡcr�+y)�
�8or�/�Q��w��T����i�����5��u�����}�׳elv+Z,�34�+��kf�1"hn��1�6�1��Qq��A�O���,�Z��ݮ��p��cs�3�,&��e��؉
�X���*FLYt4�жb���4���YB.���`7 f<��)M������5.�Aن�$�R���ԍ-ҺXAy�P�Յ�����c���i����#\��.i*2�Њ�ȻA������o3F��k6z��&527;7K��	u���e�9�T2�������~�A�32D�sZ�i�ޅU�Ț������8�:]K�3��w�	��$fGِUN����!o��@�ڇ�Fn^����݉�+D�C�;���#3<�뵺�E{:v��8���b�D�/���"����M�MUw���^\ݟ��g�#��Z3��L��D̲�35�z�b0kP_y���A ݾ�{��NdM��dq㽪A�:=�#�ע�l ~���e�dA�"NdW=u��G��-\7�l�T���0�p�hp;��-�32�㘇I}�Vv�(��AASWYZuu��Hj�9�	M�2�6m�r,&c�-Ѵ��VS�'ϕ�A� �����z�L��}��/9��[[��!��Dfd�?fG�+q�\��\�Q_��iѧ��[4tR��n��r�7�h�+\�O��^��U��b��j���gGa���,{*�*��Cn�4�]Ż��DEp�����x��>]�=s�Y������^��dgy�B������~��ֲ��r��}�."ff�eL�5���;Ywa篥�N��	LW	w�A��ԁ�K���}%`#�-ਦm)����}H2Ec1�*�a��"�!���|{� G�����w�c�Լ��	���U���X��k�(5�������v�gxU�<����dq�S��̅��^��^�Å\A��䠀�@$�J0�3���fl��
s2��%ƖL�@��WC�����~���ȟ�d/�9�/.��=�=W%1\<ﾐ�Q&�F�f�� ����dA)A�/���>�o��� A/�z��l��"�H���'� ����d{�k�LH�_�_tГnDE���B�"2��r��"[yYH��7QUm&�[�EOA�N^�>ui���qK$��x{:�q���<�v�vn��S�=��gR�N����sy���*/!�}�7�A�W��) A2EdH��-�����a�t<A�?�@~�Ayp{y��S�qRS���N�/���}|TSD�b����@� ����$W�P@�Y�����WnNf��)�����;s��,p���~��M�,�9�h��t���~?}�5̷a�qfL�b03���IV��F�E�Un���BpEb��7��@feO�f �o=���.�0w�;�"��h������A _Rd�ȑ ~2P����~zN����7�C�Fm���]WJa1\<ﾐ~;��p=����$m��x=��A|o��ܯ���+&H��	U/:5箊~�}��"E��8�@@F�Oّ@���fd�!����w�=�*�":�g��z���w��f�G|A{��F�=&����4#���l_�� B6��`�K��֗חyOD�E�2�����U��/�o�7�N߽�"��j�ܤ����i��u	���a�ǰ�������~<9��"<��37b�Qb&fhәG������AR�z�r�_�Bc�=����|�A32@���B�Q�E�J���_G�:#̻����W��Lx��M��:WM`��B�����mm�������ӥ��}c~|��s1H���Vy��~�$X�y��U��;߿Q�"g�F����̠��7ʴ�����z�w�s�#u���5=���v���}�;�'{��/` s#���fs_V���֑ڂ�s2~̊���m��U�ЯU,쥷�I1��}41��ݢ�ff�2�ʴ�[�}V3�i�� ���~2Eoy�e�q�w�Ⴥ� A�N���o�Z�{��͞�4���;�M�~2R��"H��F���X#���uw����T݇7E�zD�Nr�����@�I?��BI�$O�@�I(��BI�`H$���BI��	'��	'��H$�@!$�h	'�� �z�BID$M�$O�@!$�0$O�@!$�$O�@!$��H$�� ���d�Mfqvz��O~�Ad����v@�������                         	� �tQ    � �$
J � 


� �  P
 
RY���(PP**@*�R�$(! @T����(�� �� 6
 
J�
=�4dZԩ��25M���F�M6Pd�[�L8+fB�B� r��ԎpFdafԕٟ
@h^�� �� ��`S��4� s�T�� ���Q
��TM4G3T�d_^sJg�M�v�l^LI�j��H��Z�U�@ �� =x��������E����n��鑤�j35R�e P |��h�J�*J�@�/yF٤r�S�B�s�S-R�ЧL���x�/%����  P/���3U�����
��o
Lt���(��]2J[�ĕ�
��]iUU����@P  ;�HP(RU{Čؔ[UY�Hd�SpC��l��ƨ���1����r�]�wnIUJC� U�e*�j�U�T�x�f(��eU�b�f�U+��9=s����wJEݽz"���P� �� 	@QW���@��ԕYiJ2��u$Õn΅Wv:�.mIU��F�Gz��w���T(à wU�e=�uIM��Q\�̕]b*=4��mUTܥMʪ� .���/`4�Q�    ��R��i� 14ɣC05O��JU(       ��UJ���@ h     Od�L�J�Pi�4Ѡ0����IR��=�4� ��4��i�D&�Ii1	�&��1���M=G�lj�jO_����O��n��K�w��hƋ�,z�!I��(�$�͊*H^�$��D�Q� "N7�O����G�����k�M��� �C��	@#�
P��4&�SHB����r��������^��$f?L��~M5+N|>���fT( c|�����\����U����5]v:k7c�.cA�J� �q^�İVԏ�[0+��]Iv�P��m���-��U��9��5�BL��t#�7��bz�(��ƍZ6�Ҫ��ysF9[VK9���Kpf��0�;�3EEg/]�XuYT bn��Oe�3V��IZ�4����u���4A�Q����8�vְJ�`�r�:Ֆ/D��["�Zti�ې�q�"S2�e�.#6�=Ʉ�5B�mD��m)�3	��]�Z輆���c��/�Ke�����i5��Ub2UV'W���� �RXy,٘n�طu�'&�VƓ�&��^�UF�6�a�;�����4/v��z�����[Y��k�^P���~�X4�ӥ�WKr�:36��+jz�¦j����wv]U5C-����v�SX���y��i����[� �T���v��36�w��h�mR�NҲ���ܖL�wv�í(�Em�&�ڋW�B�Bs%�v��e�a�[�nͼ��#kr�n��ǵ1��&�d��u����(f��2�7��{B��,M��h.әTV�"Ց��R���%2��5�����N�3H,LR�^<�B�R���Ѻ�m8i�*����Z�(3�<;P�&��;��b:��QU�/0L1m�,���J����^�n���UIdbV�$9n]�pK�:I5�^UL�����[N���9�BnakEF���H���Q��5�f��:�Û�A*��.�R'j�S.;6h�v�nVc�H�ӪK	��Ķ�mi/b٢��-̗2�^�V�S�Y��т��ؤȴ2b��>$e�L��V��+6|��4sV���$�C):hՕ�Tm۔�2r��']LOw.�J7eL���(�cb�Z�bf� ��,&��}��f]���&�hړ\�T̒K�XA�e㬒���u�̹���l�F��y�=d��F
	d�yP�VR��N�m7�H���j�$e�y��XM%����Zj�7Y�[}�҅\[uF��N��6X�CMQ�6�h�uI�[r�Z��ճr�<;U����F�i^��r� C�f]�i����)��c��@I��V��A�ն&�V�f�(n@�n�㱛g4R�3T������i�K�÷u&��5�Wʰd]�eK�n�ie�/t�J��KִiیZxt<���	��z^eUa��k+��T(�ʏV%6�+/VehtU���E�L;�i�Te�[KJ捘L*���n��Xy��jBmI��)�*UQ�HeVU�n m
���ku(��R��)��;zfV�bΫ���K4K�5}���w�U�gb3�Z��6�d�z�-�ۛ�n��]1c"Ș���˶�!�#���7�{��b�`X��lLE&72�"��h���Aw[I�o\d<Cj�V:R�f4Ԋ2�Efi�{ ԕ���kpEZ��Y61�.c�TC~�q��k�Tov��.�-fl���]��ۨu����DØr��%	TCY`��nPϞ;��x�\��oj�L�ݸ��z
�¥��x6c�̚Ј��(�b�.�V���&#�*�n�^f@Mʳ���ϊ��-�(c��J�7��ʭ6k*��[7�T���N��U��fT�����r�]n��6�䙊���gVQ����*�W-J�2�n�5/8+o0�Vh-7�ݑ;�ܻ�����e�d��M�(�8����F��G���<��Yw�x̽[�)����6m��\s1��m8�^�
��Sb�6T�䩬�nދ�����(�iHk#��d�'l�iϯq��h[G�݋4㽕�4ëST�4�d;Q����4�kt:c���uuN���/�2�-Zt,bef]+:VS��c2���+V����{�O���D(��i�](&Q.�bnS9Q����b�TM�j�q0sM-�E�4�[���-�.���S�U��Ա�ssEL�Q�0��`S�~b��ٺa��j/3MGK�[P6ͅ�(�t1��^Ǌ�5�̻/ne���a�Лy�ڀ�qd�WE��W>�_LQ�V�o�{�v�-˶�,�L�1wy@��TB��?���
D�uY��)�B�A,gBq�j���BR����I�Hm��H�TM'L�WY�Y9I�����u�G.+��OwtM�����fҩ�UN�b�����X��U��CT�@J3��F�v^IU�W��n���n^N:��Bfba�4^bn����bn�J��Y�_�U��g�sbAZ��kk��ݒ^޸�7	 � �3s*'��nGu`�
�s6�ݙ�]�w3btvV�y1�N�ҹ�Z�^c��n�Jխ�P�q`�N��I�*X$P�j���U3�*�ٖ5�X�E��0k��M�Ք�)4�6��R���X����ؠ��3d���� �Gi�j�"�ێ;����OF��ޝ�0�-���ɔvk���%��-�cմd��l�F��r�W�7�6%cՓ(��[ǻI㩘P���&�FeD^���[.Ы�Y*+ke�*f�he���k��ʮ$gQW�9�KF���b���,��rW�]�l^a:��!I̊��̲�NmƮ�䨲Ɗ�m��8�N��dw��Ӛ&T%e�\wW5UЊ���%�y[�+��B\ۼK)n:�`��m<^hpb/&i�5��UB�R���W��)R�*R��Uʅ$�fS�m"ZDVM%�3,������F"�V5z��L\����E�͸�Y��jU�m�р��]�̛N+�o,�8]Ǒ�V�襑^�J����t���Q�$/,�:+8�$�)���6�]1�{z���ɹ#���L��WgV9��]V��$H�r�ssovTڤ����u�
�Lڦ~���2FpY��4�vv�fDD+Nص��f����m^�2�5u���Qf����M�Ui�(zU�*�x沲���M`r�hp拽���۰U
:r��}�ŉ��
-/~�J�]^$�ɋjJո6Aa�?L)�T�&w�{��Z�Tr�X�)1;DT�E��M�z����jd���D-�QJ&�*����f:X�1j�����\��}U���˻ha�De��A+�@��h��2ek;65V��0�6me�kx�ɂy2ڃ�&&Pɸon�ͷ�6isM�f�@�M���Z3p�n�x������y7m[c/HLfbD�̎���c`�H5=5�4�B�:���e�X��qcwe��C�ٹ`�j���a�e�7����]U�R�����ueҘ��aB��T9��:����Z�ڋ5�[b)#4����&I��Q�sQ�Œ�ȷ2�4[&����T��H��&P�Q��Ti��Qcwc��
9ۡLh��Q���ccf,����5�V���qɨ�U�0͢�˒e�7�q�;�D驍=��e�6���"�U�9�淄�۱�S�rV�P62�P�K,���&�j9b�X{�噛(5��n�Q��x6�A�,�pe�����RŸ����e�PY��'Jѻq��j�εR����S^
�J��7hC��Ta�B�cI�2��\u��K
e�v�VE��(TKl:	*�V̂�R"��ū�8�kd��D5��w+(�XoA&7�icc'��N+͛(Q#7u(O����-�"0Մ�5���a�H����-�SiMz��GB��Gw֢������#�U��Y{�MRgu�`�v�W׏f��X�9y�VX���OrGf�D���B�����R�e�5��w��6��M�&�͔+2Ah��m#/f#,ս:wj-��ֻ�ϰa�D���#
��(���qL���F�h�V�����ǵ[m�&�T���K$��u�L�Ϫ Pr������X���K�L��wc3"�����Q��Zև$uw�jn��{�����/�a�9�X�{�����~�m�;;r�+fɕ�MCXQxs1\d-)&��t�b"�S�q�xB�ZD��:�[�P$��N���z����K�
�Vbɵ.h{��4Z4�d�Z�Jֵ��춍a���%��D^�yeJ��X�@v��楏*�d�*�e��ѹ�
���1.��«z^۳XVkoHzj�UUw[[m�:n�j��Ԕ1�W�����B)�+E�:凄*�TS�(]5f�R��N�Q�3$L�4�:l��)UId7���Q�����+]-z6-جWW{�4▨滻�Sy�[)�2�Zؖ¢�GkcAZ-Ui���;"���S�e�KR�j4���Q�zf��s/l�̼�v�oت�"�fӖ���z*��T���{�U]m��Z�v���WG
��,G+Y��`�)ؼO ���*K4��.�DY�pۋ)]E�70��T9�`dǔ�e�.�oUëdi��ĞAx��F�%RV�N�$�B�*3N[Ϩ�����רf+���Y�Z�7�^LwvR�uK��NI�g3��.�0�N1��o�T��6�dm�8$v�Es�A�Pf�C/.�3B�����ŕXIL�51m��+q`�ux�۪��`��e�ɣ����-֛�w�+t�wEM¶�ϲ�++*3�"t��Uu�5���z�ە(Օ��5�0��if:A�	V�V*̳j�mѢl!�7�LA�siȶ�AѲL�32�ûX�a��@˂�D�L�Bպ���3(:���j��p�F�Բ���U���-t#-�;�L�a�m�>����&A�ozm��A�ȒA)^l6		6	�@�w]E]�wU�W\uu�uW�]�Q��uwwtuG]q]t]��w]tu�\Uwq��t]]qWtuw]uuWGwq��\]�u��q���]GwQ��q���]�T]tw]�wGuU��Du�WWu���u�wq�Tu�]�ww\]�tWQ�wUEu��Q��]��w\]WEu��Uw���tu]�Wu�tuGwwTWwpm	%���z|to���'��O�$�#�f�;���@#��P���'�ԡ$zX֏���C�=s71�K�2yh��9���uG[��0\7V��ͺ�z��
��.G�8�R9wՈ�v�T�.�fo�oe���j�������:��ө�в�<�W0åad�����N:YYd�h9.�;u�u�j�S6N��bV�c2L�MԍeЬ���`��wV�!c���ƻ�ܹ���72K�1S�C��R��x�jTR�2B�f7qM�	41A+#��p�"�;ܵ�b�{ ����>meDw��B�����-���������6v�]�|'k�ʺή:M�X��e:J��l�ɼ���'ך�gY�&�ʑn=D����s&`��Q<"�]�4`WJB{���G/y�n�I��]��/����3Ek�6��Ǖzlѫ���T�[��eS뭖�Óy��[��9s����q�J��7(Fαi:��Kh�[9���] ��%{r�^i�쫸�k���-�����ʶ��V����.��sj^��2�n�P����-�U�w�j��έ�������W�>j-���$����iđ��gZ�ڭ(><@�B�L�5+B���È�T.���˓P�X(���5�-�˻�bUQ�7-�vk�mV��u�t�����}۷�G�l"�vޛ�re%v*=K��:�KU����ve�n�ݼ
2V�/(�� �|�[�E`U�����AnU�+6Ml��J�}*�Vm%��l8:��c���F�P�j7�38/��ɷݝ��X�]��kʫ{�ur���ŋ�t�w�v�t�UUyl�e��Se�!)2���u�M�5Ԇк׵��ޞ�-;�8N,�)C([�Wi:��Ԗѻf<Kn\�r,0�1��k���Hf9��1�օL��u����S F�3���ZJ�.���5��U�([&�pZ�5�)�f뢪�d��7v�nungqk���jڋ�H��۪�������U�ق������a����i�FTV6�]��oj�䊹R:�PX3���b"!�E��{>mj��{uy��_U_�^�:w	�5C�u&�S�qL��RTur��S��[�!�a9�6m����c�U^Ur�2�^���-�Q���9�m�}��)���Wy.����<^ժ�����=��@���쨖�]W�7�xk��_q�Tv�l����[]2m��Ů�|sqt�s�q+j�LS����KFV�mm٭3��F���CP����jS���:ֱ���ټ�$�]I�Y�O;���⾭�0�o���zY�SqJ5R0�-CJT'�r�{Om�u��ʋP4�rȒv�
�$�T��Q�S\���w; �U����l�����\[����_McC����UGwFm[+v*ڗ%�|��+o�8U�eR붪�d�/s�/���xE=��&�5N��;��aٚJ߱�`�k]6���^��#95J���T-�ˈ%)='d�gE��R���}�hG���OzP����+{��-@��2sjԌ�8��9���N�7�i�3���fD�la�crd^D(f��DF?`�r�wp��۔�N������P�M��!!�P]i���Utv걪�k]-ܦMV��wr��i/�)�ј��љy����qe֌&����������}�z�R[F�ޝ���t�̪JfEP�Z1���,mG�úͽY�Q�3{�4Ց�hj�rC���~oi���OF3x҅/.�RY&��[n�>ݳ+����J:qce�e�z�N�%a#U&�k���ڡj��ٮ�P@��[�YFv�'v(ڭxsj�v�UU������A�-�uV�X�]�ueN�۸Q]|�n�UQ�"�n��g^o]7�x緮���t�g=����&ѥ/HQj��VFx����P�a�%�S�H������7�$Ind�yv��3��XՈ��+w���;�,���r��\#�h]�9W]���*J��T/����
cS�������4�ܤ�[%P5��ג޹ך7��&�ú�q$YV�wI��� �{���(+ZoUh'�Ư]����J�ٕ�J&hw���t����p1�C�
���0jLn�8�M��&fv*�4�Mk$�QcW�)��O�S"��:���k^�5�Vʤ�����lu-�5ݤ�h�jf��]m
�^�hXs��p� G�;bn��(��y(2	07�����h���i��w/#5�8�nn�.�Fe�Kq�hC�78����o9��7l�1�������*O
����8fAtqZiSxW� ��s;�4�'��B�s�,���dQ�}���V�����7��lo7*Ua�5$ͥ@�Sn��ܦ�Ck/��v�\��l���V���J��w�ni�9Fr0�֌vp��&]0f	Y�kE�X��@���\l-3����%me��1��f�W7�ug]�����9�s�=�Mh�>�e�u�5�\�^b�d�( �u�C�����ёZ�\�`һ�|oFf�M2*���A邚�1	y\RW&0p�| �Aђ�!c{�$��F�O�j]��W=��]%fn۠@�t�[;0U��ά__�k��%������7�s&U�Q���9f�vO�W3��w��l�R�h�j��wAYV�ٴ*j���p]�e�1h;�w1�%��"v��k�5��4Můsz&fQ�u-e�a<u}Z˛�w�0\�e� �[����v���feֶŘn��v��K���f��Ð�!1�c����$�f���yꕉ̜����e�dfi��:\d5���:n���TY0��u	}i5��2�	\�Ǘ�Y����&�j�y(0YWƻO��o7(-���ATn�Pћ6��z;^P�ZL�K.�aѝ���*Շ��b��b�Y�XS2%{L����nŬ;kY�^"ܐ�Bv�2�	�WA{WT�B�v����okL�RМpjY+V�O��ł�n��ov���F���IWNVpǖ���7RCAYls�۳v�U}/�Gʫ��I�u�/�fe��Ɯҭ���V	ڲ�r�GtZ��1�R������5ߦP����r�a�?QL�{ ��*�nt�mn��n7�Hh,���jlf���x%�G��Cis�n�K?^�+�-���3mVe�׬r�����C`��qrg#�y���wuN��cٜ�[��co-��0���\A�2"^I����nQ��Y�\WV<������].9o�����E�ډJ��,���)�.�w���⁭�7}��V�s�H�R�YB��Ḩ����Q�C�k�.�N�6�Ֆ��]V9+�����WpP���M�vޓ|3%��w�!{%V�6j�S&>�1�=�������՝U2��%6ݪSFrH�����v��.�0�t˕|%tv�{p� y�F�5a��ʪ$�ۺE^y�!l��c�b�Ro2�o�$+� �Q��7@���T8��xv�#VK�˔r�Uu3^�YÚh������9�4`͇Z�m��\U����Kv�n�W)SF��u;�*���UT�
{w����ť�u�1�D��;S7i��V˼��5��*�^J��$���Zn�j�;L���N�"�ɚ�@�PMlV�}���1�lsm�gk �C#�TK�T޴���<�Z�Эv�㙋5���+nv�l����*'�CM�4�K���)Lڳ��<v2��e|�͵K1�ڻ��튾=yhMZ�V�^Ь�O��;#�c$�=�%кj栵f��*����A���X���C�N3yh]Z�?U�v5����S-����٘�u�++a�iη�����9������2�V��&�n�v�CZV���]T���V�]��n<��#5��iΗ�/'�o��kl'�m��6�u��h��}���꽛��T��_^oAs�����K�i�(�/,�E2y0�}\�d���Q�q�,f�y��)�jZΗ�kMQr^d��]V��sAB��V���ʱ�Fң����M���'ݦ��H�3�³-EF��^�j��ăE��xo;��pe�S���]mY�b���|�q����h-t%�:�1:��f�
E]L��Y��НͧZ�싚v�Y+$R,��N�N��f+�J��Z�jJwK��s�ރ�m���']��C[R��ww��Uf�a��7��EUi*��UV�^d9���,U��3;��M	S���gm�"^��"c5I�#%�Mi�M�Z`/+H�R���yT	W�ᄑ�'SU��.wiH��Y�r��@��*qv�L�
����+��un__CV&�n�̨�.ӡi�������}o;+�9��#h�q��;=1��1^����{6i
R�K9i� �ti���ή+*��'����Г4L��8�׵�Քn�;�f���b+E��0s*^�-	���c�%,#)��ܮ��R2������we�x�P�Yy���퐓���8��ϯd��I�0Y�W9W!M�2�Q�&e�f<�+*�8�lF�j�J�f3 =qp�83y�k���^�}��Mf7j�[G"p�4�V7��rĪ��WYr�f;7[�6�~�ZO^@P�q�+�Q˶��(뮫�ϻH��!��r[�SQx���U���6�F��k�S[S��{N������U�c��k��}��VuQ\i��t�#.�}9`qZ�L�ed��Js	Ą˂��Nbݷ�s����/hM��ђFB�pX�^m%���ޭX�rT�]
����y�ׁz�$0cho�A@$i�h�����4�c#n$pT*"���*h0j�{4���ֶ=.�auflq�ܕC5�1[4��5;�)�al��պ���le$�ۂ1��=���{v��4LK� �Evf���@-�F	n�`um���C�7"ei��Sr�\��ǔ�s/0&�n[���8ۇQ�z�Rp`
�}�膸�c%��f0��q��1c8w�d�'sB#��� �GD���V�n��5֍q�k\�����qq�5�P���U�ZP�9������[/)
m�0�96I��\a^��I�mU�kQ<"4�CZ�_�������뙝Z
K��謷�Ʊ�����&jG�ŷ]Xǝ�i͘��1�aM�
3:�9���t�g���q+�q���l����.�w]�m�t��C��k�Q�9�4Y�iE�5HRg1�Ј(�-��ݺсݽ��N5I�cq�	xt�x�;I\󹚣e�L�m�lM"y�GBl$��<�����v�^��5��آ�
;�!�c���GF���m�\�F� � �9��g8���:���7[w2�]���(�]�ܒ	ܑۣ{sq���n�	���;��S��5�֎(m�F�Z���,bf�l)�6Wuk�6�����g{G^+#$��\ºj��k�j('�۴��vӡR7v��q��ׯ\z��]��Q�c��v;��´y�a�.:�˞�a	��XgR�XJ+�M��&�n�Jq9ɸk�OB9���ԻoX��vC��U��@��z��u�-��O�5�M��`�W8�;��-�a0�+v]GU2�>�,��7mskmd,m��]a�N�ml-3�s'B�B��z�K��ۈ:���s��e�K�@h��zR�U��f�	:Kĳ[�JÑ�,%�Z�%�S�,����b1��ܭCeZ��n�y��jX�ؖMX&�R�z�v�nF8⚐QNy̝��N�4�u�nݽGm�nc9��m���0Wvм=u� qKЎ��Sہ���V�nv#�[��Kfҡ����ˡld�,����q*���h�YqJ]��лgv�u�`���\;�;*�v;h�\D�r�eu\X�������{�:�u�={	F6�:(;`�v�򲍒�н=q��n6�W�1�{ri7�^ c�[&�J�>Q�9�����I�=�hq\o*=7I�-�7���z ���dp�f�:&��ʹ0�5�e��FK�Z)�l��̥:h݋���=��/g6Շy��<�i=��kCuW-w^���M���ᑙ��D��j��J�(ipSA&/#��C�ݲ@�17N�a�;9�З��L4d��K�p���.֗;q�8�0�z�U�Wn�v���s틮.�nܚ��N�Rv�q�R���N�u�]�;��A�J7=����F��6ۘ6��J�K6�g�Y�����s��͐��Hca3M�Ɂzƻw�#���L5�A��.͚���	f�2I��tH���7R��Jk����vs�E��2�iC@��6�MKl�&�+H��wQk�x�9�L���Ѵ�����]��6	��!vۃ���'P�9&y��3���:�9t���� ��x��)=���49��Nؗb�XCCkV2�ؽn�ꅯLK��J�-��!���j�<AMƕ�׎e�k����\�6��pG�/�=����4hXnWV,����"��Ʊ�7s�LBibIA�Zu1zkac[i�cx��+�lܡ��=mrvB6i]í�ѸJWF���p��bQ��k�q��ܵ��WWnR��-Ѽs�f�7��-и��)�]���5%�d`�
Mn4���͔���]+Ќ�����4�H���v�l�6�V�H8�
����:�K6��ϟ;���h㣎x�8�����:ѡ�nK�X\Aq���,�j���c�te�������2��O�:�4����q̔$��8���Wˈ�����5��m��tK��i��i6d��v��h�1@�u�(ø[���vݶfٚ��Q��^ �v�i�w���!���������xgg�x�8�N덳�ݫ����y�X8D��0���&���Ÿ��6񀪄�������^%��9��u\F@Sc��,���v���SF����I�yp��\7��^�[6�X�4[��)y��5m��ϲ9u�]m�nhvt=���vb��se:)x�Z8������p�w.(�{��l���ps�۟�N|�����	��lL�n�%�m
�p�źG[�:������G��� Hc&���,Mp���km#.��/	��ݚ��v9v�Xq�o9Ŗ�F�GPKj�.�L!�]mKc�LB���#ȍnF�ا��#�7(ۋr���tuN^i<ny�A���d���1z�N�/S�cܜ�YKftx�ĥ%��y�������X�s�Sc��h��:C(�9�s���n���L�nX�HPTє	�;)7��sTvz�Fk֋1,���KL�wd�.���C������G���ּ�>4Qi�U�[�ݼgkE�gy��#w1mհ4���Îl�D�q��=�/87\����j���s���=v杠wD�«ڭ���<8[��aG��nl�S��'�s\,GR�Y���]��۬q�TP�g�z.�����#�����ރr�-����Z`�I���!�2��Z�ɀ�݄�;�=�q��c�8�OPl[��R��S�����ccv6�TK���vE8]c*F����b	�ۨa����_��z��	�͸��R����v�l�[ە��qӮ9f�]B�1-,ń�c�/.ҁt1���x��vg/��brv��N�r�\�[���mt۷�.x������\�vu΃��+J�rغ�=�tuN�$�O<��m��.�檆�X�pvڍ�������V�j���r��l̮���i�������vh��
n��"m��I��9�%Vj��W�q.t��>���t[��v��ڂ;D85�ن��y�M��f$�����5����U�v��@ZD�B�]�C�;���H�7�-�\�`-Z�î�{gv뮇�Ʉ-�z���a\�b�J��hG�M�n���L�n:^]�]A�vC����`�wWP�����Y��]��V�S�۪�U��VC�:��Q���k,]W&�'3<n����qW8��5������u#���7���v:��+xz�9]�������|�ٓX*�Q�֗\��^��&嘰�WcDW= 5���v�j[n�y��K�����r˳F^����bKW�����n/��;=�-{E�i�w��y��� sk{����;k��6��f�ȳ�ś���6����ݩ���ː�:k\� �&ZS��k�$<�$��6�"y�n��y�%�EGgX��NIs� �'#�_k�%���96�:�;�N��ވ99Ӟۗm�rr��&g'ry��6�HF�h9�p�8���p��\��ٯm��׽�$�ǝyg^g��@)l�$u��=���[�m��D����I�����A�7` ��c	�\�c]��\�ݳY{Ѽ[&n*m�+�n6YM��O�@ֳ�yLѰ��zѸ8�i���5��c�p�;�Uꗎ�p��Wk��g�^SX̘�8P�f���\�{D;<�>Ɛ�M���l�n˖	^���G[�cv�	�t\nkqe+a���e4�M���M�㮙r�ܜ�ծ���,����U� LYL;\��y�\�l�]`��Ik����u��#cp𯹠Z�+k72T eɇ��C'j5�a�ct�[�>͸�|s;��]ɸ���T,����v8���X�Cx�\3q�<�֗���V���m��n����V懍>�wi:�m�=�Pݳ��������/i5�n��i˓t���ꭆ6�v�b�OcpV�kt���Wn��ݹR���/(fJ���i:�b�ݴ`GLM�1�lكr�D(� |*��k�86�����y��,��l�f�#ѡ��bL�������5啒��!r�c�,��62W	�4��^�P��B���zNv�Wb�Xn^:W��#�bE�xɺ8�oZꓞ'n�y$5[&�.�gVC�9��\Ye��Γ\�S�m��b�c�[�IAQ��Wcb�]z뛰�X�5��\)��������C��b5	[-xҥ/�J!ek	k^
�E)U���(J�R�RR��@$N5ZՋaT�-m��U���%K`�vۗ��3�ypg��!����Д`D!Kĭ[a�l��}��X�m��	M��2��m�	�q.s�`݆?�?���Ǘ��mz��6�}>��/s��yE_U��t�s��:"����o8�{Qβ�T�a����m�^�[ǝ���Ź�����6�oyOI5�ה_K�����������uN�80qΒ�g��nym��nWOe?{v_�_��Cm�f�y����o�ٶ���l���S!]��U ���� t_=tܝ�p{��xku�^���_{�2������U�e���ګ�N�����N��iN�+�g^�<�)�Y+��9J�VN��D�TH���Kg�R�]�m���U���
T�g�pl_kt��=�oo�[�t��ݍ�y�m��aN�o)n�)�5�ԛ�=8nxk~�-Y��O���o.f���O1�:�õ���U N��ؾ�>���sv4��jMt.�LLL�$O�Q�1;\(Ӫ�y��?vo���ѕ��%�h�96�3���B'ku]���������*�R1�����c_~m����{YY����?c�2���w1�յמݱ�y�ԏ�a���6��nz���:9(��Zb���˰��R�A��v�U{w>ݙoݞ�����'�R�s�񊳝�C�Q𪪑QT��Ơ�R�����j��[����;Y��ξ�=�љ����`��j-9�q��A�)�����ޒsu�ys����Q�~߯��I�s��h�cy^*X�O=����۞���s�p�����R�*��������Z78k~��`2ڗ��
�+޼?{�6�w���t��/pW�7�϶��V⻽�Nt��˖��
�l�3�z�2(lu����rf
�vM��j�{�6�!�گl�ԧ�6k��;�q����A�W�k���_~N����-y��C[�i����ɴ!v����y�L�u�����������Víw�!��man�o%�s��}�Fm����n��4-�~m�B���ͽ��U��hBu4y}'f�����>ͼ9-��t�h�n��d�i�����֤u߆�f���9����8^z�Tv���1�'0��UWuA��͔wDmL	Z�|=+�i7l����Uڪ�;�ԬzF��o?�z���c�b:�֗�0�f�����N���g�M\q���u�ɴ�?����ļ(bˣ��6��eN͕�zl����q�f��:dt�wq��(vv؜&�,'^�N��C�U���֞�cq����c�2\[F9%�ك��ݥ������3V�53͋��q� �%YUe(+�������m ��ݫ��N�[b�Iӕ�+�����R�R8v0i����;Ó�np����x�i3璾�_2���U�`���y�l�SF�x8A��T���oQ����w/V/Qǜ�]oS蚮+�fv�ӂ�r�m|�}����7�*�z��_x{�l~��ͽ�'I�����|�U^��qr��Jk�	2�R�ۮ��v�+�]�f(�|���3�׼L˱[V
���m ��5'�rQ��qG��
֩���u��r�.Ԫ:�f3*Uʙ1̖��}=;5��n�OE{�F�5m���y[~v����N;|#�r��� 6r�>�[g'>��}G�ܛ@3�i�~&V1G1|޼�=���s/�u!7pE��I����mc��~�����/__������?6�cǉݺ7�Z�|�(u�6�&�3�84^�ŒA�b����5���ͩ�p�<�x>�� �ܶ0�k5|۠غ�0e�Q������O֕]����r�BȪA�ϸ5>.��vMw�63��7�M^(�ɉ������='m�{lٷRnEw�^�o�;P���D��f�/˸sP��� �y��}���G7��6���̷PfV���^���^�w/�Hw �Ϫ}޹��|3�ěsK�!4)�4�J�\��7.5�;��N�:�*�vg-�Q{�UWy������{�Rd�{z{��J�L[��k7>�>��ﻐ٫�S
�8��H�?6��r:�g/m���O �7Q�T������7VGC39m���'~�J�]��";�0tgl�Jۺ���W�3�եPj�p�y+$�U��.��:�
�jỡ�eN����~/���ߊ��n%/�zu������[�7�h<ܴ���Ӑ\D���s%"l�)Y��Jƶ�f��$��޺']y�]���x����ƣ�s�=�y-����G[��qnzym���>U~�B6�A�:���)>�B���k�YR�t�X��Oi�Q�n�t/��c�Z/�����j=�w/˓���nd��/��2h7�����x��^]6yD���j��������mA�0�94���R�+j(F�%�L_NU�Th�<viνYj��rW�Udkf�0j�ͬ�f	Q�F�j�pe}c`稷n�Z��=��r�l%m=�/��DM�H�K�!�#��ٴ�3QSfhF��ݙ`R8e��l�6���d�����:-�pv]�no%��͛��fn��߫��j���&9fY�,��#0\it*��MX��j�����7��-���/��}]~����~Ⱦ�@2�n�Br9���~���e��˹:�7 X�����4��m�}�x�w��2<�ʯ�k�E��m]g���.���x�z����~��^f�d��Y����Y�
�vd����,�u.��m�{%d��ޟ���b�4ܸհ����"��VQ7E]Uڪ7rq�[w�3ٻw=��]�fzs������z��P��nh���,'4�I�;�j+e}�st�Lu��F����NMD��Mud;r�{S�A�5л��F�O�k�j�B{76�s\�M��5��p�j��UR�lqsR�=�mQ}��7�{��߅�j�u����Ch6�g�TNP�t��ӎ_ojz�uSW�GހK	D�#.�tmL\ZWwB�д�IUY�Hݥ�;m�ͷ��9c��Y�B���}�aݹ�O/P�3f��a|fb;�H�O#�߲������UQT�������3���/��6�Z��k���W]V�*����RŇK6j��uD������,�����]��!����W�|rNF����DSU�W��Z�5�Xx�J�\�I���v7Q�O��J}��3;/�P9êP�:\������q���ޝ�"qn��cL��´���B�i�х�ڧ��cDB�ș5e�O�)��/4��sfQ�3dU�i3x+��F���է4��U+q�9}�r�o���9���kq����C�d�\�]���S:-˽�fA��*+�c���^4�����;�wX����p��t�,����q̣DB��x�L�MV�:�+:�+i�\���s�l�H���@�����=Mu]X]��g7�ْ����j�a��`�&
ݻ9�w�=!��lD�TTU�2�U>���私���n�����ђ�[쾭8,��,ɐf��9�F��q�;9��O�Z��*���wK"��R���`�=1����1*��K�U��/lgGH���J��K�Z���5�ڕ���*r%�|?{m�����~�h��)Ip�g�{Z�9�)���R���rP3K;BGy���5ل�l�c�$PB!哒� [e���r� �	�y�C�I^jm�q�����8�r6��DD^ې��2���$���[�,���ҳ��D���/n�w�b6{��$�fIkd'�"t�f�'!���pY[7��D�h�&d�HA�	�}��Oq6���������\�L6�]�c�����������{#�������'������{���{A�I�_~?_|gǐ�ɫ]�0�m�u�]Gr��K+����{ϻ$|�?7�z��&v���l��_�Ͷ�g��[�&)�&��]�����|����=�_a����B�ߖ�7������9�m}Bei���ku���Oq6�����fϤ�v�����3?�z�&E��_�m5.�X����6^�$�%K
3Z�J0�{���a�B�
���,t�"K���]�����3�������vn�����s�Wt)�5�<E]כ=��ߗ����̎ɞ������}<�.�����7N3s�L�7�:i�9�<8[ڞ���_�R�7t3!��%:Wg6d������U*�짽��\��-
�E��[����p9B�I;=��k6��x6������ؖ,���o��v���݇�9^���5'�lb�6Va���V���ȗ�er��Y2�u;���]�W��]a���'�߿VÉ�b3�2�!��4nf���PnpM��k1��~�x��՘���vT�h��q�,�U��h�_#m�2��l]pxP)9��X�*��|�n+�C�p�;v�6���n`���]�˵dydYWM-�0�-���&�̰�nd�s��Q�ѳSFT��n�M������$�Z:�c���{ޫg~�\Ci��;���ƃ�ޒ?��w�����߳"�z�K�e�}*�m�[��ף��v��sw�̶�Ϳ!ne�N��\��h����y�sX���EZ9'��U �m�t�\�V��d�����]�6��w���s܏��a�՚�0cf����SV��]�d����[K��m�xvk��;�s<s���l弞�{վ��j�0gJ��$.�/����٩��cw|ЪO^��]�!���n���*i"'A`���?��j��ʺ�����E�s�5�Xi��R�K�K»#��|i��lf�qޙ^�T��, "��ͼ�T��ά}G�ͩ� ���о\~m6�m�AJn�~����~�9�ӫ�O^����i�n��w.�dŖ�$���LL�E�V�K�J����/�w�uy�}gm�kg����c_.��~�3�ٮ�窝���������{��w؆0��C��{�{B�q������Z�+�|A⓴����(���wf�M�&g~���5\���OȽ����
��]��o��w�9�G�/�e���〙)U�����i�Ѭ3˜C�g%~������R���Ud���7P-��$�	J�(d@A[�n$��Nkv6ʪ�F�.��@m75��p���k�w:�����m:���F�Bj��5ue�����(�}	��3N�>J�z�V�!���ݹ����\mO燽��� #B��%4!�-�!�.���v�f�w gp�+p /P4!�.�<��;��>��@4ím*H4#����?�70�o3��p���dZ	��$�sל]3��FM�LC�
G/:��걪���H@N���Ѽ� ���BV��(hWp#{�؟B60�@Fk}�o���N�7P�t`c
Z� .�	S�@9�v9�c��t�u�����.�3���J���K�0ik�'�I���{�'>��(D�V�@�+� �<���*u�Y�P�Z�j���+ m��0зp�-��hJ�KB56޲jk]�]��hUP���u	3��y�7�}7��i�F$�P
Z�9(D�V�v6k�<�h���s-c�
Bw(� �Bam >:�S��ʪ��Z��� �@|
�1 �hC����)�Wp��l hE��g�r�;�VЇ{�l@]�o�����놳� 3��%L@9��sH�J���p4%w �hC�B hWp&�3��Hf+��{�7�}7��i�F�44�#B9�B$`��� ���Q� :{�r�PUVl~�M!Cyj-��Rfؙ��W���Q�
Zc8'c����N�~BH�-�qCp�u����nS$ӍD���ַ%s���Gt��:1wg�:૮q�Nݺ��qٸ�qᎳ�m����Ƴ�5�ླྀEЍ2J汳�b���c60�6�ǡ[����ԬV���'�v��w�ǋ�\�u����m���_��VWP�)FҸ�m������u���c؀�� �hWp�!��ֹ�N1��ޜ@j�ε���y7 �Ќ�"�|�%4
��-�I]�)hC�uˌf��{�����	Bh�`g]�w��t�u���	SB�hC3�@p���:�\h	���B �p .� ]��^yGn��͕�z��tbK� �hC�% [BT4]��� ]���Ł--k:�D�Y�m\滾�1���N�5��c�RЈ�ֳ�No|�r ��1���
��@w(��\�c��dcG9 y�w���w�θ���,@ugr��wJX[@nʫ�5�΢��D�2�]8�]n� '��B�N�l�UR���І�� �!��wJ�]�N��l���@4í�i�曃H;0k����!���@phJ�G��F�B@�q��|�b�ي����F����}Xe��02�!%X�农d�F��fs'�$!r�<4/�$hCaƀ�[׍�q�x�ޝ@khC`c
Z��������2�da��X�@І4�@p�``��� ��g�����^;����3��.�:І0)�CB�A4+�Z���p4#��o�Q;�;���\hC3D4.� ��Wp��o7͑���z��u���@)hF��;����(E���� ����6�r�.�N9oY�`��*h��k<�c]�ޝ@k�����!Ю�	hC]��f�:��w'Z\�,L�Ę�;*�1u�S ee�tv���Mg$����^Dn��
���� #;�o�;���:�քb]‶ 'P�B�a	H���F�4�����|�Y���_��)�-l9p�������@4�.�*���[Au��z���".�Z:���6؀��KB��%#h�\�
�ޞ�O�T:�;b�����7xּ�gVmj�nI��ٯO���/H��d�fu��cQ|Ϋ�7:�s�����8x@g�xLb��wJ����-�]��3<�A�@-kz�"S��w :��|�n{{�u�*�.�"u�m�V��P� e�0�p4!��@\!4+� Gε`޹��?@�^ F����]Ҿ7��i���Ї�J ���`�w }+u=r��-�T��1�ǙdŖ�f�(TY�)��L�i���І��B��n�-
� ��6��}�ޜ@gM�K�ۇ`k�8ЋhW�Zw	`�(�@��p�oz��0T�B`�э��7z�9ۜww�uu�І���B/0�.��-�5hF�b9�z�VЋhD
� ��awcf�fw�/�2G%���0�\�)�� h)�Wp�.�04#��w}w�-�dhCU�KB�!	H��3�o��j��ޝ@ghCLbKB/|:w���s�Fեf7��d)g��t��3�OC�T���G1dP�b��7�|x�9����O.��o}H��xhX�-cr�-�4!�p
F�;�@� ��_/�=��~�� 6k�}q_;κ����Е4(y�D�+�S@��#�|�}��5Ș|P�ɘ&�ԮeCTf0�+����@s0�	� \`kP�$�!Ю�	hCaw	��9���<�tL:Ќgg{����@��,w 4��!�hPЎk[|�W;q�F�{ KB�m��b���;Ө��BX��Ѝ1w NM��q�j	�����@І�gp
F�]� ���w ���7˪�q��w5��u��A�С4!�d)�]�4!�����.�$hF�Ȏ�@s�)�hD��%�Wp����s͑�|�tL@na%�w���p{vu��m7����g�X2${=��c^���7A��O�5����0����m��6�n�
�DĪ�n��'U��NG)F���
W��k|BI�-b5{��{�2)�/k�euޑ��&�N*�Ӹ�ӻzeH�u�`��r���U�ne��"���4�Q��n�-۵8�q�\<��R���l+�SWH�b���C���pv�i���ym���l�\�ɐ��.�;2;s��5���,�X����{Ԟ]WDJ��JW�+/t���c'Vt��Gp[F4����6�[ZhN����[4�&-Bj�n��¹��:9�j��M)Y��>�WP�ռ�U��[��E��36J���
���B6�����Į6�=�]���O[��R\�Ž���z���Qor�u��i�Os:��z�I���Rl����n]�Xj�䶗�}��ܱH@��;F�ݖn��/�2���}{f��>!���N�����d�/S2�Ԏ��.�w}k�ȴR97Q�Ja;�wg�L��)P�ף��WH�K��S�nM��g5�t��u]����?���~w�H�=X�n�Y����C��e�oo.�^h�;���^ݥm؂@(��pz���<�C���ӂN���;�v�+k޴��Y'yb׷��<�#�̃K(f:;��,�mm��,���ٝi���YZI�6�&n�6��pq'��yu�a{5�
q�gRR�̎\Y��!�Vqg%�u�	yVVU�qBA�Ok&5٥������:��v^gS�=��W9�G%[n��-�Kl���X�U�4������M���v{��xkÀ��ۈ�u�����ij{ON�"j��\�8m����ضz�8�����e�Zh$�X�LՈW�GAճn�&ƓՌ�m�ѣ1���m�ml(,�7b�w+Ӹ��NT��/E.���2�cl�� �����^���v;"`�-��.-tn����d�k�P��\�؀f�
@���p�ZG���9]ڳرϞ�Y��b�7[b��v�$
�+�M��@˨�8�+	��bf��L�7)�6n�͹�wo����\'EDٳ2Xp7�	�
�5#�ܖ˥�B`��*V�g�h"`9C�΋LEu��R����b�����z���:=�X����nv�k��[6�V��u�ݺ���	�=nN�d$��nN�qn��3G],c�9�1� 1��u�����P��[0�|j�"���u��Ph3[�/;��m�u���P���Ua��
��n ����۶*4ݫ�t� ���Q��QZ���B��ܽ��]�knX;9�n�]�du�uk�]���I��.�N�]s� ��	1�m�X&I�4Km�!h��[7X�y�<�nHv�#�ζ�C8�CJ�E)�\�e���`�u��K5�h�Ȋ�2͸d6�ڵ�p�J�]��,W$W�zHءv�0�e ���f�M�Kvw����CuJR��ґ�aIaeMp�tz�s;I�q����=Ŧe��,�]��&B6�
�0tۖq5v�vkt�+�`��nmr���1���vWx���8�p/gf�%���.tVnTu�܇n�M�oR��0\�lrsp������=�(��.cu9��s�k�A��Q	��J���y��W��=�����[�ڎ�P��[+�U�^H�3G.R�^�O*�t'�{�'�դ���.�x�m��޾�d����5�	~�����k�Cz_;sq�M����K��ݸ�=ܰ�j�A�T��UU��NcR����o88@<TEV��l$�؋	�aq���KM��
&bO�I2�!�S��}X���۩����s��>��+�>�B�UT^�!km���K+�u2��n����۝3!�P�2�U��Z���7;��XS�#5���<��Ck���?�z��n:��;�i���q�.�U!U7�绞�pw�vxu!؛m��M���Bb~���߳��_�v��򔧆��4m6�#�]9� Y�6g����ݔ��xݺ·z������p3K�Kv׉.tf�y]��؁,(;7}����D�����	����z;8�"A��8�*��>'X���+V0Ƚ��Sە�F�V�O�t�}�??!�i�قѠ���h�LaTc�J��!-���j"��Ko7y]�����k��we,\��X��� �n79����ݸ��}[U>�����#���#5
��3�wO(o8�n�`�����݆Cm���d�~�o�;]���3/�;X~m��會�˅�F�
:OL{A������ �B��wi]1Z�5�g�ԯl��z�6n��bf,��ju
"�
��`���dL�>������Ju�y����7T��Κ��h6*���ݝ�w�ǼԿham�e��H7l��g��ޛ��]f��^D����o�JB�z�f���I�����5�5�Ɍز�6�Ý���ȅC|��7E����9�:I{W��$�UG��7�m����g^w�!�Q�������:�ˮ�6���3�xS6�IZ��JasE�}�����ӌ���s�m�y���G�n�nm�g��\̢X2�����ٻ+�
 Mm������:��UTUC������uR�y��[ɐ��ߍ�È�俟�=�w��5��e_��dh6�ӿT4�	�v�.��}ӳ��q��wj��ӈgQj��9\�z�y!�ݷ�=��\?]>��e��=R�f��V�s��tMl�4��s�䜓�J[g��L�,�:��-��+B�	Q�������(�o�8�&$uΕu�0A�1�+0;$����ͫ����I�5�3=[��5�u���8������Q�^��-�퇷.�+n�w(�����ا(����
o�n�[�+uJ��6��4�"��6�c��s�/���m��3�ڭ����w�側0��T�D<��I�cq镄nc�S�8��~v���������Sn�o��n�:ou��ݕ�G5|�����«� �w���}�j��ér�v�M�r��n�#��sj��=�>�=��v��~��~m�o�]�}�P�V���5E�X.��K������	)�Lm�V�Q�R����ݷ;{�r�wF�ߙmЧW�t���y�	i;��U
��;z�j��]Y]g
��(�x��ej�':r�N^���ǁ  �g��Y]�O{ꘆ�Wtn#n�jcOB07�۷��5��SS;}U�����ȵ�f:���;�����no{=/f�
#ճ+{4KC�������Wr����of���阆�5���P6m�W����`�v�MkZ����nu�V�<t�Ua����uz��tI��1����F_1ad�v��C�*�=T�;�5�tOGn"��������ݨ�A��[B�z�>$�Bbm������A��y��^�.���K�!�ʅ�G�-�p-	n���ga5�0$��!\����=��篦bϼ/j����:��8�^Ws���(�gsY�yE�z���t+��1�@m�u;a������N�ٺ��Q���
xYQj�oª �qu9q0y�-��d�"TI �R��3�y5K�T�rm�麮��x�}�P�P��w�.����y�����Ud�����ł�B1��m��=�N�!I�{�^��^��sw�5F�5��쬏U/V�d���S�&�L�z�Ȃe��d�̲�5�U���'�('Ft������a�3k��Њ��	e9�������M�m7�����6ݽ��%M��S~����w���Xi��9�f�"�����m�@�J�X7b��+����79f���e��u�&�յi���;�l6�����p���鼌�}Ң�&��Tc�3'�����������D���M�T��U7�^��T�DfƼ���WeK"�fF<�^�^��^��X��d�k�ۊ7C��"�����#���nj�����&�֨��Ka�y��K}W��t��I���*cҩ�~ܩيs4��x\+�az�?��G��$�O~��|k*gn�3͎դ�B�]q��5v�Iٶ��������b862l�˳4l�M,U+�L\�2�ܡ����M��z��j�� 3]�7���sFK�c�x`m�i��v:�7��GZ�l;�C�趒j�.�y}�}t��i��q�Eh��۞�xch̊"S��'P�@
�oj�/{z"�w[�hK}P�ɷA���n[cgj�f����n���ɺ���tq�B��k��(fb�nowAP������
�5��ՓDϕ��g�7c�M��S~��弛]�|��a��[�o�}�{7]z�5T�)�+:���(b��0f�ɸ�yl<�:��3�=J�}���n�V^wt��#�zTz��m��C�k����U�����[�zL	Uz�l�5���^�/ʣv"��v�9�{�}���ֽ����c���4��s9�3�6)�2ꦪ��4>��v߻/fk�}G��g��W(��ѹ'5z�;��1�AP�8tϜQ39�ƛA��leN��7�(ʼ��M�ez�T�
�ꮎ{�HO,���d�DL�"�5���6{&֨�z���u]�"|�َ{z���3]{��e��3e���g�����2Mu���*���5�X4��������^��Ψ*��z��J�;�L�;�l�э���w]}�wk���)@iU�Y�z�D�[ᛕ6:�C+g�Yӎ3����}t$��Y�������73m]��.�\�Ӊ��/��T3wV�����*��
�4^�:Y���/	wҨ÷���ɴ�n6�.�2�����\7�<8s���|�j�w�NXEo@��GFV���SV�cʼ���Z�4OT�d���������%M]e�f�n�uT�|{ ��jk1DU�mU�Y���w���%լ��T��^�;75t�.���9q�˾q��)�$�fͨ��R�f��bre>�6K�������VP�������6`B�D/f옓n[�2]������r����[��*2����K���[Zw��U[8��!6���f�װlCd�ׄ��eK���0Ȯ���xUD�)g�bxxfS�� �3�w}���J�5!��V��2E�9C�`̼���j�U�xVJeUn���
�S��י�<�Tv�|\ʜٗt4��}�P�e��/�ڻ8[���z�姐ε���g�5���
��6CN
YM�Υ:3u�f]�i��c�f��z]��6�W���Ai�'9�Qmb�̒(��[ڲ�2�2�H�y��$�;���T�����㓞ݒ��w{Z�Np�n�r�ryn;�u�/l���I�Gw�EB�S��������)�on��N�#�����:}����o�K���\QG$Gu��
�b}�|�/��$����\ �	x�w��kW��/��x
���!c�z�����^��}�&k�|(�ܮ�H�y����m����o:�#vcv�gz��s�{y��䡵[��އ���vr�M�nj�7]�W_]�,Ң���p3�6��ٷ�Y������e!HQ�UQT��s���>��˞���n�j;�u�Ut����v�UG���jM��P��jz��P��.ZЪm�z�^��χwm�̕�]�Y���O���:��Vr��1a�K-Q����j����f
�:Sb1����h۩�+���/?�S-��g�M�L��_ݿ��u�(�7a��؝�6��Mٳuj��Bn4�7j�Ş�Ƙ�Jc7��ER�S��9m��8��x��+��m�5Vw�g{w�·J��|������7��q�o��u��A��|�}�wy5�Ͻ�f7���Q�y����S���6>;S�~��hu�3���%\���kiV�t�&�6۞�h>���0�|s��<��M��U/Uf��Yݕ�33�]�M��%vl�n��.`;�.�uo��w�z�Q���ƷyEȕUl�߽��x/���R�)D�RD�K�zI��-N�):�Yt��M6��-Z�8�E#�"\Ȭ�p��K�(ʮ���9ơ�\5��7�7$NI��Gomk���䰳�G>>�>�\�v��e�e/'\�u�l���K2�k���ߏ���
���]�K��ݥ��B���ᶀƙ�%�z}����]xg����~�%���\�L�R5�/�g'�ԕs��7��ý}�WA���7Y���{X�����&��'���k���m՜��bd6�˚���ٍ��}��%������Bh6���Q���۸7;�T���\��
"��Wh���(����dX�+�p�L���4���A�UU��@�A��Po��Ez���N����=���F�6�
�V9�q����{~�Ӻ#��Biޓ���CvQ�90����]B�w//��� 
�Ⱦ���~ͩ̚�>Ъ�'��n�W��SZ,�ͱ[��(u| 5�5J�y��X�b�lc���<��y�$����uHUV��}���{�"�����hU!Qs�/8��lB`BD��q&`D�$iVVTa�n�w�<Л����HU/\�����b_GU𙧓����ָ��m�ӕٮ�+f��`�ޚ+�{g�׺���]��
@q��R�*��8]u�W�����os[�y�C�!""dfz�=J �Ia�fUf=yz#&> {��u�i��ec��օR��}ͻ�����U+�83�1����4eԐn�-��[�v	�	�ُEW���Ϻ�u��/��P�?SE����n�͖���Lu�o=�H&f
�sDU*�������u\&�I��܃n�hx&�Mb�/gw�U:���/kTc8̘0wP�@a�R�B�����=��碫���Q}���\ኔ�T�K�˷���u]�f33������q��|�}Wg2�KɌ�	�%[��ՙQqNdL�xx{.�f~�@Qo'~��y��և?w�Us���m�U�ۏ{����a2��iiP[�.ɬ�kXi�cb4�n��N�� ����y���ߠ}�7>�A�_
�vWs�V���*n{����[��8�izx[4sƛu�o��j�uz�� ����V�ww�2�vg^wm�X��؃h2^���k���xz�Vc��h�H�����q�.���w��N�����]*TxǾ�s�f7�*́Z�%�%n�7WC���6�Տ��NU�Ú���	��9'����%�U�m�kM0�0�r�6��C�i��u���a��mǂ��`�����W	��E�^(�*��j!e+�!�7������7�9�%��+�Xzy =��6�+��9�js��Z:�;���!�/�뱌O�a������B�;\&D��(@5@��8T��Θ�\��=��y�]u�y�g�MV���'z�h6�m��sf�Ű`~>���5��~���[u,Cq|��n�lx�[՝ǽ6��̝o�Qת���:�r���T�8s:��9��j��|:�U�'��CY����������U�7��]G��<)��M�v�a����=�}�غٶؖ`&i��4s�D���\��h�=GӞu�:o]�{|;�u�I����|��M��}�]��*zM"�x�����_���a:��vѫ�M���}ƻr!���i��G�{�?
�r_�x��6�j�8@o'���Wyf_�m���h�d�|�������5�������ϰ[Ck��p��o-�p�7;.�+��,5K�K��c\�VN���Z�mN�󅮠US��޻�{�}����`�[��8��ha��)���+�\w��ޫ����{���^r��,K����mմ��ʥV,��Sݯo�7�u�ἃf����߸�/��m[��ڞ#r��c6����V�;1;6�7��3��ht`k�34j��m<�}["��7����>�{�wM�ڿ�^m
"���Tn���-[����[��+���.U��*�=T�T�LB��X�NFnGk�-�tj�N���ՇY�~<��,[>�\Bi�[H���n�28�������7M��۝�ޣ����*<�]
��m�S������7��x/IU�[�}�V6��UHQ�Ug����"�ww����k��+���7�A��=�ރu�|k��Y�S�g�t�9�;��=P����u�Z]���טjWn꽵aj9K1<�CZ�3 ��5'�{»���*����,!�Q7w��O�83��>���-��V���.)X�i]ж���[83��r�뱥>J&���QJ��K��6���\����ꪨ�V���e���ԻVr�[�7�������Zx��1�0���D6݀�b��6���]�zO���m��l�y[��C]l�_��y��V�r�)�U��U<���#�����~k�< ;7�
&�;:�6����D�uu�w���5��Gtr(o#0��Nl�KhےW�d;�)���T[;��RR=��V��#�x5\����*�p�t��y�y��5��T���.M�)ɡa�|�8�/���i��K��U�.�T���q�٨���Sj,{��gt֨��Sz��c{OE`��{�V�H;y��^c5W�k�Z[�"a���nTE�g�S���Ѭ�&s��o�����9s:�r
����kJ��˯\�,�{�x�j�X�9.���7X�s�7ÖN����N��a�*�C�9{�T��L��F��ѐm����˝��܇\h�;�О�W��'tu���v�ǔ���N[�IUq;]ֺ��n,�[�Mֈ�K�(A�7*��ۛ��g7��ZʧF�t�x����[�7jLٓ��L6����u���j����ȼ�����3')��juT�w�*�n�/.�weuaq���r�hud�+�����WQu{��6�-D�� E��+]K����~:�/�� �mĕ��oz�D��Ǿ��.(�+����%���]I��ͱ���u�{W��f�m������y���Ű�iS��c�N�JV�^�vJ^{؎�[-Yy�y�<d��{[���+�#�/+J;�6�.,�J�qw����}�
_k]�$�l�9���N�xR��yig_mw�E}��ٜy��h��;:��xt����fZw��x��n˒���.�:�Nf��Cd��I��yw=����+�{زO�c3�/�B�(�#K#cyll%��Ͼ{1�\�u���L3�O<j��K�,�c1�K��cmQ���9�,�h��ȶ`,�dז��.j
�Jv8LltG;�f�ԙZ�k������y��|�E�j��ƅҲ�p@Z��+ i6jaZIh�V�;�ٱ4t^�r�+�G�j�|.�˶��0im���j�SU�Κi��^�<�ntv��v���k���,@���
)�f p����gd�唱\���7h�ԛb]�o/q��ۙ�t7Oi��\�ʷF�q�W�1��"��=$һYq�.s{�ᅌV�%�<��(i��46.�RM��_\n<�`�^��I�]����!2Ջ���Bmb�Me�іbV���[���)����K�h3�]��{N�NJ@[[��pL6:�(�bҍ����7J��v�p�)�g�o�އ]flܛ��v�s�A���[l<�9v�=aC���l\��Wa	�r�È��4�Fݭ��Bf	F�q5PF�.����&)�8*]�l��ǧ����XCY���!4S�LWYC4u�b�k+M��� S��9ŗ�]���}vG��^�n'�[�d:;b�ݍ��[���l$i��aZ����hAu�	N�J�`mu���C��[��Ɇ��SκrW�8��uv^�v�s��&e��v�N�KP���{�>0|�ˌ.kiڳ4^�ڸI�î�����v�]��9��k�i�pQ��'n�����',ko-�0� $�@�[)��N���s��i��s�T� ��Tm�bX�M��A�Q֖�hdXb��{s��A���;1֮���~����/U�gg��,70`lik�Cm�=YuT(f�̮:�*N1)����|�dң�3�^����;�5ߨ����c�De!�2@���h�l� ��ٽ��U�� �ɣ�T��}R����Q�׺5��:�2�7$�vۜN^亯U*�����9���瓽̸ͻ�ܛA�#F���h�tB��] �c�ǰ��n�:��]bVҪ����_7��}3��9�xw��1[����-�l��}��/��׃��wj�xZ��է�C�w\�l$���}3/5�l	qf�!򛌉Y}��w��� G}5�}�O}ep�+����r�؛�n{`v�H�U�^�8-��sy��=�UDҢF�*A�����U���;}gܞI�Gqc�/	8�n�d6�dU_�Pn�A���}�/9�v��mUsOx�ؐ�I�T"I�"	����ԚC7]�Yy	��.���tC��}���V�^Ve{�C�۠��̽zn������M�����9{��'�k�v�J�Q����b��U7��6��7:��ͻ����X��E	�	�����z	�>w���މ��'tZc���^UUTv:b#cw=��T��*�_o37�=�%!��=-�Ϫ��UT���2C�t�=Ʋ�0�r{���u=��︽�:}#R���b�$��Rn౸�-GI�Qݺ�H
�t�k�U�@{�n;��-�?4%��9�k��}���V��sz���z�X��y2��a9��v�j�o8&��(��T�ik��{��
 �n�=����2����1�tԸ�(h����v�ޤ�m�b�bf��DE�S��ŝ����L�\�߀��=�ڙ��{��h��u���g�����~�M��kw��)Di"(V j��mn3���0�Ҝ�5��Y5m�t}ý�l�o���-�}x�m6�^˺����<P���л�.W�e{�VL�&)��:C��T��qGmEs]<��x���T���(��*v\M����{�<ه}<j鼽A�!�߇�۲���z�E��x]����kG����Z̾��紆Sr��V5�����z�oJR��fވ3X��Ƒ���s��P��bT�N�j��VM�Q�=��.dܵ�=q�#Y�������ٜ�v���a"�����nv�b%��C�b��d먮�H�:�nM����q����/:f�v֮ϳm���M55xD�,��B�Mv�m��ߥ�0ܠf4MMb͜��\���
��F������2B>�=מ�2�Ü�j*{�:�;������J8��k��u�_uTf�w�@6��N#ib�a���I�w�K��5Ü��R�Q�}p�.��Rf�{k��{��̫��FK�[�i���7A��-��gN�|�ǽ��6g�/���_����>�O���kr�:�iZb����b-5�82}����m�{�A�^s�ƞ�F����ߞ���U8Y����%��l���&�Sɿ;�s�p�7űҲ�[�9��r��E�Z����=�9�؇WM[�+��W�==oz_X�Ur�K�}�2����X/����:͙�w&Ch7���|ǻZ��:��A�8u_2��������F�|�y����F������t��W����=�����z,���˔�;�V`��-ic����a��k���x���[����u�3�_Nu��~��У���M�v��}��s�U���[~��ƾ���jV{�i�����IU��c���u=cޖ(��������h�.r�e;a�;�=��v2�n�T�እ~� �{5�zg�yW�
#�������q����U!y���d����o!�x{���ݲM�b�v1���9�-���^����|κͭ��E�5W��[��ep�"�{IVUգt����g��%\~�L�o*��:���z�rm�ͫ�o^�%W���������vL��w�A�+:r�ST��^ꨪ^�-��f-�yw�v�[Mӹ����;���ӝ�L�uq< ��$�;5<���N��;H����iNA����b-�����TGM�����bb������q%�xx5�o�_6�zE�*B=�+��o���.�f{��y���wcc�R]���Dę�f���7�CR���(�}QT�μ�_v����8��p*��w�d6�5>�q�fb��3����&��1+�ykkk�5�i����*u���'ko9�sDUUJ�[���yB�=5�h�׃C��5|J�Y���]wu�j�ͯ�R�F6㬛ޙ��U��~sI#w.��Io�ٙ���(���h��ˬ�b�AU�nWUT���s������5��#�\���a�n����(tAECB�=YX�t�G�79�M���Bӈ����H�&Վ��0��v��	�e���a���M�Fk�5��$Kn�n�a��c3�����kR��\h�.R��ێ�t���l0v�M�_>�^�����Y����0+�i����#�����V�"�U.̛�wd�Vg�hj��K�; +��=v�����kk�g��}�F��WL���G�Ђ�z�]`QY��n�A�k�w Y�����%Q����xi��l��}"D�B��;��X �_<V�
\����o(gyzZ�	�yM�<hA���7j�����Т�p ��:xp���3�3���(G�@Ⱦ�(=X�۷��O��@�R���@Ԛ���@e�Y���c�E����[��>�Y�r��D���<�8b��m_e٢�kW��D]ǠnЂ �}��R��2��5���κ9̝ˣw�����q�jfK�"p���(��`��k�� ���/G���E��s�ګ��q����+TW�!���8~�}"�a�ܻwW�˽�����}x�<B2/�J6п:���P>^"�x�-�����L�E�As��e}�B	҈���@Ⱦ��sl*��j��y;Up3�&Z���Z^7q�|_1x:у0�ȑ2eI(�HI�ʘ�Pv��v�-�3�x��A�=v�|l��9����S�1�Цf��4� �dT2P�"_H����o:(,���/;���O
xi�|A6Qr��{v��W!(�ڠA����ED+��{"Dk�O��v�g��e�w2�0�t{ĳ:cO�}n��\ ]�Su�>�ʏOu>����#w��)s=H�'1l}g6Qݜ�p̷����m��WUޢ�vS�Y�	����s�<��:n�c9���wT%;�-��o��%I�{f�oM�O�jW:��-F�톷�a���].�^nuJ�7D���>�������ܫ���r��jˇ+����Wq�<�å��i��8�6v�����7S�̕��U��l�WyO!��Z�h)+��Ƃ���p�H��t��y�Y���Rp[�x�� �G�-��F��V�;�a�$eQ=a)�����b!�N�����[2�3\	g�9���;]/&�I��Zb�^c��(�8s��-�L]��Z/7�2Ňlo&�$*$�F��2ﯲ�n�.�ʬ��uM�3J΢���:� M�X���[N�e�y.p��۸nl�t0\���J��cҴ�;+����C7R޻��5����k�ט5�s�pj�;~�ۢ6�]�.�5L���6BAbH0�!I^�Y5��bǶۯw�Z��ד�y�[�����/||�|�۲o[wa��O*��n �k�B��-�BYd�Bģ7�ݯ,�.{��>�B�z�-XK�8Y�X����m�Lp[	l�"l𬱼B��Z�������c��d�#�;/ ����z=�{ͭs�e�ی���܊9�1�'��c�N�a�'
<d8�r�-����٬�Y�LS l%�6<��[%�@	eC��)2��׬����M����)��Qk�XM�X}�V�{��$yYjG�m���S��		jE��A#-�!N�/��1+���z�޶m�<��{׻��ф��d��Hڴ`+�D�),�[G�k�f���=�z�;�Ͷ����E/���{���?���F�\� �PA�(����B���s�Yl� �P��z���h-�����8�x�Z�Gy�Z�!_FE_\�!����r�+��:pO��	��#r��20�����S=tw{��.�ڄ�Zl2�T؛K2�7V6�an#�/�� ��QIB��qo{�Y��G�'λ/o2�%d<@K�$�@���"��1B�R��-8�;���� ���8�n�o�����dq�/�IB�/��##����K�O�^��l��
 Ȩ�
 ��s�.`7�H �^�^�w9NY���up3���V�G�P��^jZ2���y;.u�٢�2h����Y�B<��;�\��ݶ��bk��+/w>��3����"��?H��"��Y~����������� �ڀA����}8o~��τ�q�%��њ݋eV��ap�4ɜ]�����/?v�D�IB�u<����L.׈�<����wP�"J�L�=���u�����(� �9g�w,۫��ѫ�#?t�W׹B��U��d��L�l�b����f`彬E`�C��@qڠAP�!;��_F���/��+���힞
a��A�"
�v؇uQ�%P&DE�+*�wn�A��w{�ͺ���ס�r�E�+/�\��2{�h%��+��ME�o����S�ms��j����݃�����U�_��G���k�aᶹм�&����8瀞���:�KfY����þ:�?9Z�c!h��ݯ;�,%X�St���]�b���ٷ��[�y&�8�Bn@�l6km�jM�B{%1�<N�%�-��a�=���2�v��`�ۚ�m�}�>�F��T5�LRU�q7XpR`ME�w�����}���h8�^O7�V��r��Y���B9�7p�&�A9|���\���Z�')�>įR��>C2=v�T�������ܪ�"̊�J���3|�f�[�7#8 A��^�+��� �LN	i�:�B�Э���*{�%`�C��FŪ��!���Ȩ��B�	�Q #��G͹��ko����^�%xs A�Q�-���g~����jJU~"�gc&y^�8��i8on.�mGY���mdH7jhG�FY���v.�a��{1�$��h��$�FD6��u��/K�ju/'7�){��v��2fn���x [O>�h�҄"�q�2�ʰ���&�uA�6:wu\o|-`�����X2$'�X��[@m��b�$@C�nL#����~�S5�	���^�@Y�U����:: �}\��%
�!�{��jK�	|�of��Z��N�FE���dP6Gu?��%�G]��9�@��Q�/�������W�(�psM5�I�nu.+����q��.��}������#�Z����*����xb�Qg��~4p��P=ʈ&��"�/]G".���H|����yn����.���}[;u�|�o���w/P8}v�v���fS���G���uA��A�q�[�V+�t�V+��ۛ�؉�����q�3�x7�Q~���d�}�k�~x�"���c��R���5/]����/���W�)q�O��s֞�k�����D�+��A|dR�eU^�&F�@ҷ9s�[�9#9���DD�2P�kw4j�FȪ�b�ރ	�k\�ơ�r4*s�UJ�յ��Qe}"g�P��f���X��J�hB�TA��"^�PA{|� ����܆�ݷ��j��. �(Fdz�+�l.6e����DAC�2/�Y����ۮ���o�3��!�D,�"��yPܣ��׬�坵��}��	�	�B<Dx�>��5��F�Y1D^�V�U�g��J�v��7<�����v��LI�彊�4>�G�#� \�A�PE���ϧ}��_t��c�����@Q��P2/�»<|:<��ҳr����r�ڟ,nw.�c�L-��|'���gם�s����2�|�n�d��!��2U��*�A}v�v�fϧs詽�Qܽ2�Ae<��ٷ����P �B��#"�7C����H�ED2!��?7B��9���ffg�=O5���A̯�O�0�"��"�:Ґ�F��軁�/S�s��H�������ݗ�!D3��=v��l���lU�-A���_*��:��`���B���E��Cv��F�m_zLS����S
{2ovfV3*&^f�X��FWW4�ڬ���i��J������z��x�.���fb�8\��k��Bƻ:,{mn��pk�;GDܗ'E���2p��xJ��E">t�/���'D=:Kf�t�e�O5�k�c� ��3�`D�xܝ�W��XzŻy��%��\�P��x0ܙlu�ͦ��z{�"i�-,��R^�W��oN�e⶝6+���}>(W .|��ص��8ۚ���b�k��0x�|wU�@�(P ȅ��݌R0�V��-��s:�H�8�/�v��b�������m2�
H�~J��+kɷ��hx���PA��"��ر/cp �>Wp!�����v��. �(�يp�f���A0�D�@��!~Y�����&'P³�Gi�vrp@��翉;���i���ejG�hk�x��4;Z�r�7h��L�>B�7k�l��.�ocx&�@;�#�S���� ��j��v&E���v�уel�X}+�u==�ԃ��li}�n��U���j]!K�sj��X�����}�^s����^?Y_s+�/��E�0ΔF�
�bD?H�D�5z�n�³��o�·(a��x{h~����ó�r �.�@>���=Y��;��Hp7�Zת����TF�ZȨ"��n��>;����s�;����i�\A���}�B��Q�Xg�!�I�A�E�F#Ŷ<�ô\!eх]]�uV��B�QE��!^U�����Y�DƹYuU���� �/]� Ȩ��摥���TAJ����Y�0[C�G��<	��Ǝ���j�B����{|L��g��kY�]4[��\�ʠ��E0��ɍ�(Z�[w;��g�Es��S}�����v�~��9���aDI_P���}ۻ("M5軁�&��m�Wa���Az�4�#�a|@��""E􋢆�֬j6g-��h�	��A�B�dTD�nn�/o+<�.愨Z(�_S�Ֆ�$�;j���{THR�&pg Mj�A�����ϝ���1K�g+�M�(��j&�]�nЂ3���<Z+��@ �@��&��S���0�� Z�L yp׾D{Z�,��nנ��WN��msû�扮�gP׮Ԃ.Ђ,�����^�7 @j�񻁯':_<{Ui���6g�̀ʗ�>LҖ�]�䝼�5��jUX�gU�j:�nF=��VtΎ�sP�f�A҈����D!]�s�!��W:�U8��(aa�@�<E�+��l��}��{�ٮq��2�%-�!��ɶkTt�x�F��O/;�ݐ �ev9������\ 3�5�V]y	� �E�0D!�*Z��)/��q��ǵ1�)q�J��A�y�J"6= �� �!v�p#Kr�r����aC9z�����7j���>�p ���͌��y�4��'��*������v��]�^겠O�v�;ӝ��f4�.�P �@�v�̀�2�;)\�=]�ML��ct��Q[��s �����Gu���m�V�ՙWU2�N{x��>q�,Ō�Tb�:�EUI#WMb��{�s�Jḁs�O�LT��뱱]Ng�8�5ҋ�5I�41W�oY�Y�����8m�5�#�X2�L��g�l������p+Y���r�����[q��ô��Wd������"�.����Rs�2����1cV	?tڥ�h�^L�����'�=��W��m�36�����oכ�b��Ц��=ܸ��wF��Ɵ9LŹ,����90U]e�E�t+(�}���c���&�*�N��*�%��k�r��]���V���P�b��Ž�'��%ի�Sv�VE�GU�q����Y�I]'�k��r��wL0�����s����r�ϥ�Lw`���b�Q��N�����=r��'�#%P=7s��q��i*����e���f�l�*v+Eά8�dU�Wc���CTɱZd�عi9*n^�M�U0Gb�李[�� �u�8V���An��M�s���[��r�����,�|��$��E�c�n�8�me���j����lH/x�E9{6���V�Y=�֢VZ��5�_=�[v����Kﵗ��ͱ�7�m��ַ"�̓��|���R�l-��"M�gg�S͚C0�v�v�"miY��3��2Ͳֵ�{�Ś�ז[i������M���׵�km�$B�^��v�Y����ktm�4�-AY�u�'�q�D��M��Ύ�ե����ޓ��9N$D���-�Ό�Yi����^y��Bw��B���F7��R��8����������܏W�g#�'[���6;!x��A�u/:q<�Z��.<s�l�y�K�	s�8���`M��v�Q����m��ӵ��t��=��^sě֬�F���s�#�'�ex�G5�:<��@��d�.��q<Ru%�.���.����3
�L8�h��M�r9'�M�r�N���l&�i&�͞(�Ҙٗ,6mH˦kqD����L���e�nC�g
jV��t�	�cgN�e�^�G��^�mz�"x�zc9i�� ��q)-�.-rB� �Eβ�k�%Z�N]��#p3���u���@]r���э�y����s��؆ظ;6֚�v�����z����xɇq �M�b7J/[�.+���Hncq��d.Е��� a�q=ȝ��6�m;��z�+]�]����PvyN\g�)y��q�1�P%��
X�6�6;Gb5�zK��K&�Nu��ʺ���*����1�	t��/E�6�g�,f1��7:��E��6A��y�k��Eİ7b�%�ɇ�+���b�6\��6��L��оm;d�vu�n�v(��a��=uq�6�FⵌY��C�Ym�V+^���vv�����ʷa�鮰�K�4r��6���]<��ـ�"�C�]��因�q�a�K��<f�˕�0��C�S��;h�Gh/e@�5ϵ#�,Z丙8��46Wd�pj�϶qID�R��pb���iI�	�ZP�<MBSY�*;x㎧����c[s�.�v����i6a�~��~M�U����'���/�F$v���>�e��/�/}�{��y6�U8��(ak*rg�z�9^�p#�x�"d@C������Ɲ���gV<�=�G4[�oP~�`��/)������TD�Q/�����V�,�{ێ6cL��ID��TA6Qp 0��L	�G� ��r�Ap8�^�UlN{
�5��^]ǘP�j��B����¾"E��w=u2�,4*����{��~�A�@qdTA����7�S�"jKB[���՚�*�C��nL��7��Ά���N��Ǔ�8��l���S��s,� �ǫP����2!@���g���6�^��s���%0�]\�v���;^�{U�����٪(Q�ZI�;�<E@��r-��؜�(Y����m���zV��:�
 �������盻l_p9�߅}|�|A����B/a`��#�R�M!��v�we=�}�3�iq��9�N���ّ��ϰ��`v�x�!v����_+����N_/�>0׫���J���z�Y�N�ٳJ�at`h��i�25լ�ɕ10�B��^`�D��ڣ�+���2�K3D��D�P�C!���x�>�RB�.\�u���)�h@�۴�llN��2P �����:+o����	�
 ���?IC���?��S-�x5��`�-�`:����,��j�8l׸-��.�!���\v��v����kbr�B�a�F�E��w���µ�s�fV�4A�����0�)�w���&��	������6�Vvp���?9B��#"���DB:�n]��^Ї�\����S���;�#��z���wם�;��֦4�&�Z�3Kp�͆T8&6�����D_H��$��*{���x!<�W����O��!@�K���(L+�ؽ\�j �C�^�^�+�h���@2'��ut$�t�>��@"�E� �%
"/�� [�N����s�9�7�����Q�@7j<}g�s��=����� �w����f��|�zc}6�aӵ\rJ�}N�@̗�o7kLӖM�:�
�.r�2�w>j3�d��C�i��]0��rd_Q�$_H�b�Wu>��\�h���@qdT��^u����gJ������.�AXA��1��dv�;����ǿ�!�D=��c�9�������}[B�j��*�2!DW���.wU^PÑ}�=�{q!|>0נk�_gvl����P}g�k�k�l���b;7�F�w^fF���E!�ZA�Av�n�A�|����(����sμ�l��5K�d��tF.l0j�3��!� dF�1UW���'B���uO3=���嫈:�A��n���Ġ���]�k�����Oڏ��yw���;8ʩ2��>�;z�;��YH�l�g�?7��햁t��&�r��W#�t豳�sF��j	-�nɹϊ��\v�����)�Yx�mQ�\ob�ˎ�gaY�s�mk��6866jq�øw�8ݘ(�P�'����(El6Lf��V�i��0ڴ9�����tܵ#a��w=�~��8h���J�]Sh�ٱ]�5��v�N}/w�>�ڃ�)�{��:α�;T�Z@w �wx�w \�A�P}'�:=+�>�w@ד״���5K��@���V���26W�m/P��ڀA���b��=����g�$/���8�x���n׵��]�q�r���}g�v��CgX������u�{�kTd
B2*"D>z_fe����}/�_i��[^?Y�bdT~���Be�7��1�k�J(�v55�Ҳ�SD�k���{���썞�K�g�У�7�g��x��'��YqP���� �~�|G�7D-~��ǇAN�f��뫮�}y�f�7��8Y9Q��7�g�\�n6mOmظ���/w5cgX�� �� �BE�>cu��ޠ��}%�$�����y��t��-�	���,c���HN��oF�X�Fm�=�HƮ�@/&ۙ��$0�j�*��3bH��whQ�P?B�2W�*��O�����3xz�X����/�VD�N��[�C,�!y�V1�@�k��9nŵV��%bf�gi��<�yg^坋��p#U���pٳT��;�2�F!�k��]�]�u5#�b8�=�-���6�xG<Haa�#ZE�D:E�g�����"D(Ȁ� ���^��g �s`FdT�7:s2���.
d��n{϶�d�푗ΡYy8�Uĺ�����NQ����α����v��w�뎎�j��4�}wnU��x�lٚ^�d��&�.�3;�5��a@�*��QdI篱l�љ�1���7��S|�r�5 �� ��}�k��K=Tm]RUTH�(��ծ��:�h��R�b��{(>�^�\��������b3�[��$���կ]�DY�ڒ ������1�x��=��i��3I�L� ӄu��������f�D��PA�����>�cWnN�''�e��a�cB������j�n�\�A���͟v�z�Q+ܫwp��ֵ�΀|n!_(��W�؇a¹��Y����rOmC�Q�m�gQ�6�c�ep���I�W�D�ܡ}c��CsG�b�D�(FEDH� ;�~�]C3m淜<6����g�:W�&Б�~���ߥ3N��4�&�ZA.�-J:�QZ��my��2��B<A�� ����%�r����2���2�� �/��� � ��e1������f�S��G;�k� �q\�E�;t��(�}����?X��+{��yo8xmCq}�l��}"�D�(z����V<�@Qu�]�C�`��¶H��׊s[$�A|\��LA�"�E���z~�b����5���A�B>k�k����.\�K	ѥ�{{�.,�-�v��{�����l�)�B;:,1�A�٫�j��TQ�I�I�)}�G��<���똝n��%P��Q�c�I�Y=l�&q��S��7�;����E��y��'Oa��t�bv���P�]���[E�M��B�ZC �\XD�c��[���1-9*�����[P���m��}}�����hH���ღi��u)�u6H���M{�
�}v���*���6ḼGi{Fj~�B�b��?ItD(�Эq=zn�Df!�Ou�}G`��	���
"�P�rzQW���}_?H��"��>���a\��^�{_V�����B2* �(	hOH���R�0���윶8lٛ^�%-��w�gG�ND�+��A�7�����C
�\��b�^����h	k�%|m�c�<���F��vU���p�غ���Q��Q�&�+��?z/�\ x��</��[���oM��Z�F/���I@B,Ȩ���R��f�3��:U�e�Y����t���)���=}�v;�f밦x��������^��<6�@A��n�����3�>u"8�}q}>��/ʖn��	��-���y�Hi�j��~����a�G��B��PA��[��=;ѬU��fЏEn4X���͡DB2/�J��J��8�@[۫�{|8lћ^�%]��v6[����ױ�t�o�b�Mu�8�E�#�#�c��Ń�"I%F{��B��z@���`�c)�p�7�!S���y�sh��Q�W�aDO�OV�z��t�svx]{|���8͡ ����:46J��ԃ#�@���(�>B������+|�3��5����������<�ɔ#,H�8-�[wX��M��h�/�+��P�j
��;&�+q�y3�dƸo��23^Ѫ΋]IYx��}��R[{�&d-{�oa�m0�7blA�*4�	Y���6foV�r*,K�\����:AI5G
��ُ/K{R�pj���T�-��0"��Z2�N����JD�;5�Uٴuۨ�ణ�y�i�b-V�%Ci�c&��m�D��Ӝ�;�V����X02�����zz��
.C*�g�(�qcIɜS�;B0�W���>ں���5�Q�C,�ۡ4�+i��Av_'���΋o��[:hiՇ�ݗg���ѵ6���[�;��mr7�}{8S��ԩ4�\ti]e�]�����g^=H*������樽quEK�=��e�w��V�Vv|��ɻܤ������蔙�$m<;���ں���,�捇��ޥ(�ی�r�{Ԓ�Wt��+r�w*;��$���d:w��J0��&S4M�u����sq��̺��<\���$+�J_"�F���6:�m�n۵��f�gC%�6�f�l�ۗ�$9��/kl�7�g`�ƙ^u���Ժ��{��ݭ�{i�f7����Nr���-���m�P��99F��m�۱f��2�ݓ�'I��,ݽ�w��S�H��$E[X^^��N���q=��k;-�r�e۝�Y�N�D����5mbf��/lFXs� �[�{�6��f�C���Pyyy�DrP�m������`{K�$@K�Q���1�Fq|}'��z�z��$�\M�[�z�HiB=ʁH�0^��s�%�AX��è�~qED�(�%
2 ��"�#e	Sy���o-b���hA�ڀE�=��Ϲ��O><�vZ�;�9�jl8&a*�-6ab!���]���5D�P�"�%
��+ۼ3�m����ۛGe��
9ʁQ/�B��3>��(�(�oqy�P�^����-ㇹ�D5>���Ң8W�H�0�e{�L��x]�Z�*�=6�A���94�!z�4�E�o(��c8lѭ@A�.���Ӫ�b�R�f˻ЙL{���ţF�<���:�B�E�k�P�T��Y��G ���n޸+�x�/���K�A�
^�B;;���Ӂ �s�{�"��\���e�%�G:$ר+6B@����81�IM0Jd2�E��)S�_a� ��FE@�+�NdlL���*�)�էa�E��q�z��(���*qG]�uZy``�? ��yF�u��F�{��'q�ץ*�f���r�B�1dU�JOv�n�;���X󂁼�z-��E��v��݋�D�w`A�PA6V)��b'���v��
ˑZ��0i����2* ��E�6Wm緺�I���v(֯q��=+� �a�6�����/��̍�	�ۧ{9�,ݝ3NSٖ��'ZS"�g�2���c��(�H���P�d)��N^$�nm1l���ɝCGGG[���si���ֲ���ciLY�GM11��9�7<�͸�Q�����B]H��ml�[7L�����%�=4�-�*km����0�m��rv^x���6��Ҝlt����=ao������˸j�G\����2:�ku�#w�$e��)��G��|���� �
�D/n!��K������!�
S�N߶�i�W�؉��]��m�7kp�8!���Ӂ2�PE�E��.�kۜX�/}���j�	����e.�=/��(mAk�w���d<�o A���$�P:�7B�D(�@��/u×�D�4V.˼����w�3hG�#�#"�A��6�6Eo��M���T�<.���Nѳ֎��aJ�D�͆׫W�� A|��gF
z���kWv��9�v��:�Mz���
2!DK���[�3�����1�䢧d�:3f�ov'Y�m�[ڊtПw3&�{��I�B�1%>#����oG���ld��o	�� <�_x������8P �%
2/�^n`ٞF^��\�
��[�D<n!D ��P �(Q�}�O�rw* �P����<cy�;k�����b[TA0�%�&D(b�E�8�X=pp ��ǌd�pR7�&��E��wCgc��!�u	�7F��+�
��=z淊���R0�(V�T�͟,��ڠ}e����'���v���)�:��h#�Ah� A�^�.���aRd@"�^5�9v�z���v׸�D��ؖ��C�^'�9��#�@Ⱦ���J'�[�d�9�L�H�b��>:	vf�[џV�d�1�+�-J�խ��"�Mn��)G�NB��/�_H�k��˽�4�A���/Q���o/����]�n����Gb���E�dTAP�&n'�R����;�������% F�n�Y��:f�}ջ]��cJ�T��:Z�JR ˡ�3\��>G�Yo_>��2/�Jv�l��<*ƑG�|�r���J�E�K�<���^ʔ�PA<W)��f';��w��� ��s��㞘�`���1 OZ��E�+��L�!�VkX��E��'۫�jϡDITߎ#��m sU����Ꮃ�H�勁n�'K��K�9F�s���.�{�����N�0�{�a�M�ag��H�gW,�c��S#^|�v�M�!w�cpLc��qG.wt�gq�z�1�+������ƽ��w�{��~ٻj�f&��X�&a*(J;!-]��]����і�x�K��{�ޱ͸�9k�{�\׎A��0z* ��]dB��z�iq׆�Ŗ�s#�0mc�8D���1���2$¹�d�۫�AP�"����FW	�s3�#;��x��rD���6�t�yrV���P�1/���cy�n�ID)ń��Τ8�_WǊ ��"1dW��T����C��[�
F�@���h��.�\C�uҦ���b�YUZ���`��T�rܪդ� ��]8]-�
WӨ��o�gP�]\UDy)���PIC<�@&��ŌaJ]�ͺ���	`�,om�mN��sa�1�ే���X��d�[±y��V�q n�nv��:��Y�8ͫͺդ^�{]cQz�<��hj��O�9�/'V����I5ty������B��1f�ٲ
�Wb̺�.�\|�SBڀA6rU�k���-�΁�̽B<�ڐA��,�7j3��u\�a�5/n�wu�l��*���2W��B����l-���#v��
 ���YIC2�T�X�2t�V4��qr���{�E��HMI2-ǛTA6W�b�9�F>���8qA�瘾94�q��ޤ.���Sܒ2���� ]O�p�|�v��J ������^�<�?0��M-ܸ�"Z@u�/��d��n����������D�(����P7�������b��� �K�����}�Fk���*{��d�c1^]�y�f���oa���x:C�	!u0�uF�F����@��~�^��1y�"-���G���8�n�����ŀ�2W��]�^"�^7p$/^��5�^���<�q5N=jI�)v��)+�f�9��� ��PAp ���c�
�@�j�򎉈�/��p ݨ �P"D(ȧP]��:/i��T����qƅ|�E_d���5U����֠8�5vn�ˣr�c+`��]���<��F���c�g`^7p!gk8����9k��5��xe�?'B�b�	�	m ��rUC��Yr�M;8/s��
�-^�{��{���PA<P"�z�P>�	�p�����7 ��Y��B���ee}u蔢Qp�霃&�G;����+��P�=�S��lf!�)qݨ �B��oڭ�mi�5���3����G"� �({�ݧ*1j�¾"J��B�辑y����ѯ:�:�o/CP#\"ϗ��N�O��:�s&�(�]������V�j��UnC?�?K���2�PA �fb�F:�f!]
DNZ1���IL��w3���Mև�S =^��,�g��5-p �>�BL����B��_6�{P�D!E�GV>�L]����&�5� iz�z�P"69W
���H�Gt{yP�W)����α����v�i�{}1'�^�Z	���p��Y(1�;���/Fǫ	�]��jN��z�/UF�
"$2* �B��w�!���u	S��4[|�����%x����ڠA0�םZ��kt~]�V��wE/G0�����a����K6!�z������ܚ��3g���Bb�]�(� �� g�w�T}e ����l�ahf�z*o7�c�x�gG���A�ȯh�g.ۡ_��j��
"��a��.Me,������;K�d����>���3z&P��j@"�;�n�X�<#�a���~��Q��k� �aD(Q�Vf��9u<SP�Q����	�B#�@�@��_�{r���E�=����̆hv���RJ�f2{�nC����
��xE��B��
��<�7�8�;�����i$6T5��묪�Q��Y�����yfk��iv���S6 �˫���M���rV-�8L9�;5�^��ndf�J�O.�	�j%ժ���	I��H-#��jām�F��M؎��cY��$�Q���&*���Z�`xe�+�����=q���Ǳx��I�P�us&6�)�l$E�.����,��t'NbZ�*�k��T�YT��L��g|�I��P{ٲ��{�Q�����V�rT��I��b��$n*7cie�۩8�67J���U��jŵ�]�3^R�^��7�@|��e;iJ*f�L�fc�tצ��~Wb�^k��7�HP3%Δ��[��r�HF�� �z��V5���d��]��*W0�iuF��.u��f����L�Ɏ�켧��h#̓�LM�k��W�
וVc������	0^��Ԃ�g��h������Hn�x���������$��y�b�Nmb:I�cggj�Έ���Y��jdP$m�����m$N��e��Y�	nKn���NQ9 �Y�oo+1�س8<Оɧ	�)�X��3��y肏&�[g[{ݜ�³<��{g)�Q�=����ę6rI���K�Y��b�(��t�m���;���y��B�D���M����[�奘6�K٫w��ik,�Ym�q �%�I�RH�֬M��c�dg�{�(���æܶ�c7Y͖�"�V�^v/1^tj{�W�ۛl�Q�k��"RNI������Z��J��lks̫M��hh�/9����ݣ�Ϟ��Yͮmwf��x�uׁqӻZ*հ<u���k���Ӑ�#�T�Y�W,�9{�<�h� ��}n�uAn,��5��+��ѱ�T��GQ���Bt+��;3�ה�ᝆ�����$qY-�U�Ͱ=3G�m�rMV+b����i����][�=��>B�z��ę,3���}c��S��<�F�.����S�rVsԶ�*�-�b>G�P�#�Wz�67.۷��їb�k+<�_+�BV�f^6��������w!˥�ڂ�ؔ�\I�OX���<�#h�� OF���]I����6��!e5X�сx�kE�&�5�&�ʢtԮnv�I��I�C���y�Y�-����Od�X�+�q�mg]�CU�vpM.�¢R�AKK�����J�B	��#� \���d�k5el-Ȩ�#�tv�]�'��8z��ϓ�4�Ŝ(��8L
�p�y��SM�mƎ�Oq�h5q�Å��Sk��v�G=pq	p��o�E������0����]<:���{qc�ي��j�@����͵��5�Ǝ��<n�#�Zh�%�}�>��`jB>,s�dݞ��2��ڗ^��K�-�.�qꨢ�t\��v��;O^�.��[e�z�cTgW�my�I��nZ���jNpUb����H8�\�hKov�!+1��LT
�{0Ź�sίY3��v�N{Mˁ!rZm�x�\î�O,�h�^�mGG]�1�]`�L�/5tO{OO��6-�]�L�m�7]�[���]s����C��<蓮���/wCyi�-A�^W�*2�� �A�Y_@��FI[�(�/k�����xD�/A�̀+�"H�����7�24�T�&����W@��so�T=�y�8/\�8���U "���bUA�A݁a�7�x������.>����Ԣ^Ϧ� �P!�� ��h/�3
:�x��_�^У5��|=��T7�/���hk�����)҇��ݝ�5����'�u��˕�3h���s�_�嗢���[�%�Of�ӽ�3���h��ug�<��et"�(�rb�[�������{X����A�K�j����y���n1
�o& mT�,�k6�0�@��#�P�o�N.�Z����6��1z�vwH�	��Ȓ���h;�3�I]*�m�h�g�zO�́]ǣ��F�G��s�ZΖ2�� ��ת|A�P2b��q;�y��r��j"/�ϴ�cZԅ�F;j.䑗|�sZ�T3D���O��){����#v��n�w@���Ҵ�[qe�)B�Ґ+�2X��k�}�-��#׬�eE�=�]��{"�
'7�VY�A�B�!�
����&EDI׹۟b��K^Ә��Wk��w�0�7(A�=dl��&쫯p���P!�
�� $��#̇V*�?fJ��y�][�7&R�LOQ��ޔ�42�6]d�z'n�
�[��LS;�����(#^7k���h+�z��A͡G
 �B��g�7���6zO�+76g:^i�1�G������E@��_H���(�(�*����]��&� ��l����M|�y�����e��ZU�й�c	s&"�Sp�og}��{�;���6������(9K�X��s�WF�YB|�����/�B��x܌��Аs(���{�b�G��́]�2��3��wW���Aݭ�6V���_���q�ޓ4o��Т=��d�w���AhD�@!��A�|c��n��3K�z\l������*����qfUvŁڕ�<Z�;sc)­21���f�gC��������o���"�@��]��e�G	�� ۣ�ùʈ= �%x���G}�y{%��������+?LG4�Υ�5��BgH��Hm����	��I�M�|׮�jÚ��;�{�H�c+�زbA�B���!@�*�6Q<��mV���hk��;��Aƀ�^#FD{Eh7h@oU4����}w��w �g����*4�X�t��@&J�E�G��nףc3�֐e^� �ݨ��;�{�H�nP�(��$�{�(fP:���P�D��ˣtf�ڇs�c��7
R%w�#F�v�;zWv^�,��bC��������*�&\� ]��vt�Olm��rL$ĝ9O��b�ELȉ��э@�������kklGiX�@�]L����j�S�)Ќ�n�E���kRf�L"f�L��%9E�XFl�J��
$��{���E�t,����y���G�[;*��^��hd��'
g��Wm�����m+5���X��Qf�Ĵ(�t8�ɘ3TX�ӨAn=fAkْ]l���"��-^��>�@k���7k�nעr�m��˖��k�z4�7(��:WsZ�%Z�B�� ��"�U}t{'o��5���Tq�M�@��#"���!y���L��"�6Q��Gm��Φ l���@�����w@_/�j�E����)�~���:�]O6v7�ލ#��@w/Y������O��|�b:5�;%��SKֶ �D�G]6tM����}�x�:����Av��3��p��/ZO9��9+A�x�n�h M���j��u�7�uɻ��u�^�u��y\�le��IGJ� ��ȣ�.��y�^�ǲ��>]��`l�zJ �{� ��<��#<v���B7h�sN#	��LC�➷oF�T ;�
�
"J�tY���@�?01�*=d-���i}��,���iAvsE����* �{U_H��+���}&�l�{�M��t㚨= �'�װ ��^wgZ}��h���,���(`-\��8'>�Y�r�y��]��SQ�A��׮ԐA�Q������F�xc��M@��wq �>�Nl�"�ݏG���w�-�*��V�F��S���DX4���sPk�}T�-sO1���!��vUb���R�׸s�~��o�\۝��������؍�D�[�7�n޹Φ�m�P&��m"����Y��w�&f���v��n�w_e�������(@!NeD���L���@��v�g��w2�k�l8�#]v:��R��ڢ/�W����~ǪΨ��Cr�腢Q)���������k��<�<쌲����Y�p ���w�q�����Vm���n�W� �2* ����۳쵀�sT���Ҟ�[c9jP�8l�Ge܃Av) 5����+�$���f�7��mh����]�WK��T bݨv�i����~���+��d��;�M������Yr��kw"�!=�t;�jB�N���a�Ȭ]`\*�t��:4D50.��JK���z�@Ⱦ�"�_H���]^M�A��+�ܬq��60�5(AvǬ�n�E�=���~��	rʹ�8���M3�Lɍ^1�l�{;쟯t���;��#;��e8�jae/mT��ʵ����~2*"$�D(��J�0�D� ���w�^�܍�8(�� ]�U�GO�h#���1}�"�����xQ5�i���ޭc���v/Y�.ЀE�G�Ky�c��`�'�@"�#�B|���p���8���/ntZ�ʲ,��M5�"|n������q���A�o��^�ݍ�<l���
"J���?�Ý��:H���=|�{hڷ.���8��w7�s����4���B�f,�M��V3����޻�>[�jU���91q��[��f�'���<g��؋�&��U�g�n}l�v�,p'[Om睢T�:�:㧎�+��]�ӹ�b��"��y�6��-�18��o< �i�&��٬4#4(3.�ۿ|���b37`f �j�³mcR�H��5hE�nϝYo~��~��RA7j<�<��V���?/�f�|�A5G���]�#�d�q���+7+D!����ny���\}4�W��L �G�a^H�0r���]�2�r���O���j卿P&���6�%W�/�_9�vZ�F* ��j|A�]���y�{��v�#[�\y���B���e��.��~r�e�vS���f��b��*wqHDq�ޡi�I�B�V0�Z<%���(Q(J��K�}@���YD22��s�N�ZlV�8~���b�1}"�E_��]�o�EJ�gj���w��93v[}�{v5�c�KZţԺ�-$QǺ��X�	�R�A6��u�voF1�&A�aĺ�b��n�҈�
"J���Tkvw��>���Ux��6�F��VA�Ȩ�G�K3ª�Q�(�� �k�{�������v��B��/�~m ��A"�B�{{eWtu��'�v1|��؄evί}o~�]m4�Ѭ�l�yt��-�+(��u�ʚ�[���e�Bہ]��h'��:u���#)q�F���t����ʁȨ��&D(���7g]��(}�<�_F��q�r1�
���P�$�/n��r��}@Ȁ�Lb�D�G�>��A��o����wF�F*�����X&sǼ!	a�����M�CWl�V�8�\�Rw�Өc�:���+�:u��fn(��ov��.�ۺ��嬡�k���ԙ�������x��sܷ/k�U��ٹ�:�e��N����9b}6�-P���2�-Y�ٺ�k ��wtA�Ep^c:�@�Ef�Ӑ٣�Oj�ұ�Qǧ�meX�ŷ�	�A��ӛxDRt��:�a%{��q��݂���heB����CrH����2�b�]�W��}��%f�����vܖ�^���Y�I�U�`ϗi��˭�[ք̀^cB�˸F�`ۧ����;����ɉ���v��w�3L�b0��r�ʃu�>4�w��48��(b�i�W]ڊ�uC3!f�*;�L�q�"���������n��T2q<ܜk^G�C{8B���8���Q*8�R�_e�ƅ\�v�]gwt�A�{o*�I+UT&����7ͭ��Z"����g+�M�w-9uٺ�j�x�z��\��.�5n���t�\iz��
���޵���= ������3N�NKmӥH��I,�If��j;,�&ݢQ�r.۷6n����)%,�%�R^6%W�vwe�d�嚼ז2�#-m�-�˝�h��Xj��{w��-(���u�mb�j���͛wyn'OkJ̆�/k"�l�sk@��)�6�DR w,�Xۍ�m����y(OkrK-e���%J^�h��b�x^[���v��8�۰Q�nH--#7Y�N�-���������qfKk6˜PL�frfIf�N%6�q��kvݏ�'ǡooE+�=�_���B�D�Q T�
�YE�#b�_TC���N=�Nb2�U(��2�lyB���/��2!DH��֒e���mP�T(��ӽ֞�@�� �(���G��*e珡,�:�֩I�4��+�ͻpFm���4q��e�zs���,�n�gGV8�|�c�^��8�nb@X{fH�@]�F�a3�����"�y�#5����u���iA���.�24יv�.��dv�pu1==T����E�{C��D�(���A"�<�'��_h��b�����]3����_ L��29G�Lvb ]�E�3�W!��X�g�;���n�1��@:�䫽���uT���}�id�MB��]�F��Yw�1�µ�!Ewa�z��FR�	�P8��@�f�}�|�c���uWs��LR͐Ԧ�Ԓ�b�mv9�B��e�z��uc�V����+9���@=u�}"�􊈕�J�^��8נ�Ύ�qKs�c��څ�H��/]
=�@�t��(�k�-}z��7;�.]DN.f��F�A��������0��{��}>��Fz�=���i�z�6P?W�Q���q��FE@�dTD!"{��i�M��w��8v1| ġ ���$���'��ET6�W����0�ro>�P3q1r��'|w)|�%)�\=�{����<~�>~�y��$��qM6��]/T�蹞׍�ͶKu�m�f���]vM����K�8np���W4X�}i��(���˜��
M�ܻ�b!��y�ͦ�g�u�n��Lu���7=kY���Jt�Q�O���u.6�m�ޞ�܉�u8麇ά�nv��=O8�i�2õ�>�@U/Q�����r�"qyp�=�����_Q�}, L�P#�-B��aex�@�no{m��Ӱ.�@&��B��_x槟Q������"��A��v�h�q�(�fRt^wbϔ�/Q�R��װi�W�	��Gj�A=|�N7=.�'��iA����u�,�y}"�D(���\Ľ�2ȫ��7{�mv��w�	����G����9����w.�v�.�P�]sJ�6�d�a�z9�5�>��PA7j=�q:;��X��u1S�������^\wrH2�IV�����E0#R�c�3��L�ݼ�wR��>ub��v�[A`�y�]L��3%����8���qw>c���J'LҀA�봻X��S�{7B5��bA��|a�I_M홗�C7��vp��;bOP&� ��D�+��+ �O��]�k�{5z�v�:;q:;��X�i�Վ�'�}�ܡ@���r@�.��>�7�H!���N8qΔV/w���fE�"�Z�����E"���yn���%YE��17b�ͫ��Ӎ[+�lD�(̹�э��.�d���G>�C�mz-n�7j\)��zZ����Yrs��b���(��<�8ک���7� ��(�@����W��^C[}^�0��:�ڂGso��Jy�Z�veQ�5��0�h"���ʐ�i���sm7ʌ���J��$n׮B	]|*H`!�t��(Β{���%�A�	؜O�tX�<yn�k�-z�����Q�Q��1���6/���{��p Mcb��%J�$�D��t���C9���H��3"q�,�{� ��G�����N&㜨�^�w�������G� ݨ"�_H�.�m�3�
 ��(Βw���.���[C̞��ؒ�{H���AB�A��K��^f��:�=�x A���A�Q $t7&')Me��r��wp��9ʌ��- ��Kȳ���JΟ��rṹ{�F����e�=��[��|�Tڭ�9E��j��������@�dB�B��3�A���(�um�;5�$�}egP1_B9����Wf�D%��&��f�xj�;Pĺ�p�L4v}|=����v��ڏeC�F�e���k��}Sg�_q�D!P��@�ux�l�݁:����N&㜨�@D�aݨ�&�9����T�#�_v�DH�
���[o����ٮ"�d���}�"�(W�S!k�?H�A�W8�/Lk�[��r���;.&����8> �P����QJAs�0�~Q	=�l�Ύp�-q��>�V}v�	�py�T�<v�1zd��f�p��k����+o�i�e5;[s�߬P�l�a�Ef���sL�Ef-�Ӻ�]�m9���s�T���׊�lktUΣz�汑�m4\Q/`�����gh���\���wa�Ž�a�KR�z�L��U�!vl� �Y�6����f�ֲ�csx݄�\���'�����]�4M�MM�����BK���X�sωo������D�Q��}�[��!m8�Z4��?)C����^��a�cN��+�;��b��l�1���3�ܠ!�0��z��|B�4���?\�����Cn��T���\�Q��L��b�ړ�����*��O�J�uOM�[5�$]�A����f�A�����T Ȩ�"ȝ��J�S�ϕ,�:3�j�}����q�6Q�j�=yy�����<)�Ԙ���a�3t� [�ج-�ڲͷ���e��Po`��-�p�Ů9��aïZ���� ��3/���G��c7�W��yӶl��JG��QM9T�3���X�
���'*o��YDo!��f�[7�$]��I@��.���zH�ڀ}MzϮՃ뵷S����ծQ��3��P�� �@�w<��6�p�->�Y n�Y�ϏV-q�e�q�PF�l�8��7��7��^�$ݡ �.��k��y6�y�O[�[9�$�}e��$�_�S��
�[?n��@�u4r�x��˻�SR\�X��X�������7,&�I�dF>���Cb1E��CH>�G���B��v�1N��L�c+3*ص��Ջ\s�k���qz�^D�R��ŀ�B9��(�򒐶�+��+� v��ݙ��:(ɡ7JS��x����1�'Z����ƕ��Ef=ų�e�}D}9�mЮ霮C���z�u���*���K^�����Ci��m��#;�r	�m��[�Q�VWz%5J�N)*&��m.�Xh0F�;׍��a٣WWuv(#v*�ڵ>�_kL��f���U��x��Y,{(�w�n�o�걹[oփhW���ڭ���Ζ�_���F��jd�i��֮�w�_�������0��m���~W�x���;ד{*�<2?Q#�m��-g�dw��;ae��@��yi�ͭ�~�G<}��E��� ȝyӝ��l���Y�����}�������(e���/78��t���)n&�V�7���#�Ue+�E$��ζ����q��ۯD�@��f7�:�R���q\�G:���v���wm�my�YP27vn�^����K��j3-�z�RЪ��O\(f���K�����)n ���ڪ�N��$�=����������%ug/�so�[A��R�s�z��A�3]�o��%���3�=�?�m��C��m��h�HH����$}�4B؄� ����cv�!5B�ǍU���G�F,�0Ӑ�C���� ��+$�y� �0� 퇆��^�yJ�%�����b>щ�&{~��yc�w�GCاK�_�M�1�C��&��j���w�74����|�x$;�8ʬ�B@�G�G?q���}�� �$� ����a��!)>���H@��_�`��~� ��'_�!������_���� ����W���l]���4)cޤak�P_�{��{G�#ģ�A�͠k�a�a��>A��__U�\O�b�?�d�H{��
�Ǯ��lc�؄� �/��$A���7�A$c�2҉������G�C����! @#°-�=�#�c�{
�a��R ?w�H����tEl��I��~��P~��%���A��BB@�F>������<�ޏ����=_�K*��U�Į% B�/������_��^�#�,���Z��>|���3�Y=g�B@�G�{�=z|��6�O��kKR6� ���@���	@"ӥ�� �/�ͺ��>0C���*��!��0�~��(�,,��m�1~�J����4/'�Bi`�`�ĽhX`U�vO8�sg��A��J�>�jZ"���Z���Hڐ�����K؏A	��蘇�_W�F�����9�x�8{�ޡy�A��<T'��CH��z_G~��h���>�։������ B@�G��/<z�7�7�DA	/����HX�� �K��_Ҟ����G�oϧ����=H��I�g��^���A�|��c	J_�>>LX����wa����������g�5&V�f<���	q�`7��z!ϔ{�hgِ����/08����x�>�f�	@}�������$� �)�~g��?�}��Y��y$�=���z��¼X}D
�0��KCA���W�g��c`��g�@���]�Y_�rE8P�*�c