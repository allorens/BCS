BZh91AY&SY�� ��ߔpy����߰����  a\u}         C�� �4 �             �   |�[m�mmm�l���ǆ� ��P< � )�4  � s��׭��ܻ�׹�s���L��]���z��	�{Ͷ�>�;�q�=�R(���C!:��zi -�;1v��:4j�  yJ��6��uݔ�'�'xz<�[on��]�%��I�u:R���r����
���;�x�׸i�@���Ե�OfQJ�Q�F�� x Gy[{�&��wk�'p3���G��5/v�m�׽L���ĺ�@`�JHRn���OmRM��k�e7��y�oN���D��r�� �c ������h[��.pw�Q6o6v��N磽oc^���#��ޝ.��xz^�J�R����y=�OM&�T�a@� =�ӌ2!�E�����X���w���]����kK��x��eV���c�{��=�==�����{�u�j���'f�6�                      h �U<C=J�R  ��` L�C ��!)*�Ѩ� �0  �h4�)H���       i ���`     ��SU �&����46�z�jz�
z�(
��&R�(0� ��� i���G��ޫ��޷�:�{z{��6͛�r���C36��1��6��f��2�����f��ݹ���w��?�s�Î��NH���,kT��o�F錐����a���Z)MBBld'�@�A!�UUUT��-�[a����;�~O�oz|������=�x����"�ig��s��`��(��ha?"F�`7��#�~��H��d��|����pz�?x{9��"��*�'�':z!\�K��	��DZGb42xx`"�

/x,m0�z#�0A�Ȏ�">N�GDN�e���':'o�6�4�&Zfaֺ�V��۟# �|�
����I����� �3I�,���'zDx��a8?xDf���1�<U�U1�:A�xy3	">���L&\GG�b@�f�$�T�	��fD^Lx��1��$C�L,��	⪦>AL�'=0�#��G�K\ǆ"b/��c˖c�1&Q"P��̘L�Ɏ���O0�(����"&fLQb�Ŕ"dŞ8?rFh�}+�BW"��\���3	g��c�0���H�#]�F��>�R��ӑ	t�[˄�Γ%}1Ʉ�X�D�<xK#�x�ݎ߉��G�I=2G�}�t䤦RK�J3�I/�{	����O�C�=�G#�$�O�$�I�x�YfD\��8K�?t�K�N|@?v>A����GI�L���B��x�RR��ǉA�K=���	)�GD�L<FC1�ǉ,�f:a��ID}�&^3	BcS	��>���#�%�KJ*rbJ&#��5 ����$C1&1_�鏸53��"�$N��`��c�b��ç���Dr ��}��7s��KGK*ȏ�G����`�%��O��`�#1���wН��\�$�G�e	Q"QC˘D�_"X�"%���$�@��B"q�"33	�Yew��$j<tF��$�,�f<@�BH�va�P�<">�h����))<�RQ:#u2�w�َ�H�&0�<bG����3"d��=Q��'�DE���ĿT}x{H AD�P��&{�YW ��O���xD�"S;�x��D��h�J�	��BN��BtN�b"Q���0���'�?7�W���D�r%�\GD��I4' D����t��"�#Q�Y������D��0�ȔI n0�X�����&2I�83	b[q)�F! �-D�#�CƢ|Q<�Hn%��%�B`�3�?!G�В"S	Ą�Q(���'��(g"~CL�"IO"Q8%�L���"|tJ���~X�P��%<"^$�p~�����{2���<Y���4܌�c3���J�~Dn0�2p��)"J���ÏН�"kܘJ��K8/тX�"z'��2��3-z�r��G�p����&$N�+�؊zaɄ�fS*̸��f�f����3%�'��Fa\�>fxy��_c�t��f�,��D� ���1��s%�Ȳ�)��w�35���!$G#Å�B`�Ȝ.�2e���G�!��#�Qf~N��/� ��Q������O_�=��e4�<��==x��zx��SR�iQB=��G��X�y�ώ����|��<�%,�1fp��Dx����D��#`��^��$��Q*؟`��X����'f)���lDI�G�Ij%0E�$��a܎>�D��c�e#�DKcĉ��~D�V&�8u��D��}�#��N�P�S	��&DKj%3��#y�:a¢$��%8�%2b! r,JǗ2��bzW�P�%	%73Bt����bdDf0DL��Q�ߣ�T=�OH8<���J O]D�آ��O�C�x�'�Q)�)��a���Ҫ0��М�3y��E��<`�xs�(�:X�L�	g�؈�$I:5S)$' � ��BxN�:�B"'��ď�"Kq(�t����'�7 �D�ID�܄�ID���ȝ(o��b[L��ju�ڬv��gS.���䮝}��%	Q%>��	�&0���ȄNL�	e�Jx�0���N�p���LM	�q&O~��'i��y�p�\N�>1�>�p��9����'���<D�4��#Я3���R� �4��D��Ofd��q)%(~e �4��įR��L{�}BP�A���� �fhIy3BtX�f��f�C�gt�E����O|}���Z8h�¸1~��K�9�iy��|�0L�X����O!�x��Fne,b�b���S)���a"�"&�2916#�_b��GDJɔ��DtN�ꎒT�CG��89$~Dn�~~r&���F�">���Ģ=��"P�$~����B'��D�8O�"RDn�F1>(���zE��I�負Dʨ������aMD��y��G>��,��'���y�&<��,s"|'�"~f�xY'%��N'`A�Ȕ�	�'�~����Q)���8'�0K�OD��"(I.��~��`A��Jŋ$���Fc
�I�.a�"!����Dn.c�	�Q"7	K3�UO9��aÇ�G��0���zz���$$G�d�����1)"KȔ��u�8tN�"R�:�L�,Dg����S}���N"w�G�&&F�#��J�!�y,�vx�PF ��:p��ϑ<�Q|�L8=9q�����RQ��G���f"ĴP�#グ�	���>E�����'�>���,�}	N�\��=�D���tX�����a'���f:v"A���$J1�)�a�	����#�����9=����H�=�0F=0����`��6x�� ~HD�3��� Ē�(��'G�w���!nc�����9�%:P�>(�E �>��Tx�$�����9Y1�*�cM4Ʉ�M0�؉H|MP�L�N#ȁ���_LHtG�Y>��D����a>��a��"I����� �7$��y�<(N����LpF�a<�]��٠�R��ȿ�Jl�#�&o��l�N8�������'���9n���]�F���Y~���,U��,������r�<v�z�`,0��$>7�ޫi����:�8�,���y��̂��{���s�@7�V>�0]D���	���w� �`���%Q��$'-R�C�OO�~	Ӿo���l�Ǐ�(Ř0�h�ekǩ���r�����lm����<wn�$�K/��w��3��������?q�I}�l����^g��i�p���o���9 �ɍ��^�����8��;�vs�Ec��Tf<���竺���y�����?٤�\��?T��~㕇Ko_�?n�����s���;��*�%��-��s[;+1�'oC	��2x�P�OZq��O��,�=�]��|n61<�{k7�tn)�s�s,��wƼx�s��ﱙ|��۸F�2*����t����a���Gss3�b/�������.L��w�U��D��>�FN�'��>>��%��[��;����M�z=?\d�p��Ū/N��?cS�k�iZ���=�CTI��Y�p��$a�s��f��{Ėo����yg��*�pχO3�����i�!�w���M��АmG��z�½��'��&�?��l��0��\��������#n��JCt��)�k����}c\��e�0���!�)��Y���{�2�O\�f��=>���{w���E�Bi�t=���~;��0�ϋe~���8~t����o�~=��h�J~½�L;���.L���x�k�9�t��rOM�q��^`�o����K�r{xfb��^y�𳟔�p�S����1̓�罓ٷ�������/(f��z���~��x��td8O=���$E=0�qy`��u��w_)�$.Ø~;��+��<���O����@���;��靚۷��3�폵g�Y��ȓL�w���Y�.zB�x��f�-�W�X�>-MY�u���і�+�\��&�G_=�z�9��S��y���V9�I�3�nP� F5��<㏻��ujN|,>�
��y��{���o��9�9�At[z �g��;�f�;�J؍����L��N�^�N�9�R�����Ȗ� \�7�Z�9���߃]��P���3|ƕ���5�W��)�=l�?�,[�k9͜��7��s��=u��c)��S��)�{��3d6�m�fD0����#�O��1K�?m�sc�_v\�5@H`z��5�o��R�'��NK�i؝_F�P�#'�t疌�/�r�O?(���Hi�8��3��M9��$d���M����nB��7r4Gj,�^cr�$�+��~�a��e�T�E���<�mg[!�݆���M��ٻV����{�6�8��Lꎣ�:�{D��������1K����8������ꟲ�R���0q��&|@��{pO�'�ی��}43Ϟ����d�ƙ��K:]:�e�Yg�Myy�y�f(��~Z�
����'�(�Z�RuÁ�L$��Y�	�@Ε���ӛ㱝�Gޏ�j<B#Yy+���JyQS���W�4��9Gz{�ţɫ��]�����Rc�nc�}�\����c>�:�\70�13�ύ4f��q���3'g#�U�<�GH�;:�S�ߞ\�����m�X~o��-���2���ί=$�у��9�O2n��qn���f��cS���7ߒ�m��R$}��j����a�8���y���}���IFF��~*�L<|p�TZ�	K|z�Rk�i2:d�;�ݸ;<f�s5zщ�8a��o�D�����ld�q��&�;pU�U�nN(��z3�DH{FQ��9�S7i�tX��*�b&L�I�y�=OU�U����{��L�y����T��{D�~,v��e�x�"r��L�Ty/������z�&ޝ��e��x~�ʗ�n�s�^{5��l���5g�"�����9�(�L�N�ĥ����l'���DG�:�v��8�ӛ�[Mr���Ǫ.w�hU>����P�^>��+��]��e%y�q[�2^xv5�����j���+4�:�|n�d�_���g��u�s��[8,�� ����̆|���.h$=[�F�SL2}�fӚ=�#�ųN�ق�۹��L��na��ѓ���f�N{:C���ݡ-�ڡhD'BA���X3w�d8��I�#Nk}��e�L=��FӇ��F��x�W��	>��)5��1{{�
���@�^�1g���>��e�G���;S�j}ˢG߭��d}�miE��B[߇JI+�9��'�^��32w�0Z���~'�C�Q����?x�r�����CҌ��}	h�G�1��a���>�3�k�Fyg���>�2;���ssN��dE�����Rs���)��h�?;�7�}û�����bFncgc����n"�
�^U�+���|a{ָ�2��/=Y3�(��gv�����rUݞ�rfϪ�$,<�C�s�kf�:x�g8h����5T�������6g�_�8�6޷�C{^�p�}��[����;���$�a��g!�S�[��=2L����b\������d�ό����{}����|9���i]��雏�3��޿_m׃�!>ζ�گ+����"J�%�,,�s%0�=+ef�P�5M釷�;�OxyA-�-��`��{���e��t˯MbƯn�m�����?���l���p¯Ge�4��.�͗��}Y,�9��DX_�^kk��9����Y�y��2�4��"�M.M!�3�,{�;�۸����y���S��h�s^��|or-���C�_�!.3�e:��fy��>v�������LB0���e �:��q���i�3J��R���>5U�//c�����z�Z���G����"�k6)ٚx��Ǆ�G�	\�`�כ1�B�W��T](��q�6�oώ�2;���6q���V���_�{y�Fs���y�����C�x��Z���(�����a��?U�Jn\?�y�(��+�V}�>Q�絷+��?v j��Os#��n�ff�wf���#��zj7є|a�M�颦t�-�ʇ�^>���=�V�$���~w�o�o�YN?�N]��O+�w�k-��<t�S���7n�=>_R��d�gN=�S�����b���G��>�c��nHS���l���JӇiJR�q����!mm3j�D�0��vHX�,#R�MF�p��]a.�ô�%�Rlf)��	u%nՆ��h�]��L��p4�;*4�^�rGn �m�$��Z,�H���~
xј+ ��K�1�;y��;WG��.�1ʬ6S9�%�['������/���*n�0����ov�(�I>`��K�(��F�4ͨm�뱬IY��5�]��hy�F�OuG��S����|�`�F"��T�D`D���[͵�na.�\�~OM{]G�7�3Hņ��y��{b��b��E#J���͠BE9 @���߫����k�����WcRmfT���p�s"��S����Ô0DJ��V1G���W��7�ܜ�����i���H��0��h�8X$F\�5n+�[>�j��YhI�v�t�(d�J�>p��B�R��y�,�]�ɡi��l�ژ��e��]0�3=+�0��M?F��힖��3����.������W��u�^���G��Jէ�|~�,�z��>��d�nҟ�s)/�_��֜Đ�<I�޷5�p>�S���D�tz��6��
�H�4IVR~n:�eWv�G�Xr'���\ު���ҧ"�o�;��6�!-�aԫ����lwX���7_�ޗ�o�����!���� �D/�C�{�L}�ӻ�v�h�g���;8ܠ޾�Y��9�o;�4��8/[�1w /�$�h"���YԎ_�	�m(�qu���--ʎ�3�R�2�W�h��zC��I|E�~�Q�10��� �m�����_ ��*�8$F/�"�H��u�8�ju�׶M���٥1Va6#��.F(,b���������Q$�o��7���Q;o��8n=�q��]e��uS(��p��}��_��� ?���c���'��	Qi����ό�yFc�cs���06a�l�d��A�ք]1Cv8d2Lc�\��ka5��n�&��xqoX���n�[�����s(m�=��n��ۉ�^�4���vh������\�!��8����T��o"�ˇϧ(u3�S���-9�g��lY�S��}ڽ|������,�I8�:���2���OD����:�?F����q�Z�yr�m�xyw�e�Ǔ��<�w�gjqn�L��o�?f�=�٫6Vf��oO/O_��ׯg���wwws�W��^�*��ª��/�UEU}�{���^*Ҫ�aUWU_+J�^�*�W-*��UqU\c���9��� �Y� �$��}�󾲪�k*��ZU^��V�W�
�����g��y[YU^��U�ՅUU�U�W��Ux��V�W�ª�3A��D}�"���@������}���z�ڨ���
�����U�*��W�wqw�*�*��ʪ�W�ʪ�������k*��ZU^��V�W�}�L�@����w�ʪ����X��UQU_+J��ZUU�����_,*��*��ʫ�W�ʪ�������0��k*��Z��Ŋ٩�]���Q��q1Y���z7��f�D�V���ǳ�/���k��z=i��t{��G7��F�i�V����u�um�äN�$K�	E��Q�,K����҉�,D�D�(D���:YB&	�,��	��$�&L���ӭ���vL��u��""bG��DI�	�8t<���	�&	bx��b`�xK�0���g���H�X��0��t���$$I9$@�	"H�(D��tL(B�L�0� �>3������B?^��kػk�5�
5l��Y����߶�[o��2n�78��u!Ic.zl:�[Z-�Gi�6��BWϭ�&�o�-љe��Ř;,�k]�q�س=��k
+)L�L�k��݀0b�	���m&�J�Kl�
�CL��.@Bk4Z]k�؏�=y�z�#W��e��lv kc4�Y����쾛9������am;3�Ws�о���I�u0rn�Ͻ!7�w�{���T�y�k��y%��X1wl� Wf���Z:�R���nP�νB%!oP�G NB!N�I�	h����h�jB�Vjh存���ԡ�������X^ev�v4����3*K���
XEi���K�`H�3R���(�f(���� ;P]T�Q�l&-�V�lu��,pR�5)���w�-�����m�7h�S�h�@��;�ɾxg��R�5�,&�J�눛L`���XN���Xh�L�7�8̦���� �Ji��oth�vM5�1a�h�Yw6@�Y�ۇ�� j���\R`)F�	�mMc[0G�t�Hg������	5��j���u}]�9�^�|�(x��B�VY�ұ���n��33CYsZ��М&S��Z�b\ͦ�����R�D3��Sid5��+�J�MK���.��p�3���X{M�K��ue���]�{v���$��w���6H,d����R�������5��qilΌlr�^�|R���;��m��h�k4X�Z&�:�腘͎��kS-�j"�q��),��#}sbdk����\�)a�YV��.��L.h,v���V�*r D��6,�7=���F��º��f�_�b�y��tB˭���P�]����6�Y����dԛ��{�����ĩ��9�u�^r�d��mث	a��e���.]�u��%��[r�C:�m��Ƨ�mi
S5e��m�l�kg�B���1?/��}f]�K(Ţ颔HY6u�mE���43b�7F��p�t�����6�T��6E�3m!��!6��� }����������������ݻ���񻻻�wwwnàۻ���|�9��wԪU1UV�o8�ξy��4N�%a��������N��Q\�{3U�Q�����u.u��c���bf�Z���v�(�2[�6�e4��5�e�gfhXگA�4����(ۼ6]�Za�vKd3X�:�H�u��쩖���3P���U��ɮ��F�[G۽�u��P��e`�zQ�ndvv�N���bb�T6�"����mk!`A�P�
4�f���Jҵ�]It�ԅ�Х"��zOwu����.��F��YQ(������K�k�0��J�8�B0�� Fu���@�7
~(}|��O�����ZrN�<���6#��C�o��N��i`�;�j����M�33�'�$ʹ�����Sٲo���B�u��p��SAX[�lw(�����0�M:'J�0�p�8q��r�]6���QsXf)�`؏jk�@�z�=���0/�_q���#���b�њL9Y���4We��|q����Ǻ8A�;ɐ�$�e�w}�Y�>�̲��\��)s���Yff1���e�����7u8d�JiŘ�{��v��|b�4�6Y��4D�Ή���:`���$�@�,!�{U�i���^m�hp���I�����L���ղ0��bt�>�g_��U��m��Wwra�[f��4ɾT8���Cm�z��I����_St�)f�U�m2�}�k���3�vz]��rd��%|,D�����>�pL<a��D�Ή���:`���C=��Dr�WFNif���W�t}�l�}�d�}O���"������\!k{�1�1���������*��1VKll��������M5�W�]]Ķjۦ���4��=�wu�P��!�^�R���f\�O�O�Pp�҄L,DL,�(J8Q����p�Qx"����Z@�~h�F��E��%e~�`�Bj/|���{�󙋫�s�.�#/�Y��6���|���8��;�g�bo$��ES�$�4o�	�b��9�_SE6%�u)�&R�ҹ�4�����H�.N-z�C�'�_\�ލ���C`])�S��v�W�y��7!�)C7ẻ��H9jz��r�y���nI��}Si�����!CfS�%��	:)��<��iz�+�ZU��c�&��C�m)ku��h�`����%	Ft�<!�؂�f����Nf�J��pUM:M �4�6�X��n�1}��-�`���Т�:����V�o'-�|ɚ|f�Ǽ�]��4�:� s=�X.e4�7=0��@�C����至}�:��*�O����p��D�DL,��(J0æ	��~��(����t	>����V�^�+FG�K�
v�1%d�f�����7 ��r�a��;4>����6n�?QAQ�Te�X����.2h�||�S��&ӓ�w���H�Jie�C�s�͘J���i��'��[�b�A�]�x�4`�5Q�ޥUe����Ǎ0�LĲ����p���2@�D3 H~ =σ����O����bI!�"^��\8��F�y
A^�@CE2�.+�0��I�C.��1�S��^�3����<����Ȟ��jR��v\L�c���O>��d��b3^B�'��SΓOY�O�a�X�P�"P�c�
8x`���k�H��a+�6O�.$��m��j��*}�3��N��p���4�2vP�.)�i��$�L@ˤ�5ޘƮG��a;��r�	��\>���<sC����1;�[ǩXN�l�iՂBV�H�3w<=:{ý^�� /� ��_Q���li�j����.�FD�4}<�Dm�y6$û���y���"&N���5	��M	�!��}��k|�8˴�&�UJFQ�.�*C�����-A���P�\�n���os�wW~�)�=Qݤ4�8a�	�	bYBP�BQ�0N�������B�|{�D��3!�����d�}6d7��7&��5��0�s��Mh5���
"C�h������ɑO/�\�d�����{!�u�]7.�2��f����Jv��J�Қp��w79�_L���&��PԾ_�����7=���Z��G2�_/�h�'��G_7���Z��Ke�1<��6�/\���٤��t�|iei$�F�?&���X�iD��JHӄ�0�#'&��K�����y<�e�L�Ǟ_�_�a����y��������y���8�'��y�'��O�<�/����Q�<6Tv;4O����-�<���ya~b��y<���a�O/�痷�c��_�~'����_��O�m���'��>cɷ�c�/ͯ�ח�<��H���~N������<�yz�������N7ry��y<���/��/��t��Ǖ��:_�j�=�^~�~�Y���O�#��MM��IӤ��JK	�4�t��SI��~�M'�w}ߧ��#���}���/dpf.��*��}�lb��zw��v�N��EwvxZv��h}r ����ǒ���u�{�C��t��&\�}�sӜ�Fy6;�Ӹ��(K_���q�'7��PoIyՂ�"=���{�����Z��NON�ߴ�?�����ݷ�+�XO��g'��������韏��}y�www��������������l������e���������fe������M,�4�D�0�J4҄ӂ'��Ƃx����k��q��r:Vn�g=����?0�R�t��%)ڃ.�M%�Ѥ� �p-����DK��-���B{U)<?:0��0ve�Yfs,����K�P���%z�	J�Ţ8�}���k.\L-�6�Te���1�'n1Xq�d��C$��H��!<�a�Rije�e~�G{&��y��f����%R��uR���}�lI�&r���NQ<�h�h�~]�A�I82Cс�)�!���)�\)�y�8"kc2�
T���taM�j���S�u��矟6�<�<�/2뭾y��V�d�w�L�"�"$82Q#@��	�2 dL�0������$�C�(N	��9��A�'A?o~'�����#:|�>�����8V�ݹ�qaX�"c��v!� $���$�!��jT�Q%��P'�cNFD���3�L�dVۄ��&pa�E�9	���0�A�>���n�!(�L(�����ؖC�'�' �<@RX04fC �O�Q�)6+PL��$�Q6Ăr	
��d��6"~
L�,�#�K,��O���`ɱ!S��HpDI�2S(���0��JW�eZ~~u�o??>m�VI��4ҎpD�xЊf��5<��[Κ���zi	WoJ{��:P�POx��ǯ��=䭬���
�{�����2�6��K�Ua�d�ļ�MQ�Sf�Jj�5t�)m���r���Ҽ����}�+[�ch3�&<�����V���<�qۈ����s�(�.��b���ۮ󦻿I��R֎N�>a��Q��I�<Q}
l���d�#$�e��xd����VT�R�e�Z#'�җ�~r�8�1:2�~�U���ϗ��SE�c���QFH�*;���`!����Ȱ����lD��y$�2�����Uy!���r�S�����sG:Y!J"|`̄�l�5%N�#(�"DD<��0��)h�ň�]W�8���5�3�~��(��C	@�58R���ȰS])�S��d��CB&���ʿkZ�R�d֍<%�ٖ�82"D�O"�C�ج�>]SQLyt�Dr@1�L����0����m!�!�Lb�e��~u��ʹ��#�0��2�.�ۯ6���6����UQ� ��S���,&%��$�p�"2JD��,	�.�ۣ��Ĝ#"�H�kDm�V�C)Tv���`�"|!�� �	S �	t69����D:���#��M&�(��>��e)R>~00j�uN�>��2I��DF@�J!�	��($�	�N2i4"{���=fy�]H8*��A>�&��A���G^�?�'�B������!�?C�DChp��d,�}dSȉ9��������#!�DD�R}�t92C��I��!���\0�2""J�!FJ�~)SL�X�B_�9��H�>e�_:����x��-�e�]u�^m���bc�31�xSN���UTDD���$�2�a���bw�^L�H$O�`����0I�?A��#$�n?D��2��n�!!-n���ax�Ѫ�G�FIT�p�(�]��mDd���aݰ,JHH��Cc%MB�R�!�
�"}���L�i,��#=;~x-�XA�:}^�E�v6�hDd20,>�'NL��(|�Q��$�fS����M膆Q#Ҕ��B�����i�P�
	imX�� �F�f�Ue��A�_�~Mde*����`�7R�pd���E4"$DD���5	�s �ɰC�4ȡ��A;Jȧ*0�""J�d>2!��X}b�h���y��K�b���*�����������ʹ�u����ˮ��ͼqح�TjW�^w�	
�H�H�}"1i�f~D�$DD��%���9H�o��'�G�(rD@�G�dD4}��0f�ACC$��~2T�fNl�.7-����n
S`��Q��~5�D���]���`�����������d��D��%C�N��& ���@��x����1�n�9H�	SBQCF��2l�Ʉ��Ynjmd�$���"d-,* �@rSB|2��� ,�3�(a8�`��=��4=C�="'���Kd�S4jD"�{72��R�>�S�d&�~V��NO
	�`��L�
]�0�:��ߛy���ϛi����y�y�]mכx��}�ճ��ul��as_����$�	1 IE�E*M�BFDAR��I��qk��S����E�B���T�V�e�4�b��#@�Ae�`A����Y�I$�S
z�7�!�������p���0�G���XzE�J�+��3�����O���/���|tTOa�D�☋�X~=�8%Ha�ߗ�̬�'�B�h����ܥ�͆�����L�l)
j!f;����D�+j��d�aӧsM�����=0�nRx$���ÚG2��[�ǝ<���YB�DF~&�+(<��՚Uv�L~��Ô0K�C�LJ2j	��{h�,�0PDD#��bbKi��Q�zl�w�v6�>�-Os4�R�b���=<W!��
DL0D�P��)�R9�F��!�JT������'!�$��xD�?�<tA4�M4�N�==8z|t�ѧ32�FS
��N�=�C|]þ�UPFC��ɥ|��o�>ZQ�|��b!�y��pO�UZ����<�c#0������ZSQ3a��=�F�XD�J[�ָ~�jM0�֦���3m:��l�Yu_�%��[H� V/G�
'�wĝ�0��,�0��v``bK�KS=��O�)��f�c�없���`��bPM�IP�2����fg2�p�0h�Xa{(S!d��c���h��)�L�}:��h��np��0�T���l-7���b���m]J|�e�H´�θ��O�: �i&�Q�N�K4ڑ�f��������Ub�3��#�_��0e��܆�V��$|���'!i�~����(y�8۸h|)R�B��od��{�{�"}!�ðK(4����D�)C|Η�ˏQT�p��A�G�8�(�#��G>$��,���Z5V�E�l�H�)io��T�~FYk�b��"p�M	$�u(hL���D�ta����>��m����tNA���eJ��c����7�E�U��b0��y��|�?>m�	��M4�N�<&�i{���k����]Jܶ�㱕�V �*4�ȿ]�j���n���H�%I�6��"C�ęJT|��dKB����~~̣������.�`�>����,����Oϑ6���J��|�[����4�j+���6`���JG���z��i�|0���b\)|���<�����T���x��~��,��2L��9�NC�cn'������6!`�o�~�w'Cpv�{��ri���,��Щ�	���L膏���Ri�e��4O���y>mo͗���6����<O8�1��4Ï/ͯ�/o/�"��z�W��u"ēJ'%0�$�0�40�0����.�\y~O<�'�ͼǞ_����+��2��<���y�4�i{y~O<�O����x�1k_�	�G���&�Ѳ�uU�Q�S��Ik�����,/ɇ���jO=������i�0�OǮO���&W�2��y��o3��?>a��ח��I�5"~�H''HM'":N�����6�=s,��.azyq<�OI�J�:i:Y:Y�TF�0�bI�MT���I���Z<��#��Zy�̯	��i�������y��~a��<����6����G߱~�d�Q�r�k���[C��겒Z8q@�|
�X� �f���u"�:6���KUO{Y&
[ G�ϧ��saQ��k:�S�I�?�����Z�R�EɏZ�^��khO6Dn\|�I�����CW�O�:ĵ�~��h��xE�}��uO,����(����"��d�3ƽ�P��	#�kW⨚*��݌	*�4��?5wpWq\���։#(x �R^Hs������W��2i<�H�)�ON���r��}��k���M8���È��5B%��jr�L��y}�K��`M�&$9�?uI��tӣ��[_��X��=�ia���K���i�O+�{*�`�|�5{.#��mDĨ~�=��#��b��ɒ�L���b��.�/���C������O[}{s���˸�r�3��q`K쁈�&��P`O�h���-6�v�&�U�՛������F�@װ8���~�ߟ=�����(�l��X��ℳ��M�3�.�������,_^��k�0��D�9$_����v��~�wwv���UWs3337EU[�����5U[�����6�'��0���I4ҍ:pD�Y�;�f�>��*"nKw�u���8mL�h�M��1fͺ�oSF�j"	�妷�5��1��-��۶#l�l�\�j��k����J(۶5m\�K����#�֓J�������ȭ;lQw8"k�t�(DL��l�3X�:��m����V�ڲ�5�6�L�5-���-�����J� �)H����{lkaI5+(:�1�i)a4o1�l����X��˩UlD F2qI?z���$�46bJ���V�v���03.��#P�5kx7�t���1�V,3���s5����}o1]��NG��!�h5�tɝb}�������&��~���t�p�;����U��Q~��P�'C��A��"fS1|�39tf�?��B�{����ág"*��1����&3��_���W��K��y[i���T���4�$u��A@�;��6�h&$U�W��~c�ӭiј(���T�:0ْR�.�����_�u.}&k�u��4����M4�M(ӧO	�����n~Sx}�g.juUb���h{8l�?8ʧ��t'd���a�sp���bx�L�y��f���ja��=�r�#��S�5�a����{�-i��\8�[㣦�G�J�[�z�Yև����)T��2�t�JQk�vq�z���њ��7Hɂ�w��8�O9��z���g���~���>���9,.�G�6h4H@�����$��J�p���<�������<�.�ۯ8�8Ի�]�e���+]�&�-�k���G��3ZbV�-���n�M+T��;4�s��eH���űX5M2wGL�~50:;2x���<.b�3��;1v�f��W���9���7%)I�?Z/��٣��iC�
l��}�Jb�P��~|ۋ6��?{T�MԬ7I��r���u�W���.�<��Q]��qg7�z��i)m��}U��	j:�����??:�N�u��/4ˮ���<��nB�� .�q&9ir��M�EQ�����M��������)����i}4��~��4#����2�r��>�<�пNX�������2�ܧ�gU��.�b�C�=Z�8���[�����)�p��{��4K����E^ԩ�`!�ٽ��Y}�if?xF�Ϯ��i_R�J��*�I��gT�-������r���0���<tAI4ӆ�8"xG��.��g ���Bi,B���h|��h$���P�����f&M(��
�����$�5	�t���rG�r����Xg"!J�=�����;Xٳ�HE��Əʩ�I$�c.S��j��+�&�럠��̺�h-}؈��^��|«}�HZ����lh�x'�����`���|���d���U��&���'�g�O���i�f��7��b�N��e��)���U���~L��}T�[�F�S�P������Of�ȶ�p����zvD�{`��0�z�f9\j�L~g�#d����5ތ�+N�\p��0?��_l���,��2Ha�Me��OT9<���h0>a�;��^~�N�r�a���e��??<��m"A��pҎ�K4���DW�N	]f)�UD�?��P�xH�������9��@Z�V'2����҆�M�=�t�2b��/Zr��e��7�C��q�ǭs8���~73ek��  Ư���F㭥$���Ȓ(��ﵬ��y�~�,��j0V��K�<��8!����vw�=�X'��|�<��+?9�a�}^�շϪ��6���Y��O�x�$i�(������mѹU�J��t<�7�UU�e���ce�~˶��m�t�}>i���f�͙i���_6�������)��i���v�oɺ���h;��o00�3.�O��i������<��^��p���_���&ckvw��quӔ�m�g2a��'��l�)�1�ԑ�gN�M�z���/�CǑ��g�`{;ѥb�t���	"_�t����=��,D�?���H4�NQ��if�A�K_��ٗW����9��Ԝ9�f��)5�ỵ�y^�Xfx���T;?�N���S��`�{=x����H��eGH#��c��w���aU��=��_(ώ�hLɟja��&��4D2�5����D���ۗ��GC§5�"*?�շ��6Xg�T֌"&М�֗���:�}��h��t��b�e��Y�_e<��e�q�U�D1O�W�y�q�,�'��: ��i�J8"x��4~$U�R&��
Cُ+R|��$�/�Q$xh��@�شc�0�U3�D'�P�0P��D`����խ�I�i�4��!�7����=:u�!
aRHj�?"�h٨��f�OO't���S5MYX�����������[ν��%�0(w!��J���S���nG�y�/m���4nC����b�S﹗�fM�zS�o��n�Շ�l�fj읯q"�Zk��nU����v�9��ן�A���
R�}��f޺����k[���Cɹ��Ѡ��`z62�4�w|����)[>|���>u��x�$i�(���4�Lfc4�]Qє֪Ķ���)��vkK$�[�z��̫{dݙO[�s��Jn��n��!�f��ɨ��o'�"�3��FCGi�'���|��k]�A�_K�Wd��:t����A���l��C��[w��f����o�q�빜y�)��ut��M%a9l����/��c�}j�B�o\�o�|�2�1^y�o��Ya��#��˓�\���m?-�������Ǘ��1�s&<�<�̲���0'HM�IH��R0��&p�SW���<��<�|yn&��=W<�=s����NI��'�^e�O�%�8ǚy��o������|�ؕ<y~[�1�\z�.�L����D�H����������������O=so0�y���y����x�<�'�岟�����7s���|�#Dj#6���$�FI��ai8i�dD��If�$a�ᆕ%�t��z�O=s����4���؜y���/����b]��ǋ�<��0���#�F��-䶞ci���Ѥ��
�I�I�D����MpA7���v���`���LeM��@��CI[�sv=�C>��$���B
�z����ȗ8�Y�}'��1�ʪ|�đ��z�,�a$;%�zl����)�;QD��Iа���&�P��|Zޒ���c�3�ҕ(�^�Ҵf5ņaA�1�b�ڻ������4�yq{�Jon��u����!�U�zv��9U<��+_��u{�]�I�oM��0�⯮��xn]�� wo~��fffo�aU\������U�����݅Ur�333w:I��i��h�: ��i�J8"xM,�~�	���"0��U���l�|0aa�ȏ�8�=|��_�=/��0�Vڋ-�f�]3o���}�?^7h�X��BbD[���b$�h���p!�E��?���J<��8fg!&��W(�����.��Y�qw��su�f,�r?y2���֚a����$I��N]z�K�4���q�\y��m:u�~y�^a��mלy��z��r�.��.Yk��U�Y��4'��6�mhr���SC�ա��͵w�JA���^H뮎L���4����xn9��
2j�E9�T�6p�Z��-6۔�W	)�J�����hv������͹�����d�j"1�Ô��^�0��^��Z�L4��n���>�����M3M��$G�3����S��7�6�`�l��>p�f�~<tA4ӆ�p�<&�~�͐P~��!�&J��'��C$�*��F�C��~�{V�-%^7E�m��r��8��s2��=�~��m�Vn���)������"�DYE�E�$��v�!?����1�u~�����h�=0�����4�X.,�\Lϲ܍�F]���GA��K���.w��u���ѩ������8����X]ufO�o�[�{$i�a�����6���6��F	�e�u=���ª�r���?��ɭ/|�kJN��F�da�{9}a�],Ǣj�Რ�?~����K��T3W���!-�+-�a�������)�k�Ϙ�i���8mu���3��߸oƖaF	�O��0 �M8iF��N�>�y���ʵ�⪢	Ҟ��٠�_ܦ>��LLސw�y��{=���n�͘k���p����x��,l7f�R}uO�Ӫ�����OS��ۯNJ{��}�e�X��b�Cr��5�e.7%�`���;��������f���T��`�-�1�WYGQj��˿̴�].�io;y�_<�O���<�/0�ζ��<�'����)��K�y�]�x����͙����Ī�����Ͱ�0�X�ϵ[��NW�ɳ~kNg]���Z�h�aŭ�l�\A��k^SwY���֊hnU3.��Uc����~F�°��~옞*M�K?ECG9�K�{��/sBC'�@?f�pq�LT��f�0�)���3N�oڛ�0�c�Ϸ��=���OS��+�0�ϟ>u��m>:�:��/2�N���<�W{-r����Z窪�zY����u8���I ��������j�s�sC�Su�j��\MƦC�s�<�R"Fj1K����mi=�ǵ_.����?4j�%RMu�c��1M��>�7&Zi|�ɓ����đr�[���>Fi�h�;&�i�2uW�M-'r�o�b�e�4����+�m8�W���i�μ���m>�&�pӆ��if�Gbz�kN�l���İ�H6�m�����_�iK>�b�Z��l����q�P���I$�@�����#�K)&�3	�I��A�Bm�ɬ�K��V&�і��/�b�1
�e���(��Di:=�{�5�{�G�V�Q宖�Ƀ�=~��&wFk����Z��-�E�۾�M�Fk�}i��[�W�f���C�.p��{��=;f����a�8�>s�?}w�������K:��)�jM�a���6����I���և���>�`h㳫Қ��Mq�>H������g�il��i��M9���if���hC8~?q�Qמe�^i��yǚg�o51�b�Ўڵ��L�x����8~��h�)���9ԵI[�z�g��}�*I'\�bҳ�6��)�Hі��j!� d#?~�vt����4Q �5s%*P���MرִkY��hˬ��OS�Jd5�,�a���_?.���a������4b�u�a孴��ӌ�i���o8��:`"@�i�NtO	��iș4��-�������UQ	Â�����ta���>��A_iG�R��el��"%12��1��L��ST��5�����mqt�_�ɍ%��[�yq4�f����)^:yС�/��u�5u��e�z�y��N2�Զ�q��$�%0Y��K�Ğ�����*vO�R�Wp���6�Mk4f��v&T�M��S���AÄ}[8�ҿ��i�-�yן�?�������/2���<���ܫ��y����߭u��m2�Ϊ�$R��]�M>C����-�~q���t������5��R�}��MÐ������a�t[fÊ/ߗGD�)P�����<����s3���џ���<�
~��p��Ӝ)�'~E�LW���\���Է)���[w�n!��]h������x�|~����Xj���-S�-��:���~M��ܟ�[������~^�^oˉ�����ΰ��_���������RO:�I�R!4�#�L(�'FcI�׷�cί���4x���_��8Ǟ_�_�i��e1Ǘ��<ƞ_�m�'�����0��Ǘ��O�2�
|d��c��2`�G�<�-~a~b�������_��\�����yz��bav���+ˏ/���y�ww�����������<����4ӔF���LFNDi8F�Ȍ4�2�ί�<����؞w'��4�=s��y��4�؜y��.<�'S���˵�=r���yk�a-��zN.�_���lm��������2�0�JM<V�BV�Ge��UQU������?Y� �����
Ɨ��}��~;�1ʼ]�w�tT�ԁ�S�9vL��AP4�ׯt4�Ć@���5�N^�m��>���p�k�}&v��F���2$~/m����S�3u���fs��^�Ş�قj�H�I�A����C���⁻�jˆ�-�L����Ӵa�!��(N�����
!��C��z$QV��2EAR�t�>a��G�'�[�j�f�M����fN�P�'`��!��j�rU��z}�L��7�4�������'��&�p��UvD��2N��"M�����P�=��(w��g\��8���Ő&dXl�F�{/�k_�U*�����6}i����h��Y�lV}��J���qv�vn9uֳ�̳�ַD����U�#\�3SY�v�ݽ_xI`�T�=s��5��6�����/��M����"U����=�J�63�a�,D�*�C�D$y(0VS)R�[4�.��� �"�J��{�}=�����gs��/s337v5Ur�333wcUW/s337weUs7333w��i�,D�<t�D�4ӆ�4x`���h����e�D�H��jpcuЫmb9����5�Ùj����5�8�"׶�B�."�m�K5�% ]ac�rjP��t��Z۳i|���lh؋-���,՛j�BٱV��WGv��ţ��l�iq(�m�.�v����"s�Kc,���G4UìL.h�5������2�m�]�V�/z��k/� @�$F	��iRgt�I �>�~Mka���&b�p��o
�V"R�Lɢ��C�V؟Q�`C�����`�Q�Gb��m�V�Y�Չ�f����m��x���z'�D����,�������d�7�``����	��S�����ũ��~s&�~kk�����}�X�1����5��e�(x{���x�Q-ګ�G��+�k6��y�^q��O0 M4�Ǆ��3�;p���7���UD),�u��e�����L��o�7�"�>f"��SG�^j}�����tTp�t9`�L�D���H��0ٔ(~ m�)�bOOk�c[L�r�nQ���-���U��N9!b�l�]_5Yy���0J��g�0�=\z��]�#G{�K�if{�2Wa�Za�D�a����&�pӆ���|t���۬�Z�=�C1Ӗ�����U���g�C��r|zxn05?d��75OA�k�)Nz0�ګ�תS��!����8�����|Tq��Jf��?LK\y���^c:�i�ff�M�y�(d��o�_�^�ѿ.�m��ζ�DEmu�-�Za�ad2���t�i��|��|��	J�?S�-�M��:'�Śi��:`"@��8h�8z|t���w�*ªL���Y"�F�Ǯ^&���g���ϊ7Gߗ�L���4a�S��?}��Yo���fB�i����B@��G|���[Ʃ�D7Z�TK3l�H�ͿS4�*��/S-��ׯ�z�nOX�+/��u�5��g2}���و�R�L�u��4�;��7�6�:��Y�ԫa��i��6��I�2�s"�[T�c]�:�N�x�0��LH4�������w
�jP?5$Nq�Z/�,��(�u�Á�ޡۚ���.�j����=?B����(e�&v�K�,m��A��I$�@��?��4�'�&��-y�\7�~o��c',>0-Ɔ�s0���WA�8��1}o��Ԝ[��?4�G��ֳ���R֬o�^0�Z�9�m��(JX~�߫�:�J|��Ǟ�.c~��{�4�m�e��2g�J��#������?K;���B��M��Xa��X�)�v0Ck|�5]JE?D���7}չ�2�\��}x}����;DDv�/�C��%tm:�b�QDV*+��J�8�(�$F �i�*�5�����fK��4��2�/�~y���$�pӆ���if�ى��Q��2��UQ	�O�����:���d%{���I�8���em�&�5%&�a��Pah��~��fnj�C]��\'�F,�a���L�<:	�S	϶7&Ûŗ�J]n�̌�;[-�+�	u?FƯ��Ή����(�C�����9�y���M|&	��,��k�c���8�.v��o��U�G�x�M<a�i���LH4�Ǆ��+����J	��UGg��3�p�������!tn�}�[��O��ya��<���a��W�d���R���E���xXy'�F+�]/�S_�O�7���9��\���9�Ʃ06�z�!�t��k9WL�D1L�~a�5��2��ޒS/��}�$N^i����f�4��)��0O��ё|��Q:7�r5}~>�0QG���Ïǎ��"Q��4O	�K4v ��R��j��v��F��}�˜9�,��[HѺ]J|��6��1Zh��A?b�NA�T���F�8jW
(ffQq�N11�� ���~h�d�>��|b�0�����ɠL1K��Sh���3N4�R��(��l�_�h�I@p��I����rf�o4�����~�i�5�,���&��J�2p�-:��0C�O�0�O��, D�M8h�=8|t��__��&+�O�L�4͡	�ǽ��Kl���:�萖*������(�x���
l�L鳭��0��t���)���S��"���I$�)�)xx�QG�{V�١�ݳd.�	���f5����w�j��Z�I�?sZ7��Ҿ����~�`�峚��Zq���m80��f0�O~b��O4td�p�4�|1V<���<<��3՞zh؇����V�R"q2���ݬ�7T���B+������ۓt�2�LU��f��
�-T�p�}��3-ne���uj�0����/���?M�?8��o�~,�<t�D��4�xOY��H{l ,�J��"�"k���?�f4raA� �Xr��`~E�?R�֍2������Xh�ئ)�t�e�g�'Z|ɗu�9�"G|�2�ZX�>u��;�����h��sCf��x�_��l����<(~9��pU����eK���L�e�-�r�&!)���v�0xP��8V�Sk�~4F�S4�3�~~i�<����2�,�&�i�I��i�4�Y�$�0舖X�X�%�d��<`�x�G�""t�D�IAJ쐈���Dt���Ӭ#�d�(��:t�$�%�$� ����	$ ��Q�:&�x�K�a"`�&	e�bX�'D����bX�x�ӂt�DDJ<q!<ai	"Y�$	�H�Q$$'� N�8"tN�g��X�0O�衈�9x���r%'�v��u�!d��\��EÛ�r��rk��$c-.,����pЖ�2?D��5$:	��=g��}$s�� ����o�#J9��k^��@e+����)K�Ԏ�UÖ�f�#�	5���/��}����u�����<�I}������z0�ԟ?��i�٫z�#��0ی=H���A�C�����g����������r�V��&�Vo�����.���{�~s/�ff~���W2�337wgU\�������Us3s33w��Q�K0O, D�M8h�=8|t����UD�)�0N�?"��L�Z%[��2��2Jܯ��G�3rڦ�,���kn�L�:��ܚ��<'��/!�@���4�32P\�P^�)���g!���S�e���ުHӚ���͑�y�v���тD���Z'x�:�?C
h?���3f$9�%oCRt����W��m��|��iî����̼�n��&��*����fc31��em�UUK1b�O5�OC]���MC垔��o9k��r7+�.+�1�	�ˊ4��������O��!�;��h��F��l3H�mX>��bKZ9�Gz�CӾ'LɆa����ӥ5��[L�>gdC��Ԫ�̨�����OL�|E�\�}K��4��0DZU��L;oe�Zi��|���pD��ӆ��:if����g�0TVj.Y)@���I�tB���K���nq�>x�Uf�>�⃱짘+��v���z��6>gbce�v����ә����Y�n���ݣ��v��9�
���0�
(�͌f��3wI����4�^��X֪�<�S�zS��el��,f�jN]o|e/���n�m)��4�m4�;VD����Y�sr&k�хP��'��n�n�IĦ��_�a�""�huWL��>�y)�G	U�T=���B������Qusx}�(�����a`���
}�~0�.%f&	�,��i㥈�"Q��^u�Zyǈ���}2�1���i��UD�,4X?8�2���=K��I:x�R�o�&0���2�d=gC��xS332�|o�̟!���l�m�M��)�i������4��J�Vt�;���GE�ȱގ�V�X�Ҧ���8d,<�z	��D�O��:��o�z4�1�����+���2�GŲ�9L�4�~chrV|�.?<���s�	%	��xN�Y�]Wt��&xs#�|Ѧ_���m��}(|}b}�^���9[��<n�m�h�v�{�l;��rX���&�P�>��=��4|!C�~[���X����4�����ʖc>OHY#g?d�7WaKJ��ϩ���DGg�0}H��S��ve�����1K[+��s.6�̽�����l��(եn��MS���I�-��H��W���ٓ=qN�0�:Y��a�����"P�p�ΚY�o�|����p�����+�.�޷��<UTA6��{�}�N�f���y��?&{qg��Z�|�F����OiC�v��-�-�bct�/�2�#��3�ſ�O�V�Ɇ[-�#N��~H����V�?""�VZb�`�Go�����Ϲm͜F<���ȳ�ߌ�R>s���so|r�U�O~b��5YH�n۬.���\i�~|���&	"%	��%�4�Hت~���rf1-F��#�6��WȂ-!��)m�jw�eQ9ȡ礔Q�W��j�BV%����z��\窪�{�7�y�/|}��<"_n��I>��R���M��F���E��S#���y%�tܟ2����T�?ݓ�ɗ��:h�a\�9���6h��ҧ�S�����z�xw�s��X^�O8h��ա�?~�N���B��iD�9�8�6����
�WԲ���&=�6��d��~�f�1��t�����F�R��w�x'5�[L=����e6p�"&�:&	"%	��%�4���t���$��c�4�"�6�Zs�UD,�?j7��a(|��Y���urF�ak�#��u�������D�{6`vX&F>~�����畸s�09'O!thH��������]�Q��� FZ"�|���S�e4�>�o���K:!���'�� ����9ǩ�q���I���$�l�Rb�ۯ�q��Ϟp�$��&�4D���h�>ߣ�+������#��� ώ3����}�������TwKY��!�)8�|�O�����F�/�ٯC4���=�&��{y^fZ�:0�#�����c��XXn����ٰ�b/�n*/�JSӥ
�C6&�Q�E�~$���*5�>J�&�=O�u�gG�2G�W�U�뽹��Ͷ��]~a���`�"P��"Y��4�h`}�>�Y�}V���lh�}[m�Ө����y�̴�_S�S�҈6�.��2p���\��+ꨖ�����j�]2]<�柛���=Z�w��ۏf��K�0Zۧ_#�Y���W�fÐ�����3.8:�x����<��6d��ߍx�f���u���6��f�>y�Z~m�~l��8Q#	&P��?Y��h�(�(����X�%��<u���agJ:$�DD舔 �H��"P��DDL� �I'�ÄI�A���$H<"&	��DM(ӆ�0�Oib&�&	e�bX�"x�D�0�bYbY�'�B"t��ŉ�%x�|��aE@�A1b<��Â'�|E��L;ܟҦb}wU�w&�-�K;VS�N�u�^4F���2w�۝���m��	��IіXhcb�k��a1e�	������	�����������T)Q6|��Vn�~Wc(8ws�*s���a�(4`�D��)|�a>;wR�_C�/1{0`�=�č֘����q�8�4�b}�ٙ�@��S��͋���*⨉�Oez��H�PD��O/e��ƺ����%ۇ�}���=���-,�ƴ�܊{�iMvc컗$��Y�7���S7IS�WtFtM��Bs�O%>��P]�9C٧q6<�묞��M`�Q
̨��1�ߦ���IO�R�]t��Z�-ڗ����b[�l�a�U����PCO�eH�������~�%F�/�Ii��a�>4}A�J�O�*�D�B�d���0�`�]�� h�_z�~��4�t��eB!�nĎA+K� �� H:A)�>�5"d���Ǥ�z������������e�ff��֪�e�ff���s3733w�M4���i�Y�0I(M8h�f�,Ӊ�O����n�cB��@���%ֆ�.�u悵0ˠ�V޵��Z�-����9"M���<�l!m�c1�l �]Q5�8�fwx�����Kt�����JᘃJR�����m����}���za�m�Ե]e�I�Bueɋ��	]��=��kt<���n����i�Õ��*�h�5���K��6�)�����)/Vhk^����I$3g~�z6��Sm�P�V4�b�d�������λ�#K�v?^�{5|N�mm���4�C��0�?�t0����.�;�Ŷ'�iN�v�<Gr��>����{�}�[����|A����R������5��{�^����3N�/�lD2~pZ���t��C�}-�����rT�֬s.>�&���a���ӥ0588�Є��W�a��0���gş�4�0I
0��if�xӣ�o٧Za��uu�3Pꪢ?B��V�bSg:�����}T����߯Y�����{=>��V�2=\7OS�Z�=NSSI�0��7�$I�#LSo�֘>���i����m�G����Qn3��Y��I���4g2E�sP�82w�&�d���V}'��:���%$jy��Ĺ����u��mU�-��󯟟<㯉"aFh�if�x��������J�X;UTC����F\�a��1����S!�FN��7!v����M3W\�n!�q�_oU�8P����{�v��7����9�a����>���B�O��m�~�>�S��F��r!�{��5�Y5=,�W���0C��b��g����5��&O��w��R�ï4�n�>~pL(8~,��^���=��R�O߮& h���G�3b.q$�D>G����7[-�k-6�#&��h���4R?�#D�J7e�o�+����^ȥN׸g!����r��׌�|�u���gI����	�5SBkt�+Q��ɅW���u��eii�u=T뺫�q�?VQR��SG�*�v�>O?�(��f���J0�i��if����W9�¢����8�2�$荕>�>zIh�JJ�-���Z��2G���u jr����wq��OԉB����m�	k���ĒI!��څ�^�����m�ԋgL!�c�U�^����j�x��j�<)Q�0﫞�uˌ}M���ZZϑ�el�D'�`�fS/�0�ٯV��e��>�Dn��v�hn�+e��~-�z��~��Sx5NS�0f�Ұ�Y0�����3Z�S0�j���<�|yy�����'��	�����ψ8Q��4�0�X�.���̾y��<��d���TT�T���r�z�����"Yޮ�`��+[=]M?&��3p���V��2��u$�T���*!�2�gċBM���p��Ga�a�z)��=�zP��<���Z�qqvc[oO!ҝ�8ףM&��0���������}_��(i��Wi��[�.)[�~�љ%Ϫ�i֞q�Ή��&�aF0�,��*���85��P���#���!{�JZ�nD���;�5�vS3f���;�i��iن��.�ɷi�u�O�׻t�te�Lĺ�����]K���;����QM��}K��1���P�ú���d�C�6S�!��Q��̴r�+�eL��}]a)ͥ���[���^0�g�͑�<�i��y��Yfa��b%Q�4�K4��Ҫ�cf/5c��M����o�/�$#�S�WO�ڲ��֫/�Q�� ���	(Y�"h��H�|��];�C�S�S$ܹ�ၢ@:S�����@�(�cU�����C6��+�i�ϓT�D�[��4�C�"�2\Taa��?o�ݔ�Xn-��b����q�����\n�"F[���i�����8믟:�K�J0�i��if�1ˉ�ؐ@l�ғ��CI�c��Q�7��	IQ��-���2�,�%��z�[�_2�t.�ʺ�v�P�1֘E/�OI$ ��܇?�6-�����I�o�D�8��$j*�	������Ž9�nm��܂I�}�7�q'���6��x��j�M�d�)�)��5ǵ�0�8p��07�W���l�2���Gή�����a�p��i��9i��~f���0�K1H�λk_^n���U]V�4��$�8~D��	��Hb	��M��	F��&��ff7V�p�������h�fϤ�]��u�ore��|��i��%��aF0�,����=��snh�$�͎_UU�X}:S�������s��0>�Ṁ������:�����x�t��gmr�ҽ]B�[z�,SH]7��P�e��W즆�tkX�5q\5��Ͱ��2.ɭo7���O��'���nXxd;�Q=�?N[mrx���)�5᳧
�`�Ky�e��դ�1�����Ɯmo�?0��G���J AHK�8"tD�0J�0�M<a�h�Y��x�GL�I0��H���Dy�W�D� �%$",O �$	$ �Q'HH�D� DDK0N �pI(�Nt�M<i��&�&	e�bX�"Yd��a�Ĳĳ�J��`�$O	�����	�$	eI	�&	�J�xO	��&	�"aw��z��^x�gn=ꩣ�xP��J����|���â�mk�͒|�Ҁ�BJ��Ň��p�W->�"v��G��<tH/�*Lm��{P�V�y��(y�����r���윥�Hf�K����n3�vH�e����U��>�ֳxL����ʽ��)��e�2���}>ȕ��g>1!~`΢���L��X��8Ʊ�q�_ձ�c_����I����=,W'��~�w�\�s��ff�fn���W33s37wwx���{������s3/s3w�M4�Oi�X�"Q�p�L4�N���UTB�'em�Pхߔ��pFx!D<�8mm�n/�a�4Ɇ�lQlR�o3����m]Z���a��Mg�����t������n�ɺ�^=l��ml��S91K:�~L��?o�+4U-�#Z�l4hM�F)�驯b��G����[4��0�u��q�~|��ub%Q�4�K4����&L��Y�t�r�|UX�a�>���4F��~ჾ�#T��s��2n��M���VZY��C���5��b{����О|��}LLw�3�+,��R��m�u�����	�إ����,7!�{��������D�a������`��w��wxe^nWW"S��m���y�X�"Q�p�L4�K#�5'6��7���w3Q�qZ{����]4�bVUtR�\bFSe����m��Q��7�B&��E���I'��S�Ӳ�A��q�Je4rx�[������J��d{�i9��q��'lm��Ł*���}g�Ed�<�FB�&"��3Z�k3g��=��e0M	�&���<�W�M���{����NC�j�	��-4#߁N�w9������Q9)��U��\6`�<5�%n�����i+�xe��v���;]����}ne�p:n;�0D��"���чi�����r�H�Z�
n�mdF��L>�w4��K~~u�����K�J0�Y��ig��T=IIes3
uփh�L�S73c���=t����pL����U}���{�4������F�E����F��p�!�O�Y�	�=!MυuD�3�J]B�����g浿�z&��"�,7��PG�z�L��i38!$!ì.�֛�;'F8&Cp�����]-�N��-�iҝ��f��4�o�p���m�|��Ϟq�u��>e�<��>�n�I���*�D�2�NC�%�O���N�p�"h��}<c������?/���Z޻e^���fk�"������9q���y3sS��S�>�s~=��ˇL��L7�\�8S4���k5�q�t�T�=JU�A^C�i}�xrt�ҥ8ob!���W� Ӧ�'�?	��ı��?�G���ե����d��-o<UX���V���	��fQ�D�ꪝ~��[r�9��m��.C�J�
w3ݗ2��ާa�Sz���h�!ڍ3������9GД�ƾTg'�?A%;��u�����w�>�y/���h���1^r�v�aH�c.������n�#h�0�����}�;|:$(ᦞ,D��bX�BQ�,�K4��7*�f
(���1�l�\��#V��〉S!��0Z�9�>3�;���f7#�MI���`L�B0��m�e��&Bb���y����`�9��q��n0���b�LYFF��f���F6vM�>bxM���-�����n�kF�է����zKeQ�4jh7?P�5��-V�2a�m^�6ⴴD�'�e�֢#�f���\[1rG㌡�ν�>m�{~��=ӂ�֍��sN�C�4ʕ����{���j�6"2K=6w�?ZZz�"fp�H�O'�,K(J<4xt�����߶�����R���KÅ<�{���{���o��0��)�~�m����n�4�et�!�{m�CB!O��6>��C�|>�/��N&۽b�퉽�+��D�oļ��L3�4�e;��\_���mU�G�(~�}N5M��T���j��M��J:i��`�ibX�BQ�,����қ:Z+��r&R�3.��V"va�Utr'�>�mkջ؉��t04'�#��{6B���-�Hfᦉ��8d)����V?@���Z;�7���[�pLr�o�ʥ�0ؚ���09Z�i��.2���>~ì��e�o���S���0��S͞T��o�{����}��.e��9!��<mV�%7OUct�-��Ӎ��μ�,D�(Æi��Y�ܘ��ĕ�ߪ�>���ts����D��.�<!�_�hG�܇�T��t����>�Z��1�t�hJ'ڈ�$��*SvZ��)�7>B}�{�����aN��ˋiML�5Y"|��u��a�1Oi�������f���V�z%����*�|��Q��ǜei�_0ӫy�P��$AHO	BH�8"X�&t�8X�H�%�i��igD�J$M ��"Q�%D � D�8a`�i:u�uh�Ӭ�2�#H A<@�"P�""&	bQ"A��i�N��4�M,��$D�âX�%��%��	��'K<'��"@��: ��0��:2G�"I"x�$� ��"'(D��%�<"8xp����;S]:AZ��b��}��'�("jdH$Ζ�e��O�;}���<���qѳM�K�N�n�>}�`�
�!E�i���3���$�r,��1�f���g�ȊHv"YZ�mu,��ϼ�:���>%rZr��9I'��`�ĝ��[�R�h9��?G���P#P�®�����(1��)�0P��. �{�ג#:�h6[���A,�*]&��,(�¦
AF�GdiQz�T�t�>y�)���Vc�V@k������x1)�1M+%PW�I�u7��\����RcJ8sw�N�%�P�v.�a,G��ć9����[����>M����
��к�"n*ݘ�ִ����pټ6�?!��85ᴉ%+��%p��P�*���	��nI�x���C���|�.�xj�z� �~z���B�
���k�!yP�c)	+J!�a��	6�	r�<r����?�f�ۛww��~����-���ۻ���[��۽���ޭ�������OY��D��,D�(Æi��Y����=���T��Z16��3K����v�z<C�Խ�"�������R���gјD�ލ�5�u�EK����]�Ym�����""	��e��Q�b1�-�`��&$CFP@�,4_ݹ���UO��Q���z���	��kLf]�~>aH�Z%�Z�(Q�&��2{�kzX�h-��,DJ�$�~ ��c~ڪ�G~���>2-Gph���6Pcm#�;��P�����8���|뾳�E6�m��yŠ�H/����24g}�~0�JQ�>�
	�}8<Ukm�=e�(�i�YG0���RA|�}6m�vk��q�۾�t�?��u��r��~\J\�ySa�W���/a�=�_ԫSg��E���h���!���!�z�2�[k��\�#JҗS��;�y��8��Ռ���~�f�չ�G�:tO	�<X�&�ib%	G���>:o�^Ū
�*V(��z0��U��'�!�}�)�?NC�%��1�=>��=��<�SG��-L80��A���3����wL�P�}�"��A6&���.6Ŀ,ku�G]���,�<^�	�g��!������=��[,4S�'%��w�oN�D��2�Ů\���<n�a��6��o��:�8�:��_8��<�wH�J�X�K��x������x;>��ґZy��DG�ޓnq:�:q��'_��b�>�>Gʡ������!����0( �֐ay��R		z�虽�p�;�g9W��Z)�罹#ۥ�^gru���~�֕���>;6nO!�U���'B��ɸ����o�m�m)t��[����ȣ�%�xO�&�ib%	G̾q�y�~3�a��rL勹>�Ub!��w�lMM��p�٣!N	�~㇊7y�@�O)��۫t4�ӓ!f�'��?	��0�af�t��-��o�#(��f�����N��	Ļ,3��+�yo�$�3�3i�h�|�K]DDG��ה���8a�o��
tس����M0��0�4�K(J0å�if��I*�P���t�`i��.X�v�l5�ö]_,�ܩ�cJ��E��#�\[d|�¸&+4�Iok1fkb�l�[-�����z�?lDp��bI9�Ŋ1���S~�1<���kc{mΝ�gk�FPO<(����|6e�KSa=;F�xz~�6e�ܯۗy~mn#����G�a�r	��t���^�ΟCR��>��it���8����zm�-�Z�ַ��2�9N3L�ǟ�������:~�2ȎɠВI��./~1).�s�G�/�Y�͉� ��g�u�Tn��0��bh��4�P�a�K>>:|t�U^(�k�*�D�i�f�`τО�v۲��gC�&Q�]]��}'&2e��s���s��]	�)��~t�m�����W�4p#��G���`���9�Fɷ"�n񋵰�~�4�Rߞe�X4��mb���i�rDO�2we4l�������/O�L��Ϝi��X�&�i�D�(��i��X�gci����`<_n%i}MO&���=�yJV��<7:j�4x%"{'2hM��畻������`�)��������؉����y�wDGt͙vݶ���mp��<����	�MjO�#��#�=X�)��(����:��st�ˆ�Q*&��;N�5'�/�J{We�]e�qםyǛy�a��y�qq%uk^������b����I���<�Ή���������h��f���ݺ�oi��Y�z~Ќ��L���N���}T)��R���?|�H�=?ax�ot�l�e�r�����bp�6lMB�<?5&���r���ԃ=�����-r6N6�r�g��/]��^��[i��q����x�(J0å�if���"$���OW*A��E����b��m�L�XK,f��6��/�E��m[^����$��;��q��$��O�3]���Kw�\�e��m���9���U�#pZ�}p���R���H�n$�����<W�y�Gƹ9}��[�0�Tաq�Lf�b�����|7F��߻�fg��o��Fp�&`��2|l��тp�I��ޜ֦�����O1ZDe�v�e����IóO�)��M���pn6-�ܹ������L�f=�9�y�a�3�8Q9�Wǌ(�gK�D�<h�%a��4�K/�v~��;�����L�P���Ϙ����+��z	�BQ5���L���o�]>��;]�?vO�����k���n�Iu�m6�S�i%5\{��.���sX����~)h�O!���n�Z1�;s���:-�g���
U�z\�����N�Q<1򭻕�F�o�Ө��q�^GY`�BI� I:%	"'D��b`��b!8X�H�%�bx�GL:'M8Q���F�i�M��H�A"�	'�D�DK(]q֑ӧGV��:ɓ,�pA�#�	"%�""`��A��i�ƚY��&`����	b`�`�%�`�Ibt��x�"$���'�Έ�Y�:A��$tNI@�YB	�:"%�X����Ç�7�g���[K�[Y�[%W��5����[�i�.>.�d�4ӄ�����/�2��2�ج{��s�a(��6� a樳��k4�i�y���3����(�ya��v��ئ,/ea*��8���7��p$�{}R��ؒp�!��d�) O�����N��[I�O2H�|7�B��(W�����#:H�'�S�\�����{�w�(�_a�#��E�ڰ.Ȟ,��`�1��?�ʥZ{�������������������7ww{{��������ۻ�t�K,�KD�M<h�%a���,��""9�<���y94t�:[�	�)�����VQ�&���m������Ͳȟ���u�&���s3��a�~N()ݘ# �'qxhО,cN����m����ܱ�t�5rKZ%#�y)�Df��5Zc�˯���F,��4K4�ƉBQ�0M:|vl�:`��������UX��>��e�70��\�8%�z��S�(���	��6��0֌sY�k\��+�IBZ_t�=�Y�O��E}�^�Dl��MwɆ�/�>�!�<>�N�b@��d�	�9�{M̆��<�����:pO�D�t���٥c�&�yy=�ky߫|'���Q�w��L<`�&�f�x�(J0æ	��Y���t{O*fj�ȓ���� $�H,����[���
�	��[^˄ ���I�@`('�o���籄�����j9��c͙�s�V"5���}��s:}���.0��L$�r�N�!�W�{�q�y�Z����p����Dٹ���ޢ-�U��O���`T�|k�wT���-�NS�)����1���ѱ<�[�9��Q4y;6SBd7;
hО���`�:uMMC�ؙ���˙�c���ֱ��{�Ss�K�O�������s'g���N6l��fh�i�M4�(��&�idK���210�����$��"O|�GGD��w��i�PM����(,_iH�U�b!L�Um��3��g�����ngӇ�n|(�<�o'�Q7<3X��Q�/�i��S����jJ'5�E�J $��O_R{M��'��Ð��S�Sbs&Nтv��j6����3����t�>�=��l-x�~��[ͺ�>|�<�P�a�LK4��%�RIi�V"v,�Jy�S�vh��um�0��y��#�ͳŷMo�u�I�\�o|N�Yc��Z��[�N�6�1�`�'��!Ð"">�ɺ��)�\����	�C�����N��pJ~��=&�D��m%T����-�����`�Y��4҄�:`�4��'������U ����U�Hyi*�*�N����};���OD<�myxRtM���2���n��M�,���Jt�3�hXn���ҝDg�&�a<`TT�a��}���72`Q0�wI�=���y�{�u�K\�<;�i�8'N��A?s����p�O�>�hy4w��DZ6�m�3}�ש��z��Qm��p�J4Oa�af�t�J�(����4y-#�H���E�3JƱ�q����"�0J,%R)�?�ԾO%r�qZ@f;)� �)�n��+�X�#�%��Ki���.�3�V"k�}��{��4|\�E�n�m��F���>߼�!G���{�O���h�孝ki�U���]�������Y�9��70�Y�d)��w�����I����ɂ}�o�D�_i�V�>=sN����~m��ɐ8x|I&��eˉ�����<��:�S7O�V__�ů��r�xv�.�1d�:��Nw|�ڪsX�baZ<���ç�h���i�M(J0æ	�O���?%P�+�T��IP��*"#d�f.qUa�).�wda�[�vu�����T�C��k�?\�u�3����p��j1O�������1W3K>���>���z�4�����uW+��
���F�t�O1hz��o�P�,���;MS�ˈp�0��S�:�V��������aό8h�%�i�af�e�u�Ϛ|�o<�j�R�or���a_y@t�Y55Vx�><+�z$�%1V����sD���ޒFh�}�����5�����u�5��˭���r�.j����F!�G$��^䑖U�{�ĈJu+a�3���8��iQT�>�zY�J]C.���Z���1Ř0�q�r�Gy��y�_8�̼����O�m�a�&!r�I^�\<�V
�SL**�&��m�g xR��5��t��N�a��`=�˘�?P�k̸3)%�X����Y��L��>�"׹����<����s.�L�:��v�~u�ɧɝx�W~)��h�ym��Nk.p�T�=�z{�+~�#�Ɩ�./<�d�{�'��b�?y�տK۔ҖW�*��Q�f͛�ͽ������Ϳ�����{99'qÇ�6f6tFٸ�#��`��u�7�#��Ya�,��R	HD"��JBD�h�!l��H���dH�D�"ȱ,�DAd(��&����!dDYі��"dD,�Ȣ"��B,���"A�h����dMD�dDM��DY!E��"Ȉ��E����h����Ț,��m��-�dB-"b5�4[D�mE�M�h��mE�MDȶDE�5�",D%�id�Ki-�Ki�M-��B[L�d�Y&�HI��&�m"Y!-���2Y&�m$��d�d��7n6�I-��H�H�L�$�D��d����$�Ii%�ii%�k"�H��%�$�,�,�[I,�%��dY$�L�ȴ�Y$��bd���Iki&[I��4�,�,�,L�bID�D��,��m&�I��K&�I#K%��%�&�$%�id�ZD�d��$��Id�dȖH��I-���L��Y-��%�$�L��&�H�H��I��Ĵ�ZM,�-�L��H��%���%��H��%���4�M1bI4�D��m-�L�I�H�I"D�I$��%�iI�K�[K%��H�L��[$���f�HL�"[Ki4���I����im&����Kibd%�ibM-�%�bBe��[HKK4�Ki	dɥ�Ě[I��Ą�>7	���d�,K$�ɓKI����Ki�L��[I-��	m&�ɖ%�B[K4��Ki	l�bM,�ı!&�ĉd�%�ĉm,H�K"[H�%��A-��4�ib)%�E���8��I�q���5��$md�&k&i$�h"	6�A&k&iYI&�-6�3Y Y6�f�֙#k&iZF�A!#kF�m�3���7�!�M��e�ڄ�ֱ��a5��YJA)�"E�,�3��dH�DE��4DYDE��M�p9dMDE�Z-�[Y��mȈ��D��9C�""�DB$[DE�,�gDE�4YD���9F�"�"&DE�[D���dM""�DYE�#�8Ȉ�H���"�K.8n#�8E�DY,��DD#DZ$H�,���DE�D��"��,��Ȉ�"-�"�h�h��nK8$Y,��4[D"�",���X��ȱ�b,E��E�"Ȉ�&E���h������[E���m�"h�dH�",��:!��"DȐ�4E�E�HZ",�E�h�,D�4X�F�!""h�D�m�#D["ۦ�E�DY��D�"�&�"dDZ5�H���"m$[F��$MD���dh�h��b"-�h�"5��mD�h��k9�8"�"-�E�DYȚ,��&BE��Y,��"E� �DY� �DYDD�"F�!dDYE��"�P�,��!dDB",��#M�&�DE�#H�$Y-"C���DE�DY�,�4YDD!h��-�h��,���mE�"�i��,D!dX�E�H�""ȍ��""Ѣ-�E��dH�-�#Y,��DE�m,�m,�h��&�h���E�Y�2",��h���h��"-�h�-�DYE�DX��4[DѬE�����dX���"5�����,E�����--�d[D�#DZ",��"E���D�dY	D��"�dD,�dH��H�$Z$YDȚ,��ȄYE�q""�Z��F���"Ȉ�$&�hY�dH�m"�"--�"�4k""�h��$Z"4Ȑ�H�DY"5�E�h�dHY�dH�H�$,�#Ds�4H�$Z$Z-�Z$Y�D�DE���$H�$Z"&D�h��$[DE�"�,�h��$Z,E�"Ѣ,��DE�4-�h��4["�ME�-�h��E���E��Dh�4h�"d[E��",�����l�h����b&E�h�h��h�"h�E�Ћ2,�m,������m���p����u�Λ�q��u�c�?vy��6fm�F͵��U[:CÌ��/?Ï����;{=]�w��g���џ�=ng���zw��������8��i�76�[�'4�vyt����vxv<\|7��˧ɹq�s���'���t������;���^��{��{��͛6o�g���q�������M�?3��v�:�lٿ�q2D%����͛����N��~������7��8o�[~9�չ�x�n�����֝��}Lϛ���l٣כ�}|?��H��C�mɾxfzv~������nm3Y�Y�g�w3���8�3�gk�9�8�f���׵ݎ������Lt����ym�9Κܩh�z:�K�纸-�\m���m�a�km�k�z�q��kc�f��(�Uk��UY��)x.�s�ǣ����=��ϭ���Ŭw���7Tf�$l(��Q#l�F�D�m��m����'�������M�έ�w�vvy���fp[�ݼ��zm��of�?�������O���~���뽞셛6l�g���r����W���}�{���v#��������y�s7�G�������>S�xg�Χ��[�e�����f��C�V>������n���7��f�c���v߳��'�<}����w;���|Owc8��ޝ8�a�i:>�f͛�Ok~��m�/�W��>�-��#�;�kpy�=�wk��Ⱥ�3�F>��\1�n��n=Yj��䫖�s�M��[����n6#G!��=���>^��|��n��97&����8���f��c�� w�� I��4d'��a7D]�k?cv�f���Sw{*�/��;�^�f۳یٳz�_k�o�6��g��y�\1�?�������wV~���9�>9���|���~�z7��{������ۏ�9d��7���V�y���f͛7��<vg�2&�����o�3f��owS�{�_���ø�6���<�S���<M۾?bv�Өv�4��-$���}���E�%\�:�Ltkɾ���G/������6��3����3y�tg'��|͹:�r����]q�6i����ͷ�]�8�8�~z�f�o��rg�h��ލ�o��x�wnxf�;rc������6�ӻV�7���o/����7�7o>��|��gk�����~n���Q��f`�%�]1��:o����_/^�c�{^���N7͕�ל�#F��/�_��]��B@R��