BZh91AY&SY3�s���ߔpy����߰����  a> �            � G4$(   
 U 
 �P �������65�kka�x����|  �A@�  }g�����ن燇�x]{nm�ݞ��މw��mPʹn��>�p^�}y'^�������ݢ����%\���R�q�[�H�V�����R�֊5p� ^ ��J��aM��U=�U�k^3.�QU]�o�/g�@�-��F�V�R9�8�-�^�f�u�K��8Ol�ѥ
����a�x= B8�K����UK�����{�ǽ�=ܴ�l�7��� y
�7]�������L�7�q�v�xz��n����6�
pC�U� �N�ک�[�3�S�{6&{�[�����Ѻ�8(Wq�b�w^����t��8�nѽ�{�^�E�������ph��i��`�y<��;���6���p�{:�v����8�\��[��(�u��G�sw9(��M��pz��ى�L�7Ǯ�                  �  JU?@5)T���{T14چ0L�L0&�5?B"IT�4�`� � �O"���    L@   ��MJd	��z�b���FSU�51�4��G��m4����@U4�b�� 4F��A���� y��TYI+QF���L�:7��N5屶lݎ�������n�ٌg��oS7��i�ˎ>����clٿ��͜��_������o���uz?�����9G����������f����K.8q�+�պ6m�7U�y43���UUUW����l��7}��׷�>~_����{���g��ˎ\�C3����;V�Y��F�P�	�p�b�Fy�0R��$�dq�H`���L0e4�����d=P�Q�t|�#8udP��|ϙ!�D1ћ�q��"b�쑔�9�I$�Ʌ�fS����*0���Z��I�� ��e�r�1�����:\*8f��!�Uq��&aڵ҉4�dA��)��P�*e�����C1�0�dA��v��Tp�TQ�HB,+蘈&�r��CqE;����;��/b$f�.2�)�@�(����	�Imɩպ�$���d�:��ܓōB���"M��jcj�+D�D�)(���kb{�TbUmE��2[.�{w'Hv\����:A끲�M|��
S�B&+Lc!3��Q��ˍ�#���c�D{�g�H(z$�C��d�=Bz�4�XA����M��G�e!�Q���I�3�P�(��'�c6���?�P�)�ꏢLf�D|�C���7��$\�ZY5���H)����X���(�*�z��wʄd&!�چ3�v�N';Q�,}�0f��4������ϟ�T2F5QE?�,e�P�ͨ�XC�p�ҋ���������&����I}�-���$2G	���d��3!1�Ҝ�XͅD�8L��S0��,�XA��r���#��"��m@�����t�`e���2�_R�h�z��1���3�(p��f�1�2�z�i62ጢ����l������Be
� ���b$� f�L�erMj_+$�"X�@��c�����E�k>VD��q
�N�3�3p���΅g�J;
dS�|algB\�_qƾ��k�6*��	&�?�t��BE�����c���z�&��d�JBk�=T1�����1�c�%�I$�Hbd�p�CY)I#�L��3�*�}
1�c8gV����<"í|���U=m* e)"2MQ2������x��+\)<@��(�N"�)��3�-�(,cԜ��
X�a1�X�d�3�U�iic$\ȲpT��0`�h�1��I$c���|���	��W8\H��h392���+/��A$˅ӄ`��r����D��U
`�!1��e��qN�J�,fUBDX��p��!��f��4�~f�JX���!�_8Y�	�%.�����%$_�f}m+�,�i3Ř3B�K,�%C �"�&�-p�a�}��ʃ�H����@�r�ZI#8r$�(q����i���p��ZA�ӅBl+I:�T2F=�L��簤f��qI�d&H�+R(LK�y�I2F7P���r�L�����g%�L�.��
M��$�H��"�U�C�"�2Fc�PY����Be�u8\KJD�/��S	�c���dBm.�	�Y-��I	2F1��z�}
(4���.4�����j!|�,�&;J�9�ORsИ�@̧�4�p�a�8�)1�2.�f�"�l8X���2E)��5ЙCkH�&p�f��-,��`�oqa]�XΒ>.�K*D�Lf�!�Aj@�i�z�����D4�Lc��oq�qd�"����"Mf�2R�ԟ�"�;����}��2�
�[	�r���.Y\�0��L�3��Li��6+be�X�$��p�ӍzDk!q�2���`�����"�s�\k� ߬�����	�d�f��Lt($��9_0̂>k���<Zٺ��t׃�dxh�u�F�t�3
9*��VX�1�S��� �Le��3	b_1ډ��&2M���!@�6�ƺ� �Le|�Ď������H�K)|�2f�1�O�f�V�dr���c�����q���i=L�
��1����$�1�
� frђ3�B��v�c����D��`�"0�2���gJ��1�F#	�r�4�!`�_?�n2�, ���C$f�T21!��(c�ќs�1�W),��a��lL���^�3ʌ�(a?� �4�C,r���Ti�4��(�Hͨ�I.1�3(c(f�c,C)b�c_"�V[I31��P����c,1�s�C�3���1걌T�@�8B�Lќ�C,���aT1�t��9ʌDڑ��3Z�)�P�|�~ߓ1�PY4�����C�=�<�9G�;�j ���*#�mG!�nTag8�06�	$d�P�bf�!��Ƹ��G�3ǩxӏV���r�.qa2��w�0z��)�DC���ڌ(��ɖ2�(f��p�52��.��Qc0u���7�
b|II2Ȣ����&=q1��8�Z<�J��=qw�I�C*ձx�1�I��KH;�4��R�ǩ����	/��"1$�&�%�4��b"U��qM�@�x��Q���R��h��$�C��󈁭v��WN��N�� �^���%N�|ev��T:�F��N�et:x�4h��b>t�;L��S�icJ���%.0fR�����f��[��Li,�t$anP�t��X�(�:���j��j0��c8mg&Y��Ɍr��IX��9P�>L�_�D8Ld;Q1��1��x��6����G�bmF2�(c֬cB����KeQD�4�C$e6�3\�c�� cވf�qe%]JO1�|�d��u�����Qd�QB$&&2�{c0��A��QD�c��0g<��$��ʇP�D1�q�>��@�7eC�4w�>m|�!��[��:woI�:w�UgOB%��~H	��O����8��_��G�4y����~#���	K�k�^���^�3:_�vM���9Y@����d���j����Dc큃����f䛲v�J�F�`L.:6���w+J~*L�����ެS����"���BGO�����V7e��4��wȜN}������n��l�K�w0��wD��G�l*��~2�2�·|mAY$�m����Y�(l��/��ƥ������.�aD*��+������Wo��dl�������sQ�mL�D��-��*R6	�]y~�w,O�{�z�t��hm;�t�۽̆�tz;gE�\Q�4
�� �
�\0��F��0����aFk����w!���Ҳ���e�ru+b�$��wW�a1�i�ȯz���ܘsH��������4�w�1a  �7� 9������Ne�>̆�dj��~�->�m�FA��{��Tt6t7��Ӎ����}�Vt���8(d6�����~��2A��~��6l$>�)С�ֱ��89~ƺ�o��|�������bd�X�㳥������$�oO�i��ꘈ�+}�5i��2S1~�n��oN�߿}C߾g��1����*��>ݛ6��$���;Zv�;����Ս��gn��Zo3f3S�6Ͳ+�L[�"���}�n�y����9����^��;I�83q͓���@�C�e���߱��̒S��fW����e�����ޭp=Nәj%�$9,��	<�c���yu��1��\K[1nP����%oײ����$�s'��,�-���}!�^�U0n
���j�:�%^���0�257JL�<����ij��J�s���\�/��u�WHt��� ��F��M-�L�YN,X�2Pj���b[��{����:9���,��ufa&z�Hͅ�T�(��88�e'nN�F�_�����V�"a�# �|w^����]<w�%7ZU�j�����6�,�`�in��6U�+��i �L���c�S/�qcQ�5<�9�Y�ۙ�SG���w�z���$��}7X��\gLƩ� �?	F�Xu�U���?{������RF%�����~�LX�GŻ��-�n]70L_���^�d�'�E�ͨX����-������d�'d���n��Í=pV�IWH��zqznk�$�f�NRQ��B�rf:��YQ)(&%t�p�+ayV=����_+�"��0a��֫&a�
�V�v��nQ���ı���
i�Kf�.���s~�v|���	H����ޘ��3C��C\��t��ɶ��s��qg��b��A\���-� ^ί�Q��=�Z9��i��{�_{aN73s�Y���|>*&���*0�:q�|P�$Ϥ�ݝ;r����C��*b�����]���rA�,�weٽ�9נ�$TM�g�&�6B�=1���gl������V�R�s�:��/q���l������3<m�T��"-5=\E��yyi\T��e�~���tO�Bx >N��H4��qg���[ǒ�Wn�ϳq�kp�f��d�����w��ou������s$z@���F��\��<�ޮ���y��V����zw�F $0�;q̛�I9�vXU�:�����}5G?j�p0��;�<ӫ�=�CQ`��^)|�т�R�5\r`W0�����U���ßG8G}~��Nq[��a�ϧ���<��. f�ش[��_t��}�(v@ �l��Ӌ@5�FZ�vw�s7%���yT�N�Ft_;����kg�S<܄9�Ԧ�!�������|?h��$L�� �h���'l���(�I>�z���\��~������[<�qx�������%����ϳ���O�Z.��� 9:9��T�1�3�sX��~}�n�+��}^A�2E�k�Q����nJ�Q�>=�q;l�H��,�d ˙��>��:3_�=yfnI�>�x�dX�fwS[��]���v��&��vS޹� w������z��I��g� ���3{���}��U��^n���u��%�(�Us�&L�F%�e���<�̚�s0��[Rqd�e���|�y���#�q|���Ftn��@�ɮ�{9w
+��E8�v�=j7fw�r#Z[��K1���������� �U���Ku�{��w�l�ٷ ���0��HG/����v���Dg�D�:x��6G�����1�O\ �! x&�R����w�ߝ(���s��������Hi��c�!�a����i������K<��/��g�+�}ss������(��I56�j�]�\��t�`Q��'�����}!����� 0��io��>�l�_sR��G��o�����k57�ft�������os�{�����{�s[ �Էuɗ3!c���� ��_EI˞0���t��ta��� � ��}� Pٚ�u�@Ǘ ��<( ��\�<��� ,��,���>߲��7#��fj�/M�Qi����K��d��9���fq�7 |��ˣy ���N��������}�^��Yod�M��ͿD�;��W^��9U� vH
�Y������c4����w�w'�#�{T���v/v�,z��6����a������*їw��6擌����^������wZ�>��6� ��ʴ�f��2>m�Ow���>d .�+��0�D�2i=�Y�gۻ����|����~���'Lx�d��֮���Ӛ`�[V~�~ž]o72\��sY��a�Ѕ�!��]�זYO��v�׃��}��{$M��������F��  � ���_����I��ݹz�V��]���̻�;R�+���'��ux�(�� ��x�b�8���b}�$���I�lU�=5�:_#Q� LFw��gd�]�Vx�Y�eU���%��H�{��2IBHh�W#�������d�d��P���n8�vt`A��PL;;�4���w�g��8n�����w]����������$k��Q���Y��@�����e���Gvz������]���?���a&G���2L?���9�}8Q�$Jٔ�"�n�bӄ͘�-�:�eNr���0�q�k[�],�.ms��3cd+��n��u-�%˱�c���0�as`Sh&K�X��f�e�V�u����h1�\�1����x��*{�������=�z�e�P��ūăi��XrTC�iaN,���ߤ������F��R�B]1���zrH��{'�&|$!�I��h��9�{�l{ieJǊ]m��h��!�*|�eG� ��m`�˭�)��=��N�"x]q!��q�B�Um��>	�GX�mOW�/�����xJD�e��cS�����#�.᾵,|���%$�u&�;R�L�ک��J� �(ėM$�"��d3VY�g%C�7������8���ހO�;V.,e,'V��
y%�Kִ"�n	+.�m�|d���۩�ͨ�w���!c=vԁ��탬Wє�X�u,k/Kv@�4����]ɩv)���bң[s���,8�-�Ȉ�16��[�Yo�R��E�`�8nQE���xqx� Ě9fR�%�3[td�i �&�^N�J��F��T{l�w,���d��/Az��0-j�Le{-StѦ�Wb&/!y �C�hr�EH	�P����E��"b��GF�%��2,�,P�pI8��A"DOJq���FP����6�q�K�k���m5X��-�J�%�K�T����0B�u4�0	l��L����ɤԍ��j�\O=NЮ��������	���.�(�k�ed��Y�sCZ)Ņ@�^*"bΏ�1y�.�p��40�7my:�Մ��
k�l�
�JD�gZY1D��8�N�YW0���t�"�TD�vz�+�!)g��t�a`��`K<�d�=l�A�3�DD���>���#z鍡ă����g��w{v&Խ&;{K�N�E�&x*6�m�T|rEӜ��ݼ5ɶ�����i)q�mV��K��cDLM�q�J���X����6\�[J�[j4h��)hDE��@����a��d^��P� AD�j�5^4ֻּf��/�*��#��ͯZr��O��/OO�OO���y3�7�w�\[��|��?���7��s���ߢ5��6��e�kq8m��������O���_����:�6�6�6����m�M���ܶ�v�tۆ�m�i���ܶ�v�t�6�n�n[m�m6�m�m��m6�˻���z��m���������31M��6��)����Lj�j��H1χ���ý�orۆ�m�nm�km��cm��-�ݶ�6��o�m���m���m����m������t�fe�6۶ۖ�oM����	 ���|�m��r�m�nm���-��6�m�m�m��������m��1��m�M��z�6�v�t�m�m�m����or�n�m�m�}�RJ(�T��)�{�ǽ��=���1�۶ۦ�n�n�m�m�m�m���m��m�v�6ܶ�xۆ�m�m��cm�޷��o�m��a������m���m���$		|%�)�[:'�X��l��6�V��^o?c{q�6h�Z����^����(zsg��χ��ur��������#8�1�2�Ŕ3Fp�4fќ3�4gac,B�3F2�c0�GX��.$d@�|���	�,e��Í3�p��4�3`���D��$Cb8��e�1�@���8c4g8f��`�0јY(�1�1�f�3H ��!�1�1�3�3�3I0`�!�!�L���(�Ӯ�:�:�V�:1�c9��@��a'����j�����/߅݋�V�d�9Q qIl���d2�q-�͹ұ+)�э��D���0��I�h2�6ۘh�	�'�R�o����+H�|���i ҨAJR���a�[�]�Y
.k-��q5��e��L�qjc�Ϋ�k�(mkmu�H�mE���� ˝�F���lrC\a[��f��h�4vf��lZ�>��_Z\YR8l�5����+�9�0D13����O{<�d��nF�n�aɳ5�Z�h7[tU��5qe#*�Q�f��#��V�o�عkjY����4��, Evqŋ��E-&-�K���֍����j[��E8�����dc�J�E�[��Ү�kY�v���bk��&V�C��nkte��P�c��ڬ�	�X�%�	�f�X Ku���Z�S�I���ke~�z6F����[Oj72���f�P������5\X'��X�l(+U����m���5�Y��u �+[�T�[b*Y��ڭ;j�q(PQ�Ae!f��Hd��1[U�47,ͽ��� ˙����{V�\ᴷJn24�i��v��΂�W`���]p�X�T�Yl��ЬUf�n+V�xt�B���X�Z�kc�V��J@P�6�cIc	`ѽ�5�f����hUC�{U&nŶ�"B�O��x��=�b[��Ín�^K��-�)[���$"D�
cD�A3�����!�(ٝVWE%�d�-�����ke�ӬaL䘍9�LK�d3��v��1�[CVm�u�f9����)�j�6�Xs��a�k��ċ؏�=���"ȥUEbr!�FjT�L�K
[u�nԹ�lx��5e�V�M\iq�����޻�%ٺ�(�/o�(�d��l�b�l�Κ���^kIB;�ݭ҄����v��-�:�qt&�b[i5o�m�T��,7dn,fb�M����s�[b�u�]�A�6Ըŕ3aQ٨�ɋ�[Y��i���J�&t�ZtX�GV ��X�B']���)%Ĭ���-Y��Mc�&4d�i/2�,�M6c6����*X2���`k �=�\���/���K�:
[�[��J]�ai��jXZ=������K�ݫ��ܨY���l�/�|E}�2��0Ј���^�=�j:���|||���7��o��>���㻵�{��o������~^���ǻ�>��;�_���6�������|P��8�ƈ��8gӍ�4��1����M��nq2��Z��(:������-.��m���u��q�Fi�e�U�����H�/�Mj$�-�5;Wi�%��6SW.kh@�:l�.�ei�]pB[Z�lfhƴ2��-ش���5����uҍ�mM���[+);J�I��s&�JP�j����{�],�5�n+H��maY`ia��cc�1��Si�%v��f�i@�12�̯[�"p^x��F�f�5�I��l1H][F+�4UL�J.�H�*��
X�ǈh'*-�U�'!L��B��� 2�(D*ՌR����RE��'�}t�.����d�{�a)�l��IL�F閏fT���4n���u_4���.�Ir�!�H*��=�&�`��bD�聠��u��!v�/���*���"s���9V�/�T[̗V�1ܱ���Ym�[y�������4�F3�0fds��Ȟ��E�|8�4��\����E�U���.K�
�BQCb>4p�g����~��t��c�Z�V�>�ݫf��YϾ�N���u<��i����E�,Z�۵_UuX�e�F)�WX]5��+w��19����e�Fh���4�F3�0fd,�"���J��LWYa�]˺����}�4��G���*CBF�����E�j���eC�e���[7G�l�%��^�[`��ބ����#.�8��h�х���yȒ�����U�M��{U'W�ʍ�O:��<ۆ�u�\u�3�0fd�ܫF)�rX�
/*�7+G0��Nh�tp�s<�	vN��sQ�f��I"B�'G�=��3Yy��RjNW��TÔ�'��o���T�����ϙ|�)2�TJ��>w���&�Y�M1����]1LS���u�\e�-�qf�`�3�p�8ь�L���}�b��#�T�:5�����a�+:4kgv�kڰ�ڭ���T|aҕ��,>c�J�,m�&��6�4��I&W`�s� ���J���f��2�,�,��slv�#dE)b�e�S���<�����q�a��r�������٫j��+��$-�l��K�Ӕj�;Fp|�j�ѕ^�l���d����Q����J�'�*4XM� ���h�9���ux�\�mn1WP�w#�,��_}��MPf����F�7���t�K��d�p��>n���:0Ѫ��@�ٔ_���{���J��,��q�<3�p�8ь�L��JȅC ��uX�{|m�A�}Sh�Ͻ}(YvnB�V�6�2�_m@g����^���i Ӎ}LB|Ҿ4Xl<Ú�2��z����o��y�q\����+�l��sX���z�(�дj��W����x�"�U�������k�|��0�x��ֲ��>���'SNI+I�N}�E��A���88{��.{k-ٲ� ���,�N<`�3�p�8ь�L�7Ws��~>@�E�M���t��}����m�I9�0��Qf�0	�t�-�ƨd��n�ثUa��<��ieK��O�N6ku�^�s��y�ߩ���ő�#�#ܮ6�}٬Nd˭{��x�a��5D�Q+}�+)`�W�> ��2	(�a���8gh�q�N�뫬v9��Kld�;O���V�Df���W����E\$��͇1.W`Î�*�gSME	&%'�Y��񍲉�F�W���2Ö z���!5}.Cz���tB�}�/+�|��r�q�ٺq*-�rzH�1m�e�M��F���6�'�<q���8�3�,e��|���z�^C~�h�Ȍb�c�y�4ɬ��}����ޙ> ��lY�����M���f��;�l��͌`'	t��W	��I��[����
���K�Yp�U�n����
��\��s��e%׬�JK6��Dx1��3����N:�������I������c��)�&Y��))��w0����OH@IF�R�*�����K���Q}���֤�5�U�X���URz$����nBÕڐ��hꉇ��c�,�Ğ���fx����g�p�Ɩ2�1�P��& ��u�.ת�ɨ��[���b�=N>g�v����З�Eٺ7FP��-ֺ�eL�8ٟa'��2����ƞ@-��|n�]\��k�J�X4�q^�z�.Z8˨w����橭���p�K��V�T�e�)��Gv�?�-�m��������u}y~u~GS�����_ɗ��?#��:��N8�1G�dq-2�&�I�<Q�L�8I�#��dx^)4�������=,���MB�EE'��n<ƞ^�[ͯͼǟ/��	%�2xd1xdl&x�	x�P�'�^}%���a���Ǯy��y�����험��4�m�yxL�����m���u~qo'�/�c����y��y4���z���c��ci���c�%���i�c̯�5��1<�:�N&^/��ȿ#�]��䌗����--<���������ߒ�a~b���ȿ'���z>��Z�������?œK�����{����k�m�P�z7"�x�_x������b��*�V�C�s���}���v�2g��u+f��P��d�NT3|�5WF�}����&wô�J(����Ͼ{��oww��wO?/{����w}���b���{���ww{Ƿ����v���!qGaǌ<m�\u�^uמy��<��W�5TDD	M��4h�Q~/�Ϊ�D-UĪ���Vf��DDJ+�՚��Y�Je���'^6�ɝ�΋m$��14(gm���gv��iܦ���U���]��p���i+� m(�J��_R)�E�=�W�%!�e�j�A�{�.����C���Քe���S|�%Ui
w�Oԑ�Y_3Vm*��EaDj�>��a^JVwKV�ZE0���,D�WŕA�4%�B�(�	<3M0����~<p���ǥ��t�1M�����7BW]6�v���L��3�;�8nJ����+b&u��-j{v�Y{�VOn�����X��`'Ԇi���n��l����B��@�J���mDv��)_�|©�}7����5GP�Dvꪴ�_�tgL0z���r��(Dj�Ns��5���˽+���%���&�B��(�Q�u�Ⱦ~�}�iQۥy
�0���� �Um���Ֆ�˗g8w-�&��i�[��n�nR����u���ߍ��뎸c8��,���+�y
QC����� �,_bk6L!�Z�l�7[Ĥ�G���%ܯ�{�/x�A`��{�������&R��Xi�6�a�#�aqLe!4�׷�3��m�;Z�R��v;[m7�<{�� B!|�[>��±%ƻ.CJ &�tft��Xg7XJ�%f��0�BЋ�"5��K�S�jYpGYe�.M��7�uY�T+�SLUy�����|�Z5��/Z?�7N4��Ev�)*�Ĵ65F��2���s��d�����L�"�+4�-�mZ�IU��2�d ���%{���)�)_E>B��%W�""1Q]���xB5[�"�6���%�(�#�-[b�Ećr�DE\|�Ol��{��X�*�q4�iZ�-�:c�)]@Eus�������X�G-uWU%ST֓��Q�U��*mlJ$oߒ�5�K�q���<`�`�ǎ�8g�ƒx��u��w�����\����G�!(���J��2��TU�J�!3@��a5�Â"aI[�v���yhN�{��V	�MZ�R�DD���5[ ���̙��n�yQu#�}��",�,�<2�n��*C�R"%�a�˗�Q�F4�(�ԧ�=)ȩ(Ķ�=lO��TKF�D�+VY��c��b]�>R|@�j�ĜE(M�n�&���F�R]|5Y�b���w��`�+u�v]W��+�����"n�T�}IX&�s�#r��@yMWq�2�o͸���x���:�:xt�Ӆ���zB|Tf������}M.�"��4��C�My	���D��D�߲K5��A�����Z���B�$?rO���R���TV�M�v�Y��KU��"%֐P��Tj��5G�Q*8����^��kr[�Қ��=Sߗn�E}�P��_	ޔ|n�=N�L"8^�«̱Jʑ���{�dK�Z�?Nj٥uE1U�U]]��V"aIH�[���T%"]B�F�"JJ�T����J�.\a�j�բ>���9I*����<�>���u��0������~m�6�<�:�1�A��=gt`�s��븈j����K�tZ����1~��佄�W�ozK�>��UQ�,K��+�ԟk��7�2��S�? ��Dc��\�eԈ��MB��l��3~�H��;&��6[&:'u;�k�Y���9.}��{�/"%�^ ��+�$C�ZYU���|�$�J��oݻ��]���J���e�F��(�T�	F�=��u8��js���"+T���)u�#=Yg"���c���UM.�UW��>Z�x�φ�+�<��W���	F�T�.��C4E~u�>��-�-�k��wx�/��Y�)u]af�����ChƩmT���Ո�+~q�ͼ�o�3�p�0c4�Ǌ=�Ώ�"� �)ā@n�"��[�3[U�!6T|�gG��Yc{98���k+��Zz�9��q�8)->D�e)X�[�C�(���j��Kֈn�@�m�8F�3�2*7���Ʀ�1�j��(IX��`T�Y�K��α3����R+woUGQr�"��4Xj����Е�Ee	��Ԫ-�p��EHVR�ha�����hb��s���-l�ݪUG�uOTqs]%RF��e)\���[z�M�6�/�~��!���+8��Q!�C(b��wU�UýK}�%V�Q	2��h��4M'<%yL㗌4��R5��q�k���8�M��J1�R���K���W��e�L���iI*��J��T%V�[<��ş�4�(N8¾�L��{^~�^1L���~����<�o�m���8뎸덺۫y�i�Bf<�=����`�P�n
5YY���&j��C(Y�S��wpb���_�FPcK,�礒"��WU�f��Gy&:���n�)�k�>Y��(�Y�.�Y�uO��=l��>��>5GJh+1�N���c�i���ե�?q8���:I@�
x!��4y�EF�P�nq���L�HH����H�J>�3H�k���ɸ��ұIJ�Գg븼���-QR�_ij�1���Bv�UqM�u(~�I=R0�t]U�Umm8��o�6��u�\u��my弚.�\0���⪢Q�)Q�e�\u��Uy���3T���ڕ8��+�)t�m[���Q�?%SHj��E}�"Us�����N�+T�X��.��V)u*��Dl��aW*���Q�&h�;��K� ��"��Dљie����>y{��7�;�0�����C2����F6�u^|�u�At���i��&�oj���uII��j���%V����-j���;J�"��O����صj��$ j�f�/Ev���̫��R�T"�ۯI)n>��\YqN���6���~`�*��[�^m�_�a���8g�3ǈ<W1e��uU�OOHPk�V�hmo�~�t�ZYyFo
�%?TOhܣbD�%�ƍ_�]l�^dQ�U��L�� o.��y|�۵�m�J��)�b�R�b��.�^֓WA��!�1B�CIG�f�F�JaE���lӈonI?eR��a[�Jn#)ct�U"I^Q�	��D�+f�ذ�ƫ�-��H�O�a�[�=�����������>]:��bWW�d�?����+�3�����x��ǅ���u}y~|�'^_����e��<�z丏B\q�|&Yz#E�a��ye�L�Ǔo/ϗ�_;�z='����|'nH��_�^���&�Zߖ�~H��䷗�cl�ͼN �'�ផC<S<C�F�.-�˴�<�Z������N������Ǘ��<��-痶�c�/ɧ�u:�&_��y����!���x�F�F���#������<�<�qzO2�=s(��\��f<�̼���~O<�N>g����������x��FK�L���Oc��l��HzOHM�_�����Us�by~O=s�1�hz�����A���r}�u�[�u��9S�b8�E����u�3ۨ��a
a�G�C��&��F��I[�Ҭ���'�u�G��;{Soutn�n��3o�(����_������xS�R��Vie��i%�Y]��Z��[��w>���Z��"�&�xWUT㵢�@���6%�#�����z�3�v�6,��ך�����aqz�
������N�t����ō���0�Q�����������M�c1"
T�j��hE�Rg;ڳ��8�5����{^*��`k�* �}�ٕ�ߍX��N��޼Ǎ�Y��k�۸��U��*]ݺ�af'�E�Y�#V:ܮ�7k�o�+E���1I�	|�=��H�氥i�*�5�������X~�Jf��ܮ�)�b�]65��b&�m�b�QD	�ٕm��S]5�F�JjHV�9�,Z�͡�6�t��%��mIv�K�+a�p�kw3�����=b�t�/��4��#��+W�f"����&�'ߺ��PlL�T�6gF��?�={������{�ݦ��6�~�����}��o�������m����(��0�ƞ<x�3�q����/��J�f2AU���ܔ��v������kw[]�WIhJ+�.�����+�_y=���5z�m�ɍ�$ڰ%��RY[l�S����]ٰLv&م;0,ddJh�8`wv��θ�b�R:�-�-�kX�t�qZ''%s2�Ս����JA�fՙ�8k����R�~lOO4/���nnb��`\�)VU�uk��c��	2�S�u�dt2f&��&�ZS3˳VD�*����^��L߀ BK���&����-��peu���K�I����i�[��qå`w��.�i"m�Y�gqM~=�,UtZr��v^�S�im#���]Vi���-k�X�/�����S'_-l6�]aհ���d��Hhh��)�p�(���z�V���R��"!��[�����ϭ�7J��;��0WgƏ�_;�N�i�z���z�Ô��R�Q�*�Jg+-��l;K~J�C��(����W/��Lo\��J��0I�Ů�x�_{D�8��Wj6�ґĔ7D	S�d�2��%Y�,���ώ?6��獼�뎸�N�y�y��v�K��pҪ��ƥ`�r���(K�j��N��p,Ԧ��fGh�b�BP}n�͝�n�፸�~k�.Fi�Pv�,���OS�"T�4�V��/�k�u���ϟ�Z���Q~�W�UC2�+��֦[��^f?�������;U�w����y��`�.��+n0�e��X��kȕk˦+�f궼#�4��]e��K�u#��u�����4�o6����o<�:�6ӧ^yoW�۳$ջ0Ȫ��CI���蝣�U�I���r�Y���,��?1Z}H�H��.���/ �:���_�q}�I����J��=c�\Ň;�:\27}�G����Q�L�Ns��)��+�5�u��&����~čL��M"٪,84cG6]���gM���՗R��v�K�(�!�W�6����Zf���ie�|�ێ�x���:�:�m:u��l�x�c�d��� ӉgeY�iC�˯�L}�k�]>g9�!/�,I��룋"��۲A4�/�ZÓ��F��s��*%�|�9����n���>,5��>�e�����:���j�h�Yu��d֣)w禪��U$;d����z!~*��ט����ኧ��Ϟ��b�ԁ����XJ ^�U��,����RC�J�Y�0���!��٣t��2�î����獼�뎸����|��G���uYN�^M�6�Y�\!E/����G��jb�Vm�f��w�z(�׿w0ȷ�4�[%[��q4ߞ��k��-sd+[�� �8-���?��h`-�XƑK IȜp� g��Z���wz���DUD��CD�.��BH	I���)��9��P���%6�gj2�T{u"0�2�b!u�]�Tf�}`�$!B!���z�\V�if����,I��a��UY�Uf��n��hnB��.��n�Z�M���})�2`�����"�S���W<��0�8Ej�i��E���)�Č��Yk�7GO�D��|��q)�D���j��C��>�Dj5(�~�y+oߤ��&�~a��m��Θ~<p��8����(~���uPV<�ۼ�:���w�M�wS�%�:�7����DR���\8Ƣ�^:���z+wW!Η}��Z��'�{E�
�TL�����m!bx4A�$�Q�4���)��b�mm�q���u1Oے��N1U�"�0Y���N�uG(N���,���N}��I���%���/<l�2E'1w��T��ڲ���*v񥏔j�F���%���)�q�����qfP�睻���eIh��G��4Y���^~y���:m�u�\u��t���K3v�����k����,Ϊ�$<�����iv�b��$�[�NܟUfl�G�>CD������X������aB��t��ȑ�1M7κ�fQ�N�2K��[��U������{Cd�������\�ogR���'�,84��t0��>=�k!�V�n��~H�Ӵ���|�!�a(�Q�Q}��F_(��D:Y�f]�)�Ǥ�#N��O6����o<�3�q���{ꩈS1�eڏl�UTC|:]	�[GG*��,�5�a��:�$M��q�Gi�Ӎ�^��f#q��T�`��$7[�t�ʆ	K�d�'���L5O�u���q�'WQ�s���H��OɆ㔔����O%FP�}V~��J�0�f��3��\��hn�ԥ�IM�R�Chj�N�MW�D��.�O�C$F[f���j+X_�8�O�0�~4a��3�p�0��:zC�a���>�W�5��ԳC2[Q�էv�v1; �F>�_�.��D�>\�@n���VV6̳9�cqj��ۻ} 	6��I�rYi��餴m�n:�9��׵ҭ�3G��ɵ�[�6?1�\���`��Е�<�+��^�gՃk��v���UB9N5Ʃ��m��SԔ��k!�j���X�c�*��֐�#h�%C�U�TȶV�hӶ����h&W�&�mh���_I`{�I[1_<��]V�.E,�;L1#U	U�3�~�CP�H�jk0m�s
GeG��j�jV���P�Wn��0b�Q.\i)���gR�~���J��Zq��~m�:m��p��0c<A�b�U9+�2v�Ui,ϊ�U���Tgǆ�WL�a���ɚr�e��pB�'��(45_�J���s���0�@�<�W�/(�=1�@J�6��EЙE���И�A�^XĔKXlL�s7/r�l&W��bM���>.�<�>0�v]�7b^��j���r��xl�tX��J�ƑWR�J�Tx���5���Oܓ��[P�%G��<��si�f���A�Z�Lm�9s��g�!3��8�	xd3ǥa�L��ǋ�_�/�ח�6��E�y�<�a|y|}s��4������闘�m��ǥh��мC£�*#`P��^����Ύ6h�>% �(�'�������m��������:���ig�b���Q�a�l%��A,�<���������yq��k�1�y���k�y>q~L=s��q���9<������1��������>�k�ˏ=�k��<�nO1��0���<���,Zx�y��/1�ͽ�������a�J�<�-�0����+˭I�����h�$yo-~b���y�����<�=sg��y��<�~av�'�������=��޿{�_��f��cm�����v<ߧ
��юv�w�P6�dED_�����YZx��[�q*P��vI�V�ޱ�v�l�|��\���[M'>�UL�TCQ�I�dt�(��4��/����߿�m������m��������Ͷ��wwww�y��{��8��(�8�8gq�iӮ����$�TEb�J��U���f���(�4V�IElO��ܣUZ7��LV:8y��{BW�p�z	m�ZX���ݸݣ~ ��v�YfLs12�,�O�[��Ί�����\M%�e{.��n�N8'6J	�+>�df�n��rN�0�N�++>F�So�4�Z��Վ���*�!����~0�x������h�,�t��L�<�V�U�j�Mw�-��.�\���O9OTmF��)����PpL��,`�|ʼ��r6�ᆡ�f�j�.f�C0�r�Q�k��S�o�2����Q�%4�v��F�o��M�ME�6�V%�dF��DZ�G�����eJ�&�Q|6&�Ig�C�}�.K��n��GP�#�VӸ?}K����+�kM��R��.�F]��J�ï2���~|��y�\|�m:uז�#��O��z�i3����m����N� ��>�,j��	Ly2�=,F�/����e��e�Z��e�r�K���Iqì� E�]� [)�D!Tp�7+�a�D�1�˓�6��a5�IB�Tml&���h�+b���bv���k�}ωy�e���h8&���(�+�^Q�<�\�e�����a����}.�-�&U�}M�*���~��L�U���gƏ�h�	��'������;}U���L�G-u�Au�ӉB�>��UbC�\5^�(ܢ5X&z[�bH;KYR��Fƍ��{�H�����۴�i����ڗ.e���8�4˯�~u�ߞq�q���^[Ɋ��}�B�����"���j*�#Tk�<ļ��TV��th#CGF�\G<�b�>�YL�����
[�j�g�Y!4�������V�=iK���Kc�'+0G��@X�Pс����&� }W(0I��*aɇM�#�"&��=.�	}=U^|�I���\���\E4�������Yt�pOD:4��f�~>��iG��t�|���?T�afn�y9��F��<�,�����Fx�ǎƌ��bzze���RTҪ�!tѴ�5_�A�8s�Vv�К�5V�j�͒B�4!�&�E��%���0����"|}��[��72jmn.A��_Nn˗m����cL8e8'�,�*�F�u1m�R{H%C��D�U�'�B�Ʈ��ʤ�
ؚ:u\S(��	��'�?%q��1O�r_����m�~Z�]?6㌴�o<��o<��q�0���:��|����~,��c�����/����8^w3����w�����yi9�Y_*�"���q��~b.��V���%?GQ����F	���E��bT���;������2��-�uYʇ%��G�'_[n�z��o%淢��}(h����?B�ո��6E~Jm�f��2�����	E���c4��s�2s�a)��1U�՚Jv��a�찃G'�*�=�G@hC��#��M��lM"��C߆�$�����8�b����.�m�mƞm����ǎ<p�4f0c����Q
���}9�2���ᩂ�1<״*��.��+>�)�cޕ����Gvr�sN[%L�+����֝n,;��9(�EE� x�e��o][| �n����%;��ɐ�=.�Me
g��N�R���<�t�QD�����)�8�]S��%!��.�UJi#��t��n�?}.�!�-M��%��j�����1D�qkq)�@˖�7�Mqmar���8��f�����e*�A�W���T��KS��)�E`�)�a���IZ�D��|����N�F�>1<NNކ�B��%f�!�+x]a��um�)�Db��)mVƗF)��wkb���G���i�q��O8��8јX��C<G�(�awC]��E3J�H�Y���J��(�?!��qx~J>�g�Z�)���%��2�#�)���(М�M:B�&�br��%+���ײ�4�)�e+��]�Ul�M4%|��\��[m��.d��ƪ����S.Iy)^5����%]Z�Q�4e%�`pO�j�>�58�cn��[� �A<�Mh�M�w��H��
�i��LO����6�Ϟ|��8�㭴�t�==�ߍE/�2�j�H�a�(��D��+^��\�<�a�"%ӷLR#�H��U�c�-�<�t]'>�=�w�)Mh�C�w���JV�N�h6'�~+���F�:��I��jjjK��#E���f.U=H�%6�ҩh�?"�#ѢQ�TC)+5̒�Xh �^��"��M�-)V�~�]��JD}��t�]4��"��~�K�[i�`�?U���S�N!ʩU��q�ϝ|�6�?�����<��:㎶ӡӢt���=���jcvͪ�$8���I�$e_Vr�S��"���<h�*�5=�>�.�#x�9����_HƆ�{Sz{h�qsg�Yg��|Z�J���F�*��$�����*"Я��#T��,�)*�#���s.�O���;��h�bb?\��}o���z���r�0��3�?�f"N&�?>J7�tv[4pN����{^7��8^'Lr�O��<a�X�/'��N<�I�8���y|�K�>����ʃ�x�ZF�b�z�</Y>=+��G���b�h�^4�z>��	��`�����|0�0���I��2��g���?6�3���1ח�'X�'Sί����ˏ�^mo4�������k��W<���������4�m~y|q~Zޓ��q<Px�X��|&/�'��H�%>^�)�K�:�&�_��>c�/�/ͯ)�V��LD���k�����O1�y����&\yq��o1���\ylɤ^���֚#�_��0����������<��/o.�����������+ˏ/���&�L�~�'3H��dV��Y)s7�̉���p�& Na�?��<ot��f�������(��'����om��Ŋ���ʛ>8Zw9��دݙY�"�����0�DJ�� ͵q�� �'�~�oz��n�̛�,֥d����N#@�i!��V��L0QWaZ�r*�p����x��=�2�ͮ�G�k}�Rv<��؇ݣ��6Z�<�dA.�q=i�m������72�k9l�ɋ�d_l�O:x}�����0i�}V���vu��x�n���[��.X����s�[���ɯ^��J���۴G����Ҝ�!�ڍ��6N�:��6MeMw�iJ��i���k�{h݊U/�l��ճ����o;z��b�m�0�K�� ySm�]��mjVRJ�U�ËrTbʿ�э�������(�̯8�	F�:�F����;T��a����_/y��o����{�Ͷ�o�����/6�}��������m�����8��8���8g31�g���~�Kfb͇'�%�mRf٩����Xk5�\�U �J���y^�%Ɖ6���]����4�L.���.������a����`KJ6�X�J,ba��sֶT�j3Y�ģ���m���J{���iq6
�5�h.�[e�Gu�7 ��v���]-�5J�]��Z����	df�	IT61R]eѥ�B��nv0M3S&J7�Rc��@�[�#�mB�2�:��m�:�Ж2�*Ǫ�6����(�d��X��-㑁+#o3%��i���6�#ne���v'ZG��~��I�����[���k�N��i�r��ٺ&τ��4������\��|p��H��~ZѪ����M�F��n�;i/I6����Q�u�閐�Y���p���	��WٻQm}7��sWy����F�8�a�?}���9����,2�o�?6�������<�8�m:u�uIXF5K�I$iО	 �a�|�����Z��}��b]�u���!'P�O�Le���J�|qZm�'�/:��'�t�&ϓe���>#v-�]d-���SIzFax����:tD�϶�T}L�uXG+��W���+�>c:Xt�F��~�I�tgz|Hz|X͟1ǜm��y���y�^q�u��:tN���B6�����pc��|���V��[mkq�gLI6���i>�{NӍ#,&i�n]��Ѷ�U�>�0�����d��.����#�?|�ԊS���ݪ\�vH�ռB�G����b��(C?pY�&����_��8�9��̚��w�u�yZ>3�K$���(��Ozl���Zf:�.?<�o�>~|��:���GC�D�.�U�Ui�T;ʓ��醙E�4�t�2���m��� ���F�4HT�'dd/��!fa��2�~[4&�ʽ��1��~y�[GǤ�a�i�9W-�+����w_���]W��gb���$]�ƫ摍~�4�0�,��m��l�_g�#DGؔI;8]��p�e��6������μ�8�m:t�'T׆�.
�ƈ��h�뺝��$�ٍ�;i��~�m��(�|�K��Z�)8�77M��]qw[6+�፳b~��&�g�/��`A���*u�"�*T4�ڸ�Èݶ&n��1��:�ч�h�B�"��.\Ӛ�P�BΚ�/���a�|o���A�t�Ҫ��g�ֺ����9U�B%�<���@��ᗈ�&bH�2J���P��~�6��7��J��_�}�SO��Cg�k��}��Q��Rabh��uE�Æ��{���#'����3|�Z���P��z��`.�TW.�Oh�#V�Wb�%?S{��q�y��q����<p�8f0cș��EӋ뚇�S�b߫Z�S���m�EĬ��9��;�G�|�������!g� �'�zxtѱ9�>��h���8[�z��یc+�KM"#u��GU�#h�˵8��^G����Q+	^��0I�0�	Ԯ��xx$��沦-c���"����آj(�D;��e��Q��N������ղ�����>.�	f	��;D=	ƔQE�,��4f���8g3���SʖH�r%�=UZE��Ju�uX��^1��~�L��G�N]kK&���>!������tp8&���!��bIm���fa�&
�a�o���������5�S�Z�i�H}OR0�R�ԓ�i��q����O:pM�߽����z"eh��4{CG�O�j$g;Iu�h����O��i�m�Ų���M���ƞ ��3���b?B�6X���"'��ROE�	�bzt�]2��^V�߾ؗ�*@�q�W��q-�au�fᾖC�^�#Yn��ꈭ���]0r��k���a�#�G�9�<���/�#��>}�?�]�f�8'�4p��ք�%WC���%��}�,���U�(烶VQ��q�<Y��Ɵ�<A�8g3^K����ѓ@���	��!���d��/G�t�`����* QL����c��މ�S�{ژ�-;챁�����.ҍ�%Ćlȹ�C9��&��kcb\$�dB��ikUlbu�;R<�n�Sku��ЁoK˫M��-���cNyUW[Fd�?�H���<�2yh�[i��i��)��UnS�8��ʜg���~?<�>}�~�S4�.�{2��H���ܢ�m�����v��D���um5H��җU�q�{�3	�c��oȢ�� 3��o�C�#�8���M0�?S��T�W��K�|Í�q�FY���4��xg�8fp3�tn�7v��4������Y�a�ba�}���[e�FW�ቿT���G�kE�l�O"�Ǣ�]�h�,��J�f�K.��dV�,���c$Mfaߗ6t���'�x{-O��U�������,&��%yd8z{E�Y� ��m-`�هBr��{teeڕd%���2@�F]h�*;�~�`���0��0g��8����3M����h�0c4f@�01�d�2ؙ�8ьӍ0f�gQմ�V�]W]�u��ɶ^y�ox�ь�3Fi�8Ҋ,a�,e�HϘ2�1�c$��1�1�h�3��G�Fp�&��3K$��#�1�fc8e�2H `��C#C�@�3J$`��!�!�HQEE1��1�A c�`�2F20`�����s�_E~������j�7f�_sj.&��L�*��`a�γ������~{�wp.���k�s�uw#�=���}�n�p|o�+��9�Kn����:"_,}}��5�9���Uّ��#'-�v�<5-�[ۡ�L�eK��{3�{bb�6���ܺ�;=�NL���O1�WO3�.�b��x�]�j�ߜ��9�3W���[�=�$鈙�*��G^�Nc�.����C��mm����W�](��l��Ei�z��N�c��v�|�t�����E��Υ��j�b:"�/Uf�)���Ī��*��nk�֢b��j%��*�iU��v�8Wq�;��fE��d��&����]�W�����iˣ��rb�rJ��w��J�j���Z�v�y��uf���������H3z.���&�6��telD[յ��\�u��VF��X�����<΍����7;�i�_�b��`�����g������5ͻk�:{&�u�|�b�Z�0�J�nͩ[_���wk�w�^��7���6�o��������m���ww{��y��v����{ޏ6��� ��q�x�ƞ[μ��8�m8u�u��O"M��E�G��-��r\/�$6h��,��#u��J�z6�MW_4��|b���;��*�2x��Z,y!�Ȓ��)�J�j�NJ����舛J�2�H�[�FĻ,�G���#�o�[>�)È�z��W+4���_�u����_��W�mm�6�oͼ����yםy�m�������s6��|��%�/j�<�*�4ۧi��>8�'e��L��4�q;]-`��L�'s�<�ԆVό������R	�z}+v�M���C(��Oh��6��et����|3N%���=c��4 rx�G��n����4o-�z�����Hb�L����6ۭ�>u��yםyÆag�>�X�+�*Q(B�W�pL�V���C�0:�=`IY7��#�ӥt����q����o[��|�:U�p(:;V�b충�M�j���̈́�� HKE�e%�g�^Vm-�P&��c�m�,
L��ՈV�v� b	R�j�$��n1�����F!=�7G�k�3 au�n"�~88�`��u��������Y�ꯛr�z�����ϯKh���Ve�~y����_a�Ç�{r۵�Iuw��Wg�D�֦5|��P�!��wG�#8�>�G�2�5L��<ۭ�ۯ�i���p�,�C'���I$� ��i����[6�ԿI3*l��~^�x�mUu_�N�Io�}����~����U����x�z���M˝��F�>:9�L���[c�X��0�����^xIw�zhL�9�t�y�I�y��>f��1N�1X#��T�}Mv�F_<Ӎ��Ϟ|��xg�8fsI�d̤����h�j��C�5(����Z�D�8+v�A�M��=�^<�ka��~q��郫�1�k�����y��d�/��+S�$�wr�,��;�xwTz'`nZ��Y��u�Od�W����D|����-W�~����Ƀ�{&i�Ʃ��N�l�,�Y�Fi����38c���U*���dLZ�ѝKfb2�w����\��H��{���ڡ�b�9�*7};	�Y�����UPNW�P�ĩL.�f�m��L�kV�y{���Tw6�=��KU��CSG梜�D�$*J�E�����(��#7��ߥ&=$�-�i�^C���}0Ò��it�4a>��jP��a����̮$I!a��P�(���
�J�EM��>߉;E��x��x�K?3O��ǎ8f1���FF�"M~y�4��Lc�fSfc��$���bq�n����Ol�P��!�������j���3nM���J)����l0�h�~� �M �F(�zF�8�%�`��LH�i	�^'kQ6�(ڲK$R��3�����77�l��n͛��{Vv�k��b(����;FQ�U;A�ʝ��%����.��0�9_>glW����L�x�r�WIF���;_��'K;e�x�<��'�e+�BHNMh����
��aJ�uf��X�o����[e��õ�y0�yl��M���:����<㎶Ӯ��X��/��I!O�>|Ǥ��],���Id��y�9M��GϾ��ʺ����~YoKV��0�&>�;��#��|��?q��^.�©��}�VV,�of��
9F���������o,��%aX_���)�/��0���Ϛy����<�:�N���r�8>K'O� �~Z��2�{��~�|6�(�v�����8ӞHJ�t�k�mzEeǚ6z}��y5�`�x[8{�5Dߦ��Y��jc��M��M�j�&b�a�m���x�y�~��p���T��`ٷ�����O����\#�m�}����wqRv����ݨ���< �,��њx�#<x����q�eG>��U�ӂY�A���r�!�^_�{fYl�-Uc�A��V����0�j��MѪ>�O����"�F|<VJ%|w��;�����I�z��ӕ�;2�aaGiE��'��ǌ�<������-��u���t�㌲�n<ۏ3q��d��h��3�I�8f�h�4b�i��0c��0f���3L8��"A�C �@��!�p��d�e���Lҍ�<3�<Y���Yg�X�$&!�0f����P�0c4g8�gA�)�0f3b��Q4G�1��c(C$��1�1���gXq��ӭ#�GV��:��Y@�b�@��1�1�c,��3ǆ:�J����ٷ�����Y�������ܭ�[�\��6��cݹoz�t�mXD�+Z�X�fQܣy���7rF�n
W���u��Zr�
cU��Ň��F�!�� �b��n̲TJ?I�,p��GH܊�_F,Bħm!��9�hq�a�Y�<LE�j��� ǲ7q��6�Y���������7滕��� B[[R���ʰʹ�kXU�Q?7�[�^fv[�V�݋��'"��y�VD]QH�"#n��_�7w�o簶���������46�����hأ��_uoEW얞�_r�K,+����?f��mz�O���!�DO	OO�p��%��{6& ��m�=e�A`�c�0fn˶�'�"����8<�QǵU(c�r���r��+t���z6�7�ɍB��#���5YkV��)�G�c�^>��^=�Zn6 ��ph�,r0����j#��B�-̨��N��^9���q�c����W�{��������������{���}۾�����O�o���������m�v�i�8�K<i�O$g�8�X��p�
fWDN��Kih����v�in�,s�c��&�[f0cQm[aۡ�å�v,̺�M�:hZ��@^h��KB1#���M14��ȋ5�k+/�����V��u&����Kpgl�R�ɥ��˭v�l�bL�]���ۭ�1Zi�M��4C��[��B�>�'����Ki�Q��]�uG\Fb뵎!l���t�w� !,����u�A��5IN�sZK�c�&�i]��m�������Q��+�b0���P��g���Y��l��;e�ݑg!*��Le��Vre��[o�V�K6D2�1O�I&�;\�3懶;MS�֙�(6x�߹��Q*��(�~���ڬG�ܜkf���ŻO�ͺ�\��^1}�݌�K6�5�9V�Do�ߥ�#	�am��k�~����U���~�OUq������וuy��]㎿0�,�q��3Fi��#<x����233�T�*�	�R�T�����7N>|�4�o�֪e�0���7֘�2��D8j�~��������E�?J��ye��V�R�>~��'�cn2�y��<>6Vtӈ�^��h���䬿4��;�6e�Q_8��D[�6��Ϛy�$g�8�3�@ʩuk��0q��U�Wi.�9(���C�r1�bsф���>������/mSR,�l�1M#Do�������Y&����OL��E�y��_���W٩I��������Y�i�w�\x��-�A�3��4�G��y��;L��8e���ӱ4ɵ��ݶ�:��:�����Ϟy�^y�<`��	�}���W�$�@�Kq�q�����4�4普\�l���}����˭72�ve���̚ՖCZ�i�c:�S,때^%Ӵ���ʝy����񦝧)��h��I"4~�-ZE�!����/F��Y���G*O�˟��̺�rD�t�;�'�S�6�$�_fֹ����:����˒Ȳ�Q��iǍ8�Fi�Č���x��1�W��+��!Z��'&D\�x:����1�R:l����3=�a�en!9�hȑ1�	�3M��lĳ@���XW;��_'� �FO� !]��Ð�K *���`	X݁Y]b*�\,rn;��	�ޟTo�e�		F}����|p,�0U7�ޓd|F��$������6q��EvT��?J�:��H~O�(�?l�A�]�_%��	g3�0������1���[�ɘ�Dօ�R�rTfC&���j����i�_�����m��֜y����|x�#<x��<`��:S���;r�:Z�]m�$|Y��4&U�;,�nKnj z�a��6˚R��h��I$#O��"[��r�WkO�O��-�j��z}LS�)�G\��y���*���}�˂jI	(��e��J�oڳ�ȼ��8l���=�Z�l϶i˕D�u	��5�s-s&%V�n��t��)yi�i�mm!�in�XlɆ�,=n}���?2��???>q�oϞy�^y�\y�\u�1ϳ���UT�J4tK��+U{#�]/����Ma��l��+4�O��=���X#����Y72��2�f_���v5j7r描i���}���b����f.��r��^�6����{��ez(-3�Q�&u��^eưRjb���nk�(e�� �O�����'8?��wph����F�h�ӗ�}HקCT|%kjv���]�k�.���\m�?>y��u��y��:xt�gE���4R�U)T�hS�vz��	�_��$e�0�q�)��m�Դ�ڱk����rB+#+�W*�噙��M��ѻ�uW-��5]�j���ф^�U�4|r�3H����}�iOѰ�����_%�(�,����j��m��|���?0f������"�i�4f��Og�Ǎ�&.��*��5w5����	�u�b-��&�D��5�&���o�)AV�y6V?�\����^�E�SO������kP��Z�z�O5�b��֫�P=��H�L�fZ��I�����,�sf7;c��3��ݥM��JJq�%0��e���W)�3��,���&����>g��T|���� �����/Z9�S���/cG�Q��W�;G�
��Jϑ��=p�x��8 ��ߒ����W̚�� X�a���c��]-)��H� ������~,0�~ �<]��13"
<Qg?xјi���<x��<h��'��K�����J�	�Yt�Ca�/*�4f�4E�Jy�����W��>�Hs�1{��(�p��gw�M�sa���5PQ�P��Y��x�Z��C��Z+�Q��S��.�/�&&+�,�(�^��Z����l��/�=�������}M�D~e�j��D����z��y��q�F`�3iA�8g3Fh�8�h��3��Q�&1�h�ƌ��3L8fA �!�Y @��22K$c,cĸf�3�p���8֖(�y��a�a���V��[�]Q#(g1�3��p�3�4d3�H��0�ad�!1�c8c���$�0`�!��&2�1�јa��C��YZ2t������[���ьc(C1�c#⎸��,��^�y.��7��5�}��|&���k�%k棽�Z������JlwS��i���<�C��p��w_�]o};�3{��\������&=3ӗ�9JF!����tnG�qT̥9dj�9�s�����}���{ޟ6�wo����{������ww��{��}��qGqƞ4�<2�<3�3�2NQ�U��(�=W�7�Hl0�9FUBG�a�Os�,��8?Y���5��-]����wQI�ؓr!v��-�/�~,�]7���>ǻK���I$E0�O�S� ���-��ۦi�a�.5�}����H�t�>eu)��N�i��y��Ǎ��4��x��xќ1���D��,�{U����G�f�[,Ѽ.��]T��ؗ�%��ta��L�8Ifí[0�Ξ= r�̤%\�B��"� e}��FPh�u2X��ItC	D2�V�!�!��>T�����l4l�Z���Ұ�y�:ە�h�<�|m�w���q�x�ƌ�Og�Ǎ��|��Ͳ��_.P��sN�d1S]�!w7��4�Tǅ�"��RZ�2a2���K)z�+R˺֚0S6�X��-jW�� $)o	���ݕ[4&�*�Vr\��93�+\˫tV�f1Vz~>�;��M5���P���ŏBN�Zezj��c�z3(��Q�1X��hZ�}f#�5�[an�O�?m�������J��3ᆇ���u�oįl�h�]�GX{��4�����Q&�o��6��v/��X�]�Qg���z�0�ߒ/󍸌��O�|�Fa���Ǐ�ƌጒ�ig�KJn��Mf֪�'�Ϩ�zh�Ki�l��q��=O?wm��v�l��Sq���p�O
��o���,�C@�~������Ҙ|y�X�Q�4��{?�cd��SR6�=#e�[&j���2�� ]w���r��͈Y�Y��(�V�����N���]y����[|�δ��:xzp��ӥ��"&�=UUʭ��F��5���8����d#����#_��-���M3L2ɚ��\;���Ee��AA&�"�q~�9�J���!^��f�͎�h�_k���y�}i��&_"�t�O�b&̰b�<�ܗmSm�mn�]��uĔa��ƌ�Og�xg4gd�y���+��N�l�.}��e��mV[�R���s����_]��ՄJ�]}T������?}�7<�GI~���ߦy�U-]��;U�ᇅ�Ϸ+(D����~˾�2ܹ<.O�P�9Z��+���dd�iP���3�֛q�����Ű�w�WUiK~O�E֕������TM���<5T�Q��&��v�VZ4���le�)��!�[�}\D�5Z}IO8er�O�]y��i�|����<�<�θ��1�r}"̑mڴ���?��R���.�d��c�#ҟ(0-�WI67$�0OX�s�	A�����M�{:k7kfo����M��� $&��y��`B��l���w4,S:�`�a�l�b\L�ø��Y�P(�^arq��8,�����\�gŎ=�q���W��Ӫ[���u�+�~�|i�}w%���q�v�d���ޗS32K,HF���A�e�7�x_�L�s-���]NS�8�B;Y�~�%���������YD�22ȣ/L�ܑɞT,t�f	Â{.��>i�Ϟ|�o�y֞u�\zp��ӥ��<iA���)~�UB%m��{R+.6h�:�LbSO-o�%�j�M�̻�g-�Z��8��Mit����w�i�)*g[�s.ƥ���>WrA/F[�Fke��2��B�̹��ۿT��䮶�i�L�n�cb�<��m����?q����ܑ�2�v�e�<i���f�<2���<h��E��˰��u�ٻo� !{��`�.�˩������/���K$�O��v&i�L:�u�[�r���z�v� �e��9ة���×0r��4�G��=�T] �N}���Wܙy���"��3���L8��obc����8���q��q��:$u��$f��8�Ƙ~4f��OǆY�Ǎ�$���/�P�!"��*�	��'M�`J�W���v�Qbib{��l�Ⱦ��㓐��h��#Z��9��U�OS��Yi�Z�0a�OҤe�si�2��vS��d�C���V��o�櫬9re�����t���ʳ/��Kory]a�N��6׵�{OjA�8y^�vh���z34f����h��:��h��3�0fH�!�e2�`��И� �2
 C>ac dd�H�X�`�h�p��8�3	,����ǚe�a����#�e�]iwQa��8��qf���`�3ac4��Q,dd�c,c�,$d�@���1�1���o�i:�:�udt��2�Ƞ`�!���1��2D0a#�2��d%J��})̧��9�jBA�$�"	S�#[fb��Ƨ�w@������oz�0(�r�ar�ml��v�
!J�С�VY�s���a7�u�bd��}^��yj�!�n,��q��1�Z'G ;��֍�ݼ����q��#�0�	��cْ�\.H�H1<�+�5��2nľ|h{7���,�_8�F�u{=-��g��p֣q�k�G���)�>	����|w�(�a���*�>�����\
�$=�j*��D��4cSff��
�ٸZ�V��ܩ���7dDL\e��on��6�"�Uy�}�XV(�ܡ�}�}��~������O��kTwϲ���}=�� �9�&����K3�LW��j�B�z�2��A���n�Fh� 76��>*��˺�w��9�U����w<����K��Mv�R�8 ��E�"�K[R�_wlAt�+�X�x����(�o+�B&C2U�[Sl���Q����jF��_��+���߽^ow_o�������{����{���^oww=��{������a&x�<Y����<3�3�2O�d�Dϼ���α�e�GP����f.�c)m��bY����k.���Im���H�����Mc�����Y0�,L�Zd�x�e)J�7S.����I�a�S�(��{̞3m �a����[(�����+�,�eԗ��&
�v�Ń�����E-���˲RRF�Af�VX݇%*$��QHi����Ũ�-�HKx���Ķf�ؚU��m�S�E��L�j̺-0��UA&�M��D��m�"�X�t�m��[�2iR�+}=̭a*�Yx9���~��K�pOh��X�y����.����%�is;e�a�Y4ѭm.�j��kU�+�SL}�vL>��c�ۑ�������ڦ�,!��Â�w�,�W0�p��B��͖wp,_:�U�SB",��e������ۻ�r��%,�^/�E���/�5ڈ�&+F9R8���8��4�ǟ?2�<xg��xњ1�UB������kg�&�Ce�^�C���an��O�g���1��%$V1��>JW�"eLp���HӏS�s�Æ����f������BMm�����A4l��^�9�&L�:iSx|yAæ��#��~�wM��b�z��>4���/�i�~q�Xq��\|��Z|��3�8�4c$���$��I̲��b��wk�����K�Ky���]�OWՇ�WԪ�l�b�!�/�w�%��n�%�ȥ�]^s��8f�y�e�}_<����9Re�moR�e�蕇\�I#�>�b�d���LR<��f�q�ӵ(j]6s��n��{�#���a�8aP3$$њaƞ4�4��0g�q�Fh�D�\*6~�BI%�"�mk����MS�Y��Oa�L�3$��8�.[h�!�j��Τ�V��릴��[��/a���<�!��L3��0�M�m��L�������.��^�I�ghBUC�V���Y��� ��Nȳ���f���Z͛�??J�>[�4���x�Ŝx��3�8�N:$<�Tn>��K̻R�Yv�C@%XI1&[�kcH71&�Y�.��H���m�,4�16�B�k�[��Ɗ$/[35��O�� HF{<�h݌CVU�4��]��7�+���K y�8�nҦ��F�	�������*V�Z��6�[t�&����>F���B8�u�'�m㴺w��3X�-�ND��R�[f��}X��W=RJۊ�7�f�J�F0�9N�N�9G���yEن���0�Y$��,8|�m�Ի�vt�����F*�(d�P��=bӊ(��8f�4��<3���xњ1��rFV���0�Α�{��	��ճ}��׏��X:ܼ��`�����Ad��{���RH����	��TIyG�����YIL8a�?}"��j�O��-<�x��p� %���J�B}�Jqu.�n���+Pbp��UUS"�S���0���U��3�͐��*���m�i�����\�͞i�έ�+5�b���`�Ze��a��|��ƞ8�x���xь��I�UT�6ٲ_Q��YKVyCm���Z4�[�~�M���5X#l0P��,ｊ<�UMm���/�Ș��.�f����$������a��d,���j����VP�JH]FQ��<��}�<�X��������&Q�N.����sc�����ʒN�2�1U����\u�Ϟq���<1�4�3���Q3�~��y��I!�|�ۓ9�s�M�����W+¡�>x��n]�L�Tô�����*.��Lݘ��4f�~��_�}U߱rS�f׶XmL5[Ԛ�O��O$y�2�F��4�����̰���x�ϩe�%F�VU�b��6p���4�6��>T��#|m�5���4��M��뗆�j�?af�3ƌ��4��3��O1�XLܘ��\��8�"Z��7R���E#I����N�q⚞�[RƢ�!�4�����Ķ��~)˻)-lb��Ɉq��w*�!g��Vӎ��p���� ���gN�Gbp��Q6�jU)y��=�zy���0�
�&��D�v�)���ȕ���䙵Ĭ��-�u�ޥ�=L�D�u����'�wlg�0��[�&�o��P�UʔryE���F�#�~\������#x��,5��;��M-����o�e�^$��*��F�O�&�����:��/���SӯSO��s��r>a��p�x��4��3��O1���C|.�t��'s�DOM��E�yz�ˑ�#��$�-�)��#ꬿ6�c�]�r�3IQ+0���اF�4F�NV��k�*.;�;�`�������E.\R)�/.34�8h�$�Y�����ʬb��9Fm\Q�H�Fi��l�m��͸�o�<�8b��3��4f�fќ3�4g`�, e���e2�`��0g�1�C$B�`�$c(��2�33�3�p���3	0f@�$��%:u���u��N����ζ���p�3�����0�-4f@��&2�1�3�iD��!����1���c4c4eaӮ��#��u�,2��t���ip�@��1�c8g�2�@�S���o���K����#J�٣%̔<��'m�Tl�O�K����7a�r�뾨u��qk�EL�ޅ���f�o_�ڥ�V�o�(�
śGU\��i��o���owws��{���~{����{��������������_�����af<i�Ox��<`�g�<iប���̹L����%�6��un��n��%M.�4e�/��ӭ�o��X`x�=�\�]�[�qlp��ƛ���Ud4�r�(�Bj,Yū���+�Ǯ�UO�]�NlYG�o����_�%���˦���m�K[�-m�E�e�q��4�lI+mc��<۬�y���ϟ�y�y�^u��y�ή�+<�I$����]�z�b��)O�خSmkқ�L}��ut��ZYu:�.�/7~t�>D}Kh�8�n��O�ii�z�Z����ٌ����-8�l�-Q�m»�xJ%C��\5[��K|��)4�*U�8j��ᶈ�i�e�n�=\�|�I[����[M#m��e��uן:��y�^m׌f<i�&"OT�ҪA
j�4���M��WM�>s묮�F�����W��G�X�d�V�baK���s��L$�#��  Hw�.���Z�7*���1�=]��X�,J�2���3�ܹ+a�
�jh-�΃+e�unק������A�]ݑ]�G|~;�L(0g�6��
��$��Un#(eyDDf�V�ka��l�9�o��U�h�%���ɼ��n�yUe�(�4j�P��(5����~4�}����QT����h�&���kg������z3F\|��DD�G����/�������ϖ���q��>yǞqכu�Ӧ�ON�%�6��b�����Vr���4)�*�bp�!y�ahj̰Õ�X\�rbX�:�p�V��'jH����Uƣ��(��p��6˳u��]ّ�2��D�%�뵷^y+�g/R�e��}ke}���M�w�ƛ˔���P��uh։<�)�f[i��3�x��<p�3���xb��)�r�۶;�n��b������e�U�I�魛x�i�����{�/�|i��t�3H���2i竺g���dJ��+�3��2��̒`�>ϫ�L����QGTa�[UER_i�a��Y'4�f�����$�Ѻn��}ֻy���2��Iq*B:]4r���u���[l���3Ox��<`�f<i�k\�w���Q��5j��o9GKV��n
��b.��wB_� 	��0#�ۏ�#K|z������.�>�N�K%�p���Tt�h<��p<0�te{]����i��T��١s�y�=uP�$D;j"��Q_N�LDo���]�vBWh��f�ɇ�G��O>��q�uf�L9O�W)�Z8��1�~4�����8�ǌ<|��U�jM� �T��[{��$;zU�|��0�܋3r�tx�U�s��qa#,Y��
�vn%�Jފ�y���5�%���_� !fSu�Z�D��@Bhb^x���6����q C@�\�Q����ه0�n����]���(3�H�(��Ņ���/�\0�}�/��Y��'�ᒍ��̿0�������縉e�l��>m�F��i1�����!o��ۧ)�~���9���Wv�,��gO)�%�3���Ē2�4�Fi��<1�u�θ��y���{I$0��j$�N+�>Ctˈ�|���JaQ�
#��.�ٲ��ei痫�eT'M��ݻ�T���e�b���^o�GI�K�d:lõVoo���;V�m8�8a[Z���ǧ�u�Wv�Ʃ����L��o�|��t��xf�ƞ<aᑰ���о�� ����&#�B����lHψ�9��R]���-��;��kX�J��w(�B$�����j�*ꊭ?/�b�X[�6]�8�0�|r���]7Lq��h��7��ї��q�BF�WĒi��<h��ƞ<3�<1�xgx�"J�~�/Zח��U�J�I��v�M%j�O������HϏ��ti�,���<琳m���F*�"���[���Jr�t�S�R�*m�I��ڒ$u֝yG�q�`Ӛy�>d�ַM8c�������*٧�S�%�Ə.:&%�DY���}���F�^��vSJY^Ȭ���F͛7�|7��L�Y���[K~g���\��Ç�6�ٝV`q�έu��G�s(�J�˦�
U�*��q��5�$$Y-d@�!��R�F��$H���	���" �B!d"$h������!"B�H��,��,��"B�H�!h�"DD��� �$H����BB�D$H,��d$h�"Ȑ����$Y$���[D�ȑdIk"H�K"L�E�E��D�ȒIѤ�Y6�E�"K&�Iid�Id�I�#Y4IMY2K&$�5�h�d,�MdwM�D�,�AdHPI&�h�Bi&�h�ɦ��"k&��D��M�$Y�8�I$�L�)���de�L�h��#DId�6�h�ȉ�ɢkM�D��D���ۧ.	� �$Y-4M��"K&�kM#YI��&�MZmd�"2�H-6��I5��r���Y$I�I$�h�H�dH�$�,���$�Y"I&Y$�m"I%��%�$��$k$�-$��d�YH���-$�d�,�$�I$��&�$�$�,�4��i%�$�i$�$�,�d�$�R�$�e�KD�YI,�$Y$��i$�$�,�$�Y$�i&I%�DK$�I�Y"IdD�dq6��,�DY,��$�Y$�K&I$�I$�ȚdK"$�$I�$E�I$�4IMdZD�-$i-$�KDI�I�$��$�h�KD�&�%��I�Hֈ�Z"Ih��p��mi"Mh�YY5�I��E��ЛY6E�z�ף��N0��gh��"�&DdFE��6�2-�f�6���b8C��F�m��LDȂ �#�<B&�fD�,�1�&ȶg8a؈�&h���� Db8C��al��-��D�M��x�,E�E���l��ah�g8f�h�"DdCE�nx9�;�,�&Ȇ��,h�h��f��� E�E�D4M�6E�D4CYq�q�0��-���AlDlD�LY��E�F�Dh�-�Ah�Gq�-�M�l�ȱ�D�#�8b-�#D�CD�[mD���� �"b �2!�b#"l�l�14FE�DdM�lE�A�"-�!�m�a4M�[mm�h��h�E�Dmd[4Y�kl��&"�؋XȘE���4��m�F"����"�n�p�d"5��4s2FH�ЈZ4�����D��$,���5��Z4B��2�kF֊$$-	������D�B�!"���#h��#kBBD�#kBBAdiBD��H�!dH�#Z,���d"BBё�!�$��DAd""E���$$Y	!"!dH�Y	! �5�&��B" �""�! �-��]����E��!d$-�A"F�$$H�BD��u�$D�BD�А�dZ$$kBD��!���d$HZ	Б!h$HY	�������!!dH�!�H�h�"BȐD,�$,�D�BF�#HB5���D�"F�""F�ヂE�D� ��"��d$DZ,���$H�hM�"!d"5��$HZ""$[D�"B�HY	D�E�!d$HЅ���H��F��$,����F�����m��Z8xk<�z7nY�x�3p�ہ���n��Ƶ�mJfƖ�:�\g���������;��^?���s��~�v�c����:�>g���x���8���8��q�7M���7�p�|�����Ӄ�=��~w;zS�o�����OKs�:o�����w��������Χ�8oW�æ����ٳf�6zG���o�����<�������o���6o��p�K5�7�oϛ��u���g��c�D�o��p���o�3���D����_��5�W�y�ə�w?f3f��qg������#�8=gvۖ�v�����6��oI�vs�������Y�q��;���a���|;v�w㳺=��Y��^=?���n��uә-��v�]�_'�vpFٶ��sr1�c�ͳf�r�m�ێ8�=Pf-�͹���X��|���h��#8��rt�_C���n����O��^��ކ��Z�`���q6H�(�����l�C6�`�㗭������4�,�ۿ~go3y�^d[㻻�z��ށ���wa��Ã�����oűo��>�7m��o�N�6l����w���v�[����߿Kn���z���nǠy����]\x�[�{���>'��?������&[s̞��7�z�=X���<~{�w?&��ьٳz���׆߷�O�y8����x�]���>����6z��׍�f����lپ��|�̶��;��L�\.y��ruǓ��7'���|��9w�ݐ��?o>�7]�7�VZ�ɹK����o&s�Kf�b4r>���nvn��v���w��ٹk����8m��7�{&�glw��o������s~��~n��3�J���n�lٸ��oW��%_��ף���v�c6l�㟥�7ޛh�3ٽf�_�t�y�_���������{3�������#��k���V|w�����o��o�#n>9�O��m�[�������6o7zzck�m�ϻ��f͛���c�xw���7�<{o��g���=OS=�=�ĝ�����͖�{�����"�]���ѹ8}(���L��>�W�<m����_������ʰ�YU�����f�7�^��m��L�8�>��f�o�8nC���<�o[w���=�ߞY������$~ß4V�K+~$~���8Uc����L���l�[��G���{���7vz������G�t���~���>nݮ�����u���|r��9����h���c���/���"�(H�9��