BZh91AY&SYث���_�py����߰����  aP~ @   @      v      m�(�          �          ���JD� DP��}�`� �) �(���y�{�������oy���m����^nރ�מw������>exu��E   :r�N���{���}�Z7�}�`w����4p���]k�h^ƺ�Ԁtw��   �*]b�����<!�U��� ��l(�f���Dy樵��S�WA�a�X�{�oG��wc��(  ����лV�;�.$z��J�C�;���=���p���{g�5Mi{h;n� �[`&@��]�B+��t�UV�H=�(=�U�Rֽ�j�5�û{0;����C�=s8 ͨ�X�4-s.�;oG"��z�;yO'���#m��ק�oG� ��2�FʡKŀ$�m�v�[׸ywX�R��ל=�xh.�����O�^�O:��N� �B�}�}�ݧ�=T�{;����;��sNr8��z��u={�8 �(�
��
q�:���wg��˶�]9
;ݳN��5��=�Y����=�ӚHc� ��y(vc�{ؗ�g���k{N{{�{7�%��^×^��                   @ 
  U<�?T�R�2ba0L�b4�`�����*�F&a10� �24�4�)H�UM1� #0i�  J��I4J�!�0�a�L &MbST�	��e5<
zjzL���SBf�����L�)2M��C&A�C@��g��mA�jemL�X�b�Ve2�F)�i���{��|N�k|Ͷ���w<:�[���
�Z��l�SM݈��a��f��ٰ�ٳ�������8�����ο�?��?k~���|�nǠ������R��؍�l̈́Έy�O�˅ʫ�~�ٍ��x�3���*���l�m����|y���6�'��}w���{������1�����i���e���1$�F���	$ԓ�La$��Y̓���I>k��'�c��jI�D�K<�d�%��g3���M8�ǲH�<��ROR��<I3$�%c�Lz�I&�?_��I>�q>fx�)'ɗ�3�I%�m&�R|ܛx�q��z�Ʉ�-=�m��֖�I�1���z�&$�m'<x��RO�ͤ��ߤ�Iy�"I�<�I7'I3�I'�_�I4��2�|��'���_�ޤ�I�1��Ԟ'�I&��I���I&Z�x�ٴ�O3�/��Ov�O<�L�޹8�)8ΒK���y$�ƴ�L&X��L'�M����s�ϙ���^��M�ƞ���a&�|�O�MN&��*m���1&�jc�[�a/����a4��R|�|��OYe���nL����O��Rq��cL��׳O�O^��ְ��>c׏S���Y�Y��0��l��q�S�>m��~4߭}���L��3'�n7�{��=���$�x����ɹ�Ƨ�����I��$��&�m,co�2���I��'���e�d�؜�10�4��#��/1�߾N>|���}�iϞ_g?��׬��M|���>s��8���6���i��gɖ_�M��=a�|�5�c	����G]}�l��숍���u�X�N-��O����.c$����q��׉����V>|��֬m��}�&�����)����I��1��>&2�O12�c�I/q=I����O}ƞ&V�'�>�$�g��a��cL�Oؒs��g���Kx�����3ԗ12���q1�q$�=�&�'1�����e�{�O��8�e��z���$�i��d�M�Ǆ�cI'�����^��I8Վ2�=_�ğ$�|�e'�Ğ$�q�q�K��N&I'��1�y$��c�N$�I8��cl��/1$�?X��$��2�){�$�m��>���$�m7�'�%�O�Ԗq�I<_�M}��I��z�_����I>��O��x�N&��$��$�[��a�^�I6����$�|�Mg"Is[|�Yǩ$�z�L��I��SI-�ԏS��|�N~�$��^"M����g��'����<q�i�Xd�I2�i%���N=O�^��4�|�N$�~��RI=q���sɝ�i�y&��'��I���$�<�q��0��)���&�qL~�ORO&�a>=e3��a$����I=���o�I3�I��$�q�(�}<L��~���0�H�>M}3&\a-��׉�<�M<q��ORNO�I'���$�=e<��1>O[�o�6��O�7��~���$�K���m&�1�̣ĳ�s$�K��g�<O��Ա��2���I/��I��$��LI&��9�	=�N'�6�O_$�q'�&d�I�bq�	7�$��ɧ?I�I�be��3�I$��)���I���I�>I�c�$�r�)<�I4�0�gX�z�lē~�M�I���I��$�}2�|�N&Il�I<�a���$�Si=_��ݤ�a>I=�a���L��n1&Rc��I7�L2I<�<L'�?m�I縓I&�}�?I��em����ĘI<���O_I#�ޯ�I�K��y$�ycl��Mͧ��I$����Rm=_��$�0�G��$�KlO�Ēz�i��I&��8�cI$����L0�I$��m&RnL���I9�s��$�|�$��&�y�$�i��$��	$ǘ�I1��F���|��.u�Zˎ��a�;}s��a,�f�CD@؃ԠG����$xwC�y�>o��k-�Xˍ=O1$�V0I%��I5�I��O�M����N��I/�ē���SI4��.$���I��c���o�m'���8�z���OR{$���yc^��ĒLix�i�2�՜I5�&W�\OR�9Ēi~���
�K�I��	듌�ɦ�1&���I=I7&�4�c�O�Kl'	�I��Ğ��\ğ=I/15�O�?{o�L�$e�H��:���w8��J���;�N$���ǅ�?/�	<Z��&ڱ��X�i�J��q���lx�=L��$�|�a������,������ϽĚ�1�s/��SMc$�ěa+��y�%�IǶ0��-bOV��W�/�%�F�^����&\�K�bN�պ�:���"u��x�5>I���M16׉<��I��i����	1�e�/1��/�4�Mk)��N'��s��q��5�z���D���Ikx�^bN7�|�n~�I�1�׫��K�y��^�I>�$�kO�h�^�Ē�8�O�kOo������/����'�3&�ZĒk�L/1$��=I>�4�zĒ\m���I.c>rm��6��޼e���$�NL$���_�ĒMOx�I�bI�M�O_�M����<i���䕍��y�$�Mn�e'�M'������I$�kO^��I4Ռ"x��I&���7'$�q&SSi�~u�뮲�|��|���d�z�+q�i��I,ci"-bI�XĒJ�I����I��	$��<IgI.bO_bI2�~�$��cI'��I6�o,e���o���ǫ�$��$���I&��I/q$�V0�Kx�Ę�I4����$���$Ӌ��I2�Ēx���8�&Տ\x�q{�8���ǉ&lm��O>K�|�)��q��M�e�L�I>[���e$ϸ�I�,a�_&�I︚x�Ny��RL���q$���0�|�x�����6�{��2������ra�^|�z��-�e'1�_��8�2��|�ӎc|�N58�+-��i>f}�z��u��_��x���M&�1������i=a�o	���4�����\ǛV<|�6��e��&<I$�sI�O��ϩ&�&M���I'��3�$��Ğ<I��I$�1�&Ԙ�q>m�m�cSno����0���v%��������t`�:�v�q��\�f��_Q�:��}ִ�nq��Mq��l��$ޱ6ÎM2���Is�<_��/q$��e�$�,�M90�z���L���4�i��̮7�ZF�M��'�a2���'1�m��穧�'���fQ�g�x�I�cL��y���I������dl��H���Ëen�i�;]u.bOc��$�y�0���O.g?>M7�|�ľĞ��N<_��k����~�N/1��>���4���'��z�Ư؜I{��6�oz��1�I˘��W�e2��M��m���gĵ�'��%�I.bq�eg����S<����1:�����:ĕl����=p�.���><�I�g�k���'<-���r����Y��_G���9A��8I�D�6���z�r���덜�PM�%���ff.LX��mR�`�^�Ʊ�)Y�c�K'5w�{�����(�b�FEt�������W+St"���맱�֤v����f�b�db�X�mou����-E۪1� ��'}�y�C�j}��I�����-p��t�G	^ڦ-v��c��8/�;YO���a�#{\P����Ǎ�����g�����C����-��-��/{_kx*��������QYI�J4���֮K��q�B��������(`MV�|>Oݰb�f�}��z��Ԅ����K4���ۍh�w�?k�yy��4"|�e���ų4a���I5'�&�v{[��°�;���6����� ��ݷ1f^Ӕ��xz~Q��`^��Q�F�j�g]����}(�c}����^���#�������Kp�n�6�]�]�3Řu��/(��Ζ���ח��FP�bG�8�0��lê��L��3JAv��^��GJ-u�a�(��+���m5r���Te2���\e��M9u܁C:Ua�MzaE}B�T�d��^�vS�r���u��m���}m�,�N�p���3��zuk�
]xQ�	c"��~W;�'��p�f9�ܸ~A~���+y�ʆ���o�o�ow�o+�8qA3�y��;[���Qꋰ�:��l+|�#�T͊I;��=4�y���Sm�uw�νp��mu���L�W�
D��J7 �C��s��q᭥><��{E0�]U�܂ϣq�6N�~m���:)�qMG����0��~���d@Ю�l��8q��X&`X�4�M/�7�n�K�ǻ��in6l~�eV2��CSnfO�7��6��!S"]�w��:�Q֜�ӅL̶�[��Bu.%#6��a�k:N�N�'��V�Qq�Xh��r}��l�%{+�W��HلǏmܩ2���+)��ש�yQ3�\�Q
�T*��ۃS`l�e�7��X�v�e���DA�۩��,m�ɂ���aM�	s#��
�δ�3��EϞ���l��rŊ����Σ~�􎢆���Ǉ��Nզ���l���]X�c�] ��W���q1p�2�yC�&�RI)9�#yO���k[L��f,���u�TsN~�a�����o�x#�z�iɩ��߲��llW��X��s��Š��N���3�yw<ᑙ!�Oon�+ne�ѓw`�b�*���s��������rW��dd�ҵ����ٗ�"�YO���h׆�s�/\��ҽK�q��p�a�k��V��(�a�.�����T�����e�zEу�v�M[W�p�q��d�\Ȃs⩅��c�����$�;�y��4_���=&�s�7WFXa��s#�H�ˮ�߭4�]p�d�Pe�{	�Gu&r�͹�kw
��٢��q�ä�2㧇6��1�n]+R�u������,�'-��j��,�gQD��X�B�ѥd2�����9��O��u����pT����K�ǆ��F��hZ���'��}9:��	�+K��]��>솠�q���7qA���r��'&�"�9뙅i��޶�8��f�������x�~LzDdNæ�m�y�>gc���Y=��˒3_#�܍��>��o�ܤ������j�{D�:�������*�H�j����YSsK��a[�,F��V��d-v�GPm�/�?�+�g*4�U�&x��f������bh'6Ge%�[���]yAl�����/�3M�~�IIou�I���Lά{������|�SF�z�}/��T���!�?m�#�ͯ�擼8I~����ل��6u��������\U�s�kηn���o�t���sצ˶3Ҥ!��u�9m�zYT���z�fa7�9���DT_����	$�������7f{L��䦒���n�]E��IF!�a�j��
��B�#�DŬ�z��)x-u�aY<N�yJk�1�,ʃ���d ����f໌#����Ǚ��u������jC�1����q��$a�f3(@�k,�t�3�%�����BUm�	vX#LT��Y�ȯ�����߫�;���r��Qߵ�<�}�E7�}���	t'���sJ��y��/!(���t�w,��1H�f�i��`V��{��+���^�)��;V2�!��mۦ"�2VT^�=��ޮ��4�^�Yva³��I[��'SU��>nw2:{,0ܥ[���o�sU�ٴg�#z�$��:���u�n�qe��n��s���g��U"��y�<JQ�,9��N�8|S	�7�T�*)/_�<y����ǦHK6M��Shŧ���_�o\͙��Ps�sk{L��m�ͧM�3x���l��ɮ��Q�*���ñn]�g�dc���\��R�N���e��6i䭦*b����w��ˤ�IE�p�����+��}��Ml�T~��ێ[��}�Tܔ�A
͢Ib�^�J��B��M�8��r<=Փ��+�6�ԟ��=B�����%�{]���L�Y��(g�w���!���p����"~��y��=E�Op~�{JGK�y��GhAc`�l!��m?�4iD�#��p�7�N��O�owb>(~^~2F|Zq':z��7��C�g�x��nҰ��Z���~�_RJ	|o�M�F���N!�OR���ci����zl'_�}��p�l�FI�vj�D��gp����q����L���gֺIe=.ȤG�!VC-�Q駌��4Č�]��KT��l�$u�ۣQ*]���.�R�VV꣨�T�bd�\$��r7����%߱�=�@������������S��rH��aIf	{��< ���{Jd���^q���v�r=����W�������}2����X'���0���\9���&0[�_ҋJ�%M�sm�9!�(�����=�Q��g��&��!/Ѩ�Sl����9�z�K�ɹ���,"{}0���Z�g�<V������ґ]��^�-:�}�ɗ�ta'�3nL�l��}k$�|t��Ǣ��*Pّ�k�ׅ*����׶�s��>"p�]�[b��++Ͳ�e�_8ʚ�)�طZ�k�/�Y=)�>޻�zp�W�n\%�؅F�ݏ,w1���v�s���ҜOU�qu㏦�a������I�An����T�wͺ��2��W�8�Q��:7?_�;��<�ҭ��N�~4�MxQ/�(|_J�%Q�G
E;��;�+M(�vD���t��l���������)�V�V��=�ey�u��瞼g�y�f<��#ӄF�y�fy��Bc�{�Ke�C"^���ג���(�g[ow\�Uh$P^�{�a�2��oJ;��-�Z��	_ͺ�ep�s]e|Q-�rg|�:��k%��I��-�zt��S#��m�^�?�-�V^�}s���]7n2�z�
ҳ[4��eu�Ǯ�J�AKq���~4���Y���Ӑ^ɖH{[�	�Y��5��V�*u���!��u�u���n�{�eV���ܸp9��}[\�Q��]�r�n���
�n�M������E6嘃ٲմkC7<;�b���g�s���?d��Z�VLM�X9Fϵ�V��ȨM�qƻ:�!���dp�ܛ���^;�&�c�e(�ł�Ix�=+6��	,���t#=���&��9�<���J���d̯,s	��66	����G��J���%��2�ϥ���lEj���N��9�Ng7���`���N��6��푿e!�]��B,���nGs��u��^�bN�f����!*�IAL�R�q��5ֱ,44k���3o3"�朻D��F��{�����XL@���[|�i��	��I�"�J���1�>];�um&>�y�%�f:B�omՐ�V���jMf���k�q�.����5�6Y� ��1Q0��'����Hy��kc{)������g*�Yb�>H�o3F�&z!f����s�����������G���h��||��w�zsŖ��>���z���]����G�&�ԯ_�������y�:�v�<:v��t�1��v�e�����h�1֚껞���L��n9*A�s	]�[hWJB	�j$!P���0n���8@x�i��ˮ)���{���[6M";Ku�e]���9Ό�%���[I�b$��o�̀z��{�4��KY�)j)hA����Ha��[-�&�k����w����K�&X[Y��^L��sWr���P�Z�cp����6d�$�Ƒ'R�[Mպ�0AJ䡛t��γbfB�\�6�m�J��`��]]��e�ά�^q;�:^]���E�HS7ZZ�j��xyÑ&H���1����bi��K3\%-*WlP�]�e���2�Rѻ�'���p����7�g��K���Q�-;�X�]&����ʇ?^�C�@�����X׍���]E	��2�����J�Ml��un�Ta�"���T+���Y��7>]ܫշ6ki(�ͶZ�5v��:�!JT.N�]0�Ւh]\�̽�Q�8)�s�:��w�V	uń�U�ab��.1�]������Kq\7$wѵ��#���ݶ6+�J�ʽ�X�oR�r�Ì�r:h$9�$9�0��ת���xd�'9�	��+CT��Uȃs�&���<Jٍ�6q+��b꺸�BȦ�������1n�\K��5�"���ԀG2�)��t��źOQZ0��FSk�hu��W�S-+m2441�b\bir1�;����屦Yd�Oӧ��f�q����_Z�W%���Ԛ��\M�Rv����x�c����^��6�
��l]IU�`�� Z;.0������Y�>������'A��k)�����k�]ks��e�m�k,	X!wL̳7@�^,)j;qYf� �̧x�nS�f]����,�%^aͻ#vm��]4��ۏ�#���i�պ��mb*�f�z��gk��l�VT�\[hD#��R�]�6kb�
��K��5�o��{6ݴͬ��Q�i�W'VKe{�kr�63��`+��]uٳ6\�nM���y���n�C5%5]�s�b�r�K�aX˦-.p����E�m�5�[4�EuЁ���pBx�p�d隦D����nJ�M���q�P�LC@�6��1�[�9Hƭ��៯M���͔�a*QMsn��Jhv �m4��u�Hy���c*X�#��"[��qEڶʙ۩1�fM�K�uX]՛�fk)�2��ؽ��2�s�:��,��k0#J�hR~�__���x�,b[��ռ�{����H��C^b�(d���j����[Y���0�����y<�}='�~$�F��+|��-�_.�a������򧗟��y3�]�e�W.'���ݟw��߳������!xs۵e�Z��V�Y�l�e���[��d�l��c�f�������z����|<>oEV�5UW,UUT���b��努��ڳUU�UyUZ�UW,UyUZ�b��g�W�^�^�_V*��X���UUn�U{U}*��*�-�^�_U��������A"��T*���J�U`�LnXٜܶ�ۉ�I�������xs���6܅b�5r����1C�f�-�y��g�}���UW+U\�UUr��U��UW%UU�W�WҪ�U�W�U�UV���U�UUr�UZ�ʽ����U�U�b�����U䪯������f��U�U?�c߱�����i�b����FP9Vʪ"\���T�W���g9�{����{��ګꪵW�U�W�W�W�^UV�UZ���U\��U���5U\�U}U�W�U��UW%UV�5Uj�*�j�}Vkur�j�U�璫5UnUUUb�xswB�T�UI
$rQqD�j�E5j�,�ӆt�(��Q�[j���)2���:�n�ZՊ
���j�b�t��L�Z�d���9)Lﳉ��9W'[t[�����7�lֵ̈́%*_���?O���0z�g���>�v{����:�.��=\q�q��L��OI��	0�z��&Ӊ�Gi��mG��S�Z|�I&�x���I$�m��$�O�I�I��8�2��O|�I6�&I'�&�m��i�I��I$�a�I=I��L$�I�N$��ێ$�I4���I�I$�I<O�$�i��M�i�DK��I$�I�I�I��oRI�ǏI'ɴ�z�I�ש��[I�Ye&x�爒z��e��M#m0�0�����$�u�\a�/UW���ݱT��=��E/�Յ�z۵u�.3m�6&Wsb��)k2j+g39������;{;���cRreb�m�����!����\9GUc%����e�emаV�ե�%�˴ls�j�#�b�/�밞����cL��5k��š�4"WC���Z7j�LZ���m�e0k1+�n&��^�{��[�a�v���X뛚�����ȣ(t�i�ڪ���kY`��t6�W]��6)+����)���+,�$"FKW���n�R
e�vIu�x.�����] ��t!6h��Y�hq ��In�e1zVʢ�5�f=f�\4��]t�л�9(�^�����K)v�m^, ʛKv�qJHV�fc%�m�� ��B���Mn�.
�ȗk�t�iNlƖ��3(�ʵ�.�����3Vٝ��f�]Of�ސ�2��u�F�cr�\���R�N�sws��`eݩe�[Jc*�H\	2���Ҙ�'*i5��Q�C�V��F�i���[14l�m#|�&�Ϗ$���\�ď&�g,Vܥ��3P&ZUYA��nUa�Ų󩊥�cX�fס�)��,{f[qU�m1!K��"m1�v)���b��S2�5��1��ô{d�o��]�qI�_!H�>��^��a�+v�:�tp�])��aKF��5sK���eD�����	��y/7L�ݳ�I�@ֆ��@������\F��3mZ��8�.��J�k��M���&�,���gm�v���ʋ�:��6�b����:���1a�fB�V6����0v���8F:�-�u��۞�m���YD��f�4ͪ �T�l��<��ˌ����'ٳs��2��Ժ\e]�ғ�&&�!�k�%�XR�P��sR�ηq-�-u
��/����B��]�d�%�Z�Ѻd�]4�t__J�\�ۛ\m��mu�mm	��ps��������J����A��^�Z׿w��Պ�������}�k^����V*��s��?~�T�Di�d��<��m:�a8�i'I���[�bL�ǙϘ�Z<2��\5k+k����l��h�7&m�v��l��N֕�86�cb"&��in�8+�e]b͆������$���e\D�Se�X�ڗ�VT�Q�؆�G@�f�[�\�.%�k/.����UA��4�cḥ�tm�N�6�*v�K�iuMa���	�v�Z�f��wl���5B��m��� ��c?+�,wH(��eT	�kq�3KD��k
����+�em?����\�0���� C����12_|�(�t�\�pۋ���u��;���k�˗-U7[v0���r��SN����:��WQ�4iY4�����a��&k�i8˒}L%�Z[��0���a������D<�58�Q�(��$,�k���N#]H5�].F�����nH��nH��2����wu>a�?��x�8��i�]N6�I��q�Zu�u�[u����$T|�J�ԓ��|��L�eb�Ix���m��"���#-�.�i�%�>#��T��U����J�*醙b�uos��,��ϲ��!��
(�=������Te��L�P0�
b��7�۴���3��nVx/!�Z`�������������1��$�k,�6�]-uo�@x�@C��hQѾH�/9Fj'9���Fo�I�I��i8�N8�IĒm0~��e��3����][m������ц='R��Vv�۬>i��6�kA6��>��{I��S҂+O~�����cuw(�e��luM�H��4$o�~>���
l)�~���D���Ϲ�a�"���+ϝ[I_"�$>��IH���J¶ڮ�qĬ6�5�Z����7rn*�E�R6�P�I+�mu�>�m��X|�ǚqǝq��N&�&�q$�N~��c}�Jr�>$�I	���!��O���K������5�d"�����[����a�c�Xg5���#�
��v�V�	�a�������9�}��������E�M�ߗw���*Y檚^Y}^�;[q�v�I�V�|�/i�MV�u�ӵ<�q����+�[�[�|�oo�u����:���ն�FXa�&�i�Rq��N&�&�q$<4x�[A�!�N�7�a�@������ę�'z���6u��!�I��R�2A�k���	&����'�Bi՘2�f�C�c-�ZҬåÐк^3.��U�یmB��A�cJ�mjK\̙�f�w���¾w��4�ג�9�2.�l)�B���1kVQ���PkMÜfe�����_5'��=�0a���3�.�w}%q��7R���ޕ�O�_,�k�y�����>��.W��RT|���o��/��}�s��1}M@,�(��w�7��RJđn���-�>�ݥ��6��7�O�ƶ��9�
G�1�a+BJ4������9�O��zz^~�ji�#.��%�]��㙓6GͰ��Zu$�m��'M$㮺�n�_�W���$0���H��2��uݷu.�r\�6�3��c�|j���[RV�f/ݻ��9r-��\O>��M-��q��7�Lc�z���u��LZV���m��U�}��0��ᯮ�â��	�c�gK5�^yjV����|:^<�S�R�H(�	"7��m��L��' �K��}=:t/ �<ع�hc���n���m�ǯIƜq��m��'M$�I6���~�_�c�g���d���n�V=ur�w�鶬竧8����c�x�ɦq��.x+9��ŃD}ں�H�qZ-Oم�����Q��ie������/�u�u�r���뛕6��]$��r�����������i��wgWR�[<{餩+V�<E��ϒ��UU�)^pP9PO9�G ��R$�y�K�y�l�80�C~B�@}W ׁt!��I�={G�z�#7s�\Z�a7Xi�D������
�` ��g���T�s�e�x�h��=6�N�����I0㉤�N$�w��w�c:�W�L��x��y��j��a��}�������H"wn��.M����.�YTt5m����E��.D��2:���LĦP�m;M4�4�*�oI��/�%μ�n���m{|{o�L>e�=Zs������zO����6��X�8h��/>�5<�\��G\���b��j��;-�6���:�O<�6�I$Î&�q8�N'�~�?1��_���ȅL+߽�
�GO:#
͎@F;&�����=b&IE&��aQ�$8�BE�-�,A׋�`P��DU����X����}"[	���y#��|��8�@��]äś"2S�x�+�96z��l�8�8��S��Vfl�f�¶׳@i`��Msz�%��c%i�#F�Q�Ϯ�{k{l�uU
�u렘��jKt�5(i�sZ�:\R��\UIxۉ���Kq��x=<!N{��l��IW�3�J�|����=H|r��R�8�]��-��E�����S���,�B����V�c:m3x���Cn��m�R��OjL�]Z��0'{�S �Ϳpy6�\d7��s�:�q$�y:��J��ȯ;��މę��F߼�앷���I�x��7\�ׄ?N�C���s�ϣ��Ӎ�e����.�z��|���i�ө��i$�q��N'i��UHK�����-8Ӽ�O�8�U���8�g��3��q�}&6�����Y����KŽQ�ջfL�y��Iϟ=b� �eR?5���8��*�i*�JS�$�Dd�s��n|�7%O����l�i�w��|�S�a&6���vQ.u:�V%RJ�\��^p��{'8)��:v�D��fK�ny�I}���]�.L���ؾ8�:��1_Sv�]�r��R��{��f��o3M�#U�1�LG_>i׳Fv����-1���ny~q�b�a���yzy~O'�i��]��z�cO<�^_�o<ŧ������4���O#��i*ө�]N&��nO�<�<�%��F�^S͢�����/ίi�W��yo��������:��<��O=s�����1���<�6�4���0�����o>g�������n����<��O<ǜ_�2��^ޫ�_�i������������?0����/d��������0����Ǘ���mGS�ח���8��_��W�]cO/��c�_�_���G��c�ǖ�˭'^_����Z����~Z�$~_������~_���8�'��̞_�_��<ǜy��^^_��//)��痧���y�������6�m{ao<���av��<�랹o1�e0��mc�/�̒��&Q��y��O���bI��-Ŵ�|��y<����/�/��)䉖W��rQ�_�w��*J�Íj~�����~�[����H��O�d\T�J��?�VQ��|���U)��u��u�����������s{����~ֵ���{=��}�{ݹ�?~�;�kZ���}�5]�k����Ya��_=:�N��q��I:éכy�^uƜ���wln�v��YND���U"��$��L/��c*��>�$����8E`�1��7j��UWD˼�]�Eu�D�#�,}R����UU(��|�ǝ`�v�+;����y�3�WWJ�*�\�R!ĪY*�i-[m$�~Gͬ��P��W��=���+�s(��<���H��K)4ڡ6Y�~s��f��V�<�B�C���1�ޫU�2�Q^�ޤW*pd���T�8��
��E8�]c̯.'�"���#�FPӱ-Z}j���]����-���٨�B�JC��I�K>���Q�+:�"��Q���d��BUW�Z��8�MI�iŪ�r�i8��_�ֹ�]�Y� '<���?I�0��WbT;N-_T|��UŪzMV�b�Z�h�վd��O<�N6�N8�e�N&�u������q"�(��7.�U��"��V�G.�Ir�\���5����(����qk�L�V9uR�����]ec�2�6F�����er��ĹA=y��E9�֨�nȊpY��$l����4Z�S�%��m;FίN��y^�s��y�~���V�\�Ru��Q�_�*�]Z��=��UTh��1Y�n��R%���R�*�iW�I�}ʖ��V�"���,�V����V⬋�b���Q_1��w�[/��S�m��]Y��}��[EV�ʒ��W�M0>J;K�V1��%l�C�5���_�^�Q�6�Uh�"�TT���4�!�^��~̖���L*�G	U�u���KE/�*Lb�|�|�
�*������ȺJ5Է�W�ի�Un�-Eƫ�$�XJ�Q�WV�2�̛~q���\m��u�^[����:�4����b�1�I�����x�]�������3�dj��H4�i�8ĈmXعac{����`�R���O'\k5�3[$뗷w�ڨ�#5����:��f����ׅyW�r����TS����hQ�<�Xp�l ���U4;u��-��#�zŴ��]��.��&��Z��t)�X�S^���8X
۫�y	B6V7�(��A!3�Yג�394v)4�:�f�k�θu�bmv�3��YB�XarQ������sPr�#��Q�V3�+$��(�Sb�f���*a'\��\��*є9�'�j+�-R�*��;.�ͻ&��i���n��'�����]s���Sß��8�!�a<���Vb�E�qZC(���=!���}���GBW?$�ΚS�^���D��勃vZ�H�S'��7	�f,vx�ả�Tf+�R�q��Ee�U5�$d_���*�C���Gm%���"U|a��7P�g���QN� ���_����d��4:}5�'�t��M2�64���k����]�U̚�$<=>�'��y�
���*O0�^E`��z�Uyg�=P��u]n�Eg�����F9'�E0�yH����>E��Y|��I�_���m$�e��n���:ӌ��=_D�	T��J�zN0��Q�+�-�k�abF��۵��\���[�E`�1���_6��F� ~j,��"+�`�E�8b�~��{��ݲ7�7�>��ު�`��:��&1��M㨧_X�@ f��";�D&���Ȧ��0G�X�&�	�WPEg^�99#�Nc .�zn��J�.*�+~��ej�Ee�X$�hV��(��}]|�?f�.\0qkW*R�Eh�k�aCp�+�m)��aY�q(r�Gy����F�Q����U�ga5ls�8b.��U�Nf��n�����D�B�ԑ�d��ZUa��Qu��_���^�Z<���G��Ei)��Z�~�W�.�!�%Un��ұ�&1W�˩N���?S�Z��h��fHZֶY[ύ<�o�θ�m�����m�S�&�c������B�MܺdH��*��$T%Euv��:�wx��>Y�9�Ǒw/����UD��Bݽ6ɚ�M1V��:�irKUBU9Ԗ�K<�]��ک&/��Zu���&_FXi���i~Z�*���n���]��,�����~����d�S�H�UI>�<:� �p�0nm�I�	6�TĹ��2[�!�պ��~E�J��q#��(��u��"a�!��>FOW��t!����A�5*�)��4���%d���\��{]EGYa�X��W����˻�{��]���UmŌ��)�:�X���l'T>!���q�:����*���F*���#�>qg��e?��f����|�<�6���6�I8ˎ�ۮ�\M'�?{��v�긑"�~��5��1�����:��FZЌ�VE/��]�/�Z��'�e�Z�����2xs x	=��d��{1LN��ni#
�u]��Wt�ev7;����Ee��Xe��YVR�EBUH<}a�(w?=����^���P���6��QX#ʔ�VQ�&���eyD�U��UB*��ֱ��ksT��_O	ω�Ƈ�x" ��U���m��u&*���Gy���������X�Q�WT�Fz���j괊�Qʏ;%�|����#s��n����U��-ԪY*���[��4����u�0�����/[x�����'m��q�y��u�i���?}���Lf|���ܑY�ȐF�$-A��V�G.<D���b<�KV6z(��1�&6�a ʌF�qP�͎�%a9��C\+`�X��PA�7j��dRۦDڔ��]ڐI�a��u��w�x�w��QN �;������ja���Tɥ�Zl�]�`�鉱]n�Z�cp�o6l�j��	ޝ쎕��N��qf�yn%5_-��j��6��є}+Z��x�3D��J�<~aZ#ʩE�ģ���ɗ���S�.�0<�G����	���$��>F*WQ�ϫul��F��X[dTi����C�����$c�dD��HJ#���p1N�Z��h��%*#Q�����1�FSm�/�s������x(�(s��u��`l����}Kau]��%rq7���|�����ه��)�j(D	�VTh2�S(o`�VӦ%SgMȸ�x0��~�?�H��G�i����Y(����F^�����,-^RR�d�s��za�^<i�o��?���S�6�I8�i�u�mԷ���.$H�J�T0��c�ol�/�"��:E?E�[�奮���Im�έRS����j�����S�9�I�R>A
N��d����V�U�F�t�*�uT��e:e��.��|�jG]E�̗OA�Ժy�GP�_%IW&)�Z�ͩ��0}c�-�-�,Z�<8@��{<��{i9�-�=��D���y�y�fk)���S&���f�6��I�e]Ic-��M~�[/U���mF�-�a*�c�I�Փh����_aw$]Rnr@����j��Uw=�8f���^�q)Xmm������X?�u�㍶�N8�4�uכu�_����m����$�X"�DtQ��y� C�1��N8����ɺVi
��^Rϑꕪ����9s�q��$�X{�i*���S$��.��(;IG��(|'�Ϟ���{a��؅ᷜ��uFi�
)���ĥ��j�0�J�,-�V>%R#�}����L�qt�Y�ۮ�0�.T��i,Cb�"є6��h�g�d�y4��c���RTa����q�L^"��=Ż�~���j鷺�]>a��o�y*���'ֹ.\����_*�Jq)h酫�El�Jg�-�	��0�[��O�	�Χm��q��N��4�n��Hܹ�$��}�d��>GQW�/�s���>~����(���0�����H�5B8��̽�DjN[--�����L7ԋ�|K�������'gwK�I�HTy���NTD%kra�U��q�8�]w�+ح��#ܟ�/�4�U�y�+��[��i�9ZZ�R����)�]��%��Z����Tq:�Dq�$�WƗO%c�ų�Ɋ�Wu1W-�_��f��|���aԪ���jh�U��+ė�Di��\KJ�IXu�k6�p����#kz�lJu�d�9][--��o�:��/I����<����g�����^_Y~ĵ�b���q�'^^^^^_����y4��8�GS�����#�������+�y����y�:�6����Ǘ��u��-��G��^a_�_�_�_�G��e�����������������Ӭy4�x�4�'�|ǟ<Ǔ���ɵ�h�y~|�yn'_^�m�'�_̼Ǟ[�痷���<������������'�cϞcϗ���6�������%q8�i�:���l[�����1�y<����O<�'�)�'����y:�G���6�n�$yq��x�G��_���������m��1������μͦ^_���W�W����y~y~y~yv��'�����󍳇���0�L'�_�<���_�,/�ȿ:�'�h~moɔ~O���L~H�ԍ�1�k�a8�&^/��y���y:�,	��0�	O@�B�����<�	��D�H�2_���)�S(�݈.��&n�ao0�OR����OG+�Jo{�<KHx�u׉=��oU��&�xFA�������� �d?^�_.=��k�M��||��I�p"���LJ@�+Ֆ��F�G���Z���N��m�l~��y筛�+>�Wx���cB$ӑ���d��g@�������7�B�Z�56����em��XZw��.�F�%uJ�.�/[À3B:��pIM����a�)	t0��RQ���Q�³e���4����a�U٢��F㩍�1����!�{
�R�z��޼5��q�i�ìl�m��K��SB7ƅ<i���<��w�-UiM�����;�$F��ފZ�%��q�.O��[���E"J���{ �RNv=�yq5r�0��E�4N<"0�""�),�]3�S%E+t�*r���g'��{>S���k.��Z��\�'U��dZ�$�n�jV@�r"�	��r�ȃ�S�q���*k�E��i�4���=�^���a4���غ!	����mt
��kJ6�i3�jMj�[�4c�Ȧc,�fb��Y�$u��m�kI�kV�%-s�R���6�܎ʙ�"V�3�Պ�[t�B�X�Ы+}0���b��l�-V��H�Q�ո�1m�ɩ������&e������(Y�Ԏ�gh��ғr�7,�ms��pJ�Z	�f�ɲR椧gS�1�3�a�����b61f�y�ڹ�8��xϙ�m}������w�-}w��՚��s�߹��Z־�{�j�Us�2sw]�|�5U����ɇXe��<|��u�]N8�i$㉤�u:�6���'�vnL֑��1�c����0)�.34sp����-��Ty��[lm�+M�Mkq�Q�Y@5?W;�5���U(W�uJ�F�Fk,�m��	�?���hN����X���]k���c�-4Z�j�`�qX��v�ٛY�Vѵ�j�	k��c���g�-�Ƥ���ݖX��s�.�n���,7���;QE�!�lKi=�5%��ل�ŀTV�mq���8�����1[�'C�ڼQI�/��K������yr��|�9P��K ����Fֶ_����b\��#����i����kA����0�O�&j��������F��ܹ���8�][�[�m�S�j�i����8��~��8bc-u��l��?L�O�0�ݜ�"Ux�7u��떹>c�$�9$��q�u��|���%/U�����G��D���+e�K!k_Jy�L9�`�2���BO�H���ց��$Qħ��"��k2Z���yJm��n�-�cx�:��|�[M��������]u�mԓ�&�m�]x�u���Lc1"J!*!8���Y��E���,㎰a)\&����r�=k�K>J��DE0o5�|�u���,1T��lj�I�J��u���,��O0�Iy�?E{7U_��r�����zKv���(���3�õ���ś�����ӕdE�m���l�~A�R���Ї�����M��7:��`�aU��ّ0ך:P�R1�!��o!~Y�����1����˭�+�̩��e�Gp�EkX�챜g1#�i)㖦��-�$]VjV�е��N��T��Z�c)k��0����D{���3)ڑ�[���|�:㮺㍶�I�I6�0�n�m\����.��b$ID.�`�R8�'է>k��ܻ�~>��!ao!�i��ޫ3k~yn#��u���\b=���0�U�ٳ2��Hbs�����<�WP�G�|���Í0�����K�#�8Ԑ��58ڈй���6��ٹk[j��Q~�V�u,���-�&��_�w|dp�\[+H�����G7S)wwa*���+#�F�I�*�C��(�(�`�˪d��y-lvZ�}1��.���O��	׉9����j?%8����uH���a�wn�Jٻ�FҴ�[��"F����k|�o�>y~q��q��I8�i&�N�M��}��1��܆�9����?Yu���m)��h�������k��`� �<߿����>�=��YDU��B4�Ktk��̕��&���=J��K�&��Ѵ#��i]�2����9�a��� �d��&�������C������ʎ_�\��>�,���#�Z0nN?�����Z:s���O��kWw�A���.���
���ɧZyH~��?$�g7n.;ÞM���$-b��[H����Yͥ]V\�s����<�xW�Y؏˥Y��|����ԑ���m��"��K|��'��]N6۩'M$ۉ�c�G�|�
���R�G"(�#����l�wYx�1bir�K�+�*4[�$�-�9��a9�����l2U+�6\P�U��m޳�-����넀LI���"e���FUvɱ��nm�˴�[\muG�&s�ݶ�dٸ�4�}E����FU��1ٴ`�i��f��J�u����` g.�ji����Kp���~�7zl�k=]Y8|�SDiV*֌�oM��K�8�O=X��;�'D�:<>A�(r���W�{e����{�gu�d��#�I־�xt�/?�xs�<��[e��?A՜~e�/ʎw�IV��[-*�����!h����؍R#�o��*��q��-)l��L��G�<!�N[>[|����Y�X�0'f7�]uQaR:YZk��5���NC����W�L|�, ��Icr�%4�t�j7[[���h�l�Dy��[l�4�\q�]I��I8�i'L:�M��9݈��xtOD�ч�	*߈r��?&}sn�U�ߘg��Q]S'h�����a�y�qUտkȗv��2�Բ�U�c���9��ۓt�""֯�[�R��N���|�}Skbl�uSa��[qn-o�]TAi��S߉l��]߮�Z�w����c&#�ZGt<�=��a#IpCYkY�1�*��kn����ќm���خ��2!���<�/ϙc�nK�J���c��8�j����_���0z�����J[_d�|���G��.O8˟-�Z�m����q�κ�m��q��u�]<�n�R��UU��"D�C��a��k92C��i._�i�0!��������h�Y�-�[iJ�O_���U���~�b�>q��vL�J��cdw�K1�V�:�~v�s�����)ɷ�&��Tr)Q/�2�70����B�\hR����'�˵t�s%Ӹa�VH���e��m��ߩr^3��O�����b�f�v�f�yne9F���v>���JSsr�%���ӊ����%�/�����~�!'9��{�uN���gw���k|���_'8(x�w��!�(#���XppP2�P���W	,�d[U��q��U�}!Ϝ���~r��sI��6�|�cX��ϩʼհV�+ַiտT����+�-k[�����ۮ?<�I�]I�I8���k��sX��H��l�ܒ꡺��֪%�ܻ˕�n4ن�R�H�Z0���>��K�"#���(!��rGq#���a�tg��8����^Yo-�1���8S��=�:}(]a.�9�������a�k����]�������p�f��?>b�D]Z��2�Ye�Z��6�0��W�]ݮ��~z�V�}H��6Ðp�V�ɮK�#��&����ؗs�40r�Tz�-�O��?2�YV��E��U���u��a��e�h��W�~�'�R���Ix~v[O�q������4������|���8�Τ�uԜq&Ӊ}<>�����$�mE.�1)�K��_𢆩=ǘ�I��;�p�!{uȯ�B��m��ryǡ����k��v�&��$�z�:����<W��s盦�#�v���nd�Y�������̥��.��N])+����-��3�q"�5q�E����:�]�
� �mn���]R��n�3� m[F�W=U�שm��f�Ĺ�I$ÎS�=')��?�^s�^'��uYo���r��mVo7U˛�b��a��>|��V���_�����4��ś�-�0�J�0c��ˈ�ӿ�����q��Z�]8�h������KT7m�*��-�ܘm�/��Z�]��N��T�Ty�i���y.�f������0�ص`��R_9~|��2�"v|#��Y��<"�)��W[�q_����B>G�p��jZ6I*D�%�:Y��ŗ�@)�#�9��O����nلj�s�~q�|yg�$]6�#�ޜ�&3�3�%i�GQ��m�[��[�8��:�:�N8�iĎ���f��0Ī�L"�kvmoǗ]E><�����N1�,�%u�]?<�a����Z�?y�_S>�.�e�m��4��JNO����9_Su1����qﾭ�����Gͭ�����6�ˬ�IG����~Z�o�E�-����Ib��oyO>r�i\!��W���@C���)�kn���7�+�R��,�l,�KJ@�1�9�zC�S_�B4��u�M��/�ǖ�Ҟ|�iȈ���ݲ�V�-dqHa8P��S�Y�ڼq���蓆ѧ�o�R�Q�?&�̘������_��q����u�������2�'�<Ϟ_�_S�/��W�W��y��6���G��y��O'�$�q{O�ϗh�G�c�-����>^�/\���y:��%��.'�ɗ|Ϙe�<�<��"��/�/�\������y0�O<�yzu�4�x�&��/Ϟc����V�˷�y�'�y�|����N������eyy~y~y~m~yo'�_�i�|���~O?:����?/.�?3����<�y~O#�|�'$�e~u}N�s������y�X��<�4����e<��K�m��:�F���O&�o.%����~O-~O#������u~M���������y�<�_�_�̲�Y_���W����y�������K|�~iv��y��0�<��H������O�^_�����-?&ߗ������i�#���ߘ_���2��\�����N��$��D��S09\��_E7J�7����M��X+�������f�<=<�u�s�m�b�|��"�B�*���U������_���|��k���ʯ*�v��w�ֵ�w��ʫ�����Zֻ���UyUs���a�Ye��_>u�]q�]u$㮤�6�u�δ�$��Vsh�uXF�x!���vYe�|$��y�N�U8qʘs��8ˋ]Vv�FX�z�]i�G�r�&�u�_nK��)�W��|�,#��b��x<HT|�pk�u��5�ˍ�.��H��l0k���Լa�֕�Uukz���ql�)�Y<1�"a>	���VB�D3�!0eꫥqF;��WX��*�|˫|���D�{�w[e�-��L�բ*�����}Vӕl��qsl�C��%��9P�)yx#�JC�:PD�!
b�u�q��I8뮤�M�t�:��=1�D��g��R"9�#�yu�7W���Ļ��?TiJv�Q���gek����l<�j"|��f��i�;�N��T�6혐���a��~�u ����5�Q���ea��j��ϑ��Gg��|��5�v�6��T�*�Dv����1\yo#�H���g��C�F?0��8����&�럟RVpÝ[T����a��%V+�I�ꇟ�O���,�ea9��9�'��p��FR�D|c�V��߾Mem*X�O'�q~�� DDv��qwxn�m�a��ַ[[��L���'RN:뮧N8망|�w7x��M�^��j3+�>��i�\-�H�j(��4�0��,\$4�GخA���ҹ�zBөM�5�ç<<ǈ��ӤM�LE����U����~�m��jD�GL�΀M]�2��j�ƙ���{U��\��`�f��{���^�/�/����I�!IM�A"�d�
�R���@���U֮laɶ�2�����k����*y��tO���'�~%Z+�Dz�qĝ�>���wD^%e�<��m˪�eQ��m����*�׿$��ծZ?>|��c��k�����D~�Ji��F��Z[�n�����e�V�I��S.��R4�H�����|�"��FNG�&�燜��|�����J��%EDDe��^v��ua��K[h�K�EZ!���zI���)Y��s%ڪL]���-�j��A��x���-�^a��[m.�He""�h����jW:�������Z<��Z[+Z�mo�8��m��^u�\u�]N$�q#��{�g�s��U$�S1U��n(\-p}Wkn�v�wC���u��nm�u�+�cn'[��&园�ݭ�;Y�eu�,oҕ�OC��x�����uʯ�7_DJq~o�a�c\��9~]}QP�7S̙���`�Nn���.b1��3_�R�#����գ>;e�-� Բ���jV��5�iBQ�[5 5 ũ!�J��l��mm��!+8��Bq�AdFFF{��ezt��m����#�~O����j#�{��X��V�(X�9�²�(r���[A�*�K/�����܂�T��[kM����sw1(;8׆0�Ye%b�1�ƴ������B:f����-X�֧�����E<Q�8G\/�iO�*cU�/�%����7L?6��ב�8=�=�,�X�Zz�9�y>0�u��(����q@;+ؓ���)��R0BIÿ'���{;��J]����9U*�QU�dJ��b.�.�"6�n�:��Y�3��J�5���\�Z\�1$��y�>Gԅ�˓n�zMV|�ֻ|��FOu�~��ł�KA^3���K�����,y���P��hm�	j'������LQ���4�`��)��,���'���<������57*u�����f%W�Nė#�<���oRVZ4�YOYi�q���'RN:뮧N8���5���y�p���*���&W�b��yRF.c�u�l�"7Y��S����?>Y�Vѻ]4�.�/̫u|��������D��I��5��%Y��]?&j*�/��f�؛{[��]BTP�	F6�\�Fͬ�d�ܐW������'7%S�������v����Hw�H��Ը�/�M\��D";��;&��Dh�9������w$�i�M~\����|�R�ugQ��>���H�V}���+��_f�r���d���-J��$��a)�f��Q2�/e�Ϳ�q���'u�S�'GS���c����].���_�����b���/��i)h��i.���qf�E�"?k�>h>%�Pa��w���Y,���l��S��4�w�I�?!�;�,���
��|Yy�98�
!�ǥ��T~�d�&�S�;F��U]����g+�#g#dTmu_XFaԦZ��ֻ�h����wM��aF�[z��v�a�]4�ijmJ�G��"yd��ڨ�d��P�*Ҽ��#h���9R�E�ku���ǖ���:�8뮺�'GS��#��,�?����|���,%a3��m.�.�66Ř�m=l��p\��Ybm��B��74��o�{�08;5�(ނ��͒���\&ؕd��,>�z�Z�J���Ā]M��]����G��bO�^���VI�Xұt�TuٱŚ��jB�4�T�qu�Mv3)n��I[�^t������'�a��	Q�inT0��U�%}��C��er2�1d���������0}���s�[�^����t����^�d�Os��.�-l\��Z4y��殽H���'�}�/=4<�|��HH���VB#Q�b�Wܕ�.�e����"̣��a�=�"G$���W��9ߺ��v�h�$�1;�Z��F�Dz��`���?���eᓆ*�EJ6��c
�j2���y�w�~��^KD���]WR�Ci�a�^s��[mUDmZ��+|����i�]I8뮺뎤�H�|�����ĉ)V����Vҫ�k�[U�}X�����=�b㯚Z�����y�x<�[G�����?I�^���H�4�y�w��K��%���>mj�}�D�%-�V5����������C�v�i��2��T���.�
�e����K[��G�-x�9�.��-�"���:�8DZY]m1�p{�L�q��2��K�׫/>}*�3F���_�3��s9���A��^_1r|a�>�]��q���쟚u��]��9^[>F����>m��6�q�I�]u:�Iđ�_:�|ĳ��)W*K�ĉ)�˦�{��c���}�6�x�y���R��VҺ���]G�vO?7�~��Ŧo+O�ש��aڊ�K��V���;�OǙ���K����6RYk������y�uXG�\�6����aZJ�<�f�{Z7!Lc�r��'��Ydk)f^8�|#�*�G�Yc��u~����}S���[���W*���i�����x�m�M���'̵_U��}�9�DZ����p���j�d��>Ji�0�Ӎ3K��VҙZֶ�[���[�o�6�8뮧]u'G]|���Qx"&�����!����X�e��ݴ�Õ��J#�b�J2�g�'�U�v8��M�l+nW6�Յ�D����~����OL&��_�\��(�W���j$m�L���>2�Gͬ�m�W�~a�m\�`�S��qlbsw����VJ��>��^4�٪�n��Zj��E��/�3WVi^e������D3ꜯ9&��%ɉ>���-�����H�ͱ[mg���xګ��i��|�n���8�l��:��uש$�i2�L'�&�I6�x�'m����L��8���6�I���$�<q0�$�I�Q$�m'	&�I�̢z�z��M��0�ē��q�q��m&SԒO�I&SI'�6�I�G]u֞:뮶��x�8�ԓ)��|�$�'�6�I���L�2��|�ON&�ĒI$�I�x��e$�I$�e$��ׯQ$e�Qa'���I���	�RO_8�q�]m�׎�é���Ra�=����#����3d����0�o�&&V���a���q"-5qY6��S
s3H%��dȀ����<fF�Zf!�0U۝��q�C/�y��CYkC��ֿQE�j$�`�ē!���BKڝ��I'�.��7<�$lnT��¯�mw���=�x��ڙ���%�Rڍ��ҚyE2�l�A[F�K.�}yx铩���&m�}�q���
��P�7�4���(��r�q	�*`�*Z6��0�lYNT .��,�KPNE�Y0�_t@ˡ";�3�㙯�Z �D��F�F��f��(-�ǉَpŴPY���-��92�0�Hp-��kL����3U�U!�-������5!�=�v�B=ɾ�<������x|�q�i:i����Z�^��F���>I�J)7��<5*J��������$�� �$2Z�q���N(\�|�_�+)�^<g�]5��H�<Qt+����*ǆ��>�%r=i�O��=}� j5����B�j��n���ǻ�:3$�hًű�v�]�*��-�ԭI���\�M��V�m��&�	���f.��Ж�na��jrƳge��C`���-��ZZ�f�#�(�fR�(�cQ��u��[@��gc[tWY\605�S�	��&ַU.�,i40�(�GlL�em���ҙ��;
�[Z3k���[�:=�`ݾ9�m��4��h��@�m��,���A��_��>Ͽ|��{����߼|~�Zֻ�������;ac�ֵ��}�j�j��{��ַϖ���<�o8��:�u�S����#��O���g��[
�.�U&q�X�@]ojz�oI�ԙ�v�&�V��j,f%�e�Yc��c+��Mn�hX[u�F-���M�Z�ur��"]+�&��C]�4�����7��l1]	S�7Sl�,t�ДDnuabK8�|��d�G�Y4421l��m��[�艬��̮���cH͡[.3g�������|�5D֖I�l�֬�ۗ#M�K��B��CZ��������:i�s�jE�Ǉ>�<��e�����uk�\�i��\IL��)�1Q�n��3�����(|�#�a{�*LJ�U�e��./�9%��v�+�N�iT��n7�Ĺ����Q���8�ثE�Ԕ�:���������nvrt7���!�#IUd����4�q�[n,�χ�?M����h\�~{OiXy�.��y݋.ֲ�,�����}H�d��q,���{����U�	pđ�*�#��ַ[���:��n��N��u�]N$�u�}��%"3Q�[b�C�m���>�s���|�ub���Ǒ�]\5zw����H}��7���H��L.�����~nL=X]e+l�R2ɄU��*�W��m~֜qu]#uF��˼��1ƽ�/�"T���"�>ZߗWO��0�H�w<�����C8�����f�S8[8l뫤ii�6�r���'��;�2C�9�	��a! �;�=�*>G{���q)��4�}�m��kC�����b�0���qΥ���Ԗ��խ�#O�u<u�u�Ruԝu�S�'^|�߿a�oQ"JD"q�̥#���7��}�2I����+ޫu����F�];_�'�Q[G�Ke��m�&ȏ�J��{�X���*"V�ە��6��o�;X�P����<��ċ�E���^����]w+�mı�������Kn�>G�~G]G�W��\C(s���|����t�եJ";�G��n��˯��mr���߽$�o���H�.�z��1r�$��G㫤C?$[�F�n�M�w��[hq�%���J�>C�&�e��j?W��]Z������y��0F�y|�<8�n��N�����q$믝~�"D��k�6�['�;��x�o�Y#�VZ4�1uR���_jB���!�������Z�EVjE���;�\V�)��J�r*��Z���ҕm6�h�qku�0u����j��־��un�?ZZ_��Ϫ���qyh�+������ai��������Tqeu�TFQ)�&E�3)�|�W�H�P��(�r���1})����"KaƖ��C�-ڔ����cՋ�s�m���|�-�J��+H�8�Ȕ�KZ7Q�F�V���e�:��8�o8����:㮺�ϝz��"�]ż��w�t��=��CbO	����ئ��0LK&�M��D���c��Z�+�ϳG�Iu"��<M�Rg�X�-%��Mrс���:P�hM�K�[�Y$51���r����lL5�9��x簷͙����D�u���y�5�[7G [�3}���3#r��A���mf\���u�e�M������[�WK3N~���OF��<��a_%u!��%F�%����������>a0�5�1�~���qm�Uj�2����^9��s�>��:�%V�N0�G��.��[Ky۫��%�K,�0Sp��a�
<�<���~Ͳ���I�2�b�տ7_V������mu�d�
�ɳ�����a�~�Ȟ%gڶr�.����z�1�eb�s�x��2�[���H|���>�'�i�!�SJG�E�����o�$�,Nǌ�s�u�zR��JtO���6�:�u']u�\Iמ|����ĉ)�J�6�F�hi6����	Y���9�4�4�ִ���\��u#IYF���[,�����LC���b�����#n.��尊�7��m)zJDs�%�~Cn��n�W+���=in�S���$��b�v��g��b�11*�u���La�+9iW��t���{�/,~[k�<(C�Oh����	����X����}G��}X�L<������W�s�r��x�)�xcߧ�� �nY�Eq����:���H��Oq��q�S��뮺�'^|�����|�|�c(Ƴ��$IH�#{��a�+�6�|g�umB�+�Y�3]�u���&)�e�.�xC�O�O??'�v�h=��:��4��]F5��4����� h"������-��yE����	I��_D�rp�O�Hz<�Ϛ"���a����a��%��H�q'�2��Y��g��k�ةRJ�_'??h�x*"�&�o��O�����|>N��T0
��gj,�Y��������^E��쿱u��D�z���N�߲�h�?��j���k��g���/	�E��j�w����}��kq�����(��o<��6��']I�]u�N��-k�1�1�DS�=:S������XZ��s�ڵq����S5��JZ��\�{�p���.�V���`�����ВV��8�w����-_��?	�Sz���ı�����A�~�u������߫O2���~��.�wu�+������!�b��4a�ߒܘH��&�8�!���J|�m�eߤ�`�8�yű^�����b#-Z3�V+Z|��'�����[>F�8��<㍶�<�:�uԒu�ɝsx���c�|�����������:���Ж��JWlW:�F�>�m~|+uc�^�9|�b�;v�x�Q��AH��R�f�B�Zƃ)�P��KR�q1����]h�+�vRe�˫�u[�,p��i�XO�QE���_"Fw¯���R���b�X09�Kh8�Tڴ,�0*��Ԃ3Mb����vEfh=�d��}KGαL����K´�8�e#<���>u�8��q��kW%���4P�_7E�P-�kи�qþ���W/�j�>;[}X4�a�bK�z�afx���c�ܒ��J��iUθ����o&))Qq�[|�g���wؚp��mj�;��:ikr������~���;3�g��Y�n�fjb�Kv��OI����%⼔˚���,�-����b�>�9�$����_-l0�6�םx�6ۮ:뮤��RI�_:�_f$IH�حV�0�����w�l>W�U���r5l^+GiۮG�]|�^���'�㈍2�d�ħҌB��7Y�2��2�lVkKoISֺ��N6�����d���4�G�F��%�[�q�Ea�'o���m��|<�����Z.��*$�3]���K���S��)��!�(��5�~���&V��zSu)��n����5Dz�H�a��8����+4���-��.8�O�q�zۮ8�:��]O�I�D�&$�IĜq�8�e����"i2���֙I8�'�q��Ğ��$�M2�&RM��$�i'���O�|���_$�ORe'm��M��$�$���I�I'�4�I>I'�Ri:�u�S)��oI%��0�OQ$�$�&�I6�4�"<I��|i$��I��$�qL��^�I&�I$�ğ>|��$���"L$�RL�z�i����:Ç]L��,�����0���7�˒�t�~��1
�F�\?(�ެ舄O��w���T��4�[�;������O{��{���u�k��{����s�붵�w��sU_U�s�G���>GϞy�q��yǝuԝu:�I:������{�0�?"$e�������[\�za�0��f���b��:LUm��&�e���k���q����C[H�H{Ģ	���O�o�I	����jh�Z���"�]Qt.F3I�m�4�Oy��$<��[Y�#u��SMrRo�yJ�1�K��ɔn���ޟ4��fK�j���i�%ݧ��>��-iUh�W��mĦت�8����[_}�.ֶYZ��#��q��q��q�y�^yמu�]y�οVq$�A��l���ĤB@�`���C9����>q�N%V9^���b�W9���-����_~N�!c��+�Ti��\�H�n]*l���n}'=�|>�U�9D�~�������}�-"�)�_/��rGO���p�m�	�:î�#��vc���=��Fw�ţ��| ���������Β�}-��^s%˹_�U��#���9��k,6�3�o5_�6�}\-�����4����O�mǙq��m�y�]y�y�]u�:�sW130����e@�)�⎵e�"eE�zѴ
��k?��M����,��{;Y#�(�8�DR�	'Ak��[J	Hє��䚱�%�.t�-�́aȓ7+f\YKl&eƗgI7��gzٍk����,�Xmj�����]��l��]Ɍ���:��8�q��*�o������Um������%�=�����h�7�i����'͵Q�p���C=�:x@����+^?��O�G��2���.6�e���fM>m���J]ܴ���2�TGm�e�ۤp�;���F�HT��*�L⦒��(F����cIx��Lqד�O��-E��Q���>Z�<i��6��6�n�]I:�<��ϝw��ىR#��ۍ�s�e�ݙ��W���zBͣL9�q��7��2�&3�7.��#�@G����W`��!S�u�������g�N�uw:�>aI}��{|za�k�ƥ�c�縪rS�]��5���W�i��#�j뚓�&$���.�0�~K��n�T�O�Qʎ��`�C�1w���jM)�1mĳL�h��lQ�츨���%���ۣ���rQ��`�G�xSӿ���?����?y�O�ї��m���5��ӆњ�e��Ixe���[mka�\[���e�m�S���u�]u$멥�Q��x��bD����MWݒ|���������4��"���sl�u֌#��5?5w�a$�گ�8|��N�ZOk�R�&ܭ!�w	#��c��}���=�r���]0�Z �`ͮ�8�����<h���?���/��I)1����0���5�˻�4���0�~&�4�u�؇y�U7��#�����bI��~i���=�+���Vܹ#����qdE��מ�g}�u�*�uki�_-����2�6۩�RN�㮺�u���a"JDyƚw���1��q��8u�n�z�MV��S��G��1���ߦu'�c��{������S�^��5����ԗ#U�?��O���?��W��c0��f�fb�	oN���V�4�)�(�E������p�����q��j����@�i�BhkI1�7���+%�4VQ�s��;�ͻX����(�m!�žik|�M-��?:ˎ8�n��I�\u�]I�SNov�đ�T�.**rʯ�
�I2�}g��|Rz�MR�J�ʔէ��­��c���nf�3���iOAA��5��g�ͪy����,]C)aAZ\�٭b���U��f8���F����2�gMD�ل+c?x�/O9�|E�a�̊٤�S&���˨%F����Άs�QE�ݱD."�R�Y��6�e�=�*����$�����^��o�iwx�'ur��I��4�yןW_4�a�m�m��9x�\�fK���e�O���2���)��'����x���e����}�+��R2����۬c��O��X��^���5���{+�1i�ۆ�Nj׻vY�))oB��X��Y���XH�is&�~!H}8�~�e��������{Ķ#,�4�q��Yz���_6뎽q�mԜu:��<��<��:��7$���mV�&+L=[W�S��wq"ki�b��<�[n2�e���X�o�u^{ɺ�[xZ��g����Q�!%~{��.Y󌱄�u]}*W�S.2�Vݓ���>���K3�R���f%�j���G.�F4�qE$����%���ww2gؓM<��3k��n�V��y�����~a[k~���ҦZqu�k����Z�0�k|�n���m�Rmԝu�]u�S���g���QE��:z�)���m�4ӊ�-�чk�"=_jJ��S�H%G��G#1�e$0^ �;�>�>��|2'��/e�qh�It6Y���զ&VVe�َ���\ork���ZY��H���l�'f%cĩ�l>]l��+đ����&=|��!�i�R��M�{�M<�e�~�"lˍ=\G�����,�x�L�u���q��I�S�<��<�μ�-��>�IR{�^��Ԗ�a�_�a��2W��l��F �}^D'�!���m� �i!Zbn*��/P˛X�*��qPHA�c�|I�<(�s�zJ���&*}r�Mm�Ͳɦ}޹O��J|���)�>��yj�9U����)O�ӕ����?%�&�|a�r�W���ҿ':�o˚���6�f�f���j����.UP�m>q��8��|�8�o�u�ˮ�u�SI'�L�I4�6��x�'i����L����RN'����a6�$�=I>I��I6�OO�$�I���x�i&�M2�&RI6m��m��I2�I<I��OS���$�I����&Ӊ�]u�u���]I$�L�a$�'�6�$������RI�I��ē)&I�I�Ye$�ԒI$�'ϟ=z�&Yd��	<e��x��e4�I��a��o����y�u�:���>�b�13;��1K:ޤկvʘg��'��aӳW-�7�B)�4�D}�����m��ʃ9����YH.�����Bp��#Po*��w �4��eH�)ݙ�;\SY��Ӹ&�����!�*K�8�M��Q�qg�]���xlA�9D���zz�����Z9��>�{Gڇ���M*�l�÷�v:jj��h�%f(�:G�����NuG�a[y��˝>��!�fB�pƑQV�Z��3��-��[tF�&zR�=:X��Kq��T��4D��n�g�:��篝Y����P;r�6i%��<V��-�tgA�-W�"�cy�{3r�J�ev�N�*L��t�憱B�x�S�<${�A��d���i�BD�]�v��Z�늖I��D�6+���p6^p�[]Lg޾���f�)��YE%D�i�/)JPz�V�'j�`f6�9�gxA��T�=ͷ�cg���"%A���ANJ�=7�R�[_e�{�b�X��U�Q6��J�c�a�Y�뵬.�e����֠�)��,�͔�Q�ԹÄ�I��6h�BMQ�Y4V�T�SX���v�Qv����&�29r�Y͙1�:9�ꫛ.��hi�Vi|��}��M�%)�	���j��xn4(@���k��E�:�۠$��S,ы+3iu��l�1;;ڕ�tν�q���5F�&R%Δ��`̣]B����&x���h'{�k�I6Ŀ�������|�wU�\�:�>�����qUV���]��}����*��s��u�_<|��κ�>q��u&�I�\u�]u?����݋T}Fa_��a�ԼI�5��B]��\�z�pMM��2��-��B��AQMBٚG+�F)���a$�\�����Ɓ6e��֦&�)�Z��/�6Ì���,k���6�v�Y�K@!f,�W8��v�BM�����Jl#a5�;0$"5F]�)���!Lm.!.��M[lf!��k����l��Iܒ۟��(%�^ԲUv�M#���mZh6Ŋ�s5�d
*�sm�#�1ɚ��pm,H�%�I-ۓ����㌲�|��{x��,�!�Ӆ��sIo���'�=��Gƚ�����3v�K����������}�'r��x�O��כe�6�t��3rض"b�'����#�<������f��ܶw�^@X���+�n�l�,K��%IǸ��v���\|����k�r$�S�ܓ
�+[,>uo�m��8�m��n��:뮺�u4���������[m�s꟰ˎ���]�ܽ�7�m�T!�릏���1<�2�ߙ��F�>x�eH��~���bN���p���]�'�[�{0��>~Z�m���|��9���m%W��fF](�����g3T�b	�x�����[�~��&\m�-�ϫ�w�+�յ\q$t�V��I<�?�9��?���k-mT����䮢8�L�����_-���<��m�Rmԝu�]u�Ru47+�K1���"B=;�5X|�SN?|�,%�\OD�JtN���邀�̭E��Y�/>::(������==H�$��ז?yԻf����<Z�����4b�d�I�$>n'�#.��I�T�~]��v̵�������JqXsu&�'��[�>m����H�|��������8�c2��M���8���Ma�,���M2���q�6۩��N�㮺�I����ȑ!�L=Zq��H�N>�Zp�K�C�ǟ�c�}�Ć$kG�C��fk`E�f���d1�%�mL�Ox��~^��x����0e��޷�)"{?�oV��c-�Ի�峤��_U�^����q�70�.I?W����V^闓�F�u�t�Z�)�HƖ�|�ϙT>p�2��%ϱ't۸�L~�F�򴵭�yo�u�|㍶�'N�㮺�u:�Z���Ǿ�8R��k���_�ѯ��㼝�j��PpPS[yJQO�ޙO���O'�i-�Sj���,؟pw��	0ntL�)i�n�(��Y��������Bh�0��������QA.��-�Y��rG44D*�H�[]�T@Ձp�T퇗m6.�fgyϾ����V��|
}4g9D�I\*��%���;	�2�f߭��գ��q.VR��e����j�V���U$�w��K��R�G�Vq�����~�K�|��c�ʶ�2}�d��yO}X_�����_d%&gSZ���0x���L�%!��ۛ��֗��lVȯ��y��L�=���a�c��L8�)�����u8��m��q�]u�]u<��:�~�"B3[q�~~��M=����K�1Q��~m8i��,�-��yl�j��Tb$w8�Q�i�$f�6�������2�$_�����<�x��u�[ĞkS�����k�9}+�=�z��?�\[/��h#��m)���#m��V�������T��]uu�k��/p�b�K����ᄭi8��n]�_�{��s	"����$�b���m���|��4뮸�N6۩�q��:��^u֜�����=����$#���~s7_K��v�M�j���o[䯍-n�O�O�yr�]~�7Y�N����rN�}[���F�D��)��b e�����Yy �`+�hٶ��Jfg��b%q���)�i�h����Ng��K^n��P��禘J�ϻ�.���������"q+�v%k^z��A��jjD����E1%��O��A���|�z��E����Y��8�l;��%�J��f��.���2�����z�L��C��ؾm�:{�{��F�E�l��5��>����_^�|�<�]��+^<��3��5��A+��c_���:&�q�D>��ΕQ���A�Yu$]r��T�AG����~y�k,�}fs���� D�k��&�ou�4%���W6{��J�Y��_'z;MZd�Y�1�.Lu�~ޞ�v�l�^,/^	o[Ҽ�,�]�e�.��u�%x����߾�����|��ױz�Ca00�<��!������.mK̰��e-�g:@�2s�ZׄkX��G1
��BgU	�3����2�-g9�2Q���(
s��^u+ �t�9$9A8��!{9\�3v��{19Uf-]�.��36��y"�ɖԜd�䰭�<>|�3i%m���a�Zm�q�������l�t�e��l0��|ۮ:�8�n�����뮧]u&��;9ŒQF�RU���a��Ւ�ҧ#m�1����9�jm�ۯgY��ΐ�b(�oRI��+���_V��/� <�уA�Ї���N$�O�f2�}[ǯ���7�(&���cR)k9���O�������zCnW�ڤ�$��ʒ�L:��ӆ��k��N��~�}�1xTy�Z��g�K��������+�A�(|U���F��~�zm�����\����5�&�G��Wq>Z�0˫|ۮ:�8�n���u�]u���ӧ�Q��'����kK��-���/�� ��Qļฮ�!����杧�E��A��+0��D���M��D�V��iE^��-.r�Ĺ����`1�&a�#It�f:�T���У6�k�{UPH�$�[n�u��n�r!F�-�4�!Q-R큲͕j�w,"�Q�!�X�~��p��OA/O������1�����Ğ0���D~nI�8۳�KŽVG�ZK�>r�ru����=9�s�>扟�)�F�$�(y��w�J�a��ܒ睒�Un��V�y�ǧO�����|�^e�i�G����riyrgk�a2I�'�j����3���I������]���a>iŭ�F�$�qƛm�S��:㮺�y�:�S��I$#-6���̣�'Cp�㧑q����?�2O�nn�s��3���_��J���ov�˼\�n?u���$������e�"Ɓ�u-��$��xAT"S%�R�n�S�NĘb�Ɯ�1�i��.\��n4q�em�y��b~�R���<�_3ȶk�%u��ϐ��/�s�Y��<��}4����<��8�>m��G�yy䓉�$�>I��M�x�'x����I�z�|�����m�#��RI��'�>I2�i2�h�M�I�8�e<I4�q��e$�f�i��l��I��<L$�I$���ORI$����IĒI�N0뮺�u�[u�I&Rz�I6�$�����	��ƒO	$�$�i&<e�I$�I$�����̽D�,����f'�I6�=x�i����$É��:ˮ���y�Xx��J��uE�g�Ӝ�wL�Ii-���*�Rڶ���9��+jt����w�#ЯEnQ���wj�$����n�L��*��\S���9J7[j��g,�v���6��:��f����6x�[n��L��Kgu�����/�e��g|(r�����sǛ��Y[l�IMF��lC�IF"�����z�}��߿���?�*��s��q�����{�UZ�s��7��w��z��U�s���.��珘|��]u�m��O��$뎼�<��bI!)��>E����Z䶍6i+��+�\��/��ܸ�מ\�3��i�����<�5�$f����{�>+~��;�ĩ8���Ή�f�l��k���'��9O�����Ǐ�a��>+�4i�u��e��c>Ů�ǜ0�vr�Z8���I6a����y�rf�úK�ؐ����ո��Z�0�>m��8�m��|�q'\u�]y�|�z�d��2�x�8���<���F�@�h֬o�4���R�<�.�](���a�����b�Ԏ*��D��>��@�jϞA�2};�S���=E���Cxj�����l�)�7k�q���5� P�g _wh?��,t��5/����j�&��s�m-��m=X}�����u��ݪ�8�ki�|�6�q��m�S��:㮾�â�t�IIN)�0Wa*�sw=�H��Ԫ�Dh�e)B��\D��И���o8e��Ж��Ǔ|����6�۪Nbm-5ir9ff��!�GU�������ڵf���8d�F���U���&k����v��ŉv�)2�m-���"��Ap�h��V L��I:xx!H��/G��G�����p�*q��A��o@4#�x%}�?%������)�ᏇE=���3��F��%���ͳ$r�hӵ��0���K>z�������ӿű���ӧ�>����C�0~(c{#�>��	?�x:ݺ�0�u5��t(]�@���x��M�s�q��/S�Y|�>q$㍶�oβ�:�o<�μ�ͻ�LnI!�q�q��D0�Z��#o�z����ڶ�~z�q�FY��X�h��.��Us�8��?��`F�B�{'#Lk+`�x9y��uq��H��T��%W�@�c����ҹx����m�X2Ƥ�N�:�4�Ϝ#rN6��ަ���>[O��S�-(�Z�2۰س��c�J��o�����c����-�~�Lܖ�O�m��Y�u؞�~��n��Ϣ]��5��������Z�ak~a�>|�ο8�m��β�:�o<�μ�ͮ�95��.i���{������d����}9x^�rT��*�_u5V�e��>��ɦV�)�#�nI.Zb&+u�4���ͯ::h�#t|��l�&�,X�F�I�L��m*�u	���}�OϚܘZݭ�W��O�N�O�'n�']-��\v$�<�m=�
k��LbK4���Ę�1wV2�C
�Z�����1w.�nv]����n�Xi�-o�i>q�q��m��e�u��y�y�gN�9�HF+�$b�׸����\i��'L>v����g�'�z���>����4ц]nK��4�c��T\��>O@��z}NA���l`�_߿ ��$[cF����!�i�=�2x����$��;U����&̿v�?'�ܬԩ��Iqx|����m��S���g�ۉ������-���8Y({��^ >P|0t�1�I�o�i���|��4��8�m��β�:�o<�μ�͵����W�l��PZ�=n�l�9E�-��ٙ�]p���y|�Y�2хH���1z���E�n��K��$�=5�f#�^v�]֥%v��m��;EjhZ%x���̱*����m�²�*�T���dZ�aX��,h�H�ڕYQ�иl�un�QO~����?S�|��?{JRBx�@#�C;�F����F���0`�Q���A�l��L2��~i��m��a����^��Z1�0��6p�����"��+&�<�L����F_0���F�Zh��w�|@�������0\
o"B�4��F�ͬlkaJI]�1��9����'�դ���H�a�i��XZ�a�|���u�m��u�\q�[uמu�|��F1$���T�����e����1���Y]l�`�1!�%�g�n�JC����-�g�z�_=Wԙ]�$����:���|))���hKG��D�Iu㾷İګC�vjj\F��~��1[�r�˔����[��d�b�3]b�M�ֵ&[���߫�2��[�����+�6Ӭ0���#��8�N8�m��OS�$�I��9U��a��I'>�HE����T܉�)"�b�tt�F`�4~�M%�w���<��]:�z�닪�E'�^��\�Q#pĔM@\����9Hf\�M�,��풹��ߕ������1��x|w5؋���h��ϒn����e��b��>����5��Glv���9��O�?n]\�c_�UM��r�~5���[���:[̭���GϚy�\q��m�<N8�i'S����e�kx�1�4���mwX�a+V���2�֑��H��#�{?Hxx�>x�э	-b6,f�E��t�l�tNx}=:c��:_��O�4�bs�9��>�.�b}ww�U�8E��2�U���n�b�I���gr�o�#����ww�ߚ��-��e/�ļa�Z8㵛m�_zLW��ߛ��U��.�2m��il0�O[�/�i��]e�q�i�:뮲뮤��I'���m$ۏ���6�>aN2���'�$�O�x��i��i&�Ԟ��I$I��I6�O'�'�&�N8�a�L��l�M4�m��I$�"O^$�M4�	�I$�I$�6�q&�L��$�i&�u׎�˯u󮴓m�m�|�"$�I&�I��I<z�I��x��ĒORN&$�z�>|��L$��ǈ�4����)&�&XM2�z��$�M=e=I'�'N��>>�h�B}u�f�m���TBO�H�p�*~�gA#�Τ��b�86>��f���*>dOQ5[)l�v?Z3n�A15��/B����^Y��$"b�M��i� �*L�Y�W�%C��1��H�-�Z 
'EN�V�sQ�3Z�$�o;���k�i��$��%���.2� ��1��|h�S�s/S�R�R�ѕ��7��������רaR��O\��������%P�T���Ҳa$h���$��"9*�mF���J.~��BD(>l������\�+�IM���MJ�mv��gѦ��������ޮ��R�+) c[�4/���[�S*���i��(��Y���N�p���"�4�(C!E"j�`f�Y�e���2͛����M0UJ�ST�b�
������ޚ�o/��gh��/��ڷ	}��Q!\q�T[m?vDgH18��4��/\a���n��4���F>XVv�kd�M�~t��傘�S��V���j�����I�y>{o�����q�d��R�Lۓ`�K�2Ý.���݂貗��Qi�CMf����d�jc7������])�A��:���3�Jʹ�B��+�Գ@rZ��G]	��E��3m��n�(�Sg]T*؁���`��q��5HTh�j�*��Ct�f*k�7]X�.yeն\;KK�C��Vk��@��@��L��H��vf����SK��)pŅ�vM�*XKh�VDmm���5�6Aq��@���G������w�uUV���{�����{޻UV�s����w��z�U[��N��/e��ϝu�\q��m��8�M��:��?��;�%ܒ�c��3r�ڋkaj�ܚ��;���m	@��JB����-[f��%Z�ҹ�n�e-b�6ba�L���cR�6t#Zݕ�nbn#���ۣ��!������ꪍ�MD�t�L�aR��t�ZZf[s6�L^�W����.��[sZ���i 1���M6���d�EX�t����|�U麞K��sYͭ�E������@�6�<�-к����1�r�9)qV��CsI����G���t�􂬻��MW[�/n$��Q#5n|ܫH1�Q��=�&���(�E�|�B���߽�ˬ�O;w.���ki���6��0m��a�{3����[��{o��?5V�}�I��s��M1��{,K]{g&���X���PM15���v2i4�O����ԓst������n�Zt�CwFkU�r�m�V���L�|㮺�4�n���m$�u�^��g��f�I-�=_��N��9'�ť�#�c�']FJ����Kĵ�2��G蜒����}?J�V�}�VX���K�.b]�8��7_�>8��A�!����<,/�.�6��
B*�R��ͶvZ2�6e�Ɣ|/�|�6�?i~�G�fe�KE��\�n6e\r������r%8O�	[֋�'K�U
PLC����u�\q��m��8�M��O<��ө��ǧ~�HG����n?jf���,��a�A��s��N��X��-���`=��$��O�W[q�>p���b�`��b�^�v�1Q.6[��4���� ���$>sp�Q�D�>�����%��i��2�3M6���+㲛�D�u���k.|��ܜJmuF�`������0�\18�����Dg�b��+L�"�㌞|�n?�q��m��8�M��N�����I�S���S�in��\Z�bH�t�Wk�2u�L�r�}�4�o�)��{R����M%���l̦n��i\^m!����6�*���Ҟ�.^�/Rj����i����?2�髗W'�G����������+�_8��u&1����&F�1]�a9Q�w�&^�]�U�v����?�0Ry�臎��\Jmq�%y�����O1��a�e�zT�d�ao�d���~q��m��Xu�u�]u�^y��암Ē��f*c2� ���.6Qd��*&o	�d��됿G�,җ��)O�^�����Q,��
������E��$4�y"-��Qb(b6����m���qVl��ɸ�H0L}�z��M�ݛ��3c��Fi�(���UPK�{(�*hˆ�]��Z��Ě0�qe6&e���λCR�cv0l�%�՜y:�f�nnK�]k�q�s�����Z��/߭��m7�ar���^�]�,xm��sT���FY>m�������V:�8��H�<�~�x|wٻ�I-�z^�L�x��hч��4㻗.&�wT�3X~b�ކ��Z�V���&2p�j�$�9�"~��q�~'@Bj�'ɠ��I��	c��O��S�6�m��'I����]L��$�5�4���M�Ni�n/�^qŢW�����y��������ɏl�d��G��@�Kv���IR����1��S��I�cvd%��D��q���A�(`��{��L���ԓ��\��c!1)�f�X�Rj�D�O��Ǜm�Hq���h��}\J�ih�|̻�ka��|�J���i{n�cĞ���D}[d����M�yǝq��m�S�㉤�q:믱��/��1I ����{��$A�}�d�ųya�$��d6���[Y��qs�ۗ1���-�qn��01�F��7R�B�.H��2����5�j�n˼�;�|d�kq��c�8I���&/����ۃBN��9��=oY~Nz����q�$!�g���;y�8����b<�\�t��R�!@8����0�L�b�ﱷj*%INZH�|a��=��Bp��w
m�WIр@�s�Yy������ѵ�ո�'�?6�q��m�S�㉤�q:��~o�ޒI �!�~�,`���>�I2#N>�>�4����+����1��1r^��w��c��$.�׵]�)�%�䚎ec6O�;����ǆ8m�+l�NbO��a��1%��t�[,�c,��ޮ�Z7\��O�sw'NSn^ӌ�m̊�]�\kQ�%�FN>��X�/�&䍲m�뙓}H��˫�F\cG--ɯ۹�i�m�el4ɧͼ��㍴�o:�\q4�N']u��q�9�}��s��z�����'�m����!uk�{8n3���K�D�;S߉�|�}.�藵A���R6�}�-�@��Q�ݻXQ	-Knn��t�1&���`K�1�b�5�fũ�.�f������岾i��l�ЉqKi��"n�6cj8����3�8�\��1�t��Q6��|���L�-��_�qww������ˉ�团=Y��^}���G�l/��O9��W�|!�"���b�+�.\|i�]:��çSf�۬��2�q�QS��2l��c��|?r%�>?��b��.HI'6�W#i�4�ӈ#��b�[rW�oK#�e'�;đƛq�2�_2y�o8�6�M���q�Zu�]qמy��]��$���2�+���9\0��k	v�e��]לre�N0Gγ]�_$�w�쭜L剜�����3%���L!o�y����.���<�cl#N#"<��}L���b29�IM��v�g��vst�q�*�5��;��]?.��'�	&�#���?5ٵ��:�a�8[�9L]�k���'ߴ�W)ǋ΍�����~q�ռ�8�6�]u�^:�II����i6�mǈ�q��=m4�<N2���=D�I�oi��I��)<I'�$I��)6�(�Fē�i4�)$�$�l6�M&�IĒI&�I�O�I�IԒO�I$�6�4�Oq0�i$�L��O]u�]q�Si������	$�I'���|�z�I&�<x�$�ԒO�I�|�4��0�,"$�G��<D�O,&�Ğ���&�����䓋t��[SW+�K�ܕ��^7�/�c���t�O�3��I���{Y�@Y�߷�o�\�{�j���s���}�{������s�w��Ͼ�{����V�rt���:�N��q��m��q��I�u��$�i�~K��s��%���IY!�UȗճO�\욯�'ߓ�%W��z��i��3���u'��d��������G79dd���][^K�L��I���y����<���N>t�4�|Ǿ�]ԓO%ɇ��0�{��c�-���ե�^�JD�S���Z�tLy���@��{E�w�=�ؼbZN4�����?=[0F_�m���8��6�M���q�Zu�]u�^y�U�I"��=^I>��jS��r�9�]޾�j���O6� �g�9���$��W�8�0��mẒj�[KH�"��G�yC��!@�D����w�����S���8�e�OM�E�K���}.�<ۥ�˦Wꑭ�H�J�5����n��V�ޤ�Nr���I�[!��Ԛ|�_,�Ǐzq��N�m��L�u�]u�]u�Ʈ��\�q�3i*c>�\v����Ծ��F|�`T�J��ؤ�B���]�6�<,�b�>�vN�I��Q���K��׭�c.�ٔ�d�XuԈ�8����j[}�t<��S�KH�;�l͎��U��9VS���8��4�+��-���#�GBEƚ����Fb6ļ�;:�f�2矪�[u�~L�q��v��֛����F1xJ�>N:b��U�u�!�[�'��M��Ծ�	�c8I#����yu�Qg�W��ܜ̜q�vT�ԉ%0�����4h�A�o�����V1�ur��W߫'��٭S����'�(&&��9�@t$�b�[.n��aD�"9��I�����8�\I�%�yu���w�T�ٻ�e�ީ�m�-��8�N<�q��m��q��I$�u��bI��H�ܭ*V�]K�k�K�m�{I����?=7��H��U����]��D������ҷw58�ɇ߳'> ����:��P_c����^� ��7��%WA��O��`��ؔ�)N1���ϟ:�����%�.�LS�'\a2��[&.=&��Oц�M�RmY+!+v�V�,�\�Fj��յ�ͷSG̶k1��|��:�˒��h�y�����Ի��T^n��}���_���I����Fa�M����θ�m6�u�i�]u�]y�z�;��1U�� ������ ���I!s��ς|}�+u\�<�m�s)����"Ԧ<���o�\!0͍,��VU�V��c�-J��;�ݢm��ʵ���e�Ɨ�Ix��gM:�LW�6�m�3�f�ku��9�]�y_5W'Zy�mlq��R���V$��.�*ӎ+e��S.#N<z�����I��i��e8�i:뮺��1�jI"��vK\Ķ$��텯��p��3]zM]��bKkRJѯ>,��҅��L�����9¹]4&�M(�`�y��������<�Q{̠1@��4!�a	|�H��<�vMVϟ�\j8�嵌~���o��.V���4~e#��(�����r$F�4���Ku����<��.��ĘŤ�-���k�u0ʸ�4�K�]m�m��d��O:�6�M��N8�IĒu��?}���d�$���{!fW=A���d�"#���1-���D���T�TbŻL-4����=hJ_kafE�j�nm�y�~���'��z�WK�lIu�A��4ff�]IIt͕��&�����YQh��N0S(;�I�6� [���k(�,�2�,7Wmeq1H2��m�E�a��,%�8/N3�q)��xA:nw�?O���9;&�'�U�Ɯz�r�C���H�om��N7Vۇ(�9����	��m4e��u����.�kf��TJum��N�f"��R1P;�X?C~4`��Lx�и��@4��Q����Ѝr��3�u��+�$%`�g-�t��~=O�C�1�!�ޟ��f���2S���wiY"�0�����8�m:�a8�i'Iמ��3$��#M8|��M�w��?5��H��~���y������V��R]?s��r_�ֲ��N~Ě��������l9_��$��!���==;�8�����~S�0����^�L�-�aDq͹,i2������~Y���w]��-�f�$�w���|^`���7��K����H�i��_��0��S�ޟ�4��'m�\L'M$�I:���1���
� N�T1���4�Wτ��X�t!������|!���_��D:�d���R1�m�ڼq����O��KϜ/:�Qc#=ZVؼ���������bb�6��e\i��5$�4{rm�i�I��<�d�4�u��w2�9Da�5Q%y�^1Y<�imSf��_WֶY�#��]r��-V�h���׍=8�O䓍�Ӯ&�&�q$�u}���1����}�}��~i�e�H�$�>[��/�%e�~���?�wKf�L.��03qD�1�l�^3rT�n%[�x|u�ս%��`�&���<NB�8 С`wE�a$�e��m���ZI\w�����o� �i=�~1C��zNW?`ڸ�u��q�]ۭ~�:ӭVѾ�Ê����{>&�[��e4���U�Uٳ6q�7��_��ў��u���?���q��31�eJ���)���s��QY���Q���m#x;s3���!�E��"ȑ"G��-��"-$DYm�DH�dH�""�m"D��!4H�-��h�"�"D[k"D�",�%��"�"D��m�""D���Z$H��!"�!�fq	�Ah�-��"�"D���$H�h�""[k"D�����H�"$H�h�"[i�""�"DE�D��$DY$H��Ym�H�h�"D���,�"$H�H��"D�"D�-�ř�H�h�"DD�։",��H�h��"E�[i,�"D�ؑh�""B[e�D�"DдDKm4Y&�D���"$Z&�"",��$M��$Z�H�"�$[D�,�,�"D���"D��m��"$H�H�ċDB"E��-�E�D�$Y	m�i-D��mm$Ii$��4�DZH��k"D�If�h�$��If�K!%���c��KI"I%��$�$�E��$�����%��$E�ċMkbMd��Zi$ZRXZh�,$։$Z�Mi$����:&�I,-�,-4M%���Z%�,-kIfZ5����e��E��k4�h:[��+2K&�k	$��-lI%�V�d���I�a!i�K5��"XZ$��Zk&r��I"�Z$�%�H��Z$�E�,�Ih�H���I��$�m�$�Ii,-4�,��$։%��5���h�"�ܶ8�ɤֳY"-4H�Y4H�Z"E�KDI$��5�E��4Z�I$K&�%�$��h�Y�Zi$�[i$��$�mdD�E�I'^�gM�H�Y�Y�����l���e��l�kd5���{���t[H�,t�:�f����l��de�e��l�X��;�:�tm�[4#h[m	���BƄ4!�6X�����Bf��	��	�����m�Bf��Bd,B2�&���mʹ-��!a6��l��M�d�	�XжhM���lB�-���d�!�m�cB؅�d-�б�ɚІ��B�#B�B2�6Xг&�&�ɡ��&��,�Y��4��e��g̚ƚؚl�ƚm����&���3�KFF�[L�L�L�Y�[d�FM5�5�5�4d��5�4d�d�dd4��44��L�M�Y�M�[M��&�Mh�M5�M��Mf��Ma4�Mm�Ѵ�4�m5�44�m4	�Mf�[d�4Ѵ�4��[mfM5��m5�h�M��5�i��	�i����f��M2ki�Mm�8�Mm���	��	�Mbi����kFMlM6Mm�A4�4�s�:J^gdn�X�FM4�4�4��d�d�4d4��X�M�FM4d�X��2hɭ�kl�i���&��h�i�2̚l�̚٦�&��٦�&���h�i�ɦɣi�i��hi�&�ͳ�a5�Mm�F�[CMcMl�[LіF�FMa5��i��Y5��FX��i�[&�MbkM��M2�Mf��4i��LMm���A5�ɓY5���ɬ&���MfM1c��(�-���km4ɦ�Y��h�Bi��&�M�p�F�g9�b#ZbL֍#H�M��mh��b@�4���M�LDŐk!&kBD�dgn�n�5��I��4����!hDH�M��$I�Б!hH�BD�D�$H�$HKbА��4��BD�kf�hHֱ�s[$Z[D�!kl�$H�Q4H�kb"!h�!�Ȉ�!��Bh��h�"B�E������lZ4�h��m!d$H���ӧN�s8D����h�e��"D�D�$MlH�"�"D�[i$,����$H�dHDH�ؑ"E�""E����-m��"ȑ"D�D��x�d$H�m%�"�"D��"X�m�E��"E�"D��,�-�D�m�Z$H�"ȑ"[D��,�-$$Z$E�"�"BE�D���B�i���"[iBD���HY$HY���o��+�F��W�����㹛���g�?��ٶ��%�1��f�T��OM�������^��������ݟY����������8�����{�������vI��=.���GMπ�y��]���k����4��|�?���O�����a��p֪��K��o�鳱�o_���ݷ�����l͇���_��?~���������-� �zv�^Cfl?�mȄ�[��W�f�����O[�Ǵ]��Yg<�m������m�=���o�֝��>�g˽����G�7������D���·�t�to����g��nƿ�z��n�t�|s���җK��i�����*���m�4�>��׎��}��vγ��)&��������_S��w�A���g.�c�U���M�nfq��ٵ�ct�nhٵfb���3c�l�c�kcn��}�p�p�Ǔ�	��st:�/��vu7;7��;��z��y7��3n��!&��$a��-1��Lͳ��1�(H0(H�]�����o��i�Y���|�f�~9�o���|��m㼇���é��?��;>���/��.����#l͇3�n�t{��}N��3���w|?;�o��nǤN�:�ǳ� ������w��:���[�e��D�����>����~^�����6f�ُ��#^����?Q�s�����C��z���E��l�ogn6�f�Nϐٛ�{��3-������%�Ӧ��}G�����W�U�a�M�
[X}���`�l����Խ-�W7��i�,�x��sb4tgp��M��۰�Gsx[�\�5��9�6���7;�<��w7�&�:GWC>���:&xi]����x6ٛlw��%^;�zp_7]�opٛ����f�	���=��m�y���������>C���{s����&t�?�=Μ/�}'���o��������mϖt����}��m����vl͇�0�fz��p�o���q�6���>g�{���o�=���y��[��&ξF��_�]Y�����YWo�����ik�7�ד&�q�#�Վ��������dt:�_ӿ)�����)�a�YV;��hU3a7�{y����\�rφz�����8���mo>��o}���3ӛ��ɏ�S���Sv���V�~�<�^Y�-� ��[>��(�=��xpg��������y<�v��q�㇉�~O��w><���7��;z!�~率啧ۜ87L�x��������w$S�	��I