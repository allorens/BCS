BZh91AY&SY)p%��a_�`q���"� ����bG>�     /�L��TZ�6bR�*�m���ZŭKm�IP��TkU� #e�4R-��dmX+,�l�Z4��֔*�m���mK-W�묵j�&H���Rf�ՉY���F��[��ET�V����jkAdj���4�-��j�����U�Vڔl���[VZ��Q�5Ul�f�nr�h6���Qm�ВA9�8�mfJ��&�U,��v�m���m�U�f���ʶ�,�3 �mM+m�ml4َͫlAET ���	m��+8   v]>�V����ۻ�[��u@�)�zYM��vm������/U@S[Z���
ʁR�f�Q[P=�����	h=��ֆղ5���Z�km"f͔�    {�h��ݴ���¤���q�s�W���8=��T=瓎P'M�^�z��Rt��{aT�w*UR�M��x��^�Sa�ѷ-������yR�צ�E���V���|   Y�ڥ"{e۳�{�U*U^������J��N+�vލT�D�T�]�� �[jR���z�K���}���
�{�*����|�T��U�{Ԯ�Bj�}țV�	V�5�aT�  �3�J�UK�{�_=�=>�T������/�'����{�JB�Q����zWMJT���_;����U�Wϟ>��YM���yAJ�R���I(J����^�G>��T�,ڊi��
+m�L�  �w>���N�g���{/a�Wޗ�<}+�W��:n��T�T����ޔ��Ig���*R�'��|��'�*J}ϥ��
&��w>��ϟA�J��w�Wov��_l�y)/,T�c5�Z���ʨ־  ݛϢ�5J��w��}%���IU���o��JT�}�O�k�ZU)J����Mg���׭�-�T�ۤ��ޛy�H�*g�8�T�ҭ��:�����=]�]�����*��f��* liH�3�  �w�Ҥ����P��Sޞ]M�J�R=׳޽�ݕ*����%J�z�{��zP�*���{����涠�b�h]��{�鶪�Z�٭��F��c�  ��\��ꊪ���W� ��=�5=N��^������{�@�lm��ǠMw�����{g�� ���ٵ-��d�@�)6X�>   }�}��h���PE�S��
��΍V���{�@G�G\�^���D;�Ǫz49޳�ֺ݄��Ļj��)Mʊ6�k�����  �� {��P��V���*�we���4Uo/^��:���:PV�%��.��4��n=4��t�]Q��     � ʕ* �    Oi���(      ��d%*��4�@   �%J� �    ��&
�(2 h    ����	�Sz��Hy@��d�O��?8�P���������>�����]�V,ϖ�^ǟW�{�=������=��_�T?r( ��UQ_�8	������x�� TV��?�⊪+������������w��/�|G�e��&�L� �)���W�/Y��az���� u�� u��u��:�ez�ez�a�Y��� �u�:�=dN�q�:����@� u��+�W��Y�=`�X^�=ez��������N��u�:�����W�/X���E� u�:����+�G�'Y��/Y^�=az�ez�d�Y��`��dz���:�L'YC�	��u�:�ez�����C�u�̧X��dz�ez�d��d�d�u�8�e�'X��@:��C��YC�u� �EN�'Y	����DG���YEN��=a:ªu�T�(	� �(�XN���aE:Ȉu��"	�C� 'YN�(=`��u�P� ��C���YQ�*dA:ʂu�P� �����YE�eD:� ���
!�C�'X N�"d:�"u��(	�T��'XPxȡ�PC2�`:Ȁu� �*/Yzʣ�Q������`P:u�W���eQ�"�Y &�d@:�+�@����Y�=`z����+�G�Y�)2=ez����#�W��Y����� ����:�`2�d��Y���@�(u�:�a��Y^=r������X�/Y^��`z�u��)�S�'XN���������������3���Z�#��Q7ůW�I^�M+K3�ۂ���LB�:3 +�<{����d5�j�6$�X�&P�g/s-��;��c��ԈI����;9o3y�
r�"�X���"*�k#Uy-�,ZبG�����YÄ
me����a���*���:�՗���K�аł�8Ù���yw����퇪�鎎S�c@#N��c]L.�z�/6�^�NP���`"�1��͢�f�Ѽi�K]f�Q�O/}ƕb�gv�t���5�Ե���wn���=)�)�K9���_�R�jͳZ��ӨT�Oa͖ʳt�ct��af�Ӡ��X�Xh�.�]^ۏ^�����Z  �x`���ٲ�����)7�7�]bL���t)��F����)R��6�]�Ca5K�y�ܚ�ތX�}(�n'����$�Y�Crb�է�3n�v�3>,��4�e�te HѠ'Q����9�*��5�٤S�e̬ٹou­mj_J)ԓto76ں�$&���v�W!(e�Ѡdf$��X�I��.���Ik^kR]F���I�]nHX�N��6��%{=!!-ė>=��D�x��<�}\��t�L�&������HѴ�j�Oi����<���/f*�@l��/"*U��^)��:MKU~֖�,�J=�K��s#�ܡ���y���CrT��i��+[��m�rl�2�%fDkMw�.K�$��	-��ֻ٘U���2D&S�K�4I�k�ر<���cp�>:u��Ymb\Q���wZ��<̹��%:�mH�$h]00����!��ݭc�6��lMf���Il j�(���ʈ��(��m��̔㬖LM���2�ҳ�h��6��v�ܑ�L�l��ZA��,��e��b��f��cp)����z-ҭ��u�$f�J�GYPȫBKE��dK��%�y���	��b=rҬ&���``����zU��Z�Af���c�C����0��nlU�pb�F�4U2C�Mi�Lkf�y�P������$1����ůwV�Hش�q�iU�=\��u��9}dS]|���)�&�i�fXF�˄)nLb���L�P�ËqC� ��݋Ҳ��ƈ-\{f��s%l&�=X�X��hh�'�|�6����$oq�d�/i���mm�-�o@llRX�o�m�N�!h7y�Z ]L[�7f7��į-D��u���1�6K�2E�sD�Yj�+#�q�C�MgN�y�բ���3g��v�)U(��Ei�����b�)�:ٶƸ�m�@="���-
l��OƤ6(L���A�=�ye��������(�-��.Z�%e]'� FZW������jGoV�Z3a���$�G�NT�(�	�wrnG���L�
��*5�P�����9ۛ���H���^ra�ڶ����[�����	�!���mj�x�0� �1�B�J��z75y8-��	^dg+JŏC6�X˭��A�јo�R$�s@�&5*Iw"�v@�'�NS
��S*���l���dl�t㯱=�Vs*�.�뽤YA����ii���Pwb�YfQS`11f�.�^`�aY�-�C���&u%r�
I���"|[�/#��0 �қ���������왐;j����a��Q�����7T��H;U�k���-S7-�fk5}��w(эb�YHMc%[n�$XrL�j���W��݈wn��`�����6�Aj���I����?X4��j�����Q%��CD���Zѓj��R�ATG4��ܖgۻ#P=t�V3��ݟAX�$�w+&lgd<�G1�+@��,ڣY��Pdln�M��6T�}���Eze���\�/V���q$qmi������Qu0"dݺ�m�ti�bd��̊V�*�z!�S�R.��Y:>A6	�ч e,�9�U�Vq�vw]�D4�0%3�륆�[�/��JZ]\%Z��Q맇�twr=�,���c�Y�6d��x�+�Řwf(�6����u������ �k:P�V3U�#�P�SBZ���Fh�� ��gv���v�*��&N��[	Ѷ&e��F<�3%�����`"c�Z�X�)ed��A��Pgٚ�h�0ڻ�/��I���gj=���+�p]���(��*L�Fͦ`i�V�f�헌AQ�zVGDh�ja���[1:��m���7�t���j���a���7o�\U4awW����B��*����J��x(����m��pi��t,���RyBK�)�A'I�O�1�M�1@-a�JiJ��٭�an��d�87J�e��E��2m�њ�<ӑ��f";Lb����y.�SU�m�rL��p�v����X�[6[����m���M(0!2�LMQSn��)����P�U,V�x[�T���hyՋ�\�,:� ���� ���1桛[��{%��Vv�H[eӸ6UK�d$U��.�C���;�Qㅹa�� �
�����6]\ՙ6G4�J�9���5�R�(�JX��b�r���f�����	ݘaƕѱOH�V�a31�I���i��qaҋR��m��35�x�|i���De��(3U�8*�h�,��y���wJJǻIV�T�b�k�U���v8\����ӵ���U`
}�c"&��/�-mG2�U��I�v��62e�QX��ʤ��T�b׬fU�t��4wv�ݒL.íWG.����QH�AG����uy� ���Ʋ���J�Ś��$�.L��AJ��F�ؼN��Ҳ�FZz�;B���nʄ��	��N�F���Wh��E1UO	�c��B�Gzs"/Qܬ��f�2��X��j3u�@�9r�R�P�j[�̀�$�e�wq'V�m+G2��N\t�ɗ 9�UH�ɤ�ƌ�P���u��Yq�K�M��)�dLU+q�:�;{2�A��2���F� 2�m�1P0�;�kF���&5����Y�¥�3�M�z-F��B��w'�z2�=9y�����i�N�����\l�1`[���B��%�U1L�ʘn�S��/r2
���"���v��5��lS�%��x�Y%�1'�e��*���b�$.�B%[���&�v��sq��K�o0;�FF�	\�nZ�̡x�-ia��^�Z����n��ZeX��`]X:���+f	���u�2���3m���T��v�=b+n�����L�[}]��'��.��2d��);Vq�7�]!�V�Up�JZO|m�̊���K7�����3c����	�+�J�AM��9�
�L�+V��;X�ڨ��*�5M�ub
f���f$mY�y6�����Җ1�VIY4�6�8̌ތ�*"蓘ڻF���f㊝c�opl"֧��Q�vU�o`Ԗ��XR��Sjc-���uB��54#�.�Ӕ����i�e�j�V���VAON���!;B�<5.��Q��C),i�kD8ͣ��z�E��l� ����ZE&l��Q��6�f�eE�QM��l;�
ذQ�)����X�@6��uՈ/H���ˎj
��V�k@ �ԇ6	b�lv^e�z��1���'�M���V�<�FEsq�����#A{p]���$z�+-�X�<�B��O~�FV/�q6�T�twI�Q#�>�&n���ӆ��ʺ���{����)Ɏ��I;	�p��>f����Y6�*�������B I�K[��$�)�f�˩qe6/pK�*�j0�i�(�:�tl-�)�m-�,��\ݶG���
�1:�a#���a!6���ܭWq50Kn(rD�f�1=1ScA�3�RvQ��B�-fiT�G�j!�L�Y1k��9����uh"+s�f���]B��ͅX�˳R9��M�w�,��Y��ِ7=�ɲk#U4������0��t��ŷ��{K¬�V��U�Y
ߖ){(�`��M�»b"tA�����Q7EP��bb��G�^E��xV��h�����%
�Ϋ�nn��Nn�`�)a<���mѴE���t��:.��ê+f(�l���W+5Қv�aݖV\�z`x����u��VZ�)u��<Xz�d�V�a#�#C]Й6��cӷp@���՗72h)o��	��N�ȲK�#-�vHU��9�@��t�QT�hy����ikuâm&k�
��m��[�����C1���e����f͆i�4\�$�˄-��6�\�j2J�Y��;D�"H^��Mn2���mB����^eQۥ�D����D!z�܃iPV���a0��	Lj��E<WInd��,���L�7wE�������JYAvi'�-7wJ��l
Vy���uyđ��@�൛��c�]v�uS��[�Z�1	2�X!b���ʔwn�J��qUߢ�9������&P�fT�fR�n	�1���T�Y�Хw�k���ek��s*�+����� u������b���q;��KZZ�3i2S�e*5�<kb��h�d�*��1Yh����� �w�DCy�Y�RB�*���,�Z��셕	׊-w��ĻV��6- w��w۫AX9f,�̩A ��XF50䀩�i�k�>�В�NM7��[�oR�yl�un��1J���xe�l�u3i*�Mc�����Tœ�X��:3(0`:��p�Y@�)�c������[ٯn^šd��1u"u�v���{@�@KUd����)e���f��X�!�ٻH�m��7f�n�؀���.��5mm]��k=�J�E�,u��a,�[�<}���ٳOIky��;-lu/oU+�NaG�B�$�Pa����s:{Ed���ItLހN,~u�;sJ���l�+k\Es�$D�%��k݃�v"�Z(��0�"	na��T�ѽ'BXhя(%K&�)�����V*������J�u%l߲=i���Se-�ø[0�����3�͔H�{�c#{GVk�.�O.��T�x�ǭ4�u�}ָ��y*c�lՊ/�>`��e�	�U����[*3�������[Ԩ��7n7�����_�q�.T�kы2�X�J�$U�w��@�Cn�GR��)��5���L]�������8���L�/tۨbt\hw$aڙ!R��8�,ZƩRJ��� L��Քǆ5��� M�6MT,f�ra�e�$M(�M�-�F����ͫ�`E�̬u9��eE���Qޢ�4�=y`ޑ�|�k���6�@m�ݔ⡰�ݭ��k:����X̛��BixE�h�T���r�<���V�{�0���[�4�W�v	�6�N�4-�eB������R-ٸ4�V� Sh����spa�d���4k�$����㧦av��
J�mnV�ը�+),{f�&-��)�y[3&�Y��t0��&iV�IL�2�f�+�:���ݱ-�= 3`0����JZ���T�뭣Wo4����l/Ǖ��W�)^�n�Hî,������P��Y�T�ã��0�3�u�� �tiM5��d���\�V�C.C�4q�ZaS������B��I����Ys6�6����X]2�X�q���h��
�8A�I-��hPz�n�ݷ�"��L�!2�n���K֪�b�V3K3V��lZ��A�k˸�k!��tFm�d�2��y�Kp�W�r�����C�D����HJ̙��[8��^�S�E��`i�,��@�I���&��%�HPAI�kkZ���<�GA�v����f��L4�������2�J� `�K �%��X7�m�;[X,c
�-|�"�=������e�4�].gw1��R��",d"��T+j*̷b5����/i<�Q���i�p��4e�4Z���`�R�˶\A혫i���3��سC���"ە�A���؆R��k36�P��Rbڋ! �]L�p�T��ֺKd���Z���̋
e-jRn\���:�so1L�H�Ű;����U��X-6� �N�n� �a�$�V��Ti��#y�%�:n����TWm�0���M�7aW(K�N[!��Z���6���dl&i�si��@?^�t�����p�S#Q�ņV(]%�� ��j��րj�dײ�ThS���)�f�b[YX7�+�U쀫j�Hjhtn@�n�5�������o���okN��U�j�f�X-J�^q�Uȴ�h��;9���L^^����J��Վ�	�a�n���/r����E��[��U{V�C:�搑sh{���CE�.�,�쫒��F���-�0Zˋ�P�Y��n2��b�����t-�6*ʾ�0 �iIC�(���N+���
��v�.�#�j���Eբ�RP�=��ӣj�Ż�f��ܭ�E%c՚ѭ7��e�V��������4����aХf�R�b^��:�'��;hڗ5e)�٘��O7��� d�o�<�H/�tb=}��}��VQ�v�޳�['-%�^O ���m�����a�(ād
��$�2�ͻƱ�ˊ�E��-��Z�E�����x�&2�L��z�vp�j�:��@T���M���l�w;"�ҳ(�eEB��R��*(�n;}(�E)�Bā����[�{��(dǓ���wj�y5�3Xu�I/#h�Y�;02����A,�(YC�z���ܝ9���}u�&*�.��A��0�:��^��j�+�p��"�J���#ꅻ;��)j1�� .���`�;���y�q��vE��mW�T9i΂d��>����~�kN�㭉gW���*�Z]�LCb���9M-r�y�z�EuŘ�����ev|�Nkۿ}��<�G����@<pZ溰3�#�3��X���}>]�;�����	�L���΃Dm�ɤW̓Az-�	\����[A��NOY�Y$�$����>*ϑu�u�'�#!�z?�~=�6�m����_z��������W�d����!w�'�9&���k{5������:�(�U�ە�*k��>7���e��=�U�(�{��[ٟ.�-�#G�{U[��:�(��Ć�c�CF'������)�)��P�bRb=PvŎN��2�9�ŬW�,����R�d�����7f�9!�d0�=۸�����,�v��3����h�����n��Zt��Ń� R�o(Ӯ�|��)�|��T�� �qJں*e��u�k���}�m*�2f�ܽ��x�j̬T.��ݖ9�^��ͩz��Z�$��xY�[�+t��9[�!N����hn 7�S�[���1�8��i���n��6�� ���4H[���"ܵK�5��ؒN�%φT�.̱z_Y���Q+�2� qjئ�{.n�N�tN�Jm���:�,m�o[�B�&<�ΎWZ�v���<����2� �"ќy��m�}}X�0���΄� U��j�"�(�a�!i�YW��K��,K�[[�]λ89n�D�����'m�ܙ9W]��6ԙh����8c��!i�w{sP�y9���+6j�{U7%�G�Tx��=;��{�̥�EB���SǄ?��\R�H�xV+B��̂�)Y�5�;9�:̾��U�Z�_�:)�"���Ӧ�.�T��Gw�FiW}����[�P��%�ar�s)栱in:/�Q�:vȡL���*�V���ܚ9f�Qa$y�4��#����oEÔ����k#��33L�*V%e�*M�$�K�Q���w�ݚ+���K�U^�"���\���Kѭ���kQ���]Z�#�|���������W�=}��ǁ���ȬU��dݗXZ�*�X�\h �����%�Ʌ�T�osQ͢��<sz.E��IB"���̔�v$�^�gl�6+C>ɽ��S�i�%>�S�%wYJ�d�ͨQ(�s05�����_ۀ�'�$�B�O��%�K>��0(%�##W��5c�ao6t6�vq�{*e[��y�U1
lt\����p���^v�|�񉵬���ِm�O��'j�96bU$׷[��cz���_WaҪ"0f�;+�C����n^P8�,K��O�\�6-;+s	�.N7xL����hu�L�-,�f��T"Bɱ��C99��'��<�sJ�:vF��K�}����5�y�5�qv)		�D,���o��	ձ�u.�5��0��R��b��uS'�>]�h��T��a��M�{CHx��,NO��`��c�ǋ�O��=���(_,�˨��<���� x���\%Ƴ�bIا����ҥ��a��u�h��jN6��,��ۯ$�jWK(�t)�r[�X�ĎkY[J.�Ie���c����pmvi2A:?��^IWZE`��`��2͡�s��M��NW$޻��� ��0�5�2p鲚WL!`����xm
�gq#	��l�����V'�4R|[nK���YG���wF�۹%^��L[�2���u�ҧn �9��!�ʀ��Y�P�S̹Y�/i^ڦ��k3)�(̗�:����d�q�b�V+	tֹ�����\�g�1e���r�M�m��b�?e��o���9������'���r���%>]rUs�9̳��Ȕ�Վ�R��4�N�Q�e���]�p܉X,h���z����JWc�t��(��\�ls��J�I�U<�9}�G��rf����;�n��[WM?�]Nf�F�ݗ|��`�+�y#C|��Ff��;9���J��T�mǟ||�dE��V��}v��i�S>�}�N�J#�A�.%1�t�r��o�턵�Q<�w%�d�y�IW�e�w�)e
±d��n�h2��ң�gTQ��h@�Po�I�Qd������+)��]7s�T�X-,��3�|�Hu�rƇ�Сk��Qb�g&�Y˖ȫ��|��������ľ�!�a�#���8>��������(5F���@���d�O��� ޝ֏5j��s
��2s�'˽./�<�Y6��3�m���gKc+NXT����csD��J�Z��9gm,i�F�9���˝���t�+��=?ژ%������'�`z�c=�{�p�
"�M)�������Y	�
��55��]EG�MiT��5fh3oL�Տ�8h�ɚ+�T��FhG����}�����V	Z-93W:gu��o�`ɺ���;�Ξ.\ht�Υ�SX�ιӎ��.��$�4SűfݗBЧS�^&����ّn� g�
x�3es�Rx����⭇��h,�V$���YqW�������udӼvg-�\�M���V�к��b�Y�fت��)�Ǣn*,��Ç{�a��[#�6%c�X#���s���EcStLYѧR������Xa}V�oG�4��ej�WWMʥ'A\x"��uet�X�DI%�VuA�:ѡY"��E��d��0Y,�����V��⦶�˯ül�^
�r]�]��v���.����	�^Y�E:�}ʝڔg\ۺ�-��[:��W@�M<tf]�[JJ���	s�;]��`�qi˔s��%���(E>�u���E����Bۑ�V��L��S,>�S�5��"��{��ӖgW[�$� ΂��L�6t�P.�Yp�:f���S�K���ȷ��)sF�������l��u����{��\њN�\���r�e	*9p̌VU���T�_ܘ�gm�ˤƱ���M�F3O !��Ѽ�m��T��m����e����jP�9uZ��:6L�S|-u��"�ǃ�J�#zhL@�9�s�S�f���Xk4�x�fQK��J��k~��H��l��]�IS� ��xp*/��Bm\Fdra��Ԇ5i��\4ߔS�kΛ+@����	ݾؑσ���{&=���l�/^ި�-� �(�Dz�_����}%y��f�M�����h����u��>q�}�fse�Y�+��6��D�{Xsj�Rx0���,����eMi݀s56��Y��"x�
s{QBJ̭/q�CK(@`��oj�g0��ɖ����b�s)<�شY�K�)�e���:!��%�x�3d�X0��/� �]얱J�\�e:�)�-KB̝�y�.ﮅ�U�.]Hi;�/X5�h5@�4ܗ��p�LNT�B���rf�z���*���o5�p���o���A��侚A+>�t��C��㚫��P������Fz�w�7tY�KqA�����fkȊ���L^��:���"��V�ǀ�|ݱV�4�2Δ7	��f.�)�N 7Ì7��h񽻰z��+`8�!��>�t(�M&ݲ�K����;����NF�H:��O�v�zOr�C����Ko�'eDɚ���{/�$�2B/�J����v&�vk�W]��*G"�2Y.�,_(6�6"�)����p��ۺ�N�b��N�Ϟ�q�)��e�Tk{}-���YBD%�rs�p�rY��F�騯;�#�\[8�����;���h��ܯ���U�K�eh˸z��̤y�0(u{w9��K�<�k^ي���g�ݻ���eV�!�A3���p�T����0_V*%�%�^�{H�,��R
�J1L�75��<���՗{����*SD�L�xm���Jl<C2��bi���[��
��e'l4TdU�������%��I��`�JT�
]��&�܊��f3W�㮧�m*٥�����L��8��&���������;���Pn���ue�[7��R�U�x����O7���P�ߧW3�G����ip�����	��p�J���]�f�*�I��)E��K�<���E���,�.�[�'-f[��iq,@k�JC3��M]���ܖ�.�&7�U��}+��^9��)��
H�9��u<�qP��]6�E��������0%>Ҝ�X�����o������+�b��ab�T{���b�3.�EQ�����(m)��&,��2��U*011��Y���=0��u�yʻ�i��~<�Ã�M�t�*�Q�G't�Q�t�;&�'f��Ʉo��� �y���V�q��N�'{i_ ��L�B��jާ�i�ɥtro=�0ٺ��u������vd��녽�]�� 5Cҹ�X�f s�!�H'��rMȕ�J������U��s��m� �)���������Ǯ����%�ǆQ5;�nnu=9��7W*�k_Z����%�x'Ii���Ʃ6i�����Ԝ�SܧZ:�p)�YCQ��
��Q�Қ+	�%��b"i�
�Q<؍��Ƒ\���=��:���Y6���QTP�O%��'gw�_0rc�]t7N����AO $��
���B�J��2bl?����3[��SKu����UG�@F`ϴ��bcB�sU��	��j3QE��~w���{�
p�����+�\+y�΄�hȐ��ҕ���Q_V�m�����;�b��m2�4n����VY �/6�(��8���Eӛ�b�;��]f���F�j1���k�R�8�܅9w�vΘښD}���}�j'�^.V.�:]�U�oWH��&ܱ6���~��c��tc(cu��wm����`	�I�
�';ݭ�6S�΅x��f����pW<�%hj�RU��Ȫj�ˎM��YW,�W�:��L}�ob��\�Q�q���Z��mn�,m��8���ҧSB�󭹎�[�;q�fɹ:����\�����iΝ0����ҟu�k,��:�[�\.�X��c����+�6�j�*|�'xI�Y��R��և�����땭-�
����^��9�����☢=�_��c��'�v����;�m��r8�X퓃���p� ���*�gn2�gW
&��lt{N9͜��w���IKzS�[%\��q[�:�z�9Y��挤��h�������';a�x+��sWJ��h������*��RP�O�����y��L&��$�n�B��0[W�
�K;[�H�:�.��[�uhj�p]]{5���*��aS�nӌ�����H 핐N��gw{lju�����bӅ9�cU!��n�:�m�k��<5�"�5w�ZE�X��ʗ2ZC�i�S��R�F7��x����37d�un:%��
=n\	�3�-S�s�4�a��e�{�_INʫ�:����Ҩ�rl��mhTp��(���V}��·y�pC:���c;h��ʇ_N]�*u>�־W�@�N1^ou"p��V^m=\Qyr��PCO���#�H�
w�W|�]��y{Enž�NcI焸��/]ile��t&&>��9++�a�-^��@�Z���*A|�+��"�hڛ�0y��Sn.�G��L�V�ЮZ12�i8��%fV�\ɼ_>��)G$�CM�Q»������5�p��FJ1t��r*U��`��Q�a��m�]���)-Û�����F2���
͉��m3�Mut��+fr�sMnVS�]< �Vj����ddB�=�o����)��]Ȟ�EcC+,ul��.�ݼ��$������7"�MR&�U�q�4�%�

.�̆�5�Z�([��wz�U�)�j��r�2��Ω]�Kj�ə.CzàwX���+�2V�_n�w(����癎tۺ�9a����V�w�	��#"x;�oq�1�6�yn���hыDe���7Ք�]��ݿ�8&�	���9g%^c
0�S�!M9��	�+\�M�f���J7�T�`[k�x������4W+�2;���D9.�@�NÇs`�I�l��(w�)�L@�;�g�/aD���(���2+w�3L2��t�bW���4Q�
�p^_Z�@Ju���B2mHL��,�so;*�>=�Ւ�����Z��KR+��������ҍe�[��+�M����!�(OlCi�3S�F�1ŠU���ܥCQz�5��/q���ۜU�"9q�t7{#Ә�^��N��}'0�Lyd�:�L�ڲ�VZp��,'��_RII��;m������3@A��9��) jEވ��d�9�<'���b].���ŵ��n�ĳ�ޱ,<�묌;�jZ�N��0��śђ�X|�d˄	��j3��Dq�y:=�EۡWZ���� '�ʁ�g1j\W ��
�=ZYs3� Y;	"��&�J81:�8c9{��ٙ�U���0I#2t�F��yAd��ա���bU���0��[{�ږE�%�*��[�O�˫�e޳�.�Ks�L�/`�/�-��������4
9z�v��3����}0�*7�wKL���m���e���Ed׵����7j�Ik`��wc�_w�D�e:Ŭ�M�8.۵[�H,�/7Ev3��1*�������/(T<�5��W��kD�=��O=�P���<h}o�/!�.¸���Wd���{�]��y��jc,�FOB`�c�v���mn�����B�&�3�6��"���X\ǬWG.�ʹ�Vz�aTɒ�|v��]m��V�����j�me��X�$�ڷ���f�j�3cVlX�mH�:{��/������2[��#u�I�޷$`aRIް'wwQȚ�N���?+n�Kl�t\H��SCﾐ�tA�b2�s��n!� ���Ӧ�:@ݻhMوQ?6)y�ܡ�0ǎ�I�qѮ,S��/��g�C�P��B��l�(R �����G��gr*���)�r%��HD",�k�\�m T��4K�W�X0���-��5&*O
t�/����p����VU
EU�%`'A�5�9!�mb͵N��F��O<1VTD��j���>�{����*��������(��}��g����)��ꨈ������_�����ן7��F�o�@[��ES_�n8�e�/�|;*�B��B��z�N�E���h�/{
N9���W�Է�����ӓ�����)KL����]5�7�k�,��Y*�����ب�ފ��4�%|�gJ�9��gm����_#+n�A˭�"�`!՘��+WT�E!��K�*�^����xl9�5���ulZ��H��,b�Hؕ�l�F)��e�Lm9�>�����8P���]�/��$jr���]&Щ�Nd���2��F5��m��FW;Vy�T�����Ύ�R1���n$�=�p�q+7;M�փ�/H��w�6M)fۥN�t�����-���ө��g�i�� ��j�v�o�h��
���m��t��Jσh�˕d�S�q�$|�̒+� �����gn\��o`jΌ'L�N�p�	��!��]�nv[Q2�t�]���A-�'�y��yѱ��8�+'m#��(��]��p�ŽX4�9�iˋ_f�T�A*g^�
�A����FCN��i�4LL�sCM�eM7P�����)���B�X��D����e%� ���Vj����%h��}R�s����;2�\kV����e��̏�s9W�Rf�Ӫ;��	���1� ����u�63�4h�\L�������b}h�A����*��Õ��à�#W{�TUG\�G�j,9o(�ۂ��`��P[�_G���|}}x������������������>�����z�������׏������}>�O�����}>O����}>�/���7jmL	'�Ad�v�t;�:\�H��:��K��I��7+�%�J����@ա�3��&;':J�(.�[�12띌R9\�ȵ.�����|�Q{Y*V��O{o��R��	�O�^�S���wS�M�|�bU^*5Y�S���=�1��rv���ݕs&P���n{���#����ѓ��T���|.t�5�����t��b[��cj�p��a���27S��̞�P����w�1��_k�i�=I`f̗���Y�EZ;��|i�H獸P���(\{�T�5�q��e�8t�ї���;;�e�pΰ"�eUNy�Љ�(�Ӊ���=
k�i7\�ga5�6��ol��9CD�T�!��O��g�L":O�ܡZ���Ƴ*�T�c3kjMPj��FD��<����G�ʂ`�wPR&on���ƻ|�ᶰ7�ņ��h�fd@7e]��5����Q�]�%r������q��Q���n16��|�e�e!��ֈ�DwTB[oNۡ���r]�YV&�����˗s]��וyE��;t�t"�b��ֶ�ݛW*��fk���t�49�x���6m�!ͽ���e��P�<+	� ���4�=��f�2M�����ֲ����c��3x$�U�Z�����L0�ݚ�a=����3{8��&�������3��{�N�IR5�Ų���V����i��[.ɑo}����}~________��}}}}}}}}}}}}}s��������?�����������>ϧ����}>�O�������O��掊脓#�	d���r��O�W`�mSNvb �v���D$�of����{]�XF�:��ڮ
��Y�BJd�ټI
�ar;z�T�Xr��eJ��C�S]Jrd�\�mr@��-����6ϖ��}`��(C��ɏ����Y�4^\ޓ+�n�J�Z���Q�u�#�֏�C�T1E%Ż�z�3�䗘��#U�O��q�
VD��כ*;�C���Uf�O��4�TYc�cĨ!�j�	�R빅�nd��f����B�n�Y�@t���Kb����^��U����X�e�rSyl��b�W�ș]��T�y�
h]�N/�`�Ivյ��x m�љ&_F�+,�O����w��ܑ���I�$����¨�u���U��w��7Ǻ�����Tu�",�$t��,����\����f�*;�%��{4�LHzhӫ�����א����[m[�mSgv�&ػ��Y�ېf!ʌ���$;z#��*��ӏv "{�P8���[o�}�1����i�ۮ�6k��D\5�WS�/s��˄V����:�y��.�P���muwq����ys�̓��Q�ӎ��(E�$("z`�*�wK��=��T�����P����K��8ኅ��b��=tl�ô�����>ϟ����}>�������ϯ����������������~_�>�������������������>O�����}6�Ӫ���]�=����I�J�ken�������z�0!��ep ��v�0B�d�)ڱ���d�]+c����Kx��ӪZ���I�Ʒs%+���ֺ�y\��ۢ*Z庴z����M�/�7:?��lne@\����)��vk��'nR��2�I�r��<rv6����k�����u'Z�ɵpaų�E{a�u��m8�����F��+7T�2�h:�ܹ��v�ۦ��.#j1�\��6up$�j�D�?cZ��+%v>޹/�C2�%^�C.�e��x}X��gG����/�2�"%��y�%�[׳
QdC[밅M�QSW�CuÆ��:�Fу�X̬�=R�A��3�K<��@ԕCo��z*��%� �1ԛ:�z��)cj�Ƴ��{��,D�8!��2#J�8��o%z�E�Q��Tk����v�p�V��]rw�p��K�J-U����w*l(5A�Ŝ{�\��)���n��V���J� ]��R봯�����]��b�lŨ����5Ѕ>+پ�f�i2hᛍ�!Ӈ1���T��:�f��ȭ�U��[�7l�d&f��3�etܽ
8���&4Cu��d4�q���o>f��]A�;&ٖ�����ӡ�R�o/�ܢU��L�*p�㵅I:1ʃ��=�x���@����'�z���������������������/��}}}}}}~���~�������������������������������o�w�ϝh�w6��8�ac1���e����ƢxiL��5�+�6gQ��J���͸$���D���te�F3/w7[em��YH�8qG#f=��@`pw25��8	���]�Aô�%������%& �f��Z:^���+;B����=�A$�����f�[]c������7�%�*�%	R��Kv.�S{��]�o*n�գ�[mVŻ �`�f�l�*r�eH�6����l���ޫ;�%h册�x�K�b����������3j���O8�u�d�)�Y����|4&o�;4��ufE��&���7V�]�Ac�r�j�vv;�M�1Jܜ��O.��_r�x.��H�".��F��c�[̩�m�JN����͚�go���H��]Nb���c1�\0.k�I�
{��g��O U�ݢ�IZF���g*�����/��c}�pRR�0�� ��!��z����£W�`�M�m��6��͎��ٍlQ�G*d�t[[�;�w1Z�78s-2�x���{�Q��&Jm��	(���M3xP�׶T�e�s�!X��Y��2t�n�"5��ӑ� RV��V�WD�1��r�	C� ��1A}�5����&�^����K�����i;9�E<����nh�#�w({Z�M��q����5��U�	7K3+��%�����C��B���nC�N-[;2	zynLp�qе�!�ʻ�H�GvC���*��E;��!�Һ`�xz�reԙ�F�N������̧;iczd}�m��z�ew]�i.���\`��m��pKWeG5�}B�>�ƻ0���Q�n��ܾ��%0��G�uf��U_x]�2�")�*��Usq�f�1=g'،��|�m<��l�z[̚\SGt��R^��u����H�5�ҖipB�qF+��\�J�y׼Hy[3l4�N�n�ɤGv�g)j��e77)���KtW6i�]I�˴�����zN7�b.a[gumԫP��8��T��f������d|Ț��6���@�G �қV.۾<�k��Lfdɯ�|�B����t�u6�*��]v��$��GQ��+atљwk,�(�q,��E�΃��<'���Eei�u]�LIz[�@�5Țs����lS�k�s��f��nS��)��[Ŕ��3BCe�nU�D^�P���)�:�n�ED��p�[Yhk���18����.��m�<�!n��eX9{����l�RK;���M������Y��R�z���� !��2����I�{s�u��N��Z�9���y�	�t���<����Nٶ�(nu<̪���H4����՜�Ƕ��:N��Q�葖��9��w�vf>{��/U	�Tf�Y�ױ;Y5̱�¶J��Z@�U�D!���TZz�8�a:�,+4N �:�6�sm��ų��.V���`׺7��k��ؒ-�t��IN��}G5�a�Zc��Q�)X�Y	\��4���S;���v���k˺v�r�>X���@Y��e�}e�"�Hn����b�K=��͖��C�[]d,뱼�jJ�u5e��J������岥�2& ٿS��KAȷK<����0ܮb�ؼ���h���R�����9	Z�qB�\��o\���N�!{�oK9�N	']Pb�V�n��8�E�]=�Oh�Ãev+ARx:�0��`7��pfMR�.�A\��z����07��xGT�WF�Y!i�4��$�c����v9�:������9�@�KM�Ƣj^�:��2�<-u��4$�t}j͚�8���h��*'��ar��{��}���^�1Pxn��1�Im�1�22�v���mb�L땽���St�{Wv�p� ��n��w*�ȸ�49�N�)�`�`��F"�L52��F��5���;+9ɸu�Nt���B���]�Ɔu��v֊ζ�I.HQN����/v��{��E��N+�z��wDT��0G����oD'��u#k�cy�5���]�Y��m�HFշ1=fZ���bUݭs�pDu����[��Ut�g�/˸u��_Q�u5=P���B�v)���w%.���t��U|�N%eM㬼�NB]�6$�mi��
�	t@��}����hs=��ګe��z�^����Ц�us��npW�3�Zui�y˦�J�U�Y95�D�{iF@� O�Wb�����'bx����-Т�ʗ}G:���e)FF�˸ ˅���]m�@��M��֢�g"�K�|(M;������Y��\v��G�k��]�Mb׌��/��YEM电85dvzvR4/z����h\;�ζ�R����r�m^����LٸL����ҝ"B�-Rm<���,��+8�r�Y��L̜�Z�,$o ʗy���^p��P���34U2��8oq1�+��I|#z���m��sPi��rn��k�tm�U(�ԭ{��eH�Q7�u�k�G�t�|8K�s����s�>�R��O�kJS\�ke�� ���Kێ[�T:�P�Nis��C"z��8R����!R�L��pQ���˔^�W��+����D��-�,E��1]Z
�|��5�:.[��CJ6$�_3��;�5�.�Lٯy��A���;�U�Gr[�.��V^���'�Aٶ�bl��)`�]v}#���Z���B��o)����.WL�7@��9�N*:!^�:H�;|ƅ�Ƕ�攓&e�� �s����N��v�����@U��]\�}�/�-b��oP}گ1��5��L�^7R쁰�*����8m�����֚�꺺�@y�̍>�:�[��nH�l��𥓔з]�Vc�ԙ{]�Oಸ�lċێ$Xj";T�]1�Zq�ڌ�i��{����nT�4z���nŃG�1���J%�b�{&��h��0Y��X�
���t�J+����z�; �<t,?�j�&����qX i�bM�6��Y*cHS�i��9��G}X𓇒�V͋s6\}!�,Cyu����PXwT������b�xb���/$��^�F��H+u����[�sҴ�0���znu�^:��I;r�PZ��t&qg%j��;&t&&��Rnf̗M�Phk9=t�em�9�޳Ak��ڸ�$L�Q�Y����<�s���e�P�6��ZhJ�[�Ga�*�<�.�����#p��2U��4:��r���Wn�7S��u�1��FC��s���&+}2��g�S�K.ಮQZK�/>v.�rSlM��B�P;t˺�l)�m��wZy7i�6A�mJ��b2�����3^	Y�@����ةZf�xܽH��GQe�ݢPݮ.�w�Q��m�Vx�3:�q�X��Ĥ�f]��7��Yʻ��d�)��a�O2�g�A���4Y�;8V�ڪup��VC��@n�"㞶7n�B�Nf�\)D��d���$��z��q��v�U��ia�BڃYvb��.vvK\��n�V�Q��t�}�dF�5sMT8�]t�=�j���J���^I�Ȧu�X��
ͽ͡9*��Zd'J���m
/3d쮣�zf�U>���^��XU����/�ء���L���cz�N���_uJ�vEPh)mt�-�e�Ν]�1�d��rl�#��ƪ�cc!I��.�Ev�n�xG�WsO����9P�g���6K(�(Vt�벭�զ�V	��3y��I냺�Ѭ�!Qr�I�mP�L�}Ü&R��^�ZE$0+�qn-i�_J3���|_4t���hG3gM���Y�Uqw��@[��f�'(eg�����ڣs��톩�,|�f}�-��CK}FU���W�۩����Xq�:�5��eL<���nļ �����X�l�;�i�掫w�Dr�騦��1�֑��Dr�e�6ttޭ�
�Kz5U*�r�,ܡS��%��\�����1����VQ�S���Si���kb�YO)`�ֻ1uk�r>g���!�W}w�UN�E��Et�ĕ�]	�RdNذ}j�v�.���51�T�����k\�F��,=�ۘ��<V���҄!+x� �R���2]�-�$�Y��{"�: �8i�%h�%l�O�S��Uz�r�������/��ޯ*���_ϟ������z����p�q��X�����̧_��Ʉ��"�X#��Q[J���f�&�N���4У�H�Yk�rL�[&�7֮��̓�l�S�9c
��Îp�*c����R�^J���B�,Ks[������t�u���&]a�j��]ۦQ��Z.̫I��r��(7��a�&m*��PR�Ծ�ZN%@8�]A�ݎ8+��^-�}���z=��o.٭��ɑ�۴�e��wa,�Vܷ�������;#����Gzf����~D�
�5&I ��U����!���ńL=���ݰf6���ӷ\��@�:�e^b�WRj	��=��/;+��JW!L�����)\�\)�*��v�S���`�N���:�ʆs9���5��
�+��${R�me�d��lT/�JV]J���v`������YA������^'`��9[ndy���S�i���N�z.nw�@�u8v�U�-��\eK"[��V�s�o@��SQ�<�w]�\o(�Ke!X�����3����%���*I��3���ѼL!��V�f`��~�%M�����x��m��p����Q���K���S��y.)���V܂H�9�z�j�X��5&<ɓ5V ��Оl��tʂ^	�\�L|A�jeJ*j*���V�bP!&ɏY�78���d�i�bgz��u�?K5�IJ���R��Lt(�Lh��C�1�Cƍi�R2y�i�`,0o���}ʹS���**�P[V�*�,����hu��ƃ�mVg������4�A�b4�j�mMS��)b5�Fة5��5U&��4�iuEET�`Ϗ����ǄN�j�\UIE����6�QEF�\9�F�
�T[V�3�������hu�*-u�tX�bI��N�*k;C�8��Z�ڶ�N|||||(��&���'%��ƴLkl�c5DS1Eb�b�`����ɒ�F�(ň)�4F���1:���y.��TIN�QX֊($��)ڶژ�����Q��f�kS�ӍdӉ��UbMh0DI���m��EV�j��S�j"��:���VڛTF�1�V��mض#m&Ʀ"�1h �(4cgTETGlr�ͷ�s��9���յQ�U�T�Z&u˒D��8�˅R�O(�
�
6�93<�b�i��_H{��sʻ%�\LZN�K�rz`�ή�=/�0:��_V#{"M§�4w;f!bNރ�'W�6
yI�}N"p�L0f����K�Յ�U���|A�/�?S���R��tV�+P�tTC������F	@�.��m�[��r����~�������pU��3��]���y���"���)���&=q�7`� ���+���UOtu��#���:56��#�����ph�V�쿫j����p~��Lϛ���W�}&�T��
��:\W%�N�����o3��?Vs׽�:�ϰg�z:���#=}�ܟ5��(N<�{�y��us�~}"�0�{r�}�>���'r������4E
�`"o�	�ƃ����u�W!�"���+[W��M��;�t��}M�\���/,���}&U	<�+�ON�5��Ev>�uvjɳ�n����?P��n���s���ߊ5�zw/zr�o�+�3�F�t�X����=�oZ�\�+zo�߭�5��sFE9�RyG�������G����m���{�����R`�bK�Z됽�����X�V�%Xu��@�����dYX���p��:�P%��~婿c��WP���(�״�Ǽ�aͼ���j��qN��+���;b�&��c	����5S�29�;��ɼ�ِ�g�z�ѧ�_*ܼ�^���C�[��i�o���	;�͓}8z{7w���^��4V��\���*���%]_����+�k��iёkO�3����v}�S76��f�uzO�1P䦰�z�-�9���J�U:���n��j��<}}�~4��}c�?A=�v�irozx]�c�zDM���v�^����H�V���_o��q��o��E;����/~�Qk�g|���>wҪ��oW�wU�T����]ۙ�b��_�T{c>f����MHsS�(�u�;B�#�%��Z�C'����9�;:N��Y�����C����s�?|���G��֓��>={��?s�;�!���=�D�<~��ڮ�Z���c9�|1}�o�n���nviʚ��hNv�3�u�M7�5�n�FwC��V�u��'u��}hT�eyF�ϞԶwVJ߯�V�H���=�ǀmV�б����W�2k�k�R�7���[�e��Y�8��]ԣ�$+�VJ�(�vq��j�OiLWk5�yS0Xє�E�'����Yzr>k��6X�a��x~}o0�|�rG"k_Y�l�D8�֍�=^n<k���X�OW��ǈ��l�)�OgI3�����.a�dALhN�F^�yǍx���?eѰ��>�%�ޚ�^^Eg{:���/eh�����G|���:L5����X
j��h��r�����A�C�e���������h�c�߷u��9��ed��V?YN1���q識!��5!s�}yO��u+�fW���4�k�zs����۵$־֑�N�z�Q�~���aa�����3B���Ҭ؂u״�w���3�e'���k����-��T�[ڶ~�j)����n���0�vw��b�{��j��u*_M�����h}r�y����V��\�ݸ�j���>�o�/�����,����z�w`�b����Xјn�3}�/7�E��h��PCZ_���X���WӍV)��Ӻ�P5�+�t�kҥ�̥^yG�J�+�)�O8v�\��Q��>���[��0�o*�lthM�9iϚ�+����W�c�f{���[�TsW�5�*c�95�+z�Ž7��F�fm��W����֢�>��^��h�<�:�u�j��h���-I��nsfH����x��]�K���x��j�~�3��>n��q�h~_A�X�τ�nL���V���7蔕��g���[����������l�Gn��j����-�"����r��޳����:r�XA��ͼz���s�&K�'4����ƹ8��*��6�6�9c����o�w)�PkQ�������|�Q���4:��]_k��3��}�<5q'���"Y����N��6�wP虿A���v��{G���	��i�ɮ�l��)�;i����Mc)��������^78S�BFk���<ŏ��[��g���}��N��xK��{:5s����'7�������V�1]�V_�8��t�DǛ�y�|t�x��{����ɏo�ד¡�e�S���U��mi�]��oZkԱ*��C�${�D̪x�"��r����uܾ�7�j�F�-'!/�t9�6\3�-�6���c���X�,\Y��Ic٢�m�}�M�^���{��磿$׸wd&O�б��8�B<�u'����Y;ӔüvA7g�A�ǃѝ���7Oԓ�"� �U�������z^Ƴ`	5d�3�t�H!},U���
�xV=�dy����i�s1{�2�sz�������/4�V+h!K�DaMײ�r̲�׎u���ډK�ll-���(�^q���5uM��4@��w�f{a��ک\�a�1�Fy/zX4֞5�Տm����䝁l����c^�4�M�P9��^Ի�����KϖR��\�e��S�u��Yo�
�Y[֗9v��~����'������}�s�w���W���FOv������a�q��+��oVl�h{������\�uz:o��G�j��k]{s���l�c�5eNw�V{{	U���]3�x�ԩ��A�5{�x]�}����u��km���z9w�V��9�k�۩�kb�9�H�z��9��?_��{<����~�D���~��o�>�ە��8��,8�k'"q�	E�+���.|���X�:vV)W�`C2�oND0[
�K�wɋޕָv��iRP��*���h�KW@��\|�lh%]�=W���ˋ�s$	��2���:���z�G�z�*G�y�g��JB8��Z�ei�Dw&�mTE<x�i��C�6��;�I��g�V}2�X�ijb�u�s�s~o[��>��p���}��;����1۳JTv~g�S��oů'1�t/��u��6��Ϧ2Y��bA�s�t��i�dV����w�R�e>��Y�_Gu�Vc��ۺ��?/y��ǒ+�K�������/N��9��YV�����߲��2��:�M�6��sa��!yo���]%��_:���B������t�q�m_{��5x���S��]��'mߜj�L
��j�P���������.�+��!VIQ��]w�W��[��pU���f�����*�@��P��Z������`�b�i�H��d��e}�b��r�_�g����ٰ罾�)������xbʾ7��D�u�]�f���o��C�e�Ȭ��B�N��-6hl@��{��{���|�=�yq��H�+�T�bLf��G�<�&T;&����RWh%o�"˫�.`�č�R�)�{;��ɀc1�tټ)�H�7\�ʜ���v�l�fs�n�u�ʃsz�G)��R�;��`/|�ו��o|hu��?q��
�Qϟ�L�W��"	|syQ{S�O�8���6}9�eVr��}����Ktj���׏���>s>���:��y;j�3��<���Ool��m�����$)4e��	N�k�.�;����cL6���Ӳlq�h�^G���I��#�0xb�f�W��;�J�\�o��hr3&�=n��=�Ǎ�s,��=��ɦ̣��O���מ�R�ص������<G�R��L�U�37Ⱦ�/���{�re�UVA�͜虂NgPK((�㌜�9����\�g?m�ݢ�j�W��׏��Oy�g՗�����������^�K�k�7R���ɾ��8��~�r;��,����jf����{/�$�}�r`e�L}Qy{�W��h��jN��;�������}�m�����Om�	#��9�)Nҋ����ZQ<�O�f�B�y��n@�2� f3��=�d�%{k�r�u�e��5���*���q�OK���e�O�ώVmL�e���"y�m�&#t*��V��J��X�wF\�[޽[�u^)!S�yA���}+������]�=I�B��O�����\h�0�ڸ�["TIuCTo}���e䕗��+i^|Õ'�������p���~�'Y��"�u2�wޛ��"�̦o�Q�^�v��~�{�7�����{��.19??=вR��%/�������mg�Y�Vsվ�Q:o:Iy�z{1�W��?LEqw ~�%#^�^y��̕[bu�=ன�tSpQ�1W�12�X��ʬ�\���8����4J��ۡI�cǎr&G��g���}�zCt4��1q� >����I�$��[S܎�/!����.��}o��r�����΂��O�*��|�Yx�ռ��OzM���1�>bb�3�1g��{,��k���H�-�� ��y�W�=����{D��딈M�Mx����0���!�Ζ���������un���䧡��aJ���x���X��J�)�i�M�-)ܧ"���N:w&Zuβ���Pa��ے�S�&]F3�g'=��.�jGW͛ ��IeL��v��S{�{oT9�z�B�$͜�L��35ѽt&,�DL�}ۻ����r�C4h��'�� nD�E����9��`����le��.�H��B�l������v﬊c�ڔ�Z�W��x6��s��{�K'�fr{G��'��*y�����L�h�>Op�{��*i{��y��Ђ�ڬ�Oo�u��}:I���Y�BW�¥��n]�\%�Ro�x�Sl\�/��+���*װR�kO��|��K��Ѽ˛Cн�&�n5�m�ߍ�9b���q5��W�U:z�f{h-K.�/�'�i�M�f�-���*;�x�d������{k��tp���t�s���T��������H�-y�n���O����B�c��Y����(����2���&���
x�$��y#�=y�����j�X�Ի<���t��B�b}ֽٽ=��C<;��Pc>�x�r�%o��ԧ�WS�Y��I�}�Hω�S�;d��k��wj7����ޘ0�e74��- o��nhy�R؃p+��s�("3�3�j����WP;3�}n���& t$t�h1��nX��o\����|��B�/X�ՌQC�8!6m��U�0��pCR�S=�vΒ�w��7���-!����Ϻl�����{��^޽�o�zcȄ�ט}Nokne_�N�7ݖv��}�B�|��g��L$I�1cʹ�����{6�7�=n������%�{o��W@�$˂�ߥ��g�M4e^�~��#W�~��}1�}�)t�럤`�G������{�oŖ��Bʛ�UL��ϧ�8�1o�F����zP�N�<���/�c�I��Љ �R�v]��:�?v<���=�ڞ~���F�/s�_tI���|ǋM���gfU�.��U��K������=8; ��q�q̲���B7zݼ�e��zgwD5�e�W�Ŕ6����%��V䛿o۟H��R�8�K���������z�O����!n^UZ�5����m��`����%�̞����~}gc�j�&��O�0+�T*�:�?W��}�*���~D���1����@�xf6j%W�u�N���R�o����Y�i��K͚�x��� IfwS*�ٱ�f6eǞ�I�v��A[�)�����>{��֯s�+|������ˎ*��u��]ISz���`�U���ua�iR�5;Q�GOf�%�5cFks;(ʘ�@I�s�T���{M*r�Ǡs��;z\E�����v#ƹ�N�BvS�5�QY�4�=��:�A��ۚ�O�7�0a<��Ki*�)�����w9;
��cN��I0��(��.<M�-��������s1�t|h�c�j�b���^����F:�JJ��������=I��Cs���K��f<��&�e�,\�F�O�妴�>) s�8���W���EKT�*oms�@yovtDNb�h�z8�j	Ow~�<å��5-�� ��t��iǖ�|zvg1֯�@�S��T"�m�>F���f��ǝ���r�&�@M_�ѩ�n�.ʉ�.P�ƥ�.�m�Q��ɐ��w��xQ�cT���w����xF�<U��j��[n��1a�����t�:N�NZF|Fh٥t����/��Veð�.�뜝�!�(�=�����:�wmfp���#N4��}� K_,��x�рꨬjuA��e�d���6����Ţ�`79�S6I�3t äJ%��o.l\\y��(�����ێ�r.�f]�u!���)Eݴ��{IN�WS������f��V��H������󥽼�$ܩt+"�]c�%Y�Q��OL&�{�Ϸ�&�v��l�67%�����}I�i��gQ\`�m-Oxr�xM��%�c���XC�%EoC�s+��!ќ"s�m�7�y݊��T�@��4)&�z�K�b�2^���8S�%�D��7�X��+0���VF��K2�i�SV��nPl�y��+6K�4d��dܼ��7�
��{]�����Y{�OOl�H��e)�B�]Y)Zo�^��ɬ�_
��c�3:VT�jSs96�)�f�ڃ�-Im���o�*{Hc)����m$����)S=׊�.y�@&S���<l�Sj��Y[L�!ʩ{&_*ƭpnU����Y��N]{�I���1�wI��ܝ���������oY�ԝ�t���T�xo�7-�E��(�*���hP�.J��k���NFwl�n�����2�[j,��m��P��+v,3�()���6��.7�#<_N �!r�gm=�)-���A�B�Z�Y]�ӱ�o:d�p�i��z�������-ʺ�ƙ�����G�c�b'��q˻|����vN����v������
xә����Zx�7�j�Fр*��a�W�ˡb��BǍ�h�W�u��sO�vku��r;OK�{���ۛ{�&+2wV�&p�P�ȶK��J;e�d�h����r����)�O��)̧��,٢[�y�v��e� �x5΀ݹﷀ�H �M( �G�*�-rW˕AUlns���sh�<*����v�9�D���f֌�����|��Q��~{����c"΍jti(���¶�����sh�nsD�$�cm���Q�j8x�����<�����8\#�0Gg�բ�浵�m��;�ݢ�[r9�b�N.r1̚#�3\���أ��F�Q�nnnm��s���p�0T��|||x�1DE���s���h�\�9Es&5��n:[���:�1�51O&r�\Ѵ��D[cmfs�<6�T�`�������yy�r����r�-���j*�NOVe�D�l�PnN�\5Fq���͹nl�1�.Z�F�q�61�6�G'Q[s��c�q5T\�U���.�ªcN�����ګW9m��˅X�E�m͹�,4���]\�;mb��X��h�X�k��l\�m�b�\�D�b��sg�Z5�nsQp��nnm�6�m6��gI��&��qr5r�14�#0r�¬X��sd��*��4\���w�ws���1�ܵ�9�V�\��msh)�v�.�������i�v 嫛TD�ͪff�#�i+����6��QF��[Q���g�ەsjH�l��"��RZ�$��"@�w{��jG��R�{+b���T�|�T��{a-��͘`�"V�F�	م^�'U��'�����x�r���z���	�9�2;|\���ku�f�|(_�:_�\�����H���ǙUJ�w��Qb�6�efhh���0�	�1ٱIݰ�=�iۯ���D�o4����Pn�>��=2���a���	旉(�Rj��~���)��_xE����Y�w�(��z8��a E����V��������:�cjDp{��~��_�,��ii�1j.�uV�}��pWPĦ�W�Y<��׍����5uuY����evW��K9}∭���R��O�{�߱���T�U�MJ��Y�D�����.)�bmn:� ŖtK&�
�7#��O�/��f��c&�P}* �v���1�<�ַ]M!�W��$玷�����["�(7��k�MY���=2��GgIS��2eOA��c̊�^�?#g�r��,��`T;"���,?I���ӓ�Eg,�a�@s��P�ɦr���啙�������!��3���焿daF ^��5�v�BԸ�O�%@�뭞��W���~|+�}xA��{T�P���R!h8g��ɦ���F�*��&Qt�V�zi�(䠿�*t*Ƭ���F�Ɔ�^��y�N
p��)[�I�'=Ș��m%Vz�R+k��)�G=G��/@�B��0A4�����l�0$#n18<�$�s���xֹ:��Jj�|r����*غ�ұ-��1�!bL�3|���������i�� =�&��{%�����Ttq�ꑲ!�I0-�2d2�!G,�	���I�T-��۸�N{��֌��Y�����hL}:?#���"�T	�dC�x��QkM-�YK"���ŷٚ�E�m0]����-�c�G~q��u��s�����������c0��pjv��5J5��T8d���.��R�4���}��2|��l ��
c���[?l��
w]���A��I��z�=�S59W�}\-�4~&!#�{#L����ǵ-�����g��n�	�a��6x ��!DeE�7��F�8媋K�P4��"�q@���MA5~1�߭�`�xbŅg��,��ðU�\L�y.����R1BW��b-B�"&T�	���r���G��r&�K��Ν��X��KQ�p��,���1�R�eFtx������j-G���"�y3♅2ܽ�E>:��QGy�V��r@�)V~�aq�}Wj$�s�J���3����*EY���^Mg���$=j˨�G[Ϭ��
�+���`��:���"]��,�5\�X.ߚ௙��CK?;��_�?`Ӹ3*)L
��Qy�ҷ���;��v�S�����݋_^Mhx���vvHX+p��,j�ׂ�%��[�a�h`�+@��3�{Sgb�����!M}�#�k���h���3CMؼ�LA������ʭ����]$��w���2-ި�=�Ilm閽,�O���J�^|�R������U����G=J���.ǃ���gx�����='�쉣�e��N�F�*�+�̻R�7J���E�X싛�n����,�`AU�h�f�qv��y�P!h=�*�Ǳ�	u}�ڤ0S���*ד��f�-q1ɞ�s��*{��%l;��K�VY������L��7s�B}�rJ��,4��
RUYν����jT�W�T���T�G��h%*��r�Ҡ���H�@!q͹�dtOs+����B-�B{��C	^8hˊ9j��F"��y�↶}j �����jBV���̸k�,����T֦#^ڀ����@�vq�X	T�ƭ��Z��+�z4�:�5i����7{���ί���yGĊ)Oب5|�U��h�����璓-G5�]����l �;�����!�����y�EZ��o�-p��f�Q�� @�쯽x����.b�����Ы�6��O&N�u�n~�Hi��1�>��B9#X&�"mJ��E�j~�yY<�n��i�짔�=W�J����re��'p�d��Vr��$���>�`�����U������?�
�:�PZ&a�ڕ7Wm�/^Z�`�/$����}B�ә�0�ug9�]�:<�V���]b�*f��˘��Ѷo�����f���W۵�c����m�ث+�3\Ҽ5|(��3�B�AK�s��l������: �B"���\✈�雎�v��E��j�-C��,]��xcz~&�����k��`Z����5Ԟvǂ�����'�u�~�q�/�O�R��ws%����S���N�"�M���G+�`H���Q��&��5-���<KXe�5�ޥ�����3mu�]��1�d�4��ɕ�UЬzU^�[���[E9���ur|��j[Q�k��F���ޏ��#�ފq�����ftY����c��[t�=S�d]��tZT��{�+�B�TC;;�z��'����}?���rcx���wH�yP�k��f��1q�,$�����fYs��m�]c
E����uq^wƁ���(Lɽ��VR�q{�e��u�Q��6��G<����x��n�J���U��z������J �[�u������ۻ������m��=6M��6�ŪRSڈ��˟��k�X�g�gv��4��ǭ�9�.�^�L��ݫ,��������Y�+u�w����\���_.B�mϧɟ������˺������噕F����z�`.�T�Z��]B��Ty�vU�7Q:an�Q��ݻ���M%c(;K��>s�X��R��	�)��tuGΆ7�nn�Ev]K֒��+�VK�'r=��R���})ݭ��v�rղ��J��%^����˱T�:N٫/d]jd5���8�A�����3 &ް�UM�3qYllԤϝc��ܘ��v�Ύ^Z���ʛ��t<0+C�J7�xP�l,�
><�T�Q���Pl�������>�=1~�u�L-�^�tq��G��ݙ���J9�d; ��`(6�T�8�WW��f����]�u�n�ŗ�L�ջ*�>���IP'n��?O�ݨ'�t��ԉ��H�NK!��B�mz����r���kXbj�R�T�r�B��`Q�8߱)P�^�Ur���Xga nL�G)JvR6��ˬv�Y�_b/@�3WkE�&����t����G=��0܌��_o@�[��>E[���ʸ=dJ|�Yix����@3Ϲ"%���G�]W�ރy��zEz�f��ɶ��N�����#��L.���
�R��b^"[b�OSQ�a��M{I��%]\Y���::j�_Sc�O3k�Eem�Ql7��R?_ܙ3ţ0�������LDk�Ej��F+"�6�z��F���;����d�PYɶ�[T�~KkZ�ڧ!������☝1�2���S��9�g�f��fP��z%��1F:�pP�͞ˉ͑�'E���n��.(5XfR�9�&aR��h���RNu��Z�r]�Q�ꅙ�|:�%<��o)c��M�9gQW���7ZZ���8e������6�d㥙l�Y{Й���]F+	�k�NW�?����'�~��:�$��a�s������)��Sx�`���z�l=:���6y����U������H����/sF�S�}�����7=V9OE�����Y8�[2���A��5O�����[�h$fzap�W�$]Ŀ�����%��
03;�O����ˏ�yv�y��*�/y��_m���@��!wu܍�w����c-�0�b@���>(�2����S~�͞���ꭲ/�����?�{�oРm��m�sO⬋'����/��<F�]qǈWR�9��W�g{�坤�eܥK�K\T�����N��[{�����$m+
9�0B�.D�^O@Ba-�+�n���R���\YwJ�*��vy�8-l��݉�#m�+�?Y�n���;~�f��:����Y�^9h`[�]c�y�4b�X.gS��$hcU���F�����^��\�ex�{��ez���y"a������Զ�ն�u�N�N��[<}t���K{p�O.�Y�����bC�l�9g�+X_|�;LGPF�� �ޚ�h�e��flY�;�M�Y26_��Ѫ�`�X��&PTJ*��y]��\A��Õip��C[pхP�����Q��$�*��{Ԡ�Tw�ٜ��򾩖�p9ղ���x��"������#2�e,�s��s�f.4(�<�+�ʹ�{}�֡���{� t�b&rW3w�8�s&��o�L���r�ҽ��Z��`8��,�p�s���N�}�M��ڛ�W��_�����8@',�賖l+�`+�^�Y�ty�C�k�{2.�$������W^6[�Q��vO]�zqLlUVD5C��j~�|�퀾�R�R@<򛇆�:����Z4C�~Q����#z;'��P���e� �y��a>|F��tC�W]Y[^�Ͱ��ŕ���lR�.��*~�߫5��E��`�+��й�S�y]C����h����kb������9�x���jMB�k�"1M8���@�o	���:�h����<�g��g-�L�ja�f�O3t)M�z�#S��3C����g���X���G3(m�q��Tm("�^a��#���A~�	�G�Ċ9SU����Y��&]n�fW.�Ɂ'qf�92+cc�qa�)�6�cO��&�5K��ΗM�5M�i_v�j/D��^�d<�v���3	�{�?q����s�tu�/��I��T�X�ӵ D$��*�zj�O�Ct��iG,x�E`�&I�U�8�xӲ,��<��f�'��ĀǞr�}�.��*�5�A���T55��,��� ��s��Y�����K�{�6�} ��w�v�F^�*���[^�F� <=~Ԁ3%E�_:W���\�r����u]��w�:�T��s\з!�'2&T4^�x��'FIK�4����Ze&�{���ꪳ5M��x����j!�#b�{��8��*T8�6�=��q|
����|��pT]u���@�A��=8c�5pXeie��x�!�-��=eNYa��'U�������W�[umU9Z;.iU�h��tW-ā[wf�����d�$��=8g�+�Q��Z�W>�#�1���Zމ�gףU i;!��1�oT4m���j�G��<�xئ��0�Z��rxR�65�{+����pY�iW��@�e��rj��{츦�ply��(���	�cz�.��*uT����m�UB0.�rX�5��١
���+��5k�׫�f�7jT��8se�'mMp�L>��Bk�8r3�j��\2��ío���g}4�T����֗c�{�j2­5�놏�UD���G�X�0ʉ� e�D��D���!6Ֆzh�����Y��;�MȻ��>�^Q������:���x����m�1�[��i�@c`ͮ`����M�j��s�[4������
��w�[Q#ʒ�R�R�>>���R�!��#y��aS����sr�c�䏘���
92�~�=��A^������e�[��օ9�X��Ċ�@T��)�۽�y������k�i]y�Jུ��%������v�&���% �`�������sؠ]b�sO%d�vV�5誱q�����p�{�i����Ħ�S%��*��s�$hn��S� ��!��65�v���TѬ�ŖܿE�ވ�����X}�>�;��^�%���R��D� �{o�zm�^�px�����
�߂%!��Y���}��r��RD&��@M Y2{�"��Ң�\�~o{<��R�o�S��;4�x�º��Y\������m�1�����].�\�����Ur}Q_U]v�EU�2�<6ty���V�@ճY��C�pA����6��z��Vm�7�ٺ];�*4d�������"��1��W~3�<1���gv�t=1���F5o
�23$!�52�qʗ&�{�����{Ê����WwsW;	���V�Nt�ݔ��5H�P���j>[H�gt60���ڮ0���)�
����M/4����8[�۝3��L{-�|�!��O����p�#O� 4}j�=�9<�c��avٽ?VMWa�]?||$c�R#K`^gxh�,�Գћ�,N�N��AD��@�W����O1�����2|�
6Y�Q�a
�tI�ʩ?s���'=��7#4@�C����j�ǲ��b�m_oh��Տ���f�)�/�}X�v�usp&��0S�L��sX�.�ZM%�)�^�`�����1r�N����(u�����!�����"B<�G�#�g�z螽��u�q!/�E7xSm�W�¹�݇o��­@xÆqd�d���Py����qh̹��j�f��eE�ԫo���7�*����ۮ�c�d"0���0�a���1�U���^�=V�����1J�÷M�7��ع��gM?��ҥ��l}J�Mz��֥7�R��U(�o@� .oi�Sf%ص�e� y���ތ���!�+�b��ڦ�KkZ�S���-�.�k�¶~R��/a��֪�P�iݮ����� z�N���fӬ��|*-=hSՍ��:f�k5��!�lmU�˫����/�=�R�Ѝ�085ڍa��qO�i����B���X_d�ym�wNwu�̕-��������
��𿮗��u� �s���fJ�c�G!�L�WU��̵bj{W�.�^�T:Œ;��X���snּ!h8|k��KF���Zt�Ue���5���:��Uά3�;b�c+���cL�"�����O12�eh�w���qNc�2VY���B�׎���&�=�|Z����������)T��)#p.3�������#�X�e\.��L������wM�c��\n��he���RkΜ���:!Yy+RX���+|NY�h�]ȑ\ ��p!2v�En3��qwیY��f���u�%+5LPuլ����lM�VWMk%���F]�E�N`�n��j�<έ���p���g%M
r�b��A@���lİ�3F1#��f��K�ɣ|�F���a��ʛ�A��{�n�a�jF�Go)j����|2ng'Yuoi
��e�{��²ƕ:�*�����U��M�ذ��3��7:�"h6�S�I[v*O�ZFќ�ы��,IJ��յ{��ީ���� ���6�q�E���ǃS�3���v.���u(��}��Qm���3H:��{�&�d�g%�\S��nP�op%.�����JR��p�d�����<3�sD��u�*fG��&]go$x�l�tB��x��D�=�m]գb�
��^%�J�f]〘��A1I˴�P�
����u���c�}�s�9�f�L��V�F���,�I������*�k��A����&¢:q�m�)�W_�
�<���s7Gx��ݗ���=���Q[�=��kͧEmg�RRn�c�b*��\@r�@�����[���EԦ���,��_x�X9���G<0���6
��un���ȪV&���Y6�訒Vb�jV��L8u7k��ev�xV�U��@��h-��虬#L��N`<kKxm���1����=%��Lol�8X��+�u��+^�e���iǱ�*	MZ;/01|�۬�R����������[��(�9e�K.�t��#�p��O!Y���R������9�]��γ��O�L���=�"j%KP[���U*��� Mޱ8�W�G�%�T{7�5�"�N��Z�Zr5����]-r�r��G`ֹ[�.����枕��N�q� k;f����p8�eS���^5/t���cp�ם�/5o2�|jnٱV�jk+��#r�m��cWŪ�[��QXo7S��4�r+�9�R�/������b\�5��Bد*�4	����d.�yaiv(;S�ruc���=�ʝ�Y�x�xԘֺ�[MMZ"f�7u�����m�g&����u��֭�V�T��k�� P�)t����[�F�V��7q�}���#)��Ct�g����Դ,C�rڗ���!�����칌
W�næg/���5b�&���l�O�Α�QnWZu�/ �������:� i\��ͭ��&ǐw�=�R��t��%�����k2����m��9 �l�d�=����as��kR���YS��J�ҧ�V�a�T{-��8�2�q���cYS�v,7tj@�i�`�o\v�a�,��୥��T6���3m��Ǚ�V�fͅ9�umM�e-un�ܗ,�/D#	�Ք��h�(Zj��;��*�r�)��K}I������]��_{�]r�f���k��.���P�����Uʖ���$51�L��03��=)�(u�~`�E�� 	��
���>�����~w�����7.SM)��ō���SUImQmD�iӚ#mkM%�b'����||Mx��裱���{b#m7k8��5��sh����QZ9n�,İ���8�������&H��3��TMkA<�
���jcY*���h5����>>?���N�"��&&**��� #X��ڵIsfn]ەܚH��������y�ETU1IE�E�Jj��1�v�T�h���i�����54M5N�J�F���@D\��*��q�"'mch��TE��򢊊-�LQkCMEM5DQQUKi �j#lI�"&&�&�mTAI�nl�G6�#Y�9*b��5���g2�j؝�TZ֍0S�3fш5��J���(��1���IAD�'cTELl��
c��6�D�T]ت���y�D��&��A����$���A�����]��n��y�vF+�t�}lҜ��.�X[�h�E.����K��tV��Yu�2I	NB!�N��f��{�.>ne���='��4.�*���y�=Z���y_a0U��y(xD����.��/��}�x˒��b����t��df��.f���r-�l�Uk���ػ$�h�LߖrZ.O0V��A�§?4�sd��a�X��B�4G��j��Fm�,�)�h�ν��hf5�G�"'����N(J�~	�i��"÷�R .;�R;�5;��+�LC-���g9�Y���KxZu�Hނh��q���>xZQ���T����� ?99ɇܜ�VS��.��U]o�0�x��!�C�*6�,�͞J���:��W�N�T��4,s�h2���nQ1]}�ץ���v�^y���U[�}kAֳ{c��C��I-�-3r$ǲ
�v�]b�br�3�bK���T:��٪��.��PSĥk�΄C�]�t��l���5�)���Z�y�Ҿ�ùAz9��-�.�A[����[�X�����ǭu(�zm:�v�X�=�J��s����%�Uf�����*�"=�(>U���:����i�%��e[��|��=I��|q��Us�6 1l������N��qG�gNTfћ߼��=���`��c[�f����_<Wlk>վ���x�ڷ�T��om�r�I��N�h�F�;Ml]a�OvM��9�d����dǙǞ}���)�c{0������� 5wbEʌɵ���F|��B������_�uM�ZBL �í�T�C����2A�[�}j�zj�ÝL҃2��F�Ô觊c��T�d+7c`�\�75ӳ��C�\��Ѵ�|�sh�_L6�lz'��t��2�o��LS��L��A��j8�
5��_"���٘T�q�v�N}��}	ѹ�0���e�9�ձ�����YFK%���8q����hœ8�T����_�������ϝ�����a&SN�{�ݜl]��K�ݟq���_�K�LK�7���U]?[F��dַMR�	!P�N��BĂ��Z�x�!�-��<z~��ޟY$�3��妕]��U:�cg�0��(ه���fM��}d(�ă������
�!g�^�=˲���>O���
:���SeōQ�oH�3�љ�2���@��a�i�������a�M�kʼŵ���K�0:c#7U�ZC�|�Kքҽ��l�؋}3�Wz
J�:+��lD{k$9��
����5}��YQ�V������RCo�9��t��f��Sl�t�=뢙k�h�i��7���7��3g⣛���o��[+�9�ƹ���k�T
�0����״rx�	"����4��3�@�;|��+F�� ���^4�zs�-ۮ4�P� �x��Ô�4"ǰ�iT��7�"r�`m�]�s.�;7:]���0o3y����cy���JW�'��y��~�u�7ve��^l�0�l�r$�l�)<I=�"���G�� PSN]~�pZ{C�9���>R!3='h]����Z�.���j��Y��1�x���^�p��O&�Y%�T ���Y�F�Q����y��Xzoo�&#LǨft+���Z��C'��;%7�R��w�j!��@�H]����'��[;����s��"Q*˹p�$@.�����<� ��Ss�t�jʛ�8�S��,>�)�mn�~��p��X�����V'bD��Z���@�� F�<��]0�UJn�J��߭�ɛc/��n�z�{ojzf���t� ��T#f~�NO��n���͎��t���I��.�m-a��6�@��y9K�/BR���cP�`y���N�7�+Y��t3Dmn�w�9K��Sq�8X�R�M�q�.�_u���F7�_��-��D�І�<!����۸��1X̧�y�3[�;vCZ�CTx��η_>zb�U,߆�Nx�`�3��<�^�6��#�=��^��1��������,⥷�t��&�"�>ԧ*沿b�s��m_� �gi��g�ކ�dޤr
o,�m���r�m���k��R*p�"]��t]-��ɚ�)VOa�]ZzXm�H��y�Y�RT�;9V�R��:��~���0oy��v��(��Z��j���E�Ih��^�| ��j[%��0����h���c�]T�T�n�u�a�u.�?C�0ӽ����z��>��((p��\��5�bv6�{#�Z=�lԻ>x1g��|i���$F:�"��J�P��s#��&gK�����f��������u��<�DwG�!2i��K1Q��[�&�2b���E�{� #~�� ѐ��'�-{6���Z��AS8�t�3��t]�X3��ߊ��}b��,z���4b�c�[�EWK���r����O_��җa�!y ��O�.w�4��4��Z��8�׿��m�z�:o�����;}*b��W�a��PY��Q-gڲ���l[�O=;�z�>c˕"�ɞ�����m.h�kBZ��^�`m�B�l����&t���ɾ�3?WE4ψ9�|(lE"�F����G3��<,mX r�2�#�>�4��/��#|1=�9nyv*�s�V���������M]���5�Vf�ˎ��B�Ǝ�A_)K��t#sO�VG����a����ܧ�g|�P�j/j7��U��C*�*��7�=4�qR�*Ae��u�\����:�G�u"J�󹝋:z��� [FЭ\�"�t��s9-��F�8�*=l�\��</����Gc讯-N�҅��,e�
���Y�Y��|������ɝ%��k��i�)j��9 �WYt*�}w���_���(�%M1(]|�`��W1�@�ePg�`���Tk<�|��(���w�>K&�'KRݝ�Μ�7�Q\�x��
����4��/���8�ߥ�sץ�b�-�bX�SQLbfr����*S�:�KW+�]bx�##�[+��nDwpl�2\�O1]F.",e�ڸ���vX$�eB�~�*D�}݀�[As�|r�4���OQ���P��$���ޒ�r��ۉF�fo��,\��]�O\�dQގ5�;N��;O�=�8cm�󜥾�M��]y�ڋ�8��POzT|y��R��4��5#H=�q�)���^d��L{}�^������D.΁V�	$�}(��/>Sѥ�Ԯ���Z����۵r1�,��Dc,4�fk�|�"FR�6��E��ϡ��#]}����a�k�E�oئ�L������{�5�!S.��dQo�M+��|R���É�z��ڟ�)�M�/��A낹N(J�����Dc��AJuf���k�!�$>�h����B��5���C��`w��gG��ˏ���*��%�\ ��Ӛ����J����t6�
�.�&`���.d���6V��N�1�1]�5�us
�֔&є�����}G��]��/[�����U������J��B�q��;g+,���6.u$�Y�k�,��p��?�A��H� o0==�T4�DK{�M��/X�څ��Gպ����k�
���x7����i��c�į��ͺ��F��/,���g��o��+�K�/5Ws�YX�jGS�W﷮D��"u�K(�j�D�F��e*}/�vl�j2��O��b_%��	L{�C����>�1��W���Gsbi���w����=�v��Sx�ڶ����Ѿ��~��Mw#�-%�=t�Q��� *-R�'�.;*�k/9�Q�J<��b��]����_]Ķdd��*Tt�����L��e�Қ��H6\3n��u�钝`Oǟ����Vn��_���ጂpy�;��.�2���t������{�$%]f-3�ծ��ݰQ��A5)�|
*S#��ʹR�ç�nz�j#�~�=V���]��K�xjCKG7Pp���G?Z�l���L�7Ju�d�X�0�r
w�:�NNu^�.C��j�|�k!�$r�T!�ZdD>žq��B�R��rިO����*a[��͉G�]����bFy��Q�-��� ��ckA���+尠�}����"�y���X���a���ލiKޔ���n�	Ȁ/kfep�5�9$����R�Oؠuc���[0k�Nͪ]��݋C?h}��f�5}�+� v�=�gdzЄpn�/-�/(^B��6۵A�W*��:�S3gX���r8P�=ɲ�����<vP��	k���྿(~Xa&@�U�}����}=,uU�b�~�ХFE��z32��^�9��Ä́��sXR�"
��r�U���D����Փ'ګ+�Y[8�����8m�����Gg�z�6�kIy|#��\%3�ͫX*kgWB6���b�&�������iR3X�w�4�P���,��i�+D�u]%��*$�'	��;.�ؼԤD�ٟ/&�5���;��u"U��5,U�KA��Ɗޏ`���2/bb�tm�U�_��i��1��j�Kpr 4��j��p��t)Q˻�,���:ފ�T���y��g�X��Z�X�(�������'���g�.�#l
����Jױ��S�3�G(�K�%���zGw�M/_Q�15�[Q�)J�|����rQ
k�މō�!����;9�m��� 9J�k�e��ؖ[�k[�CߦJ�?kH����rߨ��Q,,?��(˕�Gy���;��-��z^� �O#����L�Tȹ�.��>�Y�l(�����V���M@��̽���!�ehi�V)h,}�	_Fⵎ5qޘ���J��:���C�4ܗ��򻵬�e���R��{�7Y�Ӿ�v��}�ު���D�9L�4ފon ����mQ�@i�����W:�Xe�������{u%��9!��T��HԨ]�7�P4�T=��YLS�����h�u�Ѽ0������W�U��]3)2�@ҡJ�b�������}����H}!x�0���ِ#Ӕ���!�8җ�JJ{Q���<�k]}��b����^n:Lwt]�/�Z��NIO�Ir��ͬ�N㮘3��n��{������Y��*�r��P��\'";�u��R���(����+-�	���y�1�q�[���3u�=��7�j�YxrS��B������v!p���1���9�)���^���{��}����^��?�C��.w׃9|���zv>&=�3f~�5��@���L\e��d��5Ї?mpCʥh�yW�`��;ڙ
�K�?D6���~8~�r���=�q�t�E[ �/7���)��R���)�|D���9V��2�FH.gXsY���C�P�g\]�h�J������(G�upZ�
"6�w5S����Zh(c������HF�r���5ʋ9����ݾѓ�hkV���6\=A�\�%fL�������K���@�1r��9�"��b9;/a�N�\���[�0;:��;�G�8a*��Xn������h��"<�T�s"rU���d�U�y��,	�sW���/��=v���.k�t��.��8���^7B�ӈ�6�;���E]���f6Է�ϟ��`�Ǻm��J&�Z�H�j(��'V�s��>�;0�r�q3���8�A�LX1�C#��
�����
Q2�0�*����p��	ՙy���[����0�aXëM�z�L�x��3k�Q-x5e;	b�p1J^ԍR�����+_�lg�g.�F#L*��C�OQ1c��*��MAdK&��[T�~KkZ�E��:S�謊Q6�0�pr3n���tx,�3S-IJh��蓏}�I�:���dSdђ�EA~Aj��s2����y�.m��B��^/y�~K��`�� �=�/呴���`j2Iڠu\�w���*y�2+�0�=Qr�����G���Ha��z��f���vԎ�!>�论���6g��P(�6_�T�� +YC`Ԉlt����r�����Zx�P���2����ޭ��mL��oK5��l�E�y<{�ܧ�n=��0���Ϭ,�끻�Q�/��MRV�����q];U�����)�v)���&^�\���7�4��[?pr�N:I�Ji�}]|�w����a'�,ߋ�򜗽��z�q�Tp�L;�6�����6ș�moEGW�_�	�&W��|�>n���Rr�.;P��Rz<hu����q#C0�p��|oN*�!N����w�y��G��Z���ږ8S�v�ST\Av��-�!�ض��������,���P��\���;���v[�ջj9�&}����J��:�JX�7d��	��iI��NΖ�V�	����Ǿo�`aY�fP���o'3�������55�����I��x��]X=Kn�ձ��u�A��1�M�'��h�9x6�C�zp����BF=����
��XV��n߱O��4�[cb|l-lv]]�ջ���Y���ϐ��L�e��0�a���3���H�	^�Bѭa���{�}���6D%-^ۡ�׬~��Y�)y����1\��Q�/I���,������@��I����ױ�ڷ����ڑs��ؤB�Pd�L-�Kְj����Ȗ����'���ʌ�����:.Ϻg�Z����t	K�,z���wGyg����)Niv=G8DQ�>�3�w1�ml؂Y@���"L�zY	��}Eo�а	L��yUC��|h�v�qj:�1]W=o'c�f�W7[��m9��"��U����[r��v�zq�<Q}���P��r?\Ȓ_���rPފ�1o��3�A����x��&�X�zY�C{��k![�ފ�~���O���E�@�mu���e!�6�̆i}+��x���x�:�
�l�7coh�lň~g��z�����'��=�%k7��=�qW��S�+r�ἳ��R&�����tkm�N�V���HrŹ!�T�Z���÷�V�^.W	0����2t�I��`����+�%9N}�;	��G`ŖG�\b�|���zP�U�;����ya�$�}�²�Xܲ��\5�h�I��ڳQ���R�ƺV�E�"+�/k���nN0�Ǩڹ9Ŋ��^QV]BJ�ܤ������}]`�3S���ݳP�=�S�Y���|����Qpu<��n�VIS���8z7*��A�l�c�.w��vk�kOB�7
x_8�����f��@ٕt!�gk{�%d�:LLƨ�X\��e��&��i�V��N6�`m�T�e�Y�C�a�T��΁q3uRfj�F�B�ȶn�A���.��{t����si��M �J���9A����K��u�6�&����<bʋ]e�zfh���6%V�]��{Y)X�Ij&�J�ǣ�%lZG�Uk���M����$]��&�m�A�������YP��|�`�g=,�^Q�`���b��m��V�}�K?>a	M�bl��:N{0(EJ�o�sT4�Ǝ��GS���l�Ȟ�Iޮ{֎�{4��*0Ω2�gL;��@�#�eh,����ޅ���ՠ	+;�^FoptQ
b �|�q5rgv��v2u���i���?��+�yՂ���4��9yD]��Q2�8f�:�Mĕ9�w�,�ꋎe0��c���5h�v�����]�ue�
����c�(�<�_�%P�y�|GI��T��~x�k'�=�{pe�}\o+�}�z�tށ�H-���Y��}۸�#6G]%֝�U9,��N���Ѳq��GgwMwj[��w���-WЭ�b������͠��O#����)w��(��q��Y$�,R���d�5ͬ0���X�c��Mh�,ӂGqkC$�^ع���Mޮ.+6�Z�֡WI��2��� V�����xF7���IH�Y�Dyô����6�V�����7�j�K����&԰� �/>�Nģ!�H�ӭTz�uv�qΜ9Fm���hۖ�۽��Q5}:����L;u�1J���+i�Y�\.�ϛ=�`�L+h�b�_�6|�;�����&j2��q��+�y��%HZE�{a��Yd��lPy��K�����;1Ȯ��%q���sN`{���xF��&�O��+kS6�}�(��!Y"s�����j1;X�@�ց�N�۝'��.�?��GV�l��x��ͣ������n*)+�F�4�He��k�\�g.b=&��
�6A*c[okW	w�������Rw&�f� 
�?�TV�f�f�V��7#�� %>Zf�6�\�ɱf��G�o��(HYZ�,V�t�Z�
���*Ӎ�6���"�bh�h�&"	(�i���ٲe�Js������UQADII�U�QA%]�*�����#sfb>>?��|y���QE��1TQ4UO3����#ͻ�j
b�i�������UIj+Z`���&�H��M3k$A5Q�j(����O�����>���f
*����+a�m�����o��kERQDDh�L����Dnq�DEEC45��p�͘�"�9j�����jH*���"*b"�������hh������4L��l����sjH�����^A�j*�(���cTQPTD̔EQ1QMͦ��kQUsb*f��51EU��"&j����*�+N�sW"b����s�<��yU_���0}>�57炕��R�a ����u@ Gt9��Xvv�%��R�Z�	g��~�����o��^�oȡ�ei@�P�T�@i_��~O~����o~o���bz��2O^� <��&C�^L,�\�����0��GZ��gf���v�������n|�7��B|r@�8��<��뼊��4iŀiO0�WO7-Z�M��uձ9�[j��D�`��5�j�i��"�a��J��r�_]�f�{uJ������7�=S�5�9ג��ati+���:�7�����	<�D;�m\�E��Mvy�ZwF�k4��4����V7<��ǯQ��F��Z�Ƃ�]�v�W$���'a���{uz��B0��e�|3V��ہ*��d�&5ԫ��`�k�}���f�o���1�B�Gg&�@i��=���ȑhv�m���G��ޡ
rM)�qY�r�M�����({J�������S��wQ�#�q^P��.��w���̩[������c�B"�7���m
�h���[�@��ǅ���'�6�{����p�s��3l��:a���Lk���SG>��y�b�89�h����^�cposLFYV,Tͪ�g^δg"���NP�X�3�C�rᗛ%ݵo����k#���k�um���l]w�������m���D��i���i=Ol���M��n���Cy�*	�k'�b�i�ٵ"�j�S=*q�.�%Bz�t�:j�t3С_L�v��r*��b7׮�����K"��xU�L����aw4ɚ7pn�����ߐP��L� $0
д�4��*������~����[.W56q��eP>Np	��CV4��U-�0�%��s��FB���H���eTgZӗWn��i�gŐ�馮�,��l�.����U�œ�o�랃�c�����+�z��;ͬ��"��B� �tIa��aS,y� �m�eM�)����[�T��4߷����x�Q>=,�u0B�r��{�Ϋ4�9�o
*�7rSM��P�V':�vO]��뼹Y.����c3MX�M�K�24F������Ud�y�4��iQOqϻM;!MUڳ���p��e����Su�L%k�_�@0������m�1�����˾�?E�á�[��Ք�Ke���OaD��j~�tp�Ո��b>+��OIq�2L�S8f���wy�L�ܘ6Է�����ԅ�{���YՇ�p�#s��M�łsSU}N׌�M��W���ة:�^����쨦MQ�4���TS���eZ�
��I�����(h���]����-N�Z<yL�P����Z�c�`Ɂm=6�p��c�VzC���ݛx�VϋRc3 �?�o3D^�i���thu*���[�����CJ��g����B��kz=���.�G�L]���4��4I��U9�ˡXw�M�j���8*�5ٽ�S]�*���V�]��_b�/R�pn�裩�ڛWb�9{Z��l�%�&��U!.N�;�1�O������Uq�����Re�@&A)U�"_�����_YU��]�'�-?�md�V1q�ֱBB�.ޯd8|�>��`��[���%�V�?\[1��NI��C��MA��D[h�HL���1uΟ_��DF};f{<H<�D�|
F��뷻��Gܼ��P�Rr�06�;��O���>I������yP�tv�VDA��ޞq�wy�u�I�{����=v���/����Qc���gz_)�)_HLE�S��Ȧ#:�[\ܷu�v������Q�Ռ�D���{>*K4�9W5�}�Ƶ>5(��*|�L/
�Q�{c����PfT���0]l��3L.�����V�t4�\K&��M�
�ּ��+c��8�޿uj�zf�9�L��s����JG�1ǝ��m�yn(�ֽ��V�Dx�i��wM�D]���x���/�b�,����k�	�������K�n(��q�L�eP�.ϓ9u�e���u�bӓ�<�gXɶ�Mɗ�v=�^�D	�1�����r������{�,s��ܕ�w�i�Qge�*�:�����]ݎ��GW\�}0���NCt��4?A�}��P2mw���sr �R��[�}�������}b���ϛ��}�-�3�+\�}��E��Y�w�EiX�}�+��b�R;f��Q�ְܮ�̤4kaA�Y`�6�e��B��[�x���Tr����2U^��D�-,�2�@�"҉������ �f���8��͕A����������e��\�j��F/��f�wm�o��1(dG��wO�1N_%���w3�3�:R�qԀ�ζ�R'��@���&^�r�4��
2Yn3�A��.k6��ϺXǓ�7U��WD����P
�-:Ót�@h/e�
בӦ���0��4'�kg�~����i�"��E��w��k^���p#i���m�@ެ5{-.� \�Y�Z���lthr���V9��y�{��GL�)�t�>�|&�*q# S=fR٧�w).C�ʞ�T���]qk-�f���'��Ƽ4oaΡK|!F�0��`��#�ek�<��{>	A}�eۙg��2�;;=��گi�7V��=ܧ��0���5����+_��8�+�LE�w9=ܒ�Nnv�e�a�9<�bb�,�`p�Q��f���P��&���D��ޖTgG��]���/쥙�Eȭ^j�P�O!�e��S�SԽc�jq~n�3����1����PFD�5�=���k.�OfVl.�`����}q.�|�i}��L��e5�Ơ����^�|4����_���XU��!����6�Ԕ�9�c�u_����e��<Ŕ�Xue����"�·�4�[�kh^v���� w��i���Ǜ3�D*�	�4۩V%���Y+���+��1���l�����j�>����̽�1��WU�׾̸۫����ͼ���|���� {��f(e
P@�>�O>J��mke,篒]b��	i��C�T>.����_G��<��T7���P[��m�T�<�K��D�jd5E�?s�yOۙ"����qw�[P�@��e��m��s�A��-DB�Y�짏��y���:�uK���SB�s_��J}ħ�y,ٱx�Im>��o|^q
6Ge]l�M����ّ]W�w��K��r��h��F�ɩ����1��*}��f�mɛɋ�;�}0�>>����껽�����mpM�t�=	t��c�{&�a�����:yzw�5��1�u�1��Fw��G�T!�]� �͢��O�H�8�'�Q�#�TP��'�W�Z�`�����Y�YX��+�7|�8��eY��Z)��?B裒7和C�[�cY�q�̞P��[D�Y�1���:�qzL�:��W��i��[��~lO�$�T&cS��]3�7v��*j]*�z�iH�����30���1����7LG7�@zZy�;KK��]G�f��4�@|�F=�Vŕ�ڸj�1�≌k2����H���Gӵ����?=R~��j74�Z ���@�փZ��4�AT���r7Qv%b���m��o��;�ͤ��ٛ�׫jme<u��"%��WϻKY���B�H�Ap-�X����םN��V7�b��&sB��B���\�[�c������($�0��(�R�#B�@�(-"���	���|)��'O���:(т��|�r���~�^�=�TZ�y[lz�{�5��9��\RηR���X�a�GE�"j7��_mSU(���jX�oA�����*:�W�&.����8H�rA���&���&�[j
��m#=�S���`����l!{����~�s�U���k�c�a�(��^(H��U��痥�!�[!85�������C��I٩J�Z2��J��iP؆�mk�%3����ozD����`L������1+��_�9�f�_��M���޼�1\*k��a5�����k����l�~�Kk[�e8��z5uD<�|w���'O�uo4�}K�����}=Au��x�ḦL���<��M��ˬali��i�c
���w��D1�����h�zԒE�Hw�'�|�]0��Sw2D�</&fٚ޸y��EΉ��id���Sp�gP� �c��``\r��8�u���i
}�oMVٳ�C_NL��ADV�>�xo��,9Ƶ <brAO폋k��Om�>�{߮~�.'����-�5���T�o�������bw��"ŋ��4oS�jƭ��	��7Y�NՐ鎣ϟY"�}޺vm#������2o-Q�[3������G5�=�k6]��<K:���	y��"��/�++)$v�3'Pr�����;���6�|<��ŧϫ�4[s��	�
U&U�h��&Ud�C0��<0��B�s�)cp�Ѯ┷�<�P�	���K��J�k�O��Y��׾4�+��O"��j��;N?)��2�;z�6�5j˪c�h�;��U,qžx7��u�~zb�z��X&���3�g���
�w��!׃\ax�y�J�"6�"Mftg,��#K���������j��.ݵ���*jҝ�[g#y���lIaWE�\�}*D#��H�<�# anuoD��g���Id�7M/�K2ϵ�����)q��\�7?zD5y��}#��H�������u��v��I�.�C{��>�t�r3��]�ݻ?ߧY��Q��d�M0y�e�=5V��$k�-{�r.S�$���<P6nQ�E�^;F�{�Kf,-*8f�3�<4ʂ�Q�0�����Ξ�̬��n��Z32��n�n�`���^˰�څ9ba�R�(;^���V�g�5�WJ=����E�O@MG���a��ª�za�Ă��'��\�e��vK)d���eʯ�R��~����^$=���LA��j�fU�=��s��;���x�O\ɱ�;}}�q���4��x9ύ>�&r���[55N�5�5t��Xƙsz��pg�؅������Ɯ?���O�o�ٝ���u�mqeJ��9�ns��5����;f9�"� �^ձd�8=z������N�?]�����M� 	�`�&�RdU
X�Pw~�_�~���*��7x��?����/�M仵�	��4�C�=�럳v�˖ج�t2�)�j���2)�(�zb�2_[R�C+�)x��M�9����VB��ǛI�s�P���ݦ��]����EE�'������s��Pc�tF0�T���߬I�O}oXEK:�×�3V��f:�����&�|�p�EE�p%@��X��\��a'�_Ph�pL���ng�^���˹��E-���y3���7����-~E�}������`3���Υ�jC��mmv5ERv	��{�@K��0�Vl0�PȮ�������1�7��.��|�F�*!�&N&f����b��WԐ=)M�I�����52�v���=���`.�0��gN�eо9��1Z�{���5��^,��W�E��maP
�ZYZ�c���?��w��lg*WB���m9v���2-���
�홛S��V�$0�D�7�]�C�r����3���D7)Ӈ��&�P�i���ݡ�^2���d��34\S��HnZ{"�BL%g�MY��QC���tv��o��Y@�뮾�>���(>��9WEg0���y����x�YԽ�6�Aq_m+�N��Q�s{1���cVr�����va�x�J�"6S>$^�;�� ���:-� l�mc�'��cz�q�c����`4>>y���~�%L����H�Ȋ1 ����~~�_]��o�!����C�^��f�2wk�;��_��z&Y�1U	��[:z�}*��Kn2G�	˜�Z;!�	�j0!zT�=Ľ�_FG�RK�3J�ɵ#�� ��W,�V�&%[?�1�U����(Q<c�j&S���_�Rz��-��eٙ���x�#y�7��ù�����;שp��Ώ$�fǚf2Z����gz�o��2�G[��S	��y�� ��n�T�5�@C���[϶�ЭFm��⹈y-�.� Jz��ZQ<�}����T�_'�,�=�HiV܄����0Ysߖ�'��]�3�M늯b^ۖ��C�{ME�3=�^$�q�+'N�<��st�1��z��sP��\��*�nU��V�����^4���������Ϸ07��˸T��{,T#��k������y����m�s�=��݌(Bw5��U�-<��7��D>�ה���kOb�Zb��`�&��'&MJm/��J�R+�������}�y��]n{��I��v��mE+7G&Ӎ9���̮P'+ca֯����z�y�Q �(�;�Cְ��z�8nC���/�����.:7�t�9L��@����8���7�3��
zb^��d�B�u�0Q���Y~�z�U��Pa��<܎�p��z���4�2�cX��o	k��4�Y�4�)�H�0~���z�q���=n���@�0
L�3(�$�@�PA*(sߟ9�����ࡗ���%)��9�a8������<yТY�G$Cv��C�[�ٽy�q�vq�c�̜%����U�qٽ<��Gs��Ѥ@�
֒�,?��	k��=����^5�r������U���*)������ĝV5(1pmG3�UM�^��^��A�([U3dT���_\��~��}�XPZ�\�s֬�����cO���8U��zmo�#���ã4�{��$�c&�s`�Lb挦t6+��<���^9u�g�xP���Q>s���&]
�\>���ܵ�����)OpU����\Ð#��	5��_��"����� �;��h�����zU����J#6<A�rW*�j�Hn���CU�Ĩ�Eu���T�O�?M�jE���S���(�΀0�^�f���}4�P3�,��h֔�{⷗����j�������������Fi�c�S[g	�iH��7�"i{��0&k�[Xa*$��I���U=.��;oZ�����:��^-^�S�ܡ���G6u���ػ�[s��xHχb��1O��ݵ��hnX~�t.�tW�m�{H�3��1�s�Xe�rr���K�x�ݥY	�F8�e2�^d��*�y.V�ۑp��2ũ��os�t� tN��7�ǖ �*R�I�Ҡ�S�:_���z5�O[�o��y�-���ua֦*�7�=����tu�QŮD��Z%���6��Υ��(=�n���JE�����AFM�Ʌ�%0��4�E%t����{��)F��־+��`�G}�Ԩj�V�Q��rMΉ��v��A�Ȳj̩�e��7(S��l�;�6�S������˸d�x��i��6��bI�'�ኴ�F��B�y��GP�]i7�[�5֌�b�X���p��uy�&�1Up�7�O������>S,��p�A��o9I;{��8�m#Ϲ1b*�8�+�vkJ
�zDӯ`��n� 5f&�\��/�\��h����/p������=�[���b٬�%(k�V
��c�Z\�X�Q�JT�#]���8	m}���7i`�v���)�')�o�W>��kI���Z��U�f��n������{M*6�d`����gz+Õ(	�J�]hn�'�'E��Vep�PE���v���h��ƫ&�k�������Q�P�&�Z��X;q�;U��8�A��u���#��:�W�y�;�*7nc�S��V�E��k��5iͧ{ѓ �sx��+q�p��:�y���>�VbO7�<U�7���&���xi�.�t�|ۮ��9����Z�����Pq�4]D�CR�I�ã�zMЅ���hq4�t�ev��X�Jh���MS0��
�q�Z�Tٌa�s���PYRc��_�� 0�+glў���s���7�wC��׵���k��DFht�u;j�٢��c�Fa�`�j�������e]Yz��pnRS6*05R���멌��8_o[ɜB-��������e�p1�C|nZ��#2���и���ҏA���؟]�[Z��q��]���+�����3���K�-��]R�ҝ�zeo3t��ڛ���1ܗ�5a�5�D�Ի6�v4n8����P}�v�ȶ R� t�X�&�z�#�r�H��� �-*�ŏ��\eV6V�
%g�7P|I�C��tn�s3e����Dl�i���Y�+/n5�:Uʷt��`�y֥n������2��#l`�eS+�ʀ�]���vE�=U�:gB�]��/k92dQ��ʚ�dG��uhY%�[e��6�؈-�H<i۱!�P�u�-P�m�]9Ǖ�gQ��pK�l��p��v/Q��o�;V �sU���R�ǆ����5�+��)�Ҿ��]�Nh��+�I�j�r�v��ΰ��L�}���<�]����^�/"��]ZU$�&�e�=�eG7)bt�_G/"�����g]�� �b��]"�̷�.�^��!���&[��i��-�\�P�ޔ�/-tJ	�BԐ򺞺!pT" Hj%P�m�ro�`�/��h5[j��i���KCUV�UP[d��f���j"o#M'�������_5A�ĔAPEɊj*b�j���ͩ�*&*	�������|mT��E3ETEDAE4QV���ͨ���bx��>>>�U3�h(������Ә������h4b(���3�������.c���""���TgcT�6� �j�&�uU���U͉�M1:�4T��5S�L�QS[m�lh���X�l4UQ<�4͢ɣZ�ө*���֪�j�
v��j#Zf���:5QQ4Q���h����*4mV#lñ����j�JH��bӤ� &���bֈ�(����*��K�(�*�К*-���TPkE�PPS1�F��TU)�t��C��Prb(����Z�C�5��剂��~O5�(
?!��
d��k��֦��ݙ�Qg�m���'�-�V�O�wcص��esIӝ]1g8M��*�t�\����U�� �z�%U �E��Ƞ����JfD	�BeBHhE�Pf9�w��3L�O��N>��R��}�_�E��@؇��}�2�*��s���v�P��r�+qW�U5`����g��y�Gמ�jD1��M-�ۀ���qx|z��L�x㼚\�:��t[k���t���F����7�4���ބh��X�	�&C�n�L�v��;&rY�uC_^u��p�cɹ=�I���smx�Z��9�j>x�䂟������me{L��Q�ʷ�_ �R�U�x�؋*y<�y�����R/�27Hݟ�By�@��؃�����',��pk�j�D7��y�~��G��өT��6�ܲ(-#�v�6�-O.�Yp�H����=�H<�^j��G-3
�w�M��y?g�Ihʵ^f�fu�b��v�8�&w�Z�>�%r;H��|�,p�jj�Jyc�,���+�oӱ�R�3|j�WO��l�T� ���r��k�6M��HF�X���eQ4��_H�Ԥp�K3��s%��W��Y��ӫG���|��C�S�z��5�B��;AhicZYQu-+�RU�yzs=9y�6M����ftH�e�x`j��;��Nz%۹mֽ���|y}��iS��>Nf�ONՈ1.�:����b�ϰ-v���1=���p���y�1#,m��]v�S/죫�{!���4��H���y�sU�8�{tVv��������f	�b�
&ZYP)�P�T������~�o���|%3_���V!�q�L�e���$`�T��|[؅ʱBVa&]����[\��X����9uc�HU�(*�������xӴQ�H7�غ�C���={���\�U譻�*.w�x�#]��x� �����T.m�45Ez|/L�x��&n{�	�S�V�oS0�U�.]�.��f%]�.l�.��JusUJ΁��I��"qz����O��MK"Y6�9���ec�d��mk��\M���=bb�6/-�ֻb�f�;�>l��#��%���C�����a��j�@?ń�F8�i��1o�_�����dSa*o�U��ϯ!�]�?�{jT�m{ ��2����vvfu5�	N�
�4iŃ&V�OI�b�Xnm�ͬ����e�h�SC��]�����O�D'q>���Xl�U�^�j;o<�9������|�	��d���<r�ڿmܙ�)�^hs����S�Z�=�?B�xǓ:}��F�:,��nV�����f,���	�G&�ba��A��v�/Ip*ȓ.�?B}�D<��u"y�	l�L�ʄҟ�FN:y��7� �}�����/�@|�of��W�+�uBL.[{�!�P3{E�p{�J�GRu�]����E�*FFW����˩�*���-��)\����eΦ�oɽ�w�'R�C�8M��"X����6�8dsy�
GR�i�S:�w@_V��:s�i�'�pM�������Hd&fR�I�h�Z@��V�IaB�Sϯ~�x���}_{�>�E;�^ؿ>C7�"(4?�̼��1^����6���8Ȫf
�Þ�:auc5������|��y�L�#mx��J��4�*
�Zf��F9p�!�w��SQ�<��1R�-u:�nx�41�t�m�޸1���v��M2�'�ɮzk*��9���hc��ͬ�ܐ�^�ǒ�oq�Z�������v���p���s�R��L�gN�(�b�+d@Y�����6%�>ЊkҸ�t��F��ˏ��ؤ���cY[l��q<��O$nQ�ۃ�''�q�֗_��uG5�~=��q����h�r�����xr�mGۥ�2�sˡ�*P���Nlf�9��꟏`[U3�s`�"~T�/~=e����<�[�+P��:7ysX���e�j�{ZR��@%6��w�"���)i?�����ҏ���rA��y`c.�%��b�{lj,�okk���;sը��`�+m�Պ�!�\{+����_@%;֚�����뺻ri�^����k�:e�AdR}���M�ݕ�,(n�2�8��+_�L�>��2�ݬ�y2ӚgC�tsyWt,�8�SmٖOol8��2ɞ�R�+:+^[N��c��	��X�J��0`u�=!�ŭ}LS����}�pXī��|w�u�����A�(�����:]���f=i���Q����?>}ow>O���{�ߟ�O���Uf �Fd ��i(Ef����7�������V�խ�䳉��f�+g5F�W5��~Q���+�Ӄ5�n�wk(��k�N����r�=p�JCO,c٭Rg�+�cA`{X&�A��钝bx�<�������o�S����zꐛU/��4�\=8ԆȞ�n��yO _ �¼MJb�GP�DGQ�HY�gZۋ΍&�
�k���W+ͺ9PB|r��8�*/�K�)��#����rñ���*�l�\���������u� ���:��K�D�*�Xgm~ia1z���2�L�>����0�(g#b���&q�6`��ύ`�,'�V�j �@	�� ��{.e��Z��F��x��~B��tt���'����b��aS30/]�F�k���8��Na���7�-�4�C���#��P��I՛�i�7�,3͏fy�^@5R[���j�97{�gM��g	دkդM��v�UB<������+��cciM���ҳY׍��=�=��$�t��g���1�V�@o��9���'�Q��`#hUSE}��6S�'Fw�����K�v���
�6��5	��>�م��}]�ZT���R�[BhV�c����M�[Z���/#T.��BӱEj1+��lD��j���s�:k��s��2�����!)��P��^�v�1Q��W+o�ikڵ��b���	0���(̨�ЩB�$��ߋ������ܗ��5��-������$`J)����FCV�[�pi������IZT��~�g�z���!��k�(p'�
��gY��H��ʱ�950��; [�Q�[��a5���7�Fg���m��:�	�EL�y��kk9	Mjc�d�%e��μ�T1eD<�zw�G.����s��'����I���~(����݉�nu�;��~��L��ַ����z>{���ƶ~�f{=����֌X�$0�b�޺���k��¯w>o���vl���X�b��;_o�g�w�����LH�5������Ir�#3q�T1�hvC�Ϋ4�g:ǈn)m�v�>�W����d�6P9=��L�d���`��z��.9t�鑾���2�?i�͙u����d��TS∤��<7#�:�Ƶ��
l|��f�8�AkZF���6p=0�X	���&��ۛ\��rD�K�(��,�(����IA�,"l��#���)�7�X��BY^#[|w=�����>>��29J
}m9�0[�v�T$�J/c��f`��$�����v�YfM�����9�{*f>A����V� 5�\�:W|�7R�i��[W��[�s�rw���Q�n*�EdN�k�7� %�1�6�����жDd]�J7Se+����bV,r^ǹ����^w��}U�����0B��D�P�^��^����o��(4�!�΋���t�/-�#gz��v�V��ڥ>�u��au�'����ɧ�/���5܁��Xv>lYaf�Pm���*� R�Q�9"���l��7\1�O+r�1Y�;$\R�Z�j1���(G�~ݖR�C,���L���%��b`s�R)]���]Qs����˼-�(:dMC�/��z����N��k�(��5��4�Ǟ��	�:��e�V:KT�����uzN�����įgf���[.�ແ��[4O	$6�%� .YJf�AK�%,�ٍ==>�zx]�׶S�K��c,�Mws0�7yS�QR����˰�\�%�͞7.���E̽���5�=�~�ټA}�<(?.�Sa��/�8�ת��'��3c�*暃���w�;��s��17;me[>\��/ɼ򖝪�ʒ`v�*1'��w5#�ܡV��B��{w���]��w5ɶ�mSm���v=��a��?(�ms�ۑ�"'��ӄ�-l�Lm륞j*�+�`�6�"�q�4��r�W�<��QIͅp$��G�{�oE�V�鿅����2�W��޽KFQ3깥g��,c�^��BV=*ap�<BYz�j�N���7�J߽&t��|;��1A�G��gf�tR��G��|+]����Ƥ8>԰�ֹ�^Gh�ֲr�Ot�t�qܝv�.✏.�B���9�y�{��Q?) �*̃H��	J��>w��p���l!��s�ҩk�J-99�����5�s���h��b�l__c7�ʼ�wVݝ��3��ωc�<�;N�TZØ��(�/��P<��m��E����?m^F�}"uy������76S�&�]��>��R�M�.����=�ʃ��wε�`"�g!e���숧B�CI0V�>[q_��S�S
9f�_�N)�bg�6T�1�)�j���3Ƅc�;;zf�����?p��WƟ�B^���H�V������je��V%N<���d�]�b|��5W5z�Ev]������u��۱���^+�4�>n�`���4u��?BZ���PS[Yk�.ˢz{�"S�V�6c�\�p$h[U�@���}���~�A�I5�cH��oVC�R��ru�akV�-�\�60��V+����<m���@��qNlK�P��I3so����˛x�\�)a�5x@\{dU�7����Y�Ie��R��Y�i\��6�.b�f�O�0V.�*����l�d@p�s���UT#v�@)|wy�6��+�щ�ȿLg�ށ67��1m7�]~R~G>��`�2 i��:�鋕N��w��>�{ذ+�p]��R��/��4m2q�F�k/6���]:<�e'S�����α��o�&�v!\��w�%nv���AgEI��^=�8����x��V-���1����T��;��}�WWv��\_�U_�L�LP)04 ����C@�4����߯�z}����������zW/�4^�To�W)���v^�Ԋ��g���b>�&����ߺ�c�u�p�;�w@�S}I@Ώ4̎�|r��1R*�,���y¶T�q��U�j�������]���X(`������2��򞽚Vخ�6�[F,���we��<�m��8.X��75���+�i2�����6r�'ƌ�>=�¸��{�}�3�R��cV�0��vժ��sUUN��Ιy6�^;��P�-�4z������锟s�O�61[5����[y!��;�"���n|[؅���$��	r''�Z����4�	j�6U�=�����t�۫Ɓ�/剬���gn������_C�N>Ց�ĊT}�\{��s���)��d�z�)�؟��6?2�������r�s��N�Xk;��	}ЋJ�Z�M����q�S�(��K'�6�,���J��;�BX*I�U�,q3�������iY�X�a!D�:9H��~h7Aj�5 �N_fZ�ٙ�4��UG�m�X3<]J�~[.�}F7\g(,;8L+S��+ \&��>�G�i�c�O�oo�B�k/&��� fѣqY��55z�C�9��竜��5-b�k�xs�tv�⦁�,R'�P��B����	Qب��D�&�R�,1��M�e�wTI �,�Ǜ��ԏB��-���pD�L�꜌��sӝ��s_V�&�9��G�"L�3B�ȔP*�H�K�2���d��Z����^�b�N��ORoW�:�n��f�X����[gk���o[�ѬO��_Np����>�����(:����g����tYTQdz{e���T�K?���7(-�8���_�r�F�.+�}jѨ9�Z�<��NW�]6q!��vw{Z�F#�_eF_<���?�"�u}:eo��ӎ
����k����&&�y{�FԕA�.�5��+�Ww��|Oz߱-^�r8�$qU�/�`ͳ���}t�%��/4�iP)�̬�7.�'�v5���������ޝ���y�9#x@���$�K"25�3Q����u+S��5�"���I^[)�F:b$��6}�f���t7#{�&���]�m���}.M�_�=B�N�^$���O�x�)��S��I2��>��L��ַ�r�dm.�9t�d��#s�����;Q>��u�^w�Q�R|a��=A~끲�D�۳2�f��g40*�s��7E�co��6O��t���?T1TTr���{�T1ǱH�AOm��<~�_��F?T�-v%~�ϱt{�E����S���ȻZԛ�,�4���]?^!4dBw�I�Kq���dv'ոGa�ذ�u�j���2A]&�J�X���MRx��׵�m�f*�N٘�x�8�f�����D����dm�=m�χ�>�{�0���ȓ#H�'�߯��������o)����%?0:�Sw)��
����r<j�C�B^2�#f@���bk�ݤ�R\w*mЖB�u�RK��U���nw�zj1���v��G0�@X�䂟�R���9��K�o�"w���_��ȖV���ɉo4Ur{�%���Gi{_�,{>\��V����}=s�7�{�l�<<8��6a<"o���&�WIjju+��q�ɄߝG7-�N[V�����b���\Gg[��c���5p���-�r�L���6d\^O�g;�{��;�S�-A��6���拾F�1�5!�3F��������'5�&�jd���i�{6����=������G�/V�a�8�[OX��j�~܏e�����[1?@�꒖�hG$mJǤ@j�X�F��Q������f�v�_T�����t����qϒ�L�Vԯ���Ɲ�@ZH�MX<��s�u7�r6H��y�7M��;+	q�衛ګv���-�n��g �����n�={�]��6�X^����������&ؾ�2K�����uQ��l����W�l-�3�J@�Ã�[-�>8}(Ū��S#	.�ҹ[9�y�' ��Y��N���LM�2�#xЮ�ʇ>��=R�� �/�n�\S�dX�۽0-�W���i	]�F8���#�T�ӏ����ݹ!miR.WKW��U�d-]sm�na�n�&Mc�(��9h�Yw	x8�̗æQ3�(=Rܘ�m�UdM�!RY�H�t�F�^�)J	���.ڡ�v���W\x��(�o��*�ؔxl�������6�7��V{D�� �����M�$KC�^a4�8�b�k2��nSR�]5�j	�L�
}.��0Xk�Ő2��Ir�P�����om������07NJ}�K�ZV����8]uo9zU�e�e�}���d�8	.�KF�[�j��+�!��j��.
���^�A��ʥE&�f��Nb�4h���D�m\ӹ���lz�x�9�{2D :��[Y�� �3ܲ�O�`+�.M�웹D3�&'��D�Um��2��{z[w��wR��j��B'H��,���|B�Bi뮄�&�t��2�N�I5Ҭj%���J�|LI��.�	G�`:�v�x�,9�˖��OyV,�V����DzQF��\۳��t'�ǂ*��%`5#쇨�,W�*8(mn��U:gPwBm��X)��G���K�4E�� =pźiW@S�>�.]����dB7��f՜�6!�j�j)���g{�knP�۵³2�{qe�C����m�˴�,P�8o_,�j�fEQ����+$|Mj�u�q�@��ҵ?$�-<��ok��#\Er�r�P������IQ�[ݻ�0[4J��/�U�os'E�(&3���r��5�J�IyMt�=y�(-�[����f���|孻j���ξa5F����'��4�vFsu�YU�`ʾ	�u���9��l ���Zsr����&�� �dek�s]�c���8Nvu�b�R�ﳩq�h�ވ#}[�&�ֹj�^�C��I.k=HTx�Q�S�4�4mˡs��72�@�@t�8%e�R�SqQ�iA�o^�̙���Q�.�vqr�.5x�T)w5�q}��y�㖲�CV�ܺʺ�0h�����P4�z{s�pl7��4��j6Ҙ���R�X��W�'�"c���iJ�un;D�.���Bwq�)T��Y5����o3�Xmp1��j�#P�RV���V^�����65�:H2�n�@�ô�*�`]f�4iKM"�&D�1�lm��T�����ZDԖ֫��X4�5գe�o.2WS}O�����6m��������iw`Yƥ�V� �*��:N J�Lڜ��r�0k��j���������}v�����S�Y��3-,���mIxh��� ����g%�?�[���;��ZW�yk�e��� �����;�Y����GW��=��+*J}�n�@�X�������:���"�}�C�*������(����tQAQ5E��ͪ����֖�s�~Ϗ���PiE@���\�.���f��]-%:LMC9�||||O �t#4���4U�#�IT��)l:����������<�ъH�lU��:��N��(�)���)v��S�ATP��x������a���j+��+cT���i��� �(����LST���nm�RDДPkA\Պ&��"F&��I�9�*�hY��I@m��5M��F�W$ܬ�t�R�F4X�-�FܹDCU�9̜�M9��F����
6�4I��DT���gmZ�U�j�-�sp�KgT�Ӊ[j(����t*�:�
Ji*�y:I���4EkAZj΢�-}�c2�	#��V\�ʿ�WI����״�+�:D�X�ࠣ��;�����>�w|y�������?(}���Bd	� �
)�����o�O���\�����s���g@�Z�?N/u�J�h��w��E�k<�9�:�%�ߗ'/�v��`7��vvuJ"+_�q�R�)k1�ʑo�%���-U�<αҽ-8D��YS��ګ�G�T����}x�u���S�����L���/A�@�����sP�&���(���TOE{�&���'�P���C�R~N��?�E4����3�c6Ѫ�X��_�d���{�6�Y.�n�{�s'CCJv�`��v�XP{2yŀ�e����������5��������Ũ�6���~zӬ	�"0C��}Y�ZH�(�ו�����s��_���H��dw8�j6�^d�^|�[� �hE	�&t4�ɧ��.�yʩ��"�3�p�h�g�u[2�55�um\D�i^Kv�X����d#���+12�f���Q��$�k�]��d�Y����Uk�Z��\�΂FS-m_�9J�$����/����<�#$��?xuh�!r�`�O鿮J~��󑢞eCJ��l��	�ֶ|�@\�u��Ҹ��aaZ�--�C��?!��i���v`���tٙ���.��õ�� ٳ���'�\���W0�k��@�fl���IW'x�_i����>�;��C��DE���`#ZB�����n����]or��-b�D\|��{Mtcb��a��z�=i��� L!0$­-$����:���hDL}�I�%`3�����gݐ�ى�;��Z�j �iG���k��y6���]|.qo;��|�ơ!�����V9����/n��y�ш��X���lj����׫f���� z!T��[/����G��A�Gv�}û3u��ށ2́�,&ִ�Z/�&�oCL������ߠ ?h�,�t�dC�㜽A}�ꪔ`]�҆X۩�"�ױk��B�� ���X�ѧ�{��_�E����Tw)�4��S�SuZ��Q��D�V^:'��jw�r5�f�p7�W��ty%mǚga*G"=q�*EP��Y�iD%�����M#���u;��4�[�� ����J���DI�����d�����{ ���#[�Tn�e.�_pZ�)�u�*�����-r�'�[�/x��q{p�
�!��)]��-vƤ�֚1��4���PH�Ic�裦EE�zO�'��W���J��b���YF���NN�xx���ɚ�OG��ڛ�F�iy�YЩL-��H#<�0�f�Py���%:�l���(s��[�od���Y�.̜�*s�uΑ��j8�����ݿo
�ВՅ�k�8�9ޝ�h��Q>�z]���6��6���iX(�Y,��,�щ����C��_%�N��D�ĺ��X�k)�5 ��U�����%\�Ev�1$=,D�N��X��b������+�>4����	�a�dߟ�<����߷����oB����M���:�l�0K� 
��=�c�=1xZ�P.�d*�2�Zo�+��v���/j�M���L�?O6�>�-��ҏ���G�x&����(Cp����d����g��]�o_pJzu���*�q@��-�tk1C[�H�l'�B�����Wco�5�0�c����2���L�'7�>S�hU*�8��ԧ���xGW �t�o�9��įzh(�+��]J�F*H$�u�|"bۨ����-��WmčF���Y���ɳ5�ts�y'�*|<#Yt����mJ�8��g�;Y=8t-~�L�\�^Z�+��_u6h=�=�3NHh�}�|�tC�cXnߵ2��U�L7V��ں[�I�ɵ�{N����v��(Q#K=��c4TZ��Y�reZ�o�f�|�Pq缺�hl������U����O|*�3��Ih7f�7��{\��2���pi��GųܘY�ɹ՗��R۸MF�E�F2���4}�-;kyp5���h�IޖD}�0��[��l��E���X���2]�e���P:��<n�wEpm�[�k�v��]ގ<��ǫ�g�%�=Ʒ;��Lk	ǱIB3�Y�;��J\�t�}�Ӛ� ��f*��[����k"<�n$�G�m<��!0���������_�?�$�0B���:{T�Ji�;o����P��ֆ�b�i��{u]75�H��jl�%t+U�=��3GzO&G�\W3فYo��l�b��:���M"�Š�x�9Cr:���wA�r!�����y�qf�������J���E֝��_��(1���?t�u����"�pW`�]�K�1��d���A�T2.p�X�ySl#y�!��5�r�{�O�S,q�Vtmݢ*rbO\*��ۺ�%ք�#)p\L,�Swg��m��G�����y�Ȳ�����-7Q6����d�$LD]�jAv��9�Z2DpmҬO�"�a�c�}ϩa��㰥�N���Q<���e�a�����G���8�k�0��dK)�%����J�^%���-_/�Vo�Jq��r)�f맰���c"�X�H!q���9& �}�?t��:���6P*9�\H~�U��]�U�]��薹r�	��ł�d�/�|���Y��/'��Ό��!	Pޛ#EEV���+xKR-%:f�ޚ�r~�AðXY�!�d/�A�ό�?�{|���qK܍����[߶ 3�蘱����N��^�5?h���	.k|���A7{�0�G���5{O s���[�G�ئ�F����>�x�rv%�)�\`e.Hܻ:��c��ڴ�BR�^�u��0h��ƚw+hد�g����
�����o0f����8��ؓuD!��NkG�K�n0��O��砥ft#ka�nAa"p��i��q�o�;e����Uȟ����o�o�;K����^����̟~W@�
uZ��Р2���^I8�̹����q�ZNl�P��_��6�
��p��ۗ�Yᩍ7���� ��.^�^.{��yJW����ܢr��JO"���P�|��|�8�{eV��
�wdBnl���ݭ��,��������f��Z�VK`�p]�s1Ƥ���Z���0�r���zG��ew8��{��*ʩ��:n7�����]�,��&vz&��s���i'��au�Wߥe��dp
y�t*Lw��yM{��O;f����tT���^6�+*�ߒ�ֻ���xi���VL�z]cK�"g��~���ͭ��Y���K����{�tRu���?�)��*o��!��]�O{�}����K��l��7~�S�����G$
|�ao�M8ޓ+\��珵P������{� ���y�o틿b�6����+ZG��a��3`��gi�J�^���E��W~�xY=��*�n��J�pD��j��O`�w:}���6�i1�=��5G4���<8�8�Suk ,�}R��u��2��͑JLm<��d��no6�{��|����y(��-J����.,n��_\���:Kb�9ǫ��&�߹���������b��ߨ�������Hͫ�w���>��7���4F8T%�sЗ!�O̚}w�N��1�r����8��dŏ��S�]��ύomH܆1$�VE�]p6D'��K�~7R'�Gb�M�Ҟ��M���'/�3W`��N�_MAi�I,���c��B%*�t�7�����ڦb�Q��t�7AήD��L-��="��J��xo���>�8��B��4#k`7d��ǥM�pO�b�ݝ9x�Gd�<!
�>�Ǵ��\lM�3���H�ơk�>���[��Zw _uVN��.�����V~�A"@�Z�a�w�6QO�l������5s�?^�b�JI3pV5j�j�����"�{}�|w��61�����]߫��˿b)碏6�ͽ���~��d��a6��U�[��O�Ru�DGE���U��UT#7�Ѧ���-8R�s[�R<��j6�y&�f����B3n�<ڏ���s��}+.����f��l�霘t�_��ջ�&�ݔ��f��z�2���B0T�G�P3��3+�����������M��K�E�[X���i�T��ph�����w�sZT�J���EH~;��$�������2N����|�YN@��^Q�	��o������׿b=N�bxh1�:̯j����{+���DJ*9m�۲�-�����
�6Z�u�MM��5e-b�%Rt��xUxX�8�����́?
�op�÷�c޺�е�l��[c�c
jLCϺ��u�x*�/�r�u^�ݷM��|V�� O���}�*����>�|{����u܏^�z���Y�ur�{��|ȻH�q���	���;�<��󳆝�N�ϸ��N�Dm�����[^P�~Wr
�.�H3@/1[�RgA��P4�`���F�6G���bz���:���+�ɁL��S����&nFT�?6[�x�iS˞�b��[��DƸ��X([��Z뾾'�uH���
S	�r��28Ӟ�Ԃ�e��9�R��'�#V�]9��״�n-5w�(SN���/��N{�ga���6;#�'�1�fUը�E�c�}t�>R&�#���A��-3�)��{�ݜl]��K���P��j;�aPXp�*_\��^m������b���n���^��A'�b�C�[�rz>˞�}ޏ9]#�=_��S�6"YVێ�n�:y�`�K��A�(R�`!k��@v}����r: ë_�	�aLJӆ�Y˹��9F�y�Y�\v�i=QC��� n�9x�It������ׁ�������u�R/Z�m�Mץ����9LU$�\�n!=��zȖjzum��)9�w���ElÌa�ݍi,�wң���uΝ�|��G�5�ڳOp!�b�}�͕������-�C-R� ٘�vCGhcިh�k����S�=EQ��Z����(�=���6�Y�b�p#�VjN��N��o��ؙV�b=��dD�S������-uGx��W�y�c����UB0.��X�5���xg�SlB3l���ց-�ږ1���6��g��N���q�n0�{���w�mz�<��!�BD�{Uc�~U0��r�z\�mQ�������pN��S�Y����CL�ps»�M�
���jBm���c��������y�Sr�~K��� 6�T�F��;�O�C%z<�3�V)�?B�j�R��5��Rt�FD��on��xGk���],�1N���Y���?kH�C�����7D���߮���+i��6"��Fb㲩k�ۈ��8��+\e�/W00^_�E�,-��1�j��G��`�N�7����uv�Crr&nt�S�Bt���۫�U����=���u�P]����k���צ�e�]ݷ|��M�1ŉ��9�ڄ��\_<b���&��	J�ֹJC�����A^u�ڈ&���٭�3,¸�WΦAK����q�zhm�s���2*ww�]eoh�����tAM�r�;�ZF��2���g.��ECX��؞�'9�Y�rt��J�V�Z�Ve�ܓGJˊW[���B�"K�	����m,�ayǂ]��62��6c���w�����g�9�Y S����_Vn� ���{ �u#���"枦�^#��omL�x�k><-RI�q��[hs+Is�ou̶�ʢ��%SN��:��(LC�)i��&����n��v��EC���ǵP�;�?.��e��#,hu�zX� �y2Q��r/sB�꾅\���L�4��f�̀gt�#����ز�̀��"�.��\Ķ�����t/sb{�!e:;J�k��:����[г�6(�W�pR�?e�Xo]�)�z~�4+Nc�Z�t�k.�H���1�J�C��̍l:��+��'툝R��D}l�f_�w%��L�S�R`C�^�1A�7�ϋ1Q�D!]��5b����(�1��4H�>�%Õ'���*g^L�v�!��ғ�>�LE�3�.�N�ׅG�j�!�w�(��z8���,�W�:�Ѵ�X�Ĺ&~�)HS�}�c��K��Ǹ��%��b��t����6��m��VT�uS�:�֡M��p}�_T�+���1J^�?5G�<�1>���j�o9������վ됕|^т_V�ڈǙ�ٻ�s�/���Y5GRP��g��%	WL{��ǚD��e��!��̣}k�O8:��1
t+4���vQ.�jItsfN��k�DtWWoU�� ����>K%+��wmsk����X�;V�e�s���VI%�;`���ġ�7Uwo;}m�#��uϵ��LGS������U�;�5ΚfG�9�^>���aj�*���V+�ݾ-l�]ڐ������蕏>���#6�k�e��
�>`Q���������I�=C�[���m������e)Kǣ���}}f5�Z��5�M-|��8�-�H��հW~c�?K��LG������y�����v�D?���@z�+�<%�d�FFwF�[q� �'ݝ����8{c;uM�rޖ@w]��GzY�NQn���SA��	̄`]gLn��u34�o�;.�z�_u�L-��������V��
jH"���"��B�
9f�_�N$��aӹ-�v�^wk��)�^�4�.[�[z�-���)T㤑���C"���w��8�kvf^kv�nvI�z�B���"�R�b����kg�tMsw���ix�z`�X�#ΰϪ�y����3�j�	���c�y�ja���1�N2�]C����WU�^J03��S��U�Z�DNC��v8�|	�jF퍏�A�9���2;U��;�:�^2��q�t��2�,�Rw��?ڷ����
�C����y	���*�rcٺDJx�������i�-|5�����ޑ��хNa�5_K�r쉲��&X��B[��\����b�.���Q}�l~��cs����Ӌ�}y��$�r.x��z��8��Q��Z��a}2�վY�����چMT+˟��}4gd�s���*L{/o���w;j�OV��\z�Xc��ehń^���4��BbS��N'7oC�6�w��J�z��d�z/�۴����q��E�b�ȝ^���jR�C��f�<���f�hf�H�J���
��K9�3�3����ޤ�+����[%@�μ�"�hKV��1�v��]Λ���r�2��;L����D�ڼ�W�{�Փ3Io,�5��N��勓)5wu����Y9}]��C����� �vtZ��}�0�f��7��h�ҐKJ�<t��	q��l`؅dꄎz}:��5q7Jcz��36�>z�7]�#���$�fW1�u�|�E�X��:��=�Or��#��c6e�	}��q%`ה@�c�IC���<Q�0�].2�C�κ��Υ�o++`.3���qX�� �<9���"���fT��նY5�k�l��'1;�/�-Ι�Sj�TvP��_�F71\'!P͛���{Zꃐ4�
����w��;�����:Ȥ�T۲��d{�Z4�^0�^n`"ُ�ق�4r�9�Z��Z�5t@�=�/��Uep�hr!͂�#L�a���^��+BQ
�,hJ:o�i�Y»�+iB�}8�(�l��7�㙯��1�����x��
͍���o�`A���D��@i��8�\��%A�#׬V�
�F�o��m�W2���nBٽ�y1]�gL2T%S��X[�`}6JRkU�'�i�ج��Bg><�[��7fD&�6yqaq��iw2>o]���'v���t��	��0��gs�J*�II�kl���l⫮y�U�E�w��b��I�f&�V��Wt�OSf�.����dYF;��]Β�[�y�W�-��.ow��ܮ�*�����2�wU���w��V�9_E�c��ͨ��V���֮�*�iJ4"+'f.&��z�|-�*l��H^d=����7�ʻh7b��T��9�.�i58�-�]�!��++YVY�\i�(�쩹A(U,���)B�<��ѥ	��1�ô�l���m�;�^E����g��u{���O:�c�L���Hr��=���t)R�J����,I�wg��*�){�j��|�G��	Ҥ��T���lgv�5��[��s�:嬤�Υ:1��o7M����]�q��׋��s3���\�;����N1�F-mr��V��S��:\�.�}�Zb�|㢋zkr�R�Oxis���؍cm(-A�]=[�n�x�V�@L�H�ս��@N��Uh���Sp}s�j�
nذX$G��5��;pAdX�@��X��?��J�M%�11U%D�3�L�"����,j
��6'>������1m�E�����ES%A��kHj��4QAS5�b6��-Ȉ�� �x������Tm����8(��QElj����bh��cAڢѧX���������N(��k:�������Q��m��Z�����J�55kPS�������S��F���PPh�l�J*����KcTK��M���ՌAZE��th���Ѧ�����KF ��'IXv]EQkD�UDU��lD�S5b6�4��M2PT�1TES��Ȳh�-bƱ��b��4Alb"gX��,DEG1�j�A��`�)���Zj�4U��.�Y�LG�5͚�j���"���V�i���`�f	��*���Q|X�:b*"��& ��"�J*��	��Z�F��   �w���"3
V���PÓ%^����.�ۧ[M�z�v���+s�r�ԯ%�+kz��g�x�V�����mD�x�S,SQ}^��}.!�̗@M�a5�UG��<|;�EP��l���\�S��zF�y1?]��efͥ�}�{�=E�L^�R��>�ip΂p�7Ѧ@Z�W)�+�"�*� J�a"&-�=�OzY�ޕ�Rj��4�����	�	��W�ޘEv9K�|k_����Q���itO��.o�]]ۗ��-�"3:�ƺa� ��O۝4��r�>-R����F*�l]A+F�^ g-�P�|5Ш�{S���^��P�g����'yM��ê�uJ2�8���I`���
x�oI�(������\�)�{�TŜ�i�?gBd���'�v���AN�G>e�y=�U�Dg��/�m�" �4{$��Y]��yi,L�����2p�ώ�����!d�ѻ�[3���3���Ū�z�(�e��������m��
�ǆ!�[�h8=����R7Yf".�{�M��˹׃�"�i⛵�>��v6����}�yJn��=��1M>�a�gW�N��̛������ڳ\� f�9�u��Ys�z.�WʹM
��0�����%w��Ѳ�i��3��l]܍7
�&����N�0�Y���XE�1ߵNT��Nݵ�K��wH��`L}��`63��WS|�[K��_����5��
���!{dxA�(ҥC�O�aY�iR�����&'�P��kJ���s�l���!JF�����J�+����K�i�Ϧ�/X�B��+�ɗ,ڮ`Q�˗�s
;S��g�|�p_{2�m�g�������
~kS�Z�3��T{�����U)q���ը��@�Iab�{)���d�e�-ç�C�f������7������e�'�>�Q��	:�n%&2��vS#�U��зJ���Fo�us`&�����!g�C�'���=8M��A{p�N�W^^,��yl��FWn�jvf4�H�v��	�Q�G�v��:�|���N'��,v���ӽ]04��C�r�jb���b�ޘ�Ao���1�V�/��a�阻�1}yyuok�����u�|űI,�7��A��}W;�iQ���4�6Ξ�:a�У8㓻j}˴���o��||��_c�]R�97s����JPn�R'5M�����������U��f�Ads#��h�]!84⦸�V��q�O ]շW��kj��MjBmAt�X��/3�_�1������cM7�g��xY8%{���c��߮����?�s�8h%��O߭�k~$�ˊ ;IQT%�p+ˀ]�m<ۗ��;�K~:��mnV�&�ꗴ��b�48�����u���g{���n�Kb��ޭ^�q��n�*io��ᦡbMy�y�ϯWЈ�Ty�]䭗6�P;}ݦ9����b��٦=x�[��fJ��Θ0��w�'0���xT�*�nS٫A7U1�2Y��nm�f�C��Mb,*e�~>]6�K.����`U��7�|?"-�C��i^��d;���Þ�<�]�~ۀ�y=��C�"usT�'*�:����r\N�=��6�""�o�7�USFΈ���!ƪ�h=q�qA�*��b)?5�tsm%+_��c@K��gW2�����nsZ�w�H��@m�"5�^(�s��{9�z7zs��Dsj�yC�ض$�r��i�d���B�X�tp���Y�.[hk+�D&��e�6��"Z@�ļ�ٔu�fa��Ufge䞶�;:	}n��O�hT�d���LX'�����^����Ɨot�y�Zg����Kd4�M�c����L��͙����@�,yCE�q����ؘj�z����v��M:Ǥ���sw�N���]�*G���=�,20#h�j�z����|� ׯ������}^c�u�EK���4�l��E�^܁q���Q�Su�fo�"O2s�V'NΕ}��������/Iux\���(��o"(�\W�]�+K���:�u�M�}i˭�B��$[4�Ű��ABU֋B���5�n�a�o��v��z���Zٜ��YpC��v)���5>�nt��̫��nceʍ��XC�v���A�7��.`9v���_y����fF�<�h��˟��ٕ�'(���t@��Q�{lOj���V����%���ܾœ��(c�o�A��~�V;����cpO��dsS�7���"�X������,�4
2���E_�Gw[����"O�T��������a��2�^n�����E�z����|ڳ3{���_�g�)b�"�4�S�s�S��������R�V���L�@��1�V��g'������ofU۠i�{�x]���t2��My�k7�DȻ香�-sp%x���{x��O)48��Ay�˻e	�v?<+~�t&\��'�K�[m��z�8�ƛn�ĭ��]R3���֝������F���,��DB���<�:z���F*��2�An�9���#��%Cd/}
E��ʐGi>��z�,���X��%�W�8|�7��y�Z����1�:օ��Q�x�45����$�i�;)7H.]������G���B6�v+�b�]y�
���^e��f�,�'�xG;5=�~U�dY���\�b��6A��,ꮒU�K���+��&p�t,��:���8;}bc ���v��7Ww7R�=[�U{�!<��Z���o��f��^�tB�_-U��)�ҏ��\4�rU٭�[�lK9�c���*ݢ��
|��R[ӭ*���I ݱb?�V���C�w��G���
K:+6�f�#Ȓ�S�yVSo�/�˔Ɋ0y���zЊw��lvhw�̟X]\��F��+ų5ђN�gFƩ�B^m���=	�ݴh]��I��[<О�\�;��6��_Fi[Ӊ��t����G(��!�Mb� ��q�<�d^ȝ�:�n'F�5�4��NѪ�z���5-�NǏfu�*�'2�u��H�v�rMO�"`:��̟#^�C�A�v�/�����)K���@�:,-3\Ẅ ��b&� ��� ���Uq�d��]t��،*|2�6V��_e�w8����EN|h�g�O��>~�)�1e��µ�o��Oɫ�ǷWϩZJ��ԟ��z�s��F��C5Y8�庂�'{�vǒ�_�5�N9U09{v0��0��d(�~��՞��~����~�<;mRޝjF��nGl57����BCT��]4�<��bV.aN�gz��DG�7 �$]Dml
�/"��$��n:He~.�dt(��X'���l��Nr�*��ٗͬ����x�*�}�%(�����H�ĉB����ǭo[�Y��w�7m�=�ay���^�;�h�u�XçH`�<ֳp��:ic`�I_�����
Ic<�&�w6��k���U?;�ab� ��դ�v\���ʎf̜A�].ï�q\�Q��W,�,a�h��9��N�i7[6+����ѹۑ�����ފ�j1q�����xnY��� ���/�|�8�>��=����l!�j!�7`t�TNp�y�Ͳ�ё�Y�gc�x�z�[��2�r��z��w�20���R�]s�Lh7������bY���f^�2u����TS.~�
����Y�rf�b���Ϟ�2�0閼j��o�rQ�9}0�4ۡ��ً�=2�H&�7�*Su��m��k���(
��,��4i�wR��~�rݻ�����N��1��O�d9�1\���������`���3�$b�i׋v��Eꎚ���ʛzQ\��X>vza�A-|r�����6.Εj�_�cS�Q���L6��B
QU|�WN�׾X�Z/nY�V�ņVK�k�R"�
G��a��;U��{rE���]�3<6$�t ����fFk��H�h�ŕ�[��T�	�����d����֡p�h͜��Y��)��,������s>��M�v3�z��i����)���y9��>��q�YUQ�T��uW�S(�7c
��ʮ�X�|!��%��a#���|�]�3K&���u~wtw���ȊB𳎺�r��
�ds�Vn�#<���B.4��u2%���;P�H�jrnՒ�_a���vMR|�.��c]j��{*F�A[�'N��pV��n�|����sDw���oD�ήh���}�ͷg�x���5xNN���$��ET#,���-KO�����} �rW+zq�6st���F��f�R�$�����*%�i���*�d�7oN�#y�m�r1u��g���9sy<�(Ǉ4{~��:��{������ηjs;�M��?*�؈S��\7m���f��۞�V����k�{�nU>���\c¢�-��'E�SYõ;ng���� �sxN-J�pb�zo���<�@>|�ʙ���]Ջx�ͯ���)m�+�d����|�/H�x������N�dn؋�W�dmc���>l�'���%�<n�F�mCh�7O�Z�f�q���u�g6��x'Tz��;�4��y8��v�̰ɞ�k+i�z.�.,�9>��g�0�f8l
sV��r��J塕]f	q�r��^�'{�wO��qW��g�v�����Zճ��冷���������9���xʩ0f��j�rZ�7r��:��ٗz�����^|�\=�c:����Ӝ���%bf�L>4��j�ъ"�8"�A�;VsU/;<�*U���m�٪��=կ[�����/��`��Ě����e�{ׄ�$�j�s�2cQ�J�v��ik�� +�f��vM׶�̗T��#*0����&7XQ��nΛ�o����q�|^}V�YL�ä�vb��i�|W�}�57��Zg�G�f����{_�{ӏ��h�Q���>�8~yX���2�[m���L���+]��W�_��1�]�^{�ƽ�[��\���Fw��)����Ϫ B��zrC��M
���6���CM@B��ԩ�SͷW��*�@ϳ&��X��N3};gڛ�i�t�nf����7f�v�LR���Y�|y��V��:��<dy���,7Y2]�MM��Q\����v���*}{�?x�SՌT˕;��k �����j���o�˺��h�lSHI��d�r��>�g���R
�4�̋T��ګXH�v��}�9K���/v@g"dF-oO��g�X$��Y+k�e ��7�d/��%�k%c��i���UO�`T)wN$�j�vU�W�oUŸ�;=K�<���'�L�=�R�p\.�p�mT���.U�$��OO�����̝c޵X�{���N�i�E�rs�7O�F���Y���#2V��:��Wb62��p=��	�n��}��<M��n��x�y�ꦷ)��*��q���+�${������[�e��Y�܌�:���I6�x�|�ٖ��z�3Ҏ��_�9��j�~��sO�f���[؀[{�j�����=�g��C�yϘú�%�u�� Й����fy�����;�Ί6��!#��������z.^�b�����A�U{S����*���
�P{�c�hUy�u8gh�y秊����2���6�f}ˣ�oUWt"�s"%f]�N5�6œ�5~[���YMBz_�}@����U���-�Ed��� �Ra�d����h��}]��Nm=׎[�������m��}��*�FGj�.o+ޑR�{=����I�Ƌ|c�д��w��1��<}>��z�"��5�==5�;]Vw�^!-��\�̓���W�����Ŋ���`ʕ$�xh�)�����QL@�Gn[k���LZ�^�vE-�GǶ��ܪt�9@�� ��Z����ա��mI����a�C;^�X)V/�09v�X�܃��G�>Usk����5�v�r*˰QӽA<m䟪����x����i��Pv�38���F�-b
��Y^��!�IyN	�j��������l��숚Wu���/>�E� �oNV�fgJ��/1fy���S�u����ٛߑ�q���Y��1; bKk8��7���d����m���ѓL���ǆ�!U^WH���"��1�v�K���:�e*�Ѵng�ᓭ�y�z��w�QVؤ=�u\�}���Xo�▁�r'�����۪���w��[7Ul�Uq>�cB�g&Ʉ�2��e�ٞz��캛�@3�4�;���J��V��[*����UN�զ6�:�k�ws��Q�f��-��2�)�m��8��n:�J�5U���m+�]�˽,$4���m���*}j��f��+UYN9���f��fD��M)��.^�l�`�G�P���uN��j���J$+�'ޱć�ciҩ����xvr�fU��)�rq���d��؜�֬%udb�i�W��=z����wl��.kk��}�
���ɚ�aks��,:Q�ld��bp�;�*�u쬦��������)��2���J3K�9��ݳ@H����3!�{�DgeԶ��e�$�U��j}Wwuݩ��DѪ�_ig��E� T	��.EWEt�ǳ5���9M��JQR!�o%��E�����󧳇��C�7N���v�������5JWP���k���ۣ�LV��b�]��Sw/n:�@ҹY|���d·�o<�eK�H���}�b��e���.H��ә�2��VqX5s!Vt��\���ʬO��uw��t�$�����sB��o%���OL�gI^:U���nM
F.�@�ێ��m9����<!R+���u�G�q;x�gR�n]�r)�c��m��NP���;i�F��v9}�,�ߔy�5Z㈴��v"�0���h3Yѱ-NgVt�i��6�c�5��X���J���)����@�eK��P�oZy�*Tz$U�C.��P��xm����]&$��K��ӍD4>H������p��;{\�c��k�ȅ�!��������J��+(��F஧vt2�+�|T���k��Y���f;��-ܕ��]��gS�����@6ZΥ�Mku��35WTIr�K��!f�,� � ������Gf���2.�[�FAn�w/Kt����P��
�6��[2E}�キ<(�w�р�y�0����]Ђ����Y�Z�o�l��<���/k�J�R���Rb�.]%}&���Z�i���1����Q��7d�w^YN�1\p�㔬wVR��Ϯ7��q�ZJ��.����M��O��������-�'��Q,8�r�c#����X�+3�B-46n���⠣w]���V�̃u��r�u	1d`m:�R\/h66�xJ�v�ý{F���@eKdh�q�e�-�������UpY��(�[�"�k�W(��/v�,���e�{��]�.*�溹k7"�B�pᕎ���6�� �*�fo.�s]
\�O��aU��� �"���պ�#����fqIfғ�\Ď��K�gN%�G��ˬ��~o@�R��et�fw=��V���Gs�.���>O��C�V���4�/2jťg���o'���i�t�ˌ�}�D�d�m�T��M��r��^l1��-�·��H�s���	�7�v��b�t�<���삋�`Z��啔��a�L�HyD��s(�Y�%t�^Z)��t�-���w'V�b���ňR{���+�H֬��8��5�q�UVTr��i�u�3Zn��j*������7[�:{^V�'A$F$�+դG[� N��EZ�9�i䛫%,�P��S+���*��˻��>}V�c㺨)&�|Ɗ��F�j��4h�a���AT�,-`��*�>?�����i����QK��E&#U��EUUD5-U1Q�S�������j*
�ӈ��(*���Z���AEIF�l�j��џ+Fj�(�b�h�U�E��1Q3QZ�$T�U1F��@PMA'�������Q6,m��k�61�F�F���1Fv�&&�&(�����k6ƴ[[b����UU-�gb�R����mEZƵTN0U%��d6���[U:
�i�E%�X�k-$Zb�X�������RDSK�t*�$ZBd�lDQUTP��f�hә�ɶ5MD�AX��UF�N��8��T�I��%�`*��)�Vǆ�-����X��-�ţ5��P[&v���v���;˟o��y��ϫE�2o&Ǹl[<�ڊ��l�:���n�6��y$A	3��J�V�{����˂5W꯵TrUd����ta�}^a�����tF\�w{�w�j��I�|�d�ȮӒ7�A>�١��Ĥ@��$�3��$\T�n�j/݂b��#�q�b������L�x��@-�C����ڄ+*V6'j3�YI�5�הk�'�}/*E*yY�ƃ@�k��Yw��e�N8kf���,^iO4��Z3b������[���(_�R�i��
����ʼ�дKCi�k�p���XM��_ffK��o�ֺ�Ԏ�>r�2ދgml���t�[	���59�d��{f���Ċ�̌��h����9Q���(��q���v+w��3绀ܪC�Ԯ3*n�����7���͔�[�i!I��ũ]���?�u�fFO���2�?\������ T4���3����x�[@����Z����1���A��v�uY������z!D�ANYQG�2M�1�v�JJ��Ǐ��I �>�X ȓ��c��������Ϥͬ�VٙQ������[BJ�-�����ӷj$��蘌�4�¤��ε�)�4qT!�0ĕ �ҋq�}9l��=
VNQ���Ԃ���T��qmSL�Eu{8Q ��Ͷ�[9�^+}k���W>�v[�7b3�`�#Z{N�w\��DDj�Y�+���p;>�P�4���.%�Ҙ/$�c'��ͣ4�ex�ܯF��O�e��j�Į���������n�Z7q;�͹�9;�Vt	�%�񞭆��ʇsi�?
F�t�������Y��GZP��w,�:zBZ�5p��b�mǋ��iq�V훛��=u�u2��1��p�٢�YG5̊9��^&x�SX�f��F�}ԔA�ܺ�=�1j�":�}s�����Y�ȣ���9�A�>��X.δy��+��od�#HjQ*HJ3Ұ�j���1qk-��cC�[1
��w����i�K<�nA�F�����<3�!�ȫ�f�/ݧjn�sDӾ���ye�vOl�`f΁d�f��|�!(���x�Ys]Q]9�)�n��3p�RS�rmj���]�㦛����>8)���Q�����"��vj�@5+yоՄ��*0p��v���-ਨ��tL�Hqm���6�ՌwtR�EW6���ʛ�{�:ᴞu��T��>�f/�T��W��=r4�y{���h z��;��v��C�e >��B՚�ާ�M��wy�Ε�
�3;1�~�F�#��y2��,�뻛vR�j�:6���R �Yr�~-f|�ܭ��v^up!�X{��!㩃�����k�E�F"��PId,Ҳr�+*�KU�dU���b�`�t{�m�N�6\y���4������VA��7���g;<Ԕ�)���ݝ��x���}7�zY?e5Ȃ�=\	W�u7BYa7@�{��u��z���8�PKg���wjC[y��5ȂH��w��Xd�UD`�}$tC���t����k��)i��o�b����P���}!��:[0F�����V2^��[�{j0=Iì�؎�e`'K��nJG%�h��8v'#UF��5�S���Ɔ��P�N���=�L�JJ��~�-
l��k��P7j���UN����+3b�\��3�������Ҙ�[�[��yl�LW�sY��M	�V�wX�ʻJU�<�II�n4�p+9\/8@K���у/S����*�4�������}�J�>W����(��('�}3<�����4S��J�`k=��u��M��nз9<5S�S��QV��VR�8�w���M��+y<����+�[TЁ�ŗ�b��df�ú��'Vg"Gk�mg��W�}L�^,3m�T�����H�](t�Nv�_b2�%�u���rm���y��m�v�12���`h�hZ=I������}�Uj�Q̷��;�"-����u��hp1�; �yt�f����2���V<E_Q�r2�R9{@6Kd�]�o6�"�D�X+��{�;���M�<#�h���x�`� >��UWg�m��7˅��9Z��UuT��v�	�Jyg�����ve��D�Q��#�ʥ�T�����l�,�H�vq���ͽՆ/zr���w��\JD���fg��c�����ؘ�x��]�prV���OP�W4i�[.��{WoŮB"Ob�4iՁ��%6�5���!S'�T����U�ꯕ\P{sx�6L+uF�g�S��ڡ�f�`F	ܙ8�JT��_	-LWC	84ww����걖�=נjil��d��eF7nQ��d�3%2yۼ9Z\Sr0{-�=�b�u���M����*�a�X�I�Ů!�)�\�E���]�J�ʛ��MZ|\_ޔ{po�u��|���y�
�Rwo���5�
�Tr�e�=�て�{?R������Y-�䨚EX�y[@-ܐ��פˬ/B%�c5B:�]�v�o�騘�����;o y��rc}����Z��y@�����kYLb�<G^�̥���e�eΩ}fK�N��j�)C�����2g��zZ,|=�@Yi�%�4U��#x_܍�?��|�h~�GUK����GO5�̥�j�ы�!��79�#���.z�~����7��~eĜ��ƌʫ�.s$liT	�n%� 30Pn��X��o�8��;R�ҩt�_�{�z��-H�f7�?f׹�Gv����z|�\��3SɿKa���rK泵�*M���"��n�`�GHc{xP�u;s7�d����d]:t��w��S�3l�����	d��7W�wr��L,~u:,t�N
w���Έ�=rmj���+Le1I}��s�Y7�' ��@&\���c��rr��+=��lOs!���='�C�E
z+��J�'[��bp(y��v��u8�d��W4�%�R��o������dRIif�E��j^��S�~c�^�ާR6[���SHϣ�d]͒���R#E30��|'F�l|�3|F;�W�\��s�g̕���]�ٖ�v���E[#^]sNם7��:���i�c�Ǉl�����	Ŵ̪�����D�dol6,��K�[h?k_)�;�q�ǝ+*8��n@�V���䫞aWU�Vf�zl�jh��Z�;Y��i��>����:��R��2�i������:(�K��W1]K=�~W��j�����syo0��"���p��g�Kܖ���'�٬�:��p�`Jފɨ���QЩ����.а)�����w����K��[u�x^��-�d4=49V�7)Y�|����;�zxZZ��j��B�;^O�@=yv�8��=5$Ok���F��Ɉ����R��<n�W �9���(�������EӠ�U�eH�0�a2�f�z�{��5E�����u����N�#����zb4\	��:��en�S2�.ы6f��r��U�nT(�&�	�s�v��)����Sj5os�Juuq���K�.�&9����ed-�ݚ���A�LH��wWU�����b
�Q�j���8"f�>���,}�/�	�.h��fs�����3��y�:ڪ����sE}�����������'��E�1YwŦ./CݿH��\��pz��PԗN@�EP��/���ȼx���L������]��u��T@g��){v�+j��إ����1��4��&�o��Q�腫��^Fo! �#�,���9S���fP2Y�@ݍs=Z��j��2���X��ڽ ����x��*w�t��zC�Iy�7�=��sI���ߌ���~��
+%m�r���nR�˘ٓ�ُ9�~�f#f]|����rG�'W��>�� �����y0��w�NC���w�ۦ:����ee��*����l�M5����=*�C��jO,]m;��Y����sso��H�W&�mW� �Ե�Z��|B�þ���<̞V��&�z)�f�������^ɷ�0X~��k��m�::�M��U�-�3)'����c��F���{�l���V�n*�|M�+�����/e5צ��Ri[�억�]�]�-=1�Jʑ��gj[(�7u=3y���{�M�#{���I4�哵6�b@[}!�-���s���;��Ě��x�)dtR���]ҧ�z�$�vw��_��Q`�Y�hGe�K&f�Ŋ���ߡ�$GwM���U�Lq�J���q����ʈYNcu�VLj6M�Vkk7��|�t�D9Fz���Ee,�3�Gv�,��eV�Ɂu:Z�g���p����G|2W?��|-�=Th�I�|�vI���0���<ؘ*�|��(u�����6��in��9Π�A��"f�{�0�y�dy�w���i�e(�Ȯ9SY��MP#���{�k����a�@1��Ќ�|�>�1ߦ�WmWn�i�K`��9��x�$�*��!eY�d��z�}x���f�Cm�3\���g����O��1U��ku@�>#(�yS�2	�J
���c�v��|�jDI�Q��{/gj�����w�_̚N�uu@��3�x�nӣ���K��u��1�	�p��GsoJ��q�u#�8ƕ�K�ꕧ�t�ot3�"��uδyod�zm�nIV�+��R��"���ͮ�->	��̷��� ^��P�g��C�GF���1!{i,������z#��z�������R�w���l���l<R1�˘Ŵ�+�"fz��[���k,����er˼������/k�����k����-P:r&������k��gk\��J(�*��R�4�1����q)KÖ�똣�N��k��[���\�F���V������
��&�5=��i�t0�n��nsYg�u[�!�� �jX-4U|@-5n�fE@mZ�e�s��l�e��^��Yظ �'�C��i���q��p2:�}���n{:V�k��y���%N+� �f�a+:!������i�)�TM�J�`M�e�0��uѲx���W˭lDf���@�z�ﴟ��>��+��U�q���}�'��{J]��J^��J�����4p��X#�FUr��#b���bo�zf����Zj��򏊡�=sF%���=*�j] ��}�r�9�r����P"gS�}�ܿ�)^�>[������(�|��V�a`Ηz�]8��rn��pG���ԍ�בh�;7��QC������0�O_p�����ȹP`�������u��	���-��UeՅN �WSXs6���d��=o86�?������i����
krl������nl�A�C4�ZdKҟ�_g~]]'u���z�Ch���������6�X�x�����2NP�m�W��-+�l�_=���-9y���MH�=���ʦ7kWh��\-�h�N�e�Ϟ2v�ܜGu*���ت�A���ى�ޓ��U{�;�9KkĬ����֥��Q���7*J`f[�am�UZUm��h���KMEE�����nI�H�+�zZ�"ٚ%�>�ٻ3o�Z��r"������^��Ƈt��4�E{=�q���6X4���Mt�:U��DDx�;��oQ�oW;�w8(���ߛc�� �O�ނs��>�MA6~�^��|/��e�t��ವWsp��֬���M��a���(vSp����+��᛼��9��w�L+A63%�ө�u����V7$�66��Q�s��r]���K7����@C�V�t���/�W�#r\��Vms�_u����r0����`os�1I(Ǻ�Q^k�e�4�*��,���n�-�{Od�[қ��p7��r���4��]+�U�,ڀ�{z��K�/��F��������	,�1�����Y��ቹ�,����H}pI09�͊�/`�:%�������g���3e��6��71�YB�{m���ҋ�v�#�Q�5uY�=����m�o���l�ȘYm\T�gl���M&SYr�؞t ���r����(q��ɣ)�饒��&l���W6����B�j�
T�9$������$�I�ܧßێ�a��Z�c���Sv���u>W;%�CjN�>����P�t�8��'D!�XM�ʁ<���o�sJ�pmL�+�m������q�ۡ���^5o�k6��n�X/8���P=�)D�{��Ŷ�o��i�c%m'�UJ�C�M�ʸ�r멝�m�lۆ�);Y;I��Ŝ��g��▇�'�%�K�cA�˸5�Ύy�C5_	а�Y��k�bѴ�����γx2��������gR�Q��+���'Hћ|0O��j.Y�:�Ծh0���)�
g�#���ޑ��sTw\� �-��h:���8v�uM���V�����`ݹ#˶l���nL�2�n�6�
�ʰ<�C7Y3�ièL�}���K�ufB�gc	&�ā,8��J�%�nk��h��b���R�A�r�.8)�A�h1eR��!R�q��k�����Yt�l�#�v�^$�Wwr-bwr����Eu\WGu>��^�B�}@fC�u�hM<%	ݩ`Ż�+���9@��R�Cz�����%r����fe�]��V-@-w�t��v+]!Zo.�T��I]䚢��u:4�mu��QWb��:+�T�rI	Y\�\��ࣸw8�Lw�����t����2U榱��OvGM�kyu��^�o\+^Pշ��jYB֠���R��7�g�.튝��uwϭ���3��xUMt��Z2ip7ի�z��3���K�9Wq�`�+,����ԉ�.+\�$^^���2�K�6d��$���fcp���$8���Utd��:*��:6xwvo���Ki�]3�<t[z�G|��Y)�y�sk*�է)�hm�TC����5��rt��ⶨD����1e��Q)�Ν���u��oa�җ#�l1وe��
���Mvh��͵5��E=2���O��Ѫ%M;4,�v��Ū_��P���>}]�ͲXR�7Y�m�ŋ{��K���1���5�O)(�m*n�F6v�xY�d�KbW��*�[XwyШ���ab���K8��wѐ;����B���*��b�4u\.���ͫ�&K-\&��2n97�������R�ւ�t֪*6�V��ƊH�Š���i����~_���UUACX�5��HŢ�h�mh4�S�Ѡӵ�5H�Ϗ�����TM$C^[a�������
Ѧ���Cl�@MI�mU�Ũ���������DTh��QK��h��
���j�:
(�ɣj��������("<6
(ӱ���AUT�.�l�t1S�klQ[Y"kTZ��1 ��Z�C�4�mgTD��u��6�[;b�
V�@V���"m�[V%!E;X��c;Z�Z�֍5m���Q�F4kE�;V�$��&��6kX+%Qmm�Z16��PL֐��mh��gb���颍�[��*�5N��jح�4[ccT:h�m�HPК�N*	�f�ъ�4j�� �m%RDM�u@E J!$����dU�=�R�9Xt�<Ӓ��]�v��90̹V���n�n����z9�wl.���9f.�֌!����3���7@d�J�͑3c..�i�?��د���IgK�U�,���\<�j^�~u�i�ɘ�W���4���a�K��>q��%gQ�g�e��{�ץ�xbj�m�g*�ۉ��3l��tu%��3əmЖ����m�2gd����}������}+	y̹�=��{������.z��V�?:uӾf��W�o�y�4]T6�ʼ�Oa�\�����/��O��;��s<�v*�)}������#���p���:�D�}��F-��㽎�b-��~�y����|h��dq�H<솫)	G�]=>�E`�+S�]9f����U�*j*��wK6�fֱ�[�8�U e��6)x�|�$n�h{�[}+��C���3wj�Ji(�'�d�����:��6)x��6���;vmE�����E��uF�Q�(o��t6��5K ,�w��A9��V)��/6�4�gL�)�5��Tq6{���bj �W>ݛ���7����KEf��B,\Ք�%���{*3�g�
��T����f�Ĳ�����sU���t���<����׮�B�I�.J/��Df	�e��4e��8	J��xrM��	n����8��)����Pmc��C�q�T�>ON�c����zRw_r� ����3;9���Op��)�7TZ��FM�NEH=׳��W� ����<3-ԏ��k�r��_��9�wdɤгrE>J=�f޻+gt�s�I�Fh�����'�v������-n��]A^��\��om���f�3(���Ty8l�uN:�&z�P޷a|X�C�P���qڷv�^Y���>�QZZ�)Ҹ<T��7�v[caB�Vj*7����0�^��gиϮ6�t��U��bA�]@��c�#���bU��ksz�{1�[�jYl��?P�R��E��ճ#3���u���Ŋ9��5�]Q�t�k�Ԭ�Ɩ���|�)��ܛ�C!s�˙��鶥��َ$�K�Y�a+*�6���M�O��c�1���]K�&��zo�wuGŖ|r�Y��\�ϻ뽄zʒ���>>iL��B������0��>ٍM��4��˜�uֶIc�17xs�k&ܡ6̇���ʥ�G:KwE:;*�^�u��.���`[լWj?(�H"�ڻn\�c��Ϩi�,Jn/3���,��VUr�T�H�?�����^��T��q깣>cA��e�6W�'�T#O�m~���l���9���e'���s��q��;Z��R��;acq]F��U-mp��|nc9O�l�`ɏ]���m�g�oX
��ɋ;WM֝�rn����go��k���O�޸�1��Z#&;�E�DW�/�r��0_L�T��f�ƞ:ԇ9��f���/^�ٮ'77N@�~���v���f*���W�c�t���.�#�e� �׶5��a��J���ےt�t�_���*�fHU�z�:��]-w�s�J	Y��'4���`j�Kۡ����)��_������t۟�z�pޥS6��WQ�;����۶Ɏ;|,�M#Q��t^�+t��������zVGz=�o=Qx[o}0�R�o]z8�O�%�y-&�V�Vɭu�D�f����7"Cpp
�u<&:%�ib���,h��dL]Lu�r{W�ivf^=C�2� :��}ׂ4�Ut,VT;,��x�寕�ήWk ޜ@c�Is��r�f�#T��Ȅ����S(کr.E��1�L΄wwTw�0��HB�?	m��~��r}��vLڸ����9=Coa����=�4��ā�2���\�Q��Ր/�����z\v����/��os@��V}�L�:8O�P��Cz�=ť������j�5�k*��u�L�`]��|uey.{�4p�+V��j���Pq�xZ<����fm����Z�Lf|.{]f��=��q�L�}�m7�Y���M���ܯײ���H���G��5_c�n��@h��@��I��(�'k�z���r�}��r�V0�����r�_O��d�x�I3Sn�Ih��4��4��&2��w�>�Wt�IH��U뎌��趹�ɩ+f��ٌ�#Rܡč�B�m;@�N�e���R��SL�]�=ՔNn�ni���]L�Ve�A_qKhs���f+w��sV�5Oދ/�ϥ�;7qn��2G�"�K{Y���>��K�j�k"���|���<��OS^5�rܝM��	cl�B���F�|�p3�:&t��k_%AΚ%��s]��$t��EL�=�Y���κոgM���2�f��o��M��̋؄��Vpku��n���D��A���~�n�'�	�AIoˢ�f(ӪP�) +����W_�\ȵivT�V�[��n�ue�]��ߏO����R�O�Ƈt��B�q]�4S��E�8Q�wW�=5P�u��^��<&c7�o���o�Q��Wh��X�74Ԍ���v�|5������j;�܀�lS7y����`�l����qyS�y`�����4��iv�K:��D�����Ӱe�m�ڻ
r��*)v�V�EIuO��%r��p���JΠG{t,9e���T�Ǭ}�'8�d���BaG������B���c)�2�:�6����0�,]�L������NoM�t����s^�3�q�T$w%����
i�L�Njl7�����Sr�V��`b���?�|?g�助���)��~�X�'���5A�]u��^�ڴvt�5�2���=��ay��,<��Xg�f'qny�;�bC���Wl�Lx��r^^<�Վ���m���m�8�R�R{�d�ոC�1]]��}���z�X��o�+a�9}�g_�����S�7
��	�Gv�'C��ʝ�e�Z���}���Q����RJi�u��|@䚭�ڶ�<�:��՘}G�۹P48�9 �f��x�:���z/-��$+3��uwl@�3�v���M0AT�1�S�إ�!����8�嶳��ӓ�R�G����~�I}�Ť�2O2��V��]X�_c3Z�z9�զ������La�79�=�?G����䭛���,�X9���0�M��'>�DD����F��n�S��}�'g9+�^�U,��<&9��1n��q���EaQS���d%���ge�f#��וO#�_�G�n%+P�{ٚae�f@����;�����QV�*�h5���
h�u5?'�Q5~�K�L������weq�h{�Y^��e�W�'c�B�1TH�t��t��DY�.ȁ�vCj(����b���GR���.���i�5V<d�}9��oK�l���\�k��#�W�F߷%#�;�����rT�f�y�,��>+4��&ά�VG���Iٕ�J�VGKX�GKV=�xsst���l���E�h�O�\ɸ{T�H�X�&:S������İ0�(��;P��&WV�]	a���b���ۮ����S4&#u_;��"�rl������6��C�����`���ۤ��Z
�&w���6��6�v���8��!,��p��8�k��������wȬ�N�b�(IMkfqmp����	�h��il�v0m���C�]";���{S�6�O�zj��$u��QÆ뎬�g�d)���t�>a��$�hlP��]���m��4ox���0a��h��=��I���M;�v��+��l��3���,�S�^�Be��Ww�#֯E��1B�Z2;��V٘�`Z^�1y�q���^�xMݻ��}��<�Z��6��&�P2�ڳ;��"6Ik�z����g泻��k YQ��E�4�L��K?�'�@����c0��a/\ʜ�͙�<,�Fh��*s��g~v����ܙ��x��!�N&��ݾ<��z�5��3�{W���/����?z�T7����~��X�{V\4���6P�j�vԽ�`�ۥJtT2�u˧OA���y[�5�s7q�>J;Y.����"W��5�����+�{CupHc���u[v�Joy�뛞�\���V�*:7�L��e%���X��P�Q<IƛM���ͧ�x�[�����WP��>*�ۭ�e��#6��5�w��7[kZ��m^����]��c�v��7��@Ww�j8T�T���v�m�r�^�{/�	"�_|e}W���s�	����z�����'wI[ݤ6wb)�?u����ɹ�jt=�u~*Z�ۜ��֜Q-��h&�J�bC�63S^
Ζ�����r��ͻ]ꈈwX����+��p��3�x�+�͝�.F�G*��j������j@� �a�$2Α���v�ٹ��ղ���wMnD)BsQ��K����E�����!��̬Rx\�ʳ^��㤠�1��
�޿���gWV$^�RӒ3ylM���]`7	�=J�ͫ#b�L�<��S��2������i��&"vf7(fl�P��u��8F�8n8�6^<��m�p�ٸ���ٻK�Q�1�'?)g��Wem��7���V��U�H��J���וg�Z5뺺Hc~~|s�Z�L�V_e�������Kl��c�y�H�j��lr���gmw���mˏ7M�z�)�β����J��R�ɉ�6��3�����n��㪺�>�s�k��盹���~��9W�ծ֛�ؗ�!a�T�U�/�/۬=bg&�b�󳩧Wcq��7��i4�Q�T��a!���qS}p�܈f3o�"�;���F3L���
Cd"�i��#M���װ�z<~�����)GfS�4�h�5w�G��ޠ��,��;5�f���g�W������n����#��G��nڐ�j}������eo �+��N-��1��;Qzb������'�])�?Sz�y��P/\l񾄲�RP�̑�s&	�������$3L�~�{�<��ݯA�y�sY�S=pm�=���$ʫ��ތ��Ԗ�D⛀��w��ų�9M�,�Z���V�J�\�qK;*���u�o��ٵ�6���H$�T�z�Y�ϡ�;ٺ�ۛ��=���ٗ�2 �o�6��Y�kV<K��+�FoV=�
4*�� �P��A燦��e���	ø�`�����Jq��΄JK�G@f$x�Պr���G0�U�����9ze����(
�����Q�3v�(��*��r���}�f�*�D,-[�2�N�%=�T�rd�>��9�P���n�/�`sj�T]�Oţ��5U:�]��)�[���Ձ�T����z�칾ή��A�\/=��.��L���?%�u�IT��J���̜hq-OJ�ff]��<�w��ƎY}�(X΢Ap9�+|�ZB,�������3R�uΏs��lZ��ּfs��v��v]���K}���/߰-�W�-\3����p���nz�b\�u�5�L�;���UZ�����{�ʭ�4$p��[�]�H�����z-��	�YMx�G�39Nl�}�;���yy�ۻ/ݩ���QK+�V��]|fֲ������:���´�Lc����{*��%;W�'����r�8Z�♹�c�{�����e�V�fZ�Cӱ3/]Ws�ĖP�@�9���m�h�M.����u^Q"�r�b�dem�C�ǙTy���ܜZ� 	�ğ����R�Euv�|����Xuu�ܮ�bYVq@���΂�RgL�m4�	�z�5����`�՝�^��b� ]2�w�Ŭ2��63����4�G�&�U5���DnR�
�qܩ3Zy �vPQ�����[���qL�ц\�{�+��qc(�9b����b��q��%����[X8л �A2#f�D�cTֆ��/����N*<e��i��\���Ddp�.ĥ�^�*[�~皑�Oe"�n
G��up�y�������v�pܺdZxi�>��H|Ŕ��3�"�7P�;A�.�m4�%���H��܎�.��[ݩ�Re�it+��YKj�]��[�+Wn�ٜ`�ԍcۨ�ĩ���wh+�p$�kV|���ܺ�`�t\���!��G�s�Z��t��a�5��xk�NnjT*�g[�{{D[�)-�C+�Pj�����T�)v��R�%=��b�͂)Oe��$�F�򻳮U�n����G�	&9�m2'o\�GE�f�<�8ֹt��_aJ
֝bx,��;�˕�Nwk��e>�
c��K�9������^ɵk';(�.�8�+K�|x�^Gm��}�_;�^���m��;5���Ô֧E,tn_
'�/
W)9 �j���t�G�71q�p�o N�g1��`���.�v���Drᜲ��r�J(9�����{b轆��)���vgRfr��%�;2�7�$�̘=�P$��v���:��J:j=]�ѳ�,�[7bU���� ��'*Z�-wm>rRY1fŤ�^��t��T�;+,���$Af��7��-���%�U�R���tR�Mf�H��c�;\d���%S��A�R���\D'b�l�ϻ���'k�I��h�ЫȦ�����Ye	#ZՕ��*�IclE�k��oB�J�H�G{�`b�u-o8��MFPĎ��ʵ�v�l��lh�J����t��v��e�Qe����>ŻC�+�B���DHajژ��Ým�Rk�q���u�4���+V+�3t\Gn2s��'W<w�]������yl�M�t�YG"��`5ҹ6d+i���m�{�½f����1:S7��A��3��(��a�՗S�L�:a�l1Ύ�*Y�Y�o��l�a2ojֺ����J�v��X�2\S ̬ǧ�F��N"�e	o=QT#R��y0G��PA+�eKVts�b(���%M�q���i���q�i�� Q�V�m����VJ��������s{���%����g!dU�(�q�[e3�M&������!+E<¶�u��#�A-�)�{ �瑡#@�Ȍ�-r����ƺ��E��/ݳ*��V��P�P��O9�U�Gݐ�6Axܮ�Yhnx=�չ+u��p:�[���8\�$yG�)�+$��`��	$��m��mgc%kF�5>Hh+�	N�MUkc5���c4Z����~Ϗ�UQ1T�^F#j�m�1;h���l(�4ljv�Ϊb"M�������HDxƀѣm���u�A����Z��X�[cdg������"���STi����clI@j�A@[:kF�`-k`Ϗ����ǚSmEkV��֦�Ń:�[jH�gj�6ɩ�5I��@F�Ѵmgj��i�Fv����b+ıl8��i�*�T����V�EF��:�4[X��B(���k��Fө��F�"f��b)-d����T��h6�[)�j��j��[4kb3��SEL[&������b
(tf�m�.\h$�
;l�m����F��mF���M�QBkEUƵ��4顤$����I���G���Mo�jإ��6m�t��`D��9(q�,gvcԞ��H�eU�"���:Wj�У������=�
�³`-Iuu��=����g�iQ�*�[-�1}4� \�_*|�!�z�.n�+��&/DY]g�s�z��4j�j���"��m���� ]���H�m�ƲB0�h=p{¶�IJ��ݲ�<��(GR��p8��F���)�ǈ�ϭg��7
+��s9]�d�>ۓv��l�y[Xkz�C��ql@u������S�u�����m�U�LI�H�ˏ���'�ϝ���f���f9P,�l��g����.و(��{�m�S��h��|�$WFb��򎳷Z8�x�Kd��͏>{D+��#	�iј��옹 ��q;�O+�k����m�{�c�1�o4�݋�oٜ�Z�K�Λ��]���떁��њ2ƃf�p+I�f��?z�Ep�=���_'�!�iOb�Xݥ�x؎TI?|*�| ��sϯm��a�8�X�,231K��g�j�s�P�{�C	��J_E`f��nJ����u��2�M�8��k\{YF�w܏�ڋ����)��td@S��^`no�M^�O%��ݗ���b���C�)HJ-����5(ϣ'S�So�����������+����m��<��)3��՚Ղ��+[��ێ�`�^��E���o��*���O�Q[���]=�t�\�g2�N�Ha��:�ѴTd�U�r��e����GLL�`��79xg{1�*�vZ�	���H*�֫ڬQ숟t�ǚ�<�����~��>ٹ;�[UB�U��Kݷ7�I+e{�����B��n�\�,�f�n��L��:�;��ǃ��>}���eqK�⬕ws,2�N���Gy�"�Y�HkbM�V����G��D=��}��Gp,T�ٳ1;�yw(f4�ؕ(%�^66�>�ig%��M�Šn�[����]�gF�KM^Y�<��=�^&ӭv������<��Bz��FH3&y���m�2�<Z2�Z�'PQ(���+���g�^0��t0�d��/}JT�?i+A���&$r��xi�׭��%�k�_xV�֣z��'���֮Ѓ��9�:>��$qq��aO�۱���"���n�pksj�Va���p��E⽝��'��7	$�օ�3�]�Y1�6/��A<�)�Ir�R��^%�Vb�Z�2:���)]d�G�;�N��;eπ���yv.�R�^iwk�0nu
nC{ω>�Y��Wn��
u\{���oy,�]˹�bH��}ӓ���^�ˆ���mY�o���e��ش�m�ܨad���~'i�q�uTn����WC�fM�+���	��&9�2��q��~�"�6/��u�{��m����mhW��9`�&�t���|��=�����4(�T)�AX��<����q'Y� ���L�s���bt���1�ey�̇����=�*�P�&�;����r�.���"b�!��Z�q7�=c>ef�����5Y9y���	��=�Пj����L����)m�r���UƠ�mY�/��^��w�6A�Q�k��]0d�8��9�~�_>���〜["��1i�0�	l�B龬w�;���6#a��̪��3z�2o����kr;�=�O�/��3�Kyh���2`��/��F<I^���al�&A8��¯��͝,���巐Х01[��nOo�Kk/c<G�>��r.�u�.G�><�Ȣ�t�L���O�JUÅ�S�E�ykg��+o���pJq�e�������z{�қ{�k�"���Jie��R�m�e����7iEuV-�]w��-qq���VO��wOz��Hj�)���ip��6�6��|�^5�V�}��Sn�j��D�r�E��픖s������D�g]l\{�b�F�cfȌ��j5^�(rS�t�ƃ�������\�]_���x�(�F�9#s5��j��b�z���v@�S>�]:ʄWr�I�[v�m�C��4�np��^ ��z�3�Dm���߹+�x#��9�y��2G�Ҧ� }�wꟋ5o���y��`d��:�ܭ};[y��G3������ͧ%r�o��������Q��>�k�`��͓���j."�D��j�������鉃y�hwN�a��p�-���gO�c�d�p��h{Fp�v�VIQ��C%�O^G+l�k����q��M2wP�6vMv�y��5M�T�]s'ԗ�������t����.���u{k\'v1L%pk��<g�O��(D(
c��M�F{F���^J��'�5ږN��Gn��4�u�w�)GBb��LCo�U����<.��;�uE��8���.��K��`�r�-/�s�l�ri;�އ�����e��x�\7ׇ�m�D�.�*�]Z2�k��w�G�G׸+XQ��H�*}u"�k�.����s��;����O�������Et����dκ�D*��U/]Wr�cY���[q���0�ovL���N�K'T8�N�ڙt�t4����aOǰS��Oe�����n����rN��YI^PU��e��%��<ul��n�7p�s�P�f��_5u{��,��uz�\�ݭ�W�'v�e��4�fmp��Kۘ�`��,����[^m%+�y;�
�]+ڽ��^�y�{8�m�o�Vz��>lh�u��q��ˇt�7��r
���`Mx�`�U���T��9��@�ʉ�,��v�����5���{������-��;�pG�6�Z�#���ò͘C{<�4���i��W)�0�R����l�9'�mH�OkG�:$m ���[,9�:?{L�VC^�^�ܥ����D�㱢�:����eح��<�7�������l�p��}+N�א��!6C"��e_34
�oA�7�:2{'��x��uw�t���i���H�vʑ��ޞƪ�h�qUhq=���GԷn��q��@�f��p��봵�f��b��=��*f��F��	�-sl�3�6��ӎ2�d��+L����v�ůmu�&{WIsyG��M;�r�ѿk�Y��K��u�������=ޝ!ĊO1�fQ��"� #�A8�4,44a����6r��p��/t�p�w�0�O>�fbo�`˻j�ͪ��hf|u�r����ֈ>:� �aC���ڥ;�a{�>q93��{p�U���Zq�8�I'_#��oc�ң�[2����.rS�E����J��W�s+-�[!+��C9���{�M��j�;�6�j�=�{U��܍����v!� �Z�⋎�[��Ɣ���*�fH/^^,{W�6�d�S�63=�"��2\���|�Y�҈p)a�����_��M���{����b�8^���.�%NՏ~�F,��6ǇYc}Y�W���V㛝e�Yd��r��B��� -�ٽ2G�~|xz�8�7��ѺO��71n�P�n��ك����Ί�^��R�H۠G)�CWXwA{Nk�qR�V���u)wvŭ�g���H�h�h:�^}��<��fxi�ǵ�5o&����K^�[d]��G���V�[�g;`�b���|�#J�6shA���w��#���Q-9&Ы戜��֫9O�T�XO -[��D���6��?3,}[�)ጫ���h־EI��wn�&��j�WrV˺}]�ߧ�, j� �e�=�TtGL�5�U��g>���y��ՓD�Z�*{�
<!-�q�o(�>8�ɞ�}���Ik��@��·���B����X�-|�"�#:"�l�w�&��3�{�(�`P�i���0Į�H*=�)�i巖�e�^>���{�X����tdC�v�t���ԁ��m�P��7���ɸAv�6v�U��z@�w9O�3Z���,h4����"����^�3�Tי��[q�r^�M7��/�#xXy��>����.~eH��0���J�����YMV��uoO7���U�;��m	\��d�u�`���)����
�;3�Ɲn�ٵ7#���(�g�خa������aV'Y��+VG[;��-�oQZ��먱�Z�U����poκ�d��5��t0k2Ѹ*�a,��o)){����~�z��b�Hj-VӴ4�v[����+��j�6�v��<��]@y�u�wsd߭g�oHO6Q�J�+U�	.ˌ�3��Yw<�y�|��Pg�_�����}�X�tP��.i�8�;%�kI�nl��<Ҵn�{����*���_K\��
Xg����;�k�����p���oGҽ����5j�W�>�eR��O%�>�1�	h�:5�FT��F�ݫ(7GeR�EVU_wWG��nSV�[q���ڲ`���t�9���;�#��=��$��<�u�5,��+o�wx�T�����	[ӹ�A+�TF��ʏ�c�Q
��g����c+56w�Y�l�k��r�!_P���S��$u�
��K�5������Ȋ$�c>�`�U�ᯘ]��ќ�D[���I�!3FX�f����6��8�ݧ''i��٭n�l�h9WW��i{ۺE�}#[�ܟA� �4�b�l�v�nڭÏ��Ķ�Xʻ�;+:�QͲv�AM�F�|;��x��kO�J�)U�mU��̴���m�.�������=��|��a��2sݾ�NJׅ�~�{���Y�|^}V�S7��틂2��8߆�'0z��Ξh;=Iَ\��
=�p:�Q�3�3��a�{���o�]���v�J�}��B����r�=�&%z�@�[��oq�H����9�(|��g
��WӦ�j�����P��b��r[�c۝����t$���Z�ƙC�ՍىvjZ����4q�yJ�B��N�7����{r�UB���Q'�`J�t�3�Eo?�5�{&����͏<d5*�E�՗q]�F���9�]�-g���J~wLR�~�5an۸i��6�-�<�
��MƬ��L^�GD�>>�����ٹ7�F���?��ox�:�^�J��P>�;,�1�sY<m�ơ�Ӷ�ʼ�wWlKx�;?GU�Y �4�YA+ʢ�⭖�-���h��k����:��׽lQ��W��5�|�#z|�	+:�62i�:��Y���ɶ�',��2o_w]"/�uz�Rb�RS���ϣ�oV�";�7���ڲ$,ZJPUۏN�������,�E��mjO6W1(G�ԞV����̧�#LN�0�MN���B��.�G|%�je�w9L�ְ��	����Z�2�o?�\YƹAly[ U�ַi(�y;��~H�$zٯ�F\O��~{9���\_끦�6S��i�� =w6�&�2�,OX��Wu�o��Ϊ�uy���G%��H	�b=��6 �/��Y��t��&��;vM�w3�;��l�����X~QhI�D�}��=W�T7���YTP��٫*�&��O|@�=Tt�2�+?G�f�WV���OLoԸ��'���+w�_b�^�%A�'���'�e�m�K>�\3��������4����W~���5k�}��%^�sWG��}�szj<ad�D�ǭ�F�ٳ��Y"�1	�e�x@J
�s��[�Ql噓�2����>��󑙱�5oR�G;>Pà6C�2"o�`�v� :h�H�"�[y5�l�fg5M�M�G ��hl1�����z������?�����{�����~�������"/������`?�w�p8p���?���A���@ABE��D aTCώ�Q��
���9�r�f Nn� s�x��bb`9�� 0��P\�� 4�� 2��0�C( @� ��3�% P �a	
d 	�%@	�a� $&`P	�@Ba	Y��$"e	�dhdP	�!Ph`	���i�@$"a`�P ���� !�� &��UY
a@i	 �B@ �� �� !
@i��  a ha hd@@HB  eX���T?����y<�O�De D�@`��@�ߗ��~���7�����?����7�������~O���?��~���QU��������(+��L�����?�r@�����D�`�����Q_���?w����A����|��?��'�@������o��@ZD	R  d�U� � )X$@$ �U� @UY	@	UYUXUYa@	aUd@F �%UdI@VVA�) �� � @	YH@UVRP �@ �UXd �  � " �UZD �@$ � � ( ��EW�A������ADDZJ�T)@�#��?o���!A�� �>�����~UQ^���<���s�?���a���x���4����
�+�?�?����0*�+��Q_�C�0���PW~�x*�+���0�P��������~����� �UEo�����������>R����������~����	?������TW��?�� UQ_����<C�I�/��� �|��`����/A��d��	>w�
�+�D�??'�����`���~��=�/�U��?�UQA]���������C�O��PVI��ja�q�s�6` ���������o�
T������
�k�Gv�-�� ER�J���&��J��*R�(��H��%#m)UR�-RQ�uH��*� tݚ��6�j5��֥����+U���vlV���+{r�j�J��
�-���,֭%۹E[Ll�U��l��j�l����c�m�ԫ�L�h׹�)���v��١6k �m�uڕV���Y��S[fѷgGL-*mE�Y!�V�h+-V����i-bՅ�Ƣ�V�T�S+]ή�bĳ&�U�[ZU��6Ҷ�CZm�   ��Wݦ�n���;���&���إj������r� �wrP�SJ����m-���oU�Q��5�=[��V�z�r�b���sw"��hi�:Zֶl�K6k3f��m�   ;���
	
(P���)BE	
�:$(P�D�
�l(P����U�[���*��E��7�.Tף�v�׮;b�:�]���խ�5�t�l5���ڳۻKB�UU&��ru�[�  ۾��tݴ;�xz����p�/LQ�5ww�ƺ5�Y{�QmR���k��Bږ��������zs��c���-�8�a�^��q����'q��jV���(��  �^�Z���z�P�=I�M�����ܻ\���y�z+ڰ�3�{���]�,�UT)�a]H�5q�����r�J
(�	T�F���D�3[�   ^�D���.&��gPP�un�v4c	]h��w  k�L����`[C-�Q@�Z� �əfjj��u���v�͙E��  g��$*�����Z�太QUh`��@�ק�^�H���t�U��ڢ��*ݸ���úе�ڗn]�-���J�ֵeX�ia�l�>  i�Q4*���6�.�JJ.m5���M&���4���8  wg P �.�  n��ٶ�jV��b]�m�������  s� �ۚ ,]� ::[\�  j��  ��` �;  v��(���� (� �vsM�Z�9T�l�m�/�  � ���ݥ��.  �n�  �u�  ڻpt ��  ��  J� U��  �6�[o�v6��c-��dU;��   ��-� G9�t �� �5w[�� ; �b m��  �� 
�u� t�D �x�~@e)J� )�IIUC#����O&����� )� ��z�  ����UOD� e*
� ������o�?fg�I�n�G|�$]������Xð�ѱ�v�1X�e���O�}ʭ�m�����l�zlm�����`����������6ɱ���}���zC����U?�����Gn�h�3j�X��O+oT���)B��:q� �N�%E�����P�u�$�j�u)�`���i n<��V�'�z�&5u���3�'�c��'�Z�I�t�	[�eϲkw���B�2�̛+�;��D�7I��b*f�D�vrQiͽXdH��U&�	��%H/h4�Q��ذ�I]�]��yj�\�MSr�Z-ڣ�� �[X����(,��6-#2�ۿ��5kom���TN�E+!��d��q�'��0'����/�.'�8��肬ް*RB�Mf�keoM7y���E�/{4a@����m��i����C�#We ��/P�V�Ң7�T�;�1�Ӓ�U�Lk�aS`㖭^�f+Y*�l����I�bF��%ER=f�46d"�mʭO��y���YJ�	���TkVRԅ�K]Ll`ŭl
4���pVM��Ip^&`++"r�E�X1i��:-ݫ�қ�i��b��* `�4���M���Ss;�0)o̎ͩ��Y��-m��N�ԑ��hmЃ�[G	/6�V���Zc_��3]�AGv��@�ծ�U����z�<
�뱩YS�e�m]k����K2meȴR�i�B궱�03C� ��B�KR��k�Z;A1�86i�����Q/�*�6���:kX7��#9xY,6C�C�T*��KN�fP��D������-&���wZs2�ƥIJ���E�-�q�rR���k V4[��#1SFn�j�^��h�B���ٚ�-r��kͻ����*�nPq���ZR��Y�w3EA�C>B�4mU$C�~�Ťa+m����L�>X�Xi�V�V�܈��M*�h��A������IViͨt�RfBY��7jP���N�˫z�!�0�-���!w���ķ�RfСK*�HP���%h��]�Vn�2��;�vm�@�������	j^%R]�l(�[JH�Mե�xdX;��j2a�.a�X�q�D���#�AM���D"��(Pw�%*�ڼb
[o$��+Lm��(����Kw&�J���L
I�lw��wY6[Ś�P�Ĳ�0�Rd�c%�a[����VSR��V^Cd�X�����S�)�E,��5&f�D�ᩓa��,�{�)i:�b��0��\�[J0��ɋ����X�>��abmr�^�����%��k,j�A��bI�yu���
L�J[ӫf%h�ɛj�d-�
�̂��΢��݋)��J�5$8�i�eMI^�/r�b��p��S0L�^�i����	Y�V�V�@�xkP�!�hC+r��툫~�!֢���0j��H�$�r��r�[�.��v�4^X`;yeM�U���jܝ��Z�I
��6�i�8IܣE��K�]�X�� u{ft�Q�p5Y&�E�7������^dІ�8���OO���^���%��]���.,V�LS\a`�3�@j��Y��JF���M.��v�n�D60���Ջ���C43$��Z��i7���H� ���y^�rV]��4���!fjV���C%ӺC]͔��h۴�f*8�ֶ\�U�	�2+��Գeb;�a�4YΑJA��3u�E;� ���B�F��u6��2J�pe�{@����!
g`b����wH�eCn�A莦�"`[tm-ֺ�.b�Q�f,�Q�Qa���Kl^�X3GecȢ�x�_�S����M-�n�r�̕��Q�W�����20ϻ1)��{�XK+X�E*�n��1J����l��V� çcF61^�IPU���аU�ͷ{6L�Ƿ���[M��#n�<��X�� �Mll=\b��E�2wxc���L��Ac6�p��J�5(�ֵH(BV�ͣa7���I��V���2ط �,�)�Qh�y���n,�j�i�H�LڎIF��x��(i�������*,� ּb܁R V�[�ʳrE	:��)��̺7hh˖�ژpҖ����:n�֗P��M��`܈�2����1�C�$Ե��6�1
�-��Y��Z�- k���͇�֣��6�92b��ǂ�f؋���ݴ��
Rv�:�� ��`�w32%�K+)�ن�EL�g��@�!��Փ�ރ����\Yt�1�]�>��q�Т��f]Cط%n�eW���5��CR�(����PaRAҼ3$�6���a�E����Q�s�Xenh*�!�i��G2hA6�J6㌂v�d�t۫��.�lT4M�Иu�1��^L�ea��� R�^�SWEkx�jB�j��R���#c�i
C!��h���/[V^* 
h:�6�oql�f��C�,�X�;�@���ͳ�BV5w>��VG�wD)�hW����LI��]��'��&wo;f�7����`�e�7B�{#WK#��YgsZ���5���;Z�*r��MLAJT�J���b!ܻlA��YMTØ�˦e�v�X�d�A�5l�0dFc�D�ʲ�Ӭ#���D��0ӵGK^Y�4�P=WF��3@�J������N��ܧt3ّ_��m*tF�kE"�ٖe��:C�1�{.��jXL���T;�����A����/d�Y.������KR�kbي��bu����T%#�ˍk	n"�F�Q�@�aY7�a�F��G:�GolY�{w#�#$;�'�T�77".2����n,���z�Stj:��s�Ń�c1Lr�4|��0e�A�\��ď
k�N%N�-�t{ǁψ��{å	)�T�E��k[zx��m�cJ��J�V��(m��{>��I�\�Yw�6��!XC�J �un�{+��!�a���L�0�ֳj6�f�j	j�ա-3����V��Ҵ�*čL�a�l�ȭ������8PkRV��h\"�t,^1��{�Xw����f���Iibpb�Ǹ&� Y���4�f��B��&�[u�b\����Q6D����h$����q��p�Vz&g�[A�(�~�U��Ө�H�ѡѽ9I�p�j�Ϩ9��Nd����L M?���%�x�f�rf85�wi��F($@�yx�%f6mҁ^�ћ�QS�>�M��*ĸ��]�"k66����cJPV�ZXFCXԛ�'xED��s�Ф�WX�o3T �vl�n�UJP:�u4�%��iT؂�.j`2*�Ӳ���mA-�+���M��ׇ*�َ͠����E���Sot*�FY� �u�i�ޱR+�YĢ8	�f�@]�ث�d�	��c	yٗQ�aMV�=)X�����CQ�A�ş��X�Y �;ڇ167�h
bj�pk֊��Z�b%V렳<�<
U��4�dWa$��0,�oiML�x�4�[��-��vH�s8X�Z2�#km+E*tD�	�
v~Z����2��"�ȣ��%C+lĮf����h@�x��]��U�xٶ�R*O��r���U�j|���3֩2�{nbJ�
��b��Ĺ��֜Y����,a�%�5����ٝ���oK��^e`,L]���v��@�-�t8�4СS]c)�;0�0B�1ĕ�x,��Յ��5h�q��iItE�Q�{V����0�M`���U�U����H�xr��d���J���x��&�FV��hM,R$�+.����ܲ1�����>������n�ra9�l��'Y���r��%f�U�Y����[�+E��!X�3)��!��n�l��$k%J����� �q�!�v3m7���y0m �7qlܨ@��h�շ�X�8Ò�*ܻ�a�Ȓ�#S4;�m�T�`L�;�;�FZߙ��I��
Uс��{i��`��۹I[�!9su��k%����E���Q�
���t^Q�  Ǧ�:̡��t��R�"�X�hS9�M��e֝K*Xh
��x+)�2��oYͭƕ�Ͳ�
<ܵH�V�tYQ�U��J��p���#5��B��FL�u�cTw�%��!��ff(~��7i���/MXW��-թRWX�F��C��Q��^���n��ok������ݩh�fS���O�{r#��$"v��E�"��i��(>���?�A�`�v1 �"�"	�s�Q��Cw}o��J*�l�NԂ^c5�*�YSe�V+�r�֕3	Q�{,�ӳ�%�;Z�^��\j�)
"�z�j�23Mf���GE��z�T-9Yf�6��ɳhS.�7cj1Z����* `zwh�3Zyw+j2�/f�2�k(c��=�KL���V-����	��"��Õ�j\�
(�˰��R
�{�e�����\���� ��^R�ue�*4�TZ
���,��(Ҧ/sW��Cp=�؁T"Z��ԆՖ�9�����tآ�޴3R���^�&���z�	�D+#�U��6\�,#Eؕ�7p�y�#j�>�U
{���f�4��n�)�9Ef�Ib�t*����,ִ��9V�^R�����"�"�3k�E�0]4�1�2�'3e��\1���ϳI-R��Ȁ�'�ɻ��)��f÷A��䰊�R��NӸ^�Z����X���b����j	-�Zl�Hޢ-3�E�nf����oq*�م�q�c2��fj�p���^��%E�����Zʙ�U�5�?�m�����%�ۊ�j�r��6X�M���E�(�gin����20oj�2�h��=eԭ�S;j�I���<��[�v���Ø�t��+��a�1WM�^};fA��(�Y��"�t�����;��df�wNV��i���Ȳ^�n��y�X�Ŷr�������.ux��j�B�S���kl�
sn�bʏ4�
񹍪H!"4xϕQN�;�kr0j��hZ+-��IZ2�bv&�/3B��Z���M�-���1#Q+{Y�a�JJm�BL�5qf��hS���u���@��@@���s�mfm�\n��e�9�WVٶ$NkCp h�5���mn n�Ut��%!����ՙ����т���E�*	�ѽ-Y�˫z�R���e�.`�����Xk�ʗa7���K�0sI�JxMIb#��z��o/cʌ��mʗ��ZER֞���l�4a�u�](6cVf ���5��2�F�)�h�QSsqmOٽ���ldѴ�An��m�AAF� ��h$��*f׵���#��Y�Ş���������ݳ���eK�v���\Q��c����Z�2 �4,�G]k�,l����m�Nee@�m��E9��&���[��al���Cr��P�ĥ�,No��!��:��a���cD����=����Y�'	��T�N:t�Vɑ�yvHZ
զ���Gq�;W��ŉV[�1�7��E����ۋ��nZ:�����s.�
��/�m�5�<j�ù�&f�J�^&�]�u*�Y�7y��eʏ5��R�%��
x�lņ���2�Bf'`�b��w*��[�*�7���e���o�+N���7�$��Ջi�BGS�ʎ:�]f\Ү8�i�GU��V��7
�,Z�l�j�r��M0p�%���l��{zi���6����!QMK.����R���yN��yq�_4BL�w�<�Q ��B+��J�K��^��K/���4sP9��V�ݤHX��ƣy"�{�Mq��ۉ�۩������-L��58Nз��k�f��5�W��{M����Z�S� ���252C�kQE�c�4��#F0p�E�ҩ��,��MN���՛I�v|�+�%t����A�����Hur�sh�`Z�^�t+\��!�L�4�e�ěb�'a�,L ��,�R1���*\$�M�{âYH�sZ:�0ò���#VL�D��QSr�֮��E7i���oФx6��s(Z��]Y��-j�n�hFP�;�(k�Z�iPș37���*ݻ@��Z�ց���j J��t|�Ytb�/N
��@�WG1�h�eMI
��pJd���6�ѡ`�B<ڦ���,���o^T (XIYz���.��}}_p�fɱ���9j�ۖ���qݧj���3w��`c��U`�U�,��.蝏S�b��<YM|�[k�y�8�T�v��W��J՛M�'��3-]����ʽ(����YY���K	@[n��i��ZI��jܷ�Q�ǭ)��H��P� ����@�r��(�e��w��t=U�n���$ֵՊ�p��5��^m��W%���30�F�6�Ήa�dC	�ނ\Q�T�r��ߐ�h���@pZ�y	VU�5@��®���4����c��G�X�nEB�2�Z�h˳��UӔѰ�L�aQ�m⎤է��{3Ei����L�X�!�_e]��A�J��eAv6�#�7/m*�0��F���A"w5�n"�bǻ����r5ge�5�R�u��̳%�~��kn�TÎ!�T؁�)I#�nk��!�,�4ѧJ����j�d�r�L@8h,�.�����oM���ư�Ej�;�D���a�+�/��K-�ь*�J�7�]X�GC��S�r+��-j�aN�Pt�5��IL���-V&�9��sTs,��:I���c0h��j����)Ϛ=�w<�thO�ӭ�j�ـd��J K��?k�9��+b`)m%���:�۶pIHSK?Hn�Kq�#�hS*�;��W[��V�1^2MS�P萗{����B�'�1m��M��>7e���+��dY���t�7J��N,�tF}(�M�qe�vi�+��E_�ᜧB|���s��oQ쁾�l8�k-�Τ9�˙�y�\�& [fӬ�O��k�wO�JUt�֑����qO�H/3[��[ͼߊ�HN�=��s�Oen#4`9�T�s]#�L�V�&MYԕ>̔��{��I�q��O4�IM�{�����T{������9>��N�9F��ho�)/tQ�;�5���T�rJ]�im���L�C\�`�J�kб����h�6��1$δF�a�F�E��W��ֽ�u+���kh
v:�]oe��ajm�0��ъY����u�y�r�0��#��[�YDP��h�A=�吣��;�D����.��],O������oQƦ��v�ݮC���v>K�r����@��{��]��R8�'�;S<�6w��ذo�6�؆���H��c9ϰo85ĝ8�@͞��Х)
��3'�^��<wE���{w��PgX���t������%�r��O�k
iq	�riv�Vx^���L,��ůgQ������Gqe�S����=r�	!���M�X�Wc���=����s�:�<T�����i(�DG��� ^�T��+��'���u'72s��{ڵN)��K��{}������y {	��=~{z׋IK)� �;7�� ³�'����Hᖅu�+� 4����������-�s�Q��f����R�ɭG�U�*���RU�p��#'x'z�Ѵ��O��lG8�m��Ov�~���x��݉4��+pS�1T�X�'��	Tu^�:�~g��>��p�=��qq���:܎�zUƬu���1���+�^
�A:���n3��
��y��Z�{��iθׅ�^���A��l�m���Ѻw�c:�>[���,M���Ia�	W�`���ڽ��Ҍ��R���\�����i[�r�b�6�H��:����B�����@\7���;wL��R����s���*���u/�v`t�Æë�+o��e�F�ƽukt�N`	���vYn��\�^$�h{͹�/F�	m<�K8W�<ǠК����LRN>�n
[!ygy�%N����LgNz�v�c�j+��gJ���Z�NjC>2q��`�NJ禿j��$��pv�^���16��I�h���N*��n޺d+�n�e;�h�A����e�prw�	�.%1{���˚	�lX���g���6ss�����_�O�&��k��w+����6���kh�B���Re�6Ӝ�쫑�vqwf|�R�]}A�M�N|��ײh���≭�`O$��fY���r�8����nB�A[pv+�r�G�s���Ʊ��i���n׃� X���t���&[9��/v���?�tm�G���wF�U��	�j���%�x�
�`-�MoWwX�Wj����%��
b�:�q빛݋;1�����G���)���6�B���3Nm@��^�O�k0���~�`�y�涹W,�P"M���q��������Zyt2�i\H.�s�]o�	qg���Ĩ�]��ӖW:�Pe�R0�\*v��R��ܔQ�;l�� FQ7 80��O�ӕ4ݺ�k�1�t��/�"��46��,��-�|�5�׻�\�,K�U��mܠ�ˎz�y��25����D^?)� ����� �᧢L�g���d���&E���kIK��ioF��f޳/�ϗ��U}DfX�e����F5���fo$��H�N�!����t �1~�G���1m�u���L�Kl��(;�oNJ���S��fQ�JF맧�7���>��/XӦ���N�����i����K*�Q}���=��o�����E��.LΩ�	�D]jmCW�5y���:^��f!>yIFK�s�1�%+<aչ^w�Kx��xe�s3��W��w�Q'd��x{��s��a� �cN����#X�㜠��n���A�Q}m��%7�]��Y\�:ݗQɇ�a�vRB}�f�8��s�)"��V*y-?���q��/�P��X:����r�Y��Xq��C��8���j53�P�r�L��wq܇�#�fc�bq��M�,�5�y�]���j>�������H֏V�=sF�A�g�w3���+���J<��af��;�K霁�dlC����M�<2p-���go��[�d��M ���&�����P���k��&s�٫�ۀL���#���2�s"�{�NO����B��p�	'\��\glSw�;ea[ �Rm2ӈ���n�[WYZ$���q8�oW0������� �X%r�{ٖ;����{mf	��%ok�ivx�T�;�'Bd����-�7��_nz�X���`�orvu@*�ُQ�GhU�+9s̋GB�U,�Pf��+�s��L�Iv]��L�B�hE̼Zk_\�8\c׫0���7��NM�fN#3Vz��%;��G&R�q-�ʒڕq����Y�溎on;� Q$ F��ێ��3eV͒&��c���q>�������`���rX�k��+�φE���:��	s���,���fos~�X���yu-��GJA~7�%,�^l-�(��T�ە������͚�2�	`��󱮸^�z�6�3;]F�\n�/hQ+Ni��ѯ�i3��j�Ĵ��$�hA4�'b\r�*��I5��t5IxJop�FW ���]���:��^_�C�쏞c�*�۝\"Bև������QK���E���c�����r�y��Wc�6��w�w%���2��au�!n��<�31�����q��<�Ή;Rx%ea��WW�g��l��9����ή� ��+PH�#Z��D�CnpΰI!�kV�]r�Ecp�����V5QjX14'���ڂu��B�&�t3E������$�BXI�q]�Ӕ���A��r�KՉ��v��\J�N�n��3s`'� �::N#9� ���ۄLP��!���Ӄv����H8�[�ճ��B����|��P��y �bc�z.���y�؄a^�e
1w3-6�1��u(﬉��-�	�yƷ��J����yi3�^��{�!e��o+���$q�%Р�Ny{��D����r�g&�VgdId0�Ҿ��q�i�lzZ�ȗi�N!�����By}�Q{p��7v���d���r��cO-b��U�@��Ρ8�zB�Z�N��G/.Ӭ��ַ20�7��=�GQ����j�CN��q434^�ۦ�w-�M�;L%Bo�����P�֦��v#����6	��� g�;	�g�I�Ho��Q��]2�!hcI��`k=q�wndc�}���<��#�3�������\��M�Ȗ
;N�"�лW:om��\��Ǝ�o� �Z�4ހ�j;s��7�[;Ϗ
ֆ��;�F���+M�N�͋5ޞ�����F�>��Uu��źj����=n���3oAL�A��$��im�ۢ�9Y�h&5ƼǛ�n$��n[�=mY!��
1��5wN��X�8+�ݛ�QU�CJ̝ڸQ�Pܾ�n)Qܚ�]u��*8^�R\�2n�g-���q:�v���{y�l�9�+���V�N���\ә�z���){tL��ӆ.�7��`���t=`����0O�G�>�9����%h*��,�a:}�B��A�����{���.�Fb�m��o����a=iD����Db(�dS�:�Nކ�C��(���y�ӝ�c�l�,'3�)���fg>X����/m�$
g��Z(��iU��p!�ɻ���o�6��wE�٫��[Ѳ�:8���R�w�~G��^ԛ̶w3�.yʰ�ݸ~��*,����53�t�+w9!����:Z2�:8���iuwp�#WΕ��2Y�xmV�����O@3 ���qK:�/�5EuĞu��p�����+���Ga�o��n2�nh*�1,n��Ȳ��������]���	�·m�tE���%?�]�ǆ�|5�e��=²��	d|��Iۛ]qc�r��?�4�jd����)�O�����q5>�G���)�xem�6���h:��x-<&�W��kO�?��-�������!��[��f���O�vœ�;f�{�S����oW^<rt�9�v�U=�!_1ɥ㍓׵	#���Ek��X]���J,��`N�|%�zV������)y�ޞ��-�L���A�ո6gFn>��Z���u�Y��\�]+���0䏟��(�\�:�'fѐ�M>��/M�%�@���>ٙ4��z����w�W"�ֶ.RJ��;\�h�2��(����gs����R��հ1����$Ut��G�����z��v>�<��Gu��,
}{������~5&��Få(�b]��$ˏC�A������na�=�\�&h��M��C�D��ө9�4�3Fx�+�v�[܄����B�KtE�I=��}p%؇�w[P�xx�j��:�Cz{����م�h������z�(�k@�[�*�Z�Ԋ��Thd�b�osh �R'{���^�O��{�L��*|}���6V�JiU�m�
��\�,��JJٻ4�,��k����e�+$���رQ�`�e۔��#n���}5uY�`���{�y\��y��bv��U9ǸB�KC�IDtV��⮜딇��c��xq�l���8+���(y�ru�~jl�xz�ݴ�f���@E�srۈ���T�;��i���rΖ��zy����2ژ`��*)�0�wڒ�:z�$|�^�N4���{�D�
���N�,N�}l��GzJ ��;C�*����Q�v����/n��sAU�Y�͙��+{Ӻ]��}ZݿC�r��ē�o$M���V1C;�/`���L5�F����p�`V{�����PJs��)�홻���t[�a�S1�R����B��تJs�=�J�}Կh��qu/.�r���d䣨�9p�/�h5ա�0�Z�(f\�Np��J*�9k�/����U�{��u4ap���ca�dMy亍S�m���[�S���{�Z;���SЦ�o�E���_f����t���;4�k���dޙ@2\=�oj�>���Y�����3T��yYب�k��Ů}w|&���de�.(;AZ05W���Kn!|^���s�i[Rl�_J�h��,����.�0���N�4����:�|�n-��k7�)�ݝ��K��p�Lr�9��1�m���5,�g�v�!��e4�a��V^�	�u��v6W��f��&��<|�
�uej�fnh�Ar*Q���9���.�Ґ] ��Ĵ�n��/(>$�����ф�[�(R}���4I��R��RfμU�����9�b�Y�f�'�p�-}-@�-����w�b�����갨��R����T���k��V� �j�_�M7���-Q�����aoH�c��>�9j�&��ob�H�yLm�]��`(���D��+���V�ϩ�d��Γ�J���n�u�Ê�����stJy셼����3�5�o�L� Ӿ�v�!��63��F"��39�Yr��T��\ʷ�;qJ���K=}��Gt�s�)�r��M���W<�Ut�N��>k�@�'�>z^}\ʒ��Ͻ�(��h@��
�ӧ���"OHn��DKU�d@@�AQ����>"A��#k�AfT6ku�z1�I��ޜux���8���O@�J� p3qDJF ��}v��Y��L�!��zNV5ݕ0e;�W�ޠv�C%��e@{=O����;���.�<�B�O��J�s�J� vꭗH=;�kd��ws&/!���ޕza�:f`A�6��r}q���zw���1.k�����C��w�:�ٙ�+�j� �\��o![ة���y��&�¹�fō:�n��4�}�t�4W��Z��=��D�=w��u�4M��Z�z.�3���{å�%W,Z,�ޝ��u%�v*@����X�-�P�[|!�Me��з�c������b�a�}��O/4B� �̵y��p˃�9��j�����4�������Oj�\�t=k�@����[�/a�<3:�F"�<kG�V�����������ܓ��[��n-�M�� ��ƫu��}jK�%�嶕,��&��>�ǲ�\�y�s`���Oˆn���}�A�%�_c̪yf�%��d͵�]�`*�2��)�S}y�V8�G��bŔ7��@Й���=x�5�����ۛ�����Zr���T �yp6(R�a���\*���V�t�9</��wH�v��&���6�1�L*�x��"��w�T,^N�+s�/�ΩB�Ϋ9��L��xΥ!|2�g��J��]�`�ax�*�J�C��-K���Wϔ�ܳz��&��sz�!U1,�x�ggc܎V�l��f�!ھܒ��� V0�f8�a�����+�;���f�l�u'`���MQ]��E��ܬ�8�����ָ�qެ��$��t۬k�L���P����w�z��v{}���8�:�m㬔g�d��^��E�o�)�ג*�WC�t�3*]������p��SQ1�pr�pe�F��ﲳ���F�<��ef�7���z����Oq!�Vt1z8u%�X�S+��*�c��C�
��ks����XO��0�raT�=t����Z���rP��,�r
M{� `�̩��ց���̛w�Ѷ���4��J�-�k��d�P�G�s�N�ׯ/�S�_,��@���O4�"is����ݸqb:E����t�\�bX0�9u��u#2P��a�_,�����P�JYηy��>��-ܢ.��t�'Gڝ^k�;���ٙ3`��B*^�G�`����f^��p�\WS�'��L�9r�۬���j�>�}��ƠF�\�f�:Ub�B��y�jNg�[{jz��8w���#ccm���cm�k�w����w���i%�A�����r�!�&�>�S���i���$��:|U�T�'׎�?KR>��Qj�7�`C��w2� ;A�3�z��*f��R�2]v�tu�;C$3��sV�x�zP���u�^�����$:�rG�G���
`�c���9;o�?�dm�ͷj��f6��)Ы
�KΩ�d>ޔ�xZnJ�ȱbYە��g Bb]��O����b(tq_�$.�S���L�I5gS{t����;3a�����܌(�
�wӞ7[qMJeon�x�W�a��e �������M�wo�M�����rno{<�^�7��r��8l�殓���"�A����qLv>Y���n�����u�5:�:M�*U�lw]n��.���.h"ݽ;9%1m�ū\��N�gu���fRo)����p[\��7�k`W^������܍g
ϺIB�)�[R�0Q���Y�W#R�yݢ8��X����b�*8��TW˸�
�gF�˶�:[|j=&���rh�f���8bEZ���X�w��"�s)��m�E>�{�%Z�e�WX�����"���V6#��M J;�oq��\@q�V�]�c���nc㋓��Rn-6��"o����)�am��-Ym�稼�[C�_oK��O�2�����%����6w�˻:X
�{z��͒�m��g4?���Y������d�Ɂe`�[�1"[��kN����n:o�
�|8�6����t���1���T�Q"��bCkj��&�+y8	ǂ��\�7-��ߕ�Y4�l[�(��˻E�u ���zpku�,�Y��x�7���4�zj[���FZ8��S�{�]ک�ÜljT�I\g���W�n�TN��U�f͂�]^t����Q��0;���zi-��s�=��s��}=7Tt�-=�b�ʞ)�b��_��Mćk��/��<�3,�"�d��ZPs�6��-��C�,Sʴ���w&�>�7Mrb�Fȶ�q��ӗS�����֜+&�}��ݧ���/@��Q��޹�;��`�6m�"�z�B�+���pA��CGK$3Gw}Eg@� �SǮ��1��![�";$�}����f��i:�mb�+�
RԮ����VU�Mg��'T���t�'F��7;�?�q�y��|�9iq*4F��>^��Ejb۝@�sHƖa���&�^���8�<4^�4���Kf����ې�Qf|1��<R��vgQ>Pv�i��Af)�0XTn��Q'�z�ďI�����"w]X(�x�D�;�.\�wy�O"����쳈z�v��Ghӧ���;�hM����RZ��� �uL�݅������Q�� ��(Kk�;l85n� z�8U��O�w�8�3���g	�4')g�cr�`�?wjhR�Q���9�-��<ѷ�x���4�g���e�@Os@�Ee���k�}ۯu��B��1c�>���B&�+��+��Wl�xHxB*f%��W�Ò�<o��/+GV�c��I��y���΁`wv�z�k��M�{;���{��_�P��B:�ɴc5�2mg���Ǔ�0���<qecA�m:�meE����;c�{Q�۽�n�}�|�|�0��
k3����Cz��Q�~;��;zЇ���5"�:���u���d�q×7R���z)NެT�vD�a�b�葡@����cr�$�{�WB�ј๲�Uӹm�#�u��5��=bo^v�k���b���\yA�5]W8I\*թ\n��ڻjǦ��l��|c�ݏ�״�D�ō��6�nu<�˼2��9�8��� ���Ť�k��\X숖 �$�/���Z��;3+8	��^�ĩ�eI����5�3gp�-R|��4켆b��اjV�N�E���v�|ה�|cxp1W_i��$�����\�3���]s��g"t)h����z �Nv!O~���.+6�I�*���Q'[`:3'u6f� ʀ�r�ځ�z,�4�˯x�83ܺ��c#Г�f�$��Yx��SG1v��o��owc�V�ļ�y��S���1�f���IM'L�7w��%�&����g��4�T�Suľtt�B77{,�/՘�s��`��h�z�7(��ϴ+�,�c.�:�m֙��g��]w75��� ��7C�Bh����(���՜��/���8�}s�����M��+��׋pwz*��qJ[2kk�`�K����)�v�H˭�$��SWt
��TX�{D���G��b�$p����Ť�� ]4�!B^I۷V�X��W9���7����,2��3b�{���T�M��&�n\ض_�C�4#�����:��jWdv���H򥯮���K�5Ǝ�43��b�P�
��J6(@qS&��M��`��6�=Cx�[�%y��I�`�\R��m��3Ͳ�ȒV詙�*a��Jz��2un��9f�x�s�~^�� 3�@�`�9�Bή�rs�]����4�{�Nz��Q�ѓj���a�s4"S�)�����/Q�̊fmm�m��BmM�f1x�f9FM2|�P�O��Qz�;�>��6������4f�Vס�pۚ�q� ]��w��(¹
좣�7zt���o-�mc��ᒬ[�&M����((T���T��0V��"���n�OQ�0?�X��aU�Krb�Z��u��i��=�x��<7����4־e_�ҋ�`�M�H�z�b��@��*��E��;��.��kҋH��
oeִOd�.����ޝ�ۜ#��Y��sGj�C%��Sڊ��Z�/N������4%���t��GhwY��l���J��1�h���#Z���|%�J�&}��s/Q�-B�=:�<�C�� ���۽��T��Ÿ���G*]�.|0���#���{�݃
�S ^㫷��t�X�a]٨ZPZ!H�W�ò��q�TA^U�Pgv�^�o���yZ���5QPy�yC�����{�nf��P�ӣB,�&tNV]�_vc�Zk��r]�^��'Ig.�BZ��!%[!��:�vAK�1\��B*M�L�@삞�ڼs~�sZ�%GS��ަe��z����Ĉ��n,�®�� O��'x��
e��-�jG�^���i���ܭ|�����z�:�<d|���CEZr�_!�shO5.ƺ.�oM3�%�z�<���w�b�0��m��g���I�3o��͕��t��2+��i��>�d�l����� 1�-���`(+D�M��Vl>�Uf�1i���8!�oY��ٿ��4OL!�<B�c�aVf��h+\�v�ˇ��Rζ�<�Gx!�gl�S���ի,�ݵ��uXR�w�!���}m���h��>�7V�,��F]I�1H��Y]��Ϧ����~i9rv�m�z�嘭y�#�G�a��#�FBa.��/��7|oo�ݳ][��h�3-f[���u2���P��\½�c�u5!^P�\��k_�Pn�w��z\Uٝ�l;M~R�hw��$�k�cEk��֩�.'��:��:�֋X��N��K�S)��\����ԝ^����hS4�wC7�=�����ا����.�� #��V#�B���sE���� {�Ya���1es�� `%�9|��S]$ 6��4n������ S�k��z�a`�(fޢ�Nv32(�FmQ��%׵�%�l���	$��)E��Q�H0�h<��p�����7���ī�^Kڄ��4fh��%@�)i�u.Yj�W L��:(�rf�	��I3��K�'�|�f�P�z�����XY�SDfۭ��L���;�� b�nv�������7�Q�\�@҆��z�:����%�^�*�6��C�y��"d���� gNj�V):�|�ݝȮE���\�3_lL�X��bݤ����;�h􋬋i�%*�Ei��oy�c�"F7dV���z�R>���ɔ��^ē`��'�`f��1�����r`�mYN�ذڧ6��'��}���;D)7��m�J��ش��+���x�u�L���/�b��_:n��99�j{�� ����$T���*`�:+�u����3|qҢ��!MM.n�ܹ�bKr-���Jڲ7�j�cݞ�Ֆv�x�l�U#��h�tk�\wU�0�d�ޢֽ;;e��;7���٭�"���Õ\���#�����3,���	qZ8d��a�.Pɸ�{�9�W�?����wEk��^}�wPA��	��Y	Q�jt�Pq�.��o/M5��c&�wu�c�w<l���U��ŹB-Cl:�<���h�ʺD[l������[/��#��br��̎>���N/+�=�X�@�@jJ�Y�3�,siS���9d������V�7ތ�7���Ȃ�A�Zw��J�g0l���yn浈|�T7�X��׽;v��&J�.�#�'.�E�r���U�{�L	�fi���W�0iw�G�p��X�K����n�vvn�ڹ����n��`�h��8��i���0GE���C�<]'��d^F���FGB�
i�9�
���;o\�a�b��K}A���} ��I�����۾E=2� ݜ��D=��u ���"��N�vwc�)�̫��k�M�c���s9=�~Ҡ�]�ڼ���^(�Ր����)�)]wN=�tؔ�7t�3j�a�\t�8��H�0��V�Ҿ��\�^���*��2t¹ئ�
6]��X���Q�\��N']6+8j���E���Q�#�v����sin�����/������"�F5 �ձIkĐA�m,���|}�T��I�]�;�`^�<�iM�OC'��B�QL���^�oT���tjWr������)�p�1��Q��s4q�3*,#ꪆ�Vwrǧ�'��Q��S�˨���ᷚ�C�O>�讗[I��V0�j�+{�Ix�Zc��<ʭ�m�eɻ���p��{�|�/�6���T�K������ٵĎ�q2ދ��(�PjEG{'�}���(]����9�^M�QQb���b�Z�X�P�}�R]�sM8�R���6�.�k&T�C�L����(�z��ǰ֧�'���A��8��=dp��w4�f>��of�;����QNâ��ظt�k^jdb�T��:m��beum#�t���ͺ#=�Lr__Hu��u���x��b������n��������{�d���N�F��eK\�R#]1�(��ӂr*=��xŻyX�m�K�YϙN�t����O��Z������]���.��k����:<qU`�ݵث�9�����[�^դ��Hïfv��]�M���X�2���jp|��`pT���/�C�l��}�y{%bL��1Ȓ�<�27vj Aٕg�.��� R����{�:�>��|��z%xc2�c�\��:�B��bJD�w�;����'̏{��R��O�؈�߰���Vg��ֲz���%��$��+7�m�j�vt�5�m������QN�εS:�%���T7-A%�����$70���|�d���	�0f�R��B��)��X��3�YYͭzf�5j�l�A�B�G���P�\c�xi�:,�G.��2��A%J�+�}�Oy�9���q"�kY=���7=��Ao�b&|d.���iB���F��1��/�BHl<)�Xn��$+8#�)���0ٱ.�����S��8;o"a\C�u�����07r�'H�>޽�r�NcY�I��P�m�SՊ�d�ˢ�+e�OjӠ%�:&p�
Ht�*u��s����/-�wW����LQ)^:�j����l��[g��PJ�6��p5R�����\w�:o�<݄wg��cf��?#���q�hIz�s��}�����S�-]6H�̇Sh�7@G���:f�:z�#T�6t��'c��;F�Ӌ�m�^3�tnk��,A�Ph�t��:�-�'��[�f��j�Si�)���Gu
����UH6j�N��ֱ�Ț���V����q}�}K9����.���ğP�c[��*m*�,� ���}R��k��q���x�;5s�;w5\d�$H˙�&U�99w_5�t�g�i
i2�9�4l�*%���%夥D%7SZ�S;�ڧ��0$՜��x)�f��2�旋}����	�v�%����w�/-7����3B�#=�g��V����FJ���cC��鈷�7Wq�Y�
m�qp2�����嶹�~�-�'�+Tr��ܺo��d���8;�{4A�xy���,���¶m�f�<wh�f����A��Y[o��y��n�Q_@a\�k����p��K��a:q��+�v̷��D�Ck�0��BNL ��5��u�D�� m�r|�^�ܹ��ۡx2�H�Μ��;���,;�e�./��U�|	�|�<:�fP�9e ۬��!¢��1����Tw'��>�w2�W����`|�.�Z�au�o/��udf*��w�l�De��鶬X��G�Z* �ǚt7�0��|e�z�6��b,b�J����!���r�u�L��u,��H��l�Ў���w.�;��o8�8w]=�c�����F���TG7%� ��!�2��&��9m��U7Z�[W���MPI��Ol��C`�*�(��1Յ�����k��ժ��\��`����U�h�Cw�m_E�`;���,K�\�\�	t�j�`�ht+k5,2�9f�^���,����%նå�����o��R)��u�t�h��h֛X���$�:�jeu�ֹt�i���j���Յ_P���W8m��J�5��GW;����eݙ7)�� '*M�q��������?�k��ُ39מ嶞U�MkT���x+,j;����I��=9�P���䀵SG��"zS��IߥU,T\;��ZoC���Ƴ�Y��r��;�zx���yN�^���wFbݗ�3�����.��q�X�=Ct�2i8.]Qe��`����}:�R�n�&o��
^��H��n�؝J�<�w��u��_oI��Q�a��>\��~���o��RgWQ��-�Vk��R����'Lzy5­�����3��6S ����=��Q�D���Ur��o5	�lMZA7N ����o�qKuHi����o�bV��bVv�hR��q�+�,�5� %t����4K��j��[Ϛ�C{X.��s@{h���C4;��Z��h��7���3����3�)<�X6�3���U+޾,����w�FuYj�ᎇ�%�}F#$�k����N�v���L���ʹ�p©���;�iJ�P:���ew:��љ�3���al����w}��C��W���Pj�W��ѭ�����n��5}X�L�M��V��q恤��<��zx��{*�nK]�ۖ)m)�.ʫ���1#��h]Y���.�5�u�&��|�
[�����)����Gm1�^`2�����t����a�Ώ��!�����G#�E1�o��x���s3.�q�I ��+sF��u��`��ߠ��(�вZ��w�<���I)t�st#�<�̂���H���QJ�`&R��P��������r.2s
-�S�y$G#�h��:�B��M�t.���(*��r����s��7n8�j��z��WJ�,˜�J�9�W�dr����9�X^�W�2��G�Tui��\���fNvzݜH:�TE������DQ��GL9z;��H��$�wE:T��W�+�'����$���pup=9��3����;���·!A��+�*�܋)�W�\���ʕ	$;����Y$�,ȴ��Qy��!�D�8Rt넝йaE!�UV�n�W����ܖz'��Z�Uz�:�IS4Ny&.t�G'"<�Uf[�	Ӝ��Vl��9^��TEA�F����Ћ.�Newg:�B�)�$�DTa����,"�-G]��N�9�Dz�;�t�"������@}Z+;z�K�x����i���=!�����Voc�TC�Sե�V��\�Y���qJ�*D��<�TC�`9*�b����t��N�?����a2g��jǸ)�O��t�^��,�ڱ;.�'o�/I��С���s�OT�Vp��s,���a��W�1�-���爼=��ϻ�`|@��y����f]��'y|����Je���/�:J�/�
��A��[��W�Z�*U�Y�qGʖ�M���|\f�����X�pV��"��5��m�~4)!�7иW��6����SUjW
xxq8Gu�����I�P�*�_��1p��nLp��Du
�vT�\�ҭ��]F��09�@�_^��
NHT��	�������:9@�m���N��t%�h�g���_1Cb��<�񤝷�����1p;�oW�{~�s�y�����Z��C���+ꈻ��	B����]�b1�ܗDr1x�����J:G>ʼ�}��Ď����o���'� �;���XJ0ň�]d�LE�Q&CR1OU��B�p�.����U���髕��q������y��y[�{ʝ�E�l^w���NT��fg�O*��@v���vL�1 �˶���d�	�R��n�k��tj�]%�^�`>��n���on�No/{�wW��ʯ���F,�S�{�����>�-��y����YKx<�����r#�x�};5g�À,t>Sv�66�^UH�|�}<Z69��i��/i�\\��}�W
�]K�g���G�BEuvVm���pL`�k�+��|���V�E����\Oq���Kv�=j�b�?,ʴ�/i�{|5k~�uT��%�j꺌QN��c��[pz�e�	�ݤvJU��w�*a�j.��\�kBِF���eD��q�pV��G3�����Ҹ�uP�3��&d5��ug��M�u���w�!����<E ��Ǐ���Y�O-Հf."�+D��-�u7���4���U/�^y���(���z ��T�Uv��>꧑�m��"�!���}���:��U�����aT%L���s��j��;(�MK%i"8f��B�:�_Ƶf�ϭ����%����{j�>8�v��Y,\!LW�ڡ&+�m��d�"�|��hF�簍����Q��*JK���.s<0��k�kr� *#zXa7��/��t�*ӏ,ỿcq3'���v[����s:q�r���P�����m�a�@��LpӀ(�ܨ�0�/ Y�uWa$���Bѱ&�������k����� r�ti�^�N�f\)�Z�Lm^��ښ��.ʧO���c�vD�*�����m9$٥IIA�f�b,kf�L�qYWW��)��|�ݧ�$b�Y��r`��Y8�n���>�.�7F��B�s=�E��8z�,e��|������O��l�o%l����1T�7��1f��6b����yd�LL}PQ����ו^���t��-�L0#�΢vz}ig�*嚜��E�����,��^�o�����,�&�,n��o�p�(���w�T�;2���>s=B�s��4�J��L��g������8�6~�j%�̂��S�Q��y���~��9�e���i"�u��q:��=Mn��׆ī;�i�gW���%q���ʮ� N�͇W��՛����0��H��H���PJ�b�V�*������1�Z�c3o2�`�'�k�\���:B�ۨb�;'��N�(b��?L�_\�/qu�F�ɟj+{���6{��܊�=>�R��ztB{���Txs��EK���;��� �s�&h	n��95Ir.0�sn�����)ˡ�dC� 'ω��mR���=$�Y�~�$z�n����ؑ@#�a�0�TBN��2��@���?0:��v\u�,H�;>���B�v��yG��ӽI��2�Ժj�1v���W�Eǌ�0~���f�����4kL�{��s�uh��W�{�/�Ǌ](�*�s�{�[�b1k�]�Z��c���ɛ� ��p�+<o��r������N��ϓ��b�����X��(b1",/��x�×BT���� �r�����65�Ӿo��O/pB�e�ՇjB�����ɨ9��Ƌ�b����TCi��)� Ԫ���wV���, �	<b��7/�69��ݨW�O�� �L&i,�bmƆYӔ���Os+��g�EG,���ex�je���L1~4��҇�f��vk�{@5����[YQ++.G9�E�7'�����6r�L`�8^D�!��B9˛�/�Z�SU�;W�������79���UD��o���p�bȼ����D�RX���M.��=X�t�&�v �3GE�)��;5SC�O�g��F�7��{�*����6d��gT�����|�w��|D���K�Q�,U�}��-úa�e�`�U��ggj���%��>=��h��p:�/�����E/��rt?����i�(�l��>9�dl������l�|��Y9 ���g��^����*`������2S�JZ��]wSت�.�4N���*AY�K��J'�9=��ǔ6*qםF�(LkrG1���71k��Z-b���i��=*e��q�W��4��g�ͷ��{�r'�=�s�%w�;�ja,�a��� �t�i��3��J��7qC�wi]��u/\����S��iB%�;c#�(��!	����N�QR�����U<��J��78n�i����:���g��Rg#O�&��	��%q_A���yZ�BE��n�ګwx�nK'�����[L'����qС��*s\��2�"iJ&;or`=ʗ���7�zk]�X'����Rӡῠ��2�zi��\��hE@VX=mހ��@N�U�������Z!d=X�W�:'��H��x*_>׌�5��a�LV�����n�9��rsi��4.��8p�@p�"�����u-����=����X3ͤ����w/:�5�ݗ�e��j�f��y��	%Wyx��+�`t�[��T���~����E�g:{�:�5hfi5+���0Q�z��M�{w <���p�6�i�mp��s�S�!��[�gs����g�r���p0'���1�J��{�!)L�F���b��b!V��j5�M�ܓ��}W�N��/:���>��e�9�4��OiN��H�C�������s���s�QzA�[u�5yo��"��F796]��]���=�d���(����}�� �>�Q�|i���F�2:�{qG%�u���k:�[�O�����7���'|5�݊��Ւ=V�x�Gzx_D�@�^�.�<H'/e��7���-&_<���6��A�h��>���Ȫ�Ō��Q�Ҁ��n_����AG�f���j�nif{�g72R���!��~��<0�,��Q��U}�f1�#�U� �j�m�o1{�"Ҩί!��G�����_W���؎���
���o�_L􅄣M,����u�;�AEi��A��_u଎��+J�{Q�٤c��U���:@��(	��U�B�����Չ*͝�ݹ6ph�s2�_&:Z83�d#�m�|mU���B3aD�:�G`A��W{�y}�� ���L(s+:Y?+u����7�`�=�q��1M������&�K^]w�����Wa�z��&��꺐���1`Hq�͠�],�T��}H^nt�f
3U���l7K��P�ّQʙ�Y �ch�$f+��[.��̤{���7�qS�`�n�Y]cg�V�ܴ���,�@����TC�1���nE ����{�0���+���7Zz�K�;ɧsG��u�|�T1e�"�rtCy`[0�1�l�®y�W5y)��kmJOD�G-5mH�t�y3��8�Y){<�z	I׌�4^
�8�Cg����5z�,Sj���ݻ=S������}G����\��
54���°=G]gV�3ӵ�8�SoO��C�pB�σ�T-;�C�I>��L��K|뮍�VA̋`�.��ԯ�
`}�7�8s!�B�*�nb���]Y�3���"�Xo�1��f�>�×k�aޜ��}�����2���Cd���Lv���,t!L6�I���rA��#h3Y�78��@(�8���|��0¼�zk\�3WP�ݔ�d��o*�4)�h'֫�&�d���vF�<��`�5����f��W�y1�ac��]�����f{�
+�p.iN嶷uE"^�A�_B7�E|ԁ���:`*�DNJ���d�sq�#�㺘/��b۫�t��.�	���nq�{|�������V+�����Z�C�t:��º,޽�����ɇ�l�b�:�쿾\�oi2�����W���(�7F�@8m��e���E׶spw깋,��=S��OTPV2[?\6������b��T7�Y��!�y822V������X����� \5�]e�K�W�=,`�z%����ɢpVY_KƗs׻ܰu��,Lq�d)��&#]D���*�n0�+r"t}�U��y�W=�Wj�'O:0ꆍ�\�P k��(�Ux�Mdi�:��RÅ�AKb_��~����u
��t���	����=[�la�#�o��`��ol��$2�/z*����ܭ�]$���{BXn=km�w(�s�8/��bo$��}�,�=��Q�'��:d��g�8����y���"�H<�t48n`�R��éf�^��u�}�_r��9x_��r���l#��ݎ|��� ���������gG�h��>��
ïv�7�=n�Δ͗1�8_��Y�~�D�3�hƩV�*��o6�Յ����˜�	S��ʕ�8C��<#��*s�)���3����4�-^�WF����'Lk�<�;�"�1#��,n�Co�4>�I:�rTWH���1PX�!f��z��2��^��/i�T���V�����¼�k�\�S	Mc�y�w�k.u=��$Y�/�\�@�(��TO�T�*��ry�ҺV�x.f��4ey?_2u*�����js����QG�%����:ٳ+�\.R^d��w_�q[Ż�Z19ލ7[{����2�6�1˨l�ĦP<i�u�p�V��G	�������%�`���ʫkblEٱ6\f��7�(��p�W�&��q��7b�r�Y8i����*΁�:5t3�d��O��W,���c�h�鞮�<�����>�����`�1Q��g�^��O�>5A8\̻w���[T��1p<�i��5v�$y�]V���n��fݕt��y��>On��kw��\�J�EU��ZU������v��vF�� j_�CT4�8;շmt�m�%�T�`N�04W���:X(�=�������@\,Ϧ�sE#Q����ܨuu���X=�V����N6���c����|47ʀk�Gn�=�	�Cҭ��������a]��K����BM�m�K1��
{�nH���	��΁�n����ye��,�xዹ^�mf���p�c�L'M�1�z�˅?'��ǥpTm�)�1k��;q�.���E�
J9u~X��\��Vxhڄ��c�)�p!�b��rP�q�EYy�&���ycSѿt����Ұ�0���a\=W��9�G��{\T�]�d؈��#�Z�`�k\��b�	0c���LM�J����v�ceM�;��T����\ͻ�Y�c�Y+���K��
���^30׆d�.�S��xg2ޗC�(�'Đ�sn��ws}��S�Ƞ+�e��Kdk�爼=����d]E���FB��h)���:o�7��zm^�fj�i^������G����:rvOm"�=��&jt�f�x78��Ƌ���#Ws� ��gr%'+���ەƯ[c;��O�Q�yӂ�/jj^Nv	(�d�xl�nؐ6�yݞ�����i���.�v��fl��eC�y8r�2�������W�
��8k�[��q�5���GX�u/8�˧��E�J���ô�3놦
0�D���<����� �5%q�m���y��Vw!3c��õ8(F"���p '��CV�h��F�����{a�[yS8:#=�j���|���� UQq&ʜ�B���#��J`�����/;��i�W��i[��R.~��pV�-�G������<����kC���R&Qn��9�]�W�����Ӑ�K�Gk�Oˤу+���Ԉ��\,�Ώ?��^�U�g$�O"�;�����W�ta8ԭ��0�ˇ_-5�l=u�<4�7�)���&Qu�`��4��o;
����'\�[ �����e#�Cɍ���U@G�$	�Q; C1m��x���*���[�S˺�'/���PB*UHv�<��Ќ�p*�~��6�O�ƾ`�K��ǖէ�S��{K�_OQe���T��	�4�G�Z���V�E�����8�G�^�HEn>�|�.P��4}#zu��ТYX%>k:��:��9:�:����:��즥 ��2�C����ua+ޫ�er{��w �ҙ(K�H��%� �l�un�m�;2R)C��ʖ��t$�[і�H�<D�쮈��1Jqs�(5B��k��|û��p'�d��nb܎KV%Zu�'�S�Um�Mk��t�1Y�Ḁ���i0�ۥQd���7ب��t��K�,}�Y�N_x�,Iǽ�$=�7��%s.sq_v(��i�_wq8 �m�av<
�j�i%h��ޝK��s��D����îa�)��*\F��&�د����հo�>�Ik�.���"�>P��M%ژk}k��[�0Q��\��%<���W�[�,W��
�ٴ�N/��4+�"R%n��T�\zf�V������U]h�{V��l%I�	vo�9���F��+n�8�a���:s�^*t��A�a��1/d���.�f5���S70/�����BN��;\�z�m[-����1]��(�mD���İ��Mx:�19*�z�Rh̲R�G
�h������*-*�e���<o�.��K�n�R�֔-C}�t]���pZ��V-�X�.�������:���I��Z�7��w0əʡ��B�]�����3����Z.�G�d_;�E�ǵ6�К��Z�z��A}6�:�6�b����;�ڊ��떩����z,A%:"�4���%H�'�\��9��}����Az�O�0{��[�^IN��oF7��G ��q�;��'/6I�9��p�RV��Q^��P��z
|�⥋*��~dh���RU��^3���w�ߡ�v�ɻF�~���=s(]��?*�	Lo�}C�Tݮ�Y���t�22���[YWjΜ�G���r�(q۹�\0trUͣ�V��7s��9G��f1/U6�.��,
�e7��A =]ٛٸ�R��11��0�k��]��";�`���P�7I�#toNۚ���^���9�xw���������d�±h&�Auϥ����9ENU��*�V)v0��'��eݽ��H��Ύ"�^�պ����#$|��bV1jN�4��`�y�8e����:���g��CID��7����c=�Ug�K��{�#����O�/N�}�pʀT��[t��g]l���QAfi�����i��nlV�����w6��ŃR+�!�j���K/7*��i�����b�R���0���	�mm��{de17��N�N�ƪryz�,e��Z=���d�9��93~N#\Q��<�=>_:˨�J6���i ���}(��<gt��S<ʣ��	ƋT�
����l�̹�Yѭ\��cj�N�}��iC %uq�&�9���X��@`��y��!1'�ݜV��"-<ﳦ����u�����xnm��/u��n⺔{9+�ۑ�{#�M��NഖM���"��:���Ξ���#J~������Py�ߥ�N�7X�
@�H'�	Kd2WQ3�H�����3�)�uhfs7$�xZ���&棞:ք�d-B�GH�(�Cd�R0�s�w�.r�@iQ����2�j�k����+5%V�QiTC��8DK�)��pّ�+2Cr	�+��]�<�1�e�,�U�**����[�Nf�z�����Q̊)��wuZEx��)�]U�U�⫛�6wM(,�]���"�9�!�r!�S<�D������s$��D�"{�z)����T�<ÄTN�r��c�UE�PB �rp�qݚ�s��B��5�E�TU̐�U�x:	c���T�̨(��j	��t!��*���S�+E����wJ�D�	��G���U9z�<*$�B+���%�	���u�3�˨)��TUJ�PS�VP�y�AQ]$"֕ȳ�U��I�)VN`�,��NHQ�
�ng��U\*��4��a�	I�'�jP�Ls��E�"�9p���n��	��i��I
��ܬ�)P�]�'t�����������J'N���=�����[<�-��\���=���cV��Q�y卾hގ���e'����o�iC맖����:��H�#J�3'f��Ϋ\!�� �����|��ߙ�S
�쉾�]ɿ�������Sט��<�&�G�~C�}C�C�ߎ7�C�?!����a�c�O���]�4��$����y~��ia�����2�ծ�J�P.>!�(rr��_ݤ��N�v�����˼;N�������0��V9$?;�7��W��}N���Ǉ˂w���=��������9�P��C�{v��lG� ���ڴݧ�fm�R�ƃ?_���nO�=�0~=�����Ss���w�yM�	9���������i_'�޼�7!8�<c��-�'�9��@����G�v]�7�/��n��%q@}I�
���|��5�"����+����Cˏ/&���������ɽ��GtS
���ӓ~Bp{���?�����q���ݷ���:w������������r�M}���ׄ��O�n��(���� }/�o����˓�w_޽C���v�zg)����p?�����8��>���ݷ�>��hz����90���߱��n|��a}�߼x���?��x��x} ,���_}x.����y��>�"��"7Q�|�[b���@�շ��wTz"(#�"�Q�#������yW&�>����i���=��H&�����&���v��x��\��?&�x�\O��aw��{o	!�ܩ�����<��M�>_E���>=Ṧ��=��[�C}>���H� �D_O�	<8����=#s�!�܇���{��U7������!Ʌ����xAw�v܇�?'&����Cϋ)��8�_7Ϟ<?�$ߐ����o.<�>�|O	.{���j^�_�����z^� ��'����ρw�i7�/??y�w�p.���!����N9C�&�O~=��0��o�_�?|��aWyǨ?��o�$�����r�z?�����#� ���Bq�:1_�Z�|��D|P��~����U�S^�s���oI��۷����=$�����|���nӏ_o�<';{y]�������s�x������Ǐq�0��A��o��xpz5��H���7��3�^��|��~=v���������99����w�}C������0��I�~���|C�a|��~�����i��������}��n����C�ɮ��x�����#��}Q5N����#�(J��El��ٕu�H˙Ԇ�%Z�\�l������l��!F{�v
�)9[8d��/R�mԚ~��N������tM���β-��}�N;j�UD�W���'hE�,nP�8;:��Z���/��.4�p�񒌌�J2칛��zV}��$Dh��q��P��GϜ~v���'�~C�aM��>��~ON?8�@���yC����o�ϻ����|w!�~���������������8<�/��?r!�z�~}��}7(�}[~=���DH����?Dh�!Cˏ��������o�=o��m�����7��^����6����>�{w��'���1�ﾱ-�
���^ߞ�z���|������ra}�S�{BC�F_����<'�6��'i�<������HI��!�5�ǝ����O�=w��_`���<��|㝿3�����O�DP�>�	��.��p�;�_n�rG帍����}��mƳA#�6��x���PS�}|;�{�90�����0�PNO���㓐���s�;��7���ﴘ\|qx�����#} xW�-��r�}Ƨ��^j�<}�����ǥw�ӏ��vS�SO������=&��������&<�������x�!�'N>�N��$��r����P�G���������B#���@SXv��I��Pe�����e�G��"(}"=��E�� ��/>7�zC�}C����>�H.��M޷�� )�7�y��׏�ޓxBt��~�yIM�<��'���x},�����R�}���\�Vj���+��{߿�����w�o�s�T�п��;�?���`���C������aw�.��|�8?w����$�����᝿����?�xǤI����;��7&�<�>�GǏ�s:k����$�6����ϟ�C�a��yq����?y�Ǆ]�������P���w��e7�'�ǟ�x����	����뷯��0���n��ߟ����7 (���?y��#�DD,��M������'yƚ�P~�x��}����;ӎNO��;�!��޼^��\{O>���nC��=��<��&��=v>��?&���=�<&����O�8|�$�P��c�7��/���}c�>�(G�J=��o��kԗ�ħ'=�}�DE����#�"������Ï�'���o~C�s�i���<�}C�y�����}X��{Os���Ă�w�=��Ǥ�&������v���<�������I���ힺ坒fg�3�����s��n:׵�#����C{�f5�0��L^;�y5ۃI��g�׉�a
�e�GX�/2�͵8@����Gn���<��&�7=�=�:�BU�֡Y�u�J�ڡ�힫�w9��Y�N�y��3��K #��IP�0�0ۛ~�����zM ~I�;�����i�bC���\Aɾ�{��OAׇӂC��'��i�<�}}�=�S~�;|t���M�>O��������~���O�O�)�_o���т"Dy)�>��o�������I��|I�]���}��ɽ!�0�Q��'�=&�{�
r.�ޜy7���|v�y��|�A>��0}DC��1怆��r9��Z�D`����P�#�q��|Y7�ü'����\����_���_ɿ�����C�}C���'{߿x1���ry�����U'���1�9�9����r��4 ~Ii��y���}�z��L�{7Jyڄ��G�"�B=�<y��ۼ��;���ps�G�o���G��7�}v�C���}�zTߐ���yO��=��~~����S�~����]�g{��Ohra���^�=�f�jZ��J�z�������`9߷�n�� �����a@��oI��xO/�&�����Ï
�@���s����c������C�i��{��_��.�������<����W}q�&�����#���S>���gv��`� ��>�o�}�����raO_��i���9�8���I���-�0�����>>\rԝ�z�<;����z?�xL*�Lc�#�5w�<>�|~c�| ��ث���w����} D��C�>���8<�����x��U����?~��_n	��s;w���Ν�����>�/)�\���w���C��䈄!��1�g�s#��>���]8�F/C�8&��Z9��{���#} c�O�zC�~������������\y@���O��}x>;zM�	���'�p)�����ӵ����:���ӧ�τ�����I<y���!(��wt`ꢦ�^��Ǯ�{k���G�F��?o���=8$9�����ߝ�=&~E?;���P������oΐ��������Ă�����v��$�۽�xN~;ro��(�Nҿ'�ֆ"(}}r?,zDxoM�yuy(�a�?��M�t|O�iI�<����r��97!{�����O���y���Ϥ�S�ra��?x�o���A����U��'<��yL/�o[�z�"<(}"!�4�T��^�0��] �WPOV��=0+���ѯ3ٟ�{����f�)�-Q�`�f�5�^�ұv!'�W�O{��m��/\��3r�C.OrJEI���kE�����ݲzr�kK�7����BW;`__;h�g2�s�S�����n��M��u�90����;�or��~��n��n���xE��;�����7�$���oJ�Syw��9~;~N~�$��?&��v��ǣ��xǗ�ǌ|��v �V��@��F�|䥾/_���L*�����}gyL/��F^C�}C��9�raw�~O{�yO�r�_4�I�Hs��[s��9]�������H~q�~��_��ۓ}Dgߢ�¾�H��
�Nƭ����q��{��Er�!#�|d�������N>>����?���O'���?;���Bq&���'����!�i�O]�Γ�aw����㼡�<��={�ʛ�=���|�<�����_��܏].oew����DCG��:��#�?��3~���_n�>�}BI~�z�P����?'���]!�u�ߐ��|O'^�����='�o���=A���xNv�㼟��ql�i�ڎW���}b>�">�1��~xWoi;���e	��q���?'�rzq��߾�<�N�������{P�U�o���7!ɼ��x';w�=����ԑv��漻I��'��߽��{+}>;��g��X\y���p`� ���rl�<B�>�t�����!D`����\?n������r��9	��U�G|8@f�`k3�$EEr֏`k���Q���R���2?�<0�:*���k5.�{�1�^kM�s��"pbwj�ӹ�{4�1�n�[���.	È�b�B�����BLֽͭ<�(�S�^K�}6%���&]���3�G�{���UR�s�ypv}�6��M^��6Z�Bc:-�9�5��2��E{��c=����q.qFe�iq?���;Y�=Md������8���䇗��� 6�D��>��׷/%�Ȍ�nލ�R�ɥݠL���� �����Ӡ�e�J�y��Ռ>���3v��ߴY���i�8����^����|O��y�#Ua�t����\��ţ����F򆶯vc���.$�ˆ���3,�u�#Q�P�p�(���@p;�T����.���!�.���2v3*)����9���V��7)���ɍ�q���P��x�\ʘ
�_K�v�C�P4O���<��YU!�4��Z6:5�Eq�^��Rw�X�����b��OԵ�Gқ@
фʞ[�ۚ�R�碃MW��q=�M��iVu)����ɼ�q��g��wD��޳N����&�zJ�u��Ё�;���2=�Իp���q�ԁ���J6*�n�������A[O	�̜��Y�ڶ����}A�ƣ��&j �����@Qn�_�52��0Pc���w�ݚ�ll����W)7�F���,)1?l7��f�rzVPm��<�i/䫴�N�c`��]"p�֧uNw^��_]r*\���A�m��bcyK51�3�d�PuI$E_%Ef�^c��D�4��mDMTwdŅ�,l���'�Pw��b���+��	1�//��h8Պ&!F�ų�Ԫ�+���]����4a��:�//�b���ދ�1ne���t�n�S֖�Q�&^eaݽ���vԗg�Go��358�+ɔ����۫�>�jѤÑ(���`��v+K�^�gF�}ׯ��%��N�v�|��?��e�}�ٔ�iȱ���Wf��z�Ug��u�����W|HZ��^i4�Kۿu[8��F{�*B����pk�΁���rzo�k�;������nE���\��yZ����B��ʴa����\f�܀���'�Y�J�����`��-
�������k��NPuZߔ���ׄ�������\H�7���ё98�]�B8YJ���	�\��c��}��/�J����/e3�W����_ϮO�u��]��I��3�ڽxڭK�"x�4
uZ����W�WX֎���@�n?x�>�����\GY�wQ�ՙ��Sv{(��vW?s�?;��U
�M�5�@��v�uQ��\P�=,`���u�O�m������7e���]�C��6ԅSPLF���@?JU��enD����{X٣��QFzigv%W���[�c ����0O��\!���p� �)s����)i0���G���-V鉶��S�(о���K��܁���n�H�ꠅ �v&
	L��i�R~�������2yo�y��h�`��i�l�u�8�j�e��$��n%�%M���F=��Rk}��ǩ�vr��kL|��%��5��Z���j�t{F��߲�4����=���ve�ʞ�c��p4%�ᶪ�F���õ�����3n$z��_�c�ә-��TP8[,���|�s
�tD�*�$ن�ky�Q�֩\�"ba�E�&b�a�\���$��T��]c����U�C/y���͓;ӈ�F��'�����(���^&��t��^��t���%'V��o0SNy���{�!B��ޯP|��h.�/a��v��?m��8�+i����S�%;��k!�N�dB�P���� ��5�u�F�7���k��؎����.���lt�X/꺍�={��Ù,������U	���(�Zp�+����2�>f��վJ��c7����qX}3gLD��;���G�Q��Cog�o(�jI1�E�և7pr�����QBBr����8��~C<���79ׅmW�]����績J��v�f�e��R��T4�C٬��ڄgXx��8��܌�W��;5SC�O�VE�M�z�d�v���'����N_{��e�r�¹"�W�BΤ'�|R������,=Hf��(�[�Ձij�F��P�=Y\3;M��}l�O.4���H�Aց�.x+c�Fsk���.����VjE�I�8��U��e����l�Z�:�>eK��c�v��t�8X��Ks���O�9FohZ����u��l��Pv�\-CC��|E�~>��"��Cq��9T�c>��W���B	I��bu� "����v�V��)x�PK#uD�q�_Te��<�v|��j��
���+܀Z�*��)L������4�E�s���䕷^�������ח���Di��ӌ��[�fQH!@��6��N��/6֧���У��}(4b�l��	R*���#�{�_��W��B�B��׺t�z�23+Z��[ ����F��.Ŋ1�w6�V�_�P�5��Ra��ܼ�ᚧ-N���;}R��j�DӔLu�+��1�n�1CC��J�|ep�ڒ��uW���{�G}�����i1V �s����d_Y�a���\v�@Zj-���]�Ab�m������zcrCn��Zie��q{��\7�l���(X��C�w����_p���F����}~�B[�3mos��2[�l�9�	�
���bϷ҉�Xk�kI1<���|�4�c�Q�{�AV�6JwO��p��;�Fk%�2k��A�wl50Q��&p�7�p��8I�ًd\�2{%�۩��m��Gu���ئ��ǰ��W��^ᵗ��bQ�Xߪ���JZ ^��(?\�cw�Z�y*�n�=�M�[�����]�HE��;�!�3~���O&v5up�q'���U]"�N'�b)��:�����7!��^�$+����g���GUwcj4��� }��F*K����.pP��,��� +��yb��B/��O�C�˾�5�z��.��fN������3 ��y8*Z�ŵ�G��;|��9�������nSy�s�R��𓡺��Z�H��{�[�+݁�G�s����j����gÀ՚��Pf��j|���}Ct�/�=�	�]�6���:a<!��Ώ:���3�>�䅾�<�8W)3��U}�ĕF2�s��>}0����ۦ��.!�R�����&+Y���}Jp:|{q��X�Ts��F���D� �K=�s��C���ڪ+f�3ncVYF�a�N�����cv� Q(��&PS����腕R�N�w���!��i���۬�
aE\tV�8-K3^�w��q^R8��m	:�yw��䰈��΍�W���f�F&�R���J[S1Sǆ"F8�o!�<�Gˎ�.5�4V���/��4 ��j����jszĲ8Ɖ+�q�O�.1�G�l��ʇB���	��Ѡ�ױ���"du�������!�Դ-u!�:�^�V�H�c�Adc7h�VžwIKQ?��X�o���޿�֧����kx�H�M��}�����3�VR�AWJB�=�����_��u��K9}(��Mq��nˍJ ����w[}ͪ���AW��UWե�t�$о�;x'��W�&a3PZ���$��]#_�|Ն��+�>�Fb�k]�k�׸v"�_��a�/��pl*<5	1_T7���\�.ND��:ἰ*-���2��5n��&��ֺwTT\�jxEi!?�v��g7��7�Te|�[��c秢T�e������7[vw�#����q/jƇ����e�k@C���Ud��10��T��E�x�}Ľhu�|�ߺ�pX�^�y!��o����b�,�1	3�ʒ�{6v���sQ�#�d���jP#��*�`{A8^|�i���]fU�_��@D:u�%G�a�5���11�����5W2�e/����tG��ڥk�����'����{y�yQ�cݥgDE���\�t�P0Z;��w�
���E[ʍ	e�F�u�m$Q�����
dE\����1��c�s��#y�2��o�ҧf�����m���:��e����4�Rb�B���$�J'�((�����MQ�'T�6���f=f
��c9a��}1��?w7��a�\�ݱ�؉,i�����5v95攖�y��y?V�ѲDgMO�n�d]֛�BT�av����M4%,z9u�Q�}D5�l�or��Ҟ��uj���f��6�ۚ`��d�S�9��ŷR<����|���]�'3�z:��O�=�{���{&-$���c��jF���{sL��u��U�9)k�B�uN��	"�h�|��VX�'>��c��kK[�e�f�B�Rҡ�{�>��V����?�'�[Ho]��I༗��=zOR�k�g��� ��Yκ�i2�ț�vq��c�\�f�����!'����C��s�u�nj��֦���`�+"��O[��ע/�%I�(�+v��gQ��~K)<�����Kǈj�,Qr�^Q��e��_��HG�9�y4�ءL�q~�	�ϸ���q=W�V\N�X�X�.�!Q%7�s�^��_Cyi�
�w)7��2��-�J�^mZ]Y��m��ǽ6�X�mkޠ�VZuz ���>;�2����޾����|E#3@�9�j{�*�䫺��T�&�N��Nmî�cpڵ� �q���m�ysc���r�>�%�6���XÛ�V�,��-#s\0�+b��\�ݸ���vF=w��*�Z���:���*,1L��5�2�+��M�R���ckGQ����Tş>xu�]�����9g�%qm:c�8U�7\te)O��9��쨇�T�;��K)����JZ�����#e���+a�Cz,�۱p�i�5�v�.�Ә� ����Z��ZW)PM0Ep**Y�4ʺ�*��>S� �W�(Ý�v�)�X�vT�)$`�X�ͻ�,�MeX��ւ'��8��g�T)(�}�u�.��n�e������O[&�(�&,��͝�Т0�}E�=;��-���G�����M��JUf���|�G]�ބ�[\�|@�e�j��R��I���Sv�N�V3�V�Y4-���R�ꛁ+n;J��e`���t$꽮�.쀶�+4�d���"tb�Cb��w �4��S���J�i�ћSYAi�	��M#'c�~kfȉ����)m(bVi����s���K�2 ��h�wR�����"���ms��A�E��q�t�Ñe_
�\"Cu4���1mYz[�<gt�Z�`?-^74w"%��o�ra$e�R�!�ݱ�!��ٸ��vj"U����e�5��R.��d_�+Xf����Ц#w�r�8V��T��`���AnO�6��%�%KEo=dhR)&�*�B��Ӟ�|M��F�)�6U���c��t|�v���Ύ�勌���^n�r5�%��y���@I�u�d�Υ!�l��m^9�%,;ك=զ���w��[O�(��1[�;��6�Ӥ�j�I�^`�]�5y�ڤc0�zt���~G��%xB�(�����[��Ve!a�YժЂ �J��z;�t��@���2wٺ�r��pD�:H��*���#�R�8��Ku�2�0��H[0�J*��ML̕I2�QR�.��tH�<-���1�Ȍu�T;���P�S��N���t̬�B�Z���@�"�D�%�.H�IeQ*��#����t���(s ���<����9:�Hx�)��N�ZE�zR(�qE��M����H�Uy�a٩�kK֑EP�'6K*�����$����GM�rʌ70�ʣ�0��YW
�wK�"��2=B��%u�<�U"wp"�r5+�s\�9Q)$V�(�P�t�#C�t=�ֳ�O]ih#���I�s'"ʬ�GP���u�.G�.�s,�(ڡ9�y9�K1%ø������{$��,��d?�aJ��&5����ͬ�����\%s�������Y:�*�G�g#.^�L�w�lխ�%0ul�X�<��2:��}	x�{��(�����5�#<���
��u�"t� ����kt��g.���Q�-\sO3���C���M�������ޞ ��3~��d��ϟ���_ػ�m�Ѹ�Srگ�L�\��4u]����ۇ�@N�pX���)��bo��* �Y�8k��Kի}@�h;����{�p��l�ި�j�O���GS�#������E'U+�@峛�{p�r��z��%�|t'��H�.y�v��i3o[���:S7�h�܌*�ǖA�A�����Y6��O\9��-��c�J��鰄�W����n��;��9�s
g��u���t滝d�<��e����T�h���v ptp��גS�3�{qP� ȳ�R(S>p��++�fuPJrLX��昞�zk�E��c��uײ`���F�����ۡa�>�ld3"������s��`�
bO�3c���v��/��[�J���NU��H��f�/�-��e��E�+�Q�&����&8\�Kì�G�G��o�c�y#+yᤱ�K��s󥜱,at��S��Pb�/g8T��4:�^�u�M}���Gi�~~޶@����{�f�jp����1֥�t�4R�s�;Z�u�����Hq\�$��'*�h�`.�kYݢ�V�b��C�NX����睊87�_�c�ci��M�icׅ���o:b&���N�%�_��_T6��E#7��=�.��:�M��g1�V]+�=��[s�.���򗫀��gHb*M���7]��J�Q0�ʜ�S���#��r��O��0�G¯eR�}��ZU��3��U��e��4M�[�].��Z��`�S��qWy�U9�4��q����x��x8��i}��n�L�F��0���U|��	�f�|s�n�u,oB���\7��vFȞ��J	M���:�m��h ��[ZՅ\;Nd�..O>��5K�q�y�wLhJ�]���d�@-�g�0uו�e���{��_�Ԩ	S#�Yh���ơ/uÄ��O�v��r�T9�lgNQE"*Zb3� ��am�m�]�ՠR�4=GWPh�|�H�S�D�$�6cV*L柰nrnkKT�TP":��rΫ\�z�%�` �T_GϩR]�رF<nka(z��1�𭴱��s���\��UOs8�[���pU><MnU
=�"�[����R��W�S���>`5Ү���`ܜa��IK�da-�#O_��o�F�NҳT5���S�25�K"�u�1��uà����ǶP�E��gF�<j��S�g��]*NFee�b�f�\oT=�Ih[Ǚ9��s9)�h��S˭�
�eZ�OO��<��z]y��'�wq��>����7s��-�S����Ub,k�@�u�*����2�p��W$Ó�R��Љuߧ����{��g۵WK��p���"a�)�o����e u|�"���a��3���٫`b����˿iv�FGT��vk�r��T�5J�B�D��%���NWj�p9�d�B����l�N9�A
�H`�T��8��v�aI����{�?��_��*t�7�p����Ie�T��X�9��+�#l�p4@�}_�����U�
Q�X2p 2;��1��m��1�&&q׀�:wn��<G��L?V�!����p�slYzP�'"=���5E7	7zwk�s�]�x�RFnJ4���/�lM��N�!�Ι����
�>�A��[��>I��f�o&)w}���}V�2P�G3y_����!����
�δ�D�y8�����z�Y�Ö�g���0��YP9����W˹�G~��/��l����=�l�#���7Ջ�w�7|/z�����7et�K�1q�9���V���L�P�cq�5{��
U�/���b��;���l�Ɵ$����ro�����Δ����)�f�x��v&o�^*0��/��Bnʥb�zQ˞t���������a.���eje���a�Y�9��^��fd��ݛ�%�^�B�kN5������5qō�����UU|nw��:qذ(W�R��L�(�96x!�U!�n�w �69��ע���[�ry�2n��.;�����#(�|�'z�a!�R�.�{�u"%���h����o���i�>�<�$��� ���!�ѯ�� l����t��޼�݋r+��UJ}��6�ӈ��P�N�9�Td
zdء�|�$Y\��*��zOnA<�c�ɋ�˲��;��5��QNf9��yZ�{� �"��Z�|��h�++xGUβ��,�p!C���s�wN@!aI��[J�s:�I��H_��&�@�C!�yn�L�p�aq�O�`�Hv/��ynN����W�S717?>/x*=P��I���}z�M��<22Ox����#Z1��U�����5�&4 �9U��=�9̺7�4��՚���L8Ǯ�n����A�=a}��a��g���5��7�pj�N8Ywk��<� q����uR�N|���t����M��%�r,u�e�_�:���F�����Gg>�7IK�z��o4Y�Z�n��0à�&���CӼs`��WfI�#���QS�k���ij�Lm!�ǈA�9vd�b�XxfIgp�����AZpn����q)F���|/k�X�\@�=6��wTH������簻YMI�p�����o' '��
��`�;e/��zX��Bp��;{p�bi�f������wZ�a��ڽn7��l`�w[��>����hɗ�5��̨�+�OE"��d�8Y#Ջ!�:5����K<�g!ƙ�?�Wj����j3;=]#�Ӓ�������0T�Z��o�QW��Iw�=�|~ɵ�ԇ�>��3�ڊ�⋆b��-�2e�2<>*�K˯A1��/����Uå�[��נ(��	�Yκ�(��8A�C���
ˈO���'!�?���5�P+��>x�z����-Ÿ�!f;�O�;{p���B�%���`h���袠��$Z�NN+�AE�}�~p;OW=��ꂊ��O�
]w���q�8.T�M�A	dU���.�qn]�ƺ��H
���,uE�H������;�u&Z�j�	��`��¢�N[Ɇ�l�KR��%H�}�Q"k�9A�;�u�:�x`�.{p�/Rv�gΩ[��T���^���{|iS��=��M�b�i��1|F�&nT�Y��C��S�7Y�7�ަH[-�{0<Ygn��L�ٲ��v���w@Q�|�@M��]öqYk.;�:�39�U��5�S��2�T�����9C��==:��|��J���U}�}V�^�KǙ��J��zJ.r~GI�G���G�C�iv�BR�����޷�R��׳m>#L�)ַ�+bD �9UѸjCrDP :�>���O��R��e�����E�װo���#�JW���q�*׳&�ށ�N2!Ԁ����c	� O�	<b��7/���q��^v0I�K�v"�����/�1��T&W,�aC��C0�`؆�¹6_�a��yg��ч�����(�Q�ԍh�k���X�L<=�J�UJ��Jy	�j(�nO�{?`$�P'�0&�9u"���FˍRI�_NSq�B:���gs�������>6j�]b�u�O�`
Z�t]��gï�%�3����0�G¯gʸEQ;<%ZU���v��O#s���*Sw�<�%y�w@8�t��;�p�_�kl��R7&���̮�ګ�:��.͖��ղ���n��������wLk���J������B��њ�'B�]��]{��2����LE�S�>{�}V�y�8�w���>�6p�VȬ���w��ZZ�>f��{�#hT�ʝRH���Y̙��{u�޳Ӯ�ѐ֨�ե��3�'�%2��3ϝ��7�T�l��u�d��;|$޹>ʌ�B{�w=��Nd���4�6���˹b��3+4�x�.S��k��RFLz-GߘU}�o�����R@._�g@Op�P�)�x���2S���ne�4�	��wr����fVnOt$��l!��������A�q�]��u�F�;H�G8T�׏�&�\�uy۩ed���q�=y]y�q"���%7Ԩ%�=�>�UfDl��u}2L^d��n:�r�Ş��R�8'n><��Ճ=t��4�q5�Q�9*�E�ճ��a=��J��RHu��t[�{�Â��+<��@W�2�\�"�\r����`�l1�QNT�K�캍֜�V/Qxc���ٸB/�LN�������� ��d\'$@��o=�Q1���b�O�B�}�D:�[&��.��1���Rejvl�j�h�Ϊ�|��R�B�a�KN5���i3:#E@��TE�|��fk%35҃�O�w�`#L��L����܏�Gϴ�)��3��뫷I�<���C1J����2?���W�z�>���W���-}��}<k����dL;���p�� ����պ���f���.���sYD������+p�%�@��b�6<�!ƍb��a��:�7[����4^�NKu
��0��mȅ���嗌뺳�J'Suݏ�����9q���3��";�8y[��4r/��8���򹊕rT��n����E֍����s��J�!@��ȨJr��i�,؋o�X�}�}��0�no=���<pV)"�:��2����_�)n
�mh��%��+�.��]G�$5풮x{;����(j��jGg:d�1l��'|"�j놇�������A�	�^&P9�9�ȹ�)go#j�vc8�p9��*�b�OJ}0��n��(!�~{�x�����f�Y���;ԣ����qU�L^����n,��Mp
�)����cDNn�]4���I���V5A�^HƢv@�J���ro'��fCi����h��)m���EwNsk��vѐOq�+Ke�/�lU³��8q�>m?��K�Y[������Mo�u���.��V,8��[���j��m���|�`w]7�ӣ�}f�_M*g�<V{UƤ�\����3�n��yq�E*u�[�@��@�Aҙ�3p�c7��T{�CW/`�Ƚi���Xp�Gw��������	��s���(�H�'g����Z��-���)j�����"4h��=;�3�S;�$�}M�C�E�������{�Q�x�sŭt�K���O�c�t}��}����k�v���y�n�+;]+�^�i]��%�<wsZ�����ӄk��W%�����%ۣz��Uf�w���痐�)�VOL�������m�h8yefQ�">�����4��Z#���ɺB-��c��7������T*�R�s*�8�=7c<b>[=�:ӶG� �P{D��咴��5P����X�4�D�����Z�������Z�Q�bZ|�c�zQhP�e}�e"��ȁ��3X����k+�[��{��/����v�nnlWQ��Pa|����u�tŏz[�6#�JK��X묳�q���JY:�v�t��ꤲ���z�ʹ ��"G'P��j��oL��1���B~���_E�8���u�i��H�S�.#+n�{�1�.�n4�KL�t:�����gs&ˤ���%�9,���!i6lC��VN9��B05�א���{N����vƜ\����?��Dmԁ���g#|��88����Z:-t�Pћ��'�� �⤫�v�Ο�Ѻ�;��ʃ�m�/�`C� �r�B��=��*�.�hZ�}��m�T�މ�ZpzX�=���7,j��
�	�ciHU Dk?(���wR5wF�i�Ht1���:nj��Y�֛�!b��]!�l70�U
���Jb����l�V�&��[�)g7wIx�H�5e��G�	/vow���j�ϒ�j�_����jNP�>^*gWF]�^�6e�Ӻ"�z�Oy
�7�6�`���dD]��_UU}U���y����N@ �櫶_�{Qoj��8^(��u�#B�uY�(��B�T`imS��G:��r��@F��(+��]pQ��?"��7 G#��t�C�@c�v1'��eo"��/�EGG:��y{MJ�l����nb�N�f���&�S�10%�3:k���֧/��<�w,�s.H��0k}q�/�x@<v�5��w���q�C�L�5Mr��ګ��N�K1�7v���%��Xw_m~H1S�3�xf3v\<og9��{�J7�w��b�M�W�s�gJ��ܘ�9�>������|v��\en����5�Y�M�H<����V��IqxGMC�cE�L\#"��D��<�>8�K��B��q�"�g-2R����[��6���y�PSf+*6�e���K pB073��p��8X��̫��v�KQ�H~���DxU9����ٳ���g#�A��p�ֲ�l�5�s�s2�3Pr�����ľ��f��"MXc�E�V�\��k��ٗ�g���\��^*��w�]����Ԯ�-�yg!�6�vG�3Z��}��W�Ry�N��
��Y{Cky���F����ա�R� ��T �b��.�'[X�0mE�V��`��Q+�=�}nz����a�3�S���;�<�s鬞��6nRD���kNҲ0�mK�Zo]�l��'��^P[A�7>�Y�ܕ���bÍ�F��]�Y�`b*�-֪_\�F)�U���3V����ZW�뤚ܬ��[1�����;��w��2�n��}��+ڮ����Q�%�y,霫3�;ݹ6l��8�95�cO1l�|^��K�t</�*����0j�Y޴)�佒K�e�`^Hv���kGsF�^і�9ab=Q&�^=ٽ�ŽM^��k`G-+;��Kuk!{<j�m���j���/'^�2t�o��x���(�V���i|�K/PQ��鬡����s�u���Cf�=Zc^S�޵u��*��J��[z�[�����IYk��WU��a�uL6A�c�������妷����9�cm7��&R7�&�"���*`,�}�3_w�A�ǹ����M�r�i�T\C�\}wwiՄ���w;��lW%�5?|�Xy�^�p[���;
�.u}�Ƶ�ޝ����%Cu��@��@ť\b�e��(�h���Gz�P��@�q�������R�c(��vd0���0Ȋ�n�kQ�io�߽a'={M��)v���&�����m~��du���X�(�;�Tr�,K
tq*Ǹa	���J�h�ls5|��fM�]ꢃ���z5���~PY��;k�E}�0H,Dh�I�-����R�4¡m:eT!n����(�5O�Ǻ��t��v��kh6��D�.����:$��c��WV�ow	rc}���I�G��5�+י��x=b_�`�R�SpÌ1�&-	����zT�3��X��h]<+\���!h�Q�J�<�a�j�;�����,t���{p�D}����MM��7��8�Z_(7ޓ��foyȭG�wJ�5��E!_�xo���%Z��rM�-�M�{KZrf9�ò�0�hT�����������ܝep�wy�"�E�v��iXU�X��s����v^������]�`���/\�9eá�]���%��6̽��Kt-��]"k�[��ZΉ̐b��e�"������Q2�ʂ'��Ӿ��^^�%�+ND"V�sn�N�/�u�vT�6ML׻�i	�LW[2��ܷ8���ݚ�k5R�>��P�u�IwI�L�������39������}	&hNƔ���[�c� 'C�ھ�[Y�k��k�2�g\��n�ۄ�W�F���[�-��I[�)N��V� J.��xi>�W��c�7]l�T��Ṁ�Y-�̢�Adʱ�-h�{=бdz��{���y�aV�Ҵ���H�K���"��[���qI=2:*N��8�pDВ2�н��*)G/q���=�GL�IDu=�9&Z.�t$��ej\T*(�&n��"�[�ܣ!273�H��X]+�YT�*R�滧��9�CirR����YfDJ�����T��UUj�-�IG",ʕ%��%�-,��G��b�*2͖AjY\Ң�Z:��ZQ�eq"���旮�r��O�C4�(�240�t6PYb�$�Č)Z�2DJJ2�#%3"(ĵhJQ�c�DeZaYiX���Gw4Вt���$%4*�R¡R�`U�,������TB$�H�T�D��Ģ.�I]CYUZʣAQ+*�3�rMRU�fURVQi�$F�u4���
I2�$�)�'��t��7^k=�a���J�/Fq֖kz�1H��<5mqR�u��:�,���Y:��LV�t��e�m���O~c�>��?l�Ϟ��u��6@~���E|�+~�r0�G¯eR�D��x?����F#ή�f㓭Ԫui
��mSD_Kf/�r��u�{��1f	H�I�+U�/���z2��Fb�����W�euh��<l����;|s[�Cr+�}p�i?+>���݋��2��r���[��:ۨ����U��Q��O.��w)z_�k�A�U{|2:r��on�fi��O����(�tP�*�"��*�LP<R}P��:l�����c�(�Y��_�Q��>]�#�|����������z��
��Bd�х��P��	���}ƆK��̋���#�.᠗j�Z�"hW^k�|���J�� s=d#R�m0���Q؞�x�ގ͢��io���9��9�F�y6 uHu��-A��D����^<���
۷O�%W�b�C���I�p�hE}V
��@w3.0X,�PG1e�0}��U�N�n7�=��+u�yJ��7xL1�&+C}4�-�Ã n}�X�N�"�����b�g9Ǩ���knl���o��]+��� hj0+Ä��C�Mt��ոE�P��4��x���!����f���"�E8w/_M���#s�f���j>ŷ;D&����nֺ��� ��b0�*�u8F������nơ����7$P�%��@��b����l�<�
V�p����+�Tc�n/UWG�G��47k�u����E}�e�3'<E��3+�V[|���N͛j@l�U8 ����A�`:����I3'I[�e�B�Qy_+8��Jfj;�'��\50Q��`���-1a�]�X�,��.m�,(ῇOZ���(}��-ad`��SXaq�5�Be��o'zuN�]׹#a9:q��:aB�=���2�*�����qS���ƴ����o^�:���
(SrE����l>��E-�X��{ UX<��[��	��Q>�y�{ʲ�b�E��Vn#O 5���m�M�
>x�w��F��z�/>�ق<,��qJ�'srGŮ�9Ժ�n{�
�O�c���r$)1x������~�/��(hW�p$��J�[���\v,M���F���J�'�xm���zX����PܦR2z��iN�ٽz�9���T!ȫP�B�o�2_*z�J`T�97����UHvӿ�T&X��)#��k���Z�b�͇B=�ӗ��U~�O�L²u.e��l���J�i/�'�9�}�r�̗��*�2�k��[t��+��6ժ�����+S���H�ܙ���T�>΀���AW�;}�v��!Yh:S띅\�`/S�`�����3i�r�]L�^�wC�*��x顈�:���Ӧ=��Ȥ��d�����꯾���d�⇼LB�����kM��;g��D ���:;��}C��
��2`���Ԡ!ob���B���'Ydƅojt,��"�S���"b��(:S"��雅��ce��jyoN��;w˜b��b.*�԰����F�a��+�T&l���V�:�M>�2�7�-<w���y��丙a���p��N�̂Bgt��J�Q	1_S}P��s��9W&a�2S̾�{�T�gh�e�W��0��9)G�ȏ3[g�|��/����k݊r��o�����c1W�1}�b����%׹x��#Z1�n�e���/F�X#m�O��О6��襑��[�z�K �LT4�I�w?{(u���v�Ӈ�ʊ��Qc�xArrP�SP���r�T�R/�R���� ��a����]'�0�E	X������S�ʫ[
��M7�U���}_^L`���ٸʹ �ΛDNa�;1�S7�E7 `�+5_%��˨{��x��Z�s��
�e��k��ܔ�F3_.�w�2W����}��"P��X�_t����5-2���|`�UpD^�E��n	�����7Pǫ�β*1��4˛�em(A�軍�p=�Xv�O=)��{͎�>�mu�h];��]�W����w�VC_6M����O��M]�^�D�_�����]')e�U��o�H~Ŋ��	~��°�s��
 믲�o<`����ғb�5�R�ЎP����1�i�_W���A[��P�7�/��%}�t�%��5`c��L!�l��Z��⚦�����Ũol����"����DL������;���͌�VК���Dεq�b���wS�h+{L�̼��w\X�_^���w�!"t{��r���+Ky:>��C��B౹������/�袻9+4�تl�G�9!ј�\��`a�����Eqx�u�F�,J���#l�����h���i6[^�Q[;=!9v�U��U���VQAY�.
��!�[�I����U�΄�"#�e�~�N.Դ��H���U�{,��r euэR��IO�xX�|��N0��}�X�Kv��кf)�^Ӕ�*�({�Q�W��Ǵ�Q����4����CH4wa7���:�j����`�zk��"�BN��-PjH��P��������.l<�f�V�W50y�凂'�Sg)�t� �ق��l/`�v>뜶�b�ѽ����1{0���K�V�GW7z/w�l���xl�UԵ�t+W7���*j�W!����}��]�:�/!̚L����ֵ�Δ��o�l��c{d8�z������\qb���5�>��^���'{9�~�;'۲�9��cG+���ƨ��]��� hI�,HD�7ޒ"�͝m���7 Met��q�1���f�,�c��E�F��o.���c���¬Y����
�Hіo�1�,,7a���`w;[7�t��6�f{k��5�m�Zq��䏋k����(�����s��(1�*&��i��|7���zx���A��F/�g�0T�dl
ǫ��U�\kMQ�'?r0�|*�*�N�	iW��v�~���G�e#w���n&;}uw5/�Z������m�c,�I��0��ձ���\����-�{���ٕ�	B
�m�v��kun;�:�]���ò6D��t��c�fj�i����_��-#�S�ϧ_���Y�J1���Roj�3u��演��`C�N�;FtS!�����2y�$gI�Ä����i�s%�+�-ZiW��C�f����(��!	; o\S� QA���_)�]@��yQ���ǀ�y���Jv�~���I��׳��>��k2�7x>ھ��[�˽
�����j鞦.��օ{]{k{'7�I��ܢF�����ɭ6�D��M�-�����,ý��T��S:���_�u�>� �H#����v��~���>�+sy�ƻ*eg��t�ϴ�*,�
��rP"�J&z����1I�7���-���v���c���Σ����Y��E$*:�W����r��*�t�#�u̆�'x�X��e��c.���$Pϡҫp[w�,wpFřf8E����`-���� ��mrK�
��0LLS��7��Cv��!ܘ�	��7܀�J�y����9(^��E�s"w�_n��I�C��eA����u<6��Gr��C+�LUCj:��y�i�����o<J�(�1��l,�K���E�8���������nWkx��s��RשJڗ_b����
��]�������in-�2ٻ
�j]W+k�\1��jf�P��+�b��z�������qv�%j��_E��T��l^�ֆ}+3g�I�ʯz[f�����H�;��Yۼ:����v�P&��mV8Ƹ��l8x|���&׸�k�\�M{q,���V
�;7���Z�7a]�tQ���qy
�\����U����Ĺ_(��;/_X�x#�o�Q#�9٦�@�i�|�� /6VY�&3�y�c��C|����λ�C��*1v�<i�g����Ȋ�.���$#��5�BW\{� �g/�o���>�ѵ���oG���%+�t-��P{��Gs{�ݬx�L�g �-�0U���wf�	OԨL�t��gV�r�'y}uR�N�
�x@f�f��⧯9�̏�|�ٱ�+�U	�O�Y�+���\�xú�i^����x���%{�m�Ors]�Cy*�ډ��L��;��.�)3�����D��Z/���<m4�\wm�8Ɇ���%?���T�c|HN/M��S:-�����MH��j�놟 ��9��[,���UWj�;�׺j����]2�f\~'꾉�:�m)�:���:ἄ7 .�Iw]m����mZ��Aq�0X����ene�O2�;�m�	��oi��EuU��l�a��v�z��zt�8��w��x��7����>؆R��`����}�S���Z��lW,�'��W5��@4�^�_m]ykm�����iYW��'X��]���<���I��/"bnM�=4}5��,�N��q_v�$hJ���T���;�߸�;Gu�9�Wpn�9s�t#&�k#���quk؎
QGU�	m�@T*�<3h�G�}��S��3ݭ���f��̅?6���� ,a�tV�|s�܆�t&X�׭Uedgk�3���3�&;����+��>?7u�o�h�k���'��_��_S��Q}���r�=7�+�B�O��xhl��JrWV���t�W�n�՛���W�q�D\�W���c\�63����	p�k�pG�??�����sV��r��&���]����v��K0!u��v��n^����C�o���sؾ{ë��ȕ�e�U˘E���ZvWmuw�rʋJ�6��O��U^�zj�0y��ԕ=���xG�81?�Z�dlM^w�{�V�����-�m�|�Z��s����Kɾѩx�����u�Ւ�ՙ�T_5��t�	c�)�p��U�ƥ;��p���7ww�Ձ�F���ȳ	p�\�����_t�)}��r���$�����i��
��v9$;�������lݶ6�Gf�(�}�3�S��	۳F�{)�Ir� 	W�V����Ը�Ww-08-Q�g}�+��q,Bm�5����o���������ӾLuW���ΦK|��2��|>��|��7��eG]�',�������]��wڝ>�g/���/���b�>�{�SU��k�	M;ǌb��#��c9�W�-�7x�8y�D���j��5���6]�Sv"i1��"؍�}W$�����S�c���Bƻ� ;�TDjN��Ȼ�����e���qR���B���u��bfc���c9��j9Pu�B�mC�K�
��ɳ\���YvmAר-��@ޣ}n��������v7S��]���8�|�^e5S`倷�В'+��Y8�^e����-eA�u�uy9X���TLE�7t�Yб=��k�)_��oe���P_eA�d(�>ū�y�ۤ�髢>��y�mw��m���o>Λ�-��y�UH�a��)C�h��o������t��b�/�|�58������7&��l��0�K|���wq�ܶ�V˄�~�Hզ��h�5!F�Pc������e�ƽO�rbs26��u��e�K���bҺ#�^���W�ӎ����%>յ>��<=���]���o���V��#�cҮ$��IxW^ͅi=m�⼷P*{���UUW�L��yG�էeYͯ��wUm����kr5�G�����M��c�,���S����?|#�_N����Vy+��GV����\���f���sѸ���S^�P�T?mb����_%\�ʸO�D}�`���/��'�۝�=�#u�ջnƄ�B�Q�� ��W�܏;�{[���-4�>r��q��k��n.T�!H�	H�H�Ϭ!���˃���7����u*���������x�����h�<::�r�TU��r���`q/;,of_�K��}!��*�b~�,��N!��5�}���}=1��%�?}������x+�LmC��tnV��f��2���Xw���7���Ɩ�E��xm[�Ջ�T2�1V�;"�Q�8KT�u=<�'p�'�Lڰ�	i��_mA�����+
��eUyx.�>{��Pt�(�F�u��S�}�J�
�Ȟ��R�Q�'Q�I�֥;�L�N\����,S��珘B|�F�j�ǳzt1R�Q����טs.D ���e��T��6� hﯪ�H@��au���N�Q�	�;�;BV+���gv�k���V�F��"�B�����9��''2Lx7�����s>���]R#,������]P*��Nu���I曓:�X�9|vq0�ςSp'��stoh��ܱm|�H�P��L*���<��b�v�w)�~�Kۛ��'�Zׅ���Ln�I1�6Z�'�̧��׌���#��i����M*E�*�z� Kg��CrV�	@��h��eRx�]^��gU�wu�"u{��4�蜠�A�/Y�v6��*Z�����G�C9��T-�<�2rTz���{޾M��KZx0��ŻL][��h�w�`Y|2���t��ѱ���'}�b(U��N��!6M-9���R��λ�\��z��T��9���6�]eka�����/���5gvawC�һb�Ʃ�+N���Nq�*g�n��ʒ�D9�%n;��V7x�՗���IBw>&ihR�lJ�=��R�홬o`���b^	JcTwgH��i��V�T�DQ.�_*DǏB���o��H/���`mGb���e����Po�F�[/]n����
Ί���YB�)�YJ �Ny��ͶOeZ/l��m�������3U\mk�Duk���Ķ�WJ_�]���Y7>]��k/�Ư�,���W'<���|��/�yU����܃}F���±�Y#	���M�c��ֱ��9�cU��lcLb\�W:6Y�n��j�A�6�\�{2VE�'��*���qZs�Γ�FPv�[��4o�m�=�x^7h�
�Z��%��R���K�t� >�XZJ�`$)��\��v͊v��Z$�W���<��F塮�#�s�v���wf��	Uz�wnfme�Ge)�����`7V��ݝf�V[�e���7A�zv�[ȼ{�u�7;9`U��\�5yAb�w0��3n�"�2�外��F>����nK[J"�������6��Q�5��p�;&�*�)��OA��qʱ���^�0���u��3��c�P�?��]1���>���܍\�mG��Gvvљ}"�#Fl�V���%�e(b:A[XS�6bʧg��nR���ܚ�Q��<մ��Vt���$�(��vx7굾5g��s� �p��:V�u��UԽ!`l�;���+��g�I��&p�}G���ẗ?<4X����N��#�x=h���*���,�A��x��euc{z��?+pA9��1��|(ރ�c�l�6�0TX�ǘ�����ܣ|��(�8)R�s#o���j�o�|w�{X�=���yV�9�$����s����뭘�Q��2� �����2V�$���r��Ұ̥I�r�p�m�K$��"ԥ^�!�z�/����p�ݏN3�zE�u,4�6-��b��B���TL��.EȎl®�e�Z������5%�UZjҫ�d�E[XJ�I$����#�'I4��2*�)*�K�I,�4���g�ZF��a��e��6l��d�iRk0��s��bJDTh]-�-SBƑΑԺ�#B�%�h�m�%ԥ*J�ńr��*B�ZRWD(�P*�Q2�iVI�J��'T�jQ�Q�\��ґ=\�"��#D$%0��-4��#)EZuD���P�/'=d�P�eR�l��8f�T��ˑ�����Ut���fBQ�
B�W
��PP�ʴ2��P�**��D���bPh�´��e����Z!Q"����r.Q-EL��9K2вB�"+�d�I��fDY�!Q)a�BQP�]&��*�j�1D$�*+Sպ��8O^����xuOO�"�8�I���n{s2K:�m��X�Jj��ڵ0��Q���������q*z����t�����G�oV������G۲].��������w5�:-��.ұ-:1�-�ٮ��j:+0y�x�q��hlי�߫�V�����_����3JE��{m�+��R��}Xf�l��I�C7��^�m�>��|��~��gZ�bY/�+��9ss����T���o6*�MoCW�=����]Qպ��Z����ae����]gD[�U��Yk�����5ӱg��^���Q���ÓKgz�CCq�T&K{Yկ܈��K'����EIϪM�����*�Ե�S;n;�}+ӳ_|�����zgV9G��&,sv��n�	>jaFs�!=FI��\�#^w�o�m�G�i���[J����M9s]������o-��od4�Q	��6�����|!��[������V�/8��e@��NL��ws���_t�)}��7�8��H���+�M�+��NHT�o1\b�ܿs;�5�<��0U��sݫS+1�u2M���_v��	}���KtcJ�S�y^pQ�uv.�ذ�B'3��2!ȕ�²lI=�e�0���:�W�����kP�qv��U�ݯb��E\�l�㘖h/�W�U}�^���L�6Þ�ф�"�f -wpfoִz����6n���
`%[ʜ4n1���c!��	��\%n^@O2�Ęȕ��9#Sη����1���w�B���}�o=����K��f����1�qF�U�mS��5&'��n�y��	��p_h����-�+�y�@t�_$�m��*��./8������tq�[�W��=.���J[;��D�rPY����37��31�^vֽ�FDwSnTʎ��O˦�,9���%�}�1%���S�����c��ʈ��ި��QQ����EbE�叭%ڦ�e�����١�v��Lm�?����^�]]��ƞ�L���������N�wu�~t��诠�N��=i�w��ZѢ���S���N#7���'ګ3~n��ϰu��ҬmJ��kASQw�R���{B�"خ���/�f�P�;>�}N$�e�x�g�/۴�^+*[���.�4�Y�YmR�:�$��.��*��}c��yn�S���td���g�⣌�xp��ُ��J��;Y\�@/Ax3���5ۜ�4y��ojC�Fs�AW��DG�}\��;)®9�/j깼k*MnC���Z�V���<q�6��Ğ�[4�E&�x�?�n&�����V������{�{ٳ�@o�D^�R:|eJɹmu㗼��p[���1<�T_5�GL+z�m�n�یq��鹼{5̔�v�z���Zl���B�	a.���~�s8ɜ='SZ�F�䣊�~�����`�{�����b�%�ڎۥښ�;3y4��n7�,�;,�%q�pX������F9�W�������si���	��c�~m�s�� <L�Aw��,���H5�}%�'�$g��x�n���R|ܾ3��wz��j_�,�"�c�m�]��蚛����<�n�^c�Zg9�YϮ��U�NZ�{�2�e��1P�<'��'a_)��{y��^b�ǵ��k\߳��#�͕�$~y�i��b|�Y6-RAū�z�����ƥ<�:ξ�!Y�^��Z�����.4A�5zJ�чG�N^�O���5����Z��s��:�r���{Y)Y������u��F`��=�x쒞s5]�r���U9��|���W�}_X�|�&�6�I^�w)C�X��yX�]�u��w�4���r��S;���0j�}Ӊ��T7�+�ܢ�(�9�[��g]9њK���\$�66�6)��g�y�M������mߴ�Y�>�,q�U�ܙ���g��{�C�Ҕ��1m���]�{�}�y�o�nJ��+b�Y,R�کQ�{׹~����/|�/�=u���S�����ƚ�Oz!Mv
�;yrz����ƶ\�������Aك�Ĩ��j��W�mZ�P���Zm)r&+3�c��r��HT�AON��q�<��%A������YG�|�5"���s�1�Bkt.�ƶ��w��W����D�;�4Չ�=���62wS��v1���)�u_�4���@��9ߜ��#��ď�Q� �#rڛ�{./�j;:�֞%,�j�����q��-ؚR�_�m�F��'��C��Cnsb�̧w�<��CUb�bݏ^�9��c1?�{�F8'"�<j��
��֟
�ܸ�W�++Q�^up"�<��(���}��vE��'*:�A��d:��jp��fgҔV4E��k��J��u�0d%�k�}��}wx��P�/�{�/��ٜ��놩[cI�R)؛�q�����q.w�v���c�i�&���y1��;��>ͨ�����b��>Ĕ�^׾�z����o��>�s+|�U��g,���-�5r}�����/E8Ǫ�s7+@Ϛa`}�i�E�*��+�������X5��<P�i&��]�~�Ug�h��C/jͩ��k�l�.��U��'�Oc��)�1�ճh�!��k���ߺ���q��`���,�=�C���O%&�X����ՆoT���>�fo�զ���g,��{�əݥM�{���/m=�Իzg����ç�p������n�%�}�ZΏ�����sy+�A6���7��^ߏ�v�ڍW{�4���MX����$Kg�#"�2�����n9J�����gP�~�"w<ì�)`�FoVf��͸�59r�*-+7��D������{����{�a���^�`��̸�ĺ��4�C�c6��|�y^�;��<8���������\ýO�ٶ�/C���;��8;�H�v�/*��]� ����EFK�g5|���������菢
ұ�.����Ĳ�svCz�u��i��R���}.
ϕ�Z#3i�]׼�*��2oj!��9��v�ͽ�4��o�
gᱼEP���da�MU��Qk�:ͳW­s��h�V�ji^���Ɔ�9n��*�2�5\�i�}yyK���>�s!>������s��}�慎-�3Q1�amo)��J���V�-0�yQ�	O]�@]�qN�JY��ɔ�����Ξ�ZjzF8�܅W��1�˶�'\/�[�p��U k8osk/U�Dr���U/�=\u|���*g��]�V�[b+��c�
��uEɲ�cԮf���w)�P�ڇ�T8���`}��CQ�Y)[��Q���zk�gc��8��N�䬻�Ӊ�z!)u`y��鼈���z���[#M{<e1Ճ�w8��ux��^�X�;���Q�F5S#K��2�g�U��ya�f�ef�-t�^�4VZ��	L�]��Z4e_Y}ud�+��0�#h�XT�T�8�S�N��+��M7Yq=��{}�����9Q��"Geʌ嫾�\
�y�E5A+ik����cُe�6�w�R�)ש�k�k3��꯽;F��=۪:/נ;���*ϭꨋ�ʁ���]J+7��:��%�F�77�u��U6X����-�<U��G>��u/mt�:W��bM��#�\;�zM����r����by|qq��V&$��uL�z�4�y2��z��������{�j.�pT7"T&���S���oy��̧�mE�c:{~�6�b�|��͈׼�Ъ!��u=;�xc�y���r��tLR��cV���'����ﾥW��R���d�괲���rj6d8�R�ĥ����Z:U�w�5K���Os�;���bP���5�g$(w8����\�@K�}����r��㥸��UuT��k�.ʙ�x�4�]�9Fa�e}�`BR�f}ve䍘;b�97���y����_j���;�;�������f�]J�U
��u�O6�}�*fZ iVp=���u.sJ���^E�BC��o��>��ޭ.�Ѥ���.oԭ�x�wq7x��[7m�43v?��X�M�=C��vq���(k�<�mQ��kgV!i�dyҖ�:���E��{�S�8����En�i���>��چ�7�P����m�kk�s��[g�������g�[��'�O��e<V��Gbq��KY8�f���eBN�����W��"�M�5Wv���I�@��9���귦c9�\���Xv�S�l�.�?Ob��m=nҬ�UF���7 [�Rc��|�����ᬌ݆���W�H�NoѲ6���W)�b��	e�,�n��Db��9ٙ�ڇ����\�8���VV;�u����;f����@nT�G�\�Sn8�W{��P�x�׽�]JԌ���-ho3__MD-����.�<��f��1����8��8�h�ڽK��!_,�ڕ��ڇ�9|�ܖ�yR�I�����%3�DO;�yqTnK���ookq��Gy5*Mg-坝��%;Ѻ�I{ƥA�u���\d󯎭V5;�L���pL=�c_X��s7��H��eF����� ё"��`��o�6𞜭;Z:�ˉ枭����U)gg�_*N�2M�78��0��]����N%uy�%>U>�� �g�.7��걬�_q�
�J�ܫ;��l���I8����b}�}��p�ӎF������{_CUjo�Vڃ����Q*���R�h� 2i�G�F��`����Ns�����)�J67�$�v�����bg����f�+�{0k�}�I4�\w+�dӤ�!�e\J`F��'�y�M���ݝ�U\�����?w�ᒽ'q��B�p�:ǊY���F�[�7�`L�j���_a�at�p?Okˀ�2��P�]p�ô;�o!vA�59�S�\�5a��!�o�ό-�����ɫ���+�L6���=�<ʘ�m���b����ђ���+6�t��1��r�5ӷ�"TOں�*Ԇ���UDsP��͸V4�˂�D�ϯ1U�9m,�ӱ9Q2�q:��Ӗ������B8����)�y�m�au���;�Sх{�������9X�3�;����hl�۩��e>s����Z���=P�*8��Ut=0u�_�x�l%�~N:�w�����#�M����t���Bk&��Ws0B�I�-nI=ר�r��s�Z�:T�WQ��<�Ѯ �����97ZTE�V���F�i��v�⾬u���n��FF_a�Ҵ,��ٟ���ms�q|��zWW��/'+c�Q�Q��zYfeN�c�ܗ��~Ħĺ��4�U��K���QokZLyu)�^�7���Pk�yZ �r�~	��zB��o�J���߲x�����A�YV�R9&��^���Ӵ���nF��ie=��y�
���V�Qy1k�,��)�>����pwi�7}������d�j���A���k�Q\z�Y7���X��[��v՛��˸o�}��>��g,���m(R���"jN��7T��{���7�I�9�T_5�GL+{54�5�v���&!�n������7g5%��V�p#��G��9����h�K�����֮�����۬�K���y�ƾNYW�0��L���.̾)�iJ�=�c�r�ݻ��9n�MS�u��B��v'�R�W.ڃ	�W��7�K�Q�x�އ;ݙX�~��6�1dkDf[:�[��.�޵tX�H_v?d���ﺣ���Z��a��F���WC�]��ЯuB��i~��k]�v��zZ�ؙ�k��X\2M���lM��69��*��G��zF��K�X�w�.�lf�H�9����U�����`g0ucx��ы��RBu��2<强TH��Gn��Ǧ��*b�j�j@�SM�\ڀ\<S���+=�3Њ�Ӷ�ˉ3Lk,x����3�뷌��{�Ea[����oR<�8jţb�N)J']ΐ���劉�iB�Z�lj]���fg4pjAǟ���t���{��\A���h�\��r�7ϣ�W�^,V;=����_�����°���:�)!�0t�uqަgg5����������Y�[�Qm�40	}[w�M|}�<cު\�;fI����J$��0!s6_:�
�cd�є����K����}(W{g)��$5�4>�З0R�n��Q'�f�$���5�w�;sX�fC%Ѯ"rOU��f�d֮����lxPy-~��^���O{"3�$�,;q�j_���S��Z�f�U�mL���/��8jq��:vĺ�����������-OIx)<�Z6����Ӭ��͝Ž\�Ĵ������Xh[�@��.��Z5n�+9�v0l�U��Paj��0i>�� n��/@1\��ִ8�|4\H�fN����@cq���q*h�r\I�v�\�G���݉o��F����ٙ�T� �w�/]T֦CI��f6���⻽v�5x❬��!�f���_	���Z�wS��t���'0�X�VC*E+*I�Me�r*�H*u�6�%!��.��T�KY���:k���k�=��!�-���wǒ�����N9P�)A���)�Ov�T��Q��=�w�̽^�.ă��xZ�i2���M�3�v�AM�v�=�9S01���cdW��\�J�
&�IX�<ǽ{�J.��ݩ�jvE���w�)�闼���Hy+R�7�v�������D(.u"*vTŚ�q��Mڥ�nN��lG�� ��n� �����O��L�A5p�0mT����Z3��[�ı��'�<6ͬ�䵣Om]
q!{�C��@��ms�r�gV���=vV��Mp��on�ɳ���1�j(G��>ʛ�;�����L��e�1�~Yf�����O%�5{B�J��*���N+�eu�	���w,�d@���B)�<��.�+�ZT1��喿o�C��p7��(�[�u�[��C+�vk�͛��A�PK�a�<E�*X�Л۶����ben�r�q`i�z5R�6z�>ȑu���+�2��<yٵ]8���k�Z�u#�Wi������.���[G����q��{��C�������o,�/.�,�M�<��y���T��q�Gq2�Tu����x�|�W~{�����k6�ǟ~���x~f��-H�+FsfEF,$�P6�P��e�fR�P�V�Z�T-�J���<P���W$�,2�"B�8i�t�),�����Y�A3PЩUwq$�E�(�STN�f��R�b�e&�URZ�8Rt"�Z	d��0��&a4�j�����鈐g��PGr��as+j�SEJ�֜�pvr���hVD�!�!$�*霕je�GB
,%�Na�e��-E2�4��%�йTHr�!t�K]\͡�p����f�QZ"�̢�p�rٛ(ͪf�$a%!I�t�j�&ʳ*���9t+�Rt!3��MfjaTE�eeeK%J��\L����_�)]T�\�TWa	ڟ^�{H�f�eB��>ٵIXֽ�B��;�:�N�8c����/x;��:�ƞ�����p��}��v�+e�sz�_hڈm+x13_���	Lh�(����q�$�ejV�ęz�%���e�r���M�|C� w�1�e�.�+���q��}�����6����,c�:�TG9
���!ܺ����V�P�biO�=:�ؗ���.�)*�{_zb��ݮ��z2���'�:�95ͭY�ono,[L�/���'ϧ�b�]��foP�%�"����ײ2}�<z�%��tSMx���m�����=�Qo�qͱٝ5PU�|����Y6���鯞�Ԭno��i�\�����t]��[��ak�ꬸ\ا����n־�����*ƥ�޾Ք7Dr��j3HL���m���֛���Fud7����fd�0%�u�Q>⻾�y ����7Ӹ�����N��]���R�]80�lU3��K�WE!��r.�����%���.��eN^�vmu���ŗ%�FTSV�6hoc��a��/ӑ&sY�������/p�A�љw�k�M���i��	�^�7��%��/*x��/D�����t��c�}��F [7�郤J��u�M~���6���)p�����ڇ
c#YQ�)p���7:~V���U|4�<:f�O^�:��ݨr�
���ᰕ}.d%¾��-h���=8&$��$����t���'�Zqܯ�q��:F��W�h����0룓��u^.y����f����j=OS���Cc@��aB��1κ1-ꬭ|T�h���}�,���k��;��2GlCwy[��/�h�2����?�1.�%�7|�ݓ_b{��r���'S_5���NW�Vd�fo�͝X�4x3�_2�t|�W˗�������^'I�D��s��Sܝ���a���ܨ5=�R�+�~|�gڻ���x�oZ��m��mO?���E�lm|Ժ����_<�>YQ���j�OZ�qg,���1՘�^C�tݧ8�43�{{4�����~��m ��1����y�+�8#�d�������(\����2f�:�<"�\�	�a�0M�yѱleZ8FX\���o�Y�N��^ۃ\�\MgE�ݎK%)��+/z�go���1�T�P����䳳T��Q}�#`��Am%��{�]�D.�6�a�}1����F�cu{
�Rη���}T�}5���׮��Ԗ-�N��ڣ&/�-�t�n!�S�7ZCv7��oj�_��6$b�:�v��8��ڽK��bߋ��:5���1����n�^[g[M��Z���Ѷ��R��}J�-���}<���o+�|��ШM��s��J�F�M-��|��5�HiP�C��PgZ���\d�:�3&N���I���t`-+�?x��fΗ���	��u*%&2�&�U��rd�3�/��N���	6�ۏ��sM��0��*�N�D�}�ޓJ^]�L��y�/GJ�٤�W�;���2b�%pͲ� BO�>1�*�|y<�WL���s�0;��|�kN�������Dnb��`�[��9�ƌ�sW��]�U�sڡS�����]��6��C��q�#
�n��v�z6ܮF'Sћ��p�j�Gu�kV��y���LiD�5�vv�#�m���YUw��3�h}ВT/M�1t�E��e�U���z�}���ͣr[�vS<��y${H�yf��5v�V�i��e���ܴx��^�Z\�c#�3;�ܸ�t�ot�0V�@C;�?W�W�.>�G�N����T���P����
��*v�^��չ7�6�z��ɛ�x�0�� ٧�Gi����>�3n��0��/��>���'�cO���A�l7]��-l���/[�Wn�*�ꃵ�S��]C�:�
���UWc=�vp��{���3Ԓe�w�ej�ʮ����hv.{u4��z�-;١�ǂI?{�n/u�@�o����������.��/�(��ک�;��a�W�v�g����5t.f�����^u��nq[��Q��t�����{yq.wʗ#��v��I���my�{�_3�&���������wgQ�bi�s|� �S��m�ks�{�����_\w�rT�ZP��W<�V���:�vv[��z��=P1��m7��\���Zຢ�����7/ns ٖ�-�M^�qYq[�{)�&�Ʒ|�.ۆޣ+4��S�\L�>�������������9����ѵ�;�T���vг����h�\����_8���N�mf"���$k#�s�wa��v��X큘���I<l�_^'N_$OpS�Q�w��ǚ��L3ssUss�����U�$\���bV�@�u���.�g�|2t�y��O�/�x���Q|�-�c��&��mm}���-/l���<ņOr�z����+���5"�eOE���y��2f�zJ��g�����ڥ�R{s"�:F��eX�X*M`�����-��˕zX�8Y�w��YMt5Mdq�q�7��pڟ���M/��tW�,o�G��ue  �9��k�n�m�m�}/����w_7s�*g���~�G��N��X9�/�ҥ~��5}�aR��I:x�>P]�z�����'���F"�|��ׅz�]����f;S��Pu�B�mF�p䰯�sm:ܾG�5�a_)���{��]%�^z���e�~��o���.�5��L�lm)�)�wާ良x�j��
�.:}��iõG���s㗧���E3_���"�[��\n<|2��[�}F�A}��:��x��]����+	3jfu
o��K�/J2v4�wW�z�maq]{�oZ��k��}*'r�m4�N�e<8s�r��z�n�	S9c�5e�m�T�j���H	�=hn�e��Gi�e��ֹ�������CR�yJ�5s���0���0U]�����"+�z�n[c/!o���Vl7��}{4����m�^�Y=�`9���L伱�[Y[2�
�P�k��͊�x�nB�����6�n�"�{'H���[I���W���x����D9�PSv��G�{���og�=�D�X�P�f��K��Û�������zwu,�߃���y�����Vn��R��đřt��.;�`dc��1=�U�Kl$�����L��\����5;L�6Ʈ�:���+;��W�b8�i*dn਽K$�{#i�7YP[]G�h�Β=��&��Sp���}[��Q���	LJb;�\U���u�f�1�r����t�)�/Su����n��)F��v���I�J�������U�|� m�i�_.M�T�C����Nv�R"�>ʹ&�kW�)�h���@�+rkݾ7���N����lf�~�4<o/�4�%��U�5��܅w;V��]u�I�AM���ܥ�̩��n�#� ��1�����J3�W��s��qɈ��bc&ԗ{�w�
��5bGAV�"K�+o����Ō�B,T�F���w7Ϛ�%��@��,�t7nehp�㪪�S_s��V�V��4��6%+(�%c':�0��]�7��S+|�}G��NS��k;q�X{��\fbT��y�5�.bP�k(F�l�)v�^����j�����[�콚w�j��OQ��[
��?�,�=rmz����w���ݞ�M��ƣ#�U��Nj�wS{�q�Q�k�N��7^�imP賜� �m�I礳����
�{�}9�-�(ﯓ	���7�O����ōFN�W�'�n���3X��]ZO\�\���X�|��/5!iV�����t���n��<d�����
{D�ϯ���O�U�}:ڏ�=�o+2��
�t�[̉j���k�W"��W	���>����2y�kF����_q�eU���[��Z�W5�#���=�"T��*z]8�Bں���NuP��ԩ췙Gi���5n[}��5���WvU�r��Ɣm��t�?9�ť8��W+�99�n�f��f]��G��@R��&c�=D��{-ۼ��-��,�ЈC�\��E������Bz���o���Z����v��F\��kc�tp�7.�f���Df\ѾʁXB�� �����[� �]b:�Vb�fl�Zٯ�i^�	\=̯��Tͳ�B]O8Մt"�����ܾ鄵�L�O���wza_t��s{�^8��\c�ت���gsz�1��bЄ8��@��#�Eq�Z��.̽�N�Ld����+=Φ�\�;���,��:�M"4����V�by��dt���f�=�<�!8�U��ނ�:�����
���"�뙾A&�%����ד����囏�L��I�`KLvY}��2
q}Wj�����=�g=��k�r�MIM�9��;
���:�]b�Kr�s.���
�`Ê*S�-�˚w��3�'��-J���wWT�9e��0�O����4��|��V%��T_V|f�mTW�%2r����^+o9���Ov�vyZ��+l��W�wߏ�ꔽ�<�v�<5�n�k_��\�Uck&�V8*vq�M�~�|������Ϯ
��t;�J<2+�t;-��6�[5��̺�Ǔy���xA-8���OM��f�P����wG�n�Vc|�l/t�vJ��L��+����d1�����9�0;�g�_q��lϼ���|�m�����>���^�tGq�r�}ʭ٦h/�_4�����{���}����nJ��ݔ2�B�Y�o��x����<��ڴ�M[���]��]q�A�J�
:;+<j<l���[�d��VV�M�������:�[����馻�,��=U&��gw9�['�`C��1��%���_5}GJ��4��p�G�7w{��WgRU���䙼��M�6:�Gt��3���zx���Ϲ�0�t//�a��_H.r�%���l����r��B���_<J����_DO�r��n����=��jc�Χ�9�]n�RB29vw::�C�+̖��#W^��[�#��/6_4�W�Rm��q�2໅P��*���퓳�YV3�Z�&3���v��g������C*tڇ�Uï�����¨�MzОRQ���Ɯ�+�����9��<K1c�ˎ�IjK�w'�ab�=��o�S�J��l$�hm�x_��3ue(or�W	Nބ��K ��j5�ܱ�R6�]�����`X��I��"Tij��f.�l�g{�z�׊���o)�F�P�C�0�9(�3�k�p�yZϨk{TR�|��[3]��TZϓ�zR"����;yb�Yj��9���am�ǝ],�{Z��^ʩ7޸�0�d-m��Ȏ)�F��ת�Z�F�`��k�N}=ʜQ��i��ŝ'17M����C�[{i<hdv���v��j3W�q]���[���j��ዋ�v���+�_g6)孿���м�j���V١���2�����ɞ���k������-u��ևې�u5s���2�r�,iVr�'�PN'�S�k~��G:�#�,��[�ފ��nr�O'�QG�k�=:��dy1Q='\��d�Y�jy.uw�k�η���k�	<ߪo��m�=���/o�+$��=����W<�^��OO4��OQ��J����L7M�q�����lpf�n��΁�Q�:��Nm�w�.���Ah��9�f�@�)�|P�;��Z����dmj� 북�_K21����P��,R�vs���=^�ҙKD��݃ ����T.�W������j��0�s�;$��X��ɛ����`m�h=+4|�V[N�\͒�=���|�c�w:蝃� �ܶ�����/�`�51��f4������.��U�箟\鳹f�W�� �Z�`&ay�>Mej��*�Nrx��vR��.���M�k���iʙ K�9� �)��z�{*ZL����M�U��C��h�1�����q(-�-���kί���)���p��9�b'�X4�:3�CivLzh�-,u���.o+�>���1����_b�=�="����x-͠V�Y�����uu��AmWOk�o^���2�z�C�W�$q^�W�h�Ўع�­���n+OB�D�����t��h��ll���̈́l��:�͗[M)����uS��w�%f����)&�o_I�`�{q�bDa�����e/^�e$/9qϞt�ۉu`:_u�(&�F���$��]YT�G�9󺵇\��:]�1}-���7�k�֣��^�k�Lg��/�d�(]�Ӻg�2�v��/��Uޅ����G旸s�B��_����ڛ�qj��sF�|�44���BR�γǳ�X�'G�>���Z��j)�r����Y�yU�qqh�İf�w��y�^dHod�L=��N)v�z��b����J�`nkOBMi75�H�󨑪9�-9��J[*�^1�/�^sJ�5��4�e�v�O�VS��/k����A3�B����^��i(�;����%F]c%۲oDo>d�8v'�\������F�ק�U(o����h6qM���M�r�T h��T<:�.�T�W�њ��-͍�_Zo�:A��<�+ҝسv�j�~�Ŋ	��#�VN�F���)�j�;y������):1���P��L|��j��)J;)�.:���iU���*a�z9Ӄ�oۥ�5��%�Oq�i\�\���u�+sea®�V�[ŁJ���`�kW'e���!==U
7�%~���8^�6++"0ݕ0Y
�6
*��꧖�xWnS|cd�R�C��";]ͥ�yX�
T���cr�^�x���L���R����a��8v�.�8�B@����ѭw(!��>+2gv����yv���`�ĶY��e��-���H����䕺V�
����;82��0�R�`>!˫�e��2Q�r��-�2���+���g s˴����`g��f�����!������iS}��ý��W|1]�2��y��D��ϥAN��fX���l���\�_e�x�K�&���u֒�BFf':�t�|@�Ǌ�.Ų��{�N깞M�Q�MǷT��6K�{���5�q��(0x��9D�ps5{s�!~��S���WgfK�D7�P3�k4L�M@�bWN%I�+@�B&Tg1	P��+X\N�j���)#
4(�S5���r���9GE�L�PT�$3�ciĥIT��#3��Pa%�hRI���1a�e���
���i�iD�PRjV�F�VD�`VBDW��ZEVTDЩ:B%#J�(���E�YhQ��TDg�A�E��E˳s ���@Qv]6A*E�5�RaȭNr�-J9E5�h��� ����U-���i�EQ����(��IC���"J���b$TU�SB���*���MM2�`YUӖZ�A/w(�n��Q^q9fwK3Q!$8���XNL���ÍΕ��y������p��٦����*T5���ٷ�Q�5,��0٣����.��n-�V�7��ؑ܍��i��)���n5���1N�t����J�F��}[����4sPs�e�ݪ�ﵺ��M�����b�C)J#��F�8N)�oPv�]F_l��_Mp3����֞u�Mu�J�G�o���RE')&�jD8��W��Q[1L[�Q�����cr�8{�Uu8sz��v��g8��'@KLp�/���ڋΧ�Q��ߤ�͝8W���G���>�րy|GcP�D�-a�ۣە��Z�oP�;;ϊ��d2�(��+0���<��]C�v���
�c��=s��n�Vcy�]���/��
>��-�	�~�^��m3}�46~k�i��C�7�Q�Ev^k�qR�S[�ټ�1�:�z����
mmC��n����*�|��B.�w���#�g���8���ں�oLZ_u�.i4�lٱ��w0AX߱�`F
E��L��!�1�{�Z�%��n�@*+UÞL�D���vQ;������
_hThf�ks�4�e��Sޡ̪�,�u=��#"4pn���@dՎOGd�o��V���hz�Ej�����*G|"�d�Z�S��R	��zQS�|�l�W4��~�[�Oa{6�����j�Y����$�\��͕ϰ�ﻛ{�H�W�x;�2O�p���8����LSu�hv���1kW�pf'���K���S\kT-���k��
���X��:�ێ&����_iOԱ{��PO5k��p����ul.�Dє�kJ={���[}WNz�Q]f���Enz��$Ҹ������'��������2��lg_)N}}��'�G>�����.U��j]ޅ���V�P��g�/�'�v�}�lqz!o�\ek�]w�5�gh·���~�^n�����Q�R#F��"�2�1;�cF�]�
rn�9�fu�����qmp��M4�|S�V�Jc�A�3�_[�<�%j�\�.9X�\Zާ�+���������X��_h�o/f;a��|)	n�{YƲN[@�����|���hj�=�Ʊ��\1�;`��s�� [��X�7��d��S������z�R�9D��ZKv.5Մ�Z�z��u��Fc����d[����"��G��p.p黽�8e/+Q��*u��R�ps�j]�m�T`��!�Is�-j�
pm`���j�V&b������p��]��ӎa�+u�kVb�˛�fu��_�߁�|敋myx����7��4�MMDW��|��}�~z�׽�o�����~�(v�n�Q��R��"��8�p����S����!Q-n�7��t����BX7lݍ��s8��]N�K��ԃ�'R�<q�{�>=��#����W�˥��z�wQV5m����'e>�;��B��x�8����9��y�R�۵�i�t��j��w�Z�v9�I"k+N��{jS�u��'���B��ek�j-�~|�8�{���ᷪ�*3g5���|�n\�S\#�25Ԩ1)p��h�V���sSW�;*�r�Nܥ�3���L'M�	\J~	TK�K�}k�-;Ӯ��v��M}���c��K@�WA-|k�Hw4�Ty��k�"��;�n�*��WW9E}R`��w%��5j�p B{c���y4��v�|F���C��o��г�wE��ɻS9Z���v�z�S(Z���m�#��@�_-��J�+�_���nw��9�h�%��e�O.���'��1N����Y�c�`7ޅp�{�����o�@.f�}Ҏ���:���[�4��]�9�V��WR`2����f`�[nY���BMu�9�v&nY
��"��X�9�e�%-O���ל�Te��lF'�}����T6��	������1��3�@��-��n��b#@y�� �zR�|�.^��糶�</��;kxmsm��[�-8ٺW�x�4]|V�A�u����F�b�:S��P� s�-����)�2������W��s]�B�|�J�����{5ėOL��Ÿ�-���.�{{-ؼ�7(�ʃ��eY��N��C7��۫]>Kt|�/��';�~P�����#�����m�C�zU����#=��:�v��G)�/V8�K�m�sb�'ګ1�ܚ�ʞ��}�}��gѱ��u����!6�v�Ĺ�O�)�;e0�R�,=7X��}˚̴3:�Q=�lx���=�K�dPp�k"r]��H�Cej'�g2�����_م-����CE�D���ĺ(��,8qwRTn�0�Q��17�Jϻ�oV�c�A�g`��\��D.ְMS}�S��zeq
�8�jɪ���Vn	�m�_χu\�-q�Q:�JηV�:���f2�]|e�ݵ��a9N#5����D)�\(,P4dcQ*ғ|��������*֪��_i�m%#�J>ʅ�u��3QҺ�G)��ͪ�gE`���&���G{>�*�f�4��bX�&�%pͲ��	ou��F��uoN�.���V�ϭ8M_O\��%#�/��
��S��pU k"kw{����K\9�����ڃ	�W���fpO�����S��"z�|���{�Nxbu<����-����sϷ�+9�ߊ�H��9;�㻢����^��o�R���n�Ύ�]¯� Ħ8�'�\��!�.^�ƽ�WV���KR�y'��hc�'[P��˨
����;�ߍ.ߊ]ي��O=:�����V���&f\�CiWl2� _v)�Vff���5��![�`	,�vr����
VT���l7��Wl��s�ڸ^r��&��nYA(�Ȼ.W_�o���]Q �!:��o�p�iٙ��;�J�t�������P��Y쓳U �(e<Y��R��Y����w��D5'���yO���RWŬ��0�UgFv,��R�	�y��y9��6�v[mN.��{u5��[*���q��[X�l'���	Cwg}Ar�ۼ�QX��R��Յ�޷KC��=�t`��ժ��Z��.�ʊ�+l��P�/����]�1mQ}֞N�b�d��B��yZ�⥮;����}cc,���M|����z��>Տ.ݺ�QÚO]U�
�<�����l�Kn!�댃��\6����8��5Gs�ʼ�)�=W9���q��U��J�'��k�<��f�z2LA��֎��N2������_�f=8�W֓��|����8]���T�}�B��!��\�mjX�y}��8���F�����pU�^���m/Smz��Wx��S�HԽ~�1��z�p]���JFBU���.wp�vq�8zK��ix�h��Z)?wCAZLU�0�WIsQ8�<<���x��P�Iߨ�4����HG3	B�R�nb}���㖟X�p	�f`:����DL��*	��!�{�ʰ�[�����J��:�8�i�Q}/8��a��3�m��uZV���xu9���o��[o�5��M:F�nYV!��	W]�ٗ�ŉ��� ��g��5GZF�[Og��5���[�LE)G��]���"�Jܸ�J��[<:)���W�뻻q���cil�Mg��y@+��{,
�s�Q�35�}s;ح��*~��lD	_�x��x��d��|{�6�Xr9������@��e�W��j<�Ľ3|��h��my~�Hɽ�q��W��}�iµ��K=rN��ή�=iՓ�~t]�Ǽ�OO�Mdf���0�R�~�����{x	��>�f�s5��6{������	W��Sws�&~��9�}c�d]ۦ�g�iZ]Y����*���i�0�I�PKG.�mr���� �[ߋ޻���v��Y��m�z�K�v�3�"�:jg]~w��~��U����������j^U�{U<�@���-(����}��ò#�����m�����9.��y�j*����T��ތ���2���go���ǲ�{�}1q�B������^�~�~+����>���Ｖ�7p���/o
�{)��˙����ߢ!_PP��ۃá�!e�_L^��z��b�������9U�;z����5��_��j�1���Lȕܙ��⬊7��q�t����G��iA:�|���ݶ_h�r�!d��!n��tپ�i#&8-���k}�g(^�k�T���{�3���Ԡ�:��u{Ǉyϙ�\���ő�w)Es�����g�Gb��?(��Q%x����D
�P���>�#�{޽�_��Cñ��g�2�z�8�/����x3a�k��x��C�1M�'t���9y��}���
�#מYs�w��X�u����+������~�W���,�9���񑅺@�KG���8��z��=��楙���>��Wz�i��"���D误��@����. ���aժ�4���'�w��5�*.��n�~�+~9��+�u����%�{�x�4�`�s.H�Vs���5'�~�`s{{�Fr_z5��&kҙх�ӹ�2Ʒ�c�3��A����O� +�{.��Π[�7�<}���u>N(ړ\�L��M���50�c)��5[F�\�wd#Lm�N��^7·�5����@�Qx_P7y����g�ݐEBlR�|���C��+t¼�t���������iUף}����՚���l�uP	dzr�xaz(���Q�X��6��n�;ͯq�/���_M�ǽ�O+8��˕D=O���&Q�[5+���*tʅ�>C}îѝ\8��r��.��P~�*��V���FIł��4+���SVC���C��{}F
�'��(���[�[�=-]�(\�����0��qHE;��E�}�pVzվW�Y�'�[�g��?&��k��w�g�遆c�]�ς�X�d��N-�z�;�<~��n�z��ƽ��W���ϸ���>�_�=��5��w�9<}���{�gJ=8:"}(o��+��[{�_l�ft�������O<�k�r=~�㞵Q5z�}�.���lP�xV���}k����#,��~ɭ,a;��w:��H��1W�Hz��u��׃ے:�_��=��]��ڤg�/r�(��	H�y3+߃�q�Y�Y���̩�=�)�t��ltq�(�2�r�e�W�5>�s��^�]��דÖȕ$0��D�0&"����)���P�UX~	�[���!ک�{��GU,>��L���[-U���9E��r�3�w��&��"_
� s^�'*f�7�
�Ӟݫ������l���+���+�~���\ #H�21�g/El{�-vJ��6�d�@�M�����j�-C~�x�A���u��k���˓�F��DmZMo�7�ܾ� B�G�Q��!��kg�{�특�s({�(��1Fm�-����R�N��E��p�cN�t�����֫A��rₚ��o��b�#Z��5.Ǹ^e����GhD��Y10���C\���l̅��i
x�7�Jݦ��;��]Qu�Ħ]�q������@���m�%�w6��5�h�]��8�m�v`� (?4���^3��bK;m�]�ڊ��L?@��ۉ���D�����%�����zR>	��噛�{r����]mkxV%����u`����W��92���&@|o��DS��:��|�C�Y�#�E�}3W�Ίk8i�Druh�:�� /z���EO��h1��B__�d������/ {#bU�Ը˫9G�G������7��`J9�UQ��&��+/�,r77,.���>�å`��%鬬���<'ѳ�f�K���2=�3.aG��O���=��؏$����'�j�qVJ���=TYsý��]���������^��b�lxk�o���y��巂�*NU�#rY��yY��R*�F�яDj}��v�j^W��q�5�Y=�����V�$?d�&g�2�z�9�O�o�g)��c��\(~��+EǞ��9'�uLó�[P���u�� k�����d�U�B���d�}|}���ޭ�I��M:CE����3$��2�����1]��w�棁�y_���=�^+�l^� N�}9�q�~�qϷ��_l{.7��c���Aq��W�����W��5EFc��s����GsQP�K��3�d�}�C0��.o(rNwOA�.�����6��qv3th�O�������L/���)��[$}Р�Nq��f���9��)�_��!�=���-�;��<���37Ql&&�_�i�oF�d��&�U���6Ѵ���O��/+�Q�A�+�����w+W��E���֏C���C%U%x8��j$Y��O	�����5_sR���x�+n�aT ��ޡ���6̮�ݷ�2�TF�f�������Zk�K�-�T�����g��\C
j4$��	��;�:�U�.A����E�y�1�p�f���g���	������Z����-����TV�-�B�5�	��D�jw�K�.����|���Z�ٛ����c0�I�)ZV��*1ż�c&�Ĵ�Dc�W^���5"�ܳ!�3߆&1��Z��㛡�n�����6�&Ö���'�1Jͽ���V�Bڎ���x����)���\���h)!*�ŉ���8��Lnȥ�ݳ�:"s�q�ae>�ngC��mExT'�&_W1j=.F��{)�g�W��[��]*~{ѹ�]��壆�1D^�v�;��|yz��b��Q���x@�;Q`�/���ޣ�r�"�rw�Sj�)�Z��w�i�b��SR++��+x�m%D�r����q��3S�������}9T�Sj[ox����<w�x����}s�2���Q�?؇��9˴v��!��������yFl^g�H9��b�2��%]q��2��N��
��`��$KI��N�\�N��Jǋ	�S�S����	9�����ܬ�����y%�U��u�ܫ|�ڂqz�n<����<���!���KF���<@x8 �����æ$Ь��gS�^c�O2
@ZZf�۲,f�O@q�طS��.�#�ȹ��ڋcP*^�}8{J�Q��{l���?d��>A�e��Z����z\[aF��0��eAPLN0@B$�8ԏ^�[��v��2������yH
�E҆N��4����B��69�I)�w�&�ʹ���Lw���&<��(4�laΨ������,|(�w����A�M�Zop�<]�!�q�B11f��T�\���{�=O{ЧF�ZR#��;/�E�!�g������/Zin�l*�lge�%��TUٛ��%�k��T�nS�Ҩ��_woR@�u)��xhe.X��驷�&����3�a�Q[��a���X��np5|���\G�VO0i�w=��Q�K�yC�_�mzm�l��;g:��W�N�4&��xi��Q��}e�eĂ�`\P�kk���E,��&����+��x��wY�P#n.����a�FN���ma��L�r��[+�B���F�~��s{�˪q�����D�C��Az��:d�GUogb�o)�M$���H��"�w	��
��s�8S��\�"L��$�U�B$�9��̗Y�AÖr+)��\��t�Rt����K�bG-IDj�Tjg(���B�"�H�ȳ�Ē�t�JJ�aB@EQ��ft���J�J�(��I�ʪ,"�	PF�y&��HH�"�Å$��7v��fg9D�Eh$ē/6:��V*RXf&s�'8��h�f,9�L�$Ԡ�B���*<�)0��L�YQ���EX�d%DA��D�)�A�ʱ)5���YE\�Y%J�$m*�j�MaUAq3�X�K*�épDS�Nw<�T�ŔdQTP�;����H�R�$�D�~�;��^�$���o^��!��ގ��w0���4�8>l���j���;fgY7z[��|���P�̎.���D�}̬t�����ޔ1u���9��\�G�/ţ��P���F�5E���]�B3��yg_�B�P�T����NM��n�H�ǟ�d>gF}��K�{��7��q�T�9Q7��C�v!=070&Q��D�5��9�T����q�^��!S{�B�?:b�}�=���������6�Cs���=�=���F(�R�G�����4=�u��u�m��2���^�����#WS���E��H�z�n|󞹐5jhW�_W�����[��z����+7ڪ+��k���\{���]6-�*M�L���D�c������*�Q�����3���u�����ӟzg�n����W~9���>�]���+�s⤓��I�#�V�8����ׁ{v�ur�Ȩ׵���2ƧB�5�����󝈓p=A�k���O)��}Wcܱ�&��I�z�������2|:MGs�zX�Bud�5'��=#f�z棲���y�«S���vQ? U��}�"�]�U��^�W�������L� 4���R~�����c�C��N���,��h�\^�L۾��x����9�Z��ղ�&���ݕ6?לϳ�Ǭj��;]�5S�]0)d����B�� cku��l��h�F�EJ�����Kx��Q@]�>R��/^Z;=���*�1�d3^�#=S���������ر��mh�!'��Ó�g�ץ�xp{����I�f���)K?o���г� �u���\Q��M|�:�'�po���U���z�Z�w�(;T�dO٩߽��yNO���oM�K�׫��o�8�v��	�<Wq��<[�<tt��=�
U�s�nҳ'D���8?�1	��c�T�H^���X܆���s��?ƅ��_T'�ym�z<�nY�>��;��P�4��`�}T����|0�~�R���wa�@������yי��=��7�s�)[�W鮽�{�;U�^�^��3
�ؙF�$����`LT� ^E(ڨNϫ�|2g��EGO�4�^���n��ƭWv�0��j�:�U �6C�!����뉨p)�D�a^/q��E�6��=
�[���ģ���*l��v��X+޿_�B����CsD���zhQn�.�:��g=;{=U;��HkVw�K �}��s��Tz�g}�:+�~��\�X 4��`���3$��c�a�w��O�U�~�#��<�ϗW�}��W�ix��w�G#ޑ��{,��T�����3�d$+Lt�e�*L�N_�wKhH_�~�n
�[�$^*T�bhÛ�/nؒ���2��Qv�G;,X���6����a�fp�	��H��[�I+�QT�@���+22�ޜ7�����E,�$�mЙ�۶js'm�KU�YH��.�峸��%0��t���Ox���Zw�����~�.�ay���ĿV��+����n|����Qރ�ޤO��-�50�c+���U�u��%�q	Փ���_�ǯ�8Bt��җӉ�ܝ��}����z�+�7�L�50�r�L+��t�������x�Rj�-��~����=�Ѿ��ޠ
�n�xx��$���ٰf���ɇћ^�97Ƽ"|\�\��̢�(�{�Ϣ/.�{2�2<ꥑ{����˸xQ��%�ai��c.�C��ˉ�2�ڲ�ɪ�����j����9��LZ�d{��L��)��ߕ5rI�7V�ܳ��Ɩ������gO�2|+M�������`uƧ�����>���nF��a.�׺��C{���1���O�}%��3�{5������ k�+ك������������r\����]�õej1q�%#r^�0�v�����2�[��I`�ꆜ(m��u{��v�}g�ޯ3����WhhϽ��ȍ�*j$���MCk�p���)�	U,���/޵���@���n�;5��&���^xP��|����^��l�����o���(2ZD�Un�P�F��!7m�l���P�Zpm�H��+V�q��=��u(=��5ފ΢^��NT+�i9����{|��i{�]�=��'��R�usF�m�(�V@{^�T�����k�[�ձX��=9UD�;�tXH��U��ӷ���d$��^���_s�}�l�.��V%o���z�9������|o�~��9E��f���c�|�^q���f�C��R�g�7�Ǚ��B_<W®��c"9����騿[�w7;��5�{�+��I��Y�����D��#e���>���g�y<T���Wz�\��n��_�NE�x^�̂*/������10�WH����� 5�����z[<:tq"��v�=��|wi����g�ܸ�_}n�m�2����r�㻑�K'���s��6	��u^:oz>i
C�gǋ���*� ���E}o�Q73��3a�͒{T���Y={��s'�WG��Jt&1���7�<�����I����N��,."���VW{�˯��y����̜�#8^'���\'ۻ~�>��8�{n���'-���x�A>y���֣��^$g���6�~���Zo\�j���%~��ȏ:׈���}K�~q�7)J�+�ɸ?)e�%b�\cWw1,߸�4��WP�x��s�PŖ̗{�2�a��6w����:Y��^r�-L�X��Z��ٜյ�&�:K��s(��l^�@����N�@�XL�׮r��-; <�����vN��_S���1�r��O�{��C0��='���N�<���.#6kM����[�5^?IEu�e�-���m��N�>�u1�ʐ�{�V��=�r$���vnra�g��� cpt�ꆷ�j�ե:���7��{�;A\G�Z3�E!q�%%�=;P�}��̱�T�l�ȯw�X�D�P��v}�Q��U׫�W���~>]ˍ�p���9�(��'����#�[ͿE4�x���;�FL�>�+���ua�@�^��⸸�O��:�q��l��P�=N祇w�ؖb����:}��@�U '�~�y(6m�ԏ\y?c����ϽV����h�bb�k������y�{�PY�ɝ0��F����L��o�x�ϟY	竅������}\վ����3�V쁉Ӹc��P��!��'�7uJ�T�Xr	h�T��q�:��9��K#�<hc�Mu ^G�	�߳�#!�5��R�&@l�֦�|_W�������|��H����l���\}�w~���=������F{,��T�Ișaq��Ǻ.�̽��nJ�����B���6��W��&<Dv��%�=Rl"k:6��UCqD�r�n�>*��e�l��vbG3;'w*��<�9�.��U���m�lq� ���!oY�Պ��N����w<Jl;u�u�-2�3Jt�Z�W/�LA
�6�T���
sr3�{���;��[=�~'�j������O�Y��>���t3�Q�<�����i%�;�=%�&�x��W�+L����F^���Tm�^71~��9��#k�蛕/zĵ�*�v�����D�NI�=q7P�N�v|6J�:�Z�c���^��W�Fo������r,K�F��8y8TY_I|t���FV釛>����f�/m�-&���]�%��s��g7�����jNCTGTG��b��碴yx�D�GN�;;��f�iw��)ӗ7�����y�ϣ6�_Fs�`R:y��E��Po���:u��&�� -��p����"'�:�\o�ާf��7�5>�׫��o�8�v��\$o�<W��<{�oh��͌����2zZ��K�rz�Td֕������{�cq�_����+����n㣧�Q����m���ax��'�o�8\U0'��b�ɝ~���A��ϼtdG����}���J��cG�f��3hvez��U���/m�af��$y;L	��D
�<��T�1�|X������.����Y��Z�6��)�W�ۻ�J��b���
������
׼�c���Q|�ٴ�v_1-R,M�RL�̋�Ӟ&V�W�=��I��l�<�Q�U���J�'#��Ov��=p�,�q�)�qn�G�����M�G���ye��Հ߬{�KG���:��<�c��@�;���8ܢw
�{�|]Uv�q��u��pQ�BI\{"�#c�����`h����V}
�2�������^�z���z�_s�}/��uAE<J��^��}�S;�8:�n�\{�^��馎����}�i�\����ʡGҙ���~7�{���W�7���Q���iw�
o�^���������9��{d�����ba��YN{�@�Xs�FX�o����R�Lg��O�;�M��{�Y�ީ�� u�_��%�%�Ʀlex���h�F���e������S�~�Ov�����Y�ѳ�'��P=TA~�'�ᩇ�9���t�����ϒM	[�Y⯆��<���6�1~uE��y�Yr�xg��*<Ĕr�e���ͅ㛓�`�����:�RG�U���}��L�����}�_�n�|C��Gq^ʨ�]G4$�����wq�3��RM�=*�j�۵��읭��4��q����~��C�ֲ��G�kݝqW�m�*>��~R�lQ�$�3���]�f�+PY�/Z���=�6Ҽ�����.�r��$(+�m�{���֓75����a�j�'&�i�����C��������F9Q"
z��6D]���{�v�}��=�ẁ�3j����y,T�JK���Y�D֊b����ǿX�b�gv��Il�V�0��!V}��Y�3���;#��y6�{��;T��sZ�v_F{Ko�R>V��/�9�ߝ�`���vK�5�����d}{,vj�x���[p{�ޫ�Zp�G}�ï��;�(�0JD�n�?�WL_�3��1�(�vi��-�����g�~Z+߫�'����x��rǪ�1X(r��=5%���j�w����yz����Vnukvw��UG����\<�s�i����iS
r�=�@�_�;�=�17Y�1O�k<�������W�E����\{!z�:�#�����+��p�(���{<����.+W*}��Wr� ���R�FAR�7,y���B�x��_���1ޅ<ˍ��r��Rn�WX}����Gk��O��� �a$���_��ͅy_�:�x���Z��M��0���������G'=�#W�q�ܳP�A|U����}t����W�����F��tL�E\�IT4�䄥hk�,t��}}��Y���ٔC�y�3�����$���*_?k�v�G�=��-�`m�BFl䜠I��EN��"�d�A
x�tb*���b�Oqxl2r�ٻ�`wgn�D"��g[ĤH��;��x�{�]�������/M��{ƹ��Z�h���g�"ˊP;,dԆj/n=����f��c�A�i�Zo�������=�.� ���dT[�M��-�3a����I>[��n���(>����7�nғQ�����/��b�n9�͟y���Tz��$��s�V�"���$0�aD�fԿ2��Q4xw�6�{�8X�2�t��<ˏg��Ә��:k�y�Ǖ��[�����[R7�ϣIG��?3������FN�Ӭ�k)��^��jq_��o���~rգ7���9��,��*�\/m�1��=�Ih�ه{^���l֛� o�:�C�yF%)�LsX|��M���X���:RCܗ��=n�w�P��xV���Ew��:�*�᯲���z��Ƭ�=}�6M�	wݵ��U���"2�߯ĭ6��|���#�-Z)�x'��Bf__���?V�I\37/�=��v5���V�Fx��ƽ~�o�����\o��ǜ7�l�+>�U"�i�t�<��[Y�y܆r�1 ׾�@M�\+ɕ��϶�x��X��������/�/�«W����3��+������E��螐9����^�q��f��ԏ_��B>gz��{��N�-��&Q]�峓 ^�[xxv��5�F���xd=6\:�ܞ��z������pr�=�5`�
�|x��k�#vF������lu*�!��v�1�/�{�����HEE� o��um���i_d�4[Gpr�Zz���?qΧe5��eC�rG����U��g�9E��q.�|z@�qU"IH�7��s��B���B� �_'{���%�Xs�=r�؏H>��!�6�G�!��7�J�T�Xp���˩��R�f�����K���k�ۈP�W�#�{�H���4_�ԁ�xT&󝿦@l�֦�05�D���s3�ǵd�z�ϣ�-�0�W��Wi��Yϗ��/�l �<���uNT���oe�'�a�/*�M�3���ܑ,����9�^�o£�#�W~8}:Ϥ�r��.�z��_�g�{�*H����f<��M�x��_\�2+�s�=�B�;9ظ�s��~�*D{7�"��D����mo,Js/����n<|O��D�qW7P��n�y>'Y�gW[����>�޻�X�&j}����澽�^�n�ҽ�C�QW���`�<��>�����=���%�������v���J�^��^vx{�'�K�Щ{ۘ(g�ਏ!'N\�gn>��xn#=���n�;��*v+y�v�}l��v}���b�X	�#Ū����uж�V���<{"g�4���o���jM�CnÖ�g��V���WL���*��|/-T�Z 5+�Z�+0:���3��[�Z��B���ft˱��u�	���I`��9I���AM�"r��<D�)�fve���s�.�
'�K��H�,����vp��N�"����?{:s]�U4p�,a�Ж� ��~�<�HkÀal���;�I�gLur���3�ݳ:�E�2C\ �ِj��e(�r�l����2/;6��A�r��ԍFyIP���z�"�Ĝl�`SvS�^�jy���ުa���Jf'���5��y�q�^�����I�f$��&��c�
��53�VG݁WdXr 4�c��K����v��W�L�]��p೬Pr�Rm���fV9{AKF@_=�֐]g^��5K��\o:�ch�����&�M�RP@Sxخ��}�
b�(D��V���]&�Wnj�n�)uobl��Gǧ��Z�}�s��8��.�7w|�KɆ�Sֱw�X��X�}ۓ��#PUu.؝\�N$����v��j��tf�	��MfA+!ȨKUԕ×OQ��=�ӕ�[x�e�����n�հ����0u�
��a>���[��K�鏩��-�볻bU��ؕ���,�m<s!`���ݾ�4;{x}t��r�wXw0��S�R]��;�(',�� �Y�R'1EY�;j�;XRN��vwU���w�s�@�=���L���oU�`H?��O.�Јk��xR�;O����c]��KU{Zp����8�]%�g`�@��jɡp�R�i}��B�d�Rnc��<#:�]b��3]�r�̣��8�5�9R|4�>�G�	�s��CR�5"۔u�J��8�@�ʒsbo�` �THr��	��Wd �nj�u���p^�|��|�>�ظ�Aѥށp�0�.��&h�zl�R�*��k��T��s�i���湵"���[:�m9�#-J���60q�&Y̟_oq$�;��J�[��7Rq��A�]Ӯ�ew*J��x�	e�|���6=�U~B4�D�e���R�{jN�t�b�z���Jx�3�n��1$S2�ffo6��盔T�L̔4u�v�aQӛt��G����v��Bv����1���)�s!��
r�,i#��]���^޳W�JW�QV�H�y�Q���Bں�/�r+�l�L��b�:���t��%�82�D�l^:�%�l��b�`=�z���q�wܯ��N Lw/k�+�\���2�#�����?���>�.�wn	$���C���\0)�H���mv�i�we3��������xwz��6#mPL��E͌�����H�X3���sZ����7���ܞ=#�׽3�|5I|��"~*��ITZ�:J�Y����:I�ib�AE(����Q*8P]-
�z�9Ty�\�	��s��۝/[N���t�(���,�@�%�DNM9N���UA�MR"er�%��AT\*�����O\�<����sP�9U�W=nN\�3�72"�

���V��ˑȊ��9��
(�m]��9t�tӗ�*#�A�e�! �!B(�N�NYӔQUy�ejNE	\���r�]�HD\I�	ER�7$��"
��d	ЙqZ�4S/E���������b�^q�ЎY�Uª2ċ�L�*�͐DvEU�Y'(I��z�"�c��L�ueDE]8�rKS�D�滹:!9(T��p�ԣ�&��EEʪ�b%ES���?��'���؝�K���)�\[�xT�cWҦ�A�>=Ǯ�ZF=9R�o`����jZUs�t!�P*{�$�bz�~��Dem�_�)\ޟ@�����^�~�Z�]�pٴ�G_��(�u�ʏ;cr����j�p�T};8�*�U�Z^���r����V7!�_��m?�a��[Ak��#HǓy|��uK�T��F/C�'�Q��8JF�Ӏ��0&�X������R��>��\�˱,���V�6�}\W�;�g������� �$y��T��ȁC�W3�'��h�Ǿ��ezҾ�w�G{4��`��KG�ޯq�WH1�)��;>rMA<x�8M�$��p�G]��73��|��/�Nv�A����"���{������_{����S�Yynh����w�xz�I����b�wF�:�j�8R>���P�+���z�9��!�F�'E}~�r=�Iz�P>�D׶��/ �O�`�u_��>G0����}��R�Z��Nq(��x��&5o�u����ަHؘ�^��D�9����:�c;��l/L����1~;�Wo>E����_�|�/�K���2[���ND��\�C��SU�O����\7��=�)zY[��Q�31�]T{u�4�T�F놤8�,���oK���u�k9]�Ύ��X�D#�@�	P߶E_�oqLd�l�͆�MD)��0g-P*:#��B\�خ�8W�{�\kk΋;Ȕ�z�)s:�ѽ���H���!N�L+�nW+��]b�ê�����fi��v���~D�{�:�r���6���"����'�a��+[��LD%�����O���w������с�ǹ������/E^bJ9q2�m���cD���O���s�6�gR���F?T���~-�ׇ�̢�����̇��0�	F��w	�J����^���L������*������Ƕg�%���^����Y*?v?C6���Qgߌq��ge�}�I>�YCO���5�^O�i�r7�gK�#S�~��x�&[L�봖��m�>�K�\>�<c����O��Ϣ����kK�;�k�5�C^����/}W����ίW=�^g��^�ք���1f	H��ت�㊥��ɝd}�+��]���][\U�ݻ��W��s�3޹�����9����
��,r��3k�t�������9�o����M�V�S�{3�Q<���D�w�Ox�ӯ��0��)W��)�,��r��&�,i�f�M�/ڡn(dS#��j��J�of��ߺ��/Sg7�<W���7���le9��[��o�*��
�8���31�mDФ����^�^�L��ww���ȅ)YȽ�'1���V�\^ɜ݂����7թ+���JS���L,Y�z�'7����E�F6��8;����z�j�q���RMVz�ME-��rmЙG� ��5�w^�\�M��wVC�T�(~��\�u�./���ϑʓ��ݶ�=��'�@h�A�	9Rr	^+ex�}^��ح��b�-j�ٙ�~�\�.�Vx{�մ˝��=�T[�n-���ꋤLS��%��u+�#[�^�:+ݷ�B����Ѹ�)`��� }� LS���l�̀����0�}��r���V/Q�#ݟG�C�p��p�yU��9�����ȯ���&�|��1���G����r�CcC�۴G��������)|n�Q��5�9�z�(ۙ�0�4ҍ�z��^{���ƱG��~�:�&��^mh���e�34�X�ww�:�s�<o܌�1ӭES�s��n^�*[(fNuz3ò���?�Ӓ|Ν�ݓ�}�D�Ӯ�7L	����^���穪�,���_�>V�x�\Н�=�pǐp�Il���C̟qaFl֝d��Rr��l��l����������ڽrFD/m4Ny��,�(\>�Z/�Ew���:����ja�.�l�:��n�t�J�3$m�a�p�+����j]�ңqhKshΎ���c���B������d(7��V�ep�z�:�e#�9��D��s�&��?1��������Nް�ԓ-���v��Z�`��]�<��l.�z�*�Ӈ�gH���]����L�������q�y�p�䠢3���g�{ў#��7}/�g�Cfp�HW�P��L���	��wq��^�q���.7��c��QT��c�$�#ӝ3��������3������M���L�>%x�sA8����v<_��{%��F]��ߢ}��vn{�X��u��2��Q���qT���yzM�ٷ�R=~~�=�O�ё��F����I#;Y�S�]�FA�G��>�q�\y��k���+���$�x��^/_Q
oo=���o׸��к:�
�N��k�M��p��~��F�j75��T�Ȃ�K�w8�'��;W7k}�/�ί}��ｖ��p�ԑ����/7���:���W���G��̀�4��}u�}�N�>�Xp�Gw�����E/�]o��������ܬn�ʓ
��y����P�J&�TD�)�;� �ӟr�|q���L��o��}��]���y�g���Dw���҉�9�t�_��!�\�2+�s�=��p�������;Dg��9����U�ea������۲�;tΏy��*��{=P׷g_�E�^�[p��
W˵j���j�W"f�߭tn�ɐ�]t~�q1��
�쌡^�lpF�)O�,��]�u��X�b�#Y\��5}G-7Xc��gi ��E�0ҷ��w>[ܨdO]E���O����<���R��՞Yc��h[��u9��Q&�����w����/�'ä�:��c�n[0a�p����Cu~�xn�U�m{jǲ� ��<����K��ו�a�m{�)[������^���ug��� z=���dG�T�'>�;޺�C<�V��x�-؝�x{�F�m��uU��sY;N32g�O�鿣:��V<!���8�@�Q�ա<��$��܁����U/h����彙��=�������ۏ^O�Ώ����5������3ݱ��G��Ep�P��׵FOc��Hu�=cѽ�C�NN�>�ɭ.�g}1q��K���46�����[�h�n{&&�U�{��\���Jsp�L��+��J*�����=uL	���c	��[R���wa���#,�{�}�Z�U�v�O����{c�^�q�\n}�m�Y(ԟ"���`LT� U�EDoo� �Kƽ�}A<��Ox�,B��z�/Ah������5LUT���:��t�p=z���׽��ѯ��P�?0?|��������Q�����#��{����S�Yprf�Օ��f���>�T�D��:uӺ���e]�v!�h$�,�ߖ�Þ-F�x\��#���-�O�̀�ڽ�I��K��ʬ >��:��'9l%|�%ռ�W�;8l�K%��8�g{�u��M���{�%]��z�u�b��k��LslX�uĲ�^��2N�۰���,ˮ]k����WM
��L����!��F�x��5^�˃��S>�c��~�d����1��q� ]�Nv{�ew(^�; [>�(:�T* ��9����|����[��OS�_N�(�_g��joE��n��}y�)\��DE�ٟ����z�&�.�3�9�}+N�X�oև��r�jU��7^��5�0��53�T��<��9�I�s�-����ו�b~��h�>�/ޫ
EKzLc�[�^�|U�o�_�6����>t<�>�8����?
@�L����^V���6:�J9���O��w�'х"�گÂt'��7~�<��s����$��2�o���oT�;�Y��Ͽ$�%Og��ﻶ�כ^�q_5���̿9�d/uA�Q�p�\�9uu�Pk�zTϵ�iH��%�g��N�q��{�N�c�3xX�����e��%���?MH�d�\�UibsW>��gm�/ē�{�JD�1��ZU���Zu�����`uƧ���d��)̞��Ej��F��,}&���ƴ���+���b`����[K+K3�7�{^�>��pd��
Ȭ.��B%n�:��B�VWh����������ۥ������W;���:�S�T�"�ާ��@�>�X�,Q�~a���t�\�j�i��w%.V���,�Yދϭ�aAݞ8��d��_���z*������ɴ��nf�AW[��j����QU�Ѫ�$_���y���;#�l��%#IxO]T?U,f�:W���~��i̺�������LǺ�ҳ�.v��י�exu��CF}�h�lL�RXJc��ȣ ���WN�v�E���W�R>٘^*'�\<�ν�#})���g��S����~�8=ꫭ���K�P����d 2);�7��v�^	g�\{�#���Ѿ�q݁{��&��������^ꠏ��GdSꑐ\�M��w>}D'��WC~��9��"�MD�Un�c��Z���`�q�t�5~�p��+�Xόȁ�:Tj	^+exڈ}^C��wL����idOK�{3Ƞ��ў��\F<�"��L�,�Ah�����]"b�O���#qꨬ�YuǷ�	{go�iq�Se�Ԫ�s��
�� j3ِE}n�m�D�G�&@|i�nOl/g��T�l��;�=��R�z[=؍G��.~�}n��#��z�R *���o�Y:��,���I���r��P�K��lp��#��d��Q�/KN�F��=�:��:��x_)�S���jj�G��U�[A|�W����xu�~qm��-	��S&k����w��ؒ]b��Eܡ�Gm����-PӁ�@�B������i��5����Wu��6qi��jj���I�Ţ��؏
�A�G����;�eMY|����#�҉������+�6�<;�;�ƙ�ŏRy�M�O�ŋ�H��5���z�h�s>kn⼤��~��Ӓ|Ν���N���d�7��3W���{Ω{���T�mFU��瓽:�І����5�{�gL_��n$�v�v���W��f�iJ���f�o�+����Dd���k�����Kd�:���\4/����=�n$�
YU�9
)��~��˭��FfJ��R���|�������~yhp��((̒��&�J�k�<��]��N7�y�5>���3��^L����	��wq�O��w���v��c5���C���˺Y����P���s�x0z⩁7޸w�)φ�^*yՇ�]{N}�K�h�~s�j�}_��s���d��U�Ưeyl�(��޸�`MO/I�ݤ9�:=��C�}�sQEAG�3��k�y!�h�ir�Q�r�0�!ĺ4z@�qU"`��~+���>���c�ݱ�]�#=}�����z%#�����������*��'`7uJ�o����+����%�5)]W�,d���A$���-cc��·k)�$r�i��l"�\6���F�C���g����7%�2���j�~-vS�]y�{�VSi�>��������ٔѥ��Cj�3K��IZ�2�WZ݌����ۙn+��x5@����3ܦ�.��Y�d{�d��P��/,��)#��ש#��R�o��p����ў�� yK�.LR[^���ЧTxgћ4+�;���>�j�k��]o�����^���}�:��y�;Y���е�ܟL���LZ�%�Ü��8�^�i�\,�*�Ϥ�\})��=�ط��3;�/F��*�>%��Go蛦:��C��V��|y�rv.4�{2�댿C�z�n�f��nc3d{�ީ���5s�V��O���n�����.�'ä�k�~�6�S�����~}<���w�/��d�~�a�dy�=+�h{�� ��V��Wݵ�[������d�u���:Gluk�K}L�5Kj����_�G�T�'#ʈ����P�=����9s-�+wo�WT����i
�j>�uT+ͪ�z_�M�u�Db�`&m<�dN���T���+C�>�+��PU��.����U,�V�Cj�kN��+O�^�2v>Y8����w:y�`]>�������B?��VnC�W~�F�0�w��է��3���Brw�Cz�.����Gw`bz�k��H���HT�����k���5|�g{�\���W,���N�G/�ʵG��a��Y��<��<ċ`(�֛���h�(!��u�\%a�2�w�(l�/5H��hA���w.�W�w��#y��Iݗ�i�J�*�����ۏ/sJ������E���{#�s��Ä�K6L�:�X�ɝ~���A��Lr>���g�W���<3�|�粟Uj�q�l��͉�j$�7�Sjy�G���2���Cr^���;
��綪<���Ō<�z3�%���xs���8�d8�F��;�5Y3�F�Ν�k��{���O)���_>�(������x��xwo΀��^�7�(���/jfYk/=��w(aT�	�s,���H�h�q��E�U��i��"��A���cb���{咭h[������n&������}�X\wz_��*�N��gu�62�\��J��ZAj�ӄ����DO�꜐-�0��t��s�:0�V�@��n�ֶp?d�.�V��h~UN��A����D�r�{.[���NIh���C���14�m&<,��&����w���o����U���~��E��l�B������C�,�g�U�u�sQ�S��#v�r���j1���Rk�/O�����'b��K=�:�!�]���E}bJ9�D
������{t�ۣ��(6�0uV%�1��X1��wّ���2�զK�6��֨G۷�Q��7�'R�/m��*"��u�vs��B5�zX�E�X��ֳ�-�Z��r���P�T����*�`��X(N�eP嶩�"�����Dv�Un)wR��ؕ�g����S��Va���v���H@xC�`�+�/"��v��;w�T��ZK���&w!�����c�Q�%��(c�Xuzv���z^�ۣ�rG3	hc�<�N;=@'��5q���Q���ݚb��P$�+S�Lhݹ�'[)���Fq�]���;;{y.������h�����>�+�=��>ƁcK�,5*}-�b�;����Ռ)�Z!={NS<GPǮxA=��#�\�9��Ɉ��k��T3$�96�)#K�	�Խx.�Ԁc���d[�)נGjf�#^����O��t8qGQ���m�[v=���$�p��Wt�fo%����uh �˾�r��K��l��(�hV�*]7�TZ�I7�c����o���:x��5�K�h{�h��:ڍ#F+�fJ�{�tn�lDq�屣.��3y�^������I`�OX�X. ��9����w_����ܛA�v{�=M�\9�++fX��@m0F�"�͗@��.���\dn~췲r��d��!�Q89x��nx���;w:nE��u��+e\�t�ܾ�Y����=ṋc�#�A������(\���"�~;��k����f&;ꋓ�Gn�
ڜnn�4�f��%w47�K����|����w��!k�گ"]��Dj:����%ox���7��СE
;���[:�k��o%u�E�,�z���gWn���|W��3�$�qÓ��%�Z0r���m�]iw���vgo:V�q���+�l��zǣ�"�W��7$�r����w�W��eixQi�:;��jԀ�9��A$���.8#�"�ma�\^N�)�(�L���U�;VM]��NG���/���*}�?N�K��Q��ٓ���o�;2Z������<��� �R�{o%n��y�3�>�kb��өY@�ܮ��V.�n�o����)����{{��x"�>�iM��Q���r��F(^R��^,Q��b�y�m�Ngl�{yt+S{,�� Y�q
,���Y��sm
��LY@r�\i=9X�.�]Z����T]�n�ؖ�Z�m34��dݢ�N�&����Q�K��}�VMe�Ն�Fb�0}�Yݕ�Z�ڻ�w]��mҬmXE�uR��s�.�r9\��MX���u���#3-4:C�7&��� �Ԍ��$���[w�q<�\�Np?b��wF�8�t�����O��S�9�=���y㰫�A&��-)QO��8�5�jʏ@���$ml��t�g��iۖ��D�*��&�L��#���(b�3%n3�ɹ6�b:��B^4��gSZ"�%fr���د��2�ΑL���s�\���l@}���xUAE�^�᧭(�����(
".F�+YI�
.BW�9p�,���*'2(���r99����IيG*�(�bvꊜ�]����g��]R*����r*tD�2'\�*�Z�;V�9�s�$Z��F%C���ARan���u<����r7w�*�����Ktj�;(���(���(#�2��TI'�NwfD�W����L ������QG'	4�(��"�ݧ�{��d�(�;��N)��uܹ<�<����TG�E�M�c�Nt��7E]�T�n���TN��� ��q<���
��(��=]��'<����u4u=����ГwC�:��-B�-55�Y�+��Ķ\��
��Ȫ!6(���$)�r']RB�̹�T!̂��wYD�p�d�����j�:�{����NY�p�%r!P(�C�(�����0��'�a<��ZXU���$�R�n�ڸ:�[�&7{��"�+[�Y����˻��[���Qኹ�Z���c
�9<��R�V��n��B_�69�0���|o�/���ۇ�p�����Q�b��<���O[q=9w�kv��ﷄ������ߣӁ�\�t�ic�3y���W�?�x���
uN{�-9�]�'�;X_����i��25_��j�>_����\�OJ��<9�/����;���g��k��g/e�^�Z���o�|P/��TrUo��(�C�=��YK���3��'<rڍ������l;�W��ؼ� ��n��5׼H����=��u��hw�QF.��$;'fax�Q[>�{�skϵ-�{���|o����m*1���o��ϑ��m����[2<�����5�/+�_����6{ô�Q�*��D�0'�]p�0��y��B�<��ƹ�o�2����հ=���(�4������R������9M�`LSw�p�Z{V%���Y�ٽ��=�������g�ۼ�[>���e�M2� ��= r�T��D��X�:�HI�����
��N��gUR�J��^�j�I���H�Q~�p��+�X�0["7��Q��W�Å��l�X���g��������d�Q'��XB�_'z;��h�5m\bP��F�&���&ƺ\����殑K���/����{z����U(n:���7�}���z�*g]c2^�l�G�a���
��@:R�m��-R�
\+�I���k�5`���-&���oG�{����lU��Ze�aE��H����0*-�P���0��H�����(7��=����U��>%#���Lz�ަ��U~9�L���=wl[�@��G�:(��(��28f_�sS���3�וmҙ�Ba���+�Ǽ��r6|�=�6 U�1d��s<��i���H�Y?���>*>�ds���.�{O�o��P���q��l�{΀�#�샩��~�+�ǩbS�G�^�I�咷 ���ܰ�#6�;��𚍖4���c�	�dz����u>u�<�n�-�۾ɹ�}�⧊�۸�Y�*=�K/N}'���ׇ���>���Zn>�?����F���O�)z��u�G�G��sʏ�vU��~�:b����q%���.2�Ō���H�z�=����U��}��U�u�1M{�G|���9uï�,�([�����]�"O��kb�V������-�>����Q�]eG\F*�;�{���y�'>�s���u���Y|���HJ�P3�гg�Żؚ���F�:0�n(���;���M�����ƽ~��~/�u�U@�to��H�.��>����9dݫ�L�{�����_�̻n�]M�ֶ�չ��W�3#dN�.l��_��y��Qۺ�Դ謁�c��e͚��e�E@��+|�ޝY�	�V�X�b�MJ�I����RMT[���w���9>+o�SQUuyܳ��P��=	�Vl�*�ς���?_z��d�s�W��4G����DWc>��{֛��������#q�F_=��϶@�jz@�\U0(����%�ڙ�&�?:�T�m���J:ތ�å3�>�pt����Wί��r�1��]��+��$�x���߽�y�d�h*��nx�/ݧ;�Kw޴���1pw�]Ƿޢ6�^�c�3Q�Z4K��&�K�����l�t��rc�R��>%#��}pUC�Hп�z�9�u ^F���W�w"�������*TU6�}�ۉuf��ڕ�@h��jhW�u{��Ba������~�^��tq���(t˩���o�;+�B���Ϥ��ÿL=_E�"i�i܀_���2��7�Q��+�O�/�"{l��L�2v���f����`t�~�����7��4v�n���Q��Zdk��ބe��9[�qS�g%iC�t��rJ
����7�>%�>�&��ͽ�2|:OSK���
��V�h���=��:q�3�/�{�D�r�q~�=6��c��EG����_�څ�Ӛ����z�tp����}7�萳�y��,N�h�[��jV�B�ͫש�A�+��[�utŪ�12SUo2�M@aY]�lC�s_o`�|n6�+ow���N��W�Չcmigxv�A�A)��8�-=nգ�c���SAh���'\;�J&�w�m'ӵU���=���X��׀���2��)>N�r��nċ��pTy	:p�~�l,�mQG�2ai���צ�`j=�W�}P���(ͪ�z}�ӝLح�	�GOCWM>κ��s]~�=��V;�`�F��g�e�s��^V�+��,����zd/W��d�/�#~蔬��UZ���g�3�K;"����#���o��V�KK?*��C��Oz�n#�|Z񳛦�}w�B���-�x�;��7�c��-����R%����7=���L����99DR|}����b��H�D�]�dq��������G�����q����W(�I�3,��uP��f����3݄
ǽU���`k�`��KG������1Nq�C��w �Y�~��x����Fc�z"���q�x�ϟ\^{�<�?Sg#W��ޭ+޿_�����P>��O��=�xoV��x��'�Nn"�4*t�ݖ���Tr/��u�H��#��^O#��wO�s5{��ʏ!�m܇�Ij���`���P�����Ӌ����kw��&8Ϥwڼ_���RJđ��J��y��*�҇������$hۉ�Qt�,�T�mπ�2�����viF�,v��Qgr�g�Q���y��}S�B��Н�0�ITʘy�8f�4�k5��D�tīFwd��pΨR�f
�aW�rI�\)'���b�ď�	��pU�ߴA�Um�
�T�p�G�&&�"�4�t�"GM9u+\�]�e{7�YK�G3��<^W�3�O� W�fA���^%rZ;su�2�L>���P��>Ь^z��=(wg�5���[�_���� �z��3�7�L�.+:�Ȝ�S��vs�B�j���c��ѥ��\5~/��dC�Q�� {��P��������ܝ£��W�����@��3���fǼsrc���7���}{p�m�����l�~�A��H���	C�Ms��|�ag�g�e/��o�|���c.=8}yU��K��:X�j�lz�!g�q�G}�v����e���>�]Q�����~rI�7>�6�i��ɭ*�|+M둾�zW��T���T��KE�������>ٶt�z���b����g�_���9}�VU1��ZXN�z��xq+�T��ΐ7�����^�"�_;�)����e����b���n$�'�8Z��S][^�Q�����t�T��L����vv��܅���:�=�{+í��3��H+k�;;&]9/�g�m�s?tR:��O���Nu��e�)h�,j��
6���#�q����l�kb��Hyl�{zL꼝���C�qq��{�����F�1a�y��w����׷P��5���_�7;��]Hl��*�1��ͧ8���y��({f检��q�2�mT/�W���Nx�_o���q�̉��x�	�N;�z�{�N�{��.� J�:zd02���2�ڱ(�~W��٩���Z�?�"�׽���������p�_t�q�׫Ô�^f���}R-��c��C�!m�iSK�ağU�W���%���y�s/�a���=�⋓���0�U# ����.���#:��d���u�3=z{��L;��b�"}\���.s} k��d_[�n-���^����WEA�z�qW[��&=쥧6g�Oh>���H�dz�_��[Ǧ�~�S��]������P����ۢ�B�Ê=�W�@�5��11O�h�F�x�b5M�~���W�|�,.� �)?L��V�lw�����Ah���,�XY�f�y�B��V�����B�M�И���6OR���}�5��y����}wq��%�6K�M�
�kC�������ɯ�K����:�MD���{�;ǸQ�.������O��۸�|Q�q��YzH�8r|??�kG����E���P�d��l��~�'�Z�rϗW��KU���F2F��8��Ӧ$"gK}�!�Tb��T�X�MR�v����^�>S���L�\D��B-���a.]6T޾r�����;�5��^�y�2ݼ���q$b%Ӈޅr�b�q����NK���n���P�U�\J;m=_����e����U�/N;@�IeG�*�_��t��=��v�j_mr�#�nv{K��X���~�({6kM�H�3��b�~��W�θuǖZ/��+E���r�m�ȿ>��[���ǲ��}U����׎���mT�͌�l�z�YI�^N�Ἇ����z�z&{=��hu�=cݒY�P�ӱG�ت���3����	��'��nC^�q�t�ٽ���3y��椷������&}�%��dC[E�l�*�g��T����ü�N|6J�:悘�+���V�����ƻI�������ǳ�8۵Q��Yeg� J5�z�S��o�'սS��g$��V�y�Wo�w��C���=��������q�ȅ4�p\���+���k��	��eMwf{����&����{��Q��_
�����މH�Do�����G�)���nfgc��R�&��\�o(f~��1Gz������AJ�l��u�l���z��V�\���>l�|�"z������}�#ޞ����20��a�%����?��n�=O�mp<���*G]
��nQ���՗��E��V��Wt%݈��F�e:�w����b�qȖ��:�,�[XŃGf��ΚV}����Y�hW�Uw��T-%mJ�Tyf2]�;8���\�"aQ�D*�:bܖ�F�X0���*j��f�ܺ�[%�듻�Lv��������� �]�E}~���$���z�HqN{N��wN|�^��׍�,��N���3�}���P�]�lΣRo�@T����Y�0�ۉ�c��C�V�����Z �4�9^滳yBc=�^71{·�����>gĬ='����CW[�Ȏ�v\�p����i�R�p�>��`��xz��'��'c��#�W�?mX���7�	XnK�Eߧ�����WoJ��%�/F��^m.7�zx�� �J�~��T�'#ʈ����P�=��o��+{���o�ڰ%{�����ӳ��c�_ٵZt?��u�ƫv�|QM\4�79���34���t|��;���Z��@�g�H�,^���
�=J��`o��j}�#W���c8����3P���-_�Wmw�g���7��?v��m��M��"�W�5��L�/�r��;�q8�׋|�w�?F��`�����q����j�(�Y�R7�늦��cn��^�Z�����u҅]�ܟ}�>
�y݇�g�:3�u�{c�^�p��������J=|���ʘ���� �X�����������gV�������.:)��Mo!�$�^��\���N\��������z��j��V��=�Kb�[O{N#�]Ґ̠�ޓ�p�+��I��{u�<�J瓎�'��.���®�����e���3O�����[U޿���c><�z3��M��ޯ.Pc�S��:\�@�a��y:�L�#1C
�����5
�Oԉ��������Q��~��F�'�v���1��zǬT��k|].�`�*����܁�7;^�[��}�	����U�ԑ�7�{Ӟ���S5˒əbJ�����������Ϥ���=�UB���9������n��(@����v�ǝ��8z�>�>��Q�zF�g�Ȩ�T�"�뉉��TFS��Жm�ۀ�=:67�ɭ�e+ͬy�}�q���_�'����S��O� W�T4�7�`�~õ�[1�'V���;�;�ʳ=�Ǣ�����_�e�Nh�����)Ϣ\�������	�t�s[�}���%�&�7�#+tüu�j#O������q	د��w,��=�˻��x�z<Ȟ�ȷ�����|�h���o�>�l/�ڇf׸�}��3Q{p�[���ΪY��ڏ(�Q�f������6�}�۪��죆���r���ZnvX�~��鿴��y����<q?&+��dc�lIz5�k�Lռ@K�(5���1f7�7��rǺ�>����c���j��lK��Y"'�����PE�L�֙�|��������1�l�x��^pY�8��þ�	�֟V9�C�+0���܎�[���:�ˎptk���<P��Ʒ�9�3�w�Z;�]��7���&�=�gM��'��D�P��v�ˌ�Ю2|+J�׵�r���OUkw-xl^x>�i�6��<����r=��7X�)�Q�碻�I�YLd��>uRp�v���>.�^�����C�2��k�7�{,v���������~�f!��F2�H�R��FSPt2se���T�W��o�iA�(w� �	�̩�M�)�^ӜS9��W�Z��4�4JZ��u{�U�V�Qذ!��B�=5%�桁1޸w�A\c�^7Ϯu�9���Iǒ�T	Uw��Ab̧a�GU��g�r�<��o�E�M߁���˷�bQ���,�:�O1�w-m_�j̗�}�8����Zk�V��#�(����9]z�Z'rX�:�f����v\�Ŏ�k��~��~~��dw�Rg7�4���w�=5�X:`�u�G9Ax�p7��N}��G����GO����Х.��!�i�N����^�n;5��ת�G��W��mV�tgw����bb�Rӟ���jD7IL������?|�'��m�o��m�o���`�����`����6��6�1��`�`���X�`���cm�o��6�鍶m��l��m�cm�l�X�`��ьll�m�6���l���`���Cm�o��m��m�cm�x�`���m�cm��PVI��v(W��@���y�d���t�Q JTT�UD��"J����J����TAU)%D�*J�*�UT$�*�-DI(�T%)^��Q%JH���*	H�BR�
���R*�JI*$��kP�Cq�"�����*��*D����J�$��EH"()RIAt�!"AT�UTQ�UR	J� �ъ�Q�X2�0h�(Hڌ�%I��@fԊ�l�V��6��J�E��EHk�  �@	��U,� SVPj����@���wgE( &,
P4�w)�@  � �4��갥J@�Z�E
*��  fS��յ�i�E-d
AUJ�։l6ִ�P��j��
XU��#5)[��%U�  `m��Y�P6�M�� �I�J
�� 4�� Xb��U-h`-@։U*G   �*�ͨe5Thث
V�@4V�6ͳ+j�f�
�ŁC[bō4d4���ִ��Q���  �AZ�Ul Y�4*��CmPhUj� ���P(3XZ�&����f�5m�����U"���� 5���mj�P���(`�U,������ڍ�0�
�TƍVh*�`ҤI*���)� \emTf�- E� �ki��0Z�hhыT
4�m�4�4�LPQ��imh%M�1U�PV1CY��UU��� �mQ����a��QVXZ�b3Fh�ͭ��L�4[m���IY��+F�Jm�
hU�!�h�`	Q5R��I"Qhh�� ]!B4ePF�)Q ֪h4�dKCSL�5�&L3V ���AUT��?M2�RR0C  	��`&���$�*z��  �CA�#S�OL�mA��@ h  � O����`      *I鉦��5OF�R4h P$�P1T�Ч�5O'��h�22M=B�5�� �Ti6�!&n<`��@�t�O-�<�� 	$����d���C�?�I`N����BI!��$���C	��������֟�t�ٴ#�$!$�J��?�`$�a2A�R $�!������}�G������>�!	$����ar�&3'�a������,��@W�+������?�����N��*W�yt"h�h8�n�{�%I�%�n���D	�y7^Q(���C[�L�-�*�v0[jd���-�����B�r�V��<�ʰ������-�4uM���I5���JMvL��Xa�M���kC(�����f,op�u6���X�u��:�i�hb{� X.�P�BɀXT��h�OiZ�&���k*�]������ZvXUe2m֬��!�#]�y�ث2AZ[�ur7�3h��ɡR�E�	�l�v��6��HO�\�o/qi����VXubL����-�i�*��1�+79J�Z��e"�X�h�m�hGD`�V.�Me�'n-���[�"z�m�
�δ��"�"c�B12�����m�gv�42�9 �t3.�[�NlX�Mdj�kAem��U�p�[V*��J�N櫩�����AJb5N���)�� �ǌeޖ��X�orm���x���]5���2��;ZdW�S�Z.F��Y��C$�T1�h$i�"�55�n��Y�0�V���9x�-.��&�9z.����d�,#�n�52a��f�	�b^A�����EkǌU�jެ&TwE9����:�n��պ
kdZ���UZ(Iq�%�z͊l�Z�i�a��:Xe���:�p�9���ú��gpe ���7X�b�2���s,AKEʷ����ugl��Q��&��4
x\�sPr�[�	��&�h��k5C��,��t�"�l�0O�ͧ��$�Y�&*YN�/i]��;5�ûky<-���ێp��ifPۻ��+scQbL�2�Z�n��z���Z��V��9x�Sn�Cik�W�4(�Sd7߲��Dڻt3 ���i(,��V�b�r�&5�bR6��4f�����j	�5�w�s�N��kmb��~/%���6
 ��
�!�Q*EW�Fls5Cskq�Vi-���Z4�k��H�(圶+j]I���QT�$bHh�dH���vLŬ�c]��.��&etnan[6�=�$v�TӴEa�m�jX��5i2)��;���kj�I��q�.Ǝ�@2l��jAË�PX���j�k;��b���S�����js
WOp�^_ɼ.����)�$�M/	�*�m7�'�P�`%X�Tǰ�-aƓvt�f@��BP���yn�n|�W�'�ڙ���`�3�-�A��Uyr�VP����hU��ZVM5��������mP�7(��d�7�9�+e\R��V�)�PqX�N�,��
'37!To7�1z�hA��5�������oKq��-�`vV#�V2�b5��SvQ�KV�S6�a�R�b������vx��%�ӥ���6h�t�H�i��j)3U;8r��W�VЏJ�6���j*�t/է��w6l�­칮�ԫ"����)Vl-��6�~aij�Er�ș�t���щ̫*ȩ��i�?K|���JOn�4�~,ҸwXҞ����l�X�� �XҒD��4X8�խ�Vl��e
�j�^5�\�b�^GSuD\�NIX՛:.ZTp=�
��`��pͭĲ&��P�&إ�axq��fH�[GA����h1ޕ����:2��攦FnX7���l���5��aRSMe��;i��hs�2�)X���j�n1V�j��"���e�̊��Ȗ�#�J�ՂEC4�N)k��|!�xf�j�J25B��sb�)�Y���Z!͠.���2=TX�=����ʱH�.�j�:'�f���:��[Gd[��ܴ�z��u�5��bĩ��Mxu���o]*w�(�A�;EK�f��{�����P]D�S(eF,F�����g�jn����3�եU�V&�0J����U��<70JJ(�K�U���6�P�*�C '��4��P��ٕ/".�RS*����hMI��OYQKM5&�R�*A?���9)���x�ת��
F�'v�Pܛl]C�h�D�]�V֕NwqE����PS*�������0L�qԁi�d�F�������ouB�Sq2����Wb<ʌ�.e�uO�B�H�)�,�L�EC� ��1����6~MR��V���o��7`iԗzm�%m,�V�-2m���d�@�%�;"�IS٭俦�n�S��F� 1���1�%M��RH�:{ v��jE��BE�l;�6�����ij�s#��#�ݲ���)(zխ/���!�����@a4��Դ=/.ge�x��u���2�c@�)�J����l��S?9[�bV��!���/���E��q1��UŖ����Dj�Wo�uǹW��f������қ5)6E��:=��W���5����'@2nhf�lRVU�+!�8"��K]ͭ�-	��-KyLb����n���mК��ѓ";�0+��P)�Qf`��n�B���x��%�R��kKi4p��]c ݑ, %�2�t�:�
�2"ׁ�86茗���.ʨ��fdq�h��E*��&��u�K?k���F.��S��{YO�PU���6�Z�d������M��#��0�N�yn ��b`Y�-�6��nh:��y���3%��(]L��Jz1-{n[2�_\Ɣ�B�(jT����Fܻ:�Ix����wH�����H�b��ڤ&Y���ת���9�j����%.!���aȂTi�MC�J�/*��1qlG@$��Q���y���(+�J�s0�V:�k%�+U&-�9����Y�if�R�1�h<�v�&]�0�lc
�Y賾��>�յ�M�X?��H��K$VF�,,7E��[t�n8%>h^�X;�v�T9�Ȝ2��cFRtUv���-���nէ��h�,���-�+�M\���չ���t��!��L֢མ����vs���/
�E�M�-c�q"_^,oK�GY �z�ke�[�4ZQ��XU�PS�+���*����bi�����C1&���;l*m@$*@a�[�#pE3	)^,��f�07�U���{33M��I�j7P�������`ܱj�հ��dmM(]7H���{�2�b���ɶnd�]�c�����"�*B��-ܔ#٥�O%E�.br��Yx�f�&[�l��gQt��dcБ���ڂ�c�u�.V��ӳ��%�x��%�ȭSsV��3W�P����kr��a�f�ŏk/�2�ڼ��J"�X�m�ɪ��w5^֭��2PSv�"�d=������Zڑ,�J��p�t$���(�nV��A$k���i�
�Q�I�M�M�	`�ifn(Y�A�f����~�ۻv�J��ɢ�8��2�X֩b��7v��&7d��&S�wT�/7
I�H�/u���%�+�p��,*�TZ��Sl���!h'�z�^�9��`��={ ��em`��sb{���< ��
{��N���٤�%�ѭ���R�s"6��lը[���C�zq��^&/ׅ�֬7B;.dV�CrV&�`Z��ׂ��v$wW2�:�E�D�/)������$��&�6��Gh�I�8�%[e�����Zs,���L�HN<v���٣\���(l� �ܫ��w�Skh�t�˧S���#��LԼYz�I3SJ�����k�:\.&���{�Q��U���Sm}��
�K�;s�{-Z��f��%�(ֽ�����
�r�R�WE%6ѫ!Ym�!��V&��yD�u��q;y@@��m�����+T�٫����tm�c6S�jm������(�ⷮ�cN���YWv���W�=6Q��X���:%e �	u����1��%<���5�{#���"d�)�7B�]�n&�YM`7����(����k
`�Ǯ�M��	U\�N8f��w@��.LI\��zQ�2���[��W/�&��۪�)Q:�y>i��G��U�RB�����=��n���i7����E5��8
$��h��h$���5S�:61I"t�X����m\̗l�]�'38�RzˡAj8�)�j��i��b�w��:a�ŀ˩ZPJ[�RA��:�6'ɦZ3U��bT�5ω9xT6�JSŠ�ׇT��e�b��u�F�#IU���Yh`%�,C�Κ$[d��豅�B��]IP���r���!Ӣ���Z&ʕ�s)ޜR�LE*u���X�f;f�f:�u��45�u�Ǭ
�I�m�n�l=�Nk�����B�m�oR�
�ٵ1룔�E�DVR3"\�,�uor��_(������,Bl��##܎��&�۰.��]D.@e�I�Oc̭�gq�j�����j	b�nS6�j�t�[�;i�E�f�LHA�Rѥ_�DĻ͉֙�����Q�i��l&]L�6�(�/Xe+�[Ȣ{�f���c%�D�N�N'x�#4$�Hw��ߠ��\�ӈK�U۫1�Y.V3P����F[�-���^�q��+�f��a�ͧw9���|�چ*��5!������"]Dp˲��Ш��ui�A�P0�ܶä��K�uu)��B
�,QQ�W.��Y�V�x���&V=�anՑq�h=ZpMj���
C�GJ��2Ri)ub�4�l+����e8��%Z����fJ��m&�WFJ<Yw�x���6�+��լV�u��j<ÚK�P:s1Ըu�@e3*��eRR�+ ��?^ۑ���;����r�:]��r����� ��FR�9O7S�)��d%����ϙb�[�T�n�XΚ�t���)�M:�,��IZ�����	�R����UA2�df�]i6̤+1Ӛ΍�V�h� ��h�i��c 7V&F�}g����n&�i����$6�7OV��j�����ػF�κ��ؔ��T����)5`���F['ᙥ�#U�.TԳ�;���]�t*6LQ�G/GjSU ��`B��v ����m�����X�	�,�DM���(�Ov5y��������n�K�yW��Rké�Ub�����I��5����b�"�_[p��eM7l�K��H6��r�I�M"(,uxb{��+9�JLè��y�s,<{�ͽ�,V�
Pb���b�.]������sWЉl��y*3$ �{��N�Ɛ���7�:�n'u���>� Y�v04�T��j� �.�2�*ѫsI��x���pkN*܋v<a�U.��L�e-/�(A�Z�uLf]��de�B��s� ɫ�eٖ�厵u�UYbV��ˎ�D$���u���_uH9��U���j���B�ٹ��q� {%�"����YD�G��D���,�o%_=����`y����0�<%6��R=S^����������o���!W���Z�D�0��i'�:��:
;���mj�)$r����I+�IX����� V��n�����}���=��a�'5���I%��A�3�S<�fFz��2�+%uc�N���+no��}��[���VS�%&�r]��0�c�:�.�R���Ar�C6�,<u�)�����h�'���ʠ��5z�1��X˹mY�Y�;�퉵xz���7�wTS�s�e�]����9[gh���XV�q�*��k����8K�[�V�W'wːn9�¥Y;#�����}o-�
2P�o>!��j[���Zqf����>.�;�gl
���t[�������R�]��S�ӝ�ڤ�(��|�U静}
nfBY�|B��PUǵ�7}YI�=77�]j���pF�X$�S0<�G�p7�u��7�W�M�;}0YLgF��cL�Sy��H[v����WUlSQ��ٴ���kz����}�f�eF�� ��&(�!ܭ""�%�?Y�f�؞�u���k38�s������s2�.�()]��80u��8`��b�poM��y�W�*t�.�\Ei	�2u�KҠ��n��K����8Q����H�9ɓ�(�����7�Y�Mmu_D��f��(��o>�*ص����NH�&�ep�.��XTvM���� �t>��@_=�"��l����㵫�%cS�N3�@�����H�� 9.=H�C��:Ve=5�8��	C^[� :fQ}_u�`�� R�_b��w�A��k�a��ܮ�H�mGO�z���-r'�ظ���#�e�vE��
����w|������9��M��*�(%iK�@��<t�f��
F�浰��5�*T�]�hl�%0�sWB72�I����h���heo9-��N�C��6�]`�>�ջ���3+������k�vGUm3g�7�EX�1�l<p`40�4*�i�����M�{��I�STkn�Q�P���s�y�t�DtŠE��ѧ���z�$��+U�sk�'��,�bWC�A|��q"����Wne�S+:��Sc�Qu�[V�r�f���n8y��Kn�E��>���-��ӻ�{;�����r�5/2�i&�Io�Ú~#a�k^m�z��t��t��&��L��FW1�C�YC]\j�A�,w:T��T���3]���(��Pm�>x�p緙�=�H΢��r0�<����٧H-�		rRyw��$����)�S,囹)7����� ���.��MY��6��4rM!�k�W%�]n�y���Qw��!�A�X��{4+�ӶVV�[]B'])-�o$N�rvXABƍUn3��x����u���!e�U�T�i��v���Ħ�/^>�B�5a�W%J�õki��-Y��:�VE[�f��[���&�b��}�K ��+������z`J�j�M��3�L��Xqb�l�j��8̗Yo�i*�W�c����|��He��
��s�if-8®�nှ9%�w�j�G�湜�)ѡ�#�Z����_@_���m����iֵ��d���mp�y�L,�K�]1*�]ICl%�ZV�Y�%Β>È���mWɺ�5l�1ǭ>�VgV�n�}ǲ�q�Vj��뾨�+&G�E����EI����*�AP���حTrӅU�ޭR57#�'�ͣ����1�����U�Z�ͽ=e��d�ݴJt0C��fjRڏufXr�T�g^PM"ZE4��V#�z:Y8e�Jt�b��ȳ��()L�S�ξ�n�e��n�+=����o�-@��r���l�;̴zIc�F�z�9���5 ���b�����,+U|Mt׽�vI�rՉ���)n��.�Su�u�����p�����sPI��GP���X��}܃�ɍ0oG�y��(�����/fV����T4�=��e�1Tŋv��ݮ��uI�Uj��'s��1�2�n^m�9^h�\N� ��F�]ٌ�\�τ"��:�uO.гDY�2^L�h�x�)�U��A��aT`���ZۙP����K�`��<����o;�;��m	�R}t�Мڝ�enI}U8��D�w�u�Yb���]-1guv+=Kz�u�`�+�E�1�x�gj�{Zm��4̼7�]$���u%��4̎���'q1W��Y��#r4�%�p�F༓�2�E+���+9Iq:�H4���������{{34鸳k�u�A�2��zR�lQ�O%M�8�T9J����[�
֩�-rw�DbkM׷�1�v��/^<pe�cZK�v_r�ڸ�k���@!�3ld|��T;\2,��p�	��c�Y�Xڶi��\��̬v�nCbY.�<�+Y�����tv�hZ��ᙦi�vXr��S���eu�r�r�wY6+{j���'\y�'ݎuN���u��mS�A��U#T�aog;�5�y3O:��h�]��㴓�_ۦ�*A��z	L��q�"B͋�����ޒ��𫄊�˺v��t�U|4�qή��h"��2�h2�1▐��5J�Sȅ�N���H����6ȕ{"F��6�Mepz��%F�s'&3����.m�F��H�͐�R;�kd���sYj<=,��B{�>K{)�W]�w8�u� �NY׊���ǫ�M}��յk�9��v�5H��ʙvzV�ʆ����qō��2�`&Ś�{GI|o7�Qv5��'�O���f�3,��}}X�k��fP|�R�,��ܝ6��:��e��xN�GdIӜ��b��O�c��Ħ��@��.Ω��.�wAy����+�=YB̩F����} 5��H��n�i��e0�vd7���LP�k&^�����]O����A�e@�:��jɽV�ed7]]�cseӆQN�#��9*��8��.��z�g,+n�:�pq�U�{Yqv��K�/��V-�kE�;���G!��详�:��R�ك���s#j6�B����D�^�i*œB�ʀ@����񥴹���)�U���8,;� ��Z��'�1� ��`��;Q�lk���5��������.��v"��V�-�n��b��۹o"��k]v��+_%߸��;�v�Az4�dg+��Β#"#�ҡ���;m6�Õt���R51Y�\5�>Ğ�:��i��ݒA����S� Zc}z�n��
�{�N[��� K�I��w}z'�p_f�אnQ��]��t;Պ������l����/Kw�/~L�����0����{$�՛��s:�5�^�%j����'d�c���X[�G�w[7�\Ҁ�a�2�y-��5��2n�\5֊�t��{�����*��<����!��G�#���� �+5��I��=Y��v��*�?U��Z �:�;vX4�SŔ��%��v?�:3��ַ�1�!�u�n�ښ	[9��{p6��lԈ��Z��t#�G��)��u�S�ҺU�ݙ�+xKGq���9	�k��z�MnGJj�`[pml�oy�i�)��^TZ�H�N�_\�7$�o���WZ�w������PL`����
��C�֭�C���lUi�ƴC7���3��߅���dJ�j7��3I�R��8���d���΄%�f7C��ht=����y���`�&HEv^�ƻX�����������kyX��xW�hhX7�
���ْ|J�$d�ƈ�ǔ�6���#(�|� �L]�Y�)��Gt*sܗ������;�b0�kS���o:�I���Vʱ�+2Q�A���s�j�ń���� ��5��� �S�=��7E���Nެډ`/�p2Z�����R��λ.�iۑb����8��,C�7�xT<2��c:���%V �j#�uZD&mQC��n��uֱMs��㚞v��'��nnR{�[�j":���w2�|û������c��p���q�y;Y,>@�tv�����F��BN�j�Eܙ�[0
�����c,�:^�'��Ź:�H����xQ<��кJ��֫�[�
�,�Q,X]�]�;�V���oY��^��Щ��:3����ӎ�W*l^����Ø�퍅��J�ЭYP�U�oj�r9�}|����[���^pEq�ҋ#����y�-:Mػ�f���^���(�Qҽ�mK�K2V���i�ל�>�9V쁗�2��d����'!�Z2!Mw�����`���H�8�;�#$S�˞���twנ��'_`�Q�`*D�C�:��\t�Ӵ�k��[���9Q-[�e����b���ɽ�N��ӭrՙr�R����E�������Y0�oY�>݈���N��k/iS��VU�	�޹]�ŌB��t�n��w]�&��2�^9�^�	;�2��3u�V#;���h͜��.����S)`�t6k�U�td�;*rԱPdFt���"�ut����SW6nt��/VD-��[�h�T���1ݯ���&ç�؝���wuk2�jH�v��ƥ�������F���YytWb����Q˼�_.�@�M���Lx��-;�;�h۹tI���u٥�wY�b
2;ʻ�U�A�A�\�7�[b��.Y����i;���|��=��b\�}���B�C�:P�Mg_D��ь��oǓ�}0|�H̜��W(fA�x���$t��[�;H��W�r�M��԰�˔��k�U9�ZE��Ñ��5�WS���bڧwJ�
nfd�J�)l0c��9w];�r7\㙣�gd�A���Qum��Db��j-�5�Dou���.�9���N�̸����)j��`[.����j�8뮭��u��t�S=��e�mv3� >��|z2��$�Π:�yt��H��r[�-y�~нe�P[�C�+��xg_1��]λ͝f��\�b̲��S3GSws�p�c�+7�G�j���{8HBz���s��|��;>[g��C-��5�ڙ�:�E��ޜ*�S����W�,E2�����6�7�)Et�����w{��٫�k�������xq�x����aA۽��#�yMb�u���Ņ��<�s�ȇn1+ }7V[�9%��e"�Yw��r��^7�Eۍq�M�f۱��G�Wײ �>z{�(�|�5�+�ax�� �{jl���5��v}e��W���wI����"R����r1�+��W3^�I�XPmI�w>��d&�Sٛ�NG�϶p!k�� L�K��k)-�7���y�&�f�s���I�)i:�f�m�gn�#��Zjo1�(�]曀c�*!�jh��3
(lXuka��-*ݪl�ͮ��`��t0���bc.�b`��됺0��o��f�(a�K_H�h.�%�b��������P<7k$�/~�O"�L�ǩn��a��ۅkdv�(���	��Q��,���R�G@]����[T��+� �#�������_������������Hu�&u���$  ��쇧�=���C��3�|���9�����_����ϳ;�<�	��أ��y-�c۬�qbV�� �5\4�:\�ḛ¡Ҫ]��Ћ�m�'(ȃ�����=sK��\�Ι����<B�F@�e�YD:���g�aU1q���iR��\��VU�eݮ��7��V�
�n���6޹B촓Uڎb�*���Hx�>ϸA��:�ޫ�E1��ʃ�[ϐ�naݲi�����N�n�f��kl�(in�d��X���Q����3r�EE#�e���u�Nd-,nv9f�̕�)<L7j+ck�s�S-��b�t-�h0�T�UH�V
���s�`��Zۚ����嵖��Ș�Q�]��ّ=���_
Ym�<�E��d�b����:[�;�R-7�́+5=����2v�U�y˰��K��L=��D<U���Xݢ�V�WGt��+.M��p�<�#�����7{�pW�V�4��Erkk�[�r�N�Ad}F�5#������B`�DJ�4��J+�Wē���O��!w�Q�c%n��x:9�r��-��}q�����l��h����Yy�a9�h!��ך�5��4��ˀV��0���!Z�";����f#*'�z7�vԻ�yjR� 
]����h��%T1�ߏa٢�qu�-��t��n���2]<�9��l�v�F[������w�͌���������V��|���Ũ+ �Yg�Ҽ��D@]Z���Rn��(ؙµ���)AD_a�+V]��e�9��*4��k��p�h���:�[z��ɫ�- �`�T�he�}�k�,�ۅ9�j*�oG���]��Z���ʵ	M�LkB=J�kw��y#�:�D��e�WW[�G ����)X�B��d�@�iK��N������ؤ�W��ʻ���b�H�e=�N�������]7rEٵ�NKĪ;��Մ�a��l	�2f�GWd����s+A��2ť\�1�8IûMY�[4���Kѵ�[)��K.�1%�w56�^����4�C������g��%�^$4J]������c`��*��8���2}w�:u��V��ޓ��YeP�{��%pe���6��/\�ݘ- ��Ζ�7�[��%ZR�x���?+T9b]�������펏d+�>��p���P��iX���`���� \�j�vG��3��[4�+H48;/s{/h�����UoO�\۵�s8��W�D R�HoRb�G�(�6�N587�����V�r4�b��i�����J5o]%�&���w�2K�M��/���X���4[��I�_F� �op�;g���ǯ�����Pj$5�6���Ml�5׭�Ǡb(V�,��=���u��4��c���Ćn4p;�*#���.S`=��^���%݋��hYX�J�e��I�\�������؞VT��|��to6�\�6���ԥޅJn��(��֪p��\�<�� �W\�4B�*���GL�.d�&1yBR��� �h�5�i���=��3�H%�3`�坫�|�:êE��o�ۥ��֢3��
YՏ���Zp��$ʐgæ�e����,�Ö�U�jNs8*��IM�TÔ�δk���t}ұ��>�]�ow�j%���+��D�T�v�Z���e�Mn⹩!���yR�Z)�HV8g1Y6vL�Yce�ќw��'[:�jh���w5��jvg;�2\�`�(��A����ٵ�t9�
��V��Vk����*�> ���H��I�X}�/Y�]s��Cw^5�7�)G�z�q�B�m�e���$oD�� �)3o�;c8�ۙ� �U;Rv��TݎQ��.��͛Њ[X�Z��g��Ea}Χ��Cb��Ϡ�;7�D+��̬�n��v�����L�Nt��}�|�V�F�n&�e�n��Y��j��&]뮮�T�\���W]Zk�d�Ûf&etZ͕Б�9g���<��W:ђ�ۤ��K������Y����`����X{MF�5��"9̧y��f�ݱ	��خ�|��-�.Dk>�cK�-=�|�w�ku�K&Ӣ�5��M�R��[;71ε�ǧ9sQx��1;�J�:��s{7lJ�wtt� s�pU}�Huۛ�l|÷A�R鋲�2*Ԥ����m@��7��EBh��[[��W�`E!MRf����Q{8o{j�P�-:�X�ǳ��-��q\��[�K�p
���\R":�6���4��MnÓ��λ[wq��WVq�8���q��9GOv�OT�A��WJ|�m�,<�`��m�ǌ>����ꬾ�$(�(�].�*���1�z-0)����͔��O��q*+������e��.[ v��x�b�m��Z�g-��l���X ܮ[WRM[�;8�tn��w �tK�g�]X�/i�*��!�+M�k���jkS�;��m٧���.fٱ���gs���U:�ڳ�R��I��h�;�>�R�7�5�r^R�	*��7!UxpT4�*�Z���wu)�]M�A�;��>Mr��*���y\#poF�v�߳���:�W�����[֬|�U���p�QDs*>�k,�ܰ�.S��p���9|
�:f���x��#�]��@�|NG�V����gf���E6l����8�e٫i����v���rZ^=��+§`�#�V{T�'�����a�� nU�.-�d�5Y%g2d]�}N�ő�ĝu��('&I��ᙋk�Y����z�+����G,��.K�J#%��cޜB�osWm�3M�	G2�jϣ*�/��M��Ȋp�f��ʻ]�ݱu��w�$��R��kȷ�8԰U��p"@Z��ۻ���gH)�R��Ӳ��j��])�9g�2�w���Y�C��捃:��|��g��ՙ1vm5y����A#���Q;��l�ϐ��&�_��N4{���Ὗ`�ݒS�m-��AQ͎�
մ�Lr�q��ս�m��r/���l�A�P�%u�3��-�k-7n����s�օͭ��ά}��s��R@�s�k؝��l۱y��^��vY&��]�ŝ=W <F���mY���8�#ҠxD��f&Lu������`@$�fS��l�+/e�M ��dQ���u��A9�T�<��NS�l����Qi�ekT��P;���W2qoe�����X�K�l�����`u��Q��Md.
|�#9���Jc�Y�Uѣ�E���{�[�v�G�|�!�b��ǥF5w��Y�}�44'fwd��']2̴��ϵ��e�T�5h���e�ø��$/dN�k�
(.������e���yA�����w�@/G:�},J7�$�2.�+5��b�js�{��k2v��&�nQ˻��t;/�;)M����Ա�-m�H��K��#����E���t�L7�}/+�-�*U��Th���Wu��Qx�)&Ɋ�μ��R�m�_P�2
�D��{���x���F)m]༣I��s�RL7H�em�A9a��ñ㾚�,���<�r�xq�#6���D��Vv�@T�F��.���E��%sj����-#ev[
��F'WL����F�;f��e�QT�qa/,:Ы�S(�k	P�"U�+L��w�]/������י	�S��<�)�z�K�/_b��scz֎���k�A��=5��1�h3�ѫ̎�����-�q�WE�-�	��Of��R{�_�ݽ�؄��g0���v�.�Y:��3�C3�d@ۗ�7:��/;�a���Bu�)8i�o*���9���P���������z�=cvFO[PO��	[�=jm ��N�LGp&�k2�6��������n���}��;�����ug3A�qDd]ZN
����|������y�*�e5z������3�y���.�ӈ�Նc��c෩^sX���}��o��t���,��/B̢��p�sI�"ۜ�+j�ֻ��A��޻S�Z���f����N��@j�j��1���[O`x�&L��Ŗ��������:fwΦN�a�3���O�,:���]O$J�qp���t���Y�
�,���9`U��(h�ݫ��N�XR�>�Xe�y��Yi�_l7�y^J��eq�N ��8�|��ӀF)V)[��]�E؉��镚�'g\e]�)��{Kr��E��^�r^U�A�B7IM�Ӵ�o�S��e� �R
�������V�qc��!�hL�s3{'e&���b�Kv�J�dQCk�#j��z���ϳ�`w�5�Ի*T��AV����a<�����w��;U&P��J���{Mv��|Jxvv�sf��,��s�:�sq=�,�b��9h9\#�U��`�$r���Y�t�S����.�+M+�x�븑9�E���r�.�&P�X���q�m�MM1y���L!AZN�Vj�Za�z�fg!(���'k72�)���U��wEܜ��GN/�0��[kj8l�[C�]�Z�T�x�U��u�ڋU=���a�����}��d/xn<u��vU���q�3��@�|�j8L�sWMN�Fr3��{�
G�A�z�y��ښBt���o��gt��:�u`.�'b�V���x���q�ڞݧ6��*��l�WA�C�ˮ컮-s+a����ig9�	�_��W�����B���w�[������+J�j��[�iՊv9�˽D���e��w%�gu���e��eAd�]j�Qt/e�����Z�#�
��+(��lZ�htT~�Z���p�V!�3�8r�EVO1nc�IT��M˂�]qA-�����\ZY���wyo���]���0�'�]o$M؅b_u�4p�49T��C_6��v����l����L�g�3\��qZ ΦWW\�5�s:��'e�ü��n�Gs��ٜ��q���O���ɤ� �;�>t�p�Q�Y�(�V�e^}]��"�pf�1�f��ֽ�W;}ُ�����i�����-d���V�	�Ц�hR���DԞ5�7v�ȝ��9R�[�~��\9����2�����u�<��/��s��������yX�8�R#�n�viq�m�o>S	��&uД�\rf"���Ք�\��%�+���T/�E�v+�3mK�{��D��	����*T49�"{(W2i�|�l��2�*o�hc8�,v7^D;F.�S:�ȂG����J�ݺ���W�[�����[CE�R]��d]4r\�(�&�G�����Fr+C2�dŸ˨�Y�b���h'6�'`9�E�]���NX�vm��jzۣ�X�T.��t�s;��SU#ʸ���卭���`(�"�B�Ypwt�:��b���ʕy�.p�"�I��[f]\�R̆�mfst�bG�ac��t��N�[I�xG�"׶-�3�6�/znTBRsc��Z�������:�9s�'$�ą��)*��kֺ�=�]{sZ��BI`���d���\�\���|�ߌ���޺������u��`���HA��[��qв��7@�α.4Zw]<�7��2R'�@���v2Աy����l|e��z�\V�����u7C��&-]Ӷ��]�w",���5zѮ���;[��%�V+�UrK����iMβ��2>_q��[)pȯ�o-�'¶n9�!��b�#��]�J�*���;�Vn���r�m
LW`�%��Vfٔb�b�HJ'_ip��fu��e����;��I���γܣ�:|����r�'�.9��g)z�\�!鬱6��$I��gq��+�wV��X�*�ٷZ��{�V����"��v��Y�VK�SR��msU�J�E[A��K^��l�v�%F�ᢧ5�B�P+�.p�� �J��vm��}D�L��B��,Kˍ�|y��3�A%�7s�Z��]]3{������ordr�W�ڕ�̺Wt�ì�Nv:(Vk�COW(e�;O>��.�\4w֋z�S̫HX���2�7Rf�r�5ukz���6G�z�K6�7YT�]��5�o��Ӽ����{��ɫ�˦l.���p�Q\\V^�Gx����8�=�:�ZYZ��פ���2��L��nuw�"��>ȱU~aX��ܵ�T�[h�҉�R���AL�C�Vڢ��K���H*�8�PP��TR�`�U-eL\����TUG���j2�T�hקj+�C31+(�lr[Z�+k\�Q�+A��Q(ьI�DƊV���R��*��%Vڌ2ڎY�EUm�:�F
t!\�Re�"$X�,*�[aR2ژ�+p�ʖ�8c+m5Q�-F*��UV"*!m�TE�b6ؤP����YV�ŀ��-Ia����U)��F�5���(*(�l��b�h�E��0*�QEU�6���Q�h�X�����_ވjo_��LWK��ݲ\����p�' P�6��n����W7{���5sE;�ۥS���+�����'�/�Zճ�����}�]K��v���#X^_���۝pk�V����eǇ>����`�ف��u�D�W>�=��~o��+�����]5���]N��4�b��Y�]} �Y��C�!z�G�z3_R���i���d�<0W��=�+K�oph��1���G�y/\�]�뎉�	S�)�_p^g��"d�)��#�vΚ�sF�{5��u���2i�P�G�<j���G�Ċ�{d�O���k6$e>�W8����PZ��m����K�����)\w1��urG�קbz���I��)��㬀�_M���y�C�L���Z?���}�~����M#�AYA`LҒë�za�J�t�ټӉ����{[�`Ű*F���X�8诳~%l��
�o��֤3-��;��-i�Y�����v������h�r�N[�K�9���:�#س;R�:���9XMWU��ϏL�L�����~[��hU���8m���z[�'_��������i�Y��}��r�X�eW�*es7<��A鸕?vu�Oz�y��]����/X���+V)�y/N���bG�S;)s��>[LE�Qp�S�~��zN����a�����h}�~��y�7�N�w��]E�{���}�u��u�r�g�ơ�;��m2*뽸[+7:t��7<`�D`r���6FL|3��}�gXX����E��t\*0��hV�N�����}��z��M�1��>�\w2W�8U0�г���q}_7.�N����w��J�==5cn�VͰ/%tY���wLNRO/{J�Y�o�ꏺ�(7y�ֶ��w-VX�y��lخ��6�	��3kpJc����':wNl��*��O�Ng �(U����,����'Vt�R���d��C3������54��m���x$VAȶ�fQ�#�3B�LM^c���X��׻�t�����c�C�*q!;��;/:�Oq�=Ό��]�u�Q��m���q�Ϗ���Ǿ�;\�A����@�GݗNdc=��*����y���X�����['�h+�ĳ�2OCټ�,R��I�=�џd�:_\��yWH^E�ʋ@}�}�=.ڼ������5��hvE3�ws�w�8]}��<*f�`�����]��<۟7Wk}.�v{zG�#�&}����^V*�ep��1���=u�^���.�7Z���v�=�f|�W�<�/���?;v�c7�kkޱC��t��ܖ��U�Ŝ�J-����ij�[]b���^0����nŹˣ��^�(S��4Z����۫G�#/1_D��gBډ�:ƶ>�ý�c<i}>���߀ӊ��qi�V:Ǎ�+V�Iў���]Ddl��p�����݃C���X{w�?�y
ƪOS����W�����񝩕���y�\]ֳP��ȶ7[��s*�C��ƇS�<*��v��xw������0UF1���qt^t�nhkyid��v�@:�z��n`+iҏ��';�Ѯ�����*�F^�d�xgk4�mN�N�{y�A2�y���bj�i�2�q-�c����wI�N��6��&����]4���s�<��o3��^T��S{d�~}=^L���x����?aBvKc�ɷ�î�m�K��A�g�yAU�]Wiv�7�>��T5�rt���d�݇�ҡ�w�Z���^�*�����Kkc����P���Ӱ�;�:����p��EHsNJ�eE�6��;��ώ������w�#�I�,�6z8��|���2q�b����͝��s�|�x_J쭊ࠜ;y�r)������]U�*�󑵋�L_��K�(/L���/\��=��X�8K=7�'���m�3���
=����qu�S��9�z����d�Œ�g��ޑ��!G`�`߭�k�WN���O;�˿/�~_iX��}������Ï�����v���k��>���Ŋ��||�>�J�&@gM��r}SҸ:iah^ྦྷ��:	fmMݝfuǝ�7�����S@p�U�"���v����U<g'.��}6S"��|Jo��*�W�O�AS��9����<%g�lԑ��c%g�uཱིIٟC\X8ۮ�M#�n[��=��^t���i�Y�����r*M�5}�zrSX4�V�}ʢ׶\+@�G��������}[�r,]�6��j�>owB��̜z��X}8c��s��3���[����*{seΑ�5�.�+� {������ހ�75s5�����O�]��oQ�o��m�־���ے�J����ڝg�Yҋ��}Ԯ���J,J���~��۞�y��4�[D�#w��A�x+3ebBM�Ÿo��~ޛ�ޯy<�6�!{Y>�==�T�3Bľ9�N��:�wm�~�k�e����:i[��x���Ծr���e/<�ұv\.ָo=�>�禷����<(�`�>�۰g.�uH<s��5.���.v�r��߫���'�gL7�#���,C���m����lƳ��m7�AU�d ~�ku �ݻ��{�IW�q���Y ��Q�=Tz)f����Pf�t��"l�l�o�.�̈́����6�a����{�
�{I�8EԬ;��8�F�n���9W|�.��U�S���M]�e�fQs����qv$�>�J�����{���&ߺ����^��={�u�y^2�!b�V��;��&D�{(VY#�K�ri�~����/��m��~���}��TnJ�A�:�\(6���
�MgB7eI�s��/l\��x62t�ۆ���8���t����-�뼗X�(��>��*^1����B1Q�Ȫ��e>~v���TFr�=N�n���|e�����G6�+��wJvy�>�i�;��uҏO��q�EQT6q;�l�)�̷j}����r/�؅˖��c������=i�I���l�ɠ���V^|���!'�F���v�bJ�x�_�\�}�ʋY6�ҋ��\��r��L!�ں}�N%Ӵ�Ϟ�ิ%"!��H�֧�7w��٪AN�q��[Q�p5yWWi�����^��Ϋ��ٙˌ���%$��zU�.:�.���O|�}��I�!��u�+*���[�ӗ�C���żv��Ηoݼ����O�_�=��!')�z�q	:�_[�1��g����5�o��O��*b���/ޗ�:J���P3��4=nm��R�A�=��'y�{�by-�}��B���p��C���*Ǟx]�S}������ō����r!?2�p񿫳l
�e��w�����y4�귇��Ϩ?�
��Rt�yC32��hش��r��V2!�O���������s&������^���B�����ۉ��Q�c��r�c��{���Ǐ��;aB��pV�s]��C���+9����+�@�B���ʸ�V�(iʊ�~	Elp�i�zC?20�J���^��b�]%g�=귷��Jo)�f%�z�.{���9�50� ��V��f6���r����Л�z���k�:qZ�n><�8�������,v�J��9m���ՂU��{�~9�w�/�ą�'���N&�����<�X��x��5������n\��,�z�]��G��Ǔ�Θ66���������>y4;��_��d�~o�>��/�d����uU ��/����6�A7�s�󳒱VoGw���_�PK��At7�حj�Eþ�5���9.o�*n_{�]�M�V��_z�a�p:��+|P�}ʟ�����y<�޼�W�<|�Cdv)Q�}�3�^B�l�M�7}k�|�fEo��سv|)?�:tF�o�~-j��q���.�s�^�,����.<9^�.�|�mԗ���C�.^�����]8�=L�ǩ�ٹ��5k!�@�0�?s�`�%!]ZU<Uze��z�/��l��Ćm9	��.�7��z��v���l���ݮB��d8s�}9�Z�ɭ��It��O�ʏ�k��Y�U�7�Vԙ~�����"jU��~�h�����˛�}�zS�z�mO/(!z��G⫝�%A�q�;}!�f�W�l�)�3�g�^ͧ��٩v��P���y�{-��;EN�{�����Pe��HP^��-�,^p�{�
����#�F1���J�=5�����<^粝����+��h�<�	����8��@�\=��m�{j;�Y�ɶ�5�Ю㹍tT��x�W89�d��^q�|���t��J;J�{�֩�}�<��L�h@�����S�B'��V%&��,p����ڇe�=齮ٟ/<��睕c��-eX9�>���>?�����1���~�p�����B�ewK	A�YgGQ�G:����T��-��]g*sY��Xl �ّ��es���R��Ey[�nj���TF��^t��k�#�M���
E��7�K��L���B��'wJr�Y�S��ȃ���D�e݌}V�b�.�����Z���Z�R�ud��Wذ��#["<��Usʼ�{���P��6��F��>����)̬����t&�n�;Vޮ����z�
���y장:��9]���Gk�*Ug~�y:���wr��H"(���R�2�]Ğ�G�k�6�l�ͨ;�͍�i�J��z�ogV�������f����$�(򘥚�
�E�E
Yq��Y%�/sif�o�=L�ݎE>�.�U����J���u{η�v��� �`	�/Xˈ�+b�sO6��1��W4it,<��Y3e��ǃ�����Kdg!�+�#*���3v|\�Q�)u�����luY�٨WT
�.X"�� �LƮ��k]1Ԯ��u4��ܮ �i��!�/;P�B��ᐍm��%��Ifk�?����?r�f�! ��Z�enf�%hM��.=��C�*�'0�D{zU�y)V�u�������̠��TU��W�H`���9^���A]��R�j�D姭j�DZ������� �J�h��Y"ʩ�5zM���&�5ʺ����v�r����w��E7yf��mEy)ȍṘ���Lo-"�2����H��I�nI��.�O梺x��D����(ڵ4^���Դ��3F��7����q��	,Ǡ�T@�w@6u�v�f�к5e�M7����g ̳Z23�ab��I�lw+f_-���{ZH�e5oZn����%oR]g�k�K�7cB+`@qVZ�!
f
�,f�0rYXe��-�>�r��`,�ٳ�5��r�X�ƪ����S��s9�%w$��"ĺr�],P������X����8�@�]G�+�ve̟d�p!kQ�Zg���N :`����]�`@B�2�u�ga����a�wR.�[�۵j�Z16�k��k#:c���K�`43D��u�!f�����c�$ҙ�rsy;wv"VQ~�OϽ�M��+}�Ul�N�9"ih��W��f�s3��0�'ܩ٬��ߝ���?�����%��KmjETZ�Z��>��c�bح�`V.%E���T*6�-�4q��j& ��X���6�s0�Ȉ̭,b1T��,jW��G+j�k-�mQF\����ETDW-�ŉ����EUDR1��U�E��Z�R.e��+Aq�m-,T˘�U�L�c��2�n!�ڕ��U�m�fZcV�Z�Ube*aJ[F�(�K-���+S��l���Z5,�kF�Tm��%PkU-Z �F\�Q�iiB�n5L���5ƪ�R���Q1,�F4�[KD�*Y[iU��*�"�-m��q�r�ťˉ�,�Q���r��\�"���[KYH��b��cD���F�J��qQb8��%�U�m�S332��)������aU�Q���s\�]���_Q�].dWܮ�ԱS�5��"��r>u���x��+���y��{����_Mˌ��y[,]��3���k)�].�v�7�)_c��|��Rg��M盵$�*�:tT�d�X�̫��/{�-򍑹�������h���7?$��ٙ���_G���V�;��_�o�~��I���ѡ����#���Ի�P9�9�� j�7����U��ܺ�4���s-�q�1���=�6CyyM����m��q�]��{]>������cx�a�����/P��Ɗ����/��|�z9U����B�
l'�����6Nխ绶��<��a3��̔䢘�г�*�|z�\}�����ύY^t9�0V�yè��K������L�ov��s}��:*	���n.��;\�_y��_
�-�~��]���>����&[����Ҝ��c�,n}���<X�M��/*��OM����>[��U�Nfk鈾��Dɯ�w�rWݎ���>�]IĹ�o��ֲ1�B�ň���g���9W^��}�֬=5�]��L��U��CϩiRq2\��~�dz�✔w�['����9V3/ڤ�ū�쾝Cy�S���w�ٹ�V]��WEy��=M�j^=����w�OݕӮ���ڤ�z�|!U��,�%�H&��pz�U�\	÷;��2xw{���;�jF�^��k�^�H�OP���=��/;��7Qs\��-�����/k����)��r�.~����MŻ����|sWl�
����C^<�p���>U]sӦ[��Vs����"��Ww�j�ً9Su�W�!��z�\�b^n�y	2��6f�A|wz_t�����Ys�U��:ѳ���(	�`����VcԳ�t��B�.6�M3t�`�-7k�����K$��>*����e��s�Y��n���<�{4U��u	���:��]�R�ѓ׺�{�ʓ���1&��!c9��+��-���.�<+U�f�s��8*m׋��^��!<�s6Uٺ3�58�����e�bxV�W�q:�;�ᵓ��3~�95�p{��*2c�;��W��jV{�qɯ�'��=��l�I�_K��F1t:񙦶��)N���N�>�R���LhsI˖~x�I�A�{3�]a��J����ڄ=��)�_������5Y����ō�5�^5�>]�uU�z�1�u���ז���v);��f۸yOUe<��;���(d���j�튧�^uۧN��ϓ�֛!���4�&,G(.�OmA G�͇{s��|�.W$�ڏ�S����O�t�2�t��}HR��se3�Ϧs5Yy�L@��o-�oz�R��)Ԗ�r>��ﳺ��<�q{���V�Y��rB�[�w}�e{ðKZ����2�h!�#�}3�8�Lf�/e�޵�s~S<�cd돦Z���u�(�Lw��>bw6��k�������;۲3�ܻ�W&��&��iЬV�����jE�ƺ<]�ң:�}�{���NT���={��{�"���D��|����O�1&�=@��3�I�靲0�;�d3�l��9��������}��&�+'��3��q&�cξ�@�:���d�a٫����2�+�N�� ,��O����h�~w�����ߞ���z���d3�+$�ui�`kT&�-����C���Y���b��~� xɞ�h���~�w����^����<��>�ePG�CԜ���gG)"�i���s�d�=5ghd�C��'�7��$�&�d���{u����ywo^�y����\�Ӷ�v�8u��l�@;���&�i��H��d��l��	�$�Y��$8���;��@�
~��&s1Q7���!����W�_�uk]oU"�AzЃ[9�]�[�^��0�j=eeg���}4<�I3fm#wum��d-�y˅�ѧ�x~i�U�"�dO;{/"�K���yܧ^k��_k�k��s�N3hN5 �'���$�]��6����"��s�ĜI�I���V��1�nÉ6��nn�z�k����������l��J|0�?n
�>I�4�(N��'��� d�2M+$��N2mOP�`r��Va�����0�/E���y��ӀQ�}����0�8�w9���G5�x�7߹!z��RC��!�'W���N�d�)&N�6��`g|���/���u����'H�ui�7�$��I�n�08�u�7ԓ�cud�y�a;Ht��1$X2i&�E�z��m��z�ܽ��=�;�k�z�;y��[��I���L��3�Y�ā�����i�V��'��X�;Ha큌�"��k�{��cs�+���wx��3�?�_}��Y�I��O�4�I��i;x�d��w�3�'̞ i�d2y�$�
í�������A}���;y��O�i$���=d�,9�L�uκ�|�ٛ�>a4��hm����@>Oa>v���ƾ��𯫇�����}��+�'��٭y��$�
�^�`��,���r�2n�:��4��u�!����&����>d��6�:g��CL'<߿o�w�����|��!R@��R|�����M�Y0�x(�N!�Y6�xZiԚjN� ���~�M0:;�	���W�?x�J�mq[�'������? c:d�p��$8����Qg��$6�P�{�d�I�����e��4�Y6��'O��$?o��o��~w�uγ!įZ�on1�
5��
^Xj�����6��h�.y���ۭ%>�w��1�B�
��%)��`��L~��֋�l�;U˷/�q�9�ͬ��YQ]��9Y��M�X���V�i���c��~�]k���hp��m��/�Cl�@�Iya��T��Xm&�1}ַ�C���m��d������8�|<�ߏ��[뾻�g7�}k�bϨO�9Agl���d2�d�!Y�P� Ұ�&�`kVCl��h��������9��o����hM���gY����5�I��I��d�J�L����0&��q!��H(cI"ɴ�}��d��&�d3Z��I��~�ۼ&�O~�k\���	�~�G���;��?$�[	�;d��0��!��N�bCi:�&2i��"�d-�!�度ϯ�W'��%�;����
?}��=��q&0���d��7��C��<g�M'a������3�d�П2VM*��;I�M��lּ�6_��s}�w��!S�V�b��i��v����6sY�����w�'��Yq��l�$���'ЀO������u���%��@��B2nӆ�'�N���T�ѪI��'f����b��I��ϰP���v���<C9���<�{�|��]k��7;��RM�����z�l�6n�8�g���n��v�	���'�I�N�j�C�C�~������^|�y��=Hm� ����$�'Ga6�>{l�dݰ:��'�I�x�i��ɪ�H@�=���I�b�o#�ϳ]��]u��x�����4���+��&�:�x,!�Z�7l��,�d���$8ô�x�|�� |��{S��
�Ϝ�~����N+�eyX^�g���{����\��h&�;��|�5�)&��݉&�+0ҝ6�w�6��W-Χ���kssEs�]��,���x 9��5��t=Drո_�=;��y�?Σ�z��}�v��[>d=��i�a�oy2O�����I��$��j��,&�^9$�L�Z���I��s�0>d�>����36���q�P;d�f��I�P�H|��a'�V� mub��P�6��N2y� m']�:I�2'�&��|�_|�{k�g�ԫc�ޞ�� gO�x����Ӈ��L�Bi�Z�4ô����,�l�ՊORL��Y�꯾$ ��%ڨg��n�"���~}��l����%~@8��03,�$�6��d�:���!��d1��0��hVN��Y7E��a=֞���y�5�i޳�p��2m��I�C�;Nˬ���O�C�CL��Y'�6�@�$�s��6�ﯲI�LE3T��D��ާ�n�=����㟓��<~��$����a��+�N��&��tw̐�!���$�s�$���$�
�2�E��m�w�����f����w��޹
�l��'�C�3�=XC����>a5lRW���P��gx�\�m!��y`)�N;d8u�+}�^�����[�E�c�ağ!:��T2e��7�!�
�����E&>$���v��|�|�+:ݒ��������i���T���,֜��}��^w�$�8ΐ��Ͱ9l�F����d�s|�HT6����'�V�M�FP�!�N�Rl7�;��u��|�����9�k�����<`vy@�'̚G�`Cl��$�m�7l����I�;9��Y*L7��!X�}�*�𣾿6�~��9�	�:u� -��E�_词[vϫ�<��R�M��e�6J]�v=N�sB%�u�ǩ�szJ��wib����Ũ &���Bl	�1�3��ֈ�xVz�u��L&$��#�guwgk��f�E;�;��}���N�뿻�Hxɤ�E����M�q;�����m�zÌ:N2sxi���=0��0���羸��}��}�?kϵ�BTOl$=B�0�O�@���4�I�(m�ć�=@�'-4�v������0�I��C�÷7�z����~n~��|G�����}���P��V��!�T�woI�N�d�)'�u�i����$��N�d4��o�~�����oZ�<��k�>La<a��CL���$�e��]�C�t}E!�C�=C�N2w2��&�;�!�[�9l���M2j�w�������7�|��=I��p�����,8�m��P<g���t�*�'̓��$=M2z�H���C�d�w̒i�����O5�I�z�o�����^𝵒s�'�;OXe�8���	�t�О����i!��ِ�0�{5I� �E��P�4��N2^x�w�s^�޽۫����O��d���XM$�OY>I����xϼ�>a3�i�Hd��~�0�����VI�=뫻�7�h}�v��s_kb��(E��Om"�����	ć{��8�m>�z���6�6�S��	�͡4��ֲO��oy}����~�;�O�T=����,��I�_�<d��;�Iĝ=\�D�`w퓌��u)���Ii��l�]u{�_y�yל�s�����6�Ę�3T&Ь����m�F�R|��<aS�N�T�`z���̒���0��B��~�����]���.��F��mWb!�&�'�M��+�gyGwŠ$���r,���:����p��b�{��kH��"0k�|��ga롛@���5}]�]9��S������˼G�LaS�e�I���O�`y�&�m&0�a�Vtr�4�cēf@�%x��V@Ys�	�!�E���G[�}y������}pu�w�^�	�t���4�
g�+$�tZd�,j��%�=9���%awE��'��a�z�o�0�M{��y=�u��{�C�IY���Hg)�RIߖ���4�)6��mX��NZ�[�R�q�-�� O¿E�D}������;�~��{�x�����!�p�	�8ɶHu���Y� y�I�'iēěL��l��S���ެ�v���6k��^��7�����Vaÿ3�a��6����g'L:�ChO=�c'Ȳu;�v�i6��(O6��9Ւc=55X�<���;6~o�ף�~���������i;zC����^Ϩ�;`f�<g�'V��8��_p6�[&��a��d�,���M2rӘ�����{����l�2i�톹a���{O
��s$�s�r(C�=a�CHy�C�:d�9̀|����m����ߝw޳�����5�_���x����H�rӾP���<x�x�{��'���RO�;�y'����R�3��$�����?�����k��������������'4����	�N�i��!�����@�`x�Y5���VN��!�I���G��5�~��"������~s�<~�O����~#��C�8_o�;���7S}Δc��]]�{	�]��7�dw��f�7�|�~Vj~X�߯*;΍�ȷ�{<'��_�M�Ǻ�����	Mk{����UoFN�]6�j��Y����ڃ�3#�͔'>�^��ё��{�������R{�w����w۪�*�m��t��һ�U}hS=o9�����wO:�ʔ~��u��[��M[&{���ؿ���5}�~���O6�{���Kz����W��T=�=�ζS�l�]k�[:tƚ��t�����v3ؓǼ���7���<���1���6��Ԍ7��:�[�~�\�z�;*����Ú� ��d���+��w���t~�v+ܾ�VvH�����+�eo�F����ooA�z��^��]_R�	���᡼u�`�^�*���&�d��f��N&;>�⦪�>����ۛ��y�D����'U_�F�옧zf��g���!s��A���5.w\;û.�r�8�ݰ�?w=�5MuܬfǓ7]i��v�GK�D��5�LV��A��KEu�l0��_s,^��K��N��`6evr�oX�U�#��!;n].H\�yj��j��Q$��ȉ�2�*Rp���1�]���D{�15d}}�b���7�R�:�n`:da�x/�/��l�V��vsuv�U}u�N�j������c��n�o5�o�F�%�l�&�Y��yս��A�����A�@�]&*��O�t�7\�ރ��Hz,_-��*�#�8�,������gV�[{=�2�pƻy^�[(�l�Vv�	zۛ�z�ё ��Ǝ��}������;>�-�m��5��=�����uG&����g�pci�O�y��\g��p�;� ư�2\[u�ov�P���}Oq���Q<��4�D�_3�V��5�R���þY�ȶ���@rKF�y�e�(���}��Dx��vdN�"=��h
�]d-і�#�K�x�����D̻�����av]���*�v���ݧ���]FН��j�������9+ƞ4��ܙֵ���E�,[]���̖�R�].�mq
�Vt����+�t|�뱙�����n�F3�"����&�>ZJ����6:l�¾:��t��D?����ʽW)D1h�aV}x��@��K�f7`�իr�p �R�P&�cbTdWko,�{��SHx��p2��-��$��*��k%ES�F�
t�bV�t�h�$�r�c��Xnì0A`�"5�lh5ڬ��[_u�u�!׸c�$)â��H�A4�M�8N���}o,A{A+8�(d92�ڳv6�vT>1��Ц.$�6�[l�(`��5r� Px�үKE+���E�s]@��W^��"?������D��:�	*���Gd�6z�������E�S`jm��v*���\�l*���+B�Y��Ѥ���F��A�Q`X�s"�C�:�ru⑊frO��#v�Z�-rh��jVs-�I]��:�9Wu��xzt]W���T���9[)\�'^Qq�+9���'gl�G�w��"�fb�=��V�%�oc���q>�}�Vc�v��Ȥ]nu�ggG�5�x[�Z�7�(�t5L؅�%�v#3u>%'l>wTۻ�����r�
?B�s��R�Q�jfjUh��km���L�E�Uh�X�*Ҷ��l-�-,�-��\�2 �J�S�̙��L�R�ʠ��əR[[e����DfR��1���j��V��j�r�8!b���U2���\m�Q��Qm�cE��b�qm�G.5k*�Dpd˙Je��.4LEZ�X�V�X�s���rdr�9*[)b��U[��ڴ[Km�Y����b����rʘ�2�-W-Em��3�0e���eeV�.ad��i��V�A����j#�ih��Q�֖4�m�8�b�j�Ѷ���m�Ur�lZ�+b+��VDDC�����Į���r�cZ�a����e
�8\�W-�E��ƹ\�.W ���DQr���[%�3(��#m��rܦ%\��[u����~��W���epwt����y��K��/��f�w6�4t�_�]�f�{�|י��?��}y�'�'�;|?�y�jP�]�4I��~^��_��Y�#{a��\��f�zۨ��>�v;����_��f��kx�~h���6�����yG��X���ϲT�����7͍��w��a�_�z�o�'��5�ή뛒��9��ϯ[z[��������lF�<Y�=��*o�~������::r��Dr�Uג��:�/Z���U������ȝ��o�nL�ڷz���Ç���/��c"�^���`kk�w�,U�/H^}Q�=��_7��F`���Σ�3꽇�x�x��>X�/�+��4i>=u��Q����5V�R�_)��α�Ꮎ���P*S�=[�\0f#���m��.j$ۢgj�z�*���e
^,Rxi"����h���(��$�	U��K�.N���Y�����a.�1F�V.�Q�d6��ݥ.�>I4�ny��w3y�k}���������O~�_϶O��_Q.�f=b��:�C����Pp:��}$+�b/�/ U�O��q���)��PeA��(G
|e(ɨ���hR��g��
�i����K���z���t����ʚ�g�e�^�JK�>�8����i�Rv��˞�\���m�Pv5)m���g:V�JĆr:-��z�;���$�{L�w�Ҧ����+�U��D����:�zs��w�[c���םgعey�~2�Ӭ-]�;���9�_���A{�^{��};������E� ���u��c^;��+~�w��v���2L��Sq�"��R;���P��	��:&����qS�*U����%��Gܝ��!٧�tq�Y:�u��ƿ'���}Æef��#��tB�~��w^�nK��*�ؙs�������ٮ���J��A����};��G����}C5��Ů��]3-�^����=����Y����`G�,��;�*��XB5{��{�������Z��/�h�s5ˑƻ'δe�W����v��{+D��.��$����\��pzS��`�ѵ�Xe/glZ�~��:���I站=:�[�ծe
a;����1)�k�E���ɺ�6��ˁ� �aN����";�f��1�:�p�����mwo�*�u�A�+��1�|'�_;�ql��Q�v6ˢ�9�Sz�k��{�����\lt�w�SdO�����ꜬS��b�;U�9ܺ\ǽ�����<x�v=�<r/4xX���0�[Ԥ~��{���"IF�fv�~�W���e5F�]�vZi�So6��aX��!���koR��?QE�v��T�Sq�s�f��Zѽ�lA8:D�k�܆����Ӷ�v�U��]?�}��}����������i_N�����{�A����&�`�v�s��ۥ�ؽ����>�:�ï�t$�<ۦS�6}�&t�{��geG/龷�/E�F|s��k�bS�.j����6����ks޴[�ۣ�ܕ'��������.�J�7���:�g��^I���vz�:������<�he>2���2� �b��`�Y�&�K��8��HV?������`Ď�f<�D��ں��-���
�/���gˑMe6pS�]N�gj/K�o�ǘ�����W�zЬ�D�cu��hlS�&L�8�=��m7��+L�`,�3�Q�:;��x����1q�G����-ƙ��4�^Ǘs��m�<�Չ��ι.�[��haYנ�vp`�����p`�Ƕ��c��F�ڝH�`�}\�=uИ�l(������-���я s���N����+vI�n{Z?��p�ӏ~�4r��J��z�W�2:5k�3���Ӹu���(��~3���{�>��ep>���R����&jv�8�S���xw=��\]t�TC�)�='����~��z�v{�S�^V���jn���f�y&�ϋ�>骀��/#1L�Ht�m���쿦���?c{�ǎ}M	���=͛{<A��~�6��l5#^�ǥ��
(����<�M����c��vN��j�mo�}��.��ڱ/�����ܝB�\��4�I��M}P�o��!���
|���[�1��띆N��h?{z��7�驩��.�t��o�޼O�Ek���h�Cǜ{rE|!�%Ƀax*,�B>Ɉ���
<�P�ɣ>����-�ɺ���uaa�'�­i5Wr�o@�G+����Jl^�T��9��fw�3�ܞ���}�y��ޝ��������;۽���\wo!��3��>��@.��9�zk���;o#]���[h^ܺX���/>��3�����Ō����W">��Wzg}�u�h�x_�(wf�؄����ѵ��v����:\�h���U5�ƫ� Wz�R�c�ƙ��9צ<s��t��V��0���u�(���0+�^I�'�o��l�H9]�юS�{
�Ӻ������g��ݯt�KվG������Td�fwݮG���>�["�]��������qxvO^'i��τ�)�N񆗲��V=1�:.i�:��S~θZ��uǻ�v�x��{�>�KZ�/���Ɉ�!r�{���YX���h'�n�쀌>p'�s��_ }7?t%\���Q�ң�xf�uK�ι�zY7T���w����y��َ�To$��s�ռ�y�wfg(����c��v�����}��_�>���)=v3�,�{�	}¯υUǐ��΄���'s8��l��wy�\d�:ƎPS��ud�2r���z3R�=U����]u�+)EW�w��uk\�b��=Olw�}cc�6�;qZ(]H�fP��d�J��[]��Ծ��*]g�a�ئyZ��t},%��oá}{|�T��=��p�q�u��V��<q��VK��q-�vtl����V?�1�U���hN^��~����}�%e���/.�Ո����/���cIõ�BU��J����{�i��3��R�0��e��4)��p�L=wJq՗oQ����籌���U���;Ka�J©�|+���^��Y�Y�%�>[6wWs��a?K�h���\1\�r.�y��Ӗ8�d�r|2�������aN�����Z�=�N%��»+'ׅ���_+���k�VWC	z�-86�*P�<���=)ӎk�մWtܹ�WKz�<M6+��}���������qo��R��r�N��U}�yp3�]��I��P�����u0�ːz�~�Gʮ��ֲ�AgR��{����:s��cxWg����ݝ�����t���m�O�&K�}B>x�{b��.	�WƑߣ�=��h�ӓ�(��ޅ	mob���~�s�/{���Z�S���'7x�<E�����z9�T���׻��{�>ع/���{�͔=-���;"�����S!#Cx�����fn��}�����s��g�ѡ�o'����a��W�ai=������V�}X�g�/_�/4nR͛iw���sO �5#����4g�C㼯R�����W�8{�v�w��o&#2�e�l�읖�&w�+��im����J���Y-Y�9K�um��u�x�N���=��oiwLYϿ}��_U�;��y�~�\�R/����t9>�ch��%P��Q}U<}Y�˓ռ/�/S�5r�j�^�z��\�SYM���bn>N��/غa��M��z���Z�hWOS��K�R���;��3�w��Wt��8����#�'Q�_V��f5�S&Ynw�M�6Ƀ�P-���U�gH���д�N�ۍ��{}�C�>�eѶxf��h{���-2�Z��9��,3���M��+��R�M}�� Q>��T�U�����a����â��옳�:]�W�F��W����"�N���,gB���U�,7�2��b�;��7Χ����۽ے���=��'c����o��^?m\V4���4 �Hm++EDt��`,�=o�g�Br�@�읺�R7�gn�umZ�>ޣG3�9Lr���q�}R��+S3;{xEܫB������s�}�ϟ?����:T��g�npV��I���|�{&����]�����o��t�k��ʾ�0�k�慱K�V�v
��-[�WN~��v%���������m�#_��t��ͫ�:^Vm�#}2�Y���_ny�>t>kG}��wo�����������>���V���rK�&M�Y>�S��W�>���P�����X�ʈ�ΕF�N�^(�{�&��ok����7�Ǎ
����5Y�{��,m Rr=�o�wx;>+�h��*�T�������vg6�/��/]�{���hȍ����s%���,��5{C��Lr>�n�>�h����]G
��^��K���lUv[�ϼ�^=���Nq��h�xʎ��]8-/8��o��=�Y�{���ெ:����g��b�&T�Nւ �IwU���J�H`��]��j(L��=Z�R���ᄽؚ:��B���!�.���o<�V�R����w�ǴKnk2��|�!B�ڣo0�Jmv�K�dh�+��8�y���qlt��]ק&��N���:�!�w@,N���<�K��#�i�)?��>�B�(�����Dm��-v\ጽOi�R�9)^
4�����D��W�+^��ĥ3%E�vsM䮥��/��)|�"��ޢ_�gQ�A�B�^ޓ��ݕ�����V>:%���#�S;�x�ӬV���_"���"Ҳ��&�!ĝ����8]��� ��i�k�sP���L�Y���=J�;+#27:�c�_��.��V���e"-L�ca3�.���n[�8fu���\6���א�<F輛r���vK���{fV��ϒ����0^��k�ަ�,�Z��Hg>�٪�U��|��-B�kk9��uC��g*�ۡ]�:�E����o,�:u��G{t%(�;e��hڼ����!z�o�:jV�`G�J�<h����P5n��B��G������ΔD"+9�^� e�2*�'_�h��~ke6R6)�
t:�kڶ�M��P`hE-���O�'Qx��0J˵�{���O^Vz��2�b����1މ��	�l�[�օGi��)�e�A�)]�p�>�|���6+����MU����$BVVZ�1e�WwJ�7�JDS���d6�=����0��!��ܮ�n��xAȯ9+��ʏB�q��L��+L��Z:q�ˋE�JD+ ��,��^�i�QI����]���o�Uo/}۸��nX����b�)b=�݀pa��P�,X}�:��K6���;��S7��ϫC��z��*t����:]�7�o�����q�Y�tsb�/�q;���^��3�o3��ٰ�{��#����ڧْ6BއM�zf�})f�5D�}\_{׭��F��K��b��j��U]��y�[�6��Vv������������L1��**V���\h��!Z�
�UQr���2ԬAVڂ����neʍ�\r��J�mU �Q����R����rۙ�T��b\�A�r�,�J�-Ej�Pr����J\��Db*�cQb�m�cE+-nZ2�8�W2����q���*��̢4�[neTV��5�U�ܸWp)r�s2☱n.c�R��3.UF�\�)ne�LF�72X)�\h9h�m�"�+(�R�.2�e���PR�Ĳ�0Q��[b�Ak(8e�-�U��(�h�VbdP1�����.Z��V��\�-�KKZT�+n9����X��J�Z�̥d��V!l̢�j�Km���s.Tb5�(�EEɔ��5.f	�.,ȫ��U�0J��1�ڢ�-mZ��)~?U�(��Nic�|yK-��n�����s����%c#{;�Oe��y�2G'^{]x۫y����}����q�/���)y��_p�1��)S��e��I��]���%�̂�R�y꫻�'xkT�e���a��)ʧ$T����L�Լ���еC2h��c��t>�y���x�߷���災�r�}�2OoB~e�J��|��'��Q�\�;%���NF<�?�����%��{v���=�{�{=��2qS�h��ݯ{��%�D�9.�^���~����*���AŤj,�����{��]��:�=u7_�X�r�V�`8Ǖ�W/�����(�����)�9E����8Z"������Rg���|�Ң6�>�r�;=�V��p�^��{MLh�*p§>�6��د���b���GVZ���T�\5ؒ"̸.̷,��ٛ���c�k;_on3���Q��s��C�tj�k�\c��r뾲�Q��+:H�3x(
��Rk�fj}��ʳ��5s.�Tޫ̐nɉN��}���ķ�/�n�)������h[��5�ni��r�ʺ[������By*��XZ�a��'�yJo6���1�[~M��z�<"p����8�����]��U�A�?W{�?>(W�pua�c�il!��RC����>�\�w���aO�'�+({��>�CGg	̬���0�B6��L���0v��Oc��Wc]��]+|4=㓐,���t]f���M&L=x�֝���Ge�Y�wl�/m�vD��dQ�BH�x�N�zg���٠��>Oz�����}:��U85����i }'�P��;]��f����:��Kt.p����n[~�v�93Z)��[�ٜ�]n+���w�zSTp]�0��PyQ�n��s/��	����\i^-���;�ձ�6�b�ޭ|�k�?�}� /9�r���֑�)ܝ�͔=�{z��z��f�h�ؕ�t�������4�U�R�t=�z5��Ϟz�/Uz�zL�����sC�J�xQx��R�v��^�;�Z����I�vy+�>i/d��~���W�a�^��}���}���ڀ�_�z���z8W���n�I��st6";�v��Φ��:е�k�ί���:�����c� �ԗ��-gg{���%y�� 2�����k����t#�η[�/:�<�K�~�Gŉ���miu,,��A�Z6S�f�)o ��&Æ�0��޺�<mg!#X+8�]a�k7Ӷ&	��j�e����h���� s:��z�����1F���]P��i���
� T�fk�מL4�Edk�<͋�ܽ��d�*p�缸�r�c�Dԕ�RWn�,wW=�֜]���We��\�vyK���]�}���� 8���oq~�*�����Rq�u�<ه=+�Ԝ�؍�[��Y���]�'xsT�k��1N:���E��ܫ��6�gc�c9�./o]��|˪��KK׻y��6Ӕ�����*��JAt��ٵ�罍�"�S��0)�x�],]b����ss�~��]�3�k�f�*2��'��U�_�y'�͹XjAv�Q������/]yf��t�]M��tb�<4)�����%�{Wz�LA��y��d���Ύ���m����[R�egG.u�����Ж���±f��.ݾ�cVvuU���:����8w��6�ީ�X{������T�����n�3�9��j3m�]��G�y�Ǵ{4:��9��ԹYA�f�h�[�Þ�:/ֽ~�Μ������,3��>��B�A�X���	�ۮcM��X|v��2�f�!9��rNw������f�G&[l���G�ٷ�t�c��'�{���oz{d��'��ę!��k�K^Ձc��T����tW`E�e��[���[��s%�ѡgB�wg�g>�����zT'�����#��8Vm���r��y�9�>p<4ަ������p�|e!>�ޞ��a���_�t�Os������|�-��cc;]Rq�8$9���{s���N�p�W�<�}j�c�c1�";4�~�����L����?<R^����Y�4X䗝��ܹ⮞����Z=��H�X~¤�u��$��a��S@{c�{��ujћ��'M��31�Ɋ���߁�r݃�;C���&��ig8aȯyoX�9�TQ��p����O�v��u�`�y"����������x��v�C��M��ޭ
a�Q��w��RI5C7b4��FU�}Z��qeu:`�����T��u�wPYO�+{��tS�}_| �f{�q��w~���;���_�{�z;�S�.��fY�������gc�3<����=�}�6L��z����{�é'�g]��.̝#�u�����s�u�h��'�����M�߽B�[�Νh�Q�{�n�T0�5��m��Us�t���s�-�0��^�4��d�
$PcX8MvW������Ԥ����_3����a&݋Z�2�,մK(1[T��N��]������Ϣ�cZ�=B��X}c+�Ua4%T;���[�hڂ�V�vn읝�p�	CD%D�>7����YQ�Wk�A��A�7�Od�ۃ�p�a516��NXO��[,���b�i	W��G6�hyp�=I��'�Q_{�2 ��z��@�s#��W�҇��(u]аl��Ȍ�T�� �M<�.MU�u�G����M�j�67�g�ߔ���-d��+��Y�S�.��ާ���n[�ڷ�Ff4�wR*��5)�Ͼ������rV��y�˴��-CE9-�`t,ҝtiG�/���	B�C1(Gu���f,���n�z�_�;�m�����,�z�i'u��P���z���"yxX����˭B�@x�C��Rvخ,���d+^õ�s�o��5����Lٰ%iWɃbT$�x�_���WSα�]3Gg��*�ܛ���s�~�AT�X���q��B�Pʭ!�i�뇮�7�e:�^�&��fY���%�`Aa@�2��o���	���ߗ��.]����~��kǯ�/�S,��rf���g��>4 uJCj/.�}�{%�����j#�r���R�yY��;Y�R�\2��� e�A��Yܞ}-��>S�v�v���/Qp���M�\1�]\j6��W��Y�e�>RZ���X�J�X�v��W�3��^Y�zex��d��*�y6J�O�5GAV{k޺�t*�S���e
�@^Y�#��O3=U�!��^y�yy�_vS����m&v=A�[m[�u1�v]l�:�|�%�]͝��ю�l!�r���Kܸ=*�-�:��������z>�ۛ�g�)� ���&��?bg��,�-|ℤ�f<�����=�/�7=��DP3�H��l.U*�����q�����As��D�
5�����Oƿ���$�9~5a0�i+�v��ʺN�_�L���ϤX����uy=������LU����o��U[�~Tau�Շ�,L:$�t���:g{ֻ����]���P.�ب�Y�H>*s����?-���2�F�l�����v�GC
��d)!�_?lV��uC�Y������3=�\�z?s��8t���AO&X�I��Tȫ���Ϭ_Tx���yc}Ͳ�B�C.h�++�~ʫ�+
փST0�T2�_ǟ��*��q�S)���Hk��+B�v�8=mC�w���=��_z=��k�7>���x��/�L�,m��x�F
��R�Vq����q�:BoV?e�'zi �8q�Ѓ^��j�x);��i7̝��(9%�vԨ��fY}��5�ڳ�;P���m�lnKy|d��������6��2A���|�,�g�z�������g�k�2�١��ޛ����Bf9Cc��V9�f�D�^����/{�Ev�?;����wSĊ@�.��vz�p�+�w'�o�~��gj����1����RP�k�I����Bl1,�>t~���q� P���3g,���s;���=���XF['~<���V�)��GJ?-�3٣Ȋ�r���ΫE��B���Au޽8&sP���L86�j~��.X�#���MAy+u)U�੼t�B��+&�#g�u<�T����e�y��Q��͡�R�\ w��b���a�b��ZVO���/Q������`��3i���8�(@��!�>�� �
-��H��y�F�^��=c8�F(��B���l[�"��AF�U�ʥ#����)�:T�eQ�2��s����"�(��ۊ�<xJ�d�8f���4&Ӭۼ���|Z�CX��y��
�|j$W�ڇ6Lv_6G�y ��^��Sa��~���Wh��5���#e5D��Ϭ�AL��[�v����O]؞ۥ��ya��݉���}��}��{_OJ~�4=�x��媫����)��4�%RBCæ�pv��:��ϩ�@Jx�~��\�dv��VW�<��>����{�w���+���g��VK��P���,!��ק_���"���$Qz�~������g�h?k5�<�j���gY�cˮƖ�>��aIy�2_���}U�͈�
�$m�]ƼD���틋^ڷ\~=վ�ڔNH6;��6 �MZ6�Z<���yq"�!��N��?1߳&�_e�~s�7v 2}^,P��a3*W�3�D����#�]x��VT�{:&�o�Ȇz�� s~C�_xB���%��k����P�����Σ~j�`Ƕ==�-L��[�Å:f�4A	?i�4HkD�7������y�6��\f�mX
/��2mص��C/���d�W�V�h�|��8��m�v������ּE&\���Z�V%��u�GƝd�ٗ��舫S�����n�M�G-�Ђ:I��g�Yt�����->BN�N����G3pF���)-FL(̕�}5��QXL��|jL�h�v+�a۲&��kxHxuP�So��w�k�*r��q���Dm�G� -��b�ON�a�kP�R�H�/e�v�Y�څ��H��.�m̔�q��c��Ӕ�#�dl�U�p.�>v1�7�e����L\�	\�M��+-���VH,��uj���4��L1}κR3{�EBX��ޘ�P˖7s�7:=w�R@��d�(j26u{(��/J*��ц��0�.[J_r��:�q �Scvnh�d_z�!n�Tlh-v��ĭ$�:���dd�r�a�Bڬ'5�맂�!b�B���
ܮ�|�.V�S���vnO��َ#��nP٪r'x�|���O+��;��P�ԂX�t1�	�JvvWwK�g�(v����L�v�"�@��S��v�NvvN��vEVJ��"(n{Z�\��;>T�U���82�0v>��nʸ��w����Vw��`⢗x�Q�#<����@A��Lԭ��5�ݣH^SWR� �LU�r�����YR��3:3�R;}5�+(�����e]@z���y���V�f�O�|!b�2�u��X��mǷ�2k�����1Ɏ���
�Q����Ѳ����k�1��`"���.������[��o0,�, �=E-��t�,a~��v�g\��$w�%�[���*6�־�S��ޔxq7��;��+EkgeՄ0�9a>�C�T�ลzM�V�F����Ψ���iܨҖ�KV]���B��k���t�=�p�r7{һ/�c�v�ЫkW-�pcv�.�!1%�n�w��3\�V(�dr�
��U;PܦW���:�Q�J���V4�J��9wЗ��_K���D¡��Ò������8�Ne��ۜ�E}7���]Ů�i�])t����[����!�܏T��P��}N���$'�k��mME�gm9.�Xu�#����ξ�cb2���+��>�vVrԯv�2�C�oQ�&�s�ź�Q�#��\����i�{�~z˅�m�Եh�2X(fV☊*�Je��T��Z`�
�F"�k�Zڥ˂ۀ�V���c�-�K\ʃi�P�KL�h���1�h��-�L�U�T�����U�nZb�h�m*�4V�ncQ�2UV-k���q\������lSE
�U���k-hَm`�6�c0�e�U�Y�ܴ���P�Z��fc�E�,31q�h��j�mUQ�)�"e)�fG3&&���+��KF�j�\��3-����X\ȸ���.3.9�D\K��4̲�2��p�R�Qm�Թ��61��pV㋈�ˊ�kq����K�1�9iC31(≅��J�cE)K��q���VZ�-�%.S\1(�+��S2U�.6��9k��-\�jeɈ�U��a�e*�8մKG3E�l�Q���-�Z�̴�婖�
��ff�2ԥq�8�\iLh�[�pL�K�R�30nmʴe��31Se��R��\%[nR�2�8�kV��m���6�\�L��)m1�E�fy�5��Q�gh<�v��p\���}�ǡ������|�\�����t�O��ë{yַ�����|>=��p8��%�㪿����u�^&[��^�������_\4Q���d��U���oOkٌT2��D ��gM�h,�Y_F�_y���wHa<K;w޽��}惣Q�uV�P�`�>'\��n������&9ӽ@��2��$�v���*=8&4x�4\;�HW�٢.�}�OD*b�yk��J�D�\h��J��Y�ʍt~�"��Kϒ�8�e��;/��.��k�<�?>���p�Sϫ@r�H�P�X`��i�]"��\2j���K��SQ�狫��U������8zU��k��)���1W}��WTG&3�M�`�J�������%�X��*��x?O{�3eգ�鏘(�i��:=��mq��W��r��#ɞ�tr�kk��Q�:��\Y���^�� ��������W�i���S86(s�Ўmz:#��\4����u;�(�V��=6�G�˕���sJ�ψ�����[�mh�i��;_N.���TAP�v-;�E��Z5��w)�v�̮��S�_7��!��|z-{|�ؔ�KĹ"��ۥT���s?W�W�U[��C�s���PC�5ٶ��|-u�p��f��WE����PQX�p{�5l
��i�:gU�_ފ����žP��Zj��Xe�� �yT�ݼm����b��,�W^�����Z���YA����h�(wU]�VB�k��Q���+�XW�#��ų��"J84,�K���0j��A�K������ևUNи��WUS�,]/-�TX�����h~�75��d��6y�
�ܡ���6�A�1j>!yh���2!�R�� 4���NO}�5۪�5>�(֟:��LՄ±��P�J�Ф/�ȇw����Η#p��Q5ZI����wʨ��,�	+-��pm5�:<�N>�ۃzZ1&o),rR �,ʬ��P��th�+�{���r1[�5Ix�|}>K��/�6Rb�ea\_5�XV�uCa���jT�[}�xڡ/����F=�aY��@fxk��D�I�[��(����׻+�:d�Z��-B����yCϗ7R���"���9�,�ڝA:�m���Ѻ+�(�shvL6�l|�I����nNjN��U}���w�d�����
�8W���ޫ5H���5��oR�1�<�Sϛ�vֵ����.MG��uY��[Zچ�R]�U�w_��m�L�>X�̊eq�5xՎw���0_���H�x�-�:s.^�j�K$����!;z�w���P|��V���������LU��4X���o>��v�x�_�|f��nuCs��uq�.��Au�>"�Pc�J�mz�۔����b�8.�"���"\Xx;)3�F��m�\���<�lC(x������s���(`��C�G�������i/`��t��997ѽ�[Xz��1��Xഞ�.���ơ���DX(�Ar����v�_)�{�P(|�U
�҇� �񡋽zp.L���x�W�W�l�_��Ny��G��q@��=����r>4(��G��|����*u��e���Vb���ŹP��n^2w�;�?w����7c���Z�ǩǚ�֠�ְ���f����4�:�D���LT���dv��mN=5n*��e�[�vuo�e=�������|�{�[�M�#���3k�:�C��L�L���SEP�B:{6�^o{wW���4l���r�Mz��L�=ER�D	��ʅU�a�\���;s��;>�F�-4U�݇�y�[�+�N�^_s�f�{�}3���1Ӫ��¡�t�H^U��eJ�������	A��)���_I��"���4���w�!q�|'��o�0E?�\2��X�3.{�˷]������,Gs+F[�\�dЅ�h�VD$���H�qz&x��g�C)�3@j�a��9�{~��(�;c��m�䑗�(��3�hA�:�᯲V�ˌ=�tG.�C�3s'-�Q9�6�����eW7 A\D���ꯢ��:��l@���zS=��f5�g'4U2��]]zV�<�ldL�ȝW�G��u�z����h�.���	+.�t�_a|�TEv�Lp8�	f��3(�n�S5ݪc"���sx9�>}``�2Eͬ��Ӭ[�*p�y`������n�xp��_b}w�d��2n�,������ꪪ���Ξ��_���$̄�b��g�.��0;���_ϥ)��/��۟�8�=�/C��i�L���pf�c���? W��1h�>��7�	^�1��IݹӒ0z��Ʊ��q߇�x�����B�Q�a�N�E����DϺ��;
��|��Vz���r�mP�k�����g�%|;s�΢�="�s��h��@�A��]v�_K�NY�UǨ]7}�ו�zfMO��t@���LV�Uƈ�D�:l���e�� �6?�����o=��ιP�`��(Ӫ���W��:��a Q�� G8"��~�~q���l��
��
�\h�،V�h���%�f���z{�_z[n��'n��'��3�jf��J���cưr��tGex��([��/x�54�?{�;��:m߈�P��0P��)t��7��,��'!�ޅF�yW�����́ ��mgf_����!͋⮵F�")u��٨���7(mk6��+���Y�5.�p�=��Q���,]�1�+�S>�:�X��:^9$�s�k���KŌ���wt��w����/ۮN�/{��W%q�S)�0|GC������,��v�Q{K�n̥�K��y�i
}�
��eW�<|t[L�%ex�5�M�L��X���s=�ٜ�>Ɏ�[-��|�tb��B㉨Y�UO�B���������T���*2F��Kj��|��T;Ň[�fhw��կ�̷Jc�;i�է�'���ŃǄHThq��U9�F[���펊\,�w�P�ߔ!w�������4�u�o�)�)���&����ũ�����| ���^v�zֺ�hf��d!�n��Ѩh����[��ϣ<8T*���
�Z��>�f�Y�Yzx�P��l􎕢����4���e�LПt�T��`��AD�9�)|o|���k��Ķu[����Ͷ��N�ٯ
��Ek�*0�<ള]U+���9���j�{Ui(F����3�zE���d`�A��L�ǽ�<�is(jb�Ι�֩�oh[���yGK�1�.���ҟ+�
e�^��1�r�躹ש=����{�oT��W}QJ��mxk�_���� |Y�}N�=z��+��4�۱HS0#�/���
����ƌ��n5�윺1Z+��!�!B�}M3}�2� 2?]x*�,f[�7�����ۼ{Ι��\˸sԋ@�����W��P�ʍ�3y�U��oY��G�6&f���nS>wl8CE�Cb����:�i�W?wvl����<>��"��S�8O�U��`�L��yIR���D�~���xL��`2V���sE�Y_2��Xp��փsT0�i�O������g�Õ��\{]���Z9ߍ�+�$�(V�6g:ջ�k�Y�D�=�� Йf���3-��W�v�S,m��ª�#�w��1������pW�C���;�{�9<6c0�7�6��[<r�v��`��p�V�*��i����3�+L�~}u����b`�[許.�T���^y��P��ڿk��IY�9�0'AF,�%�A�-�`ݙ٠[m_oQ��b{HI�̶�о��՝if���f�u{γ���(��[���3��ӿ}��UT�t}�ޡu_�j�|+�B��*��q݋�:{+n��+�8�i0lcA2K�i�d�����*�4�����aiB�i�E�:5�,"��G�8osKh��^F�<�3g��k���B�Pd&�C��P�ŧW&s>1C=T���V���v��,��i'°N1p]3Cj]X���Q�E�P�1�~�gi���Ni�x<����!�Hq.�#]2��٫;7B���i�{������K���mP���3�QT�K��6T*�1G��bG;x�i�A�x*�,R�RU�'�'j�y�XtH�0���I'�n7�$����c*���t;A��E�&�? _���PbMG��s�G�e�{M	�y,�R��g�?y�Z)��Yg^X������i�3|��Xf����%0�~��ɨ�/�H�'�|v���9�`b�JT�ӝ���~��lU����i� iy,�H�����Ȩ���sM�nԥ��U��!óV��GWN�^�{8h\�n�F�t��E�Egb�;^2�,z���b��{�ݫ���f=v���� |�|�/Ϙ��h?Vy3�m2�c�p�:_���Ju�$p���節�4p��T�|��>�VS:�-3���d0C��zd�fr��g#KF_��C��D�0�()D�L]Ƽ~��=�3WG�a�w巻�����j5�i�.0�nS��ӣ�jN����~��>8Yw7�mU��
�*�����:2]��(��^��T�Sѱ�b8�J�3�G�߂��T���n���*g��B�;�r�|{*/1��ɨ��.U�g-�;(^�X�z�g-��Y��d��0�1��k{��^d�5*��li�޸sk6�5��d!4]��(]��]kC;��)s�{Y'���QP'��<�|Ў��U�xԯ%���M��7�ܩ�2�$Ǎ�P_\4l(.�`霗"�+�gJE3���*���i�h좭���gm+�����]Im�B�";����Qs�$�x�J�oS�ѵ£5Ȕp>�9
�T�ݩ�c�c��q���}[��,H��歂ܼǉoa�j)wϗ]�Wkf���Y��T�1y���� }��V�s���d0��c���2�S
�V�Uiө�H���F%-���H��0e��*B����\h�ؚ���^U�CV��Y���/7�t�|0�U�|�����%J��58�[��v$;�K3-W��{�?ޟ�?���~�w��P���ꬰ�Ĭ,�BΜ�7��<�~�*�:�*�v���V��=A��t/�d���r��yS�:>�y����y�#/�
�/ļlܭ7"��I�םuV�7d��j]�gOt%�Bx��W���f�t�0~F3N�Z=�t7P�����z��pŚ����O?*�=�Y�1!"�<��uz,Q��R��O�{#�L��m��[�ʬ0-��q�a��lh�ˇ}�AUG��H�4�A�T��w,���fU��u��-�0�ֲVlP�T!?m�|�zkMo�����6.�;:��F��{S\�v�G�m�`;��p����W�Z��m�b]����w��$�hok�;�y�B�1R[�<`��0�L�)vں|�u�y[f��rL��a�&l���1(�/���K!}}���n`p��V2֕}���oL���N3R��0^j��(�j�ٔ6�H[#^�%����y]ۃ+'i�L1J�%Q�ܗ��yW�8�;.��)u6�t�G>�׮�g�C��{��~[�-Z"�l�����͡j,��˫浰�*f|�{,���v(�i�ի���gO6�9N�[y���:p�\mՆ�M�ը﶑�i���e+Y@�)ks>�y
�'s�\�^hk�16󱽧�~ȵ��7t�,I�M�֓�m�%P��oz��h�ۢ�ep\�ʇ�%r�T6q��[q��{ܹ���q�+4��E�Fo%�}'F�,�t�Wm��j�R�ޑ.c �3zq�����h�V���f�5{��4�V;�r�*�Է�sV��NLw��Cc�`�P���6�u�Z�e��ٖcySF�q}�4�1����G��;v�3�v�2������R�Jjor{�����32��T�qj0��V�FB�L����a~*N*�E^�'���k<&#o�1*�9.8S����Y.���<c��+y+(lU2��]�3M��@�K;1R/�e�����Q�0��g��d%[F��G�t��)��Iݿ�缍1���^�O֤�Z�b�G݋eYu�UK���dI|�k���ٶ�SN�K-Q��R���u��n�'e��)��*;�j�E]�,��;mva�b�sғ�4��G�L	�e5�{QlaՑ��)�=�7Fv����]��vו�o{kr��c��L���p�n�2*�����b����b��gk��7b>,w�J��'G �VlICW}�z�,�~�Sk�t��M�����J����=]�)u���!a[�Y�2��T�dr�yK�����0�:̈́�k:9�fci+zn��Y1V�ER�{�Z���*�D[�h��K4����Xg��� 1P4y$$&��vn��ûD��0ؾ��yƵ;�%��<�+Yt���e���{��6	k��fv՛��-i	N�\ǎ��39+�K5%�����vx�L��[��k�
jMx�gu�ڼ��kd�R�;򭂅�Wq��tS��R=��3��t΀j/�~A%/�*��(���m[�\Pf�0˒����eh�U+�ۆnc�je�%0���PS2�2���F8�L�UR��)k��pUµD\b+Q̦U­b[3D�����I�ĵ���,��������L0�"ֲ��҅�e�2�1�3啕U���%�feT\�1�Ҙ�q�
,kb8fU�)R�T2���j1���r�Ŷ��@fP�+�5
�%PT�pƭ�G�f-�*E�〪��k�G.0*���q�j�J��cV+R��+-+�
+
"�\r�����mE�Zfc�R\��TU�X9mB։�1D�*[�Jָ�U.X���YD��j*��UY
�E++R�J�m�U�  #���.w�HO��'�M�יދ��+�������-��a��\YλpNԾȴbHgH�%ӿ�����_Oz����Q0t���fvԷ~>�Q_
8k�B��xix=��Y���寷Aߎ��Q��.h�D8�1l�4X�%���!�4���3���k�8���Y�a��AP�v���K8��
_*��`�z����!�&򝙨,���C(�|����VK6�T�+��pY�Ɍ��o�W>�{�F��A!�g���8�:��b�߶������2n��[���{�P��"�A��/������L�v&U_�X�Q�<7^ey�R�Ѷ��N�c��Q�"�}P�iC���@�_lTC2��Q���=[�ѐE���Cc�����U�����u��A�Wκ+��GY[�����\1�qh�,<��U�t+4�����-T&S,p������ˡw�3�oZw�O���kdZb�3�2hTl���U�+
������f'2��{ԏnc|V_�&�|jz`I3�ӽъ[�ǪBj�]���F�uO�Q�����CY�M�è�{�9�Љ�ża�F2c�ZW>ꃘ;C�]4�u��|�%_cH��/U_9���UW�Q(%�gg {�ؐAB�y�3�\��s�N�3��N��>E�X{���~���B�y`fǹJ��3"f:���b����;���8|�;��35m��W;��1Tp�z��Co��T7:[0ؚ��J5��@-�z%5'��;C�F��%+A�i��v��=+���~��/nP��n��yfϭL�{��FP,O��C�
�t�Zܩ����o�M�ނKW6��|����x�ЙL���� ��z�ʯ
jơΫ#��W�
o;�Jnx����2�����.�_΃!7�O��w�N.L��F�j�S���n��5ŝ7���L��^������!��vc�O7����S�V��S#lb���,UP��:������#PHg��q���5DA=A/Uu�@���:g��HH�(z��
��S��h��~զ�B��jw�'npx.�!�dHb�9��o&^�,Y�V3�`��I��F=�8*��(�7�d�L�S�� �o���,��D�,͹3%����8��I�>�x�qͻk��WE�T'8����2Wi��k+.�v(��7��z{y���{�\�\��̪�h�P(lp�!��i��C~���ċ�G��&�q��]B�3�IT�ʢ��P�:^����Y���T�Լ3��۾�8Zæ��D��$�T-�K#Ti�A�z��_y�S�F=�����&����1u��>�.S1�T�ha��;��%�X�d�Bj��Zk6��;]S������P�q��ߌu*�����ο��!-���O?1W�O�	 ��_T�ﲇ�q�\\\���{�/$�M�oy�I�q]��:Y������k}P���=�V����zg�{z1F�̭�bW[cƍj�ĭ����_����A���~�ɍx�WŊ:PyT���01J���WeC�j�&Q��x�&.�_��,g��)Ֆ.<�)���_�U3�Z>��&J,%Pz���0�{�ҥgSBfe�R���j����PJd��vْӫ��0�֙Y���D�V7f�"��%hu8c��v�A�fw���� | �_�c�:��ɜMS�y��/��m��P���YY�h�8�w�d�mh����H��i��b!�e��Y�`&�[L�6�XZ����=F{���AÀ
�G	T���x[,���a۞�m�ڪt/s,�^ێu��x�A�n�R�4R��b���!*&��(h�VQ,�K�l�_�s�l�0[%�hh+��J5q�Ua0��*��%��ʊ�n�-܃�ï�+f�>��p�f`�S�E��I���X�,�W�����p�2��0���\��T���<,j%�Lђ�Tt,�N�5��ʕò{wި��}M�:Xr%��e�"�ԸY*0��s)�T*V�#m� �����>{�B�H��b�u^3i�7.�`�����yV�%oי�Q��v��i\�|��+9q��Zl��뉃bj���il�[}{�"+�
�V��<�ڬ�y퀰n{�;0���o��E̨������\�R��r�}��{st֋ ���=^��7�ggG�s�fN�?�0���9���g�Ҁ��$�
X�VΫف�Q%;�UU�}B5�����G��?m\:=9^����5�H�+L:��5�6љݏ^z3$�����Y��=�xd(1R������Y\Gux-}��r^6�<�UC��6=8w� u:����x@�]�F�ٯ��Q�o�ܺ_��`ʯ�HK]{U�6/J��.�Py�㏔3:�^���;kܣWsi���,����j�M�U���|b��nE�kC݃m���9MC	�7�*c�w$�v��A)3F�>P؀�Ty`��L2tpu�x4\-�ݽ��kkn�������D�i�j��:�����W�=�Qq�4V+�����t}k3y�<�1T2�K��p�L�� [���L����.-���u�{��~M�qUmq�)�ύbC�8�`�e�P\�U��طF��`}hx�T����$Wו�]
��,A��U-�A�4O�.t.�:�_Y����οr�[�S�f�V_idC�-K
�eԵ���3s������$�N�d���X�Q����c��8��@#����c���ٽ��:�u��%�������/9!�Y$�M�S�W�W�f���ӣg�P�U����!n�2���u
��$J<LtP�T�_���.<�㬮�4d�"���	a��C
�_	��$tWVz���f��G��^^I)3x����t<-����$|��`�>k|�nS,Z�J[�y�ㄝ�^1�Uʎ�{-@\�7�a����F*�^6}{�+Y������Z|�3�q�P�b_�C���4��5x����f@�B�:>�*�V>��ν,PKo���tu���ϐ�([Ր^��K�>l���swn�u�W�޴N��x�d .�2���:��%�ơ�^�B#x���˸W�C��sZ`��4bDq���P�����M��uwƮ;��{]�^�����;�p�<��3fi3E-�]�7s��G�smn�wF��f�Y��l�t�9���A��xʮ���j��Gj1���\�w�l����>�W�2ę�z���Ⱥ<}K3i�w�CE�h�w�}�峩ڊ'C<�M\)-�ȉ;z��z.c��p����|K���5�=���7��N�ca���uj�.d�)��_rY��qx&��w��X����I{RjWn��l3z~�7�����t�ź)�cGבּ�D/(yr�hT����]GƂv��h�>�aS�Nѐg�޶81����줼��%��*���<h���-g�"-��S����B*u0��=l��p��!��L�E��]2��h�7ՅnX����N��|��tALX֖ͪe�>>&�J�hd	�vv~u�%q�{��U2�|�P�
��yq�~���/�)�X|�9e]����Ep��v��n�T��!��>�Z]���lนt%U`�$���ӭ�p��q�E!f��S�gѪ4��b,�jG�2	����|�V��/Zc�/*�E�,5.��0����U�C�&�/`�����s�)Ŏ�����A}i0E����j�)����,܋��_��X�%-���gio9ޛ��+L�K��8,q��YN�G�u__o�^����<FoQ2�f��P��Je,��u�����k���t�i� w���;|n:���^nÝ�IC���5����ړ�S�Vv��ؒ����T�⃃��S)^���8W�5Y'L>��	#�f�D�X�E0zBv���i�EA�lؕ�t�5�=B����o"f�'T��I�76w�9�hq��nT���z����0Ba.��*���z�۸I=<��zN�0z��ì�b�Ӕ-h��1��m���S΅>�B7s}5略���Ԫr��8��P�[\o�f�f���>Vaf��G��=��{��� X��D
44^����:��N�.Dp��}Ci�����=Uɭ�}6L�n��=ZjS$��uX�z�3�W�D,=�\��hmV��{�JU��b���GW�.����n�MCF�J�i��D W.��(!�o�)����l�h���5|`�� ��H�V��P�ojhK��M
Ѵ���oy�9�ݣ�:l
E}(�^P$��)�W�h���r��D5B����.i���J1��`�%rc�.��I"����N������L΂�׀��R�L*3xG9��o�ٖ6`��.oju/,���:��&��5��L>{�Sh����:����5���&��"8nwN;���r����Q�|�!U3�(��%�P�r�7�Z/��:�tr߷�&@d��w	WDn�X��C�2�c�`�VJ�������`�sb�GG=�8`�Y-�TP�ZI��ύ�b-A���]g��1��������x��T�<���J���P�֗�i�{ZU����k��#|ߩ�{�׶�`��{�Υ���z�U��*߇�F3�+L?�ih�r�1��пB[�n�;��j,2|�ʱ�GG*��a����<�z�*X
"P��N·�f����g_���^>q���؂q�q`���ǆ�כ�69��B`�������q�6(^}�p��ڸ�P��bu*��7��'����8� O����kCݟm�+��n-�`ߖɎHY������4xy�����5���l���σE��u�2�=���<כ���j�VS�߸��Ev��,]�E0lfl���J�Mb9�@@~ٯ�k]ۮ޾鸲�U�nNFw@��|[��$��Vdv�_&�7r�p�w#؟RjF���a�w[�w��5�BUxI�fப_(���(�����w�/��v�.S>)ViC6���Ƞmr6�¶���U)5���Xн_]�݇���϶���}\lxS(��H$9e���d�,�0�UZ��M.�ۓ7���q'Q]�)_��g���u���Y�� <,��X�,��|�p�9�A����ت��\i4��2��X��R�`Ta�Q@�-�-���Ҹ&@x/W��1xG[m��K#M3:;U�Y��T%��ٽ�:ߔt�~示������D!Nt���,�	f���d�������*�;A�nVΐ�g�-3ּf���E��*�Q������D�Ek�s|���'5��6��~���B��g}�;�g�*��p/�q���w-��\�?{��F�� /m��z�W�ș��6'������_|"�p�;��W��9���n>Ӊ�A'�(��Mm�����m9����n��ȃ��i�"o�.���C.���*��ڝBLUf9ѥN���^L��ɜ���l4rЮ@��}���E�c����ԕ�"���$�Rhݰ؟re`M���a�Ih��q��9��R��c���[m����+hu�*߻���k�.���m��hJܻ���1�o3�
ϗu0�ݘ~t�-��W��,����2IB����&K�-���o5%�&�55�F ���JL9F�aꛄK��k8�$�b}�v�_��e3,Iَ���#L�"���빽�=��u�|�!U�n��k�V@q�yoa
U���#,m_0٭j�M�-R��A4�t9�p���{J��\�|�7j���u�H���l�9I�.I�R��hX�,�P�46��	�	��os⨭"�=�u.ܢ�h'^�t���T��N�+��q(y�;�����ZVO&�˔;6ޖ�~��M�2�^�)�ñ��n+����J�����igv�!nn07�f�M��m���'u)��0/U=d�3v>��1�x�u�@c4���.r]3l�u6�c?)�K.�Ϻ��v��O���hU�9E̊ VR�N�rb�!��Pg
�4k,ەbe���p>������v��e�%��N7V(�)��>p
��f<���EkXyMؐ��9O��e)�Ҡ��N�J�+[1J���dZ�i�<�j�*J`�#�dq�k��T�-�ө!V�-ۭ�0[�� ����\�ׂ��£ܒ/��B8�]�1���GA�.���#Da�F�L���%L�-b�!��J�&��n�7��0Hd�:��G�0�LZc4�sD�.%��m����U+{�W6����,/y��t�f5l;,�yf�:�/��n��rڔ.VA���M�#���1b�|t�U�/��dێ��߷sm���^�&$7�L�6!X{87�x7V�l�8��ٗ�������
��n/�����H�9nP#:��\X�³���T;�j�B�� �|�w���$쳃;xAdQeew^\�Ԋ��P9�*ĒTc��6sC�']m�\��݌̏ ��H���3�HL�񠺙���}�����P�N�h��*��5v�T�� �k�$Ҧ!��V�U����ڰ1�C-1���E�F���m�mV�R4��mKm�AAdZ�Z�De��R�T���D��kUQT�%AIKAb���[b�Z�B��QH�R��UEmT���Km[E�mF��%V�J�e�*Q�*Q��--IQ�ʖ+mb�Q��(�PQ�Ke���
Ĵj*�Uk�IF�R�+QKl���j��J�6�6�j��X�D�����D����Ʋ����E�mmYhR�F�clF�Z��DBҕ+j�ԩEKK*UF�m��J�E�
���YV�Z��EJ��cV�B��h�m"�Z��	UPI�Ē�8i\����'=,�xtj3)&\�wA
}��|��(:�5�r�P=[:�<�C�Տ�H�P�Vw�&sw���ŗ	9�S�[�{����N����aN+b�\E�_ap��Y��X:��y�~������5�W�=�����@�-0b\e��Ɵ\�eq�e��%E�$��1%�/7�GNb����&};m��
�K�3���8L�ʬ�~����M+���^i}e��l��Lཻ&���x\�ʢ��o��[{&[~�Z�; Jύ��gOؼ�MɌm�����!Wk1�|�'��ˋ��Q�f�	�7զ�g��kL�)t���(`��k_�y��f����3� p�g��&4��)T(��`��"dn&o���=X)2��LN9:[�t�W��/R��AL`�K	��%eqβ�8�H�!8|��U�-3���k�E�9�����3b��d;���Cˍ��%�X�n�(D����Tl�'���H��R��|�R������|/h��IS��1�r�w<�ϲ�F������Y�ͮ�2
��"꺚�f��gW^��`���+T/�rB��W-�pK�K��sy۽���*j�s�c�=Oor�8z�x��J(���I�Uk��FïmC~��Y�7��t�*yY`���fd^2�R�\C6#��U�;Tc�u����\�>&�%��[u{���)��ڸ��٦`��g���]K���sw����zfr$W׫Kļn��X〰Ea�������J8���'{��\�a�L��v<��x��p�5Y����Hȉy6jv9�$��fWv����{-B8œ����N�����
��=��K�7�D���H����{H���U��cS*{�Q��5s�8%�L�+���=V��_���w���fL\ ���%}kB��S�`��V�R�R��M�sg�]�P��u��fxW*�1��/lu��P����:�.w<��`��P��
�Mve�C��Ӆ���x�0�Ϥ���u^_gR�f��v�}���`ӪRo�;W;��^��;�v]�4�)f�VT�jâ����w��d������B08_��2��ucņ���W;�z���1������:۽Yq�I�/e�AWkZ%��mR�4(��Mpvr�h�6�X�^���q2�8D�h7���!�.6��b���.4E:�`��E:R}*盔��d�06�j� ���8Ԫ���,ڜ�(K��U��b�~lG�i����wZY�4s����
,�3���\h#ӂz��&V�Otɽ2;�Oyx��%\hY�U�3��G��5�ڙ�%J�FP¥5�
�^�o,��=��پ�+�c���r�{.�:��"�A�4��]#i��g#��~���N���(��6�*7���W�S<�ά�3]A�]��يŶ$��yM�)�u*���s^�ɻ|�*�Q�]/	�a�K7�eh��#�~�T���53׋�ڈۋ�ь蔭0v{s��~��9�Wfz.3�eV�/Z�ߔ;���鮲*PO<��~�w�,��ɯ�1�p`d��(��A )�tm0���g!&����z3Hj��t��%J��]�S٧#rtef�iڭ����fq�Ք��o�V�<&�Q}͇2��n�ym#�3�t�9�J>�gb�����VV���ꙿE�&p��>,I�Æ�F�yG��ۢ䠟N���P���4�I���j�쬕�/5B�qa�V\�|����g&��s��BPG��D�8%��߃ڈ������~�r�����O�D��U��4X��C��kK�)�f��L�Ugn�z��nH�7��v��Π���а'X�R}P肺��if�q�N.�<�UOzp�Η��O@�'������lV���@6.������ٻ7�2��g�W����,�;��0��	@e�ci�I�ɚ��.�ø��p��y��I�a�
�A�Kk��B�ɑ�(2�QT�S4iS�tͫ7��.��w���c�l����Z,�#�\�R�7�,���P�wS�Qy�7�dUa�!\T�F�������(/M0�xf���"���Th=���*�|Z6�P;�:�۰��2����}�G�ȴH9`�i.�+���.�F���Q���ev����v�����8�J��U��ۛ)��`���K���k�n�|qZ����t8�'np�Bb�8Յ�R=���N*��Tp�x�<�An���u�d�ܯ�J�O��Y&Ĭ2��L�$Zg�x�=s��C+�C�E.�#��{&�w�WT�͌����0��VK�w�>|�TL�3�w��&W�Q>nT���W��xѣ�<��N�)U�Pˉ�c����VĘ2��׊�JrssE��N0gj�+�"ؠ4=���W�P�D�)WB��J�o���.�]*Òd+֙�a
�3>��	#�'�ł%�]V}��jI�ކ���h�����Z7H��L���kL�f�v�ъ���n�s��[�8vZ�?#�bӒ&u�wL�J� ��OV�T���u������)T�'�Mc�2}����T�	�v���fLcn��p��ﮞucz��mx�-�^O��V�+��MX<&���`�K�P��%��*d��?]%�����v3�q�iSL�:�����2��]bMZ��%+sp�ƺu���+_�k�Ve����{�ܮ�*+��Ue��Wr$oWX�KSJ��8�'o6�{K���w��C�����L�'V�N��� >�T�k�0"�)�>%>��C��D2��,�e�a���M�yQ�`�)4�y;7L�|]���K�	��q�3z���s���.����T����xl���<���US0Ѧ*�Vk�Q�%�Jv���^�����_�o2��%1P"��)N�ݩJ�'��x/~H^S*�����%�N���Xd�f����-H�_E�a���=Ȃ��b���O-%�xw�w+>0*ma&P�缡x'^�����,��������Ѫ~ړ|W_��N�|.}���L�
�����&��Jt0x��=�u�!	����Vy�.�M���Y%�}D�ե�	z��q����p���:�i�'|)N~�v�~����|%33���ٞ:p1^(f�$�cޢ��X�ec�9�wOݝsI�5�>#KC��<w��2����Aa�R;W�Z8O��!=~��=]��Ƅo|䃨�I�(C1�w���Ir�0�ם���r;�g&�v�-��z^�O,ԉ���]���(J� �*�}yb2�ͩW�;k5)��bٽ{����{2 �sy�a5�6����8�ж�%��I��N�>ڷ���x�o����R�fw �x1Pє+��6�o����`���wJfp��~k��iA������X"9<�z�z/ܟ|�A_p ��D�^�|qE������e�w�f��0�z�0��BsV�����f*�ƭ�+�(�G�q���`�8��rc>Y�i����0�락&�{�A��D}�R�������ʈ�\1����(�x�������r*r�l�k�A��]T}ܤ�2��aAw1Ze���<H�}W,J*
'�5�l0�=XA�A��LXDp5��F�>N��L��^-<�����%��x�Ś����e�lxR+���`���#U4i��',�M�{׼D�ei�C��o*b�h��ZlJdN�u�_�]3T�}�֞�n�a�JOeޠ�r�V����_$����
Zp��V3/ּ�ZB�^�&oCB`9�f#x��&3EE�ek��0�,f4w9m��`��\5X�kGe%#0���9�c#�y�প�2��os��5]���7��)ʛ�z��c�pz�n>=�M�V��g�hx �CG:$*��/��C2رbj��{r�#�,��A:��7����+>�x��
�K�ҏ�֙7�g����d�->��\I�V�`t"���{���*��X�~�J���1�0�ic�~�K��o�2��UlC������Շ��u5V�lF�/[y����x�E�� Zo�jU3�6=8q��Zx�渷��*Ck`�'�k����AZx퀑�@�?:�Ecq_f�q���~��PP��]^�]��?xv�B	�m���;p*��I<_�r��[c�-nD7�}#�$�:�Tw����+ꆼr�{Ҕ4o���\U5��|S"��&jQb�u�w��xz�DG�^�S����!*��(X2��-,�r�,���{ә�1�3��b���U�Z\P���]L�B�
�a�5����n���ڙ*��q�i)H�w��/mS˥���]���/S��]㼻N�p��:�ׇ���x�M� .R��Db���z�m@��h����xS��d��������!���[Ӯ�}�μ�P�=OQ���ȇ������ ��i��� d�Y<����E;�S�k�ЂQ�!�[M'B�_��bPg	��j� (0x�
Ű�2�⸪���B�ta��֒VV�4�ɐ���Zlu_^����ҧD����O�z��j���NTh�V����,>�C
�d���=�8�ݱD�W�Ä1_E�XV�U`ʇ�S�Q��Q��Jǂ�ƞQ�.t<��z��|�V5H�צ
�	(J�/��`>S�C�.� c���p�={�gC�������z�|2��z���TXG�y3�i�C�W�n�=����<��3��sB�d���Q��!r�:p�*������a�����z]��+�ۚ�/5X��P�V�gʸ�l/���Co���������݁����I����g��0�kCn�R�<y
�i����H�4�������Lڢn�ѝy�|�r\+J������	;s�&U�4�]9��4��E�ޔ�{I��Ol^,M!�!�|���NwJNj�x�Ꚋ��4=y��un��kg6U��/U>ً9íd���G����ڝ��������Cԇ����+�B��1&a<���e���i����GY���-
o>��3�	�o�;���W1H=��nZ��8�N�Tz���E�����+>6�gr�+�3��M�W��??\�a�9w=����w�U�o��-0���׌��#MU8j�/}7�c{�P�������Bѳ���d��ҭpY�׼��g7�Z��}6Sl�5Z�5�NP�N��	�4s���6��ѵǄ��]�o��~��<ԓ���Ї_����B��f+��P��*�wB�!�ƍSMڧ ��3��o7��-i��ȕ®Q"�JpվU)UX2���P�:\|��Z]���>�oÝf��e=Vleae�n���-�4,>S�dj�L�jt\a�q��3�y����j:�}C���}�GA���x"�ԺW�C;��K.]�RT�Mvm?.�s�BX+�l�в|��sӱS{Y�ǝڮ+fL������HLA"&��I?nV�0��α�K�v��0��3�l�wn�cd���q� ozu�:}v��'��Sx,k�%J�lʹ�(Wp�G�9m�Sӌ����-̧}�5���Q�ݮ��wT�Q�g*��U�ށ�㊠ǮA8�F�G�K���W#�R���n�DrY�y���X'qR[�CEb�)�&�>tІ��e�Z���b���mk�N��%Jq=�� �]΢�yiWw ��˰*om�}4�ό����!�9l����غ�{"�젻X�\Z�9���]�w�[Z(jr�L˔���Z��n�MH��d��D� ;[ɋ`�;Qw�6k�>�A��v��7r.t��syK�Ȉ�C�o���k�^�Ώj@Y�go4�m�5��#x�\��:�@0��.�pR���le��m�-/� �[�ܳ�|�n%�
��Ω���y�҉�ޒ����.��o9x��	q.(Ne���Wۂ�r����v���A�dD��Y�7���<胻}��.���:	�n��gC��7��xA�b��v�0�{�������w�^ԭ۬�ELɘ�R�EiR�E^"�¨�{u����������v�r�l<��&lTt�T��A1v�Ԣ�8@Z�:;b�cJ�PU���yV�1�8�ۄ2�Y��B�e4�`�mix��Q[�DJb�T ���9׏��WH��^�_"R�y�ӈGX���1��+��ʶQP���̂Τ��٫Z*��n�0��%#J��Y.n���n
+�3"���4�ƕb��[T3�s1�0'Q��ݔhE�<�2��ޗP�|�ZK������l\�ņu)h%PI �r�n-�EyEA��i�pv1�wZ)<D(5�L���uݹNr�M�yHk��;o�E�Y�,�U��g8k�n��vg	�ߕ��_9^kn@���|�4B�w/ӝ��vWV��������R�,�5�7z���b��R��[d,�a��vI`p��u�6�4Qn�:v��SX]�5)\Y���༻�%�	)� 7
�M���@�H�v��}ڮ���-�]�^<M�&k-�=�Z�AK�>�Vi]�}o�wvs�!N%4賜;���������(��cȰQ�%eb6�-j�V���J���-,%U�j4�j֔h�DQ+
ԋ���ҰUV��V�V6ТQ-�VE���Jڪ���X[b֊��F���-kҌ��
k*�(��Vm%-��
Ԕ��miA[iiKmjDE��j�T�����ե�AJ��D��լ��R��#X�+Q�-KDb-�V�E�(�Z�P��`�2���R�A-
�EF��P-(T����Z�EV�@�[h*��Z°X���)k+clZ�� ����P��"�|��%-ùӈ���mҹ��3,��WK\о�;/�s��=���3�����S�֮t}��8�;��Ǖ�v=bu�E�p*۫�b
���0oڸ��~0�C�:�����Ѿ�E�8`�d/�m���K�ȑW�K���܂��`�2�5}��i=k�~��+w^�����`{/NH���b�����m
ba�����h{Sw2�o�$[^��_Dւ<y}�1��:���B���Vxm��d�5d���-c� P��޾'����>N��Ѓ�}��]�xAOL�{1֯wu?{�St<K��-�eS5)��8E��/�;o�)��Y�RYEc��ܦ/oH{�>﮸}t)�9��sLĴgԹO|�<򩼙�ǜs�:�ٽ+���~��2�n; x>�/Adכ�q։�?>;<�#l�:�6X��yӽ<��w^"�7}
�����
��x�+�#�ʭ���}���ƥ�vOj�hmUJ����JC����.���i��#Ww1k�����]W�u����gU�r��a�ezL��%�4ᮻ쾡Q�|�w)��͋��y�X�D��T]LeWPZ�u��s�YX��9l�3���}��'^�t�;�J]ׅs=��s��NS�'`ޫ�qW"���0�0��J�a�P`�Ptj:�T�P��VƇ�ι~��Y884TZ<��t�@�V��:��B�I����g_�w�eL�����W(yVz�P��eu^T�%i���eK^�'��|����Ot��@�߲������U���e�"�$��r����V��]T�5�LxԴ�l�fuQ��B��j�b��^�|o-�7���m��k�\0#�K�X��E�X�!�2�9���Zl���3����+AByq'ǝ:�D���{��?u�U����>��8��>�y�g�_���3�͈�㎡~�eT�an���܇>>:Q�IY'��b��������(�)W�^0���Ꙇt͝<gyi�ٽ��>v�yߟH������]3�m#���8C4���u�Wؽ+eB��E�w��Ȯǜ��arq��*}f�����Ô�1�2��kgK�Z栊��&
������GMY�:h���̫n�[}�4�l34e�}�Mnɥ��`VL�Q�7N�ە7dIs��v���g��l��p��Hc��=A, 2ts:���>y+@z3E��*9�x����[��B(q\�et5��CpW)�.��E������Qy{go9���>.덪��P�tλe:F��o���B�����S7�շ�5��,�)m�dq���.�"]�\f�b��2(t6�}�v��^o1^o�nOk�0�T+��)\o�͓�ŏ
�|i�#L�t�����]��s7��1j���{F��b[QX��\ۄ{뢩j�^P0��y~{6Qb��ό��U��)��Ü-i��9cWV�s.�c���\o��v��߻Y~����*�eR|T*�]*Vz�t�в�ւ�����w4�����8 ��lV�L���P��>���7�Y���]��y��S���v8Dt{-�L����;+����dX$Zg�W���4�S���&�M[Z��K�0��M3ׄ����v�V�ۼ(厠fIdDղ��%�CB5�m��a�u���c��&�]3!R��gP�E��O;o�"�V6H�wI��^�uNS���~B�Vٽ��V��ڙ���^�ؙ�<�q�֔N�?@м�U����c��59aw��q6�4p�G��`�Ϸ������w�c\m/3��V��qV<C]g>�V�`U�!t��
y��Z����	�-��m�� �i�.��8A�T+��|�x�t�Y��w�sm��}g#o�2���������C�O����p*��8���˽ݱ]!��b���d�̀�fa�>��U��ꝼ�G����S~U�\�Φ� ��n�Qգ��8�:�^j��|���!�|��v�ӈR��W�C�c��w'��" ��/Ƃ}{U����o���U�Ι�(ru���>�y��l�4Dw�p���4�h"�Y�Gի.��`2��ɛ�}y!�z�<�u�LgB�XY��Pc4�N���a��1c�XO��2��]^K�F}M����NZ���1�м}�"Y�jon��V����1 �~�:�-��>��,�۩��w�^�uY�w�݅��4��M�~A�k�sK�i�t�e����b�X�%f��;���џeHLv	�8PbT*V�F��P���[�ɓ�=��-��1Щ�`ES�Fy��X|�R��
��~5ٔ;�ҿT�w{7�ue��T�kC���ؘ����;�*S���[����t�$��Ѓ�v�x�|6��z����R:�/"�Ժ[�W�b�λ���:}��U�$��d�A�nU�W�i0E���6=���s��.�s�kMaW\p��=�\��3�!���IXoާZ��
�/KF\���\p�PܧPK���Ӓ&ny��Ǚ�
�Y��:Y����J�:l���Y���=]oިq�4��έ�i�.��uhU�� |ɾ��}�;bC�%�B�u]�,���ʓ�8w��3�r]U�V>S�݋��a��_���p*�2�J��L�353�y՝���֑�n=�z���a�4�TR�I��/:L:�{v\2�q�N��Ƀ�n%}��VU���Ջ�R�G�C�]I��Y�%��c�i��|�Qx��{�z:�M�z7M֞���
�,�4�k뵜@�Y��	�5&�1k;�vb�0`;>�~?:I�	p�f��>ƴ���'����*g�M���%C�ŹxGkrYb�x��]P�glhu2zpΦ%�.��kw{C�׏����/�d=K�}|�
�4Y%��\�Q+�"^���=�ւ�������By&�)	n�(.��i��x������%��4D\��,�p�e�����܃�W�^.� �{=���=�>���1.:jP��f��7��6_���i�D��Z�j����ۏ7_f��56���	������,���p_il��6� ;YV�u���1Q�/��_�0��ti��Gz��	d�����(GU0\{���5#.��`���r�6$Pܬ,�ϣv��Ӣ�e��({)�s����7���<&�4�ᾱ��U����v�Y�bh�+5iv��[f5~W�p��b㒘��g�����6V�XWT�i��Ҋ=\���(U�k<UK2��cm	y3�w�Y����1�*�����՞(G�&s�`g'�s��q�PY���ݝ�q���W�+���wXf�6�`��$��٭�}]懲��u�Fl�Y����������ـ�B���G�Ħk���Yᐠ���w�C�˼>�͆#�_�R�|(�����b���R��eÒ��n���<矯��{h��=�l㮪���G��0p�Ԥ7^�q͋ҫ�3z����>�w�nZB��㍨f|:���b���O�4&�{ٞ^��{s���<�]�w�"�f��O��h�����ϩ�],����N�M�[zB3��[:"�#F���5��`ӯk�������2���k{9�T=�T�N��7�����|PU�ܻgj�+��@����Zrc]��k�f�+¶��z�O�C�	�vx;��������^�ǲH���%vQ�p�d��ꨘ�J��%��m
�&G����*�.iR��Q�>�=�+�6�gS8H�X��b���w���K)�m�='Fҁ�S"2�^E��[G��3�_v�#�L��m����.�^��#�-��=[�;��`N�;�8�;!��h��%w�/�gy���'���:����gpܹR�͓�5�H���P��v(UD!��p������V�"d�f������n{�с����TP<eR|T*r�G�Vz��w�+���^RD�_�[3V�q�|�>^71\�1�|�Ea[��:~�v�ݪ�|{V<j���nk�%���.0ά>�Ao�,M^0��f.�Eg�-3ֽ}:���z��������tVW̠F*ί���>چT��;��t���)�׽�z�04t���^�,۸h�Ϫ�#�"`�r�Z�F��w.��=�k�]f�դx��ǽ��6�»U�X���(Ps�Ū�I���a�OY�:k���*Zb9]&A}��B����]��ӛY�s�����6��!tX{��w��O�ӅV�*�.�u������i��엋�k���K�7��(�z-vT��ϖ-;:�p��;�'L���u$(�Ji�[��Oe7q{vD���V	=/FZ���~��,x� A@��
.q���{����qL�g�M���˷ �#�nun��.r}�T] ��Q��eN^��+�l��xo�J^ٚ���l���v���*8��A|{�
��+�/�v���ac�3�����Q{S��\X0�r���^���!�GI���O�֌r��T�<76�4}�8�yw�S����B�&x�Jt��v�y���Y�vڨ����ڪ��szy7��\lz���@��>l�UZf+��
�W=;��9�2��p��=�E_u�YwD���6N�xڏ�%��!!��\_���������*p���pu�1:���ܑ*3_2b�޼��:vG���/v�
�Y�>7��R?�L�[�P��+�$���=��e)�ǌ/)�\hd�M=�[u{_ZL�S��ކ����8�V�~��kF,C�<4/��u��k�鴾/&���V2���O}|�M��s	8D�,�qdz\���4�w_=�q���"{�~4Nv�{�T���|�t��h������\2*�cD!��lߥ���3CùF�lI'=2w���P�۹����쾌=[�VP��X{�3�D͍��jJΝ�\P�Vx��ey�y�o��1y�%�2��L�h����-��{�d�U�+�
�.�1���$��������f	3��&rS�}�af��ʅ�u������y=ut��%��s2�N�A�eTʀ�Z��(m��S2�1:�Pe��ek��ד�b�ǽ���z�����C�F���k̃o�||u��G�ީ<��*��,cxS0�j��Y��; �$a��4H�m��ӳ�+s�L�s�~��0k���˗�z�ResVP��f�S$����A4(�����
4o�[�zf0K�J�,>�-uj!�VAD�7��JC>j)Awm!�xbݎ���~*%ƈA5DaӌW�?"a��x��1a٠�CZA�	O���Z�WvO)�	����G]:�:u4)��`م��WQ-y0[��6[N��fz�K#pދ�'�Ķ��[N��U7���G��C���M
1dYG�����|+&�L$֪q�R�L��Wܡ�2Wݲ��]ϋ)��;ciҠ����	��c�.�]]��)�����cq'}���*��T��H����9D��E��
�r�}�c�;�
���JI��k17�w���0yT��:�)=9�$�7kbSE]��;SC�]�ai��\,C}�,o=��[d��a�yrA>�ӊ�����壣�P^�i��F�C=��Z�l�s�l��u�`1���X���#O<�����c�pd�O�������u�r�Ot̻��D�b+�9�lbֳ˕���m��٩�y�fr*5$�r���T�4���a��a���ջ��\�enH�;�:�{��z�5��j�dn���Հ��ث]b�l�G�8�RS�X��-ǔ
Nf�R��^Sպ�c���@f>��c�ΛMTާn�ϥj�l��}Q���r��H��ar��o	 �����,��n�=ݝn;�R3��c$ݻ󓴢1��Q����d�r���la5b�KT��p�2��B#�wG4bꖸT��!�c��<8�佷Y����n*��]���
ȥ���1�(�H^��pp0e+�:��p:�Z��K*J�]+�dh�r��;i:*�Yۤ�N��AQ�7)�Z���T��{lX��ɫ�CC�he�q�Aؾ�N5&���܍��&[��:3.r��	*պ�@a?bНn�e �$Z�%��Q8�����&�g\q9k������&�җ@��:B�b�{���3J���]��b�M�,�� l!C��4N�k�ms���I�}��Iw4a��˂��MG�,���Ь���;��������=:q�3;��"r�ZoMܦ�k2����,<�� 46��� i�Z�v��u�GD�g�hr$j#�������l���Sn�ɤ�k*S�ˣ��Ra��1�`������ҭ3׺eK�@���fڗ{��#j��XpQ�쬄�|�u46��ܫ�V��ɶ�{6��b�l+{��.�2�R�N�Vؾ��q��+r9Wu��W҅1� E}@VQ���[T��*�Z�Z-����U��h)%b0KIT�щU�R����Z�mjKJ+-U��"1[k%Q�Ȗ��-�X

�Z�X���**
*�mB� �"���VEFJ�,�e�F�J�E�m�B��KJ�X�+im�*(�h�����*���U�aX(6��YF�+m*4m�R�V(���Z�Tb�Q���Ikem+(�(�1��Z [T���P�EV��СV�Zأmkm��R�����XѴ��hV��eTQD@�ڣh���E*�j�m���Z �U�**��*(�KE>��U�$�I�fm�3�a�{vogr�A�@��B�H���]��/+nJ).����trG;�y����j���2 ��z�],���Z���9��eW�V��^�Y���I�s�ר�L�B5�W�e*�]��DvW�m%<]w�[�߅k��/��N;�#�u�~z���P����p8��+8gU3��� z�OI�w&7�����ǜ0`���B�xmu׌7+_��Y�C�e�����1M�O�]F��x��6nV�|�75BM���٬�Н�cU3�+��vc����Bk�bv�j�>�AT���H��q��B���X:���`��:�_�<���K���#)�ͣ��>hZ7���XM^'�����P�O��NAu�k�זm�<`�q�k�X�x����@�_5)��2`��
��o�M� ���Q<��Byq�ϔ3�5�X:TL�d��u���}=��w3��=��T�MY�؇�6�C8���Ҕ4|��v
�׫<2�O$}0M��"B��"������o7����jy��t�]�%���r�V%�F����{���o)'�Rg��<��Il������zz𙵏���2�rx�9���S� ��m����$��nkm
i�Q:ę���C������/�>�R����ԝ����P�6*���L�F��u\��I���К���Vs"P��߾�tU]^<k�M�8�b�����X]�����lW���v�&�������(�(H�¶�������.4l��!�`ͫ/��'�������?�$��~5i����Vİ�7ʊv�S��bK�2���q�g�dTiP�Y.���U`L�
��R���pk0�Ҷ*�*�5��n�D�]�H�:C`TQfQ���.O�[#��)8��;�]��Q��L��{���ϥ*���q8&���=պg��Bw)Ԉ�GR��㲰�-7ɖ0yx�M���c���[g�:<���{��^Z��X`������Xh�:'�0�֡��؅m�����oϏ5ai�<=�h������6�4Cg�[N�J�����{�M�>ݳ��o�]ҵpS۫�_���&�J���s�N�x�|�G:��*f.$�w����P�r���� ��Q>{9µ��]i�;;��0����m�ֆ�a]�ت<Bb��4�h�l�;�gto-�O�mV:�&���B϶���K\t�(WE�9~�K�!oݳ�����5"4�]�Ő���ǳ��Ԫ�3��u�2��OE|��k�8쭘=�}FP�X<N<��:Qbi�����ؽ��7�v����q5��o2gϾCX���L��ju�,!�Jύ��gpWϫ��F[ɞއU���z+��3���Av��Urf�C�-��u��=%8a�R>Qw���8��V�,�+Z�}}lՆ�!�j����%>m���m*���\�tz��ʬ��<�.�Yǂ�z�K�g��LX��>NS�q\4UN�/S7��I�	]�XV"��ʅU�0�A0��wn	�{�/���((Y�EƊ���"Sa�"��F�=	�}������K����KN�Y���;�ɖ���� �Nj��c��H9�Ćٜ�k�-i>r�S��ȇ�N��{϶�X��u�v�P���z��}(C�N�5�V9k%=ɽ�.�W>1��Iո��l�dxl5�+L���l��<�Yρ���{TEbӅ\~�]�{�]z�ЛS�y{�Rφ�����c(\<;���f���LR�Jx��o�~�Ǯu�E�T:m����`��0��LͿ8�wՀǮ����P�bE�\���"^�;��q�e�(�J���|�,��"ϸ�y�U��0�헣�<7�έJ�,`�m��p3O�u��7�|��P���� T��
F����M����3ÅW���[�1K�50�»U���L�D�jY��]��TD2=�'y�y��owb���R���B�
S)�[\w%�8�c���W�z��@��@������܅b<+�<5�V��֏��Bg����ރ���*H)�P{z}�|��KU=>�Y�TjΖa���0�Ix��Y5�{��:w��EZ���/}�v�NI=�`8SXf�K�WuVA�ֱE��ʗA!1��j�^��6���9#�SY������^�Ņ���|�2�:f%��N+:���m�i�}{��^������G�l�v�9��g�]yfA:qp*��� �>�<Nx�����7�f�nyg	Dw�`�Y�J�<��'�گ�B%�)�p�� ��~��s����C/��	5E��<��@�9�_�J�]B^N�w�/d��o ���J�@�6�fԪ�E'b�L�Y��):�a^j���1=��{6S��d�٭F��TzpGEr��U���=t]Wt��:�����i�^(LD��FU�(aSU���"��KĲU����vlT��9�5��J�g:��Z���EʇD�,�ϧ*8m�T.;c��^��~��ۇ�P��n:����c%X<���{+۩�qFD�p)X��yo��:0���Zl���n�>
m�H�٦D������cW]�t�������g���Y����>`��)Za���8�v�/�i��qk��l�~$�+�z�e�a@�H���wr�q���K4�Oڇ`;[�Uo��n�o���l'�A>E��͉�[�n�-��x�_"Y��}��f�t�u�*�i-�<#���N+ƶ�����i�ؽ��/�d�7Q,d���f���y%��ڙ�����Qk�V�R{��3�,�ާ�`�Cm�G���V�i��*��P����uڏ��5k��4�x�͋��\j�3�m���4C�^*�,ɻ،�����Ř=ח�WU��Y��ڄ<��ͨf�Ư��6�p(TZIG�\V�{\}o��p5|����kr,��L�3_6�^7�FR���W5y�r{$���]W��qi�+HG¢��ۨmU����t4g]��#B��_�ov�����v?kC��߮�0�Ŏ��\:����+:8�
4�C�����Kѧ��u֨��@��+����+j�[U)J�~�3(��ʥG��n��Q�}��� �O���A��KW�Rt�[���*)��^^�"��2�����]�O>tG���0Q��f����V!O.�:q&����U,�"ۯsĠ��ـ�LB��3��V�TC2�C�W��F+�x��+���"bCv��n�)����B�>��)f�;��!C5+ٙ�n�NN�\v��@�H�m#W�(Ky��|ggX݄s�h;�.�F�>r��^��\c��=u�>��q>�,خ��s�T�y�,l>���y�}J�f���"�����v��׍堾�(X�ad�l�9�fVA�컶�\�)��[��yh?PǡQ�_2��Hc^7�/��=�P�y�J�B��
����&p�3n��6'��^���+�m�8"�yr�:y�Yv}�7|����2�r�0D̰׈�<���0��:��n'�H���s���u�̽��x�_��4Ж�rUgT90K���6[Ձ�ʹ�ΜP�hׁ]��;����-2�"!���r��\{}o�rw>F�z'��{��r|�Tv�8�lK���o�E��|O�]�X9;8e�\{�ɿLJt��]]�E˲`P��x���U5:�_,!�#��q�]S�����'v�@����m�߸�
]�B�V�Te�����ǃ�v��֚vZ�� �2��b9����A�מe����r~`ࣶUJ��w�R�\���j����.\X��F��nh���f�f�B�Wo[�n.�����a��V���t֯��n��W?4��Z��)t��e���+��0h�]�a���Y��{&��ɧ�D�\o��}�L�j�:��:z���xJ�LX��zᜍ�/��:;��r�&��m����*��O����ǊV���ȱ����_xo?kgADi���E_�t����I�R�5�s]߲d����wS�UB�z��u[G��pbߗ�0��,cD�\n�3<7��N��e3dT�4,9.j^�Ӟ�E��Cʾ󠮑e#aЇ�VyyT�9�9�c�!�{��T�e�=o�q��B[��9��Ayzx�x�Ճk&��tVd��w�Duh6=�X�mC�r,"����N^3��H��,�d���ږ��B�*�CV�]W��0���q�=,y`3�Hȵm���WO0���VlUq�b@��#�Ӫ߽Bc_i�|X�ެ���M�xq�u�ǚ2�ͣ%)���V�����������mw'q_)И�$���N�8�[�:��ƶ�s�&��Vz�#2��b����s�{M�"�幹���N�N���׮���6��Vq�,O����L��>,����=����yB�~/5����rn~�]�a{��<,�\xU�*���8�qȓ:�f`���fI���lg��p�WA�@�R��|~t(�8K�]�R�gy��nz/N���3%��/A��mB�1Ֆ�_c�6��q���W{ٙ7�Tw���!��;��m_ɯ��&��kVPZ���,�S�;LDP�sG�T]\�1���bv�48j.�h���������]q��������K7�z�{��A
���!	b�j*#+�eʍx�4ީvӞ��w��J�43P�j:uZp�a�KF�Q_5c����+���>�f���{���Mu�J ��4i����l+�UyV5�dq��ұQ������ώ`���S4P)Ub2�	׵�W�����O��x�AH��f�����n����K�j����v�L��A��s���m$r�w�k4/clp�����yuϋ����t������X8_^q�F��t�,�I��L�.*��i�;�x�ܘ����������_���o6�޽��Ki&9*���"�(Y�͛����*'ٮ���v{�N�$�/{�
�2W>�b��A�~���.P�=+%@�m����o{���cJ�46W��>O8s��b���;Vdɽ:�}�={T�g�����{m��g=-���":]�^�j��9���M�i
��*�Vƫ�z�o�(���F����W{�3�N^���Rl_�ъu�9u̼~J�'����Ovo_���_.�)q��UIݔ���\4N8���U,+3[R/;�F�-�ylګyػ^(j��gK�^>Z`q����sGP=�6d�<խ2��΅��k�~{y���ȝ�1�<�_S����c�w�c���_:e��+��:��F�[:n���{�K9�Y�ՙ9��/��Zd��x��jLN��ṧ�V��/>Z��:�t<�1�Nut&&��u�;W}���>�}�v^�Wځ+��8�g*肘��w�[!�m������*T�29Vp8�+9o?� M c.���p1��j�%�b�EV�(����	1IǊïe�wWu�e��&�e�'�${��[�V]�f��_mwh���رj�B����GvJni۬�≄w�-�w"�N�]�x�L�S*��ݲ�n^�I�sW�$wD���z��������bBV�S�R�ȕZ�C�|�lQ�W}�\F�܋��Z��,#�1a�%f��kt��Msw�PWn�����5Q���M.����Ս�6��"��&��b�k����7G�3�[��_Jo�
�R�w��V�R�m1Z���`�{��ї�9͈+��k�3��^ZFT�rl��h��,�k�dL�˩����v�I˅�iiP�-4�;*Y�(k��ݛM�8��Ŵz�:BCM�VL�],]�-���$)��ܧz$�@b�bq�'v:����c�d��{���}Z�z�r�j+�!ً��7��u��w]b��%���T0]=�w*�`9*���;����7:���^�<A�Qڭ�6F[�̖H��� �:��U.�V�/O�Wc�����f2�8�]X�s\$�k��*�dǚ/$}G�=z�=���t%{]�����.ܱ#c{�%���p�Ρ�w[6n��y���c��+���6�'��\e^�J�!F� �x�mf�*�#,�wli�w�P��1.�]C���u�ڵ���<G)��w�٥�k�6�4�֛Q�˨������7�j���E��O�U|���B��!��z�<aF�{��fY�u�n�9V�n'r��6$�nj�K�uhp�e�W���)[��Iqن���`��u��h��%^d�LN���pN�s\�wv�{�.@BJ���h'��.ؒ<�#��y����Wnq����(�5%5�H�-����ܵ���qt����w���Y�E��z���A��X�k��i1Z�\s��i��}����&@r�R�0���^��Qn���Ӹ��������_=ٛ94�����*�b��Ҕ�e��V�V�b�T�+ET)j�kj��"���Zq1"8�.32�Q"�[,Te��Tˌ�\iK,[[L+1D�b�`�ZYK����&1V��2�U�J5��J�ʂ�R��LXfXUfZ�.Z�&-���j���Ael�.7,�f\�9�h70��c
�#hfS����8�\L`嘙�啅V�j[i���*���9aU����ژ�U-(%��-���
ŭj�c1���CY�-)X��E�4j���U��7-b�fDem�"+�LS-H�kW,�����pQL��}޵��k�05���N���v��wO�?)���M��\穫�Տ�t79-˽VݝE�Ѻ�F��7;�Oվ�YS8�^�=*.��OU��g)�W��rg��?7�*�W�N�2�p�=V��<��q#7M�7sZv�M�n�>���h� �T���]�S��]�co�+c���vL��+�a~b�G
|e)Ĺ]ơ���k;��話³��hm�m���EH��s2Ӯ�U�����y��&}4U3|�϶�f���8g�ӨM3�~����[��E�O�D�<R{7��п5X���ք'�����kb޵���cO��ܱ=�od�2�O*��ǌ���1����r�l^/x͍�rg�oX�t�gVDe-�{��ؗ�5�wvf��R��oA����ӕM]$/�=�Wh���f����[S��SS@�=��bl�ޫ�RZ��Ⱦ�=;��	L�5W[��D����۩�a���ʷ\�^d���e$�q�����u�[+�+�ʏs3��&�
Î���S��<f���������+�N+엹O�s��`��uΞ��e-���'�|����\=s���,Z�f�K���c�Ù�մBߜ<(�6A|�5GK.����Y�?E�Ӭg�x�f���Z�J@��`����a���޷oq��[�u&Պ��Z�[���^:���r��\�8��e��h��d9�Sh��y�s'�j~�"1f�/R������PW�"�X��0U}�;l!�]�uq���gy���X��^{���5��\.�1\M��<by�ce�3�jQ��o�X�R��.?���7��{����#֘5�Rv�:eX�O<�ϻ<�;B�b^3�:��'�S�36�a�E7'��� �{VT8|O��=G4�8�~8ј�^��hT\�w��-v�[-(+�v�tOT©d�w[�&v��RX��Il���z���z���ׇ��2�k��]�t�������3WW+�s�n=un\���M��o��X�.�m�];�}�~b��]qob���~�BvO�2�Lª[w�oz��?y�����;�K�|wo�7ǞBѼ�Tg����O9�C&�P�'6w%�����5sů��͎:����"�X�u�Ы�{}dlcw���Ƕ����:�潳��B>@�����n���3��;�Wљ;G\����rnGH�z�Ju��(�x���0�#Y:�޼~��]����Xޯ���z���Ҿc��\���u���u�m�ߍ��A\�DgѲG��ؓ�t����s��@82{ݕ�v]/��U��/�UyC��<�Q�/�(Z�WVy7�l	c�ʺ�fJ����rj�A���\���b���*$nŜ���k���|�}X���G8�u��|'K�#Z��[ڡ4}	��_Ş�\��k/k���[;��xm��߱�t"�w��|+LI��u��v|�^&񹏦vw����T¹�)�U0�Vqɵ�gH�M���ŉODwG���E]��=y^t��c���}��w����g�:�!8�����N/wٰ�o��;���Zف(ƈ뢤�O�b�Ɔ�8Nރ+Ç����֎jx�9���6���E3�U�^j�=�����{b�ϓЧ��ke��4O?9ʳ7�l���%��;�Å���*���=���;��i�ٹ:c�X�G2z^.�uaߗ�����^����彳sۨc�1�v��>���lP�/��=F���F��±o��n֓�Ք����A���z+'���0U޽�:���h7�X�ƤZ��7��������s\�w�k[huHU���%v�t�K��b���)���2�ݵ��n�)�sd}Îs�)h�Y'���}��]Ek�=�u����d�!����y뿇[�V���;�I2lְ�֚vN��k�FC�f�5|�T�7��W�b�Y�'���֢'3A��h�N�gy��T�*�v�I�V?o�3=}|I���t7�	�<k��w��զ��f_��'l[��2S���X�tS@hY�^2�Ԡs����cޟO40U83����(G
�ܭ�n��eT���ޱޅE8��Gy\6�2���ܖOp[��>��^p�y�Ǘ���w����*
e�mmeDd�g��t�;�-�}x�T�;V�1��n`�������a���]:��{8x��z��VkϽ�!�g��g�>���7{��\�JY\T���Y�=ԃ.�c<�gk�����J�_P����,=��4�%Ԝ	�Qb��'RɁű%:����֞R�I�>~v�I�A���!��hѳ�@�mvw��_d��:.xڞ�����um��x�*��k]�e�N$�;WJ�V�W����T���^y1q;)Ӽ�ܯ��ku�S%���/W�����g<+��p*���<�wk�q�$�K��:�d϶L���?fJþ�gy�&���(6���=�ɂ������\���z��їQ�o_V{za^��Q��B>��@�#b��w~��ck���μ��UǇ:p]��@Mb��t<ϓw��o��~M��|��N�*�󠖲��z�7��K���޻���������u*o��\�MA�`'E�LK.X�u8�MA2�go�choMFk+��n��ݾ��f\�_�g�,�SB<�/4�r��-6b��\�ժ��f����n�5t����[m�ܲemssfl��.�"ۏ���s�u{���iN���|ćK��^���`�0F1�����JmnB}ǅ14W?VP�YQN��6�w���g��Ů7����Q�G��S�s���	�藣��71�ܗ:���bu#/�Ԏ�xk�v*W;͇���nk{���}�lK��o�S���z�C�����^����d=ͬuӽKV��:�|6緳�(�y�	����n�x+���sGO11nX�}&�c�c�<���[�,>�׭�#�ˑf��ٕ:�p�X�9���nu������w`EfN/���W#쓺-�a�����xL^��=پ��8�s]�b�jo�j1�
Thv�a��l�[8^bHe��ƴj�n�Fʱ�00�G�wY<ű���_t�Yˇk�]�'�-��At��ξ��c��31���W{���_oخ�C��c���1!}�A���Jm�Ǫ3r�}�Ӹu^������j>�Θӵ�|�틣�he:��/����o�fK�?=0[0/Or����M��p�F���\3�=��~�p��gR3�U�<��[2�X�x �x�oN��}����0LS�e�kY޳CUC5g-�t���f�B�b�	���t�Mgp�Xok�?5��R�;����h�N/�|,t&�p�a �α^��g�������7�K.Ժ��W٣�mwEF+���j*�7�r�/:�1�>���>�d����!��epZ%3;�}������ݴ�j+���Mgi�2@�:*s��L��u��<mg���d���n����/u?�xK�,���� pQ��7r��ܩ�3)&&]��{�;��";`tш�bfiFr���0�7���7/;������d��Ki������#;��W �O).��C�U
����a�ũΫ���t</nM>�w��TwҌHH������{����I�məSə۽>�����aC^.���������<j��)��`��:.Ȧyws���n������{k���[w��/�͕}.s���o�[{�5YuI\uqy�D���1z�������l���js��P���Zτ|�ad��`����~���yy�ԭ��y�с㲳zڗ��P����*S�'��v;�8�2v&���`�v�y�t�N)=]Dv��<j�4k�мb����6O5�ζ}PD8�򖵺���ᆅx���S[^��uoI�n�{fu�OYl-�깟SEgO���J]��7~�8�=�r#�ʝ�����B��F���[����ζfI�y�u���w�3����R���j�zP�ث���J:�N�eN�`��i�|�|��(={�����~dG�8��ݛ��T��~. En�Պl_�� ���0"��:V���G�aA�1Wc4������p~bㄈ/���&��qζ��%�.ؾ�kmN�Wo��Q����ƓC���Z�o��n���t��M��x�;��ǣ
b�l��V���(3$u"��).x�5X��R���eWz�y�i��N�퐨�ڣo|n\L,ֹg��oTt�/ϔY۞���^�'�o�y�|T��9��N��z=�y��jX���R���\����>��̺t[�T{�}���\B����>U��:Y��R?R��U<tn^<�9*#����P�����N����w�����j��_�*~t�UU_텠Ii���II$?��af����C���/����^�/���N���tG~m�$�0@� ���9�!קDΣ�	��>!�`�~��Bv�%���'��BI�/�����w�;������{7���<��}�FgV}�=���|P��Ϧk��{�B��`sgs���{�$!$����i�����~��� ����		$��A'�$��'�/FH��f�&�/�^U�P��9�\��x��X�@�M[�DUL� eO��ة9�3����O�)���?JC�:���I/���-��w�3���ߨ�a��u��"ys�	?��w�I!	$��ݡֲ�����@�I ��$����z j=*�k�S��}d��������wˁ�.��IUJ� ��1K���I�y��fH�Vȹ�`�� �$�E�+���'�12��)���^ 
*���Z��Kpt��jO��`[�"�h�p-��ɩbZA�k�8m(��u��r�s��0sY*�ģ�^��mUU-pc�����E���Y��};�`���������O� I!�r$!$��	�`D���V����|;������P���O���HI$<ъ���0M����>�$���I��~g��u�����+R�?����2�S�1��ק}�}�C����CS�~����D��?\��Rdk�����h�8��fr����*?0����C���a����Oڈ`���I�y����Ý9�9M	.�5��ݝ�UDUN3��C�@��д�O��G�C�?�$�$�O��<���	��9�v�T��m�Ȱ7rԔN��h$�S�Ν�d�����$��q?��惿?� ��i�9����)x����l�TETׁy8k����������!��Т~�O������S��y?�âJ���H!		$����04 �O�"֛�ET�t��B!�u��?o��w�|�O�~�����;<��"�����RO���'?T��.�p� \�]�