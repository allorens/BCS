BZh91AY&SY��`M�f߀Pyg����߰����a ���   �  }��    (|�   t    (  :    95J�U)E
(��D��p>@�2 =�TP
���<Ժnm뮯g;[�B�S�s�Ν6�ظv��ѹ�4��=������mw�p*����^���s#�;�5�7�k����a텽ݳl�(҅ �U�j�<:��h��9:]��åps�l:�v]��t賤�n��8)�=�n������0qf���f�n�w^���[y��kwnKg)f�@�7� �(�3������w\�V��wl�6�����]��ݺ�< �c����w}w��%�9̢�љ�p�69;d�{����py
(D����ݶ��.��Tۢ�M�m�ڨۉ�\��;���۽���J��#���uK��罛��Vn�x�z k*���;[�m.L���y��Yd閴�Ml�]����7s��f�K�ۡݹ4m��Jr�q��������                 
��)            ��F��JBi�L& 4d4��L��S		%QQ�& &�  dhɠ�)��������4� �hbi��ST���M4=CMd   @$ �h 4�<4I�'�z@z��@UOIjT�4`a�� &�F#�>����K*�E�	W��(�l��}��/�������C61����٘�����v�s�_���۟�����_�yG��s�(�E	!	�*��r>S��\��*�w�|�1�6?��� �9��� (&����~��a��U������_������?Qj�3��p�N0��t�bNa�'xba��,��"^����p�Ýf���l���$Nm'Rf$��O	���xf�gC{+��M��M��%l�a�1'~��g�0�IP�e$�K3xN}��k�$h��wbÜ!�;F��F�&��o���u앳y$���%�#��$���N�)����2�|���/p��/#��G�.1�腿$�2|��Y�r}���C�N�H�!�&�4J�$�J�D��C�G�a:�I�`�G�	0LHgɉ�8���f�(~J��(��dL)�ȓ���gо���t��ك�'��Д'~N|�H�ã�t���d�F��丑6�:pxA/a��pf�C��$9Ĉ�xJ/D��>JD��&����ĘYn��w��D�5�X���LN�bV�`��Dp��D���DE8P��+�4bYC��"V��"hw�KH�x��|��"n�"gĚbN'':�#0�h�$D�$D�'�l�"Z'G(~���$N�xJ��n���%�O�Ĳ��0H��������g)"o�8;!ϴ�>���t��6j��"u8e��G����B�[�"DG�:?C�l�n��Lh�P��`l�~�;��b"D�O�0�G�bt�H?.A
)Ds��,D�p�K/��ؘ��5�����zM�F�f�d;D�o�pM��tM�NƦ����6��)�J0ܜ,��'48H��X�f�4?n#r��Y�3��}��̜��ú���5��ѫ��o|w�g��Q�Gm+��R�?X�&����"#˨�gJ�Ĥ��єv�j#q��F��tΝ�?s"_�R�3ǹ��������7bq:V+��x��vg݈��$�c�b<�Dy�)	r:D�F�˗ir䡸�%����#���'j"XȈ�8k�@B�7>A�p�d6%�DE�:i�AU�DE�K���:��Ј�0���'ȋ���{���M�8O�rA�N���L�A����"mʔ'#SdO�Au:i�t���X��"�aej"<�DE��(Nq�d�#å�u(M�u���*"oMJ ��$DE�J���smK �Ȉʩ���m�����K!�O�j�"��a��Bs�K ��8i�JcQ�ȕB&�B�� �`�,�pj`��S�O��2MF�5"k�ȍ�N
�N�[&���/�N�C���>�����.���(B��o�wR��]�)3���5�6T��nG���J苕�np��J�8#]����ja�D�v��2!L�		�j�M�־���rf�1�p䐟l$>A���[>�S>����=�4=���|�p~K�;����5��!ۜ+q8'{8��(���:_�8p�$�ѩ�şgW�>�BӅ>yx�.�e�S�3�y����mG6�/h�ѱ��N^5��Z�ƺ||�[����{�J%j�;�懓g9duU�G�Q0���rt܎�V��.�|����)��5�gJ�62}I�J֪=�G2�L��v����*^RR`�S��1�3��5\�S�*%m7iI�0��X��؝����ے->5�T����Y�_u}�{�w;�ΓNg�}��-=ߚ"��N�|R)>�n<�g
����r\��Dj<�c��`��T�NF�ԅ�S|�ơ�}>u'j�r%rK�ުS�uQ��<�'��jr�Ƥ�.D�%r$'c��$�}��7ʕ#�F�oU*�����{9�o�9S��Ӛ��K��d�{�5�4��!�C�B\�j;�����R�{�0�g$�u7&�k
��Ȓ�nHp�#������I],퉎���g
�d�8�]J���U6ܻ�7������4?'D]�aedL�f��ĺ��y)��؛�V�7C�bv����"%�����"S$DY&�g�#ȉk+���D�֥|�D�O�0�H�{*�?"V���DL&��SbA��c؉�ܱ��Mu��E�DM�r"a�\�Ps�JDG"Q��
�"A��o��ԤG��d�D��l��l�B[$D{$��#�H��WM��FQ�&�Q]rRh�}6A*��H��;�������v�+�Jc"'FDD�,��qb%�g
8f���K�E�/l����N|ԭ�M$ەV'-�C��N�+W;plû�.��M܅��gG����gg�8�&��jDJ؛���Y��F��ks���A� ��f�Jj����ͤ��H��®"#م��I��K�w��N���9%�K�*�&7U��T�$L����'N3L�_t� Բȉ�"&8J�Uq����	5�uT�f�?a�A�9�Hs�������^�}�'�.ί���h��7�' ��d�%w��J��R�))�ZnVە�%t���r�y*�s��W*�M��ؗ�n�S�y;���b�I؛�UN�Sr��y)���\Y\�*�L�qܙs�;��9/��ܚ��ɩO"a�8k��nr�*����7�h�jt�N�V3�q���檪Id��n�q�����H�co�M�Y}WX����Q,=�g~�~��:�<�_᳽� ;��}1�����OJ��!E}�L��/���@�|�� \�">�:�^_���_�ur�m�nmI%�EZ���rؚ���UN��-�yتԶMZ�F�V���뫫�9�^YƇ��U����=��U��ݩ����C�c��YS/jkGy5��S�p~�o3�����׷�������-���mvs�5T���=��W�?n�qo(ҹ�������톢��E����*��84qj檵=޾�S;Z�ܻ�Ww�T��
��wT���3w�Oo�����2Ǻ�����oWv'�D����ͳm�H�Y_w;�u?3oQ�rs���Q��{�u�>MM&y��lݲ���%Q(sG�v��3�T�T�e7S�||�Q�+�J���D�z�ݣ��+uS�N���9ԒK�>��j/{����o'�'o;�s�����W/;RO��8����˖$�g����ػħ|���9�<
��\Y��vq�&98���v��ui�W����;8��޴:���u�퐧y�'���6͊�r���w�w�\�*�����rh�f�x������>�Դ����5�W�x��r4%Υ9J�ҳ���ʸ��Ö[˲/�*oyԻ�=\u;55Ϥ]�r8���oj�7���}哕$҃R�����)��8�I�s*]��ԗ�]�\7)���_}�j�O9[e�N���[ywb��Ϲ��н��Q>?�k�x���Ծ�J�m.%��*K��3����q$���b��E��W���>q5RQR$ �تӿp��>��6�o&��ʒײ�Q��uʔ�mI��Ku4��~�|����7�*�u&���:��Í!�YZǞ�;|�ވ��vr1�����W�rWֵq/sUO���y�$�≜�����ή��GbZ�*����x�I�'��_
Tm��FeGt�]�̓�����>��U�볊�)��*'2j��6���7����y$�y9~d����#�l�l/n����g9�.[�"}��Mޢ�u!�EhU����$ǰ���$����%Wv㺶�j�Gwg�n�7gYW4h����',-5+xʯ�F��U�lE�E�Ǯ��q^@���q�-ݧM/zl�ߴe[��4dEwI#�ȕ\c9�Nn���.��y�]��ݕdF�=U��:͛�nl[�^6���(�sl�X�y�L���C9�:u��)��tg�����M��rg���,x���IW5���8�$�Z"���]�}�Ù��ۍ���tr�l8�Vc.4��'�u#o�m�h�oțZ���Վ��:(���9S$'V�D�>#r9M6��N��E��h��V�i#Fn�R�~F�o8J���ݑ����}�okiȽ��[�q)������+&��k;�=��Ӛ���W^}�<"�F�Ĵ�SC���BY\�Hq����'̫/tq�1�U�gf{N��s�n!82F�q���}s��+�u��~!�pS�5���6�P<��EB�!����چ�^�\5Tj�ӟi�TQ����H��K����DJ���IΗ�G�'����ߵ��#eTq��n.iv��m�[
�����bf�b�녩���Ź�
�~�n!
����3]Z'ٶg��G1����ψ�s���6�ԝ�~�|�4=F�q&r#�2Y�r�����P�B:o4G����u��TV��'�ۧ�Z�$�iڲio�VM7�.�kG�!H7��?�oQǻ��d����M՝ӏDR<�f�)��srAMG�q"(�tn�g&�D&,j��&GK�U���ϭ5c�9xot��B�G����{��_�4EzW�>��7��O�v�'��'4��˝��|l���fօ�9M��g�H�;Ỉ�;\�l����ӳ��8G�3�mp���=
iN�N�����D�j8�(>����aj'8q#�JQ��W�,��B4;�:�x�N47MX���m�Ґ�k+J��e�Nd�q5�T��[9�.<P�Î�iv��v�?.���yu��x�¶k�y9!;��m��TV���/tbK��a�黣z^����C�p�u����=���7C��w4Z
���W���G�������E��S�+Y�.Ӯe�(�������)?3�"��S��t��'��8���Y����]ŝ���tYǷM����p㦷���8��~Ez^�Lq��+����9>��B9���:=ya���6�[ �9�.�]#Ep��9!k4q�o��F��rdTu���#�^M_B�������s���F�W���;J"E����(p|����kd�'&o�SN:_�g	���-��~�;s�ߙ��ybe���.Ѷ>�6�М��IV/s"Ϲ��T�,��CΔ��Y�B�q�������U������˹�5o9�G�݆��$���s?ty9�O��/�<��FW�)n��q/.o����o������,�l�~��uӭ�`���y��kA��R_i*7����wi�s+4��R��>����z7zt�� �q�Დh���}ө`�����e|���s�:���߻�(p*�������D7�8o�����+�?x�e�?o�ol�Q8�g$ȇ!k�*A$����Q��Պ�����CG9G(��7F��.�Y�Z��dS7E�V�A�N̻ê��E?up��ԔR̽���Қ����7��ߵ������V���}˩'Ի��W-���M5�eJ5G�Nq�R�$�����~S����
�?�5�$����>����L��K�7�/���o��v��9���r՚Ō��V��a#�o=�Wc�%d���Qp�ꫵz�r�ݖǓ���'��['94���,�Y$$�p/I��HK(����'Z[�rB��*K>������g�����v։	/v䐄�`,q���ٳX�[�MY�7��Z�0h�4�	`�`��ɈBF>������^�_	��8]�Hǈ����%�ok��RW�W#�,4�&�qfǨZ�#��m�K5�B�dPן>���N k������'8�����}^��>��{��w���A������h�7Y:�6��f��n$!%�D��/,'�y��]Ehi4���Xqn��NȾ��~Ҋc�yRz����bG4�K�D�3V_z�G���I		hU�|��o��[�O��>]���3�^��E�p����J���k%��ZN	��/��D�X�e��c$-��m��\p��8ܥ.���].YWf�X]����lq׻����ݬv5	�̪Yf�nkZ���l�jKd���d�udߟ8nƥ�j�R�U�F��岩[��b"��HG#J�*+r�-�͖��ݖ�t��KYX�,k��(���'X�����1�H����U9Uej:��)m��XCY6l�HJZ��]ݖ��Mj�=M$%%���l���R��K^G	��Q�*B�U)U����I��wMJkscs�g�םZ��n�",ku����ux����ƨȤ�))�>T6�J�Q�jl��1Y��[���b�d��[-�dTN!�[v�µRrIEH2�3�����8�I��R��Z,��$5�Y�:�ؒ�[C[S����7��>1l�)X�w���l��!��LHT�5%$��8�M	X*�+N���,,njH�uQ����ջ�9v\�cTCQul�M�6�l�ک�ź����h܄s"R��W��e�3UN')!+�lVWc�c�����H�dcq���WJ8��ڶҋI/R�d�#m"B�A�"��VYW]�5bkk���/FEQ�	�$ƣ��d�IEe����X��X��gn��K�[^{7a%�כ7,�R�>��k�D�I	f��v'��tUD�m,�F���u��J�'U��^�X���JUSkm��%mcv��Y]l��ejèݯbJ��)]����~�G��9�d]�4��!Q��3��8ܒ,�[E�����.�jD��T�\N<�k�t�I��]���Aݕ����V[������/AX�"P��#���[n�T�����I
�MYm�K'Xծ$�C[8<��9`���6�+ʒ�H'�;;+{ʇkI8H��(�Tnص�ئ��I�n̎��\٦�6����$��Ĭ���jш�%�V\ٹ��*]q��g{w�"%�qZ�ՠE7e�R��1�Dl����WW9ا	ܕ5	Yv�U&�:j���;�����3?����zከ �2vN���A���6����?[�}�?���o�?�����_��QZ���F�~���������iU^+�U^�*��t��Ҫڮ�t��Uv�ګ�VեU���J��]*��Uz���]*�Ux���ZV��]*��iUU�*���UW��\b�ե��>��|���X;,�C͝p��1�����R,5����!�*�Ҫ�UUUUU\b��WJ��]*��t��Ҫڮ�V�v����iiU�UU�ҪڮեU\��R�������UU�UUTUUTUUTO�B��-��n-�A�֛4��0������u�5lՀU>�}��E}��oT�W*�⴪�U�U{*�8������1UUQUU�*��iUU�*���Ux���Uz���:�UҪ���X���Ҫ�UҪ�WJ��iU^�J��5����+9J�@d�������K���+��{�������U�Wj���UmWJ�Ŋ���Jڮ+J��UUUUb��"��V�]���UUb������S���[U[Uڪ�WJ��]*��t��U��a�>�e�ā��I�ڳ� V�Se1@�ۖM������[j͞V�L�Y����l囓
�g-������O�{~׺EP�������ʯ�� �������~c�,��N�(��Ή�8&0L�""aӂYD�b'DM� ��B&	L�X�blІ� �DK0N ��"%���,�`�4lM�dЉ��ДA8FO�� ��X�"&�ģ�!��х:p�"%���'
D�6��&�'Kͅ � �$4&�	�>�z���pS�%�<�5��6Z�nղ�b��J�%�Ѱ�!y�!v1-tY���嬖EmI;J��1����	q�^Z�D���FV;J�,����si��F�d��fț;Gq��a˖%�H�&����Բ��4n��W!V�+U�4Ui)eHN�WIP�U
U��6��	��:��IAb(���F���w!���Y�d��$�̶�i�҃��QĬ����`���!LcL�ٚi�e!�")�̥b�וm���9��e$c��]T�"�r��(B���	B�B���DA���YȚ����4�0��m�)k��eb�b���H��M�h��oAVgC��+r%�\�8�1[Z����R�v��-��TӑY,q�8B[�V�$�d"#iTխ����̑�k��IGlr	�D��-Tb�H���;Ej���+ve���IB"�I[���n:����cc#�mR��:��)YU�����c���H[�R��H�D+��v�	�H���$��lU���)o+0Fl%�Ij�X���Gi�{�������wwv�����ǽ�{���U[����}�=�{�������ݯ���������yQUn���}��}��Μ:t�M-kq�m�8����U�����h�G� �MI$A%ki�[P�,yM5`����+T��A�Lv�2�\��1�<ZnB�2�όAwTZE��l���Jqfm�j�GK4����M��D���C�vw$���՛��R�X��j�n��>?�����4��(��څm#f��%τ�A�X�ϋI$^�B\�i�,T��%�A�pCC��)&U�`6Z0'yd6hîT%d,����.)m�zݔ��iSͯh4�W�[���Ӈ�p�&862��̌���.
4��,2�Ŷ��[�q��p��L��L�I$��>�6D����U$h���R�J��nt(�(uw�\pe�iOuqǌ�;�i�6���i�=�B����e��H�"$*W,�+U!�$�{��O��� ����w&	s-��c��๗J:vB�y�1&�tfn}2�������:&C�	�}.I$���"՞�_eљ�~�d0�$SQ��_���p�OM3�!�>2�$�~�V�b�BA	�����*��KN��aX����F���T�����Ә��I�:jk�0���
$�d�*�8C��#�ĺaWC��7�=cKe�m��u�\u�\8�8Aq	G8�I#ᜥ^�dmF�$!�����R7)�~AÞ�d�`D��bU�2K�$̏�����:�Bg�{��p�0�72��S%6l�.D�n�X"K��DLIq��FF�d�g���>+���+�Zxvۄ�xiӃ��H�Q�p���S!2"�>#�[n:��ӎ-�\u�\8�:p���m!����*�Y25��5�3x��n�Fԭ�+�%.$�TK5��H{j�l����H�օiR���Rx���qr��$xȈ:��*��m�&��GJ,uV!W,�IV��Hu����H���� �����U���$�v�C�C����4�$$�E��q�c!Kvu��K�@�y�1�IJ$�LsЅ��ƒ4�%��`l�����N�6:�˜>N����)�%b�e�l�HH(㙽g�ϼ䘩�Y>����Y�0L�a���tk	��IB�X�S�+�I1y�ì�z�{�S0�U]�F�@�z8rg�%���,�T��;3����%���4Y�s�܅g�h�JtSY��F��|��<ˈy8�v�	�À飣�˱٧w4X-2HB!��0��q���4���i�q�m�8��ʩ<��I�t��	*T��xpf�cNN���HA����b�%�nդ����y[N�թW�:�j��&������`ᶲnY��:˺��-X�c��6ݣ)�/+�b�cq�4��x��[�q�m����:p��!��6����I$���[�
�6l,�dّ��]�Y���&�
�Q����ܡ�6R�,�Ud�1$\ߌ�Km11��$߸Ig�����ƌ�b�	1�h��v���EQU�E4�n�L�n:a�a��bTL�hٳf�4۫q�m�8��˯�Oy�%
��oOb�����q]���#c��qFL�MȎ[D!��(���.8'K��K)�ō�r(R��P���6!�,�
)U7E���U?$�I	ʵڤr��ȡ)
��T�`�C�ŉ�p�{;�̇����K�O:L.�D����$(�^I#�۱��Ԭ\3���Y۩bK��6�v�2���r���m<4ذ�L�v	s���v3(XA ��ƬP��&	f����s��2�ܚ08!�����6lp���i�q�m�8���.�SU���h���jI$�Bbgg�c����$�B	EibB���tX�$���K'�\��l18gJ}�;��bkB�w=G��!��N�i�_:����	�U$!��D�j��1\�\��������Dp���p�3�K�{�h�c�g�%ci�z�LZ��5���i��1��e�|�qO��ͫ�����I�(�x�x�<R~
I���4�'��*�>O�U����VVҒ��Z2�Zx����J��[��jZmjţrZ�N&-<L�jx�%��ӹ���Z[jZZ[���Ii�֬�V�Җ���U�˩O>�����M�D�����3$���'����Z��1ii��%���д�4����FSn�h��2���Rt�Jm�x�KK]I����֭3R�R�il��R�̵Z8��өin�nT�Z���3%�.����z���LZD�11�m��O�X�j�	�u����,s��7��O��nP�i�ĉ��8���՝����çO����3�)����'�}�?&�Ȕ��)���K���q6_�ʪ�^�=|o�m�P�f�\�ߑQU�����W�}��T���y��Uw��k��=�Oz��{�|{��{�������{=�>����������l�g<p���	�tO"CF6khQ	�UTUQ��9 �D8d���sm����ab
h�Q!8�l�:`��4D� �	������D��D���7�çv�(M.lOS7U�1X f�+ک/{ё�^��R��/�H����nݤ�r��盶C$'��Z���L��.��[M-� �g�^�)�USUg�)L$!v��bjW���̯#hSǘ�a��b�$��Y��L<l����mƜYn��2���J޼�L�UUQ�!	���AG$��_ J�,��D��_8i]1�I78X�
jIZ���B�Yt�p�� ��J.�6�@�d�`���GSlC&3���H�Le��ã*a�^!�N�ۥ�8���.=i^��EL��5wip��獖0r�h��D�v���pI	�vn�Zni�M�޸�A�N�w�IL8F<b: y���Ll���<�P `�h���|�Kun:㭺�n��2��T�oe�>�����E6�kJSe�nʚ��2)����W��b��J�md�B�/��"�q�F<eX�%�����TB<,c)�ڨ�r�DM�V%�.�I���$!���M�������0�PDLCME*X������+�Y�` e�l6(�	BS �a�ő�9$���쁛�"�<l	b!�ΊխV-t��F��H��41\%.Ha�_�tQ����#��4pD������b(u��'��R$��s1�}��[&��P�:�q�00�̂��G�!��y��)�LF~4'�(!���<�:�JiY�Q��+g�`т�2ukq�m�-�8�o1�����MUUQ0&C! nCf��S�����6��(` ^�(b�har0�Ԅas�# Ly�'l�i�i���Y��[�	��߅Z���=>��u�ޔ�[�L��&�t��ⱁ�Y�@~ņr�=�_V��Ĳ����
m��7����&��Ue�\�����#Ǩ��,/[�X �`Ē%����l�z�l.n)v!�A�RB�d)�s0���i%`zžq��|��|㮺t��x�|3�:S��?_ʠ��Q-�y�Q%�����j����A��v�Ų�@�En@��
��FB�H0ևj�-�*S>Ğ���8�0�1�7�xC�b�ޔP�G��xD��R��e��de�g��pqƛzѢ	�%�7`�<�aA�!E�c�P����<�<�(����<�w\;L�#�7So�8��4D4�Ʉ�]�.8"#���L/�Զh��׻�|9(�i� �G��<x�>N�<㮺ۮq�m���ɄDLI-Z"�,�-��Uu��j�HI��2��N��UUD2�M$p<�Fw���p�z6��%@�QH> z�+�Y�E��Ճ3���k얡��Қ���&ZXXX��v�%����71x�R�`���`��(ݠ�ր���M��.�r0: 7?��^�fu`@��na|plKP�a�(\��`p�:6@��0�I2��IOX�1�=G����E��R�U��RA�� q� ����z�a�h9`���ˍ0�ґ��I%�-���ޭ�8ӎ��]u�\8��x�JO�^�?�GO�v�&��a���Q4�s�)�JA�KV�h�)35m���(:rF�6T<�d�s���"HN����(����(�dvu�ݴI�	����j^�[m��K��ZT;b!(��
W�U%Q`��!�O�"w�������Z�����$6T�X�a
c� �)�c@d�:��%!-��	$��Z��B��WFX8�.1��Z ��h|��1�@�q���P�U꾰�, �"����$6�*.@��>�KbйbX��w)�2�����A�f���eR��ꕹ�P< �c&
�IX��M:��|ӎ��]u�\8���o1�:�O+ǘ��|O7�UU3���0�3ㇹІ$(��$�g��X�Zh�9�؃�� J�!��p6�<0(�h Pm�4�)��.$d�p�!X�ؘc�R93�B�ϩ�A]��)��Ѵ�%7,�6����Y� �Ƈ$W'�!�UJe�!�9: u�z��tp��8BgZ���.sl��|&6�bc8�]mպӫ|㮺ۮqjq��-��UUUUQ@t #v,hik�.HI��l�sr�������`����4XN���CeQ4]���t;R@������}{r&!E\�!!Pn�7u���^#U*�27�-���S�8�/�^K�L��cH�i(���X� \`bnp���w�֞6��
����RU	$n� H!4Xb&�0l�֜un:뭺���x�8;8�5�`�,Ő� qH�ؐ��䐭��9���Kvy׊�� i��M ��"ѐ`�0R�&ؘc,F`��)�����>�yg�]a�4�
�nݲkbJ�bֽ���F��# �ya��Ht�.BB��	��)��.�;���9&YX�&#��d?*�$�\̆C��p(�)�����1 �DpB�R�r��M�M��$��d�0�9�E0Z-iĘ�s�\y������/]E��>V:�M�8�O�6�+E�WQũoU�[�[�ŧR֧S�iժӫS��������[6�ҭ���Z��D���~)��|�OjW��>mO��uju4�b�V�=��=KOSĴ�1Id�Uioͥ���N�N�J�t�
��K+��x��Z\�����R�zʖ�x��Z�%�)i�&-�b�J��*�$�#�"-�$Ɩ���R��&��KCn=ei�x���)ژ⸖��e��R�ŪӨ��̥^$�Z[+̵[J���Դu--�-�4�i�)iȼI/iMIj��-"ZDi1�RZ-<E�0��#t�ϛ�^E�:��Rq��J�8嬚Ғ%�R!�ݚD�IT���$-��4��b�X%jhN;l-��FYQ#o��oe�`����rK�b�uS�
>g��Ԓ��m�#��j��㴔�4��N�Pm�*)baT�� 8ֻ����M�Q�����R��B�F�	\(�[]��p��_>�5����@�%M!���G����-E�R���tC�^W���<�=l7�!t�e��� ��p��dTK�!t��	L�*I�y#E�Z#5�4&�t�a�uU�6nQ����A�M�zD�p�'q��O�ZiH+��/G�XݚR�"��y�3�7K�����Tkf?nZ���X4j�ȜޛK�84q��������IM���dj�b���{�y���/4���"�j	��O�~$r7�U앚�Kbi�J��UX�2�n,�"��륭�۰�w&��2Fn�Q�jͥU�l�,n��8��o#����&'(��㤒�[UJ+�ىf����&�)�dMl�"R�X����C���%����eڎ�JVe�m��V�G������R;B�O�%���o�2�C#�BFK��dm�2�"�Ǿ4tJh�-VƩ$�{�n~��� ���}����|�����{����{�����8��{��������{��{��Ջ�{�{߽߽�z��{�z�Wܻ������p��<t�����<<#�����C�lw-��.ڐ\v"���n�j�D�R�8*1��HA�A�j�1R�KB���w�U�SGb�uv7n�m(�pC��;)M5u��i�Ո吜�i�1�-�e�cXV�7�"��&g��s!ኆ��Ud�O��!��1��"P�C��X��#xA��*�e���!�Xe4=KF��$�q�`�%�X&\!N	!���j�C`2@p�Ѣ��� �RBˈP����.w��!4�L@q��)�H��BA��J�(.g�b�L˃�n%�/�DI	��7: X,�@�A�ƗP<�� �m�	O�(���|ێ��]u�\8�6��4v9�.{�UUR33��i3������, P�|SOV %�F0�j<�S��
&mŇLS�H@2A�E�%+��B�i���A#���v��n4��m����,;y�؁b̨�,h�Q�mX���Y���G � t�47?"��3	���A�c�e0�=S��IXWrċ�T�p���ٲ a<\���:ۮ�ź�n�q�mm��$��t���RL��UU ����2d6ovŜ�1$l3eri�A��%�S8(s�ʪ�q:��< !��HTK�I����&!5���!���8LB��,�G�&И�`�mnM�(��N�&�!�eɟRP1�e�nu�C�	fB4a�rᠣ*�s�ZM�M�8��B=�c�UH<�71#��8@��n�>������*HIf�zH�؅�6X�Ӎ>m�Ϝ[���F���{$N��UUHd�n�F4���N�� �r	���%��������%�c&pw#A�3V�śf���օijQdE3�0���O �C��m�C��hM�ѹV��)$4:L���o���\:�0vY��q�8���b�oF
#Q����1!���Ir�Lbb0����ێ��;v��Z�p�e��6��� Ӑ����X=�PEЭ�`s�ԕV��`�Crl�:��d}�z����9�� ��f[|�[[��[���F����Ʀ����6E�+t�6WJ�r�u,b�=�8W��#�:Ʈ��ː�aH�!�S �Z5G�juFB��$ZR�ו�\�e���MԳ)���W	Ih���88��-�L�E�b����%d-�u65J2�Rm��Y|�*��7���aG�:���d��G�M<[��t�3�h8�u�t4@�����,�Z�b�:�����]8j�>0a���Q	
���%`{]:�<сS%�d���qƇ��}ɲ�{J/b�(�S$i�؀��b���$��T���zr%`�	�LO%1��c(MKZe�ƒA��H:;
G\���4W=�Xh��dz`�¬�n�tǨA��Z�	
j��ln��p�K<ۭ��έ�[uÎ#km��p�N�����d�L�<'�DS��UBSv��HK)�%wK��8����7�r�h������<n� D��Y��XsM��,�J.�r7ha��{$��	P��F�K�3w�Nrd��Kؐ�P�&�E.1� �?�3���s��պ���M��A(~�J
�#L�K�]��.@���v�(��p��c��<`��;u�[�������׆�ꪪ����s�{�>�~�U�3���������M\LY�K����H�3M�� V	!P8�C��̦nfb!��儲�E!H�):����2hl���L��i��v��p�|Q@^;�t������U6v)HhcI��$f�`��
��h:I"H��l�����6((�K��r`l>֫@�ч$0rFF)��:7.6x����:���\8�6�+O���I��UUHf~�&|9�D9h�s�X��t�s���M.BR���"��V�nY8
����nq�w�trh���cC�dՇ����*f�#���q�Ɋc�JA����2űܱc�T.�J�қ�P]�S�
0��P`��p�aҥF��x)c{�Á�U�Xx��_�����q�ͺ��V���8��!庹Zm�$�Ē"iWZ�Uwb��$6��k-��Z���EQ���"B���!.\�]�D1�J��I׆��N
�n�h���E�&����IRH�Z-uJ���L��k1�ʪ�@�I/�u�i)T�Qf�Ca�$��p;2h�)nA�1��dճ$����gDv���Y(+2HB�mL��Tޒ����q��$dd�a��#?�����Y�arƐ�Oԙ���̅�>�_���i�s�!DQ���hɦ��m.�]���k��;.��;xd)�ۀ�ݼ<T�H�[q�O�����Z�Z���<xGN�yVk.��*�[��T�-I�y�-xp�2?*���?
�wo���;��E*U���L�zg8d!�s�$�~��O�lrNQR��:p䥱�M�>�^iІoD!%H�t��1=�������J1c7]������O94�
5	
rx�J(�U�𠁞�������8v=,Nc�	����H�Z<�S��h�6�#�S���i��KuV�E�S�U�)թժӫWS��x�D���+U���KKE�R����,��i�ZZz���qV�$t�\��h�O��<Q�8'��`�/R)>H�KZ��ij���ZfөoUH��ii����[6��KK�����Y'��|pvO�&�o�4����[5&*�%���Ո�H�H���)I%'�|�Gɴ�&��6��V���h�U'R8�%�Rיj���igj[L�ZI-V��[6�ҭ-8�\��h�T�%4�i&R�$�1K�D^$��Y8��-"=G��KE������OC�+��w����߯�]ezkP�0�{_�[����CWWS�������j0h:��������_��l��9�~�z�T��w���|�U��~ ��?O�����~�U�r�����W��{�U�}�]߽�yt��V��r���{�t��V��׾�w�ƞ�i���ַV�����͟*����tM���H�2&���6l���7�Ca��!�g2�e����4���9FE&B�T\��8�J�K �(�H����6��1��!&���\��Ѽ<���3$�aʷ(�\c�"\3�2���UQɱ���r'�����:"~���OaΊuf���UUHd3�3>����vd:�p|�7��X�Z��Y�͹f�est��A���V�~�L�.0v9�'���+��
�9+ҭkZ��㱇9a�;r:���m8C��۲Ʈx�f����/��������M480�`�&d�x��o�pžx���u�Zmվuk[kp��L���Ϋ9��]dz	T���`q�KMV���D6<l��6lq<�(��Pj8,�'�r���r�7���KF�#Hq�J!L�i��t4ܥ��^�,D���s���k���!F�+#$M)D�vJ�ev��#U\Ѫ���˪���UT^�Ͷ�j@��QړMm���(�5�[Sw��6��Xt&39�+��,T)��72̄$l:�R0�����nd64Txttl���b��[izCI�|�0a�273��x7<��k�~��M�{(ZI��D��j�Mn�R����ckq3����~�=���D�t�Ȑ8A��&�ERlhp0\�gϛ|����n-Ӯ�m2Jb�󊪪@��~����y�	<=�<��X(h|��"�B)C�ɐ��4V���6�Ms$�xǣ�R�#Ȑ<=�0@ޏx���
���B)Y:��D�&7di�$*ЂA�JN���<�		4�g$�"zõU;0�Ɛ���2��0��rA#	�.nv��V�kun:��źu�q�[Ư�'�52��2�ƨ�����f�ج��7�UU!��9� I�fSs��ZB�7��4��P�rq����F3W�'�8pB7��#&E��8KEB�E�R�VY�AX"V��	D�+��t9�����354�ǟ-K��]�!�4����!pΤ#	���'���;
a��P�,B�Vf.q��O],`�ǌ�6mŭŭkqn�ui�p�h�&��UUć�S��|%���;3��HC��!�x�����D-��߫;"��I#p��\a
8��i��4�X2]$($2�Y��g��8��4�!!ۚ�j��ܰ!YK%>��B8���L��!
!L�|jtt!D3ѳc���r����ǌj-���q"��RTR��-�1��bJ��,�8d8,4�+��X�����[N-��[�x��"C.�jW�ַ�!����������݌F�yv�q�q$>r�.j �"��B"v��!X�b�:R%G",	q�IiTq�U�B�W]���\J�%-���i����Q.7S��R$�wy򪫉��-��͹���
�6����l��SUI[n�&X#D�E��Н��1��J��af�! t�\�e:8y���7�ŏb(��-L�-�$!���B��km�cD��y/���E�4��|<nB��Ξ�����,C����`~8u�b$?sûj���qnҡUTIi���9��#p��u}LԬDO'�/6뭲�-�V�V��źu�q�]a^SL3:�����S��=3�������=�<R:��k���l�/ǌu��a)��dħهY;/�8�2y�a��Ƥ�K8�۞��J�om���x�x<EWy��3�W��\JjP��k�$6$6#>:3ņň<B�-ttQ �C��b��#�aO�cX�S����R���-�[�Z���:�8�.�9��! �������A�0����G�Q�FXT�[���U�E��������T��X�B��)r{3rƔ�2�����.�R�<U�\RL!%e)^Jx�֜q�a~ɗ��#�^1��e'ST�Kە+׈��cn�Ƃ��HǋN	$xӆNj_�LދN��.��D6<)���w^�co�ׯ�N��[k|�:��n8q�m�+ư\9yĞ<�扄�0�c���I���lKP�]�7_}�UUćW�z�#'�G�GbR3��;	�q���66z��o(���F���F	Z��#X.Z'�N�L�vtQ!	��{2�2�I�1�HHD��*��6Dgɖ2ꐢU��ӲVD��X��u��&�P2!�k�M�}y�ȱ��u�<3�!L>Ot�>�7��q����a��S�Ɠ����q6�&6�c�S���cKu�V���D���+	���+DO�+�RM��d�ZZfҭ-�ZZ�i��-"Z-J����-KKE��%��S��-X�Ԗ��SԴz�%�V)--Kf�ũin*֮�U�Rު���*��~�V�ij��:�GV�-XԖ�V�Q�ղ�����Q����?�g�r��?I���E$G��D��E�kW���-6�B�Ĵ��SԴ�����z�ZGU��3�J�����U��oUIx�יjej��J�Ԗ�]In��+RZ��S)dY��"�"��ԉi�G��2�\�+�YG��Y����u��N���j]����6qs�.sEwj\�ֻ��C�ժ��b\�5��8
.�qm�k4���lDWT�����Lrݘ����W/�q��]���QN.R��l9�B,���}�ܶNu������J�&'�J֞K�{�t��[o�_<q�}&�ݛ����}��T�����K}G�~�w���D�6/��$W)�~�*��E�D���̓�H�I&=��A�(��L�6��IV��$�!NiMŤ{�����V��7h��O��,����+C*cXV�2[!#���[	^Qі�6�(�!�dB�g3�r�{<���y�$�՛���ߩ:�Xo��蠊6|�Ƀֳ-�,�9��g6\�ٽ������)��~��}�I�/��:��9��i�"������m�D���Rn'�G�D����e��p���E#P�cI�,m�8��͜)P�i6n��A-�,��CM���𻛋{�u�ĸCt�.n�LCy/���Ī�#��j��o>O�=����(�g������$���kmW���i9g,�g4�������w���ھ������D�ݻ�4���[�'�?��=�&��趮�Jr��)�bP����Kݽ��_>"�%�I%u6h�ٻ��$ڤ��e�m"�"�4�MMh��QD����X��ݖ��*N��f��h�q(��U��� �c��$JB-�k9�����K����;k,�+e���D�D6D5&��o6)��!-|[j�l��շ'Q�c�;�B��ú�"�Q��%Q"OTMK��lE)S�̕F:�M&I*�mMj�;��}���|�[�.�����J��i[�.�����ګjҷ~��{����U�]-߹w�h�ƚim�kukZ�p���T�q¤���7cf�F���[MȡfLc�QƂ��AY-�E)n5%.RЂR�:��Ki[
Xĭ �L��(�C%��e	,J��B�Y7uX�V컭��U��]�6�6j����n��m��$9�c�$�fڶ��h�Z6�"�p·?a<f\�*��X��<I^��9�X�ػE�m�t��	D5�K0���6.B��a���$#=t���J�9� �0BzS277�L��s�Y���q�����m��V��Hm�!x)`����%�Aq曗:w4�!7?�3i��迉�{)O�?:�ukZ�p���^��[�VsY�|UUq!��`���Ą!����Td�&N��I4]��'��nxl�ٳrX���d�B�|6!AD6
��v��t�!��$��(�l�(��F���X%b�BC3s�:J$�!�����:�66�.8(�	
,Q
Qv�1��k��mO�z�qkukun�Hox�����ζ�m�b:чm����I.`nQ���!gM�+^�TF.�@.܏W��e�N4X���7�ܵ��kf�b+�\��a�u�!c�rIP�w:{�S�({G�B�,��y�E�8s<@H�jPܔ��4��(�t�%5%`��-Eǣr��DrAGp����nx�>�6ǭ���έ�o��V�㇇�;9��ʹ�U\H�>�OaƛHy�>a܅�3Q�΁�`�{�\�X%��DF��ĭv���l�xx�̑���(������e�!�d#�:<��.[�#�P����4��9"3��1V$�X�=#�R�&�\�,F���pLc�_-�m��uk~><x<xGN�ߝrY[WmW,�=�0�I�M���R�VBh�5�+1zA-+�t}ݚ�$v�#��F����y�t�b�6Z��R�rQ)ժ�R�F��,DKW{�ٓj��H�W�UU\DJM���IY��E!Q2���V��6IeM66�-�J�c�4GL(�xRp�0���0BY�[}�by�$4�qu[�|�O\ї�T�r�E�u��*3��B3�.��K�(�g�Ns�m1��$��@�C���0��cM̆x���]�U���#ks]����,���l���y&H����E#��ar�SǯSx��-Ŷ���ַ\p��L�ʘ�F*UyZ�U\HpO12���:4�>d3޻�TڭuC#���Cb�X�c�L7!#s��<�.X�������n�Sr5�����?>�GK��ʳ�gi��(��L�!��>o�f�$`�5,�+$�٣H)�Rԧ���ٔh�B!��n;u,Jڪ�C���\l�M��)�LZbE1�㮭�\[��[庵��8�6�=��z�UUUUb��9�b<�ĒqԔ��Q��b��x)�L��1�$|枽DGv�3�D�7���Nc!H��EfQ	檨�U�I�����8hϻ�H1��e�h�	4ౌ@�|���"��a�	f����f�B4a(��������ݏ�ix;c�+m'_<m��N:�ַV�\p�<<!�Ѿټ��{UUq!9����73��A�!`�#��z&!���E�M��m�[,ق�L4u��o�[�K��)��B��@����rǊ,Bh��Zn\h���7M%��R�̰�6m���r�G�c;�䉹?D�����4P��(}��}�%ǆ�[��u��|�V�\qÎ#m;�Ƹ���R!��cK�~�NpI����C�$R��H�"A��C��tbt.R�۹K6iHE�Wn��$r�2��-f����R���jk]%�"J���ʪ�$8iβ�)XX!F��tt�$�*�,�9c�0c�e�t��]��<�b����"J���p.�R���T�>1��yJ}�'&%SY�B)���̉��D/��5�<y�:��-�X����}>�\B�9�@H{��w�Ɋ]�a��66E\H�1
�m�|~ĳ����C.�%�n'���<`�����[u��Z�q�8���TY��ڢ6}�.!G��4�m���j��V��-Go]N��UUć	���1;�B��: \.SLe�f��8Y�w�т�F���Ie
O�$w`���)D���nL�,8#N��u%�B��B5͌Ҍ�M���$�F���&�<�r�)�	%�fz���7��<[�e�.
zD^Ӵz�H��ƞ�D��d;[�_=[�����0�0L�æ6!�4"'"tЂ$4%�b"a�0L,D�4&�١4ADM��N�D�"lDN�&	�,M��Bi����bhJ'$�>C�� �"tМ���0��6x��a��<x�㧄�䈚H�bP��""a�ĳe � � ��dM�����]����+���Ɖ��6�)��y�q���|��|.s}~�)��g~��xs���^���,�|RG>Y<}%<O��hy�Ͼ>�t�����z�/?�K��I����_�����I~��&�m�����z{�|ݝ��Χ��_Nu��l���=��qqqr4/7ě}��8�.>{�:���%�����M���M�/���Yc���R����aw�_o=�ߊ����ϛU����~���yګj�[��߽�{����{ͪ�n��~���{ͪ�WKw~���l�e�t��<'��n9�'�O�{�ꪪ���#lZ�ͳ�*�x�Hq��!��4�c���o-�TTӳ�h���і��4=s��Dx���Ǫ�)%(��M�]!Gt�(僑Q�m#�0���A��Y���*J���HY!��!����7RU��P���$�!`�c�wͽ�!E�@����\��2d���8t�<'L0�Qӟ]���q.��UJ�$=Ό���W̧a� �
C�ہ̹�>�󜟝$m)e�r%e�:Ȓ�SiJ�U�gN�gGH��Y0\Ӣ�RG�����%^C�y�eu�����gj�bp윕��l�sϊ8�`|Ɲ+�������Z�d�Y��.]!�lwq G!�φ���dbG��kmX����[n-�N�kuk>8x��ӄ�xċ�袪�*Վ�v�D�XkUil�z��ZB�4)
XQ���5��oqܴeqe�+���87a.@���֨���M��v�r�J�b �JĒF2E*V��"�nD��&285h�LP�s�UUĆ���khT���ZF��RUB����t1с�kny��b��I��r�3gH.�j��0Co���Jd�W�5��D���ی|�`\v��
#�X�hر
i(wDa$�D e�ѽ��fg��S���B�/��:cj�ђms�QFF�9��>���F`.C$ �����1�#*���&����V����ӎ8�)���*PI"w׊��$<�)L�Ͻ>�86��X��� ���ܫ���$
���r<��Qݹ��\���m[�p5�$�K̤!w��N�gL�_޻`��m+�dR̫"R�	d���:0CE�73i	u0��Lj�x�5�6�B�ca���L$!�$O�ɼh�:���-�K|�n�n��#�m�YyD��'��Q �r�n��Gd���������҇~v� ��4�8^�.qE��GZ��%pn�!%S��!O0m�p!g�IX�kZ�p���J��HHZ�'��!��#��&���˦����e��sŋ��GՃ�;0��=4J��P{����CƊ!Lq����}�if�;��<d�fi�����>u�N��o�����qSfN�w@��wUUUUM�{�C��!j�:;z> ��ɒŽ5yVMJ�x1!�bQD%�AP�v�b�i�T(�æ�u��ĳ��Í�!u-=v4��0=�CzI �-�Y���GI�8��8V���o8��u��J�&�)�qLF2�qou�4�խխ�O<#�:p����q��U6ĤTQ�I<��dM�+Y"�2�[*]t��)�lI6���c�F�V�ص8��F�ƚ���1F�jn��TV؆�bS+����UUća��i0&91&+$�IkԓlKp���y��zC�?C̒�1��
q{�*�Ta��2�}��A��h��!!�=���.N�1�P��L���$8e�rkѐ���V���$!���"I#��$U�+,I�f�08x8͏G�7ny/#ۈ�sc.�S��|�N������N8�)���c���;�*����0��,CTͩV��{�K)�}c&Bv7��Ⱐ�f6�v�p\�������&��W�$�\�ٳ���� ���5$e�R�O�I��KPܓ��6-۲�,-��q2u��~	��
�U��x���<�6�f�<�w	�[<��bŋʽ�{�rm���F̺���>u�έn����6�+������$QݣzUUpN����ݽ@�p�n��C>88���'a�6�>�$����||x����V�44a	�%�jCM��ɮVZ�H���h��c���Ubg9f�q�zh����g-��.k~��(���GN����o&�0ɗ��|���|��[�ukuǮ8�)������)ÎK���+Uj�t�X�Y���ΣV_U\4m�N�đ}��QnK����v?�����\�% �L���Y�jv��p�[����!63����,ٹ��0��Xۢź]�K����g�c�=/����8�E�IC�G�{�x�;�)�9*D�8��-�x����I�O��ѳ� I��N�8`�����2tН���:'L(DL:'K(D�"l:"tЂ$4"lDD�����BlM�D�"&�DN��4!����N�&	�,M��Bi���8lM��8Q��xD�BtN<Y��<h�b�ˮ�kqkq���[��u�\B`���xK� � �"$( �������TMh��~�(Ś��C/�MF�b�����e-���v4*�Q����5�CEwUcQJ��W]Q��".#��4OIwlUL��6%��lh��+�G)2�mv)l%�I(�չ�IY���!���4�I�eܕ-4u ��q4)my[%s!\#���"
b�eK%��
(��QGiH2C�e�F��Eh�G������x�)J�aaY��4f�st�.��(�8S�6$��p�Z�f�6�ɢW�F$��C��N��"��wFhj�f��I1A�C�U�h���̐Bʒ��t��DJ2ɌG�b=**�<�Ez&��SU��s���j�nZ�VLr֥�%R*��V�Z�S��F�EN%��Y
��ZZ��j�*�
�GP���Yh�ɛ-�덉8HTX��Ex&�d�D�݌nɻ���Ֆ$n�,E�+�1T�i��.RETN!F�l�� �vX[*U
E+�+mIQ5]V8#uGw5٭a���]��-i���TM�Z�jkW�u������]�w�_��{��j�Uv�����{���j�Uv�����{����]*�n��~��YӇ<����Z�q�#�m�9�{L�i��հ��.��-�܂8���Y��h�UٓM&�M���6\�$]���$CbB�h#2���IZ�c l�5٦�7R����5�\qda��+G6�#h�I��g]���%ٜ#�n74f�:�ҳ-6�d�����3"��O�����;
jc�����-�8�64i��bt4s�$<h�3��J^��<{��1&1n#��J`:I.9l�I�h�L����|��JIK+e-ś��V�RSa\�u���h�.;r4���>g5
�h�ZK�=[�i�ξukuǮ8�)���$O�'J��	�	�C���9�0����cØ ;��t�!�/s���<h���"��0��c1��_ �<SL�PG���(�9#HCv���Ē�79�>? �琳�rp�Q�BK�}��xL8� ��)����8�o�qk[����<3�z�6��m����3����m�Z/\�<��~�����nŭ%�KT�����ac��yy0�I�G��}���lz2Ei�u\�*�Q��VB�r����d� �jr���Z���Țl��,:��K�V�F���8�J4�jc��=)�������[Z�4���:�[��xxC�;/�8��,��������&���0q�:���r�!�~md���-�/��n%��h���1�ν����te�읆��rf"hɓ�lc��g˅��O�XLT��;���L;C�}nIҍx�Ac�>.h(p��Qq�%�J���:
熞�/�q��_<mm>|ۮ����l��8'g}Dl}���I�b�v�)����U��,�s:���4W)6��m4�K�t�q�D�I�'��ΊIU�!ԓ�IEWm�iW-��ݔ�T��:�B�ex���|�m��e���٦���%��A�9���X��M�=�Udh�D�ƚs�~����t�3�tɓ�M�9T���]	���F=p62��J�GM�`��Y�\��<=��mtM(��Gf��e�)�f�'۴$.��z�k�=o�α1:I�"O_8�o�[Kq�]qխ��q�qM��1^J�f	ﺪ������f��xA�C��]:>|`6q��m�*�/b��02�i����J��<{��ޝ�U΍02�&�pIPp�ϥ>*4ZvQچ�2L�C��)�C	�Çm;���{�M-�A�f�5p�F�Q�H�8�0u�PJ��um4Ӯ��\uku�\qSe>���9ڪ��r�L;���~��0�Ʉ!�����Y�� �,g�gG��A��� ��V[Tŋ)fbq�A��Q\� p/��ICX8�� �t�CT8Ǿˣ!�Wl��7c�vp���Y&J��Y�l���2Y��c��-����qխ��q�qM�x��4�ޕU\y��Nbw���	>=��6,tla��^�&P��3�4H�F��%\���Y����2���`�n�(/+1�<\�b�2�M�I!�y�џ��9B�4�>U����ɀ�<�0���|!D�U)r��������:-k�hB��q�.��><t�����6��q��u�\qSng>[��{�I:��H�H&���	],��^�<���Vimrx�z͵"z1�$�;A��|���);h�PB4ІXՉ׈�%j۾%��HSmo.嘚����UW�'\�2	H⤈�XN��.`e�x�X�V��d�*C��h4xp�DA9����"I�>�zgYC����k���c���ΊƜ1�R%��LEJ�X�:����9������e$��$�A#����gA�p��m�G�����	)�)��z��q��u�V�[e��6riU��iYA-�����M��c���ݧ}x�UURQ����4pphdl]���0.r���CwK�4�ǁ�%�ಘ
0����!/pd1���]	���ԓْr	TZ��ȕ)
���[��E�*J#	*�x1����!��!���Xr`)c��q���=p?<)ls�z�Ǎ-�����[n��`�&	�`�&��0�8P���:X�F��Љb"tDD�bpKbl�Bh�$b"#�'JD�tD�B'L�X�&�2i%	�(Æ��I�YD�DJ�mm׍�Z޽Rθ�-o뮺㭩�ִZ��k[K[�0��ĳE � ��E	2A����wS]w�;�����އ��X�I�%��{s�}�v{��q��^3���>��w�n1=��ߠ���r���C{����s8�|�U�ww����{���t��߽�{����+�U�����^���{��U[���{�t�ӧ<y���[���⶙�UUUUV�ˇqg;�C�ݫ�D��υ����֡��d�u�[zj)PE��;�4�������\�M�Wp�і��!���$=
Mk���g�)�e�ǀf�s��������(7��%�ɐ��2�:!��W$�#%QQ/2�lh7�΍.t��'u�|�[e��m9Ɇ�0D��m��x|g�yC�$�{�(�>1؂?Qɽ���AM{���x��ԕ<�Lx��$����%�$ni�ӎD��O1�vxǌ,rmUäx:y�a�}��#!�����HBPP]���0�2��h6�=�:�]c�/]|�O�6�\u��:CǄx}I.�blq��Ke+h�UcI
�e�Ƙ�HR�R�+
R"AR"���]�,H���h�TL�$Ǎ���Y$v�i�����#���),�;U�����&�������Hu+/j��:�E�: �n���V�#���%�n�cĶ^�kGJ�%�y�����0���݅��l���m%�,M9�w��ɝ|gyN���(��'\�tS�=�.^ɐ���%��UTn�py�������=OG�d�cP� �vU��4#h9�ヅ䝏���׫mm>|��\uku�\qSk���Ɵ�޼����tvi�P�;3~#!�ˡ�����\z.m��n�:�x�c��2[�Ե*�b�m@����=�y�b֖K@�zJ�m,�vٳԶL�DX������D�Y<>�x��9�NC�`�F{4&a�y�%�m4�D�Lp�q�6�崷[�:���/��C\�X��
��F�Ō�R�-�s�UWg�|v$����G`���g��U%S�4��F��t���%�%n��m�e�)ĸ!]J�Ɣ\!iS�$���X����]�s����GE�����'�sD�1��Iw4�,I��]�� l�g�2xᣇ\uku�\qV�8csvay�G�UUp�?}���	*��$����&x�p�	����ϊI��6�I"EpV�.	��)���oQ���t�eHwNZZ��OK�����k����� �C�u@����W<ԩrbGX��:{Lm�|Ÿ��޺�n6�\uku�\qV�-<]L�v�,́�C
��&�Ki&ɭE�d�F��Z$�k)(�R�[��#p�Z�qқ�r�FḎ�yi5��Dێ(㨶[v;-�lԵ�[) ����j����UW޹^��Ww,�!��
K�u��('1�"k����LYǂh��;����ŭ.[�dt����:�n��*T)�l�p����2&���5T����m�O��i�CL�Z�U�5HSb�±m$�)X��<�ó&�d�8C����FA~2�3rR��S�N�:"`��:Q�ºK ���UUUUI��p�NPێ�ҫ�r��`��8m��5Z�F����m�k>���Im��[ϑRgbR�� ���k�$4d	)��j�&��w�t�UT����xx�M!���Cw�Ie�~#CX�Ox㭴�|뎺��GG�{����M�k֚�K|�m���|T�ttn��aL:悰x���$��<	��b��֕^%^SeI&I!6&�n�����kI$�Q)�k�0��A�w^��U���M�ǲa�<<亊Su3YLa�Ğ��CY��*��#N:����~ź�ׯ�i���:㮸��q�p�@�� �Dr&�!l��YF.Va2�*��&u�`w�	9�{�a�N�!�x��$����n�t$%D�8:�TyR�CM��3I��(#�7t�̝$�oӁqc��%�6`&xIN�fN	�8
�ޏ�zk}�D���G�ܮ3��(��T��ĩ�����gjQTtۦ� o1>�ǋ��g8'D�&0L�""a�:Y�B&�6"""'J�(M�âtDD�bl�,�f�D�"7""&	 �� �0L�&�١e	�(J8&�� ��B �"P�6'H'D��g��,��0�<x��B�DM���Ǐ	�Ǆ�4Y�� � �"#>!�Yϥ�!�,��U���#��FAM�ͻd���┃=��\��[eE��n)}���N2}��s�3嵱�囅yݩ�����~UjJ�y	I-INOst��=��VG9��F�������4�a���6�)%9*.�k��wt�G	�3�|I�qHr�e�c��&1sd����#��6wsD�s`.��ȼQ��4%�J{v$Rx�7����#���F�M�ƛ����=�8�'��r�m,)�#�s�����B�P� E��p��B�%���C�XB�\�b����7y����BB�,�E
�i$���F�U4�d8ۤ�y��
G9��գ��ә�,�����e�kN�%&�"��;�M�>���Ԯ�o�o��|���.�{����Q���}��%�o��H���L}������X��M.�j;���ݖ���]ZJZm���5���ky\���Zp�(+v��wu���Y)��)%�VcV�K4ب�ֶ3]4Y(�B���I1�c/�Q��2>�%����h�6�©X�(Ӣ�"��hV�3��m�Tx��+���$bQ�ͰNǵ*k���wF�5��s׫���U[�����Q�{������U���}�{����uiUn���{����{�1Un���zΜ:t�M-m��uŶ�8�6��5o1�$~�UͅN5T!,��1�TulyT�7UEH!�.HA��
�ɐN7DB�%#�1ډ`�"WPܗ]�5XۤI��A����GZ�X��2���r���AٶBI�i+���/���ˊw���pq�""t�WZ&ER��G"u��g�0!�����Ĳ6\��I>tؙ,x4��}�Ԡ����v��kYã�B��4pRd�� M#���l`9���c�2J��,�.�rq��od/��޽��$�iZ��Id���I6�3�2�GG�-ý�d��d�F�4dɧ[[�:�mqm�a�Če1�A�%m���~
2���w��$���s#��2u��@d)�o�dn�20n�6_�K�,X�F�����pM�Cy��V�]M5%E,N�ʐ�$-?~ ����L�ІC*S�cs�=$$� �忼:1	,�w��릏4zӍ8�ku�]qm��#����.b⡾I$�Gc,j�cx���ɞ܍��s�t���Dː۳��8�a����,�*L�ЧХmݓvMf��i2�8e�y�~'�)T�7�y�����^zH���Ac�$��<6�C!f����zDg�q�F���o�4뭺뎺��GGe�&3X���y�I��6[��l6^��'*ъ	�"�h�R�!4q4�4�5 ���ÇY�?�ኆ[�0���A�N#j��p:a���>$�a�A���>��칣�={��'�[ˉc.1�X�|u�ϱ��#lsh㯛|Ӌmd�!�æ���F�f�uyU�۩��t�c�,Ó��rN�+'-V� �w`��c�bDT�!lc-e&��	��rE2�tR���-�jM�'T�pJNqG�d��j��.
��Z�Z�"I�+��N�qX�ڳG�M��?$�XJ�R�k�օh[�J������(��vlf��	) xi�'AL���d�C�c��6�CK��<GF����QT:���d:�=	$����iBd��\�����C,��l�K!"�ō�t�"N��|P�����c⪈Uq�=ac8d�2|4p뎺��GGe�<�U(��B�YԒH��q�J�T��./I�Z��ǤG�xǇ����4���b\��9�]��a��ݛ�4Lt�l�)��vlJ��N���+�~�� �hL	����mòJd%Tc�2k�̩�[M-��:㮸��q�q�Yy$�a�5���X��8c6Pl��v�	�����Nt,��$��t;�5~^�;�Z��4�M�CJe�1��m�R�U\��ǌ�p�8�>(:6.��=��Ә���XnQ#7�1�.�m�Ym�Zqm�뎺��GGe���&5$�	X��<%J�|��p*��.����e�!�ƴF��M�MxȆ��9La�IRK�$8?~4!4�%��-�ۉ铌�6ŵ�cg��'%T�Ą8K�r:�6����!�O��']��!W�z5�Is�#"�|�y�c�>|��i�[u�uŶG������z�U���	��ݒE]��I ��nSc�������b����*˔�i�-�h�].X�[�-i�T�vԜUTՒ�T���Ij-bX�+YT�����\�I%�H�>��VIr�w�J\�"�;�J�u��X�!��	(p����9�d���s�cRL���JEI1���-sFL�}�'���M���p`!�l�Cn�&��Yˁ�cC�ً䏓DN�%u[�!���|{��4���p�Co�I��$�/[S��u��6�:�mq:C{c��y>���KaSU�$<0x'f��$����x�*t�ɝ��v*�kY���[I���Dot�V����iˡ�a��Q	]��MU�:8x�4�z;(��w8Ŭ�BSD��K1]fihYw,�.xvh:�r\�q�htP2�n�[���=A"�����p�;㮾|N��:p��:&	�`�&	�`�""a�:YB`��b""`� �$�؈�8"`���؛b4P�$,DD�8P�$b"=�b`�'&�١e	�(�pJ�|�����K�(âQ���0�<x��"`�(A��8"`�<x񇎐�Ś(�x< ��DК4��n���ޗ�����p[�;�޹�-O��|��޷c���or3�j���Ѯo[ܮ�Uk$o}>�vR���I��.��\����[�r��v��}:��U���_}�m����ŭ�M7���R��|Z:�=��{��lyD35���n���r�a���FsW�q�����cms��'�����r�+��w��n�ϛ���}���O�˽�V�r/�m�z�=;V��������o����vvc��\"����s��l��ޞ�z�����d�����'7��w�<���=]w�f5�<�32�x��7�u�^��]��&�y��c9ß}޹��S��^�(�7��|���q.��5߆�N���k�t��O�d>R�z�O>V��E�+�e�s�7�n�7��ޫ�ѧ����N9�f8�U���}�{����8�U���}��{����cV���}�{����(��wwk�Μ:t�m-m��uƖq�q�Y�I$��!!OH!��qy1D��Z�9vO��%$��9�?b�Ca�η�Є#�ک�f@΅��L�����R�3r�I.�e��k��%.�Z�(����u�L�ã�sݨUsF��p�3�:4,���.�<i�����a!�.9	�e��4�[[�:�,��l��I��$�����P$�.ޘr��<~��=���ұ��d$�y2�",��K�-/V�Ѝ�>�va��y�2���a��������Y��4e���$`FI�� �!��O��|2'?��$S<g��H���N��f}�ȜRV"�|c,��:���q��㮞8~�!.�5#�J�[��u����W��'!ia)�ͨ"i �Q��B���]� ��$/jsd9D��IuXA҆Ƣ�Q��3n�f��+�]��-N�N9k���[,B��J	b����I��K�Y^ĄBe-�6��H��c78\��n�FQ�29�7$��d�!�p�����zy;9;'#HA��A������BҌ�؉VӁ�v����Å�.��֎Pk<�X�I	1#��7��$��Gn����[XB�j�����AE�68y�dnO!�f��2y��뎺�K8�8�.�����Z��2Z�׫�Ƥ�D�E=�I��sQ�(�`9Ȃȍ�G�E�2<�	7P�F���`:=ru[nh���{���=0��〪�^G�X�!
ZZY�R9	��Vl�d+Is����{�py��:�#`�_B0�4�g2�I1�RcX��6��m�����뎺�K8�8�)č�����h�b�l�I$`�=sf��2T���aӮ���I�gl`��M��w?XP�X�H�ٴ&r��.BX�r9Ty�Bhƽ��$���/$�E��2���dŘ(��0O��vBK8#Aq��u��in��\u�Y���C��L`}����_�^���$����t��T)r��`�����!(�j,���ZM��ŉeBl���:�2:m0x�⎖̖�%�UjyD�9O�!��i����nĔi� �ڐ�T�F�9*�ccNM���g��c4Y��nSАǤ��s�V��B�@�>QgA�=6�׭4���:㭺��h�L��Oe%mr�ԟŷq!�ͬ����v�h��[���Hˑ;H�l��&���4܍R�R��(�)GFR���D�V�u����쌱�$��I�a]��&Ǜ���z�6�+eYE��K.�g
�V9\�0p��lv�R�֎$�70��>�p����!����nI%�&
 �A!7.w�!U�����b��9b�]#$�.�e��&�SJg����g�4ߍ�=��	~��"2b�+�KY2,ZKFI$O ��v&S?���<T�co��o|�?-��뎶��q�4d�%�$�0��<9�4S��Ez�˃�t�(���j�cF�<c�"�a�Ln�*UPl����0<?by����C��A
D��F�Fưf8�H���s�&ɚM�����3I�.Q�ZH�r.����4SO�[O�m�:ۯ�6����^�d� �����%^�$���E�FM:v0fH&�g���А��;�B��hab�:z�8&�S�J��J�ĒC��5�I/-&*Y$"��%ŗs�4r�?w�Ƥ����htD�g��g�HJ�!,Xt`���J���"������8p�6IY���"a����x���&/˱bj������q����9�u$�����;�I�	$#q�<9�Ca�M:rY���k�D���P�E��aYJ��0e�=p�t{�r��!�'�[���L�:�4���;�C)�c��0��9���EL�sH�1���۝2q�sޙ���Zת�h�C�a��&��O��ҖW�UR�F���k��}���>���>���{�Z��4��T�C���od��f�@�R@BDI`_{�;4ZZ&�Ih�֋KF�4D�i��Z&�-6�ZZM-&�F��kD�Ze�i��D�$Z&�D�F�M�h�-4�h������D�i"�kD�ZZM�M��4��4ZY&�-6�-,�E�i���h�D�ē�7��#I4DM$i�"dD�h�DIMθۢ&��$�"m4M"%�Ѣ&�"h�5��I��ɓKH�ZY&�I��&��$��D��-"IbZ"I4�-,��id�Ii�N�I4�ZZ&�KKH�ZZ&��iiE��$�id�ZDY-,�L�M,�KH�ZZ4�4M���i4�ii�4�-��I��id�e���$�KD�"M$��HI&�2i$$�BI4�Bd�BY&�IH�Gni$��M$�I2HI,�Y$�D�2%�KH�H�H���%��i$$I�I$$�H�I!$�!,��M"X�I��HI&�&�&�d$�BIm�I��-"Zi��i�I4�ɭ,KGn$��Y4�$�$�BIi�$�d��Ii$�"i�ZII&�&�e��I&�X�5���M-6�DIm$ɤ�K$KI-$ɤ��"BM,�F�id���I��n%����&�I�IidD��I��i4����&�%��iKI�KD��%��4Iid�"�L���DI-$�5�4�$����%��$ZI4�&�D��I�q���	�#hA2�	�,h[4r76��!�m�,��[!m�؎u�u�hY�A�m�F�[bƄƅ��X�+ó��uj���:�q�	�Bm4#���hM���n�Fж�	��d!�h&�/6ۂƄbb�&hF���LB�&�Y���4,�X!4&!!124-�Lж�[���,!1	�FB�	�XAfBLB�B̄4&!fAfBmhLB��f�������k-�9�&�"�"h�-E�h�h�܎ZA4YD���Z$i�Ț5hPDj�hɢ"�"D"E�[D�"Ȳ$B$Z"4�d["�&�D�DѢ-!$M,�#H����D"D�D�h��"&���D�#H�H�HB$Z-��\�H�H�-!,�dYE�dH�$Mh�"b,�"Ȳ-�,����"h�#M���D�D�"dB$B$MF��"&���"h��4D�h�-��F������,�D"D"D""k9�DM!&Бh�5�����$Z!�h�h���E�4H��hMF�Z�E�"ȴZ$kE�"Ț,��Ț$kB�"�h��h֋DD���h�H֋""hMD�"Ѧ�E�4YBE���uȚ$Z,�"�dD�F�Q"єi���5�D�BE�E�H�YE�4YE�F�,��Ț$&�DF��Z"$-�F�E�Ј�&��,�E�!b&��d-��E�圳D$Z-����h�5��Z4ѭF�i�&�25�ѓF�CMh�D�h�&�4i��4i��2hZ:q�i�]��q�h�4ѓF�E��	�M4,��MhɣX�hi�Mh�F�kFZZ5�Z2ѭі�h-f���#Z4д��h�FZ$Z�hM�h�hD�DM4Di���-"m4�4�i��$�DM4F�hD�Mh��kHޢTv�yb��x�4�Z�����1F3-a�*�l�����p�Z+��
�?�o?>�>~��>_����}n~����ߜ'��ຈ��:�t�������V��?>k+D�����>
���|Y���:����lo?O�������,��wn��T|�U@���n���/������1��9g�o�L3�q���[��o���o{�c��;��qs��?�m��0|�~��$0��&�@���QT�������"�m�����@?��"ٟ��xR�`�)���?tJJO�M�U�-4�}�����ܧ��RH�;��	x�ZB͙������j�
!_+�� 6 �"o�m��m�=�����C1X��L��|[��֧�Q~u�^�~��gAWO��"�1��/e�7���"F�
$����`ƴZ66�H�+ B�� *K}��ΞQ��^G���@2?��آ"����~���O��V��DO��'�	>������K͹��U��U���ם�z���#���P��p�G��_s���S�n��K����Hw� ��_7�?o����`�eEP�~�1����d��/�~D�<?�� D>C�D��EP��?��O�3�,O�)�??�q�~?���8N�٢���l#b�2�e"	�_I!|v~�~JY��� ���`��>�aL#�(`l�QW	ID?�������^�w��1�m������b��)�äUP\���_��~�ϻ�k�EP�����F~���}�O�W����������������a��KPG�~��j������/�?������R*~B��G�_�?���'F���_=����	�__޷�l�VjVSP�YYYJ�VVVSS)�S(S+�e+��[V�Y[V�X�YMX�B�Z��QMJjڵ)�++VV���YYYZ�Օ��+(R�ej�Օ��VՔV��(����յjڵ55j��ee���ڊڵ
յjڵmZ�Z����+(���mZ�����X�J��jQYYE��mZ�X�P�P�V++j��V+�5b����X����L�V+�j���MYX�V+�5lղ�X�jV+�mZ���mXS+
ej���)�j)Z����X�����Y[+Q���[el�QFV�Օ�V������
��2��B��SSVյ�V�Z�jյQMZ��ՔV(QMZ��V�ՊV��Q�ejQMZ��P�+)�j+ejj�m[SjmEmJ�+(��S��b���6��AA[+��552�B�X��2�B�MMF�V+�l�V+j�X���V+��b����b���b�[+��(��VՊ���j��j���R�Z�+(����Vը�Z���YYZ����ڊ��V(�MX�����j�QX�e)EQYZ��j�)�P�2���S)�+QJe����S)E
(R����VVV�B����������emYX�����B�������VVVV�������Z���YYZ����V�mX��++(��jj+jj+(R�Օ��Veb�l���b�B���)������څ2�+j�(P��[(S(V����(յmY[j�+QZ��ղ�b�ը��+�+S+
�YLPV�R���R�
�b�[V+��b�[��b�AX�V)���
55b�X�V(Պ�b�X�V+��2�X�V+��b���b�X�V)LR�)�V��+VQL�����jVR�J�VQL�[R���)L��ee�e�+(�QL���P+f����+(�����J�J�EeemJ�V��+jP�
P�
5���eeeeeeemB��������YYJ����Ք�����YYYB�ee�SR�fV�JՕ���+VV�Z�[VVՕ�+VV�YMYZ��@~��������j|�D_�������?6S�?�6�I��-��q���^�H���*�X��6.K�Zױ���Cj�Sd������䭷t7�)�XL|-�`��߽0������_��Ē�D���������V�!����G����|�����~���VPlO��lt��������bf1��Y�>�&t�=	��~���>O��	�'ԅҹp�ߞ�/��f�O���r��������?�*�00���N�.�p�!0��