BZh91AY&SYm��l��߀`qg���#� ?���b<��I7�O�mEb�٬ͬ�5-�ҐQ[f�)Zʍj[�kB%P�*�(������4���-[K[l��kE+Jʑ�
�*IAZ5���5��2�m�M��h���5V��F�6�YZh��i����F��Y�mFي���і����Ke��5[0�%H+kH�V�K6Q��w{V1M�6�LL�֔ڂ�+ecB��6��ŦQkZh��Z�[5Z�jͳZf��2�ڙ���j�m���2�
�R�V�m�[jjլ�l�:��iVƵT�  h�Шj�ٷ����YӶ�- ��]B���FuY�F��v2���N@-��m�i��:�m�+�VKf˦�m���4�U�kf��ƙx  ,�z ���:t(��� : 6�\� �0 4��� ]�5��Ӣ���] Ӹ 4:���(�j��)�J�T�J���[Z�  1� ��,  =6�ۃ@ -N��t6�� � �� 
G�{8 
n� 
�� h�@t�WQ�cZ�m�5�Lil�4x �x=��� �[�'@U�Wp;� �t��7wn`Ӡ m�����wv����y�� �  �HT�Ume�ME��R� �  w  �v���t �uF:�X� ;pn � ��� λN�(nи �n�r�:tt�q� h��:�R�хT��m�c� ��4�t(r�iN�ӡۣ�  ��9� );�����4GB7g Pu�X4 �`� n�g��݅M�[-3kb��إM%MZ�  e�4
��� �C]�k��
�q΃T:5����@:�
 s��4@-9�@7`t�9à QjX 4Wwm�EZf�Ʀ�Q6�I-�   my� �'

��p�3tp ��n  wp �j㡭��� $.�� p�U �ѣZlBͶƒжֶ�4x   -ׁ@w�� # ���� �:�@ ���n�� �1�qZ��\  wu�[Zc�(��Zƴʍ�   X�P ��@�k�h`
��8�F0� ]� :�uT 9θ� c�]@���@ 5OlU)UM	���4Ɉ��ъRR�0�0 &#M0i�O`��Q@�      �~%*T       "R4h�&F&�jm54�241=M6�J~�))�*�  L   	�M�oG~<p�
�ʵ�U������kKeu�ke[Lr�W[+�8R���VeK��ETW.�QTV�(*lEv����K��y�G��<>]���!������RI%��QQ]��TEk�ǏUT� Q�� �dAp" bWw�]t�U>WU�+���]��:���]�r���wWܮ����w�u�r�������Wܺ��u�_r���wu�*���]~%����]_r���;���wW_s����DP���%�Do ���wwU�s���뫮��uuu�*���wwu}Ϋ���]�wW܄T3"!�TLȊ��̂�� *f@QS2 "_r�����_s�����}ʺ��wU�.�S����]Z]u}ή���� �����{z��Ƶ}�z�.F�\��5A7n���бV@.T�1�طӉ�y�M��ka$���S^k�cv����!7p=�-V��m��[Km�Pk�%�u������ٛ�����3v�`��H�<� %ْ`u��][�e�A�ζ�|-�X�i�+E�EՑ��z���:n��U��!�I6v!�`Õ�8f��K�O�Z�F&+pL�9CV�+d4����Q[V~�KPO�m�&��kx�pV�̢��5/,�]ӳ�M�cf L�g tJFr�e{B֚��X������v帪^�EؘV�N�7*Rn "�w0Q��3M%��][464� ���Q���mk�r��%%�D3,KCi�BQڐZ���u5�"U�72TzK�H7��,y[��Z�n�T�M�[��۳�50�.�F��9��ΰi�������p6��O�m��)��F�{���VVв�Zn�W�i4EgZ�qf�	*[2���"$e�7Nan"b(d�լ8Tb��eXO�b5��1�T��J�8T5���kt���T��u܏ln�)F���kFɣ����.1�=Ԗ�����Z�Loj]$me�W�����<��]w�&�ѡt�'2CM<z��/0
n�I�g��xN�wtY�	�2����pkCl(Ĩ%�t�b�ؔvs�[Y{Lh�686�B�F���b^����s�/�k��㠮��N�
�������^�o/P}V�m�x�ּ�\�n�k`��@ڕ+4/��cw���ZRE*�r���K˹oP,E5����(�@Gw���FZ���7��a�a6sV�6�ֶ�,Axi#J�k�1MY@��u.�f�MIbkX�hea��%�X�������{�Q����8(�8u�y���0�)��,ڬ��V6R6@��Z���ԠN�H�Q#�K<{�3َR�0�İ�S����o@��R�]F�,?���ږ]eE���?�]͗[�}�5X�HҒV�ȫ]9O0����d�m��w/si�# ���h���=���T�ԧ��&,CqjN��˱[i� ��u�A\�C�MKz�=�)� \b;�� �����3P�$�5Z5�B74�`Q%� f�2�g6dr���]����B� ��ky���ul�#f:�h�+2n��w���+4]��E�[�Ո�)ٶ,
�ӒQh��,Q�����: ��h��N�眖6o	ـ���Y��mm�Ђ��h���3��'�M*���JN��Y�� !�5�z0����SL[�v�������4�hc2K"��c��y
�[�SÃfG���� 7rm�5�A
��ʗz7wnU�躰�-��d�R�R� b��î�|�7�+	r��kmM R0.���&d
Zw�YFn;âʼX\�qc���VЁҋCfS K��4A+t�jƁ��{����s(��c6��(�Û��m3tw*�Ʉv��j���a�`ŏuM��t�"*��\�9p1Xf(�x��"�ɀ"�T����X�n����ԍ0VY�y�<j��vPc��EŢ���Z�����&Ÿ���]� 81LN���Ӭ�zn,�k:թf��ň�sCVM�tJIQ��n�;ӡ��I�+IY���he*��-���nR�Y�Cgư�w+U��[�nLn��#
ۚ�	��{e��	�cf�IG����{����:�&����a���T�����+82S4��Y���&�MI��(Y/)�V,�4v��JɃ�o�ǯ��6n��HDr�a^if֩g\���Eef$,i��Ю��:�-G�_+|s��t~O�ګzEk���b��!6C�:��E����A�Y��iص��2�n�n�bQ��hkq��b�6*!�Y&eJ7�V5��曮\�')��AkK#��i�5}/`�@+��i�AХ��X�Ke�˙���RAU�����u��M����Y�r��*YQa��3�(!��+��d�uki������w�Z�X��`FR���BU@�ph�-jlWV��ɪ
A
�������Um�pJ�nk���c ��N�c,XU㨴��B]���*�#Z�4�x��[�#K[��J��G�C�0f⊃Y�+U�K(���m�JU��X)�	��J{uͪ�8�Q)�:+G^��eְ�ѭ�F=`c�t��ޘ5L�g PM��ٷ7[u���eGf�zH��v�ޝnСJ�P�¯7Fo�Y�\�Q6b�En������-ܣ�b�]�6\On;�b�4s.H��d�����X��2n0�@Yӫa�DZ��.��
a[@`�5T�T5ƪ��ߖYt��1,tM>v8�pʵْ��V���;l�փG%L�kI��7v*���$-�1�BF`p��0��C�����?-�N�nd��ũ�H 	�ʽw5ZN�4�܍S�A\�8�)� ��v���2�J"9��Q`ͣ�[D�R�ˇ+E^hu���R��/r^�X���Wz2����a�++�ءz.�v�h&�0e�L�כ)����B�op�F�5�j�%ҍ^'���	=���^uęN%t�+ ̽R�,� a�7F��d��ˈ���;�B��X�4E]�<�$�B3��%�Џ=N(@FX��t�{L�t��n�At�3W2�X/&�I���šl�4S���7L�_a��tV.md��$3���Ѹ�e��qDŴ��#5���H��5}b�Ob�˥4�L':��M�H��y��C�1�hee�U(�4B���:�O�w�2�m��8�!5I�޳E$�s�ba��,V�K�j�=���̛���&���o]�b���96��Sɐ)wZ�MB�}S+F�z�6��̬R�#��Ҳ�����5+d�8�K��Nk�*����8�"��Ӄ�{��Э�Z\7��0�sZC(G�)3U��<[�؉�/T�͠u� ���r�F��L��@���� ܣ�n7h�-H����n �p��6XyJ�ث�XEZ����Vk))����i�6)��v�D��v�ى��f�4����{YqC4�Q��ԗn�ڒ-�]��zaaC#d�͘� Y���S��@y���/Y*�hӬf$�Y6���N�f��P?lT���jX���Ȃܶ�hx��/ 5V}���m�P,����ɸ�0���d[r�#l�x��蜽�(h� ��K��
�5�q��b�f��*
AI�^T�H72<��{lL�%�U7V��bT!��U� Ԭ���Ċ�Ȏ��JMZ�gٱR��v�hi]V��hAρ�eSr�e<�n�-mJ��yn)��J��ͻ��Qv��0%��ڗ%n)��n��;r��b�
��or"���(4��߅LJUC2݀H�EH�N�Fmu���3�:Nҭ�e�4��ԇm`ۼ��"w�u+\�F���xws5=�B1{Z����ܳUv+��]>� Biu2o��X��f�72�^֢>0�i�m�֩J1S�@,p3�&�l8/պ�S̔�DM���Ԝx�Ӌ��267.�\�]#t�K����̭
2��4�}����ZM� *����A����,5&��5�nU�i��B䗉!:�R�7#0'R-0�kI�`�ؘ$�Hd��J��"v�Pm�f�3�[�����)����*9GE�Z`�Hh�5��t��^���Ea�*�Ǐ	��Ikq�ݬ�	�s62� 䳺�+I��`]h�5ާV@fV����fLMn��Lr*��nK�J�I�ə��!�s�C4���d;m.l�@yX������s2��mTy�nX��<P��űM�M���FR2�B1����oV�k.�mԿ�w"D���Ʉ5�!����E<Ób;�i8�S�CŎ�>��V�R�7���qh�c��3
�n&,ܭz2GeLYr@��IMcҶ��'�Ȕ�D�a=L*�c�ķ��Mҡ@:ɂ��pԻ��1R.�j��l�Rႝ���6�1V\���n;Ô)�0dx5%H\%��ّ頵�M�aeаe17��.�=6"L����RR�!X�*�;��}�+8�Ɖ�е"k10���Y>m�`� ݤ���jb�{��:%��{c5K^���]C}j	��Z�������̺ǹ�δ�E�f�Ղk�VL��L�9�#�H��_z�ⷘ��$�4V+�+&k2譨�C@�'\��K%�K�m���!�5�qm�:$�rjGt�s)R3eV�nـi�:�m�h#�3"�b��'+n�P��өFދ**VJ[D(�v5�wnhp c�i�u�ߙ��i�{�bcȲ��^���p�Y�fP��n�cʷ,-���Ip���.8������`B�)��	��^�ݼHD%-EpC����v��)j�q����-w@Y��f���@���/��͛�G�X5�$ň��M�hU�Y���R<�������2�EP���v��V��{Yt�
-�DZ�E�{�U��k-<06T̺;Y���/�oJn�'����+1�{���,M�%;�+̕5@N5��덽���hص�eZ�̙Kd۔A�c���w,15����A��x���4��ܴ�(2�J{�I��u9����l����J����n�`�]r�m����F�B��kiEb��u�:�Z�rY�1S��LҒ�$1�aa��2XW�ΐ̶24,� .k�-!�Ҳ� r�eaF�20
w��f|u/��ݶɒуb�mn�Q�M����{k\e�Q��2^�u���S]��Z�ۙ��`lN	.��{MJL,�2���J�����pV|��h��A�&���֖�'V� �d� �z�V���)��7��X�li�76��f��%'mN�/6�ڼ/+�u���X�Lz�<���p��3`<Z�f�� ә�d^TKql�ubU���z3][��EW��٘so+Xˈ���y���mݱm�[I��V.�j,k�|"��������YB]��j�V^��`xrF^�2Ƙ\�shTP��@�ßE����PEt���+�ڕ�#S#��N������ ݡbDB� �4[�jd�*f$3,'��+ a�d���JB���X]yV�ܰ��B1W�SV��j�:鱴�'+ij�>U�LT�r��-��L�"���G�Ec�[[V�7aR�-��}��Zc3�͛���i�Ã)�J�XiU�!��N�j�����ʑ��� �w*�+6F��r��ZA�ҫ��h(<�7d�&$����f��R�*���/s1�
Rh���fs%��h:B��v��f\aeD��B����7;�oi�;iwV�u�s��Ԟu�e��7�&�Ksz�@hs[F�"�W�tP��h.f7,��kn���$Dj��*З��K�?a�$L�ʔ ����¯J��4�P��ݭR�+8V2F���;��G������ �*�䌙V��W���V���e�!Z�N]7��%'wt^�(�KĖP�*V�����b��;��T�LhγN�F�e �b���
0Y+&5V���e�d]�6�BR�q/b3i�SMjOTůD���fht]�J�NŃ+�����n�y@޼U�r�ɫl���Q�ap*�f+����f�(�̏KT��'6V�g��۵��[lDb��q�����w��mYw�V"�v�%�#k�\�x ث0�ѵ2�Z�-�`�4�f�1���m�(�t��!��Km���.�,���qݎZa�mcu�0�E�/i$�#2R�M:�
�A����ԧ�Rm�X�λ5!=�����L��Rr��8�;t���/
�K]b�2�.���K3l�a��KoY�Cqͅ\�+o����`\���t6�
�R䡱�SY6�eEl�Ӳ�ւ����Ưu�"�K�]B.��2d���+wn-170 m5HP_"�@MG3r�� "�h65O���Ӄ	�0 Gr^�S^ZW�B�,�=륊�N�G%勴:��v%�ެNj����hlpV��@��x&	��R^�� �9p�dT����Y���h��6Rf���ܤH-5t v�B�$�;���/4:cC��j�~��Q���`Ul ɼ��n��v�usJr9��*'D�O�/q�ḍ�!b��ЬA/rよ{4n�&ţ^D�%jd�䬆�zL��b$A��N�a��e���J{����
�k�[j��z���!'Km�9ge���̒i�xfT�V�G���`n��:J�MMF��)�ܨ�f+���%�*F
[�I������]=�u2�I��ڼ;�	�(�CZ�z�k�Ѐ:���&h5���Y.�g�A����(�Kݹ.�A׫~ȱ;�(�5Z��wMAs+~���Yb�
	QL�U<T��b�/qƎ)�1h��I�-��&J�әy����2��Nڈ���RV�k��7^&]l7���ћD��j�d��I"oM�9���*�55"/FJ��am���T�Y>�F�A��=y�9*2��e����cU�ځҖ+la�1���VFⰜ�x��svJci3(�Ds/X �aM�J��,�Ą�(,��)���w8�nE l�x�7j,�����e^�5YL6C�m��	{�]G�e�(I�2�DƤ SC���N(�:��k�Q��]��`v�f ��in��ܦ]�����	ɠl�.�2;�:5j֫�E*l�F��a���9�l�h��jJY�滶���Yl��'-�]�sb5�ʌ��+4�cuu�j��u4�P�=�p�{r�3>���5������4��X���H\Wg�Iտ&�{W`�AF��$*E'ğ��Mu�I]%7��vGF����X�Lr��;נ،��D�2�*�N������⽐3�����F �*���o{��@�}$��e�tM��[Y�l�+��d�V�íI@��+ �����Wvl(�e���:\ �;#5����v�
XҦ�Y�O9#s��	t�ۛ�����17�e8���[��
煼�f�5�ٳs��w��ˡ�B
�rAJ��ع�ҫ����jL��2RhM/_��s:�f옸�*J"sFe��S����H�<�NjY�ۗq�=Z7�A�n�ʝ�`m*�vQ�o��Wm"�42���O!�s�Y%��u�B�=�=,ځ�u�n3W9�ڽ��r>ʛ6��k=ݕ�p��gٸ.�L��u�*M�ʷ�9�qYg[�՛�y˒�'���Y��jM��̡�u��v��ր�t��U�80Q����!��WuZ�����ܺYg���5�tA&��0S�J7m���V�oKf]�>-�i�`D���f��$���V�Eu��}������c���L���od�-�WKëALt{�U�ضX�˳�j '��)���v�^�8���6�+oc]�Fuμ��9& �k��K\�{��R�hw��=��:ᒘ�����+3$t�᷅�Xi�f�G���x,f���[Ĭ3U2�Gk̓�:f=yt6:ܭ�ש�1��'e���g���89N���J��XS9pa��olк��r��	��� Tץ=+��K]�R���;���N�������?�N]�h��q�7]���������B�]`�mq�H�ʼu �(�pe�G��U�{6�7n����'/��Rͺ��#��B�M|6� K��7^�H@�m�ӽ�>��-#�2�����ks�S�۽l���6����r���`�9�U��6���W��w4�=@����R�c�TF�n� ��6����=�6�Kۧ*��}3����k&ژ�c����vz��ډ�B�5GGU
jtuv(�]��0FzӠD/r-��@�D��z�mn�����qRg��Q�GYS�d0�;�&HЁN�,�s��W1�:��-;�<�]���.
]�kt/9]cOr�>����O+�$m�w�!����vۻ;O�=+�Յg��LN}hIs�h]�L�C3�,��J���v��OHyA]H3t�4]$�e��7~�ӯf�Nb�}��^G���=)]-M������Y[J��yC��6�3F,6�$��%��u��w����7��Gs��K���51�7��[�s�]��Β��k�Rn�L��e#���H戹��k��ѕ�7�-��Aܺ�&
avC�����}�%0�sL��AP�
���<�5�3�����x����,�rcDr�s���{8ծ�ԝ:�{��w���x̩���H�Η㧫��ނH(�^��6����,�}�)F��Q4��n�����}�F��σ��Vv�3�C��tj�!^r�Ҍ�J,�=k�+�����5������C�u@�-�
��}C&�� j�̬z�f�a�;s�V�0T�f�רj�{��Q��9.\+%��`�a|��N%�����CǕt��-1cr�:��]}Ӛ���CL�U����r�d�q:��w�*؃�6�S!�pOz���x3�E��cx�1�V4\�qǙv����sy]-h�M�����\�l'��x�f��]�Ӥ�L�"��l=���&�tB���
��r��W�4���1�(������X�Z�*TV�n����֨8�Q��ԣ�9��tz&���a��������O�:�<���_p��K�,w\ҡ/c�����k��1N|3�˩ˬ-�X%M�svd�kX��Ѩo)�e�DWwvzm^�yF�\#/4�V��Qm� �Y��}�v2W[��V���Ws4�t�����h櫇�X��2�a�+yS͠�!}���;��I{pu���"��Ū�<ie<��<�F��K����2.�b0�`���6;q%Q�;v�mUg�(��s�7��
2^=�ٴ������e��u��
ҋU�ёa�;w(��_9�:�G��+�3����&��x�r�h�p��N �7����(�- +N�ɧ���D*>V�&f<�����Y�2C�D+e�U3����ڲ=|2��!���Y]���F7}%\�$a&,͚uƠC����K+67[2��{x�-�o��>�K[�l�mখ=�$;���q_ث6]�s�J���Rb��^�	K$m[�oSM=͜\x�<�]\��#�Ý�d���؛�S��**�*� 38C��M����z腌0����*T;+�K1,�Ht}�)��(�w�x8�rkot|ݻH$9'�fѧb_i{[X��i+��.|r.�ީ����m�:^�!%�y��ó{`� j�꼕7�
R����P�Ne^��9^(���DXٛr�=��:��	�B�*�2A�ˋFf��*����P��� �μ�N�+�`Fk(�XG�t�c�Yf9J�p�g^�ۗ�0���G��0L��m�|�7o`�e�Ѝt"��#����5�o�$+�uE�� m�ٕ!��k:��ڔ�u��� �*���T���7\/4a��E��$m/�#��(�X$,�/R�����HVf��}S@��f�\lV�,1��1܍$��������[\N��@��a{A�ܾ��南d��a�R��e�8^ʎ������+MB���/*+��n-�6���!`�1��\c�J\�n��2�X`Y�_Y���'u	c��/�9ܵ�T�����G$L-�Ǔ.��҈{}�f��RV��Q���3�"��2_Ӄh�u1+���i+5�dO2�K�)�a�ǹ0^��$�m���؃�v�aȅF'���O/(X
ٺ�m��lݧ
��5�h�Cw�~r���`��� ���5T[��Y�^�ڱ(�����u�ͷ������"�sS�e]vN �-��o6(B}}̝\\�������%����ٮ�j�\�A��w�\|�Ķ��)���y�Y�x��t���̤��wtGc����
}*�=��b�}ȅۣk&�k�A��!�8֗��\�5)��W���J�]���{������n8��_p�l7R����/)�{W(��a,���B"�5���R����ev���h�YQ�x��A�Keˊv����r�J���z���|�O� Z��&��Y�^ӣ�2��;��]��w}�`�椑�|e\C��Ь6o �t��dҲ��Q��)C�I���Q�W��)w\i����ƙ��^����i��S�ㅖ.�WF��C��g�ܻ�/�]m�jEz/8�=��u�hD���K��ea�U�5^]<�R"O#ǬjΎ��=٫N�w�&�DY��ʰ+&��C�@�Tx�:���r�B9`r�v�'g2iDB�n�!Z��w4M���7�2�IV�G:Cjv)k��kqN�8]d/�J�fN��OuvV��ӥ�P�]��Q�<�t�B� 7-m�T.:;4���K3Q�Pݎ5�h��	�lNs�=i0WV���Au����ظ�8�V�	�n5�q�4��F�qD:�^g\��*I6�zp=�� +;F�-�c��_uJt̋
�dD���	ڈ*��3�m��U���$.4�T�Z3o�R��]�[.[<.�3�,�5̲�@�Gho15)[��ԷL��\�j\���f�v��
��5idX�B6*|�T���$d�g(r'ŲK��j���!��a,�;�qhlI���J�;M��Sp�gwb�\��qS��T�aĶ[4�9O8�BӨ+ Vy(>Ӕ��Z�
�H�!O�mœ����6A���x�F�J�d�F@�Yv>"H�9�c"���G�)���nkʱ|Cab:�C��-�����eJ
rێ��i]��j��B9L�� �u�����nN����@2��p����iTb�	��cݳ��K���5�v��������i�zv���8��RWp8�@Ⱥ���o�D�7�(n�{�D;�|)�;�Ro�0����4���:��}t��ji���d�|�wj^�2w'Y]�C+�١.�
U-������w�ҧ��X�C�u�U4����w6��;�E��ܩ�S��Y�S�c���������N0VR��� ��kgͣ�d�-�wJGyٖ7�=�@���!�S��̛��kb���0�aI^N��L�%�DK�,�r���wmQP�����c�l��&��V�=�Xie;π��M��漩�$c�)uX>mWٽ9YJm�pu,Ķc�962�;:�nFzɲ�,�F�'gf�һ�pY�%˜ɵ��[Q��J2N/���Q7�)��|�ڲ))g���2�Q��9�݆9z��6�ǁ�GMA��ٷ><��fʨ��Fp�-����׺շ��)}�>�e^�dm��ŦX�۸C�I�n��i�R���+e_QiS}�"`=K��F#�ՙx:7D��|n��4�#SH�1%h]��p�����m��`&�֤�z@���#�;�ŉq��Tf2b�'�c���,�q��7h���f�#��!���R���訬eՖ���a�o��L�e�YD;�=y~\�.0/f���,fn��, �>�����:Lԉ(y3�,��V�n�&G_Q�'i��,��	yc9�T˚��nj%�U�55�tv�Ů��۝F!V�u��g^i�ɡ0s��u��,�ΨX�v����4��˕���v�`�g{���]HwKA�Qw����v�$�[4��.����8j���gc ��]�c�S�L�0��;6�G�^��㿲��Mݹ��`gK�2(_TT4Wp�cyt�1wS��fΤ*���!{%���M�Y��O+�;�������[h��i(�-Z �Ó�A���Tȅ��{c]^#��/�u��X�_�I�܅YvBّ��k#r��W�W���]v�,��~|�J:^p.]�'ʗ
je�:�`��M�q�9@���+s�wq<�$UAwY0���O�����S��V�V�Җ�^��'
��Jl�gSw�V�{�Օ�:�$���4��*5Q|�ݩӳH�70�]L�l	6�U]f��wM�ρ�%*�,��Xll{>c�JKv�V�g~oumB�mZ��⫥��4�G@�a���:���v�R.�vw0��bT,���2�1+�6��̽����-��w����)T�7 =}�+vBe<������L�7��9g�CR�=6wb�:�3.͐DE��f1�Ia�2p����������"�Тz��
�,�_DG+ʛ���4v��}`�ZG,�]�Sٺ����/�H�I@l9}��	 �`����b�/-�9��e�]��׵��M������H��+��-T�I���M��8���R���T���ڲ�w*���EZ5�����a�~}�*����ʽX�O�hR]Օy��e�:�C��ۍ�F��-�F��s+�'N�6{��3ި��V�
� �x����H��u���s�n��/� �n��u�.!`2�"`�:+ Pz%C6c�VZ`��W���#Ud)@<͋�r
���>��h��J��W}ݷ��:/�hP��G-4���QW�@N�Ypȥ �b��]�'-��l=oQ�ۡ��v�j ��)us(P��I�� f	����#`՝̖�j�W<ڠޢ��sM��XDTp�Yk��
�ؚ[�:�lL}(�ъ5��ѐ����^Wa����)�"'�SdL���A�w6��i�3���Y�[֏�7A�^3&��#1ɵ�;a5���.�v�H�(r��,��&��)���EW�F���Q�p�����ous=�PHm��5MC��.�(� u�LK���H�9��$w���!_cT����T��QVaIb�.���=B�Ż�ܣ�aѵ�\r�-��q˓���a�Ƥ���D]��{G��Y���ݗ���ȼ��̥�*�]�֩�7y&����ft�'2�3-�ݛ��LROl4����:�ŧky>5�-�ލ������fK�j}ct 2W �T��&���6��띛[:f�D���)7���婂��Vl-����y��H��]$7W�ب�p��v�f�+��C�$���!ֻ�0r�N�5L�n��o�o6�UKju�!�Z��������F��Z"�1�
���ۻ�Վ9YB����l��U�NO��eS�m�P�Wl9*���3��X:�j�Ŋ��6[
.�΋x��R<ɀ�������0B�_<ķXy�V�S�q\E�C�D�������x���ꆖ�G���b���}�owe��s-0.'QδT�t��y�����
q�Y��!u�}�ˡ��p�Iد�����:�um9�N�y�7�ӧ�)><	O*�CFE@)��rn{\g�}�(�Vkrq���D��KN�C2����a}�j8�R�Zᰫ$w �ʰ��`�|:�9B��]a9G�J6ݲn��.�Jh�s�������=�|���1�c;���`�:S�콽�#��J�d�Rv&��{̸kz���ĦkU&�>�ڋp��'	�G:��W����t�g`ܮ��`t��M�|��s�ʴ轅���a�(F8淚��fm�7���t��s-^�G���7%Fe�&�4�X���{c�vR�����l�OvT�|6� �@�
4��t÷�j�b�gq"�@Xލ N���w��B��X+�ec� ����8aU/�
�C>�q�"�3��p�����]��D5��� ��=$�`��yǴ{�%��{�����JֹT�����i0��+.9����؎(�wLל�mM�yX�opV[���v��\�����Odi����i��pw|���Ř���9򡂏e7LI/>H��zd�G��T�k��r���%Q��2E$��J���\�N*�n�L4�P��ڪ�5�.�p�s��=�>H	��_P�[��RE$)�M%E&)�a �;)�K,���B�
o��>y����羾^�Uu�]������뺐Uor�U�/�����h*�����6cѧ�������w'���빵�7��}Js�M��_eCT1�1Ps��a��
�Б][Q_�̀�����F6nW��fn�m�D��s���_Kq,���+��pQ���&l�VR���ul:����0W$h�
|��C�r�)4��̚n���S��bx] U�ƼF�w[��L_����KFP]{�F{V�S�{�7��&7�n���֮Ֆx1J֗ǝ�{[j�69���n���*#�M��DrK��=�vPn�L�oN0����M8�"WKe��!��6Ĵp1كsIS6Z�0�R�vB���v���S���hl媕 �c9j�|y��\�T��ff�ٔ{�f�NB��`ʗ��w1��Jn��&U��{�6��-\WSfP�n�����̵���`��1e�a��o���-'΁Ȥ�Ѝ6 �{y�&�,l�r"�u��T3͢�j��/z��uNB#�p��k�,�\��Ɍ�Л���au����S6�6f�S`�sȃ���/�(L���N�N�Tn� pZ�d�DnN�4��iRЬ"�:�91�&�RX��t��.�6+7���=�Fqph�i�
=�%V����$1X���k�+�v�7Wɧ�9��w_���h�L�٭��d�v�֚v�#͚�e坳f��]�nޢ(3�OS'T�z�׳M*N_\=ni��,uuVT]���u� ]�ʕR᝽5��N;���R�p����[�b�� �5br�j��)�hQ�ݰ����r$����'J��t{2������3!^cj��^�QA+vr�Xr��/Wo���4h2wo[��.WMnC5S�C���h�=�;�����"@o ε՘1�m�����fӖUd3�Yr��V��O+y�%����=n�,�r�o���,�k\�[��y�$tp�<c�}l�:d�Ka��-��׀�l�>U�j�,�oh>7G�f�:���]vr��"���>Ħ��Ԭq:�$%�Ւ��wIk<�J(g�J�2��\(r��V��N��-��٣�;��W%7]SJy/�=cv ֛�MaԨ�5�"R��,^��k��]B>�l�-�ҳiv˲�+.��*�Ƈ��dj���;c�����[�+#��}�,��{�mIY�g��3R���+�ڈ�A1�f�Z4z����Vl��U��)`��">C��ݐ&+#�W�(�0غª�n���U჏;���>v���

Њ��.�B�U�AwF͌	���&B��iVV��Z���y0��۳YK:�����'$��v�]N�)��>V��׆��ZDV��"�y�u�h.��Қ���3���Ra54�O�s�w^���Ė^��^X<�K�kV�ce���1��j�''��T�s��s��mfx�\� v�fQ��r-"6��9� ��^^J������m:;��8�>�8��h�Ў��999��(�^�]�&��z�bI>.��X����Gq���nO���n햢�X/�dk-f���c�qkl��i/��n�݅A�`f�͜��7�u}�h�TDov��]#���(S�,�� lu	}%J}k[;���1�jh	:��G76��]4�,�5�riԕ
7�M�ͣ���LK7ۘ��<�'��΅�*@`Z��xƑ�ɹ�Whʱ�3K-�J� �Ԝ�6�
w���1zK8p�ܥ3��e`��j�U�1ʛ5��g�̭v����]�搳 �3�+�"�Z2�wC�%d�)uӡJT�lҭo
@���f�p?�E�X2�߻+�;�@*5�x!Ƿ�X��+�o�Y7"�S{�����֥L�C�?]��2�n	�u�I�,a�Y�gK��2*(tL�h�U�%�yL�G�k��7�e���G#nMh���]A�p�,[��K�����>a�].��X�6"�eљC�)�����H�x=�z��\C��/;��I1>eCy�lȲ��M��W�k2N�2����u�P)k��]���wTi�u+;�R��PN��X�������7VN��Y��l���f�gܗ�m��˙�Y*ك�"�q�ͫ},垳��<�J:/��6j�wi��3��)ʒ�ġH����`�A�)*ix+�M��άS��u�w�����ͧ}���nZI��fmmQ��A!p�ZP�i�9�FW:�`rzX���S멯�_:}�JW�z��nj�4��]q�M����DJx�9[�xǗ�J�QN��L�55�q�{Žԭ�����l7�u<.FS^����ֵ���i�R&�v�L��(qL�m��.\l�Ε����t:W�ܽ�Ȫ'�'*V %�Yn�mG�5;�f"��Xwq�K��&�U���%���j]wF��S�ݬ�)8/�J:M�Gt����-*��X
.�D�������q$&�	T�����k-�l74wVm,V��'S�հ�������q����uՙP��j�/�J'���`��X�F�!,$��X��F{.���FJ#�+X75j�7���Čz{#,� ��RT�o��I�mu�޾[�XjN=9�}.�u#kQ���7����I��(w8'�*��N7s(N�^���"ʽ]�f�j:ƌ�uխ9�r��U����ei61��4+�4A��>P��@�3u���iN\�թơ4f\m�5·�h�	�8�cf�ی�ٙ� ���n���j�R��S�g�U�]���F�������w7�:J�I�"	���I��;iDhr<�Z̫��6-�
s��Y�{I�Z)=kx<͜��7rgtIقƱ�Z+2T�;�fe�4i0�5ؒ���loo0dT�3gn5*����2��c/�	tGbզ�SH4�y�jP�op2%;��a#k���njL޼7���pj��hn^'#k)�@"f��);	�o���l<��|�76X�
ʩn�|�`�t�k{��T���2��ţ�<U��V���[]S�[Zd�Bf^��������ۡ�	��o4	�ˁBI��d�$��å�͡r�w�]&^^��r1�LX\�#y,�n9�q7���@��j�Z!�1�x�pg�:�=�`#8����EtC~:�K��t]��¬�Is!Ҝ���>N�V`���,A.(U�s�5r�!�	im"�pWB̸�6tI�� 6��N�KX �'�o[�DW,�Hg_T���å3��u��\m��]/��P�bmbtr�ʢ�pVws7投l��z4u�d���Ӿ�|�Ќ]��VB:fWR��ժQ��l�����#�E�����⩜Jnv�,U̗d�M�YN��V=���I���\]��V���̎N�ZA��޶+ba����<�V��Wܱ��jq(3|7(K�C�$�e�5�N$���Z��N7�˵���kz�u�欘����H@Ƒ��/^�p��&�K���0��݈���+�/j�z��6^k�͗mB�ޝb�N�Zz��d<I��3*w;1 gi���(�!Z��R�J��}/�e�4܀.�X��0L�Y� �u
u(=��-
|��y��Ĥ1��1���db�|8Ժ�SFj�O���ż%��ԗGK��$����iu���vIU*K��Eښu��!�𩺸q�ޜ�`��V�o^3*n+B�-RQ:�MMK㏊@�I��-g�B.�[��L����7n\�;(���64'vҫE���5y*G#��V8����r�j��z����N�e��("(�W*��mi�!���M۝,��j�8� �m�(Щx�U����PP&��{po������������WY�a��vՈ1��F�+Ӕ(4�æƑ�kE��	y����9 ����)�)��<p[�+�9,�F{4E6�`�Z7p��m�ݷ�1���	���pZHwIK�����c(:,���8���EF��D��!����c�^#t�����9�9\s'��
�"d����+q��떄;��fUp�N�V*꘸tV�p=};��wa��}����.�(:�YB��*��@�%�]�����bҏ�5�%�(I�v���6�*� c�.�L�&�D��.�g�qr
�]�s���նS H�ȍ�6L����ˤ�bԞK�2�f���er��o�M<�U���{��]�[��}���S�i����)`
� ��.D�p���<I�Zu2��xLrQ��)�|�
����h"$�w�w�-s�Z��<��=�Z@���e�N�8�=��Y����ȻgR��=����ob����*�M=j��+�^}"�+/��짫��c�s.�Tȝ��I�n��юK��M����# �f�vu^���q�P����	M(��Jԍ������ʜ�G�L뱚����|����Ri���s!��1YA�����%巭�r���\���S��e����7n��+�hs�)nVK*�Hd��$�1����f���L�� �ޣVk0v���I�|cʾ�s��t�0�ѷ��"��
�2�G�V��e@j�ȍ
P=AԆ�f�^��՟u϶Ѽ��Y} `m�mu�����V�a��8f��j�r�8�s{._R��E�"�ղ� �m:NV*V�lܠ��ԑ0��`�l�W� �NHk��g�ʍ��\�;*�ݲE�Z�7o��*U5�R�E����ˊ}������0�5��F�dn�C�X"�if��އ��(Q�3ql
��.M�����)g�;{-�Y�k5�JP���㒉�]�v��Dj����L�A���;vv5kɏ���6����Ξ]|�J��/]Ni'k$n�N_O�̚�b��
V�+D���M��=u�S���j���������i�f�#Y�h����sZ-�RZ���d&}y�T���CZ��!���0;�Q��(V\|��{�l'�Kf�ރ-#5EwR�>:XG�>��xkt��ݧ�Aᦖ���$�i�7q8d�4���hW3/��xnn��㷫9f�:�V��b9ҥX����(�|)\]@^$ �4�ݾ�^�#�5d�˝���e_]�8�g�e���*���S�L�qz(5w�	�T����(c�����G�C��X���4\�-@7^r�H�Ԓ�:�|�́_j;{�R�VkE�+&�R�$��н1i��R�P�m�e����3	6�\�ø�n�bœZA��2d�s;��k	{��e��6�lW�ë���ۆ�5�tW�3�	X6s�% �i̬;�r�X�EO�k=�cZ�._dwڕ�_�1�,�+�3sK("i�fվ�yگ��%#mv��"�,���m����*
ت��۰r�I.�1�S��y��vcn�f;�������p�;	\��f�Ps�&8,e���3Vc#������Ե%V(/e�T�jrk(����8��ޖ�Vi4y��16�ַ�	�Z�e2^�;ѦSæ����.Yܓ�9���*aSb뎱x�n�Б��VkT<tjAvs���'/jޫ�8:y�m:(��QLx��O�,v�	j�V�/*�HNW#P��9R�Ǹ��\�`12��1�-M��c,�s���U)��oB��{���3%s)��_Mŏ����n'O�/�b��}p���Z�̣��)Av�/>ˁk�a"2�"ζ�{܎ٳ݀�O37�嚺Z�^�V�57e(�b�6�iJ۝�9(1[���cP�����ϖuo2�tE�_dN��zS���<��H�]#;��n�d`p�Y��F=�;JL�۹ζ+�1u6�[9�N���=��,�׼�%��8�a���@L��:"G��_]�P�j�K])�漻���m-5���_d�JD�u��q'u�2M����;�֒\�<C���
����._N>��[;n�S�-[v���]�4��مa��	%���Y��Ӈ��f�!hu�f�)u��d�t��5��Z�ͻ7;o�D�I�:[������-����.���j��X�m��XN��X�p�-&L@L�m<n���� zp�����[��l�ݤ����z!O7�P��t*۲�g9���=B�
�n����L�RQz�P>�[�^����mn�uw%[�����CA��hA�W��p=�G�CEk�#k��i�fCy�h�P�R ��>B��?B��L�-"Һʕ���sg̢jIX�`�o˺�y �r�˸f���j[L	p��xÑ���q8�̾�(yf,��8���BNO��"��_s���WW��2�+���Hɔֽ��zȣLmp�D:�v��Er/E��l]c�E�����&_Tl+�ۺeAذ��ڡs�g�V�E�F��z�R	���Tᕷʑw7Y��]�Li!�7L�,�$Ď[��d��(��n���v�'t*�^a������޶������Μu4f���(4�n?�[3QV�H�z�s�;/��htǫqL���7��9o+oah)��紤�7�H�bn��������E�AVd�f�kze�4�ط��mn��G��D�r,WV����Z�g �k�{z�p�.6n���'�z�Nv�Kh$��-8{�8��8�".f�%����qgp�XY���x]B���n����4�9X{ ���5���#{*>}ն9�&GI��uܻ����4l�I����t�+G�:*�����z��V6�}���ƈ^��;���Mt�J�{��M&.Z��Y",�\}�y��ԩ�,� 8U�*V��[÷{���;���,�R�7k�9Q!y{�а8:������AZ���'J��ᾴ�J��ٵ�ܵX�㋁u9롯K1�>����ݺ�	S�x��P�Z��f3�v\��0n�Gi���:�%%]���+V{x��%�����m<]!B���q�G���˻G7�]��`c�-r�)8��f�҇R?4K��jO�y��n{�� ��U��;b�u�!�Y2�D��RoeX�'gQ�8�t�b�������FE+��	})J�L-j]+j�K�k�X~z��TWpv���9���dޛ͆��o8�nC �0�Yq�-V�4��w��-Uw��rm���η�k;�w����f�o�36'�g[�1rm�R���&�=�cj����G�n����˧-m�W�+g<6Uɨ�rSQ��:+�u-��u�����ޮ=�8p	5�+�oK��Z�%ur������_T�k����qP�w�C#;Id����C[c���#�R��Ѯ��mϋ����;f�m.�e�`�{��*��sw8����{b��crmr#��H�<i��2�6q"���<�U�9��n^R��Gb\�3����PwPAZ���b�7���/�U��=t�M�2�l��wO2&�r�^<X�+�Sb��R\�7�8J��mc�\o���E���=$]��]�QcB�v�o�N:�`��n���n-s8@�w �<��^��3�_���g-MS�`3 r��X�I�D�v��f��T6ܽ��h��wm��b����������"�tQh�5R.�f�b����8#�m�6����ܤy/#v�z]�g@9��4�a�ݪ
�.k�ͳz�+�FS�if�EG�w9�r��Q�+l[���-��7�5��u؆7�O��Vru�3�	 wcm�ю�c���^�ض�u	}-�(|�+�Z��{ȹOuI���pn��C
�����Xz�r{p�d��60�F���P��86 �rf�*+A�8�u�owIwTn��?���GB���n�r��m�f�9l��Agn��b]��"�{ל��mۚbr[?:���Kqϖ�^ځ�$O-�6�;��[��t�]��A	ܴ�))L�$km��shDֲV5�m�`��E��kص���s��K2$p�4$����֎r�B&�i�����ܐ�`G^v)יm�kvV���k���aqv[��oZtD噷m�p���`P8=���\��e�����g�I6ē��y��tIY��|����HD�Ge�Qyu�=�ג]�GC����:��C���<G�d@At� q��ԝ�v!�w����3R�6�h\#k�^ےC�-I��g`�� ��dq�%qT3qӕyX]��wտS!��p��L2�r�fЖ�u�����fa�w��d�@�T����``l��CS�����+7.��T��[�lB�Փ�Z�ER����$G�ҡ��fӑ�Ot`��6>�#a�WD����)��f{3ڨE�R��ܳ��u� �9%`-6�+�f��^Y���
G]Y2��ߙ�¯Ƶ����*ABs����ҁ=W|
J¢�:&�w�e����#fko2y}�C�$��8C���f�W"utf��S:�HGW�D؏g\fJ�<=4�K�%I�����L�5�v�gqש��7�����	�W#�AG�+�^�{3�M�~��=��k}�V�����p3^ˡ�V��*���Yi��^M�����k�a��ݓ���fy����ͺ�����5-V�8���J	\~v�w��E�yD�����<���g���>�5��j�D��qSYv'��v�R���#�H����Z �G���Ʈ�-ݵ��"�U>�M�5�P��:����4JF�K	��,��Ψ�����s���qJ�#,2[R��L5���`�� ���0;Ū��Vc���
R�M���&u����!Hky<��ټ�0��Q��7�]��;4�aЬb;�8�GK���Uyձ*�������\ʩV�XU����kХK)��Ʀ� �={��=0.�e{��.dTzk���z�eN5
��o�qңSI��4B4D¬�w����-G�`���eW�nU C=�<*���tkF�FQ�"���Sp�W�l�w���רN��OOR�}�g��V�S��Ѫ#&��J=��}�ƅ��.��3�䇑�
��?�݁���{�,�w��/<}��$:�q#�N�v�m/%������
�]�aL /8�y=���s�3�le����-���RB�E�:��S�wӤ���n��=�x�mO36�g�~[�<�*�WV0�������޽'}&k~ �8�k������yN�3��;Iq��|#rU� ��HygM�mlX����^J�#��3�֒��+~�^_{7Wt�r��^y�B��@���&���J���V�f�b��;[D!�Qp�"�����q�*��V�_4�f���dt-���Ժ�>Ⱥ���k�Q����FG"	.Ը��-�k�]�����T��=v�}����Rh���4���}���TW�#�.5<f�����xn�p�oe��<���r�PT5�+�A���n?D���=ؒ~ �z��]5~���{�:^�My���|�=���X�F^y���v.��WBe����uH\n��`7f�� ����]������]%�y!��ܥ�n�?�S<�P�{�q-��<P�FQ�0�'�!q�)�S5o֩ة^��w����ނ�q�� 3c���y{�W�>��)��=6�ݪv��{j>=���B^���&�U���<Vw>�T���P�r1Z`a���[AWmj�]Pl�w��L�k�Eo^��G��M�)��??Ki��9�B�oU?9�s�B���<�X���^�o�)&��2{ޭ���L�O�s8�7��eO��z��Y���q寶�eu{֒>��{���p<����XZĺ���:��U�̱8r�i�+L��t#��]�"x־��2%�κ��2��ْ�VsD�w�6Z�M�9���{���+S�J�է��y����(��ܹ��(R\U����Eps�qu�䮺=;�,���Z���0i� �ܔ����{��W�ՙ�B�J����ˣ��V�V=�}�E�.� Y7��{W���%pH[ʒ j6��{$����~�]�k����홥��V+ܺ�@Ej3�
�\9$bQ^�??�����v1��t����(�ֳR�����>B��p#��=i#�~?O99��ji^��iN��W��J�u|�S��i^}�X�k�yt�%g�_\ /U�%^<���h�^��k��%6q�M�}[���<靮w��L�����g�$�C��ˡMZ�=��<������o}��^���N����:�p]�� b�UK�,{�}y�]'O���Y�U�~��~s~E����`T���]�����Y��?	�?3T~#�^���ɸޯWy�^�t��|�����J��*��بwO�*z��u���\��6��%�;�2^O��G� o�M�����Ѹ�ǡs�Y�mlޫ�Hgq�z�r�+(x�zg�8���mYB�(����QI:2��:�xFА��+2t����=MlKcQ#N���N��Ӻel;Xv>ۗ}i��5TrV���Uʇ��FK�ʳ�9c�ة^^�.}�5�{~n�E���Q�z���:�se2,QɣD�����-7��c�?a���r�W�����M�#�^8XG�������p@����&��n�VI��#ᣉ�>(��JI㎷m���<�L�b������m-B�$Vz��d��v��F�:��ua63��a���^�}���~�ٳQ�o�N��x���힎�=��e���V�ǻ��"���k<�S7��w���u� �$�i��_{0��7�;��r��~��%%���~u��%�������WA.3IaED�J;|W��z���7�Մq?nA��r���6��!_���ӽԒ=�� �+K1��ud^����(z�c2U��=?P#EL�C����WԹ1��-F.cԑ�{|bߟ�����w���a���AP��%M:���!���3"���7S���z��ǲ��	�e�Z�"�od�2˔���v6XU�(�Q!�%�A��J�[��-�c4e:M���+�W����Gi:V���o��9��+X|���
�
O8�x�K&��fE55�Ach����)��ugj)�ީ�=�|f��Jr�H(��{��}.��O{����.7si{G���(륪MR�p�f|J�o.�Yk���X W�lՂ8%s�ku3p��u�	B�֯s3|��H��zM����뼯:��n��]���tL`�̅^�� Vx�Yj��q��׆��[*oĝ.d;ޯS����Ѩ���F�K�ӆ%5�R��[�|1z`�&{ԏ�Q��1���s2*0��������WL�>�	����O�Ѥon���m{�!P��̈́R�B�&h���P���f�)s�{H�|"�G�	pg�������M��YZ����Wٸ�ud�����^�3ء���/�+��L?##�bk��/ܐ��n�D�b�W�9�^��6�DLW!����4d�����+��'w��u���L49���pE�x��C�r��n67�R�!�\�[�;��ֻ�k���n��|���u訟|��x�
��[ER�zW�l^�����/��`�L'\��B�U���=��.S�M:�-�,�����.�,�b���[{PG����M���G�۲/�c��_���>���Ԟ�R�@��[�T�hb��6v��׏N����++#�4vB��
����RQ�6�3є��h��q��#ph���%�֭"�>����p�$���G��+�j�볱��ܶ�!��j�	g��@}=�Ϗ�M���a[���l�V�2r6��)R�j���s����r��~�M�3֍�o}�|�-���+B;}�W]>��)�Y�Ζבqzf�x�	��	���u���V��Y�5~�6���/�2:�;F�tݥ���+O�o@�K�Ӊ��������?Sۧ����LW���3Mq�͋&�g�zq�y��<�l�����\e�d�j��yV�ܩد�z�-�|�͓4�ޮ�73ﳭN�7Q{�k�mg��]`�7��،�}x�����&9��b�=�KG�+"���;��DK�Ȣ�cb;ff���R�p����� ��8E�R.j��u	�eF����7�+c�U�e�����^�� Qc��\��:��ˆ�^wT�[���Z���V��GC����ʑ�ԢT��
�����.+���W�R�xR�X߽�w�}���,�U�#�>TɎS�D�ٌ���9�~������5����{P�␰���r�'�DFP���M��f/j�z�uN^#��b�α�W\�z�!�t�&�hy=�R^l����G���{o��.��� �c�}���*7�{�$���+�{V_���~Y���+n/";��kiXK�{v��M��������<D���>B$g�i��޽�%!����=b9��#���H݅۶:�|���J��3��6Wg��S~������<;WIq�K8�|Uǲ}�.n:A����jJg�u٠FԢ#�S�S}Tg��A��y�c��`TR�{2����=�m�A�!u��o��Vw�Um�y�h"�Ĳz,�p�O$�����Ѫ��4�����k6k�ڨt�����VG���&�{]��t����;�,/H���1$iq;��FZ�{�Q�;eo<���������^�p4�n��!�%�tyof�ҴE�drYؾ���b����Q�gt'v(�hb�:�E�һ����!r�J�_fr��IDm�[���a�!X�飵.����É�,�}ޏ7���=!��>ˠկ�ۯ;��l���yZB�����Y�ޤwd��=o��i���.��Х��M�7�����ZxR�N�<��<)(a��S}��'�P?=��7sއ�i���Ǭ�GΗC�l{��l��쿽Y��ׂ�F��s���M�eI��簝�(ei�vx����Ș��@f^��O�"}���Y��@iX���ٷ����=�N��n�O,?o�Ңٿ?�X�L�]3�ݫ5zst��DMc��H{w��eE�d������F(]7'G���0���^�������|A���{�	'P6�-+=j��U�lUuE��*ۣ�i]p�^]��d�<�i���z��܊��������^lQxu旻����҆��{	�G�K+����䕅��}�W��o���5Ql��0��ۦ��1����f�|ơyoUa�L��󊺲 i�gQȒ�����N�N�{u����Ud�kH%6(������(^и4��n��Du% ةHsb��̜Gr��ݙ��p6�K��<�ق�JBrL�;v��GyoR �|�;��QW��"��<;W_J	��w�Җp�5��X��'I>��lGِyU9b�zCD��8�h�4g����m6���S\��ڿ�(z�c2U�zh����Y��U����K	�oW!�qV�%4v��+Ku����M��#�C�ղ�׀���.�O^��wwŊ/�g�v5��7xWM���D��5=�p*�B�@��a~P*^��T}WFeB��c�C��[�'��~��{��~ɤ�� Wn�bFs��	�+`!�Ơ/��=w�g|/_����vT^r�Ն#=��2��~{s'�ꝏS�B����\�W����؜f����a�,���s_�]}`�7��lA�D$k�����r�]�M�u�_���s~�!֊*'�\F�̨��Oj�S��WG�S�Y_ԫ*WR��=��ܟ�Lt�U��'ܗs�U5��[���h��D�7�f�}�֯��
5Z��a*Gz��U��يPbRBtW[x늫Ӄ�#����l3IK��+F�Y�W�YV٣XP�~��`"�Vgn�ԶeuZ���Kء8v�h�b���Ĺd|�,�z�D����e[`VӋ����z���ɧ���N����&xVF�pFy�Dl���]z�mO�R#�/�|h/�v�f�}b��ӊg؎t.Ä���L�AtǼ�c��,��`�&Un�b2����3����i�t�������R����ۦ�6]-��r���+�W������>t������V2�3�V�:�a�j�t9���(����%F��;{B���ŝ��ã6���FgD�� i9o�\Q�X;01�]c�`�C��f�g�t 5*�1z'Z�訷��r����QNr��&N��6k1gu�EۄKS)�ܔiꓚ����0�.s{�4՜��&�557�4��w ���e
�i�\�޻�ΐ��+��"�h�Y:ե�a�R��$�Q��өu.�����gU�ems��I|BS�#����lw�;�t�\�Vi{�4����V�Z�xX7�H>S�B��w< �9�l\-�[��H�+�]��Zc��"GMBr塚�Gd�Ad=�ۖ{��/����{s��9YЪ ]�����ܕ�q-�*���p�.j�Va�͇��{�FK�y��,�i�	b3y�shɓ	�oQNS���[�5�"�J�A�դu�ݕye�p��˵@w7.�}~Q??y�e���"���.�gS�*ֲ2p����([�P�h��4ڕ���y��e���[����8�+,m�bm�2�j���ԧo�@�W3�;f�BL�ٚ�l�q���esnT���E;rm+%�n��r�$�n�m���+t����uP��]&u+}}[L9x�(*�9
��
�]�<���)G��}U�,�M��W8����ƻR�k�jt�]���5��VaŤ���mr���E^��m���ft��4�v�
��@��������%f�&=�f�2e=�Ė�eA@�Dm��Gsu��0���Z%�:��u�Yݥ �r�TG9hX���/.uv���Q����[/d3,��}6��>�M�7�U49����󣛰l��H&H��nM�wAvl��Ǝ,��B��˂�\��v���]7�b��_X�E��D��d%�������y]l�e�h�NU,L�Բ��Lavά�",�7��iUׁ�K�7]��BJut�j}{W�X���[����w��
]]!�l�5	�"/IY��e���C�ܳ���ak���	 ���a�g�h ��`�m��@
k�,?.��]k�Ji��rD��2�������Ω�:R��Q�wH�����̶v���7G4�휨q�Ҟ�K6���9aL��2F�eU���B���� ���й�>�|1cG�K�����w���몥/��A q9N��^�� ���w��,��E�q)�}mD�9���3��\��n��J�ĤN�N$�/�7��Qe>lN);�9m�r!E)r!ˆY�ڲ��R�#�8P�)Ê$�=�HQ�q	8^́ G�D�u�c�#���i9'rQ��$s���Q@P�_�G	Q!t��u�u%�Q$q}+N���QQp�ӜRt��k�s��H�l�g�t�����fw�n��890�:K���p�閊7aQq����_>|���������_�k�ne��������t-"E+�gj�.�a�c�U���	�B�h�R'���}��ve�M�>�4z�����ׄ��?���)O�%��ݞ��q�lN6(1m,��<6~��YRs�q>�'+َ���ޮ#�+���7уn����N%��� �yX��=��jdM���B��P����St�>HE:��T,��0��/�Ǐ,��Թ���~���D��oհG�B�'*�.cTz�e>�j/�q�{׮sӛ4�3�c�jlz�a�7��X��R��5�3,�w��Z"�׆tZ7��{ӛ9�Jpl�f�a��<*�?
�؜>��\M�;�h-*	������#�t�HJj�ڼ�M[�"��}gb\��L��U�����}Ѻ���c���+�@�=���h�	5n[�3NZ��m�~�|{[a�u�/N��O+b�Oq�K>�?��q������ k��G�'7>�Uc���<}��J��"=�>����蝗�r������W���J; �� ��7��t��/��pns��\��v��Ƈԥ�p�<=����i�"=2�cU�
�M�6 W�;�]JE��ft��A�y�Щ���=�\������J'qP�%r���V3�\��˒���W&�KPJ��t��o(����5
6d��Y���O� 5��w��P2���7�`gzi���(�E�f��OP�I^�yXղ� �}K_��DVT��D.蚽�7�UWGo:�ԁ��z��>��73z&p$���%{�80�Ֆ2�Z8:H��d9��͎���^��HɄd��ĳ��F
ի�@��:)z��h�>�m=}��Uʑ�8�:�8����j����k���(��tZ�1�{D�gL0#)Ж��Ww��7�O�{��eS��(��eҎs�Z�Rs�%��]���r� =N,3�:��q�O�&A�X�D��M�ٌ���/�蘢:�X�徕�66M�2~]�/[�s��8��L�j���j��!~�l9�:_�����,���QC�F//-�F�`�����kȊ�I�yg[�`�!�s5�7��M�y#��6z5N��xX�V<��l i��������8������Ö�����"�DHF|!}m!5}�{�a�FD�񜙭
����M͊���7�ͨ�mN�|Ν��3݌a�f�5H90�Xr��
�t9�8��}쭩Y�"%�C{#��!�ѱ]|7q������r5�V)�U�bv_Ji��~��9z<�z-⁑�=���[R�;G,h��UQ��7_�q�85u5����� Q���t���Ύ�P��>&7�t�EZe]���j�.��ycʸ�F�B>!��ɺ�m�b�<Z%�J�|�)�@�ɏ)�c�T�Oy��K;��HIJe���w����-�/�6�����
����ߧ����6'=?14�#pE�s7� �֠�I�΀�����zbr7w��0����z�dl˸6�)`��}`��o�-�]HCϴ�Bg��/�q���p�=��Ǒ��s�l�Wl��C(�O1�-�,@�z�϶j���+��EԠ���, �P�x�����;;-:���p/)� ���q���/Ш��b�g��7�U�6$O�����(A3�Y�r�؁������'�g�������yZ�m�ٛ�ն�ބ߇��lXk�D�}�㥚:9�2��ӷ���v��g7�'����^b�̻��-�X�ʭt�ߊx�`�lýtw����@�o����zg1Uf�x��ƇQ���;,P�pp��X5����6��N���rԃ�:,�׽�}i_��{����5X�ۑ�W���B|�ge�>����.opj�(�sz���'���,l;�=45N��+3@�BxK��W}�>�ܽ�r �=��\�
�{jw��5Y�7d��0�f�N%w1`.���ؕ7�s,)�1x9���y����\�ÐG�+��˙p��
���@Lc��vZ�C��dIW�d���>n.P�C%=ߠ:�2[�V��m�	�춵4'(^sM�^�j��tiZ��HHro��-ډ�5vkNޏ��M����7Fh�ނ�6������W��g�UdX��b<�$�>�Do8r k��5��hN'A����1k�l<����.��B؝R&���s�����u�K��7��0H�6�/X�ӣ��Qޖ�߬0ҿ���%�u�,��ߙ��AO�yh�vh�L{C��E���\�ݳ��.63����K����<FD�շH^Ø"o�4����<x�bڟ1Ց$K�F���eS}}��\�,[�A�V��k�ձ>C��KE-s{\�C�|ƿ�NO�6j.6&40�b�r-	�E�lf���|��b�p�6��z�э���~��&�Ĩ�0ô�nׯ}8:{�Nv=3B��R؟`�����(![Ϡ���ڽ\��η�UKҘSW���xX�g�զDnV۪��W�Dze�f\�����3�����ʯ#y>t#_tX�p�T��c�K�j~~k!��g&*Y*��E^�(K�j� g6I���ȳW�ߙ���xO��Յ	vX��n�^}Rƪ�&47J3j�ÁR'�=���B����k4�&�
�h@b�t`��k�ܾ/`(��vIڹZ�w��g�O����h|��K�)�P�oFbR+ޫv�uiTJ�޹�DU�V�ԡ�ɛ�#*h���:4��̧���49���]̫�����D��
|M��f�m"�5�,���ff�06��0�Ls��X鹨t�)��v�K5$�i��k���s�3x��g-��ڲ'6����l쉯u	E�?�O}�y�ڌ�~v�bFٜ|�O��a�7Weq�-�g*�iN\���� �`J�bdM��6Lt��]Dw� �7���wfw,̩^�z{6K�1%�&:id�N����?�m�58"axB"A
���)��M��p�=\\/5��o�S3\����ZRuM}hN���*��k�d(8&a{�W3A�P5�s]���m��o��᨜��<�C�������[�X!_vz�Ʃ�8ؠņ�T_�xl��7Rw�����1F�F^�i�6%ECz�eN�s�kzux#�`'�DV/[��?`av�D��Y�FU�<�i�&�Ȭ���a`����P���ϣǖ}�eϧ�y+��� ��b�}Y�Wq�1��z�@�o��'�X�b�i����	�Z��z�ao:{�Y�m��{���<}>u���!�y�Ց0kW�vٿ@�kޜ9�Jpl�e�#��W�>��ؘ�{A]�7���>�{���s���J����s��ym�q�T}>���d�ͅ?��V����y�L�O����5���s�s�Ĭ
�Z�w�p�KD��g��QP[����oXv)P#��o}��!���9�j�niE���m�q;,��;dT�3��uҰ�)��U�.����r�o0�dXhT'��T�QֈܙȞ�e��M8��"�Y�u��T�}h�	5n[�Uo�{��zY�ϢO��յ,��f��0m��]�1n�<�2b.�;�8;,�^U�u"�'7*fܦ��c>� ��"#ޓf�q���){%ɯ��@����	B�v�"x��)й�E�S�s���%�Tt%&�dz���Í4"����#4�+��	>z�ы�@Ȟ��g���A�<1�HVBξ/"�{��w�!M5��S�DˏL�
�f(�D�`�[�	&oꘗE_��2�*P�P���x^3�Ms
5�o=�%iʏ5K&���|��#�kfb	��I�_1%K��Q��y���k�*~�/������׮��8��}%���j��=�~�pT��jEnzu��B�{����6D�>�+��~�R���X(��nB���~N,3�:��6\Z�}�n�b����^N#^	�Q1/�
11AN,z��J��ll����[u�a:�P������}U'\�4���=�8:Р>z�����Aן4�r����H��_��yPg2'�+�J��5m�yt%jh�w�2�x7˭;SĞ�F�ەj���e�X�.��X�3�T��3�`{&�;&a��Uө�y����C�v��Q�n�d��wwpI��15Vz�b��[Z�SuO'u3�%��q�;����(Ӊf��<��e�y����E�����^�yPm���P?�S �x�_�������6��Љ�T��>�2���![�?C��"$b�1
�b95}��{ ������؅C���79ۓE<*�>���o���|Laǻ9]��X��FXs�~��/�*�tN*>�FemJ�7���x�1����c�W�cƊ�=Dea��7��z��i�~����/�X���� �_�y�p��?7�s�����M��sJ�4T�1��"ϭ�"tUS��B��/Ck����S��Q����1~��:�>���lR��>�a
�X�lH��!�M�!ʪ<8��	[�ss�r�G{z�S����a���!��8QXҽS욁�p��qu(1!��x?��(��b�|���X�?YI˯zϝC��N'YKGC�����73�>D�)���R�7��\,�źm�?{3��4'��?ҫ��t�Խl�Ƭ���N�,k��#����z����H���j��ƅ�[>�><�1�P0T��+B���UZ��<P3Y�J��*�#���AC��ۻ���:q�տFL>{*�R�l3IPI�Z�k�X�B1o5�i�����u׆�!������ү`��]�uo�I\7��j����x=,Ne�K�nnZ�ZÖx�z���A�q��x�Re��mZį'B/9l���j�����q����ua�ٸJ�� G���@�
,
�<,������?H%I�gS��cE�jE8�n0D��O���>`�竼�D���tL����$:�H�9^츇�6�!sx����ԣ��?s��{=���$1��(�����21O|�DJ��\��M�Pڻ�I�e�7/A7~���z���3���f���%ِˬs	�������0�NB22%I�t��|¡|%x*ӛ�+�޷��ox�R���~�c{G��9g�&E���&�PHI	�b,�d?m+�'eMT��]a�)���z�=�
vܪ㫨:2�G�fV��o�>��lMAz�S�'�`,�6}r���mO�q��y��qOQ��v{Z���N�P8F�C��٪^e	ԁܸ�`<�3>R�7�b�O�>`��5�X:�f{���2��2�*N|k"i�����eS�Y�U��_Ib�{AV4|_�Y+1K�K�k��ܖ��M��� lT^N��l[�hO�.�c4��A�oz(͕��GE�{�vC���9�毥�N������=�ޚs�g�6 ?N�R؟`�����rO0�Ϻwj��ޮ���6��(������)x܄���r�tw�W�U⳪�<��9���I�on[���kE�&�Oy;z�X=�ߡ`������R���&ծL�vy��q��7�=<�	V;j�+I�fcN� �k�6_^����V&�ŝl�)����_��g��r�?�y����r�MCrٚ�m�p�զFN�Ӝ�=�{��*U����]_�;��s��+�P/��ep���K��:�Վ\��Y<�LR�W8H��c'��������۩�cf �E8y�a��ۃ�u"�ڞ��Z����(Lҩ0s�c���U��~�F1��hO����t`�+���㗿��b��7Rx�pk�e�� �z��ɾ�Ⱥ���#L�gdM�"��X�k��N��e�sӘ���ߠ^�]NΨۄf�=.�Ɉ<��f���эڌ~ۈ8�`J�bH��BX��@���=yv����e��k��GE��p��j��-��^	��g�Q�>ۈxh��j�D�	�Ժ�2���l>y����yUs��c�����}mI�5��8QAv|Ug��Y
3㢦���yf<:�r�՛-yGt��b{dX��|,׌��V;��N��8ؠ�P�x)��W�t�[l��3��06�&�
踴=J/.��kzux#�g��Ȋ��p{a�|�q�����=]����ua�iS��C��Mת� ���E���|@t��Xu�J x��`i������*�j{v��y�x�]S&���r��nԒ�en�4E�3��6���ES!--��)�.���,ׂ��Vg<�2)q�LTͣ���fx��'X�����-���cD$}��V��ɢ�Oⴻ(:�,WK���~b�Jg����Ul{�-�A�r|����F�ܺ�J��j�F$����}�͚f����D�?_޿_�E;�������i{k�oĘ�^��4/��lC�>sx�E�~����6sf��Ϧi�C��W�W���������t�b���l1�W��&�r0WΆ��=���E{Pu����O�	���;�+_�uF����1"NER�sH�şZ3�M[��ʪܽ�>mc������o��tsLE���fs|��?T��W�(*�ؖ����!��az�H�q�s�)��{��(��������
0Ιb}_O\
���J��ȃ�7׾���,�p�=bԩ��b��/1Қ�4�5�v�T�%��hؓp+��Lh(�u\3;�ͼ�Æс�λ�ںd�u�<������ǡT�Q�?&�J�(HU�A�W*��Q�-m"��Cf�f�[c��}��v��Ϙ챐qZ�G�tm�Q�d�����\Gݪ�&`C`@(�E�O1��`��w��f8�O^ ���z�;�>GEI�w�Kn��w� �yȭ%N�z�[����Xt੿^g���=y�xԠ����ΙXV[.�=�����B ݃�-�͊]�x�m:�1z�1�S������@��n9$��%�u���T�fS������Ht���Z˧x�M&�A�m�O�[�tB`�p�iQ,/��Sv�N�.��Z;r���ꎇT��N���|�*�Nj�*�*�,w}z�!q�yv�r��H�g��+�Ձ���*R;���c����]�ΧsUb�b:�iZ�_Q{8d����1�K4�,`{Rm�|ygR��.ւ$�P묏1-��p��V�d�˃!B	եgm7������d�qm��ˍ�0 6���ao�ʝ;�ݘA����9�*�����3d���#)�'n��G��+-�J��J�*T��AS���wF���d�bF�L�6���`��dEl*���wl�P�v�$�oX�X�K^h�}w\��#.�.S��:��W5�=o*V�j����$�T��46�1-�09�^�_*9ɠnm����[*�J�f��K��aQ�ڏ{���cp�]��ՠsV���L[�^l����e8��+p�m�G��ob	�|v�]#W70��V�$��p����.���4}'x�����}���5����aB�فa�9ziq�g�!V&>�_Y�P��.��ݎ�h��(m	�U��8�87�I�\%F�Tƙ�o�n
y}��:�{g�iG'���(^�!L�X���=D�TVT.h�_[18�6����:l_i���Qу0�j7R����AB�E�,Vy�����g��(V������n�9�-��էA�G9�ŀ�$ͮR��U�急��K�9E�u2hc��кvC8�ts�����[ !/{����l^�C�Pt�X�S�Śþ#�'sxS����(�u-mT����P�����2���y��$�����v&{2�/�ۂ5��C�@�:.}��:T{]*�$<�;��^'W�r���
����Ɇ����U;�;��]�����u���Ԯ]�:M�ږ��Z"��f�D�̸j�W�KT8uA��GUԔ�sƕf^Sb.��ݍ���C#�c@2�εj�{m�K�Î�n.���s_*9��es�ٶ�q�je����7uf%ylCƬ��%+	�o*n`��8�Iu�qr5�
N�#����qɜq5�57Q���Vq-���� �w����kUrc��¦9Y���C.��U��#���CQad��5�����Җ<S9�7���\w��网�c\Xy�0r�wV��3H��7qv�m!�㜺�Dv���nԦu�Mm�v�Z)*}ҝ]u����<Y���呤�d�a�6D74S�Օc��u)nkWN�B�s$�q��)x�	�	�ݲGy����V�*��6�{<;�(�I
�.����k��:��n��u9����P��^gA{c��_l\��Z]{h�!˿��>��wӲ��eD��Eԗ�e'Rts欣�D��"�����l�,/���G%%O�vt\�E�Eύ�pqE^V�|vqq�wE�%6�9$�*�":���;H��{vq'��/#�+8�����w������<�;�׶���<*:8��DB�;��G���$������IrW%$\^ݢ$λ(��p�������ݝ�G\U��u\���,��`�p������K:+�˲��)(�;�2�.��ˈ��\9���˪T�/�i��J�r��O*�o���;%��E���D&I�wSJ�݊Ŏ�-Q����`�%������=�-���h�F�]�o����U���!���*`Ω���OV1�����}%����B�Oh��0}H��S��a_gp�C'�4�1c�N8΋5.N%��.��'
�)ņS�Q�w�и����C�����T�p���u�(K��ְ�����߉�Wxۋ-޹�V��l�ث�ǜ6oY3Jb��1ә�p�s�f�i�X����8mʺn_ r�ex��EߚN����ܥ�"��Lo��7~�#W1l�k�3{4���5���v�����S�[[������ެ��H�v���j�џyRbB��
�Bj�'>�^��Pؗ6�΅#��O�7�}���yw�u�^�+�zv����͌�aɍ]L9��\<l�D�;;�ڕY��o[���Ϸ���8M��C�
���2��g�o���Y�2�=�u�:~�`Ǣ�(�=EnBjӭ�է�d������s�.
£X����nM�oTA���2�!U[�]eJѝ4=�'j'�ȩ�C�����(���}[�ߣ�O�j['�xj!��o�^��T�Tu�>�,�v�e��F�N�h���ubd��L��ԻL��5���K#})[6�^��l��ؗ�&W"F�9���wu��>�n�]��t8�;�����p�ײ+ܑa]V���$��pM/~�F��6�j��
�a��A�d��\p���¾��7Q��m��9�a�lc�ʰ�ԯT�϶j��
1^�(99��)��Wǘ�S���9�kw����q�y�����ӜүnZ�p��1C�#xf�U�0#џ1!����C9V���M��=�ƱЋ�`_�:^�����^�f�������'j5�P,9�����Ov@u4*R��}�1�1�v��fh͙k囃V�V�F��@CY��ts�'�9>�I�����A�|}�=k�\��\�AS���c�+˫} �4�Jt��Tf�ӓq�}>�/mZ�Ɲ��V�@�+�:Le	󕃲�`�� �.o̽u>
�G��g��뮽���& ��:�71Xd'�
1���*±s4T&��Nm]���v\Cr�eO{�S�!zZ*<w؂���9�X�`թ�*�N%w1k�l,46%M���0�]�)ߓp{���9��9מ'�\���^ڄ��9({ըMg��HN'A��d:�ұ���f�Z�`��e~�?%z/׏|m�h�1�
�H���bs��ޝ��ƟNwSbj��'��a�ig�'k�.8
�����)�����=#���7���;�9O����u.��n
,�T�
{yQ�I�W�Q���k?C�`�u��:c����wH`��r�X�J��Yu}������m����ώ�M|�ޭ+p�k�c	U/8��o�6�D!�ך6��7�uR�iT�U���UU�5hX�&��Od�O�Et܏V��~ݳ��.68���$-��~���sWõﻜ��iGk�ȗ�{��*OM��b�z<*Tz�Q��w�ދ�1�Ib�{�
.I���anfO�pu߇t!�mz�����W�Y�0��^�V<)u�k�5����SK,��?dw�����f�+��&���n����^���Ozi��Lб!�n��>���q�9�����&w����|(;�>&��d)����5�񵏄���ȍʧ>'�,9>���S{�[�[��!:���)X�,[�����mˀ]�L�A���g&
�r����(�p4��w���w,EK�&+A��E�b��a���pbлH������\�nT,K32��+�<����'�T�{"�M}�Bz��_?�GD�=���Y{B����r}�q����h�Q1���u4�-�n��x� �dM�"��}I뫎g�i�`�LJ��kϹ��}�!lY,�shbS�t����v� ~ۈ8��*±$�Bi��.������73��c�Z�F���t%v��KmrX����f��˨e�H2��s�ʛ��k�pv]�4G�α���\5���������n(j;�jM|0�*�)<aHp�����=;]����Q\�c��X��]�1�(�Ck�Q�_m��3x���� }*�o����󈭟��+^<p��,��U�}8
�1�v�B��DL+�P��B�*���a����=A�7گ���7SfyK*��":�>����М����U�X\+!F���}�
���J}�ZfX�>�DO)�ǞSFt�d؃�^�U,KVؖĆ7P~��K�����N�O."\���UeJ��N��8��=J2�a��5�:��'�DW.��_�����ǣc�6����L�[�d�7�x�qvPzX7G���~�ǖ|�}�:�J��Yp�D�;?�I#k$O(�0�!�V�Q�&���^������LU�*Y�?x,X�}V�齇��S>�y���7ܽ �yY�����[��x�E�~��#^���͚S�g�,9�-��������;������@�b.ǐ�к��f:M0�g���s�6�!趱��>�F|�K��n�F�}�\�~��kL���l�)��F�"�}h�	5n[�|����ld<mc��۩ߌ�LF�X������ >W�a�y֟�j#b�7w3��dC��q�S�۶�����r.�6K�b��c����2�yoz�[��9t��\����7W�ie��)�cd%E{ՃEw���S�m�y�AS�A�Ӻ�j��r/!�Y.d�U�uv�i�gkfM嗑�N��_w+���l�QȦnh�p��a����Ƈe��3yr�8|+��|>��gxB�'���fG��r}_Ozz���(S��_Zpx��9ߗ;������b3,r(�9���V���v�eM����hؓb,E�Ϡ:1u(t�5��~��5�o:o��
����9�1��mM`�c���tL��}3�T��h5�0+�b�(e��O�o"�V�~����k�*l׬_J<���+Y��Fەj�M�w�|��#�:�f#�`C��]+��}o9�'��yz@�e���fp�A�Ϗ,��V�
k���(�Ϣ�}n�6P��[��e+�g$�+!?�~�n��s�D�<'�h!NX��]��Ò~�X(�˱�	«�ӊ���/�$'lJ}<�=��1��ʌ3�dP3Q4;Y��*=�^[�>�`�zN3.��1��g�7O�.���w� �����(JT��Nܐf�igX��H��F2���n�;%z��Ἠ�l�r}�ڐ�;��{�"�q����#�W1�ю|f�iu��<�+�4X���5��c/��~�y7��7��m���:/}�� ��LB����M_�s�{>��s`�L����w���-�D�l�����t��a��㚴!�J���Q4���]�ޜx�`yy�0���.�2�Qm������)P��O�?s}0���Z�4<8!jK�U�'a�It�]�v� i}��l�h6��&���gx9��<m���ʯ��g��Z�?���\���N@<3;z;+60L91�u0��\<l�D���cğNE�Zys��=s7�����?�P���t6�U�q�eb��7��},�	4�?N����X1�	�U`�NJ��W*�����џ��{>��.>�+��t��� ���4ṝ]�WI����\�nنzp�cy���5�<}[�ߣ���RؑWR��Bf��hbÞR���Wc�a<y��Hp�lc�ʰ�ԯT�{&�h��b�9=�>�p�۞�+f����6_u��/,����4��j_�P��K�o��	bB��?wP�����������/��yL����j�JߖnZc���l���m���Bg�Pjf#� ��7��{|t߽Y���srĉQ�&:d8*}f��՛�R�^��S��w�tǦ��g������?��[��}k~�Ɠ�?/��[��>W�߿o���e��X5���M�;t��X=�"|w�=���M)ȭ�d?��f3�DʵB�_D1�c �>r��!�x�c�J��h�\iߴ�_۬��t.k����\�YQn�%�}p���j�+e�e M�a��'n�+�K*�bm�p���c�nTDKs@-R�/C�����O�mkT�K�7�L�08#�m\�V��hhRZwR�k��ŀ�����ۜ%�̈́�3���)�>�������^�Bɦ�ү:_�w1�>O.`f���:"U�3@�Bk�8���zK^�<:^\uӎ�L����,L�8���=��.�(�Z��U�.���<�[>46%M��s4¡}I���F�`���{B�Ku�T
���+����}Z��4~N�`�s��[^�B^��\z��M�t��C��]�Z�_י�ohu�n׌�oú�NwSbj1z�R��c�K>�64>�LB#���zX�7&ۭ�XdMxR�Z%��z�K nٍ[�f\l`��3;��1iC�-��o%%������U���}�Ȝ��p�������S�G�K�T�3����1����ܯ?_��ݙ����zH`��<�j����`�;���$��,��8�%�?��Z��c�Ѧ�-K�痞&)`>G���y��7n0H[��jܴ��p���v�{�Ϻ{�Ns�L؀�/��p��s[��=���>��ubrC���� �(�Y7m���j�~��d<mc��c�L�@�z����{#�5�ʬ�w��Gt����=Qb��5&��])��:�>�r�o��/�\��x<�L
��@�ה��G�|w��m��X[j@�謁X�b%�Z��E�ӂ+�b�@���(Q}`�i\���[��+qNB�ͩ�Q�A�0kJDq�et��z�ٴ��M�Z�lv�v*�� �Gr�U����$е��o-ݖ�&��-���_UW�Ļ-v�!��q�	���9è�E���a��nZ�H���Uk���7S[S�<����=v�Tb�r&�P��~9\t]]>��R�e�.�����3k&�����=�|bD����F]���|�C�p)�G�HbL�@5�|$K�=uq�oZ9�������%y�؅Yu
<��t�>���ntcv���"/�)]�_(���]t�΋1�g�yEM����:�d"�ㅠ9����w���Tc�m�%8"a)~�å��=#�ܪǐ��s�Sfyɹ�%}�b#�[RTOԄ�Q@�Y��²z���T�eզƤq?�|k��F ��ת�Hc׏<���x�iX��^�u/橱-�Lx�xN�{.�u�s7S����e:�2xl�c�YR��U��b�\Xz�eN�s��oN�#�g��yX7��*����0j�>��-v�#��9��Y�٨��p�֭W��Z��Y��_.\����X�5x������wy�����r ��b?_�(ϓ]�s�z��6i�62f��R��������ŭ����6@#������qL�1WJ�uHR�;kϽ��
��o��ˈ�����߼�>�5)T	��?%wJRΤb��8ԥD9_AJ�8�<���A��J��%k@՛c��t���:y�`gT�$�W7�����	�Iӥ��W���ҏ���U_�j��٤�����C��q@��;+>�X��lD8�x�E�~���φ�lҜ��ϜXT�R���E��G���C_�\vE�DNi�O���4Ñ���nw���=����Q����m�����z�ZI�Y�dz�3xlvUY��`�����FpI�r���Un^�ld7/����o�i�E����]�C���ɱ�ە���(*�غn�;;,�Y�q�^�R,��NK�������9ˬ�Ï�g	��;��8��)�>���l
1_P�)�`�� �7��\��obq�=�,��ޣ�_C�](�����Jq�6Up+�#bM��W�/���@�V�aB�6�^(ێ�,�wu{=��伊��ʸ,8c|马t=
���.=3�yVL������U�H^�݊�������b:xұjI��k=�nTh�V�o~�唀��Qum��]��c�]��A���yI��C�*%9��Lt�8ʃ=�X5�un�5��J5��Xc�����1��S˛���?q1.tO���S�>�����p��u��M�9$%��}��r��^@p+�W���ݪxT1���e׷v�;���5�j�K(���9�Mc!��{M�ߣ�j_-�A��A@ʂ��R������#��C�3h4[Tf�.�����o�<��v�m�)vKei��_Na���F�j1�h�˖�Ẫ�:�}�XP��}���U��A��P�T��a�d���񚉮bb�(�^[�Thm�	�d�:hb�Y��U9y9紗�вi��9޹�	����2-p�Rb�i{�d��i�k�M~�%��R������x���^�����C�ב�q��1;�1W1c���6��,�0mM��P��sK`z�2I���(ߠ��fm��|k=�M��LB������~�Ͻ��y�����ɋŖ�s�*�3/�C�\f����ٝ�����M0�ƅ�Ü������Ή�pָR׻#\EW�+ғ�������#`��W�O~�mK�ߣ+�i���fxI�!�t��/���y��zcڹW��K۞"��w�`d`=�3��kT�x|������k��/Pp>��8��\7a�<-�ޫ!f;�Lץ6�zbr7h���}[�ߣ�O�EKbE�R�ti�~b߽��Q��v{��N#&���b��h8OA�� L�hީ�3횁c��SW��wU�}RO��[����й��X����TX>�nsJ�����b�#Vf��g��G�4h�,K����b}
.���3��"omR���2�a��NWJ��t̵x�����p;$w7�!�edN��c�}�o���2+	�Z��֣�tek{����%_>��M�/$����,�[yJ��x-�]\C&L��2v3�돴�Џ��@q�/q0S�pi�c��p��s�v6��z�9h��S*#%8���uu�H��N��b�]�b����y�9zf����t����o��C|��}�-�n�TJ��хK�A��)v�.|8l�� A;�α�Y�`���EK�R%a�[F�>�j��+��[�2ofIW,
\CkQuB�J��D
��!c��/�t�I�O�̺k0�O+��\���N7�M.�;eg�&ҩt�۸*�	���b��f�]0w���IH� �(b�U)�2�,�I�VQ��̾�7��.D�[FL����G��SD��u��34��n��1����C�Ρ�Q�"��P]�ݝ:��ћ-³
&	�����*nm��eq�]�d�n�䶵�pB^��xʍf)��ѵw�u��=��:�b���ʖe���.gkF�sQ�Qbcu(�,�OINn�ۤ������{���;w&�T�|�0F�絽��c�E�i�h]\��0�=��3l)�,�8J�GK.�L�.[2�&TaH&�..����X��V^h�M��[�q"С�R��22R�GvNT�Չ�۽#BQCv���Qw^�+[�Ŭe�$��\�7fr=aG�uұ�� ��֜�gm֬�`Y. Ἰ��uDE_��׽��zr1�Oj��Э�Z�)�z�E�3b����f����[Z*��$N��g�%k)1�߆�&r��wB�*��Et��r�I\,�#�����ҝ	F�5��Ҹ䣫)BuV�S	�V�e�,.�k���ߐ�U/�^,�|��� 	�2�dR�D�m8�@>���]yr�޳��s�o��g6�C��]ٕ�G@B�i�R���N�R�Fm��!���\�a��[5��0	5�M�ܥ�v���dDؑ����p�깄V�|u��iwW`<d̎Q��v��ag$���6g^q�����ؒ����ꙛ]��eҠ���$��$T�/��nf-6dI�؍p�w/z�%�����ƯO@�D��/0JڔhMͥ�t�Մi���ŻD%�r����pb��B�[�]":�^�LF����9�E�ݡ�t�ЈT��rqݎ�:fʇ3p�{�K�r=GJ<n�1�w�2��
�ǀX�� _^�w��u�y\�xg'I,�7g>�6�>�-�2e%�+����m<�})_<��7n�1��������{#�Wv{�V)�Mg6 sht��3�E`V��Z��wM1�m���ugN})�Z�Po_4��ک����>쉭u�HW3�,����P��(jWZk`3���e�M�f���Ȯ��Q��U�����N�0�1,�5��nsX͍��efNo��o����B���;;��.K�����������wuGgy^���ú��+�;�����;��˴��θ��+�=�y�זw�t��p�<�ӎ�㽷E�I�QEqfQVe�v=�8�w�˲��.,�s��B�(����:m��i�iԑ�S[�����8��p�;�.��^�yQ�k+����W��m�WgVdYݑGBm�:H��s�;C�.����.��:9.;:Ӡ����̣�.�QI�Qq�������+3+(������߿_bGQ��kʛ�ؿ!|�<9]�S�k�Mx3��u箂�Q8d8�R��݆A˭�˛3N�U��gw�����ݪ�R�,@�?ʒ!�Õ�V����u���M�a�Jl�0Xk��L��|;pV�V�_��>��?L�;ڟMȓ�pw�੣6e�Y�5oʭt��S�Y���ګ�ǽ[���;b�����������}k~~��o���[��>z���r��c����C�} �3��U�ߤ�Gu]r�<���S��tԌgE�Q�exB�_DHc�Ŋ�+;.!�*�OÃ��*>���E�p=�<C�yҼ��g�yp���p)���b�k�	��u�j�9V
��f��S]�6u��q/I��aw�@ϒ�S�W0�r���~�V=9U��#�����4�c.����at��x��2�:}~���k��@��P�&�"K��0Z��\+a�޿:��3v)�ǯʧ�\E:ɨLm�"�!Z�^_��ϳ+zv7ƟOt�&���aJ{P!��n<Պ��)_��vA�����.3���p�obhp��H�_����Q�H̸���>�~����A5��� �m���+]"H�7�$m�T��Țb�z/��=t,�g��uO�a�Ә�i�ޮ��acZc��m��Q
�%�vGzWO:-z��������1ļC=n{X�\����b�2���0e��Z�H2�m�Vo ����L!�pM���Ó��D�`|)�mCm��9�[�Y�vzڗ��f�'�h��e<�SsYz���_W�W������=�5�͏G�KB�=�+|��c�`��y�a�P��_����i�����L i���}��c+���9����|$�n�5n^���2�'�ӵ�>���4�>>��ۗZT���gH��N<e���}�.�s�}>W��7m��
j�~�d6ոӝ!Lz=�oB"�N��Noq��U�c�LP��#��S�̛�!p]-���l��ˁ��ԿA��^���vR��G�����˘OԲTdȎ��9u�%���.��v:��������f6��f�:@�Μ�<��f�I��\���'��������׊^����ES۞����/�{�k��s��w�p8�C�s�dM�$S`/���H��W���@Q�~^�<����O������ak��>H�3�:Jv�~��F?m�����C�ʺ�PPH~Rc�Q�Y��xx��_�0g���w�����o-h��u�zxvc ]��V��D(�5���z���座�����R�@Q���V}�b#���$5��8TP\T�´:p������3��߹����nY�9�_�f�l��ےCө�}�
і�݅˰�Q���Y$¥�[q�y'��7�tff��jE�H��N�7�ЛB�8���h��WLI�ƜA�S������._�f�C/1�O9��,��®���}_U}U�mh�yx���n��VU��B�(8O���oyO�׌���W�vz�Ʃ�.�fE?gR�[�]�HS{�f'��^T_�<6~��YR��Uı**01�Q`e��sFs�p��ڂ_��uD�v/I=6���"�W�&�0jdM���
ZX*�pc�~?�G�,�lt'F��:�X�1/yY�Kf�`��#��b���k�N{�\����<62g��5"�>�A{���]aקk��!�9�߻+>�X��lC��Z�s���|���͜٥8G���'z|���&���6�5��v�� @�<1�I��.����y��4L�����g�V&p~�`����u����'�������,!`�ќ�W�s�U�gs��	vx��G�����ա�s��c��|.��_H����E����!��W��n�3��3��]�^~�`�Q}��uXe�A���0g�W���W���
�b��B�v_Yf!�7��DC|L��q�}�swQo����u�K�;	N ʛ��`^|��6"�\F7�y�����lSj/VH��7���n�# ���=`E�k��g_e��K�������z	C��l��U���x�L|�"��$�{��WG�s�ܢ��%r�{�e���31'��'EZL�m�S��(-0�l+�k���P��b���Fj�r��m����������[R7���.G�[W�^U���n��mMg��t:�N����<�&`�D��8�>�n��m���=���(kꛩ��r�2��2+Y��Fەj�M�w�ʨ�x�j���̙������F���Ǖ$xI�A	jn�:]Xv��a+��ո��|'{��>��߳�uu���$*� �=E�������^�]q��U����ƫ8�åG^��� =�H^h�y8��n��D}�� �b�H�q�N��bblp�����}+���mgA��Gt�^�aq�����U�[�7z�1;�q`�S"��Z��٥�b�i���b��Em2jD�^<����;�ޝg/ж_�����;�m)��a�,��G�����,�3���웛����mi���c��B�oa9�f�� �����1���߭����'��Uw�oVt���z�w�܅1�>�6rf����M���t������Vl,9�?.��~�p�����@���'���':_�r}�����'6�D�á�&�����cMt8��҄�b��ױ�Wj���U}�۝�y�=�3J�/^h����E"c�}{ەwc`�-gf�E\��T��g:q�T�������9QV�&�k;H⣩�kzFl��y�Lx:�A��˛��v�����M�,�k�89��$;�;����Ұ��kð0��}_U}UAa}7�l�#�p��g��P2����+j^j�U:^*����A�߈���2b;7z>�|�y���1
T{��Un^��kט��ߨ���}[��}V�D�bD��hӍW��ݻ��.s�Ѝ{�!�����XG8~���lgN&V��꘏d�=B;�)yw�D@ڟB�p}|l�h���WA+�*�ue�9�^�R�!P1~f,v#xf�O�g5��r��;Q^Ɨ�G�G�	y�Q�X?U�7�r��ߖ{-������j�nl�j=�- 9t�jz���8|�~�Q ,�p�'���`ت
�k�yc*��7~)�]��W���:0�q�:�Q���O
u�r���4tP���tstpt���7@�p<�k���}*����bZ2B��`'IN��n���
0��AP�?_DKF/��)9�Q��-��fw35�Z��pc��-�ɼ�I���wPa�C\�S�%Z�s5�
��rBi^�}��G�}��*��і���ɸ�`.�$$h���U0�<��\'!xCbP���7��&�{�|^��=�"��f��I�5┫!�3�ݩ�vma�D�:�L���d�0m3�s:�[����T�9��}��r��FX��^%�Q�C��}Dxx��oQ�N�wC;fN��g���:��⻓��ʴ'�>T�oӃnC�$�:�����|>(�!]�R͙�}c�.ȯ)���>���o��r W�Z��l$'t�-\��O���`�������L�_�W�P�u��]1Z�X~�7>̭���� wSbj0�aO��f,p=@�;��s?qW�U���P���0�pV%e�Kr,z���/��ս�q�\vy*ۗ>���s�$(K�߲Ť�􃚠��G�U�N��Q�4?�i�F�Ȩ=/"���V������r�`[ˇ��-Ǵa�ϟ�!����Ѝ��=9�Qy;�
�-�MRs?pcԧ-���>�*��Cs�"ϝ��%�p��5nZt�8_;O�z�ӝ=�1X�߫7R��#޷o+<�k36 {&cP�b.�pE���nۗ���r��j��|ǖ�y��R��|�̼��T��=���X�p�)K��5��{fܨ�ڗ�cQG�=H����Z��}���5K%F2#���VŰ�#���)�Ϭ�P��ۃ��R3�/}�E
�B.tE��8�_8�/�Xj��ƀ�(Lҩ0C�r&�P��� K������׊\(�A��� �˷K�f�L_��}�7�"�R�:��Zb����<BT��%t�`�[�N�+�X��^TVY��EU��N��ej���+�v��2�T��R͖��.���F����a��of��'IYv�M˦�ޡk��XO)�Eh{\[�n����彩�������`z?|q�mڹC].��	��<g쉣�$Pb�b���9��~z<��\����c����l7N��6̧)N\�n�`~ۈ*r�+#h��P��������}�ŉbXb���Lt�s z�#�8>�+�z���Mϊ��ҁVe��|n�^�6����������Q�j&2�D2:������yO�r��Dw|}mI�5��9�QAp���^-1�)�T}\�R���c;EL+5s,B��p�)�yO��^2߾K+��=���⺗�8}���`����	2�TZ�?X�G�b`�Լu_���Տߊ�4�/x��A���������}����^��O���L���f��f�j/�q:$�F0��~���k�Y���y�_cܞb����n��q�LB[[ �Mv	��?X��L�ܩ��a�ߴ�?x��2}����,~������ωb�x�b=j��3[t��3P�L���fu���L-ٯK���_�\�T᧬!>vc��FWζ�!�sX$�^�_��=�1��ө4��̷6h�SsJQĵ�����c���� \�><9A\d�:�΅��:�깐�osi,����Q���:���3�aL2�7��b�&sj&��XP�u}yFYhǷi+�cP��Y�B^S0/㷿�3t_Ik݉����������,?����	\l�&�t��eU����p�A��ќ�V幅�ED�~�t�W�G��EY�e�i��X_c����1��~5�
�6.�����"}� >q��8n=�y�ў�G���!�Ŝ��Uc�N`�ǀ>� � �yLz~��
��W�(S��&S�U�(��a����%���F���c��u�87%N9-|!�Jq�6Up)��@U�1(�\$Z�m�'ǆ��:Eҫ�gNm���V��}��C�����������$L�y;��]}g��e�q?�0��{�=;�L9+,�Fw�����ߑ��F��lތw�`���F#�������f���1�#�}��1��!T�GKR�*���un���NJ������Q�~���p#�����a����~��g���ɯͿM����}�W��/���/�T98<�
5:���oY��I�Fe����'��b�rFˌ)�2*��Um.,������V���c#�]s�=��P��b�q���7�]�/@n��'S8�S"�
�&+&����� L}��DM��{x���]_�V�bL� Ø�� �AH4��e*Mw�Ix�a&�+���0���`�V��M���]�ն��C��R�����C1X�v{�D�x��N��ܖ��Vf-V9^V�����7��7q�ۡb]�nO�kyp^gW�� ���^�:}�WX��WG�߀Y~����&���jȊ��Ҙϓ�CZ��=���#�y���U��eF���4:`��
��oc��ᙷ���rؐ��1
1�[���M�g�]�岮<5���\�w$dOKrf�Шz�)���]Ӱ����ef�4Ó��r��\���y>���g��E��������=s�+�B"~a���V��h��S4�C��S2q�{M��O���#̈�Kj���5�۞���N���>����/� .�_���r|�:�m�|}܇����nd�P�ꪷ-�c04�r7i^�^��~7����b�0;��&^��NWz7���mU�V�y����U۷	�����͌s�2�-�z�϶j��O�����wGw����¶.����, ��y�Ge�9���j_�*<�P��3m�#_�!��#r��ت؟M�"}@fv�<h��V���1o�v8�/[3q��ۛ�%���V�Oxj6D����n�0��E�M���%��
�]��%�Y�5oʭt����aG�\�n��8��[��k8K�BT�f��*b_j�T�׷��_����������g@����7����=wԴe�����Z�M��f�h<����̭ꐨ���f0z�(���Nf���6*D*��jP{��uҲz�n��2>9U}U��Vf��A8���;�)��O����;h;�8P�*���	�?GA�����Ŕ0L����Y�v8e���o�
M�:�%;��jC8()B�+�����Y���%c�ѻ�Ƽ��{.#�yb�c7�hro:W���)�B���F��T�9�0c�u�����Ǫǐ��t
5v}+�v\Br���7��b��Ҙ�U�.�	]�.����D�l�4;��N��x��c"T��ng��X�y���9����k�r {ӨMx�		��1�^q�)J�/n�k���1~���W�P�u�"�1Z�^_��ϳ+zv<e�H���.8l΄8��+r�^�!t=-�XCY�Xڟe8�n������h��h�{5K��1��d��כ�Q>��B����2�;��1>~��<FD��q��{u�+VD�.=��Ҍ\ԉ��3Ԙ�u�o4�\�)��f��1�X�ߊ��+�=�to�8=9�Qc'bcg��߼�O��,�C�ܽ�����Ⱥ�ӟ1|��)�*jܽ	ڀ� v��^���}8jsޅsy~����:Cr����ݢģ���̉;+0���PV�@�ZI*Ν�K飠��H��U���'-���#F�л�2�Q�\~E�����|��r�w]>��%e�\ ��I<j�c`٥���V�Y�W�00��n<%D!XA�2-լe�9G"�;M�9E-�]m(�N��us���o:�D7(.����x9N�Y�[�՛ܒr1ͮ ����	�9�@GkFm�N
�B��ћ��9+��%Z�������0<�\�\Pͣ.w��i=���8y�|\9G�i���[�oV�\��5�)B�#Xj�� ub��-K�J�w��׵��r�3�r'���/�W�w�T�$@����먦el���Kim(�;�Nra�á�.�V�B�i�4��vw�=���$���Ϟ.��0�"�7�Di=ׇ�	z���)ڜ{+O^˸˶2���5i�0��ϣ�A(q��qmur0dx�u3[nJ�*B5Z����r�{;��̣�p�9��.�L�8��zv���'��2#��TQ�]�]v�·bY��A��T���Xf�N'�|B�],��:+�j%��<��ʤ�>�[z�*�c��{�{�#�DWE&�t�JP����O�}�s9��hB|�wK�1��N�U�sJݓ�����X`Ԣ�:���D��WeA�s��}�D������X���,�]�Bcf�u�/+h�@�MG�;b��v .�T�y�#�|��|��#��_RӼ�Z�j�3"��g��<W���Юb�\�X�NE�YNԫ"�Z�c����7���Qhӝ�0v�ʷ,U��$v_`��:���/R�Тէ�M�h���7[�`����G�[�[H��o��k��Yaej�l	8�}�Hˮ]{�Q��fSeDlt�u�U�٫z,uYֆ�8C
)/a����骦�.kd��2���}�S��`Ý*Yη[�0��ғe��k`�|t6��ִ�Ӓ���S V58�Ρ�!�uu{���{3V��m��n�mw>,��0Rz���%��-��f}������kC�b\�Zj봼}�\�,=1`���.�ng[�@hm�H�D0�ȊV�ו���;X�Q��۶���F�,3��vǮ�HĠ���])�)�Ā��^��Ŭ̐�tJb�Տ&�N]v�۸���n�kE��x6GQ��a��ʈ8�gF *!dy��K�]�\�a��Vo9�{0qJ�[�s�'&qyk��'��hM�-���Q`��ŝ\ˬ�iPE�%�;f��A�	���T�D��5��,��*��n�^�ب��,L-�IPۗr����,6�v�kZ �캄�Q<iH��Kfj���7Y����"��YH���G7���$˲Z鑭�ק��n��
�T�<�dWֳ;�ՖxV�;��u�O%��4ʡjt�L�I㩶�*9��F��q:=�wK;�S���t���zd��#���s�7(ud<�m3l�6v�/��
����V��fYeP��`Yt�D�I�t�Y6�
��*S�3N��q�Q�q���)(�4�(�m�YGY��g6˚��Ҕ[b�㬤�*��������"�K���gGD]��vQuf]�v�,��f�ݕ���v]evE�\]�QIQw��:��m��h��q�Km��q%�dt��RFۺ���8���*��ʜ��,������'�nw%�f��,⃢�\ڬʴ��rڏ��W�`_�g�xh��9���k�������V2�R��^��.�d3�3ɧkȱ�e�e�[}UhA��,�*>��ﾯ��'"�����C��͈�0Н�9�}>W���n_���r� �C�ǽsU[�Z���8b}.�?��L��ۥ�\"b����T�38r���tX����O�ܸ|��������m�α����B��� GN��_0�#�tE89fÅ��,i�cM��ilN��>���#[冧\�ɂ�f�I�Eȓ�'�@����>�+�����t�<{��8��:��z��u��{F.]�w�+�].��	��<g쉠z��Ř��>��{����~��oǇ��H��X��Ә�a�w�6�NR1�}?~~� ;w�(�o|�}'�+L�]j{��On$f����%N�×���;Ӄ�oahV��(�9���>*��� ���W_	1�W!�9��O�11� ���&��7��Y��}�ʇ+;�Du�[Rw�5��7�3�YK��27w�cӺz� �!i�����p���?��bT
�>R/הyM�5�-�,�b�jZ�~�J�zy�,�-@5>S�%!!M�0����UeI��N�J./�=J/挿߇�y�?�b����u���a�l����+���f�g؇Q9��X3�s�%�(����t]�r�ˡ��l���3̸*v#m�wVzU�_��6�-nŔ��6�ή� ����wV�%|�t��	껳��,r�A���`��3SI���YU�����Y��v{}�| �}
��vo%$�ݳ��^8Q��"+>^����]��;��>3{5:n&��F.�h+�K��S���~s�b���o�{�w>�:<��0�D]lC���k�N{�\�ޜ٦��u�)����+=
�>{�?PUԿմ3Bŋ�C~������8���q�U�6���06'�ɖ/�9�\ʿK8G��罹k�X��]����N��BM0�aup��M�OU�ݫ�<�<���t�v�a�8�?��Ku+���s싣�a��њ���X�#޸ȸa�>��ƻ3�,:�2���n2��1�}[R��EQ�7q��ȆGO9�z�[�3��A�v{��
 cN�H��cs�U�S���0%^S�O���"���|z��SWQ��5�wпw�r���6��!/VE�.wQk��ܕ8��S��%��#bJ]��a&;�+�vt{4����aԐ�]u\#&��n��mM`�c���N��zg�iyp�Co���c��_�����=]���s����Y�0䬳��,d%J�1nLj4rn`���E)��mff�S�|��H���l���ާ ੩�ξ�p��ݣ��nCiI�E>�$���N�q�C��ht���5yћ���5ض��NBQ�ﳣ3kcr�;ի���c���[8��v��L`��1.��Ē�>�諭�yvW[~>�����M�c@���Q!�0)�*lT�KS�*���4�G��ِ�ˎ�7���Af8�e_�v�a�
{D����jH�&%	p�ѻ�!����Ƅ��sp�*ӻ^��C�K�VT�ܫ�~N,3�ؼP���)�2LO	11��EujQ/����݂�{f�|��^lﮇAL�f�yc�������8���2,.�p��Y��2g�GM�2���Ҕ�`��{���SJ��ʤ?g�I/u�w��/|����c#юr�����^�Luf��N�i?��L��u��z���Sٛa��Y�ϼ�#>^�!F|߭���:	n�׶�m�J�:�Ľ��<�biʌ��C��\������3�7���c4Ó
I��%���>���l#E�P�9�L-1:�t�z�*_��D��(״�𾜶�X�n�v�b-��]�|X�zeˤ#�:�c��[V�@�gkc��mK��O��Q�|�\F��U����~~�<���&2�Q�x�C�A��N�U[����^�����(���}[�z>EI��}�1�xwf�Q�xYY_��F1�L�i�ɞ!�4�D=o��V%t�d���鮹v��g��<�g�ԍ�b2�Ԡ`��/>�kS�.n�õ-�Xn� �BA���4�s*.()a���2�u�(wp�
	ʾ��"���U�Q�����u�!��~��	F���n!��}!]�6��`9��=3c����I�S�j�=~R2�L�R1��r�M@h4(�+�u,98r�
p.�p�y�E���
����
����o8�XA��>S�h��J�fZj�۪1&l	�$36*P�g��)^X��.�0/[3qෝ@�35�V����V�&��p��*�53}3��"}p%��T8,�z�pj�d9��J��`�cjWi��/l��5�^(�v��@�;�zd�ޑ���'�Ŋ
�"���>����H�8}��>B�X�<��􂣩���%��S��΋0���
�'�mk��q�N��᪢Dw�0��`8�\݄��Ε���a��\(ϙ��T`�\���4b�<U��F�Tw�<�K2�b�Fz�ߥxˈj^�ȅ�g{J�LaW0�s��%�	�g1^M�5�q]��LLcrFD�c�%z����Y��S��WZ�����Va��*��Gs/�ϯ�Û�T��!���Ŏ�[ 5{5:�D��]�[�L�/߇Sfh�3������|q	ꊹ��6��tB���J��vDN���3��#y��0�W:A�:n���j�3Hu���BNN�.j���T
�E��on�EQ�ëu)���޾r�c�x�'�\��ʝco:��sZk&��y�;�"�F�î�8���J�y�qñe�YGa��U}_}�m����hH��Q���9��a�ig�m{%��ʗ�dM
P+D�"ǯ��R��Q8,f�3��ϰ��?�A�wQ��-Xf|��orŖ�dNq���7GU��S���ri.w���9x��^��jc>F��}� �N7�������u���o�b�j��ŋ7��P�1��i�0=��џ1�;@��jϸE������8eM[��ڀ���X�炽"��;ʎW�1�����l�[#ޡ]�zA�s����)^M\(Rs�Jg�U�ͩ�dA�"'�C�ֱd�3�F	ݺs���P��#��S���9HB��b����ԝ�G�f�5��c��nQs�=�������j�x,�&Dt���a�G�H��͇��;���s�]��/��"7�y�#0kxjpj�ra�P�f�I�EȚ=Bz��_�.:y����E�ه����"��������\���<W9��&]�{��~��{�;"k��$\w��f@�5���]�y�k�'�{/�#��sl6��84m��t��ͷJ��qvY�L���0�p'U	�C�?\��jJ�_G�I9��1��P��[u�(��֦+s(n��	环�b�!t}w�T������$9H85;ƪ��⩫���z�R��Eݼ.F{��	��V��5�;cuN<>ڨ_$�ң��������狶W�����t(��G�x�4�X��ns���o �Mϸ���o���S�Uv���Q�MFvTB�
�T"$�B}���'��*��"8����祙�l�Ww4�^��U�1����P]��ϯ�²`:*aY�������>R/׏=�t�oO민4��i�JsNp�V��x�uJRؒi]G��?Xꬩ8=W_)E��]6c}�[��u�<��_��*��gMzp�&�8Q��Ȋ��n����.�ț�^�ό��E��Mx����#����1�#a��Ԣ��~�~������c97�W[�c�z�׬I���|�_�9��ar����p�1�2f���CD�6=~�����t�vV}`�-�LC�f�MRE�[aAs�'�D�@��{��^��^M��>��á�	�¨6$��`�<1�i�"<�יw����7��3�`&o!m��7EQ��dK�d�ͅ.:���LG�EӀ�Mj���Ȥ����k�{�ny�SJ|e�Un^�ld<���67�>�'յ,��J�������w�j���o�e�Kϓ���6n��r�3��T�m�jM�x9�'b�<!���R�ܸNo;�À�[Q�F�oU����7�ڧP�(���
E��>��׉���:5-��Dʙ*]�<�"�@:�#��2��:IQ3�9�t-Φ0�G������{G2�^�n/�W��&n�R�Вq�s�V9O�lc�a�fd%^S�N_�� �^�A�(:�9ӽL��оs½�6D�c�uP~����U�K�;	Nqv� V�{�kY.�2���׽�m���}��G��`ȱF��Y��t���y[SY��C�Nd��U'w�������R�G���i����c?U�HX�J��W���Z#��e�e��	R���Fە��n�te{lo�q�c�#�k'����]�{:�f#�`F&T�Lt�8T��yn�8-n�����iE��'�J;��__j��=�~�pT�33���B�(cZ7��E��Zݰ����"Vx#yj�cr�W���Xe9�����&'���b�z�P���ޞ����J_��0D&M�2B�,qz����a��])�k�j�of�(��h��{�Q� ��Ё0��Qc/-�f�`�	���W\i��C�����ޓJ�f����x�Se��{4����)���
[{O�f��tx�z0y�bF�b|�g�l+��8?($��sI�S��Q;J*]-v|4�YG����u��|S>C"����s�R����n\B�27�����pL{�u����{h�N����ۥ;W��Z�9�rT�z�s�Vm���1E����Y�Xq��=�fX���}U_U�u�ʞ 3�j����ʱ��W�
�
����{)�Y�T��Ze���=u���e����Y���|0Z}5D9��9�8O����fЈ��j\p��0���ر{0h�s�i�2�s0a�t�s�T�?N���5bڷ�C;[9[R��:k�}��#��}q"�w׎�o��~������4�A���pc$ӆ�~UV��ͬ�<��nѽ�gձOwSt�0^��u9�{���k1��
ؘ�$mu��B,+���<p�Hp�lc�ʰ��B���&�{U�y��Hɗ�/�l���
!^�,99��)����^wQ�e�8Ud5.�3+���q�r�d���b�1c��o�U�6$O�����JL��+~Y�1o˱�ŊCs��LK�EG��yl�U��ngo�޷j�*�?H
���4pkiW��2�|�������!��>��Bk���
��Mڀ��g��}�X��3�'�@�Bz��`�q��#�G�=�|��]����L���վ�uI�gBt��S��΋0��R @��<{���7Z�v�{��ǹp��WW(��wy��?$����$��o�"^Z];*Q]�ۣ`M�2���0KBb[��_��WP�L�|A��
����f���p7�����r����<�|re�6���B ���E+'�	S1��"��  ��\�3c�����	�/;.#��<q�0��	97�+�'ss�~�~��V���]7�����h��ޫ8�X���4%	p0m]�����q��n �˽�SJc�����L�z"Ly�Y����2B�sa�s�n	�=3������1��43��oG��w@)f+���Y�Q�:�ep��6ľt��&Tc"��W�P�u�"��R=�_����l��<^?��O6O��4�ɹ�:��ޗ�:DMF|��)�;�}6����ڗ��&�)@��[���O����2���/w����}}�N^�s��%,CA�pbߓ�dNq��m�T���q�ݠ�e��Z�l�^��*T3t/�0q���_e��,S��U�>~X1�������>핟�A�|{7�z졟�W�b�u追"П
���ӟ!|�Ō��8zչ:ݨ.qG+�2�E�	���>�W�?��:�\7�u ���%lO��9�蠅��_�ݷ-�_B��id��k�_��:��0�vIp� �mc��kL�ܪs�OE}aTG���Ô�,tX�"��C���zߵ�;�2�����s�Q���P���ShU�~�x>� �heխ���O(��{A"��w�3�f�d*y��<�s��1d��v���7��{9�{�֙V����I����u���E�:fk�t;�:(I��4� L������}��0��HK����S�y�)��ymK��Y���?*Y*"t�Ƞu�DS���8Ȥ�!Q�����Φ*5����u��g����r`��B�mT���\��z����;�r���0H�=�;�x�p}
�u�nW��.^���O�tL�y`�!���❑4�<z���=�w|�ͱ!��z�_T�}*��9�9�6���@�6̧)N\���Q��N��ٜ�E��~�]�9�l	}B �@Кb����:\z�#�>��oa�
�8Zɡ�GDe#���JY��D��όB�Z"a)B�5��Y��|r���Է.�|�f����x׸{�����	¢��V|�M�f5s,B�����^K���}����]/)���~���=����ݞ���T؜	�,4��g�%�׉���/?o�R#�1EOݢ1���	^��JN�j��R6���Ȋ��p|��1��S"wՎLVMFL��|�n7z�ʿv�0�%�����t^_��+ٗ��φ����ȃ���x�~��7�&~�`b�8��9�Ok*W`��W#�*e:q�B�Lt�ݲ���K��n_@�V�a
@a�XL��M�G���%fV%4��`��eB�Gh��(�p���縢�u�A����qS>9�ԭӵ1�o ������Y�z���@�����N�74u�7�*�qXV[gL�K��;�]u\	5=�"���Ʈ�fj�k�i%��9H���w����:��IM�
y���bb��;�`�ʲl��K���҄V�#&��O���T��E�h�fʿ�V�ҭ�syb8�Z�Nk@�ݥ��V�d��Vofd#��T�BPi���p��j	`Ķ���:��Mk���$����	^2���N�s�D�c��"M�K[��C���tU��R�y�iZ������s�tPiƪ��a�s3���7��ނk�_.�B�-y�P�o�_<��b���F��]h#���1�u0���B�K�%]#}]y��MY� T���nV3��+�*�d	l�dne��g��z-�fk��[B�{(_jl�!����J�˃���/�U2q[X�콑�6� kU!y�=�e��}���jğJ9*"_yaó%:=�TPɏ壒ʾ��f��=�� ���P^i]wwq쩅���؜�)+�ZJ����C+n��L�˚�e�6����r��ZJ9m����N�w$�wՓ"6���� vDA��&��ѩJv'Sǃ��FMVzm=]��ܻ�Ж�,Ǽk���s���l�3�����	>� {/B]]ȝ��K���9�_�������+�:�m�7���;�F�D�2r�ڛ�P��љj]hş\� �g��
�/8`x�n�K�9פs܍�r���(bӽ]B/���Y��9*5	��3�L���Li%fWTz����X3��n4�/�=I<�^��{k�w�D9���Qc��+��tj����7u�`3��PU��n�GN����9��Mb�tN��f����⡣ѯ�KZk$�vo�z7�GqD,���њ2��݅u �<Q�1�dl-_]a�(7�BW��Duv��D(��B���\-���N�f��=��ʮ��e�6�����u�2��F�Z�*AD�r�Z����@敝�rȨ�
�[A ���5�t�:ڊ�n���Z�m�'	9���R`�N�=��g��6w<n-��V�C`5��I��u+��IR'D�˕{x��͜���.�7h�o�ȳ�;��N��v\.��>�B��I�q��_h`��)R�"
�9��&���hv�,<u0�X�T�&<����h����8ァ��n��l�٘Uʾ��[��3�1�0ޱ4+��@��4��m;̈́��h�4�ü���{����Qu���%��@oK��M���u�Us�s��dX�R,�+ ��i)���],�|���[OpR[z�9w�Z熻��'C1�]��]�qs����Y�yWz�����˪�ywq� $GVYSn���,���u��G@Q�q�t��#��+��I�iHu�ڸ�8p��P�ڎ�m�waEqՕd�m����{�ug��f�'o��G|U��fEZQM����;�;���V��D��ΐ�#�㓺��g]��l큕�Cn���,�4�♨����wnrQvu�^u�n켎����J���m�%אw[��m]���GZwY�Ve�g��;-��eۃ;#�{uztu�i�sڶ�I�֣�����T^�xW�Eה"sjû*�w69v�ݖD��,�����mQ��m�yDtۣ��β�.�n� 
U������II��`��]ڶ��
W��݋��1�i<�pm9�x���.��<��k�T/5qr���(n���> }���q_ �ó?�6sf�3_xH��N��a�6�+>�	b�v�U�<�M̵�3wV{e��Gdi��i�[�A��p`�~5�좮��.�bpi�ey�Ԉ�S���ו��Dt���s���{mc��;;3��.��S�/�I^ fPk��H�]�����_{܇�C
���Uj[�Un^�c!�mc��}f0O�j^�h*�����+�ރ�ڎ׾��}�ni�=�D<󸀬/[�����Uc��������g���B�8<�E��;���'w��}��O
���}hA�ױ�w��;����8.t-�r_��a)�ʛk�錃1�w��g��d��W�'\
�p��P2'���7�pH<���򶦵��u*^�L�e{��z3xSL��?����v*&a�����@�f�a�TlY����4oc5��Z��.MkRv쨂�I�.���;��]�{V��u��(I�HISu1����*�\�����|������,/1�nQ=����U�v	��੃`�$Lġ.|�߮��q�'x�(ֻ�٤����E��2NNN�U�sK�]J��ˎ�*�^~5��%y��6�v�޹�w���R]o��z��(���eH<����'�_#܀��2b�{7ੌ7w}Z��۔��β��8V����8��$�S�Mِ��.�g1�U�U��v�������
��
9��nB�*�МXe9�����M_tM��u�˯n����c�:�,y}ҽ��&�+����n��`N�_�ҙ��O}�c�����f���_�+ߪ�2VѤ?U��^Zr�r�ex�����"+�%0@N�F�D�їs�y�r����9�y]�+B��uZ��r�i/�Qˢ�R�xg���;���`�Ċ�ქ,������1��h���E��hF|R�D��a�ޡ�.l�L�Шzǅ76:�v�g`m�@fp_ؽ��Y��E{5�	���V�]Xr���������{�[R�DF��m�R㪔�'\G���oΟ�۾*2�Ҙ~6a�
�#8$��:�r��5��nxT�v<���KX�؊^�K޽g�G�mm�vE���ş[��N�
�ܽ�6�kwi��(���A�Q����]�p��P�s�?��~��W��z,T�$uJ����B,�]E�q�ঃ��P�'af�K���E�tME�
���z�&}�P/��0��&rO�����T_��m�@���[��p�mԇ�4���5��YH+Y�3��y�z��%[�6�XՍcP,���l��'r�u���,��ow�D� ��1j}:�H��4.5�j�����P���=��9�����%���䌃�N��o'.����V��BQ��Gl��!�1~F,v|��Ϫ�I��>�Hfn�&s�5�V��������"��E>R�ޢ���h��k�nm:P�k��_�jf"��O�ĉ�u��ꃂ�-��Z�t-��wI�~������|�f�աU���;P�lý�s"6��x�Ț�@�	�7�l���{n벼x>��C��`YaE�����:��@Rm���)�߅�jF3��g�tL�l��W�p_z���NY�:� P����Q`P��gò�g�(7a8�Ii���'�
 ǜz����m�o{���8��l�v:�̰�O	p=�wޓ�ˈn^�n �]�P3���E"^�S�[:��uh�3��:���U0��l46%���� ¡v8W��]c�@޽����9�ɍwU�n�g�Y�YR"i�v9���1W1ap��f�j�P���]�+T��/����G�(�z�z1���+xD��=�]8;�15��8��1��FϮ\��p��D��Ny]m�uOfh1��g����*�=g�zW�f5��F�A���LC���1hO�9��S�ڈ�R�Ҏ�����d@�����dF'9S���Ͻ�������^镝0Z��<P@��5vn����xes���*m�r�׮�wgٗ�ieL�pu-�D��G.�)İ�n���gf<3i���G!=�gV9�L��5v��9�5��:�P�2&S�����촰������]��7��7��pb�J��7�#����8��M�Y{?z�>x`p��~���XuƟ�9�.�cM��uФ�n�չa`3�JE-��馎T��87~�����=�8Ϧk��a�>�������(!`�gݞ"(�O�|�g���j�~k!��p2Mi��N�Ӝ'��*���8��!yuyUT��Akz����n�!x�/M�V)p4�Կ}����U,�2#��NE0�#�{�G�2��>��:ȥ�{�d�q��=	�ۃ���dFg��Ω�*n�,ک1�EȚ=Byvճw1�U�͟�l{�?��ȸW
q�/���{F.^��x�s].��	�5��S�rr�_U�O��;ޤ5�DפHc`@u�H��r��9��1F����ѶgBt��ˮ��Օ�Ow�&N�:@����w�	�߫��>�C4%�*w��q~���Nw��=V��*��D�f��U�� ��[7���M������{ƀ�}��Em/�/�wǙ��I����P|3L�F�C�r��B��b7�K0;�\�	DM��6d3��.�p��8����ᓱ��)��+U҄
���:��f_9��D������(ɲ�+/7*ɛyemD"��FtK��Y�Cm����:;۝UtnIӿ½LD�[�+�OԄ�QAv Ug�
�Q�詅f�f�x"�jC \�ց�^:�Y�5�i��.���4�B]������N(1��hg�՟�jQ�b`� �v��N�[���$vq���E��[	΋5�:��8Q��"+��=�� ]��7�����}=2�������A~P���`���EŐ��W��+�/�3��#Ûyuu�>~�@p�����&j�kk��(_n��%��O���]W[B��P��Q�_>�o:{�Y��X��Or��Kw�Hc�
�a苆_^�-�׽;�J}��:��W�>��؜���{�4a~��=�]{�.���\7:j��kn����g�v%�F�谩�LҘ�o�nCUY��4����ʜ�u��"���FrM[���*�r��ld<���66�2�೰~���~��i	q�7����؇�B�+�q����
���ԋ'7>UX�?}�<}��J��<�h�Q��LO��I�����m�`W��1*:���ެ�R�\���q�pZ�v���g���S?-7ܨ�`��ޮ�Z������Z˽NV���� �����Uuu�wh[��e��=�s�J��6v��'}����+���f���<�Ί߶��7���"�ϓt]q�=p�3S�uա��nn]`P�Vo����$��Ӊ��C8���	��O�W�*�6$؁^��@tb�J*}F�yW��F!�mMi
�����bh�9��ԁ��`?Ss�Ϧv
�����D���:*a�Ygz��B���X�9��MI>�w�ܳˣ|�0��V�oq��ލ��a n}�P���"4���S��KyB5��[U�:�^Z���z��(��tU�v	��੃f�D��٫���j���dm#�x=���J9ά�R|��%v7!hU��ņp'X��6\`S���C�g���M�X����Ŋؘ�����x}f���Z�2~E_��W�`��Pc�H�OP��s�9�D����B�����΍�Q�d�����9)W��Yy�Ja{�9ۋ.<���)��33�"�1�����j��Oìd�B�1^�@����|c�3U��~QԽ���/�e�$?��ὦ#�j�ޡ�.lɚШz�)����߇�<9��e��or��+��mRLh]LE����͜�
��у�[R�hDO��C`3=����S�I���Su�¥-Y�ӈyE���S��Ko�A$�7e`B�·f6V^>	Ĳ����ַ]�X�+
'(
5 ��{��3r��.���s�A�N�rF�q��mVU�״/�R�t��p���ܒ���-4�*�s�K�'�S�>O�`�Q*���wu�r	�x��^��6fگ��
�30e��K�r����@��F3����f/՟q��C�$^��m���6'#��S��%�xo\AԠ�	4�S4�lb<��n�nǧ��U9�l��.�?���, ߣ�O�j[/����i�� �UG�ǎ��p��(��n%*���ɞ�ގ�j#���a�~�z�϶j��
a��_�(99��)������*x����f�x���(�:���k#���*/�Ŏϑ�3s&$ϤO�����JL��)��Sc��M^v�k�"��C<�じ��7�����'|�l�@�ML�a�O���>���\}���3Ӎ�����I7
�e�1Ǖ�,V�F�O�lýǝ�s���8PwDP/����JB�����
����N�v}�k��~�uI�g~N�����5#>gE�[��^�]���y���m���XB��"��]	򕃲�`�� �.opj�(�sa`�����x9�Y��=47��	V<�ʐ^m�G�R����d�A�{ ����׾�1{��f�p�6Z�Ze���W%mAY��ْZrb�7�N�`w�N�t[{�u�x�e�5 ��Nf��f���:u$Ǣ�L�����}�\����:�l.�I�:�)'Z�U�'�ۛ�w�{,�8o�.�,�K��a�{�J�g�$���g�����<�>��|��_�����t��
Ep�)�X��:���w�S/1���|���8�ƺ>D�hIN�e���¶W�P�u�
��b�H��T{�j���W[���}�����Z�c|�t�ú�Q���?XcY�X����2?g��!��gP���zk+�f�����'��^��slƽ�q��.�3�ʘ���pb���o`I�us��w~���'إ.3����Ց5����R�~�г1��˃��-Ǌ�ᯟ�r�&̥ǥ��w���\��~7�E��nN��v
Bw�]�iϐ�>vb������yVw�;�ܲa��a;Pg����+�}9�ޚs��LՉ�`T�'�A8}�-�P���~�W=��#s�|UR����r���xk�Zdd��9��\E_�N3?>��}5=��x�����ŵ�U=�>�r�h/-�~�Y<�LR�Q#�~�"�؝�T�E�ci䡏�٢p�j�P��+��Z��b���~]��b�rF��&47J3j��9"~�Fk:	�n9y�������R��1Vܽ,�+	.U��{��&��/��I�%�n	�k���dtig"��Q@�\�P���
yh�[4���[M��{iQȱ3�p���d����+���!�����M�j�����s�Y�J��0��/SlM��_m��'��U�hZ���/`�	<W9��&]��p(�.�"����G��x���7�����$&�����N}}y��(�z��@Ϛ6̱�@��sj����7�1�Ҝ�y�j0/m����?:W*+�.� i�/p���ѻW1�WH\L��3�H�,�p�n|�*���]��m�,U�&��DH!P��p��Ǯ�����B������}��f��>{�"�ZRt5��8
��Y���VB��f�\��@��|��]x�=ݚ{�V�co'>��S��`�c�=�ভ�:�Pb�meB�?oUeI�������o��G_��ؗ��\XC����`��f��G�G(�O<��^��~���x�D�(F�/�E�_�
���j�&�`l��G��ph�t�+��ٗ��ϴ��g6� ��!�S�GM�}���[o�YR�������43K�;���>uʘWRܡ��Q�_>��g@o{+>FG\9�#�^�J9'�������VD8��^9�lߠb5�N�٥;��a���
��"�6'�DfH^P���TS�p���8>.!Ъ�ǘ�h�bʛ}�I�:h�Q�x@4�����e�X�����<�gG��R>�����=[��3R�%Nc#�S&խ]o,�ұC��|ᵉgs,)ӯ;d���kM7L�ީ[#5�@|�7,.��+<;w#��D�]�}�g{�%+Q�U �aup��~6��8ݪ>�Fؗ7��5��:��
��P�2�2gW{�[���Eנ=B���&��sભ��ld<�q�����O�jZ>�1~�_fת��W�ky;����;�9�dB��/[�۶�Lے�P��}�&���Š��c=���z��:��~~������	b�v}}dA�z�1N���,l��8Uk�����E,�g�*t�����K��Y�W�*ѱ&�
�T)��Ŋ���p��ͼ����Χ����ã�'.ڃ-t�}c�����3�9���Ss1��D���;SJϬ��.JR�&2�Z���&�0����n�iʍ~~�����@^�@�"���G�E5 �����7Z�^qSf_eA��>x5�un��C�ѥ�sE�������S��$J1�d;����}�;ϔ�}خ�юrna�>K�܄���8��9�
8d�?W10�2=iyH��r{��J#]�����������}+�̓�8 ͮ���c�N�w�Fe*�TH{�璫�܏��}`Sښ���&I��Q�#!�U��3��.��f�,�'Y��Z��ng$���[���x^3R�r�u�=�pܼ�ɀ�s�E��g��{X'W-���3'NkV����${���Sy �l���J��m3�P��G)ݞ�+v�1(3U��Z�9N�gD�J.��� j���:u����F�<8	�78};���X��]��;;f����]�KﲟeB�r�h��d�����ޖ�Ԩ��u��奺bmw!KZ��>4]2�S����;L6�S�a�����E*�������-��F�$�*R����wU��&+�j ��Z0�:�]6�S^�����Fh���)��-4=���p,��]6u����n�t76��Z[���l>��_	wl5� ��j��#Wu�C7y�JO��f����d��ށ�b���e=ʎ9�i���&#��U�A"R4�Ǝ���t�IX�M�x�k9�A��E�����BV�
�X�+VP2}�T9�j����3��v���q!�ؕ�r�惟"Ob�n����1�.��-�ʣ|���Y��ǽW6�<�yV�Aq<��V��\o�2n�D��b�X"�p���ìIB�N�"�N�}�-�'��r�����x���K�5{�3���e�V��uEsAO���ԱY|U��<��&��K�����t�X��������C���/�p�	.V,�4q���si�}�b��N꾗D��4��D��ua���f��L�u���q(��q�M�6O�a�D�ty,-��5�M̗2��D�xˏH�_!QT{�f*܈틗�q���3����������+C8���ur�PK�Ag��^`�te]�������^F+xKZ�N���B��S��Zoi
r�u��W�>Ύ@���[��6���l��y٧���Bۭ��H>F�GvT4�Zg�G��ʼ|�ɼ��o@�m<�"��\H���cCX#��1���U�u.)�� �d"������glV�'k�eHs�/!�}��wRv�hJ����D=ۯ�cUܔ�+�I�D+p5�lԘb��3�&�7�w��+R<�����t�Ӧ5<��X�E���}X��!�Vٳ�mk�ʙ쓷WnQʗ����k��]wg\��hm�QzE3s�J�x.��
`�a��Py6�`e�K�u�	�zd#FZ�-��5i<�M��H����Δ+���Vڕ�h�ZhV���_Hmd���Y:�,ԑ8�=`�O�k���Z��.�LӾ���+Ȗ(0��!���ܝ���S��R��4j�ՔF�!գ�_Qn7['O����s4]]�t��oSŎ����!6Q�SL��ur��V;3d�t�����켾�}�\լ��d\�z���u�"��x��hЭs,���6QYκ�Eƶ���5�U�ojT$(����)7p9W�t���jTy{7-�ܤb�Nc��hp�c����T����*#(��u�gv�\�È��K���N���:�/[Qd�A^���8�;�����Iv[j����+�����ˢ��yo7Y֝FD�ge�j����m�y�7{j�*;��¼謎���7l�i��jmI�����vv�˭;���Y��3��j��W�u�\u�vfy���n�-4�<��yy�^���]���m�a��n�n�:��-+2�����q�YE��gy�\VQ�V������efrgfLMYefgD�.¸�m^i�m�mۼ���Fٵ���U���IKh�+��y��i�]����\]y�E&��*Ҧ�g��q�ڳ��:mѶ��l��ػ(ù{^��f������˴�γ��mZz���}o�/#K�-a�NL4k=Q�,����/��
���y��l��Z�\�����)}�v����y���'X֢�$��W�/c6s|=^�J���T���\ζ���*(p�1�tܾ/�vW�7����*����sOV��wN,�jસ��0�;�!J�,l�k� ����3�W1^�_]m�57y_Y]/�r͍[[/������s�D���(�m����'�[���rb�phT=c�lv�U=w��s��簮S�^���a����͌&�rcWSp?P�m��OG���emJp��x���	�����k?�O�?�E[���ϫ�7��+���b�~.���5���#>g���S휪���sL���cڞc��5b�}J��nE�s�qX>�0I�΅Un^��������b�h�tY�u)g�"��3�G賮�~���躖ċ�!��qE��n��v������d�EP�ͬ�-�y���͌��
+�X��}�P,p��F�R��n�
W�T2��� VS����{�G���C���Nh���j_�*<�P��}6EQ�3bD����B	�/hK���;��������k�i��>���^�f�5m�7�څ�5�P-�L�p���~�We{�:���},�~���+qa�qo#r���Ȑ^��Q��F.Aó���V�_d����e�V�' Ք�Xe3����fo%�z��:^��yx�X��썶����K�J�����초�j��-�.�B���ʷ���͋���v��s��(��B�UNu�R����Uk�n��(����?M��tN6h���iLA�t�sc{79�� C�*:�	0������r���<V\ksO��Rm�ߓ��c~�MHy�����>���?{w����Ή�� `B����Q�������q�����-M�J.S����gk{�Jb����0��F��b�h�M�Pڻ�I�츆��7j�W��8��#�E������at�Ws�[+�X>.��W��s�#S��S+E=��y��ۭ���Ǒ�|� {ӬMx�		��"�J�,.������B"@��d�n���b=���OOPTd=�q�ٕ�;2�>��&��S
S�pi`��3�g5h�+3�W��DY�M�܇�/�
p�t���٪_�1�{2����}$yS��pbО#"n�ѯ4�5�����?�L~���]T�7����N/�]3�~����.`�Ÿ�T;%�=q~Ŗ���Ň�퇟�<�Դx�k} )�ӛ5��0�r-	���7�»?.����fr��ވ���.�ʑFG�b�R��f�xmw-R�(޺*��oc��F5
�y��:_c��y�D1z���{�c�]���`lu��4 �v��^��J�2M��i��2N�L���2ب���-��t����vA��#����7����}Ux�ܧ���?��kҿ�ڀ��v3��}8:{�Nv=3�bC�د
lOh�����u9���]�";I�q݄00�Ϭ%v�� �����CϛX�A�2<'v��}�z,)��G��{1�׃y�-�P.�V���ً�{M���4�ԿG�Y��:}��|!44���½N)9��{�c.�����D�~͇	vX��.�R3���\�nT'�jz:��ٻ> �E�5s3�h���P�:D�Ȝp+�P%�E��p_^9z-^�Q�.^���O�k�e�^�v�E{Gq�.���Α�XvD��#`+�k��N����1F��o:O�K2�R���g\\�{����ό���ntcv���[U��P��E���/�F���4��*��jOƽ~�[��g�}k-���ߊ�����m�,�*�
�T"R&��)�4��ۦv�E����W�p�5\�'vX��2��Dq�fx��DJE�
����Y
3�����L�pDW�R��)w�4���.��Ol�7��S�5�-�,�wg�:�j���,4��?���(����OG���`�1<]t�>��ı�+�ۦRYIP��5������	�������0)�6�R�c�(�����#W��j
�T9u-c�8�s����4�r�j�SB�-]�"����2�f��X��|�3��}�i�iy(]ʻJ�����r�����]����>�7<'���(���nv�oN�m��O<��^����c|��%����w�s�ʈ4����~B�ڭ
ġ�o��~�a�Q̿��i�����w�I�����=[7}5�t=o�o�`	.�9�s輚f�������϶��:�t��ϭ���sޞ��r��a�'ٯ����[�Z�sO�`/��zw輚S�ϦXr=�p�+,Q (|Ə��I{��g�~R�0W�Ϥ�F|]\7;�j��kl��֪����~v(u���bN�9�U~���t��,1g֌�jܷ>
�ܽf�Cm[��G�cǋ��V�,F{��g7�L��O��}?PU�t��v}�dC�+�׭ԋ'7*fܦ��c�L'b6uzVE1�?~��B�?_,�q}=bl
a����N;>�":��Y�S���X^��ΑU'ˢ��1mv��c<��QA)a�63y�l@�@_91�=PQǆ�A�Sx��;�b�����__�����y�m)��t:�	�2������������嗻�~�}�[���=�������5��߽�ե�֫�����؋[]:��3�_n-2�eI�73i�Y�ڽ�٫z���;��8:��m~�G�����v�m���w�8rgS�[x��*�ǋo���.^U�+4ٕ�lL{��P�������B�jl�g7��jc��h�擌v~�B�OK�u^g�unTh�V�n�}��˸�`[3��T���*.�����{���/�_�1��s�
{,�ոD�?�OC����6^׃�����*
��A\n9���&���,O�k�+�bǮ�q�9QAѯ%��.��-U��'��6��=O�ɪc1w�1.A�gDȡ騚Q��
�_�-���`�l�B�]�/Cw�c3������7�jc��TZ�2��p��y�.f��Q_F2���o��씉����ޡ</�ϻ�lY<�)�w�a��b8��_�=� 3{4��d�}�[�.���P�5��̝^���}�S�:�"����Foa�RbF|�LB���[��~���C����hJ�Rɼ�=�|sw�u��]�^���N@7~����Y��L90�Xr��\<����Q��=s�+�gD������`�S?M��P��EX궓��mЎ�s,�C��f`��K�r����~��B�h��O�ǵ���G[�6f���VԬ�k�6%��]Dg�]71�o\A���1�i�s��ܸ	E!.����^^�@��x�̛��#VD�����s��I깰Ұ6��]���t�g�{@��3���F-�6mX͘r<�jc��T��ލp�b�"�[�553oF�O3fR�I���V�7��M�"v>D���va]/��R����5����n^��V����5u���P��z,T�$X�!曈B,+��%���3f,*����Ch��9�a�3c�U�����3P/��A�+�b�'�)�W5��d,��>�=Z�_�l\c�����Zs�U�5/�B�c�����s%�Ux/>���@�h)������}P߻��:{5�~��nK���5[3Q�j�nm:P�]����ET�y�k��9�)7��;�<�p+aX��5�^���^
�zF��@��Э�y�-�����3=�2�q��ƺo��~�/�'�L+��1t8Y��; �X5���	�I�gS��a���DQ�m��v�?���*�T ?DW�u��>r���g�(7ai�HU~��ԭ��ey�]S�'�
3��s�)��+3@�Bk�85]�=uܰ��n
����5�=�q���sֱ�niLw�\��ϒ����V��hlJ����h0�]�8W���o����Ayvz�S\���^ڄɸ�}��&��		NC���懶����rvP��@g�B�I��י�d�$�#f�V�(�b#z�������bnYUN\�xO���ku��9�t���ͬ��i�/���`>���U�l	8x!��p��������u'-�Y���a���ьe�lo&���P	6�)}@��b-[���~5�Oyd�.����u�
5�-��ܭ���}=�ؚ��L)���1���E��d�F*��UQ��t�?��O=������Z%��z�K fٍ[ٗ�.��>T�<�?n[��[�����YQ}��A�_^�h�z�TW�_��|.���g;�n��qb�x�F�0���^��=���Cb�/�a�X}�w�o�8�6j/읉�aVŹ��A��s�"� e��o�͘�����f_!�~�a�b�)�r�v�8��<�׾��٧93B�"��>�,���������j&g�������}vܵ_Cr؃YkkL��t�8OD|��Z�%�>3;���u�p���W�+ƾ�}��|=9e�+�d,�X�4`���^A�e�x=�R*W���R��&(h5�LQ�F���v�šv:������r`�J�G�n����6#ΪL0:E���=�����H�������`(���7@I⹜��^��߮w4��М�Ҝ��s�?P�
vDפĘL���C�;}y����\{��c|�vefD�"��w���Re�ڸ����i�Г��݅zhS��f�[�x\+p��5/��b��o�r�p�y�3}�=w��K'S�n�a�G�t�a$B�O�Lz��U��(y']�2	Ƹs�Ur�;��e��������6l���7d�r���ݨ���qV��j� țQST�K����E`�ӕ�g�KU�[;ʲv��ߙ]�����;���`zy]=�@O����D�/�W���ї�7�W�=�{u�WO���+;�Du�[Rt5��8
���ϗ	�Q㢦�|]TL�䄳:���4#`?��R/�^<�f�e�%��g�:�j���WQ��Ll��#:�]��{Ϙ�#��2�*V꿢H���E���nt��ԍ��D�Ȋ��p�1���~V"��{��{�L�[�r(*����
k�
��G�_���yMb�<�t�`ߺ|OX������>������	'�G��Y�?_�6'].�8=׮sӛ4��c&k�Fƈjg�_Y���ޯ9k��xz͟fﶻ��s��<���iq�S�kW�tf�>F���6sf������a��a���n��*��_���]a��T4�cWX#+�`�L9�up��i��~��'%�pN6�睷*l�1������>�]�Unb=�Eр�H���#<$չn|U�lиg���_�&�>��A�x�#ۣ������&��
�w�KVT�����̏F&�f��b�-h9�쇮�U:�&��1l�&>!��ou�k$�U�
��P�B��e�s��Kr1�LU�T]M���W����j�A!��C��,�j��w[c)�6ܷf���s�hM�l�y��%��h�ر�7q�_Y�� >^�R/�q�s�V?�=]q�����̜����:���@1�W���W�� V�a��%
q�.���޳�~\Ȍ〻��kp�Ou������PFsҋsa)梁}W�6$��+��ы(𮫆g�{莛�O�D{}��/q���������v��v:N'D�9���Ss1��&0h/���[�&K���x�(������^����+Y��Fەj�M���Բ�#�ճ1�=�dT:��S����
�1�uM��K3�*��cunQ=���a߅����O�*��Jx�J�npCh9�e@�6�8Q~���;�ʇ'��Gcr�*�МXd��\ϑ�a>��)*#�MC�#eF:&E5\(��x:Q�WO�u��N3k�q��ƺ��G�*�]bw�{�Q}�jaCҙ��Z�pPi�2�/�i�u[(��?r2��a��ઃ'kM�-�i"7���"(�ja:�Bj�,l�k�6*6igXɚ�T.�b� j�;�h�x�r�_���3���3�[�*��_J��^�><��L��K'�>E�C�w��G��M���N:�wm`;t�u�V�J���\Jbׄ���������3GX�/!f��4im<��ܭ
`��1���d�=m�z❆h�O���s�Z�Kޗ���v��FySbF�b`o��`m_�p{���z�Ĺ�92�yô�!˫�D��=ⶸ{�{E�o��l����fv���͌�Lo˦�r�"��l�D���&�LxZ��7�e�~<f-���dIhh���.б��W����]���Q�҆��͞��EBr񁽾�g&]��A�(n���p#����M�u�n�ݕO�eR��
8Uq�}�-z�!�ln����1;^�uq]�문�lf��Y}��V��6� ͻl���o�ܕ����A�:��=�x��)M����^O�f�t�m���@�G��k��4���N}vr�ݴI�Pk�#���+IU��>o53'��	�#�n`@~�{���jʬ�q�����ޡ-�����+�Xf}ŗ��u���>�4��D�5���_�ؽ�&��w��_@�_Hm_�h�x�x��b�}c�N�~���2��$�7b�;��z�:�SM_X뵏���{*���TY��A�y	�H��q�@��I���Q�:(I�w8�M�wt��6���N�c�3Q	��� X�0ފԒ�6c�<���\V,T��uܫ���ޕ6�H� -j婻2��!{����[�����Χf��ck��x��T}.vEns���K���tb�4#�W���}=ܲ�z�9�0oi��y��'��"�oy�
�<�CڇO
�)4�YtVc����a"�mMЄ��T�b�\�����2���{�7�fuJӮ�ۛ��:�_���¦�X�3{����s�>���H;IC�v��c�>M	{(D^�1[���L���zk�[w+Ft�ۛm�9s{��I^޸hZW�ee=Қ9�Z�P��*����g9�S#�bL��z�S��]=�ض��-�,�r-�x�^Y�2��V��x,��&tu	ߒ�)­Mu�0�����.:˼ �F$8��2�f�.������aK�V�9�m����l��Uk�����F��2Qje�Wt�	���m�N��ɻ����F��,�	�Mҫk�SϺ4)fǓ��b��ԏ��r���9�>��r�w9F� 񹎒���5�<�����Lk;��;��%~�ߗ��QoJ�S�Wq���<�t�s�4����8��qL�2�����W��:Xx	��# ��� ^��@�t̔)AQ+����0]k��rt�^�ʴa�݆��9>�d��û7��>/�8���N�c��_5�P�j�om�d��t\�c�ܳ�YqtF3C9��p㬩]F�
����Cw�!�-��äA�F0�폕��;U�@p��iɗ��l�ԏdY\j}��\�r�:0�Z�K���J���-kt���	���m�*�nA��L�'�4ۉ���8㡖'<���ʄ�W���p������u@`o\�{>��N��U>=*�hȪ��V�pVrҕ��ɝ�]��d��q�����`�F�7��y[��7e=wpM�L�m*�5�e��P�
�d(M7)ҹ�����׍_9I>;�>=�u=��ӿ��;�.�I�:AW�#˗@���h+�y�Y����=�PA41�b��.\I�C��	k	r6=�-��_u�B�;��%:�m��[�Q��k���q@ъ��$�����ev�:���tz��[�ӳEŪ�H����q�x�J��ř��'I� �����\Ђڝ;�f��=�{y
�2s�չ�q�����T��E1���;]H�l\o.�M����Zۦ:�>�����ˈ���U�:���6l�l&!��L�{0�&�h�*�ז:��]Q���:��v�)ճW���p&}wh�p��t��";�[O�9����\.]s�]��	�l����!�[{Bu;;I)����ZB�36ǻY���� ��S�Ph�����e�w���O��mԕ��R��{%Y��EGE�qu�I�a�ee�YV�����v<�,��wdR�wgeef\�m�α��3sj���v���mݜvuyu���� ���t��ٶ��9�e燶�p��+N"+��fu�D�g�݋������^��;�����.:���u�V�dۥ��Ā\\mn8�J���������H��E>n�legv=��m�F�3����³����l��Pu7ǎ�v݅��Y�vV'W���;�C��|��fr]��XpQ��j��6՛,w�rYY-�c�N쳓����r)36��Qva�gIEGڳ*���{ p��8ӲĎ�O����;��ɷQ�1�vgk����eA��7]��d^��9(��l_�h�}�zI9�8`Ҝ<�擊nSz�|B��Y�ɱ�A��k����[(��::�at�]6�31��t�ܳ3�~鋫�݌�:�����W�kBǂ�)0<֏X~�����X�x7D�!������&OԄ+�=e���\��Z!yT`!D���jϐ�V��mv�:G�W��	��;k|�/>Jв�z�J�����%{�R��*��P�Y��vt�	���Y/U���k��&�)�6Ŵ������<2��>���&gν6��!Ņ,!�W[��_��^]͉��j�q�\<�k�S�u��bb���u�����C~�zӫ��������L/n(�y:mwl����U����{���y*��Chh��h����Q~�ɡlA�rW��	�ϓ�Y����7�o%X͉-��C�"�
�A�g��/+'�~��������6�BA�i�	�;O0Of��_�lP/��ȝ�C�����>�N��\ж"�+c�}�]�m��[{����N���~$�.�9\[�{h8oh��slX:���:��VNT��fK9	�0DrU� :��}�;�qum����>υ�t��0n^>n!uۙ,�GT�ф�wC�%q�`�;e�ev��(=��;�k��L��[�q��:�<�"o����f9�����>�j�d}����K�ƺ����@�	z%�r{m'��0i���޼~�˩����{2���s�����2G�1�av���-���n��Պ�>ճ�fr�oTH����#&�w"�GW�4��Aw�g߄>����S�P�%y������Y�'Ԃ��XwXZ�s�$��_r��H��wA�<��y���tx��'ޥ�$Y��YYm�8۔�_@ Ā�K�k��u�A�[�ʼ&���k��*h➿`��F�`V%EFǠ�Bg���N�U(��J�t�S^��~���l�|����B�F�\1&�~�λ���I>��8�����<�5��p|[Ј>��\�bӆ(�g��rfת��g��+���z�U�T0��^K[�{�����m~��:e����v[�geL�Q�;a�9V�3m�ܮ��j��[��]�:�A��>�Ԃ�cl�콋� ;�.囬����k���	�elo__������8�܏*L��Cw��z��!�:�xyM�4�D�z���s\D9��q)�7�T��i�:yũض�]ot�v�iq펦��˴�y2�+#���j�Հ��gHԬ代T������w���e=v6�]����-�n7g?V���e����0�;A���z�aL;�m`���z��J��lb+�ӝ����Q���zJ���0S�`�d^b5��s	�v� ڷ!�}��윥�~���̟UMUI���*!����(5�#lE4��!
�؎�m����Ϋ��g]�����=��'��S���69��lt��!;y�m�Y�2w�ѱ�,[[�j��u��1~�B��}��^Cޞ��~�χ��8�C�v~�\�<ݲ��bT}+]x�2�|�u���Z0j�@s(z���LyK��Bš;���Nv�9���oz֔g�E2Y�����`��#c.'$��h�zu1�ǆ�$w�h��V��fM� k'+>���X�9-���7�׸Y��P�\
��6��;���
y�|Q8tZ�*(8��~S��s@�J挽�����"�MJ^`������w�]�������܄3�_j�2��c��R��$�N{���W=�+�����w٣=i�rPÎ���]m1v�\jܡ����{l��v�7ml���B�mj��Bl��`Y�q+i��[�$�).X�n��]�9,^�:�1?0��܍N�=/4s�&��X.��V)=�~�F�o8#�'����l���cG�U��V����[�A�K/�?e�vo_W��زkZ�*��QK�+ �J���57ۯ(��7�83�*���[�(����^.���M�HP,'�r1Ᏽ᭕`uƅ."���u���u��<�oW�����f>��#T�a/0��쇾�k�v+�J+��3�^�R�j51h^�����w~m��Xy����o>l�O5u�}��ޡ[��݌��z��wjtJ~�]��戯3pX{��ZOg�+=z||�NW����e�����͉�Hh���#�k����1B�VՐv�`9�x�ǁYYo��.���!�����փ��ن�ll��������s�X)Ouq,�枃6�6Q�=��nJ��z~a�D<^�nc���M�(�1u:�2�V~t%��P21�����V�������xHۓ!{�tSӯ"�o����r��i.Μ��u=�Wt���⽍�y�z���l�n��1tR����t����ڲhgB�����v����X�yᬹ�ҭ�Y�
D�lj�Oy6�"�z�����K\�vۼ���Y�1ܬ7��ӵ����8���vH5��f�<<���\��ѡmo��F���_�1cu�&M�}-�=�ި�sY����y3`*�߸��&�em׊�|��8���K��19��:#��y����ÁX9~�@��P8Аڱ֏g�+47OO�r�+s�ϩY*�/Ѫ������������X&T����q�j�a�1Ӎ�|7D�����'e���5�M�iq|T�.z�h�J�HQ>QP�J��1�yl��S]���=�w���Jв�y)����e_T9�3���k��0�`���m�����y�$��6	HX�6ņ���pf�sc.w��a��zUx�����8�ë�CU}u�ށw�þ/���6��`�AQ�F%L��ιγ\�gc�[�Жhn�^�'�����sl�Vw\��[����Un��'��f�t��6��:ͭ�v1'{��IF�;�Cb9pˤ�9Q%�n�;r��h3���Qɮ^�K�̢z_R{Q��X[�3'5��ɘ�3��K�ͼW&�D��Ͳ-7�)�ݖ/*���n�,��o���KQ�1άlvV�M�#�S�O���cڹZ\0��TѲ9�gd��r{����~����u��φ�o�������J͍-��C��wUw�a��r�n��+���A����,7��4�m}�ݝͿ��.�͋��fo��������'��K��'a�&�j%��u�H��N�����֏dZw]�9�)�������G�6�,!/D�-s]��.�lA�7����|^И߲yh��G�`�W/��P�0Ǡ���qk�)r�Z���A��sW���F�D�[~m���\�����AxWZy�H
xǤ�j�ך޵7�=���5cr�;�k�ϖ��z�Wܳ���&$�ku����6�{�}>��Cְ�T��/�ɥ��ѿ���nW�_G��y����j��Q��G��R;���޿�x��M[�בTdX]A+M�9���<�2�\���y�*Z���sNh�E�%�w��3������oH3��\cr��y�J���X؍Z˚�B��o���x;d,�z��-����d�Z�f�S�����a$�܇3�]?��U�&P��Ɯ#�O3���^92��4�?Vұ+��?/]���u�|�ϔ�C
��
��yvٸU^:*�LL��f4=Q$C�������7��h{��`.�(��cQ=��)��^��?�O��K�Q,*�ƫ���7�#��v"rz������=6���W˼��ŀZ���}7+~�l0�]n�xe�����_z�o�^��a�ԓ�|�([���6b�u���Y�U�����B���z�����G�N�;��ů�u��,>�S�Ժ~~��Q1��dn�'~q�1w%�E��M�Rc�y��9��m����sꓲj��r®�(l�j�U��}��6�SNiP>F��kL�Y�dfпz&+�c|!B��W>�5��>���nK�T������!;^s�u}.c=��^�A���%7�h��`/u3)y_�=�끲�R��d>�U�0z6��O���)�KΦ3:�5��sْ����H�S�mN�M�d���T���u��{�V�iV��n俴�%��b]e�/��s/S�5tj���ok���L�6`�={o���D���c�ڗ�R�VtnT��H�2�>Jt�n�K�aڥ�������L.�23���䦾Zټ
�%�<�u���?w��_�����R�+��y��5������^Y�|�3�,͌O�bd�����H=��&�P���C��G���<�믖|m�R��96s�d�`��<���VFW�re���{w���pCr�@���G5f����5)���`(�6�z:<U�d޼�*uu�{to��h�r��Y�����R��揻���ʵ3�����6�����=���̈́�_φ;:5<��~[\�|��X�o���ǲX�o��l����U���0�f\1�[��'�W,|��5*_�6p���o�u��Җ�����P4��{e�(-�����~�߸v��'9��L�h�Z<��u=��=�Dxϯ�&�ϗ�Vޱm���kȿBw驤�o�j�+&s�{�
y>cn$�_ho��Y}���]e��>���v�3��Y���x'�~�����1a(�S��nE�{ڗ�\Y�7�wH9���ڞ�fѣ��!ݏ6�T��#-��T�۩�Ε\f��ߒ�B[n��ά挴�t����`�&�7ù��R�|�n.|et�*���_��m����d��@`��wz��/�$U�_���~������DW����j����7��;�m��]g������y�!(bM��zߦ��=S����r���{��i��j����`�e�ޯ�!�����IS�f��}�;��%��HžP:f�u�����S��8EU���������x��φ���o� ����w��J7����l��{#\��џnu��﫽�W7�v�z&z�J����5361cu����7f���uU�&���w0���>T�T�/�W���GٜYy���dY����Q�CP�Q7H^�kpu�r�ށ(q�jBj���V�b^��-OzM���E���}�Q8�[j�g��T~��D�8��<�F����М�R!r�Q����q�k>�Nj����*���^�*����ӽ��^�<nf�uJ�m�b��������DT�e�C&��/vVvp]YH,=z{s��6��z�g��,+���#K�d>�a3shb��fj�,���4 -ղZ���d���0*����X�d�KC��N�sz�X�|QZ�]����'��Y��]4\Q�~#'&�$������	Z�*�*��g�Jp��E�z/�grP6�
C!
T4.�kߺ���H>��$�m�iL���V��Mo��x���H��.���ʿ8�<R��u�ދ���}}͉���D�#~�Q�ae�φ�+@�=������c�Y4��}�*�!����x}y����wn�����T?X
.�,��'��\r�g��ݏ���V:�X{Z)VѲ�W'����{o��oyt��!{��޵M�e�������ؖ���\�]O��^��uc����3���i�	�;O2H;�=�{��Ǿ܎�ά��œ��oB����z�Q��B�J�m��[k��V�Og�݌�q�Ț����cfj�nI�H��k�M�8�K�/�-sC��zx���;�z�xg��ޙ��$TD��-1�M��Kz����Y���ϗ�߾�avLw���s�y���C�x11K�Iü�
K]��1E����(O9uzD&���T��ّ�U�^�,7�j���adN71�*�B;ѐ[7���8
��7�ܴWt�k�<������V!d�����ӯ����ψgGJ�}�v3+��F'�#x�8ŭ��e��sᏦ��r��d0Cu�Q4���3��6�x�r!�4�kUwi�3����ջ��Mۡ���_&���I*�8w>]5�^M��!H���X��͊WR��B��z�D���u�M�7�����Y�8�rJ�]XUg6C�pm0�[�*M��+�c"�Y�x�l�l��q�
���2��n�q�Pz�I-v��aފ�k�}��$ʆWk���%�v����:���ʏw8i=l"�[�'E���Q!G�,r��l�O:��֟ډ�]y�+f����ܧ�d���:������@;�`�"�i��.�wwSv��v�v��,��s��S<�����<���f	�!� ��d�-Ɏ8��wciY��;���2�nֻ��=���a��c)D6y�l�:�wSOH�N0_V5�kpY�sV�C�����r��l�J��I[�!iɂ�f��r���#X�K�����ɍ[Z��N�􍝷�"v�O6�p�Kg(�ؗ�s.���X7�s�M�U٪�0�q��s�@��4/��i�T;�:��Ai��-��1�ۼ�0�4�qx�($�Q�c�� ��]nqPB*B�0݅ ����7H�8��=�Zt�f/�6�������b5���xe!n����<Q�[�$�E�H��l�=\KX��������ھ}�W2���P]wK��*�v��\R�8C�}3:�S��B����N�o���uݑb[�v�n����6�V䘏n�%'�9nr޻��6�6d� _n�F�RRem�֮����qgQ�18��퀳�����`���J.Fd�)�(�8��m�����,����Ұi8'�1"m�V���Pd�Up����d}V&n��ff�-5�4�K:�A���hr��nǋ,tm'x']�Y�w�iɵ����GH�V����h�\އ�չ �y��N{�d�G��{*�-T�%p۽y���7��}�D.������'�mmm:�׹����Tju�{PMu��!�o��M��<��S�Z���p��Y��y���3i�7�١,�-&tЮ�X����H�
���Q���E�V�6C��l��R[G��}�a�pa;�ӛۛLP��p�y	r���� F�+W_m�Z(���I��N�6��W�6\�Zb5�ʚYJ&:�j�vw	��̺i�۬?:qͥ�5c��J,�QY�����^t`e�֧��`�g��d9�F����vj���0<`mi���'��%�m��P��\�+;hq��sT��楼C�s5�8���:�7 Ln9�mZ��Y�Y)^AŝN�q���I����N}h<+�u�s2�᢭�!�@�|��ϛ|�����}�ygM�v؄�q���"A#l(No�{�F���ݝ����=���ނ#��{vs�����QѶrvn��ˎ��6�L��ŭ�F�t6���"YZp���vZGFLj��/2e��.�r�>��N��u�6��$��:��$�me"Ts��;s�;>{��wfvq�Y[kVٶ�L���� ��芒9$�9lu������C����3meϋ��JN+�Z���+4"��f6�FVƷ.��� '��n32��Y�(�V_5���*ˎ�8��kq�*����4�"m����[n���"�轷�ēj��H���kJ��ǵi�ְ�8�H:rNF�n-�,��<�S5iZ$ێД��'��9Ľ�m�{{�+��+D�c���b!3:_=��pP �;sW��r]dpo�o�7s[���r`<P�������مK�YOMK2=2K�m�_L�	8�W]dR.�ۄ��o C��p�n�����[5{�|�Vʓm\�=P4Ѐ�An��y��>��7��B;<��~������ܩ_w-~8���'�
���<���f)����I���k�xMr��|�ZŁR�h�?&�U4x-��9K�`z<��yw/�\LX�@�5#�߬w���|��� ��o�~/g������閹��Ƽw��̝{�=����-ď�A���/
�f��{��h��v"ñ�1��O=���0�`�_P�\<�U�-��� ��uO�����e*���]�`���gO�;��$ߪRƯ����������,a�/ڽ�D{��<�	��������j"���%_\h3l6�*v�����\S�6��r��̿!v�i��ɱ�|µ�� ���[���w�F���͒27�5ޅ+���O��(�hz��X}����^Z�]�>Gޭ�e]�4���x6]_g�g����67��_^��l�Q���m�g;�Ue��ǥQgH�:�NƔM�,��c{�JA��
U�w��4�o]5�3{�?.f�:�f��H���[��K���\���Q����x�׫o��JԼ撬ңY��x�fΡ�֊k�ؼ<����#�O��6��h�030w�����9|H"�5k�����w�(7�ClE4�HЁ�~��蓗զw�u��7h�z�)��O3�:Fܲ<T�b��c��gHO���f�:�n�L�v'�ΐ�v��g�A�Elu�{�ļ������,1�Pj];��O~:�g���{�C�����4�o +z�3˭գ���Ƒ�W���x�~��xiBxy�ԭ7�p��`������&K>�<�	����nvR�oNo���v� �!�W_3J�Kٜ�9��r���t�q��k�^��s��<�D�`f@u�;�0UH�`��ycR�!O>�����3*�l״�β�.˿Q��8؃���a�ᴻ���#>�����^�%ˢg/��ތ"ɢ�&���	Ұ�c6!��b�����a��A�eխ�gs
�0ͧ7��u�z��|A�Y0�دf�"�7X��63z�����*�I�|_l��.8��{7~�U0L������t�ɬĦ:�w:ڽF���FƄd,Ge��Ӿw�.��1��<�Q�Nv�;Q���6u+�2BV���hfV��3��q��^��X���2�yp��^�aL���]BGg�}O�u���*���o{s>��6	HXO�9�1��5���F�m�0m�M���.���uu��E���>3���X�
�oX��;�+�����U����L1e���`��B���������u�y���zi#��s�C�uI���w�_�;�շ��P��)?`��3���|��*C���G�}�� ��@#|�x��e�>�Y���������ȭ��Г1V�$�G�܇����-7�i�ݲ����;>�v���!C�UD[�^��o^��}�������z�T��-��Ͷ�$Oi�3�):�a�q+ӗ�н��]�����W��d�;x���n�2�A��|<�qӪ����Lng�;��D\��.1d����iU�:ݡ����,n������8,gOE�v�uf��&�w���|���]rh�
�2��Q��c�-^Ap-wG*5�A@(^_d鹒8�Z}c7|���ײ��:3�e'1��7�x�W�[�ˇ������m���VQ�Q���*?���讱�]̢�nD�%)4�ܫ�X;Q�(2���~3.�Ek.���}%��Q��^bRv���j�_.��=�h���>E�}���9Gz���0]֏#B���8�[ԕ/i�W���&G���/�^��<�
'6�g���pQ!�,y�9[2=}`�w𚥶<�i,�˛Nj.+�F�\���D*�TU&��n#Z>���9w��Hyѫ�-u��w��/�,�^J`�W�E�}۳nw}u�b5�2�GU��i��^�ZH>��>%!a6ǽ������={[u�~��B�1X�d�q>
�1���[ۼ���sb}�Oo��n>y��&�т���$���;5���2�~?a�~�V�e��<Z�nA1٫��{�Ը�wɇ�i3����co%_\KkE!���%�(N��V�RQ�ΐ���9�����j�;;�o������\�����!�1��1�]��31���J��l���ׅz�CL�݌7� �n��������4�睑��*Jt��P���K�m1F7]E��;h��vCD�O���mS���{��7�gv��n����|-K�n��r),c��;|�Y���-b��V%ҝ"}��h�D_�|Ń�Aa��	�����=?�^��������0����O��v$Pk�%��H3���J�M���4��#�Y���+�hO��Qh�>�lON��+8zh!�%�p�����-s@��m-��2�]wvz���7���+�OGX&��:�2Xc�$�������g?
�=��tK=��"B!����X��i2��W"�=P4��$�7�<��2���[���^�k�ى5W�>�XwXZ�s�$�	�3��w��>�'"�Mr�xk`H�V)Z8�x>T��4Y����m[������zjm59��=�5!'c�;��k���)��}��`*�)�yo/�/Χ'�['Ș�c]�(y�M0�H{Cj��k��4�������C�ؓ?�uл���}��1��%���8!�5%�<�U�-��zH!lu�:+��^y�߽�}Ri��"��a�`8�$�a�2�P}3��ב�J֮���pl],�Թ�[4#A���p8Ne˽����]��jW`��H�:W@�I��A �{�	�N���<��Vr��xtl� ���/�\׋�A��8��2~4���_�������Lk
��m���6�z֧�=��幥(����_x���!6u7����)��v���:�D�)^�<����?j�=L�<�~_�5������[��E��`t;��}���{l�緝LF����hx[���]h����me.��`&�7���g1S5�/'כ[Z)�
l{�<�k��,'E�sM�p�U/}]�ؖ��]�)wfOn���6('ü*���?<��|����]Sw=9��]D!/U���{�)�K��ʸ���l6;Eq���Vo�E���FMl/yg���
R�V�߁�eo�֭{�ļ�G�=����V�R~�N!�^���wr+��V��O��o�����M�3h۫��D�]^^�߱a�y�G��}�5<��u���� |�3�,�'Γ�a�N����^������Z�m)3�2NP����QAϯo����Y�S��&���osJ2�u�]�l��;v��`����ͽ�����P�v*#�����u=������;��:�h�k;^�Dolޡ5L��7[��8�`����Ky���*5�;��Kd�V���m�x���߫��k|�{97�Y9]5>몃p��AHx��{m�/��k��8�P��_�����<
� ŗ<��ה�lwU�q����v��u��	���bBW�iw-��f���b������}3�b(�4�N��X|1�8!��x��s״*�,m`��^͗�5�y���`�i{K�bB|QAp�`֍�Sޝ�����c��Q��N�ں�'���w#�jJC�O���}��Y�>��Cm`���C����J��su�y�:�z���W�z�y��m@�\©�����3��g�^��j4,��W���fsx]a����g���7��έ�V�1b�.�G�����J������f��H���Iy^6���Z�5��B#۟i/EYy��݆�]��
����갯�Oc;&�]6mWxB�V6�U�Vɻ�3}�WjN<�8jf�y�^��*7���}fQ�ʶ_�LI�J�f^�"��J]@��0|����U��`*vN�7]�|ch��~!����:�M�BQu�������n��_.&N�4[=#Y&�[%Q�B������4�n�VVG[;��TZ�f�t��~��Y��j1�!���hvm`iQ�=����6�(��9#�|t˪[53ޗ��!C�Zϕ�^rv��X����_��a���c3BHzf
�f�������(tm��^Y>n���ғ��K�Qg�Wz��<B�:��K������ΠI�{�v@}BK+>�e��"ߩ૳�:R�Vq��/�{ؗ"���}���g H�@�>shW�{/�y\'�ꆐ+��,�s�yj���O>�Q8�[j�8��8(cE�a��oEYڋ��z����BGyY���,�ͧ�p./�⨮x�h���9{Ѿ��c��mA�g��C!|H�~�|���@�K������*����I\V���F=��P��X�T.��޽洐k��&�)
3�j'%�%Q�B�	��K���1��y��E-�ӏl�s�)���ɦ{j��n{)H�w�r��[=J=�j�|�L��,WY�-ڙW�o>}�sS��c����}RM9I�>�p��v�Y+����=-n���]vU-�V�����L�wWV8�n������P!b�;�+�]��੍Wu��]���}��zb��2OM�d��`�B�.�}���`�N��Ct=Io�?B�˾�|//���J3+[-{�9����v�	���v6�U����ȕh��7�_��V�x3=���߭~hb<^�q�?`-�F�+;��}{y*���+�*����3�һ�+��l`���ō<��=��K]�H'8�<X�½��׸o�ë�$6f�}��scE}r������+�ҤY8��4�ɭ l̉�P������Y��I���W�m6��M��z)��3]T){�uj�&�W-�A���kz ۰���	�bu?0ǫ�$>�-/���n�4��I��vl���᭚�o�!�{�+���]2���߿>��O/���="�|+o�x�]��X���_w|�������~@�9�RD�f��h	��EJ���&�2jٚ"W�M凛;2�~��.X��)��fu-1a���>�\{���:*�ug�=��k�Q�fS�E�w\�]�����r�#k�ͫ��Ȩ��OP�w*u$P�+M.��+��2;����@�<��� ��G��3�	}u���x/<������m�9�\o�r2�e���������m�����!EPj���z�z��MS��]��Mɬj$��Cb(�/u;tVv� �q ��6���WC7�`SǚQ�X<��vy����b���u�F��#b�Q?0�-�~Z(�7\�P�%Jo=`�X���a��a&ŧ2gA��c�$�a�>cWI}�O��(~��Y�G�j��s�Տ~|���I��O��=����o\	�N���=}ݮ��p��_xv���*�O���l{��
��o]_��~����ʕ���L�w��;��t7ݲ8[��SȰ��L;�m��ge��+#g��٨�qQ5Ӎ�{׷�o6$֊/�"�����_X�a=���m�Wx��`��ߪ�7�$�m���8"�'�o�{.�lH���M!�Z~B�P�ǁ�Qx�z:~�~������uWe s ٳ�R�l��G����9Q��צ��5�t͈P��{I��l^�&���ƜF�"��2l"W��{���=cv�:d+=��A4w+\E^aiA�˺��t+7㴴H�r����yL���jw#W{�t �7 � �������n�t7q�`��(�h������S�Z�Y��M��)Csy� Z�+IDgD�7��nіo2��� ��\����so4��S���%N+;%Rx)��N�Q���r�9Ye�C�-뾧{+)*��D�z.L ���u�f�� Z��l,ʙN�9Y����%\&-��t�q�9
���n�+�l���x�t���C��^��3%�
=z�Yy����{x�L���7��W4��v���+��kp�QL���S����R�4�|� �=�zeW>T�H�=DZ���(�+��m	b�G�wX=&�w#��jVV�����&�/�L������
}C��I�4��9F�m�1q�Cc���A�=X3��Ƃ.���]:m\@���"��}5������7�����
���1�s9\i��E���*�Z�P�{��l}�y!X�G��զ�k�����k�. ���:���|�Ԥ����.)�\�Q�(�.�-HE�S�Z)�[�=)��C�.�٘��ɝi�����j��(Vok���.�'�EgK�*�g�c����VR�r5��U�M] �c�׵1�%�l#I�+.,�U��pe[G3��sU�� ]��yn�#�R1ԗj& w �D�˳d�B���4��C�������n�p+���Q�t��z=t��ăw
eݾ�zMr�`	R���{0ϟ]���XA�%������ך��Yf�kwQr���c6*�zR��3����� kG�[�')����S��]Z؇��L�+`�S���"0d"gZbh�tbc���b�[C�WvP��0�U�ꢱ;C<�JD�ڸ�[$�N����u���Ԛ�����DR:w	uAsi�h!���aŌ�Q>+&Q�����:/eq�;�T���b���+�� ���>9	f�qˣx �q��,ف�z�z�uwͨ�]��z��6�!��l����b�V]���*uٓ�g�{�WL�9S���b�痍��5�sE�G8���8`X8��X�oP3���)��+nmK\��AV�&w�Z_��}2h��WҐ�Z;�� �ݷ��v��0T�8��2��Ո�H�Iu�Bl���ۤ���	�Y�I9w���~ö�3 �U�}q��Á�twFTə���tt��B�X�>m86�UL�m[�+N��`Ǘ�ލ�uԮ�;�B�sL��7z�@5ՎHL�{���{�t^���t{�&�B3ˢ�l�/�v5ܽ{2��N��gK9at�u�FÖ���Vst�E$�ף���z&Yv����{y���s-�t_Z}	$�bXa�w"�2X�Gc���[�I UhD�BtF]�E!�Ӗ����w9Rm��99�W��^b��N��Bg�jQ#�8��[X8�:�3��!ّ�w���X{�<��ۇFwh����W��o{�^m�7&[׷w�m�A8�ݨ���D�,�ӌ��m�[t�;���zے���ŗe��$=���"K�{zw��fY۾=8Om9m�#�i�]��mep&��#4@���|޻�)�FݶӉٸ�^��G �y�^hI9fJ*�vfլ�vrw8�K�����Ϟ�p�N<�ͫ8�&Vkmml�6�"I':-��	��Q	�ӅE<�Ȝ�m9{7״r+�ۏ����=�M5��,,����"e�en	��\�me� �B:u��d@���� �h�+)M�{�V��Ꚛ��:�����1e���H->�X&_X��J�}�火���cM�r��Op��-��n_$�q�j��j���f��߱�i�'M�ܗ|�PCa��Ĭ�2u�̭���U�����yJ4��6���V��	y_��O\���(�걵�.���hlOz��	�S:�l���ɿ����mӋ��\k7�[��u��p�y�����h�?Ʊ��a���ٟi��>u�����zǳ���L�[>�q����T=��Au �W]|��ŁR�ro�=����fǬ��{`�#�����9c�; w|G
��Y�}c���j����Mf{̣ҽ�0�%�һ��p�֨������@�p1!��ܳE/=��؄w7�jf�'7��y#�I��'���|-���@�O�I�u�uJ�'M��Y��&�ʲV�,��
��\�/�;-E|�b3r��0H�ʁ�{�lz�G2�v.�������޼R;�|=�Bl��v�.���������O�XZ,TZ���'3.M�����,���\�p�����*���*��.����������IXj˰=����s���Vg��E)(�����X٨6�h�*!9��N=doB��E��ͩ}�6�L�?�)�l��[��v���Ir1:��v�?�9+����]n��]��{Ͱ��	���{dm�����W]�g�����}��ײ�Fk᡺�{�]�6�]e��M����D��Y�>�B""	�
��o=�e\�b�a�Oދ�)]
�Ȟþ��OV_���#{��ӸH=�]��/Y��o��y.�lH��g�u"^9]�'K�4��g�}�^�3�=������Ц���ƨ���;>�t��!\7�.�߲����p��y����w�!GT��m3����Ê�W�ǳ��'p��7K���xy0�l�g�uSK�h��>匬��:��������D���f����!��!�Ǩ�J�����ms��i����vM�'җg�g�h�]��}�������j:�t��Ƨ�˔��Mw��Kم"�k%�[�� w�XC�@��zr�ḙ���Qh��=���v�h(�yՔ�N��V0�d�Z�<.����cU�1WӤٕ�����X"��ʨ��v��Nb�\2*�ܧd\��[FpzpG� aqe��}�+%��L��]7�ƻ�U��������S�";��<��΍ّ��4*q��y3w�J�������<���<��m�m��6B����s�^j��<^���$͇1�R9샺3ȼ\��������m^���M�Fϳ���X��z$��m_�tu����e��ZT/G'z=�
����p5�\�R�g_�ʳQ!��V�<^��H}�j��D_��4!�9D;�9A&�J}���ro�0cU]c}W�2g����L�Ɓ*g�K��9��/F$�%a	�}o�ɠ:�pA�ޙ��q4�\u��t�z�ĹN_f_�X��3��N��Lm����o��m䮨�8�P�=���s��>�HX�|3�<�z��|8��kV��]��t	�^MO����&0N	�o�z�K�M�>C�̂���Mg��{�U�:�|b+����B}��o"h5����7`�!C��&�bo}uU���7y����C��J��J�ݒ伵�˫�ukB��8%�^��9�W���U⁃��l�/��"3ם8���s�lP��X�<щ�3';��޵3w��{��5~�p��b�Ѩ�cL����3�rs�d���yt?e���d=x��	��
�6����<Y�ޞ�����G��HC(	i�vס����H1�F��a�:G��+U�c��ƞ��o��N���O�1"~�"ݜ��zkkg�ΧZ��o�Z���.m���6�OGl#��]ε�k2���r��	��G��<�|j��O��Z�G>[�ח��O��];����`�.$>V+���f���q4������;���9��U��1��nS�!��G��:�F���}����⎀�Yc�t;���0����\bG�V�y`����vr�1����ܵ��G�&�����T.�U�ѱ��`��4�TNދ���7=�j��={��B����K���4�)îf��m�Y'���W�(^F�\�̱��]bue4{U�b߂�_{X���o�j(�wՓ�^"w�t�~��_�G Vj��J���܉��Ty��;�[�|����~fe���W9 z�J��-��h��r�Iش���V�Iu/��:�L�e6R��o�8Ŧ�3��j���cX9/����95{ܖ�����+9�J��Q��M<���{\Nn+��c9�[w��}���6�� V���N��.�9�vj��u��o�!1\�FOW�q8�k~�{>mz�"��5:�ʳ��l�갱�\�z���g�ݞ���U����E�_�y؝|�u��F��M��T{ג����j��jܳ^�o��͍��tJb)��ݭZ��6��g��=�I\��J�I����N׍�m=��7/�k7����>��w���9�f�>SAm�V}j��R��=齷�wؘ����5�n{u!��cC�'�V>�@�K8����
�X}��=c(�
��-{=�"�ί��_�3BP�b��5tN��~��f^�J����F���'�+Gտ��O.�V��8�jYW�u�ύ�X�{�'2����N��+n҃=�yVN�yc�d}Au8�Mo�ϧ��o!�\���O~3�'�u��HK����zX��d�
�:�������*m����T�Л+o��:k�ݘ=�:*���sr�����g�PY�%(�w��q�.]۰<n�S	��8���ӛ�n�DT�k��b��Ѻչ��s�U���%�3�J�9M�6	�'󖼜l�V{Ю���?G}2%Nl��A�c�csǕW��m�r�EG���2���d��Bk�+�tV5�|�x�cЂ#��/��A ��'�h_�Bvڊ\1T��\.�egg:,�y(��(]D�T�B��ά��|��B|)�&��m�݅՗[H�_T/��ם[.�Ъ��s����`����a3��J�f�=^�8k��])�X�Eg�_=�`�HЧu�����
���){o3���I�"���{�G�+Z��L�Z9YW*�Q,=����[.TήvsW��!�'�W��,=�ڵ��+�����o&�*ϧ釽r{x潢��kG	\7��+����ޅ4�|�v�;��輓��^��M�Fg�u�_X^�hm���[�M-2�z���>ֶ�g������*�S�/�W%��P��W\���{�N�q�b�tI�5��N�MZ�7c�θ��&>�[�	u5,H<V_bF�X���[;�Y��(��G!XV�3�����RT���b�	�}Ĕ8��r���h�E;�*׵ɳw;����dr�}�:��^��&�!�����Kf��@ރ
��5��o�6/=�9��K�!(�W���&|�r�ꁦ0�A�E�룓�}�i�s5��K������|��<m2Oˌ�u �=�h��@O>/�ں>��-�=�]~��_W�	���%�k%�>�[�g O��q^�=��oEw��)�B�lh��n^�� �q�3��Y�Qcz�͹3��ʃ�0�/O#抎�/�<Q*�<��e���F��10�X��[
$xC[7�u�����^�Na�|8�/������<��J�������)��+�~���5��r��3ڱ���zI�ZI���-&Ŵ��}9&�b~aS��ׇ��K��U;�˸nx���D���W_rbl��Z���q{���
�%wd3{q�_�)�h~�����gr���7�V�����M$Ү�����i,�`�h'���}tk�W'�2Vګ3q�ָ�^�ztZ�)���wA"j�A�� �yo�����a��\���lqR|2�2鮃�eЗ��S��-kYpb'�TYZg1Ͻ��N�6�����V4���}�����3����B���*m�lzE������T��ˤ4s��S���ŷ�Z���s/O��	Do��*>�}�`����HA�/[�ؼ>Bϙ��Y����)�g_E�WsCO���.�ƹ��JN&�~����M��a
�*7ѧ�>�G;��ޫ@����%W��H�d鿣r]��!�i�v��v�$jT��w�޾�!��|L�M���i����N���Ha�v����D{�_��W"�
������5���c�.z�L�<�=~�Kfo0Y��T�٩L�O@O��xI����Ux���]�����ؖ�WWXw�|�ϻޒ7`*�����?]|��f��E�����`�b<�苼�U�{���X��&���0e�@���޾�Ǌ�Tt@���C9NxD�]�h��Y(�(��Lޘ�{(�n��P��\u��� ��~,/SƸ�'[�ͼ-��Wc��^�V���ϲ��ܤC'���c;�8���JO����еj���p�Ҩ�wt�2j�q:ם��0!� p��VW����^`'F����1�ǾA����t>�q���޹+V�+���4���m`*X*���b6#L0N�e3�����I\J����V'<�7=��4ؿ��\�Q��}Y'�
o��P�c��=+�<A�k����'���h\��b}��'�,��n;�o*l��&��K���=�DTܷ�ˉ=TC��s�4{Mm�l`��uLDH2�`ɏLz��7��_l�!��nB�\h����l�y뮰��A�mAw��5V�W��Hr��=�>��ʰþ(�`�ha�/:�y��.:���ƪ�G��!�Y��"<�+oV�S7av���w�('@D���v�L_���7�;��r�_o���ͬ��%�<x�y4�K��K�GU���ǟI>�N@�#���ݟ)����edu�+�������U�D�Qͳ`���P�ۛ�!q\�^�c��"��g�h~9=g
͕�@�9O��$���"�Ŧ�QӒp���,`���T-�����m8^��@Iv֥��m�F�c���Z*,;��W<̹�95)��9�{��j�:����s�q���cg"��O�Հϐ��K���gԬ�hv��
�^��VY���gt�����G�@\ן��﵆�(r��g�>wc����<V��jN�s#<��:��?7a�Nڨ��|��?eh��ҵ\�{/�kK��[��4��l��.Gr�i�yc�; H�Ї��C�		����2��V{D-;�+=U��7�I�
y��̤���8؂~�|v%�C~����q��V�����5V!䍯6p)�kBp�r����q�O��7�Mۋ�YꍻK�p��cbG��&����o@$�O�C�`$bS8�s�3����x��؆d����ӷV�ug���_{ڄ�)	��5�&E^����1="��<�Q����C�?d��I<n��=��ь6?:�`��>�/�G�XKP��	��yl�`2�g�ԭo�}&�������J	΢����
����R}b�"+;=���(`Q����wuV���Ie�U�uT�uT��T�URWUI�U%Ww|���������ww�UV�*����Њ*�
�
�����]�ܕUI�ww/;u����ww']�ܝwwru�^�W%�� *����(�
�m{֗wwrWww']�ܝwwr���
�*� �����]�ܳwt���ܝ�wr]����ww']�ܗwwrWww%��ܗwwrWww{^�Ui�ww']�ܕ����ww%wwru���www%wwrWww%�RګN�K���P@�U@�{�ꢀ�( "

!�`�ǿw�6�qm?���־�>�+�O�ĸ��.��zB��E�t�N�TV�c��݊(���� U���H:ѩ�Q?����"���8t9�<�HD���^G���9<i@�APD{���UR�wUI��ww\�( o ��T��D�]J�uU;�]U.��U_=���o��q�> ���������2�z�r�ކ�o�Qը�yQ��y�K��>������0���QEErv.��ͻ�1����b(��H�,{]:�
�������TTV��� Q�*70����eP��/)�ۆ�E�x���㷝E��9�Ppᆆ��V�;_`�`o{��(��A֢�����{ n���(�������#n���E�c#����n�P���k��(��ὩF�[�TQQZOo�ղ��{A���
�2����(� �������9�>�8���_T�UE
PTU&�541UkCX�J	(M%P��E*�R�*ٔ�J'��C�$6��f�R������d�
*!Jhֶ�ےT��eDխ*;���l`km�ȭ�Z-(ҐiF�ULv뵶ɥE���P%W���i*�M�Zh�E����UUfiZ�F��ݛK&���Zԙh��0�k6mSY1Y%b���J^�S��l�!S-��&�0�j�V���fԍX�5eb��X����kiT[5��2Z�5�T�  nZ���K�s��z�)�[�v�n��ׯ:m{e��{�V�֏v�N�n�=u.���^��4뺚�Y��wt��W]��w�i�ou.=������tꛞ�]����oG�����V�V����kD�   !�w��bD�lHz7a�Gp
(hhQ�	�=
���t4(P�������a[s��\�c�w5Ku{jt��g�m�W�CK��`۹[��z{��ާ��ݻ��ךk�ս�OMl�U3M�0�ͭ��m�ٖ>   �omW��sR����v�n�]���7��nr���4��l�j��-����[+[/<ݽ�^�=^�������/@W�S���a^����t/n�Y^�z�t{��ۮ��{R&��96lZ�f�>   ��jŶ��=��v��װ�r��V׶������/Vs�^����m��t��[��^��wi;���m4З�]��W��{�ݖͶ��{�ݏ@��mp�\�Ͷ��u�[Y�2�ٕ6���   7w�h�Aں�]t���ġAyv�]P�G4�n���� eE]�\�]��ʦ�7V�E�;��ù�
�V��͉�m�j�������  w�jڽq+���7e�T���6�h��v�*�A��8���`u�m
���֎ UQ�:v��+l��u�q��F��Z��[e6��  �܀F�J5>��*��6��G]hu�a�j���qE*�j���l..�*.6 
��lu���{��$�L�F���&Q�e�   �������Q��\: �t8 z��,����K�` {��  ^����uB<��= <� �Z7S����mVb�*�V��1o�  3x>� ��7@� � Zwxy�=
 w�e�@:Х����^4���w���= �zx҃�w//xPz���i�[e��l��ji�e��/�  ��=:����:Pn[���G���t g  ؘ .�\( �s\�4�{W�� �ދ��"��1JT� S�h�)*�M��4"��IJ�� �E?�� �a � �M 4 $ʑeU�O���/����s�����&�K�bfsiT��FP�e��.�z%Q�ǖP�������dF�?�l�}��m����`��������6m�6�6?����y���?�?�ed4v���oB���J�JĬ�i� nm��C%��J����9�"ܕ�*�v��e	�W��՗Re` �8�ˤ��N͹�um^��%-��-�.84Վ������$f�o
�hS:�jb�,�y[Ò*6��q���aL�v��F�Ա0�a�I�0�h�/SY�.��Ӧ�bʂ�*���;�5c�Sʩm&i�"�4$V�H]i܀�3 ��CKm5����N3�T�Z6n�fc�x.] �3U.Xx�����8�Vl�6T�H�T�z�:7�(�t<*�zUf՛(����M[v8p,T3(��W�.�R�&I�	;)$��[���Pk�5ݪfp�Y#��VW��iQ�Bf�":��B�p����߃�7��I�ia$X$�V�!Mʷ�M��=��k�j+1-�b�Z�d��An�[z�hK���"c9a�Wwu�؁M�[�����(�Sf4j�.3!w&G[fQƐ��D���^ͼ��S�Q Y!Lĉ2��b��a������@����&-�WJ]��,/Z�%����̦�z[�r�[sFIb��Y��2��5T�zI��!�h]�uc)��0n����|�����4�f"-�4��.�c&U3��^�#��JóFK7�fcm�ψ��ˑ^D�//T`�� ^\f�'c���μ��,d-�4N�H�.�8Ҥ���0�J�B���	Ų�g0K[soqH�q�kՔ�r�D�l)�p�"]��0�B]�sc��d(�ّS�_%t/V	>�阨3or|�1yyL��j�ӬVl���U1�"CY�Ȍz�d�S\�r�Y�w��ʺ1i�⭴��@˥��e`ˠ��U�mH�)򭩂��x�n��̢�,X�R����eJ�9��G��&�V���A�-e�����0�.�0nm,�N�*d4�S�$C�n��.8p��f��zS�\��v����J	�-Ml��и�d��.�̫-`��(-)h �v%�d7������Z-�E=�a�`�偺�Әk +4`zCА�ɫFA���iEw����tV�J�q֝�6ʣ�*���%��k�.L쿬R�N�M[ec�-�`��pX��;�l�N�k�$���hC�X��l���ՉVV�Z���u^���R�o� ��U�}Y��GR�={`F�X
L���&M1
Q
	Z�7En�+�ڗ(��i��f�SH��kub%,6n�y�����ϲ�9�P*]`̤1ݪ�P���kT�L�����{X%֩vd��7�>rM������;��+7,!uܚr�F�l�z7Z� m ��dOj��0�4�˘�ѳ�&Ͱ�.�ƣf&��ڂy)\
n��gagI��{t�������ԧ@-9lE��� = 5�MEm!� ^ۆ\���(�$��;R�n�ͧ��4U��ܸ�����K�;�Rio���m`�h�3�3�u���0:M���P�b#r�o&S E)���EI��4^��#fP�&�f���6�ҵA��2�^R@q�kl�t���P�{f�#n�l�XCO*`#-�AJ܈�G�Xl=��@N�ɦ�z.͋��o2�b���F�WצZ��i���4d��.�Cwu�VA�f��ki��SŎ��2D�ͬ���P2s@�
�ͣF����-]O�`�v!nVQ��٫�OEemj�kn�2�K�ϓKݣ��;�ZVnģ����m"R,�zY�5ARo��K���)�����a�[9*敶N�3\��2���aQ�Ȗ;�IM޺9�������z�q	��k�A�5ukq�Й��0���y�(ݴ�CT���T�L鷆�7*5��ك�H⣰Lj���� :cY���qҔB���ˏ��� ac+����5gU�RI=��l�Ee�r�N�S,�ǧ�q�{!�VQi��M�P�$ ݍ^Z*ŝ8�����������!;, �W�E�;Z�##�$mA)�{��ۦ�AF<��ŵp-�T����m�+�X��[��CF5�L��q7Kk[�m0tIeq*sI�x1K�틠�FH�w���0 ��n�@�R�+��W�0�:�\�҂" �(�3^� �<4���壷IR�݀pA�.�B�wv���:O�o6��[�b���(|��aU�0RE�Zƥ�F]��g\{
[u6Z6�⤎���V��6$%(�kNU��2S��
�Q{�l�l��6��a˭�v�x��a`�v1n؋\6�X���HHB����D7��F�̣i-���)J���G�(��/�Cشz�ŷ�ҐS+.��౉۬ �A�Fb��%6cRkn���6�m4o&ٹ[L���i�'�k2���Ur��dP�^2b	�n�$)��e%ge6Q�KY�/V9j��\J��3T�șBz��wS6�b��U���m+�o(�܀n�{�l{�M�v��8��)�O�e���;�n�;�b[(�+sH�R��f�١0��B�9����a�@;65Ѷ)���9w��\ɫN��l���X,9nPz��ݶ����f��-e�0G�]b�Mr��&2��X�۵�V]�}�L��^^ˀTZ��׫.�%�}��4�hH[ ��6D˭.,��Cr���X�n*$�"PԊ��F}�mc�[mPEذ������Ȥi��6ҫ��Q#f��w)9��R�(��F\ƭ���J�Çr�2*&]��X2��@�h�P�vi�-ĮVV�XOn6��JB�i�C4���L�EJaaғ	���tnT����*]��.���^��J��+j$��j?K��Q%��ᬫkN�G)��Wv�,!83aH��7z�J�d�D����)\!&�$��
���k���`�҅�/ih�H\��#Z��ۖo�C5��Av�eM6�k��x씊��B`C#f��b���w�0B���i�}��+�1M���/8�{s�@*��;�eq��u6�� `�L�S̎��V���J�e��p
����iBrk�W�����z�"nU�1�,��֡�ҙ�F���B��x�E�bqh�Wu�7A�աx�^nH�C6nM�b�Z4��Yn����qZ��9s1�*�@[yY�
ˬ6�"F�v2�#���2�=�@�v���/n����G��	�̈́�`�6�d֩v�i:�(�v���)��HʺB��+ ���<Ʃb��Vhl<��%凖풂���P^�U2�ʙ(�R�e@�-�B��nm�7V<.�t�#(B@��j�4�B���f
(��f��,5���Z)��َ(8!b����������M�5af| Vᤲ���Cb��1U��l���J��f�����f��!I��5��'q<
c	u�Z�m�Ǝ��$6�� ��u�`�KT)��6́3\��/B�k��n|cK��E	E�7�/i�,�	^%Cf?��l�����HX���1�.��̚(ҳzB;�'+h�(7#t�=��(i
�14���,��m�M�p�=�d8�෰���c/6�n0b�&�A+9� �P �݄��I�j�����M�����/#l̒�[I��$�m�1X�YlIz��ڶEc�����L"�J
sq���JJ67]�;EQ�yi������e����i�lH^�#���QJMSdh���d��(IR̺�����ʹ����;ݭ�e�oF�l���>͛��� �bz�X	ҵ��b�u�É? Vػ��&|<)�)����Y�-rԎ%KA\M����B�b�%�i����X��˦h���f[�y�����zQ����F �{�	:&a{��##[M�wY)VQc"ÛZ.��me<E���O)TS.E�hn����+iV-m�mc	�2ͩ�>���.�i���6���Lf��&�Ė���9�%�����&�C��j�O4���Wg!a�m�Hʡ�Sh�b��OKouFkE�����S�m[ϒ��ʔ�)*l[�[��Fe]:�R%H���w%�ԁ�5�᱌I��^D�\�2��ӑ}�
�A�0L��B����%�Z�2�Z����3P�$�l�{�%���wN5�"��%<�bx�ݖ[P���� e)DŚ\J٠L:v&�XX����U�j�u�K4sU�5��s(�yXi¥�R:���o\9F�h�۱Ss@�a`�K]#�#���Z��&�FL��I�W����n��R��ݚ����ŎۘFH�4�#f�R�Fӌ��\�o2A�F��(l̻tQ��!2�P����z��	
���z`�tc����̬GYۑ�˖ޥz�2R���$VKr4q<��b[��i7����lB2�%�l�T�e�j5�� tX���7I$,�7(�y�j0)dPCP�[��a��L�]꒙lSɨ�T�2�n���J���~*�ρ,�`�bۂ���/;��5k#̏Rͨv���UÖU���O-8*)^�1&5)
.m�x/N�2t��KI����VtH��Mj=
^Vʴ�[��3 �"�����x�(G2,�n#kw	Yn�+S��s>��O%`T�hb��0�gr�T�e�8��Z�p
�*E{pV���KF$�o֑�UaOX4��n�!wwrӊ+�ʆ���Y!���ܴ�UnV��5�6�������e�q����N���З#n��V��5�m0�%Ke���t��3*�GN��0�m��z$� fnC���
���a�vc1�r�k�)��� ���	B�~2<�Y)J�W�1���P�rRE����t��zkE�n��oKN,LՏ��\$o~[2�kES��Z�ɬd�uD�NL;�����0��[�7[�(�]�Y�i�q�%�fa�hA�6��[�F�����3+V�N&h��.sXIZ7Z:�A�@�e��k��>�זSE]�!Z)�1p@:F�@�Q�2,�]]�mȨU#�ڋ�Ԑ���|�˼�b�h����.�lN�6�k6�"��2��E�@ �Z�dxl�]bY��];�le�/+%L�#��;�������v���xݬECȳ
J��v��+���H漉�B=	 �hgufS���hH�w'��9�+8�=��cIY�м�HYP
2m�
́мPe%��O	HhFޜK��Y,�͋Y�ff��У�n�GX�
pfܕŗ2�6��
�f1O��U����hV����U�ӱ�rXr��`ou��ErZ�e�Y1��w"�QYm�J��ot�*P;h�+*�5Q퍓dPwV(P hA��[U>u�2���s��L�zp�I��ZR̔Y�XKCRD�	bM�L�{�����*�m�@EV���kJƨ�&�t��%��CI�tqH^��7��:�;pe�c�.�v(<��U�E����ئk@Yi]Ú���V'3Q_@���[��w2j$�u���Z�"Vst #��u�m����"f��{d�ʏNd�S��歆���ȭ(ͺsNCp�&�T/�*9�FJeMhkC����.�N���D*�`�V�9`,��(��M� ��J�S��f .��Z���4j
�!����v��ZWW5�ٚ�*	*m� *=��G�*�+fCLCwq�t���*�m]���#�mI�O�je\�OS7w����r���p&LXw�2��̚��Sx��Z��s��e1�R�v{�g��g����2�yI1kE�ik��l+�W8�[K6���B�-��{E��Q*�f9��%�e̓;
\B���&<��R�����[�����ke�L�Ka���D��A�̅�eT
�Ɇ�xD������n�VC6[�zY����D^%%k��Uʵ��,ӛ�V�� n��m�m����q|i�[�]K�b���r�;)-�΢�������+I����23��)�*^RW��E�_Л`۬��س��%f\J�^���Y�;x�<��u��ZYM\�3��+�0�C��InSnX��aP^ܕu�L
�v�x��Oh��(7{!r����Vn��I��t�ZN��Ln�x��c0S�1e)Q2�5��y�Rl�#/i�i�4��7K�1ģ�Y�+oji�ݕe\�J�-���y��ĩ��fm�\���%JMu-�[�m	0��^�ˋo��R�Ǌ��hW�H�ԏX��dgaT��ن�<�dU�w����'s%���,֭�81eju#�K��Y�&�먳l1+�p6�"��ד1o�
�6�wxŊX�l߰�F�PCh2-�낭����d֩1Q�r�㔐�3YzjӘ�K�޹.᭬�2^�2�����hcuvv�*M�6aY���o#n��|+3⤇XU$��k4=ԋ���-v�̇6�K�(f�Y�V$d�ˡV�m�R�C&*-$d'v�K ��(��7�,ݬ��j�K%;��u>��"��MD�<�1�pV�n�d�R7�[b��*Rytd��wp���kp]�"N�\� 5���t��2m��X\41��emҕ��ʑ���fj�.,IF^�7�V�k�꜈�uxPՉ
�U�[|�;�(em�Ӣ�h�+o]�a"|v �:J�[L�fn�&f�D��Nb�7iQ�+h>��^�6@#$�ɶ�YDŘ�c�e�J��'�V>ٲK��p`*`���>�b�;d��f�/q��\c�����`Z�#�Ax��m����,ݬ˵���e�P��35݇.�ܴ���cE�٠�{2���H�`�&�@T��Ky�di{,(����dˣY�e�J�9�������"u��lh����t��(Q�) �Z5��ws�\%@�X�h`U��`��Cak3"чt��6(��!���r�бT�Mt$MMJ���v����e�5��r���\�ev�����p��V��{��۟P���Ez[l�
����=����=��7��|��k��
lKR��C`�u�:g8��S�v�a�Ě//�d�����;�[!r%ծ5y�·WI���{X�<.�g�����5��(�P��bʹ��B�ފ�-�Òry�\���Aa�=y��R���LcKW���pVe��pК� �`R��SxQgI�䲙����;n���6���\j���Ꙏw%���$�9����P��J;/���MD��u�n�cb(ݓ�S��6��順P�8��ۺ"��:/��琻�Q�&��N�HG�ը�`+Ob���t��3����l8�G�,�:��x��H�y�c	cC���e,&f�tV��@`8���*o]��;�9�)�Fe�B�T�tdlӸ
���e|:jT�Ae<7@�}��SJ�%1�(i]o�W8r�o|�yS#���wWm�*�����V��\֕q��vDZBq6����R���g7s��7/���7���nкC��r8uR��r�JS���0D��1�Maae��lU�o�;�3$�Fٽ��؜�egB�A���C���س�9�j��E<n�2��kN��N`Q�h�Xޣ%�ِR$��0�u���]y� ��ɖ@�4�$�u��x��7�)k�Х��_.�F7���˾��h�s�e'�V<��[��Zk��]�,q�B6j�sof��m���DMU�g�*�'K�A.tpH�i]9��1��4a��
�e��J�
��]KH7�uw.��Qa7+)����������5ܧVٳ��q�!T�k��U�_*���A������n�_l�Rk:����
y&S�0@��ƺZ�3��J�*�L��S�ac&X�c�}g�gfu]*���X�kEZ�b�<�K��M���R��=��׶o�:i���Y� #�q�V�����|yܻ�8�241LSc��cfe쑦���pܬM)���GY!���
m(�Q��X��*��+77 �s�Nb�/jV��Q	1�aI%���������*:M ��7�/'�3��9Fw��L��uc��]����Av^�n�\V�fvb�N�d�&:�k���r����FUx+��"��F��lh�K~���\9օJb��q��))�TYy�
k�a�q�P0��`6�%N�s��Z�neY��%p�o���Օw���IN����V�e��dc���V��^�-���T74�a�i)Qn��_fR<vV�:���=$O�����h����زbXJE#˥l�#Z��:���KJ�&�h�
*���ѧ����I�%�!*9lw�����O2A��ێS�E�F��,.x]�Ɗȶ��`Y�J}�yکR�y�9�aj���W����}�"���&ᤱ���Z���V([�Z�xDШ>{*�kx�]V��f���J.��0�$0�̢	��Q�y>v�)�����ů��,�U�6���ܹ��7��`�j�;ٶ��ù��Hk�e]�/��a7�Y��)WvK�1l8�9�ٗ&«��,�ue=`�򸼬�
����(�"Y�	�w�Wh�8;n��C`����T�'^<�G:N�
w�<k�%ۙ��f
�ǔ��{L�7���Ki_b���v8k$5���	��D���ué�4���]��"���ǟV�\J�6i���Q��#�:���<�nGh��%�������ಣ��A��7���7�����Ngýi��E�
i�mX��Pְ���L�w+/�+BC�zEOoG����(�&�3�ვ�b��3U��H`b�9�v�c�X*X�7�!��Wm�GC��..��	�m�;@��v(T���Q:�Y�ԓ�4MI���R+/����Eb<Fm\�QΣѱNU�	�#�@SxF{,�j3ױ=b(ڻ}��*�i f^�������-k��� ����_Z�%>���B�z�qdH�7tq�2��WP@j��Ε�b��>ZێU����Z�1]��8,+_iiv�BK�3��;�h:�}�:	.�:+F�!: �:�a�f�%�t�m�A�9͔��A}!��7D�ϧZ|�3�z�U�����;�v(���Oa6Ki�����k�1��<�kuIj'k��B��&�߶�CQ�YObb���dPV5Q' ��`&�U䧓:M��V�u�L���pp��:�k݂��+�Nם*�}z���d|�47.cԟQ��O�=�M\�U��5s�GNg.��{>wIT�������rA&�F�	D:�Z�M҉\=}8
5fT��:,��=�P�����<�`�W֣���TI6����읎�r��J�>�J��t,|)�m�\�sm�<hnL�v��!��S�aL���2�&ܠ; �H�d -��z�[�g�+ѳ��a�8V�b�O�gn��bm�a��1m(��Znfq/Uh����Y��*@�i*�#�Pfq����z��-�-��F���t���f,3J��i�@�bo7Qǉ�V�e��%;yuryC���;�
-�����2PINv`���]��ݦ�)G!c{%��i�҄�`loG'y�.ĽE�Q9Uǫ�F5܃X����o�7-@�E�6p���3Q���w��Ki�ũ��k�NU���`��u���Y{���^=�5�-���Tti�Pc+�7�2(�ܓ����R��g9;�;�
����x��)n8��w@39�F��|��7-NӜ )Vq��1-)����%Ӭ��Z���hZ�(IRRڔ����pW+�T8�P������y�_;���}RZ�M�NdK�D⮲Ă�$����B;��Ѳ^^�o^R�œ�N�R4�g^�-�7�К�Z(��#2�Ĺh��.ʗ@�j���&9H��G/�����ը��k�H�U��n�9���*و���������0Ԩ�	�m��]!�{��a��c΁A����݌T�G0#:ř�����샐�6�v�PE��gS|n���-dm����i^���Z���5��m�{�:��u>v��vNmMWy'>]CiM9r�=Q[���;=�՚��W]hqr)!�:iIם0[��4;����*B��&��-%V�t3a�2㡌�1d��j.��)f���ݢ������s����Wi,\5�bo��\�>�뽞�JZhr��x{�TLL��엎�WY�_6�%etͭ�h�"(���-��Ө�5��L��Wa�V���Q1 �2�47����a�BSV��[7j��Y�֓�ʜ/���;va��d�+���8��I�ͩ��>����9�vf0��LN��c���*�g�6�Q�De�w�[��ɶLْ�|(�ÉBI�9���\�Ŏ<f-�n��Pq�6�S�ltU����>�R�,��鼏ؘ7���Āof�Q�t�)�_U��#��*b ��1y����Z8Bͺ�=6nqͻ/��n�@�+������x¼���tL��Jf�q��^���N9A-=t{>��.���&�];M�^�:�xuq�\��g�V��y�L�D��6r�f宇G��ػ�k|w��y�0nU�L	͜�hv�zY��&zZJ�<��C�|� ��{�l �X��B��R�	�-%�V�|;'n��pCe��[�,�
��Ԥ���GJ�Hj���Ǹp���VtZ,�����ZW�� v�C��L�<��L�4y�e�3�䘊�{-�	�L��r�U�,ܮ��53"�ntZ*�P��$uc+}�E�����lYT���u �n�M��]���/D5&�F�wf�.ڃ6f	q�l>0RV��c�V���	���4�%
�'���y��(j�s"�[�<ل�`��R^-�^��v�;��QÊc���9ˊ��$��@=��vY��:�jC���Ʈ9��Zg��'@V-�"��̨�WA���X���b���a���zC��rVt�r�-��=w*]��<�T� ����5݈�P7o�!�K�EҝP7J��>Of1@�	�=���)>�,��R���#R��5y��١�kl(��LӶ=9޻���j뜷IVV9fe��3u�%:���YP�ۜ� �*��Qe��f�X��Z���q)�����1jɶy]�U�F҇.�@D<P��k�ꊬ7Y/\�e�R�SN,��A�'|�BśB�uI}�7e�a�}c��,X������(�=@,��V���2�#[x��>Pe�,��gm�=�ç�H�@�lrv�P�w���(I�O{��Pb�=�µ짝�e�
V�{�@��0���C\�)���yDc+Qb�v��T4�Ym�š*�F�ʷ�_*�v�w<޳�=���``!C����*�t�k��+yIy��v�*�f�	w|s]��k���W���\��8��P�]����y��si�*�96�u����hKR���H��x�m�5��U��[�\^�l����rY�m1F;�Gl�V�6 �C�1��hre����=WP2�)mK΋J��;(�|�:�������ˈJ�Z:%8:�Sa�������ܧ��y�(+�FU2�Z}t��mկ��!r���z�WJX7�7eْ�'b���K�kJ������
���V:�w�l'JU����Y�7��w�9�+lT{�T%�v{���*\�)Ij��t;�7`��VP�A�iIĬ�xQ��P������V�;�͓.o!�$���`��yI��*�a�[�:�ȧ0&�b�f���U��K'N�]�wlZ6�K�ޡ�	�������8�Z��Zb5�B�r:k^n�.XR��×��e�|l�c3�l��#wM���Ph=lp�n�mkt
��tA�o*B��蒶�����o[���ҧ�5��,E��@�VkEz��u�T%XlX�K-���;����Ր�<�Ѷ(+���ol��4vwj�!��Z,S��U�w���a�nT�t;X��/�����k.H��� �4(��{��Q��o�Pm��2���7�Lw��r��bћ�)�C�.�VS�]���-@��$au�����Sf��ڍOV��K�N*�*ɻ*+<� PKa,�n*���̕����`��:�a�B�cy+��ٚ.�"G��X[F��3o+�;�
d�����+�S��2$X�Z��\Q�Du��@���6`1aU}�\-���SRV�Z�4��L@t�=Ӛxr���ة
A�����R�����M'>e�u�4r�,֖ҷ�V6��eq�f�R�D��j�7��d�X�u��:����I��[iU+�Wp�71�B'{��kV>�D���i�s�W���p��k��pv���}yW�,R�o��%	C'��u��q��:I�R�QV�	��^6]�5p�]*���]��� ����b`�LST�sq�n�v��� ���s��kU�lJ�/�Y�*�Fa�$
��!�{]��D�ya�23f���8sP��^��j��V�<Awa��v�[ŇV!y:���c��-�۵�-H,��;o��~!�V�^�Q�.Z���8����c�W<ͯs9zώ��C���iG�Cch��5F kk%�U%�{X�l})��{o��f�*�ݒ�?�ٷQIA���ڋ��z�k�D��VN۳x�9��s�CX��h����z^VA��%�Mw�x�_]cհ������J���!N�0y�:?�7Ni�V��p{dG�����g��@�INrP����9��@z�M��t�V�w!���y�z%Ѝ�rj��v%�������v;9�VĵqZ܇5�ݽ�2^ܾB�,:�k�|���nvS�K�8�S�݌�h�2o8�X2��W;;�N��9�;|r��\�O-�]�k�[��u�{,���N�ZI�W5��m��/�em��ch
h�A�eAA�7�8�#�3;
CC��cTc��q�+ܔ��hΎ�x�sd���K����ԥ���uo"��Yy�m��kbǫo�Bx^�N:�+U��y.u]R�8 &/jUҏM\g��B&<ǉ]f�y��XtIC�rQ�R�-�Iu�j,uN[���v����a]�+�v�:٧!	q]Aӗ2Q �Wp�Q�܍1;f,�GeYݙ WnՇ�cs+mkq��\�X�P�{���[W���z����88'�]�	G�;�1��2��Os���H7%"R}W��5L���[����@�ݰ&2Z�wݢ1�ۤ掸�SK��eXJ���\���}r�xe�T�ҬNr��tp��S��;g�C{��)mM6��M-=�.�5���3H�z��ǰ�9+�WZ�5�޻��Y�f2�0"	�ƒ�k�Yض'i���x�*f��K��a��M;	B�}2�-��k2R�U�;2�F���WL�d�*>�뾽��eܷh�ڌ.b[�$�a��n:;�c��Y���ۏ�X%R3�D�N�YV��[�ǎ�c5�����C$�;�H(9�=nҺ\�W{�����5��У��t�>���F��Rt������vd��k+R7:�ܪT�C{�|{hd�Oh.���T���w;U��6�6��KOG�ú��H�2���١�e\B�4��\vCY���\XUvaq;W8�G;Ds_K �]�T����u�+(J`�Bu�|4��e=l��^\�������*�"���`�̩�����w�!��qm����*4lѶv1
ꙙ�[�d�v:�l�gfV -��Ҿn���3�5\���.��F����9��>�sչ������4s�}��OV\�r�G��\鯩�GwRo��j[l��;�l^�:�1���ĶN�*\������0`�y-t���rb�d�F�-�5Ƥ٘��i�k�
R�q+W�ׂ���XzDN�I���[�\۹]i9`ftj�#����d����y�D2JS�������k_߿������l6�}���������������г�ߨ��O��'&RfT�d�m�64W0�#w��U���{K丫�9f�n:R'R��<M�5o�t�f�� �P�x]W�|���j�v����Z���L׽�����RB�4q�U.ϴk8�|-J{IŮ�+
�@�j1�O;�{8��z�)�[�0nW��OQ	�ڼ$۫�ǾB1��-΂Q��]<42;*E��b�7(m[�wvN������j��-��>��(�9�;�J�F-��fx���@��q6�j��>��� j&'GyZ���VI2���8�s�۽E�v�Q1S&�\3�w���<W#|�L�Q�+%_BŶ���R�.7�/0VR�|,;Jd�ϝ�w6�u	��49�B�q��X�ؠ�_zH�ڳD�� 9���P)cf٧Ϩ�B�Y1��C�0Y ��z�¡�j�[aY�g4��d�F�sІܳ��ͻ�Yt�;�/�w}��X e�	9��u	��tT]X��pƞ;�$�r�a{�˾����<S;�*�kxqι4���uŰ�ګ����K��9>������A
�Y����롉f�wKs�5��Vs�W;bl�^/�с. ��CG	�e[r��_K��X��Gj��T/qN�@0�v�U8�R#gY��L�tD�:�ڎ7i��{{,n_gg9��,�1X�S�y��ʀj�<��=�������|�k���p�7[ݽh����-��T��"a�$S����^��t鰛wij𪎲�8�y;M������RWʂ��9�+��TCo��ǧ���Y"!��hr��c.Z�h
��XPs�r>	�l-�z`�	�ʠ�K�[��%-��`�͔�:$��q5����j%�������d�۠���&�!�x7 �E�]ʼj�� ���-72怒�Q��M�B�e��F&Dv�m�����h�[�O��u��_wsP�ٚ�J]tm������=�\�Yq���+ӕ��c:�����d��˳V��k��ټ��� �Y9���NX�Q�M�S�0���Ű�X43���*W6e^�YN��:VU�5�<zC#��2���*8����_��`�ۛ��#��k��ƒ��W�[�`��q���*g�h]��Ν��<�^��Au�Lzn�����/�=h�+cg7Z�"�H�ߞ�הre��ڎ�V�Z�������U��	l[θ�}����3a�r�ȝ�,�����뮶�_+���g��P}[����e:m�
-�z�]��3!���EM�
;{;�\l�];\�8��u�Lb!J��KSU'�;����t���m�ɔ%1�f"�ec�t��u��]4iPHV�Xla��l�w���E�k3啥���-Ÿ�ϰ��0ؤ�r��7� Kl�������ɦ%��g*5J:� K��=Śy���4#�:�J A��F�e�W�wp6Վ(�y>�J��]�`�H�B�q��B�)@�4�~H��>�k�u����Y�D�,������]!�辻�&G���]%j�WAkFvl�>��s�eg+bvA�=��S�£��rk����ҍ-K�#�RSs\�jf��CZg �����W�b�#�	��.�7"��ChG��r�L�{;��6�`�0���{Jެ��@R!�a:AoGh\ŨmG}]d��Y��Ƕ�i�}��f�5SȘ9���n�����9.�wkr��tkz+[��dΧ��p�$��Y
�V���V7;��n��:�[Ύ]vj����)oki4�@`٪�L�G,'[c������У�=4���B<9e�Wnw9㢶�2S1���#k5d���Wx6��⤺� ��N��de7�9��x;Y*f����D�kN X�W�Fq��N:ؔ�{]֊KbE�q��	֝WC�;�n��9�2+��*÷��,�WO@�jn�,��N���-3L���V���������,N�m�t6�5����b�����xA�T.h�����]����]���S��De7v�
a�Q/o��{�(�g&s�2T�i�A�;aRj�̓p� ��r3��E*�a\���.s%ؙQ��n�[Sr��|�
���WJ��Vû��E���c
I��C6ޓaS����^�]d?���� ���G���������=(h�5����4q"�g5-�;!mSuT�����j�Ѽ��F<Y2g�35���b(�ʽ�NzyWn�܁�7o�]|��Z��Z���bl�7eԶEoQ��Y%�D�zUd�,bTqRĉ�w�#���d����\A���d��A�Ϲ� �]T�NQW[j�Yɴ%d}���q�緛��4�e���zs���q��&��lee��X��Y��O:�R�������t��]��rP�Q�(3�\�0u9�H'"�s�ތ����ByJrf�;F�0�^�P����_97�2��xEU��V�sBʉwΎ�G&J\6M5�ʛo��K�J)v�	
���1�E�V��f8���G
z�5-���(ǵ˕��:�s���&[5#�k��2A��m4��#ߴ���P�NWv��ec����{�ჾ��9���9��)�vM$�(���+����&���I`�*�^���^�ܻ�8fۑ"�uC�^vww�;�(<r6:�t��$�i�wA�a�w�N$W�I���7��*��y����f]k�~0(�yس�x��,��yv��,Z����U:=����v�Y����ɃE�N���e�%�Йk�jT��!�` x�T�^�����]{�fθ��m��rľ�r*�;�&VJ�A�`��Fy-��ӑG�����WQT,�2d��0�n��F��6�K+Pn!<9Y����'�Y�ѫ�h�6䬊Č����B��B#ϒ��:�h��@ᬮl�V;d�[��[�tH�4Z*��+F�msܬ;A��v�e�Eݛ�z���u75qUq��Y�n��'�{6�fûZ����;�ҰvL�<WSt"�`l�I����F�[p�M.�b*�z�p��٭8-�l
v�>�J�Մ��Ib�ER��lc+p���5;Z�Y���,'V*���f@S��A3o0=��ݰκ.�Xx��(93s;�����Yx&���Z�S�]��4`�J��}j��6�;btW׬�Q������y�M�k'$��t��	l��3�����Ma�1�p�ӥ`�}�)�N�}�['V7U��#Ӡcͧ��4[��]̪�H;%�_MP�i�55�!�f��t��9Z�b���O�T�6m��u
v���2��/2�9wsz���B��T���jYtn�=9PEÙ�p/��)�� :jm��W}a)�	ڼi�[h�3�����D*lj��X�3n�`H�Y��R�,KM��ތ�a4�>?v˭�#��P��ԝ���v�e�c�|'��o�����w�O)�[�1���T5&�y��V��m�߃�f����d�n�󚱂�%ԁìO�eZ�6r`ۖ�h�˫т�J�5i�
��Q[��暎�r�u�L�`��.�����y[(��9����a� ɴ�ZcX�Ec������|�6cgLQ"�,5�v�uLi/P�n:��|X�C�dUҤ�%r}5i�а;�d,����M�5:{UJ����ku�d�e��P�NM}�՜{R*�2^�ۯ'��<�����Yy���ץKA�+��"'[T�E��5u�����a�"�E�%=&��n�tz��..��6�E�桴��$�����{g)���tCZS"8sjQ����
G�y(�{�n,n��@�q
h���*q����!3Z�pWusv�ب�����R�@S��FX���	m����e���ު�����UNh"�_0��ϸj�D	ܱ
r�,�i��巅˽TУ�ۮ0k��d�|��]ƙܼ-ι�5q�Q�U�\�U� U��H|��͘3���6�8����ƚ	Vwcݣ�	Q��쒥�I�Y[Ij�'��S�[�B�_:}��Ŗl���y5R�{JJ�@�-+[eR��-Vx��St�59��Ⱥl��A�v�-�#K#��}��F�y���s�d����ƥ+0��5��f���EP9��y���4�urʹ�vn��\EMp|�E��ts@ͣ-��)n棧z���$4��%D�a�S bQ�FV��Tl-���g�6㥪=͙���h�r#9N�@�%����u9��]���r�26��(�q��
����!�97dqi�e8�j�T��6)2�7\"�eSղ��=5mIM��&j��'k`+�o8�`��
��	�]��۔����wóY�w�G1�r�J�X_e�NG0W;L�yK%k��<ȥ�<��kn��&�_cI�e�n�k��f�t�FI��r��te,4"�ނ�]�sR��f!P��L�W\[��[�+�-
�KeM�G;9��y��Z�u�ܥIw86�{�`�G�Os���ru94ԺR���+��I�Vs�7�T5n��[=1 nX�7�N���ӼЯ�IQ��p|��(=��-�p;ZF�L��[�N�R��Af*���ʰ�V1gVˤ��W��c��xy �*0Z��r˭ҹ!�n��M��H��w��ݒի�Ҡ�ia���܂[�к�aa�kZ6��rY]`�gD�]��U52����j��i;�*2��nm��t�9K+F�4N�a�ྣXm��C"Z�Iat!�qn�R��˕��\��ʜ�ÆA��-��������D�m��+6�Qw�$>�HT��8����I�"�8h����Iv/�R�Y2��#(B�M.�[԰f;Q�����]�̤��"�Z�5X�ְ"N�97F�M	yy�N��!J�T�*5h�h�3k��S����Hѝ0�^��I��a'�j8�a;"������a��-e����	�������SY�_c��ۚ�۹�p�4�Q�6IJ��Gf���R}{P�Б>p�Dk���D�E�='ы������z�+���b�l�EI�4塎�n�-��rp3�1� �t�)�A �rs�����Z�
�r�NȳU�J��ay����檶�pV�O�n,���1��M�~`��T�A&�ե̝\\2bZ�v�M��!���p5�o w1��x����yNcI��AꛁV;7�BLX7dJ�9�eڔBD�W���\ؓ�i����, �\��c���N8������8dU֡Ċ���v6��f�`V*3�i�fSi�����":��h�Lk:�o��0�f�����j��t],����o�Z4�5��s5c1�Ww��J����炶Y�R]f�_ch 4�S7�%ի�+�#/��+�b�bXw�d0_lEihӪ�:Y vE���e<k���	��Tzg0o���2�g*jۖ�J�q$(�t��<E���E�{ٵ�a�T6�ʕ�dŏC_2�\��X�uU���e�3�F����8����Y�A��je��p����u �����M��-��U�&��)&]`�i���IT�X=I�!�F)�R2ξ�ׂX�[�}�dےܖ]�Ҷ�GMm���HO)�Awf7�ƈC[�ձ��Ү0�֯�ņ4�=֊��$�YQ�_^�q���w]��͕�P�m��-Z�U�Q��Ѧ%|��WyX�v�6�ZOi3�]X�iO��s�����cܳ�H�I֝e�F�*��v�pupb�%ܝ/"���L6�ܡL��aw-��P��
��B�i,��Q��kfʒ�رsH9.y�����e�wb��0%3���K�����a�1����G���L�������HP�θOVbW������JtR����F��SՕ�&�rq�d+�Qy��o�q��4�k�H͝��m���	�XKTH�X4�\1PRI�,k6�ȳ���,�8�4�&�;W s3ј�����w�냑�ǝH���;y�p�fE�v���$S��V:H�W)G���bܠkuZ��P��J.��1�X�#g���y@�53e0�霛��hI4��oA��p�YL�Pm�W��H����\8^匉ʸN3�!�3c�׌�d��f_J�9�Cn��ކB���좩57�z��T�L��p��&���v����pP��v��9��Dy ��؎��ә�R�sKh������u�F���8M����ͺ�X�`���MV��o��n*6-h��찜�W]]�N��i�T8E5��e4o��j�ϲa,�n+�lT5r���w]��+�:Ӥ��e1�L�V�3J5b���ر9PmwbD��:f��yd�I{lʰ2ق^�tM���[�T�(+b�ʏN�S9��TƢOf��������DiQ���Yݹ�VQ�8�<��*�\w�e��� (&d��6Ť\x@��[��� ���Ztf[���h�N�l1�*`WV�4.��:TTo���*ު��P#�:5�j�~":���C"(�����hE���k� 8C�w�T�tw�Q��M�&���m�v�(<�ccxhW̍F��SWvAs����m�k���O���c ��0s��5���2a��oV(���r��YN�gN�ot��V�%2fj5�F�K��/�y��uQ"Ij�PX �EQ���sz5]�F���҄�9�C�t�S �m�SGsn���`}t��t5�V���T���yfH����0"�iCp�E�0�f���nҾ&��JQfҏ��-/�^���oR�t�Rt�W�m��a/T�cj�0�Z%����&rY.�d��]�
�¨�r����N���5eq���yL�Zy��[C�rR�{,Z�&k��4B�T��n��9�wttY��7��*�iWt�p�m�u�Aip_���W�U}_}���/c����줂1��k��1��R��:k�����m���e`83[���]�B<�Y�{K'�`�R��#ù2��t�v��PJ��8Ԥv��G��J4���+/Ƭ���egf���/�6�o9%j;��h�Ά2�r�ͦ�e@�(�ki��B �̬ܔ-g
��n���V�j�v��7N��T��E�u�P\��ݖ�K)��z�v%��	N��K�Q�+ⶑ��Y�I�DG�@�C��ᖖ�s��w���=�Li�V�3�s���-/76��.�mګwe�	mp��Z HLjf�<�a kA_wʰJtܸAUN��ٍ)�L�J�tHEF%؝٘����w/������ ,�7$�&�dv��(Ƈg^9t�J����GR�`<FK=,�ICQb@�4��8�M�֎31�{ع�-L|7p>R��̥j�IY���'�
q�y͌���:��mr���ڙ��|Xۤ�J˂gnĂ���gC�\�^TvK\��>U	Ҏe����D�3�r}�X�Ή�e�L����SH�6	�R�<�q
��"���l�� 6�ys�/j�����G�;�tZ̔֋����co`D婌:�����[e;�yE�U}g(���vq�Ց�˜e\���a�Ѻ��	vԊ������q�ܘ����6G�n�Գ�Q:�u��]JX������u��>w�q�A�#�TDs��U9���%2*��!^A
*�+��4S�w"f��EPC���ɑDD\��vA�9dDL���mȲ��9UNR	��̠�Ȩ��J�EUQDr��YTQDp��E3q�\.QU\���V�\<BQQ�\���p��Ʌx�*�DG<��.�ʢ��U*�#�r玕Ȣ(9QAȔ)4K8�C�:g)RQ��BQr8DT9$%҉�EDEh�t�*����QAA"�q8<���9W�"�QEY�Xr���Q��+�S3dTJ��ee�+ZW"Ql����(�r#�eU�����,:Us2+����#����s�]�w���E-պ����uң@&����S��LwZ�g$����uǮȚ\�@2���L���r�cˡB��w}��ϔ��-�B���@2���YZ"+�"��4��u'#[�t9g�\.����	:�e=�<���:߳�F�u�C�Z�j�ݢ�7j�:�;��uҹMb�w�*[���!�2&�;�Yc�˸uz�d?c�Ѱ���r�p�b��k�b�9�9h�DN�SsA쮎uVT��^`����{}��)�t���G#�x\jT�֤*��ӣ�D�����׉�Ξ�C�Z�����5�f]*�0���S�m%��o�3��
�������59n�}���\T��GM�ͼ�w2�"v\��]�*uby���ƘYw�etĞ߯�*�(r^����sQ[8G� $�}����E�N`w_�} �U�x���R��`�-հ��Q��6���?p�f�Kĕ��Yȭ~�\1�l����ksjw�x����a���؜�9�f}��x�b���v�j�N�r��+ڸ�c�^��G�wI�~{$�껡\/�j�vT���a8��.��U^�q=�4ϒ�[>*J� `D�'L h�I)�_N����Q��ѳ�R�nL(�G�bj�b�I�Y"U��H*��q�����-0`Wb����z�M��Nb95�LB��N�]�0e�̵��E[.���BD���1S��o`��h�u��i�Cc,$�.WD[��04%mfW9,��^r��Ɣaz�� �����%�g'��������S�n�
&d��wq�SyYTRC�#��`�B6�u�����̙ߩ��d��s�	� d7p4_�^/Y���D�?4��>�v�o�՛�ʃ/��B�+�;%3f\@n���%78��Z��f�[}/UYٗ�� �`�@���8�_ؼ̪ػ����~����)2���=��Hc;��<��ڛ���@%x����S�����CϴDU�@��DmTy�ר�
��U1<������i��76���Bn�矚W.�
�2|uѫ���Z��􊧳tK���թ�Voij�p:_�y�6��L�;���l��-`���6��g׹Q��{���"�=�8Ҍ��hFθ���g; FoS���d�­�s���W{W���o�P�ܻX�xm�]G	����I(�	��*��8�֤���ئf��9�������\�u�I���>�p��?t�8�}�[��Ϲ�Wr��Q�����fBoy-��35Y{S�*y^Lƙ�qڬ�%n���b�8PJ�V�����Ψ�J��uЫN;o��Ɇ�,�x�������6���ޭk��8v�]&�u-��U�I�)��6DH�|<6��t�7qJ:y3���J�N�j�B������eD���p����6 �1�S�G:���.�Use�m=�f�e�M�'��]e���l��ت��g�"��jmY	�zG�Ϲ���0���7�Ȫ��0��-Q�֒%��Vv�I��a�V𪲖f��a/zXAG�^����܌��XZ1:l-x�t�"��	!L���mr
.��T�=�����ma�춼gEL'_gzx}3���t9�:�Y�±��&����5��;G�Un��J�1Jf'Q����CC!v\S�oL��*s��^�B69����ё�f0���ʦ�y��Z��Q�r�?Ar��J��X[�_�u3qN��KϠ���{K��(�=�n����s|Ԏ��
_P���{������������!��$4yi*h������7���{���Wڀ�=�! J���n�5�*�2��6$���R��]���u�q���Ǆ�>S������q��QJ�҆��tS���0,���o+�eW=����4�gȻ�3T#�O��#�+�.�JiF-K5>���(V�F)���"g8�cC��u"����]S�-h���v�c���g�/kHx���G�I�c�&�5X�)M9>��4v��}7t�\�l�S!�>Εg��E��8Z,����Q��;��!����{����2�J�������CVﲏwU�|����v����F�Si_#�(W��{�K�ޑ���y-�$�0}`�>��=�}�ǖ=O�o*Ey�>#<[�*S��q�N};yNr
�s�ۛ,ANy\73@��U��b��p|"����� L�7�Q�u�;���V��Y�c�P��J�,�m�,��H�8�$2��ҹ�����f��*��c���p�>	jz�$�������J5yX�P˿W���f�_w�}��B�Xu�F�ĸ[���Y�1Y3�<Fu�n���U����f�؁��VG
�"3^r�t�r�
1��E)*���17��h�Ș���ܭD�:��H��:)�X��u��8:���N�/
�t�;,�;���VӸ�Z'0��[����!���4>(H4�>�6�g0|�+����t����滙]��р�J�a{PM�Y(?�W�s����@�&=ش���n���2)�.��[�Գ ��C��ץ5�;��lAj���>f��\���d�� ��K��
xk��bb����m��L������v�MV �tWۻ>DQ��H�g�O��V%e.;i�q��Q/��6�.	׷��W������>y��ռ:��J�hW�R��6m`���������������\Q�|�G��Ukx�����P���`k
���G�NV�?��SC�����Ќ�z���C�B.�C���i����,��E���P;�Dq�ْ���{D�F�4 ^»E��Z���l(Z�%��}-�s���V$M�����9��
r���G�@.�ʂBu-��[%�K�Ԇ��9�tR7`\�&�D_�u��dnSB+!R�9��s�,�}p��ߢ]9��I<���:��[��VF���0��sB�y�?3�H6,�^�z�����-��D��dN�Jhc�<L��gbD�Z�����c����>�7�$�ݏ	r�*��L����ĭ���!�V������`y���ZWp�b�g�ϊ���]o���y�]+4o�?���A�Y��%;���l�ynmX�$�QkRi�]�k��0d$�i�<O?����"i���3}�k���ڸs�!���k�����y�X�E�g�M��%]���U��u���e����S|����z|'���_G�a�+Y��X��J��C�eoQSt�E�4�r�&�f����nX�B�z��j��.�nT#1�$�*;�QNܬ��}(�r��[*udr�)�x;!m��j��ܘ�-�62�]_\�j�`yJ�����(�q��Iv�
S:��:�����=:��l�$��+�ZUq3�*�q���|+왞�Y���_b�������hl	�T[�/����S��{dRy����w-��&���K䕤s��=�c��A��n̍��\�5�a)����n!��5�6*W�?�Q������'\�{_>ze׮h��u���)��a
z����2�����g!Nh,� �0&\�
y��Q�#*�f�"���!]#�|�]���.`��A\�!����|>��*�Z�4t�!]�k���+,�)td�S���o�MW)0W;2gi��d}/:��u�n�h���p#���Q=�V\�^�RWG�'0+J2(�6�2����@��)�S��N�O���v��7=��"��
��OD5�^T���q�.��el]�_C��R�����*I^�f8bO���*8}/�~ `�`U�r)��~U@��~�d���l���1���@�'W+N�Tew����j��m&�M���׮@��$��WL��N��/�Ѽ�K��X9�y2��3`��J���h�^(nX�W�ٳ��3��WFr�@������쭱Bj���^n���.3�ԋq��v+ �L�$�Ău��skBQ)S�}�u��4n��3{�t_�!�F�bhc�K|�2㧺�p����A���4r؇�IZ�c��Y�a'��2>t3���Y*��Xzʳ���ss�r�0���{^��j����g+ FoR���d�­�s��ژZ��;j�*���;�U��n]�\�J�|���96:���ʩ˝$���gW��oE��4�]/)�Z���̬���Lzv}��N	+W�̅WYg��z��	E.�=aW���^Ԗr���tL)��9�J����)����la�fmKB�-K�O�-+�y����o;j���k.�	�֚s93���,2��s�ј�^u�}1DlJ��4���A,0u��S���aO-���̻ќqߪ2r���_�8;r2�ahL6
x�����LШkl!W��^o��k�P�L{Ϯ���t��5��9�#�;S��i��tV1�a՗�ݞ
�;�k8��.^�$�+@T��ԫ����y{�B�*s��^�B7�N�Y3q�������b:U.��!,T|7OI,������P��ަr+��0#o�n�R��S���y۬*�1���i�J�a��H�ƪC/9m��\�N9]��ΰ���é%��I��	U�ؼT3�RR�N͇�����O��A�7��s�#�v���靹��(���4��:k@j@����4�N���x�g&��ƹũf%�?8]�7®�ْ�i��l]����cP�ǒ��t���7�v���\������[0��>�`ʯs�((����-wM ~c�%��ǘ�|o �sW�}��8u�! �8�n���Ü���^��$�$QJ���{��˲��Ky��7�������_�ip�Eؗ�:3t"�I<1����f�:�
 ��͋}�K�y��A��+�qoi_#����뿌��y�8��uG!;��9n���-D֬<��eV�����E��b�{p,��>W��½����qxJ�o�Hk��u�r>�)�Hg+=�kl }�2�u)���)򻁩�v�Т2I�L�e��Uݭ�:N��t����YX�����;f����g�#8��B�����W��=�j�퍕�4��%�ɪ�r��uDW���2��7:�gɬ����:]�T�R�w�����'�M����3G��o�:����� f���P�唣��8�Ғ��Oa(�W4�b�\�<v)J�B�1��b��9�e�[���Sm��c$,57��e�7�uC�!k�^�M�2��{�_�Fk�Ѭ[和��^��o+����"�P���!��iV[����)_D�G�)��ƺ���I��2qUr��)0ìY<zba�t�H'T�F��걐+��\���ּv� �雌P��dBt�;��2�ړE���w�̡���(,��H	�i��6�����w0���c�T9�����[>���nٍ�.q!*��?W=�!��GK��O2��=��u���풩�����T�P�T�-m�[�h��cԞ\��n��w���6�˱�N� �^��q�ي���_���j�z��W����^EdU9$g�T9<7y�.t#1�5<H�$hXr�G����@����\�.b}j�a]z��j6d�'��ؑ�I�f-����Щ�5@�x)Y��k(D�ݬ�g�n�D��ˡ"RUrm�9ԅ9xqFܩPX؀#>w�]�:���N+�{�۴=��� =X��0�{�[f�[X<��HEV����T��f�놕���辳��M��-.�<���:��ə]@����\x�vԮ�*7'1X�c��s
b�{�Qٺ�3u��Ŵ�n�Jh��\b'r�G���:�����+��t\��xHӔ�hQ�=)McCf��SڃF-�n�����T��Y��ǳ�e��-�k���;)�<d�4�8��%ؕ���/69C���ܥ[�uq�$�-,�C1r��E��{�<w#kQy�/�u<�t����S���q�d����X�8��Uc�1AY>�zM7]�`y���i�k�x*1pڳ�]��]=��G�WS�q0������O��ٿmL����%�OBkG�0V��iu��bS�J�;x{6j�e0�<�6|��~�+�OR�=�k���ڸs�!��w�N��V��#���2uM݊	�iE�f��OQU��i�l�0����P��o��S��<�s�v��\8v6�Τ���W/���8�<%Ĭ��}����D�b�خe(.�~?hl	��1g�ksՆ�ꏧ�[���]OfK��s�g2� kCY����9���2�j�����u"�W���#d����������-G�g��iV��%�/����dg�ۖ��c�\�N���YA�q���䱐X������S����
�P���-�glm{$�7tߨ{7Eg�SC�]w�m�	l���@�:9?e:�0n��TfɽmGs!�˂�L�`ؑ0�	�U�
3��2Q� ���{��#�=[dS�Fx⠍V��4�(�Ǭ�l�����D-h��Z�ʂd��a�y��Xo&�܍N]�OJ���4�Lp:Y��ч,gqRk����6r������7iA`!(
>UJ�qֹ,f�]l�&�|8��G��vhŔ �}
�|i�N�c��L�*]��lgK����<5�'Qs���Z]v��u���.}ث(η��l�[���j%]8���j�ۻ��
k�vY���w��hՁ�,�y2U�fƜ�G�-�<y�C]m��]��i�smK;Xm�Ў���q�����.fʊ�Z37�6�>Z>�N��s��!�2��WK��Η�:ǬAl4�eΐ÷-=�^RہP��E�R�%�E��t�����u�1YԠѐ�Y��Sr�3���{J�vi��s�l.��RW+7U�t���; p�M:913~�c$�����x8{���R�)tz:�����⛆D�*s�pRS�Xy�*?%��W��p�p�H��(�m��:�qVc�U�����R���{�����Bi:"m+���:]�,c?���օ�;b�_$Eu�X].����0Q�P����𨉧T����<�r�mJ�
Ϻ#�Q�K�o%��4w jQ/�<��Z�;�u�V%�R���1��c���q�l�1��uuEbEL`�XۼXtK��� �a�G����c`l�A��L�7\�7؎��v���.V-N�L"�6���
��X��U�9*X�h=�c��/��t���B���d��.���=�"���	ً��4�ܓ�}�:�D�΃�gb+���:��ޜ�+�I��\��� Iʧ�+��2^*"�6qC�Y.9�m�nl�z���R����BvL��숥"�oA�E>���U���)���8gM�sp$�;s-p$v����(bHW5��T�]��W�K{�8�9I���(j�\���� �y���9�3��3�*��x�F�S�C疞�@_w;QB�56=��fɂ���s��T7��醦�`�3��.`���eS��:5�\���Z�-��6����DΡs	ۘ#��Y��%�@Ӄf^�U��;ZDi��V$�'eGO 	ѽ�(�{,���f᫶�[�K37�̹b���t`4����I��;.l�(�Nx-�(sB>!c��G�
��G|[ѡ�<�=��y�c��Z��2�Uخ��/�z�AH%��h��5|����p�Hf`����gbɩeZ��fڂ���_I8p�V�Va��|f�0��%\5_d,��2M7�B�gR��B2��Y��O��Sj��l����ÔCV����F�x��u����4L���}�u=��F%=��:kE�S�񃑀��hIK�ںʇY���ڷ��N�1I��A	
�{���Y&������O��A�~`Q����6[)[��{��:�yR�����/e���ꗷK)ZSz�[n�dsw�U@ >�p����R4"�4�E�"�����:t�AȃA*U����As2L��U�VUv��\���*1��EEȈj$TY˧.T���(�ek6yK�EU8��kB��+4ʂ������sZr*"�$�e3��đA�TFvE�NQE(�EDTEZ�jd�T�J��9��p�,aEDUd��"eyND�G%J(9\(���`UpԮ�gT�`Gf�"��h�*��ĎG*��G*���PQG
*+�T�r%*�̨#�W
�e\���\�sR�H��*.�0�S"�P��*�ք�9AQ9qZcH���1	D@��)P��Df*#1j�Fj���N\�D��)f�4���(IDT�8�DD&I�R���UPT�U�*Ј�<x�0�c)Z�)�0�5����~����y�v�i:-�����,�B�a̽z]�SS�f��u��jW%F��`�T�wItЩ���,r�����;PQ�W?|�?w����aw|N�lt��
�A�"������9F'z������L/��~�ۿѻC�|���S��o�\��x���ϝ.㴁���'���;?9��1�*<V��w|��վ���\���On�N*oK�4������g�tc�}v�vy����I�I��
o˽p��7�A�O�nr1;�u�G��ݧ|?|�t��Oª��yX�� >�+��SH�J�K��y�y�h�x2�iYx�"�Ͻ����ߝ�[��oy�oP�;_��<��o�N:�A�ב�C�����Ǐ.��v�x������p]�E��ԺwU.�UT�r7���[I���w.+�>�2$�~�~����<����q��|�;M��Ϸ<��N=�q�y�6�;q8����{c��7�'n������q7������� �l�̀8������>��;9s�F�Y���3�}��Dz��i�~^��2O�����ߝ����.�[N�7׎?y��>&x����|q��&￺�e=N���>o��}�'t�'�t�v��13��8C�@dF}s�x'y^�j���7> "HG�R��$8�x���Tt��� x��tp���㾻I����v�v�qP�����7�O��9��G>F'z�|��}���>��i���6�7�r����ʢ2f~�����+|�>�;x1���|��q|�yb�1"τ�z�h|=��z�q��C���I�]㎵q���L>Gλ��e�?�����p<I���-����7�N����}������=��A#kLlA=0|껂�ʺ�r����,����i7������>��\��oS�v�I���~��z��?����&x��q��x�I�]����v��	7�u���ޡ���o�\P=I��O/=;������r��}w������
���*�����q7w�s)����u���[�n�?$'����t��i�g����t�+�gq��;�z���Ճ�x���w����I�O�i����FH���7�>�s��n�Ϡ��9��阙�S
b*}M�щ޿79�F������~�۞����~��aT���z�~BL?����ڻ����N'n�<w�k���:x����&�����u�9��?�[y�ʜ�j�j�X�4�G�RM!���c.  z�7��*u�y�F��ׂ��nF�8{p��r���I=��
�k�����l�ch���e_ �dVo6��&����B��Jo1I�OӦ����̸��kd#5V}�� 2��ʃ�-��ǻjk+�AHx#�>u12��2N���~���۷i�g.���m�aM���{�v�]�X>�������S��=���z��}��P��P�w�Y{q���A&^'�n#�}�������#��{�������M���;�N��e��|���o�o�;�ۏ�o?w�:q��o���o�XS�ߓv�Ǒ�?}��u
~��1cs�k{,¾oN�^��{ӻw�8�SР�	7���F�N>��r� x���Z���޽&�	>�O��'|����0�z����z>���_7^s��t�Ӿ��LFx}�c�7C���W��H�������M;��o������&�����t�]��P|N�q�&�@QC��O�
�I�/v�;q8��s����ny���ݦ~v�9�#�11�M����z�k��5'��}�j�ݧ�|N����}q��;M�	������q4��O\t�y�Ӿ~�����N���G;I�g/Tz�&9���;w���?����'�詏L|fپ��8�̥��m8�]��%�O�O~~��8�i�}����ǈq���y���}O]�������]�G�o�M�	�w����ě�����7�ޡǰ�v������q���G��E����]_�*��>�WJW�gÏ����|�7���C�5�s�:w�z�!����'���~��[�whq���y�o�I�BO���u�7�q8��O,v��'x�'O��zM��8c���1S�U�zTzf��`l�X���ɏ�U�uoS�}v�>��á��N�����<B����w���ۤ�;��o����;�bw����N:wI����~q�v�Hqw��� (����;��X9��e{��5�=���g�,�~�ST���LRz`8�ym�,w_P�0���n~��&�������]��;��|ǉ�z���ݧ�7�O󷟻��aM��|��"e}�������@��yٓw�����ز�w'�Tt=T��|.�,��q���������;\��n;�q���}N��O�>b���q0�{�p�7o�P㏧��^A&_S�߸|@�';_���;t��'_��װ�1���P����V�Uʠ�M[3s�f&.9"9��ܤ�Ji�?f�E0$�=k�N�W�C���_T�ն��1N���W����3κ�%pz�A�m��u�Wo�fQ2|`�1I�Ѹ���oEKh�n�7���l�e�#�x���M�����'V��^7q�'��||v�8�<{`��;Hu�����N%q��&�8�C�¹�1;���'���aw�������!�k�q\!&��w�a�݉^���{%�%x"�}
�|f"�=~u��Rq�]u�8��ɽzM�y�t�W�o��|���0�}O���v��o��8;qӻq��:M�-����9���wǈvr=C����;��}��e>F*c�ġ�9���%O���1S�G�*�����>�����һ(����ޏ�|}pU��;��ߟSq�ۉϯ|1;�������<C�aT�����F�C�������w��z�'��w��^�>�>��vwo��#�@Fρ!���S}w�]?�ݧ>�'ӝ��ۺ��������n�;I�~s���]�@����7�`�v�O~p��z���Nw��8�]����O�~C���οq�?Ԥ�*:�_㿮��?!�
��>�*������$��x��X��N��9տ����'�����8uo���y���A۾;H?w�=��Ӵ�|�S��Ǯ%w�=�M�z�C��3��e���'�/���i���g���x����'
w��!�ݻ�x�|>X⸐�=nYL>F�u�?��@�'|?�p��i��7�N>�9�&�ۿ;��o�I��������Q�y'T��x��ۋϲ������$�v�t������4����=��\
o]�����hu������qߓ�����'q�ݜ�L*좜(�?!��X���1ۼ|M��o?wô�3��}�k5�W�]������;�k9����!�©�������P�o����]���q�}��hI�����ۤ�B~���v���M���������t�ڭ�'I�Q�n�;Hu����?z~�L�}�֨�՘\
���e�i��M��8������f''�O�߾�o�awI��~C�@��8t��4�q��>��F:��/�v{�6��;����v�ۉ�N��Ӻv�N�1�L�T��!d�*��i��x-��G߿~�q;��owQ�����t��yΓ~O�����S}O��?}��F��bw�>��o�z�����y���t��O�=�+��N;=�C����D�BH���d!cF��쩪�we��z���f��J���y+h��:�<kڱ����������y%9�&�t�����nՎ�)j�u=k�]�{�ݡ$U6�Ve�K�lr�>��TM5,Bz��Щ: ��c�0=�,
9��Z��I�H�:}*���g-�N�s�on{���`�<+�}���
�+����n! u��{x��:wn����m�v;z����9�t��/m�s��n+�M����~��oP��I���7��w��awn<N8��s�����'������_V�ޢ<	'�$�0 ����w�N��7��t�]�>u�7�8�^���G��n��}�ͺ�<v⻧|?��v��I���|��vD{�4�����$�@���������Y*��}�U�>�!�����O�Vߟ^��N�����9w�C���y�8��\�N�?�s�8z��v�]�������~C�q�~��t���#���BH�<�Dx����}��徼-7i���z:~��D9�?x���f��v�o��z:v���=�I�Bp7�����;w�i^�8\.��~�I�N'~C��+�M�'O��(x#�"�����@��Ͻ������ǵG�Z���|��1��~��鈯���}�?�����o�v�|�����t��ۈO?{�ۉĞ�������c�L+�n���v��$݇�����t奄rP<Hv��u��I�B��]?߿q��>��#���e��}d� H���1��ߐ��>o~w��7�8�������t�\z�q���x�i�]��uС�!���tc�>���=�c��0���{�c!�T���n��|��ߟ���5}�����ڢ����S��3?t�(FP>$��]�㾻I�w:�~;v�W�K��8�����>o��7n�ڭ�?��׉�SN����Ѽ{r�]�}� �@3�#;��4��>�4��p�ݾ�����RKOty����S���C���}q�t��8��q]&��>�s��a�	�����{��>�w����C�s�!ۧk�q����z�����u�7�q�;I�Ϝ7����g�0E^�*����Λ�:颶t���I�'�㏩����ڸ�������|G��F}yr�H��}���%�c�[��]j�R1%�O����ۮ7ɧ�n#ٓX���-���
�%����-�йQq'�����j��^�F,s�fKYu������ ��]t��W�&8䝤m�on����9pW�`.�k<�hL�'�b��
�Q��	[P�r�\Y���rA��Q-���s0���*+�^��<�}.T��r�[j���E���ډ�|(�t�o��%#�B�C�ِ�v�o���א�jW�?-`ݠa4��$㤸
���H�~;���{g(̸9f`���/����T3��ب^�p'�F�	F�������`�}�����(�Рe�b�b�����;8W<Hqu<|��h�Jy��.]ڔ�sIT�oN4x46�0-��w`jxE�vd��6�엝J{_b����<�t�\ל6�@z�48���*؇�r�f?F��)ߗ@iE�toVzy�ӧ��;=ڵo5�V��6����8���X��p�m�qg��x�{�r���E[����O��@��H��n�иMِ��v�g�!�WJ�Y�D�c�����&*Ԫl���o�m��hu��i�>ϳ�����L{��y��g�)  ����G�cl�f��Nw�Ջ��aĹ�n������s{��|.9f�$������8��k��)��3ǶrV��ߖ1�W
���n�
�s���lM�������"ǆ����{U�'��]C�QQ�e�C�S���F����3��u�ي��z� ��+U�'zp��k>(R�m��b^&_��=~yw	�i���	���nц5{(�^Bz+���kV��e�V�:��}�(ҩ;9BiŊD��#�Y%�oN����ν�A(�#���{�oJ��+d�Q���/#�m��Э�w�W�Tٮ���a�2�' _�9��k;na�k����E_mДE=O8��&3寔�hIU����>��7�� &'I:��B��֒���32⪯i���c�.^�����ђ��ۦ�x�'���֯b~��%n��Cstv�z�X�D꩒�a�P,>P�}᲼�Vd��
�(��U9i�]�s3���iL���S�&���˳t�eULtF�,��ȗ2��S��׏>�|�ծ�+�yK��������k�
a���n�=�H�T\�'n~?s�jv\��*�1��9�v�E(cS	�/@0x�\��=$�l�CuhyqO>���NR�;&�o8�H���5�.S1)�{99+�A��:�"<_����� ��<&P#|z�/�t��+
��<ܭ���j;�r�S6r���;�;3�ϼh���#��®�������k��]���͕;Ϛz���zȿ�
v��2a����VL�*ɡ�T˹�h�G�]��-��'ǘ˺�� ӈ"��m�sTeOC��e�OM�(U�_X�>ֱ�榵+IU���t���B���)���2�K+�����p�_�[��	+�Vr�$�ve>h!nJ�ͼX���K|M��O��f	��$�ܒʻ��?�t:P��}�Q�c>N�˜O�����>Ij�ik�	�z��9U��̤���Y�(ׯ/xK�Tbp(���BI�؈��'DV�.Z�&���ţ 5��f���l{E1�+�F z�W���~��'�M�]�{�U�7��=��f%=Ux�A׌+��.�q>b�v����\:̺��\Y׵�[�0���\Zs�82(&%���������P>D�F�X⦀*Nr���l�=���~O�yN��\;|һ �)R�u42#�9ߦ�>t���j�;f�th_0����R�.��7�8�-*5�����-T���͹�U� ��������q0�F�s����uXܭq�u����UӷU�X:f�KT�;�Y¡�\|U�t��Ȏ���gɰ�����I锞�.�j���h���^������]J��<�%o��3�9�|#n�M�*�jY�����}�e��V�R�&z~�upϲ7���H~�Ϥ���X���=p����j�X�FS�z��*)Z�JQ���Hc��p\���X����f���yfM���v�����Xemhͮ���Kj"K��ِ���}�],��r�e�;e,OKu�t��*������]�F���S�շ�B��m��!�i�V�:H���4�|�3º	۝��ZMY�ZŇR[i�v%3���AP��ʹZyD2�Q����>�ݽ�b5k���5�خ�W"�7�e��U3�ޢ�g6��U��!L4#�8��x���E �(C��ө���N\:�(�"b����^�5��g�����2/1#���]8)1��'�uM��K��ڂ��	t�D%wL�_v�p>��-=X��(Z�k	��0�s����G�pQ�*e�a�W�s�H���)���s���0��_C��u!֮'J��-�N��F��4�9���k*\�i�R±��'�����)9U���W�\M���W��DaԮ�gmh�<c��{��YN¹0/l��$����::a�;�w����&\���K�[y7��MA���|�X��+l��R6�i�\���]"�l4:
�鸎ܸR��&����>V2��6���^	QҔ��h]�Mg,=���%��F9�r� �!0��,�C�	ݖWq\�G��`Yy�.�&��f˴�-D�3*Ξ� ԯpŧy�a|������w뒲�R��rvʎ�`��_��b��o�+o�ҫ`�5v���!�"wfɲS5�Ok
��E�v+�J�V�}����f�k����H(�,��i�Ӳ��D��(7��5�|�U�b�Ją@C�?tvC��^�����|�� /ϝxT�5~9�)���8_[(&����Vv^�W�E��иU��*�/�{Ov�����><�|��/>7��|����������������^D����>�W�*8��ؼ/W��:�e%RS<��s�{�Mg.���$=9ܳ�z߅l�7��_^�h\��RV�y��=���:�#/!��K�׳�
��5#��y���zp�����Grѱ��9�9 �H1�JJ��}Zn[9�+�Jx�2��׳9��Ü]P����rV���a��>S��T�������&"gr���������X_�ǜ������r��(�e��8��O�h7w*h��ݜ_M�ݖ>���������7Y�!|�vب�\�t���ɐڿ�\�3��Ojޛ�w�u�f%#��/O��`�wh +~���ߞ�;���\�WY0�ԫ�,K7Rk�n��r���vv���| �]{���t@
�^��q߾8�Av/{2��j抵Rc̖2pA�u�eˍ�r�їB�^Μ��jݘ;���%j%gq�
������{ݜ*!f�����3y��ۋ�Wv	SpN'+�hR�l���t��e�َ��n$����v�{@�f�wR\�a��,P	�fI��ʾ30	��S��Ko��$�_ ���g���ϒ�ttd5.�����d�
�gƐ)��F�0*�W�\��	{���ڻ�Co��Q�F$�>�m]M�������/^�M� ��3ѕ��L��{��H�P�p9�V�n�����>{�=A_�4��ԓı�ʇ8}w5���hM͜6��e��}�3Z�N��r�X��Hu)42s�jU���G��}����i����
���My�1�1u����i�U�?O[Vpq7xWޡvk�7^�	��ܜ 97Q���Y7I�[�M�l:W�i�N@��'���W+��ًZ�V�7��g�7:��O��0��;/RrYa �Q�3P���*�6�_k�-WL9\��Hq>�.�^��p���S�k��8KX�;�Qn#�fXϞTCBy�ʙa��,3�s�%�1��:LgVP��h��Ic��<�{��sd^ ߨ��wNRۺ��N�Y�ۑ�2�Иl}�Mu���x5-��[�"/�t������|+��z׌��k��쨹��O��)�s{V#�eJ0��Y�O�|���+%f)���6�\�:>����d+1��E��"`�ۢz��U	�GMOz��XnU��H�
��ucܢ�ϰD]Wc�n]�
:f��"�s�W\�.w��x�>2��B��o�*sKp��uʙ��Nn�	frj�>dԳ��Q�|�J��-�o�\j��D݊R��h��m�7�9U� ۶z�ܥ��h�OI���c]�urn^������JЪ��5Pu͖��ۜ�G���S��Я�c��!t�e�<� ̋z��m��]2��-��p�c/����4��gtb�ү vdaJ}q��-�&)ـ�l��Dkv��_��k̵�S�5bǲ��+��zJ�=ǂ����
\D��-��Gˣd���;Sڲ��zA��C|��]�R ��y���o6��k������]l���)�*����
�M�|�������'J�J͙Zւ�
$*vW��Ι��^A�룺(D��:�hQ��u��R�d�2�B�ʠF��]���IXZ�0�������(��V�]�u +kRa��"�����u�9�UbF��ؔ�D�e���M���>��Z:����L�;[	�1,�
�u���Yzt�a�1�e�����FFe��M&Xjn�r�5*�4^���ڛ������e�J-�2�U���!z��6�v�2ԇjla\�;�e��fqM%R�t�[�`^��Z;�E��r��lS[Q�oaZ���s�	Hs�x��}������ҙ�2��Ͳ�<rt��֥��v�H���{�Q�	�j�dij��L�`a,�v�:�v��Zx���VL��x�q��T�t�#W�,�ҝ��%إj뷵�O�n3/��:�v��e���3���a���K����K3�10(���W�bhV��t��lgE�Wr����U�c�]I;��>�n��f�
��(�[���Zc�s��'vN��}���iy{\��
� u'p�xTO���KՅI�K*m*���]�*в�]9���E�Ή��z#J��چ�^N
�\ݤnE4Fb������^"�'Id�Ҩr�Z�kD�L��8'?�(ƥ������)��Xl��9�Ou�6���ռ��A�Iwc(�6G�9�,�_K��Z�y�)�U�N�[qƻv�u�����z��u\2�H*5�Me�,��g8(ݛ�bS\U�&;$��Ů�q=�(�" �xc�l��xNq�%<�.ﱮG�9Nڡ�N�XZ�����S�����K��D����G���g{y�����D��Vg'#kT|%��"��c��*[��չ1H�ⵋ���44m�/9;4�����:�g��ɢ��QJ��n.�WV���%
qZ�u����]S���Ģ�#E��9��r�È8s�h��|X����x��	|+�!_ln�o�ᔧ_Z�����7��3X9������.*f��YT�N\^�r��W��W<�ԣ�*���(���<�]�#��4���s���J�šf]4���"M�Tyk*ʊ��:��U2���j�ʊ�VS�yg�����3,"�ˢ�1�,(��T��Y(i9[�#Qs�L��е������p$�x��K	2��BpJW(�+�dm*��(Ȍ�Q�(�&J�ǉ��
�E6�H\�%K�s���Ir!�8�2�\)ĄEA��ʑˈ�"��H2���<Nba9s�,��&x��V(�;���W-��$9�D�1R�&��r4�*,S�Np��:����$s0�,�R�"�"�H�*
2)L�,9h��qU�tIL��0�T�WX�ɜ�:�ЕdHfJV�Ȫ��&DGS1 ЬEP���p��9gMI9�j���-N]9b�d�E�$X�+VP���y�t��.gJSb���c��/���X�4�EN�rot5�5��N��Ill��O�̅'WԔ|��3��z����_����d����pQ3<�后��C��X�<Iۢ�T�R��;#����/.�����>l�sk�I�zp��#}oN�B9���ё�ի���Х2�xL��=p  n�hz�jȷ޿R�\>�gsȬ�o �����;2@�b ���N�#�� p�C���mz�McΕ�]8��AR�]�&8��D_�w�uR�Dw*��*}�L�HX��J��'�µ*��}�xIq�Pv����Ot!I���@�(۰���Rì`=�{3=m�����g5&LJ��=�U;1(8P���ujLhR�B!h0��/�p�x(-dFIEҤ+����[:��jS�b;Z���Od0��|��h��=�|�>@��+֏���.�8_w�K�[7{�-KTb�{̈́i���3�\O�P�]���?2����\+�C�ܜ�j�L��t�Eވ�S��-��߅vy���@p��Vz4*� 6�d�0w\+��s!�iܮ��Q#���.�Ll�к�݇�|�;���j����~4C��a��=X����m�m��,���
�3���U�{��ɉn��Bq�[�U5Z��]H��l.9�*] �e�"4`f[�q�/X�Cz����Kw0:7(>`��
�h�W��Aj��}+�rc5v)���6�r*�3�&V�]S�ٮ�s	�����9N�{�="8EŦ��L�-g%�B���&�،��VZ���ܾ��E�%�]������&���׍��|ǹ�.b�*�F���T�龬��oA�
P��dU���P�7
��S����<|���pu���~'<Q�3R��8R9XU��l/{K�>�Q���2�Q��UQZ�L����^߆�P",�'OC�mc2�z��W�/VW���;Y�>�R;8!,Xu%�c݋I7n��#c:��/a4�׬w�G2))���G��u,�y
�d�)�h�lG�V��L�5QIgq�w,�I�4�R�p9�"!��@ۉ7���!ϼ��u'AN�c���N[�B�󅣹����,�H�R&l	`�u��j����S�$/
܌9Oz{����꠹�"�g��K/���o{���7�o��yJ-|�����f�M��:�9N#�(�+�馊u�/�LK;��:�"������5kd�ԫ|c:K�BC��T-�J�h���n��p�X2<U��k�j�(�B� n�2���D�o0� �f������p B�i�vi5��o�HϜJgGu,���P�C������ȏh��Pݕ*�3�/�\� JW�n���[9�\`/-���[�\���s���k�Wo�kO��Ӯա�}{�����;U&J믮Q�uωί@�N���+���R��1껥d�
1;<m����zr=�.S=�fynKj��}:�˛N��������#��,�W�� :���Fn�Um6���ܤah"*p���5��3�'��@s�������Ĺ�^��և,�^e{7=彴1���-}��*7H���La�Y�D*�|�we��fE�y�(�x�r�"��d����kG*�tM�5GO��[��s=��3��Ø.2j���Ti�D����u�U���v���C+�>��f&�������+�Bd��\�~���˲��&��O�߼r�?��:���O�j]�z�dm�-�W���;���贓���̒�I̟�B`M���u�^��[�x^ҏ�[��s踓��;�]j��(Zz�F��v���#(k%��]�$;|7��V�lC�Ju�_IϤ`_>"�S[�Zq�<X҉2 �Jf�yZ��9na�.�\Kb�+|	u>
��|�Ŵ���/9_������E�����ګ�H�B�)����k�{�
����˾����b����^Sf\�.l�w+)U��.ޚm��8�
kuSY[nd������U�/G:׈A�Ѱ���".G���ڐK�]ǌ�q�1s�|���������;[9�u��@�V�p�ZK�E���I���|��[w������#Y���S��֥�O�vm�n�>�R�8?Jm�"�D��c�Ġ�tk���n)�'�^ȜM���j���]���J{�*P�� ��(��.��ʃ/�6�*�0&�c������W\W8��=6�X�Cv���9(��ٗӢ W
���qtq@���7ΞV��Mm��p�T�?�(�obϜ�4.2}��Ⱦ����~ `�q�r\�������vOA�;O�ޕ��w�:��龁rX��!'��m\T�	�`�n�K�{�*�!����wj��Il� z�W�&m`�4A�#�?J��<�G��G,܅�<�#a���!Ԏ٣�.;�5ǵ���h�W�-��g��&]NP�QԇJ��;��Z{U�E�QM�Q��;�}͕Y�WD�pUژZ���*$���P�H�+���̡��Գ�KV:��8x�as*^���E�����G'��:ќ���7j�z�=0���+�	��vǖF^�	��j����g�W�P���*���� ])]ݺ�{�h���Wt���H�ՊiE���1atp�7�z�]�����c.L��И��{:f�N�����p�cr(ozU����n*I*��9Wv��-�8�=5�yS��]�W;�(�7dh��߀�����1m�s��7,�oHf���|u��:���2}��Vf��έ�(8Ú�&�{Ԑ�{:T�ݻ�\�ѱ�%���+�'d�rE���C�7\;�(=M��Q����m��lޢǪr$Ңps	`��������u1z���8;r%̰�鰹�Vlix�c�T�R�o��z+�:`!v��W �����v�f�W������垥���Wzק���ef+�P3$u�k!��X��70d� �Jf�A.�p�BC!v\S�kn�ɳe�K9�ܹ��om�������+W"q/��{Q\ G��5(���}�]ՙ˶��#'P�d_�u�qE��3���9�]�I���I:��&#u�!卡5?A��B�����xcc�E	�"�YN���66������*Ɂp.K7FjᲔ&�zH
��Lz�
�H���H�OA�H�q���Ü������fi]��vKy�ξb��$�48��{҆��}p�4)\#!\2!b[j�f���]�կxG���F�N���r<�����#<f��!4O\��-l���f�9VT�[igٓT!ڸ�18�D��o �(��1q6�i�d�P��eN��������yP��BU9X5�c���%+*K�
���e�:Q�Z��7�7����ky��:�U��@V}�$�o�4��Y`���](S܊�_#�<��h�3ϭ*Т��H���h�_l�J��Kg��������.����Lnv�~O��+��wJq�s��%CVo���G��D��9�*��N�1��ʘ6r�i��
vx����Y������Ƹ����T�Xf�)Ll���q�ȗΫ!;����\V���e���uF�%��3�/�9r2�!^�C�~U����N�ʬS�z��`lMΡ��k>2���Pa�}>�Vۇ�M�{��
�և��7)/a/��88Z�j�s���p�sQa���(�����R�f�q�VΘ8k��;�aB�IT��vZzf )��\E���jy�J�jfqe�Y{��`��e�B�"}���P1���s�@ܨz�P$Y���̽�����m�7{y<#����Q�jե��\T�Ǻ(﯃jEt�#z}֓VpBX������OTiΚ��{g�pr���E1�X|>���]Kٮ�W�lOg���r,�2B�k�:�;���:��)@�ݰʗH+߶�kU뜟vZ�HF���rT-�F*H�t�A.�3y��' 8����`�_t�]{J7��x�+-�V7e�+4�+|��D�)3�E.N��c�l
k_s.,�\�R�v^��!�*[����� �nyoj�ݴI���U��W�{~�pf�}^�|yC��S���n��۪�[�����`t��zW��R�Q|�\�K��a]��]t���pw��>��A:)�y=�nN�{.#�J��e4���?<��o����ME�\�WyHr����s����c5e.8ݗ���=�[�9.���'���?r�z��t�����:��y���iNY�?`�����9��Av.�.9,�S����ҶؗNd��ə	�"ũX(���oV����};���E��YP�#{!L\"��6�,d�.n�3���ɇc�!�`�;�y:1n��ׇ�������6SA��Tt���\S�#~E�˵[=��yw<�Ztc�܌�XK�Tf6`��S�v�r09���i1���~UP�9��� �kA���t4�[�LU\U��+TBJ�gRHi��N�ˈ�@,�֦n3��3-��I�8�M}�V�z����r8\��4o
�l��yu�%����:����]*���/�V_��FS�B�_�F"/�*�}(xC��y�}t�M�y䁻�8�mk�+F��|���Ү��/Տ8����f[�:;≢0��E�u�Y�M���皪T{5�F��Ч,�9O�K�V_p�� �B��ڴ�T�;܄���9=s7��5�a�c.a��  =�3��wv̰̻��&�������^'���t.Y�~{�\.P�}�3����m^1��q�Bn�2��Tv�z�Pg��؉/2~������s�s�+/���]N�e �9q��Vj;�=�ܗ�xf���T���QR��,�ZC�ç�+���g�����4�j��_��jJ�Dt�ajN���4sԗ ���M��xN�Gƽ���p]K��򞩖Ѡ�Z�i�mqJ1���H�_�˙�3D�,V}.��)��JC�&���7+3e&W��\�.��Ȁ�쯝B�7t4� 7s��B��$<K}�8\�w>��Wj;�q\丢^}�D��Sڝ����
��{8��Q;�]��td(���B���cj�_��\�-��������Mb���7(j�f�bʙ��:��pY�[)�;�HL�{�S��-�]cS`ޥ�9���q�	\:�n�>�~ `�q�.o�J��U0�d3���nF0�b���;>БVP7 Dm}"3�g�ڸ��[I�c!7s%́���	y�!��h�b�R���6�ƦD�<�o'qcyX�+s�
!�pܱ�X��U��{|`�T��aY���<qq�\�ƀ�O���w|�?���`�sՋf"'dY#=zh�߅��5 �����W�n%�V	��/P�0N��sN��h�N��������z�^�|��*��B���_	z��8�|я}g�� iM��{v
�l�R�4��m>��tY�}��U�ag�F�YVpP���x�Ga�Ԩ�kĆ
����T�Uş��vS���Dk���3KU�L�����ieY�S���ꡟ{,6+�O�/z���� C���cq����HO�]�f{]C��1�V�vX��j�{���ؼ�Z��n�r<96�����w�xv�>q֮�l���Y{S�*���b~��o�q^��(�#�;i,]���iWa���+��e���Оu2�X`8*������Fc�8���5�R�mǪ�{��ڰY@z� �r����[hS�����|�>Ǭ�y�k۷�<�M*z%މ	V���[7�(��ӂ��Oȃ����\c{��ۤ2T\������B抵��HGn�d��L+S��PҚ�g~�DT��!���@��!5*�515�b�y�n_��+��S��p�qd뚐Ü�����|�+�9�T�ll�-j����_.�
�~�l�\F���|�5��Y��Cض�k]��w��]Y	ax���shyx�ð� z��ֺ��3�=E[h�tzf��Y9��K� �������\3�#+����a|_�d�"�юJ�
r-;H�׶w���pK�]�9�6~������o���coC�"gxvy��Φn(÷�g -�GtBvgI�4^o�z���i^b�n��f����N�H�ʘJ��l�����E�����i�a����j�f���mt�ۯZ���+f��X�D�H�-�NC�Vn�5=�"�$.<3qx��u�ڏ�!E#�V��d�l����
�>I0��}(k���:�C4)\#!\t%���\u��G�Se�-��W�����&�BiHũdz�>FǴQ��{J�|���X,��i9��W�<�3����A̺�N��u���hk��j�`Y��?鱬�K[��,�^��)�3�����ӛ͈�$m�Q�:�j9]��"-Kz�mu���Ʈ��:�g�g00��ʽƆ�.��6p�&3��Îv$K�U������?nt��6di���s�Ύ\k:�9���B]*�Ge�Lڠ�� ������9�We��Ρ�]��S�'9��3*Y���̀�M�_�p�8K	}�������0�wV^~�ЀK�,:xf�<n�z��j����T��ZU��'�1�
����uVv���YRM�7`3N� xIx]Dz"g#Yw� �Z�8s��cmb�馲��7U_=t����Ը��1�C�V\jA��һ�(:�s��PA��v�H�>�ں܌b���D%�\����w8��Xq��Z(i�Р�eL]���䮉��|^B�qP�dVt!�%Ů���6�����6�̛Q��UƵخ̡�C��"���2���2�t�.�\�	��>G���6%��1zs(VA}pve�O5��{��̘Jʎ@3z�Ѽ��HހԵ�]@�N��h�\��u؍e-��/+K[R;ҖegooV��+�II ��#�w�6�ai���Vv�= (�%+�u�/�)sR7(L��`�g˥ct]+�����0pkQ"�=�+-��v(މ�3^�=�k�vg&ڷ0Yx�ᤫ��~T�����Ҧ��f��:)���H�o8�;�XvIV�<3�(�V�d��w�]��q,�=ϸb����5b�#�������]���b�SQ���'�WVǷ��RP �:0���vjkD�.���;�xn�
�ށs�B���ǹ��s��i�hp�/(r�k�&�M|^�a��(��B��j7ii&cV�"Ցު�t�����=g�wCx�$����8������Ńgrn�F���KZ��u�Z��=ne�BU�[A,���L�����۫�Q���,�˱W)>Z0t�����:b�ۛ9l��z�$�sN�nY�:l	e'�)�(�"�k�+����Q]�'Q��a�+�
�d荬3�貟f����X�Tv���P�� �]ж�0�;�U��Y�_N2�8m�m̩\��;�W�WIf_;���HN&��M�f]��R'
7C��ë������'d��j�kx�y>�z������-�]n���v��R;�j�Py��:���W�+xc�0R]��T�gҺ��ل�:m� !���,%�9�S���d�.���푭��*����R����Mŕ�/�YF���V��6�RP�Lun��vu�芎	��<�y��>��Q���v�w�x���ou���K��rY�$�rC�!w^�E�)J��!�즫i���`wYS{���(�
Ek	�+��gs�c$e�)*���jO��	�]c��W�k�q�K�K{{������."��5���L�N<�5N�8���wЕ�:1O���ь�U���+k��v�T+�/�֍q4�*}G,Y~4��Y�J

��O��
_*�s����Ȭs��3�f����X�Ν���������u���v�e�]�A1n,�mHX�V�����gv���b(f�Y��M�K�U��TjfVn�3��*<���e�:(��W���-:�z�GbЍ��AR��g�ê�u�F��Faoo�c�j|(��e.b!GBhYf�B��LT�͙��R*��S*А�T"�$�S:WI:�0�L��*�+�%�RiĒ����Y%D'#�gJ*���(����eT�H�QVf�TQ����$�U���e	�j�"�Z&�L�[N�d����js��jJ�Z��#L����f��%Qr���3H)�+RT��T1!V(��"LH�(�Ȣ��*b�J�Q�U�9�īL.!�M�%d�N��a�W,͑aTj����6���h��N�W(��%N�f(�T�K)0���V�� fW9�E�����4�9&���9I�d���9H��NU%FHUl��-4)-9�U+QaTRA�JJ� �u�F$PM:s2	3M,2*��M��T!b������x�������h��!mas��k6,�u.w��<$���!`����j�r��\H�|��0���/4$���UU_W�
O�s�Ȉ�m��a���w����+�{]�0k�����.:��
��æ9֚���i�EI���f�*S:lyfY߾�C��h
�_��QZ�N��!��Q�+�<�ɋ�΅g��t|�x���cޘ/��*���k�>�I�>/�< ���p�ў@��1���k�ݸyh���E1�X|>���b;5���͉�W(���㾙���6���@��3+�⁚
��t�Aד�Rj�r��*Z��컥��II�{q��H�*�����F�k̅K���Wx���fN�'�����\�wZ��ԮJϡH9�<W]L��Yy���u��$�W&�C�_!N\=�he�`�1�9����=�#b���������ݲ�RBu-��Z�8�+��Β򐊺�t�U��Q9΢F�t�6ӆ�^��S�V�g5�.a���V�{�̗�d�N�LT��R�Z0��R��=J��O	�9�Q���.{�u�yc�����/��]n=�ef*���,_��}vD]KV�[��,�f�_63{(t�M	%[xzVɗr���ظ05az���\�'�� �aT�5��{������E�HT�{�6)
���̨rm	
3���oV��W)s=�P���v�J�a�nl�l|ZSS��� ����{}�w1%?�ؠ*s+#��#bSA��Tt�Gmd�a���̤G���V���{�"�Qߪ�׮���g\�>��������}���%�W���Ll��j��*wi�ھ�t�y7j�%J�Zԅ@Co�þV��U������C�
s{�㍬�74�����)��u�v�w�c�?,�uv���﮽\/����l�9��ӝĸ89lɗ==3��a��������G�a��`^[XX�}P϶��, �HC!�t�x��n�WR�����Q��~Zo���s!��ֺ�O��곓�w�\�w��$�I(]�V� \1�n ��;�,�Z�>r�#^Cb2�s�Pp��6�hû¶�\E����������5`婇9�ع�䱑�԰ȩGMd	E����v2�
'��B��Y"���@�TO �j�0����o<o��hu�f:�'$ۭi�)J:+ʗ��$;��x~��B�77@��d��>d]���o�d\`fxM[0����t0/-k�U��:tl�N0��q���״_�?dAd�Bd��Z�<�½�3�j-��Ɔ`(�3
ǀP�MG��:xŕ�})Upf��5�3�`Jȹ��5
��� G7�2��#I.2-�;�皊ۀ�\�J�3tg%��*7�� յ{�����w,�ݥ=>�mdC��:~N�����i���y�s���J���Iq�p�f�������a��Ry�F����թ���\�-�ٕj�B�p;�vi�*��m��=�������)�oa,���4.9*�@�ṅ�.����������
�W斧�3Գ�U]�4<�G�Vn���#H��I�|ڨ�+i0,�dIl{��zH�����.ښM�´���S�6�S��?�=���}�����Z9�	��F�b��m��M�6j�l��j����l,�^v��Cxh/�U�*����+�;��O�ٝ���3d�OpF]N�c$�Bv��.��}_q����%&�J��.�t=b��АN��2^Y��C�6T�]nfOk�s��1�*��|k�P�9��U=Uj�s汌�κ�׽���ivEXo�[Q�¨�s2q�ʓb���}E��+��_Jf%f��|����W�@;��T��2�OL��@v�W�N�\�(�k�]7�}���;p��݌��(f��l����W-�Kmž��p�n{LJ�J�ډ�L��*��t�1���W�fҹ���dU��˖ۑ�� I΃�}\F�+3�^Wh�)�����SL�Cp���I>̇+1)]����9e��	��)C�0�~�����d�����(#w�p,�6�38�@���t������
��?����G_�6�VԬ���N����f�`q�I����O�t�>Dep
�걽���T�껮ޝ��/�,=M���]�Fӌ'�����e�Md3�+���G�:Cs��PW77�`��<�ȃ����R�5�~2s����db�9n�`0�z�`����:9����f�g�E4���S.�b������Y�A�m�ܝ� g�D�:�4�����!���ᄙ��i
�p�S=? �􎐈z���h���v���a����}�:(gv�gO�O�ڪ�̸�ɀ���T�j��([�ƷU���,���
8�M��]�W��X�V���.)LS�ja=~v��>I�U�}Z��|��:�oj�+W)t���<�5#M*	~��Y�S��`u�eR�� _V/B�<N����5k�Տ�+���Q����եa��H^�S��ϐ��lp�����Z`�_F�v��:P��3fDZ=�S�\^�c	����rN�C� ��)J��
����j	�v����g����$��fm�^��� �k�Y2�w��x 7]�u`�;�LJ��%ttd��Z%u;X�j"�+im-ځm����\��u�]GC�N]��h���� ��t�#��Z'���ӗW�j�.]/|��h�yFa��8�'o)�UN`��ܱe�0l�Q搯W�k��N����{RJ8��HWp2@qSڪ�(�[�Wpmʚ���jw�Cˊ�|$X;8�{�:�o�<���DG�p6hf|+);�j�<�-F�9�<M�˒��LA�c3���{o��="Vq��ċ��0�Շ�F��K��	}��8.��=���r��K12��@��v�8�M\����E#^[`���H��#G�a����<)�^t���Ɗ�=����ngX�D���H.I�����P�L8N�����4�lK�^��Y���'���:�7���Ĥ�V�S��;V�&��7�;��멕�<��ȫ���+��mZ��ejΤ�;���>��t��e�7qL+�ҕ<]K��ep�hN�o�m�p�Σ�Mk7�����^@�#�q�
�k���pf��MdVU9$`UOeE�m�Q�q�:�e�!��O�u�+�;t���H~�bxK�PR`�e���;t�W�.���V�Afv���}�=m|ffc����i�an}1顽YKc���]K'ϰW��J�T���H��6i�7�(P��tv��0���O�f��Q��Z��7ܛ�]�v*�v��b�d"����Z��^sp��b�\��F��:��'�W�}�}O���(��$?�8�>Ub��Q��⃭H�-}ƭ`�o���kָ
T|�N{U*�5�-���j��z{���8�N�m`b�HN�������L{�p[��A�n�|Ov\W	'_sT�:�*U�H�ȎV��sYR�%���数˧2^����B���]ݜ��QREv�۞]�m���h��H7貽{�ꮺ=<�ζ�,dN�2�ӧ3��-��d媕�
�9�V��^�����,�W��yS���Ǆ�9I�B6w�S�#Qw2�W��צ���?H��7�y��(����A��P�u�hu�Uo>�z��#�q��işVn�gh��is�n�)~L�U^���Q��4+�V�K��뛄���ǀ�9�W�m�MD�)`z��:�ן:�毎w������®�#+�*��u��ӮS�y��J���_"W2g"'e������gz|'���_G�a�yma�P�>��4a䉎'6R�._d��ơ�Tv;�Kd���#C`M�*-���G��˞�Q��wΨ;�i��_K�F��'Zw��@SU��c�s��d�j-<>6���س�۱��dsE5�c����t�}`7�9�x� ��N���E�3���)nQ����}�)W�3̱���}'�ss��f��R��e�#ur-�U��Q���.&�i J��(_�x��oqX������FS !t
)_�u��QR�Գ!i����V�k�lS�!��t����FWC=Y(5�=�U��R�`bҒ����ϲcH� m��Cb���K]�7�n3|�-*��%��R�VB�ԇ���|����&��:��;�
f,V�
H}���ΙŴ7��	��8V�pN����e�v�P]Y>���F@0�-����E�6Ҙ:r�g�΍h��n0��][�:c����ϲ%�R���3����c�"%�j�܂�,>�?gu���_4������A����#�@����(7hϥ�J��:�dV?��d�����j5�E����>�6���u;r�ҿ����q�T:�ݙb]�������*�f����C�w��f?{g�-�~>�܋U��߂"1ryo�^�5��i����ۯ�6ж��wWva��7s�y�g�) 3��a���Y�u��gZ8����@*�\,ܪ�ҳp�i.�Ȯ݂�,�#Y�����k�e����H�	�e���:��R`j䥍\v�v���J�e�U�d�����}=LC�.��ĮNW�n,�s^{�8��[*�լˣ�K�����$���f���؆�3���*�%DGRɎtd�ъ;5����\�q}o�#��(g;s��\@�Y3�s���9��q�azL�T�v���}��G��,;Rr�'��S���d�­���jao���eY���8�� ��ϼCŶ;�%f�y�˦Vui�\#]]�be�H�=�I�u�8��+����;\�B���{N^�^��[�w�$��9 k�2�^~�,Q�{�m�^WgS4��K����������F!y���Ҩ�ߧ��G-��<�������*�� s�����,34�����۝�;z����Z�Y��:Ъb�ؓ�Y@;� �r�|r���K�?Mf-X%ɼ��s���o�e\�:e����tz��E�6B�B5��zKqb��~0a�:�:���p8p��ՑS���x������s(u���gEc\M�� إ3�M�c��,��z��j황V�Y�U{#����Є�������;P��i\�xU(�� �Z���V�ΰ���E�(��@�$Kaj��ɍL�VC��g -�Gw�ْ18�B�'հֺ���/ے��H�x���bʑi�.�x�q?X���T:0�[ؓ�S0=։���\�25��"v�Ӝ�ƺ�z<��s;��gb�$3)H�.���7w!�,a��b�
�R��|��6�,`Q��x��w�3��Y�n�Q���Ŗ��d�ΐi[,b;�%rz.Tު��X�yǗ��ݮ�]����AAεC�=�y�1���}�}C9-j]�t���|����k$&6�j�uO��[�����ݍK�ea�k;S� ��N��=��b�˝��2%w�^*�^���>���
���q��[��վu���ð��")4|�n�הSHa$?�V%g�ᆄ{wzSS����6$��})��,5}�#V=����*Dc�<�U={�;,�}Y����;���\&�YʨՂj5K�y4� ��t�SGV��E8�s�l��__m�©��s�G`뇔�\��,��������aSݮ��Z��뿅c9K�n'}�Z�2�P�mVT��B�f�n)��׾i���ݰ�����������_8w�����$�Z*����^ޞ�m�s��x6�ݰ�'�}��iCO����Ȯl��j(�f�-�|��g��;�Z�l,ʱ��P�-�a��w��{#.�;764ƪ.477�܄�8�ȁ}G���jN��XMJ׾72�9�7c`�i���0��W�v��y�:)Zc��D���x"̫�\��n�w~
��nc��˳U{�R->�EWi);��jl�Foa�.�}r}5W��f%��j*$�ڀnX+���,r|E�K��w�:��5-�>ZgVz���c�ﾪ���Vgz7'x���#��Ѧn�T���܍p�녩��_<�S�":wx�'o5M�V�M��L쨿��i,]a�S|/���.���>�Ν�����]u-'�0�\Dܺ���|�I�JH��� �%*Dm�|�iq\s���K���S�(�4�&�e.�����C����H����y9��ѱk�;������S�
�3%�M%s�f�"\b/ �٩�(���$��G\Z�l�ȗ�VC�
��*z�(-�	܆��T�Q/�7����f�6�����A�f������v&�s�h�Ue�*��Ck�-�r�N�}��ݱ֗Vo.�E�������q�vuN6	��;�/RY���M{�2���}��H�%��D��ˎ�=��f5-&�/(5�=����
�S�^ÎUG,z��ӈ��o	�g�����޼*��0��($���<��M�
�؎��6�xV8����dW��42�n�^�.�Mf�+U�n��&-p��nQ�T��%]ˮZzM�1T����`o�0��V��r�FRq52��S����6�Lټ@-��n����`��K��ٛk&�K�WR\�Q-Ӽ�Aޔ��&t�+h�_UlŊsx�����Z���;E�ٶ+��t�lzN���/*پ2q�������Ѻ�ͩ; v����w+5��#�hˣXPyW���z#����|GɆ�$���Mi�WJb-q���GyK*�Ѻ&t�a� [����u�(>ͬ(�ND�5��4_pw;�R���\�
�'qM��ɷ1���֖���Y�iҜ]W�1�W�����Xj��m������ÏC��:E���4�̆��5��1֚��ODvR�9�b��������N�F��*�#ݥ�<ZW�*
ͽT�wxՇI��s56ж+stT{�˩s��7/�ebZ/�ε7`�l��n�&�N�M\��`���/C6��왽{]|团�9Ԝ<�[-s4���;J0�]��Ću}5WEJ�5n<�깨<��㌩h
kR�]ѧF�* .��+L\دV�<mwm,������o&�i6��į�]�L��Wl �j���Ez�?ڏ��Eq<�1("��k�ţ������m?Q[�/������M��q@��&�I�?(��$	�n��|���!�U*uv��;$��������jʋ������; 5j��໢����޺M%���h��"����^�E���x݇�$�̇o���z��\� �k�u�I�[��\��I�O�oRꃜ�*m�mut�Fa���ibJ�:�*L�\ͤo\7 Eh�W�k͗m��-Q��][�i1RY�r������`�c���8Jwz�3�D��3��t�y3L����X�R�f��w�S��Th���f���.�(нuD���
cFw+��o�E�L
�.�;ԑ��˺����"����*�I��a��Ⱥ�\��_3]A@[��Qt���'y*^up����>���&1r����@թ��&�"��fm���1_+��ƽi�6�
��<�6'pÕ���6�)��K��p4�֚oX��*�C��$�H��gpyl��r"i�71j��������.��t�y�"��.j強��4��% ��<"˶��FU����+:��3p��/7\k�ogv�+yoD���&P	�ǵ&�k,�jx��s��J��B�5�S���C�&��c�Q��c�#����.�wE +�G�Q�[8`2���N�k���9�X���Q#��fm&���TE�W
��X�1\\�?��v�)p��(9���*=�ِ�ܑ�G�ڱ�lD!����,8��|����W�\n��G��[�[S�bb��ʾ�C� A�+�T*jq ȺҔR�1CY��8[VDT&��D���HVČ@��2"�	6�Q�ej
��*�!���EH1MS8bsVJ*I�T��R�e�$�(�E3�B2�DUYY���(�)���RQ�i��`T�mR+.�&G""�P��i!tE�%e"�̉Yfr:�sL�3��Ί)!*�j�IBR�աȨ��"�!%#�	��U
�"Z�%2��-J�R�YK9+Yi25)UNe!�e�(�EZa��.E��,��+JL"���՜I(��R�Q���ZH�)4����TRJ�p�����dˉӑQi��Dl���KbE�.��(bE����#T�!*&gPS�KV�b��"am(�I"Q�t8iBW%1IJ���)$:d!\4J�JRIh(̉U@�]�e Q���W�Ʒ����0�3)q2����E�<Ҽ�$o&l�m5�3�pw'�s�u,=�eE��$/�}��}�Fl�M枸����CtZf���6����3~	��������V�l�	�8y�vA�)�1[��T[�^/�����y~�m��,���Ryz��{����f>�n��늌,����'�����*�b�����"�wػҳ/ZU�z��2�'�j���p�D���[퇍�v_h�&`�5z.��I��n5�7}3��j��U�]:Xr��ԭt����x�v��Ik>���w���e�W@�77&���
���'��0����ѫj�&r��M"B;w���K��ӌ���jͼ���'��m!$x�c�3WB�w[q\�����Ķs�+Z;�z���#sri|L���u`Eu��ԧCwHSӽ���8�jd�i(�y˶�nr�t�%C2�vg�3k��l"���%H�I��Er�GQAM,�l��x���E��Pk��l��ؑX﫨��#Y���S�5�������gS�d�|I�ҥ�}K��8�ĞY��hZ�fE5�a�s���]a�e'�|Ӓ�dT��x��.�P�����ٲ����(ry�,Cb��fu��5�c�"�������B��*G����>�l=�ͱ�R�QȞ��i���OY�"��f\�%	�f�|�Ij>pm�[�Ad��bx�ܭȖmq~Y��c�yy���̷9�R��)�Tj�f��sW[�NS���#~�~E���~�	��w;E����i+ʌ�v�v|۾�\��|�z%W�����;_�＆���������{�M���\gsJ�u�ϊ����Z~�i��*y_[o\;��������5�Y7nZw�vD����ی�UO�:y�mz��L�l�Na�5˴�fs%[�eٽ�ȚNTk�/�5�Kw��"�+P�z�Z�m+B�
�E��h�������a3T��ezmZ�C�z���Ѳ�{�����l�|Z[^��Cn�����<k��>=� ��8w�j)�%%��J\���q�XblχF�ʋyr�#I��/��<����Mn�J�!7��lؾ�:�Uт^���B�̎"�	pe�~�M�*��]�>��9'aV(���.i��Ҡ��b�Sf.�t�+:�E�Y}8�>��K���Mvm-*+΢i�H�hӛ�o9��A�6��&b�+��o{?����"4�cVSio���n�z~�nk���i�|-���4\��g���O�SƧx4��H���Dx{�!#��\�z�fr�#1˦���t%&ȳW�Q���uJ}�4:K]7����L��L,gO��Of�;�.sv.��,z����k=Q��Ȁ�M�E���a=%�H�)�����w��bG8���w_����-�����ō�H'��4][�����I�z&���>Ԧ_ͳ.�f@T��*z�Aw����\�i������+v0ARwT�a�״�3ǹ0�6n�NE�㚸�v&���Ȟ�d(�:�F�~.y^�Y=���?m(�}p��I�,p��	��*�`����xa7�ZFf�Jf7W
;��|����ǑS9�:9�vU�{����uzk��}h��ۃ-���p���V+Ț];����l��T���V�VWA�N�ό�w�∉h�����[|��ڏ�����v�9R��p$�p�9��I��Y�Q+;�¿U�n*=�2b�[�z��V�"ɲr;wW�v���@�f�n<J�]z�oS�K��tn��l��9�g���*�0�4�{���>��%an�sz;�����j ��>��w�>�b��&���Ӫ�����Iji�-�黑�4�U�J=���n�|.����c��@\9�gU��*q4T��n����(�9��ZP��Gd�4&�dt�v|u>A���s7]V��Y��ܘ��Bm�vZ߁YMhf��L�!��Ia�9�jy�L��9���,���
լ�os\7��Zi���{�##���H\j�D��3+`(,���Ib��{�w8��κV^�]l�=�y��<Lrx���d�����*�OY�	&�E=��Ȼ���ݪƊz��T"t^]���y��-�T:B��K�j��K��8&�w��lS��*�U��?Q]��S}Pm,���<�jmB��p3��y*L�U�����0�;�ҧ�ZG����G\ZȖ̼��S��HED=�mU4O�;�	�	��n�8+�'\#��M��K���	���v𶛦HS��^^�޺V�v�@=�ܾa�m'V�҈H�]��.ձdm,����7�;�_s�Ѽ�8]X}��h��j���K���n�6�א �f| �$���Qw��G��+��m�H��D����Ymug$�9��5]'/%�琱�s��HeS���2�9<%��]}#��NTe>��/i}���z�UF�t�v��ai�8�W=�ϭrLv��e�x&�#Q8�6��o�":�g���x��sհ�ۜE��o�S�U�^�G"`�^�Vt1�_/��t.��=r���uUe5ފ�o�7��.(��w�fl�1tt#KO*r�[f��f�����y��2��ֵ�5�us����E�ȇz�"�����������Vu^t4eb\-�K=p�o�i�Y:�,d+-˦�Wn��r챪wY���l�����䭌��[�=�
G��ʓmx���Y�[�xنqڳ{;*o)��6�����|�ݙ��ĕ�#���J�����b,"�[���{�Q[�5�r�g��)�6�˵�P���d��G�oC8�i�)m�UҒv�&5���Ұ�N���hu9��q���9�"�.C-Z8�fR��ۦ:2;rm�{�B�R�L�R�ޣ,+�t���v�ts:��.mhp�G/�V�w-wΔ�Y����Qvfl���p���e1"�3C�6�AJ��X��x{�[k:�z/nY�Wܷ�s��\-��W�Ҋ��~fT\I,];sUP~MfR8t�4��Z����Cgsⵣ�G8޸nr�#q7&�ě�4n�jB�A|��uL�l"�N������y˶!>�nr�t�<���]XO9���h��U��*����k���r�DqM%-�y/��.��)�'[�i��UyHz!����s�as�Im$S���֑ur�,6+֯wk.m��t��Й �r�U��otD�q~Y�ZUpE!�|Ӭ>�������]As�j7OS�)��.�9��*M}8���-$_���������^+�&��&{�ϙ�]	;�\��|��+U��,��:^���Z4�m�l����K��=����m��*�ϗ2ֳc���$��d�m8f�r^�8���Օ}����߯"�|���/>UO���X��<鵀s�Q�oi�9�q�)ya�����e��m�����2�\�����
�-�)t>�������=���Z�s61��sP�xM"�U�Tuv�//]@#�3���9�:5��s�;ʺ�*p%s�8m�/��ouww��W�}T?zw_��#�Z�F�-�T"���:�i9Y:�,e�4f��=����t�Y�4�s�Q��iK�*G�U�j����h;�CڧI���o�V��l<l�;=�g`�S=����\=�[$uy�IOP�v�pnn1�[��]'���n-L�����1�9���m�|/N�.��;�����M�Ds��5���4� [W�ܔ���p�v�⅝��U������ϗXw�7������Q�7����Jfy�_7�+Q�7<��\��K�����C��At��Z�SW!�H�NM���]Bs��8�D�	lK�����C��6�55�Ӝu�Vݹ�E�Kݛ��*2�����Ճ��6��#�i=����L��y8�U���$u��up�2��ޔ~�Ī���w�l��]�җz��y���>4v�?)���<Q%�8Z�𾕁�W�;L�����E(���u{t-3X��-����M�F�8���b�Y�D�R��ל-^�����[�����=j�u�v��8��[���N�(H����S'T#��>�>Ù�x^�N�U��k�!���w�f��$�_�6�B�s�y�ۿ{t�]�ūήW'���۾�^R�]�֟Vo>���Y�N��k�V��܋�u����ڹl{5zqb�[��s�7L��`�,�z�����S9�:7�SK�C[��qD�P��Dؼ�;Q9=M����ֹ�UV�<�괱'D��&Uv�]"�5co�٧�^�s�a�O�X��Ϧ���V�J���+g5�ub+b�	�9);�ؚ$�v<\�hYR8�ڶ���W<��Xog�s�h�,��n47%�|��V{�aα�����Q�t����Z��T�H�rۺ5}n��ke�1��M���υ�wʒP*���|��gA�L�D��ti��
�V�a�}��L�f�CE�j�!��8ϫ%���6ng����>��7��|���at{�~����h�Pe�$���u@)��a�sv�d�{���+^h1+ڙI��qD�30Δ�t4�&���ib�8smN�����b�ᇐ�q$�n�QS��S�µ����P��f'�9�m >��q��S=�����犯�yo�p�������nWQ�DrL���荾�mj�ꨭ8`ﱙ��RWv���	Rz�	&�O��,,ݓszL}ϒ}�������K�{S�����HQi|M@s)t��zF+���z���˱����p&�}/9-��7NWʐ�bߍ^I/��ҏ�}�S�2K�ie���d����>�G\ZȖ̼�x�dC�
���{8*��ü�����MDr���g�mud"�4�l�\$���n9������a��c�՚�ݱ4�LI�yYK��":���ZQz�!�u�]�A��ͱl��UW�\<��j���F���G�j1��~S԰��3��w^�&��ܩ�.58�ã��u��V�����|j�/=����n_��/���ȥF�)N5y�^*��~N�L���E�ˈ�;�����(�*����ĕ�֞��J�}4��DQ��?*-�;�һ�2}��7�7�ٷ��ޡi.lţ�*I9ܧ��Bu����sw	��R�v�sc�ݮ��B��X�T�q¾^sʻs����R�z���[E��%��s�GP��n^���X�+C5������V)��5���=vh}}�FL$Xm���UU	S0�sh"g�v��ٽ�Ϧ�5�:�,b����"��k\�Ǔ��I��+
N�*��<
��$��#�S�޵	dO;Y�N�7�|�i�Ϊt�BҚ�S|�<�����P;�5O��ߪ�H�2U�m���(���$jcG4�U�{��
f���.�@_2��i��{�)���je���:��{����]x����ɯ����]���=i�:�.�gq9����?@l����o[s�����W}��u>�ۧ^��#�|G��r�s�g�#q�����^r��d������r8�Z�G�@`��=2_VGZ/��9j#x��D�e�:�py\t�fk�Zwv�Wp&U���]lQr�萕�H�\�ҝ�9�� �O6���
�~v�1��)ķ��@T����Bpn���/��g������O�/Tɖ�g��Ց��u��b�ۣ.pʏ���e�$�Ю�R��r��݂�6%u��k������6�m�u�pe��Q���5��7��MmKI�[3fo)Ҍ��V�|ܝe�J��+{Eȫm^ֹӈ&+�$�;lMó �ն��宱��-����ڣ]B�Į��.�1V+Dv��ʒ�I���1 �ˆE�S5�v��P�ݸ��ܾ��x>zW|Wfd���M�Q��Ke �QV�Q��_=V.�
VV�����N '֠�څ��2��䢰ҩ��:�;4cVӻ�-ګ���M��\�ڊWe�P4Ė��Jَ�+Nf�r�
��A�|]-���$c��^�e�-�(@�U��ܒ�Y�K��չ-�w�jT'��X���K��͝�#��H��Y|;�3~�[t�ԛ���wkz�jLA[��*a�J�Zn
]u���Ig+���nN��]B�-���e5Y,\�ru3tkq��ʾi�v����&�l⬨��{�}�v�C��Jk'�幕���G�7R�PNy��X��Yf�
��T2����	ej���}I�Uy����i���4�l��Nȧ,n�B�G�z8Q�K�ZdW��B�Jϻ��t��x ����dY�@��)Vܹ2ڜ\�_�V8�hb��b��,�Y�n溛V��,1�KȤ��:!ڲ+y�����t����fZ�:���m�:�����,���>o-u��V�SY�t�]�x�X�+F�k��1!������Oi����ΈӬ��R��f�'n�1����SYȎ�@.E��I�M�u$�:U1`�n
��iawؑ�'^ø��g1VgTE���"����EW�:XĨȅd�$�䭦��h9
c'��Fλ�����r�*�[=xs�b�5�Yɘ򻉬�θ�\�<a�D�\	�=w&��^v�\��X��5������5u��W{s����=���+S�g��f�� �����uظ���_h�y�(�+�݂O`��̤�P�h9�|o���6Z	6{ �\�[�n��Kfڇga�I;p�̢���Y�EU鷏�!6�G]E1JV�D�1i�z%\Um� ���wݔ���vMl�(L��Mĺ��j�Ҙ&�e��eqܢ��e]����S�bۺX#��9�
�������۵��,�����m;*�ܷX���6�{�,�n��Nt7X�Z?
A�:���0���[��4��-�;�r��s=M��\��
�^�	#N�W
t�MpY'c�%�l,q0�L��tyԨ���&�r}]*N�M�����Y�7A΢F㎂�EQȹ�*��a_ �Д��^rմmM��*TW�F5�uva,aK��9H�^ݒcR��v���lA,
�t`v����]u`鎹f]k(�&���K1X����kL����&��;b��߻��X�|��N��Iʅ�0%c��W@���={XY�V4	�d�ϝ|�e�He���3(B��FI�*,$ʓR:l���U3��*B�(���U�3iXfFeE�"��6uiZ�D�洖K!$��H��6X�J%J'*��]i���.Ud!Z��:����:dI���$i!�3BԤ�F�ȍbh-"�#Q*C�	�"�;DĂ�IS�\�H��UKK��ZGe�.G(�Vt�.�Z�AEb�U����������F�E�J�W:j��qK
��!A�KR�J�!��
�MK�-�\��+J��8�A3����r��:HdY�ċ9Tf���DB*R�6�L�Z�Dh'S,(�J�'.fb��օ$&��0��I]�,ʚ�
��p�jT5J�
	���a��p�gj"���-J�B0��u�P�[Ë[J�r]�j)'�[*u�Z�Ax�c�6��罥IhN	�*xB�x����/6;�Q0T�M٨�wֿG��.Gi;n�Tgw�Kj����q�����h�58��^$�Ԓ/���P�E�m��ҍ�I֘��}C�!�V��[��z⡳*���N�=��%�b��F{#y;��ǟL��Z�f�m��6��n�i�b�{�/zwe���b��ӇTe�MU>c~L��b��si�VwVc�3�.A�l���5��I���Ya�I3�Y���S�ޓ��Ǜ~e�U�t�-Ũ2z�ƨMϾ��G�
2�3�{���^�Y�%�QF3':Q�����;=��n(˵o�j(}�R��롽�6����ݴ�WW¨�/5��e�zE�D�o��`N��I�#�
�|/sez��:󮧐s�V��7���nF�]p�}�-��b��M�+�)Z�-��z��I,_�B��)����q�7���_�=��)�� ���,)�cz�T�,��1�haR�4
'��%�����Ӯ��y�m/XʉiTx��=Pn�[��l&�<�����1V�S�tE��B�/����Һ}]$¨N��������ۙ��V.�Twz|���]J��:h��U���{�w� �Z#�Vm�?��(UȬ�Ӻ��3���zG���
�z��=�ݫw3J����b��H���r]7��q�x�wlE\J+���[\���<�y��̖���{I\OH�LӼ6��[74S�u��J&uɪ��w�E��?Oy��x���
�T�I{��\,Ÿ�6{��ӛ�E�i3[E�W\ra�Cf�$�6�S��΄�VtQ�"�d:�=�#���mnWciw���6�y�;6wV�ä�ܷr0nK3�2�8��E_s�{�7&1���Ot�/����yg�&�R{E:E�²O�RK7Q�Y�[��N�����#������Ft	�E�Ŭ���s[�j� �2����O'��O[g��_�1���N�LotR��m�ce��)�;�Q���|�Wd&�7��<\�o�bu*���-Ng�f��#\������CǪ6F_�W|�
.5aʕ�q|+�pC��7^>�`��b�x�$i5��B�gn��q�_7w�9����34��f�t-��h�q*
q,���-fs�g:<5Ш���'4�$'V.Q�*�ar���w�*w�W�X�\�����wR0���-͔[��m�+=���Q��W-Q��E�鏶_�I3����w>��u}nϧ�������M����CY�W[��sF��s�&7}��	Wk>� ��O ��R���\7�ryҁVCMwN�HJ�oթŠ�l��뷟	����Ib�7®�M�մP���a,�R��Yi醻\-�ӊ!RW7&���>�=f�	%�~�H�x�zws��V)]U�u'%c<�f�nr�!QI��4������.�>�&1�;��.H���Q'ig��ؗ�6��*B��.;@�n�/�^�"]�\��"J��/��Ye��.�*��t��fĀ푺%�E{�����ny{7�]Y�)�sA�f��N];=K�WE�Z���EVI�ư|]�����]��r��\�?G�����Yi���*~��ԋj�|�_����^-������gK�ͭ�[����/��5$��_�q%����@��Fa�`b9�F$���U�l=x����f�enhm8�����|�w��V��Oec���s�K]m����t>,Y���IM�T�L���sϖ]s�x�o>�ث��G�j1�����ܥ�mV�s���FW^��M��\��ϟ!�#x�������o�S�R�d���6򸎵��=���uaU={�tZf����.��)�kB$%ʳ-�z
k$n��ne�Ms���+q��nT;Զ�x��R��]j)�����Ay4��-�a��*%q��"iCY��,�U����EF5Z�v���ɿγ��X�;�_�����G.�UoZ��y�Ⱦ��9F��3\�e�+�܉��ޥ���}���`�S=�����t�PQRM\��swDsX�W���.q����n��C�� _��4T�J��W��eܛ��1�w���� �<�z�8Zc]�Ҋ���dnS�<��*�NmjZ��_�,6k�Xo����֎�8޿z�{:1��j�p���{}��r%�vM���[�N��fN��wTT�������� �\�%�����zDhsw/���c�������i��`vޮ�A/��f�[�2��I���r�֊��2X�W��K#�b:��(Q3r���m�nY!��V|��:G����Z݄8�F�L�����a>���Q瘞��\��i�2V�0�OX�#�}��NzE��s5*%ڍk]v�e͹��k!RK���tЋ�ّf�G=G�����	�qI=����w*m�j[�y!�T�HN���eV�k4�W��ڼ9��F�d���E�mU��Zn9�ˮx$�;;K8rʆv�^����L����'/#ٲx���^ǵ^X��A�sJ�-�˞g���͸�����Q��h�o&���̵�͎ǫ*�������oA��;�ݸ1�̒�1!X�&�N�Q[���Q:i�hu�V��իJ;]Aa�[���1����ݸ*%�kk�i9T�]+��j�0���o�zy7	���W%�x�O�$y�����\;VY��Tٞ���C39��T��w�
5a��4�ռ�l�0r���Z��J�����{�R��2(�ۻiAE�Jp�J�g6���+��n�-��rA�T�C�g��w35��yV's��B(yi�d�����Qi�ڊVˤQ�[� ��=�q"T��=��[���}�<l�;=���_Fv�3��-�5םuc�ܭ�V�!��ӵ��e7d;�S���ۆq�m��v�`�=`�{W�L,̧=Pq�v�G�q�0"p���T��µuq���nk�֚}SI	�
fx���w:;P\j�EO6f]|�%������|,$� �h�Y��t)�p͢�E	W]=J^����m�O��Q��V��k�a�}�V� U�o�+��O9���&UZ��N��/s�eZ麗m�T�+f��-�u'k6r�*2�p燇\6��y���/vnȯ��fK��l�T(��Xr�?>}���ѓ=UŴ�	�U�aYE�l�Q/��d ����N؜���6��xȔ�_�>��3k��6��Ҍ;���I�1��,�\7u��o��$om��w�V�L���K��Y����w�s�{+Q�HÆlT���Kk�T�ÃQ��� ��lJ����v	{1��c6m�wSWҰެ�E���L�of�5�쪑���[��I�p�f��r!���n��L�RemY��U4	��`Q�Ŵ�]�b�e�=��h/�Ԑ��-{[쵞��^��+Nf����:�M��s������Oh�2��]q;��=�H��z���g�0R�h���Ғ���p��ܝL{���j��=u|.���]�*{`]��Ky�ě��I�����yH���-dCV6��m!��s�pTO�@�*�ɨyV�mf�H=9�ֵ�i��:��.-ˬZ�D��v4���`L=t�� J4��>2�.X��f�&�%ɍ��Qnq�}�
�v|��p�oH'Z<9n�xU�K���s��W֡,��v�477�(oq6�wY	�뺬kR��f�^Z!�.�P��G{~{�a�7���J�������Ȭ�q����>����S&�
K*/�F����i]�����w˲��p;��j�\.����蛒~gB��Q��*�ب�ONj9Μa�Y��M�-�ec=��o[s���$���[|��§\T㛁�6���م��聍Yj�\�9�	�kr�eZ�W��.n%��z��R�s�\s|�*�Xԕ������h�̅��]B)��W�^�m�����o&`}y�4�Īudor�N1���O&�x�젨I�u%��I��%�y7���8ޢN@M(eI*��g��>�r�@�N�p�����E�2��9�W�}��w��:��Kf\;R�Ut��1V�V_K�Y2��{*�Cw�_e.u��шE;���l��eFl	��\K�-�N����g�ʔ�h�x��-g�"5~�.H�,��λVl�oS�ל����������z^S���؍_k(�'��,�����X�MC^W���3��Y�^��î{cU��f�}��]c	ջRu<�՝d���샸�t�jW��ªz���~�^d.<�A@�w`�V�Ն�?N[������⣸�_nu/��ҹ��-N�\Q������<m�	m��v`-Nf��,�[]�4�������9����7�>����	�3����i�e��5j$|p�2�߭x����/��L��E:W�I�wsW����v��Σ)���\�.�ؔ �e�K1�
�ab���G��K1����{�.�$;2�u%r�����xz홧�ǉ��e���ֹ:b�G$�����J�R��W�^�C
�'j�Kp�����]�<L�����{ҙ�ĕ��N�"6����$Ie�9}���#\5��8�>���Mɢ�z��A.0UR�4�ꤸY�,��>��)��$�9�]��u�+���"�R���&��-mQH��� ��<.86�V����c\��o_��\��W^mAoPqj���6�&������.���)�Z�8K%�.y����ì�Y�ͫ�Η�S�1�D��[V�P~XQ��_G]]×�{1b��s9_>�\�[v�K�x��ȨV�~ʫV*�E��fE�[�x���j.�v�$seфٗ��k�YR����bz��*-��4�ڰ��,�f��J�m�����xں���Zn9�ˮx&��7�f,؎j�����l��ݘ��v����[�J7�'Z�®>�}
;z��rB*�la�
h�� �[�얙�$�Q�0�0(�}]C���֭�`)@�mn����M��K�\Yd]�x�0�@2�񨔟aμ����u�2��]w�+obi�'6(VH�����=���1�nN��԰(XPk�5�]-L��,?Uo\ʽl��+�M#:cy;���-|���\V�����>�����Y!9m��m�X��ên2�U��Ψ��&�E�F=I�7Х�R՛�\��&�������&��u��]����)�S�QFn�3�v[�w��D�Aά�v��hMʰ�]�h?�1��l���3Y��T�6c�}<�\F���
-��l�;=̵����=��%�t��n�]���$VD��O��q����ㆷ!6�;O�_EC��)����n�Z]�F�S&���D��:���9�\+WWɾ�b��
[+w �p@nMi�P��}@�7����_$�.8$���o���f�l�ޗyN�Exn*wwo-��\r��z^��͛y>�����?N�M�k��7�u���v��'(>�O%�<���C�P�*�r %���r�*���T��f��C�cޤ�B�ێ�U�PUΨ����:�\u�ً�K��im�e���S�JS�-\.�:롇�f���r�ٴRA�ȕ�s�\� �9��uԳ�Ru 9r�@gmq�c̼\��'hl9w��`,7|��p@
ͬ{�sR-g[�a�t�6�j7[1+�%F�U4��BTL�.�8D%g��&��g��f�[X�s�"f�$P`4��jv�,oܯ��y�[:'�np���O���>�"�a�6+�	o�al��Fw�RnM�6�CXA�� �Dd�E`V[5oEУ7�V_ػqQ�������՞�ُ�V��\�]�]� +���7��:uݘ��ڻ�Qؚ[Ȏ�z��Hu�I�5�|.���e	�w�'@c�����DkK=Ś�5��u�h�hR�v�=�U����@;�=�0��mc�!&7>;������L�	�to��aڱ�/c�`����l�D�F���3#ԝ�
�v��C�Bŋab�ݎ>�n��+Wj��Ҵ�¾�7R�����[�u�B��U���H�]�c^���K�Р4..���"��e<�]�q�H��{j���$c�[���r �7�w�[�j�h��(X2�i�|8��f��ވ�:Sy�U��.�5uԱ�p��*�&	��P�
yĮ��u+��Xp�ݩ�o2�N^>�P���E���G�_0δV[�"��c�]��m:�I!`z�%\�ʴkz2�u�.�q�㴘�N�l
H�4�wk3�y�X �7aru݇��7��ڼ]����(�]�=�[�&��P�����*U��Z�w{�թ�#H�"�]�6�R��`�:l��5u�h�7s0���fWj"�s�[y��	ç+��Z����8���E;������N�t����z&؝,`u�E���1�;B�)�����E���0Ӊ��v*M��W)��[/����j�g`z�N70Њ�-���{6XX��v��7tB����Dc�ڏ1�o���Մ�M���>�7)t)�"1YYI��ܐo	�j�+U��ZGF�}�7kܮwP�}hM���M8�ZؤF=�kD��b�C=�6�����}ڷ�zغ)h���ngaG���ABf�����.�|3m:5L�s��dU�������v�h���p{RL��K��ɺ�!݅gK��Pt�O;2�O��i�Ӂ<��m�r����]K�!�S��v���5���/h�7�����5$WcM[$[{0 ph��@�g)Է�QѼ3D��k�$��1S���5mofh	c�5ɬ�sn�,��x�E�bֳsهIrq��뛥�r�W�Օ�u�*Ē��H�7k\�9N��U�5is��;,1�A��3��]�9��c��w�JS�[EK��c����_V^A��|�xx��X��Ƭ��&��x/��3z�a�����3��]��_]
�
�ZJ�G0��#S!#	3""�f�A��t�aS(���*��9�����J6r�UL��
-V��F�$�UQ�B�Hl�E��\��T�Y�E)�r*��®U�dә \*���Y�EEL�
�L��*%\�q�9r���CR쫄D.r���0��HB�W)�DEI��(Ԃ��A(�"T
��@��$�B�W*���j�F	Ӊ�JU�\�����s��"��Q9*�ȃF���r�T\�l�J���R��9f�H*�rJ��&S"���'���*8r*,�T�̹�0#0�*WT�d!����K�J��ZG*#$�sR��.�CfPY$r��"�VIuH�W&\��eW3.�BAD|6tn�9���KD�\�=Tr1OD�J�V���u
�����o�����IW��L}+u�w-�V�s2�h�wڔ�>ƻ��r����c�Ʋ:ঔ;���J7ZD�sI(IJ��Gw}�a��IN��q�^�C�������W	�/>��^|�*@Vc(�wO.��E#SQ;�"w++���[E�Ɇ٪䓑pێs�.T�����+67hK���D��yQ��v�Z}Y��ѼY	;���yiU�[�Ao#x�G+xTu^��<�Ղj5K��]�C�1�Y�����*��s%�*�/{����i����:�W;��uP��.��=�RY�80�V��r���s]�Y�T���2�CV6��|��;����<�U��S�A5���ݐi8���ƨ��ˌT[�w��]��V<�L�����h��m��&7k�;r�O��_dӆ���oCs[��m�+=ݴw��Fr:�*<����h�=�D�]A���K"y���(o8d�E\�dwa����ڱ�|��K�0]�:���Ӯ@"�cK"uR��`���Y���=���L�e^��)L�J՛M_�E�7ݍ��:�gO�V�iΥ���`T]8ų��͖��f���&�Ȗs=s�jہgl��S爘�Mű��*�w���~e5��>�Y�Ϭ8iy�$ɓ��<��T�K���*��e��G1A֚}�/�T����Q@�9G�d��(6�^��(����Tǈq]�\��p�k��#���IEI��5XFu�w�f���}�i�7x)p�'!��ȊL���+��z����D����7ʁ�K	%�X����|[�!��\I�	��K�kb^��S���S`I�:/�'%��^��6mX�j��/������E��[2޼�VGN(������tC��q��Ԅ=�H.�'���:��K�>E;�h2D8Ga�U,�F���̜�맻�^Kq�!`�Nį��*�{�Qvf^=�&���]ٍ�]e�ʌ����Q�
�n9���k���.��i�qG!���7���G�%ϋ����d����C�CʮX2�U���H׷g�G$���$kN�ȆT��'HQ�X�c��0�k�V��ͧA��EK��:n��C�~�g_��6�G�HW;oX�J���c.��	�Ed*s�5�]h��\q%����tk}:w�pǒ�5��yO���Wŏ��\�B�#ImZ!��5����ӱX� �3�ɯ���UO^�tZߙ�Ŧ���HxV�`>�	69۰C���q��V^�M:yA��^*-�;���D7P��{��{�V��� �T��j�YW��"iCY�0���Q��<{w�Ss���~�"��il՟j���/�ЛV��>8iR�6��e��/����{[K���=�n1�a�g~Z
�kG2�[��a̬b�{zW���QT��z�k9C�5;Y��5�[��9U�<���ܻ]}��4��������9}��fXw�7b�'���p���8�$[!��	Z�
�7�����ϫ~]@��%������>�ȸ�µ���\��$���u�ȝ�g��7���������2�O}���t�����2bQ8�/�7J:�]�^w]u�q�nq�0�*�a*�� ���E���"ù��y�њ�N��{�/;�C6	Gl�#�R�=����������OF�te&kx�)�,�m����3�3EҜ����NK��k6荎�t*7�|��Pg�m�=�ݢ	m�]���:�u2���^`NiӰ�@nGԁ���+�P&�s�M�
�Ȣ����*Es�_�Yk"��_.�BW="�s��]K�-�������䯚p�t�2�Kq�!d ����Bqǁ�𗝘�b���{i>���O�I�Ͳ��\��٪p�9��7���ĩu���w167.
�4�b��\�?Zر�H��6�y�͓�l��D>�ѯ����Ѡ.7f��Eo;�e罃��N3s�� S��6��F�w�� �d�IB$@K��-�o����yi��D�7Ά/m�Q�9Y�s^�c	��Y�n�n`Hq���s̙1OC�g����k9?�#S����m!dw)�;э�+-�G��S�"�-�Z�ο&9������oan5�7c��f8��un�5�<�l�=�a�g��xk;����Gv�o:��ݙ��D��t멅ѩ�����8krl�����:���ۨǅe��Q�W�$����Y,�@�>���p�,�/�K�����5n���Yފ�^�^��P�=�$�e���Y6Z��-h��gf%���|5���(#��cq
��֋ˆ��o�)ǫ6�`�2J�ڂ_Z��z8z�.`��Öj�n�z^�QLLn����.�[��*G<9�\+W\��ᭁ��Wd�Ă�ky���
&8�� ZW7&�.d��	%��	,]a�����b���t�PGEe��Z;�y���#Mɯ���%,7�#�-��9�_R�Xg�fx��ac�i�M���:B���-�3Գp;��z�{
�e��!K��݆8�ڈ�)����{�mdR��s5��Ht��̹���J�SC;���������Qui�/"^9y��C��X��q�/9�K����R�9���K���L;�y��z�q]免sSW���z�'$�c���	��lK��G��=�όga�o_z��#�X�����1���m���j�5�]N.���E�t�r��x�%���ŊX�KJ������u�`�c���8b'���i-C�y���F���wW���}�=����ԉ ��ψ
c�����in� ��ˬ/���k�����HM�x�ɯj�n����Z�1��}"]��p0��O	*�� �����؍��{V�Q�=6�(�
j�%}
۸��������ח��lr��Ψ��a�5���'q�e�|��e��g{6�>C,����^���>瀵�P�1Y{�5�NN��,�ϕ����q9�N���goQY���ANiE�}���{V����ڼ��N�q�����;o����_�w���]ͨ��s���v��,���tu�K"y���ܪ���70}��:�<�V-�)��+����˵�{*Æ���ȃ��m��op�Tb���^�Ȥ�����p��]i���7�ܒ�OU	B��G�q>Or5�|�j��<��n-g����\@I�v�Zq���6���sj��ͫ�u�2Ocq����r�E�.�9I�a�rV3ڜo[s����j&��&��d�G���3P:D�o�kv�p���K"^s[/vn�c*oj2[-�>���s�*��j�|5f�}� ޲7�-L|x�ɼ�z7��������pgE[���',^���޻}��ԖաH�]��y4��9�g<��&c��K�)��û�7�@��(T�nZ9ǂ��;\�i_4�T/)b���ԠoS�(T/]�RؒwjR��oeP��Z�ȹ�yM�a����Wˍ*���]����K���k��u���x�+�tNxz��N^D����5OT��/*3"J;9V���up��}+�#�&.]��\$n��&�Y�e�8\���\�Μ��\>V�H��4',���"ߚ~��m������:����Ŋ�ٓp9��\ՔfmĬ��<+�g�7������U=z���������Cg����G�z�"u7�b-^O[U7�e�[�m�:�nK�s�s�p�r�����z�t"ʾ�~��W�P�k�����Zڳ������	3�־���T--��V�4e��r�(~G�3��5bH��;n�b�2�r�\�[�����[���g��/���Z��Z����ə��樾�kP��򃿵+Y���p��o��񸛓fK�E�t��f��nQ�n�5'.�f�D	��%Ԭ��j5;�ݹ�^d#zR)�;��]I�V�5��Ƞ�u�(oh�|7p);���;i�⓫;��P�K_}�c�`�������3[�K 8�b���E�]����;��,1�Lp��8��9=��o��B�7Cc�}���p�[�]d+���|j�8����r��/�K_<�l���ұ������e-�����5�R�*df����yC���Ӻ�L�O6h����r�ŝ���Ԟ�[v���{[���b�?]I�j�~X~�c�� �I�f�A-8�UÞwm���/"^)j�U�T���gTl���w���i=�X�)S�'�O��:)t�-Ƶq��PT�T;8�q�ZF��b�܅o+OV}�_V|��E�ϛWV�9��M�<����wp�Q��}�4�KH�{-��R5V�,k�����^G���=�as�G����5]�ξ)��{�mB0.Rv/#L��c1t
{���;��v��`Z�h��R>����8q��ry�q��}u|.��|�e�,,���X�I��>ڗh����`DòAA�: ǔ|.���jho-)�D�,i��:m34v��C5��]�)�N�{���T����V���S,gr��|�y�B���%�1c���R���(μ���5�0]M��]U�ѥ|w�R�J�E�<�k>uO��L��_vGgTc��T��Y��.��fMwXe���Z��\N��,��
�s��vD�ȃ�Q��o�R� �jKU�@|��ن8�X�,q ������K'�+�ܔ[�8��c�z�i��wۚ��@�ҏ*��c�}#��Ӯ�'EG���[��]��2viުY�Om�z訥�8�z���S=P�Q�y�{���
��tqa�0����Q]�L���mEI�.dʋ�%���j"<I�I��E�~���-��ùn|޴w�o36��rj��R�)2`v~
$Ov��)@���?zI����}�m�S�*�J��I&^w���6Gwp�5���ߐ�q����P�/�k"���813x[���<~i�4�Z�rG��2%�O�G\]\&̼�x�¬�cj���GgK=Ȍ��cV]D��ب톣[&��)��0��r��/U�ϛW ���<{Y(�.��̒,.6[���y.��i:/q�0k@=VEݼ���)������-d���/Bo�C�A����#:�E��3�������D����^C��=�R���e.u�iu"�S	�n�*��H�\�V�ݹ7�M��������Y{�o�$g�r�ID*�RK���;�;;m=�;O�{�j��{�s>�����N�=�������p�*���׽db�k�_��P՛�[	C��=��������>��Z��ۊ9�˓�3z���O�>�O��w�v֞��o���8lB5��ز<�W�z���^c�2+�?����+@��~�^�v�$����|j�+��a=�_|-[
����n5yo�g~v�������<���T{ъxfw�Շ�������ߤQ
p�؁n�|�z�+8z�"s�׳�����9�u�ԑ�Θ�WP�ݮ�c�ʇjer_l�:�X��ɋ�����[ؓ�ɇn�P��wD��uqKq̚�'�b����|�v��ʲ��#�Hd``.����V=��GB�xZ����p�jG�#�;2���
;�>��L�2��H�2��_ʜ��⃙_D�U�>�٪�bf@ޭ�˕��B;}�c�����\�s�(�#��U�mVF�U�\���=g5�sA=V��8��+2��j&e���L����'<��K�T��z�pd�5Z��Uٓ7��
�VXG�����l������%3�
�.�;�vm�OncK�&V���.�':3u��<e���WN����B(/5�c���]O6.��`���h�،����f�cf+�:U��ܘԜ���2�b޻�n6Q�}��I40�`��	�.�7r��n����-����g�Qgc��������(P��Ağs�a�i�s��z�p<���V��!u%ji:��j�۬ҡ����`�jʵ1��"�Uv��9�r�2��ɸ1�ʊ����r�'U�"u3�)�K��*�D�K�v��s�i\�e���<w�8�N)c:�ϑ��c�>.���b���'Z�hD
��
��
�p�۲�
h��v�е�G�1u���%o�>��u|��Z�s3�ƲC.�k�:��z��d�Ѹe;J�099�	�g]cm�5��-(���*�%��'��Z��c{z���8^U��#�z�z�dc�)U��p�O�ؾ3���+�ܽ��*��Z�����$����*{|"ӥDj�^�Vx`L{srQr���wDa��SS�6������(�ӀFuܮ��E^$*������e�����x��0,˸�Q,�D�+��>�rtcI��.���1��&��	73CA��[fD๎�OD��u+4�R�w\Hwu ]��XKz��m�:�<z�ԗ�U�٠��#/Zn*�robk"�m0x��b{�I�n�XSk���9);��Ƥ6��'O����uA�5����F9'']eեB��+�ژ:_L��].�[c]�����"��s�V=U+��^�\��r�3Cԥw�=XJCk���[�I�3sى�l�I�62r
�vC���37 =N�i�fD/`����R�ƥ�����ψ�+��2�{,�O�e�.چ�!�mm��ə��z�
4��M��ZTZ9sj3�f�HeJ�u �ը��m���*�mӣ)�3��ɹ%i:��y�����	x�g'&U�2��Y��]ĝ�b��H�X�M&�2���I�M���]K{��bZ<mR�f:Kkq���9Ku�YYӭ��@f+	�)�OA4������f��wi���n��TC���)T�l�ewM��cm��ך��ä
O+�,t��i4����(��%�<��j���m����\��[1R�k�z��"b��B�����6�8����+��L׎fp�"r�4e���w���wbщ�S6���`]'[tf�kUIb'��4���R]mN�ʰH��%��;/n��:|��]���|:*��%�x����*�cgɻ��MVqVn��	K� ��[��7*��u�k�Y�%�T(|>  *�EjiΦ&�%Th��
�&'#�r�&@�3(�'@�EBHp�̩:EU3R���"Q��QP���HH� ��\ՑQIUQʢ�As�V���$��*(���"#D �+"��2J�T(�+��UU�#K�K4B���(�Q�39DU*d�DfUp��j�\��(�9ʭ�"�EG#�a���SQ�EAW����*qAD��"��9ʸs�W.PD�¸UG**5.DUG"(��I���G$��
���eQTG"( �UșD�dY��PʊAETW*��I��B̪8EY��k���(�
�0��P���*&�hUAI�S ���*�&`acJ,K*�3�9�*��UQR�"��h�g$��r�".EPh��B�K�r��e�錠z�*$���2�}[Du�&�ʋ�l�@o�ǫJ��Xb�r��d��7�,K��j��:R`.=�$@�׿����4��]xd_�r(7~�b�|�F�`��V�ϢFHAt��{r�1��>�e.�L�H3=��<E{����YC~��SY^�$#`=�"9���Ͻ끹��#Y�S�0 ����s܅N 8{�&W�Б-��א��X��*C�,{Ny�z�]��$�\�7OsW=a�Н��p��!A�u�M"�zՌYMb�>��ʓ>�o+��i���E槽��V߲}��=,:Q�4��Lڦ��T�Mg�~#H����+��o;�-�RO��8�=�S�*����_�d�]��w���,0}�B�ѭ�p�Q�Y�v��ᢼ��,�xƙ�^�{��޹�X��\���̛��mP�^����S�^ST�>,�������}���M�_�^#>=������g�~���ȣ����(�=��/甥XO�؅!��/Nץg�������çac��N|�N-�N��v�z�׃�}�φM�N��=�Ӝ]��b���B=�֌!�݂��滃�[WÅ��ߑ�3=�W霘�:��w�0Du���[N��r���R�,@�T�㙙�+��'�䉸��9$y2������"
:t�5h˛|Zv_�,�(E7qAϚ97��o��-V������}a�˝����+�K*��u��[�n���ql\���&Y�s����$��٭N�G
�L��v_ v!��Ih��낖�x����,��4[��6T[`ߟO��;
�M,ʊ���>�R��l{/��5�%�?i����S�dPz/�F���9�7��noI�G�v�z��ye(����!����g��xx�.�q�Y�;�e�De��t 1U�ߧ����<6{{�Nq-�zh�n}�W^�[wLsur��z��{�>��z��=�#�Ea	�oXS����
�ª��n�H��t$+�bZ�8�zu���ȋ��&�y�3���doz���a �F����<�ҕ��8��Y�"r���>W�3_HK�S�j�t��O�޳5>���(�}.m�=W��r/�wUo����}�
U���>2֨�A�+䄾�ĲR�|棐]�^Ĳmw�9^K|�j;�r��;�����ru��{ޡ;q��EZ�
�D����4&����ȿgxqޥ��M���F�����Dw��8�����J�P_TqS�E瓁�����o�.�IRvM@�}�⧷{����װ����lkT������ǟ������!�̱N��n�c��V�Z��q�Z����eڷS|�K,yt��ֶ3W[,U��\]eΖ+8_Ea��ٰ����ee�~�mR�1�r�����YA��۩wc},>:X��|�,�����>Jw2蔗,�6`Rl��p�|�v
��%4�t�dƄ�֔�#�A��3?[�2wl�"�~�vȽ��dd5���Ǽ�,F|������I��5�`��B�s_��%�,����@Q��hs�G��k����NCY�.u�aظG(��m{�������0��Z�՚�[>��0��՞��2�k�CϪ���~X�H;�s��c�(��wR�~�o{��3�>���C~����W5�v���UNlu0;�T/�"�s�h��ֺ�3��-+���C*�n;|�Ӯ��}U��p��|�̝�;fo}[CPr4h:��"�g����;G���8�<6׼��'W�z�Ń��ϞW�+����H�5�:E��'�=~�gd��y*��Gz��n&�ϳ�����ΐ>���=~������x/Z����ջ'W��i��:o���v���C0АlW�܊!����8���h�_�N}��[��{�y�]�Í]m�^�o�(�a݋!���E���!s���f|i�]Q�W�n�Sv����>�~:qn�h�Gn�۟r�lv��e�~�>#k=p���O�-(p8�c�.��o��K%���Ѯ��N%���`\�x?d�Z<H|�>/ �Zޓt6���Q�ӍJ��u�o���bf�h�ڰ�������G�M�=��f��f�م�X��ч���b���8U�G.��N��K�d����;9m��-�#,���z+<f�M�	%�Ո~-�������p�^���>��#<�N�;�+"$`Up���Pbg�G"_%�Ń�.Z����#�QAwx\3��Eg�ؐ���l���NxS�UHA��(
^�T���c�G��5IZ��SA�w�QC>��ϓ�6"}���ǫ��;ٟr�^�=x�nl���.���X���T;՟@���M��u�.yc�A�b��#����k=b1���z������sU�V�>��j}�ؓN�� �7��B�D����z����{�V��~ʟJ�������ڪ�����WW�}�q�*�ޯL�;ə�>˩��O�����ܤQg�OxB����F3kԲ�=�g���}��,d>�����~���>�L<����?���0�:訉)L���O�G���_�Y^��p�O���Ϯg֫�*+��.O�P�����[9d��^o.����r������s���s�M@�Q��{G��u~#�9����<ȮϿ^�}�U>���LV����ܿx�}�!�t8vEW�n'����N�W�x9���}3.���G���#�~���bߞ=��n����rI�(Υecq�Jk�7�3�Z�^�89���ʪ|O&�L �w!F�����qmU��4��t]�9��Õx�_��j����M�+**�ܚj�'��NB�'ya,)���LT�5b��,�\����",��P���I���+���K���D)7�w3�^��z�"}�_M_zLxoi�\U�]m3#ݖ�;��:��G��
���U�0FC�Q���㹖�;�SYNu��>]���;�`����؇���l{1O���<�C�"W$�C]��F\/����b]�����]{=M��|�r(���!��p�	���ep�?;����̬���$���t�Q��U�S�7������fs�e�=:�]xe��"�w�z����ީ`�o�	�ul8������9#=̟J\qo���e�
s���FM�,�r
-���W����؈~���q�F2k;;{|��~���(>H�u�@�g�!#�j"j����L�ReE?<r}�9��c�3��gu�_�G���3��ht�+a
{>��o"h�K֬b�hx���)Z�U����>K�n��T���%�G�hlD��Xu�ɗN�e*`�EJ�Ȁv����Xq��́�� ohO8#�<I��a�넇�>b�9�+�ۿH�z�3=��f��@�^'C���?�݋$3������6V\OУ?n�i�ڵ)��`ܦ�Sp66.#��k�� 8Igz$��A��L��Rx�prƹ�P���K뇜G����f�}x7xM����n�s�5��X)�@��]�����%��i��Bp�]��! �ktԕ���� f��eE�.��Et枯9�+~�A��:Î4�/�q��<��S.����2|��z��OG�a�7��.C�	=zVD�l�9h�&���?��z���#��/���n=Y)0�����J�S�w�x��Eh���
���+"z�^}W{�Ӱ�� �>q�ǧ]߻}:Ⱎb�;Ԫp\����Hg� �S�o��B7�JF.J��Xݮ)ӋVlzGj8�f�)n���ｄ�7MX�l�:��#}��~��F�h��낖�@�z,y\<Yلh��<�S��$����}�fg}��O){�7�~���Y������khu������꘽�^X�秃V7��z3�q�X��R��}wDOz�k����~�zH�2�e�z%�1K���/s	n�����sF��˷t�~[wLg��佂=~�ީ�|6;����y5���y0�M���W�ѱ7#���H6)L�H�s��~g.�2��ɬ-���z���ޏw�g"��!z4��tV1'(!jϕ�)�Ԅ�U$�/��3���MO~��T�J5A���A��K@&��x�޼i�;��6ĥ�&���?86b��V{���N�B{o�_nD�B)R̨(��[E҅XИg`�����.LЙ�Q�1)H��������5s\�Ĵz�PQDN+0^-�㕋!{Y���\�]��E)GEe�Ϲu����<�P0w��,�r�f%.�W���n�j���ý��j����]/=p5Wz+G��b����t{l�y�̐3�z�����H ��Đ'iL11�><#]{WN"���nǠ�6���4*8�����=�R<4{m��;ٛ��1V����jr���w'Y�I�#�P���8��������dA��~������b�s=�{3{��wr���z'�ݞ9US�xz�*��Y"�~�W�/Z�FC^�o��,FD>~�c3[o��6b��i P>��<�jn|�O*��=���<��M{C�8�6�x[�7�8�fˑ�s����Nռ��2�٪�>��R����9�ٹ�{u�����@���~��ґ�2EE�Y��AB�K��J�������S��~A�Q�O�+ɢ2#��o����`wg¡x\�KH}�[���,����45����n;|�ӿ;���W?\/:���l��hn*r8u�	�S���gK���U�+���������垡��!�y���	P�H���S������?���g�K�Z�0'j�<��n�����I��@��֮ҕJ�Y�4v�	�	�]�7S��:c�]d�=h�%�7��k��ƶ.�;{����hjuੁ�0/(ԩ��+S�j���G����V�Z��J}�l��%��&����h)��W�`7����nc�?^Q�n�wQ�ϝh>������������ܖrh���y��\ځ���
�M^İ�ND����V�i~g6y��y/H��D��!^�e\�����j*�������m��#��<tV��!r�L�3'��nM�+��qN:�� ]�z�7�ҽ]�E���]�����oz�Y~�?ZQ���Z�j�%�����|��s�w��<��[�i���;ЎdR�r+")����0���x��*���Ϥ`T~��*���˲eԷ��/�PsJ�3<�${�
h{��.
�Q�W���:�C�WH��N{�U�^�zD���st��w=�I�#�r�@L\BG�E4==�QC9�pr�6"}����z�g���~o�����̱��~�}jx���/�UY����T�b�\�x��u�R��>�!������o<���Y�O~�󫩧nꂖ蚨^��F���z�[���V�X^=;�Y��\���'�J�k9�9��*�=���󼙞�캑p��cD2: {n/��k�W����j�O8"�o�O�򶀢�t�,b7��oO]�ߢ��yL#O4:��z�An.B�[�}s���qd5�)qSl݅����*
���Pp��Ԕz����u͔.6H���)䡓y�Y8>g����+jM�s��W�p�DC�Y(M���7����s�g>���-��}��Ͻ�~L�Lg�@�ؼO��iTrv�{�;���e����;�o�e$<�|Ux�ח�?'w�6����lx�������v�������Z��1��X������OWJʽ�!��8j4�2b��ú���K����kɜ�ɸc��f�<�������"�dG�C�g�Nv�WKϪ�pt�*�!��uyg�e;^�H/=N�Um=�zCz;I�$�p�yU��w�Ċ!I�U�E���JQ|��q`�܍�9�o�n���﷓�#~�_�Y��ݬ��YP�L�K��R��:p�߬{е��Mҳro|�����)zI̘����NF��xv���|�v���+,��#�Hd``.��h��Qz)�?Q\7�8^YW�Ƿr+�!�̇�z�ü'����d�#!�ߤ�Ee�Y# ^�����9�1���q�˭(��^��j'U������γ�^��?Sy��S����T�s���=�=:���Z8Mq�j�d�/�&W�9�ߤdM�;�YCm���}^�$#C�b!\��Q�wr���e��"S��.��૵W/�#�s�d�� E(�sf�	~+ f5t�ֽyג�0t�J�6�:���
��̇��%:�p`���v��P�T�v���;��]m��12��C:^к���-l	� �u��w�d�H͎A�.�I���v�M�*����K��H��	�4��wCe2�I�h��[^鉟n{�̠{Em�'�׋�|7@��qV�=�u� F�K֬d,���P���|6�{�##|ۋ�]��䲤�D{���G�hl��Xu�ɞv�mS �H�^r���jj6k�[�uǐ�)���H�k!�a������mߤ{b'��>�{4��R.0�^܇�����p�:V.��<=[7��	����4�����y�Xϡ��e���\���=̖=3�T�Z�5{�p�x��
�{�d!:����Y/�Ӎg����{���}��b��(�&�w��c�Fz(��B���N��ԸR��=!�W����߸۟g�qlzwgѾj�ˡ$um��Ȫݺ�^3L>�+ɣ�׼"׶�F}���B�ߝ�|"v��~�?~�T��0L{��Gg7�UX��L�n�R�r=�zb�e�D��C)�_T;S���(t����e����v9�9���qiV����#�-\�q��1���S�){�7�~���Y�����)��.>���߱�;�htޠ��i7��	j���.�k�`�t�R��W��o��X`6�Vܻ$���E�a�]/0a��[-�z��N��0����hk�,�fP����bfK�w�b�SI�ۑ&�3K=C%;&V���9����k��9�$��B���{2]��*c��0�e� k�nQw;�(V}�*�=�sYGe'+<�MCE�y�rU�-�
ve-��M!R��+�]�]ə��������-��T�e�b����n�|%�]���w�"S�J��O�9�«��P����v1�oo���m��HR�X����n�-�v%���ES�U�F ����(V�%x�~Pz�����PФX%gTP~��N�b�Q�w���\�N_��Tn�T}S���&�f1�/�6�l]t����J|��R��㴡u5�������%��1�K%s�ӻH�VvV�+�� ݴ6I���;�Z�Ш�]YPp���եt8m�6�����
���
J��!Ͷy��v�.K�1�7�I-'K�խf�5b�6�RH�h["l��G�'9��.����6_R�z�=ו�4+�С.3��s�%��X7��CR U��JfaY�7���;6���ю�z��w1RpuR����m ��W�LLʸ�Ƹ㕴��2��7nWcy���@��6L-:y}�a�ܯ��$�q{�T��@�uaN�R֌��nĚ�I��r��v�zF�.U���N�dA��5���m�.�Z��r��6��̵�����"���t����-�O������Wp��9��F-��Q���0�;�'%��v<GAR6���3.��v�5�L>�ok�E��7�)1�r)�����)6�Z����6�+[���wU��\�[x@���
�[��r:=��Z��2��د&��t���e�?^s�e�P*sb��{n''j�*t82�:��2}�E 2H�Mw�U����=I�(�M��7�7^:U{�ܥpF�E;s�v�"�d%Y��uǂy�'���:J�, skq�
5���,�D�TN)Oi�/�+(ܼv��U�[\���!���C97�ju�.d�w|%nZѴ�u��A�������Y�	RYÚ+d�ú�y9L��	l)����u��1\Ifᒮ}���\��
�u��b��1Q]�	F[s��\]Pq)�Y;��Bv��� �w��\����i���v�m��8δDE�`���%-K�f��Y�6V��ymY�hSh:P*l�na��U�vf�!:�]y��
)4��;�	�Gn�/�U��"�Ac�e����̭1V��Q�DT{R�;��wh|��,hq�>q��d�du�P}ٜ���$Mͅb\�h|6X�+�֕����j`n6.����afZ9�l��E͈skU�v���Y�v$���ao��X( PݖZ��IV�;�R�}�vW|�9�*hږY=�g�R�G=#�SW��O�������$CB�ADE�qU��"�UP�fAr*�p�J���9Ej�D�D9"��Tp��5@�&QDTUEAUV�eDA�P�D�J�`��fM6�r�3���H�L�E��!$�DvEG:B\�� ��HQ(�+�����:�DQQ��(��*��@�"��\�\��ɪ¨��&E\�*���e
���TY%Eª#VQU&\�UUr�(���(�\����YETr�N�Dr��@�!	�D*�s�UQʮTUG((��"�r���ZQr��UQQ!DAr9G-H�W��ADEr�*(�\�Rb�\��.G �s�UA\�>w���侖�pe3u:��$�NW[�Ԫ� �J6��˸�P�]�R�sV��n혭-A�մ�Gʭ����.,�))X�~z?G��ḇ�r��߁�d=��_��t�<z=��l{zN�Y�ݙY~^wշ �]�{�٥�T.}�: ;�2�i\{ �߮����5��N�����|��^�J�u���o��F�|ݵ�g�{�'6�ARW(�����
�W��y��g.�2=�����zL�/w�mV���}�����Q^�=Υ���Yȶ!����3�!�䄽U9��L�t��'|5z��4����r�}sSyӾ�_�]�<{�Eǭ�,������+�E}M�ō��߻Gy��^<�V�E��;�B���#�V���e���d��9���E\*���̶$f/(�2���x�=���}[���Hx����������Z��m���������d�1٤��h����@��'���'=7�,�0lkT�0������X�~� <4{�3ޝ��Ez~3#��5�W���Wꪛ��R�d�m�$\���Pղ1�vG��y�X����um^a�^BwlH�Ϊ�G�­�9��T�?JiP��lL3�5�r#�t��{o�EU�txX�L��ԓǼ�y��Mk�3X?Vʿ9Y��W�4+c��БH&��4�)g)�ѝ�כWz)��zR�w������7��!�SOAe��0��zJQ���F��գbњr����0�BOp���PLC��t�.��:�1ک�8�B�te9]U��S��d>u.��<n�z�no��h����;B�C���v�9s�/%��ҕG7�FֿKTl����g=.p�nzw����>���y^M�*W��p�0;��P�<ze{�dY��j�i��ui�4R�Ǡ]x��Qw3q�垝�ww�ꮇ��[yfN��3q����0�Z���C^�q��"̂;�Uv��Q�Yلh�1�k�7��=C^R���`�;�s�3&M�qc�0�aT����r1�C�*�;q5FVA��]A�S�Sީ��z�#���'}�6oE�j�XO?Y/gLi��9�P�U{ma�A���Z|&��3>��g��ג�w�ǣr62cw�����_`�l���v�����~Ǒ�+���C"00������67��,�A`o5�+�u~�)8z(�v����a�>����e�������ϧ(!hx �T8�U�����'�Ep��9�C��D-��2+�/�9��{��u����3�y9���Ϥ`T�]�w�!������3�^��L�=fA������s�Ȭ�_�!��x"9�ّ��������b*2�}�[�����*�z�B���qWY�J/�\�ȃ�`��.��aͼ�	S�R��w��z%E�x�*24lC[p*Ա,�w����y�\ָ2f����n�����/��f��a8�X�Fl�`�
���l[����eO��&�me܎X׳p����W����aА�E4==��29�pr�6#}Zs�z_�sw �.*N-=�F���@�w�6k<*P:�P�DI�5���\��l��S�g��';��U�6Ex�U!������Uo��{x��Σ"U*�P���^ɥ�.6��X��vȻ���9O��7����i�I�n��f���ۿ
����'��ff���E�`���dg��p���>�X��Ĭ�����~hye{�����Ϛ��-���}���C�zh�[W7�n�_S�Q�
:g[�'s�e�u����C��~��+�y�����sӰ�ߐg�3�4�v�}�˟38oY�]�bo���)v�Ah�'�螮�dU�yL����Yt+�=A��8̪ql�vssQ��U8���{�x?
џ/�8vUx[��n��t_?�����ߺ~ _M��W�6 {;�����k�G����;����j��C~��	h�_Ķa`��s>{�gS}Ro}~�ȭ<�Y��;�u��k�����wJ{����U�@��}���PyS��uJ��q1b�,�=�����t��>��"��~ U�Os�Mvn��l�gi[��C�pKͩ�U~��/>��i>�!vW��YM/.	Cs_Z��<���r��Rc�y@�P�1��J��Ƽsհ�f�.[t7u�p	�G���C]�:ͥ9�b]�{�Z|��ǭg������T�fL>�z��c}����f)���+,��B;u7a�8?yF DT�s��j{I���n7>�U�YP?sy��_�oz����{!����$]\}&	?s�ᗙ���e���{� 
��5�촃�n�½���{���O�#{�,C q�w���3���|�WgvE�}Y��+�?lx'ŀ��U����ܘϕ~�5�^�)�|�̲�bں�2����_���!��xz�g���`�	����%�Bw�U�5H�$�S�r��.�v_��.�w`g�r}K�N�=�=;�ܗ�ϘxR��x���Ao�!TT�B=~���U�9��g�^����{�=8W��v�hl��X�*����R�9�Q���U���K���G�/a��{+�����|��f�`���=���̟:��Б��`ר�]���1wR>�.}��3�ճ{d���X�f�_�#��<����c��d�25�S/3�hV�Qo���Dv�xD��)�dO�ea��v �Y��5��7!��#���۬?y=ɜY5{��$!F�V�YN-EWX����lcЭRf��?p��5BT<Λe���Ĕ��x�uݣ��/��Q��6jЭ�m=�n%�[��J�B��Җ�V7;By{s�z����;Hm9:��I�PVR��䴫��$-g�/!�o����jM)�̎�I��:B�h�T����'kee]�çac��N}S���W�!R���+u�ߣ'ڭ�����u��/-��L9S�\�܀�߂�Q����~7�M���cݱ�M�vA�9�♛���Nÿ_�d?_0v�$��v��o��n`n�¡����s3�}�UM�W�N��7�y�.���O_�gW����>t=ˇ�>^Vd�����i���۳����eJ]��KSJ��>p_ǲ;e�9^�lI�CS޿��/�ې��G�MZ�^"�n߽�J}��{'���<$�I֗��_����u���+;��zG�Ӿ��a�3(���}�KĲ� m��Z`�[�E^y>%����@�W�ϗe���M����3F��(3��%Q۬y.}�ۜ�}R�d?,�d[��-	�+�Nf�%�ύSn�fw��X2Aõ�|�#\w���ԏ{ײa>�0��i_�\:6H2�(Q�'�.)77�.���$7t���ʨ���.
��'�V�@{~`�?Y�{�'o�]�!,z���j0��w7!�5aR��q�!�ژz�6�0L�Hۓ��vȖ�t޸o�䭙ZT�R�;�g��	��4��ZA�[8�n���]r�j�����
h����T��rk��)7K�]c����g,�tu�˹u�H[#�T��иS��E̽��MRV��h=_1pP�G��6'�ϼm�w�9^������y��({�݂��3鯅R# u	����ެ���j��}�B��k=c!������QF�^�Y�n󷻶�|.|�꬙�uU*X5ª=\�e����^�i�dd5��q鬺[�]oW��Jl�v#��౞�z$�]���J@��dc�AR����}�?�]�5Z�ٸ��)^Tg�O��fɟ{�u������ߛgߝ�g�����:C0;�,���z�����������
W~�8�Ӈ�sө��}^���T�{n�x07S���`FxF^Wd��<�0KU�{���t�7�i���g�]�������y���yq��e����*��{׵���	㼻|�/}��p����vos8h�!�i��j��N����W0N������z�u�r�ES�>�z�́�|���b��->��CR����W����a����u�viș��Ԋ�}�^�}�M���ER?8�hUH]���u�62Z���D>�_�f=Z��q�.����n'�m���:�S컪������e5;Z-�m�f�u�gݠ��C��Aʺ�Wq;=t�r�q�I���N�ӻ�Gi#.�po��MV�w�0�'�rZ��7�����<u�1�9�L�� �h�1ֵ:95������o�'7�����_��.=�*�E�ۢ3 ��V�=8�W���!�87}^�[�q�&2���{�^���̳���|F�YP�n�0-l�V��\��i+Io���dO����e4=��Exd_�r+"��p���b;�2��*���jI�H�yz���ڢ��3,�ѩ�_�����s�Ȭ���x":���5����վ����	��OR+��<�h��eU��/����T�9������9>��oy{�k�}����= ��3��m�1Sp���g���Bw.�EI�KÜ�>ƝF�n�&`Ƕm׷y����T�wZ�m�xz����P��M�sU����L߬u{��K..�Eg����P���6(�>/�S�Ͻ�rۯ �ޯL�o�6fj��E�*`�D27���J}��UUsif�t枥��B��Dt|r����97�q�~�����g׏��3���n9�ԅ@x������f�j�,��|�|:�ٵ��bW��p���dy�\ϭV��;qE�N+�����>��#�H�w$vYi��O���J��W^ʹ�ʕ���h��%sb`Ú�4voy��2�.���~������W3���f!�]������p=ݘh��fsy�4-#Rr���]ŏNk�^l���p��cl�ý-�M.�C��/�z� �J\p�f�sӊ�8"�m��{�u~#�!�%���S�]��"������<Ȯ�׼.!�V���%�����╳���L�^ ��^_�}�i�3=���^n��홟}�^9˾YC���9hW�ݫ%w>LK+�ZM����,>r���y9�ʃ���Q�I�7�_�NBk���x�����j*��$<辡��~z��{m���i1܊�َ=ݛ��\ϞğfL=��`�c������S�;Yfn۩y�Xb�`Z��{�0�{�=C����*݇�n�7�b�����|o{!�������W�����P��Ư�;���) T �cƔ���iN�9u�~��-ߴ�G�m
�M��^v2B������v|�y#$!jϕ�s(zFp���n��[���E��~�3�b�?_i"Z�tV{&3�Y����x����z�V�L�X����j���ٓJ&<�l��T^��T���دy㝏���a��ґ�@T���8����;��
x�PU�1����qJ��k\|�Θ�r�l�,�!���x�l>y8^�V>#F��ڥ��_�*ip���7n��Sx���K60�-̃.�^v$ �z�Γ�o��c6h*�=��s+Y�Pnn[ISxx³�flY;�R�j�&��ŧ��v����8矼G�S�l#��Yʞ���r�{ր�ϫe�鹝V��l�ݸ��b�s�WB{�IMH��#���E}��������r�G���f�`�ۿH�ϯ�2}��D{ۊ@t}Q><��%�s�$z:���Q#�����=Axm��#�d{a���W���Z�|��ΕsƊ���#"{�'��ɶ=�A�7ᔧ��[+"_�3�AƳӼk�29��3�mu�\7�}��w�}��jf���P���|>� }
=k�:Vy/�N�����w��X� Z�W���wW�ۂ3�=��̅8�~���U��&�u�o�T��w)��*�*/+�K��Y��^3�G�_�@��#�!����v�g�a߯�3����\�h���۩���Y�h�z��&�]���p}}vD����z�3+���)�/z�ǲ��3��fK�2��.詃o�sk_�w9ڶ|h�T@h_�Q�Z��fVE�<%VyWl�`w�Rc���`�j���^'��N��=
xo�1g�R՛��Id7������_�����3�^��g��#ʫ�ʴ^�vױ;��XQQ#j��*B�d�ͦ9F^�t��~��hB�0v�њV�R�߫�����!�=y����}�Ϋ��Fޫ���Ӄ�0��3�u܇-�s�,V�<OyP�@����@�c��WU66�ْd��#�uĬ�w�D;��2c���}$Գ?Y��/rߣ�}z���j����O�~y&�zL.˦*���v�U�.��ܝ��>s~Գ�gO���#}R�c��gEc�r��ϕ��3Q�T��A���yc��&�F�_W�˅��a���o�ӿ'q�-�3�6�G�O�`d�kD�Z�6��)�'ǎ
�Ïxi���z����sQ�>~Y�,S���|�fH�P��������;W#{=x�G�����&S�4&����h{��r�>������>�e9o+f��V��ln�y�?����?Ub��u���_�a�B��zoae��5O�;�\�5��;��c����/�n%{�^��u羽��V�o�5 G����-_x\�b�{ղ+�yR�7�U��>G�lp���Z�wҚ�����E���M(��K c��~�F�kU��^\��\����޻G�򴠬7�����o�|��\����Ͻs룰�w4}Y5<�Lp`z�*j'-���8�f8�s^�)�p�
��_��5���N��lC>�J�ɮڹ^ʩ���K���dy٧	��h�ӝ����A
��mA�e�u��$i)�a��J�uJ�:�����\3�4+.h��p�]pRF�+��ųi����F��F7vbZ8�0�i��2�N���+���qۦ6)NN���Tok���7����Mf���F/+t��J@����+s~2�wu�'k\�r)�ip}emA{R�Q�O,���(���⇲���ݢT~��}��F�X��
B����y&$�
|0'��b);�{�w_u��,d%�s�%u,�a�7�?�R��LKw��;�)Ӥ���Q���Ʋ|�A���kZ8V�M��H����8,|��AhS;u�Ho	:8��r��?�ú�� :� #��$��HW=�V2V�<�*vq@���0�6��\���J򰽥��ߌ�C<���P�(K��;��У[zJ��吶����RSg]n�f���U�dv$��T!��wMa#�����f.S�ח��OVf�${�mx�f�'���>��J��� �u�WP��}2�j�.4�^�m_0���S���>���\Άn��H@Ք����O1���]b���,ɅX��9u=4���m��d�������e*��-)/u^����/�P��]M�(p�r�ퟯ��7:W`�d9�=��eO��1ʾ�#43q��ǚ�ځ�w�/��ӫ��
�P������/맒I"��`�*ȌwA���$����be�z��i��"��3�ľc���qp�;����x�%��۔�gW_e�q�5>n�#�*�Jط�4j0�m��w����l����QC�g���U�m4�^z[O�.�$�'jp���)�c9"���Iw#� v�{;�؏i_lT���$d\'T��Np�R�Dͨeڨ�r��ׅ�\�axs+4;��l�Y$����Ȕ,ZٹP�FPᇯr%�8���>�.쭷���������;_j[��huEƥEj����3���B����	X. S��2���w}�Z���]Zz��ͩ	�&VV�H�]*�\���nT��i*WM��JdT���q�V�Le,}�TG*� ��⻣�%�\Up���*��N�g�&W��թ��8gp��|�t45�vq4�iz�R��V��Ѝ��a�.3���[��f�pح�z�K�I)]A�F�;�[к�ur�+-k$���y���c�7+j/�z��BĎ����Ӌ��_v�HV�ի+��F�ά7�jR110h2hJAL�E��ض-�x��S�2�c��onp5�����us�+([�KxL�5Y��b���7|V��Ŗ!Ma�W..��fG�/+Gə�&ܑ��f�#��'Ƿ�`�Y��R&�Z$bÙ�7P�_%|�w� ��:�]�n3��(+��g��k��Kz���D��]lB���X/Q���|��]-�T�]�^�����l7��N� �  T(U�UT)Ap����"��
E�ʃ�(���AQp�9Y��TUU\�r(�"����r*#�\��L8QE*�r*��Ӗ\Ԡ�J8DF�R***"�EQ*9QG+�UW.EU2&Qv'�U���(��L��*�9˗"� ��U\�-J�*�*�r*��Q��9U�QTW(��fvs�":c#�Ȣ �#�J#(���\��*(��G3\��Ȩ��ZA"�Qr�DQDQr ��*
�����&ZҠ��������AQAQ�(��+D9r�*��*���TG*��9Q�+�G#�r.�ʈ*?^}�t|��c[�/��̹����¾�0�����\\኎��L�Vet]v�vP"�E�ځS���o{y[X����������j�q�3��/@hP�9����K��w��C�����.8燡��Y)gf�8���Dt��mϽJG��P�C�{�F���߇S���~��xxG���J��'�^r��l��磴�RLZ?0�vg�~�=n���#�
UR�ϝoýs(B�S���zoܗc�5r=�3����{+�^�w�z�\iۮ���+��T
��+c��z³q���<y�GX��+��_����'5ǯ���~�Z>�YNЬ���ejK#�1�">]����7�zW�.�FyO�]���n�W�=Ɍ/�Ν���؎�̳����lVT+��Q���;yP*��u���*ԋ 
�
�CU�6=��C9�^~�Ȭ�������dy8�z#��_��{��V�y�9葀TxL��\R��J�#~"��f��Q��+#��Hl]���l�b�Z���]B|d�;����U!p�P	w<Vߏ�ⷌ��s�P;���;��@���f�x�8z���q�Oܑ��#^�P�B�~҄����ۦ�l���3z�>�,
�vn�8������m��C5���-�B��-���s�^N-N�@s3dcK 3zL�����,Wz/*t�֋�#cտ0Zc�N|[�}eʁs=�ALr�]��z���K�ݎr䆱�
먷�켼䃒�I@��{���3_s�:IG&/t�G%�'�W��X<4z���=q�4��M��75P��GD+͞w��Wf�םF�7��,���cݔxVC6���*}9�̹m׀�����35��]H��S ��=#���GǞ.�f@�\[�XH�R�7�r:Q�[����|��3�����ŕs�.�S�r2}k}��X��>���N�#�T#^�Ь2<C���dA�܂�^!3����/���F�¨}�vr�W�[����&:���tmp�,��U�zU@�b��{G�\i.��g��ʮ۫����AT�{�����/����>�,��/�C�`�M�8,��
�l��z�9��^��X�g��^�H�e�a���W�3�U����TdO�S]�JTq�}���զ�z���s%���o�^�H�ׯ����u�$l=���ј=��˲b�j*ǋ;u���]�އ��
W�J��̷�'ٓc���s�u��~�O����yVY���u~2�C,q�u��:�jP���B��F��r��=�-�swp��p��T�>��C"n�=�W�x�ן2_�GAR_R؏1id�\^��Α�Y�#6��� )����%�<s���R�ޥ�9}�uȖy�U���	�o�)?XǶ��y|Ą��v�&4X���Wj��#��+;.֣9����W��7�%�v
l�sAgm��x�dL�$���~��'��^�<���#�?���x+��&���"���I~�B�o��Z:����c��:�o�C;�a䌐�����Nj��XE6�C9gÄZݪ�;���㕧J/��s�5�q�N�{��h	��=끾�bNPB�	��z��PlЛ/bk�{v�ck�b]�]Z�g|�o�B���b�#�v��=�='����R�����p$�A�`ߪ�A\N�v�5;����={c=����.沧�?+S��Z����2�<���X���=��_*(�`\H��:��s��1־k!�g��\��������W�g��Md܎��'=�QQ�:��;AP�G��sp*�V��oc�ׁ���22�d{b=�cq{�YL�3�E��]�^�ǣx��{�̛#�T.C
�m91��
=��^����A9�l��m��k�r�]ە=��������_�-�<n�z��YVf��U�D��8&��̮��\VwF������ә��N���~Wk���W�G#�f��{n�gt�^y^�|�+S�.��.u�9e#5����s�e��Zu
ݛ�2��-��@=�7�폖+.�.��A.�m��:�
��s&�� ��'���:����)uau_
9�o�i#0�Y�����a�ZMj�k����ҍ�zC�pˣ�O��s ���ە8D{{Yէ�\#}�[���fGo�㙛��,��;��
��>|�$��v�ﲪsc-.���߼����G��#�xs��B��#`]? �'��3p���S��C~�\w�o��ԯ}y'��^��޾Z��s��J��>������S�U�(�,��̰l8�0��2�����	���Ξ��cˑ��-������TU#��]g�1��K� !��S� �ߎ]����ۺc>���q�}�a�<�خ�f��#}c=�=�����.=�#�E���F:�)���;ׅ�>>w�^�ә��S\8z��μ�Ͻ�g���}�=�޹`�?<����'(!hx �S��,Et�1<�<f;����X�U>�U"�~�ˊ�}�i��߯d�u����<z�������ff��Adx�ޘ��
S3_�@�U��j9��+>��j������~�$�z����Ay=��V$T���)�}�C��&[������)��sQ�(���������=�km��}*�C�Z{�D�3�����j��u�������S{��l=S��!QυȊ�|*��?_��u!�lKl>��2�q6�V����'j�����Ը/�7���F���ee��eW���)w:]b����4ʶ�M;Əf���@��*󥌽����C2����rQ��o�fɕ�v����Wb�&��̊G}�]챚9 Ǉ�|���:�US ��P���f�m����l������غ�^��Һ�� �'��̱�`��{���w�$z� ��L�C95�]ӳ>��q^��|mCS��jה�垿{q�Ij�%Ɇ��s���>�Z�w4Ud�����E�0=�:c&���o���V����숫�wY^C˾+=&s�ٹ�N��>�9��٢=���1��2[��ON!��-v�T�GQ�"Fϼ3��q�[~@��d���b�N�����]�Ϊ�V�M{s7��R1U���ۭ���#�d|����W��M�P:�M���L���[~Y�G��[ܼ���u���;��U���1��m��{Y��o2_(��%�w>tVx81�jn&j�s5���(���p�R3�ׇ�o���u��']�zv�``y`�;r(�>��dz]�.�/:;{=^v=��f\U�Q�����=~�ߟ��c�j|dY�*�Q����S��,��m�N#�ܝ��|=���G��_�an�SϞ=ɇ�{�ӿw�����|��ψج�*�s�r)b�݊:�+��=�u��t�R=��(+(d)�3z�x3K��l��.[�ׂ�bu
�p��J
ꉁmt/] �k�'��b�#����^�Ή����o��E����왎i̫lN����N�D�{B!W�B���|���s-���pܪ���C5»��G��p`q���U������_�r+"��p��:;޹�C���C�7dj��Vf��!xI�]�^}# ��*��*����@n�# �l6j�_[�Ȭ���Hy�#�7�E��w���pj��xz��1J>UR�J���ё�E?=�1E��(��j���>gQ����G�N?��m���#��m��*mU��D�%yU�_���Ow�}^���67�S��WS���z\���	��^�ؚ�n�e骅� ����[�Ƽ�Nos�#�߱X߻)���5n}��*}9�{�2�w�=������ٙ�캑�h;4��9��]Ί���X�����H6,��/b�@��vzw�w�3�޹�^D?g�τ�(��=�>͌���E�+;�}v�G��]6|F���s�H؃���W�ȃٹ?]���U�;[���9x���^�7��*+�h`�����/�kåX=);��s^�8(�4����W ��O�i칭�o��d9�z�x>��̊9���1��ѐ��,�%�:���&��_��J��e��K�_e����Y�.��9{��ӮJys��yt�`U��v�(�^�m-nY�^��$����й���g&�s�L���{�v�$�嬷�T��l[s���3��&^s�2���!��Lnn�d��N�jL G�v k��Ǩa�8QJ��`?C6�n3���3�׳�=u�_�$�XD��p�A�ݟ
��q��^���e�9�n����'^����y�4�g�6�.5zׅN��{=#~�_���%��c�ώ!�c�����ݖ��n�t�f��@��G�,���\�{}�0����u��W?m�|�v����A;:���g]��yU'�D E�1@�p� �_�=[w4�sy�����xO�؜�^��=���
�ǧJ�
%�%^��[��YfTM��z@3��nd�6=)������&����^-�ۼ�1�U,27�R����fE��D�����L�\@�5�T�+>"�g={Hg�n�X�Υ��ʺ����~�Ȋ��ON��ƇA�O�������'( �fR�P�'��f5[��q�)��BHMo��)�Z�+���9�a�O/���2=끢�=~���
;��
�>g����H�e�z)+V0�4�.�kjL�~x�b�hG�K ��[3�}��;,�{�|�:u���o�3� �"���	��X��7�d?�*8�k=c�jG��5F�~���v���A���
���)��\�w[t��F�}v�Lľ3�S��K������T	��!or��^���rc��6��Bf�smD�*�7��s50����	[�U�Y2�u���M,�L�N�����s��t'>�g2^��Rs}���I��ݵ3o�C� �3�*��[7�����ll5L�kݑ�>�u�.r�7�*�/,ۭ:�SF���{z��G��>؇��pG��Z�aU��''ղ�Z Μk=6���&_=��U��%yQ��=��܃�z�}�`�� ���T(�Rt�ֹ/�!�)�ﳫ�)d{;��ǩG���;���|�[ ��mϳNfϧS���G���~Us\��no��џp`wg)̭X�F�p���fz&����?Vdv��fo��,��;��
�~����I��2���7�����S]W�(7ǹ��T�m0;�G�o������.��{���fWy{*W�){�=u�r�>�e�'�Z��X/��e~{~��5�;2��x�~�F��wc����|ğT˔������dW����O�8R9��˄���d�'Mm��@U)� e���Ӕ���>���Mc"`U�?;G�J��+��σ��^�[Ǒ�+��B�
s1>A������_{NyRF�WD.ۢ2!�&�g�ΟG���A����}�s� �Z������H��~��jV�<7G�t�я�u��V��UӐ
f�,�g�?�s-H��(˾T��4,D��,��	W,���ʻ׮�:���؍f#�LF�D��Y�︛���ɀ帲%�9'�ܻ��2�m��$)�R����U�+ψͼu��܆����)%��w�g�=�U9ꦽ[��{"��3S�S~Ν^������R0w�����u[��^8{�U#��=��b����x=P��C9�dVz��N�}~@�WO���D�'�-���G�VxOmVMyUJ&e�>LSvddA��t1pP�������6M{����7��n��;G���g߼�^S�?����׼eQ�DO֦�[`��)�_�Iq��}�錌��y�������F��Ǽ<��p=[�=��f�un��K� UB�*�ݷg��O�A�z�rpbw8o�$z��b����	�yfX�m����'βg�װP
X�jݕ-b��1���+�;��LG�[��&�{��7�-]�-�2�z��K_�抬��yU 9B	�I�\��~����uY5�!�Z�ᰲ�����9�sҝW�Q��6��6h�ˏ+���x�ޥֈ�����x�)��b��BL���;lߧ�����Y�V�N�Oo{ږ���u�C�^�yq]�}=մ7 ׊�g�P_;= 8��U�~KUo��z����1�^�T�����3Uxw��ϦMuӨ�.�*����Y� ��-���\\N����Xb��VoE�I
٭R��F�u�x��h�ɮv�$�7%�j��A���.�xnb�O9d+���x<t��$��\����J��&���MA���s�)ܛ�����&_x?�*��$�pQ��UӐ�C�eS������9~�fYާ��j�s{�A���5��Ϻ}^�S����x���']�zv�F�
s��ϗ%���O�{}��eٱ��~��I�低�H��q����{�}_���o⦚�qj�u����K�K������ ��.+S�.ݺY��ǹ0����{�^���\�9��9�5znz=��W��ƭ��r�� r!ĘV�r[���ExW�n(7~�|�ޙW1�j��3j�ⷂ���1��N�;�+"F X��*�S4�H�"�Y���?+�u#�B��������;{�a��O���ۏU�W�� �T���bj��#���b��z��Qx���F�+~�{��z��wn�(>H��U�V�N��3({j��~�Þ(wo�����m���w�T���z\ϼ�x8�`=�\lK�U3�����ͺC�7�C�|9j�wж���X�ܦ�ZUG5�.r������.���y3?��#`���[���� 7���������nl6��`�1��S����v�o�0l����cm�̓`�����o�0l�y�l�[������cm���o�0l���`���L6��`�1��#���������PVI��h���������A���y�d/����v��A���DTUBD
�DD�$�I(�T�UUH���H� IEQ(E"UIJA%(�*�*�����A!@��((UBP�R����)%*"�0*RA���$*���)������Tll��t)P(�	)T�R�%�QIDQET�E �J�$��I!RJ"��T(Q)@�*%"�US��B���!�   �z�U�m��n�4i��SPiv݃P�
҅�Y�����uF� @���h�4j�R�MMeh�T��UR%
Wl����6<   F
(��R��'K4�V����n(���QE��qEQ@Pc�q��(��(��3�(� ( �tQEP�ӫ��( ���U
"��{55U)$8   �� z(��ڴ�hd�h5Fֶ �[l�@�TZ� 5�5h k`ªMY�� ˙ERT�h�4�-��  Gu���#��@�2��j��  Z 	mS� ..��c@ڱ�mV��kf�@�*�%T�H��
@��  ���ҕ�m���[e��-M�[{���;�����1�U+M�ɍa�J�
14i����Ftv�N���ۋ�l몵ê�!$�*
�"I@/   O=�EP�ڡ�;X
�MU`�]N�ʰ��Q-����a�I
���t��쭚 6ka�uՖ��Ӵ�e���ܚt�6�6�!H5)$UAP	R���   ���E4-;�uju�P��dэ��9���Z�`ƚ�� w"����n�6ԫL+5[Q��gv'S���R�*�"�ER TljIH<  f{��@6�f&��Rm��i[��ii�Z�v�&�uvִ���J�ʤd������Y��ww)j�[-�t��Z��6���J"Rm�B(�� ΝCi��m���(*�֕�j�,)�Pzζ��Mm�J���u�ج�
T��6ضѭ3Ki��Y��"����HDRR����A� ֒5@[X��v��U����[ ���RU)�a��Z5Vlʳ��ʣlئ�ڷm.�Ma��&ƫY�U@u���d]�(Q@���"R��i�ʒ�Q���Ɂ1�	��"�ф��� ��@  �AT�I�P�   hh   �~%*��       	F�¨
i�jI�M4iMF�4 �i���Jh2�Ҟ�'�������G�3Q5�@�@�Q��"�&b[�%B�@bHa%�Mq�r&�̹��n;|�a���m��>L�HI����C�B@ H~� 	!&:�������	���<?��	�����.��:�������C��?H2A�	x ��%? ���~:�			?P��d�E h@ z�W�����䞅�vn����}?=�=��w3��}y����4�l!!�H |��m	�I!�Id� m$�!�! �`@��HI$�HHx�&�B m��@� �I!��&�!$&�HB0 @뮶o{����)$�K���j��{Րb)?}g������$�$�����w�5�8�}$=d ��g>�G��G91�%D:�5���<}�DЕ�p�n�޺��G���%��0J2����iyI�U�K�ݨf�R��,wÔ��o%Ds#
��X4���d������\6v-�%3�Y�#%��C�se-q`�i�Q��lk=XK?J9xS�����A�3j	RJ���,�Xi%^S����A���`�&-z����J!o�l�ww#�
�u��d�/5�`R��Wjj����Y�9P#�ЈT��.�`� Vܷ�����k��'yv0�3H	�˭���##TW���ތ��=Z�T���4��%��L�FS�'h0­f壶 �M���[�P�ul��e�)S���*��<�zJ����t�:sn��J]M�ۉD�l����	�j�Ih��٘Ͱ�J�e��ǆU�ө���`6pF!�u{��i�R�R�2�j3�
ykw]%+�FD���� ŏc�a8h�y�K*���v��U7�i�<,e�
ub�PmR�+\�B�jY�	���/K� Y�t4@\1�k/i�e��PʏE%�:�h�@Y{x����P9��Ĭ-��,Ԋ�Ͱ�,m�`��� W�;w�������8D��j2��"�ڵ��iڲQ�wX�� t���E[m���׶�*��z��)(�RԞF�ʂ��x�MJZV���Ѣ�Д1K�Y��(4���I5.V�ֶV7�7{�[��1��T��QSq�k6��7�I/V+�Xń�
�D5�����P�idgKfe,��qi۩��M��ْP�a��fe������]J�hP� Dr�(��&ޒ1��nؔ.�:ïȍ�D= �0(���P�t�e9{��f��cv��,R%-�;Q5��x�# @�ʬ�bB�3v���-�p��ܫfXa��쿮Jh�e�vU<��gd��.DLKnۨ�A�r\�mZ1<�0�T5HZ�˥m��Wwz�וoQ{l�E��Pw�;�e��Bj6ְŘe;
�r��$��"���n6qV��&
�n�+������{Y��4I�R���X֢XS�6#L^����(�11�;���!:��fK���l�Ӑ5.��W�`V��[e䊬5!���c�(�I��1�tlS!�tt!�{��M�w��+t�W��Q&�ۀ$��zm�yiXڅS�Q��M� ��Ɨ@QJ�6I�j��{�X�L���x�yI
�\� ���h:�J�V��#K7h�I�m�-NT�6�G@�R��TiA���fb",�i�X,��?�[`���'-u�;m�܎�nd�n�WB1R��fm�A��FQ��fZ����@`|�;����[t�k�MiV�M͊+�DܻTh4�I6-U�x�(k&^ˀ�`�m�[�w�$�*����U��RR�-źrؼ����kC�1;5��&�%�+	<�*�"$\Yf�b��ې,8�a�&3Wc@e%I��` 1�s���[4�G1�Z\W���]�:5��EQY"�Z��gcc�6�*3Z�ұvQ�c�9��֬��G���`��Zy�M��F�+Vj ��7)�*�4���Ҥ4"���z�*��������Pn�82՗�1T�ح�i�y��âҠ=Wr\)���4��[�Q^�5x���j�2��r̨Ѻ.��
$cݢ٨��H�pYO�X:v5�y����`a�x�lP�骟�q]	Y&In&��:�[r�h7����-���@�`\ ��UmY�ZvE�a9�b����ƍKN��W��Eј�ǚ]�n�#�-L��t�M�:[A]�5���C� |^r��N/0M���6�;2F�V�:����T�sR�1a7f&�!�B��V�>z��YJ�KE`�sJ�n#�Q[11�AKDmZ�j;[2nZ7�C���Hl���"�[@��,H+.��f۬:�ڶr-v�y% �,���BK*,j��v�sO�d���NhU`���Dc�����dTV:�t��]MKN�B*�9�[|䂻X|��]R�(�e�2h5�����nRa�YX���j�e��
��*�2�����NM�@f]쫷�-������dq�1�J��T���E�.RvH���3sa�T�ʽIʣgM�e��Lee�,(nln�[�Z���).V�O L��;-�x�̨�R�!"Ƃ�/EfR��bB���K6بov�$���J�܌ԥ�k'j��V�QY4�e�����	��؉+HjI���u�0��K��f��w��� �o���2�%�:i�ˤ�)�Z�)&l �V�Em���)�P2�*�w��v�*5�3�t�6H ]��i�/$�R�vQ��"H�e����V��/n��n�.*͔+R]i�;uy&Ќ��.Ӳ���]�*�PD1*-����ibq���ʧ�U�ҥ���㷹��5��[����9Q�&�b^�����%�vhJk\˨8 �W;l�Ghfr��#�D`���4�w)1sd0���̭�����ɤ�����NĨ�X����t�Z����`G^�#0Dv^T5�F�uk�.敒õ�����D��m9-U�
��ݵM�r��ַ�U��,��)1Y�o-��4��n�\��c`�$�֛x�7T�	�fF3sl�seU�J���n:���P�h�F��'Gkf��H�U�[ȜY��(�����ZuH2��EB�6$R�E�,�����5��h�U�qG� v������3�.�J�H.J�.��u�1Fi�c�^��ن]ڕnSN��T� ��j�U^���	R�qP[�a�)M�W/�7�w,&�\��Ҵ��cp�Ktd��^
ɯt�Zݷ1�����LR�J�u]^ ��N٥��Йqn7h8�!��ؗ�%ż"c|̀�ͬ�e������g��Bչq]��^�K��f����U&Mv�`=n�$�n��֜�;{`�E�f�anm�U��xkoq%�-�X6]#-R�����7�12 �\�fMZ�Zd'5�s2����z�e
Ac�����c.�djb{u�7�r�ǵq ��Vja�W��*1T�]m+��w*���0�;��lt�<�S&'��V����f��\x�AY[��7w���{*ӽ��ַ.�c��G&-P'�(��`gѰ���2e�x#Uy���+U�5��Vj� �j��cn�Wv&录F/+c��nc�c�a�3m�m�B^Zj;��n�n���J�A2 vT$)�`&]�*�����+^��s!��E8�H*�Ĩ|�wZ���f��b-�W&j�խ�n�!I֔��ܤ��z(��ث�ê���:؞VB�,��*.�)c`�WD��f��Fp�;��u0��/VB�4�x�K7W���|2<��Y�1 WI[{�\� 6�ز����#�wN�h-�v�Q(��$&��X�F�I�n��3)�fe9V9yA�˼jV��S"�vG�am�]GX!ygF6������2��W[Y�Vn��NM7p,sV`z����㹸ަ��N�X(��IP�����0�'Stc͊��6�ڽ��7[��;���j� 	���+3(�xu�+2d�87V<�:�C:�^���O��˺ț�ۚ�ei��������{�Zǰ� ���J3�*5��	oS9����j���W�1�T��*�� �F�W�C�V�f%��p��R�`Zh7��F��2]�amL��nm��(�ě�;�*�]�Z%+�*Y@ѓh�u|�"N�b�!��[nQ�="��G!�Xp�Z-M*TpZ�Ҽ�W�!���f�H&�
���tda��W�]��
�V��֌��Q�JbEQf�@�K�
�=�����[��n��J@f\�؇^����Gxo����hM7fn��]U��V䣎��c���*Ŗ�QA5͆"�Xŭ�e�if�ܺ{Nm+*e�t���+
E���I��&$x��ԓj���h�'eX�ӧJ��
���Q��\Z�m#zJX�;*�ӨH�'�f�{��\q=�$��U�A�
h���n��ܦΚxl��r95��<��"^ݭ��Q�mM�ADh�J��*�*�g3/6^��	a�Z����4�yb��4ͦm��4���K���4�S9M�َ`Wy r`�o.��r��ZL�&��(�˂�1�ff�kO�iJy�E`�W��{�4fӳ��ԷX�N�6�w��O�TˎĦ���SU�$y��Kw3te�X�Ҽ;�t�)$��ߝ5�Y�a2��bZ+X����R�����%b��`�+ 40�׹J��HT���XhbeJ�R�L�S�q��n��U��`(6�I���)UыRSTSJP�gp
B[MQ���"`Vh�l�`�(�N��6Ġ�:9N�5Z�0�b���X�<���U�$pʍ9@�{L����U ��md�z7y6Ém
�<�1T�25L:]�I�J��U���X�<0�2/�\����dF�Q克.ۦ+"5�^mM�Rl"�騖]l��Z��*��
gn��F�"�WB(����f�U��mX�t��ݚ��{�J����MO�4��~u
`K�Waj��Vcy�IgʒB��J�)�u�aGV�Q55��i�ݝ���KUǭnǵy�$�f�9�J=��ǖ.R%��-�u%<�Z"��R�t]�ܦhZ�R*�:��'%<���(�8�X9XY��7f�n�:a�`��P{�h2bug%��O�W`��t����vC5x��y��]%bƜ�m��ۆ��N+QKxb+r�]%��4�Z����ꌉ�f�)Tx�aun0K��ׅ԰Ke���E,���
�v-'ؘK%�c�P�O�Q��.[��EN�e�Aޏ��պ�&P�wa
�ѕZ�ZM��8� �J�$#to�	hD��b��ո��.�1�]Հ1�E� .�X5�W�q��*��ppV�zy�X�r�u��ތWkK���EP՗XQ��1�sG�+]ՠ�n:����~Y�J�Dc��b�i/��m]�ZZ�XɒQ�3r$�Х����V�F*�j?eb+uD�x=)������"���jÂf�6S�E�-M�wU/i*ԣ���R�G�i^�d�6�m%�	�h=��
Z�,�+NoŚt��a�9���T�k.֥j�DTC.�$��[S�Y���Qdc �][IV=ʶ�I6�W�3RW���ںyP5Wf� c��V�Yb�����T�՚)��1%� �R��8�i��[� +�=�K�EJY��p�D�X�anaiɐV+�Bi*[1F��fn��LX"����A[�>���v��Xu�I��`�+�Yj��X���&,��;r�m����Jj�bb�t1�sNC&b,5�����C���͡5e���7-((K��J��5�`î�1��˭����SD�M�A�	)f�1�+�*��݈��C[	x�(�́L;J�z��͎S1L9�$�r�L�S(㳻L��d�c��w?;��Z�"Ph��:�#2S�0�z�1�:E�bk2�n�͊���Hh�t�KT��e4�sDoF�<���۔���*�̧Gon!w	Ha���	q���ar�d��
��+V�n�Kv]<bʪ��	ke
��R�2����{H�NX̒��󦕵#+v�T3#�6n.����bl��O2��S�kb졮���_�d�6ɬU,П{�Iq�9F�4hY�J���B�4�=�3�L^�Ԫ�y��U�:�m�o��UL�������^�oh/��t�h�Ne��;1�0َ̑�jU�⣱�b;�X�hܰ1�bX�̢~ �Ll0�蚳��4���q�%;�劆{A���
��㬎��p�,�S�CZr]���wX�ٛ��ZػT�Z�ô7iQ�.��z򮓫d�k@��y@D.ުIR��I�E�W��׍�����ȡ^
�{1Uʐ���NVPײt�'ohYu��~L�3?�	�+2V1�j	O$2J�U���g�!KY����]A-�ܢ��6��N�Z�T�.1�vT��Lc����Q��H�K� g�Й�-��ښ.��̴�TH����y�*����)U�|�2�!Z�sU���Ѹͺ�w��bJ�{dT�<��Q�āѷt�{b�`���k�g.��F����7.�ShM�.3���6^@��������
,Պ)�^A��U6�͢�C���0�6�U��wH����z�A�q�mm{J�1��%q��e\�Y*-�h�`n��n�w@�n:�ʴ*J��ݳxkd5�B)J`��ui+�ۭ��nb��Z�+6�2V�n��v��Qˊ���&���V)(�*ɪ��q�Wa��%m��(ݫa�H�)�{J֡j�fҼl�M�;�X��KDB��n;$�-�'&&�YP��M��r9��ͻ�yI�WzW��.�I�`���͸�Vx�C7j0ͭrA��7t�X4�(�
�]bl;��o�dS/E��JU�J9�X�u�#��!7Z��h��fJM�%��Ƶ.���\��4�Cx����`�l�ij�H�b$u�m���9R��W��M����2�XĤ ��PBmR�C�ԫ�����(��n���X.�q5�T������BG�-d��i����F�u�&�E�� ��ʪ�� h$G�%܉�G^e*𑏿�v�t����O��?�ϭ���3'懟��?OF~Z~�P�S���s���<(�����w9�����Uv�+��:����Rw/��W]����k�[i��:)��Ր*�)�kV���eJ��մ�,�N�|�v[��qps�u4�>�݇�9wSW��o�y���]�2�\����q=��}FbJ��Ϋ���[�*8���:la9S��5�m� 6�(os0�@��F;�P������4���s
�w����*�ﲎ��s��9��X���d�ť��"���s9f��]��x��f%�(���ؔyZ:6���q}�b�j�ǩ�]-�0l2�;x���P�5u�{��|�!(�\{8f]l�-\�oN��m��9j�M�W ���ڴ�7�9u�b[����l��av��Ӯ���N�p3���eH�<WXqs�p:ٗ�)*t�A��]/�v{�<zRޣ]2ذ����ޜ��n�2f�s����oz�y�s9K@8a����:uM�WJ���ZeX�ekn�>�C��*ܒ��ݔ��<Z� ���L�z:+����0��B���'�ft���5X��*[\�,�;��@�i��m	������2�W�v��9v�86Bxe�mujԏ3Yi���>��i`5j�9�Fu�$��z�`g���e좗ݛ��a�ժ�Z3D��;���܆[;PX�g�l��Ay�Y��D۠��a(�'���1����R{C:q}r��xK�;eM�uЭ�ڬ�ĠշN�Z6�ΣYc9��,]�'-��πy�D��*��*��wz��Z�tR�h�g�t �j�K�$�|h�]Њ�;��W Ǐ;ԭx��ˏ)��'S^L:�MaΖ�#�4\ж�րQ����;�uP<:���G�����J�y����*{�nIt���-���G��30� �1�	��*:X3s)P�{���x8]�B�`͙�ڽ�c�;ە�ݬ-����[ո��{D�/)��;���)�e�c�=X��ݩ�a�����qeӷ�&���wz�p������n�A��އ�_��QǳA�m����*��xT��D��_Z"�0�{)�o�vwD��5� 3:���˶�|:���I
֮T	�Xb���f�gS���f�3x�q7�G,ͣ�m�������2�Ae��Mp����oi\�g�eN�Ε����n�3F�*�If�c(�����Wm\�+��(s�Q�{۔�|�-E!r��o���ʎṇgEսӎ����R�"��N�Ke�Z]��Z��0)��9Q�\#�!�ת���!�6Bh:OA\XTw�_^:Xy�f���ꂥf�(r4�SQtĚ-p�V8��j�cߌ%�_��r
�1�����c(�0�L`�
���9��]�����8L�;�Y����lh�^*�t�숼�hv$����`^�Ge��R���xUt���u��"��N�Ŝil��b��r��s�HS��c����O��FE�cۺMݰ)[�xH��X����F���B�7GF�wh�I�=o����dR�cOjv��W^.ѷn��*qKwgb}3�ncuEP��i�8VV}�ii�Ʋf�6�J�fF��\�e�݂��j��ܜ��������c�*	�����K=��B񙕤a��x�\��,���q13�q8�L_>���6lJ�7Ol�6y���ze��X�G:shi#[�WR���"t�Z��F1vy��;9�l��֐&N�lھg�ה��ssd(��G)��@Ee>}̨�ٵ������b�#�l�&
9�Y��Z�;(c��:����hlS8q�grZ�K�bF�Q��i�5Y�>\�6��d{+�GV#�����]W�ZÌM�+EL�rdy�9xd�r�W;t�n�c�hWj����5���a���W/7��$t��4Nu�焷2���J���u��Mv�����>5�A��o�+���%�=u̳ �&�omna��2:����Vss�����n��A�P: ��\6����EVj�vԩ(�ҧz$�*���lwr�H�f�ӘgIkه�#���y�wf+|����_.�8`�>,R��x�۷��\쐺�z\��1ֶ,���ްe��N�u@KR�|^-K{��Ls0��]��n���A�t�U
�����}� �)�J����G��^ec�P�4��M
� �u��Z�Bn�G]ĸ @�A�YK�qWY��U�o����A�Jm։��Ҿk�s�y��4w ����R;z���f�YA퀦�W�u�� 9w��=y�.2����5s��њ	�SATU�K��PH
u��J�)ΤȒ��%�T��,�.�6�%3�f
��4k�-	�>�ud�]�Ѫ͌/�E�+�KVV����C��Z��UԨw�o�Y� D���ڍ3��
VHS�U���NGfeӹ�,W5��F�b�۟tam��ECr�V=Ŋ�����u�)К6��htԴWf�G�Հq@K���d��m��c�5�Єe����Tޘ+����C��/����3�_4�)==}��:��p�{vݴ��12ِ�PI[�oq�,�+Q��	�������3�<��g[�a�<��P}�%�
�<�(+U������yګs���ۄhӹ1r�^[<���lv {r%���Zg쓊�C���c����`�X�Z;��M���Η�qE;y��{ˉ��[Q�d����ߥ�K�M�E��������^�ϥ��.Orw9�m�Z�S��Jq��S��C:�X8u�	Y�6�%�Q���K"<4:���(.|�^Dr޽̘��&s5�g3���5�**�cnn��ݍ]eL�-M�%b�K�ʹU�В�b����oMq�h#C^f�R�6`��;���g'�ō�e���M��o&ju��Goo9�TQѻ6�,��rb	��M@R�f�{׼7�V�*��Q
:71�9���\���ir7�ƌ�۔Hʷ��yE��9r;s�r�����oU��w��TK�K[���w�kJ�f�s$�r�.�U�Mŋ4�}ܢ��cs, ��$A��)WZ��S��(���Z{���oW\�B`-��F�V�@�ڎ��9���G��{m�s����-q�T�9��rweE�ݪ��_i�v]`i^�ٖ�q��t(�����sPϱ�����H�=�R���Y����B�P���-J!Aөf�M��V�;ܤVN\]^�ˏ�!�e.o7�]��YhR�����jW3{�Fɕ� �{�^,�@:`���x4ٳ��+�����z��Ov^rv�.A�%��ٹ\�����p켨c�r��k5�8ݳ��WU��Lɹ3j�p�U�[���+��l���ЬnV�E�3��w
S�(T�ڍX�qs*rw{�5L�Gc�Y5f ]#�B�_oʔ)c����i�_V-���WM�,胓���RXS�����/(˘�c)�dwn6!k�I��1����n�#|S}��!���۬������3N��I|_m�f�j��|��7q�=���+r�`����b�t(V��훽����_CX1�����k�J��vb;�����_ܙwr�*�gMdi�7���n���FC�r��Y�i�2���;d�׿][V-K��S������mfj"%c�2u�}Wz��Ա+���C��#���7;pL�m�f��h���a��w%J���D�=�z�:v��m���wGZ ѢA*U�[�2ݫ�Z���"J��T����фFa���2{� �ݹ]G�a���4����X$����
���;LK�ҳ��}�h��`�N,�G��7��Z��u�8����5�@�í+r��ۓC�ϭ�����Gt�M��)(���_�+�|���;�n�7׃y�w$㉼ɔD��w-�	��1J:��]���2�Tڽ�%���[3iG<���r�Z�����bs��`Yח�S�2�s����(���:�=-��O^�B��^T{wQ���؋�CE&��;b�b��:(�Z�g��9�@f�h�x���v�Qx,���+F�,[�/�u4�v���q�u=i=�u*>�=��p�F7�R��i�B��|vX�xUX(��$���,���ȭH��̼t7u�������5��E軺-�&���]�2K�V�UԊ4j�������J9�哩�;�{x�\Ɩ�9fsh+���4�H�<n�w��;X�*�m�V�C���b7@̡���96V�gS\�����b4w+�mK���Le�6tVwa�uò�Ѹ��fԊ�\&��a������� nƤn �z�]ʂ�;��\�c�C�X]uky���z������x��U�O��Df��b��@���}��Nė^R�0�]7�K��ٖ�e��f�yC�O �[Y]*��x�E�k��u�Q��kM��e3ʹ��k��Б�[��<o 2�co�`�I�3��o��&��`��;WX���_epi�ϐ���+�	E��q `��]�p�|&�����)��a���27CQXr���mmHv���'81��h*�ӤQR�����q�pň ��:Br�9�0;U��s��u�ꙉ�<C�"X\'|-	��k���� �CS6�k{Q;�"��Yger+��۽�"��R�5N��o_Qm^�&���ws`��L�оC�
o+M�sz��J�}0d��$��|s5RK(�:5���k�%�׃�����%$��R�WAeJ_,��l�Mjs�\���݂���s�+T�P�ؑ�Q^;�x�N�X�h������
M��!�v�{c��;����q�@塰k�`�CS��8Y�����a36�Iu��q�;;�.�`pZJ��߸��=�K2�QF�.�X֝u8��NX���'[�Z�!�2�6w{cWw[[�B�9���Gv\����b���f��fd�J�l�;VB�Z�,�WW��
pKMQ�/�Ո$�|W#�L^j���ҿ�*qs(]r�A�,�i��K� 뺹�q
��-���7T�Dp��+&]J��]�T�wo�<*�R�TO.�
�vM�-�zQ��V��Eۘ5�N[D��K�/E�a#Pd���>�N:h�2蛹��	:�*�;;2I��$�vմ��W�kN��sJ�E�^ ���*%�ɤg�>�m8oX�W9��3�"���=��7T9p�, �����q����+3�1A�t�eh�wHV
=������#	�Ϋ[͛�����[y��M/�U�:_��os=����1��lis�ܚU`�\�ލd�����j�-�J��]�{���=՜0	RϦ����g�K�塼:+���+=Ę5��z�|K�i��WK��j�
��_Sz��;ú�%�Y��$��bΓZ���{ �f���)�:_u��V�ɼ���Jm�KLb�������^I�"g�bpJ��W�pL��|�g��T"���.碌/�ηwǰS�99D�ܲ+sN�y��ƨu�P$�Z�\�O\��e�F��5���4��i�G��ğ/x-p�3��� % F�q�e�ֺ�ʜ�<�6C��u	B��dES�v��
	���ۻ�ȸp�-0�x��G�x�V�^=�*ɋ]�w�T�$qZ8����
ԫ6�'��O���@�s4d;f�[���z�VhX��Sj�6��^�W�ظJ�9�hkj���J���\��f���ԍ%��V�^���:.�n�ݴ5�iф:����	�*�%\��: ����Y`͉�����|v�Gȵu�S�D��"�����w6�?	�R�t���7no>���lY��Mgk2vya�{�۷��ԋ�gEf�v8vM�O7%�T���x��4�AZ��C�^�i�ĭ��,����C�����w5a�\Zܒ�����(
r���UM�Y��ё���ӗ�z�%t��Pe -�D>ŝPF��<�&L��f�aj�w��{���ɵ+oECl���li�����Sfw!OJ#94����n��ͪSaH,�1���{xY�]�'���(Eku�qVkI4�̴iHx��9"r����VF�iX� Wrts�1�u��ɽM�K:�=z�Cm������Ȇ��A�9r����ߘh�oX,�}�B�nL���'mm.Ck�ǯ��u'ϪC�����:���}]Fqs	��bg3��u���l=%�ѽ�M�v�S��K��x�@�f�(K������X��էk����̙��bG�B����#���uZᷨ�v�����'o/�����>V���aW9���yw1���ܛ��`�Jg*���|�7�_J�I���#�<ʙ���ӻ�ww$���v��h��m�A(��O	�W5S�o�pyΟ^g^l�W9���8q��g�sx�w0D��v��ya�ק�|[>Fs�M�a�C�$�7s��"``KsBގطQ�=�I�j*�\a�;L��ZV��H�Xk�M�8[��gZ�5�3RŎ�-=V�}�\��,fvpN_oA�W��e��SF�)s�<��+R�Y,o-X/��%�9Ʊo.R�5�yoJ\vq����U��1�M ��9tkIT,� )jc��.�6�Z��4䠶�N,���'6׎����υ�4��N1��JEN̻ʺ�J��Y��Vv�δc�i�g�������F�AK,0��ys\��X�γ\�d�cu��Uu٥C�y�w0�����A���K�ȸ��2G2�$�����^���'L{�����?2�O�f a�6_;����@ M����I��o��*�!����  f��c��!Y��^六3�Ɋ�ݯ�����1橝P�R]�1)��j��6���NboQ����w TzU�J!��������}\zT+s4Y��7�n���::��}�M�v/3�ح�zxs8b�6>o�Sk�n��u��E�+��u%�W%� "�,{t��x�	�����Q�	X�9nVh��+��{
����𯌲k�*c��:)�/���g����m��t������y���qe;4&,@�ϲ�/����ݣ�r����Yx�+5�U�vbpp9�u:ݽ���9j/���4�*H�K��j�E����
H����Q8]u%`])v��|l�@���s��}wْNu��8�f��J	:��C��ʁ�b�e�X6󹭼�/U;M=�������X;ũpK��f������U��:�P��r��б��l�}��)��M��K;�n��(��%�Ou��r�YvU��K���ec@uA}B���R���eu���<�c�++�O�ՉA�P�>4gb;�.-gs�\�2Ê�N޺��ETg�ً���bf��;s�uL=�R?����*�9ڬWub�NC���0�7:�sW�o�SYD�@�kV�	a�}+r�Ì� \���aQ=3�,�Ùє������Y����il9����+���
B�b詩��oY�q&6�C������r.'�]�VT1Zǜ�zV�@�j�|��ܼ�b�V�u� --�^�F9ܻ�|a�-%��]d`ۇ�`�շ+gw5EZ#��F�w��@���*��TB�������wkT��0���j�M���x"[ٵ��YGE5Aλ�s��
C�ٔM��.J�xeq�	�ջ	h-�D�[4<�,� xt�grF�BԪ�l�oM3�O�ٻ��n�e�����nJ�b������@1�.VC5%�on<[B-Tz y�V�lq ��+��c�l�b�u��$��`="�C�4���,� �,�W�sQ���27Q"��L�ӗM#�DTt[��������H$6�·.j����
�C2���X�6�v���M����wjU�@��#��-_���e,�6q/�U��k�-�5�4���{]L���U6�P*ݬ���\:���\6�`ڹ�kr�j{ZVǻk�5�
v�Uo/�Z��9TuVI����v�p�_R�edL��J�)�횪H.���mJ���=��+���Er�S��gk�5�Pl��q�t*��e�﫯 bbY�魕S�:T�P���)��&�q����'N�2ⵅTqSĐ���n(/�-*⭙Kr��� �;(T�y@`<���&p��q����ɭZM��#�f�L�D^ϡ#�`S�K��Hs�7_�*�c��{6׺�z�G^�Nn�i�Ĭ9��wG ��:�׬�eW]��R�*�u �L�mH+���5Y�,]f��!��O����Jv'r<]�_H;)�ڔ>�\.�MWq���E<��lV�2g�}�"�9���0���хV�vH@1�mLWSEwf��`��
���W\�_S�Lӱo8���H�/$oC�[Nޣ��OYF��\�OeԌ.��ܨ��w����jn֖kb\����M_:V�7{�1�5P��R��;m͓l�垬�b��	�Y�j�gM@/��ܦ��e��6u�+#�������5,8�G�v>L���i���=ZQidu��N���˶6`�:��f�(�[xp`�Wt�(%��/�ST4���[���5��Z�%�.�gk�^��릶��lg$�v�F`�BWX���:݆a�q6g��G}�N�b�6;GU@2��l��Y��fj����w�g���5���v�\�mU�ҙD������	>����wʷ7�{���[u,Ŵ^��(�7*L%��԰va���v$&�i�wb�a.��pԠ���X��p��h�e�ݙ�#��u01������U�Y��Å��7(����^/�R�g����Hf)�D_^tyVc���y|� r�(����G�|��GO��Y�k}V�@�Ƅ��ڱfk��93���Mk2������mω�%N+|�9ԡ9%Y:E��:hԔ1vR*���{��ӹ��_<&�g�f�7|lH��OVb���m����W�u}u:b�_^C��1��ڹ���uW��mt�����Sܮ;Q2�s��i��n�J�����H�k;4G��H-��;o�ٚJ��0j�
赪�dt���m�Eӷ!�9�N��v7ʎ��;�;oB5�!ݠ�ڻ7�0�]�ltH��Ѷ�m�末��-Y�ɀ(aT>�یs�e��m�=\�¥,�P>��(D'+�uo��7��HpS)#KtX�)n:�T���..���,�v��iT��8A�/��2GI4�o��r���-eq�}ٲh��g^uL�h�I���[8�t�ȳ��9P�R�ee�d�O������k��T��ԑ6>��T�we�b�1�%���G��Zx��建e�YG���!At�X�Q��7��R3�Y��rv��r�8�U��Ky�t=#�mi�,��ו1��.��/3+k`�Jn)i����A*�N�;�룋E��ov�P��ԾCH����p�f�儶B����e"[�T2�Py�Ni�P��Ϩ>�Ι�Y�{]
�ǎ�+�Ү$��q�a|rf�pTFMu�uwVs?#ug1���������:-O����Գ�B�a=��7�uu��ι���%��_4:��_h�t�M�/jޜ��qw�B�M���:v`S;_\�6�C\U��k)uήu��ɝyĞ�adh��x<�C��@40�*�>�с�Q����8t�Ozs���+�>=3\�[[v����j�Dz�������4�xH�&B7�B��HhgL��8�M�{��
�-�g�k4K\����r��u������H��zw��Y��JXm�+{wz���7���$��h��MT�r�{�*�gqΧ\	t7^�V:�sZ��s��j@�K�J뮮[<؈���q����M�����Szs���s��PZ��|X�c7SL&+7g
+l��2��%�'����A���u�1Y=@zH�{@6��h�P�;(��J�-;j�,��:0�'������t���%����$���u��d�ػ��WB��]ݷm�)������sYrr��B�-]Ð����m�XtX(]���-�YQ;.��f�:�R嶴�6�2R��x�Kw��}��6�q����ɫNivt�:�5
:w2��2�h�(kV=�K��EW_=�U��}�u%.�R�Cz��D�Շ�m���t���U�����h|�!�vӻ>cA���jޭr]��[�GΎަ��u�J��A��L��+\V��t�Y*����[ς����h|i�	mǔUN7Ζ�Z� �V+[B��{&�n-�� ����vs���+Y[��{G���z�ڼ�n�h�X����m�![8�w|�K.^r�&l����R�M�\��`�J�������h];t:��G����/ruB{n�T4*��#���ȹ��c�6V
�
U+�=��اˋm���V��u,\��	z+4��ݸ�}�U���v�Sżd�d��)�j�SC7�f�:��j�ȉ)�;�,�B̈�Хn�Z��&u����O�g5q��YY�O.�&駴
�nf��u���۹у���]W���r�7�Dv/��{��vP��� 3Oz� ���D]i}}ҟt�iX�dCI`����R�M���v�!V�m��+Op�f�������:}�����;Qx�r�s���z��	��w(�{��ŀ�sv�k�1f�A�S�V�+`'%N
�K�)��g:��7(��)Z{krmY��+�WYFb��&[]N�ӵ�՞�#�����t�������Wnc����/�����6�97	�$4h�]�{qf&���J�	7}�`hu�-<�[$��lh��Y��FZ��S��lm�l=u�A�ل��T��]F�%����v�6�ڜt��,!�j>CEm�K�'��B�r��Z̇-7H �Z򬗷���s��E�Yn��)��� �;�"ob��x�m�s�_W��Sc�Č�Yc���̵�2������W����ʏn�5�Ӳ��&�
����س7u�d:q����ŋԲ�[�i�j�s��=[��4�Քg��qc�S���u��^�5۳kL��l�n���b�����@2O�����h������vԶ��w �/������>x��5a[\:u��,	L�WW7�cE�������������p ��a�z]L�WZ�O��SK�-��6k�Fb�J�{�X�<EYH�m?�S*��� d���:�b�\�<��)tn4!V�WQ���|���n����LJ���Y�t�����;�sP"��Xv[��Ui8��)&v����P�}l�k|���Y���n��d��y�F�00������wo0�S���㬗�,�W�]�;~&�Pr��s��p��vW�{1���`�sWR��.�������F���@lA��l�+��w�qyb����F�gig��'��D��� �%]E���ͧ�kη+[�K}A*O�F�櫂$)4� �ƕe�;]4��EgZ�9���;<�۸��X���J���\Y��t�U���؆LY�<ج3-��Ꙕ��vus �r���1,Mr�̕X*�Yy)�x���6��)fa�y��F�q�D����K���ܕ�;ڽ�|VLܨ��[{(X)�Z.Vv�z�Q���ALU�uaTo&�"Ļ-��5c�ۗx��]��uïb��0�h�؛��b{��!��.v��;l�t��I��V����P������B�y�v�p�!\Uݴ��TY%�C�J�ڵ\��_
�Y�O���ܧYn}z��� ����-���.����0k34�%���v^�������Z%f�]���j����(b������2��V���d���_��nDEJѬ����4f���2MD]\U�k��nA�,={������3�uJ�;6��]f:�b3���3�<hm�y�j� ��l��u+-��#�rf��=��ë��'���愂�t�j]�L��G���Y!�%�ȸD���/n�%��6�KwB/k�U�s�����V�6��r�Wy;V�P�r�7*] ���Eʱ�R{��eAL�WLM��ൣ�ή�5�u���,���7s��bc���>��C¬�m-�&�Ub��٠1Fdӻjcj�IzQ�<���ę�/YE�a'B|���d�Y,#K�����e����s���}o)c,�X@Rm�ap���V���+;ޚ�qR���H%sGIn�'�m�����ޗ+,z�nQ�����"a��zQ<�nw�v9'=vŁ��k��`��}�`7Q	��8H�����w�iE���S�C6�RT]-�K��e��7�SW�Lk+
混�[�鉋y�zu��T|eC/Z�.��-ނ��2����ـ\���%������t��Ƣ�|Ƌ��j�X!��hk-`{nnZ��+vͅ1S3*����;�� ђ*��3$��k�� �
nwt���r���*���Q1	��n�Z#��93ݘ@��Y�t�R���=2��7�;��V��#1��{�\$��(f�I�K:u�� \�FP�����)mCv�+��W��E����P�y͛��Q�杇���ţ��\k��cn�ZC�Ι�}���;NZ��i�{�S�}'VfQƜn[�c.�9#�&��0��{˾�ia,��X�B�J����wJӹs1ɼ���h^=��;�o�(��.M�ڨ����{T�(}%��u��]E�7�I8+5��ޤ�PK�9]����K���e�6���P��b(�{��Ιw���B�[ƶ�����ܛ���_(S9G|��R�$�tm�(F��i���#������d�YyP\�ti$V-"I�N���s�Ѳ��7s]���T�݉8�[��S6��V��"�ari�i�t0|&�:���ҙJ�	�x��N�7Smh3T.�{�J\�굕�N�s��ڹnq*TiʛR)Ŏ�m�5�4
�L�u�s%Y��Ê�/�S��5�I�����9k�]�PICy��-�n�&�V��e���-��ڴ11O�E̼�Lr���v�gh3j.S�!E,f���D5�-���Xs��S���ʙ
�f)r���[0�j�>�Ļ��tWL�q�
��8�xgk4�Fs{)_r�ֺ�m�yFL��0d�5�6�sdO��S�Y����`i���N�+;���he�����S����R _����ڈu�gW6l
��U���Z�_�ש��v�+��k�e+U�[v���u���	��v��#]W�^��܌�Wu���Na폫�u|ss�@$�}�:>ښX < ��q��f�7�	lCm�i#��F�G�a���i�/z��M��7�r�929v�娫��2X�v���sC��A��Y�O+H]!ׂ)�s��v!�EK�V�`��U��$O-�}-g=���)� A��1��A���
}0�)Ct����Ž䀮�89e𫧜I[w>F35Qv�9�f��	n����Xh 9:N0w�k��]x�i;BEL������Y�;<�٭�%�kReƙ6�s�	��5��+{$#d`�:ABw3�����.vv�j�?)?I$�$$db$���M�09��?���<$�`��j�3����m�ʇ�rD��3=����Gt�p�Wl$���
���`��\l�$c���N�S���k�">�;x����z[�ӓ�]�׹wN�]��'1�/r���5����tA��t�O��VӨ��B���y���jP\��	���뛅�쑋�V�*��W/�<t�>��ik���f�>Ԋ�R�
mo����]�Koq��V�Kt�7�I�TB͚nցX�i^�}.P=D5}p�3(�4�N�vR��O�Gy]e��/GF����S�����_2Ҽ�^`LX�����%�y(���x^WK���u%�ĵi*q�D��OTf��,�]�5-���-ӣL_S�N}m0�L��GJW�̮��;4	��^�K��A�=��7.�:�]i3�M0O]����i\���]Y+o��-pB�vC{�e+�l=y�b��PL��V�/��R�����%��jR�]B������������?d��Ř�ǤF&w�씠N,E`ڋ6��BQ_�qm:OF����0oX�e���ݸ9�f<I�vr���@�'�,��W����
c]�n����:�:]�	цc�x���FK��}Xt\�U��������a+�=�Ֆo�4zoby�F�����K� 릊�%�˻����9]��2t�sT]�^��1�m{�⤒�lN��#'�).]x�J��|}x_mI�|��(��-m�V���M�0��EE�P�´m**�DK��*�6�m�ne�PV)�E�KD����+UkUQZ�m�5̨���孰�UEX���\b�r%Q���\��6�n\�[���ä�ꑴe����i`�is.E�3iZan52�Q��V(�cU*V�e�hZ�PnSUf8�f\2e�m�-.ZZ�Dr��1Tk
��1��b�mV�#z0�",\��"�[3.R����̭�s�e*֠�[jR����̨����J�b̴V�E�ˆd�*�0��iqi�3	�3%r��(�[h��"��QDVト�m��[�.88+���R㌘�(ƴ�jփl���n��30�-���LJ�*���h�̵�%,r��6�[ie�6&	U���X)��&#���EJ��9U����X�5kVѴaZ���0Qr�Fe�i'a�wN� ;	}��D��ڂg���峱1k/���G��������;,o�^*�֮2��ܙ0�8z��-�K���ջϤ-�tL]99ׇd��_߯��O�e��yzBWs�Z�c4� �����`�޲6�5�9�q-X�^� O3����+.T:�8�:�Ø�b��d䦸
��Ew��YJ�f��Bga�Sz֪�C�j�����5.YWK���r +��HW2xW�����M��f�]�*�#�`����)��
�u;:�<j�[m7�Q-�X��!�����a����f�d�`�����i�h����ݻ�7�+q��p��Q�N1º��WHV7��H�]2%��0<��'�
��V�/Я�..^I�{�zÉ�P!��l�IV`�����5.wU�V�1��ap`O<v��Z�G��U��ҙ��q�hܡ�cV�S��8���4���=)	Ȏ���!2f5m5"=n����RܺceLu�3����=�
~��6���V�Ch�͹VPr�eK�E��繘Z"��;� �t��0�iB��ڮ�ĝ�qǎ;T�+��e,��8����v����*T��|�c%ꫜ�+����u�n�:7������k$�i��.-����Y�������v<�sU^&�W6!*_l��ի,�oj◔�~uÃ1�ӳ�X��dLi��'���:�a���A�oy����]�D��Ά�rn��o>�k���L�V�vX]C%�N9�p����dI��ՇE���_�f=�Tt��G �1���.ؗ&|�9t����Z��h�؇��}q
�@�:8�������
7���"��b�K��#N,�`"�	{���*Zq�)��F�H�`u	^����R����,��	��8���\��T"�ւ�����v��p:�`�Bf"DMD1�8��ԥ����&��N�M����4r��q�����ΎN��;ܠ�u���%ח2á\�P�^�~s�~�B&�wަ{HXO��;)U9�|U7��ԪP�OdJ�cg%�tM�ӝ���y	�#x�WU.�2�&f`Z�����d��[�B����IN��Y,����s
q��z4�;�5�+7��OCT�O��.mdИSE���@�\\ދ�r�P@��w��I�TgF��R�=�1Ov�D�*l �}�߄��>�1c�|�3�w���%g��o`g4�R�å�H�81E3
$�u�h��;d���0>X�C��~����A݂�f�՗5��E�iWV�1�gO�^�t|8�M��h)�nRI���'&s���"°��ҧ��g3�p�y���܏���ٜ>)����D���µ��&4:]��J;�cYX��֖��0�F�M3S�G�t7��3��1vo5c#e�q�':�e�\�f���f�¶Fpl^��5ƞY���ִ.���9�8���/~��M��:v�c�8ܸγ��S�;7Z�/r�0l1�y	|���7�e�9rU&[�,`�S1���)�=����aƚR�S#%�0�3w�^�[���ٖ�\!�wna85�r}�4��И��%��|���z�=�]B�j�|��뒜�ڃPa)�Gf橪�c�r��"�dCc:�Lt�4�
��$�z?0=��y�Q�ws��R��q�)*ZϛpoȾ��Vn"1j�tT�6
�$t�p��gU�'BL�m�mv/h�C�H��ɡ�qb�A��񼩣.���:��Zb�nj+�I�5V�.�9wYv*n�/F@x\�g���+�3����¡��N쮊�r+3m+�MKt9w�t��~��**91�)��H����L��a���Vn��y��t͛����Q�˝}fg��
���Z;Y�]��iu�k!�RW`f�BE�NU�O�9"�>�K�Ԝ�
u��z���G���-.]8���\1m'a�*T��ش/OL��NAifz�Ԗ�pY�˺�_]�bo&=�6qS��*��Z �,g+���`Z�ˏ׋'�](Q{Ң&Ci�wU���rI�Jxw����B:P?%JƜ�.L��qNO��	�n� �)��f����������cj�a����5U������g�6�2-T-�┘W@��c=N�b���KO��X$�bo;{Qh�ҴR�x�.oy� �\��J���LdI�VL+� {(yqX�]Υ�?b�s���M9,�^e)����y��|���*���r��ps�чz*yd�L�7����X�qո�F3o��LZF�&:A\\MI�MX��.V��{!��+n�(����y���ԵmK4��c^gZyE��ͻ�:G�F�3�dKp:Uj��f�A�����J˴UX�];�2r]V�|})-�'ԗ%�<�};dq9u�6�V��A� ��{	EjB
:��� �0�=�}{Q��5c�])+�R债����E�]�X�^��k���	{��L�ƚR�f�����X�|a�Y{�n��:A���f���Ę�Y�vC�etIP9;�QM�~z\�T����l���(wNz⭝4�t��|[���04k+sB��N^Ů����f�h�!��Ƕ�gf��z.�̵[ x��R�X�l�.(Jg��n�ȡ�:
n��,oV��OG:�;\oP6Ty՝ͺî٩��\���,x�<�8Mj�N��Ե�	�pj���O�&����𤕾굛;.aPbD'�%���XR�>����%�Q���Z{Fj�h
��s������3�^ni��Ȱ��:+�+x��zJGy�;X`���@)>͔���
��i���I�h�SJ)ʸvB%z��#�0tx
���])w��*��W糩�%�*�Oގ���1^�7�V�<�q�攪&Ҡ�>��LTA��v�Pc;V�&q��I�3mOX��� ���	�ў�N�T���dD�%BP(��u��3������n�N*#�i���B4�w���q�26%˘�b��d��@w�.��IŎBW���Œ�1���)�7A]^o�~Õ~�E	��,��S���2�cV�����d��B�.�-~���C���uQy�8o;�!m�ߥ��D�2��&A�Z��R�9H:���0ԩ1�lC��n���s���='M��~�8�.�c�쨗�(�ݣQ����յ9s���j��՞��`;�UA�-�{9}X�I��e�������s:K�\�R�\7	�5�����.�#���Ѭ�M�����'P.Q+J�b�~��f�v.��>��S�Ϛ��U�}�f;�B��H�������7oU�YH�M,��&UČ�$��Euvt����B�fDy��U����>~��%�Ib���,C��V-�$>����v\��|z/�w������6v�����;�v�e�/[un����{/'E��͓z���NoJeS9��P��
���#��n��;I1���ˤ8Y5�eq�PT
�n�%%jf>w�̇f�D̜���k\>�0n�8�9�������F �iGTNqCs�%��Ⱦ&s@ٖ*w�����{p�_Wgc$(�֌hk����1�0��vut4g��pY�޹��ԓGv�3;J�jzTT�fr]��gFT�I�R̝�(1or�[�Ĵ�j���Y��H�Ba��ee)fmq��u�kH�e8�z
A��ߥ��Xy5zˬ=��Q3�+�r{�/*��L?+���q���X[�YԚ����gu�b�:H�7�4ᛚ~u� 'jX8��^qR��ͥ�:/�l��8ϯ���&F� 8�y��+�y�2;J��D�x�����9Ϲ맼�n�}��c	�z�L�9&T�/u��4�u�3;3��){��s���zT��Nutu���O�k��<��'�����Y��R�'mٓȾ��.I����W�Y"��U<W��kW�lt{�nr�2vh���{�Y˕�U���T�ʸ�x�.2V�ú���ss22:�6kv�XVR�ݮ~�bik�\ڂ�-��<��O�����8V5yv����s��|��iL�}L��V>���c�>��l�fW��vz����ng'�k�R��3]�G���|\_��1͝ZԻ�̷y6}"���{;����@��"���h�z�����Jgʙ���8�tp�s�쪻�֟.}�r�u�H��+'
���_Br�,˛}�,��v�N�)�֞��K.y�=�,yV�\ͮ=k�S�6��ݙ�2|����
^d>��]s|�%u��>(�`��o u,��1Tvn^�(:z�0b��;sVc�}a΄�tU3��c�i�,�3:� ��%�4��yC<),>'��^n�;�&��'}S1�]î���L�[(�x-ysI�wgN��'%M�@r�9%���v�4�R���v+c��2rm�r�V`���qCv�W�,�I��q�a��U:�9B�ù��t�A�-�#a�I� o�� �k/ҭ<�k��Y�VS�]\��i�Ø/a�5m�<XytnTTD��9a�*�O/��������3e�o{��bE�<��śz_*�9,¹�����L�V[���S5/:n���<����u�{�\rgj۪n�W0pЎ�S��ߎuܯL�݁Iy/K���Nv)�}���Z�u�~nk!+�aTq�O\�tѫn��28��Q�4���Y����G6��](-�doy_fq��ҷ� �jNM�.7����l�[���K�
���d��}zi&l}/��9�m��SFm+˥���Ӕ�=�����A��}�#Ra��ר�<P;.;��0�����(���K^���c�g��#�t�~Bѻ���s&_w�:K��s�5M������SUz4�"A"&�Hk���J��r�rk=�R����S��0�<����*�5�yK���b�<��tq޶�qy�)JRsq������@#3s�] ���Z�ǒ�fr�洜W�72�tj�!�/v��՚�J~Ru�#\�}OW%~������ݛ�"�3�Q�^����^j��|R*���6����p��U}4�fVM��rP%�4	��N��\ë��}��F�ʦ_K��Cor�3 ˳�
�z�����@rYR�Y譎rz��3�O��yp�^�"�|c6UQ��FrH�N��G.�q.o��f �b)�W�%'7��Yo_J��Z���fbv�RR�����e׶�jr\TN�`F��|9)8�=��o���$��n�*7H{�1g�	5��}�m����*�ޕ����W7�t�L�]�[8��Uk�j/��Ŧ����Oj\�.B�v�w���/��ĊO{��5��$��3f9�{M�Wy��f��	OI��$]\9�H�њ���eP�qk�1q�;�tZ�u�۬���7���2����u�NFO_l��cg�N���!�9�h��f��Q��΢��qt��_��/��6ih�-G����sn��,sȒ������֧���l��Pw�GR�-L��޳LL,�s�����oxK���	������oQ�\\�gN��':�MrS/.nhr�4��,��JQ9�Nڹt��=�1@u�1�9�U5j�y�����n�+���e?v|ag�9<K��-j��9Ŏ'�H��Vj���ýq�6V����{瞘�Kq�����Y����r�P^f�Ƶ󃛻����+ݏ��Y;�yXq��G�x�w�,��z����ÅY���U.}zz/ڵ��4�?u���$�NJ���^mF����K������ŗ�9PV���ni�y����x�gV�˩&v6q����]�����^)���'*4�U3���~��F���.W��M1�gy�Y�P�y��SOd�Qp�_BRajeS����Rp��V��o�Nw��1�ז�U�h��F �iGTNqCs��j�q���@E	OwZ�������jv�%Ezu�zΑ[*�
<X��ooÅ��x���
�k�_�K^`iQ�j���a��M5�]�V���{��EU{�4�:�k��Y�� ۵�H��Ν
�Ρ��NvE!�J��ә�Ej�}�p�����vqVd�|%cu�RU�����r����p'�F�P�K�gn\*Iˍ����
��Q�'���4h�i@rN(5b�t`:Ҭ�gS�{���9�8#��W9�lԑ�i����=�6ѕ|���ۃr#��9,iri2K�{ת)]ҳ:�٣��v(+-_#��oh�}8ô��^S����%ث��q�[Z�V_}B)Ժ-N:[�/$i* ӍCj��Jĳ�f�TlK1a{���Dݼ�4�2�g5���Y�n��>?-슬˒S��3�s�̗զ�A�
�VFC�ϩ�ře�,}�u
���-R_fV`��wq��H�l�8�.��,jIP����'\�ʲ
Q�:���:���+ٽP�\,���s�`�l7ǹ�Gq1W� I�S�ɼmrC%�Җ�`Yv��R�Mb�Y��q_]˖�*�@�W;� �z�l|5���c,&�`p[�wpJp|+V 6�������Xv�|��x��0]��`����\Y�nݧ�3wYӤ�\WW|�L΁]�J�%��:�9�<4X��0��0]�Y��T�����!��k��vW��W[����6�l�ʳAݛθ����5Ү_}GR�jv�b�
��Q���q�u�{���ͤI�h0G]k;���u^�c��@Q�˓\���U�<O9N<e���S��}���oZ��m�Wԯ�$�$��ŷ�& ѵ�J�7��!��[�e���;Ӌ�y��T!��n6�봓}3�2[.ݸ�8RM=���c���M#�=E���I�N�]m.W�s���tg����&=٦ʨ���E9}x�\h����-���]�l��9����@!)�b2�Қ0:X U�1�[c��<̉u�X��P&�e:�����ٰ��yB�-V�˨�U��6x��"�_T�CR�擄1^;�E<&�<�`�#K����7]��Z[5�]��(uu�V�m���C[*ܜk 5��J}�B��'w���`=:��:�8�S�3K6n�Ⱥr�p�oy
@Xc�a�E����w�|;����"��/;7r/�	T�;go[��A����ሒ(�kq��g�h�ᚕ��M ��3k�ԡkT�^�״�膀�TM��r��55�p��CUb�@
�;�qĪ�-�oi���ggMw�;��j��:�����M�Y8��ά�k��h�.��G�M��u�4Yc����u4xus�0h��+k��hyGB��I�SB���{J�us�J�:��f��Xʻ�m�|�|�\�:�!顉rD]LX���+7�t��Wl�뷏��ݟ��J<�8I�~}O���Y�GN��4��9ɶ�Ηp�_s�K�7�7%�{�s�<��u}����l��2�,S�jX�@�\�E�ʸآ� �E1���EeȸdU�p̷EG)D[j�nch.f[���TL�0��c���\mT�[Q����- �PQr���b��\��c�b�[X(en01c�-kQ1*Q��R��lG.$̦8�3���V�s.E[rܣjT��*�)je̊X��s1�n&E%J¢�-l��Y�\�s0B�1�K�R����\�3���QUJ��*[I���[-�aS̵�VЬ�Z�ҔjV��1`�f5Aeh�JP��V���V��Ƹ�c+[ekF,ĸ��*,T(��2˖ň�YB�J1Fҥ`�l�hR�PYVҤ1
�J�U(�lR""�#P�V70�q�,QG,��TT�Z��m��"ZX��1�Q�EX�VVѢ��R���ܢ�����#���b�J�,Z�"-©�j�s;��w��iAf�暉y�3$4&��p��i�y]ٙ�˷]:v�Y2R��c�/&wJF��YZ�͝ؤj�u�K�NRz�sO�������?�-v�H��ԓEk����ҩڞ���-T�nR$b��p����x�%����Z}���{�m|�w.��a	,��}�n��[�8s\(��9}�凐n�ן�Y�N�s�^��l�Lu�✷�l}-%�q��9���~�*j.�[�XF��ԚA���]ɇܩOK{��.Z*�m�?wmDq�H̏%=4�5��;�s��C�2cw/;Y�KbrL�A�^�y��w,���چ�y��>	��W�J�E����@V�U���]-S�㻄�rn��*�q��)F:�э�r��F)�Ж!�Z��U+�M�7{{��]����}�
���|�l�G<��L�ͭν�PEҌW�h�o�r7L]����zT\jֹ�V�T7�f�1�d����䦚!w,}���ŕ�]}�Wд�Ǜ:��菻��q��/�f��u�q5�P�i.���������(\	e��K%(wWs��5�I��+�1m~��h�>�<s^���^^z���ޮC�n���kh�˵��8��U�Rw�ؾ��I�=�	\s7��i�E�']�&���iw4���n����V/�DeXF�i���Y5��g����ҞD5'j�+�:k>�DsT���j9�p�w�?����PTWCq�tb���ɉ��i��I�Q�7��2�y��m�]g�ˮ٤~;@~|�4w����v���a�W����B�|�8Zmb��!�3��χ�NBT���w犘H�| �N F)"6�K�2���Y<��q~����p���V�9��z�%C�OGI�����oG5��<ȍqK7���K�EVd��eVU�|}��օK�a�v�C�i(�Gx��)������o&0|N\�Q�;��b�a���⊮��]�{.����tT!}�A���/�e���᩺M�����qM�s�m�S�ꙅP��S�<��ԪmU�=o���)�c5zP/'i�\�2�˯���Ml��>����z����&�|{�)�ث뀛�8�ҰWjU���x�y]E��8Q�]����:�,��5^�f����+��E�K[�4�Uεp�?F��,����A^ێ!�ز�g<��l��\/v2��5��%9��:qX$!Z$ww����p�n�T�_i\�����eH]W����ڕK5��sm\K����PH��B%
=}�ց��{�D��iޞʭ%T��4�ז�ͨ0ܬ�������]W���kw+>�\c.m��IA�v�oK���O�z��5��V2p�
f��༑��:���̬y�u��V�E�F�|T:�r*��=��FjX�wF��jK��ՙ�qfK}�/f�ϗ�'Pۿ�ɇ�(���Ji���aS9|ڒ�܃�^�*������]n�Lm�����v��pvR��1}���|�����ͽˣ�jY��{B��5��s��f���r�ҍ����_BR}*�;�字���]����
>��cK��a��n����d�ӎ<��Cx�_x�����@@���{���=%y���o-_|�rq�d�I�i��rL��E!�W٢:*x�fh|����k\��y(d5��|U�v�^��UH���=u%K�{KPӡy]3燞:BG������O��W�]���I��Fj熻;(:���n��ga�nU�5���b�M�B��,�L]v��]�u�/��և �gn��H5/w�B(Mٽ���]��ř��309K�?�G#�H%��9/K<^�.bOn����q8��E����k��W��J�.�49t���u�"��X���5���}mgXI��͟sN�<[;V����C3fE��6�v�Se[��¾�觵�3}:�jMK��%�e�6����5yDve�q��/Z��B�zfE�SA�H�cZ��sx2��/�����8v�죠�ӿBY��'!��V�G�e�8����k�nO<.Qo��-�&�{��+�ݔ�J��R�Ls��4��Z�u+�eT�j����l(�m[H�gs�K��p*>����۵�d+�f:����O�oMO+��x�:���N��~�～kη����'�q� ����i�M�Bs�;I�OPٻ�O:<�x�m^Xx�N2m=���}�r�ᙻ�9ןw��2��!4���p�N'����'�O:�Y�M�@��d���N ��u��!�5>�N&�'��߸q�iP���2{�'��<d���w�:�k���e����0�*b��=�v�ۘ�ZU#pL䶳�a�zmNS��: ���c�`o�����v�Z��kc�ˎ=3yx�>m�'�6 9(�k�i6��j�6'����dtI<g}}�Zۇu.�B��1��hg��6���^�i�ʲ���)˛��O�g���zԝ2m+!�6��xe�d�%gP�$�	ѯ�C�M��jw�I�d�V{�	��C��Y8�d�3�y���<F�M������f_W��GI'���ֲO'��Y%d���O���f��<N�8��a>aS�6��38�ɳ���M��*k~�M���B?^:�����ltU�|�U���X���8f2m��t�	��'�k$�$�z�V��2�q�Ь����O�2OP�juCh,'ɯ�m��XU��g�ݕ�ʹ���Ǧc�1�>F{���sxq�$�����'����N>�}�d�I>Mf�J�ԇV����b��`z�6��c$���k���d&�.��/�n��ފ�3�z�譨����+P�x�m������!P�o_|��N�� q�N�;��Bm�2k��VI�o,�'�����h,5�;}y��_{�j�߾����z���'0�N$�u5̇L�g�d��!�w��I��w���'�'{�vɦN�>�� ��'i4��I�:d�޲����9�]���K�J���1U˾�	����)��\�Å�q'q�0��$�tk�'�d�f�{��'Y���N�P�>ɶOM��;d퇬j����zíl�o���b��Y��=�������{�b3�J���׉+'�te�I�5���'��l8�I�{;����a�w������ |<g޹�ywp�Գ�����[���Y<I�>�l�'�Y��N!�'S��Y&��VJ�����䬕&�8��T���m����x�N2m��7^�	S��Q��"}�^Vo�j�s��i��x��)�d��S>I�s!P��kvChx����L�i5�y%J�a˶��L�m$�S��z��}��x�ߟ
�s��^�e^��N�$�d����u��^�y�*�f�-��Q�鼬QJ,�0V�^N�Lffc[�H2:�����J�;�Gw4�gҟ-u��x�7�M=�.v�ۘY(l5����X���s��]�>�/�d��N�1�G8w�Y��������=�5�&�/��"��c�&}�>�LG�r�z����{�d���_s0�	�k|ɤ�AHjs�
�Ӷ ��x��z��x�Rj}�I{�M�=�Y8����~@��w|��Bsy}�T�<��}��>�2����'l8��~�3L�C����$Ĭ:7�Ad���8�h)y̞$�'�Xw�!Ğ$��d��'��s���xf%ݻ��Y"�/��71�d��#�>2q5&X|�;|N�t��C�S��&�m���<gL�b��$�0��È,��~a�O����m�Ĭ>����}�R�&���紪���b#�">���>dזE�OY>ML���$�*a=g��4�l'F����'q'���|��8���$�0���t�<C����O'�>��#;>[�/.�}}��Gܪ#gѶO_Rx}`z�a�]�Ld�S�O���&�S,'oi��6�<J�jÌ6�tk�!�M��jw�I�d���� �g�#Xy�B�톢��ޏ\ǜ�}�j9�I<C�~�l���w�p�'>}I�Nަ��VN u;����0��3�N&��l�ĩ�Ն�RL��ϱ>6�����}z�~�����ɴ��Rm�Ԭ�߸i8���f�N0~�6��}9��	��'}k$��q�k$��`u�R�t�l�Y�&ӳ���>�����6�hN�ό���3S)&u�P��iX;���&ҳF���t}̜��8û����O<�d�}I�d�a6�f�J��C�޺���s���3�w�o�ݏ��6��ԝ3�RC�N&���q3]{���$�Y�Cl�J��t�2q��{�	���ߔ�2t����q�'l���$�?$�޻�w�w�����G��\��}�l�Ѝ{�}>�8¤��Hz�8�2��|�i�����I1�}��&����vɶN>!�,�����=d铫�]����f�eŃ�]��T�{�o8�3����7��[��p�P&{.�ރl�(�^�p�N��,A�('S4�3���?�Ry��/�β%�'��m�O��R��ʿ�v���9�OK"5���l��5\j%@N��u�j8Ad`:����c��˞�ﯸN�=a�x�|�d�	���x�}�IPP��>B��
N���d�k$�&ӣ^�|�0�gy��q�!����{'��i^�����[6�u��=I9����'l�$��y'l����,'�铩�dY&��VJ�����
�Ĩ@���>Maa6���^�>��yϬT��+EgY�D�wv�@f�����'�s=��I�;3�i����8ɦ w9̓��ORt�r��2t��m�z�*T�ݤ��%d4"!O����������eP�����2F-p��Z��)<d��>��̚C^�&�'��3�i'&�y�L�0��9�Xt��h�	�<d�z�XM��}u�>�aYh���^U�F-�7r9sVO<�8e'��2|���m�޽���'8��7�+�M0���u$�T:��8Ì�l�:d�
C�s!P�O��_��G����eV��mT���>�/=�I�N{�����{�,�=�te'M=�^��&��]�v���&�����q�����I1��~��I�_T}>󘉘�_ݙ�,����ϖ*��܅CL��C�C��s�a�	���䗻$��O�q5Ն�����;�P�l�Z�Y�N�q'���=M2m�|���yL@�����r�eQ F%���r�'�)&';�Y6�	�����d�+ϩ0�ί�<Hq��GT��m�	��'IXx�4�4�I>a95�&�{��9��ފ|8Æj�z��mŞ���������O�����XOY���M���'i>d��'���z�׺�&�4yI�Y8���P�'��ML�Ͻ�	��݄��.�>.�w2���||�u�z�2z���5�z��6���&�q����L��w>�N$�+!�)�N2x���TN޾�IY6��O�>�yϘ����#�f���"A��Jf� �g$li���_WN�~�Y��u���Ɲ���13y�o��3�d��1kwO�r�t�x5�3A!�Q�b���zl��ti���;MT�^���c�]J��'�OD�`�w%S�U�9��Om�������*����
cg�3�B!��eN�a�Iץ�8���`��N%Oz��a�M��L'v}�8�����aē�ĝ����I�=��|���8���`�NQ�IP��G���>�������!Y6�2ϘO��֬8��g^�d�T��� ��&Ҧ���M���?2N0�o0�#�'����FznۡY�����z����*}����O'��k	Rz���x���6�����I6�q�z���:��	�ѯ�I�V��AI�NyC�{���-��T�o�$u�]�g�h=��B��{�>��ǌ�����q��G5����Y+R��Ĭ�AaԴ��q&٣.0�$�g�N�&>g���+z�{}���|ׯ�g;�����M����q	��x���'L���̝��9�XM�̜꒤�����V,&{O���AaԴ��m�����|�l�޵��=o��zk��޻��^t��p1:a>g3̇>��<����Hzy�6��	��xq�N�:d딜f�4ä���:d�T����}d�	�t�
�Ĩ����M^�/]�]u�;���n���x��p��8Ì�[�ی�i���9�'�;��6��N<ar�2i���a��;I���I��'�:N��!�$��Y&���y緞��o�W##���3�ɏ	�d�I:�m��	�OY�~�q�I���!_Y8��ﮦ�N;a�g0�2M�<��&�x��Y8�2x��}���w~��u�c�����i޻��=CԜ�X	�N��IR����%I�+'S)6��'�XM�0י4���M���
퓤7<�'�&'o��N$�y����>�5��y�߽���<b����
��<Af��8���M��&�h>�$�XM�rȲ}݁��M����=��&����Ԛd�C߰��N�oZ����ߒ�:U��`6���/�hT��2,�9G�zV�MO��#�c����q�yvfQh���ṋ����4l;;�=�����X��%{�}9�ӛV�ml�������2�lΧҝBs��ȶ��8j�I23����!}2�N)ӎ,;�bV��=I�����h,Ns!P�'�Xk�C�<d�ް�m�ڲWL�~�Nj��|uCl����vd����s~B����|�XW�&c�c�'>� |�@��x�z¡��$��ߘq��9C��I�*�Hq'��u�I8�����$߶Ol�Mu�}�ʯ���o6�sy}�ُyI�}�0��]��4��$���=M2q�t��8���XO��Ì�J���2x�䞲���<d��g�&�#���rf8�o�EW'�R'������V���MX|�x�f����Btk�=f�6��5�z�8���$�!�����$����2m*�^ q��)�)��ϵ���ǻ�z L{�@�z��LwI�Rt��k,����IY�I�Vt�q	׵C6�ɾ��=Cl�J���Bm'�����$��y�g[�1?W|�.���/�O����S�yI�u���I�Fk$��`u�'�I�M�S(O�N&��l'�*u�Ad�צ8�ɠ��"�i6ʛ��o�pr���(���q5IMZ?Dz�<�����w,�l;7�q���'���N�>�Y'�&�f�J��AC�VN0�e��:d�k)���8���XO�z��o>�_��u���~�������J��a�I�*k~d�d���~I8ò� ����N��䓏̚�M��%��Rz��Z2�m�N���d�l�ή���߳z�|��}�|1�|�I�Xz�2Ly����iX<�hd�9�	P�o_|��N����i;d��	�|ɭs��Y�tų^��Lz��c����
/o�E}�'HVOXp�����I�O���r&�&7�d�� Nj�S�OM��8퓶N�;w�z����
���UvR��n�u-�����ڮ���n��03+�Ѩ���B�g����:���wM��ڧ�<���'p@m]��q�Q)!��;<a��jkt��\��z���]�V��Vv<t���(u�U ��ݠf��$�lN��C[���ś�K�k'O}B����'�a*
����Z�6��Q$�'�^�>�$�4w��q���^`v�v��f}�l�0��y�l��:}+C
7bj��k3Q��ſG�}��z�O�'Ɍ�>��8�A�a*
wi+'�u��m'̣	�OS�{�㌓l�{����=�6�8���cJ-�/�y��X��=S�t�=�D��ɤ� voxN3L��g�C�Oy��m��$�XM��VO��ve&�8��T���m��,<q'6��ݗn+�QP*q����s�}�@�1�>��uGLf�o��2M��2|���
�L� �[�C�N���&�h����I3�l+'�h�d�I̦�<>�;���^k��u�s�Y;Bs^d����N'i��y!]�톧�g&%a���q��5�d�M��59̅Cl� ��v�}Y�&�{�%Ւm�/^r���y���s����s߸E���L�x�i�5<�������O��IĞ��@��d����d���F�È,���N$�
CS���M�z��RI�L�{�����󮏾8Ol>{T���ϣ�>�ݕ�	ɏ{��hN�>Me��'o���6�y���8��M������&ؽ��$�0���q�bto�8��VC_k���������\Ͼ3����:d�+P<@�μ�'���/I>d�|a=|I�h�a=g]�i��N�}���N$�O=�$�2q��]x�{�f��k��u��ߞ��:ﯸ|�d�!�a�N%d5y���z���OO:�c&���tɴ�'ot�&Y�I�T�0��a�8�k���k�9��G|6���5��ߟlu߿rN�����i6��gHhy�0�&�����8��O�Ry�����$��@�'�d�C̲3�N%f�'�S�ݽoZּ�2��/��?��d�%[�w�j��{H�;3�.��*e�M1x���)��ýnH;f3ݕxf���$�vW�ލE�	���VX�Z赁,Z��i��_	k4�["=Ks!mp�w�D��Me���zb|��;�z�)�mR�2b���K��)�+f�X���v7\�xb�S����x�����9A�\sq�]g{l�������J%	��-p�u���z/g��\r%��Omfv����kf>��u�e����Hp�\�	��*^�7��X�K�|�X���Jm(�(M�Tc��[���ľp�T�.�Z��[�:�u����F('\���A�����(m����vš���p���VU��9ΤI��F�i����X4�u*AKR4p�rT�#U�j�v���^=۫[�OVϺ%C�-a����|�V�95:��/+�5݀;`���o3d6
��fxr���:���π.�M�Z�6G�6]3X�j,�bb�5�s���6]e��&�ML�ޜ�P�T��r��J��cn�H6c"����ξ��vΔ]^Uy�\�;����g�����:��h �u�����b	�=q'K�X�{t���z�M��d�Zy��FI#x[��U���6w�D|N.8^X�%6YY��c̗v>�&ՇcP�GV��sjl솢�i�W��
���	1o3�)x.�5v|v���	���wݡ�`*ۭ�9_aM�RM�[T��s���N;j��UH���8�������$����D2�����UV~;rzط�C�#ۛ�H]�d��qΏ7�0JkY.>�s/��7�k�Ƿ���V���I>���j:�����o��b�5��l�\�>R��lG���u��Zv��f���b�&��ޗD��/;�>��>�A�����Y��4wZkB�	`��j��ٴUEh}�������<|�d�F�A�'D��!8#��Vl����o!�3EbFd���iGAП(e�f#�ƹ��\�sI�}���C��ë�)�~`�U���d��O�f�9�#�9�o�n�D�o���]�'V_
���ĩ��vkj���wXv�+T�em�gvLt�r�1��	�Z��O0a��A���[6� ̭oz�_;�L�z�<���'�,v�\w�*�ik퀂��;�*^v:�ȁe��8��\�5�8������Mp�P��X�}��֮�1R�WE�<��o�Tʋ�Q�U5i�1�b�g>���hN-���Y�z�{]{�9�uw �3C˔�b_csn�M�}MA������V��P�Xf�l;�����*#����n��l�����*a��0%����3P�Q�^:����Ӟf7)L�'F֫:{z��Q6�Hr��:d�D����W�A��c��ܟ_�K=V{���Â92w_=o�9�0��G��U|��:WNo���5�|��9/���}��m��r�Z����.e)r�X`��Rն�5*�R[�&1-Ƃ��-h�6�T��j�̵��*e�(��eqr6�-j*�)r��TVڲ�m11Tr�XڰV�-Q��'T��a:�]Z�:@ą��[�P����e�n(,�*
��j�YF޲�Z#��\��V��I�r�FТ�1��mD�h��Ȃ������b2�2����q�SB�1
Ԕq�F�T!Ke�\\iP��Vň�#i[[X^�L����˘�A�E����V҅J���$PF-�iFڸ�&W���&"����b�˘9+��m[+"�Q�X�,�"�Z9՝ub5+m��LQJZ��b�Es2LAQ�VfW,��.R���2�Y�R�F����ZC-z��.4A+q��X+�"����[Kh1%�TQ���Ebֈ	JJ�dE��*�zJ(�(�QN��E2�lꙇ��{sW�?�я�Gڸ��Y��5��Źf�i,�����[r���ODک2�*��I�ƮV>zz`��|\|g\T�{w�
�z�L'q��'���S��k��
O�6��7��N!�}a�i����d��I��2q�����ֲO�'L�IY8��}CԬ�$�<�������>�wּ������$6�:J�I�g:��
I�^�̜J����"�l�J�o�!P8�_s'>�N0ݰ>t��N�Y'noY&�M��>��}�w�}��7�w�~�=��IX|�p�8����2�>C8ʕ$�����i�c~��&Ұ;�"Ì�{C�=�
�g[ɿ)�>�{<�DG������,[�r������w|9$��'�RVI���RV�->aRq�V��2q*V�O:��i$�F}��&���i�l�{C~�L�{�k����'�k�u�v��g���N�s_`x�����O��&�������J��Ö|�I����M�q5��|�i�׸3L���<�Y7���T��I�<������-Ϫ��*�3K���	�:�cE�I�IO_<�w�/;:�MXf�峍��l8f��䧦xFUL�>��n��n@�.��!��5�5<Lj\��].��7	ZF����v�N����I�^\ݘ��!N6Ԫ^�bj9����A���J��R�f~��|��������WA1�8V��;��&���s�{�z��ݼ�`�2��E��\��fS]�	t���j�6���=�/��ZKWsg�#m:��B�p&a݃��>[�����st�p�z	#���΀�I��ҷ����	����v!	�l
p�3�D�������$�%k��ϸ=��k�R_+�˰x�Cg�����7��9N�G$L�]A����ۃ�oK���|�[+'c�W���[�e�VEO'���*�/�35�U.~�EFս�7}��>�}���v�]�}��y�VN��M��yD�r��w+�i�:�^��B�r��%�{�g�S�u1��5�\mWmoK٤�m8��욃�"��}���L�e���m�
�I1|����"��}s�L���*�����-�Y]���pkA���͡�G�n�w��n��p��(�0�d��H��8�<����˵
6��j���fmKe	N7u�[�ъgjN�NJ���#����5lq�����f��)y��sˤE,ޤ_��q�fv�T�����L1A�pw��n��8Uö4?^�vy��Ĵ�j��j���e
�f;��������0���5���l�F�B����LQqb{�lH&�@�S{$g;�L��(�B�V}���
�uJ$�[�����OieM��f�cԹwe�d}�;xҸ�tl%5T��z���Y8e������#��CR�n=�;����s}���yj����qk���$Նl�N�n�����`Ji�y���K�)���M]F��^����I�x"��%Wc�18�*���,͌-j���L��b��yB>��Պ).i�Ѓw��!\w�����x�k��)ۧU�k��^���*�=ʦ̝�[%���F��,5�W1T�gww	kZ�	����>甍B1�6���J�����],�©}�m����oqw��W8
�o_J��8�\ک\��ڗ4Ewcx�k��b�M��7����*/V���4��^�(�57o#ܿf���h�9Gj^�8��^9JYƢ�4�<��Z��d��P�:�|Tޯd��V���8��u���1}^*)����ҝnVwV��H�<lT��Z�\���=�z�k؀e�HX2��������sQ���$}Cs@)�H�
�\	���YWu�������f���μ��k����������*Р6��'TĐ�$5wc���Q)��^�G3F9ӷ$[Kn�*��4�>��qյ�9ۜ�g,�u�X�u��X�{Àg�n�joVE��ڻ�W~�z(�5����Q�{9jT���o/��jsb'%��H���p=�y*Ȯ7�yP��Uk%�'/%ﹾw�[�q��et���rT73�v�4	��5� �S9�)"JLF+orH��ԓEF�\|��f�۞��ڊ�Ħ�T9t�7;��G*;��eʷx�tE����&�:�)ͩ|5�ǻ��Q�;�<�*`wJ�����9���ZOn/Ĳ'%H����� {�\/`���.ѻ��Z:muTB0�!�	K��ana�:�F���\.���\�իyR7����W��;�V���S�P�9�V�«�<���� ��l�:�i�����\4����e��]�cwKq�WTaK����H �r����d�5��sn�&TnVA�<�F���.�s��m6�H�Jn��]6Ru�-f�q���-p*9��[#�N��Q��}u�S<P|)��ݶ_݃\�]؛� %Jfl�}y�rw`
zZ�h�i�+@` &��t˽�L GuM�����$M#��=��[:y#=�<�.\�x{�+�]qwhX/o�G���.��������[j�S��졒�'��>?���o��V�r��o칶v����7��Fޕ�Y��8T��Bw7"�����K<���~�;1,Z���}�(N���Ǵ�����Os��̽��V7�*/RŻ������-ז]}4��O�ɢ��q�qG�Q�F-j$��79(�ҙT�_��Z���r�u}4���u@Κʆ@s��p>��k��NQ����ϕ2�y��6�(�0�O��*f��K\.��f鋦|#J�a91}	I����hu��(zd@r����}����`��O,��G��]s �ܘ����RY�s�c��4J����ִ�WG�t>0��u=��.+�����	�8�'K�n��1م��5����̼�|k�u*����W�<���x�d�P��E���o���p�s�z���M]2�/GTr�f�sC�~��׳UZH(��f���������-�U4���8m��E�xn��Մ �-�؅ �K�1w�//���.��5�<�f��d�C1m��|�Ǳ�F=ۭ}�r�%NwX3e��
�IN���Ws,�ԣ2qS��U��!��z�������n}p�K���Zm��Ƴ
���\>A(*..܌�[�9	ٞ;N)��j�������j���%��dwn�T=)[�Kd.�̩�jU��Q�#���=K5���m��t�h�]T�(N(�B��ΛN'9I�{�Zi��[�U޴l�[�̚s��z� �4tu���&�%$������q�6��W��UA�v�[�v�gV��i�+Vw?BK��s�i��w������}mb}-�z�gOB�M�"��f��dF�V�9���MI�wͯ�7���z�^Y���(*��=�<��n��4{�m(�í�Ɣ�*g/�R��)U��<+�mH�G�D�c���
i��5El5ڜޔ�t��d��]S|��E����Q� ʨ��8@}%@�Nz���?��Q�iԇb��~:��̵X����F7�t�����L����e�
ۼ��Cr�q���S�O^������d��Ԩ��q��̆c8���1Hc鋋�b�W�Zh��퇏Xy���X\��.4�)J:%e9A�qu#i�����ѯ����� ~Iw�z�9�|��Z�w���Kd�L;-g�R0���S�4rS[��%�l��Qȿb�)��[�qe�fv�N�NJ��h�Gu��wc(�|����&�K�+��폔�O9S?"����Ρ0w�C}��F�i5���ր�i���]��9��q-6���Ѯ��Hʸ�؞�3���5$��.�~Jnk��|#��;W�1�;�n��n\�c�� io5Gk�0��\!=3Ϩ,؋���ש4�2�\Í��{{������H�\'��:�fBS�+]e!5�J5=��)����ܖos��dc��}r�An{ �X�.3+\u�b��`a�Q��aG:��O4$E�[Kr7x�-kT|�Pa�Y&#�T#J�����x�>��4����9L�Ե�׾Q纷�I���>��-��yXq�\2-?�����.�v��`�*��!�ֶ��p�Fm&�RWY)�E�n�Φ��#�9'&b�Zk��p�ugBB��t��헎��wkM��Ԁ0w��	�p��b�����
���Bg:�C�]#��]J�Y]|\�gw>�ꈃ�ع7�/��m�#�YU�{�O���=Oy��|�w��a4����۝�:�2w����bʣ�Tekp���}��oAC�B��e����.���܈8:�#}4��L@Y4[��J/�9�Uݦ��'9����y-�z�.(� ˯GFM"2����Sb8�{�X��mL������Z�� �\cY�G�v�rZ>K���9A�
M,�Ȟ��	�s�61��RqCr^K�s|�%om�ŕ��Έ�hP����P��>�b��.ـ>�dJO�[z�z"��RM�S�<]�����%E��]8��7^�**u�9W��sY~�n�,���t�[�:ڴ{SŸq]/ڪ����U0K�.���x#�I�2vpd�ww*������[��-Wk�锌*�f�69q�����[.$<�����p�܀�k���9]*�물����V�H|O�݉4����x�W|.J�m�cxk��fŰ����0o��]�I#m���Z�����O�XW����s�`��ҫ2�ꙹ;�rl������{;G.j��q.�]ߢ=��|�jFn⑿{u��\Jg/Л9���C0陑�M��U�RU2)Ϩ���֩��j���x�jA��K�p��i��{x��Lh^�s�<;�N=���ez���#<��f�5ͺN�l7+ ������i6�{���5��/i:�h{V��i(�ro���Z�W���m�<�9�Ŭ���k�ϖ�{�L�m+N�i^<�{��{5k����~�OϺ��Ҧz8nq�o陕�=�Z�������m7naË�陼�N�N*�UoF��L��֤�Ż��ڇ�иO!�{��1;s������Q��!���)�L��9��[��9u˯_L�5I��<{s�����%��''�ls���NV�ʙw<�6�{�y�V�	�{�U��St9t�	�q����!�]t?��CRad����!ןM^��l��9Y��;��K�L9���˗Ϯ�{9�H����rv�WG=i=����|x��=�1t�nf�@�ըc��#��Z{�!ϳ@�_v���C�B`�ޢt#�o7�_6ժ�TR̚6���3\&�M�w%�~���{�U��v�0lw|�3 ���GR�Օ��9)1�������n�.��`�ޮ��4���	�.��/pE��d�kx��̇;���oo\�[��k�o+p�)��iO��R����TUNc��f�##����]��Q���/�gݗ.�l%�95unڲ�l#	T�����r�ݮ�o��� �2��E ���㸀�V����u��p�-&{`�
V3���S\��ۛ�u�Xԣ�1�s���W�u�p��A�sgڻ'+���˼u�3:獅��!��jQ>�bk�h�=̉s7} �}��loa��q�d唍#[�6u��w��������t�D˝\�su9���/ѻ�+SPa�Y<�P}}�lҼ1e�{���*�s��=q���B��->����y^�8�\ީ9N=�������\`\�����˟cδ��e=�4Ȇ�A*���]6�]F�.bq�&h�}��5��+�v�F��W��:`K�l/ ��Η���=9�e��jSf�����驍�qt�M����偟S�#�{K�=oHk!�T1�/F��n�U�-|�J���ھ�3s���(��yr�-I��]Ԍ�6��G5f�_Y�P)��	0�B�[w������Ѥ�WM0+%Y�_a����N���w/����7+�W�c˝��>���>v����:֣W[cn�Њ�U`��z/2����.�m:�3U�e�HoWf�&j]įh���̧m6&>��J.t)�52����TB"oNyסW=�2�ք�݄��Ŋ�7JcZ9]�eX�:���։B莵(�vX�8�dL�{#�1�p�es���5�P�Q��e���OD}-�N��*}S/��G���b��S���U:q�6N(^Qwyͪc:U�ksBˑ�r��/�U�
��fZ�V]��ڛw��9�2$�
u� ��=�l���4�uM0ӦH��M`=�"pu�1���Ξ�=����s�L��KќWW��VeeL�dv\4\��pg!2��[�n샐}95�����(�[t�<���QǕ0�Yيh]ҟ(�=ɒ�7����s�s��������tU��;n��:|9p�F�J��s�f%���*�'�r�V������l: .�1n񩹮�jZ�gr���`�zO;���N��}�Y�ewwМS��{���Q���{�p�͈��;Y�.�+��,M��&�u܇2����x������-�5:���GQ���k�����[z�3��(&oC���o4��r��ިɊm�F+�S]�0�N{9ͣC�Xv1.˞9.�q�W1:kx�Q�Io�Z����Y��+��14��Sv�[F)���Sx�w[y �!զ�9vv\���t��]��y˻Pa�wXt��s���vBo*��dg%�(ӷ�D������-Vc0^n��ֶ���.�m��j^��GJ����h��H6L��Q���Y{�+����d੾z4�W1'�P��y7�
)"Ų�ӕ�z�w.!r�.r�r�Y�5��P�9��o��	.}�e��t̩yj���+vPO0�`�}��kp0�9KN�TtB�k��c��L�P6�5��,��Y��2֒�@�ݲm;��Kъٻ��2՟t͗7��h�#=E q>�G�nu	OUl�E]n�X���F���A�X�pR)[MJt)f�ɷus�;>��J�h���&�[���};��j�N�så�ut��!��IɗX{���C�ݐ���h\���fG/4�vqw���<��c�R瓑r��Xy����l���#�� ������G��\W���\�wa���+� ���;��O��:?DU@�+KkmQE�iAV"�aX"�PG��
Db�b�(��U�(�""�����%��QQ*��VbPĨ��ʖ0DUDH��AUbőG�
���(�TDE��E�[jZ�+*�U�[jF�FVb�YX���EDYJ�V,DF*��t�G*�,X+-��R,1�" �"�P�4`�*�V�DX*(!Ȍm�QEq�"���J�b�T�$PX��*1���F*0d�*����F*t�Db��`(*�bUA�Q������$����Ǫr�Q�,�IDm�`���*�������(*��"!��"�AU���(q*���UADX��"1g��;�\�����7��׾���cv�v����b�g<�۱�L�êV��T�Ի�z���
�����<�#��MfNS���諭��M��U�9L��j�xu���8�sq�����(��Q�lW���x_����Ʒ�N�X_�Ǵ����iL�S=�R^7�,����K�4��^L�|���-���&�]�ɢ�V�Q}�ʍ)�L��u{F��X���\��7K�>]�~�̃.���cd[o���5�噏j�Y
��\���x��!
{Zՠ�nC��ۅk�#P��:��̜����� I-v���Z��vpSw�g������<�Qg�u:���rTT�Ue�=�k�ҋU�[N��!%'���R��o�ۅ���*�8z��\�:����9]����7}�o΋M]Sh�C�w^u(�Cf���qv6ڕ�ytӌ���TW.19���E��d�K���;�*]d=��g�_;KMf-���U�#0"����m��N�I��>7��\�z�0�z�*����lA�+���[��[��u !��tb�_cŧ]�R����w�����srV]Ww��Z��>>׊���>����nG�v�LӝΟm�v��R���|l"v٩A;|n ¢�� ��p�|��17/��{Wu�����{��&�&���u^���~I�����5S9䧦��1HG�j�̨gp(����b�W!�j���;�\�҂��A���\fVC����VeD��J�����Y�m����Q[�M-j�eA��d�yH��%8�Ff����]j�E�?U�����緸��˜�S��;5<�����W���gI��P����`;�Ux���zT\F�es�+Z���L����+�Z������ٕ�4�d�>��,fʣ�T\a����Nf%��i�N��Q�\��NK��j��V�Y�����Y.�sPs�mvi֔��*Η�)L涱C��p�����:�����R�D��>�Cu�5ʏ������O����ۊ<������\jU��!Ȫ�9�M0%�3��B�<���ܷ�󸕽���C+�N`�V���#�>��WrdSψ�6����[}��.�uĹJ�CqZ�Y]��	x�Bש�T�}��6�������:ODx��"��"��/V��}��]�<�;/�U�*������i;��ާf�n�z�ۣ;/45��".a�<�^�i�������w;2g�`r����D�2�YÒ��V���Ks�&��A��Z�z���g�צ^�����jy9T��5��<��:�3\��R�'������}mٵ�HʨU0K���\`G:;��I�G���3�D��M.�[�n&7��&�Yu����Ќ*�3_��EB��~�W\�L�������-pnw\jMXf��%3����o]B�AW3^���/�,V�甒����2�uu�M��}��k���nk ���.7����9�Y7�LْX��k]E���uxĿG6��������>���f�¯{>��-ͬ���sl�'���Z���-c�|\����G���+t+��1$��1zE���=��z��s�i^<�gW9�O6�7q���^���m��^�0�-�����bi���HZ�Y]�U|u~g�}���{���]7���uA�K;I��Cu%A�WP��Є�� pgLnXֺ�D'r��e�x�1`B���"�U��'���XV꺅va�ݤm�F��Y
ޭC�0�s�gTz�%��|�v޴�V�뽨��ɜU$�o.�I�������8��.LI��K��EE�N>n�|��0����Ӂ�ɤ`[2jy�za�1o7m4�wj���;�z+����S0����'���ˤe�␬N�օy2�"5n��pWt�1t�Y4zV�Q��	��}
�w<�[o;c�n�;�վÆ�,����P�{6Q�)��ё�l�wI��O�t��=?Fb�7�f�t��ꤴډ�l�u#�5�dJL(n�HЫ��8�͌nn-dP��w[���]���1W!�h�C=�N�ɦ�ZLV�/gou�z1�֌�S���ý�s�|g+�`C�QS����J/:��uú4;�.[w����%��WL�OC�#
��w�y�#�K���ŏU��g������j]�l�n����vX̙�L����I�s�ܑ�\����oj�دX�x��Թ�Z�:�OEmr��7ܝ�MH���>����کvUX�Hw�zˎ��A���:��<�!�����p&^�)����בC#{�⫔�>��Y���s��r���"�Ȭ�^ٗ��wVz���+�a{d�Ϊ2&��^-NI�w+磌��w�{5���f_�auL����-t�Ӎ皔Lf�&;��t%�=�x7��tr����F:�UFúٍh������x'_-75KVw4���7Л��y���[��+�yt�_4^��Wh�џE�V��O���\�lZ}&��q�+3�7�Y�V1F��J�_,:��f��'Y�7����j��q�Ra���-�&�W\���y��Kd%�B��`v�jU��T\a����}
�ˎmH�h��TO+����ө���2��<���&�����Nn4���%lm��������Ђx���̃.��4���J�������ӎg�^�	>�pw�b��T�� �n>���0�D�GR k����H:�2:�m����=��ˇ�� ����=e�fv�N�J��<�oЅ��39�~������D#���;�q'��s��pG&5��Bu�,nY��#qݖM<�ݗg�]�p�55���H� Wa�C:ܛ�A� �I�j�uf��%;N�M��*���R��uٚy�t/ xt�W��v����.C��������BsG4�[���l���E<�}")f�\+}m�ކgkVD�/t����]0қ���|#�D�&���������ѣ��a�&���t;�sN��*�*`DwJ��˦9��F-'�[��6�u2�p�S��+�`���R;V�S0�����@������1};��l�31�S��V��yʸ�1���J��M��e�p���zek���me�n��򶈽+ik�ޔLf�g��W�Cs�䲡\fS�7Vq�a͑���mf�&6� �qj���������Q�eA�nVI�yH���C��u��ɬ�)6�c-8i��k#{���}%s�KAo̌+pjk�53�{�5V�n��a�1�6�W:���-YZV��2���~���}Ս�[���u/"s�߾�s�J��ڕ�}�����*�{J�í���Kӟ=�����`V�>�:(�ރ���
:�G���+j.ep%»{�g���%��HR���ԮD�nn��Emu�2�8)v��{-�qK��/4�*�.�B��7����������c}!�o+�������|��g��u�x�Y3�˾V_�3 ��O.3�fi��-}�v㵩/�Ã��>��F�`,��F\�5*Xe8[ܢN�@Q�����aS9q��z��6��.�&�L,��D�����sn)�g��j���jL-M�KV�1�ۣ�jw�35�)���q�^ŮPl�1t����q��qCr�^���q+{oء�� �㘟lw>�o�s\7Q9=�Ԍ�ֲ'���+oq�[�UQ;re��k���&�����h�ҩڞ�:������5�*�̛�ʚ���q]�ޭ���������+��T�`>�˦9��RgyŌ���z�5�(^���}a<����t��aR3	K���K�ݾ�y�KZ۪��(�N-γ�5a�눔�N��W�~U���5. 
�H��WkQc���/h;9�����R�m_���nk �Y�~��ϗ��9��Lx*6{B���r�>�ĜF���f4�SJ�
���&4����9&i��1�3����;�����������˨vu�z������,���&��'t�h`{R�:����X���q�{m��ÿ��:M��fU� 3L���h�w��|9���t��M�:�G����ۤ�F�Su�����d�����XQ�g9;���+�����6c��A��[�MF�7<)�쇋�r��<�Q��N�ʌ4�\�1��Q̲��)�]����W\]]���%j��p����}-����ʌ8��DnZ��u�.���[y��RU<�o�v��N3���֤��-k���U�ԯ:�iZ�y��{�3'i�sG����Q�2������=o�\�ьa:��r�ݓZFWOd����Nyjgʙw<�d]I�I�r��H�[���ΎiWl��)5�a9;��[n��E
��^���B���q��t,�E#�gjr[#�L���A�ƪ���\�>�Ҭ�Qȼs�➪��^���fv��v��EN�>������	씒���4�P}PZ9��0]�=a>��L����?	�rh*�^׆�i�?[ ��؈Hlޙ�z��R��٨�n'�˵�`�:�GI�*����N���Kb��n�'ܳ�@1�[���}����G��G�"��sR�s{�P�[ܹV�g���u����Ԫ��U�Q�h��o9�Q)�5�5� �2���
EXI�Ļ��@Krj���V_F���\�`�KI�ʤrS����:�;{x�j�7��^���KBY�ʑ.�i����(����B�@�BP�9F��<s�
�=b�!�\S��<�(���('�����e\�ݕx^���F�ld�U�l��r�旅�5L5���8M꼹%�v6�~�u�K,x&=rO�����/9!\/�*�YK�LPSyqű�Z|�4�uf������J����|��MI�>nih��L5.zd�Y��ĭoY�2���9r���hZ��
�uB(��m@t�:N��Ӊ�=2��`y1�P6���f������S��J���U���ͻr�}�k��W[0Spco؝�-�b�I���=��Ym>׉��6o�\��V&����k��O>�2�.��os���ˣ���^t�~�h`�=D��I��)�n`UtV49ԇ��]��ɼ�J�k۬��)L7Hk`´��ӹ	E֨G���./�V:).$��i7���3;����f"u�T���)q�+u9�cBj�Y���ʱWͭ���\��ן&b�Ik���\ʩ%ww-���z=��>v���$G�˝��8�20 Cf������NTNN�`A����ӎ>v`���u[|���l&�W��{��Zr_�ddx>���G���-WP�t.J�k��v��H{�A �����,�_(�T��Ьd���FF�G��K���,o80v�|��Ar@S��d��~�hK�*L�
XU�"��C�wbvO���ꓛ�Q�m=����
�F���g�-�!F�k��>>���D�Qr�]�����wy�R����]&1�"k��J�#��qP���^z���.��2"R6�7&8Ed�ΎYϏ>�ܷ{�Hq0�t�ôH��C�`WR� ){��;�\ơ�M����}#�E�F�����ނ�uf���j����ח�uAЮUʅ
�I�9�7J�9��r�<�E��tq�Ԍ�X8C��c�v�dK���0�蛇Nt�ٙr}&f`y* �����z�6b��jj��EA�y}|��t��W&�bK%D�sJv.9�ɗ*�	}�[��^���QN5p��"�mI�'�$�޵𥽛q�N��YV衜��ݨe���W��ؙ���ͧ�Wk}8�������\ ���q�,Nv2�v��Gte]��MI�c-�V^�ȏ���F��G��̩���|L�[58>�TΤ�]R���kK&7ˮ�wa��Hn�$������^]op0���տeƵ N�_+���d6h�"����N�Y]J��Z⣼�Mr�r�q( �y�6��|�x��˪R�Lx��74����2/�/	�V��VW/�T���2�nXu�Q;�}�>ޚt�p���_JJ�t!��g�R��ՠ�{�ӈ�n�|�u���뺝l�&h.=�j���c�u6Hݞ�O2��#}��b���8���=�ǖ�;C�M�/!��I��h;�#6��w�p��0���&�Q�t���_4n6mi�vr��h\X�)5nm4ҹ1��� ��0C0�w��20�T��Ҭ��x�����O�1u�qe.sd?��[���U�*�N���81ԡUܑ��R�8�WZ�\�s��pR#1K�\�3"�[�>���s��E|E����ά�rv5�-3e��.�6���z&��oQ�[�{�M��{Ee��Z�C���b�&A$7��YC�����1��jue�t��x�G�o�u�]�ձp螊' �8b7D�ʓ��&:nh�w�t6y`�ԵP��V�H�\&� r�V,+��f:F7y��F�E�Y�Qr�r{�$�5��V].̢�f��"�����V�2
��Lv)MPگ{�{:I���|Oy���ey+�Q�7���r��s�uM�����X{4&��ɲ��_�a���}}g�[I �ّW��������)&h�fr;�l->�U����H-v9l9Lc�x9L�0k��k/����W�.3��[]7����/o$]�9.�JҀ>���&J7G1뷧����5<�����g{�ڏ'']���a�;��tD���h��Z�8�-T����;���8}|��{x[z�k[��)�z(�l�yK	�Z�H]��^�Ԧ��I�h�{WLq�Z�@\_ʳ��{)3C)fvv����<c{\Qh\����<�7[���g��y��nݭ�#��r�~)t�r�������}SI�NU�f��5}���ᤥgHW��X��]�܁�{'f����
1��lq�Q�ջ�h!�]�L�g\/�oA���ውI=�Ŧ����ջB�)�wGED��kz��� ]����\/9��	�A�eWT���r�oR�@뮢W��+��	��y֞HԳHH乚b����]�R�
�9��sG�c�B@L]|Uo���������׼�s�$����KwZ��ĳy����2���wІ^v�-.j�3oV��b���R�0�3��'3�}w�	悁���JPF�-J�e�qw*+S@U�tm���oa����<�_��q�uh�E��XT�0D��E������B�($EX��*������8�EH�PX1��bȫ�DEVƪ��"��PF ���� ���(Ƞ��D��YE�U��1�� �Q��9kh*�*`��1V"�1��AA �[�V��Pr�H���Q��TamX�X�-QQrʨ�b �d�TUb�`�QKi*TUF[(�bэ*�%h��,\s)�T�ʖ��V(��L3E��Z1U����m\�m`����R�nAFکmUA��3+i�+2�\1�b`%�UI�\����--�ȋ�e�b8�*V�EY�0��-���iJ�������f8�*UU+�B��M禵ק����b�R�_��66�O��V���f���Gn�O�v㼧S��}�50p�Q��{�%M=v�K�Zn=��������k~����w��\���P,��9��/�;� ��Sb�Q6�4\"�f!�����`s������3.�ɕ�m�ὼ�y+z��s{����a鎉��L��)�V�3*;U����m�S~YFϧ*�4<i�����sǆV޹�^��v@{k,��Dm�I@9k�g��n��î��^��0=�k0N{i��!����Ndv$�SP�U[S���W�(��U�=��p�ɝ�ZՉ�z�f�lj���	����ԋΰ����nSY��ʤ�<�ש�5�s0���7Ӽ���R�ȗcg89[�����1��q�X,�l=�W�j@�dޛ���%�)��TQ�Q&��y1ބ_[�<
4)��&:aY����n��*�C�C��>F��K�Z:S��N~ ;U2܋��1-�C�U�:t�Ψ����0��^����R
�+��C� =RFӔ$t���w5t�`MƼ0�c�W7}�R���\������AMj�ګ�0J�R�3�*�P� i=C�������b���^����{>��ߛ�޽�;�fzQ[KGb4c�飖M��QV5�vuEDV�ɑV�
�T)K�Y��岸��*�7�H��F���LUr�VN:�xHً&�
�;6��P��(N]�o�|�.�1�@G����ժ����Σ���7ɣ�7}۷����#ޏR��V��Ԧ1w�����g!�+ɶwBY�H����q5�9���yݩ�e�1�X]v{��j��Q^�[J_e�;ܓ���0^\���W�� _{�f�IG�|�T	�p"��1i
����F�F�s�u�t�l0�g��S������.�y��ҷ�a����.�����\��H�.��
C�p�Y1�q�Ы�� ������I4���]*A﫣|%e�J�":��E#����!��[��
\����&�p�*�-/e47��nĸJ��D��+&��	�}e���\�u��R�p��_��uQQ�	/>�\T��!�͙^�w��pz���mx��+��9����RCF-w��k�Ž�]��D�:���z���O�ϵX�n�p�WQxq���`��֏1�����S��Nv�ÔpC����9��4�c٭���P�K��9C&�Rv���!�8�xc[ڌ=�K�ȗ%����S~�*�tË�a0���E�e��������顒Ѹ"s����.�޶#"�9�t��@~V��@����N桌 �Y�+2��7ԛӖ#��� 23-�gP@Zʶ�0��ػ9�;y�����*]oo�c��gV�P�M����PwJ;�q*`��ͮshj�V���.�]'s{yo/ޏ{���؝��{raML\���]����i�/x�����b�.�n����{�s�9�r�(���|kF	�<U�Q��
�K��m���l��J$����(����8��{��(!1���4+�l�.�|.#�&�3������'�YҞOB�޺��qc�,�-S޻� � �ڏE��>�|*m�+z9�$/���H��M8�����G5m9�|Q�˳9��T-&���>]Ӱ��M�= �O�e!��b�p.��������n|�I�y���ء�=@�����kUҗt���b����}ɫ�3�)�Y�c��&uF@�f�$��%��_��D�:�R�o�����+
w�EKC)��Q.jęH��Vv-l����f���È5�4 �BT'�1J��T�#8��P�#�!�nW��)��fj~���6�-��A���Εv�I�^��\�y��&��ӷ����ԋI����}�jA��>+����v+�_$+���*甞AM��~�s��6m
;��,�v�O���*��mc�s�JM7��]I�a����M�^���
R��|˗%�]Ƙ]�$�	�y�����s�o���R���+'�k���w��ElO�n��ه5,E1�_2n��S����O���������߲��W�L�^F9�{�|���z�}�Yԭk���ɟ��	����m�K_��od�}���r7����t��Q�6ƑS1�.qQ]��
po;3�MKP����ގ��n�`�*Y�X�ex_Uqpr����¬8��뭘<�լ�!�Ug#{�X9����R�3�}Uڴ:ُ�Äׇ�i]R�`�.X\DjǼG�l�u�-��9�e�����0Z✈���p�8U�����,]�$)������:���)���c��f���[<�wr�
���1�(��ޫ"\�Jh�~��A��Mlo;ڹ6��V�:�q10�W��](�-U=
\*f3C�9Ь��"zO��9i��7qY;x9� �����Fzb����p1T����Xz�@U�"��C�wbv]ݻw3�6]�l];�á�O�t�.*�K�<L�>�)H��6���	]x�E��'�&y�t�j��%�����(�R�l�2�����H��5p�d���^z���.��2%!�q���X����B�lQ���K�%��T��Bk���S�����3]hY�K^]�c�>�m�2q=�+���[=\�U�y-�Z4���q���r�Ӂ�6��k���.jQS�f=�.��޵@ˬ�+y��<3{;9b-���f�iV
��kޕ5
y}�B����F�򾯾����zN�b�a������Ъ�`뻥p�5�8 �o�)K7�Pw���C����ϊ��(���a{�SrWޮ�ٿJ���?2vO:dI��^�`%5��7�^L���j�l�}�Թ�#��(p�J��ݹY.�0ج�t�L; x0��u�I6�=k�3�	�Ւ\3h����{�⤧V�,�J��niNźs��.r")���(�r�7߳�lM��c�*���@챹X�����(��#����;<:�s��}��ŏVF�d&ej�����]�&/1�J��!���<�NP���q2�n��o&�+̮踗���4���]d��И}����>U.&8*r��S״P�)qh+u���q��n�p��zo���j�plm2���`{���.��6
	�J�ֆ��4_F7�$�����)轲�ߕ93�p��~z�n�f��m�Bc��o��)R	��b��:���R����enʳr߇��mKUL���=�C�\�獕9 �s�]͡�Ѩ;��_{��������;>Lu�:o�R멥���o����\�1����b˓N��^tM�����5k7{O#��2��J�t��������{hi���(���d`_d��4m���h���=$뫕0W_#�������h9���+z{$��!�U9`qQG��ě��Gɂ��s��z3B��[y��n�"��Y��2.a:2nY�p�K�Z=�9x8���J��#�r��ݙ���Qx��m��Pc�.J�D踀0:>��+�W2f�)��׆���3p��Uۍ��� ���Ԝ�Pй��qK���GS��D�JT�s���Y]�M�x��:x^�`�-wG���Y^��m�C�W�x�a�	g��1S�&�C�u,O�%+t���[��V���q�8&�/�D�3�T\��&�6v3|?��9��L�,ș���W�"�[���mkPVZ����?.Qғ��M���l�gX��%��;��O!7��^�.﷖�ەlz�B�G�ixV��R�0+!��R0�;��.MJ�x��'}e��>������;A���t$��y�eR��H��V6�������h
���6�d����l��7�t@�Y�u	[Ȋ�O����t�f���qyT�μ�]��t��.㿏X<6b�Dܸv��O^K�Y��C3n(�����ն�z��e�]؄�wu��*Fn��r�����69HB�_м�s��H��C~��;9n)�Wn�N�+1����(�Z��N`wա�;_R�Q�gWt�����ﾯ���)�"�����F�.ff�CBd�xT��8}�F����P������N�6��<e�}�w�b�g��l8�
vY\\MJֈ��+@����ʅ9�t�h���20^������/�[-\a6�.1u�9�ۥa�Fٍb�[5�p���7��+V��nr��S��\{s�r�K[@�uX��R��s���x��\F�	��.�6[�J�n��9��n�J�OC�7j�׵} �)��������)r�]N`=���� /��i���n�a�R��)�;zU���>���zS�^-����ґY.�҉�=����eQi��(;� o1^�����6WHz�r�(肴;��� �b�!��۴�"s�S�N^ں"��s��
���Ļu�OC|V�qI�t'�$OI���IZ�)��q|*�mH��)�0�%����Wt�6L=wY�'ٲ��}�M塺��얰2:�����e:�re�T0I�����J�ơ��,\ށ=b&����]��������M�X���^@�������N�u������qڒM����O7�8�8��j�OrcP;k ��U��U��ۇ%��k�j\�|�w5�z�e�2��|jKI#I(�bz�U)������Rbi	��y��o/�=�V]�>�r�j����ۡIP`J��E@s�V��<�#��ȧg%lt�0��� [ϴZX;g84�X�����#@J��Q�%��08+�"'�Tr�4����W��2ϖG��p��*�Uǅ*�J�� ��S]��J� ߉r�63�q���x����."6\oPWY��G@l1��'���a�xZ�p{ U�G���ꋵx�vm6�椪QxW��6�G*S{��[n&��aD�!`�j\���M���dB�0����Io�Y����C�xͰ�+�E�jf8\��be�.]�ڬ	�<S�N�ِ!�8�S��J��1������¬8�뭘<������ɸd���';���P6#ެ��
���U�[*O�l�&���b_2������,�EjTe>$�e�x�".��ڠ�챜��N�Ju'�#��Ψ$��d�sW	ss5��U*%��H����.�^!Q�"��;�<n�]Ց.JSE��P�#�����.��;�����6�>��\ӊ�u�N�rJ;��2�n��u�/I�iTͨ+�r�tRZs�r��&�F.P�K��p�n�d��v�e�[>�\ya���̴���j�:.r�x^Ͳ��k^|�H��No����Nz��'�t�����+�Y��_i�K� ��F8�;do��T����>��~uxn����n���J����so�@��q�ܬ�ݒ�T�wB��; ��%����%ɰ�9���xB�����U��(�R�۬��'e�aXtq�%��eRK���[N��^ǂ�A�h	�+z�Pz�v�\!T���cs�L�i�
y�:�͚
��FGJb�*�|����<a��1�ɚ��L�Kf��Ce�v�䒩�d(��Uq��4q�|I�ñR�髑��Rj��Şyڟ4�;꘽����N�&�Zus�['d��2��U�Q10���<&��~���׶��仳���^x��ocR0�@wnVz]6r[D����+�ff;����[{Z�ŎB��t7�0��{����B�Z��L2WK�sm�)ظt�f�Ǜ�m��n�,z��!U��H�r/<�?��+z����)Ҙ��ډ�ɛ�8�چN��zj��E��իF��	����*ab����<���Zτ��0?{5�;�[TѝR^�4ԇ����>����F'�E�p]��K�.�߭�߻��[b4��.���k�vyu�ݝZr����s���&Y�G�	έ$�f9�|$	-�Č��?�-���N��ƃ��vS�̹���oy�!2f_e��e�2�ɀf�p�V����g���W�	��;�x>��骯3ʥ���e��{�ewN5�Ic����j���Tl��̭fc[��#<��;za\F��`��qL��a��+_H��g?��]w"t����\ǣ�kV?q�BǪ�=Ѓ甐��SV���R�o�/�g}�'��v"��Ե׋��RyM�4g��G��.��D �h�����6b�V��+s��h��O�:�UK{4g��i*fk��E��ojPb���\�u2�V�j�F^����wRz�i]=ͽ���ؖ�RKG�?0�W���;��؏��ƃ�c㻎�W���Ҍ�3Z���1�A���m!=(a.��*�_'Ԋ��羐(��ąu�2�o��u�;R��]��t&�
{}'<�7�p�:�
��B���Nx�%����������JY�����u�����l�T�=������~\��D.HХCu}��V=����5=.�/D��������l�w`Ǚ�K���g�M+��b�>����kS�沸��J}\�wh1����d�=��6�2/tJ���Eܙ	J��p9Ďׂ�֮j�v���U"��%)�:�l�iV՝l��!�W��+
5�s3R�[��������[�uQf��*�2�S���)D9��IM݄Զ���X�����k�r�(�H��\�b���}y#��T���r-d��*������h�v�(c[v3�h�J,��9�֮�:��t�f��մk^KAjQ�����g)�d|��I����4�b�ln.c�����$�VJդ�]ws� �J�ZVol|��t�i3���tf�U,�ϞZ�����>��<_,���ʧu�	]t]N�����A�u|�)(������ܵ������G[�|K��z���!�}Ԣ?]��>lw�a�\}�&�f �rJ�
��^m�'���0��١,�����e䨥,�w�q�+�9�k�ȍ���Z/�݀E��������ή��m�{���:W��=Yݹ"�uL��$1�������d;�8�富.j3�Q����=��S�u-��pT�5�w^nG\��<����y�neL`�#���ֻ"�{�@�h�]s1G�:�bu��Kz⋛7ϥ-��3'M�[�p�:�ݓ�T]�|q:�Jt��[��t��j>)���t]=�RX��aP��ߥ$w�9n��]�Ӌ��]u��v.=!�Bu�u�`#�&��v��7Y�?{�������x�;��-�\�v�V���/�9��=�]�c3חD#�Z�7�B���R'C����
v�>Y�nS�-�͘b�Hu쓱���+
�r2�QtV�<֫˶`��յ�;���hC W�=*��ٟK⽗D<����[�+o�U�B��v�u�8|�&��$��#�� �����.5&���,l�e���[(�r "�u`]�+����A�Tj��7��l�Փ�b8�l޽Uu2�J�|��8� \�Sئ��1*Sy�i��m+]).�E@b���,�[w�ڛ����K���H��`ܵuf���X@�_B��!ؠC���p�r�'��a׊��0�Wu��N^�n���#��<�NQ�A�����t�p�t�n��%t��g�V=��qa����K�tr}��=y/"��K*�_V�N%�YWɴyv�0n/�n�̊�MYقo(�6�-�(1�i=�^l�@�P�Z�*[��9訟�X���ښK��gbgcT��u�������".����ʃ��ʼ�	y�5=;��"Q[EG� JR�V���Kca����U��?�HI�!�>���F��o�ժ�I��j$Y7���۱R�WK��k�G�lMಭSzFX5K��]��r�������������\��Dj�&�_cI���Wl���՜i����vH���}B���[JU��)*6�mU�E��+��eEQ+b���\�¥1+[�KZ�Q-�(�m*V���L�.ڢ�r�,�(���QU���AH���F
��Eƪ*�1`**�̥U�l
��bĭƮY+`Ԩ���ŉmlVF"*,X�%�e�QVe
��5ڪ+R,��5(�
�U��A�
��ª"(Uq�1�2���UA�֬�`��\�T�n%�"����UE�W�̘�q�0\�Ab���*���P[[m�(�\A�+�EE��	�����%`�-��9s,"�-�-"�m(T؈V�+1�@��m�\���R,F�(�Y�f8��*"�"1j�j�eJ�+2ز҆*
��V�,E,mh�Ĭ1�L��,�CcZ,��i(�[�L*�*������:^o\�Þ}������=��٦k�H�=v�n�i�3�o`�W�F]6��l|��o�Yt��3�wSyy���q��^��:��N�a���k��"���Xv
�u+��7�D�����;ltXWI�(,Ѯ�z����ttz�B�#��h1�m�r�"��T)r�f)����]%�$U/��4*3+�o�qI�W@��`1�է�C[�C1�g���Djμ�ܬ�^ƍ�'�*%�&.'a��&�a��Y�//�+�1^%f�&5S��-�[�^�lw���|���U	�ҙ��͘�ta�Z�3�53ܽi����u�s�T�G��M��vWX�\��+G�5/�b\ܬz�b��sd���V��Mr��<�T�X(�b�0�F�u�f5����Z���S�E.
���W[�J�n�H��	�BBl�7��%ᄺ�^�7��*�U	��]�l�l�-`�:���f��E�`�f��]��
������1r�\��>�|���w%�X���s�l�7�mJ��_��,d����0�qU��(��M����\���T�W�����7���/:Ӓ��L����a�+z3R�slv���G����̼5o�ےL�U�+K�f����. r@B�����%�aG��D�9WLWu�ҵ��v�)ՆouETZ�<��SOqޅݝ]�Ͼ����
��5=�ʌI�;Dn%�jZ�o���;U������U�֮����&�A� �$}����T�{,_���@QN^�X�m��"��ds�H\;�<Y"zD�Vs�y�u����Ŵ�.���Z ��o6JG|�n8z�= �[��<s�b��P殬�;�I��37k&���DX�������X5��59������аG&��e�^@�N3!��V�op�ó\q�A�]9*�Dג��>�Rк��Y��\���R*Z%�(rq���fMb��^N��i��,]�{T�����5	P� A�;��`p۹U�Ц3��|���=�1���r�Y*wEND�S
�B팓K��G��3��*#7��N����:�F̸���q��6��l9]�����~�R���}�g���%��r��(l���� ��m�ʔ�ߣy�P1m�I�-�-���� ���b=��5!�qϮ.�c=���juB�(��?m��:o��U���]�k��tF#$�V���gzpޚ�K)� 	���W���b���:�ן^�%Zę=V���A�l6�4e�`9|�i���T�o7���R�NCs�Z�OlGEh2�@�C���}���	k�";-�TT�2n^� �D�RIӧ*���YjE��x�?T�n޵�(AS�X�>+��ˋ���x{+m�q7��bog��]��Q�]
;�����:^�����h�v4.Y�T���P�ؙj�D��!N7x�E^jFy	~Vaɘ�tԈO[��4
UA��1�6`��%{u��[���I��
��Y���� Y޿�f{*!��0�t��Y�µ��8��\���M�%x��h-���,q4Y���l�(�/�/���T�f��Փ����㛭ן83Wy��Dh��V6|��U��qQ��x0*���K���[�$��e�U��//U��y^ �w�]%xkE��|C�t{�RJ��cb�źP�<<¯LN�{fW`���} 9ф���z[m��0a��҉[�%A�H�L
��:3���]��Qd��<7ԗ;q�9)�;/��P�8ӽ�ú���#(V!\&c��D�1�9�t��qQN~�k&{��6��hՕC�)Lg�us���&y1a���~�$B�j�B�A�?�����n81�y�����'z���H�Iт�,�`��!����j������j�%7}�Wn;fx	�Þʙ8Ѕ+�A�Ҍ9Z�nǶoJ�j.�0�N���2�����N�_n�9�*��̾��S~DZ�e�c������oGsr�Z�,��T�c��jF��:�*�9-��oΡΗfg֧N.���r��\��Ì� ���Rw)���^�b��	ձ%��ۚV�_���Lu�{'/J|o�Lv���-EV"F�F��.:�x>��JD�����7V���S@�Ǭ==�ydOpc�NvK�\���3�M:�W��%o���r�����M�K;5r���S.;�Q�c�Ku�h�Aۧ(�C�Uxi��R�$��-5��^��i[�����9Q��.w<-u9������!�ޘW�����v�3)���n-���mD��-��x�.t�7�*\^ǃ��^`�]��G�ԇ<lk���yRW/js=�8���{�7K]Yva��������R�.��BV��=t�6�������,��or=����8Y�1Ғ�z%�~�I�*�b�|�1��t��SUVsF�l�s�ɺKq�:c6���b(Ɋ��+������J~`/�� �p?§��Q�W�YrΡ1�6�ͭ��.�=��i���ySǔ���©��;�%^��ֲ��7����7��9���vN��t�̱j� �����\��_7K��`\�,��a�̝��R��Z��xUN9��7sr�/uwH_O�U}�����,!����Uӷ�Pa�PzkZT0�&��|:�:;��t���������u73[۴���ڎ����S�ɡ�*�'՞���ˢ�XD��@~
y�L�	#�s�W"�y��*�Hn�	wNbߵ��{\�����
�C�J�DµN3vy�m��[S�c���=f:T�ZE����vx#0c�Y��v��y�Iä_�U@D�����b㹀A� �� �{Om������a_�*6^�a�������PpDŒQL�����kE^����N�0㹡4���h鎐m��bD!w�R�l�ݻb^�c�J�j��~�&�o���]��EÙ$�Ď�W��Ma���1�p�X�2@z��(�L]-X4t�uP�r��'b[b�u��&����<��r��c�Ԥ���˯��F�A�qL�V7���4��:�	�ҙ��'чq�FZ"V��U<L��^7j�U�:��m��ڂ�F�m�*r_B��jJ֬M����Yx撣#���w�	�e|C�ã::�q��9�T���Od�/dqL�"�+��G)��;�+v�+V����s����s%��v=��']s�Ku��[�$&n�zJ�!�&�e 溰0����m����o�_yΥζ9�;���U|�2?^��:N4������F�3��[F2k�S9�UL�?�ll�t����%7Y�g6�*b2QW���Շ��R�V&��#����\U)�[�&�8���Z&�Td�J]�Q�%�#�J>�8z�������XB�1�+&x�\�S�
���������[�en$���ѳ2�iJ�Y�L�ά_^�E��aj�)ȵ!���[,qT��͌���P��B%��z�b�L����|�,+�=������J���� E<���x���Vw�5�*ֵ�!ãIu{K��-�\u�����F(�'n��S��纛��|Oo�\�˖Iʵ!5��"��:�8d��;�3��8��ܨS��j��v�6����X�y�o�������|E
��B���'�P���{�w�RY�'$��}���noqR��h�a])D���0R���@���:�t��^5Ws<|�8��F��uY�=z��{=b*o�� ø�F�5	P��NQ�'�bd��
@l��'.�y�e�� �n�9guЩA�p��7�6�C@���i��N�-�M~+��5zeywv;�Q�67��F�<�]��gN�{p�M���`y���;�J���5p���TU2�m�u�C҆���|{)7*Fd��(${��s
���q��t�Ϫ���wۉ<f�J������1t�Y�d�QS�%1H�B=d榺SAh�����u���*��zj-U�9���͡,�Õq.�7�-><�M�ֺt�k8E��8/��ȷ���NI�6�o�T�.���([njL�Kr�Í��Grd���}an��XB�B�;]g�5�xeU��Կ9��]�����ʍ%/2e�)��G6s�x���z%��Z��:�Uf豴�v)N1�)7��j;	������u(�-�i���>�w^�I[L���y���ױ^J[�	�m�t�sυ��\�qf�%�D����%���HN{��0�3|�R"��w�6,l�#A������:�]��ܽ����T�Xd��Q[=x6[�l�w���#�Gy�u�����/�r瓌u�(.[!�J�~���Ⅴ.J$W�X��'_�,|XVʖ��(:�����tL$����Y�E����ۼ�ު���I!�H��F�Ti���XohK�/���s�^�t�s�����Ξ����vo{�TMD�ܥ@Kzҡ	�`��#����[ީ����z1Z�_RZ��`�r��
��T--�Ϗd��.�"%��V�V��9�\�ݲ��ݎxD9Ys�[���ǜw�!�=���8k�E͒�\ءgw���~�{� >������k�G�r�_���]��#�:�t~�$��MV=����|<�����i'<lv��_�t��|qQ�����H��%FH�L_��o�܋�<xڍrp���[�$�莱2����:LZj�It�������Z�[4x�>�?hi��ǎ�כ�����l��zz��e�j��ћι��/׳����6!�9r\9J��.�3b��;ϔ��������9�Dc���a����ҩ���-�b�=jvK-�m�C�w�����z&�f
H��o������!w��J`���R���,�����W�h����	�
���GG�u�]{H��ުsưROobdkr{:[ݱKْu	��<rUr����֍�M@T��S?>�]�X�Kw4����$���3�K���0���)���.Py�g=}�h�I���Eed��Wbe�IL�/1��z�<{�Fm�#:�e�\�d�-�30|����;za^��c����h����[����1��i�^\G;7�����F�%tO����oe
�a_E���y'G����"��[�3n5�gQ�\��C���
�Pٲ�f,��.�"�t�,��HI�*^���+��u$w<���1�[мs�R�.5��������'����P�j�~���τ���=W[N^`��X�{Q�.!��ю�;�f�#�V>2��*�-�їqU��w_�b,Ø��J����߇׶T�D�*\�ν�����x��%��+�ٺ�i�7��c�t�/�h����wx	�i�N<�<;>��-j�2V�=Xӝc���.:����m�1�T�ܠ�f�Ԗ�/ -�� 5��/e_�E�};�]Sw���'�w�W��%�:��A�j�tL�gC�$l�m�tY���5$�n���42��/UC��	�)m���P�6�A[��S�t��U����RÆ`I ���9f"�v*Bt�t��d�`���ȇ��&�T3�1�Vu�����L��{x�/.�揎pxfKuo"**9�*m*x:����<�̌�v��t�Ҏ�$�%�v�jp�Y�˝{d\@ Ь��J��g��ڬ��f5+��3x!4Eu�؞''&���-���%J��;&�90�hM7A }U��1��\�� ~7y�c���|�̺,�N-�-+.�5��w��}@Ừq���Tkv�����*�<6rS>K`U�������\MY��M41^�̅�}J`�Qi�]'nַE�y���ڳGsX�����1ku&��<��!�/�i� Y��:�Wt���ވ5��=|Ϊ�3��n۸���c&�Y���vU�p}%{Ȏ�|tR�X���ҫG.ՒjδyzV�C\o���3@�0�*&ۡ1�%��Y��%I���P�X����m�9��~�u�8�ګ��2�|�.����4&Kt�g��DT2�c���
���|��h��e�F//��PxaCP첸�����p�J�"x�l��������a���԰�K*�;����4�:��ө�%p�ȶ��#��x��4}��֤�� %g-k%��%V�ok�jŌ�dґ<M��K�<|2�2�oث�-�iv3hm-�Eo!�J�;Ǉ���,��V�\:Zd���`.�0;�cw/s�f���� �l]!/t�����Y�y�Z2\��>��Ր��ي�ha��v��,Q���'Va٧쮉��	�F(���z}\�\<��l�M>�ɀhh�W�1����VwP�����r>t�������*P�9x�X�m��"�+�G8��{ц�{��ʸ.�U��3���ʠhKt˫�u��u��P'b�V$�pب�R�T%��_���F�Z�S0$��A�_М�EL]���S�/C���Ԙ�e Wwe^u`¯�	j�Z��u�uG��ڎ�e���E��N�ҹ��n�u�}};��e3+:������\c��ҕ5"��zW:&�V�F�Bn���fP���o�3�]>[K�nj�ui�,gE{
��s�t�����/��j�B��i��9���5H�:�T՚�ѐ�	�\�:����u�*#12�T޷hk�����6��v��F�9´�>�X�va�{���HU93Y`��(�9h|�Υ���ҟq�8�!x���[M
��HppDm���^*,��ܲ�;ѥs�̗����c��n��'��ڈ0P��S+�E;�������u��{D��'��ɍ���)VlRkM�m�M��IJ�%��F곤�Tx��5�츯Hp5y*A�X�%Eu���Cv�-�o�{}|u%��uN�颛c8��b>k280��ONh�����<��$����J��r����&k}���˾w��m@h��q�+���V�Y�z`�L���4�B_RL/��Ū(Ю�J��#Ou�E��X=���w���\z���8���m�;�P�RL�V�j�ҷ]���\��c�}y����L���]�M$�s���*�J�l�Pe��n�ѫL�u-T��tBDK«z�)J��3�Ό[+���F�k&'Ҳ�T4��N�Q�zse��<�[1X�X^ͪ;ݕ���2v0f��u���I#��Y ���Bq����:� 3����Ԡ*5���% �7C�;[C	ٸ���Lw�v��l�oR�XT�)���U�O��j�<hz�5��2��91u�X:���gb�;5���EZf��Ų&�eQT�.�(о:+F�o�U�"jJ�E���wz4J�B=<�᝴�s�.�.�7�vȭ����֣5��[ZM�w���ʬng>)ҩ��Rw*���QJ_����Z����oV޵�l�,������@ފ}�����c���2���ڕ�x8���e���)1��k;���f�
R�m�O7�T��Sl}[a�+4vS;K)TP8p�<>���e�ӂ�-�!�w G�ɡüo�A����7M���kx�Ud[�E%�e]�fIL
|�8og>㯅2Fޫ����u�P3�垉vq��t��d.�U�Z,�G��_�4&r�ܣpc�H�r�3�}Z��ڡ�$\������ʺ�Pm��f_ǜ���Z�ۃ�����O�d҃y-<�^s��]��$��R.��x����]�7{�� �!@�*
	��U�%�YCN��T��6-[�x���(��d�ęVY�2�3���J��Z��T�6�J�P�\��
�1	��. �T-��-��P�
J�1��PĨ+0T�S*E�11��J�q.5-je,@PR��E�[L�ER�1
5�����V`��
V��m�V,R�8�V�**$U�F�f5FAk,V
�0Ĩ�m�*�e�YX��AJ��T+-��Y1�ER�YLp�*�Pm
!Fc�E�¸0++!S��
1��dʱ`�+
�e�Aʵ����V\�Tĸ�*ũ
�m.	f3-��3
�dL��eK�*��4�1�Xc1 �J��-̊T�K%ap�⹙���8���+1*����2V��H��
�
�VB�lQd�XJŊ,0�bU��	PĘ"��YRb���*�C\f5c
�PU�&!��*�Y����q1[0}wwU�7:J3]�1�D�Y��u�����������D(=��JN*�`Z���ҙ�����mN��l���9�����^.6x{g�9 �3����*s%�r�L��p��c���מ`V���HrT&u6��쨦o'ٚ��V��8��+"vO���h'"D9�6x��59�������m�A�/�*Ks��|�{�+B�Y룧�lq])D�J� �R���@��c�NV�Aef�i���6���qZ\����A��p�;Sl2��B1�dJ@JVvz�w2��dZ:�:E&��b�^;�E�hj�L\R��d�T�y�T�I��#���"NP��7�v�J,��=XltK��)��]w#�J�Dy�l9W�2܅�{��ݽ�59Tt�����p�����K����;��9�����x��1{��[njO���k�΋�kr�vӾx�\o)@q���\�J��kέe�J��^qp���w��Q}���V�`��TFI�5������á�V��xe*aQ,OB�_����:��xx��eS��=��7�r.�)�}��rF��J�V���߬��N�74~�w�M�����Q��8u��ةW�`:V�sc��x.��]V[��F���\z�Ϋ��j/)��)cܷ��ngJ6�c7Ǩi�ξ�C����9B�rp����=�٬�l`��v�e�ث��L��!�Q�5�'akki���|P�
���q�?�U}_V�w��o�9����zD��o{y�L�_2Ԉ���p�4�X@0��F{� �S�}|�ޚ)�,yK���`�L��R�ws|�;_�gta��x�˭��]4���7C�`���6e
����l��ŏ�"�g&_8����ۣ�E:���_V�?�_���J243�~��t���]J4���8�Xw�K���w.�H��}��Cz͏^�]�W�zJ���aLOKaUT3��Z{�[Y�mNjs��7�Xz�Mx�*��T�~np�^aVrDL�GSGx�Tx{��Mm�3E�9�;��Y���36#�Ue�Ȕ�I�M^I�eM�����g�\H��1�9��K$�v� j�_�)�6ˠ�Ә�:�������qm�����
�py�l׻}�{�sy��(VA��)���9q��1�k ;���=�ڿxk[;$��F����wMLÚ�����>��3~&��69�]ƵqRS�b�3�v ����Acq�k�6�]-�ۙˏ�mk�W���v�sz�SN��hJ��ݡ�2�gfuv���@:<��:���U�gIoy�1�Y���q6���Т��חaEת�WqMw�t��an��@6��BK����䓜��}U_U�m���a�9?�M)ؿ*s��K�Y4&�}�TP�tk�&#���J��\��4��V�o=��r�>���I���G�J�^�~	�٨
�]
b'���k�P5\�kw��+(����XS}�̮qQ[	��r��3��b6�� �U2�p�+�3��w?F|���-�_����6sC���6��uF�+�̘[Nf`��=�1ѧjv��(0��ro���-�\�͠�A��;���v�c��]Vǃӗ�'g�=����LN�N}w��;2���B_��K�t��ˎ�RyM�	CFx���K��}r��R�.)��,��龺j���8�%�ľp"*V���"�� ���x1$��P5�#��Z�Jj��C*�:�*_���\�0�,�&�㴒�����������[�~�o�[7��eL��kh0e��w�UӸ����I�j�tT���jͰ��gZm�+poIg���t�Ѯ�෴&�[}'CB���+d�35|*c'��3��i��;Z�x/uw�^9+���g������;��@�4���r�V�D4��gC"Ⱥ��(g^��SUm��&�U嫞V���祀�Z ��pk�����!����;��\��k#Q�nuđ4�>����G����b�z�^�}E\)��o����#����:�qKt��? �+��WԈ��L�������<��y��o!� VKJ�T���	����K�ʡ�1�7�9�uϬ�J��z0<1�*��?�{��}W[H�i���=}�b���������� ���*�z��~���f5+��W73�I��N�������5�T���t�d��ra�К��@_���{�����2'7���g-u9بp����F9�&2o�n�
�h0��� Е��N�b��K��^��}�';/�̱��Hr� ���4�.v%D�t&2$���&�*v$=h.���Z�<��@��q���̨����f���h���Ɇ�LɈ���h�Pb�ڨч_N��f�6pO���{h���V�Oh���v;,�.&��j��X/v,�'/-7Ե�	�V���GX%eE���n).�b���w
r6�(��1�����C�GA���ךn~��zm<�D�[�)��{F`0��z*��Ý��\O���~���K8�T�ս́g1uW_M+�ي��%4y��}QVݞ��2�Fe��ұ�9���^=�����է\��}C��pw�<k�I4�"�����یv�&;f���Kp "ӇuM���0<����%Vv`�$�u���0�ׇc�陆q�����n�<̹é�a���\���������-��*�L�dQ��sE;K��ιٖr)h��#
fN*R�f�t�/K���^�J3��`��.�	�I\R���<�X�].�=�x��������y�)`��]4�[�r�ʗ޲�����6ĝ�:{��ʗ�S�F���I�(�QN^�"Yu�7�@}�rxc�K�M�	]�:����ֶF�C�!8+�"�Ky�)E��%LV��w3�O�݊�m^'{Ք�Ff�T��/z��ѯ�# @�W���Th�� �S���Kl���&+K��3^��UU��[*vv�o.6C���,ߙ� �!])D��U�b�K@D��r�W����b�K(�G8���:�-�;9798/�ӱ7� ���aY^J��#��I�MV<�	r�5
�%��F}B'X���1t�Y,�;���"T��F*d�)5��;hWn��y'�@~ܚ�>Aʻ%�z��D)�%A]_�hK0T1HL�#�O֮;�w�������z��y��ڴe�[�4��ʟu��&���t,�×�17�f�M�vb�Ρ-r�',��"�WaQ¡8��ONм[JM{n%�����2�U��Y�j'�{�{8�ֹ2�u��z�*Z�v�Z�аJ{:�`���It�;��oA�y��ą`r ��m.���{ƙ���s����<k=��ޟ[��tx�h-=�x\K��Z9�jb�I�#*f���])>�f��4�_q�`�6ۛ�X�w_87���JQ�N���uxX�ɏ�P����O�x̋�F�F�NuU8\���*�����Q7�u��Tb�x�8l����co��)�,��x���+�I�rN���lۼ��,�':��N�c7�nD[��lE��F��UڡX!�U��f�Oh?PɂbL`�'���S����
6ʖ��;Σ�Cn��˄*q���wS�)�vZY2�qh��+��m�*��m
++���E)B�T��K���]��s[Y�}�Q7I\r���,*z⬉靐�RO���-�*AU�J{����u�k E� �"7g2(*^�aM�*�5�{7�V�@�:8���*�{�@���%ws�G��]�s�Q���k�M�P�R�]�paL:���5�BT)��G�u�`���zGVTз��Y�ɦK��i�.(��̴*R��z���R����o)q�,�m;�*!FNּ9��#u���_�e�,�w2�g]�<'j툶��yq�m���k^Jww�j�v�)N�6v+����(̜{�[l���U���'	�;+����>�C��^Z8+���V�hM��곊(Į|{zR�@�q�J���G��Pw���@MN�r�7-:��ȶ��k���W���-�{�3'�C�]/U�*p<L�㲒�k�>������;��A��r[���1&��U��*ga�G�hǱ�J� V�8�w�7ݦ�Ct��j���]����p�{\�o,��]-9�;��vH�a�}��GG��V`c��>�|53�5֎w!T�%)��(	Ҙ��P3�Tx����7�>��l�}�
�X�$��om���85��/���If����p�^s�R���(:�W�	���U�Z#��=;=����ozz�)�\b��
�Q��9�vq�'�d��̵��fx{db�`�uYY(��M�H����uL�A໦cd�<��p����������gf���Nb�7�r����B�Q�8C%V;hp�^�<O��^u��u<���t�t���JQh(�������V���8{�~�P�J4�����4��� �&�z{�]�U��j�ڒ|~ȷ�7U7f��ݫ
<��y�ܜ�>��-y��@�t�$(��m>h5��K�(��.�]`x9
�/>3lK�o*R4��������y����MU��y�����1�j�#�,;��}>K��J�Q���j��#x��U*O�w��O�e��uy��/~n�W:L:Yh��K�*�Z=���ОV�f]��7{�. M o��������d��^��Zҡ����@H��v)�� r��]
�w�����'�a��4R��9
��sq�+d�3Q�=�.J�5��'�ΒG{Eh�<L��&�OJKG9��BR�?0����*���>{8m��U�R[�.��elw���DB��4)������-��9�;I��r�Y��zvsn3Y�|1������[
j��2���� 4+�J����u��`�ܳ=:[��+����;z��P����n���:s��9�כ��>���^��yʗZ,��WȋҀ�:����>����lAǦ݅+�#:�3���DIU^�#��)�KK�#��;��eH����(���7�b�y�ބ�)��m���ȅd�������6�����xqQ��EF�Ot1��C�0<��0�JɐU�91�U�Z5��)v�������B�*���VzO�QGFV�qXk��D���МIڝSh��c�ne�n�p����t9]���U�^��`��W<닑���>�]�,߾t�jQ��.�"wCb������U	��,k�@h�U
���[�*q�.�u�p��l��b�(����0����WU��y�K2������P�@�����QG^�����.u�7n�Nm�XP6mn2�(��N\f�q�=r{��5���GYN��0���pxq�^�g[j���yV��.!�����|�N�Q/ݴ�_��LZ.�7aI��\������.[-�w��.���Ky��T�Hw�f��Erx�9�1�K�Y�y�Z3���Ȯ�yd1���4��wn<�K\R�ً��(Ymt��e\M�L	�QM�p�������!K��C��T@x�&=�w}�,x�a�l*���H��X��xq.�S���ĳlơwzhNe��ܑZM���(�� Ok$OLĸ�g�dVi��zJQo�	X`��%痽/�Q��-����y��e��=.��td`u\�Os>"P5�(V��o��޳�_�PG��2����G��1S�3�i@8�k,��&�K]0���.�Z�ĩ��VoM�v�*<�u�,����V��y#t)1����ly.2������g\2�S_]�֟1r�g���}'\
◙M�6p��Uy��]��Et�}[!���r���u;�V�O)�Y�f8����+�^J� �)h�
�e�62dH�FY��)��r������}t����vrm'�t�EK�A���&��T��u��5$���d�s������w�!�k����Ju�ꊜ�0Ø�9�nQ�/O[�kd.�1�22M*��?���U1L5�����	r�r�%�Bg���z�Ou�}k�^*7�$���V�� 
��Խe���jlA�Y��o*S~�w8�S�7:�^��{��G���I�4��s�B��k�^��Mp�2���_��,mR���z��n��	#�pb�'8A�xa��0:ɏ�U*ad�=(��B�B��G]f�^�L�Z'�M�=<㰙q7�u�9�1�Y@'��t�C���k�0�5�F��Wư+��m�#���=S^�U�K��E�u�]��\�e�o[��g&�qWC��ό�#�YG�Zp��#��:*ʦ�'��:���m�.�ws~�Q�#c�;L���13��"�nv�:�+�����j�X��F1��.r΢��q��ug7���c�on�Sp��{��Fz�zApu��s�����wtt�9ǩp�\�#�B�������V����غ�=߭��
��`�����2�{Oi[��|�ܦ&:gA��7,�ZP3o��"��b�pֳ/����Y�];ޡ��fa�S�)]m��]�\�Z�`�[W׹b���Ch��&'�w�����z�DQ/ߣ}H;�й7�Uau�m���On��v�X�eQ��a�L��n��FeoJ�ͭ��+E�<��s;wV�#Z�L�2vm�h7`Ej�Ѓ�G+E���8p�@��X��a�i_�q��E��C���2h��f����thn5�j�Ւ%@VQMRW�gRĪ;͜U�I�]�f��0�<��7t��g2h������p85{Q�ޛ���n�JU�T����1��w4��f����e^�عb��/xF�C��$���ՊZ )�&�!"l�ܸ�]��fN�ͦ)ݩ��S��ΨJ�:�X�._!�P�U�]�I�:/B��:�V��sr�7ǒ�rh}�D;�e`��>�/T:���]H��!}7�
�Þu083�6��uj�#G��b��5}�9��)��}��dśmV���'[;�����]zt�@[s���V�c��*cu��Zmn�,T�l6�BV��Y�֚�F�*>%Kz�e�t�7��{s}�뀴�mIW+��f�Z���n���{8��u[���Yf�N��=P�Z���|B�r�%,|�5�l���듹�Vǎ5D_K�k8f�ΛÔFA4E[��vG���q�����;-�6�;n1-JM�pY�D�Q�.��yv�Q�q�2	(=z�u�����7��g��d���jf����I��,&��׽EN�\uu��%6N:�vF�VY#C����6�Ri��s�I��dh�0;1s;g�����\���%��0�wl�N��3yl�e��u���k�{�&�����t^��6���kJR���c��l��n�n��`��9ۋ�v�� e'���(N�I�0Q��u؈�7�\�
ִ��m�5̙ہ�|"ոz-�V��,E�W�k=)]�f�v��q��:Z�*�C#	�Vo�ɑ�E�S�Ƕ�ʬAt΅�7�N،[@��-��9H�5Uݞ}����`x��3f�T�<b�Q2���C��=8���e=9JS+�d�����y������X������|1+�y�*��4�V����Ow&��\�g|�3Y�u܊%��k6�D���v��tIv*U�U�8d4wע���K֎Y���m�L�����sl���tGo5�Y�X������O�������v5�Y5pvr�[�$��6��\��[��o�ׅ�8�-���Pr�b1J��@�Y0C
�b°rʊ&2�[d��Y%d��%`)���V1�����ԣ$Y*)*d��k��Z��Ȣ��&$1 �娡+!U�UfZEL��Hb�	��LI*6�-aX*�10d�\�V.%E�e��B��e���+3-b�P�b,kJ5�eE�+�����LLB�)��fYX����A�d�L(VLAm�f-��(�0D�
°��mJ��Im\aU2�a+
��L���&)1+�&Z"�X��@���[1���P��Y
�T3. �Wm1�3,�P�1�f0%�nX�-�﨏�A
�o'b�1��r�Ĭa�Aۊ
\���l�5s��յ�^���Y�woFޫT&�1�z��`n�s���Z\���Y��f{��rp�
��Xt>��ve���,q4Q���>,"�Kэ�ĭ���1��\��r��d�*F��j����������Hy�H�wC�S_��դ8N�;h�w��G�x'��*^�<o�[5��l�#���x�@�����xҭW��9��&Z0����q��z2!�	���*_�7é��H�ޡ*%�R%w�V����P��T,�ۻ�B�����)�M���=�dp��틞�o(�YWE`ē\����$�NX����Aڥ1�u�w�~��\��w�i2Bn���<z���r�u츚��WQ105�0c��O���9��C�jU/�x��5�{�ݲ��= =�Dؗ������ތ
T�ר�-��������!l;��S9�����۫���9/v���J��sJv.9�^��	]aU�����ypzǽ;o�ȼ+h)��M�o;� �Jb�'v�m�m�S���*���L���~�/<�ʶ�rڑ�%���T�.�m�~O+׾�R=����=9�V�M��q��ky��}o*SMGI�l��/x�t3A�+">u.x�FF�^i�H�m�������5�g�1f`(Ni�z�5�}nT��ByK.���(�4v;g��Z�e�cޝ��}8Zp�T��#��/M���!��32|���)��� �Py��s���J*nl�����V6wp!ze&+hL��]�;�o�i�kU`����b��{��]�/(3f�'2a�����s��� G����:4c>��=ZՏo/04��պM��>�߉9�`�=��jܾ�KBc�R^�:���yM�4g�����鮬�������o+�O��=*U��y�V]8�`�^�LtK�K����αU�j����k;��u�Q/2��
���"˛�e`��m�0�0�-����Myv�&�9����j`~z�T�h�@{��؏���j�Wi��������e[Ԏ�M�ϵ��� 6\Y.�S�g����?}�	�w�_���F?{&�|��3�l��␛mn���/WNƿ
���
$�a]WJ7�X��L��s���[���Qȱ�>S6�2�yz���tsf��g�"}�`��	�>�*U�GZ8:�����RT\��#BA������rV�>�h���a��<)�&dv�CWqD6�c�P
�W�T
޻�-�Vgb���8*�K��S�q
�d�i��
��MWFv�]]���؋��@�(�p���/4̼}-�8�FhulN�����ҹ�&��^�}!}2�u�9��3�{w6�i����F���wv*��wB��/�k�S��G�vC#�!�j:qY�����.������zy��xO�,Jb�rh�x}y�S���w�ھ��vU��o3�J�
\���,�d�M�tȵP�"� s��a܇��ﰤ�G!�wC�ml���c7�b����
\�N��T7Bc"T�6Ӯ�+(Ν�h�ހ��Gz��r�� xV�Sk�+N��[c���Ԃ���U	�CX\���)F2�yL������A,�9�E�
��۞�(�>�S�0=G�í߯N��^S喼�<��G����G8��7��ω��JʋÉ�/>K��D�i�ܒ�!�=Y=�m�V�$⯵
�Ѧ�4?Jce�y�>�\35V�J�Gǥ%~2%�	� �/n�	�]p����sG��7�����Lb.�;<L<e�0��[Cn������$p9~0�^��EN�S�bљf�bn1s2qR�h�p�eh�K�;"���ż����^S��ϔ�ƥ��>M�s~;�݌��·Bܚ��O�"x<b׆WF�k����EF,�����W7{�=�4^z߽�*�|^����Q4���ɒS��*fm�&��]�E�.���v�=��yz����dv�z��B�{:v"ɷ�܎��G�B�)ih�=),����]�f�E6���G7���gkkg�V�Z�=|�]u�\o��Y����N��\�C���T�ʞb�r���*�ʖz�v:��9!n�"��/G8��wDk�6F�C� �]���.�礥>[��˙ê�M
�F�SM�n�t���n@)|��)	�W������@{��~��^���ù��C�s|�_%��UT/������'��B��W�c�sm���Ғ��MBT^ɜ�R���@]S�:��]��X�X�"�����Nn��������������ws�o0w��v"0���s�߆ި7��'X�HsN˕��S�@�����RߥH���}ާ�|W'u��(S�&���<�y�o�T�0���z)��	d6�k+�=�����ðL���#��u!Z1�kn����G��^�:�/����ˮ�ފ(����h��>�-�-���H�:$��à��Y
tç�:x�:@�1S�݉�R�Zh:������F���K�A� �&�(ubxn���Ѳ�����g;�:�q��+��o1��푒���1VV���h$�ع���m��7���:�+%.�Ω��C:���r�S3��;�s���/U9�-�zI��\jf8�*+��7�)���'S�X�`����ݧ���ݑ�z�9��ܭ�E<�;\�� ���`�$/t���@[��:r!�l��.Qu��Ҩ�+�3�z*�_	���F"��1���u�HM�Y�lNDu�i�L^G2Ԉ���padݻՊC��9#���[�"�.(l�0�Nn�9Q9;)��l����̙�"o/���|7�	ծʣu�S�f�)��@���<�	�����\�tR�6FՍi�ʡu��2��J���/:�>��Z3�dh_y�B��X"�ΏO��؈�y�x�[��J�BT� �9�7�,�[����g�(h��n?\� x_�[�{�pVวXL�>�w�\OM��>z
��\|}�����/dB{�N(XM�'S�����R��;��Q�Ү2�A(򮆧ܣ���D�s�����[A�$�"�-����r�t�S�"j����R����|Uq˘�2)�������uy�R%i{6��a�ڥ;'U��['9��.�V���&A���:��pЏ:�V�h�`��c���[��-̾[A�{�əв͞�m B��>���7vd�ǖ�T��g;�\Y��?	珺tٔ2@p���8��$� �����zN뱅vN�Ew���!F�y�B�n�Ĵwî�O_S�罎�1�j&D�I띮��ֺ�r��o��xD�/~�
T�I�eR;���
�c�����g�2��Bqj#�n�/�ձ%���\2���?FǄ���C�e#���3��cĪi_	7.,^�������w�t�(�v�m�m�S���sp��!��f�uqw%�y��-�Z>�S���|n_{�8�7�̕�Ru�n�A�2v�%�m�'����g8����Na����ʥ�������8��U�Ϸ�ؼ ����{�w��.�-\y�>�^Lu�����2R��<��o�z\��u���&�m�����y���t��p�;p��09����Bc�^�U���g����_lj��s7���v���v6rr��g��e���/[�1�䱟��\n�(:�,8�������QQ�&����|�0�.n:�X1�1�d�O��å�Z><��02ں�u1.I��O��j����t{�Z�+���O��}�#v=s#׃j�n�ob ���6�m�>c�q�~~���%[���}1��>�-�wlS���j�
o��e B�^9���ﴍɹ�{�5/ouvp�U$�yr�z���	��w��`�K}P�"Ut�����6��A��rerT9tO	��6�]Ю�\ɚ
�_��<���Ko��:��ż��]��:��6^��g¦2j D��0:V�b�'OD��N�sw��m�=03Rň�]�0�=�m��Ŀ���U�\��H`���'x;���l�J�J����^��{{��Ɩp[q���0y5�����ïD��@�^  hV�F�o���>��;�&��s�Z�6��T��S�0�o,�Pp6Μ�qNL;�M�@TOtQd�ue�֧ j� �V��h�.��K�N���d�K`P��P�WJ\e�P�M��%�6���$@�i�L�(�oB��Nh�?��~� ����/�TM��LdLi���1��0.�\'��7��5Q�ۄK��1N����j��}�>��@��} Wk ��訲yR{������/��̘�ʺ0�"Ѕt�=����
����`L�#¾u��=�e[qZ�V�����E[W�B��U܇XJ�w�+������D&�����#ӗ;4Ro��\93~Ȋ|_pݫc;�.:���������Gz���^ڬ��x>�H���4��
�}�f���C}��Q^vպ��/�1��Q���W����	�c����QG\2�����:���%�}!-�N/7�����t��aFFٍb屲|����*{�*6vvp�pxq�1x��Q�I��<����FK�J���]0�j�1Ћ���j���A�S�x�'n�C)�mJ��yz��~2�,�N`'���%_:��)|�W�c%˝���k�"����wۓ�K���3�Ь���m��,����q�QO��0֮��x�zQY�6��Ttt�HZ
X44A5
L���*5���R�8����uK;���z���S�0؆����qI.�Or2��YG��̔��Q[2B������B)�x��~ ۶��
N�����4�Ǳ�cP pF|p���:"�;z�:��4�mf��ıs��1ɫ�3�)�Y�f8����h��4r��]pez߳��L�>��_��a_�K��R��S��h98-�v"��df;���C�w�rDl�|���5v�[�boX�4�\u�U��8��O�}k�~;��(�v�8�,�~n�Wv	BLh'�	,!s"�z����bԄ��x5�D�p|֚ulk�`�v%O�e�@6M��w��o�=;�wP��)s��jk�d���}L蚌t%�}J��pK�9��'X�HsN˕��S�#�r�z2�Z��p�k5A���ɇ�
��@^Jk��],߉��5��u݃�&�1-����Û�k73ںY�0_���&�]�C�:��6�j8��<��1�؃k6��V66�:�g��R��1�%q@��50}-������U��a
XC5��zϣ\-�-��_�>^ޞ��;/���TT��Gjf8��Q�N��!N��d���]mְ�A����J2������^7�������D�E2}~qnߪ�?c�ߧ�[L�? ���/�+^Ԧ�*9�h��VK�8F��r�����(N�lJ�0Ӫ���2Ԉl�PEe��M�����C���X���jO�"�\�
�\���D��`_�ʖI�Y��	�nj�\��-*��u�8�t��O�-��S���RE�.���s�����67���:�_ �\���\�P�{U��o��Q����ҩ$<�U��ޒ��>���`$j���u��=X����������ո3�߮�.�자�x�$�ټ]�9}�pko��@ꑹ�@�{yN0����=���Ǫk�׵�jv�/a3�F�͎@n�bt=�gE��O��>�B�򞙬�"T2��/�1�b�yB\��
_���]�׳}%`u]�0�"*]ک�����
x;R r��!����D����":K>�4WB�*_�n)�R#l��M�Unbbw{��J�.B[t'==)��T,��]̡��Ue��JC��Zj�K�RH���S�k�\��M�+}V٠��<\:*\<��g#��=�n��zX��=�F���)���M�Y�ŃG�t��B�
�U���
��|���s���M�9�8�y�k�c���7�)?P��</=�کln��vf|&f;��9�l�S��2�CH�x��?(����^�Ǿsz��I�ulB�d����[�:a�2���&}�j�sY���!�}k[5.��:�N�r����f(��LRd���t�T�e��<҇�w�n�5���%�d
z~A���	s��U6/���\��&c�L7X��s��a�[��ս9W�vx���'P�3���p�(���/.(��e��}��6��uF�>\�e�A%��#��
�����Uq�3+EG�R�0wQLJ��z!������"t�/;��
<*6:�a�9�Z�w\�t��M�k���ۻO$a�+m\�^*h<�V�EsUD��J�0�ft��Un%'2�_V��ו�N�&b�3�Y�鮠8#�!�F�=u�fVE\�+LsL7vᣥ.+�]t�t��U1B��,��9�ǁR���5-'{C�{��*�蚘�Уj��a\��0`o�0;q�=�@2�4��R5���������\����
<���W����=��n��LT!)k���`W�E{f�R��E���n�CW��VK����qѼl��E����w��,V�U�egvwd|����p�K~��'l�(#��Xsk��\�y4�n�ip���u��)T�-Y��.
��!RUǝ[�"ΰ9`�wSO��M^�c3+klf��s�Ӌ�9�ʕ��{ASմ���G�/�Y͛Nq���V�(�=,�pE͑�`ыh��Guc=�R�p��/�7cHv%q(T4�%m�Rd��u-b�T�O��Ź�]Ȱ�+�E�]k}KB����
�	9VN3n��4pV|"�Ў�R�����h����^�y30�[�(V�C�h��k��邱�� �;w��s�\7r�#�cW�16a�w���7��]��:u��\�βQ�&i��t'wP��A _.���06ar�Jeb�+�=��K.���J���WY�le��Y��\ޢ����vҎ]$��R�ڶ����w��q��H�y\iae=9��0۾x� �F5�O$��V��ot��R��H����Z9�pW
�y[�!�Sz����	�5�r^���z�[;v�	[#��kp�,���fw.���H�����+�l-&�hX�q���N���uX�jȩi7��oz�X��#s�v�d-�X���V��M7�g9�},��7غk�5$ց�(k���ұ��b'�'�R&�I�ں��ǌ
a�j����r�D����y�q�ų]�]��}�֠+�=-���d�4����)˶�\ݑ�G/��^Cf�yDf���;Oo�
ҁ7�å��xe�0@6p�u_a�M�Ki��07x5Lu�솾�|{~����{��x��6��u��ʹ,�M�x�u7� �x�Z�S����R�+��Xǫ��D��X��V`����=څ짼�q�5�����D�=�O�v��6�2��EF�5O�3;Z��h����@n�7�l.u��V�ਹ��K��ݯ�X�/#�q�r�>j�EϳK�X�Cm����;�Siɳ��;���o)��/�mA\�U��8c��f�=�9�o����@S��Ig&�]�A��ٻ�f�����k8�s�d�V!�޼�9�>���vN��ֺ\ZT�騜�a�ӫw��h�g��Χ,�T���t�ةZK���;#�>�d�Lǽ3
}3!�1	b1���S��(�1�� �9q��`�V����H6ʓV
UVIm�FUqP-���"(bQ"�-��(�AVEPE��Kl�
�VՔQR
,PX((�T�UJ�$-�bȰP�V�I�3,����1 Z�J� FAeIR,+*�YEbŒ(�X� �q��YDH�H�Kh,X2,1��H���LJ���ŀ���r�,SI(�iUj*����T�iFcr�f8��0��-C-Y�T�mQE
�E-�)�e�%J�+TFZZ�S�s2�J�b �cY��������1��[XҶ�XVHڵ+i�)��z����]�����ڝ�I)�4K6�"aG�K3�ҧ�"|�{\k�z��B�fu5�D�������$�#ї˹ε��π�v�`7U�0��^���Z;fE�Xн)�ѐ�O�c��{ۆp�u�U�5./R9)�WI���֬M�ڌ�>񰾭v��z
���/:��tQ��v�<y��I���b�xs����%��Ȅ���1�j⹧'ݳFPA�).�ٷ�F�|h�=lبL�;TTtI��K*�c��.M�v�ct�ݩu�U�{O������,���W�=K�4�d����\=�
�� �u�Ϸ<^�ez�KG�+�&$��tR�{Lm
~̫"�,�y��K��󻚺E�'X�c��	�)m��1L����Ocs�&t{v��*�EX	���*�Q��*�M�e���9�u����n���fu(}�y�%�7%5̿DB�HХ��]@��F���u����<R{oL�~����r�Q��B���V�zy��u���F��� ���l�p���H���ŒT���*�e�J��f�B�uƶ^ݯt|/�"2*��X�;?b�p̝/sd]n##��w�D���d���t�F�^Y�4�AW�� ������C���{ƣ=��y�s37ڠ��+y��%�H�KMt� k����sމ9GV�X~2]��X�̜�<;��W��.ۚ��g(�$'7{JI	��{�E�@�h0�A��ĈB��)۸Y,�ɸn�B�6�F��o�[���]Փ� b�+�:�5�*t�af�\�o3�.v%D��˃�^Ї�/����^��YCC��7J��'��ۂ�f�B��uy�;�����^�Q�'��N����۾8�n��Vq����O�}�J�f�t�X�f/.0�o4��������K�hݬi@+U����p�����X��0v5|j(넬��:R[�JK��g/���6��U�oI����
3lƱq-�����=§�j6vj4`QwA����w�8�)^����u�.�K �Z�'�h�~�]0��I���.�6[
]�S��FTL�5��,<�˦��e��0f��`.s|���D�u��J]�,�<A��w�����94����J�t�����WgK����6�D�y�҉��L	����50�,.7����W=�F�!O�B����G�_L�"�MC�C��To��~���
P�$r�'�Z��×�\����N�ۭt7]�c6�^aG>�˳*cr�8�XBNqm%��S��t̑K���D��qn�.���)�Y�2y�%��i�StZ-Toh���cR1�a�œE*�օZƮ��s��Y��U�0gbk;���7y��/����L�R�����G��jp�Ü�;�<���K�� �h����I���ZRW�k�:^�g��p���@)�k�3��k��ތ��@/r>#D�[C/�i]���'8VK��Y���W��oFe3�ӑ�`��W�c�sn!��
o7��plL�Tֻa&�P�5�t4 >��P=Y���ç�\R*Z�vrm'�t�EL�C�{����9f�0#�m�5΄�*r�ǉs���������.)�w���OV�<^~~M�Y���o�L�����R�t���I��C����>o�LW��%A]7W���J���^�5��)�Q�>'�	U��D?C�
��nf���xPS�|[����]�'Z���F�
����*Sq��(��ĶI�斁}Nt����$Ge<k1Ƃ��穤'7���F˼�ljDv�c���Q��M˰�E�[�������	�s��7���<����6�V�p��^mۗ��=a��G:邹�����2��8�5�>K�8��}|1<�V��%�Tn�TY��Q��1�Ñ�[ه:��_+'\��G}�H?m��2�w���Lݞ�tW�H!-��uwbד�M�twcݝ�όcip���y��һI;ڨ�fq��`~����g�d�I�gN'�_vvl�;�)�p����WK��J��8p>"�����[L�� ���A�]Ŝ�n�»�\�D>\���p�� X��L`�%�b�(ʉ��L�V�N��Ȩvql����8��s������ц륖���	��q�kMҮ�[���WZSjَ��r^��yO���K��3��G
�����r�EV��v8�����S�N� )�{%e=�����=�.T�e�	l�>d���hҗ��/'���3��{9�#��0 r�0W�\���}Bj<Wl�n�q��U­@x��X�Q-����j�1�#�%�*3�:[P�|�您V#UYx2R6�7'��������+ٱ�¡\&aב"%� �rR�u���<t�1 �w5Vn+�p����^N��s��s��i����H��1&F@㙎�.���1�[�;^�oJ���J�������f����Y�Y�Xۡ��࿇�^<�3�����k���:ǷEҮ�od��=���˞�>�u�⨳ev[@xCN�ԃl�ף��ز����)���+E�����X���Rt�gp��:�r��g4&bnl4��-n�ΡgPAv�+uh�V��6��������p�S�:j��C]N3D��et����A�y���.㛸�0�[�%��{��u�yxc�FǄ���[C���	��/A^���@���g�#cQy�����_P`��wN��N�D�tظ�Nv��q��%'�������!�s�Ĺ��l�>�ͼ��3M9^�� �EEjfHΓٺ{��m�*���� ��/#|%u�g�ja���s��T�`S״P��,G�S��P+ �������G���q�V%�%2����#���>^u����������ʹ6-u��U�͞����&vn�bm�:�7�[��	z)+񒗝a]�n�3C-o�}Ϣ�b�Rt����Fi��*]�%���A��oYs��NJ�K������t�@�����ҧ�!��_T�¯&:wnr:�Z3�Øͪ��uFZ����u·.�RӠN������������p3�o�!�3�&t]r��P��������*W��>�:P�V��O} R�?x�4�Y^@��`,]^�hT�w������ʝݎ�U��8�;��[���qK�~�b�K�������3Y�WW��w:�z��E��W;�qȶQ��cҼ;I{#��ۋ�«/�u*ʽˮ���cb{o�oS��u���ᕂ��O:�Gx;:�=ѯ����v�>�s�
kW�Wp�]A��񼩣.��P&y�$)n
.�M�&^�{�*�+)�sJ�GU���L[��bm�rT[J�K
�;���1��M@	�������Mm���2���?_m�}C�b��Pxc;<����ٞx��y�I1�ˑ�L�̚c����5�h��5���b�,�ռ38nt�:�캃�����˓&�9���jJ��a�r�79���V�6KKµ+��~/ebD!wP���vU;�#".�Q��a���5r�Gpp�)N� ��J�qN�b�V���X;��&B7�K�+lW)�JrĜv�oe���{�({��E]�n�b$�ͣ�.��K�k�+N����<D{�X���d���_f�KR����W�����O�;���|Y�q�X��Y˦�w:7[��*���� ���j_g�+��a3W�*�n�&�X8����!בgDި���Ow��9ڮj�B�Em�9�8�j1�-��1����=�
�`�d��/�֕�x������;˿u������<�#w2�x����P/�m�H��PF��9�_y.��O��9��צ'�ǯw25Т�ueV���T��͠��%��Ա��]\�m�Ej�u���՚��؅�Ctp=�]\鄺�����4�'[ܝ����.�"\0�S����'�^E��R��L\"��ra �ӝ�2lf.�y ¥�l�y��b�/��֓c��^X�fkǢ�x�K���J]�,�>�Ymy�Z�t
{���7If ���=�ͣ3�1H��0�m҉=0&��PmEr�&m���;�!��=�w]q]g���2���Q�4��U��+�#B�]���L����U7Ug��6�k���dS��]bY�f59�\9�Zz���tpR�D设\�^�ŉ�|�Qj�*ch3�wqIZdʗ�̊�}�)	]����#�זfߍ�f�R�P��|,?����
�I�ѐd���:�W�;`�f8�r���2䅷@�}ܘ�<�x���5�0R���@Sw��p�qH�hg��ɿ ���`/)�]mi�ś�*_ ��C0�����J �*r���g��by����`f�ٜ���uvO8��9��Ø�f*�J���Z��|߄���Tcܶ��v�8Ӟ�m�9��{i�^��" N�����}ecV���uĮ�.�,$7��M�k�//GF拶"ձ;B�l]O�.3�#��u�^U��]������eek��3bn=�hPC��'��R��m��Wt��cWen��7��s5*ð�\�(Lߛ�X@���pu�\�Kl�G���\�	�G�y�+�&W���tM9�X
�h�K!D�!`�ԉ�^�6!b�xV]oT�hi��[��F��s��.��Z6�Dr�b/���k���ڋ7�:�3}n�9F������!�S��:ofP���X����xe��^7���m����
�5k(֕e�r���/4�'�;8���{L���]�4�%�;�%	��;-��u�����,F\Y=�>�G,�S��H���p3��꘹�)��0HS62�A���?CճZ���������8֎�D�>f���7],��/�!~*�X�L�^ߌK��"������q�҅�ʖQ/���L�K�W9�J���٧-.9; 9q��wz�&��p.�GLWEB09�R��ĹR�9�xB���ӳ�u���ii��������8�E�Ԓ:|�)��\R�r��z3ϨI]�ҥ�~��΋��ҵ�V"������n6
��^�V�f�8lZ}S�&,��3;�pK)��4��X�7��-Y9��U�ƹ
\�geI��or�7�h�zWX�wv({a�&��qQ{��鳢h*����cXw%I���zT���1;���9��ʃ���*��7G��@����.�5��,~Ue����ۋ��w�q����3�ц���E��D*��2�L¯"DK����*�QJ]�*��1��J#l,��{�md�md�MU����I���:�Uʅ
�đ�wU.��CU,c�v��'�=�9�_���p��k ;��ȕN��6+�:s���1S3Е�x�2�zM��&��F���騵����n�|��IN��Y�d��ѝ��e��;&\���F
쫐�je�uz����*B��a����f�]��
t�0�'��nP��{�ܻ˯[�d�.��<�{n���<f]Ѻ��3��Re_:�SG����7�����6�g�Q�rM��b�(նA�k;���,x�L��mʖP�n[���qUWI|f�3�[s��%+���Ʋ��w��a���F��R`�`*����ps�"q���>��;5C�8�f�F{����|D�ʋ������C��И�I_�ivM�δ�٪�׫֝�񷧘��.l�.ݪ�R��_��ŹZ(�]m򧒮yN�;�z��2������|�Qj]=�q/mi�}�]A�"��Ղ)%�Xհd�/N�yo�O��3��7���D�f�R��.�I�[���
}Q3')��,�:���R�n���e]�N���ʗp�v6T�X=e�nDɹ*��1Nv7};g.͵T�=�:��Z���	�?yp��p�l�|��s<�`r�/n��}��a�y���wd��
₱��Y�I`|bKG��=�����{9/����y�[�r��K�x�?��<tT>D�!����]FUЮ�q���T����̅3x��"�^�6@E %�b�'<�0O�ԷL�
��B�*'I��s����b���ojOcD�JZ����E��[1n5����9i��,*�8��1Q=0�j �)�mE4.�Vv�uú.6�����M��<���LMfǌ���JI�fp9��S3�D�u{�.㹭D�Ӣf\��*ʍ��ԕ�Y��
���daT��nW��즧,}�ܵ.ܫc�!_#ē¶�L)8�l��p+��N���d�M�6n�q����z�>�C�)��k=}�~n��N�b�R���1���\�:�.���rj�.H� Nڻͱ����n��C�����K��vx鈸�\h�H��v�ݦ:lv*�;n��]�t6z�m�ƴ�V@�aѲ�f��7}k���X���{4]6�ш���C�Y+wn�����s��v�"�n>�^�
��th�N�S�:;�u"�cB�%jR��7>
���f�]���!إy� �[U��OG�P[�/�ck&��:�&�휜D�e�F�^0�8t046�3U��)��[�oK�v]	��`U�I{h�$9��ך*�n��}�G}�`]c�d HŪ��W���O�Iϋ�A+�1���8�%��{�`�(d\��WROXV�X��鑫���s9"�9Z��y��u�p����J�c�Է���s��WzyB��|��+ގQ�ΧwDJ[O��;O�P��*�hi�܊Z@_f�N�[�\���3g7�Z��u��o9^��]s9�FcQj]hk.���ޙ{�ʖv�.I:0g^5+G)D��U��Y*N���l8�t�#%� TT1�j:�R���d�+(%�HwA���$d7:�:m��٢������W7�r˗CY[�����+b/��x[K3�W�T���\XѸ��7l�냦��ln���)��y�ᨃ�;�Ҧ���S3."`2�����s�~�c+_PA��tU�>X\�e'k�A�s:ۀ6Vګe��1+3�C�f���'	͖�M+N�v����C/f�ps]ȗ�3�^s=�:�ĳ�C����о=�>r�ȴMӣ�ݘ���tVe'չݙ��5�(X��Hb����*�Ӈ�i�0#,1{r���־�YNQ�,wR��j��|M��H%[у-�	Xu�|��l�S��+,Ɉl��K6n��9�*�rթY�!F�6��o�k�K17�zp	��h#yL����&���mt���眵�3���9�m�X�`ik�݌��7���r����u^<�f�XN���A���5�38VF�U<��jb��tQ4kK������3 fv�ͬ&��Is���ե��ݦZu}�}�}}T����T7S�};�Ě��� �G��䰁v�����$jݛ->Y�ʳl�r�ө��ƖS���M��`���P��Oxs��o�5nQ����SsY��ww�%"82��ۈx{�(X{��[�%�:��כ�FՆ%���^�(���Nvwv��Xf.qu=T���Ds&��;8�7:mw`�]���,5y6�uA�:�L���珹���F�[&�ηڻ����aX]��a��q6�e�F��\� %i��u/yn�C]X��f)�A�:��\��Aԋl�î�lמ��X��en�����"r�lC
�W��:�RR��}�.�fWvL�v_E�wU�'>�"�]ԁg��{�����)�.|��r_m��Z�[��d�b���5����P\q\F��U�+R�m*�kEEm��a��T��P1��E�X���TH���%*c1R��,��E�(�e��[b��ƭ"�EiJ\n)h�`-eDAE��1��R��-!YiAA@R#YYR�Q������`Ғ�B�m�Ԫ!XV(��)RT[j+�QE-��̴+.5FER�H�Q��e+Z2Ue[q��",R��-b ��Q���b[TDU�0�&2���Q��H���ֲ6�(��Ek(�����QV+��؂�V�r��+*�0b#+X,(ʈ��Rr�`���6��T�aRč�F�nf�*"5�m�ZֵQF0<��o����^c�����N���פ>u�Ve�j��{3�#�Nd]�:%���T�ݩ�U���cɹ}��HzJ��;��qBK6�elO�r�1�'�<�Ʌq�@
O@x5R���R�p4|�����,�z�jr)j��Hԃ���U	��)�؈=kx�׏�hB��Ƈ��E����g[���]�w�b�dm��y���ˋ��Z���Nb�sq�u��>�r��X���{pN����v�͂�L��L�#�3�����.~<�{�龊����ϟ[����Ze��9.PЀ�8z�91k��N���	��]�n�\�p��w'$���Wv��u�11�}1U�+��-zU%cО8}�=�;������4�²T�����A�үF���fS��ţ���(	�S= �҉=0'p3S|�u=����5&�A�Pq�]0�>�x�,+�=�:�VG#f�I����P����>��� �j��-�N�/l��.Ý �(�/_-G���s+k�tj�h\;�<Y"zL@٧�I�L�HmsC�9�}��L}�'��"��ɕ?f33

ݔ����j���h�:|�U~�]�<�xIh��Y��F�Ӓ�p��^*����D�L�ǌ`#���
R�a�3�tS��Y;�Knm�3s'�#��q��b8��V�S9�Yy�i���|r�Cץ�z�*�僭���ÙKp"ӝ�*o(X��[�N�<"uu���t�G]�û�j��w`B��[�Ȅ[䪹�9��]�׾����%���yNb�NuR*e�|s.�r�gT��x<h�]���Ip�J�
y�B�.Ǝ�������fr�R�`b%����܄L8<{8��5��6�k+��3C����R���/��Ds� /ǉ��1�����~��')�t=��Wfc�Q��>��r��9)"ǋJH��f�sזG���q��{izR�#e��uq�ƥ�!��tP��nih��ָ���b���!%}�z��[����v^g��+ir�x:��tM9�X7�e�f�Y
%� ާ:|ԩ���̚c������� gu袁"{rZah����x��b/y��8���bv�n%�S�	�� �x^)�F��f����El������TЯ�>��K����[oa�Z��[�մ�\��}x�sԹ��@���@s�o^z�
��,�Yد�YR}cd�7�v[!,v����N�Ԫ�>�f6�JR"����cf��L\`@.(t��1�	lf�t.���v�%ͮt��^��r��'`����膫b���$D٭���m����@BOP)��uƣ1JH�ݮp�^_'�Y����s�rPgv�/9R��2�w^�%o[�����Q7�ԟuz�V�*���ݚVZ+�]�r���j���M!� ��O�>�� ��:�5=�y��qh��FG�`+�)f���b1xr���ݾ��Y}�E-��aS��C�.�T����*f2n���p����.Z�O���~�{�)�P���*L:QQ� ��%�:ؗ'�>n���j�\�g���]Ju�Wݫ�G�
�8�������T��D��/��y�^�/z=�	R1a�ݎ���t	��V�:�O�U���Dw�Gx���y���κ�k��AL��U2ލ�2��y��ߪG
�㓁#�����W�^c�q$u)B��|Uh8}�q\Ǜ���&d�B��/˽0A��(`�_��/�J}�(Wq�B�h^%��v��ɠ��i�j�
�wF�Ӽ=A��c���a�d��zU;0جΜ�52�$�Ϟ��J��pc�ۘ�-�9Uel���8�otSc����sw)��.��V��T�s�;��Y�O������bǫ,"�]G�������G��y�'���K��PTR�J�=�,���ֵ`xɵ�%�T��7� ����x���K�i(�n�U��39>�3ͧ7t�ݓ�(�έ�����WL�X�N����Ds����S������ ��3(�%.��M��9ǲ 	�f�W6L�è[���,��$���u]�NC���g+ڴ`lo�Ba�j�_G�o�����U��f�"z�ۗ�gui��1N嚌�k=�{]W8P=l�7�0>z#|E�S�o����K�L��]u��n	Z������k���v? )����vs&:�C���L�L�F�n����k�t�����6jc�ulx?J���	U��Of:�>"�W�1�|z<��������-��~\a�c�(��n'�Xqq�T�D�*\�	�.cp�M�g_'�'�7ST9t�6�C=Ic=��Q�{J����q񐏓wnsÙZ
q^8Ő��K'v�����AW���J=���RKeө�=�d�_T�R.!m�����[��.V�w�F9�X7z*%� Y>�:P�Eh�l,���$(�wP�����u(�D8�Bh���rCB���wd~���t׀@8�|>�E��~#p�	�)څOd��|oZ�2���{F��f����9�M^I�:Dt'J$D��KE��$�*p�T�}Z��r�Mf�/��%�f��v���GUP�[�M]���,f�r:� �t���T��ٮ=�徠9���bX���iLqG�����9Z��������ÌR��b�9��i�N��[íAy��DH�!�zw^�(7� �u�����PS���ѐ���L��a�x��y���feθ����
h.8���H�L���LϜ��*"����6��>p��]A��;��i�
���x�[噛[;�c�R�>ۚP� 
c�yN�`�H�*��0�[�Dl�^�T��f>x�Jŵݑ�ҠFE�T=\R����	X.)�LP
oӤc��'7^iW�K�^�����U���=
�D�t&2$�����Z ���<��}��&rѸ�H<���+
:Ul�OpV.#y�����F���x. h��:���l�JՖ|�Q��fi�U���x�BsyeGoD�1lf�m��1�
��jLbjĹ2��S��Æ�F0�#�Jıo'�(�X&C}�-q��{���#�3��.[��q2���T�f��R��	��U~l�ۿ n^���c]fz�����6�r6�^�	�L����d�-E��^��#���	������.��ntJǡ���0�����x��&��	&G��>���ե[B{iYJ3�VE�J�����˻d��a!�B����Q^�j�C�֌��-L�՗n,hV>O�U��¬���Y}�p���*wj`��']�Bq<�j�^p�s09��n7�k�����������2�I;�V�C}ꩳMw_���_�Y�9��)F|X���m�E砺��#2-Yw�9^y1 ��o���󀲨.�.`§�!
X6s˦��t灡�'dB�h��{Kuη���_f,.b,{yz{ӸF��v��d��O��c�7�u/q���~l�@0�E��:n�Wgt �[�$Wqo:JR���ea���k��+x�N���M�S�#{k2��uӺ���,{X@_��,�ѭnfW:���{��s�{�V���7`�i�--Ê��i|az未&���5JZꀦ*�0����)>�D��0nS~E����ߠpN�T���*VDM%BP�9F�s5M�}�_]�ky�dk��u�]�(��Ԭ�Y�S��P�؛��3 E�S\�U��s��['-���O[��Lգf\^U�9�+��o�,�+hy> Ox.�%Q��!\�u߻ݖ#2.Zyzy����uDǾ��~{<+cu��L]��am�ߥ��[����:��b�����*�!��Y�*��z|�\zv�*���i�f�H)|}⏣�Y�7��r��_)����=oO�O������<PXwna�g�^��C��v;�p&[�9�T�η�����u�\*�:`�7��o�N=��z�*��|�v�i;��9{n�ފ^yf�:��s�h��'	���1�\.pb�'j$d6�ԫNg3P�v�����K}Z�`u����������4a
M�.Z�v��r#�t����u�ԃ���n(宅�+`[��8x�:ɏ�V&����t�X�����p>I��%��F�:��ݷ8\�Wܪ�1�ijD=l��*�������[���%��1vny��N{� �UFz&��g��T�E���X!y�;�!ţ���~+�m�q��i�Y�۳��:��j`��E8?�F>%���%�s������rw�/"k����O{��3�����l�K�h��qQ�r�Xa��|�U�!��ݝ�]䎻���<�yJ5��5���`迎#���$�ǯ�4�.�z���g������j婑���A�7/� iv�C���ߵ��0�DnDj�t����8��� G�t5���5�n���z�I����|G���h���~�x�xV���\������:�q���Pc�;5j6tQz�%���9/:3�4�vy�D��U�V�.Z�A]���iL�t.�Q�+2J3�c�
tp���Bs��q�%��q��w����ѻ�a�8���#��2MtzBzPŰ�zm�)����:2���|���}�GӤ�ƒ���M]P�\�͇f�G#�	��V�ٶ�	���%4��i�ZL�P廒��ԘR��E)g�ˠ����#R0�w�Ѓ#'��tKs]��9j.&��o��l�m{B��z�#t�q֕t�t�Ct���*S�]�Jўl&2�m����uރ��`�}���e�ExV�G#����0��Y����:D�yxR>�OH�����'2��sm��P�W��9S��4�/�l�j�C��.M�m��!�a��{64�z�/���5P���fKb��68=#l�%u�g��Uxi�yT����U�y���&���J�+|tl��j�u���^u��ô�2����#��FK�lv���XjqZM8��X#%��
v�1ލ�7.2:�˸T����֬Kܨ���VUJ�j���Yj��cMr�7)�R�"�Xb�
���P�4g��d|=9�C�����R���Y��y�u島�q���_�D�������:-�]A�:�.�`�.��b��k�W`��4e��qr��q�;F
�qӢ�� &��vNb�P�he���PZX�rˤ����Y�˥&�n�3�j��d0p�bo]e"t4�h�9��h�:^��8�ш]ֶ��]9��u��$�*V�/��n��k��K������%�K�I��~`'��&o��R:�%�#�C�O�H��s��!�3}��B�� غ��J�V�����^�[�::���?ss5��H	q��h�-���4�t�L�
��+'I�����x]gIvA��ѸָV�e.��x�7M�� <.c3Y���x�M^IaP�t'J$D�3.A���:u�R�QKjc"_�V:�*7����$^�wQ}�ɎM]�v�Z5Շ�)�'���1�In̙�"e�	w�p��9,"j�Z�/�WV�����.��PpsyU��=�^�����W����%\S�d	�n� �)��f�8��IP@��S�U��̒K�KWoQY:�#\O7ʁ�P�+�R|���*�z�t��SCy��d��O�n�;Ɍ�������ʹd����LdI��d¿v�� �jN<|�=)�庽=�<к7�ᶇ�b%pV/��ԅ���¨hL�niL�K�'^،5Ҿ��X�XJ��Vϓ���Q�LV�JQF�N߭�
sL�
Tp��I��6�d"2r�zl�i.��t9c/�ʸ��.���w�:��Tb��JX�9�M�y)�[*T�@pӕ�Ά�p� ��+V�]�2i� ��So�����I[��Uz��3���y�-�ۭ��1�9qq5&#V&����/�ϧ��噢]����)<�]��'`�s�fF7�=gƩ��)�]j���u=��:[������A�HwJח��5գ��*��a����<})-�"\0�S�ύ��q9�]0��I��F55�ĩ�[ܵ@��.�c�`����50��K]��b债��{G�#�8&y> э����2w�ٙ~�JU�n�K�.w�{d0bc�)9A�3�+���
�.ַCso�K��O@�������=���K�s������� �AMB�Fa3m������tS����Rl)@QN^�>�.�F˞�Z{FF�^�*���&�M�I����y�h��WA���[��zJR���p9R�5��T�qR�}u���"1��biB�Fv8��*_����r�ę.H��H#x�+�����'�f��2=�ɏS�{��j�b��3ն�i�e�C.a�xd��� V�Ӣ���:���Oc�#�(C������AB�PT\�� ������B?�!I�II�����ga��S���;2R<G��bG��̖�����ZA���u��m� Kl �oXI! �I! �$��ZY$��ZR@$��@�� C޵�A�́ �ЁI�%hʋUE^�QAt_\��X�TV(�,X� ���ɉ�O�D�!
���C�']�-�h�Rw%Ű��~�3��@��d"V�?�쿓�}����\���,�Rh6��,�M�J��gH�����š�4p��-a��T�0L)���Yߒ�� ���"�Y�	�������RO ��!'�'�Ԁ$$O�@d�a0�������
������0�ˌ�2��7�!�����>'��3��=C��#O�h BBOC�I����\�?�`�@��C��?���I!���hH{0%?G���I4�æ���O��?��������Y��0�?/�=O�ٜ)��G��=�;���XO��)	$�$O���g#lJ���:���!!:�B �=a��]({e�$�/�!�,��)�!p.������w��;����5�P$������x%@U��
�ac�~���>�����zy�Y��1�;B�_X� �?P�a�O�C\��d?�5$�s��?�A�?��M�~��P���x��8��n�� �0{���o#��~�oxǙ�`�A��A�������c���>Q�)�X~ؼ쟬���H�?x~����~��O�����������		9�D��	8~��������zp088��������[ ��H@�������?�?�0����d?bX���0��~�i#�6�?hu�ŝ`?H�pĀvN�~��N��S��D?�=�'uYMM����'�?hzI�l�"r�(��$?�@��Od���!�Υ�ă&$�Bny]� ���� !!"���w����?������� ����?����I"���B����~�����������c�f�����������f=����Ȕ�����������|��=����Ga�O���8�˧�=�`k~�����B������;<�g�d"��@?����!��`		,'����ه����?�@ޞ!���> zy7��W���o�䇝��C�2	����dp�������:��@�����C�z	�� >��}.��߁�xx�I����=�Ϡ Ą�~i����;���C�~��C������`��C��z��z�������`��ge?Y�?��{�#����a ���`�?��?an���	����3�M�����D 		?\��?�?��j��Ƿ���3���&�^��3G���,!���0@���?"I�~����]��B@�a 