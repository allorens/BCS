BZh91AY&SY�6��r߀`q���"� ����b)?}            7                                 � @B� ��>�MeCm�`  �`  �           �(               [<B��A����**����RR� J��*I("���! �
��%�APJ�-��"   �IUR!RJ�$�Th���'����{5{�R��� �9�ANt�� S�Ëѯ{:�I�t7��:�cOn�^��   q�IJ �*�����o}�
+�|x�*��P�(����Z�$hK��� �;� 7�҅^ �z}����9���y�<� �  A����)P �UT�*�U�
PM�ʔ���Js���aҞ���i� ��w�� ���S��v9>����{��a�` x�ª^ X���`>   ���) ������{� <{�|��| 6���p|v7��`�� 發�7^P*� �w����ǰ<�t��  @j��ꂠW:�)B�	��J�jU#�l@@g�n`�r uRMp ]a��è��ǣ҇�����< 2B�0   >R����!ް s���W ���<�{ y@;���@ݏ/@;�{��C��    7[ϔ���H�� �	UU)$� 	�A�&�݇@@�e(^ -a��z�����'�r�@�!Qpk�3�8   ��( ��� -�iAN 6Ǐa��Ԁ���� a��J�z`�`s�����X <P  q��J� V�Q�� �UAB_ f��}�}� ��g�Tw��J��@@�A֞�����%pkk��;��  �Ģ�EB�>� >�9 9cʊS ��`��`r �2 0�z�"�l<��z����=^�� >  �  @   �L�1JT�G�dmCFA�`&i�S�"RUP�   �  �Ѫ�1IJ4412hLC @6J��TF�4 � �#C	4��*R @    TԆ�*$�D�z���h�z@h��~?��}��_���t��DG.AA�]e���3y�e22�wn������B/�@9��������@D?P *+�'� 
���O�����~������#���UV��U^�Ѐ*+�0hJ�� ���?��~���?c*~�0��"�Ȯ0����"��.0���� q�^2 c
2 c 0"c
&2(�� c �0�c 2+�"��ȡ�����3� ʡ��� �0c������0�c
�ˌ�"�0�c0+�*�*0Ɍ<la�0Ɍ�Ɍ8Ì0�c$ˌ�c2�.0�0�33�Ì�Ɍ8�c2Ɍ8�1��8�c.2c.2c.0�!�8�3��Ì8ˌ��c.0�0��N2�2c.0�.0�.2��0����c8�0Ì8ˌ�ˌ8Ì��0�8�c�8ˌ8ˌ��a�2c.2c.2�0�8�d1�q�q�q�`�\d�a�d�Ld�e��2q�1�1�1�1�0a�a�\a�Cd�\dƘq�q�q�q�����\a�\`1�q��q��Sq�q�q�Ɍ<e�e�Ld1�q�ld�\d�e�e�\`�	��Ge�Cd0`q��GL`1���	�aq��Y�a�Cq��Ce1��e1��d�1��Le1��\d�a�Ce�q��q�d1�i��Ce�\g��!�`1��q��C�0�q��q���q��d�a�a�	�e�q���q�d1��Sd��q�L`1��1�`1��Ci��d1�`1��L`�2�q��Cq�	��\`1�q�����\d1�q��\`��q�q�a�a�n2cq�d�L`�	�q��d�\e�Lg���\d1�q�q�g.0ˌ0�Ì8��2�&0��8Ì��c.0�L8Ì�ˌ�Ì8Ì��32�!���c���c�0�ˌ�ˌ8ˌ����^0�.0�	��ˌ8���8�c�8ˌ�Ì��32�&0��0L0�.0�'�2�2c2c.0�2cc$Ì8Ɍ8Ɍ8Ɍ8Ɍ8���8Ɍ8�c&2�&2�.30��8ˌ�Ì��1��ˌ8ˌ0�2�&12�&0�.2�c.0�1��&0�c.2�.0�2q���8Ì�0�.2c.2�3�q�2����c2��&0�a��0�!�2��0�c.0�c!����c!��28�̆08�c#�&0���̦2��c)�̸�c!��0�c���0��c	���!����q��)�&2��!�2��c)�2��aq�8Ɍ8��ˌɌL�2c&2�
e��0�c�0���L+����
�!����ʯ8�!�*�"2�������*�
�0�c &0�c �®0��0 c*2��*�
��.0 c"�1�`G�������� ʮ0��!2�� ʎ2�� �.2��*�(���0#���
c *8�.2#�"�*8ʎ0#���(��.2��� ���8Ȯ0��*� �0c
�2+�
���.0�� ��Z*������asu5R.�D�4�T#�����6
�Z����\�:%ދV�i$�&]sy�ͬZe.�][�'�~Ꞝ<�js��+t������#��\�o��C����a�ge�`1�^�'�z2��^+!���!�֎�k�f��ަ�%�Vq؇q|�q$���nR��"y\�8o��Z����Yǥi��6s\��e�g:I��@GwG"QM�	�x@��u� e�%h��	&W�[9�N{�� t�nh,���&=�EZ.��;
�;�3S�.m�3�f;���1�vbUL�4�ͣ��7p]�h	��b��	扳��; 9t�p2h8LG.��u漍5��LaG���c"�*�ų�UzU^��0��H�Ĉ��Sҁ�;��(�s��T�B!>͒�wt�[���J`J���m��W6����k<�g53`yN��hi
�~���i�cy�E{�iG�TŶ�v�u՜��N]/E� �V���ۻK�d�8v�t�U.����N�-˽��ԖwX3���#����sV��a��wŵ��t�%p�ňg<��}ݯp��n�Fv�Gm��"1��/�ǵ��Q�秾
:��f�G0��k+ax�m�qe�	9�˼�bBj[�n�$�[\��q'O
�w����⭢8kSMV����آ܂Y#6S�|Ni�`�L{�֞��㺝,Ѻ�M��eod3��+!Ik�.G�d75���=š�*Ғ�OjT�;��$Lh�4��V���rSga�ܪn���1�$(%��
1|�_J=���#�G��m�xzwr%���(b�����[X��C/bG]�8$�f3Ӹ����o��p�ǫ���4z�o0�[����C���t�R�=48���cGA
���[�����F���F�0�n2��|��vWE�m.u��Qڔ2E�܄U:��Oo�N�[�3�P�)�����f�ζA�e�����.�d��n�"Ƀm��|47�ܬ�Ri���^r	�\�6�t��.M��[&ӞD�u'J��k)�@��Wt}w-}uNA�c��"p���;\�i�FAx+1��qOjX�dǬå��'N��7{&x7f��i��Q����OM5�����Gl�8t8�w�#��h�T� u��	p��i�ݼ)fr�yv7I'w͸H6:��㗵��Pv�ng��L{��C�$wI'r����ҳ�ۺC�B��wkx�[\�5�ٺB�G�d�T3u����mGV��
:[i�E�Q�/!ܻ�Dp���صn�	d�A<���k��ڬn�NU3�+X�0w@�5�����{(@W��WK�5�Z�n��T����
hNd	3f��d�ryL}��0�I��:�;rY��.1#[�!�����ۡ��9�#�
n�M�dWz͉K[Stg>܈����.�u Ղhν��o("��>��3�$�
/}�-Tn��T0mɫx�,�����l�%����4���*b�X�Ț�NT�"�E�#�e��.��l���v�
׫��ݓ]���Ui�
ɓ�x�^r���9�u��*Fm��@��C8vŅ�e������R�Df�@�C|U�����Y������	K��-�v�ܣg��!�9۳M���l����۞�Ǳ�"b����1%u�K;Poy;�����8<�����՗.sr|�� ����	y�9FΌ脝�ν�|Ό��@��0�Gk��廌hyp��X�2J'�`!��v�����1خ$�&��7��Vᖑ��MX'i^םp�Xa�I���ܪ�䘪K���]2#ݍ6�l���hWcM�NB�8k8�=�{���I��ó�nm͸$Я=��e�y�pw����ɡ��h�t����ւF����!n<�aE��mL%��Y�n^W��;����y���3�c2F#6�=�Kћa�q=�k�znoL�Vc�݀��O ��;�g�gj�
��m1��a���Y����Ni��N�:�%>����F�n�	���2vT7>H�;�k�#[�>\��s��{���Ӏ��`�>n��s�ܺѹ�<�؏�,�9��,�t��P8�7,���`p��ۦT�:$�z��\p��*�n�XX�>-p��'�ɚt�n�YwI�ǨCF�9�0ޙâ��b 1n��62�-.���v��G˥��6oL= (���N����V�:^.z�ø�Ү"� *ۭM�K�(�p�c�uf��x���02���S@̈́PWhX�VI�$�U�/k.[�(ږ���񣇳�s�R\�M�*� 1�mD���h���#oiKV�!i�u�E��M�9�.�Q�YVY�C��h ��[NcŤ��ag
��`���p�Wm�1��]�l�G���>�c��*Yg{+����j��� �=��lM�1��t�e��wT�cn�61n��gf���D�[��s��/�n���r[�}�-�1yv��
|z�/l׸���4v�d�ր�nC�8��NԦڙ� ��U�E(
��y�sS�WQ���=��OmVw�it�ضTx�;��wW4�;ݧ�a=�ҷ/ʷO9U����}�W���(���Z��P�e+7CXWώɸ0F&�jֵ���
㖁��P�:�͗���C����Ϟ]���;L�1-�t�Y�f��u9E1iG��Ξ�<��P��"i�s��a{4r�G�d���݌J��/,ZoF&ֆ�f��nw��fV��i�jҎS݃��{���G>d��:3���Q#*\Hg{��	Slu΂N�*��ǻ�n��[��N�7EwGpUhG��b�j��oA�v�Eq�J��-mM��Dg�uՅE�3�4�"�5�b{�$���ێ�������k;��g���<��8�Źf���ں{ 8y�J�s��!�v芪w��+;{5=�fMY5ua���Hp�Gt����b��kn�xk�@vn2��.�Lu�l�ji�������h����N-=�H��z�c�#�e�w%�A�w)2�7'>�ڲ�Pt�`�ك�I{Xi���';5uF=/+�h�~ݤ��u�Sw�
}�٤�數f	RY3G�����r��B�"�[E��ӣ7��5��Sܦ�[�Mq���-�#����wb��95��[��8N;�3��E�X{:���o�薝^*y6�,YZs�ʒ:�s5vT&�ws�8�8�-2t�>9$�v�;�+���ӻ����3��Ĝ��7�ηM�i�|�,�i#�8�D5�w6�d�k`���`���
������ ����k=��8�\�rQ��D��+��}^F���M�;w�x'.VA��t�����v��Y�k�O�$�a��/7�G*��{V����n�L㵉��!OJ�rU;D��j.�#Eͯ�p=[�qi�n�Wot��Y�zb훳H���;w�=@(�1�5���6�ӱ,���j�9a�ל�\�}6-/Qۍ�c[򛱢e`Lع!8^����u�F=γ�yT�u�/
��+��%fgeG9^�����T�vJw@2�NӔ����{4�0��8�FJ)�un�oym�ՠ(��3+M����ϲ��9���<D�Gt<���;�"<��y_Tjpgv��ئ��2ܻ����x��l4z��4�D��_���i�ym��Z��� b˝�i�拽�H|�-�Ƃ1혵�s\�7�H����p4r���þi�*m"�	�^-��^���_:�<h��k.E��WN��͛���`�!vq�-�|�7����ڽyJ�ƈis;0�˼H[�m�0u[�6��!��T�Ι�}{Z75ʤ/���c���[��^� �h�Ҩ��lH��EW��s|��.���`�2n��U2�G�������t�F��ή�ǹ��x��J�Q�uv�vV����b��'�W����͹ٻ�Ʃ���*w�4�R�^����3H���L��v��K���ۗ�nB�t5(C��>x���!��U�>}�hx��7r���$���&���Pq�,cs��]x�.<���|>'�&"Q+�UI�s"b����2�@�{��8;�v��Ƴ[���`����Eޮ�wklQ�M��`��M��oU�C�Z9��^�n��w7�Rr�%��z��*玙��ԍ�_�؛�[��x�H��sp�tj������:K2�3G���务�׍G.��#�g�k{�ē.[�	�R��M1���p�`1�c,��~�VK��,���������:7���jǮi�N�rk����s!�;��b��a�5a��P�%[�%ِf�˩bEJI�F���9��v���GӖ��i��X���}�n=�N,�yQ��}Z���eÝ�F�=��.�1�{q�����b�*Bv�:r�����z��ǯpঙ�;��!�!���L��-}2&[���wEGvIvQ_6���VQ���߮��ġՋ�HЅ�ɬgUB��(��\2tZ'�t�Z�MW�gK.�����[�ี���'^׻k85�u��b��#�+cN�����=�VGMO.Ά���h:���Tk���l�z�y��q%-�p�в��W4ع\b�h@7��`��ż����S�Ǜ�oQܶ���t�^��Ԛ^�I�̙r��r3��_��	�����ɭ��8k�t�� ���F�Dj2A�kn���i���	o\�79�s��۳�AªN"^��o �v3���.�����Z(��4|x�ܯ>iی(��Ц�r�����Y\W�3tJm��s� d�7f��%���GH�x�sY�{5�K��;�B9X��SZ���R�A�3�z�qb�k9�s.����Ĕv�db�Z,�r�;z�ރ��r,��ǈ[b���8iyJk���y���]T�SW�{��^�๮�6����EC�WQ��C���nw���(����񸯽�f�i�u:G������Z�b�"�%���9���������Ô��C�hx2��sF)��zmG���qڒ�&ΎA�y7���^��l�z���Zn�*n�(O��!=��h�5!^l�6V9ۼ�el�&�,-�aegG)�v���� �;^��]�1�h:��no��u���i��L��"f�_�ub����o�L$��a�nV�8>䉸m��q�_N��/K�ʬ'�4��4���2�f�fo�H���ƽ��l�;w4�����ϻ]���k�Q�v�p���8���
�7dY��ib-7;۱s$���G�j�$�${�.0��nЉ�*����\��qbs���H}���5�ĉ��`g���d�)��"/cʣ��"n�s���;{�bk=Anm���3D���诘�n���w�XñM��}"jR�49�;���&ȅ���*��3f�G��ׄ�pK����8݀b��^״���鋡ĸ�Ŭ�]/�_do6s<��FWUZP b(�E���D�ڀ<z	��8��4�{zCu��D��;#��� 1�F�+F�����܊!/�f��b�z�B����
�!� ���(���R]l�t��Ը����m���D�7{��[4?{O����h�l�7%��Evݰ?�����㿉��b4&��$r�����P��b��p��2�턳X����z9����Dpu�,�e,Ø�A4��R|�o��!�������@I�=����	���`*�'v�{��.���&t< ���t~�_����� -�	�YG�y�&�����D�$��Ս��
��R����WN+�y' ǃ���ӯ���ü��to&tdG����qoyh�l���%_���NjYV��د/g��s�6�g���F*�_uVz��P��%Ð��}:�g��#�}J�VG��:r�7��N{�f�	���>lQ1c�Iy�#J����~�Ň�0���}�K}��0*�CڬH�lٳ5_����_3٠�ŢM3��r�F�X������~�X_��<T/�T�N���"k�ؠ��zV�����g]h������qAa�z^��ܟG�ļ
"�z���u80�=�	|e�f�NI��yw{g�+�!�{�#�<-�Ҕ����{����=�;���3���nox����s�w<iז~�]�
���pw���;���]��o��c:��_����p z�'_H�M���q|qETL�B#��Q}<�:- neD��=��Jų�~�NmyQ�s��IwL�!b��H�B��dD�P��(Pd�V�?z������[[�o3�J#��3�ݿj�F�:0]�Ν�b�GX����+m��sb�F�N9%,_,#ݲ�������iykٝ��j��
%c�~�w9`�?�ߥ9�xx�e�}�i��w��L�[�������y�t_���}��ڷ���w�fí��C�@W�#"��)���rM'i�H[?���:t�L���{a$U!j��?7��[�����'p�q��n4L�
���.��0����J�$��������绮��̹x��zɁe��Л��0�O����v��L�|���Y��W�����Y�c��)� Lr,�۰z^)e��)�0µ�]��w{c9̝(�wU����1��q�"?�.�m#F����o[����V�%~Iz��[����n�Wg��%�������C��4j�}��V�� ׸4�,x��q���zu����+�nw��3���7�=׿������G��L.H�Ӕ�`�C0~�@9 �4Њr�P�*(� C��^H���"R 4
�
�$9*�R�4����E�9�O y"�K@�P�"�ҋ@����"4�J+H Ҩ%	H�"� � �( rG�����B�B�B���!�
�%	HR�J�+�y �B��Ҩ- /%AH�P�- ��y ��*��R�R��% !@	@��/-�V �B�
�I*B�ZF����C��Q��Ic��3,H��0p"�qD���ApT����7l�	�t���E��/��[<:����|�3�Q��|�y�=yy��v��v�.�BW�rl_��Մ,���}}��D@��?���`�c(
YI��BpU ��U
~h ��0�HE��]�1��ɡfM�Fi�pLݒY�K���F���y�V�3@1���g��_^:a34ъ����4}6�3���,"
V����X�>D�^�F��'������а[�a ��(��b8w��yw1�%�e�����g���%�1j���H���z�j�7��m�J�:>5�P1�n)����~����~'�HgĜ_��2��N��!������$��ֹ54�#��,�I��"�@�M�H�m�~7��RѣM����ma/kPU���9��&��7�<DQ��Oj��D�U��9�㊸j�<}k�ϗ����#1�aV�i�$���� Ȭ�H�,FG�&�����b�km���k4�P�|��b_p6$�!���8�� ?1�c
�TxuĆ�a�ο���Zy��h:~قg�Q�l������dA�È�gO��f<�C�8٦�V]-���,�G��{�z���w\Ы5,�4_wϫ	��E��D G��O��:@�����}=�?�� ��?�A�O����y�}>����������|oϛ#g���0�hB�9g'N3���ǟO]�.8�Ḁ$p�*N�o�Ь�==���0���������>��Y�1��Ud";i����÷<&�9�p��Te��=о>F9f4���\�����{�x�d^R!ۢ@��>�s^�7٣4��X]� "gY�3�StM�n��x�nv�r�����	���vx������x���g��k��6��A��.J�.��y��Ś�{���{ɔ[�ު�i��t��ڴCC}�q����w��Z��y��,�������F�������j�lP���jw���$�����g�Ow����L�}����`�j[t}��#ʌ*@�g��U����`t�N	����P����;��X�j;
z6���륭<���{��f�ҀJm�� �H�VS������W_s24��;��O�t?��vp"�٫�=#�̕�{����Y�=�����z�g��ג��6>|�uɣr���BG���H�����=�%X��ۏx�d3��� �w.Ղ�G�{ZѺ�&���Cd����F�邎�d�\��Z�.��D�7Sg�%�̳g]��LC��X�e�1tey�������������c��뮺�u׎�뮺뮽�κ뮺뮺�뮺뮺�۬뮺뮺�۬뮺믧]uק]u㮺뮺��:뮸뮺믷G]u�]u�^�g]u�u�]u��뮳����]x�뮺���]u��]uק]u�_N�κ뮺�n�κ뮺뮺κ뮺��]x뮺�Ӯ�믧G]u�u�]u�㣯�]u�^�u�]}:�u�]q��������ޏ4N%�Q>����Ҽ� n�:6Ǭ�Ng��/e�kb�� 7i��[҅�������jX�5�_r����ǽ���#��A;"c�yj�7�<p�t��-��߻��׺{x�9�lDf�+|���h��{8�"���y.��̼��3�N�{h�^���H�:�o�iG�C{ȽՂ���Q�%�Jc�H����;A��s�\���ӳ{oM]%���K2|�U����@�^G�+��1�T�:�������ë��x��!�!z_������33�L&j�V�^#�͛�N%ط]�:(5i�{�φ˹�2���E��̵�h%</%d.y�������>M�>������^��8���~-��qv����w�uE\3X�e$�AC�-��Gf��2n�6nM�jd�.ܓ��m�ASTS]�ˀ3~�3r��~��������'�ѧ�M$ٜ�+��뙙��_z=������{Ьu���l�9Py���Q�Y�皑�[m^�{�]�=�R��y��2�e�d%�>�cו���oe���Mi�|P_t����½��F���������C��������I�Y\�޵��˝6��X�����Z�k 5�<�e!��j���X�gQ�B�@�{�X���v�ƶ�M�������n�뮺�ۮ���뮺�ۮ���뮺�ۮ���]u�]~:�:뮺뮽�:뮺뮺��:뮺�뮺����]u�]}��:뮸뮺믷G]u�]u�뮸뮼u�]u�_���뮺뮽�κ뮺���]q�]zu�Ӯ��u�뮺�Ӯ�믧]g]u�]u׷G]u�]u�뮸�뮺믧]uקG]u�]u�_����]u�]}��:뮺���.z�7���w���7�ʻ^�\:cӪ��P���o�ˁz�1>���Ҩɯ�������3��{�}�y "�V����[右1��mm6�=���)����"��-��t4Ǵu �	x�3W����_o�,򧗇�����Ќ��t�Fz�{�3=}�\/�V���8vn}��ۢ���#��77�tܓϞǻ�d!]j򯠾��	�#{���������x%�vO?c�$r��b���Z�������a�!��8�o�����^��������KǟN�77��{�oK�}=ggz)��$r����͛�O��7C����<��2����h��R�0v�ho{�f�<�|G����q�˜��L�q��#`������y%��n�ټ<�ޔ
�Q�o_^�W��`���[V���ǻ���<�ߩ�1���N-�H�}�r'�ϲ��O��z9�����{7�a2}���}�>/{���ᇠ++��v-����;��=���з��U�3��>t3=�;~�Ec�x˨��h�L�����<1
=�[����b�{����c��i�f{������}�coFOtۧԏVY���5�n���c������t�G�|]q����������뮽:뮺�u�]u��]u�Ӯ�뮺�u�\u�]u�Ӯ��Ӯ��N�뮾�u�\u�]u�ۣ��뮺�u�\u�u�]u�^�u㮺뮺�u�\u�^:뮺뮽���뮾�u�^�u�\u�]u�ۮ���뮺�ۣ��뮺���^:뮺믷]u�]u�^�u�^:�u�^:���]{u�㮺��]u�㮽��뮺��]u�]~::뮺뮺뮳����=��)�������xq3Ӟ%�������ޔ-Շ�}�t�_-��,+������,~]�y���_n�_<��mA{��v؍�s��0{�[�I[}���-�����oc��i(j�ݺ�<��j���i���~9���p��'��;�7���޳���g�ĸ�͢�u+=�\���y�"�/�CD�5b)Y{��Q�s��<�S>>x���\7:��C@��J�C@�^���?}��9��.v����j���L���^4�7����W�x�u��{�ԩ���Ɯ�O6[>�چ-���w�+���ؼ��������_Sx��,��x�����}���ڦ�^��Wv��Z����낿{h�^W�S�^��e��%��Ɠ���{�a���^���x�>]���8��^::����W����Ow��X�y�K�Uţ\i�f�赍�uuŅ�ޣ�g�HBo����,��x����=���c ��F�/��g���c9^g۞�ݞ��-}�R�'�5N߾�����㇄w�՞��^�l�����D�M��� �͗�N�y2̵�����ѽ�<6v�����)���z1�����,�D���� %b�>�<׾�n����o`��4r�p췥�M�ք3W�������Mվ�<��>�;�)s��u�����mt{�$�Ϸ4��9g��W͠�׏AѪ 03�W_l��@�5�x�~O�v=��Fzݯ�E��t-X�Vh���n�a�ի����i������W�=�S�y��{�x����c3�� ���׶u�ކ-���Q�x8���r���f��nf�:�x�,ّb؛�B�W�x�;��,�;e,��gc��W%�v�7��JC�zy=�wk+�5i�S�aqNl��h��i߅�dr�	���d��Cpo�Z�Ǎ���-~�-�5ܲf�r�}ƨ���d�+�{�g�Z6w�m`�_��{�!p�-�;�P'|��+�̳n�=ݜ�����~�	N�b��y���!�3@~7�L�S���Q���6;QKǞ�\l���m������K���gY�K�	�;���7ۅA��z�~�,9��z����	��%C�71ti��oa�eK75<�|��|���Eǅ2�GY6y���i;�\ܪ�w�8_J����s�,;��z4	��5�'�܍��r�|3>VFN�+i|b�;���׏X��ͳ���������xĻ4*�Y��.�����\�,ϲ��*��LϳwW��4�xy�>�GU�� ��^�R~\����8�S���دxL�������<O���u��
l�8����փfK�{�8�Ip�о�ʓ=��V-��7��M����f<��`^����t���������x{ۚ��w����o�|�w�  =A�X����br1�	�c&�3"�_��{�p��:mYBL���Q�-�ｈ��q�7�ֲ���f�{�s��x�_��{�I���-�9M�淅��v�K�s�z��g�į����f&�'�R+���r.;�g83>��T��{��(s՟>���3ü�ֻN���;�+�'�d�9����^��xb��ZD��H5��<�GiA]?fe�����'v{R���I�۾a��4�/<���wu�\�^:",�A���{u��:��{~����`�t'>����S�����Ϫut�5�9��xb؅�_����̵�8j:����o�D��9��-.��X�>ېoH	l�����}��j����XlӵA�h�}��� 7�j���t�ϳv�jλ�����v����u�9��E�p���iY�}�&����_�+��J��>raoN� r���&�B<O�%�sVff��à�'��+��No�Μ�����,����5��}ž��kb��� OQ:b�;-�Tϳ�?O8c��/��l �հ�3���XȻC��c�f�]_}�����ߕ�
���*.è�
�6%�=�;�{*ϳ�qRu���р!�{qxOe����òз��M�U�{���y'�6�u�2�RS�;�w9��ՙ�x��2��X��Ĝ��͝��m\5ӷ�>^�{�+���u��d�7�\�y��q�^��Uz��ϲ�w}�b�~̉i8�ew�N��t�ý������r��gٛ<��{_`�"��Hx��9�����Xn!�}�,줌,�p"u�S����6$3�Wz�=����K�t������|����W���s��ݛ�5����[�C��>ɓ=����-v6&S�x�4l`{�"W!�8C����ʭضg<��;7��97��}�M#}�n��7�0�����y*nnϦ/g�n�:��������?d��4���3��*���da����2|w�}����ϽϽ�c�[��b�#�=���� �}O�+Z�f7�ＳQ�`)=���zy�x`�'������K��K�O+��f]>��y_"�y����X�9L��o���]�^f�5����[��޲���3�g��	��:6��	��9�wTy�>@4�wx���%I�ؽd�}�g�۪�[�{OU�_����<�q`�	�d��)q��3Ս�O~ڹE�r��s���xlż��Yh�J�9ϲ������jQ���{��W$��VL����w��&���|�4;��s2tS��Yӹ������n�m�9S��ܞ���{S�r&Jڻ;7fG��������A|(�F�W�q�~9�С���2��rњ2V�1���V�qo���}˦��G�a�(x:��}���}G]�'|��$��a�7o�.���WK����l7���帵��%�ϩ]�s����ۗǰ��鼗���h�^��ݾXy{��{e�K侏�fϾ�R�i��	w������9��C}��
�/^r������c����ż�_}�ކ6�&/��������||�|���P�����������7���A|����B4��;^k�k�c3��>ۇ�p�P0�?G��6����}7�8u��w�c=ཥ���y�|w��x+��6S�u~�#tW�}�p���o������dY�m�z;��vG�M6�H����S���W��;C�����s�0��,�|�+����`�/�L�~�����Q�<���Ou���O˟������Ε>�>S�1���|���pu/9�y+�O	�L7�{������v�]9��p
"Κ�6����x2L1�v�w�������7����9�lo��(�ɮ-��1��p�(}�p#bg�՛�q[�^��J����. G��6s��'�y��zＯ��b�oC�I��e2xؚ��>�,���=�5��|���'��c}�0�{�s�MV����"��>�l�n�[�}�;~�^8��M���AW���:,D�{,.~�rV��n��:7���s]�hrH�_o���z���t�6�ۜ��G�k�U��G�~���}&�ws��x!��W� p�����M�s��|q�r���x����X흷��3W,�w{�؇��Y���A���]��=֭��ŬX�c̑`����M/U���|_!ts��au���'��Ͼ�Y�Ϩ~>
��('���[v���������6{k~������|i��&��k]���������Ͳ
��D:���蹖�랽���Lp�냱����b�b��}읞�~������p�O����� ����w���ju?yn?_Q������_T;݇��&���4��ۏ���Dvه�( Ѩ�<ƚ&	B�gU��F�،��x˥?��釕�dtf�������vqo�o� |��g����͝����(�?�ղ�Q��0�Gu�N���j?떯<�N�cg:���s���6b�X<�7a�_n'�W��3��ݧ�Wɼ���j��{N/9uUsf,���g���q)���'����NQx�����7�O�6s���g�:Fv�x)���[R��R~�͖�ø:iP�U�ֵ{�'�b����}'���r�/w�F�<�\ԍM��n��I����ۯ�������,9��O{$>���l>��Fq���v�p �w���'��Vy��=�����G�Y���+Y�x%�w��}�k^˗��]�f`�w�s����yN��k;�;Y�R�Ã̏x����Ok�y��uo������9IZ�̇�#��^0bA���9`__?�����4�l���\ל���;��YZܾ����;�?E`��S�ݥY,���wo�dk��$g��0�C�ʲ��@���uU�s1���m����;��s�O�]Ï|k�ٜs�;�f�}�pկ�}�<v���j��(m�tU����a3�:=��G��H�n��r�釛���w����������I�O徜��~O(��e$���Tb��ݕ@�������*�+��O���o����P ���T�~_^�_���1s�.ˠ�D"�����a2��T�Y�Ā~M,�(h�hc&����<�b(��m�y�k�_J?��l_=*����¬.Q�ncZ�W7d[C 4�$i�Vҙ"�֌��5 �z��٭�lk)EI��Aظ�"˓&�/6,vt�D	a����l��ق1Z���F��ka�F�k8̥��V��0�9f�ͦ����ɬIB3n9a
޵{a3jĖ̷u��pr��u�\���:݋��ѠAѮ��jK��m�1�����
`�3,*as�`�i����R�
�-�iRM+���XC)"�-c�6W$���7դ�5�. M1�/6�����&!��l+���˱�����K�2�޻v&�1�db���,t�R�ܦ���0m�˱v��CB���� 3-���)��J��k�f+�itK��`�%�̵��İ��M]�[`��\A�Hm�Ba����XIr�Kq[,��� E
]��*��.v0[����f��i�AƳZ�(����lf�<��0Һ.Ѧ�F0tc��l`�16c�.�tP2h�I��T��]e��c+��J�ZC[P��H�q5�ZA*�K�a3���L�Z\�AT�J1�j�vy�1^b�1՚XL���-X�`�RQ)M���2�P׷]�v@��\ݫ0՚1�[�H	�l�tih�sWr3G$�Ü۱b���f�ͤờ����"\ǔ�m�͍wX(E7\S9\�	�M�5�l)˥��.��t6�e�-Z �Zd��X��<s(,��f���RYBTԅX�V��jv(�.r�4��E�����Ĭ�51Y.Ό /H�Yu٘�EP�t��4Y�����G%ں%�[-f6ᔭ�����:��'Xi�in�X�f���L\58�p �͋#m[�i�����A�̴ҹ�-�:��j��@���9�vI�β�[��l1��r�kp�Kŭ՚����4�vXR�\��p�ħ$� R�7�kt�@����h�ث\;RR�)3)�X�Keƅe�FT�]�+(�P��#A�-n�3Y@����ƍ�������1l���X;k��Km�a`3dã؄����3�F�o��7m��n[��A�u�4�m��!X�d5��E��0� �!-����K�C:62�[�F����%6Ț�<i��a�uxL����0��	5���U� <kL!��Ͷ[5�y��N�K�Į�"1Εd;Z��]����!ͬ��Z����ƙ��v�("�M6��c:aF� �@��@��Kz�(l��9v&���chjK�T���- 6��DD-�V�G��P�1t����[,��GJ��m��
B��ƴ�fz�f۬ZC�)Jkt,��6����15�0�M)L
��VL�ҧ7.p��l1�nE�!d���jqi�^��ۛGi�#-/�e��)a���9)\jR�ᗩ���^��ģ��E�Z�;���"�2M�u�]�v�4!R�YWg�5�X�%�@��8�0e�V�G[�#M0ڰU��Yp�tÓB�"Mu(a,�+
괲��YkQ��E�e��]�h-�̷, ]�	t�]r�$`�2M��������A��+(FJւ�2ZFʹhڑ*�6,$��V�r�LUX�J�%p<r�qÕ���n `P�
�c4�lC���K��Q8��R]eK\��lXv���c�SR81�͠[�K��:��c��<ǷYx�+cZlZԍ�Q�ҭ��
�1�h-�v�Z�JiCkp4rD��z�Հ��
��^��f��-���������"�B[+�0�W&&uA�K3^�h�q����qF��XWsvdm� ��IMf�ɳe#��#.���+,�Q��G\��f5n55��Ά�Ѻ�I�L޷V�٤U�7��N�ѕt8���k*�gAX����ת]�1m[.-�-�ZV#�rE�pqF�a�)�3;<1�\��D�5���֨LY�/7��b�362؂]k�ɊM���aZ[e�)X
��uSS&m�-P�e��6����B��K)��0n�[+�l�$��3:�Jh�W�Χ�-̩Zұ�m5ѳ2��	�H��]�K1n�f-;Wl+y�f26�U�P��a����m�٥ ��fEu3�,���3f��b�,!�Jgg*ل{��Ywi�id:����mz���aε�ٵ�9�[%]�ioZ�*T��Ыյ5�ҴѴ��B«Į�q�-6�e���u��ʲ�e�BS4�ܻ-�]c٦t]ufeλ\J��R[E-�K��X�o^46).0m	(��4��M6�f�e�l��4�����l�	��i�@v4A�,�(K��^խ�،X�r����ˮA�j���JU��Y������kZb��΃�BX`ʙ���@+R	*8�̝��Rh 6�D(u	�5XX�q��f�0�iQ���4H�Ė�]`��7K�
�YB�stGe�����]��e6��0��� 3MX�c�9�8�Ԏ��m�7U\J]�Êl�Φ(:m�;+�AK�[)QҒ������$FS���C$��,��^���V`�v,e&���Q����F�D��
B-���iH�;f�"�J�R�v6CM�YD��ƀ6Z�������sk5�ړ]e&���6�9�ʢ�mV�[��PKL��i�L\�ƽf�K+�����*�ٹa�y#Z�p�Bf�*pA�IlHUnD/-�����!�� �\�6��53�Щp�$���p�vq[F�B�٭�J��(ĸ2�.%�2%��Tс���%C��i��!���Y\L\$z�� n%�օ��s���#�[M�F�h�LZ��0�YB�.- [�-�E�֓�l��nmګVZ.�;vu��2�ZW��pm`���Q��6-̥�pT�C;Ȳ��r��@��T���ֱ,צh�b�a�f0�9u-�ո��ґu�L@)�k�b6:�]e��܍��Έ��:e���e���L�ѕ�����KpWq2�,,��Sm�8X�+q��3�u5��i#1��M���\�B��Y��0&�h��8s��!�bAɉ����ѦfԪҹ5��,),[��X�ݴc�7;e�ivp�%�dͮN	����eI�3H�(�n��`$�҄�cnЖi���t�4�յ�e�\
ɜ��up�j�XBSj�p�e�m���Bik&b���,fG6�Bfթ����e.�ڹ0���YaV�������70�יa�.U\�M���ұtpM[�V���R2i���P�ʊf�v)k�cn�2��l��h3�1]Dڍ�
��(�n�T!��b�@!)��8�\�@z�
���æ#r��;m�)j���.Wh$�u�.�j�oV�0-�#6Ή�������.1B�3�M�q4��[ 1��6�$RVl�R�,��(��j���˭ؼ�1\�y@�Z��Ѕ��Y�[`0����ɣ�ݖ�Ҵ.�S ]�@��43��N�B�7��(�-tڰ�Vڗ�y��@�PЁc�f6.�щ�l�6.����iuZ$�T�Z)R�M,L��/-�H&n*uktQ�[M[�v`�8-�̭�K�bU(����dwh��n�pu�Y��m���08��HZ�	m4ҨU�7v��Վ,ؚVUfҼ�q��RT���l�l`���"�T�cS]�jK�Q]���m�i0�ٶ�UB�
�lY�5ɐ4H4�[��΍Z�),qaX�M�\$��h$Q��tmn&Y1�4ն�m��1�v3At�1��!���V).�����ʹ�JR�XX��������[���Jʸ���
�2�+4���8ͺP���ѥ*ǋ�
�8 ̶j��KBa�nZ2�A&�I��X�D��1c�27f��gF#WM[Z��&�A���w[Z��D�6:l���AG`&oB�K�s��4�TQ[�J�havj1ͫ�W]�.�B�40�jњ�V�"��t�àp�g�GkE5�)(s�N$u�e���6e�
-�u�˫�-�.X]-L�� ��
6a�5L�V�[�r�&	�i��2ͥ�͢��5��Gm��i�X��%���*66��e���3��\5ڷGfق��]�w/Z�u��ytn@�:j�	�ZT4rmq���ѫn�b���:�+��HUm� �΋��-E3��\�-�n�m*�����ʻ*���l��4�b�v��3:#��v��Ҹ"�������U*�t�g���Fe�]������iUUv��3*������l�p@���[P��n̲�l�;dZ�Մ=Zx�ष�6�4�B�T�� �Q�FFp�k
Y�c("q�H}37�ǐYV�j��Q�C̳�#��Me5�WF�P�� ����,����5 AaA���,:e��TV*EkTQDH����h�1e5�r�D�T�44�A{}��ӎ��u�_n��뮺��^��ꥅdX��TH��e��S��֪�&R�yaR,QUD`�X��*'yq<��d��jnrkۯ�]g]u�]u�^���es�*
B�(���Ċ(����J
�j�h�h�q�	M�8�����u�믧]g]u�]u�^��m4�Yù2���h,R,�]R�ݳ�*(ԭ��v��E"2):B������告�v�X:�0]�LVQ#�F�hE�PQ�5�b���,(��%�+�&�*�DR(Ŋ�U��P��PX��m�HZ���F�)U� �,� �lVAh-�$-�Y�&4+ Z�-eZ���i�[�2 ���l�\�'���5Qmk'3z�-��n6�Lp�
�V�U-�E�6�LL�Ґ�KBT
�A(�̸�(-�eE� �ZB��[K#U��Idk9�)\�bPjD�(��%1��Hd���03!ul\�5-�L����0��Q*m2L��D�X��VW�U*V����%T�ciF0��ʚk\��)���ms,�/xTq�]�8��������b*T+T�`\�.E���[iPbQ�mm�O\ʲ-��¦(�Qm)��ui�������Q��hڢ#�(����R�-�f�CK��Z N[�O�pi�a1�P�vӀt���iH�[*�]��V3#s8Օ�f�!1��������Z�4���UY]��8���]ݙ4`�f%��j��A��[1f�f��Ļ%c`��#u܃�T�{��ʁY�4%���,1�1���Q�f�5Vi���]v�W�f�@"]\���B݆-�nu\��5���He-4yn�(k�[N���b�Ѓ�JY�ŋ\\G���R�֨UՔ�u1���vA���]��:驍Hd�+�[z�aZ�3.&aX�x-�U�&���e-�ґ9b�IJ�ST�kg�*t1�
.-&#f&���ba3�fb$�9���ZEc�t J Yv�%n�a"����;T`���Ku6���CB� �KY\G2�b��S[�vb��֚��`��q\Q���m�;ZKz�;UK�Z�8n���{-�c$��tf/i��-Ɣ��#u�m���p�,f�F�A%��Q��G��b�$ )Uhmz��f��r���+s2�yZJ�WLG3d&���R��B-�1v�9�h��d��R*�Q�;m"@��e�,nՅ�cW�4D�İv��ⵗ��鱶�@����.�9�0KZ r��6��d�4-�\�Wie�e����c)hP-X>W���c�p�c4�K"at�,P5(E�]M��s����ō��-��.m�FYF]�-�i��fRU�&B[n�B�5��1(i`�fv�tF4iTb�h�1��.�yKM������b�������-m`��[��8ب��B,X�L[`����k7ah�Y�M(��#ra�4c,Cd�HPe���Ã@:��`��4 c8��NY���քnE�nvr�g*����Q�5��l� �ѻ-��n1�c$� :޹̵�q�P��)R�@B��61!lx�jE
�@lj�Z��R�h6F[c*/ �*�+bӄa�m�լe�����5i��U��iXU��
T:�R���*��u�Q�R�[l���`���B�a(Z�jţj0T٨g9�b��B�lB$H�j��`Հ%��!X�*�R���t����o<x��}��0ėb��ZA�bs2��������%��l�}=�[��oOrϾC�
N\ŝ��Rl$W�d
jD,����TN�Ɵ,��m��@E��N�(B���KHL��lQ�A��ěbN1�����Y��;���C��y};�#7&pz	;��K��;;�NR��U�)S�c&��ٰE%0�]�C�=�H=���E���?�y��f�Iڴ�'-����zǷK���a��v�7V܅TJX�d�]Hl��݇p޷r�8:|���K����]1�TCkH.կ� ���L0Q���f��
�L��(զ�lG7��O/ߍ�}Z-��߈I��<?&q�����!^����{��̓s/��b|��ȻYo8�_֢pW�%��Oof��l�͇ܧY��������5��dc�@�Y�w��\ܹ���y�������X��� ����-&QBuA�&�i5�u,���7ri�T��>�$��`�m�۸�xI�%
A�d�uk�~֌rX��_e`���
��� ���M*��S�:���+ﷂM��cN}�-�4Fk�Oi/��nu��L.bLd��{0H$K'���P����"��)RE(��hR+.R�s��vlc��h��F�G��&�3�ڞ�?	�;��Pb��4�/�Ȃ'W���ٔ�%�����m=m(��i���CC	���k��v]��"�P����!4 	�ݙ`A�S����cem��oI���@r�B;JM�K���W����[��y����^�!�H��{%i�ik����������Tn~jj���ӗ�~t�g{��q��u�i���n����f��΢d�dﻷQ�O3=tj�݊�Ƽź èw���[����R�?�I ����I��wdI�^5~^�������\�ED&KXK9>5�S$���!�с�^� ��u�k�>���/���5�����g�Z���n� �ֺX��c�6$���B#e(�;0�Dmû�����\��&|��g~��"YN�S	$�H�}0 E�7!�֨8�`I^ܙ9pE'yx*!C�$��.۹�"+׳j�ڃlI ��D�%��q�#Ic�0wS^�9���"�eh�b!Ȁ�-L�d���Hެ0j�=�6b���<i&%�v�u9�$�����6�
xf.�J���~�r�l��{Agb"�&I6�f�$�VC��Ґ~��?0��Lw���O�̾�5��燒�C˴���P1��O���?��S"�B���7W퍙y�y�=��	��1� ŉ��Y��o���4�]\ծ�VkT�%2M�"�����5�q"c.�I$W�q�k��0w׭��;�e��6*k��xxw�eXM�ò��%Csn��e]�hf��c.F���������+�02g���#m��[ �@�H�}0ď�~y��ݦ���Yk��H�浉��D�������ݏc�{՛�$�H����O���'](���Ly̹i��>)�<�:mJ�"H8��evi�"v���f����-�'�-��t��a��ϰz�r ;���[Q�o���~+T&@���Q�y��ɦ��2[W�W�p/[ݟ#L�,��AZ�	�9O*��f�[�[)x[���V�����D13�����ߟ�7ܗ������"��ݺ����˲hV'�d�x�\X;s>Y�l�;t#t�w�G���{_hk۞>�����|���F�H�����:[�2ɕE�?����ar�� K�N���e�r�]5VWK��O�'t8��/�� h���%ܬ�̫e60�<e��	�]<v���700�Ս�J��o4s1-�u��e`q�7gM�d�I��t�.�d@J�.J���K[�V8�@uc,"[��BV���	��e��F3m3�dX�,!��V(�h��6	�)ibv�Z"��A�v�U%c�V��c!�VR���1�YTtv�A�R'Y����F��mW��%c+lh:VB�1�鲄�1^]�3��{�?�]a�w�	��2�-x�1����6d�!�aʽ�*4-u�)��W��a���q
A2Z�YɁ��\��_~U3�����.���ȀS%��"ڛ޸��y�S�6)�嵯;èq$�|0	bN����\�NA��#�zdH��gvfN�塀ON�^!@t��э2��A�J�!���􉔛Vj�Lzr���V���ҋf>�troG�aȇ/
��ْ���{T<N�!@H&u���L�i��j�W�U�=�7}�y-��Z���n.���t��i��,�C��ku��s�fqR��q]i����.���>�z"�2��H-%�N�3�5�Ưp����*� ��C�߹�(��)9pP�43h�j�ߛ���k�fKc����;�\�`�:�E}]�=�܉_L����>{��{#����տ��]O�pSC,X�mI����D�	՚�U~���/ֶզHCNN8��^
��Kb�rZH$��}(��������j�,cr�I#[_]A c>�Z�(q.�E�x
X��&/��"���� �U�u��MG�������������-I��x�n����Ů��Odȹ�{��xr��d�m��2LN��yf�;'ޜɆy	��y�<��\]Osq`W\�}��>�5�ay�M�b��(�34�ѳm�2���~{>�ar�g�74�(��%�>�q;��2є!���2�X�}� ���cD��������������9�Y��Åf��$���P	#ٯ �>/4�elߤ�6g=���	��I�����V�{S ?_c���q��_����'pc�Lbv��)Գ��7;ދ�vqzӇW�w9~��R�r펛��{_�<�T�j����,ms1�,d#cg��T��ڀı�x�dk�N��'p�	7�����˨�k:��,�X��� �FN����}[��f�Q5��6��&��O�7��=?t�N�Ue��4g������Ǧ�* ����"}�@�/����_FS#B�Lj�P�,���q�$�"�(�[v&s�����k�1 ;��kj�q��Lvv�O�<r.J�^�6���� w�<}p׀�4���l�/���qy�qF�	idA�k� S%��q��R�R(%ݶ$�#c��ǿ/�z>�5J�l��6�4�~�N�'��=�,�ybK�ْI���FT>��T��X��ɉ�����+x{�b&�%'3t��2��T�]d�N�,b��X���5JY��x�ǧE䘨q.�};+Dl�|rT�y{,�'�BY���Ö�����NoMQ�w��'��}Ԇ{׹o?�������<2b��b�m+m��F��Bw	�	cs;)�1 7�����VXt6��.��Ј%���a��	)ָc��u�m-R�8h�K��%�8uKCW�Ԛ�f��T�v����cjj���������!�H��	�����D���R]�ӆM�d���&={-6��N����d����헷��}��Y��_��iŚ��S���9{����/W�`9�u�ʶ�	��3���y���R��"Ă�X��^c)���D'.S�V�`��s^�͸�2��YS�-����
b'5�+r���zZ�$	�l����9D<:���D�A2B�^��f���	���$k$�����v����`��i���uLq$q�C�yo��{����aj�>�3�Y�˳�l�����g��n�����<|���L��J2O�s��7递^>9����&���9e�C�R<I��C�=7��V.�*.���(ij�i��]�j
�I�*��G9�n�\0��tف�*R����ai\��7[��,]��3E]2ɬ�wYYWG�M�L�`�њ�T��
B��5�bՖ[��	�r�ӓMf�U,1�!�3	�M�[�M�	�����e*ƶ%�����a4�n����U�f\몈�l%�2�TImM�4��JV:�q\�
F���(�UF`�����WE�r��^�� ���$�@;��k�>�Ƴ�ꩍ�	Pj���13�kA�K����1��Ro����^0�;8r�c^�%묫å�{t���ؘ�*��*
��u��"Xn��$C �7��;Fv����d5��1 ��[��Ajڵp	0ú�4fwLf��;�'nh�X�)�D�gD����o��|_s���@�D=w�e������=�o���d���� �}����	L�^��,I����;x#Dݱ)$z�"[-

��W-�s�meK�YL��B«�rm��$�8�e�~@�MJNg��Ù��0e�OI� �w�H�f���vMԻt��?�Z �S��@��g&�m5Qcx"c��{}����f
1�Ha���~����U�)���O�6�6�%ǜ��n[�i]�<�\~i��o��^ۧW\ζ'=�;Q�=�bH�rm��u1 Z�^ �cٳ �'t�����M�~���ߜ��ڍc����>�d4z�1�'N�r���A�B��/z]�hD[��G�^�4]*PP����^��4�ҭ��ÈC��53$-���̄���Gs�Rۼ����	-�{�<A�X�I��x��G�<W~��Ym��7� I�ׂA%��ȃ�51!L�8�߿'��E�3�i	����G7Y�#�D�Vفb�7e��L��D���
��{�=����1�/��	d���ʷ.$�F�kK:�A;Q9�6&SS��rЉ�Ȕ�=[��Cè)�.̝�v
��s!w���2@���I:wT1�%�+h��)
���vsNa���YsI��������� ��7�(�WNþU�n&Ѹ��W=]���^�^�������E��v/S���k��_r�_���O�{���{����m�j8�Cf���+|}:��Q#�ٯ,�#�o�r ,�)����h���b�w�XQ��$�o3��vM�:7�V�?F7ܖ�Z����S<��"��X<�z�`^�.Ex�n�:=�欀�t+��<��O�Ӱ�Ҝ�#&���u�n�u�n��I "mqO߿OO��>��27mC���"�Gz��)�I�������._ �*�O9���8��kB����y����9��+�\�f�]�7)97ު��7�=���Tor�:���?xyg�m��s����,Y�S��h��~��}����k*E �OmA;m{��>���Ibc�1�l�o��&�C��-���������n �0��i��ǯ�ì���j�����;�x� ����`j���ɚ9b�qyy�|��d¾<��u���{���tȖ�@7�n�Ļc�z��\��M��x�{��ۈ�b�{ҥ���y�ضV�Y������g$���a���=wsB��u��ɾ`���w��o����=�۞��}3���=p���~ÂCH�>]�wv�;*���,�8쨅㽐��חg�!�a���^�6�^FI,'ٔ�Ou��
���gw=��;�"q|����p QN-��pr�!Y~��=]�ȍ�����Ĥ���ʬա�)YQ��.[+P��T%�F,X̰�f�̫6����T��9mK���ɩ���������u���������������uDOiTDQ��Xi*��}KȰMڈ<Z��)E�):K�QYR��MΦ���'O���ǧ]g]||||||u��ܜ�����*7q��r(��ǓB�(,Q+E��)kX��f�pc̞̚��NMΧ���Ӯ���]u����^��q����
*�A�DEU�F�;eE��VF"�Od-Q�X�vٌ��^�	h�&�[��%F1�j�,X"E��m��`��Xq1ȑx�U��b�(.<sv,�O"V�"!��(��m+<�
�+��5U�բ�,r�A�`���E�*26��V�Zʑ�i��,墨��E"�]1�1P�
+�!F(
(��*
*��,m(�m�[h)[lm��X��ȫZ�uj�U�X���jшaR
�����AA@Z���bͶ"��d��[lg�vFj%#,B���!�Y�O��)"���RƲ�}�oD�����N�umӫ�[QGD}�{5��v���\w0�e��;O�LCJ����&���S�t�BJ�����1'#
��
�D���5�5��\i㛬 �X"*n�@�4C�"�G;���	�Ȧ�C�˿��L��c��y�Ӷ�g�z���f`	@��q^ܐAg
�'Y�&!��P���}��Hd\�El��t�B��	?'�Zjza26T�v�J��s��V�;���+�u��9$���0P������U�6����0�ʴ�a�ך���F u���ޒjC�q�e�[�$�$����P�9d�
���&&Е/���r�ϴ����6�� ^�-,@� �1k�۱�������s����Q���J���=�1&�T�ح4��ɗ�kI�À������'�q�~�@�8��X+Ϟ����5�M�����E�/~�M���8�o;﬉��h�!S>�;�Ǡz��!�x�#1��YS�5��T6�SQ22bC����D����yt��҈I��bCa`��]��}���!�*CQ
�b>���y�VAO"�ćsY���!��52W!�$��%���Tt�t��3P눷�w �>Y�b�w��6��~01����[���}�O�a�w5�ie��H����N�rƑ�
CQ��!Z�|�������]{���umӭc��c�CY�i��VT�$�Ld����S�'d�u�����H~a*H�N���}4�߮#��Aכ��D���+/Y<s�S���Ɉ�� �=.���
#va��k؄u.�4�sPRW�4َ�?=��&_][sV��!�Xw��Pی��[Hy����d�԰12oϾ�'X��Y�s���[��$:a���k��Y,N�ɈQ'��f�m%aO�����o��h�Y�Op<I�0�Ϻ�P�Ì�g;U�d�RΏ�?0�L>�<�
���?FLϷ��7Ñ�G�~���9d�;�=���T�r�:}���� 7}_@dX1�g	�V�s4g i&�'���g���8ɸ�CC%L�}�q%�22V%a�w}�]g��C�����VAL�q�0������I�
�,
%M������HY:�}���x)�*��Q W=C�|�纽@?0Y�C�l�-!�;�2���
����d8��1�SqП�����������]��VC�Ґr,��X�E�����
"	w�J �b��7��jIJ!S�y�jrrC�G~y�w�]j*B(#�E`��]ki�a+Y;ߟ�Cl�1`M�>�>�ȆbB�9�~3�N�]��ܥ1j�,�왖��Ӿ0<����'����{��Hǧ���g�&�]�U�H�⪏W���m_#���HX��ƻ^"���X$��k ��)���ng�Y[���Ą㻦|/��l^^�n5Fl3T���U�%�+,4
�j:�Mh��B݂8ʰn�HQ����a:P%����u6�	��SmY`�Yy�4��:,K�mh�\g��-R��Z++-.n�J�VV����#c�G5�P�hL�W0[�[b7��2� �	��)P��ՔK5%ݯ\&��
�����N���Cc�b��k`��-*sl$���\ 5����<��n�AA��i[�X<���6�D
�)�7�m�Xq%N�3�w��ł!������j�C1b�,�δ�(2���"by�>��������i���Ϋ�Go��@m�Ad;5��淳���I9��/c	R�
�����q8��q�+,O>��$����!�n�Dl���5\F�x$�=���ޮ1�eӲq'L*{�^�0�B�X{Q4��3�N3���Ŝ�0��<y���D�Ѩ�28�)�7��s����$+b��*m�R��*�u�_�ծ�3B�x�<�p��â���Q�V�%	Y*}�\���D*Oc�0IXy�oD�7*J²V{�}�d���y���pw����G��a`�!���!;�w�EYdŚ˰��桱�B��Yi�_k�B�;���Z��|�j$S�Jy���NJ�)��O�ߺ%Cq��25}��儖�ٽQ�&�!�E'�0Y%k~t��O+g�q
�%�S"+�SCX��+�9v�Kh�M�\����	C��߻�]�O�ؔ�\�4�H ��D�	 9��@$jU���$���$��,�@2f�H���[� <MQ�D�gp�^�~����m1�]��e�ް	T�އQ���jϲ�E�~ś|���ӈ�w��_3ǬcU�)�kw'�~�\��>� �����/������}���L�Ec8w'���S$��w��l�W���k���^!!�)'P�A��l���-ə���y�r�΅緮�d�w!��H	�7~~�g�$��y��+�`�é�+$���o��HG~<6~�zw,���d�@7j�i�y$X$�t:�Y V�Γ�m���L�2 ?��(h]^��y�D�$��%Ky�v|-�Hû�R.l%�o2�IEvHƣ�k��/��mD�d%MH�mw,��y������"� �-�]�� �A$��:}�.���4���ЉQ���i8�r.��f���Ñ.��<a���Bu=��Ji)���C�M%{��kY��@OeP�T�U�$!�Ȅ���K-��R�I��ɋ���FZǍ�b�
N���h��5�{�M��`�m�D`t�@&�xh��k̄�!��)��IU�+s����`-�p�$Ó���{������x��M�;�L�)�U�>!f?<��F������IE���'���O��wL�LA��dg��3��~~�k���|����Me#a�籎u�����G��ZJ	�P"B��Z�����$�!�Y-��QUw�BN@$�b�$��t���$?x�Z^�$�ɓ�*�H��wv�;��u
 K�d*�k�����C$럭H,��V4I1n���o�� \p��Y�9\Hu"�m�=z�����)S;�G)��	$�;��0����M�
R��#n>�ߍ��mZ��߰Ӫ�\��WMuy՚���0q+e��6a���s*m�Z���}�m+��Ŕ�]��M�MH�%�]�ɟ#a몫,ҹ^�g�x����RMN	7B���O����j��t���;Ԟ��q:�h`�Z�	>I6�m
 ��~ Dn��R�]��0�{G�cْ�]��$��c�
�bx�#l*�.D�I%��! �"o�E��*=~`l���	$����#,���.L������
@x�.�Z)�{����\�;�W�wV�A%���@8�9Cv�>.fv爚!QS�<�Zq�S����,�/O���g��ȃ�r���!/kw L?��tu�>o~w���RJK,�R2�,Ad��+��yÜ��I�|�AG�RN�8-�?�@�!$�KV�L���V�]�29�!�;B�.gG�t=&LL� ��<��e{�t�V��$�I����P�]��(��.�ލ��3�H�s7WK���Z��ul'����� ���i$M�Șvwt�Z��@%]����0"��Y�#)kgxd����	!-�H�w��i��j@��w}��ݒ��#1y�MI&R�����  e�|�QA)�����&��p�M�D��:xO	;��N�z)c8����ɋ�.,Κ�`.� {R���A$��~2% /NԈ�w��� �S}s�Tuž�`a��$�nP� �8�L�R���u��E���	X�� �C̻� �	<HPb�
�o��"R�wֆ�{�$�=Î5 ث-k;��&Z��{}�R0�}�Դ^�Ż�p��q>}Bn��{�����^׻�i���C�p���I-!��R�ϫ�Ѹr3~N�h0��,TaO��b )o	��U�e�6�v�aj�~��o�eRYd��Y,�@�᷾~X���J��ct��6.������͗W5C*Ʋꅖ����3��i�`�䷋V�ktc6Qn���8[&Hv�]��j�#��L����qZ�+��?��(��m�LX�s5	i��S&�V;�K��I��])��Z35fuV�13)�k�	C�p�٫- �tΑ�~w@�<n"F��ke쑬�&Ym!�b����*�U�IrMw��������	������9 H�Q�o�r�E�Y=�ljų�Gh��\����e�闔�K:t�.0��e�� 煛�;�Bw��'f�XN�����!�ɝ�hH$	.��I$�]=�$�I��?��8�>TC�@k;��]f9IC�
���$X}�� 3���]uM1�H�N����K�Nd96J�<��@�ӽB�'�% ��%���"w������[��5��	 �,[�4)I0I��@$����4J�nbXa(.{�D6�P�	�<#�$�uO������}N��,��fX &�;ʫQI$�ɼ�$eN�-�yHW���z=2ֆ�\9%�t�7��-��7V��0mZEm����l�fp��e]Ȝ�p\D�x�!x*(V[)z�ҋ&)2[9�&��w���� ���O��;a��\��e RI�Nu0�^�A9��AG�RN�<�e��d ^����=b������TͶ��}o�����}��[��DקI�Nz��c��W�����US�B��	���@a�kd��<<J�����
Q�@B��������[B�����x+gE���^]�Ґd���F�P��Ko��tDxb���#5ӆ�NΙخ��8�j��M�-SJ$���\�$E/Nt�&�K����Bll����C����֐v���3"�x0�$�^��
�L�-[�Y��6���g��[ߓ�uf�R^e3�BM�k�ⴄ�i�����G�#'0�O�32�]��0h��諡T�$�r� I2_9L��\�f��$�wN0��x�i�ͥԗ�9��#.�������:<�MX�!�՜��<�b ���*�ME�.�����A\�L9՜�k~hx�3w*���d.��P�I\����PS�	
�HB
���g��R�2U�V���ې<ƉLC��^BD��|�2�)+]�b�LNGH��$��b)E:��<��'=>j�|�ã��2I$��}�p^ȅo�)���l"ﬗ�egݲ��=�1L��DQ�˞^��h���l�P$t���l<'~�}�N/�<d'Ĳ���
�J<<@HHiF��@P����֘��y讱�6}���6�PK��!�������]����w۞�7϶��|��0%��wu��&IC;�Y��<�I �gz��^<])`,�|Mˮ\�lu:w�ss]hI��D��IEfM��@�����(�dJڗ��N�^��H
#A?OP�J��bX�W�ϯ�|
��+��{��/� J3Bݝm�6A���[�q��*U�MW6�~�>��vr.�[ʌ�� �w�zy�R	����RI�ό,����a�:_�*	Edr�������ی��&ClL����dR����e������d�I~�̳$��ց�4(W44<%syv%�n���z�Hg����!x*$��σ��%}=4�x��η���LØW\<�I$�vk̢�LJQ��$�5�!h�bF �1��s�+j�fLxH�Q�o��1$�#^x$�$�{�@[��$�-�xl�������ߨ^����.�11���n*E�̞����'�������������"��v��6Ȼ=��A���
$�(��<g�#�)B�R��D� (
R��/���v�Ro�I;�{>x������O׳F�"�J϶$B�_�g�2(>�I8%���dC;����B@&��[WD<�5���{��z�r�^�V�m��	��">dV�b�f�i����6��+Zʇl��1K�*��@�;{��xw0�/>�v���S[�@ӲN�n]��e=�K����T�P���IMfP�^n��D�Cü"�~�wkU�P�SO���>�����h��ƀ"B�6�cXw%Y��$��7ʡ��#C	���)0�30�<0" �����E�vD�H$�Q뮽Ⱦ�������;��$���U��P	"ɱwC�I ��X�dਛ.���l���������C ^�Ѥ�%��a�$H-}��t)ת��0M|�j�R�$������Q�./̬�d'YS:�R%<������^����ݔ*�I"�w��`�j1�����ʶ�`��30{ս�Ц��@z�D��HG�%������o�FgH�;��L<�G�k%�C�vڔ��\�A�c���9�s�i<.y��!���7�W"k�.s[�n]��#�(65��x���,�mT�<��:�@v����ۋ�G%6�����:�o�V�=�7{_m[7{��v{}����g;���c�.^�v,�Sfd=������%��Wp�:2撹��J�
á�W��B����<���G���%�tgot�΍�
ɾ�/���0�x�R����;�&�{h͝Z݉�"�������R1�f�3� �����Ř������2S�~=���=��u�����k�����
����4�sپ����b��Vt1��ّ�gs�_�Ő0�´ h������iU��4���Ł<m��o+���{m�`��&�������KƵo>ǹ�V{5�W�,�t�g��ow�2��/`��][�2�`�3���듥���ۚ��\Ͻ3�������t��.9���{�OsT8ߺ��L��4�k���=*A���@Շj��)�P�=C�h��Z�7���z%�8:Mm�yL멒w�B��}�q;�u�3=�}3�mҸ�~��@�7�na����CK�`�H�7��k7��E	}O��ˡ����sܩ#�s$5��u�c�ሩ���w$7i�����LD�g,I�M0<�A V�A`)E�&F�M�:�t5n]T��B�%寎��G�$�/cM,�,6�g� �ɫ7�O%���Ɩ�4#j�P4��L�+�Ų�����w�G�����M7_E-��n�>\�=m �J9Z��7��hl��\q*M�;V�e�]�͑�e�Q�ut����yꯣ����v�&Y\��7*T�q*C3WY�9���Խ� �^��X�*r�=YAUQ���+`�`�Ƣ��M�Z�o���������~��G�]u㮺뮾:�ۦHD�Oig
,�)�Y4��������
hi��ǧ�]}����>=:�u�]u��׷枪���Z(����G���Q ��>�p=);MES��ۏO�������㎺��]u�]{|vw<Ң�L,TEUN5��(�Mw<"�����''*��V
�]R�,��F��
�EPUPQ�(�5h�X����C]�b��Q��q��LXQ�Y��(,U�QyJ�S�l-Z�(�Y����ʔ�En"�DZ�)QV-e�#l��J�L�a�#l
�TX*��,���t����k"1E�D�%EQD^�a��X��1b�T��#`�U]%V
*��*�`rA��T��gn�1�o"W]�W�||�CS.���i(K��VZjZ�����c���1%ɍ.�R�����Δ&ֶ+h��L�f�DA�.ٛ3ih��."�[,��E��ڵ�ꃻPļ��Q��Qа�5�^ckm÷E��7,{1���;VhM�H�ykY�lD���c5�%s+�����`b�˒��A�j��:�,r���뛜�Ŧꪉ�٘�Xju�EL�Eе�lZ1JuV��uT	�B%^6Y[�������p�b�Ks�*�i��Ĕ&S/%K�����5�\fV�Ij�h:�Q���)�rL�a�t6�(B��B�Қ�*4M��&��f�k��
�x5�� JS-�]K�Q2h��bF�zi��)��:�	�Z"�IjQs,��쀚��z�ր�p��36�
�H�]°n�Q�`j�����38f�٭����T��j��\BR�:Xb*�-�Z��h��Ǝ`"��N-G2�gk�A�k3(�z�&X̊#���)�z�f���4[e쥭tR�5�&,w4�[E
�f�z�X��q��k6�Ć�<hsӜB�1X�G%�\gu�[f#- �6�;ė*���m�`��CYu�l����e5��c9 \��+qlڀB���4��k�&%�0Rj��iT�2�یܡ��U1KVmZ��+n�B&U-�b˛��j%��
��,q�8�ؕ[���k0,����C��0�a��/e�Zr��iW��ʔn�t�ƫ��n���,4mVi�(-����f�*L����h�Վ�f/a��m�bʚ�)[���X�R&�,]a�m�1#e�H�������f�,9Q�Z˨h7G1� n5�c��%̳M,���\���r��;6f�7*�\䡖&ٚ�5�R|�En��r�fP�9�M�Ͱ�		>����3�Q�3��*�P	D��q��/�pY�V,�Ia�S7Y��ZM�����L��&�T҇jA��%���Wa�y!2K�-0�	��WGb����U ��mv���o]KlȐ55A1�5��V�Z,��Y[��T
�pL�\9ʹcR&�>i��F�c��,"Cl[F�p�;L°��`%��@%E�0,����4]>�O�˽D���4mWMM*l��0%n�%�-Vm��ظr��ɐ�i~���b��ߘ���3F��G�:�I ���^j��f�3�r�tk ���T$�)$9v�� а%�b)�SK��L�;�sDh:�Ⱦ�y����	$���r��Z��D�d��ƫ�Ɉ'Ӹam��JCv����I������0�����I���v�z&��01�a���'g]��! �b���L�L� ���,��<m���%uܬ���Zv,�薄��whhw��2H�
;z���������p���S�O�o���;�c.fn�_����t���>Ɋ|Dx0�@-=�m�6jI5���,PI2��T�z\W9Z8y|��,5U��]'�[�y)�sL\홳�FL�!T��Ιqf�(��pY}���ܥ�R �����H��K��e�$��N�	�K�J�z�0�	QR�	3$���2ҕ5x��3���&g�D���e����}�-����U�0%ܣ{p3�Z7�{��ճ�h���[f=��M�q���U�I>�� gh��*��o���}���~3��3����Yc(HB��?o_������[�2Ō��I2���*� �x�xg���<��%Ҕ(x0��z2Ҽ��;���&� �IO��{VL���,Q�h��������(���IC{��P�i����4O�f ���Kg�߳�N�WJTJ�vLO�y�;�4+�n�HyoK��ﮐ�ړ,g^O�D����m�b������p������q�R�A:ݭV�.x�d$U��H����/! ��/yQ�+C ����*�g-�P�q(�F\-��:�˖.k2���&�m�j3B�,��d�k8w&#����(��vWM)$	&��/�g{�}��>ll+~� ���w콡T�=�XEP�!D �k7(��D�ߗ�o6x�:�])2I ����4@6��e�%��,�����eHU������҆t����]��I ��t9��I[0]؆:��<{���g�y����o��^�w6����ǳ�qj�&{P>�G�����h��q��*#2
��|c�7�|�����,��3�x�A��x�� i��v��U��ϒ$�4\����%�bH|8R���Pim.�\�Gk�[��JszhH�3��ܗ$�\��3���\w��,R���t�%��`~�� �������z���y��ɊM�YB��@$�nK�H�H��eh��fP���d.�@� �x��ʈ�mjs���WE�2��Yd�����)x�J{nK�H$�Z}�0�	&H���2^«���݅}^�'X��	,]2�<��ILie�q�;��7�� e(iٍ٘���2{����^$��E�t��I- =�d#�eA x�r7To�V֎�^!AB����f\zfa ����帥�]�H%�ԟ�FUې�e�+�]� R��� 	As��iiwkk<�a�x{�뾚�9='���8<�I/El"H���S) �	f�V$������II�ۿ��'f��î�M��򻒰o^�6F=�uzyR�a�~{ٻ=\��؃�����X��˾��a�p�		�u@*%�2�Ic,�)HB>̫�����%��A�<E.����W8�߭A��H�}Y4�^n������pA����y	E >r�D�uu
�A�ʱ�J�����~�o�b�WY�J[�IZ���¹*�	���\�m"�hc'�����KM�'���BY���P�I%�]"i-�>t!jk���2�N��yf�R�;S�D@�s�j�H�vz(ӳ��9*���E�>�is,����X���H��H��RN{j�ٰ���2�� �`�9�8p�DՅO<�y��$���H�̬���;��h@$��z��R���B�&��6�����D�臚��7�j�.Q�D�����
��$1wO�7;s�qS���Z�JAX,�y�!(gOU~w�͛4�@$�s�D =oV�1�њ��+�:A$�U
��.��l[���n�k�2J��5B��m���?{�~��E��(`��8��,;�v�l����^ִ>�z�����G��)���������-����<��|7�o�N��}� FX�	*B�2�@���֖�2l�k]�f���L����WP��@�En��pL�a{h�T"�	�-�;]���-���L7�6ᙰe,���K5s31%Tasf3\V�fnŢ�l���a��Ra�֮�M	M�̯'#YJ�)4����Ѕ�Ď�@1���2�@�풳:Ya���u1-����m�r�]��M�➒89�lݶ�"�݀E�[fi�Z)�e^q�&٥����g�.�tXMN���<�RkgwK�vh�I �e��/!,��b��MGUz���b	��Y=�©!�I9ݚK��a�˼O����UD���7����,@��u|��MFl�ԓ �/!$�L�r�����r �6��v�2�$��w�BTL��]3������4?Wu�����gQ���w- �w^g���E�y��=���PˆH��zD�J�M��/!"�u�y?E�]g�"�zrQQ�:�^��	9��e�9	� yq���$��Rң��76�o�1<�,�ۤZ�z��>���q�)"R��R%�P��J�~?�ֶ���h_�X�ug�7����	�K����ͱ�L���fT��c �'��|��U����g̕^tѤ	�{ba%�ϯϰ�BJ2.�8�Ymש��ԡ���-oM4T�t[zmA&S��qE�����	2W��ޏߧ���R!\lF�.�������w������ˌ���o�w�Ѩ����"(�NJA��xN�f3�<5�wmEנ{=V2}�o��i,M�?����hbɀ�(G��(O�*�7Ϯ��4JKt<�d�?,�S(�	<O�)߻��g�w������H���2ВF�c��I���cI�H΍���u�/)���P��!H7G-@%��9��'��f�4^�q����q\Ȏ�K�������gv,��=�I��ޠ�}>��T؈���2��#\�3�����=r�)$�W;�D
Fo�=>R�]ᙉc<�m<��	%�~R%	 ��H�Q:�$[��um�:�+r8�4LKkb�V��m�bk����)�%[O��{~������^�堇N�
�K7�)�ܻ��H[@d)�yH���CK�/9bO	C;�<��J�:Eճ���u��XYo<����u���1��@��M	.�]
jN��*6s=��s׮N�H�ʁN�!�@>��icJԐ@.��ӳӤ��#}w�ȱ3�j%u:J��Ԛ��+���<Vt�ßO'[2�Ba~�_���vV1_����I/gڼf��s��P��������֒�u��2� �B �a �@
H'����-�[o���{��]�u�Ʃ _m����Bx��jOT���c�z�
t����@J�($�I��t�4���.X�o��|8�xH��RҠx��莓��(Ql�%u� RH%�� 93�8�c��Kf3��RS$Ol�R ���wK�%����.K�IHO�Fԗ�RC&�i*�+0��@��W\R�� �B.T8.=���zp�q=�kTW*���~���i�%��^R�پTw2 )yō(�$�t_*��$����Ñy�6^�ϒ(z_��هǄ��ш9�k��r[o�קJ���e*XW��%6	.�q��.=���җ��{N�Ҟ�:x|�X�I�)�����Y�2	��|�=-~�~l����?�^I����/!%��"W�U�9:�� �Kj�^�?f����t�_��\%+7�is?3���oK�I$������uX�W�d��#w��t�����X�\�Q��{��:�y/{������;�����?ym��	��Oq�Jw��Ap�/� }>���� ���$�ŕ�����ؙ	�$�ݚC����!<Jmד�.d$I����+�-ÿd�x�.�z*� �vw�h��H%�烍b�_<�]�l1>�:/#]��g��.���I� �]mt��%uc2�q?I�~��<C�<9]p�i+gwXcà�'�� $����)�Vs��=�$�Hb7�/T�I RHZ�RC�	3�ǟT ��0fgz�x$���MV��6�y��wu�f^BI�L���ZQb�$za�`��d��9�uol`����$��་Ð�>��h@ �'��-4����3�}=��lul��'B �e�엖�w$�~y���i��^����H�_lL
zE�K::k�^iw�����$$�I*��S�^�ˑ���Mo�!)I$U��G'Q� �J��;�y� $^n��ӳ֫��s��i�$�*�yHPJ��A�L�o����8	��%�(��{pi�+׭�����規\��qhf��͇
���̀���weXzl� pE���f�W��:<�x����=�}|�>Le�*kYEΚ�&�y��՞bCP��uO R����V��|޷� �HΣ)$���N���Y��'o���꒻7#-b.��ź9ݵRU�����6]VeKe���c����X���%���#��t��;;s�X�^Ue�K�X�k͵#btK.b���XmHe�^�7��A�iT�\	���h6k��U!�vm�� E�k�:�CEi4�)�:��V�$�Rb k5��Q�5Qvc���vP�5��*5�b���ث�˛�ai[��J()����{���Q
"G~0�u�	 Js�3�P �=]�0fm�v!��4ɓ�{z����w��T'��TD�zD�6���⼔��
�f}�~��@,A�oL��e��$su5��)�HoDE�E>7|F�������@ �#}�2����U~hjpW{&z�8$����q ؾ^Qxr@>4�rg���>�w.F߉ �nķ� �^�� 	%�7�ڽ�Q� �}= O7p�~)�3���\�H�^	%s[��]G�V]N����+Xnl�� �!�b���ɖ1�ǻ���=ϱ��+.r��[,�Wm�1ݩ�X]X��a*�٫ZіS;lƖ\�cU��}��$�N��a��M)�5l�bƖ��I�SX7'�k��0łc�OD�뭂T@)�&���R���Z=/�v����M��?#�y�0c�r���\8�-�O�e&�y��w��_p=�r�}�w�6�g����W��<g���e%������h?,W�u�GS�C���	$������V��'�t�����7�o.d��O~�-�*�+�l�����H���0ԏoT�[���C�(8��.�;uIx�8��"6+$q�f "��k*by��{�ڽ��1� eg@�n�Vx$(�d{�:0�cu� a���ɩd��{эH�d��fCI��x0k${&o^�:mZ�/�%�Y],ڪm�M[��X�Ĳ�5ٛjt�^��n��
�.�"g}25�� �A ���O���F��&f$	��Ǚ/Vh.����= {-�.�_��w�Gד�-{��A �[�8Š5"H_�ZA/���΄C�1 ���u��@)�$[�T��r{!�a���0�f��$Q�%�GJ|��,�>�:��ˮ�SS�����f@��)#9{���ٽ�v���N����c�S�����e�͵��ST.f�X��p9��R��3��ھ]���6���[��Ob>��ۍr�j9�z�v")�U�h��n�f_v\K|w�q�^R�C9m����m{�����9��щ�f̥�=.��v8���:��|�*�CԴ�������cۥ������ ��}��Ϸ=|.���{۹7�k������G�{:t���%��+�Z����9�w��PaM�ow�0\��}�!�����kV��I�cΫd'�ur��}.�{uc<�����v�C��|��R�q���]]�}�i/@�M�G{�r0�����F==��ƨ����[{ǻT���bܝ���s��o{�Z8���=�2O�?ڡ���=������·Ǧ�w�)�Y҅跩���Y>ߒS���~Eygڻs4jJ��S�=�{:M>��|�<'V�wx�{�����پ�yw(z{��X�GL�\65vTVol��>~FbK�Di����Ǵz�rf�����(�v���D���ۋ�;6I7��2z�����F�Gw^)2e�1�o���Þ,k�S���n�5BO�=Oo��q� u���Gt{�����ٗF���8���)�Y�|�Orp�Pg��5F!�မ8�x��n��ݘ�.s�ô�v�Fu@��8a(O/R�QF&G���Z�����޽p\c1���عh/]SI�Iӎ7,�W�o���TFq��&&�%�Ǥ�1�M:7cG�T����3��$��$�	��ŀ�*h,�,��(�\������ǧ�_o�ۯ��:뮸뮺��㮸k��(i����z��(�l1��lP
�����^:�}==��~>��|q�]u�]u�^�u��n�8�MBE���D5GIJ��f((6���m:�NL��M}����u�]q�]u׷��]z�(;���DE#�!ʚV�(bT��
�� �J��Y@m��e[�#��J���q����c�R<˒,U"i�X����B:�fXq+YWt�jG(MZAH:�i钺d�%a[*P��@�4�M2�*��+bT�T�Uh�(��n�2���r�ɪZbR���iZG�>�ʂ�"��;� nXQdJ��O\g�����x �A9������$�o��,$���H������Q0��#;&Kև8�	6����$�EOt�6�K��lmyxŏ������fH����p�}
�A�xx��L�y�1�w\�y<���TvC3�2I&��e���tCH^�/����kjVc�l��bM)����	IL������)J�gP����������u�w6L�� 2��P�Hb@+��mH�)<��Gg���� �S�,&��W�x*� ���#ĐKD�}��5]$@#f�d�`�}ށ �z|����� �3��9���u�\+���]�?^T�_�3Q�H�{��hl59�!�~�v� ��}.� ��xx�g��}���Z�bvCP)�b�nv4�8�˷��|�9.vXG�.��l��'�}�i�5��tE��G���/x������O�;}���:M�钳����}8j�^u�����<�֨u̼̹�?NFR 2�P$e�� ��u����;4�<�<<v�B��d�ï�C�����#D��ᬓ����A�������~��ϩX��O��p���M:YE�k0޺d�	�0�"CE�k&e��K�����O�򎰡�s=zc�e]�%��nwP,�lמ�R���)��2� I{���lu�s�ІQ Ƞ<�3�-̑��6�N�˪0�X��ށ,Ke�L�X�2�zG^���&��O�x0��UE1�Ά֯{b@�Hy��د^�{e�\�{�ߥ�y�"��&Z*��:F«=5�:J(�W�C]eĞd��ٚiTGw���M^��,�(�}[OV��)�"$]�޹��Ic�^�ދ�؉�Z����Ҁ �g�d
;����{ñ��
��3~l��;��sf^��%~z����/Y1��Dު~�jؠ<���w��-9���f�R���h,S��Ɖ9���<	myc
�>4��}x���3h��[���E��h6n�L�	����{g���x O�	^�o�R	�̶���=]IC%�M�#��%t @.)m��X03�����1�jlt�װb�
�-�LٚXF�.������c�J��f�0��W2͝���t2��3T����Y�n[6�����w.������c�[Z9%\n�aehk�n�����X�|š�)�lA9T6�V�f9��u�rv�H3tΡrj�ɳb�)3k3���3[���YVZ�T�4q������~��۹�X��bH$�����@����g��v]���$S�x�|u����܉-l�(��M�`A��� �y�j"w�����t�^�B�"�g/<�	��m_BN�2x&G�ޙ�I�1��MI�����{��<��7�~�$	�퉖��i<Bt�+��{��~��p�G��Y�ؒG2D��fIdS�<�χ''��WZ�N��+��*!�V��$�$p�e�{g��Ŗ�2�ݩ �r=�$<v:�.���&z���'㡣k`�gGl.&�+��lk�k,k�MXF�3;��C=z��A'��}�Ɠ�T	��l�@H����]���H8���	 ;$*o&K[X��N�A����h,S30�������3����AYT����@���B��լ��~�l������^��M�D�͕�����>g��3�z�}�����@;a���@>���x�g��y ����"}]4�LH%�_O�$;TC��d�O:�X�m�C��;$�Ŷd�4�&��H�d���`��f]s�	�>�Hb>�zdx�s�%��4���N�3�#!xQl��S��>V�qm�	�jX"!I[z�����@/�r��e*�Ym[(�Ԕ��XZ�HJ�hض6²�~��Y��8.�mzCy�'t���f����w��7Q�!��̀�'7�H�O����ta���ؤ��%��lJe}�[wS�#�#�2XI����g��Oe˦�ٗ�(@!O^��`�,�9�g[مl��ݮc�A��!�VQ�b;4������k�_'�>�MFȐO��H	�3�Ή�V���L��^L�D� ѹ�d�@3�v"��
�]�I˙�
|��FŽ�[I%��s�����@ �r��������/��a��Pm��t�\�$�_��n`mYy�#n"z�%���7��DG��=X�u�w�{ޞD� �}����<�K��{4OK�(X�\޽����P�1�@�:��,e$c) L߿s�A�����o�}�r@ y��+ó�&,[[,ڿB�ȍ�����!�/� �Ő9��&A �۲�����0i{��̒Ox����B<#~؍�$�׳4-�މzb_\C�cryz��7ۓ��h3�K �[�2���g/��^�55��F���p����$��c�<��J@��t�]�f�����SR�������IJ
Q
G� �Ji��2
�r$���*���O�L���C�@Cnmų,H�ѕ��t�xr� ]VȐo��{���7�z	$=�ْA�� ���6��O]�r(۾�b����y儂=7�8��v�s�O�q�H�{$	$�v}�$%��xC��ݛnW��O�������%2מ�$��3��:���^V��=P��P�x��Df�"�X淵~;}��kd��1r���WX������1s�z~���C}�q��{�|�뷛��e?�'鑔��B�����n�ֿ
k�#<��iX^��1��e��$	����=�;zD)�a%�@�H#)d�����]�?��V�	sߒ'�@�j�+���t��M��j�T2�5��fcoX�B~�'���cՄ���v�� �������p�4X��32I ��{$O��D��J
O
X9��-���}t�X�;<�Bny4�$� b��O���q:;Ԑ>�� @4�M���G]�N�<�×ޑ$h���c�h���͍�@ u��������Ħ�"�ֹb����duA���P�C��jv�O22Qx�$�oO�	�v��m	��\C�O��"��xp�
��/]�4��:$�{r�"�O?�$b	���'���b�pz�m�⬎����v��d�����~\��m���f�'��!wإ��
����و�<`���l�u�4����	�!�<C<�bSU�#nc�45Mhˬ�I�n2�2�Yc,	^��Mꐯ5s�i2i�FPl-�G`\�m��R\s��m)B;d�#����{�Mx���m+�r��.9��kepixD@i]f )�i���[K������f����\J�cD�"Bcv�HlJ�+p�16��
ثR�;gZ�^�����LE��F[2n�עv;Tc�rȭv�s��t6RkeLP,ȋ���)sc�@3�-S]5�5�M���t
�~Y�/�xv.���zzD��Z̾�$o{���k��#��+��V�jnL4��P'��I�M�Ï���b{��:a�2 �.F�Tq��{���c]1�,e�@_wD�ngze�]>�~Q���Ʋ|�%�`Yڷ�X�_�f����~��u�D��l��@o�����ݳ$��rww)��xs�	� ���h*��v
;Qfc��2Q�,� �!=�G�:U�.�؋~�sli��̨�,k�{�s�K�w���=sDr�$H<7�s`ܫ�2�� 5g@����D�(�+u/��=c�<Y�
����XR ;����æ�u�u��Z�L���X&c�7����{�����k��&�:$y��ӷ�T�{Dn{c�VИ� ���#�lȇ$�t��YxpK�x���� ��k��y	�z���C��X�o�D��F��6b� �?_k 	4YGN��A��!�.�=)ř�B���M�a�NO����R�X���I��=�Sq
u��E�2��dL1;(^WY��=FA1��;��*
	F!׼�2@ ���@��|�7�\1,Mvt��RŜdz�/q�r�At�Ǧ�Dt#꙱�:�,bjbhIbU�%�����Gy߳�Ӳ����-p?���� �$����]3L[�	*
hꈐ�Dp�Q4�V�v�Z �����&�A�D̰$��qqǽ��������y$a�L4�8�,h9F#uv^L���Ua�ˣ1�����K���C\��q� s	ggyd==�D�s��� ]ߕ��;���皑$ef��[z��(xDB��V=�&��L��h���ّ�	$�r�&X�=��d�@T����eweH$��C�#� ���F6��ˡ%2a|��p	go�aq�m��5��x�th��-��`"{/z�$z�ä��^ؽz�]�kfu��W�ޫ�п����`��u��x�����ec(���f '�����^ĉ���� ��Ӌ��A(�:�������7�����p�y�D�#.5��zf���J��v���떛� ����҂��X.����?2d�*%��`Ǐ9q.�����̓LvL�I��,@�H��1��./���ʢ�YO�u8SM��L�A�!�)r�)��,�vظE8�	��,�Zû������X��Ȗ�d�I^��|.ގ��G��P%�{e��0�8E�Z�������� ]�M��jd�H�db�<�=Vă�&��љ�� xHk��E�A���Տr7�萙7���Jǽ��yϾ,+a�&�d�g8�W �p�B�gZ3���@�
d�=HAH�wHҡ�k���Q/-݅�^���aUL�3qb�c�X�x���w՛������F��k���p,<£~�{"2E%�Tŵ�����FX�@e����{�<�L?{��j��8(�:�Y�L���~�K=U���`'�#�� Fo�D�'k� 0 o��^�=y�y���Xm1��Ub�f�V��BSf��pa�.�1�f�B���{��5��o��j�EZ'��X[��� ��q&"����l�@#;�CВy`w�CϘ�V��1��E���ە�"�`���d	$���2	������VA��� �N���z&<	��ޙ" I�p�ÎA�R䁯>x��ws&H�%��2�;���<:�C��Q1����D{��A`}M=�!�� �Dq�;�ۯM�)zI�38���Q$��2q$�Ĳp����D�63�u�mve>tk��d�FV�,{�8�'  ��B�gi��?w��x�׿�z˽w����f��L����z��9a	�_��N��o]�\��	�������=�D:P'��L�^���wR	W���u�[�t٣�.�j<�=�Q���)��0�V�vJ�h��{F�{���b�OS_��w��?*������FxЍ�xс����)0�Ѿ�M�'�!�8�����%�G��%�7�%����^��?v@hZ|�r�����9�lqb�Y%@.O��w���|�5�xK�Ǹ\5l��=�k���I�/��Ng���D,D�ɀz����Jg�{��%��z��z4<�n�YI��>ٛ��W��;e�@�F�̗�׻��	�����1ٞђx�Ѝ���lY��.ozm���z���=<�g�F&��ߟۚs���൐3����G�{�|/{/!�g���r�͙'i�}�d��#+~����Rw��o��u+��4:�;5h6�&�;��^ ���`	*����c�l�W7�uwo];�=��%x���B����i����*��=���\��S�1`�՜=}�?��ޝ�;�ޛ�����-��첥�a���f-���Rm�R���N4�B��:gM!Q���Q�c�0��5���&[�V���r�dn<\�7f��{B@c���ۜ�x�!ԐG���pd�%ބ罇ŭ�0H۹f9ũ�� :�w(�F�K1=J�L�8i����݃���xD�{.<��'��޹ʱ�D�;�+n���a5���^pko��v;�� .NL��ټ0ܖ�"��Z�9��=I�z`!�� ��ّ�z�f[��d;�X�(���e5�O~y0�t�<M.Ar1����юD�Ș-�_����G��!|xqM��c�0 -�c�#�A0���A&8�"��.���g@%�+���oG��<��x�����ʹ���<��^L�M�#�'$hJB�����f܂�(N�O��MM�'&���u�]u��]u���װ�[�@��d�A���P��xp()|{~8�믷^ߏ��u�]zu�]{{|u���)")JR�_p�)j��R�)��oN=?����㯏u�]zu�]{{{|{W�˅r9�RC"� �C�,��"H�ղ)AIM0@�dp���AS��Xi��>�=��
��R&$�J��x��i��YKK
�ŝ���PD�X"��q )*L�$�R)RJ��D
���*�2c*
DE&�d�)&��TQP�i{�%r"j�Ow"�QQ�oM�
±g��[T;�����ن��T��9b��p��f!�MY�Bak��]�L����v�`�kE����5u�6��`݋�̡*72���Ʒ����is��n[J��bb�F�ǚDU��T#��ɝ4l�Ƽݶ\Ոԛ�v���n�\˙��srvF��&
G����<����&b��f�BҪWJPc.�`��Y�����+�C))Tԕ�2L]��4�R�qW����a�vBk�9k��i�i�5�h�Ŋ��muaU��-���©�������h���{�Ѓ�ia*�ua�m#..Z�鴵#��R�̈́���Ghi\$�JÙK��;b�盡�\:T��!��D�EcBc1��֩W�'�ykV5X�#�M����y��a`����ZGl��%6rU�����l<��t�ہ��-���8ŕ�Ae�Z�2�m.d�̀I�k�4ġqnP#�q�&��.f԰��1�[(�k�fR675ƙ�`�$б2\�cL���V�Ņ�%�:�q3L.�����n��V�:aGk�X+'�1����aqtu���ц�i�&�0K���5�4.���
���E��R6�a#�����U�r�`��7T�m^��5by�f� �Wf�.Lbm��Mշ�b�+�(��)uk��z�����4]���6�*a�)�#a�n���%���WF٠�������AuP��iX�k�xZb[MB��	���*k�PE-��hcb��Z]1h��E�&ƍ����	\�n���R:�nսL��e F�+W�d4"��Zmaa�t���q5	(+��u%��M6Js��Hk^	�p3KN\lT��]h%#�Q������7r^VkU�.�l𺵛��|˕Uq��%9<�R�Aڍ�xx���Yu���Oc)c,e����knǬ����R;G(�HLT,�P�a1�эh���%̣�AV���Z�d.��n��e*ಱ�]��]*u�0F=��4���n%��Y�M�Hh4Ԍ��˕�s�e������.�:����ãY��62]�Csx�Y�.���FB�鸡J:�TY���9�u���*#\�rm�.�c6����%UX�����+u,.���*&؉��h�ne������?"�T"U1=���ë=2@$��MuFU�z�=X��]P�j���@p׾j�](t�[�~� o��K��Ͻ.��1��'k�e��7f8�el�,��z�����1�tRH��w.��<��˕�# o��)�5w�O��L��xu���֦L��	��3��^`&67K��x{����s~��8����7{�F2LH혓 ��&%����gW.=��$J��@�I�=���<:�|�׳ �$��@ǽ���1�!,$��L��Li	�;8_wK���y���u�ܠ�4��Ҧ1��F�1n·�%�$�L���i[�f��i�g�)�@��u:|r���P<a�e�@@�k)�Qb����'x'�&�XY�z�i8�S���o�̂tѤ�èpP�u"�GtH$�uZ�2���l�"�Z��{0?��g���e���z�g���x���?�^�ܞ*�.sʎ�y��!E�r��&�|�51ddœɋ&�bb��	 ��La�I-{�@��������F�ſ�L�B�A���q�;�r��Z:�,m̂�I'`*�oHȭ����#��S&�� �5w.��<��׾͔�'������as��.���$�Z��rWk�^߫sD��~�TN�$�i��A�;���a��^� [!�tsӱ����z�0�g���I"�2e��:��&��|g+���3�y�m��­�~lf�f٨GA`���ŋ�M���A��Ҩ��Vj�T�����`�:����{2�^tH$�z���eHOV��׫��7}4d���"[Cg'S�Vp�bZ�;KI7�ai�è�3�:9�Y0$���L��QU��M�끝�7�#:��H,�Oht��"U��;S$H5[�iv(Ų}�`y�ԎE�R�)����0���+�}����]�݌����<$^I�=���1���fgK�u�o��B���4�U+�~�����οk�Ա7���PL	���'_E��h����9O�=6��<����0r �.��k$��@�ʘ�_\q�WE[=A��$�(O���;�xr@�bk�$�r�@����h?�0�޶x�t
.�ew@i͘�_��������Q@��%�"�m��ừl�b�QIf����0G\�0a�v�9�Y���m��A0��nEG2�܊ � [�b�UG���z+'!w�N2z�e� ��
���v����B&��87*+,(��e��g5�_dQkb����9�(�n.�=1:��>����{M�ÿ�H<z��1�i��R@pn��,�$�u��'����ߓ %��y2	���,@8���r��B+u�����+�Ib=4Ԋb��FjG��+'N����j�i��S�?���r=(����(�O��R�Q�N�o��D�T���y!mM�8�@ǧ����v���9���2��R�췻�?}�o'����\�0Ô�,cwO�I;�dM[�b��vW\b ��v��E�:�����H>Ka)(_�#��j[�[�&A#J���m�(CF�Gb�`8�����7��N�����z�fL�7�(G�zKHP��o9��K��z��'�SDGjE���"�aü=�c�7"@=79u䑹���@"թ��I��֪%�W(�2{t܋���bz}�H;�*è2=� �ɕ^�If��P!�O�eV��Uu5"M�ę�; /��T���V�w�
1/4^/ܬ��m�����e�%����]�C���l+�
�r�M̔��ǅA����P��-� �O]�z�/=�\��r�}�ّ� ���D� FI�>��uQ���=4�<_K��q|���pޔ���+�[�
G��P3�"����@Q�����q,�u�yCJx��+!Q���uK ���<h�	��׈�Ul���J*j��,����f��4��?��u��ש�}�ɥϰD�ݑY(VfW��f�p7]cQm(mc�MjĲ�v2��:CM+&�&��^b���Z�d&����r���q1���k	�7��:j4��GS�in��#3]s�l\ ��R�3nGD.Te��E�,Xaۛ��X�\����κV�-�H�ІI�h\�ݪA�٭ي�������J �'!#�Z�p�,a6um��D�j"�b沺��#�x�N��Ô�$w�o%�i�#ϙ1LO=�� ���7w�ф��$��tH$�I��t;�xr��*�"Ky�f�E@Y��<����ٖ$��u��i`]�����T���V�(�耐*���s
���$�{/�,4 �N�+��LM��$����%��1C8p�6d�l�I�'A�����C������f�<[�W��x���s�	7�q$�A �ߦK�68���c��̈́1� ϯ�X�0l�;� �M�& ��.���"B]�y��r����D�Ā@$�\�&AL�;��y���K�����?.��O~�f2��(j�mt�j��4��a�=�+v���t�,�*V��Җ&����Њ0���d��u�̰$��a�$#:�9� #n� ��d=��ݳ��'Eܨ�$y1o1���59.Fб���Q�Rj,ݡ���پ��g�tl������t���W;�5�������3��)5Q�^5YQYW�8a���b�1b߅NT��@ܽ�%���� �Z/N���~��y�t�]��y�魖�	+��`NL�u�^"��IZ�_?SSPb��&Avz�����ü<�>��ޜ���R������
�G	j��>������諢/3m�1�Ȁ�XN��(2+e�$���SC�dwWsԶ����>jX�=����	�=����c�}.ẁ"q	c�K_ ��3C�R&
q�EÄ�li]3x�
WC�O��ݯ��9���)p�!H5��+� ��{O�o+ ���dL���L�*��4\� �P���Ꞁ4�)�j��8��κ0���>d��O���X�{�$J�I�����g��&`=��K! �H��U�҅1���	颐�^R�3;�3�ڗ�����4��� ���?5�+�߷����~��
����{��TǶ:�m��.?z���h����.|z�&�).�TDs[%�ŋw�q �gܞ"� �^�K�S��C�r�C�𹮺[�sö[��^� H��C;�w���=�7u���Y�$E�B�׉a����Ă ����*=�/C�ҙ'� � 1;{��1L{��>�����b*t���(�$�'.���1�C�����ô��"n���놉QM^}~{�K�R�5j{��s܄%�&�V�bI�R�e�fd"r2�o7��bL� �o�h�P��!DP��.dy�T�ظE��-��R��}��f���Iq�j�b[Q��.�\�a��G&�QTz�^r���W�hy�P�
E��A�_L�Q�U���L@�m{8� �gt��R	��i���;���H���]]9��D2��u�Ke�b��ȐNlG�3<d�iS�8Z�5��+�|�ُ`��&�AJ��Z{����7U/��DwT2�M=FT�z�d��B1X�,X�x犑#��b��K'.����zf@,I������ݾ�܂G���� �齆�	#�#�)7<��<QI^���-!��i��bQrf�6�����ڒ���їE�w�-�iwC�xu��鹐I G��2��v�t��oW���j�6��ʒ��Y'{�W��uxI�J��ǹD��ѓR��跗^E�<�>ف ��}�%���a�3DC؃���@���� �#�,�$I����=J��{��]NK	1��iF;�!�����
�O�wNz����7���U�"I �kڀ��������x��O�~lT��i|�<L"�a���
�GK�%���
�^ד ���a o]̍b�8ѱ���l�ɐO=�}s�8��ltY�����W�e�{N�g���`�V�9V1s���{۞������c��ٞ nEw=/xҳ�ə㟑`���<yI-�rS1a�p��Ė�ZV�i��(YJdZ��Gk5�Zqϧ�#Û�3��h���s)�)h�o
3U�T쒚�� \�9���^4v$4�e][�H3��aT;[a��v�i)nf^�V��iF4���Ԫ����/5c���6B�S��\�i��M�鸮����r��pl��9D2��˛�3))j��L�l�p�Vh��b+�n�R��]e�-kvb��Iu�zӮk�Y�`]Լ4���k�5e�7.\�a��\��������p�oۙ�B��.X�jof�U2y���##^����&����WɄ��y�3�w��ޛ�!`�fw9U^3�$AV���A�wD�K��`�����b��Dq��
Pa�C��@Q�]�g%����"�%l�^j!�_�Y�j���s8p3c�H����N�E���i���W`!�q�^���n�ś��i3]��ʹw��~>ܫ��I9�,�� �P�����B؁q2{�T�C��m���I>e]�۠@,D��"q���L']E�A�_H�+xY��2�������\�u���ujg0Iq��8L"�a���j��\�1dw�"HYwM1�F|z��׈�Iu-b������C����T�*��gn��}:�O'���fhg�Tɤ�~��|3�Mg�/M{��g��o�4Y����v���%B�֏�gR"TJ,�؛��b�X�УsZ5���馪� ����J������v 1���H���r��U��c^�$k$_;���fsZ��XH9y�$�g{� 榋�I���y ��I�xu?��m���ѽ��THᅀw�H{= K;$��_�������dF�ŏ�na���	<�`(���AiD��㏭��mwlu��,-� j�fY��!2Ks١�y���������>���\ڶ�]8@��L�U��l�Zh̗&�[p3�ￄ���W}��`�,I%����&��c��ۂ�8��n��˨�A}y2g3�<L"�a�9�x�s����}�Y�20
n�٦ K�g�I�K�c���5����g�^_��F��j+|Y�!9Z��T��H.�]|�B��z%sf&�?:��צ�Ѻ�^E���/xf�������83��'��&�WY����2���S����ɱ��#�J���������d杼��snY�������?`�+��Ry,>�`��}/�XjXF��<z(ݼ�'XGukye�4������M=6���X��8�_U�@�ܱӘ%+=����9�w=�u�3+� Wf0$?>���,�yyXg��\{��L��p��=�zz�G!|�\+Q���I��g��7��p������I{��I���6{w�]�����Յ�&��-��nu��_��L}|p{���e�Ӛ$�K�}ݾ�f�;0�ޓ�g�l�w�X��%���caQ�ޣ��]�-�dn�}���޼��yv��,��Z=O�iy|w�9@ߪ���:��q{�0���,l���ΛW��6h��{A+GM���B]�.�����������{��ǵ���=�	��d[���"Kճ�����^q��_�����p��x)�x��6۞�0��Fq;ⱜ8Vi����y�F���Y)4�h�����^�ybɷ.��ݳ�4�@�VY�sn����`:-�'^�L�A�{�=��w��^�|0p.��xL�;�zm��j��P�F�˯�y`����Ӆv�f8{h^B/\�0�u�i�c�����6�So5b�J|�17T{3�����$��c��b���Hg/�r���=��i���o݅�u���yJ�=��/xL��aZ��J�ALj���j�%�{}�ӏOn�ߏo�����]uק]u׷���I[ �r9�7�	r���օ��Ĉ�aP�8���^>3ӏOoo������㮺뮾�u׷��ّ�0��m�i�j�b �D��k��C�š�r��=8����~=�:뮺���]{{{}�K����$�'�.�Y����j�f�Z��̰�`其�B��F)
±EX����*�*�J�a���
����x��(ł�*���U����ʐ�B�EՖ8ը(8�1"ŀ������*�`T��c�(�
�IU�V�XUdQ�,�RV`�m�Y��dVa�֩KT�*DRAq2{2$bF3�|�z��R�z�{�O���d�Ɛ+[Y�w�T[c�:z��Xց'}3!��d�2Cё&I ^wD`�$yI ���l����!��`7�{���q�b��yC�d8��̆I�d	F%���GL��s��I�Q3ޞ�WR\��2�ƨ�W
�el���z���s�Ԍ���暓
m��	��/��Z��o�u��A3��aX�L��D���#�_���m��Ɖ@�}~�DP�`�yp9�<ċeBs�^x����J�H���2	$0�����V�'3J��	[���E�����f�:Y I6�d�!�р�s�>���I [�ORv &>�tK�k���AC��NU�g���<��r��˜�Ab�:E:(�f��,	��yqä�S�z��:P�o~����َ��f��?�9S��Ȇ�R�ռ?���	xR�N��7����_�+��r��� X�,@�$�: �&(�x|�\��S�*3�ހb;W�*�\�nW�y�tI�:��a��"I��"@��[���gxw�Hտ>ԺꎖTJ�j0��3��Eڙ6�]�1�km�5Jf���~��(�3�����u��q��1d}1$�OWt�=����}&���ӆ�&�쀮JD�H#��u�$�G�0+�s&YE��}�I��6���;�,��$U���	ۙ~9Z-UW��3ݢ",@0T<��������{�A ��`@f�q�Kpp.ܲ���$�r_�d��H&=v�L"�	���7�;*�~��VR6� Ȩ��Y& ��L�Ws��;�I]���Ј�Ι����� ��D'*��]2Ie�K-g8������	��ĉ�L���B�~2O�<-�VN��O9<z*��MNЛ���OW�)hZ���� �{'m�k{���m�Z�9����US���ii?�����g���ޛ.2s�1�x�ϋu�Y1	bBOWGH�E�����������:���)VR�P-㵀r���Z�*���V��yf��i-��<�O#\-TZD�9�Vg��p�I�ٴ��c�&V� 裠 �l���wb9�����ԕK)N��F5��8�4�Il�h��:�01R�0%�t̊��p��,�Ԥ[���k�\�QRl� \�h�Ҵ��u킬�V��
��#e�ѠJ��gJ�\�Cbbt@CZ���X�:aZG�����]������@$�ɒ	���8v{}3��_��c�>��H�L�o�&C=��F����
G�����Xq��[�6����k���Iݼ�  H[��AM����o��Z?���`8uB�̩I6�}H��Q�>��'{����&u�bC��&�|�:!�%�VD���ɜ
W�+=�$*���jdB�鉚�jB�z�Û�&s�g�[GG�`;�wp�y�w�����%��ni�!�>��,螞�$�otH�~�����y�lp����E��7�Ե2�����0�	E�֨b�XYJ�1E�ζ�<@�wqd��Sw�s)�=�)1D��醕}1�zF]�l�!����`4�ւ��]�û@>��S�(X�ng�TTV�z�慹>uU/�R?uc��'����5xr4v7����h^2}B�K�B�9�̛lq��F��|�T^MR���!�ŋw��\	as��A,K{��!�,ݑN0�ޮ|�$y����0���xW`߭�u��&$�B+�)R�~�W}��L��φ��A^��A��p8�ļ<P�*�s���oH$�=ș�ŉ ��Q!��qĘ�9�T�My2���[���}��-��r*zP��C*R�D�|�臦0�;�P��� ���ە�v�� ��̂��̒'��D�_���ā(���|��ғd�ٝ&��CY��,L�n���8��L�T�j^������tΊ�~�]|����LWf��<����%P��8��j�'��S>�����x��[Mt�u���T��sN��Wd7����j�ؐ�H�ǻ�o��\"xه�E�E/6��bEZع��� �{&{A%8>��p��K�;����0��[�{ʔg2p�z�{|{�I�vjgm䑒.�<�TP�{��p6]�:}�ꕡ�׈�9�fΧ��6\_�D�H����������=7,�5�zdݒO�	�& ��ç^��=\��I�NĒ���Sf��蘒�zw'�����7��$�l�F�b^,[y2$�$t�H[^�	ʚ�z�.�K�ѳ6�,�t�9����H2��j-%�Kʗ��BOw��.[�D�K.n[Q��٠�Q�m�v�em�V�1�9����.H��P�}��ܙ���K��ВK��X�����[�u� �	ܼ�$g�=�x�^.��HD��s���;x@����q�$� ޗ�@��������>����FUn ������	$��|"X�3��K�X�Yr�v֧ ���@�	K}Q�	��E.mh)��Pދ�����uwkdπ�0�d�#�1�@${�3��W�Yz��!R���(z|¾͹2���ە�;���^O�b���=�jcm�G2�`�$_�\��U�;�.�9P�꽼���LC!�����i�I���a(w0���{"X��ăH��� ⫁4މd��&X���ǌ�b���9�a��^yԞN>ۚÜ��|^Ry@�IZ��,v/HX˴#֎)�j�m�ՙ�,x���:�R���-��^�(�����}.�$�t�bI��d�}�u���o9��	��侙2��E��:j�ތb3xZ�ϥ\Lߤ�2G:_% I%�ݓ �u�ۧklc�=�?x�!�;��ȽcOo�ȱ�;�ȢA&��Eǣ�7�2e�bk�4�vB���h�ph$��w �������_y������8K�|�%���	c�x,�wp����֑���G;:g֜I)Ht��U�G�A$��_�Lf�ͫ$GTY�	���`H$�^Gzd I�;��z�~�C�g�R�B>����Lϊ�8�ϩ=�E�=���Y��G����\&�x	ȕޏ@w�I4'�� >�� 60�<VO4Kc�u��Os�����G(��b�S��/���q�q�o^yq=fk�I��  ]f�Ƹ�eҙ5�B���� )L�p��k͏gb[��k�Ŭ v��G:ՅrV�sy��bM��5�R���96�&Y����q�F�
6m��Zr�H0Z�]B\�F�X��R]�v��R�)]��y!��M��F-����X6-�{eR�@�#q-9��&M�M+H�ʁM4�u�J���r�sjT�fN��)Qu�>�~�߂WQ�M�
��Q�o�H$��ɖ>M�U!.\qƅ�t���I��$$�(xs/GV5и�29nH��u�O=["I�vD�,P=ђ$~�ԲzI⪽ |6����+�gf�:����^�qrZ��A&^8��{`�Ͳ<�l�otȖ$�^L���h@��]�D�P�{�x��#�wZ����]��bI쾝bµ�8��J���P$��vȑ����8��Q۱5;��\>h�wR힨�����l�v%�Y��$J[��d�u5�#	��@(Yc��ʚ�%�&�1bU1A�X�l�k��X;;hK�N�"�ˌ��Ep�BI��7�Ē�f_�Q9�d�N���e��X�e}�'�=�{�D:&�����y�X��~�xvj#�	�D���q�iwKV_墭��B�p��%����r�JD>:�3�V�6�'���uUT��x9c��dbF$}�Z�T~믷����}؎"B���x��aj^ru�h���Ċ�&ZI��(�%��台��oFo݄�X����$��q�'Ͼ.�4 �0�JytMm!����39ҭ�8$����R�9;�w!W,�cU=2W��W��E�*�����#��2^�n�G:�����[h�3�d�	�<d&X΍�t����=��σ$�"��Af,g�1�lh�h$6�YH`����0ݜ�2b�U�!�����YÇ���FXpɯsK�S�����$��t�5�j�(b�O���wA#�#�3���i!'r�T1��X�鐴�Wh�zw��44F�$���� I'jUp�Q����9�=�@V�9e�9&!���o��ȃ��+��d�\ܓ�7�+�k�ECb����wB�@���o��螞�����e�gk�y�.��wHB�J��9׃����Y�#�F��|D�d,@�#��9�>2�&&��I� rl����vL�/X˱����"\
��,�d�W�cLF��+d�s�{v�`'7#�����r\BydTtȐ�@.�L�9�������	�Z��u�$���7ީ�uy��ӼB�#��
�WZc����du�Y��fZ��T�6�Ԇ�QC����&�3�q����p3\��Y"4���I� �[����a]mlh���@[�0�r�&Ijo_fp��!����"H�$�NoeF�lm�=�'YG��d I,�]{RHT=k/���DSL� �a%^*��8�%���%�_�fv��<$�D����	;y�$�A�ڢ�ٶYt����:��]�\,�����H$Ez�2 l��9�v�8�����M�y�����n5�����}9I3�2ǯj�Ԕ�6����{D^Y�Y���E��=�Si�41X��i�bI���[@�H�<P��L�bX����͎��;�:���Iͮ���d�r��<�D$�r4���a"JE��}K��% �u��E��;A�ĺ%VW(m���4QB�	�����-�"h��}lp$����
�N���Q݁�^��G2@����v���D"��${X���K��i��<��G2[�i,d6:8�.ɽm�"�ė�~��ۯx�"!�+pKs�䀉&�:'�c��1����$�ؙd�����$��j�W��J�{������>U��u3,�$�o��I'���Tl�s�Բ�m�;��-��`����C��݃~��A73�v����0i�S����/��j�2�	gM��:1���l�*�B�u"����^-j�?��"]�H�T�US�0�M�g�=����6�5�/c+������GR����q��7��E�t��ͷ�Ǡ��W�NǿqQ{G�|Fz�bN�����,g/ge�M��&���=�:��x���]b���3BԀť�V*��;�C����I���X�=�_�ǦrxS[�#؀.�gW}�w1w��`>fܝ^��5r��x*���{�a�;8�jTͤ`�Z��%����w��� ��}�qu�=ǵ��o�qM�-�{�+F�[�u\�b�rJ!���<8��x�Q8�3X��6��r{��%Jot����o���7���z�����Y�/0!��I�c�r��,q�΢1���jygoz��P+�N����|�־,��7'yiغ�7��� �ρ�(3&������twi~�����Ņݪd�����H�V�7��A��^�-�3�Z�N�����'9��CR�=�p�v^�}[Wzv������۞B�ܡ(�r�mg-{��Ԣ�}^7|����w
�p�N�������Q�+��j^/Ǜ΂�s�徾ݾ�.�o;l욧пw��Y<��N]`ـ����D�U�YN�>�f�*��0��N�;�M3�`[݈�l[\����Z-�JQ�/@�Y	ox�� R'=~+	~%-oo�3Uk�J�4���&`�-�8�'7F:D�3��ni��}=U:��zD�d��s�U-)>
�9܅��ap�1�u�A�*9ZCNь!���:���s��4�>@�d1�
g�5�s�]�r�3ߌHs卉�OR�%�zy�S��kN��g�lDe�`~y�|<�5g���c��>E��؁ z1�4|M�Uو�35��Mou�Ԟ^� ���R��E�J�Z���c+Iγ6�^��:���ۯo�뮺믧]u�����x��r��zƑC�Qb�#P֩+�;��O���ǎ=��{|u��u�]u�ۮ�����6:�"��3��J��d��dy}&K7:�N�����{]u�]u��ooo��.�<"�OXґ���Q@����%��ڑTX(�PĘ�����8�1B�e{d���aۉ�[g�P9���PR)��%J TX6���l+-�WMTX)X�E1�R���R���h-1KJ����f�n�i�X�ݶ��Q��JD��HT\eV�v�C�M�eRi�-�1����դP]["��E��4Պ
��kEs-�ΰ��f����f`
��`M��-�%����͉��L!+�t0��ZU0�]Z^F�Z
]�[��EJc-,��;06*�9sL\Բ�����d\��̍���ȴ1ja��:��v���+�
&ҖR��;������k1fc�6�Y��v�.�bQH�� f<F]�+44���s������a���hc5y�h=�L���:۵���*f�l�BR�<`�V9�&����e6p�5����qd�$ump�m��!h$&ɍ�չE���X.ʷX�Y[*]ԭ 2D�p4hٛ���Q��X:�V�4��XC�+2۬�]p]v��F�5s*#i.��-��2�8��j�n�;j�rj�n�^�S!m堲��e@Z�R]4�]0 ���)�P�Y\Y�h�7��`�nP ]7�8��l�b͡�&�8�%tN5wgavY�#v�(��n����MZ�6*�f�IK\i	R�Dt���RU[[��T *MGF,٥� W��:Eγ*:-��l��v�n�!���R�K��e����Ҕ[�ݬ@ NҶh�� k3�%�hTk5��R��\B��T��Lb�c��n�w�e�Ԍa^�����&nl��L��Tlf���ܥ�p"GM��͗
Ĕ�h5Տa0jjfV/V�&'�|��/�]�)�i�]I�K%���*e�	WQ�k[6u%V��7���+�qcݳ��1MŔ��"�Ylņ�f�A#qyc!X$z�W��%�c4!����ta��6��n�VT-��l4T0��-q�h��#׵��9��v�؛kv�3X�,kIv��$ɢ��mi�j�m��\�3.����B.�c�T�v&`���m��ҦuV�\���l������Y�eh�c�o��]gN8�'��74�F\$&�˰v�0�:U�0ن�[B[�I�sŤM4`
	3˔�^���5� ֛Ce!�j��ဠKH.fCW�[,��[�*)��j����u��3f�B�[m��>��o1f�F#D�1�����p�ن`ҽ��6�T�b#F��kJ��J���!j�Z��u��ԅ�(XehU�ۆU͛J^�̔Z�Ye����`�*m�s��;��9�L�l�12$�M??$�}�,|��{vw��{���HB��q�E>;���'��]��AS^���QÑ3��&�K@���	6��I����S��$c�����ݥzC��",)�【{��$$�a�Cu���qS��f�$�-�4�"@�ޑ>��!��kL�o����������)�y��A$��޵�Dm��&m���%u1	8w��lzd�%���h�7<���A�b@Wq�H'{�"Ic�{2��ǑZ�c�XN�	%�\ԣEt"���(�FZj�:�l�R:ٕ)X,�%�)ɮ�{A�I�DC���I<���VI.{�0˺�)��/R���A�Ŝ�Kb��2	j�	�P���'�(���AA���l�w�m̞mu�o^�������Xr�����G#<5.p�l�Y��Ψ��d:�����SO���L��dg�z�F��:�U{�>ggq�ީ�X��w��Ϋ�n��������'���'̇��M $���u��+y�vT#ݙ2-�hC��R�Q$Ǜ���C�.b#�O>���n�-��@�"I=�u�SM�GJ��s{�=x}���s�\���8���m�qz~�� z-�S�z_/� �xx�c~�I���$�}�2�p�<�ĈEIR��tU�-z®8�mnU�j萆�{c,e�Fikv�:��������:���$���� y�eͲ���P=�'/}]m�
�N6o���P��Mi�^�ߏfx ��W�^���} jd�2���L�Xy�=���&�p����Rz��4AP�𢅞}�����Dt��}̸�?e{u��D�e}��lڳ��^���|i���0��G]��g���⽯�q�7���_��ب�3cb�1b�e5s�Jb��{"X���c�w!+&�O"�����bB͌�	3��@6��dk;��t��Whf������S��r\�E�3ף�%�w�,����l��7�p$�|�d�	��;��3O�ܧa�}Bv.J��O��׈�Y���v02�⭄ֱٚW"[����X	��	�����"!�1ג�X�{|�X�	��5�er�v++&儂	��� �U�������D���zD�m�
��[ޏtP�A�ϰʍ1 ,��S�|O�{|��1��گ9�ۗ�H4�<C���{2�,\=�tK�#���{�6�X��u��%�7�!4�+{��>�F��h�JxQt���ӑ��}$p@��� �-�Ȗ$u��O��]
0$w���S�D�>h���1��-��s��Ͼz�'`N��on����('���9x0�^8��&�7�!�b� )��d�_G�;|�w!+&�OP���ˣaYs�׹�^ޠ|�^�4�̂+{&A �{<��ԫ��'Mga�0���ʆ��v�l4��������\�4Z�;]F�t����t.��JD?~��>o��0���{�[P~d�'ؘ�d�2ϱ'jQT&�e��x���l�8��.�@xxx�n�m�%�7��t��S�f����dK��3�(H`w�a��xxI�+�M�W���l��R[��P�G�=�c�����6H%�ٲ���2u�ѳ&�WC$��F��x_<;�w0�~o ���E�ִ�nG��6�n`��Q$�A8��l5QltI�ݡ��C�42�ʁ9���G �I0
xQ����Սb�c%�͋ͫ�/��G��$AS�䴂Ķ��.���g��v���Y7����Z�1�����|}������7�������Z������:��>{����[�{j���
���*Ё��A�߿s���:7L��k�\6�/�y1#�f�ӫִ����hV�	�WУ���V�M�Rh�:��*BkV�%� �4\A���֔�+�y�Z6�نѺ,.���f���r9�ZZ���.˴�p�,˭�ι�TM���7PB+��U�tڒ��3iv���V�2+e^oК��K��lj�khA҂��F��ցu)A0�mK���e�j�X�ʀ�7aci)��JM��e��ֱb\Д��B��|��x)�}1�2���罳%�#�� ��b޲��ĂA޼'�H5�GJ[���Ј��{��!b#�)DO����,H��K��]ِI5�ӄRgg�y�<���1�~�/br`D<<B2/ɖײ(�oϲ��/3�I�m�m�|�Ȝ�l�ƲrE�Gbz���RC��9x����<6>�l��@$Z�de���:n/��|z��G������� <<;���ع`��A[�D�)���׈��ڏml���?�0�,k��l���>ߟ�n�޽հ
Q�Y�o���y-%�#��Q��SP����+��Z�����Q{�C�Xi&Q
8p+�3$�,��D�E�t�z�+��f�^2�1W�H,	ތ2M���[�৪���gob�o�.W��c�b5�1Y�<��ڵt�d�y���LM!���v�=��w�%���zV���-����� �)*#���1��}�|m;������ڊ^��勲]}~&�����e�_2cZK-�ܺ8G?N3�,i���`��H�6��Z��[�ı ��� �X�����y����]�.4?���:��@��Ѧ���.��,���A�v%��s��$��D���$r�{�q��]�˴T�E�.ˆHtǌ��"�2|Ԋo2q��"|�.�=��q&���@X�
ъʂ����s��h��T�u��˘U�K*lҘ��߿�I��]�����
�{�AvJ��$IbF���{Y�}��AV��1��6�0<���&��k�ӿy��Ng�i�"H=��.<b�s�!]����q9VB�	���c���&�!K�h���꺸�U��O��ҝ�u��ψ��\jN9�ײ��x/�N�	���n��t]fT��w��m^X� �S|�1��_wtKR��H�m�B�;��B"*��]�a�tИ��� AL�\���0Z�k	]�2��'ۧ1s�b!<##1����"�h�y�s� ���Fw�2'Y��+	Y,���@$x䯻w��|���t\�D�3�&ڍ�:e�����jJ��f��-\�Z�&������9x�7��e�ˮr(�,��?r�]��{W��+�xXw��ڂ,H'��4�-�n�C����vS�! 7D��Ɲ#f���%2̼� �	f�$�iI��<�H���G�Ynhk�<:�gf:9T���B9���@�Jɥ��ħ4�;[��XԠ*��2��훃0XM X�>�9f�Yp��������i��Q�e�A�i�w6(��oI$W^@�H���6�� �2�O�������C�O�2���["H�$z<�(�	��i�x��.�NG��.��y'~����6��3�lٶU�������ק&���N�[̬�=��%rp[������܁�C���-$HR�Aϝi�D��@�ITQ6��B�5��X¿�|���ڟ��X���'�DXS���'>�D�.O��ZܕQS�@"Mǣ�� �w�%��zkN{����9��-�w�ڇ3e�7�f��m���-u�R�Ś�ݕZdԶ9WC�����넠DBxG���l�G�("e�7}� ؑ$�?�q������k�c�q��$	Ѥ�^.��zd�מ7��m��:J�"=d�Mn��<�R�eK��9޻a��?v�$Bx�i53���t�I��c��t�f��1�5�)��k��C`}#\PF��<y�2�����\���R�1,N�l�6�{�m�b�����{�2	����tC�QT"3��ݕ2���;��Q����%2d�w��N��ǟ9���`���78r��x{��X�h{vSFQ�d�:7���%2"j����Tr�p��2^���O~�^<z��Ox*sL Pp7��\�Hc�a�6�m����.n˂��y��8��O6��B��F����
�@v�{��]\g`st ��6:���m4c�^�@�J��j�%��/9&Q���L�3Vف�v#Ɇ����nŎ]Ve��֫sR�-���\J1-�Eu��l�[�Dv�˪n�V�`��-j�K���4R��*�A��ˀ4,��B�F��@���M�Z!B�\�rR��]J�:T�ڹ#�`�L6�J�X�R߽�ݿw�nŋ��!�}ޖD�s;�fĒ9��%��̂h���)�֥1�&[��2M��|p��O� c/fH3�{׃���x�ۇ�5�_lI!�w�fS�E�fG{���U����I�**�tze��`I˼�jLF���l�1-�[��q � ?��$�b���O�M�N� �D;������#Dvb�2����EE2��2I#_��g�m�ՏC%o	���#�F	���!�=Ϥ�m��@Q��^d�lF:KKg@�Y�m	ElG �u]M����=�s�Y�+Ht9����R��r͐n�3S3r��D���e6�J),QB�	�������4s+��_ϾM,���< ��O�M7�Y���u�Si��3�%y����Iܨ0���o҉�εgΤ����S���P��G��޴�>~�+7F���޴Vx��nR�U��x������d(5��i���r��o�&,X�
�L�'2��$�菌�ہ�j�~���|�u����vg=�$�އ�dX�=���;+aRPj��aK�"u�z^L�i�Iw$Õy���na1X}1Po3�Lm�p= ('�Q�I%���:Bž��F�>n���.D���lz�9:x������V=��ؐW�G\A���9���Y-ȩ�q�N�f<q�	bE�d��׻�����Q�T��ښ��@�Xe�@f[.�i�3&(�,�*K����h�;9Y�Y�={�� ���h%���K��H5��(� �wD�|_�t�ƏY�ܑ ���d���B�qE;�G�$䨮��g]1���&�MR	1m�qؒX5ot�$׮�g�8����p�-���]�$�(0�=�� �7��,I �#��Ե�"�L�O�n)�+&��gݷ��ȏe#r����pq�p�{yb�{���c����o�l97�fxVw^m{S{�ȆPc@e|�m��^���;a޲˹&ێ�7��T���yz��?�m���
�t�4�R��}3t�����3{b�{���] �쭋�T p���qԬ<�a��{p{Vq(���i��w/G�ɛ���S�����sW��,o�\��AT�#�G�f�_���܃�@+�|�x�;w�v��L����qՔ�^ݷ�9�_�Z4�O��ψ��a[�a��MN�ڟh:�E����!��D�O%�q`��4?y'��Y�=��p���w�2g��7!(��}�fRneɨ,ݵ}���g�7�ۏޓ��h��mgL8:����O����u��d˳�;�4f�|� ���s���O�Z������.F$:�9�g��Y�#k�oh�/��n�~��C	7�����r��;�WJ-��^�P�	�N�s���>�cE���y�7��ބ��&�8��v��l�	n��T����s�0�'β����^��x�xp����f��g��K�o'=������)�;�����=.Էj]���:׃�x�eV30/b�v/�VPa���i��;I�q��a�i��OH�+7��0+<Oz��}e`�x�m���f�d�P�a�Y;@�t��I���ؓ��=���1˘a�'�)EAEe��DX{c1DP�,�
Ki��2j{<~:���g]u�]u��ooo�j��CIQKl�$^HL�)MMVq�Aܜ��"|x������>>�뮺���^���͞
ǢR�2�A|�X��Śj5,UF�� ��dX�ǌ����������뮺뮾�|���sg�IIm��F1EX��3̦QX&�_&���(�"��]�ʙLX�,�ՖGUV �V�(�h"�e�X�+
��h��X����[e�QTET9s����5
""���mFiH���(VV*�ˌS�-PQUD[J�QE�U���R�+[�r���eQ��E��ED�X�V1l��"��"(���DB�QG
�ȉm�:�"�UdA4��'���2X�6K;������=v
Ċﾑ4+��9x���/׾U��_v���>�|M.X�[s�d��{|�x�gf��5��&c��M��~ �E�tzm�2vn̕ާ�3�����2�I���@�@"O^̉YgUt�F|$v�~b͹hi������*�Ů���!p�K.mjl��4����Xd�%�<B?g���u�<<;�U���ȏ!EgdH>b��|&�z՚������2ĂKz��#Y!M�x�:B	�
-��~i'eqm��~�'�CwFͲd�� ��H�A�9J�2JK۵Vx�=���=B!��<M�2	b/�bA,oj�A/��BVnvr��
d+sjA �{�fL�7J�$���� ������W��jY-��� �D�u�Z����by��^��M�L�d�*�<rp�gL&� w׷6-�o�z"<�y@_�oVF�X�4�{)�o���7�n�[<�Q?��K,��R�x���m�^��!��v}H��2�7A,z#}tk�`�����=�ќz��������ϟC����c`��h�~u��6˓��kr�M�I�H-�kX��4e8�9A�JK���8���ޏL�]���	,I8�D6ώV���>���dNz2d���DBxxw���<��(�Q]x=�0g�6zh[̗��Z�;$�~y2	���{�{��Ůݠ��k��s(�z�� �}~��2�&n'�C��d�%��Gă���(���3Z���xD'q

���L��;r@ ��0B���%���z��]>�x�5qR$�O�)j|E'���߱��An�D�y�b��JZ����c^��2����d{�1x�rx�v�dH���n}y��C�zI=6��|Ϲ���Ѭ/y)n��7罳�8���?B��ו~Z�ߢ�qQr�=��úH�N$���D����G�U+m6?_���,e�Ye�A��CB�E�����)��xh�JL�If�h�� S�,)5�������{B�.��t��HT:���v̀�� ��5V���8k��Q`&�tÍn���\`�6���8���;Q6C�l+�GmI�A�W������+��.TG$�q�*�u+�	�����x�����,,ѣGfdhL�Ek�bm�M��8Ë�͹��H����p��\ie،J���C9B������)��|��o"A��d0 ���+7Ϟ!���~�u��$�	���,H���Xt���k��-�H�Dy�z�Y{/���e��NOML��� ��:�U��寮	3�o(Q��${�����/��$����cn�TnH�I��ȓ���L`L�U�N	��t�DB&<%������sk�|/�i���6� �ݝ��`��v�%��Y���6.4�3�p��xN�!
$U��̒I�w��!�>��\�7��e@��]�$���ξ/7F^8j��D#^&�]�.B(8l�Δ���jG4v�݂ܘ�B{�|�[	$�B���^��4�q�v�H$]�D���[�H7g���Y� �H��bhP��� ���5@�o�H�[y�!N� x��s����` x��I7�}�Q�?+�RC=�����p�$��v���5���ao=ݻ&�`
�,�Ut�MP�?��f���)Q��`�0;���(d��7۳ �C�}"Ab�����3�]殢J^8NI���zZY�u�	 �ddo�c����."�v��̑n�I=y螲A�5���M���������^�7pO����k��A18�ht�	�sC�]P��eC�8���������`H����9���a��H,ke�T>���T�UO��=]	}~��} H$�� ��-S���Ͽ�K_UR�����fU#n�@��hl��df�yDqi1b]ͨ��}&n���C��.�+�i,I=�d2;ݞ=���� �e�L��m��zI8�w�co�Bd_�;b��J��$�َ21���]k�s�� nv����a%�����판Oz_H��X�;��W^X�)�;
|@*N��M<<n�y
}e��M�r#�<��w��ϩ]�ׄ�=G��S�����w�B�R���4�ɓ,Q �s������Ad�{럭��e�H7�A똗rL{��{}����>�̕2��PH5��Egt�����>�]�X�l8���'t�s�`:"DC�G�V�����o��=׷�|P�bo����$�eGbI�t�e:��zH�ėp��]b��WȌ���JZڮ"��it��	��)A28j݄���D�c�0�{O�$d1wL��{Wn��`/蹐X���#��3��@�O�{�@"4o�����O�KS$ٕ,D�P";�5@�9�u}�1�86�4qxB%8�w��;����{��D�S,�n�-���=�A����Av�q�ޞc�I:;ßb �so��v�4�=OU�[�K�J H�͙bO2��n��e_vDQ�F
�
1F���~����TY1��x_���ٛ9�w��3��!{O*����V�jN(�	3bx�O�;�t_-��t��Ǔ�K,���Pܳ�;���$�� �u�K�&/�b�I���P����Gzdęc��=�3 �H��d]eƬ�5��Q@�$��y��D�ĻZV*U�A���2�Z���ں�4*dl�f�\搚�z�.+�>|=������/߼~{�ߞKn�bX��!��#����y�AD��L�'=�"v�H����tDB&2���H:�@����G<�@����H�#z.)� pMr�����:H��Kxr!�"�w�e�G��I�j��	�W�L��Gwl�PE���[�pa�ՠ�)�;���U�U�n3]Z�A,z�����f��bA#��nJ7�>9��D��ɖ&�3�X��x�#�;2$����O��}��\Z޺e�i��˱D�}�2^d�5�bqܕ\�6$ߟo��w�>[���8ڳ��;���W�{�+ߴb��L��\���ru߿o{�b�w�Yw�$�Y.5���ڑ o�V���]W�ڧ?���^�q���}B��N�;L��.�5�k)�H@f�BjfT���T���/i���JgE΁dD��[��I�B�9`ܶ�h��f���H.6$��L���ۊ�]�;p�2�2�-��V�%MaIF��3�T6�.�E�m�r��cF�6y���5���/l�g��)n��Ƒ�i���� pK^�ʵJ���f�\�T,F٘G���6Q�շf����>��C�� ��&$w��>�%�5y�ƤAe�KJ�[�lhURQ�7"I=~���:��bi��)���}�k[�>#�_��k���Q���}o�I$�g�q��4 �C!�s)���j�\�՗<�l�	c�-k��1�@}pg9����E���z�?�c��Z��Ls�&q�W������8�����q�חG� n�b��#�1�X�H�ޝ��#1�q�;"��X�Hw��)8����~�A$��d\��������UIa�Q�K��H��#���������+�M-�3���ޣ�sA�h�J.R�4�C��\��1k��A����$�K}/��̽�4a��-Lnׂs���/&<e2�$��h�-&
.䘑xݓ�$��h�W	G}�g�16"�Rm:�;2�VWT�I�ay��>i�>ד�f.�|�R/w��d+������1��w��{�y�X�����?K���O������AX u���m������\&�����|j
]�k�g$��_��z��N����""1B�t�x@���id���ɀ�Ț�ؐA;նn��a�K[y�ĵ��>�I�&���.` �`zg�-&��ZN��ۍ�S��AML��솞eʲg�j'd�����]MFxC)���f�f�#(�%j�e���&��r-a�A��ф��J;�u����ݯ� H�cP����<��5��<e�ٯ ���P8��:w5l_k2q����P��{�Ot�2�{�y��"�_���Ax`� "�tEQ��(��]�s�(;�c��蹒X�z�儂oڼ����
6\��?�{���	�ɾ�ͺR�jŅ�����*燐��G��;&��ι��vwW�aRs���de�e���=�a��7�2�_{}�$��u�(�O^#ŏM�Q�${���WT�WGP#f��A"��$�	ݘ�+��KzI՜�4;�7��9�rb[�/$�@5��!cFד��I4D����������ޑ2�wS�"{�32wvɴ�I�=h��~�<�e*@���h�L8]�����5��-Cub�"�<wL�L�%���Y�c�1��_.)�Cf:D�[���ϛ�M�FN!(�1��(�D_���Q����I��Iw�)���F��-ۮ���]S�u���4�I%�0-��0����G�	 �e�n=H���TA͝:�}�s�礒36�A$ltq�M8$��:�8��ܓ��{�%�dױ���!��q���Q���j�<�$.���bz&lm��7�~�� �v����.yo���t�g�Og����𞏜�}^�@�����̇��Ѳ/v�7K�IH I'��K,�,�E�_=����_s�/�Q� �G����H�A�����ՒîvdEG���$�_t���t��-}��~$X[m)��� gXK��(�ᤣ��z:X�àJ�A��ȶ9Y��>}���7-��SD�H&��d"K�ޙ:�vm�9���总3�8���g�QUh�V
��D0x�o`��<�=����?C�Vzw�I��F�w�3' ��Q�#�v}|���݀RIe7{��$�BQ#t�}0��=۰$����<���fh��	 �)kɒ$2��X��@��D90^ ����:[�abAM��!d�g��X�v߬J�'�y�c�<����I�ZԖ;C�D���u�� ��Y3��>����u�&q�� ���t$�_C��T�!t��1�-W8���5�P�l:��D��_d������qwu0b�D�0���}Y\������L���Ԣ��i��}�.��>����}������y�_y�`�9����M����wl�/N�0=�P�ϑ��B��ʋ;o�eL�^� ��)��Ol$�9;_��i�=��?	�;��=_�#��;}�p�_9�X�
e�rn)��_yw5�2/v�ǯlO��8��D��G������rl����t~/�������ӨŶ���n����<���Ѻ�a�'��xh�ri��zZ��g]:��V|E��x���sۡ_]�v�#��^8t/�dj�܀[�6C�}��b|���|���F�a�M3���{x��_�5�n>��2�Yb�~���n^�����X �+���0y<���>Zrrµf��x?z�Y���-�X���=����6����+|��,w1�뼋��>7� ϳo��W
1{��EV����{��k�h��r��/B���h���g�s���~��~��߽��خ@��Bvj\D׾��6��{��-�sSx�u�g44c�Ri��gzի�Լ�vo�d�����+6=����4��Oq��Vb�9}�cQ�0y,������픍�a���'w]S��[���Hc�U�wm��w�}��Y�on�o�q���hw�&H��l.o�r�	~���Z�i��Y������X�s���Ԃ��td	CÈ�m��2���=��!Ak~x�z��hC��}�����X�x~�س��3#��ct0�0����(Ki�f�)�)��J� |�>�\� <C���׏�� }W�vՂZ�cv�΅�>��ԕe�kQ�y��OAsHK=:K3������H�ڰբi�9�q<���ޟ#o�a[���n�`�33ee�G�m�՞|q�riu)j޳2�[�ޟ��*�堪��iAZ�&"����Dt�
��Ȧ�9��fx��}?G��~�����뮺�u׷��ё����$�.���j�yJ��V� eSO%�D_c,�S��������|u�]u�_�����謺�MN5D1˧Qm�[miJ�)ET�
�=���N�糩����|u�]u�_�����k�8��UVѤ���TVEbڡ�h�"H*(�,�Y"�s�*"�X�:��"+,Ͱ򪘂&�*J�.����
����U�/0��
�X(�t��3ZYYcZbStJX
*��pUDQR�mY���kmU�0U#*�(0E^䖊*�t�(ؠ�	iDQ"J�����"�mX�혘DUUT���a�����"�(��P+U����*�*0UA1P���Z��%�(�����j��*�������TQ�Rڢe%�����M�V��;k�X��b�3*������%�!G����ф�)��E�M��v��k��bя4I�F�\���ն��DTVQ�.��cQ���Pm�B�l7An$�V��Uˁ:�����ܛP/yB��1���iY�m5�TNfծn�ư�3�h�]b,2�1z�A�QSB��
�X��G͠hkbJ�#]̵����W�U �ڔ1���鮩k���[Rg�3t�k
���Zke�m��*�m!� -f,e�iv�cVF,�%L�պl�5�lŀ�pfض%��-W21�5rR���ڦQЭCl�t˙n��FkŲ��s]rVi��"Z9�*	
���.9T9��k3l���l,H���R�B�W&��44$�鄕AvHƤ��SM�E�fhCAf&[��pVk���j\^�]1�aY�ҒŹ���M*5���Ķ��
Ұ�Bղ�՘��(�"�h�y�Ŏe�Љl��7X��X5R^n�L�d1��օΌȡc��XK�-LXK�tr%kױ��ˤ9�i`��S�ft�/@ԺT%2�K�ŕbڑ4av*L]��ܰ��c��E�aQ�H�gP�c���l�0Ս�H�	tF��ݝpB)MKT��&�i�g<M�1	e���d�����B�У���ֽm �R�n��v
FZ�����ff���їdqD��M��l2�D�.�&bg3X��7L��5���p�m��f,3	\�ְSF�֖듶�ٵ�F�r[�$�(8�	-/b�6튰��Y��`��`9c�X����u��"�qm�t�5�����Yj�4t�F��6-��8���#�@��F�ku��cC\�$K/g�Dw(Ki�I������(ַ*��Էmkfb�mK�4[����q�w} O�Z��ci�J8Y�k�e�ߣά8�3LFU�`��V�R��]H�,��]r��`v�\f�+���M�3R6�S�:�M�f�JT��fl�;tH�\��[f4×2jjSl���r��҆�Cc �j7K5��&�J+tôe �e�DIBZ��{<���Z������i����Z��2�Z���Ұ�q�5q)�j7kY��f�3�r�ͭ������(�b"G~�p&��Ή�A;��,e���
�_��4ΞRF�@�{&A"�AIqO��'rc��t\d�� ���s�O��X�#דMH�,{o�F1�[��~�h���D�t4���v��[�LI o\�M 9�{��ɸیä�^g��$k�q�����`��y"�x�W!ږ�X1�Q �A�mćd��~8�g���"z����]d�5x,ǈ�&D)lc�$I�Hn�	�zb�b*��ڂ��@�Xm��H����9�x!�.�#ϿI���mxQa��P�D!�� �L��f���n�.��`�`�9���5�g.H�I�bt�;C�D��͹�<��ne�L�$o��z�X_�U� ��2	bM�\�hom�u���a�ݬ.�Z@U����!�˝��%�u�Q��0g��.O����5�֏dlt*k��}e�1gy��o�rُs��A�.{��{G\��oOU�L����/y�}}Z��2 v}�%� ����L��P8l�d�Ӳ���	���LP�rg��KkW@X���� �r��eĜ̹a2�K����	lX�Z��D0x�G\,��\G��<z�!��L��]�1-5�FL(�o[v#�ؚD�-�}Q�1�H���}�^���D7���L�&��`�';�C*Ϳr���}������U�Ю���a��� �cmf�Te�i��*B�^�p�w�" �����}H=kІ&DS�H��5��ǃ�y�ށ!������,v��1-w��%2�e��2֣b�y�$׃�'7���f_[�����=v@P��<H���5cٖ%�_t0�%�,���H���ެ��M�O��j�e��/��{�KȀc�,�=Kj�g�a�,S����((�������D~��
��7���?:����)�}3-,��$�v���t�X�y5��
�l��֞Ra�5ݓ'�"v�m��ڜ")����򁁕
)Ӎ�QT.k�T	$Wt�����sEKz�ڲ�ۑ�	�ޑ=R��ې�Q��#e%
s�3���`���ɵf!2�у��]KZ��J������/"�;k��$
�ȐH�e��L�O������|�T�����^4[�xt�"Ex��L�&]��U���O~M��,$�Zs�2H6�߽�	��/C�|9�Bv|��{�%����2�N1���K$|�^;�jK��פ0��� ���9�2}3;`��԰q/��x��+չ5�YO���U�@i��o62��r�sd+Ԕ���s�S���YK&�g�\N���=�W^~������;#Z��4�����ڥ�Wg3�;ni�(}�Q�?��1�c*C����wξ��,��E>7��N4%](��?tךj!̴�K=��}�ȫ�e�kh~�M��OL�	��X9M��?�Lq0@�g��8PX
Dݙa���َՌ��I��mKŘv��)a}~��-B ��K�y�u�so/dI$y��ܠ�m�Y{茩�ٖ-޿H��	=ߓ�4��h���޻:y�������K�yu>
_�5���#w��${�5~�w���t��DU���o�9:�����R�i��2e�쩐YѼ�+͌��S��q$�f8K�(.1͘�7�8rZ����i�/����U{V	��m?���ނO{�����B	>��q� kǫ����������/�A<�DKV�D���TA�f��P;_H��ӧ�o�?�W0�zq���^Q<x�JEG�)�o��[;�_^��V�� uk/L JH��cx�,��ˏc1�XT�����D�MV\�l��ǜލݿ��,c-��-�K�.����iiz,�U���4��:8m!v�Ç��7��a��E�&�6hm�sV�hl�t3w0�t�X���؃���0�N��6�Ia3��a��3ե]+��#�c&и�I���Zꃔ�kB��;D�͌��@��Z����ĥJ���x�%�%e�ifMX��*$.�%���%�]�B�!6KZ�M��LV�lvBje�Ũ{�|>�O�Ƶ�?��TKsW�1�K_GL���4fF��}m'�2D�	j��!��)y��/o�E�g^����c�S3m׽	���u׈�	i��u��p�$��~E@ ؓ�׈"<$_ٌ���,F�lI$l?��;:a���9D�ٌ��>��-�Q$��	��#FX�u҅�#�=��G�B��D�Y��@�=�q��V��=��c�����Q��2��M�"I �^Hi�N�TL�q�=��$�m�}0���s}�>t��PIG���.Ź��۱�ъ6���95�l�f� ����W�z����Z�Zl����<��A��$s$�˕�H7}�Y�2�ah�� �d�gt�$[�<W��˥(�T��@���t=��=�S1d��<d<U��!�ș��t�.Ob\��� ��{�{bg�`Vy�8!&o�J�'�9��l:X����5�,d�6d�h���L�u����4��`����~yq��I5�s�`�%���>j@��s��b@2�	$yЭ�d�w~�c�	!ܿ{&I$��E5�@��/Tc��Q(J�:�!��}p	�riD쾄�N�@���y1��w;M���q�6I ��(�P�#�=�H�y���ow�F��w4Ƙ�y�ked��W�x�u<��LC�6���-u�4fB�6��˝&6Aڵ�DsDqe��n�u���ר�5ד<�F�CLu�	f����H$z�2}=\�<#��P=4�Kg�^���$��y	�K{�@6�z�ѷ�w��g��I7���h�[ �K���m����8$�z:$ �l���O8�t���7p��Qs�|��?
�{�3R�߸�y��_'9+��w��y���F���״`yk x��,X�b�"nG�̂ �{�O��1s�W����/*�k�vFE�{�k�}�R�A&��@0ƻz+���z���ޏL�l��D�/vc9�o{"I]���T�k�,�S2ă~��o��X�_�J�#�̼��p]=E���@6F��0He�.[3�����.��:Z��׻�r���x�n`^�8r��1U��'#�	���M��Do���̂z���	IG����0�c<����OO���&��,�#/�A�Ay�KΉ���fܹG���\W���~���s͕�Բ:�d�.n��<"��ċ��$j��I"��k���\\ܶ�㝮 x2@�˻"I��ǝ@wP亊_��\��� ��10���	��v�A�;;�{��%�`�#���w}|�����l��;4�4��f�Ŀ�Q2��!�f
z|[��=#LmIsnS���g%�3
�K���e�[�\���͟�Ct����x	"�@z'�dX����.6�z�H%�*��.��}"sr���٦e�4�c�2��4rD�L�5�謱\k�L:6iD�SmT���F$?'�x"���xe<A�A-�D�d� ��t��G<C�ob���C1@m��2�Յ�:x!�*�El�cO��u�U�l���	N����CJ.�w��'���]�g_	V.��|��M澟8|.`�%���z�i�<��-56}��깇�g�z8�W��҉�H�j������}��Ĳ���K�n����پ�Af}`�d)��wH�����8�P�9.���>��,H5�1U7�n^3�j�{d��kT���3Ӳ��6�۳���&H� S�z��z��"���&�Oc��aA@�V��w�yH
�����ϳ��7"9{֭Ľ	�G�O^�!�^�3�у?��2B��jm��vQ��b���J���8�0c�5GFm�W�z�8������p���48�Yq�U����+��!+�{%ursY�ZT�۝��f�:.R�.�h�4фJ�cF��n�ɣ�뀷0���5�,Ԥ�P���n����l�kQCU�������2fWMY�!��m��JV���+(�jQ���&�0��I.
�Q�	rH��#a�H�ҬkT�j��Q��Ƅ.��5`P�M��SQi�6uu�0LV7MP�?��}��33Jg���52	bA����ށi�9�����EIc���L�uG�C����t�w����.�8�H�H{�2$�q����uG��41��;�>��"����f�fu���I'+�y�QBI`j��A'��@��Z��DC�)��c:}0�3�x�Z.�2�Ζi7�����:3ڹ�8f�$�gKId�o�8�*"	���K{�y���u�"szbM���^�Ot`7]S �H�z@.Ƴz(%��^����~��ҍ< Θ&�HP5Z��9��u�B��B���.��]�Bg�߲~ ��/�>zxb6�� u�"-�f|���u�1l�O�_= _p/Ō�}���?f+3JfG�5�2I�����~��!f:D���w����u���9g�s��5>�5S��L��` ��~Y����\Oܽ�?:u��3W\�ٸ�$�Y�5ֿ=����&v+����%S��l\���|H�Ҭ��<�f;�	bX��"IĒ�bI5�N���sފ���@�VwL�Kt�A�n/�	���1u����C�o���Y�q�J ��D��=��v|"����v%��	A���>�
�����vϨQ�ٓZ%V�@���	5��$�X��E3�V�d�k2B$��?iB�|�M]J쀳k���cd�h�����kD�)��Ş��=�u�\���;�?`q�n��Y�%43�3o�Y���fq�ף{M}� �$�ޙ�l��T9F�Qb��mąl�%�j�d{Os��}}�$�}��2�w�X0��t�t��Bj��#�}���Z=x���K�*�t:v��RXj����V�VB�1������]6-R�D2��9}��~��G@��ix�R��cs�S���q�$��zzo�}pb/7�k��3��;m�z�퉱���o��,=��_��K�^�{�>�r��t�����o\��[V�t]3�JT�#�Bz�H���Ǜ�ڤ�f�ۥ��vc�!��e�_��3��e��/�=s�-�I�A^��̶HL��g�1,�	�k��*{��o��������/xk\���%�{�=�/1�ףd<�!���͙Zͅ��,��~n_]^�< X��O���OW�J��[;o�O�����g�Ǟ�-�X��ĕ�M�g#������i��v뻝�٣(�i,�3.=������?0���7����a�.[
��Eβ�N��8'��%¶N�����=C�>�<7�!�!�>~v�t��'G��pӝ��tmΚroB.r�����o�Hcww�ҍ��̓�c]�k�S��,�9��x���v2W���-�϶��Z���"������b�/jׇ�c����Y^��1��M�=���5�nv%|B7��{F�IW9o;�▏M�%<��{�.�F.w%-����v�	:�|��gK��R8�nͫ{�Or�<_�D�̨w��sN��	���!�>y����ݛ��W�w���ox��ɇ���hG�K�u2b4 	"�j�-U���R�UX���d��������9��&�3��|u�������]u�]~:���謁�&�
*���TF�û*)<j"�Ŋ�1UM:L}��S'O�������||u�]u��oon��gy�
��U�$�5PQuKb���RD�e���;�2*1&5
�{,������v����>>:뮺��׷�^��
�Y^�ezq��%A:f"�#**���)(�b����%Tuj��F
T���TX�{��]Yf0�Y
�&в(��Q{�L��E"1�*1|ID
�&Z(�N	�����`��
*"�(2�M$Iwr ��b����"(���*���4�QQ��b+��
���EQJSG#�2PM�*+J��V*��ʂ�Fq��ʊ�m(�
Df��X�fZ�*��DX*�PG)QFJ�h�g&�������"�E"��b�x�PVvՌM�
E�z��'�:�'�׳�M(�}D�xt�x��=َ��Ǎ�Fz;�n�%��b�T2G:�$GwCP���^F`���r|�	'�LDEQ}��jD�<;4�}�� ��푭A$��ɖ;}�x{�m�D� �hYH�mw$�%Ԍ�M�A�7l�6�^������C��v�q��]��n�ٙ�Z6� Ud�� :�:��/!��S-"���4�N�:<A0�vz����DZ��e��H1]�����",�wt������`#b�[.�٤��4�!'Ò�,Y�ː$��*�xL�,f��k<���lQ��ȐA-��b�݈xQ�
"Eت�WTj'�˙�U2A ��id/��p{=��T�Ji+gz��=g�e��w2K�O���Ü��ʹ�����3J���.`�BxŦ�|n�g��n1�c!���[���������� ���]�>|��2��D��>/z�(W�/�ڙb��[�2_��nYz{}���Iĥ:��JP" T�(<깖ݺ��Ca^V�4��X޷r�8~{�|��m�"x�D�I������B�jY&0��c��@'3�<f���@r�USlw�Z�>�)GN���CKJ�}\�f�ݻ�LT�Әz�(I�	���r��H1;}4Z��+����&�{�71�]�2����8F�Q"�F_����⾔�2l��:�Q+��4�V���~���1���M�#٫ėQ�
#ޞ��$��闷��W�$�W@�X�7��,Km��3��6�h��u����	�y_~;�C�(Voݷ�t�������fp�
�{���zvy:�[�pg	xS�ȉ-X��߁����D�{�|,I{V�͊���Mh8�k�&�c�en����8�N8�Ǐ�f��@f�.]���6u�d�LRl3�N�j������ݎ��c4s[c��V�Uq��HԮ�6��9�[���0WL̀+�u�mrf���Z9�Q���Z�Y�-��D�e��a�	���lL�P2���u�@�v��]SB�N(N׵�cT�:�\�]�3Y�BeM��+m�Y��,t��M��o�qNI�ܒ��͊�G":���������|�h�ɷ������z�]��r%��!�}2O��}&����'gD]�L�!����E'�1�l_�e��}�>o-w�."��l<�i��*�"��Ao_�H#w���%yR�&x`$UΠ�A�]���~��Hu�L�I�3���z��o��I,{��4W����(J"���eͭ�"��~���G_�sCǢ���b|�s!2����n�{�h빒p7f�Cp�9.��^v0;s;��<����!z$�v&����S$M��ZA	����4�(�	�<�5Q��L�"<���l�UhJD��4zݓ3a�5�Z3F�@P��ن������ �v�U���ׯs,K1�o�]��z����Mx���֤@$ع�kHZ��'��Vzy���I��}����\��H6���`xT,�{��FȾ����B�z����fE}�h������?��F����8���7?�,c!����Y��N��$��H4:'����S�̀[���ӧ)<1����~˖�a���$��[�:�P{ٝg�S�޹%��%��H&��C!�@r�_+�{��������J[�		'��Z(���X�I�	�n��X�^j��a&�׸w �(J"�����~ؒ��{���%�V\���q �w}�=]^{����%�~�4KJk2�V�"�Q�b�Z�A�v����9v1j���~޷f��z}��e���Ss����]���ɓclY�r{,���닁 �7�)���]�8I�xNQ�M�[�&�4��bzH�>�Bd�'{� b���CS/+ۨy�ǉ���$h�K:p���	��'8y{m��W;���S������cԼ��۹p[7���ܚG_�Z�����p��o�}��ʇs�-Ԝ���ywygO<a��y�������n��O_}2	�_�D(�ADCȻc}e?����Y���ǂX�q�ە�au����zzBY��Ǜ�0!��y�ІC�����n3�d��@��frO9��O%���ݡ�7~�H$���A97��9qP0v<K�����>�6\j��lن�l���N�e�m��+��fPІf�/

���㇪\p6�+�lKlU�t�vK=�Dn0���d��d�<�{��b�#è���X�7שk�u#|��	$�W��$':�yBų��1�xǫ�^��6ϵ��B$�{"H$�WN\K�������}��Pޞ�2޾"��<:p���x�y��5ϧ���I:޼�{������$��}�.xޝ�z.쪇K%x�+�9��T���uۧ:�N�#�2��^�G�u�ikx��Z�;w̙p����Sq~�X�bňa���L�"��$U�:�P�����/��jA��>O��%j�=9�-�����ȱެ��A<�2��Y�QGt&�İ$-��I��`C]��hisCuŕ�]*�K��ٛm�3�翗�)V9w:��&#�5ђ$�Fw>1�4սء�Y�re��}��KSzo��(1���]<37m;����-{���d�9�I#��;;�U.�c��z���»�P���QB��P6�^��$s̽,�=��' ǻ�I �z2OޓD���p�<U���/��+D�$S�"��8�X����_�zG_9��X�fL���6W(��<z���=��ro��T�/��,-�2ݙH-��!������1hs����&�L��J� �+~!oo+��a����]��]�TK�f�{��g�ï?j�?~�?�RC&A�϶J1�3kJ���$�	� �"@�
q� ��g {�[\�]�ѐc���o}�eD��79�������Ԛ�ͪ;g+�j�Qu�B�-H�i�v]��*˦���DcY�ؕ*2�[�-�3�l�a,4���(m�	���H��cV�Tі��i�M�\ᶙM�YZK
Qr���VmFn�5p�d@��m���ު�(�k�9���v��%����&Ƃ�R��T�m��	e	S:h�\�hbmu�
�M�*k�lȚ1Ո�]lC��������!�K�|���zD�%�#~yi@�s;�>��ma��L�H��������q��]��j��32%Uˆ=�[����}��H�醐�%Ov���͍�f_���IbA����" ;�{Ǯ� J��F�P�1ɯOo�dZ�>~�l��a�-p�zch"�H9��Ct!IG����lZ}ܨ(���BzDM��{����$�FN-����t]��[������������21�@���e�7"=b;��H�|0Ē=��&���qiiw�5���<1��z��=8ܱ2ǶȗL�H��`E�[c�t.ͱ�mX!˘w{FK�Bp�	߃�_�dI�s��^dG���96�Q�Z�`�����$��rĐ0�����Q}�$L�{s2�t�q�+�L�Ն��^���O�;�)F�.�;ߊ��������o�F�֑�߼/�_�^�ܨ�ߒ���+~��1���W�˹J�;�^l�'g�D�(��@~u��09������%��=��2"D2ȼ�"Y#9�6��5o�s� I�fă�v��>��;~��" ;�H� �+ȷU�m��n�x"��N60grX�Q�$;��UH�NFDx�Zۯ����A�� �w����۩�H9k�'z�\�*�I�;�$���jaI��q��`�n����>7���U����L[j�L�4�!7n"M*Y�3�� уl&��b���'����G?��|��$���HH�~0
�c��u��L���L��"R�N�'�=+����3���"����X�$K%��L�q��0E{�}t� ����6ս��a�V^od	-�H吇2�^ߺ��G��ܤy�=8�|=�y>�Oi�|2����{O�"�_���lE�>���E ^�^�=���.�݌������1�H��FK>1}�^��"P����vķ7��ƸP������|��8�ڜ�{�I ���I(׈��{P��`�5"H��$
�ot� ;�f� ��fD��S��QZd��{=��H��s ����mif�59��"�w--��>�J�"�b����s�,����%���B�p�e���t�v�l]�Bt��մ�2A �w�Mi`�g�0�t�|��7I�̐$$����`�D;���ޏ��eu�l�\硼;L%�Ρ�wyuQ �9`���
��c�v�ĺ�xt�D����H�l	�Ӌv5V��}�>�\(�W�y����A3y�:(�xA�B���g�X��f9ۛ4�\�@ry���ܖ�k��o[W���dO5>K��qP�����<�W�BL���D����1B�f����ճ�cݟ=�� �h�"��x.��,���q?]�?N�� �O�ޮ�����O?a��S�N�z�dH��&J~�^ѯF����Pău�%�2Gz�D�Qq��r	��i�
E�轇ik���-���`ɮGi���l�A�����-G,�>O�O���;Hq{�y�%݉}��9��/�<��C �]��>�Ξw	E�;�߻3=��.��#�6D�H;��'Y)��W�?��er��I��l'��p�*��l�$z�=j�|�a�_:��d�d+k�I �Hۢ-/C�w1_�x�y�f�סNvw����nz$a�Mw"N��*��'M�u��w�PD����95�Қ���(��Hƚx����F���i������,�H�`�����������  ��?� ����$���TUP�C�����{�H!�!
BBi��@e	�Ve`U� 	�f�f��Ef@�`U�Re�)��&Y��@��D	�� �i�@�&DBY���a�� �� �` !��V�Vhd !�Y�d��VBTYBBT�d		B��$$		BVhd	BB�e	B��$!		Y��$%	BB@�ed$	BB@��$$	BB��$%e�	�$	BB@����$%d$	BB�ad!		B@����$!		YBB@�a	BB@��$$		B��$%d$	F��$$	BB@��$!	B�`�	�#�$
@`0@`@���!!+!H@��L��!"�B�B��*�!"�B�B��a�����pHBP��!Q!	HB R�D�$Q!�a!	L�0AHBR�D�%!	HBT�P�! hl�P���q�
�
���%��"��
����40��@ȫC�
��b*�CC�4��40*�*��ȫ42
�B�3��*�Y	Ef!�VaU��VB BBAY�i�V& 3 ra$!U�!� �i� �� �� �� �Y� ��VfQ^pC�M��2*!(!0 ��� �����/q������� ����@�3'���������@~�����O��̿�Ƈ�����������0I���?__O�|�����(��?@�?���G�@�ԕQ_������ dG蟲_�O���~�?���+�������7�bAϠ|�������N�����m¿�_{�*1*�*�
�����
�2���*���
ʒ���+ʋ
��
,���$"�2
̊�������+!*,�+ ���Т�H+"�*$@Bд�Ј�% J�$B�	H"P��B�H�@�� �B(D��J�L"H+�Ă�"����� ��+0���
� ���2�� ����"�"� �B+0�� ����+
,$"�2
�ȫ$������+!�	������� ����$"����*�B+! �)��W�J�H+(��?XE�������'��TJ�J�����g�~����AA����t����� 
��?w��~����Q��GI��#���=k�UQEt>�?�?/��}�ܠ
��TQ_އ�C�����tb�����sBEt?��C���d�e�!�P�����٠�:�UV����P�_v}ʪ(����s�|���w����~'�w�����$����� �����?�UQE~�:���='�~i���|OӁ����]��w�I��zUQE}'�jO���N ~�������?D��郁�}{=" �����_O��È~)���e5��+d�B�� ?�s2}p!��� :� P /�@�d�� *� � (�
(Z� �[ � �M#F�@

h��� n�T�H�TT^�B%ET�PB@�I���*�*����T�(���P�J�(TU(JT������
�w�                 �                  |          ��r����]�j�J9��V������ �6���*�k����n�������-� ]vմ��R�+w:�1T�)�   ���:U��ꫩ[�uS�s��� =� ; ����� �5����c�� �t� Ӟ`�� �;�!!UQ|   {�        �@ 2�c���S޳�^`Oy��g���< x gK�
 ��� �` <�{�*� �U{e֧#[e���(*�   �p��R����*���� u/[ks��޳�z��i��s�ڒ6\�ʚ�8t3��nmp���ܵ.׻�kɋ�f�n��Vh)U"�T�|  �        z\�W�;v���)�ԧ���݀ի�q�p ;@���]���i�e�6V�u.��ˋ��ˀ�]���n���9�鴊D%*�#� {�W�;���sjUv�n �-[W.�u�k���V˖�\�ۙԧV-� ��km�ے1�r5�[+s��Rf�Y�k�P�"��|  ;�    �  �U�����Zjf.wt��ӛ���� wW2��n�Z�.��[k���ښ�j��ۀp�ڛ��嵆�LJU*�U�|   ��ϛ�Ud��7[R�n g*��evl�9j�i��7]5h���ٵn �ڶ�u�m��ݫe�\λ[rh�UQEJ��           {��ۺ�w:�Yk�U8��՚�]�pP���st���6t�����^�� ��S[�N6m�����5IU�  /u{��u��Ϊ�� �(�v�+Z��풡�Ϋ�ks���j� wWU�\ִ7[���s��T�nv)ֽ�T5O�JR�  E?#)T�1�?L���Q@� �?h����   ��%H�C@ �	
1LR����a�_��������O�$�7Y��1��?�Jg�ɿ���%�Y�B���HJ���֭��ն�m�:�֭�ְ		������Z����U�ʫ��U����3o*��K�Ӛ�:Ss2����*�/1�����ȶ��8�Xz�u��m���l�u���rDSЬ=ll5Evl#%ٱ�{�5^ܼ�f^fQ	�I_ץ���jV#2-�xT�KoG�L�,�F⽸,��7D�yFY�Ԫ�4]Z����5͡�@`ec7v�Vuk�O�(`���J,��wiaXR7v�@�%\j�EL���4���MHh�n&�`�%2I��9�4cԮ�!8vJIɮ-gX��eЗP<�m3�ͳv�1h�Fh8���Kב����՗(���jA��
m�5;���ñ\֮:�NMYu�)�#�6���ٕ&#w���ݹG*��)K`��Sr���{2ۺN�(���le��?�w�^�ܺ;"���C��7��Z�&�7S��\���v��T�(�*Q1�:������Yi�q�5�7��!v���Pi^=�&9[B���"�˓t�5���Xi� Z�:��l���ͺ/+*�:�,�AYv���+u�ԃ�����ln	2',[�!����x�K���r�K��Y��j2���V�ŷ��]U�e�����!��>��e�NYy!64�l�5XHM���r�9a�.��j�ɚ�Nf%/7r�fԽ��X�m��R��	��*6���b�E+��Vixf��a<2;��̏L�{�Ԛt��Z�w��+5���d��G�f���C<��e^M)��F�d1��Ce,�H�^2�V�N��˒�0�-����Cǡ��8+1�����V�Zi�~{j;�1TF�f�4��y2�D��A��f:y���2�$DҖ���D�����nX蛳�+ۨ��k_׸l����X)v�#i4t1u�[�Vt��-̠�GW�2(RTTX�������ʣxTo!ǋc{�˼ŋ@��z5a۵1���g춭d6� u�t@[��hce�����ڦͪ�D�cvY?\�Sy��y#r� �Mޔ�����Ou�)fᰤV���� � 7J7M]��G
���n���Ǜ$!R���[�r�������{Yw�4X�Ɠ�=�-�Z^�l1w�@v�'u���-�l7W��J�N,3Q�p%j��M^=�
[�W���(�FeV�w0��z3,�7	/u��e�)�W,@`*��A�^��{���{�E;?� �CI�8ԃb,�d�p^m@�Rܣ��{9�.j�u9�qU��nn7�ӷ�nV�̢6�4��J�mfN��h�C
X0Qv�ݷ�P�R�+�,$�� ���7X��๐e<ƕY��e�ڻ�dv�����Lͬ1��P��ͻ��1<��X�=ݳD+dV��(���)��E"�!Zh"�p8�Rwn�Ch �a�A���"�� ]�EX�[3mVE�.Ч�v���=�M��j�c�E��M-t�����c�ӷN>d�iI��ͩ9-��/xU�7��C\X���m;T{��l����l5+^�0kko`��S/)�����[]m.�	��V��W�3,��KZ���m�8�i�i����TRy7�#1�oE�f}���I��MM`��P<;Tk��7��������;�7EC�e�0̺��N�ƍ�Bп�ԡY��W��3i�;8u���'(R���j��Ym��& [VoY+�1��L��*��6��sb�5�����4(m�m�AXV�sU�;Z4Z�n戋������D����wOn�Ɋ\d�ªJx��$�m�4���i�5c��v�ӑ|���q��ߚ7�rʾ��^����ӳo	��i)7�d�n�-b����Mh�g"y���eLßsnn=�3WO[[�>.D��g3�rcn�� w4�D� �c�eei-ǶH�5�'�k8��+�8~�5d3Z#Y��W�ʫܭn�R��t�|��c��ky� 4sy�������\t�FJZ!�$l����x^;����A��[���+S$4vh0��Q�n�vY�Qo/���p%�'X�q���S�巴pv�}�:|u�}�C���he�CLA��n%[o��9��l`,�6m�T��1R�4V���*Yۚ3v[r�� Ԥoj!��B�{L:X��L������l����#LQ��O�l�
d5sMљ��6Z�i�v��e�5�Ớv�)��S2�n��j-嶭d�cݎI�w�f<92,ś4@��r
�s��̶��x�.�7JFާ���-%{D�`;#vdzj�rf4�{�ee�fnT�����
B
=�s_�xgƒyV�/D���m��*�AX�Nᥛ�������$����AO��n`�p�!T�TK��o��q�{�Qi/c���3oF�(L�a��}���cY�E2�۪��1��Ȭ��,4���Rk�[�m�۠��TP��uh�V�U�<4��Mw6��bKZ���m��{X���jV��N�Fs�1�N�%8a��ά�0'h2�^���A��$-nðUrN���3o/md��\sSى��B�`W��T��w��X��"+8>��a3�.�t�<M�n;�#�n,���R5�vY�N��ܶ��/5�YE<ش�{iI�;����|���Wjhi�h���wme4���`di:4��z�Ɣ��DЬ/wYz7/�`hx76���|�,�seN
YN�#�g5B�9��<֥��%�����"�S��ց�1�D4K���M"�[�mX���L���3cZ�2�d�[R��%8�l��`X�Ne�q@���5Q��R۲Ū��6�Uu&�Ў�JU�k4e��m1|������I��2�F�[ő����ǧm�9��X�U�q��f�Ӛ޵o��[�m�Z��D��Mԧd)�F�p��q�1{�.jVh�nVVI�S0��n��`V�ۖZy���4��5������7"p9j��gٷ����Yy���%^�R�Tn�� ]�Ql5�<����\�/6[��nڰ��Bne���D�d-���>́�*
���;U�V$�QӀ:G s뫧F�䐰���w�PphPnRՏm�.b2���Zt�i�q`�Z��
2��ҵr���&����Jb�2��Rp�5��q��49�����j�Q��7�>xq:"�[�!�!�����5r=�v���:��+j�G�L�Qe�Mx-d	n /T�@,�^}��6����D�{zwd��YI�(�|s�K�W9.�4f˭$V�$n��m����&��lȆ���1ݷ�k]M/,`ۣ�^%ciҨ(���ͳ,:�h1�B{6��^U��٥���Vuu�c��jݰ�0�vH�_Y�M
��'*��׻�����b��z�������o )Z��X�}���ʃu��F�� ]�T�w4��i���j�*T���ƃ��ǔ�$�e=���2��nL�
��%+"�1%�EP_A�ګL�Z���p]YR���`#��X�P+3r�eA�;l��i��Qg��a�I7��5�^��պ�����R�v)�5��ݫ�)�Z�s�[-3G��`O1��k(d�gZ�tXV�R��r��(�Y��U��|��T8h�5��h==���1e^��md��Ch��
,�B8����ٶAց�`	C����膶�E�);�6���<��vᡴ&\�̽��#�7o�w�T�5�mE���f[+��°��V3�`$%����a&��w��^;�����(�ԛ�+'/I擤�<6�J��o����c�ofUU�!pS9�k��/*	������^��Ӽu�d��B$��Ղ�,f4LX.� /*�
�+Z��*0�,J��� ����٫9Qf����c �Û��j�m�yRY�Fa�eVd/e捭��}��6p!�HY��5 ?�ڙ�3&�d�f����K%�Ts�P^������M�_�.�StU���+�$G.��m�j���eWf���P]1"�ksu)eZ���ә�GI�o`�E ��b���i����R�ee�	Kr�ͳk*�l�S��E6L�6VH��j�[�[��D]V9�����*n�s�|�V[7xj��[tؓ��Z��aKiа0f1�S<�x�akz�q��x�����h] (��x�*�m�䩃5�Nh#��WN�[T��Ս��N��G ����	�ݺW�l��W�ȶ����xy0;y���Ur3GS�le�W���gs��\
�j�fq".��5 
ޱz��x�=6���f�wk!���`DG�i�S(���y�k��%MwF��8�^�*{�0�e�k.�񤎜�}��$iЕ�H���5��d� ��J�ٰ�ܺW$˩�ex��X��h)�3j�UYr�!��d�tA�)��1�\B=�Ė;KH~)��&�.A2���e��0�4Z�D�G��oiBr���2P��X���"��̿�K`�$tji�GJ�"�ѷs2K���n;9A��,R��zYͧ��6���8��pwx(Y��pn�46�� ؍��ɹ�[Ʒ0ک���ԍǁ���3%��Hշ&�{N+Q����*��ؤ��ZC8�DmJ��+b�Q՜���WB���mn&�V�Ʀ��ѣR�Ci�h �[�y�=�X<�����wG����Ѐ�m9u��Qm�w-%6��B	x�]e_[�2����Z�&�����Qŷ����5me��ڼ�!0ʏo7oӤ%���;V�";��+Z����v��-��.�q�ø(PhayoU+k& ��3w%Ն�Hb��z��Ř�K0�2*K.습����޸!J�7(��*XL�:v�^��6�U����de��f��,9]�KkL�h��\�!VDZ(�*�S��mX�M.�c������)�Z5
T�0�BY��-h��N �\����Y#+�¥��-ډ�ֵX��xu٩m`Ŕ�ګ� �c�L�L0UA����h)�h̤�����2�i�o �V(�z�7`.�̸�F�^���̸�̳{��PH6tT۟d5���&-@M�@���:���$f� �5��{X>3���L2�m>�&�XL-:��^X��q#bͪ�ڈ�U��՘�нش�vb)=�-��Z&�!W���}ҹ]�Y�V�*hx4lh�eM��pLj! ����bG^��x�H�YʽWLiZ(by.]���L��YX7����t)�Qv����#�q&�Sj�e�H5�2�G@�8rU�ѥO���fj@�����JXQd�AP�)���U�� ʘ�QV�N���9�6 ����n�$�Ok]ط&�-k.�X�����t��9�����Yu�oV�ɵ��4�y�#IU�(s��b��7Djݺ�f[�u�<�[�C���k'{��*j>�oV�k��ljse^�.�Z�{��#��/��9�m���U+��J�^��s4��aA��J�߮� (M�tjwr���z0���x�9�қ�$,�$��XD����&�\�umɗ)�).H�{Y�~zf*ǣ(��2B�<f`P����?-՜j�����p�f�iw�3t� �g���E'��e�m�n�)����θ�{��6��,Hʔ����㧦��+&�-��
T�ٺZ?:�td
Db��P�Fc� �-frH]�s��|w����/,�����3���-�AUÖZ�	�������Y�'�T~l_�V�O�b[wx�,�ݎ������[�ɻ��[Me��Ļ,֦�=�F�Ψ��+dW�2�I��Ҟی��1�˃G�Z|��aht;�����A�έ;Jk���[�WW`ͤ;U%3b���u ��Lk�6��D:z��uW��5ۭ�gr���+F���´$�Q�������eY�A�n�Ei"��f�\U��9��k���]X�)&��%T�u6�E���E�"��Gr��ke5{���yeZ��i�Yg`�鬡��̙WO�FĴ�1o+��E�q�E�A�P�u���s��%Y�;����X^�̲�޽��"Y���c���[y*V�!Ʋ��l�Ź��n��F�D�2��G���Z����']�%�UfL�z����X$�����e^i�<z�ѻ<9���U?�E��S���ލ�7��٬QVl;�!f�u��ɖ�44%�̧R�!�����Y�q��뷓@X6ZxNm��
����֩�!�D���MSI��X���k6��*߯0F���,�L�5]HwCf�C-�[�`��S�A�m��[��!���t.��]�NXV�5���0�������"��\C+-ҙSc,,Q;{��d?7�b]�i���)h�U�u�W��2;ea�G�m�lJ�d?X�e���-�!V6���Y�x����T9�ncZ����V��F��	��6��+@��6R�e�uf���<���v��{ޱ�jH����4�j�Z)�
�s&�1e��7M�`EI���(��9�A.)1�n<O��V9xFۃũ�+]�z���Le;���xJ���̵���j�m�z�������lc��bd;)�{T��ZW��)�Ưu}v �SW�[O]��f��e[��pй��=�"�5�*m%���ЊVHV�ϛ� I��MZ���H]i����뿯
�F&;�F�T���Y,�$W5n�Z2^L$ ���mԩR:w�B��X ��G[Y�2έ��0+���f�wH��sVB1�t�0f��a�vM����(�LP��cL���aͳ{�V]僡長N��3�od3��Ѫ���{��r�L���R؏ 8n�f��^;[��[\򭻷J�k�Ui����IZ�2�̶F!P��2�VЊ6�5gۘJ�i�VkW.��5��:�sZ�Sm�U�[Tkm���mj�W-F��km�m�6ڱmW-\���k�ZѵU��Z���kW-��m��*�Ū�ۚ��U�m�Ŷ�kr�lmU���U�*�sU�ʹV�[W5��lm�r�k�msZ��j�6�Q�+ns[nkm�m����[�X��-���m��TmZ(�ըձ��Ŷ-V*��W+[\��m�U�ֵ�lmm�jܵ���*�5��k\��+m�ܵnkW5k\ڋmU�mh�ck�ۛZ�V�F�[mE���*�V���[��մmTkmF�����ѭ�m�mmnl?�B		�	!J����޹��L�
�+�43���n��LVGr�,%��	���+��z�+��;B����}گ:di��1+6C�)X��ft����#٪�`�a��:�N�5ӛ&Y����_�E�S&7Yv2���;[1��s���h!�$5��e^��m;w�d'+�����U�]/�WA7W��pe ��VS���=Ga�o9o_p�s7X�W3�iR�cp�@� ��hf暁ۻ!F�D�v�y2���j3Qi롆��Rt��q�8D��'U��SO���Ű�N���CRn�S��2?�Qʻ��YI�tE �\�w���R8n��mӥ-&�3��t�Մ����L唯_`3;udWOw*J���*��mn)��$���|�nnRz��c�R��n�����U�6��VH��Z�V�%��yXb�)�w٣�,��7s���"��{le�U��s�;���
�c���,Rwطf
��u�>Y�8����k��hR�uZ�����8ݨ.�0Ќ8`;�TL�he�-US��ǳ�x,ث�귚�ѩ��j��V"���8��޽��9�sU�6����1L0�Wt��圴��R�]���a����|�;D]�#s��O�+(8q��K[c0oe�OfTz�é��{em��j�]��:K{v�2T�Y�����\��y=��=���P!�h�df�E�qgYx�>ǧ�fB�]��!�����	�Qke�k���#��J6��wF[U�sF�7�a�ǰ<V��B-�i+�r���4o�t4���r�švl�����].�*q�[øJZi�H�i-���1f:�F�*̥����jR%�]n�&�1Z:��2��t����8�+�l_w}�ꭁ��,��ZY.�j�YEU^rT��1cű�P[|�"ԣ�t�8��I��w�9J�x����Ml��7��(P���ګ��J;U���nq����'�,R��D��BuM���Y٤���Dfl�Q�n���\�Xٗ�b�.��+;%�Ί\V�g���
�N߇w�m:T1�%�՚z@fķ9hV)B]ͺN�Bծ��-&:�q=Y|�Yv�b�6sy��q��<��]k�N�XζJ��+�����z�!��3�sv6���]AM�k$SY
���/LSh�'�k�@�/(V�Ĳv] �V,�b���E0����>Ök���.�]C��e^�YY�K6��n9#F^:��W��!��g�&�*��I7�ǋ���,+5{]̵��ޱ��D�V�V�#B^ W�2��SYB5N]�G���F��]dpau
�Gs�Zuw�G�͵1�ܡ����r�.<Nu�V�,�u*�-��J�l�8����4Y��e�z�!�	PQ���b��1*�m��h�`�ȫ�η[����bZ.<�8��R��[��T�]�`��BTB�Ս�zG��n��|�Հ�NU1DU��.�����v�ff�:�jݚ�θ�M���1��o�v��VR�eeJȺ�<Y�87�%��:�6�h�I`���Py�\�V���u\�p��Z#k%� Jڋb�݆I6���N�([�K9W�#��*˔��@�6�+6�g�xWQ%ǲ����:[F��YW��;�U=��c�]��f��!�2�4������bw��NG��SS�xɯs,�xop]w��'sq��Ȓ쐾x.���p�����wv�w,9E6,"�����mm��C;X��3�mom�ƒ�
c���O0w<w����V��a�\�[��B������I�N
T�A]Ѳa�6h��C�uR�(k$k{(該�9\0c�ڳ�Sdd[�UX
$wK��[4b��b�tC�@_kT�f��U�����̕{9�`���%��Bۘ�wq����,�w�o�^����`�;U��miя�֕v��̕r��,�ʴE�
I#;7l>�{�A&Cjq�̖)NY�\t�*h�gH�;zsK�I��˕gj�&[3e��f���T�&�;0�d,����^���A����b:ru�����F\��ѩ����Xꑺհf�I�7�Qe�L�:�Jj��o'q|�U�u�l���'(U�Yk��;-'���f����$F&��U��)�uČ1���q�$���x�0G��p6Q��G�o�ͬ�|�q����N�S^�P��3mK�*��8�tcxc�[�cf\�=�_d�t�g~*�8�)م����������ڮ���)�e.P�ͥhN��`[���X��Mv�2*��]��M+����Uf����Y]���eXu>��o��O���lg�P\�Y�vL�r��ݐ�@}��:�FJ���hȚH�%�#i�����I1O�GO�q�2���}G2��'�tIN�^JB������S+������݈uS��M���PT��ᒹ�;��(m�6*�!x��e+u�R�dR��k��Ɇ�*ָ:���9����.jZ���+U�\�����|�^�J7{�����j��X��y9�69kQߖd(.���!Sht<j�^I�`7B���!YY
�ј�D���R��s)n��츛�I5Uc �4ݡ��i�|��5A���;6�����c��%zr�%��Y:7J����9$C�J[���&����-L�������:��uxU˳w9�ۧGhѐ8D��UP��X�W�G��M��p�R�j.�<=�v]�8q�3J�S��A6�����U��)
�����t��;Y����,l��.�-�J���ֽ���\r�Z&2�ے���ӺdwlW}\�м��`Sr�tΎ��S�NW[+�Fj�mWJ�a��f�V��2��6�uI-	��I����vv����pP�.��oi���gw[��;����e�hM��SJp�`��E	Xf�d�:�i��T4�x8jy�nǍ�7!�qf�'Y*eT�+U��R��{��<��1�*�h����}9���"�9�!�#r�u,B���w�ר��h�uJ',�o�����{c+q�;��hP#]���#�ǁ�s66�<�t걤v�KxGT�]]ڣ�%f�] z�32���)v��O^�:
�	`������S�^WM�h�K�l֫57�\y�Xt�w��ChR��nư���f��=�D���-����i�lFeG�;.I�+j�up��mv����f�B�5V���Jvq.v6��*Rm�9u,���Q�.�Q���@�Et�I%�]i�$�4�us�-��*�4GpJ��+�Ӷ[���ڬU� )'&���"���1�ˬXJ��R�9�d�QzA]�Y��7�dCi��'h��u�4�<�9�����f�5�l[㙁6���Mր�%yiM�ǳj��+�N��5Y|�ݽv�C�u�%D{%�(Ͷ[z��ʉ���̖��fU�Q���F�������R�K˱r�!te�w]'�l�)#`#�z��c��讂� �*��p��l�@��Y`���3J�P�lK� �TeF�e�T�W��:Nң���`M�G,]�l�F�$�7���7��q��#]�5�#�Ր����:b��SqC]7�6Ȫ� �J�cRT޽��t�άʾ��u7jI��}�¢��i>=����]o��XӼ��N�
�nZ��8P[���f���pT��,<Y�:�t�C�T�z�lC�3�0P���f��u�-b��jK��^�/�V���X�Mޭ�QѢ-�95@k�
�m:2��r�w�J�Z䗠�x�p��r%�[����	t��4�6�35���[��s��y��t�_EV�S�\�b�]R�i�La�b���[��_3��j�Uo-�z���25������Q�9Nە��H���b����(�ncS^D�Kv>p���h/;_]��:5�ky��Xwr�N���B�	D��nV\q�������)�P�'�ޥ�}}l���v��y�V��+n��I��9riK�GL�v�m<\��j�nJB�]D3]>�[F�퐘%��-ֽ�J�˺5��s�REX�V��{1غ�ή�Ne���g�xs4q]�k:7��w;0�� 㷙O�'����X�j�և�B9B�1��)�{/�-�ł�$5����R�@!Ѷ�){n�ݯ�ٯ��j�aY�q�J��,�]��hqa�чm��3���֧ŉg��@S1Z�r���t#Ô�p�Lh�Uwi���t[4��#G���7�z(�4rҕ\��g
kt�N���G��e�in�F���J���}E�W��^ظ��	��Ɨo�������T0��3Jºo^�^1��o�<��X�(E�e<qۦū�+I���.o���{�����jY|k03����gS ���=��^谣�����H��Ug5S��:������n�HpQ[��^��q4�*�a�#/��ս�z�t~�6�K�|z�vWr�߅b�.�"�������o��ץu�z��J�Ͷ5�mmq��L�|E�7�)G�r�pj�u@�,�5�S�Rv�y�gd]n��Te
��u�I���S6ݓ��Vq�G,�p���J�g3c��e	�;��3pj7&�˺�b�fm����I5�3��"*�1H�3�c����{[�@=|�u�%��=W|̌�w|r����҇W^b��b�]�v�-��ǭ����`�\�1�V*Y�;S獡η.e$�%�
[*ݠ�jW�`F�fcq}U`��ψ��h=��2g}R�/:�"\4V��S�
ڗ��b��u#!w]͑%��R�p�^�]�]9F��`��G���|��zrk{q>#xf�]vjҏZ�ސ�T���jd>�w���7�/[P�5D���nt}��m�
�ky�uF��%�*��F��8*=��UnڱiN�ܘ���WK�������Y�m�h��דQͻHୡ�e�%�
�MC	Y4ev>��w�h��2U��5�L8o��Gt6��껓�o&r\�X׺i驒[���3w̾�떨		*�]WKBn�2�1��T�Z2�듹���fk��Q��j[���Gw���#ܹZ��A�!�r�),O�Tö�\2�iе_��ѯ4M���ˮ���e��L<���`�W�+n��ܨ�V��Sm�ݤΙ�d�1i�Iɜ�.�,t�R���홴./�U��kzv�h:��PW���ݫM�hL,��|�;�k���8�邃]���dף�6�39,�7�dȬSo+S0�sC��+ʰ%���;)S�G�
�m�h>�����j¬�.�6��%�4/� ������cҞ����ˌn���ʎ��aez9,��}�s�%A����5���vBAK�K����t�w�����FX6/*hgE���ݫt�ky��v�ebt���b��1��]�K;/Nm�ˍJ���ꐸI�QHn�B��dQ�g'f� x*bCe��}
��p�]��80�Ȯ3�^7WZs�ml�ؗL��t٭B<�nQdWahԆv�N$��F�Ÿ�c0#jU���J�dK3u�Ι�0n_G՚s�z����p^��`}}b��,c���tFf�ɣ
U�x��I�� 	ǀ�r�Vb�/G�� oٝ՘:�������v5J]�����̣��7x4�gi3oxmV��Y`���M�IIp�m�+5m�s�X�t3_lKBN�4��Y�F�����=��>x�5֟`7����D`��b���/�l�b��t齖t���Z��Nf��,7ú��5��q��FI�j�=S5�sk,���6�# -jU\�)�,Tצ�s���w$�-[���9B'X4��K��T�]��v*X%��(��U��-L�Ed�(4�v�@�U�Ko�ѵ]��'�� A�'`���g5}*]^TLƨ�0��j��.o��+)1���v��?��ư�v�Խηk��[���{E���[�1n��XGe��!v�A������K&�AG�Z���ʎ*黈��}mt7�׽�k�h�#X�;�U�N��+�>X�:��u�a-�q���3�m�ʱ�.]=�κ֦8��Gz�7��w�i��N"��պ�'\���]�`�f��%f�ۗϳ��c�rK�qZF�2U5��8,�%N!G.�B��S(s�=�ɝ��p�v�D�v�5��R:T/Mw\wĶ�8��7�p�4Q}�Z�mֶ4��,�Hjgg>�@��h��c/!8��#�wdR�a���T�T9t�u�ﯜ]MU���5K`�تU�v�����a�՘��}�����땲SU
��eAm���ƺ���;���!�����ɂ`q�R���,%Eٳ1qr�D����T�
�z���d��:k]-4�6�ۦHLj�}z���p�F�ś��!���S��v']�c�c�*p��¦u25���,�(ͳm�b����W��c��bUtܒ��0��]��o���M�rU�� ���tT�:Z��5���������K	�HW+z.��\M[xrI\�V�^Jo��ZF�۱B��H����3{���c֠��ٖpC}�U��z)��]�����'s�b�د8�bZٽT�,�y_tW�	��hF�t9;ϳ!����Y��7b�'�M�uH����yCs1����8;Go���M%V[�����:-퍺�6#3a:TT]���$�N������%��Ш��@�г7�5�.�W��F�R�V���������e�P��V�E;g�J],b�+r���
��*�N�5t�׃u˚��VG
2���lbHUs!Q�ٳ�U����(8Z"`��*%�(]l�nfyʟ4��݃wٸ�[���=�����1�j��zC��a�t����W9v�Ѽ Z�x�7�
AQ2<�U�7ݵk�cwֳK�m�2ζ�a�z�[����eu��8SrG����6���76Ɇ*8�$µ�Z�a���o�e􁟑<�oZ�)5�k0N�2�ctzR�l�L0C�/�$ I4$��s�����m�������|��܆M�[�U�f�;%��Ýq�n�vh3�I�r�����밂m �*�C��pP���5�T�b�wCF�ɹ�QK��ON8@+&����&� ��p-���,i��:����{&�`�`��ݶҦN�<�ìpm��;��ɫ�nG:�nU����Bmt�X��i�&���c��G�����w\P�:t�zפ�Z��έ�W8���n�GW,��݌=�]+ڄ<㛝�-�fn����H���]F1�r<݇d�9��S�s7��#�͏7��x��v�댝�]�u�
°�ɸNۆ�� �m���ly�,P�B�tm3�9�w�ڶ��׷<z�� �X�N<�������$�ٹ<�`�m"\X�{�g=f:���#���5̡��%i�v����eR۱tr�vMڧv|&���;An�-5��P.$�wZ��[�e�r񝽨�d3��y%��m�����1z�`<�O1VбV�.ۚ����^N�\��嫡�]��t�w;�qƔ7�l\��l�뮋�Zlհ�Ð5ta^XzWc�.��gnpe�c��$�]��ƕ�]�fp5ٟn����/P�g0Y�T�N1�-��ny�Җuv������h�cD��㞹��6M���7d���l�l���:��n�AtnTѻ7gYv�[���Ϣ�mήwck�x�vՉ7����aַv�W��#v�ny݌�pz=eᵕ�Y�U�n�V�۴F;vƻ��[ˆ�u�$�\A�x�;kK��ݺ��,x�n�3��������(��⇎�z�独���F�WlT��}�h����-U���ݫpu0�5ٛ�(��pR#/u����\�N�;vǭ�6���:m�Mַ\G[��]K�G�݌qQX��k:�\\�;`sCի�vw[.n=lE���=gu���Qۍ����#��9����W6�.�%���۞7sSź���tr���E\X��e޸���Ǆyٵ�ԯy%�n�d����̽���Q���x�ty��.۶�)�,sQW]mO/h��NSh���Ǟ2!v'������1n9Ƥڣ��qѬl���c=�c5�`Ս�l�u�|�����]��_.���6m�rwW\��H���%rq�tu���m�|vڨ��ݙ��5�,R�cn�{��{q�fJy6ʡr!�b�Nʶx��(8:$z���5u�xD���K�[�)�8$��nyν]gV5�'O))�mk�]��#vD���J�dh{�v�+�e����t�ی���wd�ʻ��N�<r��Ѹ�Ò��ǧons��k���B;v�Vq��l�4�)���v�����l�����m�Lf�q����s��G�+]��s\:�������rO9C�旚i��x�D����F�a�ny�88��S�a�G5x�#&ӌ�J�\�1렇y%�%�|���0�u�]t�躻q�V.ף[�n�hۍ��Z���N.C�]�l�=�sѧr�ݕ�F
c���7Q�û-����ON�ND�ն�ݝpe��Y:4����;���4�	�X��\<���%Zڞ��щ�ɺ�vFӆ�&��v���[���s��<sb��{r��+n'/��p��1�l$�	����.�n��W;��������f��'q�R�ٗ��q�quћ[���4�:��aٖ��7�M�SH��]���;:krjL7g�:�'K�
9����:�*��;��]t�{i�v8�h��i�ӧ��pv��l��!�=m�cN�d踊�>H��َ��l��«nۅu��k���a;n<��Wn؟$#1��<oJ�����a��dI�&�ؓ\�պz^j��ʫ��oS�' v�ݡCƜ�;\��ڍ�َ
{��/k�݀�9�i}xy�:������o:�c��9���9Zݫ��W=�8��dc�K�x^zx��ϷV�m�W'cu�q�׎��\�h9箶L�/Um��Y�L�xSF�x�"��N��-���I�[q�teN�)��ZdۨQ����qC�kۃj�<����Q�'k�}<�l���H��u�`=l;\/F����{	�������7=�vW�Sl���]OTd�GgYM��ۨ�v�;�v�`}XCgnD:+�;�v�gm�	��g�Q�G:y�Qv��H���f���8�wj�윕˳nsE<te����Z<tN��m�W���-۝�#m�>7n����n%������Q�m��jb��S�m�i7W-{\p2;p�;�����`�s�����d��cK��n��aa>�ۺ��=���}u�]v���Of�n�g3a��v�ڍt��֭Ş���b����]���y����G�(a�(i�;����9�a�؄��ɱ�zz�j�|��=�ȶ;l�����Mwa��҅��ǹx�"j�6�v{lN\sv18[�.�:�y�b�3�[]��V�j`

�)j�*��-Q������6����tv��E�>1�'0�Czv�����;|-��a8������qy���[�&��\��퓃8��G[q���E�����	���v�5��$�����7kt^�"�n�m�+k�!N��r�Y�[��&����l7�nl;\��]gڶ�f��dÞn�"s�E���]c��Շ]���Nyx��.���<磓;cq�C{[��n�+k�����6ƻ=�,�uv�.;8띺x5��!n����.u���6^E�n�{v*������;���F(9 C�Fޞ�2e6��!�WB'S�'-G8 6.��Y��8�;5�g��+�����Eɇ%pQ+�c�;88��s��{pm�&J�[;�a�]��6��(-�Ixp��7]�^zC#��v$.4�����gsћ�Y�E[O#v5ݭ���Լ�E\q]�Ƈ]g��TM��ݣs��ۧ���x�/$W q�v��T���c4vv �������G7�{%�^PC;�{R^�^;۶��; �\���ƢJX�s�5�\�oL��t�QV�øM�_9ʱ�7qu�Wf�`{u���@�j��i�]�6�$�X65�<;�G���2[o*�$]�n:�;��
��ЗO��w�&9�"��T<�SF��ֵ�S�mW.�����:^����vEz��=�Ca3�r��뭫��{"�>�̝y��F�퍷�\�k;o!����IE�eΙ��m�"�"�s<c�m�$�{B��=S���Їo@y�����y&a�M��nf�kGl[��!uX⭱�v���M��py�{�� �����'��v��[��wc!�S��*u���\k����D�'�磰�&\v�R�C7H��R�:C˻�������v�.�	�!�;�N��z9Cu�E�ۗsT8�[���;��\�1�g�1n������o7=�9���WA��ϝi��j�vӏ�ܚ�4�4]���׷+��7kdB��u�c��y�z�`ng��BN����@r�4�V�j�l��e�\�x��:����������+v��%Fwk��<)l�)���J�I�'!�/��ud6���l��m�M�=ٞ�籴u�5�DOfM�t�c���@4&74\�����n8��aLn�꣑��m۝�tޖ
�I;.�5=ң�J� SÃ=��;��{[q�'[n�b�N���l���g�[t�oGe�v=^�	�v�k+���<RM�d�����6�[�f�^��lp;q�NMM�c\�ͅW��:]�;R�LA:�	�i��.�K��1���[�Ǎ�Z�]J��i;-�pv�0��1�_<ڋn��S��bnwT�@�a�E���9_e�N��G���aC�<��|reڄ5m��HD����m�zS��c9�]��DU�[�[�9ۻ<^\=v"����3B1$�vz��kL֎�(���sf�ㄷ8���pn��<q&R��qm�nm�8�q��
�r�n�n8uvNn�sv��,q�qU��};��# F/=m�;�u�l�C�y��� rv$)'���Ɏ�z��6$�79U��pFe܆;s��cq�\#�G8����m�[�{I6����v��%�k�G/i���� �&9v��usĊ�;k��/g͹�QƸ���W6� '�nGe�{�{k��{���l������5�i\�lX����q�j�����v(l'v��p��nA;Y(�6���w�f�D�;U����hd�n7p��-�9��R[�ʹ�nw);����8�m�,cq��N��m�z��N;tv|�ֽ�^�Sn��'9M���ǣ���q��$f�qq�o`�f"�Ű���d��{�uڒ���I���Vx�3�U�Ǩǋ��1a�
��v7kI���4Tc.��z�]���G&^0sv�9�9:���$v�s�f��z+x����m��kQ`���wVM�����A�J�J1���2:�mX۸��[{n9�;���ОN��:\f��s`��h� �ܗl�F�F�v����:��!��ь��UdG��&��.�ˤ�<9Y�m]��AN�kx�Y��s�6-׷�r	ny�[a��2y&p��aʜTqz۷<��P��u!kQ^�v�^<�Wr=���
i��/��ú�zl�v�D�elc�Y��7�� ��5r�l�g^Kγ=Yz��$=�>]���%ۍ�/9�7�ݖ-�x�����Stym��O�ut9�h3���rjI3�h���ϵ�t���H퓧nn�f�6.q�GW�77Sn�9;lyf��W]�ǟYǅ!�8���Uq�=�bp�������,��^� Mw.='����l!ua�5��9ƞ���\#�m�mM�㎻[���X�6���k��Q��O�o]NxΣhl1�[yxJQ��n��Lq�7Q��S��(:<݃�/�v73�d�yf3G��\��=p�Mb����4R�)�����7�j=�8�a���ˮW+��G7iI;�
R�)�PHd���2"�wS��)s�$h	ws2�$;�Ā�D�C�2"s�+���9��s��1N�,]�SL�@b�d���&X������0� ˛�r�;sQrHPQLMN]ww;r�)4���2ffJ��M���B�B"f.u)�'7 3(����c�t��7v�#�wn��F@AF���XE1�wR�]�BH�wv!&!D�"��P��s��МݓBwgp��$;��4n\�XcF��N����ȂiK��4��1�I�B1^�{�9Ļ|��'l��>��i��!gv;I��p&���zޏ\:�+���7l�<��ͷB��`��`֛p���6e㞵qWm�m��W���N)'+d�!{v7\���5��P:��͹:���ͳq�/Jc����q��<���ܻ��A�V�����[��m������'[�=�l샃�6]sa'�b.O:�Qú亘��.8��qH�q�2�1�q6�ζ]r[��z,Wqq�hD�m��n#f]���8n:u�^ێM����e�b���0�x,s����vR8}/r>�z�ѧ��H�v8ݕ7���E�7���Z�{7�g�#U���t��tKz+������ˋ�[Ѯ�c��/ <Pz��g�Ф����kAj:�M�i�p �^ʢ�^ݦks��՞0��3���Y�{h���؛8ݳ���j��zs��{S���Ý���e2T�G7\��WV��-5����^,tu���Π�GXu�-O�n5ϟvg��8����m����=[�Px���v��ڞ��p۷Ltmpp;���u��V�T��P.�u�n�c;��+�6�T�y���nv8�NT����Uq61�a{`ݻ<��0�ܮ����;�9���.s�����h]���0>َ���;q�v�ة�\����j�wZ���N,t�e�^g�:_F}�]�v�-f7�<��M�;�ݺ�&�[n]��n���N7kp=����/=LЉP�	觘+ݼ�6��K��x�9�53��q�O[��h��৓q�ޞD�2i��j^L��	g��ɓ=	���&x�mcv�Uv����V�r:=�wG�8�B���)�<�Y8�y�c�7��k�4�*l�F^�=��oMq7\�s��c��uI��:� cb.j�]��Ň��ɜ��k�s��rΑ-�깶�W��F��m�㍮ك�:��s�wNܗnx]);vs;�:��%�:�{��۱a��웟n�'s�0�p.ܮx�۶y8gnwg� ���nv^÷n|ރ�s��x��݁x;8v0��7��G����n��Ǎ���@s��l/c ����r��ɜ�y�w �'��v;"��n7m�U61�6N��;d�/py7d�3�N��ݞ_lm��'>���<g>ۛdr�@�?y����ڋ,���̝���L�H'�d��>)[���n�S��>$�n�~�5����^y<Ϩ�\f5�O���=�Oē��� �}�s}�zҮA�{����X?Z ���ߣ�	���~$���i��}�+N�[�A??c����+�>�I�(@��d�}���g4nzu��3���@O^x�潭�*OP�j�z]e;S�e�4��ڊT�#�I��I�7tvUc��O�^L����3���w<�t^6 {�.]xq��RD���E��^s�G�^,i;�����Lk�z��D]��%іI���Vm_���{��}�~�?@5�n����/;î�}>\��L�s�S.<�ڋi,���=����������2{C��s�t���jS���U��s����+ȯ��7o�9ܱh�ywu]
)Kܠ����X��u����;;�&Cu)>�TmW���W^���p=���+5��|�1�T�� ���w��W@r�i�C&�Y�'+[/|��Չ�}�!����v՝��Ʒ�V}��c���}w�n���<�P 59���|=弖Q�F�ɋ�_ ;��U\��9d�UT��>��g��k��;�H.����#�A���@�S�tU�c�����U|�9<2�=X.q%��Q�̐m�n�Ӷ.�ֹy��m�^�튼V�]j���5��}Ln8TG���M��\�g�	 Oc���oy�8��Y��7#����Z��,D��^�s���k�s�<[=λB$�&s��	��sw�@;�u��s�ά�]�����Ǜ��\�[Iuz-zH4_��4	�qت����/μ���$ٜ�V7ؙ��g�+	��7�q���[܂���Qי�i�n�v�l�S;���0ڻ?zc��A��0u���#TQT��g�u�׫il�����6 |��?��_a�� ��������禍�vX?R ���zv���`z/"�����~$�Κ4�u0��\�����lq�ټ	�
qvK �p5�^�^�ݥ@=��֧]�z�� ��r���|��$[��o�Z��B��O*`P�g�v��9��-܊��k��:��h]�X�wa����H
�w�2#��'پA����A���/�I��o�ᵎw��c 6^*7m�,�z��$�{=xI'����3��od�ɴ��3��m�{]�I��:n�mr�m�u{�~��sF���_��I���L+��X�k�/�T�O%]
�7�ޢ'��/m�����hJS9���\=U���5�O�X�C���#櫔���QOC2��~�{�t��{��H������� ��n�����M�>�>�'�߉�.^|A$^����\��[w�o����#�=<C��b�QA�nY��Y#v�gsv��#�%(,�?VڃN�~��>ߴw/	 �� ^����;��������_]&�;��@��Yu��n7LP&ktp�{�;1�i-�(��v$�=��Y�|0_]�Mmx,>Z�$"���k�I�ӹ��c��y5�����V��ݮ��]X�7���D�ؤn���cڕՐ۞��;ω�o���H$Od{��`P��	;�8�s���*����$��w1���{������3,��\���yNo�sS~�w�J��*v�guw���t�K�޾Qy��˞YN����yጿ,�Q\y;�A#�^�d���o\��N��/wp��83#�1� ���l-:�̼������83@�<b��m�/�;�n��i{�m2v���:�v�p�w�4uMcTvp�k�Ɣ���S���S�Cb��j���vz�籍�՞v��vutm�f,rA�v��!��������\<�����t��=�껓�.2{#�t�`�h֬�۱sB 	ȳ�6z#�W"G:��z1٥t{��\�l������Ut��u�q�mZ�%vF�%@Y-�f��u�i�UX����A��O��0KA��=~�N�B��Jg�󙌝�0��BDZ?_׻~��A��약��T��O��ͺ�{��`��z�Y{sf��D�D��Wc09x�K\� {[��� .Z���87Վy�J�+=9� �ũ�W��U�B-"��ܯ9��l��������I�Ӷn�A�W#�e���b9�On�ٍ�X�k����e��Θ�{���×���l��ߣ��7�����s��^AR��]&� �p�eD����v���F��:˶:{e�s�w�
,�oޅ)QU������>{y�bg�I���-;�V:��x�ʚ�A�_���t,��DϱP����RZ��}蚝��[ϝrZ]ـ��C����8���8�	�ז'jc�Aұ�����[9�K߬^��ʾ�6�=��s~1�����vs�^Xy9k���I	a$^קn0H$�)lc5_\m�N���9�ck����m6�ﻪ�w��b���,�O&��ri��T���(kw}����X	>���o��y�T����1<�F�F�[$"�8�r� ��m�))h��Af�{�j��'��X?�wO{�l�G��{��pv|x�ٝ����9^-r��7Ӎ�"˝7��r*�3�]�VP�0r���w��'�}�*{;Zt���b'��TZ�� U��y���Q�k��3����}�#y�2{��zYފ 3޴�{;[`
}��8?c��$�䁤hQEU�c���� U	��`
�X�\�
�}��M�B�GW����虲��M"-�'U�0׽|'^���SA�{�Xa��SO����5D�<��a��X��$zǯf�l�A������wA9~aK$������vߵ�;������Ϭ�}욟�|<��:á�z���ak2��X��`�=�@��Wc0yx�Oͱ�=���J���&b�>Ӹ� ��P��3~8���{}�bf�uWj�ťw���U��&}H�h(4E�c�[
f��Zܾ�����o��B2�\�-����4��s3�M7�s�۫3����������j��^m�FDc�Vз�)a����30�^L�]jx�
�[`?tT�{.�t���{���rG�rn��Y���9�>��[���|��E\�)C���^�NZ����>��GNL0��Dϱ�;�}�v��t&�� |�ӣt(��s�r5���i�bq���6��Fخ�[���I,q���q9�Ul=��ޜ���JhpY�.ˍݜ߅�w�x_'�J-��p��vo��w�%Z$���{^��� �0.��rsҭZ˲%H�̚4훤�O�I�꫹��k��9lng�Dd� �W∻p�nS1��7	���܃�s����}�}}�C<��&�����w�$�[ݙ��IU%a������io��P��:oP*�����Gbq�vi�c}�zUr9{��/=oT���ߗ·��,�ߵ��V{�敓�9N���dF��Q8������&A5�e�`��mm�/{��	�vn��i���J���ٻd���!T�I�k�ܽ<]���z���^N� A}־ 
�MlR^~��]<��}��2`��]��U�b��mǻ�������ɺ�����P��[��|S�͟av��XA��i����m
�p�M[A�˭a1Q:�b����<������9[���O^*�Iי�wb����qխ����9~p�*i�!�t�ҁke����m��� �mw�Q���Ѧ$G�DT�h�`�,$X�t�h�v�h�&�p�Ё���;yn+�ni�8ް�����k���+�ծ�y��up����sɰd�v��yL��:���j�t����l��;��i���۩��ʆϤ�z�"��#�v;ql�^7fݞ�t��</Ag��w=�O>��ػ2g-��.x�ι2��1���v	���:	�[��Ww�?Z6����w�����0K�T�P���(�\4α�I׽�fci��'�u��{�H�GknYu�;S�t�ah1~��w��H��&x"_����kL �/�����Y�3t��C�mE$qf&��t��~��k�e �ʏv{i	��`P�}�P�d��lȋ��)Q��^��s=C�bɔMt��F���	w&�@'��ٹ��׺`I��^
�>��*��˻�6,]R�[�Y&�?_�}�E>R^+6�u`�]s����74�g�f�|��q�sKδ֟�X��]j)���n�Cn��Ó�!c��z�n�ϯ�~~�f��U_����ǹ����00q=1�!�h�I2�����;0�@���1��v�LU�s�8��9���ņ�������ƞ�&��eֿL�ק���G<�H��V+����쭐e�m���ϡ���ltG�Ҿ�U-�Z]��{EI�T ���`w����y���K���;���F��Q�$һ�^�ݦ �91B������#w��
��ٙ�m���o���J?F�TRG���C^�C��~��~�{F�	�:n�A#���Uf���e��&B�W���~Yg�nW,	���;�6�^�����eg�!nWb 	.��4@#��
Z�ȁ�:����
�s+/�de]a:��A�i�����۞�q�GS%PrAϤAeQ�1~�WI�U$*��毽��I��~�|�o����`ק>6�߷��c�� {�f���`��ӈ��$�O��^i���ߞ(%�ruLP T��o�����`��w�94x�~�&ֵ�?J3��P�b���4��s0'm������=����}���6���:_]���6�q�M�w���_�슋4��:5oXJ�Ǯ�=��72�_`׌���/�C�*���(�0�+3����]�:<B���]:�򹤋΋P�˱'J��wK^����O!���{�����+
u��]����Q�E�x�m	�<֮�9�#���W]���F,�v6�9���80�bev$W�x㒲Vy�c�?6�����|��¤k6�;k)��.GW���y�������(p4����ѥ�w��*��fH+c'���w�R�޸(8�c���V��$��xP���՘n����8a9��M��}v�渊�n�+���n���R:7Q�dZ�a��{��C-+{�sr�,x�����cJ{.�y���q���E��-�iQ�(�)�/��ꍌ�I�b�ֺsʟ,j�}}��@�dD�{6��Ji��V$�b���8��WŤmV��7�o��C F ﯖ��U�4�-5�X2��b�YB�SM��=W���mMT��*��*�D0k�d=�P>a"Z�e�xN:֙Ϛ�\��;��w���=�`���5�1<����E��A�2h�5����d��t)^3�m��e�]I-C���X�(�R"��ӡ؎wM�C�L�l�0UhPTUw���p+��lĶT�{�olUژw��-�T���:R]]�N5z4ַ�`K&�G�p7[���`Y��W�9��-�RWf;s;`ү����R���\ K��Ý���(�)�b�+�"i4��r��Dh�)LBûnQ���]ۦC;��wn.vF����4��PD���%&!��\�9��˒B���$i΄���Ȳ�J	Ή"��%,�I�K��Dd�7t�p������[��(Д��4ē"wW.p�9�I�Fd���wvBP�K�d�&�0����4���9�e˦��S;��$�F2`1$1�9Ĩc��d�I(� W;wq�dI� dġ�RR!�˔l���\�P��Ĕ�3HZI��s�E$b���t03I,�l�2dP�����b���I(�IJ\��$؃e
�=��8<z��4�$�s0�[.�]
�vI�w��}�pw0b�G�k������{_7�q�O����Kg��:���N��]6*��T(z?7N��xgj���x���fO����W�l߉�߼�>���֫by/
۫g���]��6�m�ͧ?���+�؂��G=\�Y@��=��kb�
���P���w���t_��}"��cmo���/S7�THꙉ?j�����y�gv4�
 9v  �>n�	���E%�KP4]c�B�ݏ��>�+�Ԫ����� 4O���S�����&`$��w@'3�eZD,�����6?<����V�
ORB��=�ͺ Ǿj|v��oI:�=۰��mj�����!rU�U�d@��mj�Q�٬,Mۥh i{�oz�F3;&��S��UyJ��{�C�k.sK]�����)��[�=��bi?c�N�����=�~Y3< 9ln���+:fdVκ-�n����$~I�c�D�N����V�:�Rv{v��E;�7PrFp0y|U�t(U��\���띣H"^�`�_L�����={>�<�����cfE٫����K��y�ۦ�ż��� ��ϰ�	����	2��4��O_��e��y����7�
Z�#�f'�^�~'��g�A$���Ӂ�N���	$M�o1��}��f&�����D��%�k�=]�mR�ޮ9C�~3<��4�	��5Ъ���=�Ōac�|��7@R�W�$AP�U�/t[���$�:d���}yFb�;k��{=��@W��6*���/TM��m��-�4��6Wz޷�n�eK�7졋E�@���{�$��-˘3$��s�e�����5faS�oS|}߃x��E��;d�Яm�Ζۧ��x���{z�t;���.M�Ʒo@c�5\c�3�95U���kԎ6G-C�g/<�mm�۷]�[�oo`xSv^{n֦	�0h��������q�`u�m��!�S���v��k��"ջmf�cA�Hv�#�.��on�m	=g��l�9�m����rS���㣷��Z�q��t:�mn2��v������c*�\�����6�k�9;px�u���:���j;3�����uHK�֜v���������&�m7�>�/
-7�-3�gf��6h�^o��<[��x��,QH���4��[�}��#Y3ճ��$��{t�<m̿�=!����^��љ�|ٝ�ev6[PA�5�s���H>7=�@$r�L嵮�o��ă3\�$���_a���J��*�X�^^ξ�!ӂa[����
�w��>g�С��۱�]X�	�d*��~l��|����־<�� }���<���<�ؠ��=��� �|n{�H�;��_���"���4m�cEn4�"�q���O��c�nJ�ͭ�Con�sE��L;�U�������܌sC�f����*���1���A��(����cJ���Q�{���cF!�4w��y�|"��g���1�F��C~���V�L	��#ַi�lz{���Ѿ��A�8�?~}��߮��R���N���r:�PHc�f����V��_��z��#%�8���ņ�7)z�0�;�}��F��|����IGAj��A�[2�g���F1�M(gs�с�꣬:�'����޷��hƌh��{(-�������F5�(5d`{[��ֵ����Y�6�|��!�h#�һ�A�!�F�r���bŮ�F�Nls{�&�ޭ�l^�w�c>�Wz��k ؆�4����*aa(�;��Z1�����=_s�c�����y�ޟj����i@j<�_RV2����5&�͓F�j�``��}�v�Ƃ1�W���D�o}���k���G�ﾴe�bPg{\�F1�iF���z�a�Q�3}���վoz�])�i-����y���T<v�X�M�y�yɥ�ʱ~�T`�%$�~�W����}����X�1��W2�kP�������1�����}.�����p����)������ ��$��+�HǃA_ǻ���41��n�[11Vs=F3��Q�3�{ү�K��g(�iS�F(���r�lCh���g~�z�b��m*�}�Q��j���oR������}��5��Z{6٭�LCh�}�A�<h#�DRﯽ����&�=w.�t�e����ך�����m�W�T�㉣+M,\3�w�une��i��uK�#��~�?/zhV��W7��4ʕ� �O>��|@##5}����bX(�0�����h����$޷�֋F4`�J�PNo�9��J����>b��1A�h��ݤ[K�20"���Y�L�q�oҹ�A��_;��ݝ؇�#��#&�9�e�I�M�c�oz�e�w��Q��j4�Q(�+��ƕ0�����w�r߳�t^a�(���hƌh�h�Q�}|�Ń�6�j?J�i+e09�]m����7�o��T>�����;��xc�.n��-�$��`�x��[�@�;e������Q�~]`xdh��;H�����_}E�IF!����m�c1�c��=Y=�5���}�F5���(�>���1�&(�>5�x���MmZ6�m�}렱����P�>�r�����[��H�������>�v�`c#A��7���!��|S|���#��}H��2�=�l�CnoLݠ�cg���bXҌCNWh��0��0��4UV�>��wr�}��Qm�&�����h�,aQ5Q��;]��2����ַi�mkvS�#Go��ܲ����c��h-�") �;��yH���h#�׽v�l�d`F�9���1��ћ����S�^����������E,��m�^lS��P}�nk�ݚ�@�Y}|��rI��˭p՚����|�����F�N�� _���4�÷�ݣbb��\��޵��lf�Z1�#�~�)�0�Q0��3�`5�.^�X�-i�lw��-��#A�N>���؆�6�zﴋb{�����*�>쌞zg�nZ�%��Gul�le��p��Iʐ.6��f�e�������gMsR=ǽ��o{���_w>��`F�ҍF�}���m*aa�D�;hƌ#F����g���5�q��V�yF1`�4��iA��=�`Yͷ���I��dѭ�����1�Ab7��ֽ�v�u�ށ�Ve�$��}�v��i���g���F1�iFhΏ�{��w[�gB�\�bGzj�bz�	5�h��g��4SF(#Fw3�bkPj1&�S�rM�����?o����I~M�8�D���n�YPC�D�G���F<��ǻ��i2oLݠ�bb���Q��ws�����7߹]��������XҦ1F1F�w���cF4F���=��ьP��m���/��)�ƣJ&���e%i���_|\f��������LL��_ԋb��{+��؇�_��tz���tכ��>4ԫ�A�[2�g{Y�F5�(�Q�a�v�a��4n�%�����̍�7c����t�nSֳ��=�o��K�m�)W�ii�j��g\x�If�ح��n��k��̲Lڻ?�|��kڢqI����B�s�'�w�vy�m&�kt�So,\��1�칳���<C�ێ���xth��:Z|�۶�r=w����6Q+�v���^.�lY뱇��^�Om74t���l��G�X��Rntf��h��-GI�92�ϞK)�����=�.ctWG'c��^�,Ǯ[:u��c�xDy����S�;l%��G�^����륇6W�OƷ������[�&���V�ՙ�y}/�����wJ3q�����w�-�� ��a�ў�e"�X5���~�v�`c#A�{��]��h6��e �PC�D����HǍs]ٚ��{�#�{ݠ�,b�3�ьCk�j������{�Su����Ҷ1F�D�+�hƌ#D#߯ݣ��iD�iKo��㚮������|���ƒ1�.-���8�W�Ki��_+ݤ[،�}~��Db�@Fu��T��<�g�?w��>�@��gݮe#Ɣbÿ_�F0��!���nh$�գlC~�o��eK�;�y��=�RWQ�+F(0�o��0kQ��6_}}����F�8�A����s>�N���W5����+�{ԋx4��{��&�&���f&*�w�1���4�PiG��v�iS���׵ǂl-�4K��-э�&�����ьX0�(��(�~����o�a w�_�������o#�Ut��H���8
82T�����ϣ�����\�;cH���s��V����>��H�~�K妒���]��ޑm1�Ϲ����$�#�A��]�b7�o]ن���2�>ƺ3��e#Ɣb0���Q�0b����OCz&��3z)щ�:�}���LQ0�[̽c�wF��=��i�_L���Y����u-���r���1��n�W+זj:Nw*j��1�w(뷪W9\m�:����2r��n���H@x>h�;���5�(�`FF?}��f01���Ƃ8�N�i��:{3Y]{�g���w����_-���O�nc,���{ݠ�-����ь�bQ���ԃl,�1F��]��^����G:4F��#���ьX�4��iA��;]��e0')���m��z5�vcF��w�}��q���m��") ��E�$"8�G9�v�؆�6�z���k���ݮs��̾{�q������ܣbb�|j�bz֚�[V��X�����)�0�Ch��Ϩ��in�fO_ƻ�j�/8��#���E�124Ƃ?Nv��6!Ȏz��#&�9�O?�>\��:���3����M�V*=�z,�8�����ͽ�[*�w��&�$ٷ�g�*�w(�`0#Q4�PiG��n��1�m9��֌h��4e�~�u�J�u��j����1beW��Ń�6�����%l�{�)��nh��������}�<bٮ��\t�{�]�"H"1�{�H6�`FD��Fs�ϩ�(�6�ھ����}E���4B�}oS�7�k{���hƌ��w2��)�lQ0���ԋbU[[�����^?7sUB/����#�qZ2��+�����!ț�^���Į���Cg6g�y+1��g(��&�O�5�eg��k[��8���q��>�޺Au6!�#���R[{O�OU������*�_����g:���>��ի���(�iG�u�,iS���'�~�э�#����-���_>�;�t#K�(�}��RV2�����!���ѭ����|�v�Ƃ8�6>�z�b�<qz�����"�Ƃ9Z��A�[1���ϩ�4�PiF0���ь0b������]�^���SӍ���wVܰ{^��m���u�ͽCO<�Gqv���Bޣ�7&��ùө�7�I��#mM�o�PX�LQ�b�#G~�}FX҃Q�l���1��#A���[�g}ܚ�{7�w�h ���r�YPCb">���#4��w�{�d�6��7|��l���A��u����|������k�m�n�H6�6!�Z;��֌h������v�b��iF�K/��{�K+��~�%�SW<v���O[�6��)�m�e�|�lD$=|��D�Dq����W����}8���^A�!��5��}HưiF�J0��;~����B����V ��Qg�o��=��}���Y���z|Cb��1@a7��(Ʊ�Q���h�&F!���#��5�Vw��w=��x�B�M�������b��2/8��啘�����UfG�;�rnK��D�+@��*�!G�G�&�^I�9:k#}�V=��}���C�A��z�o�9���j�Ԛ��Ԛݠ�,b��}�1��6!�Ӟ�,T��;���=��Ch�����6�M�3=~�Ń҉�҃Q�s�IZe07ϔ=���u���G]�wk���l�th�87 4BP���v�\!��c���~+ߛ���L�H9U���_�/��P`��!�3��QlC�F!�=�ݠ�!�w�x�y���+�ˤ[]iF�Ҍ �9~���G�k���z�&��h��߷�PZh�(0�N�̏�׺��+U�Q��4�Q�F}~���F�4���� �!�nN���)��ȯw�H�!�e��t4���=�v��Y|�Q����J5Q��ۢ�V�&(�h��?��*Wy��o=�y��Dh��1A����!��m���AL�~��:+deR�K�M%���;��+�g~��ngX��E {��/ � ��7	�v�2��mD����#�s�p޹W�K�!��a��v�a�h�o>oZ��鹭��-щ�7�fP[E�F�&�=~��McKG^�>|t��ќ׳�[`S#.g��1��#��}�n�S��#���Hǉ��������b'�Y�}�?)4���U�6��0���ܹ-T��
=w���[��0�j��oBww���D�k�
�u�}�m�����Ѵ�b3.�8X�I�HK���v�ot�em㘻dXE���ژ]BBB�B�l�ؽ�|N�ay.t�:�1m5H������ejý�D� �e�v�����VI��7{����[&V�;���\�'���9�PZ�u���6[ݮ�b�/-��8�:Ҁ��0��܉��X/"���y��]5ے�ŵ{� ,1 �����8���^T�U86�8�7Vd�e�ݲ��neIr���Wal����Ý�:������7�WT��=�&��QΎ�
�����9�{��e�tr�'�r�f0��t]Jgc�`�ڻ�8���d�M!�h6.e���u*�/�e-�B��$.jK�b���f>	JB\q��'����:!C���b�6��m�!o{3b�%eP�;��^p�U,�Q�UoA�2T���Ґt��f�h�WXi��2�v�͑�2�T���ӯL�F�s3B�f.����3#�o�d��k����u�N��(ٝ}}��%���{�]Ua��31�*��P>]]�C@�g����S�����-��c�g�d'����8%��4��Q{�s/��:OT�*{|��Y�V߰��&�e�@٪,C��)}���Z�=v�.^��YnB�|��]��ohx/ᴒ�2E�e����;r�K�Y�M�u�9Bď/-�����_q��{qW�oc�]�����@�I$~$��D9vEݸba��,�1��r$�6wu��1�3b�"$�!�DcH%I4s���\�$"�$�2#L�bR$�3%2�R���,�"h���a�)�Y�0��ۻ�Q�̄��P��4�)2a	&�30�L&��330a���d�H�ȹ��H�SL����v��P����!D�!(1 �Q��w[�(�3I$��4L�;�P"f&#4ҝ�#���.��&bɄ�a��2IC(L���ƊQ%1	1ݐ��̔Ѕ&�@Ȅi�&�� �]�!DE��d��9�J�i����E�]���B*A��\k�m����U�pU��}���c]n�m�6:��"��qp;�M�yF;���2�L��m���f9楺r�F5=8�p	�ڗ�i�y:���Tz�����p;X��$q8��m��j�5t���h� �]n��F����vۢ9ݧ���m�-dN�y���+�\����l��<��r��K�+����l<��ӱ<h��Y{]V�@c�k�@�j�u۷d-��w ����Nm��)ǭ6��\ח�jd�S���듗,�j��)np��^M��֬me�*��(�d����k�\A���@�<�磗[	[���U���gn,��ɺ�㓐z�Ak��sö��<�rn�b�nك\�Q��w.3os����k�t�n�Y��n���Y�l�ݭ�,�l:Q����QW�nT���A�sKϢ�WZ�.��u�7@U�����Ϋ�ٮ�p��v��m[���;7���;6�|qs0A����Y��S��3	⎱锪��BȄ�g�8	�#Z6w�y��'���u׮�:�&���/���v��Uv�^��3�3�os�Ԝ�\�r��<�p�v-s����q�e���pm�l�|'���S�5���n�p\;3{;;7Ղ����{��l͕�+���͈.���^`����c��z<�;�����c��;m��m�.�)O[�ہ�.��@���9���,�t����ɽ`�nκ��N�E��=��ll��Y�8��O�MS���.�38�9C[[v{&�ع�1b�!ۃ\��*u�P]�۪ݞ� �i���<+�:���ŋ\���v�=\�x�]vt�L6����v������]f�<ns�Ml�.�x6u �:��&����D;6�ݹ:ݘ�'��,���\`�<�YGN�`��܁���nz�Й��lqu�	Q[uv�����8-����Zӂ��kt�Z����5���kI�7�{����3���侫�B�ͻN��U�}]c��l늞Ԋ\鍢�n{8������{n<�Vw\���������w6g���:�`8�ʖ��z�;����Z��el�v�ncb�Ƣ�r�)U�6{�t����ͳ��H�H�[��rf��)�۲[vs�q�]�4�7A�#7%�'D���x��Y�\v��5�ڏV��=���mpF黛8�v�F�ۧ{4�\�\Y�)���`�۰�gɦG.�;��m��v�9�@�ډdQ���I�p	XHI��V���}�l��M(�Q�s�E�+a���DﯿZ1�mپe����������c�X5Q5�;t�����~�܈(RUqm����Y�_��[A��D��o^Ӛޟ]X�3(��$ ���G'���
bڱ����F5�(�iF�9^oZ��U߲�1��J��c��z��ڴm��#}߹AcE�A�b�#G��}H�!�1���k��k�~��k�]�0:�h#���� �\�I�_~�c����m�C�ͻA��ŗ�e���=ɿ���6׆�j4�{����V�61F�r��"�0h�h�Q���h�+�38����W�X�iD�o��RV2���Ƭ��jl�����F�_>�x�D�$=|�����<�����A��yh)����5�_��cX4�Q���h�Q��V��Wq�=Տ��~l��5��f���
�OmƱt<��u��[�;t˰�)g{������]#�[{d<�h���s(-�ؠ�1F�9}��kP�20!��v�`c#AUߵY>���6�}���8A���F<A��MX����5�k[�e�}���c1��J5��N�ǚ���-�~��g"z�;��$Hv�B������:��iT��U,�3V�B��"ӫGǆ<O��ZV�w-��BI�X��̤��Q��D����6�#��ݣ��iF�K���\��k��o��R]L���ɹP����Im����{��c_��@/��QyF!�4�F�]����q3d�ﯿR-�Q�4������(�>/vu�7��kjѶ�h��~��ƻ��b6�6!�_����XҍFF��������4q�s�H+{��u�|!�HDW��i�7�};�6�ކ=n=�A��ŗ���L�iF�iF��n�i[��3��:5=�i��h����F4cDbL�s;F1c҉�ҍF��n�S���u��I�}�o&1���\l��ɹ׌�v���!#nGn��n��L�����z�U�¢�K妾M����4�<h ���g�� � ��4���v��l�VÕ���ew:�f���Ck�ag=��bb��p����7�l�"�0h����M�F*�������N}�g��*��Q��4��`FF��=f01����!���t���j���{����}��{囙�|����osZ�K���-��fz�f&j(�6����S�Zb��]��U�;����Um�ǚun�Mq��rE��a� ț����{�n+M�pF5.T�G[��N�����Gh-$���u�[[�`�}�B�9�#��Dh�Db�����c&��(5�v���wc��pAB�r��m%��������1�=�뛜u�GM�LCb4H�s�QyIG�8����[-����}H���~��������M!�Z�v�aT|ڄm�*L^�~�SHi�mr��
����o|��6�����8�A��;{Aj��"H����#�6���sRs����,�����UF�����8ݸ8J�0�oV��u�
_
u7,dx�ߟ_]��@)������g���ܣ�5J1����V�&(�1F����"�1�4kx��j�[L��=F1cҍF�������[{�z�=�oSd��e1��̺�4�#��+3�։�w���6!�󾭠�y�0#Q����F5�(�6����,;쫢؆сx�oS�7�=�f���cF4G���ALCb��=}��m,�207�w���;�����[�l�1����;{ALC�"4w�ϩ�k^osZ���%������Kmb�|����|�J5Q��͠���1F��_~�cF4F����v�#�����c�,����t*���`ڪ/EM�%�=�qu��Ю�T���B��0ɩb5����n=����^����cֺ��I�cK�5Q���~�%i������j�֣���ldh�W�A���I �~�Qx��������u���Du�s���h6�L�6�ϻ|���`4�PQ�~�v�a����;ݴos�޻�Q}T!X�n������h�9�:�%���e�n����-��\�W�#z��{g�Mh��}���b�#F��}��kQ��6��;c���:^_)9��^�'�G���Z�!�"#�_~�cƂ8e�{����H޷ݠ�c{;�c0�ҍ}�}�&J��W~�{�m��&�0�Q�b��_��cF4F�4F(�{;F1baPj4���^�췽�z�����~���y&��B�9�̎��U�r���=\���x�6"H}���D�Db�e[�[��sS;]A�t`FFj�;HưQ��Q�L3��ь1�4B���'�k{����ݣ1�=����w��|9��#XF(&�7��"؆��������bA�4���� ����~y's��pD��w��x��=�e�95�G�jn�i������b`F�J1�s�E�����wZ�������b�}^�Z1�#ؠ����1���(5�:��:�U_-^�߃�`e��w[!Z��:�Y���63�ۢl3c&#Ik����ݧs�],�O��o�nC�r��Z٩�ނN�fo�{)���G#�}�������~8N��s�Qni�����u��u���؈V���+�:�Z�a�ݽ��^�u��4���#�$y�m̦k�g�9ڗ�l���;��	���]�wUٸ�3��vv7SȻ��crh��'dk&�&�4�l���밓�!��I��jK6V�����ۄ{Y�ۢΈ��ɷ�%njx�6�kq>�;no�r�<Ѱ���Շ.q��]�O8n�η�������9��9J;PKtJT����w�i#���:�����h0x�6"����bDph#���ݠ�-��g�W3uߵ���e{�r��`ҍA�A�}����4C�7g[#z�{��h�!�M{�)�lU�M����/�+�|��u�[�r�Ɣ�20&}����F�'��9ۤ�r�~��V��ϑ=Ͼ�c��G�顽�R7�Ƿh1�Ş�e�L�M(�CJ?�{tXҦb�Ch�Fs����뵈����l�o�[&��(�~���V�`E^���S{٩�zq�vS�#G����zk�'kƍ>�1�lGĀ^��QlC�"84�k��A�X�����A���)�_z:��j�Դ�(�0����`1F���܇eV�ܨu��m����t�7��4SF(0���эcJ������G�������c#n�ܳ��D�A'�t��r�Dwٜ���ɲo�����E#q�
�o�6+z�����渱9��;��uCS���q��?�\o��G&�BkRo�4�1v����5��(�9�ai�0��4C����8�8��[�nOؼ�T�2 o�x4��0�(��J&�|�����������H܏oq�lݘ�6��+��#�S�R���.�����.�9V/W�*<��ۖ�;�ˠļ�}	�Z�v�x�������Y��;�BŊ��T\U��H~�ﲋ�F!��s���6X�����E��ҍF�a9��~�Z+������1�1F��.���zZ��{��m����-�0�Q�h�3;F5�(�`A�����ʵ�_�� B�Q�Q/ݺAapC���g)�ώu�ozԍ�q��f1g��F3�~�w�ߞ�'_=�:�4�PiF�^��S��!�frэ4F���3��ь^����w����V5Pj7�w�������M�f���#��!�z�̠�<h"q��@3�_h��!�}ϵ�ZI^��}׭s����)�{���!����{��#Ɣb�g�}�[������~��"��;-���W<`�9&»r��'g۫3�����y}/����y�ooF�6kp}G�h����-�0�Q�h�}����lC`Lﯶc��}��r��������
b��"=���F1�]��X���h�ԛ�e�_{3�c�Ɣk�O�m��M�Zn��J�A�0�Q�/��rэ4F!�Fg�}��a�ҕ�rߟ=�qS|���l{c|̑�7�q�lݘ��F��/���I �z�E��lCz���W�߾ܣ���n���Q�c��=od��ߋ�\��W<���-�Wb�9����)��E���U��߇M��N�8���|�5���=��!_r���S?0#ڀ�~�?R1�lCa�3߯�cb��wL�����F�-�7�{����u�rs�̟g�!�`�4_+�R-��F�_��248�A���� �ú��s=A�~�}H�!��w��c{֤o[�n�c1�/��1���A��J7�v豥l/���5'���\X������m4F�4F~���b�aQ5Pj7�v�+L�l���߲�f���u��!�'�GD�����]�c����3�nݥ�{<�nu�z`��__}���-��~)�mV��x�A�"H>���b"�rsݻAL������7-��.M���\��>���F5�(�Q�L9���cb�1�=�{�ѢoO[��cF4F�Y�&�b��ϻ�Y��lԧxh�{��汥�C`EϹ}���`���t����/믽o���s/�G�^�����G
�c�m�Mͷ5$ݠ�,b�3;F1�iF!���t[J�F(�&(ѭ���q�:i������GX�����g����b��b��t����}̑�7��zٻ1�m�Wh�O�;�z�y�lE����E� ��7'���6[5s�g)״���3�z��'M�6�A/q�`"����<]A+D�\�r���� zm�ɵ��9�Y�b���oEf��7/�� > �y�ɥ����6����c��{�ފF؆ߵ����&����cK|��=Q����.� ������[F�8�A���� ���G=��F1��ٽ�檭��~w���k�r�m�x�5�nv֕�q�e��ۉs�=����~��fs��M��9G_�K�~M}���Q����(�M(�ݾ�`Ҷb� �!�e�ьCh�v����#LZuϾ���iA�҃Q�v�IZf4���s�,$�K\b��Kh/f���4�#W�k�N����QAA�4�}����X�����e�m`ҍA�w���s���8�{�y��(�3�~o[z5�[��cާ��>h�!��=��1�iF�&F�������W�o�L�Cb��r�]AADsٜ�c�*��2��&�ۚ�n�i�1{�ߨ�W=Nߧog\�5I����Y��M�۾�m�=���v��GU{��S9a���	��V/4�y��H/���/����p��߹nz��vn�ؐI!ޛ��9�>T@K}�Y"�:���
M�������ue���|`�~<�a�:hz񘯫_3�D����\�r�[�S,�%��		$����z9�"�sQ]��N���2Jܬjٌ��u>�H��nےZ�1��ҙ9��=��p���i}������7l�uOrsv�+��v�y�����ڻ&禳�s:�tZ�{N��K�y�2�l<r�yܿ�|Q��Yj�����î47��0�Wy�۶]�<��lBI��s��c�N��n6JxW�v�ث�<�p�<�,�p�i�[����u#{�0�-^�X���|�Ҏ�����з]cH����~���s�:[o�:�;�����ǵD�$��m?���:���U~�'��Iɼ�,&���Ɵ��9��5_Wh�j�I$�잒 ��ɲ���'g_���+}���)$�1Ksf���l> �������r�Y|��}��`�g��`>5�k���3�Qr�������lh�{�;�$�^qϡ4H���'��M٢���:��W��n�~Al��
X�u8.f{1` >>{35���|�Z���o��I$T��� >Ϳ���J����3��0�˫�9T�2X�B�*�F�{n��ݓr=����G��o��6N�*����c�@ [�����I$��7��]���
�ۃי!���3� ���%�4�E�4�����>�X��=+@i�~f�i�MK.0�>Ǜ",&�jQ;��o����2��-נ�δ5�.�̍�hh��y�\��E�����f��uJ�|>|ٷ���I�jy~I�I$��;�" �_)~ֻ�\�`O�wŜ��U��f�f���$�;���&��w�9�ؼ���Ʒ�{3 ><���Z�s�,�Q���gF.v0�������I5i�� �Hr�v��I}=�;��N��{�������|+�����R(�,r��n>�J��$�I�}��ͯ{w�,�g�83�$�~m?� ��n� �� 	-C<{��������%,�V���hڥ;�P�\���e����l9(��e�Э�Gs�Gg�P��̗�F���|7�`����&�ʵ]��^�RQ�΍�� p��h�� \d�NB��E{gI� u���qK�^�O�@4I��o~$���!$���X�����yb�s�Vŗu�w>h�H�<�$��}�],\��۳y�*) ���:��.��֖1D^�2�7������\%)���fYCUB�7�y`vȞg4zc��u5���뭮���@���9+U��j��B���%`��F�@�j-�v�=����7��25��,�<ݨ�J�	e{ѩ_!�<J]���n�V��r+ܚ̷��t��X�+����V2g�]
����9�AR�<���:m`6��!�zol���C*��kvS�q�M��O4�S9x�vfv�e��X�����%ob9SF�mILA��.��C���VBǲ�����F
�ݒ�|�g
k3�8Y�����	�e�%���l�X'�U������&[�a"����[���5}N�Z�|w:�#��ǵYPhX��U�u��� �b�D)� �;���)�=Jrh�2̜�Y��f=gP%�v�j�ߡ�M�O����OVe��*�]�R�[�X7�%���v1����5� �bಔ����b�Զ��|R�X�I�(w2Ł]�����u��J�9�w�L��c;V!���壌�N�& �u��I�}c�]�v�e�M5�dR֫9
+wR�[��۔.�T��s:΋��͜�+���b�:��[�fsj��Ӥ$U�em��V�ffev
W�I�P2�V�tsZ�.�j������*<o1��㹫!d�N�F|������+����n>��8h�6���&�S�߫��@���]�r�%����wr��]�18��"Hh#�4�pC)�r�FF��N��N�ܺAgqĈ�"!2H�L�:@�����2f��C)��X��2S\�wt�2(
�7wpԻ��ۂsp�L�@�d�e�sv"�\�r�$�`#i!"Hь�2CbdRX"M1QA�@,FJ:n����PPP�I�h3"�r��pL��I�I9p��I��A��$&��"�F�!�u(�!�d�Q�h���Jf�w!Ԅd�a�Lb"An����c!b��L�d���d E��˯�G���XTmϽy���"ڲE�4UZ���{���,c�o�.=��<97�@$�<�H$�kڹ̦-�[W��t��z�5=���̲r�]^ct|�쐒O�����dͶ�����p����d�'��6$W�v��b��p~i{�7�Р���1���@]��P�r;޹4�VTړ�
�Ɲ��!���FyAE��N�W��>� ���7����I���{T2J,OF����#s0��˪�滮` ��<�x�j��q,���?o��%I5F���d}���U��4�.[�&��-B
7Q%Y3�^����>�^潬X �9��-/gV�=D��MOI�%Q'�{��a�=Ȼ���+�j�A�}�C��X����Nq$�s|؄�MP�^y� ��Mں�+=1��몑�,��?w���W��z��;��{L���)$��[V���iֿfO���pkΚ��Z�tF7���GIjf|>��6�~�7��`k��d�����3�|�l�@���j�b�}2� 8�Y�'���I>$�~5�y�ď�7�,w��|�.�r��1�#-p�Z� �6ᶠ�U)��,�Bu-j���X;��l�nV�W����y�bQ V���d�$���2s�w�(���$$�Mz/7L��BˠR7HJ'3��y�o����=�t��o�ߪI&�$ �y.�h��W~����繙���2�0��˕��� i>��I�O��ŉW,��� ���ŃlG�;������lUU��{u��jȤ���$��ǘ����f\H �s}�=���U��x���{�Z�=ؽ���X;jˈ<3�� �O��9	y{��	��(��&���i�k|�I	�{ӌ�N�o��[3���]��'������������o6|��
�ln��!�Mf.�M�,�-8�MFn��p��G�����+��琄�޹�d{ֆCa�kE��F�[5WoK��q�]���7�ڰc���m̙���k ��'���:w�<maH�m=n^]�':�9c�3pk!m�Ioe�&9��m��\����e��Hg�9����l<���gw<u8�y;I��)�4��]��L�5�g\[r�v�#a�SL�GQ��f�|��D[tI���ދ&1�y�]���r/\�MF۷[���eٯ۷�^�yl���քź9^-����뭋��Jڱ8�J#_�6�������[h� �9�)y�hF��[��n� <���KA���J&�nV�R��{9�	�&Տ���UǤ#��&�$�k��x�|�7	$�ʤh[�eV�k�Z�G���n>�o���7�l{��$�\5��y�ė�%��D���{��)�e�A�*�r�ύ>>~�׻��w��j������TN����I|�x���g�-�T��3�1-�/'���S�IVW{��c�^/��U�L L!��$��t�ԉRNrBI&���n��>uz�Q����nm��մ.�A�i�Fn:��炻�#��ݢ�r����躐�Х�����{�䀢}ޚ�$�<6r�D��Nm0�+�}�f}��.{=��`k��_�N2R�n��zn��K���_Nav��Yw��vr]*ޣ�#îj�*W7��Y
-ڱ�����ԏ9� ��e������1���=�*#M]�7c�iz��> }�7����u����������vTh%�a�F��D�����8�U�.ɼ��1���#�N�|�?�P���\U,ūQ&��[��HI$xGɢ��c�
�(�� ������~y�nt�]~%��l�� �k� �5e�}�k���Z��-} /��+�5�h^<5yj&�$�o���ft��!���~��� �O�� �ӤN<]�7�l�ژ�� � �e��D�/k��ϴNSvN9%��amL���"K���W�e���+�jS_���I'�?'�&� ׎�x蕫�R�����ּ�~�I&��3F��R��թ��}�����/e�_ UEKf��߉ ��� ��swF"�U�}Η�3�>�%����X�dv�f#�}̯���,�a��uxe
}
t�.|t;*���!�K�-1n,]��	'����\o(E؈���8���j��<�(��u5V�����7?|�|>����������� ϝ�f�k��Q�[���l�Γ��W��pUa�H�I4��m��/����#����a�O�o<�k�z�h,����nx������\�ϸ�&�^�(��,��}�I ������>��R�
q�@��~.N��X�;k������W�����U��t�V�j5�qw�ب�Br����1hI �kݻi$_?F��%�w�[��i�}�oC?p�����qCF�ep,d�i��wl��ƕ1"��<D��D�J��߂K䟺=�	$��ٚ}T5X�\���5���9��=gޛd���y�I ����W���$��tZ$������[B�V$*�l�d׋��{v:�\|I%x�7���&���I� �=�P6$^x]��=`oq�j;�cH��M]v��Sen�L�{o��Q�A	]W�
���}���d']*�u^���j�~����o�zs�bT���)F�nV�R�Ϗ�N��M��a�zy}Ú�~�zݲMQ'���	D�>��ر0:���sWu�elR�喂w�T�=
��\���9ܼ�w99�Uޞ[��g���~~����Ok�ۆ~��� 	��r� �'�}��l��[�.i���Ol��	-<�b�N:����N渨���7}m߆H��g|6�K�}���$��z)۶�	����$1�؞7��������:�Vk>/��oillA�voY�o���ee�Roex$�HOw�w|�I/I]�sz)������=O{�ם���P�א	{��7� �����|=ǵ�~�u5�V�I���%o��"�
��Z��G��3 t�1<�^U���d�Oӟ����D�w\N�I%�ݴ5���v�j����ęƇ�E�o��l�ɪN��05Yb[���(I%�:��fT!P��2N���|�CƼ�W�|> =������dڦ�<�X��vȞ�=�M۝���Y|�类b]�u��wm�������;ۛf��GS����n;O��l��Yj`��U'RD���=�����]��;�/;y���cFun
S�s�����Жy�`�rJ��8�ًg���ݭ�[Q<�|x����v�n�ok���G��t<�<�j8���œC6K�m�5v���m d��s��:݋x3��t�ڑ:����@vy���2�s�����C��[QKu�9�߷��@ �{7�� ��2bA�e�5�?�^׳��K�����G�UA_ƪ�5�������h���i)�97�$�	)鑖I$�q�o� �5��Kfx��g7��]��oYz2���U	˗>5�M����=��)�=Mλ_9ⷼ���� ��o3�0�wz�C�[��7�]��^�'o����-S<ʊ��	;�Ȁ'޿Gn�$��N�*u�;Ɂ��x��C Fs���(wz!������o��{�H��f�Yh =���$�	5��'R^�w|���O��~���z��y�-��ӷp��'\��X�'�h�V�_��Y޿v+��}�9�}I$�qNݵ�D��:>�S�a.w�ٽ|f�;� w�w��}��{Q
9[�/1���I	�l�� �5K^��ᗚ�R�1�+�Z��;|�if��b��wC�kd,k�؊��!,(�ϯ'P�0dn�H�����[`Ѻ��*���{����b\�=���w�o{@��>�;��z�����\�UAX&��w0/��S	���7����̩��b�b mOi���A'�;[�����lQB�W��,r�u�Ϲ��=+�H�����	&z{d��MN��=����}q ;�o2�\������ӹ�)�ӻ�H$�^�Wf�J@<�������JV۷�&����ܢOĚ>�q����GW�3���נ��X��8�u�^���M3�Ne�7e�kc��ε�접�����=��-,��|����������=����� ���1��_�����'I(���+hS�:Q�����y�����qƙ�<$�$���>$�N�� VT�����6����~^�s��l��n'-�3��7���9���(	 
�)�e�ޯu���O:��r��������Q�֖�7;�-�pDT��"�ⷅ���3��N�۩cR��ce���l���ys\�B7�>�kĒHw���� ?o�3!��]�$��ԔN�'8�FPJ���y�x�7ѱ	���� �^�v���l<�ǷJI���������b��UD���;3\� {��y'hυ#M]�kޞ� ������� �t��'|�7E�NUj��IѧU�j.ڶ�s�8�f%�wm�=p�t�.^8��
�s���27�t��7���ߦhx��vwy1���NI������I%~$���۲v#��.��˼��>�x��
lP�G�c�$���Y �=��	"Ǹ����Z��|΁��_2V�Pt�3oS�� I'��"[{�����˭~��I>��� t��>����aF�GQ;�l�.�{_OWK3}�h��~N�$�{����NlgI��Q�Z�/>�v���V��S���R�s��x�{]m��v���b�	��w�	�sF��+|O8m�}�����}���%�~�~������	$N���w1�oy�P�~�9��o��4�`g���$�$��F� ׺N�|N�ji�y��xj�`[ZR�<�#q��Wi4h�ݴ6�p�w8��M��j���{���X[#"r��ߦ��|�K�{�m��IN���)yFw�\�ߋ���A�|;�ϕ"o�s��X�������K'��6�P���O$�I�;+@I$��t����%3%���{]\�Nd}�{��B��'-�W�p���I��zNs�MI�H�~�3}=�<r�&&���E��t�'��6��L�"�#3��5̻~�S�;�C'� ����K�w{w�I�^.n���G�l��ў�J���;��UD�c��$ ��9��U�o	}|��큈����I�'I>$�h�Nm�H���SݷSy���MԴu�a�w���W��'�9�l��jT���������#���� �T�VsW[2������3B�6YjP��z���p�ټ��o�5�0�V.Kuq]�nffX���u*�V;���p�|�X�'+ћ�m9�^�ש��t��m=�BI�05�ˡb�#�`^�zVѰ`��Xy9�{K�$��Z��t�2�p�k��U>Y+�mӺ'�V�Ӗ���ZK�W��f��>�O%�9��C*��Y����c�GU��e����]��3܊�hni�E@)c�v�b�P>�����p7}t^:ҳ�ˠ��	n�*j ����t�X` u�K7oC�9�$k38�L��;S*!���n����X�]�C�w��m՚xN�r�,"mMz]����;�Λs]pY{�US�*U����.�XG"���N����i+I+���T���Yk�i��vm-��3�q�uu6ۻ�^V���U��v��9fk�rm�[�Ej��/�,�M�Y5jt��)݆I[3��Jۇ/���h�g��Q���-Ť���+P�{��IHq�܅��6��n���͈e\zA�ػ3hqf[˷��6�e�Z-ؘ^C�t��,�{r�Aa��[O;tc(@���<�F��ռ�ةr�ʴ(��a�F+��"F�p��2�s��.�ͦ�a=�L�'�lM.�Xvs9Zt�y׼	�/$V��Ԁ���)}jY�u�zD��5j�T���^i�iW2�\��{7`��4B܋��7����51�~����|�W���P���O������?o�I`5�BI"A���X$)", cF�d�3F(�_^�VM3I>Wc�<�!���z�����bM iy��i	L2M%"H�2;�Ӯ��CE�	%y�lb���^��ך�Qb����a�Ds��LE0�\ѹ��D(��llkr��&,&'uȹp��%��F�n��b���F��<�$��;�I��RX���ab��%E;�$L�F���[���#Er�`��H\�-�ͼ�أ2���GwIS*$i!,̕�4���・��<�?:j;�w���}�<��N�nvۤd��hƌ�B�g��rl�[8�M;�����y5q�����n�nx�c�#�͸x�;��u���Lr�F6H��M�]��{y�u�Ĉ�W�H�Z�ۃ��ݸ�Jw�c���2Q���OC:����m����g�M�����jx�T�����Ae��Y���s�3ڹ�ݸ�t��b�^0�n5=�� Y|p��ðj��;w�Q�qs��x�3�/h���O�c)�l�{�r�f�r=k�0u����:�`�	;خ/�|�m�m�������u�ܛr3����u�ێ=�E��Ö�sɇ���m����q�V+a�X�+��7;�C���qg�5az��a�Y��ͮ��ۜ\�,��8&N:ه[p��n+���Y��\�%���ʇ"�v�-��w<�rv����v�'X�烐�V�y9˺��d�݀#����ҭ���<E��N-�!�9Ƭ�hz��^�]8n�P�6�֓�4d�1�b�[^_NK�!ٱ�銷q���YŎ��1�Y��r��Ǵ�Y���k�Gm���iy�n:���G-�Ge�7h���ۍlOg���9�b������"�U�7�v�6���/Z������9�uPlu��ln�r1�67GQ��q�ؒ�R���A�@����+[d��qn譭v�\g�\�[Z��T�.{�68���u�u���*nۦ��ss���^47��Wi��ۻl�J�l�gu��䍹vܼ�o/,"��\_2�z������ɹ�çO>m�tt���e�ȕe���Bmb�3ڑ�-h�v�����G즏��ݷ^۷<ۛ�E� �8x�]�Ŧ�8�Ep�s��4��DR��]�T�$����ͺ��z�d���WoF`�J�c�;.o]��#f�5q��1���1v�n�wb�mZ�����&(�v�N�m��͞��y�qh��m��V���]'\���/Qc<��nlf���@���wv`�>6�du�z�f ���\�u�FM�p<p�їn�c�>u�m����Ф;\��q�wLS�n���pcaY����N�[��p���Ų�u���l[p��䋓n�`l�笮1��"5���+��mqv.݃�{��6�f�	�;k�ٰkk95�a2x�z8�=y���j�瓂�ȡcn
���&���j*�B�]�n6����ג:���C>$5��^�������Pq�UD��_���n���w�[�$�9�MI5�9�tN�	jل՚����؜��I?{�� ����vVKc�D�s�O��ŠA<�ݙݳ����sѠjl��|I��|"��h�+f�M���wR&莂�	J����~έ��{X�6��.z��c��y���� ׽'I	?��޻���öX�N�I^����n�o'�����$$�ϡ4HL^x�A$���UopTK���K�$�'��:�iR"��h->:�Ē%�7w	�G>Y]ϙ��o���k}ܒI ����:��rΐ������R��,+���]C�����]E��ٶ�,K��͌�:��A�sG�_�(�YTN[�#=�sx��Bg�f�H$�K�M�ԓ�u8�&��`���X�zzH$�s��R���d�j�e��+������zѻ��oZ��X���,�̩�����DU;���66�]U;݊�X��~�����{LI�����^:�(I��ҫ���;�B}�{�}2I$��+��D��O>q��?��0{❣ş[�I���H���Z�K�.#O�������oF�.�]��x=�}D��?��"	y����J!�#2(��S4�y���ҽ�v�?Ʀ�$�I����h�U���J��r�?��'��ɨ�(ݶ���sG�$��9K�jj��f�R1����D�57ͺ��I?{��%k7�yWu��1��n�o~�\��JT�{c	��m��sɫ��a4b8GNz�AV�6��-�Ϟ�8A���x�� [���� ��'H �ꙃC�+��V��-�ٙ��?jR��TN����c ��w��l_E�I?h{|�d�$����BI'4W��@������2_��w1k�s|؄�s9�+�{�5ލV��zjX�f�˗��]��\���^�Z�&�*��:yo9b�BL�d�5�~����g�`�r��51�sB䖾�W��ꪬ���i 
�y��4I��:HJ/`7�f��]��,5�2�[�B]� W�Ͷ$�6N�~$����@�~�T+p�B��f,�H(�%Vf���w��Mh�^M�.����Һ�	!I�2M:Nn|H�>��{w�j���9�{݋�J����+ ��Ɵ�ֻ]���QE��D;f�.Uߟ�{�����q����y�h�D��s��$�x�猧�Gul��{��IG�7y$-��ڈA���~y�k�ho��/Y�+i+X����$�l��WĚ$ѯj��~&/W@j���Q]����5�.���N���I�kurl�I�A������[F�� �3�y�TI$���m�Ǳ�6�Y�^����.-�;G���H	���В@�j�$������Hs�/�jѝ<�S|��z\�����N���u�+5����ɬy��[,uy1\�Wyw���E��鷽<c��r�U�Te����~�n�H��f�]eRG.LB�3�bX�=��+���eԿV)p$��{�ܒ�$���$�G�{��h�ړ��^[]֔V9�hƮ@�l6d�çL���[�5�����nڞq��ɢ�*�
�y\nwH$H��k����2��g�zha��.��  V�������7c/,^]��M}� <�����BI �[�'�G�sX$��u�^8��=��:���}��l��ƽ��\� 9ӹ�(� ��{��ï۫���=ݠ B����x=ӹ��]=�H�c��ܷOگY���X��s�I&��d ���v�L����nkA���$��|�=Z��$R�YD�/��S��s1�}��~���$��z�${O6� ����(���w�d��q�6E&E�5�º���a��^���o^X�:�<�FL�8U�l!�|��v���p�f>���Ă<���ݛ���}WН�y�k���$�{3�I�tn� v��=�\����A�6�mA����5�KŶwv��\��z��j�q����7l��[���2�"���\�X�쬻u5�u�����<��n݃��Fø�CN ��G&�E�p8{v��1׃���+�֙�{'g$i�su�z��Rz7�\x�����I��n��	�ә�v�ct�ͶuoZ9�16=����'�Ǚ�f�m���k�\﫩ߩHG.O�
����{O���$�j���ID��7�F�̾�����fb���=��R&�����*&���f>�]���FkXNqL޵Հ���N�L������h �ڽ�a�'ܻ��w[;5\L$�����{��@���7�����z�ɇ	o=�;ٻ�|�t�f}F|�w���\eUTMY����p��ސy,溽�j��,�� }��{� ;�k(x��#��N$��~�.kSj�.��U��6|�l��$
���1JlVz�0�*��Ē{�sr�$�W=�cs��k{��3�<VP	dm�ߋ��o�˲/��+t�s����P�7H�v޳��ߟ���^S���;����V��oٵ���N繦J$aں#�q)��MO9�!$U���w�)���滮,^�~�k�[�7�|���3C>���ľE$��e����x��%�/j�7=��6�!�8k�]��K;��-{����3+�$��=󞺊I$�/=��Ik=˻�H*�����y�k�#��bM�LL�t��MY=��?Q$�c����X��m�s�@t����A�Mߵvt�k����r���t�H����vt�>Oc����I���Ӣ@��uS>��.�Io������P��J��vh��m ;Ǜ��k���׶�q&�����D�ɼ�2�I��O6���6��x�>�آ7%L�-��S�ln�s;����c*�(Y(�,��>�xp��+���/Q��Bh�*-䃢@>���~P��ѵ[Cu�����M~5���)�d$Sꬰ�;�Ι�Y[][c�V���T�~�w� �I�75%�G�L�*3�x��u�}�^ʧ�{�k���ԖB;50\�w3� {��2�ފ���Ь�o��}�
�\�����q�_��QjM*Y8�/��'P8�U���jK��-�׫fݶ�O2fh���S�:^��ĒEM~N���p�df��ƃI1�Yu�=��NyX���ʷ�/^�� �|;����%�>��������$���7L�߮�:�IIG+���s({;���;����Q,�75$��8����'���7�{�s�}­�v�w}�+lw��r@�k�ܻv�-ˎ��5��7v�r�۵�:������v.���ⵣ�{��x��t�b�$��t��W�2�iǞ�[� �5G�;��>�6zb�+�W襹�׻����M](���}�I'�}��[��D�yΒ|I�vzz�#��t��>��rH�M�i"w0/M�V��3}�� 	g�钖Nx�H�jno։({�����uo^������.!s5�=�#MC5 l��  ׹�d��)�� o	T<"�o-���0`�5�������9C	��w/��\c6U�X��R$��
��\�e���ukx⛲����&? �l��>���Ÿ��/0i�.ޒH�<�Bv�ݏ�2�j�$��#�~�۲J$i�sŁ�9=�GA��6�G/�j�|O��UȴFj}��s�W\������x������m]���r����Q �y��� �=��N��h��x�'����I9���aj��Dл!n�7�w	9&3��!毘�I�N���I|�o�n�L����Sa�{9�}�{����y��5:1	5D��ɲI$�n�ve�}.��~�O�I)�I$�{f���X�r�bwX����Ӽ�8��Oy�9�'�O����Āh��7Og�.�Lm���s7�	ՙ9\uZ�%�p\�w1,�p�f\��㾊��I���H �N����5�'��<�ìچivp�����h�S�����mҪ�������a��y�r6�ua+�L�Y��߽F�g\r�MI���ro��1��^7:��)s� 7;{N���O:��;n�����¤c���)���s���7�wˮ��Ht��XݶW���̺��c����mvq����]��Ӻ1�m%]+oQ.�B�	��N�-V�;�sɱ<�d�5dx4Cl�S�����Ԉ��^��cjAT�OS�}������Qs@��C�Y�^�aC�2�t�ѻ]��ۭ=�l��vzWQ�I8˧��{p���p4us��n�g�d��!���p]C���9k/u������P�I����d�$��n�5&��tʋ���~�!$��ӛ�u���̢M��v��z��}�A��gvf;ۮ��K�G>��&��D��<��5IQ��kV:�_\sbK�`��!J�&�������| s�sS�d��gw�k.�y�$�F|�"	$�m���b�X_���#��ozo~��黨���>�4bI$�����hI$����R��j�m��1�k]��$��x%�b��
W
���3x�� ߳�����E"|��{Tb�>.<�"W�E���3�&�|�ʡ��I�N�Q�%	TMխ�r����	��s��(m��gS���GV&����|�{�C�¹f׳>Z ~>m�@?w�t���ݾ��uG���@���T>�P]FY'�B�.k>9��%B�cŐ��u㡅c�,J��:ӈ]�1fj�#���	_3M���~Pf��*���9X��mWv1&�H�W+u#Vq_\��}�ȒM�|ղM{ϺI�'�d]����Nk`��-̞���[	JSF �7�� {ݱϡ$�Q8��^�<���g�>� ���{�'��cqK�f�>ǸAt*hd��$�&�l��^�Ѱ%Q&���"��½�x ��;��M��I]%B��Wy�=���	�Ɲ#~�������� .�_��D����I?Qc���Ә�/*e�U��@u*;����ՎIucO�	W�¯f��ԯcl�Ma�ʁ��.�p�+$j�
��|���I n��Bh��Ϲ�=����[��Q8ky�9���ګj���me��ɻ�I�S��	�cWSM{2�}��3` >F>{3� �2�K}�E�-�����& O�)'�B�.����шI%��N�I�U|�lX��Ư�3z��B�wcF��{6K��w��B�x�Au�nof0���e;�`+�K'�^��aa)Ż��Bq��N]A;nT�W�18f:�fhzC�]2����j9x�mva
���V*Ԝi�1L�Z��9R��*�Ɩ��X��ˤ���GX7��>�|���D 2����b���6�u���z�!eD����y�s�C�O���7f�L��L�W��6�S��p]m��&�Lɝuwy�Pƕ[Ά��%�J�t���,�wS�}��޽���w���J���p��tT�yZ�5�;7��2!Y��_E�K��7�Da˃9;�e:�f�����CEʼ�Or�Q�������]��G�hA�ve�[ݺ���)��ܩ�5����c��*ɏ}�˧X����ǖ12�vu�(ǆ��F���b�V���qh�a1���iy�n��g:�b����-t\�����Vt��)�gn�C7�$Xk1T����ֵ��d�K)��q��ّ�[P�"�F���uc�i�}�*�X.�mn2�⣤:�>{vi{���i�g�i���*�����)+\�SQ]�tS|�ꆤ<�|)C�1��
��sn=���H�yrYh\�9�;hR����s�9N�ڛ�9�n��`e��=#v��#\ު����A3}i]Y������Ľ��'j�
����b!��$N�N�᫭Hb�����/.�]5�3k�w|�vn�W"�uy13�z�k�p���4Z�8C�>��z+��f��]*/:)����M���q�3K��;N�|.O�ۖwy^�r�r��776K!,�4�1��b�s��h�JW�s�sE��k��7z���ӻs(nj�\����r��/.Y+�h�s�Mr�5s8���ɂ�y���st�ĥ��\��^�k�v���75��\S��A�Dcd�5y^�tcP]ݻ��k��������j�wQ�wMs;ݼכt�wy���lk��F�*�D�c\˻W7����y�9���{ފ�����E�c��Ș����M�k�H������x���-3UvQUKa��`z����Ӌzg��eh�߼�BI?Y�oĚ�I���$�����skr����I,8}o�I.)�G��y=�O��S�I!&�o��h�T�շ�Ǜ�B'���Wi���ӹ������խX��[�9�v^��5��h��-�}��v0�2+�R�x׽��=�yù�T �rwy1u��ŜA��wٞH7㹙A}�<��(HՊ��Κͬ�L�S;o7t҃�rz8�ę���$Iy�۶�/l�?M�{������t��Z��q���� O��:x��;�׭���}p��晴H����e���K���I�#���j�9;������絖�	_����	 �^��d�.�}���62u�SpY����u9���g+��2�U��4�����i8���F��S�\������
;v��x���;{��l�Ĕ{�fG��U�J�-�v�a��sز���=���\���P��h�~�ݺ$�h���xA$�ޝ$�Dխ����(�v���}�]�u�Y���!t��:ۨ���u^t$s���t���F���F���/ƞ�V<I����[�I;�ѹTO,�d��yOsX�����}T��썑_�^c56O�4M�$�)�t�]�I��q~V�$��I!&��zϯ�9��p���Z3���;������>���OĚ'g�MȒ�[�X�G�3ٔ`{���������FWm�����<܍/����3�I*���(%ϧn�� �ܧh�R=�/�}'�eqA���O����G��쐀h�C�a�`~T��ٸ�l��$�&l�$�Oē�z7��خ��
�2uk�C�j�j����q쨨��k���^.���@s�X�X���3q�X#:�ᝩӻ��NZ�`� ֹ�ዏs��`ES�B:K%��<�^�9^GG[��n@&x�[�%j�4<�����:��7]�7.9�ܘ��<0I=V�6�6�z�;rм�-�y���T����Ƹ㱛v�t�����x��R�Mړ�vG8z_F��'����ݜe!-�j�Q�yC��v�R����vr\�ڶ����h��9����Kc�nÇ��0y���1����g�:�ؽTN�� }��P:-�|�֓�\�-uӭ�����oȸ�H�n��i�g�D w����@/ntv�y�=��Vn*ٜ_�F� ͝$�
q>���_�Ϗa�fPA�w/�h�m�/L�u$$�wq<�^�;tE$��+��ח���������NG~�[��{[��� ��;�b��i9�z0�a[��Q&�;Ӥ�BG���(-���mlv(T�g�:o~�-��ԭ㨹�(����I&�>��ۢ�Iz-�J5��t��A�w����T�B�-���/�g��g�l�/�]�c�U{̟���I$g)�M� �L�GNQo[ߍs�b�qK�ľf�ڎ�g��I�o�C�Y�q\��P�5n����L\^�O���׎�;��`�=�xMI>�\��%������NL�w{���f*s2����)!h�'�w��}��;'�Jy�k7�$q�\ Yyo1��\ؐG�Q���w]�9�;m�1��WG�Jܱ���b�U�/	yί,we��ޱZ.C��b\���2��ml }������̴I�S|#�@��ݏ�@\�	�H(���}ɭq(	 ��̢ 4��w����dbYٽ����:�	#�y����ON�9U�nb5�w�;�-�^^@ c�O�$�I�|ݿ�?kޓ��;{�5w�3g̖@�d�}�+�����b�N�gMf��~�����}�q�/xR���~I$�M�n�PK�{=�}����0@�6�T�\tڷ�S<c�\/����6-Q��9*��_�ajָ�s��B����<wZ����{3(���};�-����a9�;��j<�bK����*F���2����]k��;���g����Vyމ�C����/rw2`6/{������j�;��=��C��Բ� ��L0/Ow�$ w��s� ����B����.���J���Ic�]����+v̋2�iu�i\��N�g�[x�lM���jV;n�$��Xpix-R[;+f��/�Wğ�׷4Z+������$�"P4*�-����(�i��MQ$�x�oI��>��I/��d���=���Y;_�Gs1P����#r;r�k�ѱ���^����xo�,�/nʢO�[�`�7�k�C�\���2�����������vZ*��lhm7��|��ٹ�`6���v�b;Svs{oY�����߾�1<������(��s~����>�Mw&=v]E�/M���h�]�:I�4��z;$,���g�4k��P@��ܘo�Drm< �����$�E��o${o�U�oY �[�����L�"��$5l��	$⼬:$��hw��-��$�'��$$�j��\�Z�vY���-T�W�w�Qo�uI�;ծ�V���=����Y6�$K�Ϧ�_�]��Q�^�JWv]!�\SGk<;�p>�'Ez���_'{�Z@��5 �dɣ��5���q4}����f�V|z�|�Ï\�%cސ	����qF'�����T :��Ś{"���'�KւHt{;�'��,���t{�h����B%L� X�~tE�p����8�щ�E��r������V[YV4�}����Tn�5w�y��I�����$�k�v�*���M���;� #<k�-���>-,eE����p��ؽ땑X�v�d����I ��  G���hbAƸ˥������z[4uR+dd��&|sF���$�	lSR�$�!c��n�?9���UK{�� ��f*3����BB}S$���4�y�ǵyt��{R`w=�=�j��I�}~n�'�O�����v��s���e���Z�{�g5b���[��Q9��t�I�l�*��Q�d�K�����$�^��E���;�|_cd{9�Zk��5Q��'Alf�\��ﰌ�$i�^�v�]/p;Z[�d�k/����u�Í���n�{�I����3,k�������}-���#�I �O]�T]�^�{
�S��
�0��:�G8F3m�	�g��������=���l�Lt�v��ݺ�m��u��z��ڑ3�%����pRe�n1��-�%��6�O���q��G>k��8÷���n�Ce���g^�5ڵ�� �rH%�qˮq��ç��[am۷v��"U��T��r�c�u8�zۊ�;���;(�����.��7;7�,=�۹���v#��:�iV��:���1A����׎�g�7ޜ�<4I$��l�!;q
�ix�;N�k;ַ��;㹙���}�24���-�\��KS��~��sV��I$HI|ݲM�l��'�}�����Ĕ��|꠶��\���2��i��o>��9 �Kk.��!����uI ���b�������٣ʒ�6J��l�+�Ih��˳I�P�^:�<A$C��wpI|�[�o�.q3�*^<�4gs(8ޛ� 4Ed.i�[9�$�D����{DŇ*�4���I��y��'�$?+����}�!���q�8�ݻLv;)�r1ι���.a|�Ed��y6��g*clp�;�x�Z0vIeGg���U����rĚ~Ý��1y~9�^�W�!�����xL�RLQ�Hݐ�Vy��I*�$0��8U�i�[�*�2�����jֱ�^K;n��T�s�oVu.{|\�¦����-�~������MR��lN{4�҉��y��Y��ǅ<����I�Ӹ�Nz�d�	5��wR�}�,�2g*�����THʣ-�$_k����y�v� ��Nӓ��sH���� �������q��j+�ϋP���3��3vs���?J� B@�&�U�4�y0�$���Ǘ^r;*�qf8���$%�GU��%L�-��� ߏf��M�~mxV�$�5��BMQ!��'� H�;�����fl�ݹ������1]��X��sGhN�]Z���-ź�����`c�x�[��/t��o��� �k�X���s&#��y�Ն��������n��gMRZ RJeo�s�ܭ�<י��yq�8�n�}�@ ����� s�s1Q��=��ܻ����&	��%$���ug��tH�����I&å�Zy�œf���X;Q5{��u�{z���� 0���b��qv�%��f����y�,ʎ ���w.{$޴�o���buZ1���w_Oy$Al���s�x�f}Amr�t�O�cE����I�ThHw D��ȇD�g���ğ{gH����������տ�T���;�7���{��s-��\r�ں��D_Ě��<�$�h��6��H{ϧw%�7�qњ��/�viŹ��^.ɍ"� �����Fu&3��f�9�w��?yRZD�S.瑽j{3� �6��{gI>'�}���BGc�ܞ;�N�(1 �x�f*E��F �a��?������Ո=�����x�~[I�I�Sv�В��N�	<��͒�9��IF�R##sǻ߲� ����$@%���/��>n��p��ff�|�7���曽L(�akFa�rf8��e�;���#�=��$@F�wp	 �]쩵��3ֹ�n�9~�0D�9C�můF����Wu�Լ���������r-�����=��=���Ǘ����A�~�F��{F�5��<�7��W+�H��#,h�o��F%Q$���?��<2���Q({yc�O�L��$�h�+�B���lSK^uxzN48A��T��V��n���V�O#�d�8�9��eR�+\*qys����*Brz�ю:h�h��9�I �\�	�[[��Z�������$�z@ T��uv�V
��OM�h��`��O`��.��=:�PK�}7{�K��n���ܝ&��k�D��@zðI"�.k5�s���|�׵�� =�D0{���;���K乾��%.�ɺ(.kf�����L����M�w[����H��9	$6�;d�I��n�5{xD�7cp��R�OU��N`���x�o	�O���m���3m-Un ��=$�M'���	&��so�]T0���+ż�3�W'.+jWl�CsS؈=�ɱ�&\�ԥԘ�v�;��w4;��]��by��j=�}����an�ydt�1 ft���γ�4*%��%�}�#�^����=���ۣ[����5�R��6�:v�8Wm�����h/Mg,.I`��]��S�s�n�r�5}on�7���Ê���UR�-n�=O���vtn�g^Ձc �������L�^g<���^e��m�_L�2йl�[Fr�ͥ3B�jj-=�j�|r�\���ܬ�+F�X�۸��W���x$���N������F��*Cw�ƺ�[�R��a;�}�g��{�*�J��Ƅ,���;EM.wQ�r���׵u���4ʜ&���e�/�H��)ᦂQ�e��H�w[���*����=i��j����z�hSe٧�΃��`�)��X͘R�V�3��}tJ���#�xn�w�A��7E�8t�	��,�y:ͫ��y`�}u��>9�����!*�aٻ%K��̬Tcn	yUE��g��T)�o�͞��q���dۜ;�!]���0�)2v�	@H�X�/]V��X��9��ʪ���.�_H�-�)����m�l;�FY˒�w���(<��FW&qc�j'�/m���8� O������Ҩ�s��u֡�hN��y/w~�|J�nVu�0[�F��l��G�r�4$B���H]��K��!����+�nV)��WJ!����5���v�����T�n�-�u$�k���<�7hr'Z}���'��V^d}5v<4�~1�Z��-rѸnF���D\㝱t�s��X�9Gws�9h�Eͷ5�:��E̛���Qs�)(�����̹s�¢q���]��"68s�������:sWdDS#�#N��AnniB��+��s���M�]�k�nr�u�2������W5˛�']�r۴��a��u��1dws��鹸E˲�]�#35ˌ�P&��w(wn���k�.Qbܹ��Q�:�.t����7.m�����q�� MDY��K�4m����nw]]�����bAwu��a4�C����dZU����A;=[.�'�o[��R*��CcΌm��h���p�\�q�����-�iI�|�+�Ux:�o;xy��b�Ķ����0�|��<A���V�����c��N�q�vSh r�z'��q�Tt]F7�x�*V�v�2]��e;m�]���.EW�+��V�\�a��˶��vgs��4㧎���p��m�vq��1���nmݶK;[�OZ�[�&�y�8ܸݽ��n:y�٧�u�壛y��.u��3=$��5���ݖŲ.���M��7.-�2`	�ۘ�ε�vaj�Z���w|���y��N�ŕݻ��G;q�#�������i����f��l�����bON�w	ۇ��euٲI�n��{!�C�͂�{q�oPkqq]<����c��vǫu�G;l;�v�>v���]o<s�.��=N75�竜srV�Wc�8�xr�Oi;]��qr�܋�k����G6Gs�v�p�u��)�;r=��]�xNv�'dڞ!�����6�A&ݗ �֢���n����64h�nػbR|c��c���ѫ��v��S� �㚇�Ө��k.N���d��yÌnѻZ��ϙ��rt�m�9��0�l��xw�x�殶�p���LX������tq�6���͓t���b�i�ob�2W��s���n��.��v�����>��n�����eys�q����|n
i'W\�O�������緮y��Ʋ/\���HcA�ED
�Q(DB����#������ê�2�u�ԗ�ںy�e�u�s�ݺon]l�����]�nn:yޭ8�}���gv���Tݸ^;O�Ʊ;�=k�p��r�7X�n��:�{t��Oź��r:VV����ɸ^K���v売�rp8xX��no��[գ�=�箓����V�D{l�7��n��jَ��������R�ʗ
�s���^E�z�̎�h����,N�`ǚ#�Q�'#<�V��5i�mȱ�$�v�%\;\h5�Z�"7j���7A7Gk���K������ϲ\�ls��紉p��utS�sV:�����5;Fts�:�KF�:.qed]�u��a۶���V��7��痶'Y�v.�fڐ�o1��b;t�F�l�Ѻ} ��6��6���;<�&�v�X[R��:�xo\q�&�{�,!tv����5�6�v�>��(�1����H��M��S�06�`�t�ǋ�I�����E�;[�֖߽��?=������N�w3�H�3�\� 2O�}��%P�ݿm�;==���@?��*R�.}%c,U�ă��x�4M�{���W�����$��r�D�M�� 
�׍�b||�{Ͼ$�U��6JZ��˓h�s( oo���I��Jm��=�䵋�I4f����A~�f}�ME��0��.k{��.�0���D�'ٿZA$�i��В	�Γ��w���۬�}�sa5zRV�;-"�0+ﻙ��{��skf��~1��u{v���H����($��};�,YW%j�L�Z�!

���]jd�ƺx��Y�a�3�Z���IP��~���+Z�}]G����֦��p�f* |}�j�ȓ�'�����%,����+�k�8���|�fh��>�Q��~-�=�wr}P�����̫Az�.�j�t��\��Y��<;-���3�_�a�S��MRj�mC3�Y`�H
�8���%�$�i���I$�{gH����&�q�F���^V��"�X�#��>hTL��9��{��s�6��3-SL�Oē��m� ���'�֖��)+S.�$sZ��o���R�h�0zk���&�=���Q$�Fy_;j��'s9����oY�MES�R�7��4��ތJ$�3����d������}�/(��X�N��I*�4H�Wɯ�����J[b���V���N�y�:�i�)ў�n{�Ԣt�JUE+�ص��N�*q��H�g��{س@=�󹵱�Ϸ�^�uD�
�>�Άb_��" ?M��O���UGc!�Z��^9�h磼W�a�o�ѢO�I�7��D��4g����O����f�`c 魣*_}�WDB�>9����T&��&����%G��;I}���"΅=�1	����5qN�����9^��*Q
��ԧ�ڽ�YƱ�����U���l|�)Г�^ʝ~�l$L|���G������mH�
*8\o�ܼ����sG���� ���o���5옂I?7�Ҟ�yݗ�� >Jt����F�� �P�V΢�� `�7MKTd���#}��3��MW��I(�H�+�Q�����h���n/9�P�vE�!M�<'B�-�<�Vn�r��/UuA�787nո��cG�rՊPVi\�,��p�'�W��I$þo>�^�̼������=����~5�g�ޖvUeN4Ya����͢K^�׮n��;]���B�MM���Q 0o�h�+��dx�Z��6����V��	 �kS�&�> ���k'�h��`���rώ'�j�&yOf}�m�ٙ��kw�̉���[����]�n�\��5��a&����쒐I�7l�I	�s�F��W��o&������/P�WCOR�����4EfeMԐ��s��uyF�#�Zu�RZ��5��%#ѫ0Y�m�طJ>	/��{3�mX��܊��a�=ky��6����×���L0o��K�뚉'@L�n�:��9��V���렼:"�1�6��j]�V��K���|1kt�L�[�3r���N�~��L�Z2������b��H{ʹ����n��ʏA��o\�����b��ZO�J�#ep�O�7����2����b	3/ȍ$�H=����$����$���_�deI���zi�4Y\�e�W�K��7��JK˥�06��ڸo�����$�{w~�W�!=�wpI=]�Q2֦;�Mi\͙L��������$���]�}$���&��u�HL_%���H]��f][�^r7F�1���I	$	��:�=b���ܽ���xd��$zw�tI��[�$��	�W��Vlb���g�a�� ��^0�d[��qu��D����~�s+�޺W���y߱L�N(�c��G��ž�C�Y��q|]�`�\��Ğ��V��J+�X�TMz�4�92&�;g[���It猰�^E��∖��:9�GO/;=��.�ۋ6u�ɭ�.���whJsm���X��y{tݶ\���Ϋ�z��:,�g��x۝���Z15�]��ٮD��U�������9���G[>�%�m�Q��q�y�wd�^�Gr�����X.>Nz7�ƴ�nw;h	N�
���X�%ڻu�hn�;�S�s۾Z� |\󟛏X.�{q�h�g\nQ:3P��qR'{���7IZ��$.� ^��K0�&��{�! �I�Y̿���S�ۮ����,�]�s����Շ�NK,E���l�+�@��u�R��nc�g�IK�5���I|���7i|n�X-�e���(X3mX��e+�ߖ{��I-��v����Gn�o�����o~ ;��ٛ@ {��>�����D��W(V�4g�u��,���'�I-����Cf�5였 ��1�9���X��w$���J��ȭ�y=��$��n�����'�e�0�qM�|I$�g�����&���Ȯ�f`��?/ϵ�n��v��j 2��g�ŵ����Ԟ1�v7e��pp���.w�쐃#�n��S~�I&��W'�L汓�m=�VT�}����O$y���ӳC�m*m�n�&O���0yb�CZ\|d]ݑ�3/�w���^Y�xE��n��k��d�1ʧ۽�(�e9u2�D775�}�-�Br�0�;F�2^�+��U���X��˅�L�����H$�C��v��?7ʹA�}��s6U����IՇ�n[h�*����o��4I?�j����-�hD�8�n���=�ϴ8�O�J��
�=y�7=��������h���z'��~$����2I'��M��K4��a���fg�>ޖ�4�Y-�E2�A_}��~$zo9U�dڑ�xgi'�9�D�G���H�D��M�%��{�pM�<�Ŧ�Q�#v|�RdM�$�����ʉ���3m��>�-v�$rʳ��w��D�Z�}Ӭ�|_%��n/�K����w$�=��5�}��~�4�2�s3�1 �>{2�����@��/ź������=���m_t�:���Ԟ��% ���f\ �|���>Y���.mBn7�Ps�[�M���'�Q��$�=7��N}�3�5��Eў�̈c�lGj���x�j��U��������u�iW�*$5U^���Z��mHq/{�����x2� �S�®��9��7�4A$���w�����7,��ʂ�ĉy;�mB���4Osh�I3Ӻ@ �������W����~�|�zn��&�YaPD�ό����` {�=��\}L�eޫ���'JQ�@5=;��D��̝���nI�5}�m��(�ۂݵ����b��g� �1��&�jy�y�Xd�sε��|��+#D�Bv�+�{�� ��޹�>ל�����=�����|x{���0�~�����'�ܬ��6Z��G�[n���Zύ�U�&fq$���s`jH;)�E%�
÷`�^�cS+��p�F��gǵ��{�`�A�d��&���S�$9���j[D�L�����@|{�;�r�=h�֧l$.bBnr^}-ߪ��ޏ!В	U���I%�'��d�$T�5�;'�~fߒ_$�C��O=c���=���~�w��'��YIz���+��e״vU��^f�8��w'p�[��d��M����i��֥ۖ�B�bG.�px���1cyN�@y��z~$��[�BI&��}̃ B�=��I	8ތ9w�юX0t���S�|//Zlgq�z��
�s�xރh�Ŷ�_:߸��Q�9X^��s~��ߝ�;&��*o�L�kYU}�Z��=�fo3��F���Ϡ}�'��edr�82j����*�ӭ�u�O{{S�Գ;�� ����0 ��fb���������u����e�\wݚ�>������ �y�����y� �n{3�1 ����i��[W��p����t|�I\��u`�����X��Ir_'dTI�7�N�$��t��z��v������NM�O'~�;a!t��ӟ6h�O��9]{��!Y~{Lc�U�x�uD��&��m ��t�!#�#�\��7���9���
���V�؇2�f�J�a���Z+�^z:��x��~�Ϊ��ֺݝ��3=�.u=zXW���﩮]Y�8����Y�/m�5��)snN�'O%��$��1Si̢m��k��1��8��u�ϟWk]��08�%�/fJ���̝m���ںN/`n՜u���]��՞��ӤA;f���{v�V!Ʈ9�c��$=�����l6�y�!磢e�}�q��M��NMnJ�z�7���j�Tz��i���nuh��>p;��N�ضw�r�����n^`�몝�����n׮wN�s
v�=���t�nQ8]�9Rhq�S����ͅ��eaw?��'�$
��m�M{�:@���P�zo��ﬂH��4�4,t^e�t/8�^}͎�����ʞB��:ҿ.�h���@2O���$�@��6p�������P�B�
�{�)�s��TI�}���'�I.�%ft�m��-"H����$�=�w��IM��!-j�#^�\�w����\=; �Z���$���nI4g�c���{�f�k�ׯ�5�絋omޯ�" w��ϟI'�	��4Lޘ�4}�r�)*��&���tI�>�!$�g�c8��ʈ�Ͼ-&���$�XH\%�����-��D��"d
����EG���u;���	�|�7�0��3�ͭ�@طJ�:^�^��d {��$&��0�Y(W^��� �s�߈j?S���!�J3}trg�;E�۽6�n��/�j�78^f�{1��I��c�U�����_z��>V&et��j�+��w���	$���ӻ� ў鍒�b˭:e,N�?���TD�r���F{~���� ߽��$������j����I|�od��A~��7S3�P�K,r�L@���{]��d<��Ē^M�!4I$�މ� =��ע��C$���@%V�$�tlݛ �
����o�Mwtmߥw�%�pǚ��U��(��Ll�~���zv�(�o}�����G�U
�EѺ����c>P�ѮŎ�uC�v�#m�����	���im��A�TM�v��}��r_$O8� d�hOth	=<��z�{�$��=�ܺo�����֧,r3�]����2��kh���f��yt� �~��0`W޻�����w��t��ݵY(.�ˍ� ��oca=�x:z�O���W�>��Ϻ]uN�set��w���y91=�>
�;���^T;:�n�}R��+�n�>ב\W2ا�҆
��$��6@|6�o�t���Ι:�X�Ɋ{wuU�����}�jPǯ5>�������'�u���D#] �e^�#$#�n�Y���[�A]/gu
�}�>r�l�nv��@�񩬼Rg|{Yے��[�r"��DE��[�\����/s�:h�
N��h�u��a9S�N�˜��:��없[�u�`m�95��F��w79�Qŝ.,2�렫2u54��ڡ!���w`:im��I��%[,X�;sG;�Ǚ�#�V�-q�2�Y�J+�j�1���v�o�91USܓ`�w
î�����/d�T��ǵ��
W]�-櫋�Φ���=���{L%[!:V:wբmں�B�5{�/l�2��Nc0��{��Rww״tL��.��P�
���f�}��O�fu�)��
�(��86x�b��U��u6Fp�ʮq\�
3v^�kO1�ڪ\��|�{G)�'��ij�!R��yv�l�������u��{M�����[Uf�X��:�רd���5o\oX<�쉮�Zj�Rմ�����O�D����;��˽��r�m�Dmkt��l�,�p�×*�;����1�q�)�+2R+6**����c������f��aUٔ�ç�쬌�50k�F;����l鷵Q��3�g<5_%���1<�m�zOkܙ��s�tq��mGW�1We0�}��V�t$�晃����n0#Q�6A��H2��IRcF��n\����N]��٦(�Y]ɮi@�c��5�p��1sp�S"�gur�2%2�!���̠��w]&��w\��3t��릹�a�͒�.%4gwL�J��!������M�J��;�JQ"�
�nwm˚�tH��@QdJL�%��� �����:�K�e���.�.@b��k݉,9ȁ���,"E0Ж!9�\���E$��P�wC����wvl	�9Ҙ(�3��uq2#��.��
�܍"i1%�T���ThH0�wi&Fw]2�\���2�.v0� �uرr��I0HLR�I#�A��7wA���H������򲾻�$R<��n�x���`'ڌJ��NV4���s޻S/E͗NEN�0��)�w��K�H�nhI$��N��vܻv��7q��No̱HI\�W�>;���l�}�9���������k=`�"�z'� �;�ܢq��(�8�M/��ݡr�a9�+��6�����i��;���<n�Z��6�Y�V����HBFZ��ޮ���N�7RD��ӻ�Q�W˨q���ۺm�o��b��ӽ�Dn&����G�HI5��2w��q%=��I��$��&��:ITH�,w�%y瓾 ��G'S�Z�*p���sx� o~��ʄ�h�a�^��n��Q$�k���X0�w}���	�=!�Ӷ�%���n��X�*���i��I�:n��$�^r��})�r��b��v��ūX���[�����y4׹�j�)p)�P����7{rJæ�k��k1�������F�gx�5n\h�y\6�m+��̣�j�6|Ǔtj@ES�䨉����{���A�zsC!{1R�ϕ6�4���$�'�Ӥ��#������vN���[+�Q�����S�����	7U]�ޜ��U��铥ﯴ���!%p���;�b�> =�ﹴ� $�;y� .����v��y�� =��BMj��ٲn���1�1�I3˦6_w�+�c9�q$�K�>�h����@d�ǽ��U�g���������E"q4_��G���������I$�B�V����n�H$��G��  ��;9�[��E��S��B���$|�^v6L	>�{{�I��ޭ	�gӶnUp�>� �[띤��k������!7vUd�.LH�3Z�����,{��������oejܝ$�I&��Z "M=��E�9��']J�D��q��+'���9�w�׻.{+c��HH�go8���
lW��R����s&.o�^�o���KQ0Lq�v�]�+t�[5ڈ�����n��}�&�눠�8�%��1�-kq췶�ۭsbwC��̺۲�Dz�q��V��ý��urt�����q��e�y�4gݸ-��&^�#��X�S[ON�n��=���S���|w�M���i�g���{c�um�Zy�sGl'd^���CF�����N�Z:���k/=��pq�ݴ��Ns�l�ͧ��^���w\�莐|��P��E���]y9�KUD�5i+y�I������@$�-����H��P֮䥞���{߽�t�Ngb��Uk�& ��Κ4H����甩x���Oğ�?{�_I{b�}�<^̬�3Oj��ѝy��������� p펚4I'�nV�◩��ʺ}˶ �nkI߹�ϴom�>�Dn�Qϳ>���[��^�ܤ� ���~$���E�?��wkx�M�0�/�t[1 ��k_ ���<���S��A�:hTL�v��<�T�:U~^�AQ$�k�ѶA���{�d�������� ����Q��R���vZ�nN�aL�
Ʈlp�Wc]��do'}�~~�0t�mry�5� @���}�|��{�������#�7�v������M��o�C7E� ��i���D�8&�~�C�o�����9�-�x�r�"�N��H\�#����8܅�%���}�='Bj���x�y�j�ko��� ��oZo��y���}���p��9S��QHKS����z����*H@&v7Ր��DN��������K�q��Iq�F�*��֞-��^��:Q�� ��fa�s������w�]�O`��Z߻��3i�?Dn&��1��F'ā�^+0v�v�ԗ�p��3Y� ��{��� y�5��n��_=��q��Q6��m�)�( ��|�۬��<ѕ�ϳ8Y��g���������*����٬����=���~}̴J>�d/OE���4�|� �j{{d��{�M��*�T&|G�֕��OW���V��d�7��nI?ia(%��K��vo<�ϩ�'hm�D�j���5�{��� ~˯� �発�}��a4(�x+k;9g�q�qȝ���t�L�ŗ�I��u�Jڷ�5K_E>�D)ٚ��H��ٮ<���c`\���Q��$�I	}�A%���=}�'1r�@��m&�)����j~ў���@$����I%L�I$�����`h��s�MIs�I>W�q���$)u��5����16��r��j���6|��$��D�༬ ��m���*�j��w^+�t~�w�3�m��&���s�^�s�W\v�]�;����:A�-�[����DD�Uw^Fs3���_$�K�K�H���jBV����Y�~������u��ң��$�w�Uen:�5���Q9�����(o��6'ĒE�^�o@|.{���x�߸���*Hfs�@'��@���J�ra��P�	|��M�'R���3�x����`I��Q�s���A�-X����[^}'�X˖��u��KOz�I$�-�i� ���"T���=�I��wI��LgJi~=0N�R�:�YDط~>�V��7�Ґ��G�X���Z8�q��PL�7Y)QhV﫩K!�6�s��wZ�����
�e�����ıI.{�ʄ+���y�TI�J���u�H�D��{�I�+6N��=~���>뛑É��k����l���qЄ�Bͥ��u�-����*�>!w�F2B�W�G<kZ� :��ϳG�$Y�{���V�^G��E�fg֊	��8����I�"_��\�w{Ka�t���ה7먮��~��I/��v�$J�g����Wy�0u����߭u؜w0<�oi�{��c���w�ɿ����s3C Y�{��k������ڽ(g!�����}-��L�<'s�%�H�x$�H+>�����Z�����3�8ǖ!�9@��G��w{[���$���קy�ݙ��<�2I&M�j���E��J�ޟ	c�7��:�v�P�ǧn��%4�&^Ҧj������IK�Nt#����z;���{��)Z,堘��f��:� ��a=\�1�:7 ���ZI��=����97hڌ�%�8�mC]1��m�8���uvWp����d���x�jWYs�s���b'0����8� L���D�N��^(��vU�Y��Pc�l�;�9�9ۃ��m�q��v�û1�Y��z��P��/�^��tn��oO��K��mO���-�]-��Y�l��v:��mO���^5�g��O��:0����ի�mj��R��yz9[FJ�F��並	2{��'��H<3/�ʓ4����'�I>$���4���2Ƚм�fI|�tĿ{ڹ(���I+������	 ��b'Un�ȣ��<�ד���N r�u�׳���D�=��$�N-zquEA[^��@z�39��{�=����7�$�w�,N�6M_H���c]��mM�r�$�I{+ذ�ALz����m��0�A���}���S����J�2b&�" UDע��w�{��[�����o��I♔�$���~;�f8�0���O�"+T���P$��Sk:a�8�j\k�=�nY�(���
׳�οX��
Ü��ޞ�!$�'���D��#ܵ�K��W��x���>��0f�����#Q�҇����"�2Wt`/^w�{�	2/+&�s,�E��Z��mq�v�Y�;/ʑ�5
i{Ֆ�����xWD�r��3[`�Z�z�&���+pe٘0H�}�'{[25l�Y�׳�`�Gi� B�u�Ńo���'k�ں�*�r(���QUH�y����$
�Z��^`g�>u�P?��ڄ�m{��3>wkc�'��k~��=����&'�Ԯ��@�{&�7�������{�[3u6�߆��%����9t,b��� =��`Y��L_j��ff��S��(��������N�9���陙Ǵ�J�/�GG[gС����A�8M��Ν�Q5Yh��`���u��������C{� �?E��@}�|��/�VX�oה-����[hO��Ѣ�'ELDnN�2��{sV������dt�{t�	{f��I���'^^�2�����ꐌ���\��/;�m=�;� +;+dDgK�}��v�)�pj�Y@��.a��k+RǗ��Y��Ar�B���%�w��ʹ�>�f��5�4z�'S������:��:�ch��� �j�?l����ͪ������t(	����;��jGT�ysj��|8�D��G�w�4�{�i��7�qnDg��4Ho}��G�;	�yU]w���/'9#@�N�XJ�J�&�[��r���/�'"�V�MAo}�}��X�[����T�Ѥ�7�	>�͂���˾��h�}�n�O�WE]��t�=�@���V���OxO'�1@P����	'��N�@����a�B��b}�1��$�-����6�o��H`P�g��,���h-���w�*���B��Us>sם�Z�w����ռ���@�^"�&zc�}���C���Z�Y��;��4e+*�<{y8��J���u��5��#W|�i�K%�J����+F��f�Ƨ5܋�"W�������O=�],i���F��pD
�Z�gjF����<�
p�O�1��B�ѡ7{^/o}�2&}WT���Ӟ�g�ͨ�q�Nҷ-�	����۳q� )��Kt�.%@�4R���=�t�֥�I3��ƍ��b��%[�z4�ժ��xc0U��=�#u�>	4C�'��gA$��O���{��x9k�dyn��$@y��@��Wa*����X$��n�Ktl�&o��s�Y�~2l�?���h���,+($����tok^�a�7�`^G��	5�� �H��Ă~�<��hX]��Dp��z�?��'��
�I]�b�^����I �E�Ǽ�F�����PM�k`���:��!L�qx�W�6'-{3��ٞ�gqC��Ϸ5�od*�������U�{�r\������]o	�f��J����f����}�7�zj�P�c�;��N\���	������I9c�3�G�86�k%wtQ�A>���%,{D:2��6`h����ݻ���ʔ���%�����褪ڭ��fR�;��1�.��"�7��&q�-�LPS�J�4��PχY�M�n�z�&�D	�m�ڜ��O�h�qǲ���P[;lu��g����[��L��B�t�ʔ����ָ�"������]���ϩ<J�:���NΞg�ɔl�:�ƻ���e���z�C��T��I���+Fir,Z����<���9-�eӼ�y��W,������z�[h��+h>L-9��U�pY��e���z=|wX�$��6
�1�\E��U����x��W-��s-uЛ��6ح^��r�$mřz��m9E��H��;��͑�c>�pr��2ou��'�[5η�Juy*-�4��[{j��-��>���׮�)}k/�T��,pS�n��{�,�U)�IS�Ɛ�?��sI"���e����Uq�*�7�q�����je�z�B�U�3�	�e�R�H�vGz\��U�Ӯ-"cG�K�+n�����T���4y���j��S3%W��%��Pdf�=�F۶\�כ�"��ZkIm�*��*v���g^ӌ0V�r���f���i�;�J��Y»u���=��/��=��|_?_|ܾ��J��CA��lTlh���wWD�v� a�D(�r�F�I�#b���`�l�#\�Hܘ�$)&������DBM&�t �� ��L��@�	P�h��wt�Qݮi����e�,h�\�e�)�����2�422I�J6 �)wk�D�I�t�k�9���R��C�AJ��T��M�FH�Ƀ�1��M�2�&�7B���vP�$��;��6[�K����`���2��A #�t����u��(�U�#"N���J I�r%2̓RK(�L33D��Jr��0�bJ4awn�2F�1|�K�����u�m�{u�Td;u���ۮ�)lw5"�a�]�����l����Wv�J�݀���z�q`���9�p��U���0\I�	���0��9����j�j��;����ł�Iٚ�����^��S[h�s֎w]����Mc\k�Mԯnw�]�����On��N���L�g#icko<�ҝ۞�X��6�]q��u^�T��ݞ�t�G#9.�.5��=����4��ۊ�vL��wn��Y�rva�q۵<u͙d���W���v�Siy5��q^��n[���5�3�������I�n�3�:r�0����ѷb�*�H�@�K��Cp��/&�r�w]���M��Ŏ#s�q�c�����m�&�jwF���k�g74�v�,n{c1�^������ݯge+G�V��bvJ�8�:�Ŭ<u�i��rI����	J#n0d"vwk�)\���Sg�ut۝Ʒn�ы�v��;Q��C\Y�u���=g�Y��i:7]���+Cy��&��c='ON�ۖ)����U�z�y�9��f9ۃr��n��`Ń�t�����]s�G����-��h���^�ر�uR���Y���e����g���=�9���ȅ�hF�[`�c/(Wv�j��8��˶��v��^�;5��\8�d+��n�m����W>�p���+q��Ʊs�q��C;X�mZ�8�nu�kv�.qW�/�+cfǴ��<\�'f�y]ֹSZp��n���5�nT�Du\k��Ilbv�O/�k����ۊ�7V��*��L�\@`v���oa���yQw`7�rXJ��ps������n�k\yָ{��<�&�]�ō�O���v��[vz�����n;s�!��Cs;�<���L]��������M���+��^�Ɏ�]�<C�g�Q��s��7]n�m��z��njݫ�]��g�-�k��\2���O��n͓Qnm���ں�Fwny��=\Vq�����"':�E[=�;�m���3�1�G;g�w��1%�M�z�c4�V��SU�&�4͇[Gm��+�z'=�B�{v�E�6����귲�!7��NĜ�q�t��n��.M���[7=��uq�n.�n�6��g��eG�݄��7&ڎ
ٗ��Hڑ�`�\�'�f�P]��i���x���������*�4IpvV8:� �ٶ۬�Ϯ��s�D���˶�����Ĭ�E���2�Z��Q���H��W��C�|��@}�͆���S��}=@�v* oV�I	:<n��*7����2M�q���<����H��6��W��Gθu��GͿL����=+)kPU{�3cMg���c^�һ˫'7e&�_o�m���Wl�G�3��k~|�m�v���{%�xw����y7I$�N���h:NP��W��U癉�5ѭ&IXK���s�����}ן/��N嘼�I�>{������� �<Tr�΃�{_��/0�u���9�N8�z��m;N{q�
�Qc�����&�m�E���/)�T��3|�?�O7�f����0��n�Y4e9���{��OӜ�:�
�f�UUF��+��|F��Ne�^M�ׯ�',@��+�;�C�n��ޫ�pf���0`�r�Q��B`�'�l��Zi}���=A;�l�-L��M�IZ}�` +�sn����Pw��=Mu�w}������`��;�b�f=	.M���H5���֩C=rx~o��1?��e��w[$������+���/f�]���Hg����� ��R�P�~��B�_f)y�7`�����M���匊�f$�]6�O3��b�Yn�"�|	���~$�zL� �~��=���u�٩s��_I��Q��H�v�7[�Gk�]��u$"�e�;]LnEI�U_q��p~aB��Y��l��
��P ~�����C4�����]0(oye)WM�Ԅ[�Usd�;��]�]���s5�ɀ {|�/������:[:V���zf�˿z�"��$�����8��{�t�5�Z|���@�eڴ�~�.8�ͻ0�&�*�M��V>�i��s�bF�>Өzn�:�ȋ7U��~{���Y��Ov��C�ފT�ې�����$g{^�=��R%H�9�~S[7x�Æ|���) ��́@{�s�s�k��g����!~�����9��]eo��(
�rt=~'<�U���@|Զ=l
�:��oK�O.`B҄�:��J�j�I�9���f�iGm�,؊)`US�9/ծ���𘝱�Q���nA�f�$�H�웧�1�@��K�@�����"�|�D�Wg���':t`��A��׏�@P��?��{'7�7QayTdJ��L��n�Wd-��U5�Ns����ico*���G=�cw�#�� �|��U^�Nt�V7� ⵫��}g&�����q^q�}~٣H'�L����zVZ��о�f�xG�~�Ty�kv����(ίZ�ێ��p�WN缟;�݉m��/_7�ٛ�����<!�u��}D���<HT�۠���$�*�!_۷��F�AnV`G���#̫r��}{�F��[���zV`�^�.�uw�\�	.�6�v����m5d�@�����i-�箝�5�R��7{��rC�l+�����y�cm���h'���9��E�vqo[?U����y�ck���`������c����P��d}^���I�st3ҳ�k��ǵ��j������B$�T�ҫ�-뛿~$�/f}DvOy���_C{�П�r��$a���7CJ���X��
�9j�pǍr�$�r'@P��yZߞ�C�[0��@��n���X�A:���/���3f�.���9�7?o���$�|g�2����j����C�r�Kf`.�W)�4��R���m%��[Xy��l��o���H휵8s�2�n��/�,7�b�7cV]�Ǣ2/�:mP$1v�*�h���j�5P��4ʤSUǇr���[>�R9��]q���[��݇���cn y����`�!�^.��ZӨ�
�X�%�6=w�dwev�v�r����%��������j���Wo ��SvͶz��d�E�ݏl!�Se�wjg�Gu̷A�vss�$��X�=*���*��V��9��`�t.w'b-6Տg5��ɧ����v"���77�N��6#�#��S�&���}m�����sS�t�|4o%�P�����8�w[��=I��qcoϽ֪�ےT���\WI��7Lz.��s��A��w*�W��Z�G��=\���җ��P�=,��t3,]�"�/�� ��N��^v�����P <7�e
������({��$P�ViUמ���Ẅ}��I����^�\���:�X���}M?����X)��Uټ���/,6.��L�ɇ��-�����'_ ޞ\�	��kכ�Źɭ�����D��m�+j/o)�;x�b��ĜoVbջ��� ���U�����}����Q�/�}s�f�y�� N�M�x�}�����^�z���Q���	!&�� J�HW��^�~/��QH�ix�s�*';,���:W�C4YA���>۠�1Ee�긡�yv׍�X���6au�F�>��+�UR�p��o;V���7"S���d�@�z�I�w�n�H	=����a�z�B�~�8p����#�di��˕:/�|���,Ԯy/j~$=�4����7A�=ԴP���U�"�X<��}�yf�Ķot ���t(�\��}B�{��r��v�/J�&b�X���oKPb����=�?���j�.��i��E��C����7I$������w}��ͶЈ#�},+�F�9nW�;*h�U�gm���^.&rNۢnO��L�t���ݚV'�T�F�����H=��d�Ilg;��qy���#�͉���hСvE����y���{�/��R��פ�Gkɺ	�}3,���w�oہ����k}` �(���=o~$.fY$�M�X�U��W�<V�ې�*T��V����,� �ۼX�f^�k�M��R�P���*DL�W�����w��]�m��ym
]k��Ө�)^�L�v�(G#� �דq4���u��v���(�������z��*��t�A�q�������}��{z������s3�Y��H�,$ts0�7(�������$
�w�I��g�$g���mҵf%bSQ��n8C�{%��\)ǔH�
׷,.9�ɐ.(�W\vyn�cO��g�(�_+�o��6�~��`����i������&$����H-��)�8�]#WV.�c4�\�4-l�l�^�~s=䶀=��*�
{�=$ح�y�cݖk|��o�'�YvM"�hP�"���+x(���n��*���OH�����=�Bi�WB�^ݍ��&��@��>N��sn�yV.IV�^�I$~��A�ݛ���{����cfMx�c�c!��io)���9ى��K3"����4�
��n��Uk5�Xy�W�~f�<�Vc�j��I>"E邨�Uz��]���&�R���H=�قE�Y�mj������Ӡ>���YnI��<N�ҡw���%p\�h��\q8����\{��չS�촋s�8F����l��"d���ԇt}{ݿ|�P�|�Uu����9] �9�T�7��A@�����so[z|k}�����}����y�@^�|��X�����Jm.T��u�U�
���7���&�=$�%�/:�V�O�o�n�{vn�8c�Q=E!B������%���fm|מc���ovn�H�9Ϟ�f�U�/.m���5�X����v��~#���DY������6�]�]���r�cco�����vi��"�m����ܐ\�f�kh^Ņ���隐=�ԎnDx,�'u�h*�ѝz�U�y��ÂZ�����k..W�o�N�F�OPv2���T��h�!۞U���K�XƮh���]��^8��u	�6��pq�]��n�{�������^�q�S�4g-{k�ȇp�ܔwNC��볚A7P捴�2�
y'���������{f�u�St#�����xva��Ý���Ml%��#t��g��U7k�@u<�6{	����s�`�$潶��kFnk�n7��C�.s�m�u���r�<�ƞ�pt�ɡ�96y���Ao?���~SZI�B����4�H-��߉�	�\X}���|�u@P���
}H��l���;bv��i�禹�����yOr_M$�@����?g���{7�����q&���f8�]_f���mw��a �X�?OC��{! �7H'�/M}�=su��`f3��lvkGE���T$�^��߉'�O���,$��{�=X꘰�/�c�73<H��d�l��X�{�R��@P[9�⟁�0��j����3�/��
���{���S��\�ٍko����RIkR�ӑ7fG6�j���yxx
��_�EU%�����|���o�y�xI�;�A�ٻ���a�3��K�m=��Ҍ��l���e����;�oZ�i�k�*�[T�������.� �9��!P���wd���.�S�V�[��'�K1��5��{��x�\��@[לP }M�6�>x:��u�KL�P����y����H^�F�i�sًm������-z?h�����@�F�{w~�A�6RTi+4����yc��(�O4�����5���nծ�|��Ǩ
�j�}�=-�B�k��1��w4�~�s�Ϝ�+�o�G"��XI/d��~��7Oc{���t��O�Ԕ��� �]5v�;�ZI;'<������D-j��8PU�o�M��%D�vE����$�;��A �{���._�n�t�ub�_c��w�@��P���*꿶���`��۴2�蜐�� ����M����{7�ݻ�Oo���㒒����~��g�m����$�f֋��n����4�®�b���QD�ƩP��_:�Y;�i3�ˣ��B�q�ުtP�p����Q���,�D]ʸu��v"ꋽ���׋%b[��f����y�ϧ-�^��k�f-�C������	�o#�8�TV�4hι���W �K��k�Kws_I�}3i���Lu�uK���pW)2�m�&�N�SF�O�����ƥ9�p��v�I�r:,jT��K �P>|3M�w,�bOQM�f����&tp.��.On���O ��:z6Szނ+u�Sj�9cYwu�P�,�[�Z>Uq�T\����ia*�f_I�O�*Fa�7!W���tf�`�b�������6D�C��3V�����`[�t!W"(�DU�+�(݋��*z���n�lE�.u�N�s%ņs��;���ӓ.�m��y1u^�c[����Z����<{0;�����}����i�-Q��*��/N	L�.�T^W�:��c�l����u�������N��/n�Iv�|��t7W-�t
�3��͋�B ���c��xYל�i��*�g��<tyZ����,!�#��
����=5��h��K�y�;ws+�	�j����K1j�r�<�G����ƹ��9GL��,Eww�efε��i��H!���MzwB��X2�(1]r5;�ǫi�F���=�5�E��+#��	����80qo*��o\��F֩o�n�뼈}٥7�S���oIח/#3VP|%������33��[��D>�5�jn}KCcb1�����s
1&M&H�(R�uԢ$!d�1�n0��`�&)9�ݙI&;�]�k���$I��I�E$I&�s��v�	��,҄��[���Y� ��� 9�C��f	M	s$$�ݹ3)��d�M��J���t���K�@Cc3ΤQ� A	tX� ��&"6���K�]&���uی$3���RFf�';J7w).��j�k�H��$52YF��2U�]�u����K�L�C0e����s�Q��n�"�2�ݹ4�d�w]a���&c��d��2�lPc)�D�)) �H�"���286ƝL��>f}wcm��.��έ�RZ�ݏ3��5�lz�\�j���I?�9�h�\le��;�ަ�����m|>����1��/�?c$�g��+�=鐍��@Kٞ�$��y� ��9��??>o�Aka�ee`��ݭ]��;�Ɏ��<���sԊ�\q�p���O@zY�J�]�
���ܙ�߉/���G�U[��([h�f���)o���9�xb��:�TJdX�N�Mb��^��O�߼4�I!�stA~W2����_$=s=�.ۃµ���A&����ݿy��$ڹ��$��!�`�J�����h'��>~Ѡ�G��0�U�,�X:�'u��kr�/c܆�=�pL�~ɚ	<�b�A�}��{M�}�ĘӇv?'==���{�.Eh�&���x�1�򚄛�gr����ӥ���F�M�5(�x�������x$j��+2��lf5t�lo��[�@k/���\�s q����ؼU�S�}wM�Ky==���nZ�$N������K����@���n���}u������~�����Nk`P�|�X��ة�K�#�U�/�(��S���ug3]�cE?\�A䓒�
U�z����|{�̠�ة����@Ot7�y��I*%�/���A&t}�@.�ۗ3}��&� ;O��@S����n��M*G꿷~�c�­����o�q� h�U`
���
ޝ�L�y�1�HO������5P8/����Y�^st����ܑ���.1�;�hD�N�	���f�����NfB�����#�
�X�5B�B�ޫ�6#0t���3\�2�]��*�V,���j������Gdǎ��si�eһ5Z�֎$��ɻ8u;d�ڳ�m�·���l<���7c,�
%e;v��{/oh�ە��Huh�Ϲ��8�;�����w5km	n��cQS�^����:ئ璭�\nt�n�9�k%�ۢ�vˮy�^+���5�m���]{;�y�3���n�O	�8	�A�۠R`ҍ�&S�q��� %�p��}j^NOc	\�v�;7ncv����`�ݽ�8*�\v�\v��u�c6̻��5��L5Z缏y�K]����u�{_V����mР;=��P�����p�W���y�(uA l�FX�U�������8o$�4�����sI&_���g��N��FoTvq�4]٪��h�RA����٠�N��Խ}o��U�w>�t�[t�g�7@F/�P�h�.ȼ<f�g�׽�`�$��ۤ���t��Ag�=�S��;O�7��=�Oמ(�iR?U��o�th'���U�Ǳ��p+g�T��l *���n��,��u�y�߾S�	�5`��Q&�����q�Uׯ=&md�^z�7�$�U�g�����
�YIdw�=�fck����M��!�\�%�����7��̀�cΛ���"�-v'#�:�4���./W�{�uj����gw�T�w	�FGF�h�~xY�G�(�z��|��ε+��u�A�m�g��պ�Hm��Lxn�-�^`P���`CG�*��9]�+�Sʞ'@		X<��ѫǚ����ٖE ��P{d�=�<� �k�t��'-�E
�{S�~&�u��rǉ6��؟����ր�<�g���
�=������Ƈ$U"��<|� �����s��>��`��:t+��e ){7��OZ˧`����JrHAB1������uݳuӸ]]��{.PӰ�K��kn����w�� M#@U��ϳ<H�˹�@ �o=�=b�%��>�Ǽ� =�_`�^�T(V)e%��&s���|��Ś��j�u@	$׮V	�{�H=�s�*����hy(��G2�0eл	��+��>���� mwۺ�Q�ш��?�!�M����!�Ӊ��,��P��[���q�UPy��\�oN�p���eZ�Q=A��덕b���ۯ�Y���{���`�I���w~%"��RWW���~R�s�Y�� ���@y��ӡ�'�R%�R�����,/�̤a�.��e���
�W����O����{g���� >��m����6�x�����Z�Iʢr*6����	H��b�v�Al�nv���`x�\��7~����~8�77�|}�1/#�I>�N�]}.����yI���ow~9��ꯍ@]���r�����ގ�6�V��@�)���{�;t�I��k��X��"�&)ZF���]�@�M� ���СC=�w���~��$���n� �읺	L,�A]�]
9"��^��]�mY���w�6�;��I&L��	��,�_�,�s�AT(g��ާڪm(�g�o�2�2T{A���Z��;�.֙�r"�B�So0��.����gmf[��x2�;�������&
 *�J�;��� {�y_Z�d��Y���^��P�uz:߉ ��&}]Č�脺m�|�@}��zl����:�m���.�h��=�����.�&�)fbߧd+#�����3���X�{�� ]�\W��7~�N��s�oO#�s�	<��	�4�4:�T�^��Xv�������1�	��S�Wx���j��q�w�s�r(z��D�df�~��I�[Y0Q�k"��y����2�/42D�;~�g�L��ba&��H�9g�L��ťl�WS��6& w�x�����9�;@�����sZ�md�4��,��!#�N�]�O�9�}�����Q�5����y}t(9���8Rs%�u����Ʉ�2��x��o�8]��D�V�,:T�]���5����*��]t� Y�m�E�o+	�j��� ��p�Z���\�qu �[��';�t.[sf}�P���V�<�����㵣x�6��#�����3ѝz]��N����󷇣�_�㭌R�a����窸�n��8�b�<�k���碃�wV����ys��չ���]��\<�u���w�殥}��7��*G)��gcq��㎌mϖ7[��.��M�G=X]����;�hmێ��n.�x��W]���V=��Ba�W-��.ώC:��wd��B\=���綠���s�t�c�`��T���9�������@�5�By�ZM�!T�kn��/�2�vn9BQ��k�$�3��o���B÷�؁\�:>ܾ
��
���)_��	�<^�o&a�`�
�T�X��[�^ǻ�@%Qb�������'�װ ~${y���_�+ ��V��}�ff��9D6,ϻ	��&��r������s�sZju`�+��m�f��B��I��fg����>~;��ﱁO.2��z�:��|��Wa�o<���]E�uu�$���h�uI��� ���=�K���cuh�&3t���/���������:����~�;M{J}�޽��m���qg���ڙ�ד�NM��S|���`0z���]/k7��I��;�/ok��%���N5w��Fνue��.9�[%eS��j�ɀ�f��޳y
�̷�wm�x-a��,��G���/;�uIjw��	���M�	�׳F��%Ov�w��^��ǗO�vX�Gc%�1�g=�i$�^�4��$�Pݖ��^S� ���sP W���	}@e$�&�}��'��D�V����W�nh$��f�$_��Ow������S�w~'��L��d$vF��7���ڹ������/�=^�t?	/}�@$�+�V�m<.�,���F���������8�);FΎ^{lb�mF��%��UT>�|��ە�,]��~�7to��fi �?OUş�5鞘){�3[`P����΢����	$y��k��'�g���s{��������׾���A�W2��׌c�A=�Op޳�7�sCA$enY�o��$'��%�u2����󯓢���q�.
�ĳ��+��ځ��[��v)m�5sdѼ�
y��3z�#�3]�x�;�}��A~������s�/���UY*»��W����L<t�%�� E�`�H'�긳�A#=���~�>;Y�=8������r4��6I��+�Ǽ��?9�&m���,�W��'��^���s	�=��A0�3�'U}��#��,]bU��<j����:�
Ul�9^���&����Imz��ju�N%U|��y��	-��	=��A���3��.�}�o^������K��;ա�+ Uk��Co�LL��s��Kϳ�L�M7�0��c�����N���{������1�9S�G�!}��z����'�ߴ�n;�|<H�H$Es	=�w~��Ў�i�I����}�2mq���.�EwW<�N7�� �=�٬+�Y����
'��=�z�v���H<O����f�za/+�|f=�Qhj��U�ʾ���]�R9���X4[�`n��'K�ד4oZ�r��v�T�;m3>�s�� o���o��0*վ4�o�w~$~��7~3{B���r!�H,��0�+;��`�]�hwDn�uV:_nx�g2���x���_|�����!~�|��i(�2M�4�A?{���=��u٪z���Rm}�=7t3x�,! lwo�����fB�_*N��fI���}�st7�Գ������}�|��d
�v����wI �㙠���'2����牂Ig��O����#n���*�򁻰شWx���z�;ʀ�}04�I.c���'�W1��37;�0P��{y��
#jj6�%r�]}�g;����+�|+����je(u��H�g;�����+^$ I���%���m[��Z���ն�m��mj�~�m�[o�[kV����Z�ߥ[kV��U��m�歵�m���Z�ߊB�P$�	(�$ IXHE����Z�ߥ[kV��mj�~*I_�H@���IXH@���(+$�k9[z��|�K0
 ��d��D'|�  �    �     (       ( @     P     � ��
*�(  �E�@H  �J�*@ �T� T�(*�U �B�(
P����                                     �          z�+6�ؒ�f�*�J�e�һj�� �AU3�).l����wr�@�:�JY� s�ULڊ�,lT�%J��<  ���J��itԬ� Ԫ�l�L4��Qf�cV�r�tp 7:�����US�
�m��EK����B����KO  �        �CB�i^�R��D�ҮYT]ŕ*P� ��Z:Ԫ\���eW@C Ӏ �@PS����U�RJ*�)X   \��llP� ��P�]�U�hU��I��^`����8 ��6��t��(�`J��6(��Ҁ
   8         �
(خlUR�ses4���� F��� 42 ����d�
�B�Ix   ����4` @� ���#4  	  z�Td �j��W�  �         	��D0&@�  2 ��  �V  Hd�`
���[4<   `y uL��  �hQ� �Ð 6 ��NEr�0�iU]V��%����	 x  �        ���*�jv�es4�JY��Gf媔�� κ�\�]bJ�j�Z�q9tY�*Nٜ �)U�v�RU�)���@)�  ;���5Eq����U� �u��]ԬҮ�;֛jW��ƚ˛ )�� v�nX�jZnF�%Y��t˙�k�|5Oɦ�*J�2�E?�RU  4��M���@ت�%"��dd��T��i2�J�40�J6T�  jW,��h[z�D@`Vnг�����L�k� IL��g?�$ I5!���@�$��$ I?Ԅ��$d �@�-K�s�ؑv$��7w0�8��R�x�-����gl���##hA�~�z',)q�N�Ü-\��#�؋�.��<���T�M�u��V{s��;��u��:��',��G8����1�����B�D����o T�Ms7�~�B�uz��sˏ��p���� ;c�ԋ �Z�	au��z�8:=�ݑ(����̴�wL�ǣ@����.V��vۧ[���R��
'6w�dM蹣N�[��+�.�W��&�)d���7^1�5(1hɕ�	����gF�:���th�u��eƌ5���l0�S5���^�da�GRvk���sW'���o.L��u�x�X+rGS;��[���3��&2j�˚`�_,1��5�O��YwJ���x�)��(P��7F�9n�	�O=f>�'c��$�w"�3��I6�еAFZ'o��f��u�8!s�7����4w=�훮UyH5��W��b���ۗ�͜�Z �����l$�Ѝ��掖rcz�h`Û7��Ov�;;�C�Q�2Nc�p#���q�d�6r��WL�ј�e�I�Z0ɮ�]���ݲ�_oo\�z&���wJ���-禰B�<b��۶ב�{B�[�؆�go1�Wr�`4�Ntծs�$y����vl"q�=�I"AMT�' F7ێ�n�z��4�&pP�e�.�:K��2EA�=Kݴ,����oI��Y_�{��wiq>�q�DکA�y�·`�4G�U����E����"t{V��Ti7����cn��&#�lOx:L���)}�d�ל`f�Y;����j֛�� $���G�wq�i��Ț�d�ܫ�q��ƌ�9��9��2�8�Q�������lݗ9���5Q�U�H�:4�L�5��"�[�.p6�)H1Ƕ쎲4��绑W�w��hJ��H��)(}�˪���W�=��(	�twWF�V3�}�&�Ǐ��s�GR�"<k\]�zw4�nL["�?��_M'6rEBa�80V0�o�f˥vާ4�]�)�[���gr3v�n���s��n�{Db��v�v�a��$G��	g�ض2.-���5V��t'�1�?{r�����0�90p8��8#ƭ��A�m�l����W�2>�ڜ�{�l�ڙJ��/u7`g80J�;�Įρ�!��$�� 蒯&��Z�^=ϳh�#��:�;q�Q��;�l�9���[�u��i� �(+�sV3�� wE����J�&t�$���/��� =u��K��=F�y�=,�*(H&�%��ճ.����M_cV_	�c�3-�{y�Cy.S��J��Z�3\�S��'h�:���\)#�qYQ�����
���$��$z��r{+�U�od���`�dw;Gˇ{Du6u�@��QBH/%R���!*CDyE ܖ�pQ74/�6m�.��9������l�סMP�z������e�p��kL��I5���v��n1܌���٭7͕�r:N�<�@xh�����	�W�va=	�	e�,�2�r��S����<y���"Qn���dL�Ϋ��rĻǻbR��hbY#�tr��΂��(����j��`��s��}v��u�ϐ�q�w������e�
��@�M�ysGj�méұEyN2L��m��7	b\�6���ԉɲ��u9$m���9�� 6嬘�>��~'5��.;z���ԙjf��m;��R'�Ǩ,,�CZ�*��ͯ!�G+C.�]6�Ы�{�d�y��yn���7�u��-&wu� I������p�m|Q�����oE��Y��O���ʪj�ծ+����;�"�n�w���\^=���3���9)�\Z��eW�|�Ĕٻ"�)��!LD�٣���������:�C8�y��>]���ii���ssq\Ir����ۛf��C�mC�UY9w(dM��}�f>��9�DС���,E�4��n���v&�f�\���� ���X7���9bc��p\y�A໳�%�D�����.�4���\RN�����d�צ�k:I��u��1a�D�s��gb3w'Y#�i��o��,����G�.�˫w�{�ҽ=K�>3w)��d�S"�v�Ob?!0|@����S�^M�귚y��e��鳌+&ΰ����[� T�+�����i�-��KF4�1a�r�\U�^I2�rȬ�%v����8������=�\z&wuy0˛��B���{�O�-qS�ݛ��L3qU���k�ǀ��e�����Z�ö�oo"�g����Ů��gmބM'c��5b�H gQ�S�݂k��w��m=�p�f�< ��*�(��q��!�ջ���7;\����:����k]�qM��ˀU�j�d��[X�-���i9�m��D�v�9V���	&��Ӓ�p7�9:K\�F�г���j�� [�������+
�c[w
�p���uN�R������خ�'Ú�9��J��{�k���v-x���׹tx�jYF��-�9���lT�E�a}(V=�|(�gw_C���Nh@n-��:�q���%ٛ4b���c�e=uwݫ�)���@�x:I����*d�3T��b4 -D�)c8ђ>�@F�r��=���u�n��
�c<.՜ŵ��>MM�5;E7�����_ѣ��t)��r�}[��
�_Hu�^ԋa�s�dĻck��cXۜ�C�;�d[��>��h��w���"�ܢ���jǗ��=[d���՜��T����2�v���ǻ�=���4��'5�T���T�B��ͱf��e�ͣ]�0Ne��rT�X��6u3����upZ`|f�y7�GТ�b���m4l�:,��$8�Wr��P��w#�<s�v��Dr|�Fm�EsNj�[7�C����r;aڞq�ot����8s�h�;���!@�����_r�ǑI�w��0L�uQ
�,�gn�����~x�M�cF�C��]��$��#7iV���~�#���ٍ�yj�f��!ǆ�tBϙ�s���3{"�Ea��Y��h�;�i�tPi�#����-��h|N��]e�{�f�Y2� n��q�sz��8�Jw��&�X٣��մ���ĵJ��/��|.-R��y>�v{���K�L�z��g�аW��͘`sq��,y�ru������Q��#.:�BEF�hx�}5�S�إ��H�l�;JYo^�{͍��*���@\� s�wQ�p�&BU?�Xo\�ov�@��0�`������՝on��B&�����edH�%��m��n6F�"P���F]�UH����.�ְ s�8ۜ�������8��s]m�T��n�K�� Pjy�!�5��#Nժs'`��[�[4���N�f]=��C��i+H��6���� �A8t�i9�o7h����ٕ'��[�ySxl�j�5wk�l۫pHD����#�t%]гZvq��S�zb���ť��qgvVn(eD8N9d�|9
�a��w��ά�5u2���N�N�����Z���ᧇa�Kj���4�vB�{��k��p�;�Բ2H�_jm����k׹0d������$��@��7�'ۊf�qC:ٶ��J�<,iy	��-~�D��0�OGy�;���n;�`}1�Ý�#�ќ�g,散{p\y�.�t��k����Bc:.X�n����n���Vqn��Y����u��a&Nr']�t�2Os�N) ��KE��NnD���%�S��J�殤O��rk����ʫ�j�I]�'Z�ɇN�N�0��h[�-�6��-_k�("��R5C&��4k^��ZpņYq�"��1�Xj�2�WE'(g-��i��2A��%�v�sV�1�)���O=���<ɭ���KU/���鋳_v"�;�Æ@�!������x�E&\��B�=�ss�I�P�؞1�9��T�pށP�ߖ���&���s��%�gpYfHu\�&4�=5���P�FmN��Z�n�	��ȯ>����}z8vއr-ܞ)拊yyI�<U�9>]��#�ٴ�Gq���Y\q1�S��\�����"��HyiN��,��M|�[���H�П8cN)��F�0�v�)x�X_Q���t�8{v�����y��7u��;���5����u4K����c9���{�f�1���@a>�sh���[B1hz*wc��p��C���:�;E�-���p���Wjq��b�'f��Cݨ�i�C�nW�N�`�p�T���;�xg4P��)y_\7�������k_c�����\j8�):sf�
���L���Ζ$mڠ�[�	�.���_G�K���ӸSb����;���j�m]�U/:�nBlz1���*-�r&�_]��3J" 0I�p���1�*"��5N��{tUq�n*���S$Ys��W���3sr�i�����v���=j� �D��a�����۹R�RY�Ub�/�ܤ�Օ=�6-�H��.K��zb�8�M]v�+���I�鬤/m{�:��`Y"����e���LW J<A�\�#.��x��_QۡQܜ�����'�.���%��n̺qȞ��*���wX��.tU��Y6�U�<�m�q�dY{�:�չ�H��bܦ���0�F�Z�tB.9�	lŲK2�G����uc������-SuJ���L������p�b�w�O9���ѯ�1��M� ��s�e��z��t�h��N��]�'�`�O$o^E�u·f��viV�f��A�__n������' �ţ���mW�ތ>�r=��<`�I�gM	�v��u�3u5�8���NE�f�Ն*�*��kl�1Q�{�����s�Rê����������cە��wK�4������w ������i�oWoi�d�+�{�G9��eٻU���,jNbPDqm+Wp���Ɓ����88�,�n��M�ݻC�4q��n�ך�+߈Zzw�s���%'Sp��ݓ���d7�۝�i�9��{E���0Z^�M�ؖ��CMz�v��0h{$��ޯ���+GvDu$v�8�t�q�wv]�<)uL�5I�h7YH&�偅�t�è��΍���%��YT�ވ��!���]�nE��.혉oeޜ�ll�ź��Мl��ЊF��Bg���[˜����R��6�ɷ�s��[�gZ�}���h�܅�iȵG�bo
X5�.Á�Y�N�v�׏�ԣ�/D-�m��O�> K"�R�cx�ZJ/] 	<�핎�jq=`&�XW'O�	y�{en���쮫Ư��Pri�r��E^�:N,��N:���kݫ�n��ڂd�s<rwv��T{��^�/\�r�=xG�x��f� �;c6^�f	N�̬�a/!��D'�vW9XC��kD3�Eu�9�{CIN3��_37J���
̭l��(�tE�*�8F����77;)`|������N؛W�]ƪ�5�q��L��N\Xib8�8���N�9"Gm�nK !2��Q�p.�]=��s�NPP��&�̮��E�r{�٦PF147Ք���s�ݢ +���:.����o0�`�PxZ�Sg,�q�F�oC=��^��#�rf�,gV�V��J^��~�k�ć�G^�
�I������1���l7L}7e�E#r�Qn>�rn3Nf�� #MYʍݽQ�� �2l��B�j٧�]g(Á���s�f^�F��aaS�J���V��v���
����ˤ \��=�h��"5�}vT5�>��Z �>k�BG���D�:x4����B�Í�Ȣ�^��%�9����u�Տ:M��Q��qqY�c�3z`��&j�đ��'��Q��Y���֜��%*�IH��Ӌ]�'m�Yϫ�\�v������E�N.�0���4`Y�M[.ѵj��7����,��M���^$���92;�&�Z�i�$�8�[��d��Q�2�]�A�8�ʎ�d��)�&�ߑTp�����ki&lڱuS.�CX�*���A[r]9�)'��s��9�Ju��qQ��(]N�urN�Hŷ�.ϭi$Ɔ�
����)�͚t��Ԯ��3�8�@�X�(l�.��gt`�a�@����_a�O��qB[����N2K9�kx%�5sQ-te����Xpj:d�띵�(+���K�*���	/�Is��%�����|	���������B��;=���d!�M!�ifȓ�Nwwv���֎��UN>�P��E�Ց��3��r��n�:��FQ��%�*��:��.�#�E���ʰ�vr�8dvT��]���GN�ŝ���´���}�8wK�}ԒF�sbz�jx��9��%ge��t,�^P�2��Y�I�h�N|-�'A��Ø�����OO�չy��Μ�d�8�S,K9������ԡ��D�o~&-���XL��_�cB,��j���u;l��G�Rĭ[2h���j��+o1!���p>���%��J�v��r-��!NYl[����/�g��H����,�cN���j���SY7�خ�ߖ���p9v��@$:��a!R�H��
 �dX��HH� �
�H�IXd � @� ��H�%eIR�	�$� R@P!HAb�$�@X �!"��AaE��d�@�Y!$���	"�H�I ��B��
�J0�� T�����(�����	Y$�� (AAI! ��)!%BJ�$�aP"�T�d��@T��@ Y	� �$	P ��$*H��Y �Y�E!XI*@XP P`@H	T$��,��@$��IB %a ,� �!P�
"�E$��B!!*!RVB�$! ���$�	'z�����������۽�=�4-<<:<�W@�N��N�V�̞�]D�vo_-�^��1�1��崛���c%��^^Y��[��0��i!n���|yT7@���*ܞupj�����b�iKb�O.Α��&�v^vf��ճYE[��m��q�^�cM12�^z��ݼ����>����dqjK�ɾ��+g�^� �BOuyAƵd���"Zg,��j�v�ZEeOP���x]n�XM2y��oD��B�,�#aӞ�d2��K����<�0�O!XƘ���i˕_F���o|s��0����<VI�9B�򋵠12ټ�e��F��Ey÷�~wщ}�m೽���ˁ-h�2b\����b�8ER��h^��P.-�ؼ+��`7��<����xM��C�M��x�{,c�.��^�uM�K�o����w����ݱǦ����j�e�L�G�/�o.�z�k�?vY�`�2Fߞ]�����R�a�1�]ϱ��_d�Rx���q�m۠�E��;�.�x�B0�4�p�4x�{��(iI혶tW�yzI�N~���3��}��`Pq��w�=�U�6b�i�2�P�	��֥����d��)C*�P��ZK�u�u@Q�t�7W�;�r�3v�*�l�ٜ0Y��3F-�
|{��<O���n���!����0X�w)~�yj����ם��i�ɒR빺L�q\F�����sS�*�Z75azl�B�S�ќ��{:*ͯ7�������}ٻ=ݲ���:#=S�j�LK&b�O���Տk���7wg0�)��4�BN�w��o��u̕���˙n�x!��X�}�Ձ��z�l��˞�#<�;B Ǿ���B~u�ǻ|����[¬<3M���}���kF-\��5]�6w��'|My�{�����)�_z<����H�f·�����#��W�C�V�u[=���-�л�=��}���y���J���lU$�V"��˹��d2�/��2A�#{,�>�~�E����EO��y�Ҟ�v2��֗f�{fyI�t����QH���d2�ʐU�q�CO����JC>���ė�B�w=(wm=�{�Q�G�U����o3�cǵ����R��� '.��^�=s;�����oj��n%�P�[ˏW���Ň�i�\#�[oT�b���x�V�����7�Ѕ@��{�Fc7�@^�N�M���o�ׄ����_����;Wh	�q�!͚���ϼ�L�w�u�����3���N���x[4г^^U�z��]sɌ׭{.k+�1<�9rR�:i�]kQ��2�|2��5����<t�B1���pԴ�G��/��7=���#$��Ww�ok�ӵ�U`3r�b�^��H��%���X~���m�nG����P����n�w`�]��V_vhx�n���X"�v��uLa�����J=�[��0ɕ�#�Z"���ʞ�̧z*�؊�n����r�0j��z�n���w{���C�ǻK�������o��Rѻ�vg�R b�o	6j$2���9�[��1��}��1��^^�� �5�9�&����n��	tg=�.�ݬ�zu'�	ћ6Mמ�0dM�Ƀ6)������^U�bg6��m��o"�tkN�p�|��K�yr����$�K.o���ﻱw�8�Q������;����r�.;�fq�f�"�ظ���Ż���Wz�d�|�������]���N��|^i��9���vK�q��#V���]��j�L�Z���_���.�����+de���x빪I��*DwS���t����Ѻ��χ����O�7�$�׽���_g�N>(ܐ���#�};v�U�ʞ�U����;w˘�^�r)h;tz�jػO2��m���J��Щ��E������^�[l~�
�<hd�.�7�����OG-?o����,���v[D�V-]6��+�����U�M	�W�-�T�����M��̋L��R��vw���wm��vm:=�co���ti�9�<op�}���ŅOx7֠���9���#�M�K�֌�iGz����q�h�J{���+���e���Y�f�I�P���7<ǒ�����R�rd<v�ۇ�Ϙip�MwM>�p�~V#�9&w��#�&{_��f�A���\�.��O�G����5��+�>٫�&1�5���L�����q�����nD�GS������!���y��^<�.h9.��qUG�7_3����������o���Ů��'g+���r��=� r�5
��=���=��a٢�߮G�*Ų�����Wx�Eئ����\������}��=1���f��f�s�ɖ�[W<�����bͽ��p���k;�Ns�rQ箉�n��^�}��j�#���>!}�}�����O�<�zLߎ2�N���]��h�gb�w��R��Z��O�Cܝ�z��G��1Ķ�]��ӱ��;�qQ�"��cbo�A�Su��Y�o��X==��g��Uf�OfoF޾;��ze�Y=q��⚌�d����8o��x�2<G��wl�I���*����״Wή��W5�wk�=�W��X5�5c�;7uG^���M�zD�M��㾳��xf����~��%�M[)����Ţ�V͛�Z�� �פ.f�{+Z�׶-���3�T��U����1P����棐f�̞^�#�7N���Vީz�4�_{=��Fz�(hb��zcY};k�gg�>c��w3#-���/W�t�U�����9O�⩹�n��1�������y|n�k���I��bc(�t�K{+>~�����ǂ8�=`F����l��X��y�N�J�����L�r�6�i��sM{%�"��[I]���x2h��W�@������f�Fr|�T2���x1\�m��RX���He�H�ڻ1�ǎ���S��\��ox��-9��0�ڂLS��!7w�c �Ҵ�3ٓy��qw4=`�����ǚ��OjjK�;���R�%��m{�`'}1d�˫ط����LJQ݇~86xK��~x_�ލ��g��JÛy9��ag4{��h���������<=E���X}3��Ԟ�O�f)����Ï _���ܨ�2PNr�;��cH��x�wޤP�}�6ݣQm��5����р��Њ�	�QΗ�F>�&�c@�v=ׯ��K���d*��S�]��]Ž��γ\&����{Zd�/�S��Y�cC��`;�~�W��=<i�I|��S|��`�S����9I�x��z����)]3v0#.Ϡ�fnh�XEFȲF��>�:gf�عy�z��c����3�+���N�oz���8*���O!��Gn{<�~7#~�Y����On�����^e}<x��b�,9�wv�����w�ŉ��7���M�"���'��	�#����rm��TnYy ���O+Fꗥ[w�j[=O�m��x u^�)J�MR�21\��<ю�L�4du�->T�=ݫg��c�$0v��f3� eޏ���|�{z� �}us4�yۄw��ZW������CN�}O��n/b�eAO�ǋ�9ۡ�w����h�-���+��/uC�#��[7�{�N�è=Մ�tգ���y���S��Pv���G���u�,	�z_x�{���m��][���El�`�=�V�������Z&��Hu�"����;���7��|S�E���u.�.�x_�I�2<�X���ש�3ȼ�_{ؑ��������
���R$�̖V{�k[�歔����s^�� �����v�Ms�h�\��i���7Y�'��{Vs����&�d쐙�u�qѦg��@'mC��ຌ��O.�'�S��3�{�Ću���.՞�/ճҗ��o�%%�}�=��@�o�Ĭ ��@�.�CkL�[8�Q�zY��^:��]����㉽hg%���� �%�\�w)*�x���� _M��p���({ݭ�������\�{�G���Ϫ���f��I[�{��6�J[��R+*�ϧ��$�.,��|�hU�*��%]UM����� ����>c�iW`��3E0�¾����2��^G�z���e�XL�[|%W�ɹ�ssLd�9����pW=�»F-��B+/�s!z���d��P�5KŃ����V�.K�yb����76���\���4}��p~��.is|&쳱�o��3}2l���6����������fܚh�oc>^�2�PR���zM������2��GZ+��I~����w{ޫg]�;E��\�e�.�����En�8f���O��v�r�6�բG�we��� ����ظ�!��ws�KB0�>���,�`�~�PÀm����5Ūe�L24و{�3�b׮��vu�o��j\b�xv�پ��e��f1y{jд�;���Fv�r���v��G������5���Z���2���ѳ�����D������n��b2��'��;�E�X�]�g)��y��D��:�cܲYp�Vd�Mzv�3T��J���kך��h�H���[�gQq�7�8G1@%��l����oĴ^��ݱ�^&�i�m�=[=�s�����<P�2tG6�C��ǄdS��6h����z�(n=�������:���Gv�g�O�!pMʘo�	ˋ޵����T7h8���y����|�"����2���L�<&��I������]~r��r�;��\�s*�����D����pQ�ݽ#Yx.��6�ʍ���{E�;������>��!f���{[D�
3CY��2}hM�z8I����-W4VM׺r��]�;@�MNrz}Gd����.f��>${g8G��Zm�wo��ڏ��G;p�e��9��1]���*R�Oa�p�@�f�G5MW�9�l����p�>�ղ�A��j���<Œ(i��ڬ�>K��C�3D�[�-ju���G,e���mۛ�[ui����ݗ/C&�Q[�ݯ=u>���?A�B�>P7���x]{�}���7&垗T���ۆ��F᝾�C��.�����(�{N�Uo���I~�&M�'JG�b�٣�� w��t�Ŏ�?{F�t�A+�5L��<-��en��1�nD���������|�}��VK�S��������IH��o=�sM��A��hG1=�2����f��/y��H^ndb���kw�ˢc,>�����$A�O���o������1�!Ż.�|�.��-G\,����,�1�"��>�\s�������g��;io����L��4��[s_�u�<1��~~W4{��׈�Cg��r�v����nA��s�Ʃ�N���	���B �~��^r�"�[��rj�ŕ1	�"��C+Xa���a�ZtR�绻��Ob�ל~Z���n��P�G`���i���I̭�j��F1�$eW�B�K�e���f_eBY�!]��+�6ֽ�����nݾ��]p�}�����o�D�G���'y���T��ɞ��.��7鷞W9r~��lW��򯗃~>~����/W{ò/�V�)�U��GZ������ռp�=�ս��ޱyt�r�7G�o�1W��|��/R�]�2�N��sT�0û)�0�Ia��G�'�vt;���z��pʙ�{�����&�-xfۛ볋e�ס�UQ�}��ּ���9�;� ��[{��^V$&��Ys���c�`ʂR/Xa=�wPw���Foa��w���~Ӟ�,�^��:��[�N�fOU�}�az���}l�3�<�Ϳ�6�4'O�/@����ѥ��:�g� \�j�`T�s�-��d��p��_r�x�
��V�K��|o���^��$��g��J�yp�;��:���ވ#�ӵ��mXOGS���j���g�{����t�x{L���^��j��đ��cɱ7��D��Gc`dy��ֵd��=�j��-�iv�,{����ػx���-�?"��En�X2i^�5̫Z3�0�6��q�Sg��[E{���c������i��a:���U�O�{Fn�2����;
&���ޓ�{G���c�-����\����>��/� �k�ݴ�I����;��7��rQ��qy�s����ў���;�Ænl󨭧ӗb{�.;�=AF��"�>�n�_T�ׯ���$�,wx^�.{ջ_5y2���&�nQ�B��_��~Z�X+m?^�'�@������U����]��$T��^ �0�s���^�U��:�y{O/xl��~�]t������t�;�c��oX���ze^���\���:<xO+�����=��togv�'=��U3l��(��;5�M�NP��)�[�oД6Խ�Hi'��i��M�C��>�F�����oݼ�Nǀj������O����M���~4]�l���͈�-��^κ�)��`�z�=eگ�A�oc뻗�-~H��I�&�	w�����j�n��Q޸7Ny�����7ʝ�i^O��E�}4���U�o�]�j��_!yas<ȉ���٨��lt��n���|ι�h�N>�&�E��zH�G����1���<���{о�w	C �9�d��4c7�l;�f��*�u��V�gc{#@����=�>���;�!�yMݙ���^�F�>lX������#:�4x!uOUJ��>�y�����ef��)F=~#�.2t]�B��M͏)丁���W�u$����$:�C�M�N����6��g�4��SƂA��Z��|�;�l����Di'f�_Z�z{݀��n���G�x��i�g)�\}��o�^����lx�z�5YOB�/t�ť�����|>�;�����?}�[�����خ��cC��<]����-Gj�ϗy��Ǟ1��zWq�{n�����;��v-�7g���n�e+�J�Ֆ]<X4\�<y�6�sƧ'�=����7n��9Ay:M]���;/��g�ǲnÏ1�k��-�n��Q^%�[s	��s���{ekq��.�"�r���6��wFv����s�S�����*3�<�%ll��v�4�.���:�m�z�e3n��m�tzA�+gC��1
�ҕ��^�ٳ�����I�۱j�<v��ZsI��}�Z4�>5���{f�e�.ѧnژ��{k��A�!��۰���v�kkm�3w�;�o]�#: 8�^W���-M���+��lp
�=>`w\�6��h]@[���v�5�.-�&(j�ps�\�G/��,d��ħ��q�NVՙ�i}��m�H\�an#�V�f�˄�����Y鋜.���W<�v���gU۞n##ٍ��>�"�ĥ��li۝ҹ��Ml]ˋ��d���LF��۶yomϞ��vE�8�:=�u���w܁�g8s�i�f�cn5�����W�g]�0��ضΫp�붓W[�>qs��+����9�:�1��m�7��H���م9M�Y�a�S�}`�G���a��pձ��u�E�ۃ��;{��ŒÓY�ۜ�c��ʽ�Y�=���)�\U�r����l{>�l�=��	=�l����3��\�OFۓF:��u�4'��j�m�^ry2�Oj���m��ی.Ƭ�����u��hs�yc�ۤ�\O�6rJ{�y�k�l��f��;G=��;�ka;�h���f<ặ[�F��v����ms�9�����7$s��A��ѭ��gώg��=n�:��yݝ�Cܙ� ���������\>��ݞΈ�
���\�6�;7b�ױ��� /]���[!�N��9���8�X<�]vٮ�6��U��͜����k��3�h�F�%[�:8a�h��v��V�v����+q����1�`'�¼U�x�י�Uۇpt���cz��k�9�q;n;n�[��Zwc&csەSG<z�[�nw�s�vnvH���q��v�=�]�v���x�x��������S��o=�d�����<���8�M����j���,܇3���to���S�����>�/u�]���n=�fD��'>K��h�91lxB-j9^mۖ��9֒�=��;�5�8S9i�}��o;���W�s˒�$�ͩ��շ+m�R�!˝�Zw5���<Ҝ���=�N�s�ں�ggs-�Ѩ��:L���Լ����qٮN��캺�N��I(cA���-k.��w<��#��[qR�-�WnA��Ɖv���vϧ�Þ��x��.vX�;��箶Ƭ�;\���
qpO�o��T8g�nˍ�6�=��1��Ҹ��ݽ{�C���p���5��Z}9�lvn��c#�Q*Y��y��h�{p��vtkls�3qW�e����\N��9�*NϹ�!l�u�����sS���b�O�.]s���۱ͣ�Lv� �uC���i��է�,�N��X��+��@nm�k����cJ�`,��Oi�᳙��nI�*��ܘ��\��p�'8���<��:wP6���[�v@�:�4Wg8�;��v�vs�����	��U���]���2o>�!u�7�q�5v멻Gyr�\�.M���-�k/Q���Sӝ<.��;x��Z��Iq���=p�&�n8ld<�t�ՈW>�X�b{v��]��s��m��N�ջ;������,x��MuJu��9�ܖǙYj�0nf,��]]`�m�$Ƌ6{>��W�m����L�9���j���v�E�֌��빸ɱ�q�i�����q�h{ꊸ�経�ƌ���ïW�҆�nZ�s2���nKq�n��=;l0�U�օx�W�#�j��'rg"�K��g�E
��cu;n�:{O���m�ks�WO.�����v-�����D�S]�εr]<�����i�1����xn�۵�����H�(ǜ���q���Yo`l�[m�nJ�qF�ȫ1���x5vS/�t�1�s��gZq�����q��5{{'࢓��:��\�	:zz#f�
���\�
���nÛ�iW�ճͰi�{sŭ�1]�v�s��\\�&�w5�c�{����\��3�����Җ�<��W;��s�q>F�7.�$��ǔ!���t��#����m8���-�6�l󇔎Eǌ�z��gj�8���Ƹ޲��z���.2��aM�����z7�#�ݷV��"�j���lz�1��s�ő�s�=-tf}�S�x��[v��m��͍q]��Y��`.�΅F�pH<=]�����Ę=A���:�b�-�m�:yl���+<����u�`ݷl�kn�{��9��M�:�ĩ��Ku����)�]r�+�,����e6㰼vw��s��'�w]�S×M�%�w<�V���U^�tr��n�XYp0�p����a]���u�Cݷ�n����c)cQ�'VƎ��3��;���T�z�47��#��v�V�u��s�R�Y��Çۖph���B�Gem�mq�֟sga�<�mu���n����V�ֽ��3�ch�t�n�r;v���m-��^��۶*5�$(]�m�M����7 ֻq;�Fx�1�.�%�
c����`ԛC�c������0azm��\\���ͤ-]�N8�kb��=�����w:uƽۘ�Rt�:]�������*V��e�6iގ۷nq��ރ�Lչ�����Q�t���'l��\u���"v�۸bεۨ�:N@y�Wgkzg��s����n�U����qm۵�ϙێS�Wt�%��Q���Y�p5�>6���n�v����#��\�]<ڹ穬z�;Ѵ�m�\Q��Ok�g��=��s�N]�uY����u�v��g@횣�˒�=�=s�2r���w��袧1�c�J�n�cy�y���+F2�yn5[��Q��N����ݸ�Ga�/I[^x�V`�H�w=�Uz�k�� sy����7c�]��N��g'*^����𼗻%��mD����{	���m��)�,ll�ny^ݷ+����ܼ=qÉ�Qv����v��ݹ�bG�8�pkZ��Sb��G5�h�>s�v�wft��n�x�.$΍k��M�mv�g`6�/\;��E7S�"R�^q���K�\��<�h-t�.�ۯ����弲s�v:�6���h43����W�9�X���B��3��<��t�A��N�Y㰏n8��t�y����;{U�sC�;�>�1uWQ�t��m�7�3�ΠE��ֶZ,sݗ�7v�#p��N�hGƑ�U�wv���D���w	��T��zGqcv�먒)
��ݛ�ʝ���R)����G�����۵�:ǁ�-�*�[��	�\����g�Cg�����vψ������t�OMt�=tnڹ��[��tWD]����h蚕�Kq�ͩ�����:݋�y#p�5�Sh+q �M�vǨ�v��Þ��Kn�Bu�T��c��J*k�;�vˬ\�Eڂ��qq��tq�j/=��eB��'�-��ʃ�6��^�lN�����3۫�tnʼ/G��:�.+�c�tKy�շg��on�=��cg�*���<�c�rL��(������ܸ����ǌ<p�/��St]"'6m�u���=�˘V�W3���gYԥ�9�,$.ܚ�t���@���k����uy$�w�9U\ןGZ�`�9�L��"�]�K�ˀtst�1�r2�@ň�2`��^�(�=�A�-A!va��)&0m�\[h��ݥ�t�F�k�o<:2��v�ł��sH�\^th�C;�ۺ[��7��:�sJ���⮱�@7L���n1�YXU�.���(���qmz�;PPgr�y��;	�{#���z��#�۹@X���h�n�ccl��[�ֹ��3�aWVQ�\2����/f����2�H씙����%kt��Ʀٻr��&�4�#��m]�$F&�۳ϮnE%�g������i���i�s�qЋZ����Xˆ�Kع�]3s>�=v�GKb������^G�����l��q�K�3���s��,؇�o78Xq���S�n�-��ͥ�Z�{������ώ1�W�h�q��ns���`�t��<���d#��m�=�(�rsZ�3��#&n�;g�b7�E�u�V��z�4�c^1�%p�-\ۛk�<N�d�����f/��ݹ��ƶ9�b��fs��,����b�F����MG��̸\ո�s���}�ۅ���v�{m��ڗ������vvㆳ�.�m�nAwv=�f��<��+���rO�{<l��t�0,����zv���[�x��rmϡ���=�mӋ�
c�۪��V�P�ka[q��p��>�ۣۗ��	�q/E�RB�R�g5�rY����z���FW�֝�؉���v�mh����s���4,�sQ�{����nL"�O#��B�K��8�w3kq�W�:�N�7�{���U:�(�������X�@�·h���,��s�\�,�F��GKgY�P�xٻ,�E[`�Rt���y��{wi���[�؇�zLvp��Q��]9̳���M<n5���ۖ�m��U�G]M�g��3�l�͛z���ͺGZ��0��#���u�u�y;{a�x{=EN��]�q���-���ƌ��q�s�:��1���Ju�e��k�u,K]<��n�㎒��ڽl���>����4�]vN+���a��<���KO���v#��*uKk����=��^KLF�b�k<�N^N����6�K��j���5U1ڣ��mի�u�-ƀ����^�݆,�j��
�+*Զ�%�J�IR
QV�jm��E�-E����IF�1�%eF���m�l��E��"��J��J�YZ��ت�A��X��EFV���X��Bڌ�ʋ*
�+
�mR��Uk+Q
�
T��+T��X���A��eEm(Ņb[*V��B�
����AJ���h-ID�e�V�V)TB�*�(�U�-��(�(��`ŌT*��Z5P*(�*"����Kl��T��"�+-�* ��QE%d�"�X��iXVQF�b����Q*J[-�U��d���,-(�+Z@X���UH�Z��������iV��,
��I+
�X,+Z��+%eUYm�V�[KXJ����,�TU�HT�2��1DJ�b±EĒI���1��_T�gvܙ��`�c�TfG׆���kbpL̖ܡ�X{7h"8˶�7�ݮW���W����˫�{p.+:\�u9���nd6tr=:�g���C���N�y�����6�	^�lݳ�Nm��;�-�=a竞���Tv��
����x�[e@K�o�_��dN�?76#��q�B�7se������k{d�Иa�����7d�[&A��9
��ƍϯH$Wv�l\a:M��7�|^9:ܯ�5�G8/\�]�׬��8�N=՚�^'nx녇���M��˘��{G6{#�5�-K������Y'GU�kn.Cb����Ɨ��;�u���w:��3i{k�	�q�f�ݓ�b�.ͱ������(�����&��*��wk��V<��X����o\��8w�؝��^&;r��vu�aQz�����p�]���֮^�n�b��a���`���c"<���,lgx���{;k];#�(��i絽<��y��c<i�����x�mp]d�lm�i炈ݰq���UH�ƽ7�3���n���n���Y�e�[�v�|���ncv3��x%-�.s�gg�ۀ�Y.��j�t�qٙ:;mWf�n�웖9*��p�#:v�ζ�M�花���y�������phܤ�	�z;N�v�*v��Z��=�Ǝ�\�:v�s�	-���r��7�����.�노v�yc�i����8:��m��{[p`�g���Zw�9&ܙی%��g��ٺwxݮ8��1����A��]]^×�`!��kt���W|������	�.��N`D�u3�G�����>M����^x�Kd��e�Y�qY�[�������W��1���&3�N&�����ou��ݹ�=+���;�IG��sq�mz�ݩ�#'dh�kw��?>a�S�	�Ê��grc�T��I�@�/n5;���-4d7l���ۯWv�uǽ�{ʇm���}��<��Gs�Ȇw�s�	��m�睜���܉�ǝ�{����7�l�0烷8�#�>]��2��oo;�/O���*!�^�8;	�W�\nW��gl�/nawd��/;>7(a|�gq۸��y�v�<n^W�ɐx�2��8ܩ�� rv��e��N�vM�7 9y�wl�=��qö^\r�LF_���_� �j��_��=�`ľH����	 ���V�}��g+���J�ݽ�1/o�Y����j���a�(5�~�-��!�S+WKkd��V� >��i�0�m�C�ڼ��U.��_f�}���c�a���Ԉξ�o���[�� �mr7����U����W��i2�t�ǅX;T�l"�n\]��f���هޯn�d"=��p�"+�� ����ڻ�Ǎ���DI��l�}��Z�7T�Sj��h����(��l�Xowl����n6ӈh/��@ ����X�t�q���:H�6M���u�aѹҎ3�n��㘬�m�V�qj�vo�����H��)(+��T�մ�E�۰�:�3Om�b����$E�_u�3��P��B�TLT�6Mg{3 :�����ђT��_߽���w��Ƅx��jĺ������+϶rH��Q���fL>ƻ�"y�Tn������;�l��xFb&��'��|ї����� @L�|�w����׹�Z�:�+̨��2J(l^��i0Hw�1O��/�s��� @���&�]���ͻd:)��j�R��Z�^��c��.��No[d@�w��Ă +����w�^������;hX*�ڤ0h���wٝ!'BOv\��D�Y�qN�W�(��!�����$�d+�\�NV�Dm��h3T����xpu]t��q�x�c1�:}�D�'�m�qT�ˏ���d�jf�MQ3[\���7� e��� >�]��� �z���j}�vI&7�谽�N�6St*�NN�[� ���t�����T�m0 ��{3�
�m\C�*h[㫉����2w���*�D�Sd�w�� ��``/E��{�Yy��s�h�s� Ś�Ϸ�z���"o��ٗ�ו��=�%�o a����}u5�5X�r��j����7w�阊I*�Y���4����*	�G=���.=�����h��~n0 >���h���r�)s';M���>h"ﻦK쮋��)�tSTڐ%���0 ߺ�e>ʌ!�}W����1��z����w5�^&j����Q8�ᜎݠ�aMRr#� ��X�c��kګ�Mg<�RI��<:�L,&����nbX ���m ����q
#�LD�x�{���	�H*��$K��[�6j��'K3�8�g���L���)��M� �:���5g���z��e�$��-�N�m&�U���]f[� >@��m�D[���
W�=]��hD���� }^�m :}�B����EH;��E?8������o�`[�����j��x�W���^���WN�^��tPD��!���^�oq��8w���y'��~׷S���X�<�]옮u�2Ǩ�>�"��<��'� /K��*�J��P��������/��;�n�_��M�u{]����W��Q1��n�p��([�F�,�k�8��1mmg��^E{Vq���@�ۭs�ۏ/����ӕD����(�����p��  �z�٘��_Y�j�@�ǻ.|���a��H�r�
w�q� ���U�΂|�����޻�a��y��Nn�]�ɩ�����qlRM�骧��d��/�0Q t�V���ۿ2k���GW��CW��Nd�w�e��mb�����KK�o_��o��!�u�$�϶MI :�Z�͊��1�܎(�o���W�cS-QN��c��ϱ �=w�.�w�Y��U�@��c�� $N_vb���]�;d�5Z�2�}t��;�P�/���:z�֍'\<�Mb�+}~��O��W����}��R��F�M�ɇګ�/>�͕c�l n��&^I�twN���ܲ�)�.�`�>;>��om�V�k`LW���M����;l󎼥�m��u��Q��v;��g�	�E�����x�%��Fl��W��[��0/�t�Ã�A�^|����7a7N�lv������W�%Ӌ��w���@�d�]���ëc!��ol�sx�=���V�vt�n�=V���q��g�g�k��m�!�1�ۖv��O�q�F���c<���˶�&6��V��C�f�V��H�f&iM�����_���!$�w�H���ʕA�/�ż�p$I��t��J��UN�e5M�\���1�p�����y�ɑ 
z�s0 �z�L���W�Z��Nm��t�^�k�\I4��ES�>�nb�� ۽� ��7L�݇�w�� ���f, @$u޴��f����b��S�><��/&�=���w{I����� K�z�`]��{/�{-m������3����MӠ�a�a8��P�>��W�ͻ��i 
��s0$J]} ��=}�ɾ��s[��,y
Eh@�i�4�$�Cc�4�ώ�c��s���ܾ����X�������ۛi
�7���f}��A����4u��`��a�w���c���� 7���&��%��SE)���ך�a�;�=��{R}cNz��]��j���ա���t-��+��綅&��5���J�yO���)���W�wF�=�+�h9��9\��7��R	W׿d N_wvtI$:vݓ\0�v{i���[Nl9�Ҫ;Q2R�����7��P�k���O�k ʗ��sü���#��"�H���IX�F��
a&�4v{ݙ>כ��V�U^�>
��`�~�q�>:�w/)���wu;p I�z	��"���b��S�y� ���Yw�3@m+ʐ��݂H��w�w���w�'�PV�{�%��WP\=8��'MlY׫���ܖ�N���\⬡�\��P%4xfx�Zn�O�͸\@�*�u�� ����s".䊿w��<�>��6�4�d �{����"0E2]�Ԋ��ك	_>���b��n��e������wۙ�!�X�+֪b}7�����B�H�E��Ы٭�@ �sŀ���U�����F���Q�w �q���K�u.���v���{u�K*�H٣�ږ��ms=�.�ꮟK���ٜ���e�f��7�\��$�_ݳ�G��d9�φj���l���|�;�U*y��e$ -���|˾�� WshժCލ��q���~�M���\(`�n߀]��d9�I���[/g7ڽ]�S����ݰw���PI'� �E�������r�,T8�:���� V�����W1�s��Dp�7c����%�X1�����	��_�9v��h ˽ן` ��\A����,_l�bIz�ې��h�)�M�@�Æ ���&�x��.����]��|���~�� >+���dm�7"kܯ�6^�Y6�AVѧF�U���� 
�v҆$ s3�yT�]�>�w�|�{ٟa@��i��9���(&�.�7}����h���]/=X4yn �s��A�{�N!�
��w%�ujF���k�x�F��䧨�l��M���\�e��wA���ﱟ^Vi���AV����/�h4�����c��H�䏤<0:B�l�M�q,��$�{�&=v��a9=�ل�E���D�_{eč�Kg�|sy��+��w��+���ċ0�[N����h��#/�|��r|�g�� ���������=��q7��������v�0"���h+%��fS*]����a�s��`�o|�@��A��v�?v�&�mj�����z� ��[N!���o�M��yfG۽�Soۉ@�&�j�m�!ҧ�yo�` ��m� ��e>�i�=���s}� 
�6�!���m!/�z�AV���I�U���2�L���N�*�-��� ��+}��������8�G5xO�wL�Z��i���s+�D�M]d ��$H�:���a��b�V[�v{Zo� QY�v�@|u��8�{t�!���tn�|�lf��R �/a�����믂�4������k�d�$�V,��S�y�| ��o}��5�;�hc����1 ���"�Fݦ++l�'L'G��9/v�GM�\K�<��kZ��Gb6����c:�R�s�����	��	E�z���Y�	�0��g;�۷�"œ�9��-UV�;�tc�A$�錸�xn�n+`� �i�U�<'%��q]����Ɏ�s�@[GQ+:�5�Pk����v�yU���½u��c�f����w]dm��]AmVÄ�ۛ[�L��d��8,�����'ߟ�g�~���t-[�F��C �}��d@����s0*߻����'I����i�A�
+;���a�gU*�)�T�E��v`ľHN�]��C����p��(��v�@|u��2I��Q�g)u#�~"�G{��"�1S5rв�`H2�u��� �w�Wַ��w��x "�u�DC:�w1a`苃T���-�f��Z�_Y&���qQ}1 -��0��n��ĀA},g����tt$���zY3'��*�R�S4D����f, ���fϻ}��D�Ӷj�����t�%,���b$���Af��<7q��V�*�"h�Q*��xL�4���izc�cXǘ�X�j��Lw������J�**b��*�� ����0 ��HN�K>c��*��ܖLI.������<��S4�QSUP��;C ����d��ȰR��l�H|VQcɜ�b��ܠ{��g���c���E��q�m�°�絡CYV�7}ѯi�P��n�ܩ�]� �>��nf �_6�"#*tO&w3�~�̾I@�h�UQ)����r�7ٝ���>�v�3�>=�U��Q۹l��۾�� @#��M�S�w��E$�t]S��·7�ޜ8��j@w��^��ۮ��^���G�<I|�r{3���gT���-�f��\0��}�vN�Ko8������f@��m?�+�]��R�������w���KźK��Y�e��G+���g���lt]s����ۙɷϿ�����呫�O���D����s�	$>ݻ�&�T�u���{<�G �km6	���Q$�
�jShU���l����qu�ϱ��@ 7���E��|֬{C tv{���xx$�0�N�e�׶���[L ),}*6�����(� ���9F?)�����SЧ�,B�\#>ַVޏQ�ސ̄��6����ֳ�:�Q�s|4�zw,��F�|`��q��ǕFv�~a�C�}&`���/s�T��D�3՚�#;�Xd�=p�ۻ��6��.��~9��Q?y�W=������H��l����4��t	��3Ԅ�w^]7&��N�fJӣDWF7~�ݞ�恳���K �_C�_C��;ޟ�m)��.1ئ���:�5z]�ʴ��c/x�T���6�7�:ǵBV�_�E���Uc��nz���4xYSn&E���~�1�ul�z&Y��n������)}��š�_��w^z�-�����Yv���8�q�5gOr�@w/����Z-Cc��ʞ q2g��< QB�@���ڲ{$�+�ݧo����x���mo��x��fԏ*yz�S�?���`s۳�n��}��I��tUC�����~O0���Fc�Bcw�=���۽����^�1���{�s���b���ÓO9� 3����Ö��C����{U����.������W����X/.V�Vly����@ތ��=�!�F��˯j���[v�d�_k��C����N��*c&���oq]y��lOw�4����7b��kS�^�Dʚm%^��ZF����
?������M@y������������{��Z��.�6��Ƹ5�_��d�
1���t� ��j
JsT�M���ݞ����[�z���|���-�k{f�y=ۛ�o�v�t�}�w�������Sr�Oo_^r�銦�Uam�*��)j�Im���R����YU��d+
�k����R�Q�" �V�mF4�X��PU�+B��UQ-[Z�X��[j��k-� ���eA��**�X)DaU*%J1-,U�e`"�FFZ�
���QkKe�%a*"�,A������(J�h�
�H�����"4kPP�
�Db�,Ub���R�J�)*�X���FJʱ���H�H�%�EU@FJ��X��"���EE[e- (TZ֠6�2�,�*Ԩ#++P����Ҫ���
"�"�jEJ�J±�FJ��Dei*
1������,X����E��"�`,D�`���UTX,R*Ȩ�((*�)"�AaR���#Th�mXKJ���"E�}[!$��k������n�[�Th��b���:@�U�on���6J��7l�I$��v��I?��D�h�/�N�H��]I�躧u��H��*�^,7��}�&u`�ݿ4� Ew��@|:�ۙ�70*U�.����ϊ-���C�1{����Aq�d���5$��'����y����o�ޤj6�����'s-�{v�� �����>�S��r��sO�@
��v�_V��J!��!&B�����}	$n������/�r*�wj� U�u� ���c���գZ��1�<�d��D�s�I*e蚔�®�7� u_���ջ�ޝ�dwy�p ��۷�	��~܇5<
N�4�a=��(H�)k]��w� 	��p���o�ְV�Um�]s�����,^k���ʹ�Tgõ=������̣��c�5z��W1h�Y�~>۫��xc�ή�=�
��W�.�`*!�	#3��@Fb}�LJ��JJr�~��X ���<J�/�v�J=wuh��o�@/�X�{8b�==�S��v6�MR8�z�e\Q��F'ۇ8.���[�aq�4����Hꢷ�}���UE�uT����H$N;�y��H����C���.��k�t�3/�ɟ$�۽�����t���-�f%ne�A'��т�����Gé�@��w3DEv�M2 �)�o���r���s��$�D�BL�܉��f, ���i ���LWMMT?O�}��� ���x��"�]��kYI$�U5N��!׾��q�z/�۰w��İ� �ki��#�u�F�x�RWs~$�&�KW�I�a�m�Y�,Y1!��pD'��ji^SĮ��1 �+��l���vÚ<��#v,�kŇ[�FfZ�Ome�U�[ǜ�t'�.�o1%��N�t�&�=3ݺ&?o�=�yIw�wy�j^C�n����"��j������[A��X�� �ۡ���;�su����q|LW=�a�fn�`���vN�1뵮���=0�sl����×�5���>��nd��%�Rև�v�;ZG.�x�s�+���wf;:��ܷoAĵ���v�v����{6�X����]>ñ��.y1�Ů6����l���}-猸m�	�s=xsF.��xٸ:{4�k�)קvlqlݷ3�p]ƣ
�h�pi$�p.豵�{pc�8���6U��=w��߻��8�;L���fvf [��0�Q׺톾s���+v=��?, ���������
�.�T�D�gIi$����g�Uo��<� "]ͧ�\^�\�p��բ7ҵN�[�v���7t���-�f�̹�$�K���� �ˬd� �[M� >��]1!9�*�X�L4j�5
�읳���{�:����}n����D0�}�"��\�_�Б��ḇ�ŔS�`��3R�:�� ��x�ި���`)��C�E��4 �v8��ޖ"~<���F�`��h��űuB�g'ayD��tݳ�"{sr����~�}�?�4ݎ��������n�n�� �vf%��ח�~�~*~�,�x�u�[$/x��b��E;{����`ĂQ�h���ΛD�7��Q.��/r{�o��$a@�||+��ԇ����A����x��N�m ik���d�xOg��TS�s'tg=2����m����$�����I�߶o؊K�e���SO�� �
�]�B����U9P&s� �$
���}*�s<���/` �;nb"����`}�^\�I��UT1��_�g*ٕ`�A��m* �����|��j���d�{1A9<�r�'�+�,\����DO����v���'��Zs����3��+��3� @Z�&wL{%H������cwnY����=`�C���ˍT�]�6�\�h��i���~}����[�0�|���w�T �����"�m6�^�׶I��}�U�=* �&���$��E�H:m���,\�-��rR���ɹs�Jr�s1A��ͦ����_T�{�u�ɵHF	�Ҋ�
j`�M��f}��6�ڶ�
c�ut�-��/7o^_e�Ǘu�l��"�[������e�y�~BX����s��x�W�ua}ǯ�a\���Jc�l��{��0&$�K�5��M~��� �ͦ�O)�!T�L�QJfi�2���u���
�P=��<��"�lH�	/�V���s"`>��nc�t�ذ��зJ�h��P%W2�1$�|�m�=�y5\���~�Y�T��7� GW6�d }];�_���q~S���9e�����&��J�\;�n�櫴�����͵�z�e5�p�ɪ��5MOo�ֲ��o-���X�us���"
��r��og��4��s�4b)#���ḌMSg4?���.s�{Z��u�׬ ��j�
��r�H'G���7�kv��"ۓQRSUSJ��;V�AZo\�C�/\U�����毷�� ��DI_ս(�#��@��N�r�Ȭ��n�Dnz�|c@|�;C O�zT	$�>��]i�]5j�>qt��{���gz�bb�Us�6��U�wnLGw�w%ҽ���R��̝�-�w�~����~$����$J�P��5T��TUS�����4�D��l����DG.��[֛�����h >T�ې�l"�
��m�b���F�A�}���kN��:�V��\��]�P�����t��:h�����*���$�I��@����
={����)dǷ�b�'��ޕW޲�m�F��R|<��q-�篺���e�Ē	=[�D��~�q��d����Q��*���kj!���4�&*�M�_��` ��` >������k�[��>�;�_�|�~�ϰ��w�*�)���M�v��œ��ܽ�Y�n���:�ۙ� ��m��{�������1uF���Q%lX��XT:I��};�$N�ˀ�ڧf����yWo�'��T�$H-���I9�]� �!����ǚ�fv<��֟�;-uc���G@�����Nj�C���	޹¦z��:��// ?�s���|����e/e{��ɧ"�����&N�|�N��A��7C�S��������\m�ZX6�Ee��:�Ϳ��w���;�=8���[kmr��c�cQ�i}�q�x@�6{L���	O�T�ro7+ݟcn}�M<�{vDB존P�y�.��PauF�|G�p[V��ۋV�I��L�����x�s�w	B�ֈu�i��딳�r�q��u�b���E����t�vx�'t�u�hy�v;-�.��=�b۬�۔i��p��(���{u�������E0����^�d� 9��!$v�i�45��3�^��|��ۘ�>�#˚���� �N�L�s�G��o��mqS/kio��D��^�x� uki� Ys���/R�����%7YJ�2�aѪ,U���=�$'�K�Jg4K;s�-�t���䀊���Z�0�����5*iLUP�u������������y� Dխ��@.��r����8�@$nn{1`!�@�f�i6�}���HO�o|��ދ\�O�l�
��3"'��i2\��`呑Օ�y{�9��'7�&C�I'�m6��C�{X�j��s��|�N���<v��=�������{MD����s�c��	�v�3��:���غߓ�s~�h�os 	�m?�\�ZT��TS��)�G�%4��Hk����o�5�SR�>�w��٘xs����J���ܙz;}\��Xػ��+^l�ݘGfٛ�s��U�NL�����$�y�����H';V�����C ��*F�Ӿ~��#U�,��E%LK�%neρ����mσI /*��v�����}ͦ� ��e@���4��l&��Hy����{#�غ+XDm�[�Y�r� |W_nvtsE��f�5�� �X�b�N�R$���7��w��_ ׼���~��:^��!$�]�D�I��s*�u��_��au��bD4Y���
�����:��s���ܛ;$�\`��R�ŋw�����v� U3U4���|�� �zڠ +��LH��XJl�.�X�D�򽲉�F�����7�I$nj7�<��w%$���T	�����I
&s���z��^����}�h{�eIT��LӦz��� Y}� DVR�|��.Cx���p�ki���X����U���~��[�z�{�W��2/�����h�j��&In���?fO��<���{}:���}�������!{]�Q$ϓ�}�D�Hl��IS�v��?��l^�H�z�H$J���fb ��XU)~r�TǾ���堜�"���h$�Z��\��I%��l3��}�{�;BK��eL	��fD���w*#Q��0�Z�T�4��k��r�L������z� �b�Y��H\z��:J�4�&*h^�Ӽ� u��$���H$�$�z��2I��{Ք��y�@ 
��fa��(��S*�[�,�޻��X�����e,]/>i|�	/�^�a8���b}A"2�Cy����'�F)�,&Eʟ,����  ��nA�2p��Q���>� ��s>�&����ho�ʤإAU9O�,�~j��^"�=ꨯC��n0S��m �m�n먣86�z�ͳ��.��p�^}�pA[�P{�IA*�=��ޫn#���'���<�\Zq�t�D�K}��5y���
��>�3�����~�ϰ���U@I�H.�[��W��Tng�-�u�U�D[~�x� ���dDWN떃�ꁳ��?��N����m�$`�#q
�{.N�nM0O�V{j���d�����������"n	ǯ� |��[H +�vQ9��i�z�=��7s3�E�ʷd��a�R�D�1Ql�7ͪ�jr'�V�	�y� ����DӺ簓��wZ�E_t����r�e�S5SI����چ|
�n�
����f��|���i�@thF(-�D�)�A�r�˽;ً�e��9���V�eϵ�DC��nu�����G$���a��JߎD�JID�:h�3��@ ˿kŇyz�ݍQ5�@y�ӈh�=�Z@ u߷3	_UZ�����4�m�!~eXk/C�7�I�}�П{�p���[s�E����8!����6�R��J����]�j?>ˊ!�w�F��05}�zqM[����'q;����%�Rˋ	ݕwb��D3S�!ܷ��-ᢙhi�x�X�p�l%�����7멲����n9;�P�����²Rc���L�.��.���,����݋��o؉��b����n��7V�OX�o�8��4�=���>�g�/m�A[��7 ��FsZ�J���пF<}���ƀ���J'��S'2�c�.�{]A�rڰi�ڱ�䉵���#�ksx�׆�x�t��/��]'I������:e�[�wN0�3F��sw�4H��tcKb�Y���y!�Kӟ�n���¯.x�����.U$�&���.�����A��ɇ��2n�ͬ�.uX:v�p�l�[Ѻ���^�/:TxD�*�!}������H �����&C`��w�§i�ٝbO��3��پ���bS|~IO_�B����]�r5N�ݱ{��\���x��A3�Xwu={f��$���l���a����]��H��b�G���%�%�������[��R����z)�f�A��D��f�*�s��2��=��1U�?mF�^�3[&��ƍ�l�/���s�O��w�;��2:�5կ�O�����V�o��b�0�9YZ����Q�
�K����ҷ��//K���qw�(�L�MB��X�b{K]�D�;4���{�\end�>�k7^^n�7��bY�F���`#b��X"�YV+]�R(�(�UEAJ�R#TPb
��++i(�T�U��)mEAH�Ȣ����TAAH���c`�
�(�@D��TPX�
����Q��`��%�ADQAb�1jTU�b$Q���"�AVB���U����QTD���aQDJ��R,���j��1AEm�c$DEUT�eJ�Ŋ�J��ej�P�X)�-�������E�cVVTPDX�m�i*
"��Z,(���J(�F,��IYX*��l� ����`�U�a���(**�A�E:ݿ\a1��(�N;�ۃ�]39��4s��{S;�Jv�g�jzv���-�S�<�\����(���W՜^�6Τ���T=W=�I��m(�"��nN�k{�Dn��۝���'8q�f�������:ⲃτ�g����۩Qci1ۉݑ27���=�ӹ����hd�n��lu�sƱ�j��=�J���b��)��\{q���u�]��q��d���[s�t.����۵8�1��u5�C^9����6��^<g���絳v���y.B�k���6��E�#�x�6=���u�+��am�5�S��Xl[�����g��R{w!<[���w+���L䛠�A�9Q��q�2q��<]��.��;=X��x�fu�����s�[��pdn�)��t��w+�ˊ6�˻�c�����r�o9�/���t^���s�oV��oX�<�G����C��vN2�q.�g�K�A���Q�X��$�N�ޮl W�r�T#ۧtW�t^;���ưq֫qǃ�����ƪ�6浻1�a�ln���)ƃ�y5���sӮq�k���ጶ�8Sv�b��k���v���v���l7;"��r\t�k[����ƺ�K�E��zӷMƌq'8�uq�:6N zqq�=�[`�wi�u�s�;�v:68���d�D]��GO�+��훎�;������=ǑF�ЕӚ%]t7gvn�og= b��:$y9籓vua"��`��Ý����e.y��wgs"qڍ	�W�&�k����9v���[��G�ۮ���1Ns�	���D�X�+<鱭�O&�Q�N	���m{u�8��B ��q��g���í�>V�v{g���9��ػu�k[��+<v��W1��ٮ��j8�\k�q��؞�kg[��zV��su�<�����mp;T�^U��E�X:WpZ��t�cu����܈���y�۳l:p�h��K�Ѷ��lgBv���<���ӌq)�m���g2�{��������L�Z3ɝUf{{s��ڳ��O�6-�ܻ�l���8�T4�0s^�^^�lF����`|w'of�Sg]g(9��n��k�q�<vR��	���Sӛ��3�V�]��z�%�v��=Y�x{p�8nإ.��������r�Qԭ�ir;�z��O	�����χ|S�#\/km�;V�w=��^��Ȃ�)�<qAg�����v�s���tޣk��v*�9���<&�v���y	�TZ(���I�?�,6ZIc�� �~��0�v�  u߷3>	{�er�Э���-���Ȭ�i����[�$�#����xV4d.✞�&�DD��j tW����nbX@�jny�qvk-����"jjB&eT�C��ܿ+�A�}�0 ����<�@@x��M �~��!ᕠ��A�7L\.����'�6�w�J��$��[��-��f`�����}k��B��wz��Ҕt�$�QJ�����f`�m��J��{�����g?;aw��K��"�U{秷%��E�]UA���;7VT�E����\5V�=v�cHc�ا��`RA�y{�Q%R�Q3[\�]��`��2���� :�Zm,�W��W�{&�]rY0$�]��1Y'�{��f�@�+����08���޼ڗ��v��k�
"���jq��=�۵�Fw���s�_8�b�������mQ�b\�W��[g�&|v����SnÙ�� ��@�oF����Kl�ϵ����[b�w�A'6�N�[�R��'��k���D����%�����XD]�� k��L(������� ����� >:�`�(YP���5M�L�C��vuZ���)�wi ����A뽵m $v���á^�d$���ϱ%0��Kn���6X�.~� �"�z�V��W�}h�o�%���""1�֛ k�eč�M�ܲj��*謢h0(�F�T�=��\��A=sA�]����j�<\�q�T���ztQJ
P"�d��}�ŀ�A�{pĒ	Q��q"}���`�j}�1�`	w�6rr��%R�Q3N�Xo:3�8#w�]+���f�I�����l�c�n�� �;�N�ؤ���VVDm��U"I�A/2����nȁ��ͯV��49���'��w��9��x���7��+�(����nY̕c+��G�9���懿+�2"|v�����ݐ�����5-j��i�~�O�u}�_$�^%�g�D��6B	*_�c�/���X]S��Tѩy��;^�x���K� wc�m �Rg���	���/�t��༖�"қ�
2�*&�P�\	���K䉮���>��Qw[��0	�m7� ��s��	%]~��[�7\����e0�?�,>�N{Em��5ˌ'`6�[�0j{p�y���_��������^���Tw�ഐ ��ۙ�Ju���G<����d	=�t�w0�J
PJ�4�����K5�Ν�fQ��� �z���Y� @I�Κ "z���DKq����W^XϢ_p��4��*���/��	��<� �=��k����9;�XD��vb�VDm� �U"�N�.o/�}��L������� ׻�����+5���[�x�sT���\��*Y6�c��a-/z~�?ĒJcIGW�	��Xw�ϲ���u���|}^�Goy��$��?�|>��zIٵ�(�����:l��Qb�	����������s�h��fV��t�ޛn_� 	����=��L������������6ە��Tᲀ�:�Sx�{��.Y�`g��'V1Oi3K�����1߽7g��#��%@�A=}�0 {�M���u��^��޺�y*|�)W^�C�f^���[|�we��%;0��{�R�n��ު�����=ͦ�If�F�E�z�2��(��H&
`��S���}�� w]�i�O���r�.#}�e{��� ����/��Ot�E���&�b�T�k������Doyߡ��7��	��W�@WW�UWU��s��j�nfbB�;}�L:����e�	A'��s�G�c	9޾�f$'��i�];�X_z/R����@��v)���:��CUz�/&Fk�f��Gc��Tz�?���{.�!�-���C�b�GV돴��{�M�  }�ǣ��_i�ARlq�3��i�g^.ۋp��n.ι2�Z93Ʊ�t�n���X���m�vvw�(���"�޺^H�B�X�
����:�b�l�0m̽9��g����tl�f6��;���c7Z�l<��K���;u�c&j�m��;z��F��E�x�cYGgvH-�6���ۃ�j��A���lvL�ݥ�u�λ�19�w��k���\v'��v�&�Uv��O7����lm�۫l��iM�Øt�4��o�O�ٟb@$�J����"P}[���qݫ��f��5�*}���I �Y�+!C���o���6�؜{�sڶ>�?_��� ��m �ݹ���,y��{�0�_�-�J���bD��.D�[����m�G6z�}�|]ͫ�`}];��J�%{R	��&���3�@bl��]Yh ���8��'��G]���D��B�nY�y�#u�W��A5H%5u�fst w���U��n��Ow�m >Vϵ�@Ju�n`��w���]�oYHAH�v�N���8zB݌>�GnεuG4i*l4��[�g���+t�������6�䣛s�D�7m��#��[�I}v��&�>1�}%|���>�3�0��PthS
���H����w�f�ǟ��gK�/}�yN���Xڵ�=�[A�G	B����⌯[+����|�����]׳]���2���V@�*� � �-ߝ�P�U�~r� �Wۙ�_L�FQ��!̮�"V*�!��b�N��6^��1ê���|��ޗ1�'3�k=^�ů�WN����s$��
j�J���b@��M�~���߳�r 3��t ����!�\8fI�б�(���6TI
�J��� �*�:g_�� n�il{��j�'�Tjk�nZ@ ��fb+��p�ǫ/���꾘N�h�n��l����p2B[ێg����9�u��6�E.��x���AZ�i�j����Ƴ��H�w�� ���p�s�7�*�N��=Z�����2��3CQ���� Q4���[�hbR��YV���iy|�> U��b u�����6����w������X�Fh�S%�	�-�q�� :��C A>�My{��c՛��,�d�޷k;畢��ȶ9Zhf������֎���^���2��Bi{��b;{n�*(j��|��E��pK2���J�f��+�_}�������#�#n��0� ~��&��Q��Pj��ԁ_-��&c���7��&�=�>�I+׷��� ��eU�}gw�� F����>20�UD��URJm-�9����끯�٫�:�6!�w��������m�L�����r�J�b�Sy������I�,���M�ڴ\s�A�b1���5�݆J$QUT��Kt�A
����"��a�wno�${WaI5����p$l��E<��gH>~�6	�Ey���`�M���� =୳��fz�zI��`�Eov� ���_���^n�/}��};�j�Hb@U�e�� �{��?	�V��^�Y泶@H>{Vl�����#�%T�A�B��.��H�M}��s�t���Y��$T�l��H5]�l龮����p4r�bůݡ�'*����}nz��z˕h��ǌ ���h빪����;S����9�e]K!��|>  ��5��lm�(��A�f��w߽!�~�I���g��b�od�=A�1ٿ�"���$U۲=����|��|I^�� ��Æ㮺1GM��z�lgOe�	8I��T,2<=���H�[J���D�]��	$EWn��<�.��aX�	W����;�����iUA"�4w>�>��������Ų���"A��l������7X���U֛3�pz�;@���T�\�Uf��� ��p�{��fqU^�$���H	"��n}��S�	ِ��76�\�x==���@$ ��h�%!Z��`T�Ͼ���p@�P+k�ޡY�w㿳���7��:��A�߿h�F����9��Jf�3�p�AL�>��I`�d��=�gz7�N��~��w�����%@�g~��$�S9���9H4�+A���a�E߷���+��0meY�wv�e|���m����%�/e��s�U��Y����W�[�������⯂�2�[|V�Q}����آ��ڵ�˨����p������1qj��+ױ���$�.�q�TY&1���ۧ�8�*K��&������!��ޓ�	���{v�w=�9�[/��Xy-<n�F�u��]n��/݋�nBM��մn�6���:�=��;�݌���^6�tr�h�[�S��-�8��ؓq�s�9�W��u�:�v�b�1����5������G�&w!�0������^�[Ń��g�v0��������i硲_�w���y�q9++%ed����h���Q%H,=�gz�a�'9���w[��8'�{���N2�Q� �3���8�@		�T�	��U@��@
?�����8HR��z��;;}���:5��ѿR��0*c?{�i�
�YD���� ��IP��{Yw���C�����:0�.5�����L�a�3�����Ad��ú�;Ѹ�2XʁA*5���~�>��Ͻ�`pk�!KLg����� ��=��/���'�^����[�T� 2!���h�{8����n3�|�J��S_~�4pI�(���+k���XlaRT*J&}��G?oۗ�u�gyv[~� ��~�D�8�O��?-��	h�.�085�7���n8HYi
$ ��X����l���3~L����h�"H,=���B�c%B�*!������+���_�~�;���~�}�n.e�׭�q��u��;.�nz�L9�����eRo����߷a.:3տ��{�§�׿h�N2������`ʁD�=�}��`c����g:�?$?Zk����R�+D=���B�`R�r��A�f�� �?z�#A #�?|���{��e��ݕ�S����պ��W{'=�Oޫ��Ω�dދ%}}�u�zE0eSgk#�c�=%��Z�a�/ �T4�՗�>����G��w@m�%aXV������%B��3���h�'VKY5����A�w�B���}�0��A,r,��m�.1��65�߻��!�H[@���o�HV�+FO�y��c>9��Y��6� T��=���B�q��D�
!�{����
5���1�-X&�|0��"��~�;u߳���3��N�T���<�+&�R
�w�Ѷ�R��}�����c��{܋�!Xk���P��J}��c�90����s�2�I�>��ND
��YFJ����Gqk�GV�����ߋ�|M��
��<�w
�q�Ib%M}�{G9Y(��`ʘϻ���Y�=������^�ST�x��tB�"s�׎��<&�v�t�RY{i�`O���߿��b�^��>`z5�5���ۄ�H(���F�)
����
�c>�v�L�y_�z��g�{�?�|	�s]�*AC`��P�?}�a��a���̮1��3\˨e��T����D8��VN���/W�]n�W|�����~�������~��8��X���ϻ�Ô�i
��v�U�_���^�~�+�J ���
��L�e� F���aYFJ�2T�}��pI�*J°��~�`��0�w�^���ޢ!��m�A�Ca<w�^��裥Ex+�]�*fi���@�>)gy���מ�h��]��T]�L�n��w�N���v����#��7�oݹ����YŋlTvB��!r�_0��$�*غ�ҭac�зT��]�/3�n�<4O#���-L$�����c�le;>�EkR�=��<��fɠ����,b�qv�w�Yל=Ԩ}�s��e��È�=4sR{�]8��w�dB���2W��MKtc��l��OX�Z}v�iI�6��h%=#پ)����8��ͯ;^)��Q8�&>(Z�ƌ�f�;Tg�����!�{��>1a^�Vr��W�������gG�?;9����w|�ug,uP[�����'�g��5��9��S͘�w=⎠�w�tj��7�7}�(�ٲ�SUV�L��Y�nyy�=
WN�Q4*��=���pj�[l�Kt[wP�fd���x�@f���	�|;�۷w-e���r���{�u�o^���zw��D4�W�Xf.�|���s���1��PSۆ����ct����FXX6�K6�5_Vo��@vu�U��x2�U����}��a���=���wSk@#�z���s��\!��kOVu��vW�	9��i�f�@̭ʍ�4	6C����מ����F���j����ߐ�9��_o�ł�����f����9*�z���oL�ɱI�a�`��_��������J�Ƽsp(���u�M��L����B�H#�b����X�X*��((���EDbX�X�Zʈ$QEU`�*"ŋ��X)iTdU ��`��TH��*(��"�����*��E�����,R�`�)Q`�+""��E"*Eb#TX�h*��`��b��AE��Q�V*�"*�,R}h�FE��Jŀ�[E�F,�`��D�b��@U�ɋ`��J+$T����`����ZЊVL!Pj��*��"ŨX�1��S���*�(,�ŊV����V�#���# (��-UX�E�"�.#"��J5��"1e�DQE""(*a,X��1F��H��1����I!s���
��aR
J'���h�'Y,ed����w�F���h&˥Ua��G����`{�v#g��w�Ԛ���a!�I /�o�7�h��q��݁��K+wyޡY��W~�O:��>C�*k���8Ã
���d��ۑpd���T����i9+%Xw��z�d�F���/ܙ@�P)�o߶q�ư+R����8r�m!Z!�/����Z�مxa�\]U3MkNy� �sպ����z^��i��u�.Ɍjj\ji����k�a"�¦� �����h�AgJ��S������Q%aXV=��{�a�¤����������IS���q �r2��}���9�ϯo���Zf���Aas���~p�Rׯ߹����9�{�7��+X �3���N T�ʞ���B�l�
���o|�k��\{�������2b�&93�p��*sz����B�VV��f(ʐP=���;�i����g�<����S���6�yG�@������\�(�n�2��s�6��=�{�L]��y��ï?�y���T�߷�Gq
���+�o;�+��(!RPN����2t�w������_��)�?\Sp{3������^�f�6b��i�����U3�S&����ct�YO���:,/�K�&vs��7� !?��?������w��8�@�q�����%�\��lXÿ�gz������h�%![{�^?w��c'=�@�AO�����p@�P+)����
��J�T*߻�a����_\���.;���1upzS��d����b���g����8œ���nsB�2���3UW$��&���H�+:wA�8��R���F�a �T���}��`{�w�{�8.7�8�o>�C���}���R����B���+�L$S��T� 2 ^���m>� �X�u���ן����w��q ��+��[�+����}�i����?sx������y���=9׷��gs-�s��`p��j!�H(����0*:��c��_�����O*eN��oP��d�T����h�Aa����U�T��lσ#�H�}������Rq
�YX{���6�2Q��@�7�wgk�!KLg���?�K�g;����k�oP��Jl��Է�f�g6�`q8$��ߴq ��%e*c>��8��g�3�c���߉��+
s�k��Xm�IP�('w�����R
ALg����w��eŷ���~۞w��R�ʲ��ѵ���)�<�#�S7/6=����x<�u�ݪݻ��B�������&��o�}�}��~�~�M�����)��Nػ��`��n29�vŌ����f@���^��<�K�ƻN����)7n��t��X7���N�m���FvW�r�㍞�j��M��{v9ܱ�� ��5�x�����.�E�z{i���\
]�4��V�q��P��'=�������x�g[+�n�͂�t�λ\��zz�S���&��֌�8Dk7e�p7\>K��Jzf�'�^��6v�t���F��vj�W����?����i��]��5���y��� �-�}�w�7�HT��K1�w��3�u5�~ֻ��q�[��+6�P�J����h�
��k��v����pd���3�����q%�VOc��oݼ�Ͻ�����Y�A�d��J�Oo���085�Z���ϻ����HV�z�s�?Gys���G������Tg:(���H,�����1���	8�IR}��y��[�ߡXm�IP�߻�d�+%VJ2�3��D��@���o_�pܷۘ8����W��z�i?;�޽�C��@=���򐭌
�K���v
p+*{���
�w��9�z���$0!��o�8Ñ�a}��c��[����]�,6§7���q$�VJ2�������2o��=���׿{>�@�	P.�������!m1���Ô�JB�k�ޡR
oy��<��滍qo:�M��ks�2�1�a��y��x.Y[�cc�۴�pT�'T(��HI���T�U��������e++%Lg�{G"N!`���+
׵�¤�����}�wZ���M'>��h�'Y++%T�{�c��� ����t�Q	��*���,=����	- �c_��w>��~��W<EF�ϯ�k"�>�_�����4s�DY���Y�����l��B��9����jS/lܽ���������~��HT��K1����8�@������Iĕ��+��8�o˫�}����0�)�_~��3���\3�q �?w~�u$�VJ2���M�B>��" H\����I;��8i�5�Z����{����HV׷�i����V5��t�۰ ����FC|׏�1�\:�Y�1�C�H ��5�m ��g��CL�������熽�}�}�o��%���S��ߴN'/=����%�c�8������i
ZB���}�����s�c���� �?}�w`q8 T��X}��0�6� �g��m���r{7��5s�m�w�l�h��Z(�XKL�����=�ug�ឱ����:wV��h����Ơn�7V�{����~��q%" ��f�+*�S=�}��`x����9]8�N}^Y��x��Z{��t9H6��(�c�C�"I��M�Ҭ��l'"M{��G���J�s����>��'��7�h�N$0�>׷�i��
��P3�w�6����YY)��~x8{��>M��sD�@�1���B�l�j�'� (�7��0��H|[@����7�R��R
w�����9ک������^A蹧���ze�ѿZg�z�����{���q�[�ߓ�^�{����pU�n����yf�s��HI�ֵ�S�@�P+('�����*IP�g����$�\�l*O�A�~���?X�䮼G��3�e��+%Xs��n2�Q��@�����08Ԃ��i���`���u��U]�9_�x|�P M���	���u+�)'MP-� dAs=��ND
�2VQ��3�{��8������a��m�XV�\֠��
��T�3���$N2�VT�}���@�<��ث�Z������h�n�ݭ��ֺx�6�jKdxv@��/-۴V}��ϯ��|d��L�q�F����h65!m!m>��ѾR��Z0*Y����'"K��}�k�~g�M�[ޠ�l�
��b�}�a��?s>�+�ی�\d�]�,60����pC�,B�}��}�������}�����@���`q�
ԅ��}�t9G��>�H�
�Z�W���~�=��'��"����۠�T�U F G�~��8�@��%e*c>�tq'�+
0�1ޙ9�ko�*J!RT�߻�H,�Y,eLg�w@mZ�j��_R�(���G�����¡��y�w��-!B�5�w��!Z0+A�R�>���*a�kz��齧�����9�����=�u�jS퇵r�z(x����$��e��r���$=�{�/�5�Y����Y��W�s�HI�L!�T*�{��$������&1s3�m�хL������!ĔB�VV}��F�Y;����.{���>H(�����`q�
5!KL����)��j���Av0*q~���?��k��8����$��kv������Y�2�DV\d.��z;��}����8�q��s�2�Iϵ��8�++%H)���t�����+{[���¤{�^����v��m'ɞ���N2�Q��������@�_\l��*f�s�`v5�5���l�R�Ʒ����ε�w��F�R���R�>����
�X{�޵ �;Z.��� �wv<~~���4����7&r�H)�g}�I�!Rw[֍���eH(�s�^��c���c_�k�!m3�����A��j��a�D7�E6�"�1J��Mk߽���g�yy���ױ��|�FJ��S����8�IR��z��*AID���h�'�<�q���~d���p|Fl�w>� ���vy&�?"�,	v,�a����Ƥ��w~����ޯ��`m�0*Y�k����
�Xw>޵ �6!�o�ч��?f�{�z��g�\��7�Wf-�k�=��p:���N��%�_<�`�'�*ӝp��lnz����M���v�:^�%�n3���~Zkt����}��q߿<�&ΜՍ������{i܍Ơs�.��6[n�ӻ�r�rGv2���.��G����۶�mp��I�YN_D��mtu�:s�9�,�=�8�m`�+�zGv�g;j�nż��
>}�+�^�MU��g��\�3@yqd�/����]1�9����[u� �v]��u�9���4�ۨ�ɫ���r������M�:#թ�����.T2����ɫ-gnDM����P�wy[I�h0��~��}�~�q$�VJ�����h�eH)�{~��085���o��u�v�5�R�ӻ������؇���P]�
�{����\c���`a6$ǿ{�N VX�Y߻���?x�;%Oo=����V�aO���pXm�IA
���o���N2�VVN����_wZ9w��B1�폴��:��-R&nG8Ѷ���j
Cv������o���`V��z���Y�_c7Y���J VT����Af�*$�T=���8Ì+߱��8�[s�nF���O����
�'}O���wpD���V�ߵ�q� �X��w�6�X�H[L��w@}����w��AH/���oPR
l֝��K��sq��ֹ�O�ed����s�wGq�_�0ןo߉X|°������
�P=��}�i��+%b!���>�F�jl����)|��r���Rڝ �u�&���cm�[.0�v�'�r3L�ٺ6���	�a�#�O�;�v����)h{���|�*Ak�3�}݁Ă����_~-ߎ�8���?k�ޠ�c%B�����ѶaXS?<��g&1s3�q�#
���~�O���}��څ����UO��/n��8#Qs��3�~��+up7[��Z�Q���=���<5晻�{^�=C�v�4�M�J���&������}������kG�*A@�T?������F�,jB������9H6R�q�ܙ�M��������+���D���1��:	���}�G��2VVJ���wGq
$�(°��Ѭm�/�����`��T{��ѶNA� �P~D7�z��� _�Ov:M�TYL���Q�[��y���ԙ�W��
����h�%!Z
�K�{`q8�R��?{[ޠ���i���raD�ƾ��q��aϱ��g&q��nL��2�S<���6��B�X���kzѱ��e�y��~��T�{����XjALg���99H4�+����.�K�����~�9�T�uۈm��6����뭰��v�Ķ���]Ʈ֋q5q���iN�������O:��ww���n�w�����e+,d������'�J�XS�k{�����ض��8�[v{�y?k��G'Y(ʘ������o6^�8���Lq�`m�=�뿁#�>	���z���bZ_ k�����*Ak��~�v�@��=���Af�*%C��}��\���s��8}�}�}����q0��3�m�T��{����T+%X}���Y,e@�P3;Ν�۞�ox����QLä8���k|7q?b�Ya��l2���Ex�n�
���nNqLO��I���o�S7gK���n��BA���`5�Z���3��hNR)
���oZ��
�_b��&�	� �!W���E�����w��6�Y��������$�%aXVw�����%�T�;�w�8����1n?�q���������FTn��X�>#}�	��I���)��~Xc[��AHn��=�>����;���^{��$�5�s`q9*T
ÿkz����T,C��}��0��W`����~�O�^�$!):!S�[��糶�1�K�Di.zu;"���P�q��~ާM���-���?������`a%ea�kzѶVJʁR�w��m����}�{�s[�y�{��R
s��tg)�����P]�
�;7����ˇ79qq�8�I�o��q9++%g�e�������&���tu'�+
°������%*J�߻�d��#�O�U_U~)�W��{�����F���"*b�u?G���h6ԅ��)ho���#~����R������}2��4� 
� VQ>���Af�%B��X�w��Gg�}q�c.f\3�q��O��=�η�s=�L�1�?$��d������F�R
J����h�A`p
#�H�����y�~^�fl�Vju�IU�2H��{ٳ)���ߕ���c��?\[�Slz�{e+�2e��u�q��AC=<��`su�e|��?���!�F�w�������e�|��:�pg8��;)�I���ߴq8 VQ���~�t�η�޹�}�����,+
��w����
�RQ>�{�d�*Ad������8	��>��_�K��ytc��6��:j��Tk#����18�at�����@��S���T������UE��o����Xc[�ZƤ-�-�}����R��Z������ND
�>�>���s�g|��{��Y�L�߷�,��P�����a~��6�N�-4ِ����뿴�K��Ͼ���r迧^wz�ѕ���*wﻳ� �8Zg>�t9H)��hY��x3~>����L�	��Ιx�nr��@m8$�w��8�R82T�}��pIĂ+?�ݷ?�o��7���a�%�,Mw��2r2�VVJ2�s��D�q[~�\�G¹ƅ��������˟����>��$��|�=�i �`T����v��R,O{{ޠ��kY�~�CPIP?{��aXY���ߦ3�g)pd���#
���{A�8�� ����Z62�}�>��u6��*��|����R
g?}���AH-�����N���7���ޘ�������M%��� �F�6�v�-6/应k���K�!�t�=�zys�]��-���Lo��.���]�iu��zjܘ��D�w@�B^뛏�R�$����|{ye��|/����i�7;p/#8{�5�K��e����Ԝ��<碽�W=�X�������;��Ў<+Y��v3���cEr9g��D`��D�f�;��p�ٺ��5�0TfVx1�^��D�=��zk�yǈ��%����f�K�^,� )�vkà����"~�������U���n�F�|F��/�D��{	�1�YW<7��Ku�h�].�4�@
@�	�7��w�'`<���p�����.%� P�I��A��T۽B����ӛ���g���3�~
�5��3ے#�9�r��oU.��|�<�A9��T!`٢���w����|�{u=��˿/���GƙX���i8W0&���q���^]���)�*��3�w�EJ"f%����ڗ��JTgtO�9[��(�{���j���N�2	���o�E5��y�����R6h",�W���W�>�#�����(gq=�P�����~UOF��d������j�՗���^��F�/�۝�zvo��-
'	���]��{��ܢNȘ��NU�'���t�M�?1���3]�5\͑gIs����{̯z3���w��f�S��˼p��n˯��zM���a��<�J�%u���i�=��#�%�x��y&"2,V2*���
�ȣETmW�Q����TI�DB�E����+�*�(�I�b�[KeZ�����Uc"�A*TU0�ʅm�d��b��d���0� �-��1E�
��fҌmV ���Z�TV
(�FإTQb*

�,UEQYb� �L%�1b�a���Qb�H����d�`��DL0�*EX�Fa�PVT*�
5�S��b#b��EF,ک���QH��*���F�QUm*�E�Pk�IX��#"-L2� ������
�QDE���-,��T*��ł֨����
�X�Q�V(ŌQ�*�pʊ*�2ڨ��QU�VUD@UFb�b�"bʈ�(�,Q�`�A(��QQU�b(1E�Q�F2�`��"���������ы���2���0���`Vz��}��S9�c�N�o\-[�����[p���uζ��)�Nż��ƃ.+�(&��Q�v����uh�����]��I���,�ya˹�}Hrq=���9��a�
0��"so)n�.ۦ<���\#��[wf��\�a� ��e���%Ş��'	��W�Cr;�<G�� s�l�����z�7����L��u�";�N:��^��]�C�؝��n�\�tX�!�K۞�g��`W�5�^�zk�j�d���֪)\��OZLS��{S7���=����Ai�!�ڕڤy7m��Bv퇛���۪`C��箹�a=�M�s����˻��hy8�Ľ�h�q�-������7U8�N�3��ZdEC�!�[�Z�N��%:����_<o]J�r3�����#��M���p<v�lw�n&����-�������[H#�7gv`z���[��=8:RU��6��hƊ�Yvv:Nvyg���0x7\���I��긶������l�3�t���d���^8�{Ӥ�͞�w�u|.��=g:8^��iD�]z��V�x��z�Lq�p�i�����Ė<���ݛF��v�n#=��Vyx�@ܖ��c�P��t��:�6�=�n��cXM�cq��n'`x�1��y"��zש�4�3�'v�Q�h1��g�n�ݱc�8ָ�8�\X�j���"��u9��۰���Ȃ��O���!��r� ��v�f���ng�X�po�g��9+�	���w*�'F�ܛ[��01�2٠J����N���{�}S�H�k�9����h�ݶܼ*�e���۷q^\槩ވ:�n|`��ݵBv��Ոnt6RK�ǎn'�V�/Nwˆ��l���m�	�,gk)I���<����웞0����Ic��V�'�u����Bn�1�ۖ��a�\zma	�n8ςyUӞ�scv�A���g7<ӵ�8ݝP���`x��������?p���ƺ�7�K�N�ݳ��]�m�l��`����l�!t��MG�ZN͎��,�!���\�!���ڍ�w\�Le��wz������ǋ��M��e�z�����7ޚ
�E5{AC�L��akN��mhb�a��<v�#Y��γ�0q��^�s���������u�w��e��j�,w]k�:x��R7��`�p�����t뤤�ubu$G���d��h��G�˻r�,���L��*�p~�����\l\������D�Ͻ�G���� �s����N!`���+{{֠��
��s�<��g�w�m'����8�Y81�G�C~� ��w��&Ҫ,�{8��kk��)���=�d���\s��x���F���k��R�>�v��R�VQ=��z�ͲT,IP~ޱ�q�\�=��oG�?0�,�s�6�
���ٟ~�/�`g�"Q
�YX{�޵ �m*M=���>��7�{��jAH)������i
؇���PR
ngf�{3���6iT aG����0��y6 a��++%M�]��$�$���^����
��*J&{�{G/=�~�=��}�va��+%S}��N	�
c��e�qs�U�6)�{���֐�h����)
�[�����?;`T�3�w`q8�R��O����,�%H(Q����0�
Ý���9�s���~��ԫ���\'3�ڷg�np��yy����yx�۠S,"��(����-�l�A����aS?��h8!ĕ
�FVk��F���YP,J����Ѷ��q���c�|R��=�h�)
؇�d��0� ����f�LS�K� 26	9�{��'++%g����{[���?O�<��Ǧ�b�w�#���p�n�g����Ò=<����K��z?^�h0�#3Vo����ڽY��D�A�Ϲ���_��$$��L��G�I�*J°�/����
AI�
���������ed���_������۽}2�:��'�@�N��&Ҫ,��pa�(�*���R��3��{F�HV�+X7����]�{�oW�o��<@������,��P�%B��{���S�W��6�T�n�lσ?~��ްg�~�ۃ=���������3�}�eH(J�C?���q �8ԅ-��� ]�_�Df���bQ��/�,����gs�f�..6�3��wG�e++%L��{@m���N�L$緽��%B���׾��2ped��3�{�'��߷������2���ۧq
�Y5a�x��NCn( �ȳ'a�¢���V翾���bݹ+s��Ѭ=�~փq�
����w�Ѵ��^
�9���8�*s��q~��c����lM�{ޠ�l� �P�]�tq�V'vߌ9�1�pd���3�����q%B�cz��c8֛�����2�VT
��~�tm���
5!m3�{�i�HWƿ}}k�6-����뿁<�"^�ʚ�ܘ�2�����g�Ѵ�@��� �3����8�IR|w<�����������=������D]�#g.�h�I���W5m���9��d)L�O��Ս���~ޡu����5k9�\.~5������w��%�,O����G8��YY,eL���� ����Ν2��(0�G��������W���- �}����򐭌
�L����q�@�3��Z������(i%B�o����0�
�^Ǳ����c5�pܙ�2�S�׹���Ad�+��֍��k���|���D�~��͜`r5 �)i����9H6�lC>���.��S��~���K���mA��B�	�fĐD��㝒2B��;��qu���$�}�w������3��Ï��Z���q8 VVJ�S9���C�+
0�.}��pXl~����f��D��K���'_z�2v2�Q����s�wD��@��w��2�b�.8ذ65�=���ljB�������.����ӯ�� =�}���>?��Ͼ����wz4
����\\��n�$P�ԽE�[ �%���M�
��� �q�I�f8�^A>$�gu�	]������MQ)�t�uV'>������:@~+:1d�[���C����n���dh�.���fU�8������,g��������Eש�w��%��W�e#�W�,I�x�[�z<ZQ��KswQ�|i%���~�{�7L��7p��vA~������>]������ ��ł]����{��������)�\=+c��&�*�EX�Iks���v�4}�yw6MtS��ɲ|���$�V�uρ���+��+���;'�u��v���m�F�ם!$�v��ޮ����YzŒ	�owHSk��	��4���e0M&��_�t�d�W�����yR�Ume���A?,������!���z�4[ �%���ofy9�{v����Ă^퐒~5Y����]Dɀ}{nh�T���I����� '�*��$��,#]D�w%�$�v��H"�;��>��Gճ֏l���5��{�{����yE=e�zu79�y]d���oۯb�S���vf�Ez�*s}X|s%������_�J�s&����;/wͭƹ��,c"�pv�mr�s[��c��k�ڭۙ뮌�<n�'�m�֎�֮03�z�^:���dW���E��;ji���rOr��xj9���[��(�P/Wnt'qvu;g�	1����)�w^Dwnz���
�D��,�.�k���X����g���̜� &C�qw5Jխ7���Yۗ6��7,��r�e3x��k�.��ہ�S���	���<�k�j����~��N�4���u���{�b	Y�����2xې^9v,����",]t£I�LRa�\� @�������%Y-�I=[� $���'��{:7�|�vxxn���H6ˣR}��d�j��O��GE s��vg�	��]��]�vpM^e0^ �ak�����Eӛ�rM�\��?j�� �B��ʔ�����O�+��@H���X�2\��{ ���~]���Kw��s�A&�{���_��	���#��qU~!�������m�:��.�Ѹf�n|�93vL�<����磾�����-&.GD����  �U�ۄ�
���-�E��O잓�'�U����eN�
i��G`�*�iV���{{�177"����F�ɥ\��zf���礬G�x�ѩ�p%[O���۩�Oy��/�z���en�3��H�/��MV��	+���$�ֲ겸��5w����}֨!TZ4�X\�ВW^�?[�޵~����ѹ�%/��� m߷��~�C�SA�]�}�y����W�\D{=� ���Y���>�a��2�k����4��T`��	г=9�'�O���0�>��Oi.�����/��}� u�,�7p��hn�êl�E�gXuց"%{�W�����-�Z�wf�@��J�t
h!C���K�"� �K�o�_�A^�; �s���+��0G�n������	���ˤS���_˳�	�%�ڮf��ސBH$-��`�w�u�x�){jO,�7�o���'vQ���A��^�� ���X���w�c���aWS9�V��^^�}�F����ԉ�Ú��nL�mH=k�@�4g�/Rt*<8���Wvi*��k��_�
����Ho�� �{���H�g]QB��i�L:�e��R_���#�I�v��	 ���!?j����1;�$G�b�'���N�a�*N�ΐ�~5[�s�uؾ�ݓ�rŒ	�}�I�;������"�߶�suc\��%H۶�G`���yۜ[.��8z�u&�U�3w��[S��$�|gO; �G���$�*��O�����,�b���O���CwX�	4\�����q�oB����o�$����	5Y� %f:��`�\+k�7TS���Z��@j�� �:��������$���p�&�;���l�M��e2[�u��Ul��b��t�	��U�t�.�a��f�a����߳��垽�d�g�*����cF�ں�H�}��o�^�ԇV~k��G�~]��݊x�~�S���g�ʟ#}�	.�(PltS��.N�W_;�{��Y��^n�'���ݟ@@+�X��Ȫ�����b�F��0"!��(M����Buv�^ᶤ��3��s3���?�G���L/p�����@I]}b������t��U�g�d��EV��^���-�)�uE3`�_;����ϩ��;ν �I5]�! �����,ׅ����nׯހ���/E6BMp�wd�}W�d�ێSs=�����u+wĂ~5Y�?u__�+Eey�tU�U�}�0�*����@$z����B�����c�$�쐏a>�T�m�E0[����'�@+;�p�4��@�]�H $e_X�!wwI���3�6���/ia��ӫ�ȩ�T>kD[=���g����'V2���lֻ"Ŀ*Ur�2����� o����8�Y�\'Z��-u�1t�ܺM��kn�-���ҋ-�g��zoR���75c�1Yw`���5�B��狓�[��"[X�ܾ�B+���9�r��#vx�nB�`�ҵ�F6�80M�	h��������,ͩ�Kwc��5D�7� ��ݰ��g]���W����Bl��h�WNh:����Kh��J�'�������x�^�ŵr��\��z;`C	ЏU:!�[f�秵�9z ��4N�{�$�2§E0�c���C� �_;~'���'��v�;�姠�˟@A?U�%�~�h�e��i�%>Γ�@*�c��+V��!����ٟB	'����H%wwHEAB���{�Ez嶉lQLRb��>��`�I]�� $��]�)�Ź�� ����,�+{�.�3la(��৿M$%Pl� ���I$���  �U���0_�9IϽ�G�;��,��]\�N�t�&�T��x�g�CE���W/��X_�}[rłS�� '�U���G׀�~!�MSM����[��n3#��4�s�P���nlA�Rն�}�>�A�Т�-��ы �����H&�;d�������oK����q{��OĮ����$*tS�w{�AV�����=���I�j��� ��n3qFp���W���0Q�`�y��;ԧ:O�z��Vx�~O��=��.��bJ�Ӓ2Ľ���A��t��MVvϧ�N��e]M�&��av:y�h2�l4Ѹ��d�MV��I+�ٿ�����G���Y�0�"�wH	j��Jˍ�b�b��X=��}�x�V��	�������U{z@H'���7{��������!42qK�&����z	����n��AT�����;�Ă~����'���U.��噗��D�l�]��.�Yw[;kh̻U���m��lq����4��v���$�*���}��$���t��ы �x��4��-�}�H~���C�Ot�E�Т��]��ĀY��e^_�m̥�/I$��n�H$�,X'�uz�����{�	a{��Ya�N�0�̹6ă��Oę^�Ko���d?uܗU[bOf����VAa��r���u2��S���y{O���sG�&I ��'��	�����	�c4?l�@�{z�q�)�b���w܂��-׻�^{4<���
U�͛��6<�?M�@�i$�o�r�cy�)k�k���9Ԩ;��^-mS��eKo�w�ũh������?]����
ӭA3��[�W�����D;���r!o��;wR�OOq^mmk�ӛwi�]x%n��n��{}�U�{�r�c�Q��#hA,A6�.�Z�{���.��\����|˟-�7���l��<%{^-G�Ǜ�����h�F��*�v//Wmi�h�y��)�A�>�>3Pҁ�A�g0��̠�Y�{�)���7�^���T>>�Ƚ�Y �|���uΞ���6#�ܰ���>��L4s)�^+<V��ػ}���F�z�:G&p�S����ֽ�<.����jҋE�6�{H�jn�͇�Y|��ʼ$�dO����a��Cp\�v�^3�m��d�^�=Ǿ+�{�z{�]���Sv��8���Y��Y<i ���i�߮u���u����-��)����a�:+��K(�L�>�Vý��k,lFWg�x8kn��cW�Z�w����������~�c�녖)o=�Ý|}密�A��n��o�]�=����{�3�Sfz�K����K5-w��f�ɳ/F�ÚM��$om��l��^�o'0��u�^�R/7�&Q�:��ϛ~��?}��~����6"��#E"�,b
�	���E+Z�"�+�AG)DEE�1����UG��#Z��AH"6��U"( ��jUU`�2�05�iEJ�.��"�(,Q��-J+*(���QIlkikJ�[X���KlL.1���U�5�QTFb�J��1U�6�dX�("Ѣ6��Q�6��UIF�����
��$����b0DF*����RԶ��Ř�Ep��e*��U[l1n%��J�cR�Չ,c�J��mPk+T�EADDT����S��
�����YZ[[B���R�EQDFңh��0cmqja�(�V�("�5�J1���6!�()KV��J�)H[[PU1p*+�PQQ���j[U�QX(Ԥc���0R�Z6�A�ƪ��p�*ZT�JU���eŭ+J�KR��e�w�w�b�����|{��*ǻF�4�tJbO�vt˱���M��sݐ�A�q���H{�Ӗ:�`���U��e�e�آ���'Vw��H$��ۄ��f��Y�'�$�r��o{�C�[�۞���;~�p��!��ֵ��}���]�gd�8�<h�h5LТ ��K@M�EU�5�� �y�`��$��B���Y�}�n|}�6�'��������N�f�Qtj��wd����{���>L7^����A {\�"����[ԕ�AΠ�y�!���"�t�D�'�	������Vf�����Oy�,�E�wI��xd0§F�t#����0�y'
s�I ����I?��G���|,J�����
�]�������xh���\�QY3t�N������j^C[��u6+���>���ݞu�����}&a%w�\c��9f(3M7D�7�l��I���*6�w�2��{��ۛb����{d��VvޓΧ�Ճ�z���6��.:5�;��_o<��ͳ��� \�L��Of���t�e�=5w
b�b��.���v �o��pI"�;d1��rx���}k�;l��zhz���l�UE��{ �R
����1��73�BI��gl���g�u+�ڠ���D��A����w` ��p�m�ͮ�������?\��	$��C�Ol�)�HQtKrW�1oo��M^L�I �U��@H�r�X��`�R����c�Ě��aӪl��.�\#y��F�Qt��T@��΂|I���'��� �k�X�7�x/C����{&��Py*�9b�O�u�^ճ�aC���+(�_M�Ey�m��[t=���^�{N��~����9H��*����F�(^��C�.�vW�����v�1�r\m��dݻu�h��ckl�97�X�G=���ٹd��Њpv��t��R�����,�
,�A��3�mŪ�l�{���`)��?�6�|7ʹ���|��<�n�����c۶��gr��s�<�q$�O��+�h�94]��`�H�sʥ���gq��q8Ʒ1t��ڷgQɳc��1u�Ͱ�n^p���|����,N��I���������D�7����j��@$���]���*.�+�z�A��l���T)&.����c��7���,����^��V��>'��,YP�z`����s��◾E�YT)جޗ���8�E/eN�/���(]�Rs�đU�� ��v,��|�i&j���V2��c�>Y�)�w>'�nOA���eزI{�+Ǽn�}u�o�D�홰C��'�(�m4(�Kr��A?��\�׳h{fH�4{���̐}�ذ	��� �%2bTb#��`#��±d��A��`���\;XtoE�Z�m�xm�]?�{��l~��:�ˮ.M��O�v[�A$��������W����A����?+[����m�]�!%��v�ڙ[O
>dm�i���=炝���ު/޶:��de�M���.:Ӓ��ʵ�%J1?Xt���߰'f��ݬ-�)f�a�X�'�O~�0Ov��	{��߳�¢'��Џ1P��I0�t�_ǵ��!��n|H$X+�1|�~���$���Y?���&�^���-�ʡN@^o`=���-z�o��A?{�'��I����{p?ox-��_���p��G�I2��:*Į쐐	5Y�������7	�V�X
wu�?j��I|��:V�'*��4e�*�D$Q\��'��pЗh͑2�%l�#Ͷ�E�<�����z�!E�[�*�]�I5����Y�!��
��!C�CY��	���	���tY4:m�V�&τ�K�t۰�x߽�dE{�����5Y� �����;y�@�O=���]�[��!�m�]��[ݰ]�UƏn��"UܢГ��3�x�po�j�f�S}�<�x#�2#݉P)�.{���ũ�e�^��k'�ln#��(]�]
���S?|5��! j���AY��I0�t����7�g�� ���Uf���v�[xǧH����	2���m�
�����N������g�K���,�$�U��@I]/귪����u���n�9���c�/f�:��7eL�;;g��#=���TKC8yxQ��L��N�{$��MV{`�GWK��u� ����$�U��;	�S��dQl������h����t.h��޽$H]� $�tYW��Ax��]}�E�'�,e�n����$��сZ�%66����I��l��H�rłE�Xܢ��e�����$Ѣ�Z��e��X'�Uw$?F�/�~$=����ڹ,�oޕ�T}�q��cr�����ߞ����О�V���:�|��ެ�����Ź�P�<V|����Yܪ���$�쐏1BT4�RT�m�g���yݶ3���\�W�UrHH��A��C�x7������������;t��]G]K�>ˌ�'V��4_��=�6���=�ߟ�����6��O���˄�yۿ���C��꾭6S\�VL�$w;�d��Q�-UR�EgWK�'��)��6Ϟ���fgBA������!�t�w�h_���Bw�|�l�-��㿈 ��m�	xǖIvʹ��s��d�����~/�H�E��h��o{ܣ�D��]�w��v?	}��$�Uw����|l-=��O��lX%᱕�&)���{6@~U��{Ɨh�Ϗ��6X�A����|	'⫽�]^���J�u�G�K�s��aLyf�,ct��,�ѫu�ɽ���jHvt�x�9�3י{�b���������^���Q�Hx��Vg��an�zj�۷����n�ɞ�a��k�lxR�EwE�T�}�w.��	Ύ["M���UqYn��W��sѺ��j{!̝���X�y���av�xoj�b�xp��B�0Uqͺ''��aq=��,n���N�UxaB;:\�v����j���t<�`�l�c���qBѸ)e�5�w)]S)�on��j3sf�*�ux�;�3֞-�=�Ų�q��z��m�TC�F���TM�i�\w��Ă/}�s�~'�Uw�B����++�;,W�,�7�(_���4]2ʡN@r��Bj�ћ0[��m�A �{z�*�l��9 �L�[�Q�Z,��N�ͭ��^�� ������e�W?W�)vO��s;`�����N��)�2�[%��;�k��Q�]�h#��lB@$]��;��k�W����y�2k��	�����I�i���\��H�v��u����*/B�vH	�Uv􀓼����3-�,��~?O�/�"�e���lnܼ�a�r��f�ͷp�VcK�a�#����ڎ�"���4�pU��I*��A?���SR���O���� �Un�e�G"�A�2�����O��e�߉f�m^d���e�{e��y\�Z��j��'*�`��]������cЯ9OX�Vq[lP1ݾ�r�>f����{3sw�%{%��B������v,�C~n���w�|H�~áU �U
r�쐓��;vH$�U�k�F�����=���I ^݂H�wb�!h5��H���1JǺ�$��u��nޚ�$�$��	��ރ��Q�-�A��A��ϩ�Ȣ�-�K-�$���{�|U�nۺ풽�ּ�	 ���v,A7ݽ 3�g�a[�N9J�"�!g��q�9��^������[j��M�]q{;V�4h�n�]&)4�2�\~���ۿ� ��ސ�7ޭ`�nVU��BF�݋ ��7:LSI���ΐ�������y����m��d�}��C���\�vp����Lf��s�}����)�V޿;$o��p�~7V�z�)��^B|�/q���z/_��=6&�o+ufzM�4n�9��B�z��^��T�c�[:nL����Ϫ�3ە1��ܵ]_؏g����ذ	$_v�՜á:A�,��9}�2o����y��
}�I��*�լ˝Y��ݱCZ�</݌X$V�^ȚD4iSX��d�J�{`�o�}��ʿ{�7��]wb�$���H��d�������|��;Uv��I.m�8�r-͐G�R�us���m/��t��ߧ��wS�ټ��ы�y�m�H�v�2�2�|�Ykݞ�I7��'��t��T�
e���sg��oy��a�������	��{�b|IU��(Wz�<4��0���:LSI��Unl��IU��!�4�u��K	��f�ω��
��ϡ`��b�%6AL���~f|꼏�x�A���Uf��H;���wQ���~�=@�%��懮W�,���a��'��ӂ�혥�;c0��.J)q��=1zX�hH{7�����a�����'k�����'Bte�B���@���;v}����I����ݶ!%Wv������1���O�j<�C����X���Ub��ƭm�U�y!;vy�cƦe�XT�*)o�ΣĚD4iSp�� �{��$uuس��]=�~޹���B�ސ����CtТ�-�
ˎ��O*�?gJ�o�wv7�U���'� ��efz:��ٽ��Xt�ShS-5`�}���b�"�X+kś���$Uf��?uuز~�r�&(�Uvt��{r�^O�'�s'������	���6��Wo4�\�r�k�H� �]X>{�d�]��V���۽u���z�v,�k{z��A����d>��ʫ' ������nJ+d��}�y�-�$��W��/2d����5E�g�i�s�RyCtt{���)���s�<��n��(���I8�q��K��~[�9Ǉ��=�@`"�y�ҵ��瓵Y'�����*�۞kb<nz\*vMX�3؍�+R�cb`� ����H͹Y���8gN�I+��N8_?"b�,J����V�͗��=/�������;�+����;l�$Cn�',z��^�*˖��*$i{䟩XQ�*q��߈����g�Zn[|@��lى2wf��%�2/lS�*�ҝL��l��f��{!�w�����W���Vh�l����-�.n.Q%H�O�3e��l��kn^�齱k�x��0Y>Ȇ��ٳ�t�B���塴�͆�{Ks^���ww���o�k�xl9=g�9n1�N�W�K��uIem�'� m��O�
6玻�4�k`��#+�^\����	���[�/���y5G�ݥ�)��6@�ǐ���y/od�r��V}�����a�G.��Ef�/pZD�v+Ō���|��Qe�Z��g"v�Y}��]��SXD���Z=�t�ш q�x#�ﶰ��o<ؕ'%�l�v�IyCe���5�{|P�C�R@v��7���T��x�~��{����/Ow��;��{��dV,#�ywFzH��t���i��
�YBx�{d��-$��t[�{SJ�yz���qc}g^8+�0d�+S3wU���OF��=�=����2nS�l��?V��Eգ�R؍B�����ֵ�f1Qp�AP�j2���*P�(�KZ�X��B�p�Y���R�U��B�AD��+F-JT���E-Ç �iV�%ERڭ��
0kJ%VT�"�-�����+(5�%�X���J)l�Dm��Z�mQJ�JRŨ(�J���4��T��P��Q�R�-��X�+QR���(�Ĕ�
�bգj��4�Z��X�mAEV#E�����Dm��FʍK��*����U��m+lTm�� �me�JEm�ōAQ�RթmH�UH���"���QF��F�2�)lF�%J6�J�R��ѭ*ZږQ�ŭDX�R��iQm�KQ�[,mF�Q����eQQA�2��Q��m���VԶU��#JT����,X"[P[[QQ�F����)RڴmQ-h�*-�����*��A�m[j[X����TT�bڍ����Km�x��n0p��*;O��W�x��l۷V����*7!Żn�����E��>wϘ7ò�/y<��"����h�\l-�3�%g�[��nm��OYH�3H���Տt�]l�l�u�pi���:$]B:��)`�y�&���xccr�=S=���[���z0�
0X�8rd�r�Bp�k���x�t|���u��Ggv��m��@���֎�Z����k���W]��n7�u��h5����1N������YꠑlJ�pn��Cu�g��؏V옷lnNG ��7 p��Hvv��u�VOn�[v�˷��c3���F���q��<��W������tF�LGf���v��1���3���u��ۚݎs�'��Xb�}�trK�� k�&%#��f�v���u���vwVѸ�����	�\��̆�9�wf�tqn�ɼ�p�^˻�u���`vzh׉�T9��8����f7n힧v��.�۹�#�V>c���֖�������JN�*�qn[���չa�Mn���ܞ�\vv�3c�ƒ=2@�Ț%8q���4��a�^��1j��v��'J��-ϫ��m���M�S��p5�u\<��m����DJ�IoN�����R;a���;t��^Ie�݌�K܍kM��xs[mڌ�����o/��-��kjy�v��4��Y9���A�K��dw'k�Y;�ʧ*(��v��۝�<ku�)x�ڶ97:�ۛ�� ��pX�p�.1t�jۤ���e�Ѵ7D�>��]{Y;5��;B�-�Us����s��<wnW�y��غ��d����
uW�Zk����h�sRu�����e�.�.��XX5�!w;`�	;������B�v�,���Ц��ֻcYٹ�|t��z;okn���2�s��3����8�4�+������m�s��v����#�<hڏ.�Ż[�x�O9���(\u;��98�B�7\in��ۋ�m�uO3<��;|�|ş�\��j{��²7�����g:mj�\�=��5��k#WW\����F�,�����x��Q��sb,,��m�*u��\�\t�k/%=t\���ގ�Wlp��"��)��3��瓪8���v`�n���aŝ��2��U�ܧ|79���.|JV�M;�Gg<vՓ�6�T�m��t�'Q�]'Y��q��ۍ�]P��[kf·;�;���+7=�{E��.�kc>��t�C��=�k�zТ?i���	�i�U
~� �����}^�O������\��  �W�Œ�k+P&�e*T�Yϥ��׾�[�_��{��BI9]v,��뀓�G�g��k��}������nB��A �w��?���tO)3�s��A#knłA5����|�lR��2i�/s%]���sy��~>���$~���>����SޡxO���/�E�k�0�1E�Kf߉�������=>�n���|H{�b� ���>'�AU�۔B�m�X}ޗ[�E�h�k�N}����q�:��8��s8��vA(�<\/+�Z�6�N��)�
e�=�/�A��۟J����o�vg�0y��d����"�X���4�*�9���3���:��q���PÄQ�M�'��n�8n�v[�����p�N7�z�:��R�]=�
����[T{��#I���n]un�w�[&K�z�˖�����>"����;4[�)OaD{���U[��Y\��IUSw����A����OǴ�^���q~�=�G��!&���:�>n�[%�>+.3�}+
�Gd� ��넒	���>#�m��x��U�5�w����>'���U5J��L����B	��m��Ʒj���`��ْH5^ސH�۱dW���{�]�P���>>�-�D�g�aQ!:H3E���ͽ ��:��m�cɵ�ԻN��:}�w���㮒�I�|�w��*�z} �m��ߴeg{���I5Y�!f�k@��0��??W���c|��{�G�hSf�	5]�A^�ҋ���G3��8T��|��,��9}:	�����iU�����]�6z��E�k��0Z�f_���>���c�dw�6x�p鱊H��i���<q��h���L���	�74:Gj�|I?Y�>��H�v,�g�QI��&�+��=+��=պ�>�� ?�s�	 �M�[�j��]���;�2}6m�7E�,0�G`Oz{�u�S!�t	��#���`�M��%��MUG�^�ߵ��K/��6�/ Xq��m]��/k/F�]kV#���V0�mk��~�~�翹a�ڙ�Y{�N�,@���C2Tǡn�˪���	�;����H0�1D����I�?�9�m\�n�~�U;$�O�݋�_o\ �Q�I������Ic ��2��=��`�r���Ē7{�q�K^l�O�݋$���W�-%�*�)�v*u�1�v��Y��=�;�~%�oH�j���74�<;E!�}Y3��}��ԫ aS��;��z�=��hm�{%o�M�oE�QJ�Tݒu�G��3B�~k�@P|]����Z���F4�7�����~��/c�A*I��c��>$MW�d@�{��� �2m� ����]���&[U��:��};�9W�����t3f�=���m6ٗL?��^�[T{��j�7�O���;�b~&���{��{�\�>'�_��{`Xt�*h6M3f;܂V�l�H��/+�v	��{�@H"��� =W�̶OY��Bn�+�H0�1@��[�'�U��;���[�w=�ٿa5��	��l�j���Sd˫���9R��[7��D{'�� ��W�d�z�؆���yq��7=����\&���E��9Νp@>�[��^Uwm�%ogH	��j��b:���[��b�����W��t���H����҃4v�.&|���4\g�����t����_+�_����	�y�rx3ݚ�v�j{B~�y<>�N�M��,�	��i-ᤃ�7F���m�܀n|F��7n���6�NW[E�|��gs������zN�#u;��y��9��.��[<�/�C�h���n�]�u���U��]q�zs��S�E׎�n;n�.���K.l�orq��p;Jq�K��ԣ uOٳ�z(�[.�l&<!��[�\����	I��'cyT��E����vnL�qZx���a-S��	�$��l3���u�a������+C�U%I0�O_�O� �{�B	������Vx��s�q`t�H	��ݾ�����Xa��V]�,�^�o=�ͬ��/I �MW{d���WW����+D�a��s��~/�f�R��d�6c��  �u2I-b�/h�Y\���O�Wnτ���0O��+�a�b�l�WN��XG�����'���?���%ooJOսy�ݣ�,�z�!��,d��S.��Wgz�e�],����I� �z������*ϴ�Kk ��8U:��Re6�b�d0Ka�]�g���	:�W�x�iw�KqƎ{�����i��7��u�넃��?�$V��=0����m|rwl����$s��hlѪ��&����^��<(��+=�b�E� �9�ܢ��\K�d�G��>��ٹ�,S�� ���Ӷ˝�і{���� ��]���>�v�m�K��@A>�0�$����$�V�xw�u_�������ϋaҢ��
˦	$����G�-ۯW�G�� �W0�]���񯭚uJ��L�ƥ��n�*�a��,�W��nJ�$����IUݭ�wwT�&�|��a�_`W�Qa4��a^�~�EW{�xk�R���v���d��ސ�j��}=Z/a���a�S��:�[�<�ӕ�0G��=ۭ�ñ��[�7Y�d_a調�J�AL����� ����\�	 �U��V���;�G}�l?�_���4����Qi1N��N���TO�s�8N�VV�X$V{}p	5[���8�Y2���~׉��� ����j�_d�OƫݰBI�yy�oASx�D�גssۻ�(֜��s��z�>ܶ���z�2.כ���Y/h�fA/��3��dд&��4l{M��4Cۋ#j��uᄂ�{nH���!��c!�*,0܅e�ɢ�nB~�L��$�5Y퐐O�\��*�;��q����j�"{7 ��h�t�%Mɦo��A=]Cޥ�0$�{��ٞ�j�� ?�W?���T�Y�yX�_g���e��cvvl���Ʊ<�bm��ut7W�bغT�l���n��	�-��6��~$��O����W0�;���i���o���t�	�wdx�}U*d��vy�?� ���f���/?fX� �U��	'�+�K��Z|5oo��ۘR��Qi1N
ξߠ �z�Ă	e�\�S�18�X���I'�U۲O>a�u�^�ƨ�I���:�%H�Ly�~�s��= �H���+{���n�T�ZShm��s��P�j�$%׹�F;�u����#A��wq�����#'�c�~��/>�)^��;���ov��!�<62Q-Qb�r�L�~9]�s㛜r�Oz��ceU�^�l�}��2A�����v�}����F�4]$*���i��@�Kʶdy얱��j��p�{;5��=���~��ߵ.�ɦ{��s���}_2GWwHY�~���ʧ�W�$���o��d&K, �%yU��	��z����}�����?�=]�p��㢪��\�#�5�m0ESD�[[XOĞ��\'�M��<��о�W}��|��	���Ҷ�M���b���vw��^l�=�`�n�?~�;��V��V�t�!����<�������A��_�QT�n>��NJ��<�Ѭ�f�o���_�+/pW{���JM��U{�Ҭ�̸�@��M���`��]��=�_lWW����L_o��ne�x�c���.���Kr���+)Б>�X�Q� \�O ���Y�����h�$ �T�*0�A�l\��9z�pv.�
�	�;��8V�q�/X��2�p�9'�v�'��q��pdq�Ʈ��75)Fں�k�Mf��������'/O<��S��v�K��k�nyc����O,�Ւ��I_Yi�s{v�6�\%����x��a�m�km�;M)!�VxI�Lvq��bqʼ�Y�$��y��j:�ͺ�0�pu̻puŭ��g5��Wy��<��6���\����}���]����tY=}�$I]�˙����g�����VoH	 �U�ۢ���4̓΂��w���g�����t��A���>��#
�0Hˀ�2%��ED�u��@$�w����f�ךܫݾ����;[� $�UݰC��؅�d���L�g�ԱQî��꥟�� H^�A>�hf��]�͏xf{d�8���ePi1NO�͝$��P��݄o�О��^�O���BA��l��z����g��a�-�Si��	[תa���7gm��DH�ݞ{�u3w\3�!ɨy��J���k���}>5^� ������ӟ�G��h^ɲI��wt�8h��N�j�4����xר��y�wء"f]��M�l�����7�����]�1]� ]�I�fl���hf�ً��ڽ�9�d�;���3�kCo-��y�-߮�OĊ��=`][w�'���<'Ǭ/Zt�M��l˹�y�?�"�g{ר�0�˟'{o $�U��O��3w�o��A�)�W u���Ѩ:H�9W:�$���wt=;=c��{�$�+�:l�T�I��=�	#�;�+wE����]�.��$�wt�x�z�l7"��H����F�l �:�%���k�.#s��N�SmN)noY�a�w�����^���&����$ ���$��i��9��+$�|~���̊D�?�QT�t}/I8]f�������q����Zo��(�7&O��4_2��-SF�r�A�FWg\����<��{��UJ���L7;��sV��P8�y�&�*2��Pl�׌�/_9�ūw&�x@����kS�n�;���4�V�٤n�",f�� qn��U�|l�;�F9P�]�\+�wj��3!����'�궯/]�Yxb	I���/�킔��/���M��Ƹ!�ȳJ�7bP/,�*���}���Ԇ��07ݗ��C��{�|���v�����/P�V����J�+Lc�{��8V��W}�`��j��Mپ݊ovl� �z}��
�`t��̊g��Kt#��sƆ��΂s���o�^g�3|�ӂ���0_��w��V�笯8w�R���ueƒ�Ίh�/��%��2|n�[�g��{ޒ�jU/���/�E=�q_�+���7�W=�Ba�ss�Ty]�ɫn�7Y7,U��+�e�[�م��2.s|hC������}�_v�{�B�;��/���2[�<{'�L�K�4�J��O �]��s�_{���k�ܪ�|�]������Ѝ�g�7.בYy�����G�!6>iw�5z�7�Z;���o�Gz�]�rJ9k��V��2��ۋT��������m^�ZYs[cT`�nl��.<��׌��^��<������w�����՚���ۓ܎�����;�NIZ񻃫^���"O�l��oLڧ��:�2�����a�{�t������� J�qz���r�|�D�}�J�ٴ�$��ⳝ�ô ��I�e 񂁯��P~���Z�͙0�G��[KJYQ���j���ҕ���m)mm�e�UZƥm�m�E�Ej����,QE��V����ڴUb�h5F-�FնQ��j[YP�*5�,YR��TKQVVTJőek-Q�(*U��m��kT(���������)Qh�h�Z�ذ���5���ʴ�UUj����V��kiZVƪ��Zѱlil������[m�hƭ��6�(�YZR�E�-���D*�iZ�Q-+DVV�%��m%J�mRȣK-��cR��-#JV�%)F�1Z�ڢ�ֶ��X���
�[j�RЩJ��-��J5�h�֕�Z*���ګh[KZZ�[*XԴ��`�kP���Uke���E���[m(�*�Z�,�JХ��Q�*���-b�-l���Z4XĨ�*UUmm�Z�U�ѫU�E��IZ��Eh�[Pe*Qi[�Z%b+[-�J���Yl*�im�����j�eci? D7�$�|�$GWwHI|W�:i�m�l����oc�	u��]�p	���3��Y���:�d���!�h0�0jF�6@	'�UݰAY:.���UD��$��t
��A:�_��'�{�cZE:a$)����D�#����<	�8��[8J-���e�0�x��������"���&�m��~�\��I?*�t��fg���V�s-��Ǿ� �qڦi��iѧ 9}�p���a�r>u����$�q�� '�J��H2!��I����h�d�TU$�Ve�HO��U{� �{s�����,|H$y��!�VoO��E�(:��5H� )����y��v[��B��I �]�!$���X�_yw{~O=��d3U��js�g�ƾG!�j�Ό�}�����,���Yth>�+(����X��K��l��唯Yx�8�-�$�!��{e3-����#/�޹���t���la��_:����{�xW��@�2��,O�=g�{gh��plyv���J��#GsA���MZ��}�?�{d$��6c^�԰�;m�����5+L�4Bl��7g���I�4�5f�V��3o��H'�@U�t�	�0�"$DE����q"KŪ���a�F���쐀I͔� ���C��#׈��n I
��>�z���4[Id�TUë����x�*]�p'�&{$ �״$����\&�d6
!��"�h�e�5MR-���d�I�y������6oud�ݗ	$z��Y ��z}A�U�g{,�?8e�=�o(:8��<����z-X�'s�u��C>I���*�[���<�8�!Դw�����}�^�T�.��R'M(�=��7!۲A2Ap���G<9�\:��kqG=��w7���OM����8ٮ^ڛF�g�C��O�f/n������i��ίGh# �^z8�0�&�R�p<�ptm��8خ�լ��W��J��ϒa���ه��������[d���2;�c��j㱂�	��&��%�;���G�����X��k���S�8l����s�ݰ]���m۔�&X��F�h�6;7m�.Į�ݫ���c����i�4�T�t���WQ-�t�`��M����I������
R>�;����z��L~82�4B�5 ���~6|Ϫ�+�֌�;��G���'���\$ڥ���K���*�Ӣ�dӤݟ>�`�����	"%tS;��������:�l_Ğ�z�'�/W�j�$çF����������`�?�����J�ޘ^`���$}�,|L�a���)QTS�w�rB~!W��G�ݜoǼ��}b�Ă}�@H'⫷��j���n�> ����A�i%D��������e�1*¹mk�����]m���k�����}����j����[Z��I����HU��x6wq�B�Ԗ���?H��d뭢[��M_�˝ ֬���x{3���^���CN?w/�O&'��RKR3�6�n�uW�.z��uE�{�Gj��v�����p����	�ѣخ�d3��A$�-��	WoH	¶!{y:�ӢÙ�A:��e�h0�2jO�<͂Uwl��>�=yu���=�?e��[�"]`�Ti�E�i�oB��E�~��N�ǫ�� }�x��{�L�-)�Q��Gnΐ/�I��$çF��{�a�k6��L�T~�Ϻ`����>$�Uv쀓^�`�^AU��?.����7~����ǳ�I,H�qWAaT�û��ͱh�m�{��~���nG�o���$�^�@!^�g��b�v�Jޞ�AU���/�D���:)� 9o��H&�x4��^i��_ �[�	�vذ�����z�����d���[��MX.\��^�w�a��ʸx�=m�wl�׼��'��"�����8���F�]ߦm��:%��f��~���B��;{eb[���^ނM{�Œ~���4B�5d�F[��4�h��4<�'Ђ+w��~$W^��v�ܗ�3�\pz�ސ�.�JT)�E�[���j���I���>+|Zoh��&L�����y� �M��@�$���	�j�6�6&RK|�-D:K?��' q�x�(v�ާA��aӣN~�c����	��7��.c>��ס��H:��X$d4V�E*(Ra������Wg�oD�Ҷ����b� �M넕�eCգΏ��D7�����j������v	'����_�������~��Tސd�5�������9j2�SW�~#����A2�z}	;��}���e�Bdճ��0���p_C��6��{��UF���w�9�H��b�Y�^����]຿�ު��n�B�o,X'^(�:�MH)�:B	Uݲr~�~F���;l��e���D��'Đ����zп^��g|n����vܨV��i؃�9fѭ����;v
܃;����7�*�"�-�o���vA �N��I�[�>N{ŝ�~���m�d�Ot�&^ihSi&:4�/�'ЃOR�U��y:^�����=�$*�t�^5��?SP%y���+�"�)0݁�� $����ăL]#Z��rYPx�>���*��!�l�,'T]E7!��s5��]w��Vm
o^�$�B��3�l7s���e=�Vz����Id�u����N��s� �s�Xqͬ�W��7~A���@H$���>νb̦�½�����Ǜ����xe�m�E�4{��[�G�Gw�S�+<L^z�w��<�\}�tz.����*�-,�&�����k۲{��7�{؁��_ֹ��Ӷ�p�*)��p�%t�Vrv	9�z���y�ە��G�RB[8�ع�T�l�-�t]ҽDc�.pt��
�W����b���α��r���v��.7Ȼ�v�����ӭ�ʦ��,�r'n�y���ӡ;xN�(��v�0x.���Fa�<���a�*\l'V�ݝ�F��<�n^w�W<�\��<v�^Fۡ�ws�È�؇��+��`�t���
��`;���xW;Ob�I0�����i����{` `5ݰA$�^ذ}�y�</Ɗ��=w�! ����%�F�"�-�n���v	95�E�Ǘo�^߾ ���� I9׶���^��h3/�
m'EӣN����	 �^�$�<7���ϯ�  ����|Fu��Y4U�n���tmd<��e�s��g�A'6��'��7��r�<��`�ނ�����uE�tSr�Gd}S:����!��Ƽ��:BA?{olY?:���м��3���I��MP���R]�9��3��Z�uX�q�{v3jw�vx�����6�6�6����X��_;$�=��#\�]^"�op��>=��,٠��l �Qhկ9�=�6 �8#�5��]�s���Σ�NN����9.�����=G݀o=����n,�4�_MY&�=7V.�̓�u�r�a��h�s�$���H���! ���&�%���^��\��Ѡ[%�-�=/X���}�qp s(T̥uy���`׶� G;����w��5AST�P��+;�l~��L��I%;��$�K����)7�i/'3�xIp�IN�\1%��%���*�L9qm��3H��l]��*'r����7�ကE���0��]�A�^�C�T�ص��A�Rm�I��`�[tt��%s�����j�K��m��\�߿�f���:��)��W{�$J	z_�`�@U��h<��o29AnjA]��(Z��&	�L�̓�v�3���/���9~ݬʿ �>�wۙ�Uv�l�����əܯF�7�~�� ��)��A����
�!�I��q"za�aܓ�Y��g�d��3�i���6�#�vG4 ��v{mS�6^���)z]Iy���B2�^��Oz*�.{��u{i��

j��C�w�������ϱRo�	o��A�H�K�-�d����ܺ��so�$�gs� [�6� ]����K��P') ���f,3]b�UT!T�VwZ���;�j���3�q����"+|���� ����� �u�g<�������߿�o�74j%�K�vb�on����c��J�v|�s�7S1�=���￿~�m�9�2��o�s>�JI�mόI$��]�nWDĂ�DF��^>�ϰ��*��1�y1ͣMPb�n3ձ߂H%�_�ٯp�c̾��$I/��D��Mv`!j��\�T���N��9=T�t�m��,��>1$�Κ�$J�=��B���x�D^�!���Lw�m�ɪi*^��f�����>g��@���D4�}����Wx �{�Ϫm&�S�u�D�~��%�׃�I������i3'a��쓷~����gm<˩��ƻ�s*n��^#�b�/���x���p��?a'�� �}m�2�aR-��p�޻�D����^,=~n�����=�(����g\1$��阕nzWh�
'(�_7��^Mq\I��m�iu۝��w'FQۙ�5��baO��{bT�R@Q�
��pπA���!���}���u}0�R�/l���M�g�f}(��M%J�l����ې��=a���zv^ bI�l넘 ;/�1a e��^�{O��u��a��K��h�Jjbj�4OnS`|�<��0bI�73K����pq>	oMvI�/��}ٟb@��]mPM�Cm'9r\�3muj	h"'uհ s�nf _$�o������^+(��d�I�gx�m�ɪi**���8�	7�pP�4*�vɧ��	0$�K���	�� ����8-_�x�g������yNx�^�(=G\v�_�P�|e١=)n�t�D��n�]3�̵f�jG���ssO��f�,�)�S=�=�������7}�?o�I\�<
O����<��M�u)W��O�y�R�+[�fF�lT��Lu���$y�/u���r沉��Evm~�L�{�y�*�l����ܼ}��=�캢��sA�kv��ԄD�@���u��� �����=q��O�e:M���t���u1���j�����Z6���w�q��xe(�1��u<�9o��/а��_���՜��FIu��{��A^R>��#�NI�`LMl�^�{L�UԸ�V��F)GH\���,v׽�6�M��w�'0�> �/��#'{��E����h����3�%���§�|����׫�w²6����wb��k]ϩ�'�wy��ܞ���n８��F���z�`�n��S�I8a�{�sk��^� �s�MN��x>��p| �|(��S�/О���G�_�������b>��b�`�)1o�\.ʼ^���o��Ř��b=9�tf��1�f��E3�h��D�p��{[8��ebT�S94����x70D�u�V�Ƭ��_Br\��n��*W�ܛ3Ƚ�@��-C�{��OU��g�m����= ��sΓ`�ܹ7��o������q�
`^sW��7J���^g҂�o�$��ȧ�I���f 	ݹ������s�!���>��pu��^힤:y�k���;���֛�^~�}>��m���*���F֭Q�U,Dh�QjQV4��*�PQm�l�D���m���V�[J��iiV2�YR��ڭ�D�KK[UVڔ�E�h�T�4DiV5%)KiU�k(�(���(��Ѣ%�Z#J�4*�B�m�5�V�������mU-P�m��hYRֶ�
��ZU-��ET�E-��Ш�Q�j�
%��Z�VRբ%�U�Q�V��aQh���ڕ�6��J�5�ұ��,R��m��j�J���T�l�Z*��VԥK����������h�Z��*��E��V����B�J%-*Q[JR���Q-��Z5)DK)m�� ���UF�[m*,T�Z5+m(Z[AiiK)Z�h�����
��b�T����#Qb�F��-A�ԭ�ZZ�A�Rլl*�)k[E+YRU���R�b��/��߿��oߎt]���{��;]�ŻOu�9�
��q���i��F�u�"um��싻�<F��6��xy�*�6Ck;a��<�7X�����e���5r����ӭƸ�]���u]GmÁ#v�^��(�'�i��]k��}6��9�sŻk�[`<�]�l�a=�R��oC�Yv�[B��:�s�vsq,�wn.3����+vK�r�N1�d���L��w\��/U�Ϥ�&��{ϵ�<]�RI�>�Z���N��Zݛ��z�t=�l�3�3�{��vg�0yR{ ���3����ӶM���vT�R����]��Mn�gc��v���j�� q��	�y^ئ��s۞	��w��T�2��5��τ��n`-e��:��Q�H��x��{$$�l���6�v�c5�.��d3����s����{��(ڲ���(;���[�.y\�܇D.��gͰEÍ��v�1���}��p�i\�kx�:�1��t:2X�FD.��v�1���Ϝ�x뀚��ݍ�9:؋��{��+�s�h���ϱ����Y��K�cv_]���l��%�֎7BN��^G\q�M�uÜ/��H쭫�nŃX�=o&i���t��[5u�:�`�{rf���g��Ǭ'7P=�s�st0���j�vSe���a�֢9��<�	ǧ�c�E������l�TgGO^��&��*�'=�n;&����z7n�g���{�Ll�ȝX�V�w�T���7Tv��&��Κ��$��Nw!��$6�����^;Z4-��r�uom.�,���ݎM��GsE��C�OF����N�[]u����=�Ŭ��S�{�a܅�x�t5�Đ�UN��ֺ#[3Ggv�q��s�:Nztv\\v��kSa�`{i��\��B���op�ۚ�83X�kմP�ySKBn���x���7]�6���7��0\�q�������r������s[ū�k��mX�ƪ�T��9�C4���\ݗ=�db۫v���w�g�s����P�6���qx䭸υ�n�xv�S��z���ٷ��ZMi�ݏ]���C�n�5m�eݺ�B�v����Vc�G�:��i��2Gh��qmD�����N^�?9�ɟ�V�+�����`jH5���n'����Z����
�L�&N���w�����Yr����e�l
�oK�����Xt�z�a��뛃-��;U��@ٓ.�g����`3���ؔy2N��c��??M��J@�J�U^����� ������PI7���4T׷H����%4̄�TS��I5 K/z�0�8��Ʀ��~j;z��� ���2#&��Y0%��&]:ݳ��˳�.�Fx*bBIQU���c�@W�چ $���"�3����D�I$��~�RAS�A>�gc	k)�A�ti�������"*6ڝk&k) ��<�� ��i����k�q��*#�#kք�\�73���ڠ��e�tK�/ �ڷ�`�-B����b�{٘���]�nS{���u�~�;'���Ͽ��VB<�.Ǔq�;��rogf�*Ѹ����nIv.�t�w����c���٣|��}y٘  �޷۹nt�}�=����vfb($�M��f}Q�����1U������	*�2$�R�����਷��/=�^�_W��ǲ�-�]���e鴯+����M�:�I
ŧ�#. �h*?z�������s[_��K�Q���� ^�V�Dw�*�$���iD�=�}�٠cHl��h2��� H7ݕl b��D�']V� >*��6@]��q���my��%���{����;���Ֆ��"�D_�ڶ����i �����Ui�Bz]o�<��E��
����6����I$�����Ϳ#��~��V�D�� 9��İ��c�e}�c�{쯈ꦘ4�o�L�WA�����C�e�@�;�t3˭����:���������:����(�O�e�g�|��l"������ޗ��7Hv�0�6��\CH�ˆ$�g�N�����B�ݓ�H#:�Kڬɫ���:���1  Kw��?�����O�����v��%V�MQN�ePu'�w��$ĺ?s� g�U��[(qݶ��꒗���{�!��{�	���dU���f�i~9��,t�rҡo=Y������R���0��m����L�;��+;��&$�I��1,�w�Y�4�&�T�AY�w<9�Ϭ�ܷ�����	����@�ݙ�|5�UflCZ���ZK��p�:��j�"�P-�.|��ݘ��k�o�x����Қ׸]�<v�o�F ��sM2=Y�d0}�\)"C��P���"�4Ƚ7/l��d=C��&�N���i���������i�뛚��'�W� ou�  M{�m��:oժ��^��r�$>��gؑ��J�D�`)9S�f\ �=:z�b�s&��z� ���0 >&�Zi���Q���bw���RKs�����d�H%8'ۏ��]�� 1V�;�=�����ٟaA]��`��F�tRa��5'˷���8�v:��� v��ϰ5�j� ;u���W�E2��t���sFi:�ܲt^�EZE�J���ݮ��Z��b���R�^�L��ݢƊ9�/��W�_����Y׏?/�lKĜ���$��(ݘH&�F�
��W�o�հߢ<��z�+ޠ�ǭ� ^�̀;����f-��nCj�I�m�~%*-R
%ָ�k�]W�<��^��>�\�6��=߿[��y�0�e�����0b$�{�>0���1�O6�SFS�f, �M{Zm!��'���0�0�rʮ��K0ku�������k�����W$��{��衴����C+��M�Z��Xcyo�`m�[� d8���=���ɥ��f{�D	[�?��}p���wx��e�l��J��c����%�Uä ^wZ��u��`$Ȟ{�4m�|��t��I*�F >΂D��*�&j�W��	�$�'����1�^W
�=71'��:մ�f�ۆ �{ىa/'4GsóSܳ[~	/dZ�G�FϨ=�ux�s�yy�c\��8n��y�E��������n�ld�S�D�^���,7���]F ��K[�<v2nB��n��]v��M�g6�v���q��s���D��Vk��-�m�H�u��Y�.7Sxܹ�5{���ӳ7���}���m�e]n��@��s�P����>�����3Ã�7'7d����L
랞��m��-�<��Ɏ�s�V�.�#-ݘ��v�l��e���glp����`{m����v�D�[M���H���5��(�>m�����+q"������n;��ۏO���߿��@�d����]�n�Do��� �{٘��\��W�ej2��?�z��0��6��
+l��_��8O����W���gu�C��=��ကD����@��sg{}�E��|�6�)�ۻЪ����>	���` p���G���$�޾�I�$>U�{!�p�SZRQJJr�A����Y/�*�{��9d4m>�����5LF����+v�1o�I�2�6Jl%B@�/��� 5�j��X{Y� c��0�I|���ϱM>�D���c�gs�'Y�[<�q t�lnr�I��8�06�m*&��E纎�¡I�٠��]�Y"�A�����Mvڶ�쬨�9�"�m����\�I,wݐ�-�ZT)�N������P��WW��;S�Y��bOY����V��/z��#s�d�샺F�����N��w��d��{�v�)��Lՙ�0�/Wצ�<�p��͗wX��'o��N:���#���}٘�]�\C�����;�� ����H��TT��^�c���ݷ �n�h�&��]��I>\�3�E�ʟl����4ۦ��n�X�Aͬ�]Ô���˿s� 
ku�����x�B��Fv�������?Nj�M�X��K$�I=[[z)k�&��S��|�~��@�5���0�����K��_ z^߳����Mh��W`2	�k�g����N���,�z�W'����N����z�t�I6Q�
��٘�I%O����T�\�� �=w��{��������a��I�٠ԁu��(>
�o�𻋥�����{���	��!3��r��>H�U������snk�Y�w���J�$l+;�����ڠ@�t��GT|/3�2�z����WO׍�C�0��ʬ<Rd� W-�פ)�
(�����M���Vyy߶�v����)d�2�M�+շ��H M{�i� '���+"L�=12J.��z��T3�P��m�w/�'�z�����s�:�y��]�X��G�x�I-��$H����6�)�M�P��D@�*�^%�q��3���퀮��l"'�m�� �~��<N�{��W��~���S�+w#�N2�vk`����kqk�+��;�C+��2�b�������;����A��چ ��;m����٘�5�k��i�`�q��@%�;�x���� ��� ��;���'Вh��W]��%���w�p��~�_r�$���f, A�u3�5��k>L>����b�R6h5 ^��'���~�$�
rm�ן�uc�����9@u_�3,ػȊ	SQ%P6���}3�w�2=�Q޶�� �_�3���9J����)�?��O��a�x�^�{�oDs{;7��q�RZ�id���Zxx�Lw��et�L�ǅ��{�CY
�	y.������o�~�.Z�q%�:�J&
MO��J�@�Ը�{��$������P�N�J�� :��3� �z���f�}l�>������������d�/C�ݮ�txc��QݝH�E�͛�Cۮ���:������a��ꨚ��'��`U� 
z���=���W�n�Nn�vW�Q0$�\�ۙ�$g"��S`8�Ys,\J��QΪ���v�TGU���������sw�>�*��t��w��)�T�R&b����XD'���b�3��i^s� �:�u�� ��i�~��6O���]krr�`w�D���$�J�t�eu{eD��Pg��,T�L�Ng�I�ד+D�IgDNw^��� �=����m��Q�l:�6LH���������[���o�5��f�F���ۙ]n�2���Fן~'W���<;B�
���3W����wх��<��Z�q*&56q�V�:�]�`8�nwf�/li�۶ vzݙ��8��9v9t��)/��V�K��bt�9�;Nt�۱���V+��uQ<�{��Hw`#�a6r���/�rV%��ޑ������|�2�g9�|7ڞ�WRќ:�=Z��v7ph��h��[w��|�S�ob�t&���&�S� �C\\i�x�ㇲcۗS�JM˞݃OF�[M�و�fisRq	r��;,mx-v�I;>x���D�e�H�C�!.�TmK����3�I"j�m�b�OO��@n������;�%s{31���bD�/{��t�f�u�行�j:b/������H	�l �(s�l�`Kz\b�"��Sȥ�φ$�v��Jlɧ	e̱d��7m� �=+�ֶ�^����4�lY0$�:�ʁ.]�N6]SE&ª7���7�Σ���-)��,���=�X #���c��
써1[n�}2	�N�L�&�͖��k�F��~�e˲��Eu�Cw� �X�zT�"R�{٘�}rj�׹����#��}}��lpݞ.Qn��cGD�7� #��gW�Qh�U�C��iH�4s�SuٴH#�f۠A�{v�u�mz򉺞�u����sM|���r�VD9�(��p6�����d'�e�մ~�\�榼rr7.�7�1mBVg����X�/��������s�v��[������������ڰ�F������;'j�O�o��$�%�;�Z�>G;���I}0^{����}������M*UU%S�N��� ʾן`Co{M
}�/mz1~I$��v�$���vC���ki&�,��VL��]{پ�69���<7-��*�s1 �*�mo�u��}>�nX�ވ�l���M�TdU����JI��{/&�z����倀F��c��
�� �Ku=��G�6Mn�U4i�%�Cz.����D;`74���\�l��Tc���{��&���e���m��$�w %U��h*�2�,��۝@ ��f%��kQ((��(m_u�`xVv�o�U�n�_r���K�fN]�6A�qO��:� ^�$�52J��.����3��*�m�DO��G�\N�	>����w�ޢ�凒w��d�����=�\�xx3���|g�{N�og|��fT}}TȧO�!w�k��B��{���v�G(�l�ٖ{��M�Dy`�ӆ����۹noZ���d"�ǵz*P������W����Z}V��d7�0�r�T{5������sU7��M��Z]t�^��R�;@=�{�R����[�����k4�Ԭ���e�K��M]h��զ���ٹ���6�2X��"�\َ�q����=��G�}���y,�ތ�ئ������8��M�iGM��h��3F̏�_3=����Qs��)�t/H/����w7�oS��&��I�^�Q=�oA��NH5�����JY��x��z��<�sx�zh�Q�Y��]������{�|}���&N��{�%��%%T�R{Z�����ox�t��R�-�:�i���
�����Z+'�$��lJ�5��Z�fɒv�e|��16��N�5� ��T%z��Ǖ���B+2*�'p��ṱkһ|c�9#��%C�17�'a�Qm�h��_��Ӆy��:�J􀒇}h��9�qI��Ё-�o�ܞ���)�9}ܳ�8?%��i2�7}��u}�8\�qn�a�ԎG0p�3��d-�wt����}e穯w���e>���o??t�e�Ug4[�Ιq��K��-����w�c��A��¿*w�����H�O�۵~�����P��pH���{/��^��;�<�y�����}��mc�ɹ���l����(�EYKj()F4��c[U*�T�%B�-*,��-Q���5�am��R��,QAAd��Z2R�UkkDaie���h-,��-��VVQ �ڌQAR��IY�E+PmiP�YR֢�����Qjm-i��Z�VUB�5e��*�b0���[EE"�ʋD
��F�[H�m�T*J�R�ڢ���J1U�bTZ����E�j��1�,h[E�`��b�-V�ږ���EX+��h-QPD�
�R�UeH�j"���PZ�EDcH�eE*EU�B���X,�[dP�J!Z��ڊ�(V-b�d��)kd�
0�b�dX�V��ih(*���X+lP+-����b�Q
��T�-�}
>�V��  =W��� U��`9A�L0ۤܨb�
��=V����s�ń@���i�T�\״�Yi�-[ǫ�l$����C�úkd����_%M��8�H���T���R���.���� ���i�A�uۢz����q�Oq؛�۪t�=�������=;]��=�ʓ�+�c�f�؇��F�4v�"v����1}�>��b�� ����� uO����gmHJ��b��0b)$��$J�>�]#D����R.�q� ��J��y��=>��op ��	K�:��&|��������ہ�z.�(�PQ@P�g>� 6�u�@�����7e�_�l��G��^������`}*�EDJ�IF�m�p.~�c	'R~I%Nm�H�w\�U�����-�����lKw�;���TE���HC�h���P[�w�6���9q�P�pY�8e�w���j�\��M�7u���C�$�ېH���M�6�m�n�W��@���x��;=��hWW������w\�?�:��1`_��kʅ+�����ۏ�g�i���vy���c�gt�0��m��vu�]h�ur*ݧ����O� ���~=�T�.	�n�I�s���	^����߲�_{�4� [S�rÏyB��-��xR�T��L��)�����ww+�� ''y�DC:��3 'r��ʮ���p\�H�4��jD�v7D@W�y���U>��{���lG�N�k��#��s0>��-b�)T�ϯ�zg�tc���A�yn�����@ �]|�J���v�x܈NM����J�I1**���k��0b$��.=J�^�KwT���DG���0���m4���Κ���e��P7}��UK�ӛ�|vz� bE8�S��s�<��x�<z������r�y;�R�d��h����o.yJW�F�X4i|E?�^��c��h[�v�P�m�k����96���m�v�U�u����e�V�	���L��h6n��
�.뇳<71�&��-f8�z��޷R�l�<�+ۂ�L���vκ�dm������ّ�{qum���]�̄�ۧ��i��g;�6�.˝�^:]��h�.�%�l&Un�9\ݼ 99�[�x9����m���U�ݎ�փ�)v�=�;-�����G<���<��ѵV}.~~��m:i�j�n�{\���	$����0 �]ͦ�}Y�t� ��gNϯi�����}��8(*h�*��?��2�y*fǪ���W땷�RA��sy��]ͫ���1_�����}�Ɠ�fQ�[A�Ho7�L� ��nDG��zc��d������D�;���I@'� �+��#5IO�a��	��N˵_U �$�Uw�1K�.|�	 ��bf��[x��<3w�I�:�	�tnL�%��%�~��^�o���R)��ژ��k�������[|��0��kA���Z�U���pH^�n�%�,ݖ9���u<�[O[=����5Z�0Y�Ww�}~����G}_~�f, ��چ ^�c@��y��m`�1�d��I=����v��-4���|����v"p��9	Ov�B1{F{=b�mͻ����Y���nl'< �� N�����N����V�}�c��>���Z#%��ʟA���.G���wؒD���	>H��Ϣ�~&	���q~��zKA�� Y.h�&�,i�e�q ul��A�+9�P�\�� ����h:�=c@���Ec	6�Tʪ2���	�'\��""yx�� :�����H����ۚ�����Eu�M���*I����I����F|�5��!��JƳ+�^>�m���s����X/^#;d�՝�AQҤ�H�l��3HQl��ݻ΋��ΕSP�Q�u�T��cIf10s�|xsr[���(����`6�u�� A=~��ਫ�>�=���6��i� T��b@P�IV�F� �N\O�ۙ��z�d�n�z�m�$���]�$��~�阉$䧛0f�<�೾V7�n��tԕNZ'��D@��y���=C�S�j�
��y��+S����5��^-�I�����0n�����=ш-�>��px4���V��x��n�S�W� 2���@O_�32;eșN���MDJ��{��,Wt��l�`6�v� 	�|=�֚�<oRyei�%9N�&u{���e�TҪ0�9��b%%]��39�����z7�Ԑ�O� ���,  ���b�e9�R���6��h�N�U:�a#B���X��ۃ��Uț=�ɍ�<7�K���������\7:뚾m{�4I5��!ĉC��H��)���^�79�_�|'�{3�Db�(�L��ĳ�,\	Z�L��)����� ��7� Oki����g�_��/w�Ph����e����!В*ݗ>0�|қg�m�����$�	��HN|�U� �.,n��S��:t���X�Ffx���V7�	�fL��� ������^μ�b����K|�Y�OY�k1ȥ����Ad�����o�8��I�g�������:�Uׄ%�;=��0�s���:��^�d8p�T4��M|i��0�yn u�����׽���w2ȼ�x�Ю��y�D���d���夛�����}���4�@��2A�=���}��Og����n��r�����u���ݹpZU3A3���f%��=�چ ��]@����Fo�h�^5y�o؊�$k�,A����QT�j�~�]��켚�&���=��{�M�t���A[ݛ�,�3 �ɶ�ٺ�;��TD�Q0T����m(`i *]�t]P��)߫n�@��i� >��s��Iע)I:�J�"��v�}��m�'�{��w�̷ @V��'�ݚvv���2�r�K]y�'�-O�]2��:t��1�t r��si��%̠'�l�U��9 =~��y^m���Y=ط��5��8P��
�Y�;�.�_o��,�\cږI�w{���ߕE��'l;^��jG�l�\�<�����۵Ůp������.��1�Xմ�ͻq�R���u��0�����cW�m[����N��-�����u�95�jq�n{t�g���7h�tq�q�cBl]n璭�}����k���@�۶�^.�!Бɪ�&�͹�N<nZ�ٟ.�d͹�F�.����;�^�3�VIh�����W����+���Ѥ4U���͵u�]'lp�ua�k�9��-n�Ep;)�Trr�<Y��[}�~���&=�/���4��0 �=�興>��vf ��>����~����o`��I �]҉�����&XuM*� X�;0I-���}�g<�e��%�"Mu��E���<���Vg�}�y��QT����w�� '����� V�#!��!J��,�
zw��=~��=���K�)��ӥq,��ֹ���u�cr�A�/��A�D
v�s0"O_5:�G^���vO�* ���ܻ	9��@�U%LDU;i���X �N�ۆf�rD��
�r�����X@�u�E��Lv��t�b��j�l׳�]��E��5���gk,9�.
g��b�Ş�ɜk���n��I��^k�(ĉy~��5��h&߮(�^��8����=�Z V߷3�lt�����>�����r����
'��d͸�b�Ӊ"j4o �u;\M]���b-��Х�wS�@���[ݜ�����;<�:���lSҲ�� z�s1 �&��A&k���ĸK�vV���N��L�Lų*�s>�A5�mC w{�~u��>	_�vf"JT���9�:��Q�b�5p'�6�T56���� ���6�	��9�#t?yt��3��O���ax��mWu��� �=�1]�I�/<z3��~o> ��֚d������n!�B+D�{��l$�j�������45g��ݴZ�#/=9��J�r�=���������(�[��+����I4�n�I.u�/��'Cv��d$�
�l.3Mm۪t)�Mۊ�N��Bڽ{P���W��, ]�6 �}�b"SB���v`�/{d���ذ�ڕUT�
J��	��V��n��A}u�t���Y�p^�Yeh���d�`��n�h��2x�m"�y2:����J��bG�u��M]��U����j}N���ܧ����	����"J��(�:����)2êj��9Nt�)�Jbo<�"c~ s���"�;�Z�������z��j ��i�S�Z��&���\^�ޓ�IW_lϱsݞ���,�M�4��>�- ����n4��v�=��8-�W�TU5@�Wi�V��8����;jp#��M^x4h�}~s�gtꨙ&��@�֯�A�{��@�@O^�f%��0����;��|�� �"�X�u�I�i��E�E�ܸ����ľ��fޱױߒ�|�uN�@���n`�PIf�fs�.���+��V`�)�����
mSq���D�Y{��$�dO�>����y��_�0m�- =~��2<t����B���	X��5�c'Q�EK�<��^�h�Wշ��ĉAs���oi�<8z�V��]��u{\�}�:ŉ^��g��k?�=��7G�n�0'�Gi)����QN��tolw�����6����ǑD����XB��L�3#W���A�}j�fku?�y��` 	���0���֬�Iff��-Ѥ��JҠ�"Ca'TM{C��-��8�Ӹu�y�W�EN�m��w�������&iTR�G�}>n@�z���F >�i�3aq�����D09{��|&��S��N��w���xGfI�Ns;X���]���p���I>$�Q�z�d/����}�Բ}��4�J֩�2T��U;i}ۘ�>��A{��s��:���9�u >��q�U�M0\Y�Ҧ�f�MQT�<S��U{�׉�o�D���	8%�|ӈi ����K�Y�/�D��v�>�O��4�e5��_���ކ|�v����˸Ɉ�]�vf m��h��m�y�8վ����$��	!I����$��	!I���$ I?�	!I`IM��$����$��	!I��B���$�	'��$��$ I,	!I���$�RB����$��BH@��	!I�HIO�$ I9H@���PVI��d�z������@���y�d���X��                        �        >� �      F�    ��|�H�DTRB�J*J �J(�@�*�(�
���*H �S�el���R��� C�`��/6��L�]��D8����sF�P��S��I�^���v�� �例�����)z�t%�S�>�92J֓��e+�
�R�<��Yu�����몘
 �P�*�I$*�)%D�U�ϭ^�w�:ҋ`�{wz(x2t2�{�E;׋��{n]8E� �JMj����ꮱ�S�.����g�.����������  � }�BED�
���	�>��Ӣ�Ϩ"v���[�����������5U�� �uIw@ ����@��    ����b����y)\�U:o���v��,���8-�\�]C���l��6GP
   >�E
�U"U��:�J��Z^�.gv%]�U+�I����=`��S�t�`�퇚 �� ���1�/cJ���<u�QݏG��.m�e�`�l��̈́�ڒ�h�� +_|��O��J�U�^}Q�iY����У��w�'���z�c�\�twi�y%��wwzc�@ �UH�y붥�}p'=��R����G�M�*��\5���`����<�W�      ��h��J0 &�   LC)�`��*z��0�`� �C �OF��2�(�1` i�T��%F�d`  #	�05O��C*�2�d hA�4�L@4�H��Mh��	=MC����4l#5'������I$g�����y�_�N>���@$! hyC�5
~@B�>���,�h�@I��@��0���'���0B䃟^���4�(���?��;���z�7$�! 0�p�t��!�`�$��!!	�������g�#�o��~����� B��'�s����B��-&O�������7�XR�"����>_x�֚���wv���z�6�u͗��<��wqG����#-2�.@r���Y0=�喪�<b�\nZ��0���"���-��u�:r�ww�C�^�L������� Ccj��U	aT��/��/F��5��K35��K[��:YH��d �H�"l.�� ����3x�Fto:����{+|u"�ݵ�ٚŝ�u+�5@�uyb�ېF�s/[�j��f��񍲝*�Cʤd�_��N��-#L�-��ܗA/LE̾{��D��5��7d�F3�����m�Ӽ�\=���>Nwn��X�]��`@��z�tj�˙cyLܯf��6i�ٛF�X3*�w"��u��o�'v�rT�)����Sa���	���s歓m����5=��;t����	p�&8l�WZ��r���N�� 3vj�AoTҜ��Y�z�y�ս��">�i��i"p�ƭ���}mJC8/b��GE�3y�����R6���޹w�|E<�$�<wx�����4q%ִZ`�3�}����,�;��6V��E���;b�$F��F ��H�᫬D��q��>�B����X1&����,Y{6p��z	��U�4�nkCu����*�3E�8�b�3���Nt<���<6!�Vl �������>�>_p7qv�Z�L	�����Ԭ�J�b�D�A�ԝ80�]�a�u�^�7w�m��s˻7Y�l��o�,�q���j�J"̶jӛ�2C��2�.hHd�e���K{���k���Wh����wqj��4�H���LǾ�hْؒ�{���on�Y*�N^��
c0V���Єs}�����˂��t09��
�u���9�Nx,|�&o=�{Q��݉�����fTEd^�{y^�$�	� ��w��ټ%ҵ�,3��]G���`8��9�!�3�]�+:����i#&ۥ�m,��d)���Qc:�v��z�w1��wW�b8�9��`:�(1�ǋxg<Z/�`ӳ鬭�U���#���ӝ�N'�Uu�e a����aT詸0�]3��"��2�}.��,��q�� ]�ۼ�lwa*��ۢ�Ţ�����h�	R.#��؎��:֕M�����MUods��j��3k)T-��J/e��q=8�!��o.�d�s���3u��v����/!��s^��NA�ˬí�[���n��{4w���y�Z{�w!���;��J����e�u��KsG1ܐ�w{��ݽ�,:H�j��X:�*�ٺX�kN��,Z"�3lKp9�#����\��A����yq_h�ů!�5��
���d�	�Y���ƒ�vR:�r͇i{ǹ�KZ�#3DX���"C�;��U�gK5h����\�(hοmλ�i��i�p� DL#�z���AL�x^�2�fM�z�8s�����P]�T%[ >(���N�-|��nfF�MŰ�o�����u鶾׻D�s*=ٹ1E��当4G�`�e���׼&�_�0 ���tBݫ/S�,9�VA]�x���)������%�N�ΐ-DI��_-�	k��P�#��qwN	�B�&�����vsج<�{1�p3��<��+K����Ö ��ל%�ʎݐ+V:�n2m���'7^�Cm׸؊P(��w���ġ�]��.��_Y;��S�K����/��,d
���UUچsV���	M���7MU��te�5�)��xt��/v�� �M���w�ߐXȇbi�t��q�t�v�.ר�(4�N.��{@�~ߢ멩a�^�5�`'�r���G)�W<(�[�q�=���Jfe,4�X����wqH�;��[���ED�)�M8���6)o/��9Z�%�@`���]�z�r�	��Xh�IN4�����wqq
�*�ɭݵ��-'[���}xj�F0u=�5����%h�;�-Ӷsah'��лwxt?ndexw&�f���O8��0��d:����Q�!D���s�ˑj�Um��Ν�8��5�ڮ�kہ��9����n;OW�8/מh@s�F�79eq�.��t���I�xv�F�p�$Ij睠�\����5����
9��V�:#0�>6���(n�y��U�nt������5ۗ��-� ��N�NL�/��䃎��VZFp<��;�Yz�wrWC���.\TTӳ{j��@!j(B�B��;#79wq��޳�0�rݚ
�Ǻm�z��u��{lR<����3���΀�k-��<�#�C$q�q=�(��nL�gHN�rXƒ4��t�nj��X�d緤�d�4k���;��:|�<�_TS��i=ʅ{XG�+J���N碓z�뱾4� e��sz�咅��=^k^��
�G��� q�JKi��N�d�9v ��k	�������{���W	&�Aۇ%��rZ�����֞H�d����$�Y4�����v�D��	�I�]X�]�t�?J89�v-8�I�����n"7���9_(��i;z��v��l#�K�����T��jh�,+�53�lKL��f8wr�b�n���5�ݸn�}P�"-�Ǹ��Ԡ|v|N�Q���)��a3R����k���БѠ���g"�e������)*���h��;fܝklN;d�JM�g��ǩ���n��;.0�v�A����.m����nl�cN������%��q͓Fjmٯ�wV(yb�Mj��q��6S��qQ��tu�`��ŧFr(5�PW�βH�g{Jc��;a9��=�ҵ��<v��j)��>Nt�mĻy,�=��^��9��t�9�n��q)vǤ�齓s[���;/2�r�Fq��:LX8�{��7T�Ǩ���~���N����GXr��[ßN����{w�nuC���q����p� }z�����(�2���T���\yAٹՁ%����C�y>P��7��7waB�Ƚx𓥸Q艏	+��y+ZMBv�'u�f��7�?䛗��ʙ���	���uk�7��r���H4�"Ž�@g3��B���Bwy����lǫq̅�Oj�v�AΜ�������磩(��L�'�%��K�;�:Ocy�"顥R�\{�t�\�Fw!��@X�x?{ާ���d��}��b#,�2��wj�٠�r��^�{٫nWb�HE.����Ihڏwd�EةFex\]��2�13�v�[xt��枛�l)^w�6S��N��bݺw�؜Fc�^]��zM���h��C7V�NGh���}����8��0%���7l=��w�V�T����-�u���դ�MC�q]�;�
;'^�7N=��%a���q@�Q-: /�.�F�8�}�sE�z���]$j�z��*�����n�����n�`ǰ�W.����O�9rV)���}����ria��;��as���ś���&h�p](����t7���ɺnCY��3���K�f��`Ʊ��������:VT�.��]������\�wE�8wA>x���T���������`����m�\�PI�ߍ9�\Hfn�Bӝ��Z㩬���<H�&�6��c���n�=;�]e{wNA��^:/:,��ݲu}@-�=��uڡlR0�=��륪/;,p��"��n)��j�b���qse��qk�Sc[����3�̌�ݦY�M,l��Y��#gs.�'d4\���haM��).j�v�M	��5Q8�9�Û��5��K�K�t��=h�K�#�g���8ǳ؆�1�1{�>��L�x��b��j��>G���t[�q��v������#�\s��	7\�1��L���y:޷ALۛ*aeZ)����ͭ��Y���¹geR�z�+{�!��K�U9c�V��a��nd���ʮ F���-�T�&��G�G���"�\X��/���6�Bkn�d�n��{բ��=+�X�6���J����ux��͕�c�	b�Hވ����sz"ӻ�t5B���Q-CMN��˷�8�����z��C�Z��Ñ;c� L��zO1Q���B*�ϳ{�H�ņG
�XC-I:msGv�V��p3�ghk5A���_[I0c;
d`�#G}�`��{�Eۛ;yΛ��-Y^m�z���gχf�v��MVf�G]�sr�&�NoBi΃7��c��Ի)�itqS�L�N�&����}!���g�~_m
k��βS�23'އ�|}y�(�Nm��k���?����N�����IB~�H���) �H� V� �H�HVI(BE �`VBBE!R"� ��"� )J�B$$XAHE$�E�X@�%HB�"�$�I�	��) �! VBB�$X@I%I	R@d�,�*H$�@���R,�I!$�T�	RAd��,"�PVBBVHT!��
�*BY HB~_�����������8�s�G��$B��q��p BH><�BO�C�����D�Hq�Fvs�������k��kg�^�&�����P�+[[ט��w���_1�d��08���=U%��WJCƦ�Z��2p�F���B�<���'�{��ۓW��(ᯮ�D������o鬍.�ի���9�����s��`�r���}��tX~{�{7���8�_M�����'?��Cc���g���Cy���k����Ķg�Ef�	��[��7�,����-�ݽ���=��᫯>�ף�b�y}ǒ\;I�w��5{��H��ە��q�$%�ݹ枯l1�|�ux�i:g�]�|������{l����&C����1����_g�g��pۆӻ���
�ˮ�u���<�4���������	n�=�Ð��ě�25�]���5G��_�Qߏ�j��7���{���ԏk���ܚ�;���!�k�_%%y�nS��F��v?{s�.��U�QW�y��_yX�=�ƹ7g<��ww%����9�n���V�$b��O>�����5��f��D���g}��JY��^�B���������p��d��^�˒`�~�������m�d{Ӯ�w�����^9샯��S�,���Y���}�w�q���_�:n����[��*˻�~���Yؼ �S��6���aѸ����"��V�ž8[�덇Ǖ�
vE�)�ǁ�����x�s��"���{�;<Ut��7Ʀ��&q�6;��ʩ\T���;3˛Փ��sٯ�Ʀl]�$�$Z1>�nY�|p
�P��0=�Ů��m=��W�-�5ޮ��@�A�9�ڽ3e<,}�d��8��3��J_l��C��ť���;��>�{N���� vr�.A��g�D�.HN{�c�OY^�M���K����M�g�es��E��^�JW9�����3��zz�7K�Λ<7I��
!��wW�m�����dv�w�����Н�3Fx������n+���Яq�t�}���Bk�"�H�ǽ�<�Cn��}�nۯ@�t��*��ި2vPS��V���.�h�#�'�J۾���ѡQ�����b\�.ݏ6
b�������`9���j�YN}����΁���3��q�V� �G�6ǫY;�T�;������ܚ늎���F�?z��k4��,��{c~ٳ_I��8���.���=E����E���yE��N.�j��7�����YQ����`�w��#s����{��|���w/���\���Fק}��z��+n�Æ)R��W�?&�Kp�u�����MH�к���G�lw����M�w��l�Vx��ׄ�v��4]�mhP�7gJq��\#�h�%��)u;��K��i�u��r���}�#9����}ˎo\m�"
|NC��M���p���r�4�g*�_AY}p��{�նM��vm��ݾ�#��xz�� d�E{�5�y��Y��=��U�F�����I���O[��KȺh0r��;��yL�Mt��^��{7�wA[C����
<4̞��_~w�Q�w�Eg�{h�/k�w�<�g.و/x�}2ou7Fm�+|���;ڷj<���=+�A���»Ԍ����m�N*{d�]���@�vփ�1�kxQ*��YBY�r"
Z,#�xrc�cۃ�*��Ͷ�F9�m����yg�׫ç�zxxW����GN]�#�	>Y�z�g��6��3�ov����:���M�Վ�<{@�-��Ѿ|�}��1��O���}�,���x�8&�-���z�5���{�����D����1ҵ	�v��3'�pv!=�z�>�Ps�'�{D�!I��{�0��=6?x�����/��n�{��s�6@��}�o������y{l���po�Y�j啀^�oޚ=���Vk����=�ir�ɼ�}��N^=:h��o�� �hm��c��qgy���2�u�U�og8�h=���G�R<'�+�q�*����e��|5ĺ;�\]���n��z���x�qg}=�a�7^���ǩ}z���ɞ�a�Nc^�t=����Hl���'���l/hQ9=���<(�tb��V��D_�ic}�$�>ꔱ�Oq���� y�dh�g��fe;�W���H~�R#�}wWrÜ�7�W�;o)xӏKp���$%%�7&�W^-�P	����E�cn�l��OԱ�o/
��~���I�L|�:�z�G���sx��g�l���x{`}+:,I?D3U̉����� �-B�����������ᯔ>�APE��#�D�E��4Gt���0y[�)N��/�w���==��h�*�A����O)��ۍl����s�ѴS^7w�kQ�O?N�����t�|l�{�;h�1��9�����<\����?�{��k{�NA�٨>g�Toپ�^�u<�������M�}g���P�}� =��n��ہH�"9�-\��|��׼V�f:�E&Li��=!W��\YEgG�nwq�"�Z���}��ϗ�Ӑ;|;��{�-���׏E�[�=���{t����,�Y��<9(F����B2:��!N�+}���Rh|ԙ�]̳�5�K=��&����MsOk�������.J�wxp�~Ӟ�W�Y�-Y'�ݰ��G�����������8������g{C��囇1���4�I�" ��_����l~qx�o{�%�ͬ ��_k��>�l�΋}h'�|�|f���=ýVp���0`��pK��A=mӤnz1�7�E۞Y���8G���N���*�� ��6�A���.���U�@���`�T_x��H������XV�z�g��ޞߚ�Üg��0�Lپ [��+��p�0�/+��{9z�����{O��aS;N��l���C�x�Ȯ
6OqYF.�i۾Ü�[�=������W�����oI�;_��}��.�{�ѿd@�.g������[��}O����4B�����zܩ�.ݾp�k��ܙ�6o�ma½=/���'{�d��Q��h�	�b�H���|�͞^*f�{.p�[3̉�B 7����-u�q��-�n��/�#�������^�14�ͥ��7��,1ݾ�0��k�XuC�W^�dg�k[o���{�lᗫR���{��w�{�j���V=�@��ږ�Ҧ�p�^x4�ݕ����n�U�! �xO� ��m�)w�\�[�G8����}6��q�9��=ݾ��ͰwO��xݙ}���J;�U�1��g}�i�{�N9b�y-��r�{�ML�����]�Ix��U�1k��񻌍�n��n!����5�)�.�����ω���Az��[���E�^��/`�J�,��M�e�1�7���o�t�m���y��`=��;����{�U�TN�1����{���ڍ�:LHAnv�#R���]��˺�}WvG��v�ŏX�vz�tXqr���Nh�k8�T*}Z�'�KĄ��,���;ٶ.=nr���!z-�س�¼2�[��1���(Ʀɼ<��L=�Җ8�)�+1�n�_�t���^K|QN4������w��Ԗ���p4�,�p^8�;,�z�}p���<����:����=9��yk<�����y�>�d�F�|| f��K�����ٯ7x{��Y�H���L�Z]�{�X�q��O5�yo���c��s���i����A*Uu��kգp/v��z�\�p����e�Owqe$L~_q��e[�W����<~[�WU���u���u���Ϣ��&� ����z�q[�~�姸rp��{�M��9ķ�e���Wɍ��m�ƈ�ҹ�\��[F���O%�!�w�ǗK�Wo�ն��q{�J>v۩��ECb�����M������B��)/�d�(y��鉇����k��nH��oo`N�a��!�d�N�IȂd�v��Ŕ��y{n�Sn_)ot�d�oB��ym������w��be�vq���H�4i�����w�no���h��^��}��$9b`{���y蕡nr�#k!/t<Ĥ!�G�WNҫܬ�>�t����{���u[�y�܁k㋷q:b���7����	��`��}=�ƣ�u}����œ]+n�(��pF�{([��^����d��������I���&�oi�r��o����YH͋O	��+J�ah�+�c������+%w�ԝﲱ�9I�:�F,��~�t=��M���-��D��!`��֓�z��O��A�>h�콧|vM�9����˷�vox��t��/w>�'����'a��.꺭��~��o�vQʘy��M�4_�Vf����1����>~��nz�l���8nx�q�:wN�wc��3�Ậ�����y�Y(A2IB*�����QRnuJU=����{��@A��d�9]C����XR�^,T�h�|'˳�BB��'͚�WC���2�v�H�$5[e HF;9�s�����L15č��i�"l#V���B�Z'���+�`D�s�����0�b4�thФ%fc�3*U�V$���Q	I�Ѵ�(Z����'�3-�Z�Us�ۆ�����0��0���aβ�V�\�j@�a�����l ����f8�U0e�N��4f����Bg��sui����I�Sn���HT�96��R�6Y(-�)@Z��V��4�X�-(lK�E�mTjf0�n��Rո�Q4�3]�K��[�]d`Lˁ,ݱx#�gJ�oU�]I�j(W���F��.6@�t3�4������*�Xi��7i�*�a�u]�V.��6)��5�kU��gh��
#SSLZ��Ȓ�u��dt9��֤m6	&�28�6�]�� �m)K����бц R��e�R��Τ�� �s�݀�W�Zeā�]�,u"	�e��t�[���l,�Y���b[r�X�\Bثm]����u3hYIm��BkR�E�17
��L�K	H�-�h��-�e5�� ��	�[�� �\\����F J�;�[�kJd�yܳ]����,�B����)hs.Ń�X��hsL�]Gj[vb	�F!26+��X�騥M �Mm����b�qS(���˝�ذ"ʂ6F۶��˱uz���«���kSL�ܜ���v�,;Cb[k����R\d5���-)sP6
]����m�棠�IB��ض�5����"1�[̦�h�Mn�K�a0l	�Xd4�zc3H�жb�x��F*�c%��f�%ṋJC,1+6������0���0����d�5�3 �]Yg	2Bl.��8Kv�YpS.�ԹD�515a�0�]�2]����#l#L�%����cw#���nL]в�D��Xɯ�7e3�$�X��e�m��[�Ke4B�k��j��,f���[דRы�e Bb��5�����q�P1�6��%ul4l)�
p��0�nQ%#6�-�ٴ�m�F����׆L�jVk�P�C&K:�ڻ5֊�66iE*K`Fm�S�Kr�뛱��vh	���b�McB�mц,kTh�\M%^55sk�^f�C6��d���a�䪳3G�#���4/kz�-�n�c�f� ��l$���ֺ�ĭuB�&�:&���:����:�j�F�lj�6��ni�[���c��*�[tm��q5����歮;[41���ݶE�4$�XX6-BQ�R��YU�m.R��%$#Lܰ�Mkk)nG[�.��Ȳ�� ���]�-�mj�`�4��b��]�I�y��J�[�K�c�� ,:�����%f��ٙ�Z��殶�Uݫ�,�C5êV%-�ݒ�Ri���v`U�\�ً΍� �Z�sa��Qy�hذN��an
�͊X.�q�n s3�����/�@�I�1S8�Y]r,@	�p�v�4�c�Rm����-4Q\�IiF��!�D����!2�'[XE��D�$z��-3�3�hժX�`I��TF;�����`�[������#Į�\�8u�Ѷ��.*^���.��W�h:�G�lٶ�K�2��Ch�lKf\ d�1���b�ͳ]mj(�BmHԂYZGB%���z�]�9�jʍ��A!�V�F�i�P�Md�seLBhKy�(�<�%�7�Ÿ"c5�q����aj.����+�f`�iR�/+�K���A
������cD�ݠ`%��4�z�2���؅���X�Jh��+	� ��f�=uר�iI�+� 6�b�H-[�'U�4	���t*CM�5�J�y��`0c�f��vx���5�ڐ�Iua-��-�mK�*˘��M���M(�WQj��X�TYL�X�J��K�đ������� q�8,M�X�*"�\��[�]al�+i����]�;�V�QRꦆ��c����1B9Fk�p�T�b��t���L�3����&�l�e�5&ujh4��=P�t`[��,҄��+�h�tִl�ݩ)�-4lf& �ЧupV��Il�/d�C�(�l�b�c��ǦR�͍�(��a�ږ!�4�f�����[��m�n�4�1����E�i�2�5a��Qɬ�cy[��b��K�����3S��b�Ҵ�/%Ҙ9��M�5�ԁ�bh��.,��B,i��R%�!��!��iH��T���:꺚U	������̱;Dجu]��j&�m.����iU���^е����nL/b1k�6�-�ԃ��,]^���H�b�h�0��Rb���8W2�M�Z0-�p�M������,�6�� �KSgv�(���e�����^���YLn��9����Me�b������j��XX���M��6�֤���@�`Q&m�K�M��qA��J�]�6�a��қ���!�1H���Z֓m��a!�J�`�K�q�)e� �m�JU�@�U6��knqy�	l�m��m�8h��s��df�K�;@��A��c���8Φ��̓6]�,/5.Й#�]��K20P3*\d��Q�M�#��1`�1��ň���Q�:]�5�F�A�v	�g3%
;#��V�7M5��]�G+��8ٌ���P�^6.q�c���T5�\�hR���������ă6�RfTK���v�ζ�k�׆Q���R7�����R�굂�Z=��.a�뮫a���,#�Mm����-���.�,�L�琕�)��u-���-Ch9є(�k(tZ�Z���P7�M��P2����ͻj��JR���4���\��`1\�Э�i@)������g!�4��30��ȵ��a�L�r�t\�1Y������T�������M�6��mţ`ȸ����cK�i�F��2�e�����������l����c�6��eV78�U\��k���Ъ���Z�I��)w��`�+�V�]u��-��`��\9trR�VL]*ݥՕy-i3��%��
�ma�G8RTXh�iv&�Ԛ"�A�q���\k4ZL��h�V�kc����ײ����nX�F�kv�\k�3�m�� ����
Krڭ6�b���������(-q��(��`�iR��j�h�0�P��T�%id�J%�aEAJ5+��QE4"�P�Vq�bJTQaXT���:С�V�qF�+`��E1�:h�r�*VJ�+FV�)*
E%clƠ�XVMی�VUeT�I\�ga�Y&�12�ҥ�(v�m��K�wZ^oF���ݱo[���9�Œ�x� �[�KAV�*+��J&�m�,��i[ѢE$�.;�Ԧ����!%f�$� Rv�*6����X.��f0QeAV��fc	�SV�2�Zu�I/��:}m��{7�>-r����R�e�����5�]k4f%���l������ڄ��R��M2�X� ��#֕V��a�R��i��t��	]tX.2��(ő\l�K�W-)�g*dK+�\�c�fkP��H�a�i����aZ�Iu`��b��4�hL�4�5�0�M
���u�ɵL�f�cE1X�r�Ð��#s��;+-�����$��,y�
Z��2ɱ�&ڀ��tK�����6M�����R�[j8�ڗ,ۀ�CMmp��&�T.Vi\)4֜$Cf���5X��*3���X/j��-1�3�J��[��:�)�������Ԍ"2��4.r���ͨ�5�Ջ
l��9���j�J4D���v��v�]�R�a�Q��,Ge���S��TҎi�km1kzTf�F������p�ҽtk�
˃S4�(ћ���	J蒰s˫<�O
xhV�ss�C�4�Bh�u&��JM�&Zɉ�)o,[2Xaؗr�e����f�3[
ZG!��Gc���&p1ʹ&H�K��qF��&�������ڳuWq�L�:16�]����̹�VhD*��f����l��W�AJ�mu�Vf��7��m��A��B���%Ե�֮��wK���#
�-`��
[�cciX���ؤJ�Kxl%�*#P���p`-���6��y��e@kִxH<�9���R����mKU����y6�X���
VB�
�_�������5�d�A�НH�O��}#��5Dn��D��O�,�={Z����M�Q=�ze��	r ��O��my�Һ,k�h1�ʾH�	A��� ���00�5�����
��A0��sy���R%I�vU6��}[�0ɓ��n��ʹ�q��APȝ�b���F��TI��M!�����li�~$����ȳ��1 ��ϐ����e ddbf��l�&W#5v����<���e��{x*�=j��6&^��T!_����EGB)%0�6��eg}��y�Y�Gp��z��/�I���Q]�s;#��]Y�«c�T��Rӄh$�ה(�r�:`��θ���T�R�»���{5� |A�=5ѕO`�6��s�^u�IR��CL�7����Ea�l�����G���U@V5��RaU�U4���^�D�Z�U�A#�R �Ҏ�>�5��Q$@S`�"��jsA�F �n�Go��^��H���ج��a�u��[�5�Q��ۡ@�ޔK܌���&�ř#�O3�]�����=�$���N�Q����$��^��pҐ )g|�ޣ;���y��o��"-^���n��B��3
���\�}��%�ϊ�ߧy Ap̓���d)Ja]�Osg�ݽ
�ͥ�E_��o{#o�����_U��3(תI����ݷ�H$E�屆I��B�5�w2�D��E�gk*M�G$��ky�2�K�lmv}���c�u��M�����b�u@��1�3E�t�24�$eKrD �4iӡ@��*7�h��A$���ha���iC����&��v�Q�⒗W���Ϥ��Q����RJa@mj�����,� �K��N���}�w
(ǽ������Z�k<[x��f�x���Mz���w���<pL��Y""L�F<�SL�*�w��9�!nb|�6	� ��
-�@�,d����5p�Y�˛vɲ�C�Ff[F��2۟�߾�E�6O/� �w��ܣ3Y}l���(�U�H�M�s�j$�n�\��� 7�v m":"W��5��ܐ���Mб���15¼r���0B7;���԰[��Xg���rފ����~TA�k�Y릠�i�V4諛��RJa@�S�,���Wv����>�*�#A3 ֜�ຳ���Q3wy�a��7���k����/l��o����%�<�A�|�?.��,�+t�ιk�2�e�h�ƅ��Vf �,Z�4X���@u4B3��f�1�m�1t114q��/	u��]�B��hQqaV��.T��kvՕ��ՠ�˒�[ML�Cg�TҰ���[���B*�Գ0�h���{ZY���1v�cgϿ|��;8νTI�����adV\n�N��t��(��"�&%B,��ċɚM� �m H%�>�3ںӕb�iS$�%�Dt���2�_Q[�:N�:�sR �f|z���!II	�G��W��\�$�D����p��=�kr3(�^�}�f�֮\�� �|�n�覆/�n�N����T������+r�5��.\�}���eJS
�Il�F�t9ӎ�ո� �F�m)��T�X[�TC���m�Ϊ�����#a�c/\�WW�M>�޺QY�;w}NE�S��1E�:o;� .8ω��hQ�v�(�z��%*GQݽ(|Ϳ�=%ז�{�-�_>/[T9��$�U��	�����p�p�$�z�	�{.����bjHRRDB��(��}3�[��7E�$N]�z���.�m���Aў ��m�&�@�B��
v6���N�I��pE��|(�s����ځ������!�[�����H��լ{�ȼU�Pi���v ����(��͉*eIUe��@�sZD��y�r���D�8�ֻ���J	|y�m��Fo���U3;Ӻ }�&��T	>���}\�%*LJ�Y&�\e�a";P$�{��^�v��o����7Z3$�
�]>g��TDM�Ea��Da�$s�r�N��p���9��{Gf�,@�.��ЉҪTʧRf{Um
Q$��`�2�$��d�V'eP�w�	{Ҽ{23(�_>��Q�=&����i��R�Um�VŎJaJ��>S�"�2I&�-	���/��<�HHp̜�ٱ%JS
��z[�EE�;���fI#�o%�r��!d�Y��ZH�X���'��Ξ����ig���i��p�X�w3�[U��#�&���k  �<�t�B*3£H�M[t(X�;�����p��ͻ�(��o�s���n1�����jG1�e��0���9_=��hf?=3�>�L@'��-.iE���йH"C�d�CrB�$,�ͻ��V�<.��S�P 73j�;C}W-�i/63	3M񣀒K����$=�����ID�����k�S��v�yΠ���@�o�k��Y(����d��bJ���mNk�*�"a���o*�|�K��~>�5~�'���_��T^6X#v{;d�y ��9Fs3w�2��������y�?���f�(�si��fmi��t�`�*`���fz��`K1.�1�tf&҅ن�go5�G0q��Y�����<\ʥ�l2�nvk(�,s�8b����mx`͚G5X��.+�Sh5Fʹ˂�E�tpZ��]\�k�8����P�v�f[�t��H-Pܕh�o�_$�4\}x|V�o��TI�i�R �T�2�cUܷ�EE9¦�#��pMd����v�-��%^��{��N	�!II2�f�H:���{��p ��Ea�� �u�@J ��`�/S����8��*�I=�y�R��e�4�[UUq\R���6�A�Jw#����۱s2� Z����I��A9�Z�����$�L�v�NT��g �D��O^�T�0�j�u�֑�C�B�zܪ"��m�ӥ
�Q�ω>�g�:��64��I�a�Y�!��a�}��V���F
vz��v��|�2A;����̃��Knf����n"��u�PO�+o������7D���^@t2$uK�%$D:rr�MU��/j k�B�n��[P��yӽB�R��,����ߨ�K׭ř$�t*Q�����t�Ԇ�2Ͱ:�n���Z��ƻf�������Hܨ��ݹ�}H�sTC�"e���$gn͈*R�Vx�˫�J�y�C�zP;��h9X���kos�>�ΖGUQ���vZ-�O���������h!]�V�����$�{Ǥ����ۯg�{�nw�y�/gkx�����1D��d�b{`(��ބ^�~x\���a�ˌe�:OzVq�7�gL�[��v�󶱡ﻆH��Ӷy�=�̜WN�yg�Y�ag�N��s���q�z���'x�������,�#a��+t��t�*p�q�ɬ���v��&�<7��FW�]~��l)���KJj6w��ڤ ��]�y���d�7��Yڸ_(fS�KNb�-�q�=�H��O#�e�f!+��Ho1��{�
 �!}�T_�h��w4�{�z���C�x��Md/�}��y���=$�����'�z��}�2y`"w-�%��	���~�sa�D8�׮���/y՝�������s��|�m��G���Ҿ���F���/L7�����/\�L��w=�/3`�n�E���<����-J,��������2<�k�-���r�����U���1d�����4��1E������2�U��*fV��[Q�<�F�P��k����QHLK��$f�B�Ŕci%��-�J7��y��4.8�9�%�T$l��IlB��q���b��Lr��UV�-����XK	e�Ѹ�^ ������w��BìD�B�[H5��J���[U����\Ū�b�m\n�Uch�%�-(ʴ�"�X:�����^���[qH%�$B���fe���1(��EAG
�bU��S&ư�lU,���%мKh� !b�MYoZR� `B�%��ZYi*��A�4��-��z�A�kJK, V�!�m�RX�KeV�6P��\K!ԭ�(�-�S����FՇ џ�$���$���
>�∘2��2��9}�=g
$�V[U�}�ŭ��t��"�"c� �|3��yI2��D?�f`oѠ�I�n�@���*]�y��6�a����H.� �F[9�Au����}�������}����<�pV8� �K{�F�očʌ��ۊ	U*���2��ٽ�V�H��#>	���sbJ����ͣ�|s\�H9��y�޸��d/UΫ�[A>\h�)	��x;++���H8ꗫ�ڂ$8f:�^�U;����s*�i�l��9g���mJ�d�/��Ձ\��m]�'g�	�ݑ���][U��ڈ2%b%�D���"f�B�s&x?
�ʡ�Ƞ4nW1EΚ�IP�����c�%���B6���P��>����Q9 �fo���OC2�v�0ܞ��Om
'�R�a�LJ�7ař!d�E�.y@����zP�%Q�vu_+�$nTdkvw�I6Y��O(��@���͛�RP��w�c�څ�������^�J��Q�n�gL����Q^�dI|�q�~���d2$���}�ٻ��5�}������oW�'���(�Vx���lU�JlP�L�e�
7㽧�}Xb���}�7&q�#��I���!*�i.��k��8���1� �pTn3t�gA�%�\�íl��W�u��<ᎏ:Wfk]tmv�I]��9�����i�#k3R�
�k�%��`�n�Zt�����(Z⪋s�.P��T m�II�;]DMe������T]�����
�M��� O2	$�|�T��T��i.0���@rB�EM�V!�:��Y.�v�}8t�>��
\c��i����&kM$�[�U�"����}�g�_6�_k�$nTdv���,O[��
�P5oj�-�oc�
v��⌃W�6%BIJ���i'5�����h��2I�P��=�>����=l���ov�e�1���3f��9ź��n�s�ϞDH��m�@+�rZwk���;���(�	;��(��ځ%	�2���.�U�rT��1x��V-튙�'�#�}��%+��-�p�d�5"yN�PCI�~�8|��uQ'ﾔǷ���O��3+C���B�*{-X����?L�+�������;�;�*r��ۋ"��p;^wywU1��8fvx����JҔB�@mH�e� ��sĀMcH�2"F^U����/�>CjX��Ѭ��v�m��k)r�݋�|����������!&�$�㈦�NI�p��ޥ�317VH�B��f|H0�]��wu=���9ڀ��;�:o/K����7��iҨ��*l� �� ��g=ȆV_<;���������Z�����3���`�+biF0�?{�����N�^_��@�n��$c�Ee��;��ml�tT���*����:s�ETe_Vő �m,���-������O�F�� ��V����M��R*�)�`��ImE�f�H�[�\�>}����ۨ��
 �Ȧ�,���v�����d��6%BIJ���Nd��z���]��oJ@sdAg=��#Y2.]`�D���� ^v}��}3����� �'ĝޝ綠D�BhD�e$Q�|C֑>'����}��՟��7"2r��I�o�,Y���4�|�ξ����� �މ/���}����#��Ơ�%"#��}�J��֤zEwO��p��ZJ�Ŵ�B ���ɜ	@�KLR�N˵j8��T�����UY�� 7�Q��R&��4ӧ���!q���S��d�ڙ�S�YG��To��"Ѥ�k.��5;�*JU����Ƒ ����g�]���Nڰ��HC��������ը��� ���@4°�,f����6��(Mu�y� �F��ݠ�H�ԁ �ɝ��٨t8>W�}O���w`�k�ݺ�-��LeV��gn�H��d}��]�3&:`�L�hW[Qm޳bq��s��9�ιR�"q��a�������܆m�I��ּњ�i K	�(�Mr������X�j�F)��c�[��d6�1XF�١Vc���-MsR����l5k�Z�M���� e�K5�.P��$J������ۑ��?B�E 3� ��JF�q�Y��۸���Ay�8�*�+�����ռ���� �ω03�mL)�=W�#�2;G���4� 9VT��ۢ����2	w&�(I)W`�:�)�� ��H�N�}'��lR�ُu\�Gr�R"D�v��H̠coK漃�d�H/��S�⹅w$��*�v�h�9+CE�&��sDYGU6�����v�e���N}>� s䎑�[:�E�/Q�/.i���ĤhM"�$@b/wٓL�n>�˨n
�g8ڰ�}�J���N�n��T}��k[=��렖������>�V/�8�$�_ߤ gt����l�]���pR�ͳG	��@>�+V��x:Q��H(�~!N8��2�%v�8RB>2�S��9�m� ��2q��2�9�
JUX=֑"��ٗ��A!F ��H����s�}�<�?�:�<�"ݶٖ�gHJF*&�G{|}|����5��R�M^�@��H�+\�(�$6�y�m�TE\On�z�����ҋ� >�l��{vA^��V�z)�sA��R���:�A{"���T��6zcNq��^{7bm{7m��)��t}��D?�[y&gZ�eǀ �>�o>�/�� �Νh�J*��H_n�Kw��g��A��+ި�[\���rI_S�2;3. A��\����O��(�YM��?>Y�ֹ)\��:v�[5���W4�p�W���w��W?=8�P"�$��Lύ��7"�O�����H�q�E�qmJ�K��v@,�I��@��V�p#���@��lB}�#O�ǩw���m_��.sd@i�#�y�c�*g����yK�>��Y�M�5F{��N��UfوB�u�5͋K�z��ތUS�WZA�8}*0������x����@��@!J�5�Ϥ���#e��*��%�H%ř$�/&�=yӘ�_�h4!x��"A��E�Un��+����9EA���=��B�q���_��W��eDr�N���8��� 0{A�w��$��ݿ@P��WW׷ xP ;�_s�b*VP��Ҳr��H�B�Y��[Hu���T�}�>�dSپ�iԍ�Y�r�,�'��Q�H$�Z�ۼ��_�;N�(���@���D���-5/ol�9ًx'�M�̙� �����º�ne�7G�St]�gM����	�dՉ5�{�N{Q$�=����ݞh�{��A�u^�xǆ)��fɈ��=���p���4��_9���vټ>t:��5�_��6��L� ;{^����!���;����N���Iv�o�����n̰^ۊm��ʊB�{K{�<K��"+ըR�����{��bͽV���o��f�t�y�o-����I"/�s�Tk���������%�����FZ̓w�M�Fuղ� yy��[��"2�7��~3G�TF`׾L�z�wۖ�S4�(�V�6"���YǑU��$�N�hWx��ͱ���l��ɻ��x��`�<Ł]�t��|�ݳ;�yii��ã���Z�S�N��qh9����y)��Ԇ��(��,��==9K��l&wiڧ`B���O�"���yM+r����[ў���
x�:{����*r�3rh�wƷ���ݨ�M���׀�_/w��<=�F�����w������(�e欶���Q!�1%���4j���%�,!m�~����z��V'	ļ��^���$eZbe[�)��q.QXŊR^��e:���j�Է��V���,�V�+*�Rq|JjYD���ڒލ,�l�P`=@���0(7��s�֗��+r�
����e����eX�����\�d�[5�i@��4j�����^������Y`��6D�N���1(1
�C[��E�����Zq�[
"�[�m.Z���A13�)Z���Ye�FPH����ձʠ�+rҥ���{��8�t��Z�jv�r�D�e�"��u��]1H˶\소4�)��.ҋv��f�6�	�65��qF�&�睑�.����'2��D��]�͂�J�E](CRM����SY�xWmQ.�g:�f7X�������T�0ՕD��X�-m�.M1���j;-6�N5�;hKj8�Yn��+D��\Kf��0�,�Z.�*A�
[��h��ai
�6������i��Yj :l�iNґ���24Qi6a��4���Vi�ZEy�CC 
�l��8��D�����Q ��l� Զ��rᕱ�.������mG���j%�j]� 4%�h��b�J��1�cA��0�U�\��Fd�Z�U+
J�\�s�o1�t�c@��&��դ@�K��A���CCM]�F�D��M�8,m��6Y�]M�oh	����`A� ]+X����-5EXkz�MS��L]`a�n��i]��V�5�P�M���Tخ!-)6��F� �5�/R7p�C#��b��9�)a�WbS	6a���[L��E͘�`&�R8(��9�����a��;�ѥ�J��]eW�p�b��B�H��UYs�f���b�&rk�5Z���U�]�p�Z �̬Lb)e�ĥ�6�,Sb��X�)m����m�:t�qZ_�L.4V�-P[�<�)�+l�7l��k�Ά�Jڃ�;u�(\��ʾM|-]�0Gf��K�d���js��SWAr�N�%��u����[Yq�˥5�Zb�L�lV�CM�Tf���«��M������%�oV�(�ˣ��p2�%4:ET�'��_���*2�?S������J?n���M��>"A �rG�Z�&aB��sR3&�����A�ā'� Js����@@���+RH���Lr� �cH�f�m/�#چ��7��ע)Y3� ^e@<ay��uF�:K�^(
R35fi��t�-���^gj/_*�_� ��
.M<�x�^��4�+�vc�6P�94���4n_��=�
��%�� }Ԉ#O57�e�y!��$np� R�+�X�n7�M�Mv��R�/�)�_��3|��������	��h�Ur"a���������� ���$���$u�w=� ���P����Y�g���e�k2P$��2vl�J%J�V]1[��r��漈q�7�6��nF\�:�HD*���K���n܏7�����^�S�����Y>��=ĵsi�EK���������5�EK������X�^����ә=	_�`Ehғ>g��[Z��W��a�&\c.f{���3��;r4��<\i��ˍ�2��)�'�B��Rlzv83l<��<�u1a����]"������鿿 ��~M+C&&(*��Xh�N�lyӑ����s���>yhL���C���}9����[���7j��nn� ���5i�)$IX
ۜ��ɣu��ܰn}����!�'"�'��M����++:��m9�-B2�Re��_3�F�݌���qo���킥A�J��H����9�uX�6�H{��z.�!J�4ݩ�{q��x�}��#P�UCE�D�[�pm�r�v��¯�ށ4��q}��������)#��������r��}*�p]�X��o\�﴾�e{�'s�:�U6ȢTR���u7kRq�hￏ���J%II������`Bq�*[��|�E��HD*���V�B6�o'[��uk�����$�I�c�ϯ��D�1�e��gt�+��)Q)W��7Z��r�s�����x��z�@)�ԥ������u��s�]	r2�����'��?���|j��|�Y�<�x�?!��c��%?L�����6��`��3e~��?�U�e�����Ӥ��p��Kt5���؄V���*cL��(�%6�I�hAV!Q1(�Հ�Yb�V�L��bU��X	`���-(֛`Ե5K�ZH�az�xvٹ�13e ��	��d�U6��b�vD�`9A� ��k��ؠ�h�Z�A�����]���L ��]�{���ȸ��z|�����}�D�Y���H���	BRR�.}�;6^�rwHqoUa����y# R	K�+�G����e˶� ��zݤ��T�'U��$9�n�o�j��s���W�!J��J���7�q�6:|+�{�ϳ�<a}���Lb�b�f��m
�V���ѭ�l�<�y�	T7��\���Gk�{�{�.�<ۑj�3*]�]]��Y�bӌ�
�ɲ;�]*���9s{��S�{��+w���Yg: pү��م�~�o��϶@�N�����9C�tu�))8��s�u��[쮐;zw$Y�
B!P]��@�R=]�7zUj��Ἀr5�rH$��=`7�퉋�ţ;�(�ӟ�1�`�~�7���4�+K͗M��D��	]v�͌m��>��g2�S�d{u���"�U����ފ�	-�yq~�.b��.}��쪜�Z2�wR���+V�����N^�k�
N��&f��=�����O>��Bw�N���tnz�b�ڪ�B�BSQ�g��%�����nW�����dm�))8r�:���S <��o�tf��2rET�<��b-�
��[��Nߟl���o�M#�j�&�0�7l�[TP�Ȳk�ٙ�Yb�6���Ͼ��{%}�	��{dE3��F��B	�%o7��R�)䂋�*�Hn=d�kۮ}�NP����� I���;.w�<r�&��E̎��{$B32���5Ud��U�-
�� s$���:�y7|�K��
!�M⁵�`(ȗQ��ˁfȯ�s.D]j�ʜ�:>�OĀs:q���I����,��O
�������H �5-<���Z��?J�2;<B*��Z�@��X�n�&%_�2�2�B���H�/vB���	;Q�[���in�H)AI����LE��I�ԁ�t ��eˋ���[��R�ʓ����<� {\��o< ��� 7]|o<�h T�w�(�5~r�"I'\I ��ՙ��Ij� ��t	�c�V�N�Z�c�^E�H ��ɝ��=YtFp�fFĴ�7�y�\O��ۙ���Z�;����<�V,�#�C<�l,q��ٹ�[�����=ޚ�P�cuH�2�k�� Y����bje�a��#0��%��[�l�������h��(]�[6e�n:j��9]�M����E	r��b�����gvE.���j݃Z����Gb�jl�`l#��]�ة��V.%t�t���e���i��Z�����3U����'�p��TC��l�˨�ƫ݋�q:�ja~42����t�@ ��0_y/���q^���y;=�+{y$�␲�Ѐy��[|;&Y��H>��{bT�R��]��h��P0��ϐ}�(�Ř=���ȒC�.�%!�s�<kʱ<L8�HBG{�P7v.�V���m���S�Kh��حՖG:Ħ�Lg;]�u������4c秭�I�h"I�#���]���A ��N��BT$�Q��� ٣Z\�ta�ʧu�wH�3�zy�v.����p�p+z�
�M����+����ŰgF������d{�Mo$A��D��U�,��'�f�7T�O%��$>���jM�|Gvϖ�!���A$'v��}�����˒ �eD �c]�i��*�� _\(��� _�Y��?\�;���"�Ax��D�OtH<��1����m��-h�ι�!�A�n�q�Y�u���������aT�~��wg`D���-ʽ2q9�!^]�U�����Gu�������t�os��UM��=}
��I�9�D�E�	�~|64N�X�����#.�nmZl5�Ǥ����/���ŶJ����3&�P���{�7���؎{�����}�����Efn�W;4��*��\F��^��v;�Z�9�|�����Fi��W�r���<ۺ����:s՝=G���������J�����71�v���0;�NO��9>�k�D�^�X�5/�{��?�+gy=C�h�&Uø�_g$�}^�6h}��h~Q�ݝ�^F� �4{�RB��#�����9�O<������ޚE�5�����G���;���,?z8mi���ͭ���Ǟ����2=���T�}�\�FX�g��{}�sބ�8���b�4�y;���
x���r��KL{i,\I?t�m�+�Q:4�����;���;ҷ.�V��'9�2���@��aF��({���r�<���Q��!D�;��^�;{���<��1�ٻ��e�y�x����@v��d�d�۽5�H}k��Ԗ�ͯ~�S�x�FЩ�TX���ڃ�+Z���[��-��ZV�ef]�����f)ƪ��TmUV�[e����1̳����(��ɋ-Qb��	P�*�QH�b#q�]o0b�e�F0CV���TXʕ�F��A�Tݕ��V�V,Q"�QH��"��iEQTUH� QA4�*�QTCUJ1�EAX� ���TDQ�`�#U��E&5P`����cQJ�ukV
0b�r�Q��*bQ2"?(I��
-��$D���g�(�+���]�8��I�$��P�7�|O��6�FPAIcO���{&5ļA
u#���݊?.��9�H΍uE%E]ɚ�c���LKXtdu%�}���T�U�� ��@}��_.�{sDvD�n�$JTyJ/]���@,�H �Ȣ���]M
�E��( �l�OW���l��y�:��s�S΅A(I��i�ǙS0
S�|}�Ƞw2[��J��G��
�%��*/2w/#;~2I�A27cy�����?$n>�{��,��� ,�z�d��A��s:����-y�$e:��9_L̐��w+��Έ>���Q�[��[lѸT�%�ꢨu3���R�/Β>���5�C�ޑ���I%VL��"��-V��@�6��)>#Bw6D �K�L3Z��ᘢ}y�h@�H�#�v9D*��أB�G����9
���	�c� ��.)�TL���C��N�1XV�&�)$eE\� [�3�)O8����Z�/�(F�^��dԄ�*���t^�%7��2�R;�򼳜.�A���V����{��|�q����0��\��ɡ�;e���I�ۭ.R��@l6�)K���ZDķd5���f�e�q -)�AѳZ,��A���t�1),��^�s3�+J5���j����+��dnr��Ynaf`W0�5��ˮ��\���k��j4k]1H��w����7=�r�(��P,�Hy��u�ҷd@.�d@��y!QE(�^�gb9oٓ}�� �zO��|FX�;�ɵZ���)]�؂'�΀>+�}��~�,�H��c�y�4܁)n���k
�� @���M�	M0�*�'�ˣ�&T1��n��H����܉>m��cܨ���Y��a�F�M�R��z˻=Z6kv��}���ȕ]�<�=Hw���H��o�Y��A�Hܺ��B�Iȯ7ʂ�f�Ɲ�#*P��	˞ W[�ڜ�u�^Q�D{ Λ��r��kz�1-���|  �r>� �� �ͤ	����08Y��R�<�|n�����KVl�u� :ܥ׸(�%+��#�S��7�ۤ =����]��!{��gs��p�*F��x����}%�(��_�b=��fgk���� RM:Q�H�5��3:�M�u�B�e�߾�UU��� �2@>��x����F��{o%΅AIL��y4�+dD\��^��m"O	�NV��@ڴ4ȍB!X�؉ڼ� �m�H��׵+����a��wcRe~��*�9�(�u�����g�o;�F�*6M������+&����@���G���P�	
k~���k�y	�ݐ_{Q gDN�ݶ0��"j�*�`Q1J�_"�B޺A����(f�7"�c�(s��{��Y�Z���?�D�V^�أ/"͛��~~����	Z{{"�H����9��"o�!���j�2)|FF�Y���:�#��L��L�M_e�G�za%2�t�����|b����:�>�@k�}�C���V)r�d<�F�iǒ ���>1۲z�#��x�q��^C���2��_��v��(�y,=Y�#dj���}��$	�O�*&Q�N��ڗN��K6�E_R��ݬ����0[�2����*��Լ�%pB,�ԛ�?}��:n*�ҷ�(�g]#�{�.�̐�j���� J�7�2�>�{��G:�B;�_W9y���,�UQ�Nq���d�w/�=����@�d��PrJ��7�V[���@��͊�e�%w{�o]�"u��uD�D�3+mN�>�{ix��B�T:�Z�Zج���cj�crd�O�a~�6��?W|SʺHwccc~;w��
ȃ	y�>� �Y$���*�03
�,(C�&��s�ש���Ř�Ic���%f!%m��pXh9�`&5	ti�b�ƚ��W�YMV�nki�q��*��c����&�g44��d%�Qr�ij����WT��3����PR�7QYmf�ʲ�t]!VXUcDQ���o�|�BD�!t~ ��AI/Z���P�I��=��b�Bj&���{��YןH_$ ���o��}y��vj
T��AI�k�Ζ+WI�j
�$A��\��UG/�G!��P�$��<�"�[����{dm졻��(���.A}nhYݎs2w(��$m�D�붑�\;�֡���~�}�#���Ϯ�2�H�?��x��Z3rV#��}z�WA�7�͒>7�(�;�ֆC�D��wI��fy���*E�'��g�<��D��}�d����3����d��9z�tuw*�޹'��Zj������5�?	߾A{��G)�1�}��L���g�"}�@���r"z�ג8��	���h�J$�n�a�� ��o�Gǵ�I=ܛ|�C��aT�]ج"eB�����9��g �D�ς�P��>��[<�jR�c�-KWM!mلչ�i��W/�吏@V�j�6 ��j�f���o���w��u�̺P�F!X�Ӏ����ռ�H'Ÿ��n}�W�R-`f{�H�GMtI$���?^�H���ʮ,�Z^KQX�X��F#�bgv�=�91��.f��8�ڞ��l����	\�|� fn|��$��|�Uת"f�vg�r��:������/������n��t�{�-�(��ob���_fs��+]7yB7v��Ի������SQ�D�LG���sU����3�UQ�LO��͊|{2B��m��$_\�cUT��E�D�����C�ʶ}�ӄv9�G'b�;u��t8�	�[�t���#�2�y�!��/���se@p[nOW��=ڂ>�� ��PQ���B���Kl��\��|�j�Ҝ+Yx�'#�aUo !4sU^��M�,�Q�V����<����uꈙ�%U�����LH�� �X5)"Im��/�L�x����7h�Ϊm,ʷe� g6nv��*�����6g���́��%x�_D�����^�Yb���)����+M�5�w�P_=J$Cq�e�G8e�%	JP:� �H��z��ͯ��X��f�@����R��&	�}Ol����ª@`�w��I�������/c�z����C�� 7�\�E��;�� }��F�y�����UA����ɜ+�U�7�[�A�:��B=/q^��pb��=s]F�[�9\���f�LF[nzm�x�ƴ�]��Oly��h/Ѻǀ��x��{ʃ���0�����x�1�,��[�k+��u�+�<{��Ű����90��'<_o���S�x}:9��7}I�۾��=�$�T�>|�*Q�qpE�;}w|���6G�ᣕ|������x+fvh�@a���3�y��cZ�kl�Z�Te��.��ҫSs7ƥ��=�{ӫ�������'_��z��=���}G�$0�;��ï���L���W��:2'Z�v�.�9.:�R��ő7�ɬh˺�E�u�6�����[���o��|���9o��=@��q�o�^^1�S�����Ϝ���������o�Dx�f����yf>c�3��i~���lݺn�9æ�;�ѣ���wg�l�kq�����n������ �5�R��=���Wh��zO3�J@�����t3��Q���U�<�(YFA��� �x�UE`ŋ�*UX �O��j��DUD�iDDU�Q��
�TMYUV#h��AUEUEbŎYb[QQb-�E�*4�DTEF"bU-��x��X)l�1�feұQ�(1ATr��Aݕ�6�k%�]�(bi*�-�V9J��b��غ`b�郕@Q����*���8Ȱ̪�1�l2ܷkt�`#� �U�\E�E6�9QECVfh(
*�Qb�{�Ư#����Jgu�y�6Vc��P���!�R�d�)[I��6Z4f��ʉ�E�x^t+.��Xй��k��T�a4r���3�l���G�kh�l�e9�ƌ����
�fV���2�ͤ�&�3e-H:��vm5�Q��L<מ����� Վ��Z��ҷj��%)�'�x�v���j�%�7c+�d����49 �I� �],-��i��\�"�� �`�ᛃ��)�b3YR1��XjY��ݑ�,���),���aA�9�t�ַXݮ�MH1�V�^aK�ɝps@����%���r�I�v���.�ʃl�+��I�h��B�ʎ��)�+�͢쫃��{&��V�R�Wu�â�F�;@m�al��A�Q34Z۸�.u �IX.�<H�m.�����+���[i�F���.Y�Gn	�y|�6	�	�6lR��[v*=4Cb.���N�b�����R��i�R�Csn�pcYEn��է��p8GGXk�2�]��ɣ-e�M0R؍�U�A�W���vv:��Kə�]�CJ�Mk���*��HA#]f�%�Đ&�mP���V�fh�V1���[�2�ˑW*��U�"����lћ���n��fd��K���b���.�$��bP?��W9`�,�2�0�&Re�WmcV�бՊ��ؔ�-�Ƭ�j��e�loX�*%�)ECk@KΦU�9�;uH
��@l��M�ldcH�1Ҭ�����` ٣t�9b��0�e77[pʹ��,n��78´D��l��.�j�`�5ki
�XКZ�FGRg鿟�n��S��[�� ��
�:��$Iq%�
D(��E�J�6���v >7�,̊ �`Q޹���SU%7/
�@��� Ew>��+�� �G��z��"*��l�_y��lt�>�� �eC�z�DI�+.Ɣ!!�WT����N&_n����I�/;�##TFq���	�����цMVi���&�^t�>�*�S���l�᧸� Fw* ��(޹p��Qb�$�I[���ϯ�3J�3����C_l$b���A�$�J�'c�ì�bٛ{��;��h��D)������NcH��r�%�7Vp�B�*J��H��ҔgNKsi��I���}8M��&R��v�d�@}����G[H}���#=�sCp:�
�P<�C�F����I�KHk@��u�.��?k��������y-���۩Ͼ���eYk�����ou/�H&�ŨD�/��z�!ӄu)(;�z�@����re/"�����u����y5쫼��2�Wfv� CȒA$U֥y[�@s3yZ%2'��]~��r����.Ç�j�������5�	Y���xv��$�l�	��ע�*$�
kż��ͬyJ�%KH�K؟NkT\7� �[h!��i�J;�A�H�O��7�gs�s=6�ʺޮ�;[��AQ|�T��SK-4�ơf�kn�?>Ͼ�A�����$��$P�5�o2�H�/�Oe֐�$"ߍ�J��"{y��Qx��X�S���4�R��OO]����<	:�#dZ�apN#%��Ă�2T*J�{����l+�/~��!����+%K﹉�L�=��&�l7�=����Aa�s�Ǽ���o|��R��}�1��`T�/|{�6�@����F��.��r�����ZU2��݅ƳC�H ��e�{ZGwmL�#[[	��={pFd�^WW�x{��?� �.�3haXYǽ��:�.�q$�����VVJ��޾0�6���>��M$7�5�R
AO8� �Aw�^y��m��w���G����.������![5��5��mM�s������\8}�~��;���1�d� ����m
��w�lB��u�~w�A���;R
J�y��>��h�N�5�H,=׹$�>{�޳:���1�Z��)����+,d�:�̆��=x�k9��3'�τ�zB��[�	5Ǹ�:eH,9����
Ұ=<�}�t{��:�bA`tԂ����t��Z��{��m���=�.��8d�{��<�o����s'I�7�Xm&Щ+
°�rI�
��X~�2k\��]>�Z{:�����O����X��[� ��y�i!դ�Y��w��竸'(/{�6�+(2VT��2Ci*%B�/��$	��狾�wm����Z��p:�G��'�����)wN�X��țt��\�PU��;���y�%���[36b�
et8؈�"��+i��0�)��T��FT�eيƣ�X\],٢�ZXX��Ul�y"9c�6W��h��Ώu��B��MsI5�"� ��cJ��Y��Tf7ҙ��Z�Mt�r�m��3hYtR� ,]om)�1��l���d��D �x"<	܁��Gރ��YX{טm�@�*J����`i��w���*C�Mq����`V�|���P�� a��4�� ����s�\�bwϘx$�%aXVs�CI&Ь�<��O��@�rг���z�|_�r��:���X{�p:����ۉ �Ho;7y��y�=��	N9�$$�}�bA�7�au��q!�Mw��6wo���Y1��;���A@�V��A`hjAO;� j�ѹ�����O�|���H���)�[�l�{t�2VVJ�IS޽�4��]��o�q�:a�°��4�R&ӏn�4��YP(�=��&ț`�??=��O�E�j��r4(�"*�$P�Kf4&X�֣�{z��3C�9`z����H)l:��0*AJ�S�|�4�+8��s����܆�
$�Q���0�
��$�S"W���$}H�O�6�1)<�\��4��\��$:[�BY�VM���+}Kzb�����zNe	�s�� ����{��J�R�-��cM`Xԅ-=��I ������+���( �3�^�!J��da����42T��S�:�4��V�a�<y�o���+�� ��
�z�1�C*AH)��6�`s��;WX�Y��Aa����Z��r<ԇ���}�t��(�S�}�4�@��%e���
 n"�ұ�#�� n�H�'Æ^��f��r�S^s��H,���>w"�����n�Y q|ۙ>$�-8�I�`V��~d6�	g���ﺖ~̄f���J�ٰ�F�f�jE�n_߽���j�`;�1����d�Q%N�� �IXX°��rI�*L燎�N�2l��c&�Y(ʐS�}�4��ƽ��ksC�9`s�^u���B�B���<ߜc���y`V�K*q�8�h�����2H)��������O��������h��*�Dz�N=�q�VVJ2���r@�Tx�'o]ۙ�	}�b�ì��A�Ү�λa����G�,�F��u[qP��!4$��ُ��n�I���� ԅ�㞰�Z��Cߏ���b�;	�AV �0���d�XZ�z�FJ�T��!���aX^|�P�M�R���O��:�d�T
�=��&�l�f�讱ֳ\c��=߹$��z�1 �z�:�Z��p� T�p&�+(�Xs�$6$��3��|���o�}�f9-͊��ZS�n-�*U�w%f\�}��ۆ�Cu�8I�;�����YXs�xm�@�P(����cM`g]��5���Cv��I �C�}�m �������u�+߹� ��=���pJ�[�4��V+
{纆�
M�X��2hR
����őd�Y|j��L�
�>���H)���c�k�qW��[Z �;�x�#�O�(�T��{�1 ��޸��fF�$�"��@v2�����2<	�m9���T��3
AHjZy��]��F��5��Y�8��lZ�ܣ�L���o����N%�.�2,�}��3��`V��!�؁R��>�ԷZ]p)��x�1�++%H)�=a��C������$���8߹$؅ID+%��c&�Y+*J���i����=���_�|�a��m0g0�4�cl+3E֮�_�g�ǒ�n�^�Ѭ9߸v�R�Ă�SH/^��6�Y���89��m=�Y�6$�V޳i�aϜr����9�Ä��S�z�؆�++&�����]�:a�����H)���cM`V�)i�~`� �0+�<{�<㾃�x�r� T�����xr�*q/��3Q�������6���+��ys}��^뎡�AI�
�y�1 ���y������;2�4:�-a�9��'�ֽ}9�C�H,:�H.�*N�� �AH,�O}�!�7���w���OD�ACL/�f0�
���xu��.���
o�p:Ci ��p�͠n�8�s���p�Е���Ă�R
y�8&���C���Q���^�P��.^����OYP"��Uo:f4dn=�U�
�mK��e���7��;���ǰ������m���mKLm�n�#��75fWj)0ݕ*�#e��T�~ѥm�%̸�i�ðj]�
�.��C�F�1lRYy�a閶)`:���49��p�u�f��v��3*Pf��k۲�]nf�4 4�����n%��B$�4����EUz���>�kw�I�g�^��s�J�2T(�����i���O�7>�G��7r�g�	3��{�]���R
��^u��m�x��>5�j�5�08kw�ݤ-�9�Ž��߹����R
AN����e+}�!�6	*%B��|���ƽ�H,5Ϝv��պ3\C���T6��(ʐXs�xm�@�P*V�������X�R
AM{�����X{�&�Jk���[×\S�K�9�|u�Î��I �~�iV�a�d4�b �T�{���;���AH)�``sּ�+sC�9`r���HR��>f:`U��5I��R����؁Yc%e��^d6�ĕ ���a�����O=z՟��$Ve4�j���7 \ݡr��������}r�g
o�02z��YX{׸n3i�`>���X�>��x��7�p�Rb��Ci�
��{�楺4k�9Nc%��Ă�2T3̻��޳�o\{��E�۰~%�a�����7�3lٿ��8��B���� x~�>{ D+>=�i&�*J!Y*_~34��YP<��vp��'I��ێ�WY��Aa����B�B�`>���Z
� T��{�^�g��z�R
Aa�d4��*%B�����@�A�˽<bB����$;����߼��R�7�
%@�X^�$��-����fu߽k��s�u��)�C]��AL�:��˭�S����c4�R
$�Ϟ�C�<=�}rLH,0�<�H)6�d�_}�d�ʐP(�=��L�޷��vzY�)`Z��J�h4�G[Õ�40ݍ7/�Ͽ��s��N��<�!�����=�$��@�|�����g>��~;sYԝ�q5���� �9�H,:�ysZ]f�7��&���z}��0�z�i��+������R
{��H-�o͆�S��y��Kth���9����4�R
y�X��J+Ժ;���=���瓎t��iijY�u�N�]��G^V����s۫��C�;��{�{=2l��9=�D�[z'-�m�.:ǽ�������=ܱ���w׮�˹�v_>U���E�}G򛽃�������&#���o���h��޽�{�+����7$���w�ݔ?^>}z��4dъ���>�Nʲyծ�ݨ+����
���Vy���\��=�w�N�!�t��Bw�#��{��̪F2�︥�c��\�����ʟ�����:��'��6=��3�}׽I��>��X|�h��%_�L޹��ȯ��<G^
�#���}=��l���W3ؽ�\sӚ���k����e��=�Ew���FtF���K�^�_3G����﷤�ڇ�=��Ս���鶿O^}�����in�@���;fpA8p�1����q��e)� ��k]�Wx�����R1�9���̻��[0/-�wM��yϮ˅1����DP�,�T(��b
7V�2�Vҭ�:J$�j1����*�Tr��TV֪��"m1�b������T1�\d*
0EI[
��P����e�c+V����� Ċ�E��,�($Rn�(��	j�F�R*���"�B�%�T�F�Um*��ֵ��h���
d��KJ�,ZZ����,�+DX6�Ul�R�Z$Vؤ����aR���Lh�PF6��T��D�)a�U�J*����(�����Z4EES31�W���]o�0;I�B��VJ%�|f2i����J�/����|���fkZ��q���~�vs���~�ԇ����sy�� �@��`M�
��YS�}�m}�]s�{�f�&!�+���aX^y��n���qRs��=`lCi �����6�{z��ǃH�X�bA`i�i�>`���
��k�b�$Ş��ϼ�\���(u�e֤z�ٻ(���V���g����r��+��z2VVJ�T�0�M����ߺ��
K�n����}�8d�.��H,�P(�7�M����<2�4:�Z�^�i �s����o0k1��`T�JqϺi��T��rCi*�A/�~�[�~��t�O�>|/�[��b�[�$�
�{��6�Rz�!���X��x�~s� �6Zyט�H-�
�<�̆�h/���Kth� r����3ϻ��޻�N�FJ�S~���m
����CI6�G����O�~����|��|�c���U{��.���nE�=���; z��oܺl֭93a�t������}T���&�m�Oz�'y��j�5�$����B�B���1 �{�璹߼o�
AOu����Y�u׹��@�|!�2G�>�:r{_A_L$Tʒ�4fͶ\��.��66�*SN��5�z��۬�3^ä��S�z�4ɶVJ�Þ��pf�(��`R�ԟ ���,7sc"�T3�ķ}_+�&'4�� J)�$�q/��3C%ed�<w�l�;��:I��+Ϟ�H)6!Y(��34��YP9���{���qǸN�l���3�o�-a�y�۴����Ϲ���
��>��|��9N�*AeN��!�6��D�
0����Q�aOy���-�.��1'8��;><l�2�Q�����ĨJ�y�1 �45 �^��g�\y��������Ci6��G5-ѣ\�߹� ��p�&��޹�|�E�C
��w��M�*J!Y*^<�d�+%e@�S�|�n&�O�����_I�dg�։�*`�̣F�H�{�,��Nuj�0խ�y(��M�G��I��J�W.��k`,�:l�  u�6�ݚ��A̼n��Ԗ�*�T�K�a�.l ��&z�1�u��R�qFhR�(�`#@�]�*1�SP��P�[QL@t�Z��ƪn�m	��5�e����f�9솶kR�\�%A��
�� �gk��m�}���l�s��:O_��
B��|�1 ��N�� �Agr{�����!���(Z��3.����v}�!Y��G/&�(�/Z�72}s����O�j�(n��C�(�j�m��:�ͧ�,�WI����W�UC����=]���
��nt�H�巅̓l\VyTY�*!I*;F�*{�t⸤h�@���Q�nw}��j�q�R�$'#"3`�Z�؎��;/�y��qEW��t ��d>@��nE���pp�aW�z� G{��!�U$r��lh"o��ĉR��/2ksr�Eo���N���`f������=�yYFI7���P�O��}�� I�~�cS��0'�t5��e	W~;�!x�4$�E\W@@fz��e.�����nm�w=����l�D�� I}a�3�����ľ&%�B�D��O��[�W��Vד}�����ۮ�H�haQD��n���K����<�f�����c���L�P��TA�#q�ʖ	>�K ���r��V,2���ݫ���^od"|w�H�lD�N{�72~���Tt�Y���? �kY��"t��	�n�V� �{3�NI�i����G�7�&=%���ݮ�ܹ������f9\w/�:���>��wZtFP�v{0@�{5Β	<�I�&뢻�ay���渜�p��u�!s6)ڌ���n�A�T��sd�qH��ф��KD�1�8@�����d�e����1�|���c��?���܁?q��ȹuyfe}�w~-87)��"vE)�0y� �^D�A�B=~:�Z�'^`�0a&��Hw�"��skn�P
���ڑ��u*:q�n��J0��Mf �no��&���?o���=��/��/q�����'�4e�0%�^\9���[�����.�����IϢI�΃��;�D�x���꓄�.$�i��s����dLAɐ�6�a�ζ2�"���Z����u&���no�sޥn�^d���T���&b�hb�k/���v�)��	�d K̊�.Ou����C��5=�ؑ!#��c��b��|G>K�y���z�CQW8^:7����t��|ב�#'6V�O,AmA|bT��P6{ �D����ːSr����$���Z؞6����Zr��yz�]��\�0^���n�)w]tA�n��MtAo���v�n�C&)���3�����멝�.���jC[)^
S[+���*�X���4[��ms�\JV4�]�l�[p��,���I�MJJE�;�N.m,�:�l9�GBb�3�6��ҵ��u�b?���<�Z+|,9&��)5rY��]���0�
U�����I:�+�E��s)C�ꀲx��p�xҾw_�VwU����� [����9��;�wɑTD�
���H�]�������7ŗlЄ!*`&�D���(Kp�۩�-ˁ���H���0a&���Ax�0�mt�R��t �ʯo�����+XII�ЛQԭM"<䕥p�u��*��'�}�5��~o7�	���羨;6�ޙ��<	�&���Ӡ�()We�A���x٪8#w,ˡq�Q�&�<���|���C��8\�{_��yS	XΛ��Bʐ1�Ē~$	�����mT�/-��ąJn{��ͨm_v�Zt���-��A��k�ЂD�8�΋�+���c����H����rwq�+�{�n�Y����R����݊]�.�B���t�	�� ��'ǋ��W��]���I���*C���),�f�Ǧլu�]��|����O�%�O��G�����A�"�KىP�aE��%���f����Dn�D836�QAJ�;�(�x�"k:;�c��=�p��]�8F�G�x�����;��Z�7�}G����e������=���!���6uG�#*b�]��㜹ݟju�I�/�I���!{���{+%=�HH��3|�$��Ɩ_�=O��� �;  3��Y����&Y�h`�*]]!�ƍ��˗�~e����y��7�" ����j�6� ��H�oWhc�*�1����p��V��/���ȀcTb�g8��eq\U��D�B���I!�I>"�1άm���E�X�R@�VR��p
=s��DK�>7� �O�k7�%��s]��r#�p��LN�+�����nQ �%����.ۛ2#(��ޱ������ٍ)S�t�_���2�ns������(��Z�{=y�y_����>���v���8�K���75�4Ζ鳆���߾�X��0fܠI�>$���#�m7��u���3��z�Zv)T,����PE[Uȁn���Ȣ	���M��+��r`�M0i��G^%�-��lʧɀ}����U	{1%#0�6��:P�C��$����{R�1�0v�H�̸XRHP_%��z��:G��/wt�cj��J'���/J��ff�v�t��� ���jC46}_g�|����K�{��e���χ��F�p'=|���,z�\���{V罕�S��5������x�|=od��y)�w�r�j3��g-/��2�����9��e�!������g�����.&�����F���Gw�u'Ӎ��q5G�g}Ǳ�>�Of�tJ"%�j�:;��&{��H�Q���掋�ފ��������d��o�.TL�A�Ы�h��hB�WG���<��{"��5�H�%�ôx����&��H8�j��}�J���y�맴�n����n�xo`�t�L9o,з\�l�l�j�@%��ǈ�-Yk���5<�ǟ������{�zz����Q3ۃU�M�%�����sw'��z������+����-bwOE��5��]Y0�F��~�������<��Ӕ��q�~��w�~�s���R~���E��\#���'=�w��5{V䋰B;���NG����x�Xآ2[E"*)R��QV����0Ɣ��D�X��*�J��*�"+Y++b�""�JZQV�*�[[�0�J�jڲѶ���b6ԶX�Ze����c�Z"��-.7����4�.6�[��F��J���6�v�b��1e�Q*Z�-PT�Q�Kh�J*6ִc
��)��E�r�EAV#XV1ueb��Ah)m���֢
*��YmiJ�D�V,Z�b�-�k1����7�՚Lb+3v�	��+m�l��[X�ZPEX�TU* Ue-n9�+R��-���E�X���x��L�����h�k���Sh�$�*��XF`@��p�����v��f�	�6�u�A�%b�Ř�tĶ	�FK�
+[�$�6���lҥʀ�u���Ѯд����0۳�m��p��.��j����)0fe�ƣ��Υttn�A��&�6�UƮ�if�� ���L�i�R$�4�Z۹�3og�J�	-
��V�K��3�:'=���SeBg�ՒՆv�A���[IM�AH$�亄�d)�� ;^Rݬ6�Θn[̭�k��;\�Gu�Vږ�\��,���:Y��n\�1s��ŕX��q)0u���ԭ�Ա�U��E#tz��a��٦��b57�Rb�����&ؘA{	)�#��-]��qbh��ס�Md%�Yi4��R�9/l1`j��0Hڣ41,�����G,X�XSmk�M�e46�"�k�M�bVQʂG]�7L�B4њ`SFG2���1�n.�˫rBc7h/��6Ҧ,�5�(J�%i.M�0s�)]lZ�6��LF��y-�2X�,�GgufĢ�c+�Yw-as�v�.ĺ���a�m;[�m�Z��%���@*��-�Te�jV&�6��a�`�cfWgKQW*�Uv\����d�R4���Ԁ�]�@�3-�a ��n�D�02�Oĕ����t���ڮ��VYX�.��=6�f�,���Q�6��	RiK��Z�X�T��/Z�
���RSj:�X�
�V�jͦe��(�v��5�u^�Z@�a�F��R��,ь"j@.�	�M
g�q�L�hZSLF�ȗ ����HVٹj��__g�ڹ~=��s�Pܨ_Y�Q��S9�LϥE(��+�K;����YQ{�����!�W@x�
A��	� Kz�%�몳xhC縣H'z�"��We���U}E����̖��P�H}���v�sU�{ݨ�ڭʪR�Y��E�t��ځ��i��d�ْ A����r����Tr����n*�QJ$�����7jTe�����
�T�y��w�#��e��8��wjt�r�S0�uGn��gd���� ����_ؼ2�;.�8q�12�dF	�����{y	~���D�$��6�;�
���J{�()&@gC'��á�y�>I���_ w�I�hT�)�@�w6������ ��������D
�ޮ��vk�A z�\Y��3��}[|���s��k���w�:c"���T�5
9[B�@96 E�|�Wפ������ ��	�}�нƧ8����[>@�ts/�"H�S�.�n3��XGĒw����U��N����Tʙ�hq$�m�	z��y�GB���<x±q��1���=�^�r.�,�jfV���[��y�I ��'�w�\�ϥEU����;�
��)��|�ĉ7�F���D�I��HȈAL��Ԉ!�A)["s�aWA\����w�ۓ���!ur2������b͝��B�e��߳�R���]�^%��!m�V\��$���ڣ}MJ)�fm�zgw��_qD|7�/	���>�^��p�"�i�R@�Wg���A(5�<fv��n8�j�	:���(��1��:�dml|\�=|�!�d�����ȵw��ޞ[�� �!�0�\E����;�,F\d�=����Uk����I��"2V���W����T}n�E
�h K�H�_D���ֻ.�P@ �5���d;<h�u��j��9�7JC�:4��g�� >���&����'*C&�P��fb ��p$�	f�����/�H�A�"��p�Yyy�ף��(Ԍ<�$
��s9��������}<���]����`�$�u�>��B��=A�A>[P���!��>$�4����G�ê��  =�I ��s�*.`t�1�|�\-������h)��D�+���1m����޶��R%$�x�>~�t�>jY��73m�����m�%ch�6M���']�"�
�p���5�m��UQ,�-���ڎ������S�E�a�ҎuY�s����ڲ�!Wi��kK�&8!��ג�b��)�cے�\cL�L<h�31�SbdD�HŴ��kCRFMA�a,��Gz�������}����1Ѓ}�{V�n�����p�8��I��>�����w{B8� ��Ψ��6�l<\�f�0�v^: Fo}v mjuJ���ݻ�����#�l��EhU�_F�l�F�';fv���֜R
%P��^��_;�9k���E�I �����|�=h�����=��Ȱ�6�j��a��Kb1�Kr����lQf����v�UI�D�dglӍf�A �ﲨ��?)A	��-�r��]�↾<|7�xa!�S'>��O��7v�f�]���0���-@�>��D��"Nqp�Ի��@����(迍�d�=�P�|�kiT�����^�xSc�*��N��T4�yTA's�	-�uD�T�3�MP��ܬ���P��Hy �d���ƽ[B�{��p)�%��l�?X�eR3�#I�-�#�w��T�ssO�T�:��=��A�ʈ ͉;6��@��T'ϵ;+jE T�7��GSU��ڰ�T Fk��÷6w��&��DО��$�n$I�z�;�EE�r��6h��t�8�o]޽˜��	�z� ���:rC�����ۭ A/�z�P�ah��":��DORD�]ğk�[1f������̳1�_�B{��cN����Wo��r|�f��uezy�,�;^MIR��M�Rʷ������gV���'8���Dzrm@u�H79��,Tٷ"��A!�Y�e �U�M��=&Ƥ�	��O��!F�OD��d����!"�2�e@`�x��HW5<An$��A�U���BA���"����$E��M�t+��ݢ�s�.�����e�0�����nO:�X3y��?{yN&q�/�R�1*�~��s��� �
$�T�!��t��$�'�U	��>�����������"�%�-�Ø��[��{�Ŭf�=��ok�$m/��+t�A�mP�⠨*J���!M3UY�xMg:�5�أ�!�TEfnD	)�RF%]�OU㏒>$���%�>x�W���G��fT�wB�#R�����}�P��f`YّR6w��K���6'���N�C�7��uV#wd@-�H��|���Iv�NeӦ�"��|��&f��E��/fӐ p�MY�6�ߨɕݬH�\%�Ƀ9EF��0;JͰ�-��-�6�v\�p�]1�E����P!)�f�T�CA40]��M�Tu���u�\V(%�h 8�0�5��չ�ephP&��U��j�ZL�\8V�t���ᙨ�x5�F8M��٢���˴332:��]����ɝ��)t)/���ȀF뢆x�b[�P$��Uٖ&���q>r|Y[���FwdH�5���۷������l��G� }�t �����ssX��:�y�Aܡ�"RF%Pn�q�Uv	.� D�A'��^x4M���QFa eHڋ>�m\Ѯw���P[����WT�ϦfxW)0Ķ�GZ;b�{.�31D�T�Wy�J(D�*��	�<��ι9ۃ^j�,�m5S0��5M�+�P�ٯ`�"�w�[H�#SZ��#��UYѴ�G	�ѳћS}��ޙ��W�����I#I����^T��7m�u��ThqD�Mk���]�
�6���D-� {smY�w��FJ#�v�"����t����B����͋)��C8D��J�-��H�sѨ:I�� �M���t�z����b�I�M��i�T
�f� Sb��Sꢨu=��(S�)vޠ��]�<����\ֳ;}ݝ^��� �(Dؚx�l�)�}\1FI��$�ͯX���&dC��b��)F���Ds� �&��������-����w�2מH��	�\�.{ڡߩ��{_�&�ڬ�G�p�ؾ��7��ghG8᭕��\��W�_&r��e,m�L��Ϸ�u�ɳ��]��59���jx�=&�tq]��{������ѨEG�}�
��}���2]w��_�Z�w%����
Na���D7%����"�w�y9^.���lV|ķ����ۻ?JV>�"��%���d绤�s��YO�n������x�Ѩ��=����_�'bG�x{�/��u�W�`��}'���z=�Y�!�]W8�WHv���C������d�ye��XmH^�LRBJ𷈧�n�k��{Le������s��?g��~����O �sV��@�X7��+��а�]����?z�-��ay�k'���/jc�j��W]|9�ه���uJ��Ͳgd�UaxPd�T���G;3{l���%�3{�w�����v���e��,g(�Y7Ӽ��Z��>�����,L@�S^a�1C.e\��ZΓEEt�W)EV�Ŵ���Kim���J�6Պ��.]8��KcIJ^��Z[[�@���^�a-	e�X���\/YH� �+i&1%h�RҕER�R�7j.Z������YkX�TFZ��\��c0�m��E
�.V�DUhر
���iU�"�mj"�R�AF*"��0֨���D*R�̦*�"R�`�s)��[kD2�\%%im��V6����*"�U)-��M�3� �	H�	�����z�-QF�i\�cl)�d�z���&��$�_���'�|�.�0F�O�kՃ�>9�r��_���@,�oz������_������Gh�\PoZ��xw�R={��;��B3]/���O��|�b��e�q3�dl�7V
�U5��0����˕.q�w�P7��q$�<�W��*�
��(��T�H�PE�z���~n������$7	��x�qw�G5� �H�"s$�� ��<�{Ϸ�X!�A.��2fPR�M�S���D��@} k�m^Z�۰�x��9]x��Fe6���m!»jlv{���7�*��,􂎒&�|=�����d}�����A��$�_ٵM�踛$UZ@�Ǥ��S��=��u.��r�Ui�C�'+B��M�@w��?$\��Hp�> �w�Q�8�=�&qZD�Nb�H̪��hP������r&�	6�
�H&D���Hz��S�*5�����B*9�g^����$��l�B`�֕o'lU]�E_��@�Kת�m��y�y�D���w���uQ9Sޝ�R��^���:B�u�^>m�U8$`ֲ`��s�(�n�{�
�;]���i$�/=ܪ�u5=�U�XU}��H?{����A$:�#Jֵ��3L]���e��\غdb+s@v�Z��C�;G���c6/if5��ʛb�ö�pYb���l�)�!��@����Vǎ!H�1�Y�6�-t[�75�ʭDn�	Q���iI�īi��v��d`T:#6#�6����Ͼ���(��|s] ������R��٭B������_#M�J#�r/=���M\t����� �c�h���B��H̫�w�D��+Ė��;IG��yw�6@�˲⊣�x�ץ�� �����"A���f���	.��^-�&�f�ӑ��q$^s��5��A�K�	8�|�8��v徺����{�AA���ҷ��;�1XQ�WZt�M��Sm�D�����72(n�,P�{��iwYB�$si�3�0�vm��F�x�/�5po���}u{X�4YFX����]��@ދ�D,�t3s��b9]ΈBo��t��D��x�>����n�-ʨں>ޛ�(*J�<�Pz�	�x�6{���@k�ӧ|�I�A��+3�a�U�D�ؐ}���r�b���$��H��TQ�A	P6��&��B�D����� Iy�����������}�z�h�=��sxq��������yj������D���5��/�H$��uG�Mk�8���D��4""%��i6������@=�'ă��yƫn6q��w�1DDB5�=��מ<<wW���k��n/z�no�v�J�N0V𩫊g���[sy
������٦�ͭ�W~�G'4�v m��ټ�IQE��y;�}�9��>��mZ���L������$�pBI�a�͢FkAOm^#xj$�Iz�^#[Bs�r{q1�D���e\�Y�,��Ǖ-�Oq�"a%@]|j�j�[i�3y�p�}�VĂ	��x��0e5e[AzX�2��`�m�Q�Q�'o�V�j�m�	+�Ĭf�Q̪��Q/y�Xn쀳��clqE\�ׅ�GF,�]B�Cz���=t����'��voM;x��q|�ٗ�5=�r����)N�E�����L���KE�/��}��~d�;3.(|(~��f�l`$d����D�fN�F�=��=���y ?� f
�yZL�pc�Y��wׯ����Z�_�;�B5�I�+�yq�ݞ�hA������*qEQݽ);��,�Mh ���Y�F�v7�v+j��;BbaA���$A ��O���ս�ۂ�v�����l�m:�!h��_g��^P!�K�ƙ$s�UZ���Ѥ��9���A�����Ho6�iu�TC�H�,��Ϋv�:gR����qsg-F�5�A�yqS�L�}<��Ut\�F��ȕ��d%Ց�R�,��}������C�&f���Q
m�.�BMt�+����hAr�ږY����B��jAu�������7!em�Sh�+K����Z4�]#[�4)P�-����1���G]qu�����#e��S-�c*j�[J�J���:YWn���F�Hgf�\�>���Æ�~��~���ڣ��;sd�d�8m�JP�We��8������p�$���	s[�2vm�gVR�0��6H$�j�==�n�V$8�$���ո��10��YO`�:D�B|РKmD�wV'^��/��c����`g�)��p��cv(�$���^m�1���eM�7��Mڤ1^��!z�5S���n�3s[lqEY��W�o}+�m#N��p�K>�n�U��ʒ���ɤK�<:#���w{8�n��t%;��a��Dx���&�N��<�G*zrnMA$]�W�r4�������Ԩ���#s��w"�&��k�8��˴����˔��Gv�$�L|���HB�l�5��ȗ`��v��*ݕ�!p�R֛�&Zu@���$�d�-E�*,���\�����$�е�Mt�V��}��X,�����}�0�e�Ç���B7}P��Bi�d��ﮝ���H��>�Q"1��:F
u�Zw0�*J���.H��,ψ&r"�[w�̀��muƋ��2
B0�8�u�Sz�X�����f�m]���M�i�zV>c��}��a��W�UUS�v��ξ�`�{�҄#��ֲ�K�ضEt�HQ0�(��g�.s6���n+@�l�8���ݵn��wn����|��m&��Sm��U)s�0#���hZ����� ̕q��B:p�$�;[�;���z����5�A���$D���۴�\D�Ǔ�6I5d�m
5�z�c��&�����QNaà�o�X�H�Wsw������k�;�U(�Gf̓�����>kϜ�;J. ��)��A͉���I���
3���������J���fI��ӿ��]<j�⪜�6�k�I8�)�y-*0h��<$6��������޵��UQL�i���Rcr �cvįjll�y��m8�z��T����V� m�{�7.<e���1P�O3%AV%�M��&h���7�۰=�Q/��bk�Orr6���N{'P��߲��~������g�j|��i���ӂ,B�"F��j�_jD���*��a�W9���^w��Q(�͙ ���T���΀o�}=(ϕ�o]�^�s*�F8_���|YjUrE.��x���G^_BycC<g-��-콦��Q�A{���{���'L|��
ݝ��v>�"x�w��p;�4߀�˥��.h�"]5k��v���
Č�ܨ/ܘ����=�!�d�>9���힕<�v�	�/��H�&����^ݎ�.ڇK�.�%D����^$1S���������r�7*�����N��{v~�/����Cr��_�����(^t�:3~X��S���Vo�\�n��5o�ٗ����<X�����ze~e|<z�y��o�=�w׎��3����y�y�7c�ׁ���Y@c�-�+}��I�jN��S�i�;�}G�����}����(1������]Cz�.��g�=��#E�����I���vo�w+�9/Z���x����e�=�xh���o����c�Y�c]��Oc��/��j��b�b�����v\e�Ţ(F��WQ�zF�x��-�	�6���u��x{��<�Nk|�㮫�S��f�#KL�J��r���J,ke�������Y5�Ņ���
f70Řʊ�����Z*��h����ȎLiR.�N�E,DեqY�Z"��E��ӡ�DA��-+Fڋ\F��9�G*�F��&
�l��SY�Q[[m��Lm-�m�Z6���*�Q�1
u��TaD� � ����A�-Z��[f!�ZfTV���B���"��+zU��mil�,��(^%JK�ɰ�d��e��e�E1�)�(a��d�u�дFд�P���l,	N�(��Z^��|��ǳ0�13��ie�H��;j] C�a�%5�m�v���tX��̖��3:&�H\��6�
@T�@����-�`3eJu��6.�A0Щ�2��i5%n�-�҅ �],����ģ�;7-�� 5ʖ9����c8,fͦ���XY��h��#�8�:8������Ґ
U�����Օ)��d�6I���k2ՆcpB3l�!�lq��6a�e&�F�Bʼ҆adl�*�x�)��KM�l�]�Y�5�R�"	-����Y��9L�3����&��YvM4#�3J�N�i�G9FMvY�\G�p]mд��36��LM�R�Tc��%]7]2h��]�a�f�y4��vT��L;)��h��وp�l͝��6.X�KQ���-�gKJ��	3�h�3m��hX��a5t]mv���;s.v�I�ĤE-)��d�*���/.�Q�ԡ0�EJZ�.�/&��Vi�h�&um$P�ƷP�J�I\�E�ݳaX�hBb�R*B:����]Yuɉ��36��� ���mbE�����jvf����#CH��z%�WF\�n�� ,��Rjf������������U���WeUUvQWcV�L�I�yt�5m②).����i�1M(�n�ɘ�v��6��r���ڍ홒�Mc����5���k��$�m[r��ݝ�@2؎��6CT�̰��Ĵ�f�1MZ�Xi��e��:1�F��Y������V&f҆!�1�vn:�X;,�`��J��\�ƦG6�X.3�v��fݴ�tC-�J�}��	��w�D��HK�d�V� �/�^>��|��B�Y��K�ݻ@-͑����¢��7Z�n��LI(+��J!�2A�bG.�7���{��z*Y����DJ,�o��T'|������n��[����2�|�� Aw�D�Ky���d��;�ƹ�lGo5�ã1C���[�XE/Q�i�kiY.��ݵ��W�߾x8p���ؐ����$�Nkt1:��N�$�fM�d�	�W���]�0��w^B�I��i)�D��Kz���9΍ۼbi��E1����!}��.Ɓ'c�F�t(�x���>�d�t�qڷ�P�گs�j�i
��I7� �^�T{Z1vU��wu����(|Nm��ͪ�r��CHR7�����Ys�,�ϒ���l��I!Ƒ>$O�
=�Q>�ߛ�=�;C���%�$!����l������%t�Cge�Ϟ�RQK���w��fl�K��)�) �������J%ٛqD�uϦ�K:I$�ܪ�><ܠI]����'����D��ָ%B+0���Fo�" ��/�ʫ�g�؎�>2$��4!+6n�8;��o~����<YÚ�:x�f�隚餲ڶ}'o5{�Β%Њ���v��;��gpWWv�7�"8f�3ܯ�1�Q�V!vU�D�Y�'q�t.��P$�9@�K�g�{������=�^�"DS`
"��� )^զ����8�/��}�h(*K �7T	}��,�AEH�Ƿ��<��?~H=EуV,R~�0�������
$���D�gŉΤ��=�H�%IP5��,�$��U���˫Wd��e�27;�4J�&U�n�ٺ�M��� ��H$�Ӻ=��x�Q�{v�{x;߽r��4W��ŀB��l+ɽUsoCf�,�Ă�Њ��!ETq�	��m���{�e9Da� �Nki8��8�Yɵ>1�2��\9�(bD�4�j��-Pw{��R�qW��@Xt� ���۲�N{r�3����#ǊA���H�E�U�݆Z9^��}����zP�f�ݠ�;[���� �;ӌC�)�,�k�T	4�rђ���$�����H�%IQ@��j}b�(��I��TI��X�0Y��[��BeU�w�B��P�c�D(��jЃ3d&"�ߤ��r�t9q�ݳ/s�|�i�^��a���
����WwN�**w�ߢ'����ɵSZ�� �V��6b�!�bT0�K�![3�Lq(YV��.LE�6�s�f��X�&=e��,e �Z0�B�Z��tMu3�:��]+�H)5��B�X�B��K
[���	�h`�]�pj��YSS;J�kX�e�ʦ�9L���r
�D�>�uS73\#��~ �}v��i��}�q8	� �|����*�x�fN�$�\�u�@��u9��c2Hu��I�9}T=� 74�7�u |N�b��wd@��ӌC�vYQW�s2*�KOj�^��C�s|�.�g�muq̲D�
J���D�)�?w��l3g�Y��@z}�;xNU-:�b��e'���T�+L��B\Zԫ]5J�w��Ϣ}C2����A';�"\3$���X0/j�F���;��BeC2Տ�S��&�Z�ҰM\P˥R6
�W3�!��<��yatJ%u�j�9-�s�: �ޔI�Ȑw&�k�5���0PU����:P /��ޛ��C�� -l���-%��-[��^�'�4�$�o6+0ɳgopX%��� ��س��{B�wV�<�B�i/{v��ٜ���\eD�S���c��D�!.u̲�����}	R���o�@pGۙ��V�xE[H�Y��8!B*���Q��}Qsh\aH<��^:*,Wc�1zڜ�TL!
+¡�>$x�Q!K�Œ09������ȷ�&:4�˟��ݽ��ṝ}�Sѵ��+�;-�z��Z�Ig���N>u[��(3B]�%�;���$��'ʹ�� ����	άt*�ȹ�D�?^��F�k��{�lɐA72�x�����1��A��o��@&��`cja�iN�f�m��?�~�{HV1��o��~j�I��"�}WJ;��P��T ���Zr�)M��*�AיU�Im�	&�an<��dR
�w�(�1�Q�W��ڂ��ա�d˘���8�SY�$���|���E�꺶=�����r93`Shrؽo~�Z��y�FBv�c�*�Ω��3��U��(3vS�@�^@�����f2�<�!�I-ȓ���ch3�~��ݕa�9F�a-A�4ۊ�UP�:�;��ȅ"%	��l�ޔ	�<�I��cd�`˶�{(�<8�8����A"�e����,�*!����y�Μ�	\�sx�R���-��A5��<�v������	��� �&`.�p��u\��wI	��p$7�ܳZ�M�G&-�s���㿯iR G3�2�1�r��k��r��Q�s^�Y�F��.�ܫ.���}Ǩ�E���g�.������~d�4����jD����ی�.a�)�!u��K01cm������!e-�Ѭ[h2��n6]],�i��^�iu�L���b.�؎*�1U�Z���`���u �ev��nj�tA��-�����2ۣ�b�ɒ9�7)@��eɘ�E�X1J��~��"X�y>܁`�H$v�C��0-�_�#�@�H��-I�.�z�5{��qCfi#�I�ᯞ
�.��}���5ۆ��!5a܉��W�L�n_�#u��G�w6Շy�dr�[[�;L= �窉%��g)�>Y��f!@�~؄�M�p���wrJorv�(fI�m�U%�H-��U�~��+Z�ִq����3YqU��^������;`�7��	���H{�e[�����n��v����S�����<�D[{׬ު�B�ؙѾ��>�m�V(q�w7�k޵�� F;u^$�mz
�z��P��C�B�! T�3Zמ��N�eJ�L����,ݐ/�ӌU�,�J^+{뿏�r@A�O����L��v|g7��Tt�&H���c���;���$	OI�|-������j���ep�e�t@��*�ne��n;����"nu{/�`#�� �JH�T�{��a�gv,@�2@Y�x)
q8��gęnN�]�=�O���ő'��j�DC����
&!IV%��>�"A��''�|zC�4��Ye_طt��+�
� G'|~�˨�A��w���Y]�F�ճ�w�5�Su��GV���\�R�ç}�U�y��vN�[Jyz纙k�~�=5
gg)��0\�}�炎Q:$���^z���w��j\��M�����p�xaW7;Ǵ�c����Z�J�/��<��X�sy}�8�H�S�A�vEW��5L��f�!�Ǘ�⽩�3�|�^��0��{ۏ���9K�5���`�|�{'oZF޷�ʧ�׮�T������\<�2��d�೉9��}�C5�CW�7�g���9�����ә�����΄�nY���'61�=ˊ�ކOE��\E����[�{6Nݧ��o�Ƈo��	�]vI��7ϧ��Y�6�=z�=�;��/x��'f�����c���HsO��bx>x��� �V��/D@vL�X��ٮ;��LY��.����b�?pĳ�IGFbr�J�qmq��a2ҵ�)�a�.RԂ�؅5�!ᓤ�
AQq1��3��U�YAT�KİElx��y��[!%�Wc�mmP�J��B[#z�ز�kdma�Y+r�̦ ��%E\@˘���(�DAL��ˉ��73w��@���)z��b�!8�� �<K{^��n�ލD�km�%HKŒ�v�Rؑ� �UnZ�Ƹ�28��l�TZ��TkW2�����E2�Z��m|	R���l3!cy�K�q�֬J�Y-,R�Q�S�(c.!�f���1`�1&e4�2ؙk��7���{� ~?���B����]u�O��f�B�J@�o{�Q�&�[Q��8��w�d�T
ڪ�q��	��"��P���{���SD��RBq5�,к�5ZP�)˰-�u�����P�Z�6Y����W7!���+d �>^i�M�p���d̛����At�K�kΖt��C鮊B�N;�����fϧg�����$	�� =����j:nQ/țם�5d�>>�Тy�K���LỨ����|7G�L(�E`F����[��G��%���~V�Y��A@�="��';���ں�Y=�K��	|��>��ysr�y�<�R�����V.��ª8d��"�UI�o�hN(��h#��Z�m/ɽ�pȒJ���]�)Q0��&��9����e��j�I��x��5F�L���(H�+�mN>K������E�i���� _G_�2��dkA�`��G^�xQ�$�4e��:�S�4M��갢b�bz� �:Q��'����œK�Z�Kے|�Jo�;��;�Y9����.C���{��.U��7��=����b��>z��6��}|(��O�\�w[��d�~m|/��l؎�,��U�p��iDX�,)�	�Yp��-��l˕�j���[R[���V1�k�@��e�uVܐ�6�{kS�	�i�6�Qv����6&Jk(&��^*僃W`r83X�[�X��sU,�	�WR�X�\�����$
��4��y�J�:��Tʺ}��hP6�EgY�BM3Do�f�������I�>]��5�n�ʕ8�V��8iH�wؘ�k�DƑ�2+9 �T�*���JA.�UבD ץ ��~��`���UrB��Ϥ*P㆜@������Q`�IY�$�q���u�5V	�.`e�n���mi3������*�T�fꎇ(��L�P@�:dA[�,u�3�}x)RD�l�-�@��Rhӧ^�c��jWE���|6�[��t;y���_ ���M��7N�����ܳ7�����%[||���NG$��^>��Un��"�!7}g����O*�D��2A���2*� %*fQi˕����$qF|A�"��z���Ȝ1ЀND�$
��H(�1
�{B�$洄U�x/<L�"Hw�T/���;mmD]���*P���\m��X�9nC0��:�Ңm�����Jz��_/��V��{=&���$���uaD�RU�O$X�[Jx��
�yB���^�F��ǲ��慤`!*MOhQ��"D�ݺ_~pa�������h�n=����fS���I�9�Rr":�]_��W����-Z7b����BqA6����������s� �d9��v�j}���W��Ja@ֱ,�6���z9r��3��8�8�0v�+(���>UNg��Rj�K	12fV
%LB��u�
���Ipȭ�uS��y���PA��y#*L(�T2$�kO��q��ͅ���5�����+�˙�-GD�r���@>4���Un���� 1�w�rA��P�n��#�wd8R!�<��ֻ*(2Ģ"�O��.�H��u��=�۽u (q���&�u�3�w��5^c�����BM`D�O<չ�Uة��C:d�I��
Ȯl������弔�F�UT�)	���mL&ڽs�e�._~}��s)Ư&�0T�.�v��Y���q@�dHٽԂ��!Xn�i����ϱ�"H�n�ٰ3h�nq���FT�Q^�� "��,����-ݬ�����Wc�
��UeS��91�ĔY�O��s��nl�b=qt5�y��"R��4�^o�V�R�<Lę$�O��[B/T�.���Ê��gz��v�qVeLw%qq�|�y��c�&�m��7�j!�
�b �1"1hş��&���V�'�0��.�ڬSjQf(�Tf]i�fMoP��i������������Z�[d�d�+X��6X��h(��eΆ6cV�PL��,��WK�qU��z��,uۨ�M3he�q�]�v�K+7P<ehV�ٙ`]pV�jr9��m����} �QVag� =��؅�����=��)�G�|��Y�IN>�n�A�s����B>	��V�>��+m���I$ns�o=Z�b�|���Dm����7{v�Y� wk/�JpҮ����]
�ҁ �ᖻ6t���X�Q���IC�U3� �:Q~��]��{�{v�m@��J#|~���"��c\�aeKtcB'��ڪ�T��N��f3`IB������D���ˈ�5~0ݯP�i�#0�!&�;�$1�L��1x��u<T��3�ze|�I7M�s�vŞ�=)?\�|k���«��^g'�I�� �>>�-��oE/
)%0��w�I�O�����(�9ϲ/uJ��T���75�*s�M�-ȓ�m�20G��(�>�^Hʘ�	��}v��$�@ɫTl9��I.�	{Ϋ�v:���lԴ�L��siX81���JQQU��߾F��~L���}>A<��q����!Ƒ��j�H�3M�n���6��$gĂN�hQ���݊o�7��!7cb���Imh�Ȓ'�c��%N����N0ɞ:�2T�F�* e�����q�1��c��K�W���W�9=K<ʐ��l͵^˓zQI)��L��dA�fH$�^��J��ݧ���LC2M��IID+��{T	�ie�gUf�� s��۵ξs��f���#z��h�:��m{
�Q+M�V������S0���O���I<܊�)��\dY�	yyT{`P�
ħ��Krr��D�A|ڢO7>��TKMčF�رp�F�庠O>H����.���wn�3b�c�8ȝ��|G�Wˈ����mD_�����@��Y��/;ݦ8u#љY!oyv�9��""+"��^\�;/�J�F�Z*��^��wz�^���	$�̔��R*�wyV�w��a�l�1�Hͫa��}m�㚰2��n���D���i�1���c�Ͼ�玆ͯ�`�������(	�Q�f7&`n������^JaI�QdX;�dJ}I�ix�,����n����製ա@�&�O�8D�O:��:�R�+���P �2����M8���yz����$� @m�\���I���I��s��
��|�g~ E����{˽�sN�B.܊,y����}��?�*}��T���!hH��� ! ~��!I�H�V�0Fq�
h2�3��j��/����h��ׂx'iI��͈7|�CI�Ǘ�I	,d��(RO�����˱������*�6K%���O�d�$�H�'����:����IH}p��=!�J"d���B>�F�ãR���rsJ�3�èR�����N~���|�Ý�4�!	����~��D��� 	'0�!	� �̒���Ra ��a�C������(}���'���H]��O���O����������$i�� BA������C��C�� g�?RhHs0%8�g�!�=�2�1��u�[�L�H�W�~L>�~,a�����!���q)���?�e !	:>{,�2o��m1���D�}��� ! 0`pt� w�Y���NY������rh���������~��>Rq!�������!�	�����	�?3�B��c�/�grl>a��}s�	�I�O�������l�����������S���@!	�,�xa�?�����$?�'��@���
�>a�ҘOYa���������a�"�O����~����gē�~��?y������@����=}���"?p~��rtuà��@�y���B��&�D ��&C� ��������A;g�0��Ai����$��N���d��n��p|��!	����	<!�꤈�ԟ(������d�pN�d��}�ě!����H0�+RP?p<�O8�d��%���2ZC��٣��_��A���<�����Od��!�I$H��g� ��$C�?/��?������<�?���������!���A���j���D0~��$���y�0�0�2?l>����������$Hi�O����� t�������A�rI��?L��ԇ�����!�$��|O������<�Ù�?�t1d&?���|���o�~_�g�'�!������W���C��$��>��Z�0�q$�! g����q~��� �|���c������������XQ��N~�/�Ѳ�(	7$?O���F!	�!�?���r������������B@� �O�'��A��~�N!�ǈRN�|����3g>PX�0��D��������9����"�(H%�� 