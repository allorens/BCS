BZh91AY&SY��(��&_�Rq���"� ����bD^�| T����kF�mU$�b�l���e���[a���i��Jl֛fM�m��i���J�5kk)e��"����T���j�&C	�ZU����Em�2͓mj�me�K,�36���JiB�*[3L��3kY4��jk���YB�ekFcm-Y�����V�V���(��J���uU֪leR�;PNZ٪m��y����J�d�V�m�@jkk5���6�ɘ���kb�Z��ĭ�3
�����f[��cT�e���Zl�S   �>�^��8;Z�WXM@:7e]�����wj��@4��gGUC@���*�3�i�mQ�a��)֭�ե��m�ѕ�HI�<   #�Pz � j�X�8 4��  �wu\P]�mv� H v��    ����N  t{w�X�Tkj�V��j�Y�e�\   3<  h{�p  �)�F���8� g.� @���@��th� t4�ٍ׼�(�Xt�s3&J�Dĵ#RPjT<   o ( ܽ�O@(x=� ��W��z{�� ����m�(9��  {=� E�  :/W�� b��
�����15m��!�   �� ��Ά� �� ��  w���4��  P�������p h{�@�e����;F�KU��ڒV�����   �x ��mƀ pz� ��  s�n� �.�@р
�۫\  4�:�� ��  ��!I��-�*l�Ҕ7�  u�� g�� Pnp 74 K��h �8� ӹٸ �]�[��:	�\u�$.F  wuFڙeJ%m�kP�ڦ��  �� ����F`�A`�U�� �:V  n\� ѣnÀl-K j-�˩��+RJб��E4�7�  w< k80 e0 mS(���v���� ��0 r��4j��su(�Z�b�IͫZ-��Y��  N� Pݷ���  .v�4�]�� &6��r;� m:pM�\  �� ��P��  S eIT��@    )�4b��*�      ����R@      "��	J���      $�5b2)�1='�z��@��(mM�J$j�R�h�   ٻ��]�D�]vQ�-1%���;���YV-��
�L�}5��f�Tۀ���������\�������H�
����UU�**+�,���������/��;7R
*+A�$�k�����bk�A=��""+�����U����cb0�b�L)�$ed �m��k85�5��gm��k;md ���p�`��`rv�g,� b�`�,��dr`,��gm��&� ���!���,�Y9��;`�lCmdY�C�1gmgl9�Ŝ���;d�,��1g`�Ck&,�;`��,�8ɶ��v�gc@Ő���v�Yi��0)��*��QK!������� �C k (4�E� ���SA)����D`(�0R��)LA�-0PR0R�
)L T� �Si�*4�QJb
�0
b�`*%0QR�*)L�(!L,��gY�k&�@��md�Y6�@8���Yv�0Y6,�9M�����G�ޫ�G<���/�AU3������J��"�8���V����ʻB�p� s�B��<{&w�E �a���)��	I�j���x�1�5�D�w�*�P�|��yO��l�h�t�I�Wϐ�E�"U��B��5]]Ef��h3Kp�#>�8qd9E��U�6���I���#��d	�Sp�;E๻�PVS�t�.�c�0e,�t1��BtI�x����]�D�ne����krj9�tP�*f:k&bj�����)Y�nme��5je0�M	mJՊh�dZ��|�5�[o;��.Ʀ�q�����Q���ōn�3v���= 2�\�|U�{t�Qw�#z˸���R����*��%f��p��CFFŸ�YQB1*mb��qD��[f��)�^T�\�0l��	א�%��'��=��(q���H�4֦l����Y���S+\psa_]%�l�N��XLG�ֱ�9[���D|$4��cֵ�M嵋(Ь8�����t"si�)۬�Ӯ�phr[YD��I��6ʩL�77,$:tH��JK��U��C���&|��2�Q��b�ˤ�.��ۭ2���<���)���}� ����DQ�m�+h�e��#76��N�F�������:qo�lW(4�p%4V�fЫ֊4*�S�^ctbf8�DT
�v�e(4�j01�����&�s7.���cBf�Y�m���+Ś�{R|�lXN�8ۏ�/�ŗ�š�D��f��2� �ݽ2[�3�C0e Uf;7M"��۬Z0�˽�F-�Smw������	�}ڈ�·U]���\U�8c"�V���J6��h� �bE ����i̷�)���Z�EXI�.�܁���Wj�V���T�U���9�nWy�8�z�R�od�-��3"X��&Ӂ^������Y��GaAW�!���jf4�dån��rb}�k���h,�J�=��31���E9��̉�j�!�c[Mު�c�NU�sd�w5d�$�N��HV+x($��ØC�. kM�0*�W0��g�jַBD�H]%�R����W;n���V�\�q�F�;�0U̙�Ew���jG@�+�Ytin�R���h8'�_{�.���Bfs���<�Z�R���cR�zѱ�~�3-� Y�rr���c�#��h�A歧���2��|U�œ���)QW���)��,QOq�����v���sbx������)�hX��Pd�,�3^��M�;�te���dTk)�X1��'C.��1ڸ�c�Q�ag*�5޵�i;2:#5�[%]��w�I�I��m�4*K-�^m<U�5ۺc�YV�����(8��~$�1-�[,:[�ե�Ŗ�x4�����v��B��`1�ŠޥY�2�T;�Äk�z+�km�T�,�e�z�80c��m�`������Z���V9f�J�d��S�����Tkv��[��,
�
�wP"☂�%����pe�J�Q�a�X拢�a�okU�����J���q����sv�b���2Ab�B��"�U�M�+m=b�o�ICOj�Vc�p޲��.��$�g%�UkTHGVb��!�tCX��6���3`���Mͬm��F�ix-:٣]�E����FV
��4k��)�G��Ayr��pLm',N��fa3c1�)kR-*�ܽw����ȈWAի:����=�Ѧ��.��}��!"3]nҤ�3k0e?�	(Gx 8��̋f��X���'#P  л�3f=̛cC�����lc����ff˧�2Ѭ6AerM����P=ո�I�#��D�-b�MÙ�f^㛂f؇0L̠�4�757gma ��\r�25P�RO�h֬E��L^���VmՔ��[�]5b��I��ԫt�2f'X(6��
f�w�؏E7wJ�U!��M3�
��(���E�^�NF���E-�:b<V��ܱ	5`��g��*����E�Ӗ�uhRܸ��k���:��Jx�^��;0?�Q],SV �+.ձ~��U�r���pf�dދ��պR3T���Zg�1��3Z���+9Z����wV��*����Y&�Y�J�ԛ��E��8Ip<�[J��-��Y�v�Ƭ-ųQJ��゜�r�(�1�D�˺u�f
.��W�&�Z5^���S�3$"Ќ�nUИb5�zH� �U���.�J�a`�զa�Y�l�fMY�k�h����̺h|��k�7��-.��W�����R��N�Ѕ�av��>���43,;�$��J�D����5�Ve�PfnHi�D%��b�ܭ*k&mͲ48o0Vn� �n�Q�	A�&��)�.=Te��2�d��K�%�2�����˫�F#����7�*�cV�r�$��c��Ų�*c���!�C7��m^lv��1H`v�$�{n�&����ҢosL�Cv�H�GX�e7�%���n�0^�̏����l�ZwV�W��I��+(8���@���AJ:��T1Q���R]���Zu�n]J;Ko��&CF�E5�x�t�fm�C]쐋�
i��#�B,HcM�6��5�\�X�]4DXBv@�ÔUf s@�j:V�j%�e�Y���Z��v6�4�8�lE˧J�-R�nm k>�0R��Un�����8x�k�t�E�ÛɊF�7]H۹��F��벲���^$�[`c�E+ñjyz�ű�1뛥^�-���+&���͋r�Y�,hq�y[����%٭���PY��I�@O.j%K�f<WՊ�$ƺ�޲]ԓ�_��o2-.l��#zj�dN��Wh�fky&SP����T��V� �2ғE��ԽA�n�kVP�a��\���Ǫ����#���n�!��@-�hKۇIb[HW4�۬.P�#�d��r�j��P�B�v�QFe�����0���K��V�o+��<dV�F�H �JS%��R 7�TWrΉgi�f��o�3������Ru���I'ylX����@d�m�dY86���[`��-���K1�{K*`�X��G/h�EAV\�5t��D,�j=1��63sA��w*;����Z��2�Ga���@s
�;%��fe�����C1h�(E�:�N������7)e�����nk,o۸���4Td��L詢VV+7r��i����C�՚nf�4TȲa�iMnB�9���OwN +6��̱Q�4���0P�kRe*��YfG�N��ŕ���&�I�֘0Ҋ�H�pQų4�>b�7.�X�e*�X�8\s4��tlKXa:�i�2��Q'����6��-�KMY��(��-�V0�B��&qj�j�֯�Jl��gn�/6]Æ΢-x⩦*�N5����3`"��jѩS��سp�7Ba"�f4ڥ��jT���a�ǈͱ5V}�6�ˤ���ugJ��9�F��qj��9�Vpv���{��"�,��cfS����h8�e-w�Mf�x�@h��Vn)Z&�%J�I�[)�(��i����������VBe?�
��ި��;�-e��cC+���;�<��v�>Pb���-eو7��4")���]cu�,��b���Y�!�hGlhb
U�����d�stZ�QkHګb	����E,@�j`+�NF�i6v!�<�lS@�Va��=K.]�"^�k0aW����[���{��5�2K�7O2�T��)���æ}7��kwQ�W��g�ř�%�u����m
x�٢�[�!����e�#7reܺ��ozVkG<ж�!��U��/��Z���7S�e�ȵ��۫�K*"*��^���$��{�j�#h�(���cwX �D�H��Z"�yKCy�r�s�N2�ܟ]�a��Qf�w�Sˢ�e0��%���6om�Ø\�C2��36J"y�0m���y8S:4�N�[�[��l�������r ��A�Hkv��7F�`T��SX�)km���Qh����bK)+��,\�7"��Ec��l�Fn֜EY�L����*�h-�z���,<�GWU���p�!��*���j5r���t)��KNޕ	3k�1\z�ǳh[Vp,qh����(+֜�X�Ru�f�X����,�,����Ѷ��f5y&|pB�I٭��n&1P��</5��[x�4i�����Y�:XR��o1�µ���u@�ٹ�7V,������H�����1�`�*r���T+,Z;��N�Ё�b�C@2��δ�XI�q�[/Bf�*sh�W�V�.�*TÛ��Һ�U�{F=V,"Q���ƨCQ�7�w�-ۙ(��nǃv�`F/
b�)Rpi���7��7U�5��X�;�ya�DM�Į�"I��Nnj����V��;,h�y��w(�F�H�2�Qj��^��>�Q�k.��v�.��.Ԛ|�����m��Zfi�/������l2h*�ګ۔�]e�`R�ո&�s]�.�+*<);�U/���~,�Эh5�ö���V�*�Ȁ�2��/U:�Mfv�GM�y���T��L{���&���z?:�����H�*���8�\�����^�YGhX�G��&�HU!u�T�@+�6���3*Țh-�m�[*��t��q��G���RVV{`[n�5�n��Ekr��7�ʧ[�:�nM�z��W��t�ՙJm$���j�3%\��0��'U�Q�
�xu��q�k�t��\0��9�e��xux�^��ja��	�V�~�$�4ͩ��b��ţK��¡r[Ss+~�r�G��c����B�R�5- �o+JŃ6��֪'4�r�����J�Af��;O>�4��9�:��L��s'�+m^������S�T��ʟ����D�hgs
��Y�E��QP�˒	7Q�CN�˚�dl��*V�ͣn�kA���᳉	H����wv�bS	�e�u"�� ��Ym����I� ��ue�YJ��^bw��U�=qb[KdU��&���E�(�zm'x(3�l�i�@�ìP�^f�o�����e1���. �`zz���M�� 	�X�M��$B�]T)abX���	�}wL�B܄`&��:�]���qL�&GL�W�πӌWe���?D^�ۼ�Z�gch�ʚw^m�y[R\J���HYu��Ո\VnBR̼�;2=��܏cɉ0��6cv��u�次��ݱ�&���IG��$j{�,��|5X���b���`��@��;��R�ѱ�h�&<�tq'���Ҙ�[��crV+��S��y2�HW1b:�&�{i�A���u܄�Vf`�3H�6d/+Cx���Y��u��Lє^&'�y�325e�T��^���h)u��TZn��+S�hT�͢�c&��wN'tpi��6a��
)K*�@��-�n��WL���n�ԨM����m��([;6:�C��pej�"������81���8�Q��F	c��h	��#�*�o׌c�Ci�)�r�@���`[Z�0��_5&%��F�H��݆���6�P,���w.��Y&kx��J��%,�hSGb�+�0B����˱q��
M���`�����:���C�щ�H����/]H�a�Tُ�֊q�D�e*4�J0�m�ɫsLm3xŃ�q[̵>wr�#Z�6�כ�j��ϴSZ�P�04�|ī�Bm�.
:o2���j�O��1c��n"�E�pi���!kx����ZՀ����̼ɵ r���[�LZ�$mk 
Q�ˆ�3S�j�i�^��3�*h�e�����eKˤ"�B�%�Z�l���*pFf���eޕ��O��yL:ұ'/^��H�Ux�³+&C��P6e%�U3Z0��Q�YXz�i�V1ֱ[� xJ���A���ے��e�J�۬u���Jl���h��Y�l"����Y��Z�&�(���;�A��[�%�$KM`X�R�9�5����Y�r��+L�vGX �ݚ�jm��{�ƗGov�M`�1�n�cJ�V����/c��6���E��q	,"M�+,���+Z'3PMe��ᨚ����Y��t���K��+��!����~q��U�SXM�7j�ICQ��,��j�{k4`b��]=y2�A��\�5�A�S��W�.l����vm���4G燎�k�m'�k��.�[�9�A�CX��V�����7x�hjr�Z\�m�Mbk��4��Y��� 7A��4镠�Ѭ�I��"����*�])1E��U��uso(��]�j��ͬ�ȓ\�^�����G>c3(�*倨[X�Gqn�7XLЛ�ɪ�;�&H��3j�T��V�W[K�e7D;�V�s3%�sZ�M�S[Y�-c 8�Ǹ@Sa=�	�x[���TԲ�}+�`�hue^,we6�iZ`��>�e�*�ƚbE��Żbj5$;�\�R���HЛ��9�
D[�cm�K!��0n�Zfaq�J�ʶ�=�p�����V�W�(w��A i�
�g6��u�!|]%��}�0��tt��J�A�H�Ln��EGkf
+33q�O,�t�E�R�O��Q�6֜*�O��\�� ��}HVU����\�&�u����S�2�F���4����^U��l8b*��v(��;RJ4���[�R������r�D��!K�S-�VZJ8�p��('g�Qˢ�̼�7(M؅q��w���Y�$�1W3S�x����m��ĵ��%Њ��hIv ��[�]bXcܥ�rt������8U�ę�Q��̶���&:����������+�����ݶ�y\t��C������1E�^|n:���O�K�B�P|N�3 ��U�ef_O�6Vo���=U�5���v'҈V�����1L2kve3��˲�*�	wd�pm���SJ�E+��~��Ec�ϲ����C��7H�hƭo�N������ ?��=?@C��<����Q�ʻ�-��7[��׷=ox�c�n]��RW"���']���d��KOPT�>5���÷BJ�h���g+�����8J� �Z��'Z��������E��P�d���oo�8���^�`Mf���XT���"�K���+�6�/�GU��cP�׵�����ޡ���ͣ1��o\|����ZS�������p�!΅wө&qt���T�V(M���6:
��O�zP��C�RI��9�[�z�,m�rIA$�DT�*iCVYܘ�8Cu;�����gENg�{�i�,���EOaQ��i_3����,C�h[��,�h�!q��$�P�-[��(�u���hf^d,��u7��/Z��|���[���cs�k{�|�b�FHI*ÕnVq��s ǣ�)+��fuu֢�Ԙ�BW#�5���vy�@�0)��;��sU�|^Z�Mi���l*�:�3u�f��E6�:8>�h02l?3�Df�{`�ީS��"5e�!ov�N� S,`q�=&����m
�溹�PZL�·5wV�E�\�辬��sq>{|HP�t �JRU�<��3�܈�7A�ƍ�jj�MIz*q"�6�9G�i�ҟ`yPuM����q4'`��:��r�P�@�{�.%��^�`�\��c��j�Q��:E^Pb��,Y��P����;f�LK��[z��F,SE&'Qx!���-s��=Ԏh�4�5At��]����=�tI�v]�͛ �o�!A(f�JT���o3�Z�'�R�G\�%β���Z�;�v�g3-��ݭ� k���M�>�dLSCK2oT�5�PK�1�`� ���u`8�u��6A��N��O<R[���{�����b����8����S�����8�y�m�>ɧb]�
�\��Y�ujۥr��a����;E]'���46IR����)h�u��Mq���Ǣ�w�s�]Р�k'<��+y��]b��'.f\�Q�T�h�F$	��ŷ�
�ApTk��b��v�A��7�,�{�X�*X�
�h��������`�5JX������R����t����ŷztF��JQ\4�V".�&K��cd���gH��8u�;w��ڨ�ԁ��W�'Ov�'�.�H;P�e]�bB&�FHX�',����:��d@w���LQ����Tr�`
�Q����#��t��f�P�T��#��}2Ν�\5�Ep%����\.�<٪����yJ�(b�+g�a��.ei����L9�KYlqŝ�b�n���5���]�Į
Ad�l#<<s�2)RXp��Ip��Ν���-�-N찒<���Ӂ%ў��o+u�r$j3i]�"�w������er(��m�2�j�{�ת�Y1��Y���d[�+2ޥ4�r��q���/��U�siT�7F�H��!�:��S�\9��/{���P�K( �h��Lb����뚥*�������6gRd]ޚ�Hn�ս�A���כ��]����٣{�*Nm���RU��Ar�uj�r�r�O ,b���4v͘�ܫ��>�*�Ү3iJ������Qg����4���N�b��9�i\�LE��;M(;^�I�e\�3[����P튍F�T�F�'qn��,���Y�h��h..���ȎuG+���F.��1gi6����w��B�1ۭ�&����'�ط�K7@L����u�4kw�3��l&���v��#n+�F���B����m٥[���1$�ٮ�tj�Q�=H̴�B���P�Y�d_��HF�˝ϫŶ#����I��-U;U��a��JY�Q���NB�K�P������w%��͌J��_LcC�t�ӯi�H��m��ŗX�չ�� e+
Ԡ.��Q����t
��\��v�jL��A8�o��a�]�X��QF;��.���h�A��n`J8y�i�0Bt��!�˚�1`�ս;7d�:����of�`�s��MVvƦ�Q��{7a��+�L�]�9G��wk;5.���a̗�8㕦V�t�"��EF�v�7�K��rb��P��m��"��]��jB��zTV�v7�E]�;�;vn��fK��o�;�����݋�j-)����a�s�5j�X��I�t�=����� k(�K�{1�3Z���5�Fð�\�W1.q}	4/7&%]6}a=bTޞS�n�T��AE�f*q_���ȁu3�ھ�Yz�l�t�c@�� +V^n_�Cv���!/c�N�55!z��D`w3[��s�k)T�I2{H�x)�\���ѽ���z�:��K�
���r�|l�u�w�R�M�=q����Z�u��a����m(�����Q�6A�DX\3�gםՐ��5�֢v��m���<Vq���9;(1N�goY�j�G����\�ud���b��>�7��6j���r�܎��ox�x�tYiVѱG-e��̏^BԽs���]�|!�3ewH�]��f��e]�ӮfJ����+��md�u�#�<��:���`gm0�P5�&�,cy�η�ok]
-���vu�pW�I�7��}f��ݼ�J�J�365*}2�/�А^���V^4��9'�]]<�Dɹ�Iu}0�d�݋Kf��k,M��X����x��n�-񸹵gq��H#x���f�!�gc|:7�Z{Vh�U��2����vNoJ�����/Z]N��"�dkvG5l�*\=Zk�z�|^�4��:�уn���O������p�I�.s��K/����WA����E9�w��]�d���=�]1Y,����n$|��p�c�lv�9��s��s"�(�Q�|$�5�G^̬|3�>��K��Ċî]˹ܪ
8�3������tH�8��DV9vSD��u5���y�F�w��I�p�oheg7���OV�:ء3_�P�i�í�CC�S��ɴ1�崴����*h����7R�Yǘzndb�3]ڃ�B�
7'h�ϵ��z�1i�56dhwb���흏���mcb�w�X���o�v��e�K����vrkC�e���ծ��g<�/nL�O�nM��MR3
���H.����b���a�\���{Mɮ�4��>��r�5���4����w�ۡ�TO@�]t��h�ٴO$+0j���N宽�on��ֺ�{"mPǰ,��X�R��s8cl�GրRZ�TE�Nn5��K̠���ߥt�U(����v�q�(Ղ���l�E���x7ь�aڟ^�6��wvԍ����}�!yQ��tN�$cM��_v�˶�N=ߎJ��bĎ4�IIY���˷P�I�*\�NR���"5�f� o<;���9��w�j��[2s�B�(��L����;b8�4j*&0<'�u����
g5Nì�_j�Ck9e���2�R�F����Nu[�B�t���sC�)��c5p"ݸ�d�ﲎ�d1��{2���X�:�6�A�r�wH�ȮkZ]�r���C[�X�x(nN���W7�o�2)�v��;�W���2��z&5!yg�q��j4�;��$���P�<�o;!I�\E�Y%��z��.�+���;r�u��{̹)(�v0��#�I,�g��E�ғ'jL;�UXŗ�A;HA�wֻE�S�4`!�n�t�0y�0�2Q��Kf�>�AV���:��7�qa�W����JW�[��o[�jr��Z��t�l��%�r�t((�f�]�o٢b�Z�z2�_W�jM��d	^��h�Q\�8�È��`�+�8z*}LJ�N]>͖�:���]�>}��G���v*.Y���u-���7�ؓK��aWc���f=�����n�J=�7�ƕ[_#x�J�CVr�8�V,Z��}GC���3��T��τ�]�}�������Լ��u�kڜ�4�-����.��w_P���Y-O/Xqy�� ���|�6y$ף��vw	�U��\ S8��j;�y��E#�͚���RF�A�XR�1`�{.A%P�'�`ט�kGt�Z����3s�K
��N�m>�g��ͭ�ũ^�i�׆Ff}Wf�ܝ��%��VJݹ�] �쥕��i�o$M^����N1|:rP�	UA�<�O�vV�6C�n��H=��ה�f]w�-x;&�����e��ȱ�%���vb�gm��ZuӋCTO(vք������Rc���~90

n��f��D�HU��p%C:�"�aw�����i��d�����Dz�^��,�֒IX����s�9�>�'����+;c1gz�"
ELԂ�}n�J-�i%��4�-KWi�m&m�$E��~B�ȭ(d�����/����AQ�XJ��/zd��V�2}���-��,��v[u
v[�q�<�샗?�iNf�B�p�u;V����Yم�۹W.3��G�Ƿn��&�k�ᴡ��/J�Pp5b�)�x�aʌ��ΣC�����\��%]0���[��v�Q[�=�frL:so>�ۡ�(	��N-
A�-�����:�3�絷�"12�G��aR^�vQ�ko�c�Ë�>y*�y�b�E]�(�ip���,�y�u{�%��bRb>�4�QU�Jm�v��g(5���O��J���5u�]s9�P���<����t����콹m�vc��ԥ�䬫T��[3;�;���BfU�N��0^P�2�����,��{���T�0�ާ��WR{p�u���͹(��A۰Lوq&��j%˭����sV�.�\_U�a|i	U W���1m�-]y�䤰�Z��P���qM�1�c���s,��JQke��O6��{b"4���'��15�{	���c�Tu�,Γ!����T��\��Vf"�-,�{l��n\���Kre<lm�Ƣ:�o4���K�ƬF��u&�H�.�^�_�~p�醧*C��q]�Z5Q���>���{��z��ش21�
�&M�A��f�ۑ��ޫ��r�ą+���!4�ԉ務V"���0q�ۭ�|ր"��j�n 7j�FD�i0�'bM��9��F���#+le��m&D�\/>�{��O4�-�`)@�{*��E�J����Q���\�������tT2��( ��F^P*��Z�YMD7]o9�Պ�T��H�Bv��Yݚ�LG����m*J�N���e̻�9���;�6�{�U!�6�;3_f��fbw�˓�j�Y}���bb����Z
��t��~+��զ�XP!N�Vp�7a����A�O>�nU����� �L��cw�z�|��y�ZN�f��%uj�^ex���!~�x�u0�ʳu�ֵ݅2�D���+��R�����c�⽬�y�E{V�fN�ރ�AN;4�x$5��R�p\�3�a
W}�8����c����cȯ;�uJ6Ҙш��1��'vE5}�c 䵠������S �.��rg�� 5�a�${AR���g���Y�R����]�M]nRKi+W���5$K�qm��N�{x�8:qwWLN������(�I-���b��_=���C{FD;T��f�ۨ��\Vtf�5��G˝A���.hL����-��ԏz	`�x��,h�d�T�V��͆�m��aj}��@�:kp�*����V�����n�_;�&lZ�m�{3�%���]Ԋ���S�O	]���B���4�T1V� ����+���G���L���]�,Ꝏ*p�V� 3"�^A)��BY����������*�b�t �*���]R���U
�j��6�����:��鋬�o0E\��,�0��yb�)x�x�&v��z��;[�0Y�� �7U�7)���Ҿ����o��fl���N�woBMo���b5dFe{uX�B�]a�iÈ"+sy1��WM�:�A����<��a�)m��_n�0�SA�55:XtM��}�%R�d%�b�Lfq�ٓ��So��v�iF�Ν!��i��&KZ��Gc%�5�70a�KV�X.�՗8/9H:�5y��.�CZ�;È��D��Iғ��(��t�Z��@i�}s4)��H��:3��U�eZ���\4Ƨ�ωif;Ц"����sg]� )�*�ʇ:��2��xy{+JS�,�-߷+�Vӭ��/��U0 �������m��+�2h,���J��s9S�	�M!ot�Ն��C��U�aq.�tx��F��9ےt �o�i�]��Xw��8�͋��AW%)>o�;��o(š��{��mi��^oT����Am�����N�4ͪ���C��+��Z���byJ������9eu��IP|�Vx>-�/d�Ή�R�9e:���kz
{��$�HIK���)̺�r%8���^ ��e�{���Sn;yaRB�vo�4I|���mGZ��ܭ�*u�����hU�����O#����Ě��s�wV#fܑ@�7x��)���祷CX�pDf�*\�i��,�r:��;H����΂n6e��,n��t�淎��]��fk����ick'[��]2�O:��ә}M��Tq� 
z�9��1
]im%&��B��y���B��<�3,@���Ċ�����9ej̜��ln�F�U�{��*�~xd�qUa��r�6���yԌ��W
���0�2Փ;��J�V�K3y���M�WQ�`7�2u��u���:�N	���b��f����m>}���lC=͏�s���,\%��+
Zw��}|$C��l3�wl�/�W��j��]6�Ps��,�rnVfgH�Og7%�e���m�������-��I��=��d��RU�h�5V��5x�g�gno9Q	���4��k��:�e*屘������Ez���E�AdV����������A* Q��2C@S �S� +�n�� &�.�	�A�>!2��@�i�hUx��Fv4&�J��B��Wd:�HR(�!5F�Cs[	l0����YLL��_�TPp��_�ݚ � oծ��v��N�E Wˎ���{]��������kq�L�i�5�9l��I&xJ�b�".��S�f[�ܧC*pT����(�#	I�����[��I�ɛ�&�f����ɵ�ЏfJکBGf�䮬��	(�3�f�V���ۄ�����^e���X�,\�b�SoP�riy���Sܱ*_[&q��V��rb��X,ӕO�6�k���<�ِ�!����]h�*аm��L3$�%�r���LEJ��|'s��K��݉��sb�3��W;e�.p3�����+>��]�k�k�'J�ٜNl�vҦ����f
�Xm������ܽ��w��s�MaM7�24p����&R�񊚉D�{{��;}ʺ����;�^�ł7b�Xn�|�enٚF�V���*��l��9��J;��s1�ɶ�����p��`��0;�#�oE]��y�,ɡ��17�����z�9��ލ�Xr�
���6isq��X$�zke���H��n>E�]�y�ދw��g%�OT5,c3R��Z&��N�����$*F��-.�a�q��+wH,madfp��PFl�,B��$c�﵄N޽�b��ρǁ�[�H��[鎈)%�;0�zn����j�:3qh͑euё���ls��n�T�����"}ND��\y��ӎ�mʀ�R(6��ރ�*Q�p��6�����{���y�v��w��}�w���7��}���������}�s������}�w��������Z߻���ﻷ��}�w��|�w��[����������_^< ���]��Vj��*���,�!�u�����S����f������V�K��5�u�ed.sab|ޒW}��q�[7����x;
&]r����S#�`��r;P1C������z�8�����m���Gx�6�3�C��-��$��Jv#���a�;~�P�8��z��@s@����v�4������xoh�T��e��Kx��02���rl�99��2�o�S���IǸ�ô#��f�1t�; =����T���u�,"�n[���ۦ[��ckqs�I:3�ISwu��+����V�VN�R�+� 4M�&�bnq5r�L���aj6N�EONe�(��\�Ü��� Kz�ⓡ����}�BX�[�8Uc��8�p��էY�z�	F'.w�н9�k�W3�yxk-X� ���_5%���WAK%VQѻ[��)�se�\GBx�Za7;Z��qj�Z/S�X�����y�ȳ�T�LV3���>��x��G�M��i:Q��ER�W׻t�c��ܴ����DvLm��|�uk��Α��ļRV�.Δ�t�2�tJ��
0��֝������v�+y����ڂp��ΰ��l�=��x@�e���y�vT�:��A���F+d��7�FV�(�>�4�:]^ �M�C��|��<M�ê)�4�⮶���3�0�-�x�]';B���-�2�L�W��K:��>����|��?����7nݻv�m۴ݻv�۸�nݻ�v�۶lٳq�v�۷n�ͻv��nݻw�����?���GZj�;�/mM�`��o�+�W}Ӳ@�)��2]��r9J���l;�=���+��εD��*F�w�d�Xx�����4�bg���;�=s��:����)�5Wt�_wT�E���#����safk��n}�����a�S��e��e��Hurz�.��S��z�'�jyHn����]3��[[.�jT�P��)��V9�T�R ���4S�vqsN�]Ǹ=�˓slr4�Q��4�h���ݐ���סg�)r��زƒA�1KwU�TΒ�XfV�5�NE�����&�3(ի�s�v�5p7xWh�n�)9;p�w�����ӫ��W��݁�R/�WHkb��w6�u�1���w4�y�e��Cu����8��"p�=����HE���'{K�mYy�7
ғ����]��t�Ԓ��p���M��̤{7���dS����>�_}t�`}��4��2`{h�ͮ$�� v�i�rR�2�_�Q�]��b����5�]��9}�CI�1����0FLn4)K��a�U[)�*��O�P욦M��;� E�.vT�5E��@"�U�%����Z��Ӑ�*fm�s�] V�:��С�msLwJ�M��h_u�I���y�z{Q-����#N���wf.�[���!d�p���)
����0*ݨ(�:�<
��+��wx9�l�1Y��9p]J�zȈK81�4wR���l�I&vu1�B9���\�oYzJS�"�}2r�(��O^�;,��5�k��j=�[���
Dz�\,��w	]snL�S�X{jvm�C=�"е�c-t�	.��<�e`��n������uv� ��'m�)�r���K1�eY��s���À�4��7�Q#uf5\��;�
���F�]Ʃ5r��bۛW9�}u�K��\�L]��f�ɶGp&��2n��n�)9:��genIP]y5��I��]/_6����Z��*Z:j�b�n��ЊO����if�+q,����[��1�AV��Y�*�/�l�i ��Sl�ӎ]Z�2t:��BP�Pe��O^>�
�t�4΍N,76a<P�\������&��(d\oV�V��S�֒O<�[�_n]#>�^�����oaܦk#����.Lkn�Cs��Y��̌��t̔N�9b���;�s������6����~�ڍ	�d��ˍ�5��k���.x��k-N��z�Fo�L\��MD�q跅=�}3gp�"�lbP\Ց�i�{
�`I�hrN��m�b�\�_b��#� fSvd��{H�:���  e#c�Z��Z���\�Z�Qm�Ή͎Tc�*ꆅ��lS�ŠTu�mkX8���4�r�:�m�ɖ�)An�X���ܕw ]�Ue5���]v+��%2�ŖsB
�=�J�f�mJ��53�v�u΅�HX��wrwF�V�z�D����m)P@�g A�X�0$�3(�}�mh����F.��'*I�"<toR�ǣU���6���t*�t��Y' �x�A�P_u(^�%]m3ّna%�T)���XX	���+���+�&vG��r`խ:w%�+�؏PEXݹ}-��%z�	Bgm䙭#��lY�0X�+�W����3�����N6�
���P|t�G������)7��S�$s��Qf�"�A��lqK5�p���P�=�y}�HM�,��l�$ �#/�R�T��hT�]��=F���#�iur���\"	��ɧ�!/�Y��8�i�ӪXM��6j�ghҐe*���K(<ѡ�JIA����]@@��֕���i�b�6^tB�d)��2�s����`�c×2�kV���IG�K�)f��Ee_)C��������a�Q?(�B�N��������/�NqGSn�VZ$Tl�ca��%�{,���$�sfI���W�d�1(�C��S��d�����aT�˭S�a�'Z�Ud���-qh���ޜ�o�
W+Q&��L5HJ�ő<冞-�v$��h�Iڲ��r��]5�S����uݙuC�n�1뿅fԝJY�B]�PΎ��^��z���%�PeK7\��������vvl	� v�]^�0G��g�3q-}w�#��qv�9�Y��ֹ�GKW,s�+$y��.&�cOV֔F�֨=\,P�xkx��w��D2�>���[:k�"��r����ť���F����r1�EԻ�|���h��`���t�n�(+���36x�6S��	�VYT&�2��h ����3F4���MwY}�Q0��;�C$�-u+�D&���ϋ�tD�ڭ˛�sLCV-�=�.��-Z�f5z��kh�4{�t$R<�0DONKfƅk��=�I�B�+�gT�jU�"G.�����i咤 �G	��l�5���(�S]vM�z�+�,d��/7.�]�v����q<
$��Y�������w���!���<�ʴ(�e�]`�K���� �6���5����u�.��<}�C��%d����X��,ճ��$:�:xp�[a��Z�/hNc��Zh��CC���P!�,�;�������؛��ܛ.r���Y����-��>H�AA���5�!��;q�Ob���˝a���}�^�Yd��G��&(�
�XYG�$�X�YJ20�
S��8���/g*
��0�	�7�D-X�mf�Q�p�5�](�o�^ދKyo�$"�Cܽ�����d�ϗpW��2�P���µ�"�dt�X�f+��ɩKp2�zZ�8&d;��e���c�h�ŧ�-8+*�]�p\a�*Yc}B��Z��u��[��tӢ��qU�\/�v9�Q�n��O��W$�<����B(�9Z��K7����s= b���C�oc6C F�7�t��H�ٽ����!��K�.W�̲�N���5H&e���EVʎ����ɘ0Z ��p��S7��z
n��Oo3��Ι��4�e�zZV292�Kx�P�-���=��M��
����cp�.B���hq�ɂ�;(�b�!��Q����	y<dC]r����=g�K��MQ*Hܜ/���%N�6��uV*\ue�ˉ�Q(�;�}c��n���Qo`��9�Ӽw)FxJ��y��Ӝ�\���ZO�k�<�.@
��/�ܛi�U���͎�D>����F/��U��IS�^�$��y{����Ni�-m"+	9��nC�s'�feu%���P�̊��M��6[��{�9�,ټ$�5�P�q���4�b���2�^��ݤ��ě}�t5J��>}�B�4���fW>�:4J[v�:��`^�Q�;0e�Sh�t���:3vԼC�6ƺ�z!�$2���h�)@Af�
�1^*F8������r�+D6oCy�.|1b�zn���1����D��s[�M )G��!�M[��+�K�b�T5�K�v�+`����ɛ)mDP����r,�t�W�jK�������<�䲲2>`+kr)��]\�I1=�כ��	�]F�2�Mɐe���e�y�L��(�6�-<N��M����:�mb��&;k���Q���l����\��xd��E4����ƶ�j���3h�dl�9�@Kr�dm����ḉ��&U�CBl�:7�;wc��q�u����Z�w���LӮn3�7N�dt�c�� W^7�=��#��,���E�zTK��l*���~�p0�f�r뱐@�:��������Z�:�U#�B�.��JS���Xs}��v�|��D[��{f���L�X�ĝ,�xOb�(������^�T.���ݬ���z0L�$�;{^]찤�'�35^��t�{�l5ǪY���]1*5ܕ
��9Q�2�_��%�c��q 1�ۀ�*鎝�k�=���.H�u���n��*��Pv�r���JJ��3Y��4j4����!�V��7��|����Y`��YT��O��Y����J�!,j��b]k�̾J��ڷh�ڹj�{L\�Ӿ��p\�3 �8�Y��UIV�*�Rq5]���27�Sbj��4�J���t�˔fw%�z�9������0��z��[�oV�(���M3xr����k�*��5���Ww]�tGm���Dȇ׫3�k;��S���E%#����cf����4��S3-T��a;���:�WV��5�X�яh��h�n�hՌɛKQ�QP�v����h��%uf��M�/�b��im x_d:yvX�,tk��SR�:ɤx�&�ꭇv�xJ��ؼ.�>��+g���>ˏ2�R�v�a��D�ʾ���I�����rm,��7W,`l
���&ҽ���Tq�bzz]�Rs.��N,BȒjn�{��sN�M�_m�jN�	;܏X�ݴ ��f]l���6�{�V3��Κ�.���㺼�HmJ�]�Ŝ֭��p���n��p�"+3i;�*o^�T�o���P��B=]t�Wk�cyJ-�ٻ��s��7�ɝ��XX�1��@q}&�2��/��h�)F�V..ʧ���ӕ�%��n'�v���6��9�qNO�^(����$(�����;O{6��+�N�NED�n��������['q@�Rs`ڝ��� ֛b,6�{�u$)ѽS�b�<�$�y�\ �jMʩ6=��e3���4�]'����ф3����r���E0��������BNV~�z�!i��z�v��0�p3�O ��M��.��#n����pS¾����5��v2t�9#(f;\{Kv�$5V��Z��^_e�*�����Vb�'p#fR�-@�QҌ�L����u�O���}����4����F���h��˸��{o��**���έR��8��OL�pE����e=��S��י55�S!m��\<�T�#{�E���PQ=;�p�����L�v�y4u�E땤�gtq �S��R�R���+R�{�*������]y1_A6/l4;�X�����6n��;Rir������)mm 	�;��ȓ�l�����G����Ю4����
�S�!b���n�yAiB��a���V�7����﯃�$Zh�b�o끭u:*gWlP��� �n��%j�;��v�ѻxA�K1{�i��]���t��S
}�fp;�,p���U�8R�Sٲ��N���2��|`5����Tx0S99h�D�y�Viᮡ�8_ ��$�Y�6�u��Ƈva["��MZ��[̬Ar��S�ֻ^�:�[M̱�z�Ͳ��7�3�lK�]�l�DCH�8����]��(;-�݀!�}&��7Sԅ��m��J������s�vF�r�n��!E�V~RvoXw;R�ֲY�s�	7�n��Y���V�K�v�0��T�6|v��P�&�Y�E��[���48��T�PSd�[t�*�Z킋���A�N��2]f��>�77z�j�S�%��������kbA��Z��PT����"; 4�.�g.\����9]%w^��n�)�N�������~�F�術L�f����k�qV����a����TOj�+/�����'Jw*�o��5�	Y���1iHSe焓����L1�M4�?����DEEc�s�:�:����9/��18�T0ȶ灆%`ZV5�E/�*�9�����<��3E�U�MM
��Y���PƝM�Jl��S3/4�������[
�Fs��N��q]HT��u�n���_]��<�H����
]�*�/B��	�+nk}_RnY�-�����U�h�ʉ�T�n��xJ(ʛ�{32�U+5�4Js��o���Ҹe�)��!��W.dg.Q��{�c�S�f��o�6C(SAk���Q6�ī��]���͆�u��v>����d��3^�8ӻ�$ȭ�0NkeR�J���/�7���	mD�9���`�x��s�wX�4#V���A�4i���g�;X���[�@��ym��|��eZ�+��(l(�n�-|�u����3eA��W�c��z)�m�����B�H��&('B<Q�v�+̚�ެ��jh�i8�gIѓ�A*>7��AiZ˥{����w��o9d�����/��;'17y��V;��Ԑ-A��	�!}�u�f�m"���'F���-��S���qn`Vk�U"�⢃��)��Ų��;�Q�6:���[�l���ǝ!�Cۖ�ݹ�C��������Lq�d��$�u��u^R��bM�X�"�[]��V	K�����;;�[J�ٴd̨reY��^
M75�J[ڮ�N��r�*V�av{��2ARK�C7�詘,��du����N�R㖄Nf�n�1�M�w/�4�����y��y���?�W
.���*f�QOλR�:%ғc���2I�&����~o��~#S̋��YdFT\��\�T�%��"�ܩ�D�
X�9�7����o���t#���t�ʋ-h�D��e!�p�#�;����_ z8I�q�6<j'%��2(N'J���N#+�;uI!��7wT\�;.�W�NNBTFm��	\���R�KJ
�Ow���C��MV��.�ˤ^gl�դ�O2ef�)�AI���:���n�9�P���
r��$�{�y�Fr��Ȱ���$��N]���B�IȠ�̑��͕^���Y�#�����+K��p�J�O�9fAF�9^h����t���F9��z����T�P�8K�7�
)D�:9b2�a�g4.�Y��۞BK�D�=�:Y��8��<w%\ʗ$��(.����AE[��D���V�3������Nu�|E�,��cʙ���H���4�[|��Fn(�^+uڶK�A���j��[6�}�D�����'l���VL�NN/�Iۍ9��F	�#c�k���;Id�^�)G&=��MxnJ=������~����۞kv4�G<	������~�3�7��7��+���>�r=�Gmk�I�<kV��M���d�'n3�8�_hm�O��=]-�}͂M��	7V�i�^��6��}�08���s�������ʕ�=��TU��]vy]5�o���3S՞��>�Rz�0ד<����=^����3�w6_[�w�_�
�������a/3D�Ȯ���=�w�K����a����t@�hִBk۸������K�uǧI�9���v�����f����(���Ҟ��m5�d���?�ϳ�Ḳ8v:Isg��w�t�'@5'5�(�@�yW�qN�=��>�� ��j�FeM]�����������{���~F�Sq�O�&���5mpD� !D@�f�ʓ����b����m�6�%JǤ�2K���7S��_ma2L#�{>�A�0Q�ڄ��f�tr�h-�����;�y�e��I9يj�mf�	cY�^����5vh%�S���0ڭ��4��jT0&;Y�F���_Υ�U�at�k����^��;ۈ��N�q������ގ�{A� �g �|�ߟ;ɞ�;���Z�r��ﺺu;��M��ĉ �Di֏v
�0�*:�C]@k����:���='�@�ϲz��ٗ�;�ȉ}�8�{��
�3�P�F+A����=��k��N[R��	Q�f6r⎒/Ga|n�|OcO�,��{�j���c�$�I�3�z�ӵ=��tta<#" � �$6d�l;�>��9�g�6����7��x��B5�b�{����z�̪�ݚ}^93�Hz�����=�ۉy���=<_�w3~�2�g��rvۃ4?Vhz5rǆ���y$�w��	�vx�3���|�@9�k*�2k�5g��^�v�pi�kX����l�o�O�����������r�B�?]���k�۴4�K���'\����
o��n���top*C�)&� ���ꁷ|6�Ǖ�5Qew��t���9�Z ���.P{��N����ݜu�XgA���Jn7O�A���G^�CVu;A}��7Q��ŀ3P�`�3#��S�s]O�n���M��N�<������I�b�=��F������6y�NO=ZX�륹uSř��{�5�|y��;�c�������Ư��yt+U��)�]7u�:�/��&'mV�����*Y����r/��o���8���К�_-�X���1^�.���|ڛ�{a��%�=�K�b��=oϷ�[Y1����f����N��^�D���{`��!y[P�ܡ�X������>���d5�[�6�1b�S�S���N��<�f��1�u�a��T��'o�LsJ��>л*w}>�e�^y$�/k��|�.^�<�'��(�9�C<���l��������ў�Q�2��7~��(~Ԣ�	��G{�F�����N�t����y�Evx�G'�c3lΖ���d���)�b����K�^��^c�K=��復R��#}�\;�s;�֫��؉��գ-2>��+t&�zY��!8汽q�p4�=�f�@��� ����pM�ʲ>�u��)K�gm��*m���R����d�P���s��]��i=����]쬞_^�B�R<�ֽ�ѓ8^>���J��<bP�馝D�v�C�SndPo`5#�Ft�����=�7s6x�z�q=~�	G4�<4 ��.�f��[8��۝u�+�K/�9���|+]OY^�]V����'���8�5�z����S�<ۗ<K�MM�q���$H�~����灝$��9����4����vx����0��E�cOŹ-��l����o�Z3Y��\�O+6�O�Y�������l�;�l�ʺ��J�τ��S'��Eλ<�z{'��@�p�)l���>�:8ƣ�P�����t)u�U�,��χ�5��}7�krdU.�Nӯ��B�/�꽤����MI��d�0g�fϘ'�0��]r99w�Ϝ�X;�}�׷|LE�i�{���@;Cg�7Gy�X�9n{,�s�n5p�q��H��7����I~g��W��.c1�賽ۙto�x�}���n���٠bV���nv��J���N4um]*ں�	�,��N�q;Ũ|����Jf�Y[��!;�xF�J�Q�]�v�p��ޚs%\G�2��wL51�1!����M�W;�V�r,W^'���i�mS��"����չ,�N�W@}���Q����Z(}J��Z=\�Ǯ*���F�ӤpJU%>/͌�����D��՞w��ʎ`���+o�K,J�����>���&����\s3J�~窚2��5︑N�`�cb��X��Et=�1sm�ǽ<5�i:w�h�9yd���GA.G�iK�{ځ�\i׼��Ɂ���:P�;��ܞ&8��Qz�=�f��vi8���u�V��V\�Y���vmg�� � �>���k�1�5�9ZI�fMAܪ���/�!�l�]=��	[�m�#��Ar�H���;#���s�<I�k�:���cV��f9������p����;�]-���o�6	3��p�d_��Oi0sh�l�̊��2dxϛkd�s�bbwc�p�h7ٮ���u�pqb*؈�����U����q�n��菽^���ʖ���WN��f��gɍء��_UK}P��ji��%)��U�v\������n�W^�Ū�n)p�=(o$�4]&~?%��b�Ld��qV��,Waȱ�%95��\�|/`��b��\�$��,.�p�}5Ǥ�*�Ʊ��3`�'X|�g]�8�e[�/T��Dw-���ۑ��`���ڞ����.����t�yN�'/5`�R��zvs�<6O��\gB��Qk��ړ9��Y�����]�N:�_��l���ib�R>��.��������<���g����h����35*�=�؀��}���wޫ� ���\kS�A�I���=6���{�K�S��N�Om>A�809�`=�Q�3��w���	��fAqC)M��}&dU����_�r��=��Zo�_CPƙǾ�&d��Vf.�P/-D�$H$ӭ� c��P#�	�m1w\��^y��?�&��Ӯ]+>����ԫ��]<~҈�qh�ez�+��W#��~�//ҦemE�;���f�?z��^�{�/z+;橕/���I1:k����4�>�k47���A�'�#8�X����w�Zhy$\A]�Pe�跒ܹ��YW�uY�'����W��!�fc��Q�Ğ�O�U�2nl�w8��`k{iD݄muEN���]����*�����[��oy]N���!�k� �[A�d��7K����qOJ��e_IM��{mw	MI�����'&�c/rj|CM9�
�rň70䍼ᣳӽ���^�`����]��c�:~ˍ5�ɡ�P|��csL�Y~�LGMk<�Jv�|塊�z��$�2{��5�<�A<j���Sݹ�>��³�g��-{�m�0��ϙ�k���>�5~S�2�>��秽L�ۨ����W�Q|M�%�y����Q�r�#)���j/��a����!�8\>�^٥3����e���OE�|����j�Ľ�]��k�zx}2o�����W]k/],^ڙ<ęqA��e�&]>��]�5WO0W�,��	;}S�z�y�ג��$'�:�g�I'��N���=���ۮ����)��R�yMe�=z���ݘ�.�[�fG����jFP���k)���몎���h�T�P�eZ��}��r-����zm�l��g�:���a��X��ղ�/a{�7A����9'[�sܰi[^�)�b�]+����a�l!���Bf�[6��VZ��e���*�C�Vd
���i��ڵ��H_Uې*��Ngr�Քdk9VaT�t��k:;R��Jw4��ej���dTi���b<"�smӿz��9�"�5;}:b��%L��U��<���t�B�4�\w���nX���ٿ���c峩=핝JGF{�Y���C$��U��.9�a}���5Lإ^������W��2����Pǭ��Az�)�ܻ�y|$�$ou��Q�t�=��C��6Fc��,��`z�Y�:I޻�R.d�ճgWy��w��≞N�z��_G��̔����Nw3mע�ܣ"�X�y�{ν�^w�K�&�>��� V��?�1�$ֆ%�l��	-���ݞ�l[{�S��O*��%�Gl�?sy�z����q ��<8�᭷ϝ�Pz{X39��<ǳf�s�f9�Fz����
�}R��2̨j,��Ͻ��E��x�k9�ʠs2oL�) ��}��Ҩ�?[��Z=^X%6i��3rtҘ�� ��/3J0��y$Kd���u�9]�r��z���Kh���L}��r>��Xޫ�ԉA�mV
*qU�Y�v��_Gt9m=(7�M;����4����V��n�hT��ԉ*�M�%VTK���)�_D��,�:�x���0�:uM�펗ۃ� $���s:��f���T��;��!�C+��.�ˮV+�g���n�0�������s�W�ɥS���sp��ʯi��֯��&{-L��_�b�u��
)<�SS}@�͠ݧk�uT�7Pn�M�v�i�������������W�4�y���t��w7�[��Z����H?VYY<l������H,��C�N��$��m��S�*	�'7۲ޠy�gn���?�d���Fv�����:#Ft<�ޑ;��o<^+vf����\rV6�H=�~����~���c�<Es]�_ e��ڇ��zL��TYvP��#���l��@��#b���g8��\Y���ݺ-@�oj���V��Jױ_1W+�ڢ�z{�͞��{��j��=�e�39���1s��pݏX���"|w	��#�����f��Vmљ���/�Bm��7��6��z�	��}}G=�~\��
�,d�=G�����Ty1���.`�o����SOS�K����a^��f���L���E,J�Ӗ��.�jOm�;R�p���ư��ރ^6o7]�����,&0q�g�ʹ�٨��"@�h�.E�$n��; h�zl�*`L����o��WZ��L�y��̇S��ץ�z���u]S��V�:h������,o}Hc���f{��޳{�ƒR�*���2��^^�.�Zj�}�6�Z1������CL�=LkɆj�0�t�]^�WfX��F�}�E�a^�hq�=Qq�Qx���w�w�� ���R:�2���(w�Ei��]c�Qu"g���k�[�z�n>l����Y���}�/Nrk�H.�370��a����p�3g&p��Q�g�q�����n۫�}��!�����R�`Mkʌ�_yӱ^�0R�
]թﶫ��Ҹ2�/ �ms�)˗�&�}��<�t�j�ڇ�s%_Υ����*F���/5�c����#�L�;H�F�M��d߯d��Y�V��ڹ�<�^�tW������>U��J���8_6ջ�x�m]�(�7��ڷ��NTp�ws��72�b�!�nc�>�®�#+�֪�V@c�!1ő�Wx�=�ٜ�t
�ћ�U�Y���ч���-p2�=�
�-x��QA_IJA`�����w{H;G��1��ε���n�\8.�3�gmZ�D�2�z�|3�_;w��b��E4-�n�Wwk��N�������b%c��Ě{�m��C%��SᇔW�$��J�ûbȀ)�gW�^%�����<���q�&2��Y{|]ɋgY($�1
;�@1��q�9]�xNn�'�މ�e7˲�U����NI����5%E��|��9�����]�v�Z�}�㴊����v��E��)i�2�N�7�q�('�	�钋��v��urs��֦yu5q�6�<��?�y��cc�:����5�#6�Aҵ'!��T�4K|дt���Ǜ���r0��c�)�j��Ò9F�tqN|(�޵�[\�
�(�1�Ԭ�#h#�x��#���m%l;8��_h,�dv��������T
�23�#jy	��][)ù�2M5.���*0M��l��f���9[q��a�H!��Z�n�Z��gJ���d��Y�%!��ݼ���z&���PJ��	�&��E�l��M��5�Zd�s���ce��+���o:F�b"
�@�z|�^�!�1�XFp��z�>�x��J�sO3ryds�`�&u�P��rb��X=�N�����&:�t%��}Ջ�W�����s4�n�5�A]���;y{��Կ�3���}Y��Α������v#w+�Vn�ɼ�v�\c]�kM��UN�uː=Zs%��$�R���`�AL�6���nv�)�1}�H��	�]��"�u�8��g�e��0"���ja�y)��[E��vWB�,o������ػ[��pE���i����V*IY�;i�Ȯ�2�#�r����D۰��w��4��� 5���b4֔ٹW���6��d�a��Z�uì��
.өK4�iulIQ��rn�5�v�LP�eΎ������כ��m���"�1��!ȵ�Z��v�(���U��j��U��/+�|7lT�`ˉti��ׄ��L�%��6v�!���v�I�K�R�I*�ف�8K*�3-Mw�**�oO9����q�{rh<�n[���u�����a�����$�	J���of���-��}���l�Ѣ�μ*�����.�m.��1�
)A��p�g(E���vh.n��
�˂-y�E� w,
�64�Z�gP)�V:�Wg^P;��=Ҵ$��І�p�4�8�����eGK�j����T��3�L��ͫt����`jxi�Try��CV�^vk\���j���	�V�)2���]��-Ϋ��M������ߴ��p82�,�qZwr��H�>�0��T���~~���ϧ���犯��I�;�HvL��N~]w.�Z\����uΤ��E��I�$�\�]+^>W�U�����o�����(N(E�Ts���N����4�@QBEH�E�Cל��<rE�v�ߛ���c��J.%�-_(x�.��!��NT�TB��A�#�y��+���$�M�O#R�I$�M#�U���$�d$'
�W"�E*	RBAL�2��P,�#'qM���S��Z�FI"�(�#*��ЪB5�q9p�f�\�ӭ�mʮ���9+*:H�9�]"]r��pեB�k/�x�<��N�E��9Ni)��)�4�Z�H���hD�ÑJ��"��rV]%��G,��a�x�'�����M��q$�	<�s�ӈWtw"*$(2
x�<�*<+6Bs^\���%B�����@�%*y]4�"��#����W�����p���`f���Ke2�E��9ՙG� ��s�|�R��ܒ�n+�&���(��#]�4�V�̹���W���~�<	��6�|2���h9�f�0R�] ��]NŴS��"���D��V^'���l���f�B��H\sL=�OS��|:/�sH�i�{ ��qYA
FL8y�i�sc?B�/2�"R'׽U��V��kH(L&)Պ�����͵ y*f�;(2��q�g�Uz��h�k�1򞄉&�?|�W���o��t@�`q�ǜ�τnϨ�UZ�����҅&��vJ&6KMW������mn��AoM'�mt��V�oV�^���P2}�%��h	�c+6+kO]�|]������[/�8�1,�ߊSL�M]p��q��6Ju�X�'�S���Tn5�)�h�W�!	�r=`��{O��Jt��op�FSm~�<��ȸu��ztu�d����GV�q�����r�f87/�`��q#z�$��I���"���a���/j�=�ǩ�N
[s[���;��|���G6���n��8�^Ω��ft={�Z~X�A.���4�슫�؇vá��&�<d?K�����q;1,��n%�}ګ���/��M���c���P�f��k�s$ ����-a9�;�3r�OA��ݓ��~ۉ>�P��<X�����xGN�-�$�nF}�s���w��u�>^}�`��ڋ�-C�ۦv#�,�����}��t�2x'T9�U�+s�l)�Z���ܹ��r=�_$�K�w����u� K������K�G�1��6K�y쟍�ίƤS]����UD�T�K7/Dh���|��ֳ���i�3��lia��8>�����v�-J�S����xš�^��9��A�k,{z}[c�LW5�y�Pb�݃P�݄5\�@Z����B-��M����hgՆ�pǒ�e4��
�-A?tŨ;�X��K*~ʪ�Y��*��"#��c�jF�	X���TpК�4]���f- ��pφ#M��f�*�tk���<���"]� �����������}���5����ϋ�]�>A����̻��k�C{����&�
�Ƶ�%eySu_�`�FՄ^�Uϫ�۱@cWR�ڶ�QӺf9�D�c�&J���Q�g͊e�����x�`��F�n��Y.@�n��^�U%ռ&��������0B}ka��C ��g��|l��s������^c���R�ܯF+r�A}1[�2a^1�����U
P����qa�r�m'��!��m���3����go�Ґ�����:tM�^�_T��=�n.���n,�!�D�B��[fz�cҒ�E�H"�!$��y:��U'$}�r��)�5p�� y��]�����Ҕ�����i�ǻ7h���RG9wK���tĬ���-�ݽ�^�3� ���Y���S��;p��%�P��=�)�E)��)��^�зi��f_pճ]N�4r����p��C��oK��b=��&X�LV^Y�N�i��v5�Za��n��U�~{/�=z1�N��fƘr�L��ʀ8������wc��׍���vB<�ݛnN�8��\�6��s�w���8{d-{�!����9�+L�_lVVi.���u{U&V�g�%��$�G),Qن����܇ǐ��̛��-�Q���K�_w�-�n):�7B͇2q��⨰��<ƬR�`����7��۔_N��bKڧ�`��r�"��Y1@0zb����Tn�hZ���е��%�J�\.��*ujE����kckt����r}ŇfR:9�@|.hmK2��u��)P6˦��;�X���ε���H3�3\&le�����dȗx�`<�C�m�d�0	:#z]�F��#�ٸ��H��<��wy�㨙vX�����lhtg/>חx��C�|aQ�8��r��E����/�*�P|(|�t9��٘z������IL�2;s����S=BC�*� �Ȫ�� X�a��j�2t�#\d��e^��T��F����ȲB�nwg�
ԟv��q3Q��Gi�gk��o�G��#�����WC�{y�!��  �=0��-��6�ƶ3��2�Yqn �f�������[�L�B�-=��N$���Z-@��K$ ��6�m:`:��tS?I�U�zR�[�;��hV�������Uձ�U��2=���fP�eQ���&�a��|V�dc�e\9@�3�r�c0����s��Ezv��WB�,2%�D��W���Dc	g���1t���R��;�C�ᩭ������H|�`%Lݔ<CO��W�Є�0;BU�Ya�l��[�{{����MP��v#'1�}Ǆ�o��$8X�!��� ��;M�l�#�ū�zC4���l1y,�\�ĲoX�ƒ4�S�_8���OZ�� �6O��ǉo�j�o6��~{���Oӂ���~%}}�0�ʥX9�Kz���:��p����a;��Z�жa�Z��QZ8�QB5���	�ۑ'|҇VUt=����T5��a��8�����3]��T�S������֡G1�uMk�1ln�.��0���殕�~��?�uz{�ĭ��������3�0�/`�.�x�ױ{tա���Dg���pt�6�N��*��c��X�Nћ$�X��=E9C6��I;����իm[���+m�.�e���FZ�B�HV�b�2�in�.-�Ggr�r��K�xF�<woF��}�F���EK��n5� �����g�����j��E���8Î��h�[M�K+�.�qF\�͜��玲���
=ʅ��G��,���-�׽6�X�2��n-yUInnC�]�X�s/�>�zfy��Ǻ阗���Lg�h�^D<끅�Fvܴ�71���X��nMhvHvS}$�Xc�C�"ex��`��y�ސr�o_G'|��n�?>B�͈�8pO�MIO`��+�s9���q��ג�]N��4c�}Q�3�?\K�=E�[��m[:��Z@�a4��rz��ǳ�ޡ�;��4�-��d@��� ��p�Һ�e�:)s<�ֶ���<�
��O6Pa`��_��W���,�����}�ݵ.J��� �i���&�^����/�9m�\���[qDh~��@����(��P�%�2�1|����W�ץ|�X�DC"%�4�̝~נ�j=$2j��4��UӬ(�^=���|��q��X,�	y	��4c+�˾��)��kzN�ٓ(`@)4X���rxeμR�ebQ��b#PW�X�� ׅ'MxG�O��<���kxԝˊ�|(V٠Nn��&�b5���1Q�?����(:�����f�Dx�.%Y�m~�K`w8]?��}�3*g��H�(%��i�W5�9��ՙ����wX�����ԝ�;9_N�y�us
����z�=R9Wɛ3�گ�C���/{����پ�8�;4�K�0M��ƀD��Qz)�|"S��SH�kk�<���Uq�%������ozw���"��umOU���P�zT���Rr�\�$�[\Ù�;�ô%��'Uef�\�t:TK�Q��=��8@�yȄ�^ڞ���Ƣ�TCp�	���~P��&-NDE���F̗����E:��sx���zC���`d0Q�>�"
,��C�n:��l���9!���3���4���/�]�־�?d���*?a��ь�#������D8��uP�t��2F�Z9k��7��AnB9U�߻����6�t�ʢ��Ż�l�0g!�����(�+S/���һ[�K�:��N��P�~�7�Pc��ǧհ^y�e��wm�����2�rr�{yy]�۽��4.m�$&�3�mO�چO�3��i'���0W�SH;@���&�p��M�����,α��p����^��#��0�@���ojF�V7�?<��Bk��v�e����|8��.2S�kO�3D^={^m�lw�q.9��0���`�}�uT���V6c��	���ّ��]ʺdy���gAnW�O�JSӂ�:����d����]�0D�y��U�ߩm�w�
RU�����<L��B�_���|)���nL�Г�&�c&H��;�*��JK݌��\m<�]], �� \AS�����Ce��Ď�Bv�wH�:h%A~���� �yDӲ�8�5Fa��֤���6�hl�w�\E!��������u���U�D�"g/2[��A�RY$5x�8�^͛eCu��hO-.�U�'$���&�i��k,h�:��WPF5�7���vOV�K�]X�@�[�PQp��3��CD�5A^hΙ���Is�B^'���d�2a�tc�(��)��,)��[9!����<v�Nv�=3��W�1�$G7�(2�u/	;nC�7�S��	�{1�YJ��ʞ�����[������ӌB�	�d[A��o@�i�H8��!��.�7a�liRewg����;����fum�C���I���n:p�6S��F3��݃�A�OH�Yӌ҃�gtQ͕�si�PݓW�Ͳ.���i��m vk��~����8{h:�6��r��
T�h4�.�]nV�h�K��VP�gh��̮xj9r��PX�v���������cv;J;��v)�`�9�.�[uԘ�����,ߜ��|]QaY��j�V�Mr[��=Q=ѷ��j�f?��]nI[M������qƵ�݉S4?J�6ԭ��KVs�Ή3��,�F=;��y��1)"7�ܠT��#c�]�^��Trnһ�KzQ�~���6��l��\����������降�����g'e{����%W�d�:C���`�O�(�T:�smg1�i<,q���{*	{k����t��a�49��5�$*d^ÿO�G���g���3,���X�J��mܭ�p����ּƷ�:��N T�����rL�w���x�	�!�6߬eK2N��z]�lcS�YT��b;���쮂��ʘ z$�Q2����fA�ƺ���ywo `E�ݡTcU�1�|�#�vz��iKc{7a�U���:@A�za���Y�6�ƽ���	(��m���w���p'�/G\�{��Ƕ�u��6-^9��HB�&��q�髦.dӋ�t����
���\��L�L#�q1w4^�TcW\�K[Q�!kߎ��fP�`�<��ohI��h����צya�[x(y�φE3�͍����lQ����K�Є���{���[ŋ�qN��>K�k�,��(]�{j��b��z�o4���A�i	Đ�e4���v�a�sd[���i.t�O����G^��Hk��J`��B�2s������C�p�w�6ڠ��5c)��ݲʞ�/g�x�%)]L��{�q��iN����z�`H@A�K���<��^/pM����P
X�Fe�5~c"'3gS�����h�=[�j�A΅�4#�B�1�49�u���"˩يu��)Rfh7�������~���Qfr.z���a5�fJtY�t����F��8�_X_��������TPz?�e�2��fۥ�8��B�� �kH�M�4��_E'L/�J.�s�1�����g��A�7;EgFӳ����������vmd �L�:�&5�B���*���,�'�T4�0��"޵��՗�4��?�B�:���a0�����nىN�S�V�.��Q�X��iK�:3A��lu���7��u���{p���~`o�:=k�z���U��E���U�X|\\+��O�O��N�#���K�R��<�w,�C��?N�`�8t�Dqy�;k��v����es�v�Y]G�(�g8�;��@咩1	��fk��3�׬3<Ǫ����ĸf�p0�E����^=:�n9O6�*:���7�K������H��Kώ�-�b���wI����Y���Z����i�й�8�D��}��tOg6����0��������E�[���螊�ƓCv����쫇��g��,�9l��=OE����ӛ������Ee7Rir��L�h�(�	�[�_�
�X���=b�+�EIj��k��Y�x&]ܢ�� N��I���s�._S��M�c]������Jրt,�����5�67�Pk��˰l��v���S\D��6p�;H,<�1��������6_n��f:���E<5�yg�����5z���Nfc�ϛ�6Թ*f�Hd�H!��0-�VR!�g&�r|}�6��ǫxT:E;ǆ�a�w̏OUZ�(�(UM&���8���� �	��0�&>���ڮ�a^=�Bޭ�o��B
H��d�!�y�[/ȴ��6�A�f�C �f�3��!�%�{)M2����l����9�=5��5�s'��Uө�$ֆBQ:��R�XI�i�2;d��DJp	˼'GˤS�����e	眫�T���u�T���y�C5��FY����#����'z�$��I���"��v�El�&���:72�7��{x��ɳ��#Ͼ{aH�7��M�6��u{�q���S6a7C�˭�&f�-��B��Ž��y⢗��İ�����1��
9���혖\�:�@��=���LH��?WDO哿V�!���x{J�P��0�_��[��b]�:1��������I�c�<Ke�]�FK��)�A5mw��I��i�oV)H�S,ٯN�������/���<0cW���~��߿}�����_ �~"�K���k:١R�5�&�)v*�e�4���Wb��N�"w=��t��}�YOL3[��-VxhW2�^����6I��cCj�S��K̍������+�ޥ�L�w��^��5=�_e�z��m�۪��rP�(B�i-�[�� ����`a��(p�g�G#�w�6V�K�{e�,j49���Y�iVv�PK�Z�P%��i������b���9Ea� n�H�������F�F�� �NeۋZ�aЬY�s]'���Zwm,�;R7̱E���"er�]6>]�]���L�s^�Vf\���+��ܺ���S7 [\���]69-�v¨��djؔ8���\��
	�*\��+��J���v��$�b�=3f]��Ҳ���qI*�j��swQ}����d�s��1s�[C�@����Ws���L�oS7�r�"���F�H���#�K����Y�}Ȧe�c��3�̿���ݹ�D�b��tƕ��4�H�]:1L!�ԃq �:�ā��>����ɴ�ʊ�HM)���.�O.�P��R,=a�v�(\�u�)�Y�v��=QS�}�� �*��7	rl���ZsQ�D�r����Nứk�Z�I)�w|3O[M��,�wNwaQk�㖅��zr�	�����xQ�ʖ.m�Uƣ�áF�>���xb�+x��}]���Y3wB�"�.�6�Z�t�aӈ�E�*�Dݧ&����9k.J�Ӵ����m��?}˳���zM]k�36�"�Z����x\%�^�.pf<�Z{g�V�jZ�f*��ťtU�C��<$S5Ue(e�n�e1eew^ΐ쩗[�hGBΓ5>1X�F�g�v]�0�T롶v���C�#M "|�p�3���&�j,��j<٦����of���CyH`�xZ��펉F�N����:c��x��^-��k&ʮ�Yp�+�3(�����j�\8�A��y��j uuJ�0���Uqn����9;�N�:�D����2��3�g��3D������vk W.��ź���[q���໴D�[9��:��6���PBw+鑱�ou�Ub����8n�/�0�σ�z��'�k/�{s��=5��zݛĚV+j��0-�����G4����ȓa�;i��t������/fm=��hf�(r�{e�N8�'bho�[��1ﳈ��3}�4�2,Z�U+qr-Dՠ;:u�A4���k.Ա$w�9-���B��`�-�{���6��s�:��vA@�P���z<�d| D�Л׮ˎM#2,��������à^)dڝ��w+Wm"[����yZ���-b_s۫��]ؗ����Ν��B��]��Pnc�=���*⮮u��]\�;�6�¦��.����F�LJwN�wJRo5�I
R[8R������~{��(���7�w=7�7�Ҋ9���~<x2U�C�r�!V�Njr
QT�AN��LY��u�{�o���>=�%[K0�*##Yq$��~]͑�i��\SJ�Q	:
��(\�As[�|��B�o���|����0%J�4iG��5
��e��Q����M���ѥ�/�/D�I*MSZ�=��T:�)���I%E�$�Y���������ӫ���*��LS�P��J�!P(�U&TF�S$���V�B�36P\�DT�FE�At�$��O��s��I��{oEʫ���2.GV�Aghv�P,�%��R���N��Щ��x��T9<T{YDE���y�ǝyXQp�XY���px/d�\3�4��C�|N�$UQw6�T�s���(�AEG޻.�$���4��y�/XrN!Fl�(��<�	PEw��Ȫ�]��Q����P�T M�Z���am	8�.j�2R�+x����@M����m;�U9���.0Nee�U�մ���6�U%e�����=�X4���U�O[��0r$h'�v��}�b��v��(�ë�cYk��Vߤ�sP/��!ݻZ�������_^�����A� ���C��9�mC'��4#�a���#4��p*(��� ��M�QB��ξ���|d�ø�vy,퀹k0���H�J��?<��Bk��vML@�������v�id�:I�sͼ*"]� �4\sH0���6۝����&�:��R�rCv�&iD�'jJq�j���o�i���Oȧ|�PF0��ȼ������6T�)jOsגy���{5�X��A��A�rY$1F-�sf�c�gO����j��:*mU��ٵ{]�����\�c��[C�k�6oB	��� ��j��WV3ю�Ơ2���pͬb�VDە4�W�{z.p�e�:O�D㌩x��^]:ɲ΋�D ��E'Vϓ
V%QaLָ�w��j��Q{g����tك��h����h�r���T�����GW\&�=�'�D�S6���܂�.f6�ޯ;�t m	�)žŰ���k��|k�`�q6eC2]�i�3�8�뱙�`�{19��"&��6{e����FL�_5�Lm2!��3�VJ1�½�ڣL�7����U�Ư},��٢��x���7v,���fú�f�AʑN�#��Vڴ%5��,����.rn+�������^��K�E��e+�1�[j�^{w�7� ��*���d�t;#O5�8�'Z����Ӿ[�	����F4Ð���A�q��:zEV�iix�!�&��Y�)�S"����8��m vk������<��]L�8���1Q=�yJs�*��)�F�D��0�0���"�RXבچ�ٷ�ꄻ��Q���������b2/Bz+�X5t,���+��`oc[�L���A���Qx�f��J�����ӇR�8����"�ƇT�m�v���D�q���{*	{dj��K��t�u�54[�{�W�:y�Tk��Ħ�^ú����>f���4�|Nk�R̶����)P.�j"����L�m�k�=��7o*�Hô�R��@��^�90!޼8!0���~�eK2N�N�z��w,c�Jl7�#�;jX�0��]��f�z�3 �cC�[9y����Έ��2�慕--}��VX�%�G-��EܦGz]��zA�2	E@A�QpjZ4=2Ή���j��Wz�Z�Q79]�Hb�|�fXfRO��3^�5�A��*,q�.��!y^i��t� ��յ��7p̕&�I������L/��*�+���Tm
�Y,��҄:	�,\O�����n����ic����4SF��<6C����s6�-)�n+�L�rSi˦���]sAr���Q����'P��Z���-��I�
�Wdl������`���8hE>��{�?�xk��8{���U��'*Zڼ�HZ�ve����x��ߨ�v�9)%͛�'�d�t���똨}�lS<	����g��ڣ"'jX���M~��3�ZnC�?e�f�Ձ�]_.�u'�y��,�@��i�q<(�F���0b��R�i�Qo���]���}k�T�t�)����S���o�k�<'�o��$8X��|���ι|aVl�koR��'P�n��@S�kӽ2���Y'X�Ƽ����z�tdW��:ָu�w�Oһ��u��5��a��:��C�i�Y�� _E'L,r�E�s�1�1u;q~�-�̷Nm�:e^�#���1t>�

���9��T���ȓ�;JUYU��^��w����v{g6T�R#s�w)��C�K��a�#��`���p����SEՃS�P�v��F�tT�hxQwjj��ݤ��/V�E�8�}��ǻ`8�J���������Y.{�z4C�"b��6�w+���1k�XN뢠��7���?�\`l�b�?�Р~��E}�]�"��(bb4�b�SM��-�z�$]�<���N���>}�8�"����I���fŢ�&��uQ�H�湚��9��tϟr��r��uzǽ��=�X����get���]N#rG�y�� ���X�e�3�����ؚ5�������ysShX4��2h�q}w������y�R�Pܙ����f�\I��������6=q��z�ы�dX2�����Pց�L]�gxpO��<��{P���l�m�_J/�Ǥ��H���%��[&�lC��ʈa�Z�1)ɼZ�3���50V�"T�{Q��gdf�0R��IO.�in?9��Z*�����s*��[���y���,����c��{d����ǳ�#[�nf��d�-+[�t�j˩�l�t7���ɇ>���Cai@�J�~���ʫ��})��硹3lϽS1`c	��[�وE���3j&He�\N0-�.����zǫxTM2r�@��*�b��r�R=}��ż{b�#/r�K]ʦ�TW���,r�5ZSI�*����馞��x(,6G2m.t噍�&η�"a����ׅ��8VJ���'9D�/`�4��Mn�om�����W����[�ݏs�����D�f���u��B��I�<�>x�Jt���$i5���i�!�U]YVH�ٮ�R��\:������*Y����*e�#���oR��E'*ܘ�f���u���7Q�ߦV�3x_�½�P�u�x��[��c=Y\�Ϟ�{/٢��@'~��]�����/���N,\Vlޤ*
��FeY�{%�Y�Y��&����ьm��%�V��x�M�5�#�10C\ySs�o@�J�!�]:p�'Ob��9�G�B���o?����xz�:�WrP��gQ`Z�F�X��>�� �z�M����C�q����a�fn8)��g�6c*��T�b-��ۑ|�`O ����r���?HN��X*aQ�"�q k�.utS:�Ƌ�U�[��Z�թW5��*<bid�e/EGs��q��wh��v�,��W�+��6�r����ɥ���IՉ2)��4՛ғ�Z�&ެ
S�
�Y�^�ٷ=���)�!֞�=�;w�Щ�<���zP��C�еaD��,}���ۓ�^���PW��UN�r R������}xBd�͉�j�hg��4���`�h�ݴtA��۞ּh��� �΅���E��5q|�����0(-10���d����zS��n��������"�����^����.�q�q�10��Ӎ��,J"�u]�3kC�i�k�3�|���i��<�EN2H���}kO��sdS�{�2�c
���ѧ"���a�k?ݭΩ�����e�ƿ_��A�c:[�Y$1F-��)��l��Þ����֬���K�2�{��e���*w(U��:iΠ��Pe�R��̖�n��ĹPCx��l����\-����>^�N����3{T��˪��mh7��H�y��^�옱'�nm"D��5����#�ͻ��&���3���+�W��3x�ժ8r�Q������f7^��V�J5�� �Z�vOB�	c@Ռ�c��$�e�Xڰm�n���Wy�5�qHX�N2�/��N�jɄ^�!Z��QI��"SP����F:�9;{������|�Op��Бހf��nK�	�ŨtBd���_`�KY�{w.�6�{��\hZ�TS����;"�{�� �ƟC�H��vC��U�Vk��M&;��\����C#����x	���"��\hӅٲ�_�dAƟC�����i蘮��X�$.�8�I!�P�n��K*�5}0��������xeK_��?,,@%���[���ٜX�ϢWp�W#B�����F����F��L*��\��r�'�JK�;P�Bxwf�)Q�E��-�W�$T�.�?5Ϙ9m�D�_f�Հj�Y��N��U:9�U�0j�-U���NnS�eX����.{p�1� ��C��p�1�:�sm�^�D�q�ǥs������=j��k�q��w8��'��^ù.P�f!��0�R̷:Kc4���aϏw�x�̋"��^v	����x�FW�z�P��1T�ͅ���^$��4!�N��ui�oUm�������8��BhB�����0s�۷knWq�x/ZSf�lj��mdH�VR7(�}�)*�N���7���9(������1���͕7~y��a�<�o,�	ۯ��r�Ǳ��!����=ʯ�x���L�]^TV�L <F���=���Q�v��w�[͵=Mɚ-�v˲�9F�7��^&Y���i:"��@�r�.��U��⺘����'�y�S�ރ���Bn+��括�7� M��~� ��� ���e�2"�P�xcHSЉk�iͨ�'LT���A�q��:^�꨼{k�s�6a ��r/@%�Dϛ��KMUl㰫h��/;s��V���b�� b��:aV�w_TcWFL56.R����WS�4�E�W&�����bh4y����	1P�)�<���Ý�`Iv��u�_�jX��6mpUq�ȩ�h���ۯB��vAeAb�I�J�63s����}h8p���~4�Gu��YF�uSMb�[�����#%�L�"�,On���L:*E=�����{^}��(8�|6u�,�@�Y+���s�.��`��c@"Gb�N��N��K$�s��F���`@�.-�&�"�v�cæ�f�Tm�ƽ\��T3[�`����h�Y��"�):a|�Qu��ǽ��ۖ�є���syrU��n]�v�a]9�vVev�۲�Jn�V֜9�$�c�0���+�{A�蔺�kWO�Q<ɪm9m Sn���<�9H��fn��:��t�f����;%`��|��`q��[�cE]���������-c��˸j�͝���}�o7����z��j�(���q噃S�io��f�~[�`&=�"x��(qT*�{/I����NlKo'mv���n�C�_8R�ym�!ã�����<c��ZDp�nى.�����'hXќ���Iy�N�1�KM�@w�9T�c��]*�^Y��S����#�����������jF3�H��n�b;;+��y�,[�ʭaǡk�PKܽ�J9�]K6��b�:�B���TUW�w��;���FE�z�ukq=<���fI�^��.T�$2���c�o�fy��f%�3��c��j�;�M��s�se�d���"��B|O��xf�vپ�_��zHz�D��'7�:~�/�f=��ѰY���w���TK�X~aA�8��6w������Ǎ��
^��q)��B�V�����6d����:��x�:���թDJ���"KHC ���O���ǳ��9�p�4��"ޟ:�Z�՛�\/-�e+�_���]�2��(:��Ut�0�W��:�f-����]�*~����#��-e��6�;(2�,�e�MjN�z�i�cռ.�.�Sg�:/ke9u�|��r��-wP���B��f�,.��\L��rR�T�ٺ$��,�ûv��qq�H
�C��9�H�u�s�ص�@��J駧+3l-f!��[Q������*�-�c2�eL�gG����3[�q���"��SR�wL�iO�J�����_�����������d���B6pO)J:٘4�M����v+Ӽ���P�&6��{�aG���ޭྲྀ;�4��4 NX[2�C!)��/ ����TZ�D �rxd_�)M2�J4�����=��/f�H�wT�x}jw^��2LO;6T�&
�A�K��N��1�X]"��EE?����Ve'��ӷ��0����h�W/�ӯ00E���T�Ǝ˰G!C��R��HZ�����o1β3{cݯ�)Q���z0����l!#����~��C=:�]���:��4˻�;NZ�8��-?,O ���n]�+ǦG@a��`��a���y-��QeD�ti�έ�ަ�X�l�R�(�,�����Gs�|w>L���)}��WK�b��Xt������Fm�V�K�!ڟ������,tA5mv7�W�s`
��z��S,�Cb�ٶS�kh)����E@�	�$�@��ò~OC��h�B�xL;��Z�8����&+�ݶ�8��X�`���k��<hC����,��ŧ���_e�>��4#�$��bX!kkeu.��)6C�v	�ĭ���S�l��KZ�&9��q�m[\��ڢ�]+��>��(!x�T+b�W�iz�nr̶Czt밖��(��^WW9�+'
K�U�Wr��Q�����uf���j_<5`问Z�Sʜ��76�0�iF�=�4'W�3��x{����xx��;濡�d'?�Z�_��j�p,;������0(->���lmH�KzC�܎�'s+o+\�v��=�<츷���/������6�kdK��h��xt�h�.��e�������m8��=>��,Ӧ�
�d��4Y����J�P��eySѭmuZ�۔����s:GX'ئ�y��J�y�ж(� Ũ�Hb�[>��6ʆ@�t�w�PQN�/�e^-�:��`t���1���h��	F�����Ђ|k;'�P%�Ռ���;��V�	������vX�b9�� }\���~5��O���u�W�L"��,}�Rul֭��X�w1v�:~�%���R_���߼�W�s����
�]/	;nC��������&*S;*{y���d;7S�lD��kR����}�Ы�� �Ƒ�q F��o��w3�0�*)��a����[��ۃY1��Q��ax	���"�ג�@�E�����F��A�6^_q�r��ξ���tC�L��X�8�E�JO<b�K��i��#h��=;�:�q�x��Pc�?�חY�_f�N���]�_dn����`�y�'��vp�"�	ɪ���c����J
X�Q5#A��^��t�LۥW,sr��Yz�!���Ɩ(��oss��S�R]��.5�2�M�bm4w��w*7��+�;��q�����y��+��aR��'�۵qp��".��}3��g>V��їB���^�����ĭo:�e�ft��b}�r�#3�<t]�D���|�T�E�=�qt��+��t8�1^o�C��@��R�$A�bVtM��W�z3.V\w�A;챹b:����ܹV�;�[�j������]�+J�{X�E��oSϦBzoCT���.��n���9���ӑ¸�T�Y]f!�ʝO0=3�ܣ;���6�5/7!tx�^F8�h�L���f��*��i�8QD^⨴J��!,���	IK�80Qf�ܩt�Qu��D�m�X��Y5���p���3w$X�T3fCa����.���)�ftY�'��!�BK{���NJ
���K�F���\�IyD��ev�:��Y��-�Q\�������E�=�U���y��n����X�Crv��캋F�I �7�Q��-�I�+M�Yt�d�%i�V�Ҳ]�z���י����3��s�T�&S��Z`ׯ��܀�p2��o'+%;��n����f�w
�&�[�e�6L��B�:q1���w��2Wa]Nr������\.��lI�Y՜�sy,w�E������o���'.�Ԩݜ�)��&�NWp��u����;�� �8�Nш�����!0�g�l�C�Y���>
���:ط�IIsܶ+Tue]��?�e==�(���⍛u����љ��qk�o���㋎.��u�T��I|�""��fV=�4 �N�v���grA����M����T�rol�WQ$21drjAg0 ��"�Rof�X�i��ʛQ��g/�n����e*CP��u������u%m�S��M�����;�����a�m�<����	��U�8糞ۯW[dT:�6��J�7���U�ޅV��R�κ�b廝�&Y��v�sU���ɓ��wXH�ۖ䛼���k�m��ԗ��Z�ԩ,Y*˼�H�[��˝۹ 4^��9�t7#q� p�Ovc���sx�E3�J��n�h��䷰VM��B1n��$�n�!�*wiX����t�n�p3�js�e�|����-����{������� �̡J�v��D#W%Vn���R��}q)�����Ѳ����vPb�ou���;`��؋�2T�t��*Sht����ü�����b2��l���ri��3.f`oހap�a9#1̓�]�t�Z��%f���Y�o��f��K�m>�?mJ}٭_y�f	;;`��juX�'l�oOv	[L!VN�9e��I.�TPA����U����.p�<��9_#�*�DuW���j��ʨ�Pzl,�|c���7��|�\�������^-�DQ�(��*�2�B3�8��m�����%�\�"��ݾo����²��-��Gnp����y��ٓގF��w���-k�!z����9����	Eť^bi�f����:b�h��R`\���+��׏,u4�<�\�Vf9���9Utu:e�'<v��*B�\��G���"��B"��Ź'z�I)�R��q8Q�ğ��(�E��
L�NW'R)׽�zl(3�Uy�;��e�Rfer ��u<�tI�
a^BF���p��p�B�����ʫ��%Q���\��@���Ԫ+$#�ȇ�U�(���5�;�뜂��z��:e�Y)�8]�Q�e\(��P��"�X�BsB9)`���1�GI����Bg((�Ԉ���Cȅ^ar'$�Aώ�#72���"*55��
��J^Zn��JǜYU�J���/��	u	�(x^^y���������ϒ s��V����I2Q\W��|^	J�^ML�r��J�f�3�4:�]�¯���|˭n93�?  ����oxx{ػ4�񵍚7����C$�:����F��aT,�熣�)=X	IcH�CK_:8��;x�n��%���N�Ѯ���A����@M��OEs�5t,ۙ:�
:y�)a�m@�~t������M@��}`�������
�G6����Q+\v�e�"ل��ī��|�=]�g����8�М���'���w%�
��3����9ͩfMuk����)��o�ѽ���'�V�3����2u*�.�ǾP�9^�R��z�-A��.���x�	�k5=!����,���P�U/w0�K����t��,+�Iv�e���"�UK.l�`[:yח~��j��r��]�|�c��h�0��u%�ۜdw��u�Y5�2	S�B=0�C�)9g����F��ŵ�U[�j��f|e��DfJO`UE��Xͅ�C6-@��K$!��Fp�Q�T�]:�V���|� Ӗ�~�{ ��Xt�O��h��F5td�Sb�!k�fnTsD�C��W85am�+-Լ�P�`�<����e�T9��g�!64��2�{T�%����g0*��)\A��㛕��S�� �j��Ż�gN����܏1Y�%�,�Ы�R��p��[iM�}�V&-�d�����0.b����sT��c��L���O-��W���ȺRf0)v��6M��G1�����?�߾����������83���U�|�ܤ��kZ��'�,q��W�*��_�]I��n����_����^���9�Ll��E�9��3V��y��g��B��xN��J`��B�"��w�0��}w��b��{�)~�y]&�����:���� ������^�oL��<^%�u��Lh$i0nz�%tvp�4-e�-��}j%�~h����ϝPCZD�2����I��Qu��LWK�{4�-�s3�hR����Н�{!S�3������3c?���b�&4w(Q��*��].z���ɲ�f�WW��m��-�[�.��Iĸx`>ϘG���h����������W�6+'M@�w%�2��H.ә�Y�=�Gs��T;��@�z/n;`8�y�[ã��ֿ@��p�[q!���4�����kN\�51JUk=_��^��R�i�m��`����
����6g���z��/͑�u�v�枘f8��ޛd�JbYG?�2џM��m=r�h��ƮG2����&^&so��O�3 �@x�<��yO�����6C�ϯ��c�C�"a/>�^o[�ث��
�1mn��!v�S@jܠ�5��(GI� K�)�C�F�O�����7���]���[��K�Ԍ�;�&A7�n5��Pu��)1K�9����j�d]�N�\��.Uv���u�,Ȟ�u��b�T�����o��󍳝��|���}�������~|
�[�C�OD���円�~��*l��Fk��h9���
^�J<�y[��ti��WЯgz�c�w$/Z4�[A�ǹޡ�FD�ǁZZ@C ��{d�9���W�5������걱Yq�Ki��vw&i^&y��������i�m�k�=�憠���##)˰�Ա�TB�/��ՙ<�Q�ٯf"�q*���;(2Y�������6��=[ :E;ǰ8��lr��6��Uz��kuw7����F��DN�zw����d�ҚN���h���[��D÷k�ݖz��z�U���N�5ơ�%�ʗ��=x_l�(d�-^��O��bX�(�k'L����ƬR9ƓQW���;����������Y��&���P�>O�$����'.�F��	F�6�!W�}�@��gMmq�<�"��?��3[H�����u��C��p�ƃ6��L1��T[�u��'"���uE�;ι:�'��msk=]�����[�G�Ȅ۳�
홡�r����hx�Zu�ԦӦ�}����@%�s@�����?KF0>O�@b\eóTT��2�����w�dQk������af������Q-4p�7^��j�q�Z\�P�Du٘VM
����N�°J��]�wӂW�%�<����]*����j12��J��2�wd�꽁u[���(ӏr�f_�w��{����7�� 9����^����^q�9H�z�%�{�ɦ��:��e��5�#��t�Bkx�#LW�9���l矍�:�%��wf�G:�W:�&E1�&����)?5�2m��O�T�6\>Cb����!��ӻ6!S�p�a��K�7:/���kݦ���w1����z}� Ͱ�3��i�e�65��,~�����_ieu/U���{W�)l΄�5ZP5{����pl��%�%�!mx����M@��q�x#��0(,��綤k%}I��꧚���h>��ĨMr�.��e��/���^��x45�%~�H/��p9�v��B������P�$�Gb�~Brq���oO�)K6֙<�EN2^D�W����'�y��C�S�+w쇆2�s�oT��HbB-���)�
��u�mK! �BZ��!��8�Y�l�Q�WTT�nƶ!������E��,d�S�>�����	\�U�xoB	���	ȵX��4Mom���e�f����T�o���#�7/�.3��%�T�O;W�N�l�E��X��l�7�~��<�Tf �.Ԛ��ꔊ��}����oZ�۝դW\<�]����
�tb�Rθ7|�f�9eٙ;q��ɷ�mcC^r��ֺC�$w�5z�܂�3r%��f�:��˥
J�4�P&�R3/{|��_;:�����?|��������?����y�ϟQ[*�{k��q�JĪ,)��[`ꋇUq��"zf��v܇nADS�u��-5:�gy��L��M�˼'\R�jĪ)�؍�a vE�*����zA�" �vj#�ma��?_F�wV�m��_K�>�3#M*L��8���h]-�Dt�z�o$�IJ��ᚮ+Gl�=}�A}`K#�a���'�f�X��b摴�s꜋auÍC�<�EZ����T�r�8}h��k� ����YB����U2��T$��Icp�ދ�v��}����9��O������L`i�b(+�\�~����\��5t,�s'\]�*��{�ECĻ���ųU�äv���UԘHOt_w��_����_��2_��Ï뿏���|>����MY�b��Kc���l�^cGjź�7)�{A/mbT�X�b��p�xG�<�;�T�䲷�s���њj�&h���-�d���+�5��ݢ�q�nc�(�j�"]���z噕:^xȬQ�xl_�gx�+jY�u{�G?��<*w����a��m�cҹU������dq�}<^���J���վ\�{��[�[k�	IYR�q���T#�l������D�M�F�]
�]��Ѓ�W��1�Kz�n��U���S�ƩVŗ*���45���W�lf�+)�wy.��g_n� X�J�ˆ휞�� ��<=�� ��+%Z�+YLڷ�\	�K�<��#nq�ޗaבd<�� ��Pdz!�e�ұX���FV��7?@T�^)������L�"ˇ̄�ET^=��6�f�A�� ^�^����8m�Nc/�[�c�B��5�R����?�[(�S�G��J�D�c�W���}y������0������s�b�e
7��ދaP�tlS<!	��C�����LRv��e6��ͪo%oȳ-���RŨ��,2*
Or�h]�Ӻ�1��E=������)�Q-��M#����܇@yA�!B�z��ا�����^%:�
��5B*��d�>���zz81�����B�K��l�ˉ�n�o0�����ƀD���BN�<2.Pn�cA#I��������ދW5)~{�?"*��x~�ᩗjDA`��c@�H�^�I�o���*�]?`Ż/rv��N�����/�k]���NZ�w��P͍1�uuHLN܉:v�8�VهCE45SG+�S�r�u���ʂ�t~n	ĸx;�CR����h.���ls��{��<Z����t�ELo��~��K"�̬8(�p~��C�$��;�N�T���FJ���7!��;��
ƫ���U���b����]le���3�q&�r�V����|�Q!���$���fn8��U��m�t��,�����^ͩS"��a��K-�5�ntS���t?����ɶÝ�>�������}����o���k}�m�Ta�,��T��Js���@��G��`d0��9��Tq��.�\��a�u4����B�a��u��sԽQq�e�7Pȶ��6�O%	D;��׊��z/��!�y�vmt���ۏW�6��Lm�u>o��k�93�z����e��m�Z�yz�kT�v�*3�X�A/0��j?W�d;m�"��c�C׉;�ZK<2���A���D[cP���� �, h|.&%M��mFk���9������瀖)��f���U�$^�4xb�OS���o�P��xg����!�Za�z�x�Fo1�Uv%��VZ�&vж^X����d�@���/�2���q=sͼ4�yg�b9���	��zi;/�$��2��Ŏ�:�s3�}��dy*f�;(2��q�j(���6��=[¯t�wh/Z2�^�-�.��nA�F4!,���y �H^k#�0�cӱ^������MV��{
�q�{Ǣ��sc�s��ųؑc�Ϫ��/����0D�9 �}���p����'Ĳ/~)M2�%��玥-�i��F�J��q\�1Nz�+z��H�K�)Y�ޖb	�����/��m۳���g~Ե#�a�ٚ����L�h�(��nR�Y��^`H���T�[�ڻ`p��K��{X�E�8�gmǊkr|�K���2�� xFF�g��������o7� �1���SOoB�Ͻq����[��
HQ%ٲ�/	�����vI/�N��A��=��U��f���ź��H�T1'�cdv�j|����G�f��JY��T���za�ΘQ	�"���c�}O\s�ͭ�����E'+=�"�-�a�@�az|�>�a�<��D&��,t�K&\�+�Q�w�>�j�q�=��a��a7C׸ŧ����E�u(�50����ь�DbzĞ%� fe��qZ8�^�9���\�ՓM�;Us]�^(�5�������:LK�@�j�R���7j��g�N�g`��@�`�^}����\�	c�M[]�J�(��FM�X�>g�Q��4T�{��xM�i��_�vc���na����v�E��S�~}�2)Xp/����ƧVŋV@l�f^�5<��O���P��M�L��N���!1i�>����hv���͘:���=ۭpPnSLM �Y7
t��^ø�v}��9g�V�m!5�N6�5����EuS�وv�t�	�]��f- ��q �/��s�"]�ӳ߂�:q�؁*~��"�ۭ�r;�m9mK�c�ʺq����9+wgz`�rr
��ց>��ƲJ�iv�n���g=��  2����eEӃ+;�,�C9Vc��qGbY��)�ok9L�Q�f�.^�m�֨swo9��̡������վ������6y6��ccc����ݧ�ơ��7�1E�ę��s�z} ^Y�i�2yڼ
�d�&a���>�6�Y��&�a���詴%�	�兽Ŷ���z{=��Al$P!-@%�CQFq�Mg:j�I�m�|�
ېP-��@קx��d�S��n��S;!"'b}V�΂}b� �ިP�L�gd�AMz��{���;Ռ�u�5{*.P��P.lD�R�<�5�pɄ^m��$Cdi�fL�%Gt1��K��%���+��,)�-�Ʈ��u^��y[��Y�C��d�p��)e&�ӆ{�6F'lb�Ũ�I��N��BՉTS��#gOd[B�Ӎ�DcX�ik��Ț��ǵ��u]�8�
*e]��COb�m2�2�^b��EK����G���B�EF45h��l���8ףPHP�i�!9�� ����G1T�z��'��6Ⱥ,㛆.i9����b��:�_A���_0z�v���P�/����QR����Uz̦�45�)=V�B��U)�sW��g�C�b��/MC	/��7!��8|m��� &���<�|],`�0�̺����S���Y���!�;���ӝ �b�\ڔ6���5s��\���@7�y[�n)FlW��a�[�{v��%��M�f��g2�Jڅb����E�w�n�Ax��j�g]�LP{p8�X�S�|-�yR���C��rW�v3��u��smގ[�����}u��{���=x�AM�r,�o��������z)~1����F�M
��tru���͹֒�N�^/�spy� �ؕ�:�cҹ�x�%�T���@��s>0p3@Cc�pP�/D�Sӱ��VSA8ݬ��K�ʖe����&��)P6˦��;NW���,���dȗv0:�5��m��H�LV9'+��j��am��K1NloK�N��$�Q2����i �b؃s�3�
����՚4j�)�
yw�X0%��%�F��#�.À��!��$=� ڣG;��4���4�iS�С����x��X63��@��e��d��꨼{k6�f�A���7�e������������X�B^i��t���u�o��~4�
�s�#�sÇyC%���L3X���� �ߎ��fP���p��l;�1P懶)������K� �;f���ڹ�Fm�e}<���K�B^�5�	��T)=�;B�t�{������!�/q͠[��g^�3&�2�I��~�����Gb�m�BS$���0L�|Uy��^��wJQ(�ыU��6�@9�����w]ۉ@�N���˛�f�w]y�Ӽ�9���i�+7F��6j���Ʋ�.�/mw]�����̵	�ΡV����Ȏ>��Kn��<�;2�)���z��O9q��/Q�bc��D� �Ed��3�"Z�9CT`�U�|�1�y9�3֪!d�B���n�.����r<L8�-�u���D9�j�ox��<y!c�#x,��5��6����⦳�!��C���{\R@k�Y/���]u�]��d4I�wgM�*ɗ{��%�0ul�[c�Po*>5�׸՗Nv�-�Y�V`�:�j]RG���g��X���P�t1��f
�}kC�Bi�]+Vif�ݭ7t�g�gXK�:��� 㫝Z�wS��m
�@�nvuvYwײ*VpuL�.���]����lʳ��-��Ԯ�j��9�*�*����b��p�"��Iea4/4o@��R���i;ǡ�u�˭�`[��~82f�3Cz�N�ov�T�,��_5\^2���ɛ��+�+�Q��'d�:��J�2Ƭ2�/����V���ܗOo������J�ܣ��b��W÷$h7Q�a��e�[���w+6�Tϱso�
���n	Q)Mؠky^�2e]�m>�wpZT��6�_uy�U���|�#����B����}B�,`��qǚ([��;RU]�S�k&�Xmq��R�fGe�e�su�a��U���f>\4�.��Q�Q�=���.��wl�n�x���D˶�y$V������L�|�k@�9�$	S�
��Oo+_Υ�\mm�I���{���`ܝS`V��7�|6n�:��vii(��̏{4,g.��c92���<�pt�^p�z�u�-��׭�A�1��Ƒ�s��ݑ������HB�Z���F���Z��R+FA`�ր�O`ݭfT�� Q�д���įZ/���ٕ��/�7E-�I�@^����2s5�9��`8;�$'t��[v��a�<��*9*i�\\VU��X��$���n�t��,���nÄ=Z���x��^�c��t����D�nWk<��||�ߍұ���:4���w'>&ٝ��MK^���Io.��Ê=ײ�@�]k墹�X)"2�ł<e!��m8Щu�En�����U֓9�ȥ��f�����,{�����
*/�^Z7n��F�x㓰��\,���h>T�c�ח��7��'�oi2�ƍ�7�ö8��lrɚ�p�u���L�ں s��T��:OK�B3-�.;���9Xk��AҒ�bDZ�1ʂ��K���Q��r�7���E5�8гD�&_\Kkw�sk9��9�-2S�9���/\��ʋr�+�s���7*�L��[s75�D�Q�ufe�*7�}ػ�_�]9O=*y�kPP�Y��{���yH�/-|���$��[�r���I�Ymf�;.�æ��TYܗ9+��l=K����(���>P��w���>=y�w<�߻ࣗ#�%y4��s�
m<�W9eȨ;�;��Q�!�+:s�w�L�	Ԣ=��o7��|ޫ���Ǭ4�|�r˨#TVm(�)$�V��9OAE˕E�,I"��n������S�uܣ�TkYUUTU��$��UU��:�*�H��̪���ʮEA�R�K�����V�	Ȫ̓�q9�(�Ufh�Dr�s��*��\�9Z,)�Q��m*���E�j4�)U��9UfrN�Mj9�d���eED�;�f\�r�$��+� Q^�&UdˡuLȢ���>��h�I��Z���B
�"�Bˡ_ǕW����|Ny�Ӡz��Yw7K(�6Q���QL���"�*��1*�"�"�+x�s�e<`��Nt$�2�;�*�	̣��C��tJ���(&Q\�R����
��{K�K�|K�C���s�x�ʈ����%�r���(U
�T9����gڔA#�Uu�$�Y��򜄽�3�9[v�t�I�`g<�BJ闙�c�WZ��Ts�����K��~y���￟����1��d��>� {��S�����#���|w�!�ǘtC��'�����^�{ze'XĲN�<��͊B)2�א��v�s���n�*`��놺�/�_Z ��͓��s�TƎ�ȕfS����P�NE���݌W����)��L��T7W�wzേp����!�͙�<!5W��&4w(Q�|��D���rү�;N,��*�z�XE���ҡ��8�u����{�0t�g앎������?;b؟��!qΰY;B�Ê�2�;�Uҡ��@�z���sz��0(��M���;m:u�������SLz�U�V�V��=+��T�/t��B��m��l�).���6�[{YE>�����B	y��HɆmǽ�=�*�eO�Ǣ�x��'����//�im!�����϶3����ξ�vO����"�Q~�1�I����{�7��%��[��N!�+�tE�j����` �� ��\LK�6^@ڌ�K8�s�m��z�-���/-+�c��Q>p���� ��]N�_E����~��g�!��Ld���_�0O߫��4p?b�zbsLu(�,���tS:�Sʔ�~�_\�=�t|۟O)%,���P�*DZ�Ȏ�x�ysQ#x��|�T�׽a����5���	��{�f.�o���r�����6�*�/7g`w�,��^s���sNR��t|&
�9��o�����_}_W��_��a�xxx��'��������hsf�i��,:����dÇ��O��o5��
�\K2�?9�*�f�}�O?p�լ�O�U>���ɛjrTͷ㲃%�l�!�l�zǫxGh�>-��H�n���%߃ea�^}���AL��|}�����)A�W���{
�q�D�9w/��^iJ��P�����u��fU���`�����ׯ�A
Kh���Ƚp�'���z{��#,R�L��*��6xO�n�6���N��~O��������vI/�(tu9�~{��n�y��lD�P%�y#I���7'���gG��ki��m��ʙs��/� ʬ��-bv�0�L�I��NV�"�-�a�^=]��y�s]�N0��D`M��^"�*U��u�j�PeGg���0��0���q�O�y�o)At��zC��l�&f����=G4.`W���3�	�C�"�ud�u��W5��(�R��^��砟�vr$	�Mɛ�ʍ��z���}N����� X����<����U
�V$Ȧ4 ����ޔ����&����x�ئ�
"?e~QW�Vţ�o��(*졅�dW1�/6������E�*X�k�XӽH�0"�q�G���<���|�̏���������u� 5m�2ϖ��N�1\J�Ή��SVqf��۬wm��8g>ݬ(�{\�)�'SwqV����>������ o7���<.���j	Kvr����2���<�P�Q�J�G�Z#O�U�;>�4-Z�L:���m��w��ӱ��\ĺL��Ĩ�j/��:�;t�0g���C�-b[�'��Z�"�~Z�ur}��xC�J����l��S@9Êq6��:m�{�9�=�9��`PY��`��m��m��cu��˘�-��8pКf��0�[I���^���l�wl-m�T��y�NC�f�sCY	���ON6ۜ����f�L�v�T� Ș��[�E��
I�m{�V�\�w�`�(F0���E�U\���b��l$P!-Id��S��1�"fR�O����z3�3lk [?<�zw�\e����n��X*��W;m@oB	��Zg�:檈Y����:�
u�%�ǫA�]g�����@�W�V��?�L��ˣY7n�+,�[����/�3���r�Cn>��rpȓy��ˋe����D�Y�����_^�d��8�<�Z�ݕ��!=�[����9w����*�Z�TS����=�Ы���=N��]~�2�p���]D ]���S
�fEt�`M\��|����B��kM�\yp���.d���Ob����j����;�[���p�Np,{��;���jG��k�{1�����Z�%ð��7)���h�_"n��A�t����`=��=�< �E-E����S|!�C��tƇd� �a�iiRe���_<�/Iq�o�Ӆ��-��bl���Q�k��C�@��c; _��A��,�)��}R�͎3l��/�&'L(F��~��]��ކC��5�Aܳ�Ϝ=�-y�!�������w�i0���\��7��`+�2k�h�=m�ή��)L���C	O�ێ���������qx�u��г�����#%$�l����\�����}�n���׺�^���p�����6����*��g:q��Ǫ���!�_�(��8��S�=2���X�b��x�a��̺D��j�;�˳�����@z�U�R̶�����@e�"�#�;NW�Է5�,�j�~kՈ.kw��ʵ��gP�t��{XS�+~�2��'V7�ۧ�r�
bK�,ݏ\fa��Êݚ�}�,�+<9��Ġ[>��˺�Pm`х�S�
���G7��E�Y5�A!�.��{ghE_n�i��C����a�i�:"۫�ok`3>e��DfJO2��M������S�>����%̻����q����6sL4�ggG*`�E�-X��z����|�<��-��nk��uyM���0��es�UEy�3
y�R��p�ۮ-�LV�8�뱼7dR/�R&c*���Z�k�h��v���}�~^y�~��w߿�o�����;�����Ll9�����i�c�[䠎zK$!H��H��t�u^�x�, Xt�O��h���)��)ȩ�J��$UF!�l�*������κ��e
6�p�7�Z,z�SW�_���th��.���6$�1���5k=8�vGg[�l��Є���!2X�J~��B���{��m���YG1EʖL���q$>Pi��We{�C׎�,_D&=��)���L:*E/z�m�+��3�v�#�?-��Z8�o���a�����5��q2K�/Ŷ�l\�5�񆲲a�m%�{kYƓ
~��u_5��	�DB`��{�cGZD��'}�g/ǝ�����fm(�#�O?0Cv���<7o�mC*:��
E/�~@`.��t�����F��J{t��o!:�R�^X����Z~k*]&���p�v���z}�d���|�8՝��ڲ\�{��6+����58�� t���Q��j;�M�T;��������l��gBU��uM�����m
�K�����4ںd�2�%:�x��{���ߩG2��m���	��g����הn�u�j��Fw�p��
V�v��'��J�����`�}`�X7+�U�Ħ��>L�ٙ�����{�{�l��1Y��W���a�>�sA�#5:-��#$�JU�\0�,�~L=kZ���i�+��w���)�j*w�3sv:u��=
�͝����}�� ��:�t��U0|����ö�i�L3n=^��'*S�Q��~F}8�ݦ�'��'h�t��|�X��6׺,3����p����<��{��2~�3d_���t��[����}�[uV�}K�C�"�&+���-���C���w�����e��Q��fn��d�	���6�Tu���Ra���0�z!	�.�i�[�F�T?c�=������Z��غ����i���^�xj�͛�Y�{$��+(!A0��b���xi����V��X-\�85ft�X[tcB��"������O3>�|�6Թ*f�eTN0,Q�y���a�%UC3�:-g���o���"��-�X}O#''��ª�	X����BSe�R�&�h���`��n�(Ő<U���GO��L�r)h��V���ޚi�[��d�,T����l;%Qj�q;Ϯ��vi���m�8�n��4��Mn�om�L��SۼH02@Q%ٲ���ۦ\p�Y��!��v\��ki҈��_���ƩƼ����������� �5���5.*���!<�^6g[	��\��hءҹW�ot�CW}F��"�Nf��E�P&�5�Nu=���0<L�B;�P i�w�9�ݔ$3)�2��/�M���5jZ��z��Þ&�|ei��c�t�}�è�?�}������Lwטl�{E�}����o� ��c??>��������������}�);9'z�$�W�����(ז�0��,�q|uХb���4����:�f���p^O"5�����ض��uL5�M���-?,O ��P;��3���")��]�}ЅN�|��֘t9��Ĳ�ՓM���\׆x>Y#YK���cm��uBS�:*�Ѭ&��N�!�wh��!����;�'��"y���ƄV�czR~fUQ����ּ˙�Ny�ye=N@��lקv`763��#�?��v�E�uCs��B�>���<�#�e_cF�իXa6�����I��_l��#��
���Կ�:3��/�v	�]�.�ͼ�knԩnMk�ƃ��I86�
�M � TQj�~�Pw����Ĩ������;�
α�#G.d"b��ꑬ��P~yÆ��.�2�ZI�����<��hH���U�)E^��-� C�j�D��t,��m�;���i�kL�v�T� ԉ�l��%
/������g=�f���N���Dc{�d^�Uϫ�6+��@��/�<��>ڿźX���R0*	���B�guA��6>wݻ�I�K�K�Enn-��k:+t%mhԂ�b,�ۧqԗL�B��uE[I.�]Ӱ2RUܳ2ޢ��K;���
Ɠ+4�[�w.�^6K�L��]���+�W2��g_U�86�{�;r�_}�~���7������e����T�����m��mޅ��d<��#D$���{`��h%bv*�o����S���4Tj�h�}dL��@�4WV��1��Օj�38A@��C<s�]��TDN�gk;���>�����2��c!*��rc��\��P�r����-�ơ���� ���b��'P����=J{�k�iA�9;Q�v�=����D&I��N��&�j�*�qw����ȶ�-�}	rȝ�uչ��'��B�[H�$8�P�b{�N�T�`�&*�<�/Iq�k,��`�8������j�K�ռ0�� B#a�O�� ��\C-�8�o�Ry�ȺY�����F��,��E2�-#�{\�	�x�F¯Q��_ԏ�w]�}`�l�&��9O���@���Za�xe�s��(,HGj&wvj���>6�M�@Mż���t,���z��`]�ܪ�-��>�J�]�J�
�ΞcV)V�Mrl���V�`�C�w��v����]��t���]HL�v��yD�q�ǥs��1����'��s�j�*'��&��nܽ
A����äH���������34i2��ܦk�ʙ�5���G�.�%���q��i��̞�3F�z���)��d�7$+6���\i��j����g<j�>����� ף"����.JР����H׊pW����,@
_ō��;l� �}�}��|���{�=?O�_�Ai�ݘ;�ѝE�5=�,�WMc�wh�j[��z�*]7��]���c�/Yݎ�V��0!�z�@x�X3���L3$��\L3�9E���L3m���퓠�w1&�#2b�v�Gރ�����U�����_z������(��pT[s��{z����9�x��_��L���[�]M���P4Piza��eC�m����	��Yq>��I�/ٖr��Ǵ��j���"Й�[���,q�/�d�+Ț�M�Ӧ��������I��He���s5j����d���ձ�Ly@X�� ʼ�(Q�����H���46)�!|\���^�-���]��L&��{L�%s�,Z��BSe�,R%?zWm�Ӻ��rF\�"R���|Uo��`趐�I��x	
��}ؤ�t!)���N��L����:�>�����b�iͳ��_�<RC<7�|w���؇H>SL��h�!�a�oD$���V;\MRx
Z�{g3h�oa��|�	L(Tt�8k����� �6;��e�n'ZD�T�4@Yf�+ꥄU�w��%���m�L�{�r?��7ng+��jP[�f�j�ɨ#ל�`ζֻ�X��Br��l�A�A��	q��Aw/�Y�Lw�/eJ@SR����wmk�ܜ,��Z�^b+�T�J�'M+��P�Q�Z4�S`齹�_|<����xx{��S^�Jv|����I����J.��)�-��:��p���PP͌�7*��6j\;�E�=��H����H�q&���������]&��q.��#��k�3��w\^�X��}mF���5�`Z����%I�>�Φ�P�z�&"��8u��m���G�I:�8A�,Žk��Vںd�2&Uk
�ҹ����{��^�����Z���o���S5 [�!�?���k��/b��Hنnǫ�6�ʔĲ��̽�˘���kv��4�û��:�\�*,3���8>u��`,/E��P���̪2�΢�[�=�GZ6�y�zt=D�^}��b��!���t���𸘕6_oy(����c���ީ���^�������K�H=�$r�v��o�؊��Ȗt�5��vh�l��q�yw��\����Ԙ�{9�C�sp�4׻$��B��p�/f���xh�fL۫�ldqY���`��R�a�ז��d=r?��݊��m�vPeAd��Q��z��v#�{�*IV�eEy{�}x��]MR�Œ�g�a3�N��Fʹ�@��oC��j�Rn�u��; n�ũe���b�ת�l\�w��F!�Q��&btܱ�ң�f���Z��@/LDf�u�5���C-�@��)�4b0�'\tWeu�+�'�ta�pz�m��F��湔�m^�[�F����/��YT�e2�A��s���>�8�3Yf�앀��sB�y��O�@I���d�����)c뎥�is�j���v$+f�)�kxlw�^*�N	��uWX��ݩ�V<��Y�'AH�a+��ݳ%Z��^�f����a*�}W9]��w<����A����L�/Pye�t�!Q����j�*im�ޠ�a���:�S4掫|�d'vn6�l������츫�)M�yHR���;����S��m��f8�u_�������F�E�R�M�Xyl@�:3ϓ"g1,sȚ�g%j���%p�SehՋב��`��)��ͬ2]j<�H<�W-ʾm��WM���*�5,T��u$�;5�μ����W�Iy+6�k	�wՂr�u����qL��ٍ[���%ԭ��P�z,9�C�qk7ݸ�ˏ���U�scG�h��*&�9� Zg�f����pl�|%Ȍێ���V�a�\��!��E8��{S���VִzG�]�|i�B�{5VeW܌D����u'Eٓ}�J��X�'^안�qs��xo��f��ۭr�[���0��h��V��Ďܨn�d��.P��y��y��ԅ�W~پ�o��Iڬ6f�m0^� �N����F�v
�kG���La��b���uq���#��r�aƆN�WK�.��)�9^�#�V��%\YڐrC>�f�W�撮Y7:)yO���nQw\�������s<N`�,��e�$���\�lob3��e$�Z���NB���v��dt�a�v�D�{f[HQ�Fz�R,uf�p����|K�5���j�c�5%�j8wX�����-�R
*��.d%5�G�iLԙ"V��O$��&��܍dZ�c:rNCF�@8��@!Լp3n4���s�sMͷP�&�Yz#?tD��fJ���"j��LO�W|��	`rv��ǜ+����S9��U�0V4�a$9��H��vy����c4[��|_���[g�����3�W0�����WKzp@��TÂں����Es2P}ts����w�j�Ϗ�\D�����qZ�8`�5��/Vȩ�m��&f�7��3��yk�t�ڠ�/�&��k��I^kzZ㹷w}hm`Wk��ɨ$��'����󦕫�tr���o>'#�3�̻��.V�V�i���[��M݂�k}���M�D0/�� v*C��f��k:��TB:�]ݪVT%��c�Ʈ�Ok�h+'t۶K��+��Cnɱ�`�OK
q3;��ɕ�Xy%��˸۵Y����q����32������(��0��B�>Gt}�\�^��AU�ESؑEG.W��=�þn�o����>HH��94�Q=Kԑ���]�9N�i�PJ����=>N�֩�#�Q.'�#��rus9�+X���GVh�r�2#�-���z��
/�9�9�^�^D�L�F�r�L�{�H��twO�%�~xw��yH��(��x�N�˗L*#�Q�;��9EUEQQW)L�W|���!��?:�����B΄�VDG �Q=er� �M8r(I ��9U	Ќ�(���UAE]3�Ĵ�'�?)ȎS��BQ$*�#�U���p�^<���(�-e0�#�z7ya��_#�%�D"�*��+Yr����*y�Q9��2�><�eȂ��>��y����]���<9�l�]��'��nuФ4eoP�c�1ne��0��z��QA�j�=ߗ�???o}�}/�ۮ�������6�Cg!������f��~�|��ռu�)��a�������~UZ�+���7���|�LcY�hٚb���1�w��7oӱl;^�ս[�z��;ǐP3�����dY*�@�|��k��1F�:�Z��6�K���(FSS�[�p�t��{w�\bx.�{�xLD�CE妤2݇U*3�͏�`���]%�r�	��"��F�[_�ry��.W�= �5��^2�D��9t�rn�p�t�H]J�a�-9*HޥI>�NW4	+'Xkх��<�m=��J��m�q_c^����AȄ�fn�;g��QL���-?,�O �������'����f[H��V����?!^˩���=PS���5��G�e݌2����^���2*�CO
��ц���[�p�ûWF3�C\u�~�����"y�ĊI�l֝�b«��#��yl�u�"\� �oWJ}
�Y�^�ٷ+P�}G�/Q�����WD8ꇳ�m�m���%���lJa��5��������'���JDs���~�<��P�C�ɶ�_���{�?W-�o���5]@��WCrd�@=*��M�w|�U�ʹ"�_~\�^;�}���y�����G��b��|-^�#=�5��U�c�����u5�"0]%YO+NM�7�Z�汎P��b��;y�8��՝��.�[<G^���4�l����>�xx�{���F��4��Z-���N�T���I86&�+4��<�П��j�{�����uu���g�͞|�׸�GB���v`k#�!��Æ���4]��bľÂtE��=�u������MUzY�Z�j�xՒ%�Cd-�dL$�:-����輳L�CL�v�T� �Dq���1.���[V�#��C 1�Yz�<����c�	�#C�["�Us��͊�Z��C�c�¥���Y�&��CS/j�A��L�=v�c-qL��K�XP2pAO���L����p�bJux���	z�X�l _Z��	��%�]8Ϧ:�����z�3 �]z�Iq�9q����+�֕����mE;.��M���B��<�G�U
P����-�ƯuEê��q,Ќ�M-W�^*�m��Н��l�u4�.�7%�	����'.��2(�%Q����"vi�b5@QԶC��;���7�'�����i�+iĐ���.�4�sfw�Re�HLVsȢ��Uʙ-�4����e�����P*�=|��� BF4Ð���R/G`K#�a��y�/�*	������!��-Mc��J�i��e>Wf�6���Sn;�µ��.���O(LG$��"�cX�Oޥpm«(K��eY��l�7ȶ���τ���+.�޻��Qu�b6Y�#:�'��9J����dW���[�4*�;���wY0�~����r�������;��?����(�]G����߆W�?/K4�������� �kτ9��:�����L�#\�Ӗ���hk���r�2�˔���Ib��0�'�vh�2c�cn0t�17e�-��t1�/t��:��K�WBչ���w�<�����m��Z�B{���z(;���Z����8�q����O�����
�m�� ��i�j�J�a�J�T��%A��E6���]��|B��B͞��$S��gsLZ�CjY��΢Ú���&�}��+ÍKs6�֌�qZ�Z�6b�T��.n�+y=�s#dK� �<{D&��~��fI��K�O��^�畒���k5����ؙ�\�D2D[.qL��^����H^�^a�>0�s�N�v����J�h��ͣ����I!�#�t� �醓�-����5���2�.&3%'GI/��_�ÿn�l���\���{6��(<���Y!
��H��t�P�Y�� �!����l4��<�k�sZ�*���T���e���A��B�Ru��ޜa71P����0�r�R��C����u:k���GM�QABV�[`v�jT���m��0�N��ck*f�ܻ�;������D�r]r}ZFխ�8�×5.Im��E�l������l�$�(�� ��i�A��������:���qc�U#������`�[#��j��R��G76}k�d	Nժu��u�.���!)��T��b�)�Wmzܖ�q��ǺV����Y.��V�����Fŷ0��h��<� r��H8d�t!)����'Hb9!u�z�o��S����9�����C ��!�Ǳ�|��'�v4'݆��U��C����e�tD�묹O�òs��-��y�)�FS~���s	�}iٲ����1���pB��	en֑�ь�b�Fta�.�`;R���cHoT7P1�����54���f��Gx�'��ض�������	�x�P�`�(qT*�zb��_��Ƽ�L?5�\9��l�g�ڹ�J��p�cf����~[vbK�jq�c�$V�Ta��w:��w=,�|�b�����B�W�xK�ުp�O@pށa��������4ڬuQkejUk=\��z��}NZ]������e���Q�`��7p��qy�;k��vm��ޛe~��1ۤT��K&t>��~y�����>�zL�P=r�h���|`3?�D"�ѯ��mC'���4�;��(�w��Y68zZ#��K+�ѻ��~��R���V+ϖ=��u�}R�e1jV�M�'�c~��"ӛLu9�-�7����r�Ιt�)��2<�Y$�I�(t�w�.v�)0�m�8+��h�!J��a	�WDw5�Uۊ���N5h����{�y�<�`=���C�~�G����}�����G��$8��LW��b�:�;�xA��cX��s�GvU��;��%*ǌ����䁛X�K��	��'�S����gۙ�!Xl~`h��/&��<��{�c�����\sH��=OE�����3p�4�d�^+(!Hɇ7�i�1�����l��F�}{�X���άF4��a4�FS�S��ɛe�K6���a�Fk�GL�,;Q��������Pu�3e�;�K��-�Xt_##��L���b�;�JlT�z���8��d�E��kCS!ڍZu&-��x��z���-�� A@���d4��d67�4CH�g����lv�B�ƫcŝ�S!��8�q�d^�Ji��F�]�n>5s�:y�� ��Q%ٲ$�яƲ��έL�J]k@!�Iz)�|1�ީƒ4����C�\:����h"B��
����<��MԳmuIh�'%C�ԩ'�I��sȣKk�sQ���)�|���.�f�����^s��
��A�`mK{���Ƣ����[����1i�g��%�gQ�ܼdyn;&ү��
*f^�C��s$��k��Wc���2��lӵ��Iy�d�cR��r��-��m��W�|���T��5�I*���,�MbI,Ǆ����C��gF�3)�����Zi'/iV��T'��h���&��GCk��v�l���/7���{޻�ckQ�C���ｊi�q���#/'�r@Ȏe�c�&���W5�E�mP�ɮ�f&��or�.��z�|w Ļ�tc;l����a�?�\��Ȧ4��D���l!�f���ZsT� ��~k�Zd�ՊS�QٯN�ۻ�����K�F��6�Ṣ̶�!o4��~C����h�&�,t8�����s���P�n��3���5f��合�We�Ylgim.�T2}��h?P�I86#4�_�M �Z��M^/b�� ��k�9�������)��s�\LsoM;��I��c�`���\�t���Zܶ��X�Z��s�X�<�Ƹ}{�-��&u~��m�9�>��4�5�O;MR:׳ohԢ[:��A�Nz��ӌ#[9���@�{��c��["�5��y�͡M�ʭҹ�ڎ��h��5%�CP(�3�͛e^�ΞG=;��`fI�l���7�-ۧ�Q��l����!>����O��Lhլ�u�6K�9�p�N-'��\l]�z��,W���ۏ����]�e�<��7᪊�w�NB�P�ߗ�V�{<׀J�cP��b��z:��q������o����;P8T�i�>��Ij"��U��@/���sd���eF)�VL�4�̾�gu��� �	��eBŉFb,f����������禴��kZ��.���M�P�:�Փ��A��,�,2$��a,��'��[n�^��vi�[��\�t����k����ۇvInj�'�)Ղ�W*�qo,1#7ј`VdF�ᝓ[Jzh�o)#D9A�Ð�d����fzT�\^b�2rp_;�U�.����������+Ӆ��-��>ѐ!"�@�!?P�Az;YP8��*�tm�8���qe�G�G�V��ru��i4��vk�����|��`����7s�M��=3Z���L�߯5�Λ��#�@b�¨Z��G.Rz�T�4��0�� ��8PV���q��0���L_�";P�%�)�@�l9��.��Q`�g.k��[��GC�����ee�L��mF.ƾG������t&4T�m��hZOw1�\�⠗��J�\P�O5��~آ���*¬����C�����������mK2��XsP`2�{�;ND�լŶ�1,�z2��<����c�s�g2dK�p0�g��@x���R̓���Ӈ(��5�5��㷍<��A�7��"j���j0�;.Vw;���8.�v$1p���[�Y�n=��t�vv�v��m��&;�k��kW���A�e�wfя~�ج� ���g��vC�8f9����7�E:��]C��\�vh��f#�����KL���?�o���No�Gy�_��G$?�?y���o ���:�I��v��o�q����-�xtg/:��q�D�y���½s��i�6�|��5�:Ȩ�N�p�<׫y�C�����I�ʺ&��k�P{.6j�+bU]Њh�u���t:��ME���Q����(<��@�W ���W��s�髦.Q�g�j|Y�-p�Lp]Uѡ[��q".��TcV؜�kj<d-{;2��B��G�>�[�d��5¼�]�ts쫇(�3����C����	�m1����b��Bk��BeK
O1W�5E�Q�����[�KOwE!�L�4��]=��	�!�}/!�>!��sЄ�2f���Y����*��:��{��T�	�T.�g1�k�<'�|w���4 ��0O^�h�ٓ �Cb`���kv����x��ɕ�p�K$�tS'4�C�_8k���5��H0͓�.}�C�O���]Щ�(�i��z��J��0�}�0�r�E��z~ވt�.��CJ�F٬x�u���K4�Y�?�>6 jBbv�IӴ��W�*�z�Z~b��!t�~jN%è��+[���c�6'c�b6������m��Z��b��3Ƈ�� W�����K��\��if�ɵ���{˂�D��w**F�)��*,޸�'��Yŕi���͚�RB�_\�m($Y��s�}�^�YZ��:�N�նAov�}G�]���2�kNJ��,�}_W��U����{ؕ^�(T�������ƟB��6��� ���t��*�=Z��Sb�眳Y��S����{6�gU��T��� ���a��p�_�b[WL��F�ǥs���ެJ����K�k�6w��3��4����+y�:W**����v>�M[0���|f۶����71�����s���K�S���������,Ɓ��d�f~ƈEݣ_ŔpEP�,�e՗�V7�L�~M/�ݲ��2K��1�!���LW��b�:�;�xA��i��g���6+5k��Џ8x���uFk��h9�3k)~.�~�B.�i�[�F�P����ݤ��L�����y�V�C��@X0�a�=zz/��ӛ�������dÇ���Bʳ-Z{�U�QÝ�
��O5VPxX*�~?W���,��R?��ݲ䥛8�q��]�z���!��XS/;A�پzǫx]]�`qm���W�Z�+�^�+�DFj6��ӯ���m@��ɭ(��v-�=�V�o��
7ʹ��a�$�gyf݈f��c�k�f����;��BM�P ��kX@��$oV���[��1]�J�n�p�vwS_r����]�{pr��8:=D	pT����{Ψޮc�,�Y�N��)'|�jsI�^,��*T�����8���������xx�q���fL���&�Q�!8�Q,��Ji��4��Dn>5{gO"���A���ϐz������]6s�.�f��x��@#{%���'�b% �ƩƂF�[_�ry���^2��m:!�/���sz��W��� �f�S���`��q;ԩ'��NV�"�-�a�Z�{���w�WiW����B�u�Q��a��!#��B)����wl[I}T�[&��8ŧ�T�B��f�eR��]T*0_N�a��|�S��@���L"A��F03�
9��q>ىe�~�ɦ��U�{D���\�Om�K��5���I��t�Ļ�tc;C`t����D;'�]T+��®.u� 'sk"����P-��5U�ߴ�O�kL�z�J}T�6VŻ�n�����ɮS��n:3��i����񎮡���"�x(�Á}e��z}[~������P�n�t0l�"�D��2�[�Ɣ4.g^B)�H�M��]�����e'.�`QM �Z�~�wB�4!�=E�h��k{B��Z�;�gg^���H���ojF�W�A���pК���L3�U
߽c�/�e�3�{C5.|��LeMo��D郷�e\0�4�Z�j<j�r�P
'�%��!8e�U��ވ�b��.�QXۢX���.&�Ģd'*�����V"4p�j�2�?�F��Oh�YN�����b�.	���=���Β��R�{�<���P�����l�q�O4(u�D��P���Kt3je`�/f�2��d�9�y�k�)c�f��ӱ@���N�$�l�_���5� �#c3�u>a�ǆ��lJX�lݶGn����:�ӥ۲�k�̑�;��6�%�Ŏ𬹲m,c��H�O�gu�ڔl_J2F5��X5��w�ǽ�մ��U�5 ��v^vVMp�-)��Q�J�o9,��/�I�si�	{���Yj�^�eV���2�r��x|1Û[��T`���j���Q�(� ��'�rQI��:�k�E�ƺr�{BL7������Fl�8�vҩ��)��p��ιq�4�׷p���h;���@+c��@ӱt;.E�*3e
�o��W,��6��S��Em�
�Y�$���#������#���g,�G�ݾKgv�I�f�Qz�Z/{F�*�g`Z+V�����y=Mv���%�ܧCn}&������6q��i7��S*�D�B�]ݼ�T��ٱ�Y'bw;%nPn��7�Ov���%}��>!��z�ݕ�k���c�J�4$�)�`�9n��⻜�upv�ݛ|�;�Y��}z6-Wv5l ;�c�b١Q<u�[�5)��ʷ�&WLbC�YZ{�D�l��P�3[�j��$�t�ml톀��3h����wZ�l�-k:��4�lN}N�N�G�B����4:���M�tR��9!�(:�F<�s�>7�`$�)��3yh���=�PewA~��&S��ډ<:,�c��%"�Y3mY�>pá��w�e|f5��L_%u���`}�T]8��3�`�t�,�kt�1!W2P�U�+�GݷH8e�L�G�[S�>��	\S�m�h�n���h��
�l%�����e�9I�=��>r��1gZ��Ruet�j�e�f��T�|�^�䞪�ڀ��#ǫ!T��[��ࡸ�	ץ�*[��xM��:�+]�7)��#A�}�Ǌ�.���E�2Z���Zd�Z�t��H�K;��Y-�����+��|@Lep@A{��R��2,愻���٨�O[��`Ңݭ걜���:��k��^�L��tyH��_ئ��xv���;W+�dԳ������M����ek�ɥC��NG�ݬ���z+�W	WN�qک�mg-}y9.f�Jn�Brj�iߖo����^����xm=쉆���� 0e"��sY��3�3_�Gް���N2���jm��6�3�p.DkxA͇6����;�z2���n�\����T�6�]�})�bڍ�a.�W8�����!���=AJ��h�6J��1vvܬ�O3��G�f]�<?����>�ٝi���5#�$w;�ch� �6�_@�E#�Q�T� ��Ϗ�jW+_P�?H���EIm(���a���QUh!�UAjEA��ow�����z�!2�3]IȢ��N�i�Dr�(���.ar;ԇ������7����;�<�Q��BÚ��*�r"�Ǐ��e�ˏ-N���*�BL3�{^P�%���|�*)�^��.c�""��r���A^��wB���&%�>!�y�(�"��u4wn��'&�!U�hI=�c�U\�*���n�®�D�������}���PH��OE���ˇk>�z�|�psd&�c��+�,��Vy%U��3�S�d!J���DN�(�6G���2�G�{��e�����#�U�\�򖴪�QGV�Ҫ)����׷��Q�h,���Ԅ�$$ꘕv��С��w��w	�;�<y�ZI<w<��u� �ּ�G���TXTU�rO�2(�:T(���(�CV_y�p�{�3�޻.TE�AA�U��E�����:{,��+��n�U��8՜��gG9.�}Ϟ�gL�dV�.�B�8�x=��S�����w\lg4>�\���ˏ~�C������&��҇8���T8�(��z�o
��%܆Ӣ�ba'W=8�nszG�זi�����;s=���K�Q�E�#N�� ��Fa�}kO��sdS�{�2�c{����|bx2VU�C�߬~��WJ%v,e專qG!-A,��Fq��f�V@�t�9��"pL�h��=ZבdhM���&�nQ�,1z��.�ثjЂ}k;'��|��Euk=�|jQp���;����7"�mF=�V��=�A���7ON���M��;��r�N�j�JĪ,)��[\���o��F�;��3��W�1�="9�O��5�i���fK��Mͽ�'�)Ք�Zӳ�V�)�I���M5v�q��	�h4N7�A�" �@قP�`n����T�=+�CU�B�7�K[{ƫA<�O@�4���/`;�0�� @AƑ�~�As�!���#��W1]�H�V�!�-C#�+�o��"�x�1sH�f��;�?<���^D9��D�NEt+@�ݗ'+�hՒ����+h����\��r�'��*K�C	�O����!��n	=h,���5�Lp�b���8��Ŏ�Uu��g�(/��&�V�`j{��c�{�L<d��g-Y9����zG?+��^>�-ė���:��$攝�N#��NY�	��mJ#u�YS�f��!om��L$vam�R_f�q:7��Dp�����o7����������?�@��z���5t,�s'\]�TX,���6��k\���{p�;�-ٱ��4�[�{�§P`����is*�����Q+\u��\�9/LeA.;V�1���'���v���4��������!���>綥�m79�
T�˦���l�&n�d�S�ؙ��62�Zz/a���^�`<�3����*Y�ucz]��S�{O��n.��.ݼ���K�,ݏ@q���冉�6:3���.��	��_!�>0U�/r�`:x�geUWMl���v/"�y�2	@�4�za���XD���σ�DKO��ğY{��r�]�����;^%�ޙ�\���yn9��B��S�m��uH�'e].�ܴv��ꋝR΁X@��\O�s\�X��j���K[.P?x� ʂ��J�8~����ӝ���4~��>�
a��Y�B9��C����ժu��ږ-^�BSe�2*���YV]�r����7��F�h]��ס�V���{gh���I����^!�v)-�{��WR��4�EOE��&��\=zY�Sv�^z�+R/�����	�GM=3
��hݺ�B��r;}/Z��Z�f�$������žf���aK ׀��Ck	pg_(G�I~��� �E�%�Of`�	rӯV�e%S�1�e�m��{�~��T�Ę.]����ί�J`��R+cg1�}Ǆ�-���D:A�`���;�#k�)��<�񌆋�-3%:��,���tS���Z��a=}iٲ��!vY��g-�YÖ��t.�U�֑*�R��yN�r�\�k<�%�P�@�S��p����F=�i\"�6������H\�sT	� jBeGr�;JU��^��~n*]&��<�2	73ׄ�>�ξ��o�-ì���<|���F�lħ[�S�9"���B�w:�ӊ�.L_��dR�ކ��"]Y�i轸x�G��`e�G�2��ښmV:���P�VN�2�dD������h�]܉u�0I�n~\?[@nr�G����G���TW�w�Dq����UH�#=ɯ�Z�~�g�[��U&7N�O[�1��3<Ǫ���όg��sw09C���d�����������n���P͐�}$�[����D��1^�tE�j��gâ]��i0�K���~Ȥ�B�5c�"L�=�Fk��C��X�K׸�A�!	���U�޵;Z}������;���7Yڛ��	�8\���b���j^�T��y��vP���5=QM�M�P+=7�z���M�t�����L�h9�7���̓�e�"��N
ܴ�uͶSk�݌k��]��A��q����m��&��rC����;?�����މ8w&e�{*�����->C ���$��=�g7�sf�i�;$��e��7f��g���;\���aìSk<��;(d,WK�����KC�ύ{rfڗ%L۝9	�L4���y1�n��YD���`�����ٴ�=[¡�)�08��Ƚ����B�`��=7*�\��xK����l��Pd�iM'�]8¼z/�i�5��
H��p��t���������s��{��Њ�6B�h��A8�9D�/c�)�W(�k�Dn>5{���ȧ�v�M�@��N�Uhd!yD�t3�cHC�	}%0�O��N�j�Lh$i5���4�h�
Zb��K�6v󟺦�d<�qC5��2͵�<W��v�(q�ޥI>I��yq�4���n��j���2���9�>G�e�[@�� �Bm�Lpm����uL4ل�93���4���]��W�/��[ݠ�AOCQi�%�a���1��
9�އ"
,��t�v�p�!˥����?w�˴�k;��H�R�Q���qxwm{g`�8�������%�	�U���Ơ\1�!hQ(�d�]���� IW��[Cy�8z����^L��7�*3�6ApȄ��
l���״k>-� �2m��ܞ�N��Z0	Rn7�������=�3;�뭻�c���:�VɊ�tp��L/TCY��| ����zc���	C؍Ci�2���ƭ�z0Q�|�ɷ��Ъe�5�7+P�~�G�M�z�S�����dZ	�B��^����u��B��D�A�k~c���_f���>�����O��t�+��jݻ�<���1,�P����9�]��a��p�N�3L���QE���5�8.k���U�����r�O��{�=���v���g�X�6�k%{��p��U�`���y�C^���k[��,��lt8�����O6D��aCFG3ä��Ӎ��=�>���;��c7����7orf�	�NԔ� �3"�Z��瘸��%��C�
�!��["���9Θ�x�+��b��f�y�^킃���A�PK$�(ų��l��3��zw�`��N���-�2ŕ��y�.�@C�06*��+�V�7���]�,�,hլ�c��)�ͱ!����e[�ݽ1�`C� ���0D��e�S�1��p��B��RukU
V%QaLݸ�r�����U��]6��Qp�1�$F���K5�L$���&��Jnj�'.o����Z�W4x���TK�R�T魯Ѵ�*XK��Ko�]|�{�kE��N�{�Omj.
u�����A��K�ؤ�4�ړ���\�ЙN^��(�x֫��*[�%����n'&'Ze�8sY��t(�Egu[�I[}X�B���p��������Kօo$�Ё�����]��0������7�	F4�t���!�\;���0ݽw�O�j`ɴE6L���\�.Gdj��d�sȢ���t�z�o'F@��i�!?WT��q�C-vl=��v��2шCe�L2jJy��m�u��i�.iv'�]����[PA��˱Z��le*���p�A�]E'FnD��;I�PeOD�x��OV
�Ƒچ	�ݚ�!���R�c*d�9�c�F���#+B�)��s��E�+�X5�,ۙ:��qTX,��5*q��Ot[a��>%�x�Ytw���ӇR�Pbʃ��p]1��#�k�еj%k��=+�ʂ^ږc:8;��=Rm�j�#�� 7�N�@Y�)����a���lsL�涥�mgQa�XR�DR�|��P�n�j��1�L=�n�]r�i�*����e���Lw���x!0�#m��'G[���	eTd)�����Nڼ�RaC�z$�Q2���b!�
ǥr���d���Oh��s�v��}����c��y`�]�dpoS��{A���)����I�ʺ&����꩔?���e�q����r"&��)��mӾ�׳UY��9�1,<0ޱ��k���w�һ�o]��N�aSvSϖ�9��4-ĉ��y���-;Ÿ�e���?g
������b����&c�2�4��qw5�iޚ�OF2׷�� zg�W��0��,�OÕҍ�|�_8�����^=����f�O�ij!�\4"k�7N����R��ln�戕�w�\��Õ����q��q�3$��3�q�F��K[W�2���P2�m{ܞ�lH�U2ךLK�r�p��	1P��,��!64��-"2�j�d�f� �<��9��NwDN�-;=�hkRz�'3�"���	�{xjkgk@Ŵ�_*^B�+�3�e��NXS	uR[��s;�z���P��W�j&��	O0MP���dtf>��:�eY�W΍~�����n��@�:PΎ��mU�N��_4'�קze'Y��,��n�cC�p��W����y��־�x�|�Y�9I�jpjf�")�c�����ɇւ�i�<� �cC6F����t��<q�gԫ7_��Hb���E��G7WT�Ǝ�
��P�x��^�����,j�u^����mn�p��0������a0��kLp�n�6����'�8:v���0�ó�
"2������2���J5�?}_�WA�(g��s�0d��sm�`uQke�E��W�*|3��p���3�h�spͷW�:U��[{}�d�"��L*{8
>C�-��)GP� }3%;�UHV�CC��ck�17j����|ǝ�vo�3�"AԂ�i�[A�mq�t�`�n0eJ$o&ei�;�`t9��2u�{s��7�����yVzЂ��1k˔�=����{�(�i�]3m�c�!�p�C�wf�M3;O�V멌7&h�]�m��T��eO�Ǣ�G�j �f5���0������MWY��4t_ ���:���{�n~̀�}(�����l�b�t=1lb�U�x�����&�2���tΫwD=��a�q1*m>�޺[��ͬ`��$�B9u;Ge��8���l�e��-��E?����ȖxBiid�{d�M��Gw�sf�i�vIaǌB��1�)��ɶV_ս���v.F���|geWK��������mS�>3�iA�����j�~{��;�u�&m�R���v��l���p��ʙ9�j�G���X�}�x��eZu���vQ�<&�԰�R��ĈM{�2�&�-)����W�E�ս[�z��+�~�]K�����S�W�������DzP���=a�(d�-Aq,��Ƚ���(FSW��ơ�l��z��F��c�f��G���07�f	x�����K�蔑gK1*�*���.�{tT\�R������i��Pl��u��V�n��u��!s�c���vh�x��x�"��ҵ,�W4^s@�{��#��� e�]X��1�hckl��(��z�݀)�쒅3]0�6�XżͲŚYG����N���`c���ڮ�_���W��s��W!�f�.K��>�r���ৱ�8�z(y\MC�9�ݷ/ Ъ��/���y]�[1�ւ�B��V�?N���=��e)(���oE��b=s���Ӌ�fK�'��g�x9g̟�{pv�mO<���xwZw(dx�K�{B��Z��~��ύ<0�l�7��;� ���n���q����|�8;٩�k�ʍ&��[K;�jJ�H͖{��y��.�dgk�RB�F�H��2��\��=շ&:|v���X��0��cB�ݤ[��`5>��#�n�g݅�l����~)��w0]q����m�5
�t�E�_�3��_O�~���k)���\�w���V��q�:���1��|�Ý�H#$r�Z)�R2ƃ/�<$����.�폥�.�lk;磳{N��*6�
ֈ��xIVD�����t[��g@B̽j�ke4N�5eL�ዼ�����3
�GL.�������,��i�f5�WT�J�
/��sM� ��W�K���ޯ?s��ŪN�1����}�	i�)�Z�GkH���g�hX��T�e�� �E9p
�\�E�A��Bv�K���tԮ�6V���y�޵��Ĳ����}Yxc�@�VD�W[O��+T롃6X�Qq�z4-�1���F�WL�<#b���,���Rh��U�l�k���Az[�9�i�S,��!\�x� �#C%d��(�0I�1'�W_L�ޅ��{��NdU���A-	xN�p����$FD��뾞�����l۾���ƨ>Z��n�ó$���P頤v1�e�x��{����gy�rnN�H����kmj�]9ї��!s{Y��tO\<�.pb*�����;"��R�讔����̻��Ͳ�m�¨�e͜�5�	���硻&e3s�ؕU�� �aIE���:Nû.y�&B.|ˢ�/zH��n,6��;.9�<���Ѡ粨o.T���J�ݺ�3f� ���к뵹�Ai���CO���FvOmv�I���1ձ�-}�E����k�nO�rҾ\�&�S}Q1��]�������pk��<ٽ7&�zQt�ǝx���A!�]����3B�N,����u؇M<P���튌̘Ƴ{nMe��5�w��9��6p��tz/����77@V���R@�$)���̬����kvH6�bS�'g�:yuc�x�P������im�#���y��؂���َgDN�!��84��DR�#N�&��v�Xu%��f��c�o
H���n����M.��S����=�.�E���t��Wk+Ƈ*ڽ5V9�ьJ�;z k�bT�2ӹ�,=�م��˚���%��+yYu�F���Wug1�|�syf�6q;6R4mV����"��:W}&��ې�w��r�V�ZDu�+�s֕#&d�q%�gHRK\���L;"����4k+�V=���z�]^u�'Z�E�L+�:�=�'m��b��i;�̗7�i��k�[[:�J�[
���*��V��qQ�%WL�U�s5�֚�˥[6�w&曼���eL��;NB�~K�/������%�QL^��$p:��1�r�Xg;��D���ֈ��qԌu.��7��p ۡ�e4�wq�[�%٘�C������8��2��V8^���i���4�EC�K��\�Pۓ%��:��LJt��V���r��}|�ƻ ��d�u�e,�uV%}�v����X�ҲR���ˇU�p`N��:/L
wP[���OQ�3H�����
���/�͇��e�t�T��9|.���� ����Ж��:��|K�x�9�y�t����
��ý{$W\"���kH'^��$�M*'Erm��z�5ޖ�UR_5�P �l�>�2��xҵ�����z��0�=���ѷ5�nܠ���sD`���$,�b���w�W
V�B��,���s�}�>�6e+�ˀʧ�e�{�/�:���L5�W��Q3��4d�c2�j��̞݀#�@�@rHg4����G��C�h4�P&K���8uC��j鍔Gf\-�x�Q�&���T����ڱ7��p�`���.��PV
�(�v���lz�d��nU���X�厳�/n�S��w_H
���V��KJˬ�oM���8�l갯�8 ����=�:�'g1�#b�6,<��	��]���ju�f�b������pJ�I�|���"�Y�^���^�I��\�W�Z�|4�Z�4#u�8r\2�^���:�گ)��d���T�EV���;���8 `ͫq]\��Qt0�L�%���l��
�r�e�.=����<�+�oE��m�n:o�l�Ⱦ�H.�}ĵS�t;�چ&�u��p٘q�Ҭ&.̘�ւD7�>J��^̵�vru�gdP,�S3�MԻ�8�Ɓ����{!�Ę����'���3�Y�/m])l[h�쌕�ܷ�����Հ( B�� @���7(��r��?/?���ع����8j�û{�o������&Q�ZL��xʝ�����%E�	Y;��s���Ğ���AL��e�����|�>*����"����wg(�(��\�I4{ݼ����s@��:H���o��(�>$e_DZO)��H��:r噢y�4�:�:I䐝����=�^]�#��.<T���I�t�:M2"q�ʍz:�}��R��U�Wr����=|g���78Z���o^:hU˼JI_(��$�3������[�	�g
#�/	��K��ox��I�<�����GԞ�{�]c���wx����K��<����'���;�Rw�B����ו�=,H�G��Q+"����է��!�֑N�r������
GQZi�]�����:��::�R�9:�Z�ݗp���-�����q{Y�/�ϯ'Q���w�y�K���(X���V|N{�ܼĂ��+�]�uuQHO\w$p��)��]N,T����(�Y��cՔ�z	�7	Idx��6���R�i���s�2/��%u��ueF��Qs)uen1�6�i����ZST�9=;�;�y�y��1����Tf��z�I��;����q�ϲB���5��:*:�8��:,�{<|L��9���Q �c�i���&�ӽ]��۽�*[�Ց��=}|�q�$:�0��+��M���p����j�}ua�r's�o��G^q�n��"$i&Y�R� ˛�Jz��i��U�E���9�6���T���H1�P�}�W]~�=>�HD�ht�l�=ɤ)����aw�l�݊y�'H��g%��P,w&�nz�\T�j+l�
L7L暅p簾M���ˢwkNm���:���
��}<+�Vϒ�9��,���I��f��2c����=��X�W��Qڼ4歬 md�!�����"�q�:�V�l�XZL�����IJ�"���vd�۩��x�tk[%����5j��q	����� m��	./	+��	⛫�/T>�
�Lom`�J��v
��
�us�m;D�M��R&���0���Ȥ��m��ːrN?e�}Rڢ4�CU]��Q���x���c�� s��\�Ɯ��3�:`o|�X���!��ޫD�yM�,�w �n��y���cwFNt�v��Ӽo����P�~H�QAƅ&���+G*E_<�Y������{��k��l��}2k�F������h�I���M���un2�ҥ�-�.1Vd��?PUu}�j���+�ӫ���kp޽�+���;P���~s*���r�y��{��wt�'vM��6��X?�`��or�8��5��O�<��F���כ�d:;O�*��h�j(J��d���=��G2�smq�EE>\<���i��¨����i�=A��VX������·_xJ{��a����>�;q4k$�x6k� ��'پ'�1�"��Lt�t��E
y�i��s�8b�Ϧ�CR��١�x��w^YS\R�ֈz�8���F�}RL�}���~���Y��ҡyG;*��q�;A\���X;(���r��pO"�Y*�6)��W�t@A(w&�zx�m	�CVҞI�6
F���D{CU�"c���YIr4	��ls��Ya��/"E�4��8�o'\��(j�&�� 9���ghB�"m��rĦosÈ��j�^	�&+�_
�N��`V:��7���;�XV�s�N�J��fX;&�	Dҫ������-��^��4
:ٲ��N�8�n�]��\��k������=
l!=�ף#gy�� R2h�T^H5��W�Q�fu��v��X*dƆ��!oW��څ:�d9i�ȥ)���va޲fh��i�e�Oa���oL�h��P��b#����BG�ɼ*��Ҍ፪��ɫe�ڻz&�~��5��O ��!���Oc �xҒ�;g��cfum�{�>/'�Ww�a�ُ�p� 9g�<;���v��7}n��si�sؖ�q����O�sl�쨓��f��k�"����5�b��~��gj�{.z(��;[�y���5⻗c��������b=˩��Svh;f+Gq'rzd����ɻ���K�,&��%%P2��n����.�@�b�ݎ���0.S�;7� �]A���=ն$�f���ݛ0!Ć��OH�:���7t�f>�n�RT�e�!�]�sm�M���$�enս��W-� ��%Eem�ۉZ5f�>v,ɇ
A�*�V=��yM�M�ӽ�Hgh�9�5��
��]t�����ص1Hkooaj��J�"v��٪�w��5�$$��� �Û!l���e�ǥ!=C3I����cf���|�d�d��3�@�g����0�ײN�`o7^�-uT�0qU5Ts+c��z`���>����:,��3��Q/��]/G�h�}�e��=U]5g۪/-��𒬃���[j�-̍�]{+��뵨LB>���J��P{�3WK5�|� h�R�$���VV���Ē��v�X��ɹ�^_�T}Q�ø�~�ğ^o8���A6������۶t=Ln�S#b������rA�}�L��� ��q(�:(R��٢���qt2.��Xn�������>�9�k�L("�4$'m�F�����w.N�Ta����bX���K��ʁJ�xA�T��v[�� �d�d��DnÅ���7O.��5��Ѕ���ls���7I�H�W���˛���G�A��9|ks.��ے�@��RQ��j��]X6�l��'%�І��7�h������ogMT�7x$�W[5�d��G�u���M6p�P��T���p���39��܀)��ϓp)2���Nx���2�Y�՝�!Ao��U�L��<]1)���=R�밎��N�дOҔW���|�sn���ۂ���$>�l���8٣I
�\���Q�f竱*�es���A]�{lf�	Q<�:��Sp��`��j��a�����ѧ=�Cyr����V��E�������~2ݜ�AF�>�7���8H��=���J�,۷���8WKnK��;v���n��"����D���C��Y�1!c�VlDZ����<3+P�ꕨ-H��X�E�>�<������2�	���9�����u�Q ������W"|H�q��v
�[�|�lx�ű��h���&��[���� ���Tm�67��^Y:I
HN�E�tR��뭴U��dNn����_^�i��I�`؄,�{���5uך�FjB$hq4F̰#6�GI3[��xM���&�'^_WK=��a&��s7=QqR��U��XM<�ߌ�83��ᇦ�ؓՅ���o�S\�g\������K��-�a�;Y�ҩ��)%[�[� ���qCkח�I]��s�jc��;HI�N��՝V�}�+(G/5�Zn����1�'c��!�o5S��9�X^*켒9&�3�\��²�]0��I֜�SsN�Y�Z�8^�I4Dwh�3u��^I�ۭ�,R�OeQ��4�}V���Y$cS���OM����k*��#n,/Rd׏2�/��E*Y��ɼ�SV�.ŭۉ�W��bMhFZph~��d6��ޔ�gI��'����d,~1w��FG_v���x ���.΢�hS�m=l��"����HMS���\+�i��}"��v	��A1�-��F���MO2n|�pk���o7�zb���T�җ�a�ca�����ْ�t�;2C?�w��7�	��r���Gt��<m`l=�~��4�p�����θ�!�K���K�m��.z�'ǖׄ$���U��#i?H�7i�N�5t�<ۋ]����C��>�'׽J��x��yNP� � �n�Usycx/�.)�k�N�Ѹ�z���\s6�OA\O˔[�Ӽƞ� c�;��z���ek�l�#���@�Ī�kw��,ծ��bF���S[��ˊlc��^���!5����h�6M��������Ļ��)�bq�z�a���n�w%s�c�b��N�&N��S/Z�[³^�f�>��=A�IH�c�^yj�E�����<;�M􆣐�G-l<+46o�n���)
�A��_)�OYYS|�c�v����J}�NqڼA�Ycidu���r��8l�k������F�"�� �v��S�Nge��B	5TT��f�hx�UY���Q�5b��q(e؁��4
:ٲ�\ӧ���'"qȷ��m'4�O#�h�p�>��D\��|}�����
i4gmW�Z�#�y�{K�۰�`�ܣ���J~�N	Kh	s�|"�Ƒ���Kܥ)J�B���*�"����ۮ��T��V��|�]�tU�#��gK����5I�7`�A8cw���w�O�Y����o����`t��l�S��H8�:VT���L"_�v��~��DcΓ��9���!�d0�A��-��}�m�ĭ�0;�j��A-��QyR��=�:uD����T�ym�gm0c�D�U෫^2h1Z�1���I*rg�yYH�h��qUb�Y{Vs0�Yx2�±�ַ�hsb2��qb�3�}�]�6aiW��8���fhDH[6�މ���st����1{	xR�0��/�8y�|�TI��`�.am���f3����XG@t�*e*7=^�[U|���֩�ܻ����	��.ddSUfe��d�>a:�O^��G*,MN�gt�f��磜�M&�߶��7�U찳��z�:o KF��;7�
�uf����놌���E�j�Z����d7_�ͣ���0�!@��am�(�s��S��9�|��v���T��[ �2�R�uQ��4s>a�Y�:���Cb(ǧԳ�	������tn�Z	�:$�˝�C:#E���)᧾�Q���~�9������2z�yҪ��F�;|���,�R'����\5�+�����|% �iT�]u���Z�2���	������7m����cw�_U�Fk��d{P�s��*����B�� �ԓM�fW�����R���**�Pr=ƨ�8qE��w�:�=1�]7�R�!�7�[Z�T"����QGc�h���mMZ�����sfP���̝FA۝լ(�n{�2���ő])h����+#;rL�� ^�lFIgM��<�oDם?U��>H��B� ���	[�׷6�#r�V3E��9����cw.��m켮͎0yU �2}�N����'%�f�V���ȯ������+;�3y<��"�JW<j���Sْ��-�+�4j���s6�kx4�^�b#o�6	;ΑW��)q����sz3��?ujڮ�hUCz�g���^Ff���*�'�+�(�4���]��NF��]YI߻�j=';����n,1��]��L��k&����-�f�N�yN����ضl�+ �ݛ��8wt:[f�@a�9�v�~\k�y�8��v7�'�5�L�73T�l��޺�8T�t6z�>���ha��FF���i+�ZY��<��Un�G&j��>m;�8�R�D��d1��h,�0n2�h��<�����p�����o��u#L�r�����6h�c0���n�/M�~@�q��ĒWƠ���ll�B��ځ��G�+s��[R���:��I�r���ȵ,�1i�a���j����0�cT6U�@��ɇ8�δ�����HS�	U&�gBs/k#�_'��o�'z� t;Je\�w��I*�42V[{I���Δ�~�T0�^�	*�m���\d�GVq��;t�<=m�ҙܸz��~���7p����~�&�F�{��y��&	#AI	��z-�b��M��T��n~�:@1O�����af�'������f�"M��7��\�h��0y��ǩȍz����=��h��	^� W��b^%;����;����̂a߯���w&�]�9���s#e� �,Ak��7fz�v`�Sw��6��\\^1��g��U�U)죵ysNdU��y�4��a�TOq��1D�í�bT?>��;΂�0��%'EKeVK.� �iӆ�qǹ�bB�bF��u���WԸ���g��X3Y�!���ؚ��1l�E�n�3�4T���߶�)��(�ǳd��QZ�Rf�ʜ׾��Vgs�_u��;}!�l� �������$�8�|�Gr"[PS��o�~�	v�E<������͉%q�ԙμږ#FG�8�.XF���&+��E7�%���' �UD)�4�<��9�a�]�����a<��;�ˀ����)
5{�����JԻ:�p��ttA�f�8z�
7���n�VZq,�����pt��M)p�`^Rqb}L/��ffsz�r����mi��'$��C��!]�L�
�wmܓ�/kBW�{Cދ��>ْ}�qѡ|����2	���y^^2����_W}@�j�킖k��~�	F�ӯvHc&-���<�p�mX����b����i��wm�Dн=j�np���<�y�sT0A�eXu���^�ǰӌ�����˩��Nq�.�I���wWG�@2�1�ڶfN���D�gf��89)Z�
�9CfN��t�!u�i�D4T�7�DOyC��6��!I���^\��%G��5Lp�q�x�^Fdo6�w�Aq���3" ���%Yc�r�fW;�\"=����H.��뾮�ܓ����7��5��X�UǼ{���jJ�Z��vd|̲g\妒v���ʘk�霙N�J�15G4W}�RG/�]�Xu��z���;\/�`m��-�ed��Rg)%����,n�Z�in6�P�r��'���7�G�y��Ћ��ܫn��Y-9�xz�'S�2�b�b��̐�����xrm���Y�8���\ã\��LU��.��3(��/7�L͚�(:B�P촦��F�l'/*`�r�/�����NuA��Rȸ�	SΚɔ�
Ɛ.�M�AO.�u59!��2���l��s�xo6��6��L��:�MH\�f�1l'ǉ9 ���D3P	����c3�q�j��I|cX�t���A���&� d��־�l 7)�a��	�X��XX'�@ѺBכ�ݐl�����'Hgb�Z�3�&���n#��ƃ��Z�4Xɛi���'@�p���6�^K�ܵ�)�tRE��6��xl�}�d�C�t��.G�C���h�G�%�0r՚Y&�SF�iԷ-wl[Ӓ�ѹZ8�!�Z� ۺ�(���T�e��:U�Ҋ���F[��FZ\�>���9�C|a�b�:�[�w"�>G�eVQ�l���)Qv�eb���M@�gz���9�����˶���hLh�tmt���S2a��\C/MJY��:Ջz[��'h]˟M���ʂg^Ҽ3�ulwZY�����wFЈtu��+�y�#��9��q�|�^n^�BŘ��us��ajt��=�$DN����n8��RU�i�3�Vn�x�}ƊїiSG��q����"�mG���l�ɯ<�z�8���1,�6��r6p�1=T���90P�gROoq�
d�5�Vl�C�*���+$ 5,
`����s��2!dN��m!�Q�9���ׯPZ8�R!c#*��{Q�|��7m���3u]�-�C���{}g����h��RL�7��_f�hE6Z��)����!�E@���}�8
��]Ȕ+#�iDuƋCq�/\�Y������q����:g���9�^r�v�{���>g�ty��<q�p4n:&�z��N�ۜN��9)u��
�W]E�==��Z�o���{�)��0�(/q���|Z�Y�����{��y�O$�x����7]B�^κ������z��ׯn��8����x�=�p{ޜ^ǾK�'HH�=Ǥ/�w��ǴB�1trISG�e۬��j��뛔��}E-'��9\/���^���M�Y�J�I�%�J'��O9�I��
,�(��u�¯%]�;�!����s�sw]�3����I�EEP�����I7xJ)�c�o8��(��P>Ğ/���.)���UP���u�)J�p��bE��Er!��y�XR����!�����)�z.�
�x��HI4G�<۽�y��ԇ;���9%��TV����y�T�*z��y�c�5�vz%�.�C�s>$��>>�(��	%Ыߣ�wx�5��7����6��
�ph��������z���*�Y�'e';�r�'����
yblnٴn�khBhQ5}r�svl�������\RD���܌��m�0��0Z�6� ���R+�]Wg2kPԶ�rE���vM��6����q��K�ݿ:�%M������xp��*d����w�ԉ��)�� e'��S�[�M܊�'S�n5��I���Po/z����b��1�z���u�n'9󟑾v�[�+΁0�g ,�/�/��zM-�҉�Ѿ���[4ǳZ8wl$,��m��5�����gc����T�5�ϋ1�ɫ�����] �d�֏v
R6)�rB�����#�(�<��^3�,�ִ&vɣ�$f׹u��i/������W]���v���X�pU���fp���!������&�"�w$$u�x�%v1ͤ�ڂL�=Qg=ؿ�Ykk��-���B�|��u*26F�+�]I���g���d�����0�X����a
p�w�t$�d��N�������NX "6ںܗ���u�ve-��h�87R#S� ,8u1� �8;r ����&��zC������,3MĞ���Ȋ�_[卮c�3	�����*=!$�������ۻC%Z/@{Sz6�s������T
�!�]�}p�F�P�(��m��ff�p���v�.*��4���g��s�V�P�h�.���C��q�@�κF�KX��,͝�Σ����A�J��UO���i� p�##��f�3N��Tl�]n4������P�<hk�H'WP=�f=�E�A�!lAC^�SN4dU������26��RQ��.W��ֶO�%D���a���_]�HU���h�!רkə]]7=]�k������]һ�]�X������i^��Sa�h0=��l�~2t97U�)W��RQ��O�����'��6���D������F} ��3�òF�\��2չ�}䎽]|�q����/{��1��ޝ�!]/؍��ä!=�yם��_O�)X)��*
�Y�@�m�����v�����u�e�\��*����TdS#�֚dS��˜w��d�h���.�ۍ�*�j�J�{I�30�3�0�8xA�<�ܥ�%�N�;Gn�-��c�^��!�NVެ���a�+�<�Yݲ��g_�51n<A\��z
�3���9e뉂.�{^���Fb�ef�i��4�x �>�c��0ZK�m��w����cPif��C�􇺽��W�Di:	D@��r�T:-ȝ0�.E�,�����ފ��D��|��jf��ׇ$-(9~@�t0�Z�sZ׾�f��sהz��+yS���g���
j��X�F�H�K(vI�u/{Uf7�^�6E�Y%�lo,�����u��U� ��
q(�M�j�8�Lܸ��1z7g̚uU���T�dR�.ZEj�w�:[�{e͑����:(�t����Qr�:�;2=!d����>�l�'n����	
��	�8o�Vs�w��%`7IK������C��)�a��|��^��[{O�xt��*�'��J��+��#6���Rp��c:Kٲe-���/�W��G���FN\�v%U�+�|��%5G�Z9��9����*t�\rT�U=���F�[�����k���5�VQ�o�;zɊ#K#V&�*G�3&�w/)m7wEֽ�.���I����q�#�y�n-si�|2�}#x���镬)�s�sN��9�q�Ƿ�p}�y>��E�W� C�m���:�d��6z�!�]������ȝ�k��}����f���
�{=N,n�r; �0+�d��XLY����9[�qnB�{O�Ht�=ԬJ&B� ���~�=>�����|�)�������=?D�B�];ѳ��f�l1�w��/r���^*߻r���b��١�
�iW�	���?z��Ȩ�̮�Z��<պA�Z��T3��b�����w����O��$��7��\T�j��~���VEF<��L����)�m^��?Ч��g�tj�Z��ujho��C�\�&��S�Oa��o�
Mw�c�m�*�jxamwa2�&k38QӨ"ٔ�E���,�S���v�����C���&��E}Ⱦo�4����T)T���SNg�lͪ;W%{�X��΀gC{���&++�gg�AB���U{WS髎G�02l�<�:mg\������.)�e��')<���Z�C�J��:L��N��%�+���9�m��v�<3�m-�I�Ne��v⫠�n�Gq�+&�����/�=�u��T�YÌ���[&o;��{��}"G��	�F}΂��q)�l�j��/�V"[յ�^����}[��K��S��锕����g�U���l���������)7��s#Y�
dV����2�m<f�+N[��l��Jp�`Oe�:Rq���}n��o������.W�Q�}�Gp��~{o:ѵ�K�+� �ǐ7��(���de��l0���t�#�4ÿ<:���L[����qf�ң�j���X^}�v|��6õ�=X%
���c����v�V�H8�Έ=�	�h�o%�&���.�k�O�b���>�Q�϶���Gp�����k{Crwz�+Ga��r��1�F��t*��V�4Բ�����t����� �>ّ�H�/�/��c�a�b{�/K+�u�E�0��CV�9���gc?~�ѿ�Ǫ5���s��c*��vg��\���J�={}D���]Ld>�5W4714��|+C��p���iu蒥;�	/n��7e�N��-�+��p��o��cY,t���;zਦ�՛d:��0U������s@��S�Ö.h���"��a��6仛���<�� �j֏�Jv)���;�+��M�=����j���騻C��WDD��˨��y�YJF�9��qc�o\�c3BkǨi���{����;�2�V�\�HOZx�4
:�Xu=K$筣�L�1�x��M�[�t���h@b;c���JԪ26w�Y�)�;j�ؘ�Ǧ2�2�p����:s�����|�A�mG[�����}��^Ȥ�׹�G%�^��B�Ї_�OXn�V6L]Ɵ�޾���Tâ�ۍñ��"de�t���\���l�kp�٧�Y�ЀJ�iTn:���s��2� >�ۙ�]�o;g�k���5�:Z1��s�2R�s�5�=$��=�[1��-�B���3��{hX���Z�s�Xy>� ��t����ԔP�K���Zٝ��}�ݝ4ڡ�Z���"���]��7�a��2��M�P�35�^}֒�+�}_�
�*�������v?d|E��&�J���* ��@Q�ui�xҷ��|�n�̽q�wX�Vr�.P��nRd�ڒ���<�,"<0>�xʻqk�6�<ے�<����ur^8�7A�x��t\�nV-ϓ��V�avv�+�w��s��
���,�����/���}�����@`��n6uW��&� Ҕ�^�O�?8�~���=D�=qe�9W@(`�<�fǸo@3��#p�.W&m|�枪��Q�o����{�ܪ��� ��0sa�}>�����E�n��O7OG<V�TH���>8O�� S�TiOPe��h�!���
���NMfs!Zq��.�٭�Y�#Lp�᧏>�y�X��{/j,sX�/閹u���֐��<rm�GFi��#I�ADG�k�嶋Դ����z���5�m{٧��1��P�h��]U��Z�4 kԖ�y=(�Q�O{���z��|��l
@��<�S��V#^�����0�}B���Uh����{b8Vމ'��kI�Q.g ��A���"��l�=U��a�N�祔,�sŝ��Ir7+�ě0v��w2zi暐<���Pݪ�Y��F�����=��y*�:
5��0$�z2d����F9] ���KGl�ʣ�>.����W�n�̬ʀ�:�%�x6F`[n�u*	n^��K�e`դ=ج7|�f5���5B{�ڗ��V�I�]^`t�[�2s�ع�[V�	�[���#`�$R\�4�K=�n��3�Uev���;�K�OV���	�cG���cٰ���t���&R�-������<AѦ�o1���t����C�ӲGOa�Gǫ�*�+��7ݜ��W�Y6]�zM���8a/�����D�g��v�Uky��UԴ�7}кo:Zɶ��'8�:]J���k��dy�oPm�*�f�����[B�5�����l�� i�Q�pLz$�[�����{q���8`Qi�k������y��2\�r�Wƕ �d�:���W(��t�c��-�*��wk:�4u���:�R���r�E��l��f��9m�7]ug^a"_Gb$r��hd��׍�+W� �՜b�6C�uYȹn��$s�	�T����i�Q�x�����Y~[�z��O�˰�]E�DgB��X,��}������usv�LQ�ޑ�zMoG��)6��7�6�@}�)W����^엩y�WX��/�Z�8i�:z�u��xII.v�kB�Z9��x����|V��e�W�����h�T�&.Ѩev-�H��f&��[�;r�X���x���S/l	?u~��^��̈́B�J[W]y���B��v��sҋ�4���;��2M�!H�i��=��(wB	@{�0�HHfvK�+j�8gH�����N�%�u>WfR�i�婹�;@!\���M�>�f+0k��n������}PU�#&ו+
Nϳj�TӘ(�Z��0�wwwT\�7`Z��?!=xE�::
}�W�B?�A��Էԁ��[��7���ߪA�	��܆d:S�"6���)+�%�F`�m>7�O;�gQ��?_Ht�i��������F2�m?��w�:�ץ�Fd���~og�����?G������:�dj��L�z)�X�M���{��f�R�C>�4����}=���{�g��hBr�Vq���0�'0���qGjϦ �6���&}���'�;�m_P6��Z/���vvP�&%�����t�����V�<C/�3J��Ge�+ʱ�xh���΂%J��߭�*i��Z�� \��wI![w�p�-罕Έ|��!��onJ�.���_D��ü.H���n_�o=RQ]Z:�g�2�J?l��E�Q�R��v��<4�.2����}�O�ݯ��yx0��j�ٝ]����o���}O��Upv�r��,^�3�I�&w��O��Gr1#rF�Rb�[��r�鵒6�������5�p3Ϛ�o�l��ϣ��B0�frBɽ/�/��~ş��N� M��}-)߼b���λ���5���vm�Y��Kz��O^r�l�3݀�m��]48�$$j���nh�e���~��G�̬B%������]����t�gq⬄�x�e)ا NK����b�T�pͺ1�������S�7"�.Hu�w��Eiͥ�Q7�S�G�1���GKPWB�P23)AԈS�'��W��
iGL�C�L��8�����mӽ-���й�٠�!U���G�V�ٰ�X8kr]w�Tǳvz�{/)�%�F��N��l���T�^��Q�U ��U�I~{L�oY&���i����ik|Dy���Z�n�'f�6t���.D [>4i�b�[��J��]�L�$�T�{�/;��(Wmn�I���f�k�������V+i\F�:�I�H�����Y�G�q�H���۷���!���l����s6[ۗ'ڢ]R���7C�:>ۅoLT��Y��l���ں�!ׅ�H38��2X��&�Î]lC&��aJ�D�*��d���ײ}��..�}P���ԓ�����v���v٪v�M�¡7So�2]XS1��&α`A�w���ƅ(������3��;Q������ݽ�ډ��n���$T��k��������9��dP;��$���P��E��T��f݄���Ė��r+����H��'&XR���v���y=�Q�U��4�����m	\��$��#O2��V�D��I�>X6X�8wJcE؏���ԥ��w���%�V܏Uͩ�� Y#\�-yturvB�dE\�=:�-O�0R�E�7x��cr?����G�:-��]gJch�hz9u�'m�F�����
Kz�
&G��ɗ&*+|�]2����;�N�O�D�צѬ����6��UCp%2uĮ*I��p&ڼ�uё�V.�C��8s8�`�]�Wy����xs�v�՚��!(�����#pf
�}`>	(�xt|mĕ���Vd*�8�c��	<������%�_�I�:�ñ�2�9�GGU�\
V���m�Y7�Tm��<�6�J�{�o��oO,�<��i��Y���uxM�UE���5�m%jӫ��P�X�f=�-��C�bU�b��kIX{�������AҼ�o�B�l��V��d�w7����yp�SҤJ�.t�n/�.ẚ�q<\�2E�S�}n#���U�.�ن��ܳo�[�Ӕ�ͺa6��}��ә�#Ԯ�eG�X�#���8��E�S�s,%r��qb圪>�{�AX[�!�J�blC��ڈ��t��zݹ`vn���uN��+f3�՚�	D�uj��f��d}�M�.�kRn�76w=�Pc޻4�Nj��C,^^VVbMξ�X����,j�W8��z7�J�|a�ot�:��z2H/���gl�����$zk(���gI�p@�J/�3v��7�|��"����7�;2��	L�'��aeN�]�a짖�\�:���T49F��8�tj�v��jA�H��J�8	5�Z�!���{�!k)V.�f�!���8�2S�l�5*��F���_RH �`�Ck�g)�Ŝ��h�ZI��8Ou�� �!]0���Ѭ��7a�Ek�1y��Ga�s��ݜe��K�w*a�d��ubŹ�����꾸q.	�WK���[#Ӛ4G�p<�QKOO,�kf�kᅻ)ј��ĳ�3���]�/f�b5i�w�s���P�a};M���.�ݜ�gK2��J�F�@R!B�|��G�u1�wc�;�v\���S(��:ev�7�����WY&������y�!�Y\��G	L(�Z�B�8U˔N��|�7��|�>u��x7�q�\�Zn�2 ��$]�<��m㼺㓄�: ��"��xP.뛂t쪌�U��<v�|�<�J�DM�\��udZ�$��M�L�0=IΓI�
mΐD�0O�ᅯ�M��N^	�,�i�h���n��w*x�:]Κlל[)�RI;u4�����$�|+rI9�!&�yL��,���+[��	��紙CǞd\=d{�x�U&j�����t�s��4�RO����<��B�ny��蕈#�=��c]*uI*�d��gry���D�*.'l�>�(�>$%I>{��l��me��n:=#\<]5���+ y��)�/������0�j�wM.��zl˵��Ԅ�8i{~�Ù+�9,���߹��?I�*�j����p Q`�t��sz^�[��CEĉ�y�r���z�����4�J�:�C^z}�uux������SMҫY��A���pI�nOI#��q��+RQ@q����xZ���+7�E��f�Ek��j.EN�����ǟ��̮���S W-~������q8(�v�Dr�;xGy;��v�ƸC��\dFΧ��&�96���.��n�>��>+�W��f�}ғ�Cz�������vj�op>^N�������x5f"�V�q�{����Pn�����w�ɚ�l���>J�ͩR����ϯ��c����d|����2�i9��f�!�/Zo]��lB;��8h�Ϝ@�I+��txY�>�'�i�<�㢌�1��.�Ok���v���m	�c��ϵd��Di<7���GSg;�} J�9���1�wne)Nx7\�PP]�㩮f��5,�?V�bv���[�#�:__k���
�:��f{PN��[����������F����kyM�IJ7{r�%��4l���<[O�u��bih2��q�d�r�ywss�䢽q��lЏ�|��œ5uB�d�H8�`�,��3�Osf1#{�A������Ch�\z�MU��}y�!;����4�����ï�v� ړ@�֐z=SSNdag�
�9���DĶp��DR�:C��ZJI�\����2j��ZFv���{�ҭ��W����~�|��k�-D���vu�D��Q+�x�x=ڑ�n��.��,��s�7�3{��r��q�rE��=�D
��f�'�$�t���nl��=������9�U�\1��*���8d+��$t��*�'�WJU�Wh�l�}��j/{��9V_6�vz@a��\��_��(����J�s��ɨ�5E.��z��t7+{�q�u�v6Pa�Y!�oPْ�L̼�˱5�����Y��'NV��^�J��!]l�0y�a ��a�;���x�%{6��f�Kh�#E�\]�Z�]�16v��F�����jh=f���^�E�F�n����'�%��tu��Mfe>B��Ռ���RٖHL���͗K�^�n�E������-Fی:.�XӅ:y�vN�a}�5�r��4nV#�W'N��8�R�(�]C�Ƙ�t�t�Uƞ��ۓz/���G 㕸7b��P:��˧+ˢ��pv����ڜqpŎF���vB�Q�CX�V��쐕�d��G"}i t]��f�������ó���x���r�5�F�/ޏ?p��ȫ�w���ta�E�t���B��G����/���� !f�O�s�X0�q�̋X�a9yd��:�H��ܚ}{K�^��g��  �=̮��z�]S7op:��fb�*@�)m�:�^Y�)v4��R.i�첊�"\d�77�|�c�WF� �1��<(�����(+��%^X�(���U�Wf��9����t�m�^�����6���!��d����+�t�0����N���B
���e�����6���i��8��K�2D:S�"��)"����L�<$6n��75[4��U�ٙ��A�������$��Z`���^kj�K=*��,P�*��Go�"WH��ַ�y�#��K`���30n�~�r�o^�㚆�)n�X{�w)��� �aX�镼i�͢C�� ��%��9�/JLN.N��o+2�I�d�ũ�ۉ-�K������:�u��E�+��� �-|�{L���n�U�����qؗEX�!f�����An��w��67�g�B�)/��^F�VQ2��>F^����"��^��gq���7���f���k�v��(�Kϸ�ɵ|i�vw^���ʽ	�8��ZX�H��~�_��S%�ߤʟ?u���[IS
��w{��N����}�<�$�'��2�C������T��C���Ն>Ꚙ��*����3��Xk��KcgǨ@���ϣ��F }�99�[�_O@j��R�}Tm������6�5Ż$'E��Pg�gC�`�e'�WA⦦ED�B�s0�OW�s-v��Y����A �V��Jv)�G����k�m��ȅ
 i���S��?o��i�g=]�Ǩ�J%�VR��r�����7�l��+7,e'*��(�k���$���d���hR�}J%R��B�A�\.�7n~���k�7UR���Vz�(��n�!yԦNw7��Gi��7V1���L�B�%Xy˕�0��ft��^�»?�#�ye��x|WL=�\�:mC�#��e��S3j��6�~��z��	�>&ѯq���<ip��w�\PL��#ck�g�S�KQ�Z�FF� �G���Y[��UU�������S���j��:�*����"�V���ֽ�k�ʴK�^��0�:�jۍ(��]g�+V:�V� bb*��P�b��:�o�z�;��=-�]�����hqTi"���}r���.���C��"����=��밎�8�	Obx�=��θƻ��ei����[(/1�=f�kѨ�
�dl��;!OZx�(�4�XO�=k[,?\Y�� �3<�yve��_E(U͐�g�;�9g�fWW�nz�b��Z�֒�<�d=�=�T2N�<��H���`�mpFl0\ˋ�j�h�9u=�x�S�kz�S��"�w�ޘ+<�FN���#6��=1z���#;���6��Ǖ��l~}��J��@���Э2Vf�I�#c����D�u�����^�N㣯,e��E3'f&E��Ŝ;�X�BޫTk���h��6Sڈ��S�;Q��7DVc}d�-��r;6�����Ki��t2��r�����~��=:�t���:�wzw�B꫻{d�e�욗�si��nS��Jo��G���6S�Tm)A�{���1�ca����*mĉv~��\�����6sLp��4ϸ�ǎ�'*�59�/36�3H �^�Y�gBa㔾գc4��4�
 x�,]����/;�uv��}?~���u#Cz(�{�b&���ũ��@�<E*n�1���V_	#�;� VI�N���q`��>I��V�j1C��'�rh�sF�����A6��]� �SÚ�p���2"Le;mhg`�,4DK^~�Ͷ�����&y�Y\��lɨ:��;��/^�h�chF������1�5��
4prF��v}�R6�T
JC�5A����Yb��Ʀ�����T�[��Q!d:"��d���`�03a~�I+�h}�I��U�����
h��.;q!'5Z-ڋ|�f�C6�[�yb�A!�G*�҃�
��jn�nۨgH�6�lu��ao�	�&*�B��ʵ\���ڽmR[D�<&���]v�Y��c�]f��X�i\�#���:���SS*35��@�9#�wt���5�<9��w�ЧZ����rV�V2]�Gp�1)Ŕ�])'W�M�9���;���}�ݯ}�!ґ��d���ЁW�?��d��M���@���v�������9j���4i"����t����5��dy�o9.��;���w}���3}�T7�*Y�f�����F�v���];���m�����tF�=C�Ҡ�d�ռ{�\��Mۧi����v�5���)���ă��lz�+���GR4t��s�`M[ӽ.�e��z7B�4��A6Y��%��<+W�$2G2��!�'��V�tw`�'c�A�V�}��:,�xTj2��n�ji��F��ޥR�m!�w?F�p�D/r����/�|�1Y������i�ޝu�pɚ���H-ؼ�#��VA�M>���o���,V҆?w�<�����݅��cy��,�g'ջc���ggP5��������][�Pu�3���E�S���w*nXڕc:�U��	��GWU:��W�Z�aι(�Z�g�J��A\�ͽ-�8/�Y��U㫔Z���$��r����<��?�OҶ��)WfR�i��74�0�z=�7-��g�j��:b�a�qCr<��
]�Ph��g���,R�Oc]�E3C˝�[�Ps�����u"�����+jp��"o��t�]:^��t�D֊�]���t*Q�i��e�f����Dd�.�#����J~y��||����vF��h���x���u#�8B�����w�OH��ܷ���h���r3���(��y2l�CW�y�֏�W��8touw~U�:jq��Bl䤫�rI��Ek��W�Q+��0��l>�����{�g���mlЊ��N�C"9V��v��QzX_x�ɵ��"��[^9Ǭ�Yw���},�g8�P-�ٝ]����%��52�2��YT)��nף��*,������d8ÌF}�77:V�+Z)�O���|����&��_^�c��cR�6��C��.r���w�~u�}/F[Ź[F���fG��g�P� c�lG��#��c�I�f�~�WCpI��{N模��Q�)X���]յ|�ö�<Zt��c*Eؠ�0��G#˧Y�7{uѬ<�$7z/��$9Cy��v����Qh��=C�6��m�F��dd��1�,x�w�4f�� �����ﺀo�O��1�D����d;�>��E����J�:;��&(�䞡��/�F�#I4�G`�>ا�Z+d'ӛ��Ƌ$N@u�W��(�s�����x��"^e)��/���U�;Kk��VB@d��ȏh.�H�tvnE����d�DU�3�D�U�IL��&a�z%����t�e�PW��dfQ�JԪ26w�YҚE<��73v�^�KءH��Ǫ�术P��p��!�ڮ�h�V��ȓ#Ka�w��%��\e)J�]3�r5[��pq9�:�C�ַt�?Gn:�,�n��B;	����x&�F�*����p��&�{��i[.��GV��p@}�6�)�/L���h�	����Pd\��c�N�J���L�؞aA� !�H�E���Rm T�
�|!�#��r�m���������`w�>u\�����;;+v
�ӏ.K�X�wk�C�M�t���ڛ��`C�+]��bk���.`�O�X/��Kn�����l䢡E���q��w���No���Z�l�g�Od�Zx�(�q���}[��;%���j�8�v�6�2�-�[�ǜ��]�7=أ}\����Vw�1�2k����ܮ� �)]��?���Ͱ�O�D.2"�U�F�d0,��}�����+2�;z�6T�
�d��3�fψm��G��n�|z�O�u�H0��kz�9]����=�Bt��6GPn�N�aKrn��l��"���GY��f��(�y��W&�8�I�3��oM���Z7�7�H�,G
j�jH���f|_D{ta��|]�.rLc�m�����l�i� �g(���S�Z7�o,��t+���ylfSl�N�l1�{�Y���9m�=9��B��F�j�xp�5��*��D��_Tb��.�I�DTm̈aC�H&<�S��a�<;�Ó����vn��`0EEm<�_s�z�ae Vk��b�( ������L��Ƀ �`&����L��8s�G&�˜m��{�޹����`.Cnɀ28ز���m�gm�8 � V�*�CU�6; �9��g!�&M��3�V@ �U�U�U�U�   �U`�Umjl�0�U�U�U�U�  �U`�@1X0X1UZ���   �U`�U`�U`�U`�U`�U`�U`�U`�Umk��� 0 VVUVEVUVDVE�e�4"����iA������P'˻���`6�g*��$���K�nׁ��O_Ë�^�~T��Ʊ����������1�I�5�K������m߯&����|�A?��y ""�F��(���ֽ������7��A�I�/�vg<O��N��`(��b{���~�w��[��E�!W�_�.M�Z�c� a��w@�(��Ĉ� �};�h, �81��C�0`��!�m�
 @`�U�  �� *�"
����44
*�X ��EEJ �� T@��$��c`�D�Ζ���D WuP   �3��x���Ƿ�&!P6��*֠yX�3ħ���o� ������0�5�ᨆZ���kC�n�?�F�w0?�L4~�;�r9TW�Ɇ;�a <S����q&�lUEEw������;�Y�i���XA��6�2�j[� �+ ��ӗ�,��!�@��*@���x���d������2@�%�02AEEd�[b�X�.�&=h(����;�C�jq�s����g��so�5�=|�g4Ν����� �?�{�RלAEEe�:�=�b
*+���e��4,!�Bk�C�	A�����s�4Ԑ�Y�e����B&�_�9����t� ˆ�hЇ ��\祃,�f���.�k�b;~�aԼD^�����b�� DE|���>���eXs���B��� ��b��L���x� ,� � ���fO� Đ��wޒ��(D�R6b�f�J�U(�-$kRP*�������6ʥ�-2��TA����"J%6�	P�I(4L6���}������յkIa���l�clZ��M��CU��U���v6M[��RƖ��̪�+V-��aff��SYUDЦ��5SF��f�jDڳS,���m5�b���*,�3Zn۶���jő�b&k2�fҪ�eTU�f�cV�3T5�U���m����Hm%�[KR5�Y�ݚR+��3|  ��ػwکg<�os�۞ܼ^t���ۮͽ����u���JWm�^����� ���zz���N��[wu�u͝��݅=:�\t��]����M�M�ҦZY��5m���  �>�C��Q�ء���<S�:4(_|:(S�CB����{�xQ���P�lC{o�>���z
���)Ҏ�����=t�9ڧm�K{�\��ۗA����w��ۛץKa)�m%�F����j(��  o[ ��m����7u���x�^�6��.��Q���������AEV�ܫ���[�m;l�jP���^ٯy�gZ���mԽ����6o3t����A��yeiX�Ylͫ5����Ͳ��   8x:J�K�����ދ�����t����O]�h��w��ts�����릂�ł�4�w�t=:�/{��y�޺u<�j�*�^x�*�����d�Yf�	�d�4�X|   �>���@M4V��j;��Uv���tAda�mh1� �Qg7m�A#�v�]h����a�5�uJ��5��[km,Z�������   ����_mtv�䃶���t�Wuc�*um]������׷8��wkcp&+��]3��
WZ��:�@Q��C���f�ڶmV�2��   =�X�mc#z�]i�]�S�v�Fnm8�֩���j�YA݂��]c}Σ�lj[ښ�h n�  ӣq힩BMaiR����:%u�   ]׀ C�� �p �`@ޯM�  զ� �` ���
� �r�`�M���  ;MKR��5��5bv�t�	��  ���  5�[^�5����p4S�  �u�x /`'��h��O��1X(h ��@�z��  �ֶ����fH�5�Zh5SS�  k��� =�.  WN`�:�p����t=�^u s��= �^n  ��t���[��� => �~@e)J� �����hdi���d�R�4y@ �!��*   "{P*���@	2�	�T� h3S�����?����/
8�=N�?��v:kw�gb�mZ�6ԽQ蒓�|�5~=�7���������?/���6��ll�ll��ll����1�q�ll~���B~���t�?Ρ5����Mٱ�v����Y�vЩ.����3E�k
�t�IB�7N&ջ������XJm	YX�	�K��E�Q����^���B���B�8��b�kEefc�Ջؙ��6�;?^��)X��h���D�Aᵎ���֫��F� �*-#溺�#l��Ih��ɴ)<I���K]��vA�Z��/F� *�o�lA�fLV7(��Jӥ�����A���D�F6���ԇc��$��7���׽�*�MY%#�qE*Xb���V!�O$95h���7�j�����4ȴ��!��+F�I����ܧ6�۔^�o��*�0����N�]nfS �-g�h��h�
j�1�Y��j�f��Lף�/��j8T -Mm`!�B[wS`rd�4��#APX��El�0Gz,��pbӇ�%t$u�9��Iۊ���K.L��ݡE�n^�ť�ǉ�ݩPn��N�F�)
R����*M���kQ�U$*�k%��F�%�E�9I**M�0l5�g-�!YXql���^ѩ𫉻\��Q�e+mq�={J�'H�A=��YV��f�D��n�H��5*㲅@ ��v9ETj��J�����ܨ	l�Z�Ǫ8�6�G%͉*�k���4鹘J�!N�0�� 6 ��ɢt�]K*��!Ų��%�z�9�8��m����@�2[Ֆv���,Rfx�WC	[Bi,���������V�����H�3+7i�,6hn	���0R��%�jhwS^�2Dh�۰ TV
�bS݆�9st�eJ�`g! =G&�u�J
��)���������se��:�d���@S��T�lkL���gMmn�.x�ܢ�EG"���^��- l�2���7Ru�)PZ��Sv`�m��F���'���.��'w��;�t1�h��"l��^���Ʃ���� ��؛x��c3t
�f2��KSA�̥F-7k^��N��cou/�Z�ӇF,�&6J1Y%L״�B&!�h<�h��*��l�e��=���K4��Mj�'�R�P*�Z.7O>�i�į��X���c)�5�����X�F�n^��0 6�õW⎙iM泵��j�m��kV�;�6�'ɔ:�[vpbDG��;W�N��Kʕ��ϱ�w�#�ma%�-�3�Vf�&��Jo�E L3%�x[q�B�H��tV�j���Z2�B&0�]q1���Vp�i/ >V�U��0��I���t��:��c�S/�su8@�0�	"�/�&�6��s#4��O?YZ)�֖L�o.va'.�i��}(�Ot�����]WNn2�݅�o*ᮦV�f�ôE
�Y�9�0	0IXCAM��ѥ���T'� dL���CӔwt�oil��K�Jkc�B��V�8h����]�Ь	��t%��v�T�L'j�EX����ͬ7C)cSq�7(5�E'N�z�����U��R���3��J�D�x�m�����%l	���M����s[���Rʼ����ԥ��lX�Z02l<(�VC����[DJ�%+"�I�*�۰��D bJ��%އ��Y�w����dЌ`sE��y��n��+�t˪Z%f��Jo�*��/�h��LI�[���0]��r�˸��HAP���An�(���"^�G�4<��/UmCHm�Bw��*RGN�n3���:5�rEa���9L�7lF\�j�m�:]����Gi:̤~�!�1�Xn�H��u�wZ���o^⼉�lda)y�l�mވ��Tv
P ��J#���J�%��B�Kxf:�K@�t��Koݼn�ڀB�J^ٷ[2�̺@�����PX�L^�z���Z�,-;,b�:%Y��oaaѥ����mX�OFހIb�q��ԭ�w��a^;�ƍ�JkZ�̍����.��u%{���η&n�&����k�7�3�;mٍX�������kh4�ڿ�%��j7cm���@��N��׹�G������S#����A���"�74cd�x��u�W�^8��R���K�D$-��
w#-$�M�+!(��E��7�N�b��L�z۹���Ö4�nA[t֑��nlB�CE#�J�w�Vj�[zsdz�,��`4��,�*�Kdhk+6ay�ܠ�%��8N��='�7@7lP��X`m��˴�7V�3Y��؛�Rv��5�u �[z�0 �����ڒ���>����Z�-Z�oaD4,
�]ی�i�Ht��$�ԯ4��7V�t`�(�wZmӦ�7t�ܡOjX��{� ��2�^�@��W))X�x�h:�NdT�����%���l�O-�?2��P.�-�d[Ů�"YAa-��t7p� Tɰ#lȁ;�������,��r�׎'�f��UM�"�B��0iF����+�����y\���-a.K)}b��)�d����5;D(�aSEX��Z�V� Ood��I��j�8�h��l��)�i	������z5mD��7ҬUֱJ+R�(�;���us\H�R�^f�F�XјX҅^�b-���`�:/Z����g"�������N�^�И����!%�:�ڙ0��ԫrnǈ��9c*��y1v��:�B���]ô��H?i������@8N��k�3��q�G^�V1�z�	���[i�7Zӛ*�?B[�2P��E�tNU�?C� t<��*%qnTz��9+۷��]]�)E��B�)�{F�{�w(W8*�h��uրG��|�1C��PvㅨiJ���]����B��,ǵ!�W��[��.�6�7V2�
��z��t��e��7(Tk�b���-�r��v�"c�C#xD��^��j��Ts6�x5m�A�H�M�s��� RҎ����i9����'T�˽��OZ�
��c�.�	WQJ�h�v�A���jc����j��rٿ��;WJ�
ak�2R�nR۸�X52(z�v��Y��iŘ���Gf5N��M
GIێ�Vj��L�X�͌����m��] 6*Rڡ��}4^�40䲦�v��C/vku&5WI
V2��9��Y�ۓ[�-��h�Kv-8v��m��^E��F���f�E��;n�0SU-�J��C���1ޗCL�7��'����,���C]� ��
�"�ZN�Rj�����A��--��ꧻ�k�[.�*Y+F޶�z�z���F�]�.����4��Y=�5ۄ�x݂���s��,��q��dk�V�қ�m�O6"Z.�ʹ��[-��6tև2:ze�7�A���o۽:ӄm���ݲ�+�E�����5�U�ڨi�1`��4��
@��*"�ї����.�mG����V1$��+f����!�L�4馵lZ�"��'�nd��4]�^���N�@��fj���Z$^"�fe��TV-t&R��EeCv"8 ^51m����Ns!LVӅ��%c�т�LM4�6	HJ ��%-�f�_7��cY25w�>#n���xj�`@���(��N��6+on����"���v�Z�@ �A:���{��9��kl����N�B�/�Y�c/S"�fͺV��y�������`��{t	[�y������P��2�6E�d5�#�$��|b��AYw0PAhĬ�Ĭ�t�#lF�lL�NEE�LhU*-�Fp\���*x4EnD���e[J��C&�U�<.�;�}wՐT��!�GZl�2��Ch���!lޒ鈀�ŀ-�B�ߤ��6�%��ԫVńR��V�-��8����+BH�R�!B��Cb7/5�l�$�:����ǿK�MQ�O.ي*��Ϡ����2� �@��zn��%�חz n��y����*��f����L�u�qVŁf���_�jJ����x��6�2R��[#-�X�"pf I[���Ņ�2
�ޫ��� �hސ���F^'-Թ/�i �#���]+{�fd��W�#B|Q �VÔo1�����A�fm��ͶJ�m@Ԫ�Hh�Ww2P��mEM�7H�:�۬��� V%n���v�u���Jlrca���ʒ�ꙡ�50۰U�tJR�-�/ �S�X�x�x�;@�k[J�l4ť�\2����/�Ba�R[�d�.���m�IMtD���v�	�[�i�[ ��W�35�Q[M&L�)��G72�rH�nΰAđ`�)�����Z!ݭ��a�����R��ǊJ�^�/pw��:�mgm�Q#䉶wv�Wh4,*oV�F�@���u��^V��F��洕Cb�A=T�{%�pY;�{0�BhM����d
�ڭ�*{f0�ߖn��c�R��Or;[Eܨ�e@�ͩP�2:�	�D�Z�n3�˱w-Q���5vm��$�j��.��i� &|��SkQ�W.p�H[4�ٹ@Sg� �:cX�t���y%'���6\�m6�,��1f��M���54�f���3��QlN�وD���jT]i�OB�%����G0��^���bMy�YBk	�p<۔v�F�-��J!V����r�R;��+vM�e�&�YM�5�Kpbw{�%�j,�fUaN°�"Bk�KvQ#57��O�:'O�j33u�;��ie���cl�����'h�����Úla!���P�8��*�R"�ݫ����)���`��8����������(�XJ�P.�v-�^�ѓq}v����aqq3*U��xU���$7OV��p^�`u���-�VkY��ۓT; �Z�*�4E�5�V7��V����Ņ���i�%'Ae�r۶�Tş���u���4�5mfJZf+�đ��+Y��B�ĀD����wb0�R'@��eś�-oQ��ڼj�.�oVɶX�ŧ�3"�Z�8T���iǔ��9VJ�.ں��O+����t�.у��xvi+P�E��wN�y��fm�-��Ы.�d�%�Iɫk1K���u`�
�$uI��HG��o4s*�̵u��nҼnh.V�9@��khS����K�sj)��Ms0�Fe[���+b�e$f�t��/��Cw����S�+
!���SLfm��۵!�T@bC)
��/4}u������s~�ɒme�Ġ-H��`��PE饡��l��d� �%a��ۚ[�R�^���Nx���X�I�ͽ`:��EGi޹u��9�7t0[�j�^����d^L$TحV4N~gwk1���j��Z���̖�J��aǻtS�-1�@:��69$`%3K���6���0����'�Z�n���[���U��e�Si	*�+v��͹J�َ�P$@�عG1�՜����Dcl͍ܲ�d�)m�����A@�M��4l��l�P
o	@�P����;�^��6H�I�k����&�ľl��z+t="�ƳK�h�t�׆�9k(�i��j]�K��@��:���≡�:������K�:��:���1���b3,=��e�n*Ҩ�f-`6>�v՛4�@�d��و�+&��q:g�U�j����m*�ZZ�ie-�J�B޶Q�1j*������#V3&�I�If�ƥn"���
Q!�b�B�$ҫ�Y��������S{-S��w.��K�F�nj�N���Hf�T�0]��l���-m;'v�H��A�Cri�����sCMƳ!ǀDU�e����x�{l��%fT������P3���M���ƐWm��"���ʡv)E�����s.�IY%���I���pe6�����V���&�aOI�+2�S��W��m<%�4֫#E5Q05̇U�0�)��4�P��a�D�&cٚD�����tƒ5��A��i\�U(�``�`q�A<r;�^��ۚ�%y��7PPс���+/��)A,����3����q^C���-azx�*�]���i[���� �S���	T�r�RņB��sB*�7���Ŋ7����n�|�M^�q�X�z��I�B]���kX(�ˍZv/%å}J��b)��ZkUk���%��`{i��\ڱt4g+۝a�
uɘ4��Q��<+%\�h��T0��÷4��׹��4ۀ�3H��34k;SC��-*���J˹s.�)������v�1F��ha�F�l�g9���1�A�<fm��~6����,�ѻ{��i��D��X�(Sïv��4ȍH9�jA:`�� �\����̽���L�bC���Mԑ$��
ͅ�!0-"
 �x�v1�K7�v�!X�ۣD�Ccݥ&���4f �6��ϭ��>@+DGr�W�nn�F�N�Zk]�S��0?��ʹ6�m^���D���8���bF�6��2!�E=a��;�@�7��`r)��Tr��W��״\�
�3 �M��^ӂ�H����+ma�?ZT����F��FL���`��v�$3�*(v�7v^;�]�6ŀ�j%�N��ar&dhm^]kZ��lU�4��J��Rk`MM�X�&n,�r��a������m[.nr�գdP|�w�TN�TБ�{G!yv����m����,n����x�<�]�8��YemX��S���/7	�ۚ)�7�>GU�m��#J=_�Qjj�!����R�Y*�4���f�R��%	R��J�`1���
;�;ń�l�sZN�4UÚ�ڙeFZ�&��i�8��%[�5�:cr�3/Nc����Jb� 
���Yf�r��v˲����iAA0-�Gk%Ț���|�U��{{t,l1��&1u�n���Kn�k�7��z�-E֦Y�q%��/	S��`c�&j:;(To%��t5ʄc՝Ŧ���u�fDhnp������:��#�մ�ۂ�!O��g9ڻ�:�K`�<�ۂ�h��gD�l�{�V������i��=���u��)��o
���܂MD�j�e#x�_!h����Ɩi7�s��e�Է$�oz�pݔ���Q�O+R2��t:�, H�V�Ch]A��Z�ؗ�����۝��u�B�	Y�N�H��[j�+\�o.��������9�Հ1�ĵE��s_/�cV�)��͙t�a�cR����ᮔ㤯7t��S�θ�j�@��n� ��3�	�LaI�s�����V¯3��;���Kh��H�Vz˃���#+p]d1��oQݮ�I���� �i㣜QMW[�9�Y7xA׹xb�K;6�sG9�H����KU�:6���Ʊ���93l�i�X%Ҩ$���FT�%��2�XI=�ƫu�>]����������&p9��j-ĩn�Ⱥ ʷ�RTć9{k�8���C%>yit�: �tgF�Ö��B��s:ܰ�h8�8�.�:��s"s@��e��{
��%�f�54ҭ��ܫ��Q{�u4��km��5�@�W{YCeLm��H��n,
�
ʔH�T�Ŕ4��kwc"fd�ug�2�B��ꗩm�U��,�q�Ot�`ˈ�;�h���,͕��Xp��]pg��=�n-�՜'�� ��-ge��h�kX�eɑ�W���R�bT�b
��g��hfж�Nuh�g$�M����@v7/�����41���e*��n���Y�ڗvc���7d+]ƛq㊺�խ��E�5�V��^M��Ů���%�u��Z�A��QNYV����gR���n�7N� ���s��q��_�b
R�}kGAYR����	�����`����X����٦���h$'5�*Uݍ�:�7g�:��5��S�/�e��7yYs,�C�U���oI 2q}vE΅�U2��ܸ#׹|
�^J�J�O��D����^��*�tjRst.o\8�7��V�>�^v�>P�t�|�����:��1[G�wN	w�*SJv��fwCAZ�φ��}���-cCH9f�P�T �V��*�*m��ԛr�l0K�w�C{WH����7�5$9Sb���!�\�3�Nr�wY( �bګ����e�(ퟻz��U%�ˮ ݣ�u��ײ"�u�*��J9�{o��ƹ��s����(�'i�/O:W�u�xj�b��s�VS����I� ��|=܎K���+^u���Yv���:Ӣ%ύ��,��\�H�Q0GfJ]z���O⯁N�t�5g*#� �
ʰE�W8P����{���{'J:p�#��V�囧���] "�]1�gA})�p�A�րNb���Ǽ��>ۦ��j�w�3�s�mH-�J�n�e��_$у7�����oDϱ0pѡ��}Onk���1�sI�e�bֆ����g  \\6[�C��^=�{Oi1:u���cnh�f����תc��k�'Y���W^�U_sum���2����1�e�Jus1�̰��B&+�ʚje��0ލ�·4Yf�6uJ��[��M]vP��\WKi]����e��y.|i�șwt��R��3���ꕫ�V@f�+ㆵ�r?�s�'pR����|}B�SV����z��t#�Df�-D�q����3�i�1V�Y������b�=�Q�.�6���(�5��Դ�-�k�81���5s0ɧz���$`-���%��=jns�Nnc�m�1Y׺��{���.�X;�E�V�x���\�g+��(m�أ�N=�i��/�o�pN�����н��J}�ǋK�]9����V��cʹ`��("��mVJ�% a��ŴV*s7�j�ANl'�U�
ǝk��#nZ����Av>�bS�+oc����3s��cIT���V��Ke������tl ����>�l��������E%t�9����Z�4VS؞��.l��װ�$����$�ζ�7-}ڥ ��孺t�k��d9�k:�å5q)2twt6K�|�f*Uko
�{�fJ��9�\�v��.���eO2�묱��UҳU=��;��f�㺊�ti��YCu�����l�����"������ͷ��{yƌ������t-ƛɰ�&�Τ2��ɿJ�{���g���L��&*��H��X]�Tt�q��͎h����^�۳�����7";Ʀ�f��]&�i���(�W�K�@M��>]�P�f��'���"�PI5�����o9�3UJ����L&�8�2��N�(w�����f���5i��/��h�Ȗ���0uj!J�a�\��3��#�����U�*i��ݡ����:K�<tU��﵌�=����,R��ޘ�
�U�oh��G�a+�ht�������Y��4)��خ�e�Ң��\��S�Ġ�<ެ�
S�v
�1��_bZ��q��Pb�Z�]�U�����|�vwR6F�{�R�9|�T��C��7Z۽�aS1�i� s kBxKA���u��.�d4����zr�o�I�M�z-�_��L�cfP�3wO$޲El���@H��p{QJRJ����)��(Wr��ȴ�1���u�r=��b��l({�Jn��;�q���أ��zJQ5L��5��.��%5J��U�je,y}M���&7�:��u�&顃F@�0gYF����A�u������4�[���
-�'�#4���o��'�����β����z�w.���2 �9s�bmG}[)e�����:�d���
���Eu�AB���jܻ?,�HL|��OCuʲ���q�-9���]#ӱ�JL�1���=z�hH墕�n��j�m�xBo�J��;�Z�]vu
۹9U�b�ଘ���4�`W�ﲆ��9�|���Z�H��Tq/Rs/yd�ٵ4l�5��W�t�*���K����y��7�K^\���1ubvJo ھ��� Ԛ�̽h�<��>Ҭ�2���X���ms�Ñ��Ǵ`Gqߪj�-�"g1=�H�u��P|5`o%7{7KdrXnK�*$��}�)o\g�*ˀ�ЊY)e�jٱZw(U�N���
.�g��]z�V��j�7j�u����b�7�\z�����n�=h�W.�?)o:ʮt�'r�UrP��0٢�DN-s�7*rv0H���ysfgs�!�����Cn��jm��g��sW���t���w�8���>�=�z#��9^AJ�~��V^�oGiœ�p��r���*��Rw�mg0���mە���Ww`,��/~q �����%��h��Un�)�W	N�7&M�"�(p�ۺ�@�ܟ<���P;��6�����jK�Z��]�riۖ�C��q��sp�&I;�ν)hr��.��}S�d_��՜u�O�Q3��K�8����=X#�I�t7W]u;#��b��6*S�8������[O1u����%!�{m�B^R�prsg�kvS�6����U��p�t�q���n=��ƷZR��c�>��&���K���>i��ֹ�Y ^.�(�]ܨ� �\��
�'ӍՈ��4�0 6]Z��|�mբ3y@V5̢r��=p�dYs>�fỼE,X���w+=�+�s���b��d��X�N����#$c�qgR4�Qgb���;��f�؂Z���K�5���JB�M�S��Ҽ[6����^zr������]I�&v�7��6RV�� c�`�\�4)n��ѥM�U��Ɂ9x����pCz]��l�����֑��+N#�|�v�y�tLh�� 0�D���.�P�o�ԓ #+�>�.*2�'=�0�O��DL�`RMS;FEˬ�2�.7���+3��U7:ڌ9��W#G&B7��v�;�:�������7���4�Ӈbӵ$�He��u�5bR)�a�}Gea��wknūB�av�V^ʼGZϘTP�\�&s(�}����; 4+f*��z�^�%$��i:i�/�`����@'m-<k�б5aHP[ �G������l�EW�6+�'�Xm'�ve.Xr�5��{*��5��Jo`����a����"�ڸ8�43���[��m�B׊hT�
����9��8Z�X�.��_Y\���3'0��u�=F�c���d}��Wmd<�⇣�|�9Ak�t<����K��]B��wK�+]K��SE��B(����BH���Et�\�5��9x���K}��q�X��}��,��n��n�޹��6�$[h�f)���9V8��B�k��m��+�,d�P��jn�GF:ο���H�Z�E���sjV�5�{6U��	JBL�������fd�]��c������[��Y���y����z�]_9o2!��g#�E5�W\��E�ˀ̾k8�&�ͺ�f����TŘ4L���6����q����x�ٌ��*D9�e���O��{���dp�뢵a�u�MB#N�eY�V�QKV���ŝF�T��ɑ:U�7�8T.m7���kN���.Y�ȹvR�S,�^ /Un?�r�i�Յ��H�oN�]�7e��ƙ�IF9Q��c�F*��ۺT�D�D�ex�DBҵ�^�Ep��ooj�Bݻ�QZI��v�C�"�֖6뎄�|mMs&��E�Yz&�b��f�G��y��,	VG���e#V��Ƭ�6�ZR���-Z=U8�$P�eꙴ�B=�q�T���'V�X����֣�q\1��5&VLu|l,}�ۅ���w��F�qf�DS�X���.�7*bj�":�rf��I��"Z��Cz�xyk!^�%dn@n��R4m���|��Vx@�d�� �Ю�/GV[���=��%������y�Ϲ���qٲӲ8MU��~��N#�g䉫��z�(������SV�빻�n��@���ɘ3y\*ѷΥ�}ͫ�:Gj�1f�b<kVԮ��>kzk��޷ϖs�2�{\��:���D������t�μ�k\�*/_Z�1.�-E�٭�·�F��8�k�Q�e��*C�{�kVe�0*G�	)q]���1в�|�"�<n�}���5��'�EQE�nh�	��6�NZ:�$�qR�7	���;���v��C�|�Di�Q*�H_]5�m�r(L��(vN�);�Z�v�,ɨM�w�d�H�i���2��S6k�bӣ[�L���|�[�0��:+	��U��;(�7K��& �ݏ����X�D������H�1\苵��a�5��l�fWY���#��ȲWp%�jj@:�eT+�Ɠ5V]�J��;�!�'�����̢7�`n�u<�v���{�N8��(��Z�*�`� ���X�=�K���z��u�Do4 S��f��3UU��-uo���sy\Ϋ�φ3xx�����#hi��M֎��ӺX�����[̫�8��2@�1Xv=72�s6��Yw+��ۢ�!H]��q�	oM��8:�;��]!�Eu�K	B��K5�#֖��y*7t�m���eY��]����[�n���0�Y��P&f
fnqyƍO�^G�iEJKI���đ��Z۽.i���P�kA���R�*��w(	�~�ujć2�ǣ�EZ�w�&gu1��!)���:�g!}�h���r���_j�l��\�f:�dT,���\C·��<p��)����cl$�ͺk�SxM��;iw �A�f�h�����F�7��򥈾3'u.Y�we��]���Ǉ�ݪ�D좷cr�?-|%f���j%茡�Ⱦ�HZ���Kx��^�'Rd�}�#�w]�#\�c쳐�Ƃ]q5+��-��W�-o%��E+/����Uf�R�J�srȅ�Y9J6>���z��v�q�C`U��=���5h�c�ye��u�]��B��8�guLN��W����l�}�\˓��Si;*�,M\�.�+ѽ�M��cr��D��B����f���Ъ�X���� 4=#�V���ɉ��2�]kΰB��+1�t]sVlT�Hk{HAc\�xM���xa��N��Mt!2��!w6��M�۹\����JL���i3Y��K(�liۍ+����� m���F�^��yS�TJic|�$ݝE�Eoz�f��}�k��'agӛT��)Xz�g%԰�e�d�+�ꆭfr��wQ&S�v֛z��x��mN�j��w\c�+��Ղ�_���P�y]IPu���z:�*�6�ַ6b:�2��r��ЏM�tGu��w��v����//X�O�罷x�;(�]2����+T��qNH
Yl4��S#�7�9�n�]�\�ט�p�Ř��s�iv��E>�3T۲�ܩ9PԱB2�^h�gh}��jM��N$nl�t���j���3VH�N��Ю�jZ�Y���.Z&�"�ڤw�K�W�Q��I�7pn홽7Y��y�Fbi��s����`q(s:1Li���5��k�p<��[����Db�A뾗�jT.:
��Y3j��[*�L�S�ZMJ�z̫���Rs�J�#y1`��x���LO]�����]r�E�>��+Q��ʀ����[]�GV�{�.��Y��K2�o'ƙ�����s�bT��� u����j\�W��ٽOA�ށ��Z�3�:����b�]3���F��1�1�J�glh���]N���Q�Ӟ�6�֌�sk��хT���t(K�Gw�Rq<B!����/Q��3�u�5ֻd[�V��+/��9H͠��r���g��4̥[zP�Pv��4jI��V�ԝuwp��ne�$�����+=���h�y�t�j��D���(D4�*��zV�p1��,����E���Q�WR�v$����7�]��n��b�mU�j��5#�`ŝ�o�����0t�u
�oN�t��n@W�\�S�I}̛EJ3މvep����@dw�9�1ʱ�D��~��������7���{��o{�_jϾ��Q?]��^��pe%�b�$F�u��ʾ�VP�{�\`�˘�:�Ӧcyw�f3O�x�,}m
I-����2� ���&�3���o8n�:�����AޒB�{W�/�U�b_+���cJ7�j�7R��j�MU�CQ�5��h�Wͩ���gv���jDRvŇx��}��;�u��1,gӁ�4��v��
�wI���I�sf�e.ޓQ�8�W�6m�1���In⃯i�\�Yz]#��*���o�B!���M<�n�z����wD�]69��i3��[LZ����sRD{��slk��P��0Tđ��M�w�N������b����\�hEU����N�k�s"㗴���� yz�4����Yv�r�N��p��� �����f��H�VY�5�aC,5x�6w&�ՙx�l��}t����Pə��-�����>�@��̰�����`�Y���B�Ũ��&ե[�i�����i8�6��0���jA�@�Y��цbC
,.͙'Q�J��nۊ�Η�v'˭s�n��U�v*o�%��o�]�S/�3@��IW%�6�M��j�>�׽�Z����#��F»f��U��S
8��_�Ls�t0gG����	խ��ת"z�=lr��P�RA�:+4�wv���2V�NR���H�E37Ҹ����Y��w=�[E�"�t��;�G9oM���rҽ�[�ӡ����muk��tyK���khs�!�!?V6�8M}+��Q�ʚ�CV�F�əΌ���N��δ��Pt�zuԃ1�]��SD=��!�(��h��4R���w�n�Z�;\+R�iY�뒮U���O7N⓴�,�vo�d8q�cX:����̘Ÿ�v�l�B]�6Zt��r��G�m�Ń�Y�BV�@�`2��5d�B� ݠkFbf�_4)����N�E��LC����a����8�B7:��
�2m��VKta��+R�k�/�3��	4ua�.vK�.��Xu�n%+��f-�CyI�yS��yL[��������Imu8;Qz�ή�o�\�Yΰ�]VDįGY@�� 6W
u,��Qb\/5���X�v��"ʻl�vH50b�78�IR��3�2>h�g���Rp|����V�aV�:�)��qVSSd�5�Gjf���\wx`֛h*sv�d�q�c_Ì�G1�y5���n�][n� �ņb�_n�ҵ�gu�V�I��e�w����-�b�m�� (T�$.X�J�D��	ʁ�x��Mk��Pe�����Q3y��iH;�}�;xqz#;�Q���̭q�JrF�nY����EQm�}��T����0�H㹗�v�.j��9��Ɣ�KF���K�5B�]�����;*�Zw�w�d ֜�Ov�ndTe��!<�T���9<.�:��eu�(:Բ]IC[+u��XPv�݇5�w��o�܂�6N��Y�m`SP�(Q��.�]�vJ"�U3(��]jwm��Ue�>�`a+'M3���_ڮ��)+����(e�m+�~��/��ёK���͊��i�s%CY���nkF���`��e�^C��O^Ԥ�n]9au�´质4�u.�'�k2�_s��9;��YuJ	�7:�j���VR5���Y�F�g�`�Y������!)�]�T�WDY���fZ��O��Q~׉88���<v��Ȝ�Ԧ��t}��e�QM���ך��v��9�qqv���5���	�!Ò�ҭ��Ӫ.�Z�f��|[�=�-X�vT9R�I卧�W9ű;e�P�`Wk�E .���t("�[��aҒ}��'Z\\!˜�fq�e�:۔պ����v
+1!B��s����=��1��ZQ�!�.�I6�uwWt�X��v��kj2�'udT%s�ҵH�ꚶ�IbÖp٘--+@xc1m�6��=@G{lX�;}j|ɘj%{��!��ѝL�p��]-oM�Cdܕ�֜LX�3UhH
�^pZ�1��q��:��������,�/�F��5�bz����2>����9wj=:���&ob2���*�U(V�C��JS^Z�e�I;"���f��(i��\-�|��Uf?�!��m\Y\�{���* .�&rr�����u�=AV��]t%�(�F�'ءJב-mtV�2��#`�R	Q9v��f���
	�a�.�v�f�i��%�[��g���F�%��U�o�m���Q�}�-뾏+8p��Ѯ�Fr\И6e�&�ouh�w�W*�{�M�/Nܮ��Zg�6"A]��v]L�X~�]�nup.�\�y=r�����Ƞ��:�Str��ۨ��Y�rk�%�����W	���`��sh�ea4��wM<��k�f&ݨ����k��z^>�,�iWY��K6�8r`g65փ�oE��*�<I���b���Ng�R؟m�Qt�IT�����v��׻[hB��*7G3��{����f�3�-���é���B�I@A�u�f=K�!�v���[Xp�����p�*���3�,��h�j�#!;Z��q�x�a�թ��]5D�U,�Ew&SB�Y׭`f�!W�g`q,I�69;1J�)w׫5[�w\�E�%u�t��rv:VQ����t\�TN��s�n6�77x�(��j�0�u�p:М\{��	�{!d[�x�+��r>�}{�9�:��3�����]��B>ttQ�jk�J���ԋa��j���Ļ�λ�&�`�1��Q_0�	�6t���U�;T�.�GU��e�D�;~��`tV_1+����c�����s	�w�q]�Vm��ۈܳA�S�=Yݒ־s\Vմ����f�]��FوWG�#+�Xb�o@i�eu��۾�dt4V�x���6u�v�6
���{�D����L֕GR.]�;�m��q��iK4��k(X���x O`,jjL�#��.�I=`jv�eg^�F��lS	d�M����,�M�fD��tK��㠍Xh�?n��v1���4���P�b�I���R�*1;u��.�c��R��N*�(8�돞�^=Qh_p�E��5/r�] 5b����N���j��W�*�d��]��Po��-��0l�u�з��[K%Y�N�8`r�Rz�+����� ����!�.�[�4��Sq[�l���d�[,l�wA�
d�5���I/���4mp�ұ�,Yi�=;�khl�,V�9��e$Vw�F������y���7X"�u��ەɋ��z8{�]��u��ȁղ�*<�:�$��{��5�վy���s�,��RsC�`C��N�YJU��,���h��#5ܵ/T��vb.隵.�)6�8��+ ��xN6�.����|q���dN�EQ:9��Y©m'�G�խi��4����
-�����X&vv+��%�rT5i��ܕ��r�c
��:�2e�	�Hsȥ��V��o�v��y�����Ds�[����l��u���8�˖����&����,;���zn�4Y���/O1V��
Ăۜ��9}�L����`Tѭ�]���iR.� 6�^
˶jfk��o��\���d�.����) W]54 ʖ^*�/�QƱW:�����#�s�T���A�Ef��y�e�}ݦ��$m��^��u�y˶R����j�ά��\���S��͆�!X�Ŷ��f4S��雵2"�!q��vgE}:�[1��ѭ�88�A;UˌT�A�,pyŋw�ˆ1���5|GS�Cv�R�s�^\�Kl�+�z��h�iٷP��廤y�R���Yu��Z4B�x��Af�V��&K�l�|��KZµ �qH�yw�.�G/ܶ�sia�U��a�ҡeM��[("� ���Z���v����O�����Փ�/�'V�����.��:.�ME���t�&�Y䕫� w�����oi��d�r�+�[����(�p��ۮ��d���M@m�e���9�v�&^oM\�B����nm��q�V͇u�9P@ѷ���16\���6j;,`�Z�o�nb��"������qܐ`�شm�.�[�+�n$u��U�赩�ܸW�����b�B��@�fP2����i16.�*�`Ϸ��AF ���>��+]q3��|՝�Cmb�Q�RJ*	hu�+#��pw+
�7X_vv�u�t�-�5q��7U����p�y6n8n�ˢw
���:�o��t<d��]�.7`���(e���9E��h�@�2������t^�v�ݢ�x�cȰ��|n�]Uz�"0�0����)�ʑb�!9�dGC3wV�t�p|��=˗���7�9���%WO�LN�v��@�E�[�d�/W_����l2�qFt���Vս:5oj�Q+V��Z��4v��Om�ǚv���9�WBfS�N��R�a}�v�մ�q��uy�nś�l�$q�����7 �ͧt#w�5�yz�.
.���6�ZԞv���%'R��v:T��Տl���E9Jn�2�0mm��\�
�w`���e����#5<٢��x�]c�}Jl�^S�]��ڂ� 7+����z��������S����+
�#�'zNngn�$�끊��u��:��i���J�kI��5z�r\�|�~YF����r����u��&Њ�����LCϱ�P�0�֬�w ���)	Fj�v�J/��\��:�첟b�bݕ͕ɓ"n�sC���L��Z���|��w��fK�:��%j��c!�3��^G!P�7�.H�^���d�P\�Q���;���7�..Ķ��nuH�h[�����+޻���:�!�-�}oaH�3s7�zs4���A�2�BUL��g3����E�	���+%�+hfgƥQ����.k9I�	���:v�
o*��6`ێ��eG�*�u��QJT,s�\�����?'��t����=�wQty��V)e3�%q�*�wby����+��r�U����,x��C�tԊ�j�r��2���Sͭ<��8\T6�,��K8D��<���s�λ���+f�N���e;0w�n§��vk8N�ޅb���$]�)�Q5��Hup�Jv���c��XU��ۥ�0Q���EwC�O������QI�b���j�`)���j;�u��I��w�"�F��C�o*��f��(�ea�p۴��u�p�EguM!��,�m]ݫ�z����r�cЍ*|��fF$��U^+b�����6U����u_m�X<��{V®uqCuEw]�6ڻ��j�0�j�9g�� �NNn��ζ;<BSI*�  �Yw�DL�<�nl��z��%NĀ�I����jU��F��#�Íjâ̽��F���T$gm�I��.��)��b=�5��h�&�ݪ���kV�L�Ą6��Y�L����*�ۭ��Rd��nS�]6��ݐUY4ʻ����a�16���CA=jNw��>�WN��Մ�vf��oh�}Hj��ۭN� �5e��Y��5���F�L���Z����F�5!͠�T��X�gW7Bܕ�;�C�s��\�քN(cO�"�\�:�����B�m,�������l�ە�-������rk���,����v���k�J��V>< �M��oP�)f��>�5�.�X����{�oSOhtSF�����.x,<ِ^�-�,v�l�;Wuc���/l�6X�VH�v�XG
��o���ĺ�[e��V�kl1f��̎=�md%fD���wVipg+�I��M1�s�J�@v�]�ٚ�' �������T]?M�Ւ%y�4t��eq�B��y��EȄ�v]�3�rٗZB e����+O�B[r�R����k���Y����e�K�\��s{8,�[/x�U2ӗaQi#8;��]�N�A�z����h�О�&W�:�Ci��,�]�g%���n]m_p�5��a�L�d��j�C��+�B,�Gh�MJ�״�oj��'n����8�wiS�2��lj��4@��]�9|�D�5,fɢ)���9�3u�( ФZt9NG�,�"�:uwNؐ�B��>R<;�� �5w^m�1R;�p)��|��wB�S&�=���]̲����o4η$F�fl;��t.�{��)�V�gf��#�]X�0cJ�^u���<��sӌ�L��bؽ!�<q�ݸ���X��K�ndT�5�e.�6�-G" ��7��qR�wJ�^��Шu�Z�h;�r��W���
4z��L�M�5j���nw�ܔ�Ă�o�V�,u�]�M�F6��������XE)�D�>�-lH�voAѳiY঳�@"[u�\�4e��IIbw:��	�R��C^X��5 �[�䫜�gk{�nb(����An�$`�Y+:gQKjؽo |(K���i�f��ew=�sm��a��4%���d�jʎݕ�$�r�3��D��&WmZ�=1�&��y2���F�)Ij���~U�}�a����>�l�2��Qw�����Z���.W}Z��hݾb��{�h�)q�lv\�C�c���F�J��bo�wL�E�D��Зj��%e��
 `�S�����\���B�r��|�f�U�\Cb��mubFgV
W\�:�6̮�<�%��C�d�KZ#.��.�M�>}�$�S����O6�hs�ATV�eh����#/�j�e2U\�r�cʙ[�����T9`��{��@J����t�*%��
[��4�l�5�}�OYN0�F]o�"����r��'ei��-�C�*��|i��gi�Ģ4����fs_t�[�g?�F�X�捷֤j(��W��(՛%�p��&Z��M�7�1��Cf�1��+v�u�]���9k���i3��e�c(1@��pC3e�	�2���Lt6
&p�2�R��駯j��9�}�����������uy��i]��∷��4�6v�q����fbky����O�(�y�{E%tח��><�i�>@e�� 2Wö��<uK�&�z��0q�%�q7VV��7������DS��^<@s��\��]�u�w�e��Nnf:cK1Z���Oa�Ih�X4�sT���;��rSb�.䲃���Ψ\�n�t�j�渽��]B�HF����aRu_t�&�%W�'iW��`�R�^'��̤Eݕ���z�#!�-�d�i���P�V�\ٶyP��ml�
�u����ciR�ר_(^��.LJ��H0�=d=�d��g�����	
��[I��T��g:��T�c��[e��N�鮎&/w.�kU��[XA�YL���v�ocU�m;�r�v�eh&ە̾=k9	���w�� z�/��[�wY�Yv�Z��S �m��p�%
�FF����wJ�{M�T��=���3�iU��n�H�g�k��d�@��A�ѨR�N�f�T��C�d����/N���<VJu��VE[��.2ILK�Pt�r{Pѹg�ڈ4e�`^w��Ȓ,��(�qI��v��x�ᗝ����J渍/Y�\(�.GC*�A�T��K���Nk=OLɬ�ͣ�2ˬw�!�2M�6�V�Ul_J��P+��/�"-X�@�sr]�	p�J�������c����-��e�o�=ۖy��N���s�:i�WN7+�H�vD�����U\�\Q�qV�{�0�*EmʧP���iZ���M̍C�Vzݗ+�壡�.k���u�w�Sԋ�N�57wT�^f�����wv'/#�W�#�S�{�8��HI븺�^y�Q�����By�rw0�8ui������w;�+qĦ��&{wV.�s�E�']۪��;�5�&]�G��E���-:VrGt:��T��y�y܊
uYj��(�jt̩̼�ˑiy;���Xq8�S����w吡�:�4���2��s�'�u�wJ�#L�E��� ��[�Bt<ʯ2T4���I��n9{�y�q۹g4ODu<�<��]Ɓy��#��,Bt���K�\����B<�{��GS=#u�]nJ�ǝ����z�:�nZ���;��*j��wvSd��LU�Wt�ꔷ�Zg1���근�h�mu��R��*>q4�^mLq���]�Z��Ҩ]m�?���6����s�f�buY�PS���]�!*��
��]�Jr��QW+jOx(�˶8�m������@��F"��:�t>�¬[,V�d�a+��5vZ������Jr���e�d�T+��d#�[?pG֟϶0g��O��೯��^�7Pq�n����1:�������i�F,5Q1�s'G�O���`}8Bk��?8���R��}p���;� ��'���i�z����AAWd�[�d��ڎ�&��U֏P��׎��	�|�+N��:���+��J���ᢁ�K/q�pf�=ժǐ�'/�?�;��/�r.vݬ:ezh�Ӳ���yLG9�5ձ�Tk��V�Л�{��SK�4����۷ɉ�&/�\,���g��E��Z��o5\�p�k�j{YEb�ם�	�>�W]T�1�
�&�����,����N)4���l�4%�o_q��!��!ZmWY-�Bt�fD����?��MJ6kOZL����R���<l�a���T��]����V����f�۵�"��V�-���멹�YO�2M�#yP7Y����u��iPW��	���`܃C����t���>D�Wk�7��s-1�MojKt3S��ec��+t>��\��jxt���P����G"���Al��q�]�w��<1��a�!
��RQ�� w
�	Dԫ��rY{��qD�!�\�s���놌���p졹�u�M��q::�����T;L��Q=�Ϙ�U�� ����be:�=F8<�1���pF
�ա��D��,"C�Η�;<�T�.u�מ���<�\M,�@�ȍ$lJ������^r�����Q��UH{Q�*�U�QK��X��e`6�� h�R�}q����!oc��ۊP�g�Ry��el�מ���ҺOv��y�����<K7�y�=����$�����J1AeOa�TV�j��මS�j�+P��;Mk��Y��F1������������
E]��5�羍cՓ,���֎u�u>�Q`��:j��,��X��s����!����:��a�cXssa[YC5����}=+��~f�6+�骎�pK^u�}���e�Fq:�bښ�����s�)��>�z~w�R�m�.�v�k��v��x0K�];������xG��xf=��=����z��r�>ޕ�� ���ߜ��5ǹ�Z:�,y`��{We�@��������:���+���⨗x��P�uL�������,sH�z��|{��-��"0]s��+[�㼊qo����j�Jb��<;ֲQn����-}�S���`�ե�F��2y��j:y�I޹�h�r��wI>ڊ�V���q<�g%����^_�s<#3kΠ�-|�4��<�Z:޷�7�����9fa]ˈ(I����zU0n���9l�N��1Zxh��>�$ ���{�p.�ծ5����@�������Q��k�([08�m\>�8��(G�%k�O/���W��W>|��N�8� ��E��h�+�.�)��"�\���SF3\�:�p6oYf��)Ѿ|f��9΁������.K1�,�2�R�	f�6��cآ��Y��lY�:c��wv��i�5<\��7y����0E��R	�G��ƕ�r�lj�}�H��]��/}�M�[����G�Ԓ�c#�e&�(�D�t�R��I�����>bt�&�4;�
t��tn�9��Q��z��c�W��-&2��[�َ�.q���>W�!���S�#�'5���"��J�>�p�����\�D9Ol�nxT��i٣p��k�X�˳$�qD��AH�z�!T��`�-�r��q�wŌo|�1��Y<���)��h٧Ot��#�Y�v�g�VY�\�r���#�X�\+b��>�he)XF���0�nW)�Q�7������{�*��M�grmt��\�dX2��}v�+�3�w�;�r�hJ��s�ӹ��9G�>���[X��o�؇�Z�S��/����L�$�]���F�O�=]a����z��$�a<����-��K��}r�>��cE���b�U1��f��]����Q��r��$%S!��
�J�%��m�<T����5*�x_n�[	�4!dVE�N����t�ޯ�-T���/E}ޘ"��l�f`�p#�u7� sُ}ҁGo:0��Ux�;��e��b;m�����B��\��ˈ�C ���l�W���S\�����iPNsfX��1�S,�[��
��������+�z$�d��m����j�"5�2��"��VF�Viu�����g��ph��9�+�F>����R��s��30g�	ٞ�=�Y��J�B��`Z�a��B٧X���U�K�^v��O^���,��@���<�J.7E���Y�/O�Z������\�Uպ��fb#p��46���Ɏ� �h�
�*����{91��k��b&���F��`���0��Z7<�O�H�wWy�U��8����jZ춎J�2
�j��&q9�{���O���y��r�U�N#J�S�iL%]m̴�i�t���G�Y�J:�����FI�P�ƪ���Ml�gs�[F�F2o��e�jz�w�h�m[	I�8�z&xo���;NCrDk�R-�FR�D�"|��]��}I���`��[��y9+TxC3�c���)�f �)\�
���_��Bd]�k�Yo<��xS�;+����\r�rV��p��E����˭�0����ŢU�_D�U m(�˕ o{�Z��9��7D�߂�i�#�I�����A�U!��O�ҦKϙ�;Z�sVkb�lr���w.4#���DW�@�4�Z����f�1f:Bڞ�ګ�ծ;
��9Ш-�ʭl��*\�o�Y����v���G��8�K~{����}�{�h��u�B#&�a���[��]�\�],m���wT4r%1]u�?z⪶~�+=o/g�w�LU�f赻��*%�9L���j����zPNg���Olޔ"���Q1������Vׁ�g���Ր��Ƈ�ON^u0+q��2S�b2%Σ��M�b��� 3��e5v���(=^�!�*�5/f�&�l�З)j�v���2'_�#��u�im�Br���c(=�%�r�C�!|��7���n�Y�����X���U�b�۬~'�1��:����[?m$�-Dr�-�9ѭ�G8�5#O���z��2
�)m'�I�X��Z�7x^�������4�;|�1��^��*��I�n�R9�z�5�vߊ;�w�X�o�u6�Rj>�TY�ݏ�d��Ԧ�s�w0���R�������O}���r�����gָ���<Y\�t�W���bWp��!��yY�v������a�[S]-�1����-d�A����(	�>�W�uR0�N>�ƅ���iH�(��q�:�=:�eicD!�:��mp�ƺI(o�x0Kٚq˳sx'�Q6�ˁ���c��r���l��w�F���3�T9�!W¤�#r���9����8��%0 �$90�"��jw`)�����ڿ���eϓ��^�����.��
- Q�V����~v`2�� N����(
�Uƫ�0rj�P[�L*�v��t����a�ױn�@w��-)f��g��!$F�.%m:3�#��r���h�c�6���X�gV�t���񾨏�s�������5`*���.'��#�]�T{^
9��]CX��;YmU-�y��˺����D�Y<ɣm��ʡ�b�**����?�xX�tr�8O��xh)ݧ�n�Bx�j�%<��o�\e{+;	�U��ĲF�`ĿvaKᕷV�R]w��Gͩ����WWƷn5� 
��ĵQ�΂�޽D=,s����9n�Ljh�&��rvT��N-wmwV<��T��b6�l�n��c�(t�}�
 �ލ}�>���^l��Z�.$�ь�}?9=oj�뛒�G0XU�����<h�XW���&��"�/�a��0���s�����١���s����!����:��a�ˆeR���{%���Ny�#�0��?X$T�ݯi�P�r� 7�����|�s1�ۧL���V��v�n���V�����]���<�k���ϲ�y[h����r�����T�p���/�5����+�ݒ�TGo)idV`�=m�j�G_���M�\�4v�iqi��I��ݓ<�^���:MG)L�ߞ_�u�yA[�^u�V��D�XKG+W�w�hm�U}Qy���̯R緂���q]0C�g�N[+>v���i��|�;o�}��]yuӥ����T�8	�˭��_ee�r5;c�p�f9ͫ��g��o;IH�엓��ﳤ} �'<W ���񊻍�]Ar���.X�|�1��a�&oS���L��ٻK*(�T����@�I�BJU��1̬�?p���_�-�u�qw]��s��N5�L���L������U��oM�I��^2ݶ��1� yd`�qھ�u};:X���γ��ָja�)r��m�Km��*��J#�bsuR"�F�Y˔񄓩�Z�.�Φ��ǅʴ~zi98T��/���Y�KL�+zH1��I�"��	D�9@Ć>%*�ll�/w�"3�:0��X��ceJ�:���+�ܫ��.pCg ���w�\9�a$OCtZ�7�4w��2Wn�$��Ngv:*�����q����}n��1��.q�Лbڙ�H��&f9��T֟�űFi�;,�i���+�,=1oK�q�ԇp�I��i٣'1�Td�2MbҕH@An�&sI�[-$2����P
�=�/��OM�|t!���Ca'wB�E��i9`IudNAݜл0S���<D{��m�����b�����,�u������VKʩ����e=5s�5S� �v)��#_�mu�6
����O�<N:��;���~�*�U����=��X��\�̟���������\Bu�E������)t�p�@v/�7٧�n-j_�&�Z<<���TO&"�ڄ�U&Y9c�m_�}ї^B��O�TO[a��ySs�nu#r��mD��nn�Ҡ��l�ޚ�"���X8�=�����a�p��/+)p���^ńn)#�ƌ�(� �s��ckd`\V�ר^um1(]GFZ���s�vww'��v2��E#g.�*K�;v7]�j���Z7�۝p���
�:�_+ȳ5eʂr@�AGfʔ�ɚe�Bc{����QۂpZ�+��:�m�%�v�t�:^�rXޝ�(�k�����P��Ӡ��������:-C�"ۖ�g��O�2�Vά\��7���qOLn
3�0��4j��x�*>O[��,�����{�}��\1�Sb��Aɞ�y�N���� ���.ah��e�6�����D��?I�<�_k�hnv�(�s�ĩ2������-w�w�4� �h�
�*����{�Pz�~6�P���֠��FR�q2�q���9ܑP�܌�sH�$ q�D�v�,���\���ѕ_%���_�]\;%;l�zR8\��m�N_�o��${�~VhZ�]?yC|�Uɜ���ld�?I��R�c8)a�|~�����E��1h�3_D�Z鍧��F쾨RW���f�>��ʲjr�1���9��r���� ��j�1pT�ҖKN��˷'Q��Ρ� u�"0	��D� [V2���5��@�.���Kj]?�{l�*����5S=����jF��ʬKT6��VumD���<���G��:�V�R�#�lTs��c��"�bU}'>YRܡ��<�$��כ,m,�${�;l�Vl����sx�I���\�\W˱�ud@@99�;���p1��p��$���ֈ�ڨ�.^s�Q@'\���Ձ
�{$	���Vb�}����Z�ĺ�#s�h�k�Esx���ʼ�~ޜ�9��9� �Lm�a�P�+&r�����`��T��%�w�(�C���R7*w���[7���*a����e5P�{늲4iD�f�V��&��>kf�N9�}��:�,�bYD��u 7�aC�wAg�n�ogV���랅(bP -2�cmB��.8����0#��QyW�*��	��|̌V����nA�u����[�h��~�}
�C��kKOt+� h��;��u��0;�:��F���Ar3���M:���y��1�T��pxnR��֐̵ĝ$g����pC+Z�&�'��)L^����{�ή�q�Rӟi����1r�1��Gw��1�N��bꅊ�Ycm��ج��n�Lp}s�Q�[��C/���θ@
Eo��Ǡ ġQ��%�vy[�|��Nq�����Uc9�|j �x`�z�#��i�8���!m�Ѩ�t��)4�ns]�x����"�L-$W�g��߂�X�pђڿ�>]6���z37��u�����Q�:��["Sx{+��?n�ƶL۲�6p� �)�m��[H��r�um�Ÿy�N�kgskxڢ�Qт=|�����Qo�]�\#�A�6�]���i����ִ��nn�ơ���-�wmw^<S�/��ӥ�b�w��+��2�lt�Y�۩��Vs8��so݇k�؉��z�Si�Y�����d��w�wZw�1i��:�T]�w�Ԩ��WiI����D9�[�d_\�	n-D&�ˆe]�[�"9������;4Y�
�b�����|�ʝ{u>5I̔6�Z �r�]v��w=(����.M�d}�4��V���.f��E�Y�i�'��1���*�&b��ޣ�5���֝�@|6�7׺��C=��Q	�{�s�)���ا:A��$���6.�
����D���_bմsfQ{K���;]W*���b� V1�lV�mQ�bk3/%����˼5����)8��.u��=����t�	�c�]X�
b`��g�|�\�A]��{z
$�A�\:���,�ـӸ�v;����:7.5xTثx�7{z�a����K;c3�m<�{ ��R?<�����Q0Սh �ޝwX��iڒr*ĺ��w���G���f�Zfd��y�oF־��X5�Y'�XU��Nnv��8��&hX�V��"K��O7��7n���e�Gm�&���U����z������f�S^�A��|��"M���er;�iR7��Bf��D�j��:��ɾ�e�����l8�`Y�{����i��m�go;������3r�6�n�,�iWD�t�^�R)t�PhZe��ݷ�/��X�T�Ӓ�`l��v5wˋ*��<���٨Jb���;��Η��n�*�! d��6u�����PWW�b3���%�hZ��>��Mu擱�͉�	�&�S]i�� �n�alH:�b�c���=�8Vj�L�����ąK4)�c3	�x[��)D]IwgR�ʄ%ţ�]U�3E�	�n,C��Σ���	�79b �f��cf���v.F��U�>:��g�̈.n0+��X�Qe��voF�B[��2�Ȼ,*]z���\J⣷��[F�%eڴ�A����p�J�zԭ%!Df��ٽ��H,��P;�j;cc�X�)B`�I�v�r��u������\º]X
Z�Z����C���ku�.G;N����(��m��J��2Ŗ��!F��ےI��IVoSr�=\llPS2���ZݮL�{Ck�
��d��vUwcF�i옺��F Yi���Q���W.Z�ǴD8.� �L�:h��V �y����WeZ�ٽ���!��9G0��Ǳd��;�庂�z��G+�'�תvY}F:s�lW�]�P�]HlK{�����Q��ʶ���x_m�c[��a������}KZf�˃��M��?V��J/�7G�ӻz��Mj����8�RWv��"	m
�L<���V~+ľo=,O-��y纺z���r��=��]r�sn���D�9�::#�[������)L�F�vtwXk����p��+��Yˮ�&����Nj��	Df�3�w<��6;��wtND�a�W�듻�8��N"��'��Κ�lʪ��Y�gGS7]�%C�$*C�i��WGdYʦR���ȼ�K(JT)֝Z�@B�w���� �*�(�p��y���.:����	sd��{���Խ�U�W�C�E^Bfg�ʫ��FiA�I.�G�q���y	U�'
�O<��㓛��܄��9�]�ćDI�Yd�.Q�r��T��:!�s�QNN]W-hA��d��\кI�d�R�FY)��ͬ2J��np�r��Fe"L�N���=Y��*�rnz�$���r��u��5TET*��|iju,����Ë�#��[�W��*S]�u�/��a����e%���ׯL�P�b�r�Z���,$f^�RI4�@�gs�ǟ���8���Cc��L*�>��P�����:�N��CΣ��ۓ���?[y�����7�O����������>�{��s���$��}��|����";oψ����߮/j�WU������'*gդ�P�nܝ�����]�ڭ�?A��OI��pѿ<��r��~�ϐ�����>��ǔ���roG���>�����oy`�� >�+�5s���_��-s�ɓ�����C�a��<�2�O�����<;�����xM�	ӵ�O��p
oHI;�}����os�!�܁��.�m��o��9�z>8�ǎ��.��m��
�:����x�󦦹�/T�hxw!�)�������P��w����7�=&q�?~��<��������|��N|�s������q'����c��7�'o?-��ۓ�s�|�&�;|O	?��DC`}����B'"���y�P�N���M����=�}w+��x7�{}&����ǿ�墳����=�'���>��Ǘ_�ra�x����;��m��bw��zߠ��;yNpy��w��}4c�#'��>:�̟%T��y4��=�N׸��&q��NWzv�>�����󿝤����<�ݹ9P�{������׿|�bw�k���Ͻ��֛̗��~�zA��ג�/_��Ґ� �x���nX��{n�Eg�r.������S�ǔ��9G����9=���pxL*��<W?�?����=x�ǔ��=�r�wԝ���!�?�v����k���
o�I���<m��1�>���ʴ��w���e�^������o8]��9��������c�ǅp.�[�zO(xMz��w�9܇����	��P�w>N�����®�����Г{�>���'?S�q37Ʌ��M��ȪV�'yU�ׯ�����P��!P�"#�<���G�"Ss��㲘������ݾ�x@����=;ý�N<�W�<[xw+���ro��~B��x�xw���:Nw��]�}��<#т�D��<���w#"�}�9s��Ϟ�>r�(��>!����`��1;�_x��v��o>��￭��o�����&O�������$��=���<��;N�W�𞝼<��k�o�s�ܜ���齩�_&a��6��질��p�k��[�_����H�"+���<�Gv��ۑ��̒�Zm���={+����c��$s8H�E}OWU-��z�R�Z9�{de,��9kB����ݗ�E*�s���q�X��9@]�2�F�FU6�YQ��r�7w���F2�삳7[�	��Ҽ�CD�(M	��}���ސoBu�7�G�)��7����V��u����:O�9>��N}}��<;�~q��?�޸����z��q�p|opI���"c~��/M2���vJ�������^a{����3R��o8oh�<w����뷏~{m?{����I������P8���S�o��;��4��h����>��"8@��2�o.�籴��m��t/j��gM�I�iL�oRfx�cw�܇'?�u� }I���.���7��oI�p��S�z��ސ�z�����=;㴁�/�����N�}�z�~Zf��{��7������lh��|�_lU|��/Jt���{a�|7�^t޷��xw��]�P�㟨ro��@QC�|w��	��bI��M������e�?[w���������ד����"0G�(�׽�~�ås�������|W{v�~�﷤�ݾ<�n=�q�7�'�'z?{�c�nB���c�y����O�x�m������s�j���/�?;I�	>��ý�]��þ�C���`U�7����s���j�I�ޓ�O�Ͽ<!�0�����������߻x��L���w� '�;]�~��ޓ{Bt��X���rx�÷=�7�9�÷ }~��'�� ��t��
Q��j�=��_��C\N���xM�>�!�5��_��}C�G���990����v����8>�w���~BK�z��N'��v<�$�O'�xOO��	�!y�z����)�)�1cV�D;��c�?N���S���oi����������N��>}wc��on�z=��&��o&�{���y���7�����.�_??q�����(r���x@QC�~}o�G�4�y��0�哔��|�����MχnNO��;�[w�u!�0���Ѽ�ɇ׏���U��ӽx��}O)��������&���v���S
o�O��x��z����~�[}|'�>�$y�N�Å��У9#�K�C�j������w�i0��>z�˼;]��7�~Nq��ǚ�O	��S㇣����G����s�[�Ǐ�I��|q����?$�nס���;xM�D�#Y"�Z�7%�^B:�`�GUη��5o	A�3�	�u�IK5k+s�qv k)W�5ƻ����=�іz��v7[Ã��'K�s�էyY,1��Ũ-%���}����&q���k�[X��S]q2A�WJN�^�\�j�H���Di��=�����|���=�7����ޝ�}���8]��C����yq�Į<��M�99�k�F'|C�$����]����.��s����¸��D}� ��=���N�L�^aV���O�����{����oHRq�x����i��xO���a_������7�<�����i7����nt�N<���o�]m��Z�&��/!��?���܇R�}n\�s���y�x}�E��'8?w���n>'8������Ex�������o�{yw��n;rw�0���n��g��P��U>'��7�9�C�=;r��������������^���iC���4}������;����v���1?�y�뷚���<!���ÿ;Toϣ�y�~v��|��}�;������ߓ�O��;�o�Ʌ���z�o)���90>���xU�$U�F���5݋�o�|���!��V��$��>�����N��K��ۓ}B�����]�_ܙ�0��O�z���i^��	��[c�\.N��=}�)�<���Wzߺ>�xG�H�C���?r��ޡد������1;��<��>�&�����ÿ!�=z���BM���a���w��P>��^}��ǔ��M����yBL+�������oHI����x��MKؽ�z>|�۩\|]K���Ko�Y������
y��;�{���7!}����^U�����q���N��+�9���:w��㟮�L*좞�?'�90�������_�������jM�K���<D|�L�3\��ʼ���ԇ&O�{��o>�!ɿ�}��G�nW{q���<�rI���ϣ��>;yM�	��[�Sʸ�|�|�rw�ǝ;U���xN@��ڠS��]�؀#�,j H��
F��?���LD��{�z�j[�/bn^gM|��M)��ztG�����r��i����~��ǎ�L���~���oHw�����]�7����v����I���B���.��ظ�.��wq��pn�i7����p�]&���7�����_���I���rO�<����x�����?'&�zC۹�]�O�p���;�������7�z?�V?�B���%~ؐz{mƜ���lY]��ئ�W73����f���Ԅ�ʵ2�궕���v�5tj�Ώ+ ö�*ԧ۰�5s������3^Hz�B�ĺ�u�wrZ�e[#j�36V���״�;��ܚ��f�;If��zp�v�Dc�e��Zx*y#2�R���j�����CC!��
���¿,y(��r��o��ü�O���m�<�ߝ;���ɿ!~��߾xܮ7��~x����ğ���&��q�����;��8��㟬�P�ٕ�q�Y�|�} ��@�9)�)�ż�����&��B���]���Z�#!Ʌ����~��w�׮��������{����I��׿���{��*c�zSBK��3f�tq�9n��zrg�V�;^�8}�?}�S;þ�U�����L.�v����×s��z�c�}�9��]tbw��㿎��o��]���>8����8�=��В�ɼ,^hMM��I�ˆa7��ﯲ9�̉.�6-�ew��� ���N����]�7�~����HO���o�I;{{�����]��C�����<-�7��������ӓ����Ǩ���?;���Nv�~���{��6po�߳ݾ���|�E��}���D���^xWН�����)��o[����z~;r�����ˉğ�)��ݏ(ra_�{����oh_oN�ý&���ߝ'�קo	��|�����n�/D��3�����@����}�/Q���>7��q�������þ�����=�)�]�w���L>���o4�b�7�ro��JiM�Kч��3M��LΙ�xgI5/xq�I��Vk��l*�c���9{P���$}�>��1������χ;I�;�x��_�oI��Q�>!��nN��������m�������L.��~����>\������nf"G�Fǽ?EᏠ��BN����9���ef݊Q|��GB>�>�^��B ��1�"=Ŋ����%H!����3#��J�+j6�e�䌶�Vea��1�`�mWP�B��G�an��G���ݐ��}�8�boPh���p��XHq�/����b:�W7"n��هU2���q�x��.6��s�d�|�I' �(��%t����ߑ7�O9r��$���=�1wa��.�hv���Z6�°i��WJ/�?��c��6�L�+.�^�MɜM����.Sy�-�/i����f���V��kq\[��:֕ZWk�r-��$Q�ڨN8�zt|µ�1q-W+�����a��}I�\�rLޝr�tzu��)�eR1�!��f�6hN�OOG9�1��{Q�A6����x�m��5��SqK�R1�`q��S�͍��ئm����E��<t����-���4��
no��4����\�XK6�?�m�P[�k�iI�y�`rڿ�;�CT
17�2������޲}Se��t��(q�@�t�J���u�p{
cF��0%�.SH�i�(<Q�Xu8��	(�ۡ��H���5��.;���~H��"em:3�#��'���S�#��K��_ �զ�/�uM|����� h���~UJL�J'�w��ؤj�'�L՚|�h���f�n ��;GQZ{�O��mT��O2h�n���m�uY%E\b>�Ũ@�*y�����n�f���B>ڬ-t�?,������I�q���%�Bs]e�v�^ʰs�	�]);Vw��q� QfA�~0�௺�i1{������S쌈\�!]�@��t���u�f=���Wb淪��8�zƾ[:�9����)�t�;��3h��d.���������4r[+:��Wөb���7����o�ޫ��*���땖oLy�Ҭ�c+��B�euut&�8��ҹV�@�6�C���]��z����Hw�C�%�>�Y"����@KV���뮷��:�2rh�5�O.=�]l��^�m����W�K�x�@�1���'��\��]���k�j�v�'��H��;�d�F%C��l�5\"����Ȭ��p���c(ʄ/w�$��z�I\�;r_�s��l�Y<�2������<#v��p������$��'N(��pOi��N���u�7�b�:�	1��˴�`�`2��Br�Y���+N<.j�7���]�Mo�b�|�y��<+���Z�˘�}1@�jv����t�d9���ܝ1�BQ"-�Mb�5�ܜ�@�148��<
s�za#���o8H�r�?R�>��]����W�i~��y<�L��!�6e�K�B�v8��݋	�5���Y=V��iTq�;��8�YG�b�.�[�;��pBoڨ�u��'\���10��J�����C���t-�5b�c�#8�>5�rt�ϋ�����w�[�eL���ƥ"�6�����%q��T�qX�*B�U��X����s8r��w��1�d��H���3�}֥����s�͜R1�͊oY�0.�|`CkK�r���鹴�����M.��7)fju��c2�ZQ@y�L�p������5��M+{k#������@�*�y<9Lg>�G���Ys����`�S2;f\�Obi���M˷M$*�fX��t�(!�c��i��N�6xL��杚7	�F���� s����b>"9ƾH��5�GH�ϹH�~�q����ڮ�B�'wA�]�B{AWv{chY�u=���2�e%
\c��k%�.��~��9��P��w[H�0�7��ތ-<����3��A����X:raK_L:jZL�Yıw��=�;+������-�mD�9�ov���2�����5u�X'�s^��ω�/=�(��`s��k�u>Bm�pjS%�������!U&Y9cۯzwϩ�Cj��(���5�������N?�P�'�gFDt�ٖ���1�)L�r�g�q�ޱX'j�|��3�����FF�BTb��(H!���TY]XY]|}j!	˘'�ud7���|�VMY�\�*���vhT~�T|.���U�*���)֋�y\:j�vE$I9>��Ǚ�٥�;�bÖ��*e�O�R�3V�.|������MSF�dg���6����-Ӵ��^S��B�f��d�r]�Jr��\$��K�t�-�S�-D���=��ɕ�_\pnV�-Ꭲ[��𒵋�t���1��}ϋy\\[j5mp��C/�B��燾V�K�.��O�:�������:�+���S�mH��E��?��ߪy���;M׶47���LD �U% VJ����=��M���QB��z�1U��I��%����1�q�"7��mmx��X��Қx)f˾9��r���E��,d/�s�:�j�x}��Y���N�1�zR8\�
��Q9gTm��Q��/���Hy�	H��z �/���"d��u��7���쨎]l!��e��ٌ��:q��Z:��"_���s���:�	T��0Ӥty��\boz�w�\�2al`(a{����8��5�k��Ν'�(N��S�"�C��;NQ�:k��:�xb��ѐ5a��{٭��r�W]z�4�\���,�KT{y�+;e�Z�<���!� ���L�T��q�p[)q�jB�\WJe��Lh��ʎ��;�9� �N@�?mC��ZVL���!�6��}�����MC{�d��g�s�Y{�` ���xuS];��n���5w׵�M��,��wZ�Ge'%�b�b7|x���@�4T��W���5���hs�u:WEm�^V��@��!����s��r�{{{���z�S>��w��*Gڝ�۵�Fn�s�v*Qp(�<��a��uz��ڠ����Ƴ����菣�����\p8G&2�pS����j���'�'/��@Tn5��|�׮����ekٕ�@ԫL�����MLV�a�C�
�'FT����K��y4�/0&"��3#W+��<�ڊ�nD嗄�~òj�o�������އn�J��/�r�]-ڻg�r��b �������f폜i�$TZ�����*_�n�o�Sm��V����<]��%a�<�T�z��^�4�'�j1+�Y��Ӛ~ae����1�9[o�p�İ�H��/��L)��Z���*�6�R0����Q�[��2��@�m<�.	�R�-�+Fھ�}y7�5�.<
/�	�'@�y�����V3-�ǋg���;�F��waN�"��)�O*�ˊ��,�t$uG�
��$3ܲZ)�gy��*[W���s��2�H����<�Ԍ�Sھk����z3�����LIn�`�9�*:�8=�j5B����P���l��G`�r�C"t��XD�n�n�w�Gƣ����!R�~eL]s�"6�<��^ՇƞN��e��@h
A�^.�ۮ׎�z��I�K<N$��m�#ޛ��5��oQ=cɬ�\��V�]�eE�F���bΦ*�A�t��r_1����i1��{,�h�d�Amu����.�ɗ�6Ջ���jqN���}_}�n�uds��<���}��ѨĦ�M��:`�X����};2�&������-����ӳ��3�HP���;�/��}[j�TB��M���>{v+�Y&�}.7q7w��Y7MKIrYs��(<����}8����ʈj�z����W���'�K���ۓ��̵����'�pm�f
z�\��1�Q��GZ�&/��A��_-�4��1�{���p_8��>6�?'�Q*l��Vh]χ�:*��x���h�j�Ԑ&�s>Yq�!���ݭvgY�N���jhn���Ż�}(�ۃ0����y�ʂ�o�L��L��zO[�D����1\�d۟�l�sU�/�kE�k�|2��$9ծ}�#;���-sQ7��"�n�ڹ�H�l�
�e�Q�2�^_�u�����1{7'����7�Of4'X�wgI4��rԺf7�Г���K��X�)��(v��<n�e��^W7�3ӣ��b
6}Oȃ�� �¸?�k��\�x�ʘ;ަ>�p�}2��.T\�#U��NI�ո"x�4�T���Nվ�Z��W�6�]��lGx+n)}�� �s�!(޺�k��D#�%�EF�?��q�&u�RHꂭ���պ�*��5s���n��������T_[@�����4̻�H}vZ��[z:�r�d5���`i�����|��C;�4��鸥�%�7{#�&�ٕ��-<�i?�x�2�wOJ��opEQ4�,��nmU�Ṵ�enh��l�ZM�\M��)N���n3��t�Z�H�����]��)�f0uJɷd��h!�X��KKS�ـw�����}h�����)���y����Ёv���7�Gc�)�Wo㛻׷Eggp1m���7v�F8ơܵ\��íIܫk���`֩�̾3���]�tvs�P\�!J���S����R\;�c��a�*y[�&p�ǉ�t7��Y؄v������>[m�����V�n��}P)�蕦�YB��4C��un��B���U�n�0J|�
&�����;Z#��Z� �Pt4N�݊v�"��5��-�u�f��W�i�ͱd�3�b�*�&��=9+��"��ؑ�4vs:���;�z�v�5Y�+���(Z%�g��53Q�&L���;��=�w*�}w�֔�Q{RP�h#.�Y+%:�5��tSYR�A�Hn�ܢќN�Wt�����`́d�h��R*XiL��Ko{p[��]��4��>X�]1i��b�ʋo��u<3[f��s^T�:�`�|��F.j�B��{""T�U�y;nN�Bar��o^����zW6v��@�;��T 9zlKll�X�{g���
�%�ՓA�y���C9��#�����lnwб�9��n�.��]8�'L��T �-���%Ē�*!ա�m+9s�![)�$u��J�*�u�ܝ*I��~��^]�,��޺�Ju��r���:��q�����v�r���i��ul��s���S��HV��E͜������*��O�X�Rɢ��oˢj�O��@4����l�>���6�]����x�	�!C��؃��f��T�WU�}��VL��U�Wm5Xu<r�젴^ y��
���1��t��N4"��3�b�>���4̱ګ��"5��=�Gb��f.�׭JȍnQfa��˻������E�̥�Fػ�KQ�K7��y�7�����[n�{\�� ��>�dD\�.�ov��[Yu�a���:�t:�ֈ�8i�"������v�k]=p�=����st�~����e�]<��>�R�kw}f�
�i�����-���[�Wa�y��)-jC�M⑜Vv���Uc�����X*�>vp�e�f6\�e���n�7��a؏�����c��q���ĆjN���t�K)X3@B�Nw���/��o������<O���jQq ��+Z�Bq�w
��z!S�w9Q\.� uH�<R�Ĩ����rwwIȒSa[�G����s�4����͎�Ap*i�C�z��"pJ��wK��*/<���\HV�UM�P��s���J�y]z��#!���Tr�����ù䓥u5���i�Bwt�v�'�TĮ9XT��ww'++�$^�W���j!V{��vP�TN�q�]�/,�(�#���IQ�̢�<ts��\܍5"T��"��Լ�����)չ�hF���r���S�wetws�3�z;��4�4��G<��4���w\�)�<up��Gv.^�W��CB"���y!gu%�f���s�=�GJTC�����5
)R�H�v^�YM�6��W����֚8��;Ȟ�5����M$-�wڕ��i�L;�`�׮�����һ����v�l��>���%�M�uy�~�w��3��@��&2�
y !���g[��~�m�،hh���Ozשwu.ۗ5�F�v����R�V.J5�}&a	��ZM�1̬d2&�L��3�*͔�@ߐq�K�$�QË�|wa:���=�#���J�����8��v�kd㖹�R�%ˎWX. l�^�"���?.N�!����m��.��0�I\]�,�M�$���E�m!�V\ G2�\OK�tt�o�<Lg>�G�9���W����
��K8�'�O+��"���:+����BR���.U����i�ޕ�S�9�Rb��vh�Lc�Okk�yX�P�[;�c6D�Ok���:����]`�������z��	��m���fw&��)�-��Ӡ)�NZNb���lâ�ioݞ8�2M���ZgDIl{x%�r���j�f�C�T�Z�A��Q`�f$O��A�oþ����� ��5Ŏ"uس���9X_Ʀ��en�[z�m����LN~����.�X8c6|�T���v�5t��jj�%�x(��N�)Xj�t ��7�:�u<׾��/�I�Of�Q�����ɿY�M��$e�ni�K�
�Bp+���;�Nn�8eNu�K���('2�w����u^9Q��鋣.j����6�[J��yy#sⷎ��W���OU.�%OV��T;=o�Ornz�I�*z*������S��{��B�rh�b�u�
�f�f$�Ȯ1C8�6�-�	}�K_Yх�啩x_�]xW"�`�t��v^�)�t��褷}V5�6�p��%C&�ݐ�>��=����b+iPEf�Viu�ʝHp�Ո���齦���X!��g��ph�1�,P����U����f����Ӂ�xN��y��P4�ʝL�+�8��U|�ڪ}���u����0��@Tf>|a_�*����z���{��.��f�?Qj�d3��M�=ꑷ
��@�=Q� };�����Ny^�>@h�B*���V7�DRj�ne��e�1�r�#j;���37{c_��S�4�<Mv�"t�+��"g�|+�)�#>g�]\;%;l�A7�#�1�1D^ƹ!@�����ў���o8��W§�H#�M�0�G/��Q˭�1y��ד5�x{-�m�<(U�>�ϝ'Qq;D��0��F��id\<����ix�3H�ܤ2�|Ĕ�Y'��4��
�εs�m����z�]@)�)�}�bg"3��x�Л��ݷdT\���v��ʋCf֬r�÷$Z[�@���q�cd�T�۹�$;��Ƒݵ4<Na�Q����7��	�?����g�>���to� 2��V��uO�)d�̰9�`buD�D�P�7��:uK�����	�*�����f�$)ި�[�cUto�\%�7����^��<���2�3ޭ�=�S[��9Hm�Uc�f���R1Y+g]���q`c�_rAVih&�ma�t��}:p��C{�O�y�U���eټs6\��X�n���=��گrTbs��O�9C�Q�d�q[z��I`5@ܹٕ=-�x���'�'.#:���C��ح�B�E�۞��	�7�3���o�W�U��|f���_u�^��Ҡ��{-��lk���k-A��f��!¶��q=�׶c�d��ګ�{.M�Ғ��%�K�)�y�6�f��� ��;�l����2EE�M�k�b9��c:n��۩qg��Oin����c(R
�x`֚�S󉹎&���X��,����ϴ�����f.%�cMΎ�l����sO^Ԗ�{�x	+�X
��R�o�xb���}�BkZ�Ǚ�CpʈY�tq�g��nf��][��.����,����t���wg
Z9�$o��I@�u�c*�6��/���Aϸ�<
��w|�í;��bY�39Mz�V
�z]�LC�pK���ܭ)�"c�ՠ��qj�Ę�L]-Z/)3�]�~��������ۋ>h�^]��s�2�#��X�ԡc�*�t���b+�������Ǐ?V(��:zݼ���C3�sO��W
�A��� Hϙ	�$3ܲP墳������Sq�^��b�����{<59�'����p%��q��BsI�<�9��P{z?bm_����Ե1i����ڤźD��b�&�u�[�q51�>H��#�S��1�x�����3T\VKG�9��W�Ѩ˄���M��:`�X�����Q?K����s9��N���G�0��u����v��J�|�_ͩ��y�F�t<��b�3.��� Ŷ���q��{ԧG�	,֘��pbz��~k;o��WhϷ�Uλ��
u����/o��%ɪ��n�F�^Be��ӣ`�a�w+�t�
�s5�8�zM^���L`�L'cfO�nR�{������'�+��Ϟ+˞D��p����m��s+�l�4��iE�����ԴujPW r�.�uNu�_CSCt���1n�o��@ꡕ���d~�y����t�bj��F�!Al��z�qt����ڽo�Y�gM�u�Ӂ��+x�1��AX���X�Gs�,��^Õ�7�K��PGy�eA�wS�N�$�Nch�C.�Ș��&:�����2�}�rwt�+|������y��F�uqDҴ��T����U}M����+�	��! ->w!Q��n~ųq�p����W��b��%�Pk��]v�P�sp�e���ۦ���\�4t�A,�j9Jeͯe��/�(+v��5�)�O�-J�M����Ǒ���@h��%�����1}j���N�Z�x�Xo�岌���N*Lw*j{1K�;��3肍}JH:
���u�5�%�S}��Id{ �yR���]l~׳����j���ͫ���1#��I�e �9�pza#x���L�J�*9e�7�mqӚٕ�$9�у��F�v�s*aE�����'�i9b�nHx���y�Ո�=n u|�c}q7-�p��ߗ���j�1כ��$y:�Ơ�v-N\>�6�ݥW-Q��S���<#��q$Fq��~�N�9�l���`-��9�;�Ld��7��NUJ���m!����^�
�O)���.��	����y�8.m��VMvq���*����C�����+� �hiE*���IL1"��(v���Zu9��9�Rb4�ey�Ԗ�f��E�|wFR���DlF�F��5Ư��hek9V��A�(�Y^���]��n��H�V�R�p��y��c��D��p�H6i�yٙ˵�[������Ij��fR����%.�O]���@�F����#�n��l�DDG�D49mN�[l��q�骫e�:�>eC��C�C���Ƭ��7�GG�*i�WOW�N�՝=�{�;U�E��j!9`I��c��u �\O��1WK�-��^Y�ܱ��P	�W[�8!'	�.VKʩ�����e3t4���_C�i������ٍ`+A��5ؔY��[|�A����3�]L C�2���P��N�~���0EN����:/��SP��*A�^�B�;���6��8:�&�Ҟ���UI�L��s~m_�&�x�L�xzw1z�b�c������
�`�Rp�����;NΌ�Ҡ��̰ƚ�"���X)w{���I���@��&���k�6�`��J(�Mɻ }SC٪}�M-�pB���-�!W�dO6n�u�Y����r��u������2�٠+Q��U���冁}��V���{y�M���#�w�5��p���>�u�痵�̥�#�h͍�P��ݪo�"cY��{�q��v���}w��z~��<9�9���!i{�#'7�0Y0��+��Ky՚�������v.U6N\\�9�i#lg �%Z��Nx�J�m�]��(�������h�K�y����욮�~
(sb�t�R�����A���%���d���6�]��M8ԭ�9tu7��2�ܧ �m��`�kOHۏ����ܩQM-h�6}' ��L!44U���oMTJ�c��0�il���ݖd!�'F�x�fo��O�H�x�X���Η�	w?��j��8d/�����%;l�zR.v�k-��y��s=׎S���ĸ��H� �ݔ5D}42:�C�����K9Q�2�5N�YѭI5e�"�+���~�Γ�����
a�4y�CJ�!7����ܕq��{���P&�q��B�g�iS%�X�sGNh2��a�%Z���N�{8��nh�qq�0����!��ګ�q��YR�ˤ�|~��%��<9����W��b��d�BՍ��)^�8n�S��`�~`y���~����=������8�O{�b�K`�0o����j߆\�Иr���Mt�L�!]�?{W�@^*o,�Aȸ�E�ӷ�Vi��b����!�'���1�&�:���C��M�w(um>�I/�J�Ջ��֙��u�ƴ��h�UpB�/�����.��`>��v�F����V�<�5��kC�Y߄�e3�o�;� �"�ض ���]�6�ԧS+�1�ɾ��r�DK���Z�s�j]ڇ�EΩ������S��|S��"$��E,[]\{쵁:����{�1C	�v��U_U}�6�=�[J��o��U�����.���6SR�Eɡ�0g� h��]R�p�W�LImsMIe�˂�tal�V�7=�<�#��pw�Φ�6�R< ���ΏƏ��d[6顜Ŝ,������&�h�Y�J�/
�O�,���6b�Z�7>���̌���"���mЪ�ĥ�D��M�J%�p;��]T�1�+�,��	�j��r|cD!���5��UY�N;y��v����<t��1�\�5'���U���j؊����x�1RT��F��-Y��iRl��b�W�}��T��{��K2<t	�����׬Z��c�D;�(�e���]���rUX@�u|ý�6���>��g�Y���і��[�̞���q��q�'���rzzʤ%�K�������r���b�&�mցoĈ�@�"��c�7<�>��ý��Neug���W������ri7\�,��*�&L���ʛ�j�H\��
�1��.�'Y�A~�}�7�=����y�F�m�W<�kr��5;�w�X��^�P�v��n*p�ް�3%(��G�	W��$)����wM;0��˅U�o$��`Ֆ���Ķ���wP�{��#vbRmr�#��v�\*�c�7�k"�`z��;N\��#��PNg%�&`Q��M%,�ܨ㓿��������j���I���.k㒄W��
����qm;�**�����C�����RW��T�F���.�P��U�t;3g#L ��.����u��b�e��U��QQ�����'�+v��E��5�୮��qQ*{:�赡U~�슡�wg�jj3;Y��ww�v;;���$�� n)�:�uNu�MMӟnO�n�E�t�wl�,2�m&'�������u$��~syPř�D��m>y#>W0�,�}�j{�ѷ���$ҵ~y��߫d���o��2��W/�y"F��̰��Y5�2��|Ƴ�37)o7�͏h���VJ�7��k���D;� d��3�\V�9��R$��u�.�!���6��w�]4s+�ork[�Z��۪4����8�u�\�|+�Z���J�lk���{zԥ�Ժp����1��Gͫ���g�B8OI���`�2H�X��Un�楜�q%u:��.%�.9�4c5�÷�P/�:�h�c��EW2j�C<w��*N!�u\�)2*>��f�0�ѳ*��V��w����>4@|�ڻ�uh�i�o7~-R�d���D�#���ռ�~<j!�dt��ߌ�epyj�*7������jX\���u@�ɻc*l��\n_+�El"�t�O5\{]��ޛǍ2�\���}_WٴyC�w�m�@~�#8�B��wщ������.����F��ڨ�u^o�u�Krmy�_^vd�7*��j�fj�7g�� E��\k�NR*���/+��w�C�f��u�t�ڔVn��&9��;	b��d���=+���)��������7	�p�unx��IG�[7����cM��W�|hiTR���k�x ��	��d�:��u�����	�is{I�l�%��[�A-���Ӱ�g@�8hdyS����ze;E�{B�k���
�79���9�( �o]���wt.`)��N����M���k���>�ifs�o�F=֤l�{s�wS��c����F���KF���Q9�*������P��n����Fr�"L`��)���a@!ꙸn�h�CWQ;��Fx���m	�eQ{�aet���+�U�:��Y�l�����4g\7w�#x�uW�%��1�lu��'y�����N�����,���R�`s�Ö�a/���ti�A��X�~��bI�M���Σy�:Ăy�,�������2��]��Ĉ��3,ގ�FvP�N����׹tjڶe�i�2��Ք�T-.��/����	�`�Y��7�&6;�.^Rcr��a�m�3lML٥�� 0�T6�Z�jJt���ZoQ��@f�wq��'`�b��8�%tZ��[��i���$`���ݩ� �$F�w_~��ȹB���2�;��e8pɯ	ub��e�Y�6���]�(�&�˲٠����O��w��O�
��֥J�h��	;��T�\ͻ�e�b���W���M��R���ĝmXe�+n��4�[��b��5����ԔRV:F"s9m�lL�(\(V��z�=׹+$�@b�G��?:�zpGV�� ��j!
���0c7�Q����t)�u��YMVE��e񸕦tV.^s Nz�l��*����0Xe�3Yq�$�v�L躅�Ÿ�i�4�ſ]b�F���"��R�tu�e�E�kz��^A-����V8����������ً�cC ��4U	�\c뾸+U��Mr��r�i�]�z�_@:E����c�q�����&�u��F�αB�Rr㖊����"X���X�xֲ�1��1c�]Z�l�kweŘ�(ѹ�;yab}�(K���5x�MggP5��Mؼ�veWR�M�F��9��|R�C���Ӳ�0��
\�p���7V.
#�Ͷ��-�j��v��>�L�SF�ޮZWО�~Oqk��gcT�Z�\��•P��(^������_[Jz��k�펤S�9�՘q��W�+�t�M�08�.rs�e�V�@�ko�Tuea�@F��Ç�[�{�6j������einY`gr\�`Q�e����1pJ��WN�1v����%Xܬ�xvj�����qhR<�z�#n��J�E�n�-�!�Y� `��#��}�K@�v�|��㽡�-r^�o�p̖��նm�s��1П�՝Iӭ�z$ڭ���ʷJ�^��n�B�e��ՀJ<�^�`M�#��ٌL=w[�))��܂!��tF^�ۨ��@���?w54R5�-Ÿ�r��UZe����W"���;���x٣6��[��p���'0K�[�vl�ˬm�9��f��eӗ����:���oV�9;SH�63��2�U;�3t�ˈ%��A��v\����/��`�%���V�+e�Q�	�;�,%�= 7���,��rgk`������۔�u��N�`������`>P�b�CK_ڸ�ZNl��|��5w@�e#c��|9�Wms�$�ݙ���V�@G�F�e����&M��Σ��@ө�	w��N��6I��Q�*��w��!�����C��;rAbFg�ױ]t8���PY�Z��@8�/��lu�7���Ҙ��p��@�x� ���Ԗ��kq|Y��WA��VJ��*2Fl3�wh��
gǯk����x��M�qWwk��;�4+�=�'wC���V��D�g���I�*��s�B)I躲��d�	���:���u��2(��{�̑!LJ��]�su��*��JZ���ԕ,�Y�䬪��䢩�\ʌL�::�QJ�g)�%a:�&���I��!��șd��^Y)�ҲD2�ITԵ8R*g�y�]V���	�kB�J�^���<�JP�LR0�)���Q�45�M��<�=\�R+"��$��44��<ĉ	�FU��<�C��[Cܮ�[����qgD�`QF�t�v�2�g4C-
�.GQMLZ��Ȱ�DN�&.k�v�Q��N�!*�=���]3#�"��4w"�j��T��"��bHd�&�����rs�[I�q;�K�TW�Y���Y�T�" ���A�H���Yj;�xD�M�Q:'�V+43*�J�$Yij&u���jNn8�!��ԥoK�x������Ta����g-�>(��$l���4-9@wb���'�uj�=����zu]�7czJw���^��UU��^��H����w���K�@��).�ib����!�(W:P��!���A��v�61;[r��=�{2��顮4�|Z�HE�r��w\ȃ7�*eJ7`��f�� :��ye�P��ӢT=\ƚ��qf��R�؅�[����C.!��{��h6��"�8�o����jwn�o�!�C�6cj�.+]ĳ!��`�O}�C1�h����T�S?%Gi�$��w�{B�{ϳ�N:@�Qx	����hH��X�2������˘c��rn�e��DZ��7|��'U�����D1�d*]���j���5���dJvى6Z�x�(�q�tv���3ۇl�1b$�'.S2+�2W+���Ƣ#=��9xzj��]�r���Lmv����t��v���Ֆr���'���K�:N.'XJ���
a�Rt95y��>��Naڌ��R�1.#:�-j�0�ꟚR�i�`sϨ��%:�u�@�c.!Z�+��-'�O9E�;���C%�����1�ګ�q
�健�,�����()�_��V�6Ha���+3]B��pLԍ�m0�Mc�v"�(��u�3ij��`Jɾժ�v����]�aؽ$*E�-�W�^��y�����V9�8臜����v�T�v���%fVVc�8�8�Ԩwю����b�m��ݙwE?U}��}\� =�s�\`?�G��)�t�E�>h��;Km�kP�OI��9;�8�������B��K�a'-�Q�or+d=+&r�!,v��D�1��K���S.;m_�xb�:$�t1������=�
%�'�%F-ǣ8R��W��j��s�z[/R3pM�djJ��;UzY��n���QY��f=�t ,�n�ot��yS��2�3L|P��@�hOmu��vI�@ᢠ����d*N�
]6w>W_f�W:+7*tݔKW~����q�j�OBN�暉�.��p�P	g�]��d��Ԧ��1R���+)���G��U�r��lTd����R��6�a�=n��r4�J�GONF��Y���
%�cx��1Y*�v.�`�ϫJ��a	;�2�����]uR0£��١5վ9�2��U���9�9滭:�C�ݎ�Q��%Cc	rv`ԝc��n�ƌUX�E7_�������e'{��F&����/�?c�΃G�����!6�)�o��j��.Y��5V��ҚB��Et�b3�x�+z������r�Ct �敃���-���Nӹg�b�`��26S���*�q+���.l��Χ��N���[�5�ev�ոT�����Gka��V`T6�гY���|���=,����}_S/���G���:0z"[W�e�븛z�'Id�y�e����y=��{m��z�]���gKiǇgh�ڲ��k�h���:��MZ�n�1a��mր��N�,���lR��G�t����-~���:7]-��1ZѨ˄��M��� �qŁs�p}�!:&r��򗈯b������^�8�����r}\Cj�E,�dч�ו�2�B�)֮��Y)d�]̨m@v�m1��߭_�.y�R��h���sH3$����e��?<�3���`������!+�<�Z��AVf�����I����ܨ�y]��Z���dX��zet����x�0籬:8��+�*0�qUr	��^��d�;&&�4x� 7��:��u���546�����=0�pЪ�#9C(�(�N�ݐ��Tno��yQ��3-��H`	����S���;�g�,�~�o�����N�},���ӫ-DiN���nEk�]r��u�CF�e�d���S/T<�����m��S/(NX[���8�f�(����n]*�]�g��A��ܲ]�{�f�� n�/k��%�q�_ESF�98��"�V��6�\%Hi�P�N�E�}+�Yx�Q�z�1B�bDs����*=��P���LoUh���s��P���ﾯ���*�Z�?y����u��Z8.��&�0y��u�m����b����t��P2�T�f��w)m��(�/6[)ӯ��V� ��|�:���\�-x�h����F5.e��;89Yc�=�_�z��m�������=�6'fÀ�jR��wf���j���3�%e^��Q�S���i��]g.�Yժ���P��=VE�z����i�NxS�S�P�m��c8��@U�
�뉹nㅗt���'\8����N�	�K�^ʊ���5��{I-=��oE�Y[�bM8cnd{7�"�	�yX��ט;VBd��]��]] 8؂�S$�7�� @x����\tn��L�i�c9�:3����4�5=w�x�����թ\&g�q|�\hiE*���t�W�8L5�[i�ʉvi>5�J<��ՙ{ꥎ�m9=�	�vk��l5?��D��V��dt�+�0	�A�Z�`����̤m�8mF�������X
f�9`I�6>�WSc�=LWJ�V�2�/ur��w��O:I�\E�E�'��-�p��[ha�!ңӚ�]Bթ4� ��7w9�a�xޞ���HS��J>���Y���u���r�[�s���v�,�q�<p;Sz�V�O#�!����]�s��c�qP��x�]�������j��5�~�NOaTX���u���Y,\r�b.!k��v:�KE뺑 I�k��m�e�z*�o�N��n�>����Q���:S;����L��g!���m]D��om���.�CΣ�M����b��ȑ���=-�<T͕�>*��/�T>UI�I����n+u�J�[p�BŶe�M"������p�{O� �pOݳ����4�59�̰�t(ܫ���f����%���nJ��u-�PFw>ج(�Qɵ7b5D��R�d1KUu�`�릞��C�D��������*�:B/����Yo�T.ʔn,����355�(Æ�n��-���eR���c�R�؅�[��a��B�n�znntu�.OٻV�q�x����%��j ���.��"��޻�f���|Z��9�f6��M�ީAX�\���B���O�I#,�ޫM�) oMI@B0�XБW����B�K�CuGʼ&��ro�wi���d��@T��L�C/��r@�R��5�B]��Z{ǅO���G.�q%�Άn]6�j�5��r.��h��X��2Nj;-�])�d֕��`��������#Z�n����I��l�vm�Y�!���V�!�VH���a��#-���lP3��*��gl�/-Z��D�FQu�r���O�n�&諭���z<��a�����x���Pۨ����2�{��k�$=_:��8�[���c��XN
��Ts�a ڢ�\L�x��s�I�\N���OQ�it����ֽ=Ӹ�sdT�rщ�������>����J3,yDF)����$���x�sq��U�$z�;[Y=�N}���7�p�Tj{ld6���@�@A2���eX�U�e�`_o�񌌗O%unM���iz�{��)�d�t]��o�v�&R�G]4绘?G���>�>�kb��B��^�:~�uB�Ed�Y�!�e����dk�:eH��k�Ts�0TWۀ����Ų��*j���N���-6Ch҉"��W:����Rz|�ZD��|)J��p��A�{���;� ���Cuc{:��W��M� f\|P��Fo �����{ܰ��"z@�b8����;�\�l�|���;�Gq�C�^�Iz�NΉk؜+j��Oڂѩ;J@k�������EE�M�k�b:�W7"n�)�b��8��nUM�+�=zr�����ǖ��֏j�k'D�cХ�ɤ6�sz�(p���S)�<��Ve� �F����i�_Aʍry3��_Bnj�{ǫ��b��r�fWs�^q�%�qEXi�3��:�:8��QKW����":���N�m�VC�����3Hc��n�+Z�"����]=9~ae���1�������V%���ѭ	�NWp�$�({0�uR0�E)���	�j���.�.�UԎT�o0zE���h�P������� x*�x"�*Ʈ���7�����"��ړ���ԦU�Fi�a�-v��r4���~�sB�%��{T=���@\�;s��=���)'Y[Ӯ>
tEcu�FKj�l��	�q7\����i�-׹�������Y��H�`��Q�a��j1^��4Trj���"b�5�n��x�%x4�/9VO)�����?��i������F����^r���h�e�UM&�x0�)�3`l�ڝ��s^���*��4����-�a�cn)D�8�&��	�쟽�4n��Z���5��+���������;�؂�&E\btqp�<,s�i������T Wuo��v���4��R�nNQ�~y����%�_{N��6��ld��K��j[u�h5��a,bU�f�$ i+ ʎ�n�R2�|e@��:���1�ۦ��K{V�L���a�ב�$\��3���gO^�y}�7��R�\w��j��q¥-��F�]k7�2an ;T?<Ԋ��WĤskzf���2cٯ�U��^�Q��;�Y����������u�%�������9��f�9Kێ\�#!�|\TJ�l�*=z���P�v�1�[-�Ur㝤��83|�Jї�'���L�G'�����,���:�}��E6�ef�5��NJ�{+n���3*M��X����gv�Ί�������圞
𫟁ޯ�]�iCW������u30�˸���<�[U|���ݸ���\�˵����YᴶP�F{fC~{^�A�(Q�<��8��J�ԕ(g���,���WԀ�*@|�'g�3�d,�k�;]�z�D�N{�ִ��\5�Bچ��Mos��b����Ft���J�����A�KzCN��5��f�,�&��Պ�`Wf�����}��C���mf|v'�7�
��OtT<g.mm��y�;��y�o�����+�R0R�CW<�G:�q�M$�srb������x���4� P+��\{.�dM��,�����Z<�8d۵�x���ȕ���Ivv�vh|�2`��F�l��p����x�q�j��TcQ�:�xT��j)�BAg�E=.p�웧V�}�s+�]WW[�TV+����"Y���着Sp���E�8�{sr)[3�!u	J�h1>���۸9=>`��Ϙ���[�cl�Ԥ�ٶ
Q=���XV���]����|ڤɥ����s�9��z4���}5��!����#��_ ���,�ns��яՉũx�SL�=�K)���7�����3�L���S,{����>{�'^��[��t���еÞ{G6�Q��`��3z�!O�	c����r���w�VEgK��u���z�7�j.�1�kX�9-1ܴ�O��y-3u�fWب��A��¢o�����y+iW��>�߯3~�Z��Y��u���;>���/j�+үxGx��R��x:Xebɔ�^ƽ=���Ö��֗N|�������S}c{c68�k��E�tr�ҩ\alU�koUW�zY�5z�h���p�D�&QR�v�R ��g��hτx*N��R����J/�jc�1�n���s�\,�[}-��yu��Y�94-&���q����U|!�-�)QZ{}W�D7Z��W�"-�-��Ń5�²p�Oz8��l��i�ʊ>�9���������[6B����x ���*�J���X�,��ۃ{ԸD�w8sQ=έ��y��=v�O���I�Rސӽ�p��=y�Ꙕ���UM��i�K(��Kt(t�|�`�?���N3K�?�{��A)�r�#��CL�|��f��z3ic9P����1PR�_=	�^���`;>s1Ξ{ofvJ*��%Zpyr��;ԡݍ���Y�B��ի��jB:��2�x�cr��s=o�W���r�7��v��n&!TZ�~Ѷ|��u9��7$�=A)�իf���h�����i0�q��ȘN��� Ije�y���j���C/�Z��e���f�7V�jz�S=)��klGs_f�t����OC[�����?|�̫��?g�/&�Z�����E�U4K�r�5�<�ͳ�򹟵ٺ�1��ɛ��b�Ԕ����`�W^�S����w+Iĥ**jA���׼�Н���L񕲃eA��u��2�h�'ֻCϟT���ES����"���+W���(���xQ)'x�7�lm�VN؇<z�֨5��KT{�ű�%o�ꓝ`�̆���5�"�ʘ����$�ą#Zr�ES��0�)
�}ەgp�u��q��i]C{'bޠ8��hQ)�ػ*�#��锂�K�����
�%�ej8q�ʊn�Y�g�l�����:�m���q2��D�K!YdZ���j&%e�Uۗy�_P�;�[��0�u�0<ތ��NeLp����W2���y���є+��'�YVЬ�k|�ض�skAu��oZ����Q��őꢓ������Ө�K�c���`X�
���úAȁ+:���^ލ�
����W,�JTꝘe�Ғ�W��_d�v�u��M�n�k�A�T `7�E��Iu��,�0֗�9��%�rInɫ���իQ1�4Q	�:��f�K�U�G&��u��X���Ւ���P���a�l���V.�J\��+��g��c)�A$Y�X�n�h7J����ݮJ���Lɡ:{�C0�M�ۚ�ᐽ�ʵ���v��p`^��!�C�!�+85�5����)�o��\V]vԸ�Q�ObN��HV��I�b��LcT�N�YxhWP�ji�'�����f:ԝ߯�³�j8]�1[~������,=�(X9k�O���VM�A��tcyAZ�P�و"� @��CPI�k��,�0d�j��<�;�|Fܠ�Q����>�=��e�(��8S�i���h�]����R�K+vh��I�CX��{*�<�tZ���h*���1�ֺ�U���b�Q��d;y��<@u�S��F"-[�L�,e������{Q���!�݃�vU�5�C�k����8Mu-fu'�
Ν��#C5SXz��i�}[��6��N��]��w���@�/#*nvjt�:,v�ܠ,�K�-���MWZ>G��(SG������S*���N�7[*�E��,c�tM*�qK��"L5��O��p���˩D��׭w��t;��XJӕ(QW��&��z�@V�[&��9�tz�;��l5�:�س1b�n�A]�i���T��]'Wu��[Wģ�u�4Ѓmg6M^�SY��(5di�g=��狑��H�E�����R����S��nZ���߅A�d���F�Di�/�η����K�f�O�u��x�^�}�C6�hd:K$�����˕�7J/	4֕�D��#�t]�Q�j�W;p�J��Ч���^�M�R��qP�Ro7p���VT��44�n��o�}|��2ȩ��rwLI���B�S����P��u��{C�.�&���ݰ@KX��y{QL���4>+ܐ2�q�B�"�G��|+�*��!�UT;�k��f��PuwH�)ْ�	�"uJ��^���"C.p0�s�-��fYu�H�'��U�	U�IV��J������V�ZA5IY�㗈b�b5n��ih��	�2w]!2��������y�V�����j��U�z��\���52tv�D�ԥaX����aANg�)IGR�������VJ!HQ�77f$dd�s'V��!�(�Y�*S�:�"%f͙ZҲH�a�5FI���"����Y����DDA��3�WJ$1i�KR5L��-k$D6Xu
Ҥ�ʃ�ias%�r:)��yZ�1�*#h�EE��e����(9,�0Y!]hIA!RB9TJEE�t+#@��	fd�P�2�i�i�����r�,��p�RK$$�HдٖTV��Y�*,�j��bR��j(��ZQrSt@�r��'sw10���w	B�k3V�m�L�LOwtBST�)�XI 	&�������������K�Ő�����ͽ��52��|:;���7�+�ӆPfKQ+֙S�V�v:�/]�Ҟ�}U�}�ԛ��!y-:���zwn9=k!���tk��;ƭ��c�7j�<�[$���Bk�3�'�O�k�M������̼��*u���(o�u_S}�4���qYNĨJ𸟯�3p�6/�m���W��pR����.IU���@��U�+N�9N��v�ZM��C�{����Qg�e%��d���q��>A�x�)�ʾ��N���z[�p՞�%�nvה��;��Jz�{ڪ�l�ˆ��A��t���TDKtcs0'N�Ғ����
%|����?}8��+�i�-�6�D
�> �;�����ŽW�;\�4���Ԡާ)q��������r�|()��	S�3R�k�bl-���Z2�1�ݐ��1>�-�aޭ��E|�r̢�yv5a����.�&�.��6��ӽ�r�Q���&���8t�n�ե}���ގ��qVTvV�3kkio�qF��s���m5~�����>o�n��D��km���+l�+8����mEْӌ���������\�Or-�T����ܗFTM��ݹM�Vq2��������ϙ|��W*��uq�s4���G�k�9�꯾���\;=:�I��paը~�	Z�yv��o'Z�Ĺ�&�1Q԰�괄�:!8Zέ&:�F�Tɘ�c`'c�~+rny��Ѽ�����r�T�\�gl�D���f�K���k�mƻ��1��5:᪵ۗ��4��b[�y�@����.K%[)�(^�b��n�ָsO�w8��� �����1
X������͐W�����=ɷ����q�c�;_e�S�,��߸��T�b{��nW��kb�ћ��e�(��|�L�G!>j�K�(��s��'A��r����mU�Χ���Ja\aq6�2�6:ż]���]�}����kk9-���,�Vr��\��u��P�F��0�6&WVUT;��tէ��[��u�{g>Q�@�?��Z��X�]c�a�$�T�C:����U�k/���o��nM�>U�=;k�S��e��^��Xc���
�ٺ���YjJ6�nU�#���ڻ{�F:��y[��[��u���=�c���[u$|\�|�%<2vʖ��ٹ(KMK�Q�j��u1��y�)Wi0�Ŵ�@��C-ƈX�����q�6�%�3�=DG�}r�D�|��6vr��%�5���cг�On�Q�O0:2��\�0:4�-���6@��P�x�:�[�PZy|���6�q�R��q2B3������z7o��mS�է�jstS����n7�:oHj�ۭ�w$k]�7n�>�f
{䡊������b9�ci�I���V�}w������� Ɗ�c�d?��1��R���S騞]��O��ފܱwo�x�ǣi���N��t�ɾٶ�<���Ac�����K��K����ɞ�H���k}S_sLM|��j��tG!�K:�X���L�o��ꠔ=��[�%���#��X�Jno\�+ �bʅ��dP�]QZ{�CF��3�/2����x�ܬw�_-p�T=��i��]Wk�<ʢ��6N=M��Kf�{����@�EV{l�sڎ�p���r�w�Zb���,J�Tr� �d�d?;��e'~�~���������ס{U;i)�<z��֭M YÀB���*��j�o��]��q�z��FS�t�R�4��/'c�t�m�-��I�]Pc@�ѶoZz5:F��sd�U��3�ȳ�}��}_W�H,����_�+B��9�v���#�e���?\Lux�:���V��gk2�֔fο�W1Kŷ�����ݜu<3;c�o��j������3N�mw!f>*}��_rM�t��*�۪���l�=��0O:[����ʞ�%rJ'$���R��4�W��E�k/���uϬ��m�ת���,=O9Jɲ�z� YY?�_N�q]a�o��5�B����M�S��'�]L]��ܶ��\H��`t�p~��T�J�[EԷ��^<�^����T;�.f�7�����r�H���QA&(jJ�1Vu�J|chX���ީκI]�Z�ѩ�+kŜ���(�=�t�`%�Ʀ�n��i����t�@��v�Ŵ���R�0Sl�9fa�
YGgW4��qI��'%p�O�&��wc������5a� ��n&!R<��DQ�T] 4Θ�D�!�t�m>��qQIK�J\���0�����I��]]-���m�m�t��_� ��md��0�8ɮ$�-�]+z ��U���ov��(K��)cLİY�ܶE�Ρ%L�
)J�^X� t��T�(�������+ۚ�M�:n.���殟l�o'���M4�vˍv�A�/%��a�7N�c���k�N�-0�ue�e�sٽյ��mT�|��ה4V��Gh��^�S<��!f��ծܫj4��G�I�Q�ӏ�o�w5 sk�����G�'�Iױ�yp^��p�/����ɛ��b��T�X~����֘�b�{$��E�=O4o)d�����k�LKٲ����G5�	�p'xe�Q9o�%6��{��k�K�<��ݞu�5��������nD�=�aq1|���I�D��1�yl���ݜ���{�y��l�7�� ��F�iBZ��-��-&�>v�V_f�48�*\Q|�'������U06O)�U��}:��JUF�9�onl��,��έP6&��o��I�����@l�>GJO��s�3����4k�5�ڿ:V��*�W�˵Z��r:C�#Y��LQ�<��Vd�״�(�۴��:��Ʋn�VwJ�
鮦�h�R�ٙp��
RB�`��8e�մ��s��*��Q�b����l�b�j�Q���f��ogpZE�F;�
�h^�f���)�����M����5��Sk��E�W����6�m����P�|�<�Q�\Znf�H]�)�{7��o��.9�]�/:3�������x;&�M�Ȝj^�Y���R��gW؟m�m+��V����|�=�׏����t*Վ�{�0`��S���j֜\�V���* ��z�{/���7�r���j��,�@>UA+}5<�j�y:�h�B\�_�d
tgr�Z2ɽ�Z�\����S���Om[����{�j[o��*�b�ri]o[�U5,�%��eO�쉎C��kj ;U<J���ǭ�����E�ó|�[����:����;N�c���]�)ɽ�t|N׳e���+��vlV���H�;�9K녮9��}Gj2�u�53%d�!�ݡT�w.CF��c1ћ[h��-�S/QO_/�����Nf�c��+���=n-�7M��+HR0�̆ �ɤt�J���
����.�{�jŒ�R���\|�o+:K��>�OX��4�Z{�)j��k���U��&��Q�Qz��6&N�:�u�n�v��w$�qȿ����[�oer�o���|/P�Ȃ�`>U=���¿����>f�/xO6��՗w� �ܬ�o���'���>Y\��_�Н�XOq{F����5+N\�UD��1GR�rQ������|�u۷�/l�Rg�<�j���wv�>�����8�w�ʍ@	�2o��}n˄��t����Ҁ������/�P}6�#K�qg���=�v@��qVI��7��ˇ�m|�{pm��P�.�=�'������O��5��r65��C�oM�s��>�8�+�!�w6ޚ;i��v�[��	hѼ�g�gV'Ơ��p��7dXlt<�-Q���s�����As�e_�W�E{���L�-EŞDYc1	ީ�)�]�Z���`m�k�P��P4�o��ۮJ��n��\��P)>Zr���i���8ø���R&~�6b�P:�I����>���*�[jR��x8����'�"�뀦�C}}�̣>K)�s�d�s��E>9�+���ۻ6��TΗEW<Ӭ"m<�LvL�mK�(t���uM�y��u��R�u��s�@���j�͙��@M��|�ck^�����f��_W�_V�1+h�͙�eolޥ���]C}S_sLMBn5�T!{E��Z��XIo�6�����9D�UY���aqjP���I��}SOz�z,�-#a�g;�k�{�l���W�}�K<~{�~2���s<��{��ug`�n�v�9��jk�<������~��OS}��EV{oW�w��y��j�37B�����/�Z�j���Ɏ�7\�eAw?b���e����JZ�c�3զm�s���q��"�
%��mou�:7��fQW � C����(�����5n OG+¡W�[�b�7�c{��������+6Й�i��fmsj@�(�q����K�x[j�m�ｯ��6�K9
x�c��$ǐ�*ps �:x����R����\c����[�542���/ʜj��f�T
�ϊ��I\-��[�_�9pb��8e�ʺ�"*�|[�X�Ej��˷��2�><V
|�N`�"�\���;u�\�.��B9w8#Z.	�<��h�Gι��¹r�ڔ��R�q>�a2vq�ZU�+qL������V����S���� =s���Uԛ�_)���W�_zzb^�=A�����V[o�<��rz��I:���u��-�=X=%�������o\o�!8ͧ��C�f
c��,��]'�SjZB�MX�댽x���
iXw�g��
m��r�t���jdD�t�9ҋ�]8AX�η��x��.i@o�����/���u$k�ܫt�B���{(u��uME���ִ]7�4�a�C.5�
k"d>Z��t�j�^S5ד�y����m_�D��囫1<It��}bNEٍ��u�&�m�K[ձr�[�,���V�s�ja�x_o����d��79;y�Y��}榸�^�=�n}�w�b}~���m���gF�A�\�q�x�6�'�>u���S/n9�kЇ>i��AoZLw� ���{s�A�7���:O8�e��'-��ldg�}�i]�"���5=�V^b�ReD�Ս
�� 'U�]vZ�G}%ci�Vq͵��`�-3���u�UFj�fH�s� �m��4�^��@��~�(�"	���ȆN-�[�,�W+��&�:�he*�;}��Sۓ6*6�����7MG�YN��������LN`�+4�,��興[Yi�I�e�܄�NN�p�F|��)��[{q
�5`����P�]��\��'��lߩ�ѕs�:�']�P���Ҽ-��I���c�+~9�N���~�:��)�v]�'�U��t�g�z�vv+�A^mf��Co����Gtr���\:OnoT@������*��I�މ���/&�%�.�.�S�(�	��Q֞w��zw��ݵA�>��=J��ڹ�s��S��J����u������/�5�����onT�y��o�G�w�LjA�c6HP��d�_b}���w�rJ��|�e� Q�P<�]�6=�ʍr4��f�W=B�}���&��o�Ò�J����:)K��W��2���+fP�ur�b�^��:����^��[[=�gn�9�c�����6�^j���k�7K���5�t%��n'n{W��
Y���~V�B���n�����
�	�po��b77�.�l�v�#0R׳����Κm]�V�	L2̜�H�cx; �x΅wK�2�m`�]kJ��n"�񠟝H<Mr� :�D:7�pC�oi(^�)/��UԪSޑ����tUt.����i��]�tV�:�������L�:CX}ȍjxxZ[�#EJ���,�,v���z�h�n�uǇ#X��v�Z�-�؆������T�/�R������s�N��Z(�F�Jִſ$���-�sZ�iј����Yޗ��Ŵ�%` -�T�O΄i�� Rל�'��"o��b3F�itM�^�=V�LW��{7�!�	������)����݉��g��6��#�}���:��t�6M��5ы��N����:��y�LH����2 ��1F�Ġ��7�IwS�j��p��T|p�2�{v�h��2�>�����.f��Kx�p[�rz)�	�ٻ �
Nc���_wru��6�Y̓of�*��4����>��p�*������Ebg[穒�z:�FG���C���0�8;��3.7�͌f�ܐ=ڶ^��K�%�`9�+�3���\�ז�j��`i[�y�ܔ�Y��ubs ŕ׎����e�v��fl���VkE_^��������u�����|z�īV�J�w��"}no�8ƶ�
�s*Aj��弩'Z�2Du�r�:��y0�T9:�S�u�����m�-A�J����T��k�w|�fLc�� )Ŧ�B�Pk�BwFZ�4�X��B�e���ovܘ���RT8�$�'���d8틽hl���&��HY롪dO6nd�`�r��M	�2�L�5�>�7 �u���O�j�<�vV�_r0ZW�'������'���H[:��6V �o�� ��IT���kT��>�]�糲�����7����gb�F"�igpH�\{����uȸ�%(s��<��DR3�+ެwP�+H�ԥ�{
ҪU�C���)�h
=��b�j��ň*��r*R�����-b�W�P�i�GU5��ٮ	��W�8]·�J�t��Z�m�cvcw��R����s�"��a���]��!�mp��aŊ!zn��H�g[@��������4�KB�����o-��%xt��u{�S�n���9)Y�	�y��Z�3f	�+�QWkN6F<b2bj�e+�Y\���g9dN���4@�N��up��5��_�[���%�$�|���O.��cH�[F<λ�oi�|DFS����qUy�ڙۮJ�Sm��ʴ�w��*v¸�M��ap������wrYh<R
1����s`��n襠��-M�ܛ�\��w\�<�e�]�I
TP�r��V�4B�6��flJ��H3$3H��<���+4���h� ����hQ���&Q�>@��g�ý���<�s�ɔ�.U��#�ݩ�e!h(�UE뜩Ʋd�����fYТ9���R���",+n�x�� ��j(�!��"�H�L��=]g��I��U����Q(Z$%qH��I.�I����R��IR�""B�gMR��ЮQR^�E�#J8�m1�Q��8G�:�!HaD�����ia��*%\�R��ҍ�W0�n8�kT%35"��Rj�Ta��Y"F�D��8�)T�:�Xi��.����ԖR�T��YYE)�a��ځ�h���e��@�(9�"sD�f�$F�ĤJ���*��6&ZUJ`���E�����$¢�*ٵNu�+J���4�I)
GX�D�TST�0�5	k$Q�N�J�D�*����i�Dm8��Y�S����u���f�bAsC�҈$�M2�B�K��&!2d�/ �l���e��K,��W7Z�b����au�T��xzW9+������y���p�F �L ��={��º�A��4r���������fI}	�(ߣV��MB�bi��T���:~���+��{�[�g\�gq��N�Un��U��u�\9P����*5x�����6��l��-9/Kz2��1��ƞ�ZJz#��������з���l��p�g����sP/M��s�� m����/9D�[�je�)��};�V��\۩��t:�w>;���f"՛��3* ���'��Ħ��2b�D�[�*˔m:��S�֡�~��j��(���>�z�;�|�����-mu��5̌�O&[Q{�4��I�P�s�������О��Fbی���uj��cM��z�ĩhlu�k-6��t���V5��l�I���4�ط���>8�f��oj%Ξ����R�Z���cг���S]X��Ш6R֩d��ٻ���y`l�W���Ib��xB�n9�\�^d��D�V���) έ�d�]��FCdݼ�;����.�b^1�+�^���t��y�O���̩��rIe��=a�+h�X9��R�GZ�X�q�����i)A����R]��C��O6�T��Qޮ$�ǫ�-픉���0T�",Ʈ]���"#��Ocx��W��_

{��PKE|7���,�O�o�>|A]���w����Gͥp�%As)�%z�H�j�~&�,�a�V�y�T��{��)�.P�[b�?�{홈D.�)F��)��!9��"v��]�����wZ�n9�����l>G"U"g����r�u��.����ܒ��5t���=���������Mƻ�a���.3���i��G�O9wpb�=5�s���=�a�[ԔZ���{sa�Lڞ����Q�e�-���$z\oY�AE�l���'i�^e�-�t���׮.�z���
�Sw/�����gjΪ5q�d_<���f�X��o94!�|F�E��V�j�[��γӺ�7�_����ד�n��̨.��s�*��z�uYZ�R9��4SaD�[7�TzW�yS��N�(p�� -u癨�z�R���~���lY�й.�D��t�����9ݛn��6�֓���T��t���?�o�d�:mw��o�4���݅_Q
��ӷ��VWs�}V�z'R���Ղ��w:��N�N�,��j�/FAv��r�6�kmWO��U}W��OF�MD��"s)�	P��
�b��{ֽ����&��-A�W$]��pRVOu��bT��AJ�g�}N��Xl8�e��\:��+��t��Ek/xT��s��+;T�ق������+�"���-��8k!9cq�A�\u$6iv%W���c{f��G\G 8(��ԗ-��zgS����ĻrywQi(������k�7�R�q�>�+䘸������ϧ��-�z��{���Xv�s��5�7�Q�D)ﻧ����FV��3�6���YݿUY�ߋߌmu	�;��R��l�Öe�P�hd���鐕��(�]�_]ņq����s�M��n9sP����p��G�Zt*p�ݳ����=hj�갥-�{;#8�N{~֋�o�k���!���p)nAzЧ� �G�ܴlE���<u�gR]�������^KL�7�GJ�j�q�$RB�p�o�w�a������JN�ޡ��l��|��F�;��מ�A��$�4.� �+�.����!��:�&�Y.]���뤜�Ǻ�s'Y^����}�p��仩�x5>�"Rt�:�sPt�U�UOOcYz�jf�ϣsaM&�]�+��vD�"����y��m*3ڭ®���2v�o9@;�7�9�녮�����g��f����;���+���u=K�X^��ZK�R:� �~��z�8�ö��J����D��݆��q�-�A���н�9F[�ЦS`�[��m�j������fU[^r��3�Y:g�߶��]y+Ө�V_>f�&��o`��t�x�h����/�/=?���.=���(�[*E~����OMߎ�.R^��}��/;������Sl��4OJsZ�]-��J�>�ވ׳�lk]��9e�� ��+��g�����^����մ=9/�������f�F�mr{9�]AT�F�֞޸�]�qx�X�7��x��$�T�'���K���6�o�@}���X�[����vR�����x�^zo�Y�A~/5��M��=L�k�e�mc�b��_��L]��cەA-� d�Qo�t�Q�ó��,�������f�)�RÔh��-^������fvq���$>c�nm1aۿ�_�k����L��8T�ئ]�e�͹�q�?���{�2���^��_w`8�j��&��{��i\@w�q=�Z`].�c6jrd����x?T�%��I�Z��~Y�X��?@a�NzL#Fˇ��`��h���f{0S��¾I�W�ٟ�g��R���U�5����P=Vb��G��v{�ҟj�m�w�w�J�L�?�|:��}�m5�W��֔;p�6oeKԶ��wک�Y�M6�]���D[���-���Z�wJF�#�zE+��ء��ҋ~SL�؜^�g�W�0���+S�m��$�ѯ���f:�y�KF��u�X�9K녮9��q���p�j����V�s(��7Q�3* �#1otJї��c-�2�u�50t[nT�.-	W�4_��Ij\�v��d�	�#�;�%0��I��{ՕS�A1@�3N�~��V ��~�i���7��g.j)��W0�D�~��h�/{U{�e�)���f�]�ε��58�k+�wSqw�^lu�6�ɫ&�j�)�Pf�:�:wn��	��s[Y�=ժl{K��z�7gcy�	R����T��{��"&�rKs+y�f�:,� L�ۇ���J-��Y��䊶�O_���'!w�\Ř]��}�1Q�7����n���@l�y�K�ң�M���{[Q;&�����1:W��Qn������l���sё��W���OxPT?�oT��w�u�R���q��z�6��D��cdhN5Od��:�0�����hjJ�Puޚ�-<�x�T�*�wM��ǉU�}��-+ۙO�<�ȯj��&��fy��o*D�2����5�:�(�M΃�a�!ߤC��ɢ�N�W}ˤ���x�>h�{�-@Zr�siXw��9����٘D.��@���L�Pږ�Ժnj\�[��i��{Ϝ�6�;gv�T��aV��%�΋4���^�S�GM�s�M�E���[Q��M�KI���e��<��Sɾoq��b�[�_ymU����=�a�[Ԕ[Ji�'�6T�pe-�
0�*��cRA�J�J�n*��|��ưRF̺�S+��,���Lq�����{iެ����Ы�n��u���]��#ᔤ?��,�8�'�����|0^p�q���ŀ���%�VZw�9MF�R�n��o*gM`���u��u(�QA��=��뎪�*%��;X��?S~H�{��k�c[]ڰ)�E2a��)^���Fy��gB��3�W�th����N��pd����Z�:�z��*^��޵mQ��ד�F��c0:�Z��yy�G}}��R�!j�ͱ;�^|����c����vl�n�W��f�H��5�kCn��p3
��T5ap�#b�&źomWnھu�ٷgfz�k�hm���!ʏ\�:�vY���%z]+��د�CYm��m�qp�t1ST�`K+�?�9{eU06Js�<��/k�*�J��o/L�ε[�SP*��5IA֙�J�����N�ۗm�B��RHpyV��M]t�8a�N�=�M���]�qmx���(���>�+�N����*�%�:B��nu��8�����;}��䯽�8�����S�/��X��.���W:�}�.j�4�W7���nLTh_u9hR�0e�
�J��J gi�{�%�P��I��������y��tEr��W�H!������o���ڝ�k\�Lj�y�q�Af� A�#h������{&���k���Kɥwb�.a�}Bl���?x���1�s�(�,0Sl�9fd��.z�f�mb�K��0J}=+�pM�c㜹�kGxz�w{Ζ���XRW�VoC��Mt5Zf0:rV����;ɯ����9#�o�:�+�s��f
iT�T���^9j�.�v���;䢬ʫ��f���Z#��4��ZN��j��X�MBn5ں�vD�"���ꗙ�zI|\#U�ֻ_�z[���ɾ��_�\9���tuQ��AŮ�/'�ܒK�톥F7�E�s���h���ە��L�����}Gk/9ѩ����^X;�n.��܊Z�|Ϭ�c����=T\�=��
l)z����=`U+eX��o����D���y�쩏5Y��/��SћT����"{!)��k*���ٶ�f��TS�
�U}:��F҄�K������|b୹���hȨ2F�ފ���G(��4pS5e��Ǥux�T�Jm��S�~yزT�:]u��ǎ{��*t���mX����I�-���rDA��y�e(7�<�2&��dG9NQ8&s���ڥټ�:�i*�mk5���r�QJ���[��`{���;o�s�5��r��9����Ş �k�]o[S�����-����e�o���kz�P�@n-^]t�L������J�����t}-�֞tk��ޅ��KE������mUЬ���r65�q��ܷ�7׼����!�A����[���@֚��(9_rW�-7�̀��>΂�V���+Uj�U$5�4�q�N��{~��@�����JW��f�(��X�����3R��C7��������
��E}٘E��R�A[�3�� �.2���Vl�t��^�|֜���[|ƻ��(��6`�"��P����ϥ�}�}�͚Uj[Z����MD,�&�mƻ�Tƻ#�|t��Vꤹ=������k! ���un���$��sP��r�k�X�ST�m
<O]�ޥW��|���ь!*No� O��}pU���}Y���z������Է�F��/%�g�g)��o}�w�qC7n��>�yV�? ��{����7���ДT�ڱDYӼ�h��γ�Ŏ��S'�Z�+1Tځ�n�=o�90}�W2��l���^EeRS�H���R�D����$ρ�t^Q�hy���d�7�̣�`f*3olJї��c-�x:���\�F�h1708��7�ޚ�.Ҽ����|9W�3j�޾��m��=�V	k��j'a�w>7�6.b����>���V���;,'l����6u��$�|��7;�;�alW$޺oS��u��휯����ȡ��L��c9��{��sƣiAu�'J�Kb��5�	��S��֚'"���F2�����Y��{\T��0*��.�¨���o1��qB� e��7&��ĮN�m��C��P�f����TD���O��ݴ����s׍�ݕ�IYq���
0�Cy�Ȁ����t5g���cx�ݡ�u)�e��ް�����F~D.�(`%���N�����7V*:vk�0�����^2�0��B��[�=���g���X�8"�6]���oZ��A+����|[��QT��3�V1L����q�mm3q��@뤕���J���w�� ��)�.�<f]��Wٕ�h��K��ޡ�^N�v���G�mp%J�)Eg<iKz酧,N�3q�R��!<�6�Ǣ�R8&:�캼7l]B`M�s���2m�����r���'	ŧ��a};��NƸѸ�	u�ܣV���BJoJݾ��V�(��!���]H��.�HG��T��xGV�׉f��Q��m �t�b�S �ps�9�������(Ө�y|�@\�x�"��s����0�x.w�ѩټTH8P�* 2kkp^c���kvԆA��[�w
m�S����:t]��yWj�(�T�h�����RN�z���Wl�	֙�ŇlCFk[]Ւ���(���Ӗ�I��^���벀�N���0�1�{C���ȚD�0�f+Q��%�e��ջ�
&��ER�	����G�g���/���pτ�76<a��D� �w��Y�D�R���(���L��9��ʯܥ"������D́�YEͶ�T��)������L�:q��C0M� f,��v+6T�j]Nm8��"��µ��
�q�h��o�MZh9���L�@=37�9�t(��v%�l^�e0l�}��|�>wW��c��}�����T������z�I|^�c��Y�:YS9}�q5{E�õym���iSU'�o�b!Ne�o0z�0ͫ�S�Bfe�+zF� u�*�$����%�ݪ0��O��L53�tE�.�Jjdǔ����t���`�\᝙�S���cQ5j���a�.�Lӳ� M�S��-��
J�7����xDࡼ	��o6^��;�\۱�Y�	�Pͩ+9h���r���IǝC��C�.�&+r;M��MN�EgZ��]�r�u7�p����n�:�ҩMf��-��6v��
N�;ֶ���D90�4�n[��#�8%�ⱌ��_Y�WLN��gk������tQ�r���a:�,ň�E���ŉ�͞�\�'s/[�@;=t-l��l�g@����S|��)nمP,gG�Y�+�nղ�P��%�ʆq]�V(���!^M�ZU���p����֋O+���Gq�tA>�6���F��5������^�4�R�ap��ijf�e��D-����Е�"���-V�29N�{p�0P��uՓ9��tT;���i��\�]������lu�`�K�����e�76��,�:�N�of�Pgfℾ�k�4w���,sS&
vc�dJ�2��w7>`�`��IGwI�T�LcZx��xݼ�s�@Jq�����VW
'hЍ33*x������:Uo-�����9^�iĵ)h'�o8@���I@Th|h@|��K+eAhmHK2�$J��
�4:��E��4�6��AiK*�4٢��%�QQ����gPP�*��+S,奚U"aX�)�THer�gKS�F)�b�IH@"��5�\��#
�E6+1
R���,���b�b����(�X%YV���Ģ��$ɬ3�m,�*��9��Z�"�DQΡH�J���3-H�
-
*���AB�.jQrM��Lª���E&�U�0ӡ@���:&EQZZIT�j �F��­f�[��*�\.���m3"(�"�#�j�ʍ2�;L��H�U&Ur�J�ȹG2ڢZ�Y�3-)L�#�PR��-D9&ͦ$�-,E5�6EYЪ��DIX]�MPͅY�� a�ᐳ"�&�折r�Fr�o�c�E�v�tĆi�&�̾��ٝf_U̼���L�I�Kk��
��7S���xc���9:�|�z|��M+��[�so!�<j��(J�݁B��1/K+es�e�z�s���>9\��o�b�NȕH��Ն���!�Ǔ��I{}�C�o�)��5���S-��k�/��k'�Y&F� ��w��?OA�ձ5޽5jnU��ѴZ{[�;Ub�IԈ��Vazq8�����aŸ������(-���/���U�[��ǚfv�:��y���!,C-�GLN��ߢ��/W��h>��{�mg*����6�諪ՎGouB�/wS6�'��ە�"����j�ׯ'���1�P]����0H��y�G\�n�5t���5�piOO*����>}���ت=?/ ���$�Ū5ŭ���rs�ׇ#V:a��V\5x\*�خI�p齵]�X�Y�^�U���;�܏'�g*�}_p5\N�;*��4Z���>��.),P@�D{=s*4� 5r��ki�ԓ�{,�~�����R�?����OL�_�m�M10�_ݘ�� �ƖW9����zu6��r[/����.�Z �v"8�ZT�N��Wh��Юd]ؖ���\K��F&^J��V�S2�0E��JM���{y�닆��<�e�GO=A(��m�	zD�^!˕���;�F���.�Y=k���7�P(r�pu1���[�Ք��N��j�ӭ�S���E���P�-��q��WO��WG���a?z���.�h�%��g_ҟ-�Xv�S�·��C�f�C��=Z4����o�|:��/m9�_F.�iXw�C���g9źx84�v�g��<�������	�r�.{�7Q��W.j��4z�=#j*�:�Q���;���zE8�q*��7�C{>{6��5����R�>��F{���c[6�\^�
�q��Ș���6`���ne���e�y)�/�e�Un�,���n�MT�,p�7�J�]��vG�����1��|s�
�'Yy=�w�_���������k�^����{G)��:rr�%[�$CfF�U���6�&]�ð�4̭�JLm�z��0��M{_[�Z2啚;fjzO����)��u�����SH<��,�;�JR�Z퉽�,vT$�@��1Kј�rY۷���WV�ܷ[���6��u��l��N�$hJH��ѹ�8�	����T���:����N�ܮw
e�7�ʯ=h�i�X��;�`쵺�\=�ݣ0r�����A�/s�e�}�M��z��u��\�(A�պ��Ť�I�F�Ӱǚ��W�1�+�<&vƍ��Ej����RYx����k*j\�����@�5�e־�ࢵF�s^�7��<�^ָ��*-&��z��=�[1ˁ��v���Xs<�׶�Ҭ�M����s�TbT�7}��޹���@b/���B����֢�{=�xg�痗rϩPu-ѭi�놶�z�<墒76�I!�ڔ�f�= �g׋��D�hjK��o�Ao���]��3Y�y{V��;��39�M�yVSR�@������Y�gV'�I�\��A��$v���)6Q�&���ʽ�̧RR����(�]@g�qm���e>�ա��`L�v���k������o�̛��SD�.[�U�t�;�8�����T�6`u��w>��c��֜Z`��d[���Ra�fpS%�݅�ϵ�B���@�K�ċS��Yb�PsGiLs<2�"b�wby|���dw���F޷v\sB��+�w�W��霄Y�*��-s93�*z�y����,厌ʧ�ʵ���9�m�v�v�ĪD�!� �J(dU�Yj��:u$�s����.�ٽ�����3�9��mƻ�YS�ȓ�Z\2��XJ�%Wt���l>�T�{0��Y�3��$떸g��H�ON�W���rl�8z�C����=�&nx���Z�J{i>�s<�l^��S�����x�x(�v=!�扜��}m��6�`+ڪ�m��SU�����VoK��OjG6u���)��V��.���,��;*���:�3J~~BI2�VEr��܆)㊉�o�R�	�-���Z�=~R�"�ʳg�(u�{}
��J&��e�R��KU��Q�{���7W�Qnެ�,�G̔su�����Pu8*���Q�ઈ��hlS���o�'�.��L��yn*6d���9n������q�K��7��FF\/X�6�NLyzF�}���ue:�v�7�l���ȸą]u�lQ��nQ���G���%�'2I����NL���B���hm%`��m�����zB���I�7g=�ԌDk���{�ⳕL�.@|�vx�����R�_joo\5��S:�j�L�[5��U�q���j���`t�T��@Ԗ)��1[:��
��x-E�Qky��9q�X�2M�ۏ�3B
���T%�c��Ej��+it�������o�����(���L�F���/����k��^��qʎM+�;����اl�"�:�UJ��ٛ���4z���~<������Dc�Ϝ�;����FRܵ��bQ3�a�o���Ѯ�_���}t�f���je�7�5�`����$�[��,�
�cLu: �T|/*����m_�(FOV�B��l������x$��z4��ޡ�4�}~��IIG���v�`���nu�Z���]�Pgsf��ֵÞ��ny�AeS�f��U������[�G���0�D��#.����ro�ܾed���{dچ����m��J��ڞ�>����u�����d������%G�^�"Ay��dtݤ����ݫv�q���v̦kE��}R��H�]�xJlpg"� ��F��*f,]�*��P'�6wR4f؝Cq7�:�AR�OZ�j�Tz�{��s�:�O?m��w��9���逬jϺ�:�(�ڔظ��n[�٪�MR��7&v���,�2�������uV�P�G�\*�b��l9o}�Fc�p�쳑QW�x����[����Щ����f��%F�J���Cc"�!���L_E�y���y�m�^��f.r�y9�P��r�'ݼ��u�t"=Gܧ�.�����<T5�B������T@�܀�*�{�R=����K��os�GmQ>zjO/�5��-�y�*!JU(t��>���ϗ\��!�t�@z����S�E�������m<gF�D�[f�U�ؑ����}�ݿ?��{A�{V��71��4���R�v�z*�b��Rf����YVy2�]BR���}5K���7_c�˚`���5<�Q���gݏ�@^ue���uXd��.�^�Y�̪+�����%d��$q�E��܌���к�A厙�T3��Ϟ+���n�)diů�e��Y�6��tS�b�o`n���Pv�v)�bqw�\�6���*��Q2�� �M�V��Y6r�[�-?����T������-Nʢ�S-'U�^�T�I�2�]��BtE�r ���
��TQ��׹Q范�L��E���#�fW�ޔcE��O\���+E i�i���I`�<�s^�P���鸷�t��������}Ol�q�����٦��5 .QWL��5�����m�GRѷ��nW;�S/y�|�Qٕ�ـ�ff��r��=��Q�(�͖�z��@�j����Qk�ʹ�{���M�w�A�JN6cZb(Qpo,\yO�q߉�v�d���㛌�꼔����!�l>�@��A�Ҋ�=OW1r��Uٶ�oh�E ����'] e���nmw+)G��Q�y=TD���x��}q�{f�'�"�9���̺Oe�a�)�z񣉥����-��+�-�8j��{f��P똚9��+h b*bן�������&�Mj�I{Z���˾X2|��T�k�<b�����4��NX�+��*��3���b�
o�xsmrkn�|8�^+���;'Ap��9HL;�dv���X��Kv��xh��$��>Ф�^ݏ�����d��!��F�Z{z�zt<�5#Q�S�L�x<��Y�^�O�"P��)I�}�K|j ��q����w�j��dWmᶥ*�}�����d+���x[̡}jL�M�zS�v��(������{��x�W�Y@+���@糿D��T&�eP���gR����si\�;Шm�T;fazQ���\w�e��`ΞCu�5/�ƶ�5�Q��K��6�;��k��n'�H���5���_N�nP�٫XR9L�Z�<sk�ŝ�qTjz�SK9�m�>�ej�=y/�R�W,sc]��냗���z�ҙ�go��iM3�����쭭�>�]k_1j�D��� �G����_G�L��/"�L�GO��Һ�X�V����5��(��)O�צ�h��Ae>��J���M{~8����N��*EU�?/���	���V��=w;��]0��:vԳ���k��_'tr�����t|��UaPJ�q4+"����8�>	����Z�ӳ*�L��R)�oc6��7v����=�a�R�R�X�]���ىݤw�	F8v�-��ډ"���ꒂ���C����u��y�y�p���Q����
X:t�dyL?M����ˡ@�ǴN>�0���5<�g>ٗ��_��~>'�q��^w	)�7����r|wm��< N�&|)��+J<FA:7��w3n���L�;���)�����x�R���V#	����/����?[�������d<X��I��B\޿U��}^\g����?W�U_d{|��Z��P������3l�>ʖn�$�}X yK�*}*-eAwM�������"<Eߝ����o�=�/vH[��c�r'=P��F��%T�JU�6z[/5�����P	ؙ�I���#*���}�<�3�#ʈ�7�U#nS��� yMIb`�\��dm�(�V\[t�����g�
�Y��y\M�O�i�~+O��������f��,��Ֆ�ⲷpn,`4yl���ħ|G�]��zW���s�޴j6���`z�����;����z��c�J�xQ�h^W��Ax��|jc�p=D|�	NV��,{ѾW#n���_������;�|�(1F��
n&��������a�ug\��"��ޫ������1AȻ#�n�O��rǙݑ,�꿓f�Z����Π�q��ǣ��ܘgq�M��S�j|7�Y�7��d)��z�b��N�Yi�7��Ͷ^�v�Yd���'\{��:�ǝ�#��-*5�]�\ͤ�ob��(��T�c����^�+TK����K�gܩ��~��+���#Ui7���U���i��Gl�9d3q���RB�OT�|o��-N���~=}�ƊQ��Q{{/��W����Ww�v��+�����'��Y4+�yRF�'� �|n�B��V��U�w���c��~�J��E������^��9�@z��*'�#�t;���l�t�(xȨ�3�m��̟G��Q~����L٩zN��/Ƕ�G�K��'_��^y����+4����`�%3�U=㟆���[��|t�g�C:�VYц�x�͙`Tb���r�^�^�g�=�q���������?W��{�����N��,����P�B��|r:�4׀w���Bo��}ܮ��;y^F�����ד�Vu�<���K�~@ó�g����������q�؇uB����ٮ��b�G��y��~�,�]��&|���c\nω0�}��ʽ�'��j������ʇqE[�/R��}�%wAϰ������xvNW`�*��J��K}�eJ�\�#l����{/#�ES���p޻��6I��sp,�ҭ��!=[r�E�t��uIz_r�Z�p�sP�CZU�>��f�K{���E��rvK���\�l+wU�kt�؉����M��HEV�
�ڕ�V��iP·+���l���.B�A#ԛd��V�F��KZo��0�n��WҲ�z�MB�H/i�������Б����[���˦�e@�p��\/�N�%[KA�����[��~��վ��ejn���b�>����1��B3t����CZC���M� 7P�(�d��$��,��e�����/�4�% k��MH���KJդޣ&�_Z;fo�;m����@>�T:4��}K�6�2��ywV��Z�`�f�YPV(���J�}�Z�#�%3��E[���ޙ\��+
���&�QlC+�y[�X�����ե�)�%A���:������M�쀍tq1��J$�>�6>a�g��j.�ٚE	�M��.�-u�4]��ew(��M%nHT(v\\���v���8�4��x��osT���O�k�;w�j�����2���v�떔us��1[C��^�ŋ�0��L�10��gv�D�Y����\6ƍ�8�u�����!.���\mԆ����V�J�0��G=�����1�SR�����>��߉������{ܖH�K޹�sN%��u�!���)��b�}�p��ӵ��ǳ��x���r�r���7���'���k~!wx���&�oU��qtOm��l���L��-��:�{3�;+��,�`��m;��uPӻv�HlL�0�9�m(�
��ؕ�A�pދ�*�{�;���/��F�J�N��6������
׃��c �~&��&2#��9�n��#���B窴��q�s��c��ue�< +M�U*�X���SϦ��:��.��E��ds�:�k��DZ� �����q�Ӑ��Y�WM㬥���CG���*YD��%N���d�tJ�:wz��j& B�e�%;3B6���Z'+�z�`�{����QvyK����%��`�PsB͚Xz�K|��%�تg�[� K���hͱԀ���.�B�eF�� Օ|�V�-YO�,GᤞW�c;u)�IT���nʙp������ŔWWv7���n��-���i�D�PO��*�������S��X�qV��8��Qpo1˛����ӒI�%�F`֜��I{%��2���d{��5��2�%��fUE[�ֳ���pU�7ִM]��]�N��Q|�.���:',�S�����̌n����Վ�G**t���*F�c^�Y(ݺF����׎e�{Lr,c�X�=5�&W��@��'Z�/���O&�6PO.�M�օ����E��E5�M��r�R��aQ���
i�;�w���BH�4���@�sR�I:F�I�J$��"���-R�E\�.I$E��\�P��H�*�P�����9U$�F�B�˔\��Ud�U�3�Ӆ�IW-։EVdG.JU��bj%r�E�Zd�l�K!2SeT��#.T$���S9Y��*.d�EC��RDFfe��
چHd��T%Jiq`�������I$���hV�#R(��֊b�.�Ҳ�U�*8����4�W�2�%2��5�b)���[R��*4�EI��aE	��3L%(�3R�Q*V�(UԐ�-i�&&�FU��u�*f,�D��2­��L��*��Pӊ����%j���+�*#	D��m�%CL��u��#�e�B�3����D�"Z�E�UZ'��U9e�色�JģHӑQ���8��'V�b�h�mf���v��u�:�w�25�x��ݹ�8Ա�u�ͥ{ �Y'��̳��ړ+��\#)>��G#�si��K���V�V�����>7^�\Mϝ�N/H�|r#�%��j�ni�`�(�zn���xK�w=�;���7��'᎘1�̰��j9�?Rq>��c>>�Z��#O_������>lm�N�s�z�o��ɓ�P���|}DLIo���μ��s�\kV��~v���6w_�ƌ
��#g�ױ���}�q:\�bX%�P*a����+Ԩڹh�������R0=��!sw<	��T����]�<���.|M���JR��/��QQ/��r�Gk�����l�W�䯔E��|i���WF��xdG�x��k@�~ːiK'�%����̦�>��,��o&��9��G�u�g���G?uǳ�wtn��to�{�{!�ب�>ɓJ`q����nH���E���`�@���R�迢�u����묨]��ь}�QY���������և~��h�;�t�������桲���l�C�ŭ�|�fG\v�ǂs�K��T&�R{����6/|{��p��b=�wSf���ۈ3�'t�7>Ӧ�xϵ[ Tny_���P�ڗ��e�Yᙱ���w�B��	6�'B�\]k(��7p�7��r������pL��^
x˳���H���v�9��r)}B��}�75��[�H\�$(s&ꏮ�J��[��.��PT�zS���ܫ�Wқ�k�f�o��]�.�r~v?S��V?U���x_�d$Y9�f>�t���?v�������3L���䢟 =j^Y!�~�����ϧ��³�$�O��A��Y��b�8N=w}�iw'ѷ*g:]C�>�'/�ݾˏx���ʵ~Y/+�dm���kS7G���o}��mT�c9�Lo��]3����jua�W�x�eC���z�G�A��Wg�Ec;�hU?cR��}�d�]A� �X��W�J�t�X��~��z=L_�K;�QW��M�����i��\s�����(���`O���g��9�����>��s���z��{���veΚ~�֌�{x��P�����J�X�(�ʌ�D�뉿�J�{c/,R��52^pӫ��n�� �Z:���}���#o�PeL�5��IzxRvAe�:	���>��.V}TV{�F�q�F���O��ȃ����}�z��2O JG�=쭛��+,a�6}�ܸ����W���r��q�F�W�z���ȟ>��`l9�3 ǧaU#��Ew�zk����\���/%Gq.#>�J:�B���;w�T�W,���[N��l� s+�]�kK�����)K�[}j��$���풰?����s)����<�v�����3����sFtI������0��M7���̙�����I�9���q~)V:�5�x�u��м��S�q���y]ы���4o�z}��nc�|�;���7>>C��Y�j�>�0�D�ɱ����y�Lu���~���ZO�nИU����F��ڟgK��
��T����Y��'tº�n�W:=��ǆ�������y�
��=�/{�zU$_zG�{f����hT/eH��d�^92�������^���}�h_�Z7�D�����j���s����9�u{u���NI�R�ӷ��������:��ۆ�#�/(�G��|jS%'�:1�_�DI^,�w>g���X�8�a�p_K|h�Ņ�z�f����L��e�WS���s��5��W��N������W���е�$z�
S�3��w"������Y�Pe�W��/��I��t�~�4�����7�g��l�mW�`�C�9}ʫa_�mץ�S�N��P�Y�LeW�?r�Q%>�k*�����Dm�W��z�E�Q�|���L�}�_�l{�NL*'�GI�a@S��}]-�#�f��4f؛���W�
�{����a����̼��\i��P;8Ojoc��T��4�xZZ'�7������enǍ�mF�3u��5h��e�N��%�Q��/��R�A���zk��3��0zޖ8��p�{ܵe���)εb�Z]iMu��3�;���<?gtTU������G��|n=��mêa���3��ف~�����q�]통Okez����VF��F�_���O�i����cޝq����fv�,��޺�2�6v�"�zҨbϠܐm�4�,cu�j�n��c����s	��\s����|��^-;�jr�Ϛ]~HȲK����GI}�EW*��
X����^W����g�<p-��@�:Y���P֨���C[.���6�06�L�(h~��
�(��R�~�=��H=�5�k�ޡ��H����w����� ���a�먨�պr6�x�y���e�����;�IBy�����ld/z������~����
ו �K'�0>;�م��i�
$��uns��Fp�+��)��ʍ����9�@z���bw��]
�d�d�|sb��5��U���^ތ��>
���b�U>�t�/���j��.k�X�����w���N�{�}냃��Ͽ{��� �֌��#TL����G�&�,�Ϡүq�X��<Ο��ϧ�~��{��X�9]i(?�,��G�{�n��+�uf�6��\��pSZZr�W����z�3`ꤰo=����Vc��
N_iL���|�ͷ=�'+$���38<@d��V�$�S���s7��3�fT�����X!00�J
+n� `�sk!�d�L*���7-�����4��;���U���s�B��F���^-��~�~��P�cW��3�����l�C�C���&&��p�d���,5�;����tc���sY,ON\��W�+�3�b;Gu��>gs�����R�&�.ʑQE�tԕ�Fz�,q>��(�g�T\j���4�$����#_kwp�W��o�x�ȏu��~����\d��,kF���j3=�m�Kk�!��+*:�M2]O��{������x�9��_�\m��_�!��^���L�,��zo>��GA6���r��):5]o�}OԄ��քZ�z�~����M�N��!�{��ʿD�:���r|iA*�艒�I���8:�z��_�1ܽ���\y����џ:���v{��zwI��q:n=^��fK*�n�Ozz�G\�}�C��d�f3�*k<b;��w���5lzQ>��D{ӀS�q5
Y=_!x�1�_W�����LuϏ�q]�M�z��1^�.���3�fa��Q��n��<k��C5�S� ��(�fW��=��bvw�Ѝ� D�������d�Ωj�7|���C��W�nJտ�t���t�vF��j�ah"J9ks;�L��)9���/H��"��jzo�إV�V���b�֎��3�$�|fn�ҫ6��cp�u�A��W�u�Aet���0ݹN�u�i��#��C��L^T��h�F��������;�/O����P�C~��:��ޣ�#՗3�q�"n�����}<6Ü�������Q�/M뽸Y	��}�Q�l��<}�H�{�F���Ϝ�}��6�%��ꁓ�I���[�'���c��q���n=�����Y�B*3�#t��}~�+ܪS��Rgޘy'�p]���2{��y���J��F�`7�Q��1�%װ�l��L�0}�s+!��o���Q�ʑH�s,�<5}�
����yR����1�Ww1��ב� ��y{$d;��IȯT=6��GdC��_gNI�,���e��
�F
���OA��(��w�v�M������z}^&�N_���Q��uF{�]p�Ӓt(�W�FH��䳖;W�
�&}2�T	�U��WL��o��q�Շ�GW��zG�Ð�>�Y�w��wy�ܘq�O���`�˫��
ϟ���g�L�X���~J�qMՉ���о�G��W�D�Uֺ��t�ݚ޿*��}q��9���F���)zd-��S�O�|$W��s�V���:(7\db�6�R�'+��9�rv;�J�o3�u�M%���)PWb�O[�^��F�4me��>i��</��6�ʗ�vw)�@�-�m�,)J�]�t�3�(���Җ@Np2�Y��)ˮӚd��9�+��!JC-;��s�Iz-E����D5��[�z�����:U
�\�k������Ҽ^�+ݼVUzo�|j�l������ڸ����>��=��\8����o�`�J��F��H�,�L*�#z^����zǢ'g̽��F�֍GZ~������n�G�<f�̓����7���beziE�6��V�&W�®�y���o����y_�߽>D������blO:���u}!��um�N�«�K[3#�QR	�c��g|h])��\����{ʪ�r���.v�Go��w����\us^N:���E�цl	�����8��6��;�V	�>�c�Ӆ\�k�8�Ƿz��_����B�^T��E{�wL+��n�W:=��1��ړ��F�ﭗZ�P��W��/Uy�ޡ�=�bt߲hT/eH��d��fL?V�Qq7�����FO������'N��+��U^�2�1�R��wԻU���a�z�z�
��H��P�0^������,��}�zp����F̸�?+�Ϥ�Mӟ3�ΣyB��?G����u��<���N�N���&�J�%*fY��ӊI"���ޠt�(��d�NsSm�Kxb��-�B}�
�w0&�	�㽶�Y�5�4Sɜ�H��D}��T�X��l����y���Ӳ�:�-�����8�s]�k��$qf�Q��'V{�c�O#�m(2���8�f�7C�r6g��i�x����dz��=���`�0�GEw�"����γ�*3��M��({�,_��^�}n�7��a��}^ �C�sy��/����x�W�u�]�ӛ�Cvxʯ�~���j}4�`�w���@ի���s�����g���� ]�����	Y�À���I��M�Mq>c�f��}�z5]�f��뉿����>^�3���ڪF��|�1����z��SE��Χ)_Nwx{���`�����5�j7��z�#��{O�������#��M3>�T��2<7�EM�{<����Af
�&%:�ll��ujc:!?[f3���l�t��A�w��$z�2kTס~S�dT)��X6����1;լ�A���#o��"����}R`�g�j��=Y�6}3���ӫ�/a��e�]��B���?`M����=��W��j9��{�U��c�ڮ�\6���?O��g��h�~ʐQd�� ��=S/�t��R���̱���vT9���ފ'v��^��	;�L��������裾�lf��w�F�(���V5M��:��lI���54�gU`ާ��Ū������x썖�GqK��iN಻e�(�Ra<l�D�quY���ӂޭ��v�G}��b跼�*�9��f������o�Eד�ѾyLt7�7�=� ����W4+^T�Q,�@����P!�&��y��Ģ�o�v��s�>E#�/��ۋ�~�#��@z��{��{�R3��r{|o�V�;��|��>.X�:=VW�*�����/���ǲ\׸��?Ox����a��_���8���{Ws���F��p�#T�������j�Ό4��8����᎟��Ǆ�qFJ�r�70_P��=�W�To\uf���e=���w#��#�5KF}�1	}�d|�J�s�:��w�������p#е��/��?~�yg\���f�RՅ���@k��3�;����2��vǝF/��`� ׾���{#K��q�|οO��Ǯ���g�Ź.Ꙡ�,�"lzZ�q�w���Ɗ��J�W��ɥ%g��ηU��{NF�G���\>7�:�Y9\� �*Gf8�s/�O���dj�9���I�8��
�i����|TW�Pk��i^#��~�,���W»X�#��^�p�.'���-9���Te�!O����C"5]o�S�!7�Zk��\f&˽YΌ
���4���z;M_����w?�37��$�Wz�ʕ��]"8�F���W5Xz����o�ŕDRx���:�I:+�Y2��43���4Φc�wɇ���.Ⱥd]G��ɪàmc�k<�WfW[�a�I���!sI��^[��Ꙋ�rY����"~��Iz|�d@S��z��
��r"�<3.�_���Qk��m�pL��{����ꉨfK*�n��1?J�u��Z>��#���瞭5�n:z�z�둂��lzQ>p=87����M)d�@2���;1�7��N��u>�Z�M�t}s�z������3QP�W�ߛ�����C5�:��҉�lrX��7[�Q#�������;ۧǧ~��T�v�������{�����to���Ƿa���
�[��ȹ�jZ���S&�|n|6
O�������/N�ʅ����ފ�j�V�F��=�^�>�+�FVQ�Ea�:<K�0�2p7>ӡS�'{�������ƫ�u���ovI�Û��N��G��/�Ubz��P���zY;�f��w��_��\�>�f=8߻���1+R�� os�˭FS�ez#άw��{*F\B�N���xk�>U}���+(����Ve��0����Sȗ�X��{$:/ޒ��Tk��^u�dB��Q�9'n���Ey�b'(����tH�κ���q��g����a.��=�`ջq���e�����4���!v��`6�;���^:[�3C�k+�F�Y�\7L��t�P�-DggRS�h���D/D�����K�;v)r�Y7K+@gC�FR�F/��A��vf��r�ѫ��2��e'��ACj��$S���]0��ǅS��/p6�V�]!-���l
Q�v�"3:�9Ajs��]a�� �	0���4���B����e�Ф���� ��s�St���8�Q,��4�f�g�����\�[�D�V홭��3{�p���o�R"��+��_a��vk�l�Q��	��\�%�����4!��`�c����K"�g���9ǧUv����Y�R���ż��͘u��Ѝ?��RrU!X��V�ǲ��Ԓ���BZ<f�W9�f��-�oF�5 ��U���K3��|$��Uʘ~D�Xi4�]���ʌ1����OU�>�Ih0G�:��&�2\	����m��Vpkb�Cd�X�,ua�x]�8��s8��c�b�Bs�T7W�!۬c좍�]�i����w�f!}Md<w��]���H���E���zX��(s��R5k�^���o]$B���Pƌ��������5�]�����F>�F������Lƴ��;a(��/⊝g�]��F\qԽ4%��!�538�Ԩۓ2t�ę}X���K�{6��r��a;�#�lq&����g�Q_%[��4�dDQgX�(B�0e��ë,/��RǉL!J¥����q������j�o�i�u����l�󵤃)�5�F�y(�;W�]�CTr�ә��X1�S�j��A� �	��>�p��QgE]�4*u])���tkٮ܄��t7 ��l'V�P/��M���_
϶�kn��Ya��W;eV_V��nq�z�� -|�p�ha�'c��9�#�.�Kz�K�Z�S�t�t4*"����Yy%��љj�M�(�t���s�F�������C4#z~	��.��	�I��"V�7&!�
`#�I��Q�m,سbM�\p��k�̭��tF�����t�ww)��˛�p��dM��<�B���	)7�xp7ҒX��Z��r��v��ɯ�ټWPh�gu� ������0M����8��'F��gͥ��w:-+#-����ą�$��g2��ғ���t����1Y�3�=���L���nT=wb�^5��$x]GY}��X�B,�}��<*.���gZ�qEv>T�����t�m>��2���)���K��S1#GuI-�Ր�a\���5���w�.��t6�3�����Y5��1�s�j·���qWܔ�ʗ��R]:�*��V6���2���<���"�H��,bQ��b�9��S��w_f��T\�dp7L�oy�\��x��ݼ�*�HjGNh��B�X�c��=jP��+��4��N�	F�� B �A�fRwu�bY	��"**�$�5+��eZI��Q+���19hc�7hV���U�R�
S,u��9!!̬���mGwT�Ђ�\�f�L��ۆUԲ�SԜ:���j�c�\X�ΈF�z���](.BqE�Y��Թ�D�2�U5�e�FEW��jr��!J�胉�j�!j)DIJXU���M�q��9�&�s̵P��Ȩ�
���춡�(hsTZI���QZs�D�{�Iy�-�R���$��M@ڎ�N:��(Q���∕Fz���+s�HG-!-($�G]�L�k�3]�X��Zn��c*S�������+0����ҳq�j������wS��z皴@�J0��YU�Д�K�u*s��]
N�$�3;�Ї�8�&���]1t��.��yԭ���\T��ᇾN^u�N���r�f�XR����^����Ԃ�%�}s�{h9���wGZQ��Q��U'z���9��ޟW������u���W������I����sU9~I��):+I'�<|&x;����O9,���N#����x�)�}␴���\�T{z��R�Y����s��j�2�Ź �`L@>E���W>9k(�-�	߹��8z��U�YeE����������,������Ê%����~/L���ۜ��u���-QC�f�����	�K�F'��V�ޡ���HN�t����" yQ� �-�K{2��0(��+�66E��>ҳ�Tk7�+�>�A�W��~�MǷ�#o�LM9�������^�s�~��Y>�+V���{L��^>����F�Z5q	��#�����mh7��@��Ӟ3���GD��<=�H�my�<�\}j}�Ϥ���B��M�K�|�F�/+��z|���>��>�Єz[~�'n�@���M�gծk�kfdz��3�`���xи�t��G*|o��G�=�wF-e@t���v�����Z�3��4w
���Z�O��4�'������lV����c���&�_��T�2$�Ǧ1H�zS���4�5�����AԂ�Sf�7ݑ�+U8����u����:F!N6��
�q�om��̬׍�
�D�0����1����5��IDs��lёk����m� f�*��GdH�������sx����ݘ���Y����=�Sp�>�
�P��yR�O�3^�����~��)�]c|�>˿��Sqx߶�i�=����ϸ�}�4��i����{>�uSo�q�Rߌ�9�ˏ��r9l�џҸ~�0���04�{��m_���k�~���wQ;{���Ӓr�����lt*����C��'l��
�.��+ģq�.F?;��������=����xz9tL��h�������j:��Ns�Xr�[�I��GP�'��>�i���;��z=c-���q�-B��?R�����+h�����?K,Z�g��uW��9���a���Q>�759�[=���7cen[=���T<���ʇ�d�1���ё�=?��;2^nƻ�j]^��Ie��Ձ}���;��_����9���V.J4�$�3f���0�{�uyD�Ps����p|n��;���^��=��j�Ω�`�*D.�<��=�íUM�o=h��>�N	8�}�ֺ����>��r�<W�ޓ���둧#ns��{����6�����i:��;��V�7Eq�jI�NX��f�a�.��]�CF�] ��Deq���cUv����M�\����7���+�W`��4�i�J���U8w
Y�ѮL��p�Mر3���2�(T&�;S�9F�T�K���8H,��2�'�Dķ\�������7�!�/�ٌ���l��
'o��zm��^z�畓����u^2+�2Z�50�t��%yM��x��>��+��/vu��ڇ�u�i8�Fא�莖�����K���P�ԁJY1���_�L4�^��7Yk��h�<�U3ֽ/gw&��+����\�.��7>'����C7*!�*A��K'�����Q]���!燺u#��4}H��S=Y�p��?u�g�����P���i�yV*;�RB��n���u�i��i=u�YB��_�}��Y�
��1��.��B~�G!��R��eD�ǲ�)GI;�(5'ho�Ζ{��z:xjK
4�}�ᶮ��;���vڸ�f}���]��я)�s��tg�\��~�՚j<_��G��ۉ������j�΁*�����q��9��t�6=��&'�����Z�f���L���i�w��	X�q��ȱt���A�@yՑ8cc��ϗ�J�
��ԯ��t�^�-��;�;�<��3��'ܾ3�"�Jr*ؽ��ws�G(E��l씅����+~��$W�F��h�۬��"�$�6�� ��5� ݒ%��:�n�Ju�}�6��,殕-����gVF"�UɅ��Xuެ��S3ۮPt
k��$y`��7"��mc�����(�]�&��h���?�O荵@'�]؇�}�"��z{}��垻Còn�W˲�mܲO�]�7=�r<�@[J���y>�9Q�^��*��,�kwp�8���7�<^����S��^���mշnD�ت�gzW4K�l�$��g�HJ������}S>3�M	�w���x���J;/5u�v��ٚn���g<}`�_B��D`B+�pt�X�w[�^�!7�Z){ʏ���{5�e�W��ٞ��i�r����{���S0�\�iA*����-��pzW��:�����x�*�h��I^���ԇ����~��}���>�z�k�fK* ��c�z���b�y;�]�eE��B�QY1������������8�Q(�{�!� �I����M�)$�2=�J��zy�������31��z���� }�5�{>f�
wNL��(��y��֪I ��3�B6t஌�L��/���\{�uT^�4}�z��u�q�~�B/�orc���G�VL�s>����\@��wR�踭}~�wS�q����~�ѕ��(� '�n���	�)�<�oΔf���A��Ox!a�bɏ��v<��U�6j��غ���fe��x	��E��2`�e�9�N����K|ze�t�F4�n�wK�)���Z���+�t]-�2��D�WbRKɷ� �e��핊WS���r躷D7���r�\�5�B|��!����}g��&�����T�N��n���<��'j�M�'��A^.���S�� ��RY�Լ^ǕX�ٱ!z�l�F�N���^���wY~㆗���?x���]gur�@�B����x'U��g~~������:/�2-)d�������g�}W�}��FO/(��w��ۿ�R�/D�я��#!ܿzNG��_N|���+�Ft��s����}��a5[��C�N�D��F]B�uRw�}���>�����n�����{ǽ]Q��Ѫ+����;�3�v�s�c��$�OlL��<�Uzf.+�n5��<�>�y�/O�2�[���ج�u�W����~��)��#�e��8���'G�z�L��G��{�zQ�*���H����O���S�{����;�vA��J8��*��`�2.KnV�מ�ɝ;���q���������O��r0��HN��N����B"�, �JY���w�QbƍwX_%�+�O�΢��"��\M�>���|��N�'��T����9���ی"��5�W.(��������8����
�5�-�}g.�|gB��Y�H�Y�"�s
nGdT�;��w�s^8��������]���=xƦ�ɇ�ut�4m���bo��d�D�6������I�߀�	Y��P��d��$���Y�K����c�dY/��
�����E}Ѩ�O���>��������n�^a��_�g'�FJ���t�2O��5=�8��K�!W��á���#Q�ʽE{��O���;K�u�"�����~�M`��3"��30�p`�s�4/-��Y��������Uy�X�<X�f�I�?M�z4{��kއZQ�Pd�D�}b}�*%��Z��n�X7���8����CY��w��ކ2�wB��������z�V
�,�hɇ�����4�榺�O������,���{ŭ����}����ϸ�ޡ�K#�x'����{*F^�'w��6RwPLm�&ҏ=�����;�sYm�S�'Nj��vڿ�U^�2�1�R��ۈܽ�����֦(�:��R���'}�E�,��D1�k�h����~(9�����C�~>'+Ӭ�;������1�Y��ώ�9��q�+&t&Nؙc*�=>�àӡ�9�>����=^��7��U�i�U��t��j�!�#�LkK'�J+�*����/�x�����_�� {�t���r���#%lͷ��}|����ҩ��\�T�6<��{���6�n�P���=i��U��6�X��ձ��+�y���ՆPv�ղ�ad����t���P��pס�)��3m[�E�8q�uy�]�]��-#��F�k�dr����DqT��=Ln{���=���]�(�I�d3��c�6A�s�%���'����0���ۘ=��,C��z�f�'��}�_����9��E�|�$������73֧uc��=Ʋ��SE몃⾯{�&�|��s��s��!�Q�R5̰���	��.ieХ������Hvj$�>�x��k]X�s�~Wq>��r�<W�zN���m� ��"w{6n�e[��k�k� ��(!Q>�s���~,n�:�ƵHvD�[f+rä���<)/6o74|��O1 =��X�~��$S�-M���㤌�����'KǷ�����������Z�N��W}E�zgY/#ƣ`TC�RDB�OA0��{TD��Qx#��m��3Я7���T泧�֪C�Uy��>����n4T?eH5
Y=_!����{(�ʗf��öV��3��X}�>���������2=�WF�{���x>O*�z�A0�1,����}Xu$��z�a���a�/K���onD'�_z@�t��vTO|l4��t2��?�&��R���Ѣ	4�*�c�t2���j�V�z�xt֋U����L_0g�:b�KV�>�EC�����^�l4o�>ebfঊ9�Qn&0m� ���"/+ORR�fV�Â�;�nj������t�j����nb�N9	��C��n	�/����=���h��+:�exmº|O��~7�j�ř��:װ=7<���1q��_���7�����z�Vi�|��G�gng��@���"j�΁*����3�l��\��5W�'��͟G|���9^�g�ޫ	������!��K�W��y�_l[�dMl���;�w����,��4���z׌��o��}S�u<7K��£;*tݖO���xin�p��Q=�Oy5���V�ܗN@mq�؇�ޢ����޹��?]��&+p?�cC{k���n��i���ۛ;�Z��L�D���Y�JO�L��7U	����9����"7�򜈯:��a��gӆ&擲�u�c Q7�>���?*�q]M������W�V&���r;�<_,�(��؜�˚ݿ:�񲼷��9��P(��A�"�g>-�5�犯z����c�>D߅��e<�n/��^A�Ը�;�4�����f%�������K}$Y�^s�3
յw
��e��r��ɫC�D����>ζ;~~��}���=��D�K+`�<Lg�XH]~�@HΩ?Zo���V9���q�ԛ�@N�ʚ������e���w�����xO�׳�0������.P�R�	9F�].���[�/��%���L.��aۺJ��R��Aw��5,2��F���X2���EM��i�(�&����Ud�ta�g���'�0n����tF������G;ֲF�O���>�"}�=8>�� ��z�j��^�Ĭ��N��ح�䇐�>��A^�Qȥ>W����j6�~�oޤ�<k��C5�l�	���"i�D�SL�\��8�5>�������פ}�j-�c~2
�/���\{!���x�5po�8��I��RE��1,����(�*vKp=8�JӢ�+__��u>7����<��Y��2�$,���Q���Gr����=~���ٛ9����o�kC����
�q=�����/l"f��CխA��+�b�ydgϽK��X���){*pޖ7l�/T	�0��qϐY����z�-'Շ�k�����<��W�����^/�hn���g��e�d��vx�2݌"Ď>C=�ֺ=���B�mW5>�/#MxX���1ܿzNz�5���,p{�/��h =�W�]�핗荲��΁�֫�7�ܨ^�`r���)�u0����P `y�{�����G?{/�y#���"Lt�����q��Tne�~�	��x�Y��-������}���§���͓r.W�*�?{��/E$v�dm�T�a�S�����SoM?[��WW���yV;���k�������EJoP��uhL��٠�6�
@,��C�ף�L��i׮R9h΁0!it�A���޹�G�%�T���g�oO�W��{A�)�(����X�b⺕ώE���~�}�$]փ���:Ѯv'�o+C�G8�1��,Ｊ�l����B>$����$�25q��r��&�sl\��%!���F��.}��#�|�z2�����P���'MçP��f�<��w���������kG� �wL������j:��%}>��2���k�p�n=��~�b^��R��ތ]�Y���"��@�4\�_���-k��h�u�~��Nq����փtG8bf(Ǚ�Yۿ~����s�ә%�pj3�&"_�B�KGF�/��o����^���/�zbs��ʾH�{t�>���%c5�T9�3"�E���3Ц�}.{ƅ�n�ȎT��v���U�Ǻ�/������H�Gj���o�h�?O�w�!ց1��2J��0���}�މ�*c���Y���
���s�����]�c��{����|'�ؑ�kʐt�?*���9��#���Gߌ�����j�n��|���m��bu^E��x�8�N�
�3�?"mm}^~�?"��n��5�%��X�뻸�pĵ�'�J}1��ͫ+�V����J�hf�`�DP��;7K��H�j�vfJ�g;���"#,^�Cpb��9�rzC��i�6T�n���W��Qf��MT'�P&�̛jřm�arX��7�R֓{��:�R�V9�EH��$��Mm�[�x��#��*M��E��]$�!9��pU�73f��Q�M_Ev�q^+L��9�;殹ٵ�P|�gk�⽎v��Y��A�\���Sïo��*,�����S�W.\[H՚���tΏ˰�S�wɋĲ�]2X��A�.�W7FGb�Q��*3ܮU��V�H��9yh�,�1\5;���F�{����,To�t��1W]�k�K0^卷ʠ��{d�q��t��$#)<��-��r��]:�I�t�Ұ��) ��d�Vv�g�NS`�i�F:��[�i7�N�9R�a�z�j�:���t��c.�����>�CѾ��'�'�Ƣyb�7V�ނڧa�J�N�O�/ne�اk9���ӽ��ͨ��F�CUkv4��2�l�����^e�]���#��1ԝu�ҩ�Y�9�(���S����i��s�(<=���]K2ZP�	�9(�:C��Z�l�.9j��x����b��|�e:��� ��Du��u��6�;m��t/8gl=����N��8�k�R�f3'�z�Bqjcm�2�i�I}hm�ʝ 4��3#z3�Z𓨔���FU�����f�+G����+��#��\��F���Վ�������uµ�y���hS�����q�.1j	�R�6t�����֣v�V�7�����Vŝ���i�f��u+��:sa����AGw����j�>Dm+1�j{3v��j�5�j�[��to���7Z��@]�z��w,{��];��0��[��Nv��`�fSgf0�N�u�råJ����.��w>��z�:��$:xa��z7#���n.�ed����ԥϤC@l_Qp]��O�p���ӉѺ�ÊVƶu�B��Dx&����Ԋ�����`�ʽ��'Z5�|�j��mʜWW �K��is˗��T��-���[��μ�M@��~�!�RI��ۆ����j�$n�+xoQ�D��R���Y�HȤ�Mh�]�)eu�;ٱm�nc��'p�J�W*}�fAngU�z�W0gZ��tR��N�Ȧk�l)�G���d���F���fi�1�̢�CoZ�D:���&o�e�8�v��0f�c���<�����K]p%\����z��1r��s�]�M�ŵ�]��L���V�YE�����G�i�Y;;c�"+��w�Z;e�+��#�75@��ȁ�����#u�Q�;oћ� �ţQ˦�����G�(oT(������`����c�*�q���*V������!ow��G�nB9'��b��|��5M#̳�v��AR����.���GѺoU��:F]��c�Q��o ��,�v�K� �+�J�y��:��q����-EsJwSӚ�#��Xd�BEji���gUW:zJ*C�9�w/I-3JP�wJp���\��*��͔�X���^T��NI�ES��EL��%Z�Ĉ�j�)�EzN��-	$��ڙ�jE��E^�r����f�u��%�P�9��K������eȲLwwi��J��D���2UE�nN�Ĕ#�k�]Oqwu��i��*p�68TQ蛺������;Bp��tEP��D������uZ��w<�wO:�R�����stY�y�wU=7(�r��\�u܈��7LD�ДGtsԎEz������u���NZr,�1�uu��͋��F�EU�G"��GizlH��GL�"�ZNR���9:T�z��N"���yܜ�%V��H��'s����s���N�AA:����Q!u�6Z���-u��NsY�j�<)�_M;e�)�*���aȭ]�f9���{�ku����O~�����G�k/��|N��/����c��s�~��)q�u�N��w�^w��]~�Z���F)�58��.|}C���t�T��>�U��*�~W�1�??��Q�����g���M�C�㘯��� ����s�]z��4�y�F��7^��>>��bh����HIFk�}���9�x�;W��YP�L�l�~UC��������n;4�b��1��I�ez8����K�.1ǩ�����+�({����e��$�|f���`ٱ�Ꝟ�(��M̩����.鼱��FDo�|��G��}q�[�NOb䣘�f�����^��Gu�C�I~3 5,�����wp|g����iϡzG���HzW�T��2˽t��Хt2�]����ʇ SRX���x��j5ՍF_�D��z�9Ӟ+�z���P�>�s[��W��^�o\��4��9�Y�����2�p7:_��Σq�R�P� ��BDϻ�.�l$��Z`m�r,��}��'�#�^2%��S��&J�����j|�V����N�F�^�ylL>e��B���'F�)��w1��:EL���^��-�\�����6O*۶�+7�J[��sQT�uO�h�NW1'��j�9�t����^�9��Iq��\���pR�B�04���vv���q�:Z����R���]ݹԵ@���M\���~dz|���N�^G�F@�n�
�,��a{>�bc���j�eR;R��������鬎�1��;��q�+�n�O�#�|{!���R)d��Q��w�MK���G��>=�/պr6�3��P������3�y�ѷ��?W���sCj9O��ܲuf��zuW��zA�N���p{���
�պgK��))|o���g���}�ԥĤ�V��v%�jӮ%eԏ2�g/g����a\@��6�]>'�}�/���ǽPa�o�uo���v��>s���Cܪ���UD��.>g�3���'���6t;�j�Ό�ү��	��?k1�w�<����J'��;��LW�Y�����uo�\ΝE��fa�@�"�N����d<B�h�K�0���*<�L
�~��#�_��O�u���/�³��M�d�N�n��y�/�׺^0��uz�!��Y��3�ǚ����<��Y�_�=��,�]���J�	dW����J^��Zmm���s�Βx�$�hʨw�tפ�S �ѭ���>�iϣ}#��F���SYX z<�p�~.�x����6�U�/��V�ȶ{i��ej�|���3���O��l��
Z�C��I���x�/�o�Ax옓��UujҧG��R��GY��^.ţ��2�� l�U�mU�/�sX�U�3�tf�nB��ɺ�oR���R�Æe�dnsm�%�����蜤���!K���`H�w]M���S�q^�X���;�V^�ufs���eH�����=�t��J=oU��3���P@�,	
W����s��$]���}&���W�Iޭ<���;�z������Lÿ��f�A*�>�o��S��z�K�G�Ē��;�C��޴8y�״���������t�z�Q5̖U� 7��Բ����zp���O��+%Qtu������d��~v����Ӂ�q�z���z�o�=j#���y7��C�
�����'|��&5��&��-���56��n�Hg�x��)�u+d{׉d��i�z漀��3N|O
���*pTK��YR�v�r�����=��;�9]Y�*�j���u�f�ۤ��R��݊��5�)�T��:ǧ��Zt\V��Z��F�?�#����~�9�ؓ����;�c>}�QY����5���p�id�0�[�����N�n3�ႏ��+��B��3k�K�/R���ᐝydd>�/�Ubz��P���q�����{FK��P�"�u�����2�^H֓T}�u�Ȉ�Iӛ���e����W��5�yEÎ���Y@Sf)��\�����U6j��<� ÷RM7CkY�}�8�ԑC ����P0#��d��{�u��;A�`E��7M�l
x���F��v�J=�c}��Zg:�w#U�_ny_�C���2�=�yՎ��xv{*FL�b��+7�,l�OV�%�C�N��a�9YU�I~%8�^ V?/d��ܿzNG��_J���('"� ��ڡU��}���{�͜���\�Xۙxj�B���ܛ��p<�GO�i�x��������5�s/|=�\�	Lq�ۜ�k�xW�\�G^k�,���@>'��Y2�dϦc�̲���=�a�)�����W�;�4�C���g��{��;�=����q�#�9>>��Lm^�-�2h5h�mD׋>�J�Oy׆�ޏS���_��=�ߌ>%GĔ ��-ӧ���͛BW��S���9:��������"��ף>^��+{�4���'MçP��ff���zni�g2"Rɫ۪Ȭ�G��� c�N�x��1����q7�,C �+����p�o�ꑦ⃮K��9ٽ�~��{�'�l���"3G�Dķ\�:Z>�f�Q�֍G_П���Ӝ}�i�Ojv�Ӓ�}y=�ݽzÜ�I-�Rٿ�I�HU�*h�퀥����}��ڥ.����'�k����+�.��k.Va�[PE�{U������چ��Lx~<��6zm�ˣ�w�����#]�W0�|�6]X�����E8T��^>yُqb��
��P��˽����[!���]*�����͔����).e#�(n�w�I�1g�n�.1P�)H:~�?'��x���f�
�͹�3Ӱfaz�*�_K��q��q�.���ok];y>W�_(�ul�^��wF���O���u�OO�p�82;vJ�m�X�!S�/�OH�Z��w���W*|o�|5G;�c~����J�~�	��V
�����d�=����5�xϞ�c��@��u��7
����J�8_ݷ���yޑ�\�ׂx߲h(�y�Z%��o�,�r3�<N���ӻP��y�R��:��ܮ�C��s����4`F�|��x&w���}���C7sӕ-�Ȳ��Ůb0�!���Ip;���~j��gqH���G���+�H�>��um�o/�o��gB�8sfX�A(:����E���^�^�k�W�B{Y�K&y(�ý�Wp�O���z��=��\wc�F+���A���c(�u��"��#�܆�\�m�����>���#zX��W�W�P�#7�*!vT�qe�{B�q6���,�e%k'�=O��W	��J�W0\�t!p��D���IW�l{�D��M��gLx>9�~=v�eA�Jg]L�Y4�%`���j�[�*���<��i�����]j�t5�-��ancK�)�ꔖ+��J������2ģ��\�{�^) u����o1��(r�����6�'��[3��&����Zf���m�=�ٓrE��ZQ*lo���Hڡ��)S멲��A�Q^�\M��ߴ�/H��k��~`K����~^g�� YC��:=!��xz��U|��$1p[����ucQϩ�\MϽif�{�2�N8Lᥕ{�g�����p���m��f�̂�(!_D����끸/ō�qg�"��+a?j��;��r{��S��_Se�};�߽��L��d�Ҡ��w������g�c��}s�h^���H�iAz7��m�&���>��ӌ���Q�9�d�	�^��G��3s]6Yi�=�Ǣ{���<�k��1��;��~�q����<g�w����� ܯqsrm�>�)�K� ��m���z�+�x=okȮ~���y��{��~���`q��:��c�<��=��2
(��p>7g��V鿢�_#�K�q�{p�?]�c���%�B2�ny�]l�>�쨞��C��f��|T���Ⲽ5T�'OwK��Gvi�����j��s|�6}�Mw~���U��f�g�3����ۉ�ѧC٪�:+�C��ý�r��&c0��^.�����Y%�lx�O��]�Z�:�v�+]�s�jWOz/mđƜD&�K��.���9j�*m���u��q�SU)o�ډ03%A{���zINji%v
ކ�'Z�%���i��Ý�G�w���4^���h��pgz�|��Ʋ<2S�x��W2�ޫ!pT�����_^j��S3϶�is��\�:���{W�i����ּd:~��u��wHw����ʝ3kӎ-E���c��ᦱI7@³�.����ɾ�P�]�y}�"�1�����^Y�����GΧ׾��˝�R�{_)�5��C��4��`.��a����Ɲ�C7��<�>�iϷ�<^�L��D�^ź�ɮ����g���'+���H�I�Xʡ�uSs�<�������+��ww9�ݱ}�׹5!�#�%��j�|���QP ��,	�)^3c���z	��L��|�):w�{R�~�e)�>�������=�0�������Lø%�P@J�>�r�'�$n*������H��ԧt9Ю#_�>�3���c�����o�'M�z�Q,�}�A%	�U�\]v���_�N��F�:�"�`:�w�H�i��ޔO�|=87��@��K=�#)ó��\�Xr����O�&Tʰds6zH/��r��z����31��z����R��=
�\j���1�nr�j���m،��q�j��t�s��-5��^7�6�h56�(O�m�%	H�N����I�H�uust�4������;�LW-��h�ԭ�I7c[r�X�w)Pƞt�ǂ*�ڷJ��.�P�]a��\شj(C�ws����)�zL��|O
3/�#c%�h�˥��s��7��q��}�Z����vuH���3k�Gݲ�4o���Ϟ݊��4�R0��=8���V��ɼ���㾾���e����ܯnB��чމ�q�=q��5^á��0Ս�o�\ה\�{ݺ(�io����֩���^����זC�H�J~Ubz�k뙳�id�O��eW�{H���G<��v�Nx�\�Z�k���j� ��+�s>�fS�/�yՎ��<�ݙ@���F}C}�B��H�B�N�0솦<�m�5/ļ�5�?/\�Ey��z�5���>�� O�qy��O����|�Vt䝻�Kq2���z�\Wz�M�\�g>�� �z|H��YLn�����q^���w�=���:��{-
Μ����rI�P�	��f~&�E��_���r�xc'DJ��%~�\�w�w�8�@�c�������g��{��;�F��� �`"������d�F;��7��0ߧ�m���άM�?_��G��ȏuz���ǻ�;��|�K��S}�P�*��*"���K��IM�Z�^����I(�I�<�� ��/h�YL���:3��� A��%�����z��\�veL�}QMܭ� (��Lf}+�:\�W�Wmc]�(�vux��Ԟ�Ԅ��mN�]N����ڂs��9�{7ͭr��@���>���k���{8H��|�z1{k̭��=q�'MçP�~~ ;~�B�z�w�>�"�< ��u��ǥx���5�~Ws�,C���k�p�R�� Z�����V�u�y�⛶����xMzd�isG�Dķ\�:Z>�&1Ѩ�O��~�R�v���;YW���=��{kA�oנ_�<f��-%��zH���B�KGF�R�}B���ƀ2�E���ީ��~�����ȟ�'��k �7�u��'TR��t9�uK�~,z󴵦��ٴ����e�{P��3^�t��{�#��+�1/?Y�p�>��ϝh>�$��큓��E��p�`�N|�KT{Q����}^�}�����^��羠�m�|���B��H3��q'%T
�n�"=L���{������z�M��q�؄�Å�m��d'U�s�ޡ�K#�x'���l��I�U�J��g��ȯH�nT��(��p{���C���#�j_�Q~.;m_�:��9�T|a�]#��ta�3�R�7ގ�?�,������Ő�?�h�C����T�]��R�J92�t}M��*��=yL�#Y\Fy��j]��j�6���p��h��z�e <%?t[��w6�܁gvO��װ,X���%P����e��m�e�JL�5s����:��"
f9@�f0ghe�
��$v�Ǽ�\̝��Qp��{�)��f��k��*15�$�V~w�����N���{��*�8=s:5zN���c ����	w���v�����D���쟭��e������'O��箽���\wd<|+xt*C�~�@�߽�A����f���Q<��z�Л��*��W�������!c�S��{�g���Ϡ��]�(�F��,b��M�m��L��=5z����S��YP]�M�x��z3��O�܏u�����q�b0�cG��}7�s�����'}>$�3�<������������n'���!zG��vM��^���ӽ��sʯ<E����mǪ��d�R ����x-��hb*����ʿ����sЯ�i+^\|zs����W��#n=4̲Ag���Q��s���X��ؚa��}h[�g�j��gК�8��ه������wI�{����_9���A��㤇Q��ٿIXC�H{[����m��=�������A���|����je�=������2�n{rnF���=lNY���7E��ޘn5��ŷU"�iS%�3,��Q�~���o��6��6�����������6m����1��]��cm����cm�6�����������6�����������퍃o�c`���6ލ��cm��c`���m��o��6��6m����1��n��1���6��1AY&SYj5B�D�ـ`P��3'� bF{㞀I**�H**��RR��E!J�
��UU@��!@())$�PU$��"D��$U
BP>�J$RJ���T�]b�*�Q:h%�!������D hjD�0���T���l4IJ�*��E� �%W�(QT��
ID"��HP��E
H�UBJH�����$!UA$��ZUP�X�@��YPP:Q<  ��v�Z�X ::a�s�ݺ:2,r�
wY�80;�t�V�t�P�]Z���N'R���*��-GNV�u�չ�5&�UB� ]`R�/   l�k��.�uJ굚�ݸճ:�����c���:(�Eݪ�  P �X�:4Q@Qn5pQEQ�8��4  =@[��@ �th;�I����T!�  �p K�fx��k[Iꓺګ[��R��kv���A��ۻZc�7v�d֦w,q�Q��B�Zݎ��ӧZ��e
���*����	K�  ý%BT��۸GwYs�Ьw':�0�N�+�7[�]�YvEmM��qm@`#V�]��n��ۡ�U�;�V���C�����!*�t�  Q{j�[b���Lv�Z��+�ttwA�����gZ�-�wR��
Wm��ei]��(�uN�κ�m��kN��-�B�PS�TR B�D��J*$�  <�i�u��[��wc�ۭ��2��\:�4�k.ۭ���m��:�7m5���7*n��9��[v()]�v�E.���)]R�KT ��"�E	   ���mJW�5�� �Ҙ(5�;��F���Ό�
SWm�u�ht�I�@4[GE��4kls��wv�C���K

�R��HQ[e ��(�kT���  �w�@�ݺ�w!ˍ�R:��KhR�kmNݲ��w$��m�vZ�p��&�t�k`ӣ\��.�F���e1���[d�����hv��R&�T�]�)�H�  ���M�Gvػ�Hj��V
 �[m�wWMP�թ�9uN��m�����䝮�ЪC��ۻl�u ���f�ivѡMȩ@*UE"�TTU^  ��{ڜ�H��.�ڻ��0 r8�[[cm�@�R�[�]*�۴9� �@u�SwgT�n��6�B�`uEi��5�i�w���&eRU@24 �{FR�  )�="j  ���R�h ����5US�@  �J��2�MB ѓ�,U��3)���U@f`�n�M	�����/��z�����<޷	!I�؄��$�H@$$?�B��IO�BH@�$��HHy�;�w���/������2`��m�ur͊"����%ǟ9Ma��`�'���97Wt0S�j�#LBcUl��`hc+E0�e9bf�0�R��X��n��E`��q՝{2�6��"Y��k$pnc#3.L�����j�~�vj��x�	Y6Ƚ;G&ʣ�R�v�oTLTӧ"�� �YF)�l�y���iݸ�c`�&�J��hm�M�L�2�#��e�U�#j��2�;qdl�2�][�j�X�H ��V$ơ ��T�w��1�ӕ��˺�?�촶��ʙa���DL��ђKf� !�љV\jV�S��Xto2�#��"jͳm�.�vf�ݫR�R16@Mݴ��#W�E���bb�K�m3�2��w�w.Dd�v����ǈ&]�ee�pH��F3���]�nU�e� �W	�C�/Zl*&�q�]�6pJ�!�+/[�����&M�6�I�7V�����=7�Q.��=���4]:b(�A٦���� ���6�G2���uop[��ɗ4-O���$�^�9%�{tbs�o\1mAgs4"7Q��!�N����T�]ʹ�^Ҽ,�,�R0��V��Ԧ�x)�ںu	.�Z" ��pU�
n6l�4K(3�f�Wj���:n4�4%fjYCS �*����L�YaHK��R<Tn}�5H���F�X9�f`$	�#I��7��M�{������1R
aL��淢�5O�YFG�b��"��n�,p�R,�X�j*��ؼ���D����.�5��um��t�݃c(���t�W(f
��n �d�e��`������$�W5�LT�ѷg0J��+e�1���2��T#z�ó֑V�ѷ��G�[8��5jl8��o&쬘���%�Ô�M�X�ۉ� #n
o�7h̸��r���N��S�MJ�V�h�Q�N���޽���e��Vj���x�lVc���O+p�Γ��c�e�BB�1���(!���ԧ���X�<�Xz����*h[U�������Vf�i��!Vc�Aς�D���fg) ����zku��F�����Ii̷���za��͔��j�%�"l�%�r��e����T��n�m����Kb�k%��z�k�,p@9@aY���%�ҥ��#�vN���Ţ�WE�	}�#�����Q�Ҏ���#�Q��pV��|Y���Rh=70������T�~ٶ@�ݚg(�CHy�E%� /v�Y�N�Ԭ̗{��y&nHX��`����a�
5��7XзBpiB&�I��fVE
XmeEؽ��U��[�{KY0L�I-��
�HZv@�/ R����f�V��J��+1-Q���wrU���4���M�˯,e;b�<�oC�iB����Rho���q�Om����2|r����Rڔ1�KK�*p�����՚)ͥo�P�x�u	J��l-Uo&��D�ckElݚ��x�x��0�LIl�,��u�E�h��{��*YW�Ѕ�V�	��A)n��$]e�c #Z�Q���[��Q�%G�R�"&�Z�0 ���F��E	Kh�F�XEV)`a��,��"�6��bQ]�2;�b�ӌ
IV-���B��-�⬴Jm���Y4C�!u�-5Z{���	vj�q�Mܑ]]+�*�D �Cx�=tu�l<���;���҃�!��L�3M����b��=D6!�,קfbq��CNBt	xB�V0:��jƺ��2��$*#CT���D-�Z��Q�d`\��-���d�v���`���P��Zbԩ�(T��d����$Ǹࢠ"a����jVT��*��Zki,�o1dwS]�Gd��X�z�ʎ�$�V����oa�rŸ+/ 0;�����W6�XKh���"&�եPܬHC�h��2Dnl��m5��C$u��X Vɕ�+�cO���)�TF6��ԃ�vkv��J#h3�T�+f+y�G���K0�\���ZrFt�k,ފ-I���2Rܱ.F8�,%�`�$�X���6�u���bdBm��)}��,�t��F65jة饖~�Y��X��Yz$K��6mї1��w4�7���mY�r%h*�*cۨp⠠y�+����S����O
�v]lGcl���J8�ר��JJm�ˤԀPڂR��An���f��fR�������r��t�hx	ߤ��3�������5�n�큯F�t��-�R�x
��2��w2��C1|f�kj
�s.^S�A���T5�,=�e�kn����a��J4�����-It��n��t%�K6�����1[y)�۽[���hkA3X+u� �5�����BB�o�ɨ�b��\�l@�Q�W��n���6eX�6E<��l�X�i{�:�"5Z**W&�e��C&�Ӹ�]�y�a�SYN1�2@����wS�ܘ2ՠ�RK�Rb��֌pc���R��Kc�ƪ�0����6�ڱ2n�2r�-�fM�����Z�����o7J$+^�{\�,c��.K-�P^ݍ�5�:���da�4c�*�k&}cIum���ƛf��A+����͛��ڳJɦ*lml�	��]�R �V9�4��N�1nVb�z��hY{��yy�5�� MR�*V:{�ySmh���w��#�Ե�t�(]�B�3JQ:��I�����-E��V�Ĕ�5xطn+Md9�+l��+>&(�
5d
�v�X��S(So۱X`�lp]��J�8r"���y&3Ym�m��Tݨ�a�f(�
Z��E6�Vն����K)����7Qҷh���,���oq�t���wJ�j�6*�Q�#�ľ)]�u-�g�v����k�ҩ���*�D6�F��0KH��d������/RRT����-�Dk\�N]�j�pT(彬�����Ǫ�Q�;v��@�AN�ו4�V�6�0��ӕ��bA�7BK��a�.d���&�\�)���=`G��f�t�����,aKB��*d�0"�
�B�uT��	,܇D'okRo	��9�T҃c�U����'ҷn�-�e��
8�X3j��	Yu�Tl��gRRi�\#�:����z�gX�8���q�&�I����䨋@#j����E�l=�&� r�B��P7(�G�O��W�}u�`��:O ΊJ�A�m^�f�Sˬ��yR��q�ʼJ�#j�Ux�X�m�t��-U���efZ�
��S^dgLC�5J�,��/)�V������S�����#̛gf�*bgn̬u��Jz��q��s+4���*D��4� ��0�i�� ^'��;i4V�[f;̺Z	�KZ�f;9�ɥ��� ��J��5Ӳ���ܢ4V7#�s�-�v`C&j�T���t���D�����[���,���Y.��u-�*�ʳu�m��7�����"�RX��@P.�j��KRbY��� #ʄbum�"V]f:���H����t�k���˲�J}�SN�T����*��[�d��A�v��d����x��߮�M��HS:�^A����5˰f��JwMT��V![�H��87;9a��Z�����ZɎ�	ѝ܈�TP�Wr��-9��8�6X����a�V^�9IYN��ߐ�7 B�E��kcۥ�D*D�F�[�]n�Km*��`(0�i�q����$ѭS�{&e�b��_�[��]f2��b�sF4��*cĶ�\w5]͠0��GM
 a�AcH��ofD�n��[�Y��<��DF�^��U�uf���9��].����8/iU�E�:U�٬�m�t��`ձ�v�<��G�ՠ����H�YS^7p����Y
��n:Ԯ8K���"�O�W���)�ZH��d�YY�3�^��H���8N����
`�Y���/FX�jK��,:�h^e%N���(�J��2^�-��I��*�u�ڊP�5`�,��ᑜnP�5��������<��9Mi��fݹA��[x��:�YF*��н��;ʚ՘$5HjQv@��i)��F��Y�n��J�h�w5-Շ~nTr7R/�6����&y��|���W�R�)	w����@Q�FF̙K.�����\�&�X�jɶ����í�b�X�X�_dB�6���'d����&p�3rE�{A��˟O�b�-c�~WH��)�B�EH�j���1kYV��r�R��+��Y�J�ò�^�4���ֈ�D�F��`�1�VP�ٗb-lʄ��*U�2| ���J�eEI���i�4�n(>��[8(Q{F���&2<���6�.U��t�խX�L6�"3�-����[��T�a$��Q�1A��.^���7J*��������j(H�E�y.��v���:�y�Y�Ud�ZZ!�JJ�Ra�*��QK�Y�-��Gn�Xm�X��j��°&b���XkM̔n���B�ق����K˃��z��0���>o^֚�O(m(�-n=�z3v"�����*)�FX3)�ۻg>��e�
P����K�91!���K+Yb��	K�	{E7�;^"��`.�j����:Yם]��U�	��Y CN�K;��̗B��n�T��`7R�PB8�e�qK�'������J�������馩���k�����lI��E��Or]�ݷ[Ҳ�������]�m�	�R
;�������{�A)��S�(A���ن�R����1�51/~��ڳBE�B��p�b'X��3ȧ�l��lMZJ��Ik��Z���FыL/L.U�^�ƀAMwa���N�Z�,av� `Ւ�X�"� �Yy�⭁U�0`u�Xe��J�*�s�xe�*]�dP����d�xw�����h�^Eb�ZwY*#ǣ!WYmޞ4�]J���n�Xh����B+%���$ζ��i��C*�m��c�.�H�N�-Mke�[���u��&���%���j���X�iAm�Z���75ڣE�Z�%�D��_��� U,Z�
WV哔�TNL�_abE�Auw׎������=�-b��B��������rw�(?�f��L���Xf;W��&����ڣKSN�]�i�ˆ����TʹRU����~ZRI)��R��h��Cnٔ��I-7�޻�)�]�7c+-IykVV�U��q����Ft�wp��St�X�//+&����-���T  ZÙ�)6�]��V���*�VU�OHI-("�/+/��D7��Yٵ����&����U,	w�*I�M�-K�d���a-����D����ʵE�����U���E�5�7[)i��/k��� +"�z��M�.\�(R�߰��a��n�2����S��&�m����N�6( *�d<R�G#۬&�G�J�ۗ��,P���Y�Y��������s��Z�B]
�X�o�6�;4K�V�Vf˭��n\S2�b@�3�$�D��]ŷwI�#!��U6��9O�uF�D죢Lõj��u6u7'�Oؚ��^EhLF�l!�<����.��8H��݂ZƵ���оҮ��D�6�����a��D7���"��X���y�p���Y�<#,�ڰ�:�G�f�plF;�R�G��WJ�i�sb����N� �Q���݃#Z5Y��0�QXj���$�Rm��&�i֕�q��k/	ӥn���s-3K6��܉;�&V�r͠�Q��^G*�;�_L�S@8+q$�iۼ��*���޲2!@"w
R�Y���������3i(�&�o*���dcl���iV�J��^�V��y�^ec�osRv�Q9��� �sa^Vå��b�����A�e�Ck�ե�n\�Ks*m�˗Kc�N�Ӈ6AB���8/U��B|YB�\P*ǎ�19{JL�Qh��V�mR�.bH�2��=ؕ���zeYf{4EM��r�<۪u���6C���
�H��u1���+ �4fn0��*b��FiF�&�������i��,���� $e�V���X� �7�V��[�@�Öm,4���u�֪mc�1\��oh�kV@���2����*M�\/F~Po3n0�Yj�`��iC�^�ue�R�]�S0:���.��I�)��c�;�*��+��)��oYe�ܙ�ZQb@�R�md�4�e�3Z�v�hEwDB�j�:��Wm�,��Z�Idd����t5a���M�#��L� no ��������I�$�eQÙE�,K&�xwq�Ud�D\hXWa;�%��U�p���#(b���VJ���d��x�Tzƴ�1޽�� �ta���8(�Fޔ�c�")�ڒ\�j�1�&��,wd��X������f��P��ڗ��y%:Ѹ��5b�B̬aj�#9�XkH6^��E���)\k%��q�X�;�,ʖZ.}��Z�9�7�@H��ns_�At��@�����ڴ�a�����qU��JL+{'Z�q��+��%��cB��nLZ�5�[6��Jx��S24�cH:&�̳Y�������"6��hZ���a��FB5��e�^4@J����5z26Ѡ'$�4qZ����l��0!�0B݊b�Ӫ�87-�W#)�m�D�x�09��!�v"[��!=��`�.��t�Ws+	U݁�-�1��-���bJ�MюVH����r��������cU�:`:�d-����p^I*j��MRՉu^���bR)$j�х��|9�j:r�(ΘzU��W������8f,!�s�x���p��y�8/�9��[������/X.���i��]f���Y�TH/E�[�f���g�/n�uX��Sc/������Ir�ݸou�]��n��:����#�6��e�;��hr�{O���h9}\tu2�0�|@;�w`[ըM�V��C�5WS�c&�.����{-�[�vc�/��n�z���+�5���N}�M��G:�Ć��5�;P��-�n֪W�_c������]����,*Yg�C�rc���B�Y
^m�����]��=ۉ1�bWs�����H)�G�j��qЬ=�a���w_p{Yb�p�y�����/rL�-�ٴEΈ�%���z�_w�J���c�[���n�_V�r�]�Eu�,��.Gm�ԷV ��tk�\m��� z1�Ht<mmͅe2OP�,�8�9�_<�ڟd��:��z fit��̳�e1q�C*1S�l���5�'V�A��QVf]�s��B�9��"�̾�.ǃu]�Ҳt-&u�R�� ��8!�{�Ծ�!QC[]��C�<�K�D-N৪gF!�@�zP<F��ã�ŜrV�E�[�Z�xª�W����|S8p=��_So�0��dM6�V�L��Vk��T.�[�Cq��d�+/�x
�W8؛ۘ��.��iu��9��I*�.�v|��@���u:ܩ4��!��.����I���|i=�·��E�Y��P0d NթlZ8G�4���:6�^tĪw{Ά5S	��
J����c��S�)�0+uӰ�֛�ƞ<�
4� �6�ɧ��d��v��<�Wlm���#��]��l�T����e"�C8�YW9ku���LrLR��Y\�t+;l���h�/e�s.�-���ѕi|[��e�⟯\2��4�'�������{�NV[�dJgal��8g*Ҿ1�����R.-.���w�f�isgT�l��F�T�A[y��ub=��
���ŏQ��J5�h�:{ɳ�!봭����#��+v x���r��ۜ�h�|��-���xK2�ӟ6t�v-+�Y�,*���О3���op]�z1��v���VXr��н�Vr�ݩ׉�8"p���*%�V䢶;v�f;����#�B���Sy*����C��ه�bec�r���R�Ҵ�
V�J���n����7m�˔~�ؾ�Y2 �8Z>���ܳ݋�޻����s�X7�;�u0>S�츜Z�N�caUf��#����^VZ�^���Y�A���'pV���R���:�>�ݙ�uD&��}P��>B-Nm�!i4Ĝ�=3�-1mn_v�D���5�t�}ɣ���>�4殶tgd9�ZqY��V�Ķ1o w9v���~8%�r�],��\�Y�w.7�f�Vd�P����_f.�7t���h�w%W\�!J0J����ڛ$ǔ�ܺWsuU��f��87�ب��i�%\��	/YY���C�������-�����/�Y}16k��HL�u׫��ϧvְ�R�!��4���xu����.�{h��5j}��ջp�ܹ�x���J{�R�@��v_f�'A9{�⋚/)�BF�rF��i>�r�1U�h����!�u��:���+z�sRβ���J��Z��-��*TچɋEZ�m1%E��Z�gPԓ���p�̭�*�Zf�^nP\���K�C\î�^�,:�U��&`�q�|p՝{%wغMW�c���mJ�\��G2%oN�G�'7��u�c���޶���J��)\�h@�;����k��Qw�!Z���ɓ�0`��H���� .���̴�pC�ك��_��[C@S:��&��:��Z:������C�K`H�Xs)�����1D�-�\1������.�<6쉚WA.3Vo]�l����V�����)���]���剄Ov�T�Gz�E���*�F�v>��R��r�Ċ��}��n�V˺�^xpO��eZ']h|�!��h������7&�S`�n���gO���C��WkjW����ʾNrB��Hµ�%�jE��b�k�ڼ�}��_>���u9gx���(��t5��k2�����v�a��ץd9�t��/i_]']6'���WA�l�BM�ۋ��?ei�E��.��H��;����*T��"Z�AdԤ����oN��˛��e���A=Ɩ��pm ���Ѿ�.eծ��F�o�$�S间�6�R��n=�������di�/1�J����91��|a���^�>�U��Z�J�r�Lv��K�'R�75gL|��D��l��i��)xf���3��\���j;�E��a�Ʊ{�'k`��\ Vs����櫺�j��㕍Z����;��\ޞH��S,�/&EE2����~S����t|�p�r�:�6��
�L	V/�d�ۻ�a��t;j-wg�h�NS�w�r5�@�>�����s����1V�O����YCy��E)�'��6T�n�}It���B�>}�s�D���ۙu�ܧς��wN1���,C+yHu�[NJ��p���WTu�Z�v�U�;�+uwȹA��E�9�W�p����@��ھ[O��|�u�2�NMdrˌu�Jm��d/v(k0�w�xS�o����Bc�GLY�"g%��kC������o,���s�l�,������r�uN��3虘Yt�&h�6rZ3�j\/3k�ve%�2�I4v���+d�Մ&��5	�����4d�LB
�]�JNJw]Z��%�� ���(�v��8�-W�;��3L� ��J0P��Y��A�:Zqý�;;���R]�&�}ø7R�c�5�+<�h���i>j�s�kc��j)�f�if׃��:�=�KfŤx8@|`7�� �u9ۇ~�[��=+�i���ᾣ%p�ښ��d<<��N�a�Ә�v�3�j-9��fu��E
�}F��#�C�!�[g��Q������k�,�M�����B-\=�X�lW�]m�Lnus�c�kdl=���=7)΅AM��Ѝ����Z�m�SX�<�*��v;�r��˔R�=����-L�o8s����1��8k��X�v���ơ٣3�Ϳ�C��E�{��5!��uso�8'Hn�D���u������&��uۼ2�q���V&����f#Wҹ,te��K�8=̦rБ�af�hPb��˩ ��><nI+��$��fgEW��·�%��F��k���G�*FD�V밁�z�n�]�c���.��5Xz=47a�P�揵��U��w@���Y`�37�+�q��Z{u��lw�N�}�r�X:�b%pQd�,��@���}�8xdnW=�<���Lf�ݓ+�*�a�g���u;Y�όg���w���{�53��,]�=I�l՛Y�aN���6�R�O����]��bXh�;�e,"p��	*X�.��Q>��W<�+��V��0���ڝ�p��vi��%ӣ��t�VgM0Zͬ&��[�P���)���Z:r�l�vn��L�y���t�`���9��\�L/,�67Y��+��YS��M���V��tE3;B�J*1�A�n������4�-�sowPMRQ)�.�]$�l�ܷ��JӚ:�3'f����tp^b����K���}�XGA��7c��n��o�,�|����iչcG6j���}�.f���{��V��K���x�.��{Su�ndh&�4s��u�y!ޚ�9�x[��	ز����2��T���X���wkO7R1v�sml���̥P<��<�%
'��ŷ3vQ5k��WV�Y��<ǠMzܾ�Jﻷ�[�&�¹X��_a�f��~���`������ė\}����&B�
v+&�Ŋ�}�\���<gՔn��/���:żL�Ҽ,���J��ˌ)�
��ЇRWKQf��hު�y�E�5��huɜl^E����|��6�9�3�ª9	�2�1���<�8��>\gM��&��6��Vd�X�%�\t4e-���d���DJ⣝vD{���٤��WSj�fN�
�L��f,�h1�������G��2O�آ�]na˝�٫t���rF���WY��Z��ϖM�A2�VT�Ⱥ�[�W���vޑ
�
���}l\��P	@�+���zDB�֠���:k/i�yD�|ƗR��XZ˖�)�[B�:1jvR��ڋ�mec�����*��e��ԭ�ؾ�G��]$["R�8ٵ%�
:���s玬���^�-V����b�ӣ��s�ꧼ� ~�
�1�O�d�C&�:��u9u��]7RҲ��?8�CuN�;2�t�/��e7�1qN�\)�t�J���J�d��&��I9B�:d{�o"ܾ��7�9Q�|o�7���6�&Ю;I;���bO�q|��	!{��CM.Uh�wT+�!�{�+�t��/��(-;�/\�Ǽ�S�Aw�=��� �]9kq!W�XЍo[5�<:���Ï���� /+�7]�r�u-t���V\(%|k%��o[��_v�L.����w�Dz�'R�/9�'.�SF�ge��{^e�F��V�/��˫���e8�V�(e�N!�
Ok:��f$�+nb����ETOM0E�l�������(Ҝ{�B�M�Y���O�}�J\��9���Zj9�W��2�5�����E���kfBܻ	P���!q��P� eb��Q��=a^�z/����e8-(�k`!����wΫ�\⢫�7RQfP}؁��0��eWE5�HC����e]��]X��R��F_X��	.��q;L�����7C��g�wk�ډ��Z�=��.p�Zth�Ö�;�{2 �'Ng�����q��Fm���K]-�� #mN"fQyC�k�$�p��0Q�,��D�sM�SCze9��6զeά��8�WmN���A56͝�K��
���=LYC7���8���&���c��t�D�3(�[�wɥ�"�Щ|��� �N�5�3pI,�P`�=���x���=~�vB-��W�V�K�QFB]nTZf��r=�k�ᣜrí����1v�YsVN���]�˽��\Շ�¤ /���mj�Ń���<Э������Z���ܩ�qk�mťj��pmǝI�޺�0 !�0�3��W��1�(��K����I�im>�:�CY��n�6�U�o��-�)^wguآ%���tGU��yD[ؠ���[�s��Vt=wN�&8Y����7\�\ˁw��V�N��c�:���X�Y1�S/�������wt'r%���֚w�D��m�8�⸷tw_un��w9�ơ�����֣�� �ɞJ�uE�8�[��� ��U�C�7 ��M,�t�E�P�Æ��NF�Ǚ�]r���kO)�gr̳�Ҿ�[t1pb�ecC.p�ys^:�f�$��e����O�� ����ݱ0��gh��!��̮	��t�dH;w}VE�L������]wfe$r��H$SMn꒙A<�˺����+vf��㡔�[��^^iE���x8�/v_�AU��[�m[]���X�&ܫ�M�X�`jX*�vþ���Vu�g�?�S�� �c����0�Gy�����q�t���P{��'Qh=|3uN�Q�u5��zW3�!�,�k����xZwr�ǜ&��r�hqC�ݜZ�C�*|�j��m�'��۝�1�è;3S@��pz�yw.S�n�l+u�!������#�-��]V�,�MX�ᶅ���b;�}iX@9w�Wp���pQ娶ە��k�M�nT2��7aH�������G7R�2��K���$U��1!�Wup���d��XKA��ہIX����aO8Ŏ�����n�N�xm�$u/qY��yJ�A�����QSVR������⁄�04�ޱ*IS���;�!���U����l9�t���2U�s�l�$����.e�)�s�F��Nӛ���ԭaJ�_er���3���-�E����4��TZ�3��LH|.�L��Uoc��AP�2�=���]���.=}ܩ`��qf�0�F��)��Ml�w\��8���	�w�*+ƆS��sNRC)�Ѡ�������eۖ��#VK��X@Ė�k������K������Q��8�k["�����hX�\�d�Კ����w�NS�Y 4r�
�ҷj�����D�@Mڜ �w$#�՞y:;��VIt�ׯz�v���坛b��uAx�g5��ۺ���"�OTU�(*n�n��a{��,�4��ڽ���G-&�u�k(v�;���8s��{Kc�[vp�p�k���s)&��0�噓G_:xQֻ��#�(jP��f���XY:�����*�_L��I���-��羳�x�[��Y�f���Wf�%�ya�������Ǥ7K�+�'f�\��Z@�Y������,���X��W;��Z8��ޣ:�4	/w��K4#�u�LWkhr�*^k碒,�nmC�0k��us�ȉ���]�>�H����	L��u6�;6r�'��c��\4�'|f��W�+�+��(Y�Y����0ul����mt}�ցs�[i��k^%��G���&�tw��4��"��:�uyy�{�-�y����R�s�
,XBA0�g4�́��&r2�^��v)*7�m;�ҝG��+���r��'�o9�a�b��]w�`z�oM����{�.�w�p<v��������Ņ;�+�=$�9�u�n��T�F;T��W�L|y�j�7�����W9e�`1��e��vV�:%�Ȏ�K�Qv"�y�.T\o%���F�;�7O�I��\���e'V_m�Gd��.�u<��@	.j�Dۢg�Q��iږ��z�QŇ�lZ��Q�{��&�keQ���������}����I���!$ I;�u�����I���R3��F�0���n�*#�8`*��p�f�.!!�SI@-F#t5˺̼{a��9t�S|k��}�on��.h��f�lDN��p�SG��r�8p�o�}�	��̺�X�B���G4���h*�C�Dɛ�g&4`&)��9�v,|S
���sh�[ʳX6�P7��z�o��+s��k���KW�rȱ+�͵]�vP�u������N��l�͖GM���4����af�M_R���1��
�����ً���43冯;���w�o,�X�W��WBnѾ빆ފi�Z��m
�,�Gm�a�j�0���vRͰ��kjd�i�ɑ�#�4[�\V�o���5�Rar����������o�o%i�l)����i*GQ� �i�]��'6�+U񑝳+7͙I7ki�9��8M��ȹ�uLU�E�sV�)U�[�yC��P*�໩.N�8��λ 8����=���JK��vD���J�=��k��AfVl�]9%NM��D{�Y	F��`�V�ǣ�`�����7m6�u��u�Ô�f}�|Y=%<[ԛTI���}��띎Ź/z�4��8�r*����x�pA��yrOS��[J�yI&�>��lp{o^C��,4Wk�X���R�ۿ�Rg2�Ӧ�΢�H�`����ʸ�,��J�+z�p�)֍m�9���׷u���Q��'3�u�lp�b�8�9�7)d��xV��WAVճ�m�ˡ]�7�6�7&�V��i�jx�:[��;y|�kkVЮ�̥iLO�1O�h�w�#���VNcz�b�V��N����k��ޫ¬���Eڂ�q�n6Pd�H��.�A8���9�噔�k���*z�
z�9�X�a��5΢��Y3^I(�o��^BMG�����݊�#�廱�)��o�TE����fϐ�}4�| �b@tK�����Ձ�E��uc7,�]��Tܵ�����	�mS�q�6�����rT�%���W�WE�v��B_A��T57:�=|W[�Os�E��޻�h��$h侧�VM(�Z���\�P� S��]#n\�+��=g���V:�w�FF���KM����\��JNm#ìU����%�ڻ��JN��������5Ú�cR�� ��W1'	��a�s��nwe�W�p4�f(n��]�1�c�Ս��Qʎ�u"l�-��]����?m2�-��:���e�Ď�޺���5�@WR[��mԽ���v�J̽��H^o�hi�9g�VF��rк�\iR7N�U�2^�\+���x�A86K;$@����o��;.NQwCZ�9{��]�1C�٦j�a���8��47�m�Q 8�V��8�gY9fO��g$o�KL�p������f���\r��Q"�խ�4Za�8���Yb�ӓE��[1f�ivd2!q���:�n�Y����� ��m�\{X�WLWE��O/;�S��w�	2`�V*���2���]�w�p'���oEp��ϱY1R{Svj\�t�\�Fp�i��h%���I�ɕ�f�ֵ�er��nQ�5�����m��8˼w��&�p�3��l(��x�W(j�e��{j����S7���!熵R�D�,�r3n	��ibD �jj�[Wcc��뾽$>�5�s.�*Ƹ	�~�n��G�r�5��<�a�A�bW��(����D�g5��H�ӗt �X�E��bH�P��xG]\b�X#ὕұ�4��̩�5�o9!�e��؝��%��p��/9t�"�֍��W�Sw�,/7i��;��m:�O38Fn��7��C��˘gg5���l-�]��8���Z��.붦��	�� �����=�Ԕ��ɍ��9� ����j�T�U;��[n/�*������� �<C��w�gx�eb�i�Kv^����I��T�զ䮒�EX��e3[=�Z��G/�I�Ge��C�̂��s�4����Nц��}�CD?����t�c �� ��JT����S/oa��i�]J���O��}���`%g���!6�1Έ��G6�>�vXC^I�΋ �y}�%�p�����۲4i�B���`凜�t��\ 9:M��f�V�M�ӷ��=�x�x"�r��Rf��AT%g]fD^��B(�|k-WZ Ҭ�m��]7���5]��kn���I��ᇺrTI6�Q�P�8�5��'ԫFF�y��mj]�d�B�습8վeghЄ}f]��.m��=B��k��m6��Zk����Ѳn���@N3*���0�iR�9֣W@��@ރu��*�ѳ*�]�#o@�7L�;4�ue��*mdAI��cM+���w]A�5�ż��)]�WI�k7T�ƭu��Z��0$N��z�W^�Ca�9�Ŧڂ���0gr�M��`s�(9�\���[)�Rk5s��нȵd��mp�gK��p�ȉ��勌Z;���j#�w�^��=��r�3���l�.!1s�)��X�W��wٓx3��tqMƵ�&ռ9 ���h���#ֆ�o�d�Iձ�C�փ�6�����ّި;�u�+j�Z����:�Z$f˫�����i)�P�I��rᭅu�r���ּݔ�����[����*�v����噒�2Ĥn�*P���v�{L��%f���'4:*�-v�����');����8��6ƺcuLx,�M4�M׫ ��+h�]b!ͧw�o)�v��Z�ѭ�TWۈѼ;�}����I^��6Yj��IQCW��:�wj֤mq죷YQ+�~vcUd�i��^��:�'ָQ���N�E�YըvD��V��vD��w�n���mf[��*bo�V�{y:���Ę�ɦɂ��*��{5o���
��i����ڎ9��6,T�;���|�S��h����j=���$����§u-��̀\�.쇩���{__r��V-�c�J���V��v����or�	�"���ƤʴtP���yQVfRoV�ҵۊľ�z�-�zط��u+��p
U�6�.�H��B;�|��ǫ,��D$��SB��ٽ'J���IT׊�;�j
w*	�
��f; V
�L Ps�K��U��m��;��uڏA�m�0�;�����K)�
�е������bYJ�2.q��w���YdW$oj`��FQS�9-7#�{wLR��قRօ�2�k��-��Y����J���.�[��TC;�W*��3�:CXjR�tk[8�y-�r��o6��+�"mV9�iE�F��{٫����κ��(�=��b���3���F
l�{�+<�L�Z�0���)'�b�f�2Aջ!Wʤ
��3N�;fǡ4��g	o���"f��̵�kE>ӯy$� `��*C�>z���D.��>ǒ�`�KQ�U�J�:JVj���m]��P�u*賭e�7�V-U�s8iR�mrXvv�A�������ҹ�ifU�wh��F�ٸ�5=�S�Y�T��]\y@�V7YW1��t%_T�ynG����)u.˱��U��t���ܳVk�=CU<��嗷 ���
)�z�b������
��/!4�h����H��xq'�X٘j�J�=��J��-`(�8�n��.��P<�6vf6j�7�	�dj�8��yt�x:-8�N9g �M����mM�޵����ʂ�"GKx#�a:2�<�x�eݧа�GTȥm���3qvk@��T��Xq��QlM�{�1�m$Lyf�ξȓ'39t�7^5ƅ�^�	CR�k,�͙Ǿ�����o��.i�*��b}�.��7[]��[��r]��k�>�Jn�N" H,T���p�*g9�!x��jb�7��[bT�au��[o�2�W��ِ�WJ�� _f�ͷ�gSp�[u�kY���=���n�I+.���o��	��vubp��]m�9���A;3�n=�Oz�B�3�R�J�S�β�kÝ`�V���Ǝ
�(m��_X�S�"�i���uWL�r[y���W��-Vl>Z�����ڽT%aԇ���±iY��܌QK�2`��gd����DqG�E�P�A])Ӝ���և)].��Z�.���v�%NC��@�/��:^��ce[��������4)��B��U�n=�V�[u�5�އY��$2�:��{[�a=rrxR,^d膙+�޼4�!ap��2(�=�}C3Vq�D�a��a;�1_E\f��dY&��ٳ��	�ڔe)��$e�v^w$�:Ѯ��A	7b��i�2��!��� �/^�<(?������QNK�S[m)�kN�
x�ɽ��yj����<f��6��D"����J�W%57qJh\x7���Zq>@R��8��ۥ�<�T�dN��0���M����]=c�w��	el�$wE�S�l���{9Lt�YGupS(`�<����J����RkT��f�;]�������f�\��G�
[���R���li)�*:YE:���s��Ց�@��b5r.��iB�#�S�2�ޚ B�]ݗb�.�`�[�֥b��d�����`�4
�j
��<��n'��9f���^��gf��1:y��2���i��-cP�1���VDR��^!�\��D�ɇV��������wsvWY�]��7��ֳ�(۬�h1F�ᚆ�Fr�]l���j���jI�+`��RF��Ҳ��&�z����pzh��\���3_Mc�Uv�n��mC��F�j����C���K���2þ�u":�����}%���x��k7b�H��5U��9��Z���Ǒ.�OSc��Tz����YƋ1��_G��f������ކ{3F�c�+@�f�[N�)�!P,쬮2U#Lk������x��tKi9��PU�@�c���ɚB��S���4�:*���e��pS1o4���
MZк�ۦ��;Sl��q��Z��<*�N�I-t�u�:�	(��[P�;t��Y�.}b�����4���6g,�t����X��FS����}��0�y�컳G�׳3ʭJ�W�Q;9%!��0��u$�m�YVIL�w+��Θy{,urn�їJ�B:���!U�0�b�Ӑ���,�:u��'���\�x��n�/l�"�4ąmMڶ�-Ւ�*y{���I��ϟv�ڣ0O�Ap�;r�ԭ���͚�����ޒR|��{q�%d�����v	�9�J3��V����\��!����9����������0G/IY�g0n>՜��-����f������ƦM]M�S�(Qd`�ē�cd���Z����C�V��V�(ܹ��˕��t��iG�o�bξ�ҧcu$��<���8 q��V�RCm��cw�-WKpN�w8%w�[�G)�i7hG�(㱀l]L��2��杔�J��]��t��A���uph��d�1m�$�N��u;��R2�t�f��8�Iv00�Y�W},�wp_r�0�|��K1���:E��@�Js������µw"��[�+�'ҝɕ�Ѧ�"S�5 "�Y���5�̠O#��4�(Z�PgnE�u�j�#�=�l���QCJ��4+6Sյ�oi�;��g[��Ѧ񗖺�؎%ug�{gJK�n&vK��-*Y �6��Y�n�j�S5�;�-#UZ�9m�*+�|2���^��`��T�1�]��T0�|��u%��`�h{{Hwf��̘�z�F��]`l-�J�z4��u�lͶ\��u��V�v$�Q�j՛���u��Vz�	pwM����("�E�R�*��8D@v*�[��)j�my�6F�WX)�ݠr�:![N�蓂x��3h6
�65�C|3�"��³nf_]:Ɋ�I�T�p���F���Z�����Hh�����М��r���m=൝�W��]���M�e�$�_T|TETu��`�g�ڥ0�MQ�r��#����ټ.��ͷ��������o���LS��h�cfîT�e���S��]r�M�W{�e�qCV��\룽��	�:�
5�����y�|����m���a��x��њ�H+l�i��V��y͚�]O�]�L��y%"�Q:�έ��8R7�Kx!*�)�P%�-S�,���Òp��U���zw���E�\ ����ɦ�7�õp�1ic�m�ݫbX��d:���˵�8�V���-Z�.��%�]][��ζ-k�q�*�«��t�(�R���U=X���O��W�����M��i�9a�a�y��Po$��v`�B�Ӻs:��Z�L|A��x�ܹ��{PDo��X#)�ju%SN<W�=�Na#aN��QE��KO�8�3�d�/nֆ�u1� ��4�5�gu��b�H;[�sG�i�|m�]k�5����[�z���٫�]�Gsd{��������\�M���^_X.��tz&�v��5F�WV�vX��x�����
Y&�f,u}t6�"B!1Zޑ8��� �,�7Vҕ��p.�!�v����.�Z'V��������v�]r��I�`�x����"m+��1f�f;W������ZK��@��OZ�M-ߛr�N�{��]Y4�`N�F����6�7��];�o��VL�]���ՈF����Ŧ��c�N��!<� �r<i
�y���5�\sneFWL�9�P���7dʺX���1��GmD/\?-�
�u���Į��Q!D^���v�܊���Cm��歩�Q�ʐ������~�7�P�����M�N�+�޸*����f�]w{λ���}3�X�X֗���aڔ,'t.�h���Gfhh����9&٬�i���*�W`�;��&����OZ��*���p��%�w{.������������[�ћ;8���y�t�w:�\��V�Hk���/{q@(QamJ�V���]�2�@ �V� �y�nTS�Ԯƺ�����+	a���b����1P���]�}{ݮ����3r�gr"Ҳ�H���HB[è
]�
��.k��SO�.�Z9+�^�8��e=h^J�d7�3h))Ѷo;!��o�[sv�r��Z�����əo�`<�vv!f�9��R˝�t��Q#��{"Jj�D�[u����պ��xd#7��i���A0��2-8*oڶ�Ѥ�����=�Fu���9{|�˫Qq�����QZ3*�S��	c��S�m�F�^�4�x�r����9p��.��{ew|��S�fAk�v�B���e\+��Z8��v =�wܲ�P7!�O�F^��|�j�6q*������U���̇��7�$g_.�Xn1�,9ܨ�*�rۂջ�B�g�+ܝlR�`Gܚ\�F������;Y&)V<���x׋� ��6���4���0
�(9����ʾ,%v�B���+Ow!�[�Mwf丑�m�n��WG%;s�s�iN}�3���t��}ozӻn�"([n�t��EiΆ)���/]�;��|���$ir�9v5�E��nwe�mD�7ua�E��B��æ3�Ih�.��l����v��v20b��{�[3�̐1{�{)r��8���?
P��Eb*�b�T�QTƥF�QQ�$b�q*F5�0D��W-�X��DUTLe����T�
�m-�б�Ƣ�cUjXc
�(��d���2���j(��*(��[b5�%�p��X!�PP���(���T��X��+��J���,*e��b���ʕ"	(�b��"�(8�J�9eW���QIPl���J���Y.R�X�&%nY������8�X֕��n5�Q"�)�*,(�"�70�S"(�Z�+*��1U�DF�(�*\)U"�Y*"VVTYr�*,X�,�F ԰�*��,2ʣ�&5m�ĩ�E��(��,�m��-U��U�%ʤ�AV*�TX+iDX�"�A�m�h�m��%B�V��j��Q�R�Q�eE��� ��~�nz�)�y6����I�wS�;�:vV91���o���o����
j��	��w��^���uhi�e��NΕUˇG�%A�M�n�g'.�����ҭ{���D���U3��5]ޞP[ƫ6=�k�@����w��[]���/�Wl�BR�xL�E�w�$_��zI~�'�q���۱��w.��uf����޴dVa}[D䆟#��%Q�Sb��O'^e7;�'FF+�WJU�q<�Ȼ�23t����j�}��=J�z�,�Z@���W��p���]
����0�{��L:�I�^�gR{)�>}����R�^�U��۲�k�3�]L��d��*�0��(/Ҋ�6���x{"�G��*^�M_N��=�\�̺-�Q�} ����/���מ�T��G�jk��J��R97����˵�W��{�-�x�/�D}�zf%����(g�\��~:^��,-*��."�o�rS۱�G6�2�K����
��r��/� ��ļ3���=C�q�o��gUЅ19������ky�
�#�U���u|%@q�Sl3��	�����w��;�Ң�Br� d��.X\|�Ԧ@ss��_'�����N�)�e��uKvHe�L�B����W�W:���Ok�����s���&Ӕ�ԩW�wv�|6��|�v,�͜tqHi����LV>ÔW-�/C��[G}���m�=�t�=gU�8b�\^Um��B�(.\�J��QE�d����dݲ��˸qx�����8R��!:
���g�V�u&���"�U\f��[e`,�SQ��qv
�P痾=��D�ӦL^�cY�PdJ(y�v�X]H��āfo��0ׇ���{{���^�v�mhE2�miqq��xs����/D�"D�H��@mu2ǆ�
U�nX��Ku�,�^��	�֔�a�R�dQ�<}�fq�O[ŀ�!�t?qX��^�g��{R�R~[�)����҇�.C��b8���|�L;N�+M\�N�ǆ�ٍ�N�k��|7Y>"�"��V)t]yv���nE襤�`�`Fܬ�?}�Ծ�">�x�ׇl�'K�v��a����˳�H��[�xg��<\����g�O�}(�E۔Ы�Y��{���G�r�
t̀�n�\0:�M�2����΢Fj�����R��y�\a��ͽ�Ǐ;|f�l���TDIC:
���q�_�f3�J��0m��!��}����DTrۮ>&ױ�:1p���}�n��s�������������ޮ�����7NW}@XӛB���G}���3$�[S���h�awa��iX��.����.��k����S�m���\V�Ƴ���:J�M�&�k��m]���3�h���|��ڶ�CL���%Xw	"��-�\}�sl<G�i�B�yJA��77�O2��JC�i_
��R/�^<;/L��Vt���bn��2�2f�xo؅�4ax���7���PN5g�Uz,ʖ5eG��`��A��޿�hW]�6�WB�f�Ep~�gh��ŉ���	��c>�xa,e�b��7�u��*�=]��z��w�=�3��ҖTj�_�8��chM�7�Ҵ��MmUq�/�c�I~{�5��Ι5�Kv��)�-F�!3�뼷�X��mu@ꠗ��euYjľ��er��@;�].D�Nct���ܑ���M�e�=;��C����]��C�*#I<�]�ȩ���P��3�UU���f5r�3�-��E9S˾Q�A��Ɛ���8������T��ʩ{n`��#[�q^���%�y�P�
�`$�]�:X�=i�v�j�Sl{��"ۏ��2Tś B�b�Wek���=���ϞY0�a�hs�I�Gօ���c���s�Z��Ols޷���W8�u�b��gI|7J_ط�ꎅ��E��7J�/Jځ�aiꁲ���:뚫�Ov�rY�ҩ����y;1�j�y���h
W������o��LaE���|)���)�U}t�ΰ s������b��8yZ���k���g���.�w�Cs#�&��S#�|��Cz[�]��,_=>�ɗ؎�����_��/T�KɁ�5v4�mh���'�Cs)%C�"��T�"��?a��1y[���Ͻ��z 喰��\P�2탁�$xjyXyv}޴�7�O+��	����U��Y{c��<e�g�P�=����h�r�Zf4M�2M��XyV&��4�s�����e�N
p����	��[Z|(����nV����wF�ǈ�^/R��'�����6`�dA/�3�o��K��o���ƽ^y��GQ�nÆc|�h��f૑���g{�Xʄ���J��c+*�e&��	�+�V���lc���+��	w��٦��<7���wc1AZ������;��h͡��&+��t��+�.X�������S�{O��*RM�Z���`��d�t�ϩ��<\��� �ye�X��E���K֧��ET�a�F����I�ʒ��_\�#�b�K��/�����{L�
�������Y˭����jeH6ܸ�z�hx5S䷇)szV�=웾\��Cƞ���/�=�5V[�%�N ���L�j�l;�`{w�$e�R�6�D�s)�7�t���4�U\�I_)ڂ�z��s�T�A[j�8^�����b�q6'[ۘU��@����Ȥ����F:���~�(�&Z^aC=�d����j)����)�����'=����eA����]��t��\D$�k׳0V}\񥚰�7�0�O7�Y�(j�;Sv�^���{5ԣ^��S��\�G��4Mt� ��8�]h7R�)YZ��ﴧ/ْ�B<�Iꎽ�,of��ׅF��Y���4h*�GĴ��e���A�?W*4j	\o�������x� �|v///N4��^*bp\���A��@��H���B��]���MkY�Z�������'Z���X�.���	BZ�reB/還���Bg����A߉�z���+{�-}Gk5[I�1�֌��/�Um�CO��B����BB�{�<r_g���+,���hu��b�>�r!�ys�FwK	c�ʌ+,�V�׹z?kG�Z�����攕�Vh�c���2���Zah�e/�����Q�=� \F ����,]�f�'4�B�}����3�W�����'�
�zU%�|W��qpu/$���7�/]Ѓ<��E��-��j7:+�oB���v)��.�9t��r�n�b���:+���b�k*gOP�����U��ꊻk�5!�Ct����uf�m�v#x�-�#NQ��j8�-|>3R�Ġ�,�w�y@eڝD���{��{��j�ݚ����pP.��� ~��� �
�/}e�v�����ǐ
��6;��L���!�~���g���?#�/L���h��\���-=n��T �&��}Tku��w��"��j����E��yqq,ܶfS��c����S��vRS�8�����C۲��v�C݁=1f��ZZ��|%@w�T1f�f'S�<���W���J��u�&�`N�3�>��3e���PĽJu*Eֱa_˚�=J(��	�^��/�Tm)����W�8�y���<{��\mm&�<d[U\}�(�]���;�25��ufzn{�;�<��#�h<�Ǟ�`�_���Ύ����<�9-�*��\�K��=U�����=�u��yx&oe�륙BQx�{�(x_Ռ���]��tk��?P~���9�f=��	'{XR-�}=���7hW�ψ��{�{���֫����_-|C�nB��o�y*������<����]�I:CŹ�n�v�+i�f'�1�y�i{k�vc>��8$i1�oE�`���셬**�o2Ћ<U�=C�oVt�X|������']*���:�Q�.��v��7P�y�Lr�gى9ֵKxCr��w(vb:��w2��i���oz�k��7��W����1�g���e��G�s�W��R�ǳg��Vlp֋�6�T������	쥮��o�e^�V"G_������s}/��3�W��p?��Ӱ;;�3S�xd��n����Ӫ�z^�=�y$�}Оp�/�1�Ξ�]K�r�8S�:�>��<K���o_�s�ҡ������i������{ǝ��Y�O�ߏ���>͍ܾ�8zj�5\�w#Y|'؜S��vN��Ѱ�:}T�����?.ʭ��X[tw�/�ujv�J�~����a�D�@ܷico���^9;gc��G��� y�</b�8Y'��q�����fs�׷>�����?r���+�Ӱ�N�Ke�Z趲߲d���L�0�=]��o��?R��%Λ<+�=c z��ܾ*�:�����_Tf��]�%�u�[b,�7G5��h'��!�!�|c�� �K�̹��'uvNU� �����z����^��KX{\+��.��;�=<�Z�����8��mvqu���T�^�� B�zs��#�{��$	���fJ��\H�o�q���78�=�z6��7�$�	�P�5�I�3탺ĳ����T�q'.x̵���$��4\�^9����7����S�R��d�yG�N��*g`�B�,Q����[c�e�j�r߻��f�κ8�ojmd�V��u:à셼a�����nmr��ۑˏ��3_wm�౽[�k:\�9kg��s�ׂ他d���X;6��_f9[���n7�b�hR��d�'������UǑS���Z,96�	M�k8l�+���;u�mwP�/̷Vsz���v_G#�e0�x5�v0��v�i�/���)����'ٺnw��3t&��5bą���5\���^T��������Ý��7���=1�nm�}8��~��گ+��dG�>V�]~����/��C��rҶ?���}[�ŝ��S�&L�R��U��; l"�����ָ��~Qlޘ����M�xWS�Nn�s��o���� �7��8����|l����2����Йi�Z�ӥ|�4��Y����um��@e� ��nmڢ2�P�wnZ-Vn�Jlިolu��S����VȾ��7ٌvf[<۩m#έN���f�]EC4OL��H�v1���?}�u/���Oת�������Ǭ}���a�YՕ�	�J�f{�&Dh��N��ۖ�0��`qǵ�fы}v�F%I����Y��x'ު��8o��s��0���ݽȯ�Q�D��5fL�=h�N�t�Z���-v+`4/�6<Ğ�A(	�\�3�]������	&��w!��z�m�<���V[�'�����sf����"�פ�G$���nyUk�\��H�>n�[Ŋ:塽y�]��w*1���w�ԖY-	bO9%]�cn�j=�/}='����*�47�:>�:�F��T�z�3�?/a��I��ˏ�������ԋ/�D��v}�t>}r�'-����Bk<F����>�V�yᲀ����WE]�$��%�_�`���~�f�;��j�M����6��x���k'|p�9����;����.L�}ϴZ������1�86���ؼ�`���2���)�i��,�+��ܽy��+�tX��KW;8)�횓:I���;J���_��(��Z��+a��p�t�'�ŭ<��x��&K��n�<�Z������\}�T��^�d0�-c�u��#�^-�Wnsۿ*�k�|ag�r�t&��Z)i��R��'7:���ԯw��=�\�=�s���K���9=:�7TS���Rr�$w'fj�up�����W�;i�����_���92%^�������Y�L�c϶^��Ԅo��ͻ|۩��^�m:��R��S[����r���}R�w�c�:�E��R���M���y>�[�Ι����a�SP�Hu+ؽ��/n��],'/�:=��z�C�ٶE�=z������*��W��36�pah�/p���XNt�%�YT�ZCܗ{bj	G�<�^
����ϓ'g
��C�%d������Eݨ���{��^d�]�Xp�²uVs�#>�O�d���5�
�}���w��A��h�����[���$"]����]�p==�2��X��x���載@��"p���`oe�������-cZ���^McA>;+Unu��g"�t�sT�oo��
����WLڢD}��[��Q���0:����\��]e����qWd���E6tn�V�]��5q��W��W==+��>���љ�����U��=���&,� �w�]}��>u���ŭ�5����V��G>h���:~�X���שL(��:�LH�u|�S9���S����q��.��"���H�J��{ZM������`�3,1�1��FE��{w�VT�Hss\��f���*Do N�c��plƇ�<U)PR�mH2z������5C��U�{:�"�y�`��&��{"�P֌��=��2\�͕c~��:M��J�	�Է���
I�ukH�l���C��J��	��vs1�y2�T�ƍt��ꖄ8bՉ*�����.2�;4�!K��\3�CXJ�,.u3iKX1�>=�h��zқ��+��'�9�w\�Ӭ��wZ���F�)X)�(b��I7e�� -fNN�cf<``�*`�[�1j_E7+��@���]惯�� C��n�bvc��m��@�3V_g"����54Չ�u�^:�m8z��+��S�642��^�ݕ�HX��]`�%ҽ���2�kJ�`��\���41 �He�y���` �r��MNn�=�"�>��8�ԇ��5���՝O�_]��ݐ�� I�,��xO\�<KU'&���<���y�8'F%+8�>�R)!�;k~���G��W��.�6���/)���
Eڬ4b\�j.�r�|��;mX��>R��� �en<����RP�R��Դ�#�VX��}]Zu��uu�gd��(OMQ!�LѢwUʝ|{�����AA\|����jٷz���>T���5`�,s	#bʉ	3�i�f�7��϶��UC������i�i"�z�j�*�0��'��o��%��/�)b.X�R�8���JRtG76n���I.���OD%��������-�|��@f%��w���	�g�Ļ�6�1�s_C���P\r��T��ӭ��g:��KC3P����N�b�Q�v�v���SK%u+�e��=�ne@��n�1��*RҮ�2'i7W�VN���i��S87(�\�'+���[��]r���gs/���1�������	����N��X��q�K�[%;�5���~��]���>5��S6����[������t����%	�}ʌ4z�klU悎��ݧoX��䊴Ɓ8v�8��a�}*�.�U�i*�82���Q�'�ܧh�{8N����k�s��ˌҡ�\�K;Yˤ����;���g;y)	vw��W;�byS��|�-��	U�eDPm�ղ�X���"��D�Z6�1��V9q�-j(����X�d���s2*�s1�˖Զ�3
���1qT-��F
E�����*����F�6�X�e)h��)Qҭ�J%�Ҩ[E�k�q�QŹl̦+��X�Y�K�+jی̲(�5��f8ڙmqŰm�B��[V�JR�AA�e0D�V!ZQ�q���\�V"7.
1DD�ˋcJ�6ʋb�\�.Zf)L�ģj�,��������+A-���*E�0��̪�c�6elZ���iDp�&[Q\LA��*W)�*�)hX��I��ƥIF(��GX)�EC)XT�eD�-��+jԊ.2��mi�T29���Q̷
ʅI�̕U2��
ʕKek*[PDR��fQm�X�Y���amQ ]U�]p��P�\A�V��h�	m�j���]���E����W��M��3�Z��E����We^�Aג{Lk�<j�u{Ͱ�j̓6o��&v��6�,�Gh/�p{�ִ�?}����%��1f��w�62M�y(�%�I�]Hhyè�����v;��9�Q���oۜe�9��o����H�R-���5�Sܪ�'��ǽkۓ�� �B�4��A��/F3��|��%_�R�?Vƞ92R�ߩm�*?_�a���CY�IΫ��7�c�3�o����WQ�.��A��&�Ob���l֋{ދ����c����Y�^>��ϱݱ�7�\�״�Ϝd�r+�KbÁ��r�@o�܆	�<��cF�`K؇XkrzJ�s홹<���П8�q�-��=����6x�[��i;�"�s�;$Yj��y�ۛlf���X�cӟw�\�I�����_={Bn��}������a�n,���l��[�ړ�:��ɱ��{�o�݄���^8;Q=���U>����X��m�����p��ۼ	nY\�&��ؘ�S&��q�����mbV��F�b �s"�ó��5�5�����`�[�M�m���[}S"�!d~j��h2����ẫZ@5�M(�������q��0><�\sx13n� }�XS����rAዣ��y�a�ޘ��O��7zq��t�����s1p�����wV�1��u�-��%%���i˘N�8��+:XWR�ܫ�w���+hQ�ozz�"N��	��W�Θ\~�l�v٣���W�{����^d�yu�w��{M}�#�������(���;֔�w�Q�Y3rs){N�}ϼ�l�vs��G�TO5A=��W�Qt�ܗ�7�^�5{�g�z�y��fo��5W�Y�����N��@�7:x��\:e�����aӲ�����f_3����h�n���"~��>ǲU����Ϝ�ׂ��tM�<h�m���4�w�{7�[5~��R��G�*{�
�aɶ&��{���b����WG���]�[cA=�m�뻏R���{�!^\��3�P�5k��$�
�����^��-N{���sн	�V���?V�.K���mf����F�wnl�:m��Ӿvz�t�]|�[�8+�b����������Tb$7��W)gsa01'ݣ���'�{7���n�j9��,H_�����?�l��ŏ�E~W�#����.׾�'��;�����t���_8}bą���b��P�l0�]S�;�<Ͷ�z{���&����{�;��6�΂��������N,ftUmT�e{y�N 6	�>2�=<��-{�&��>������rS�Ls���NR���LK��x�0�H�m#ά)ӭ1I�����r�vT�^o�kz�:�bm�\��H����W�e��8ӿ���JF:[g;9�=����e�X+��^�3>�p�S~=;��}��[��򞾳7�%ģc��~��u��:����</���1!��X	Θ\j'�P���O�;ɕ������pS���ۈ���
��Ծ|$n	�zgC!~��׫�u��������z~��twΎ����@��a.v+e�͜v�������҈�
���CҞhΝ�j_�y�jL�&8��T ��,�����s"��~��������n��a�Җ��Sf��-��½��թAj�}�9hBS%��]��u��H�������<����������1���7�k�z���kt^�� sy�<}�$�	gZ"��u�C�ηϯٺ�oo۽óֺQ�o�T{�^����N�v]|�7�4��q�*��ɋ7�x{T/k��Y�E��L�.>�:{XR^�}r]�����D1YYG��V����6���+����L����7��<��d��T��'�EkU�����cpl�NC�*�;�z=�v7x˓#ȩ����w{��D�.���-��>b|�������ï{꿪:�����L��	��u���I�W׃k{�ӊ��G��c+}|�M�s�+�;��S�Ӓ��*�:^5���<ԝ`Ŀ��u_�{?_��0�k|è,��=�Y8�����z��6ʇ�RI�'�u��'Y>Ւ�I�6fBx��Ԭ:�i���;���>�߳?~u����~�><�V�vy�8�2m�R{�2�L�A|��	6�PѾa��5���N%Bjwܞ��M�����2{�ԓ���ֲu�����2��'�=��{�s|��'�~N��N&ٯ(i'�O�_a�i��P<�Y&��'P_7�$���Y���=f��d�T&�}� u���~`x��'.~����vi�K��V>�;t �F-��9/���f*<���F�Qd�E�GGM��S�_k�Woe�s�4=:�wn�d��ڌ���ތ|�Z�8�^�(;�, �֤)"�4nEb�C34u����X��ή�5kw����	�\�'��c'��=jLd�:e��>d�k,�$�+?��ԝBkϱC�'Y5<�$�2u+<�q'Pќ���$����~?}�������/ޯi_��ǤEg�l�d紝י&�'��Y%d��Ԟ�'�f���?2u+8�|§���$���Y:�ɨy�"��:ʚ��Џ���g��W{^?��������k���6÷�|��ԟ2{�a�o<'�d�I6��d���š�+'Xqe��?2q5��I�:��� ��?k�2u+���zf���/o�7�~}��Rm&�S��2Ad���ï�'Xx�ߙ>d�{�$�~d��N0�%�d�6�������R~��6�Y8�+��q��g����B��n��w>D?}1�P��Ԭ7CH2s�7ܐY:��w�>v���I�{�>x��O7�!8ϙ;�²M����T�H~-�!Y8�ú�|���s���ow���4�?'fIěO��2M2Lu�`q������2q�����p�'�'}�<d�&�>;���$��{��M2k��V�?e�v� ��w�#�/����?W�UD��u
��i8��zaI>I�ߖ[$�7�p8��i8�ٝ��	���������s�<a���p�d}��c�����H~����Ow:�v���:I�q���d�C�ް�	�w�+'�~2��N$��0��d�~��!֤�f��a
퓬9�8�:��_a��?��i�M��~������oNv}�}1�Ğ�t�p�f�>b��	�<d��`,��~�J���t�
��VO�)8��O�SS���&��o܆ړ��B���G�~�v+�<?�v~�_��~����p�'<9p��Ğ�w�d��w$:��4w�?2N���2J�$��0��> VN2m��������<��1�ו=��7o���:�u%RH�c�\6P��Wtn�t����X�c�%�E�L�'p�o��ض�o6�2C5en��(a�Ͻ�:��l��.���*�Z�c|�NA~�t~}�#������7N��| m�R�[4{lӭo�V�L���=���&�Z_ϕ���wU���}d�����Y%J���0����ퟒq!��(|��9�!Ԟ��sY?$�I���VI���,�|I���iח5����[������$�	��>a�'��My���O|��d��N���gY%J���0�$�ygRq!����N2m+�I�M�u��	�Ng;�9�������>�����J�$��O���a�I���<��'��S��$�f��f�8��)'�u����PY%Oǜì�%d5��xÌ�J��|�w��)�|���w���;��~�鿏:@�'Nk��d��̒�$�'��}I���C�&���<��0�����i��:����|��:��޿z�Xk�é�I�7�m�^����}��y�=��<J�w����Y6�'����&�?׿���`h��ֲ~d�ja<z�L��$�*{���	�k�!�'P5��&��'P~��>���{�薹Q>������w_�W_�u����2svûÌ�d㴞�́�	룞d���������!YY��J�2O���!����m��/���Ng|�w�������i�{�Rm��Y���N$�3�u�a:���d����s����LՓ�I���VN�6��Y1'�,����ĺ>�ϲ�~�5��|o���7�~�̓�?39C����(|�ĬO9�Xu��Y�;�����߬��<��u���>d�o�I=~I�k$�	�h�d������-��g��y�6o��䬛I���C�?2z�2��u3A�xM2Lu3�8���y�Xu���xwy!Y:�������&�<�p�2xɾ�I���/[��~��gƾ�+$�t�쒰��-6¤��ആ��'R�a>I����>f�Lt�C����<��N2u���:��O�|Ϳ2q�I=����q���}�_S���?�F��,_���cӬ�<ᕉ��M��>��;]�mQX�����OK��iS�;T�Y��m��\��r��y�5�?�Zr垺��W��sB�&
�CNm���º�5X�n�m�t܈���=V��h������s��|d�&�a8�̟~�����N~�*
��'R~d�':��Y'�8�����	�y9���}Hx^�z�x���;������{�~��o�2m$��s猞2i'5d�u�I4���?2p�,��~9����0ݟ!Y:����q��	����|_}�?><�?q��n��~�����i�ǉ<C�d��z�;�2z�|��ì�a�9ܓ��O�i���~d�u���C��J�$�w�+'�Y? ?��-����� �b�y����2bt�r��2|��y�+�&��ϲq�|�'a��d��̜a��;����h,���N��Mw���OǢ�����睩n�c+&Ƕ~�;�=+'��;2�l��m����0=���q��{�a�&�k{��%eC���:�9�n�8�����*I��|?���=s���XNp����-fk��'�;�0������E����Rq���6�Y8�nk�Y<d����u��}�I+*����,��㲇��ЀH�WW�k�Oj��j?��s��߻
���J�N���������j�ud��y"���N���2OS�?2q��^a�:��$�~d��:��}����@D��x��?��e�^A�o�o�)%Nü��N�Bk���N2m+'ԇXz��{���u�_y�_)6��T&�Y?'�,8�<z��q���0�4��I�;��}�|��\����<��~�q��x��ԓ�8ç9�PXOY����N2�;�ORq�{�q�OY=�|I�2|{I�Y:���P���i4e���Oȃ�9�v~�}��o��Ǜ�x����	��p�i�h,�Ou�m���`N$�g0�i�z����N2��q���v��P=a<}���q���>e���Њ��a�V�̜m���u�gQ�tx�6��B��g@������[�dB��ե��v�l1!/�+���zr��;�,x�*vs��7y�d�T�u�&R��Sv��7��s�&w��vao��8j�Z����4n����wm=�Ʀ��k�P�C��t�=��ߩ`���{����~����#�*~���Oƶ`|��MO>�>C��J�oY	�a��é����'�XO�w2u���zkܓ���5ߍu��m���u�{���Β�c�P������YS�&٬��'�T���:��~����'R�4ŷ���J��	�a�9�_�'X<�Y9�&�7�o���?��t/���ݕ\k�w��������?}?Y<d���%I����z���?�k,�~I�hˌ�hu4~�C�,%k�q���y�Ru����{ܐY:�c��^9a9�4�6zW3�
8G�~�/p=d�O}�$�����+$�=�쒰�C���+'X~����N3Yq��'_���i�c~��N2�	�a�ֳ~�����}���[�����~����Y	�k=v��&�<9���Oy���q>d�u��&�̲V,&�O���Aa��C��Mad�0�9����r�}�O�[5n���sVg�(�~C����|���C��Y:�����d�	þ��Ğ2i�����:��'����&�5�a+	�9�J�������Y��]9�Ƕ�l��x���fo~�o��2~N�Y'z���0:�I�ל�q����{��O^0�w�d����ÏRx��uܓ��M�����a���� ���<���u݋1��������ȀHN�^$�<eI���q������g����R|��y�2B�2u�gRN<a���L:�9������@��:���못��S��~�1�y����iH����N��a8���*I��*O�Y72���d�����q!��ɧ�N�q���0�xɤ7�>a*u�ӽ�ĝI8�����/2�4�|�=ߝ﮳ޘ���g;��u�h,�9�:��5�a��u��y�T�'_�YO��*N2m�����ì�d?y���x�����u�AU+�js�o��-ze'{���@���k�����E���z�w��	3�`鶀}���j�]�gy��Ÿ0:�K�mgvOA��2� �PG^����\8Z���kHs^��%�N�%���˹f�"�P�x�b��K*���^�\�x��j;�;����}�<����x�*V��aĜa15>�d�]�B��M�a����������<>�$����7�,��l���"�t~C�7�޿��k�Gɰ<N�qy������&�x���@�4��<�}�a>aPѾa�IS�Ӭ�A`l;�Rq&�P����OY?{�I:ɯ��+�M�9�	��'SF}�w������~ӟ�^��}�bI���7CL>a?�Y�M��&�`z��8��ϰ�hu��PXOP���N%B|wܞ��M���,Y=d�{��$��Ǻ�5��s�5���}�=����!�Y6��V��O��,6�z�3G�4��O����4��(�$�d�������;�:��'���0�'�;��Y7�'s�g���s>��r{��>s�g��y�����}I��0:{I�R~d�5�g4�2βOR���I�&��?2q�^}�|�:��oX�:������$�����?}����ֻ���3^}w~�ޘ���	Ӽ��N�st��d�$���d����Ԟ�'�f���?2u4e�a>aS��q�k�Y:�ɮR):�����k���ev�΋3߸0������t'���|���:��ԟ2zo�q���O?k$�I�S5�Vd=ed�!�YS�'YLd�C�����}�[�/�x�����������g�̚J�����I�T��2Ad���~I:���o̟2x��'_�4wY'O�S5�T�H~-YY8�'�`m�q>����ߵ��vNu����R�����G�����L�gp>d�V���������,�a�����q�I;��4�ɾ�	�|ɮ�!Y&��s�IRm!�����^��y����s�>7���g�+'�,;lP�ԣ$�'��4�1�3�2q���^`x��N�C���|�k���<d�'�|�6��Ě{�I����5���nhȨ~��B�|�s�g�H��ㄮ�签��|�y����q�ݑ�[��.�	��{E�����B�%���$�Ryu�a�]��6�q+㘚���+�f�1���#�Fͼ��V��bYK�j�j&)�ZYD'�;��N^���I�}�7w�|g~�B��a�'a*
�m
����N$��|���ȯ��8�{C��}I�3�a=~C�~��OXM�u�'�>`s��9����	{��j���G����>���c�Oʤ�i�S�`,��~�5��(L7x��u+'��q'����O��!֤�f����:ßS����s[޷�������]>ӭ�c&�Nt�Ì�I�'9��4��x~���w��qy���a07N0��%d�2��d��5?XN2m?o܆ړ��C������s����}���w�{!_i�y�6�Vq��;��:�9֘�Ğ l;܅C�&�Y�����N��:�Ӟd�*I��+'ΐ<�'6��Ի���{����}{�~�VM!>�}d�'�t��!^$�oy�IR���a�a14�M$�
C��P�'�,�ԇRz����#�`����ﾆ�l�b��]���������O^$�������>��,6��!�י<}d�zo��4��<>�:�*V��a�I_Ӽ�ԜAHk���N2m+!�!Ԟ����}��t�����6Wn����V/��������>�Z����<}d�h��OSG�d�!�^a�u�Ĝa���f�8���0�hu�����J�r�d�+!�g�g���]��t0���O���
??}G�� �z���{�I�'��WI:�Ԭ&�~eC�'��p��L8�~5�M2u'RoVO����a'�u�9��ϼ������۞p��$���d�VC]��d۴����&�?׿���`z�ֲc'ya<z�L��$�*zj���C����YB ?f����]���޶�����k�q�z���~��N��9�Y���<�0�'7a<���'Y8�'�� z�z�VJ��|�����qL���'R���ԩ��׾}��{�uD��:�XX�&��D�樹����Q;��ò�D�SN����h�bQ��u���(b������ĳEJJ�X�FD>�&�f�8�^���ȧe����W,�.�"Ι;�[�=�r��L���\S�{���:��W�D� 5}y�9{��7����׎�۪��l�hlVd���K@�M�ZoA���6�p2�kA��9:U�K�����X�Y�y
�0 �d꤅Uր	��(��b������gvȰW2�k��K���a���:�o4��ޕ��%EX�F�!/(����nr�6%�/w�TZ�;K�q	2i�9�彣@�
�Ge�tfU�A�j��yC�O�YsG�5�:�N�-�:�q��;��:�/Q��B�e�8N���W5}���5*E>����U�f��
�@chq��_U�7�VQ����n�����B�n�JM�Qp�ep��n��t�N��u�|�od��U���ػt�h�mZ5�d�{]�̮�u���t*���G)ou�ʱ3+p��*�Zr�W�*,j��U�r�
'G=Ц�kz�)�&,&���E��y����|Z� j�:ɬ�v,SZۊ��+^P�L�0����T�ymۼt[X�H�1:�Kn�ʒ�@�C%��ת�,b�.�*�z�
%h >'$/��\#�\9��T&�N7����օ0�Tgk�W9|X�/ld<�4�TX����)
U�x���XV5���l��H2=z�"�|d��W���O&5X]���
�U݋siuk��e��]��[z�C�{:.N';4g�����Z��AE�=�������%�'=��
y���Mv0#Y�-�X�0�
�,�҆���ۏC���]�QbWd�O��1�pu�QR��L�"�S��y�!�ow�l�z�O�F?o���ƒs�tWl���\D��|+��I�"�v	�{f��������ݨ����W$4��k^4%ow`�ۏ�U|0N�8�o,����]�쏛���67�-}�.�7�sh���rݵP7i+�S[j/�}+t���Q�ʭ�S'j\@噽����}��_ nh��
�PTL��:��X�; ����+��f�a�屵%�� �X�hI�b��E���=�ٷ��J��=[�DD�M������ڻ����b�",���g�YZ���R?�f��|ᢠ�N%��v�I��O@[�]�͉�e9۰��Գcmo;�۴�(ʊ�gqU����Y�џwWI�� {�x�N��4�M�ǽv���P�-���Nޕ'F`�.�w�Z�#FiN�u�m�C2# qM*UvS�%�`�ڳWb�r�`��'%��[KY�e_=�������j"��Fϋ�E���vlT�2�}��N�ֵI��ѫ�m:�EJ딢�E:O~��6s��
M���9�^�V���t9�̜�^�O����Qy���<t0��o�rIΆ,\�ע�U�ur��W�b /�-J��\��ZԨUX���U+
����-lFEAR���3\ˈ�)�EX��R�D�erت6�L-Ƹ�*(�Yim�(�-dEYiE�+YTm�C�F6�hŊ��iUTU*TY��ƭ��Eī��m(�LsJ�����* ���b�*�-��&3b�iPQb���QGF�U-�PF�Ur�ՙKQJ�X[\�8�#s�R�Uť��[F1�j�h���Am�&%dr˔̣ڠ���e��䱴Z.e�q�#�jʭY��m��1�X��[j1mAk)kE��VcI�m-*1)m�XۙLfTq)�0-���-����Y�*��F�V�+m��T��Qq2�C2kcJ��.Z1b��F�)�[eTe��VTe�U���(��\l�b&���EFұ�[+��Q��l[h�%DĨ�bL���S)U8�� BqL��+s{'�܎ZQ6�%˶���G:A˶���r;5��]W���	���1ki���(ef>�=՗��w|���n��$�n���DG�i�qC�A@��r
N�u+5�p'ug0�4�u��:���	�;�a=~d�~�$��u�k$��`~��Ҳ~I�{߼gW���<��ٜ��>d�����x���RN��P�'R�<�"ì�Jϧ��
P�w�;��u���u���>d�o�I=~I���8�q�s�������[��5��;�|��Vd;hz��ğ3FR!���єēhq�?o��I���!�N%`h��E�Y:�����
��?�'wI�M2w��2i��>�ϯ��o�?w���߼���O�$�5���i�o�IXm���aRq��Hm�u52��|���������C����x^`x��N�����X	�~��u������9����˙�x�d��I9��4�I���'�MwY
�6���$�(M��*N ���>I�N���O�q?����a8�~��'_R�׼~��nq���M���d�����>�O�R�����s:��M$�d�N�x�O����3L��b�8��5���z�_���)������Չ�`o$�f�Ӧ���#�N��%�ޖ�ʖ�Z��K�U�gV�讉;�L�e?Y���pY��K��}Z���Z�(���^���	���K�Q���7�gq=��(���P�͓�6��&���Tŉ�<�m��X�>��Et#���0C�|�o�v��uZJ<��&���R�U�^��n�? �]M&-_$�c�!y�i��4�g��ud�cҍEG���ZU��]��*D�ڋ��7�����Ww>���)
ή����o�f[�L�9���22���G5Q���W�8iY�Z�JJ�um�,a"�����u�y���_P�&��\s
�X?�3O<���u�z2�W��+Ǖ2�Ƌ"�Y��<^f�Q�Ǫvf�W^������a��Q|A[�8���]�׮�t�?_�g6bm�[ՙ&u��&���{��=��@m��_�(%��\,X}Qo*�/�{�/�j|۰�����/�D��u(�cU�̾=J��Ŝc�=��ͭ�süj�^���s�6ܿ�r����8��mQOv]oӫT�}zx>�>*��ʽ>O�q��X������$7���9�f�)v\��%O��ptqg��{�=�gh��o���W�U��	9���B9�at�<�v�\f��T��d��k��������5����]�҇Q�܊��]n�í�0I�7�XA߷�>y;0	�G|��b��:��������ʭ����y�;�}:����$�ϟ���9W!]U�y~�#A�4�M�`ZWR�X�c@��=gf&Qw��m⽄��vr)�.�[j�Cg
Tz�fͫ@�*]H��g�Z�j����}��V�M2�y�At�s]�zJ�&,٘<&��-ZN�:m�Պ�w^Y*l�����9oO���|��<�:x̵w4�H��l���g��������E�r]-墸��A㛸�����"�	Ϋ��7����zX��ë}�or �Hu<r���-�9nX�-[�Gٹµj�\ȓ�z�K8!�����|�Aa��I=��XxLϥC����q�����N��Ѡw�z{�}��9ϓu���3���;�8�h���q^�G�ϭ�0�z�5˻>Z��t���/эO=9�Oz�=�a�l��a�3�z8fv�͗�����^k���.��"�5�:�o���6&���X�z�R��ջ���mfֻ`��&����m�������3~5�S,�;	î<�k7_��շ�/�5�/)p�,gs�6�2��vT��~��ws�ZR�6dΚ�{�*��u}L��|9h�3�G�d�wvS�^��
�\=q�;�����eu5�Zӣ����ɥ�(uw9����ݵd叻;q+�g!WB�q0y�V�:��aU���2���Ioj�W�0L�B�;��NԱ��_K�J慔��Bʰ����I^�������~����.s����a���Nt���{�^
����ϓ'`ݻ�]ܙ�������̤EI����t�^�y��-��;G��|�M�uMu�y=���]Sr��G{�ޓ&�������������1��hk�le/i�aϹ�8^�����{�&����5"�w4�j1�nNuֽ�fW�h�6�>�C����������y�g�+���Q��9z��O�j}v�:vB�a�Ϭ ��!v1���o+�����S�x�ǟ������I|0T��aӲP�x�NuX�o���xo���ݑg���Fz���dy����IW��y=qw��έ��hSץ�b�9��)���g�,�>N_n�~����_�[�z/��;�՘�>�*�5�����(���{�uo:ro�����T���쩷���WHe�=y���������1��Y�'�xp[V���Q)��E]��h\���m4g^��S����]�:��M⓬o>B��+�%��:v���q�ҍ�V��j��6tR���U1��*�룇��٠��8�����S3��}��|�vtr����܍�~��Ψ���|��N�ɏ�gl���N]����dwj�I��U�||�p����q�V�~ߎ�l{�&f�w�_".����U������O���kt�nf0&f[<�n����ǝ_�q�����vx��,�!kEXou�����#�f��w����P�v�R�&����G.��sI�c�
����G,���yǚ�c
̗_{o���{͆�ځ:�c�k|7��$7�A(G:aq���z�%�r���^[�7�;uBu��Z��6o�I�dɮ��7Ⱦ��gl�WK׎t����XòXK������|^9�r����x*��w��=��7����ܳ��xeoDF��t��4�*-�M�pެ�����[��S��yy��2��]���C�/�s��&��j����3op���2�Ub����*��N�����iK��R0���-�M�+;/w�e���X��+�5d����]`U٦��M<��K ������U��	�v�pp����)��r�#�2��:�C�v�_E)�t�]s�����m���_}U_ߴ~����գ���y'l�<�J�t2�Ix��/�|��~g��}��p����K�8`]��������|�d�� �����c��y�ꓗ��[g���M?K%�a피�gf��t��&�r<��wC�>�Ro�s���'Eb��}<�����^7�O�ݚJ<��2z�C&��o���࿛/M���Ժ�'<��t�\]n_�Wq���.���e��N�HgAV9Υ#쭞Ɯ�K;��s�Y�p�p+�||�{w�jd��V��A:�d�B7ٜۿ��G]��w�i~��^�9ؼgOu�.�_M��O�d�Q�̿,����nQ�C��,39f��Fʶ�ԏ:���1y��϶�.T�zw�\��e��Kb^�#h�v�V{"�(�N�^�g�(_��Ho#���ٴg��3���jg����Q��X��QTv���B�u5\�Y�mk��\�oXs5أ�'�k�����H����2��̡x������T ��`��g ��C�8�>���Y��P�k8u��
���Xߖ��v�b�f?s�����M?���6��c{\�Z���q���_f�.�N_���r+�)ouK��x�[���(aMN�a�d��^�����o6��ӣ���b��is\����VX�0�vw{��{��ި{�|��o^��$�K;A�x��=V,g�`�i�T��6�ۨ{A�\���%��|�>>�Ӿ���}�v���(c'��R��'C���|�M�.۞�*>������ԋ.:6XĎf�k2�{��}�v'}9	c3kj�ٶ��^8y��=/�o%\b��R4�߻�^x�*�l�g��=w� w=b`�����%쥜+V�r���b����N��nZ����1�S!z,	&ؗR�(p�{���W[}�A����5f�{+��s���wBhyƤ�4H^����;�}��`��o�N��V�<WnH���N�����n��f��:
��pR>���`4��_��q��z�g'5�Z�!T�ަ�چ�nn�lfq�%��pWv��Р�'�Ṯ"��qRy���f�Y�=$��oh��[��x]n��gmվ	6���q�b`�u�6�7�n�Z��ýhv�T�DV(*�Jq[�ePS5�9>���}�|�׾ys�����
z!G<�J�r���]�>�%��G��	�u?bWYw|��ZN��:��9|�g ��8����\<Y �����9�������N�m��ˁ^Wk�q7`jg�u|�ȗǝ)�|/;\5��N3��_d�3�z6����������	�;���U,k��]�{j�Y�g��8{�{8l���8�hA �N9�΁Ǜ����飣�>^�������+[㱧ۉ�s���$7�A*9�vnh|&�j���wjnzr"w9|��x���_�G`V�V��y��8�;]���f����+~�;������%����p�~��Z����ľ~�߼�cy�fK/0�'�����Iv�ʔB�}ψ����~s_��uh�����T���~V`s�ד�Թ��?d/��is�A��.�x��Ygv,8[h߹��RK֫f�[��JT��q�i��sc��*(�؆sm=!���Z��Wqح��O)�Zw)��)l��z�ek�ܥ7��9���#�����;|�lE�	�`c�*�"�@Ѿ'�]tokEk�3��7����X�d�vu������rө�	٧+��oL�~���{�K�'�Xt앬��U.^��[�(nw���n.~;��j|��rdx"���ܛs*X�7~㗗�yg���������0���]��	���ILo���x��9p��菡��Xu{���^/~�+h�C���=���ל��eJZ�攨�^�;W:h����j��{��8�=�c-м��Ṷ�{|RC���6�yiR���[����vbYKWo���^�I켷W�rR�F��U�]����y�rq�ݓ�}������u|�3�u��n��r޹���@.{��X!�<+���cۖr��ǹ5ǵy���4��ʧ��w�;����wQ�2���s�6=����{~��]�r�s��Z<�|ϥ�c�^M���Y��bCc ��y���sj��N�Ο/S�/����=�a{Y��]�"o�]^v��]��dz�3�};C�U�G�Mn��[���eY��z3���H���}������˳n]���❖;��b
���)�{�#j���m �;�z6�� ]n�z����=T��>��n_E��:Y��~��+;_v�d��l�asg�I��&oV���:3�u�vǊ�U��q�϶���tv�(��\�
޴z<y��#����
��{�᯦o;ɝ�y#��v���y�s�7����!�����ߺO,��]�/w��n<��&]N�v;!oD�W?��}9z��z6������\�ݹ�zZ{�Y�E�RV��۽#����ٵ};'�z,�&6p���O}���3�o�L�q��*{���c�tb�8���Mv�A�(����`d���Z{*��t3�d�l;��a4#��=T�o3;!ճlzUb�3E�Z����^��=��s�s�WgL^UX~�Y|s&��oM�S�g��5�ؐ�o���<a���}�gs��-6�*�o�ƥd�t�z� ����Ӎ���љ����ϖ�l6_^��ՙ���lF?#Ƚ�����WgEb�����n����jl�8_ �*�ڲ>yl=�k���녩�E�/c��A���]j�T��}LK�Pۼ�c븸gN��C
�	����e,9�T�L(z���Y��r�N���5�GZׁV\9����p/0���p6�I��o.��������Cz��Ag	I�n�V_4��ɻ��[N�]�p0�o�>:��0�>V�vo���k��'v�Ơ��u��y�ƭ�.��4�g��[XD�x��0��oCѴ:8}�!.#F�;�N=�Y�tr��R�8�Y���R��|��61ڱ��{{���i`N�X���iS������p����i�x�n�ާ��"ߑo��i�!%�v�ƪ�Bث�4�|@���[Ֆ{-�n�e��`N�
�!#B�����גG&�,�Ԏ��ۜ�v�|Lrʕ�����{3TS����ZJN�������	�a����߭�8��ܠ���mS�tb7�T�0X��-��7WөNU����6透t��i��]ǧs�k��7wz(+��<��l��*�l�~YՑ�B��.�{�W�G�n���+�.�[D[�ލ5.$�v��Iޫ�w(�j�k�v�C���Z���p-�."K��g��3�C��{t��Y׷��F�I.�V0(V�aVك��h��,R��NbV�p*�u
����[�s��P|M�g u�س�̾쩉[�P�Gj��9u��l��$kp��*+�<O�o�Ƽ�n�%�r�/u�=�%��Z,�ۏ8gV��!���ś귧^i��](��\4�!��ͩJ�>���h
��6�涉 �(.Sz>�5$�C��WC�+v���RWn�аN\�t�\mdT{����5�|��uҰp��/wi+Y�S>K��I �7�3�I�8U���Ph�ݐ���u�n����Vp��yS��1����5�լL�q�ѧE`t�qྒ�`��N��u�r��������lL���1VU�5�a�[)�C��ħA�WjU�R�O�K�[҈YC(��OgZ����J���7� 5`7�JXf*��nr�V�g�TA72K��1���J��}w�ˆ�r�Nv���rw_j�)=��׽��dH���A5f�����^�;�3g��Ц��}a��d]:�����vR{9o0t,�`]Mr�ӗѡ��z�%�����ev,}���|�E�8�c)p�X9�����X���&�\��C��[ًy�
�˫.�9@�CE-u�:b�M%Vu]#f�C��W�xb.��Ӷ'|�"d��H�4reuob�Ed��`f$�ٱ������:�u�X'.���(�)�����4V��j��S]�rBq��]=K,�_u�ƎV�=9\����:o�E1ܤ�U���|]��<9{�75�����C�YmAݍN�"` h��QER�#j�˕Q�ڕGI�
�j� ��aXV��2���U�˗%b����)X#�66�EA�3#�R[bʕ�֢ZU��j���b�A0��J�ƤĭB�UB�2����c��b��̦V��J�Ң�1
��j�W+��Kps
�*a���&%�-F���IZ�aj�*1��[VjUE�Kj���Z+J�W)\�QLh1V3)�cr�G)U �EZ�`���1[E��V#2�cYRV�c1�P��T��alX�+E\ˁP�8�-Ƣ�[s*2��Ʃe-R˖�j��c1eq��ҹ�P�\����#�Lep��f2��UL+im��k��ҩYVТV�UU�̩��E�U��m�������[��~}�w��了�m#M#�p��UwS��d���;L�vw*W�W0&��gK�>������Ys."9P�����W��W�C�$�,�W��Z����37���A籙���v���k
r����3��;�D��b�ľ:����n.d�����#6'���C��b����W�Ǎ�g+솙�)�WLP�1y��ϱt@�Qs�l�Y�+9��~����흍>uu<7j��T�aghp�1!�l�g>�r����g?E��d�X���M����=C�b*��:��;N�[,
��7��ҷuR�s�:�Y��ϼę5���`�%�����c�|=kG=�J�y����*Sm��9���o^��@������kn-[~�&ŗLJ~k�7o=�x��
���ݳT{�^�OI��5NO.#&R���γ�戼<N����.��K���1����˽W��^,b������:�c���"Ƴ���O���~g���oǤ�9�N���-�m�J$��c��x�+�����\��6�
��D�"r�`�|V�霸,\�\��^Z�T���ok7�Ʊ����樭��KiZ:u_1 [�ZX{n�_��%��Æl��זR�����ItuR�1���GwpCg~��ﾯ���3A<s�?�5Sp7/�	s�&	N��x��h_Nw�`b2�t:�X���p�yMo:�$��C|�W`@I1Eq�ymlG��ן8G���[����f���y�wB|�[%�bB���=A�v����/gx�G�8J=��e������n��ٴ����	=γ����J�j6��y�{����� g����S���\<nE�}:�z�k1s���
����x����i�ԕ��4yu����5�br��-O��I��g�a���Ґ���M���Ñ#�5rU�3�T�U�Ge�Y�����v:��#�9��3�e��S]`���\ʵ�"�e��iwo�t�y��HlG-9����ǯ>�{aY��3��a�JSs<%���u]�Sn���>bC�d��t�^�`���-�
>쫭*I�Ik�F׉^�� ϼ]�/�G0L�F�M�|�
�u���m��m����8�볔���a�	����S�V��Y�6�fi�K��\۱zx]��)��xy�_l�E��o�Hވ><�1w)X�U}���b�� V6�=�������F+>>3� N��Vk-�ZZ��G�/�$�N2�v�Ϥ灘���Ykz�|�r7��c�>�h�e���޵��l�`���I����[n�K�K/�x��׮Ls/$w(�}(������[�]��5�}s�N���������s�;�侬:��aӲ5�O>���݂g����ղn̋�G��w��ϥ_�R���eI�A��(>�y;��eu,�Ӵw<�}���v3��3,I������
�nM��T��۳��{1�m��/x���_�>��:�ލ�/v�ȯ�-�p=���j��봗�������wNǰ�6�<��{4�y97Ƥ���U�-�L�����vS%��^�eW��M9�����{~���5��Z�����1�{M�t�k����n=�W��:���i�T�a�K�����Ss�Y�пP�<��(�G���1F#���h[K*W�
�KG��&�V���@��Y䷓/ ��@�p�Ť1�R�ID+9��yE��;��6ʩf�ɹ�%�WU<爇�Y�)ݦI{:��������»w�xmZ\��7��|=(�wV����&u���@�^�{��M�	�x�����>�1*���,8���a�Y���b�^v�3m�	��G��֒��~�����r�tH$�Oc6��b�:��谰N�h�IΈ�xV�~��_Խ��%G���(��y(Ⱥ��N�Agm �Ju:�����s�j�o������EM��Dqg�s��20��������͖$��V��q�5~���þ56t���y�v�v�����a.voZ����,ݮ�N���[V��f�{�p��w/v���Q� 腼_��y��p'�C�c���������=���^L�/λv|���.M�vL���h�=B��=TkuVM���}.>����Cxt�W��u߼��yu�����;�Id��a���W�=�����3�o�H�>�*{tu�]�+;~�i��v"�p��r��uG>��43����m�@�o�;|w�����k���]N|�CZ��ԎM���ZN��
�W�C��m�o��mA����%���� ٺt@��a��Y,�#un����<���ՃS����ڦ�+�I��| ����󞣽'�V�1�H��tM�=��{*�^u��a���	��t7�⃫P{7"�Mr�U�^S���=����G�g�|�׈�we
�rªœ\K��dr��q�+�`������5NWW'�z�K��9�7�nO}�����z�4/uＹ٩唵{j/�d�5�w�d�>s�9g�2���+{�37��5��z��?u���6��f�5L]�[;7`^��mf��C�ί�9n_k$��w����b�I12���Kn?rfuߔ�_��"�@u`+�`,��zS��wl����;�YZ^wN;�l��Og�8���fw��_�q�/X�����ۅ�)�A����~;='`	�7��ӝ0��l����Y� ��y3Y/���}ʻ̄�L��R"��s)�����Ms����u�;N���c���ˡ˷]��Pq6�ݎ���R
�yp~C�N��LsK�crw-����ˠ��j?�R�
��"쪥��p>��z��y%���L��n���o\�o�sj�6�t^j��o�|�\��i�-13�. �����7�S�}� j�V߯yƪ�~JmӖ�6q۞�`A߷�N̐>�v���.%�AǼ<}ް��OY�t_
�y�]�zG�zk��G���)��HU�ɋv?W�qٔ6�_l,�˟XC��.���)<�U�(k{��Oě��n���7�=������;�!<;��յ`��W�c��ձ���B��m{���j�KS���%��(О�Y(k<K�^����+[�%�o�+&�<��i�V��ڊON�7�J�3�&K1����0k��ρw��63�����xW�C;7'����MyƮKbB�w�t:Va�ߎ�Y�Bs��=�[r��}���uy���c�q����'��ꨫL�s²W��]�o[NK}n��|�y�.����3ظ{�"�5W�����J���Ju��0�=�wO`�kvӍ��:�<�]-���5�}�̃��zJ�Hk\�Z�tePh�%P��(%�WzW.37(��"�� a����a¦kXS{M����g���xyr��M�Ȩ�"I���s��9O�9�l�3שPkZ�9v��$�Sa��:�&�9��	�Β��:n(iQ��Y���}ﾯ����~>*wd�/�F~��Jw^�w��T�;~J�8�<�HU��{�7�/6I\X� �vW����?M���gN�����z��~<cti��L]9 x�y�K��|c�(\�1!�G/��L.?w����[�G_v�p������{S��Yډ��Q�լ���ls���boǫ>063FNj���p�Q��m���r��J����E�Ծ}�1ͩsۜ�<Ql��"�#^kfvKo�'J;���|v�X�#z��E��.�7��=amm�Z�����{σ�����^H���e	D!�`�y��:WۜY�T�YZy�,yU����}x�)��%OX�<�����[����.}��V��y�X"�r�+F(���<�U��5/d���O\���!j�T�-�
���t�����X������z�>f\���|��[��h#��9�n����+�xѡԻ�/]��͗C6��S��|��t��9>"ġ�r����/r�'ڌ<�l����wB`[+6�8�����B�I�O�p)���X�W";$�Z�tVbΧYZ+/�7��33��W����w~�������_<Â���L%C2�Oe-~�;7��2�}�-%`����L�	��Y�}��_�����Y��H����ym���^L��츃�bV/_����n�&V�qP�c���1{D�W-%E����[$�i��~�'��Y����<�^� S�<���Z�S*�ӆ�i�^�P�������az�,#+(3�r�lU{VeS=>uS0j�=��inN�(�T��$��r�t=E-iǲ�Y3��|�Xl��y����PҬcn�ǟE�ڴ����)��.�9�]B�	�pK��}3��Ӟx�'��gXS�����v(�}�[)+]ZVT�|p���d�M��L�������1v䳖.ߘΆ�c)��	���V�*+�i�Ze ��	ĎpQ�=,���fcO���M�	������6���9���\����6GRv)Pן^��G)2�=2xU�QD���{�rw��e7��t���j�_�6�锏\�G��j`%�KH�i������V'8^i��m/r2�կ�\�kͻ��VGR�`+�5Z�7��88>y�:�7��Kf�z�rNy�����xJ�/�z��^촧��Q�<u3�f���:՛T'[�=g� �t��u'Ǘ�iq��欄u�YV�¥�+��02��9iΉ������UUW�n-˿tsUZ~�S��^	af{eă���L��VxIl�G��f��t�8�m���=T�m�(�A�[�hN�Q�2�*��]Ӽ�g����1�Y׵�>���/u�ˈW����r����1������,��F��Y�����<������VT8unٖ��o=~�j<%��i*�H��S�]�C�;lOΑ�\g��yp��c�VOO$WS�M�}|���J^}Ρ��BX-$(k5�YN���w�_�{���}�����(�7��煡8��o�PJe��5V�9!�ȑy�͏�	��`�ʳ��!�5������V.�s[�7~�=�h(7g�(>�jT�d4�,�mY��������e?7����J��r��M���/�����A���p��ofD��&uuC����]c,���Y�5�V\��˧l揄�>>�+��3ר�P-�����=��Ϧ��ܱf�����Ue{r�I�<S2f�5�R��޺���%��M4t{/L���٘*]����MC0$�Q�-���5��0�/|���7���}F<>�~� .s]<ܕٕ����K4w��˹�"iv�����skV��	����@T��12kй�ת*7�
���*euֳ�w�ۮH=z�*�ƍR�w���]x�No����M��ΩR�;V~�o��ʇ�����W�#��,�*��抅��ˋ�K4�';f<��0��v�g�8��¡;ݾ��Ϻ�х��-�R�B9]i`����p�;�R���u�^ěKS�XfX�s�>NX�-�a�yl�G�ҡ�����H�7��5g\�ӀpS��M��&��ъo��&96�^�)]Ʀz�n��`s@�kn��<�����g��Y�K�G��-k����M<�ǋ�ᜳ$��Xu�G���'�vl~T�3C]R{i,�Ŕ2�y��X�C>S.vֆ��sӊ��_Z�p�'��8��=�^�c�!��Z�(���e��)�w��=*�I~-�jڰVX��s���O�s�<|1��7�=s:�/�^@�	������sР��X�bQ�Q����	��c�Wp�[\|��u���&D�`k��_Ԟ�`�J���:�.W�x�3���9J,��VD��탂CP����ne�J��Vjo�e���s%m�m-��ցw�C|��M��6� 0��:ji�Y���L�/4�q^�-�w�j.���k�)r2�f_onfr��G;mo5VYb����O�混��Ɉ������7������ɿZ�v����)^VEL},�5���/�W5�7]v2��Wj�oy�Ta�ǂY����Iԛ|�=/A�	Dqi���;B���[R�t5�k�\	�����b}np�A�st��Tx�����O���1�;&pПnc�W��<���R�A\�#8��]8��HN9]h��]�h�k;�|e�3�m-���r��v�w.J��� �!������Ρ��h���y�h�U�W��o+r�^�L�I<���L��ǽ�Z��M]}[B��|��L�]֨f�[Lq�s�w�Jބ���u�Q��L"�Ҷ�3i�\��N�W��C�k����4].�"�}2qo�+����X��tk����;��
���(�w`� �6�w�mj�k��!;�,����A�`��a��z�9e���Ʒ_�D�Tn�h!u�S^�XY��s�hU9��ig>�w�[s/E�1�m����j��&�;�l_>�u(�0�d�[�L��2���;v�L�yufl!T���]4�U�-��t�LJ�d��[���˫�eq߈��pBD�:J���U�1�qX9��VGvvQ��������r�z	��ᡏ�U���t^:9%a�M mwe���;�X�8�rF��n�b�`�,�(��.I���#Z���y1�X�;�RA��؎
6�6�ۓ��'oq��.uӔ����/�c��b��ʳ>3��=�7�oR�L���Q�������Gn�-D��F��L�*l�/�%h�NlU��C5{�|Q��o�Jq�Q"�t�������=f����Vm[��%�g�����2lA��Eά�&�t�)ef.�w��`ca���I-��ۣ�-��M�j�N���l�bI7���BD������gJ��;��>��S�\�4������v�
f�T��7�fHzd*���5]�[Wݴ�`}{��A�-��u&�����f�;8�lso���.�&r�H��<��y)�i�ǟcZ���ս���[�hY�U���sn�<"����}9}�f$9�P�����c��ԩyr�-��n����{:_P�%�8T+m"���״1s�/�4AC4r�k]��z�n�'�{�-[ݙgye1�ud��;9�tf� Dt���2��e�6��/�+-�&�ɑ�Æ��4u#�s������ls.�+W�.��9�����U��E:i�NNᨵ%�s��R�d��0��D}�+t�ь(�h���ק���nV3��F�X؋-���6�`<�`U��8�,��S˫T�C������95Kxxr[m�it,l�Ǖ�*���ateg.���f\:w�;��������>?FV5̮&RԹb�\���j�.&1VU�DA�Y�TQ[ZQU�ң32*����Zҕ�jQ�pl��T�Ys2�J�kI����[[JU*�arԣL�F`��T�ȥ���f\q�iSQK����2)�1�e--q�BV()���1�q1��L@�T[qr���b0�TX��k3,��H������HfS+ZR�s%UK���ER��9J%�D�\E-���9b��3
�0��e
ۘ���c.,3�����q
�㊕+X-����V����`)V�A\kUX���Qb&2��q1ʒ((*���B�e�Q��Q�1�1��WJX�Zʭ��H*��1h�+D�YZ�8�D�2\��f�"���e���[q�,�U�"K���,Ʀ0�mKK���U��̱T ��)��Vf�7�t�W}Fg�.��)t�Ƹ:���^�o��r|&%��-�/�t�E�h��7����%�:��+着���7����������1���`ߕS�<�� ?��'��{�8@{}n�.��Lj��Jkپ���zѳ�P0��Ƹ\���ٶ5^�i;�X;1�O��gjIsyZG�:��:� �ޡ�����s�����>��s�,{mJ�%�ȋ�S0�񰄻�}�޻���;����Ɏ�b�}�>�{�/:��|]�Nq��x����#9���^�>���qYӞq�3e��^>�ۢ����J��X{r��]�|�]�tV>�.����nc3;�����=S9xU󏅉�xn�w+��O��\%���Euܭ,-)��1Bc�YP�s�	˚���x.�#mq��dH[u�ם��^	�Y0�6}IW�_L%^;��Ή��Db�!I��t͟x�G8PM���J�Uf��� Y;BQ�å"�t��>�r$ve	��N�b���y���Kj����O*�V��������hqDiϒ�6��3���S�GE9sVܭ}���(SW��.�κ����$ŗ��CsX�ѝ|���y&���$�NSWc��W}��u�A(f&>u�}ںf��h,���Fv E9�4�L���*�q�����QD�m)����6��HK��2�.x�ży�����}�D���9��w<G�;��o[����y�K�R2U ~� $�Z��C��as��j�]]{��aIq�u�(���bU�$y�{�^5~�l�L�a�0�5ґ'��dS�7�x��g��L<e�E���)�v+���W���T/V	*b��r�ӓB�iQw�� ����v�,��L�3�R��D;C}�!~�5����������WcK���]C=Vמ]�wL�Wj}R���$��f����-��5G���a�{v"J��U�N�=潉:��.t�F��*IuC-<��$;��g��A�������ϜR�p��_�=�4����{���S�EO��	V����'��g�=k~G6�+��Ǎg��+O�n���R�x�㼝��m��ȴtO��ʋ9AF�ϧx׾���O�۠���a�j_,����{^�����W���nj��f}�]�}�cbϢ����m,��AJի u憗���賶K�(a~�.�"\0�9x9�ߨO����J��ł��/��w��;6f���VyӖ�ˮzக+�T����r��c7�.A��`������qu#gsc86T�{V-1f����f������}V�E�{;�����8�|��`��'N��F'�Ǆ��]��ۙ�8���d޻�֣�d	Q��$x�Ը�;7�[}MN��W�W�}M���e��|z�1P~��ZM����������d�O�fp�/����_uW\��٥����r�α2��VF�MX��O>�Zf]|)Ď1R$Oi���E����p��D���;���i�kX&T3+-r��I���ܘ�����y{=j��~�ʮ��0�h�RAZf��c�5�2u<O���L�zĻG�������ׇS�c6|�g��y������
��W�����ّ��:c}�~��'�#C��Rb�KŞX��dc���/#L��2��DN�Q�2�{�3�w��ܡ��B'�N�|���=
���9M_���W_m(�Lƶ��P�l<	��S���~q��|�ÎR�.�Ys�,�ZU�u4�Z��Pw��IP�H��S�]໇�hO#��L�Z�Β�c�N=�o �s�as����K��r�O|;Ȓ/�W��;QhKa|}�C��������y�{*V�>ʁ�h��/�h�
~GB���!���v4T�E���<SF
�w�ʓopV�B�.XzՉ�gNC�MغPބ�Πx�1b��R6-̖W]�5-�ؙ9 f,ةr!�1@��ڇ���o/M��I�9VVM��㻝ɭw;�s�e�E8���psW\�׆��B;S�t��u�r���� g:�����Ow�}U_}�~U�6/ݾ�lW����tMI�@j쀣b(X7􆞥�o��o���y����Şǻ�t_'�^qpu/z-��C>},rY�
�ّ,��&uuC��U���|��o���o_A[\ȱN%���8�����ͷ����OV�G�`{1�|��9�]g$�{�5zf1�z�2^��8�`W���n
��l�Ŧ�>��"/�ٝ��7�:s7\�zO=�{Y�ȸ#�
5��[�->����&�ł��w�L�*���63EB�V�lXQ֯��,r~}�N�]x����t;�c���ћL�
�F�^8�3OiW96��/���zI�J����`p\�|Q�4���y�V6t|6(��0yZ��A}o�z��:��W>�A�c�lXW��V<��7e�96�^
W46;zf#��KE��7�Oz1�q%�/��:;�Ip�zآ�Z������7O�w�\\<B��~���l�r*��<U��"|:�ڤt�W
	��wfp�by
e��f7�g�UqX
�^ѹ!��=��5)Y��.� ���T�n-n�:ۛzt��oa��q�u�f�3NE�qXss*����6���`����̃��	7[�hpt��]pQ2��;9B�̼��-��dN����ﾠ���l�n�����=}�{�V$7T�����_���A34w��=*搷��ڝ�m�oć��|��m/T�W9Xx�$��~��� �k+�ϨO	�w�i���rr��<d\x$pjII�c��߾���SZxȯ��2�ٔL"�#u�R�Ŋʒ]�%V��O������i��s��(���Ev��C���2��gس܂�������C��p�]RţH(���MIƀ�>ϯ�%Z��<�K3,��E}����������h���)�χ-ԏ���oګY���o@�Q>Z�]��"��_o*-�S��p�4�Yr�s���l<!|e�8����<xg�z�����S���.gX��)�.o]�o���}���g�Ä�Mk+���R�\|��se�A][�U2�tMi�X���ۨaqQ��<G�c�xZ���nQg>�5e��[2����}�:=z��3A�X�-��q֢cs�Ե㧢z���y���bR�xu��HẨ�a��h���/�k�2��.u�Ǜo�z�Di���ԭ�yk��"�굻�}��du-4"kM`�+�;S�h"�yk�-����;�C�z��s^B����;9f.&�c�0��@��������8ZN�����_~�������Y͎��^��*���*��^t,c 61ъ,qX�;!�r槫��1�8�
�<sg.cs\���K��Z�-5�W],���M��2�J1X�r���E���3+�o�8R�{�~����:�P:�/$�:�����0�u"G��X��޶���a��uoƺѨ:t�9�C�ßl�d�C�#N|�$����0P�/:��=X�U�Û��+�S�o�u����O_�k��>�����Os�0�\&R2U F�@h%�w^�U�+wB�����n�hW.S'�)����g9h:
I��߲KƯ�%��&Y0�(�vY�w/�γ-nGǥ��g�q�XP�W��b{�b��;{�t6��Caa��<t?�P�g=�繵V8՛�����üd�H����/�V��p�Yx'�^s<d:8W�9��B�ʫ�:��K[ƶW�{�[GɆ�v��wORJ�JE�g�+�Mc��Ð�����$��y��=��_4�KƠ3 9Ή�VF�m�g��>��ʦE^�]��9~|߳���=N���*�'a�.��]�Ť���玱���۰��yE�^��a@��ǯ�#��-W!�:��ʚ�}�/-W�@�è��HLj54���X6"�gU��8a��^RJ��u�
��췸���tI��bD��޵�q�}����q��8Vo��~�Ih��\�U��h�2�'G(}c�V&��+��ǍV{i<��eW;=�\�@h�=��ە���L问�(��q�8"��L�b�����/��t��i\å\2Mٽ+��U�w����>ܮ��,lP�^:�i`��v�t�<�8x%�s�9�<�z�D���Yȕ��u,��.�>k����qe9�7�T���26k�r�ý˥��^W3 ��Y(�^
���O���e.X�� ������ }~\<Zٜ�v�$�5ێ��˾W��j�� Ϲe�X�Yj+��"���z��J��A�WH�{�G�o�:���9󤽡���Id��`�.��g~�+Zɕ�Yk����6I����8k�Λ#I���\�ky���w�j���R��)���=CZ��u�/t�ɔ�\�G����e_%�ͪ���ڧ�T�"�������䰳=��<rewz��[9�-8Q���չ��eR��&t��l�.� ���^�;×zaf^S��_;����Z���Դ���t��1�w�
�*䡊�깑u��4���^nj��w:�a�t*L�խ�v������Q�sdc��:vʚ�N
�9Y�n����8@���؂����K��7���b�Y_�D]��zƺ�VvԬ�/�3q=�����\ v��]�>�z�~�=�߃��;��/��E^�Q$��m��A�^���gܠ���򰝌�{�+'k�݈甒�!g-��, �夹�Z^�yw_ݶ'/���S��+ؼci�1�y���9��	yp����	K����-J���2�-r��yZ��\��X���>�e�������W*^	V�7􆞣�!����A��S���/X�ܖ&���{o���}� ���ʋ��-��+��
7�P�o�=K�>4Q�7��Ę液�>�^�o#�Kչ-0�u��~+��Y�]=� /�[G���ס�f��fZ҂��)u�����E�1�9��3SϪ��3�L�,�S63ۙ�j�i�C~����Y�3w�����gu�;���bwqx�!ٕR�x��l�-6��֙ynu��y����'�wlv}�v����}5��V|q�(��U���v#���r��6'v��j�G3��8�k�:Ҁn[19vgC����m<�gr����x�8�קb��/n��JEO��,�=��$#u} H���ټo���3�ǯ��;���8֞����KgD�v�]���M[b�b��I�T0ϫy�GקQ�ʝ5���V`짵�5�Ý����m,����m];����ZxqGܲu�-�pE�7p�g��-��}��2��<�L���#��pu���T1g�3,S�����x���`��xߖüD�[g&��a��sM���
T!+X��.i�:1M�d��M���hf�C��[�B�!d����������'�j0�.,��euQ	u6S ��M^(�7��ŋ=����$����.��O�%"��䈫Ͳ_ǋ�h&e��a�,O!�L��E�n�Pi�(j����ؖ����<�E�^�:մHt��5���X��^
�ط����9��n�^,�a�I+�w0��}S��z^g�|c�����38߄��B�΁k+��]]",uS�$<����ղ��W�l��2Y�6K����_�Umq��ȯ��P�~��a���D"���N1�`e�mN�����-��v8�nn8�JQf�VD�Wl��;�m�.���ʇɘ���R����F�?t$p�ix��3z�,70$�l�B�3=�@Ӿ�2���r��^MIp�˸^%�o�D���-��9w�c��U��M�=$���xq�a�⟸���f�f��;�ְ�v=F�Q�y��Z��9��\eZ�%q:��ț�2�=4U�$A�/Q,�Fg�nՋvt��|^����V����R��x�x=ӛ�f�C�CU��e;M���V�]/��ç5�N��b����\��}�����ٓJ�<�� �;���X�0�˕���v3a���K�&8'-�3����PRfƮ�o|�	�2��'pk�I�O�kM��^�x������{i��GzI>���<��};��je�׵��/L�⳧<��p	��j��=�f�pn���׆�SUc�%���׳�\�Xj��B�]�Gj'��̧s�|z'�&��Mi޵u�$7�Y�Vz?Vj[�N��1�=�[k����t7����Q`�C�9�'.jq���ؕ�(��%Ӽ!�	B+T��va��*�ʪ�+����$���!Y�F rL+�����~�D�;3e#�����:����C��T^I�amB�qx/�a��D��f��Ug�7���a[���S�#,Owy����a��,��*#M�&�֢��;]�acp���˿k�U_STS��(���l��oSŅǽ�^c�+�Bz�D"DP��Sc�����~�k^tm��5r��XbP����'�;�J��.H��:2KƯ�-�ϦY��Ϗ�r��`O�Z�F�k�dKZ��)�#��:��ˡ�@TW}���Z�&m4zaM�x�Mw����w�p;�!�s�"#�k�٪�pW[���ɝ�ͥ�u!���y��r2h�m�ݻ�4�ǵ��ڀ�\4X*u�m�����]�V��#�%/�L��R�v������u���08�=0+�W��af]��!�P�Fx�@�f1�p���#&p|-��El���g�OH�^��ǭ��WfF�e7;����-)�ٮU�C}�MKp���ƒ�Bc��}uo���+m|���7�u`�������
G��-*�������dVZ����%�d�OVL���*�%^��ĝ�jݧ��V���k�]����uۄ��h�:t�gS@N#� ��^N��������R3*�cr�ŘTS:8���Z&�<��ZD�F���G.��ٓ���J�h����r��є��#v�o��a��6n�p���l��<��i��T3(D����L�Tx�-E}����k�Զ.���y�������C����q��n�
�7H�6��p$j��ZvpT��E�>��v�@�Ō����J
��-��)�M񧫒��e�!>�;�w�����gO�%�'���VU��("	�t�R�]�:d�;�Xc�ޡ�Ac�N4����pfw�]RP����|��Z������sx
l�ϰ���#����2�|;��L�kH�!��Pa�^�R�x\w���KHZ�z��ݝԑZ�F\�-VgB����JMK���s[l�I��7������뤻tU���b
M^�}�@ ����n��D<�[��)(%qǻy����	@��\���֒��{:iWK���/�-v��b���oUP�!�>�[kRt����=�).R�Y�����\}���:�x�KO;VN�������:%�����۾�DB�K丘������׽.P귽u��8���.�,$��TQN�E�1�U������q�n��V2+�B�W���P2�h����hEe:H��s�9�YP���;�k=2ؐ�GO x)ΟY؄;�k����+���M4�V�W֦�`ŻS����Mp��K'�5Ե�սҊ��U�u��3G.��W9$Xs�h���]	[+��Ʋ�%K�wx���/�{�B}Z.J�׸Z��ڐ2�Ы*��4r��_7A��[׫ "ī�xI��>�ޔ*P��f�jv�ˡ��N�Ӭ�G|��9"f�����"ʐ�X�_t�inJ��Qa�5fYLI*枖���>6&K���to��Z1�f�]]�uNs��h�W{`�Yӭ�l�!�ЂZ�߉o��DD06sgN݊s�ί-N��8gD�Y,�+���uMt#;q���x��=펟n]n�O��}��C��I'�	�}W��D������ގ�a���������~�<�����{�cP�(UI*��P��"�Rʭ�6��eQ�"���E�,�XcZ�X(�ȡ+UmS32Vҥ��!��\k1"��3\E@���`�q�U������ ��T��m�8��kX)1*(aZ�bakU*%LI��Q�V*"�T�b��dk(�F�TU��ʤ�[��PF�S0�%kZ��*�TQf0+��EX�a[JIF&Y,H��*���S,���4J���J�%E�
Em�D�PE�c2�P*c3)i`��jJXh�˖E��Q��a*�Fڋ*J�Xւ�`����UJ�E*
[bҭ�eE"�Z6²#
��J�(*[Da,�`TR��U
ʀ��eJ��b*,R�TQk"���TUU@��b�L�ُoT�B4:	E+��w�r@&���=�5��Iq��.�:���$Ʈ��($�*�/��{������^��ݢO�:D�#K�Pz���6P:��b6%^j�P�Y%L\&{<����mL�Q����XL픎�\�P��d3��Ӑ�t����ʊ�����=/���Q�V����ѥ� �brϥ��=h��$t7K�E#����!��5�,#<��v�Ԩ���sc�w��P�5�탮Q#A�S��]��K;�O.˛I��_�1Z2�ݨ����=es�^0����-c\�U�1�o�=l���.�G6�j�Ѕt�W#���j���<o���M,V���	�dz��q�A�����86����W����_���A���-z��d�ƕ�B��قnWb�ۖ6(e/e����KI5�^.{
;%��*���@z���GI|V�XJ��K�pJ
���f݇S��t�v��(t�Y-��n�W/SXD��v�ӟK�Yࡲ�JJ�����K�"�����<�o/�g9n�����\���/Jz�أ>,V
\_ԍ�ґX=)���],r u٪�ǘOg����,:���z�����i*�S۱K�3W�R��gV�v�F^���>tE@-e���f��/��Ổ�tф��[<����fVm	QL�EH�D�ȧKj@h�j�Ǻ�Z�'\ƽ��������T�vHxz�"�Z��D��G;�u�:AZԵ��\��4!�GRu��ۆUZ�Z@�����î\��E1-��};��3���W2��1[�#[[�`�~4�Fs��=�t��2«��;��]H7\&�>�x�e���7�Y�+�ՒS6���X����gp��8T�2Y�h{�Dl�a����M��bÜw��>�t�J�
��ڋ��{ބ����&.��v�=ΔJꙍe������}�%T>j����ޜo*y��n؞9˸�S7�9��,��*b�0PvZJ�:E����T;�v�<�o@���ћ/��?kGؙ�֠���Wl��w�*s	o-$+Y���u�[-F����7�u��YkW�>7��n�EE/��h�|�|�>��t��������W���KE����e�����/g
ڢ�+����jOW�0�tHi�Y�珎ǫr�	�[{��{�P1���!�x���>\\%�D�z�ϟK�k�·�"S�{ԻW\����I�EK�dY�N:���3OV�Wg���-����WW{h,iʺz����yf�Pk w�:]�-����oX�����n� �k5�M�[n�x�p!4�Z������Q���,�K1���-\���r��}��z��aw<}�Z�.;{Le*a��(.J+��ʸ�:��x{+m����P�^6d�7哰[~�{;*�);}	���wNM����p��8H��wl
u�d�p馎ߢ����Lc���q�f3��/�ʗd{:\e��w-��)��F�T>r�@�j^���O�Ѱ��;��@���}K�Жt{���3���<]����ɟ+�am���)Ѡ��=c�gN��j��,��0_��%��T1z�1:�����,;�<�y�%�ޖ.��(w�k:��y'J�ҩ�y�*B�(#�4����fɴ�jW4=u艥@ǋ��+w�+ᣜf#���5��[I�`�2,������
�u�Vq���(��bԯz������ΞUZ��(d��"ĳCmݠhoR,Y\\Hf��ި���dyk�..d��{�J����ڀ�w�8O\�ؼ1�a�C�v�����X��^P�`w�t���#������_���"���`E�:��a��I���=s p�� ���\��ȯ#��Ńh��')!�z�W��]��͓|U�����c��x�F�����3�F�+���K܊�G�ٔvPX�XKZl�jZ5!֍�]^��k�W�𚝕�i���c>͐��&0:�U��3��d��mw.�٥��ҙ!FivlB�"Cw��w*������������]�w�lv�Iű&��,7�+2����dW��.�=d�W���%�J[���L~=������0,�_-�؆�srE�IJ,ϻ�o�+"�+�!�xK���g�7�v]�ɯ�za���tlp�e�G��aH��jS�ύ��o_E����B�P�鈌P��uϟ��^�09J.Xæ]T7�Z6}>�L/��r>��V��eY\j���L����}��o�Dϳx P{a�"Ƽ����ۅ�X�pT=�_�ʥ�Lp��k<�u΢���y_{ܖw���	�h�>3����w	"�ޒ��W�=�w�xL��aTηꡗ�Mz<�g��T�r��6�)�ub<+�f�0x�zf⳧�x�6X�J�+[P����Gy�x�|C��%�4�"q�r�3�J��W�mgq.���b���=Y��p��Yz�&����^��U��`�lz�cbX�JKÉu�����tb�>�C����|*�ڤǴ�ن%�8�� �#;��P��&m���$�yo�>�� �~��W����q҂j8Guaϣ��l�Ы�I+�����W�2����3Fެ���yB�,&M��ջ�')�:wԩci�=x �y��Xl�����`dN�T%4���m�ӾW�0�T�ڗ��d�����,`%�L��w~����8��k���k�.�pkyo��9Cm�T�	y�0�vU"�r�6��8��1M^�@�UZE����R.	��3��9�;z�L48�4�\��֥����fz��;��{�v��\�o�ׅ�S5(7��3�	�o��w��ڹ�����:`G�����_�ز�1UZ����_�I����i칾��h:
I��a����}�f�/g��3]/�x��h��O��a�kґ&�fq=^�l<��!������st9��zuךf߫jt�-�n�'�.9��P��H�)4�UB:�����NB�5�k3�ŕ��g�)�����Y��T<g�����	����9��$�t�_�
��R�du�Zfe��78nV/
I����Ն9-%e�\����$h69O+�<�4Y���c;�yg��^8%��.P�6Vo��SO�Z*��%_�3&��5�U��h?Z�Z,��y{e1��R�fN"Q^ZxV���L�#�P��/�wFǜx�}�`^"��+�����U��|��q���M��:�Z.��Q�/^ɖ�fe<�M_n���k��R���C�c��WO)!8]��v���[���i��ʁB�es�X+g]�2��㤮���$s2�r�]�P���0Je�[l�pjvP������UU5kq?�Ǜ]��k���LP�Ͻy��bܮ��卋>�ZӁ춑u���
:��vO��.��Xl���,�RW�"\0�<�'`�hA�Ht;YZu�(E��e5ѷ�ldu�jɮ�|�=�7>XD40�k�V�\�Q���^�&za߹��tc�}-��In�>$��i�N^�����^u����VF�M#�M�]�u�޻�\�v����R@���j}�*D�zY"�s�@�~�,t�KP�Vx?�v��#ڵN�ԩ�^�Vuk(Z:4�U{K���G>�Z}��Ͱ�������oYʤhׯ=��1�I{|����m&GGE����WLz�@��T�|myN5�|rE���)oβ�{�S{���\�h��(���(�����]K��h�5���/��Z�}y�(�����VK黓�u�x��+�52� s�(��3�
_nq��/]ʃ��w4��3G�y���g/,�te^�r�!g.Tł`��夫�"Һu����$m�J�ױߵ��2�7�M���Pzrk�r��;�5�5�����c����y��U�y��;Ym���i��|	pqOW#��@�/����q���jfڜì�F�S=؛�w˶�Ɔ,o�3p��1̛�b�B�p�*�W2��q�l�e6��m�����!W��ݢ�}s�U�="�g�%/�ʄ_�	a夅�U�6���������"=ה�߼�VjϚo+7e����U�NHi�8��Q㩃.�7���j��̨��Y�X�m�,���.�!���޾����<�B��!��r���ϫW����X�I{�B�:�6ף\/���y�P�ν��'�g@�8�MpSy�4��)�����~P�ζt��C��W�Vr�E���ۙ�޻2�(��?g��n���EOc�\�̺�r�����ax;�x�Y[��҇�n�{%�-�GWy~-�z�S�"kx�#���vX�U��Gq�3�c帴ӺQaiTH���־�O�ǎ�4�!��~7�1Zx�ˋ�gۖ�N]���!#��O��3�Yh�u�i�z��?o��z��ց��i�E�0���:�L�:�vQap6ϒ"Ǚ�2��Or[�������������E#y�
�[�%yъ`�L!ͧj���^�\������t�t3S�"8�$��\���w\3�����}i.�z�+�K �Ȅ��u��u˘��3�]�m<i�׺�v�;B@WPn�c�]�:\9��i����_;�����h��i��v�9��d�3U�����jk/L9��ް���VT����Z�x�@���U�����trχ��ܟe��r���.n]�y4O�/�g�����5�H�eqp�Txy����t����e5����,."<�e�Hv��{μ��uyB5�C���45rP��e��m�Z}��g7Ã����Z2�@��O��5�T�=�;��9Xx�d��o�z�ٰGr��wjI�z�n���}�g�V�3�<��g�w���lI��Ia�+0v5Q�"EZ���ƽ�%��[��٧`�d��4I딙V)lR�>�mȼ$��gӦo�+"�]��]m*4̱E�a���������g���0�)��<\VԾ�ϰ���^݈j��ph���/G>+W�Pt̀�t��u��e�8�yL�$f�Y˔��K����W���0����G�>�3�@��p2,k�h�5Xܨl<��g�T=�Zt1o�a_;��*��ce�G�����=0��w���2��:��bL��x5���Ͱ�m"�]����p�֍�.�9o@i����&��2�����L�jC�RnO>ydb��M�=��{��ʬwۻ��ȱ�%B�u�^e��3�^擐�a�w�cCz��Y4��P^��H9���R�*����#S޳�����a��>���\i��d���^�ܷ���/}~���8'�/c�g��R/ee�4�c��}�7�G�1�hLl��^ue�p��|�b���0S��O�q=Vr�ތ�}��C_�+5�����5�����S~P�{�A�gQj,qk��=ut��JI���v�V��;��#;���T��va�r��'�b�a61�$řz<=��;��9�N����T��L�Bqu�s�X���9 u���/)W���n�T���5��م#�;y���:�g�,�B9�g=(sXpl��aQ4������`�:i���5Y�\�g�w1Uz�)����<���>�{�u���mxఄt�[=K2��^Kq�`��C�Iֻ�(tXx��?;�����KA�RNl\�4��̬'���^�=������x��&�v&�"I@�=��k}�z��a�����A�89�]�<�x��7#�g��g�S�޷p�ɂ��0�=ix
��/�� ���^�M\●9���:�R4��~��{s��f�ش���֯5^̧��)���,�Y��{Ov�c��!����.Q�Ƹ%�O.��m����j��%-��+%���_���ݫŏ#�7*�r�U��ۘ(�vt�J�yMCl��v��Ê1���������f�x�mh�,NY=PؙI*�H�L;B�����0��Z_w^t��|�>�*���r� ��ėlQ#A�����a�R,��-)�77յ,�v�I���U؃PrV�~n��v,�,�Y���q&P凕b.uc�QV.��tc��r׎�N�?5�B��=��<c �eDr�� �<GX^�MӮA૪��wY��,_}�h�ط��+�%%��'�O�%p�]i�7,lY:bo6�3���Uc�0��	�wc���U��d��Dx����Y�L�W�J�TG�q9���\'�_���w�݌�k��Y����ڜ�V�P�i��g˖���{}g�'*V��Z���[����L����WE�e����B���eҬ�g`�g�x��gQ�Ѥ�5%�
�ϟ���:o�g;�����@U�B�2[k�S�y~�{���E�,����G--��֌OXֆI��{�
��i߭)�<�C}�.�l�W��gb
mZ/��cQ��X��7x�!�b/7��Gm�܇Q3j���A�L.���(��k���}�zk�1�}�̆f�`r�k+{m;2��$D*�Q%@x6���\���h�i[i��C�N	�s3�i���;s+[���j��eb��/zmhJzn��GtU��U�kW�%]a.�.(�p��]�LXW[���\\�
7{�o{�T�fLSc�Z��m�C�^
Ԭ�4�5fu�idX�NU��i�٥(���+=��ОoMq�9���H��-�ͽtir��\#eǘ�u�;k4�鮛�:�5�ާ���e�9*�ŋ�������2�.[��Z�̔Xy�
�.˨��Nu^c-�.��T�J[�Yf`�]ˬ.�.�8a����%@�wH�Y�o��)�v�2�ÛNٓ^<�ʡ��iuft���<�3�o,y��S�
��{��$��0^�esy]h���ɹ���v;�y���vQ�
>RN�����&��7'�rW��\��p��ep5��)�`n�mb�#�P�B.5�z'��q�r�'�9��؋��, ��u�)��vX����tΫ%'�� ޥ,>�nvbQ�]`�j�C b��q=��u��Uc@o���j=մdA:��g�fL�)Y����=��^������K��/U��3>���'-I3m>�}94���L���f3�|�P��o��Ntz���, �\h�:��OhL�0كL��@f^�M���OBMޢ^�.U�vx�g`��`�{J���k�->׻4�����⥍H�m���h�4k�#/kn�n%��q�i�+�Y�
��$:��Y�-u��3�#�R5N��r�Ծ��
w8.6�<ͮa'��U^�V��P\PUL6�l V9:����r�:��d�C�.L.;n>q̺K�)����X��)mr����������
�@�z]C���vn�S����l��ږR�u:�ۨ�pv�n�Y���3�9
��1}v���`_pm�'����̺
,י����n�p��.��Sy��|޲��lԱ�`����g0p}���4�
�Wh)��������̏�Epє�Yx����OE����L]۽Z2��gqN�՗�@S�N����f1E,رRx2r����Y�5��:m���Nr�1R���������n_J�2e���ju-�r���,P	fd�n�,QZ��j��F�fi����Xx;�5��������j�>:5��2���Q(r�E?�3E���YO���Hư��4/�c}y�ʚ�W5��fU��o���]f���d�kdz���Y7���o@�P�er��ű�.�n5�h��<�>
s+��Ѧ�t�|�N�
�4{�'OS`���R���.�Wl���U������$���o�dWj�Rn�m㙯Gr�����q�1Q���>�q�(�x��X((�Z,YYV�+
Z��E
��,������R��J�)*aRX6�e`�()YD
���`[J�ڢ�
2�5�,�mkA,�V
��TR�IY��
±���-�Pb
��b���BT*�F�*((6�Kj�6�J�Tb�R���X�TU���F+ �RVb(�j�j�FR,"�E�b+
�K
��ʈ�UE��dX,��YX
�%�Kh,�dD)QUh���P�V1U������m��(�(�HաY*V�RօE
�EZ6�J�k*,++J��QB�U-���m*�j�-�m"ȱb5����$kJֈE���B�+*J����D��,hV�*T�*AjVR�Q<�����m�HJu�ʇ�c#0�<��	яz���!�-ǲ���HƳ��Q��������4�kmho(��
��e�tr����1���G	�'�?�$F�{3`���XY��ّ!=�ŗ�h$g�������s�U�x�t�\�G��4M}ΔD	i�ն�uK�\�<N�d=wUyhyu����[B|�<�'�w�\�ر�3o)_s�I�֊�=zm(���R�t��ޮف�S�oFE*��CPެT�,�R��0Pv�ѯ��-$�.�Zpe����r���r��c�u�3�`�������:��OƲ��q�Ĝܞzz�2�#��v63��Ȗiʫ�zk��܇E+1�^P��EV�2���;kcW�A0��vy�CvI���Q���Y��]e�<}�D4c��渋}�W琣b(X1����S�'I�h���x}ey��q��XC5�����\/���/����A���nz��V |�^��ƣ�\��#y��՟uçojd_������\/�\\����m�/X�G[K�hm�wEw�Ӏ�+H��=�=���6�.>�e�/��\9XH� �ڵg�6Y�͒��:Hέ"�K�<��Z3.�-}1i*�ئ8�'Sv�C4����J�mR��cm��hc����L������k[���d���n�v�����L���d}��6Ԕ�.k����;P:+{i���Ь3���n����Y7����E���^F{/L���ı%���(15�|�b�_;��14�.��>�|`8-�M��y����|��2���ĳrٙNf��BN��W��M��5�!�	4WrSԖ����o��i��`V��|ßy��-������rǹc���τ��V������D���ޏ�����!�T���W�°��J���3�ɇ��=��<�}۴�Ū�9@�8��P��3�q:�G�q�`��,
۲��)��߷�0	�o�(����v�Hz���>�7�`��0H,2.Y���wh��ԋ��q Y�=�U��k��d�-[0'Cq]��֗�{�x��f�tC�Xh��;�j䡆�s���8U���֫f�
gm��S=.�(��xg�9Xx�d��o�O]�@���a��׋}�1ǭWp �٬J�-k����޸�EᲓC���WccU��"�E��y-�F���ƽ;u����؀� �W��-�.�3�ۑxII���6$��=Ý�seI�Ijad�[�ǎ�zr��V����\��7Q��]ՠG%�کw�SܚO'��+�՝���Z�>9
:B`�0*�V/������o�rG����v�O帎ub�VŸzn7�K���\2���U8R�d�x�7�2����iг��&��hN�=`w%9򵺯�8j�f�Ta��h��
\}.�\�|oU��o\8��s���P��M�O{��_c���!s�`씚���s.���^S:��ȳ�r�;&oY�NҗVM����Wa��P�L��M�5�aIA��JƵ/r��nT6�X�Sc9nYt�g��9{��U���Y�>�u�D��rɟy�$�e�+�n���ҷ�D�]竵��t/l��)=Y�V��c�`��L�n=�e�qYӟ=���b��e6'W�c=���K�Ȏ��D0L����\�-W
WIm��b�7-���b�^�W1����.���३g����t,�熡��j�Ϫ���U	4/`�g
�Z���W	��u'�fM���Fڕ���t�w�r����\�L:U���JK�Z=��2��������d��u�L���V:1_�NB`.�5q�C��uPK�Ckjk���s������GK^i�{vj
��Gb	���=;��k��ܳCoਏ�>Np����y��c���0�ܚ�G� Y���J	�By�lc\�����_��9�H=~�R�r�����W�k'�rb�&}�5��R�W&S�]fg]��^��1T|�.�{�>���;��۵��G�k5�r�T+Vd�k\����P�3�Ԡ�g�ż�'.q��:��B\��e�����<�Pld���oS�{μ�2�*�}�������p�5�d�@��8Ky4ٗ������f ����wN����-<b[y�j��7Y0ؘh��'�=���^�>�2��4s��k��z��t�u��a��iY�ռ�{��*#])4��U��@�>Ľg���|��3��}���/ou'Y�K7��0?}�Ӂ�6�c�')�)%_t�_�
��T�%=��>���M՞�^ջԚ���\P��7�%w���}e�Ѻ�������fvE�ܾ����[C7>�o�(x�wKEX�0�&cDܔ�<a���J�^Չzk�[HtF�#|�TB��y[��dy�~���z��E����(�ղ�#/��E��p�K5�-�zҼ2U%��蟍?����-����NV�nUby�P�w���l���Ħ����(i�_j�B�̥K�ZL�.�P����'x��	�rnJW밙纕�-���2��������wcZ{��m��	�ݩ8,ٔoKt�,��w^Ɏ�k�ˁ���3;s�މ�j����κ!,)�{���o���u��ջ����"M�E�f���[K����v�;��/#.��ŧyk8�O��wk��G�wcb�s0o��Y��p���6��Y�.WV�"�N��+�lz]7Vd8v�#q�VN��Q��!&ǥ30S��x-��A�6*��WJ/��ʞj�y�7����|�y\��o(@h�N$|&=/�v	�]G����V�-C�m��o���y�= >Ե↟�-��u�
:12Ұ�1�7Ƣ��G���_k�=7���v�t~U�9�&R=}v���'Hx������WLg>Յ��H�Mv������̗=�lf�:�U>���ܖ��2��K4Mt�6P��CO_ޭ�;\ɨ���7!z/,��t9]������<�/OT#/���f��@�:Q+������셳|��u�y62ٮ]Y��|"R����+�U����B�\���A��y�ZMfM�:��Ye��ΞM=7u^>��+Τv,i���yJ�!K�Y�u���.P�/�׹�����5�׹��\������.᯳k5y��۴L�P��*���x.�: 5x!t�ļY�N̳a�s�8e]��^2[Va��b�}ޣմ+^4SR���%h�v�x���˙P�̒�-+}��ؒcy���vg��#Y��^�dN��[�4qwC�,!��[��$�*�oYu�3ʽ��k�H�g6�c3M�ث(��X1}ԯV�6�y坹��M���Q�a4%�O�}��"�o"ָ�c�`J���Q3)�	���W��{]��Ub8��u3��,!Kf��hzב�0�\\%�?��E{�rmu��oZ�.�ss{z��PQ��p�ά�M���#5_�+Ҋ�~3닇��Mc����v�r9�]9Uzm�'@��d��2���;�V��0���E�%b�uw�V��ո�]vm[v�x�.4��t5�o��H���2�Ms-��J&:C����پ���Hgc����n] �se�uP�pyqq,���Nf��y;���_�'z��}d���:2=g`��YK���e�2�/+EDR��\1f�f_��r�֫�q�f�͉$�}\��|�y���-�WH���P�Te�J����w�I�ъr�M�g;*�]{y��fҸ�����(Nɘ4�����x�@�����y���㭼�̑T���:�xT�Ú��|5�/:����9fH,2.Y���ѭ�E�+����w�#$&u�/�<�4T�Լ9^j���h�AA�,qI�����A!��X�Y4�*�>,��v7�w�$&ϩ�A�z�D�A�V�9Lu�	3w��H�P;����o��z���M������q��rm.#\���|���w�pGqæ|����T���J�O��À)A��[�AŦf՛�e��XЖ�$?;�������e֕�/[����=����=]��<P�kԬ����r���I���'����Қ]X2��s�{q�fЩ�*(�м�..�T�w�%zR�/[����9��G�+��~�]�=KoV�`�l�e<h��RҬR��ﶤ]%&��/�"^w�f;z��s5sƷ��9��d�����2�À?F��j�q��˔��a��o:w�.�3�B����ݯm������%2�38�����:o�p�Լ�u3U�,���Rŷ��[6R��������7]�z�
��m��Z��~^,��t�{������;ާ����7�E�3�VBy{��׍.:e��a>jFɋ��Sf�6i��w�nk���:K��2|��M�ь�[�������	�gK��b^�).;
�K*�q�o&D<&bc�/םa��U����<}>��x;k��
�[�Xg�����º�,-�OK���?�5��x��6��C�s�L����,>�� �ľ킣�WV9؆��D�!v�_sy^46�:b�Mf��=C�o�x�Mo%y�%j���D�5�:�O@�ս���W0��,<���h����s���ņ9MS]B<��6���-/R��T$��X�0m���~�zW!�����%���
dlG��ñs,
�C۱�; �H^;0����m$�̯k9Y�q��2H�*�9�Wj���I7������3���u�|�	�E-#I���L�#�V�Ȭ�~^��5W��+N�s0�}N�H���&�2����r!�Yc`�7,��8]�e���~���L���i�D�y��U�gS�GE9sW���G�K{o��3��ŋ�O���^�W�]9�v�M���F�[�`(t�Xx���yr�c��#��oNu�,�.��:x��p�Ʈ�3|�&C�$�F��P�V9Hs#*S��s�˛�`�o;�A*�P~P�X�L]�C,�g���g���h�$WZ�<�+����縶i�}�t����"�v�R^�F֌r��OT72�U�JE�`�^����*��S�v��"�z� z׵O�i�8;����K�(���S��]�1��U�������Z�o�/&T��oš�/r�����c˦E@�.����o��%I�dx��,d�γ��*��iuL��,��f��7	�3Yо�h���wݷ�Q��}Ͷ�*�Mu��\�a$���	utضt�_N�UmfjWz�Z��zwAv�ޘ-_���וK��qK�V3�g۾d��J��h�S$���y���H.��l͞8�t��7=g�L�ʈ\C����ZS�0/��G�e;���U�k�ϱᣘ8^/J�j8�;5��Q���`��U�*�ſ�J��Ip�+ƞ�u��Ƙ�q�I��Y�qM���*��Λ���>oz�u���|���������MS:�E�]��n����[U`Ϥ�"vYNf�fu3�S6���d3X�]_�a�Iᒛ�{lY�.\��g�R^�7�W4py؄���f
r�O/��GVѽ��#
!��e�>�ǰs����R�P�A��|)Ďy��,���G;�.��gGAZ�ݡy�/��/`�q��\񘮖!kƇm)t�d��=(����P�ʘ���QF�q]{=����L>a/^���Դ�l�G���$�#yX�0V}]1�Յ���xv���mi��2���p���zq��i�WIL�-7,�5ΔF��iN��Ǣ�/mח?�ѽ�z�É��w�w�{́c���X0��^p[�*���{&�}Q�_/bB��%�<Ŵ7 �4�Z�`�u�:֖�^��ӛ�y��<sgJ�K�$)��u:�o�3���K՛��4��m�h5C3O
Kr9j��E���q�&���qy��g�[q�LP�����c�f�yH�D�f4b�jO{=޿ߨ?ߢ���ՠ������S��k����jՎT�,�ʘ�L���
�0Q��Qo��b:�=���E�=��̗��<�gR;���yp����(Q�o�*��|���W�t;W~m��3��L����j�33�sU���E�`ݢe�P��*���\6�}��3^>��-��=����[TD7�a4��b�+f{´�ex:��td������]y���Ƈ�<<�N+�`3�٧�q�,!J�f����xL1�/�x��}e��ǝ�u
���+6��$r�%�బ=�<�՟uçoj8Fj�6ψε�;:��c�+D�{���&ǠÔq�ޗ;�f��H�=�f4�<~���L���a�\f��p>U��v-5���O�<�`�Fd�C��kq߼/n��]���(g�\��qi��&Uܩ�}�'5΢P�-��z�;���Cx��<����fe9�cC�=*n�n�l��3%�E���=r��^絝E`X!ϲ�0���xY�إl��G�Z�5Ά�U�����v�Y�7���$��ի�0�;\��L���o0�*�@�R�i-��]��B��G*LXJ�	���y�i�zt�{�/�7]�ZB�oA�W����ҳz�u] zQ�7t���j���E��ne�Ҷl�`E��WZ~̧��'�\`�ZgdlA|G([��7����^gvtA������cMa��Q����g�H�2�:�r%w26;n`3���y]�4bGj�-�y:��c}\H4�u�ieX��fr :i��Gk��U��.��ՙ����F�����QD�6��*4Tn���<�R<��Pl�U�$w�g�\����f����G%��1�+˻!U�<��ɜ܌t���&�$�/o.'��r��V� ��+0�x�"������v�P�[�(��yx����ә^wY��1`�Y��ӗW�9r�7N�u(󹈎����u����ͦK�1�E�a���z^��ΩG�ʇM�x��J��&D:�z1����K�Z�W�ggM[�^7n��[�^�@[�y@�<zd�b��K�e6 l����Yų��jK�:&)g����X6������L*�귫��[w!��f�]\(7ۣ��˄�B=�0��u5�`(����q���X��xފ��Ώ�8�J��C&��X�T	]vk�=��
�TF�rv�Tk�h=\�椥��GP�p4q�=�֔����[P�]�α*|>�V���;�>Sp�!�(/�z9���̭᭣�3�[�'p�D�����R�7PC��y)�r�h���l+�3�Z1���\1]a����z��K\�\$����CO��1�6-9)X�#�z(lά��jb,��H|�5�\sJ�J��7�bЛ�]�����4��.����sћYկ��H�5�.�U��+����R���]r��8�7��4�!�ܩ�ˮY�5Ԫ�*�@�Ӡh������V&�;���ߝ��[�X�td]�%MX{���p�\�	���&u2��54�b6�h3\��mk��#O���lh�i�b�b�1y�Cz�X���a4N�E^����Xܪ�Ԙ� �s�e�wDr�N�=��w�|k�'<���	bs�;�����hSr�f�������zl�^R��l[�A�8�P�ZVD��U����D�]b#-͵��'u��y@+s ip�G�x�V���P:��{���\P�e+��r벟f$u�Tz@^K�E�@s��iU��5'�+W��r��4q�LR��̤��^�@b�g6�YOn���Xl�T�s0�ˮ\���9rt��b\��9��fN�Gf;}۽��2�<�٥��*+��wM��MDS�w֮�#�fnB��3�ӷ�����m qW�|E�P���������W�ᒌ{F�c��͢�z][�1ltBd�0I����)k못���ث�U�Y�KF�Ҵ-��Z��dUVA�mh����Z�*V(*�e-��J�Ң�@P*��5�X[ek��T�ЋmՕ[[��+
�V6�j(��+R(T
�«�,U��ch��D��l�J��dYi�`)m�T��"���J�XJ������F���d�V6��Q���D����eT��KJP����k�AT������eFҪ�b����R�T*�`1�
V
IU��Um-,EE[TDE�V�**���IZ%E���ŊTJҥ-�(�b��#!A-lF�Z֥�l+mQT��ZKkm�J����5���h2�
�J���Ŋ(ơm�*
²��QH��(�?�%��yv�>��$zm��@\jio�X�'T���2�.���&����[
��9�+N::Z�QV�N������^��k����?{Y��5+�X����+���Bֈ�ϼ�C�f*������^��V��ޕ{]Z�����^�^=�-���G�ҡ�.c( -�@��i��5����}௲zs��QՏ��`ͨp'[�y�&��l<5��[I��E����7��h�*g6�7�U�d)�;�+�M^�D�y��afr���hm��w�,��Q���4����V]�v;������'��{�[��5����?d�G��rF�쓣���KK�u2�3/�����B<өX{����}�fq�нb�uJ�k��o}�ȠC�"{�rV)t[뾭CZ���rΐ�w!9���m�ћ��h��v���~���LA߯�6�}2�e�d����Rqu��f��M���G�[��4�Ϡ�ɹ���t�#���j������>�!ۙvaxR> p�����R�.
+�m��2����s���T��>������($��9%&�c�t�˸q����:��V�qq#�(z�M*�pn�^�G��vݧsO�uehŘ_ͮޱ}����N^����h�R
+;o*�.��m(�Wn��o��uZ~�b�z쩣H�<�FS��M�wc`�[���}Vp�>��yM��sl�6��f���W�r��I���j�������n�����D��t�p�
��ϴ�(�R���ge��돔�Y��~��h�E;�+<G\�i�hK�/�s	W�p�$�~)H<�ؼ�z���l1�&��:�ͣ���K�f}R���<vԋ�}׆v^��'�4����ӗ��r*X��ԓ�,9X�dC�`(v�W�%/:����R���qؠ��KԸ��ͪ����������8+x���g?
�qر:��^�D��D�0���Bq*�â�G�{`k�>�����+�S�������q���h�:L?�Q�l.+ʞ�$�xB�X7������`z��p�@z�zQ��N.��}��b5���P:��jVE���E��w�1�%֠�Vw �P̾���S�9��Byg�is�.���S��T�Y �W\��9�bN�ۦ1�:*# ���������o���}���J�4�ż}O;�]H���ڛ�$�J�����C-;H�@��0XK��(P�`V�˧S��P�^�J4v$%qT�T��5$��I:ΏJpY�@]]˃*�|ue�]f����6�vD:�"��@Ya�����k��`�x՚V�h�\�=��=�{.���9Y��9J���2j���+j�tR-�J&�ş��F�� �M�QѮ�.����|z�jO�㜆��{3��+�Kg2e��@�[Ȁ�+Gk�Ү�yzts-�giQ:�Ff�j�zƹ���A�*��1v{&C�XP�i�4�*�K2Sߜ�!��Dْ�a\�oN��r����d��5C�~r���9g�¼ވ��z.�Ϭo	�٧ycD_
��*���6{�<ݖ��JIqqBĪ`��Q#���O+���҄�{q�ul��{��<6�����K��qK��꘳�Z+\�V��h��켽�;յ�;4��d]�j�*�C)���;�kE��n)R�y�^D,g��5���S�:��_1�m�xp'pg���ⶨ`��!<lv�¢��7l[�֕�.�O�^z�3q�{}}������*�'���T뜽'�b��!Ӭ���l�f��d��a7���o�[�g �y��X'��wzܮ"�.�`�	P��y�ӓ[,WP�k�˶�y>CK����k͗jW�c.a63�8�;fsn���9x r��{��X�/T�+��ɢ�V�Z*{ �g P�ٺkz.N�vN�(�8hl��5o��U����t�����$H
׭�u`�ֵ�w�\	y;w�}x�q��4��w����z}zά(s뱴�t�i��k�|xӷ)�ŊwQd�OmX�x�)�[�܉.���Τ���WY�`Z7>�|U�_
q#�b�K=.\��u�$s;h�ެY������g���i�+-r�І��M6z� (�e��b���;���H6�Jv��NZ��q/���r�L�zU#��i�	<C$�j�.�-�䤼늙��8�7�·||}�(<��gʝ��y2��r��(�����{��f��Mv���]�75f(��%�v� �i�/�T���K��k£�?J�g@�?��AoR�ۚ�Ǖ�u+UV����֥Ȯ�lL�2�����Z���8N,�qKB�r�)af<u�O�aS���o���h�8����{Gm����z,B��yp�Ev�D%-z����oU�u9O=���l��W%�u�9�7�0�5�+y�}���O����+f��h�C�ë{<�曯Ub&NE�)�hJ�TD�E�+�=N֩O��Û��<;��=M��˶<qǫ��3{��j��4�.P�B�E������|����LG:�5��f�W���2�9�i�H{�nV{���+����5+�����5�Ӗ��]�]n����\-��vo;`�����=��J�{��T.d�r�����g���<M��[�M(l��l���&:ɺ�mN��b���
]�P��M�&����Y}ݒ��Sk�����8c8��{8�2{j��+�z
ǩ��N�w(*	�������vD����}��m֣3���{s8���PG\E�pX��m'6�%����إT�ݢwM'���˃�2ɦ>�K�����p>"U\x=�/c�0IvF��P��������6�1O5t���VϾf����H��W"�p�,.$���g��B�vi�暐��3�A\}[�z���цޚ������ե�/��0��QWs��\�o�d�Y�8@�ƛ�W[�E���y�x:�|6(���8���}����gS����=�<k6�q=�z����i6��S�	��s�N���1Bt�g�����M+��Ho�ٞ�u�K������:�/�X9��Q/;m��W�(qY����k��Ϲ�|��]<^An�a�`U�󪋽�^�s"�_Gz*C��{�u�#[����k�\����]�\�%��-I�.�^}B��;�Ҟ��N���X�=����ڨ�<��د�R7����;�atqe*��Y'Mu�	����QXAY4�=�*u('z݅�ݫ-p��w��	�|���4��["y�����Z�`�����=��S<+W��=D�_b��.��H>�]��\�	�n�%<B�#ghxOU���#9՛'�m筛�>���@�/�f�V)s]��3�޸�8=)r5����)gP��$��r�.EO�9r��tK:�B�qW�'^]�w�jC�*yCy��ܴA�k�Q�,���M�Y~]�RGG}(C�˳�dv+��˭�~"Fr�~�o������0�Vޤվ�%bJ�+L�Ig��u��_O%+Ý�g���4�/S�y�/���	��g&m��f��m)\7b$��*D8T�qd晅g��%g��4q%�3ox[Y� ��=�{ό��)1��^��LO���gz ]��/�2W(9����f�Q�l���m6��ڱJtb��;jE��f;/L6�#�\u�T�����z��Y����&������,��5e��j!�y�`-	p�ٺ;,yF�Ğ^�謿V�cU��|��S����g)C�t�>�^�O��}>��0�]H�iĞ��Ö�	�P�o%��P�ә���]���C��Њ�)Kr�=��c�Eo���[Q�XbVS��l=s�{�^����߼�c���ЀȣU9W�t+����RʲZ��SO�W 7e]}pm>��Rhv����J�/^�����>ܓ����7�*�v�֍`�tΆ�3.�o.o�m�}���)$���d����XS��5����3��[�N0�&�&B�����&|]w��}[^�oxWf�d��솖5mz_������3L����"�t{����H����2	��g=�9�6y�>�Vy�>�{5���Ώʸ.j|���
��LI��lQ��S�E�r�2��-��}N�Y��Ԧ��犫^_��s<p��KH��v���`�\�Aj�Rg����H���n\����zG]=���,q��}�\�d�s�&C�"O�_{�(8�x�����_����y�٬%�g�xNrװ�b�\��p�邡������Oq��}x�m�����~�*���o��3��Mf.,�Y����WcN(�юX��W�#�}�牓 ��H�g]e��6{�<ݖ��t�����]�'��]�,a:����;zys�s����t��I���וK���'�\3�ܦ.�H����Wf��̗��U�5	<Y�<�;ּ�έ�. ��z��F���^ZO�����*�u����^�c�X��ݝ"��h�p��̈�p_zWf��5yuhP��ה�y/G�Zٓh\x��٤�@��ȭ*��U�m����]�>�pj&�j�ך���8������:뇵��:Yy�t�ۢ�����G^/R�:�����2�żuI^O	�<hzP]��k�ם�6�����㥽X0τ��L{���)�9zOL�ջ�X�ʿ��z�نeV���T���z�WH^F�x�J}�Zof0}�\DTI˱�*��;��_��D3�9���vo^�r�����@��.X\�����%U����k��:�����/D�*Xv��ҝ3�;�T�1���֫ �"�X��O>�|V ���G�H�z\"�Nv	��j菣ͺx��ޤ�7�T�]g�� �k&T=���!kM~䟀�Cf^���K�(g��b��m�27��}���bDς�m�tږ��h���\C���k�5���V0��r���b�� ����N���郐�wVK���v�pE��u��g���@��5��ֆ0ԕD;��E�i�/{B��ˆ�k£�OҶ�.��A)��۱�n۩�L����PPL���b`L���.�ּ%��ƜY��d��Q�r�;]���.hu)7Ee��u��5.���3NWu�g`(O.��+C]�X5�"���K\n�oegY-etj߅v��uY�5���&,R�]7}��U��v%x��]��W[���b�r�7���=t+}�]h;��B� )Ca�ܩ<�G����=����F%
u���y>����Ek��_��g���{&.����'�����L&S"�!(s���W%��8߂���{�tY���Wf��]�Zqao��14�#�Ϛ���l��s�BR�z��Z/Y_Y�v�HB|��~5�]Q3ٵͺ^��290%y�j�Ee�bCORΨv�Vh���Q�N�W�����ʯ<āH�μ��{�o:x�}�,rX5�a[ِ13����ۄY������q�+׽��yǯgc�o}C%�#���O������E�pX��Y6�.K�mi�B�h��ٻ{sqM���{PC����ݱr�O|�ټZm��2"�e�U�w_Y�*��5��y�9Rm�msj�5+���%C�gh$z�6�H|�Z��iğۖ��J=:�:������>yw�0�:�?u>ڙ�gpVZ0�*�Gԁha�y\(XDPT�;k���b�����ޖK��L��eE�SL�z ���u�u�U�:Z�P���mL�C��3,N}�}���~�]}��۸#��L��eN��U]��(��Vor���L�w]�C����NSJ�F���"��u�;[��ic�18��hκ�~�vc��ʒ�c{x����i��Hw���Hw���0fb��s8Qv2��H���!��qΤI='!�+�~�F��-E��L6\ꄵ��1Bv|&c<s�hG�9��5ᚭ���qY3�\z�Q���XYȦ�l�h<�ǋŘ̕��\)��Y�%�*'�Ν=�	�kT
R>\[Hf���6��jynm	��ׇ'���{��Fm*f����90���C�v���$�<�{�}Qk\L�P�/�:�9OeV�*�uϕY�鰌O��ι�[�Q�/Wܵ�À�N�/���X��vP�z��\J�җ!wl6�|������c�>�`����R֞E|�\�v]΃d���⮓��>a��J��Ʊ#b�]���|�bg��*N�����
]��Y�J캣���Dy3��Y��-��*�N��iۺ�^֟�fn���>�R(Bߤ�`��Rk�P��w`�.,����Ome�V����Z��"�l��3 �{s��èu�s��i+��Ia�bJƵ'�
��1�n�}�7�G�ލ蕖��i����*�>Lpr���w����5�%O�*��ÃoK��uüA�NbR���(�)iL��( �G~�}%(8��+����=O�A��o�8��.�-6�����X�Z�<f�A%Y�XiKэ4i8i����`c�jX9���vo0,�њFs섀��f��|j�%�Y�W*6)c��&�ʬBL��罔V!5�Y�$�` n�S���EL��5w1�[X��tۖj�AGF�x�dɱ�{�ۥˡ�Er^_�۴�1�q�}���;���%���[c�P��
{Z;�l�Xc%h���e7��7_=�N�
}2�tg}�zR���>\����<��3��E��}���E-N�S����f�<�y{���t�4]ef�tH�ޘ��� ���R�]�39��oj��,�=�)vT(v_r�B���]�-䳪�H�j<\]C0�%�}��7}(�To;4e���IW>���bY�q�h�I��ѥ�Y!�6�-ٸ���ly��*؞�7FU��w,\�8%��0�Z�$�c��2-SMYR�-n�Ѷ�f��2�_0K� ��qu�]9E���[��2�Xx6�9���I���6c�ئZ�ڸ��t�]4�䱖=Z��O���H�a��D묥]�gs����t#r��7�b�7i�T�`��[�dЇM�(�\�Mj����ysSk�
7����ek�-ʺu�"�P�=��Cl޶�#�O������.xK��LE��"�
�c>��pD�Z�k�Do�� Ֆq�j�}�D���MC[&ڵ]5ŗ}���@|s����Jʖ_<)�sD�Y��׼R���A��S�z���z�VZ��Zܜ;N$(gX���f���s�0,Z�j�On��6��������U}�EC�����u3Uyk�0)X���v��f�`����狭��5��pD]�O)���i�-����i�!��Ւ��6����j~o��뵻|1�k}۳h�λfU�m�/jsU�2�9�[j,�����ƻgh���[���s���&�<�ifދ��	��{���s���YԎ�~�hK5��]�KoCYI���{: �a�Լ]3zP@��4��|w���Y#����Cmڦm�EPPNp)�-���Y�l=��6�_bwY��N��\�n7g��
����͗v5m>�1�{�9�5u1�6��8��RPY���4*�D`�P㜁��
��K��e���t�!�V���~|+̎�.��f���P�F�:�E��
���F�a;X��dqnD��D�������Ԫ�/q���oy&
*sf�<�#ʅNԋ;hj��������Ug<��vIZ�&f��(;����>�`LZ�)]tV6;�Jq����wq�Yn]F#�GY�r��5n<C�`5snp�Ed]n�w�Aj.rd�x���q�ryY]N�.T\�`�!x�KW���;�g�2�_8T��� B�=q���EDglYYb�H�����ڄ�!@k�(
�
����%B�E�`�V�l�eee���+!F,R(��Y*6�*�"0�%kZ�5 ��H��XTl�����aZ��Db�H�A@E��+PTb"�ʂ�Z��
T�5%)e�JȰY-�+�b�+Y-E���T��*,�`T�TZ���PZ���mJ��(�(�YY�m�QR*���%DTX(�եEU����ն�YZ [d*j[`���ƥ��%V%E(�Jʂ�26����E"V�%jJ�JѶ�b1T�PX��+VF��(֤QbȱdTEQ��"ZQ*�hTYYЬ
�bֵ(ȱ`*���aP��J�,X�,��1"�m�̹��AX�T���Vc
�%T��ص�
��fc���*²�.��G�4;n�(}�ru���O/m9b���Ɍ(�S�Gn׹੭�ղou��{� mɯ�e-s�Ys�@L+����g.�Uw�- �g�i	�eh���+����Xǫ�L����>u�3yߨ��o+:r�>�,�����m�ܾ�����^ �cU�A<��j��s�M�U*{y��S�`0�(3��f`�s��~S�L�>^N�xs���yV��w��b�F��Cu��Ѥ�-(����8΢�YP�r���B43j���7���6��fͧ��<���S7�*��_L&��*q�d+�(�b)�L�yn�Br��ch�cv�[�P8�/%�`�f`�\]t�5��D�l'�}6��G5�yɞ�?z��3#=�Z6@K3����ڨ�4�$���)���ϖ�����L/�cR��,67�4#�6m��ؼ��η��aB�X)uH��K��!�Y�L���������.������|�KA�C�?{�����l�&e�s�I�8�J+�۽9�L2�V�δxz�sM����O��U���T/V*b��ɐA>����	�n�PSզ���^J�fg�t�XF7ݣ���4��1ׯ���7vy�r�ISL��
kv���l����MZ?1��g-����_�����yi�dM�MҮ���������pц��#5i
������.W�9쩵
�KBW=�X�y5%NXɄ��-h�Z1e�=���7��zxt���:]#�âJn�Z�)�����/i�)%葘�\E/S,ض(����i+��.�#�<kwu�J�c������� �P�_��/#u�m�S7�<�
�3�:�7���΃ܦ.�H���')o�q^{�9�r�TP������>��zm�f�j�>�ί'��9x�qQ�{Bq�Sθ��N������L�Pk�
/c�z/�r�h����^�諾�2��B�����V�gk({N-��J����0nWb�׶6(`8u추�S;�CN�W�g�J)y��lgZ����ky�iaiL�������qf݇r�z(y&'��ܴf�c�tCqj0��-�M��㽩��5��Sԕ��.X��6��D����	�Ļ/�.[���NM�[G���F*����-�JQ����h��h;Q}|)Ďy��,��Fc�([���ǜ<���G��*_L���}=p�\�����?}J�̽�
8Yi�Xo��?)��#�3�f�~m]�yP�<�lV���$�ԛkr�mnҰj!g�?v;�͜�(��#��:\}{h65}�*��� �U�Jb���F�H����7Z���[.1�a����GNN���
%8k�l�]�s�e�X���Y\��G�wRq���>��E���&u>[�PL�zĻG�Ҡ$��Ds^��8<�z/=u��_?*���ޥ Յ��0��zŝyS�^
e��-2�'�Qk6_�R���gf�6��d�8�:����d����AU�y[��Q�=tt��55�󍎩�w�:-�5�ԫw�0)y+���	�[�l<�2�����k����iŜ���!E;>o
X7z�y�m�{�m�1�
�-\��j{��=}�'����([R��||)��7ۇ}Iu�Ϋ�ݲϸ�;>�:�ʄ_��C�\��u�]T>ͬ��t�WaiC��C�x����_�;>���5V�8$4��P�l	TD6��Wx�=N��#^���M�=�#Z=�F�{ՙ���#3��+��#Ta���!��gT;j�lr8��6��i�G���yp⻷b��M=yK�7<��DfK�\�� 8g�:�uæ��ۆäB��v��8�{��nO.�ن�"��?\��������L	״t? �iM^�Rfrw����7��Ud�)�y[C�m��g%brr���Y8d�3�v'��	ova�ǣ�_y��ZR�̥�&#}چ���ޮv|S����:=��R�A��f��֝��|s���O^P��eieK$�V���b�;.X�i�-�O�	lue�t�������jw�0�#��wl_[���f-6��֙ۯ�Q|�n�h�4:}jf_EJ�ۢ;s��9W�&�x��."���򫫑g��VX8�{�k+�n]��#,%�໴�>�';��z�MwU�g��Xzj�Gi �Vi`�-�KWȲۊ�~�,[�$������)�z ���u�ut�+�t�Zj�ҁ��x���ZYÂ7��w��#(K�(�<J���Q`��a�\ꄵ��y���<xV�	�L���ut�zC�Z�`q���/E��	u6V��E5xl�h<�ǋ����GAX��ז;��'I=U3Cg��yX[H�`�.,�����<�yN���[�[�q��xr�:<wwn��f���{<�(Ж�4H���@֮Jk����3;�Ҝ=.�)�����Ss�^�e�ǆx�'�E�a����72�� �!ӠAk5�\�e
g����=��3�N��ѓ�g�A&!���5S"�F�C�2�dQ$_��qV�x�}�)��p�N����^4���]j�n����9�ҥ�;����i�6�z{��{�ŋ��h��ic��Mi��S2m*]�9��ķ�[�2����v;�̴���4�=��b��Ϗ;���M��-%�3G�@o��B���d�"!��Y�b�ݍҹ��O���̎`Fĕ�S��Hj��P�lL�0��k7��ol��m^�{=�;����p^5*�.=���ɽ0$��*�L�II��8�"M�w[��q*.�Շc�W�:��,��J��=x_�֡χt���(-��C|1׭h�J����7���2��d3
<��s����xB�y��uX�Fz�^�q�6�T��<�^�F˜}µq*|�H����>����x�>��)yև��h�}�F��Y}��ӈ��լ�>u��qYӏgB'�f��"%V`LtJ�d��5y]�<Hh�����Dal~>,�L`ܶbu-x����������フ�;}2씵,E���x,�l��i_�lX�����E���+���J`�]���C�$6�8��6��z��p���ۈ���K�Z:|��M�1����
��F+NB`.�ɨ
&�z���YҸ4���y)S��F��C
&��3婎 �짾�#��$z&)6�����Ox�V�VE��o�1+Չ�Ķ�V]�.{G�����;ܿ'=�4T��f�����������[�
���_N}N���t3h��P��Ң0ǵ:�V�ǵ;o�I{����ʚ�wJ��Ϡ�ݩ��M�oA]�b;��g�}���ʫU�8��͂��	��XTF�K�`��M�\^_[�E9S�����lj �EE'��WK�{�E���ڞo<s�B�X�H�@�<C�K��!��P�LW�7���R��z���)�d�[����փ��t��LGg�E��d�,�s�"Hg�/vm����]<��Ʉz�C1A�����w������A�*� r�.�d�p��P��Ő�^�l�=*���~���.����[�s���i�<Y蘗���x��Q��ע؃��ڹa}2��<8���ݔ��ґ~X*WKi�|bا�n�Xs��i ���VkĎ��,���k��iWk|�������a�RI�e�<��V/_�����<mt�y�\��S�ى���Y�3{�E��T�����2�#b=h�;�x��<�zy3�0�O]�����*ޡx���OΡ����x��^��P����9�>�t��.=;�'v���]hc�c�iy�6�z�����)�싉��0Ջ�����ԍ�z^��jM��vn%]mI��]]�� ��2֗L[�n^�XW�໘��|7jt-p�mGX.�9�L����ڽ�X�|���`X��(Ȼ�8�n8rWۧ���6��C1e�*�vS@�m+mՌ��}�{5Zt�(NE���yc�S�A�1�K@z�g�OB}V��u�4�ił���P��O;��>�)�ݟn]���걵<X�C��D�t1y`.�[�o8T���0��阜��;�w}yB��[�0�U�:���mk6����0�E5t�j)\U���|)Ď1R%��,�K��J�u�M�unvӨ:,���Z�2��t�-4�:��J�̽�(�ʯ��.9��vl���n�$�o��FX���C�:�^6�锏\�G��5���'��w�Ft��#)O�n`�����e��ل�y����;�� �^L�xܳD�h�7��ʚ�o�GlYvY��N���vȘ)�W���������.�z�ysb)M��>��<r��N<�Q��:�*�T=��I3@�8nq��2�ӕP�����9�N,��Ľ�������U�l�Q�R�{�Q�\��>���s�ZWN�w�p���<�y�=Ekv��ܫH߯
�7����J����U���P�L�D����I
�k���:�/.���5�������m^�k��n��v�}x4)���^��rw�������|�I/��Z���0n����0�N�W��6��E�ؙ�
\��}%�F��M�ÖL9������*�YV�i��f�L�ە��Ǖ�ؘ��5���śڽ�$��且��=�{�O=�Ǉc���O�k�S�:�x%a�����rCO��(C�"!��hK�]�t�Y�2�����U��rg{5�+��P�9�"�t���ƨ���B�����UյH����;��&���v�}j�i����R���(�I��ޭ�of@p<����&�_1��c^��o3�}K��P�������^�U����*`ַ�
bu���.'�D��A`U�8�x�ujiO�֝��w�Z�y���uK��K�����x���L��%��ر��.�_g>��AA�t�&t[���W[���Ĩ}gh$z�V�E�=u^�wQ�o�JK��|���)�þ�;P�5�}[��w+�'�)f��`���,��F�үv�0ݔ��ރ�106�2����NX�/�ޗ��g��<N�ø���<5�����:�mZ(2%H,+�.j%�Qp��auC����(Nɘ�W�"��7(��fu�i/i|g�iyx��\emQ	mw�9��Q4v���Y�`�*߽���ӆ�2��5��T[G��2u���Yn�,DM���y��.��ؙR;zq
�É�.W��i��Q�^�=�� z(>�� ���-Y����v��M��7{�+=�hL�ۧ-�y�1k,eI���A�
G��m��-�m�x����ݭV�"ŕ�Ŕ2�y��v�ϓ�sk~2.>0��mR�N_%S�kxn������jD���Z�(���ϨS3�M)�m�5���o���ہ^;ݞ3�}��Ϥ�7�Q�:}�G�����Y��@�/Y����
g�fO<b��t���+zn�k��K�JM�c��fx��U1q*�z�ø&Y,ٲH@k��;�4�)x,��k_Ii��w.��o��Y�G0#a�ȃ�����ڭĬS�T��l�z�c����f֑���|;Z�fa����|dݘW��W&c$��}�y�Y�m绽�O-���]�2ѳ���*ac��^������ZJ���t�=M��0ڻJ������x ��ᰘ{ժ�4��S��g�V�|.}U�o'�e�o}��jQc�9�/<�7ciM�ϻ�b��lmS/j1z:� п����5Ȱӻ��Xs����r����mf(�/�0�����c�f�U���&D8J�	�&�Y蘆�}�"s��v���.�yX�v2�~蟆���-�����q��
t��(�ׇx���ߠ�9���䳪�-�S�4%w�ډ��Y�u2AY9mj"ڳ���ְ�|�vV����RS�Ѿ�Y�(,
��v�ڵ���p;��]Ew%��G)�Gyݝ���9�u�pYF��[ջu��0S��O�.'�k�G�ח��ơW}W�^k�q��[s�η�iu/%��]p�p����u���BI˸t.��xƇ�����h1��T��VPV=x�:N�-���U�IƉ���b�re_����W�~�
^��?	�Xm`6�wT�K�~�-LtEh�T��?x�+=J�f��.-�]X�s[��굞�� ��i@6lr�!�Y{w,�hqDiĹ&��)���Ҟ��
9q�(K*�Y\�7�\�dh��# �#=��as��yB�\�Go���"����5#��<]��o���hᔙ�\]u?"�C6:��,7~�Q�1躽��U)	꺯>�aəS}�<�7K��$����7T�q�<�����*� �*��1v{&C��e��t���^�7ڱ���.�Fy҉X��u+!�������Y��=��t���G=9+�ZĝGQ��<���< ���¡��Yґ~J."����lS��k}�-$G���m/gD�piȶ��60��E��il�x���b�_�wP�[�\=�2�%9�n[nۧ�[B���j"���]����Vec��{é���c����,�]�}g� Ѭ�iW>�����;ع���q�F�O!.!LudP,nW^:-��`!��P�) ��l�wz��v��ע������O[ٻ�,L���b�}�f��#A��W%�z��I�(���(�ʋ��a&<�Lq�1�#��O{�/v ��$]�:!�,�K�Cx�K��C���ُq�;�d�����DWc���;�5�s2��uZ�����:���sQ#��::4�(ȜkO�V!�YP��&�e;.��W�Eui|ۘ��8i\���.��9��56�����@.}�q]�(��ⵅ@��y)�r���8�*s�7J&Ns�wN�j����H��9n��,p��ラ��r�+{�y7k|^]�q��Ѣ,���V�^<Ҧ�υ@��H�j�]a8�(��,O�kU2P�s�]�gFIv5�Ir��4�,�J����5�Z��g4)R�Z�\� �t<����'�4�m�.���
b3�[9Ց�K���%�K�5�&�Kxe�X��E�c��u��۝�3B�ON�r�[l�j!>�p��:�hއuRhgi/�+}�"������͡tQ:®������e�I��uf�V.Y `�����_v�㭻d�t�^U���7��Ȋ`����Ō�����6t�]��`�'��$��K��	3^�6��j�Cz)6�b�e�OK'����wԾ�n��ߖ:�0��6�]��<����jV�*��݊i^MH�Cۏ��mǸ2=�jl��,��fq\F#iPZ$��2upg$#�*�]�:��GϕkN�Y�b7}2w�NctP�2#GEf�����L|sZ����z��f�殏:�����ZS۽�¶�`�w\}:��ZI.N�-�R	��}�3;�Tf��׻�2l7�e(�����I�W	6*�yIx@�S�;Fp9S��V�v>=�(�v.U��$�v�-�{�L���4�R�9����&;�R�$2�rڙVt���N�X ��V�5����:B7�&-�ځnM���]��N�HؕU����a��{rLwxV���63��q\C%���s�����V�����J�Y�V�/����{j�+.s*�ԩ(�75ҳ����C�UX}�S�}]gtM^�*={~�	R�5]ZU����ê=ìs��^��r��Ȩ\���n�˘HS�V$n,�>I�:ti�u�}j�b%�b�<�Ra�õ�[����7�-�b����p%���ŗs	���N�;+RG��]ћ�0�S��}xܷ݈���,z���5�n� lyt]^ڒ���`0k�P�L�%���b����;���^�Cwܮ�=qh��ض�K�p�ˣ���RΕ�5�ڳ���F�����|�Prʀ�Z�AH�KEX,"�%k
�Z����
���1�r�e���� -h$P��TQEA�b�cR�TU��PU"�1���#H��+Z*�X�X���C�
\��H�UEE�AE�",q�֑+E�(���*�*EQ����-�Ȫ
)-,DQcl%E�krъ5AH�bŊ�*(�H���Y���ذU�1�@\ID���*
��R9`b���B�B���LeTD+U���� �E��,Q�-K�UAEV�jh�d1���bV*�Y��[B����b$G,�V
�!�TT�(�U&!�VCm�2(�UcD����QLB�"���
��+ �;F�]Kao&�v �`��k+sW3��9*֢;"r�lC��c�4w��n�t�;j<�gw�Z�x����y���/���s�G������v�I�G�Z�r����@u_�m���f��
���(���5�%_ɘ�2�:(}<�zא�Z�ϥ?:���b����(=���:��=��ە��P�]��(�{#���'�m�hJ��Mewn�:���Χ�q�����d��l�n�\g!J��ł(����Y7m����+=�粛�0�o{d�Ӏ;�՘�'3���C��2��� ڠ��s0o��ZY�y\���gq��㢳kK�f���f�C��D�z�`1s�����χ��OLo8����5ooF���������|��O}~F�|W�Z3���X��'/Ώ��-g���z�m�m�^���7ZD	��<]G����V��*ϫ-r��g�I���}�r���{�g2��F��+	|Tz&��Q��e35w�_q�����H��9W<��vMv|���yN�㑪xE@�U�nf
\��Vf��H���,�yS�^
e��G���_7b}�ý���LY�b�*��z�U*򑬭n���A�0��Q�]��n�|詁�^�aܮV�[��ڣ\�yv&:dز�\�( 6�G����7�&HC9mn�
e��$�hU�%U`Wm���Sz��%����&wH׏;�K�h�:R�6Wl �{]h<�M^
V���:�����ئ(E�t��9Nvk�ǝg�y���=I�(�
�cX(&E�6&\�~�]í{�x�q�|Jc�,�۽��o��]���LY0Pv��49�-+�ywl{WYv�)�X��޻8T���ݗ�K˅�T������ʄKO<�H�3���/�j/%(�8�&fe���k��ݴC��u\��jB�Wh���Hi�8%vĪ"xM	|+���K��
6;�z�����s����S&9������^w��Y`܆���hVh���_T�e�����η����^ܖ�?#�{�K�x9��Q�Om@S�+�z
������G��z��;�w���E�}\g��SVL�T>���}^x���Z�)�״΁���[��T�JoW7f���S��b������a�k���k��K�����%Y�~�DW�����w���ݳ/}N]���l�湏��Zi߮��&�ł�
c�Y���tL����U��>�p(��J1�	�����l/Wj{�o���k�z��3��؃:���#Oj���e˙u���F��xs�=�n��8�r��BO���YI5��3 ��J��2�t�����g��U�6�u+Zfdx�r��|�04���Y�Yӭ)�l��a��=C&���s��଴a���,��sݭn�6>�N-����|*P�:�8��b���jd󡚼��z^[=�����=�=[Z=@ԯOT��k9���Z���\�K�����`���y��P�����z�޼.9�.v�R�Xtq!���bKG��(����SW��D���x������W���n5 ��x�����f��wkU��X�����f_y��v�ϓ�sj֭�<�%�{���KLs�x�~�kء�$��3�\��]L�)�w��7;9Z�2Q[�:��u^�M���a��ߌ�/ǄQ�<}�fq�	�x�:t!k5��s]���UDp�9H\���גfJ\��n�~�<y�-i�"�G.\;.�g~6I�3����H��8�φ����4�Z�SR�\�x�t@���B9�R�2Q���Ĭ&֯L�eR��0�[�~k`�V|`�4�D�b�;.�^�7嚰�oZ�3�`I\�W&c��Ao(j�s9�r�������}gtT��l��IZ��'��[6��У���۴�������N��@�Ֆ�M�)�d�a�'opB�:���J=��V�Wq�����m����X��:�/V�1�]�Yo�b��\m��]����s�1�g�����J��l�}�
�_Ä<����U4z̞�v��x3����� �K]�5�q�]�w�^S:����r�1�S��g�9K�vu�iV�������|����/\�W�BH�2ޕ��/k��#��F	��ԽO��d���rc������5Ñ�711��V��0'�/c�g�C�R-;nnQg�.�џ)��&�}�O�����P�>�E�`���b��2��Z|q=Y��릾Ӫ��;�GG��"9§�Xh{�&4�Gr�ᄿ��:u6�uSh�T!�t�d>��W�h�%��9*��w��kׄ>�B/�R��ܲ��֛kUq�}0��*o!X=(Ž-K.��R�o������^��\/A�,6�h4��O��p��/)W��fυ;�#^��6�sm�G0�ѣ1O�R2�~��r!�Y�uA0��ӉrLKb�*�ꏲ���[y�u5���j��j���_j/*��Ɉ���5�cw��ږ��;���:rӬJ*���Y���ΩX�ϚI
�2�����)V_K��hV�n������@�]���>���ڟ__c���~7�m8�����^6v�.���4��b�Xz7.6����y�ӊc/�gU��ל��3�N�B�:=���a$����g[SuwbR�w+;������RŎ�~���r�0�1�u���3�OO�[9�e���c�c8!��nwGԫ��gå"M|F�օ=����g_!:L���Xz�z�J�����r�����o�����"V�<K��V��W��z:�-����d���;zz2�+��T}&�>�X<`������¡����:R/�)yh��>�Þ>��8�un�>��^�u}$ڗ�y� �q��wl�$xq����OR�c+�rǟ��2϶��x;X�]���g<���_'��R+�����3&���$�ܡ�BvR�;�غ(���qr�瓮��5��,g��r��n)�C�X�pm�x��u�N�CM	Szx����Ƨ��l��-z�	g�o�J)�]j��G��2C:]�q>���t���yL��|c�����W}~�`u�|�8�6	��J��P��nWm�qg��`�#��Þ�y�t���r�W��L�J�9S[,WP�k���r�r�b��2#�\a'�<����fN{�<�]����6S8|��Qّl���鳧%7]*�Wܪ7�k�{��e�H�N����i-1m��l��ݪ�]o��S:�5M����!eG}��i�‍�K���or�f�S�AB���N�/��i���Y�gpK_��	[��v��/x-�3���α3��QYE5b��LT�*����x!�U�#��í��MO�����.v	�]G�Ύ���jWKP>(2�#�=w�<�-��4o�/�[�:�3�F�qiX��N�d�j6������e#���G���-�K�����h3丏ZD6�ט)s��XY��a"�y��˵;*@��geq��X�/�5�x��.�&{�Do��h!���ZԹ��)Z{������b��;V�6�GwMɊ{���W?|�+���6��҉]S1�#�s����6�)Y���I�G�ˢч#|�G^Ӽd\�r��S��*b�z��5Αi&�w�]��;lO�ц�K�O(y���񓖠�/k��_��g��-p2�#G�	a夅k5�_�댲�~"�������tᒽxd���s��n��"���'$4�P�nU�&�
��ϴ��x`��/iћ��]+h���k�¶�(W��vu�5'� ��Tz+,�CORΨv���@g�c��f�T�~V���IS���uԥ�}��U����E���\�:�f5 ��r�@�ٲ�#��`�`ٰ��qv����+��\�e�t<�+zoX�4�VKs(���憫"W0"�4�9٭e0y�Хy���-w�|��@�x�k_؇�dk����:3ޙ距<Ct��k����d����5��ͳW7��GM��J�C޳Vn�s��z�G[��>�:����E��϶zQ}�:_:���^B��dK&���zmi�͸pjԃ���m5�ǥ���vH=^�OCX����G&b�c;�����*���;��7��}V����_��tS*�s-��ɗ�������tg����D���;���d�q�h�gpVZ0>����l~�ԵsR{�M�������"�L�E_p0���e�N�(K�3W�W�U���Ɏ��[I]��ɝ����x�Ƽ^
��ȡ�xV�aZ�V<��za0�.uC�'[�vw�t����:�ջ=����L�<r���4A�"b����d+����YȦ���ǣ~D�`S�n�'3#��U��qC�0��"��hm�����E�+��*�_�.&��v�!D�Z2�&p%��g9J�u��O����s��\�bD�%}.�5�����e�L�T=�߃f���;�'�n�U���ð�z�-�*���謖n�xb����Α1U�!T:��*wh�5$���M�M���i�-�S6ҕά�0U�<q��S��9�h��p����Q��J�]���;5\:��	kr�1YO9KW M��w-7_9���ym����_ܧ��!�}[JD����!
ìP�@Ϋ���~J��۹�9;m�P��kP�^Y��;��
^��U1q*�z�ù2�d[���y��sz^wGjVT�]uBo�܋�II��������z���x<+<ѓ��2��k�{(Y}uG���adv$Y�u����嚰��j,��0$�IP���k�/�E~&�:}��^�09J.C�.��/)�����p�%C�g�*�̩��c�r��^sO53� �`Ϸ��K�/�p��aC<��s���ڪ��<�YC��	�����cE����Z�u#��4��TC:z���UBEz��um��mH�ԻVlw�e�t4_o^e8�*�#j2�_WV#�^=^�5[��'�8ǈ�ݱ�������,��ʑ��0w$�M��G�a�.�'�]ar�"��l���l��Z���z���,݃�&e��J1�;���^9���OT:���c8 �ѝE���+�d&�!�U�ye�7��/L�\|`�|'U��A��](P�s��WmZ�m^�J���5z���[�ٷF��W�[�n��c+W7�IF.減�a����*�xC�8n�.
�y�z6Cl�b��@V�v��;�9�q��Yـ�W4�	�,�`L��iug����վ�|��.���*M/i%�A}0��c	61�2dC�wd��N_{:_S�D;>.��u��6�i��R,�����\^�j��^�X��[�j�H�x��'�y��9�9�WrɆ�Z�4�K�`��d3��v��^��.�c��|n�u<�ʄd�d�g���.y���(]��F�H�X��3*1'�u�`��A�>I��B�v+Z�ө��m�sT0�����3%LX��l������.oI��c{���H��܅���a����g�.�����s	�9�^�u��37}^���U��O&L����R8:RiX�du+!��7����V�\Y�od���{o;���9gWcNs�kF,NS�@�I*)傥q�c��Þ>-�I
����9w�9��:��t�����l��$xf/�C�5�OR�c&�M�R�n��v���XE�:Vo�H�R���W����	��6��&�C�*��޵���2��3N�f�V�J7���]q���Ծ��B/p>��j��I�j�+5֨&.��i�j!5WfL'6�u�Ru�usc��FԶ��p|��</I��gHt��G�ub}A�7+�����;l���	d��r��_�;�|7Q�H��B'[��x�od�0��k�Mf��xnV�C�p�pm�x�E��,P��f�y�\�ܿ9���VՆ^��11w��*��¶��Mu����u/�!��)��vEğ`5�)�-o. :���&s+�2���,���va���X�:�������� {vR�ѹց^f=��k�WO���+��J�*�L��\:Z�ly��r�\} �G�#�]1~�(mW�[��R[�Ӥ�������-�3��^u�����GMX��SK�)���k�tj��j���SR>�H�L��sp?��������-#� ]X�Ϋ�x����;�]�ʠ�A�}o(�e��y��o�ل��5�|�[k���X&R={Z���~�X�%~&� &�����*�]M���{3esƖXY��6a!���:�z��i�:���ķ�n�v��G�QD�J#�q��C����;�5yLwV��*��+�ù+ey0y���jˇ��_4��2��Q4%iਝ�������]����HIO��$��IO��$����$�$$�	'�!$ I?܄��$�$$�	'��IO�!$ I?�BH@��B��$�	%!$ I<IO�BH@��B����$�����$�$$�	'�BH@�zBH@���d�Me�.m�c�~HAd����v@�������x����U� �B� Wf�)T���(��U Pf�`�8(UR�sZ+��v�v�L�X�amCk�Ul	�wc�@ݷQu�A��� ]�mV�6�-e�ù]Q�ƅe��P�Qsc�[bM��2��Z4��m�#i&�8�Zmcl��Z-��*�;�l2$[j��1%"��Z$�T�h�cm�Ap;ulX3f֢-�k�     <D��ԥIM�= d0� O�T�       �&d`bba0�!�&�O��R@      �`&F F&&	�bi��J(��A14Ț��OS#FC�R|��=�B	?�`I H{�Id$�@l ���C?�?��Ā�Ԑs���g�O��2����������$�Hj@�$Q����$=XC`#	�J�*H$6���{��Mh�_�������{H�I<ဳ��=�d��LO��g�	����f)`�{�k��}��o>�s��b�̼��1�z���cSċ�V��$�Ue��xskmJ�4:���*W�]a���K�3.����0h
��6C��y 7��i�{jfL�lhw��O�
�R�h�(���W���B�ӷux��m��p@e�&*E5�b���v`͵c*�aXUܔ��8��C�S���+0e�W.��G#�ͱ��u��RY[�`�&�d�M�ǎ+&��_��=X�wvĹLR��c��<�ǻD��)�Y�y�>Ik3y�f����c/v^��!(۸]��.��qp�4��eB���:�F�p��0ǩ�8�w��G�VV���n�LeD޲�5a�-���ᕷ[���6�쩓M�Ӻ3b���h��,Xzj*���`b��;cV�z.}`�e
9J���״>��,�Y�)��R���p#��k%���̓NǮY���8��t�޼�H�S�Xh�Q�F�m�t���M���N����<M��(wW0:ݍP��Lj�@�D�v�85����Z0�����ͦ����R�w��x(��u��ݔ7���M(U�-�N�C��/�7m�[V(mBt;1�?7hm���	�-��2f�qU��3y2���I�1d�tf&�nD��)�*�a��B�s�W�*%�t����F�L�֯.������ڽ^B6MX�&�f�ړ�P�(͚�����׋q+��l$Ixz�|SѷVtܢZ�Q��dC���賷Yniբ��P��-j��ख���̫̼�T)�XVZ�h�ZR�v��=���[F�5���ף8�ۦ�ۡ�Hd�^ZvA��q�3�*U��/��V/�v�t��&la/i��߄���z�ևE�0��<uy1㺐��ِM�#J��R�;N���V[�a��q�3�a���L9���i.�e��De�݄����YȢQ�Nvu:�:�O���j-��*C^GjkeX7�X����[�\k��o2���L1a�	Ӵ)��WG^��+l�	%3�u��A���LX���Ym����kU���ʟ֓�������ֵX�d�ŁC5��2���j�u"5ҫ{:�Ӻ�5��X���5�����ė�"�䵚� ����ѥ2�V��ܔ(���ڡ��i�Z�䫠�n3��1
����Z+Mok)�Q�f�����QF��UO.�.ȱ��/^Ő�V�{����dy:�Ր�@a��h�Ԡ��Æ
.��xC�}��Jς}�g���:ħ �1>t=�����F)�a��{��5�0x|Lk}s���m�Yr[<o�:޽��Ll�6kB�ޕ��M�ND���{�WvX���)U��Ww2�lG��^Ν7��,�}r�g�VD՚�Ï:\Ɏ'�Qr[�T���s��m�-a���{7_,F�e�؅���Fn�Q��E�<�@8���rG�#�^��G��yk�1V��Bk���o:Mb-�����Y]���5ui�7��Ӝ��{T=��(�ay2���c'`t����D#\�^�Xz  Ը(ǹ����!��.���ҳv+�ε%�;�JZtJps2��y�G��B��J��_aR�+���1t�M�₮兴��@�������i��2�5��=1T��ZV�mcr��R�;�c/el�.��r�f�a�oVfw08�L3sst�1>&�3�y(���ӕi�j6�;7�TlP����f�rhr��;�)�@�wM���Z��^��/�я����[d�y�o2��= ��B�-����SW�V��;M�n�{|e%j:�t0�n�[&1mv3�9u���<�����u�<��1�Y�ZԔΚ�0'@����)����}h�[���3�I���(Inhz�E;��M����%<F�}��G+c��֊��w�2�7XF�Q�!��d�K���=���=ͬ�}�u��rxE��A��Ǽ����gD]��a�3ie��1�}u:�μ��`f�!ǎr�Kjj�I;s��gWYCuӑcfӥ*�d0mE�r=�.o[�eu+�ch�w�,�]�H�����c���I���b�"��_Sf��N1}�.�	��]��������X��<� 0������ƽ��Ue�)�u��8���猭��G�X���C�_nU�D�Ԡr��ވ���#7���/���i�ʗ�Ʈ�Î����6��ƺV�.��|&;�E\� ܙ�)=t���72����p��r�y�y:�C�1�{�m��wC RT��̝�j�P�s�q��*�a����!ar�L\��g(tR�{,�rѽ;6mNR�Q������F��;�
��=$� kNoK�S�+���K�i�:Ɏ_
[9;�(s�O]b{��9l/N]9w^8I�1i�n\�MQ����+�-ͦ�Ø�#M|ַB�F3��'*��6�"����R�xy��xE�흛GI2�;/����%o}  ��Z3ʛ���d��Ȍx_i��/j�D)3mѨ(SWR"`&U�� TS���yH)Y�ivĕ������Z��AU�����3�}�T��l�������@�} ��<΀��C�{�$'�C�=*�}�2�$>c���{��z��}�Y����B���X�Qb
����6�0ܗo��g[���VX{un���a�y��%g�*,�)M�Mи2gH�9��*���r&IY��B�h�v���4n�V)�b�0M읝C�z��\9�iL�f���0_E�Ӥ���ze�˻��ƙ��!6c.$�o~Ӂ��]{ٍ���*V�6U�dPr���q옻n�[��Dq��4F|k�뭥�s�'Ckp
;����t94E2v�:��5�
�e�WO�z��&��5֕��%Y��̽��GISJ������!l��6I��]����Z����F�JWV4慿l7���1=:h�dn�Q�0��5�lY.��7f����ܱ��m�R��db;��{
�r2� �kE�H����Q'5b�t-Mșb� Omc�]ܗ&I;[Z/�ݛ�;*�
���4թL��؝[�{��=��/4�D
��)��9�,�/�U��um 1�i�u���v���&#u��X�#.��t�y�Fu�*ni�38t4�J[Һ�v}�޳)�w`�IJ�u�n��5���-F+g(C�A7{��!��^Ǻ1i�zZ�l*jĶ�=��qĕkNL��C��|�O�ՆH.��	��B�w"�؈<�dފ�lL���QV��)�nU�\���6I��%Xr�d*�N��}�d��eN���$�������D�bZËa+V��,���of��i�ǹ�u
���`O���DU�vjv�{}AV"�y�,k�G��;y
��E2gTϰ����%��2�s������U�@����  ��b��|��\�w:]��2�>8���	�-W}�����=}L��K���1B���fcB��n�m[u�w�M����a��b��3�Z�I*�������I�$<y��Wd��0p⬻:s�q46=�e�E=�V��'p˗�mv���t5î<-j����BLPW����l�
������Ѩ�Ԛ�Y[��ܵ���Ɇ�Xz�ߛG
��L�,UH��|pJ|WZAuf)�3;)3T,���,�5b���м�m��!��t��'jɳR�Ypq���砛k���U����\uA����l�*Qh=�����.�m�)�t��\����k��5t�|3��6->t|�P�P��Jfeִ�Y����/b�V��Ɠ��� 3�u���	tH^�����y���@ru�f죊� ������P��1Rd������m+�L�yX-��2m�5����z����H������H��7���f	D%3�諒n��l�$����^S�@�d'��lv�=%EC������yȝyo7�Tw��2N��"g�Y��#c;1B����oe��S�E�ђ�H՛��(�MKò&����e]��F��{�R��O������T$C�B�b�b�W-�pҀ��j�0U��Q�1�7�5-i�J��c���L�Y���XE0�b�PkJ�,\b�ZUm�U�1
ZR�pb���k�3��{����U���`# �V�}��������u�~M~�����D�բi�J7�NQf�wd;evε�ѵ��A����ө�἞$x��M��E_��-�d�����r�Vy~�Vz�k��ѯ���-���Fu��C�λ��&������:H��i]<b�����~��]}� �k��m���uyބC����F�ѧV�����k׫^o@sPe��F\Y"M�K�xU�u�zׇR�ӆ<v��mgl�a����_��Y�Q��^�l�����E-�yȏ����4��z�|Kwd	��޽�x{�U�|�y���.s1M������� �jԷr�5�:��_Fh'��u�*".y�<�_[��9�ϝ"�>�p�-�x��q�(lw�/v3�DT��}�޽��Y���R���	�<���+#S2��/ã����(݋t�`���	�u�\�h[�����^�J�ٗm��X}���f�>��36�fLT@���%����Z3D��Yp�LL� �n�r����m>u����G۴s��D�ܥg[ԩ��e�~�N�8o���G:TD��^�w�p�ma��n[�t�)��.��|�ݦ7f�{g�2��<�Z��9�.���sܲ��[�I,ι$N뇉�\=�z����x2k=uָ��GG�ƽ-}�T��Z�U(~�YH����X1�z�2�����^�'9e��N�!�AJ����/<֔ה���4ʋ�V8��g���-���W���
����3���x�QLW
B��T�K�EZ,!^%&P��3�u��q�8��@�T���z/^���u�ӥ۝F�!g�u�7uf�e;C�0�w��O���q�+��E<Ǜ���2�yN�&ޙ�틖�;;�4����w�n��Vs�w�5�öm�s���\���TX\S�{O�7����ݰQJ���8�˥�ɪ�t�a���C�"�>w���;d�;{�W����J��N���; PpWdT�"���t����Y$�C2\�c���=���s��6�u߳Ο�L�Տ(R�=�d�ϖ<eg�]�A�o� �٪�L}HWC��#���N��,�<C,���=oi��6�4^�Fuٮ�a�yL�s9x̳Y������F�=Y��g�M���;L��~o�1C(������9S�msO��S^��Д�pn�K3�8Xvk��U!H}U�g{� �)�zg��z�I	�X��9�f:zM!��a+#����m*k�e&2���m�<L�3���s����T�L'���.h�}u��'<���N�T����ɖ9�Ӵ�ŝ�����4s�"�5�2=54���=u��)8�IYƧoL��J��0:�ν9��_Tך��y�S���͛���g��,���j��鈣�m�0��R�@�qd��[N�ϖT�ۡC�t��4䧊�pq��*� ,&a�tS�Q�;ͺ �tC���c�5��Kp�.#PӼ7��*�v�A��4�.�W����g�%���Hߙz�~�����Y�cw�g�f�n�K��{����h�7��5�&71��]dp]�H^h�ò�f䭫��es�/-�oM�!���s�K M�Aȅ�6�&B�oXu�kYɝ�p.�2����+N;4�R*�"*.3	Q*c#�ÀX��*U\�*��U�eq��%L8kJU*��l�AT�4��I� �U'_,��u�O ��̛_5��]�)�z���c�Vg���[C�*
�"�Wי������^�T��P�E}@O��*�l5h�8����4î���IS���Iյ
��t�����C[��e/Ve3���kt�;�|�x�j�{p�Wβ������iSl�)��0k�v�SI��q�������'6�[�[�f��U�'�Z������V7��iw{M2cX�����}�,��d�SVєڿK�?:v�oS�k��4���;1�m�&\1ES1�oni6�ä�)X.�cٖc�;fP�KWn ���]S���=3l:W.��<�5�&ޯ���Pͤ��v�7�e1�:Ci���
��u=�^8�f<�O�n0��8}�����s4̌L8��������0h"���A_P�ۆVc�qi�0�b�o����L��)qL�o�]�k��ͳ�0��8�[�0�l�:J���. �v�3��w�k�M�M�+��%�qT�gvk�4ΐ��ܧE��Ӵ���-Ѭ�Ȏ�	ѯk��\k4�o�^�o�w`Rp1hf>;y?����������m�8�f�*
u����X�'�<@���8��h��X0'L*R�{���U=k:+�)
>�ڷ��㷉{�Cz�5�B��3u��Βm�0�}b��;��UQ�+��!Q�η�u�m��a�;jq�޳7�w�U G��|����̒�i�QC���z������a;��Z�|?������&�a<z|��pa�Ӵ톜�ͧg}gz���֬�e�HqКߝc'O��C�;J͵ߝk�,�:�0��5�]c��7���*,�E�s}f�)�s�,��tu�i�n��,�w�v�+þ�`e8�1ְL��k�M�LǕ��������V��j�y��f�����a��3MN	`fOS~^����O��:��;���UDp�+�?p��MX�����h%����V�5S}�)�z&ٶx��\�{͛�=)U�xɋ���3�i8���ewў��̳	ǏI�L��3�3��L����:N���<��f�u�^���]u���gL���2�j�pZlW�����K�Os�5h-4̪oW�urKFG<����	K5�3i�t�x����}3���,��4�5�g��v�aX^�];�WY�t�4����/T�6�:�Ӷ�z��i���nү��k �X�C�ٮ���Nǌ4��20��9���Töx����,�w�ΐㄮ�/�5i���/soiX�/87�^����S�Ɵ�v�c�w���z1AzM��IY�����e:�&XTۨ�4^�s�s�v�3]Sn�'�������0e;x�zk�zNus<N"�d�8��gZ�Vi*C���'���v�O+'�G���2�7�0�H)×��W�o}o_g�:����!_�>�?��u��n62�%[ܼ\��}z�Z����/�I�D�Va���M�\\o1e��<f�HԳDb�e
��@p��鬝��g��H��3�[���Ӝ�-܁�u�����f�����`���Y���K��6���~��N{�F
[)���G�k|V-�<��x����X��g�r�B���3q�璽W�q�X�6^Ƕ�sO;��e6kU�}}#L0n�OT�7;l��0LCnKV��}-�!F��}�?�n�n�,C���L�ׂ�u*�J���+(b̙1,�����u�>ƶVOk�6�:˨�i�S��"6詧9K.r���v@V"����YB\I'�"�
7��9����2�b��s�7\���B����<�:R����$�^Ӈ��?d9י(e���;�(�[ǹ�e�'f$�%]s��M���.TG-44���w�Α#+��6.�����I4p�
\]�
�b�6)1"�������,iO �Y��۷tw���o~�}0���.\V�ն���p�
	h��0-m�[m-�\*VYJTm*��%���lkU@���<ڵ�������y���ҝ��r�<4���9�V�kBk���<|��(���<�d3����4���5 �����L00���Zי�8�x�,�8�`J�h�Xߦ�	��!��$:��q��B�d��oW��d�L�+v�d�L��+����sݱ[���J�b������O/���/p[%`Usy���3c���vfoLXN�0�H,�ה��$����I=2�D��2C���@�[$9�����Xx�OFN�!�HT�L2Ci!��3$;d�7I
��I'�	��Rx�OD��$<3���;�Ho�Hq!,)�I0�OD���s��[����$4�^�I2�,	�XC�$�ﾵ �'���j��L=I�Iy�u�M!��B ��n�!�!�$�<d:��w��a=z0�$i$�_7�=4�������t�Ol�)������7�$�.�������'˦����~M�%�S�F�|��E�#���+�X��V�۰�Z^_u�_�6
�̓xq��>SC�>����Wմj��k��ZX�܃lL���5�n���Z P�Ƿzy���.\[��1�����g�@k���9G�tWgxӫ��l�oml��7��B�����י����{ � q���q���,���ҡ˳1B��E��ˬ��b�J���W`�-�_'���M�ΗhD��vȽ���p^�<��h=�~�H��c�};0�]t�>wi��F�佑�ˊl8�n��*3�n	l{�%���xU�;���o;;���&p�H�i�<K5݃�~����3�����43�e9QL�ą���Ȍ����`R�@Phe��EI[C�����������o]s!�L|j��h9��g�!�=v����Fdv�п���cM;���N�/��xVgv,�#<�k *q� �c�0����6�#�G9Q�B��ĝy-"�*��h�^�e��_<�Vg{�~r1��GGv�p�<[��*�^�Ą>�:O�����4�LW2�+�ֻЕd���jpFh%�n��\�E-`w<�"���A�!������eY��^2���5��4v��0gv�/ɉX�{������P0u�}Xw_���Vͤ^v�0\}���z�z��p�,�ƛ�jݯG�$������6#H�܎�q�4[��x[��Kư.��ǅn��ϧ'�Л\�]b\���ס~�o�?�¬v��+3|q���L|�k�Ch�rݭ����dO <�+����4V��e�o4�r�6 ��
��g�[���X\f�u�ñ��+/Y�n�y��+<w�Ch����%�+����2�!
gF�������4�Y0��Q��Vɽ����d�{�����G�w)\��P0�7ܲ��k�^��|�q3��+aǒ�9s��Q��;�Ŝ�P���J햫s�8�N�yvXD�[ҴN⺄�Q6�$=r[u}ժKtZˌ�O�A��7O+�Μ���l�E�mkUe��m��b[kR�YP�ee���+m��YK[V�U��6�+X���NR�B�ʵ�-�i,kX� ��&�4�
�(�oWw��������p�2�����V���j_����;U�s�Ĕ�\D:3�W9�������^�9��O�a^�{�Wuws�L�,C��^E�����^�{�&�����U��`R 2{���EWJ�|�&�3�<5��{���͓9��tEʭ�K)Mt5w>D����"�P�A�;��lT��i��,·p�q43�S�pàX��*�ŊI��zR�n���6o� kY�f��B��]m�z�[�z��(G��,N�QvO;�(�د���m�f3�NC�`e<	�85�u�o���7c�7|��YQse�-��v֠J۩��7�?��ȇ�i�?~u��ߣ�i>]ͣ������:���zpk�#�vTR�~��Q^k{ُ�΋�{�<g���ᰋGE�#E�t�l��	���;����aC�,�#�=B��Ttߖ1汥��p�{�ϧ����v{��.�Y�:BK%�#^��%��r��:���_2�<����i���\Yv�v�7�)z�R��$%5�0\'�윷o�{�x��2�n��������&b4<ל�����C"�=k��Y���׫@�=G�z��.R��44��,���
]jlt:j���`����F*��`Q�\�!,_�d#C�<+/�گi?X��x0в�2fo�4;�g�,�|U;T�ܿ_,�0�'�t3s��wy��N��n�ocԷ���F���E�����e��|���kv��].���cc��2.��{Q���QZ�����l�t@�e�d7�R�3�Uz�t�A����+Iy���!dT��R^ݵXn����ֱ\��d[#O�_R]S�P�W�׽�>J�~�)jx�˔���V���-t�]uHi�(w������1v�Wcr��x�wV;ԳƹY�.VZ��������Ws&r�{^�E��oa��������}��s�'o��H^6���������ϱ��������gSѬ��P�ۣk�����-�����d|2���V��je�e��R����9b�#0��eR�h�ĨY@E��o���f���#��Y��Y�������>��'
N����r�1SZ8�y�N�F�lv���Yo!����K"�f��V�p�e£ȃ&'Y�7WX�&l�5�.��_Ɩ; Dt�AjM�A�^2�t�1�8��V5tk�n����z��&1+�qάNL↘����:�L�:8�3�y꣊��GrK�Wm�K�Kw�f�7�F_L|]����Ւ�8z�Ū�.<Y�3�'�8�_ƭ��C������lڊ�QDEKh���s�9߇�}�9����'6��KL�?²�i�L�p�z�5A���Ǻ^~]�)�Y'�$��#�o��E���b>�Z�6�Vz!z����c��Փ���_�_�s~���~��E��{M�>R��`# �V���3j��}���7�:��~��o��j�A�tN�xʰ�����g/$s�v�I���s0��}4ѱE�<�Z5z�E�W����X�[cX�t�>u>��^�Z������o3b˕�)���H��AUH�����hG��]�h��	�����p�v_�p�\O��G����"���o�79e<F�'����	{�oS��9qM��?}_UQ{}��$����S�.Jby2�ϧ92����Ξ�R�h�x�7<y�6�_������m��6ę���w��V�/o[���yR��ҏRɄ��ԙ�n����������,�{?M�VS�z�`F����G��P{��c��{n����G�n&�a|�n�3<�FJN�a��~!�����}�==�קiv�opCXj�~=�{̔���g~���Yڭfs��н�֭�:�z���l��7a؛���n"I�|�����u�c�Ri6�T<�bK�ގ�ͼ���r�L6�>*g詷b-� �d���_}_Un��Ғ��3�&7X��԰�]Ԇ�׌L/E[���=z��_B�J8�9lk+t��v:�Y�W�h/{"��cᄼ�Jgg�Ees5��݀�y[���9�����8�����K>��f�5���r��g�;sЮ��"�˰4���M���{U�6_o2��6� ����d>�^;�L/:>�o}c�q�'�[�Xvu#s5�]VBK�A$�(�Ne���}�%�~������ֺ�����o^�Ƨ���P:/'=���1/ʌ;��������Ն��ot��ו
��q�9�6z�k���]a5�=U;��`R�@h}�o7����x������^:`ƨ�O�Y�n0�y�kw��1]s�޷�n�.�V�Jp��B4�^'/4N3�A����,l9�*��O૷߱��ر
��BUL�=���%�y|�8ꊮ@oW)O(�����s����X�b�`�f�Պ��t"�\䀩����
���t���<U���Wl!���a�Sk���;�Wt�2����B+�&��
�����[���<5)��*�~M��祻r�5^�{6���ˤqrQ����mX4t�2VX,��c���gaj+��p̅Gv�6^'$j��͔�׹�3�q̂��q*<�:"v���Bs���'뾏G!��[�L
̣S}�w�^�y�0���[JmKAj�mE��QR"
������j#�P`�F��iR�Jʶ�
[kh֕�Dh�6�[mV1D�B����q����Ċ}--?/3y�V�?�կ���}ʢb<7�a)f;	���r����1�8pp{�ƾ�g�[ڜ��n�xPtwP]v�Y��{��S>�Z���7Z�ۭ�7%�*rl-��9I'�W������{��@/�Y�,�y��n�5<b]����Σ�v�B��k��=�J{����j���`>�뼊�A����XuV����A5�豻z�sf@@|��y����f�C޴�J|{�������oE�}f�ׁ]Cuy:���kw2m�S-��ܫJ��O��B���,[T�K��u�g7���u&
}74�E$���FK������Ş?��+����Ɏ��8�ܫƳ�����x���^b����۹	/�p8��"Ud�iwNed��tGvxֶoh@�L_����]M�=`�p_Z16��`Rp����%�_(瞉X�P�Vs����9e���\)�G���]�Hq��=�o��2^���iF���g�Ȳ�^Oy�� ~�+�/y�'p���8�R	5���r~������w�^K�6�WCF�`��Lm$�ZyG
��v�������%997խN۴��{��EF��X��n<.�Cr�f��#��ܥ�͜#���9 I�R`� �i���f�S[�����cV3��x����Xal�v�On�e�ӔX��]��f�r�ܴ|S���]��{�x�|�A�ӂ-��Җ�C̙X=S�3�Y�L��[B�L�nH ��{��2Y�9s5T���H��D�����N�V�;{��v�$��>�u�v�qy����n�����K0d{�����Q���\3Q�'<M�����7x+�(�n�<��C�N8
tda������-_�h�u�������#�o�*�1��t���߳!�o�e�|PS�~��Ȣ�T���?(�-%8���]mׇ�E��j��+;�cԟ�d�!�-
����SpȀ�a�}�y����mX��^3":TTq0�j:Ey-ғ��7�����\�����7�ªkW�ۃϝ"]춢��4�r\s}��>D�����~������0�CG=׊q�h{�Ⴗf�,z7�*R�*"Gq��@w$�Ě�V���k��>��f1�� enL�G�� #QپWLi}/W�Վu𛻠��[�n�47n�����{�V�S�mb
K�,�d�+1(wYSt����("�D�oh p@����|�XjS���a 
ޭW�MU�D-�)+,���v�A�YhM/H1u!H<P�Ny�L�&̭xxi��rL�e�B�X�'v%X�&d���8��)�'�N�]�N���N͋k|���"��ZQ`�le�-�Ҡ���VR҂,-�QE�DE-)m+"��mR6�*j�EEm�-iUR��e�����U��KZ2�j�D-��ib4ZԢ���DZ�Q�hֶգh�U*�F�Ym���meV�kl.7����k5H��|����j�r�}yf)�9z��LwZ�|����7y����'wS�c^��'DWi��� k�Y�9�흑���ʲ֨(��?Z����KN��{���
=�F��x��_�8�AI4UЮ�-7�3wO�����|�02������[�Yf��Ĺ_�V�7�Ih�#.�EY�m�OE�Լ�`�R�^�++փ�D��L�b��G���ю��|�Q��r��<�3LҷIX���ew�t�U���2�e_��c���gCja�������4�9�D�ם��Q����Xʗѝ]�c�$9���mB�aa��n��+ȫ*�/�=`L���qQ�r]�^�J�\�
-���74���̔��_ܦ���{ѣ���tH@���(gv.
��ƻ�5��u��(m9����dC���fe�޲�N�5�`p���in�~g�Fw���״c�XfOVo �pH�3+n�>�z�Y<���G����7�]ն�����,$��͞�6sWLo2'�e�/"yԃ|�uߞ�%��~n���g���[~����Q����wGhιn����.��z��~qdX�JW��1~v~|g��\e�k�<�9�˴S�w�#�ع�;�����A����i��`���0��T�4{wǳ���&]��V�
�R���?�O5P�s��D�O���mS����x���K�f�J�?9�����]Л���4Vd��C59�� /<����2����G�N&f��G�ؓl�A+��ѧ^ m��Cռ��Ok��w�r���n�,���7�����T��%������X�̼P$"�[z �'N�ز@��3"����[�4���ҩ��7���]�L1l�/(8��:Lr��=����;�7=�~��s6|}���~���jh*u�͹�磌����?� O˔1�ʲj#*춢��ӭ�Y	��5�0�/z��yz��)`;c\�YEqUն.u�Ns��A���l4M�'�ߺC�Op�Κ߷֙؇̒Ջc��@�����������c�/ڑ ��g�y��^�˞���/���"pɦ���~�c-ބ�����7rkp)�����mh�j�K>'���M��Ǡ�����g0RTک���6C�/U��/�� �����6�GPu��{��>��m�	� �{�Sb�i��k`z;qꖰ)�P L�rZM2Ï7�83$��b��Y/�ќ�,�ҋ�SU�"���|�!ƙ�#�OJ;5���s��Cグ�ɖ��*��5�/y�q��c��K[�l]��ZV��_�G��=�Ǩ�l*-����·\;�Ͱ�9"��51.h�k�f���w^�"lήa���ɒks�	�*h�/uF^��b����)Q�ض�_\�:菉"� �h[iV����iDD�Ա-mj5h��m����ck���[Q�,���kkj��Ѷ��aYK���FР��m�������h"ڥ���b�lQUjZ������Em(^�B�X.7�VB:�s4ـ�7��+u+�.�����o��y�7�U��.[��ޢ]{��PS�&7ך�d�{}���OxV,�hމΞ���@7�����u[��37�!	��+�� �#�uݍ��ׅ>$6�fl�`�S��i�����?�:��瞨U�?�_Cź^�������q�G|��t�H�Fd�=U��Ǚ�b���՗�kmx�;�sכf������bӓ9�R2(�RS/��g��Z�� ��쌽c��T�2r�L��'�����o�=ߘ�»��w[:��v���V<�3���{�R��̛�R�2�f�eW:~�R��1�*�Sk;��� ^㭹]Wh���+pE�bgP��*��I��[�9?QC��Z�{7N����oPY z��1Coy�]��J��n@w����3FqQ�
�%�WD��#!8��	(��]�-{:쇭5�h:�6�Zk%�k��U���҂������.< ��F�V|��}�u��u��G_n71/�J�"7�6U��;�M�24�6z)��X�����/��1gyg�=y>�s�1�%��5xi���^���듒lW�$�[�RNp(�ݑ��<�U3Ï��e�d��Տ3�ۀ�'�9ޜ����'9:#:���S�}i7�-�V����iM�!�}-jEV����j��_����~�:�Y���v�g�D��U�h�Ԓݩ.�'�v.��a�<��o=��}.�!�����2"^��z� ��0N=���o3�/|ֻ��7�(���[�ܰ�۳���x�����κ������޼�|���V��g��!��T�"9q��C6�ڕ�3_�*��G��������&���tir?�����^��nɖ<�O'�m��F�_vU��.芈ܣ�N�2%瞑y<w�-�^`������,��wT�܂Ne.��q�@\�ɽ�Ǖ�Ǹ��d�eԇ�3[/"��n�p������:�G�$�G���}өb'E���6�b�~y�^�����b���5�(z�z�ʵf����P�e�%��2-��p�h���k�Ƴo3[ȗjE��c���+h�R֙�7磭��t�$��Յ�Qx�D����̉�ɢ+�KFR���/����K�{|����S�(�77��f��btuy��7x��Y�U@h�r��eq�bG����J�����0]5�I�Foh�� ڕ//��	�hi��j���K�/�����L�rx(sT�pM��k#������]7.ja����\6�_+On� 'Iy�m���I��\����_meK9�"N��I:�9�Q%�#��:zqj:LIۧz�n)yGvi3z�����$)q�g(�����r�(Нc\s!�޲P����(N�֒*�uq2��S��YP��EUKq�0\&-G
ؕm��p҉jUcF�B�*-�p����c-
ʖҔcjV�Ⲗ�h�[mkq�8��QT�1�mZ�������b፸W��Z%2�H�QT�
$�����y��z��5s2H{������NX������}�<���u����]5B���%�xđ0h[��IlD[���󧽦�8���8牰A}���1����ui�#[�1RB�)F@ڄ�r��{m�e�|!l�|�9k��92�1�Yˊ�	����L�^'"5cҹ�<�z�g� v�,)e�3n�ͣ�/1g��&��u�;�5������W���JB�p���;��ue��,�`����V�6��.k��|Nx͌�����܈�e�����k%�Ã���i�1ڌ�~&u��`������e��Y`������w���Ha���k����N)��9g�ζS�M�Uyf�vT��b�y�Fy�6�/�s]}r�yVs;۔D���>�@^�G��`��]7��hqݯ����N�Ϊ�����F\S`i�p/�����1�<��n�'��|0*�-���w)z&ic�U�q��jp����7_,�0�J�����Ca˯a���ӻ�,xg۽]�\\nҾ�iH\�b�:f�\K|��ك�K�#[.�l��>�
 v#yP�X�>��w]���c_��w��W#ӷ:A�˝��h�FFO�=X/�5�����b�Z���{��/=���FB��#.2t��Y��զTYJ�3�7�(z��hŶ"}-�e��I9��B�}u~֞jf�)���Tqx�|��b�*rn��X� 2P��ߑ�L�Hcd�	f������gv�N�P��7n4q2rnɖ�,s����qL{ɒ����6��|����~�ʝ+v��;�;b��=�sգ<�=6��{����!��6�';$��H^{)D�T���ӥ�~�h�+۬��+�j�H�o��bw�*��3d�vp�U�n*y�`��S`4�H�^ve{C������L��ϻf�F�R��7��1$�&�F���9:�1�x�w��ïf�5%�3t]5u�oV�qU��|	}g�k}���=go�.W[��7Q���}���h�'k� ]������?�۝y�R��oK���4��G�B�·��@�<s��B�z\�ϲ�68S�sc;��0,��Ե�T%R�_P//��$iCr�] �7���N��n�փ�i��̕�u�3�oe^���i�䝜z�t�'�Z2i�����q�hb5Þv��ԣ��r3jff�S�s�s�JL�� deG�A����ӕv6ᕽ�ʾww���zau��<\�S�n>x�z����e0���.��;7���2=�>j�5Qm���qh"��eDq��0V���ThZ(�m�i�S�iKb6�ʕ[Z[qp�c6����V�e�ѪW3	emj�bڣ�[j��-�a�T�É��,G	�����ݛ=͡�HI�5i�k'�>�[��pʵ�Y�ؼ�J�!�+|�����g�,�fj�,��ʞ�J��]l{�ɣ��'�,�z3ˌ�۫��T��{ܽ���}���Z򻞒藦��N����i|��!/˰���H��o��\�ydkS�]%�Y���hU�ߦ�{V$����g>�3^��i��b>��_�<-;断�qX�$A��i�"�����M������`#]�;�/�E�n׳=��3�6�Ki�)~�m�4@w�����k�0{jZQ�4�|��x-�M!�Š��ήS~:�T�@̏6H��R�����Yz�XN��,��i�^Y��R�p��iղ<��C[g������[�7@��m�8]V|{:E�h�䶬dz��r�f�L���j�eBQ�jE$���FK����x�J7�5�)�hy�鵜�iO�ˡ#	V.K�c�m*w~���qFS�]�C�6�(w3��m<	�) .��h��}·lT�����Vw\��W!��@��g}��K7���|=�6y��:��E���_^YA��/�Z:{ב��W�;���P����Us�ϭev�7;�_$��{jR�s1�Ǖ䎙I8$�R��	ɀ�\~!i���N:�����C�we>�[�`k�o�s^UR�t��ߋ��w��{,K8ոpXqn�ʿ� �V"a���y�g;HU��֔�}/3��4�0Z`���fCu�<�*�ڮ��?>1�����x��)��8N��Qk���V��Y�g7��e� 8)�U����y�@���ۭ�:mme��/�rȂ�}�A3RD\-F������*#�K�̘�U�6�=����˿�V5�/K^W�Yuw.K�HC��j����[�,����>��;>]w������k�Gy>�UN8
�B�t̋���S�JSC=��"�%t��(����fy���F�o�d�M��~Ȉ���h�����®��!n�gu����{�v��\N���7��7�3y�O�>4�TUI���	Aŧ�����Xw H���0Fl=?(`�d,��������{L��I���O�.XgT2��8Іq� $�)�SV&�T,�������p���=c3�_e�5B�}l?�=�@��ċ�x��w����߷^���� �xO@�?B����F��>!�J!��\��l11�`�R���-������k�!�����!��?g���铻��D��H@��`�� !!�?� ,,�>P�����Cԡ�?��l'�C�ԧ���u�!�}�O�h>���4�XB@��=�������0|��]H`:�2$���}hdHr`%7�_xx@�$�~Қ0���[��ܑ{�ߘ=�VN__��`>��n\#�	?�E�$	�����]���a�s���5 H�䘒N�ʩ��4�8������2C�n�П�d�?PB@��I��VJ|&���	���{M{{����B��w�gd�{�����l��	��� �p�4~A���O����|��OgȌ�B@���K#<1������!��|����fB��Oho�L�B���_��}��o�>��'�	�C�ހ�C���}��|���q�H�����=���!���=�'GA��0" (�p}�-�϶�$L��$?�~� �v���|�b� g����I:��:5
�@���H	���aX ��10>�H��:d^IBB��E�D�	!�>!�4>�2�@a�V�� ~ ���p�I7�g�&ZC��5�'S ��u��! Hw)O���Y�	�� H9�>D��	$C�>�X�~��z�������?Ȟ�������	�����i�>tC�>��?�|��c��	�������C?���$	��g�^���� ��!iH����A�R�!d�t���`��� ~�v���o�������!�}���6Q@�'���#&a�h}��@����>���=P�p�d<��|���q�!�vxg�>�Ϩ=��$	}A�n�C�8e�w40�O��D��a���������(s���th�`���!�}�=�D	 H�FI��O���$<BC�9�~g�w�W�	 H}R|��O|l�P�>_*M���$�05�}���c7!��A}PO�)!��R��96rE8P��� �