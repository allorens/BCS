BZh91AY&SY{9���߀`p���"� ����bC�|   |�_Fل 	(P �d6�U Y +kf�Z�A"�i��i�T+M�l5Zʊh3c U ��(U4Ud2��Z�E���R��;,��P��h�%�V�Kf�
ղ&����jYZ�B�f�Ѩ�MZ���15mkV#,PR��U4K!m�e���cjhj�w���3SK�*�F����#I�6e��TkEi�Sel��,�����e³Z6Ԫ��,Ԗ�ʵTɖ�Jf�5meb��M9��Uff�5-O   ڟ{�;��Y�QU��:>��{� ���mZ2ـ֥UTl��{m�k���{&��[9�T((�V�65�:yoVM�R����A�k56ʴ��  �����oo-�;=:wtOu.ꤩRPp�骥M�[�/z�J*Z���)�ԥ&�{��^�m�^�M���Q^������Ik*�����i�j	kI�xժ����m�ږZ�L��f�|  �����P�nSq�ʩm������kJ�ʕ�=ީ'ON�^��>�h)J�>c���j_mJ��[�y��)[�>����T�{�O�Є��������>T �ԣ�=(Z�J�ڒѢB��J>  n�}
��o}�]��RkO>�㞓��f)+��y��{��xy����m�)F��l"%M�V�WlK�׸���F��=�އ��'�3���wn���*��h֚֫66���P��  n�>��W�QM�Oz�]a@{�eީI{j�����/M]��g�d��Pv=:���ޕ[�ΜF��w��ңZn���^�����^��������O]��wV�lx�$5��l�Z�[L�V�[�  ��Kmi}ޭ{�kn�Q��5-���u���A^w=�n��NݷI�{ަ���3��[�)R))�)�r�[eJ������R�k�<�%T�M׳C6���4�HJ�X���o�  Ͼ݇R��>�t�^���u�v�JUJ�����͍):ەn�*]iv�Ə:U)R��sҩKm��ݯ;F�Ƹ�w=iJ�W��
��[��3	��I��+�  ��=|�5�뗭�vz�z5wy�=kn�{��kʨ뮻D���wy/^ĠR�\T���=Ǣ��q�e����cl�JMV�k2��  ����AJ�I�N�p���x��d�5�Gz���W����p�C�z�:��۞��ʠY�y�kF��ҵZ�[m5UV��-��   ;���Q���ÕBޓ���'��xz�Ux�=w`=pwJPP�훇�a	�^�<%W���=J�ކ/j-[>    PB�"m ʒ��A� hh44i��)�)J*DG�4  "����P �#  ���J�  L  i������A��M�#b=C��I �T$i�'�4b�h����W��������A�}ޮ�ݿ�k#)��+ƚ�4�����Y�<  {�T��>� {��ڪ���u�����kUV���+_���������U[l��8�^V����eΛk��ڭkm��_������9m��Z���L�|ͫ햷��k���͵�m���sV�*��[ܭ��k핯sZ�6�sm�kܭ{�W�Z�+^��ֽ���5�r��[�[��^�kܭ{�׹Z�+or��V�9�ܬ�kܭ{�׹�{��r��+^�kܭ{�~r��Z�{��sV�5�sZ�+^��m��k��{��sU�6�sU�Z�ͫ�ڽͫܭ{���{��sj�6���{��sU�Z��W�U�m^�W�=�kܶ�~r�[�Z��-�o�mjߜ�U_������o�kjߌ�սʶ���սʭo�jս�j������U^f֯r���+Z��j��Z��6�orխ�[mo�jսͭ[��m�6�{�j��Uor�[��k{�շ��[{�km�m�W�-W�m���j���[ܭ[{�ګܭm�ʵ���m��j��kZ�5V��ֶ�6����U{���ܪ�{�V�sZ����mU�Z���mm�V�^���-�_|ڽ�׹�f׹j�6�sU�Z�ͫܵ{��sU��W�j�;5^�k��{��r��V���[^���ͷ��V��k�ڽͫܭ{�[ܶ�͵�m�w�u��kn�k�ֽ�kܶ��׾>���ק��|T�`��8W�S���5���ޚ&YS��YX�&Pv۱E�rd�����j^X�X�Cb[�T�7�����-o��`գ���i��	���K�	�۽wr�F�7Ö���5��&Ɛ�Ҳ�fݥ#��Ѣ�mO�ѱ=+~e7����A����/��@���}E��K ��N�A����@.�X�k�nH�5����HS����He�kpkzR!��Y�k��A�x���Cw��6��˖�⌠R.�Rd2T��wł� �G��U�wY�c�TuZ�w.%���հ�cL�V7i��ʱ�6�ڃ5� )�[cr�Z1J���l��ݢ�6k0�nL:�I;ank$n�B�W����[�e�Qc�x�0����kyf�Z��n�h��Y:�(F�cVE/;m����gnɼ�w-]��4]�2��ܭeT�:1��*-j���,�ң�6!�%���xȊ���dRQb�2˦i=���,z��Q:7�Rj�`:��ٹ>%
��ͽ�������Dٸ�u�Wg�*
Aݣpf��X�L!K�HsM�@�;b�v����v�5����km��֎E�ҍ,��&��4����7�P^�kP��k! 7��>�u�P��E��u[Y1B��33.B�10Z�������Zh�#r�X�ĩ �+�d�Mʽe�p�E(l�V���C���+�E�Š�HSN�&U�dاb��B�A�y��@�L�r��cR� n�`���%ԷWڼ���
�^li&�-�
��4��d&�^&��,@Ŷ��]�C��]��4���N�Da�-�۫�j���ƷV*h{w��Ln���5���e��M<̿��(I��awo]hܩo.����nJ�t$70�י#r�{w4���ORr]�&Id��A��ъ��.��]k�h��2Q%�V���գ��&��
�
Qa���W��%"
p�kh�[H칔�xbQ��S6"8*c�[6�,:�sZ��}0��3��z`�J�I�	fˁұ<0�[�dz�֛�x��8ٷH���s����*j�ei����E�4������a{���$�V�']&饸����۔� #H�2�:ҁ�U%,��%cb��̟��z����TN�Lu4�������-��Vm��ͷ�2�V^��	�0T�D`t�*ǲ�ݧh-�|޸�UdR|�h��;
�6&���c��w6��[x���W��īb�q~�"��UE1DIA=͒0�E�&-���^��wl�W��ơ�d3-�ƻ��[�m�J�Ρ���|���ky�'��<ᴅi8�ڳ@�]-<E2h�EEmS�����A�͋b�`��/ي�����ף	%�ua�QJGz(U7RY[q��F��n�lq�m庆�M�a���L������J�����)�#vY�Q̵l�x:�N�Ē�.��7���w$�:���\���ӈO���j�ӈK��,���i;��	��Z7%�%X"��w+*=%��ѷ���V��ڴD��*{6�c#e]���m�g5K�5�$�a�*�;a����[X��!3�#���D�Y���Ia*m�3� ���0�whP��bP�u��ʺ۫�	�ü:)Ś���ێX��"��m����.]�釷�P���E܃.'F�ܖ6=�1R��E���0����ޔ"D��rP�e��An�\.ռ��-'x���u�oq����-5*������ZֵY�B��Q��X��tD���I��Sf^���l���e��hT�')� �az��:��R��Yf=2x7R;��5�oW[�%[C�//r]�Aԗ�9Xl�X�b��橗�h709��df�7/��v��m1$�u��*�q�y���JF-���%�Hm��f�kmҦ��)64�K%��o�Rذ�n�;Oq�;��z���+p\sh�ס���P��ѷ�1ͨA�0m��+�wLE�U�T�2F��%q����O(��#Z�X4���7ݹ�76dU맮�kb�	Q��,�L���J�FA�j9y�������i��UyF��n�7�C�� &M�ӷD�ú6 cM �W���HN$Nw�L�4a��`�(�w"�2]wjkE�x[X�%+�ƝK3��QUkK�3Q�M�/Yv+^P����8�)͊�[4�J���oV=[z�RvhBN�����٬C
��m!��Z3��cvFdիN������ՂWQ/�`���sH�d'y�t:q�Ҡ�6�@H��jgs�k��{YMea��!m��;�s��4m�P��rncV���ZH����Q�N(#ƕ�+w�q`і�D�XX �Q�����46�5N�\�f�5���Z�.���p4tb�{j�.��u��;t�m=[�c���f�A̦��e�@�0���t��<��2��
� �w�C�$��+su�����eY�aڐ�:�����6%;+�ɧti�M�a'[n�ਤ����dӐM��lkeE*� �`�.�B��n��南h�P'0<�Ld��F�B��d��Oj`ڐ��7�ӡKڀЃ0Gv�&֡��;Gm�3?�uSj��'p˥7�wctm+U�R�sy�m��_u4)Y���!r�FcsZv�1s˥]���>;�[2[x�5i���V*�^�f�ӼXFࠊ���ְM ڬl�����ߝ�>ZӸ��^`Bn�.��z�����X�e5�k�mß_ieeֳ�C�В�GyW�^�l�v��z�'�ε�|8�|i����Zw²��e[�Uvڑ�Th��\w��2ȫj��(F�o�� �l��^�N��p�W&b�����K7Hy*���S�r�soNP�m뭛�Y�	ؚ��{�<le��"gv��nrά���Vë�X����(�Bm�ܵX��͗5�|ѹ��U����H)�	�4Ue�Tl+c�Q{/e��J﷦T���k�Tl�"p�X,%-jG7�f=��F�+�hR �[�5��[E�J[��J,��
f��R�ה/%�E�N=�Q�c��J �	޼*���
�Q,�
����@�1����9vB�ԮL�"���K�j�s
�d:��ޥHi��g���YO.2K�L(9�q��lШ��h�װ��T��'E�гbʃ�,��M�T%��}4�+.�Y1�B�V:x�]=�&;ژv����1Vk�(�i:�+�ZQ��l^���(�lؤ(j���+v��KI�Ϯ�X��Zp�UɌ,�g�M�Vز�kx�3�Ԝٙ)�f;;&�mLVf����8��l;��07-$�X������m V���v�N���e<��#M��"e��G.+n�c3i�7�x���MY(I���2�FoH�dU��R�Pc
u�-���(ao*���m�rD썚�[�ҭ��A�cܨ����l�^X�eSʘL�c8�Y7gS֙�b��;��ͼ��z�ᬐ�lbVH�ǒ6�{�5�M�۩
y{�l���IVsC�76դ�;�%H[��5(Ti]᭡M���9�e[Z�)mř]wWX�v�a��yP��K��n��Y�	�9EҲ�L�1�b]H�i��'�n�������@f��7�Q̭S�x���D�M�JZt��6��{(dͥr��UF�|\�-�#r'Y���6F ki��U�5X�Z�V9D��r+���[%X�r������Xy���xa�VQ��`�	{��:=6��*�o�P�nwl�i��x)��|�2��4^���X�{��ͬ�4O�+�oq܈c���N��;�f-�k�T���GbP\���/@�Q�˷(ƣX7���6�;M� �e��6��F�h,vr���l�X�*TInm����AǦ4�	��m��a�6�y6�Y�,��śY��8%k�M�L���!�n���j�
�8���6��S]�	h0��(g&�0+g��q��)��\�g ���؞�[��P��Մ�$f�e�̧�C,8w^d���M�'�{h��������r���\m;y�������*Ѯ�R�=r�m[���L�;�5��T�Vo�K�+HૠQ�,�.�:V6�p�x� ����[�����'��A��¤7 :Ֆ�Cj�wZn��,�( 7[:P6��G6=֑/onZyur�FUi��̺a�������BKL�d�������i�KQ�'v��a��":�j��:E���
$��Y��JS��Cɔ3t�ܡF��n�	�5����0���Vѥg�<Z4EA�D,4�D[� ��솨��:9cn�W4��1�g�9�E��/)K�m����fEK(Jw���(�"2ڠ�X2�U��Ñ��n	0�hݚ����
��CFp��K���̹3RT�-�a�R�Z[���h%�"1���nc��~���Z��l��&�e�4-�/v=w���7j�72�a�%�W��2�Jt ���0���<I҄=	��p`oѭ� dX��S͎�^Qt%�h�ŭ�7	-�1a���|M��wNC��;,൚-���ܧZ+L�3&PL�F���ډ;�@�W���v]�b��H�����f�lM��*=)�فԽ�b�e�.�Çn,��d���0^@��f�&������ω�יkD���-#72=J?�)B� t 	�Q�"jc��e�<���~�mXCY����XE��1���⼫D��H;�tQ%�F"6�d��Ae]�Fi��Ûzˡ��v:�
�1x_n�,om�����&]�$fb�eёb;a;��K^�eK��f^�ۥe��&8�;JQ�]����kSQ^�-B�rJ&�����4��=u�e��gBшc�2�ӎ�3�f*r�ئ�-�p�&�f�l�SN�z"N
W�a�Q�tks3/.i{�M~4�蘷3�Lb*t�m��7#�|>�j��r����/߰Z�m��	�7�՘Vի��������1õ-���i�QVXc���C7o0\��I�ȝc�]��&��,k�Zㅋ�ͺa vh�U�E�,��Ѵ�enV�ed�95�T�#$�����k3v�<u0��n����M�xt�$N"�P����7�=,
[�%�6��S(\ �H��Ϳ���U+{�X�͆[:�э6@��T2�oA���e��O-��;��,��X�Dm�3X�؋�"�l�v�ޗ6��U��g&�J��Ta���44�-���2��6��¶!����[:[;%!.�u��-BLݍ�T�h���XI�u�Fd������iN�H��l��Zhz��C�_���EqH�b�n�4,�CuON��	B<���w+wmU�&�zH��b�;��TCN��n��n�Z�v�
X��f=,��w]T�N����-f�b�ܶ�69 9���Z�Q� �N���azn���mi���%^CLq��Z\ѡ�`��XS�;�A�U����*�#�׻�YmҬl����gove�i��6��zaE�ބ�VYC�MR�`��z�?��i*�f*�hfT��{�<���|��9�p�r���j�S��:
�u+�DGv�eշ��]��ry�'�|��.(A�o%��@h2Y{x���3�f�4�.��-��`��z��F�ObX���W�U��Xd��sp����;b+���QaݡJ�۸RZN:h9n��3�1!��j^�)`ōX"�kU�F�V>N�뱠���B������b�Tw#j�5[�w�EÛ{�������Z�Kb�+����0Z�%�EǋsYȷ	m�֡�	�K�FaMGr��td��2I��jf�f�T�Z�elƝ3bk�1�R`EZCH�b�r�5�ļ���V7h�ɇKi�
:�����XY������t��@�ZFj�ҶN�iõ���N�;�2�T�V�3��%�F=ץ�O/%�H��q`��j��cUeXS��(VC%*QP,��I��[�4嫏^K2R$���ύ�`{���C0�q�6a��6��"�%'�h�heL�vŦ�Ɲ�Ff�4B8R�u5����,��%7h��G����1HPg`؆�UQ�^	��lS����%�-��%�(5Oof�ۈ8c��[��%�)H���ymKJ���h�4���l�UB�+����ƓJ1hYۏmV�:sXc)a��*3���$2�n��-��56^^�h ��մ�k� ᢅ7�����a���ߵ���V�*-P�)堝惖��+�d�ݬ[�W�+��2�w���09/Z�2�+�z��i�`n2Ee���m�ysf82��7���/rh��A���ٷch�͈�-`���[}[���g4i�U�(wLv�n�bc"*�[�rX�)�e�u��A�[Z��y���b��l��v �V)L6J��a�lm杖v�i�AK��f���Ӥ�]�(�I�m�
ՆU��l���XɃP��+7kk)M���+˼�Zkc�+2�դ­��^��,��4�L������X��i����|�
�<(1wٓ�p��	���5�B�$$u�K+�gq�45�NՇb���
Žډ~p���1�۴��:18U�U��v�K�)]�Ŭ����*t��(�	l�5	0�A܋q��ܭ�u6��F�۬��kKxq�uw4��>�/\�!��*'�S�f��Z!��h�TX��czj6��6��Y(ԘUB��5%�\��ڂ�'�u���]���&Z��27ĺRG���X�����Ɨo����
�����8S�klӗPO�&#P�� �j�V�b�����y�����3�q�dE�)œK��VSͮ뇰�2Ȳ�f���-�e��0�A�U�b�هm�G�3D݀Q�껢�l�׽�	3&x�>.z�R+����Гٸ�:�S#E�@ˍ�w�I��F�Ի��[�^��e�g���y�<���B��v�g�����$�I$��R.g)D�X�0%��K2���9n�{(U�J3�Z:�x��J5�n�c�;����u����tY{��.s������k7=y(���r����3zS݊���T��L�����5"�e���e&2UvB��gMr�닃�*V�ʇfb�'[�"�<^mZ+�0S���ENt�!���˳�\��{���c���q�7�Ԛ��G*us�s~s�ƀ+%�U�R�(7kA�_^l��d��I�����Q�[.��cmvK�A�D�K�w�⾩����.@�����[����'A"�w�k���kr_VK�Ngi+��h���˲Q���q���uY(�C�m����*m�˩��6e��Y����F��goS�ƭ����К����vZ6s
�n�aע�b��K1�� P�m�x�}t�m!�fe�OOn�*4��-��{^�Q�Ӻ��-�;��gl��p�T�-N�Y�E��k�$�������PR�R�%7Qf�+���w<�#�ި�ӯ���#��!^�m�5"I	zٹ���%��k��e�1W:�٨��(�"z�o:�[�>]�ӡ�d"��|�ܮ�p`��V̡������c�n�WGZg��>jDx�	�B����q�f��`��iS�j�Ú���>U��fDl�F�&d���Ҹ8����z��©u�M���_]��	�\�ؤ����)ί��{/2��)��άua���#m��z/�lt�3x7�o4޷S�|�fa�M�]Y�9'b�\�Ԭ�d�D�U)v�Nא��FU�&���P��ؙ�N^g6��F�m��˜$��eJ��)�vl�ݫ�ˉm�{�E�旲6��
l�L�9f�e��8�N��TU|C{ݙ��-�b��O`ӣ�_�2[h�K&�ot̔�ȵ��xʲ;����}ݽB;;:[�36㼾��V��R�m���V�f �����;�S��O����D2s�� z���掬��M��Ew;������Y+�!��;�&᷹��X�`A��`b�yچZ��Q�,9M�]�yY&D���q�|��an�{�uǛs�^*&�c`���htn��
p�^�r��9�K��1̫qtW�{���KY�����Nz���|) d�g��x�6<游�Y�T��|�ܛ��.���8\uՖ�+5^���q��ى,{�߶�z��o�z���V��G5�rzc��E���®����]c���Ū,�m���[arI�Z�x�̧:��;��ͮ�˰�1��:f�2�̸��Z�Î�c�0�V�tw$	N�)ov&�Rf�RE���|��o:wuϷ^3١�u1��$QZ��,eWR��[{�o����܌¹sNf�:E�+Z��<B���YÓf��|0؏���+dPX��d3u<��%;���rT�_$���l���æqUA��ש=ޱփʢ�k��*�ұ�	�еC1���򬍫��-�|J�-�E�d��6 �X��ut5�a��Y8F���Wd���܅�Wa��ݍ@��1�{��|���s{k�F��ڸ�)b���;L��A�v��&�0U�-�"���}5}Dӈ�2^39�޸S߶c��sJ�|�W�nҾxN�F4*bo2&IJ�q	�V��C��Nňe�ֲ�/n�na.n����ܙy��l.�
��^P�HR�}���{$e�b��_k#�Y��wM�q*��t�*ţm�2!t__v�u֡�o�Yնm+y��9���wG$���h����j�Uml!�]q�D[����V��W�ڝ�L�ã����r�7��GS�8�Pw*H��3&��f\K��[W.�
�`�l��ڒ����ū��Lk��FN�Y�h=�|�ll�soX9u�nku�j]됷Xmg����<f��P8�Kb�/d�E��W׈�Ze�d
3���ӴAj�ګk�X���գ��$���z�=ck'�`V���7�>�m]_�y�&�Q�9>��sub�s]��ٮ�Z�G���b���֥���u�f����'P���hD�7Z�T��c(�G%�iеr�>���JLsvr2���#wyI%��i��gI����mZ1S��-�a�g�g=����X�L����g\S�79�s�����w�-����P��=&G���A�������>��ސ}�MI�;W����QK��ѥv�1΅5�B�c7J
��*�MMֱ(u�;f�뾡��,�)�2�c�OtKZ��
W��l�c�x��Ɋg��_k	�؅(R�E����BĦ]�q�//R����l�2i��-�=���h�a΢��Ը~��/��P��CS<�S^t�f���V`q�{Ք�'Bue�pr�UL�wF�h>��A��*2���[�ѽ'UX�!Pw!I����w$٬=!ᓴԻp(#���Rŷ,����YO��s��u�P��m�}�4;d��f5`fh�cc�`�Sn�v(��wS���;��7�S�m�G��b�vq=��7|��X�Ԥ���v���H�R\�\�c#���G3r���ӲرVc=t������Ω[�ֵ��^��'hn��ۺA��P�=:���ٹc��/U��,X�f��\���6X�Q4�Ll���s�n:7}���R���q���݇���:������%���rVk"&;x��L�͇a��mu{YqQ�̱�Vc�Pۃ-�=p8͞��ʙ�=��Q�vܬϺ��-���X�WIf���z�<t�����X�ѱC�렮�m�q�_	&�Blo!z�M��e�ۍ��6I�	W�h^��rS/�Jx�ב��T�Z#T���%zR�	YK���6j����4�{$����jl�y�k��Ϻ�7n�Qa�tX��b�ؽ�8����]�QM����̙���e���M�ɛI��M�C"��_�[����f�5ʑ��O�Ku�#�]���V)��qÐ�7�]L�E�ٸ-�ʈ�D�-X�ө��6<�K�Zm�O���S�އ۩�WgҊ���A7��P+�u��M��fӯ�ڡ@��fk�i�)���K2+�R�2�ݭ��ws�T��a�W��x�r��}�S��%�L1].7��=��3`�n�W@FM��ZY��d/p�,ch��]f���F�jwP�Q�n�pI�ʙ���JxKLr�7Nv����!°uXR��l�,e��C�5[� <�����U�Vm4l���k�Jȭ������>v���[�A@�o�.JkS�� aKt��,y��we�i��U�P�E�C���ޫ}T&	�*�C���%C���*m�L��x�1O�i�����r��Pm�&�m�C�;
׭"��M��/�&^����dr5�~D\�A�w���hUN�aF �q&��%Bc��7ȻQWM�͛�u�x�5�,9��E��w�6���8V�|�dMR�%�Mcl��b~�1I���11�Z�cYmN� [4�t"� ��̮��+fb�wa7��7�m�����.`_W_N�ܢ�Q	��˨�[����/�d����#2b�o��ݴg0��-7�*��9�3]��9��O)[���&9,��ۮ�ڡ�:��%����Nu��"�e2���}�S���]MB%ڏg������� h���
����.���zx[ܮ��ɓ�{{�eg8C�٭���56ƻ�,_>�"7�Vg��Se�Y��d^ޘ����P�U�����k�;/ǭ`tI�a�e:4�+����V�j�Cv�J}w�� �e�:��&���W�R|L[g �຃�������c$����ݎ2�k�70�E䳢�B��[�[�"�-a@���m����<�����D:�9n���3�3����1沚#3Y�mn}�e�IN}GP�7T�N��[�>��]c����:�X:��)C���1���u����o�39K�;z�4V�IX���L���pǫ-U��㫗�/��t"AHX��V�kŬ��
�㉉�=�'��	2o�r�ׄ���dHbw�<�R��۴N�/el�󯲭n�
	�9QZ��{�R��uoF�YpP���yq���q�s9z�T}M��5s�h��!Ǔ��V�%�@a�yѲZu��Nv��Eی�ƕ.#����ƪ��n��o�-��&2q~�%��L��ϴ��⅍�&[HY8��D�%�\ت�K-B�Q{�!3Ǔ������r�]M�`�x,��L�����\`�ȸ����z�J�k��?p|�
��G2���U"�3�X�נ�N��:�+�w�4=�|��ɾY��8QM�M�5\����.ю
{�*�}W�u��t¨�%�fX�\L$�K%XZ��`���=���hX�om5݀�ל:3'
>��|��έ��k�\��e�RLc���֫ͭ�0���Lyԭ�C\_L�؁�n*2L���j*�t��.czN+@1ZḶSZ��Lٮ�������|r�U��f���U�������Yy�O���E8oT�͗S+F���eNy
EVq����`�]><��4�l|&8�w��/�;}@ZK�|ሶP��E��Cx:���3�{G)pK�����#�̷U�5��qd��"t/,���������E�Oc�Z�:�D��5�)f˗@��姶�R�+�x�:�?><���KU[�
����i������v؃c�Ԝ*�^���v����3S�%�61�ۭ��.�� ���P7�,0v!o�<e��F��\hk)܋�"L�v�1IF�XsgM
��SR|fÕ�Aa2�K�b��Kva��ܼ����ٖ��@
���PJ`��p�37 /H̓Toy�'p�6�\�l��\�9��D���%�A�⸱`*�4��v������Ҏ��v����C¯0ZI���u{�+p�cY�b����A��OO���Oc�g[�Q&��c&��V��َ�rf�d�ե���[�F˾oB(E��d�M�1�aP�f�W�͑�x��;ZI��\ՔM�s���[f�]8�?oP�-V_Ct�[�Y�[{|dᆎ��o%���m�0;��7�P�gL*�vv^G��ͬ�b�~|���<ՙrb�=R���>�c�T�]C�W�n8�>�J�ݗJM��ϝL��mmZ�77��/Q5�Al�X7I�]��q��x'L�85��J�u�R�E���{n�j�;jJ��V:�
F������#����-m�/����y����-������F.Ǹ��V���n/鍥b5B��K2I@Y\��uޫ	��Ԗbj��l�)4��ۄb1�1S�[,Wu���=�h�9)�H�=�j^�DH.�B�͗�T��'�NWՀ�c/m�std�\x�G�O�i�*vr�(�s�8`�Ł����ƅ� ���Dd�2�f��J�6U8�Q��M��TU��ȇq�%!��%���n�8fp��i��q�vSý+��`�N��qlD��XV�t��d=2��!�ʿZC���XZ]�V}�x�WR]���ewɴ���ۅ��a�Ɲ��8�2���q�3��u�u����QI�K'�3��j�=��/m���Qc	 ^P�������7��x�-�\_�z�T��k'Ee�y��P��� �j����I�!pa��s���6��<�oT
HXR]==Ϻom�+wBq1�vۊxl1`�-�)�h���ȓ�ȥ˻��Q&��%۔��K�jj��94��ȭ�x��\���Fз�g��̎��n.�pc�͸,�T�#C�Ti	�O&_Sw���KY�;m����Ϧ�D5g�|�9q�A�vv�#���-�hs;X�G�S�x^��&�$�}E�fн��5��&
o�-�5m���Q�3�=�>�t]Ƀ�[�a��m�K�.I*bU׵��;2�5�����Y��:v��pJGN͘8+� ���]>uyb�Xi9}|.=t��\n���՜	��Iq�
6��ٙ��6�#�<)AO�][�}�i��J`	Zv�P���kK�5+�x��j#v�����X�%i�s82S�Mޚ=�.�^�k���tB��F�JZq�y�;�� U�h��i.����B���7IQ��2L^�x9��Ĵޡ��P4e�Yz�f�n�f�.�����I��E_�U�)��Xys��a���U�jHI2�Z�̙\;Ygw9�4�{&�֮��y���4�+Q��L��\�' �$�3%j��v�»������\��I���&��]�l]e�,s������˹��ۢ�R�X�;;��RMrחeuHF�C�3So�զ�i7]9�2�
,�Kr��lF0vgU��(�Dm��MRl�\$���9NݺvQ�xᝂ|����k��M��8�fX�;�6�n5R�J�G�;w�)�M��F��j��(RYٝƚ��+ܶWs��T
^S�30*��3�����(�:��Z�KvH���8�C�o2�g��+w�/.Bl7E,[k�)}� �jV�ڝx�t�f��y] �r3��tj��)�.c��W0a���2�(���mg;JA{ؚu5���f��.K �"/1J�H�I7��e�Y� �M��՞B�ky��9N��rk�nM�}�p�=%9��ή�C�Ru��7��L�\��3F\}�w'<\���Cr�%��s�I�j�hx�J�]��Ky�:�=�F���k��z�ԣ�w�sz�rLu�v��#��Bށ�@�<:��Gc�H��I'9rI���Iڤ����N�2�mӑ��i�Q��
�h* �~���9}!�Ջ��$п�4@�� �H�����F�#��J�r�)�(�t�B$SX� �T,�ǔ!p"���TD.�e&�F�.S ��\�,�2�I��󍫂	C�^Q��yNQ��)���rF�B���������C���mj�U������~~��Ŷֶ��{j���g�����vG�>���ݾŲ��P���3���P5A�b#7X`v��]f���;^sO����3>;Bn�ܳķ�K���-���!�.���C��2��Z�*�z���!�|r�z���<��ո�!&�VmN*�g^-�a�b�]��q%T-��3��汪��{ύ`ݍ�YX�n�E%��vE3da#�*�̹Z��`t��X��z7R����A��4`6oS���b"�a��S~n�o0n
�&,�[1N[o]ԬQP͠��;)v�{�V�9��k
B,gwj����Kj�_s-�"9v���.��e��oLj�jTl5�j�]��&�5O]��Ⱥ�.��g׼$�]��e�jb�*æ�`�$�Ն���\��GM��ç
��x��6�
����̹f��`��o��a��6��B>�X���-����'
7b��Z\լK�������K1�º��tY�edw����#0a�8��
w>k��%�Z��j���+r�=NP��fU��\�w�λ'GҝsX�QL��.�c�7NZ�e�0�̹}���;4��f�D�ub&�xE�����Gl��s�T������
u��J��v��E�}q�9�Pܼ�³u��pCC
j�Q�Z�T�5n�y���q��.ٍ���e,��D�b��iU��ut�� �lO28��!g �Rž�NV��I�^Ҧ���XԹrMT�Ų�fgiMo%(�d՜��G�XgFڷm���V�O'r�8�>A�U)�"k_G(�����)�H��Z���3;����ngϤ;�m��=ݫp�u�󳐩�l�̘���(l�i����U��Z�����XN"�Y)(�<��H1��� Y�ek�t�Ѯqȭ�ԫ"����
�7}����}h�6Hr���|�<t
��U����C�r��d�G��n�m���J�0�}�wʘw���I�=�k!�2���m�z��4��c1}.f>�����P���S��H8�r������XlS�av!�gf���X�[ኮ,��%;��L�
�ƙ�࡭��++VͬQ�tP�mܚhG�!�&br�۲�һ.����qP���>���ja�6ܤ\�"������ve	��lF��h
y����U�q)1O��l�A;��Ȃ���LE����6�����_[4*����zbÄ�w���N�b���og�V�86���u�DU��N�F����٪��%N��E� q��j�n�;a���v���r�T+��p��WJ�[Sy���%�z���PY���B�+�D�<�IC�72�c�L5���f��Egj')�#DQM��\��wm��K��P�������L�v#u��ruqx����5>D�M-9���H�R�홄�s��d�D��]���".dAI��]����1�t�r�N�6w���e�u+���Z7���ⓓ ���˸v���&;s|NѴkTAf���6M��L
�C�Ui=}�=�]a�)g�3j�,I;6Anx�
 ˏ���_]b61%u�ʬ홹n��������,^t��C$����ڛ�OS9c�ܓ��e��w���⻘�+�g��bGGҳX[q B�D�%�쏁@t���Rׁ�[�tR�lQ��4��M���ފ.��D��9��J�6X�6�u
yƓe�6I|ETx&���9��T��ح�I�v��A��j�F��[6���}�}+0fAo���5a(��8Lx�(�òevglO��8G��vԸ�G�6VV�96pa�:�#U�KX�u�OF}�ό���Е�$����=��חgb�)f[����.�wr3��YJY>D�(�Hĉ�ߔ���6��k{Xq�>Q8�L[���wMi�߅���KH����7��y.�� ������E	������%5��|	J�ǭ�x�zM�3r�QQeoM�4�4[��u�F��t�����a��� �na8��l!n�xg��q��[z4mα۟beR�G� `�dZ����K�V��Τ��f����a,T�p-��8t)оNTG)l�A�d��t�6��Mvg��	cLK;�:)�,6���y6�ج��u7v��!܃|���q�t���)�ʕ�'��S�����!�����z���K���$�����J�K��k�@�ty��2��ު���a����i܁�iC��M�k%:�iXpq�3�|-�E�]Xo���
�����ܥ5���U��K��9����Ϋ�p�茆�!e8#��ky1�����\0J�BT��Y&40T.�s��G���h���WS��1��U����y�7��Ԓ�x��˻��Z��@�9W�nn�JsƷ���a\�OAsV;Ct��p�
4�	p%Cw�yuX�i޲gS:���OU�-�y:�IrM\�nAp:Ms��������꾷-�:�N�iWs�G�c�K�ڮ���7n`h쭭C�|�ʺz���b�V�s\.$d^Vj/&n���f�o7 �����e�l��xC�{��e��t�>Ta/iv"n.$�f��:�\k�!X��>ﻄ����.��42v3:����W\�,<.��T��M�ώT�}�Y�Sk��%.���]"�L�`�$7H�n�޾�l�s�h�Š�\;��_p����em�u9m6����.nԧa[���,3���+���DU�fV���v=Tm]��R�ֽ�u&m��;8�6bY�V@������CU}�c��t��o�����x;.�)���ڡ㪔b�]Ƴ�#d���(�a�ʘ\Z5+�mk�(i=/i=�$��sm�7�
ڵw��g��[�Dt2�Z�*gU�ې�wٲ#n��E�3�ٴum0E佚���D-XDe+��un*[��a�"˖�-=�K������t���ŀ�mHܾ�2�ih"��L��##��4g8S�w�����a4+���@��6Hf�'{Sc��/Q괢�-� |Ʈ������M�_\ʢ}a>`�ڤ�Q!���'M3�8����3�ښG[�ȡY\\���lr=B �v(lɨ�W�/��\�uc��%�x2���Ž���:��w��AY��GW,qP��wv�ԥ�[���ק�����n(�㭶�zJd�����<C���*FR�\��<咶T��ouD��ۢcՉX�p��j���!�����a<���q�F���
GT]�f[����9��Q� ����h���L��R���e��vu*�V#+8�oO7�cV��r��Wak{�]��6�K;]\U
k�2={FmJ�e���ݺ�JYmՑ_uJ��s+M�A�ƻ4jZJs�(�:_;�Z��v֫��+;��JNi7x6{'V��w.o[���Ɛ��n]_q�vL�cg��.	*����ݫ���*#���hU�ϡ�N������ofգxU2`��f
�fXI����t5�i��(�C�#�����\1�r��ö��"���u!�)GU�͝��r���%�� ںcd%�=ظ���l�{�ʗ}��ɲ.�u�'b����8as���S�h�w&�z�q+V(�+uG]s�Noέ�m:|2�R��\r�ʆk���38���y�b�`�tj��-�GvҔ��ǝ͊É�\�y2n�W@'�n]>͛Ga]�f��ն]#+%G�5"���޵˩јs����S��,_7j�����L%��s&�Ԟ(���M˜s7�����[�ԧ�.��]�o�칶ɭ���`�k�_O�����8s�8�NY�zn�$;&Z�f7�|-�3r����p�zӷ�c���eBQ�=���@^����|�.�d� ѧ��+��f���-�|���x�n;���=�gX5�/,�@�73e�1Ɖ��X�S�6�N���=���pk9ڦժל`�v����x� u�R��up;�iTή�`��oRj�M�T:�ri
��έ����\�&p��Y;D�t;'K}q�����51�W�Uf���dnn
T�4С|�B=�.�M��v�/R��(�}`F�۾P�7À�G��q�o�w�*t͘@u(��Zt�c6��=�V��K�+.X;�u�n���|��X�]�Oڗ� �;�	�/�u]<Fj��f�e�Í����;�Z�sEҝ�I�e�7Oi�YZ�ɖ8]�\`w��c�l�z����U.�a�����We'*5��@;ƥgEY�;�����V����2L2*�,�e`�}�vS�ެ($��PU��N��Z!}�B�f_c2S:Mܤ7�R��ek��\g1�Mkh�Kb+׭7Scf�(�&���m-ˠk�\⻧ǟ�V�E�x��B���D2//Q�F^�ַ�
�Ҳ*�(y�[��v-�˓�b�<�͢gCto?,�٥�dT\�˻C�t��G�1n�>C�y�S }|�V���ׁT��2�D�9��*؀��֌(m�G1�Z4Ю�H""`d�Y��b�����j
��T��^U���uk�0z�GI�e`5�k��k�d=.v��Q:�,�G3�nK!�oM��F������GS�ށ�]�������M� 5�Y���^��(�׷)>��ڂZ�Ql��t��e(�ϭ�=C���/p=���sY�p��ĭ��+���o���_2Zu�w�C'V2������4���6zs�v��/-Ⱥxޮ���C:�*�Gf����y��x�X����J��lzb��]��אb9V.����h��SE�sM��a���O_2ͧZLA����+cMz�q������:WO���䘜��v��S驒�b�b�FL��}ܒ"���zYJ���^���χ8~�O�e7���g8EN��sB�͝��W�q8j�'wyF�3�81�J�`�OX����h4f���T�L.�� ��*�-��W&�ŃuJe�wt���]gY���۵WE^�k3�W:�Gl͙^��
OKK�f�e�U��nr����aI�	n�WYz�o-V$"��'igmv`�<�ބ�ҍ+��xoo[}�+�N��2R�'U蒮7��U,
�ͣ{�	衴[�a�DgV�cJ�h��ެY���m���^:jj��{�e����@U�tܾ㿕��Ce9�KT�s&ظá�|x,S�3�qHMl�z�qLxp;tnk_^� |C��:���w�Zhmt�6ݍMwP��'b��c����m���VQ��O��n��N����-:�Ob�dpub��������`��wS��6�*SV9G���xN�����g`<���+dM�3��l Uq�gpoB4�p^�HNㅴ��Qi'�FHr������+q%%�(]A���5���/�6�1ã��_T�:�+�Ϭ�9gzQ�Õ�(!��|/L�}D�S��yzj<P�-�Gr*
��CCɕ�ۉ�W>���������k�n�
7e,k��3M��*jhM��e^�޻Ynjx�!o��°S���bOwWa��yIP��ug2� �S$<y��sElx� }�u
��|�r0���:��N��׬0�'��;����H���eъ��]�Q�3���;2\Ţ0��+\��.�/��|/�f�sT��EU����=GO>g%�ooQp[-<�"rTΫ�պPX��'	�{����4)�8���Z6>���mؐl�����/��tJUˠ�ۺr�'�%G>Ȏ�Ҧ�83��r>���^6r{�v��u�0���Z��Jõ�G�kG4�N��]U�W�%܂��M"]��j��#z�L�}�7i��si�mַ�K���=����F�[�B�c��[]�E[A�P�VID��L7��'R1�Bo
�:��)��
�\��j�rx�[S�Ky���2edd���v�]b�����%�^�ud�Cm�����]RZ��=F\X���Sů,�ٹ�s9��v�5)uQ=;K���B:q1G+8B�9��b١� {cCX�v�>��}�Ig����t��N���@=�,�k�-��d��
��t^VEzR�B�Y�8+��O�*�Kt�ʶzK���Qԕ�Ƣ��W���3�R6y���F�_^� ӊK�����Mr���>[Vksw��4p]���Y��G���X���v(y�xҜ9)��d�Σ�GC�-d��N��NL��5�Y.��p�{��zRV�6	]V�G�s��&�Q�K�n'yw�Ç��=�1PqY�1B#������m�Y[�M�wu��ƍ�p�Ф�1T� t�-f�S�]C.�V�tTK��֝���w)-j�2���:2�����3]}�v���:��l��q_/^��s�J�7�FMLTT��CH�O,f�):8;��_d��M�7��ŰL[B��̭H^��34v�[M� ohU�U�D���p��Z=���N��ń	2��O0��t�(T�}Y��㎸>Vx�Tw��Ą$r���i08���
^tט��+9����x=��̤ƹ��l�� ��ַo/��`,�ǲ+fÙOU�ڶ�dS�X�]ܾ}z{eo4p�k+n�V(�Hm���M�K��F5KpMyo��Շ�5�v2�X)��*.���,��a�"�l��r:�佷�m>���W�&�Ou$OG�-�?���]�k����<�@�S*��s��	��w�)M�J��^f����F�p�|�3d�w	YcC[�⎡{���:�\vݍT���c���֞��S�0�
3�Iq��F�ќsq��hqQ��]�K��:wN�ސOa�-�t7c�pc��u AbK��2�O�q,�m��e��y
���m�[ښ!�Hte�F���J���#m^e1OC`���¬rZ2[{�9nΩaÅ���j��A��2+�J��$	�_�Z�i�& ���vA�*h�C5+)����?w��   ��}�'�������!￾{�{����Ǿ��^�W����z�^�~����}�	{ ��
�����٢cp@Ce`�Qt��U����j���_b��~�Ł����a��P�����;�°͍�Չ��.�}��?_�'���Q©wv�+v�gn
d�
�0��z�]�æ�mUk���Nm��R<fq#�UD��<�4
�|�c�6�ͧsrfv.�h�+n�'��mÑ���z��u[:���aY'J����R[��|��۰���Y>��ǋE;sZ��5X�RDS���uE����)VҠ�-�k���/9�[t����ZQ��f���e�֘����<�U�p��4�]u�CFK��u�{�ڝ���W b�]��H��-�u�����bU87H���[XVlP})\um��{f'oHM�y��l��Ko)}��|��2aW�\���*&�//x�;�����#�y�qX��r.���_0np;��
��\ �D�kcƝ���m��s�tL�'�ݬ���AJ�K��.&��4��������M�rii�+۳�N��������ΌK�&��и쭭�F����p�a����z�|���x��3(�/R1�e�:q�&����%u����PYq>W���3��C���X��R�-ǷzA�i=�ɸ�j����j�S8G��K��Co�3�t扪�i�{3�kSc� [�$��'�a$
�g�D���	�gGT)A	28a��&CFbI�w�����S��M��4�Y�MC���M, F��q�Rd ��p��$h�����h"׋�B��M���E�R��h�d1@���&D1bF��R��c�u�O��FLh�ZfA"��%3$�(�E�A�Ȓ��"(/��^~:��m�IE�\ĔjCC*K���$j�C4�d"a�T&��B�L$Ŋ!�Wv�Q�M1$��ri��DDcyݒ�Hj$����fA	IL�4m3뺉,�201��%b����G��$`.�2�
E��� :�|�ݒm߫�ewF��Q�<罳��BP��=�+#yP\��6�f��i޺VC}ra{�����|�{9?(���;��$T����A���p�;K�;m;��f��c����nY��ׯ�j3:F�i�6L^�c����+j��%=	�Bz�;�Xǫ�r%���'�9�o�_�뉟j�yE���I~��{s�5-�&r��Yd��n���1�}~���^�\&S2�r�׽~MVN���=��7��j=�,��g��e���s�ە:��Ъ���+��R���؝��n5���ٳ���������QT�x�G��m�^�%�s AN��j��m�أ'�=��;��޳��o��ˢ|��.]���븫<���+�&Z���ix�<�4Gq�oX��v85Bo�N�
�s�9t�zMW�}P�߳��a�"�]��G���6�7�g�d�<˥~�Y����T�"Nw��#�dͪ�i;��y�h�ߋ^���&�[3`D����N���;][h_,�Ȳ˧}���������!���V��w��+�w}ͧ}M�2���m�Q����s6'*]��{d�bF~���=�6�˳D��Q���em�T��(t+8=��W��%�L��s]y;	��-9y���+7o�y։>qQD8)z{-�k�M�IW���>�����zT��C�pYs.�ͣ6��
YC޲�e]{�uw�W�]J����9���ot�vhU�t�|��*�MTk���_�0��3�·W�W�ڝʞ��ۈ:�������w�¡�`V�ūU��k�
�po�#>����s{��uԖ�������g��/���OBNs/�N�==�{�ߍ��0o�Z֫�Ny뿷'W���w���^p����ߔ�Aƴɤ���Q?wg���\��9W5ۀ�;�Z����[�n�U��}���X��Ln�{	Y3�T��+�:7+���yF�ɾ�	⯝�?Tof������E���۵=��nP
`�<���?{׹�{�R��~��Ф�<����=y�Ք�Eo�iV�۟f�OZ��g.b�ɃE7�ݹ��w���'k�r*ghy�R����4��^�m��Aw�hEF*�e�k8�{�e�[!�<s�+�ܓj�D�9kwQ��ݭ�q��X��ڪ`�S��ɚ�c�S;'n: �u����`�j��$Ëw��E7us[5w��=^�x׈���q'���_y���==o���������sfv/�{X�r����`]j~'>s���/Y��)r�{�O�雓��<�M[��CQ+�-��Ec E�����5<^��3͛�;����߷@�r/HE�7�M��f��>]F�c��;-�mf ����ᙌ$�//s[B����
�!���D4]pg������u��JY���b�s�o��I�{�uOM{�z#�~��S�G��¸��������7<���W����w5�8&'Q-l�̐]+�cY	�[�}��ͭn���4P���;kn6�78=(6��]{������!�{��+<dͳЎ~6��x��ѷ�)[uRY��3��%^A+����x��đ�2#�K���O�����?yw��U^s��q8�XY��5'b���R��{ι��a�DF�V���LB����Ys������ݺ�Ӻq�d��y������{����v�y6�Duu*����y%~��j�հ�������f:�3C}��v��`�]p���7{�`�(Gկr��+�K���۳<f%����/R�r�����o烦U"{2��޷� �۷�P:��q^f*A����"$��5���帍�;>{�R����	b�w�:W7	����S�C`��9�fNW��^ߍ\�Y���;�X���t�(<�{��I�U�U��9��k2eB>�E�ޓk�{+}��W`�P�܎oW��JZ��W�hWBA�;��^yҍk�i����^9||9�X���/>g*xge����r����UWպ�b�����.�2��e��#�b��L�mt��~�mg����h
��X��G�_��KړXՉ���`Y�ou������sf�����U-�y��@/�?{j�k6���׶D%����鋢��Y�k�W��K{�L��7�S�<���9S��,�|��:�)^
x�?*́��N��7�_���Jqo�z����$�j{lc��r�<�b=BVf^{���^j�ޙ��ń�@�"Q��hf�I�wYf��I�'�c���1�m�uShUUwcym�ڃ��oG�iV���!��z�]L���F�r����2f�}��]���\���=��譈�	�I�&;h�:��i�/��tik�ܓ-��w�ÈK{�gW;`���s"�p��vz�2R��Dz��.���k�]��)����%�<4����!è'��nm�����fR���l7���K<�z��;۪<�=��))/�x<�7�=���}��s�<ԯ�m3��9W�<��>T=^ÊM^��m�w���r�p����rb'�����e��K� ��¼�$���}��6�r��Ŵ�֩���榧{�OBQTO%M9�68��|sFX�>��]P�l���뮹i߹?W���{�,��qV�G>�==���O�Лy�mS�Ү�]�-��<滸��O/��i�\��u���������y�|��Ii��#��b+��}:�������p!�/��3n�]��s}�^͝���蘆V���ą~��U���UՃɰ�S�탦�vwuAͳ%wc���J�/n;.��u��g1..Hz��W2T����J
�2� �|�h�>6	8f���.������&��ꜳ2�m]e�&5�}c�L��Ʋ�DX�\��V�涺,�\�HԽ�Q:WJH�2r����<��Fmܶe%��L�s�ޕ�o�mO{���%_���/��/~����u���ʏ����k��Ny�|d��>k<�����ur2���;*h����P��<����Ox�����}ҭ�&1y����z,w���U�C�X�g�o�U}��o�������1Qot7����i~��D��8�gS��y�F0w�9�W�; ��r~�f!n���/1�i]�}^o��5\�s(�����Y��	Gu�x��]"��Ot�~��X̆��DT�M�D�0�A�n@������7���(��l�j
��2���~K\�u��us��~A�}*�0�4�e����N�m�]�ۜ�n��/���'��.�{�߸��Q0˦�s�7�wXޛ�\�}�7��E���a�����yo*���E��j�t��d�b���xv1�hͩ�oU� )��/�w�[���H�7~*@�zE�Q�����0W&�F��VT�x�������Y�v��X1^�@���r>$s3l!�k8�,n�s�}6r�C��bB���,w:�ӟ-�������ԝ�3�HF�S�I�zk&�Pٔ{�Oh������]���&-8���̊bLLnu޶�q����q�����t��/��׽]m�i}6��kG���xv��dw�X���`Ḣ�j��E��/�S���1F_��2-�jW�y·�ʸ߻%{�����C���%��-U�qw�[$�'`V��a�o�io-N"�5059��{j�rr泥�����HzIj��{��;H��<@�B�n�Vʥ�3Ib�7�P�w�s������[)�g��y���aۓՙؠ��4���ʲ�>re��\��Ox�K*�WW=}7^l���þ����^�cS $�;>s*�zoَ]$��{�����3�jנ~�eo�{�1|��".����4T'�����UОx����?VZ�<��1Ξ��9��1}~Z�Ώ���}8<�ᘛ�I�z���`�V-��yW�&'D�:K�¶���`�����܃'I����s[�
g2F���������z���zl�8u�i�]xKu1�m����u�t-�]�-�[|ˡ�VN����tcFw�&�Β��r��U��p�L�Q3mAqʄz�=59/��Q��r|"ю>ʣ2d*�\�m���z��߼1����߾5�� LחR{>��tҺo�=����86NW%��מ^��k�s��9��D��Һ�{�+O�Ejf�&�#���3z��[����9��g�k<����K����~��ooxV�风�j�{w���t��,�q�O���O[^�E��7Z��C��|�Գ�Y�͆��PJ��\<:��Z����g��v-~��`��=�I�aQ�]�J�h��y����^�9��m��]N+x���'T�kW��ty�ݧV}ϼ;����w �ǲQ��6��7�o�t���-�̩�w�Ϭe���\�N��f8/f�d{�)�V�y����v��y���=z�	[��{����-�g��j���W�Z��@#>�5R��� �}���u�������;�|M���QlcUqv��Z�6d�:��<�wI���F��H��ǡ�@/9l˂�\Kׯi5�@��z����Ŕ8iZ�م��b1k A��zNr�rpc��x��
Έ��M�4�h��n�� O��a��9.��G�	�]��fn֫��,���9<������ȰL�{^���z��y� ���@����;����,����?t.�<�j/���>t��ue�O>Y�����y��ڬg[��{�oy��o���{�y�'�v��{��Z��F_�u�
�"���;��'��9���W���1PzL^��T8��s�my�/�D����Dz
^���B��9����G?V�K�r$���vg1�}�:R��5CЕӪ��k_V����[���֧\��[�{تÚޗ���u�u ᕣ8jm	���NV�y���얽e������u�o��ϙ�h��ӄ�0'v�-�go����!t ��Ķ��/L��w3��5�]��ꉫ��V��y�����(ׄ���T�'z�{� �t�'�:{�+ו�������>�v�}��r	�#�+6�a[2'�Xũ���'vi5"mJX(��z����̆T��K�t;n܌6aF���y7*�n��k�ʁ=�>��s��,Ю\�ԉe��|xRmѤr,��S8.�eNW��R���ܭM
�:#��;��swj�s�ٌ�%>�A�n�sG�<�</�Mg����=��u�<m7�mh��]��U6c̄�7)����r�M�gO��Īܱ��ݴ�罊o�m��U{y�����Z��\}"u'��s�ګ� 2d�`��z*�ޗ�->����L�������w^Tܡ�Fx$�n��륮�8�|�'em�x������BΚn�woI9��$�ר����`k�y�q���ҩ5��\��'g���[��k��w}�\�j���K�#��舨G��_��U�O��֯M�=��#�K��U�W�݃*r�����R�>�xh�J|���v��j����O�۞��
o)[Wnub�2a���c6fIZ&O����p]�O�vy<�Z��Ǖq�2�2�?q͌KK�z>��ʸ�x�e����{FP��x?����z���W�޿_��������g��d�9���Q]�к�����"a�K���m�;nK�sɅ��L+X��-hOm��B�����kio�S�zbx����R���Ҏpc6�.���7���.J(K2�]�:�ˌ�PK���S��"a�b2�6���;ܴ#W���/"}#w�1�3N��S$�y�v@wN[p̬Lѯv�l�j��f��[wcpU���}�bˑ��W`�a	5�JV�)A[}��;p7�y֭�H1���1=�1��E�pI[Z0�&9��uv�n�W1�u1f�|�0�	�)�Q�3\��ǑI���</nu_V��>U�^3��٦�ڌ��jR�Q���a���Ʃ�v���,�ⷭ���V*Sc�K,�Qةjee���җ>��%�'a�n�9�2��ǜ�wkn��˅�si�eV��	��-oXTrp�Q5bq6��F�Fu�=�"�/R ��H0�;�)t(�eEq��yc7�E\�u�戦��ʃw�΀��rn �R������xj([�j=��j�,͒oS�fj�[��u�2m�j2f`�;�:�>�X�&R�`�������
�A
KI;C2��I9{�j���}�5�-J�8��8-k!Yo+���1s�m@.��S-'3[��I�ov���k��؅�5Y�����g�b��;v�!���V ��lg]�;l�*l�1���Y����T�q�X�1�����]�9yb�6�R�m͠�X�)��GSA�e�Zv;�f�7X��9�Bʥb�ty�f��V��F�T��߅gY�ld��� ��u����t���� U�]sUī�5)��R���v��,,G{�gZ�ē��Wȋ+�]�8�\]}�,L�(ۇX��n�\�͙YN|+6*�y��;��r�rř)��M�j���#�ܩ -�K���Ws�ݯ�܆x߽+o���M����D�z����)7ӓ���?WL����|�W1E8]�!,�cӡα�VԯϮ\ݽɐh�6k{��r�-[X�V��%�����������Ei�TB���wN��=�	��mu����g��k�VQ��� #cjay\8	�-�D�rV:��O��u�%!������wO�s����P�z��m�(0\6�`�g����y����o�6�����_FWn%I�K;����R$��k��N�oR�kt -4(#hL:f���DsJ�2�Xd+W6���qOMV���K7Hv���=�_&��n�#��K�����;n�]ۧʴ|�_m�εi�otrA=/Z�(EH{1�8����:���g:Ǝl؇.�H3� -�t3)�㜁��6��nC��u���Å�8)Ѧ�j�u���ԣ���i�1S�0`U��?Nꗃ�Ԑv��PV�j^J��v��ݭ�D�x�p��W'4��N��9/�����ܻ�ح0WF����t���s�!ݛ]#z�j~��{�$�����ݮE)��nI(M�!r�9IEx��Ld�(3(�\�!($��dN]���D%��&Ld2���ě�"2X���wu0`AA�;��Q�����La�*~]FK�1B�7�hֈ`(K뮱4�mz�<p�C$Q%&4\�ۨ��wv��]Ѣ�5�]��sw]u#���s�L�W-vc��.vh��JI�v]	wnl��;wE!7:.L�ݗJ�])ݺ�0�Ѥ뫚 ���t�.ݹ9ӗ]�˻�0�wv�厄s��u�N\�;7t��]7v�^<����g�t���;��v�w]�u�Ќ9wws���.�:i�s�F��5wV"M��6#�q�+���ux�7��\S]݁��}b�?K�˷a$V�V�7t6�<Y|t�{�z�e����D�7c��8 �ҵCu�-Vr�
�!���>q������XT�i[_�1�� e�[tG!k@(�ڼ�@XQ4}Zk�1�b�{S�����c�!����s�˟/�����:j�K��q3U3M:���訒�*��c����~���������O禣�4��ޚ��07��c��}�FC�?��ݛm0X�^*�<�{����d����@j�i�#!��.;�=�~��7Wڦ�L݆]	FX��.��{?p�R���������q�9!�[\DK@Y����~��h٧e�R�	l��/�\E]fLB��y�ܤl}�G��>��.�9d���^�T�p���jJL��L�	_�u����7yn�ά�G\rm|]z�ƛ�D������Y u��Q��Jw�YQ�H���a�&�Z��g}҈�O�!�6<&q|�����w҈k`��QщE��c����Ic�v�� r `�{���������?3�/�G�<�Z?�i�'��\>�|����P�4)�#t�n�͇�*���@�[K�_;������O��v�4Ρ����}B'��ρ㖙���1�}L��~�� ^>��ׁ.����h�LS1v�SeÛwN�S.c� ��u�.��o_*�,淘�u�9�����O�@����z��O2VA�L�N�����`J�ۮ��4�3����Z�����yD�/#@v��^Sb �T��7��gH���&�Н��0p�U4��{WU�J��W���>�I���g��m��'ZHXF_1�C��P>,�`بN_@���ͩ�ȩ�S5�%�Z��T�{�n'�~�����ok�H��xT��_��uJ��Y@�^��������A�i����S�C���\W(�}��񿶥�˶#m����p�a�Yٷ�?o�#����lش}�t�|W����k]LJ��EE���3p�~������)��`��8BN�)O^��`�$v�\��ym�����bg���h�3�	9y��I��"{曖�(|�	K�}��`��\'�3|��l�|s-۵����6��L�Tt\��.�v��S�~3|F��3%��X�V�#����Q�0���v{��V `���N���_���'9�޵_�~��;���7���~w�T[����O)�
��<���ѝaM���E!$f���;.֠ue�n�6�v(���H�ϓ�e��yt�(Ϳ���u@�j#��KS�Cs���T�k5U�T�i�pԪ�k4�D]k�(�n>'�@�h�s����$A��r���Yq�Uﵴ��ML��c�-����T��l�SvD�����<�;��jR��� �����*y����*k�\;�ǭS۽�9�S�~��{����Ӗ����2֔��$�+U��8�<��EO�(�6�sT�|�9e
�a�������ǃ�cX�k�
�f'���z3]��D!���|�"�b�b�Sg$6[Ɯ5���ئ�����kҦ�y���3Sv+�L8���]k��M�M�Gm�9�I�䖢Ǹ����7ծ^�z��f��ZS��=�kf	���8<\�L%Ջ���ᒻ��H��jU�%t��0a�ʐh=�)�g��e��ͼ�̚j.a;���0t�R�P�u���U�s�ݓ7�ÍJ��E�ˏb�*A�T[�����ȇ��v[�(֫�L5\�jdjS�14>���p0��Ӿa����F񡔆
ι�l��]��1�!ߡ4��<!�x@�s�Uzɣ��ڮv(�uɌ>㭔gM��II��
ӯM{m�':�����#�z���]G�=}��q�*Poغ���Z�{�6[8CS.{���ojR1ٚ�P���9YI6��1_y�`a����z���q��4vˍ>�a+m��"�j9��Q~���4t��X� d�糚�j������L�\!k���Y��/�ǟ;}:dmy���ԗ�&�yU��[_>༸��6��VT�wm:�3�`M�Dځ���ڵW�VC�
Oj����ƶ��ވ��/:��b��e40ݥ���r���N]�1ٺ�z�cWR�2v �%�&�s%��P��o�$��J�[��\�
�>���5��At�w�^�ɜ����jC��±�nJGǔ}���2������<a��I�n���U�}¾������a)Zɼ<�6D1.����q�5;Ǔ*���/W�K�m���y暔�f�z�M{ٵ2s����Y�z�9�M���X�-n�ݥć�$�x-��F�}Mç�������I��w���Gx2k�G�v�iQ�w[|�-��W�\=G�"����觼����k���2�����
Ļqs��"��d١��G0����� V�~l�Π���4�@�Mi,��-��&K�ד�AS�y�3�K�?E�R��wJ����]b��$�Er���0�d�T�'���U%|��T�Ԙ�#5N4&���>���:c3r!�bh��J�H�%�]�V�&e�%���:�q�<�ꇒ(o4Ӱ��G�* J��5^v	�jk���l~��In�sV�:�;L+Ѧ�@�w��O���S5�U��Z	�ִ�!fBݐ�C.O��C����9���<�q�qƵ��H�͞t�Ɣ�-�E�m�9��T��ҡ�8f�ي��4�SE�V���!�|8���D!�LӐ�:��%��*�$SG<�L۫��\�k������wpکJHZ�.W��*��9�}[k�-z �&-��U��˥�gQ��Yn�����bFҏi)Y`Gy�����Y�EI�P7Ηn�hu��r�-��}��|#1�5,�t���k:�"b���1΍A�6�ٲc��y��ղH֋꾱Ͼ������Y-��T��O>b4?���y���.C`:l!%��"�]���5��f��eԪ.��*pv�س�հ�:0�ٗF�����	���/f �l�t��í�,0ٛ@��d���E�"���G,��z7]jȶ;ŦS�y���<!��������e{`4x�v�tqV�bډ�N��Pv@�X��z�u�К1O��6��z��V�q��|�r�L`Fֿ��� �i�����I����U�Z:���2il��e@���i��-��S�X��#_�]ipQ�y���뭟rvg�فgQ��6�X�\�c�t+u�
D�lz��1|mB9>:�n7L���6����V�\^�'3�b�T&��8��X`�ۂ���ګ�Giz����yw/{�C�P�����'��-/E�k�|��2  �ް��XI��]�l����MHI`��ɝ{"e�H�|�=y�������X�%Z�̒�IݫÎv���F4���$�cz�⹥��|P��UI��T��Mq���1�ܶ ,g�b�e��u�j���xǺ����q�z��Ⱦ{d������@IM\Q�{0YM�%%��y��� �&��������(�k����h<�ۺ��E1�$�N�I��j�{A��G�u�8ջ	�A~@.����N�������d����3�C���e��ہ��r�1m4�V�S�����h���q���7:u��#^�W�>����'�^��R���C�[�0�f.��3�I�~��Dc.�'�[-O�T���df�!?��{S��t�e?U��D^Ka��;6�,���yڇ)D3�Rpw��@��սj��_��{�y�.Z�gM���v�z䒨���-���q-������^�J���EE��#4yi��[F�z��m�Ga��M�4��r���v4�y���X��ܪ/�L�`�b0^���?�b�X�6�?hx0ϯj���[���^�����n���9ē��.[��������t
ދ���7nn�)lu\��M8���7)�T�{oѧ��z��BUԒ6��6;KB�!���&����*�j���Yc�*ش�і��I�o��������&0��)+ρXᚉ>���S2�l�f;҅<I�;��sy[����H�,Q�$dwn�&q��F��a�
gAb��� 2�K��#�����_k� ������y`�K�K�כ#�e��c27'��A�3��l�!d���x(�໭˅2��-۫P�s@v�y2W�`m2��5����t���˸��k�X@�Z7Q}��\�O���G!��g�k�yR�I�7���f�5I#�=02�(�4�hpm�c`��_G��m��m6hRќ�d
Ȭٝ��/(9�r5&�w|�:���͚����d�&#�ԭy������d����4O\7L�Ry��aXdMy��|����#����tu�owF#(�bR�/̗� -h+�J��`��k7����Be'9@E�b�5�YTN�fj#8ȹ��S|�GS�$b�e8�-���b���1�o��N��z}�����&˚獚�Y�4��A��Y-٪fC67d&u"�&�o���ǖI�k�L_!���g���|I¹��4��	�nGl�����TGu�e�[���NתUv��ΠRҁ��"�gE:�� 1�!���y��^�䗷��߀/¶��"�����e����^��a:�x���[�ף�Z5_�d��������M��-�Oچ ��#����d�u�PyZKz&�X�ŭ�S)������ꦬ�5�^�v�>���6ׂ��(m���بbԨ�d����X��=�N4�����A�v�z�]��E��	�L�y�:;�m#tۭ&s&(b�R�Td2�ؘ�9����=���˰�f�ˋ=��Nʴ#�兞�N��a9BٔT�7��d�dz�*y͢�"5��h�a��r��v)~Sn��`�'�<������F�k��+4]a@n�PU��$U��o�`(�=!������H}X�0��=���t���>�P򞕘��KPh(��֯�׽�˧�fYS�5�+:TEr��e�z�g�����E6/s�]V�D��ι�svJ�ٹյn�ֱ},��4P���U��Y�-��V��!J�	�J��O�<<<�����	������4趻�z�bO7�֨�E�q�¡@k6���➠�eN�|x�(`�TjXvZ��g-��{Q���!� � �F𶙍@�E:����&���S�!�i����n��}?6wz1�rȶe�h/�ڣ�ܬ���z�$��!��)���<%�����@^Qz����V��F��U��F�y���{ܫ�`30_[L9�	�V��`�\3��jbyY�};��\в��c�Lr�[�%V��j`K�l.+�0�_�#�kC�]-�-�m�?�It�����Yk�GYi�Xc;��_�>���2;�@pr�ƥO-m>Jm��L���>�z`����3;[��9��G��'��� �^��W��{v����F��Qxh�eՐ?�3���ӫ'�v`�s(;#0r�&�%�-��)t0�o?�C{�4r�7�a�����]̳eP�����#�7,yj���vWNL#ߔ��9�?�^��k��Uc�u�s}Z��;���S��̭���]�$�>��r&Eu�2J�����(bv��UJx��D����m~A�}���X��/�la ���j��渱��߃:lػ�j�k��Ѳ����e����V��:���<���=�ױ�%cy�s.,�)���x��Y���7�+C)Ias�8�v�~<KLMdw?�r���u�y'e�U��[X�j5Z5j���Y�	Y�K�]�WPX��1%ڑ�Nx��Z�Gv����o4㰉�],M��F���7P�VT�[���֚��/v�g���<�ƙ���v�J�?e4�-J{؝0�T����ե�:�A��g~}Vr�Q�C��`��!������a;ƑD�(s6F�y|��`�f�A����`u�����*x3�s�)���f�f=*GVD����a�M��4W���/� ��{�+u����!��Q���/,WsT��]��[T{��X���Ch:l!���o��	��2gս���7+����u=�&##t'!4(/+^�>цwޖ4�.�?>�/�Ltt�A�߫�s�2bγj���w����j���7A~ʞ��g=#P�G`kp�ae��p�n��}L[�N�/��V��.�W{� ��)n~.Ŗ�>�qVL��1>��Yi�`Fֻ16}x�IL\�C�xR{Z-Ko)vP	�hd0���e�y[l��,��˵,��#����	E�G*�>��f1�W\:҅z_�l��qfOl�����D�n�F���|Ǎ��.�Fy{:��R{�i&;{bV�������Ui�;�?������'"��Yp�:i>��l�/��HA�j aji�l\3n���Qͽ���uK)\Ž�p�O`�n��G�k�o��N�Q��o��`���X�G:cR���|�<,�������{�z���j,���Ŭ�o�tT5�,�	1�*u1p���<�hyv��K2Ƨ=�`�%����ׇ��6��eU�t�=��;�X)͘k�4����0{F�r�v���$n�nNE�?E�����7o_D\m����t&�O;�ﾹG4v�" ϝ��*J��5��^�	��z��D���;�1p{�&��U��I���3��W�͕�O��(6]����L^P=�L�i�W*6r��sJש� 
�^}u���e����C��@�hzҦȻc*���7I�{&m�y`݉��}i���o��<P�-�t��U�u؅�s
x�J-r�u�p� SOk:�m-�pݝZ�b黩����H*��7i?�X��Zf�QF'8��L��g0��xᕫ^.��;2�l+����.�ie7_���m�.��YX�O�?�P������h�a���������B�ov[p�����6��}YM~kj5 f���Nq$Қȳ .�5�H���R�+jU;���ƍÞx��a��x^�Bx#���<�<��J�ӎ�F�c��������=~�g����z�~�_�������y�bVfL����cz�`���q����/9us�n��pr�&�R��������98��z�Cd�na��kC�t�]��e�g��///v�X����ivŇ�j:{S��T��ۛmʚ5��nwN�ɺ1øi� ��v�,������u+�{�4f�.�e3���92i�zJ��ZW�eh�k`�>�}n�(lݻhZ�s+\뇳:tT�N�o�٩���'5��U���7;�i5vn�=�y[�͛Hr������ �`�{�>r�-,��W�K�U`�=
��uBݲfk�d��dZ�K��c�nlΆW9{��r�kG��F�{��ͱy��;m�MeN����e�
�p��ٖ7u�Q,��n,l��)^��;�gm�*\m:k�*�m�XLl����嶉�x�^���}-�y8�ɝ������=�B��,��We$�%r��п=�{p�$>�> �o�������,Sc�C�]i�ޛy��ۤ�f:5��x5�`ŕz#Z2�Ry��a�&T4֫գ^�J�:D�l@MYݡb]%uh��,)�u���a��֠sa,+ ӝa�~�ES�;�K	0��qR�P���er��*�uգ��K7X7
���j®�򗂝I��
���O7�<5|����!4�Y��e`=j��n���ՙ&s���:ݮ�UolfKT��s�.ÐF]�z�F���l��=a�����:��C2�SZZ�����[uo3;u&���⺰��xT����uxÑvP�7�;�\¾�M�|�m 9�����`�m)Y,;�K��-��ee�j���
��AD"����h���-Ŏ�Ky<]�����VY�U�f�x�I�� ���.T[c��x_b)�L]\��ۻ���h�y�j��eM�)�)];Ϙ<s���{(t�Nr�ef:]����G�m[�z
&6�z��}����yѱ�o[��[7��sd;Ҧ��y9��X�3,��S���9�u�9��ܭyt��t"г��~��b�3�]��G�q�ha]OD�<NN��-�J��b��3Z�dV��[@���o4ori�pc�ݙ�˸X�V��l�{�܍[���y��e=�v؀��V��_#{)ر��qy͓n,m�j{����j/�4P�v�o2�:�5�]�0kM�gi�q��*= ����|�l��w.R�J�+t!��[�rޭ�L��Ko���|)`��^`����]�u����,vn�x�]c;����ET/���{r�y�U����Y!�M� Y"r�G1p>�mn�J� kV-�&�hísh��\����;s`y���;s[���:�a슴��vY�R���@ 4�cj���X_���%m7r���@�P�V����߬h9�	,vМ�Zˢ7YZV7/�`�,s1�|H�y�*�СBQس�۸��m���"�W5�ٮ�d���t�0!��yY3�n��3n��K�ie%�����Yc��q�Y.n�F׼���G��i4޷t�0�s-!��p"(8�`��Zww|���|����g��� �ƹ��6��]΍%˩t���5���Ţ�n��c'מx�w]s�#2����1�����Ѽ��.s%7'u�Ѩ�ND�#D�ʸk2#�4Q��&��,F��ߟ;>�]��lR&��u��Ỻ0'5�,H"�ͳ��F���фۛp��F���^]�g7KA�t����bѬȣ
�)"Л��6�I�J,Ȣ��Di�&��E0эDRQ���u��a4��,��_Ni�'9F�b�#���M�#6�p�Y1���ۉ1�b6(ƍ㕌fX��Y�놓A�Q��Q$/W�8��4�{--2C�L_B��Q�:=�l��A5�jJ�����i���>�	�?7\�;�N/4�R�-pr�:'kq�`̣��:폕YvN_�� x -*�N:t�I�N�����j�2Ս�Rv�f�<��[��0��e%y�����T�qD�e�S"��u�wL��\j�����B��Lm�ҜA�
4��x�0ڕU�ز�ta�mBn���4lиr �`��M�c� Z��������k��:�n`:�* �'��ʴ۴�'.;ۀ�ۓF�hh��ܠbt�a06�.`�y���8Iʸw�=�>7+b�@&s*���D��֝�HH���)l��z`b�!\$+҃Z��k�~k!�KI�G�;i�
1�P3r��	��#�2�옙u��5y(DҎZI�b�9��]�����3�(�r`��+�,����5Qx�"�5�5��Y�&_[�:�EL�~񆇹���!��Jټׇ�f��^�z�~��j�Ջ�3�-@Pמ�
��)�[;��H�n�@��Y^.�gE������TՅ5��Ѽ-�DJ���#�ŬݕԽ��Ҏ]IX��G#q�a9�J�[	�{i���U;y*�ݱV��K�)����d�u�P��Ϣ�/|������>z�z�(tmdҠ�h]���A3�ݥ]@�r�'��v���gM)lylQd�srLY���zT���
[���=��]fm����Q4-:���
���.�܊�i���읦���A�TU3S4%�QZ�����7�@�e��ǃ%v#�[��V#om4���潋>  �v�vu�3>����.+i��*�l�[[#@>z}��aJ�Y��bΥa$�,��R�پ��%�;��U�-L��<9(�J롞�2:��I�(�~��Vv��k��O�<���Yk�9�J�I�8�\'�4���Jr�֞�E���`i���dW��Pݥ���s�H6Lo(}R�@vsU�^��0&k_m���a�FK���'���`S�rz�R�jh���u���N�W$(�񶳐����u׻/��]�J����z��F?մӝ\�Ң��|�]�]r�Aʹ��p�\ys^&e|��[��l}>|���ˇ �A6��1l֗��kF����@z����</ʇ��`�k��_�8�ȗ�ܹ@���+y�E�Qs�y����5�S\�����fڡ�tw�4u5��oo��*��7������vZ1���,;[x$6��:�y�q��y�UI��*^�7D��@��*锶�l���347>�H@p!S�&�m	�n��m�HY��䍗�yM<!�f�iXJ��jg����?�Jx#L;&FGׇ�^����i�fX�7*ޘv�/]۴�4�=��L�4+�1�":W8�9j�wZ\tQ�y�}b�o��@r�b�h䅅��S���>'-bsuv����C��ݚ�5��6�5ˠ�k��m^�*���h���{�n��廦��_,I�|�`�O�b0�j����9�2���ݔ�E���Qyi!,p7Z��M
�V�m[�g �2�f`;#[3�ܤ�Sl�t0��DI٫胆kCq��Khss};o�XI��ឭ����]�t��Kڂ�yf��d�Ca{��0��]-wZ��W�}��ܐ�u~�2���;��L�\3)4�b&e�c�䪜#�����-v��UO
�)�/����x�'�Je�A,˦�k�.�ڌ)����ڳ�(ޜ�t�C��s��$�
�g��z�Tr�E��@�ZU)������>g�ޣ/עa��+�h�{[q���:�gxӂ�I�,�]��0��@Ì_��QD��F:mQϻh�foH���*�ɮ�d������P�5�4���Vp�YR�vs�P��W\��8<k;��Z�p��e���8n��:���[�M�l,8+���3�q�����Չ���nk����S�_Et��d2̔s��ƅ喽�7��:a`��8�8�٩�b�~>�̫Z���/�͑[uW�Խ�4].��U���n9�oNFg����	Og���ٴ��C[ܳb��H��|��=u�V�U��"�辨��s�u�LS/��k5eFݝ���n���)֪�X����眅np�0�hLyH���M�Rmcd�S3lQ���| {��xx{��y��SG94'��6�>?ѩU��_N�Ҧ'�Г���f�GcX��Ro1��X]�t捥M�<�1E��`�X+S��qf<cΪ�k������/a�,:	��x����Ǎ��D�D�a�ߓ9�v��d�a��*��n.a��
� Z2��Ц�\xA�sk3-��
#���:�X��>��[�y�c��2'�Ȅlbj�!JV�o�};����f7�	#�:r��{��Œ�(�8���o&uGf[�lUTCVuf/ZU����7ȿ�����!�ÿYaf}t�Uʒߨ���(�o�Mײ-�m�IoTO�lu:�W�#�FkL����u�^H��DW(fi�"�e�7E	R׫_��:J"�^���p�s��98��1�,������V�>�ת�)��������M�8U�u�����8���,j"x;�x���%��:)�� �.�������]b0E˔��θ��T�!��l=[�	I�?s�p)��l �7b�FZ��E�N�=���b6Ev�QW�7"zt���z>��+����%)x�Wl��u���LlҬ�~����b�=���m��ۢ���=W)o��̜�T&�αg�������\yG�gi$&s����4�FXBPl����u�湻k�r��k��ɷgC�ÖP[�)z�mm���I���[Tm�Z��| h���0��'�G��z(�1�Nԣ�m�5m��6��sM���4���C��e�9��	J{�͎�Lv��3G-��kD�T���F!@�~y�y�����K�&~(Y�U��W}�I�z���5�!�u��	���lefo�jF�8��U�e��q�6`�ys�Ɔ�h��K����~��]c�T��y�Z��8Y�O_�2]n03�X�@g >���$N%9G!�1��oyC�h��)�J��z+��2��O;b�<������A���*�n=Gd�����N4vS����f!��6��qO�͇�7�6s�����	�n�sƗ�a����c���DK�Qr��z�B�ܢ�mZH8h��^$\*����[K�z�[C�'6��_t�kz�Ud*-��Au �λeG�F��� �CF����ki��&�l�@׿f����Ǿ��s����h�+��&C�<��/� Z�W(��^�Lѭ`���j]�����c��8z�g�J?;��z��(?sq4�p�������ye�l3ś�(J||g��i;rz@�*Oi�?Cm����,ޫ`KD����[@�K�s9��6R����YJP�\��>&��{�t2f�r�쳿Tf�����ͽCl��ƞ�L'�*9��7�+���A7�X�nάn="�{��}�ϟ����ֱ�F�6ڬZ�A.&����M-6�:�BL	�q���*G`,�G1P��hz��p�6:.pu(>V]R�Pq=M��{W���U4E���C.b���)Z/ݰ�Ԋ���YM[3RPjd鍼��#��n����_�q����_����~�L��z�LJ}{�	�q*VE���S�;�9{w�3���I�VS^��վՕ�y�S&���엢Ǹ!@J�Z/�Γ���U�	0�sR�*NG�#&u[�HĔ�q��J�R.����Q�V��H�	�,�9�{/Hh�����M̬�S��l��;�$q��B�d"���d��H�[��/-�������K�~�P�.�c�gY|L`�%�t�	���6�9A	��OD��1R�0�:�x:+6r�⢺%�k�az'��g :�O�������o��Uzɣ��mW;YFK��'��U�-��
�[��ЮP��V"�K��g!٭a�;�s��-����ωT�6��t��.��V�\A��@kb�oX��X��ot&���4@�E:���/���"Q§��)��E[F���Ʃi�Ǖή�X�FO�u'ٔ��0f#]�6�;(*3����,���x�4�lP��|59ۼ4t��vs�BI�󴔯M>ͷ0S��n.���K��t��/{7+z�u �j0c{�5�Ww ���|'bv`��c|�߽�7���G��	 {�=�m�pny���?^�~T�<�T��6`f��~�A[`&�,�	�6�sŁ�O����I���M7Qcg_]����<�~��PS�_]w����KLi�``M�vF��ᳮk��%.�e��C���Ύ."A�qx�s��Y'XV5���wDq��Ytc9V�[�f6rX�����Ua==��Æjd�g��I[�ޛ;�J �`>������Aܷ��D��1�[v=�۷��t���_az��j׫�n����Ͼb�;�;����Y�7����&}/�з�<�!'[ձ:o4C����X�Po]" 9�'�l<~��5��i1��_�H4=�~��r%-�]�2�U�V���;ΘJo�����fO�P���Rd��sɀ��9�W�Ʈ�Z��'�m`����V=��z]l�f�m�����WMY�j [�]���ʿ����)Bܣ�҄�J���^Z������)���'n1	�2�G�|7Sy���Fl�Sf�RwZv�ۤư��'���ֲ9��q�Tt���0��T��1�v��S�aUo��'o��\�ҌddH��r�R���/Iʻ��x�m�!�����˂f�	)�/2�v�Cb�����􍠪[��k7���۶�������Я� �(y���j̜i3C3]�7�&���"U��  �����g��)[pM��ı�ܕs�K:��;>��|���~�b���ѵ�mX|<	� � ����=��x�A�_�&Rc��0��@ËNip�ٖm@k4��j"���Q�D<e��}*8esDz\��/m&:��G��B`�6�)��|�G�ᛩ�m���uV���6��^����yf��x.�("P�_b��o$�������=Q>"6�;���07jTD\��I�P�녏��R�w�)cw�Saζ���@�0��z4��P��w��ViaW�O���ULR��K����W^��gP�P\\ѯ;��Gzpθ�GoX��ض���3�5��a4W[�2��!
i1<��R�Nَ,�Y�dfq�n8��������K�/C/QV�O=�M��*�bq7cI���̺��K(�+�9�[���e�0Q������s\�l��X��������AY	��g>S��f+B�����\Bw�)Z�n�"�fm�8-��(<�g�Dm���e�Mp�.$8�y�k�7(����Lm�U����Ϧ�QّO���]�n���f����uy����Py�n2Y��$�t�
�rq�����P!�J�S��G'C�5�w�U\lY(1(�}�v�Y̡`����;Vm��`�)��h����ٌrU��t.���֤��7-�Їf큂/ޮ�5�)���I�[��.�������V�r�Q��-}G�A�-��m��X��u�O�y��Xz�/��)=�t�G�˴�B�?ʯ�����hڣkE����mku����N�):��R{����-�_<z<2��LT�}TK�6���TD_
ȦeT�8�4�6�K^�țcק*�W�z�C���à�~���=)���q�z��Ⱦ{dą��C��rKT���o���b����2�ËLv@6�1'E��R��P�ܺ�}���c�zF4[��\�7��)�n:B�l맏i���!��g��v���:U-���8�g8ܱEv��s;�!V���Z��lIc2��B�EHI��m��v�<�VBo!\p#�H˕#s�����ުr�M�f���R�D�9M�')��?C_/Yf���Da�	��dU�U�/�����O\����X��(��peoID,���_�#k���c~��a�Y\.��+��F��TA�d��r�Ce(�O���	�2����r�(�u��ϡc��0 ��.�1�֗&�;6�����#�X�C��j�:{�6�{Q��e���+Nݛ��z�υ��V^S�y��6�w�X��m��|�_��<��tKm)�Z����V�Y
9Xǵ�	3�6�F�����$��f���n��9߸�m��~qL�U�n�[�8�3.�775��J5ү{I,�
��R�o[�x�Mn�i֪�尤�]Í����٣\��dI)��o:|��x݇.p}/���.t��:wF�P�1��yd��NV��C�U�r۴��� ~-����h�h�I�R�x� '����=OǮ����6�������Ɛ[���D�x�p��L8K�d{�{�4x������MTG[cwu���^ɮLS>�X�y�)����(;j�N��@ڐ0E��qG�.;×����3����u��a��*��ob�pj��3h}td�t����C�{L��u��DV�{CMO5񍈮b;��f�H��qT����J9q2�����a�q��ˠ	��hʙ���Sn��x#�ak�ń!�-q�HkLV�����^�L	�du"���ϴ���R�����8M�*v��V:5������-@Y�kƨ�ĻV)T�s�u ��R�5X��3)pˮѓp�����վx)�]����/����������t�9�����,�+��+�H�&-6�Y���3z�1s������ܵe%XCL���b(���}{%��u�P���tM�P�2���¹n�cK^�됧n��ӳ}��J&WTyo-����[����ԃ�UN6�L77��N�L�
2&�XZ�Uj��3�����/$�!�\���Τr�oh�����5�w�����<�|���g������||}`�w9wU]ң��+FZȰb��X�P`bG"�ӷ4G��;D���Ǉo2���L&���/�����]��������>�VQ�uNM��
���,��b��pe�[�2jJ�=�$��%n������OVL��Ԏ^@s:�x�Ժ�<J����m�'����$Va�u���b+HW u;�rs���������w��&e�wi�ᝊ*�]�%p�)�%,�fK}��F�D[�6^پM֔��3�;��AeZҢ��vV�j:Ь;��<�!;lL���ͮ=���j��=]��{����E��NT�8�V��z[�α�F�ʪ:����ab�d�e��wJ-=�mP]��V�z*��*}���ɶ�0�ķ�m��n�Ove�+`�N�;���/�{{gL�Ic��ng*JTn��qԽ�� ����ɤ��{�\M-�Q��9������%�XW8*����P��q��a�x3K��vp��v:�L�]s,q�R���[����:8��m!�&E�u�0:�f�=n�&��&[s)r��`RT�U7�޳���qϐzl3�V>���ݖ	���4)���e���-]�5Y�LC���U�Aj�m�ɕ�
W�����N��˽��ڧ��%	�Ioo6�Y�/gh�Z���e���Vt�i��ޡO
�'_\����a�um���v��&��8Թ��!��U�2���}��C�&�+��#�ík����t��Y�q{)q���-���;���o��uI��6dZyYc��=��d���O�g��ww�R;�̺�w���D>i�� �!�\]��R��z��;,�����aiqt��M�/Eή�3lEƱ�.��IL�f���c�Ґ�9u'cF�ͷ�+�>�v�G+�趛��2<w����dX�s�*`�h+e��h��n,Dis��S�V�<������rkй��t��9r��y�u�
���N�;����b8�QHwNa�n,}��4����[%��ϱ<->�8����˧B<��ajn��G�M��M��siq{1	�pFsz�\�7�Cp������35�Vۇ4gŮ�����`��o8),b��v��JGtAV��VY�*H�N{�)Z�J��E����hI-Vn��á�wy7���IitN�a���u��[}{C���*�\��w�d�F�aTﲹ؊���ظj��޽�.�f2֪�.c���|z��R֋����:�G,x�s W)6�2���Ṝ�����T���P�&ac�ty�gQΧ�T�;�p�Ҷz��&�CYR��6s��\gTǡt�in�	K ����rț���θ����e�p䱺�i#���NA5��d�!�ޫ�W��E�vt�xdB�VR���C��pj�%gE�w����{nrm�{_�x>� ������&�ݹ��%����1AX�A`�9̀���|�S6�:��%]�&���Q�X�x�刱m$X7���%�sQK��K���4��4���
�\���s�Ί
���vl����m&�I>v�7.|ob�UҞv��nn���yk�'��y|W/�m��6�x���ƹ��wsw.ذ]��μr�F�5�x
����m�Ѣ/�+�qs�;���wE~~�ןL�}t�.b�uە��u�%x���n��7.�s_;�M���|�u��\��Ƣ.x��C�\��4$��t�^Mx�7,F�\���xs��x�������FBW'@��--�c8*B_YG��ˑ�,�!ثR���e�%�~󬠞d#hW���)l����e6��]<,�������}�{ā���kF�حcm���������d�ef�(�������	�Nl�k�NP�<籛�y�(V�gS�2�:a�[�3�;K%˚)�� ��;9�'��\D͍j��g#7���㊢�c��v!q�g��E�xg2����z�$���9+XY���^���&��P}�;DEge�)�5�!�x��y�P��d���iB�p�O+Şwm@ȗM�]sm3�`�l�y��k�+���m��֣�Z����1�W� 潳��A@��{�ziYP��k8�~��U2H���K�3N�G)��3z�j�5�Z�P�L�ZC��@��a���6�./�y<��&�n�����I��d@0r��Ř�3��A��Fkw�%T��T��לE�\D�v��Ӌ�ڔ8"�G���4!�w��vJ��D�c��n�uO�7q�\H�6j�c�霅�t�Fj�g^=4�`|��;�>���[�|��(Lm�M_�����N!e��2�z������i�3,��n�"1�5���/8M���T>���i1�U��Π5Gхe5��l�U$�yX%#��_��Ap��7��%v�tٴ��uoowj|3�Y5�g�Tuȋ�W�iɝM�e8fVd[h�:�,M��?��x�7<��ӽ)Rݡ4A����T˹n������!�f%��FFz�� }@� �<<H�b�Z�X�4V"�[6�_#��[K������L�S'�0�C��֗RV�wex�p����s\�n�G������Ѽ9�S^�Y^O&�׷���%�,�g*�j^ŵ&� �S�.L�Ά<��^ c=�^(&��Y,Y�e��|��籘��<6�M�T�y���=�@��+ʘ�8�ds�+�&�oK�Q�a��@�m�*�K��J	ڒ�O݌U[��w܉P���q�j��kkI�\!&ŚK��]0�n9ËzsK��3c�	��P����F�>����U��
�c�=)��B��R��8�n�񖈄5駡�vs���a�!v����`�FGjhL�Q! HZTKv�]������v!�V,���}I��Pu����p�A�1�I����T=5�m(������_�ãq�y^@L,Y.ɞ2�j�g�g�s��~L�EC��\0����΍帴���x��w��a�$ó�ox�L8�&��i���`�4݊ tqV��(�q��]f<r��뢣Ӹ�Sk?���3��WC^�ۗR���]��%9x��-I��u�*�M��nn饺z@Rۨ�-W��N��#E��y���њ)�{��\A�{>\2q�,n�`��T����,U��H�u�v��S�y��W=�;�\��Z2ؼO'�t5�}��J5}i�r��a���V��R�GQ��W��cZJѴZ���QF��جZ�m��TmR��Xؤ���g�Ke����%'��)?\�n�M�<�C�2��j��-]�H�a��"3���w��S��zG���k��j��D8�dka14�[K~���o0�F�2�Q��	�g��UK�
��}=[s��9^}�d�j����M����!�$y��./�<ʂ�����j�?P�x�ք�v+咖���X~f����I��i��tF��,t;r�T��I��,b�ڻ:�nL�(3��ê�.ұ=t��k�i��z�:D�w�_����{�DGw|���O=��5��u%���^����kx"�|!�jzxq���x�T-p<zS3C:��Kъ�l�M���ʹ�ڨ��s�,>K>\�W� �C'[콦5�SGF(�DqK]��ub� ©��;.��Oc��{ݏ4����h�mNyt`���(JK�J��M�����y�0�(�US�2��R�oF���g���l5r:ȴ	��ڶ@��,��c���5᷋��kW[	����q���}|b��Gl��Q��eDf犦<*��n�������jC\��O���V�6Ψ	�p~�I�+�|%��sp�
���R��VNe��=K�W;+J�v��К�&������;/��ׇ���匭��z�3rQX�.��=��Ap�\���^e��/�A�=;|@��4��jqj��P���b�'� |�$x� A�4�clm�M5�cQQ[V�{�����y�}{��Os�'
:^p����f���⽝m�6=����)�$�x�"��3ٗ՗�z+z��kR#�T�#��G�R���|h��P�).�<�c�6��{+/�KWR��V�4;��>�H��߁~�-d?�,��v��(�������.��y��<)�9S������h��;Z�J�aR�%�5�"�+5a�:�N��aXc֡mG�c��]����3"�6pü7*w�[�-7����v��X������jNt��J.L���;m��d�Iz��J�t���{�=�b�C��h�o��`���"��|�j6��)]=ҋ�$J����X��s�]��ݟCw�7��7��C�:U	܇+�{�zPkW�w��Y��h�U�<�	���Ч�;�{yE�L<��'H�w�^E���+�q�)z`/F����~}�w��y��@���k�NJ�^�X޽k'�k6��n�@��3�de��"�0UUd�՚��=��`�lyځ>�7�:R�Qn.��K\�;N%+E��gR����W�����R�
	�Bk�ą#Ij��ͽ7S3�P���a�S�7xs-Վp<�̈�<����$�j�ɴ@;��]Г�C �XjPc/x����I�G(WM�Ef�ŻO�\��"�R����U�0�K�[�Yj�[Z4o��3�N��w��ͼ_�?IQV��)-d�T�g���Sn��^u�#�8�SV��8�/+-�,t�u3Tz�� ��⡉xn!��U��9�q�����p�evFD�j��.�As�}Z��箠M�tU�3}P�?�����M��Ԃ�2��f�q�EHSCs����|]ծ^���{c+��RA�ˎ3)���W>[O�~{l�Ȳkĥu�W_J%wai˱�PM#Ѭ�b�8a��9R�m�	l�S��T�g�Hݶ���Y<�'ԿcZ�Q~9���Ù����eGu1�s�~N'4�N'68�͉NP�(�.��sს��w[wsh�T��>���X�������M�xM�'��l2t5Y�\�y:6Ҋ���U'2��&p��3}��C��PU��h�	
$r����6���g�������Tb N�r�W3ݚ"#]e��0���@͘�N�֡�ˬQ�Db��0��� ���C�_-�֦	��}��.ٍ߰T_��r]��̠��Z�{�UR���b�j�AͰ9��@lGy��<1��StQ��]�����A�/�C��u�Ќ֣* ͌*�>�����V8%j�����-׶�R0���UX�k�@�f�.�K�i,�E���R7�
t��7��ǵ[�-}EGRr6���n8'.e��\8��n����Z�&j`lb�S)�`��]3'�˃��V-�,�˃i�˧�#�|A$x����#�$x�|��*h��f7ǧ�P��HR~l
˒_؆�X5���K��*���w-�� Wb�8��P�&e�A��O�Y�KDɝ��9
&�����Xw�ի���:��z/��k�I���۪�g���D��������E1��#~���)߱�,=��]{�d&�^9[�/M���%�Be�������vE2	�l�##[I��;��6ʏ:c�=m�%�*��b;2�=c<s�'6 ٟ���	�n���R/����ve����%�-'7�+�h&�Ĝ�8R��N!6�j�dO��ʬ{�R��-�CV�?�J��5�6-��>��j���]�ybYa����A�L�'���N4p6@lg�#5ߎ��ض�cɾ�y!��M/-�������G�-�o�=0�8vW���@�k1�#U�9։�Y��I���H���S	�Wl˾D)��6p��4Yפ�d�7&r=ys
1$�j+���a�7�8М��O�gV%��˛}�3Uaa�5o#�XL�+���l7y���5�,a ��{�ӗV`b6����y��>��b#����\!�-��Ot��cy��|���F��ae<ق\��9mi�®��Η�}u�K1�5�ݝI�"���޲���l>�]lS��^�}3xv���޳��^���:^V�b��7�c��	��L�QT��}�6�#Ds����@��ݬ�;���tm��w߼�<<��[�`�mb�ϯ�ǟ���AG3�r��Z	3�~fQ���.Z�b��B��+���dBg"�?�)g��M�R͎Or,\�{�7�"�Et���)T=Z���Qj㟖�J��^���{�g}���aZ�-8�ga����.n�&	���=H���4���P���.2�W��ξq{��c`��l�5Cr6��ˈ8o�0��9�s͜���Z��)�y�d2��P���+�8��kfת��8[Q��4V�%y7*��\����m����ְa�ug�[����Xծ,���j��xh,��q���m�\3n�kƨZDZH�L�ZX矩��p�TS6�;�;�PCEժS��Yi�Ј��F�4��w<�
�Cr����~p�
�L�����7�M�S�ù�e�錅O�ǵ׳2��ټ�<�R�����7�X)���}a0{J��u�n�"��Wd��tYT�W<7�`K<��:�d�kL�Ϥ�7����T"آ�!����2 {�ō!Q� i	�g	a�Z�ђ��&��5,k��ip�=1��xԍ�6���
�S;ll�휻�mA����4n*��b��\-��Dӛu�������*��2�L��7��m��!7��hy��HXy6�{�sU����ϋR��;3��-�Y[q�U����s�ŭ̖�V������Q�-`�	�,��H����>�O�G�A��������|b:��l���sғ#��%���ËMO(>��b�� �]3��W�s�l�};��5Y� �1x�j|�Sx-��d�́ATG��L�s�g�Ka9τ^\vj$[5u�1����\ʔh'vQ=KAB��,���'�H�v��m�LP)����o�y������*sP_o���.b&����z?�Awx�=����7s�S�K)��#�1|�=�Ag[17~������
楮�.%1����1��v.3e��\��Fz�K$rۭ�� �r��W���n��Y'5��"~�B)˽F{�[�¦��;ѹO-����q�� n9C"��j��@��艡��6# s,���K�J��4�#H��
���9�"���D�EO5��El��g�ςQz�;����~�l��Z��6sC��LIV�S WϋLyк֊Q��fl}n1C�EEK��Y�{�l�W6l��˕5��
����f��ڣQ��o ����`�<�3���������:׮+�6�Le�v����P�2]��h��� ڪ��&���t�����[]����N��wK<��V-i�Ն��b��g ��F,��T�0����R/ͫ<F:��l��M�kb
x��+��|��m��4�AE��I��d�7X2�]�j�p�$���=Yw8��<C6��oA5�����;��t;�tF�#ot���7F~��}��>���ٻ�V(����Ő�v��c@�g1�
���.;���Z�W(��^�щ�5��T_	��µw�K�p��C����"����i�����(G��I�����wuK�\�*ȷ�-�c
kɂ��Жw�7��>�E�+������5���<�/r���{����)��Y&z"u��O1t��p�yI�:T�/E��}2�%�L6Jv��v�JV���M�+2�b���M5�wK��\+�5\�T��DA��N�>C#��Ns��
�Z�"���qvs^�)�v�M�)LI}{F�/آ�Ի"�j�s�!/����#� ����^��Lsl��y��n�]&��.�N�fuˎ�%��U'�m*����j�4����NH�;OG
g4���d�c�m&K��*Bg]M�Ş��;��C5��L���GQ���v�t�LF�)��6s35��e��3��ᫍJ�&j.�Nb�\b�N��qza^�)�y��J~C<b�pWVlL�>�d:5��J4e�X����8�-��&j9�q�C�j�I�?�8����}���'5�bq��[PF�54Ų���;���w�_i��W}��LR�4V��w�^�(1���a�%t.��q8�b�>�^ʌ�G(n����6&4d8��)11<(.ӛ����hs�����o2"�]�$e@�E.���+���c�J_b��<><A-�^c�o)�IgIf�������
�U��$(��泐�h��0P7����Ɏ4��E[$xu=&�sU��ٽZ�{w�b��K2קV�ڈ7���	���0�Y�\;[�OHOQ�;O��8��*�t=/�������b������UU�k�ׂ+���ͭ߉��׵��v���Q��B�����^����+Z-��T�V*���C΄gٟK�-��3���x�|���}�}3ʢ?-"XVzX��1�f�d��+
���Ic*cv3j�v����V/.n�Nŕp��Z�f����B�!�n
հ�}��og�9`��YC_���w�hw�����	ޔ_ʇF�|�;g�����(Jw�w���6�NL�Ҟ�Wn"�Ҹ�R#٭�����;"��a������%�-�ѐl`���8��R���S!x�>�uu���&��4����Zlcj�T����Uœ�U\�7u�ue��б�R�v���!�T��1�=�M��X����W�]V��8��b��^Bʘ�oD�=�g��x��}��o�������>�~C��侏m�^*�n_nB6Ԁͳ�$��k��1�w�4���#*�
�1m��Na�zֳ�.2�b�˸�0�vʩ���[�0H[&j�[C8U�e���mC��8�x�rV[�����%"x^D����-G�)[���e	a�$М�vc=i�6��1o��F\��f��'cT7�ɿJwK.���C�^i�9��0�P��u��G�u��J:�_%b)�fYvإL8U�ht�
�Q�.�
P�:N�o2�L��K-I��� ��� DLn�S,e;r^��:���50+1Z�L 3F��V٢"<�`!�"�r�cN꾬���:�2�I�Z��8"/oX�AKwk}n��\S�4_o:�]�KΏ�FaG���8[�4�\�횓j�9��au5u�T��^��_L����OdZ���2��VJ�j��I���fʻ�2(��Y�X�Fx,���I�՘�z��}Fe*���gczv��P�n���٣S�=���.Xv�Ԯ���^�n�h��ی1�-J�tPJ�)��.a쎑Q�z2���k]���2�w�J�ЁWLsP� MW�&ep
=m�������4/��	�w �2�a�
�� pS��Z�-fy�R�YY�2>����	(KR�+��B�˥�Dk�yʞ1��68m���F��V3��)n�|���wuJ������Lm�:Z�9z�v�����(����F�8�X�ӑV>�HU��ik���L��f��sD�j�����z�ba.� R�~݈e&�w�^4�8�9�.�k�]]J�۪q�7�����r���ɚGdΏ�e8(��1��+:�/@Ɍ�}j�-^Qȱ^�G���91.gY�]wa�[βɑ�%E3��eWv��=b�CdѤ���.��d6&�/��[��׋{]�ݬ�Ӵ�|��o.uݪ�X���r+�$�����
��o��{	�Ƅ��Gw��qG@��5Kwܨj�����7�[���k�WL[����
7m�{4�ik ԒꃩtPu�ʗ�Ь���y,����zM'4漥��%u@o_:��w/y�%�ЃoV��^]ȵ.7}��U�|Of�p :\<�
���z�ܲB�q�\�\��P[vz1�25/��ފɽ�K����-
�֦��d@[��������'j�]p:UյnF�cfS��oKU[�:r�=�Bx���%�Y5U�����5Vf�W���#$��xU�ـmLA��9�� �op�8or`����U���ίhb&R�3�͋��U��)��QVęe��!���=B������A}Co'` Ц�<�v�[X)!��\<�0����<�E�M�f^Dr��*���'G���g.H��FFe�z��9��Dv���YkH�]�JǸ�i��)m'��B�j-��h�zp�)��Xt4c5��3��V�2�;7yԋ���G�u��}՝��܌������AL� NC�wq���#�/��؍K����$��H�yܷ<����/�<�ݹ�wZ�Z����_���;k�>/��6wQ�+p���I�_>y_����7.�yv���澾|�\�����W+�����ֹ���ss9���b�\�|�������睝�w�/-yݳ���WŊ�n��⼚��9�⹣;���s�<���i�o�s��;���5��s\���}|���4wls��vܯ�`�J�9Į�0��'Ƽ^N|����+��o�t�m�םĚ�;��<�%�x6.U��sO;x�b���������v�Z�;c���O��>7��%���u乍�Er㳑(��(ƾ�/�5�\�s���^�$(�}���� `Rz��y��9Xa�ȶ�qctM�iG;a	9{�M��N�m�{�6b)�*({uB�4�m��7ָLo/lI�Je�^]��)�A}��*t�v}"}e�b&-��e�T�0�XL�ˑ�6��q�O�<US�M���z=�׹��P7��w�#�Zi�D�+�&���]�;=�O�A�͘
����T�r�!b�D�9����ʽҨgk�,{�ƭ��̜�Ce�ͺ�2�)Ғ���l�]0�<3�+�\/�/~�����g���l3����DQ�ͦ9������*ÉX�. )������md���cͫz�7�sm}�P��]!�5�S�R�����Z�v4�1z�"�n�mo�T��^p�:��<3z��6���R���G[
U­Ch1EF�?-�S�kԇ��÷o�"�����X����y^�N7jbش�cf��"L�s�,��Ҫ-W��ν�N�VE�z�ڊyA��A��p�p�	�07bp_j�J9,�h,ǞU�ީ+���#���7/�'#B�{x��r����py��h���a���)n���*��~+`��*~t�Jm�,O�^e@ZDZH�L��ib�M��	�m��dK���F[��Ր߆WAg��E+�z�P!~�SP,�Wy���ٕ��y��==�V.,e)=�ۛ���o�缘B��kT����Sr=W�v���ƬFD�NW8[�����k!�s2A�gf��ձv[���z�[HA-B��+�n���/{���k����e[�8iߘ���ۥĎ�AV�Cr��Ҳ�I�9S�c�,��ij�Pٷ]�k''Q����jGY=������ބ[s���PD�,nWP�p�#Wn��9�4���bجm:�j�+a�f�Ψy#�}���Z����6�����{���{�����~��#�m\D&"���e�d4�@lҮj\gҲW�GS9�P�8��T�t�t��_`&y�����ٱcPJe8[.*6BFy5鎸��i[�,�]�n҆��<U�#�y���J���2��:��S�1J�F>7�F���cǸ�����<Ζ� �MY�[��޽.���� �d�^t �4����
#�.�9�$Y��zum�)���[݇�{Jvq�&���z��'�wWƃ��⨽��2*-DQ��*��#V�e+���;p�v�&��m����|f��n ��ȇ/-}�(=6r�~5�P�r趎�|�$vؘ=��jv�ک���{(9 '	��Gt���¤Jn����)j{�5���E�FN|<&Oeg¼�Mk5웿Q�D�7�����y����Ķ1��U���ut])7h:�Fm�k�jNQ�z3�So!T���R��S��R����:ә5�C�v�{܇"�No����l�I�rһD�.N{7���g3� jFw)�N=s�$)궖�,�`]��$Dt�6�=U��Ia?{���@D>~��X�C���Q�O��H�i��� f�Jv�i(�$�;�U=���Ћ�ǌ�Lf�a��RW�`F�8f�Xl(���s`���5��]��\8󽍫�M�ϊp���$i��t0�S8;�[<Dp�M9W�Uϧ����\�p��h�|iL^��#��ػ���?�6{��f�E�B�H��3��[z:}+^*��pl��w�V���p���D#G�-��3^��5�x��0�/�Lb)��tA1R��u����Ƙ� 3�11E���&���	����1�4.��B.&S����4v��|���Q&ގ�OS�E@��}1-tO�Y��z}��RT��U�h�;Jrc���1oFb�]mvuwNN�����4=�\�%ҁ���ڗf]ҏk���5�Jw��(P�!E�ϡ��n�w����	�BgDU��6�VSV�*�jz[� Ku2=�Q�+ey��x��ݫ77�f�`6C��\�gh�� ^Y8���}r��j�;r՛�7=��շ����SBޏ���{n��Χ�/"$��d2��Z[�ù���H�؃W�ݓ,����;��_]���[2�U�%���|��S*���*+�2��kx�ٍ�&�EԨ�溾ۊ��0��N�̋oAy�*-�������#�6�ʜ.���r�vQ&��7'au�O��V�ب�u�PJ�XGdY㭨9}~12��*|�ߒ�l�}���mk(���iUc2� ����*ni������3<�h�u@&9�!d���5�7�ݫ ֙D,d"����
y�J����G�G�G��;�_1��ϣ�nz?����2�~эbP�Y/,&ɤ�\jS�&�&�	��XVUv,|���i����dy;(
کG���@t�r<�8�-�3�4�\lk�V*'5R��%���rQ���'��wk�j��C������h��B���[�f��x�G���?t���74frc�[]���H ������fZ���x�L,1XA&�-%����5
�#/;�N�V)�(��)��u�3q8����.!�)L���ǎC���m��f��j��&+0�yZ.
��������:AI�}ck[w��~3�©y�ڤ*�����������[a�_�9�5��G��C�֨tyYAQ��e��EX�#J�'7�ƾ�M�R^�=�����v�����ɕ����k�?=j�O���B&Y�/NQ�@��������
�;��)��C��w�#ea��u���V6ڀ�:J�ds�#��.�dDu�utg�Wt&+N�aHŨ�k2��6	[��ɑ��׽zx7(m���H�7�z�f'��\�Ĩ�vtͭ�yhq�>R��iMRF6�R@���Z7u�n{�- ��Ϥ�56%6��ܦ���:<����iʷ�C���Sj��%T�GZ�E�Clp��2\ȵ���Ǘ�ip��L�y�B���H�c9�*�IWS�XEuP�_,~Ψ�&��/SS4꫺ ّ����<���T��Y4� WT3'%G�fp�v�}�A�(�b�+�̴��Qp��0ͫg����cל�H�x=s�}p7��N�u��4Y�1�v��s�s2�IQД�$ �%�\J�u�u0S�~	O{t1l"O�-4��=� ������E�CS^@U�1��nC�L2u�4}���Ԁ��R�]�cnwL��RF�/j�O��i�����'�������0?}��/�h�d�4�*�e\��6��h��L��w����eHkި���R�s�4�mb�c�W�C3r��1�k�F\�˶b����7D:W�l?��NSE7\��������-v(8oV$��A�U��-�F�{��퉇���KD$���z�	�9Y�����c�Bֳ�5��j��#m��+oMmnv�U2{�LDQ�\�/���N���J{�D�Z�#��/��	֨�1־*<�n����[�.��X�3^��p �X6I(}���*�,;:��xw�o�y!y1��LV�m��9m�:W�ʇ�6��f�N���C:U�|U���f����>ϭ��ż�@m�t���C�.�yd]�t���A~��^�/H��_�����r3��A�4:�sza��� ��fX,�	���v��8�U�6�9��ʲ��%�O �p��TgF�jm���^<�%��)�My��Yi�������i+�a�5M��%���Ve�<��[f��gj�&����t�QiW�rmx�u8(���Π�8�??_��u��9&�@����~��澀S=[��{�y���ͷG <�.8����Q�ܫ�c����iyt��b�/���Q���PRc���Yy>/��P��ʃ�2R���畼�>5!v��'��Ꝏ����/��D}Mw/�1F~v��R�,���k݆	�%�E1Y4�v�z}�w�����Fn���>����Ċ���ɹI��{����0��/��5<�8��stY����޽`�@���{�Fv3׷n}�Qfg��l����>j5 �8������]-�7,ݝ<���dr�`��-�+�%�H.��ͫ!��1Sx.ʜ}�Y�]h�D� [�O�xxad��<�XhU���H&'0`�Gg*�-5�t���J��)2�0��v��uQ��s'�L���}W`����[I���Z��9Ժ��b���
��D��:�Y�5���'�bZ�6�ܽ����
h�G�ݼ,q�%��/>����"�����\�31��A��l봰�$����aQhq�.���4��ݧjQ�ި�SQ�mr{5wU<�QV��*\SY�,�1ռ4���N��/lb	"�J�<)�,��eN$�Ӹ��.P����U��O��,؆C�۪���&<^/����������.�h�<�oc�<NVsK=�"�5n��2|7�Đ<G��O�TS��ڶ��V(iy�2`Y�O>C�:&^�	8�=ͱ�9
��a^�YҘO�k=x�i�EzD�D]
�1�i�u��CUR�{�9�:)]u��Il�W�k�Ns>���X&���Kl-�pu��Ԇ�0�p.;oQԦyW��^%lsǛ�
��r{S6�Z�֐[Tj �d��o7y=T���g�]����mj�ެ��o[j�`�P����E@m��+΄~U�%��e�Ǐ��'Y���\��,Sw(p��Ǯ�����o,���;a �YҨ]ᝉ�DF�pPגo�UF'׮rԸrt�`&h�0i}{!���s��^ɪgs"��J���i7�������fU_f���O%*�J�C�{N��C�.s��;�5�T����1��7$�Ԇѡ��b�#H4��0������AQ$z�ݘ�Z��
��r�&W[��F�h��/D�rpT���
��-!��,T_!�m˶�p;�me�+oc�rs��f�5�tWQ��2�$z	�0�e��qx�6y��z3ʣ��ߋ�^��%��^m�6��Q�!�[u���k*�A�]<�Fk�5��������D�{�l}Sw�c.�Z�N�*�%2�sz*�J�#����jA�,�EZ�Cm��j�nU����"�T�QA/�����ܱϲ��sY�&��!��0��n_^���u��1e�VotU�3��!����1R�KfZ�c�������Z_:�8~m%�:0і�4^���#q����kl=�w-�.m��Ҋ݅��*�q��pњ�R��A�N4����ts��ںG&�<:{u��Mj�xe����h�怽+��TYh��`�A(����$(_���)�cA�|$ùy����vG]�E����/ژG>K+S2�0���� M��?�4>=帧+b����t�y����nӦ�L�6�]�.�f�D�Z����(�d������L�כ�Y7v�e�tގ���l�r�B��d�#��
���GYvV�Qf[�'����/����ď��T�g.{4��d_ݮj�8��u�@����R79�m{��%s�yc~{w~Y��"��K[��*m�f�8�za��qpt[zx�InIڴ..��\X�M�"�k=36����n�|��*�'@���Ѭ�l�pT�f�\��ʫU�A=�m��;�b��q�24����m�T��Mj9�וU>�o;Ud��k���f- �pL���p�l!�frYΝ�D#�N5�"��Tb��qƫ�)��C���_ٗ�T��N�$����Es�V��&5����N��$9S�N!�VY�m�f"��k#"sDG�7^0�wq�64�e8��[~f���z/9�P��}�6��9p26�r�N���[de��G4X��}�n�v�Q=���ܠc����w���li/�*TLw"��z�*���B�0�*8�wX��n:�p5�X4u���;f���g5o�U���/\_쵅Z�\0��+��ѱ����S5cz�E)�\D
�e��T\�'QO�K#��+<��8�4# �k�����_���1�L�k��G�imme2%g%;_xPj�Љڈ�p���ɖY�O=n61���gD9�ei���^+
��b+;"�:92�|�wD��N�&�G(����F��q�QKA��p�����4��8�����Q0⒏ �WO����VqC��2���~���f���w.L�g�_�)��CI��=�0*���4Y3�Qљ���7�5K����%b�s]���Aa59����oP������P�X�7J��B	�o$�h���'CG���~d��7S�P A������O�D������:a����B���~�#����=G�_*��ũ�T�����-=0��c$���\��C_P� ��gM*���^ےp��8�s��x7c��u��Y�8!��PK_)����r�B�f���`�xBK����g^�3��s�No���^�p鸇�3a����uͥ�aJ���,���!)��S;��7=�zb��F<�k��&��a`��c��[5@t���cr�w�&�]saS;����(�8#�G0�|�\�X�A�G���8u!fk���v�tqV���5f@��uu�\�L�����鯟������F�����p��=��Yi��^����_?�� ���6ߵw��]��'L�OZ|�*b\ƻs�1�{�P����@���u���Ř�˃�4��KL��ߦ�0}O��)�a�~]�x��οT�m(i�t������<���&��qD��ߧ�~�0����~�=�;�K.������#w���JK>�2��P����������^^�_������~�o��g�x��b̺a�#��AD�S�3�|���Ν�=dޓD��3�jؤ�����A���)|r�
�r9qԊ�dhmhe���j��&�ཕ�-).a{l>x��q]=��uw��RH3�T0_'�q��yI8���;tL���"U�P�N�$31,�s4�+��㬫����m�2�_.��$�N���T��(�m�F�o[��.�$c�(�67G4�� ���.�-T���*���E�T��N2���/��L=�ݔ;����#+q�w�en�Wdns�(����f�k^&{���nE/B�;:r���i9�1�7����pqРAiD����{������ѩ�k��"�$�XM,�}a��ÑKI��Z\���h}ծ��9�[O+\A]�w¯��;mkƵD�w���X@Dٛ�3��/S��Г$��w"G�Ǡh�Y�K�˄��\�����;3,���VC06-�f)�Q^��R6�֜�f-�5<��J���L�Ѕ_C�1<�ell�4�/m}��ɺ�Ot�ZU�3z�Kv�	{��"�)[���Ց���˫K�&�C�,��ח����N�KoZ���M�"�`��i#��s+�b�8����9�1��u2�Y!�{�� �P�E���C��\���Gc�ޞX���;T��*(��Afj[���]f,�!ѱ�h��ve�oQщ�f�4UwXD]#ϫK��mj	�[��y���J2��۲��R�Qh6f��h���ow�glL�
�ݶ��}��[1��pي��Մ����v�`�nb��f�Xqiq���qYR��nL��b$LT�Ќ&qdvY}���*�ĉ�wz�rZ�*.�	͏Vuˎ�C��@�KY6�Ի6O=�8U�-��
�9���>C���v�|TO�,��Ź�^�n�vTU5I�M�Y�p5^Ë��fbtf^�Y�J�6�p�K�����|�p�su�ɽ�n �-��
*o��o������wk����[�Q���t��&�[ �[k�Y��q*|J��L�)��o�mung����m5ϙ�=��'�jң,�w
�9ާǥ[�*��ͱ\��Ջ��户Cu����Q�GD�{E'ŋ]���i��$��F��5ʂ�J�L_D�e�wA�:yV>7Fd�Uv�mn�Xf�{�@Br���Y��F�h��W.�cࣶG j�7q%��[�+2��� R�v���S�W���Y�3Y��t��9�ib<vԳ����}w��<�e5�V�2���o^�I*�������Y��Y�ID����2�F�[Q���6m��OQ̅�|��X*���P��ǎ��j���"��kb�W{:VΥW��Ÿh�ÕU�ˎK\��cr� 2�3�}y���L�z�����n76prggaQwge�^tR1D
>#��>$�|��w�����&nr�α�g�s�>y_K�\�t]�y���w<�G1�<䋗��;s�Ⳝn�d��sκ/<��0c���+��wqC%o��<t�s;��y�eӻ�9^w"u��R0��`�;x�ӡ�iB`�<��w4owc�2K����Ǐ����KwW0o<W�+�s�.U˚2bF0�&�\����	;�s���k���҃s�H�<t�k�|t��w��t�c+���:���"L��J	�����3F<�!"a�
��r�Dʚ2$o�k��ӝQ����J�w�����?k���I��n4��s�U�p��Pmá7�ep����s�jn#�Ym�㛇i�Me��ԅ܊ܞ|��*Kt��X�jqa�Q�v�j[j����%܃5�jq��c�P3oC����>%�Eb�f�b���y�Ru��c�N �!�)MKp�nt�(L�V��[6�ݮg�ot�Ĝ5^�w5z�L�sӦ6��t���aT�3�q[S�M3����d�f�Վ�˒�4:�@��W��gN�N�EZ�Ri�JG�o!�Д�ؓGU�x�L;��̓�R�%��9�cp-�5�אe�!O~J,�X˩���[�������oX���e���N=T>n��6u�������D�7������ޒ��2*+�WEK���;��=��f�y\���Ƿ�M�,Ԇæ�P�����q��x�Ζ3�ݫ��z�X�G	��d�]F�3''Fَ��GtR81���z���|��������S�0pT�M
��l�f�
�<�z;KJ��~=z��:�9�5�Fݚ�`�s��q���+��L*y=ؚ���M-:Pڱi�T���O8"��υ�)�}���W�#k)���S{X��^>X�����	���t+7��nC�l�&��+�����F����+s0��G�9m�v��.�^�;[��B���m�ys�vh������R���c�y�3t�](u蠇d�f��Sb�x����#��h�N:H��|��3�L��`���{�
u8"��U�m6�"Z3���Ό���6=Z�a�Ҧ���;	���<I''�>�[���.S�������ǩ`���)n�m�M��r0j�Y������׍B ր�Q�*�C����z[���WɃ��e�_��wN�NM}��8��NH:թd=��[[�W8WZ����u="�DSƪ�ߊU��	��#��|���^,���kz���KS���w䢵��l�����b�5�@��gd��N�����H�O^��'����Cm�c^��&�t�:�D��&~�0��,�n �f������G��j�3�!����N���X-�I��� �S�nPpSvB�@�h�r7�\�E:��-��Ƕ�-f렊j9�[m]��5��,���`|���fQ�N]O?tO��'f<,�#ܦ�IVhk���7ьI�9(��<���p-g�7��=�
�m%����ߨ�=�L$6ي�"VԷ��	MGL<�)��=��.e1L��Ȧ��5<��KN�}Q��&ri�Y3�P����=fbQ
~_�O�h;�׾��u��&����X����a��Ӳ�۾��5��9�顟<e���G_��,�)��͆�L��n���IH�;�ި�͝�жͰ�(޸h�i�9;��4ܘ�Ngvp�s兲A\�����N��Q�ͥ[4ocȃ���Z�*�!�r�D�t��nǶ'6�d�m�(yxוޘ�ǹT^�PT�1y�4�˧��B��7�w�F`uK��]J~�*S���T׀��`����!?SL2~"�.Ĵ�Fݽl�V�z����u�����0�ڮv(�}I��v�-eY���LB�c�gt/L�UC���٭"p�u3���u��T`6��{�y����0u�쿵o6ͺ�)�8��=<UP����E�Q���3��E:�4wQSq8���"����B}Tt�h_n������[���I�\V5k
� ��'��
�䳞;s�������c���Z�UrY�_iK��\��ǵ�;�	�X�%k<�96g���I�`v���i��5�:_��/�`��,�/J�4�t���*��b���꼢\h5�|2�-*p��i���鱅�l�c�Oe�R�r��i"����D�5��.4?s����[����@�m���2�NM�;�;hf�4��0���t�P�z��2)i�]ˁ����WV@a(�nɈx1��AZ�gEB�H^ǰu��=����)�cI�з�b��Pt8��s{�WB�r������cHI�8<��s� �������Ϛ>�0��0��<�L���O�ܭ'7�KØ�����v5ie�,���䑸z��U��J�L[�h�/z�DĴ�����ŝ�z�i'�s�8<��d>�t8�39�]�ކ�����JE��7�2���؆�G�����kl{�f\5BT])2]n��G9Q#X�/�r�ߙ�C�idӭs]������V�����7+�k�ܩ��Ѹ���2`2�Jc��AoLu���g�"*Nc�\́\�P�x��_���ؑ�u��أ�P�C�4㰉�]-*7���y�q\)�z�(���ab(��{�^�;*�S���O+$ #Av�%R�{��~��pn�Q�N�)&;�#g����s�OM��s�t1ǅ���yᅮ4�kf1J��){��^*V{�aĎ����Α�S�K�Z��V>�޹�M�#��4�rdK�k�A�7Ċh�qU�[2�$.�Q-�)�E��-�������Z�= �j+�0�e,Ch��2\o"�8���/�)�-jA�*9�
i&zh��m�*d*��RU�����3�1��@�҆�]�(����/�,��z��|��=��r���|�j|��ſ�W�S?g�2���ad�Pl7j���Tz�r����"�	v�\.UФM�1���7T��J�Ŏ�l.���U��Ws��4�*�>$쾐��u]]ԏ�X0:d}rg�byj�gj�	1k�][��5�E�������c,�Y-rb3�m+Q4X)�}�7���$Ե2�\�j<wd��MI+�s���<�sV����JȝyG<b��-{���s
���ӽP�Ƽ���:���@�硢����څ[�G���`�CG�c�ڜc��l�XթFn@����M-i�[G:�'<~�7sSzeR��K��y�X��I��V�E"kr�9�N��:�M��ć�<��x��F,Z�YB�z�-���� s���CϤ�"��}��ت��s"�\�q��@�tD���O�|!s6ܢ�'.�*�NK��B[B�qߋ��$�?��ҫ�L+�ߋ���뉷n��k��e�v����32Uk[^���N�q�a �޷-g[d|3��pT��vs
��ʣ����G��SuӉ�x���t�3�?T-��d�r�ã7� �oTY��l���{�3'e�W�L��+Κa�V��Ӥ���M���-�;%ڎ���#;������M��L���dz ���qOq��o���bXx�tr*�AqZ�E,��B�ԭ	
@�]M}V�ݵ蜜�����	�Y\�툭����� �L$��禞�C��1�/z���o%E�̲*1
#6تc�>���������Z,��u�`����jD�����8ʮ�ʻ��dkV|&���K	�|��Ϊ���ʲ��umMT�p[EXK�Y�]�Of�ψ8��b8�* ���9nX�x��"b8�K��Ҿ�`v<�(TΏ"Z��g�����l�v���d/�8�8�M���:�1g0���HlMءւ ��1u��(��q�D+�[��u�>��w�VfWJ]�n�ƣ��r4�Đ6E]n6 �¤Jf8e�W�(l5� ��q�R�g�`3�Am����FK��1??���W<IKA��� >�e�����:��+���맣v�>n.��R����<FZ�:�z�KFsF��)+ρXᚉ�ؚ�:�Fp��F_)Ȋ�e'�5��)	f��W�&qҌ��-�Zz"�j��M���!x��kna��7D\��`�]#�X�/�<�]-�O�z��e�%��,b�JFc��g+vq��D'Һ��eu0�}�C��㽔���ug���kK iԠ��{�S��Q��������ш����H��l��1 �L"8������T��
���kޞ��k��aC��I�4����S���ˠcx�2.��뉀��ɋ�m�[Omѝ���6Tpۨ�_��_�v:�L�Bg�F�.��3�́>칈���yk>���"7�;�o�����Kv��9v�Lz՜�ެc���פ��]t�̗�ː�ۺ֫�Z�ci�p�H�bü�wg;��Vo0j�S*ܔɴ)Q�w��u���'��&*W47����Ȳ�����җp�	De�j�
�J&{s6s�`{}.���W�];$��`�v�gR)�j)�+)�oܫ���&X�R��Y�}�(�˰\e7jY��&��T`�-�S����^���1	C9��?��Ҭ�֪�7�����2��[X����Zz>�%Q��PaIV����:M�12�jQ�}�N	I���]�;����;o6�I^Su���</G �_�X5�:����h-9�	^s��S��\l��|]��WG��F�������2._^}E�z1��(	���1=�h9�ħ���IV�f��ؑغ*O�֫����NP�(�.�:�P�4�(�$dW��!?Y���V�J���=5|�ni5>hGb��P�\��cf�W;�}=��a��
�V��$(�u��CZ����ͻ�\r������apWP��p���n*��������Ғ�+^]ZU��U�f����JŴ
��1�5gy�``V�I圥ݯV�s�ՙ:}#ue6YS����\��Z�6����q:�t�<;ZJդ��i���f�Nm���*��K��:0ƶ�������iv��j�B3���\~q��Q���-�	�ݔ�����p����yN��uŋA}�=wfV����H�㾊�D�i���U-E�#���֞��jq�6uM�A�Z�wn����P=��d����'�s��m�,__[�U��fu��E,�l��bɛJ�M�D?��ˮ[�����?�{X(�OT����;�?4u5��o^ydF~�#�E�����;�k6;��*��Ȟ�]�]�|��G�Xa.;�0ǵ��.���Z�A����>��ܭ1b���b
�VF�g�/*:1p�u�c�.�9)R�����C�<��Y��N^���K�mB�M��Ƽ"8 X�b.���zj,�c۬�ʧ��	�	b�3�E�=v<�
�fMI�BI��3�V�M����N��� ,�x��B!ƥIG�j�}{�-)�d�}����B)��i�����X������BT_�I��.ד�AS�oG��=������<�=l�T0����܍
�3�f�� �11S��;f�L�W\3'�I_$j�y(2_̷Q�RŞ.��9$5��S�gN���\Ӳ��-�N�)�Z8��}�Yu��
��Ƽ����"�]��8�)v�\ݩ*o��j�b�~]�MT��̋"P.ԕJ~�b��K&��O�^�Q��Iw�f�Y�A��]^3j������O�����7�D�y�g���4CS�\�x�͑��s��?R�#��3>Ok1�#Dn�D9jO#жMw���<j��N�Tʹ�;������ŗ2�i{��Ѥ��m�(Eۨ'wu�%6������M�C��jz��� u��s����#��4;{��������䅱�5�\k}�%vm"�~�����5һ�t9�}Y�b�XW��-�Uib	�)n�z/�%�N�]r܍��4���-I3�`�}�z�|D����]Hv\߯�J���ц[���닑ѩ\I7�2����t|g�i����	]�AC��9f�t��ç6]��$���:����U�eTg��5�����1t'>�^w��Uf;L�;���l3,k��6ݪ����ulh�z9�ڱ�I���v����,��@Uf��J�;�)������r�LVR��
c��FB��/�!S=_g�����8��TM+�큐�qg��X�	�����~O��DO��9޺,�>�w����4c�Y�g��ǝ`>�aЭֆ�&�c.A-�ͨG���K�VHa�1��X��++{9��!!a����-��0r��Lx}�O�^fU1�w�l"����m���П���o͚Ir"�)�ˇmU����=�H9�����{%�o;���y�h�{�wph�}Y���JlO0�>�nY4���n|��%~X�b��C�r1�O����e��˄w
�z�gLc#��	-e��TM�꬯��kv���i?�^ޞ�]��Gi�� �2�!ǋ��R��h�FG!Ea�:6��Y7��MF��t��9��4�j���
q�4��n��sZ������UL�Xݻ��9 GR����܅�ڷ���	[{�mU	�a��AgNmD�|�%Cnc�?�m��9ݜ����\6E,Ԗ\�[��b3;�����3��1�S
/�ݖ5�i��[��@�l4���нjS��+6R�a(�9��ez;��B��Q�}��,�|���r�C
g�#�)��7KV�R�v�WS�N�yڦ)֙�fnR��m�R�5�z�kW[Ij�dd�F3��Y�g6��4��/�-Kє�#�c�p��A7#���;[Ś��t݊�h8cԘ�FYgb��t3�5��Sd����3rU܄pYp<�{c���n;��l�8�b��'����1@q(q�����*�"@��
�)�v��M��⮑yP_�(�u��1>��p��f�ZX�|"<�Ѫ-�1�,:����0b�Z��5
Bc����;m�pT���g3��m������R7�oi�.��ꓣ�s������j/����͠�u�����c�{*�؋Q�֐[S��W��Hf8*^��c�H8y"f�|�zi`����M�8��7_��P`�^{�>>�O�������}��w������P������z��m��G��F��80�0�i�:�bMsE��̬�ʋT:oMY������#�h�u�u�26Ϊ:ɇvj��ԓ_��m��:��b�f��owa���j���4x����m�0�n콏��B��pJSt*�f���;��G{{�c�u�36�Գ����5lʶ`�W#`�=�Ռ\��X�V�^>�Beب�bҏU�����/n���Ŭ��c6F���b[�=F�G�&�V�@���^^��U8��I���/�3E2\��Ky����l>WB�bgh��*F:�?� �X��Y�&jF�N�A�߈a����6z<�,i�FS��/9n��ͳnk[�\�k��"�S�ɜ�ʹk�L㬨���%����@�P5$�M��Z(%�>v��D����]����pz�S[�P��Σ�x�����U;���q<M�C����8k�+`��
Ep�uяT��cAт���Jk���˕=P|H�LR;��ֽ̅�{x8X��{�OE��^<\���Y����Ofd4��)�ef��vO�Nخ�ij��7�kU�/v��Tђ �i��D7W�\�f����Y.m�k�)���a��w��P)��FwD7eI}���:��p���udVՅ����[����Q���C+[��U��7쉚gU\�ݝ��ZB�R�hnvf�\؅"@^ڸ�!�t��m�4M���ᆂ���哶x�Tͪ����ٿsX���}�}��YD�]ݧb^)}l��E��9)Ϭ�כ � G]��5���S��̥���h��v�WiHnF�N��P&�:o2޻G���I�����;�䖱�z�[.A>"@y����{
�ɝ�,a�kB�,N�B�͕+0[�Z5��Ln�{�#M�Zv�Y:��$w�@&��h#���^���(���w�Wa��o��ue���R�\�_tR�SnJ��o6�gk�DK����f��[�k"yvw���]YBn�Ks��메�㖜`<�.1|���r�`�Y�:�mbse���ݪ�@�:���}.��ZVS�=�=���+�N�ݭ駑o5hT�r QՎ횗QB��d�x�x�U�;$u�Բ�Xy��gM�����[�uғ�kK7�6�f�,�r��|r���bڂ��UF������[s-�{qt�}xo��0�͹'*�f�۱��+ȅ��:�d���@"���Kv5-%+������5Ƈl�v0!],,��md�+ �����7y^���%��)��C; ۳�4�աҟ��"޺��n�mt�U�� r���oka�t*utV.�u`Ĕ�o�T�4^�E�]CySa�Ω(����%��(���$�����0�2�tk��h:᪥�5)�*�-�&T\� KS�mU�%s�E�����ط��h��L��uo^���'ziT���:�'s��mq'%�{{{�� �k��+k3�Z�ѽ��f��2{d]z�{�����iș�FӯɄ'�JL��s�ڂ%�ҟ��[_.����(�4)<�#t˷#�~;���;ˆ�]ۓwn\�5�q&�&A%!p�$�(����;��rL���끔�F	�v�����B�F���#s���C0a#/:�9n��\w�W��342�����/����ݍyu��ɔ���dR B)�������뫉RG��E1��^8�����;LMn\K�;�����u�(��s痁�#&I�����w	;�����#2(�IF����d��d#W8 h.�q�N���F�(1�˛�I���������t�h�s�u�ۻ�(�'�����^w.\�8�I�S�� !F2A❻��\�\�%�01JJQ������
�7����}>y�������o��bA3�SH�fb+qmv���vb�
WJ4��[�:�5���}���Uq���,��	QZ�{��7K-"QW>�!���Gʆ�����`��*����]�6v=v�n�5�p�GAb� ��h��l��GA��4<���%������@��cl�P��ӂ�}+�íL�K_Cךa�()�;�q���J�O)�
��Ϫ&�fZ�$���� �OL��6��S��W�0yUH�	��(&t�4=�.��'�́,�P0����O��^6�[L����Wn��}�l�aR*6���M�V�Z+�:�^��#���N��B(�3�ݙ	�P�^R;�∞�z��;-s˜��j8�.W�&I����j����B|zn0��x���[�׬���K�억�k!l�ٵC�29���|�φɊ2�����&#:,��w��>	��ɪ�ا�zR��`ڬ����x�^&�4����f)����bJ�ʓ�����@J��	�bs]����\�{��1��y��B!m��~Њ�O��֎X����;F,�*�Q�c>uǱC�1�M&��C�x��5�v�(kJ���tM��5ێ�h|��16�;��ߝ2&mC)�G���m�;�r�IP���.k��m�j䵰&��3�']��-4šW2[�{����%��N�fnX*op��<��w-�Na!9�kU�%�z����N��}*Ű��S
���U�Zhq����)y����ECW�Q��l7[Ż��֘2�m�4��-�մ��*p;�g^��OA�NK�A/���NxS`�֓�U_0�f�s��FK�&'���yq����19�9֤�;Nlp�xi5�	�ɍv�[>��7���]�����P"��|��b�;���qU��ꗂ8"�L������	�2Ak��r��y��q���9 {E�犒25��΂d���;��[ݝ )*��Q�ꂹ^�k���e��86�h�c����{r~�<fL�Hs�V=������*��M�ݍf�k�J����B3��;�?4u1�>��<��a���'�e���J/cX��Ǎ�:�x�XN f��\wDq�hr.�g*��f���pѩ��g5H����Y]`�;�����J��+����Ff��%���5�@����ܱ��ѹ$+�`�b�K��=��tZ�8Y��<�Ӳ�)Q���r������H�p��)�YS�F��>[��(r��2�_*#�����%@M_�pO�oдk)�?ߒv��^Y,�s��O�`�n�������_��a��ge6�İ�J͘},�7S����ȟޅ6���*�[��u�]!��]���ӭ<�v�m)���^b�����u]^�!|�K�7�+h?��qg�P=��1+����;�֑{�l���lʞ��3,mr��3&Ǽ���U�5�۔�uǘ�l42��0.��9��+����z�}�pS{�o7z#R����'�6�����7�e�Nv�ֿ��������)4�b&eZPd��TH��A�FMř�M�⭴���!1V�k���qUNP8˦�i�]c��W��0�m���8u^4酫L�n�a�I�]��Ş�aMi@��S��W�W�o͝'A��~�$4�-G���ů��jʛdp��m9�K	��@�~�#��шa��5�ts�x�Z9�o#a�����8yB/��Z�*<S{���Y��6����A�7Ċh�n*�Q�mR�Pz�(����C?num-,5E�m�+m�6����DTA��}0bo{�����I��ɽ������,O�e4�Ka@/��0��{Xx�X���\'�y@r�x4P�n;6�72\��#OB��:൯�c��R\ez�y޹L��q{��x�Ɠ�{��-���u�����]=����S��� 3L�?sDR\gݎ(N�P����{6`��������Ml�]�,�Z����y�G2ͦ��{eN�-���ծ(ِ��)�$8��x�E�?�����,�[�}ɟ�G�"F�E�H��fq����z��'R8(n�
B�:�E�V�=�7�UF���Ƨ[��{��W1�j]�J54�t\�uK�;��t~2��t6�a���:�ǝО���r]��7[w��n�b����dL=� �X�6Mڷx�u3�=?�2u�|Y�Od�dg�vC#[.���'h���K�r��;�Fdv��;��s�5�,��&4��a/_����^/�o�1�{ȍ���>Z e�_�}�7u�4Ѕ0�����DYV�4 l:唡�u���e�4����U\M�^��N�YW�ا�7v\����a����}�d���vџ;m�ʒ�*f(�����(��;=��Q�4(���5pl������9�m�mU����sƤgTA�2-�-���<�J��Y���%OF�_)k��Hp7:��m2�Rf�f*+��]�O�v@�|� O^�z8�����c;s<V���v���[�o4%&���Sc<5�v~P�ni3J΍d���Z��ޝ�P��i�%{UX�\t������{���@5�J�G������|(��y*.@dTLu�6�T������AV��ƙp�K)��C��n���H�
�{���~�_����٦��9��˔A�B=ˢ����c�_�l�01�!f �fǛϐ�yMMW_��O����O_s�*D��PW
�4�i̓;rax�ڍ��]�w�&�߽\�^�o�hy+t&��l���p.��T�38z�6<�ǽ�x@o���>Tm���<��C]��{Mu[��W�S�du�)�� ��k��u_K�8�,�<$~�z]nͭ`k�>���?R����&Y�OYFN�y[�JmD�T	�d>N�ר�[��Nu_X��4��x[P���W)���+ֶ|/�O>�����`�:�-c��#����خ_��ڊzL�a�Ga��HKGi��&-�륭��aw��+���E������sh�4DtҖx����V]"l�0���ilxU��׵SsɃ�m��cl
������%E�6��]g��G��nU�ҽ���e�f��L��&����=���}�(!8˳�-;���S>� )�H{g��S�n��W�Q-�A갳�9>�Bj�|�_c��ʇSʭ���S/^��u��4�(�y@�-$��S�<���7��8d��2�s]�X�M)�5�w7l]ϳ��E��w�3���g28�L��4<��yd�Zc d2��n��B*Ո-�iu>����|?r�����G�/B�Z�O�P�WFJgT-��C
�i:ܫ��T�ɛ������*uy�SG���9?��`�@�0Pq����ی'$b�Ϗܽ��"����(O�n9 ���3˲8��Wv���t�G�iz�x��]r�5�l�8�=u���7�μ�!/oa��T�E(���Uu�ۖX��K]d��Qdv�nX��H��ҟrʜ��Qn���ti�A��
���3�U�l��f��[[+.���rAv�)?
�#�*Л�v"����E엣��A�Iq�糦=o��%�y�q��_h�Sw�s���p��|��e�ׂ�T��gT[��+HA2�z��R�Z9d�O�Ƃ��E�Rr�0�o�Ū*xñI�j&Q	8�87��l�7m��g2b��3QG�b�z9�و�/�P��\�A�L�!(M旦�S���J~CC�졌�n=��H@nl,��mR����e�c�K���{��pt�i�Ӛ���y��-B�р��j��أ%�����`AV^���2�t�37��ǵ�$/SY��k;��Ɇ�7�3dL����C/�-j;�=����m��q��zZ�%9�e�(�A�t����N��>wk��u1}�_�M�lhZ�+��qz����4μ"2�Ƹ���}rE8#[L;���0Y��� n<�X��ܹ�m�Fn;���pS���k�/���h@�j2��0�Pa��p��[�Z�FQ�`�mZ�2Y0��Tk�둃WTG`Zy�+�#l��Y[��I~�KYزY�4< M���{}-���-m���x�L�{�TSp=Q;�M��e�8��
��Y���ػ��<�u쉜ӓ��n?	���8^7�܄�F���E��ȶ��;DI�2�9&q��b��͊g���q����*>5�5�?sݦ�85ؤ�{.����&�F=���u��g�~�+W��W��/2a�v8���}�^Z�|�۳�xC�e�����F��\`<�'rի<�Pť��b0�"��`��ݙx}�\�>*>בyi�+(�˞���w���i���p�P�[��
��Q�
[)á����|9U>��v����X�y~�=��$E��p�7���v���fX]*2Rd�槶����1X#���-�n�B~U3�DsD�z��N�j�@�r�]����*�D�S�+�.�Y��d�ԠO|/V�*0M��i�0�����c� �g�̧�Ī�p8�m�eM�aQq���ٲ���}�����:�&#�c.��ڹ�a'ܫ��{��sˈ�B��޸v�;�t[ۚ��#B�-��=��Q
�d���S#��x%���	�6;S[�EQ�����fٛ�[��C�^�خ��5 �[`��J�� ��g9k��>�͉s��m�>�$SEqU�D[mD�]�3���w�B�Ʉ2�+b�^�!&�˭:l!�fn7�;������}n����t�Z�N��F�\��)��&��\!Y��W{M��*��i��=��9X��JӃ����o3Ns��ܽ!*��~�`7��T�{���.ż���we�Ggo8�n(BD^�onvf V�mctuV#ٖ.�'F<u�)eGPC�3;�WV�(u��tSY�.Q�f�o�0��`N���9��L[���&�B�\��o�����~��~�V�=��l*#�Ε�5�i�G`bp����@�7�z������Y���{R�V/�F��U��@���@.�dfq�n8�Y�a��f�<j^z�0};*� ���`s��]p��,M馒2�a�[��BG��=gf�k�������ɧS/w��[��F����`���Hl�������p��~'k�����»���e���R0{}Vf8�k9�F5��g�����t�y�y�S�\�ь���*�E���+FΆ�oL�E�t.q�s������/�]�����˙�ܥb�{o�vPW5��n��:��<.����I�Z.�Y��1U)����XY:-y��
効�b�*��z�(�0�e���\�.�S�h��p��O3#t�����e��v�*>�f
����
�{Ekە���O��F-n��$9/�T:q��䤍M�;�y�_��ycrW��&j�Ѹ��-pЧJ�B��e^�� �Af���}/lDD/:=�E�or{�9i˱���Xѽ�]�s�z����"�.����bM�z��gk�k��Z#�F��0��A��|g!����ɨ�qĿ�+�X9),avW�����FI�;|k��x9ҵx�'w*�d0)�Y�� v_U�`߾��r�����n�����]R;�R�=p�����)3����6���ѐ���N���d�b牳�	�p�Ȇj\��(���(�Q�w���ZC�6���k��F��M.q��f��0!�zd�Nu�d{:��_Q�S���+���*���1���/��вSD-4�=7US�"�9�iY��L�ח�+���B���f����5>��^�`@呷�.Ge��r{q�,�n<���`�\��V;�͖����!�k`,���M�B�+��çe����A��9wL���0�Ƿ޼��Ѣ��\���u@m�p58Z�Ũ��0�
B"讀mpn���]�H����;7�s��f%h��g��%���A7;w�8ﱝ0�Mէ�β�w]el2�`��;'�l�(���_����܃u|ª��6��N�5|;��2�J8"��ǪV6r]����uA�tH}s��/Z�ݹ��K��i_t�s�:[QU��sU�F,��n��|6���í9�;6�g������
��9��ҿ����y?RQ��H��%A�>����k̎<wl�q����-ך}�Y�m]Q��R2��o��c�r�Xxdi�d�ԋ�!tGP���'��?k�Dh��W>����-���%�I��r�i�v1=�ս������G�)�9�2F?��1�7�V�����H�؇��������[�b�����m'�:ڷ�-�w�o�	6M��Zri����ۅ���3/�K��X�7U]���%���5��0[���)�.e`.�bm;����vj�4̴<)��>"�xW��+e����A�}����5�&��ets}S�g���l�f�df�CWxj�J��"�����cs��˦8G���r�F 6�I�b���k�y-5Z\v�=m�l��kU3Wǅ5��Ew$Gpػ�z�{�,�"��N�\[��6�g9�x��OC_q���W�k��
��}�_����z�~�_�������_�<sgY���^YF�rʱ@S�2�U�Ǜm��ʒalf�h� �ΡS���Q�Rv�����5iZ$[�[�����y�-'�o9��5sj��mq
�vpR41�MP7���5�H�h�Ω�>�r,��t���+��.]�RO{.ή��@fޞJ�锄v�C�fw�|�mⵍ�v�-�wl������.:�h�j��λKZ�v��qVlR<w�ݫ��u��+U�v���+/@g#�y�֤4��[9��PsJ ɻk����i�vj��;�Jq:d~�.�/��3�����4U<Y�ք�c�:AoH�=4{Zkn�r���)*_u��y��H@Nܗ1�o�5'#�4͇�
��]2ƢN�Ai#fq�`�xj��>ŏ�)�=�s)Ty%�@Ӑ�`b�dJ�XM�ݡ(�keq+7��)[�
$����I����+6�`�Lf���n�h��r�$�H�.��̲0B�v��]�[|�����]�ݣ��&ai�S;���-�X���E��י#o���k�����b�n��U�tBnVa��P�Jq=��)GϪt���SqZ|��/i]�8��m����I��-���*μ�^��iEYRc�!��D;k�)}��nqp�KPǔVՙL���o2�$�g<�-`�.�[����t^��/��i=��_j�|�꙰�/iG�s:	�ާ����r��i}�;���n��u.�m�6K���Z�A52~c�����6ۨ5<�]׃�Z���z�3p8���e)_��7���(xV�t�kC�S�^)v��^ �$��)�)P<��X;id&��>�sw4Х+.-Yʻ|���*�Ǜ:�����ӗL"�&��w[O�>��Uޙ��<�b)|�V�hr���q�#L3�r�-��f�آ�4�fw���}Bf6�b�hGv�`b��:Bs�:lP�hв-]5�V�qFz[�]T�pB8��ڣZHOq�Y�`7˔1q�zS��% $U4�e8l�r1���ɵ%��T��	@Z3p
�v&*�@��_Vig�7J� i�k������5 *f.�Pҕ�C���KG^d*�J�b�淋�hя뵫�|���۰�n*}@��n�5�,�Ҩ႖u{P�ސ	窺�>^�<ol����G���|rs �x�gN�I��/�f�i{��%WU�y�ՄC��u���W5�i�ad*kw�p�,��eokK�4Un�m�������[z�n=\���	��T��B�<��Kr���LJu���AT���ͭޭ�r�}-��
��ZM��<�8裯VS�&v��m�_		r�5���5� 3��Zr)xʖ/"�&�\/!nKº�FΡz2!�w�x��ۥ�>3����jU�L��;��q�E,cw(,|�.�C�RH��}X�m��hg/�ov�@��l�b��9�T�v��hZ$p2s���r�{��'!Y��$\ZN�%|���MY..��s�^Ȝq����ZL$�� LL�Ɛ�}�&c��0���QJP�J"W9��W3J��/�y�$��B��4���L)ew]�O��������
9�Q�.��RY2H�,TNk�9��$:.u% Ҝ�n��E4�u�ba4��9�~藝]��e���.�6 �$�w;pd%st��u������;��߫�RC,O:�Ј����E0d�Cw9u�y�I1!�I���J,��9#���,D����n\�bP�F��67N��(��]�I1$��i����ݐ%˱3�F�D�I�!!E%�R#cHY�IoD3F(�Ĉ���ȑ�L�H�u�,�!ڳM��7_��Dօkz�Mǭ��h��r��z�q�!�BX���vX͔��/�Q��a���;L��	��7 W���^�O�pg��|�xGe@��i������kh�M��kҺ��>��j�z����Vq����xK�S�Ii�ϥf�m����~�ӆ��vZ�;O<z����:����k"9G�D��[U�U���>�x�o�^���|��eϸ�4�%JH�
z
̈TփG-�)�"{x��k�vy���M.�N�;��v������q�FF�M�g] �v���z,�FC�L��Y�k��̜���b|Rd!��
�|��{��*�$Y�]�,\|s\驎�?����W6kڢ8+�;h��31��^���bz���qs�V�=� f�]�?*�����h���78J�p�����D^����,�-�����U�j�!���D�G�������p|x}�xwfy�����5U��\aq���[Y&��W��K��'d0�SM�O_")��c%�a��VXa"y�>�/�3 ���M��7s��r�58:T���U���mӈBe���Ca
�^y�|��d�I�BӁ��0f��㱰IK�����trո��݋fJ���b�k�]����[���X�'Φ�5�t����}\�������?�Km��=�j]~pyS%GU��?�5�w0��r�1�{��^1��]K�|/�	��,�.���(�<.4�OWu�����|v�$�1|���m����>�ʸ��L�S! k���嵄g�$�D0�x�,[w}s�۔:�x�'o�'�+�gA�%�?g�[ѿ��=��n���ɩy]6[(�M\^�D�QZx��R9����|�x�_���p�RxaT��y�q/4z�� n5/L�óm����{�)�yNϸ�9����:�;庮�  u��f](��r��a���硆��~�YmǷ���1��i�4��*t��W��oK�3lrnx{A`��)��+6�q����:�����Y�n��J;���L�}�}��\xK-���6$CB�-
���ѱi�c%�fT�w���2K���Y���G��r -kXFC3�R��|��Xj�2{��:,\�#.����n��P:ik������iM�����ޫ�q�W�wr�����{�Q��ڟ��6�|��|H���?��\�)���Cu%��H�d�Se����y�Hbޮ�Ox��w�Q=ͧ�r�}z6Fm:|+k�ڳt�g>@�2���}�E��izGٗ��T4gl�l�h_n�2��}���n��,�Qa��]��k`kaM�+/bs��P�Y���ļ����7�ܠύ�1>E6O�����	m8�z:���j2�^��5)�ӽu�f�a��7s�d�)��LQ�+)���)f�gcݎ�3��F�qp&�*ߥ��{����ʹa����6���	m1�$�ʊ�=�m���n���x.��[4�4nǗ�`ˆ�78&/�ag#LD#�Evd�������H���5��l�7�,wk)��=��s��*���<�L[�X�Fk;^zduF�!.�f"Vm��4�����c���0�@[ީ-Ӳ���7�yun?���}Cb;��RsO!v�~ܖH�Q��lk-"q�۲i�[/|��W<$z�v�-d���({���z_��ofmHY�:��&Ԕ����E>¼���Ռ_9O�R��L�w����5�u�#���6O�Ǻ��i�t��f�d�f�o����r�nՉ�U�5f�n�V������[tE&�/)����S{���2;+�9��T��w;M+G���od4]R��u�/����ںÔ#ow�a�p4q���f����靓{
;/C���x�x���]8lFq��!�������"��(��a��;�77J�8�5&�R�q�qJ^���ē֗�C����'�v�m�����}���ڦU`pf2�2�sЩ�3M�ɏe�8m���d��*<{� �뜀v�n
Vdp8��vtmD�m��Y\2L�lӁ�lk�Ct�w�=`ߓ���&����𬙺.�T��	�uH����0����n���<� �|#uNAmUɞ�ϣ{��mUz�u��:y���;8���G.˂���SM}����������{M��p�HW�KUq���;X���˥���m���v�]�8p��ȟ�͟��w��Z��U�5�å��S�ٰ�����F�ތ��wk�N�bd�v��je��R�x���id�AO�e�4�Pq�yCf�f�WQ��t���n)q�[Y>jUrܮ�j,���M^�ޠkyd�����V$�Wn�]7���k7��]��IS���2�S��,�S	�@)Z�[d��>m��̃v�աp��X�+��	Gm�[�7_<���Z��T�0~�\�cwm�y�̱���-ݖLЩ ҧV�KZ�<YU���hP�,�x�6tw�����P�(A�|�5f�yf�~4DB!�Of�q[H���ۃ�G=g�z�<GJC�{�������#ŻSa�.��n���+b�ʴ$�W]?��z�����,���\���|1��גN��>�ɉnh�,#w����ɶ�Z�eEDeVe�	�Miy�/K'���?�^8ed�d��i�؁�ܞM�UoB�v.��������+-#�0oE]*�����7N�u�k2���k�6�Z^:����&��f廕��q��e��%i=h5�",#v�Q�!�斋�����0���¹]?�:?e���7��u��~��}Y���}�-m[_e�����o�Y����H�	z�L��M��_���4����0sS�&�7ұ�ks#	m,�}����9�*ƶ1�{���Fm�㾾0}olm�R#r|ۨE���뻑7�L����,b����2|\�u(��&�7�e�訥�����x!�!=����:�,t1�4���l��Ӽ���+�w7Y��쩎Jo�B�͡Syi��{j����2^�ؔRw(����̥ifTѮV�,���si���;�g�5�bX���z��'Bg�-�8�-Y���8�5�������f<LQ+�Xڨքcz��9�A��m�GW&�[�5�=��d]�?*�rlo���:˧�h����źkx���o&S�Wt�qmyTذ
e��T�B��,������b�^�tWb݈�])u�+��&�ժ*�<ʮ4ѓ9�{u1/K k��@�s���g���p�d{o+fJ���[Sab���l:{_mG=�fD6�d_��=�d��;�MY7���O����n��vNF�י�Br�%l�]Y�V��&6�˭�`���@����&�w��ZS]���/��&�u3�(v\�Y�����@ޖh���w�X|�:gE�|���Ku����֖+��,V��>����|+�9mS���k��N���,�.�e\�@��vJ��}��q�N�qzx���g���Vv��eV�����\v���8Nu=#��A�s��V�Ұ�,���{>��`�与���e�y���;���M���� �J30n��a�^��o*�����,v⼉�O���Ƶ�;S�&�yt钺*�̽}���s��\�d�5�@���J�啧OyU ?/�z,k���8�_iĽ�>du��7�ኯ�_�fI�{�3����av%
'���C�c�e�7f��7qަ(�C�B1c}o�D��N�d�V�/6X.��+)Ԃ�t�n޺���0-S��94�	�w�e{u�4�u�r�`�L��b$.�F5�
��@�ћ�2�6���r��{=�y4�$[%���s�t��)�6]�����-�a=�޶��΂�ʨ��Zg��(��E��7��6�솖�W�n���b�v��8է8��L�d��r�a���͸���+)��ª*;6�ĵ��Ÿ�; �3t�'�#�\(y��]e�s�t+Ӌ�L3#��gVT�ӄ��]gj_�䦉>�[�^��.x���� h��;�+*�ћ�5��wS;�|x�Qʹ�[\�"N�K>G�|�Pz���̼���uq]��팤��ʰNT�5�ȄC
���x׼��6PU�}v�u�#|'kz�����އ����C�U�&'��d�TUWoiLm-��L۽%�6eҨ��1
7�[���:����xsr�j�u�}�6�c���Yވ��8�uSލ�����t��-8ė��[gw� E���h�zv�l��[},� %�����<����� ܵ$rT٧��*Z��I/(�|���.��'*&��4B�Jr�U�z���oO�6���_'�i��o|����"{6��Q�J��Y�"=KB� �����܊�Z皖���'�ȸ����yH:��{�z��po�� 6Z5�������nN�Yrr.-��q�FSۺ������k��)����!H�Ƹ����3���FE�$�U�cU��꛷ڧF̆�����r��܆D42D�2�٬����S��ߵ�GI�h�F�����9j~��D�3�j�%�>��ӳX�V:9�N;]lbn��bW���{ ce^b��O��&RȽ42T��R��g�����ZG]Q�2�]	���r^�[D�]]�|�#,���e�)��{��9�j��~�f
�<TV�06�3B�e9�
;�vcI�ݳe���>��,z'�q5�`�=��A�s�w�m��Zļ���d'��fG.�̆���h�9���)����ݚwA>�EO�S�[�{�o\����������~T����7t�>l��{���)�`�tK4���$�xae:;�5�yW����r2�f,�ڬ6C�N���t��Vz㖋F��A̴���Hdi��,��-���wv��[L�1)���a^:��6�aS�r�iŲ�M�J��#/�ϛw:[6g����W�E���jU|�TӘǽY���w<�i�ǵk�l\3eNkY�^l!y�3����m����.�i]y^c'2F�S>:���{c8��ǫ��z͵Wyn��SƗ"�oqn
��l���Yp�v)�f3��y�c�8�Z�.�}y�X
�O5Ǆ��b������:�T��5i͉�|V�K;��]i&D�u�y�����w���mcus+}���=+�/s�lӍ�U�;��f������x��(�/g8����5�'��p��UqKv�/SI�^Ld�r�i��δ�1y���������*��#H�u�)�4�S�A����8L���~�� 2����y�{v��!m��*�~-��-A�rl���<�J�-
λ2r;�^�Z�8�p�����9[����vMnP��ɵ�:m$Cc�d�j�rK�w;��2�܀>T���l��W��f��rcL������z#��h���y� �6�a�_H�⪮b��x�Ru�a`i��T&}���x���p�<����mF���ݾ`S#U�	�E��R�g��J$��Q�ynM��]�z��߳���������t����QPW_�x���#�����G���"3��C��_G�+f��L�px���d&�r�����G��l\^��}2���� ��P��\y��y�Z@�ݮ���B$Qm��i��f���,�ޫ��@F�іq���V�)�=S;�׶��;0�_�M��r���-����)œ�lmaJ�km�[J�l��ͯZ�XW���s�tx��5_��+lG�(���P���n�r�b�T��,���""�c�������/RЊ��s_��ix�~D�\����x��rQM4h�P��9#kzsv�W3��=3e�Z���Ồ3�?�����{}~�g����{=~^�/?�..z����b�}���VQ��m����*΢#t ���h;�I���)u�����o�6���l�B���n��y�fc�S�M�"�Cc|�S�Zn�Z���5���ʏ6�����΁菩�]�S&ǈ^&R�t:j�^vF��U���[�����2b�7뛆Z�& 7qn��H�N4h_�B�4�-���om�We�[h��O�+�N2ֻ�ǈ+U�쾾��3��q�9%w+gan.�*�w�7�7ǔt�c�[ņ�ay�L��[��u��t�G�cUM=����n^ۺHn<��9�Y�	���7��KT�6�����T*n2�b�pH�+.�ø�8���)F��˚�/S�ƙ��<;x$�(�
��l�K�k��,�=X��/��R����a�c�"!g�I
Y���5��d_T��R�qm�k�+��4;��{w�C���SN�9�ƭI\T��.+����76���q�n���"���j��� �%9����]���Cv�!�3)Q�(0�A-����ϝwT�GA�Si��-KJ ;�"�֬ :M�h�f�����H^�]}z�KɁoQ�F�vK�T-o��]���,)�͜�L���p�8s�W���+�1�9լ�U*b������=u�в��ݤf:}�S���V���JB.��ھ�V��/*ᎴZ�<���מ	�sP�'�Jg��X�wi��
10��d6�ZoZ��f�Q˭�L�,�k|!9v�Ŕ��"�)l��Gh@��$�*M-��u.�ŷW(Yaj�5���qM
�.9�<��N��(U�h�fe����/�|�v�ޒ�7�jgb�C�Z|6�/��5�&�#�5�3��=��QP%���j�Y��{.WSxه.r�W�лڂ=N�DZ��9�B���H:��~�}\���|ݔ�9�t�l�0=��R��6�[E��&�Gfm��c���1�SCxJ�Y��@�ün���>Ou�oo��_,�t�������|ާ�il��q�)!�n�Sò$�Y�K�Ym���[o��Č��p�������{{Mj��K*I�3��U�/�=�lϮ��Jk�н�y��ǴV�@^��з��r�Qa���RT�6�sG�{�|k3��s�8��6�����rE+|�uj�3Yt�j'+��E�[\YCA�;���ǖf��TϦ� 2�X��6�ɑ�.et�4�o1�T��Io.�������p657��A�2�c9�dQfSN�.Z��^��[Uvr�o��vHZ��.���Z�"��Z�F�V+�sU�yioSŔ�t-�����C[��V��B�W���.O���iˌi��wEgK�s,�ۮ�a[,��΃��kK^�KG�"J-��z��5'Gڭ�`;`˼��c�bЎ#�����}��̻�]��/B����Ǩ�[���gvgn����FQ2����>wξ~�{��	"�Ns!0F��\�:0D����F�2b�"�)"a�D���F���s��E�t�\�9v�>˘��x�~�D�2F��̑�n]2Cb���$awn�fIcH
@Q{�L�}�f(�$Hh��A����T��EwFdS��Rx������\)	200��2bH<\%����Ł,k���"!_g��2dA�3>y�
^urf����.v��wZ��BL$"�II�)/f��w#x��f%2RM�IHLf6;�8��i���2fe��LȄ!�ů;Ƽ�21�]i4�C�VL�&62�3D�&�IF �.��M�tc@�O��$����!e"^"�p��~�h�~�:����4�.��B���}�X;fG����ӓ3��G������'�`��_@�6lx(���,,-R�I"C P�x�s�6%4jl�x�_��ҕ��B �N���@Z9�hJ��&���8��q݌h��K�x�y.R�a5��^�n+l�m�3x�S%�!߼�~��Z�|����S�qT�)����+x{����5�L�NL��I3Es>�^Ub3x�Wp�f�#;�Dm���3^�4��+Iٌ��jE���`��<y�)��7*��g�Y��=[g�+��yV���okGE��)3r�d�a���6��,3��2ط�q�n-p�*�����Uh-���9n}�y,ç���R����Y���ZmM��x����e���>�78�kDm� �e��2r�$HR���5�	0`s�<�>���u�kk|X���ڝ���c,yեA�H�+�&�X��Gm9:\�Z��W�'�4v�h��W�i�GKCu�QL��x��!]n�@풳�ꁘ������a�W2� S��s6*�A����W��?�bn*]�01,�+38e��ړ�KF����6],;��Ͱ�6^Yw���]��eh��k�=� T�2i����,N�k6��Ҍ�w�x�d��<�ϒ���1�� ��J���#a�}�#|������SRͩc��s6UGX�V8e�lz�5*����^+�]�lf�神��3�<���v������&CQ�90�du�guT�n�m�Y^�yD*��|�L�ס&��a8���Q�jzf�oT�����l�槫۽���������>���堲ݧ�<MN�M��(�l�G���*�	�E^�����]���	���ǪS"!d��&ރ*�3�)�1�E�+xϷ�<������#��k'v6��Dw�otL�s���xρ�Z���ni&,m��*�$s5F��]ǟ���e����ռ�2�K\�<��4��{]�߳��ڥ���#-9톾�\R8qs��.�<�[�m����~f;�-O���o��y�������;�vc ]�v8�B�3w�j�먝+)�s���cv1���o!HZ8Z�/.��g���*.̲�ї���w<j���hɗ܇GnghZ4m���6\��w)�ʚyV��ȗo~�k�A��>�c��;�Qs�Dr�\Z��7�j���	5Ol�GGW�p�6��L��X��^ktEvZ��a�+gX����4 &j������pӺ���ݲo��}Q�1�ہ˭9/����іb%��Ý�k$6�f�gN䧀�M�`�	�ya��SVCe���χ�k�2g��H>�(�}��\��6��@u�$DYR�7�L��5dn�}>E&��d����ν��t�y;{r"���g�6�*Z&���W��
����/:�B�b�E"�gR��,@c�Iu���@t=��9UH�S��i��Y�y"d���RقpC��Ȧ�f�8������u$����;c���r����::�7U���Ʈw/�F�JT�3%*���aO�t�=�{i`�1m�d]����
88]T�7&�:x����\�����spܫbZ��͟.I��UY-�ܣ�6�l/��N��
������ĩ�
�[��F�"v^�8g�1���2�^�`��a�3@]�PYu��.����E^�����W^�|~F��;t�)�p�"&�I���~�3&d9����*[�gM�l�k[�oof���@LɘܻLv����,��k'X�6�dܦ�&Ғ|8ݜ]�(͕x�ˣ��;ӹ��]A�|�s	�z�☮�q���g�������n�I"h�E�v��4t�w�r��@��oW�dͪ����fB�XldV����ѹ=I2Ⓐe��6N���ǯ̬���l��Ԫ�L����d1�ޭ���8QtH�D՟���x�V���m�T��z˛�f��o
����u�L��Ft[�8K��G\�;L�
��m��Q\�-I���*¦^�V��y͌�Y	�z61���΃9��;-��8�q�"�r��u���}d5w����澙��+���Kd2�)���l7�f=ϻ8�{�x��{ٺi99�0�ƃ����YxO�|�aYN�-"�l[\��c�,�x����q������e޵L˨�����0����V8)�sqFg:�fUV�{�su��H���ċڷF/au��*h��j��ѕA�p����/+9���T֙a+��r���3�J�R�f~����F��X�	��[:���]��t����uR��,����,�N��=N��a.������� �8zD���f�TS�:�+&���'ݙ��ϧ]	���#Q���q�}�̖M�.�[�[Y�"�
:�{iG�3���Y�r�d:k�KJto2`��z��pj�����
��}un���fS^
�������R�гy2�+���y�d�Z��U9O�ގFߚ�t�^5a��z��J�U�g��q���2��M�U�����|O{��^��KK����F`�M���޹,ƾ`l�J��u{�S�s$Z�F��e�����רØ=�[>���i�.�x������xJC�:I7GH�mWq�H^D��w��l��udy�V��E��3�G[���:�Uk:pf�����6��:�^��ʙ��O�s�gS1na���H[�<�ON�5u��&��BQ�4�V�N�\P4WgT��t�2�ƭ92��8��n��̼c|�y��zg`nuV�YV��}����H!m�;�ū T@�g��x,�:/�f��y+<4�wj�~={)K��C��Z�tc�Y��m���᎕'i��m�Xu�&]�ڐiþ�0�|�����ՙ9��i��q���=�wgj�[���W��7\;�ф;�o�͜kм�^�}K%u됥i�i�[K�}^�0%�Hgs]O�'���N��=�Ӆ9@�&���Ei9��)`�N2�P:#FY�st����^+�XN'jm��y
��o�O���H��W��ar�����	`m���x������'* 3Fd��Y�kl�k���;e�_��/L���"B���5	��Sc]�\n��a��I�y��FQ���&7I}fH�uX���!_6. t��m{s��:�!�]�b���*���ht7nSE5�y(�e�ՉËt�n26f�AV�cT s����S��R=�+�n&*�Ԭ�p�)=1�z��=so�@LO՝�L��=�I;a/�9�=xs��9sCr�*�v^�m�K	ϻD���YL��Sb=V�e�m4�,�ţ#ƌPX+d�ǚUУMX[_���U�$
=HB9lQޣ�ten�,�;oF����ʩ�L�Q����wfێ%���im���.W�06m�YWFTu���.�]:���pu����^ɸ������ܦ��o;�o)m�\K��<c�%�����������}lg�{^{���mC7@U��d٣Z�S�i]�#P�M
l����c3`}�s"��^��3}d�AW.�z}�^��ʴj:�4�����q�ip����q�FE��l8�9��|ZPm���N3Y47];f؍���TCN͔�>ةN�I���U�'7���������~��Y�6�*���b��Q��ƳZ�����+&�\+���O�1���Y��0g�}�{ �S���M�r+�B�z#F^Â��W�gn��3gV�7Y�(���v;ev�+�
�����)��8kDq��yY];E����i�9��aeg�Xy
@��ȱP����r�\o7T��h�<�Nv��k4Խ�i�h4d�`g�<����J&7scF�˶��cmȎ�P�b��2ɞ�� �����Ѩ�Tu	��Z{�@���~�4u�,G50���9}��Uߜ��n��j/-Fc��,��\�㑆��h�(n�Hs6ط(	���3f�Ȗ�=�5q�XtϛQ[��/��՚��,J���ad9U"�ϣ�&'f6�jI��r�"Ѯ�q�׳�|pÙ�Q�q���j��`��("���ޟ�U��5����ui�[+P���,���xݡ�����z-%�v}�z��qNH]8�N��w�GmL��r�� Ep��[��[�ǵ{2��(e�\��զ��]�*s�7�຋]1�t�F��r�S�N�����Ѣ{?7N�܍=$T��m���ٿ$V��fY�,�]SY����K=�sýv�Vm�Wf:�:3��v�<�<�Z��p��лm��\mmd�*��w{W*7��j/_����#g��j ݶ�������!nSٶ�Į�������"깆�W����m�kv�T0]�����v
�K���#{��MM^d6��^��1u��n<I�
�s�;���[Րb�=g٭��][���&(X�RfX�E�3�8���
�͎[%��c�N�"����W��qZ9�_%|Ա�}�vղF<����s�c�>d��q*�143WD��D�:�:<35o+Y�Q{����g'�X4�}�?�śQ5}Â�oK�3�1S�f�Fk��:v��~��26�������x�qm��L'��tZ���u��H�2o��enI�þ�}>f�����<~w�����}�����r���}k);b/jI3��yz"�:v��5Yjk�z�
c/*oR��tqI6�fVJ��vr�r� �]	n��3/zY��k��vN��\��	J�t#�;�3��$CR���OF:��ǒ����-�:�t��:�I�>?�����O��^g>�c�d`���~�g$��,�kk����ZY�0ѫ{�Ҙ��miΣ��|�g�K�G����uclT�3o&��x�\�ӆ >NE�,���;=1>�\��M��^�m�i��nk^Y�sD�ᨣr,Ș˾�����-�^�4׭c2Q�֙M�YTt᷏Y�!����jTF9��,c&����ޗQ�����m�Y^�L���o�Ŵ�^ST*b���gm�/t� k�窇Ur{���m��6at�R�6��Fk���Xʪ8:\��j�x����S>w�/R�H[Y�=U˙.��~�}�ò`�ڣG�ݺ�M�i{�� �_�Tł�������x�1`��k�ط@zmr�V�ݙ;:��iS�>�s���\�[����*�r�私Uz�����.Z��ίJ����YQ�rJίo�(^��?^q���$�[I����az<ʔ����:����>��xW����&2�iD���-f��d�]%`u1�2�Um,���w�퐄D�6�|%���c~��9��CnKӻ�2Sq�A�oy�`�r��帕].�B�`{\ѵe��u�{ft͒��9�z|�ɍ�j�2���3q@��j|5�Ic*��f��1����&.A��\w8,	�Ӧ'T&̀�[�,�!]�@7���u�$��|�xI�<�5�f�Φ��^������֟[�X�fZ�@�;L�ֱL��C\�,����~�������co�03��[.ሆW���ibx�������6K	ޛ��՜��]��^�2γ��@1��$>�aE=V��ͽ̋{���0��1b�2ݖ<����;�钔H���W
�$�;�[�[��̐\��f7�0"�*Ѽȋm�N�k�ήY+ʇ�p?{�7���d��[����z��mh���},WOWae�b��_R-��Ю����M�K�u�MNgL@=�c&�t�D�$��q1Efd=�|~�9�#r�Em�cQrIʦ�����m�~h�=�nV�3W������y{=��g����y{�XAT�`�@��/+��B����F��꿣�p�f����٤�WS9S-��u�0�ږq��<�Z�+R��L���2�4<g6��r�n֋�	"���
���.Q�:�>��2��v�i�P�������d���R�r%n]�xh����Khn3�$��O�5�Lr��D�7P쭢����n�O81w(v�	��(�w\�g7m%�ӣ�5�
qI����!�Z��j���A���;��eMf�U�E�Y�i��V��m�����*�D�F�%����A��m��4�K:�<�>2nλ}u�w�C��� �����ʵ5(�nB� ��(h�)�0L���y���,}�0^8�]�xX���j	[����m\���s�K��e�U��ͧ9^��t�yV깺N�:��>�v�M(]�]�3�iZ��^�h{�t
�#(>�w���E��=/W9��H�ɺ]�7,E�"�E�U�
Ɋ���WVt�R����s�L2���S9s�naN�6��;M)����<��w7Vh���H�eh���b�J�[��!�kU+mB���ȯRLɳ���is�:=���ګa���g�y�QIv��wUk�8�P�u@�S�m.��N�T.WGj���o��@�(\J
:!��p�]�Ĵ�_ ���cY�/#��,纮bzt�i�� oC]���
�	q����Q���;�x�e��v�����^N�E��sM?�y��F��*�m�mp˰ޓyJ�-ŵ��Rl��HN(�j�x�Aw/��s����R�Y����,bn��2�g�/	�����k-�V!淲�(��޻��I�X�$�P��RW��jH(Jc"�f\U�*n���r�p|��1c�S�o"l��WW�e���5bhRv�m�9y�*��&!J�z%M>�,]�2��;���.���q�B�̃���>��x^���# ޑ�9�*T�194's�� W̦��d]Z4����=�]<�����XU��%,�dV��&
*9�k�0l�����%>]�n[�Dڷ�GL��8j�_p�@ͺ�*WY�O]g���8�6�I�t�OB�3���n�y7p������kz�<;ɞ�e���#yh��\#f�͚���ম�i��l\���˩�J2������6m�
�Nd�ha�)�S���gVnV]���t�qu�y7'؅]�u���\ͣ4kҴ�
Z5���w;��p��vg͜��ޣR0�/�V�v��f��Q왐wSS��vJ��҇a@kJh��-��)"����Dй�W;��8�{�%�/k	N��m�*T���
|����9	˫x��jǋ�(`�����ڔVY�⧂�~��#k^G��̷y�E|�Pu��h����Ôr�t��8��悫a�-�s��S�ӣNI5�F�|0`�.�A�c(�"`}ܗ.�L�\��lb�v+��d���n�!��� ��Jk&���Ɉ"&��>���fS#��u5�\� x�hΉ%&hL�I@��2#yݘ-s���6#2;��hQ;�`��F�RG�u�r����xBd��Ff�lF�Wsrd�WH.n"BA(̱��u2�y��؃]���\��ݻú�v�����J1�2�M,BI�.ԟ���$!.BF�Ӷ��X��b��2E9q D�]ٹ�"��Ź���"M��1��w1�2�	ݮ�L��F�� f1��DDdJ,�1����Rs������;�����߽۬���jk���&q}w���-}R��Nc(�*���&-��^'E���V�*Č4p�:z|ܴ�����K��5Y Ak���̊;Zv����Vj���$��P�#d�n"�T���B��ʭګwd��l>m�xNͤ�"e����U�[M�Iݙq��sY��E�����v]p�J+���aa]���o�O�Y,�J��h�Q�X�-P�����Yʮs�l<9�c^J����V�*�\K����t�8C��L��ݝ�=��5�Y�k�?NK:^�M������6�*k�Gz�#Mr�/k�q��]S}d�� ʲ50�0i�Q(�p��K{m�FU�훴K��˨ֽN��]uZ�1��4wo�v�j}�o`�������D05��T��s��=ԅs�d�w�|y]5��,��}=�g���>D�?=_��׺ͪp�js��l�`!��Z=�I�'o�_{	O,N(M���
��+'#�ˀjD6��5�c��e���92����/�W�+���ڰ���ȫ]�{�[��t��t�`���qE�W��g�7k����^p��s�S6Zښ�y�K�V���ʯ��>g���XRƪh}r��w���[�r6;+3�;�O��A>���XU��7k:��sqg��#"��&����f'r�8���C�~ЏA�}M5�g��j�N�O��(�ͅ*�=��/3��V��_@=m�L}� Χ��i�ǅ�-]u��l0�Jn���l�^���'�h�"	&��DN`��4;%��XΝ�zNö>�tj���ݟt�M.j3�+.wg=�G�9T�6l�G��y&�x�1�ˇ��<@G::�lJ��x-�b�z|�pn�RId%�Y��jS9�s��O�Sȵ!�_3ގd���ϙ|էMtA�ࣰqG�ٹSJ���xS4�I�r݌lhwm�=�U�V笰�����.O(�=T��7�DF+��/ۣ��r=�j�:�N#�t�D��o$�]�g�5sY��T_]/'+͜{i��3+�������%���3d.4jWV
�\"�76k���VK��:㨮�wS-���]����	��g�⚇<�<��i�`���!��Ę�ی�}e�	�M-��"A]��ln6Y,�R_��T]�|>����b�n�qZ��.m;w�n��Ǯ�4�f:7NS�����Iә���"5�eJ
��e�x�����Q㎺7��'m�>��\Sy���w1��J#��t��ӌ��a�&4�t����j��z�uSrHK5,~�q�Yi�ק��͆�SL�9 ا��1�K�N�J�D.�͍�U��tq�84�ק��Ciz��#2��#��ۄ`���ŵDm��}W�ױ��y��1L�xjA�clS�Ղq�I�,:u>�m�%���eF��8�}n1enN�\��˶I7����]O�Y{Mg2�=���DCB�/z�K�1u��z�CWf�.�oݗ���f��G��~�V�>�8�z�B+���m��b�����-'c�p#׉�.�3σmb/����$+�|2#7kɰ���ݲn�����3��mP���e��(�Q�b�sU>5�(N>�~aϸ3N^w[Ȍ�-2���l�=tȫ�o{ev�Jj�pMx�:�9�˝SFc�u�D�6��C��E0�v�!�z$��܄?V��l��ۇ��h3,�i*�����t���؊KS�:���w�{��,mXPd:-���7�����k×{�Ke��Au_l�ľ��d����+{��F�x+h��[Yr�b�����������©�0c�������_���Y�羷����)���WFz��O��z��9��9��V_`�{�����qؗ[�Ul�*�꨿q���=0�X�A 4�q[
A8��t]�]E�7I4��q�"M��8�}P�2�լ�wZ�*��{�j�Q����U��5W��e�>�.ʞ���ִ��Ƙ�<�y�˽*f���䷠,��S�e�W	�(�]�\���N��sOי�� �������@<g��zg^�z���8�f��p&��rl�w�z7$��_���o�xS�g[�ϼ���r�>��U4��ʀT��hQ[��X�W�y��q�'ځ�O��pl,��ZKd�$�WcԶOIt6�4�N�l��Ĝ`dϸK>�|�����癦�ZBLS�����ձ���?W�_:z���O�Oei{n�TY���ӥ�����k��|�a�Wfm���Q巸�kjf�;rӒ��.�>ޣ���~��[W�s�w��gF���Kڛ;6agk�b:���ܵ��ϲ����nr�-�r�dhOd'u4��ۇp�P�
Z��T��ޱ�"[e�"n1�T7 jyc]��f�"�j�OK^d���%�g]QT�bZ��{�������s�s O�(~wށ˯]v-�]xsζ����Z1�Y���gk�ڞ�g���d�UA�ߝ��5>~�A���8 �u�V�[�kL���jw)�Y[j�\��N�]ߙ�G���r1��\ļd�.{[���j�~���X�8�ҫ�U����p�w��ٻ����Cc����˜��U(��[w��*�-�Y�,whS�.z˾3�ɣU����Y�S	�ϯ�V�Fi]M�"��Iʹ�=���fD���ʃ"�D�t�̈�����6lQ&{F_�]Q�K
�R�Ҹ�감�جl0=P}��S���<{�X'֗��~����Cg���<'UH��F��{|'.��^���:�è��D�!�~sx�{]�S+߹��^�en��+yJ,�vHb��;��v�[�ӝ��'C�@f�Kv�1�%����x���O���~�fܐa�*����\P�y��i� �G�S�U��(�9N
��ȕ��}J���1)����7]�omR���{���&���s��&�o�/ۋ��j[�L�ӕ����^2��o��|�Q�i���z[�f_Kʝ��S�	�9�8��\�,�v�=\ptߴ�>`�$em����Tm�>�M5� ��r#�\Vv?����{P_ח��$��1ICZ&����bd���[b�Y���SWEf#^�-��w�[�7,QxB"�֨ݒ�����]x��{"!Y��単�vbwx�^L�#:��<�-��܁-Y�,s��zA���f����鶺�֓h�Y�zoD��&�i����&�Xxdi��e�[�R,�EG�0�G[��>����,eE�9^�L�i�53�z"��lslk�<WK�A�#�2���~�H)z8r�FnJ�)q��J��1)��6-�Z�$9���D�;�ayg�ݨf�>�l���v�-�t��7�v�Kx���g��܃\R���+�2�l��7V����n��ã�gI2��6������
.\��SRag����J�1��`��ؽ�.%9���ݞ��^S�̝�=����=�x�͍��"�W�qЗ��rFw�;YΕ�Eo�2�}�6�hQ��36�W.��_= ��!0��+�<�w�G�X(�>j����%���5�6|�Kf�U��Hψ���(��`r_l=X��ݽq��N]�TM׶�Ndp�`*%�ǭ]qwڽ�Rs�X㚝7{�ч��e"o�I���<��m��XOT�����(��d�9W�-�)a�G�A��� *]�����f��1uʽ$�{��͸��YR��e�+�z�WE��b��J��Ӻ�Py|6Y�^K�hV��M��ָ�5���;b�h�وP�s;�R���5&��8�Q�~���M��ڈ��Jf^��lio�v8���\�qw�3jH���H�Wcѻ�b�@����&h7���
�^o�׶(v��C�hH�a7�XL��5E����c�X:3Щ�nh�������.e�]קּdy�a��+�Uˉ֘���[/��ֶHYܛ��d�=4y�����t)�eP������>��ݶ����|������7^1Ba|`��o�Y���[��ur�b�&D߬n�Ѽ���_����:����P���;:�qɇ�A׫�9�Q-f��4�.s�W*��*r�ɨpV��;;�\eʋ�r�q��YH��<ǩ+��ϻIk���;4v�׬��������x��>E�=���M>m�·CU�jx;��Y9W-����0���_�)f]�G3��ˁ�/P��M�.¦����e�n/]��J��w���B��	~��XMk{q�`^p�-�d��>K��N+��dd�Ij�TYGOg]s"ޒam��#K�WR��6�q�3��L��d6�+�ڌΫ����#'h����Z�b�"oT���:Lϣ��N8k������ŝ��s:��A�l�-�f)_S]d7ulo��r��2�xNaV���!t���y7�j�݉O���qG�q�;qc2�b��Aॸ>�փ�E����d���W����l�:q?g�y�]�.d3OXˎ*�	��g����qF����|桟4��Z!oF�g��Uy��QH+���ޥvjڞ�ު�4��M��,w8�_����`O�j�SI\���So%��䭜U�˲�鯜���t� �ȁǵ��ꦡx�NƼ��4�Բnt�j�Ak��wӮ���TG#W�Io���6N��c���ZN+6��	:)��r��p��Q>o:LWٛ�[k`E���ˉ�&ZLs8!l���=��뱝�-$��WE�}&�u��L��8�����;Ɵ���m���h�3yP�z�a��͢�[{�PsGd.L�h��.��:�m�`e����:F��L�lDS�ͨ~�7�/Z.��+Ӹ�;��s��z����ű�t(��K��;Lȼ��k�{�ۘ�wݝ�����=M�_|ʩ���	�@�x}ǽm�cEƶu�bC,�M��>M���&����T�W�,wh�y���b�H6�q,�њ�v��ll.����9ɡ�����ӄA���#��)/�E�{xvww<cn�[Qތΐ��ۋ�Byh{�TZ���|��?�y~Y��Yx�i�����h�,Wb+;ʮr���Yn5:�g��5�.��m�Ll�D�I��b�b�� ����j;��*�J��n�Y�؎���!;��T���[�ѯ%��s�s	��W��b!q�aG��4�I���2���-��H�	Q/ph�iu�ga�D"%��d�v[�˩;Fᖁ���]&�dt�;\��:f�g��u�2%���B��uql����[�_nN�V]�	4�V�U�$&n`6"��sl'�@�vk��.��{}Z���4����|���w��m�z�X�u�0j��q]<�^楃@�w���ҥ���eq��RU��u�pO�����y��>�ZD�_wJ�J�]�D㥭��o_�7�����R-5��#,?>���������[�j���T�6�Tv&bwO[t(X����%�U�׎ͽ���A��3Q�ϗ9]��,�]��efVi�Z��}��f�>��%��sX��P웱�q�.S�=k.���E���+,��1|���6=i�MKA�%Ι�
�x��{�5{;i�hϚ�eL�.Q{�% ��s��IlS�2Hz�[��j���#$Fv�fٛC���e�Y�Û��1;_��Ъ7C�!��6!MfZ&�V6���^��G<B��C�CK�^�:/L���i���Fm �5������������� U����mkmm����ꚿ�Z�kj�_�kmj�~z���o�}�;�mj�-�+fUL��[2�el�ٕS6��lͶf�ʩ��6�*�UL�̭�ݾ�Ͷf�el�ٚ��ٕ�3k�k3[2�o�S6�*�V̭����������o;x�m�+fV����fV��̶��f[f�ulʩ��+fUL��U2�f�2���Tͬʩ��-�5vV�-fj̫2��ݹ��eY��5�5fj�ՙ�2�f��U����3Vf��Y�fZ̵���j̵��3Vf�ʳ6�+fmY����5��6�l�US*�j۳UTͭT��S6�l͵T�Z��mT���ֵS-�S6�S*�L�j�[U3Z�eV����Z��sm�ݛm�f�T�m�eUS5��[m�*����fm��eUS-�ٛm�f���UL�m�6�lͶ�3m���m��m�f�TͶ�2�m���fUU3m���l�l�T��f�3[2�f�3k2�eTͬͶY��[2�elͶf�3[2�el��elʩ�l�ٕ�5�+fmfV�گ��ݿگ��]}���5�Ve��mF��j���?�{���������������]�����W������A����_�O��   {���������ڵ��������*��VUJ��_��M�j�*��m��������|��n�������忭�k���U�+�.�����j�ͫm�5US[J���m�l�U4�m�km���m�V���USYm��eUSZ��l�ͪ��6�l�[m�Ͷ�--����lͶ�mUv���Z���]:�����_���[ՋUUb�l�-���_��]�~�W���_6�5�����U[m�>���_" xg�G�ս� ���������   {����j�z�e�M����kUV�mUU���������+m�[o:����SZ����R�߿�����-�o)�򺺿�]�Z�m��{�W�|�檪�g�~�_��������m���<	 W�w�~����� ��������Z�������������_��W�x}��ǁ�@O��������� o�`��������nf7�?���_�_*��������{�M~}��mm�[o�o�]_���[j�۟��_�������b��L��儯��<� � ���fO� Ą7�^> J�R�DI
h �R�P�k!R����
�D��J�QU���! �*%%"lҪRT��U ��������J BB�U �Q%RUR�eUTE"���($�I%"!���̉UD�HR�@H��I
�Wl�UJ�J�DR�))PRET��QR�J$$T)D��T��DJ�P�E(�UPD�AH�*�R�R�5D�Jc�  c����h�[K�:uh��P:�W5�n�U'$�S]ڝt��S]�V�l��`��5��� ֕��m۠ �fEݣ�5m��!R��@�5R�"B��  Yaн�ZP�+B�ѐ���*�3!Fٽe�.y�B�iCB�
7�����P�B�/K�E��=i�V�6v���u�]��:�F���w�7wuG3�s]+�)����+N�j�Ϊ�P��J�"*������ ��wmR�4��λ���[v��n��v6n횡�U�Ӷ 
�\�v�]m��p���[�J��nPu�q��p��:��Za�;+%k��J@�(H���#���[S�ap�ӭ)ݎ�6�*�*�:��[�R�:�p;�j:Q�s�u�@v��[��� Zm�U-m��J���*�$�RA$�U�0^ 7bJ5� ��\�T���Td��v�SL�X�MST�Q��¨��N��s5U�49��*T:2�)E�)@�  c�:�TɃF�1�� 6Ս*"��h=��۵YD�`����u�ڠ��jM�]c���
�UGm/   f� PMT� Qab�5PmC S2�E -(�Xe��0�� zr�� �a@ ��D�T�)@�T$��%�   �����n� q,� ivF�Ҁu� �@ �0 �@s�� �WY@CI�w  �lȀRI"@��    ��� wEn� t`t ��  �ur�  kJ� @u�ƀ �����  j( � ��%B�K�  Ӄ@ {��    �9�N�W+� �1V  g%� ��e`�4l���7�"��JU@24 �{FRR�@ ��z���  ���R��  4�U�� �Iꔐ2�L� 1V�kA8�	M��H����$�BO'"s��eME8�)��*7n� ��0fk�����mZ�}�k[mm���km�z�խ��mZ�U�mj�Vݵ�m�3��p�w��<�w54�"/Ľ��-1�"�&�w�o�E�����,��S�%�-e�Z���wu��z��X�;�Drc��)4]��m��,��R�\�1�F�����8nЫF��a��,���-�q:�9#�\�V���3볭\�&���QiM*F�w*�ͼ���x-�زI��j��Y�Y�[���Pz`�ˬZoa��mǵ+fD�͔%k���4d�{��U���q������H�)�M+hd(����P�]�߰������w����4�ل��/V�oD?I� ۽�"�+�*Ҫ��+�S̼6V�D&��ƌ�ZK%c��P��ͽs	FXRch�QA��-��R�i)Z)e:�i��5u��f]a�~�[�YVAC��-�M�
���6�!��IZ�������-�vJ�$ڶ�1��pB�+rM�n��R��ލŦ��� ����1*+/35�3DW�$���P����p[����n�&���U�ayX��#%f�-eM��T.��Q�vL�m��*��7u[dy��L9� l�͐�I��(�o)˻z�ۅ�tL��p|�o	�1hkr�E`���b
�K��t�|�sd�v���ni7O�P�~j�Ք�*[�ʺ�M����uCf�K�QRH�G��Z�i��$�H(Rz�x�v0spA)�v�R[�i�jY�VZ����`7V���4R���2֖^�9S�*$�G-���k�	)JD��Ĳiu��(kPI�p�9�%�E�ٴal�%�)'�,]\�ؤ���Ij��*�N �x7`D�k ��Ӂ+��9{���b�%�"ӰLt�-��,��;x)��Z�ˁ�X�qo�@��\2���E������Ri=o.�mcs"�B����/D���+�^�boĭ �������Q	u�#r<A���:}�{�m��Ɩ����d��-?�-LXeL"�TP4m�&����af�u#$a-����2�
l�(�m�W6�������[M�6�vr��+�zv�d9�TJt�LY��/2a�7r�wC��W�e�3i@���T
��ek@4�{2	�D'z�@��"��\�1b��6\�+4��pXGT���o2K��u��L�{V��Uv�1�լu�k*�e��Znئe1!�X�5g�:���� ����n2�2��P���$c������L��|�33n ��Z���[�t�C[��JF쌠�q`���
�VpG�C@C���op�6�]�ug�����6��wn&g۫T��� FV�X1n���-H�bu��&I��k8�l�ܑ�v�T	訮��e���5Z�+vd�T����n۽�9V�`��5���I���ML��m���7N
6�k`�e9���9��i\�xN������0^,�J����"�P�y�h��%�&�W�c��1���VS��6l�V2�9��K�&2��U�cu�m�f��)-MX��S.��6�-���x�h�hܽ�8ܦiV�H�2�ŵkd�9/0J+i��I6f�n�|Y��&��젴�LJ�(�T�"6,��hh�V�k�Lb �H���\J�BU.	ᛪ^�{�����SI�PA�#T6!��'��`!��E��)c?8�Զ���#x�E.�ܚ_���-U�m+Y�V(���t���4�I6�Y{NU⵲�6!��ݨۥ��Z����[3i*�`3������̎]��Z��in�v X�.�5����w@���8��ݠ�ib��5�^�XVUM$CX�5��ڛnf/��Iu�(����<�J����w`Z�Y��6Km�����f\F�Gq�n��U�wQ���O.n�<��%�֜e5� 2��r�G2�V�XN�^Y�%s(�KV���0�Fcuq_b�I����k�z�yd�Ҳ�]Y;n���G5**r�R��!�-׳E�6���轱��کm%�@�v�~L� o=���7hי@�B���N�w�$�S!�u�+9hz�f�a�6�v�^�U�(�J��-�L��!+q��.�|%��b�	����O�B�1��0��Z�v����Nk���N�E�Ռ�;yW*��gs�B'u���Tڰj�8��q�5���	��h-Y{@*Fֱ��aK�8i�l�paڇ1��-f���X);��m�y�K�~�V7yHe�7��t�B�$]-b��T�[б&/i,�;E�b\��EZ#S�i�;Ur�M���dŖ!mZn�E�6�s2h&�m�ɲ�y��N\%J�^7�nF�C�H؆�~�+I�
��i7��QoH���;(<[ELff
��i�]m���B˧Y���n��s��2�j��a
�6�T4�A�w4�-�mH(iM��/"ˎ�9B*��1Mɗ@\p	�����kWA"/���.��`��4���Ye�b2滼b��+U ��m��n[��II�V)8V�ˈ��lm���9rVbG Te�Zr��t��Q��!�!E���6�ݡIb�.�q�y���
:fh�����W��V���G��a&Ր�x�׃4�x�N�, @l��1���ۺ*-VG��
�*��|1j���[��:s�/i�G�K���l��J��{Fa�"4�0PC.S������BY&k	�X�bU�F�T�\�	N�ca�.�M�x��BSFb�nd�����1��@�����6��u2��R�����z���ٴЇD�8���ת��^`YB�;W��ҭT�����]�Sr�V���CK� ���LF-l�,�U�Z'f4RvD6d�:�6�e˖2��6�h���FoEf��I�Ku���!���C*Jf��[TԐ/��۩@Ř�N�.�V��7E�["���ҽ�wY[E� jS^F"e]���ulͷA�佬�A�!eJP0�	.RݰlnR����kn���i�')\Y��%B���I��Ct*ǹt�K4욶�š�
���Y+r�d����f��.܅�5-TVwbf��+qE��Џ3���YjSא�e��m�H!yu�["vr�"j�rĳC{�X5,�m��l�Beݪ��� Z�]e�kH��,��-�qP�"�b��::�fY�3)�e�?EL�:�^\94���VXY�kD�t��[%�t�+f��5ܗX�9�T���7���ͷ�61ޣX��֪��ii����s2�$�:���V�n���"Ԋ�ʹ"Қ���f�ԫpP�S��;��Ra��gC7N�¥ܳh^*�ߢ�21WX@[��ӟ:���(F*���V�u�Z���w�@�W̹k7-k ÓUn���ٶ���t#�`7�v�3%*6;���81܀vv� ��1=2n��7�
�&e�I˳5��Su�Re�a��m�R���m�M�)�݆t��f��Yxt�&�2ֹ��	n�.�R��E�c@�vb�h	z�.k�4h���6����sQ�YMT��0V�b�k�l����nc(�J%�z%n^�˲$�ܬ���L͠�Tz"�2�L-�W��ɟA�ҕ�ػX�Ο�,{ �S� �[���o"
�;;/i�
�`M�Fp]l���0Z��"�n��-��d�f<����
[X�Z$W��#�Xi�4�l+FY!�Y�+i��eGc2`�����^�m�h�j*�$�O;��[pB*8�wn��˗�{��D6`�bJ9�iЕ;���k+A�����(��5yB�2�fmi��5�QkrV�'��2��;��M�3c�a3FF�3h���U��XH��CJV��q�q[Uz�n���;R5m�J^��&|�N���i �b���){n`��'ț�V�f��RÉS�N�����*LM�6���$�Kmc�P��&R��V�gu`v`���A�I��0I��k+BU�tP`qT�UҰfb�ʫ��9W���/[�g{3��������C��AlV�6�b���+p)�j���b��������C0J�L�j�22*��t�9Sw%���nQ��E:Ҩ��I1Y.�Ǯ包*�ubhp��od��=%�QUZ���o�ɦKcm�x�t�{R7 I,�L�������U;����$fV
J�i�bB@,��E��.�;&�un�ë�!��+������4�)�-e�,\@1-#j�*�� *� �7]�,*�Y�nE��̏BH<�/U�z.ٰ�V�\e^줞��㬱�����759��+HE��!*a4����t��457d���y����X����:�n�@vo�V�),Zf�ԪՕ*�jY4^���A��-]��O�� jaR�����0м���ݶ�6��i����+E�d�M�r�0	�rZ��PWI�
"�+i�Kf�4h%S��ZrI``�����k�0�+fɂ��m�oP�JU�8I��Zb�fIGFҼ�{���n�4����M��U�<�a8����jv*ҷA�Ƿ0%K�؆7sl�)��D���OV�gv���kp=ei�H�lj���@��n�,ױRT�y�o KLd`KkE�yz���PF�{�{Ra� ��8Mx�X��+T S����1[Y�AkL&Fn,Y�'kS]%�I�+0�3���ѭ/%lƂh������}�H��n��u�Z���4�4Đ|��-�ẫ7��%��\54���.t$PׇZ[��Z��+�w��34�1�˨ªj�{J�Uk 2���U�ɯwU^f4�B�Rr�6���ƒ6���f[n��R�ôӨJ�2�M�ʫ�S��6���>m#(�(	hp"v�#IJBZ�7�m�`��H�zHD<��Z�G.FH���ѩU��c-k��w *\fB���n,�ݡc^����v�V %-��m��g���E�*�
�PJ!V.�cؙ4���J�A�ZEV]Z�%�v#�f��,]�[X�e��X[���vQ�&c�5�Mo]��@l)�0��nܻ5���I���i��
�tF��+KU-8�TֵbF�e����6��ٔ�jN��1��f�1�~(]�z֬���6�&�c�#4VbYi�s3+.VFsi.MwSHH��	�j�a0��9��J�E�r�zMH�ivuU�Cac�"K���a;"���y��P1���-���O/4KĢQTpMy,�V�uq
7�F^حJn���J8(��[���;�`���I���m)؋0C#;2�X��h��1S�WJ�5[�u�ĒyYn�;�t�@U��A��n�S$�����D�X5�$J�x�阊���Xr1I�釵t�ڽNJW7���U$P�r�ݻ[I�+t���3�ٴˢү|VB�V<�ۉ@�3L���`����۵��H[�S'l�����E��Y���̭+E��TfXNѼ�Aʗ[i�n�����Ǧ<�,2�m���0�z)��Emn+6X�X�Pn�ɀ�@��XhV��:���u2�7^���u$4�(.�Z�g6����[[���&����a��Lݭ�هJ�!�lh�����e&)��� ��[4�����qb8��Y������y���5x�
	z$�*��{���++%lA�Re���]G OtG�٫D����{�^];�*��!B��5,�I���Ի_�+�n�p�����a��/�1E����sEi�4�����}�(^G�n���ͤ�M�W���6���fF�>9p�wSc�u�S-<��+u���+:��>��#���NMЬ�F�����,�a��*K/q��Z�y{ Rͷ��{�r� �u�a6� �u%�Ked�ƶ�&�7E(�q���
�tә���h�����)L�X��dB���Awd��lǆ��z�5c^K���+X�ܑ�Ya uP�*VDX��\%ô�ȄD�������S!��W��Q(L0��x�X6N�[��n���Aj��ú��#ʔҵ�&��f��Q���ڢ���/)9e�՘��D!L�-ޱ��-�{Z��ŉ�*����0��n��mL���I[Ŵu�=�����Kk U��*=�i2�e�Y�����bB��L�,��ʰLx�Դ��ͪ!�����
YCu!y�Rކ�{�MYj[�Me�lК���X#�B3Q�T�87sJ��[Gt�v�p7i�-���6�_.ݬ7E^f�F������- ���$R��[4�K
�! �\�a+zMM*�f��HJ<MS�k	��a�VEM1��mKB���JH��)������t��F3ki���3w��!vF	�(kP8,Hޘ�B�%�1ڻ�ݔoD��wW����XE�ZXN�4^����oG�$l;��w,��Px@�1	l��*�8aӸ.k�6(�76$������b�hsfm�F��'����ZsVݱv��GC/Y����cWwu�%��;�M��ȃ$J��7WI�{YiPW1\����
�@G�&㉤�9wsN�Ww4��	��`��Se��(�G��F�+[H�n���4E�xN�2-{�
m�������a���ޔ�-Q��1*`�_�n�T�A3.�A�� Q��ymjU��>՛ji1W	�̰t͈��x;Yl�Xҷ�=�Tqm����5bڦ�m7Hl��������T��y[�h�:䧷m�#�m۴��*�-![F$�$�	�N��v���M�!�3#@�4�F�N��QZ)�.����R�'U��(���a̼���r����̷	�x7���˙Dò������iST�{�
��}f�蘣�x�Lv,�4!�m��؛z��b-�mU]������W�sls�ݝ����y�.�Zxn�}�p�=7��Վ��Y�ԘA;s;�㗈]����]���l�(D��ܞ �&ޝ躼��Lյ������IpC���Qw��x����U��v�G�19^��,��ͣL쳝��K*u����{e`�Iܼ�y�n�H��䴫8��J�ç(��	��l�w��sR��H�۽��.ٍ�e���F:�WL�s���ͻ�;����Z��'��5��m:��!*�r�Wl���q7�J\�a�.��R��&Q��7�_a
���(m`��]��b����^Z)�7�ӛZ�-PMWe^S���eƻF����,��e��@�ec�7Joj`iN�閭�oh����}�ݚ�>�b���4�_pB��EPt3�+Gh���!�2����kx��aEɑ4ձq��.����T���ϰ�Ɍ\�gUڇK��
�}#[׵���/����h�݇WC[[�o�JC��A��+�T���x�:8���W;�Z�j��1>���qo,�-���N�mQJ%%[]lQ�[���^���̝G[�� ˎ��e#r���:�0��d��w[�9Z�7��JT��=[C3���첞�)�t��`�u�]z3��5��#h�%�A+�iu���j���K�ýk�m&�m7�\�"��"�P7����tMd�5c-���`[����9t6㮡��{U4�������k�s"I��fA�� �%VH�M��ZV��oVs-��HP�>��j�2ğ*�����N��qh�|z]��np�P.��{��f88�[	�H�Z�ˮ[qf>2�ѵI���)+�onܒ����U����2+�\V�H����A���0�&�ݼ���\+�WG(��=�����	�8��*7tz>�R�n�c6�T��1��qD1P�mu䧭�r��`�'�W��X��u6k����p�LY|���)�Q�YzR30^<�*lfk���+'^·l7��Nu�}�I��FY�W�"�;�W���E�1+����=2����D)�Dj@-]]Z�rBv��Ѯ<�8�ќh1�LH޳��]��#Δ�w���-�w���V����&������$Y"���i�������3JIM�ݡY�)�1�)��Ь�IT�����E�Ѽz�[�f+a3z2�ˡ}�Y���:��[���3s/Yژn)����ʈ��q�%��7w��"�u.�24@�[U�4Te��J�Q����g>�ܼ6���K�eZrv:��Q-�n�$ c�LuZ�(Cr&H��mD����r��~����p���0�R걛QJ�Nek�Cm@���dS���mX�t�yx�#LkcQ{���Yb^�S[�&HW�;I�0ܘ{E�t����[��k��C����9u:�v.��w�\x��=Υ��	�d��m�'�ͮ�H��k6�!�����2Nrg�J��z�f��Y�x�פZ�6����]�J!W2��J���C�fAI�ۢ�zтEsy��{�37�!.�e��>��8�c.�9�i�Ϛ��\hiT�uJ�ɶ�����w�Z��h�I��B���,�� �7Y���{���
U�VYQ�c�r��������ޜ:��[t��w�Z-��dgN%x��y��Du�ϝ�\�#@�7��#yo�e�;m�Hk�Y5�@���z�u!�گc�n-&lI���vҥ{��j�U�Gg'$��K��u��\7	�)
�S�/_,��'!H��7z��|q y�� �́ႝ	o�[�.alK�d3]�j�-���XB��{.��F���r��H�3���p��'��M(��΂ҧ��"y���w/��ٯ#&�kWF�L���۷��h��Q�0T9�Օ�d��ɯ��v�9���Rwf��Y!���s{��4}Wp'��s5�$�[ݣ�h�4%��N�ٲ<IJ�
��GW:}�[.M]f��Y*�ý"Sk x����C)�'!���W\�oJ� �}�m��Y:��̔ݬ�	ot�ɲ��kqN��n��H-�@:�'6X�ۂ���!ѱG���N-t���̓e�i��.C���W���@w���vD]n=��*�,��"�Hͫ+[��Ԇ�A�uM��j�s��#4)#QΡ}���z��9���>��p�='m����qkYt������fZ3�)�6)4��ҹ>���	��㸷R�Ko���]{������S�~��^����{i�53�E��z7ѻ�C�*��:"ߥ�`���XT��1&���r��S#��j�]�w��]g]�.;��ۑR��:s��j���O��z��&dot��r�",�H���$0D3����h��r��v�E�E��Q�7���h^�J�\�Q��fG�us��]p)R�]��]�p��=5;U[�K�[S�(W�]Z��쮨>�-M�GW�/QOd�5��ģ0$gd�[Zb��w��*-�폳�)�s�u�bU�t��]�l�:�}0�*��a�pخW#+��,Qդ-�S�Ŭ�x�[^Vi���:�SX��r��@8W61.��z�*�ջ��/O;]��̜v�Ft�S��o���h��`��z�޴��p�6��	�n��E�ꜹ؝Ԥ�;�en�t5�ki�LA�],ݝ:�{2��o�J3��PѺ�,Nwe�����̤�eֵ��U�&芜w0�L�9��eio��s�wR2u�E��0u�,W�>���DN���!ٓr�;��R��IFLr�����V���/���풰� ���ݺ�=ҸCޜ�5�+�	�"���� ��8;��XV�/���Ւ�G:�Ν��f^�M�C�:L㧻���J�鍛7�d��d�������{�+�x<3Ur4���缱��x/Vі�c|�3 ׋����6�)�\@���Ru�����)Zye�x���O��s�R��1\v�G���j��K���d�U�V0vb�]J����t5e��^Րz�<b�i�Q_b�z�gh.�^��U�{.r�����ff�*�%o�4(�ZZy�9���`nhQ��[��퓕�Η�l�ܮ�X}ĕ�����S�u�ũ[׷�7(ebxa�.��a���?�]>Rs�`���פpV-=3�� Vu
fr8����)6rи� f�z�2r�/,�s��uح��_�LmZs[�n�ޒ)�w�:���d��S[��&zﾹ�lX�r���vj�v�˧�Ꮣ��m��8�ӈ*��W�>�ԋ��5sYh��L���G���JMǓ�p;�B�r��Lk��Ĥm���}� �>�Kn�Bn8��-�V?�q� ��:K��؜9ʗX^��}�cJ��é�vb��67z��յȷ]�J���'��^��//1\��S%��J�b��L}G{r��[�dU��ԃ)Wu������&h�K����%jj�ck�pLYG��'P\ok�gC#E�]�s��d�w'1���p���,P�ңZ�ojmm[Y>;��r�(pR�F*��G���)��c�&��:^]s[�]��1�1goK�����ѐ!EYw����9�Ju�^�q
yWé��!0]�SW�^�%f2h���U��df!N�R��Lk�>���@(N5�������`V�Q�x]
\&�p[�R�WT�h��i�eJ��I:�*��Z�T�&��u��q��w�g��M�<��_S�{��]��̫�z�nb�4A�����`	o N�ݢ�]ǟ=w�ΘjlU�_1a<|�f;tP�mp�����%f3��ޗu�7���eDo��:R�w^p²k\�aF/�w^�/�6^sķ��9c�xh��8(�L$�j3UAA�KD�����/�WN�ҏ)�%驲`����v��2������U�N�@�����NР�bf!�,���s���aZ[ç�Q�x����z��9Gy4��̴k�u_3Z��@�W7��$F����2 ���̾��Ѩ�
��'�CE*n��:wV��t�v;�MW׋:��(\T"�vvP|l��r���$l�˕��/_���5W
{��1��
i�ڛ��[7ش����}XXw�6ͪПI�ԭ��Z�Sv�{��E�*c%�T��@��ϸ��q�癢��Mr��D�
co�n����{9��X��Qf*�|9���7�����%hť×˻ym;���^4椐ȇ]e�gָ
��b�
8qJ�*V�u/k�֨P�U�gu�9v���Z�ܫ]̝Վ�h�b���W��u�/_G����U�=�Z�9e����z�@ɲV>L�V%���6˓i���w-���8"��\�Pf5�c��]]u�/��&�\���]��hN�x��n	���`$��Q^�Q��^>[F�WnA΢��Ƴ}c!�9��V�����ǉ�a�ך�Laz)�;Z Q"@b>��y�h/\g7�4u��xP��]���(�0,�i��ua�+Z#TOkm�Ǫ��{*�L�+��U�Sy�+e�R��e�[�av�J'F�!9{�f�t�$dMM6�N\\V��4n�\:B�WU֒�к��a}y���S�ji(p�m�C���_��mgn(�ޮ���-�s�$��u�@ڗD޶����
+Z�vj,���o&;�Kr�\"�)�q��*�8��g�[��d�U�M'e��(�W�gi-ђ���|���ﺭ[݊r�	��"�{Lwp*ܩ����Dm��v5B�7�3��ݸ��0�?:�*92��Y����҅^�.}6��0�m fe,kp�u��x�%:p-]��z��8�az��
�f�ٴ6�%�v��Mۗ(3}O�~��l�*��rf��K��Ȇ jO��ܬJ���&��,�
;WQ���F�>|�ǅVZ{�F�f�¬��'z�8�d\���8�pvj����c�l�η2��T:¾1:ӗ|�h�*��6��<��C7(=���@p��Y��n�w�5���x�ӽ�B�.�kɸ�WQ�#��:wPKWf��9�j�i\�Z��T��n]�;Q����7t�~n\Up'�%�[���f0VY�;���'xz=(�9k�Su�(e��U����;������42�!k5Q4��y27��O�^aԖ͎��ۤ57�e�����
�.�h�r��':ʛ!�W:���K�)SĞ�tr��-.b_A$G/g0��-T����[���8����B��v��9j�d
�mn�~|5w���̟en�H3���5p^w��;��įH��y�0��#�j�;� y=E�d�6k�nW����w2nS�S˫���]Y��M�.̚7v�uƅ.監0m�ls�؝�8�SJ��@��ּ:�%�	��PSݠ��9\��0>��/Sl�j��U��>+VۭJ��;kdW���ֹ���M/��ݴ]��5.V�8IH(8��<�UΏ����M*���R��z`uHํS�im���V��|i,�3~m��`m;|Z�3��F�ؾ����q�Ѡ���^+�g	;R���ұ��K�6Z��&t�A:�"&Qj����f�Y���鼍$��\V&껕�u���^�/e��㹦��Z�l�
�%�=c+R����.���"�j-�z8-�#B��ٓ���|e�Qvհ���+��sj�dKs���ͫ���}NM<��as����j�i�\ws8pɧQ-T�2����]>彥]{�&�6#4�x�$*uN]��#խ�5';V��R���}����mπ+����鋡�:�h@f�sH�m����Z�W��X�y��꬘I�:���[�LF���^f�U]$�CI�X��|�gc:�L+f�]7��e\��A�t�l�͆�;���\�t���k�ީ]����|G=2D �'4`�,������� T��FmS�P�0_���N,I�Vۋ���C��f�N� fL�!���hTOO$ͧ�[�� �0h�O���Q��R�n�V�d�|хu�*v��I{]�/���t�i�����T��r��7B�[XI*�sϊ�Y�޳��k_j��H�n� ���`lt���+�m��]�õY��5��n03kyϜCj1lS�s^�)�;[�"�Cdٮc�XvE��Y����K|V�e�B��;���V�iҨ�tqo�e��}�'��CMsFQ#�lwP�����|�@q^�)�PM�ۙ:M�5qb�P�G�1�	5;z��I���g�fnl�E��˯y��n�^�'���Ƭ��/�!��K[Չ����pR�'��!0h��+�η�+4�l�[��;'qK������f�̫�{zMo�ZT��W��Tn��e������,�hl�Ϟ�L+!���|��b��h�:�@�U���t��f�s��؇�;"���H;V��	�������c�Csf�HjTm�!y�J�y�������V����{kq�V��=��3�����{�bJ�o@��#>+�u�	]�ۄ6��+6s��;���+/z��2Tw�����((5���x���� [�(V3��c��wF�n������X�:�a%]j��y��ŽH�c^[��AB7{x�&���:/{��ZA��b��m����s�x�y0;�;��)s�-�q)����M��J&�1����u0<ɗ��jh��Z�H���`!X#Kƙ[�H�K4�<n�'Վ�_Zo�p��*�'VB�f�
�s�Ew�_^j:	�> ��bO�,�yh��W���g�z�)����f4>+����;��7�t6O�w#�t�*�P�n�+GDt̑����x-@��5ظ����iJ�׵��v�NQ�v��v�p�4*7���W(�}ۛY�c2�O�Dّb����&`��30f� ��0fog�<TOޢ@�x~rUqYj[Ӻf�X݊:7�s�F����sJń�.]��P<��S��X!'�Zs4�����t��q�e���>o*Y�u���to.<���M��K0���ȉݫ;�	��J���n���ECU��@˃���ڼ�x�VPX,aMY�OEn�]_\��g�-�L��ԟ�)��s6,��*\3����%�h!�p�h]%|3��ݮ
�A�n�]�A� -2�Z�w0�d�ju����[�5���{��>����f�It����a���ㅨ���$�[�A���L]q5t�H�<���Nb�
P��"�S���K��Q
�����Vb�Hu�Y�
�a�r��{o�;Js�[Ƹ:
c�7 £s�[��"St�S�h]�oj��X��V;ku���	ї��-;��0%�8���_qWV#����\(��ٚ�0ۻJ�̈́������}f@�!GgK�q�ʕkW
zo�]�Q�=;�L Q܈�Z4�׹}>��E,�o�ސ�T�۵�]�4��L��\��� �\B�l*C��|:�l�$��S�,q��+3�M���vx`��,�v�׻7/��+[uc[uc*��qQ��u$	!ګ',�Go+#f�͡�YY7[,�	�ƨ9ޑ$Y.$a����	>{RQ7�&ees S-ܨZW��.��M�y�.ȡ[�������C0i�#�m ���2���$2���1D�m�4�ӫhe�6'Ī��x��1z�VpE�s8�vfΫӼ�2)3�ӵ(�}� a�F���T�­%�R��+ ��#7��ͮT/2ͮ�!�\���-��yx^
���om�� ޚ���B�����U��v ���;3�[����oO�P�Ӂ��D'l���o�*W3s>o)���Oya�Ѥ�.`�t�0�XZM�#&�Q��F���>*G��i��f��b��Ư���!��pI�q�H�W��xgQ\X�
��X��Bg�0�^����kZPem+�[���'� ��YM�ysD�'YN���mn��"�]�TjV���r�����5��C�W8&�n>��Lέ|	�hh����%����8��L�P��a/��J�����J�bT���=���� {Dj�٘����]Jjq��2e��t!��#�e�U�lZ�_e��̺q)��s�4Z�*�Wc�����Ͳc����������d� �-fk{4�뼙�>�lg���v����Y;������L��0kݦ���x���ri���X;���S7�Ci�2�t�5�YJ��^:Q0��)�F+��'q]��"�\+��ٍ��΁�g���iSJA���/4w4�
������'Wf����7P������i�zL��=����z!$�X�R�}���L.T��S�|�8w+�34��}ܞ=�y��e�]�x���`�M�&n��|yU�5X3�_C���kqD/w$�U%FU�����p�J� ��6�i!Ap�l�nQ�rS�W���[&�ض���"����eI�n��ܧi���#� \!��T�:����k4r���׫mqx�����Sq�T�~N����N��v�t6�Z9R�IB#����Msf$6��'me�S�q���:	��-����k9���M�8Ո
bs�;k�S�C+f�Yu�]DyCW\�M�1�s�lw�a���kәv#0ɠA2"�sw��Øf�o%�����T���l�w�,e6.wt�Z��ذ��|��E�ADc��[W��t�ӝ�X���/����pּ���M�}z'
�-���F�j\+��RWG��l�6�[5���"5� WT��Z���nm�E6:������ukH���az�=�<��F�]�먬c�%���{J�9�*&����q��]a��l�k�-��%s��2+�6&Ό�MG�� R�ʹucN-�|�7y�{q�8�\3�|;��'E6�#Ժuޙ!B]Dj'0n!����.wF�����HJ[��XL�1^^f���߭N��% s�Xr�-�̷)��>�q��a�Z�:��Q彬վ�KzH2�Q�!�v��`�L�w��.R����-����29R>&%:��|�\+y��W�cUt���+(����C�m���s�s�4AxU��K����ĳ�����8���R4�t���{J����l��u�n����o*l�p������C�j�.8r�pφu�Q��n��R�r���묮O���tjZP�,�X�w49q\��7��YY܆��;v�!F��r������E��նV�l�M�t�2m�oWVw)a��J��ɼڂ�+��z��#��;qc΋4��L�Y�[)(
��YK9��1��s;��U��hW[iSB¨���Q����;;���yܪ�&N�)Q|�%9;�\���5r'	W�=xS�Ld[��U��(Š#�ܜ�|��p�5��Jӄ�/��[�P�/���f�D�d[L��V�gE���,u��V/0rh���Z{Q�c6��2>��pٮ�i�$�*}�#Lߘ�w3R�#]jn��˹[|�}L��s^�bu��a�@��!�,p
1+Ac��ˎ��9��ۇ� ,�˦�΃]e�ީ��s*Vⷅ����(�n�\�͢
��Ac�J���*�{�lH��#)FU�ؔ��#��}�-0@V���I�Z�����jX��]�۹.�3���l�Vu�Y�Z�,_I���)ꕘ�M��E���ˆ��Vl��Tz�*��@��.Wm:#j�m^�,hF����x�5���b2.��Һo��G\��zQ����Ί�{�;�J�<�:��,�ˏL�G�����n&Յe���U�Lw{b�Lj(P&n�[��c@S`�w���8�`Sm�.�P�i��-��Rh�k�f�d3��Ǌ�}��f�ph3/��y�\�k��IfX�,��*�����ñ�uݖE:�񾧂���^ ptJ�q�[�ѱ@|'\X��󺔨�Z�۵���*�;��������X��`Ap����3��v��t�>���omq���&a�n\�kX��t���JV;S}֌�u�(p�{����R����}�Л�uv�U�E���v�m7o)9�,�y�p�S���`��%���V%���)C",�EHr�]2�#Im;�:��U'"��LD����M�����B_��r��؞�,�kc�=������H
�[��.�'t���^�4u���(��^1��L�+�U'�9A�CIb�8jQ̸jT(f�'�$�~_'��m3���d�nֵq���a;t�sU����s�y�,]��7�6@l���-k�.�c1���ݛ���❅���:{�Z�3-cWSF]�)��cW݁<;�wL�6*wg�m.��'o+����` ��B�mK�$�q��X	ɇcy{�n�J��K�}�8�
[����w������L��|�{�&="K�X1nmq35�B�f3F0�U�gE�̉^�����}b:�A;�t����*r\;V/�ňēAi����qoI��������h��}��(}mRl��mgT\��b}l�wN��bՀ$^>�9�W�壦��J��%��R�$w��6@�S��
ATT�؟
������w;�6/���j[���g���ܺǱ�V`��ܨ��K;kTOf��f�<N�%՛l
��9.r#/i��	*<�\���Մ.��Sg[9�8T��0��tM�8;���ݥ8�$��u��0k�6m)aV\�N˨rB�su�r�x��X�X���PN԰��0 ��`��V�����T���[e���>{X
��N��4�m<��9*�P�pK�ɭ��N�g:�S�8��v�O.8�!HU.����W.ذ؋ ��X��Z��x�nY����-9�)`�b��$�̄իF�I6���L��t)����k�ZB��v��7�%[�x#���\�8L��e�q݀�6�j�.G{�,���{��	���7viQ�y�y�vS�w�b8���㗻�&t�����/��OW�t� �dj����
�g9x���P!fe<oI��K�u�<Q�ܶ	�͹A0r�T����q侼y|���wK�6s6��4��#+tc�bjW}6�!�{ƐL+A�݊����⎷c֥%��^�3�h���V��Y�z��"��st�Yo��\��Cӆ�o^'�wV���5��\���h�����+/[�]�3ih]�R�I{���/Sq|~�E�y�ʻB=t
��>���:</R���qaiʫ�湙WO��Sj�������q��[]�U����.U�ާYA �fn� �zїF�؁�u��2ȳ|�x��u�ݮ�.�<�n	�����
s9u��4K+J���u�{ЕolTʷ�b�7|c��]K�U̢�n��G�\1+���ص^"���vW� u ����)��t��m7;1��}�=��x]��52goZ�:�ܠ�	���ـZ�HZ"hތ��4���V֎TV޼���,��}:���ʱW:��4pcz�/jn���9�p��a"������hd%�crZ�"�v�z��g]��.TӶ��i��ͭl\���I`�dU�rjS�c5|,���.;�9�j3j/T��مεr� ý�I�K8�2�kRd5d���yn�Wn�95�m|���Uq/��'	��ŗ�w�ГM�٬ɝ`I���ԡ��nMBdb��S�7��VE�v[�b��n�7�XQK� o6��F�h`���h�V���'3kLDgJ�
B:��)�g7���#Eݛ�i4�v�ؾ��]���W�z�jV�����;��Y�<s��_4Rtu�5��]!ُ6��HS�ړ\xX�<"���|h����Z<q2 te��n�f�C%	p�0a�V�����[}�4�M1�	������ ���W	�8ĹA��/��[h4��涔����de��NwՖv�p=�-��Q���OUuL�g�I��5 �G9��]�K�<8iη[\�01s7->h��RS��zJ�R$��*��B��$.��v�"�N���]�֫�g2���kGTWE���x��|YYʎv#wL�U�X��C��ʑ�=І��o;XtȀ!�Dr��Y"�:_�96�b��ʭ��O�MF�P��@ �]�tr��,<&\*��&�t}�T��8����k��*Z�$�I,m�cy-(��>�p8ezh`����ӻ��mowd;U\h�-:�Cq�iK�8U�ӻY՘��X���[���L��Ӧ\����	Ib�$A��i:�[X�/{��P��*��WUU�T#,�6�q�����B������sͤ���>T���i�,��Υ%��gF��g���ڣOB�3�:��MKb����fY{v�7�v�A�y��� =�+^4]c�7o�*P�Q�ѭ��ǔ���@&��y�/��1�s4�/^�],SzS��h�	�@������ˬHS<�6�Z��6*U�8��Ec��Z�7�LdTy�;���٧��f��(�PA��>�I�ۂ�B<�f��i�-�7u�7M����Mm��"�Afh�JA�Z{	ڵV�����Q��k�V@��:����}��}7��ݣ�%%��뽜��Xn�L�
��at7�T͡���J� m�YUw���(�!>m:�gZך�0���VP�53YH�s�J�Z�J0;g;sH��H�랹�ɐ8�6>ˢ;�PPd��!ƻ���q���ܫE���ܦ8Vwma���]\�#�sQ꿬����ٓx���-�a@���#K~�r�ѧP��mlh'��n�v'۽,r�S+m
h�M�^�DA"�ip�ʹ�G�*���e\v&W��v:;�(BWư�a��]^C6)Y��v7P�^����1�'&6q�����Y���9l&�v�kսG\噵��s�lJ�[��Z˩y�CRb��N��j��-��At����Y�\���C��i��뫵���C�]�1�J|��x��koj�=7h��k�]�tY��H�����(�`�AUݙ�B���><F�RQv{W1�Y��5 �cU��k�J�Q��R��bq�D*�\�91A�R�u�f�u�or�Ĭ�O�1V�Vs]��7�u+:e���d;hs�_�^]K�$�]a��^3\�9�vzя>=�-� �Ykz��cpdЯND�h��U��ƀ��κ"�w�k��5����i�b֝�3�K�nm�*P��4Lo����u��rL��3^�J;ջ�՗;�T}&n݉����ʽ�q�nw�q�ru�V�5��T��A�������r���}@���V��b�mc��I\ƍ�h]]oN5�(2�Qk%��A�[x��i푐5��X�N.���[��0Lk
�0I�@��B�+��z�
����L'� \
���[�Tgƴ]�Z�R�d2��]���O]kU���������C�29vcə�5�SZ�V�N+mX�s~(��g����j�jvʛ]/N)�U�ܼ�E�����`-�݁� �،�����L�w��\cyʻ��qĪ���@j��ꔡ��d�]Q�η����c���]3}�^ �#p�e,юP���$ҽ���E��WV�t\;Y(�wD&zG��+Ŧ$Ќ|+��5!�ck�85��[����l*.�$M���z�L�
�����;��RUm�X4S)M���9W0,V����'k���z�\�5��[��|8l�����Oa|M_&��|��JTN��Q�`HK/p+�{{��C� Xr�4��%$s��DV���ËŽ��TB��:��SM� �IX&k��������3 �����Td�V�fcIE��̔�I���$�f^]G"�Mi�D9��䫢{�u@�[:v)wՅ�n��L�x��3�=��/�ӳ�rR<�-�����ݓ��]��c�:�v����:�ޢ����9��`Ie���]�ğuIuan�j�q�T��.�X���j��>�1;sn�{��m\ʉY!�@ـap�٬�tu�����(D�r����e�W#����Pw��]���4X��n��]��zV�'kO����hK�f�òR����V��u�:Y��}jQY��
����鵐hOh��u�m�I�F�V�:4:��f&��8���h�6�k�(sӿ(1��*�.��2���t:](e&B��Í	ed*�7Y�6�y��w{�`��2���wu��Na��.:�z;(�]���5��7���T��0^�BWZ��n^����ő�rӮp�����X��y�����'r��mD��S:�j���]�5���wؙ�cQR�p�ss��԰{:r>�Pڱ���yD�ǯz2\�R�)<�󣌛�����V<wJ��:N��Ս,Z���\�
��ln�]�����]���]X�'�[xS�|���S!�_]j���H�Ȳc,E�]/�6�B]���m��V[9��sSz���g2��e����w�����,Pv�h�Y��@}ԗ�S�{�_JV�n�; am;�?��޾�;��߿�h���I�d�nQ�"�Q�	�H�Ѡ5"F��%�QRh��4E&(��6#@"���*,���I"��Ё��LY)(��Ũ����,�H�d�h1�cFK�,Y�,m��!`,EI��FS�Y4m!�h�ƋQ�Q�l�Q��6�ƊJj �I$�4��9�(�$J1�`���L*M$wtQ���J!�JJ4��Ȩ(FTl&
H�bBƋ0�Q �Hd��"�*#Q�`"f(�%��0������Cb4�4F�0Hب��ZM�cl��� 
���z���>���H�	�\�����;L�X:e��+��*둝L.7�v�>��溘��ȸ�gV�-\y3�5U�paL�Ӻ���A.�ea��Q�r�P�	�5�M�(��fR/-��Ŧ�[��7�h� OV�D��DPF�7]Q_p�-����"��3+�V\@����?.~�%{S���P�II�4{T��Jʯ���$�4�Oe�^��c�������V�aJ��^�%I�zJ�K��.-���q�O6�Cz��^����t������ �e�C�W*؃ekNZ��Š�?�΃5�eCc��C�n8FG9i�U�5�g��t�Θ�[{��vn���+��q�,`�5�@��(<-9"���B7X:����́1�ekN��;O�+�ؾF�>������Cb����H@[�X�ֺd��f���D�A)?r�q�}:�<�"���N��vo�<b���c;�LH���RN���S5�bm֖IȐ�����p����zO�8$L�fP��a(��+�&��Q>�S��gy��/ ��n���۔�G~y1�	����#ג�@W��'��o�v�y}��(7��+��E�S{NB��t�󓗙rnT�zԳ�cf�'��u^�+�L�R���~%�:6M6��O� ��O9�V�R�v����-FQ�d3g�<:��vᲫ���D��ܨWt��c뿅ct�ڦ5�Tћ	�8�Oĺe
��<s����y�-4Fp��GZi��FGi���,���#J���F��`�i�\������]$3�^ ;�
#I����s��DL+u���j���{N�`N��q��f��8�ӧ�Y�����O���Q�ܫ:LpwknT,��"�[����@��r
��U�һn$%�;��<����DҰ��;k��%#����&�D���lN�ؐ,���>���	{R:�F��*�tB)�;2��Q��;�3�S;� Vs��3�{I�ri��\�%��ڄ.�j.N�þ ;�I+�|(��D�p�OA}�1�~
GV1�'��uű`�q�
Nh�U	S70����8��&��.Jӑ&8mMT.���{�L(�c1�gbģaI0����%�d)���ӯgd��T���l��=ژ�#ԝ�i38'��.���0�&��:��� TwK\)�JND �n���rΞ��z�h�N��vm{� p�fH�ͨxoW�y1���vsi :R�KfaO}z��w]�0��H%SU���9`�!^$9D��������58)PGa;�	�x.�j����'%b=ד0
gnK���9��Xnc�Ը#4��10�0{�Kw���,��3�gK�c�[�'�3`BV�ۻ���;'M�n-]d�Uk�(8�������a�Vc�Ȩ�n�uM
���̲���E��4��1Z�v���q��<�^�z�z��ǆ�k��$�LT�%�1�{s�_!/�n*���P�H�1r�C�u����*~��{��BR7,�j�t�}�����nH�)��e��)2�\f�9�d���`z���NڳD��:x�*�ǻj�t���W=QA\gM6~j�i�>'�T��d>?J�5��Z�C�燜�lM
Z�x�rL$n]U�5/�&�0�e�'�i��t�/Oi�n^��W\Ӛd�aa/�!;��&�L&�:��b5�)O�y��
�|���Ɔ��1��+s�R΍<�U��rU�pܩ��d�V]5���?HH�5r���]pQ��l�Z��y�-�|�)=�:nn�s�f��਷j�\7U+�L��H���vU�B΃Ri>�z�\WF)NҢ�`����耮T�I��1�}u���6��'�����t�0h��J�a������V�0��$�wL��it&Z����b��@��KVPilH��2���[����C�q6����+y�2gC��9�/t��n�z���˄TS�Jzqc��5Վ�;�7��K��<3��� �x�񑧡�5��AӹH��G퉰洔��F���"�f�����zp��S3���q�6�#DbN���@�؄���Z��e�����wnK��n⬻ nT~�kc�=���9��Ƌ��b���dB�j�}�U�B9���6�.�S�<4��5�Ѫnx�����@D�wCVWxl��a--]Hq�qN�LÇ=�ݹ��jK�,}¾���&����B�e���$�U�A��Sڑ��e��ZE�2��av��`X�FoE��twA�n���J̭>&�:-�|.U�+|�`{��Fmc뉳�Gk�и����U0;!�1No���n�,��c4�q0Ԕ!��ݾ�&�G,έl�5�M"���1�X����b [t��B����p��G�7��X���ռ�ep��o]x3p�LWy*���|J���I�J���ˈ�;�h�RÊ+�ݬ�),��7.�O{�G�g�pو-N�ἢQZ��c�U�۸L��|�K�uwb�'����F-���R�(������3�3�'μ*��ʘ:s¥����K]����g
��7����r�� q;�1`�Ժ�!f�w�k�9�]�h@��c�t7����j褋�/�t�ޚ6���7�M�g�n�Ԗ+z�҇Vg+�O*���F(>yq1W� �#���,�*�	dY��&�a㾅�-��D5�WY�?��l��Y�;�iB&!�;c>��(��@����g�
/<w��}��rDePyѸ�Ѳ5��\9�k䝤c!��3�~��	��'�0R=s���n.��uK@Ydx�P�]\���&a�8T�p��W�_Ř�xs{\T��� �e�D¹Rc��,����S��>���hX0��B��`VZ�E�b������|dF�a��� �]^�u$m�'&��:�{\�]����jDC��s�R}��k�2}��
u���J����� ��]3i�K�4sS ڭ��C��4(3^n���c�[#]O<F�Ҵ�7	Lh�U���9�N��t{���R��iu�6Ԁٿ�^]�q�I�NX��=t�oo��s8�35��/�1��<�n2i����2�]<:��Ϯ9�B��l�u̎0d��K�@�~��Vr:2h��]E���E�s��eB���1�J��g���Y�C.۝1��C\Q��\�a�{7EҾ���D�(X�8k��)G��$\7��xm?F~���q֣�jn��/&7��I��t��;\�����A��vJ2�W[��C�5����{��+��iѩP:���5�Τ���ok�E�WZ���צ9�Ed��XAv.�S�XX���	 ��'���8b�ҤQ�t����T�Dq"�R����F=ke��ֶ3��J�*��+�0/���!S������:��:d�C�}g��_=T���G�oOK�S�e�N^2�8�B#^�Ąq�[2�H�&O>i���ԥ(��욫��L�-��6��q6���0��u���(h��G�dF� C�ٔ��XJ0��B�1�O�w��P�n�^zn!���������	Zo�K@--b���-�j��n�z�k,	��6PbL�{;��-���v{�Y��=-!�H�,4F���9�Ot�Y�D��G;&]�z�V��*_c�Yˬ��V�E���}��Gi܇#w��ZF7v�,�^��:ƲG�Z�n��	�ވ�"��[F��26��C��T��}H��E�\�h�B�ԩ��y]�P�k���L�,3"8�0��?Y�K����}�۲�,tr�ՅNT�S��5R�p��?�� E>D*�(r�e%Å:4xy�t|ir�7��3maSB^�Q��;��P"���_'�t9�E�+$��dSɂ8ј\r���B*-��v2�v���p:�6�R��nZ�-�Y��5�;���&
�%@�Q�����|чhL:�y"F> �R�+�;�+{��s^>�q����g�y�CG�}b]:����nfu�N3�\+*�&+A���S8�}�[����j�oind�*K�*\�ԸŹ�� t��	�٤��a#���q�RPۅB�)*f�.���]Z@yXM��XH��AR*�.0㧚���	?����P�0�;
r�%�d)�mP��W��F�AB��<8X����ʴ���|���5��U�/<��:���~�b3���8�,���?c�y���T�C-y��L:W��P�j������x�Z����:�7��=��J|O�y����(=�E��4��}J����m{��,UW�`]��5�r�g�%o:��]ԉт��u��|�S�yX�b"�����Y�*�f��W�R��s.�5�*c��a��.t���9gD�VP��H�d�0�l�;і�c�:z��K�ֹeD��cNr�����LH]e�����݇���\c*�,�r)\��UEѥ!e��su���|q6��Yǉ�f�s�˺^��/�X���ܱ��R�4�r�������h�o����-t?(LH�ms�q7y��:>�*��4��v����V
�g9П �l>{.���k���2'(�����F*����v�:o������.�{x�WX�������w�i�jvcɼ�E�� JQS]��]G9K������ c�t�˲tj�f��ݎ�4����t�s:@��yq"�&�XJ@���s��r�qz����DՍ��C���g�a���i#�����E��i�A
�-��s$�|c�	���uN�Wcvx����U���[���:S6�cDp���iV�.EBʥE�I�Q11������'��k���To�<JF�4��[K���aS���9N�m������P���Lꪦԣ�dEOS�S޸E�=�Q�n��i=�H;��̺��hR~��:�CRJ�LXˁ�N|-�rja���W$�u�Vg@��v���>�s�j7esu1��	c��;yw1SfcT��6�y����[v$\"xQ����s�������];��mw�vE�S�|�5��t���K,��a�UGN��!��Hѐ=��,"9����.�6\�lͭ>9+c�VZ�������M�;#�t^�&Gle��i��qœ!��NR�y'QMZL�5����0�F7:+���#T�:��1���t��x�X�*�p1\@�;5'5y��x����9zv��i$y�.��(�#�ˎb�W&O&/�=ۍ���媮Í����y.�C�l�'Z�ڣXOל��OCD��f�|��L�l���q=7�G�f��Ln�_+�3o��/���3�^Cy���;"��W�U��}iW/��s�����/��H���^����!��{�hO���c4�A^�W��pQ�h��FAס1��+�m������u���x�) j��\&zk���t�e�9>�*��=yIit��r��Eg�t�ɎE^�Bf�>���&�;����r1e��1<+���c����=ԅ��"9o�tsQ@LR�b*�"�W�OF�r��_�#\��&4+������|4B���Ni��TW� B��z�����(���Sj�0�s�{���� 8���/�]D+��F�$�#I��s��y,C��l�(_�
�-J�'P}Q�qF��Qi���qn�����1wi�x��jƣ�Ὦ*r5���Y��<�Q7uA�s|�+��1��v�bc�]"bh�x@\b�#���m�6%M��t x�F�/�����CJ^��n芇�h�;�$as�S�Y��^��A��S�x���t�k��W9J�eYp_P֦,��9�Mxm�+��5�<E��>g�u�4(ڸ�FȢO�� ��#�2JEV����YF�&�o�t*u��hԱ����\����(�_v��f���B�_Y�u˫�t˶B�:�
ݙS+�lA�tЊ�����\�`ce Avi�-�v����^T/dV��f.H��Ck�lxLp �-}�:`�E�M�sb�"[���c�̇qI�{���@zKU_?��H���J܃,F��A��ߺ3�.�d��=oܲz
�����J��ϯ��F+�j���}�N� u��/1;j����k��-C\�.�pP���@�L 2;��1�璴U�[�Ι�L']�L��lE��M�ܤ_^j��u�^L���'��cᣊ��q(�S�1-� _:���;[&�U���V��fٛXY�R>�����U<�H��Wm�?Z�L�[/��ԏuP�j.}�.w��碟�ɣU{1��Dtܤ�YĆ��I�I����#+�Эoz��՗*���o�F�A���r��}��m�O%7�*��]��|Ge����?�a�L6o��V@,,)��q�cC�o�e�j����!�k��D�--U�hF ��N��YU!��cϞ#-�����^��U�����j]0��S��lgл~<�Z���p�@�q]Dc�ȳ̭�]dD·Z(_�ڿ�	�;��0G���9��,|6�\\\F	O%"�q�̩kȌGwS�'\���D*�y�N�ϧV���h�(��Y�Y��iG�n�RJa�N�dQĘ���x��d_m�!�M�r�	�؇Wxz�j��n�u�ŝ����U�g���T��Ƿ�V�;@	��'���2-;hM0�7b�]��ʽ��p"�f��5mU�Ȓ@5C0�� ����b�n���-�2h�Y��CW�u�uM{��
�蕇���ս�xHi���J�5��ٮ�au\;�8�f��Ό;߰�;t"X�����˒�`��G^�ܫl�j�q;��쵅�s{-5������4��Vǣ�v��s�����;S��Y�M$�_�o`9O��5���+uzM6]%y(:*	(��S����cdm���a�j]Ν��6�ٻhͼ��8�屍��+T��в;HT����}��
�s^+X��/�6'`�1p<��u��
���,kǆ�1�w�e���M!4��\U�8�l��p��V#91il9]���2=:�Յ�Z��Aͺ�A���=8$�P�������w7�eb�l5{�{Iќ���NY1+x�u��+����.�li���V��|����y���ݲ�s,ryI8��B�>�*A�Y�oK�ۃ!���udDa"��xa�5�M�t��4e(��ϻ�t����Eu�ک-7�ջ�]*Z�7`���g�������<TFS?+���u�����/Չ���7�[hާh3+����	�y���7*뵀X]H�]�4�4��|:Z�����pٱQ�1V`�H��Wғ��Rפ^���`�!�Pj�1'z�z�vv��؃TՍrM�]�'�e�gF^:cx��Y�Y��� �or�+iN���4�4N�cVL��U� �.QMt�^�N�`C���h���+Sj�"��}Y�e�Vufl���6�fg�|.��Jҷq���d�k��b+��n�k�뮫��o�[�M=�X��]���\�K�gb�+^�ݠhn��%K4^LM��[pC�;mʬg��Ot������K�ѱ�M�S,�U�z��xթ�T���U��,!I2M>+����ͺۮ�v�O��^t(��v�]y�V4�� ���b�+]'Vfbs.ttB7�.�צ̧�s� Ӏ��{rݰ����_b�O&��L%��,�C)fP0wKWgU��y5�Mx��:�����2�"#,�Y��B�{��|0J�bLIB3�q��ŕ�Fs���;�=ݶ��S�R�mX.��t���B; ˕��^�k��^
諯��(A�skO*V���ݬ�q�黼��κ%W>�P�A�$��BD(�oNЮ��(Q��N9~�S�$�ι)�z��S�zJ�e^��b)�����S��V�M�Z̪j���[���t�:Ob�0�|��J��fu�}]����Z�jf�)G�u�wb���fWL����N�M3v�h�M�޺�:d��xcFMgRwZ�T]�U�?tgR�}-�NC���� �݋�e<�.�^�x��`P�W�X�D[X��&dƍ�b$�RQQFM0К261���b�a�PD�h��Ff#Q�Ж5�&�	��,�L1!�"�F4F+(�Hу%�*dd�u�f��1Y�lh�R۬TQADF#b��$��m�b��1b��$�4�+DZ#$�0[�6D(���i4bѠ�Ԙ,˛r62c��FƱ6��`ؤ�Ԙ�sr�	�,mA����\�b4E��+����cc�p�^w�N�ܡ\�}�1 �Α�j]�ǣ3�Nxu�yg�*/��4���nŞkf�s8�N�/9�de����fwQ�!Wd��[��{�_Ҽ+����^~z���oKA��d����oU�W�ƮW��}�믦�k�x�r�o�����^+�η�����_~�|����k�_W��>��[�z\������/�1}�o�5F_��Ɏ�#�h:�9��W����[�y�-��o������Ư��ۛ��ϯZ����ok�^.W��[�}^t�{^׏_]_�z}5s}y������ߋŹ\���W��2hG� ���zl�!?�y�2F�c֧j�6��K�p%�Dl��ݵ�ᡷ�;�z[�\�-��|��o�ssn�p��a�!�~E�'�"��{\�m����Ž��v��u��@D�"+��h�F����G`�Jb�3��߿���^5��o���|�~z����߯�=�@���O��	�y�.�Ot���x����~_�<��}6�����<��o��^+��u�r���z�w����f�"�4���p\;��Gwj��K�<������}���+��m�zs�oo���-��Oƾ+�����ͽ+���W������^-�~���u�}������^�%�?����m���~����}7��^5�4>���D�b#�D����r��x��xfѭ��/�;���q�D������~v��nU�}W߯+���^�x���ڹ_�w���~��K{W>6���"�;�1��iv��჻P�6��_���ϟ?~��j-�~w��_~����8��GB�1Ț�)��p�G�#�~��x׶�^+���|W�x���z�򾖂���zW��W�G������|��W����z[�\�zW��ט��s\�~�y��[�|��O?�o�"$M��mL�2�wO����DD6�~~}z��ۖ����������5�~��A4=;
D�y�kÆ�@��{[��������h7��W����o�s�_������گk�sr1n�O�m������{�z/���X�$Dx��_>z����w�[�����h�~���y_�x��r������9�s__���K�ߏ�^u���϶������^��1{qVXNN;��P���N��
���~�h[�IFUX/������wvÆ��o/�~j��j�~�߿=_���x����������W�~o�<�Z
�k������+�h�W����ָoչ���x����m��-�^���yܼm�8�� ǮG��k�Tea�}N�6��x ��h�V�1�ݵ�g����I�]`�7<2\���]ٮ�㵀h��BI� ֌��PU`�;wxގM�݅"g�gX�KK���'u��	f�ܧ\`�^��ʻ][��u�u��x���ȴ��Q-��f��s���lG�/;򿗞u^��KG��/��K����?{|W��ߟZ����}��x���zW�|^/�W���<�o�~���{�������o���+��������Q��ɡð�����XW��������/����}v���U��-�����+�p͎��P��v�&�;6�f���_������{��k�_��ο[o��?�>-�wSR�|���e���}b"D} z<~��o�r�wX���x�����������ޯ�^o���>5�_�W���{�}{���_kG���߯~���_�W�ߕ���o�o���W��1^��o�{�������0�����\�mp�Z�B����n>�o?���o��ſ��žy���[��}o\Z=�r�z������k����o���[����4^LxDp��@�Q��4��8��5�W6�	wv�]����	��_c���ዀ\p�{�!��o8ڛU����~Z�^���������μo�ܹ^���_��_{�����h�E�b(|�ЄH�<>�6+tC�}��'Edg��F5��Y>b>�>���#p�{W���W￯[�}����~5�7���~|��o�r���}����oJ������\������ƹ�{��~/O�]�x����}��#zm�~{�!r��|�1��g�^�,D[?}��Dz�-����~7���j���|x�?|�/��h�J�:�x���^5W�^zU��o�r���Ϳ����~�z�گK���SK�<�t��6�k�8[���; lBi�>���B�b�x��^-�[����6���mϿ;^��6�x�w��l[ڹ�׿}|_Om\߫LK�W�N;�F���CyӲp-�!U@P���?�W�T�5Wn�=waR��,���#�p1�p!�]�8����_������k�}}�����^-=}y�_�}�no��׵�_���	`�78�� ���np�wDx}����"G�>�#��x1B>��Ӓ����#7z�)��@p�� ��z]�\�z��y�k����\����_��k�x�^���_��~}y_��^-��k�zW�����;^=��>7�}{���U�rߪ�{�}����ϼ��F���Wz�hݼ�3��y�E�q�[+���H%ƽ�c(����OT��YG�}`f���/-�>�� �;�6D�Z�1�z�{;zFi:�2�.��Z�z]w��wn\-��'d`��0���l^��a9u�0iJt^��'����q\���|�_Ms\���ϟ����*���]���ە����z��o���^-�]��~.x�j�5���ߝ_��}-����~������o��������]�>~zyU�GlV��mS��Bx�_�<��}����ϝzoM�����x��tZ��~����o�}��{���_J�[�����6�s}��z��������ǝڋ{W>��������\����Cr���ՙ	^�.�41����_/��6����z_{��ʽI^��<���h��ϝ�+�{W��׋Ϟ���xߪ�|����~�Š������_Kҿ⯽�ן;^+�_�w��.W�����w�=U�gv�T����)��B>�\����W��������M�}w�W�܁��$�5����!����\���o��W����k��ֹ��|�+�^׍}|������Ѿ�������x�@C�&z	�;�S�o���}���}+��z���r���񢯋��_�}z_O��-�\�W�x>*����7�x�5��}���=W���_���~}>6�nmϯ��kھ�v���ߗ��-�o�?}Dj|9B��+yF�y���� ������Kx���E���Ź�o~��k����m��o�׮ޖ����ϧW��{\�_��_M}7���|W���}-����^O}o�x�~}���W�ߟ;{m�{�no�_I��;�Ef���H�>�>#�m�{���_;�y�5�W>�?=m�������߾[ӛz���o��n�����o]�����W��}-��y�+�{W���~���{o�������ygB�՜=�vb���"�����/mx���^-�|��?���W�Ͽ/�_+�n}����_;���W�>��^��ߟ��+�sn��ʾ��J�[���|z_]W��.^����о�� �0����qSKwϔ?�G�#x��_>|��}�r�+��|����Ѿ/}����kڼU�w����7+�~���=Z��Q�}�|��үk�����/ͼ[���nm�ڮs^��AA��s�[��q{'���	L8�#�_�rܿ��܍�|������ݯ�x>���ʽ-����������j�zo������ok��i�|��r��K{����߾yPm����}�^��m�wߗ�<��C�5�����r���/u±\|���K��:^f�c���ڕ�v�w���s���F�1���g��Oд�V��L�ObY}�uŽ|Sk)n�Yj����N�5���0/�iZ	k71�g�"MN�S`��Zz/�$A���ơ�T��l љm�]}��R�5ϛ�oO��`b>��H��� c����\p��q�f� [������#o�o��޷��+����|���~E�7��^;/ڹ}�:����8��(����p��=��t48����<���� �ѽQ�}kG�����^��o��z�^����������x�z�ֹ|Wڼo���ǵ5�ߋ���U�r�5���<�{^�x��s�|��{[�﹨�_ϯ�w�����mzr:����+��AP��'�}�N�W�����������h�6���~�W��7�n���x����k�}޻zsW+ڿW�Wߚ�ܽ-��W�zW��W�~߽��7+�~���<���mr��Y�=|ߪ��.��>���DF#�B=oj�_���[�y��U�s\?[{x��r�\�������n_j�nW߾����܍���b��ݷ���w����w�_k�o^u�W��_��^���}~~�k�5�,̜h�Lr��C��#�f/>_�ޭz~�o���1^��ƾ��/��_mx��{����ۛ����?=|����}��������[�x���ߕ��x��}_�~o;ү�����-�\���po@��75��1+'�����޳���@�[����J���ֿ}y_�n6��^����o���k�{�����o����Է>7�O������Wڽ/�xߟ>z���Z7���{򾗊�W����ׂ���B#D��|6����P����W�^�y��zU��_��Σ�~6�om�}��~-�]�E����^��n�ך��?%~��ϡz��dw�q��V*h�̤�\q�{��sZf�U���kE�U�^�#��b�!�F�NHo'�	�Lm�q3��墁О����]͋�0�}g�m�����3�� /�_��o\�k^vr�}V� z��i��zh�sZ,{,/�'ԸY�)�w�|�
^�2v�=��jԄNp�������nVM����w�Ů��Z���,�R���R񤳪�tx���j�"�e�]��c��o��ey�J�am<��H���x�^�<���w��4}��M�ҙ��*M�d*�[��w��U��הQ|%+N�y2�W�U�Xmm�8vr��1~n]�;��h�s�4{b:sk�Aĸ���nV�1 �gws��'T[ٖc���L��ά<��Ӕ�Gb��
F��j��FH�ut i��<����7��:���% M>rn2x1��C���pd�Oq�^��I�ڥ�l��1����[f�&�]���u C����Wt莅n�P�m_���=�dۥXE��ABQ���\ �S����Ȫ�09ʳ��w���ʎ6���r&��:��|�52�amu F7$hb��dm3��-��4�N��]F��7oqP�8�������
�7+�5��a3��v�� �OF@uʸ�.�ᢅ���9���,.�P�s9U��Zu����Ԙ���b���.ND��:�o�P�:̮�wC�����!�	��~��d�X~ǒ�oCmJ��ێT�U*�~����hic�v�X���OAݽ�G7<ʴ{O��i��ϭՏ:���5�C�l��Y,C!LlCj��ݣ�|�%��eeyr��V����#tq��W��Yj����y�������̅� S�z�+l
ݝ��h�b���Cf�����:�w�qhn(t�u�o%A��1���|���2JE��]�R�ĆnȏM�Xhcpn�/xμfS��R\�IbΗz9Z�~�꯫ﱻi�X��*����c@��ٔ����c����+ɇ��΃70��L1��+���m<碵�Ն�Ip���b�熾�M�N٬-�-]����uGx�l����{�!zsz7�v��q���=C]�'x�{8����هC6ӦɃD"vπC��������ֶ7�2񢣞��n���U�s�Q��&�ь�k��E?^�sグ/j6lJ\�u����H�k�oj��.�g\�Ϊ����총�n#6W���U���<of��:�t�Ѱ���e���.�@�1D�s�[u�d�n�g���h�C��T踔�EfM��S�Ɣ�8���ɨxq�rK]����Dk�m��O�E���X�B��u;���Wg=�_f�^Szkً�J�&��0r���s@Dk���q89��'G�.&�le��N$��+2n]������
��0,�-|]4J�s��/#�Mþ��3tϹO]pC��Ѓ�H>�R��'$G#q�pW��\��ꠅ`�݈�����2KT���J�j��w�}l��N��uɏ�\Ɍ,���<�p1mwd�[)S�tt��e������,k�[u��oPhp�2�oun�u�S�*�R�a�^�J���b��+�r��Yۙe��r�إ��gEq���݃��nK����`�03Πv�9�Ԩ��1�0�i̍��Ī+��l�9Ud��HJ�M+R���.
w'������XN&&;.t���C g���Xjt�d:�nc"	���˘���l8��	W]Y��xn���ȃ�l�k��M'�����̺��8m�B�.�9��A��=��������U3�j�>J����I{N�v��?d��]YB��cB�R�w��Uܒ��( D`&��ePc��l��9<b��7,a��i7�Ɠ�A[V�0w�p���4��#�q�Q�[��a|�K<vb8o�ܒ�c��3ƴGT��)�;�u���q�ؔ!U�>�ӡ��=�1�NGP�Y�I���p՝J(�$S�Y\�T;�-EhT��d�t4���Le��B:��B����j�k�b2��C���*��}|���ݜ�a�B��̱��q�]R:+v*�N�-�q�W�X�]L@mS�
�cQ���^JM��s���u��z�r2����ª\%쑼i��:�MoF+��7Q����ќ�̠ӕ.���r��T�2�G
�AT��[9!�"[��>�u31@��8��'~�1OKN�VqA��!B3v��k	��5���H��P9�9mñ��8IWH@vƧ�r���ٯUo&TC)�o`e�"��wZ�w�P+wj�-�LIB���m8-p|�Z�[W����p�N�ޅu�
�o�p� ��D��?Eκ�#�JZ%��9LNZAs�zsbQk�}P5������mף��+����s`V?� ��Vye��C5R���|�ŌQ�s���[t�#�ă��r}p��]6ph�7M�"��o$gݳH�B�m�x&2�w`�6$�䢥O`�V]
;(@��a�I�q�IS��c�����L;�9F�C���ʹs�_k�*�O`�<`����_���*a����
���9�G�y:y5�1&���Wh�.����*|����� @�@J�B{~�@�EN���އ��:s�ư�6'��\����cAv� ��y�E�0�_Į;R@vS�R��񙆼3�ʵ����{[xj�3\ٚ��Eh�����.�����5��!��
׆�+������bGu�o5�.y�ԡ.��\�U"��]��Ð�P�9G��I��;�L�;�^tu��Z�6�V"���C��lS���&
25�w����}#v�f@�8Ҋ"����s��1c�u�x܃�������:]�|��6��`�3t�Ev%�")�Ѯ��{�+6�8���)���%s�v���O[�v��u�h��)�dr�=�0g-�)*mu��� �j��v�3lpYT7�+��o��#\����/��  aaef\w<�P��}8�E��80;8$F}�X3Y�
��yd)ڄ"�S����Z�Dª{7��V��+Ss�	���{��H֋j�puP�	��)DnR�NH]�w��a�8���"�u~]�����{T�Vj+���+Y_X�ɅV�l���U6�9c۝Ĝ-�f�Q��<7�Y��Z"bH������قY�~���n���_;�ˡɈ��\J�0T�^����]�9��]�3�^�Ge#�(\< �/v �,�V��=t|�[�7�Nw*5��3h�ʝuaa(�7�Բ�֦���c*5TVi�����z��gWi ,>�r��� ���FZ�[rN�k��pd�n_�V�.��u|�g5J�F�Ī5$늦��|%	9�n�v���oOc;�Y�E�wG�2���i�E�ɝ�̀��p�}K�s�9�2v�0N�성��-�D���Qߵ��Wr�L�`�Ov>{�.�p�+��}H����FCR�G8�C1����(��^E�]?Z�B����z��%D�D�1��b����\!`����@� ]��n��J�óV�C��V/j�i��)`Te3�F��k1,Vt�EҔ�//���G�G��;��*�����t<�_d�z�&�4gZ�Ӡ�w��R$�4լj�f��s��30`��t����L���BM��ș��A}Z7X ��tE#!OI%�`�ٴ嫚�݉��I֏�S���wN�����6���J���$�ɂ8���7�l��jT�� ��;�%[�Ӱ_QE��q�l1�d4Lf%L��<'����vY�ȇ��T�?<�o`o �I��X*[��-�
�'B�(=�VK�S�W*���l�����o�#xI���n�!��b=�/�̆�j�{�<��B Bx�9u�W@��fnu$��
!�#���%�7@�/:�e}��F�q]_�����^ugd>�QF{rI{�ȭEKu�	JY)cOG;�����"���l����|�p�~�Cj���#�qw|� T�8[N����c7����Nx�N��_t�?iXB�ԅ�"^�Ȭ
s2t4$t�EgF�QJtB����D^���O�H�]-{��̜ôzH�)��e�M�ie*�0�L��׳�j��d+����%�]E^�+�+����Z鎕e{���/a���M��c��(zL����Tw��W�!q�J�|O13V�b�$o�A�A�o��RMCd���n�m�۬|�7˦K( h��������O��P-ӁeIe�JY��'��aU�[��gwb�f�+~�����@8�9�n�\n�6�eچ��xj5���f�ѻ��y��`ۦw5޻�-Z�]��dTIT�b��#W�:Y�n����&�ޜ�%N�q�!Js�I��Vvx��KU�f�wm08C'�HÖ����LW��[x�/�oT�g)���C�LQ�>�ֹ������*�B8E��	�Hp�4�Y�kM5����7���=�u)���b:���S=S>Z8NqaB��AH*:B�3Q8�-vl*�� ��e��i����W�m��_�=P�^�e��Eќ���yw\�_S�2��N�L,�m��b�-�\����l��
Q��s��;���o;qtg*t���G���-�%2e�]$U�uv�Lf���b�,֍��_��:,#��iC��Q��qQ�WY˜�/���T�v���'{32�s��N�ݳ���j�c��A�ն��:ƎL��T�e.��|Mo36�+���ٽ�[�4�T��vn��l�N��PJ�yA����`�[�]\�w=�H/�TUwtFn�5s^=g,���KK޼u�>t/�"���b\�ѣ#J8��<���c���b_GL]���ɯ�=2��/��L�"�ȥ�"�)i�s)�W�&�O�M�h\8�H�`��;Y�Ѯn�S�<�ćN�G� ��j�:p��5_��ʖ
�e�#|��ꔸ���4���M͔��qa37Ep\Ϊ+t�gܑo{&(�<��x�Z��0N��6k��N��<�/���3������t�4�9A�o4ջ���l����]��nW�E7 JsU�
R\�K��CB�>۹��F�� 7m���:�V��� ��/eqie�GI=�R֎CM^��wPC6m��{Q]o�3�x�
|Ӛ��wX౲��v[8�-}M;\����e.��t*�a�v�d�3�2v1�eō���Lhil��_.�p�ʱ\�Дn^[� "
�:\㕜}X����F �_˭�o�8j"�o0��=��3�����3�E��)����c�ۚ�^՝L.U띇\ҁJ��Xw �uKP��,X���,����h�ñ�������]�J��h6-��h��1��kL��qƒE����C�=�n�r�>���>��-9�ZȞB�=�
$l��⣇śi�v���a*Ky�m�Y�9P׏�Ƹ�+?���/�2���r��+p��H��}�FQ���q�u��UȀ|;+yGy`�v��Gp�u�X�C>�5Z�J�l)���j�v����w����b�z�ά��t[
z�s��X�U:����D�5$�]��LO7�> �X���(dQsnI(�b(���n�ֹr1���A�h���5!cQ�ƍ�wWJ��"�����F��1EEn[�`�\�Qh��ƍD��4�	�QA�L�*�\-��4I�b�n\�
�����ŮQ��4��s��[�O;W6�ŮF�,A�\�",0,��]�6��-��r���IW(6���(��b�ܢ�I}g���֍��wmc;F�@*&�.=��Z��c��;�[y��d�_1J��H*�oV6�����m��˟30`���TV����N�t�~͹:ZE1��a�A-wF��2�t��cp衵�{w�54Q�wD�0�XA��ii�	������Ud�9�MVy���~]� ?!<9������ڏ����0/����e�!qD������P��1W���ܝ�q�K���j�se7�}��J4�4WoTr6;��	S��d��b���Z��� ޴7>N>��Fr�3��!71"~��ً�C��;i3p����:S7f4G��iV�.D��"Ox� ��fh]�}�<��Ep�|�G;�#"��,��1{�m�����0��gd����F�)�{=A�+((�fP�N���ىMjc����^��2��B�`I�C��9�y��rެ��;�wK�$ŀ�����5�ϒ���(�[�?9刻<+�w��V��2�zR�;ͩ�!��l0D1��@n�
{�$d@� nO��Cr�3���u���2ip���ڽ�����Z\3 �eG3|�-��K:TLF�+��s��W���Y\�?b_�!��Z�Ti��>�=�Z=�������*��Q0jP�n�jc���\ \f{�����,���6VcH_��Ѷ�=����<;N�+�ʋ�oi�a4�����>z/��.1��^�M#��Flb�Oҭ䛍�� ���+����0���6��p��?S������p�)��Q,@�{�����2�J�fx��ՙ�Χ��4��A�f։um���
�q�j��sT�:��1�#��t���QE�+틟OV�u��������!�+�k
�0�i�@՜���i����X.�Z`[���xkz���֎�Om�ʊ1_Z�"(F��&jQB��q��,u}��/ৠ�.j�n�
L'��q�n���c�U��/ް�m�bSG�r+ꔳλ�o��v��u�]��8�ӯ�p��-�����p�y�t�T�d�Y4#n�<��\�����v��Z��l{*8EE���LP<k����"鳃D!�n1�
u��</�[<z��z��ѝoP��=����V�@^Jy/
���5>[$r<4N�O1��Rg#O�*_@�軭���p�T,'�A�ܴmG�����*a��[L+�Ư��j<�e�{�c���eA�H�r�E"�a���Q����bw�a�5�*���Cft�˕���}��g\�)�L�טp:���eB6B`��@��x u��SH����1��.�ȨFi�\�`�A<�:�Ѓ�O��o[w�N!ux��U�Zd�WW94V7�㚢]ث�X�;����v�^SD�`���J��H�93QK�`���nv���;��ã���1�P)D:�[Y:yV���|���J�kB�]�h�C��C���NO�7\	�)�L[}V�9tu�0��"�:� C`��tD�F�>V�0#an�.�C0�"�����t��@U������i��MV]�A�<�BAܞɇ�Y�N�loA�(`ڼ���Fl��g���8�T��"p�]�ّ�s#�!Q(푲��䕜�SE�� vH|cK�1�U\��X3_eB���ζ�9i:�b�WI��l*6q�*�5�8c�0w�kE�n�:��xAaYu|��?��S�.�E9豴+{x���,��u�5A��eϐ_Yv:�q��o�pB�u�M�bW)����X��� ,F�e���M��wr9���т���Dtܤ�Y���}���4�M\��N�ء��s�pUt�^���:��v��+�GOi �ܱuTwAj4A'��p�Bq���&-��y2�1p�a3D�	eaL�t(�5�C�S�W*,�L�q�4"^�� ��Fn�է��U+�`���mp+8�9M�d��)ȫx붷��h\%Z[YKx�!r���yA�8�Ya�m����7�-_=���c�P�� � �}�Y�x��'�P��\���g�M/�˭�g��z�rFvX����u#iY���0�4+~̷��s�h:=�� ��k�.|�o����n�I!�����|l\@H9�4�O`�ś����tZ�v��p{~���t��;F�@f��l�ᤸwܲ뵑K��!�����ِ�s��R�>q�'��A@�N�CӬ��>H���Jg��t��R�Kx"��V��}� 
�⮽��ʝ$Z(�����	�Q��P����ێ"��>�y����z︡v��p�|�iTO:�L����7z ��wDT#!OI��8C`���*��m�1��c��NKØGt�!a�����P����5&��:�yd����暜������
�H�[�+b��a�{�����`H�݄��(!i]u�}�����u$��K���I�b�
B�SLs��{$!g_�f�'�H|��*;gwC��Zg�b�B�6��5����s�hA�71i�MImP:��nQ^~Kt�)v�|;b� ^0z���4ǝ���C��u�_A�$���C�+�~����X�yĂG�=X�6�N�`��J���t���D<	C`J��v8J㽊Y�5���s~���7t�P��0Ka�Mu�J�f��I��-#�����Z���W ��H仯 Am*5��k8���/cب�1��j��6�S-,��8�nU5Z��U_U}����s�(���ӳfհ�e�M� ��j��#�u�� !L擩	�����̌v�S�FF�UeuK���f�],mƧl����������Zkخ��NK�.��v����f�c��®#&u�R��e��iK�-�¬�qR�
���t���[���߽�l�*
�.�(F��U��i�}[u�dD�Eq�Z?9��UĺI���|��'n�NS�bk�1�����c�ϏN}T���Y;a����kuQ*^��V5f*�*֞:eЕ�/
��w��S�S:LF���)WCp<��s�BN��hp�s���%�ۇ���Bމcw]��;�b�:r�+>%5����]jn:�w��{|Yaw�f�W��
*�O�)u�s���n18�J�[uPB������qֻ{Z�k$k��0xu}s'�ҸňC���u�sS4&y���m�҄.e}��U�es�z�f҉r����e#Z-�J�o8���W��|��J�\-�N��uJ���:����l�_�s1�5�A�;R,7��a%j�Ҋ3*-�Ö;��}��X��\�O_������ԃ+�4�6�r�)m�ֳyS�q��Kճ[`�o���yY�vVn��g'I���V�lR����3f��դ����{n�r��*3��U>T��=P#^&#�F@�l�)��A�H�7�?�V�] e�|0��R�;�W��)%�p�|�UѸ}!���%߇@wi�V9'�մJ�Ԯ�)�xS�XH���.��N��y����]q��E�b�@�CST삶�1��&��'^�LK�tf#��B^�Vo=M�u��8E�0�7����s�3�\�h�n���p��L!����Pe��Y��/R���b$F
v�ó����6d��wtV�'��<��1�f��-�Wr���=�q���0j�-�&,1�E�o��LV���ٔw:�ʮ>q�!����b��l��*�c���^��_2�!K8���
�!aw�)��׶*�N�	��^|@����r�3�u	8f�0�\��P� �;������_ƶ�1y�R7&,F��&hu*.gr�O�G��|�ߓR�؍���q�a��t������7'G^ȝMȯ��sT�V�V��Ov-Hx�<�8�\��4#{e�=��2:�4���~'9�������D���.��yDR������T�������z�n*TN[���\���΍�F��-�����/3zf�ȝwv�wC�Lҡ�Z��r�U���4�aW9W-6�#GmǙ+�%K�[�$ح�]����2�����!�32ڃ�[���P�|­�;�Z��;�ǂ4�
�!9�b��Q����l�;0���xR�����j�#���B��]�M4r ��s��t*
� W�(4b����$�#�T��S�{;Jq��m�'�9���rP�0R=s򘊞E�r�\j�B�SOd�x��=H��R�k�t�ܮ�o��C�� 6�ٮ��$d��7-r���Fߨ��Oo���̫���f/�.������a�ҫń7X?��A��5��=��$aOH�U�zs�e�I��U�i�7n3��L�[9���R: L]���L1�Թ�簵G�C��}�+�9ڭ�Q^�E#9"�ڝ�6��9���F�%F�|05�\e0���'V�[����4k���}s��FJf{�������O��:~�bBq5�;�|�T���Xm�3M���4!��Rf+���O�u�LGu�����Mt��Ef��s9�\+��!�ײ�w�,5+|�֋j�!V^�#��b�!��t]h��]�&7�P�ӥG��r+n��(�]B�GS\7wVi�^L����{�6��oR�K2�]G�����w�i��	�wY��z}��T������d��n�:V n�h7K�`���Vq����ԧ�@|rެ��h ��Wٚ5��R!M�6�ôP5-8��¤��vEؼ f`�U�8u�)�w�Y��=uj��my��-��W�����}����8!f���O�p��3�a<#^�/�@��Q���%�1�܎w�+殥�U����~&�Z���VxV���M!;���T)����f1��C�!I�ԝ�9�[��w�q�E�=�<{u\��Rs�*{,�j�܁��N��Z�vJ0�K�7�h0VS<�q�cD��]�����..�<�����1�z�I�u�%�*k7��Z8WZH{w��-{w�Z���uЎ_m��zDrOVFᑪ'�b#\V��^��\GA�F�����\wq�5���UX��ՎoU�U�É�W��:�Y`a�J��8�|�|�BYU�`s�e��[���s�B��`�k�
��$)s�z�@�d�#!�f�@�(1	\�X���I[�U�iV�
�xr	H�����W��>�L�s��t�1N芪↮E���Q��v�vKyޑ!�!�C(���N�̀[;� ��LW���grJ����ù��\ʆ�U�Z��<��ʗ �-�#1Wg`��,�6XD��s��cHط���!I� �=���ʎ�kκ0�LV�H;���*ڛx�u\���}]���ɵ����}C���+gV;\��i�Y�[�9<����p�@�⏅:��G3[g�R���<-�d�m>�ಬ�i:iߩ�s��Y~��XM�s�։03c��F=�HnH�(*��cd�C�(7��l�7���r&�#f*T$�CY_;F�A�Oa!qÓ���
�a�B�����i'|��\h�J"i)=�GT>����������0�ȝ����d�� ^�յ���n|�L`���vn3m F��FY7��q�0�6ӡ���8T`xI��ם<I�\��׍,�L Oa��zyq;�W�nM��Ӓ&'��^2u;�]�뱂�z�"=d逋�|9�����ʢ�c�O�y�r��<�6W���7��=���ȋ��c��v3�
��K^PK���Ã�mw��Z8����}��M�Ɲr�a��T��ں-������B��-�@�x��@O�;œq�M+�M�FMN�Y�W8D��'
z�c>�0^8���*���	�ck�RMA1�~A=w�|�th��=jъ��lK�zwϞ�1\~���������ǜ��m`��_g\��+�dЊPF���K��FX]��u�!��#�:���foNC\�`b�L���v�_��I{�]���n<�cE���Ȼ����sɆv<)U��@Gc��9v��NC�������k=n�f6��O��[��|�E��w����/N�o;����J+��6�ka"�����T�H0h�Z<���{��
4/�~�.��d��W��pW��\�������tNN�r�;o#.x��_9��L�\Ā��!�}��xR1N'i3p�cDp��q�0�OU�M�����ҹ��a�R\��Mc�ariXL-��O �e#פ۽:��3�$�ŉ=���;&3U@�M=�A�w$�#��G��Q���M/�k���̝:/�Õ4q�5u�&�:uA������V&���Dp�>l�s/�ϔu�k,�պ٫�=��A+���fr�=%��l�.�4r�,t#"MHx��~zd�xa�D��:�(�����Nta���<��hd���da�¤7�Y��D'TYG%�73������U��o0���_�0���a"���O���İ7�Ȋ�X�GSn���rx�����YK��Jb�g��S�q�j��xh�k��LV������3˫�:��p�_���΋p+��(X�T��2�s��{��>Ŕ�7C.����5C��9DcG�����
�.��9\��0%|�0L��ia�����D}���b��س&g0n��z���w�$/��+GXKl��9W�v�hG+m�
:�n�܅�,w����l�$#����G�W��X�v�+3BXۼ*bR�.�Lm����ɥk3.�7��N����/�G��\5�Нln�*�h�(S�N��Z����f���gm�U��#Fv�����^t��i
䚢'���C{�����r��	zl9X���Y�J�p��"�T��QKB��^��f+��7ip<y��V�l'&KX�wi&�=DL�d�����Ā�6<��e��n�u/�}�p<f:�'xľ="WJV�WN*��a40\����+�)P���ǮC��{x�9���h�Yχ�zVA���"�{���/��W0A�R�S)�!�%�*��#z�9��a{�o:�lR��P̵�a�+:�<�����DsGh�}s+o]dQ-�&���)�jխvN�JK�2g7ZLӗp�G]n�C;2ښk��=��z�i����ou�u��,:�/3N�u��v:�ͨv�&ҭ VV#�cEr�VǶ��+�5V'���yg�7ʳj��O3ݛ��s��r�z����N��{{���y��s'^�ذ�[d�Ѝ���D�v�|�"� 4&F�	gQ؛2��	v�Cz�-W�c7��o`�J潕��n*)+�V�ݥ��C���z�9t��G�]�˸[���]�Vl�@����f��$�2f�4y�*��q�)�ہ�(��6w�+T&m!W��Mt�nʉ���6���2�_S��w; 6��f�bCl������vC\o���(����]P��똨�lK@
<��:�� -�g��0�V�!@�q �;/��p�oO�72��9�R��j'�ՆΌx{i�7�3K����:p���A��xNcݡ��}sx��G�	Fٵ�g-��J]�G�����Ĺ����J�ήV�l��8����S�Mpt�i�6���f�\�v:�V��]1e��ݦ_K�{�Rc2��C�V/�"U��;϶���ee
�_aX��R!�h�tV�p��Ѻ��|e��$�ja��ס�V��r��X;M	ݕ�ҷ�Bԫqv���s)�Z��t̔�Q=���	�pw����Q����ߤ���WU����]�A^P��H��T9ҋ�ś,�a��:�7���m�Y�Lom���|B�4�{O"���Ն�='���x�C:Y����yP��� I�����΋5U�؞���pδ�᤯C�w��QRC=V�^�˦�ѭ9���G�yv���{&��x�v�i���UՓo����c�Y//�뉀y�]�R��hw kS�<��	��ؙ��o����|*��m����p�͹��ذTPTE�F�,[sZ�K���sm�F-E��k���]75�
,j5�`k��V�ۅ�Qm%ͫ���I]�nb��nʌTPnk��Q��F�뻶傌�۔X���lnnk��&�����˖9���kf���(���_���y�GS6�����ﹰ�蕮�!}�A4E�}��0�^tk9K��.�mS)�{o�4��9����LzJ��30fiŷsDuv(�G\�٪��n�mT�6/= ]��
��\"���үV�]�����P��w��R�^I�+�Ӧ 
�RمG�7u�W�m�b��H�+.���g�?^]�c����k+ɺ~���v���W�R4�Ǡ_F�Q�s�t�Z���7bxo}�3Ą����tbwWtrz���w�t�\Ʉ�DJj����#\�c�*Xb�^�S��W����^lHy���u�Ӂ̳`l�\j�S:��ׅ8w�J�T��\�\<�]6ph�7N2�K�xc����įw�|�M����@�\@f��(@̔0�N��<4M%o1Vg&��a��˘��so���+K��Mǜjn2�� A�9"6�(�P'8�*a�[,"��a�o�M�l�<����p��oú������H�KcIpՀ�V���Ҧpz��i�U�s]*{-Ţ�Q��3xΎp��(_Ϧ�Tr�����e����<HKXNT��������]ӭd���Oiѽ1�w���Ɋ�m�[,�7�����B_��n�%�*�WU�A�]Zf}��Lxw�L.hw�n� ��Y"es�\��4'��\���1�N1�V�<9��V���!�.��<�*�1��c��c�Qu��@��j�j;���.df7�,7�bmrאҚ�"�ʂ�-*�(�U2�%ZP���2���[��%ЮN��uE�W�}��ؘ+�:Y��W������Z��Q��tm)�����N͛���Y�fWm��+3�����Y�@r�κb$1�y_*�����4��D'��_9��s^�▬��GK�q��TQ�!�$�;� j5�AGd�É��c2��Ɯu�:�H��ԯV��-T�u]�j��G��8����-WӕW�e�B�`�*\m��I���]p�N�s���S��䋆���q�U�^�����V~��k!�_n�nz䮎�L)��ЁB9��vn'g��\��:d�C��=�'���~��:m�$���hġ���~��a����
�BH�*&9�MA�EH���4ݐ8-�_n�e�N�/�ur�1Y���[W�4$@!�Oo滛z��L�Zل��O'x' ���r�H���+E��xN�<F)]�_�S�5�e.- �� W���o����o[hzW���R�/J�l+pm2�E9Y'^�"Q�0���V���a�I@Ιr@�J�̭!>ot��͎	m	���i��n�us�Dh&q��(�s�E�Bz����H)����\h�\39jg.�#�j�mA���Qr�1
Ѹ��`�v��}A�+��$��X�B����7���pt�]`��r��Ϋ�z��z̥�������))s�'H�D-��B�[o>��ӹ�`�N�C��u1Q�G �	]WQ�=Z/��\���X�]�ġ���<�	�j^[�N��{(�X��2*�n���ˣ�o�Q�I����U�=^8���h�n�)����#��O-�oδO���"fv�P���jc�\��@��.g_A�������9�����V���ن�grg2h��;�׽ϻ)�;�i�F�@��RI� �07LJ�	�����-U�\o#������陮�r�_���:���g
���0����"���l�F�c��vϭՎ�������;+/����2�#�C[U�9�W%��b���5��B�A�Oa�+�����s�a\���l-f�i-Y\���(�\\.�k�`��Od�Xf!��9�ϓ�	���Ň��ɳ���!��_^��al��f� PεL�Na�o���,e�͋x1S�*WS+�_M����:h>�Z�r�J�k�)T�Tc7�X�N�(`�ws���U닪��/*�ֵ��!�x�� �A;��6(Q;�3#8�� 欩��A���p1��^w�a�����1}]����b����]�>6(ᔢg�u������u	m<���UѪT��'<ɽIw[������"����u�κx`��".�\����U����/T�b�6]}���0HV���t�Pط�C��W{�8G`Ҭ�FiW��(Ⴀ���r��o�Uxp��yo�&�Ꮞy�����@���%yw���Yy�Q������v:�a��Kw\�-?]о�:�|k4��U^ctb䈦!�<J&,r]w�.(_L���:V��ȅ���U{D�&��|���x6o���j�
�+KY:>�*��4�C1ƻE'u\t�Vv�J;���ж �L�oi�bj��a�KW�<}r���]pQ��i*��9H� Wp#Ն��3<��V��v��	��\��j p J��Aw�1"J��.!�n�i3=n�Δ�c�{8��O��y�=#�ޑ���n\���J��Dp�h3�Vlzy=Dc�y9�y��0���=�5�tz��y.fX��Ϥ�9x�q�<Z�./O�R�"W�n��ڨl�l@\;_��pX�*!'V�|Z�ԑ�0��6k���|v�G]��RT�2ߩ�c��!�&�Ц���տu�:�_H7^^��Ȅ�c;����F	��
��;�L6C���Hys�z:V3�:�(�%	��F�����J�_W*�D�k��'*� �dC&v�VӼ�)-������]�%e��m��k�[z\�j_k7N9�kr�>fFP��9K���ouGAMw<!��1��X�8l'��kK�"ƈ �9<`[ڨ9�×T��g ��6�Met�Oz���
��>������;�dvɹ˽,�Go^�[h���(?�lǆ\L��ܘ�V�����"dc#���:L�Q��n,��Fzz�(��<���ݜ�≌�S��^M�,M��#\��,��MĜ�b�&��/qP��ޝ!:�3�})�ᬭ ]�H�l�\"���y32�5�.q=0rtSY}]�k�,s�,@
��-\��o/�c[e�aw�AXҮ��wv���AN�4�b��y3��DV���6aQ���iƦ4cwLu«��[x+�dFȞ��8#4���ȴ�D�vޫ.�+�_A�i�Fqշ27��-/|z���O�e����U�h�WG��k �i�5iMh��� N��oL�DR�b+2y�bFq�O�"�!»�잫�)�}X���#9�,ʤ����B~����;�_|T��XH�
xh��=	��X�`deLO$�Ҹ�% l�_ l�E�pr��)��/M]s;��Uag03�N�3e��u�*��r��*c��bB���r��Ne���.;k���Ȣ���fnU��sfu<1t�ֻVl��
��]�d90>z�r�c�[!y�z��RF�Z��}�юK���N53�Zc��T��s��B�gi�Ct���b(�r��9�PB���W��z�<q���槇�Nu�z�����p�I�[(Ӓ�*�8��ˠ���挴3bJ����.�-�a�)�J�E�8<�`���t�1�1ı;��;�஻c��2��l��|�ȿ�`�����7a��8�!Ɋ�ɪ�7��`���dD�9����M[� �ׁP�J��Dcʃ?!��B؋U�t-.�|�Ɗ�9H��ٳBj�h����oi�=�h���9����Q+Ab0D�7�+�QyLMd��f��&�w��:�/L�0��lw�#"�w�⣢�N{Cݻ^>qk!�d�p�ƣ_�TuLS���īx�[��=�|�� ��28bu�*��i�Dþ�E����F�[�n�8}���*k1���v�q�8u�:6�e�%�#>\�؁����[H��B�;��e��h��N�����PB��8����q��w"�6�q2��s�M]pѐ�E|&x��93�;����'1Y�S�޽��.�3c�����ީ9���e�8�n]��c�utFJY9��kDی�c�Nr�}���ʷ>�K5T8YӺ�HY�Ϻ�3So�ԡ�E��˷/,ֆ�΢�e�դқ�X(v,��~�DG�J��nʴl�m��x2<���e��q����T�1���o��Aڈ�.'�f7�q��5x��%˗�勄b�[�:�~��&/]¼�F��	����Xy�,�9d�!O�u{���D6
w�
F�m;*�K�X��4�s|�:8Wu����Lt�J|^:�eoܴ�G���qa��Y�>�b8F��%Q����q+&�[Zk��gq����qY1�h�|ڿ�	�;��2S���GN�X�#$�JU���o��q]��ҥs�^m�a\�7zU�M)}�	�A�F�ڇ(�r�:�'w9���lA�\�>�8c8���0;U�ٗS��HӝN��o!K&.v�s���3i<ٴ���X��}�a��q+s/��e�J�Ld������J�oe;VW3�jB�/�<�:��I�wQ�������3��qX �{�;��gc{+g�����)5B��"c�=���]ykm��r��J�ch���bl�)�J����g�q'��X��ws�{�Q�����+(d�~�5}�7{/o}ʝ�AOD��g��bY�����s��νbic.�c��j�N�/�����+lޱI���}U�{���T������Ӡ���"�
���xyO��9�
{��(d3<��W��r���̖��F�koK|��\l�wSQ�V��|��BS������kStE��O�z��r�=5�'��-��U�C�<1d�����N�8vٹ.Z����kV��q�-�C6��qM�k�v�V5�/�Zݲ��I�\�q�O�����6��C����m�?��^{Uwh�6�f�A8�K��b����qMl>\���÷#m�Vu
��ڢy��f�]���)�+��p�f��)�����O���S]�p�>��=0^�Q�X,\Dk1��F`o=�;3;7�s�9���Kyx�[x�Wr��P��0kK1/w(}��S�V�:��w#���SJ���q�Γt٧�*�].7�v�"���'069TK���
�\����g3k����'[���?+V���Ռ�.Քzn��J���r�!)��q�hp-�ouvm;�(��6I��f���W�cޫ"��r�ꜳ�i�:p�e� ���=���4�Zz%ʳ��̾�T�4yXt�f�����ёGV��xB�*����"�]ǡ��j9\��9�*�B[F�����]��w�v�P�����@^2�K��wE'y*ۜ|sCp�;�=s҅�]�c��p��*��-p�,�q��T��{���&���{��:��*��^[V�V�`*7��L-�L���/��g���*Ru]T5p� ����sg�A}���Tr	�¶Z��Š!��iŭ3����:�r6���t�!!�竴u\q]����;C�bq;�Ux��h3��(O���z�y/Q��J�J^��kS��Y�����-��~?���Ļ���ʾ��;0�����j.��Ng��p�釥��y�����Z����~x����Z�%ܧ!n���#܅����O�Vu^��\3(�|Ud\�ַ4�/F�S�R�V&^�m�U���V���W�M�m���v;���z,�m������"�(e�v�Q\�=��� a�U[β�}i*ًhͲ�):�^;�#��ko��u��q�P_5��dWq����u��Z:�Ng]���h�:^R�B�����Ģ�<ۅG�7���������GC�KJ�#�}�%P)�5��uʻ'��d򨍕Yx��L=�k��oe^�m�w/9���6M�
���N��{�OO��"�;��=oψ9:��ky��N�F�-�pzNF��TI���-�W�|�G��Yw�'��A�qs�C�b�/T,��B]�����%â-5�G1���h֙��n-��:��l��jW�r���Rߙ�U����%\o�Ϯ��Ӯ�m���Ȟ�؞l@����ۑ����\c�T���)G�.�1��@�5v5���Rs���<��2���ioC��k�u�yWO����xy�	�S�L~�[ww"��:���y��eG&6��o���J917qQtby�У�r�j�p�K�]���^���c9��[Q�e}���܌��%l-��WQ[�-
'�Y]p͑)0��/��.��V�F%b>�}\����X��X�Kt��q��R��X�*�E!��n��t(Y�G"�J��RN��s�/���lr��R�3�hvykz[]��3��)p����$��G+���=�
��yijf�j��濲��\����z^f@�J�M�ó���'u<�Zn�;WY3d�ֆw+W�|�ıu�"�9���OOu�=�i��"�v;¯`�`����wg�VN8����Ә%a��Ew��}VWʕFw1�ٛ9��؂��7����\���P2�L��TŃ�����%YX�GM��juEv�(�����͢��T:��Ļ	a7�_h�Al����ګ`U�6�z���Ir���7�Wp�ƥ�[2�nu%�oY�ܲKe5�ȶ�s��L��/'�i3;��E�J��������Oks�4RT���M��c�
��[J��	�����K��d��R���+r����g��>f��ӂ��Va�ݻ]yhD1�%��a���T�e�:��/�4��}j���G��Ɂ�n<�+:��S���.�(���=�*�}��	�y�o'7��.c��7J��tV�S��t]������顤o��7����"�*1��U�t�J[ݗoh�-'Tu�]
�[�r��^��Ω�243yA���6Nh�33��f㈞x����v�vQ�����v3���ɷ2�p���#y�G���k���I7�r�wE��6��쀈��&��F�}\�z�G�r��3��̹Q̪W˔Π�o�w2w4.2��T�K�i�û�ft���Iu�f��ΊJ��B�=ǟ��s0.���z����].�p:���R���؎2�oR 7�1#ɨ�]�8m�ӕXt�5Χ׺�d[���}�^0�A1iԞw_�]�6���gLo������u�r�{�<��v<�|;zk]�\��ݲ��GTs�v(G�Y�-kD��m��������`Ӄ�
6�X_wNH��u��z�ⅼ�Ӗ���A 'D��1K���e��K�|�=�Z��r�tS�!��ޚPA}�Ej�#��ITF�u$��0*��SF��p�"�/�b�_hn7���Fj����CQ���7F�;W���/���c�
5NӨ�C�[/�HUo'FٶmL�����kVp�+�	��};jK�4͞��G#���dn��4b�L�*	W+\Y�ۂ���l����Y���egR[:�J���+�5�r��u��mM�|���14�ڼ{�җkep��LCN�22���4)��<�^�4�Qq��%�Uy$8#�z�1�H��pΕ%�&��t�w�n5�#W��X���k�˗�FR��a��m6+�Z�,{�J�ڹ��g6�f��2h�mY=���5�4�n�٠�"�i��]�(�B$l��v!��T��1��ig"/�bZb�&aT������L̙�V�i�U�ɨ.Qj���s0�sPZ����X �]��n��������fNt�,$�d�FǴ;qo�*��t����1r���Z�d�cB��N뛜��ۜ�G,�I���wW'u�r�r�*�n]�sQ�W6�p���ڐ�wcX�����.�:��E]�F�r�n\�]�tۗKE��]�k�͓]8k�Nnn;�ʹ�m���˜�k¹]5�sh*w\�I��2�Yˍw]Q����\�eΌZ$�H#й�r6�d
�˛�	�M	1���2�)~z��������;��ׯ��[=�c����w�ybwϻH.�%U	������<kQIq�עk@�+MΆ�Y/Jm=��g������>���GV>Pz�y.�7�ui]�q:��W��*)�U\t����p��(_� �t�Ʃ��>���nÕ���1V����6�PdQL�.�F[��V�{Z�ȏz�����{�i��iwA]W���̬֘����s�Q�Tq�+����˛��y|�W�_kT[�?i�\��p\9\^p�<
��KSԪ�:�n;�ڧ{��sWھF�9JtBYWڌ�9q��ޥ����
�/��ΡZ���5����ӄ�y�ʬwu�6�h�6�Nfs��k���5�z�.����cYQu�z���t��b	�mzo��-� �����qŬ��v�{Ji���m(S##z�\�eHǫ�dT�c�ԍ������L+{5�K!��o�)N��*�r�B��ԣk��{�z�sڝ�H^�J�I�`�W�(����
��?;�0f6�O2Xx�oFNߜ�Kvc���V��l0�v
�&�DɊ��u�]�F����(`l]+�9�n�umS��-���9u2�ގ��<F�4y�p�z��H.z�s���^ʘ]���¼�5�uY��v�v�.ڂ�^7�����D� �)�n9�^�ǵ9�WL-u�f\wJv��z�@O4$��[ˁ�M�!��:9](�6�Pҷ��s�*��F���9ow����š�>��9�B����U��.�4����a�X�V
�\�3��SS��Y���52y���lOCP��}����/�J�W4�V�h�F�r��\_����t�̅����\��l�c�,�j��)}��W�گ�����׏65h5�3z���Ahϛ0��G<8H�۝�RN�����HI�y_먵���së�UE��>��f���R�M�Z,AK&M�����Z�&A�d����.;G�>��1�Qi�#;Z�7�֮��O��R'���)�ѳ�2��_O9��_I�LkFn��"�s���k��1IUŎ��eJk�
�m��+ͨ��m��Qv:_m��B�����ƽ��@�G��q9c��
�˃v� r��)V���1�Z�THDR�")<}�����tL���ʓ��[%L�S�\+���;��vڤ"��S4wS܋S��n�����#a��Ҙ�Y������\�Q�j]�Z%F��]B�6����UW�Of-O��ޝ��㼬�V�.�KUkr<W�T%�@���}G}B9��>ж�8��B�N�K�q���q۷��S��������|'Z^������_R��2�
�k�w�[y��obI��r�ɫzm����n$t�Y�LBQ��K���
��.��}ҋ�*-u�ݵH7|in�[Rx�z2UӚ��p!-�0��t�@O��컎�nY�3�#<�r��r��;o���9�t\�J=��o�=��nJì��*5����D��erZ�}N��6]�7C˞Wm[-�������a��Q�ǻn9QA�y�Yݻqy�E��:w�j\���sg���Vb�+�ݷ��&7�5�ykb֜x�b�>���F��9�}ee9Y3kj�/��W.U!�n�unTn���=��h3��T���á��/����`��	,�-����ݓ�τ�y��w!@�:@�P�K��YI�������;ͣu�D�1�'��s��gB��:�u��p��S�o���*�_8����$���t�RJ	����ȏ-=��:�C���q�V�]�Z���x��������Q�u�uy9Q���Fg BNg��X��G���r�L}�J�/*Õ��}b�o�9�nq�V�����)����z�k�j#b���7�_z����ioÏ��8��=Z�e����l;�/����u���ζ㷛�����7���zM�l��Qg���r8���QKt��Y��"r�_�*��[p��F�}8d:F�|����"���9��8=?�j%���j��W	u�Ϛ��\g4�P�#t�@W��G��eBw��4vl(;'�]J�I��J�Q�O��F�n���ʫ>�q�m|書�a/�����i��}�^�#w*�|��$wv��K��֬8�y�r���ᄦ+��1x��5�T��9��X��]kZV�4�W\C{�\c�O�
��.;v������x�i��^�A�<k�k��C\�����e�k�9�CR�į7왍u�X\.�oF�~�Ke3�}y�e-��fk}j�2SOh������.�ÇDk�m��
���Qb�!��k���%<t;G^c���{�N�m���J��x�}+ng�p�S��g��/�)�ͥ��[b�I�S��̡��j�N6N�r�8��&#�k��P�o]�a�A�1��}N�r��i�K�FF�z=<T�\}ӎ�}��bv5U?YU/��g)�}��6�F��wE�~�}&�y��,/h�- �͕�_mA�ז��\�O��ߩ�Mk���YU�T��[��{Y���;O��P]�L�~Ռc��������O�%��3�f������U=S+ϑ����moâ;�;y�ך�U\��0���7n-�n(���L[��fy=�E3~\��C�/�Î�Oj���&ފCi��e�}s��ȵ��Z��Cǹ|�DL�TZή�:���Њ���g��ۣ�c[�5����\�Wy`Ǖt#1��5��ӽ����^�'ko��;�# ��\6�A��j�'ж�!gd6�7�"�ER�r�Øm�|�S���N���;Ɂ��vh��e7S���#/&�}����wAm��ϒ<���;W�U��]՗j0�)��������]���.&������shR�m5���F����&L�).�PL�˱��SR�����$��mS3&�����$F�{��/zgd���}
�-Ƽ�Pb'y�ې����U7V�(ɚ������ΨM���^8[��oiM7�����ÇeTtꌼB�4�p!K0����__sˈZ:U���ҿ�ݿ��m|�㬭ڥs������[��L�s�к�'f������W�6�O���d��x�)��l\�	�R���X٘v�:�	eA���韂�w�]��>m)�:�I҆�ǩ>�ۺ03����j'�g��Sh�7�vK��-�3�U�%��OӀc�D̞���v��Cj�?���&j
��n�����.�4���S]�4��6�ˡxr��$�ok�M�ʄ��mC�*��T�g���K����1��Ѽ��ԎܫE�����!%r�t��H��l���#w�r��X�M��+���Ѷ��Qy���{Z��Q?oS|�X;\l�wSj�8X�n&�,ˬq|I>��TiJ$]<Ⱦ;�e勥�҄mu��oI�:�r���b#��̖u5������_�T��l57�4�t�8��Kʀ��Y-�t��Vl̒�bz�kys����sZt��Iӆ���]�Ka�r�������/�v�0g�;��-�/�Ҋ̌O(���ƥ�J��U�YY�ы�!��M<�����Z8�B�B��n�qF;�s���J�\�������o��
nv��ޓ}�f����h�m���Gm��&Q�{�0�\2l��:���Ҟ�o^��Ť����[�ڻ�PҠ�[Q�.8�{j�Bv�]s���eR���[m�㷨�[v�힂a�eE���yW%+&����
���YIڗ����׋uD7�
��Mu1ßaNn�8Uް��t��9�Ѩ���.|�\-*޻E�p�=۾��;�$9��Hk3�R�c�����r�~	p��\�73�2d�{��ݏ��1OJ�^�ɇ���i�e��e\@�[Pa)��	���p$%�)�Y-��M5J�
��s�s���掿���_<��u������a���t.\u�8a%�[R\�"���y�޻��c�yg��'r���2�EK�/7����k-Y��^g�$������f�L��oYJӜ's��ܤB�Ao(�^� �\�m���!$)�!���UH�o6��=sC!���j4`�j�`��_*6rg���p9f^��M`y-�Vٸ�����ϑg��f�w{#V����9��W%aμ�o3x��T2�t��C낮@U���G)�*�K!���%�/-�o=)v�y������Fq����n���	Ŗ��rS1y�/��T<��6{h��W��v2�w�U5B��oh��V�Qu��pR!���^|����y,��X1�z�Y��^ӑ�z� �VR��6Ն���ܛ�)�.��s��Al��~�|8�gn����2�9��S����Ψ��F�g6*ݭ�m>��Ňj#�fO��{{\����@뼍;��ȮqR������W�m�lW�m=�K7�����R+���79U�j�\.Ua!�Z����O����S��&��}����]Z*E����{[<�W%/�p�� ��[ƾ�'Z��r�N���p5��1ȃP���;T*�x����/rc1]��7�iQCEe��+�dF�ꂏv��Ɣ�=�3�V+��D\]W��ff\=Nv��p�'�wƯ��hd�SsR�}�W��I�}��F�:�R��O_������&��6��o�u��>g�voc�s��v5�J���T,��z����d���
��s���������!�쯭�ӚO���	O�cz��3.� �銺��[3��Z�Y�1��k�V�w+�0q�p!-��	;[������%�\�s�y�p;���Qo�:�%ބ�.�vi*V]�cF��J�<�LN��L�mh��Ր��x�M�����u�yWR/�*7�{�c�=8U�^k{��-��D�ɨ�O���L.MUwep���ۚ�G>������9B�c�Wtm Vښ|���5m9��峗4l�=1QzD�Ջy�([碩����#dO��Xf�iuE�*�f��}��}�9k��4����n������l��rE�.��\�/�4��NI90R��3�1��糕���Q�wSw�9��OT��;��Am?[]"���
�߱�(�sX�ުp�������J+�ꢱ�oT������r�p��e�RT�;&+��Tmk3 �a	��޵�(��3�kY�r�K��-ђ��e��q�Wq�U���Z�&��4wW+Z����ă_X��@9�̗0&�h�o.�<���Nwf���t;Gϴ�[�ꍎδ�|�4:��Y���.2���^��5���jm���!���H]�Y�b��:�Zثx�jG{;�,��yhJ3�־�8[2+�nC��<����Y%ո�[*�r�(Ɇ��l���Ǯ�{5y{�Ѫ~�����pҡ/��Y���NoY)C���.;o�7bn�j5�NJq������o����P�� ���u��}QYn���\ٹ�yP��E	��O�9햟5_e�({���Ymƅ��N>�m�������s;/�])���r�w%��t�{5ͥk�ݼq�	�xa//.)jΌX�o�~B���U;�2G>���ݭ0�%W�}���Gf����5�c��N�q��,���Jk�`-wٗS����:��CQ}�f�47)���\��f�p�B�AQS������w]�=��1`��ܽ^��tVk��5�@����:�)od9���P8뎬 �O.�)]o��Ӥ�(^��5�30���w�N���9�"����\z�d
��w�`��+��;�t�Y�]"��I܉Q�(�bZ��!ev�t�N�e�ۦŚ˭��Y��&tgg#�xN� �p�����6/o;�E�F��z�8�Pܾ���sN��>W�v�TH��/����9Y��n7��z�c�����v�
Wh�w������|�gK���:i��Pe�^���z{�2��X��EУ����u�V�;v����$��]��j�ի�>�}(p����|��x��7R�WM�oUq��t"�w�
�� T�����+��������0����y�_&�HP�D��iS�d�{B�yر�ƿ�=���2�k�A|6��.H�P�j�(Z2��55*̣��^-�,��Y���^��� 6@9/��̨��)��;v�����
x�&���c�w�'��2����whݨ��u(����yL�f���;(�&:F.�I�v�x��.0V��������U�
��vjs�Q��̼>w�=���[���C_��Y�iCo��m4[��I�s��ƻ�^��/�!�&[e����DkW��t�&�4s��;��^���w>�r�U��1S��=.1�h5M�s]u铻���m�i�|(�ޫJX
�d[���'�����,��/����i豼{�qG._(P��U$��H��k�\��#�i�;35��P|N9�V:� �]�a.��hٵ�.�M�m7;�:�͔�;�&k�o]�]5B�d1�(� ��n�go6��L�[�]�Nlέ��tGL�6U��� �۫�_|��5[��ӫs�����]e��}��:�}�:s{p�h��{�p���L��,��4�!w�����P @�:�W+��p�pu�Szq�1�{3rj�һ2^�h��.Sm�غ�r��g :dMn�ں�g-��;�FpXmvp崢ڽ��Rȩ%�g;C׷�⮶��ĸ)=���F�{��Wt����c;���!+[��d�l�G�5orL�|��4��vhW/���kL�v�]��D��;��t�lV��'��)�X������uf�J�����Bgi��ڦX�w#I�C ���&�wG[g\���V̽uM�ڣw[u��s+,:AJ)��,˺+\�������'ɐ�C}NkC;�IɠćK\�����hCnu�X]�#���*��,��.\[�L��	nD�P��n�4�;ģ'�d}���T�;\މg8�wa1��tf��S�
�0mE|��Z�`�!�
�:��;`���������k���9���;%ws�-�t�_灨}=�F����(8)�9Ɔ��<t��.L�.�.:[�Le��He�K��EN���q��}����e_3ZsgǱsa���X��є2-R�N�H��u�\�vS���m!��ssׯ��������}���\�)(#HƋ�!���up5wuK��wvM:�9p2D�k�4.�-&B�wvRD�sc2ݔ�N����+��.�����v)D%����IfN�ۺ�%���w`�	��� �JI��wa\w%ws9��X�w.��P+��wuˢ������B��.��e����HwGIwu����tP��!'.�6HВ���w+��bQ�ɻ�`Q���w) ��˵��fI�Aݻ��d9һ�$'u�����)t�t20����㹄����}����&.�t�n��|��٦�t���-u�z����YVv�k��!1�zUѷ5Ԯ
��PDm�����Z�u��V�݄� o=�6��M[����su��WeA��¼dS/2+k�� e��a���۷��|�����mC��@O6{쓚��fS�*���u�|Q�I����-i��X����̎I����u���73\�@��s5�b�g^Q�u��*���@נ�(?oSw�=��ٶP[yyN�\�p�L^���AmIl��.:|�~��j�1��eL��Kpu�^wkTWR{Y�s7H8�o+�Sx�6�P����P�c�.�㓧����� ��~o�N��{�zL�}����^!���߇{U��GJw��t���vgm�^&_C��U��
-����b���uE�l�@����m!7i�J:<�_Y�W��J�ٲ��>o�"��S[��}k�o��eq��ˈVm���c�:�ضx׳����v��rF���s����"1FMW*S;M�AR�Zڱ�X��/�3GSQu�p�ոRʇ�d��`=+�Z�s>��;z�q��|�>��b�
�p]�����k1<u��E�jץɴn�ȳ��hru��nIV���u�V��D��|s�;*c���ڣk�;T��[P��dkȕ"R��b��o]�R���b_Ly]�M���$�	�q����ߠG)	T����
��/�Z;dv^wٍ=�Y.�u�;���2a�)l���	mJ��P�l�a��Mz��V+����M�}I����6��P��������|c��*�fj�C��_ml�p�<��ݙ�ޤ�Y}N����]�Sv'�r�֓��z�J��CϽ�.D^�^C�,DOvN7��VTw+|�KP����(��ɻG�j�����j�˳�n@���|�.^ͮ�{��o��|�spA����]$�����C���E�Ӯ�s[Cg��]�y�>v5w�� ��s1��KuZJ��9}C�8��ҫ����>X����"����p��� ��i'�,�5��㽐��v���4:~{{5�������ؾf�E�����C�T��W7s3vLv��ީ��n�i�7�z]��HX�j
eQŢQ�}�Éj�1��۬2�ц���)�]���z�^�9k���������m��U�+m�`��iEӰ+[n���'����F!�ǻ����A-p�
�e̮D�Z��_P�Q7n��T��m�...>{�,���N�{9z1�V�jދ��f�˱;n��ҵ����夼��/R��Ļ��ͨ����W�m���my.Һ���ma*=]��C[����΋���~�C���{��h8�X�o���op�㍭��̀:_i��P���z������_q*.u���Z�Ls��MX�V��7Ѻ-wGKT6�����)�W�T؃���D��}|����ufX|��;�q:y��y�%-��ջq��C�no���%ŗհD�RC�@���1j��}��r����ҷõ^8ɈwI[8ʱ	D��N)w����WJ+��JT\�p��-j��iή�� �6�TC�5TWh��sٔ�x�5g~���9���a]����}��8�t�̓�c��>��iޱ�ҚQo6���T�Юy[�g5����S�jj�$Ƭ�V�<�>a��t�y�]�-^+�һ�8:>���쇴Spû�$��; �wyi?v�A�9�!N�9��Ѻ��Ca��o�+i�i��/������t:]�f���J:�k��Go�	���;��o��FGs�?x��x�m������*����Xȭ3�,��;;�<2���ݪ��&�yU�7�
�P������h���SՔw1LM���Z�"�����vP�P{^���A~���tA.���N�gfhќoZ���_^NTFrkO��m�q���3�͘�Ƀ���9�]];ϻT��|��ɏ�X��R��}Y&-�\/�y�4(�g�3���
�q]���q�m-�x��8qv�Ẻ�t4����rx�<����M������[C����ʣ7����}S��;S�3�(B�O��ctT�r׭�(�w�\�m���d���!��z���O-�+Z�V]�Q������اO>�.��~4	OÈ���%v�ϼU��aC���i��-��G���ݸm�B�o��2F:�t7U�b�{�j��Lc37Ʉ�9�����Ty]��J[v�RϤZ�%J�<9�>)΁+��wع��,]��'n��*݌V-[@�DL�g����Hu���Ŷ�ϫj!�G����5m��o=���p%2wj��
1���.��:��j/�Q�D7�W5�GJ���
i\8Ֆ�a�)+�r��S�6О����Ю�B빭Ho�J�����n�\��f�6�o�r-4%eH��z6b�3M�*�C[F����-wpfpMp��nN[�����ZwβU�j�<gx+n��c�7ⷪ'?W+s�3�����r�ݭ�B�8�M���;��L��`��)�x㣹H� (�ʜ%���9��.�7�����**�b��P�C��0�͞�1�=��#�ەw*'����ɚ�U��,�=���d$�(k)��P�Qg7�M�˗��X��wE�TA���^=�נ�f�������.��-'eY�����[O���B�>�+��0_V@���יWtjK�~�r]I���J;5]-�y���*���q���N)��Gʲ�!JY�V<^�f�U�X1�A�H�{vD�u�K5���u�m<�+�T�#��`���C�U_�OU�y�L\���ʥ���Y��N�֏�!2��i)|f
�'����9� �^I۸S�S���$"���x܆��6�`.D��k3�Mߥa����p��IMِ'ڮءQ�]����C����������Ǉ]ll���R��s�V��z;9��Z�[�˶]e�rl[o3���v��X� ��:5�B/w��޽�s����W�V1�s�OX}m��!���=�h�y[�#^���|�;���nu
�+>%Ȅ�����y/TI��}Koy��< �oY���[p�L�65��*J]{����o���ի��d���5��\mN�>��
��%Rg�ٕr;�',t��Ә�=v�*+���ܽ�ѵ	�TBcu^8���)��]ʈ0��t�vr�������m��?�,����M|�S�4u�q���eLdr�p�aI�IoC֌J,��ٗVT$�L����������l�@5�����g���(UF��;ӡ�Ǣ^�bWd�F'�|Vr�i9p��"/�*Ԉ���I;�g�=����u�XpR���:��4���tt�{�c�¥D�=�0�jT�ѫ���n!��1����ή��,j$�У-ŋl���=9�JW ٛ��-T��]�x1#t6�^�W ��@�еts�����OH�� �/��n���}F�;�
�o�
S���?Y7y^��z-����Sj���,sK��ܕ�6�ۂ�ݰ�=;��&�Sͮ�/U?�\h�FȘ�:��<��}x��V�ґ��щ
uj�&�
�Grm���뾴�(���L5t�Q�5־-ewW�}���@��q-Z���{�B[3�����J������Κ���̯�X.1U�d���;O�0��-TE�ʎ��3�mF&źX�O���aىyT��k�
���^����)���]Q��q�Q�t�΅͊�M���t
�ݭ�V�;	~����\�䦓rmP�ok;���B�!�&Jw4���ݒ#9j�����U蝔�+}_9���v�A�+�Ԩ?N�Qy+�m'D��c��O�Vot��b����[{��}-ʚΉiA�=�"TI��;�!:��� �Y.�W����|�J��[���9�x����v��}٢��V���V�A�Ȯ5��jI��ڐ4��M���.HxY\�<�5k�m���Ѷ��W�uİQ�Ӽ��m��=�T��ӵ��'sғ�:Z6H�M���t�gm.A4չ]vE�cc�*m]_�~�h�e���=�{������_�]�����1s���}�\�V���E�+�3l���1�!}������oLZݘ[3�o���v�������������&7u�Y�&�Wb;��0��_@��Pc��p2���ٗ�t�p��;M0�Tj�ۖ��o0jB�T���7�B��u\<%�Ü��7�3���w�5"��£5��7����e6���^ҶT=
�!�U��>��4��v��hU�&���Tj�)�_�q��P��ۄ��&��c��J/ _qʐ�V�O� �O|�D���~����ܻfՃ����T�#��P�A�o)�6n�X�땼��btf�.,����]��4��V-]�U��V����N��z���泰9�(L�F�Kӻ�nf��H�/���V-]K�_VvRb������z�q\m��\�ģh�{�|�mR�-�m-���s�Q��|��Q�`�Fd��v�Dn-��o1�� ���O#7��f��Z�	����T]��W/U֢'��]�bd[�����mr3lK��7���ᩬκc���ʻWé ���׹,����[9��T]�C�®���PV.NY��I5f�����l��y&����?W��f�H6���)��7�m�2:���=h�u�(SSpm��9P�{oS�������+���[U�S�-�tt�;�ڙ�q���B�av�{I�t�wZF�����yt��*��ӭ�����Ի���F�Ħ�}|�D,��M�<�8]|��2����3��ݎ_>��}t0Rl9��Y$����Z;����m+�q۱N�-�GN�lL��F��Lc�]'#���Ѱ��c�\.uдr�Ꮄ`�^I'�sa�/g�<>�]�P�D�F�jQ5�a*�p���2�-�9�e]�⓽,r�F�7�c���w=�](��g�xK�Ю��,cq��B���Su��u����:�I�Qͫ��{����>�L��)`�M�7*U�\�GBo����K�<{qVRTr�&*�P�ʸuPr<s2(:����䫾��Xl�9d�y�@�(�ͮ�ݝڏY�ů�m��*O���;�<Յ����\��k�eӥ�X)`��A���ą�����JX��k����d� ��#;|���me����(k��+�iR�y�ن�*����7��Ϯ�s���?r�m񳮺��m'��>}�����i�^c���~�X�]��%�Z���۫NB�Fޒ�t��z�ӻ0�^�7%�,_5y���k�f+LoSz�9.��J�8���S6)�Q����<9Q�m��B�|�H2�y�+�y�e�5.�%����W�DeyN.���f����M?r��ۣ���G�W���z8��tr���t�ȼ���䃋v�rަ����ڈm-���U�˗TV��v��BlI�yG8�%?�G*��Yz�i���o4��m�Ak�ڔ�:�hZ9p��h';�д�r�_Ѳ�\ak/����oT��yL<���B�<y:�gL�?W�ҡ2��#Ax y�f\����,�UV��/���m{�Hr?,�(M��u��g��(S!F��TJ\2/�ˈZ:f�Q멝3n���kU������x�'�����BS��J�\�����N�XY��>B�Mu��ܗ,��d�!�ސ�_�v֬�Q�I��C��������왂��Y6[A�6�1��\*��g���0�/�����&!QR�b�=��}rf'���a���#ަ���T��Z��'5;���sp��C��Y{hҊs����鮕�P�[�D-"77��az��:�X���G:Z�=ճhC2�����0��Y��Xtj�W=="���Hab�hX�m���_5N���q�v,v͝=˭m�����0� �K��Uxr��W@u${&Ak(1�k�}��P���q-��;�)��b��U�
�+�%̠`[H
�^�+Ss�#�9�vZ��mASu_p�ppr&D�}	���eF�lߞ^�m�9q������t@*�v��g����sqFj�Il��M�b��֋/)x������,e�y���UrС��;V9���T�q���r� A���ىu.C6b���zq�o�RԽ%�ߵX���׍�&NG�:Ⱥ�b���Q['-�<�Y����X�6=�@�bn��.#�9S�oY��9�5��D���t҇�7�^<յ�R�=�@:�wn�W��2N|ƷM]��	V�m�k��P}|��� �����eXR][�q��(Io��.gS5n{`՜�}�&��&S��]����l��X2��4�;��ݵ���A.o=�ҩ�[|	�7~��$ܦS�;�-�:�d��*Hu��F+�����s����%+H/�V���6��"bT{���_.�X�Y�J�J�*�1��|��4h^�N�i+L,<��K����5V��N��I�kj�/r��[�-c�qlǓ������GW1��mCE�W��a�'��Ox��Q7�b��1���v�S�v� �M�m�5��,
�`H��r�Ɨ�'C�������m�s�{��f�S(�Y��j�uj-
9�\릤%��'���<�qT��i��'�ѭ��V��meυ�AYPыEڃ�(�+,҃����R;@�]�B���8�L+8bF|�U�d̃�\�Jo��\�����W,�^���ob�<(�ֲ(�i�"���˹�SJ�Y:��}��l�ܠy,��&�̧,�GI���f����m[�T]���sO<ShXX��ݹ�3	�3t!�9op�Ҷ��h+���TP�K�����1��M#v��ebʔ�=�6{r�m��T�7{��DLj�o��T�^|�n%�(^WD���7)�bs���z�3ㇴ;�x��_��MWv8h��W�<� e�S���ÑKe�u��t����VM-]��(֣H������[��egbNc��w��I��H���ХER���
�����gǫ��=�ٸ�����əe*��v��>��R�<f�M��"��#Z�`n\�;ku��z��p�Ծ�?0u���)�L���'Z���V%���b�ͺj����V>�(p��\�!L��waD;���cLFu���B ��n���F+�MM�B2�G7\�L�D]�H�`�*d�;��tD��ܗ: �]�ёD�!0�I	m9�u� a.WD�� ��γBfL�a(��reݻwrwqΉ1�#.���`!H��Q�&�ÜF�pL��bc2F�f���7NJE),���wn�2P�2e˙��.�Fg.`�)$I%+�;�B��XJwr�A��w]�QI1("�H�7	�'wwk�����%�rA��ɲc5 �$�� ��nW�������������}#x�v��3L{��}\hN��A�F����m�mm�J)��*�\58����nn��vh������{�8�;-o�Z:]����ƥn-��5�+�`�DF�q5:�Ƹ͝��+�{��w��CĦ��vh��ӽU�;+#�?$M�

��hk�����5�Z�}��5~����w��ո����n�-92#�mپ�lF`�0�_�Pim[�]�Q�����bN^�1�cb�'�i�z����jn:��&93��/3�"ޜX�~\�'6�U���wX��Υ�)<%����z��9.��'��o"s��1U��Ɍ�8p[�{|�8��lcԬ��}�'���2Z�Wl�}�Yk*;ce�t{8Hŕ�1Y�NV5��TL_Sw�s��CC��Ϋy�Q�nU�+51$[=���V&[���:��9_v��g9��˛w�Wͭ��Ҳ �e�WR*i���؋�2��&�Ud?g����Y�=�E�{Ӓ�����Ef�c�7�h�V��j����5���A�b�v��vj��i��/�CF��B���Lo���dCU�k��ie��پ���}P��JΩh�����(�'t_���eg:�'Ot{�Nآ��+�-"�]�,�e�9��o53���	߫��~�\�nK��Y��3{h��@㆖M\�~����a@�.�G�^��r��5�ݎ�� �]�%A�j�,�W:3���K�4��O�y�o/�i.t�Mr�0�aA���k�Q�g��4 B�sqP�����]A�ܚ�������KKw����R���QrM^��b쾭i5�R碓����
��Y-*�f��ҷõ^8�r�Iloa���{��g��"��#�\.t�Zg!�W6oB�I�څ����\*cj��YU�A�s�p2��ٗ�鴺J�q��nj�M�<y+�6���C��<�*����j-�`�+rk�Ou㨬�Df/-O�Tx�7Y:��9֚��j��B�vT�
��Q��x97p�P�ZG�tr��Ђ��ovj;��ܨejb�5�
�P�?kg��հ�Fр�y�>��(:��
t�Ia���sv�v̔�V���e����f��;8&Å���YZ��&wyl��M\������+���x ��0Nέ�t�3�;�)N��"�{��ͱ��D��>ː��9s�9y�/'ed�tm!،Us������{Q���:
�M�ꏚ�Hٳ�Q��;[�\+�bBC�9��1���&�b����Z;�M�����������/3�Zd��_eWoW}y9����u�cD�i�㬜���=z��y�(�z�����O���v��>���m=߂�\0��G7����S��;H~�G/O.nrs�c5�i7�6�'����"�HF5�iV.^���u+܄�<I����s��W��ҡ/��	+�z X������b�-;�m'GK�q�����Ȧ����}v��w~�u���Ѯ��j��c)��`�C��J�Qm>k�����m��ɻ뚂4}P�.K3��6T���{N��#z��v��_`��Qͤ�\]G8��N�]���/v����Ʉ��㌯�Ѱ�OL�����h��p�E]�h
���L���(�M<����K7h�Js����юT�P����C�f1H�ct7*i������ϵw����`^��C���(u�mj�v���3Rєv� �U�<��Ūe���d�D�t�+�ͪ6��"�*6^�٨t��P�Kz�%�|�=���2�s���o�{Y�E:F��eX��BY]3�Z�V!�#=P݀�P�\h���o�j�w�3�:ὅQ�L+�<,��	�pvwo��ĺv�]�<z��ve�yP�P�Sb�<R�W��
���GQݸ��ۍ�)85�Q®�n�^��Qʄ��
�i�*x����ɚ�N�9�4�F���K��
�4����[ӋȎ��*.�9�]��y-Va�S�%�0�Y\���u��G9�E�*�ǵ��P\
|�lM��p���<��!h�Ζ���6�
���.��r6�c�e�n��|��/V���$b�v�.,N ��Ҿ� ��^� [�v(��� V%�ob��s������ې��:-���ii��-</={^��<9��J)h����mY�Qr��u����Uy�7kV�FB55�$��11SO٫q�{[�8 okb;��&�WS��Sh*K�8N����v(Ǧ����0������r��w�}��/p]�2Z����;VW&i��Bm�.+gµSbu��ɛ����^�G������W���Z�L=\�*�b�9�WǬmJ�ֲ�'s�ej+���7���3�y�����&[UŤ*�'�gӥ򆃿t:�9Y�k�b���g��Y�@�{O����^Q|��ν�y����w�k���P�~��Pb%.�Y�kX+y�z��H��5�ni_�eE�P�35җܲBU��l�ٔ�qN�x��{o��G���&og�\&;��8���)l�� BZ^�u9Yљ�Ɗ7�`�U7s1�}u��ju�Ħ�W'��pᩆn�p�WV"`q��Z�9����1����5�ĭypf_�	5��9�v&mN�QQ7ӽ��;)��vĻ�<.
�Km����>��+��A3U6���=P�RR���pP�wa��<(�������:��Ŏj0ú���ȋ1�:ʆ�O?��rd-MC�^�6D�Ѵ;A�w���/c�ݥ���P�����&��N�t&�T���m��9��x�y��X^�6%��Dy�m{ں�`U�2�mQ܂��k���׽�K�;z��;X1�5}|��1�,����Ӕo��ɬ�	\�a�����,:�[!�+9�&�`�Eln-���O�����UN����q�Z�w^ie�뭓 5~3>m@���c�5��/'+��+g����78�ds�{F�;7
�v~ 슧M����-m��U����[S򞎽M�+��:7aGR�Աkb3T���*��t�~���ɧ�b�K\�Z؊��i;�Ʋ޸9��e>�+�<��b`�RC�����<�ᵞ&x�۾~�4���^��q���=!^�A�+��'r�ϸ��ź�,=ݝ���J�-�}��}�;m-���)����am�='c]\OF+�(��u�������>B����Ur�;��Uf[j6��t;J��tw���*[�;�������T������OU��Ҩz7k�qoTt��{��6%���7��cT~�֏1	HK����as��Ի�|���LS{�N��y�hR�B��Bg_jb�<�7�T����4�{��볏��́a�#�/�D��=��Fw���꽷�;2�qJ�#"u�RsG@�1<*���Q��]QwV��P���'c�u���&5��z�J6T�ͣ�ah��4���%.��k�S�Y㣸��mG�9�t�u�ٜ����)��ݛ=m^s<�3�_!��7���xG�E���Y�樵�X�b������_&��|�UB<��Y�����9�=��"Z�������s�p|_ћ���y_r�;j{wہ��D�Gn�L'�Po�fi�����x���j3���S���:�r|ڃ��S��.������W);��_ہ�{b��Ɋ��10qFwSwܩ�1�4~��[9�t����D/'�5��K�}���4�K��T�����{�e��{��N����Ny��y��SmC��v�����7:�f9=-����%t��ſy��]�bm�5��+�بn}<��py�+<�B�`�Nʡ��7��{*��6񼾅{���}����eb#*��qVQ璞�|�>�r�w�]`{�7x�����{�_��:'	�r�W���Y�T�J4����*h΀���ȥw�Le. ,�aG����\�Dp�\�ءqa�9\��R'�����B�t� 	�!���V�ݾw�-�d�q+��:0A��Ad�j�JB�M���}e���O(ín>m\D�0�^���K�X8�u�q�|�O�&
�*.'y���*YN�|�Kyx�n��*	ȜYYKwp����J����韆ƺ����o�Żҭ��h}�D��e�hNs3ՏZ�>׺�{�_ޘ���Q.�|W����el�E0�)���E��<}�w�ԑP�(&r7�<*/��@����.�a��

�dTz��=!���=��y^�K��{�t{M�U�71����r=3�J>������Kˑ�G�{�����ܔ�`\�j����3Y>�ѐ}/N���m���U����@�G��Ep�uZ�����k�1(�f�{ �%�xD��4��1]9&��,{��3�w�xdC�����zjE>�sޮ�*���z������dM3H_��50�r�L,���=)u��7f�0���8>^A������	f�;�G������xc�4E|�%��;l�/�ʇy��7��3^�i��X����~�
�k �$���R���᫁Y�B��!K�V��s^n�u���"���E������A{�Ŝ����w�&ҵNC�R�*�˥h�#�÷�ަ��/��<m�c��=�9�A쵦�i�h�����:0\ˡi��怴��-�輰�.��!�w��S��g���g�wqk�k�ޒ�\D�M�;,e������h��X�E����ux��@`�j|��s��YN�:��:{^u����ΛDi�Y�躨�����9o���X�d�/������r���~�3�߇z����!
��'����L��_mD��>
����ɝ񿺹�;�C.�2E�u�=�+Gs>��1_-ſ�Ñ���c�OӑR6$ !ڏ	��S3��"���.�tc�=*i'��⤛��Mo���[9�ex+����{v���ӲX�@Mw�*�"���f��c���W��9���ܶ{��>�v��x����c��*�~�(���	���7�tP�x[��"|c
��wZcݥ��PQ���uǱ�Sg=�Y�9������3�;E���٣�9��t�ĉy�*u�h8;9���,/��B���*㟭�����=�q~{NO��n����/5=y�.|�Ǳ��&���PKf�
�gKq�v��z�������� c��eQ�+�x+o��N���x��{�9n�ܾV�ǟ&��ϔ��Y�-1�VH�P�S\��u�Km?��Ի�G)Y{�R���]i#\���*���G�9�/7�L�$�`Đ�.�s��;��d�!p3����Cy���:}7 ى����F�����vҊ����W�Go鉄��O��s�ở	C��y�uv}����W��t��[ɜ^�w� �5pC���~�l���>5�1O�h�1��E\6��w;�Va=z��#Z1o��J�溭���@yc��G�����T�n&|��l1כP�Ӳu�Xj��b��gi?�QT}�h�ј^7����
E���/�NH��FP���C�����q�lp \m�Nwz+�G��+O���[>�o3#��E�\o�i�����p�#�^���+��W?��tq%9G���\6����d�7�|}{L
Ig�<�}h
y��{n)N#T!��c�&�t�Jn���y�i!#��_\�(^zkM��@w�5_���׼H�����[���d{�o�W��u���Zj+�bs	�eFV�Vg�|o\����Y��K��~ݫ��=�]�+�d���w�{ס\y�${-�=I:l�&�Y!Y26��B�^�CƘp�b}�\;>�G�:۸̈^��9�x��eƊ��W��=���P,p92���>�,;�ǅt��׺o�5�3�����-ed�4�
�4P�m���r�{�fF�y'S�d�&bc5U��5�S:����-;K���w�DAǼ�g"��T�M-Q3�������
w;Ĳ�Chv�D���kv˾o�E���m���	�W���J�#�����Lݢ����ZΦ����.o��g`�Y�k��%F;X�TQ��
G�L҃i� {qo}�qc���}lK2g`���-�f�.5 ���;u#|M��/u9���qW����Z�1�k����>۵�G2�L�PsSш�^�x�nZ���\)�QJr�T���0h�52�u6*H7��_aC#;����CYi���������[�_)��zh�{�N���	��,��gt	\c��Ug뻒��t�R6hi��k2�R]��=������$YO&����\����P�J�_����bs����Z�$����f:*��aZԝۯ"�y:�]�b�ꁾ����J�T����гp5x�a�-�:7��{�h�,R��N���&�N���y��c�����]�Yh}�Iޭ��Ρ�n������<�1d�` �s���F�Wc�5v&[���ٜ�R��LGn_S�dkF�ң\��B�b�|Y���ͨ��K��G?���tց[��-�#j�uoj61M4"�����F�Kv�������\�����=<��j�U�vA�%��n�㊙�\���{}ߊ���i�rx�g�x�zY�x8�+-V��x$�v��J``\ie��;����~w�+=���]6_�f4��*��P&��oh9�� i�ڐ�_|��s9��,�(��|C:��-feۋM�hwV�bQ1��}���X3�.Jguc�{ ᯻n��,��Se�k�`dXZ]1��ܖ3���Q�r�]>Qnݨ��u�!�J��^Ix��lG7�gJ��xtcK;��p5��OB�&��v�d���8n��%a�@u��J�u�B���U>�F�k�p=�hw��]If������bVAܮyQܙT	z�L渔�nrfl���{�1��rN�B�-'��s���ڶ��o]qO���#F��Z��2V7���EJ�����6��*]�c�N�в;aF]�Av������YZ�r� 9#�����Y����^�Ibh���_(�V�Z�&a�n�8A�e��Sq�!�+.X���M��%�sJmYm=��\+'���d�����o]��4�3_���z�w�1Mll�HZ�ΏnX�kv�Ij��w��u:���5���*��HH�=cb*�4��]3��6����0�U�Y&��²��T����Ӎ�4,��qՖ��}1ҕ��!%ȭ��,c/��&�ɍ�����������PԀef`U�Q��[Yr�Qk"��n��v�m]H��k1�+�m>U���3���V����S�WX�cG��-��}�O��=w"!$L�9ȓM&&	�,��&
5 ȋDE4��d ��J	�(��\�eCI�1* ��&��;�
#�3']Ɣ���ˑ��$��I0�H��Dc*F#&H�%1ݮ�ɂ(���� ԉ$s�]�A.u
��k��wvL�c��r܄�2fBdЅ��H��@��ILbE�cR�ܥ۰�f�+�
L����q��Q�AHLFI������s�wH�A&DH'v�)9�2dL�H�DL�!M3.I�R0�����
��2A(SK��!1��d�b;��2$��6LS0���)@��vP�R��b(Ԍ�(��@� 	��"  q����%�:OɺW)�j�`�|O=Cs�7�S�^Zg�m�0���A�=�Sc�a[Dmui����f��W��ǂ��S�}�/҆y���ϗ�=����{ҼR;���`4��נ
{.��_��d��)���:��rOx~��jy�Qs��-��������`��/�z_�U��ޘ�w]��f�T{=+�mLMzlǡ�^#���#�%���௖�K��X���ۮ�/�Eg����F��m������<��D�t�Q�+԰�-fC�nR2� ���3���O52�X}�r�@�>������u"�雅�jz�d�Qjbb�W�����v�ԳD-�w��j���.=��=ޥo�Y`���~ ;�n\���$�|�B���_6*k����;=�fx����kxgvg�qh3�7߅G?*��c�s�{@+���4�}*M���S�=�W����� ���v^����H�����n|jc������Lza��'��+a{/���cw/=�O<�����뉺���+��=&�;�p3q�Ǔ��z��H�����S6Rӽy[�[SΆ��T����7���N�/\�輟i�|��}	_��V}cK'�sb�(Wu�^�7�#Ҍ7�R����/��c����ܥ�c��ŕe�=Q�k�i������L����S`a�o�f��m��[���
�mN�U�n���}ų�έS{�u�1>,�������Hg���;εe�Dh�8rM���+g/BC����v���@uC���b��ռ��(��R"��3^�6Z�+2���@��c��OYiW��w�@w����:�7޸�^��q禴Z�:t�/�bKWYp�N<W&v� b��&��j}.|��yLm}����m�n��Q����Y%.p�\���»<��*=#Q��S�T9NGS��ϯ��}��]�F��W#�l�[�73��N���ǐע����@�����x�nL���H>�T�>gF{ޯ#�����b{b�V㻽�읔���z;�<a^��5���*�S���ݔ�٘���J�������[�g�F�U�[�G�wܩ��UTGM�qؤ*�'��\��%*�n<W�܇����2�9�b�c�Ş��eo�_JG�o�|;�7��~�_�9$.����%;�Ez���J����=tu´�x�k��"Y��B����6��Ù؏xJ���Ϝ˓� $v&
�xxs��nz�ex�����O3� �-6�}��7QK���r=3�J9��<��ˑQ*�N�a%W��N�h���k�|TÛ
���Jj����7F�E\�8_�������<��O�a~[u�VTdL��zF�w�hۭy]�`��,SD���%MQ9�]o�Zr�[�z��+�W
7Y}N��viI]��u���E"�qb��d�`1F�z{����ޘ�ɩ�f�u�}>ӹ����G/���L\yK��ϽZF������y��d�k2��=싃�K�M\J�)x� ,��X��r�w����m���_��ehO$(�ʿq��:�|)O�� �z�+��i�	�;su�+t��OI�8=5��c�ޱmx��䢻�[[(�}m!\}C�y���D?z�M̏s�����r�X����T;���>��y�So'ok\�/}�Dϒ���S��z���;��G��qp��8{ģ}2��t�gjsk}P��a�u_%��G���r|;�r8�%e�"ҝg�Ϻ���\U�Tp� f�_�ߘ���m���'���b��?}>�����%���P�NCS�;_����V3�>~����;�����������U�4z��x°^D�����Mib�&w��u���~����$T_�?U�)�Bqv��4}��g�~|R����(�y4ϑ��������ZY����u޺��{=�MxE����;TjZ+}�}��4{�>�]����1��d��!��٨@Mo�N��=���ٽ�������Z���6�e�:����ں���9k��K�b���,��,�Ws	)~*������z�!�Y{k��4s�dg:�z}yKP��a4���~ή�b�m�F�*Y��K��7J%�p� �b�f:KHԷ���B�b����+r8�\�N^!ܡ~�ϕr�yW��v#����x\:�lV*��[�&`}7���:������1K�kRg�/h>S�*��PQO�Q�=)���}��O���G$��@ 6Y�Y��k�Mt���n�T�ɿ�|=���OD�7�H�?x�~;�t�{-�i�$�\�JƲ}���K��w�#�`N�t���L�J��ݎ�=W�hM���{k��Y����zwg�a����y���vdH�ezdN�ӄ��ZH�]��hr�H�����̡�/�KzrE���i�J��i���p����,o�+�hZ:L=5�a�S��7���z�w�l�5t�D��"SYU�C�\+E��Mx����k �(���T�I�Y�f�q�P�y{�(yG��$�>e��j_��Ts��_���>�{wb�IߑeN\���[u`�/��Zw=C��b���kB������ɥ�ǭ>�����Q��ƹ�n=�C�6{���W���E�[s���~��}��$��n'k�������������3{LJ���կ;�A�����R�kG��ث����Ua�!f%�3i�uǴ��5�s9Y�OV�Z{��u����D[_�ӥ��
ER��٢u�rM����Z�a�<��1�V:�MY�j,w6��= ��qWBqԽ픱�9.�r�L���jP]Q�iZ��wvQ���R��}ב���q�y�����sL
������Tb��zH,TW�#��O؟c���2R�;ܩ�Mh��wMė��ۯYv�ץ_��Y�y�_���s���Vs���ղo���v���W疇�-��IGn&X��!Z���{�'Ά�X�y#�x��=�������Ds��������K�]ｗ	���~���@=�X`��l��~��9=ڻәevn5�`=ʎ�L�φ>�~9��U�f�SӞ����'�\Ҩ��Y\�3|l�u?u�ۼ���`+>�\��u\��rn2Pl�=���^~�'%W�ў�+M��M�y�Сs�u�ږ�yW�k&Q��މtj>; r����[(��
�{�����B����En��[�t�ڠ=(ߵPM߲<1N��<�CsPO�*��+԰�Ĵ}����Y-
�{�W*6��z��;�����1��{,gޖj=p�s 6j����\�:�lݒ�[�G�S+�N�����U��ߎzv���_ �r�T<�t�����ǡ=}I?t��C���\�ʣ���9EA���B��〈�{3�4�vΖ�0
9�6fD���c$�_�����qJ��������cwj�B�k�ӫ�7K��Sd���K�J����P��o9KnI��f�Z����G\U ����!�Ru#�#�y���F�H��'�i�
�\?+��g�O�@^�ʉ2�}%'{Z�V�=ҧ��$�)�jtg����i�Q����F^��;����G��yN}.pz��׃�k�����3���3������>�M�䈔;den�y>&�΃5k��c�'�+���<��ۖ��w_�	��?u�{��1+ė�N�/ten�w�^�qޞoi�3�`y�����ܶ�����=�=�}��=����I�-��j��T;�ͪ�Z�3'S�c�]Ǡ���\�9� +�jǞ'|y�n;����g]OMh��t����s��o���Y�*ba�˾iX�5�/��z���7ӍO�k�x��g�c޸H�y⸫�m�7$�����ڇi�f	��==�U�X��W��W��d֞�ɝS��s��걹�~�q�X��;�q���n㺷6�'/��纖]���8O���Ӏ��Ux=����U/ӛR��uA�����{��;;<j�]��W웯OMo_��u�g�϶�\n'�Y��(��T�U0&*yq�77n��"ב�,�w=�c�B�����I8�feo6��2в4
�V�Y�xW��G���z�ͱ�*�T[��,S�8��1�;z-���{b�}	 %~�w퀁dJ�n��1�<'iY75��y�.���BA����s�|-�ĳ³!�&ֻ�X�g��0�^M���Fh7H�ѩ	���\{�`u����7��u4O޸��&��M��x�����z7���/�n���AG^�C���oO�vo��z�/�U]��'@nn�42맕J�"�QN{{�׬t��܇���\U���s��(�w�pW�ԇ�W���Y�́<;9��g{fw;���Ǥ?G��>��i�]O����{"�=J�F��q(߽#K���r����so5	�i��`粏蓾=s�jȚs�:2>>��r�6�[=T�����\ߑ�m�bul{s4�!�׸�]P(u.��ȃ�nZ%ɥ�B�Fƹ��FXۈm^Q���?n�V�9q���V�X|yP;7�(P��/x��#�n@�C�E+�6k� �=g�*Ю���o8���p�Ϥ!�vi���=�ePc�p�ģ{,v��f���چ����L'5N1�=�0��� �{����~)�ׂN����'p����'~��p�w���,-8}
�%�Ìֿv��o����d�l�iL���Ζ-�d{=��Q8����:�n��J����^z����n�����<��J�ϗ�E��Wʀ��'��B���IGD�����X�������j�[v�R�s0�|'#�6��7h�/c��,�Dri�u����U��>�<���U�K�FpI����hWCV��QV.��� v��jv"�h�ռdq�1��۝�̃:�쩗
��Xg�J�蜟;,^�֕��ð���ND��{<����_�^���%x��p��jhM��_\��<�H��.��2�&����� c�롾�^�#�^g��Ɇfpno�xg]2������hv}�Q���)�P�k�N��[w	�H^�3��l�/-�F�KV��z}�}>�z�c}�P� ������z��)����mUa�%��wǖ�BG����GW��g��/Ã�T�B���2]x���8��ڂ��]�Z:}�Z��e�7�Mi����~^��ǻ�>-��>�r�^�(��?B{1�=��^2�����>�r��H>D��c���!;��M�[f3�*L��@؈�BŔ���g���������4�`@B�K�������m.�(gC��x;�b2 �_�׋�z���#�~�9��6�0q�q�a� o�H��z��n�i�=�5�����WA�	�Y��G�]W�=��J=��� ����L�z�dƢ/�bi�m^b2׺gҧ�ȸ���ƣn�iڻ�]���moWZX��8��FE�zk}Wg娈Y8�R�rC�����Yŏ[��;r;W�7mA�E��\�m�5���%��7�:c��=�j�e4K��z::n�XH�`NE*�<R�Ƿ����خ��>T��� ���d<��$��l1�1N�O���e ��w�;��?��~[0k=��o��N�F��/�@������'����0 �O��s���J�d��������3��3)t�O2���/]�1��'O��װ�R���}���m�4/|h���iϤ�����?a�>�'Ei�5��P��#�!z���:��U��t�T�Z*n���g��F�U����nt����H�9�;P��ŋ͚�k����~ ���G_�Vc�ɏP���vڷ�<��	���<���BEF>5��	�$;>]UFV�;�WY�`?	�>[�^��ΰ{殄m�}l�g<wyz�/;�4w���K�x�K�ΩT��r^v��(?,�uW{O�k^��'%�}���r���{��+�=��ׯpߣ�:���V��y�w����[z���`�́��w�L�O�|����C���y���>��~���OtKw��'�!��C[��vi�5�6[ 'Hފ������%ͽ����Z�F|ΏpS�sqȴ�צf��.lѥ@���]�p���k;���K�Im�%}��E���/��ΝN
��)��o	�E��Q7[�[�l�
�e�@���r�N�u��{{����E��(${���(��u�E��GK:�Y94��궷{���~	�]�$ŵ��m_uw�A���k�~�FP��!�6B^E�t�j;�}$%�X^��ޯo�Ƌ�6j�xN$�K��S��{\���~����y@!��s*Lt�Xr	h��9��*N�z���K��׸ć>�������8W������p�s���؋SB��j~�*�깝�}� �z}�L�=�c�*=�*۵���}H�5�~TD��ғ�,>-b��4�6�a^�Y	��#�?C�"��Nh>gt�Ц^�o£��ߏ��}%D���tIg�ë����δ�V6���IG�f3�nn��TC��ZdV���SLsTj3�϶�;��+�!C�ܾ�#q��)��7�;+	�e���I�*����/�'äֹ�eu1����&=p����w;�Z�8%Ǣ;ޡ=6��c��T�*;�V�څ���k�{ǁ��+������w�髍�,��� z9<�ca���I��Ъ=�n`��D���8Kg7�ڇ��=�}�h��Dc�����>/=>�Ǹ��u�D-�_�Ͻ��Qϗ��g]��֋Y'N���?D'Fկ?f�Y����Fi�RɍO�ƻ(t���m�]�X�)]s�C����F"�st|om��ϡT6���q�U���;�q����V"��ż9��RF9C��m�M��޶)E@#�,*B��[�u�\�sW�t��Ƈ%@%y�.f���`������^���􎇚��6Uޚ*��v�r �]Ε��GE�ͽ�X��\��8�k*^�ǯu00�;�!va���aUkL��x�ɏ�ය�.v����V�*��fd*���0r��9�S�yf�=J��T�����J/n�����җ������f���5v�[�ֻx� ���M�S�����Z7f^=�y�Ck�<�5e�g�J*Ri����R.�J��.]fk��r��B��ι�+�GXK^���u��T⍓��qKY��pnش8�M�i2F9�C�N>%�`��6�ڵ�]�cα\�+`D嫲8�j@��掭{\������{ .�cА�u�o���0����n�k���1%Ӻ�#�5�R�nK]�+��&�t����Q�3,�0�]on��U��,!
�omd�E)`˽$�c�r���&'|�l�ej0��9+wf�8+�b�uY�>��5��3'dU�7�����1�-�G;��U����� ��0V7;��j�$v��������j��r�z��\�^�Α�*���ʣ��v��4��r�I� ��L��g0�p#B�Ćo�q�w��ۭK1�n6���{u��D�YYks�ز�ڳʢ�<��խ�><��P)'Cv�j#v^Sj���|�QI{l�fpE���絙�È��1I�cK�_�S�Pu�S�5�B����i+v���4^0����3AǍKy��4�\�eS��YWX��JOح��}��v-�5!	\���vi��#S�_��v�װxة�0'h���r.�$vw�K���e%N��^Me�Xv���X�c�˸s���ՙN	�)V������)�k�����ʲ�'��w�S�B^��f ��S����	�@nq��<�,\�hi��z��b�������0_t�M��vȨE�Y�l����;<�v�=]��u,f�ʚk@R6bB�b��Ѷ���Ƀp�ct�
��z����{���:��
p�h�{������5��y�iB�-�;�`bY�T��F �`�lC�h_���*���k�we��t"^��+����Z�bC/^�h����V���n�p����z�l����G�q���}��z��N�I���04��Ѹ�'4�x,���ַ�9��K�r�-��ﴼ�܂%�k��8�� 1��8U�7�,���Yi�O	)�;c��_:����$�BI��D`�F�NHI,�\��d�����]&h1�a��(�9��1 �b�Dľ@�I-P�)�3Dfh4�A�5"d&BPDFNnbDL�]ې�� Hؓ�	��� ��i�0RYL��r4Dc��w\!�$�
�LD�dH�ĦS�PDhh��)�$��XK4�I%�61�M���;���'w!�4iL@�(�C�Ŏ�H�1HF�Fh�ɒ2HDD��2D(B F�-��Y"Ƅ,� �4R���Dɤ���1��"P��L����P�%	m�$�R7.@�h�%�"&1�F�0j��!0�M��"F$J?/^�����޾����y���}�M�\�MC,\��]��
s��h�t�48���p�<�d��;���Z[D�\����;�w�r�乩���|n�����7���R���7�j�n=�g�dn�2���\�	�w�{���#��6�W��:]���8�s��M�����}�T[���Q��xIP��nf mf����w�O��'tȇ8]Sn{Ō'_�{n�=S!=3�t>��p��=s�ȫX��=i�S/�[��6���<���_�<j$��3,	<��XS.�{w�=P�@���5c=x������n�do�W����n] �)��;�R�٨bb��MT�Y�<�Ԣ�]�;�w����5��8�M���7��~�_�|�h����<s�^۽8�gM@���2J�^��;���d�}���P�+��u�H���S9��_�܋���%���e���Cs�k}�����}���KG0�]/�ؕEz;ֱ�����ǽ#����gl��d��{;����9>&�O��غD���tdA��:�c�!�g����
�K�w�2z�&��*%z�g�*p��P)����3�ܴJ�$GlR:/�û!caU�!fc�dw����5ws��m���vjl��-aH�O��6u�(��5֮SFr�f����K�)�E_V���IP�*�⻷�����5|+]��\^�ɮ���J+7��Ax�j��!:��A���̽�wo 	6��s����!u���jf�3sz;�za���m=��g-pD:>z�CioQ��G	�I���U����y���=P=�\�}�̈�i�(vH�vF�yd8"�Q�v&��t�z���=\Uy�=�3�Ψ��?:� ��p��%%�̓6�~r���cs���W���7��L�^�{��̿^�/��z�q��幑큓�o�%�̭�|�]�e+��(�s���1��������'kf��ʗ��z��8�%G��5�θ���]o��Agq�\�pk�(a/�Js��^MiW��ZW9�_j���~Dg��z��JEZ��Ƣ�i��^��}�z�5m���	�$zϗES�t���;�u�����:J�Kәq#'��v� �Ro	�����s�W��_��Q��R=�����?�t��L�>��%7mw�a�S�;y�
�z9��؍Ϸ޷�}�������Qn�ȕ$1�v&��bU�j�"I��߻QBw�~�����~6��p�'�ߴ�y�}=��a�R�S�Yy�	W-%g3�&6v//r���$���Q�+U0w%2�ՉF�O�����9��K=�7�����~by�@~�꽬YǠ�t�B�վ2��3���U߭�5����Kn��^�e^�8���v1�Q��^����������3W��q����^��@����.�k؍s-�X�@j�a�-a�}��m���x�|ʢs���C��6�v1Z�XEx�^�G�sꑐ\�N<�&��yʐ��ُ=Z�l{�td��ccގJ��u��GI�Fe�LL7Qt���V��x�>��t��������rFL<��>�|���ܺ���o�w�̉)���9�9"��� .��4=��h;��⽶�5��O�o�I��cc������`����#�p@�w�h[8HMx�=���3�\	��������g�>F���+�Ǽ��p��X� �#��d<��'�|�w�,z����=��J�=a��������>�Д�7�v*7y�͗� N�7U�g�tK7�OaƋ�~�N��������7�ܠ��ͭ��}�ƙ�ŏt'���^�.c|���h��,�ɘSK7���S��};(���¢$����v�?_�;��:+M�u���`JW�	@R�4���*�*�m�f_�>�{,��dЭ�Q���nKgnv���{��Zo�΀�_�>l�ٷ��j�!b۶���RF|���9��h�+�(tk�Z��vK��UN�:�:�/��{�$�i��F`����ΥJ�<Is{��ɂm�ȫ��L�ݎ�wu��xv�p�$�zV��d�-���!�����F��Z��;)NY���QX��$���d^�@��B�o;8�ӌ�_\��P�(nw���?���n�_~η�;a��M}~���l/_y�b7۴��	Co�0��k�U]�Qqŕ��M�U��/o]�a:�rXL��N�7������k�e�q�����-��B�%?�n,��5���K�t0}qU�LE��=y2��d>�~%zhy}��o�ǋ�\s�>�ӝ�	�OJ���ϵ(��B�|�c�^��N��XS��o�7�۩�^�����:+Μ*���͋�}y5s����fP�����:�\z̳�%ѣ�+��Q�[(�¼^��{���L��]o�*=7w��:9��H{�/h���t�����!N��<�CsD�neI��*ϕXW�0�b��v�>|���u�/֑��ґ~��W��e:���W��ρs� 6l�TD��=�y��>������B5�y����?���V{�� �nV
yT�I��F"���M�WyUԇa��,mE�"��9��wNG*�ǟ�ƯuW�������[@+�����U�1w�ޮ�Ppx�G�vO����:jX���27\�b2��v.6�񹀴R��'�M�5�J���� ]+��-���6��\��Pē����vy�[�������S(2�*/]���:ҽ�'r�J��(�����c�7����j�[���V��uu^�m+�7��.�h��T΂�^c<�[;�}�Z��&�E_EB)7���NciIce+�f������vo>,�|���e�eA)���v�A���"P�Wg�Txt��s��|���:��1޻7>�iu���d��T�ǔ�s~{V<�̂7�%a�=����T]�*װ�>
A�wV�f���h�r� {��×���9ޠ:��˱B��Eh��I�-��ڇ��<�����_!PM�B��z�q��Ui�>G��:���<�;^�jNG�Pt��V��=5��Iӷ>�rNԕ�����e��emÿ�%������Ϛ��~�~��{����}QWgƣθ�Dr��qU��=�H���8_�^�kK���L\Os�.{�Fr~���~=ǲp��`��Ob�V��B[녟r��YD�n'Ӏ��T�����c	��Q[t�Χv���\d��s���F+cs�s������SG���{���q��Q�Q�2�I�*n*�y�S.GW�{��D���8�|��bA�z�/AH��}l#�&�*u
��SD���j�W�lY�+�����*//7��d�L�=�<U��~��Sg#}�=���4?W����pnvk`�%"GEψ��q#l콗�)��	&�M�D!k�M�B�Yw���õ�:�����+�x�J�K���^d�j���KF�nK�Uz�f�I�Z��J��Vu[e���F,���E�o:V;�
���v���c��X�PO�*�J����>zz˫S��s��9�dЯ���7��}��
5�Į*�߱��O"����pW�~�	��d�<���=��~�=�@^R`1�U@3�o~��1u?ku��W[��L���la��������Q��e�o�ݗ"��T�rKG�baz��4�tdl���������O���׾Ӡ��O�dǏ�Zs;>�ߕ��u�(�9�u�|Lo��m�s��}��W+H����=A��H�j������~8|�yNK��=vA�4���|���}�[�3�~pi���+���|�\������j���s'���@ya�ك�U��Q˙c�ohl�k�U[�������+p|���I��q|L�^�?O2��K:Wz�q�{.���iEɜ� ����V�x��Dk�ɳ��h��d�lޖ=�7��?vr�Ǽu�#�����H�>�9Je`|�~o�m���ܶ�M���'���c/&����
�p���NF��z��
>26v�����'n�����������|k_��*�^6o�/�ESQ�ZX����@�����+���Ni+�Np��Rx�4k���0��E�R���n��P�*ށ�-���|@B�mr@"�	�sj=IN��%7)u��kˣ���潉:5�f�E�����:�4��Өkmd�BD�����^m���uل�G��ԙ"�1�W��s��>����[e�����𞺨~5�+�&+�K��0j2*�V�)��`�(��U��ӳ��~�o�^G�s��]��#��H,�be��S��S@r��u��Ĭ��(�0�Gz2|ϯ��p�r_�ǳ���w�3����8:R�B���c��4��/U"FN�y#s�|�`oL�+޿q��v�^
eוG�JE�>;��}>�l��	��s��g�����)}*|�{���5dW^����ǙŲG?�+�M��1M��y���7��}�@->�9H��P�2}%g�ba���F�^+|\��}^6�`�jhz-qO�����Us,dy�.s�a]�ܑꎄ7��� @�!+Ib��ܸ��å.r���q�ޜ=�'Gy��(zT׏�J��|��=�T<�M�Ih�D���מڏSթG*�}���#���=�Q�ґ��F�鸅���ϗ�_�A���Ps�"�z��Wo���TELj� O�pX5�c��u������))|S�1��F���@y�<��t��]o���1}���-���m�kk�Owr�O0f�7;���p�Ô�u�ߒ���#1��ba�o/]>��ڜ3���\�G6mg���d�Xf�b8k��.�-�]؄2��8�EGO�㘺��ٖ[�����[d.W�fA��Ӥ��aq����8d����Lq���Ǫ���BN��a[�q���{5s���hڟR>��븛򣆿2��3�K��������/�)�2x+%5n�uͫ��{0�RV��X7�=�ՈN�5���8c{�{MĖ���w���,^l֚�U���xn�
�\.iB�����/�W�I�ɸ���%7H`�Z��vK��U͎�9���K�5A�Ⴝ�]D�5�^��}��7��t���pW疇,��<s���5Xr���}�=����E���;���M�O�g:��nC/��;S�uLg�D7�y�T��:�RuJ�����^����P�=�^o�p�2e9�}R�\�U�h��>�L�Wu�;ff���)��=u���]GA��ﶭ\n|��edl�(�OH����G���� ��8=�~�=x�`Vxg\[>��j��������ǔ����G�,�fC�tG9o�^�_�D������������%y(\�	���|(_��lg��ǳ}@mC��#�qW�C�Cs_���&7�Wq���g��_H�i�JƩ��}�ex�}A>��CAve�&��t��֡��R���l�Co�ͳ�ΐB6��u'b<��5�R�z��I�|�����^�2���2��zO�Ϋ6튺@��}.qKS�;f�mc�ۑ��(:m��9�Qr�O��ɕ�ؔůק�A<���ķI�I~�@�~�8,���g�ơ�#�Y~LZ�ޡ}�v's�qW5>���
g�ɠ5Ϭ�>����p���\z�ߎG�k�Y������{MM<y��/؊���$�z}0X�Z�'�s�w~;���m?��yUx�x�}$w���8@�}�]�
�{�,�P�\�l�4v���;=$>���F��;��q�vn6�߽Զ�彜���`�^������q��yIg���}�$D��,)]��Q��+�s���6�z�׆r}��~���9lˑ�����W��z|���C9R������~?R��z�ԏ�{��/٪\R=�&��槁��/o�
����ȅ��Nw��{.�<��N�S-�E�Ew9�]��P��c�~�ڭ7_�M�u�|�������G!{2�gT�M�����iD��v;�����8_�at�p��v��5�Hr8���'ad�;��w<5����>�k�t�V�Ez�<m�#0ϗ���p���O�,��,��z�;�����K=9鹽������ {H��7(�<�2�M�����!�x��2�9��g1������/Y�<�u��2-��lJl�����>���B������y�CC���H�Q�v����P�j�X�r�*�r��n.�1�yA��u�Nq�|�F
h�"M%k�E��u�W�u�����ב���V%#r��}s�,a:�3�<:�J~.=;>�[{�}yl^�8�#���O�܈�W�ڬW��|c���5'ȩ���S����JV�^��(*oTvy}��ޏu�7�>G�O�`������5H1Ч���ĺ5��\��S�0��Mh;~���C
�t���\i�yd{Y�{�NO��z��?{���Ν���ǯ�VM�i��������b����Qޤ�KGۏ�
5�+�s�H�~��g#}��R��'��U���q��}[.@�:D��<�n&�U
�.|�h,-8��~>Ī+�����V��}��S䣧����V��+'��L�����uN��Cgzba~��LӞ�чҴ�|����NaC���\'�yW�f�{F���1�>�~�>7{�P\<�ID��Z;M�>���1MN�>����^���;�<[=÷�ͱ��W'��Mx��@�������,�gȫ����ӎj�yg���_a�y.O�J�긆�Å�v+��z����r/nǃ6d���(���&����W�g�^;��m
�:��qk�$�Q`�vpBmπ�n�&��]^�c��뮳�rғ�nڋ�k�SҰJ�/ �%��C5v-���m�c]"R�۹gu�߹�˸�^b=��  BNǝ�͑Io�%YN-w�]��w_܁b؛i]:�Ӫ�a33�l�L��\�Y}̊�.yJ��ʻ�M�%@�9c6�5�n8�(+]�%\A�g9-��U����P�� v3�L[;�T�սK]&������Y*�J�#(�7f�[謤��T�ִv���[w���P�h�+or�-AW:�\r���6�op�D9�޹�ňPzFS�PA02���.�(n>9RG[��ĥJ���TR�v=�<p�owVc�s�]zSky+r���+p[j�s L��Z�ڴ�=��]H�#��ɇ!庩�*�e�3p=:�*u��rM;d�r�<���H�f�mcVk4nq�[Q�-�fY��Wq\"��펺`�I-&��ז����re�[�y�X��L���)b!�����g~Lp'M�{�d�,��}���\��[���0.���V�����=\�S����,�]�Yݬ5av)v��z�.��3��u�g:{�`�BP}R�,�2��H�I��/7Q���׸��˖k�e#h4�W;�m��נ���.��5�)�3���(�݄a��.���\$vuv%۔:��Bnn�DO^��͞o5����b��5�����)H75�,j;e��sb��x�(܍◴'�.��t	'x��6#�ǅ�k�s9\�J���3H�%�M����k���e>n�3.M%ˈd�����B�[X��w�r%Y�ye�K!9ϵ7���'�#��jo:t(p�[V�زgRs27��b���׹���%O7a���p���Z��7 ��-]wy*p��:���[��8�X���Hގ�>��+�2��,�df|:�끍ԯ+��iܓ�J�>9��Ձ��QrԪ�d���T�ᐨ�*��bq�����wa'����l��ٝF�$��� �����$���`��MϧP���+����\�JcQ�`���wN��9�!��|y��f�f�d]̝�٦����X+�x������S��A	�5�ǚ/��l��(�]s�<�9�L5�4�Qp-�N����dY"���)�[W��WsⶆZł�d��+�Y�kk�����fS���D2\�EZ���J�j;����sc:��^��xa���A\���ٙF�����x	X(��}FM��Λ2��Vo"e���礸	�H)�Cʶ;0\6�[��i�8
 q�\�Z��-��K�t�e$a��=����we��tm�שB�����E̻��h�{�I4�<̉�K{�V�Z��SkeT\:
Qy�M��)�j�=�c��M�ׂAˋ�-���[�d�ڮ���t��fg��x�c�t�ѣ�P��U���e,����:֝�NN���ʔX*��\�x*9˝q��`x����Slޤ��3\����ș*(4�
(���#DF�B��"$���*J��&H�RIL�ɦ$d̰d��Ji`�4D�$�#D��Cb"��`��H�@�C�$d�L��a�e(���b$BX�#�Lc%��KI�`bD#c�S,b��Q��f��6L�c%�������%Ԧ�Hhуi6ML5d%��2P[2�ѱIA�Ql�$�i	,S&�@��X�&�b(ƌ�ih��"�1L�bcd�R%	�ш�X�Q EE$hd@VLbLQ�(�Bl�ьEQ&��E�A�!�I�E,j-��jVta�aT��d�ߴ� f���YV��ky�W-��p�ken��iVf�F�,g+�&�"3����Fe�Sޥ�r���~����	��JO_�/���ۇ�i��xk�Q�G:�Q�{ۙ�-�c-�{��r��Z�S||�O���p�_���.r�n4��`-�\{�ޮeM{=�ʟ(ٿ9��;�1¢<Y��sn&���J������e�ϭ<=7�4�o���U���+ܞ"����ܥs�}�z�ޜҹ*�ו<c�`��r^,��2�ɭ,^L�}�__��>��y{N���k,v}�x�q��{�k������[e���n$�'����F^���J�Os�o�	�c	�{Ի2%�S�k��9��ב��z�W�����!(u��ū��l�u96}���U��Sd���念 ��xW�{Uħ�C���{����8[�VÜݓ�򽹨�|{�;�*����� O�r���i��7��of��Л�Ȝ��l���,�9��j+ܧ٭{��a�z�<��&�x��= r�T��.Z&�X�:�HJ+�]��;\�u�}㞨Kr��jS+Ն=�T�r7�4�{-�<��������J�S�;F�=�V��ɮ���y~�Mm�Ա�NO��K���\4K�)k˨'��c�T�#%�uݽ�w�"1*[��d�=gt.$�[���ȽBM�rcw-K�w}�}h��N�C�3c�õ�	B+]���t��*k�諭$�n�^�����R[G��f��Mu�k��9�%�޳������+���E����<�=��0*!�5
�h�����E�&2�썞�^�k�/n�1�#^����G�U��i��=��z�ו�L�yӖ�R����n���	�G�LV�v�3��F���+��ʯ� �����{�Y
��9���.xO��P��TߥN��6��!պ�5�l�>���5	ب|�F�?:Ȍ����1�_pIL_O�}�*I�r�{�|E�����mxM}�ƙ�],z�<̏`���/fP����.�쵦}��9:S�nϿ̽9'����x~���>���Zo\�sN�vx���g�Eu�y��_d1��V���P�Y����=������v���W�����cn��9�>�'�������@r����7�I�m4J��ޏ-�(^�5��	�7^-Y y��S�I����1�*zc�����5�^��O���o��Wlz�:����G��B�L�.�8��B�������7Ǎ��˟EX���;�蜟�K����~�����e�q�M��s+�cDL)Tv��	��=���;�t��{m�@��w��ă1c�,U�Y�i�o����|*7�*ռOo_�4���#�M�)��+gq�ْ`�ީ�k�
��ۂV��$�-��D�v��-*�x�N��{�j�jQ�r2�:���k����=��,� �e�L�2>��øݪN|7�_�����ȍ)߸�܁��F����r�{�|$�;�q�JUq�l��6@�jz@�_�L	��^���{u#ۥ�o3��15~��y��e{��q�Ό��:�9�����G�,�f;K�_�9O�F�D���HE�p����z�����gz���L{��i�~�6������{����q`m�?�U������|KG����-#B�z�9��R�F���Q�wB��z�n+N��9k�-%ܺ��c\�@�>��hT�����ϡ��/{�Ȭ�R�Q���W�M���8�0���h����͛�� z!���|�F���	�]q�5l�nΓ�[��}�+��Jz�ǸD�p�x��qU\o��#ʎ����:��,�O'Ҥ�L�Gn&鎸���27^ׇg�����#�o���j��=��Ɍ~�	�X�G��.�cĻ='ȫ�n������2|:M�ߣ^`U�<�N�_k@ϒ�:��������Bzo�jǘ��F���ܗ�nv�zs��J�X�Ge�@�"n�_�����6�wO�F�Py��Wi�����|̔(ʔʥGnx�V:39J��Àl�]@:5t����J�=fv\��|�ʇ��"�vw{�,�	��k7�);7"�z�z�f�%0�b���ƀ�o�[�
8�_�g[�ñ�7ڨڧW_��o��}�?W7�� Lr�_�9�퓾TG?{n���ޓ�8G�&��z-r�h�]�����'��>�w�U������`
�����{�̣��p8׻:�g�A������b�4�G�I���&P�o蝖2�+n��\��7ӑ-W�?O����H�nZ"f�EL�Y�����EG�(%r��Af�튤=Q�Z]�L�/�t���X���3���q���}��r�˨���m{Na��^���em��"��dGE��Sb�X����5�^��Ԛ��sw�S�JN{FyW]�f�י���>�����p���G�c����${����ώ���DӶ}��J6O���q��g��>�z�o��:���î]��6F��m�_i�o��{[�>�-�&����7�2�!��F�y��3�l�{���:�h�~�_��\��|�)��F��j�+Ɗ������M
-�vZ>��Tr5���&�׭#��%��z$i�(�(/�c�r�F�������3�. l��,:��P�����ә���G������W�Ч�k�Pbۍ��op!侱nP�6�M�%c�ՐX�����Vi̎�ir�,tP�`�ե��e�l@�	:��ak�c�d:�Q��П]�`�v=�oi<[���̝��@S��(��K��Aq�ݺ4����av�{�/��4'rCz�c��9ߕ6�^���>�r���K��hA�93�t��s�:�Ët�D��>6���a8Ŧ}�}�G_ޞ�LYy^��D�p~�d��(��-50�~��0*����"=���W�0��G��n�N�o�~8|�yIf��D]�EB�� ng��r��y�U\�ϔz��M�a���]&��O�ڿ��ȇ���@��yv<3�8h�8<h\�]`t�o�=ڨ���L�����7��6}�C�eE����/���<r;����%o�:5�p����F��Tῡ)(�̰��N�q���/*��ic�3�X���lzz�^��z�J�g���������ӽ��T�H���|P͝�2�kJ���6���L�V���P���Mf��Uߐ�,`�g��sޭ��j��^���`��rZ�}��[�,�=q�I�����):{�,������~V$�F(�^�"�u��+�֎��{mr��(���/	�_���u~I ����]Ǣt��x^L�s;S	��vcs�~��>�z��o���Nj����h�]}~�J�w����݁LBX�h�͐y�rR�y]|���=
wYf�f��3I�Sx��q�2�sP��HK�Z����j��ۏhe��jW����U�I�bse��4��w�>�(p�Ͳ�}�m5I����뻶��d24�s+ aM�y�X��AP�R�S��F5�!�Df/wtr�O��R8=�Ru�'���Je�>��㊟�E�uz��<S/�}���lOL�R厺�[���%%��Q�@<�}��7~�S.�{V%��<�Sg�Xp�[Q7;��#�^�����2^E��z���
r�/ #��+�@2�6X�8������'��!�{3���|+���{�6
�i���a�{3�F˓�fE��10ݪ���V�,�tN�����^���tįUs(d{�H��1��ndH����@h�LL/{���x�V�V����vm�%-�>ٖ�{~����I�R���[L�k�w����6�ܯL��ǆV���=���/� =5��11K�h����B5M���p�yU���΀�fl �������mm���3ve��ٛu��D*�Vɯ��>�x�4s�Bc+��ٚXa;���Uӛ�����%��!��֒ǋ�����
�3kC������ɥ�ǵ�X�/A��RW��{"@��6|�޹���M�~��i�����v�?\f֏^N����MV��Wxo�W�^�2�`+��s���I)�o�Y҂7�J9;�)��1Q߻Be�x�Z[�닔�F(l�J�����uֶ^Qc���k��/(�V3�*�P���]���XQ�i��xn�ɼ�g��{����+%����u��쥺�kYE<�&�HI}�u��U��~o���Gz�5�ʱV��:b��{M�h���C�{^�$��Lmh�4�3�,z<���������*��#��|J^�q[hP����N���y@�u���n�ӥ��;>�څb��u������޿-�w�Npj���5���3QT[P���9�^!�|v�X��#��+�w�U>������wq�ׯ�r=���Y�G��Y��֔�c���}���!���͑%���`_z��d�s������z�y��k^]��y󎖢����S�R;��mڨێj�+6@�j'���0&����A���)�a�o���Җ8|���zC�+�C���q�=]�=���W�PRY�p\�����z�5R�_� ���r�j��F=��8=���d*y��B�{��ȏ!+�dF�����ǇB��y ���ly�����~��{�\���nLx��p�#�ϡ��U6ld:�6|���X)嫡������r����\��7���o��x�Z��{A-܈F����w~������ى����#�@T��;b}D�uڵ\y�]�V��9qv*e��O�Dw��^Жt9�u㛝ٗa4�V�H�fǛ�X\¯��������B��5�g��ݮިr�n�ܭ�W����h���5hH��Y����˳��}�㡨7�a�r9)�0�#�,�dϩI�aq��,z��DLS�ӹ �Ӑ�^�����WBY
� �&|���˻�O�L�5&�T{�d���Y�3����I�V����Hsyut��,�|�%2�r�Q��^71p��yND����K��+NI�=qu_�[���ə���twj�K�6�/up3}Hz�:�|/��쌏s��}�L-�2[�.�)i�¶^����(������;|�t¸ͯq��<�׶���~�E���P�]P��y���32�MFJQ���l�O�+�3�:vaY߱�G�fp���Fu[ Z�w�|1�Tw��x��9���2�-�z�I��c���偆j�?Z���֖=����x��|5k���cs�ޕ�+N�ο�~΂����{jA��ˍi�q����=uHz�&��'}1Ӯ�sx���p�U�V^��r��� }����Y�k��k����(�YD�n"\�=uL	���b�o�A �H��Fkʻ3ڽ�y5>���yN�<�3�t{ޟq���6�3}��#be�O�SF�8x �x�*����������V�͈.։��6-=��;ǋ9�}թ��}�A\��zn��a]��w�j�v��ڳ��P<�L�y�*����RP&T������H��lK�2l���{W��c^�V�r�#6����?%ueeZ�F<��ޕ��|�.6���{��K�����[�^J��S��.�8�k�i-���w+�:}�5��R&�
�{��
5��uǱ�Sg#�'û"7����(TU��)��y��O�^L�\ ���%>�M
��H�h�s�mdK7�TuïZG��h�~���:���%i�7�z�tzg�\ s��V��>G 0���~7���� z�2R����Ƿ�&r��+��zgx�sޑ�߷.]u%��4�{NL�;%��Y�;�W]�UF��B���g��5�g�ٕ^����?L��pq�fAy>����ۛ�}\m�R���ū\���>��+�b3��\����y��J�8���"�{Ɛ,p=r%\�=ػ��ȿD�BW��a��c��Z}���xhN��{�޻,省�e��ຽ����,�jm4��r�&G��D��0~�~����sra�O���/�������y���E�+7ެ2}"�X�{�F+5�w��lzg��;#�*p�s��\ς�s��x�z&)dH��9��'xJNG��J�GJ8�u��iZ6S֊s�j՘:�9TV�����lģv���-���� ��2���.Աq��S�=X���1��G�hml�,��[s�R�m.��J|�Z��q#ՃxS��<3�A+.�<�����3a�)��:.�=|L���_�6\��� ?��ͮ��t��{	��'i����B���7q���pr���_C5=���@mg���s��2��[!H���#e�Ѹ=G�*��;}s���}}~;���nwe�C�͌%���@k�~����$\g�^G�V���z����Z�\f	H�*��GG�)�NǦ�ж�W�~�����]1q�;�쭻��:U�1��~�������yU���Tͧ�Ed���}3ݎ��?zD���K	I��޸w(*Z��K��q�{NF�S)>�꩘�Ӳ�>�}��ױ��z6�[r�=��	Tg��M�X���L��{V%����j�tx��B~��=�������1����Μ��� ���+��] �D��,y��|8k�h� ^��0�B�϶�S�������}#M{-�;��׉b�����Ңj��;&�9l�z����f��J�3�|�+Bn�^,lG��ϧ>ٜ��wLz�����q�q� u�ԭV���K}�B�&'��ONA-�&|�$x`���s������A��f�6�m��j�V���ն�m�Vڵ��m[j���um�[o���V���mZ��Vڵ��歵km�}[j���j�V���m�[nն�m��[j���*�V���Vڵ��J�խ����V���Vڵ��-[j���Vڵ����
�2�ɮ�`).�������>���������T�R�HB����*TR���J"�U��<��J�BIJT�$�PI ��J��(���"Q%��**��J"�P�UJ��R�AHD�*�F�ê�)�AX� e�F�(�)i�i��J�S@#�8bPl%C�3`  �  ;   @c��s����1�CB��-�J��l�j�Ph4U����*���dmak��KM\�#Te	h+֋b�3bQ%�C *����4S�)%d4� -�kT 6�V�[t�fh��iF!�+S` ٴ$Х1U�l��J� -G@Y`�hԃ@�@5�����ѥhZ�4Ҁ*Q���m�::k����Q�l
Ҧ�Ӡ*�4�4+�@�f� N .:Ql�62Jd�	Jٕ�k$�[6�ւ&���E' 7.Ԗ����*��XZ%5Z�[��IZ*�[2I�¥	C��6�I%�h�֠���T՘����P � "`�%R       )�IJ��#	�  	�0�Q&Bd C)�M���<���6�
m���@�)d#L �4�@�2��L� �LL&4��&�&"��Ѧ���#C 24�&L 4ρ��n����m��/8R����P�
/��4@]��"7 ����Z)� ����>���������A�*�,�?9UE��@$#%�*�h]-�r�K�����ފ��|���4���0����i���)D_����q�_���x~�:չ�.3�w�l5�/�f��kk)�.�FhE���I1�,�N��8�'rĩj�v��U�o灡w�����ĉ���EXv�SX(4fVS�j�ӄ�H;Yj����.�F�H))ͣ+#����i2�f=�7��	�����xJ�Y�Y��2�5/*��5�,ZrMb��s�F;u��i�ˢܚ彄K��6���f0����yݨ���^�V�5KYL(JǢ�=�opM��ԫr'�,��Yx�%�s�#��%*���Q4j͋-�b�ʡ�Ci:&�\̭��w�KwFBv�7���mn��r	����vuܴ�6m����nG����Ï]�Ѻ��C-G+ie�=L�(nY�L�d���;�)�{�^��*��8,�T2;�23�[ʘp@��m�z)�PI�^�U0��g+vS�ݨB�aPbղ�q���K2b5��j�>z��M
�A8�rۗ[��M�����Q�	�Э;��&�thG���pƉ
�h��$�ZDww�
m���W�xr^��
X���V�<��p2��/ohMzIK:*�m�GH��iWr���R+��sK�@�Ǝ�58���6L	�r�6��D������ �Q�
�tŪh�tGzmɪ��)(RIY�&��v�pn�jT��Vk�]��}29>c���;[kl��-ʑ�"r�!oET7�@-�H֝�H�^7v����%��V�*'/n$h�d��{hM�M����${��l�72J!C+$J�{[t�B�.����7JGF-fE���q	[�����2��60�]��؋�?V���YtŠ
� ;+\XHӧ+ڏuJ�g^�R�l��f�Ʈ��zY�X)������(2�!�Nh��Ɔ�tTv�������e�X��z�]A����t[�Y+5�;S�OW�i����\���u�VTө�K*���3C(]��z0��ɹ�\6��:��E�]mȮ�RC*
�in��(��XTgB�i�����`0Ǩ]�MV���g7�k^ȃ#Vb�:e$pV�St��ԃ5;Zb�b^JD�V٦,�LwBP��	�*l��-b���X�z5n;p̺w��Y�T��ckc5BM5�]�\R�5�X0-ʢ�cݓrK���S5�p[{��R�2���˚X�����%�a�j#CN|
��eW-KS�4꡻�7c�h���Q�2ͺ7��]Jyn�JҶ��!zm�����#r,)i��f��H�tJ�cHYQB,���Y�lfj��
�o�ȉ���K
���)m=�����)\��#ɗy��H �.�̂�8K���:uh-aP���r�6�u���"�(��D�h$�&�0=P�b�#��&�^j�X�Ĳe�V��E��pCrݢnJ�+۫+��T
rE�/0mϲ�*rȠ�f2M���m�m�V�3,�f�16����ކ��M��̖@�qR5�,�M��4ӷ��T��36��HUGq=U��<�b��뉍v*� 'w{M�	��a� [�j�kfɱ�;[Z�h�x�����Y"��Ij�&��,nn7�k-
�kBW��Pl����$T�i֨}�r�޽e����m�Q���0f7u�\(�~�3!�RLn���rS�xK9��6��v.�7�cUl�����1Vƨ�h߁Q�$�gZsnz�ߔ����ն��;q�,�`�4d9x*7{�� ��$B�:wA��܃Hڑ�#�{��s"�IǐI�Z��wT��KD�*���2�4omU[���Ɖubl{�b�㡸�B��ݣ�w�J䫷�b�4^�@�ڃ`,���`ڙ.)�wx��j�O�᧓�B�6�r��lM.ء��Ѕ+�+`u�h�NDB�#�)�w��N]Du8sr��)�k)��J<
1d��זֻ�卛E���[*���0��)�����2��IHKrdV��5�6��h�4��z��A�Aj�W3lMcx ۽ӣj些f��<[��r�ő�����hըXʴխ����;q2ȩq=�2��6�7)�)-����@�m�4dF�xl��4�Làݪ�U,��ˆ���oZ��{�{�6��TCe踖�u��ɓ3cb�)�)��E������gԾ����{�����N��zsh���ƃ$�O�wr��j*OH�����.b�c���0""��BΝ&�U�bF �kC"O�5�lml�M�Y*Pup�<Æ=;�eQr*,�@Z��[hݣ����ar[:��\�H��b��{A@�Nkb��;�jw{����0�nf�Ifi�
�SgQ��)E�[-FD6��H�f˙V��RMN-�r�aJX�NF�h=4t]�^��8Ci�6ꦘv�bݕO%Ȳ�Owd`�#)QRcr�Ӈ�
�tu�hiV�3)��#�*۬(�"�a�����*K��fP�Бe�J�:,��`��Ҷ�E	ѭ��FT��Yf�<���WgQ��k*�G��Fj{QXb�rkB�ܒS?�ye�ٽ���OI�X�S��s0�+M U$�Kl��^Ⲷ���O2���tN!+[f"�<oW�A���ܥT�[�#�{eD�6#�r��6f4�U�7�u�Gn��2�@���&GfU��Y��(����-Y��c���AWzf;ܭ�0�)I�ª�e��'埥���G&������ś��ݝJ���2����M�q0�Vw*������]��N��l����#��I��m+֮a�CCX�����Yb���W�*Ie�� ��F�����4m��m#J��4�47l�dˀ�Q$뭧�E÷q�r���c�U6Am���^J��EJ-�Tw.��	�c9+4�����*n�kM踞J�����)����A66l�:\ٹ���kx�hdT�x^bwtf����*��H6���[�xcs�tX�������)b��[Z[X[�7r`j<m�B�&�i#ZȒ�I�u��ɬ;:��g- �aQ��0����6i�X�w,��iVĶ�͗��eԂ�Sd�ya6�r�pY��x�Kۣzd�&�����T�lmcP�V�c�Y�%+Ťl�Kca����;bĘF[��m/�B�b��V*U�GyE9[�"���Td�%dЩ��r���[��8�+�a���D�`S�Rw+��u*�b3B��t��v���K�f��)��#����^s/��7O<�b�ѮC�!$�)��i�8�C,@�&��o����MZ�������<�-��F$�I!���)$�I$�I$�I$�I$�J��Ŧ���H̢qQ5R@ȥ�C���I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�K�	$�I��I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�G(�h"Y�f�M��zg��QQk3�`�!l�A����"F���3�����sS�*�V�!�4R��3Y�J�pHZg��'I]匫̍�`��r�-��{���+f�ޫ�^�m�o��2���v�U�p�қS����\f��bv˵O;%�g��3Uuq��T䗔�3's-��J�3˳�q����"���I�Ʉ�D�y�g6��5�lQ���� Ψu�����ms玷P(�ƻV��:��t�QY��!�玮��3�P�M����s�aߡ��e0�����H(��:�[?Y��$�di��f]��<��ؘ� �eT�h�8V*��*=�49et��!��մ�4�!Vsm;��Kă�0�`����.�\�K�������8'�0��9Z:�:X�z�Y���u��4�ݔ-6z�īX&�Ňim�'uB���@�'�Vi�M�G_"�d�����ݭ�:�jet[����iHv���Yϊ�
A#2����un����m�iUh]4+s3�8�nEH0�����YU����{)oT��9�;J�E%,	�
��U��w���T���[b�5e�z����s�ksr�z��Ϊ#�%�5�zK�f`[j�u�=�
K�����`����� ���]���l�u����НӮ�M���Ъ:�E������oF)����|hu2m̨*�б�_31S�Qk�r��c5{��;YE�
`�י�ͩOd�NT+���=��Yx7.�/�L�ݮ�����/��:u)���&UY���M��ߺ���TL�B���2�Me���>6�M�[+c�/K���[�n�.�f�d��z�V���3p̻x�ޔ�\tzm�����Z�e^t೭qU�%�y���Y�u�]��MXΡN=�x�ఔ���>g	��+�ƜD[�_Klm5me+L����gub��x�����E&΃t��v+��{w��T���{z��)��RV.wZ����5�;~/��OvS^��42�;�9�7���z�d�"��;(���ir�c:�"o�C�b��٠���<}���}�Iz\+;�5d ˼�\�Z��4��t�K���0�0�r颞08p�};h���9�A7k��jg�'Q�DK�ջHK��+!��<�v��ȡYE&���O9]�E�穣j�4��m�GK�E^�۶A�ҭ�%%	�$��+��U)�'6Z��;���ՙz�D��Uq��ҫ�(�����5��k^mE��[S��"O�8���o�_e
�%�r��g�� �M�d��î<�F���۹���'3-��Z[�n�������X/���c�x�Ջ��ѷ�WTw|�t�K ��/��;��H�ʼ-�aɗUȲ�!1Q�Ggz���o���֍���iX�ؓ����5(�WD�&�(��r�|��u�(�.��Ha��Y���7�={-q���VV�YzI�&�Ϊ��E�LBf���aeo]_Qwfjv4�� J���w��$�M̦o��]�wݻ�Q�t�*�+���诏@uuc�*6�,�ڸ�	�9W["�!��'=���L��d�K2�fL1Ӎ��!܃��[���%�K{Y�����ԉ�W�k��u��&04I���C��4�Ȼ�Y�ҳ��%,o3X-[��9�`�]R76��xi��Z�"����8���1�ƻ���jd��6wRQ��)��ZՕ��h�:���μ��FKr������Ce_L������9�ta���=hj�%^�C	4*o>��sDH4��lm2���������6ã�{C�8#f�$F+ȧM�xr��0�awyA,��GqQΡ9Ua��F��<�1R@q�,>',;��f�a�cD*^X��9�u�7Y|OL��4��е5��p�ew��{���J��{3e�ɮ�o�L����(2�!\%R���[t1��N�Nr���hꃦ�lۻ�Ug���wv�̵�u;��X-���q:Μ��e)\N�^%��f��,��i����ǦXwL��,.lG� +2BT��X4��4��q��,�LG�[�a��ͦʍ�̧�3��u�p��Z:oY�ΗU�E�(鿮��֦T��E��6�^�[:;��x�}a+�7��<;m�4R���]+S�K޻lu�x��c��Ѩ�b��\"�A��V�=O�LTm���t��uױ�i�N��ե�4���D�Ma	nV����JP�iz��obv6�&$-E�� }���ot��R���*�'�zֲ���Ⱥ�T����ۼ�Xa�y����MJ�e�nV	z��:��P�;n�.��P��Y��R��5�zE=�]�+.���Ii#9�ۻ�^\��$��ϑ�(V�#M_�ju&�ww'yX�=u�ګ�3�!5��N���m��N���O��S'&Qg�A��1re�sz�5��m�'yi���,5Z���]�_m�ε[Xx�>�k/��P��
ȩUMj\�t07��E&���Y�y�e۳�{�F�s����i+�GVngU�`�՘&Ar��H!ƴ����rm] �}�u���0�rmn�o5lmJ=����L�E�snL���M˱
����+�V��s��l��W,�7�f!+Wt#A�YY�̵�%����3���֡������ �� r�;��k��FsR��Ww1�nZQ2��U��<}�b�p���Ѡ��n��p@�¼5wo�}	Pgf<��A{�EJO7vr4y�֥��'nJwɫ�sƟ�)sjhl���e�m�^�Q����RJc�"��1��f�X2��g2�֘��qC��s`�J�upp���-^v[Ӂ+��j�)�	Fk��I��J�����#����5)�6�O[{�Eh��|~6u;S�����	�J�on��4��&��9���Q&�,�o&��Oy��ܜ���Ot�NZbj�C��P���L��e�W+%�o��U}�@�=���v�o�<�pv�W�m)�`jjN�e2�I'wT�Jm���I$��IM����$��RI)�Ҡ�N�'�y���:K���t��$��RI(f��rg���s�9-0����k}��W��Wu�\t�	����]݆$�L����e��A^9�mtT�Ncw|;�z)9'��m����:s�VGStխ�k�����HN<]N�u%;�wF�����q���I$�I$�I$�I,zl��s��RN�e� Qc��j����jQ7��B�  ��=8�0�����U�"ySCd���F�ur�Ae�n���R��W9�ͭv�*�\%��un�*��|e���Q��F�u��-�389g+�o,�Zn�H���o1�;,Sև[�뙶l�(&���E���aR<�&��e1�*c�]ۙǵ#%�xʫ�!�o	�h-b�w�4vgu���M5�(��l���edU��C�n�^8>��Rx���-m�O��I���ˊg�����0��F�!%��;�a��V�O/���e}Tޖ9e^��&$7����}<�*Է�I��ј"���_Xl9�R+)U�t�����"��
K9�m��n�#����o�r:DΦ��I\���%a(pJ�f�L�Ȼ�4:��}M�v~��Yh����W=}��Ώǻ�=�E� �0�X��[�D�ʌɨP��Q0��z�*�|�>�k�lL�T������}/�-�-�Q���/�u�J��{���a��R���#+����Y�r8���n��mA�����jT��(v-�`��#��ܖ4��nfH�P�e=��P�R�n��>�oXb�.^��ZnYm]:Golݔ��3��l�r��d�z��c�/b���7�S�{{5�(˩�\?v M㹻x��,T���8����}n��v��7�ѕ]/�W1�YUg-6��˽a�/.�s�sN�}�_Zy�����";g ܈�'I�͗�f����B5���v�#Y��k��(�4�Ve;쬆泇��7��\u�KgE���K��tp�ي[��P��|�j�q����^a���9�{�����ِ���@�|Y��<r��졝ɹ�"��9��n�6��N���,t�n��䆯�w	�����=��d�Y�HY0E�eY��ܠ�S�q�0�!n^�ŵV�S�����DQ%t���r��pՃ&n�T�r�7�8���
Au�!n�U�أS:݌WY��N�y�A"��-:v��!\��p罏E�]L���|�,]q�4Բ
R����+2�x���8�X��ehɲ�J���	��˽�p�O����}�(�٩u�i��0�L�F�[µpY`�a�ר{5o�v%U �3�F�9��Hb���#.�t������6��K�AX��ꝋ@�!�{�'a؆�v����U�������Z��T�s��������wJ-Q�t=:n����6J
R���o76�����<�k6�<��늝j���C� ƽL���5�--�Pf��g�R��]#�Yj��%���+0<��qf��eK|nc	�su+5�W�9�js2��ؼЪݪ�����7���AlB֊�SJeF�bV$˷R��%ob����x��.��'qؚS�<Y���3��f��μſ]�ݩFs�R�:��K��f�y�]yW�������)9�&�.�mg��7������0����8��*��s�Q�ܶ)յ�Nj�%C2:T�%X�\r�]2�"n���[�Q#%�*ԧb�otZ�Z�~C<x�ܨ�o�9��}y�C0^�i�i��ę��v���c�v��ED�"����e(u�%�#��_ss&]]r[�vir�z/�^vi�\&Qq��2�g�ܢ)�:�O�z��]nގ ������S��6�������A�9J��io9V!�a�X1��V�Mu�d�F��u�E��N�9����h%�*��K\I����<"Y�pՎ��no=S��-4mV��h�z��Z͵��T�ʹ#Y���2�#�ޚ��銞>�gF��e^[U���A[�P������ܝRT ���M2e��z��):ŧX� 78��YkB�1w3}�a�CoK���it8���l����h��=�6�| X�T�ʾ緹8$����]�(��^����Rv�g�f5Ie��c�����`P᭬W2�>����EX4_����C
�Qhs4%��/	�7������ꎇz��<#3"����ʓF��*�W�"�K�RÆ�kh�ZU�Ac5*�B���.�E�kord18P��P���QR-Lk�-[ɴ�f4PH�I�=��q�J�_E%��1M;�:Q�:�VղRF�JC7z�4&NʄT&��^���q��"x����*6d�St΋6l;�5�"v���Gl��g7n�[���m��E��oz�洞v�vR�`ٛʐ�n3�c�J��r2�l��2�4���,"T��Vǘ���B���M�s�yIڧf�]�3C�oU!l<�(rI�e�^E1���ͻ�0e{iЂ�r�� �Ӎϖ�5�Ӫ�i��
�q;8�iT:3�u�U�H7�;n؋'!K��v�9�;��X�<|Z.����׸�M�ڤ橺ꖘ�@	x�`�tkqq�;�%a��*�qH��7]�gH�T�}[{���)��X��֨hڿ���G8�8�e���s���i�Y���(�y��~Ǥ���Q��yn��0��{L�juŶ)or��'0�V5���I��+z)��e�r��o{l7�t�F��g���CL�#���u�Q��e�[�Ih6W�MMhZ��nb1�-kU;�����t������|������n١:+q�zX���uy��]��8a�S�,5��\�1�nN�4	������DXe���k{�w1�e�W'܃׉��gq�eЪ�BAն����[�����z(78mX6���d�jM�*�.-��;ކ��P��2����Ю��F\��W¤9j.S�.�쉃�^��m��, 뻼�.�t���3'T������܍P�r�)��)7U��$a�+3W�q�4��|��Ĳz�Q^�j�Cn�o`��I���M�R�k���.��W���F·!SbzK�cIY��핤���^�Yۦ�T���g˼����,�<��Ѻ�YW�ON���]̛��Y;y:)hX;op<�x�Wkn,��%)�����ﶛQ;l�z��v�Q͉p��b��]oP���S˽#.m�4r�9J������p�P\*��0N�!���6i �GXs[��ugo뵶/�P�N�l�d�j�;Ȍ��줞W�K�UûZfh�\,�p;b�V��ʔ�f���p5v�G{�l�����z�f�]"�M2zk=��(^���-��|n*��nlI�����ǟ1JX7�f�s�f%��2-}���hF�i��˽�xu����R�c��3��ì�Z��'�I!	E����1 ���a�I�F<����������{ޤ�I$�I+��ʾݛ��ɭS&��
��Z{f�v2�C�p��Z�e���X�4��*֌�o2�e���N
�.wq뵪g7p_.:��n:�Z7�s�Y�wmfhC�e��[G!2��wWf���:q��B\cl����_
�aF&]M�O�vu�{X�k���x�һ�l�*�&'\{R�/ Ӈ�����ڞ�t���z�u���Ť���PT*��܋^�bK�m�j�g\����c_p�/��z��=�6�6�]��[A��\Xbʼ�V����:��9K��r�;a�����{Ka���%^�V,hk�I���f�R�7Q�Q�`�c��kI��s�i�qb�L���B�!T�gww�1(�qX��s�MI%Գ�����u�gk��w��~w��Y�h��@ 
-���6�)"�E8�0X) ,X�Y|��2Ȥd�aFV�YY��Ȱ8�a�J�*AB�Xm�X�AD�8²}��V�`�یC��U�,��I�J�8--��"��"�1jAeaR��f(T�R�R�����ޑ<U�	S�3��N�����j
���{��S����>'�VQ8v�w��3hu�>�Z�,�Y�k�8_�y�
�A�ΣN/�=��1�p�,�F���WOr��U�qꋝ�@i/2�\��{�玠�
��E��;�� v�D������Zc2)��'$"�]�~�LT�^�����B��x��}j@f/���5�y5�B��#;���?I���x���-�Z���t�?�){]����(�av�.�LR��v�X����5[&�9�ϟ]�\�i��Q�w`2���M}.��Q�_L�K�XH�P�t���3�6��v���uO;) .���5�D�v*թ��P�{����Bf8+���C�l�zs��7���+�ӂ3����C�~ͳD��z�TSP�;��imz�U�G~f��īq{#�dN��br��=���^"1�[�d@��"��g��i����l�y��!�CK���tcE��Z�ɜ�=�8�fwEC�R��<v_��	�7�9q�2�Q���~�ӳ�J��h{0�����Is3!�e����9,�d�Oso���Μmu�*�Ëdj��U%^rǚ6���y�1�ݏ4�*D4�d��$�ib�X�$����:��|�9gm*G�@U�*oɡcs���O�(s�e��֮�*g&%ۡ���)6�Ȧ�Ϋ�I,���_3}��dŬ�b֔��u���p��}��f�5��2�2���I�Wi=�P�Z�Ob=u�ć�[�U�� Gkܝ�n/��Ԇ�[\{a^�	��4�sc�P���v.,�BN/�<U��7"��ϧ���KNG������י1�"�J�2�gB���q�u��i��X�n������y�Ȩ��D���`��瘨�ee�y��L�j;����
��>�7{@�����a<��gA� ��6h�����ս6�[�·^·�n�+�.�1�/g"6�t^���*S��-�kh[�A洷{!�Wc��6��,	�����]�։.�섮�9V�Q��*{"�T##���Y��׸C��a'+����{SU��]ػ�|K9v���"�h�)�}����YE�%��3/z���7�?pp�sA�����ٸ{�<sUc�&u���ߟ���Зx����:�@�/�������E��΋��nf��]��#��
�(ɞ�	#K�Gwl�v2+��G��u�5+���V:�P��M2��\���!����H�X¸=�e��zN�i�҂EK��lGB�t�NR�{�ri(nuX����O[���L:�m�3w�{���+��gwkn$��÷�};�n%��U��4���9�qNn�3N�������������Y"39l�@8@]	�-gA���/j-��ɻ�<zW�NJ1�9�f�j�;���
�w��j�G�&qL}�{�s�꺥X{L���#Lְ��[=��˵^���������R\%���,V ��`�]X;nF�wD���w���+ZE
�����7�l��<��A^T�Ŵ�i��J�����)7�]��>����-Vpx�A;�哵�籩5[/1�w�`
���+���ث��.��Ĉ�a;�ƨ��&�vE
{�J�:�v6V��EM��MY&h������-�Gt۱�s7�:�=.�x��6H���:<A�.��m��u�xrxz���ur���;=y�),�|"X��Tҷs8/=Q�''��b�.�����3>�g�FM\l�/�b�H@W�nfx����Q���dv���ы�o)\�=!m���T�8�7�!�S/AE(��*��5��;T��|�0r�,D�7Na����]`�ǱP�m�A���Y��ge;�'ͥ|ej"�ۦ�k�����BK������k�gh��zL�:p���С�v�C�n��U���hE�&�kI���Բ.����j����;�9�W�h}�:�E�u��ȷ�M�]��fk9�Zp7�y��H�����%��5��6D��wG�;:0�!��B�5�L������|��ȗ7{�Fm��9fPo���E���n+3�%��ӌ7���il%=�(،�x6���ީ*�od�AV�z�y_���S}q�]y���;;�H4��qf!�S�\��_I2����
	�|frln�b�kW�n\��w&��y�c�Ӝ��{�8lOP{Ӭ��`��E��Ld,�.���x�sJ�⋅1�>j��Z��C4�.��\k���]�`h3�uw5T�+��Y�(�����v\�n[Z�K�
���5X@�5y��wL�yU��	quP����+� ��]{/���C�S(2®�6�IL>-�h���cg�T�(�O�������";��hɇU!�]�M ��c��y�ף� ��]������򲐀c���5S�l���:b݃.�a�x��V��W=x�al����R2��l_o,�徂b��y���z2F�c
Iw��-���]^�7P��QN��.|,�f��ͨz�-�0{3}y��r�{u�[�ƁN�qhM�`���u�ik��}�{w18��)�1�����р}�Ċ����jôd�(X���ˉ�0�&|���t�E�,=�u���D�u�QOt��R1��oB�X�<���Em���p�wa������<���)���3�c�}�9��j{�>Y��\��"C7L�R�(����ty�`C��<�|]u�C�]Q��\��|Q��I�J����W�+]�û���T��"6ء ��*��SZ[�Wf���r����4�z�f�#�,X��x[�]��0��D�W4�mح�,eY��C/t�Ѣ$������*'w�� �Έ�E�I;ow��k~���������:�>�;4ǳ�.�[�)a�ˋ\��K�:�F��--�9N��H0���'s)�vp7ت��d|���:Ϩ�o�uV��VM�[Ԧ�ՙ p�K��ee�U)�پ��E����b0z(\ـ�<jM�$fgs?�U�WR���C�{�����0�����RI$�I$��9
/#2�lR?��VUώE��	8��|2Q��;4X��)��������ʏ	�^�x�.��koln[��v��!8��1:'.+���ƎE�b+��f��dB1�j<t��-]��2َ
�_/�a��v-�L%�6�ePx��Q�Ld��d�~Pdx�eb���y���r�GB�rR���e} �H����"@���������-“k)�pݰ̵V`��wwhT��#���j���Q�wS �F�b�w�Z6�v�!6�*�ڧy��)�V��T�F��,�l���ז;�7[�	29�O�� �U���������V�V�Lj�0̥�#q�J��k%aXUER(V�e��z��X���S6QDJ����[h��0�V|��LYu��|��,�W,
�p�a���őC�si1q��'S
�)��PX��(��UT�\5dX�������cY�a��ԬP��EH�k�gS|���
��
��Py�C9��)��FK���&Y�q�+ٝ��]Ah6/�-�S��j����컝�p�P�O05��x�E�ɺ34�.����M���j9��E���G���f��ϸu��q[���N�햾[�~�/��F�!��u3N�>�Sy���o�F�ߚ:~���!Y�_A�!m���(5���(�d��,�VOݑ_O��F�͌����������c�G�S����w+u�
0�����Ϻ���7�;±ۻu߿�3��dt�?��H��ٰ�{�>Rf[mTd��G�2R���Z#���mܟ��u�d����X&
�۽�[�7~�Nx�J�{{�}���aػh�w���X����A�d���:/����>�1Y�dϪ��k!���\�?�C3.�~�wN^�E�1�\�%��㝙`��W>=�������[]ѳy�B��[#��^J��N/�@��ݤ�Y׫���Q� �ō-a�w�h�����U��QS�沢�>�m�����כ�ηM�H���?I�9���58wO}�����폪��Bn3�>N�F&������NEDZ��v�A���=��&��A���V�o֌R��;��I��0�U��j)�,���Eb���ޙ0T�v���7#Doih��S�L�#���f&���p\}�N���g�>"�KB�6z[��Q��r��ۗ���V8+�:��b��7��Tq��;h�����o�f&����lV��'ڦ=�h��{ۆW)��P�JsjU�X� e��m�|D�9m�GUGD��N�f���z�����<���\�����a�j�]Z��
�Qz]��6]�4(�����c�&3�oӱ�;FW��Z�~������4���ڵ9� M��z�]!�ړ�2�� �uj�.������O��L�=�㫾�����Ԙ��Q`Uc�[��m"�`�����1ױg^VRin:��REߌ��=k ���o�>���I��o�����q��/�yk�:[Ot�f��Tx��A����8<���J��t�
04�Ē`���!��>@5�xo�G|�w9�w��|���z�
`��E:�u��'Y���u�q`Ou�sT�K�,�uʧo�׋�C��I�CĚC	Ї��):�<�����̠u�C������皴������o��p���H���̡��ROP:甑I�m��ì�!�Y�퀰6�볝�Ҹ�aR�����O���r*0R2��Y��<ۤ{ ��Ү���8�NS]&w*]�:�캤���(%�#ލ�D{�>��k\�����a	�� �d�)L13�m	�vH��e'X!&�VIY�l:�=��Ǻ�]g�y���=��N���
z��	:�0��L���@��bH}�O�d����&=fK�<;����9a�a>�4�m�{I��!
��Cha��d��C��M{I�������9��;}&P>dS�(C�� e=�:�`ݒq�0��ɦI��!Xi$��N2N$��y�~��y�W�C��$X�u�����6ϙϨO>00��d$����>{w��3�!��~̋$ۡ�����I�g�$1�P�d�@�=d1�@�}I� �<<߿k�Hz�z�|�LY'��3�$�'(z��CHq �2�=t�2Hx��]{|�u�o���&���'BI>@����0H`��!����'��3��ԇO���_k�9������@��O�!��L��I�M��L�Hu�?XM�3�N0$�>��>�>��e�i�{I���:��B�4}d:��3�$6�Y&�0�N$��H����]������u�k;�u����6�V�ץ\�{b#(_t����+��/`� 4^'���vĆ����{��/�˟3�y���� &X������I�d4Ͱ.�C�C�'���u'Xf��:�d�x���3�iu�1���d��$;��d�Bz�|��4�eI�Xu���>Hu�VT!��滻��5�oN|谆;@4��\g6�g�O�&�
�5�>Ly��IS)����÷��~����q�ԛd��a� �=�2C12��i���E'ɿ,���s��Ϟc���z�d;��C�hI&�d�?09�$.>ć�d��d�O���7���9�;簆Ӭ���P�@�	�I��I*x�N3,$��^ٶI�5�$2w^������u�Ì�̟0�`^XO:�7a���:��2�q�C���'�|ɬo�oRC��8�z�&��Y$��x�0�����	Ϩ�m�(M���y�������o�Xu!� ,�`I�)!����E����x��	=M��@���	欓l�:c�Xq��_o�I�XL2���&���!���Cz�u �I�C��ChM��@�^�W��;���x�\ ��YpT�펂�-�K����ጝQ���Vio��`����kT�.�!d�!a���#6�G�����3{�k���p޼�_�6̲�ԁ�v�l���a�(���a��`8�M d�Ƞ�N ͇�S?o�/����Y�'�:��!甓�8�>�B�h2N$�I�i>jH=�������y�}�σHHs�u2��	�)�!�&�u!�ԁXsV@�0Ͱ�,�&4�ė���<�}�~��u�}�����	RI��l�$�:����`=d:�!��	�8ɞ��un�}����^s�Y:�z 0�l2q ���4��C��(d�n�F,�L�H`�|���1�3�|��	6�XOXI+&�����\��C�RN�&��+$>a��5����/w����¤�!� z��0�O�XI�b�uBm!�'�X
|��}}d��q�߻������Xi {<�dX`�!��$�'I�'�Ì���$,���C�>�=�5�����I����OX ��P�9Ad�ԁ������ha'���|߻����u��N�P��������v@Y~��"�q��]����w���78ɾg��g�o�ګ�}�~5-�N�fnțl�U�����3t�*��t�G%H�=$e�ÇBufT���ԿL��{ވ��#���=�����|�V�R#	�3���!�������760��Voe#ؚ:��Mf�)�y����1E�_��qG>_n���S
��E��HD�V�_���x��j�+l�O-qR�^�ƺ�Y^SU3��4&n�H+z�)3�"��< H}һ�����2��읔�G�r(�ne����vc��߽��w�d�<b�;܁� .jz(W��W�S�ڝ���O2�u)Ĕ�5,��;�^�7�PmU��f��B9����p�?0x�CF�}gG�:�a�E@��a�,|wׯ}�M� "��� ��s�s�^�����Ⱦ���O�Ԣr�-��"�p��p{��Lߴ�4�4bc�q%�"�ǃ$2H�ٺ�j�^�+�>B��7�64 2�bZ�DⱮ�*��)�A���f��r�w[��6/�1��nȝ^�4A�u�5�b�����؁PvY9��<��x/ٔ㓛���ެB)��o���`��an����y06�Fߛ��^��l���'a�è]י��oF_���¦����3�)4���w��ݿƸ�,]$>���s1�;Ow �rA����i#V��/����$�,!"�P RX@P �"�E�,H)�b�QAd殽��ן���u���y�ί���Za4P�Q�qy��'�{۽S2����/�/�p�"~T)q�7�q��ev�|x�C��1��
:6�W�ۆ�ƣt�u@�]��qλQ�[��TW�ʾ=��Ş����\�b�y\oQ�Ӫz�Dy���E˷ѢLRz�Ri�6�]��*,�PW�����y�����C���ԥ\��п��^h��]S?qC./�}d�Vr��gu�Z�P�B4���t�1��z2V೿N�Mm��D푨�:��X�t�N^�w\�u.����"%n�.ec1m�6�zj����p4�|�����="�eks.��R��wrn�a�EJ#��'|�����#�Ymt�;��������1��ً3*�۱�aQ���7��*��G��Ou:��ט&�4J�u��V��t���Y�M�v��J��0�rMe u��vv��nF_d�����j��oeh�:/��r�Q��ےv�NQ1��X](�e����BI8fnK�:��Hc��F�}Y�+�m�fQ
���P��2:uw̃�':��7��s�s��I$�I$���m�e����.�wyLU�h��aDТ�`�j�b���N-��,�͓Q�nK�r_�E���M^3U���c�6٥�3�2aN��f��M��M�c��J�yM��N�4Z��PY*�:b�8�+2�yi����1�$����.	RA�Չm˕l�Y�U�D2[!<�j;���M� Y�L�˱vU��6��	���P���c�o~W(4Bw>%�?�2л�r[���sʹ��&��{M�oQ!�m����b�i�:���)�iUӫMzM:�;��olb	'��B*�.��ܶ�ӫ�~����??Y�&�H((�|��a�Z�!qA����8��w�cV�����c�����A)
�&�J��L5Xa���5C*�"h�+��a�͘�"��fR(gW.|��ΤИfc�0�b���pf���1l�11\-<�&3e,aP�yi1���\��ݺ�T*�,)�Շ7�I�S	��.�҇�}_}��ю5ާ�6f�	�@�vD	����YՌ���o�����	^��'�P�&��}��V�6ձj��n��V����;��s����q����:BE�x�j�C��2�Z�0�4��N�a�V|��i��w&��a����ɝ���W?'�^(
T�FQU9\n]��n�3Y���A�x\M-R(�-���b�E�<x֥!��WS>UyK&�^W�[e��{��춨��{0^:z��ZYV�v ���v��gu����	m�֖��%0�%ZŸ{G-��8��ZԶ;�eD��p2��(Gg���G���Ԅ�GXbE��+Vb�Tn�}����"�)��'Ӡ������.�B��/�K]��X�W�:/�=Y�*�7�ɋ�`T�F��h���-��w�����8�p�=KS����;�V�-9W�[���|���O�\�O���&6�b,�.�4������Y=�@�Ѯ��L���o�s�m�aF��C�Ʊ�f�{�V|�Z�ʕw�2{
���cY��U��'�-�)hR��u��қ�Ou]��VJqZ�e�[B�7T�(K�S�?�z����{ގ���?D����W�Š��AJ��w"zǣ�ǫ�{�M'�2����x�;C�fw2C�^6�9��:�)��DMn�(�&Y��n��)��Ш�3j�erU�^��Nb�Q1��h��=dZ��e�nz$��"I����1O���l�n�讌F+�v�[��o:0Ӿ��(r_!�z>�-�>�S7�e�O�=@����c�Lۍ��˚�v ;�yvz�0L�Z5~�vf[���"_��K�o�8Vۡ-縙�mua{8F���{:�j�is�W�}Q�Nۮ�Up�}�6�YS��R�eC˦��w�3]�dv���cv.2^F�ñ�q�a���]9��x\J�+D�n;7���Z�*D�ߏZŽ`�d�Vڸ�9��َ��8 f�ף&g�Bi��C���(V,�g8��4�Ҷ�Jms�v��,#R�$@������ԙ���a����<�֬�W�8A��qt����&��^y���j_�nM���h���	��]v��Q.�|IV���GY�,��Q�2x�S0 h=1�B��Q�%���{�p�O}T>�3�>��f�gQ�ˬ�;XlSPÞ�]MS6��'�!{��0��;�1`%��f���w=y��y���#�"c����E�
�Liy��
P<~�ۡ.��q�غ�=�ц��+�34M�������7�V{�fs2�
� Q��׏���d��;��oFp]�Z&��P�_���0�DKȎSл���Sv�	�DJ:9gӮ~W6�T<�~�*��Gg
R���0�;��#���q�2L��1�wi��S�öqܾ��> �\��g��qZl��ϗq@7h�����H�yH��Nc��E�^k�G�l�ޖ/��ܬ��,��",cx�X�6{N�HN�Fnz��z&68z�]ΧJ�1:��Qc�ߡ����$�x��f���]Gʣ��؍F)�d��5�<��GҔ����aq�9nq��J�V�{��1>z�����Tizs�5i��������x�xr�f��u7n�̼�\�<Yt���Wßs�"#w�S�϶�9���$
Wd��D{�,�y[���j�&&�L����p�&kҡ�yÔ�U�W���z�b��p��X���:[��3���t�*w��
͏���ŏ������Y���u
z�Vr7�f�k����OO����¡{�-��ܩ�bwN�|�s�4�����+35�i>�Ux�*Ik��R�<�b�%ً�VE����VӲ��>)5�q��3ۍ�$�d�@�m�E�#���WKV[*�vi�*����/F
I*;�Q�e��u%�r�+��ic/I�3v�,�j�q�X*�)Y�&�E$^��j�ٕ�����Vrݨ����z"=b��o>ښ�L\J�����101ɲ�waf��u�MR�����W0R��W��FU�j{qͫ�A���'1໧�i�FK��3Y��&���*yսl=2q���4:���{u���0ya�<�{�^vte�z�y�6�������'&�q3�N�kV�Z������^\9B
�����׻�����{=i�Zip������8�Hv���#սsڒ���~�k��&���8&�����O1�!0v��xFّ'�M([k1��{TN�7|��	�g��F^���"��|z�Z�"����jiZ����=>�K��o�t��7�o��u���s��u�g*��R`1��	��r�[�o�4uVK��LQ��AR�����w9��[*�%��IF	��B�=}��.Uˀ��Y� ��d��yߧQ�lN�{�4��p��/R�c�>�*V����T�H�n��c���
~ߔ�򵧚���R�`�*�Ⴓ�al���H*Q9<���{��ϧ�c,ƁW��)q��q����5�TV��h\a��f4�䊧�u�{����q՜��ū�0�g��P{,�����;�~������G؁�j������zg����0u��f���q5���u�m�2hx��o�,T����E��F7~���˞'�w:ae����j�f�<�i���3׊7-uGF.��n?��o�_]�	�|���;��R.�|�8���M6����n�Y��M|v6��bC���x��g���hL�a�k���Q*�|�c��F�����;>��T�R�;��'^�8v���*tUV��c,(+gXm��$'u<���5�B���y��Y�3cH�X6	}�*�}�Q�ʺ9VQ̰e����r,�Hv�f�����0�ۼ�G7�(��U��AU�7J3�7ܐ����Y��s=VHϰ0�ڗ�8�^���*Kgg8�:��EY��(eG$��Q�$ul(6�zv�R&:��5ϩR[;z8T�\^Y��B:E:6jł��gv��i�@ڷIb���u)h�:�n��3�29U�={�w=�u.��%y�
7F����Kp�SI$�I$�I)��b�~g(\ّ�NC��a]��1ۗ8I,8��vb���w�iҨq,�L��XMjiej@N�
��@�Ւ��C�n�Et���i���N�ɦ�����r�ҨV]|�e5�tp��Q٢1He�A+�*˘qg���3��c�!� �A�,)8򘥕���$E�M&�0e�s%wV�@�����YF�yg@���]��4��kv��.�5�q�7�4�:m8�[�u?�:ƭ�1��������-N��nomgo�8qEI���(��s=���Sm�}�0���v�9�a�1�L��Y4�*�,�a*(�X-L�bM��@�<�E�nū+��-Db>��S*8k�aYR�0Ԛa�1B�q���f�-��D0�e�ŸŇg4P��*�A���Q�#�B�ѳ�Wut�*�';3�VKV�M�ӗ:�M�Yq�:�����[�?���d�CÑ�R|����.Bɭn���3�����9ڢ�p�ݜ�yv�u�D�VK�&qQ7��j�ݺ8�F�G�6�;]b6�|��X��Ӛ��&��9�5,VpY�%u"�㜐�Z�Ľ��)��i��_��x��ae�T�7�������/��x����3�K�A �e������7u8J�����uD�NYo��*!�ks6�Zk����03����$�V�[e�&*9a��srn��A�AH��)lໆ���gS��]�f�-�_*�W9ec�ެ�/�~�������{�?�V}�gô��üE)�y�V�%"|���4"���v��б� ���9Ue�&-��]��Sw&S��8z�丬g�P}ƀ�����kKYPf�� ���2.�o�[wj�����L�[���"tQ�]`�<�4R�6a��j7�&ԃPr��zc��.l�
PWt#�j�ɽ�k/���s�<��it��&r��@x���
Z=3�f��Z��u�Ùa��k%�Nt�9�8����y�:��0��&�9�!{�H�>���Ζ�f�Q���:�uO&�"�욄*&c���֖LMu��T�ĕv�x�����f�*�Ci&��u�=��x�s�\J��_dj��/q��s\���a��Vϗj(pR�5�%� ��3R�tJ�ۜ,;� ��F�_�Hcs���t<����2&�x�����(W�,F��GKT�������\:�Ƹ��IפG���e���u�<���tsq4)��8��5`�g;.}�غ⯵��JU]��Q���8Pw{�*�}��#��b�=��Rs��Pxf�t��W`�=���%j&����R}i� ,�vq��y��%���u�=�MV&E,�����~�{�)�zߦ�B��_^�:f�SYJ1D'H�o���]Pܑ{�=�9����-��.�4�n�v�=��c��Ѭ֐F��;3,�M0;Mᙐ-�{Z7�-=��˕d฻�Y������5}���-�QX8@֊�]B�9i쩿9L��;z�]k/C�HW�ӥB�ٛu��'���h����Ń ��IM#��ވ�%>��+���T}�T.엲��I%o^�Pϻ�nBv#C�5�9"�u(���4˱(���a0���p��[�{1��+Z(.Jn4�b{%E���Nz:����WMv�ּF�� ����3E^�%ܣo���}���˔[�/>��y;���4j)_?"�:"��H�Քf�s:ʬ�w�hS�+�}S����wPd[���Iߔ˼ӊ^=h�]p��j�Ё���v#6>�f���.w�m3����C���F6�#�������+���VIZs�w'-R\ea<d�\�s���#�o��D����#]���jp��4��:�ޙbS�������bJ���y{# =C��,m�so�or ����Wu!Y�X��=(=�y��)�Tu�}���GO��;&�jU���z��0���(��۔��w�+�txc����Z��aj�Ǜ�&�cz	�m�j��c��n�bi��6bU�G�ʇ
 {s��[4�o�>F/PQc"�P��++4j���4x�
NWj��ު���b7����䳚�	@��������{{Eg�e}��m��N�6����f\m��ͥU����P퀉xR��˻�07k���by��iD̆���̯|�����=�u�d��&L���EgM�)3�>��oTȖ�2T��ST�l��8���|���q`(�#ڐ�&ύl�9�˃�w,T�iۆ�O`�8k��&2rvA�)��ٞ�~I��"S����z�F�kN���uo���6E���;8t�g>,��C�|}9~�ۦ��uH��n�U�c����a��@u��}�Ŗ�s���.@�����o1�Y���gP}߾�����t�>,�G��tݠN�:֙�˲פ�%�{�h�~޶=��p��a�4��Ŝ4SS����^����Z�Ư���0��m���쨗����&�__a<�<���Ƃ�0�>__�aB��DՆ�n�!jM�v�K6Q�@�v��M���Q��}J�_�$��֎_ �ӍW�B2s���.B�q��=f�b���5x�*1����8�򇰡X��[��H�o����Y�?TV` �B�7�[/�v��{�ɥ�l��~�m��
��o��n2s���ٙ%n'�{�{W^^/m���4�YE!�5j�oq��Vٓ��Әv�
y����nB�7\ʷ���Lذ�<ѻ.���I����ӪJO�]��, t�Y����}7�����|x��å֦~1�a��h#G4�MRO*��n��hO|���x�g�y{s���Z~ӈ�:h��G��s�ڡ���㚰�[:��{�:n�TG��_2L:|��:I/V�p�^8���qX���I�;����l�..#�mX����l5Bm�̴+�φ�Y���3P�D�̓���¾5��6~��}����Ŵ1�d3��)Z>����ǆ�(�/yr��y�1%�8~���N�6��ZQ�|�vV�,�+X�!C��\:�޿vW����؀k��NHx��@ھW����i�h�{p@�Je�кݤ���f�;�2�P������B8J��)t�gpX��J\c!E6Tr�~�s��~��	����|g1v��3�pSW��zO�n_>oݞ��ѽ�E
@!������_O*�_oyYq�zJCM��nZ��ό�1�����AI����߼P�D�����#�=�,�7�uAs�(��.������0ߐ�k<���N鸷DV{�����|Y���wVp�A�%��-��7������UY��m O���y*>��yq�Dx���oE�ڰ�#N:a�1�Q����-zL�.��-��^Tqqqr��r"�����f�������b�0�u����]}:wˏr	3�A��zz�iR�u��A���3,��8zY&aV��iÕl�mZq��<�eh[ܱ�:�'�o�c��enQ�l��&۰S�2�
�ꭇKK[J�ޜc��hAb��ge;�Z��L�l�{�M�نW���\��Q�`;CyZX�RJ��>ؕ�٬��X@����94Z�s�nG	��S;
e��s8�ַv��8�V��g�hX��r��`J&���}"��u��Y��^T���mV[�"A�z��"�cX���k��=w������ˌ4a�1�mh;����݂��FM���X{�+�/n�G�O��+�LD�DC2���A�S���TX�Ժ�4X���4ؔ�V�����qn�r+��s��+���`㜙�i$�I$�I%7k0�ܸ�uVQ=1�E,�_rB̭�*�p��o��|;[q�	ʝ��jr�_^ Cxxc��JZki�mu�Z_j*o}��8��p
wǭ<�˃
_+�.�l|���8𛥸7xK�L�'*��:�ʓ��h�k����Y�}tTYD:݉k���'����.�*��&��(.�Ep�]�[V\���|9�0*���b/,� d+��s7���V=�5�N��ɏ���xzQ���@��kDo������&n���i��,��k�����aT�V�gcmэ�}��uW-�(���eJ䂝:!xyq)$�f�i>�Kpȣ�:l�u�B�Wl)�˄��4*[�Typ�z�\��keݸh��g\8J���a���(��mE�
�.%a�E0���kX��hr��a����S	���T��E�L��b�&1,E-�
j�Xb�mh���f�Qb�y�L_.DUKlDF3�Ê��Db�R҈�҈��KJ�D��aU��e�Q�(��2��+QLZ:��y�oQ�r��#�j�l!�:՝��W�#��%�9-��@���.��']��PW�0H�ܑ}Z��;�ڍVfߔ�8G����/0�,{X6��CN|�ެ��=9]��ύrDQäq�
l8��L��<Ƨ�\�f�m?ρ�CXCL?[S���W�����V�`�}�OZ�w2X���nk><D����o�t�^#R�LP�B�(���\{���\x�vd*v�'��7��r����B�#�����|��Co���q�l��˗=�$��S�{_\����D=���"��2a�B$�����N��o>�˦7�qf��-
��$@oS�6}�?������l-�n�"W��������=E�Htl-0b7ET�K5��V<aεg(���S�V��v��G�0���U�'�}qf����yhq'�#jlVj}�{ۿ{hN�����NxP��]Bc%�3xVeť��;�#+=4�)|��9}��ӽ�׈���c~d� E+,� �bEg�����YGV���2��#\G��p���_�x�0�����;��r'[�}y�VF��f/��/�ǈ��A�㶹�So��|�iC:t�ܴ�-=b��@/��S���]f�/��s�&�R���y1i/��FX�L��/T�xO���Ɗ8A��b&���,����Iu�||Yη�x�f&adg�ݘ��1x��s���c���>��_x]N�oe�={�嗀���i��d�%�[}��t�-͞y���Qt�v�Q�����@���'2������q~o��C���P�:�*�3Ŝ t�K ��A?;3m�֒i�o^g^���.�ڇw��S�	��~l���1J�λ�UQ9Փ=���^3-��48A"�ܣimo�w��΀��K����.����!F`���u��Ĩ2�Y��《#Ś:k��Z�y|�
��Z�u'v�Z�~5�s5�.*�8�
���G�l������w��e��'�x� �N��<Tק�0s޿�� ���;�E�0Μx����]y~����;zX6Y���f��Uҽ�n�M���{q�;�2��t�m^��������/���3V�;����q�O�����U�J�2�>�=[gz�i�]c���T��B�~��4��.<Iӄb��o�GW��<Z���]{�yL�n��_�i���>%�b�?z,(�c����D����|-�@�%�z�}h��.6pѣ�E
!r��L�<s<�o:/��U]��+Q����Ȱ�<�k�!K�ۆ��h�W�l�=�5�0.-�C�Qd_O)V�������1�����q�7���HF���K��u#K4G\~��
A���I�����P/+_s�R�?q��NB��O�t�'-��!��w8��3�٣��> (��_�m"��J��9~x�ngE̳��,wY;W���A�I�6
N@l*�yʮw0�V���/���ƥ�*:9h�)q���9�;Sk�	���"����J�])S���H�b�h�:SG��@����4�~dLV?��+zz���ҍ�R�:�\t�&l��aE�W>a��ŕ�H��B��
qY���}W�#�hy���,���׵A���Q��5��,�<�J�ח���:��#��g�|p��=0�j�*7�����T�YN�뮷} �0K�*�.1��L�5�=yY����Z�85�5����؅E������:Z"ε�־��lf��f���0����{�83�d�&6S���(�P��|�ዉ"���LV��0��o|ˠ��-:�������$�o'����-q�E{{��"zMޣȱ�0��ũ�r3-�e{������&�錄��!���>_h�zv!�05��{�~t��i�Y��<t
Vt#����>+�z�b�Yaz�!�hq��,5Sg�I��.ά��r.9��4p�B�˫��\%�b�X�:�>�S$��R��GM��܇0��H�0�7��@�a>�v���93��Z�E:Sӳ\o��VҬ�\�	a�������^|h��=#i}��W�Ӯt��إ���7/�.�2��J�k�[�%�:�oe����	7�ȳ�G�`C<�#��Ϩ�u�^'y2���a���C1}qY�;�i1
��u{��X�(�Z&��3W���8����u<�3P�z�����{T�v�*5���4Y�[೰�M�����-s�QU�=��y[�]K6&g�ٳ��ˎƘf�Ƽl�{/g$�~��z���'Pä�}��*����}���r�<����ƭ3�VE�XIG�v$�r����(� �L,>k���Y$91μ�\KW�@A7�I�t�~qP���#�b�B���`�8�(z+}HOD1�h�=.L�Ƀ�ӓ�Y1N������ӳ�������|E!\��X�/ə��T����R�į��d�O�׏�?/�ǵ}���)/V���=�9�x�6L��t�yT	[F`�w$����{B��4(ɡ��@՟�AE��u\��-�� |���ݲ��	Z�빶�6�%�^VC�D�J3���sP���V����3]X�t���ڦJk�ﳙ�?K�
+�l�;2���t�B&#*�JN��P�cfq�=4a�q��KO�\��<pT̹��������9�|t��3�K�9`�;�{'9��^�:y�P�+zY���H�B�h!Q�5�ݼg־��~�!^+�r�8��jD,�f���rz���e�����y�l�����V{V��z~𵥑�����}�㲘e�$V��=��Ҳ�V�����Շ����h[醩2�9�M���+���B��'���C�/*IDgyf碣������l�ouW�@����;U���aO�����w��S���u�]Tr��E�.�yQ�=���e��=yO����8)e��iªus�`D�����b���W���ی��3_X���P�>B!�K�3 f�L-���;s���\	��G�����/]��H�4����e(��pVAFuf��[{p�B��G��׬}=�#G��D������"����zp\TG�^)�a�؃�%ero�z����5��xy:���|8�Aj�
!Q�W�=B4p5ƈۿA�;��?b�FQ���Ys���R�,��?�����_W�1GN�q�~U��v��$���y9�.�\�
�����1��FԾy��b��G�x��x��/���{U��[��g�瑐�6se�dvl�����ˢ��߽N��w~��Dx�v��P�ve��ڞoo+���=2cO��=���+�X��Cg�Sh+Zv!�d�x�μ�ۣj�{�W����������>#p!�(B7*�uû/O�n��>sJ��	vne
�3d��D��6�-9��"|�{�����NT~�H���U�;>�-���,+s�Q�TX#�S�l=�0�� +�k��]���U��xx���0�FV��
 �4��Ԣ(�-�|����Y�������ΪUݙ�~�gk�!e�8X�*� � 7���⻩j��2$�y�(y�l�29Z�1� ��Ys֭���X'�
�U��+X�_U��<��/P�7ß{�Y��`��.���.�+�MVO7�-�t���a�r͛�D����Mѕ��m0<�ݺrgIF���\�����ͣ*I�q�����q��8�m��Dra�{.*�s]�n��V��w�Lf��w�M�\L�3�҅�����u�.gwP��ib*Efu��nwr�r�@��{Q�z��cZBq�MWq�z_Wh�d+�i�sb����l�X����t#�c��b�Dɝ�)S�ޖ��M�y�k���s�����3{tݴm��e<�2НvV�tU-��㻐t�6b�2�=C�#r�Wm'�������I�+%����7yv^�3q��⹀��X�ܹ�=��.��4�6��b��̼��F��J�mF�:7��$�I$�I%j�.����ݛ).�����&~��p�g���駥I-�k��>�v_��Z�*���S����t��o�Xĩj�n��@C���bn��!{��c][��SL1r)q���+N�:�ř�+5h3��L�YJN{+R\��v-�U�;��8�z��}�/�h;[�wo�>Z��rj;�N�"��\�J'663R�D��%�X�*��_b�u�[�oZ�.��%�����_;�#Ӛo�)k�Klkޔ��6݌�s=BE��ﮊ�eg^൫8�{k�>v3V��Z{�qjۃWҡ�"
��2���(=z_L��^�H��×�m�]N�G�y��-]�N�wp�^�ȭS��;}ݳs��E8��B��s��s
mw��y���y�w����F#�í|p�b�+ET�(���x� *�AQW�� ��(��"`�b�KSL�(�L'����iD����DŬX��""�*���X�z�WM5F*���ڌL���EUf.��Q����"d�U#����"�����͖"3V��"�1fP��EE`�TUb�L�U`��Q\҈�|�n�P`�dQf��w�{�*۬�Iu���?� ��|�����ɡ�o�iy����^�zY����yb޽_���V��7��oy����|x�% 8�g�Dj������֙����z�Q�;�d�,�8���|iz�l�v7��(��4�3j �vP����ʴ�=:��gj<h��yiӇO�E��y{pgzjv�9n�T�^^#������^ F+�S�.�V3a���1���Mo>N�@�%XXgnz�,�0�ӕ���
/����`��^�Vk��~gN�GZ�_x�(n����W�6������&,�����������&2��	ݱ�����z�Ӻ'2��w@�xN�=��%�wRAv��P������F�t��=���i�ǔj�WQ;�>�g�cv��Ό͝�\��H�tƇp���d��//��-i�k��/6�r�A,�}���_�DN_p8E�1B����9�=i��l�=�������a������X?iF����U�>u���ڽ�+VpѢ0� O�Z5��d�`k'����ڥ122�X��%����z��E�����_!��.>?.�o�	u ��*g>��mh�����a���Y�_v[��Ck{X�7B�F6�:�t��HJ�q��v�Kn%W��S
x�ho�ov{s3�~Ԧ$~c�ٛ�:G���%��<��4�۴<��oHR�w�9���>���=�Mv>�ND�*���k�G�`��-��{�e�tqk|�b��EHh�%��<�t��i��[Cj��%}��wC 8�l���O��3 �?Ud��?+���Ր�#�aFO�A���I׳��{|z��b:�姎�4~Ȁ>Vo��6e���{�0x�Ǟ0W�	W$�c�ń!�F��]��5-:z���!ؑ�@Z[� �./�Gt�썮�/�g �	�W'E���8����o�`.�g�> �=�c|�0�(Gz��.$߉������TaF�q�]��h�+����;D=��[�3��Vt��O 9��s���ѺXEb�^�-/�!>6y+4�����e���
C�a�. q����B(�$Wej�/��������&f^�nm��N�EE������)���/h���j���1WO����#�{��<,`���#�Sb���0�:.����g��I=j$��wO��r��qzܯu�^k��<�?Cg'������o�*w[��BqC����R"|-i�<l�n@�3r��҈� �Gx&^S"�~C�CM�����X���?���OR����$׵��jp��S����\l��L�"l1�_�,�-i�J4�K�V{����4E�~!�H(�6"�>@l
Y�y蟏z�ُ�RÆx����u�W*�n�����ҼT�Iժ kisB�3�՞�oN�"�:n�n���7�����X�Y���e��]߰��6ۚ���j��T�ZA��F��~�!���X�P�K�Р~&D��Y{5`�u��Ww�_�����J�۲��nO���;t�ם��5hh�Ǽ�Z��|��<x�eEz!7���pgR���}~N����S�r1ғ�,N{|8����/���e�
8q����.y�(-F��cg֑�]0�u7P��5Z�5� �=��Eg����g]^t���xYFC�O ��B�N2�>8��H�S�U�>>hk���x�8�Ǭc��Yx�e<�w��uC���
HI�N�ǹ$� x��5�S��s�"
��~�GWԇ,.c�N�~��KL�K�;qS����zf�f*����;�`~�#��&��G�/��ur���9����&j)��;��+�� �i�)��&3���w녎i�x�?'k�$�����ٸ+�l�l��=����"�dg��]Dt�®�fԫ��HF<���~ƾ�y(�(r�����B��=E�j��P?4#�>\�@����6=�&Q�.#��������S�J��x�ąj�ȩ!*>�P�?[��I)�:F�l�5�H��,�5�O,֒������5�t�}�<�,�������G�z��B����MāFr@�k�!�*�f�z0WL=�X�G�3͂~�.��<;3�,�<9���嚴���_2N
Z|~51FN�����������0C��nL6��W[�|����-b�N�^Qר��L/O����\���A���]���S����u
G�iNÙ]J�:���ޣR��ɽ���)�j��re�L}t��п=#H��!����*�Za�<x���ˡnٯe8*rJ�C�}'>y~���<}���)ᔾ�+Խ>|��<~���^����!�������sj
#�� M����;�L�Ɲ$�6~�Ky[���e0υ���ve�GR����P���qf�#"��g��}�Z��mJ����cց��E���NV0�qa���վ������Vt�\o�k۹3��1*�d��E��o�~����`� �<&��ܸ�ڶ�ޯU癞����0(�Ay2,!�x�\�ZoT'�&l3�s���c��;eiM�pݫ�[�a���I?���'2���şYG�D�߄�1�V}Di�W[��䩻��0ݡ�����1�:n �2uK�n��5]��c�t���� )�}f�b���֟:� 8|\C�aiO����j�l���`�0v�����4���=����̓�V�eSn�z�#�T�>�\���Z~��z�
�t�[�W�n�8t�D����D�Y�^89���
���4)C�[�40����,���^;��;������������Z��:t� ��Q�u�n�88�.�ִ�.#A�|v��tS���� ��{h�Y��n���Ӄ����wlg#n!����[\������NQ�=;y2�hU��oug#Ws�D(%�AK5��_>��W뉵Q]u�.����Av �Av�������̆�}�>:D����T~�-��j�eǨy��L�ʏ�Kiu:P�/��h�����z�D/W�T�j|D~xx�s��)U��F��n�����v ͝6!)N�>�}�]����o�ob��/X��`���"��G"�� ���g�_Z��'M��:^;�*׎�ǈ�(�\.���I�Ydy�Y�=ʌ�7E�mC�#���D�KhM���U�a@ѶQ?i�~TC�<#k�ok=���W��b����$��Du�Hv#��fKk+��AS)�2�r����e��q��J���)��T�yrI�Lm��-=N����]Q�_���3vOx�}t�̗�ŏº��g?i�G�/)y2�1�7�G
#�ޗ��#J#3X�1��y�7�zv���cM ψ�$3�N�j����-��knJ�$2��q�9}5.T�t�B�a<�M��N���X`���s���馅�^ |�����{̒|�E#���.K�7���P��u�J����9	\�#������k�Ѧ��{i��d�>�0�(}�
��K9�q����.�zV���<l�����1"�A���ǻ}W��x�K�s�}s9���!Jayӛ"ԫ�9�y�:̻�X�n�53Îf�ú8޾z҃�o��/N���H�c���d*��B�j�Y��Ă딱VS�c;B��p*ԇ�B���f1����V�+�7��aW�L֩¯.oCp��:��vgL�`uCe���붺M��_
�죝m��T��7�B"�5�����N	�B��{�]c�̣/�^���=;��1�K�68S��*�aWyUHi�y)� ���w�cE�d��r0��z�d.���kS+\�P5kF_�idqUm282-[��ܡ��;�k[���
��\�Ü>R�<1P/nJR���#}�+��C�9ǘK����B����]y��y��]���9�v�㇪+ߕ���虒� �HLwGp�G��I$�K��������8�x��$�e����[� ���WK#��20a%��0�w��q,�rA6�`)��;�u�)�)䕌�
�J�N�N��$lV,�FEE���V\���S���	��Q+2�aFRTn�cJW�˱�1��ZE�P�U�LO��!e��E��,F_�r����3/�����VW�Ȯ�������r\�� �n�7Z+A_+�t�'�q���ɐ�c�%Y��_!���gʮ��4��%��$�
��A�G.�J��
��ˤ.*��2S�������F�bb�nަN�
h�A�m�h�A%i�9���{�w��{'R
��K����R��0[P�Z�����Q�Wh\�g����sGU���"+�Ģ�X��Q�VVJ��jEQ��V(
���f1�(����1�E�E�����(����¢��UAAݒT��!�%�m����*��3�*"�S��1" ���6�VAQ8�@\2[z����Z���,�G���*�B �O��I`���a�Y��\�j9�ǖ֘�M:+D�o�BjiJ��l�cl��w[�w�m6�V�+.�^���9w�1{ϡ�o�=߾SĨ�9O{fG�6
:u�����{v�߽&��qQ���C�
.��f�g�W*�,�5K��A�ۖhb�HV)�,٘��i O���܁?Q�5U�����;�I���4���훛�G�S�\ק����AZC�a�ܪ����6��x�X��liv�5� � ͽ���ɸ/LD-�OЋ5�1�~�!\W���T���a^w���襦���ȶ�2q�u8��k�֧`���&����#�xQ�B�x��f���~��X�đ�^a�1��:x��^��z93E�Lj�쇭�E��d��Ooy���_�\{�}�!�Ck~>���i�:�<��x�����
7���\A�-x�O�����m��	���{{Ț=@�*�(F�`�A�d�=(���q}:�����8n]�OQ9M��g���n�)׮{��9�g\���./��V&aG�5��9�],�x�(��_���s񭲃B��Q��r�Vt��{���q�'�b�^�"��f:GS1�r��zM��<�K��^C�4G�×��Dq���t��]���ȋ�d-Xp�G���<p�&T���w=�y�D�Gjd��׈>!����x���P�a75C=��<.mt6E���I�zyP�=���Y4W��\ԫ&*�YƻN:�V���$�V�u����hD>a;������}��~1Y־�C^^5��g�^yt֑I=��/�o��dㇽsӺ�6،{�Yw��<�p�>;����8��ꢃS/�寨��/�z���<F����4����r��C���X�����qԾ�"p�PN
��{�%D4h���y ��;��,]��k=�q}.y��	y��x��/��}La�6�Ud�ڋ�U��pT��k���?��Æg܃�Û.��fZ���օ�X�g��P�(H3�F���坤8R�K}�G�/`c�Yp���07�:���!�d�f�[J�7��n�����Q�\%���y5�����xq�30��Ў�-�i<'������跷���^����bI�Σ%I��򞐩IUlQ�EޣsMtJ�%��8�q�S��yi����������7��s�5}C�aj~\��~EiPͱ����ɺ�g�~��R�	n
f��x+��)���/{�)�C���:������;W��,��Ƥ�{�P|lB+�z�
����K�ᗑ�F�p��f/�۪����p�i|kㆊHqӧ�����ϊJ���g�ЫɆ�_9,���N��x�<��>�foJ�L��zn.c�N*��f@�p�嵾�*���$�6f�e�Ap��/���MH�߫%\f��{sY"���,�T�Hn���Kø�,��1� ����e�$y�(����e���W��u@���F��	Иw1�}~�t�x�#>��E=���ן�'��{Z���\c����&ŧK9���Ň�������\��-"����<�P�xfJw׎��.> �:����d�-/�s��x�xs��;��3L�aX(�d-��>"�T���ʸ��Zz"�)J�T����=�(ic��Õ�uo?<��.Z{����р�B�V�ٺv;2��z�d%�ݫؾ*2���զ��t�b	4K��M��{T��8�$x�X{ɐ��z�/�.�I�x�Џ��Ԧ������"�vսc�c��B:w����Ω�4�l[�Ur�A
�n�Z�}� 0@1-x�C�w.�{�gQ/����F
�A�#BS�@R���zo�w~��8�8�f����&��Yۦz��1="�
�'�~�z��ָ�2l��"��k���d˥X��"�ԍ��sTI���u��.$�:~�NbťHd��G�{��!�\���K�6t��0��H�O}�6�L��}H�ٺ��S.�����<hr';X�7Y�~�Uj��}?(�q��Iz���V���/^�u�*�n���?�_�q��r�G	�g�c��,�.W�x]1�Ύ�"�j4�=KH�������W���,��K4p��p�,�&~���9\�M�ڟNڤOG�{��P�y^-����N�y_^o��!'�=T���]�� ��F�Y��[85����.���Z�2�R�ۗz�I�Ґyi���:����ʹ~����wt�}�dg�� O�~����^yY@T笣W�׬ֹ>:z��Jz^s���ET^��ͼE�����N���5�;�x�F����yOl���8l�b�X�����T��Y�*fl8�#q���ŉyW=���b%b�$SB���h5:�j���r��"}�ܺ�cO%����8F|3lڮ�:}������0�g�bI#Q�Y�+�#�@�~?x連�w[�b|C<�݅׽���u:C��Lo�q�yq��'�����~-o���R�{�/��'�|<oVj��A�����Č�V����<̹*-_q�p�.�\�+[�����i�r�n��1�Pwg`5(T�����p].�^;2�;�O���^�߬_��++q��P������ѕc��}T&���b!b�D!��r!���R�!�TYt�5H\jJ���񳇁�;�����V����k�7�ܑ9O��!�K��EG�guLB����>�}+��	�j�A�&��8R���7��٪�����zx/,�D<Cܐם�1ƌ�Co�*{I+�^!.\�Bo]�H�5�{j���7��w}=��.Wepo�A+�����g�F����$���䡾�<�&����(<���Ƈ���j�B�6a�9��?n�{����z�mZ�^�
:F�hf����+8�k�᠋탻x�'y�cS�\͘�w�R��fX=��+�����+�zm˽ I���.��r�Mr?G��^�x�x��|n�.o��ykSׯ�>!�9ߪ�y��,��5z�G�x��'�`��+hnE}��'����^����\�W��L(���AnN����ܲ[�d1ȝL�_-"���\�N�̢��ƕ�r� �Lp�5����Ǐ2�G"�<g>R�^����y��慥�L:}凴�z��,�sŤ����5 �<��b%���-i8�C��CF�xHw��[���m� ���fcY���j|�)m�u��;{8���<�0�,��08��2�-:�Fvy�񑽺���w�*Od�b�ˆ���ܥy�����W[� X�Dϭ��d��Z����9�t���|�f>Yޖx3�-����+�%��]�����k:��`}���꯫���&�Y�����r�$Qcb��^0o.����>v2����<~�o<� Ro��8�.6Q�C��f�ʜ��x�փ����\�����+,�-#�yZ^ۗޣB��>6|�R�v��=k�,�"���ιE����X��~f��?���K�^׹Ew_fqP�%���N��6p�ӝB����r:��4ٛ�w���)Q�'և\k��t�(��=X��؎li�a43���d�đ+X|��:��#*Vnt]�ĮWJVU�2R�b������5�n��We�D�=0�����kx�,��Lr��	_G@���́Bp��"�r���ym΍M�n�%�E�rJO��a]��z���j��I�im�gA$m��XM]����[�m=�IQ�u0�i��N�*��>�˰F#���T�%i9}Ρ�b��eu歧S'k�u1}��]ԃ����:��ݾ�Eyk3��-P݁u`����l�!씮\���f��ǳ��Z$
�]�9i��N��K0w yLA��':��+gq��c��m��[��,�Ζ�z��8�pӵ�4��E�g*�+����o�v9ڦV��x�a�:��b�M֘yx����*xkUܪ�TƔaR�F���(��A�0_w[��X��ok�����JI�Sgw.����������y�OE]*C�]-x����L�M4�!�V�R��R�.�d��f�,B˼�p4%K�h]Ւ��:�#WH�g/,������[7x�eأ� ���
��(�O�E�vK���
�ӼK6���2���ZJ��ZL�3Dc@���lc	a�)Z1�A��m	V%ZU��`�@�&%NJ)�p�5�Heҿ�'F�IY�h*8V!(ٙnP3#�b���ę*,�!��Řn���ٰ�Gr�4/~f�>B�P�ɺ(V�l]�k��b��M7�2�k�v1!F�C
�bG3,��Q�1�Wyr�d��:�tr���vwwVk���	#��jeH�Q`�X��H�j�)/��(6+���1��*(�b�L0�ʂ�Q
�#�+%@QTX��ް*�*"�07�E<��(� �E�V"�i
0Re���:�<�xʂ�x�,2�`�<l��`e�����%IƫDĬ-�U�dU��6�J�#VI�I9(�>X�>9��g�����F�F�}j<�r����*Q9$%�����>����:�b�]�9Ѫ�++��o���p�੶-����}��jp���_+b4
�6�aW���<���a��MG��*ٓ�J�SsN6�,�/I �>q���X�[N��ny�Z#Y'���w+��{�(�R;�=���w��͙�r��,̾��qW�d�ڃ��^=e�6ѵ>��=X�Q���XZ��MwA���g�[�aI="����З��uy�:a�r�Z:ݖk�hp���]f���k�ȹ�)��7�OY��Ҿ'2Ν"���%D�{}x�k+�1���{�h�Ad�Qr�މ��q�=�ze�u+�����0�xߋ�g�n�ͮV��G����`;�V�P�`5�����t����ˌT���9��o��A�/3J���D�l3�3�g�<��f����/��`�a�tuG[[�����3�:*�+s��7����l���͸n�o���x.l�y�%�M�cTð�u����D�Ys7Y�\vt}��qfh�fRv<Nᦖeɺ_��rK&�8���v��K4��v0�3��\��������V���E�f�0y\X��&8�(-�F�� �B��q����jV�BǬ<��ʽ��<]7 ^�: ڧ�x�t�+M��9�U�/�.H�s��_&��C]�j--K�Κ{�"p̽9�n�l+�mEj��Z�c�t��' L��Vxvy�t�ç��[��~�T	�Q]�#;����+3)�ȉ�a-�]baTw���Jy��a���`�v�1�<�q��UNX��<��Ӓ
�B�Vv��2�%ǚZ�����N-��:��P�xJ(JB����Se.��+��=G��\۬7?gj���PH����3'(���`�aL��I����T�G���\�� |/�W,t<��m���%�����,^1J8��RO�0��=)HK��b�~�8G~X��u���ؽ@�]�p�ɧv�Lr�K����EH�]���E��ȥ�"�;��W�τT��r�\Ѯ����`���G&�gOS
�������D�ΩQ�P�S�����|	a{�v�֋��[4+DtJ��w�k����H�⹆���Ůzg����v���Z]3��݅�Q������g�
���:�zګ���"pC�ht�ȴ�U��)�ÿnf�u���S�Kp�M��1ۻ�M���劅;q��Hz���+/;}7��_�O�%�!-�L+��shTE��ZEL�Ҏ 65a��qۈ+'sCIY=��Y|atw�QS��a�mj�(Vv��bZT���������k�G�&4-g�ة�xѼ�y���X�[��%�����Q2�v��)�y��ц�:��:���W@ɽ��O4X����n�WJ�"�!�����R9}���>z;����#'D9'�S���L�ʶ����߆��d-��k�m�I���ț;��|m��/8��[�x㱯ƘH�:�ruW.7�A�P`�zj�� e@�~��WCv��s�a��*v�{3ʪ�_.�5�cQ�Jl{�ь�m���7�)���Zt�I
���5
8A�h=]1���H��Z���.Q ��=[f�6ÇZb��=<;;]��;5�r�P���y��4u+D�=n�@1�)+a�ٌU���s	���R��S�oGkgI����{����\����^�&&��%�_`�BˀU��k��� u��/R���a����9��V�U���'	<��7�l�|��a�2�OX�5�#"�:m��ի5��V�٠*}��Vk|:�5���Λ=���q�p��F�l�b�-C��y����g��2h�uxyq�êME��D��@�$�뻸�a�[)#{��.����iY�Z$��m�OL��:�X܇w�(Q�&�n����kWT���u� ��]�w*�Ӛo^g�c뎆�]Đ�up�̔S��P4w�U��J�׹}g;L���[4�&�F���S��="����R��#�ajor��H�|I&����ຜ�	f��p�讅O����ӥ��iO��9Gss�{νԟv�&^E�[��&sp����B��p,NK~�o+�7���u!b�����wV2���M5P-�n�.etX<cM�sԐ'� ����N�Q�1��䝷�߻WV�P�(�-�W��)�#���]e+	&�A9�N�wޞ�7��<k����#.y�hx�u9/^��)����P}Bb@ټP��U�R�6�5���)7�uD+j?h����gJ�!.�����;yM�����}죞�>Q.Ÿ��,�4b�{i�X����w����7Ҩ�]F��� �bg'�+˨>��^�(��|�6����<����@����4?dKOl�-�G����Є[0���½�˹8�g|r�
��Qt�Fa�Cv��sY�'3��������P�RV��cE�.�v�@�j�E�6<���P>Ĵglx�}��U�$�r��z�)�]��o3��h�˹D���.K��T����X@���,Ĝ���^j�R>�j�H�yY��G���J��S7�����fϚl�Ǆ.}W�VO�,J.b�W P2��X��T��B��I��������i�{���]�aJ�����AN���b��
��T�hK���3m��Z�U8b��,#�E��O^��B�A4Ꚛ��3j�Dq����<箆>- ;n'�fz�IU;C���S;��*{���x��f�2;!���������h�.�:l�8D�d��rn�������q����w۷���+��f���8���:3�Y�������#OfR�Cnΰ�]����ܨ���78v�읻����"�N�m[m�X
hh��W1z��v�|�k��U��h[o�Nה�7`K�P��V�����GP���}[�E�}�V����!�q��B)�J{���������cq�U��pe������9l��R7`�Y/�7�mi�Öd*�}$֐�]ɮlyj�A3;eS�_#��J��������1V�g_S/'WoIͬ����y���}�
CBum��:�t���w���!�J۩y6����R�+P��I$�$�I)\�m�ʸ���,g15HV��h��YV��� �sY��ߚ,�ܷ����xN�qVEm��}a
t�O^�[h�V?��b����E��Er�L�/�C �SB�4�1D�����Jݜ�H�ܩ�ϰ�MZH3����$0����n�H�i�j�5f�F�#�Pw�G��9S�&�2�Y�A�.����ѥqJ�$�O2]�Y'�*��B	�ckr��wksU�T���j�2�t���P�m���IZ�[��s�ܒ���m	R*�B�
AC��+4�d���@6�4�QE�ֲi��D
�T%X�Q[k8�&^$5��R
T6�8�X��P$B*�J�PY�H�m$���ڦ�J���(ȱX�E�RES	DPR�0�
�
�ET,��"Ƞ[KhB␬��b�ROi@$Q־�7�T%=�Wy[�+}���T��J�P0we"���		F�!���>��=�c;�B���[]��N2ZC������x{�X�P����OS���i�um)7í��@y׺;�@V�^:m�1Qw��m7{8h'��])
�����{�����S��؜�ñU�����N����ϭ�+���u!�5�.0�=-�ue��h�������٭�w�qY��\H�
��-d��L�P�Q{g���a^ÇV8b���у���I�5Բx�w�W9x\�^���5��;����K�}ځ]�m���Үg����[�;�г�+���mK����8�3oT�5�ڌ1�l�r
�������Õ��5���:l�Q7}�֞7U�v��#���yD�b>}��4��b���|�h>����������FexwB�a)���"�j�^.��73E4��J�keW�M��zTˋ邂=2���C�t�0�.�"1�Ұ�$���x%�mErV�w�ͬꝚ:9�����5׫D�tFvE+�L�� jŨ�� <X#��YRc�/�q=��-�[(����m�2��(�^��*�˩���m�-�������,aDնO�Lv��=W7��m��ݤ�����D@U�xs�}5�[=�C=O�{\���,x��ٯ|SP��dK�6�l��;����Y�^N���hH��d[�X���-{�>C�?H]�AK
�8y�.λ��&�ϳ6ʴk�&�O-a�Ī�M�ɣ��B0� ��܃��EeԵ��=�]ޭ��'#�2I�B��#mn��'ݑ]4��~��q:�w2e\�t��CY.}-v�x�¼�&�c�v�{��ikPt�v*U���ITI�ʹI9%)S1b ܧP;j4%��o��{;g[����f3QЫbd���R\p�6.���m�<O�ŬbNs�k���,c��M['��N���Ke%��oE&9�Vbˍ] iF�=S����6�#(^��� `���r���ё��f��y~�خ�1���1B7��%�׽��Q��U�iprl�ۊH��V��]��qƉ�l����	�x��oy�!�O�q�٨�N�:�S�����k�:6��5�V'��ݹ�����ꁃ�ܯc=ov�s�(ʚ��z
�?C]���+�&(Θ0,�G�<���ۚ��]��<���U"�epue��K�O�z�CN���G��Ő����dk�9��Rao���7۱T�ܫ�$K�9�ϩU�;��<Ǘg�	u�B��<�p�Q��45�C#Z�l�	T�Շ�t�\�P��ʾ�VV�$�����KV�r�5�d���v�*�(��y:r�D����o�W��u6�����:�3Z�0׽&�o}{b�2�	/���'+Izf�TrvWe#0�"��]�Bܣ̍|Wn�r��'.ﷵ&�r�d�5	�f�C��t���5�]!o�r��r�w��Wy���;�$/��_@�0��
���E�~�'%yx�m�r��r�<�x�oi�G�d�^��z����Ϸ;�(��l�J�A����Wd�W��׬#SM�TX��O�b��x��4�IT�r^A�����8�C:/F7ѝ~E,.�w/i��Fw�q�CM׵m	����Y!�jw�A��$��KgM˙�ơˆv���x_@�^|�eҥw�����5�y#�м�w7ۅp9[؆�sæqoMD�J���X����_@��qǹc��������W���י�,e��잫�K)�A��rYF��q�Yo>Ր2}���7\�v���v�gc�UZ�p�����%n�<вڮg_�e��F�g��x�j��<Om%��m�i���y�C��B�ؓ^�ZR{����K�K���f	t%�h�m��&z-�S	=��-]���A�I=�����e6���
7���d���l\9aɁu��Y�˛�q�h��s �/���"�ۊ�=c)�|;�qXA�o�v�i7�v���k�~��|Wx'�4RNCE�s�V]ar�|;'�ak��rR:BӘ� Yϟs������ި�'K$(�嗀#F��5y��v�hd
Le�]1u�# �7�����,­���J��(���(��歍�8Ǉ2lSfzyҖ�tײz��J�^L/��z�+����ߎkcg�P,F��	,�5Y�k��|鞦���F@w�\oEFz,�`��CHؾ�;R���BEY�t_tpXZ�M\�>�Ur������5Q��ʥ[�ƥ�N-B巼��GÝ����O4�w���q�\�} �_��朷����ˎ�L��p&�d�%K���X�!{�}��/E:������䚭Y���M�H�b5T�U�3Ɩ���fXF��J�n@�ݹ�'}yڼ0b��*��eOX�$��pupBr����w���~���d.�;�1�Q�3������vmŔ��=w,��|���aח��Ö=^�c0W���?|��j��2���#n˜�k�wP�X7��� N���Fe���i,ܛ�� @����p*�{H\J-Ο��Z����T��֮!%}l���������{â��0��<�a�97/N�:0��XꋫI7�i���YUͺ�u�+��zw���{�������5}1Nj�#u �h�=A�Ll�g�q�ؘ�����ш��qn;G�k���Ҽ���B	�8��4�ÑsLړj-���Í���Ҽ��:;u�C�}�-v�%ǜ��ILgf�r������Eݗ)T�P�t���T.�b���oy��ޔ���|�&"Ǽ��5yh�z�S^�Q��Bk������b�P�E9WƆڌ�ڈ�]� 8���w
�i�=�+t>4��O�9Ͳj�t�G��I1�݄훁�5�3� �730Y�ͼ�mS�0�����« ���©�x^fJ*|$�p�pa�N���nB~�,^�X�G�������X��M$�����]�pY�>��s_,T�js)nNK#A�W]�Iw>y�4�ve�]	�:YQs-�g��Du�ˣ�F�fP(�.�f.��7�(�Y���g�ċ�o�����k��t���77Y&U�5�mi��@��o�У�r$�����I$�I$�J榮&�4��+'��t�FBԣ/9c2j�	���V�E�a�{�{�݅v���3׽�y�:�ڐ�q�T�Q�Gjb7�_K�V�X*s�r0��z�����1�|��ɜO3�ݚB�3�xr�ڢv7wcs7a�;c5�c&X�>7��t緑�� c����]5b� <r{)��;I!����[�{��8M⥆�V��|��0�v����U����G9g�n���nCG���+��9��9ap��{+O9hg&�V
ʵve��6r.�c�Մ�.8^�owvq39Es��^.�Qf�:�"�e��[��w5����\E��RA�ea
�J�H��2�L0�QHb�kdT@�[��E�L5
�h��AR��(��bԑQ����,"�1�	
�eT�
��U���P	QT:�͡D��d�*T�"�QFi��aŀ��R
�l�,X�D"�/�L0�R�*���RJ1`�,���q������,��E�5%iF������L�@��C�{���c�m�j�5���][�O�\�ٚD�E3z+6`�;Tt���N�q��1����;w�i���j���f:4���t-j4Q�t�]dfƫ��9@(���
���w<�a��E�?au�tsA��/yk����x*A�h�7Y�x҅�nSg!�̒��e��O]����i�%;C-I���c˳�z�G�R�/ȩ������Vn�C�շwZۄq9־Y��G���� ���+�˾����u<�:��^O�oL�%d���+�v�f�,��t���ᥚ��Z��+,U���#��D�L���-������;�m�oC'�e����5f�Uw���)��け��n�|���^Ղv(<������n&ˎ �]����:��S�D�6��iERq��:�l��x��h�ǘ9� �����s���i&&;���m�{*.0+WT[�Yw�����f�#Y���WwE�)���I����"��̧�9�p�t��Bu�����6��6d�Y�!�{*P����.f��`�~�E�5|�}#�@�q�7�ȓ�e�'�f���	�:�\j���e�s�2�6�LXT�n)�Ľ\9��S�x���{��O4eYӼ�3�C�k��j�MR;����oE���.�5�u�v��3Ũ�yAU�Q�+ђ�o�V�k�����u���ڽ�n����c5}�+Z���4M�s*1O���,�`���;�pwVΔ ��L[�O	;�~�Fc�cӽ�����;�qJ�2��[�}dd<sM�4̻��u�neo����eI7N9���YR����>���P��3hkGp���6_J�T8k���=I����=j�-�01t}��|)ԡ^l�5Pd��Bf=�`��і���3`�eH�@��tʿ����E�S��J�FB������nJ����f?����/d��Y0��o˶iT��~�f��Wv�u��2f_v9���͚Yx�շvWr8W��<G8�pV�Lkn�d�B�5�<�_�k�����ׯy���q}U7ܡA��.V�X�ɼ�q6dWzS�W���Mah)�z��Vb���q֔�!a�{I�n�0�V��rs�n8�j�^|�3+�C��$m�ᵅ⪗�����L���즀ޣ����;}�ə��B��N�fK�ק��.�d��=�w���Xs�:�֚ȦN_΋�	�]dO"0.4 ����K��ftf�kGu����ݯ+�ޣ!���zC5�ם��!�aJ]�!�h�t)��q9I{e��ڎ��}�U���1P��]��r���M���sp=� ����2�5�yd�n�V�=co�k��g����M�����o��Q���k8��;�nnr�~����Q
����:���
nx��kĪ#�=��=���T;�	�P�냑�A�O���.��:8�f��;��%do�����`,;�uV��h����j�����ٔuU��awvkm_����E��e�9�ә[�%B���727��=���k�>��=}�PzW@�V�S�vݝ�Y�)�E���T���1�����(�RK�|��Qy'[�ܜ��bxutCU=�pR���%�D�/s�>�OhjG�s��2����r"`y��b�{��P}ߪf�=��H�����{[����*˩!�-�u�����n��Ȝ�h���T�&gHp#��#$]:��+�l���[��7�����`��*�yަ���˜����3U��Tݞ=@9��Urv*�΅HO�k�1Ox§QuPZw��L����n��Ў�Od��kr���]��0Ɯk@�u"��\��m�<M�5zW�SES��s&�f�]熱`]�;�jf�o���2�Vѡ�~�^�r�S��/6|�-+7]c�b;�T��H��hOd�j�h��aN��s���n$#6�Q9��HcL�)���x��q�7�Z+�J���'������ˠ�d.f��z��L����1�/3ld�\�;b�b���׽%[���u�Vq�V�u��r���*�X(��k���|g���C��(e	^rgR,)i�{6��!l��C�����5b��[l�Ӷ�薂%vi�g�3�~�k�v������z�@�[��̚Ͷ�Y���2��SN�ԛ!�ެ0^1G��lXwb�i+M�	�)u__v�v�e�����<�9���9�G��3���yv�]FvQ��C2i��J/QŮ�fm���bI�a�,���r:c��]_HyS�T�sҰ��e��w��q�gJ�4��hFCv�:5��ᚱ�;lc�R����>�~W�Dl-}tE�D�J�C�W�x7^�YH8{CxP�Uz��DY3L�c�7�57�:P������]1�|�;�p��-sm+䧌�~�4�1sQA3ѳN����n��l���r�u�eO��!ve�ɩ��Y�W���C�����;2q����8��%f�g꓏�pR�8t>�yȬ����պO�s�iƬ`��䴂#L5��/�)	wo�ˢ���=ǉ��������81f6�$��I�(�V�U�[ͭ�mvk$̣��]�������Y��zy|Wf����b�r (��w_+º�n�>B7����.�}AT؆j�7�Z�<�޿u9�ܬ���0���q�a�#�@����(V������!$���O���I$!'��K�*�.M�y�gșa��	�s���G]Wn+b�ETUR@C����voZ��	������^Y�7WM�U����ITE� b3��1�q�
���/�dZ`��X+]�Cr�K��a��y�
��Ƀ�����Y�57[ۯ�Q��=�<s��&? �x�
/� l�����bV�a����&��������'�:a��8���^:^h'/UD\>�u�����@�Q������{�-��G\R1Oa5�?+�	��Yk�i��a�0�7s��fM9�>"�"�5�k���Sʗ�EQUn|"�A�*��)�����\c���a�#P�>�d��ETEͰ6�w��6�f��7$���\���@d%ؚv+��uz�����H�ŷ�&|BTE�k.�b��=i�ܓ���Wޅ���`�m�GB����zq�[kȈ�lZ��{X��f�B�]�'���sETE�� !�7x����3�a�W
�I4Y;�x��UE�{�U}��E��N�&%vPn����BA2*>E��@P[�T��!����B>��/AE���K�i�,�x�ѡ"Ԗ��~�����<����al;�Z3����UQ�۸�;�jnETE����}�5=ڀ�	�{�vF��`|M���bP�f���c�p��l9/��Ԟ�I�)�ۙx]��������쮳dlA��I�U����	�UDY_:��X���y���̏���К�7`44��BZ�y��I��%�@Qi�����>��
ۘ��~b=^�
���t��j������T1��nH���qd����X�v���俍�nB�d<�����HE�X���lu}MM���E�;NI� ,g`��F�jř\B�ӥt�K&��xE��4r����w$S�	��`