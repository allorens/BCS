BZh91AY&SY�����߀@q���#� ����bF^�      �                                 @ Pyl��T�T�ma���l���P�UIU��4�B�B�-�٨46�V��MQ��hT(U*E�)
*$*�*�l��ѡ����mBAf4[I�MV�6 �j��@�kCE�҆�AM0������jѵe�D�F��ԭ�!B��h�B��(,   7b��
�����V�GMt� b���T2�f�:����ڕEQf��JPw��!�ʀ�!5�ZV�   -הPt�v� �n�%U���F��7m�JV���]P`�e4)T�gG �Q��w +� ���JN��U@ڃMA�AD�   v�z�v�PR�ՀQ�m����F�7�y�@v�(ޕ�xt[e4�9�]� ���{�2�
�y��7�y=�Zm��;ݖ�4�9�=�D�I�̫l�EQn   ���ݵlh/yὅ*�l<c�����+�z)T�kK
��]�-��<��� �m�7�v������m����pt� +rXw`Zy��f�)�F����[�  &G��Zhil�u:��B����gn���-�hNr�t-��K���֨���ҭ�֛��v�B�T���::�m�S�CL�a�爋M�5
�D�Jќ  ǯa ֚��҃@��v��M���Kc@JwE�J���1жmZ����A��ì*�]jt9��Ն�ͧ\ 큡�޽�)��,�������  w:�{l6��wE�-���+�:TZ��]�B�]�9T5M��( ��fr��wd�UT�wNtْ�7\ �{�(U���An ��H(6�pݪ�Uu&AH�EP���

�j� UUmT`

���,�r�*��ݜU w��P4h*�P�JB� u��U5-@U���
(v����9�9T(��ê�U��R����Z�T���PU{���*��UKF���MV�� c�Z��C�tUZ��㪪���]@�
�V4 �n��ER�s���!Tf�
�;�8%A�5�         �*R�0#  CLL S����H� �@ �9�&    � 	�S�"R�SM0 &A� 	���jxI�j�����&�� &C �����OM5@&I��z����=5?W��e�?��y��~���-�ѻ{+�ݘor����������������pW�*�
� ���QW��D��*�gk�q����?C�g��������T�UDV�j���;@S���D!Ԟ�DD�����= D��	�dOL)��"{dO���?�*q�=��S���E��'S���T� �x�?�)�C0<e0'C���P� q�8�2C�!��^2�����(q�8�L	���0�	��*q�x�<eO9Ra0� ��x�<`0C���T�*vʜa0/�+��
q�>0�8eN�����
q�8�<dN2�S���0S��D�*q�8�d>2�`N2'�D�(q�8ȜdN2��8�<d2'���8�`N2;e0'���q������&N0�C���D�
q�8��dN2'03"q�xȜaN2����?L q�x�=0���Q����q�8ȜeN2'�q�8�<`2v��8�`N2��	�8�<e2'�z`0'S�#�T�{aN2�S�L/S����q�8�e��(q�8��#�� q�8�e0�G�8�d�/�	�D�(q�8aN0'�	�&�"q�8aN2�W���D�e�(�za2���T�*q�=��xʜc�T��T� �x�<aN2�S��8��`2'l��� �x�<g�"q�8ʜeN0�S� �x�<`:a0/������`}0"��� /2)0�e@x��q��*)�DS���TN2�d8q��"��E�PN2
<eE8�*q�A�*��@G����"��T���2�<`}0�`Qx�
�E����ȼa^0S���+��
q�8ʜeOl����2/�'�W����(�L��� �xa��`N2������r��G����@��Y��p�j �։҂�ð<ZsČ��Ѣ;{�M���d�H�m,\S9������.�#�p엣��F�[{R���7&wv�Ƒ�W�;7C��QK�/^���qI8���������3��ԟBH#~��v�q�ez¸�5iY��à|@{3v���M�ڤ����Tb9ɱ�lSٖ=�o6�\��Sa>�4��7�xc�V,�:MˀSÞN�e|�f��C�rY�>��u�7%ӿ�O���Ylb5�3\�W��/e��Y$7z�B�����C7e�Ӓw\곇�v�>���k#U-v�/3��B�罂� v���\��nr]�6���x�Ptr #dNu����:��[��g8�M���"��ޛ*�pspj4�����\������5pa�j��W.ͰjsS��;�	�^��îeT5� �y�t��zH����;J��Ȱ\�[����(��b���,O5)<ov);��#�-�z�qw�4D����i�h_k{�w'�^�`�[�� �JV8S}�D�"�]��{����k�甝�MպN>�D^l\�jh�ѯ��/oni��w�bX .}��D4M|Z=��wqu]i.S,Yc�`���"��9�"R(*�x"���qCv�SL��;{�̓!�A)t«�Uᣰ�tE��gn���0��ȶ�h���p��ȱ�P�6q�q)�l�Isqqc���ө?r�+XE?���<�*i���v�;,�����qd�Ȩ���F�n���R��p�OnF���c��:�}��m�׹ж�|��s�P��m�eȳVnv�C�>W&^�`� ��0-YXZO��R��6rj�;G��`�}t����]1j��\�ot��<��eV^�$ga�u%��w;wj�<w��[����=}ӵ����C�I��ſ9�gf�R���1pI���e��a]I���]���lhI�y�n��S� ��s^�6�уxNj�������{��4����Lz����\��:w ��hLn��e�*��3��Zԛ��E*��M�~LM�Z�,�mH4����������s���V��5�9.�]��u[���{.w�Y@��Zx����1s�7tk�tRn���j
��w�hN"r@xww[��F>F�G&@�됖����sѼ;�i�����vI������B=��wK�`� 9����Z�&�Դ�C��V�-�tYM�<c�>zٴNN����V�������7���+��#��A�1<�pU��LF�k�wf�͗v@�%�1�<cw	Y���wLkb�Wj��\�@Q����ލ,X�d�
v���+�P{k	s�]�:���b�3��f�KMH����P�Kh�yg=N�C��O���K�4�����]X������;ЪY�sh�Wx��{�_y7��b���VoB��v�$��WJ���;Yۯ-M>k/h�;�f)���0���Ty�w��ݒgwnZ��ݦ�q�R��#�#��F�Dnwd=P��[�UTL�#��u���#͐����S"�wAOw(�c�5�I�+ʇ��Ŕ�'�]�ݺm�Zsm��6e�N7wp9�5��C�&gGK����*�On^U�Ց�d9��\ӥ�[�/�����nR�W/M�>й�dzgOI�Fr�rI��$a4 �%i8��[�"��^��/(��sw~9s��o��֌�� >�(�;6c�{�e�<R�{hcN�F���iZI� H�1c��1�#7o;���{���tњ�B�����l��kWt����l�Ã{�.&b�؀=�Z��oe웝ʵӬ��Kv&����5>9�+��=�d�j��k�0�r�{vsi�����܂���պRSx)�v�"��O���w����<�;�x�8�p�r׵nD�ڬ�qhZ�r2����U�3�Bu��y�����KK@^�Su��L��0����vQ!���E�@ܙr�)W�꣄���r����1Zk!*�� ��;CԎ�ٻ�^�n�3���ΘmE�ݱ.\����S��]��.$��s.���-���`ޏ����:��q�d�Kw�3��y� =�]Ǒ(���n�2� ��K�m���9B�v�ի;�Dj�"8���^�F�մm���s��y��0��q��x�D�1aӷnC�����7�`�� ��x
1�4N��׬hm�;b�Fd��w�$�9�,�Ot�	kt��'�n��E�C;�$��J��4�ȫ�7���wEZ�v�
���x�s/.0�}����٦'�������u�%���d`E;N�J(1�A�k���o\O�j��A�'L��\��9��O��QSV`�T?UI��PT��p$�d��`�6r+�V�.�q�@��8��k���iō�а�xf�L�.��C�p�$&��(=�CN�A�{�� �ѣ+6a�X��!C�N1��&XԞ���N}y�z�>�!��xe��;�^��a<���o��2\�u3�s�.=ӂ����ݘD�7�Wo4ghH��`$e�˥@���{9X"�˪�j�M[��jװ���h�^J�I6v�����2;-}fУ���e^��)���ٷ��i����C��%Qr��e�;�W�6v�H<�D�E�L�;�:�'5��� I�ټ� ���/"�>���X�۸���/kjmE��Į�,nN��:�N�޼hӏ�����71\:0�
(����g�3rav�"�z��]|�	�8��	i r�Mg.K�;��l�񙍾��{�@n����Z��U;�⍹�T�5�|y�R� ���`�r}� va6�q�!9Y��ǑŁ\�b��;�nb|��<3j�#���{�DՓ7M��ho6�o͐-~����f���;L���7F\�,���j[F=�c��1�gvJĤ�,Ô�z�������浸�P>�,�s��$�2s����댫�%	�kqd�v2f�E{Aǵ�V��	�pK�<�58�g&N(�C�hȆs�X5k���޾�Xe	#��<c~S��>y�ϾFoA�� p�h�޹N�p��g9OQ���z��c,��f��6p�ֳa�Ov�0��;LQ����j�&�n�q��[��8��8��X��Z&�p�B5'a{�8��X�>�h�5M�I��:h�H�)�SƎW��!�@��ܣy�CV���g����a���
p��cQ[���x���eԸ�I�]���R={u?'sZ�<0�6J�8��iB�#��Xi���]�02�Ovv)�����}�N�ۯ!#;��+/��_ƞ|g��0���<u�Ӗ�3~���ܠb[PɄ	]��ʂ(���n�!ָ���:��|�X�bΰc�ō�ɼk�9����k��>R-�#����)ۻ�R5�0_�ws`6�(���,��"jN��4sr���r��r��ܳ��E��ڗK��]Հ&_�+N���ː�s�q��M���#��h�qek���%0Y�h�-z�J���c��rL�9�]�j.yN�э�s���9�f���2��wV^1�q�'��@nтI�l�H=���e�P�^7�j�Ԙ;8.bs�&�Pn�7Jغ�q������W����`�ɬ��w$��木`Ι��2@G+�$s5���9۸��H��鑴�������T`�V�pc����r=Q��9��+WN��Arc�����̠��bX���U�7N[3�+;�Ż��%�殽�������L�ћ��+V)�ӺA��U��64V�,�Q��r��Y�9q,@�!�YHf��c�qюv��Rb�OG]+��K%����o��9PW-�D��/@�ըp˸��fN�����9�`�2-N	a�.�1��%�gb[9L�I�m�qL�#j"}���|bO^��=���q>��ܙwo�ŏCΖJ闗.zIljX{���cN�б�1�.�ڔk�%M���������Q�Ōh[�(�	�'̄3�Z�7d]m�L}��i>�mױN˹WC����h��rM�c3	ǚ7A׆��u���5ɰ�]8���cnZ1y��:�o@Ά��rP�3�&ˢ��5��գ�8���b�8�Y���c�y�s�r�8��S�[Ӽ�)sXw@��Sz�2��F����*æ�b�.�0k���!��$V~��!�h�&���ˁN�Iw� ���˺r3B}x�
%s	K��x�{�D(2�kMq�P�2r��:��<M�왻�v��'��x昻J��� �C�Ҟ+;)��-��$fҺ������ovv@���p'4"���Wn6+c1�+�i Y��<�{�	�����2�Ǽ-8�:|{��W	��;ݚ�cP�ϖw,`v]�-+p֓���]�,Mj�I˸,�R�l|v���\t��WR���G��&�g��r$+�)�7to]��7w�\7k��۽M+:�����$���	^���a,:O���|���p.��(ԧ����vM|Q�ݪ�1��k(m��|�1��j�����r��`*��ZýuZ��w���ۻ�e��b����6B�:�%�SN@%&.[��6����}��3KKOd�u�ˈn�S�4ۓ�G7)뽻Hy\���M-�$�1��t��{�if�~u1�]�c�L��G,��k�É�;��lL��<�y�'��"熞���/u��ݟҴ0h3�ST!+�:~Q��n3�lLm�����p#�]���w��l!�����D����c�東�E�ϲt���.�5ѓ�(w(�m�\��;�ˠ�RB� V��zƦ�'n$S�W����6�:����Ǻ�{i�_o̒1�3��.�Ӗ:�xln����nwp)�
\��*�kB��L�\�{GV�����t;��s�=�&�\�=n�fh�F�}���� mM�9�'	�,G������J����v�Ϟ�5��l�a���Q gn��'��a�]����9�Im}kJ�ڮwR��K���
\��Mk�C��X�r;7倖N#����9���[��9�FK��F}����Ǖ��xe	d��ʆh�d\�X���b��q�[1*��Hp]Z���$� =ᛊ�C8���N�9h|y��
&�{�<��D��q��E��9����6(��zSCn�����x?��>݀v+�^�����m �@mM�ٍ9����Wj1�a����)�X��U2yw[h��j�|d׶v���7u�G�3� ����n�e�0��[@�;@˷*�c�7�&b��d3�d�1��=�\`�/-�\|^�ah�۳E�pC�hODӏ�C&<����[4BI�D�{��N�M�F�3�j�	0���6�3�?�l�����&d��kFG�n���Jj�>�H=�$� �#_��3�,=czŜ�f���_�ԖF�lm�T��L��w{e+r�õo^�Ơ�>�S�rvt/f���p�����8;;xB��Z��zkX�Q�� �j�vl��϶i��ë�A[�0����tj�������q�����, ,y'H^�n�^r{�j=Zy�i3��{�8����DL;{筻'v��-�M��:w�rp�5w��p�z�,!�݂�ه�1\��ǰ<k#�wm$��gmc��ꏸ�cBX;�-+.!ٯ��٤��`�[�8��|��&�1+��M
�p����v���S�$���q��N�*(<
q��ů��6�d莞z�I�a�w�����w���p��xz��[d�.�ۅ̙iYȾv�of���-B�,���\�]�qK�@�=qf�e�QQ,�.�Hx��9��=�-4���p�:�4�ޙtsar��<�j]���^��Z#�L\בQϟb���l��n2��;�܃pD)���j�>����[�4��ơ���c���T)��6�V,W�<���7�98�:t���0_S���A"��گh�5C[�ʚ[�+ӱ��<yw^ըn�0�r��eM�	$�,�7=���㈼�Ay�8��E"��^]� ��v`���/�P��O+�jƚ����O$F�!iS^%σ�����?�/9�a9Vxw�φk��S,
Mt:n��c��Փ\�vp?Mq���<PO�њ���G�1.)a�oa]ݐ�n.���z�l0�f�(���O�o�>��\B۠`��@34N^gb�zWvHq�5�;M'��l�_hR�cŽ��R")���͸�qs��>�c�;F�Nsh�X0��� �N���Y1�ɜCOh�.�͢	����o����#x����{$~>�3ďL&������� ���Щ?������	~��wdq��%Ox�6�S�E=����̺oO`��'�P���&/7	���v����%�x�3Jfx���4�Yx8�Ө��F�	=��#	d��N錌DO;6�ig�R��0��i^n�-lOnܑn�k]X�$��'gg?�f��	t�}���U����$h�[J%�Y�Z=R��x�,��x�-��"����}d���F���'<5RlŉC��"�F露�R
x���G���o�,������O�Q��v���=O3F6{K%°k?����L�>Ӵ�,���N���t�|��)_*�%.��olݣ^��N�fS�5g��z�⯶ˤi��yQ���R��%�izv��gĭ;��$�<I��[+���z�I�	�Z;�ad���p�=�0z���v�l-�I�t�I;�`�F�bl_or�:�dM&?�X����g������׾���}3�{�=���m��m��m��m������qE�S{6��Ƿ�0(7���\���}|��B-�~����m8g��jj]���9vxq�����љ��;K\��7z�V��Y�јfe�'f��qWE	��9�r�r��C�����6������ ��|���%�@�/�P��|�n�Yf,X��>7@Up� )��˝�g�x�� �,7��wR������۲{(�^�Wzq�w����E-=��}�ٰan����{M���� e+�c�Y#ӽ�Ǳ�h�l��|�A/+�����H�hnrH��Gu��Ub�S=���7��F1�r�7�oyvΚ�{!��c\�#���c&wt�jaa�_wlҽ��`yNuj�uҧk����7������
��ǂ§�B�Xv^M^�X�)"&�^�	eh7f��r4�������V�ځ�8)m������C�V�IX��a���0�z ԡ���f)ق�97�$E7����O[�{��"�}�޳� �%˻��5��՝�w���!�RFN�zœwe1�o�r� Ho{�^�۞���M�G�3�k~	l�%4Xli��,#j6��u@H�U/Տ.de{�c��gn��M��F�� a6T=��i�(�.L�Ĭt��a�bbc�ww���P�^�����ޞ�ȹ�4�D��o��{�����"d��AعV\�3�jAPJeF����U�{��
y�R�X)���5*���|=�����LY�HJolՓ��y&II�bø)�"�F�&T���_b��h���K��sی�5�a��z��{,�����y�e�2�-xa�}l��kVKw4�Z��lf�ՎecD�l�7�Y��	��,^]�Fxe�	�<���%ǾRx��*�w��	��5࢏V��Q�,����DD���݉L�#�,w�\/w���;M��d\4�Kx�bRL�fCZ1����.f��Vq��hګU�@��Ua����6- (�4�ON��I���GM�/�w�BZkW�8z1�~˪
4����0�c&�ʹ� �ġN�Ec6iF����������/��e�W�B���/��;�F2����glk��7�{�FV@np���3}�d�?>�<�l�%\�W\;�"E��V�\y�L�r凖[r��s�Z:�U�;����G���!���]����j�,k<����D��u��ʾ�u/tOnI�l���(e$�E�ѷ1w!*�/�v�v�k�`���R\l�C^�;�Ӌ���5�)���)���X$T���w�p�Bӥ9|�f��v�(�U��ꙃF�T4�C�V��Y{�-�Ţ%��~Y��\���.5[�,�5�.�Ͻ�=�����"�^�Č�*��
��L���j��2�w\���ך�TH�$�]�Y�Qj���.�ьJ�˻�&��3CI�.�ʱD�Z{Jt��gOK7����{��y�ꇻv�G!��y�}���k]���>����Ӆ*n�tS߷�Mi6��PW��¯!�"�0[�\5�k��iU�B�]Ť��N�{e�w���ui�u��ˍ�v���|Y�X��{D.��'Iu�@h/bsd��G��೯(i;+���؝C)Zd���n��K;��.R���;/�$�03kh�����r����9�� ���27%�:ގ�X��L�fn/-
�f�TSFt�E�Z|�(a��8�c	g��]�t�U�h�qj��0LKv
SsÜ�M���i~�X}�z*����)}A�0�h��^嗸��i�$�3&�aח�����]� �D8bS��<^�|�;ڑ��6`L=���*������9�z�Y'|`Ǽ}��I3|V([8(	@p_l+��� H��z��o��Q�����2�04i��3�/j귬�e�7��>ӣ�A�=�`¹r#��o��H;�'��Gݹ*[��V5<�Wxz��^\���魥�T�jw�ld"aXw6�/@8 n������45�	83Qk �/01S&�W@}*�@��֡���5	W�;[���3	��Aٻ*YíVA���]˺Iܙ&�\E���b��7x8�p_#�����'0-�SK[[��ڡt�)�l1Y���SگlEǾMr���D�K��M�j���c5OF�\�	յ��G^o��	�^���QӢ�i���%Β���jw�0�v��3&�:N��
"�7��;��r��0�J�R������ҳ�cyk�|}���d�ʰZ���@�P~�~���^�͆�_l� 7�^	���u��v�^5��<}|N���uN+��8M��� ��8�U2���̉��m���3��KtY�_�!:�����feEyݡ�l3� �R���(#˶>uN���-�y�r�-b�G���3��e����CT���}��� �J��9U��p�v����;�}�ދ�&�{�8Ů,�#��w�t=qcѿ������˺"��ߥ�B	t�&[Z�w$��2���k)�e��u�����фE}�'|�YEc� ��n��=��"I�@���X�T]�n���-k�dԘg'��T�T]���X����cӗ����;{��r�c���'r���B�o�b�y}�ˊޏ}5��~��U@Jv�l:z,��x��Jp�*�B2��Ƥ�ky��)*�戫0f��I~av�K�9Vo�
΁�61;Ou�d���(�J�\�Z�+�ex��g.���=8���糔��02 P���鶎N�P�^Sm�<���ּ���ϘǺn9V{M�����F�^���3i��\�w�@[���%��b
��ifC���ѱ�>��/���I�+��.�<6^+��ٱl�Ʊ�j���X�)F[1pq������~�QW���ɷ�M����#Z�s��=Ox��r��C��xn��aɀt�7�oh9d}�p`|�xT���b���܄�&M�;�z [��Şc��o�`�9���b6]��d���gwpE|�l��-�� �ks�����3��T����ػ������tg��V��oV=*�/��U�8\)�(}�H�LeM�Ė� .%3��X����M�ܴ��ܳZnwA����xm
��9�(��Y��VQ����[�o.p`F��$��m���E����}��"hQ��qk<~�v��<�=����3�{k�t���.�zv���w;����=��8JX5G�9N7<<�v6��÷w9E:�^��ᚌ��Dm�Y�ku���� {5�".8[�.gT����4�TYKAs�m��9�N��H����3�3{��p�.$,K�Ю����(�j-��+_fL��Bs�p�Պd���!�-�#.�˰ڈ(�E�,%ds�V}�.ܹd��9�w5�N�|:{֬��y�gvV68Y
D�P�/15�J�Pa�کw�)����lfe�Y�M(���k��xS� �F���{��׳��PГ��n��!��p�)�
��`�:��EE�	^W8b���;���*�fs^���r�@xJ��G��5������!�TK0�Y�w7'*��X^�P��AܴZ�Zۦ�R��K���[�0$�q����)�jėew'�{��(�7��3좕�1����^N�#f�jV,��ߩ#}ؗ[%���p3Sӈr4�$�a.�����(�n������N�ܰ�}�i�b������C���c+ؽ�wo\��scׅ���!ev�,x�Q�d4���o��HV5O�G?��k3(�H�+��i}$�i�TD|pa]`��p���㽿�75ۛ�b=�s����oD�v�6��ś��.���CެU+>}�h�Y=0��w�����ׁ��/K#{ک<SW�1����v8�u��Y�%�-��p��Se������"s���ד.��a$�cK2�W���j�
׌�^Ԋ绉/q�8�\RE|�`�l3|���þ�æ���a�{��/ݳz:�p���m}����w�؏	�8b�J�<@��J�E��*��!i��TL� �ŶO�#��!��ި=�ۥ���e�N^�"'~˔��P�R�kA�ɲ��ެ�mn�����B�1������(�&��f���TXSj.v�0ڸ�\A�v�r���ې_>G#CPmG����P�����P�M�{��U��p�[rw#N
�Y
_�9�,�X��37�ɳ�.�ݾ ��<��Q���$�s�E��eY�Y&ܠ\���zt�����<~θ��i��2f�)�a���	��g�����O�)ݷ�&^�c�je4��siL�ӛ����N�d�>��u��n�4�('q��4�����RH܌r�{�Bz��_�V5��F��Y��fi7q�d�RV�=ޞ� r���@=�M��?U�K5	B�����t����5$-�[�ҕ���R�e˜������Z6zg4��7ԣ�ɾ���~\<�q��-%�'N��~��]ì��Q�t�W���(�l�B\�3H���H�5�,,�"��_#Hn�T�!)�t��~͹�'�h��)۝�<_��q!�N�uܴ�L ��<����Ǻ2\��W�໽�饌�*�]vV�`��YN��燺����(��hYj3JJV�lVfɈҠ:��o�b������u-F��T]ŪJ��,��.{s��g��is��-�M)f��:#o�R'g��������gC�H�C��|�ɕN^�ُJ]o���do�t�D�?������|:a��}�oD�|�#8��>��yD�7�T�na�FU_P�Ûm�&�y(�m�K��e�>g��$}��3��C�=j��kܷQ�K1L�M����Ɠ��)�����y�nP����X� !Qxk0z�'�����,~���o��g	t�蠙Pt�dz�x��L^���caeۣ���} ���m �sK�xo�gM�u/��oX�ef��[����=���RL�P�<�ѽxU�O�����.�h���B� rƁBfFf���E\� �A�;w���w<�^�g�6��6����\NI�!��Hڥ긢�5!*uR��K�DC�K��ǺxT�غUx�	�>�c���}t]�4�)}G�C�x�)��~�	Gp�3���1�/�f�޽��y{���Q�`�����~3���V�2�"��I����L`�����3�v:'��5{Y�n�x�=d�f{7 ]� ����u�&v�^�%�[�n��qݺ�~^�v�����E��ox]W�������G���O��.k��1Z�t\G2ᆔ��VU�]Q8���w�j��:i7��֊ �{&{^��ٜ�r��621�޴�e�n�^p���uJ������S�wwM�tv3�6����-�{;����yvm(�m;gN�,��L�*]��8a��f�ӽ�nh~	�%���VS�4;Oq�ꩭ�sY:����ML��vj��Z�s���5� �.M;l-O��0��䳬�4p��g�����za��8wJ��z?V����7�}O��`E�y�V���D�3�D�:f^͘dֽ���sh���Qy��7�+D{Y/�ݼntp��p�]X�:�ƤZ�(�d���Y.,m���=������1�=�܌�cۺj�J�r ������rөy���4� Is+'vZ���'�goX�Q�uX�w��9u]�Z���n�L>�1��6�I`�H{��r�m��QʭB]��EY� �jpΒ�6�N�����`�V�GM������{E��	5���Oo7��6Z���8c�	OF���<�^3=L7Z���<sV���/;��a�D�+���kӳۭu<����Bj��K�*�9,U������zl��5����۸<s�S���q���qVyu�RMs��0g�p��o�=����5s�4}��*Ov�����qY����B�BY�g9���U���m���-\X��&ܭ�����u�����ꃐ/��=Z����f&�YN&�C[Ӳ��fc
��噘���"�2��*�Ӵp��sT�7�W.��z��`=	�{�Ő���u5�;]f�x��܀*��b�Λ��j�Fl�8�T�8�8ګTf̖��i�ː��t�7)��# ��	LUe @N.2��B�=�+	"�kCrUm�Q����R�M\hzi��ʙ�1����%��Э/���V[������8ٚ�g�M����
gt��n�=��cC�x���<�Lb܊ŗS9��Ph8S�P�&5N��{�8R��_8k���c�����ys��:��lX�S���۷j12>$5J��z���37���d��g�Fi۵���zu���5b�7���͠]�v�~X�Ϲt~�;rO,"�y�6`1�͸�.Q��\���%�"P�@��'y�{���������h_p�^ܗ�0�!ƹ7��y��w5���u0sPN��oq���t�Y���n I̜�pbj�&�ĠZm?��2`�Y�6�x�-���M��m��m��m��m��m��m��m��m��m�ږ��
[qF@�&Zj�����X�#t&�m��u�"���6b>���R{��tԍ�z���u��W��P�W����}��^�:�=�>JJh�O^���4 ��RQܺ� z��k�G���@}B���hOp?.��4:O���I쏨Opy!�����߮�%��@�O��/˰@�y�_����'�?#��q�!G�?���������������W����of����W��s�vL����j�4RXW�r�J����t}xT�̕y�'7���8��%�[Mʡa3 ).œ�"��I��P�M���N�cv���ol ��``�B��C��i�L>_,���j�oE�!V��S7�V��XF��w hԏ���7�t���۔{eR���jw�i����m�E8�<�
��<�Š/����:�yv��J�{�������׽��c{���<��x|�Q���򵩸V�^V��+Ƌ����[9��=P�|�{��;�R���6�l�ԕc��Y�4�z����.��$u ��nj��"�WL7�x���SYb�#V�+����N���^���J��3�MX�u9�È#�M�X���]�M�+�0��u�-᝙ި�,7l�5婝����E¸{GeW���[���'ph��fq��搚��c�҅�60��BQ�e��[S�4���4�7�"�m=pYf7䜣�Km�Rf�{�����oD����k���H�Il�VY�ȹmĿ�v�K�a#��}�P��x�=����_hm}ҭި��{9v*j�� �0~)7l,+Q�l�EklC25�Vr� ����;��+6�A6$��ᬷ�^�θ(ٽ��9�<�ۮ���S�&���N����{�zr�����~j2V��ѷl89xA�Y�;ڕ�D3�n��ӸC���x��п/�vg4�Q��׷ݠ��}���� D�mzW��%OC�.��h�> mm��8{z�@:�1@z�0���\<7ʗ��6fG޾��E��xK�*�%�T�k�n�51=b��Ӳp�6�>R80M���.�%��1��+,��$��z����\��n��,I����-��2�������R�S:�
��հ����x��zLU�:hh-�w��9�5]��l�͐�ʁ�5X���k
�o�h�dٛ;$��k�9k������'t��/Ԟ(��8���6��Rk0�v���T̷e�n��M1���;�Њ���?_��{�c�����.�9O&M���ɬ; 6��Vf�y�wQ�o)������\�}�����r��<�7Kp����	@CtF��9�d�����M��L��1�;,�3r�
w�;&��ə[Q髻V����_����;��Sx͗�������ox����{��� �mp���ǖ�m�g��x,{��
�χwx^�VV�͉���szs�,m�&(՞�v��c_����!j��҉��()dC9�nn���� ��"��˙�Ej]jH��@�F���g�={��*�!M�Q��z�SW	Ɏg#>��r}<T�sj�q$.����r�h�s��l���3��;��<O���n��e·V_B��[k�x��s�X�sl�xmX"�ٍ��	n�f�٤��4��<�7b�`T��{�빡��<|�W��-E�7��OG��_o:��'oEѵ`����.k[x�����'�v�أ�6�{wY1*!��;���L麁C�v�VP^{��ٖW�L��W��nw*A����v��o�:J��Һ�{�]�{wD�{u,՞��r�+VK�hX4ǥ����2�<>��n߸�����Nį��Ny%�,lx�4e���nۨ�S�����Uk��w�B���%E�N`Az��/&F��gF�������V�j�^S��F����ؚ�qv��8,S��bT(������L���W0`���꽠�w+���`����^�Y��L�˰�Rm`�Q������)��n{h8&�l�թ3Z5����Һ��$;n[���ԹA�g%G�'�d�{�yFO��F7�8����1�TfMh�[�U��;�~��}O����Q۸�#~��>pf73�GQ{on�йA!Yal�R�.��z���ڰ�FzS�ӱKx�uسa�D��T��:����{Iѧ�o�8Mݳ����Jaz#<�]�]��6yg�vF���"sE^����\to;��Ϳh�N��R��eb��J�$�����&qV�����W�ʆ`����^�-�n��������U���ېM�@�0	D�-��ڦ��eиC���Ƞ���|��~���1$�T:F1�swއ�,鳍��[}��U2hy�}�� ���=F�X�H�7�"s��O=�%�ό���DG����j���];��i|S?yX>��Z��Q��~�~G~�o���mO����pJS۞v��z7��w�\&�gvl7e9'��?Y���~���>&v�]� ����9��;y�-�	��7j�/���{X7��,��X���t�R�v�bX���׌i�5�=���2��^�\M�eN��m�݈�.R����M�zJ��ty'��w}]~���C��z	��5���
�@�q�� L�8�Ð�g�G��_wv�E�i>���w,��`�����~}(���J��n�MY�e�m����uG��[I����:�����=���i��|;0���>��Zd��U�kv���e�{���7������|�ek0��iu���,��DĘt5Z
��1��y_\t���ލ�by��ޫʰ�i��%0�i��=����ۼǆU���ޮ���V�j!�+�����(C��'4$�~H�����F�h���/2���^G��9���U�r5��I�8�^�y���ߗ�����o�c��l �٪��~͊�<y��s�l��1�P����Np%پs��{#��sȞ�ޙ��
<�g[��or�P͓�c��=�e�%s"��d5{	oe�z��~�8D�8N��5#q5�!�3'��&���l�;d�^� �c}�vk�N�Ş��qK��i+�Q�	����a���*ܡ%EO�{F��p�����(q
��"2�b���gs��84�vfѨ�R6��OW�����>F%���n�-��7�N�^�'��wlc�����֋�K7Mi�^DDɾ��Q������������LG%NtD�R���fo�t�d�soQ�3yQ�f�Z��R�8y ى��wE���̱�-� ��`9�9�}|�H�`�^��rNR
�\�qM�E������l��zԼ���θ��g/p�¤Tj�AzD3�}8dB��8�9u�~(u�theŶ�������-)J��&����?����k&���}/>S�y٦�M9y�9|{^j���3�u�@���z�V�*���{y��Ӣ(L�!��𳭯}� ��(��r��ۓF�z�12gax�d�:""}��I�gD��l�k��:�L3rË7W�v�pyu��������,UXA���y�Q��zð�
���2ns�֧�.�Y�qa{)�9�9�@F�<��>n;|����]�/9��m �
s�1*R&U^�n��2���0��Q�{X�y�.F��v��w�7Zˣt�0��w l-2��U�?%��y\)$U]�7��y���6VO<�����Z=n���}W�|���+
��s.*��Q3���$D����@]���@��t���Y}8��\_ng��2��b��n�V���: [�1���w������@�_nG�YF��83�ؠH��흖�xm9����鹲?P'>�1�\����X�1�b�@���H�݆�Y�(�Ѹ���������="9|"��&ٶ{������ޞ���[)[U�{��o���[��X��x��Vf_-б������S�|��eq�"��dΦ�~��sd�` |s��re�T1z��ޒ��f��4�}2�����m��6(+D�b٫"�U�ңH�X�f����D�b67Vkh�ޥO�P	��f�-W�n r���lҽnL��}<�AO5��Y+��f<�+q����g{[�{�A�8vet��p��G��uL<�EkRAd��XF��� Δx��p9�t�5O�lԾ��g�����u���3f�� �U���5��_dr��V�Ӗ'�\L��.�����FK�n�����=����uv�w[��Wk�<Z&�==����h>�����c:Z�8N�ݥ�޹�%b�0 Q�~�׊��`z�O���P^�Y�<��;<U}�Z�K��^EYK9^zpcI���1���{�K��e�g_{���gC�\��w�T}/(�A�Vt:6QϺ��<=׏�j���E�(��9����˽`șz.j�t�a�}꺗���\�z�Y������f@��k��3w���d��7�t�e�Xb���6휮�vI�G�F�p���j��J�$^��8�A�lms��ὦs�}�?O9x,O�7K+r��=�U��+���=����W��;F�#Z��!Ɗ2Tv�%5%�=����R{$	%M���cp<�=y�-�+�3**[܃0���b[�Z�`��=(y2���3;��9�"��h��^]�b�=ű6��MJ���<�c<�{�q��}��ɚ�6%u�%�P�
`ЍC.�S�E�>�ŭ!���2�/Y�`�rH��	����We�˰��_s��f��؟F�`ּQU�i�0BU���VAU�ƝcV��\��t���pc9�L;�rhͺ��R�1�wz{+�K�Sx�6o1���]A&h��t]���w��s�^d�uy�[�zQ#�B����dʔ�����Ӂc�= X]�F!� ���;;v����n�Ue�J���ŭ�hl��)���^S;T���Y|���,�ȷ�0Lb��b��[wդ:l�.���ē�`jJ��.�	fu]-�/�D\��N��	�����	��N���.�)F��_�/1-�Q܂�v��F�(w;�I烉�Qc;Nj�"O&���Ok(kέÓ�bY����Ly�J{���h�]zܘ`�]�۷m�쳴�(}h�͜<�p���N�	��������B��͛���K+0[��]�F Y�`����@VN�lsF��"��p\4�̪Ql#P��
���{���Su7e\��`M��u�����D.Ⅲ�J�����>~����-ۂw�(���Nd�\�����G{沍�!��KJ���L���/pt]�K;��B@VM�*��i�b2b>G}��[����H7 ~�K�ᤄ��}ÂQ5&�_@��ҙ�8��4���h����� �׳C��k=)�a�X��v�}|p����{�Z���^�Ca������ �t�	���{@��{�kM䩀jC�ԥi�⢂�������&�RjGD�ӕ�Q��3s�IV�ǝwv��]�3He���*̇h%6�)��,"�+(��J���m�ޒ0��m�<|/���Cs��{� ���+L�U�2ݧ{�Y/6�-u���:�_!sE�����"-�����/{:>;�8���l�l_dP�C�����so=�2��R5B�1�y��u����wwo���VVn�rT�Z�5��~4g�!T��9�ٻw�I�r�$kފ�|�}���A�K��A���7����m�M�s�V��=�F���[�1^WB�)����j�V8�\��O�dM�p�О8�KT�/<Zèγ���cE{<�6�''���"�M��J�����:({��R��.�R�Ϭ�:ƶ� q(���NS��ǜ:.x={�&^�r���G0o�m�_t� �X����7���}�JO���=Q���Ƈ�{/�N+�K�}S�jOc"��^��9������{�X�H6{J���c �K���ձ�I����7v}����;�W�=ñ��[�x�k��G���Y8
"!�s<�]�m�F��y�q���zK}����L `ʣ
$�Nڤ�u�Q���ޣrJ]B���}�o�נQ����"����
�Q��3�%��Z�F>ի1����-�ꓪ*;w�0���C�_�����K�R!_=��Wx�f�8�Ck`�B�wnV�h���'yYڵ%�V����M�_��P�4��>,�h��������.3�b��Q�x%-P�y�֊��y*���:��NOgW��s+ǠǬvzW��p�f��X��/w7"�9;��[9�I���-���j��z�@g��^�������U]5��	� ���4�~�2��_����g]^mJ,*�c��0V����.e⡷�i��-^����Iޣ!a��?l�s��a{&�M�+�S�Z2��M��S�j���؏��&;D[	����״��{�ܛBƚ�$G�>�ţ&��:}��`~�M~��5ƺ��Ӻ���� ���ql�K%���2�v��,�*��[	1���1fl6Uv�h��M�����U1��/g�qn#����R�=��cM��9ۋ�;�<z���i>�v��Ov?��/���l<��س�O��f��X�@���po��+����B�ɡFu+#E�0q;���F�ܷ*��z�N>�A~ؕ(���#=�k�5�{��lX��Spf9�c�<�`xc?nO!�����= ��x.|=������"�7k=��杠�lHԕ�����sN�sy�Z �C.;�*��ۅ��ua��;��������L���J����#�t�Z8`䒳�<ρ�;�9y���c�Ǧ��~�����K��h�Np��ҭPy)�ٮ��ǻ��L�d���e�=����G
�k�D�[y-�s۞R�����+x'^7����WY����>���K�]��!V.�oI���.<o��C/;�a^��A.D-c�<�����Q U��?��?������ҿ�~O�'�����������Ϗ���������������NNNNo3���?N��p�EHD�!p��P�D�F�hR`�T2	��6�4�F9����0b8c��h�b�� ���kJb±!^ �#P	R�"�I��MF�K�2�H�H ��LDbH>�*#���3r�i�����;R�WwM��z��{Km�	���'��W���~�{l�'��a���*�,�Yĉ�o���~�W.VWV�r��$[1ztJ��u���=����\�.�#K���J�h�׸٨-�kN�۸f$�a)d�����u�lw��}�iS����e��֏�r���|�ڇͮ<]p���}��qg'���q /��o�Rw�a5��>h���QXlhx}�@OVe����U\R��o�Z��A�ϭs�n���F�������a�IsY��$7i�b����/.ͼ k��q�e)Y�2�M1r�5����,�͏��v�#�jW$z��н�&J��x��g�x�m��Cٸ0*�Ų �p�Ɣ2�:�N.��*e;����n��{LZ2S4���نR�j¯+1�Je�Ǜ���]���Ud����MV��T�,T�����}�G�ݥ����25��(�/ahQ��zQ�1zI�پǚ�ޤ��� �p�� �UH���H�={�7cL	���iv�y��=�zJ��s���{���W��'y/
���0�ƾ��]�0�����P��)�w�ҷ�����~'t)���-���\]����B���`�5�������:�V�T��TfȭR&�C2Z�h�۩Է6-f��\���ܼ�������Q���.�iFI����(\M��!��hEA�])3
P'
!�$���IȜ�@��I06�B T�L��@�D'�,ĸ�e@!���D"�N��iđ�4P��d�B�-��l@�2D��2�F J�@��Q�HK��.�l�D��<-4��Q)9	�� ���9I�0�!�,��1�@S��m�JM��Z��SD(� �	i�I!$E�D�N8�q4�\��g���
J�Z�,�'u�s�OQ����뮺��7Y�I��&�u�tg��M�SE4��@]c�thbz���:��M��:�������g�����XԔ�PbPu/_6:�j*)���m�U�h-d������g�1i��z���CD���w�[4����)�����z�B�tcB�GS���
}l�A�F����h��A����SER�:N�:���N�QUEPSES2D�U��"��M�߾��bѓM���HS]u���:�F�v�l��N��GX�覊(��-�Pj�(hbfm�V����i��"�CUOW]d����Q]cW{Rh;��S]I��:(���fh���PQUԚ�`�Q3.ت-��詚��l���T�[CF�TAE�����!�*�*+[׮��`�H$�I"�3��F&:L�i ��$�% RF2W�v��h��9
f�b&񐴉zVQ�C<m�%�{<3�u���J���qy��!�E�U�%��;�Vk]Z����`�Ȑ1���D��)$@�8��0�"KF@Ap�	�DA����A� ��Q�����7|���zho	�����^�5�r5�y��X��U�@��<�Y5��k�t�Ot���\�5�Ul_ɂ����J��ܻ7�us�0�83j�R��0�j+;kN��eR���F����b�G����h�,I��|�DU�{"y�s�.��5���D�\m�.Dp1���+z�G9�s0�n5�]d�;�I�Ĺ�ȕ�"wk��w,�
�	�ϣS�@R�3.5P�Ĭ��.��s������������WG@�Q�"�k팾��s�N���k)��>�-3n='I�'K����k�q���A=X����ԛ�t\E�v��o���$�c�|��LQ�uq��Pwq����bi}�1���F�qv�6�os{�8T,����{�u�-��q��v��1~r+���`8�9���OQ}�<��>�g�C���W���[@�t՝�m�}�{[S�묾H�Vޘ��7;/�}Ha������4�v���M�f�c/0(Mڄ�6f��`��+�Ype$͍ɊDhf�I\$�h�Y��qrݛ�Vچ�\ir�N9I�X3z�j�#I	㙛[����i�ѤAǱ4�Ĩs_�qVC߮8���<��ӹ�2������fi�F�G>O\LNɍg��\�t:��_k߬���AS���l����ݕcRo�>,n_7Eq����Ӷ%���;s��:��cը�QW5�p�t{y��<����GE�jk>}����i��W��Y��8�&1Z����+d��K�_p���Mzf:F\T��FP� ȣD���u	�3Sn�I���e7�.����"�v�[�i�oY5��m~  ���]�ͬμK3u�]�E�sv�����sf U8��1`E1s'��\�J����B�yr�����JV�����[&&�%�u�8d�0:؇ʈ�s�[�-��X{�u�-=�_w��>V�wv����T8ۮ�58�^۞-�97�?S��m,}�"^s�+;8����$�ӵ�?�y/��`r�
�Y�8ܚ߹o���ün��'<վ�P��4��(�L�7&�VE�ɦ�p�4N*��{�hx/%�<_������a��^�r+�
oU�9�*;o0�3teP������D�;5�%�����䪓G2�d�Ψge�x<��̻%��Bn�����j����v�	���˩g<HU�-�B8�;W2���=�t+���Aŋ~
~��;�z��ܔE�x�%����-�&L�F\�#5��	\Try}�*WjR�_%ܮ�{�݃f�vf�lSE��z�"������UН�ypE����\Zب��|����96N�h���#�!�0}�Et9�'�ޙ��vHm���.+0l���>�e�G���vD�SP��B������-uE놣O8U�U���M(J
�vh��_3t�ͱ[�-F�$�X�O˩���Н��E(�5˕�u�� ��7�z1s����@D'<u�0v�oj�l��=3���5;^��"@�!�;��n3w��:A��-�c϶�pG,�g0fz���,6����/2f~�?:�9y�opq���������ثv��Ѧ�V�Kw#qH�N)v65(�����S]���Ő0��'��F���0�D��1��"�Y��}����[(k$�1�L�e�gb�RnX(M��K
���N/#1��߷o�`�kᰦf7Y`���֡����C����Z ^SlLtv�ű�v��Srf$��O�4�oh6�k�tq��`s��&d���s>���H�0r6i���X��:�&�Q11��/�%F����؉w�~�w��۴�]��S�p�=gG:y�x�n�r���aR��{��/�lJ�ϻ�c/7����$��N�/�m\1]�8�n��Aա��y�}ς�?o�Әgr�=�Q�kJ�LmC�7NϢ�,x���<�Z�x,ɝX�p�3!.��qf7��sx���LQ>bc��c��1,�3�T(�\����)���>y��i���^�QLT(�q��G�+Vae�Up����.�`tZ�k؊n �t>\�wa����ű*�D+��&H���D�x��q�U}<�BӼ���`�n,�7k|>��<S`ak��,��'���>����(X�:�&�RoP����y�.�����no��4|9�e_\Ա�8Md-��1�f[��NYK��K)\�^躷��\�W3�Py7�ꊗ�H&�����۱�ޱ-7z_z6�h�%�
��&�T�hnl51S[L��{�o�L�E�/�}�`!���'@2B�73KE���6/Q��<�NA��moA=��3�"����tcY�*�e��F�v��
9NpJ��7a���68�	��c{>W��<�!�F�=��������1���m�kݭ���4�4D�<+$߶)�쵎�P&a���`�ufnͨ\O#%�L���^<(備����|{����m�<��`ݎ=�+2z��Y���=C똱ú�#���{�:��2�մX1n��Gs����sF۶+�/�\�WG=�|��"]���iO3��p�f̍��}"��T�'��G�p�V��F�n��O�+���/8�n�u���=�9q��[!��pkۮ `�'o��c�mH�yQ=y�U�:y-vՆ��<wٯ�_.*�7�>;��6�r���5U�6U���d��"�%�Pή':J[׹�R�܀F�D�7WAM�5�̆V�����{Wm��Vb�e���վǄ�����}���|�a�)�L�{C��	�;h�s%V����K�����T�=��7&�Ќ���D��0
V�!C��\(�yY� ؖ�凹�v��̆9_�䣹��]K:摓�b��\��ñ:�s�yԣ�]��X�G�;���܎Գ�|���rw��S�K����1U����'�/~�=�Lmr�o1���;�Z8�D���z�2w�k�M��`F���oC�,2�oh�}'���oz�Z:��ЂbZU}��!�bb�P�s�!���ͥ]��[��ͫ�#y.�o�Vq8G��c^Bؗh}�������j�c�z�hK��O����Ҽ�u����s��N'���3�B�zփ�A�n�w5Ԩ��WEmDp�z7���:/So��D.wUQ�{!^�n�a�\.ǻ�v�廨���h9>{�왍�֊���^��
4d�d�.kal���zzWX1wѹ�r!W���b�����l�C��6}�Ao?L���	�ߡ�3���-�2� {�B�!��_��=���*�gg����v�ͧl)�v�j0/b�eE��*�YG�L�L�/[��lL����-S��V�2��a�Ln����#�J���Iƒ:^�f����L`�@�(�Ƭa��4�$*�A]9��1�tmK�E�r��}SNdU��A���°׋�7�p�ZS�h�u7Dd�`����nC�巿[�|o�n� 2�͝�c���B/3.��l(������*:��I�����j�oe�����.N��}[�  {�8]��ྩ��"��"^s�+;#�Y�y$�o�U[L��pS��&7���	ь����=6�+������]O���J�-<�X����q�S�0��� �m��c	}r�L���U����[�k.R=gZ8Ki����'/��Ƞr���a
����I��Hl�;��'!N�+E�,�!�����`y�3������<���&1 �.l����}���Q	�Nшgb�D��SN9���9�Պ"p��r��o��c��]�c��Cp�t�5���R~ϻ�pR�ɉuu"�vμ����Q�KH|�=��S�Ae�5o_UZ���
�*��IZ+T��|�V���N�e���0�,����&�wH���+ o3���č�����"�AډP�*�䐨�uƶ��ɕfP��)�u�*(�	)㯣g��vk��%
�9
��q�ô���Ƴ�Ekʻ�����{��n��\�Etj���ZXJ�\V4�c��|s���`����PҞ�b���������>95�����T�����N���(�(jn��].�Ҵ�D>�9�/�����ɨ�`Gp�3>���*��ur�6��t�{��r���7��;���D@�[߄t��nFō�0gAUQ���L�A�U(��\ؤ�Ҝq��b<��=?n��f�dh��i� �0��iT��3U5�Ar:}�=��"�춒j����k����
D\TN;�bt�Tͬ�g�:���~2*�����$�q�^m���[���f�|��i�r4��q��]8�N�}� ��}���ۚ��tgu,61w���tZ�b%J�r:8�8K.�d,x���/(ҁ�a�6��=4���C
2�Oa5<s�<{���(�Pg`�0����N��� ��O)X鼚�76'VV�g
]�?�ϳ{���fA��M����:��4}�+��K���tĳS�uJq���黶�bPN��	�H�|��^���/4���y�b���n�zz,_<�z0S����.g�LO��ޚ'�F�h�v춸/!�x��N�4��SY�'��m���Y��7��=&�zh� �(�׽,:�>�����H����j�D"83	tTovYv9c�i��q؇���+g`�-�U@�|�LI�}�[���'�����������qg��)FuGLu�Qޭ�k��W@Xn;�q�����M�7n����{e�8)���A�9��1�!l�����w���I��|�VV*�#�|��e7Zֻ�4��H����Iח�c���=�5U9wV��{�y)�NlX�3R�����"t��VQ�y�)�t��3�ۦ�4J�Y.*�L�\�C����}M����-��{s�����wk;�Ί���9'E�J�:Y����p�ߢ���_xO�Wq2=G��Pz齞���اv���yE��?3|z��� Of�3�B�wp�Ɵ�Q�x�̐����o�4�d�-��5+P�i'7��Bvs�����R!�!8q{���yh���8��T�v���e\5t�X�;�l��nL��P���jFcݠ�n�f-[Gg�g�r[��kw�t�>Qƙ��ٵ@פ��"+[�"�춐z������|��0���=5�x��C*��Q�@ω�4M\/�u�u�ϵC�N��{7��i��U��dM�����"VvwwH���Ns.���#��7%��$R�Nq��q����j��J��&�����ʈ��Y�r��V�p�w(������4K�MY-2:�D�����G.��u�2G-��6��W,c�6�����]���������O7��M��{:��=�cK�`��10�a��]�Ï{~v�k����-�LN�"�q���Zy��Z��2C�g�P��{Pg�Vq���bQ3�A�\.�4�h�Ǭ�.���?;�b��P�G;�!��e)���,k1Y���vײ�����Yɴ�e�n��)sf0u�(1�����G����}��Ǐo�����Ǐ<x���||||zzzz|x�9��z9}zwt'�c:1F�Gh�E����N�I�����>�H���`k��(��٫x��(�}3�t��{_�'U�=>9�w��=Uf{6����./��:b7{g�O,#����ҽ�O\�}4�兌y�7��˶�����u����S�d(U�p�0ȯe���,َ��^P��c]k7w"f^D���GOo��s��,���.��o����KFރ�c���wv-HZ�$x���qx8����˻ԡ�w�<$.�Z;�8w��G����u�u��Ԥ3ݘf��+TT�m��ɏ:�NKЮ���=���zȹ�2��;(ǐ
*{�Bw���[^�7�p��y�m�n�t�s�hٓ'z�ye��>~��LO�X����b�+�].�������5�Ŕ췸������ф����$̘"n$�f�^��7��oqƀrkڲ�APj��Cґ���W�u�d�5���Y�9�W�m�]��f���nuOC軷@/�^C$�e������9P��.�Y<�=�vw�-~����l���W]x����N�xMz��HkcJ�޲���ßo� ��Fs��Oo�k���׼����@��_�Z��+�vٞ�A�������<����ElV{�#Ut���FXϖ��^��yA�g.vݶ�z5�8��5B����E�=�	Z�w��A-�%�[IYGLӑ-�5"Vnk7�3Q�Rc�u`S/���a>�Þ������q�}��,-��=�n�+�X�	�!u�Cn�-��;����`����=�N���8-w������KXM�%8��a�y�/D�����7ݝ�gN�I�4z=��.]ג9����"�eZ|5��n�����+�3T�iN���D�x%h�������f'Ee��Wm:Zj��"�tm&�MU��cv��S84̍e<������P��`��ͷ))�\�����K\||���N��{5�:����A���F..]Px�0��;i�rى�^�ͺ�
��ѭ�&cM����Vj�2/oP��a��l��%ì�U5�XW�m@��,L�r**`�� �)�N��5L<rX��"�aˢ��7�uC�s�jc^���:<G��o{�0z�վ�򙷋o�Q߭���\�5�<溙�� .�k=2G4o�`Y������yU���kS�p$Sx��ʖDO��:#�,`n�)���sf��4�H���1M'Yk�mi�K����xdy�\���b���p���n�}��x{c灚\�M�b7.!� ���
lG�&�?�K�J�Ū�
>��I���������a��Ay]'@��#ݼ��S]5�f���ՁxE�U�L�O3������un�&�� �ɷ�A
�$}2f�@���oY�1���� 5��(*�[׬~�ݝraQ���ρ��v��ԦoQ�bْ�:�V�����	�o4������s+06��\ �H��D�(�SDEyh����QDD��D�O�����[�45SWQ�"���"���֚&*��&d��&��������Դ�DL[f;������
ZfH�'��*����
:�]ET��Q�b&k�$IQUD�DĶ������QQEW�>���D��TSS54UUE2l� �)�ֆ���	�*`��I��zآmij�6t�5QR�kD��GPt�V�u|�ꪁ��ت�ξ�ISSIIAu�DT�61TTG�ITDUQE?6�����cF"(�d)+[8��[i��=tc���1`�1A��$b �lmilVccF5�Zխ�4̚�1�Y��5Q.��5�M���g.���mlUg/s����&ΌE,g���DV�m���V4Q�Uj�lb��`�[[b��V�8-��[��]t`�zj���׮Θ�rN"1�ME�ɭ���g��b�+��4��3V}��Q]cD��t��o�s8�����������}���ڱ�h�mf�Y�	�;5L�kN�;��;�� 򂗦��r�_�e^���A�{=�}�{d����|��c����hc>ݬ`�y�Hq��4�%�7��;P�^Ȗv�z�Bb��Պy¨���`�����Y���o��o!K��l�Fl���*�!��zȤ�'D�Y�j`�P�#��]7oSO����r�y	�||�8*���Cۓ6�5%L�xeG�	��|�{�:n�ݧ�[C����G�W�����z��]"���h��"������mEzGq�[�V�ښs/Jn~��CL���=�Q�`y���[�{lw��,.b!�T{X�t����]�.f�+V���9��Ĳ/i�W)W�{��ڳCWg�I����_&mo_4��jMMs���i��L;��<�֤��DJ����x�.�Li%I��l�5�^.�嚦xE�ݶ���'Ӭ���mBc�%�+�.��F�yF��Z{Xt�Kd���\�ŇPΪ�L.eu��ͱ��c��8���B9��~��<Ԟ��K��M���yكN'+Z��P��	��@����j���nC{�<��Κo	���l>���֘r9ó�ױ��M�3�q��.�����y�|�T��=���=�&��P��0�H��{�����jb6�
�%�+	ɭ)�+*vi*`"7p7��Ӷ�!A�u*�20:-x�W׳mݥ�c-��f\�u��0Ü� �V0/���Bz���ݞ�����?�o��u�m2�Tzc���v��gac[��XpL^��: <v7�ߙ�R�a>��ة����K����{�a��Xw��cB��ƅ��8� c��֎�ߚ�D�}���p���A:[�]�ހ�x��|�Zߵ�f�U��6��0(`~`�ǈ�j�����c���E��������s䁸�>�ί�po���
��LW0��-E�;�q����O���:���,�{���GК}���^.vF�˺Cs���u�oY1Eچ�f-#�]�n���^�9�U�?��o@t�wA���n9�D��:�ON0nsc��f����;y!ZSOA�s36�\+���>���j�v�}k/�����c�g��ol��Uϫ�n�0V����xqd^��rӼ���� ��� ũ}r�RFq��g���಼����Rűr���]�<c����0�t�F��v�����&P+�*ڂ1���� �ӈ`�k��|l��s���
��с�Uیҥ�F���P���bu�A�u�W�as��|7��yN�-�j�	m
��w���z||�ȩ�����!%>���)�t	������˰�3zn�2N1H���ݩe��l_�%��|�sB{���t�����^��9y,������h.�QTԜأ�ȣ����i�J��V-M#����k�9�Ӊ�Y?��:��*�ݴؿ}1�=��pk�m�K��;e��M�t��ɭ"�/��3^�]�>��=�G�����}��
_����r��dR�$��؛/y�Y�t�J��'U�E�a<��W��zA|k�?���rMl�pi�.�O��J�,c1O�x�M5�U(f�[z�M-�4y��磆G(^�g�K-2 ��۪�8=�3J?*k��/��)����0�)FM�f36��qTq�/o�p+�S�1��!iyC핪�]槨�g�{T�kAuP�ysx��h}ĺ�j�j.j�l9/��Ux��a+ג���(�%������٨n5j��!x��pu�Ρ ��ex��k��@��B^S�"��̖����,(,��5j�XI{�֠9���9��C�ޔ�W�g��ר|��(yi�q�{�hZ��N��/ҵ�r\
bG0=B5��D�7�t޼i[�0�1������+��@�ʏ(DO����5{�P���eZ��2f.ef�e[
����+{+�{x�s+��kQ{���z�����C	����O�^�y G �_�dԢ]@��fb8���1�_K7k񌌮}��:~��,��������E�t�ʋe���������E:���<�U��`5���S�2cD�y[��u��S���q���UN��c.b�w�(���\�*);z�0'�c4�plė����l�}��<F��M�o��o��"P��L��pvZdV9���ut�t��� �*9ﮎi�۵��c��d�Q���T	�#.�tE���z�%�tg��`L���J_����ũ�����u5�m`��u�&
-|��B���\m�	��1p�Y��yMM6�����&�u�٬.�s��q".�ľ4�*���J��� ʽj�RZPu�׷��è&Y��,J�{&���^�����͆�QQ��Y��ɕ,5?)�ɐ�Z2%8��JW���Ln&��6��/D�V��W9�И���[O��I|�����/��S����E���3�7��a��#�:�P���0�BJ�������xOV��C�d�̘7�H�oUR��i�S�򯶺�w��/9�����S6��ȺP�4��T�R��B���K�X\2n�G� T�w�o��u�Q;�|E�lRW�&�f���EL9L ����-���/��0Ắ���.F_�א��`���s�C!�"��Y`�T(߰��C�8���dZ~k	@��,�T?5'�ƽl��%�A���ە�5���s����������X����kۅyu�J�˫}��5#u������V���]��J�|A�~�=m�M_G�_8��cF���߹��o����ѭ�7�_'�T�B�����];jK���,+C!������jKN6����µx�7.uiɽj�0\5a��܅'&Ⱥ 7Tn�v�T������Zۻ�Ŏ� �Y��+�ަ�+�~ݻ�C�T�{l ��#_^Ŵ#��Cj�[+2kXW��s.p-1�E˞���a>a=4��*ݧ���L��ؘ��44k�o˭@x�4Nu_u����¹d@��Õ�woJry�z��!�
�,����3<���,Ƽb�;��8����� �^��
�o�b���ٺ�ŝ�z�D����S헏Iz$@��>U�y>��~47����t���ŭ�1�L�p��s]�M�׿I���L����`/_�?pq�{�����N7Mi�յ�7_i�z�}�u�
���� �4�ۓ��x�{�k^7��4}%�*�!����oh��cr��_�;�r'1f�l�W���P�(S�~<�0|>~*�K���s�&m�RT͸b}�Bz��Q�ג��o���0ܦ׌|<��o�ah	���l�|��K�^�G�ɵ�깏p[{� kV���'�. ws*=�|�Pmj��{���la@�ǫz���-��
`xaw	םf�E����Ř����Џ���UE��N+���E�#4ɽbR��b#��{gOMn� �6x�\\W��P�|}�'�e��-��p,�KT���ul�3��.w�ɜ琐9��r��Y�����P�W��%�~sڗ]�נ���#����4�-2��vom�T�ԌI��N<������yc�;x[�tn��5iF�R�۶�Nİ�M���F��Թ�>��nXb�Ƒ��>�D�I���Jsk�S���v���s�\:o[�]��V��wJ��p�m1^;L�������2��t�Iؼ��6�����FB�`����j��"f�a>+�5��j]}[��#��M�1��F��Q{
�c����=[�]_i>2P��w��8S���*�@�y^7�V�r�-��0Q��G8vv�,[ ����i���=[�2�F���X�ػ^� ��%���,g�=ׅ�F1���� �o͇�Ǜ;����+r_Ov�ò��k W��c]����Z�&ޕG��3^����3n�!��0�\M��� R��Ftn����K�>R(� 0�.�9�?����Ưh8�Hwn݆cMA���&�0��
�ך��lj�M���]��w�Τ�9�aDǙ�mb���r�"׬�yڵ=�-�kM�k0^i�V�ggHAghtxs�pN��K�|��;�B(���@�f,�Y(OuT�U'rʣ���HN�]^�>9�=�d'��,`��sA$OyN���u}{���Q,��9_.���<n_k�Ga�p��¼�6�ĝ���#Զ��]͙[�W�oA)
�w����d��� j�S2� ŬϪ&v�J���B[�\�����j�b�m�ٹmч�b��x.��캐vQם٦I�o��Y[��lf�m�q"b���"w��Kە����e�a(�M
���T��vq;�؏N����܂��1'����L��Ɣ}�>ޯ�^�=�W�B,�������0Hq^�1j\��3���8ʆ@�����3�H�	8�Hu�^��<G~��Sn���>��a�Nm@�T5�ю�Ƭ��sW��Gj<���u�w޲-!�]G2q��-�i�5W��1w�'X��FU&�]���z���CJ&V���u0��ޚ�0e��a'iܗ>r+�,���I����u��O����"˽�
�K+����^�����k�g�A�8����>�d�$��͈�u*L��Q/���M�(W���\������@؃ az�-ᄍ`#��ٜ��[Q�������k�������������P��jRz���"�ǆ���A�϶V��ZV�],x!�S���w8
'�˶UU)��wj;���8�ԨR�N-�¨�yj9r���%%�-����T�F��TQ�?hl�a�Dh��Ff����1�1��Oy�ә:��RX�<Ƭ+�a%��Z��Á�?���?f8=:񬪼f�N�j�ޕ���Xt#�U��j�U�=y�A�9F�F����n�����j�Vƚ0J%��e.n;zrC�м(��zgg�Ŏz���/�� D�q&�ZxUc��8^����[F�ͼ"
��(���p�ֺol�(AɄ��w��C7��������{�k���-�9b� (�0�[3pе~s&=�:�~��iB/maT���R ���Ŧ�k��޼�����s �`�G����4��;2����3��86��8̵sv�R�k�wP�=���Ե��R����轆s ȗ~��t� ��a�'Y���Q�Z;]��i�[���y핌����Y�^��v�tEח��,�������0;�@��q����䜩1|��Wf<�7��Kf������Yy��	E@A���i: e]o~�66�!��[�a�Q1ܷ�-c���=�����G���z3������
���*�!\�y��n��b��{)�k�&܄��ɞ��4�)��-��{C�q E��8�Ʈ�eT�5jR=� ʅ��Хa*<����Iؐ��?�+~����G⣦���Lx= Y��ǭ��gӌ��Է5?)���L��)S�vҫ�N��B˩[�.�N��ǫp!����� �ҜI|����vG��5[�9��6�r��R�"��{��cB�1�.�}^*Kx&�IP�ط��k�<*���y-�}	��	�Bp+����mf�a��P�F'��F.�y�/4j8]n��C|)�S�T��7����t�&��VQ�U�fv��1����~�m\$���\��у ���z�3�{�U�u�BQmdț�mow�&�Ly�<i~K�a��?�x����1t���Ju�ȳJ�zO�i�#�y�#�p.n�����p��H�2N�1�d]yd����p�Q	�_Z$f��@��2�2�i�w��;+k{��ν.���+D��Oފ��Qt��ʥY��T����r��\�G.�d�[��r��F�]���[!�!�΃�Y逛���:0�wqK{��'�A.��uС��.ޓi�|�/B6�1��t)�5Õ�a>^nhj�p�n��ޅ�����;�U���u e��#��?��i)΀1����gVTw;�l����:`*Ae��x<#a����{[��&a�Pڢ��̚��3���ުӥy����yz��6���p2�Dl��̀��Ѭ&>~@@��q��9�UվD�{[��v�ܘ��X�W2��9�M�L�u�3�@�K1�b�;0��0R"G��l��/;O|u��d�����N���̐͗����Ǥ�D�&+�tE������;xw��m4�J�0y�� �n&%M����~$�b}�X��O@�$_���S���n=nu���8S!]m����=%~�h��kKO��-"�^�����{�kp��L�}�⮂����|����C��X����Qxh�C9i^S����ڻ8���������b��H�G�sj�#a^ӁOl)�4����ۻӇ��VF�c��� 3퍲��X�{���F���wX�(���U�h8���3�C.�{����_]�����}��"P� P%IKTҔ%UTDP>�JW�H�|������d�z�p!��������(M>���f=�oM�ԕ3c{KgK��=.��Ks�(���ޜag~��,���fR~��RLX�c�н��W�F0E�]�Y��_S6�y�C�f{���ؑ�5Fi=�3�(���)?�:�����Ät����gZ8�T�V^&���V^�dC$�5�!��Q1,��~H�2�(I��Gc�W=���S۸����gP�4[]N��!h��Ʀ9��v4�'��y��xN�󘕾��
j�������;�{kVLCS�3�dz�:��Uh(��ڽ��jc� {!ټ�/����I;��&�5'�C[����an�����,��9�ϑ�H|��>5�~9Q�99�4����G�rt�4�ե��%�ٕڃ��8����OK���bXp��"�'ָr9�}us�Q^l��d������3��6)�2Բx�����	��X�8�;�lc#�ǆ1��Th�o˘ý������n�JA��:�S�6՝�S�XH��W>�T��l[�O�k�X4���}<||~<~�����������������<x���������m��^��������װ&~���)�6���Ih�����=�u�͗jK�x!��8�_i����kW��o��9��R��C���pB��oQ8��.~%:��%FLSb��̓A�%0�۷����/�����,L���4��)̴����bf�7�����,�>���.>r��8�s ��F�4m��J(f䌛t;��Żq����~S/�Yc��'�S�>|6�|K"%�I+�O��88<5qz��uyLC�׾�� Ҽ��>��؀dw��!G���羇���dǾ<�k��]��vs9j� ���#C�x7��Q�hI�z������v�c��^�6y�	&<ޖ<H1%�o���#���ܒ��,��,���z��\w3��ݡsCl�B(����wI�ql�۝!lޅL�,ժ�ql��U��٢7uY���c��c:T��>�)��k\w��˩MJ�c�����,����W{��5b]�F;I3of�b�b�Ú^�I'��h�������G�ǨQ���d/)��Cb�'���u]�,��g��mH����sI!�ޭȶ������۵U�`}�Q9�r�;f�
�O�g����3�����b�d���1�U���mT���'���nK�2���o�y�a��8\܄i���|��L���\�co_-��(O�|ڼ��v�;�^�j���+E�c2ȁ��`��} R�kH��ݦ��h��/gg/x�.{=P&N�Xe&����S7Iֺ�[*�w��nB�m�]�>�nV&;ķ�����/��{�;��j��x ��v��K�[�L�5W���E���\�Y��B.�賓���ҝ�����UZ��|����Џ%ڙup=���K�)&G�K���g����Ճ��L�x槳}i!�A���<}�)k8���B�?'�����w]��ҷ(��Y%�QmX���4�.���4�63V�ҙ��u8��U�b�l�&�QI�$̇!,���OM�}�֝ō��Wѻ�������L�A���rj����*k��i�lڤ�|P;Y�I�36z$.�Ov/=C���N��To��%E4�D]p��=��6N˝�}�;�ç�9�R��7��.�;a��v�&�#�#SaKw�Ȋ��z#g1h���hT�iHd�惔l�k��:�~$�NlL�	[����e�{��ް�iT
��"��9�a��:�W;���V`�~�.n^Zwx��#��O��>BI���ahy�A��|n5Ɣ�_	���;�d�R�B��f,�?!��`Xz�D�����z]}�r}Q�L��:��(ȱa�A*!Ү��8zߠۛM)��]�-��f����[2����wH0�j�2�}�����(d=��1zL�s��׸�����p��7ϴ>����Q�پ%�7�+�Lh����3:V�dZ x嗅��r� ![�4���ԓnc"c�>�����n���$�tuz��u����X�q��j��7[$���LX!�]�A��b�1���l�i����h�D��f���b�f��S��h3��ӧ3ե����X鎨֪�=%�S�|�`֗Zu��w�U�:$;KMUP���ME4T�UV,Zݘ�ѱ%�6��;�u��]j �L5��bv1QI��*qj)*��635w�]1mmOx�c3�;��,�KT��պ�Mi�LVƨ�h�[8��(�J�"��Y�뮺4���N&�1�MU݋���*(�����Q�(�:�E�PWV���Tj&j����TTF�e+F�뮺����d�T�4h(��H�H����j�����(�"(��������US5MA���jH� ��`���*��(���E0ELTQUPQ�T��&H&��)"%*����h�*�bjIb�*)����:6H����c)��zs~7Ϯ|����n��ƉeY��ȌD�K��\���Tz$Т�7Kv�N˥{EF�1Y&LL��n�EP�ҏY1��b�^w�Pܬ��6·��һk7v'd#֒�*h$\&����e��@��(a|�!eD�fDLI��i�ϼ=���������5(w2U����=�srm8I5���� �-~CL_1ᙼ[0nu6�a�^5�?�N�����GO���a(��w�~Y�8�nt��hgZ ��!�ap+��'p�}��I86��	;Iy��U�XrѾSսKE=�������Dw��O�T��X��dk%�!��Ρ3]S?IO]�����1jӞ��!���G�_���}�S������zc�IՁ=8�m��wH�����ƺ��ū7���s����p�.yب�A��(�Շ�T5N��d����x+!�u���'��^y����úw�Y󕦱�:(Y��r�W�Fq��{�h�c�yA��c��xl���\H��>���r��p��0��w�QVս7�sX�'���.�g&;�ʋ�-�-�
}�ڥT����Ѓ2(#N8ʘS��d�9R���Ѓ*�~1I���J��_��(�ZϢ���n�7�r���`u�W]����Z������vx�A�$�^�<Ž�'g9��
�;5�҄����/�N�Gd[B�Ӎ�ck�N5� zr����؈���&��̱��D=��e��["`��f�5�wR�,m_̏rrl�LU��Z��>f��������)<�;��y9�d�co�4/S!��ۡ$��qXسr���2�w��л���{�^�O�	سm���\fh�j���2c��}@������Z�IYj��7|<�b�ߨZ{	i�n�z�[�'rA	֨r��_�8�F���m�Kx���B��*���JOV�d]��9�a���~g�l��]�ԍ['����U��7��pcΥ�=ңS��Vx��r�W<��E�(,H��'���@܇��#���
�MVP��������p[�З�s]F��0q�h%Q`����
�XH/v�k �C�7��_!��:{�f�2���0g?2��c� �c�{��;MVJok|�>s?s��BOl�'Kf��ӳ����i���}>��"���L8�f������^�r�l����u��<y�晚e���ח\�=�U-�yŗ��90!߁p�0m�F��z`d�7�a�I֌�KoF=�f�V��^�0���	���zc�)������>��/��KwfZ���������X_�?Tso!�L��ȵ���Y����yt�I�ʇD������{��P��u^�Q��$#1�&3'{�\f硛���D;�^�}��B8��H��t�o������s�m^�v*(Vy^��=2�S}s����&�T���oL�V6�m�q���ƅ�b2��f D5�F�!.�\�Q+Y�L\��͑�	p,6���!㩂�l^t[�ןr4|U��ط:j�UQ�Y��ykUrV��P�%md5�����_q����ЋB�AH�3{�7�ƍ��ܕ	�p�^_~QL�>��Xr�H�[��/3Q�箿��ƭJB�0�&���)�����d��6�h�>v���}�dNv 鬬tS�?6����K��w�*4�߄�8x��$e��ӾD�U���H�,�U���@Q�R�_>�g�M@]F>c;3�h n�{=�Q�3���q���7D��a0L��9�C_q�=|w�$?��'H>7��⓳5��*#G���e��C�	�Yơg���2S�c��'�O�GU����1��O�cb�ȋ��T�!4�ݙ��G&׎�,53R\-y��c*�.�o%�ʥX�ʂިn.e�-���%�g~�f�w��'��@ҾN��[�z�У�S��jv]ZoE��I��d�O�V���E���C�V�]�����{|幬D���bK���uLa'#Ww�����O���9�p��9�C3	[ώ*��Zޮ>*A>e���xY�n�0e��&%�D�M��٨W��8���k�箎�R�YR����zK���{�Lw���D-�xH:1��(8�@�N=8��V}�Q���iؾ�Ww�:R����Ϧ1�����'�j����=����:�i}��i`���^c� �A�_���si�bW��ɵ(�/`����%�Jv{a��>~��e��=�^��L%U�T��*-�&-�@��;��1�#�O�D��*4���(�%@P;Ϸ>y��=ﯷ�����g$b�e1>OO��gӯ^%��z�?P��~��+�>azT��}#eAs���/���K���	v���ق�I~�^=%�;	y�:"طPwb޻�"2w�������a�4����xQe�v3],&�ݬ`�y��� ��i��eW�z�j�g[ְS�Qt5��C��# �ý�O"yzs_2�nb3qS4��sy����#jUS�
���6G�G�c����1����M�C�ٲ�|<�����I��\���O�����r����U__f��y��LZ �!�Z�o�9A�6q=cռ*��[@���ǧ��i�P]���wQ����o7s����*���Jm�eMhħ��l	��z������;�
<1�\gwAI��Y���|��ZzB�����dp��k���≉d]#��T���Oc�X��t�],M���T��W܎�={��c'1�D�<ZG�m�|?
����'I��%9��}B��WI��ډ��l�ts;���y�r��b���<-��f�O�%�)���q=�i'b���~ϲ�ޛ����2�m(�\3-�[������z���u+�����㍎��Tm
tdT�q�_�C#3�:5��<L��w[V*QU���18$�~���o��)ؖ�Zd���b�ز��5[4��2�Dnjt��Vw�>��ґ;GWWy{4���� s�"Z
 B�F��a@��D�@�~���w�sy�>���msk��m�!�D3�\�s�f�b^ˁ��<��W�B=D&ژ��;�����EK����WbYh^�"�.�E�KO�/K���Fi����,"�)��u&�ʢռ�Vr�OyIg(�b�*����K$kp)(�E��q���{���X9/�e��H�����������)��!2$�ѩ�Q�X�c�R~kZd�ի�AU8�zwf�vNϷO����lզz�(`�z���z]��wV<�@,:�/������W4���t�����JbX6���p;���4<���x/�	�=?!���K�|��A�:R|��f�v8�܆����s}�v�g�}���WBCJ*s>$O�0`���v��<�wPny �uo2���|.ad_i8��1��f�8�wC�x�tUǡ�l/���צq��/tM�s���+w7�-�ڤt���	�x��tv��]���A��F]���|�=c���x	��?E�ǔR,���s'��N��G�m�W>���^��]-���Ri7k��q�eC [:y/N�/7��+���;hHyZunTO��	�"��[��D��WZ�IS�U���Dk:|�}��>��*�v/���Ϻ�c��fw}��1��ڗ�&B����cfU���x#vfP���jٴ�=�veD�+ǣowc�|[ö����e5�c��뿞�����i(Tb@���Q"PiD����0 0ox ވ��Iج^���F������	d��``���A=P%��c;z��>0
E�N[�LL�uR�}i}Mg��`�
y�#��ϦՓ�
~�k�`����#B����h�|o�0���T�����鎟.x��[k��벟 �<���#���ˈ����~�~�z�2��o�Y4ݸ�CZ�:׏k��f��i�WOM0��Ы���1� �؆W[,�	���j'2�3~˸�Zw��7y;}&K\�6�A"h1eٮ�n��F3�	���y�1L�)�^^�̈́H�DǄ��5#����Ͳ.�q��K��=5�N���.��OE�scL�3Eb�`|:��!�<4k��"Ii0>�|��-G.Qz���5�i��Sÿ��.�K��o+/��ˠ��`�bn/B^u�u��7�2u�߼L�1`����
�[ïˎ'<1�;T���-c݋m驩á�2�i��sH��1oW�ƶH�4-X1'\u��\�p�B�J�mu6v�:��/���CWB[�4>�1�@ߗ� O�}�3����{��nc�(���0�;�t7��z$NmO���2�$!{,�z��.ӁF��|�L*\:�J���Ϯl��E4��97��Ak��4��9SUA�=���Q;�}	��nwyx��8$	qh�0�2���.&0N��p��N��^{�|�����" R�$�P)@�F�i ��s�>y��}���y�������9N�L�k O@��O�n���9�l,�Wyէ�H�X@�KǕ������>/&{W�w���LIz�7k�&e�|tE��tg/#^]��ޜ�j��g}TmV��Y�C�CͺaB�6����8^E���	��7#���\�O[��b��D)�vwۢ�SwB�g� ���l�O`ME��Xݍk�D<���.U@C�H�7�/g|o��M�.����\�I ��i�SWᮊ|��Gw�,�㻕��O}r2��-牷18�8B�
���?JmA^��yTRv&/Jn�C����`xپ�z�z�����6���ώY�b٪Uf�ꍊ��%�x�	�F�)<#r(�f=���p��v�[HN$�P��H?�h��-�+��W!�t��������nB�Jr�	��%B��;YNY�!ī�V���*U�n��K˛�FNj�}��S\=�L5��@�>�5��t�	:�t�myb�T�P~���a8ghyh$��qʻ�[.�d�B��=ˠ�AƑ m_Qw�Ȣ�)�]p%�͘mo_���Kz2S�>m�	�;Z
'�U;6���8�����_�)�/g��F���f���3���3sRT������<�B7*4r̯���n��0��D1q�4ջ��6&swV%�I�X��tu�Stނ6�� �� ���݅�E��l��Qzr��E,����މ$���a�iPf�!P�R[���0银Ĝ*7��<������s�cX�uzc�7M�F��wqOM8��s��	����ױ��TsO�O��֯��"$�0��������}4K�0��m���oF)|}�*7N�ٝ����\�
�w=�9�|���A����C����-��.j���n�b*�R�v9cs��WJ簔�Oj�M܀͵���L�����/Bwy���m	�����i��@/��ٻ@6�۬G*Lo����3���1�z�����ǻ=!�xvC�lI�C�gus�o Ȉ�y�ؗn}̀�`��_��zK�$@�b� lX	�l-׻I���ѓ�/;��'iAD�����L/R�GѢ�qr� �S��T�__tS�迣�~B=Pa�gB�6M6wv'eO����T:ǆ{M-(dv�I㞭���#[��f��J��xBj�d�ROٸ�;�,aho]�Kנ>��j�L�P��C����9˗�pUO��	0��ox�����L���l��$1��0	u�s�8����t�w�`qm���R۹�.�N�l��IT��&4ld�y�B�co2�C4��<Ҏ�%�h����=�;�������wo�3d�5o�_�K�Zm�DTZI-U���Rs1A�Ӛg"h�o{	�N�q'���m�3{�.��׻�^y��~�K,�� �3(�	@	 3�89�G8ycM���ܪ;%���{���g�>�����
��摿s��� �;~ڊ��%6�2j]^E�^���Z*��Q��bz)轩��a�o��;v}hZ�,.D@��`!�*���N(��e��d@��0p#��uŒ4��߶���B�{�� �/��5mx��� ����A�%8	>9�NoˤS$�C�B� ��OAi��S�G���s~���ڽ䝛a�2��.�M��q�&Rvtκb�ij97�c������z�X��4� x}�q.Y����k�s����E�^嘔��ΦT��r,�z�����	��y(���̤��<�F&���3�%�]s��r��ņO*��P�����,a���Ϝ�B�͞�\�e��5�����3��b]��0��X���e��:���Q8G��c���8��g������'浦M�XW#��U#5�ݛ]���Jz�~��eu��v�	�/ ��%��쟋�6ǣ6̋O��1�:�ƲǾ=>��U��l�秚�C�>V��i޳��Uv2��9g��&,�}l/R�$n�3�'ә��7���H�טy��S�י�2ٟ�:��g��s�~��|heu������x)�U0�pT*�g2��-��l���MP{�e��	xU���H)T�]��J���.n95�kU[a�ċ�����Q���nz�nT2)����Qh��ܙY�����CZ<�����!� � ��R��i�i)"
"PhP�X%��x�  g���lHghCk�ڢ���^5���Ho��t4?�/�-�@���_<�S�%�*�b���=�o	����t_��v�9�v-C�[��tE��9��l�w�C�q�穨I��Ⱦ���H��Cn��D��HU���$=��[�#���hs}�G�x��:��AI>X��A���nf��]#�򤰴�ĺ½�#=]~��9АqVa-^*�Hų�E��F�Oޑ�<*�3.�H���^O7]n�`d��;�c�f�yQVժOͅ�Nm@�U�c>�=rګ/,����@Y�i����J�k���B�9�Ω�MC&= �2���L!Ad���e�e�B���9ûgѾC�UO5����������b���Op�O<CX7%ڄ��M�U������^�m����tD���BՉT��~�a��m
�N7�H1� C�H�!��w��M|�������M�����Y��4�2�0:�Б4�3��|�����3�w5Op�dr��ZzW����@C^m@�����&
z�#6Ⱥ��4�/#OD����y����O����><~�o����O����������>>=�}=��{~�/����s^{0��&-���N�'�7�9���iM����Ӟ�s�_j�o���9���F\u�*�,F�i���ɓRW���:��"�#aa"��B�͖ѵ��M����L�;j��7	�-��⻔;sŋ@z�x�,�DԼ�u�4�e�u���9�#b����wR�-m๻������a���p�6��d�m[�s+j%XN��&�P�{)k2��wQ"�ՙ0��&�sNQ��ݫ��|j��އFvE���8��_l���E�0O<��^|�QvL�;*���w���ry_E��4
O��z�<h*ڧ�e�`Τ>s_�ܫ�d����6]-�ù�`��/��J�; _&!�ܣ����/��2��>�곅t?o���z��Z75ǲy�K��s�vF�q���������g��D�����n��ƂdO��C�]^��o��,$)��D�9=�!����hc8&�ٚ�Ѡ��l�!�P�E�sv��V����lKlm�郭CL���G�uŅv�sY��݃��ƛ\q��q���q��-�-%_Ṉ�(Ù�Ä�,�Ĭ�m��Ks5i��:E�����gV{q.�S����b e���u�V��blk��ɚ�5��Ga��z���Ά�M����:OU��ϔӃuM��q��n7��V��sg����˜���@��~j��a�軗6��0�y6�e-詭�q�Q�^��)(ײ�P&K�B.Z�;&��f��6�LN���79,h���s�̶�(X��]<�rI��m����;�#9�b�Mw���e��ez�' )�/`�nv�}�Sm���=�7�n�%٥8N͸[�]H��n���$��7�C.�� ��2���(��F)`���Ŵ����	d�Ws^[�12��5j*E���('L���P�j)�l�_o��IKmwg��u��o���M&h'E�ۗr��o&媂�9ۗ��s�=,B��@���mIX�X�͞lI^�gk�F|�X4�y�Z;��8���x��Zڈ{'��-�܍{��fj��V�E:�#5���F�jzS0I7Bc۹��ON�-�e������+ԩ�.������*��*�&��NJ��u��`��HJq��R��&�ù�ƌ����8��.�7F@�-eT����a,q��聩̽���܃������D��=˯Nؑ^3��	�n��J7Æ�>�5������7w:�1p��}oxo�Ɯ��^���vvr�K�6Z���VQ���y�5*��Ѹ���}םXJ�^6K�SG*�%8fq΋�Y�Ŵݵ�����y�&�ey���V¤��%�����q�j�{����^����ކ0�j>��V�Dc�x�Ν\�U )���-�J�5�	�M��/wT��ݬ���=и	$�A �HEQO��MG͈���J���)�>F�"���QELE12^N���*��:覨������� ��
�	�g��.X`��`�j��"(� �&��(��(��*b�:" �b�Z���*��j(:�DTޣ%U51�EHSTI�QED�LUF*��()�&i)�"h��(���w����[�3UD�6��J����i�**���(���$"
���i))(�������A55R{�CMT�UQTujY�"&��b���j�(��"����'mD1E{�"j*�������*�h(* �f���������*�`�ջ�)��(����((�����f��"*���)����������LI�}W�9I��ɋ��r]�1�b��a������������ղf
���C>�Y�Q�V}[���oz��;��y$�� &UX	�P�
�	�� �{}��=�����by�:SԼ���4(��x�yc����IcC�ڟ�F�T6�*�ݷ;�A�N�*��5�(�$2}_���.��/}60��N�� �E���nc]�-��Eo���<�m��A��"�#�B��8`΋0�c��-��c5��Va������!� gX�m3+C}Ƽ�~�贌�z&�Ж�`���φ= @|o&51^wY=�+��u�)��/v��7nL_,a̼��
�~�ǰL3N�7�������̙�~��t�D��CƎ�sʦ�P�3�`{�m��+~���y�s^�&�^��v��-��l�ևuB�=w7t���&)X˼�<�P�s�2��!�=��s�ǺY�Ȳ�@�C�*o3H�e�A��,�T�=CY��°F,�=ׁ�c�Z�Hv����{�I�ME��^�k^:/�im���P��m� &���J�|��^eQ����mk�����C����]��[�uR�ڔ�Ojy��5���-�\�5!���׹ɽG�=q�a"�*׶)��2��?T���ˇ���;�NwB�{���PN��yLEu�<Nk���w�N��ʗ�p�u�g,���jpG{,��|.�z�7�b�P�Iq��c�mpz��x��;H��;a��LX9��d��e��.����t�#*(��)�d�V�8�p�{�=�u��7���O�HD���* �B�A(��<<����oOټw�.���[�<D����d&U|hRxF�Q��p;�ᦞ��1m>N$�,������݈gm��L�C+&y���ǘħ �JK��d��XMl*F�տ
5LF���6\<�}���z�e��H�d_<0���^�c�m����x����):�1,��n�eA%I�?E�55
��;C3.WC-c����'ր$f��`y�\���i��.�;"���J.���L�4�=�be��0x����?R���$&�<>D��z��#n�|hQ�4��Pt���k$J�f���ݷ�#��Ǧ���]*��	w��'|�B�����G>^��#�U�vb �����g�%6>�J\
��5�{�7U[g>T�|�a����#_��*fv@mt��*n�q;��%e��L��uN5��3�7���{J	{���9��;	���̀��W�}O��Md~�N
2W�)mc��]H�NE�����M����LS?Kޓ>�z�1�b^� �Un�fRUE���9�fA	��s�B{/��d�#2C6O�e���/��������gB��}�It���cz�^n����˻�cuo�|<8�0�!8�������>�3K<j5��e!G{K���ݝ�����zK�x���[h�pn��T%W����he�ì�h�^�l��Ɔ懪����E75:]'K�!	jJ�#�y�������i�VdR�J&Z��	�
ZV��<��o7���'�
��ܥ��׽�B�r�I�U��K�0xB��Y�}a�p(�x��,44�5��J�/���&����A!�i�PڂZNWh\:����˴������b*�D��塨!�O�K�=[���73uh�,��k	Ld�v��7�Y�ɘ��xԂ).����*�:��b�>��<<�c�t�/=� a�1�����.�Ŵ�J���>AՁ�6�5 ����q��t�o�n �@�����&p.UxjlǏS��-zMc66��>�BSm�(2j�f�ߥ���ǫz���D�d�x�T��sy�y�c����" j:�A#sS� �L(��I���+�&���f�]��,�&s�e=���t��{w��2�D�f���)�l�`u��$Y�����t�|�'����.��l�u$�$��CX�[I���fǨu�@1�m!�М�#�}�K�z��!�q�}��>^ޫ;�ׯy�'Ts�QI����mĽ���}��lA�ND&�FԱȚv�XP��������T5�0�Bn��b���R	z������50����>���ϸ�6(��ϭl�^�����-�q�{3�m��Г�S,c�2���v��֞)>������?s1H�V�q�q山��pHr�.aT|���=v��3�8r���
�*��Ҷ �V����"�<C]�Nw-~.��r�YX��1�Hy���f�o'�G��T)i!���R�fP�� ihV���B�i+������˞�t�u��;(�^�0�{�uP�PߓH� �����y�tf�p���� :�`�^}�t�jdN���"��;��wJO�`-2m��W>��
�f�\��p^�3�8�nz%��w�b$��=t�&�Ds�aS�6�/���jÙ,:�ƲǾ=>��[k<�}�g75kO���!-WN�Ҟ�� wT?�}�
�6�pH��Ș���egj�~���r�δ��E��|�je`ZUE�?�}ߧdk%}^ꓮUܭ�c��^~KlA1%��3sq��$�/����"O�pui���_,�=���3��^�p�fD՟p���kޝż����;=��iڀ*m�j��i�ִ��O6E%�el���5��M��9�"�'��vA�����*�|hvʹ�0�qV�-@��c��3[a�m�歪�|������4�S>:	��q��9<���½3r���oP�'���'>�Y�ƺ�5�����.�myLE{�hѝ��-}s������ϐ��Fs=0��^�5���}����r0~비v
�H��"����V�f�*���7�efc��{��ћ۷f�w���%��+7e�?X
��QF�I]��J����el�Yi9;��^���^�d����T��a�]��&C�gF;B1Vre���G|��n���y]�y���p>�ЊP#J%B)
R��"=}x��֔s�+׿��nU&�d�Pꋅ�벜�������q�k-��O�Z�sͽ���a2O~s��$hZ�)8����;"��oD���q�zɳ,Ont�+��y�HmAf!��v��4�`c1C�J}�D�6 ����ky����Ӄ7��H���c���񗩆�L��O�04�/��)��xӳ�xdIOW�f�X�敥�m�\�aCU�=�m���i�/�A�����5�w�����"N�¨�yj9r�ե&xF�(Z�_��to����^��s��>�+]AY�����P�_1���hY�9��,�%�h�9��b�\R&߲��j���D�˽Xt�� �x,;8����L`׾�W����L]���@
��li���;.9c�\�
�^�K������Ж�P��O��a_���Y���+�z�C���?8����M�X&��ʯ��k���`��nc�,���̃"]぀�_3��X��8��te�� �{�WS%Sif�T�[���{�e��̻I�ƺ���~<P�DM�MBu��?�0���R�=�y��̋��L6\�@�W�F�]!+�I��=�ɞ��V��9� ?/�ËS�r�^�d��m�c�i�����Q̩�k۱��V�WA���Wl�?�c��e�ˡI+�  Đ
�2@{o�M�y}{��:��߻����_��$�B�i���J �R�H�f�{���5D����z��*����y�(�����+��a ^E����
��H�e�=S��ٹ[uV�۾�Ю��%nb�mᲇ@f��D�\ON�$�&���_��x��Va�aQ�5��k��9-��B�@�N@�)�����/�ųƈ�'sE�MF5u�����#V&�1��+���+��n�PCU"V���U�,�;5�c����a��!j�i����;����������K�gl�f�!5�1^�hR{�r�ߏN��ǫxi�O��P1�|��9a����׭ӽ҆����Z$�{�O���W�������Ғ�5BJ��l�=}Ǆ�;�e�+p�����̺]�Z�!�����ƽ�����E��TT�l_fӾ��vUc�ª��&���K��.�p5��3c�`��\���cH�W�]�ݑE�fu�+�Հ����9�ۜ~;��)��?�|h$&�<<ɳ��^}��K��^��7m����{4��b���K�Qi�:
J�-^N%�l����������^<����ߊ�Dnyw�L�i*Mn�䧩�in��;�|O�{�5X��	�~Z�9��9�Ա��i�)]�-:A6l^�3E�V>V:�JX�
�E�<,�͍i�0ú^&6-|�W�\\u�
�t��n0Bt2�nj$�s�liJ��\/=��ׯ;�~y�cϣ�/t���H�M"P�)BA"�T!���ջ�Xo�ٛkr �@��:1"7!���F;���]B�)2��#��_��o	�C�ƙϕ ��C�e!�F�e<L�uQ��M�������xn�RkcfMk
 ���iA/t��q� �f���}�5���v�#��[�<�tDV<�vO�0��o#,Ͳ��I�g�{&=�Җ��^�|\�.��)[��S~��	@x|�c��� ��.�#哗ps�(�Yx���H��v����U�yWצ�{z���^��֯u�vRb]� ��Ĉ�6^�;��94��kh5���)Q�|���|������ӱm��n���S���5��*���C������K8a���w9�z�>�w=f����׊�>d,̗��O��ۯ,�b9��	���fvK�+3v�[+k�,�{US�Ǡr-�������1��7$r�׳g�ǫxU�)�7S�ڇ�u#z�b��f��@ ��".=9BUc�^}�D&��eMhħ�(�0�ј�`�n�5FvUFoc���u���N�1��}R[��М��?��&��y�C�S������� >�^�g�P�7��LM��M�i���ࣷ�����J�N�'w��	j�!�q��&#f�~���ܬE��jb�I�����T�v�L���Z�R;AA�0�Mڲ �,����d�!9�.f6�F�}��vX��=���p~	 ��G�0��S������m�Dv��k�9S�����_����=��0| �ϵxN��6_�VKk�H���ގ{՘���E7QY�i��Ed�S�\:��?�Δ3nLpe vK�H]C6��)��w{p�tv���4�'d��R�������j&0�>G�e�� ����	��g�=3�NZ�n��A�e5'��K����������K�.O#�#4�O@~��ln��ͻ���T���d?�a�=��n��\�ge�Y#X��Q�����C꺩Ѽ^����eF/p�Ɠ�yG�P��揖�\�L^��ov���{��yvp��RiWV������H�x}�yH$����OR'���|� �\^D;k��ͯ�7V�aşY[�L��50�� �6e����Gn����Њ��H�d0/��px:?�uϜ�%婣�J꺅�Q힋�U��K�i��|��SL(����m �r��wɔ�=(��־u��������8��)�[�\��7��������/b��f��0�[x�w�oe�Þm��ȗx2��r��t<߳�w�Ǜ��V�m}�B� �ȳ��B��D�Կ�e������&�5�gh���bD���ߣ�%��Q����f�V͉�{Xy}ܛ꾘9s!iN��3(���Qbg���ww�.|���(S��i�8��M=nP�]�Ba�f�/'�G��f}� #�9��
����Ko���O�''m�wO�2�=�qSl�W#.�-��=y��a9gǍ��MŲ;�>�7t!�g�&��K�W>���X؛ΐq�� Ũ���Fq���!#!����>ۙ;���+�I1��.Xy@�ڦ �QX�5A	�� �g��2�E�X����#{unV�������/K�
�&���;C�(mr9�j�L>5q�W��K�rm,����ۓ^-o��
���:E'V0��Ja^���:������L.
O<��~�5U��tJ*��uw���7o'nǥ1j~��=��Nm*�����8dcB��n�	�c[GT��,�`t�������އA�@�,�oL�H�I�0m�)=��lA�&�F���{K[b'�����z����\0D�Ñ�a��}YW��;H�)�ћd]a 0L��+�����&פ|�bKe�g?oWK8fWN��=��l���Cw?	yO�:�
7��
�g�s�_�ܤ��9E�*WC����/�����������4��j�+9��l&��,]�uX������G��c	��ۏ~�������LO+��,<c1�j�.�G�����*�����%r�Vv��/K�L�q�*Vʕ'ו)���*��LtP���FsF�E����l�)��h�7bc0]��b���1��V@Ԏ=�y��+�ݜ�ן�R���͍y뱬�?<����{Wb�N,n��\��˥5�^�l$�}njp������`�����\Ka����i7S����a�y�むOҹ�%���Q� �z&��@���J�cӓ>��u�Nn{�R��M�&�k�u��.d9�:3��l'�{&�k�Է1����3��.�a$9�^99ݣoq����D��+`��0�۲ͳ���Q1 �	�n�&!�<��9��r&������q��yt�]��(Fv����nq�ޗaבe�H$=ۇ�ji��L���M���N�Ղ-����T63�
�B,������^=���֛�$89�ĩ��N�͚����< QB�G��^i��t�:b��tS<X@��8����#������;�}xK��IutGv���*B籆ej�J�%G\=�dN�M}\�E?�fr�ߺ��،�1_n�o�����j[������O�&z��RԞ��~f��׬z���{gc��(�뵝��n��i�q)��d�?��k6�	�1)��%%�j�$��{��~��������~�������������������������������\�w��yU��?^��<��у�6O����ۈ�Aާw�_!�G��\�4�^�����H���y�YF/:��r"�����"���|����n��W�!d(�vV�&ܹ�k!\�^�m���ӂV�u���=Z������1a�K�&�n댖i�=R�{��y��k�$���������a���f�p��tg�9ޝq̦q�f��yQ��ϒ9=��&��U1F3]I:�c�u��{����̘��JZKj�6V\�۷�yfN#��Xn�D�X{�טnig(����u�~�d�;�r����*�U<G����WW�' <!@��\LLY�3��&�6�S8d�QHP�}��E����Q�xO`����!s�S�����toF�;GTQ:j�g(����%y#�t��j��4��z<����j�Vk8��C�� �<p�o(���n��B�ؠh��6���h�d�"{<�t;B*�u�U���=#SQe��-��VL0�ZȪ���wqX�Λ(�7��5�����>�ww�:�+4����)�%��/�7%�ԇ���fp"w�x��a�rۇ������Ӭް�NV0�DU=��&��$F���R{7Q�βbi(�-�Xi�M��*t�bޖͧS���Om|m���H&�dB�ڱo�,Q[�5�غ�ܳyb��e��ܖ�Bʴ���6c�������S��cg�Z��'�	������^Ʃ,�i���ҷ[;e*��G�ǫ}(��uO:"�n�^�X}�I��ݳQ������r &3�s��Wq��WVy拂nx��-�gw���s�V`��꼧�ZT�E����jt�e���J�6"�Az,��N��$3��A�D�K<�����0.�c�ө��k�dQ1I���0_p/������sIUo~}bd����7F��`�z���\����v�6ªc���������Z���w�=�a�3Gvӓ�w=˶� ���k��X���z��� �|�j��9<���p���Q��0n�7Z�����c2&�͚�m7Fi���9�sfVr��8��{"�l�}�T���_�fj��z�'�N�t��@w�sol@df:��*�K�hR�5B�s�\�LNMd819����&��U�}��yg;G��г�ά�����u���W��<K.�9yA�H��{w�Z��{�Rde��_w�cֆ�V�������ho68GU�ܩ
pꖝg�8�Q�Oޥ�X�S����·����xl��[4�Px7m7�.	W��,H3���g�y�n��p[e�ctt�sv��_�����0dsb�O[ç����C��TQ99 �Z�x�2dX!&�&��]����n���[1Q$!	 *����"���$�h��J&*$*���&���(��$��4T4I5LA��TAEQIT�$�DQQU4D�QUQ4OS�&�j
vqQMUQ0QQR�r`���(����j�����bd���
* �&�����M���k��B(��MQLW�DQATLC5US0QDPQ11D�-UQ-D1TQSIE,M53E��1EDEQQD��SQ�2DTTMi�[�( ��I��a��b�X�b(���Y����V��j��gTԔ�U5I@DTAT�4�S$�@EEQ7rh�cTCQEla��(�����(��!���" ���>H�9�\\�M�e��@��AF�,#p���3
\��\n��{j���Z���&��e�Z�i���J��u^�V� ���&���j�N-JwD�q�����{}��k���-��d���Dp�K�2�,�-�ȁ����QA�-$�Y�CL4� =�e�̔��eGc�� ;�
�v�a�c̿���w�!ŷ1�>g�	籠 _��L��Ĳ.�<�r�]�{���Y�o�����������wʵi`>d�^#ڙ�ݳ� �V3{��L�{��(Hw=~o������E7P:j��9jw��w�����9[���ˏK�3�bH��6�w��g��<�]Q���U�.��-?5���]kO�ifsy����g��xv��pEKN[�P��~]R�&��mx]�Uu���WC��di����_��9��W�:�{�IR�f��Eo��^N*ڤ��̚��zW=��Ӫ~m�Y��E�~[Qn���\+tT�B���!�8A/0쟚@�f�y�_M���1L�/{�gӯ^&9�p��Ob�WҶ�sk6�x��@��0J��	���51Y{��:~�n�f�ғ����/.M=����YSWx3���� 3��E	f�H�dl{��s�|о!�W��zw��Lw��?wlO$V���2e	��S�M�E�3�6�������L��O�P�Y΃���2L=�N�y�K���g-���r�4$��1�h�Z���aYͰ�H62�{�R��zu^�mBF�L�9�"�?��m�?��n��:D�}�t�*F���Ƅ*���\V�8v�΄���=��5�A��@X=����n���}�DQ$�U�����v�O!O�l��@y����!\����{6����u�,G4�����-����b�p�����DDn��ե,-<��^�թ�	�#���8�i�mi�*%yQ�I�̇wm��������B��T$ְ]c�Q^�"f�(2j�7���bc��Th�!^�V;MxU[ƽ���9�X��� F��EF*�?B	��>]�vx�b��Y��ء+h��Gc�P��^E=�Ǥ�̛�Ly��V�F�<�YaONn�v�[v���~�b�_��H�I)MM�Gd�P|��U��孞�m���&Q��V�����ݝ�zi�y�JweJO�b�ARt�U�Xs�]������B
/�r.�y.H�޵[��x��_��f�z�\=�R�>9	�^�'Ӊ̄}!��iR:�3L8~3�ϓ�������Rt^l�c�#=�-�Ƽ>U�B(w��v�q�k;��,��e�~��X�:%����rM����;����ޘ�������s�"��L��U��M�խ}���� ��z��9܊
j�O�d6�WT/g�g���3��J��?�o����rl�1�.�Xn�TA�)*PeX� ��iE��pb�BɅl��l��4�-sKiY�9E=sj�$Y%�2����f4M��.楍[9.�7u.�w�ӥf̀�j3N�NA��Bx��������w�s���u!WE��l������7���=	v����f��,:����FK��riq����E�:\���j����\�m������P|��5��T"��q�Ojbn�ɋ���4�¿'3L( v���[E�b�w9���v�
]V�u:����"��������o��s���LIv�L��q^�)p�OE�� U�%ܿsi+cSe�����2��i0����m�X;��G�e�^=$��6� ˵��'�/1�,:]n޶7o`K�C`J�,��E�j==�n�4�P�qB� Ŋ�A�G��覨�yd��wa���Νe@lg/ �x�'�!'���{ab'%y����N�r�G�����]3��S9t8اZ`Km{��g�c��eEÚ��P.��q�����S��4���Bn�kn��f�m��x�;��ny�C�J�W����鿙�?v��_-�L	�����2����S�N�t]|����r��U>���p�2[���$�ħ7�P�'�3>Ű�zhG�լ<��?�X��v-���g�g���f����Z� ��s��W��Z�o#ْ�Z��}wOs�F��8ڄ�#����Q�S,���vw�� ��K��!NE�2���ï�(*ƞ�UfS��9��ξ%R���N�ݴ2�Z�Y�Y��1-������gq�GY�3��z��@���Et� ׽�;��e�c1W����&��p�	��Ŧ�Ќ<��ၷ��gd�L9���%��;O�*Jz�#6Ⱥ�1��a��v�B���c8����{5�A/��]/�b�k�wS.�����W���q�:�"��^��zT%E�a���VS�%8^�g�9m;��(nC�ˇ��2n�D�^���F������:�o<sI�lS~yQ��9�x�s���0�����ԸK�?�h�,�ZX�x��>�>R���r��͍!�*�Sr��,�D�q�_�s�J	{k���F�s�w��@a������������M�qH��(�_L̥�ᬾóm��E��xg%@�~�ǰL3N�&���8���g1�����v��{��^xߘ���CM��Z'�^��N�vQa^&�b�0���L˳f'ͬ��漌��ZoU�Mt��ּ��\Ek����zO�*6���#ד��~= ����gu��V^�ï����iC�����؁6>A��}�	%�{��X�ݫ0 y\�>�X��_z�{#0|��v���Y2<�&�I��[�p�m�>.�A�����}c}�ߖ��uҗ|f�=7��=�� ��1�Qx»s����n�^&�ր2�j��d��s�++{w���WB��}��vl�&Ll����DBv箖5�y���֤)3"nbā��~�6+g�y[�z��r�9�[�:l�.s�=����IĈ��.��d73����U*�%_��=-�U-�^<�.{aUj�R��}�*6Y�����`B������rT���V#7[�'v��E"����1����Ks7!	�I��P�hR{�r�����z����htZ4�j�����6��&�_Yq%�;��ex�8\)-�hJb�s�),T$�Z `6{f�{�S�{[9�;k�����f
]K�f-�.�4|��+6�d�|�>��?BH��S!6�I��t�V����l����(=��z������b!0\��7gcH�W�]��!c6!����Ӛ�Yٔ�9G?0ET�Vq��s��g� ���Ł�±D�Xd��q~�����'�CZb��g��#�SN�RwGt�Ǥ��䠱�ҡ���wY��^8O%��~�G����*���ЋbT�iߨԖ�'h]������sV�=C��*�� �8x�V��"�Ú�/#��#� �5�:�ژ�Ρ�E��1�4zV��%��W����?�, �bÙ�E��j���הJ�BCT�q;��+ ��a��&Z��xQJ͜S�H���jx)s�(�O�/܃��ɞ� �wX�;��?Fƃom�����N�e��ꎴ��wy�影�cen͹58�D���./l��ć�,����Q%�؜�8p�QϿ}MH�چ_	�&*�{�Q7�'���8�Q':�����O����&}:��i�CSe�-��b����\ʲ��P(���0�0?|�jb��y��lMI���O$�����{3C�f�.��I�D�T^��-�P��dtK� 円���E���t�T�4��˗3�5\�f�TF_ ܽʓi���h�i؜��e�NŽ�8S������o��|ku�����T��F;����cv�3Ez�K@����K�y��OC�mᵡ��=�B�z�Z���٬^\���i�����^��[Hҕ3e�е6�5�Pz���1k�c�5�r�]Gsk6$��j煡I1a�:�@_��MW��YꨯOq�l(2j�F�;l)B�}5^�v4<������
��
�x�o��P2@���DC�ղ�>�;��Lz��l�E{�����?[m��D�)J�]�v>5s�:y��6���۠Lc=� ��/p1k�yoG>v�n����>1)ͮ�L�$�5��d�պkׯ�����{�N.N.h��}w��c�_�ix��0����c�<����6�E�Ħ·�"�HmI����lL�Ŋ�99Q'N�z�,$��u�����SNC�����>~�c�����՝ �!�5�،��Nrh��Rؽ����us��m�*����[P�t�����ᇚ������.�Ϭ�w�F�v/)�M�)W��a�K�}|�>�h�B6-��f����ֹ����Bl��K3��-I��T�I�M��'��ZT��f�-�-�{�f�����:K�>�H�F�3�xj��]��r�~�7\�ge�X}C���~osr$�w�jE>��g�D���gaC��0r^4|��	Ż�RV�j�z7g���f20�{e�l�*�QG��wwfe��\��j��T�9x�(���[򁣋�'�&&�զ���`�zr^Iމ�׹��X×���;�^��i�V�_l?���#a�>��x�����7���(��ˊvٚ���;s�������?,�)���i�!�a/:Ŀr��w��9���0Z���jVkFh�28j�Q1i�����u瓸hA1%�I�b�8�w{D�yh��ڵ�n�f�5�&H�n�`�k��^�;)�j�͖s����}���zIv�Uz��k�F��ZB�:��]9QS�vcȨgX�u������.��	�N�`���_j�G��۵���40���4�YX�C����,���w�g����@M6�ºQT'�O�ٷ&{����|4K���1���*���w^��3[�AX�� �n<f=���:Ϡ�/�)�;�����-�7�MZf�6Kͧ���[f&(T�VB�Gk;�̇�t�G��<Bs�[��C}�=8�C6q�����zw�\e���D>c�
���߲���c5^�g2�}V���j+��Ȩ �xZ�,�$k��;��}k�Oy��;:����"�ơ�B�F������>�ww� �����Хr�0�]qm�uEê��3Ǆ������X�L7��+cc{�9S]�C�
�-���*P��Js~Hд޹T����a]��	w!� ��л�g�y��벏� ��쬅q_4+z�ݞ�ܼ�b���mi���OM܅L��:#�u�z�;�z(Ժ���	 BF4�C����R瑙YU�i�)��E��pAO,��VNjn��x����=�7�WʂZV��K=�q���TS�v���=���I��a8^�i�R�:/o��^�r���),hr�v	��V�><AY��gc�~UȦ/W�����'z&lAW[�7�_9�҃�Z�����f�?W�a�ެ45u�g<�,:y-��־@�U�'��H半`sl����1'\u��+�''=����l(�<��]	l�<�*��΃�s��e����w ��L,�w�u�5f���E`=��/t:q)��B*N��kFt��Gs�}����wӑJ����{+�F��'����e�gI�ݲ�NQ˵�� �zhj��"�^'[�E�8�y��9�o���9��.n=�o��~�ˈ3����D�U\���;�����0ژf9;�XkP�J������j�֒ޘnn�0/�,!��FaWL[�kl���7a�yAH�xC <!�<�o�&�u@n�w��g(��LIz&�\�l;mHs*d���K����;*�7\�J�Q'���Q��dP{s��oS��{/;E��̡N	��2;QV{{Z/���^~����L�O���\�Oph��cR���BN}5~�Ƕq1��}-���n���&k�����ƫ0���U�C��6�\m�j鋇U�MVb�b�^�B*=�p�x�"d�!�SPZ��UKcP�d.{�2�WB�G�&��xf0e��j�����걉z=�v��C$}ҏ����F$R����;�����Jm��BeBѡI�Q�~=;�ٚ�]��P�}�c�^UϽNjn;��6�(L����|���M�1)��),X�dUԒ���X���A�n�>��{lw�-�H>P�'�ƀD��^�I�6��vW�!�'7z:/�6[�b���&���=��z�� �6H��=��5>�Kˏ�qq��"�Oש��3ޑ��y)��(�I�r[���2����r��<2��uiC��{�ڹI����
/觡]"	����c�	W�gn�O�f�:��<�<��Xİ�TE6�)�F`��KUb�j�2� Ê̹�kl�Z��h+��4��ﾮû��c�3�.����3��yc�[R1�n.e�p��;�B
��GM��Sb�r�3E�'6�6��b�x�y����%U���ɹ�����T?2a����C�SCCU��5���}�H��ke!7W�'�P���'h]��F^�Gs����z]��CQ{p�{��ݴoCC��U���	,:|�ǣ�k�4��lW�E����a����iA/t��ܪ���N�_k^��2w�;�bb�;t:��^��]3�6����O�T��g�|ő��dj�/��7n�D��j�i��'�>}��	Z>a`^�"�w�,��oݳSL��
s��?fjl��B	vc��Y�� �y�I�Ũu�v3�w�����D���{u�sN�Vތ��<���*���Zy����j��l!��7��
\�7Mm[�0�����hm`��)�Z��i�P��������C�w�F�I`h���R]�Ƚ�O��C�Ӻ�x�KwB�t����F����s3�|��ƮKi�0�M��	�$~z6�=><~����z||||||}>>>;����y��NNNN}���\�u��u{{��g�lBI�����ΩM=2Wӯ���j��&Wp�u����u��}�6Ys�/H��S��A��T'Xw�#\m�2*+�[�ȡ���.^�Ocl8ִ�R7!KM����Z(&jբ�	�z��Xd�7Gc��y�c���{�r۷s�w��������Cn3�dy-/v����/:��v��:b�	�ɃQ��{�U0�wXE�j�SN-�2�Tѭ���8�h����v�M0�8�ݥ��sd�p-���wB�4�=���捛�ݜc�*8����񺻼9�z�HK���}�Bac<��3��)ӅHgN�-�.R��0>t�*��G�.�[S�;�ۇu<b�KJ7v�����c>)ޡ�P�����=`��V?cZp���u�D��<�v{q�\z�9��=�c�5��$x��>`p�N��a?��N���J�=�r�+&
���B3<���Y�b�	�״��T=�,����Iw�8���`��"��X��:k{���Bf�6I�D��J�%FT$6�T�\�/�w�'�O|�mU��~z-�T�%�OcC��S�&��x���H�؆�pohG������Af�)�ɼxQ����Z�Kji铔M,՗�BTjS!��m�UQ����yfdc}�y���w��M�.��E���S�l�uQ3�f���gb����T�>���1zݜ�����{c�^�ʧ��]�FR=���;��p�oY"�C=������,�&�"s �3�MNHg ���9���u��վ���7g}w��\���A�zy���!��fz&��t����) �7q�TBg�˄{v���qV̍�z�Ք�QrkQ��'�$�!�f�s��L�ZV��i��`��Q���%����4躋� br��.�&F(j2Ě������!,j���m�W�1f3=�}N�3�-��f7죏H5�#�W����e;>��2�]n�=9^����8@��7�蜸��]�Fm�i:f��ݸ�P'�WiY#j��[�QL��*�a6��uu4ta5���͐ 5{��>�''��n\{}ґ���>��mӣ�/'�7��K��f��t�Y�
��p~N1W����foOy摤��[�3��s�S7:9������sg.�i\n����Ս�1v�ٷX�1$��a�EX�����9�b�#F��5݋=49G�#&3�{#>�k�7ݣ)/+e�N�<yVF��S���4��S�s6����ϣ0������帿<�qonv�鸆���t��܏�,����XI�Lb$hVs�w^+��>R�H�=g�B�{/�EI�,��w�.{ՌLy�(��[ۓ~H\��G׀�kڛ��6'	����	�bHՠ�"[��Z����T^)_6������4+Ce��	��m�;�}n�u�Gkꩤ�h���d�։�*���
"J"��WDQդ�ITb�����b�(*�C���=�TMAD�MVH��j�*�������"��5R�QEz�D�HU-4M,MARQT$HTRTlhb�����))��4`&
h�*�*�"��������� ������*`�JH����w]i��4�mK%�Q{�SDL�4L�QQAETD1URLM,IRE�CTDR�PP�TR��SE������ �)j��)��"�R�)�d��

��"JJ����(�"��!��ӥ)ii
Y����>z��ߟ:�����W�|N��m�
�����Z9�LfޭF��/ֽ�h�*�m��p�Nm�-D�	��x��V���2����p�90=���?�<����T	���W��ҫ�'�6��>�"Sm�(2j�wM����u���MKj�_�_<J�Ui�P괟��s�#�6>�(3��Z�b�{�s4Q3�w�9���Ă�˞�Fi��J�]���Ʈ{gO"���A����vm�1L���VeV:/��y���=+��z%:NC�Jsk�S*K�����Iܭ=Z�|�����ݧo����=ݼ��u�P/��'Z���&f���4���D�(l	'$��A����}hLz�m伦�UZuwJ���;�D�ٽ�jOxT�O��jzŧ�2�^���:Y��7F�.Y
l���5�sҦ��
E�^/�p�s�����Z��k�9g��|r�U��mܻ �ͭ��!v�t��) Ļ��3���7uF����x�{PQ�v���&����6*]�յ�Y�;9�g�/,�lʷ�Q�5R2�-ݛg��� �e��J��>ʕS��n��W�f@@{�3��5�H�Y�:��WX5\��B���ށ���-)�y��8����{LniZ��z����3G5�𛍼��9(˻�8v8����M޸q/�!CY�������iz�{�-�����h����L
��G�
�Z���7��㍯d�x�Y��9l�
A꽁ĩ��le[�`�C]E�.�f�C]o_u6�=3�8�=?���s�İ8|�Gh�X�$�%�������_�;x�j����tT����v�зp��8V�ȋ�g�X�ԍn6;�79�2#I�.�	�n�z`��DYt�qe�l�4n�N�n�O�)�pz�2�����)�t[m9���fY�zIv�T� �0E��|���)������?4S�̂�v<Ğ�au����U����U�/� �
Ɓw����R�o�}�����S-�^�g�f�2�S:|�x�`d���f<��蛐NwlUU)<��d�ǳ�;�����A?5��OV�K*�F���c����sn� �\�b$����ouǃ#(x�3���9������Ң�C�����4)X�I��m~]��^ꋇUq���m�?T#�q�q�=5���(R6�����r���LZ��W�'��%9oZ�"�ʤ���t�	��Ň9��}�Y*u�F�h�%�sz(��tD��!�_K1"�˱�R��7��֝��6���vv�p��G��-7~���T[	� ��>�I����V�v=�'��������}�^g�˪p�(@�rU������e�x���t:��AW������;WAMw���IM.��Rj��Ξ0ќ�ñ��Um�td�Ǭ����Y�%�h��˵V�b��i�V��M9ZiCN���	P[�(�7�t����s!D����/���ޕhru.I6L䨨�̭P�?).��]�3٪����A q4���@փ�U�W���ۚc����B���/^�|�R�)<�ʄ_�PX֥N�Bxw7!�FW^klx�=��R�g��7�^^���9~^�O�
�)V��RX,��5a]k	���<c��>6����|�5t���/���\�	��2��B��ĝx�Q=+�҄��¨��B��T�=�Z��2���Ӯ-Wk��HAÇ�6��u!ֻ�2�u�W���StM�.#Է0���N�.ǹ���kz�
�V�ԃ!��
��	�<F[���d�1ٳ/U	�/P���)y�V��=�&m�^�2��Y�-�<�˼!�`W�O.����}y4`�u��I��
�ތ��Y��֙���`��˴�m����y��{.2.~�����g�o�(ϺUZ����w��W������9ם^46 ���
}H���#K���wtd��K�S@@�W�-�CyH\�]DZ�
�Rq��Ű��鯏/��ߠ}w��2|���m��w�q1�g�W<���J��y=���xpVa�s�;���rY�M[�ZsÞ�kN���ݴ��Cˀ2I[6R��b�"u&�4�����Τ
���s���ўXU����I���j@;���ML;�͠п�SX�Mu����=�F�È/8c%~��a5� �M�vBe^�hRxF�eu��5���#������+_}V��]L�K�l[H��1 �:��4��O3r�����zb빝-�hv��1d&p�����*�b�j�R�L@�O��9�P{�#��(��ʡݯl�J�|�aVs��Y��)�JS~��u�5����-}�����5��K<�vkZ�}� ��w\b���#R���,�t�>0m}A�8�TX��$}]���ꁛ��k���A-��+F�'q>8���#��҂Ƃ�P���h�y��>N��#�f�]=�t�׵ ���H�#a�W���sP�[B������3A*�K s=��ٓ�l��_��T���<!|�x���Ý~��mU�������T�{	A/t��\�0m��[��jv���UB}@k�'2
���ˡ���p4M��}�������:�S�_m�[�Fug"_R����(�v�y�3����a?���7�����Ï;u����y���Vi}��벺���)�B"*c^;.��=�3�~{y���AC��v�;JS�w"�ѵ�W3�8{Y�@�Á���
�P�8�v���F�_tt�]��Oh"tst?W}{�5�ޢ�:�"ws���l���0���LF�t�L�~�f������T�?�Oߑ6{������\��y��:h�h�bi1�H`X^���ךz�o��I�;����;�|!��x��1S��C�"�&����[�}��D��7[���sN=�R�c �ųם7s螌׳���3,�4Q�,x���r��j���J�N�\J��ev��<���-(t{�Nn�}<�����T$����J�`�.N��j��T^����c�q�}��k�l�)'΄:X�^�A����H&򢽨�M�e㎂���F��7=���1:��[���z�o�ݙ�A@����B��d�WAX0g�B��K�wL6�r�A� �W��d]#��R�yT=6՚WJ���(|��~��nӑ��lP���hn��R�P��8M��v�,��xO��H�T�����$vE��C����q�W{���g̽p[A�Py�qz\�ƴ�؈��MHn�Oyhs>��ct�IJa�����)����1&���AF0�@>i� �T��}"y��K��d���S)�<�����+"��0�?_
+Mc��@3�|���=���4�EPi�PYW�13R��j
���6m/��tKϻX��w�/k=R�/h p�Ѷf-pܚU�-|���	�+efl\�S3x`����9�dL:�����N���*�ARvg�c�7N[�����Ȗx���-��\(�v!�~e���-�3���1+�_�|�ӡjy��wv��͓/�h[L�<����ϓH�o��hgH^��q�2']P�M��e
������n.�~���-K��gG�Q�w�t6�-ݚ;����{�b�=�oY��z�Y��s����(Y��,:�/�^������V՝��4s��}��
|���n�-�ٙ�rf�O*��R��>�[�%86��
$@��[��h/a����ɚ*gl�c���1"Y�0�mgE����S�{��sQ��	�5l�ӣӊm{v�ʷ9���dL�5?
�V�/|e�z`q�ʞ>������������t��uR�6�j�l���v]���Y}�@f��F����'�Ctgۤ���1���.Lj~Ioo=P�PC�⠆梮PjH�i���*��	�S���'�!�ޘ<�S�6�xH6��M-L�)�{����s�z���4�0*#X�F�=�+&.�ky��}����-��y�(ټ��וOk�"���^�ǧ\�=��Y�}�x|=�����Y��l��<�|�ݼe��2�b�����e��3ꅢ`ڬgfH��U0Hmeڹ��Ή�F�P�M����9z�g�=n����C�vix�l�0VO�x�Ac҅�=��y�,��Į�KJzs5�g��ܝ>4# �ן�X�	�ʽhХr���/ΟT�"��M�l ����ǳas:BoFA�tƧiܑ�E���?Bd]��r�H.`����fj7��^J�꽋4�S�AFq��$P|h��j�_C1��Ȟ�T�``&+In1����u�=r|��V�P�8�A����@��gd��Lx�=�%�z�ӷd_��#��8�H@_`u��u�Y#��=2��7@�j�۸nvM(8�y���=�b�55ɑ�w=�=w���/��Q@�&Xu�'yj9r���ԩ�HO�7!��0�6��X�>	�1�0�m�s��C���A|F�Xd닲@TXW�t������ �t�U ��Ac_�+7"o�w7<�#�!Q<��ŝ��4-Y�:�=+��PK�Z��^���瑞rᡜ*�Sw��G��!��0/щ�ve�6�&�JAM�6��[^q�{}b||IX]������\Zˠ������:����#'�P]��7��x?�ӳ:�d�[G>{��<����W�>Y5�tf��V팧����`����p?f��v�lv�Z+g�0�ݠ�T<���0���T2���Eݦo�8=�ch�����a�᱖�R�w�ǄS�����o���}��9�����0��j���{�&��0��z�f��q�tE���-��4;�\`��^a�=�|��G*�r��.�w}��Pkf�B��:z�3�;�<��Gpz������;�p�i��M���ll�O����=��s3վ�ZyEkMO����7�:���3ePyk�%ʨ!�ךn6�6��Y
�k@����N^�~L��isi� ����DfM'�UM^Ե�iR>A�����㇡�8�os�Q���۪��C�QL�Dk�G<�d�f`�"Se�!2�Z4)=��3z�B���,%uQm���VM��j�FК��P�.%��/Ux���<���%4kb�ܡ���)��A�T�0���{`��k�|�Ԙ!�Ǘ�
�1�(3p�����z�ÙjF��`%�n�O�}^t����ͱ,��Fm��T�7=s�����s#.�1�N� -�~@<ؤ6�Ť�%�GtQt���J.��)��#�8����ޚ�F�|�ޚ�,�;4����
 Bl�遌��Хxi;���=.��[�7%�ҡ��'�O;�ǟRo�*V�_z��NP�Y��ݔ�Bh��,�eF�ֻ�W7aB��Z˳+���]G��}���ul!QqNr؂��B��`�%� ;u�LۇS�uc̓e���4�b�/j7- �T�fñUZ�B2��!I��Z��u���l~���z�����>|�߼��ָxNk�S�9�9m���זF���w=Ȯ؎���˗Ė�߄>���	��}�\��mG*j�2�Ռ;�,~NǞ8'K+H����mr�����s$+��dL���ߔ�G����yN�լ��wC��U��:���:��5�'�J}:��;	��w&�k	��S�a���h�|}��ƝK���&^�}K��a�gwT���t��4p����%�O��}ޞ�U�S<: ���y�G��g�����!��v����z	M���t�>/���6"��ۼ�Yz�&�Α�Y�!�'-`C�����Y�V�s%>����<�ҘYU!Q�聓R�c*D��7�}u��V�s�u3�S�~0�|>y���S�/���ڊ�j�11g�.�2ĉaG>C�:-��>gb���A�5썂�|�C�������8�:G�\S�f��̌�V��ogTWh%����^���aG�1��fA8�"X\����g���N9�$֝���[N�twsB4ÈU����|ۦDM�a�:��W��Ed[��uIz�M�0v��k3�v��Lm��ƫ�*���e����7|��w�Ko��WM��{ky?��� h1+1f�n�5[��Fg���<�E_wB��UsP~���&%�{	W�[(JD�Pq��t�)���ƔuA�ln�u�}��٭	��g�G	���z~��=��Nl%"�W�T����et���.�/�ed
ys 3 �uzu���%��24��4��c#mz����;�ԩ'�0���u���J��z���
l~g���ս�] �r������"m	��� ��.�-�$�'�8u�-�΄6Tm��Nݼ�םz�Pe�Qu���C���k�A|�|���/�ī�<����QL3!�_�(r����&�w8X�3��ݣb��G���6��=�t�hL�N��,*�Q,�f�m���[��/�5�5@3�҄\�at�q@,���aZ�y]@�}��mf!�6��t��z!t�����xmk�2+��,#�E�Y[�z}U�3�#�,?����1�ݝ��p{}~��<���v�C����v�����t���"mx��j/��nj��=��q��3�M��� ������#���c*Ad���8pТbK�x�f�>�z}~>���|x����������|||z|||||{{��}>>>oo�K����baȦ5���i�}�;���GZ�0��[�+��R���j�g��h1�-�k�fbaS�j����=�����й��?S�wY��	h����HN˽[������z��I=����Ni;W�p�9b�IV���D�
س���f��1諷e�j�ҵW�l�g�
.�`Ums޺7�D��˧[=�^��5�s�F�vape���v.�<e{��v�=�gOs���Fvk���R8����y�Vlm���g<����p)i�f���[�E����}%D����+i�/�g���_`�z�/T��i�J��X0�
�;�b��B�n��tpki�usf��֪T7P�/�u���w���掺w��t$��	���t�B��i|7����aJp6�ٻ�Tw�P�P�76b�bF���
m�w7��yY�F
��N���\t�g���w������<�%"�GX�迶��GJss���ΠaM��F�Lw��u�|���2[�b�p�BsOZw����X�T�k����M��y.���>����2�M�}�a�y�"��f��~*i><Fu��k�Og)�C;~���j�Z��%a��FEBa�ə�ɱ�d7Y�/i��ч7K��n�,`b�b�Q������:��U]��G���o	\@2?
Θ��	�z�%��vP����K䩊����ɣK�7��w ��p�>�윭ۻ2���t�Ƞo��>E��R�@y`�BNT>��3��Y�rL��~��㗵�wNŕ���6��ZE��]3�x�����^W�|"��Gŀ�:&0���9�Gyo��7W��<U܀�x�%+9}�O�.��ذ�v^���M÷�=�.ϝ9V�0w��.`:�Ő"|������t�&�w05��cct�,�Ti�Αuݼ�>;&2�W��Ú�j/���G��?n�����ǝ�,s{/��y٤�z}Ⱦ�����k��Y���}�������{��lC�ܫ�<��lL)n٩Zv�����QOS�O"�5�U��PwE\�4��J�7?���>��3e�ݚ�-�@:��/qyxۯ��A��ݓ4� �Ǫy��M���=�&!?A^���>3����G����;��.U��Y���L�ޒ∴�Ĵ���\ޥ�I��z��~ʻЋ��V�j�nt^�W����xA_N�u���YP�������b�@�قSU;���P���`ǔ$[���FM������B�,YN�j�v��nȻ8�R�f:�8�ۓ�*t��K@���2��]N]�	'n�lD�f�)ػ�6�/��\�=�K��Ǟ�TV��Bp�{_�U�`&^\>}��7ݣG|L�Nq�H�zb�� �۔�ؼ�5bCx&+.��,N[�:+Sr��uZ��ok��	��M�B&�c�S��⪒�&�(=æ���h��B�( �(����TM%5TЕM�AMPi�
�*���LL�UALE)T44U
RP�MSG�4P�KI�T�DLA���������EQDPD�Դ�UQKDU0Q}c!UIH{�H�16�-%%PRU-T@E�TL���DHQQ-I|�(�bH�
ijH��"��!�
Z�(��@�X�(/W}8Z%��"��a����(OPu'U5JS4P��/U4QA_w�qrKTG�1�#�A�B(�A����� ������Mi���:]�ɲHtI��������4�Ok��({MK�I�H���w����oTT��\�7�� �nt�H�Aa�a. d!�	�"PDj(��l88��(`n6!A4QS�I���wO�������e?�����
v�	�%O�[���x9a�殕�0үv:���I�^����̳B&y�d�2�j啒���k��~"���(�}�S�Ԥz�j�O���|(���\�vC
�O�]���D5�#�7����<�]Z������C�r�RFCM��*�Ο�]�,:NTU��d������l7۸��0Q&Gu���CL��0�	��jE2�5�]LTm�]r�q3�)3�����ƽe�$�/��u�i�0_����Y��L��ѡJĪ,)��N5��_�o{q�CTfl�S��ߦNY�=�����0���})��?Bd^��ʃH�y��a����!(����n��eƨ�dM����g��O��t5�>����oo�B��Rl��bK	�m��*��X���2+^��M
~��{���6��O�ֿC�9��U����i�j�0�WTU�g<��vY���(���@n����8l�T�8�4`�C֠kA����E_��^���Rz=�ܯ0��*v1o�0�;(���<]',N�H��&�|�j��a���r�|���N~�z�3���Ѕl�޿�����hU}b���,M��7wx���&��$2��ѻ'�o]T�ŋB|�7`��9��ق���d�!�=n�Ί�R $������i�l���fdE*�$i�O!��9�I�ĸ�n��9�n
�#�U,'1�n��i���ﾺ��:_X�-��kԼ��48�������w��a�N5R�k˸65�R��#��`�-�,'��q��pд^8�zW=�(%�Ts	�jޥ�p�>�s2������6�V�[�H�|�#�p� Ǧ0�� �>��Z5�~��z]੻��ߨSP}z�����E����֯��轆s&C3���x�	�U��F\Ͻ\�Eԣ�c�Puڢ �ܔ���iy��za��虑 �c�)��yw����C�{a����G��f�Y���m��-���|I�޽�t*�>o�Dg�L��3��`�<>�	ʦ�(�ǉ�Y|5k�ls]Nd-z��m{���[o��K�+$!Z�y��n���h�ͤ����,��?qn�P΁X@��\O��O���T	꽩kjԤ.{�2�WAPJN8~�/�\�wZq~|i*���L>1P�Cb���9�\8�yϣ+�,$w)��L���,���5V_�=���/!��W�d{��t���<55���-��ĵȈ��^!��z@�>��,�;4Q�zlX�&,����~���eZ����w�(;%�S)�y6�̣y?K������W��n{�;g�ˁ�yAg��3��LV����7�����F+K'�A8;,�vɞ��\�C�_Og]��l��vbi�p�M��L�z���х�j�m ��n/��sߐ��v!�sZ���S�	-����&N���N(�ܧp�3E�q��p^<��L���E�tS*IRaO�|���'���k�}��{��EF5�5�ҹ��R�6�X�:}})�@�.�#0���֘&2;���t���f('[sM=%\]!���
�p�fC����ٽ��/>G�M'pV���b��_��ƗJ��V��[d�B�H<�1��2#��>y��1�xgO���ͣ9m�MyY���1�D���f�N%���n{y�W�H3�;��:|ã�:��x`1lȖO�6���T�0�e�;9ole�#n��=Ӫq�5N#x�B�`�G�1�[򁣋�4M�o�M0cj���[��K �	3�{��rb�}���S'�U��`�0k	���E"\ںP�T혶;�ӸdXïK�w��79ݟyo~O���r��u����y��b�kþ;g1���v��ԉ�`��A��H�Se�_[���v������$=� ����n=ޏ?���;V�bh �]�HZч
��2�n�e�W���s3���B0]���k�f1�&t���j}��'����Ss쿱+�DµW��/d���9-�,�yw"?������8!�ǟ�q����������x���.�f��N��E�Q��jL4շqƯˇ�Ş����!���!��	��z/���fY�h��X*�/,Q'�_�.z׶KoΪ0V�y�
��5�B(�5�G��ӛS�硹�5%L�җf����0я.TX]���&'��>�"�s~��*���B�J��)'Ђ�z}�`�EG�}
m�9�.1va��Y�Wڳ��yy(Jm�O�v�-D��$gW�Fcׅ�[�z�f �\��K=m��B%A��V�}�]����!X{��k$�5?A�9 D�/`$f�\�B��Г�׫6�Wd�o;'�a�>�܊�:}�$��ư���q�!>���OЙ'�禓��R)��T����LN5۝��t�l'9�הzql롛!�1�6��)��w�Ji'�9��[t�\���i�G<Ehj}	����V]lQ�"&f�(G��s8�?�K��T�A>Tw���,�߶��񙶛������z��Ai���6�M0����B
5���s��S�ꗛvB%�{ݬ��;�
��^M�-��(�z�,g�ݧ"��<�<1�8B������||\q�-��+�w5���Y	�z�y]��e&��;W�%�a���=M���s7��PlN�HL���z�aAK��S0�(�35	��J�YM��`t����X�Em�S}�r�K���;C�^��鴼k�<z��b�
:{?i��P�,������P�{�h$H�v���N�{Uw� �[M��D���ު�L�A5�vzJqAgO�W>�U#+b�٣;����֭�:kh��D!�9�������JNB>��Ia�^5���=>�g_�>����Њ�3.�Ӿ���#�/^��놧�'����sP�M��>m��:Rpm?M0�Ky�v�1\�Y;`,ٵ�t���j��[Ol��;��x";`.)��_��&J��7<��5��.б�m[I��Z�n��\�C��3k_>;�����l�A�3����A�� q��F�_nl�
���f��$MB��k�+:�@�<�T�C���9�=����V�f|�BĊ�gͮ�Q��Ԗ�m=���^[M�U�Ũr�ZFC^�2&��s�[=p�~o��8jq�������K�
7#�Ecg��W��TpOV�K*	�r�n2�*�0k�������9�W���Sa���C�l��O]�bq�Td.v�!����E��b��Qa"��I�yM�E���鮋�l��\<�����F���H���Nۇ��	���Ʋ.��9og���"M^�
�|=���o�*�1\�Y�g���YSq����R'�Al��-Ԥ��j�S,�b��;b���,<�?��v;2<C&���v��O4��a�漡��p[��øi��:#V����ԓ.��w�i�N��0ҪnR�ZR/��,1�Q#�_�~�������ht�z������|�f�@����*�D���&��گl޼���ʝ8���j�I�$M
~�>1n��'v �cH���O���?QR=���wp��I/[�P%4eΪ��\oͩHZ_d��S	@�H�MV����B�m���O<�ocY�9�yU]����v���l�T�7M�W��l_wGt>a]��g����Tr�^Y�f���{�0�pr����֐�;i�XSr�HaˤGb��J��ڶ�Osz���e�va��Ό��q��/pT�7F���1�b�
��g$Z����+*�	ӝه����6Gj�F�!��g��	@F�ި=���D�wFE���x�3�Gd�!�׋�vC���r��R��G���[!Hz�z��ʕ�D��>����F�����8�|�\o�և�G˿dj�Dغ�;��nA�5>��Z��έ�����b���3���-��.�l��v��Q�:��ꖩ������d��s�1�����y�����."{���"J3ʍ��g�O{�¢�A,vqi�mR�f��D���i\����?}T�Zm��YuQ4��3���$T��g�ܨ��ɧ׶�X%��͑��1�OT��ȵ����t��N$V����O�*�Қ��yv��E�L�i�����S��ae��X�ȁ�*n�{��N��3ٽg��� 6��5U���Ϫk}��Y7.HՄqƨx�+r���i��ὁ�ك�g�M�`�(�W�%@P}��ebi�uג# �����w/B��F�>�6gܫ�ʴ��l�$�^~���u#s�U!����{E=��{��[=q�ɥ�y�>K��${F�t�^�4O��mRǛa1�pv#q�nz��U�����갑&zxN?^,�ל����y��-IM�y��~]�m�_��{�Rp6�O�������b�wǚϘ��혠��?'1���g�$���qs�U��B�u*�,�u�(]������C�g���V
�^7:H@;�W7��$��	��u"ҵf�m-yg&��ԁs-��1"�a���<�f�0͔i^�'�fW�����޷�ض��WO��um'���и��l��7��U��
؃39��������GߘR�	SAWL���;�#��N13{*�%�E9��՛m����F�״��G�~������y��P��D�Qp����i�e���H��i������nn�3�ؘU<7�fVO�t�l�u���pF��J���u>q��˜қ�̡��!���%*�y�׶X��p�����yG�}wD<�O�0@�ʫv�}�8��b3ѧv}�N�d�����F��OnT�1��[�fi��'w��{[�����)hH�f��+���p#�}d����������Xz��{�7�3
O ��(%m�8	�G����h*��eUy�O�M�����P
��Ӛ����L#�$eW��v�F�u�:ۛ���5��yW�wfƲ���<��@�=!�"9�h%R��U�o/?��	�C�.U`l���6�`#��H�f̝}]����yÈ�}�n�ݧ�g��%�X�_� G�mѧG��$j�2onvjf�70nhIA�M��w��{�m�n3���'����KY�fN,�{ k͜�:��Jk5A��ЊY����@]�Ԏs���\��5q���~r����ǝ!�)�^���y��������LI�b�H��
È�X�g�A����b=ǲI�C����|F:����,XO7������W�������y �`:�|��O����	|Lt�9dD.�qs-u���bo�RY�.���vd1�������SH������qg=F�̼s�uR獊����&�ݕ]�HW��F�������tYu,d[�ħ��5]Md�p�F���yh����؎�寛޽ϓ#��T��2~��I1{��4������dm��K�d$H��A����=�٧՗�:�(�g9�`N��Wד�+�pv<;,�٫�����l��]�u�qq�AI��7�02�1�<%>}�Fy��c|��8�Oma��޴�y �� �4�X嶫��t5�����{����c�}��-�}�y��&:�}o޽ɋ�`��gM��G�M���4�����$=�P��%��"W��od~�fh�@0��.�t�~Q���4�Y$��臸�0H�����I�G��޲�����L{V����̕��h[l�z�ˈ�w܁�:���3~�9vJ���T��p�YJF�u=,�g�r��Sܮ�F��a��E���B&ҏVT��%�H2T��e%���C	�^��7�O�o�EL�S?���(ކm�]>n!]x�h��n&����ɼ��ݫk.�%Кg!tyA����6�G�V́��%�I������w0��[ѯ[J�wHI���ۖ�)�fD�p�1!>����u�����7�M���Ԭ7MyRD�ut���df:dy��i�óћv�����<T�I�ܥ@�zW���P�d.��黌f�*��_����smy�Z���OP�J��D��k�wO���|��sS�i�eږ6g_F�7o�-���]&����ʖw��wdV�R�YSX�fA�`��?�����[�V�8{VO��=�_��������������||s�������۟g��G������.f�lm�;EeU�M8d�{��M�]P�ڔ��k�"�2�Z��!�x̨���ܨɆ1��F�sUc�3Q���V`���!5E�����=��s__f�%#^5��FZ&��҉k�w�{+���'��,�+i��#1���a���.�� �t�r�z�m�}0v�W�B?S���H1�o���kfo`������s<��+\�+�����I���y�S��H˷i7Kx�<�z-�7�*E<�x���K�	{#w�_>�v��9D�nԩ�,���,�N5�ޥ��>�8?b����{��b�f�|���Y�������;�����0�/���Σh���99Cļ�����v�YL�(�F�V�7fojlڑ�`�����mɆ��@��BV�Ɖ[�wWR��I�Z'�������.z� ����P����x���ÙU��l=��<�r,�sݥe^S������T\h9I��dI�)����^��y��f/BM���5�{�E�]]�����oW��TN'AL�n���Pӫ,^���0�����ˎ�!o��/Oh����X�ܫ��'��l����^���\��k�Z[YY��ꃬHp̠�o��W�v�'���>0x�л|gĚ2Qګ�t�v�հ�e��p3�O�qhB�P^&�i�=��{��l}�� ཋ�p}�t��?��e�{�vWjƠ�=������b�Q^��<�<��<���4��-[gް)1���H%��8��FA��6�~���Qں��i�s���weK��)�|ž�۫��E����##V��`�m]� �x��K87����'���������4��z[;u�<�q���Y�r>��ME�kw!q�6J�Wfye�J��M�+��0M���M	���a�t��Pga�l�ѡnqv.20�R�Ķ���X�MJ�M�n�g=-�]�İ�}��(��i����v�m�2��x��&�4�X�MC������1�x_S`���8�Jw�]�Wx�f�Z��S䏃�yU���'��b�Vx����v���`�}�t0��p{S��~�Tɧ��Pf�N�m���g�x��E=m�,�+�;�n��1���gT���yZ�=Cظvw���Jy%i/3x���KE��ٱ�s����G�f��,E�lD����smI��Q�3��P�W��;����3i�?MZ$�r-Z�GT�=Ǧ7�F5����m$�UY��7���&���"rM��4��LN�N\i�;����m$І	Ӆ��	��хd� ��2���2�S���g�,���߯�����Z��=�����
8Ob�7L��mM��cro/>v��	x{���rgn��`Տ���c��_H�j&6��T�n�eQO�I�l��Ƿ���swv�7v.�
*OW>$�xO�E	KA%%P4�$t5�B��u4'�)�!m�T�IJ�R�)C�Д(D!K3G�`����K�������Rw5BT@DRĽN�������*��j����
(����td�)N�q iC�����:NHu�5EQ�e��/���ƐӥP?%:�������j�ii��CIAK�B�����}��>��[o<�}���"�5J��Ծ�o�6; ��m%|4Znnq�.ޛ�A�w�[ȇ�%�EeL��9���P��]�9�В��ߝ�F_A� �v�|4s:�10Sq����S�N[�oTז���s��F]��2Gtoj����@���`<e���3�Ë|��3/%J��DV���*�� ��$�{�WN�s���K���Y����QO\�������8����#6q���2t�r��U���D��1�]�Y:\���'^@�	@z�>�z��wo�ǧܩy
�i�����@2qu�:9;7:}QO���U��L\ɩ��t���Ċ�(.�L��k�Of��7�Kov��O�v=n����˗UR����8�z�]��"s˔���I'��[�;�}�v�~4��ͻ��6*��7&ؐLѷ��#��ӣ���7�g�
nAu��O%BUO�s��=4���[����	�Ν}];�g����7Ґ
��4�z|I*��}-t�<ޏ?�
��M�l��C���*�������r��'�
��s0�����5#�G�G.96��˂�7���O��~�`웿A*Ei��@G�V��٣��
"v�Z��q+$��f:�7L���8d�y�}'xe������Ǵ�ޓ|�gSݒw��U������:�sG]ҽ��@~�MO���\Z=�<��H�n�#�;UF��v��1lg����ލ詀��j!��q�n��=�laMW�Q�ۂ����\�5Z�*2�n��+�p=ś��Ï�V��|F$��q�6_�A�Y�]�_�l3,�����bx��6�M0p7�3�f�..��E�+#+�\��%����l>�� ���K�2.F־����#�ާ����V3d������kߩ�dk�}�v�OA���s���v�5rK���quuCf$U�p�yi�/I�.�>n�n�CPu�OrS����쌝=���ڃ]��7�8������J���՜���:��� Z�̀���3�lg�;˫�;�]�'��=�RC�VP�<fVJ��*��m�<=	��tʽ�s>�k�N�H�ts���Q���N1�K��&�Qł���2�mato���9�tr{wfk�}���~Rp�i�kN�©BU�����������(Sq@�`��彬`��f�+�c��MryA�����I��(fĂ�T��\ɶK����)ܷ��תE�7J����D��ǚZ�.�y�Y���UQ]{������$m�6��+��?��ŽH!��#4wm�ܵj��B�%"�'�Q�ˉsb��t;ز&'�q�:�z���W";F�X.ϛP(�E.��-�=��bYܿov�/��vs��d)z<�@��~���/�O�R+��)l�pj{Υ��n+���8����q�Oө�q�H7S�{sp�{�\xGM��=�o�wO^�'�yupϛ1��nB��Bَ�O
j�b�5a������z�L��r�2��Y����]ͽ����o�}nb���i��n��6L�jəgb@�H�y.�Ս>�a��%���ke�4���!g\P��!!�E��~�b�;�߽���Ε��$m0�M���o��e�S��Dv�� �P:��,�oiWG�������[�}W�s������t�VdƜz�(/(�M4Nh̀���z�ni���nf���˺e:���D��vqA�1*
M�)86f����fg]�ӗLj$����4�7F�8��GT��)���J� �+i�^SY7�J���͟��՝�k��^P�d7|w�y����F���H�K���вc6�o2��<����s�Yg�9Gٱ>�w5���WP��p��r6�2�ļ.�cgK�l�тw��K{��;H@��_��D����TX���'	�,�P/,ăǄ��#O4z�;z�=9�h�hV�Y��	'�:Jϓ��c��3F�A7�����yA�k�r��$;&�P�C���;�,{�؂9��0���Q6z�L\�Ko�<*�G	"qU�e�Vn�Ԙ£v`���>�B�"�w��hׄb�n���Jٮ۱��j�[�.U�����\w%ה3f�,��H@�� V�g���oǹ�:�7+�������qEs�i��{r�O�2$[�B�A��n�b/���o���������I�n�a�T�N��5S��@x|/�<�.^�"���o׾˻�0L�k�Һxr�݊�\	��/�ذ��~Ymٷ�?\6~#�X<���`��!���Y�"�	��c���!{�ܛR�Ó�Q"ƞ���ӝ˘J�`V��D�(��S]��Af���L��Ұ�{ڹ��M�/ ���������7�ڒ���������+E>ڜW�Ot
:&@���+���rUKw�B��#A.��Uch,�^����6�s�>7�nC�ި�����v���Y�fY��v���v]A���%r��,e�t3a��`WH�Ÿei���7kfy����<ڥ��: �v�{]��ac[�{}��ހ��e_���=;w/�Ɏ�\x�A?M��;�pv�5�a�$����F'_\�pm�ḇ��'����Fd]ך�7�2d^n� ��x+�Ӝ��}ҳm��e]�,"����Hݚ��	�)����?7}��Lr��%��y��.�)�,h`��QG�3�:��;�ǲ�e%pt^�j���ͥ�^��G.���h�ח���#�i��F��!({�53�����y�o[jg:�߿j�P�-KZ��	����ivv-��Jn���R��`ٲ�;7B)�:��~�/�T�����ˆ~$\}�s��`=���:����USJk�O�8�h\����M�ܼͯW�T=�r
za�a�c:�-e���Ǭb�Ò/)X�b�p6���ٌN$Bl�˞7��\F��M�����������ge�
qA�:qbVEۍ)�k�s�o��8�g�T�
��ۺ�s~��<Ǖ͢�&gj�Ǻ��"��C�<z�@��O�� 7���O%P��}��esMz�١�nF@�ݹƷ���)^%"8�[![�7�%~c�����������x���˩��ڸb[�6^�.8T�]����d��o7�wI�h�*ۤzaC��ԃ�[����{{x�l�@d���!ۂ�5l�ޓP;�|<����B(:e���)��{�?%!r~�fkl0��0Y�aܩ���V_S�>~Ln��i�[�ޏ��y�'t������7���xfIs^A��U�|����Y�)1���������"�S��˽X0cEu��m�h��%�Q�����#��?''ڝ��-����������e$ʧ����ܖ�fl=p?d�s������:4id���@]ݝ����F�#pEV��.�����ۈ����wW}�3�cy�Ž��"n�jbh�t����W[��bu�����uY��zAnn�^�hi���D���N��)�hXP��N�Z�b���r�����ɩ3�Y����0f���}��x�x<��dt���:�d|�g������%lӝ4�&&�1ޚS!��p�C0�XlGr�à��|����6���FM�`$u��"�;)�FC9�W7$�:��+M�TV��z�9�{s��+:�9�\Ub�H���s9,�����{�X&����&������q~LP�p$$W!�ƻ�\#�#6����34�m���-*Ĩ���n�����4���T=�(-%)��֫�96���}�Ȱ�1
��Qw�����B4ꛅ�ځTL�A#*�fdu=T�/:*MU��lt�E�R�Ump7�
�B*F�p�/�HmH�tf%끮��!��	�'�f�33.�%j����I�y�b����NS{��-eI}���H��k�%�E�K���+����;�xכu��B���}�?���Z���ﵰ����$��jЎi����tި+A�R�m
Ob�J�y��Җ+�0��vQ	�3��t4�pr�Z�V�c�R�'�_
�`Sf�P��ۍ�`ᬳ��p�����m\�n�_�t+�[5�;	-)jjwi=���UnD���]�S_�������ءJ�A�׏f(��'�n��-蝜g���98�%:{�G%�A���1�j6x{݆=����7S��B�bUO��ª(�#x���`��0���DFt�eW7u�w&�w��.����a/�L͂�{X1�!ŁD6�,Ү�=@����4N32s"۝K�[7�zF���HwӾ!s؎�Y�s�]S��U)Q=w�7x�f�l�\"����쎠�;���g����V�c�P޸�U���c���	�����1h&|^N�2:���g(�0_/TʝL
l�L�A�������}`��ME�qe��"��7ʶ��:�[Gr����[��7���>#>_mL��˾Dv�d�^���5	�1�ͭb�����T�a��C�UG\MǗd������)���?���e{3�n%����U�#�Z�(T�ӯL�!^w���׹~��,�U�/_s�u��&���,�����{S���X�|�FkV�x� x�6�f�ܖ�8�M�ނ����F:K�y�w�ԓ #t)Iՙxp�N��7n�wE�wY"��{V��-���E_r��/�������t�D�N|�B���+}1@�ŵ�Cq
��=j!�j��&��ݺ�|�ű|���w�y*#���|2�����	��;v���sͽ�E�$�1�i"�=,��;e,ܷS�ْ.���z�y�����.�=�ƴ���K���T����U9��Ϙ�׋+��-j�}u1*+���0��=���n����<�}+��.����R[`�٤Z��N���
|�|�wL.�
� u_%U���3ܣ�m��u9�d�<����TUC@%�<����olAR:I�g���r���*�UuiԼ)�c3�{���D��Řty���8��>�4�Q|�ʛ�)���
$��_vӸ�k3&j���{��_�t��:�����އ�Ur�Q�{����0�.(�ݥ��~�<�V\���gM�1�p�W���1��S�Iw�����p����ӱp�pc��g�C���.�D��=b�F�jN��D�>|��N�{ż0.I��B���H�¼���W]$�i
��ܤLm�����Z���!O' ��:��5���4���x�f�/�߻�_���x��c�,�߾����ظ��kIqM#Ď���]:m˫�uR�H����lZF�CD����J�`>�	�&�>i�~}	�I�._v��V��<n��Y�ba��LByYjI�k'�I�����w�(��W䶆+�5�v�x�j�����~�T�[�thP�p/f�v���Ev�hA�T�.��-\K��gB��-����M}h�ܵ�n3��{a�i(w$�ѕP�ɟm���s"��s�`B�BcD5^�(�K�������2�A�Y�=|zCr
A�]D�N������2�$��SӵY��ѧ�cX�#������3�)+a��	%D�|�2�l��R�棇gu�ELw��y��p�䏻E�l������E*�����k�#6*��&���v�G6A���l5?�Aۂɍ[#s�г������������|x�|||||||||~�8y��o7��������Ù�n@U9�S��ymG����d�w(�H�ɗ0��g�7p���!�S���є�gF9�1y��(P��VP�.p;0��wo<��Y��,���٣�#���d{��Ff�6'r��F�J��$Pqn^ɳ���kb��)���b;��%Emy��o��;���r{�nP��}�=���k�� 1˷l�s�wO:2�uЋ�9�rI��,�VM#!��ר��R1(җ�V��8�	рpz��,�9�<���������7���ރ�ct{4�#M����Ox��/T���|��o����fh�Lx,���Lk�Zo���A����&��5�Kz&���w8�_=ymXo���͞��x�$n����6�{H�C�}l������z�����rmI�ֈ����F#�z�k�j�Y6t�7��Y��^�M�8U�=��Ǽ/�咨���(����f�{��vn��[0�&���լ�Y�
Anf��V���.B�y�7-���KmPr>��'��W;�U޷4����̝}�u�w��ָ�^"�6҂&021{"�a�񈟗]�ـW��x�P�s�^\<��S��Pvx߶���9�C$^�8���k1W�����L�͏7i�
1���[���Cr�J�s^�r��χ�����C_s���އ�5k�;̸�c3��Z��erփ�[�RPMvڼܔ�m�ĩB[DdީZS��$���Ï(/�[f�5�\7oͶ驂0�ځp�a����[����s=������?x��%͌x�����އh`�"4L����vU5F���P� �s��JSdΗ���w'#�+&
�4���m�G��LK��C�ZG��8�(�6��w����(І�徘���������9���=�OѤ���/y�7'Z�@�/kdw.y�/{<RX��бj�S4�ZaKJbck`�N0��yS���V����_p��w^!P�.X+��{��=1�-;�
����4A��y��}׸p�/����7�=N��;-eRve�����24�I�m�XjηHae�sU;��9@�[�xȎ<G����/��V��2���^���K*��1�.R��|�T�����O`#�ܧ*T��odܹ����zj�7��@�ͳ�����c.���`��Y��\A���P��O�C̋�/ދ�"�ܩ^O�ܼثz/P�Ș����b�[kSaNE=l��ˬ��S�������T�@7kb�)�]膲wr��|�l�bP�S��v]�p��:���AƣN3iE]��{v�L��9����6k{/o�@E��6�̣�����r��W��V���z�����,�e ����� '.`W�`���x�Y�/R�`Z��QS�7���x}sʄ���Oɟ�
X)�n�)�\�NN-��޹������ӻO�|I�� H�
h�����A���cy��Ҕ�i1�BQ��4�V��tU#�����RT�-4���wP)CE
PR�4�P��h
�ih"h6�Q��HP�U���ք�W��Ԇ��P�'d��@iu���/[�jJ�	�EPV�h�MUAE�E�Bh}�KOQAml�i4%i(1	�F�F�j6@�5E=]z�w=K�l�h�:��O�ۜ��r����-	�
7#LĉL��N�L���D�E���TI5���o��;G�_o�u�z�z�[9�L��`�R/r�V��i�+��2� ͫ�)9��H'	rA	E��(xd`�DQ�( ȋ�4���% !,��		
0�d c���7�A�{�����w�0�8�r԰2����?X(����4y�Q� ;���tSS9j|ɝ��孝��Λ��k��U{� ���>�8Cz�6zf06�mI�1x���s�dU)�s�}�b�ˡܖג&��?L��O���H�\��3�^�,���J��Tr�\dv�~�厏�{yD��v��v���Z�i�s�5#��)�?�����We�����n�w��A���φ��{i�}�� ��g�g#� ��zbVڕ{tlvZr��7�~��Eh+����B����3�b��!� �����G^QF]�U�8(s����q�g��#`y��F�X���Ee-ysy,�:!�{��؍�Vn{�-�h�V3�?��șS�+x����u{�i*H�f��]2�e� �D�O�w��V*A���́
ҫ�����IAV�'�h�+������(��B8�un������v���x^�������Q��荙�[�p����tf�eoF�V�8���L��*s0G
>�<6k*\۰9����ؠ�0�Pe���F8yw��lX�X������c�zY�{�z��[��R9�w�����V�n=��d�v���e6�iw����B��b�\��U:�`�
^Jt�XNe=+#֎f�l�=�1r���G�/
�"���!�R��ើ]!�'�����r�;,ݎ�5�����/,�Th.Ji��p:�ԏip ���pj͠N���2�kqb����>��M�<h6ɐO.�pϛ ǀ6�.<�-�ع~N��gr��u7sd� �t���ZAĳ�$v��n���3� �]3E_$ä��#��=|c�dm#Ғ�X��tC;�St���ɦ[�ϡ�y�y b��2�^���MݕC�%z��4�-޵IHf��*3ng5��2�U0q�`F(oG�$f"�#����u/(�S<�+���Zq���Q���3d6���g����؍@E"5��<�E��]ytbzQ�~�z�1�v̎��C89�`O�u]��7�}ȟL�n�l�f�[�[�6O�oQ:�1J���'��-#��u�e��
��x���un�q����V���������㣹��|��@��:��'�YX���ܖ�6�����m��25C����:�3&z��=A��n���_}�+e�Ԭ7����l�Mf>RʇU�s�����?�����g�ܾC \�U|,��mG+�h�<5�g��yך�ז��@�%y�mO�t㔹�C�����z�Ż�ãAMU�"jw2�";E�J�Z���o�����~�����ٹ�T��KXU����=T��=^ɋ�Im�i��o99[����N숗fu��m5b�]H��
�����\�nڣ�N��O����:�OM�^�ʨ̞�y��B��G;�r*���e�Z�ѭ5�,�jH�cג )rMP|��N��#�-�<����S��wvu��}��G��Zoӻ)X�M��T�3���j��E}"Ǭ<�y�{[5>�2Zt�$=���G�\�^=+�Ը-/�β)Z��i��&���oEL�K���>~�u��u�䪂���=��z_lR��.�;^�o]���C����^*L�q�M���5���S��c]�*�8��ہ����铲���E���g���U��~�F���B��St.�v�Z�2�s3�o�FBv��$}���)Xޘ{��V쇺�UT=YrkIE��|r����Ю��A��l�0�`��o;��vwb#ǷY���a�-���Kk�~䦼n�7�����?�̀�\t�b����s�w��kmjQ���2�[��$�\�:t��EW@=Cg���������*ߨ9���s��F���C�������m�:����B4�l1�
�-�5tV՚��Sp�άߠoEظ��ɐH�%���lT���5�c�u�E�,������b`�4eG����oy�w�"Zn�_G-����4�zJ��x���ߍw�`	���>�Z�4<�J-5��.�r��Q��~��b��W:����rm���E<�p+ú A&��bf9�f䨭�^�<#_Y�]٫��ҭm�(*R�%��/-\K��gB��3���.A���pf���V���^Ɉ��grH�FUz����.i�[?���F�>�^ؠqVB��E!nܴD���ͻG�/(Kj�qW���*>��=]��ѯ��t�q%�w���!�����+&�(2^R����0�6L��B��sD�U�FވK�ژAJ�n�*뇚/p��?j��ud��۪� 6r�o�f6���Ɖ"v(~�܇��XD�|�Cr
OB��N���}�=q����ю��9�A�x
̞������������"�ݗ��e�UNM�b3���(oe���z��[S�G��Eqm���J���Cs��"�7ꧭ�P젏Ca�O�\N�ީ��\K��㐋Α݋GH��n{^�O�W��I���&W'�F`v����,���k��G6�^:Z[~rޣo�;�W�F$+Ή ��=k����o魅�s�(�-A3s0���Ϯ϶ �o�}ܖpH���p:�c�@�O�c���t�:"�\WU��u�H�Gt8:�.��^}���ߡ�b��nh>��eUdT��n��ja���L5 �g# >�p���dޣ��ޑN�x��ww����;J�
A�j}�����³Q��n�>o7����>���aZ�����u>&NƦ1Z�'�^����|ǔ���=SZ�.O�>�!�תç�����П}�u3u����R�e�t�F��٢1ai��OQ��[ڷ��FVIQ;��j	D��s�X�q�62R�fV�D���/=^��F>����o�c{�<�G����Ic��U�Us
�?I9�:Gws������#��*��r-Y*�^������������kNNٸ��ܸ�HMr�R��4�m���y�Z���FVH���W}R��ǐ�]Y5{�D-���J	=J��สU׸aUlXS�h?���H�s�j�n�<��A�0�WWP��e�}��ݜ;u됃��Uz� �m �NEO� T�q�X~q����9�fT��gCօnW�]'�1[^�W�J����u#Ll���UWQ��`��؍���M�(�&�2��I��N�f>� �{�
�g}/�G���e�O�辇o[�c�	�*���<�S�a������cE�jW��񻍯���~Ȼ+o�X,惘�y�������V3����ތ���j&W�T^$�7.tB뵃I�Į���z�줿��+�1�3�g����6�̡R!�r�Z.�9A҅S_E'�B&��!m�]��)MfF��
�k�ٗh����#6��X�Zq�X��+S��&ˌ�83R(���c��;�r�p)��|ߐ>��9�1�ek������O��Ęݩ��������s��*J��8q�C6|F���#���T>l�:ƲY�*hck˚fz�����U^3��졒6�nz}�op]����ƳfҪ�yޮG�������7g��UGl�'l�Pc�9�&�k��3]jj���Q�n0n��%����,ٟ��4�$� tQ��~s13�"��UE=��n�`���]��>�_�i�^Y�<xF�n��r�y&��\&�i��j����"��F�j�2�wB���� �*ϲ���O(�p�3�ߧ������g�2.}�,�|�z��p�m=|Ks��%�}��kܻ|z�\ϰ��AE�3�S�}Ky�xo��i[�qN�ǥ�p߹���7C�yQ뾉}L������̈��{��b�q꽽�"�5���Ƿ���m*{p1�����}�z&ո�r�$;����(���C�����Sײ_7��{8�[��l��Y�oo�7M,4�`҆c�i��XUh�#i\���n�e�ی%dT�P����š�,8G�L{D����6�������ث�ۑ;1�qCK��/;t��8}��ա��e�rEXn�)���\Q��t0z�Yܘ[~����9clʯ_��*��\l6�}k�M�j-A�t7�����w���~�/���=�?{x��I�X��d�'I�掭땤����B��l��}�YA�vU�{!�w���@Ħ"���>�⹊m^n�����x*ݓo��l$�5���Bf6�8�u8{�cxg`�]b�4:H�m�S�=�P��St�h�V�t�c���t�ό#1���?�F��߳�5��m��������8M2jx��E���ׇ�<)�{u͒9��|D����/���]���M&|H�c#q�O���3�ޫDR��A���:�cgsQ�qc2�op��y�l+�il5�T��A�>��f����x��.C�����/߀'����.ާc�ڵ�̈�ye9�c��QwEd]�Z/��rF#|��zK̚,�,�	�b�"6��û�0#u!SI��h�-�-�ܢ���{�� kT�G�N�5�s7*v�/U�O4��V>�BQ�;��^ѹ�lOpb����>7�V��kF�	(W�@{��{�y�o�����$!��^��݆p(wB�}ުGҶ\e���,cКi�{�����()�JB]m"�ԋ�s����Ã6�=Ա��ʷ��qu ��@d�v������\�b۹��6s>�<�-v�n�{c��b�mCU�Z�� ��~�&R�IVL쥁�.T�n�Vvut�E�*���<}�fBP:؈�k����%l@�m��<�����v�Q���Q¨��e츉��󢶧���UŮbV�l��¢�z;�����k!���S�v��n�I��Ju�x6�Xmε�Jb�4\�^}��so�S����a]��h��Y&��+�V��N�>w;=:����&�A;���L7��o�o��3��OZU�.����ڪ��^d͝QT��r�wp�]�]����2e�I�sk*�[7nFT�� owR��cSæ���;�l�3�����,�7.�e�h{��ڱ�����0r�\^��8M���uq�e������g�"4�O���?�3����UE���[}^�Kh$MM]0,3�h{j5�m ����mI�/.f�y0��.=�ԛ����O�x)W~���znذ�X]����:Clbm��[l�ǲ�d��Y.=Y#��Ԏ��e����8��Q��A�k��0?��<�5��0��bƶ��3Ƭ�=Q|7;��	�j��0;6��������6��2J5a5J�~|�=h�>�Πu���{x�
�7�`#Ք�lS�-q���x*4�f���fa�A᭽Y�
�n�����8�U�6m%<�3S>�@�ݦ����L��B��ֻ�:ѫ���ZJ�G%S9���3=57��ۗA���82�f��`�ÛȾ�`�[-�ݒ��D�^����zw�x���39 �����xӑS�En7 }����>�_������=������������������������΋��{V�S�]�Q__������̙t{�i/gk|��k[�ѕ����gwЃ��؛�1�zj�z�{���zK����mƻ�G��w7���.�K���/;��L��\w��T���"ޤ�T\�&*���j�0�Xj��5�{:���b�$��j� A�ǏH�=^����0
8�i��ز��l9��nk9O��~O�n��ƅ0����g]��r�Zo�M�<�>�13���:�r&͘���h�hM`(��c+�U����3���t�φ��o|__6�T�Nev�Q�&]֬�W:��JS�"~����XEG��M��g���=Odɞ����."D%�QN����H:�	4�5���ӛ���<F�8�)�Y��+�w�ٰrx=�/�tŻg��e�V!vs���r�tةFjf���WSd2�/u�����р�/6�����5��e�S1�ׄ��L�vp��T�~�r�57�+d!0�L�YuI�4 ;tՓ�|��o��bx��凸=��\Iؿ�7Yұ�э���%��nExL\2�8�K`][N��?
yS�����azԮ]C=���Đph�nk�J��a O�22�h!��`�@��<Pw��zi4U�&��� ?3�θP�+6)�ۭ6�H�]U4����䇷��7���}�n�w��v����FFE_n��M��#�EY��X�7Y�u'T)"�q;0i-��UxۋAFw��ߵ�4�v��B�m��h�(b0����� 'R���Xu��}�Mc�~rv�_�,&v���{�U�I��q+�T�[ڂ~S�OQ/��P��;�Z����הql����+�p,�yACFs�X�t��N�=�aD�Y����]��u@�_�7�9$~c`+�¯��m�R��}FR �OY�lh��6���E,��~��o���~zn�]�y|��[�i���`Ub��w6kb?l�}�����#8���~��N�,�����D�P�(n\�V��5йDb�:(���-�`��6r��k	���y{�$����$��Ĥܻڙ�K5m�a�ә5�Sn������|����@;�;���z���;S����y_z!O{��H��ٜ�վ=����w�#��ŉS��T�&�mz�`D, ���h�[�U���Wk&���IVV�eB������wKz� ���΁n"�	T���d�	�Y�g]����V���|�5��{n�ѱ0k���r��X���x-n���8�ٝ��������A�.�>�M%����]��XY�]����������OO,��<ŤvY��4z}���ƚۓ�� ()�s����G3;5���4�4��Wc����RV�A�?;�^��6L���=�U���;[�u��i�[W*�����KL^i{�����T��fW�$�
)!�'�D�Q�Ѥ�i��+Mb6ɡ1F��)h(z�V�iB�IF���ޤ�߳'D[)E5��4Һ�04�X�td�4���ւښi�����i�M,M�S��m�����[h�T��R�@Dt��ܝM!]F�Sԁ��-�i肋`��
��i4kZ,cIlLQV7v��:6WA�
Z�)JJ-b��=u���u��Ph�M+��fO�]AZH��-��Gr�@{�ĝ�JPiht����ZZPSJQE=IԔ�{��I�.�����4T-U:ӶuZ���)����Zkl��4m��4{ء�����;cF��k�.�Q�X��lU2JD��>G[SMcϲ,���=vD^�S`c�o*�YҦ
;:��8�9u&f<�&���`cd�X��8�L��BISr�{�_wlK�{��*	%T�:�ԍ/ �za!���� �{"k�ooSgsd �Fl���Ƽ�&I��N$6c���A�hN��c�_pЂrT`5������%M#H���1��srz���cLD���t���=�C�9�!l����_)�[֑��\�-�{Q�U��j�N��{��5p|��:����`z��Fɮn�������X�}�˽K�1Q(23��Vl���p̀������H4ff׾�m�h�/�K�'��懟�W����c6�[x�������I6���a����0�9qC�	��W��ԏ ��c��9�e�J�\ϵ5�z���;�Mg�M�T�<�v���`p�%��>�c�ɡ�&�����;�[�ؐ��7�����Gx�^^Ğ<$� i�_/�!>��ɮ~˩хu|��TK�P�`���-	�m.�XW����	&�-��(��n̻�ń��鄵��f��]��s�2�P�dH^�Ï7��&�.��9�w��zf�@#6�	�P% ��Ac�)��:5�Bf�yx3YYR@)�k:�,>O�XNi���ݣQ5uC2�����/� �X�����sN���ؙc�P�mes=�����z	C�OW�l�FE���6E@[Q3�������p�׽CH���GA맇4tǅ�0�,�hW�Z�.r�c�3��R��r
�f�Is�t̟t���g@��#M�9��Y��ut�S���
���j[�q��)�3��G�~B���M�u�Y--�p֔sa��!{cc�Ȏ
�p���Ҝ�nH�з��r�m)�bN|t?rT���Ɂ��ߧ]����s���*��h뒨��!Кp��mD�Vq\p��_��x�����0��
�|�H����=^�J�p��t��.*��؉�4��:�����>m���<|7�����EsYmo���{�j��ƺA��ƹeO�㺟?o�-��U�ozh�`�f�a����Z����9&��Y���=�9l�g�&���J+#ۤ����Wv�鯫�ѯ��x;Gzf˶V�k'�ɝ���y�|q"s�O>��W�]^'����]ڻfUn���:���*����=Czz�n� �˵N7`�7�ۆ�,f����Q}�b��x��M�0F�ux�՛ULg��H�r���ylGs{�cQ�a<�!}g:�u4"�(�ޞp�Y��6�M�U��y?M��a�Yq螤���/<pse�C�v��sA�<e�Eظ�D�2d�f��n�ɇ���.F{���S���Y>�n�t3�Ah�
���oy�=�O�z�N�4��7�^I��E�đ��II�����/ٍa�ILm^�����1[�){�k��i���O��h�y4��S�O�;��$,K�����v�b�[��QF�*Fw%�[�)T�o%��/-M�9�ZL��^��Y���3�}��~�.�gV��ƈ�!ew$�֌���۱��^9�LT�̺�'��o[-�r.�{�w
�.og6�@�=	����,�Fc��K&{k�9[�cyUe�n��_.�[�	�����l�	J��d�Ig��ՙؠs�w�q�wp.c����c�5��o����UW�"������0�^ŉ�r��ukC�5�OX�E`��H\��[xc �ux��x��ї����x���t]�;p��bg���+.�E��������W��E&涕�W6�����P�]80sv� 7�zvG���?_K]:�����`�萸u����o^ܲ&�b�>�x�n�s��w�M�EXn�+7g�����S�����=	��19��v�۹�0U�ܔ��@V�$wQ�i!r~���w��@au1m�����ڲ"�FJ�A����_A�����՜v��bU��	ݐmq����e*<̆�n�?m�����a�����eM$3�߼����m{*��[�XR�X��;��ٔ&e?/!��q�Ϡe�}I��:> R����v*�c	
�2�w3�
�@]B���s�g# >ّ\��M]�T^����1;ƛN�����u28������:�k2�0#!��=����۽����'T�����g9<�$I ƞhv�(�ſ8�a��cX0Nn}7��o^M8��
����ض�5B���J�"Ւ��rz1v �k"�����9 ��P����R���h�Ħ0�y�]w�>�ˈ�{g��[�<��)�v�n��R{�m��mn;�����_�Vm\��7;|F4�����+�{)�F�F9n7�1]��;zH"UN�	���s�h/X���p�,n�ިv��������c�A�c�V����r�JB}\�qRԎ7;�e.t;�E"�}G[�N��̵�����qk��B�h\�N����Ώ��֩���.���p�&֬g}��"�Mo��
��.c8j��Mp�����:�����׮��+�$eW�;UcU��V� �NE:6�ML�ּ(�f���<��s���@�=!��A�}'���)�?Y�z�c�V +�/"������ݝ�];��ȸ�f��z}�I QGͲd˨�21�Q3,��Dօ�]�X(�o�b����6�ĪFQ���`,�Β+E�1cp�f�g=J�b�[� v����zz��kbGZKʆ�
唱��]�s)��.o�T�!"�\L7��i�Űg����Z v|x�yZWa����>Ӥɕ�5Y�³�Fl7�n6������7H9�|Iq�V5}��y�CE�
57p�lex��e�W�4uv��Y齾�Q+��{/� io����-�4r�7�G-X�Pd��!V������P��X�{����Ӵ����򻨡o�{��F[�	r��6e �j�t&dD�
�!t3��0��w����/-n��/m���3�8N�}������:q�)ymO�Gd�.������0�w�{�X쇱=;������oH9s5OL0waNGs]B�C5�/��=$w$�â�wRƞi���ƑY|/{����b�B��)��ݏ�;����{�X�� ��f*c��Kl��i]�t5��v�D��cs36_�<�6�r�W��
���c:
����4gU��j�_���qm]b'	K1>�M<���7�Y�:��9W�*�8��3{x��}'�����Cַ#(���g+�ݚ�{����W@�f�I�<�y���j�6^^ۤ<�P����u.�;�E�?`WݨP�]!�>6�4\ęk�[ԖE�������뜍��u@��;�� �1�P�E�V�{v
<�qC�W��Wbn�Ll5'��*�c������eח���koɕ-�]�����b��À?�r���öA=C_��F�@	��y:�w%���w�n���3C�����i��'��	Fv���L�;��n�a�հ/0�i�U�
���J�s��'	᝕�r��%iQ!q �fJ��i�Jb��k��/M�Ab���f}+=Z\�Iڠs�ԗ���ߋn��cD��G,�����_H�!����D.�\g�����h�j�X�Tv�\%4R+��s�5#&��_x�Լ�yg���[hH�IZ�-|�W��q����ž͏jY�_�&�Ϻ
���᱇۴��Ǉh3Q4�&}�}��k�՚Ou+U��u��4��T���4N���[�/h]��p�&��gG�6����tl:�wg����6�t��b�Wa�	!�L�]�#5�=���������;REwN`�ʹ�/��g��wU~��d�£Qdp����Vfu���|��/'�A{�w�8��I�p5��}�����zJ�@Y1��d\l��y��uͤ4�^"���TD���{j}�O l5�3�,ͩy�MI��'����N}��tSدz�"+��'j�雅D7����h��6;n��@�z	��ݞ��\�Sp�թ`��+--�e����*�H�lc{���'&1�A�6�U�hTY����U�����0�V�o
�p�Y7��۳������b4�����R��S`��ő@:��F�b�|��vx�ts�`�'9���;H�&�w$�]ݹ�E���nl�a�=5�ss�i�q�7 9"�"�v���ЛS=V�R�2�x���^�}~=�H�����8:�FP��u�+���nA��O�օ3�.�z�򶻻����t�F��*��8#2�	�Y��n�i����/z�y�����$��*ۥ,�v�_[��RL��a�u�
�{:tv�	X�Ք����wY�|�\���;[n�����e�ocv�'���QA�0��OwP�;D��:$�muR��uS�:��vkSU�N��#Y�}ʃ��"#�+}���q�m����\�,�=��o�.�8�*A���g|�pG��r ����������q�>�b����oL^6��^�Wu��kF#����n��u�10_b��n`�ӍW]�5���P�8-Y76_�H<KeEՆqh6�lDQɹq��Y1�)vĽ'�f��sV��eH�T�,��Y���7J��L~��w.2���?��~w�-�J�.k�k��qO�{n<s��b������X�ӟ?ߟ��K�n�n�Q��JU5���{�ܝ������:+5��G[��4҅����x�H�4�G`�;�#!��3Hi�V���uv��ETy�K���(����o,
�$r-��F�l�@�oi�M�vឩэ��Lو����Ƥ��o�ii,уZ����\4⵷�9�'�4��eY["<D�3/ûbY�^��M�n5?݄�t �ˠ�3���'OZ=w�4�}A�U�����4�R��	ok����p�3	�)�!8~�G�Q�$eW���r5[�l�t�S��FVq:Ϙ��tލ���Z�ɸ@O(�t�U$��~�t�M�<�I���Ƿ�X������	`�����/@6�'�p'
����������}|�R�y7=R}]K�%3�y�w;Cm?�Fς�/p�|�ג��؞A j_�o�Y�y[iLr�s
E�����/l�5�NƸRͷg�ɴ����a�s��ɝ��V��7�hVm�e�Ǩ�eNQ?&]â(d%xTZn��W�j�:�"}�f/\J�E��*i\�O��D�C,�5��X;t�4�<�?K�0��F��y��l�g��_(�kb}Q���e��E�{&����YT�H�Ӎ	0���c6.�닾+�5�2��qar�j�Dm܉^<zM��׍(5Y#i�z<Fl�ހ�������B[�j�f��=��A�i�>���D,vz�8�%/����ؖl�<�1o8����Tq�g2�'�Q}�D��_�m��j��]"����nbf�P���Q����u�z#̩V�	@�ۖ��zL٭[���:����Mq��0_@xI�m��^Y�I�!HiRn~��]Dɾ�G_f]��sӜ��X1 !F�5u�}�wkE�|�s	��y�Ј��dq�t8��>m̎�z�ĸ�L�]������� � Wj*������B��	?�E�tG��=ϳ��"�	F`Y�f�@�`Y�fE�VB�eY�f�FdY�fQ�B� �eY�f�Ve�	�d aY�f�eY�fQ� �VB�`Y�f�aY�f�FB�`Y�fE�VdY�f�dY�fE�e�f &�FdXi�	�f�`Y�f�VdY�a�Q�eY�fE�Ve�	�fQ��f &�V`Y�f�V`Y�}����d:�aY�f &�eY�f@&E��`Y�f &�eY�f�V	���Ve�fA�dY�f�F`Y�fQ� �`Y�fE�eafE�a`Y�f�`Y�fE�D�VaY�fE�F`Y�	�f� �Fe�fE�V`Y�fU�eY�a�	�fE�V`Y�fE� �dY�a�I�	� !�!�ϼ8@B Uz` "0Ƞ��� �R���=�Ѐ0�0 0��ʪ� C"���0�:\�*�2��ª�( C*���2��ʪ� C�XzV@UXaUa�U�`X`XdX`Xt�VFF�=C�,0,0,0,2�2,20,0,0,:2,��̫03��Q�d�/q��{�=߯�j�(Ш 2̟�����Ϸ���A�_���?���?��<0y����|:?��&�������������
 
�������@D�?I*�
�����`�2����K�����?��@��~���?�����{�����@�!>�~��?@�v+�UE�Hi�(P�T�D)@B@��P!dA	�� P�IBT$	@� Y B@%TFA ��U�!Ua	UX` �U�E?j@*�=������~��?�@�A� �@)K��<�������AA���v�)����P\���=����u�O��#����z?������*�ȇ�O��z�i�Q@~��C�����>�"����G�@|'��I���_C�OǠ���P�I���<{1@vJ���?y���?����v��*����'�u���>ϯ�����w��~A� }�O��(p|�� �����������A���>!�)2���?`��8?q�?��=����	>~�J����S3��~i�?�v��A��c�~�O8��AW�l>��A]��>}�?�~�������e5�}��Pl흘 ?�s2}p$R�]�2M6ڭ�-����V����3Tkkf�Mk5ll�M�l��Y�e���B��̰�L�iHե�������֋&�[j2����V�٪56��T�ڙ��m�L���[j�m����eL��6fЕ�V�m,�6����L�mZ�Z¨T5h��d�-%�(�m��&JJ��z�C��a��Sf��5m�j�V���f�M5��ie�(ųj��[kFJ�F����mm�5#J���J[3E�Ō�"YK&��ڥ����ڥ���Z�d�>  j��{n޶��oW� ��:�����\�Mz��V�ǝ����m+ݮ������yܼ��e{�׶��ly8��[jo8\�]�t��/zm�ݎ��Y{�ꇶ��By{P�T�֭$b�Ykm�^�   �c�m�%�Ĉh���xz>����B��-���g��ƅi�l[a�C�}����C��}}��z��ox�Λ��w����;z�㽸�=k����ݪW�{��Ʋ�lz�w��ۖݻIM̳AK	��'Z�i�l�e_   w��������w�@5��n���;���wz�^�tѓ:R������{�5]��+]7j�PUo^�m�{��]�������u�z[kׇ��a��o ��֭�w0.f�A�3O�  �}
izW��'v��JzU.�����Y��n�������s�z���Z��@������m۹݀�u�\����6gj�*ڨ'VJZ�jͬm6V�ڵS[&�_   ���:4-,uN�;:����;���4hL�m�\R�� ��k���5��8��A�� 5v��t� .tªZ�֦�4�h�fm��   ��w8���n�t��
� �c�WD�f�+U�軣��U,�u�������+�[�un�@�um[m2mj�X�,j�l[I��  ��U/CI��� Ws��u�Z�k���*��0V� �}� �ԸT��]z�@�U�R��W*��&��m��k3-)k�  3� ��}�� ��p� ��n  4X=  q� z z�h  {� yׯ ���  r�ƛI�VT�Z5��ڬ�w�  �  ����X wkp } <<`� {��@@� @q�8 s���	w` P�&��@��,[f�M��kc�  �x�  r�  �� =4�w=: �; @8  �P�ڻn N  {�m�@ ���R�D�=@ ��$�E  )�1	J� �@S�����   i��� $�JD��T@ 5?���������s�����Gh����.��"̈́8`�{m�J��ˌ_��UU}_W�|�����=Uk[oݪ��[_��Z�ݪ�km�MUk[ej��[_>����;��?�
_��ݔV�_ɷyK2D�(cSv��)f�$N:F�e�>uVڳ�$���;m��7��d���b���MwP�{����:���02�h�ݧ,^j���Ko;�uj��.��y�8om���(�Wj�X��5ʛ*�e!h��M�H���$�SL��#i`�D��`��[���YyPKyZ�:p�峔�9WABw)d�(A>�d�HйW�~��;V�{XC���V
/)�O5�m�!&<8�|֒�(;R)rP쬤.^�kMIJ��!�9�z�HT�n�(��Q�Z�RҢ��B#(��i�;]q���Ei�y�6�Z���j� ���n*�Gلh4�-ٻ��)�fu�������4�0^Su��יD^�wSpԭx���4�t%�r�#c���FDJ���fQ�`?�G��^��N�� �E�����t���3o�m��֧�0���A�{�N�%�R�2�f<n%f�jٶq������x0d��e�1�"�HѤ��-�m=��mLܽ�)�i�TZ+C�(�+/bZ��.-��.� �D -��,^��n��vYL^douػ�GYW�n�ŏ�wP@el���� 4���J-�i��5i�弖#;��%�m����;֓�ܣb��/$lvJ�t�����M2�j�8
�1�7j�*�5˷LE��	�-I�[1�Dirl�"kF��IF�~�pCq�e ��RU*�Ô��ý�g�V�K$��I���q`n� "���^�r�[.� �j0H�r[� �N�̌�µ]:���4�-��a�Ȥͻ�!��+*J&i��/qf6�E�h�hX���CSP:ߘGw�u��袴�͈�JFf���&�!��\�Xi��aS��5��r��l��JyW�����-��^���+q0\5�)�;
e�b�sr�(I�*ܣSIR%���*Ċ[��_�w��x�p�1�@��z
����ZP�Ê�+S�E�w��o�䊄U4�� _�5ӡ�Yf��E���Ch3"j������v�2Q�Ɗ�c.�J�b+yC7�5�N�ԕL���ĮB�s �yn@�T�OH�9��#Ke��Y���v��b� ���I�-\˘�9-��Y�'�Kkc��M�eE��V�0�e��r��A���&K�hKR-si8k][�u4�G����ޗ-�A,k�X�kV�(f��7��e� �a*�A̻4R
�zV���a�	`^�s	@���l-���̣i��q�B��
�[��[7�^&�dM�j�+�w&cc^
a�U�G.ʰԛ`V�+l����d��R���1�W��O3'�bgx��.�j:w�X��\�s2�Mi�1fl�(SsY��X^��m �RP5-?�H����M�ʻW)+�R�<z�!1P�:S��1��7u��r�G��Ji�x�ۣnՖ^�"�O�+ch(��HْL& �D�D9x`���.,���C)ˬT�V�A-ϣ&��wZVIp0�^��l�J;*�MwmP���٩��Ҹ	,�h-�rRHS
=m�j�~����bJW���T�G�C��J�p�%������5�*�Q#���r4��5�4wQz��F��Klw������L�)���4��;Ƅ>��?;fb�G"K75�P�ں�z7cCl��dˤ��̻��nS��2��Nѫ1�Dt�7X��+��F�;i�e��Z�A�j��q��LeVm[�aoq(0*3+{)b���4��1	�X.ۭ7�ˉ�Ņ�[���贠us ��[� pm<`�F���OM-��sU����4H��@��3A�H&c&�%5���V�+G;�J���YYՔ���,'�kp:��mk[��`#AU:�f�M$��0�����g�Sm�M^�U#L%D]ۭ+�w��I+C��@�Zb5��|����i���3�Mg��D�p��Y.���wt5UH��U�����(]���v�$T^�*������� R�W���Ej��fR{uu�QX�[��l-�6F���1w��	�-�n��5��u.Yi�[��D��=�jl�lv��,�Ĭ��Pd
-�raf&f�vR��x˽ӁPQ�lѹ��Vu�љH���4[0�+��㡹>�;�sV[.�B�t��ԭeM��D=�������w�zRW��q�A���5�� �`m=�@����A�Ɋ���Un��
I���[Y��Kw6T�3����`�t:; cX�{G)S
:��'�oFm!����װ�1V7��n
[,s��D���b��\7&\I�@KBcB�R���V� `���wlPʲ�Y{H�y��c�d�3mc#Qչ�m��,��(Ŧ�W��3w2k1ɪ�8�l���a�E=�LhznuI[y�*��yZ���7�~�V�H$��3iJ۬�Uk*Q
��8n�*�e�رʖq&�
�«-nk�,8�ql�x�)���-*�e�[P�i]�u�t�h��1��!��m��׬+��������J���� ��Vط����m��f�5&�"�$t�jשT�ÈT(��r�ʷ�'bn�Z��-O��TYu��԰ѕ�ң.S"�o�Rt	T.M����פ1�Q�W+>-����t1�Jf�޺�����f�ݑ<�%-0e\��`X�͹%Z�b��8C�z5 NH���
"����(]n��n,j�Rm7sR�Q�WZ��md��N��ԕխyJ��A.�v��n	j��b�J�q�J�IAv�P�Z�;����>�(%.@��ݲ�zf��vy�G(k6JJ�պ��՜�xeG,����V�vg]f�4�ٷL���Jĭ�h�7$��ot�XڌU�u)ƾ6�d�`��F�eca�ܦ�q���,��ڸ��`���OsMc�W6�X���UtpGt�p�l6N8q��S��˫vw-�Mm�d�5��CR%y������f�vwT�%�� LL�3�KLXz�RP�l���)Vd;x+^C��\��YL�X��MwI'�%\�B�ً[ԑS�l�ʸ*Q���ծ�5H�/-$+C.�^0�\nS���W%$L.ͪ���tr�#�� � ��ݓ�r���F;��&��-�ָ�- �?���I�G2��hMkoM����6n�r��Ӛ�j'#�����F�T6�[���� �6��J&k�ݫ�U3dmL��u��6m,w�|f޷V�+u�+��J$S�#`e��R��e�e��˜�1����Y����1�kDr
�b'%��h���ǂ��*�RuC��x�V���L�F�B\q��tAsK��'@fl��x�;��*鼤�7��sd=yn'�2���m'x�Iܖ�#t�{Y.���ܣ%�2�(��-a��C]Df Fݪ ]��^�h�1�#zoT!�����	N���M����L,W�ͺjVj�ٷf�{&�J�5�u��%cp�1L��^MmɈ���l�Tn����7abqڙ
��0�q��O�D�i�����Tu�\����0���8��i{b���T(i�lL�Xy����,��]Cm�;khU���{��uDZ%k�q�LM]�+*���J�:l	a�нT�J�dQPըl�u��ݧ�`v� �H��5�Ƃڎ�!n����˫Z*f:4&�S��nm��5��R�#Q(P��ŷ.%K&�Ve�������o1Z�.��F��VQv2��vSo5A�N|�X�{#�*6s����զ�T�L4�/E'�"��e�L���{��#-�߁��uG2QKj�-+i9��rf˻X5	 �l1W2�ܫsti�d��|�U�%�U&�q՚��:��dF�(���,V$UnU�,�ݱ��M`���1Z֤RCRSV�/7��rޣ�ے٣�K��j$�f��V���Y#���EmRĹ6Ej3��ʰ�j��,��yXJ���Ev����W�MBk�h�w �n�!�Tn�%sNեA%LIc�f`f\'U�Mʊ�;Mò�\3�>J����z��Xv��A�%=B΀]:�z�Hq�6b���B����e�R0Z҄if\X���L�8ɥV�H���#G(�VT�)�����
��4FFM���*x�:d�*M+`PM�騥��\/]�����"�Eػ��4N�
ce���9k,LGE�32�,탬�cRMD�0�8�-������e&�ek�bQ��KeZQ�cI�H�Ҙ�u6�n��m$��NlNMH4��q:�K~7M�oɂ)
���dA0����j����k�x��xM��l+����T��Z
*u�f}��L��#�GQ�
VS̭D2ɽ(]BJ�Z��EP��֒�YsݔT�S{�ƀ���m�k��5�G{6]mh�iO#�R�!d����R�d���3���tACi 7iI�"@IڹWCA`kt�i�V��N��:د)�fԽ��H����X��6���8�d;�nãP��KSY�%�0���Ƈ5�KQ�􍌙%h���6��nc��3��bD�^ʍ��,�^O��GC��k�fi�gc��`}a��㼭Ksc���4�s`�S�@��������/SA�	b�]:�j�A�Eͩ��ɩ,"ں�ڙ�*bJ�9V��yn��QU��^P5,T'd�3cd��"�Ϙ)���(����.H67Z�յZF���5[v:6+��x4-�^�ݼ�&�Eҧ(��ed�S��	�u�!��{d����"ՄR�%�60�+�r������ܼ�i�W%b A�������7n5���l�*6�5��s#�c�J'!h���h��0�˕q��h��ib ���í��w#���'��EdS1<�z�g�@���(�7�9}�����zh����$����:�Zg�ݽoM+ŚE�_f�vnʹ٫m핋P��)� �y{��Z�S�
�df��"���:�K�D�S�&��w(9I��VƝ�R`#hP�Bdk��E�p�v��L2܎�e)6�Z�(�jY@@�Q�����)L	M)0*4E��ˇQ);n�n��Z��p�k"�J�Ɍ ����՝a�͊�sCrS+��i��x�P�Z^
�b+j�{��i��=&@k�n��NGh[��l�d*{�Y�"kr�q����ǌdla�)7�V�Ikn��
�A�N&J���#ۅ{S8U�E�*���������T�FƄ��P�o��b%�i쳯(d�p�[��������N	$�fQ��5��Q�U-�ͼxoa�wk	�	f�j�S1�yV-�u�BM�vn��6
����g�z�Ԙ*�E�蛎k����x�YT�Cj���XLjR�`����x��SjZ�渆��7^�]��J�W���XF̛{d�Z/#�l�K.̻�k�osN�YZ��&��bRaݫ5aV�Sh��M�Yum�l�@Ns�r�O5�%�J�n*��I%)�����QV����d���D��e�ڽ��)`宋�wB<���J4n�@�O�5R�}�T��H"�jR����2JrTc2\
�b��{���UMf	s��e[�-u�H�r�;�Z�@)CpڃU*7���ăD��r*�ӗS0#�1a�/J����V��n)�e�v�ֳ��K@�;F�X�t�v��s)�t���IR�n�#q��M�X�(ݝ�N�g'�`�{kv�<�����D�蠮f�#.�=��{jS��L� �����b'K	�C"̷{�R;�8#��)��-(ێm5x�h/(�1�H��a���f��3��fL�/M�W6��i^4�=0�iZ4�D��`+��;[��u�X�H��Z�ʶ��ͨ�e6-r�E�7b���7)��YGv�����%��з)a��p;�¨�J��Z�@���hݽq;�o)�3E�*-6h�N�׍B1%��v+2�]��Q�wt:E��Li�4֧�w5�xm��7g�غ6��TRf
��w��ظ�i��yH�$��3TN`Z�Ɛn�Ii�v� ŁB���Ygq�b&3l���G��9�������K2�M�w�k$'b�J�đa��H������[am�&�[v�܂�Ӥֿ�5i^��[�9Eػ�0���ˈ��Z�z�:��wh�m�]�D-����:@�0���A�R����Ơ���g֥ ^͑S�y�ko*!x��]4J�;[@	��^�6R�b�&XO30�yL)������IIrݪ��[i��"���7tJRȳu"�rҽ���ʒ�"� �J
��#2YK�&f%�EЃ�6����$ۄF�K�Z�M�e^�Jt�R��gi]ң���Yt�]*Z��(�w����l`gK��
M�!��0�$�,��*V՚�w�m�r��5���ٺt�%���PXmJ�b���Bc���o!1R�F��3Kbn�Su�\��5BSp$�F�w*e���H';�!����EJ�����t2n��쭢�Z��[ �qQ�v�ڦY�.���S��[��Mh��*�C�n�Ї/5PL����2�*��y�rܠ�\XحI�$�+ ����g)���c(�9r�F�V5�e*�R�y1��	�V���{m�� ����2�A�#u��Uw6�l"��j�]Fh!��f�@�ͶpJ��M:Ƴ����\Z�7V�c.҈Q�d�.�L���7g(\��nYp=�CjS��bҳj˹Y�c��Խ��b��.��]#D��̗JY{�ko2ĥ���X��V`֪�˶�hȥ�/N���66'�,���Vi�s>�K�wt._��{�}%--��A{�|ޖ�w>��v��S�ܮuu_:���+���9�諸b�H}WC6�*�R�m�.]�"R|�k�؜6�g��^d����;׏^اl�m���#�_��R��0z]�5a��{]7�9O(v��_r��n���j�3vd�`��V!��nB|��c^.��$U��u�uμ-���]��9N޾!�6�`c��'�p���l%�nt�W�EXl��;V��Q[Neʅ���u��g[��`YN����Δ�^r����o,�ZPj�)%n�.���H�z���ףp���Y\�/�n����]��8�o+*�%���<���U���R���J�l�y��F`K(*��uj��X���W[�k[�̇�wyQ9ʬl�.�\��v�+��(�6�M3��e��fh�a�]��Q�1J���{Ɔtǜr�`mG�u1G#7t�O���uۦ0�Il���b,=6�8d�ړ$�@�)���p����z�!o7OF�N5�Opk7�7`��볷��g>0H�|�������T]��te��Z��Xq­qj���V��yøU��U�I}.�r��FK]w����蘫�>��oz�CHu�H��m�U|k�]r�D���qN�jW�^��\�t�1`R�R�=Zh�gw�C&�Xe���W��ެ;���0h˃�6�g�'r�vw9��T޵ɑ����X���Zc���D���*Z�5��'|~
3�kw�θ2��T�ۣ��s��;A:u;(ңhd��Lkcֈ��Қ�{�v�c�ָ�#��t��huh|!�P�0f|�J��tw���I����V�Z
��;���u�r<��]Q�p`�ۧ��n,���ζ亽������4�PV�z��9,t�,A"����lNa�.��l�b�a�k�7�t[4mۗ�����qf�5��ILe��(D�_:���6�T�%��x�������-��H�L���W���c������Ҵ�oZw�P�����h���O���R53Q�}PU�p�C�	�sz�m�MN�Z�_M�;s��ʯ�^�W8�V��*�&�Zm��+�R�s�7�i���F�v�=�(�j,{m]����s�驹[-L�)��˓v�WTۭ
�һ
��������dř\�q��Ne���(�)-Z)����4�ӎ��3��������Q�O�R����
�����c�-r��VBMㆭ��&��tMIfS9�r�9670��H�N���wXe�zzB��vWL�r��d ��5+�����
�*Cd���h�,����nU�RR<t��VmS�ȇb*�����O�^`��)8=��wʐ�Y`�� (�� P+E�#ʀ���e4�ǣ�F�T�ۓ�F�������(���l�>A=�$<��T�q��'�zz�}�nT��c��ܬ��i߭�΂ڑzQ9�'o���6�
.}�b�	��o噇+E��U�K�q��u�}�����z��Å4��M\j=��l��T=]T�m��M���%#v�i�gG0e���ռ:�d������� �i�Ȑ�'N�wŃ�u���qf�j���8��v�m<M����x �:�gvIq팔�82��Xo��Ʉϕ�A�4J�g,��Y�ʩ�E;��`��귨��!��f?������Mi���x�ל�C���h��+�����u����1��{}�̶���_��5A�����.{D!��lwSv�Z4�}g���.��s�����9ܝ�m����kU>�tΫw�eX�6�'��E�Hj*�ڼ-�cpX۵�Е��K�B�ÙtJ&�+Ʀξ7�'�������w=� ��]����Ý��ے�8�t��V�6�qY��(��#��۽�njI�ɘ�lӭ��Uzj}"꼓N7J����j3jե�.�N��t^��}f%�Ф��5��Ru{$^�!��C6��J�-�m�r������VNGpC9��p�l�j�u�]:}�>��}R��w�.X�wt��>�f����p��[��]�<�OI��j�sZ��H�+�K��؄��KGp���F�󝋙��]m�,��Z�����1�{��)s ��{��IT�J	$��X�۪;3�:�o��Ǽ)eg5E8Zr1%�f���:���θ�h�/_s����Il3r�������2���rH
V^���s��nob%v��ӯ��D�X�S#�V�{q�hn�t.���x�U��w~Z���gt�g^Չ��*Z��|�	_ޙsy�ݮ{��:��gԚ��;U㨡��L�i�'�3g�;nt<��7'�e�`�y�;Q�N��r0�l����J�U]]og%jj�2����C4����֓��E��6V��;E7��؞:\�j������!p��C���#�v��<&�ŭ�lg9�N��O�#=����צ�]tsq��䄬�*���j�&��o������%N鶫�ؘ�;��t�*	�8i͝�^GG�x�(�Ot�+B�
��k@������-��,=�_vSu���<�!X���;y�}ճ��{�e���]}�i�+n+����.q���ޙ����Q�5���X������Ad!+uܩl>!�5��$7�Y��D<,�f��}��kUм�jX�M���.ݔQ�������;[Oo4�����b�w�\��ǘ�73~xt�9�k���>�Z6�pޕ7Bx-�.q=J�,SS�OW!��ޢ]�˗+]΄R7�R:[�-��g-c����Ǯ�����[}e:a���d���F�Td�(�L.ⳝ�9B4�+���R�,;�����̾t�
���ʽ���[�wT�2���l��엶������˖�q�1�b�hq�Ne!Vo@'Sƻ9�0?�w!���Woq��9wcw�R�=*^9ש����!�f�pY��_�i����҃��U�&�-��<�*��	J�����rͶ��G���k�D;1]A6'J��G���Ejo6mj�IS��^�������Ua��3Z�d��;����wm,�	���HwU��H�=�<�{���}�㼕�:�����WB)y�h�֨��-�!��b����)�������hf��T�w����wyG�mn�Q��Hwi�,}�+���ŵ/9����Q��Pn[q>�b*[�;"_����n^��5�)�����[}Ɇ��v���3����-vJ�7(��5{v��	�p�m���B�Kt��w�G���r��{5���7��0���%g1W��4�{u�7Agqv�8D���us6��.����b*��eR��p�=b�p$��j�jS�V3�.��87�̝��⍰#����o�m^��z,gZ<$�)ݮ|��hZ@�YJ�S6��@��^XZ�v�Q3{
}.��V���W�tF��݇JebP��%e�(ڦ��9˺�{��YJ��a�;E�O��VV�:ҝ��B�/e���h��y]t���l�ۏ{����"���.��$�z�S��v�-�"��u�-U�>i,�t9� ��<�-s�E�YG%���%v^�A���k*U��.������73N$��rV���L�3 
���#Ң:^󾡸C�h�m��_"E�Xފ�pf���T3�\��Vi��z��HN˳rU�';��y$;�Y� ._
�z��0U��PLb#���-v��ZR�ǥ��� zW(�Qӂ���L�ox�fJ,�243�ү0f�%�T����sT�}�.�c��;���٩��K�-�b�'���]6i���6٘�w�NlE�b��)�<�ޜ�l�]F蓇�¬�{�P�۵�8V���\]A��Ӯ���m��(�n�����\g|֊c铀����)��w2�J�n^ga�E�a�wpÏ(��. ��;m�}u�]�=I�mI}�S����v֣�]�R����.���b�Ӥ;\x��Nα�*�T�}^wv6^K<op��il���Э��멨���@[�������I�8�`g^�;Z��l9"�5�����r���A`�1ϟ[�1��״v57):g$��}R7H��ڎ=ׅ	�Dg*V�ج���ݑ���르��I?��*\�hƖ=���G�{U��K%�؆f��5���-|�;ʑ]D���$�M�ո�4���:�H��Nq���ŗP=i�yE���}�]���H9R�-"{oXͼ��$*՝E(��f�Z��J�����h��f�y�VQ��=�O�9W���5�JEv��r��T�ʰ
K�VWLʃV3��̥��[$��N��WEPQ�z9G�0�Ӟq4�١YW0����~WN�=*�y�
Ҩ�,�1��=y�JD��f�������k"������4���:f���S��Ը�>�[�6���؝6�;�Y7;,����N��(��"OZ���߯.��:ȹ�{�:�Ky�:�U�k�J�;��ҐޡMO���]�Oױu�1�ع� Y�3ipw���p�=�f�\���k-۬V��t�ޘX��Vv').����[�A
�|���A�G��3ˊ��a��l�#S�#�+�1)�w95S�e�ܾ;R�YsU(�b��e��[a��`�tծ��9J�{t�ӂq�r��rsMe�[[���ޛ]]�m�[f�"�f`�*L�ϒ�ZF�"Q��m3�r<�kQ�Y ]�ghs0a��"D^��������7(�r�٬SH��
���k�mt��Q/bt-�%�h�¶ewgF�� f��k��7/Y ��,F�Z�v��G����-�MIn�¬�ΰ�Xp*t+�F|62�!w���*����R��31!�ͻ����N���."�Ypt�d�[����fZؓ�5���̛miq �:�W�p�
�Xӧ�\MZ�w�ȖKSk%ŗ��=W�-��{o��v�vp��:��gX+H�ٵ�W�K5�F���Y�j�P��4]&:��E�Yy@G�Zw"����)������}�)��Hאָbz������Os/s#���^�J�mp��ǌ<��*���gV��ujRK1r�[}@�T��i�3\�-%�Z�K��a㎏P�ɨ��kWi詥B�չ��u�ʤ�T�F0x��*٭�g�.���+g1L|2&i�*�P���a�#Y��w9�Э�K��@Wu��]�ʭI�d���N��V_	.v���^:�3y���k�T�q�RV"��>ޥP�umG�Zesj�r�[7�CN�^�Y�ٶ�u�5�Ֆ�rf[�!�j	���uE�:L���/$�Ǔ�>�Q�m��j�ߌ�'�f�s�
����T~�U*�J�<
�|���J���VQ&�J���iv����H�6�c��mZ�W �zuQ��R�pߕM=r.$��Kk�c���:��W�:�iY$�vE|�<,�����V-�:^��V��uС�UB������7R�=7��gu2�ue9��=�tJ"b���*�U���dbp�<� ֫�u�����G��)����dx�Gr�=|Ha؂M;ye�7l������9y�;�_T��u�2�/��pIƦoN;O������`���k\U�=o��X�Z�IG�-<]9�Q�M�gv�c��˨��{I���W*g.����y�'*w�8��������N�_b�:�X�4��2�'�����Wf������ӟC�d�8%%�d��z�V�\{�]5w4V��1�7'Um�̫�]�v±
�1�se����ݥKLv'y�^����g��6�gn�_E|B����1#OV3E�ţW��h��_L�#����\���2��y�����rgM�jAs7�JަT��o�Օ���lp��:�IE��2�6!v�����O���*(FGvm���ۣC�P|r�>�7��Q��T�yS�m�V��Y�Eyܫ���7#�\u�f� �9<�\�����0��i��6��u��x��<ⶆ�Ƨ^��r��J�a���\�b�G��t����-=�n6J�7{)�:��s_K��L�3(�ܤ�$ҭ�a�Y������:�-����6I��(����3:��id�fɏ"a����m�-P0EfH�x!�����j�Is�y�����!��*̃]�{ΝZ����S��WM�Ok��M*��y��F+�� �sC���y9��Vt�S�,JY<��I�O9�IֻU��+����.$�t�I?]��ю"�۠���/�����ŋj;��`�49ڵ]�������Y���X�d��]]ֻv�,j=G,�Ȣ��gf��.V�l,r2MiC7$/:��Vi�˫ڒ��mթ�/Gb铬:�z)�6w%�t��"���E�v41��<��(R�~f*\Uj���q-�w�-�01��v�,TbֶK\�w09d�Q�VMwen*���5�Q[=g�3]��R�.rh�}�ZȒ�n^@�����ִb%M	�p�;,�꼙����ax��pe���ǰ�?����)�\,u�� sjS��sblɔc{k9P[#�Ŭ�
�+j݊ �E��`[�ז�$������(���_V���,���{�����܃o�(�lJ�J�36#W]K.��xھ��]�r8�ES&ib��:r�Or�����AH��$�=�qب�Oj<�>�w^�<t�����Ρz�$&m���Xݹ�S"I��X�Q��}ۣ�=��=�#�k8X�ͳ-V*7�[y'P��u������ut�Z>;DK�Nrrd-]���[/����+��E��_^�0qX fc}�]�xk�[:��S�u�\SZ��VX���`s�o�����B�2��?;��c���:n��58o��sT����9�[I����~i4%)�r�d�c���`�]fP�aΔV�O����ȓ�:�Z]����+yWr��5!�kԻ��aؙW}}\�M�T�a\�Ii�\�B�}kj�<��Ԟ�->������_UW�30f�` `����޳:��>Үld�����rPt2˷}]��B�y⼑�\S]�F�.�v���po�g%0s���,^wC�qꃯ�,��u:�0t�4�1�"řIY�֒�-�{��*S����9�5w1���<v;�A����{$�W����KlF(�<Yv��z�mj��kj��	-�"�\CC�{��ѵ͎H���(��1�u̦h��U!ôjhS��"�Z��)�3��U�I�ubq�=W���n������ɏ_�l<Z�Ѫv���ʑ���jdzv�<n���Q�"kb��칯c�G^�u��S׋�PwYQ�θ�9F�
���n�<{e�)ҥ�][G�P�����F�}(	�tT��W�P̫�1Z���uz�m:l�����҆��z���;�."}���՝������ �R`�i-$��.{ع%��;�v8\�y��h-�V氶��t�j��9l>�(�t��t�\W��XaT�_�e��g��+��:���BN2���2t�oZ���%Ԥ�O��E[kY'��9��3�j��K�,���k�5�;v����ҝr��nՉ����v��b�J���3a!'h��S�%�6�g���hj�|e͟w��r�!�]ҫ��u�3��/�NY��2�i��54D�ى��U֠��eqܢ�`�c5�h8ݵR��\$�Ƣ�<��e���n:7�#��Z�� 6����iOr!k3������F���r��������<��
\5B���}��Z ӭG�|9y�ȣǂ�n�54ƌw�r�|��-҂�o!�r��Pw�X�M�4�(M��J������м�wo#���+A�s�cڗ.�,�v��#�ܜk N�C�U�f��j<� ��Z��o�c������n���Mf�:����ׅ���7*��0��T�䜎�Ja�v��*̮�4�jB*�����=ө�A�k��o��p	��#��ݎh�����P��ۘ2��w����99l#1J&����ٝNYw\�"���3�^�a\��>�����jQ���P���q�	%��x]	Es���r�+�u��w�O7�wi3�rO��V�L�F�E"��C��|p�f`���=����a�f�n��U�]�2�V��A��������"�4�c{��68&�sx��;Tɐ�rio^�
��a�Y���`ūUM��4Z�vt�U�L��Y�H��7F�<]�ۇ����b����U�շb��V����g��2W�y���n�
57���o�Uζ�>�V��%˨:�ÕSknkd;�W�w5[�Cg]��bn$3�v�Y;q�!�M����ժ���X�Ow�]@t�䜭]���}}Zc%>NN)NR�i�.�U���+:��^��,���n6�7��f��;c�m�sR�V�D,��ܥ�u=�
�~vWdbS�z�6De�b��5��C�]`�=$J���C�[�vUw0��\�3nn��_%�5�K�j:3��SWΕ_P۫�Xo�vV�V�r���E�XfrW++�d�]���ã��ݯ��(�HoQ�[RZb�_S�]t�ty���,7*l�)V����{9-�]l܎ƬM��ޕ�yV-�6����T�ǊѫS=I&�ќ��0�n��z����kM�2�oEN޵�0�Y��T�ij� �y�=��ܙu�j��s�D݊o�x�D;�����˾��
Z�X5��i����Gc��iY��<C돦1N�<%^<gfP���A:�aý1h�j뮯�t*A�k���<S��%���	X]k��m�&�yf��G)ΐͅ�s{u˝� �f�D[|��f��Ԇ�
��rݾ��#Fh��*"���� �u�PB��n声��t�YY�C�5��'(�6ƽԜ����s�_u���&�����řR�bWf�D{1���N!فq��
w�B���:�I�ŋ�N�����6KU�r�-�^^��U�e\�Od��\�&n���x��b��Z�7Gn��v(�@pU4k˘`Kh�]��c��ؗ�q\*����.�-^Wʿ��%�q<c@Q�8��;!H��2�[Z�������+X�JéU�xǑ���[Ǖj���:�ï���:3f=XХI�B�;���\@)��eጼ��B��tr��	M�wjR*d�Z���t0������ؔ����Ų�Չiu�g�B:���n9H�;��b�dh�G$�S���{@*�	h0��P��\5*ܩ���/�fq2�	u�.�:"һ�00e�Os�X��k�s���̵b�ė� x7Z��k��Z�����d�8�4�au�Sky�9.�3���K��5���}�z[Ыj�Y��e��^e»�����:�}���f8(��$��ŀ�]<��a�4��������!�s�$X8Iڕn"kO���%�w��l�e�:��s&vc�k�޾t��Ӻ ��`�w�u5N���WV��m�*�ʜ���\ �܍:
���U����J�F�y��Xȱ��S�x�1�7v���PB\N2�F����¹1Ӭ��.�;`��Wbna�ҽAؚv��1w'[����ii��R�o@��J9{��x������t-��h�K\�\+�C���+��
_7�7����u��v��b�4�7;7e�y%c-}����r�ܓ�6���W�R4,��)B��Hv�`֮c��8��7ԍ,[�oi����o�ި-�S�|Yi
�٧���f���U�(GMf��N����������3�&U��Fp�𸰫q�U�� ʲr6ؐp���F����Ɖj�f�x:��Y�E�ۆ+�3r�� �(-nn[t�=�l�]�_3H[=���5��)}P��W!�GO&rYQF՝jRh����b
ʍ�o�Ϲ���u`b�(�ܱ��AX]���Y���Ii'Wԣ��y�eY��i��5�SK��b5ul�
dy�u�l�"`L�xof.W��!�E-N�<���ESt�j��U�H2��!������Wm��.uuJ���#�`a�k��
�B�G1����tT�K�!۬C�v�!6w
�70h*�1o�@�o��91�n�"�-i�%"��;�s���wR�,�v�Q��}�Զ�nc�~�@�
�4�9M��z���K�J@�@��|!��6ѠO�P�-����q�lV�k�p�v�T��n�@�\JR����|%( Y�؆)+�FOb�w9ڽf��(jj6½��x��
�*��2�pb��h��n��1/*	c7)f�Kw9�n=��ggM|�M��:�1&��é�Ӡ��E��
 ��D5�l�نɖP���x��H�k'
�kF`��<6+2ә:�o�uhL3�1x�RcV��YZa���ْ�Ȳ���]�c@Lde kE9���eڤ�:)9OJ��4t���
��k/q�-�� �D�*ű��Ink!�)3':֒��}�T����;�{�]�boI*�r>vF�-T{�����[��OBe�ї��DھO%0���Ի�w����Yh���B��}�����RTN�f�7��������元�I��˟[a%��Q�i�
�����&ç�&�FY�Xٶ/��[W�*@�;ĵ
V�秘f�'�Na�����s6�fT}Et�iT�Pmc/j���X0N��t�w]A&����lv9)oM����6�z2���r�|�W�t� �	ko��&���.��<` �8�PŦ�e=��>��._7����\�4�+'�wf���A�Wٕ�u�:P=����X;y�-�Z_X������$�R��@2�ݾZ.K����+$�Ӷ�}��Np=n�5��k;�0D(���n*��۴���A��C/B겱=P�.�X�v�5l��G�ẾQ�GN�pauÙ��Uv�R��=�ė�S�Of
�T�=`�u3��1;h�|�%�E���t�h
�z��-�R��$�9�Ʊ�*K���m�܆$^��ˬT+,9���'8�뫾g�-[�ćs�]ɮ�qR_p˛�s��v=�[]�����vڸz�� 6�9���Kk��û}ӭ��3Nc��rv�s��syw�!�ęh��RjU�q�#4ڶ.�=v�E$B��'��	]�t�1T���"}�q��۹&�M���YJ���29�yWe�δ�[��+:)C��r�빭�=	mp��/;��]Z�����B�:n�ZΥ �W\��*W<VKTr���ub����a�n�*����&��a�lK�]>���\�������a����9�i��WwJ츃���vLX-��P�<deqw],�I<��s��fQt_=b��
Z��%:�����D��#[[�n�G2��&fΕq u�s*V%*+���	�A��d�[R�Z����\˖���a�������Ip�0��uy�9N�wθ�jA��8���D��|]b��Ū��������8&���
wL��*-ݧ���U�@WuvK��Wm�K�N�v��z��L���3r���k�qR�K�"Y[�>+.�x�fJ������2�W�lgM��ha�\��c�u^�V�c����	F���X�����b��ǃ�j�y�y�/�1Ē�/y��-vY	+woU�Df�����vz��N�CT��VM�]bE�Z�VE�9���2�Wf8��m��SN�*��f��fr}��0����Cy@��?��u�G�����&t���ŃlPCo,AZ9H�3�v69�v����]��&�['�z�f��Z��}�Ҕ��q)���o)m�5�X�8��H8*��`����t&���ٮn��|�I�=,�5!�d�wN�,�:}�4�4|+�pyN� =�A�*�WVͫ��oӕ|{e+{��J_$Us�=�M�n�]Fp�S;eu��oAY���w�__3�'��^Zn�D3Ӭёj��g�YG^�G�\�3E̾X���e�u�c��F��|��p,�9I��o1gdp���1�m�n�`8�fr�i�-[;�0�& �bF˕:-̻zD��E���3��ܶRT�kgu�9[qW-�U�d7Mss�	�+�SA��H{0�.-�/E�����$KMĕ|{D�^mj�`Zӏû|�r�����rN]��b�>}dRv�cB�ڵ�}��P��.tl�P����΅�K�뎆Ƥ�h�z�ǍZ=�ӊ�㒛���_/��Q3ZS�M���ƍe+bP���)A+�uʾ���S�u1.��S��{7b�ŷ�޺y�U�mW2ȝ�K��oN�^�{q�BvNI6j(��u�Zf��Ŝ7��� �mf���	<�y���U��a3EJ�b��&��O��}ɶ4^���59\�ՄbG�o;/�M�3�qעg�W�����;v����;�h3Uyj�xrt=m��OA1F�ͳ�6�T&B	� �咆,��4���VWU�{�� &GZT�jԡ�'Yz�f�Eb��
Q����s�h�C�)s�1�q�
�Z�Z8YT��ʊ������y �,9K:R˦1��Y}�J��r�`6��JwM�.�gV�����\��Xi���zC�2��5ms� )��5�F���[���վ.��2��+soE	F�1- b޶b�(v�&�1n�&R�v�	�7���[�/� �@}���,��ɋ�N��x#�{�樟TX��]Tg���X�Gb��Ổ��(���b��X���77��m�]���A�.���$���t�/�.���\x�o	�R�Jq �y`��ڻ��H2��њ�����=�ѷu�-�-k�嗉C�r���k���c��n�[�-��l��IP�9��1�M�	\�rt�g�9�����5�/��D	���}�dPC��De�M�H���7���e�0�j��;�\/LJ��,���̬�3������e]��H��.gl��� WY�mM�V���¥Zn��5�����u*l��I��]����C�i��gu��SA�x'C��«��ߦ5��ut���gs{�n,}(ՔTr��I��̦��]��B����wsّ	Qj���j�ו�~:YK6�)�7��+��2�A(b�����>�t�Y�������������G�kX�xH_6Nhh;'gAI抷�V�f,�Ml�z�6��i�ki1 ��@ի9��y���-��Ժo�L]��EZ�̹3�aDf����}wz��tMmp:�M+�"O�d߀BXK9bҵP�Lr�T���F,� �uv�TF����)�1pD�iޣ���a�ev��*x�:�ӽ�B(�lG�i[���D{v��`��Vw:�mY��7N:����^�^Շ�^�۝�ob��J�'�]ժ��Ĳ�6F_j�ܝ+DW)��Q�֐��0���	R���g�YU6�f���D��Y�5���ݔWf��Z�+z���2(v�םE阭�]ݚdMVK=]8GG��G���_8w��{�s��x��F�g[/4��[��b����]��c
�GE&�ok\ru�`�X��:�2%�;������Ǧ�)����X����QN�@�]3��SGk>���n�Z�	ĸ���J�tc0w,�X��� P�]>kWHpm1����Go(��r�^-ݽXfF�ļ�9�y�T7/�W����#T�jd�˾�Fh�[w֤7�3�l�m�P��[�B���jy7`kٝ�e��@��[�˺5i{��G�	�ݕ���n�Pmd�� L��c}���0:�
��*�]�Eu��ҴWp�+R�:�Gm������o��P*��7��ʏ</�n���Z�{*K��k&Έ!m�r�4�Շ����P:︫mb�)�X-��r���gO�]��p�>U�M<]���UU}_W�}�T����vg]ϰ�ڷ���7%���P�����wP=e�YۻK��pWn� +\ �4e�4��8���C_k������y�.�K��.��Ww�#`dF̟�+4����;N3fR�;iQ���G��>��%{(9v1Χoc�z3�TŊ�U�TAI.��g�KL�vgU���m[	�R�E5Ε
�p�F2�R�k'��x�\��/n�<��|p�I�ُ!��}���1Ib���:u<�{�����kp�n�6i�!އQ������h<1���3��.WI[G�8�.��c{q��Q��]�!H���_ft�K���k�Y�q�[rn�15MеQ�֢Z��X��G�rӫ��+JZ��H��h2�o\[�d�:mJ٤�t��߲v(6����6(60����Sd�
�5�J�4Q�KNZ<�V_A����*t'7���d��&�P� ~LVRy�ѭv�G[�(c]I����V�\��:��rA��5S��&z$�����;\ D�wkT�φ	�BS��x�4�l�8�ǽ��u>�폝rnn��8�u/�$Wg��!�%���tWta�:�a%{z�g\�+3�&Yp��j��R͠�z�(h��|��=ט�7���V��]��](�wx
��rՄ��d��.`,7�� qdr뭩���-x+��Wܷw��Yi8����j�a��U�7��tM*����ʻ�������_�ߟ��E��DQQW.���gK�����;�7 ��������:�ss������Ger7$��\�r���؇u.����Ź�s�ݝ�(ܝ�t��]ηGN�\ܮ�&(��p�Mwv��K�y��+���I\�\�ypW�9��ws��p�\�79��u��ɷK��N�h�w�.��o%xc)(��N�w;�.k�n��\��%�c�H#C��^r��sF����tC0677s��]ܜ�Jaw]�v�y�x�d�7�uΎ���.!��Er�D;��;��4�E�۰�wwy�M^+��8V+�wN�\���\�!HL���H/�m�E�o* ���.<�e�ǰ�˾���,�B>�jrT-�D�J�\�0�M����u]==[���]���Qt�_}�,��N:����L�l��.���y�
�iۨ*UI�u:"%� p��E���AEdR���D����g��x0��.-�+�Se�JTt]��}�ڬU��b��)U�tO�p�Κ�]�Ri�s���#n۱|^��b8,v��}7Le��K��v[��ֵn<�Kff�������0�Ť�vF�pU���
@���5p��䣞�<DӔA����iw�S�5����������^ʨbK�g�����s�F/o*t�Ќ'`��� �ܺs����Y�)�&�/�]Tθ����q�MW٦�=��OZC�C\�Jw�ҳ|a�sJĻe�v��+#a��s�N�1���ܐ��S�-���Ud�x���C��3||�,��0_�So�^����^�V��Ek���ؠZ
.2�dm��g;�W.\�l�f��os��F���Hh�\6b�=@�4�㠓����=*�L�_�sQ���:6��a$����۰���Z_�Ie�ȁ�ڇ�cI�<�+V�D�p��1aW��&�]n���j<����k��H�fއ�s{9K��vX�įgf�G�����CYR+}R��h�s��+����3�C����y��^�����Q��n�C�B���:��fu�o�J�s;�R�J��k��2�ƞ�P�_-�T��J���jH���?8[U��+u�Ӗ8`厗I���)�B��F�ѕ��u��W	��-`\4�-���/��q�"����51zX�n���n�����>y�G�Q�n;*&���0R���cCˎ5	\.�EBMZ��&-���;��T�N-�NL��N�c�^��V֪%�<jP��:�=��9L�:�xJ�����^&u-��ڝ�� _ �أN{C:z_	6{��\�Ҡc�Lࣼ�+vt��U��ѽ�\{���"St�9��{���W�r�"�ܦL�m�ؙ�ʰ���1:8�S<�ja��y�-���ݤ��^Wr�O�Һ��lrw|c7��)�����Rغ�Җ�	�c.76/��fƉ��c��l�e��z�{�j����a��a����'#Ls�]|:��|�m���՝�ַ�kN=�;;ݮw`�J���8*��q֠%Ɗ�l��E�bs`�U��Ʃ��KùW��T��)�u����E۔N���Xh�_:�j�?�]�f|pUL�d_�y׼H�ģCiRα���)Ji�JəK���P�*�
*��v�ɴ��ؔ�ʇM'Ĺ��hu�|hv�K�;��[|�M�N����[�R�=��5+]�	V�˾��r��S����<lç�5V�]�|e7�ᙕ��U�ަ�k�
!w��D�>�X)nߪ��AWS��ȵtω�.�.��+]K~m���h��p���X��7X�c���#�p�W�n�a�/5��+:rN��D�D����T��U�r���s%�:���{۝R�I������`2��7)��/y���	�q�G�YdTo�玗1�K[�Ա{9d�W]��cj�^��&�9;c����9���ͫ��Uk?_��!�#�H�F�Fs�<ާ3}D"Mx��a!ъ��.�/_�}�1|׆y-P�N��1����}��7(��f�Z����cN�@,/8�N��T�2�	��ǵ�;�ܾ8�R ARZ�̶�ge�ӫ��>A��ͺ%�k�ּb$�x�[�eH+muS�7�o<�/��f��Q_�j]x�}�h�g�`6۾���?)�P�ꔍ�0���%i����Xx����u꭬��]�6\�ci>�&�nc�0ɶK�^��_Z��S���вg���B��]ێ3x^�2�����:'��b�Bn�Ju#y���P(E�Rt���x=
7\�ޕD[��w���VU�F���������D��,g�
��Ժ�˚�J�z�&�<��+.Y��k[��R��3'�۷W�_�'_v+j
a��H�
d��ɉI��2�n��ӂ[�tt��X�4���M��u�F�y(o/{hǝ�W֟)����w���|�/�5T���+.�b����juR!2�nX�6>�"(GP�Y
peoA�G:���OR5#�m���i��P���Ƌ�VX���b.1:��]��m���;_����ۤ�V)C��@��,�*�J/qtU�ܾ�u1���V�5+��wܣ��$H��Uwg
�U�0H����t�Fc�R���e磮�K�����އ��cv�-��]v���k��K��Y2"�ވm_��s��S�XO#�-.D�+Q�Kѻ�j֞��������.�m��Y�y�E:L����f�'z�h�t�b:+��;yK�{��{#�-H���mO��AdwU��!	�Ϊu����g���+��ھΡ��J*l�4j�����!�e�
���]�n�c�0�\=��u�ry
��̺�Hң�P���OSu�V$���Cf�v�Ư����<�N��}+z]����	:aj�7��R5:��@6J�� 9yUg��5�U�c��̿:1L�eb�s�����^��<��_G�����բ�W	��9ry�����-�gm&����ag���h�~���op�CSڛ�ս��w:tZ��2�K�5�q֑�Q��RK��Ts���pEnȇ*v�Qŋ%u���J�o�D�=��+79�^>�ș�sZ�`<q�a���"7�;���ѫS ��LĀ?W�����s�2��c�d�=�,G?��L�-��ة�f2	�-s1�*u�ꙑJd���
!@ ۽:%�]i���:n�ri�и�0�_a\)�����	�VY�c%\3_B�1=0�S��J�X񵆔rv	�N��:�����wR�P�Q��T�l�x��u�w��ɽ��@��:"��%�c��>YY}1��ׂ���
�����'f���f���Tw��ܲK�����ܞҘ�����P<������}��r���[ɗ��Ƞ����zwb�D����L�Wu��|�
{�u̙���BFe/�&��Z�TS7�VR��z�{��Ɯ&ϫ�w��K�iZ��\�� ,�V��	*TZ�c(�����hӕ�_+\���S�t~��J(���@U�Yd�WFK�g��	��ki��eJ��/���x3-y����'�r���U�
�|�����`�L뀃'?���q�O�٧�"��8�p6��n}g7ʠ���d�X�#H�;uwN@����w,�Jm�X�ǥ�ص���Y]�3>�u;������*RC��4�#��{e�|Z��I�Wt2�B����sx�'�!�Ԝ�qwN�ͳ�%;�ӣ�r�\Uң��U�������e������:!Qbx��j�J:d1�*����n��m���a������b�Ե�p�K�?�cCn֒t����T�|kL(�����GN��q�vu��œ;���[��	������[|@8M/��$�K��E]���^�tŬ�����}���{�n�$KM��:�؅�ƺn��u1TV�Љ�� �I6Kz��3�W�q{�������&r!ۯ���,p�|��GZ����?c��!o�䣩�?bܰ�br��&�^�j���@Ԅ�_=d+�v�A���W���X�n�������EwN���1�e#���{�?y��"�J,��S�3l֏e�뻣�0wz88��ۑ����x��m���D��]h����[uH�}��R!n+��n;xg���We�-8Wu��^\O�����%�4r1�Oʩ](��#O�m!���X^-p�������M;qyEh�wu�p��"�L�=��#7�0�?E\btqp�����":qL��m2���T���Un®�Ratg^�Op�����uf�m�Z�{4Oz8���nݵ7F�N3D�	����3���%����j�չ��3[\�^0�6��Sƛ���&�*>㲤X�f�z��B̐�����}�_Sb�N7��K�Pe	ۭ�� �ޮ�M���3�/.G'w�5��*ܸn>n����p���[P����uNo1�]����:͍��&l���l1p�>�����~τ��CA�o�$H��;J���8=��Ө�y-�q�[�@�k��]{M����z�����iV��x߼ji���{�]�pt>��_*��38��܀�m#��O.(����.4���u�R�I�&�������D���lS�lyKvjǉ�U�#�yR�w��۪�{�V���	=i�6�e�pM|��/���r��1��W	JZ���M�]�޹���I!ծ�����ų_P����c]0o�]K�o,���Mb�5aS�EZR���<�G�{|��5��˹�k۩�}s&�;c����`3����U?�{�BdpQK�g?T�*ǡ�J�2����$aqߺ�]�Y�ō�ь��p�0`ea�]i�y�y�d�
�Yy�:���CA���9�g��}.���@�Ϯb��vz��M�c����(>W\_
��hR�ך�s�V/P���Ww��H���g=�Q�[\k2�c����};��!���ʴ���a쎟u�RϮ|W
�[��]m���ќ;�l���NQxi���up�F�����N��Yu9��� ���Or��[��ۤ8���k�Br�S\@Ć>	N�`�.J�+�����XӃ���b:�;#�R�\�9���;X�8 �)�P�)�`�L����|��ꜭ������@�/�j]NO|��b��2^UqXĉ\�Mo��K��'���ʍ��2����LX��F�>G����e�1I'fM�s���ȭ��Is4;�Pg3y�J��:��ʾ��D���FS�������B�;�!̶X��Fպy�j�^.ד�h}�s �,��צ�l���H��o�z*s|ߑ�,ZUL@ܔѼ1;N5��n�,���
 l�4���B��a8��<l�WYM�S#iL̗�0Ƞ��Z�m�Yz�gs��#p��|W;�=q�np�;����S��G�E�7"p~nww[�ڞ�N�\�,}P�%Ms,�|�v�d�E�"%
1��%�f�v	ښzx�}�2^��E}~�����+P�N��P�W�O2�ȧI��T����;�b��:w�.I�e�r�S�8��-��&Y�ל� �x�r	]/o`��x?>�m�~���Z��rQ��2�'����l�3�ݸ�bW��#�+�>u��r��q�;e��ζAx)��h�g*ws{8�4�m�59�� �W�n��7_%������hN�{����I���9f�W@t?�趗�Tm*��#�*�
��*B-9L�S�[;dp��U6��Pxb������B ���f~3ԅ�L��A�W�]�X5�я��|��W���80�.ƹ�}q)�r�j_�0�u�5bKa;b�T�����av_����쐟T�wU�w�o�7%�� ��ީi����l��zH@t0�TH�٪�pK��	���//�����E��)�bi�yS������r@�U(�1�$K,T���M�=�}�����/�.+zxj�I�(��u�Ꙑ��h�d�՝�:C�n�W��Bp�N�&K}4.������S���C"�e��)��/cB�c�!*�W�s�\L����sq�Jά󩅸��wR�L��R�c"v'�
��SS�;��Pؘ�dV ��J��:���ʊ�WV�͹�6n3n���-�A��)�L��ʼ�x�OX�U�p���6����GBc6���M���<���W	q|l�\�6�HP��}le�,;�]�� ����-!���*�N���)�u/�K��rw���(��\�[<&�ZOv[\˩4����Q;/��F\��Lբ�6�GR�Kq�Ʉd�(�Е�*��r@]��{|^��]v�V�!}��9�t���J�s��w1%�b�[6!&���@97h1p�ܙ[�HC��eq�)��K#�4��ͷ�-Q��7����7�3y֯낦!���h�!l�
��IR�Zԅ@��\����k������pm�NQ���:Q9q�L֮R�\1.q��n�os�F�moE�6g6WY�V�[jrQq���!qBl�4�,`�&s��7�×9�e��*;��Z��?#�St/6����|R%y-Қ�������TY��nH ��4�5�쏧�L%�Ul��~�<!�>����J�9ʙ>�C�ء�jݲ4#<��{i�{س-d&SӃD0���&b�Z�8��	@8L!���(	�|.k{C!�)�|���]��\�f��Bir�����D1�:����\�� A�c;�s[��1c��)ڏ��n��.l�Q��9�_MC�8`�Z�"�8uDg�UB�fӞ��;���*���<Z�td ��@�o�B�\8gΚ����Ʒ;���>�5j߀�NȂO�&gXJ��x-�*�^*N�6ln�_Jr�7Z\]����oPV����)��R�/{��L+/��4h`.;�U�Be��9��m�Җ����:O#?u��,�S@e�f�Y���JwM�uӧS)!3@�G�:�s���+k�\�PD+i�ۣ�q�ؕ�_P��B�Hn�#(��	���gT�f�y��4��X��/Q
���b=6�k+	���c�-eAS6�3WK[���;b�yJ���E)fU�gmJ��\>ָ*NJ�J^g;襕��MBУ��,��j�tsSN��PU'f�$�].Q[ZҬ��U�9e�/VZ%�����l��O�eN]{S�id[}�-h,���+��V�* {������-b��k6�}|jif\f���_ZA�}|�ǐw<;a�C���]+�g�
��O,�"�p�3.��;�o�`�ţ�Gn��сJ��B��A�f6�zB�=|��nqfD�]H���{vT�E�z��1�)� 6����0�H�bP)�����;�,�zU��(Ss;���e#e��kd�QGV �ܰ�Vq
��pek��>q��E�V�S�`�<�\�r��������.PN�۬B��a�xGeՌw6�e�h`L�����t ����ڬZ�ƭB��R�J�X��Wt���|��NԴ��/�#�;��iu�m��[���Й�<ᮬ���oh<�EA����y���5�iU��"	��0P���*�!��A�Дi�%u�o�I�h�p�թ�C��7ڤ��K�k5좠��d�p�R�[�z]�wϯ�!EB�=4V֙p����Ơ*�z6�]���g aO�I��rԚI�w]N{�pe��w'�A����[���뮍Z�T�*]],��F�@*�eI�X��u��W��W��.��DD�E������>�S�[(�<���1=�%Y|-i��&K��[`{Ӑ4f�9m
eU���R�gZ�ώ�' �\��9^T�����,Sɐ'4L��f�6.˱w��α���H�LW��*� �܀K��\�	��Cb�.���r������'C;m�.���ˆ�{�]]H/������v�Z��JєG*�U�z��D�cBp��b�_:D�W@��r�X4TOz�:�����ST� �8�h�U,���0��]Ԙ��Zco5�eWg[���H�pq�5cV QQ��[z,� �E��V2-�T4�EJ�u���u��C��v��o�-��Ot�wz!�yQ쏰��ʦ~��ؕ/�ǔ�W	�}�bA^Oc�F��:��jØ����w�\t٩ne�>&�j���Cdժt���W���jf�2�$f���[�H)��	�7�|���Q��4���})u��S4�����S�4b�{���y��گ�a�i�BqY��<�y9�A�@�P^%0[h'K�['E�����+�V�ی�bd��)���&$�] �"��w.��dw\d�����'F8�����nx�!I^8Iӻ��.������]�x��8����t���;;�Ic]7�
�\'u��Ηuĝ����!q���r;�]�r،�#ݺ�ػ�n��s�r;�k����r��w.�K��N���:�9���s�	;���M�s�/�.�.\��B
��ƍ�r�������.���.� �;��\��rL��]q����W+������i&�wu�Ѣ�x�&�˞/�u݈��J1�ӎ�sw��!݌�^-�yܱ���듸�&Jg: ˻���.�t)���\��qΔ����u�\+�����7D;�fRf������T��s�u˻�fwwyו㎻��Α\��i�$
.�5�F(f�١�qmn�Gr��+�x� ��C�W��{Wo�|��ċ�8gk*ˮ�����V֨����T7m�([��>�la]���wL�S��+��R�P?V
�h/_{^"�}W�z���cs}|Qx�m��h�}�u���^����}��/��>u�����F��DG".�}�>c��
��w�ջ������8}�}�3����8m������v���n�ߟz�ϫ�hޗ4�׌o���x5��ǻο[z�sz�|��k�����ߛ�W��5b�����+� �
����z[�K�4�j�Y���~���@�����}�o>��{o���o�}����ssn��|�ʋ�˛�=|�\�+��U��ƍ?s���o����u�ס��*"K�,Dh����u�S!+�Q��m�'s���#�}"#DE�����"��E��7�ϟ}o�~-�5���U�o�^�Ϟz�����M�~}���W���_ϯ��<������ߟݽ�����7���-NY��"C�,�@B��=�����j��p����"�Y�F?&k,� �\�l-��m )Mo�̋q��	�[�������������^-�߾�lE}^+��_�|������?W�߾W����r�P���3< �@r������7�jޝ)w1�����㦨
b�
���_�}��mʿ�����o���6����������_����z[����>L�"�,ʇt�7��d0%���Аl.X���3��XC-B��R�����ث�T�ZK2�#�IXAC~/�}�x�W�x�U��y�zZ�]�?�����^��W�o��W�k,��Y���@E�fSY���E0]���Y�}��}�	DM_Wz�nr_��$�r���A�AfDo��^}�~���^ƣ{�������Kw�[����|W��U��痥�|W��{���|W�������o�o{�^W��o��x�Y�|\�5���=Ͽ���g#���/A��W�UU���}`q�|^-����7-?��������oJ�WK����[�6�?���_����m��׋}o-���w�^7ſ7��M��� |��#�(}���B��c�I��]���������߃b+������5z���q+�g!�6w;Am�f �[+�F�_[wο<��+ŧ�������so������6��[w���ߪ���H�L�Ci ����`�u�1.�3�]]�=�ï7+s��۲L�P ���ݪ��S���9V�t����4�[�Xn����'���8���i[�sv�k���X�m�3)VV¥�����"��}�����m�cL�C�z��Б�V��7z�T	Á�W-�u�y����5�����%����������zx����ﭽ�����}W��ۼ�_��^�ּ_V�/�߾j��ּ_�������o�Ϟn��W�^���W,x�6�5g�=��^yt>D�f�����E��W�b�.����W�:���[��߿[o�{�}�W�����Ϟ�������r���ߍ����|���m�_��ן�}��Y鞟+�
���>��#�<LF�[�^�����x���{�v���湯[���6�o�޼��ޟ/+i�$00�Y�ut-����t�3x�-e���;a|�����FFz��=j��1>�g-%�j#�d88�Y��<{���_��~-������5��[�u_������ln^�;���߭�^+�����y����<�{Z2|_z��",G�,��۬=�n������\���6�[2,<:��#6�-�|�ץ�����/>W��V�-����{^׿�k��|W�v�>/J���^76��|x�}m�E{�:���n��#�#��"<#�u���{б�Mg���շ�#����k� ���{�߾�����;y��叫�o>��_��w�}��ϭ��W7/��k���r�/���o|�\�����ү���Τ} |G�/?l��t�����;�w^�3^�߫ƾ5�_o]�����W�n�w�~��M���⟿�W/��W�������[Ҽj����K+���_|���}W������5�W��{���/���-�p�#}BG�p�W�Ρ�߆}r<U��t]�u���r����M�$��d@�f�ȴddS��l,�uٽ-�^-������Z�����x׶��Z=�������}�x���#�|�~�@���E�_��Oe=7��¹��U�,�g0Y��"��Lϩ��/�-�^����[�^-=����m�o�no����/k�o׍�~��-�\�3vK�!�!���o��H�A�-�]�ft��P���]����my�s�EDP��ۻ����~�y�͹h�|�}�u{oM�ί�oM�x׋��{���-��i�_��W�E��u�oO�_�x������>��߿�_���o���_���~6�}�G�S��{���ٲZ3�[�����q���_��i
[׺��-:R�'m=��j��8��B�>P˝{���V����vdOq�au��5ڣS�U;��rޥ���}�n-a��+�}�Xb��{��t%�`����C�[Np��3��@N�<�sɛ�_v�w5��������Ǟ���Ͼ\��r��{��+�F�ە���k�{k�\5���[�x�W��u���Z��W��~o:�W���o���������g�s� >�G�"
�^�.�{۾Z�b͵�á����Tif� �ab!�__��-���|����q�����}�o�{Zy���_��~��~u��M�noƽ��^�����7����^-�+��ǄEi������yUj�l+�w~��Q�c������^5}�ߞ��_�x�W��y��^��W����W��{o���׭�V�������yh�ｷ��~_~�_���������+�_����m�����LDxE���$}��{��м�<�������������s���ץ�j-��<6��`����f����@���Y�V�������n{�|����z�o��ο���*��ּ_����.Z7�~���~�"��@睑W=s���Jz,��������}���x�<k�^7ۻg�W,}_��ץ_7�^��=v�m��U�K��}�j7��ߛ⽮m��η��|�M�*�~]����F�͹�k�����>�鏨G�G�H�C�{��XG;S/�מ2���P`�Y�N���Ţ������{oM�^5�~v��r߯W��O�o���痧�oj�.oKƼ_���5�^��ڹ_V��m����
!���`y[,�3x�-�����\eק��Q��j]���A�}����ކ�/kx���W�Ͼ~E��������+��Z��5�������7�^/���w��؈���x������[��t�eK�!�-L�S3p{O����i�{�g`X�n�z>�B>� �=?o_�o�x��ί<��o�5����ڮ\���x����6���s��}����E��N���^|�_76��_���׮���ۻ��<c}m��=_~|����o�^UoVo�^bC? ��l��l_�}���վ/ţ{_�篾���W�U��z��7չ����_~���ήX�_�|�گK��~�y^�;|m����ν2t� LL	�E��k�^��\׷����o�Gp��g,�2!�hI��ѣr���[�/����<�����W���ޭ���s+����[�_U�x��o�~����+���*�5�W5���Ϫ�����_�z�����W�ޯ����g���t�X]ϋ+���k��E�|��#O���?x��G
ηq?v�틦�Y�3[g%��4��;:�aK'�z��ٓ�輻��RzA�ٕ�y��G��"]]G (Ի2�+��N���e�zX��V`��곳7obލC˭f�Ìr��C�ռ&�l�O��_W���x�m�}���^���}���oʿ=u�����zom������s~?��ޖ����|����Qo�~����_�}W|�\���>���׍�x��w�k����>�q�!8V�2�-V=Ƭ��ִ���{_�i뷿�^7��z[����h��{_�u����W�G��2�--T���ifrKAjm��_/���|��xۖ��}��6��D�8�}��.`x���yI�r����������m��oM�wm���{��Z7��w^�ί�lop�W�kžy��~���Z���Z���տ��ѽ����׵���x���<ס���ֽ/�����+��Z��)��kȢ�4��s���_�����ﭽ�v��ſ/��}W76�ʽ�~��o��Ϳ^}���<�齶����F���߽�-�x�k�^������^/~u�[��Z��_����"8Dp�|%����ǿuϗ7S���}�_��~��^��_}Z�5��o{�����k@f>�o��0p����pHb3��mؾ>ٜ�G	�r�(���Ύ�ԧ7v�E��8�Z3�W�4�ok��T��	8�eo;�*�ڌ�P�X6fmb���V(]bZ䭡�Lc�:bN'$��%�Nv����]+�#%�3��Xެ�C�KW�����y�8kS��� ߊ�
�z�xo����c3�������ceٗ��;��E��-_L[��p^\>)�-�	�I�6W�q�Ot��G_�1�W���o7&=���r��§/8<&|�o�]1���Z�N�s���bcl�p�
�Gi�m��-�=����
��u �!R�c�/ӂZ��U:w��T�Wت��N'y���k��׺s�9�{��%�ݮv�JR��4��+�vF�9˔��SӍ�(<z���4`ǔ���]ջcef��2�M��WCK��8�ٳS����r�J������S�j]�P8}'m�ȁΞ�!���ۄ�\�LqY\�\$�W|����+�!|��:n�ܛ�RO���5�Bj>\���jK/�h�3�u��e�8
=����S7�j��֔���@cg��u��UReӟ��4XG-v�֤��8�ٕ�))BxPI^�jSx9�E�J���9]��L�Y�B�Wo�%y���U�0�es�d�68�t�����k�ɗ��/����qwB���td)hB�T]Һm �]�C�+0د-��e^
����R&/�c%�8�w_,�T�F��l�2���{���'�r�κ����?Pp�EF�'Pɯ�u��f��`b�@��(��	�;?f�v8u��孾�q�����h4v��t�)<��TE}jS&M�n���P��$�L#өB�6]qv�R|�el_P��b¨�X~�{LWAд�к��gܝ��~d��.����1X ���p�j��h�>�@m3[�]A��C��	���&�	S쌍N�F;OK����Y�s&o���;{C�+���P�G�IăG�sP��y��;7�8��+�������H{豸α�OG�U���C6�(G�\z����#4��#�J�����ں�d�t�gl5�l�Uy�YN���U�����ˠ��C�X��}��"��ٺ���Y�e�j���J��b��هj�ET�� T^��.뇛$B��Y��i��$'n��YƝg�	�gj�DՆ�o���	�҅��Q�６\b莱i^T��h���Q��zȹn��r����Ob�dZ�?��0e�]��V��RwX���'��<�hwм5Q��P�8"ZS̾ط0����kUvt�{$��]�Vz�����:Y���m)&.:�	1Q]|�k���/�7)��M��q�uaZ�/��ZYC�u#�W�z���	�۶��j�O��>����r{�m,N�Yv{w����*9��E�i2t��IaZL�Y��.;wQ.�Z�-T��u�M�5YO�{���q]f5'ۘ�p�v�u�5�2q��݋JY,嵥�
�ÄW���`LSz�'dqR�.u��q{N�<4��`��T��J�� G�>��h/謚�M�U;�U]x�K(�#��L���$�#�gD6q��m��-�+�'���q�3W��Q�t]�c�(�of�Q�0�J��0�8U���֯�z���&��g���Im`�Qsk�j��Y}+����V��fhu��
?�:G�uo9�4�\[X̛��bP�WG��1V6��1{�r�,�U�=�{L�[@@r7ܺ������ے)ts9��>0��.:(���2ѱ�mG�u�6��.�2^#Z|�� "lN���t0����P*f-_�kD��$U�;Lw��:!�|U�U��fˮ��g�RK+=6&/j�����{2$sc�'K�%�i���Br�T��F�!���B�;�KQ:Ù�>�G���i[!]�P���h}�����~&`W](�~u~���¼��o�(]Û�~�[��iD�CxX�L�+W�Ǌ9Uܩ�M!X!7�؜l�S�ѩ��p�u٬�t��ɚ�ɨ�A��L�m���&C�n�!��G;�=o/E|�`���`�%Y�W2����_[�M5p/U/%��}��.��g�ץ_Z�Y;F1�mW��η�������л}12��ټ��I��'��(1�K�:������J��ò�V6��H�,N�<���o��v�f���y֧��<�Va����!��V�B�e���A�CS�g?�uS>=�ԟ^r''/7��ݑ�꬙���}_�M���+�*>M)
xWs��E��j?Q�}���.����y��=�V�j�M��~X_�o�X�ݝr�t绬���!�z�<��;+� �2�rT(m�iP[ɫ��{\{���b���;ÙDgw[��fp�C:��r��k$IÅ�\C�M��/w��K2�Y���H��D�	���yq|�m�zg�|ؘc.�n�����epT:��%�v�6!>��{*�Q��ʞ�fN-]�}E�+��P�Sß5%��� ��Cީ�Wρ�UD) oM}%Tˮ������=4�7ݽ��1���|������f�8ܑP���u���{/�_yt�����Ro�0�Y zz?��{�
�k�}���N�1�斋&,kn�v%T��vy�޽𞳲�����*:�T�}4.�������i.�Ϝ�e��ž�a��{�b�M���s����&��)��#���=-�zs#�4�0[��.z0�4ݾ�w����gIH����.�)C���g�������=��w��{~x�0r������{V)���ቪ�7X���`iy�
���.���C��*�G���T�gO8��l�.���c�ۨV��ӑ��M�Px��-��ޤ8�$.qX�Z��+���6'�_s�o�]K}	�#zS7�u���
�xb�qZ��wpU�Fiڄ��{��y�M8�#�}'Ya��ݓ4۴H�}{kjoI厞����8o�M���3�Vi��[\�hݰY���@����Q�o+H{o�*�����þp�;k�p�~�9f,'{.�v�-u6�鸩gA��B��m'Spc���յΕu��G1�4W[8{z}��B�/+[A�^ă��&0BNqS�~�<Y9�(�k!��t���\�=VMO�VL���nf�hZ��f��Zw��ʮ
�z�xB��X@wb�s<6�����'g�T��ϝ�Ë����1V{>L�y��.'�U�@f�x[��;��ř�,4,>��{��Yس9��$T=�n{b�1
�y��1v�κcCn֒t�Fx�����av�<�a��&�m6�Usp�����,�v��Y9�ӃD0���&`�,oD��9|
&����rv�#���e�b���ut@������/𿥪<xpA.T����,�9D1���.q��{����C��J����rA��I(	����=���]Rg��j��,t���p꠼���[!��k~������Ġ�J9���-$Ϧ�!-y�v|ވE����߶7��H8n�������Ҍx	d@�&�y�P����w��j�{�7y���u�_j̸�om ��&1��M��$ut��Ar6�n��~�c��qQ�)�{t];M_;�,�{څ�W2k�i�i�7*�)d���P��R)ѕ��3\����u����3;�smW^5])���,lr��ؗn`�3Wvk��U�sf
!Fv)2��j�<��m��}��,�ȩ9��]EW��9m��Ɲn�7�����*!Q��-��Zf���1�J�@��6�~�BfF@����b���͌KN���Z*��n;���֚�*ԦL�܁�C-����H�Z�������lΛ�)�QwjW���.����k��K���
5�̚�.�͊���l�t�vג�ǖ��>�1�G�mצкC�בC&�2ki;�����Wvz*yQ̭�W&�vR�soi������b��Wê"y������ޕ@�k���O
�8��kpz����}qk�v�W�-Xy{|���Ll9[��x�wQx��F�T}��n����zK���oF�ws���D�0���sΡ�p���{�=�	Y�Hx�/�5�	J���,��!x����]�nE8�T���CF�ˀ�0�ߒ�e��n�aY|c6����b:"��a��X�.��۝9',�$׉�Ψ%�o既��|�4�|���k���/�)�����j�i�n��$�]x����c�[< ����u��/���(��ן)ة�����}~�˄��[K����7�>��cYL0J)���m�g�]M$�=����>q�ܱos��%VJ�\/ha�(�	��զ��=Cl�"���h��W]�r˙)|#�l�{1��k{O�医P�]M�{+Y7��y5�]�Q�uӄ+�S����.R;Zк,��E�d����f�|�Eh�S����N�`�k�Yve�I^)"�V��s���h"DL���p�ݎ;G;Anl�4�����F�kG���N.�ZA��Ryҹ�/5�g\�*]s�;v(^}�&��t�JA�M����&�C;��U�������Ω��׉����D�w�/m[}���7��
,�6enk���u�(�)�rp\�Sh]�Fغ�\�fג�\X_Sx<����ݟ	�륏&TIm5:��C�Cc�;rX=Z�[�y��mG��>���m"٨6v�:P�65w%�"v_n��1���ӥd: T�%�N�uc�Nn�J��VN�wwˣt�_Xx���s��k�,\a����Wv�QCY��*R�66�;�X��;��j&�:���l5�t*�c!4\t�L^�V!P��1�%v�;z*��Mgu�Ԣ����ٴјf�(6�S����_�Ɠ�U|^Υ�ΰ���)+��.��O=�d.��w��>�#���V�.���k^��l�� 0ۼ���O�o:@�u��n�*-�Tw�>����+sU�i��<C�
�;�����,�>�S{�x�,���\��WB��y���s�M���w���� ��b7�7�60�/JZ!�яp��Xv�S5��Y�"��Z�y]q���J�Q�����iz��}a�,�\�c�]�y�s����}�.&G�X|j���]&�k�e
�7g���9z�1�0&4u�[7v��8�P���񅺾���.]\Me���m�;)wLn��b����p�c	JKƚ�5:-4�����)FA�V��+9����N��["M��*ʮ���C8��x�G��|�l�w��@(6�lS���;ޱ�о��A�r*�b��x+x�R����nP����
��u�ʚ��1E�2Ř��<�E�#}q��2ͷ��"��䫪iǐaLU�g 9�\3��f*y�;0��_d��bm��+y$^� 6�r7�7�Q��E�K���U���ֱ��9�{z
�I����<����s����u�d�n)��P�ڊm�{H̺�]%]�,��S��`�--5*���N��맵�q�<�5vw��s��C�-�v\�Q,9Y���M@Z ��$�*P��Å��n�v�R`-RA�Oz�ֱ;!<�()�{v0�0�S�N�nI\&�M�#]���OD����4�bYlcC�2�!R�X�Gk���i�;�%�GpN�Z<�׊}�Γ<Q�ؖfm:x|6e#r�V�|fȫ�zv>DV2-`wHR�֋�۔��0�'_�ᮧ���2$��:���C��� �<�������"���"�9�wD�Di���ܻ �i9�+�;�ӝ�����$�(9u���p�:.�2�:�`���4BD�wp��Gp��y�v�#�s�..u�܈s�y�� ��Ss�;�!"���w\N��u#.]2��k����H��ݕ�̝�$����9�Wt븻�Q#��^�	��xI��]۳(�ь��wQ"`�BSή��B�Ĺ�uus�q�y�vJ4���]�2��v��n�%�s�M9؎tS��wA���1��@�B�!"�	�BN�E�sK�7"��s�n;]���������w(F���.�www�ۜcfG3�tD.\ƥ�̻����4�&H��"��r�R�y���wd������;�!$��wv���Jaa�F�y�B�&�
�B�T4'p�1c��d͝�����m]�˪�&�j!�Fm�j��<�WKG+M:��|�{��=����֍7�=�J�6����":k'�g뫁F�0�����iѪ�Y '�]��H�5�r��W��>�/{-�/��R�g�^b����3�Nf8:����ӮA�('�݋H����$.d���9:vI��ʗ��δ?����ʆ�&����	D�9� ��}Ys����o����F9�_�T1*�+����NR,��p�k�m�npA�2J!�.7�%.��n9�u�T�`�xEĕ�f�L��6�K�ɿ���_�g/>F�%Q�X!Z��G^v���$8�(љ���X*%�1"���b��i\䆋�Rb�N̝90�PU�Ky�����B��[頋��Q{
&4b�_���5��\����\7�p�U�
���h=��۝;}�H��v�}��	O,=�4��c���X[��.s�\��~�pHV�Smvf\�=��y��ʑc�����T�^'A����߽t��MX��<LT��b����9,�\�%�z���$ƈ��vy�;�0��*b<�`�~�����]>]=r}��Fnz�rш��R����j��Bеc��_o'X[�v�����֮W�+q�h`�R]iHg��Q 7��{�������Pس��GHp[bj�[6w�\�QR{V����Xh4�,����]*�+������E_ʯ��������秺:���u�ZD�d��f#��C�S\�&D[:�W���[Ń��mL�z֎"κ�*7�A�'\�	6%Τ�(�=�A[�:-�m��ˁ�˼yQ.�\I���/[��l\��z�@��
�0��Y�˿
ʦ�=Z�3��c�4�BW�������բB�H�S�d���*Q�4j��x���m)�ǅv��I�s�˵Kr�P���8��a�����[�K>�a�)j�Չ-���`{��D��.1B�W�)�4e����'��{g�R��Ƥ�=����R6����d�� �f�.��+�Ɲ�HqZ1b(C��;*�㐭���2�q�S0�iϡ�":�x�F:�F��7f2�'*�%}!(�CPC.�d?��@�xG\z�p�.�0�\[���r��ܓ(Y���wv����TM�������H����H�DžU�P��٩u��!MBḣ�6�e�:�պ꺨��k��V�O(`�c`<O��X��pz�g�'C�Wr���u ���tw!Xf�B�H!t!��o���w�*�s�J��__s��fVa�Y��G�m��*;ՠ*5��汱Y<�n�������^��k���'��fg��yp�v�w���[:�Z
���W
����}"����wg2��G�
�>��ﾈٵͺ�[���C�I��ɪd�fX�!D�ހ�q�R�9�R��-Ǔ�5qg�%cUR�����lp�p��K�[	��+�, �D7,/�e��O�-,�)�ְ0�ۚwT���I�����p��T�e
ջ͇�M�Yb�
�]͍ie���%��L	l��;��+��c�ۿ+|25�N�[x�|�����V��9��Ch�,���S=��k���K��$�\y!4��z���,���^���D�WD�1Έ�Gcy6������3vm�걽ʵU�,���u��W��nEr����tH	��O�vk���z��^�$��RY��t�Y�:�4���p�ɞ=Y)_�~�$�<Uw}����]�����eX� uPB,crED-�n{b�1
��8���r��̽��@��{x�=���Ly��\�瘳��|�d.�J��o]�dt���ˇ�	��j�숕��`8L[C���*o�I��Q�	(���B�Q�7�`�P�&�+|Z%�

�:b���w��6ȸ�iO��)��Ay��U��V�����̮�~k˱�x�����T r�����c���8����� �'�r�ԫR�l9��[�{࿍��d?\�����/%I�[���!�%�%l�/��s�+�ۄnRCo�.%?�">���I]���`�;��Y��#�`��뎺��|���_C�8`��Z�#w�mZn��R�]��l�?eD*�b����D���<���C�g�̅p�]�p@�N�g����<��9�♁���!:��!b�V�u>"�V�Yϐ��<�oy��Jcl�Z\�Et�<��{���.�1l�M6�@��;����~�(��	KR���1���{���3Cب�;�k��c�\�F�*�KnxĠ�W�s|��/�b�NΏK����Sl,�� �˟��V
9Gb;�qI�}�&��S&O|۠9�C5CrF���ߞ��p��,��a#���å{�.���v��oy�53�����h��v���rOk�*�^�׌������@m�u�����zk�Ө�:<>w�5>�K���f�!���w!��Vy|5T��8�L�To�P��Eu�(�Wo�k�Vo�I�|�V-3`��e̓�S�1��hoY�_(�����2��B��|�}S��E�e���]�'kG:d�u`6d��V$U�P�թ0֓r��L�b����v��i�a�y[������A�K�Q���iݜw�Z�t�sgP�+ō;Z]Y��9n�Ӄ{yF�N3Cؕ��֫�S�Vd�����j�G��"#��˼�ĵ���Q����v0�غȹ�P�8X�}7󂧱A2-F�>&�������KԸ��r�Ls�UH����\�&��e�����|c6ڸA֦�X,�A������d��t>$�D���_Lu)cV��X�Ls�����hģr�1��Y.��,����1񂏋z�:�P>���oϗY��]����V�9f׼^j`qڄ��삫Y��X�'�t��eBF�]t;7r��{Q�i�:�t_R\�6:ףoS%�4{�y�4���/}uF�;w>%�F��a@�)V�c�eG'��+�BWF��k����t�8\)�|wa�C���mC�BiL�5@��(P'�ܷ�:�>l|�˫��+����BN�9����;X�۾���$-�߇`M�
�˞(��*<2W<�@�j� :�Tj�>�p7���K�ɶ�8C�d����K(���I�팻��z*	淝H�K�jL�8鱑��QX�1�V�s���Y�') =i��X�1�'O�?eM�.S���u�6���ז���rc�lo�~�V��E�8��|�JK�5;n��C"[�o��QI��X�(�&�n����v�%�HWQq�d��/�x0�ji��΁���3.���x���.������W�UW�~^���u}��̟%1��j2*6^&��u|%����4���T��
��L��én0�� ��Wݘ�w���v�T�!��w?�g=��r�ߒ�cN7$�Myf��󁫧X�����t����ڶ4\F��S,GF'A���;-���u]H��:���E��h�l�����Z�\��{c]:�D��3���mu0�	JX����u�����p�`�W%ل���y!uM�s��.�^�s%R�,z=-h��KV+p��$<�5̲v�c=6��͌|#&=��˻��u�U�1(Q��uJ�	6%�V0Ҡ�r�Xچ"�)�X8;��j��>�(�C=�
��S�nB�*GEp��+O���?��{(jc��p���R>�OeV�<�{3� �p��	�Ψ�\�1�b�]�(Ѐ#p�����!�1�R���^Ӿ�؍��s�֮�,���|&����������eG���	<��w'|���5�I]�������y��fL���tj����9Ԗcn!����z�m�w��MK��+8Y��j-�
��
��\Q��Z�ټ�1���~tO�`���I�c�՝�n��%��]�:0\%\�qrfa�}�O�.�w+�Y�����d厨U�o�=�ֻ�nU@rH�cl�"����:�<�z�&����Oj�e�N����FTu��N�kG�-��DG�D��ɹ��4 W>�<3PU��1��c����];���%^N7$G<u"�b1PGF��B�4�?� E*�#Liʇs�:�`���_9�E���������l�y�p鑪b���-�7�$��h���E�=�x^�B�:�j��K8�tw��J���x*�hjR��1����'�J�8W#���
a�H��.�t4�^����b��yK+o-��"���z�Ԓ�Kϙ�<�"0	N���(��d-7�GH蚻�a�m��{�3x^겨���p�T.ylbj�M�`)�`ix���/�~��OF�5X[U�JZ�6��*�p���c���:ϡ�=S�hw��$�V�S����A��on�(Ź�]�h&h�=��qy���|kE@�6�K�d��n�ˎ�\Oޔ��Z�����/�c��=�K��tԜ޻��锡�!%J�Z��i�4�va�@/�����&�r���ڷ/us��%��Fe���͕[�i����녊��
�O��ܻ�<�:�� �OV��E��)�brZ����K���+HhS�]�Yr��9�������������d�=6Mh(�>�-� 5oo(]�{:�sS{�"U!�K�;���+pm=1
6�]�'ZN�����`�j���\���.=`�~�����Z�M��\�(`�v�.[O>.7��t5Z��o)�K3S��J�܉�/j���)W�z���>A����0�:�1�nH�[<��źb���|��v��Ig�duڮ��i�Od�·QV��:�-j��ّ�s���!����3�1�+o��3p*��K��;/y�7��"M{�N�����P�Q�.#�`�H�BW*zz!�,�*�����Խΰ�������(Kx-z���QZ�B'	:L|(�v��L�_M9c��\3�
#I���l��#�բ�jN�������V.J.�62���I���2�\+��`W[�M^��unZсæ��g4����S�Z������v{H;�FB�(V��������2넞�U�u��	5H(r��`d�n�x�&�c��/V:�ěQ�*k�3tKQ���ζ��l�wW�t.B�yL2y�\�f��`d*�
�1	Hv\�LX��[�J4R�v��q4��bT�p�������"�L�=۠9�tAyUHnlt����[S���Wu�vn��׷��hoDT;����%Wc3�6���&
�s�t]٩.����N�ʠ��Y����q�M˾���a�\��"���)m �:��Ґ�Zm�y�>�vt!�RNޘ��Q�䆤������>��U����z�t]�}a%W�C�����Ϛ�~x�o��MB�˅���m9�c��}��}��9�V�D����/{���C�nZh��]�9�0*�|��s/���/�N��ckފk�QĚ�6p1%�#����W��"�hɖ٨zR-jWe7@�0�� iɒ�@.`���m�U��C����*��1p��m*|�9��V�?�c���^'vʮ�	}��mE�'�6ծu�u��s(̴Od	� ��Y<�'���U�.9�p���d´�k-Ք��V橚vg	C\L�3��R7sѿ�ˀ�5	O2�b��¸/�f�|'�k�qW�e�T�����I�w�I��%�_	�
�e���Z�&*��\t��0xd�eoK��v��on��]���ݯ�p�-Q��A��\
�LPnݿ>Yة�&f�❋��1މH|�Lc0�m\<�[�#Mj��C'�\�Č.q���z�=����s}x�=���'�=�����KFϤ��s�;w,�vձ]@�ݑ�o�]7�r�.NY��[|<�v����8v'˺�5ӎ����`�\Ю.����+:q��9Sk2�	|�鍜���St�.�Af���,o���˒��ہm퐫L��tf��|K���2X|�n\npySyO���F�,n@r�x��U�U}_�[�-���٨��y��}¢����Ӹ�p�)�݆�&���N�	�2T�X���o�u�+o4�@0�!�-փ���"�'��'I�s:!��v�m� !.ov��"��)Y۱�Tc!���@�w��ړ5i���xPԺ����8C���Ǘ;�'��-i`�d頋�8�$eu�:YJ���xSH��a���Zn:!��2�$�h����D�x�ԛ��8�gz���z���U��ڇ���=�LH�{
n"���ɍ�]s��6uk[-�������\�s4ܰ	�s��yRl�z�L.�;��ysuN�>��cmQ+�!v}�hh�5e�J���N�3e�vn��HU�'w��������Q�p���W?�]��WPT�/�]Lz� #К�*b9��\G�npw���+�\��7�<�"z��i̯�\�D��P��j�n�Wd��}x�\��<���t!�6��z��+Fh���[��U��|K.U�	D������C�r�_�<�
����j��,t�<�o������QvMV�^v����Mobc��*�p؟[�:��vթ΅vF�q1J�/��Sn�N�w:W҄��qYW�Vn��C���1V�+�*&���䘩؇����w�np��b��,��gmp��N���,�u�n�].����y� ��-�&ټC�k8jdbu�%P�|��N�]�����a��`�RâX�7H�*ڭ0L��������NFE-4�޹KB����g)��-�S`ؚ*�xrX�WO��MT�8 ڐ�\�WV�ܲ�Zu�)�����2՗@�sd#_eM㖵���"�3"�R�q.�N��1ٗ�;��nx� �̓�-f��s]��_Z�"����i�t��5�ZO]]��; *�y��L�B
�9�#;he�9R�.wd.K�{v��1=��T�H;� oe2�J�ԥ+Gxj�1�ze{l-°gܹwv�ϤP;�{��}��-ɖ]:�+���r>9�#���#����1wu�,>y���:���j�V�]:l�7Om6�%�%i��{8+�����݌n
��������a�"�v�@�l�a��*o�w_Y�����K�`�Z��J����<���Z�:�t��r�]�v�gc����CrwE\8���g����Œ�9N�얒v�=Y��K&���t
���Oiq3����N(�aD�?6䂹Ȕ��ʫ��ϊ'ʼ�g:���T�:��gP7 $��M�$5�i
t>5F�ݣ�wWS�!�GY �+�!��X��m�"ҍL��w���K��9)K���T(��T���Kcg*%�ԭ��uͳM��@�*_^�F��(c��}��Ŷ�1QL@]Т��2K�U�~KPW��s��v�۳�X�� �ƫ��W��G%Yi��[%j�ҩ�<�G�{���r�W�n]k�|d0��L7[Q���n��հ��RH�qp�i=��_�}K���NQ�`�2�tZ
j�L�>��Z�0
 ��qP0e;�z]f��MQv��we�J�m�����5K��`��N����s����Jdu�ϑӖ˱�W̒���Y�\��	��Qv�,���m�G$�����c�=غ���Kq����u7ۛLG�봇M�v����������<�t4J�W÷������E��om4�↸����ؠBs��|m_uI�V�P�͓�eѻ+�I�����J���e���*["�'8KHL̳r=M9�5�^.�[�v(�Z�)��}�K��;H��	7V�1����l���	�t�.��9�K�q�Y�z��HѠ�*�=Z�9+������r��6�|�b��M�&	���C�]�����ē��4.w�m���w"�#j�)���u��,6i3Y6խO�Y*�eiV�����#-��|��l�3{x��h��Jͺ�c�9�Q�׃In��<aP!��c�D���������=�{�L�}�$�
��Ѥ\�;�ȉ��یf!
I���Eˁ2�}tx�r�y"Z$�7I2y�s��bM#�H�w���y���HOwh���D���ή�:Q2��]���/r�3y�i.���y�Ԉ��<�ǎ^w �IIDR��
�W]�y���x�.d�*$H<v�(�W����$��1�nJE,�C	�#.n񹧋�w�qd�˜�×M"�y���9�Gu��" �wvwv"bs���FX�):\ĀIs���wn��t�v�����QD@	"��EA�H���$ �']�!��L�����"$�#bD��� y�I#��gw9M�H���BwnJ�S��Y��pL��	�$�*b�ۥ��������?��������=1h��% ��m�yI�-�ڱc�M���n���*�|�j��M�0AU����Tp7�. ��>���\���y��r(ԩ��*xFm�w�ŋTU�#�̀�L�OkK��P��:�
���#:{����fj�m|��t�_��g��u��3�)vT�q`ك�f`�RSc�J��i��-6��sz��48C���؅�[���p��{#�[�H}�ô:��[�T�H�;n���'/;U�P�d|�ź2�}uQ(�
[?T)T��5%�ۇ�C�p��F�w;{�J�a��s램�A%z� {��xF�����|����,��3v���X��p��������pvȷ�]^�u^HK�Di���w/��C]s�]��x֪���Y�d���o�\�3�T:^�rU��{Ζߛ�A�$x�戮cQOD�>U�
��#��*�jk�t��?'����#��=0�����.|�?�\��5=FY���"V��Z1'^3u�����Zzj��\<���bឣ�|��K`�5�`s�"qD�s'���:s��&b:�C���8�0���9�G.ylbj�M�a`*�������?�2u����yuN��U�Ɓ�	uj@/��랃�C��ᬦ��8�ϰ�*ڊ�2FY�a�@Kl���6��8��P '�xVv�������2�kZ\��]��ҍZ(�F7za�4w��;��\ip�NZ�'>��WIɧ�*u���P�:Qv3T��ﾈ�؜ZӠ�D��#�z&��������tƳ���{u��@r^F�mXit�Y�SB�;�5�x�s�ܻ��^�3�e	r��#�Z�'�DoJf�:��eL<0�q�ѐ�TKM��NK�نw%G}��\i���QQ��`���^�7/�k������ySg:VV��ڎ��WFK�g�Lf���4��x_E��b�����a�fnM�ڭk+��w��w\���V;�E��O>�2��}�m��دK�|Op?!*�ٹ{T�=6����^N���bQ��@5�:�1�*�7=�n��\�c{�[T.ʑ�L�d�|��ݻ��Y��2RԖ.gW��4s�i� �KU�(�/
��y=�L��-S:v��D��iƳ�7��S8*�gI�e%ii2{ l�w�8�l�T"�	���������Ĺ��5�v���ɉ"s]܌2=r�`U�4"p�������J~�L����҃(�5��&���#�=�h�|ԝ=pq��: i&]j��y ''��Cm#	gKZ埳Q׶}-Tw�]x��ظ=��-�llB��g��@�\� �z���ٴV�e�R��u�PO�㭺�7MDT���B��oI]����M���r�$6��I���B�:��\�8ݮ�Cc�/\�Zgw����ƨj
��9���J�U�諭���g�ֵ/y����Lpr�|��Cu�M�w��%��������+�4�y�)���n��;չJ��1���CW� �P�V�D9t�����ɦ�h��q"1�gg�$+HQ����;dd}�||�Ky�n��;]����*6�T2i�\�i�8!Zז)��.t&kL��^49�u@f����6)�h&v��t�)<������ӝ�o�����{o$�K���!Z���r�4��c�OD>Rj}���X�s��k������d�܉�r����a�	OȚ�r���l�qzg��-�u*5�`U��@y�������v��dZ��:5, ��C���>�k�?/���p0��p������6k���������`u��� +i��>�UXR�����c���{_W�WR.��d��jz�^B��ޢ�nz{�b����?�ԭVE-�f^ *��Ⱥ�Cd�#M���\s����j�Շ޾��r$k��'�.��YZ�[�|oh��p:��/����Ϣ&��iU�a�K׭K.���or������Ds��_R*WW^�wX�����l˹���x&"\�B��5��a�V�Ǻ�f��<�Ģ�Wh�˗כռ��N�v:ݖ���u��;)�=x���z�q�DGIG�;Z�pO�ﾈ�>λ
��&pI��Gz�
���t]^�M"`�	h�O����#O��?�h?g�n�me�ܴ���{r�$~��qT��}յ��,��(���"�p�p
�������j43�ym�r�u���Yջ�p��k����t�c��Cj��Z���!0��z��&�HUyS�=���u�ss�[F��mR�U����iY˴Ӯ�".��YU���S$A�L�]����G��=�h�u 3N��_���t-}qW�Ν��NS��{���h��x+d�Oϱ8��EJ 0��J�iy�$B�K��w�uSw�;�7=�B��^��[���zoq=�s�{ �N2�Ib��>O)Q�XD:�Tj�>�xP�܎u�fٯ[qok��w3�� 5���u��}���/�]j��E*���x�^Xc��iXO �\�Kdl�mW���)f�ÜE3�Ԙ�iٓi�F�F�#K�bԲ�\�P[�$�C������iM��n�/+���smB뿐�N�E�L�3Pܰ	�s��w2F�'���mbW�G�'���:�qZ����>t�0�5Ooc=��nO�nc��.����X�;��l���,�sU-dA��g�&�Wp�FtF�����*��3�)�}����X�֚�q�J�Y0g��d�oF��6n̷_�� ˳1���Q�yX�����7*#z��q�����i�F_Ŋvm���u"��8��ݘ�Hj��u�61��ԟb�q�HV�����|#�K��!����D��5��ѻ]Y��k�����?HХ���ي��!C��l�lv>�e�Y;Nc"xS�W���ҥ�e{�o����4���V�H9:j�9C��������Mm+��]w^��86�:m�O{ϳ�y�a�Z����@͝��e%v����*+��cb�ho.!����௶!v:��X�c.�?�,[�������W�����W[ˈzˇ��D6��|���S�e��2��4�73}EL���s���-�R�4��=��qɍ����B��h�Z�*g-b×��qP��u������_u�����Ķ��U��z��M?�YʈUNj
{��0���]�����'sN;I� �X0!X��������:+����)ߝV�����`9�zsu�7��!�H��:.��J��-e����n���;Whbv��Zkx@)�=�6�bw�gT�\@�ނڙ�b�(���`���=�rU�+:��j��2�@ ���#��;�W6�f����Y���I�k��U�r�wV�=��얣��Ң��2������5�6�>j�|�8�ciWg���{�j�
�^�ݒG�3x_)n��o�7�>���BI�2�^�qU}���`8���<Nx������bne�7�y�is�p��Qi�-��Ќ�V����8���Ѹ:`^�e<������o-��I9���w\�@��Q���M���B���J�е�xm��_P����ڻ?�w�ž]�n����<��C��57hOk�Q�dk����ݚw���.W��\�N$�cr�����=���?�g+���U��J�3��Lż$�o\�˕����N�o壬j�7�c��\*>ldKMך��gaڈ�;�0�59u��v�s�R|kz0{�ͧ	\��cb��{��W/�_�gd�������4��[,��Uz�v��{�ՍeͶ	c&5�ӧKxb��;�5R��;789����7:����������yN)�'���ә9�)���]�k7����V��p[�<Ȣ�}Ҕ��S�2��:�bV]��"��ul���������8�Gbn��;�`t�S �/�iAT�R����=�O�L�U����ŝ��?q��c�S��5Q�:����c��\�y�`J<h��������"�q^�2������*|;���_]&H
�U��*h����Ł�n=��jV�x֧�6��9N�+�w���p���	2�s�6�f�8j�w�S�k�r�b��|�h�lm9fQ�HTopк[R�t����a��sSܲ�Uxm|�J�|��Sob��.�z�Qh��|�ҁGE'@z��V��n��mr�i���2�_M�7ф�u�V��<��
u�~��&�<�������5DQl 2�E3$���۱^�}�)����E�8EB�]_�)��o��okngG�����yۛkL�5ʶ�f��M�Tkï�:�\|�}V����C-����¥h���(�-�Z6��:����J�u��)�[R230����_t%]v�1ʊ�u;��5\-U,Y�d���WZ8�N�vu�Z�͌��A����[�Η��c�㧜��Z򺘥�v��-��_u��*�-���|�wlS"��2�UU}�}Sz֩=�K/����7���w_���Vy���|�je�����htm��f�[�)�����aY�z��t?�;��࿡'�g��z�^�Mf\���:�W�y˼�9������|%��1D�ظ|�.ָmo��ݙ�Ko���PXnҳ��C�:����T5�5¡��K����vs�4LJ�x���n'��կw���yt�v�j����>��������QY:��Y+u���=����p�}q->�+:�]�Wՠl��A�}'�,\�Vm���=.�އ�}��4���;u>�<���zt6���cwZIQ���7Y����}R���ʰ�5�u�t�lҔ���]��k�7��w�g�DB�P����I�S�����D}wWR��P��!o����QЂ
��Ἢs-<�).�e��Z#Wϲ4�_��໡o��W�(�Л1}5�l ���sApp"��;�G�ҒY�a��v�7/fj�n3J:/�M�[Y1E��2Pr۝P�yn���T�N���$�h}tnu�5"�-�j�g[�K���k��e�na/��������=t��P���,\��'�着�'f9���L~��m?_�1��}7��̸ҝ-��r�������EaNn�O�]�.!.�ضD#�1
���v<�u��k����#aZ��e�IL܎z�ysw����w��D$�5�n5�#�1�ȞCg�kaԞ;��5��F�JA���{=����t�W�Ѩ�ᚆ��r#]�?c�i���QU�ޯ;גN2V������)~~}�j���R���ᚋtη�����|_bhͣ��d���c���+W�ڝE�s�	=i[*N�\Ø��g+S40[�����]�v!�U79B{î(��|�-��,5�1M�z�n�a��K��l���������g�P;/,auzc�qbr�s���NkUO|#���%��W�=�>�yY�&|{l��Py3D�,�5����Zƫ�u�6Z�lr��6��|��ί�aUZܔ��Iu=�{3}�F���6�'ͥ) x\oU�ݿ'W����b�/㶱�A�5�#>f�ZS��nIH"is��{���1�=z_�f�ս�ݝ��&h��]^���2ۤvB��p�Ցá,�KL�� �V�m�;���B�Ҧ����'uC���">���%ol���=�'�좶�W[ˇ�����|�z� d�ÐV���������=���G�_��u
��)O/�[=iU��[�h��&���Ob8!yw��U]��G��;��H߯�_���㏹�o������v�C:�c9P��!Lw��a�Z,'�qK�X��z�o9^lk�v��o�����k>g0RlmC�e�>��H�b�췏|��-;�p}���\��L�	���H�qGhe9�T6�5Q��y�\��tν���v;�|�Od�r	�ˍv�Bu�acq�\��1��:��̖�o(\��j�E��͸�9�]8T��ܥt����[�BC\{K>�y�K_do-�ڵp��z����E����sԋ�}]������8���~��[�Z�:���'� ��3h�U�y[.:�Zm��c$�I+k'>�׍��F��f�a�:�ثg��EI�:��F�$��#���Z@�/]F���M��ݭ��h5�i�d���t9��.SÑ#+]ʜ�	��V8ST���>�gf�,;i�j��1���f��Ws|�ud�˙vg*o7��ތY���R]f��w5�*�el\^�$�t���b�.���T����GDz��ʢͮ�w���6�L���7��g�9wd�x��A~���O��:y�ZX-Vy:S����|�4鎱 �Nͺ'P���ʞe7ͭ �Ñ�v�U�,�bT�o���ũ>
�J�}n�� ʾ�s�����&�
K��Ԗ:��wn�Ȝ����D-�n�}e�V�YO.A���Ί��Р�dN�Ђ�47�M�.���@�rn�xZ*�|A�W|�0^|��;#Qj�;����)��Iwc����D��.��[�~ǲ�H
��:$�LYƔ56���	ʂH�|/��4�/�j��{"�)c�Uxs�3����CW�>܇����J���FqgM�:=�n�\gh���\*ĳ�9�o�)�5�'v��6_��k������%ݗT���9G�eTR�ޛ�V�Th.D:W���c�����C��N��F:d������mu��XƷ�����Цb�.�),|�#Pu���.�6�:�|��%�b����vͷ�Y���[��lr�Ӭ�TyjK:`{���������Cy�s���^vqk6�G�n
��e�I�EDp&vٷ@-��q3a�n�[E.��Ș}�XGj�e����˩�)F�03�^����0v��&q����W_9� ��iJ�n�g\���߀p��{������T�[�QW��,@TV3*��Sq��lQ�� �t��+7J.Tȧ%�<;Y�����֬R�`AQ��HլёV��)��� ������,�g����ۨI��j�֯�9Z+�]�����w)��n��r��B�{����Iٰ�a<�Z�7r���[���9齫�>҉cU�>�x�f��"�P�R�d��'���T��8r�ʺ�ʗ�hk�ګ�/u��Ҍ��\$��H�w�Ai���'\����(a��z);�;\>�Y�}���! ����ԉar��^c�%H�ub;�^:�fLP�#|{��k.7o�\R����f]��Sw�VZ;*,ӆ�v��ov�
���/p�ѕ.���QY�5!#�/�����/T��It��i�M�uf>�oh�*��W��W_2�/ov�].$���Mv"RQI�@��[�wMV�P��o�P�����!�擇���OQGlާ�����R��eB;��k7{�ī���U�{�6�K/!����V((%%F�n��{m;k�ӵV9���8..5����v�o&�.˔0]te5|��VQI�����&Q�Tܘ��g�]>n#�R|Y}أ�f��B�
��!�u$��!�Ď:茑\�s���wa���
,r����/��fl��vI��� H�F)� f<\I�1$���#1"yܒ4�hD���R0���wt��λMΙ�l"���x��DɒJ2�Df)�\��� #)$BG:a��c<�d1(���E!�CM��G��v䄳 @��LÝ]��ĔR`ġ�DHBhP�bF`0��)RȔd�s�Y��,B�#4$�s��J9]�I D�K��t�bc%���2`C���F$	�;�$�D�����l��`JA�I�XWv�10aI	��L��F������n�Lw��aط1s&�T�p��Q��oj#���븪�E)۶�,���S��o�vmٗ�:Aeh*�o��>������Y���w˄�kY�j�銹2�p�}G�bN,�4��B�9�׉�vd��'X��S�. �[k�7�O�iYU8%������Ψ_�=|ZV�VU�˗;���Q=��|y�c"%���}��wgaܨ�@7V�ai�"L��i����z�c����#iBV6Z�lt-��)��_>�2�7r��R��/�꠰�%gՠl��U%�ʂ��V5����wi�5������=���N�pwˠX��7Q�zq�Zю8����<�Lt��T�;�<�69�k�y�o�/�a/��
�;���D��lNEh*��әY��&��4��rƵ�V���=CGO�Tk�CcC.g����\��s7a�w_W�_uÖ��9�s��E[ci�3�!C΍�I����(K6x���	of���/�Kxf�Ҹe�w�8�|��|��:1���D@�}�z�G��w7��T�4`��f�f��R��9+GwJ��v�2���Au��<��}��n�n9JMg�\�')���&Y��R�Ydun�`�utY}7��ml�Bwrz��v����.��<�-7��Q:��\��}�|�۽�;;V}��d�5�'w�B�6��3M�7Jɓ��2i;�MG��r:xt�� �_��
ܚ���{�w˞8|::_Z����],Of���.��Mƻ�g*#^o��?*��}g���N��U&�㮖����l�dִ�m�p�[p6��f?#��%oE���?zS��L��{���j��}
���ټ��ڷiK���w�a�m��w	dV���}�X��.9ú�+�j�o����qՏ��T��ֲ9����{'�_S�F�����_#��f:=ht�T�c���XΥ3�tg�������'�2g#����[�fhn'�y�e�m_�e<��o���(&���0���Om�S<�建7�rJ��}�mj����DV���[����҂�ٺ�i���zVv,ģ����_ɧ�������U}Z�AP`>R�chgF\��Iw]7���:�t<��Hx���_Jꖕ��LKi��١��&^r��b�&п��S��,�5���qt�.�v�}Ӻ��ε�o7�o�<�6��$T�-���e2xݻ�$��@�I�n4v�YWn>^��KdlOR�V����j�G��!�̞���W4��*��u��Z��>e�jOn �nŅ+@�1@6��Jm5y.��>�+U-��Jy|���|3k�r�:nhAl[�wr�=J�ډ��� ���T}|t-}5_u����{k5Ѫ>�M��{���V�r�|������P������6�&���=���9��c��ŝ��g��{��B���Jۼ�ҟ�,���G��Y�V�n��b��ƾM�v�0��R�J9��ak���n��&��ZiӾ�f��w�R�k�i���I0k��k�r&5��������+������r����ܸ����Y����rtjӆi�j9�ƻ ��3���M�K�tJT$c�W*���ٕK_o<��n����5?/U�K/��+x�f�����^�˯�� f*���V������pT� }��g�,s.��zx��ջZ�L���Jlxm1�5/��0nށPuc}��<9Pb�^f2^��z�z`�Z�9=q�����2-�*:�)5[ھ��F�V��gR�)�<�*sU+ʉ�ĦY'�;|ÃMJ��b��y[ �u�S���8aD��ꪋZ��-j�.v��H�~�mGΑ���.�{��g��]F�>�����|��]��/\6��9�d���3(��z��fB��y�s}���Rm�j�uvP^�p��t�]3o����u�	�6����}�e����λ�Y���'G�]X�j�6�����|��+:�a@��Ub���Bƚ������]R_W�:¨Z�X��ކ����m>Yy��wqn9��L��C2xh�\����*�'�nT*FW'���%G/�#�z�7�V*�2�G<n�XR�ޘ+��Q띪}7s\�u�¼on�i�%�ژ�vͤ����*�l_�����x�2��׽�n>]��!�J���	���D.��EIq23Qybz�6�u%�w�b�y����٣*;�L>3�Sy
����}0���no7��t��!W�Q|ԻG�VL6o~M�݃��foK�R�P�-i=u>\�:��ޔ|W��p��c{� ���gpo_+��Sc�A��6I�v��Hdk����[��M���z�n
�I���9_E���S�ﾖ�6��}�������j騕�;��r�-f�$ÿ����q�ɛk֤��CR7�XRl*�+r�;��[K�;�Tj"�g�S���w[����N���WyFFE��*���<�tU؟?�fu����sV��kK�lf��U}��k0/b�*�yd�a�|�j�sԽ�sc���+7���ܝY�7��;8��p�f���(z,ͺ ;��<������\�7�X�|�_�w>�]�c���7[����=�~�H�}��b���e^ڣ�V���
>lg��7ך���u�V���뱴��Q�پ'�ps�uĹ���j5��cb���"�jcy�}T��]Y܅:���������'�J2x�N�R�z�4�ݮ������7-�����}��l��G_�2tѪ�B�x�֭��^�3Ɉ�N���f,4fj*����8s��i <��OWm�h�Ghe�~8��@g<#aص�ъ˷�nP��+zk����T�W-̧&v��ف�}wSv��`�j�nY��k6uwV��-Gh���5}b{v��uƤD����W[I��v��ڟ|�{p�5Oʈo��x��,)Q�?p���'VP<H�:�$r�[WN���Ҕ��9k]��mC�s�%w��ԉ��5��tV���>m��b��w�r��=��8޷�)���r2��ԧ5�2�cf�v]:|�\�����p1-]p[٣M&5�-����;k�׹߬�ۇ֌� Ɵu|0�/MD���\�s��t�� Ke-m��W��Ȣ~�$��w<�eu�z��Ֆ�;=j��;��ߐ�=�Sӷ�/j�My�WN��0[Q���Lk�9�kj�����Z�ENt㏝�����r�\4��uZ���ӆi�k����c�R�־�v�V�v���P���徘��~�V��%/q8j-��K*�����"������y�c܂��7��e@�{T���R�_�=k>�\�7�Ȍ�BL1.X���r�(-�'�vQ��+�7\�az%c�9�IX[@���)d��ЀA�ި�Z�ǩ�9�K�w�OD=�=gQ:u�*�W�����(5�r�.�'uI��[�R�}��]�{L���&#��i�滺^���*d�x�NU+O�>N��{����ʬ�CC2����wh\�{AJ��/L�OOxa�%m��[��{%�ӭZ�o����e-
�X{l�Ҿ�M�����s]�#}�s2vŏ��t����/�{�|����n��u�qR��g�I�X�=�ΩQO����[C�%}�|[����m���6K�C�1�f�9C:������K��3U}��]µT���zǡ�Ci��V*�C�j1�"����=w��3�2���R^�[5
S���[p�=�y���4�8��zL�cP����}�P�B���R����B���B���}]h�fY].�aj����q�e �����!�`����\����iy*wylʼ�����ਆ�ӶP
�%P4��1=�楐��뼗Ֆ�a���_'ξm�l[���*����t��uyTv�"�ƞ�=qY��Tx;��=�Sk��vl�+tѫ�����Kxc�yS�~j�e�Vr�p^�P���O�r�|�N%)ut�ZW��oE�HQ�׋.��D��.�(fΉ]��[��ٕgTQ%)u���cg�7]�6\�o��r���_���?G;��'οD:�;���B}E$�j1p�i��!�!�,�bp��ힻ��9��y�S��ˌ��so��/�:5�3M�����=o�r+z�g��{��<Ж5��/_���{��j/j���Nu�7�����~!��՛���8e��T$�o��m�ڝd뺰�Fc*��gKI�י�Oc�IjY��Q�ٴ�����[s�{�X	��C�Qp<�|��V��]�����v����k�9Z�e��'���z�Y��%���h|�T-Tt�Oꋪ�}�o�C�S�;ץfx6(��S��]*��o�oBN�;�Q��+-\lT-o.M\�|���Y��R�s�UH���{���-T� ky=�{�v�m���r���6pvS+�a�- �P~z�Os��!R2�<�ڹ8�|cVǎ�=nH�z߫3��4��;��6jQ\��u�e��1��k��	��9L�Jp}CT���������E)��]�d���ak�`Nw)�D��ޥtV:���F��LjP���Iյx��g�_���Y���y{�m�4;^u�x�PY�鏊�:ܨ�\鮘kc2�mp��c�Y��ǻy.������63���J�߳x�?@KEѪ����sw]��	]v����yKJ��w7�)66��(}	Knt��A�M�����a�eܕ��8�f�ϻ�V��ض6ȕHѾQ�e�49��lwv���Jp���=rV��F�:\��-e$�Pˍu���h�7�;�jvy�~v�W��W�[@��� �ʹ�}�is�&���VuT��H]�Mv��v4����t��6���EԦh-������<����[�,
-y�{3m�3T֪���m���7�_k�u��P������4��y��=��ܕ�n�'{/R����k#]�y
h�b������s5����Sw\�͂����D�>wK��J��%Y���*��V�zKy椵���p뚪�j���5�u{�0Ol�����U��N4�5��ީ��\F(}<qʷ���yA*��ycҀk�s��c�9���a��w���;�;�;�\�6i�7l�[��T\��U�V(4�Fyp�����w�f�=9�꜏odvS;;9c�y2�~��+.rnf�}.`v�g2��1D�.�6���k�n8։���XwQ�Aa�q������qgrz!�TlWt�����h�Qpʾ�v�m�y��w�����:in����=`��O�,�f}�d�[�m�ض���Y3�!��O�Oz
ΨV��6`�1���ˮ����՚��[�sF\*��6���j�xW���/�aJ��*'u��
�)�j����sݗbn��u�Q
S�X֯�ڇ��:J�XZ�.�y�Ts�6�t�=e����3����}w�Ե�D2����>o�T[ckvzf�z�X�7Gh>"�[00y�Z�x����5&�g[�������ܕ�����4��׳�� �2R�����cs��]��U����GMu�k�x)�pw�v�D¤'��\l��sr�K�$�D�yފ_�~M:V�Q�E�%�����`���:$�a���v"-�k8��g��ӥV�d��r�n)n��
�:x���zF�r:�f�2�������B���X�LV8�h]��SF��y���H�rSљ]��jΔ��]�z�\�έ�*�-���P5��.-�}}N���F��w"w8jpn�׵Z�z-U�WzH\O�:\vU-�Z|b�oE����	�6�l�R)�:��� �M���w4n�
�9R/gM��J�����em��w��
8Q�;KeF:�|q��1�<�i���7V��'Zvj�l�(��koT��^��K��v��|���+�V.X��7J;��#��P}B��M(G�֛�XN��ˡp>�5'�2����1H���o>���ጆf4�����h�������vh��
����mU��yS��V"l��sW]��J肔���V+ws����H�x_5��з���I�K�"k"�Gۤ�.s�f���y���g]��֕B���/e������N��ŭ���h��]��'t|:�.G�k~��j�k.�ws���Ew3�u�Fb��dYkq�n��JФ���+�!/�����2sG���@s��Kg[�����0ۭZ�V-Ԛ���7������ ���cz�+\zr����J���G�L�.
et�ks9�U��6,l0B�'@�|��5(,��z������ծF� H{Yauwʭʘ%d��i��+��Uۆ�*,����5��w5\km>�!7)5*+V'^hH^���mg
�.�ft�mkϻ��san��O��'�uݻի6T9���ӂu��M%k��\SQ�T7V�i�kwz,M��>\�V�A�jφ�@���Wv�J��[Zw�n��uX^1�Ut��ic~�E���@�ԫ�0]�gv�X�.i�e�v��V���rE�L�=&YH�!x%#��º�v7ۮ^��gX�P%��G��V��9p��������uɮ�r�qܥJ�,�w˫�yy0n����f�e;q�D[ϞWFgU]5@��y��'�- :G,��K��uĖ�R�9vi]�RqGUŮ���P{�_J��8�601�	��\��=l,���<���ȍ�`�uwOp?��P�����G�SEr�X�}�x��˩���g*ڀ��	��"�}�b�~"���Ms�W�1�
7If�ӱw%c����B��4�\���J�^�׵��)kO&g<���pzV�ג�Vag۱o-��s�̳�[�R�J��F˗Ց�Ҟ���M>�2t��Gm����=au�:c���<e�׋�>re�[��=+-־�n�a��o����m������Ze�⧷SCy\�|�>�i�eh8gl� �4Zyp�u�_
I��UoQ�����It�Õg^��BX�;X܏�Q�LŅ�ҩX���u�;Ye�p���/L|Q��CW@q 
� �U
��@"@�I�$�$0���#�Gu�wt��T�J�Ғ�J �dȰӻ�(��c�n��s4�r��f2��Ii1���.��J�˱���RJic"�2�f�Pf��1
2&@��LJ�f`� I	"�I�]�&ILؠ�"i���C�1��!,I $D��B	1B�	 ������#	A��
0L�2ʂL$���K$���2�2��ˆ0ܺQ��Pȥ$�(0l(H"�&��!�Z4��R%��*Fi� ���$̄ɠ(�(�H����~P7{ugu&8����W0��2k�f���7���G�42�R�i��c�l��,��4������p[{V/GD�Gﾎ��M=�{���fo���$�5ۍw�ƻ"c���Z��;��ts����y��Ô��Sy��]V����8f��i��׆cX�ySH*��Wp�љ�j��hgWE�8D�ʎ�[f�W�n��/n18u��_CYQ9g���.�1�iΣ��^���[�W�yB�\v��|�
���I�W��Fp��ԶV���~�B?Vl�Z)��H�<��հ����K鞋7���{S�1{�7��l�4����l�KB���C�~̿]����N������m����b	�jZ}q�6�=U�v��vb9W̳1.4����ަ�IUͬqհ�;g�ZB��%��}q-�����zV�J�^�7s�{�o<2	�責ɳ*R�=�[������i�Wľ=g�32l��T�GJ$K��RT���RZ�Ke��X)Ycj/�EE��4�2SxQ� /m�%����`V��U]ݵ��N�pV�44.Z�Yt��w:¸WL�Ԇ�c�X�8��Cn��8�,�Y]ǘ�;��e��Cy*�.뭱Ƙ{�e�yl��M%˝��"^��]�@�1�݀��(�3,�&Ζ�����۫w�yYBR�~�;��Gs�Tv.�Z�Y}�h�#@���/g8�%y����^/Ǌ�:�ЊzD0O{`��\]y0�zyk�ql]a�jܺk�;�sZϙ���l�ȅ?t��h%��y��9�R+]c�R�,��CS��ڄ��o���q�l�OʗJ;��CW=zEB��wp����:�j����5�I��c�r%;"~ xɯE��\��r���CU��H�2�ٸ�Ɏ�j㓣Q�3M��.��y�m�vH����X֫���ln{��=��󟣜�^nI�;Ц��52y��i{�o�9VۆoK�լ)�%ޤ���CUG�}c��d�ξV���x���Ӗ�z�}��~��F���0=��ns7ӹ�5��ڗ���ښB�rqX���O62%��n�o^�}�g+�̢�ȵ�]�� ]����RNY�N�T�v��{vP��K%�>�*�5eg>�&��yS&:o=6����v�9Z�5���QUjR�d�ژ���Sj�Rå�Hn-���P�"��]�,�*h�Z�I��Wt:.w|�Y�V��v����u:����}.vC�U�@#��}��O~�8�����ܐ4��׭��Y��m@�秶T%_(د��{->Q/�Y,�8�J��_gU���T���p� �/�'TKU+�[��_v��[9�v	���������u����+@ق��ʢJO�J�T�sz��c��ĒP��3�՘�D�69���=����n�XS�ࢠw	��'�L�F��ީ��ķ'-������䵮ϡ�ί�3��+����a���9K.�֊oO$;{;a�w��|��2�_3���m��r̢�wtX˽{wo9�%�g�ڜ	od�w�qJ���I�2�;gm��jₚ�W8�L&+j��ʠZ�뚕�5��:\���y���C�t�T�9J���Q����Uq�Q�8nP=�Cm|{q;sڮ��U�����%���ڄ˞@V����R�Z�+}����l��1݋_^�e�lXVj��i\q{������4.�\��y�̘1[v-�]}�K�gv�W2 (���e�]��9ӏ
=�QP���>��k��t_i�5]���X���%c�..AB!\�m>��xh�ud.t݁�菾yG&�U;�<}	wI��h�Tk�9υ����Q=�Q���j���S�j�kIi���Zn��T[p1W��B�g�����'z�$̭k_'���w�j��Ṽ�&�J^�؜kY��S�/�2��������m�J�_q��==�Z��o�D�����E�p�����3��	k#��3e��TU��s�Sp1D�ظT|��x�g��Oz��~��^O{:��W�`U`�W����P��p� cb+%\��5;v�'�L9�'wo����eR�����=�:�
���Ng~�Ƨ3�,���W�y6�_��낳�vU�l���NI���j�_%*�*��i��6��|�z��m1aJ�88f��3s����7x\w�hp1�}tR���)O9�Z��ͨy�):o\e7�"w�7��m/0�����+k���t�J��\�����A�U��+h����^� 8�gd]y��w0��������^'y���nB28<R�D)����{7�.�"fP��w�e�Ӧܣ.�31=��ed�����%	�h�A�㴻U~������ۉ�������_}w�uB��_C��h����F�0r+.ì�]��ں���}F3�=�,q�%?�W�k��h�	4��t�wN���#*.�_<՛���`;Y�,8M�W��D)���h%>��[�q��t6t�d�ۄ/��:՛��خ���hO�q�#�*���^=S6�?Y��m��j������H��N�J]�0�!>�P�`��B9�Ș�6`Z�%t�����1a6�:�.2��o5m|��_'F�ӆi�j9�Tk�;S��Gb�辘%���N���axd젔ˉK����כ��/o�j��\"�Lt�yosw-+;K�ɗ�(=ꓲߵ�#��*��]�/ 0j�Tz���z��\�忚���h��*<d���ڠ�48�%˺:�ek���r��k6UOlu��:�����v5��8�.�^H:y��f��Q��mRDo{�j�L����g��g2�5�ib���{.c��X�M��L,��˥W���G��':� ��ˤ
�ɾ0}���V�[s�@RjY�l<��K��f^�Q�H㋗Ѣ��1f�Mr�vv�8:�Jқ{�w��w��t*�cb����O�%vm���;�S����*a��vxG�-r��瘷��9ζ��=B��,�M>�|��+:�aO�i8�=x)�nk��9�RuI}Q�NR�*1�oCy=[OP�I�뒃ҫH�Ȟ�Ӫ�Fq��d�2Ѓ�RR뎺-J�E;s��H��p{#��mν���U����*9�v,)_oLG����tsK�~��FIoC�#ۙ综�G���_oU��!��wF�H�N��gy����ڜg�T|�[����J�ֲ��l�9fQ
b:BU�c��gdwx����7��}pG��N(�6�.j���3�+g!J7Q�CM�b}���y��d����e���Λ7�ru�u�}F�$ø�\k�rV�؂w�Ԟ:���|:�n�mQ��esٸ�[K�;���N��=�j��;��6�96�Q��f��@^�SF&�R���F�M����}�k����nd�Ȓ�%I��"�5��5Ĺ�u+��غ2%ph��.@����#���mL���ݬ�=k���	N��������qyD��˽��̭�JrƊ���a�/y��;�Z�sx�Y?T7��5�v6<��g�~I_?9Ns�כ����%Yf�$=�7������(�oj��xn���o�b���u-y:����j�֞��|�i7�;��yi8ֵ�ޏ{6��7\�e��f /�u��O���5l�o��X��<��x�޷'�mD�������KM@=��l�F�R�����.�,g�L����];_�}�{6�H9ܲ�Igq��y�����r��f҄��ՌlR�or�iF[۽]�[=[܅�t��s�;8i� �/���T-T�ky�4���fw^�ٚe��u�O�ⳕ�,)��hQP*���뢒���aR�U�ع�S��nԶ����OC�y�n��X�=DHz���؂�d��I���%S����ʟM|��%�k�z�x�S���1׿f�y����%&}ʰ~̣��7jϕ&�����m%3B�aY�vP��P�).N�oX��Y�k�^�X�(��=Y����1���Ό�y�s�v.��9!3�NKy��(����>�O���Y��е)�YT�_o҇t�yS�\n��!��vlب�-ܝX1lK�A�⺾�����J�׹�}��-��商&^�ަ��9�Y��eD�p��#A)lԭyq�*�o��W��c5>*Ol�ۦ�9����8�@)F���sQ+rj7y�B�}S����(:�]q�H�;C~���k��ȕHO܆���WnME�=��Z]����q�=�f+�Ǧ�˕i�͸�p��k�&9�[���v����Mo���y���>���څ�j㓭���nl7���f���p]�*�oA�䨤SX�M���{��Rѷ��^ջ�����Ƶ��uc�SF����X�Qu��C�3끙�6��y�+0���,]�o9�Щ�-�헻J��W�F��U��h�|%1�1Gb�9�CB7�T���֔�݋�|����y�xE����s�����1�╇������*��t�$�ƛ�i�|�IpZ��ѤW�-�^�4��-��ѫ���4�Z�z�x5��\�D�S�t��C���U�s@!X��*U��Omc��f�ʯ}QV^V��_�l9�U�	����ju@x��6-�Q�䱗l]J 1�z^NQc�wq�}:z��=�ݼ�a�O@�Fy�G��[�؜	��+u�{۝R���T�ᭇ���O�Zz�M�g�V���{����K�s�K�E�ڢ뫪y7����=9���
��t���K�8�;'��ޣ�/|v��'����]��>��-�y���	�)V��*��8����v�-p,l��ޟ���C�]��u|��ӗ�p�>ު}��%U���Fj���}��V�мC)fa�;��������⺖���>Et��sS�v̫�]��y�;��m�S��:�A�{�������&{rH��_n��N����m�w���R��|u�3ξ�H�G��W�m^߻ێ3x^�R�%�=�\èO��I���}\U?a����)	z�L��}�R�[r�8;ٗM��jڈ]V�#��_Zp�C~��ya�rvU��6�S�0ӣ��9�IμԷ�&v�j�����Fh���3�Q��*��9���ߘyJ�W��a	��2f��M���ܮ�8�����r��5��|�����t��v�]>�oa6u�4;p^'.�uu��K�}����sӼ�r�F�����愱���|�L��s�+^k�^tF'Ĉj���6�v�m�r�"�1߼�j�h����~�B�	��狟#`D���Q7:�����'�?�Z�}�CT���&^x7*�:��Un�{�<�M�ѵ=����[W!vr���ldK�M�{���2�iS�tv?�p?N!��w��^�Y�ޅcV8��q��C	s`�Z�vm���;�E1݈�(b7t1&��龹�	0{*Oum8J��W��������W�Gtw�4�����
�N)��z��R{�j��V�X���z���{�,A�ƕk;�sn��p��V'qß���A��TIK��-J�E;��65�V5̛E_-�j�:6�hv��8�|�7p,)�����LXK�����\�������ǜm�H����_ą���Χ��9FQ
{���џ}<�;[������H~��bv�fѻ*�Y/ZА��c�K�J�&�E3��&yAG�ظ�3�2[N��f����t�1��M�L8+*>��n���w���c�mV67캖�i.�愸�.f5CE�b�[���ɪ�P��R氚�-Q��Ay|�I@�寶P;$�wv8�Q�]cN�	�J9k�*����vj 70,�]���_0��h��7�t�߻�ɋ�RP1CJ�B�1�Ư6���Ԛ�n)�ˁeҶbQ�[:��/4�Y9��5�n�%M�%Y8R�*����[�ՙ�h�]4e���W%�L���T��f��3Ya��)�n�(oH�9�q�x�C}q%:�ܬ�U�:���{pMF�����&�)�M@u�{�n����A��0~P![8��RU�u��++8��+�8RF�k7/idN3t��%[H�����D�� 0��V:՘���&�ZE<�Z����nJ�D�U�x�e���=4 ��5�N���e+�dE��#�u���Vy�}����칮�������z�˜������"u��K�ddtɫn�T,9���B\�k��-��;�Y/b����˩$�Zt82�ݫ�>7d��Y��S:��K��N-���#��=�,�)�.]	k*������pm�9ǹs6o�ˮS� �vR1oV���dU�0
z9q<�kN%��[VyV�[�k"+T'���Em^t���"�A�vwC�E;��o�%�K�	e��
�7�N�Dl��Fd���r�!�mEoZ77��r�3v��&tv'2U�+smZ�¬S�t�
���9y�Johh�]{�����^��]���6�Yz���UJ���^�m"M�HC���*v���\��m�j��PV��%��q�]Y|���A�����T���P�AК+�tiz�[l�^F1��ï���e>�Z+`���'��7N_-�hdJs_qq�����;�݀Q[z�^Ɩ
C+���t�5���x�n9XD:��;W_=�]%¬�-�U�Y�Wt1Si�{�	�� �e䙨Z4��*#w�-��j�T�t���}tU{ใ��:.435I/1���%n�&�C)K�*�+pw��pxF�G���m>�Ʊ��.Ɔ9��l�.N�%!Y.���N^�]�|�wS�u�[���
#v�ZWv<�:�Ȧ�3pX7���mqlgٔ�;�ɾݜ���t��լ��]։p
Հʉ�,��BLh�]���w&�}�mޗW5X[�u
�i��:N�'ׯ*dw;���.2vsy�Ȣ0W.�l���}e��CI�� /3����r+�Z��"����W���ȹ0�3GA�sip�4��)e�|� `N]�O\ʉq��:�.c{y����b�E�q��zl��0 �����ug�Ǜ����X�u&��b �bˀ��@j�W6�RG�!5ڔ�0z�y�ŀS�xa��m��Q;�����k��2c�˺2�z���?�?��4���DbKCA  �0�I�,��Ģ%B9ѳ�$\舙�A	�aQ()��heΥ��,�4�" ���E#Hfw[�tPȐ��:@H��p���2�N�Lf0&d�"dspd��!�0�d���#I�̀w]c%1��Mˁ��$� )D$d�!�dD�ę2$�R�Dh�d��f
L�D��2E,�Nv$I;�����QM%	@�Fi��]۳""DI�F&HF̄CJS!���dP��0����T�
��`m��c����9q]ơO3�V�&�3�ݨ��O��YR澾�d���r�ކ��o�c��c{�}��$ƪ�������g�S���jZW��Xߛgj�?"����g7g6md8���x��˹�\���-R�IsV��ضD3�*���52�jI�:��v�|�{}��:�� �>�I&�.5����qٕ�������o��t9���斬�w����j��[�gY�N���wV��J�#"����H�~�4��|���s�u�{ƺ�o^��ciy5��g��f���3V靸oj�9��:`[��[6�N���A�J���{����~��:�s�K�IƵ�k���k�k#�̨/���������S��r����.v��3�D��ʞldK������z�ʳ�Ԏ��.S���ER}�4��Z�\��u79BT9K�o1�>�_N�����P����H+6[Ӯ��v�õ�u|]����V҄�l�p1�P���w1
q�Uf�'v�		���+�y���-K�l'�Y~��=�ã;�.�/-�NlQ���Zz)H�^���:�&��������m�7>n���u��9-	����9����Ƃ���]a�h�K��3�\jF�ΉZ[ �W3{����R�\�bf��w�oNo'D������2��/>��=Bq��P�}��;��y���e�s)a�IV��}KO� ��@������RR|��4�J��Z��ɶ���˅]R�y��5������-����zb
�֪��駔���m�p;v��I�},���Z�c�QʇT��	8���rQ�Tovs)�E^���81��ϫc���k�-+��׹�}���lm6����ʎ�"�H7Gjˍ#'�]1A��f�k��-�4�2�7omR骮�w;R�N�\���h5�b��2�=P
UA+\ԭ����.Cbt��)}����s�x)�]��2�]��B�/�CfN6�
ܚ��{5� e�8���Y�6u��6�n�\&��L����ׄr�[A�p�9�i`���>��\�r��|�^s�w��.�3Qm���s^����ugM�"�5ᝩ�=i�y�Z�b���~7��WRs�S�T��YҦK��j�:�;�]`=�z��k7���wK94 ��DMN�y;�V[K\��Yʛ���s:a�u)A�(ŲiM�A���1��� ձ�HV.o_"я�n����$3���_9Y��Rѷ��^ջ����t�����aѶ����k�xubvSb��R�����	X2�TMc�pT�	gMY;Z�˝�K�Lgg�v�&]�<3U�ʦ� �:-Gv.m�M<r�,�\���z���]�sjy�4��͠\�s�*�������[OSx^v,ˎ����"�h��ߚ�_gaڭG;T���۫��g��IUͬqհUGݮ��5�Oyp�|Z{��K����5��9�i��er%G'j�	�E�fL��{��s�M����\=jOn
��0��`����k%�rT~$/T�9Q�?	�iu�u�u
��D)O/�z�gφm,�'��vu)��ui��6�N4�V����
��C�]��_OC�ݜ�0�����ޞ]�9f�;I��h����9FQ�J	`_��.�������!m�ی�����M���u�z��o�C�#ǧgHC7�����)ڪ)�f��ꝫE.��
�r�Ur���`����%p�Z°��/o�����170	80����};�r�Ý�"ݐ���n���KM�v#�c�Z��'s�n��Pا9%�z�V�p�s�s[�wo#~v��9UE�Ƃ{�A�1\�)yj�\�nٵ��g�|���\�Co��q�p�D��s8�z���t�꾕#崔��e�u���[�=�:0�>�_$�5	��댬�"��ҵ@�^ٚ���%^o����3%���Z�ioܝ��m��[��9�7��y��Q�5Mn0����fuK��Z����{V�#������z�����V�L�c}U�X�mR�V� �5~�.��7���s��"�7����y���	�|���y�h���U�x����N�N�����*�6��ji�P�c�pT�c%�����l۳��fW�]�B-7��7�͔�f^V��\���1GW�11Isb�Z}J�ۄ�TFv�5�u�#��I�8:x�TkG�ֵ	F��H(�	e��\�}E���A����2��R9]v���#�tc��b�!S��2��<L ���y#9�}ZR���B��|�>]:��9�&R
�Q�-�+��B����]���b�����U�r�%�*ti��칏�ډ��Ìq>ۓ�������HoK����U9�uPXn������{�j��V�F�|�7���bv{Z8�]X�{��e�+�XK@삠�Ȅ�~�ԭ��];1�e�͈�H�;�Y�y4��=jq�很�����b�i�S+m�[���Z�+1��4��Z8�r��<gG>D)���1E}uKg���S}�c�&��ɷ�u���ֳ�wl��Y@!v�֣�Ah̪MBy�DN���z���P����(�_p�0�Ș�\�Mh�b������Yq��PT6�>/\ܮ������:O���j�+�\n�s���㌊�֎D�;"y��V�w?��\�o5m.x���3E����7Y�����8�n5�#3쉍cd_levD�̕�nrt���}#�1���n��O�}���;�⟗�?{�}Y��	:��Y�y�b#=p�XJ���v��j�eKBhm��Xv,Rػ�&��f�ۥ1W ��*�:�pQ|x%cG'��+�֊�5̉��Eʵ#yw*k���2��)hN�]��fs���B��VP��W(�AV���Z{�>�eLx��=����E��1N�Ƽ�P���#�nh}~�p=N:���eKĜc宇{׻��b�no��4"	�cg9�%c��gJT-�[Q��|�⧛/\7Y������uF&&g(�k��U����N홏e@���VMi�4�,����Z�."W;`�:L�xf��W���sk|�͏Hvyl��jڞ4<J]�xh�T9��;���uP�y}�#n�|�įS;��w�sG�)�Z�Ϣ�hx,����[R:�x�ƾ�+Ơʨr��.g'���hD�iu���ŗk���{NG�O��#�p��+μyH5����<	<KǕC��.>�{um�.�-r���N�]9��=�S����U�i״��)>/�}����W��<|��Yp ���/G�a�h~��wm;�p����@��>�}��_�
�W������'J����w�T�50W{xa$@��V�܄�|Q�8 {�d0�IJ�ϑ��R������_�lG�K���������uiy�Lgz�Du:��>5�px��^��t_j���q���t�z
�}&;��t�2��7�ٺ�XVm�%_c~�z�Y��<��}�h[�䖝�Y]"U�
�lt�.s=s�opĺCş��W�@�T��V��4��;���޲U&,K��{�H$��9���C+�߸�]n�[�t���ftq6���g���y�l�H�?dz��Wٗ�c^��+�v��r�{E�杩7��@�>� ;�ց_;�B�O
�3/�q����Ui�3�����쫵�\��>Gh�V�w���j�N#�%}�z����[q~ԋ�U���^�-����3�=��%�����+>ާŪ��П���k�W�����=~����3��q���L��^[����'|.a;���\T�:-_���ަ=q�w���vFF�P�K؎�X*�2)�9��]3��ή��>�c�;�zR<��ܧ�^����b�U������+�.}X	�鱯����R��[}s�B�[hL/:�(����n��j�u�Zo�R�X�@�:$z=7:�]K�UԲ��3�#�Κrv+��>��{��S�z�.|Jq/�>�EC��1Y=�|����oYni��,;���7+�ݷ���7�ϱ�G8𸾒OT�����lkJv|��fO�?Tι���B}7�Vw���mi��������<���nZe�
;0�cs�9�r�9fe\���W���cUc�cj���#�tZ�6�v��cn)�s{sdSl����Q3ڼ�֍���:�H�A�W�W�i�b�>��D2)��ړ���M�+��M�L�܆���iQA�˜X����G@\��X����A���g�x���H_]ԣj�X�^��p��1������;�w��ׇx	��/��3c��(�Y��U�
D�>���,���÷�(\C��џ/uy��yM�t����ӯU��ѿwW	�p�~��|2O�-3�n��%x��F���ʢ�wd�`w�'ϒۛZk�rw��<4�g�Du����s%�" nk��"e��l�ؖEp��>�NVߌ�8�1n.�F��HTu�z�9��>����h7����<o�v�,)-��ȁ��D��w�z-�zO�&�Vl?x4sN�^7���m_���ȟ��>�^���ć�Z��}���=�G$ŻEƿDV
����J�]%O��^�=?+�1m�Y�o���j6/Q#Rj���P�ë��3^zN��K|i�d��Av�`߶�{�oK���g���F?H�����7�FV?l���C��V�����V
�d����W^��j����W���μ�S�B��W���vߪ�FS\}���z�7�c��E��(���3�v��O��R��4a9���H�8��f+A�%/��M�/��W���ˤ�̘�[4+�*�*������ػxq��0!�V��ځ��[��Ī�>Q �uw<���ֽ��ó������;����p2� �W�*�}ǘ�;Z���.�к��K�j̻��1q;�i,�z�i���W���ϰ�n�;�uz�
��np�s�r���:v�^��v����0}�?I��g-q�c|���R�<rϠWе��g�族�دN��y�o(U�j0�&t/�7DbR�Ҍ�ʩ�/�t��y���e%Iѿ��πV5߁�n���ϫ��T�Q��C��1U��F�ϻo2��1w��<}��O��c >S>F���A���
��/�����T�xzy9�u��z����b,��1.?��L^�]���i$n#���t!�����v9�7�۹-���K�8�硪!u�[���qd���%Q�p&�C�2�Y.�|{WN:��~��=ݸR[���*�G�#�{�${J�����^_�����Ԗ7>���,�%f{2o]y�;(�f�f�3�~Wq���r���;��'J���g��-̂�B�F���{��O8^y%+�.|���`0,Z�p�Rz�1��޿3���o�{�����Q~�ﯱ%��Ii�Ǐ�U$g�Q%�4.����3��*#zW��G��ώG�wĻ���T����W��U(�֓ズ�vu�#���R��*&�
0#���_���w�Z�#W�yJ˭}�i�r�r��۹������V�`��,gCKXw� �!)q�YL\�VWn�+GN���U�]������x���P=]wo7{z��t?K����f��/��n�[5�,{�N���w!ݏD�w�;���V��U�������{>��*���,��C�c���{�6�~1�u�2�Gӝ�tv�VMjֲ�sqi�v=:�7��鿽�����L:���������Ճ��{�ތ�>
���1r�q�9�ޙ���Gp��}��3�.~�ҵ�����]xOd{ݖ�%{�x��/îW� �t�g��翐���6\��|���#z}�q�j��潦�N��w�ૈ���xߍ�8TH�>��ˏVg�O��*w�3�P���9'F��x������,��z��V��zhfɰ&gE�N�=�W������N�������e@�ȱVMi�4�(�`r�hJ�lsJl�/WΪ}�����v�uxo~�B�V���R��=P���R7���uP�q�+�j�F�o/ΫV,������RӞ��1��C�dK�B�ڑ�<I�B�L9�yg+�����v��v��l�;�x;��9�����\?)�����y �.��O�_}��;�i�H�U%ܡ���dS�iuyo9+�kthV�t��ֱ�'�������rZ��I�� ����]*��]2�E�]q���]�&)��''c�����R�l�]�Z�]���umڭ�6��EfBi�4��gZ���e��$�ct�G%���%$�ν����a�6(t�j�j��u��eu����m�d�)$WI^̡�k9�\a�_0�Eka���+#�Q�['�mc���h�����t Z��_e�nA�(k��֜���q�d�Lk �ǩ���CHͳ�ìX��*'�jw�����y�;�6�Ů��\�@"���������#��^�k�㮁�׬�����;:�����_jy�f"L��e�wώ�f+;$�/�����`��3N�p&����6͖p�onҹ
U���rpU��������D,����*�v�-��t�<�gR��n���s�w�ǆ����i!��\q4J%:�+BN�ܨ��e���{:�gP��k�2�y�'���vmw=�X�5����B�ڰ�������i��m�:Yo�.���U��O�
�6�*24*Ç�I�Ǖ2�
T�"���{��Ew\uϡ�i��hm����pa��w����tg+�V�w�"��N�إZ�C��XQ�w-7��4�Y9�Yk��$�;naYJ]�77�-�;bw!��,�!e=�� �N�s
�pb� �}�ri�\ӝ�"v'U�ofݵS������{D�b�����OK�����}�o����z	u��Ҽ�WzJP�yMgZ���|B�����wnu�Y#�r�MD�YbN)��f�(4��.�v�h&�k�V�d�������+1u��b�Cx��8��^�Ŧ��wAә]��Z�W!۲N:��G����(e`z��Ev!�=��uهK�-֩�R�Ur�Τ��8��N��U�CFs)�1�X�
��b�wI�);�3��}S!<������AӽpΫ"ю�Ӳ&�ƪ`�B&V��� #gy�[:��$ިG�.X��w����݀���ӝ�;�$\(��7�����0nKt]&�d+�2cʶ^a�ć5vc{K�U#��������-z��&ㇸ��VR��D�Fk��-�O���cl�*f�O�I�.������3LH�tn'{�����a��m���4��lO���i�iV KL�.i�2�^��ӱ�wEd�y#MN��\5��M����q����y������yAVS��=�5{����s�	u��XV��K����+�X�����վ��1L��N��x�!p��[�Wm�g��m]{OK�	��y�_3�r�B��/�d9e��}�Z��,q=VW'ҷ��(^9oA�!��6��Y�.�sD��v�rwm����<�5�c�;Gu�YU�5�9#��r����w��^=�6���>�q�<4w!u8�0:���l�8D�����.6zL�R[��8�V���8��۰�Q]7�d���+⨾�;�BT�03DRi���hQ&14�E#�0Đ�I�h*�	�2�@�ю�fd��R%(��d�&'.F2F2A�lI��iJ� �F�l�� �2BX�D�A��H��Y0��6#0��NnA�#�@
i$��QA"I&L��L�CD �4�HIA�1(�c#1H@!��D)��*�"d��+�b10�!��d�dRA�@i� ��D(�Ԃ$6 (#�sf&�(�D��,d�����L$Кw]��� fJ4b�$"��(�I�L�����|(T T{,MOy�[�][�ݫ����n��3�wM6�w+��E�fS�q�p��,=�q���%�xLx��l�������rJ���]O��4+Zw�9�'���t��j�}�V���Yy"�ϝni�ݑy伦o�ǀw�(	�(�g��~9��ԅ_�ֆ������_���L�/4�^�C!����2Op@���H�W����z�C#��lx�W��utD�J{.���k���d�{����N�%�D@n�]FC���F�����S/�ju�=^���1�nr�%�>����r���&���p���ә�ʰd6o�=$L��Q����b�*�.�;�~̯^[�]�&Ͼ��*9�W���xİ�C5�T;�B�O
3/�����-��[����f���u�z�D%>�m{n=�?;�7�_��q�z��123c��2iL2�g��H�����Ѽ��v3aIXpz6���Y����^\<�O�|c5�+�o=>�z�޽��}����s��.Q7|yEy�=/6,K`N7d�Y���N�V��ަ=y�x<1��ddk����:���.+o6�Z�������X��^T�Љ�����+�D��sau�E��z�;�\x��Q����=�����׈����%���E�g��q�䓥�UǾ{�p�e}}amW��71��7�6�[|өf�'���=&ip��U�N+��9��n�.�'V�k!If��:��+V��f7b"H�8w<�,VVʃ�P���	�Zݜ�\�&~`��������48UOL�=Yc.�wn��P|��YU�I~%5ɫ��d砙+]����^���VEϽKޓ�����pK�H-S�z���(m�2�ў�^�:���N�ٷ��N5`�4z�@\|z}��|Kg�^�����y^W����ꝓ����OM;���(|�g��k�Y�a�L��S)L__�K�ޚ�x������ޗⲼ�<��F����/�S������w���ɛ>���z��AH�\T�B��Q�j�U�z�8yK�Υ�E�`�oU��{�q��o3�z6��$�P�UA���ڜ��Q>��o8P��?^�����ס�i;7t3i����W���e�Ύ�����߯��'ƙ9Q�p'��q /|�CGmq�9�B��U����U��r��^�����Nב�z��n3ޢ;�,N��d��@�I�p6"��I��>^���uu���Y�3����>B���[g>������z���|�zs�i̒�B�l����&bjl�/G�V���=ޭu-�����
��m_��������>Ȇk@u�~$x��{���ZM�)�u�E�1���6�@�th�Y�:uD�=Gr�J*9մ\�ĝ���*(��
��gISv�6+������ۺ����x]�t⫂̖��y�TB{u �� ά��[�Y���W)\y��ŵ׷]}kd���X�pή��V���6b}܎u�;>31�:ldO��h^_�q����k�G���Y�o����ʮ�$fz}�kVN�EǢ�&�ǉ����TK[z26�{�f�1�UXc�O�rl`>�ثob�V���չ��3��=o٢��{jA���d���a]z�M¹||�9_�y��&lyV;���_W�b���k�=Ωq�zG���U����j��^T���N���ӻP���Ց��9�Unw��9�̟Z&ϣ�_��gZ��u^�q���9�^�d_���t�:�^*�%Ҽ�f�K�1oҘ��}ή�������l�p���+�g�g�Y9�9������,�^�F�M�΃�W�uw�o�7%��Yؔ�*8�=艔2	����Q�t<� ���~�n�����?����=��82��H�,>�1�{jx�d��|2�x�u3�o��e����,cآf7k�r��g=�r��]�Þ���k ��k&Y����0�k�*����H�u�xS�x��:��`�]7I�����9��͏G�%x�H�����q�{H<�d�X�J�0�I�we��G�l���S�ؔ�ZȜ��y[t����(R�x��8�jM�X�7�]Cyέ��ݵڳ�N�
�K]�j�q�N������lۗ
jR�N�wN�|ؠy���J�1�׽J�ݨr3�>}tY�L�u�w�gJa�:�u(^���.N�ƽV�����N���y�o�i_{UHۇ�@�[ R���(E�Q��i��5�#}���>�|ʿ�Տ"�ʢ�ޯZG���;��*���q�f��,��n�t�+�\^︻��<�L�b�p7 �3!h��H,�׭��޿3���&��\O]kd�Bx���e條����铦�U$5c�����s�;���;|���m_�>T|ro!d\���B������'|�F��j�j�'�L����1R��F�定ĩ�_�N��2o R����>;�=2V��.�W���zT��xπ�d3q�?]H8����!��/�p�ܯ���K3�eL�7ٳ��o�p��m������я������q�C3C�s ��;�Ҏ��wm`V��0�]φM���ݯ�����s�Z;��Ϋ�}߮����/��ׄ�G��b�G�3��O�E{/���}^��=�Wr��~��=:�Ք��+����/����މs^�ߢ���w��߫8�_��3�~�W惊�u��vv�e�CgC������ү���{�q���x��o���~����|h���r8�m�`z�A���i�^b}���U�v�i=b���vKc�n�~���>�:v!r�"_,�:��B���q:)����R;*`"�S�k���ۚ�%ϥڮ���3��7�].�v�ȍ+����u6wk3�E]�x��g_Mb�I7�y���{7�q���/�����Fa�	�,\Ed֑.@��L
Z�=~������*ܛǝܯwF��}鲲+Ԇ���/V���R�0���u�z��݀�m'�ƽ�f����Y�cC�}�#�W�;^��z��Y���.!��9-/�,P�|�'���6o�W4xRl��ũ%*����r�]�y�^��'����\?)��^R@8K���$�ߦ����&�f�g���p�yTm�Ϝ�b˩f�۫ӯiQ�'����I��j�z�>���Us�~<�]��勫o�:��G����P; �xw�_������W��z�;���+s{��j�ݐ�m�&�N�M�#��L{Ie@�����I�+�s��Rz�팃���{Ko�w�{��������.&��z����bX%����|'�����7E���5��É��Mn��u���X�M_�z}H�g���7�z��g�&���e_��l�$d��Q��I�s.�x^ug��o�f��������LTrj�%D{ޤ�<k��C5�S�`�B�O
3/��kn�ĕ��>������v���tvv3��^��譺f%w��c�KZ{6�׿z�=������T�>��'�;>���]�2S��)0�D�]<7�ڹՓ��Z�#+\�H�ŭyi�Z%r�m2֤D4'ˇU�/�ޖ��ݛ��x�n(Ĵ�`�Oz�U�]r=G�q�k�q��w&���2o�{�{�q>ْ�|y�V)c�yP�I��A�a�@S�\T�:6�W�(ާŪ��П���k�W��Fz} �7�����s#*�33в��e�6}>%Pɏ+����T�N��[�'�7��^u���q}/e/ѵ��N��$��'XΜjh�o�E�w�8n4�wA��9���J4�A���
o>}��q���ҺVV��w�z%W^��?V���X�2�ڸ<qX���N`5�a�ʼ�K�[�P�;�U�9]�k�����@�x �ʈ�^��IدTo���^�Aj���|J�/���;�Fv���w,�����L�\�g ������^>�~�~/"��7�ϱ��T�{��x_3c׉#5�W�+�<	�$�Lo[�.nz�<�ޯq���>�~<��<��4�@�����r��T�e�x�2����z�2��ȱqR�뺔mZ�k޿�=Lmv�y;�����3��qƺ��lφfHܠ�������bKa��.
�HQ���!e�O��o8PWK�(N���	ّʐK�~V���Ʒ���-TMf�f����}a*�ܔ�[��8p�mN�S�ZN�[��j�ח~�D_D�1��X4۱\��}�v�1��p��W�]�>��.t�\�-�Wͻ����ٝ:��m��Mm 8*�r��Y�{�z����W���7��`�>,��8��s�W��GeOخ�%@�}���KZ����l�~��ޯ,C!�ב�z��o�������.WȀ�>�=�9>T�{����չ����a�[�cRt�d�Ͻ=Z�޾�9�5d��<��>�Q�{������"by�%���
�[�c_�ڿI�z|���L��C5�Z���5F�8����$z:�����ǝ�X�x����.5��>-zH��w&~�$�U�Z��w�y�ky2=p)z�بs�2M#�z�L>�>��ތ�u�5�oSm]�c���\�2cn\��f����{��3�~� yz�P߻�Rt��C&_�wL+�V�T_s��e��[��y����ݞ��m]h��u^��<e���~{V:�d^F�'j����P߻k�۱K�Թ���kF��G�jR'NGt�ε~꽤�>�-z�
�����s�r���Պ5L��ӭ���z{�ק�ӣ�"��M��d��g�+�[�q�x�U9����F�^�F���l�㙹�}C�r�����1٘'Ү�v��
�)M��k�U����� ꂆ˓�I���\E�:�ۧz���T�jy����x��q]����Ν;(*�hs�����v����UͩM�\}6���2&`��ά��Ȫ-M� �qg:�:��j=��e��rǢ<��ۙC(L�W>���:S�vX
ƻ�6�/>�����0�[�^�
��ɜ���'|�^���q|JW�2����ϑ��tx:h+�:`�V~=	���x���թv��ы�#ޯRX]j1p�Գqg��3ƌ�b�*e#u�xSQ�>Q^��r�]�GWn]��~z�g�O�w>��Q��޶=�>�����Y��x��Á'ʡ�>�:����P�y��N\ש�˸��~늸t��W��o�q����m�]�z��� S��{^�u����/�h.l�}kj�G>�uG���H�s�iQ�Iү�둷������uS+�3�KݒZ�P(��x��)��`�3!h�ϕ ���0�ӽ~g���ۺj'�2��K��g��'���H�#�X�A��r��|9��#m%l0o��B�umk�度����D��5�v�%�������b�_W��e�]5�S��=12|�5J_��S�Ň<E|ӻ�����ǌ��|�Ɠ�+W%�
sؤꀻ��Q�߯׸	Hkw6������m?U�j�����-��bC�螭'
{�#ý�]�Ov�@^ө�O�����T�D_�p�����JgU���ŝ���g�I�]Ӄ	G���^�Z���7�.w�j:u��Q�;�JLW�8��^��r���{�z���߆?:�8� zW�~���������q̼*���/3�Sr����>����]�h��G)|s��~���~�=&��]xOd{ݖ-l�^E:X��[�yt��z���s�ƝՔ�����O��~7�j��.k�c�Wx�������ݕ�V7]w�:�]?O����fp�����̱��·T�iW�w>�����,��K��r����x��O{��}�o�Uc{�j0�o*t�,��3* O�bpΝ4�,L
c���"a��	���u{/WL��{k��z�+)������mO���R�0���+�H�k�Mt8Y^͜��z����{2^����q�{������R��mmH���$���_�k�C��+<�>���9�d��"��7�*��ϝ�8�O���I�����_��^%��%�=��y��vw۽��>`��,		�+��W��]K7�X�����yI�|s�'ǯ�j�|��H�檘/Ft`�sݚ=L������ 9i�?@R��R</�t�}^�)z�hh�����B�O��+c��H���M��b��
[e �����i� M�T�f@�ԭ���bu�d��=--�5Q:�YMx5A��B2��<<�ھ=��E�������-���Iʵ���f>� I�^�e��-.w�>�\Uy�>�Ƙ�XS����홹Ԗ�j˿7��\N�;��$�P��ʌ�����H�
�����۸ҽ� *��2���{3KMw�z�Z�Ը��z��W�%�Y@@m@�&&W�����5j��ԛw8�3�=����4���tÏO�������z���z�j!��eX27����T�������n(��|�Q�;W�Ŧ&5>�I�{ޤ�<k��C5�W��P����7Wnۿv�c�rw`�D3c��Z*�˯x��R��^�c�c��d߽�����Ή<�g�9uf��������>��e�D�aN]JӢ��_�oKҡ�ˇ�����}��^�]W�AMv�g��(;�o�����>�8o���Q�ѵ��T�N��n��ޖ={Uc�&{ѻ1��Rkw��^��r�0Wo�ͺ��w��[��C]�N���ݳ0�_	�0�'�z ӭp^W��2e�6n��=��^��Z}��ԇ��}^�!��V}άo�ԅ��H˅,�ۃ0��*���/�(���n��ױ.z:����\Od� +�ZՑq+Խ�;��y���h^��:��xEUO�h�;��
&)����e�=��Gt��J���թ,�wD�fw'D����f���0��cp�� R���ֺG+����.�5ϩS��
sA����I2U0��f�7��,���>:f��o^9�m�W���"���D���mj�Ҫv�\�+�Ѓ��&�㕚{3�R���R} n9lx:��ю��'���e]1����q�ř�����s�/�lk"(�j�4�_7s��I\��k3�#ܱ{u���J�v�<�rP�z�ݝ5g7�#�E`�"w�c}f�B��u��j{x��?xd�ϙ��[K!���O���WR��/�����B���*�o���V�i*k�]I����z���F���,,/ui����B��W5u�/��xT�S�6��a2/�q��׷zQ�+]��tW-��	��e���A.��݂)/'#vz�P�!v�����ݺ]���k��N� .����Z�Ő�!��. ),	{���f�pBk1gL��]�KI*66����'B���%�HL�G?��k�)1Z��<�G]�%��fJZ%C����Sfrd�un m\f�pTX� @���e`��t��{��Y�gF��g
X&@��p�ˤ��ꦛ����N���KnjA��L���J�ղuh�n����w -����rǂ��J���\��\��$�ө���L��4\%jt���7��&c���3P��3;���r��u1Q�u��|� ��r��s�K%�)"��[lpMNw 9ʊ�J՘ C�I��{�)�=W��Ƕ��{L[ulJ)w�/^��Y
�oVGҹ֌w���m���5Ү@�́�r]9#���ͱ:�;�;�Û��n����`3V�b�w:�����̌�em��s2q�Mռ_Q��ǚn�-�s�Z�w9�e�M�l�mV��Ne:�{{�E�C`\�2dY]V]G�A����Wu�Fآ���퉃��[�
��S9j��]$���:|���F�4�������Z��e�ѶV����q����F��A�ޢ������vAc����Nużz��]��؆�P��57.��8�VWM�]�W��m�r��Z��]u����'�!�=Ϩu+�1Y��.�c��ZS�
Z���ӓ�o�uΦI�]A�]ι9�IH���T��3���m�P9��M�K�ȸ.bi���w��wݽi�j����.S�8SG��̚��pu\�&�)R|[��}�u��].w�1�S�o}f����wm�t��#��3��%bɍ��.�]3����Y=�@b�J��X坫39q,鬭�ɞE��z��s��z怜660�X�PWϫ���;�k�V�C���,�,�D���8,�3�1Ʋ�\�&��^YIƕ<�y�S��� ےr�	�ix��Y����]]������`)�W�t����AԿ?+�-�s%���2Lg������8�&R��
,h��e��`̤�b�<�E�wlƹr,k�f�jB2i!6��j1AIJf@L�3"ى�5���I�]wO:wRHG�t��PD���&�t��wx�
"4���fC���U��H1�p�ѹ�wy�$� �k�����ΜFCe���nE�k�r��+��x�DIE�ӝ�HI;��ȈĎw��)H�B��S���ݻw[�Gc"Bb�q9�"�x�
+��DF)y�!y܇�v�k����c���Dŗuvx��#Di�:m�ۜ D�B4Q����ٖ�g_�ܷ�N��5����Ȋ�l�2up�&�3�B� 8@
��
1Ƥ�9��;��R�=_wL����Ʒ������t������|z}��x�nW��~��p�^}^W����{�x��a�����k�2xz�$�J><=Tϔ�S�.zz�<�ޯq���9�K�S���>97���Z׍����u��,3���A���`"��J�.#��Q�j�U�z�8Y��]G���={G/;yu��Fz!�(����d[�φIf�g�*��AH�G�ڜ��Q>�D�yG;g���9�wm��M^������*:{�(N��C�%��a@��������Xv��;k9�WG��g����ʢ���g'��z��o������SP�K� ˹��g��o^ϻB����`7
E��&5�~��G�w��|vp��|���<���Qo'3�Rk-o�Q�N�D*���D�>t�]K�x��m�����ȟ�L��U����[�]��;�WKw����M"G���OM����Sc%�xп��K�d%O���#��?+�1~��:rg+�hgos���;�ɭ���5��2J��0��O��K[z3�^�Y�Lw����;}8v�Ѯg zXc�K��g8Q�|~Inˡ�;a?�n^����{ML(�:�,!�)�݈H�W.�Y��Oj�f��0o���K]j��\�
�Fy�;aK��FZuٙ�gr.u�:�%�vC��(��u�7;�����ɧܴq�w"aFv�K3�w�����܌��zg�,�^�.;�Rt��Q&X��
��V��~�[���˳�,�5s}�L��4����y~�W��P�S�`�u�ؘu�+��8���p���L��j���������r6j^��q���ε~��	�n�;�v����}����I͟ "Yjp��m�*���ӣ����ᢧG�&t�����l-��fW��u���:���k�J�}W��`��*��Px}�}�y3�̜9�>�YS�:�R0�:1ׁ�t�|	�����j����rU��z���լ�vL��{�B�3ŉ'��[����AFҽ���i�n+����<��Cs��~++ԇ�Au���{��!&mQU�ŕ���]�̄k\6���۳������T��
�j�G�|;��F{���}�G�{�Ǹ����x2K,q%i�p:�Ǹ4s��\��Kv�*��e��e�O��;}qW��NG��9���7�R6�~���@8K>����z�∾�����> ;�D�yJ^)l�h��TW���H�9��\}�p����o	W�B��y���B�Mzӣc��!gŚX���fA�[�w��a�;a����WE���M����{��[��Y/>��^��\��:4K��l���� �{��]�O��xAuk�����뀮'6���G��E7(�;7���f���3:�;˄��	"��c�[�ٟ��A�_8!Q2nx��d#-��|��ٌ�N���qW�)rܧ��Vv�����Y>�����z��9��*���Q%yM�=���9yf���	������/uJ��8z�g�"=3�%�F���_�'_q^FXJ���0ӥ��3yk�uxD���˻��J���wݞ�~��d ���sn�O�<g�w�!����.AE�����>ʉ�����{���wn���zݟz���oT{K�e1\����q�_������� ��=�.}>��b(����o���|}8�N�M�����؎R��U�>o�|r5�����]xOd{ݖ<�2A�,��w���ss9��䰬l���W�ں|O��~7֮=�.k�c�Wx�Ǽ!�_���:��[�������Q����Nlχꁳ���:��N/�S�|�<]>�����g{}����{���QY�c{�Z�(�ʝ7�wn���X�3�M:�[�����r�ڷ�}\�+���@��s�}N�+)���e���ş������T??&�%y�t����7o$�ؾ|��WQ�+S��%�=J�m�z�+����0�Lm�Z�6^���>����	t�5�ד� qr�!�2�DS��n�_�Sգ�(dz�k����/X�\��KOve��{�/v��[��w�i^�Fv���!�v��)Uw���5h�=?�����C������ҽ����������%�mmH닞$�ʾ^���W���ŷw���[g�y��*�n��o�p%�|����{N{���r=��g�|8����i��[S��=S�M{��I�@O�*�I-χB˩eӚ�;��)>/����W�.vVl��m׵��z6����@85� X�`��K�_G�ԅ\z�hh>���g���ݾJ�׌�<��O}Q9�f%��A���-��d�)̄e���~ˣ}^ ��Z$ד��:�V��FC����:�5G�K��z�Z�=��ܝr���� �$��ܝ����o3���u��K,���G�C��dh�o������>ȏ��n=�Wq��Ĳ}2����Z������#��m!���<p߈�D��h����uǙ��b��5~��zP>� ��k@�t��}/�K��FTp:�rxiG���̦B6�pWe׼z�"������w'~&J����m�>Y��u71;j[�Z�tz��Olɨ�L"����=8=%i��o�³z���.'�0��H7Y��ꏎ,p�MT�;/_btN]"r��G�a9�G=�q1:oQ���*|�G��Fv@�z�l�T;ꏨλ����;u���طmj<�[ݵ�_wH�}R��z IݕƗE�Y����ոx���^�]w�r٧']����əMJ<.��c�P�@GL�]���z�u���^��\?^ٸ��3����C&�Z�S�:.��{#z��|T3�>�r�s�7x8y�]��������X*�ע�ü��q���pf��wY^��cW��v=d�n|��*�̚�S z"����V�ֳʧ�C�T��6�j��-��#ԙΣPN/w�ý�|�*�}��W5>d������"���^����{��S���p�F��=tncP��Cוf�Wt�zϴ�;�+ڏJ�Gc�\3�A��c}^&�^>����y�y\o
�}�~�W�Z��3�Aa�X��;'��I'�"g��O�3�1q��K�ޚ@�W��mie��#�]}��\�*�a�}]�	a�j6��,�_I��b�,]J�:�eV��<��7��1;�I�:3{Ә�D�,g��|z��q�Ϡ�����IZe� �H-��//.{�do�ܯ2���W�o��g��S���^��+cʎ�����߯���|i��A�p/�������Wv$tǷ�n��{{;<���^!1�T>�O����y߽�C��zH�L�.���z������2,օ��ĵ^@���C�S���E�j�7H���Q6��@;^��o V�u�M�3��ew`N���!tc�xÖ@�R2�8��>X����nk��zN�f�k`$���f���b.c�}l�`�5�iT�==��|���={ױ���> s���z��}��5�Lo}��9��>����h>��@�'��v��o'%=:/�^�W��lwJ�����F��HT��lG^7��*:�~��"|s:�����k{y:�:���M�E|�\���^�
�TK��q��\k>J�k�G�;&�w��^��~ܝ�I�Ӽ�&=�iY�?O�w��j68�̒�'xd���0Z�����kԏ�I��ookV���z]�C>~�܋�������^�6;�Rt��C&X��8(a1�Pݯ��G�.���{U���?�ϙky[/:��1��q��2��`鿛ڱ}yR2�e�E��2�>��NOd�vq&;���1�az��"K�p�/��Z��U�'!���9^���}��
��I+p'�ڇ�U��M�_J�it���LTE�	o��*����;�g�族���<ڭ��/�����3@�z�F��L�^��n&X�<��>��K��=e��]x.uk���z�B�����,���E�M�>U����ƭ��v|JVe��g�O���tw�|n���ڑ�%5�N��v���VQ[̒keg���3�u��묃���XS���}����Ő	�u�= �U[)o7�
�����@�7k�r�p�uhe�n>WCf�*���-��6	�}J�腩�����g-���٧�*d���(�/��{^=X���V}�C�9�a�L���'���K
�G��=�*ww��W4ޟC��+���e�q��`Q���I���l{�y(8�YCI<�YUW��<��ϯ%B���>UqF|ϱe�K.�TW|�ߴ���:��P�q�U#n��=Kca*��Q�9�+��W^�'���^�H�H`Cs�zl��A���Q^�z�8�w�q�zN��q��]��;�wܖ���E�3�L��D(!H�끿�~(b��*Ad:��`�~�G���%���u�<�}|}g��������ʒCjQ���4/�s�;���9������e���[ٻ��~"�Ӵ<3�O�������.�����u�yD�~�,�^��*��Y2�u �\��{N�h��O�l׼�_��<�T�m׉�����7C�\�JY=_!����m�N��{:3�I�A�;�ѷ<�VF�Ǹ�^���~uro�~�=7��~����ʐU��y��f�^yw�JT=D��di��Na荹||�"���ˆߪ�����3�^�Z���k���+s�N�	�f�qI������ڷ����+�2�0y�gn��w)�0�v��57,�Hs�8L����<w�+����/̮����T�C���S�VŘ����#t�_�m�̮�'y��:\T�:u4˓��]e���w����v�f_k֓�9m��ɛ���|rXWgC���WO����o:�ǲ%�{L��33a�g�uS���̝�f������g�<m��p�����>�N��9GE��_����v3���x]NwU�c�=���wЇ�SX�دV���z�ogz������B,�ۃ0�����R�rW�_�/߲e��ou�~g���T=��EĮv��t�R����H^���qgĤ;&�\A�E����l�O�e�^�f��y�� o�d\>��Om���������C�����I�~�����u2J$j>2��Q�#q�>�,��wz��=�|}���9�yׂ�I���`W������
����C����yL<��[�u2�C�V*�~��O�җi�tr��>I���~���}[��f�p@�Pe�!J�H��T���!V�|&�A��p��;�y�|���_�؏):UǷ����aŒʅU@��I�)ɞr`��Js��ٻ�K����u�!���3�N��vǽK���޸<}>��fK4���|'��US��'��j�;�Yfk޼�n��(�(�6�H�ke�d������x�(��M"K���ڮ�M��؊��M�ή�J�l�7�q��G��C,=�yPB���Z���Da(_{|��nLݛ�̀/$c�-{�S�RdZ�m�:�x�sJd��/���ap�_q����pߝ���R'�3���{ޮ��뉧3锰6N�@l�������g��D��F�5��6&7�5~�q�z�>ϼk��3Z���4L�������O�b�3<����R��U����9�_����j����%,>�K���c̥W������x��>ٓJc�M�:ǧ�"�i�qo�³��|o�.vnv\_>�V�ٙ��m�-0�D�>�O���(�i�7�Ī0������iЩ����Xl6��������H�C�1z����;���@���m�p��(�w�B���:����ȩ+����F�o��*@�ux �Z��]z���YYάo�}Hm\ȼ�K'vs��y�Y�\���V�*�qYU�I�J�� ;QW�{�v�Q�S�{θ,^�C�1;�Χ{�7���5��<��0�vc��Wە���*�iJgr�BeM]�UKYV���	��ߣ�c�d�$�%(<�S>S��K�}��w������s�U9�^���}���;0B�+�\��'I��OV���-�u�t!L����ɰ���ԐY%�{y:��c.E���R�0;�y,���u��naQ�:�:��Rkˬ�*�b�%5fU�����2�Ӿ/� F�ʂÊ���&��� �]t�rԻsG�;��5-��^wY�u��2��7}$�,	�|�R����Q�����z}Y������.��4����1�w���dAu�1�%��x��>2��"B��(3�Q�&�=�G.kԲ}.�}j��(9~��>G�Tt��P�<�~��Y>;����TtE��^�W`�.6��^�&�	�>�F��o��*�^X�9>GTG�Hq7��ޙbkkc��ztw��d�Q�*}�3�"�[���؄�E>B����|Nq���OV�>�����ZeJ�v?�to��t�3Q�|+�S���=$�B���F�+�>B��U�9�|EI���Lq'?<������ϡ��'��Z}m�+�r��30�
lg��h^_�q��*||��x���^n<7�+�ӻ���d����C5�O��(2z,���1Q�ށ}�)�w��c7j�S����-5�z�:ڻ��~������n#ޟ z׳E��mH5�O�T2a�x�B�;������YF7�^��j�qkc��p�������5������t�{��beUb���n6�e]L?�l+u(ℽ�*���skn�:��L1�F2oT����/�ds��4Q��%4T�q|bWO�@�"�ln ��-�c�pok.�s�r�Mͥ���3h��q�qSB�J�ҔZGu���f%bT���z��}DI��X���7n�j9�:�v��8 ]MΝ��y>v��䦄�N5�I݃90�Sl�v�{��'t�CUuzh�6���
ܚ�e�H�Md�������y�n��}�e�J����1by�EH� �S�)�\�,����e�m:�^�c���.�ж��H��r���WDٶ�ƗS.ue����0��{}��wIr����#��'[�[p���+���I�c.����lAR8���z�fJ�\+��^V'p����.8�p�OH�_6k j��Z۵��n�Y�	i���K,���=��tZL�j�mm��}������>��P��k�9u)���KO��A��6�,\��4���-.U*97/^��l&�pQD�ϐ��v[����K�<��:v�sˡ��S}������:���xԹQI��4�bv�]7���9��`��0\9�s��܈�n����u�te���`�#��]V2�pQ$`��l�3p�]+51[��D�*J����e]2��N�+4�\\���Hn�����|�1o��J�Bz���5c���&Ss�˶�Z�S�&�Xa�=��Ъǣ>�Ü���wE�㥮ڴi,6�K<��$���0�@���M"����C(�j*7B����3ml����=�����w��K"�M݊b�]��^fGi"�8�q=sn�۱��	��˭t*2Nw[|R�Fu�fm-�1���`#��9��ǰB0�P�(����C��RP�,N�=�ͼv�ƕvB�|T��WsRouj<�L�qV������"�����Wn�!�	=�Yo��oP`'�z�'����E��w�O�*Y�h�;�*�gR�Z�n��+�c�cu�A�\����iM��4�/��\�sP��z���,)hn�7\����p���1������y��彊�}HلLԍ�Qw*����!D���Ç�m�JsS]p�Vp�UKB��@;�|�F�.J�7�l��n��C�Y\%��g�+�r����/a��\�Gg�`cK�d)�xx!������/�#m��f�[��]�Z�H�g�ou�j�{s(]^���ͤ.�[Ր>M ������Y�RE��_T�w��W�MD�Է�@1��Ҩo�n�[�Œ��>�@����z��}[*�3��7��U5��l�te=U�:�n���|A��8m;�����7���u8�;9���U���Uٷf�A&�*YSC�y(�A����j����� ��AE+��ҫDmd�Oha�[(�7���ҞC|;�~�;�b\��E
@PH@�o�ӻF��@�W`E��h���W(��F�wwa�]���)[�:�ܺJRJDFut�GwH�Nk�RP�DR�rb��Ik��ۛ�,ns��L���QLgu�H�2	#wuy�h����!(�wb:r�0��",Y$Ӻ�]ݹ�H�1]+�E�҅D2y۫λ�I�&�w\�E3lʋ��'K�sW2c�q$9�3H.[���8D�Xwt�؈]��d;�y牼�!)(�L�㻮낓�.��Fs�nk�H)�]r�����+�iB� ׇhEӻ�]n���b�	�tB���\:�Dp�[�aN��R�ɓ���=������5�# gr�=Qw�QT�.R������F��GNKDI��.��y֯�"%�{Iϛ���(b�.�Շi�b�-�{]�k�|�/N�@��V�WR>Vz�TF)P����e���Wȗ4�|I�Y;��l���n�j\VK�7�q�>^�F��y3��^��n&Xʈ<����4�yH��Hݻ�	��g`��*ڮW�}3�
�\P>�S�R�FoC��1jڞ7����c(���ϑ�c��+�\�M��tywnuJ�
h+��z�"�Z1��O�g��C�>��Q����f��Ğ�3ǨOzXyow�=s����2q�$�G]��x��<�����p�x�G���_�l{�G���y��,�ώ�
j=^�w����2M�1�B�2�R���v���N��#�O���@���R4��AźtN��������z�}Q� r���$7^�ʵ�a����*�^��|�w�q��$peU�=�97^�����7��\�u5�[diAUD����P��h��H,}U.IAfE>��홧���ǜ�Z��;��{޸��Uxȯ��f�T�ݎ�&J�N{�L]2����O��L��h�Q��t���0q����ݽ]��Ŷ�C�{حc�;�ٗF��Nu���:B�]b&�d��ݖ�4�����=�ziqr
����[S�:��� �:hi�S��V[|���/[=݇�O���S��`�w{xα*�P/�_v-�/�-n���~gޟ+>9��/#ƣ`S�Q('��^��c��Z!�Żx��Q����>��.�JX��vG�����[n�O��|y��_���,���ע=�G��T��ͭ�(�s6sQl�{z��k�~ήM�?P����q�|������ʖ읩���hh^����U|�gg�+պo�||��)|o��ˆߪ��~�='+��ro�{uV�_��dP�`��G.�϶g.:|
5'�\|6t;���ۅt��;����Tz���|#OIy�����O��͸�e�����՚}�l�G�gI���6t;��:,ү���K��K�W�9�U���z�l� �5�!��R�x��o����ow����o*t�B,�ۃ0�O�`W�?T�r���uחcִ+��khѳ�:!k�����2�3��ip�Ԇ���C��O�|2)�!C�
N���Mq���6A��*�o��x:�x<�Y�{���c�+և�/)y�1>�{����O\��}#�s�J5��f�ʨ���7r�K6����ޯi�t�n}�V�%����ć���Q����~̧��}��:κ����������T��9E ��or#2�<x�A�v�D]7/��x ���ö��f��q�����4����pn�%�jV�a�Ƨ[�Y�,�!�zo+����;���.�4�X�Q�Ώխ�rN6pw�_���ǰ'��$�̰$yT;����!eԳq�X��{KT����g�3�7|��{�fo8Ͼ�\{U��>�������~2��P7 �xw�_��g��^$��˿{��[���N�h�~�[G|��^�TNw޻�a�@�,҂*� z~��9pY��=�� J���������CϽHp��R��_�{��M��O�^���d�P���zH�wM���o�/	�Mz���Z/r!����8_�����"}��:<O���;�뉌7��
s�T�^z�h�.��)�yJ�E�?��F��/���\/���M_��{ޤ�Ƽ �?Jͯ{��ĉA�m7�VΏXK���t~����K��x�~:̪���k�q�~wrr�uT�1���o���g'ͪ��x���l�FR,������������;�����k{�X�{;sm��_�i���}�I��=>�z�޽�q��g��L5p6�9>Ӂ̩��f��>�3��Mo����u�����O�V
��^��*p�d�l��֬�9�1?wEF���������q�2�����%��{/��b�w�X���I����Ṵ&�6�=v��l:o�k���;)�GR2�)d�yK2�	���T!̷Yq��N�R�-��8��],���"oe�.��)�;-o��?՟�q�N��]lQ{�~ϫ��YY�����ԅ�m�Hʌ�
&��W�|�f�yLӣ�%�1�Gl��eV�5>�+>LP��"�z��&}1��^�
�����SJ��M�zޱ�`�)�y��B��^��z�O�Qߺ���8z}��x�nW��p�u9c�U{wv��2��=\�7�����Z�Uqc������ȟܪUK���}��6��e���Y�Y8�e�}����?K�Y^wA�#���,���A�X�b�U!�>[پ׳�7�P�Ow�k�g�;ub��~2<����u���q�s�<�Ie�$�2����%zU���w�2�ܮ{�ل�KJqe�O����V^��+|������߯��'Ʈ���&kF����:K��(��H�_#P�}�QK��g�v��l{ԇ}���k���E��w��v�ĢNϾd�4}$LKu��/��!���B���[g>�������}d֯j�}2^^�]S�]��z����2�%�%��I�P��|to�S�*9QJ����3�,���}h�¨�ݮ|��rttb�6�������)�5��_:h���.E��=[fe����D�mo�@��E\���{������E�b����_E� ���6佹&�a��$&��{C������16��k=�R���,�]K�uJ��'��D����>P�h��!Qs�	���U���xм�R�K��I��^���u}������������������6�>���f�b���d��Y=a�Y��Na;^zo��X��ʫ�o�uFw�����|kzX�]�c�܋������;�/f�����:|J�X"�o�^7՝Oy��E�@�i�.w��q��W���:�������<g=4������˚F�����mzF�J'j�ٳ�Q묯#������n3�_�K����ׇy��{�+�3�R�7��<��43�sܷ��s�r���:t;9���w�\lԯ���[�q�^P��,��餷V�p�r8O���+��,^��i�KE��t��^�Pr?�����e���݀�w���t�q<4�ng��.��R��9�~+>��7�!����[S������ �b��,fr�9������~z|�PeG��.!ht���?�^�<���Q��e��Ğ�zy���93�[{����*�]L�n��y�ǖ!���F{���r=�G���c�r%� ��I���5uD��35|�B�OnV�_Y�C�,�y7S�J �կ:�u����"�7R{�Tmu������H��U��Y�m�V�Q�*N�儖"��jt&��Vc���7t�Ma̬.�#K72T�ٔ�:���	O8qM)��f,i��S����zj����>4}��K��Á?�=qe���q>6���\:w�9r|�7���c8�N�c���}�mr�8;�/���{>	u@������x�����uE{��H��7υ��>���W�=<q�}�'J�{둷�����s �J�d7<Ⅴe��m��ν�A����t�_kܿh�*��6�,��[u�e��2Y�U$7c���J�v��Ԫ�G����R�7�}2��+#�U�ÏO����;�^}�Q�+�n�j�'��^�43m���+8^�3�}vc�Oz����}5�BU��'dx\C�۟����f�@~��e� ����=��j�V=D�	�+**"}պv��v������~urn1����G�~��oϧ�����o:���\��|�*A�O��p{��alS��m���w��7�yp���
��6X׺u��Ɩ�a��}�p�~ۡ�#����(��r|�6t;���ۅt��;����@��4}��N_�K���{н��Ld?z+�^�z�
�����Ǎ�8m���g����r������*��%+��X��}�F�2P��R� p���7bk�dJ���	�r3R0O3��94�!�I�3V��!pЁC���2m���j�4�:����A�:i2�Ni�3��;TSNm��e]H���9YO��4�nL����kQ����e�w-Y�Y^d�n�^�dxdK���;^��Y��V7�;�������E����=-?���PG��-�Q?=(~_�itW <�m0�@����:L���Ho~�B�mO�M:�욼\�k��%������z�R7���U�������z{o�ǜ������s���W�S&�v��~ք��BL.����ʽ��#q�.�q��8�O��I�y�6H�΀m!w�m�O=��4�۸'������t�'�`X�rKs஦Yn�X��a�]���T=H�:�W�|�l�/K�Y�G�\>���pj9T`B(�R<��I����N^^w�'ۇ��W�_ޯZ3�����'������U3�%� Zd{nd�<t%3��Uϥ�=���rG��79�ς�޴�W���������q9�T=��D�2Y�g����ۯ{c�l�b?@�LL���d{��	���p������>��&�=�W�.un�gͱ>�WB���>�L����l��3�Q���v�/�Lk�W�7�~\�Md���c�<�ة�m��;EN���r�N|\5c�6��1��pDuA�,�,'Z+��CZ����˸�`7�އ?����L�i�
��L��:��+*�.�4o0��M*a����vaN+�u��,c�ָ�wt?\E�!J�w��A��[��uC�� d�^8�κ@���	~#M�/�E\e���9�_���S�����k�sԒ�w�|�����oޠ;��P���̚�S�����Ӄ�R���}^0��k�K���^N���p�!���~�V���'�����^پ>�8xx�a�Z{^c�~���O�����x�����Ng�Jn��d7^��5��z^�z�F��X�yS�C'2�܌��a��Z��G��=�'�a�J�ƕh;��� ����u��r!��yT�hp��zg���[�{�O��Xׄ����N���xjU��ʭ7����i�*>ZՑq+Խ�;^��)���c�ʟ^�/�;>�xZ{\3�I��?�Cne��W�o�p<�D�@q��u�t�Ź��u�m�m�{��h�"��j��7���_j��¸�x�<�<�L�L_���K�>���z�}�^v,�l?@}^�'��W�/�dEy�yg�֢��,�_I��,	�"��x�qV6<&Z�G�]�JU�w�{�wS�}~�p�����=,g�K;��q��.��=���C<I\������P����<���jPU85j[��t�� āWon�k��
�z�^�Ԕ(m�[r���ʍ� �V"w�vwPqO~T�lp�r�z�}�ޮ�����^6*I��iX�K��9"[�R�Uʹ�"�o[F^ �Sj��%
�iG�ge۾��.8���w4梡p���ȑQg�ӑ.�]�y�����^eyIê#�HN����Ǟw�=QQѧ���D��|ȁ��:�l���h��+��W�!�v��{��I��I�����/3�x��1��/�U�k�L�( �>�s��/��	��|�G[~��+ӕ�n��q� {o۫7V,��7���޾��e�K
Kf�I�K�!WR��܈�+��rHbW���$E�oz���6=杩7��O�}��>�k@�6��s�ff�*�Q.{Ƈ���N<��������N����>6ר�[��Y�o���f�c���8�'�>q޸�*}�j��oXK�0u�`���5��c����'��?P���{��Z�h�}�l[�t��;�6}���Q;c��N�t�t�/��z�48μ�n��u�G����`��������j�Ձe�;w�#<|No�͝ڇu��n Խ'J��\gZ��}���Ϟ�1>����J�.}�7'�y�A[����^*�r�N��=;��KQ���
W�c�d_i �.��D_��4�X1��e���h��{�=�ש����qrb���C�ej���{	�u�I]�ɉ��f,w���J;or�ǷOv��]����l<΋�޺�V:�JqR�
���wùwR-	�qȟQۼ�]B�Q��:���g}Ҧ�l�zw�d{��/_#��gB�T�.2�����eV��eU���=�r�͟Ar�q������9�~+")���~�f/�[S��������Rܗ0(�+��u��W=S:�R����
1�r���~�ⲽHydZ�5�,�b�)��K�s,{u󙮣�I@ƣ�2�	'��W]xKǏ,Cȁ���Ͻ�}��#�q�[�y�*����]t��Z8+��d�j!�$�3 �ye���q>7���\:w�9�'�z=[�\�-�kf��g>��v}��#mz���� r�������@-��h4T;��3�y�!׸l.�[wogˏ������<��둷��j��,��ؙ ���o�_�T�O���将X��c=W��{=�Wl��]$c����w�;��{޸��ό�IeB�!���G�*�9ύV�N{|������hz+g���a��du�j��O��������Q�9�ϑ�:�"��ȱ��e{�ۛ�PUs�����]5�T:|��.>N���IS%�XЪ0�DDG�����UZ������km������j�Z�Ū����uU�m���Uk[o��V����UZ����Uk[o��U�m�몭km�UZ�ۭU�m�6�����5U�m��UZ�����ֶ���V����Uk[o�Z�Z���������������)��?�l�l�0(���1$���
J�
���XD�Tic*�@���4�M�Ռ�jKlm�d
�Zb%H���:*�$�5(�"U[Bj�E	T�a"�YiJڴ+URm�+m��Ֆ1)k[KkY��mZ[6L�2�Z�4�԰�F�J-5���]���f���km�wPT�VՕ��h��mk[v�Ԡ��J���UP#fjb5�mX����d�U���Z�V�0t�m�5�ZڵPH��V��2��am����̛F�w5��֭i��E�l���hٲՕ�  ��ڻT�j�>\(ꕵ���:�v�́�=ڢ��⨠�˵؊ q���z޼k� *�m���js�T�j�����m��R�kF��7�   N��z֎�v�B��u�UR��(x�(x޸�=4Q@h��� z   -���E  :F�x��C@  ��p  �7^��(�@  �Ξ�g��q��kV�iI�j�   � �5G��z��sj]�{\n�����n�Z� #��4U)���N��Z�� ���ƪ��X	���jə1�2V�U��lR|   3}�jG۽[ހʊ�y��NV�c��UUveWg�1�t� ���V�ݎ�{��j�C[ۻvr��{� �������]��U�kj��[M���ֹk|   �zխ�(}+���:W�U��5��utgg�=Ӆ�=�N�ݵ�S����,�8
��۫nWmV�@;��V���M1��E�&$h�Ck�Y��6UD�b��Zggv�|   <�/Tη^r��N��۸n�(�F+ݪ���Kh��Mc=v{��MR��P�on �^��@�λiԱ�m�Q��ܵ+T���7n٨SJ�f�F�I�
g�  ����lMu:�} ��Z�T֛m7�;h5��vwM%�rn�]�{5�z����]7�m�����t�k{�[��ځ�������vk���ٻdWb�e��1,�K^��  v��:7�]�e�؃CC���릲=ݜ�Ѫi��.�n�ѻ]%;��kM;�@�.����N��{�<�h��;�{��Ju�Nնլٶ�j����Ѭ�*π �r��l4hW.T�G�v��׭��禚C��㇫��v�c{�oo/`6��uo[��i�(ct�l#�ng��:z�Mm�{�S�E��:z�ؚ�Z{hJ�N̦�kZm�  ݭ�l�˟s��k���^�t�
Wq�ȶSK㝞�����z�B�(���͠�{�n�dQ�[�vu½�Up==:�����	�T�(0� )�IJR   j���b�J�  ���U"i�  j��UM d��&���
��� ��O�ߘ�����Gm�?K��/Y����u�7s:����<����x�Y��IN�� ILHB!!��IO�$ I?�	!H��BC����������Z���Mh9_�k)��?+���Գ��%K\��n�Etb��~���ɵϪ�,S�B�ʒ���L��WK�Ĭؚ5ۘ��4h��/[(TM���`4�V7-!C^�T���n�c+@[���ѱr��+dbBKi+h���O�&ք*�M�v�e���/͊�BMJȖ�vi����Ehŗ��$җ�T8��oF�wJ[���GTR]��R�%,Q̽i����=��4,��Wy�*�+AP)80^l�;�Z�DI�h�J��������Ƶdw�0�(ͼext�Ie�(�Y�4ֵX��o`��-��+v�D��8�j�T��r<��e�*�<���ӊ�o7�"Մ��x݂tN�kR�,���A�J��4��6�5P����9e���n���#n���6̋Z;�U�HG�l�%�E�D��.ԗR�e��Md(]&%Gt�vv��q�f�634�F�7�-t"(�sQڐm�6�h�5�%����U��&�v�İ��͌֒c��g6��*�p�vR�M�L�2MO(*���/~�Ʌ�j��5��b�UՀ$ n���'#�3v��{Lk��1[`��i�dx�#���zfػ�6�	��"3~�s�4\�N�f�>���=u��e��cѤEC h�Nҭ�3����-D̕���4�įB�:31�C,�4�H�swb�K>�Mi�oO҆%V��y���[��˙I��9*��ɵ��С d�ǂ�F:H��H��9A���R��&�����N��:&X�ɪ�.ºr�]�%b�Q�UCl,*}���F8/2ۧ��ƓY�h�^�Aڻ���ۿ�PZ�o�J�Ьŷd���a[4������ͨ*���ɭ:N��sJ�u�*5z��u��H�;���)�8T����J�WDʅn̻:��zN��ѣ��2�39J)LS�|�{��A�,���ㄿ!uam�d�ˆ�FA�,%�P��n��*�!���ײķvQl��Q����c�՘7n�j1*L,�X��ё�9A�9.T2qZ�(�f��l�i�2���f\��+�k4�fe�`�h�\F��3�&��V��jd/^����q�n�9ePS4� �zbӹ�f�.�5�-"�f��Nc�S)5t4�`JE�kr�p�y#B��߷&@FI�ݭcv��-(Cz��R��FHۨv�"j�Cŏ�`Å�Y[�����x��D�Kj�3,YuL[����v�6�C3�rYٔ����b�������A�X�ր������l�S��*�f�Hl���c6�=�Z\���K?1�+v���f%��ӭfY�
t�gR�o0lU��*0&�SC��5��oF��JY��E�=L����N�*p�k[!�T3(�n�VkkI�!j^��+�hB�0�D<j,x�����=�Fn@��+Dz����ǈn�!�0+paĤwr�"5h@e"(k޳5����zF���E�Fw"(ll�,���
�Y"NP��$Z��iV,�3�Vs&��{����t'��ک/��h�(�Ҵ�cvU�m [̗��BK�,��մ0SM��HZ�݌A�I�ihM'`-�^�o2�7��
������N�	E�e,
����Jk�Z]QgFn�kjڔX�����6	YIe�b�ح4eYX1���N@��J��)�z!4YC6z�-^��T�#E��c�)��U�<tY�.�E���h�z������T������)�}�DѤnk�pop}��=�.�$5U�b�o^e��5b��Ӭj��6�^���D�1-՗�f���-t��&f��D�R�o.�5B)1����-���N��:0J� �3B�Chv6V߳aZB�D��Z8�Y�93PG��.wf���BTԶ�%�G�GV�L��Y�1�#w3cq���%��������A�r�n�m�CO2���oA�Kr,��I�4L�aThBX�jM����-Ǵl�.�h�m^�		�u�3w�T�O�*Bő|�Y��
Y�E�d-�.���ݧZ�B ִ84�Ӊ&�u	VK멵x��ۆ�O���qXKf��<��(�:�5��\kji(dj���y��ݡ�9f;Z��Y�R�D<�WM$��n��=�iێ���s�6�VTk�0E�)n�f���y�T�����gAzA	����l5":��h� �*k����)���]R�w�6tQ]e��Q3^[ՙf��3fY*B��C'��I��Js�17|5b;�4�LC�m���V�z�؀ܴJ�*����3�� �!���/]�ogkm���v�)u���A��5h`wWDAN����%�pm��ۂ5gTc1�b�������f0���a�5k�O�Z�կ�GQ����I�]J2��VH�J�'�c݈�jPwZ��W����F�M�z��4�k��rdIC��1��{&`��ޑ�h�n��f�� �*+a4�6����[���S��3�LX;0��<P��)�E��P��h�����KS�����n��vdH�U⨚�7)��FH�\!=& ��&��Ge��a9�.�z
�P!�5	ˁMm6UdWy�,	3a����s
ںsw�H�E:�4cI�T�ۙƎ�!}`0fh�E����DJ�F�;�V�5�tV(��%��B�e˩kZT¬1LJ��i�+l��^[֮����T�6Y����fL�8jQ�wj<HI�-�����RR1)���)����81�9���z{XlfJaj�Zm�th�Qe���=����"n�[5nސc�7qћ��� pIB�����e�F�����A�tk���t-��8��^�R�˽�"#N����V ـ�Zzl�&4��x��Ⱦ͜`ש]X�lɁRLn�ء�J%�a[�Efҩq���^R��jjV��M�M�Y�e``�ܩf�V'��H����F���ٍ�;Vs-�(6FԬ�J��m$�	9�/塅Q�g��]㎴���&�֌3t�,�m֠��b���F>aa�K���Mc7�]�J_¢��ܷ7 eY��C���O[��6d��I��2V�N:���"d�q�;ؓ������Sm����w72��ޘpA�G/d�D�D�v�%`��ORš!���vt)B���4f��R+K��J<=�X{[��$3!�G��|0�8�T�i�vP�����^d��5&�O%إ�a�7�W�]i��ێ�S�@�.�p����J;,�z1S�6���QbD����lum����vkvĺ(����g b3.l��G	�u��4�<Ie=H�J���m`��Dt�h�IM�XYF�Ծ+n�:R&��Y(�xHǰe�#x�L�W�Hus��O��Q�ֶf���۾炑�E	p�X�i���=b6���$�+��H<�{ONG`:�
�>ш`�'4�C�
��g.�����k�`��Ime�{l%5�j��0�VF1&�!J��5��Xv�m��!L��#�_]c�L��(��[x�r֩xL H���C-<+].��FpM�N�0v��4��ֵ�Y,V%� ؽ&�@sq�G-�S�;35�\I����� �6,ѿ|�B:܄���Hw+ ���@S������[KAq�V�n���ᨥ������nn4@%7��(O������xX�/�Bs_��{D�kGDE��%D�N���E��z�L[EDJ��r�:"c;�JS��L�e��SɥT��tۥ��ʻ'�.�Ҭhh��x�.bsQ��3R�yhcy���[�����7Z�lFb{Ceɉ	$��� �*D�%M�+A�j-����&�5���(R�^^l�4c�&'��]Jګ����E��`mP�9�cS�$6Y���͖��[��n���Bm�%<gC�Uie�ǉ���)��w�e�r� o%,��Y�Ӌk6�u�R�oU��!owMÂ���+Q�ĲKFv�R�,��L}��il�**�)\�y���S��u�mjf�#��Y��&�'�
!8�ADB�;��8�2��;�WX�ym�vcT�r�B4^�lEoc�SH��[1�p�Zb��kt��>!��[�Fs�?}��h�����!�u��t��*��f�\w��
u�@����j�,h ������.���5e:٢��-܂U�z�E̓�R4ow 3d�`��3�!�Br��d��,}�(c��-���PhRl9/�-]�/Y�!�pV����F�6˸+-nh�������� �/6�,-0�������L,��V�W���'b�ˌ⃙i=윩�wN*�CB��?�ٖ-�J���')������K[�E�[ĝ�pZU�y�V��H��!Yr��)B�ͨL�4Sw+T���r�2�LS-Ƙ9h ����Ҋ4E�N�4�\Ъ���߳�yZ��k��@֋z�����7I��"	u��R���C嬊�l7ۤ���n�`�����X����1݊��c�L���y�����T+ea���Vg�\����fa-��s+.^��b��]��yk���V��n(��1��3�-܅��c���
�unM�R�ߕ�D`�R�a46/y��`:{���(�>�4�d'�v,�8�^*V����Z5��f)gR�&��Ôe�b�V�b�^Zu1jxo*Y ��Z�t�z]�X�UL��񩮥F��+?:���դ���kZ񖩪r͐�l�M�����+r�m�Ff�D -�"��7
�
�����fK�,ɒ�ف�����R��{[I�&��-7��G!v�7>��4-k���.B�C^?���;�i��Vk2iv��&�ܰЛtta���ĭÔ7/D�iV�z���<�J�6��ҖQ�;;Xn��f�8�PL�7i����6�d���hU�B!�R���-�N,Z�2��(�{ y��g]�瀫�Wvj��XC��EZ���'r	HVW�gs�V���tX�	����(�u�m1
HɁa��H�ĺeZ/Z
��t�$�`�J�4�2i����@ C%4��r�8��Iڕ��@]ؚ �����!J\�?�`Z�5�ň��w��ZuJ�����mM��\�o�B�:�e՜� �Ǆ;�%����蟦� u���m��jہ�b��{�L�!���'���nls`ݝ&)cqL���qťd�PKqk��f�p�\qٹ����u���XUnA�E�cI;���^��[����j��P%BU=��7U�� �ӷs�����wY7脍\�+5Sr�-��^������܈9����ݟn�Y6��Ciђ��x�y5�T.��ssM�yY��e [��L���Jv�t�j�b�]�r�fXZZ�w4�6��{}���S

��b�&`Fh513�B����*t~�`�*B�U�L6�A{A�jD37h��/j���K��gA�N�m��M��iB^��N;�Ol����ݍ��������Y�AS&�E���e�T��(i�2�ݔk)@[l��4;n�����h�.��ѿJOoZ��kL�V(�u7�#�
�d#p�tlq�+]��+%-�N+.L�m���][��cMzaYa���r��h�96��Y���#��	���� %��!fܫ�y�*�!�n��6���Z��t^��X��/��u9�P����+#2�L���۲��hlgh��u�Fh���8��fP|�����iLI�z�.S�ԃ����7-ޭ	���B�cj��q�ɳ#%����F�O/3n�Ć	���7(��Ǹ"��m:2&��֩8��*;�B��ʓ,��){�YN�̲fF��nۡ�&�4�kZ��i#
�W�7	�ű���0,3;ӓ�։ahZNøE �ī1�c���[%)��W�LWl+e]m�ȧ�@m:���܃t$��Ǝy�VÚ����G�m�ʼМ-��s2�9I;�M���	FF������{�q���2�������`2����٭�K9kF�Y��X6������1Z�M���DV�{/m[�񳴗ʭ7yMZ�Kzӫ�6Ӥ#4�iR�Q�I�yq���$P.��x����&Dv����:�Z�(�P��7W-��n�i=�>���<�f2�#{�̙3��VN�+n,���S��2����Y�b ���!nf���� ��[��p�iiĲ�^��5EU�z��Y}��À���Z��� hW��֕6	���I�4�-_(�Y1,(���T��l|�5��n���9{t��ej �r���i�"u�l�@w_^�ME� ԨQkJ:�����S	�Cn��M��͕h[�u���V�V��l3+U7��J����Ux�Ŏ��"�/N-8�J���N�O�_3�/��#D��I�S Sm��V�[p
�ޙٸ�Ey�d'Xl�yl�ce�Rc��n�#�m�� ���ё���T��x�6M�����U��<j\gJ��
K)CI�d"�}i�/B��6�ӵ��x�5A1�P�2��~�eּ�E��u-��qmYr�Ym�Md�g#vT�Npۊ�K��v�c�l�e�a�LhV��|��6�V&�A��ʳ�[B�l�v��N��� �;6�kkgw3V:���{��w���{G10N�b�Q�Z�0��{�+4ZT��/3H5kc�wV�ك
�H=�9���5-vNv�A�]��F���RNu�4ue��QV���f�%�q��_D�\I.k����p��@�T�C���1S�Vݬ�7g�ƫN4quJ؟j\N��Z�[�ws��]����p��ՙ������t��}�u*�po�<�>��Q�h<�fqU��>�4i9��\��܍�Zދ\)[sc�}Xf����+��"����{�Q�W��n)k*`�c���OcTRk�u
���T���w�?�L��i���2=L�:W�Us|�=
�r��[�}��;���-��R�[�
(�j��P�C�ݡ�>����L*���y������ɩ;4����~�+sa��%L9䮓���O]�5�C;��,��oF]l�����Y���gZ��s4���Qt͖Exu
DZ��Y�=��7BƎ�A����6Aב�Vy�X��)��,�j�X�w�U��}ޏh���=sޒ#�ג��/v���:8��/��:���������9ɫ��̧��e�L��ݲHATJ�}�V�W���\��賤b�Hӽ�S6�~��j�	Onfk�������)2�^o�o;\�9�V����Y.�Z�pj���4b��/�u3or���D%b�zEZI��ɖ�!Z������~k��x>��	��*�{��I�����7���7��yi�(�m˥q.�˭Aݸ<!�.ξ���e[��z8DE��Y�N���9�*E9�pp�oze��ۯP�
y�w�&�d蘂�}C:���H��I,�D^D�r�U�4P,Թd�C;,����q�Kq�&�{bg0*��9y�ҘN��Ѣl]�բ�+iP(c��� ޛ��ILb;�t�k�a]w�U��u��e�Zl�s��#{y펖�s.W(�u76�q���뮣�����Nٛ��Ñ����gur�<���r�T �/⸟��]��`ۏqм�ojmsHM�g����:P��V�J�M�Gn�y�g�ۢu1�_r���k�X{�]�����[�L7��
dwx��ը760x�����fJ�AS��S��>ݛ���a7
��s�d%��dF��h���co���q�4e��ܮ��&�G6�i�uy�(R\u�T�@��LN��6�p���7k�,�;��2�YJ�I�=��V\�C�"��p�lH-=FN����ĩwJ*A�aގ+I�wGa��H)충ZQr�EQ�{��XL��9�>�S�@��ǰ���Fg\Ac1<]����_��z	�l��B3�A�*p&�lѽ�0���fyW���ł
/XG�A�KՓQ�n�D���%X����n���G�-����v���dsS^�4:��5�3��=C&��m��m���e��ݴ�d
�|�̓d�>X�l���_.���;��!�S�����Y�"��s�$�S8�U����::���VmY��E��]��F�3��>��ݥ{�3G���a�*�_<�oP��2���gZ���݂H��
ky0�W�V��Ms�뙁��8f�Xsm@���l�u��%�$�	k�K��oX�H�oN��k�����̉�y�W����m���H��ǯk�����+8@��rK��X���sk$[�M�g7�Y�Ux��'[bR�쳠��b��Y��[��d�	�
<��ob�s� ��;6J5��{s��� ھ�R6�>�_���{ܚ�o���ʳ�=�58L��ֲ���.c^`4h�oӽ�Q�VH�w�0԰��Hd{�҄�}�{�\��|'�h��^���)�{.d	���5U���.�|Fv�u�a��f��=�L���B�S��F�c�k��5����iy����:��3D��,T8��:�o(���^f��At1�Cw��;/�Zt��6nb�1�B�t��˺��w�N"�D2�S�r�83�a>.&us�Ij����58��E�у�f:�e���H����i������˵9iz:�I����@q"����+˒r���Ln�p��[���:ZSϱ/'7e����s�-�BGNб��ǷkV�ۂ�56�#�`��7}p���o�_C��J�!��qp1K���)�㗀�����L�A�o���yP�8�֯1�X��ofm���j˩��U��⽭�xu&ﰔ=}w��rA����G��;{!��*	�ě����*�k+rj�g.A�S��)C,���v��Dt���kMq�U�@ˡ���4�`T�Lo|�����4������o4*���!e�r�^�5�]��=$����g���G+�l�$\Z
��c_x�͛�T�LK�UY�*t�-~m���6�>�>Ж���f�䝞�GyAڃ��=f�xY��|��P�E�Qʃ���h��`�;��hyM�1̪��v�׸C���Z˵��o&�oH����rV�f4��n^-���u��S�wW��RG�kq�/bM�B_]�z�:��q/^W�W5�Gm��R`��72��fI�fH�rb��V(�k��R����<�]���u-pb��D��E	8E]�%i�a���8^�G�ud/����-�{�����J:c7������*�?>J�4ǌ��Jr�%]���.����n��89���^��=ܖy����Y�cyKR+sp��'U]���u�WXl�[1s©}v'L��S�!�ķ`��콣}˺	{�v܂T��=���b|�/Q��jQ��~�q��F�g��6��C�,+��WS�t�a��;O:�[��v��sg%8B�͔�b"��x��4C���}���DnA��I���W�'t-�g�=�I�D�\:;���������\��di�xK�t�%�ץ��9;ncu���(p��-
{�i��f�5'w�:jG��Bݩ*���[�R���!�����v��3U��v���<��|���±���]�s�!�����;�A̾�&���7���؈�<�E�*|;CMP�B#o�Wo�&�L��r����/�h�:w���Nt��'g�y��Ծ�� eˬ֎�AmCv(8�Hm��n�<�v��j�QdR[�km�PwX�4a�y9����B�ʛ���=�5o4���'+i]��ٜ�\�����c{��1q�j!ô>0_MU��[���һ��v�]��4�}Wm:h��L]����{�_q�O jb��M�7���FK��;��l�JWY%ٻ�ppj+ZY$n��ܤ\��%�d11k.\ZԸ����.Ɣ�6�,����q�����S��}�׽�.�ߦd8^c�����O:}4�w\[�[%�����IudІS����I���K����n������B�t�.�%�+��!E��BT|/pN��&���9`]u��P��n��z�=�pE�IWv�z�����Y³�V�&��u�_1��m�A���{���w;`&pC;u]8�nR��\�]��Zy�YU1E����.Sp� A.��[������s���{�+�	�y����P���S�"�����w_A�r�{�.�x�6�m5����lTG�pv�u�Cs��u�"蕞8:�Bt��M�{+�55�7�U:�w�%���YF�{�w�r�
�4�
)j�o\1�����r��1dÕu���a��)����ݕ0�MM9YҸ�xI�ξD�4���W"B񖹣P�[71bmo��!Wt�L�ݞi���&�tL�C�˾#�X�ɇy?^ ���ʱ"緬��5��^E�*����ɂ��#��(�O{�&��K��EMX7�=.Sn��W;�,�'�V=�kCA�<M��Ie�u�R���1�7}=[;�9����/en^���&F�[N@��Dv�#x�f�0��
���'7�O:k��Y�ϯh�����}�eox�<Exk���VWY!��]��C�W	D��	�m_n����`Z�)���F	ČQ���N����������-��[����Z��˭���$t/�Q������hd�&Z�Wf䝊Cc����ђ�i�s����Pd���(�iK�|fa:����T&��N��CZub�n���^�t�مpb��u�%W�����O��6S��^:
�՗:�%�����L�V����ַ��`�d��*V��V���uۤ��h�]o[�9 �f�Ͳdã�����e㥌Y��n<���ϺE`\�Z��(F�$d�����v��p������}�s[4�E��Ŧ�����q���څX
v�9�}�[��dUoXL����S���+�m��{�I +T�Ռ�"ׇ��:��Y�9;OQT�C���4�Ӵ�:���LЍ��0�Yj�xH������-�%-Ӓ�k����G��0E{��0�{^BrS!g��2E��k;2gZ�&�P�7Y`�N��n�)�}���1��7�wB21n���j�+-�Ke�ҩ���t����kˈX�8T���*<�m�]\%�P�+^f�T�F��Þ���źu������3�T�W9g�A�c�z�C��n]ww�B�0�;dK�6�(�v5�����U:���E9�b�-��$n{2��7�v��޴��i�z,� �t;�����|}���Θ�Q����r�^7�.aX;�Q����%�]�[
K>��f[[�P�n7d��Y5��o�E֍U�rTjt�+l��n���෽��ȩ�����/��𝗳���j��5�CWT�T^����}���M�{��V5�i�q�AA�ڝ1�d�l���M/�B�8�t{�i6eS2nw۱����]%�Wݏ!C����K��T{\-v2�n���ul���hX]�G0_+cr�1�;�U��WJ:����F�z��3�&����*�X�~�<T�K׮=����}^Lx�{�==���C����[_17��C����m�..��9玥;6L��<&�aU�,G�˃�kS=����zۛvN.��xy����D�얥v�kr��]�/�9�Z��lm)Q��<���<0N?-,�֕����y.pR�U���Z�6��ݣA��%����cf�C�/0]7ci<�A�w�@���;ٛ��^��~�jKęYǊ)漻X��Bt*yyh�"w�����ËV��\�1�YB�\��̋�j��K:���Yi���fQܽ����&�V�n`��Y��b����[�c�gH|:�,��g�I4�������ۗZ|����]�L`q�O�:AbOe����GC�������]�L5����
��;��W��W��Ώe���.�Hg��8���ЙA_j�-�sYZ������
TJ�.���FБ+���������yl�.{�I�����H"���m�����ziR�˜�����W`S�9r�OE����A`w0��yJ�wѥ���tf��~�16!��+}S�.K
�5�2��!�7c�-N��L��V���H�mجR��8����� �7�㲯f�%�[&�ju�=`MUyPK��#6;�f���`�\�u��L��+�݃PNN8z�#�sԾi<Gz�Hwk��ܜd�h�ކ#�q?Ua�z��x��8����=.[Ei������b�۸̾��m/&�w�F���:��w�0L{�Q���{� %Y}q�ѕ�U�{37���>�;7|���8�=���eH�=z.�D���|<h�*�x臦h�x����AJ�컦�j�w݉P�<�Nt��n^�� *���Y���x�d��\q�6,����H���s��ļ~�rt��ًk�Ӻ����8/��|փ��4n�Hļ�Gt��I1�L�g`��*R�L�E�{��tƶ�֒�Gm�<�r��"6���b��')n���nc�; <4�Von>�gwu'C�L��L���⩏���re��W�y�SY������a��	*}�v�����_j�|�k�
kw�ӣF����b	eҹ�0"�*��}cX!��cI�9�!���ۅSHRr�_\כ�[xC�6�$�H������+:T%��,���m�K����+5|���/�@f���()���{a���I�G�g�^���R����pf�h�f�I�L���$6�v^qXd퇹6�tb�����^� U;2Fqы:�u�T�:�Wf�h�f�ye�^��yu8��]��%�+@�V�w�Vo\��{S]�Pf�\q��}Į��u�p��
�/�3�њ�<����0T��aX���)�=Od���9=Jc�c���0�;/u%[ْlp�Aa����>�Dn��i�t��ޮ1�������p�V��fe3�� �|���k6m�f�G*sz�z�V�ވ(���ʵ\�Ntf��(Gb���@�]m��O_/���&�'�5��8���r=�(`��n%�枑���%#�y�S�c첋���k���2�ךd��շm�Ǜ�39�e��e��@��M��Z�M�j��+ޢ��6������:�*>�l��F���wV�=�7�����EduؚFĖ̓EB���?YoE�$�!����xz}c���o�+�ח�t���J�[�8(S��R�M�9��Ӌ+k�T7�}�����Bk���)v�ΗzV>�$�Yс[ӌ�R�Ҳ�I���p��w ��M>�nw�A���/e���-���F��O_ma��vP:����P]ѩu8��8n�=���)�r��I`���ŗo�κtA~�.�ߨ�a)輭��ʪ�P�^�f8K���͊5U�9��h/%'|s�����������@$$?�$�	>H�����^1�n��3�vmfeN40h��`���#Q��xY����������\��g�ŝ��vlx����"��~c�:�����8�h#8T�yRF��s�)і�фշ�J/QkJ:�LB�<�6úݷs�R��2Ж2e�%+��bmh�y�G�A<�q?y�%��,%���Z��$@D��e�dP�3�s�|A�:�vV�GD�9rt�5��(jq��I6�������A(l�=�7��[f�9����Y4�l��A�p��уVK6$/��3N�X]J*7N������8YGƆݥj�q��\�������s$���ᄞ�%"ž�wX�pJ�՝���o�42��BW=�,;�:��m�+�Y�qI�"��ZU%g�`*)Yx�Dh-�6+��T���Ƈl�O�i�'G���ͧ3+��.�#`S���˶�uޱw�T?i�{�Լ�
R�����p��o��-un�C�Ք�-V��*pU�u��Tuf�SJΐF�/�@,����:*��e��k�� �>V�^���?i��t�}#�h
��;���rh۵���\ҷ9������:�k��:�k&+��ح&p&}(Hy��v�oY,�@%�x�7Ux1�~	�Ϗ����Y�cP�ZC�$�}N�;k��=�@R�����"MfD/H�_s�v=��\I���Pvv�e�����pω�}1�!HCΝj퓝�]Z)�G��{|��|�{���ު�׶vЮ��
��ye|�0�[MrZ�=�3{��USq�W���R�پ�x��F�|*
��"��bS5�/�rt���8��S�B$6jK�9��Kfϋd��s3/#n�̖*3j�Cm*��������X�Ci���&哻6M�W�垛6��ѥRl\u�4�c��^�s�ȵ��+�=�a-9-�j8N���u�U�������_V/���Z�#��X�`-�F�u�Z�,vƌ},ܧ!�˦�g_dKo�[��\�N��x��aɁ(d��/W"�#K��gGSRRb��׃lG#�("���aD�<���ʥ��z����n�sc��IiҴ*�W$N��d������wbGif(�$匵-­x�������YGL�wIQ���.:&)�p�Dѡ�j];|�o��׶2}�@+�^q�-Q�mjX���띍�ӏ&]���8�E=3X���^�r�{"�Z���=<ht6��n� �7�!�}�F<$��$]u�� �=S���z��V���f�`�Ⱥ�
.<)���͋�vŠ�����~%G{N7��y�_̊L1\��}yk"������I�_2o�E��c@�S<m�y�)	���ǲ�V��|W��Wj�(Eso����`!v�v��6�K#x_Y2S=��{�:irEea��S�1L~O4k�0Y�k�6m���0#�"�IX�&cMޞbԳ�,
ʖ�^�{E�XE���t��G]�R^J�Soj��\��%��鵽��<l�v�dʳ��w�m�f����׈�nu�ٌٳL۴{��Oq�ƻ���^��k������fX��;�gL\Wbpح3K�z�v�ɽɁNLy�c��dK��U�����x��� S�u��ï�,���<]F��%>5��5�*q{��e�9>}�/֚�k�3�t�)��k:�%f��ł@�ؖ�8��1�*c�\hgt�i��8OQ�;l�0.�#$��R�vLzΊ��e�.�p��{r]��7g�>u?;��W2	+�%LiܥVHx6���Һ��X�t.ɰ��V:|H��lwB&vASWsU>y��OE}8����W����A@H�7w�
IV��W����w���8mc�ڥ�X�`�3z���M^�Za	�Up��׸���
<�ӫݢ�;��&l#�d�CRl3.>�Z�3��Nǎ�7IǴBA�U��b�;	�y7<7l��y��^\�9����z��IsG�Yh��)��W���I�	T��%��pF���+�lk� cho��h��ޣI>�f�=5v��뾱��n��g�@��ѭ3���G3���Ylu�ѫ�=s�7���X��w?B����HS��,<Rif�cKf�%;���l���hk�h�|�X[�㗧x>�&5;��Y�!{}ټp� �mޛn����!x�ȶ��g�|6T�_C����.�51E��K�V8����6�s���<����gW,�6�>�DW+�S��Z�{�U�y������U���K�`'�:>�'p��‾��xm gt�r�[�Noi�R�,�OX�s�楙��q�V�r�u���:��V0�ǜ�dj�^۴�e^��9ϴ���f"a}3N���1�8k�ڻx�2
�w��u�JU9�}y�m`[�����"�fj�a�za�۴
��I$�Y�l+VT��I]�;nT�ŃD�F��-��ۉ"�3�yَ�s��|5��Ny<��0��,����u��1.E�lvb�aoεYJ�ݲ��
\HD���*V;cR}18���4�w�1v��ժ;y2v��
X���%k���J��Q�=��`Jr��w!��kJ'F���
���Je�J�L�$��s��^��cwr�Vu<� ���Mz]��y�:���l-�)�ƣ�u���c��$:���[[zN��C0;���?_!4$;�y�Eh�������.hv�ugU�Gu���5�K��\���N{c|��\/�:n�R}�իh��^�`�J]���3f�÷����8��r�3*��ā�Z��C �e*���Z|��K���{R��Ϳ���\ӎ��w�-�y�"���|̫�o�*Rqu��O/f�y�"�	�&��B16��!so)FF�u�\���u|n�28���ZD�M�H@c�=�W���՛��ˤ�S  �������rשe���Ӯ(z��8_o�;�up��S^-��jq���ؗ������[(d̚�fnp2�Ҍ�ϓ%H��M�!|*Y�����.q�|���,���]aq�l���
s�K^5���7��Bu���5�hƄw,N����![����m�*"�J��5,+eS���r�;ye�O�l�G�8�o/FPPv���kD9ܵ;�r��7]�5v�ǌ- Q�7�̮���v��r�I�_ ;�e7�A{�5y�T#���+.c���X�m?[m���q���kS8D��s�G[�3��c1��}{�[��td�by!�<f�ھ�Aj�CkG��K�8�v�"���&P����vMp�Yd�݀��w+rP��1.$֖t%�k^�#��E�\�����j?/�mj"ccIc�_`O��}`7+��w�A[{Zw�����*ՄY�E��^�K-�
<qN� s�S�i��xHn_JRep7!wxb=_y�����Tjӹ�f�Zuo���-���9p��Ke�]�w8��җF�9�Uö�4���LH��h}{��Q��vq.K����X:)XU�(l\�]�KB�6��:.�χk�{&2m�=a�P���)ܬ�5P\�Ƕ�c�v]�1׺�w=�� n�݊&e6��N����L4i(㾹x1����"�3-��	k��x��v<�>�E��16V�r7�`��"s�b���F���\����57�d| ��[�:�Tz��b.rÜ;��L�[�c���X���B��^���v,w)52uf��xNzَ1�*��i|{X�]{�dm�b�㬸q�M몾���e��r�\�nz^ �1�Z�n���0+Z辝�71�؛w�)�ވ���V�W���z�$r��ж965����;cTġ
�mBګ�hSSW1W�;�l���.)����R>�%��s��g���m�)W�h8"�J�(T�h�Ib��z쫭XvtȚ���hkv��N�OM��1$�b`����76<���W��IM��M�\�byNe�v��u7貛�.,=e(���@�1v�ݜ2��6��*����_2XD,�n��7��L7�쮑��A�o�wr���Ю�Ui���*j,f�#By[1E�S����+TGί� �d.f�W��v���Tf��V����� %Sk;�N�p0�|�I���R岜��5�TlLF��YPf��L�2�:8�N�aD��]�p{�КS����v���>Sd�&��V)�u�ͧ#�Yon_e�{ܸ�?aF�(V���1B���9v���H���>6y�n�^۠���/�w]N�x�m@P�G[P��'[Na��qà,o,a^v�ñj�����B7����m3
bj[�L<�&!v@D�o���gE�L)NgU�X�����n��;�r��8N����NQ��Z����v�u;	F�s����Yծs
���R �5�w^Q�7Wt�gr�2+��.�Ll�0<�Sv����s'�&ܘ"��f�� ���W[��Sر�q`9�;lKggo'#Y��g_v�V�[Ze��h4ϸ���t6���d�|��ʝ�J�5�]r��_����l��1֧3��q[5b*��m��p�偻�3T������t+;X+<�%*�
���2�o*�k���,�͠(���Ɇ+�b앁�*:x�L��wzbf<���Z��Z�$�őq(g�[�"��/�`����{�/�����
4�l'd�(��Vs;Y�H���Fq���M���:�C3q���XD��{M]n��5��T����4��1�MH��؅�K6}��4ӧ�s��>�3!�t�U��xC�ɑz��Q��v!���tE��O1�c5i��<1:#v��2m)��S3��=�;�v��j܋�#���m|N����9T|���dp�p+�s���E��i"E��t�`p#�.ښ��n���c�0eA��N RH�ݐ��Nπ��颱K�a'x<��)vW�(�0oM�:�Ě,�+ޫX��T��U�a[�c����@h_a��@�P$M5
B�p]�q9{KDO��]�!��q.��q�/�H��Q����(Z�,���Nc�P� ��P�x�!ß����Ru���rR�YZ�:t��P��ռ���xRJg�EwMՙ6���\BRD}��4��n�&qKZm�t��؊#t.Y��X=b���˝�"Wϵ(iG�c�v=���a�.U�C6����ỗvw�#��y�^I!
T��[��k�:ݚt�H�����2�T�ru�7��6S)ʂ3��'�.��j��E3���CuE�����23W��`�纾���2�7o���9��n7�����S��f��0~tNYb=�WQ�c,>��f�S��5Ws� \�}���H�KN���&��>ڻU��:�m�.M;�c~%��Ps�9j�A�P�I�}�'<��t���ޣd}�V���v&���9��_a�0.��w|��ى��ɳx��8	�5�tyWU.�Z��6ܸ���p���]�]"�N2W��8�y�+��I��>!&:@���k�A���N3�<�I됯	��3���->u��(p��.�nLy�jξ.��{AY��P��1���Y�'�p#/+#T�đD`�Ǐ�ix>�m����B>װ\̦\�Kƭ<�l��{2��� ���1N�Gf`�cb�[$�0��3r�ǟICZL?d�3�!���;�M��TX��w�����J�)�m\�6�z	������x](���\���H��;F�X�@��l�&���c3g��N�:�nu7v�bA~��%ʥJ��<�����;�?b=�N�P�`�p$w��|��⏹��DgZX㽏�4���10�-�m��K®�D
���X�dPj�^Cz��.�
&mZ�K�t�=O�wH8��w:�C⒧J�6�)F n1{>uQ�eS����ϔ��q���P:X(�3�f=�z�R�+����Y���J��и��$��
D��o1�ni;���C�ܴ�«��C�u],�ŃX� �U��
ŕ`-$��WdhIbHލƙ�$��n�%�w#�Lv9v:ޣ��V>�!��s��&M̵�𴭗��ȏ9���LA��t�� ^�;�sE��0��m���6� �U9�%*��ۼ0H|���6��՚�[�Y�������(�&����9�Y��96��7ɣ�oRjh�OzG�Q�deN%c�LH�͂�FWcѓwH���E�]4e�E�c���=ݯ���E;i]�n������B�O�n!�v�MȞ�s&{aG����D���%/�X�o����w3���A����4�m�w��v�fW��M�ґx��;���|�ei���\�1LDXd���3W6�y�i�(+��ٙ����g��k��B�S^�}1K3/:. N�2>yl���+��zw\۠p��\�>�A�I<�#]�Ւs�Wiaj���X��pV���IsKy��m���5�cᙱ�VT��Z"M������?7�דH�Ԓ��]I�텰*���;#�u���A+Y�[$��Y(���SJ�ː�RJ���5!l3��z�4�`�)(�n�a+Xq�˗� u�����"�ţ%m�f��/��tR��@K�2��&��f	�X�<��H[�P��|�Ia��l��Lך�:��f�X�˱ɰ���\��5�>��d����4g�Og���7E3������c��%�nbT�'5�JI�]��I�C��d����,ǔ�鍜�}��6� I��K(}�j>�>�����f�z�%���)�}�_���*�B��tD`��'\ba�˷u�6f�2�yJ��\�`[ʹ^a�AiA��y�����?�	!H��+����nO��~���EEf�����)��.��Y�ltG���b�Ѝv�Ū��+U�֋�t����Y�l�aBAۍ����Y��e>!H�R9��ޘ�)�8�\�/&�.�X��K�JF�)K��		V&L�������窼����l	��sE����u{ϑ��nQ�Ƚ*�˗;;P)�S���ǩ"�_��+L������8zm���6�՝��b>l��.���M2�_��i@��m�c�9/=�o�T��N-��yӘ�b&?wU�֯9�G�xҽ�c��r������G�g@ov�������Q��"/�Ac�W��qM�)�-aN�c�z'�i�&]ʱ��އ��U�ɪ��*�ڎT�yY�K���Ӳ�}��!�}3*���n���7�%�����[���3+:�:S[��j��N����H��0,��̰�ɍ�N�?��mY�8[��[�5��EfN��c�A޷�cG��p��xJs��Q���l��;��v�`��]e�al௕��,K�֚uag��c�r]f�u.��ن�`}�5wח��9fL|A�k�v�����OEq�8�\C���lu���gq
ǖ{m��1��B�*�Z�z�P:��awz���lލ�՛���
��aL�Zir��m��yӴkTp#�+l.M����t�ʡ�N�7a���Q���QX�mTR�Z
��-���L`�F�j)�QL2�U�j�)D��-6��5lR�[A��R���DKcQ�[m+m)T���FZ�F�+*��֕�lVTPiE�R�mD���R(Q--�bZ�mm���[F�[-ja�*�m��-�KZV�F�J$�mcAmKij5
U���5�kU-jѴ,-�JQVTKH�D��-��\Kl��Z*ն��Z�J[j�V�ڢ5�j5`���Ɣ���Z[\&ZĥK-j4j�mJZV�X%)Z��J�����J(�b��*)R�mQV�m�Զ����ZYhحaDZ��Z)m
�-j�(���Z��
�eT�)T����Q�DHե&0U�եjUA6� �D)EmV���֊֖������kD�e-���6��AkU�[mV%������G� ���!ǉ�T���;A] e�����mu�'SX�w�������n=0�8N�.��[�+F��;�vī�Ғ��O�Q�p���!A_�����)���CLJ|�|�V�F���w�\߳:�CǸh�~i1��S��ol��1�2&5�|��הs�1?}2�%��$�}��%�^��:��Z��ѯjs�k����}��\ܔ۴f	Xap�h�
|�J�TD)r�ɰpu�p�trG���VyV4��q�
U����EI��J%�Ox��w���$��yլ���G��kl���V!�DpvoO$��㖃�ƥ�ఽO�e:��x�宦�W�t=�;̋Y1�AAεoЯ�l�˼���S^C�>!z��,�мɑ�<�eן�m#�<���x@+��̘�%e�F����+�.�ޥ:�vv��M���،���m��U�<�2�G1�ط�����J�Ϩ;�����o��Z�?4�3����<��^�3)���Ga���m?����ٻF� ��m�(ݼ�/N�����BӠ��`�Z%�s��-eif];���NX�����n%)�1]�Vr���+�n�f�B�,2\�JV��d����
�3�:=z��=��4]}%��/3����{W գ��u{��O0�xw!p��3�>ҡ�Nۛ�^�զĻ�f�o�p;��(��s��0�������)bN��:aů�}������>\k��U��R��&��D��QE�qC�P�^瞴ұV=<o:�w���$���6{̲��O%��+��Uq�.����l�FE<���#�w������<����ݿU��	]V8����wk�iqqe̱����y�)�aS���sd���#�\{Zh<�����/D��D�r٠�O��ØAS�:{e ��b�[�ЦrurQ��:����~�3�sXt_����%�<�
��*+�}y��e�N�������+����^TJ��!�7,k���<ʖ��j4�Zo`���r�����1� Vx�+)8����L��Qՙ��"⸃��F-���Z���ƴ���Oo���!������[	3�!�j;pvv_���4 �{�9���g2=~��
}�2�s��	)�L���X���E@�p�myx7i�m瑛mK�G��{�V�{���^\`�֒��
Jr�K
���t�������M,�r�U��w����i�K6>�W�1����������4����[�w��gٛ+�P�1�]��E{vh�BAʷ�_!�wQ���IVK�/�L��(K&�f$�xcXқ)�g���J̘&,� 	��CW�X�HƠ���Ҭ�3��tx�r7��y	lǧ�З�,k�J�<�E��[ҽ�u����L�kB�:S��g��R>� B���CmH��׆���qY����"���i����'(�ua�<1{���=5f`��>�cVPd{�ݰs�ؠ��gS���������Q׬�=���wrԮ���U����e�ǣ�3��܅K<�jyA����u�.��u�5�������w5B�>��a��g��`|e$�zU?0�^ c�o���1]Hud���ۨ�+Z\�jrrޯ	Ƈ�`3�@�-ir��U�%���	pF���u�D��r%[�ݜ�����x/���V��S��������XuСZ �r��e����b���=-﷞gj�J��.��pr�}+n�	֌��谹�y�P�W�֏!05�o!��w.k�wG�"C�J52���֙�n樽P��V8������	�=u���q��[�ڻ�T�m�Y�2m���ϭ/���{�<�u~�gb5��G� �0�Y��X-�.a��q��D�wp�uy���s�Z��k��>���� 5n󸝈\]LX@_[�:��*��g���n��T�],A�)p����D|��M�٬�V��s���/uuv�*Mn����ۊ�����1O�;wݽ�-,N�9=�J���QI�N���.P~��x�˧U�{������z!�S��-t��>C;�����~�m���W��e��R}v�Q���Z:Ӽ{q�v���N��7��{��SE�!���~���v��X��J�������.�sn���p�-���џPwS�]�:HkD�����>�,R�p=3<�^<���w��c�ۘ���^ڵ鸥l{�/��^ͳ}הe�2��\~��c+r_���Nݟ뛭������{~�x���ʩ�ڊƁ[�9^}���Q�Oޭ2�%y�y��t���-����۟)ט�g#���]��)��^lw�
8���y=�^�6NG8O�鱜�r�N[p�Ǿ'�Q�����ԡ��S����������1��:p.z�L�>�C��,�C��Zrs���[�;ٙ腳ZI��tp��	T��y���:��6�]L[wصm��v>���l@���]����;���5�T�c��1*L���|�s�g�%�=pd]m�]�!�4�<����؋���6�a��<��֏f��={����Yk�N_�v6t=2{�)�ـ���l�=�^Zv�s�[�w��^6�u�%��E|u�	s��Wrl��8�z_��\�ә8j�֊����v����^������!��>Q�y���>��t⣔"Ӥ��}�Bz�(t�=�x��v]:!}�a�ψ��/���m����>S�؛ʷ>i��_���3��}u%h�d 5�5��Օ��t^7�x$vo�q���f�׷�9�پ�=��Rm�,GD����{x)=�g�ޔ���>0-Ϋ��_��]�̒��1n�I�-�7M��n�ܹ�c�	��o��W!u���3��C�E%1��<����,�j�}�=�L����{����iٽ�D�R=�� .�2���y}��6z�3᳘�o�gV��`���~t}-�|���˯+��KM��F���yeo:pJ��{�˞��"�0���U��k\��ѕo� k:AG����߼��{}�N�E^h� ��gy�������&e���ٳ�ct�v�����r��-��2�&,��A����	��ά��eX�驨Mp�����y��z��7�LzrOm�oȠ����xV��s���๱������x�uz�9��3��j?.�^��z5\S�e%y�{��o3������(�y�܁O�� ���p�rӗ�G��w��<qݺ���陏����g�6��a�Z�u��leh�_x�m떜�]��$�П_�2YގwDI^���#OQӮש��l�Lu���`�1+���{�9Ud�G����uz�=�7�ٍ��t��:��u�6nL#���&)�k:�ޝ���8eL�o{3�wk����|Y�G\#���a�����r��?fl�+g��^sޝ�oe�y^H�e���YD\ҡ��~�M��׹�Cs�|]Λ�y���u��;�%��λ��z"��^j�{���ޏ�f&s�j�u�g���U���Խ��^5��W�k��g����
9�k��z���\Q�O|'b��5b��/�b��»/�g�����!J�����0�f+�v�z�F�]����!��U�Չzd�Nb[H����J��F9��	��w�Y�M��5���o��S�r�*0�љS�m�w7�Km.��GP�%k<h):����<z����ǎ���;����o��^�t�+E�b]Gd��^�ߩ��y�%���U�M�\|����M��k��zlV9���ϩ�;���('��%ٮ~մ��#��J��t�]>�m�}�	�871��#;�S;;�FzS�q��E���{c�W�w���}{��K�41�l?w�)b�1R�=��D�������ߪ-ޱ��nO}{�
ܖr��c<|�9�ܲ״��ܯ��w�a>J�o��������
�-9x���W��Q��Fw9����{��M�X��X^�`'�V�ٌx�p�v����3�^9��}��<q���G��9����P�q�Tl�Ҕj�ҸR'�B0ʞ�e߇ku�4ΆCo�G:p.?`�sz[}�72ݾ�3�M�<zT���3m�O;�6n�էg+;��L��:�Aqv�,���nw��=Z��Q�}�I�P�Pvm�=�_5�M,��Jk�om��1�����j�P��7|˾3����zRE<;��y���;۷�?9N���:"j���D�*k��"e�i�o�<�E:��s�*���w�eǯ-/L�<g[�@#����l��Lo�Bqb��<��wvگ\R��ɒq�=����>�x�t�ݵ*f)}�&OO~��[D>>���:��������jl��ZӖ�Vf��,l�z����o��O|셼a��>���������O:�M��j���+/��ۻ��6�i��r��J�a�vJ�x���`S����yX����eh�5���t�`�q�T���4I6�A�:�^'�����F�m����d�9��W��z:�n�h7#Ϣ�/��rW�����d0h{'*��y۵~s���vg`��w�y۳0wBh8|�c{����~R�|]��b��{�o=���ח-�ٞ��{�M7�_c����|��U=��Ia���I�Wu��j�N�j�=<�>U%�u��5�JY=u��#^+�J�	cՋ���d��v+�͜������h~ �^��GP����r�Z:6�&�]ϴ��:cC=�n����$�77Vt��,��l3��Xfm��ge\��,e��R���^�u�X�HT-3Uv��\��Y�~~�<y��9�M~ߩ�+o��B��\7� �n�t�w7�l@*o*ۜns�G��������;^�'⺦��J0��붤����}^;���8+\������}#�ẽ/c�ޞ�#=���;�|��jO8�
3@_Z7�x�m���N��=4߶<qZO�u�������[o�ۣ�/N�䵨;ݍ�zd�M1����͂iԡvP���ϖ�#��T߾�f��{.e����is����Sf�{�6q�u)ۓk��M�����F��\�s1���a��S��[�h�ٳ:qBnV�h�=FE�X�Y+�S�nۻٻ��r��|=ϭ��O��̫�<v7�z}{�s��g5Y��3��}x.K�a��CY���x�2�^Խ>��>E�B�{�z�%�N齟:��*z��I�%��g#~p�����mK-��11�s�%�P�R]��y�Y�&w�u}z��9J{yu�C']�9Hw<�/�N͊'F���/E�AsM���0���!�.Ҍ_[�21ps��U�p���x[9��n��N�SsO���w^"z]:��*A٪�����l���#�=m�˵���v���f\�EL_��qڇO��_b�2��Okg_��u�d��S}K��/�zl�̚�>�䧧7&*^�'�׷���ӾÏD�'y}}�D�R=��U�]�x|'�nۤ�|�u�A�3�Ǧ3���_a�c�zh�G:���v>ӽ����|�z�ɕ�ޗ�_�q�ɏN	=�6�_��^P+\��$'zҿw����߸���M���G�P{��a��u�w�\S�֡D2�����-�6׳ݛݡ�v������)�w�ßV�a9y�����ǽ����3_+���q�6��qQ��Y�/S�����ͽp�ӫ(綴�{�ow^X}4�ݗ�wG5�f����ӯ���-�Lu�C�!W�mݳ�`[o۲x�>����}�3g�1�Y����@�v����tz��^7�:��o4�o�b�8v��2�o%����r����+����E����kgg=En<�J*��a�l����W�ye���([ 6��d)��DH� �O���(��ɬ^~��F蛾��ը���]�n�]�N*��/c�]�ÂN�W0�8��9J5z�e��K���V���D�Mv�Z���X3vM�\��m(��Y�I��@1�x�h���G �YV3��gf����t)�n�.��va�e7�7�u,i�2�K���������(�꺉u+1Y�b�M�u����q(r*�˒��Y\�����a!1�f�N���W\֊�(����RRK%�
�8b��ܓ�K���Wy�tŔ#�+��h�ߵ⊲4ý%��Nʫ齳��lE(��B#Q�gv��1��ԞU�*qa�U�e��A�D�SV���AXGw\�u^� ��9@V԰�`���)���-k	�q�X���1n뮱�6T,�Yθ�v�秌y���}J5G�[�*W�%.7�Dj{{4@��(>{�����eF�s���LҪ�on�y���n�.��u�?LA���ҥ�p���
 ��:���%re�� M�^6J����sѺ�(B��;{�b�s6sz�4��o�q�ǁ���(U:��:]�{0�H�Տg
�'��Y����ǩT���8��[��ˬ�v��<#�[���ow�Hw�/�ו���u�.+�����󳯻�̝�dN��%���Z�iu����kt���*wo�Nf�Z�a���o�������ӗ�����qT̶LS|fe�'gG��vn:Q��]�|V��՞��8G�u�Y���oya<�ė���2��Aަ�gwq9�^��(kf�Y�xzHr���Ϯ�s��M�킟<�1��rS4�<��gZ�9�w�� u��ݢv��J3���Sr�G�UЂ��@먯Gc>o������<���۶���ٴn�˧I!o(���:6볷C%*�B��uܦ����x���噫���.�����+�\�@u��	Y ~#��Z�((2n�V�\���pKl@��|�qP���-�ev��֒4Ḵ�k��/�:������wr�qy�O��}X%��!r���(b��C�{��t�Kstf�yr=8�`#w
�ԗ�.�C���3I��m�]D����a+��*��|z����d�z>�.��#���yJoTd���@��i�o��v���� :�6�	�W�y0��Í>�_5���cìVvWݳ�h��"�9�m�V��(ভ���K�I.y׷���/S_uǺ��#���fVT���_T��hb@ 7�G7�V������ImZۨ�#���׹�V�~���t���(������׊�q��}�G]j��ˣ}��]d�<ںN�^f��5i���˫s:�5�v5�>MX�Tkz�N���(�kbR�T����Q�UT�OؕG6�IkJ�bVȬj�DQm���DD���A�6��T��-�iB�Z6�Z��ш*��*�i[j�B�+Z��A�Z��ڔkVV���4�%���D���`��
Х*�	�R���L��*T���mm��%m�[V�j��R���F���eZX�-�ڪ�V�QFҪ[(�)m��*-�+`�J����J�m��Q�\[�ijŴ�kTiKR�mkQ��Ո�*���Z��e��PbƵm��A��-���hP�ڭj�6�--�m*Q����V�eX��+m+K�+F�(�����fD+Zڪ�5FŖڠ�T�	ZQER҈�B�#m�"�R��ƣQUUm)j�U�E�UF�Pm+Q��e,YTQ&Ńc���Dm��m��b	Z[*m�l�,�D��8aETb�᪖�U�h�*%�\b��Qc"��E������mB��Z�*�(�ֱ��"�Q�"��eJ�FڊT�Z	iYaVXWvk"u>��s���H��j,�����<ȣ�K.�܇�~���)2�����3'��
:f^�o�t�æb�Ǣ�WK�UxǛ���G���;�K]���A�r�ɿ->���P��y܍W�K�qsu�/$wcfbQ���nr���Wk��p@g���W��t����jo}'<�}2_^�w�uǞJy�6k�����*|��CƗN��{p�vqٍ�x��cR��f��;���?+�zy��� ޺�>gO�R{����pz���.�t
�NV�S۞��O�M��h�$ۗR�����y:\Z�������7bp훃z|�_t�\�Ň�b3�wN�a=���B��������{������vﳷng�К��1���R��N�p��FOK�I��ݴ�ߪ?)<�V�1�����ۘ���t�^���6v�Ӓ��f��kn}�r[�]����vm��z�[sCr����N׾�|���>�|AZ�(��uT]5�\�}\�U�̚љRi��cqsz��H�ƷVZ�k���P���5x��e��Q�L.��k�2�oEu�P�=���ӆ��/�pGx��3��<���l�s��t��G�P^k��+�+ZH�6�����.G��)߽�6kZ������vc���k�J�:�ҩB�0��͸�=�UU��*��W��<���+�E��|��s9l�ץ����z;�3f��%�=�H�L��
�P�4�/g]�_��l�4-Ԗ��9;��|��[��y���N.?dӛc�7�P:uʀf{9��{f��y�".+���ɵb=��1:�a�Q�����'�p孯]�������|}��\�T~gΜeLޗ�L���6q��5�Ful�]�!t:+������.����.�Lu���^�滽��.wܶvl�υ��A��d-�|�����/��E��׊.��c�K!�zk!�}yr]�a�vN����S�9UVnV�o����ߎAz����Uǂ*{�
�bI���+�d���w�xθ�߇�0�n��cm���>��t[!���e��y���W��P{.+*�N�nP�m-�h��D�΋���mC9z����a�&rä��7{�`�d�𛳒qݛ���f�q(�4�|N=�</v͂��y%e���^�{[ꂹ�_���:�a-��*b�p=��Ӡ�:��{��k�;�������e9_]��o��t'����U3�o-�ɡV$�Μ��l��R7�Əe|��n�g�:ܨ�x��<�J�=���??v&m��}S���W���U�O%��C3��z�ީB*��C��U�knx��S������ǛU�9�M~�E0,����*źf��}⤿)9���r���{hw���u��z5�7�e%yֽ�nQ�B�{fܽ��*/r"ԯUxw�p�ծXN[�z?d�=��'�Q����&�����wrNo����5l/�C���͇��;�\��&�٫�J�y1?]�F��\Vz�:vZ�v[,}Puv6m��Lw<�e�/7�矎7|�^m{���ه���:w��s���:�6��m�R#�ڡ��,����{w0��w�u1j�q��Rwa��M���^{a�~
�C>؛Z}S �}�y���[����534���F��F`|�;�:������v����qy��^k��һ<!���2a�x��=&y�`���T�ܓ2'<gT�Mǚ� �{2@�e��D.gEp�~��W8��w���9C���t3��ƽ�o
�[v��6��t��5���c����8�<����{�w]�k2���;�Η+o��w,:ȫ�G�^�[z���~��}ㄼu*md2���s^J��EOs�%�ʓ[ڡ���_��I�鳛�7�龼q{��l�9��'P6��Y��O2u���^2e�ΰ�<Ç��I<�uױ��'X�3��������}��﷿g^���N���y��Cl��p~d�a��T�'��,�'5`T�d�'����'L���&Y8�_{ m�g��wg��B��.,�����W�5���:�L&���y����:ɴ�=�B��'��̓�3�bJ�w;ċ'�`~��L�N0���C9���}�}��g�s1.�צ�����>d���	�
���Ad�5�y��,��Rq'̨t�pB��'߾ē̟�$��'rs)4����Ň�En�r�Y5�Z<�����~x�r�T�a<g�>fY<É>3�@�2��]�	>C�g}���3�py��P���Iԟ2��Xd���y��O }��;���}�����{�o�SdR?���4�ɔ�ņ�O��Ψe'��6�̞b��Y>C̞Az~�	4����q<�d�3G���N�Bdױ�2st�N�>d�%��������x�;��y�߲c��H~Jgk�.&��~ݙ�h��9T���FE��X���:�S���Tn�m0����5����J6R�X7���y٩������Уk��1��J ����x�4j��D�s$gr.�}P���͂��&3�o���XO�����?2u+!�8��>1gY'�Y��$��5���N��s�&��'��P�I�<c��L�����_��r����^�ynw3~Q�&��s]2ɦO�I��:�4���IY2��n��I�'YP�&<�LY��*~���LO�0d�&N}�T�I�T��N��=ߜ{�߳����k������Y'�=�d��	�ӌ�I��N���I�n�3�+2���m�Pɋ!�~d�d�0�6��u��}3���B?vm_���:�F�~����|��$�*x߱!Y8Þ��$�`��0��N2}��4���q��x�q%Ić�hm��lR~���d�g�$�U맄E�f�_`jA7H�W~��bn���zO�&�k�l�J���i����s��?�;a?$��qoi����'&��Ь����ĕ'��� ��މZ��%o�S{w�����L�'Ru?0�a�m�?`:���CS��|��O}C���$���xɦL�k��z�I2���'S,����������h������n�Y�����7�	PP�����,?K@�N��3��q'��l9l���sX2y�!��`>d�O�!��؞d�	�{zɦ`?b~?Y��?+�3}G��۩���U�~�w�~�&�M~��M!�y�*
n�%d�VJ�ĝI�|`��d�~3a椝g5a��'�s���I��j{�&Y>a9���7ױ˳k���˯d�N {��8̲q�5��	�6���I�>�q%J�`�:²q+'�b��d��d�a:ɴ����q�ޱ ���V�uni���&S�����I�V�Ĭ�r�a�I��?2u&�5�b
�6���ؐ�dϳ��$�L�X��I17z²q�LY:ɶO~�g�!������5�����vI���VMiNּ]�z��0r�,r��x��p�����|�B��-��W�.��dH�wx�Dja���\js7�X�n����J_h����fy����n�7Y(v�ӂ�6����*<֤��˱�V!��*�#��o�,+�䲝�U��m��������~t���H>�$�2�{�d�+��a�	��be'PR��m��pB��'���~I:�'5�.���wH�y���Yq�����y���s�sw_s�쟙6�/Ɇd�!�ٗ�L��M� m�d���<�*V�� �J�;�O$�
C'}���d�V=��6������y�|����3�[�﹍�~�����9{%p�i���a�l�JÌ�/���y���`�<ɤ�a����e��]N��!��� �J���d�VC'}���m+��ޒ�n�5w��o���}�D��ο��3>�$��N&ya4��,��0�g�&�2ì'��m2��I��N!�O ���i0�{�ɖI��}Ѯs]��=����~�����d�VC�=��2m�Nv���l��w��O�>k'�N�a6�'�Vu�i*l͇�u��$�
��m2y���o�z{?���}��cZ���k��>��N��`�2�io�<���O�N�y���=�L�$���bJ���>k'�C0Ő���<�ŝd�%L��
IL��i�o�k=��o.��n����A@�=�T�d�Vd���<�f;���	�)�N�a9=�u�6����$�$��c8��i���6���N�&,������9߱���������u�������m�u���AI0~�
d�VN}�Vd�Vw�B�y��'�d�a�{�̝~a=��2��|��I��эbJÌ������gz�������>�9��VO�e�RC�'S3�I�<�!��$��?bd�V{���'����d�;�On�~dϻ�6�L���$�x����5�kߋ��~�����g����y���<J�:�=�Vd�
�h,5Hm2y*V�:�O�8��'���y��Y��N�y�r�VO0﵍�d�&R~�3��~�ŉp��3���.}Լ�x?&t��u�;���ޓ�|F]9���B�� �GPd�u�!L�2�nf�i侳oBs[��avf=,Lܕ�����u��6:�H�� �=.v�!´�j���#���K��=�V(1���'�m���c����s#�� 
8~����|>g�̟��u��q;�%ABh9gP�6��d�N�y>�,��:����?0�fC��d��CGq���>x��:�7���?~��<�[~_�?}��K2e�)=�bO'�4�.��b��&N�d�C�s�*
��VO%d�b��d�g����͇-�u�����^3���*�U`�������Y��G��u_FI��w�ɦo-:�����'�,�I�Y�y�f{8$���IR����IY8���(a�N?������߳}����>�3�O̚O�ݰ�a�����(g{��$��=�~I�I�z����`k��,?$�3�`'��'�PXO$���++	��٪���)�}�{�ck�s��RVO�`zb�l�2q��a:���T2���O!����&Xg{��%eC�{��d����'PR;�AC�6��z��4�u�����_߳����s�sw�'R{��++	�㘑d�ؤ��i���C̝d2���O̝C����̚a�sI+*v�1d�>�py��)��[�wz��������}��{��(~d�T9�!Xi������%Ւ{;ċ'ΐ?LXq�e�g�2��C�`��d���;��,�~�����}.�]S������'����ˏ�{�<o�8�ԨL�wI:ɴ�=�B���g��̙̓k]XN��L�2~O�d�|�C�N����,�aԝ�x�x��>�X���2cf��o�פ��):�㴓(m��=��,'���q<����M{I:ɽ�>�� �'9��y�k��&�<��	��L�f/����~D_�����y=��7c��??�;��e��,�?}�6�y��N$�c�<�d�g{g�u����d㴟� �l6�6Jɦ�R|�����t�����I��}�Է�h�:�J%��#�n�n�Gv�ն���El�}�X|�v�gg[)��R]��@�QQ��5��m�%D�s@܁�]��_�W_��v�xe|0�P�(Zqx�5�R�u^_t'�����I�Ϥ/���f�;9̶����N�� >{do�Nַ�����m��u$�*Fl6Œc��<�ɞ}�6�Y<�5�x��0�;�ɖ�5/1<�߬&��d�$<G�?z����ﴚ������~n����=��/�Y>`zn��Y?0�1d>O̝fqgXN!S,<��j~ـ�'��3ϱ
���J��؄�0��py�'߯�C�_��1�|(D���$Fk��/���ߟ��No8������pJ���l6��l?�dŁ��u�1p�6��0��,'�k�N��2wx�I�O1T��Ͼ�}���p��� M��;\�7�Z���\����|���$��N�ߪ�i�'�_�Y'��ĕ����VM���i��fL\0�I���'�I�'?bI�V{߻�>�u��j�g�y�g:�o>��i��?}?8��" �Okx��L�{4�d�N{�XN�2o��J�q�Œ�a4r�B�m��Hm�y(�8ì������0c9����~�9��L'�~�6�ﬆ���|��N?!�Xa;�|�&Y2���q�d���XM��N�8%a:���ĕ	����Y9��s��wY�{���������$�&R���:��ƲN���8����2M<a�w��|�d9�|�I8����<�d����Hy�Rd�p$��=���i��޿^������󜾒��<j�%I�*J��d��}��u�l�MP�Y'Sz��J��s���I��5��2�̓�����:�h�'�,�Agi��_�u��|��]���ƵϹ���I��	�Oo8��I1�ԕ'Y?b�̛d����	���Y��O2u���^2e���%O0Ͻ�I<�u��{�g;�q�^������}�׍�i�C���(y�h,�hO!�&���'�d�%J�y�"������&�>9�'��I?2q�ޠ?~?}�	v��0�<^�o]X�U��X*���\.���4�̗^�u�kBq�5�����^*{%.�"B}�^.3��&G�:,R�ժŹ�H0�c�p��3����xh��2��J��l�-�v)4�Y@�$N�D�R�*�d/�4B��g-��9��_W�}_o[�볝���c��IR������a0����u����:ɴ�=�B��'S��8sX��d���"��X�OΓ\��'Y�9�g�y�}�v~��o�g���L��O� m2��5�c�&�T37�Ad�5�y��,��$�M����'̛���'�39�I]2N�s)4����=��<��.���?}�_w��8�~~g�C,8�~5�3,�aԟgx��e��.�y�O���<��i�w�:�	�{I:�l�{��>d���$���i��wMƻ���{^���?zpɦN'�a4�)�a>N�&�e'���6�̝b����I�<��G���Hy���L�O�����'R�2�:��Nn���K�h����?\����9��,�d��LO�>jƠL��3��L�βO���I�'��C�'PY39�$�d�Vh���O!�wɖI�{����q���:}��Ϸ�]6ɗ�Ӟ��O2wt�Oky�|���IY2���q�?$�2b��?2y31gXN0��:��5?l�y��,�����N��=�����U��ﳧ_�o��4�&�u��7�$�K�d��	�����I����ߤ�I�Sĕ�š�VM��1d>O̝L�d�@�F@B?����w�l�������7��&Ұ<�	Ry'�S=���?�<I<�W��aǬ�d�ߌI>xə�k��a:��q%Ić�6�ɶ)��'S�l�߽���s��g_~�7��l��|���8��&ܛ���'R�;�@�'����1!Y<������O�2w����4��K	�m�����G�dJ_|����?�VZAi�]��������������2q2`�M��~���~d�s��2u����`>d�'����1�'uv�,�d��`=I��u�`���M�n��>���۟mq��O�&p�a�����0�=�6�S�X��މC����$q>�;?��Ҍ]���[��[�k��D�}Y�7U- ��	�C#�/J�,Pʾ���q[|I�Ot�W��ݮ��}��jo��/v����o/v�H�Ĝe"p��*��.��U�� >������c���?��!*
�v�!Y6����$�N2�'y>���N���d�CGq����>x�qg�6�s���i����D&�N�7_�����������a�g�$�e���,��}���	�w�+'��T$�N3���Oٰ�RN����
��8w�<�6�g][���x���R3���z����}���Y2�h�pO3,�b�~�y�d�p$��s�*Vi���Y5�N�y������u�i�Շ�a8�3�N�'��p/&��T7���ﾫ�u�_�;N���a��,:�9���N��}`��O�Y��ć��&g���$�N��R��z²q�1d�&�=��}��Z�4��}��g�����P�ퟝ�e��k�Ă�&Xd���IR��;�a�	����N��3�b
d�2{�!R|����IԚk]Y']�랻��Ͽ{|����7�,�t��Y8ɤ�x�?Xq�̇�ٗ�L��M� m�d���$�Xk��$�9gRq!��I:ɴ�4{�!Rm'��8Ώ�n;�;u�����O̟f�\��|nȰ��'�&,:�4��ՆY:�~5�'�4��>���e��]�	>C�37�Ad�?k�<�Ԭ�2�}����׿o��_8��������2u+w���gy��'Y2}�I]0�N0�~I��b�XM�ɘj�,:�~�m2��I��N!�O ���ĚC�/s��.����׏���o����:�d�C}��:���he�Y>~I���q����M0>���~d�go�e�ŝd�%O��0���|,�� �.�U�ӗ�7��,����}�q���w���?!�N�㸄�&��ǰy�I4��{�̝݄����O2u�O���2m&�f�Y4���k&u
�i�d�pŝd�%O������י�	��ګSO���ؒG\;:�2:O�z���s-.�+6����+8v�%�{ŭ�mc�sO�g�g�JX�[H�H�W��Ju~W���@�&�V��ۋG
��v��:����b�dM|�u�m��WX�L�9|)Y֪t����'.��*�F�p�Js��o9yN������+8M4��gc@)	0pGc�O)�(l:bc�v<��"5S�)���A�tκE�u�#�/��V���}3!��.�ȅy��aC��t�w;c�2r.�SR8�%�^�#�(.-��k8�����𵐕��YU�����ӽWpu�1��:u��
✩��,�tP��<��3����o-O��v(5�e��L����n�H�',72�qe.��^�pU�u�(�DU�:F��Y?�o������MC�J5q����D|X��͞�X�<�5��]�:�w#�-4ln�o��	�0������X[o�(]�d���#QX���f8>y��c��{��T�f��;M�s�*�a�[0<��f]�{t�GVR��6;|޻7Ռ�\��e
=@����e��6�70>픞E����&�����;�s8�4��S�d�݆�X����z���2挩zf����"oy�nf[�"��v����Z���`��E�t"�'��X{Jp��űl���{����M��عJ�H�M"�J��'�=� u�`�08QZ��蓚wl�P���tϬo�Yp��Տ󜚳{4�j��}��� �#r�hQf�ͱ�W|�&��hjd��Tf
?GZR`�:��d9�r#�Ky�ǃ�5�浜>3e;��8�ux�]���)�}c�x�!�3�c���V�1q��}���f?_`W%\ע���Pybb�8&���jdbk�t��Y��4�ᒍ[��S�Ĩ�U����kû���>��d�9��Ir��][��Po���-�6�9l�0N��	��_��Qr��Wpb�v��V뢬#�v��<bgcה.��U�_W.��pѴ��eΓ4ޝ��ԙ�78� �#"�ieX�t�󲺋5<�ck9K��e��"r>�8�Eu������Q֮���w5�Ԓ�I���h�_^��e2ƺ���}��ȱv�[Ld������Ѭ��
�,a_0:�F&�@� �5n��םO�u͂�}J�p�)VF&3�;q��oI�qS�i���X�a�mS���`�
ӊ��K��`��L���O��T]�T;
+��{rL�*h`K<fX{�M�d���ۢ!<�k\�NT���	Q�.vW!L���v�Q�)��1�˖5�0q�'$��w��fS�u�z�NV��2�󩇠2��X��V����i)�[��6�&2��A�g]��z�wZz���t�̝7�2Y��{c�9��09�#���i��?>��:��z��f�[XY��S,�I�٭p�t�Zr�گ*ʕ�XV%�Q���m*r��b���EQ���KD��1�Jb�E�*T�Z�ƶ��QkE-(���kB�j��j�QjX�P��Q,Ke�U�b#��h-�*"�`Ҵ��eA�h*�"
�2��+ITqp�k*(*�k@Z�b����
�P�֕���TR�)kj+��"�UU+m��*)j��V�UQQPUV�Ҡ�Uh�m���e-�DEU���*)ikD��#iR��Ū���6��Q++��VV�Qc�W�\��Ո� �K���kV��E������-�*��������YQ�b[*
��UR�EDUD\4��E��iiie�,X�0�j����U+iEQT-�Q�U��Q-����+QPTU���k*
�P`�`ҵ)F������e��XT�"
�[b�iLR��-�E�#l�1J����"* �m�`��,Um� �� " ��"�UJ�b
��iE�E�bE3_�w��;k��`)�.��[X�Z��v�2��-ہL�ΩNBeRP��՝���4��d��Ltu`�?���g��1��:���_�4��cV��N��[��8������<�Lw���4^`�'_�Oz��>x���u�|�c8��i��r�Ҳ~I�c.os{�~�߱}�;�ｭ�{�!�|��{��y�?P�
I��Y<�����%a�N�f{�T!��q=�$���']0�=�M;I�gu��4_�y=�_{���~��s����P�VN$��RC�'��I6�Y��C���q��؇Y:�����+2y��$+'�=_~�������ז��;���v�\��{͟�{��J<!р���u����5�=8̫�f��/l�G�wsw���c�x��f����y�s�}N���칟I�z�:N��<��{}�O��yy2L�:��aӲ�0�|C�{�+�سL���zv�#���J�%��A�U�prw�侼��çd�5�:n��z��w�)��1�Rkڜ�ְ9�����[����"����`Ko�}��KWuߔ睭�L�r�m����/�v������ELXp=̸+[�p{Ǟ���z��\VW���ʎ�߭�÷fgt'�C��P����t��m�<�d�f�V�]Ľ��U7R$#l���Ūڮ;�M���7'U��p��`�[΢��#z��O}u��F�������VWԘ��^C��b�os�%�B�wJ�/�Ħ�F)95���sUq�����ZO�?� ��5ͭ�S:����`�o��;�p��t�U	�}��D��s��r�Lyj���FM����g�4Ό��c����/�����X�|����V��E��y��[�c+r7o�f�L{��z�ߵ�+L�k6�=�q&�*/q"澡���+���ޖ��n2�9���Ǉ�ǁSH�	s���{��,۴�h_Z#�p�Z�-��8H�јJD'sG�Rݾ�q���Tn�ơ��|���U��`w�e��	΄��'��J��:3�9�;ͻ��Ϳ�㘬�|t�<��[.���l��'��g�v��#��"���q�9�}�{�f�G��R���N�^[�gjxi���1�T�lS��gOG������y3{0	�ه�:!gEq���>{�竤Sם^��C�=�=�k��t�\\:x�5��n˯���C��v��9�b�����{k�V��6�]����S�O�-#��c�W]����Qk��i��ޝK�v��K�,�Hw��9���"������]9����\�&QWZ�^�o�Q��76�m�هM��X�}s���j�=�o�/�� }�o^�Sco��3�������jg`u~����}�s��n"F��֧�L��u��5��Ԟ�������[�Wo��~� }ؽ#t����*eL�v�x#��������^`�޴�s�-��ԫ�=�x��P[a�&��k���ֽ��Z--G��Ek�����c鶷��MzH�IlXp=1��}fߴL���ݩ9y���D�x�䗻��ow������hc�[���}��K�8�.����ٝ5����fm��ՙ��^���ޗ�_��3c&=9"z�ٸ��ޱǗ��&�'��j����v�������U��K^�\�
���g��'wM/���{^ֵ+�m�П���a�/�����v���o3{�w�z=�[�����G�����N�Qҍ��Qk�4Ut���z�U��N�	i����<]��=�A�!L�w1,<�
!z�Ƹ��L�1U=��䅬V�m�k�_k�a��3�I	�d�oh��ü+g7N4�oe�i�G:�Eݠ���D݂��Mok'5Y:�Nj��=���픴r���}���ץ��{:v�g���):`.Og�7ʼW�s>�v�~����� 3u��O*���~������\7���s��7��`l��Y�:td��C�#���3���8Zsɵ�� ��5�5^���7��WT�O���=�7;��y;��m����|}���B���y�5�.�����lr�{��r�S��E|�&�o=oϣ<�'���#�р�����u�?p\���Kٕ����-���ۓ�������mυ���tE�f\��{C}}�C-�<���^g����Z�I���W�r����`&ܰ��+Y�A?Lڬ�9�"��I���(p]�gm���' ��u�۬�dy=�h�$��=�4�� �0�۞�?bs��V5��\�A/v�j	-���Fq�}W�����|�}$~�,g�3���U������ngt'���ǧy
�G��{�2TP����gg�f�׉��')��5����7�0��C\���x�i��Ig�h�.���hȽh_]��7��F��Ơ���Ha���w`�=\F�+���g`yX!��b�ښX¦W)�]h�HVq�ñ��~���t��G�}���6��=֦{)�3��קּ�8k��;�.j[�i�:N�Lߪx���r{O_��l��m��?�혽�x�M���].+�vZY���6;��5)���^�yɌ�J��~5q�J=e�����jl���61��Zr����q�{w&W��|�^���5yߥ������}QO��)z�p��p��\������$s\����)��������rm�{#��� YN��.wL/�C���ͿQΘ��M��9��L'��������u�O��b�u��ٰ���L��M������y��̱���m���#�^��Ί;%��r�uG�k�x��YL��W�n�^y��Ĺ���^��y#�0�����9awɋ�-��/[��s+Efsfuոק��N��痓$��s�ð��a�ϱ�z�,�2��Zw2�c=�l�M�gp�L���}Yf���^�s���x�[g���'@���nXcy��Ѧ�^I`�5�'$�
�S&�n�t�9�'q�dU�t{(��=�zڽ�[@ED�rSl[BJyR��O+;.&di�Ύ�{����i��/����� >���e��SJݧ��ǻ���ϝ_�9;�r_^��Xt�T��S���|��
zU�܅팭�n`�q�8+E�&���ZU4�'�Оz;;$��>�J�^_�l����_��\7Y4��T����=���y�I��M��OxS��u�u�<����Tt.�����=v]Չ��L�O\z�k�����c�~:#>�u,vw��a�̖�3������y/M&6otx������e�~:#;^�K��z˸h�Gb�D��4�m�$����7�~�}�ޥ�q�1��I�}{/���ح]j^�	��)�oD��(�7�!{�?V'�Q�=����/�v��M�dS���u��6�M�]a{l��1�V����µ�	�x�%*mp�N�?}��]	���)����j��i�|��O�[�Z6;ų?9��n��=��u���L�'�<#�cv�J}t]˼�S�^xΜ*�^(]g+�B����青'v�wtZ�0�u�ĥ��7�@Z�V��tc~�&bBYo\M��r���fv64�#�A�d������.�6��׃�������|)�t���{��t��~ߣ�0+=@��y?|�y�P�\�����!��s�Z�I���Aк�<�0����{�l��t`���'=�X����EG)��{�O�+Y��|����W�7������ه��WC�n��h��H~i{�:�~R>.o�{���=���tr��t�Ǹ�ޛ��G�ё�}O�h֯}{���)��>
9ht�/ݝ7S;>u~���K�w�$ٹ}�Y�~�y�g^�:��Yk<O>�����;3�渪<��t�I��?[Z5�ky���׵�
se	����4{*����_�ϻG]úu���,��rο9�=�\��$��18��m˨�]V��{-5���S&��������;{��Vg�� ���\�Ň�b3���=���o���<�o�LS������\~��1�������~���e���g�i�/���R��X�ҝ#�ף{�W�Ik�Cw��-�4��]��x�]��dcj,I��.n���٨&Z7Щ�u��Zs���@��{h�sX��ɾ��*z��~ʥ̽����t���\��Mrz{7��}��UW���N~���a~�QshB����?�[zk�1�/&=4�ˢ�Txǚ���ܜ�����E+ty{~;�;6�^����YO�*��p��O�}=&'���^�����a{w����6�T�'޽�׹�
�17�oyn��l���oG�={.gF�x�>S�'ƅ�x`��]���綌���ӑ�����\.t�\��Nz�3�p+<4�8����p��}�.��kޕ�`�6��l��!��*9��߀�=���o�ܭ�i���-2p�<����m��<蓖*Wrl�d��N2�v����g��{�6F�n7�������\�X�F�_�s���Q�>k�{�wS������j�i�=�j�tp����}�5�(�9�y��҅�u��p���j����P�����ݑ�7��{K�˝v��o��7$[s�l	���ڪy�ޜ��>9C\E�K;Zy���e� flhp��v('2eM�D�Cj���+
�'m��EC����S�dbV+��̯r�T��N;��3>���|H�e[�yd:~Ҝ��<H�yB�]a���wj���]������}����G�s��?ү݁�{�K�&��>gO�Q��E�؉W-9���<����݃�`n�v��*z�^�o�n{x��P` ><o(��s�4��6�fԨ���}�%�u��l_��2~���<�q�
�vr��{���P�R���RP����۝О��[Y1z���
W��$�V��k�s����Ey����R_�,��{o�Pke�W޻���ߧ�k�`͜��ǧ#��l�a�|V����B�ޅ$V#R#;+Փ��s{Vĩ�}%� ���t�����Ɲ�����{���sfL~��SY���e�/���Z�/1��>�qﾙ����9��~G��"�~>�I�5��z6�A��.���0�~���zo-����|Nеǩ���l�wp���_�����ٰ�*9�rz���Պ	+q��qK�\d�D��/^[.
a-�:���<�}n9�9w��5���spug&��[Z'<巳�{#D�ӥn���:t�t��ܴ=���mK!y%�M���|9�ŊK�YԴ�V��f�W!�.�Ǟ�|� ���zwG���yϏ����XKe����`=2{>�e��޹G7wck:�����Y�tz�FN򋻪<k*<^H�w��ї�7�{�}̸&oK�&of	_�0��#�џ(!�Cվ���et�����/'<�~����������X��^}2L���]�y]�B��]��9qç������\�1xW�2�|�a��[Rv����"�é�/gu^�L�ͩroFрf9ש�d+�Xɺ܊�H��9Z7vןkAoV�]u^���_��ck�u�eu=����v���W���W�J�M<�n˕�S��5��6	�����%�K-���Ӽi��`>nC��W4��\L��M}���Lg/Q��	���Ķ1�~ڿz�¸\�����?[}<xk��8��1������_a�o$�����5/z��@yE�����£�Ƚ��hㇶH̽Y2=��f�Fr���2�kE��e��ޥ�Y�V.���3��@_e�L!�����s;V`����U�c�n����L�4k읝��ܑ#H���� �ľ쓃x*=�t(�?'}0�u���dݽ��:Ԡb����	���yb�}l[�l�#�ՙ�� otA��w"Odg'r:y�ٙVбl�B�b.���B�D��̥�gj�(���yzƵ�OW9.4hb�<#Sti�G)"�V�B��qZ���+���N����rLn�"��:��iulTx
a�Հ���{�����t�3�v�b8S�컕��3!�s
I��N��f0�5\��g�R�]'x�Yfit8�Z��;L��]^:�[+gq�0*X��f^)��j}չqQ���<�����7�v�+����t�ն�G{[X�G_e���BR��90z��Ґ�VX�#02���c{�gY��\���v�:��V�6t
1٩[N�r<��޼����1��f:M�̹L�r�D��k��o���յ���<]�v[����X��x�b������ޕ`��'�Z��)���n^ ٥/�� Ȩ��n�*Ζ*�M��Y*,Ws[���߳ c�ڻ�Vh_�RK��F*n�z�k��=�������w5���E*�i��ݶ��v����r6�k�F�b�x/�:��Dx��nI�N�;{�V�(�������,�G������mދ���%_9�j�B�u�4��;"�4��v�i�T�;�'0�-�aD	V'�S��D��t˲(!5�_GW1*9tj�-�B&E�i��e�T�������e+�� Fkco�w��tyˍ2��7vn}:\�7��*80KW�/�wL�S��r�0����0�LhvPVh���׻=��1@B��K�K|��4�n,�%Y9mҏ�2�1�84��{b��K�I�&��]i?�C��</�c�Z��tշ.-U��ٚ�ǧ}�>�"+j�n<21H-���Nzӂ��C�Jzi�[���vL�}�X��Z��_p-&�e��ׄE�r7�9�R�;d�KB�g>�B�u��w����cts8�>��U0mᨚ����u����#�!FE�.���b�EvVW�|v�Ry��!^��f�a7�(P����a��ٶ��~2n�����`�dV{g{6�{��{
�.�YS5�	Sx��*x�Id��e<��CF�d������!�;d{m䡒��K1��M�a�\A�s�J^Oa����'E[����ε�*��{
�֋䡻��b��Q�����u�W��ư��^��{V����ny�Ý��S�>�Ŋ��X͎��t{/���q�҂�x5\��R�Sx���Lǅg�mw[��e�b��Ӯ��9T����Ř��*)mD��[eH�U�Ã�Rł�+��hYV�Q����f)PH�lX��U.0\U�
F�Q����Ip�F�V+E����TE��j�EbEUQQ�E�p�R�E X[
��
"�E��Q�hZQ1A+X(*Ѫ��*��8K#Y[6�[e)eV#"��
DURT��Db�ұ��DDkP[JV�[*"6��k��TQ"6Ԙ�TT+DZ�-ceb�X����X(-������Z�ʴYZ�`��mb(�X�ETUQb�l��b��YT*�2��(�R���UFV(UmZ�m�F(�[+��8J"�j���	D1j�U�TQQ�)-��Q����jX#l�[AX�E���TEKh�б1J��b���Db�[KKm1e��B�h0V(��cQU&-%��Ucam�0�UQEb�+��T�@>>�$I�<��y�A��^ݛ�cb����;�م`:/s��t�x�x#�#z�?�=9�49���o'�Et_��f�c˻+���|�#S'A���S��?����|�ԗ{�g�O^�y��#myywj��v�g����@�}nWf�+� ϫe��7�����3ŎC��7����z�� 9f���X�qV��{\.��	ˬ��H�{�s������������	�Si�������;�Et�qܙ��߷y�ۉ��.Od����
�QӬ�O�c���x�i��ng^�ҩ��y�:/��)���߾��ٝn�P:tW�cz���Tw����'o�T�Ӄ>���5�k�K�L�V$�̐>�g�і��%�Q/o{�o�f�}��j�qK��fc���K��.<f��M�<w3jz�Ц��g����jD'ǫ�Ϭ!҅�}�<�{���������0rl��kܒ��\궄��B�Ӌ���g��s]��U�D�e���^ͫk��TUF�9��Un�������O4�Sc�'��4$4�rܱN�,N��G[nT%�ƓfY[s�L�XL�v�Dov�0ؚ=�.\K�(oq:m5��w`�?W����ũfjZK���k)n��,��3�}_U}�_q�߽�>ӯ�δ&��~D�������=L����֢":��hx��{e+���-̎�|�z.I�.�����m���h��Tܗr׻7�?>^�9�݄�r))���;�vc1m��ÕM�x���;�m���*�͙��o��s;�����[���̫�qc��{������A�oף=,3�]�H�^��ϟz^�(c��U>{���Xu�ٰ�����%/���=sQ�ׇ�����؟�F��}添Â��uj�G<w���t6I�Ξ����v�PO�[��d��x�ɠ��ȍa�O����y��Iy���>�q�e	F�ow��B�Ə���\2�#J^O]4�N���+�`����a9Gz�����VP�Y~G�Ƿjbҷ�E'(��	��%
�޸���~29Ӿ.>�o�&6�_��s����G"pF�����Q1T���uҡ;a�ޚ�����!C;[kۙ� ��x���w`z���R��tLlt��DL�Yo��b�A�����n]+��wn�Ǔ���'/��{�z^�`��n��w�'v<k�y6#�+�O�OW�����zs�.�n�����b�w&΀�Od�(|�mX�f��=^�j�^�{�}~sf�gFI�;bQ�,�u��s����uG�q��:��gp�we�������2��w��,�o
zX�쭝�����Ӣ��tMN�?S�� �']N�vdh����m�l��~͇m�z7�/v6�6%_�>j^��I�����(k<a�/q�g<�lK}"�Ny�=Y;�e3Ku����q���h�&ܹou���c<��t���m�`��ۭ�7y�v7Y4�Ǽ��w�����=��b.ɳ����m[��5}��=��{�v�]��w�+�P��y����h��Z�M��׷�4�3�����':ʿ*<㏕I~�o-����N+��>�\��g���y��<X�4>��m��k�꩘�z���x̰��Qypɕ��U|���8OVv/B����Mi������VJ��<ޗ ��	μ�W���<���z��@���̎+��N��Z������.̔�U��RE������]�=�O6MY�܀\2>�����UW���=p;8�Gy����r[s�����l��Q6�C�����Hf�k�O�<�`�չ\/���3�ޅʿ㱑���{w���	�uM�So�y�6͊΁?�f1c��z�'-�=�s��ܽ���&�J~�=�P�9�w��PY��C�S�>f丹�N|������ž���Z�׫ӏV[5j���m �EN�l�bL>��~\mܛ��n��zNv9�w���0��G��}��Qp�y=Y��:<��*�7�]z���|d��}����#�0��!s:(G��![�2���}�P���o�=�xy�|�t����wOjm��M�\���׃�O����;����<�����S.n}��`u~���s�%���%��j�Y]����
(���y~�z���Ŝ����>���	W)�����s�5n�������~$A|�e�����w�8����W@���P���p8wYu����م���S4��=)G��$d��gH=,tu�O�,׶j�������.+�z�h�u��#�w��.(ӻ|F�5Gv�-k?������><�|>� ����_���? ���t���x=���W�W��Sv��ms�v�͌΅z{i�Ҙ��z.OS�v;	u������wYN��s�|5�ګ��.��N{k{���4�b�M�}@;�l�_��u�x�\������{����O�y޾�JW�2,,�ϣ�t��ۇ�g��Տwa�:���ǒ��2�;��@i�`{ۙѝv`9�ӫ�Xn��/b��;��Y�/� �/ۊ�l�so�����ס�[N����������">��ı%������o����Q��O�V̹���}y~j=[�'���qjje�3�ڎz��uiĲ�ُ�۲�d���s5�:<��`�By;��b���GE�^�,.���p!V�p�.C.A�ۇ�u7��M�j
�O_�.r���96��zN�{²�f�\k��UFX��"�Cucm�����M�ϲ�L�<��ҊM�a��P�N_463{g�8�)�]K��X�L-�B��+�9�/T�&�'nL|�:�ȱ��ݝ�S�@�rY.�9Na"6˳�ט�7�8Y<C�8C/�e�ߺR*Qs�o)|�n�z#k�(�z�Q�����PV\�F��N�sq�VW���[۝׵��_� |>�=��I����ӾI!ߪ!����^
��+��8���zE��]�F�4:�i_��V�T�W_g�m4g�Ԍ
��e��T}�C�Y]=L�3S�g��΋�w	H��˒�:��S�g��1=�H<�:S/
f^SJ?S#�~uO:�����;/�nKNL���׋0?vg�;�`�#�u^�Q$z.ߪ��Q(m���7V���!�����Ϲ�Ճ\���"��(o��P�fY"�B�ZU�]�a��%�Pu�y���᮲�Gx��u���� �g�pT<0(a��eه�#@�З/�Ь5���wz:���G}u-i��^�\9�wL	+T!\��kzKGM��p���^+�ϪI<�Օz�t�w@��ywF��h;����$�U�\v�=҉�pXV�6�kRõY��n����5����`cԎz��pCҫP���s������n9�Y�c�;���� S�0��{�U� W���؜��p\�
�{i��Do+�ڇ�n,B�c�S��^[�7Rj!kn�
�c����=��u�١f��iS��+�rYΎ��W-�T�/�7��Ye{Eb��]�c�K�W"�O8\t�מ�0.���Pa��1�;3~nvM����v�H�ɅErڬ���j����D�.�s��O|������}���T�n�r���g����b��x���N}�j��U�KW�8�Oƪ0�F�J�I�-��8��Cby{ļs��.'�=�7�:�>`�{�1Ғ�|��Vrf�c�N�l�yxI�������&��8���qt��踳��{#pU��AP.�FV���.{�ݼpߒ��bK����x}�E���(��!0�l����V^�ﱚ���(�$m�� ��|����e�\^\�-�H��:��ɴ���;��o��o]��W���d��V���r�<�g�j��(/N{~��_�}�aW�ﮒ��ϸ�r���zO
���9�qŇ�Ot��ڰ6zѿ�RQ�<���:X|Y�q���q��{��ױ���vl�E����.q�Sτ�z0<ށ �H �`ܧ1��'�,�<�/��t�P�hu�kLnX�`J������qK[�����R���]���yHf�TW(W��������_ϫ�f�X�}gVb�śd��:�mh�%��u7�S̺�^�,t.�w<c��c�8���x��m��{��6������z��%؂��+��������LF��X�~Y���S�n*7w(���
oT�E&�v��k�)���S/���6u��]Lt�Vju�ܽ\U�ק��}��|v�>���>T��2�U��H�,�\EX�_*9��f,9��%`�={����}4�w�{���e�C?���=�Q"�	Լ���v����2ׅJ���׵ו�Q�4¿x���io�~���fZ2��Kٳ��J�(y�ls�I�;��^5�+�~���)f�SI�HS6�����4���)�w�)\���(ߜx� f'�dw���C�����LL�g_����'J���߹s�/�v4ϯk�A�lz&aã�[K�)�ޖ4�ZE���m:�vߧ�I�{}��z
�u+3o�pk��m��)���}�Y����Z��ǰ�����������=��Zd�zbՀ���¤G~{bm�32���˚�.˻��,��<u���HW�+ƚ��}m�m�[�^�Nq����Q�E�y��+ۢ���_V��S�C�N5zeW82��O�aV�+�H��K�C�À"�
�m~�]���qΎʾ��F\��"9��>����H��h�aӄ������G:��ǌ��Z9�|w݄�Q�ڴz�v��=:��8�Wr�Z��񋷶�ť
S�`�VqX�i:K>��b��:&�BCq����foL[�3t�\�Pҡ����[�D����2m.���޻��RS`�ȝ�tlco7�|>�}�t�t��T�ז7���F�fgN�a�=��+{��%2���Y�Q>r�"�ɜR�t���8�(����.)��혇�é��y7U�3�N�bNy�^��F^�;��¤>ݤ0=���z>T��&���\YA|��4:��ͬ�}���^���W���Y�o^�R%�.Ժ�O��w�(
��G��F�=�%3�'�P�*b¸���|��}|������ɖ׻�
%s�CƎ�c�B%'��I
�k��댼��6�+��\9���
�
]��e�Ӻ{8�6��1����������D3�J~�S��>[�R!�p�*�W�,�ҽg��Ϳ(�q��`J���Q����a�OR�����M!��3�*{U��gX����"�o͛���~��>��JK��a_��pE��Y�x���ۄD�kk����rJ�d�n�FFמ*��Y�l{s!��uـ��^"�pJ�*�������y�$�R,L��ڞ�ޙ�5�h�m���D��h�_���">�%�vFz�s�ORJn�跸�Ƃ�(ئ��R@΅�%u^g=<�zP�bXiQ����oi��mެ[����<�Z����ۤ�})�5[���t���lufV�E�]VӺ��v�*�_�s�����5��L�.4��7�� ���>��>���Y�_�{�z��A��v��*���T,ڜHʼ�?b�}��s������p�*<Ü�?!#���ּ2&ȁ��Ѷi�U�����)��i�>A��-����{�\2��)���,��r��:�<rm?-��e��h:=�$��VX�2�wj4o�zye�����A��J��QLml6�ϓ������xqvS=5)�Ǽ��9�v��m��g�C�g�T%�UDn�w�����%����Aa�a1e�k�����l~�4�]�BJG�<dHc�vy!և��}6�x<���:��l�7�?'���Uk�uv���<���"W��@j䡰��y�
fX�iK����v����L��鞿=���x���1�fq˕D Gw�@��Q�<!�3�i��x�QF"0�)��y|���,l�9�"�5�˗�
_ �W��.��9�96g�{���坓.>~�(;�E5WϦnJȃ�]���P����e�^��h�%w�&����<�Umr�$�ڻ��B:Y<����u�X�v8�.��>ү�$p�6��s7�0�	�ܻ)�x\A��Ŝ �{�'�<x�Is����jZv��X���
.�cĂ5+eH�u��%2��&��v�m]�����В�`hn3��Ҝ����\�`�%�%!��^܎��{���W��j9e��LloN��Ůѫ2��g�F�>\|��Ը�IN�'O���l��x��ڐ�
�VMx\3;���HX�Jdՙ�l�{�
�J;�.��"5��.B�ˮu��Y�.���%�A�(���k������nJ$�{�<�=�ь��n���!�����yS@Y�6�HxٻR�u6mݤ"7~�J�?2��9le\϶��҉�5��͸'(�I��(�3����u�&�'Q����h��R}t��^�����p��P���jV����ͭ�����u�ڐN"��e�٦m��D�B�I�6��"� �L����h8»�o[}�f)�ˆX��r�8ecoE��K��2#D�jE��;��O�Ь��/�xI3->�D6�ږ��!��W\�n�1��b�(0n�:�þCќε4��s��B=��ot��_A/I&�d��������*�@�2munm�ޞ ���D��nM��V�ܕ�m�l�p*��P[K�z��N�h���,)ll�����/X�ϕ�ې/��I��V,S:J����\�ba.�Z�p��n�,�!���Z'G׳9BM�Ň�9���3)�OEt�+ևh��p	��|�m�<�:�ժS0z��zU�J��%p�b�6�`5g����b_ob��8�紾���Avz��c^g/��3���t�������|��uwtWGw���ɻ���۴\@Nuy���!:�L���We.qGz�<9A�;��E�xiTp��ۤnHV��1&�W����V�*����{l�\.C��e����}��@�&���ha�6�Rw������o&*��OZ׼�X�K8�N�;驺\Z��`�S�VZ�W|Q[�M2r���mM����b;f�u�W鷆�j�8�ds�c~[�xuv�OZ�	p��n]��c+�p�Q��XP�}Ѧ֮��6z��B�Q-̊.�4��V�Jq�ݤ�[yo�WZ%�R���-F��ùN��<�RT/<����h�W6ͺ�[��,ژ=�7�7G���cv,,e�,5�^2�^<�Y�}��஘:1,נ���!g\"R�QF20�����yoa��_l@��m�-'<3���������ڴ�p�8��>�S(�cZ;nuw��S^���0�r^{��N��M�C�<�-�v��{t�f�d�����k�r��K�δ���@��1o:6�+��T����M�勫Pb\�r$�en:J��b�
bC��=|�^N+�k0�@��7[���e-�DU�����*��H��*(���fҠ�hŸ��X��KFP��8�V�l�b"�[X������1��Z(��Q-�0`�TE�"",DF*
����U�`�
1�+(�P�b��TQ�E�YF6�����0D��X"
�U-�`�f*6
��+
�b"  �*���\R����Y�Q8�EADQE#+Up�QPb�E�Kh(��TQDQcT��`�1EU`*��j�pʬQ-�J�[e1J��F*(����E�X�6�E0�
[Ub5��Q	TEb1\%Qba�*1DF)ŘC1�Ն**ł��l�V-lU0ն��"�DPX�"�"��JT("+P�TUPPU%�b���l����*,EV��(���b�lUQb�i�*�*"�QAc(a%�R�U�b�AH�(+al�R( �
�qj���U��ȳb%V��EQVb�5Tb"[*+"*"�A��_�?���sx0����_I�5ط������!R1�5@_٫���tXQz�Z׽hoaKm�k�|�����v�y׿�����m;�{�~�$tMj3�;pm�?	7}(�bJ�+�1��Qk�Ih�����Vv��"�ש���wt:��,8.�mQk.ݳ{ޙ��.;j�ɽpXW����f.�C�1 �x�'��D-��ӌ�#�j�ӣʥϓ�^��ֳx_	j��V��]ɥ�;�(�=|L+�"��*E�]��&}��z,��'�ΰ?�zXь�z�V�޻�<�ᢦ���������)���<GR�SBx]�i\n�o����=��\����"������� �7p��/m���b��.'���#��{���˅����@2�Vy���"Ry�az�<I��Cp����(���$�BzWbb.,���F���:�^2�'^�龺���� �I�ʭ7K�߮Y4�BOy"�\Ҋ�S���gc�탕=X��}=y���8Wgi��xRAanK�/*��U��ȑ����M�f��~������:���Y���ՙ�+M�xeg�j��(/N{z6M{D@ǝ�R�+\��ᅒ�:��n�%^=Wty�{)�ێu�����O+p\Vzz��p9�+su���0�w�3�$9�O��+���Uu�z���\�MW+tt��tޥ�o�7�;/h�:j$4��>B�]%��ѽ���O=ep����������\2������;�$��E����
kfR>�(|x�A-�2��8�.���w���wǌ�;�j�u���c��9���d��{%��2Ɇ�&�Hٗ��
��s'ky?rr�������8.�r�1��_��y�?|"�z�9Sz���|k=y��.��/o.Q<p��ŒJ
��*q�c6:��uf��6�L�Ev4��/}W��6j)����ڏ����a�š��I�$t7���I�U���׻f,=Β\\P�4��=[�Q�{u�����7��4��/'uA�w�oh��fU7\.��a����ˠݭ�鶰7��ө6n�q�nS$�l�H]K*J�[�MR��&��UϞ��ٰ�y>�K����G.�W��]�Q���1=Kw�z�b�XyԘ=��b4^u#X�n�9��N"Y�L�B�ۘ�]j/lz&aÎW$�=l����^�����w1:j��s�ZP2|�%�^��C��W,u�`�3����������Ĭ��K)sh�����z�9���{4d=�3��{�ywu�&&�2�j��y$^����D�9�V�w´���D�� +w���n��
�[n�Y���9�ַX���G�$�FTY52�:sV$`��kuy�:u��W�V�׶[��ߴ�da�������T�*��4;H�=�	/S3�9x�دmZ(c�:�9��}y��Bˉ���U����+��K֦Ui�S��/l{�H���g͍%�}Ku��+Ｚq�ZwT-K��a姞�b�)����WȪΔ߆���⻅�Qy���n�S6T���^��#/��E��mh�+ZΞdt�6Gh�N
�
_�pw;��tZGyA}v7��p�f{�N�a��ƶ�x���|g��}��q�m,L�Z�&ey�oؼ�#� ������.y4����.Ny�^��F^}sba����o��[���g>}N̙H�ixR��1Q�`5�g�MK�鿫�x+x�7�O[���G]�?yN�4�Ӭ��*��H�A�s�Ԧy䪄تb¸�Ϣ7�=�\��yg}ۭ�'x\���|���ܕ�b����B��k�k����h�O�j�0��Xk8tQɸe�gz��z:����l=G��N��lvA��S��z+���o��ԍ�+l�z/_���Å�oyŷ�}��Ine"�*�t&7���S/%�}���U�MKk�-GSܷ�uu�,�0,<GBr�)�����9��9���zF����X��u�.�؛��Ev.�(�/qJ]*�s?����Q��;�'?,h�y�W��t���琣5������Vh��m��m�S���{�:>o��T���j�ʆ����^�>��1���f�,/9p��,.�>�-�j�{VB}IO#E���6o�@��g�^�*��w��{����	�J�~��m%��N��1y�:��y	6t~�b_���w���i�x+��Y���2[6j��_�L��P��c���l_7���ޑs��P�=��g�ydκ��XOPcS(֨���}�%�pY�����-n<��oF��k�~�x�K�a�5�}[=P�F�|٫�>�����Cъ�s[�g]�V�C�����߇�C����\b�ZY�;���c�9������rĿ�5�E�_Og?o���ղ�E�b�X�f%=�Smx��	r����Cݳ1�}Fe�ZoS<�Mzm����%�#�(`�����uDwU6V�������Q\�옄<ի
]J7Hq۝/zlތ��DA=����k�i�āfh�v[��^�6�!��]�iK���w���n�*�1��L���j�;�9�rCB��ae��]��j*�v�p��}��U�e��z۹�т���j�:NJ��j䦕;��(L�G13�,�����か&���7�.��ʷ��fօW��Zו,��Z���]^�:;ݝ�����Ys�dk��;���(C��e%�v��94��u2�P�f&�yL�ǽ�ɨ��靸3�=���N	sȹ�<}=38�[ņ���f�V)s]�)��[�T�N$�y�ļ}�~I��֢�5��Y�{�T���(o��r��,�l�7C��0gx"�s�N�R�2��}ڧ/jޚ�W�]�k�S��������%dA���'�����2����t��k�U�w�^�U����:j\'�0��੸��#�߳:Q%�r�.���.���(
�]��똊E���=�do�F�J�@���q��]�pv�oG��'���[B6S5�g\3�k���T���Mn���+"ԽΗ+�pO�ѳ���/4��Io�xd�s���je�
�5�������z���uBHr�91o.��8o�ytH��*X��n�{��Jj�,�~��n�f�p�9��Vxe�0'������§��54�}3'�y�ˆ�ԭ-��װw��p�:�[��Ϲj��ىԵ�8�ɏGp��X}�x֖��
x�t�>����j2����Hu�+��yW�:�W���*!,�o��6m���{ݗO�2��d�P��Hm��f[������S=���l v�e`�;O%A�'݁ʏ��m���z��t��9N�*���1�#���g���Yy�	;�hǫ������{|��sl�%���u+�
���`��j.�qX�3!�˥�^3�\�]�q��v�����m��i
�xo��V�Zi�U�e�&��	6;ԋe`{J+�)�LHnSO#�<���9������.��cZȲ!��Զ,�e�*���e㻑#�N4'�)���q	ȖGO�|b~�����ʷ�86�5N�6Dq%���Kb�J��N�"�I��q�񈽅*��p}Ux���#ϩ�����}=�<s�j���G�R�G�Թ���k��?a���u�Sc�C��֡��.j���c��9��n�~~�/���OF��� =�;@���ڼ���_7��0�}օ��r�S�s�����
�aʘ�=�!�R�}�g��ݷ���k����H��)4���Ԭ��4��άϖ�\Y/!�U^��ǳ����of��)'�K�Ď��	����������R���U�7ᶼ<~�nfN��`ޫ� ~0Uk͝6���ܮ�<�#�씼���xz�L�������W�s|�[��a�ܢ4�6-�<��ʟZy�J��t�C��os:rwy<��#��M߀�7jU�cF���mklq#8���|�k�C�����[�n�N�	Jn�2�`�+�X��@�}��]+{Νlq�"*��gX��f���vgm1�7Nv}���� Qt�)���y�N9�m��t�E^Ʉ�LƉp&I��XyV&}޵�p���	ӻ�˶�<�@���<o�5¼y��^���5��
3�<DKO�GH�}n�xO�ź�}�r�l��oxQ����}9 }�c�Ɩ��I2kֵ��ǅ�D���-����Kx��8O'al݀q���{~�V�Y��^��*�"�:,�`��C�o��Z��X�wS�;��V��y=�,�VY�ק�X�'��S��{�@�I�[L�ei}]�p�ɝVk}�����������Yk���+I���~�Nq���/<��V�z�wN�^iA���
N�=�u&��Ӎ{�|�fVZ�-i���GRwJ�����O#��-�y����ߎ����)�鶌��4É�����t�E��E��p,f���E.��{2m����i�"��ݎη�,;���֌.{�2��W	2�m����� �����&�����&����A_�R�[�u�vc��;����qD/,����o��?c;��S���fբ��\�{�zK��]۷:�����<&�E膖p�ǳY)X������ZFt��(���vgeg6.�u܀v�F��:G��J+W4��X��p��j<�R�ǹ��{�Ŕ�E�tWw.O���Z�9��$�{����{���Iѝ�^_�{i��H�J%b���PL�ƃ���i�r�yzkM��ڑm�ݿH�7^j|�]�Y�n�,�9ΑiX�P�˸zǨ�n_%�m���}��3�`�ͽ�����\;�[����;B?(E�,P��I
�Y�J��y��<m��jhX@I�����s*��^!�f�F1+/�h�
z�J�H�]݊���{�lw�&%qN������б��Ƚ�\Fgs���Ȩ�Y`�
z�Gh颋"nx��su�ݵZ�����)���:s���UUw����LwK�k�¿9�l���t�����J���:`�mÇ����*���ڤ�>�:3Y�U��t�ՔR�v�U��t�LO4Ob��+��S/|&Z�k����r��k�	���o�DN���A����}/3�C�Y��]�����l�o,�g]j�Z�Ŕ�����w"���_�h���lg��x�U���s0���z�MwT��]�������f�CR���/�
X����9eZ�;�>壷x^�[�u QCS�պ���L2=dQ�oo�>�#W�j�Ց',�VJ��h�UݝE��q�U��\z��C�U>��b���y�E'��nh���^)��/�s�DT�7�/��W^W1���>��;�oOf���B����g��if];��jP��o[�W�>��边@�k}��/|Jܬ�����m����U�\�B����J�Ҋ,���ꇓ���P�s��a�m�M�Z�wwc�@�p�;������]Q�M��4=��:�W<�&#�9�]��uO9���Z��b�#]��;�ȴ����,�uE����zߞ����^���}��;��~|�<s��Y���(�,	v��ɥ��˩���3,e4�)�m����*w�p�{͖��`u�MԾ,��<}=38�Kx��!�΁!��J�s]Z����g����M^�i��C��|rL�J\��C���=�b��7�Ԩ}�e�̀l�/v[�U^n��ޝ��2�����7��t+�}�]�w���.�����+"�+����Vxa��3ޛ�wn�n�ϲۚ�,�̞4��x��;.��������1fwL	+��k�'��ߨ9|ۣk��稝zF'ۻ�l3���F]�:ѳ� SC���o�״�e_:ޏY�=�S;4�x҄J�u�y�;��`�Q7��
͏cٺu6�ƫ�|Ȯ=�ҷ�{P��m]�%�oR�غЦ8X���V�#��o�Q'�7M���Z��	֐���ݰi�V��;�
˜�:쩊���R��U��1T���B�D��5��?��8���k��D/���:Ƶ/GK��T>Լ�u�Bӡ�ʲ��\�g���Ͻ��2%P���{���4K8w��+:�$@�[җ���^g�}�0Mg���3f��j#���?@��"���mh�
��o�d�aqQ�>��OX�^�Z{ ��s��V^*_�؁��
&�oo{����<�;�,q����lPV�3�;��|_�a�_��V_���J"��o̷o�{���F�/L��՝�*��ʦu,�|;�ޤ�X��ә��.��nzp������vξܸ��Ǉ{��#ʍY�e�&���}�OKq8��s�Tu�OiDw��峯���p�{ҏ��q��C��:��͍kY�T*�-Kbϫ�Z:S�c��߼HA�]��vZ�9��K�ޝ���"�������Þb�,<l<QIih$�S�*���n�NL{�B��-������IW�ї=��a��<��|�v�l�����F�w�2�z���ˊl��zs���s쾴� ����[p��V8�N~�	�s�=����e���L�Lcs+5w����,�D[V��|���,�-Юe��Z
�4&���`l/hT��9��]�[Ud'e=�1�@�d���w1�	��ÛO������Z�"��|p�ŭm8𼕤��ݷV�Y�(j/�D'o�.�b|���Β(h���F��bp.��ܰ��A�̗��ؕ�6:�۝���c1�(+�/�wD�Z=���/�|����ަor�3�"IΒ�%$�S�z�ʹ%��X4=A�p���	Ձf���K�a��4���8��f�]�hG5@v�3z�ҩ���Q��n˽�P����ٽrT�Xf�˄M�����¬�og@���X��}.���o_V2q9ɤ���e>O4����j�w/z���]L�dg��6UB�k�y���Q,��N���bփ����{�=]�9+�s�F"��s�_qٰ�7_H=|��aon��(��E6𨃮��q�b4��^&CpY4{�\@-,ڙ�im2�87H���,����zLU�h�hX����)m��ܴ�0n<m�2>�|b�Z7
lY�����/G�,�4$������7��Yw9�R&j�J`�z�̮�5�/Ĭo	�21E�r����I1� ��w��ȗ�Y])8kwƛL��;�+�
��qo��6޽�RL�.��w�o���_)�i�Wѥ�9����:5����dl7jb���S��^�Z粴FjlwW�2:xw�W�#}Y�c��.&a[�3U��)�(� ߅6r^��jǻ3i�ٸV=����_7��Y8��֚M�=w	<n��?��m,oӊ����{�h���SY��.7���3n�^gCy�Pq� ��s�y8ne|�<�Q��v��n�N����==0�v��elی��_�Ϩ�;ym�z(`�����H��]�R�$%<{s<X��񼏹�m֡��|������+�C\����A�'\��a
2�Dp�����P��<3�*�[�4���ހ��u����j+�|��o�]�ͣYK@|�d��^�C�4[�b�w/t�+�S�V:�ܨ����5**�m�`�F.DN�]a 'kh̑�٣��o�X��V pW^�-���6&!�*=��ׂj�>9_���Q�1�B�Py̽s�ʜ�;�	�ϐ������)����x��sE��Y�/V�o���V��aȾ�iYv�*e7�^ˠ�un̏Z��CD2�t���M�7o����5&/R"�<��������)A���ze<�:�: �q�F��7��[��#v[�N�^H<]$�*��k�o(x��'��������#���y���;^Ѷp� ���5k$��]���wW�7�x3{ŔM�g� �=���x��v:=�N���u�.LGq+t��Yͼ�����*��M�n]��8h�������b��A�9�5�8��>���&Nse��*�ıڠ֢#R1DUb�����TQDURҪ ���"(�*,�[AQUE`#�$cTX�QG���1R-T+-�YX���(�DQ�,�ALZ�`��Acb�DeJ�Tb�,X1b*����T���b*"���AUQV�Q�X�ER�E"�1�PU�0TŢ
**������V*+��(��Z�UUQ�0c�"����1H1�����""�2*
��0
�"�#UQ���DF"*(���Ab(����("�(#b���QF1A��$p$TXVUDPU��Db1(�,QDEU���F(+E�Ab+EAbŶ��TV+�����H�֊��AQPQX�ATTE`�DA(�(�AAEAdUU`�DE���Db�۶R�[��Q�v�����d��k���N�[���&$嬨����6g�7�{6��?}<ho�w'_9����ֻ�z>G��:D�B�A�c8�g9o��_�^j�*��1vUxM�I�W���3��3�W���9�i$��^��w!��7�uf-,��KɁ�4��A�W:=��m����J6�s�5t�P��)%_t�_�
��U�T�XV}ϻl��&+��뽒��;��bJ|f�f��8�4J^6b�ʐ5�؎�����Z딻��y1�=��u�9�8���|A�Oh�`k�J,Ɖ��I��[ʱ3�kʸԬh{�/�R��
~@�8'�P֩W�O���1���(�>+����~q�9񘞥�Gh��X��M��MT�k�
.��c���@@�y���ROv����a귎��q��\L�Z3l�����N�*�|{���w���"���+�"\0����W^��O��O�:�Y�&����vT�.��<C3��z������q|ҼA�5Y��A��U�{
�{|a&t�\�jY<�jU�����)���.\���z{f�IG�ѥ(*N��:q�51c��{v۽���Ęl�͓�i�Z6�W�"+2���%oн��Yʜ�L%z++qQ�❍�k��nPR��P���p�2M*��e�@�3cOr�R����0�ū-a	��C���Uy��:d�<��G��
e�!����q��UG��=x���>�:ʗ���f�}�ԉ`�p�Nv	�]I�<'�,af`���|)�&z�=m}������S{�~Z���`�q������:юzƘs��ckz
ְt���K�Y�>�d��������m�Z	B��J���x�ώ�37ӱg�س-{r��AL�cl_�R�s�&{[ΫE�%�&����+�6qv�A���4�������K���O}31��*���ο8�V�7��ga�]$�҉]S1�"��c�t��U�/n������[{��ۭ�'�`k����bp\���A��ho8�\�9�o�]�����"hW��'���%�qg�A/.��=����ʄ_��	o-$5��z�q��g(���F�9vZ�a��g�?=v��+/>���q�O��(C�"!�tW���J'�N-��w����Hغ깡�궧uq��%��T`����,��ܾ�5�
�==U�{��"/���N����s�#�>�!��ƥ�\��2�R��׻�Q�n�$礪���a���������P�XjI�4%:���Xk`7@����;;�j��5�������!Pɪ�j<�iGݽ~Ϟ%�/,R�PV�5��`��x�R�lm��`�V�e�|d Qp1}�m��ս�;���~��K�ޱӛ�IY�h�kVK�f�ߠ��g�0�u�I���3Y�^�wMt�À~�5+кAo����cE�Ӳ%���/�oj�X�t����.V=*�������y�Ɉ��Mz����q�._�����;����c�ռ�g]jөT]K��	����+{p�7��[��e�V]&=BP���e�3�s0��;PϦ���~��w]���5q�xO��7��}�wM��"��(p!}Z�s��L��V�bu9C�:�<ro[��=�]Ӫ��}����o��+{~�rdX��XϢ*�S�AC�3~J(��ql��'/�Ϧ�?k-�e��z3����a�Ն��Թq�eUq�.����և���'R�2.�&�l�+��{�u��׽�\Y�l��ϝ��i�<,�.,2�������������(2w�������O7��<�5�^ �^�$IT��94�����39�ū:�X�����S<�����.��������pE�a����=��,���AY����M7�`76��\�JV���<�"6�'/b+Z�yg��L�suuʻ��P��z�.�u�)R��y7�q>B	�[Z�B�S�$O[nd2WhTi4��[ۇ�
¹��bl���q�8�ŗtnW�U���$r�V�^�z��8r�n]�U�?�Pk�o���w���zs�-�)�yQ(m���1�c_���=��L\|"��.ɖK.�3ӮY�rL�Si˝ʹIfR�V)6����i�|��,�����+"�]�^
��m���*u_�_�x`�v�=Ya�
�H��5��Qۅ�k�g��J�B�U���է螷Y��`�F.壦�˸q�����@�����uwy,vQь�}<�ЧVny�̳��wzj�IO�p������Ak�'�~���(�,����ST�����)���)ڢ��+y>�N2%���h�q�咴y�$�e�+�G[�;;k��"xL	��a�X��{�Jo��
0r�V���{7���aqQÿ.�k�)!<��i_bÅV���؇3��r�sL��d�K.���ݠ���^�3>�s�����u�Ӽfl��S������\��c/�1���T:�����h0{�5��)�9�����=�G ��q�n����>��u�	r�+%&qx��$�zS�� /��Dw���U,�-8���v��3�����g�Xo�rk2q[�$���LVg�u�j޻�gl�����.�7���(���r�;ON�� ��#'c5��&��sc..7Y-�;�knt� �D �"ũg
�Ux��3��s�UW��C�ɾ�8+pS�V�]��N,�L@򠖥�`�eϑZ:?6;4�Y�I��V.e�T�f���Ԍp�~X�2ߧx\CyY�<�NX#��Qi&��ilQ���U9��~���kgg�N��5zV�#ޝh�۝��5�cg�ϝ��}��F��iŌ�<r�o�`1)��(P�y}i��۹��V�:�J��X�����z\��d�q�]��G[sݹ��s�lǆ����~���!A�yƃ�r�Q�J��&���)����rS�jɚ���Ÿ�A�ß<������I2:��ghd6���Xt��7�wm?���7;��vz7�y����ӟ��џIbrɂ�����:R/�*WV*���Y���Z�Jeճ:�9�lK��B�Ev��(����R�wT�֒chz�Z�hR��9]����-�C�����-c\�U��h�
d��>��U����� ����v6�Y����}�;�2���m(ii��'�|1��s�t����v�|f'�g��"��k<����V�ùq��0�[�_�mm��[��Gy@F�=`��N�����;e(�v�i0k�!�oOӤ��2�f��yaL�kR����6l�T��M�v�ܻ���A��"u�y.��nM��yy�zn�O9�)ݔP���Cc������˽�V�6r��b`��Z�µ&Mu�y�_k�^���z���S�E��g����.G�䊹���<x�g}����W���K"����O%ר�mO	g�H�hcwեs�q�}S�r��]Os��9�^=�.��k�Vf,�ZU�k�Ԉ��N8�%E�ެvZ�[�k��L+O)*��\���{��ޮ�x��Q)�j4���8��f7�l����.��ܛ�{A�-��匈����	�f��XY��|�����5�e)+)���&��驒�H.�\���t�[�p�U����[��;�7�5p�h�-u8�t|ڬ����T��
T��!$s^���}N�\wə��x?�{Ҙ�^�6�7J��Ny�crv]���΋��o�rY�k�)r6Wm8��c�c��굧�OGCn{g�e��{���d�:kx� �f���:Q$��h�����u��/��	n���w�G<��|n+ίT���Y˕1`�(;-\��j{w5��(`�{G,B�U1X~�2��Vc�!�ΡŊ��oUs5�cns��K,��*4Ug/�w��a��-9fn4������-d�u����7C���ǂ��u:��2-�������තX���ۥ�Ѧy,���O�+Z��Uw�٬pU����/.�������*r�	`<�gϯ 4C����^~��k��]�w��B���u�3�0�U�N8)�1}"k3׽��^>sGݱ�J�w��mm�qٷ�{���ϻ���$Ts謰\	�-�Y��yQp��Bc�����o�o-^���S^�I����f��L�M��t��`��{!1��(�)�:�W:z�{_���xa�dXϲc�*z�7��^�\]{�L�_���U�m�!74`9=��[��<��������]���j9�X�t?Ki��c�����J����~�Vߗw7~^�0[�-����%��<�2�G1򘽪^�y1�R��R�.{<kh�e���7�;Ͻ�%>�|�f�������{l����>��;P�5�}Z'�ʻG���w����c��|�=�R��	�j�����.���kif_�P�:�<s�oWt�3���*��rVW��o�=���x���SE*E�LP��f%=�Smx�T'�#������ZN�u1.V������ :���qQ|�WQ/��P��\���pN�>]���[*���Q���]�{�7�'-�Wk��KP��O�o�m�se^)������+T��K��ݺ��Mʲ9�&��;0x���,��}2���&]���&"]����*l��{5����y�}Xi��r �0���M!Z굾�eq����+�o��x�������4��zsɋ���f�A��f�����a:G�����PL���y����U��kq����#�\{Zh<���~�ױz �^�$IT�M<NPtup�S�:���Z�5b���L�\�����4�[�����s蹬<fK�9�-�~t#��Ӿ񒻳���{_>ұ$^'
����6��Crƿ	Y�{�T��kQ�P�Ƅ�sӞ���{�;ckI��HZ�qV)8���>V=��Y��<�>n`F䬂�qeϺP��QSxMW^f�+�����:����"�[G�y��UQ���ъ���J��˹��=Ԥ��{OSfd>�E�%���]Á����Mm��#��^��W�z0���+nc̈́�cޓ������IM�XV$�����e�v���G:[PQ�K!��=�;��OgR�@9�$x߹��r�Z��~���s	W�p�,9���}o.��;�!</�VuuYH�!��ެ�v�gx�u�R�7[���I#s<d�f�1T�.���m��}�rv�6���\@fb�7�r����Q��l�e9�,�5�-�{�"�Y}���u�5X/�	��V�P��9.��Ԣ|7d��މ�ѦYJ�Dlrޏy^�Y��_�.*8t8�����J��v
 Ǩ�2���w/Vw�m64Ǧ�̪�J�,2(v�r�����ؿ�x���.����j�s�2[�$�ܵ+���Ǎ�o�n�o�Vc�0UC�_�
���z�Q`�q;�望�i�������_S�D�:�.W�d�Ãp�{*���ʤ��G�{Y뻰�7\v�>�Kt fN�ѱo�z�Rjڜ�ϋ��v�͍k"Ȅ�*��N��.T_|)W��w�-v�f����m�3�g޻��Ƅ򚑏&�(o,9�*rϣ��#�-/xՊ�*��v'����7��Ԫ��Zg˚�+n�:ї=��a��<��|�v�l����թC��A��?_=ܜ�,@�!�IF�tї֙�����C�"	9�_y{|�3W³���3��G��}��7,�6;])~���\3�k9n��s�	W��}�}��*���ߜk8g-kmnLy�*�i�I�b���_�+�O]�.���-$��42����s'����c����eSh!Z�fV��w]�5Uޞ\L#�E��}{��Ş/��j�GYE��E��0Q%�B��xx��<��C����Ӟr�nw�x��#q�w2�{����k�[�Q˛�J�:˗����h�So&	���Ӂ�6�d�',�J^�%}�Du�㢖%�]꠼祌�Rt�ൌ�o4"2ZX�۾d�;��]�\D��IK��yv����%!f�9"���?b}�$��[�/>ѫ*Zf.�H���&cDۂ�&�`��sk�'L?����<s�E�0R�vvQg7¢Oh�_k�G�g���Ptyǈᘞ��2�y�$���s�����ŕ֍��鉂����T��5����z�*�;\}B��l]�6�/C5��ӣ���S�}r:�r�~嵇�I^>K�꧗�^���h�W5��63���Ix�~)��y[���M(=|v����qP7J�78�+�1r�]N`OH�Ӻ�
��mg����5�����+ˋ�S����sR��}��/'�QaЇ��pX�}~�O�ѱ���/͞ޙ�ʟL��G zjD�m�-9�'��6���,��=~5�D��X�՜����k\������.��9����4ҷ����b2�i�>Nv6��U���5]ה���/P1i��*�2y�Z�7Q��9�]tz�Ĝs�b�9��A�-�-ce��4�r�Pt�T����3@Ol5x�Z�eeD��qK���4����)*�y���1r�]�1k('��^j� ��rQ�;��!yܬ���,�)�{��tA��(��Y���Jf����]Ī���>���5��k�Fe�i&��Ff���� GI/M3\���N��8��WV͢ڠ����<�:=T�l>R_f��-u|�t�l�50G�i���\�*+*�H����vfR�,%�youA�T���$�yI�h�˔����g��U�a���c�&�?�9�n�@��A���]2����آ��mX�\�Vd$�K�z��8�tzҠ%h�2��},�Y�`.�ui�p�Lf���a$V5ϵ�:Z�q,��*�sx�:�ص�7�̵��Q_M�lܭs&\��z(F+�ź�H
��dh�)��՗O��VF��R��pn��JĴ����S�'�}O���4��l�c��=/ukV+l-�m��1�V�kͼh5M�{�u��7�iA���[�y��#Cw7��˽��b�_!)�컽�b�Q���P�I����0̬E��R83{����\��+/�����k3�M7����X���<���V��D�d�/3���F�Xf����<�s3R������3:�}1=��2s���ҹ+#�I͓&/�tˤe:��5Zj���A(�GF��C�������?`���9�Q�B/�3w���\�3ѡ����"��V�L�M �kKT�׽�K����4,S�az��V������ (,ް&�Ƶ`�ʕ�]̓zDy�F�B���N�*cʔs �����o}krڄB�mu�{QVNGxV����.c�)�=�d�΃�̤Kѯ{�Z侹�G�]��3x`~]���;2�
l{O���u��'rZ��J8m�St����Ax�dvS����Ly�Wn�N�T����O n��َ���{C���z0��$oZ�S:V]+�n4�����k\�Vx`9kmG\�<�Mq��8h}2�!ihv�n5p$h����|{/1�ܿ���/r�x�i�h�A�W�K:�,��\1_](�]V£i}���G�_$$�MК�[]�:��=W3��{e ��b�U�v�_<�Zhd���s����pW`u6���7C��jO���ȗ��pv(� Yo:U��9�J�,c�( B,5�֬�����o�w[�ɘ<�V�������F*��=y �7r��uf���NK��ۖ}4_z������7iӰ�8�s-��Co^_�jV-:&���r�u]�]�m� \w4�QNkm���^�+z;]8i�r��2��!��q���H���F����UC�vM(Cu}Ne�9�:�_���t���Rw��������Y7����f�'a�����ׯ߾/�����v\h��TDE��"+���_��"**�X1E�[h���*,F	R�cQTEUb�"�1*ԬEE1eX��)U�*�"�Ddb��j�0UFE��TUQb�F0F*�25���dUQ����Z#UTE�`���*"�Z�.,��Tb�"�*V��EQb1
"������X�*���DXᢨ�ТȊ�Ŋ��)��"����Z��U1j(�TQQ`��b���UTTU�b�0V*5�QP��F*+Z(�H��������**�(�6��F"1TUH�Ҫ���
���Z$UPUD(�TUATY���P�
���e9Z3�-v2i2N�p�?Wns����<��X/!s#O��'�K���W�b�����U�uq@$�8��O4��P��^�ע�I��#��r�v��!����،3��Y��u:vU	���{�7y՝M��N��Y�Q.%���q��qv��v�7ǘ]��s��TeH_x{��?&�A�^{�����ŏ3n�C�(��T�kȾ(=���
�ǗJ�(+��M�uS>k��^�����=S�QKR�������-+�P�r������<�)V����.�A�	�츖��ְK˅�+�{�(e�ʄJGt���7!����{&��koX�'զ�\��v��+q�3��e��U�N8)�9�����J��[�� YW�N�͚�$C2a4=c�w�Ҝ���D,f�E���3s����*0���G��l^�������]վ'ua0{H�����H�el\]ߥ���T��@t�������9������~�,(6v0q�,���7���,�|:�/L
���ZgG���ϟUO�J�X�X&�s~����l�"�Ac��1�i{��B��/}e�x+������~o�5��3,�o��l�ƨ�]�U��3�3��"�Мή��v7Ӓ�b+�w|���|`Rf��K/:���;���e��#��4�x�o$ט#o�%���%�k��[
�D+�<*��G8��a��zbq�*�m�yg�AY� y��pI�}�~�ho��V����$�#�uA�s)�uKy�uS�ɑW��&)�z$�r�=#ʅ�r�F�ڜK ��fS����z�	��꘡�gN�F�M�V�8�����d`�
��q�gUij���.�v�e�����r�Υ�Z��3ݠ],s�{�w�KH?��\UXt_]�5��[J"�����bW�{J(��ȿ]��x��1��5������F �[�{`��٘�,
�L��r7�1� c���7�e�̺��S����۾���=��G)Esϲb��k6
�ن�g��r��#�.-3W*�Mu���;����/��<��[�P�.����ƽ��kb$M�\�Z
a�M`�ϯ����{�㒅C/)�,?[#N|����]�g"��.����,���+y{*�ӧ��Ǽ�@� �5�X�9<�L����/Η �P�A�&�+����XGv5aG�/޼�\���ΦrnY<l�$/��⑑u��|��jE�h���xIYcE'�f�l��Z;�gJ��W�*:ܷt��%[}�p�ͩG���@�*�֖��ST{�����e����+[�C�s�g�t��Gs�}�]�	�ɔaO��Wsp���t�ܣz��K1���w��Z�G�T�`� �n�\�8 ���r��9[��wpS3��*��3�˳�H�őؑg|�S<v���<\ų��������ٖ�ow��u���W�1��Qk�	,��F�'Z6}>�@T
������o����U���Ɣ�znV��3��ϻ����pXRP`땍jQ���U�����Nj
�cN᱒�����c�y�������fۼ%lC�яO���KW������I�oJ�{W}��&�x�>���Q��9��Cc��M�f�|x��U����N+>9�#�zz����w����m<N;��k��~�c�f��K|d��X\u��P�k<`�{l��b�.�yuS<|^96jcP�Ov�骯V�^W���n�o�c�2�J�AB���5xa�;���G�b����?��O�4�t���D�9���Y)0�n"�D�>2�Z<�����5���e����M��SWv�l�Ҋ�S����v�lkX�(H�(�'<b��]y�*�+`[���.�����v����8�Byg�ia�w�䡼�瘩�<TDi�դ�.e��0�#
F��M�qnu��]ZD]��˪��Sf��UgU���t�ݡz��m�b����w�V~�\/��oI+�j�0Б�fT��k����/�b�µ�Hk�ǸZo�#�}�ۃ��@�ZB��PsB-��g�r�] e�77��sf�rd��v|��Ѯg��.j���G��FX۝	�y�P���$]m8�^�zO<�v�b��^�@���p%�L(s�2��8����+nqP�8I��æ��S���'ݍ���~�Y;g0<�a�Q<�$�_XB���q��g-�<�`�[ԯ�2�1׻u��m���P�X�L]�ɐ�:&F�Ri]S#�|��!��#*y�>u�17�q�0���<�^L�]�8�Z3�,NX�P��IWJE�eJ�(�c/%�[G�}�������nfOhJˊ�Ev��(����R�˰�)$̍��;���:߇s�nU�|�
�S���^	�qp�8=�� ��� ,��L��GH�=��2����^��o����"����o��4��V���Z�<�*����<G��<��W��5�i�)�{��X�mu��mq��'3�yf�SI�]x��������L-���'�˻�i�Q�{�yk�p�r޹��w/a���[X}%xd�K�痃�������Y]�#:�Q׬ܡ�m����a���L����h|"��w�j���x3�%p̙Yo�/GڒukVX�$��"Q@�3����v����C��a§�$x��!қ��P0w���ccM{���(�\Q����6H4n2g%a 5;��RGt8��M�G)�W��]m�O�X�X*L��:��y�ܞz�fт�+6Z蕏C,b�fZ��;w��{b�o����]����9[L���9S�C�w��ك�+-y_�q�T���f�=�(��q;%�Q�W��)Ď=5"Y6���5'�9ƽ�XY��w������z6�V�44�JX�C^�iXzj�����[N�wޛ�n����G�s3."�d����[�|����lƸ�.!�H�j�˱�N�\�&f�	،.8��#�c�tc{9���,��s��2�t�"�},�4�.F����k��|y�K�wa��f
��ǳ�**.s�ևA]�+�yN(�^Y룦�ơ��3a� k�(���cY����&��W�,g��	Z�_Z���zo�x �+9zz�!gʘ�L�@�:E��Z��$}��J�"��k}��B��<�Kb�P�Y/.��=Z�p\�E�'�I�&^4Q��]�;�i����jW�P�UC��5pv���ј%a���U�N8)�5�ٻ������tIϷ���ӷ�H��ܰtGF�uz�35['3{+��y
���ٳ채7�wb�����ţ�Gy�v�˲��������;�B㳅'!ã���n	�Q����T,��}�H]�}Z21�2����6�&Q,�3{e��:�ڢ4��&�X+�����A���Hַ�@u.>��#�����b�Vt]�״�0l5,������f�"�^_���C�z��^�!%�#0�//�������ZZ�PY��2,,���676��p�.�Q��T>Ճ�L�`�y6�On`��o7y������:�5�C1����E�	��w6�f�ǂ����Ʒ;�&�f��O��q���X<&�Gox���ǥ{͊�W�̡�\��D�w)}U���6��]E�sջ&�w�g()x��#ʮ�+�����N%[L����#����>���7+���^��|��W�UHكY��-�,)C��`�+D�iL��x���3�r�:�S���渗�����1�>���=rc�}�rpōWѪa�����+�k6�h��%�={���m09�N_463{g��>�4����#eq� %� ��Ǫ*�\�1/?���y�螯>��똟�k3`�ȱ���ٓ	F��O�ǼO���f*���W�w��~�LSz���ށa�Bh��Hcs*�5��ܫ�-]b�L�G��̌�z�����J��saI���Y����4�3:�t��6փ�����4�������2O;ڠfp�ȶ�7���b=*�#��c��B�]X��ȕΒ�t=�����u�skDC�<��n�r�\Ж�l�D�H>f��9��K��|��^|�iy�
�/즔��diϖWb��2.kOL�9��M�3�nRU��s�s�T�� �:�R�
g�eD�~t`�-ޕ{��<�t��=!�ɹ�&o���iƌ�ݳ��Ɇ͒F����Z�Su�]�^�i���(����-Ʀ"��'+5*�ͿVw���� Tta��va��H�dv+��˪,�*,n��;M:׳{e(f���Y��ǁ%aʄ+�1���-p�%���˸q�>��
�P��}U�<6����y���X(آ����)�����F�qzl���ª�ᬑײ�7�إ�7�����p ٯQ��8\��φ}7h�.>2��%y�$��̷�xG[��W�s�ٓ;<���w[��?hBx*��"�ōϼ^jc��]�C�,X+��[�vsE�s�C;|gI��>���6V	���K|d�^u��u��Q��lPV�1��L��!�Wg���ʬ��s�I���N�W��o�XmU��T ̔{�4"a�;�ԓ��4��\�>X/>RN�Te���*�+c�WJ�K���{��"�X2��jda��+���.u2�&q�z�z����=�=�����v�6��Lo��k�o/��MX=�7�	�㺼'�iu��})/%�R���P�N��8&C�7����y�G=7��{���[��0����f���I�V�k>��3���q��Q���?{������H�+�Ҋ✄S��Ƈ�?��B`@�-����K�U��oK��������3*U��D�	Ƅ�ɴ�����Vxy���?+��]W�Jt�E�s=Y��T۠��Y�PF=���� �\��+n�}:і'�:,39�hT��w�����_�7�|�ҵO��h��h�|�50P�����.�O(�P�x��Y�ߵ�V �-��lN��w�}����%��&Y0�\�h�������(=9n����X�eMI�1�N��4�q�9,�;�4�^U�+XqK[��!ÀL������V*�J��٥i9M��%}�������m��>ZYqd�����i�(��%	���*)%C�"��6��j��XX�MY���y��`��KG?���q�0N�i ���탎Q#A�)y[˰��v�� ذ:��v�
>62d�)�&�Z�=��8�����pE</��z��ĺ2%�T���5v�5��f5R�!�H��Z��n�c���V���[���W�7���|8�]��*��,ѩ�Tk7����n�twu
\�˽<�����$���Ԝ4�j��˅��u��w<����]gz ]cD��
d���qa
���o75 ��skŭW�X���L�>�=��a��yx`.�����^��^�ި����� 3Գ��+��ਭmt�u�ּV�
I��\�y�Q*8��Wt��<��������~S��^[�'����;��"���L:���ಏ�&����n��E���w�Aq�8@+ltX)���P�����Z���o�XUf�]��h�3�T����ۏ�}�w��;+]76�=�0������9x�r� aq=^�ك��e�%Nb�
"����68�b���N�[����N$^�"S�ȁ9� jOP�VjIA��{r`�hu<NU���a��Ֆ�ZhCdu'b��w�i�oMC5W����w�y��I�^�E^��'����7QX^���dz����5�f�����m.|��N���vi�ʮs/��(�{���,͚�Y�V���
e�Ob,���NR�o��` �au ����	��A�1�)3����]OM�c]��л��ۙ�pR�Ѫާ�,J�5�̓U��X����L��ZJnF�r�C�&�;�z���.Ŏ�@�a���P%L,v�Z؉r����)�fȑq#2v�}��!�-�]�2h㼱6R������s7�p�z����離�R�Zߞe�@�:Q+�f5�K#�?o�õ�Od�l�ø�|����r�8zJ�^���Y���m
�㢭MNok�pj��&6�wf#䠩Ze�C���+���/|�:�	yp�Ev�x����*=�x%���Ogv�� ��$'CM(x�۸zǫ5{Q��u�2+0����o���哱���j�7_L��h��3�"�xB�=��_���r���[��r�V���ޔ�y[�=�U��b���C��9��2ۇ��#(9.��.���[7�%A�Y���<}b�nRn����XKD�N���	���5,�l�¿��@pE>�E���� ���Z�7�|&��O���b�#���rEߌd���f� >�����`���Y��yi�ڇ~�V��(lHN!t�G����N�=u>X�l��C��
�x�z�z{͊�C��(d�1��=]��y��+�w�.���[ۦ�Q�XN�Ƣ�5�#��r�Y`�ڜK>���NfxGa�}+}���wIo-[�-��^�������_�8�c2�=�nכ{\���OVg�Eo���`2���f�F���捚lK#{�7��}%�!��9��j�`;v���*.��[�� wPoS2.�	f\�G�Y*���48.u�8d�up�]����o���0F'l¥ /%/�J��yq���g��-��{I@�z�,�"E�jUm���ּ]r����������I�nCF���L"s���=+�J��D�U��ٛ��_&7�t�8E����չ;�Q�S�1�L�b>�兊KR)2�w&F���}Ǻ�<���H-C.�7M%ڱ�Wfn��[^��׼���t��>H��kb�8v{]�9N+��z�Jc��0\<�8��(�^ӧ���䴍��m�ʗUrH����������|9Q���C̅��r���X*�h.�t�ӡ4Y;@.����v]�a��f�l�q�Beʎs��+��\������t:\Ka%SU	�e!�v�cf�ۺp�!��*�X-��{+X���Y��� !�&2+��җ�}�A��*ҞK���ԩ[���_p7�_܉bLd������ut��=�V��.����h�
VT�b���zl�|!��L��o�Xi]�Ωp�sU����ӎ�0��Ղ5�����{,h=����
r���ynD:ώu��}0�d�|c�H�̘l�]�:����V�63�:�87[2;�Pa70r0��QY�y)�m�Ӹ]e�{9�u+����1V��w%��s��4$���wHj!n����D�NP��v3s|�@Y�<;̑�H�u��y��&��[}�py�5�:��i� ��c��y�P\�;���sj60�)�Z��Y�>ұ�ΥL���q��opc�=����K�_3���	�5ثF:��0\�O��<���1.��x�N)r�z�qʾ�V6�>��;���7�B6d�c�3����y��XNS<�Կ��!]X�;u��M#�o�)}���&	֮�7�f���Sj��w�w�����㬂�W��m�tt��tvgwd�v��n��R��z7m�,�n4���*e��������F�D7��iȅmM�Yj:w���.us�-�T4<�/D��}qXCC���fLv�U����,�)�{}��gt�\Z���P��C�L�m��r�G�)�Z���Y�P"o3��mᛔ��Or�O�֮��}b&���c.�r.�f�[#�������h��9�1H���&�;�@m2��e@V���L��`�U�������O���fǝԫ�Fv�_7����7���0������Y���$B��*�O��J鳈�ۭ�rq�����2X]�u���8.�]����k� �c�i���p�4�YT/.܋A�n7�V^�QxL|9[�t�m�%�NLj��
X\N�|���} ��(����0R}H��`�>�$zd�"B��=���A�E�-b�_֪�UH��Q�TQV#dEb*��A��hڵ��UPF ֨ƶV6���TV\\V��e�Dm���b�DDT�UjYkJ"*��#1ZщD��DE,[km��ب�������$T�A�EQb*��eb�E��F�UF��a�V
aR�Z�mj�U+DÌQ�QTkm�(�"�֢�lX�Z�kX-�m*
)R�0F*5���*#��J�2���,m*V���J�BZPV*(��5+Z�jUQAm��(��*"���8h�j"%�cm[J��b(�*�UF1TiKKU��R���)j#-�,X�R ���F6�
�DVҖ�-B�5�Rڊ��FV���(ԫ����>Ћ�K�km'+Vqά�W���v�]�z=�������,}se�����7!j<8�Vv��bA>��t8e�NpV[#i:媭\��{?��7|Q߅�.,���hr�!V�pҙi���F��^C*��s�T���;�v��Nǎvk�;���t�#���Z=�}>EV����.j%�/z������){�Mgm��ږ���1"N�{���C�vo��p����t��G�bKG�M�e<��{�I�ʧ�u���u^��<��9(��옄<տ��0��wk�`\��=6˺�;+&s��H�u�#�PP�uE��? �S��4og�y��^��v�e%/#�b����N�No�@�&��R��
f_�M(�L��������x�4_��h���F�z�n�'���u�����>�M4^8��9���XʉB��r�5�J������,s��U�ug���Y����2�dQ$kK��I��T-�R,��\��U�r������f��<�u����j���pU����f���4Y�v]Qf�_E�g�3����{_K��>�z�Y��`IH�~�1���-uO��F�߄�Fϴ�L2�+���W���j�W:�6>�Ggw��QS.���-P�~'1����vj��u��!2��[�S�gue���nخ��V'#Z���˅�#�ŔӦ��Vb�kxM��X�m�tw���L���6�
��F�YW�:�9�'�1�o�m�ս��$ʾb[�wKIk���%����[.V>ܻ���^
��h�1�f�.s�wk L5㪥�</�-����qD��@U�;��ne�)��{絻�]X]N�9�0��Dp���綥��6��T\�~�[5_���ri3yCY9��~{7��b{����
�c�ji�v���+u,j���"��7l��ؠ�p�"�U�yGo��犲ӭ���=^��L����ZwJ���mLP�W�P7[�}�ݾOk�qI�e<>���J(�;��S���t���D�:�X�{�a��J=�`|ev�W��w+}���qٽ+m��ݓB�S$��1���(��!0-���ֳ�2P��Ef�r�]�Y&��%���*��J��.]���D�N4'�Ԍ����J�1S�)f�j�]�s�����+�]K�-�[�J���v�ϝ˚�%m�=�֌��谗ewG������Ҙ��s��|r|.ּ�{~wh�%�L�C�WRg~v�j�����t�JxVs�8��W��k�����'�:^c�to�|�i?Y+��8N�a�Wb~����4�4ev�^F�dk9���M�I��%r��Azv;����CGdk ���)f��s����SՔ�A�x�Κ}�o�83��v�B+��e�
������O>H���Y����e����'H��Р��A�a���MT�1�,i�;pJ���T/V*b�p��0T6&< �:�`0ENR�"Y�_p|w�ͼr�a�zάϖ�2)W,>�+���kFIbr���P��I]���.v+���s��~�Ŵ=Y1�f�u�k�`���i+����H�;=�����ȳ1l��?tW{����Z������Z�)&����33�e��a*�1�q=$���9�^���wws���OjG yV޵�&p��.X��sƝ�:�VϷ�^;U�Q����m��ʹ�Fl��/Գ���KV׬�kk���gZ��i�I�\|���c���zh�\#��������k>j�c�[K==l�h�4�Za��[X}t�ᒒ�ھR����hٺ�z�߽v��-!�m��9�<�-�ζǹ=�/n��Aγ��W�r������);��ǳ���j��U�a�����N^�\����臨`�u\�͠{�����^���ߎ��)�3h�z!�w{����'ۧ,��Zy�6�H�$ɯ�����F��]�{���Bʚ^w1D_}9������:�{��-�w�MƑ;�y������z'�>�	��W�e�y8�wF���Ӡ�US�u�.����m�^P�EjGԟ��|U�@k��N$q�Ϧ�"ӝ�x��hk���^�yV�͍/N�.=P��â
߆��#�;�CeT��i�`=5�	،�$�%w�.������p����i���s�G�=vc�N~k[k4��]���� Kd��/�:'u�=��Ϸ���b0�s�g�V���AL��h���A�\��WH#�٩;��W�!��Ax���~�|+�Q�1 ^�\��,	�y�^z�y���>xi��BvzYfVl��̾��{$N>�\"PP�ƃ��:mc��ܼ�/N�Vr��LB��1K2�Xٸ�4�T���t�>UP;	��}1��os���_�:�K˅����|���
�ڵ�߮�T���"
z�����\e�wߩab��7#}��}��|�Cp�|��z����^��L�l9t!ەDB�'غ�巗r!cٷ�xwW�1��a��u�䥙-`svt���ٝj��pSԲ;Go�f�7��Q�^G��+b��w�Ԏ�׌ў��S�x�ދ�<}��z�7^�ڦY�3���z.y2�AȲp;ם��[�zC@����Ɣ��s2+�����iȩ�hf��rQ������@��n\9.���C�����7��6�v,�#�w7�c>�g9bƔS�λ�<�pXW���u`�B0?�&?	B
��ڄ7�u �:��x������{�Kԙ2����U������9�,��/|��csn=��^ʚ��'k�t�7���� _g]X���E�SF��dF__��%�ϼ�2��/�`�i��b�n�m�og(7�1g����Z�c��2��F�R�ى˳���I�h���}�o^h�A�S�'��Wh�٫� ����C���K��i�Z�T�V���J�=Ov6��پ��g�����G�'����t-��3芭�R���}mK�|�]/^��+�jS�(�Ǹ�6\���l=�3e��L��\���E��v�1/�s�������TF�ݶV|��SW�R��d��5�
D��.g��b)s#V;�����GD3�e�X�v^v�����ӯ
���¬��o�"�v��Gu�vsw�;�$\�ݠY� ��yB���SJX~�F��׭�v���<՝/f��C3z�"U�x{��=��ڵ��)^�v"*�/.���̥��TW��̐�ݼ�આ�p�Ssy�T�\+U�X�ؑf�?���u�8��A�o@����6�e�����r���.Z6޺�_����F&��R�#�k���y���lݽT�z�b�պ��W�+�{�D�@�5��\� ��eD���k�nP��^L��ڽ;���m�:e�����P�#R����K6�F���H����u�]�^�,�{QN��}�4+�-�ή������dA�T�8C���c�}�p�����S{c��{����c˓��0;��<;-f}�0$�IP�rf0\E�$�t�˸q���}�՛�|�s+;��tm�0ϏD5�}{�I�~t%��'��>�m�,0\Vג�-[W��.��׬5��;��c�h�ɨ�L�e��x<�m����0�~w	!�<Fl�\nqJ>���p�mx��	�&	�h�x���ڑxf�Ⴚ���:y���߉s���zm�����LG�({�7�͛+�0&:%�0�V��*�.�5��$z��oxR�=�t]� �z{>�s��������/�u{��ZwJ���)�P�Uoޭ�쮓:�z'l~����Ѐ���(�;��b�̇˥�^3�|'�B7Y�6;iZ~�FLuCk�Iڳ)'|��2L�*��J��FVФ1s��;[�M�=�#u���7ֲ�S�nb�K�j=w>��x���{��ܞ��s��ۃS_�kM5�^�,�@�=�Иq�
�(��o3�%�(.k��#߄���o\)!A�h0[S��w3WW]�zt��-��fS�[�h�P�w��z�]�S���~[�FlkB\�=/���V�S��۠|�Q'�+j�Eqz.]���ȑ�P���2 �;���Cyaܿz޻�C�b-񳱓u�כ��e�}D��c���Ӑ�"+��t�2�T��[p�x	֌���7��t=Ҍ�}��:~Xg��3�<�v�g��v�Y���/�n��C�^�^��AS�xd~�Ͻ���V8�s����z\����`�d�c醉�'���H~Y}�h��b��H}�߼Ps度��s�J����z�R��}�!�,(w醑�ғK&�s���̳룎W\j���K����=J��4&�+д���/&P���Z2K������fx�@�-����b���󵶱%���)N�`U3���v��>�v���SC�H�O?E{c%��g�=<y��l�\���ܿ7\|˸�]V��}��Ayހ�a}'�y�\�[���B�Լ {ȅ�\skƢЅq�X���m&ii𭤞�iJn+���a���xʆ���e��T!}�m��ؕ�ʰP<�B����MK���۶o:����8�K56��ɶ�����LWRεx ���#����r�i�B۸n^Y���A���۳ec�Y��>]��a�<���)��lq�����g
ί���<G����Gh�W�C��>�����5�ּii�i3�h��9:C���Gy�8�-����>j�y�i^[�'���v���"���10]�P�|jʹ�'���x�vu��'���� ϫltY�9�=�Bҿ�;��hi츁�W�}�����|�zw@	�PS�*��4;H���	/��f&�v�v������VרkV��WWn6�fe�yFl�X)x�m���Aqu�.�G<�D��#�s�K��[��v^}���Ք��i�NW���P�:�7����u&�=w�`i�=5��;����n�jn��3��#o�h��ӱ��kY�OZ/%�,��\���&�H腂�����P�fXE]r�*�Q����/S�����!��yx�p���B����}��=z�c��>�'
C��!����uZ�է��b{�{�����ş<4ͻ�iN�%�y��+�s~��T:�P\E�A�u�X��/;�Ӏ�����bp\��7Lg2wL�u�n�����9��9�C�{f3ke�x�m�F��85��iV|Dp��@O��C��&l�YOJV<�оe�v�4'ú��.����{��q��W�#�,��˛��usX��S�{Gh8�Wܷ{.���7{,f)�<h��R���uo�:;g����4:R-+�P�Ϯ�� K���[��Z�u���԰�*UW]9]矣�;���dX��P�i!CY�I���7���\&���dz'��/eǵ�t)�ʩ��oi�/J����O��C���З»��n�D�m�H"�ה0��:]���x����G@x��+,
z�Gh퀬�f�A��3�t��*b���_(��9�g���c��g�=3�hn��<��s��,,���7��|p�-�Ǆ�g�ݏ�{��>��w��
9-'������u�^�,{<�4�E�q�ZZ����X�)��#l����ә��+�m�9��9~�2#�}~3�d{<�2��-ֶ��iו	���{�����^��uFaӑ]�ǔ��ƵD�qYN,�pjq,���o��1��]�����i��bj=�բz������c���)m�a:�P`�Z%�d�ʲ��z�d�Վ��}������g���}7���쇽Yh�`.5�eVڙJ���l~��ua��Zpk[�V�ո����wh��%�}4�{�)�f������q4�,�����B��쭝�(�Ų�2��_�qz��a{�ٵ|��zZ�8�d�Se]n�V|с��2��/�+$YS�qֶ��T�-��`�������;�܍*�����I��M�a�\�>N_4<6
�����6�[�	d������Zs�i�)U\^]Q`u�ecC�M^�J+ϲb��k3`�Ȱ6a��ףъ��b��􍦵@������e̼we����(�-�<~/8�U��}��%�&xlu�w�<��<'�����5ɥ��]L��L�M)�?[#N:��.�s�g��[�I�N<�mckŘ>~��9��ņ���Aʉe.k�P�z�ʈz��v�)-�=o��)#��<�|�ߏO�U1q���p\�w&Y,�$���,n�]c�4܃����m����S�E�������?��'���0�̻0�)��^8m'cd��R�S����+�ksա�Qզ���g��J���
ę�Qk�	-6&]�M���V��T��폗�+�؀�ÇCq��]�K�F3��I󂂒X`�V5�dmeК36�utFNGw�j���AvX�C�E�ष�<3��=����@�����("K���հs�:8��/�����C��Q����x��*9�@o[��VtT_d���-� ���j�}���c�FQ�\� �۔v����<lvٙ�\�ˣkr=���(1L��^�z��r�V2H�O<Jd�ݍ��=T;n�tm]���J�N�f��-]�)�	B����)�{(g{W{�i@[�Q�R{����*�Y&I˄G5{�����O��J�\�b�39��V�q�:���t$�]㹻!r{���c�
33$JY�sb�/F��7H5��ϑ���u�Pe�T-Ka��m�A�&Q]c��|�5bE�_��,fn;s	�]��G�N`��q�n�tOn�?��+�+�ٸ/�|y�(A���=6�;2(OS*�}ʔ�ɺi)6_.���.�p�3i�3B��-}�:��dZ�ԣ9��7�a��d|d�¸-O��βw���'7���C��WeR*>ջL-a�M���E�j�*pP`#:5s=0U�Y<{�糷-y=��JӬ��/��t�A]U*w��Α�^���V��1p�ox��.�v�9Y�#��X�GY6���e�SRm`d7r�2������ॖ5*3z!9��3	�
�(_1&�{��{)�>��6��ғ!>��9��Z�s��ڽ�ݠ��G���GM�Y�I�|�+A1HuA;:��&�ӾT6��+3��X���ϲU�%�L�!��ѷ�Ow6���A�3J��Uv�P��Y܇H��x۬���w&�
WP���U2�'���G���"�/`�%%�图ݨuCqE^�u-�d��}�+���q��T���kW'���okQy�}��ƺs�&���d�em����vf|rA��El�?�b�v�*�k����(��/iF����,\޿�۔ر�p��2�'><������i�g5���)l5p)|,�gv�J��3��o(jnkZrtrZ�ɮhIŤ������þ�R��p
z�Z���=x�PeDU�Ӽre�vy��7)�î�xD�@!�@ۤ��:WSnc̼�4�8�ٴ�)3���͵oxd鈞�n��om��	!Ӊ���Y���gPY:�n�{j����1SzA8�skfڀ����v&Σu7t �K+ 4gp'�Y�p��'h�r��E�ǘ����ޚ5��F������M�z�#��
n['$��=��Ӥ���7�vrB��S�ќ+"�8��톯��l�߷A���I��1B�����X7���Ύ���:��������
��+���5��ܧW똫��ƽ�W���6��������'&lI�!bշ�ek������8��`q�Z�B����I�Fx���ɸyn���'W*8U �d33�}��nn[�Ń�z�wk~��B�8Δ�!�O}��c�`�7�4�knk��>�1q����V+K*,���)�b�,U�1�D`�+Z��UEڕ�Ҳ�1�iA`��%�
�Jֈ�(���*(����J�Ҫ�-mk-��p��QU-��ҭQ��ڌ0�0��KiF�l���EQ�-*"�KU+Z�ѵ��j��)Zֶ��kb��DTkE��h�Qm�kBڍ�T���+
�
�Ŭ���*V�RѪ�F�JѸ�UYZ�*Em�kUe�1�������**ň6����[Z�h��
[hԶ(��ѰL8Ll�h�Eb+if�m+�W�1�J�Z1�V�U����j���ج[jV��Q�)kJ��AZR��D�Ҙp�h�
�ZZ���*�E��Kj
VԪ�Bg�ctv����ny�^W��eu
8��S>��a�=Xiz��t=:jq�0k<F�4�y��K�b�7�H�� ͘��F��7�m�;$����Pͯ��O�0Mg������������n�2DTh;ؗ�����_xz�g�=�Y���S���;�Ҩ��+u,j��9d�[R�XN�{�6����<�/m���b��p�~��Y~��a�XX`LtK�'6վSʃW�CҢ�tށ�r�����W�Ԛ���NfC�Kz�Lîe�G���l��� Xܿ_o��7�j�^7US2��|*{��索��!0-���֩���`.�o���Θ�}IPҾ'	�2�jc�+GJ~ltwr$pN4'�Ԍ��;��h#�췣*�wӱ��+\db�,o�����5�M-��h�\^}t�3���^V�#�%R����x(WO+B��>g���|s�kfR=��(�4K��B�<����',5�`�f�g]{����#��������x���,�na�y�I���W�~R�I�_L9w�����A
�i�ֱ��<�`�_�}Ձʘ�=�!Â`�na�Fg��U�S)�}��Bo��Ebs}�/�U�-: X�������ƹIj�"�f��Lt�q����9E�,��p'����[CṶ1<n�p�)�
�̹��*�^o�ƩLn����7�x�_ZC��;�7��·����G�O��}?2�\�/j��'co�C� ]v/��Ca���:�>ZYq`�����i��Z2K���r��t��YY���z�!L�2�UΑ~Y�\EX�g�Y�S��+<;�����y�Wl�s2L^�����ߧ����^]uC�޴��pS�E�7n�5j���kvR+e1B�V�O�̿T�}=Oĩ�&�1L�{�Z�^QhB��+�e�Z|+i'�xHJ{- eq�޼
�}=˱��d�ke@Q��#��OR��+���x��,k�3�yv;h'/����r���0q��ؠ�׶=5��-�����v�cO���lg��G�]��ζK�w;ۜ�{W�S:�4�ͻ���k��>���e9�=�������Z�����a�����^ݿ8�#��+�K�mhե^;&�a�Ϟ�IZ��N^5<��^l���e�ə�y�g1z��j��)G���h�~��GN3ƧY�$q��6�=��j�^v̔�.���[JIݛ1Ӯ�W���P�#��2�!ai���GRv)P�U�i�GO&�Tv�>�^�Q8���qB���ݵ���A�B�f�����,ҳPIN�X�'��y����é�{g;*�\WjN���U�X@[�s�C���+OJ4+�*z����B���qCVo���uZ.�[��r��aaw��Y��KѼ�ͽ�e 9CSA}������9�˞��	���@����}���c�M�kh�->���4Q����w)z������^�_��;e�nS�S/Ob,�(�)r=N{�S��:�f��zOwlŧ�2��B_\ǫ��kOV�GB��<�/OT#4�Bq��U�=2meZ�rrC����H��J���Ŕ"���t�h�r�w���+9zz�!f���R%��u��{MU�:�O�ѝ��|�Pn���"ҿ��.�]����n_%�y�u��^\.����v7����+y�w�z(v�-�"ıB;���f�+�\e��p��'�J�Y��9x�t�l���u�_er.ma�2��t8)�8%v�Q��hK�]�b�巂�D+2z���B�fk�u�~Sz����/;�Q����,�;aY���8���g�r��K�D��� �H�.��;C�RK��uݐ���ƥ�\�9��:�G�鿶c�Hh�x��LY����b��C7�+G�`�S7��������֑c\=�p���0͌I�!�O��y#kד4�*��x�-�RÙۈ;�Zúְ��]�2��XL�p{�l�
�V�/0zh�����H-�y���2$n!n��X�+�v��Z5���ط��ιl�#�;G#��#��d-��o��w�M{U�60s`�B�,=vNr�'G�ɏ��X�l?Kh���k����/צDk��.����3�?{�u�_\��{7
����b�]3��`թ_PcS(֨��{�K)ĽMU��.�7+�/]���w���pTy���=C=�ճ��]���3W
[h�M���R������X�{W��k+��t5KK3��s�>u,x�޷��{��Y���R�lJ�6��WW�//6.��bw�顶q����?:����h{`�����e�e3K�c���]��wY=ѷ�Q��u���f]Q}v�X��SW��J+�O>ɋ���f��"X�U]]��vb�썾����F���4bG���"�	�x�����B��,��R����9�٩y�dJ��f�w��� �X�D�	v����|��x
f^SJ[��4��o˵q���Ն[w�/�_G���������fq���`6t�B�j%t���B��U��P��.�]��I������t�6xJ���T���C|�J��&Y,�$��].*�'^���3GZF+�N��YM�ǥ^���A{uz�P��e'F�ju޹���γ$��}`vj3�.��N�6��Bqۚw:�hȱF/mڔC���岓������f�4�ٌٺR;N�-���C�LQ�<�q�}��#ǁ-�-�������Ub�K�x<�	��w%dA�+����Vxa��2�ÏƑ��9y�~Ĥޔ�u��Fb�R���-CY~�/]���%bJ�+�1���-p�-(��d�ѕR�z�?s|�k�(�%���\�J���*�����w$9�-%zమKW)��Q�]�����Rhr݃	��3��mAG`߬V�U.WɎZ�<6��E��c�;{�[nSh�ݑH����}���ӎ󰾯v83kŭOU�0Mg���Q¥�%2���Λ�ꌦ,Te��{Ue���U�C�j��.�k�) ꧱�?C;-�m��_������;ϣ�5��o0i��w��o(0^�3)�|����c����4���qn��Q�eY:�3��JN�^���6���h@o�I��8�S���t���'~�ʼ�z��h̄�R`���M�� ����YȖ�Z:|��T���d�����W�&�]���/6���t��[}���4=���ʠyPKRֲ�����Ϯ]��H�(LRm#<t�A����m�EEyJ�,��r[z��gq�/xO`�EG/>ƛk6�4!=��n?#�VFJ��`)jb�Y��Ư±�O�z�_�NQ��D�,u���o��+U�V	�A��$v]��^TI��`T�0TW�+X�=��ݯ��]E%<"�cqᕷm�F�	}�؍�����|CX��д�/��`�}����-r�UyElņ��z{�H�t��OntXfs�8�.Ս��y� G�#A��52�k�X����R�V�si	~[7�/���?fԺ�zrP_���e�>z0<�@/�� E�T�j���]����z!C�����r�QԱ���y�?}ՎT��r��B����~��r���m��`��jV*���gr�o����ie�*��+���moҶ�6�߳�w*�wn�w��v
�c��T:E�`�\EXL��g�L�ya�t�&{z{�(J��/�,�b��\Uo��*�N������Z �=���y7\.��i��u{��<\y3��[4:��O<�,y���r��w��m�l�H]K*J�/�b��Mf�U߯s5Ӌ:��l*�'=	u�{]{�u�z����"%��Gh��j�����mq���<�;g���=��N"^���{�5֫^B=K^��<=W�c�[K�)��ƞ7�-0�i1GU�i}P�����2�Y��%�hX�C�=���H2�M�墕�|��=l%��Z�	��"n�3�\`Z�{0q�E�Ȁ�#�z9:亮��_7�=:[�����~�<����ѓM��|���͈I�Q==���'�f�<J�W�D�a.�/ײz��=�"��E�S����i^Gp�*�}��}�Z�䃳��;��N���ߐCr`^3�J�D�݆�E�q����O�����rj�M��z��ޝך��|Yq=7��=+n�Fl���F���砸���y��;�x�-j��r�#+�|����'���'�,��L�t�|�*����Ug�~��fzrn�Ó�J��gN�^KYL��ϱs�4À';[�AZ�|#��r�uq��\C裊�ne����W�I��D=[7i��x!����;�����L��W�����/��b�1�կq����BqN}Ȅ/�Z㤂4���u�z�굧�~=	�w��z�u,u�W��5�L	����{"�τ�@�t�V*�� Y��C�Ѯ���v�vj�{�`���ѥe�ּɷq�Gy��Y�[��
� ps�ZW�:��]������.C�J��{��׻6��n�~N�j��\e�\�D����-$5��&�˪�g�5|#�����W���&׫�h��:�ڷ(��ͮk5<cg[��;�|�������\J��z��u��G�%�%�ޣ��j�uʒ9QNXf�A�*ۀ��n������ø����w ѫ�
v�Z�1F�+�:Y�Xֻ���4��:֎vi��E����,�T��h��V^}[D��
|�t.w��:[��v#<R�p�LEoT]��L���x�����3O��蚒`J��EG>����,�;j�o���=n��7�/m�F��sVnT6=�<�[�u؇t��ࠠ�Ȱ��#�t�Mbߵ��Ŕ����f����ofY�g�0i��I���3Y�_{��k�V�4�ǀGtöI]� y=#�I� �A޲�Y��x+���ƹX���:�0�";x=�-����p.�B�NG��S����wZ�'X�y��A}Q�{��LYn�8�52��Q1�R�	��@��Snt������_�秲��>���z�z;��~��w*�7��Ď�N�*�ߴ����Z��?2����t���bu53>u,x�zޮ���Yh�k�q�}Oe:Տ�԰z��-�D�.��R��gVTڡ8y'�E�����9|�����,�8N*����ge�˹��G<`R�D=���0]Qu�e`hz)�rQ9��1x��g�5pb�U
�����7�7� �Ʊ`�ː6vݫ�����+�,�9Yװ�y��Z �Ws�/�{���7j��R��4���%m0�1r�_j�W)�0F�ig,T�Ov��ӭ�Ov�-��y�a"J�z�[����q��ڼ��3�zOTl��n:奄0����Z�t���.,����uA���z��qg��]�,�ǒ�zl���~䲧x���/��Z]2'�BӤe2�L�M)�di��{������f�D7�y��w��Kf�sXt�wzr�u��|�F��X)s\�g����v�m4�8�Ӟm���0��ܱ�ҳ4�*Z��C|�\�w�%�6I�O�K�Ż���Yo9�1lM{S�j�z���{M8������VD��|��<3�;L�0�N^�X��~��a�����!�X���ù�ς��/�]��;���*�L�9E�(�mfp]A��>�W�gu�k5P!��~~��%�ã�[�d��, �z��K�����u��eO&�y.�7�И}���4��r���g�n'�mUMz`y:]��]�EH�ſ>f�j�U�;v+�83k�FD�.�*��Os78�5]9<bw�6.9��L�xX���g����+�i�<��i\n�o�����Ѽ۹z�ʗ��\�Hi�Ae'�(2ؘ�]w2H�\!D��]�N��Fr$a\a��PO�������U�aK��h4&A�m ��u;9m�tu����>����&Vr����jE��t���}���I}[��B57+�?I?��Y���<_�e���u�$�Gy����c��5\��5�2�ٙN�
���0W�}t�x���v;��/R��ؽ��^��|� pph���n��Ԛ���.�d'�?&"f}|5F�Ԭ�3�ص�wF��w�6��ǃD�U��Iq�rɠ/�BM�ޤ[+Ҋ�S���V�\?I����Ϳb��~4/L�t�\M7D�9�|�1ґZ9y!���H��Byzz�E��f��{��G����x���瘩�OĖ���lS)WI�d���y�˪����K.�陧�:���/�^L�j��s�kfR<�#�dh5�\�#%Y���X�v�@��:��9�\��Ҷ��"M��3��s�.S7.���D����t	�X��2a~�ċ��]zԴ-�q���g�Fʬ��>�e}�)�x{C;�����0�s	�&n�E����Ad���09DkY�����m�;&�ZYqg��`p�O���Sת��|�gLA%��&
��RJ�JE�eJ�5��;\�<�6 i+��SW�Q+>�K�m^}n��c��M�W���W�b!9�R��P�U\2��K֒m������̮Ǥ�����u�id�.���b�*-0�!����,�ӕϘV��}G�5C�\�C��R�i���u��(j�wVfOe�:�-�u�Kh�2g �nwV�fCŌ��7YpCrjj�굍w|�^=��:ވ�xf48�������������vU�N�*e���I�嵌����u�Ou�WJ`�7��|ؔ:W{N�U��6�L���_�K�SK8>vW_����=�j8��v+�4�������&��hG��U`2�$˛�� �����w������	Iג���uK���,����暜��êT웋xS�j�Y������V�ٮ�*���O����g�o�R	=W�;h'�t�3�! ��ͩb�"bE�<��Q����f��I\��Oy��.�`�F��yj������V��}}���y簑ם��O�b��B��G�˅�̃pRx2����]Ci���~�2J:�U���bƀRż	V4�S�D�x,4�w����'q���2�P�&�.mӬG�+���~�z����6�\��Ɲ��Z�Ռ�@�o�*\+^��LK���Iw��6 t!�յ�.|�O^�/���zi�Nή�{o+C�i��ė�Z�Է�v����Ⱥ3{�kYn�숎�Or�m`���xE��IY*�Z����$���ЍvV.�w.��N$^(��a3sY������Я)[�l:���Ew�)W���n�/J��n��-̮\��.s�� w�r*�n�iڸ7��(�}������[O�.��E�)e��v�q�0]G���kw2R�:��b�Wt�2�X��t��%���׉R���&Wp�y��7I�(S~fǯ)���C�l
C�N�WV4�\�6x��)V:�N������!�g��#�l�T�j�CA�6�9�S��V�\�<�l����{�j�<��(N��Ek[���(�K�S�k�Ոr�ua���g&岵��¬��k16(#a��v󻰔�')ii�q	�w�Rr㋭�4�%f �^��˖6���g+Ԭ��z�ī������[�$sn���]^O�F5ݘK��!�CA�\�ٔ	\7�P��^�n�"�!�тݾ�НO�~�n����!TĢ����8�Qe
r��K1\�&�lK�=�C���U�`���0ᬡ��{[�n\˔�{/�envX��soo�aL�	󍾷5�ɛ%��is06]��og���n,�W5ݽ�.@�6���i0�h8]�q�S��/vc��c!^��
�	�#Q��+�vR�����u|�81kK�֖;;�j@ܥ�1<o�0.��r(A�	�|;����r��oiF�Q���($
x�3�q��yvU�]�/)D�2/7(J|/�,��@p�jV�F���aq[F����mm�5��%h6�ض[KmRŕL2�(��fU�QTT��QjZ��R�kF%E�imc�X��������h����������VV��m+jDj�ȶ�*���Dm���eS0��F�-+�mjڴ�[j����-h��+�IV�*R�K[*�R�`,�h�n�[KYAm�b	P�ШR���k�Q*,Z�JQ�iX6![lV��մ���A��(��,0*Z4���-Z%��-�[-V��Um�P��+mF�m��e�m�()Z����h��b�Kk%������F�R2�[DR�)j�iQ�-h�ll��R�QZ�m�KQ���֬ŸeF5�*V-,�U���҃m)K��-m���[.��w�fi�,}��>ڮ��g!��0r#�/gwX�-��Ӯ�s[` ]dòԈƶ���4�e��U�N����S���F����P�	��F���t�m�x=��-yh���
��.5%�<�$^G,tC�s�n}ޚ,X�0�Y��
d��9�U��w�yecC~�좠�k3��ߣ���\+{�/T��SΡҵ���񘞠}�.�,�Z�+[][���p��{p�8Ĥ����f;\�xSI�^�U�!U�2&`8g�r�X����4��DD�	|��Yq.��l�;=u�z�ڳ>�gR����ِ�� ��}NfR]�����=�!��N㨹'wMj�x�m�*ª�e�D�zK��0+�Ԉ��0�����o=�y�v���jN��影��j�0���OK���#.-g�s�]E�}�.� �;~�MV��$-����'Gx�S�˭��CS���h{�ƽ�;Lά��(3�GRv)P��M�Y䠪Vک����t���N�L���FX���Nv6�t�G�E��E�\k���sx�-����d����i�"�n�v|:�4��L���Os�g&V��@���؋>�j����`�Wt�4$���{2޷O}EVc8��"������]��پk����X��hz��{l���4ҍ��f%��m��"��w[�,C�m.9̿8����g>��vL>�[w�^���\�]��׎J����u�u���m��麰��-�ɐ-����1��*1R��Q
�g]���w��i8����Cԍ㹀U��`���k>���ﺇM��9��׉t
)L��S/e�6���P?Wbp[��XA��@����Ө]��=�	t�,�BJ�,��dg}�ot���Pm��٪gL2��.T"��$�f�+�\e�A��v7����}��1���(jU�+�fJ�Ȫ�'��;	TD6��
�,霻Ha\���:���^����C/בlZE�s���䊎Ee�a�OR�����,��;3]�B���o���,
�U,��k���=ii����0wK�pXW����>\̆\�ed��]�`;}^�楩{K��Q^�\\�I���P��ܰS}��^�t́V��b5�O{�'��x2ka��c�k���m?�r��q�b1�/;����3�ͧs=��)�ز��e��u�PϽ��g�ydν:u*�]�dyPq�?3^m�OwwGם� ֌���&l�աO���Q��e>B�p���o[��"��T,l ��>O�哟���˼�\:�s ύ-���c�,�����~!>�����^�c%kPպt
)7[�q��[�K^��Fr�>�+���<}n��>��`3TiV�3�9�}��=C/��ڲ�k�'ɲ {�?H�5�:����;�x��m��<�J��lҡi֖eӹ�|�X��7���OvK����'xsB�������۴�ҕE�LP��D��(��h��Ψs���C�`����s�]�޸g�yz^8��|YVWR�l�Ȳ��̺�;��)��O):�V'�e���%�O
��}�'_���1a�c^�-N��`�.,2�;��;���|���מzd��a�:�<�P^K��T�>P�*-�^�胵l�D�H���l.�Z	��M)���3���`�?l/��c�\�{��\�3%ޜ�[ŀ�!ӠAY����*���<�W�{-I���>�:䙰�-rܱ��J���j�.>�E�9�ˇp	�K6l���/C�hrObo�C�X���Q��q�G����6��?Ev�{�Y�C�կB�=����V%�̷��(��C!�ϩC��-3@e��}��Y�wL	+��
��1�]Z���U��Pc��}�7E��c�t>[��A����3����<l�ky*�6�j���!ψUi�Ai�Д÷�����uk[���
^�u���H��{-͵2��w�jڙ}Fnƥq�ǉ��F7���{�<�.rӷ��w*�׭�]�����i�Z:]�2�,S�Q#�b���m�gO�CúZJ�O��;O��^��͞�0(6X`�:Ƶ/NGK�߄��>���4�*�>LpU%�Y��{.?y`��J����2��||,u��	V<�E�����ygݝbnR��׵fT��s�e��Uk��[�o��P����ٽx
��8'������=��vj����IL��o��}�Q�Sݥ&R��.���Y����0S������g��F�e����K�g�zWbfz���{�h�0?��m'�L�W�P��y&�����p�Z��%��x�B��0���s�Ǎ�/c�~�Á��,�8Ih����P�ؑl�ҋ�A���q��ts�_GYԇ��sW��Cܰ1�i��-'8ũ��"�t~lt�����sz��N���Y�&��>��H���/��7�b�,<l<TGZZ%�L�qkۃ{�)�X#LN��	gr����zu�,OntX}��<�� �v�ힴ{�P,��}Aˠ}7݋�������7xl+��c&�7F��O#B�����S_��{u�,`�����9t=`;z�n2)WwI�μt�{ҷ���u������\��i�'��-J=�j�6%�h�\*u�H*�ĭ��X^���:���u{m�k��w���+�P�%��֙�n�Jۇ^ʱ�X�������{%��&Y0�Vt�<sO��Y�����:NrD�����ߌ�����������E��`�w��COu�kY�7�uś�i����w�)hu�"�<I<+Q�\1T�u�-�9�K.,�`z�7.��N�:����m�w�:Q��>�br�0T2�KJE��Qэ@k�D����.�{�@ڳ�o��s�x���P�j탎Q#A�/��+}�T��V#�8�뿦V��a���7��)�gs�ڱ�Ãa�n��q�%hLƉp&Iߣ�}c�bgzאr�#T~ݕ�Aռ�=<�(kW�L����5Z��j�
3�<G���kݢ���^�'GZ�}�-��{���]�(��
�2k�V��uc�ȹ�����zz���j�P<���҆������V\���3ĸa.��m�� >����3��}Nf�����U���b2s������>Oe��`�
��k�V=�r�]N`l�#��	0�v�^���(�Wd�:\�N��P�V.�w�w�<��s���\}��	º���l@`���Ԕ�\E� �����E��W�ɨt�]�C���Zl��a]��#p�����r�MFLw�zn��-l��32-Y�X-<M���4䛫K�����-wU��˚����xOK�Uم�+.-gҗ=�]B��^ �wh��r����jF�ԉM�G|���RmN5�Y�x��+-rJ�ԟ�l�Md)�k׵�7oӚ���4�zT3�;���0�:�-�^�ؐ�W�#��y^�Fa[L��72����0$��H�z����x�þL���s��Y�2��^
e�]�Ӟ�r�����l~�Y�Y�jJ\�<a �,�C��<���a�r
���D{���s�͚�/)��]cmm��R@Ϲ҉_�LƲ�dPƃ��:m4��Y�^���b���9u����x��?o��g�`���:E�t�yw_��`�&	epx��,�93�:���Wl���Z�r�B%'��I
�rV)�b��}���;&[����:�Bh�V�c���T�.ڋ�;r��]���>�{�M�U{=�~���ďb�p�/׍xl�#3��/;�Q��=J:G����A�˴U^�B�ku���M&�N�g���t��1�WV��Q��N�&�03k����Loo9�^4��:�O.����R��,�ɣ.�L�S8ܻq�Z�]�J��a� ������q��V1�{����s{m�s�SW��e.c�����,(wR&>v_F5�wAb��PY�eś���aδ���N�Q��L���.L�Ei�]Uk+�ۼ��}���c�LS��!�J+��ˋ���C/�֠.:�7+��S����yţ��ok[k��N������� ��`uY1�O�-b5��i]R�c�돃�0�!1��c}��Im���_��-��z�_�����;����c�OV�����3�}��n�:��aACW�H;��#���)�j�{WD���f
s0��;P�Gq�LP���G�f�/9]C�}U��_;��{�����C�C���y1ZY�N�(|�<ro[��OvC��g���q����^��F���CL�[Jm*E���Z�OR�.ql:����k�d������ݽуv>���Ն�<�"U�`��:��v�<����+��8���Q�O+p��E����:���5y�>׆�:��~N��eqq`������݇� ��T+i�|�1�������D8�y��8�Y��v��H�.�5ɥ��L���3<���m%�ɡ,i7L�V�s'G.m���4�m�^�p5��-[��9Kᘀ�NPǒq������ػ��9�7vVX��5<C$Z�X2²b=&�'b��oc�t�橪�X���s@a��r�E��W2��Td�%�Č�����m���vw����'3��Ӄ����~w1�.k��N\��(��@�5��D�8.��r�f���Z���ʉCo��!��c_�fi��b�5��p�L�Y��l�[WAfn�����$��K�X��wT,�L��Q՝��<��?��'(e��b} �����6����^�q��VXD*�¶T��y���:��	�ƀ������k��ެO'g�u��Z-h�Z:lL���yL�u0�g�{ �p��������x_V4��TNV��swy��Ik�AA���r�&�܎���	֍�ia���r�E6���cdܳ��r�^wl�!��{x��ˏ��s	V��H��[ҽl�f׋Z����:�,���ξ�ǹ9M��U��`ڷoDਹ��Kf��	�g�>�����åi���Ik�L�������{��= ��Y��j��!�n�9�lPe�3�w1x�����J�v) j�D�-o{��o�6��3>��O ��R��
�a���$�\��r���,/{�t�p���ċW�|��3�0�k(Z�2Z���g�@�ć��Ls3҂w�ko�E�u��I�yٳ/uofgr��ˤ�j�q^Óx]bT�QWd���6�v�Q�!�T瑯n�}^�x�xhsOO!�k�S#�"�6��9[K�ܒYR6�7s�&a��=��*���J�ʭ/���Z=�h�u���J56�^HG��u��]oۮx�jj�arޯN*�L���T4�p���:"�t���{g����F���ҩ�u>��H��=�e��;���Cya�1S��6Dq�I���[�}��Z��H�������浳����u˚�%m�=�֌�<��ה⬯���k��s�]ZP@���c����߈�0%<�(P�y}i�v�j�Ҷ�עU�"Ĝ��>��{%����\�.��}l�4�3O��&x���}4VWxb��06��Q}٥��b����]�vH�n�r��|x��5Ɨ��@�[�x��
�X��x:��C������m;��/}�g��\\�,�)���Ӎѵ��',�`�e��D��¥quL����(F���ުJ��3�a�����Ǟ�J/>�탁�$h6$��o.�������O%��c �l��y�����u��o������h�r�Z���L���>�U��*J�I�w�v]�GK���PL*��l_BJĬ����/���O��c�|8N�h�՛�s}�s��c��;��)� ��>��]!������ŝ�0��*�3�K'���^�n{g-�r_G"b��思��Sc�=��������-�2��>���dJ�;�2��Q�7$������#ʻ=l�����#��OR�����!2m���Y���m;�(9�j��93�_������LV�ȸ5�9m$a��x�`�#��wv���x�Kx����=u�%��ES:�����֮̀"[c��3�.~�O�T�y�<��dk��s��7NW^=Q��/��k�%cز�iW�;&�H��۝�,\�;�Z�S��kÄ�*V�ʒ�?��^0�����W�<JjڍPq���PT͙��w\���p���x/MF���iĲT"����M���q�r��1U.C�W^����^&�b�ԓZ�i�T�B�k�]�x�i��MC7�v#.zƘK�n��|'���jyF�|�Ue�(Ƿb�mR>%��'�9�H�j�˱���,��]{a�׽)��m-l��If����}��ΏQ�7؏�h�R�l�0�qvR���y�kOV�{�ʪ��Bư�{�nz^h{�p�m��k�gX:/Z4��tv�J��O�z���z��$��	!I����$��	!I@�$��	!I� IO��	!I�@�$���$ I?�H@����$�$�	'�IJ��$�H@�xB����$����$�$�	'��$ I?�	!I�B���(+$�k4��� Ri�0
 ��d��H�_=�JW�AUUH�R�)*(EUJ�$AER�(���JB@֥(D��"�R�EB��"JR�B�P��J$*���HQ@�
T
I(�QT!@[5�T�
ք��D�HJET����$��d��U
R]��Q(Q"U`����RR�QI%"J@���R��u�JA((lhT�TAT� ��$*J�*��JR��R�T�Q*���PUT��< ��4 ̰h�� �a��m�MwuN�mSq0��
r����mkJh�L�:h)�i��u�h3E���]	UQ$P�
�)#x ��^F�v�Z�Sm�ݝ��rMtҺWK��u�j�w)[���n��.���vt*�A�v��c�m�k��E��Tt�!v�P�R�ED��AUU   �G ht4(c����B�
=��(P�B� ���(P�BE
(w�P���B�����`�t(P�CCB�;�
(P���U�)�� ��P;m��K��@ku)T!%*JJ�k(Gm'�  �i�@l�㫘��t�S�5�T��
��ӥ;�]�N��87V�)��:�ì4+�V톫�ݚ�sf˭���wK��T�w*��UIHQR� E�
�  �ޚѣ'M7[NA��N�uM@ڝ�w7wn馊�7�iX���P�n�\���Jj۝�]���n�v��*""�%�B���(�  gm�uٔ�Ҷ��avhU���B�m\�GM��8۪U�ks�(.�9U���
i��(�QwEnt��M.�Z�;��;ri!R�"*���J�  m;�([4��	�p�5��0�2kCX�7n�R��7lv�CMq��`�����M���
u�����ꂀ�;Q����m�BH��IT��JUG� &�
([�� u` ��� U�(3e���� �,V J+0 n� nT�$%R�$�<  {�� �� ���Z,4 ���զ�� ��
ݳ�TQC�� �A* J�UQ���� ;������EfL��V� �@��1@�A@&�h4�X  � ���eIR������$�J4��)����  S�A)R@F���UJ � R"cU)#L� �%[� #A" ��FNI�V���ce"U0a&=���Up��t��{��{��v?��
� (�� TA_������D�D�y�?�?���3P��n7.��D9��TL���r�1�$��R`�JMX��Rp?�ɷ��bͱDIR�B�.����Y&K �o
H�L�v~״"��	u)�f|��س(g0e�����T0ޭ��2��m��KA���EV^݅t��@�0B`Ҩ�҂Ri+�Z��J[{V5��,�I��J?Z�'f=��KM"K���ޔ"�J�,h�d�.�B@#�л7y[)�1�
ۈcz�q�,����v���l�]�[kĭ$������@�ԠEm9�M[�0��B`)����w�k�"��1����	+:�AZ/hTC+]n�M�Ҍ�{4D�p�vE��+VU�/t`��בju"��/(S"5��E֡WW�̀�u��P͊j�ѴKߍ�e���A�q�<�Go%aPX�*�Ђ,�'N�ۡ��i+	�h���w%Kv�aVVu�#�_$�fb;C�-���*PU�h���ͬ4��rӄawZ��k0�jZɦ���������jmXM�FL�o1��x2�e���j�2[���f�]\(���xj����GB�= E�Ճ%Vj���)em�%F`կ2�[6U�6�R��%��N��+Z���֯f�c�m�3+)c�詎e�o]ō�b���W��e<�N$�{n]9�;6�-�i�ڍ=�w5�v��k�u��eM�h�%֯�[)7�j��X�fҺ� �1�Z��ݫɸ�k��Ȼ��\A�ɖ0]-����e���bh���l\Z�F�JQ�r�R*�c,�R�{eBJ�J��(�4���&�KK�VP�����-���^�V�!nH�����6�0��!�WWx��74CEd�y�ޣ�:6�����$�i`)�˶�[P��g�/�Ӹq��.d�>8��/4�`^*f�Go2��},�<��{���Hl���dȳkf�Y���ڕ��S�Qf���x'%���X�"���u�X�D�H!�mde���Lђ���y{#��4���.�*i�ZX�@惖ݽ�)F��W%�+n}
�[e��b��3HH��ɯ*`�ASVIYvr�w]$�����+5���w��T%-�v�U^�)LA�p��e�� L��[�#��F�ۺٯH`�.��r�����NM$�x VM���n�f�q^;"�wKR,�l��Y��K�ȩ=i[I��!��[i�d���z^m^���d�y �1����J�f�:UHMH�쇖l��,�7TˀӴ̎�&�^�I�yy��V�CyG,|�(
"o*	�Ja�f���wtۊ�wv��)�uJO�̂9��;%ZCj2��yv�wS*�c�\e��j1z��R�ۖE�ǀ�m4��K��N|ki-̰�=T�odudٹ1�y���r��Mke�%1��K�1���Z$�m�*�1���'R�$4�72�U��%hͩIӣfEՁL� e�W6�0�V�E��,CB�,a�J�#�j���ӄ+[H��j��Ձ�KMc53(�jn��DI����*`˹�@(��!v�Mw�Œ�ѓD�Xs���_l)InT�&��iǯ#T^$�^�$(0�sȳ5	&ܬ��Un�w�
�M�$� �x�)��2�;�̻��6\+R��`ѕ{V.�V2�.]Au��il�T5o�[V���R�"wIdGQ�1�W�A"2�ׂ
1�ʁU�c0�e/�nԶ��B�R(Tx�3I@LN���4x��U�J�rг[���++tK��Z#7M�qeQͬ�u�-�*�2;�gj!>��[h��`�Z�V&���+6�4=ի��*/a�b��-8[m�iեg�̏별�=tc���d�ǥd�2����#V謍�Y�����E�SU�R�[�6�i��F��T։vN�vs45/�w䅚��Y7=d�9&�du�f,ʺ��iQF���Y�'B��5X2YoA��WZ��V�ӌ`Q^F��n��+����I�5��G2�*[Z�c[xB�ml7%kJ��]�у�[קU��=�+�YM�� 3eE�;�7\@�,"��v(
���-G���0iqw����q:�!��y*��]��]���Ҩ�jt��Q�eE��#*����X4;��6<^�Q�X�V[4�]�@�����*ae-�*՜v��w,�\��w�A�r��Ҧf��Ы.f	F^��r�1&�{FLIZ���f�WYU��i�:.�U��Rmd����v�A�wz+&j�,�K)/Vǰ��Y�Hi72��-Ӥ����˺�2ն@�4\Q��5�r�-�7U�Zo�W"gYP]e�҆�fnͺa1��އ���4K�g#V6��2lW�ZU����,�i�.����MP�ZFj
�ʕ��6BE�[�����i�͡{�p=��V-��\L�[ �;Gk.����t^3�=,��qS6�%B�V� �v����&�ЫĄH����X���\$�
�0�d��Q�V3���D�6�AI����߃��:P�*@[HVX�0��@f(*)�xRC���̻�ZL�_e=��$��\�we�u����O.�R�1���FTur*7�����$���´��,�%@&��ӂ�죻E�R�4����'{�[�͍0+'�ȶ*��϶/76&����tmY���c;���=���pE�5a�K;�PϦV�1����l[����՛X�p�P:4�S�df�k*I� �U�w%�nAW�h�-5��A��X�<��v��nք�]�"A��V��v؎Qt�9oA�jYd���d��6Љ���!h�nAr^�kF�a�Z�:Ʋ�U��ڏp�̫�7g�%ԛ��ӵ����e�(`�^���U�A��z
lP���� ���p��]�:�{-��սlJ��)��r%�i����(VLJe�ښ�QPՖbS�&���`"��{Gjݽ�+*Dl&%��,^�Nm��R�5��
ȫd�!�a�2�P"I^�yXK�k
*܎���)ګ�H!s�ߎ�6�Ϭ�"f�N�@�Jۣ���@!��fۑ�I�������f$Mޱ@��̬;��D�i����F�5b�6o��$��JYhm#@�r��as�Cv����ɳ'ڦ"�PQ�a�3>v
��Ŭd�x�d8�mޛ����$�zd4�*��1��ԠT����^e�֪�Ɗ��y�PaW�C�[,:Yq�o�i��l<w ��n�,i�0�F<wl*4�B.�R�]�e��|��cu�����;�`�j��=�g	{�=�����!� ;�i�̼�w�h�F����Qj=�fU�D�l_n7;�fA�Vh�j���,�u�B�a��96os,*=څ��(AGN��U��X�N��4�(����
M��ͣx���+q*4F� �u�N�In�@� -�O �-i_ف�6��X��K��q�[[C"���,]�Ee��5�M@�d؀ѕ��Dm�)�2�V���:��*0�ܰ޲�@�wk�M=N��-��e�]��Z�Zϳ��z��d�J�,-�$�)*KA ��x���t`�Rv+n�}�ցr�����"u+
𛺥�[��Բ��t��f͌��KR�G�if������;��K*��hz��Q�4GK[оXPN��ӹovط���Y�[
&н�}��Շ�\��b^K���'i���a���@�ܤ��vL/b�X�lbV�EEm����K��Q��ҚJ�A�vB�1{�4��.��.��6R/n;D��)8e����kT����9t1���s2 �9���Y�tQ��d+����,���ț4j��f��GM���R�u7/2�,@��z3>��f	XD`O����Q�f�F#f�6
�ç_	����ojU�1^�\$nh`���3��a�*��eӈF�6���R٤R�Mbl8Te=�V���ۢ�Q=e�/�b�h-�^D�������Ck ��G(c&��RÃ$��ɕe�зM]l�r��̵��NL��V�1`�FV&��Yn��"Y��6/A@��3I0LB�b�Av5N㵵q���5a����ke�U7x7pd&�e�e�(���
n��JSFޫ����������F���e-�c���d6Ѱ7i��^�h��՗M\fb�&�14w7Mdm�U@��$,`�6�B��;F�iɦ��Q�RP+Jٸ�bո�в�L�l����+QǏ~��8�BB(��Ӏ�����&��pk�ė{s .殺�� ��M��M�W�F�˫����YR����5�����ˎ�S`�Tu���&�QlT#-�)/C��,��al��e����fdcj��ЍS��v�>�(��Ѹ:6�}���pL��yQKׇ!o����\H�)Y����jV��W�5pLJ���z�Uf�����S5j*�R��U�$�b�րۂ�]#�J���P��X�D����?�H�k�v4LT���wW5��j�0���![=x-���a�`�y��o@ Zt�@�e���rR.�_� �4,���*�2���X@Z������@&ȎZ��Zn!+.���̃�oU�n�EXhA�T]��H���L[F�!��[̥*�lE ��kMh��F��Z�R���w[���v�u
Vtʼ-��E��A�{�sh����n	������j����	=�ؗ��t:�Y�����T]�Oc�;�!���l�.b��ossH��sT;֢@n|
�z�0(mªd�ҍ�1��͋�u�%��,�b��
� $��^�t�(#+c�ϧ�E2����<�r�'�u��]�F�M�ٌ���'ac����q�{�R1�$�#��?43bܫ�;#(����ީ�l���ll�ɋ1ҫ��n�qnݳ�5�Mݵ��[h���V���{)Y��2��jT��w���,ʸXw��Q��fa9B֦j"/0jN�q���{�О&ӻ�e^ne��s/��	���nA�*�i�C�R�,U����{"N���	�X����J&n8���bf9�U��M]:hYö��C&��fB�X_<�X����G>j�fM(b�CL
l�g"�͋�Q�:����ź�"���[FKJ����6f�@�5��L�U��:Ajȯ�[Q�(G��j��8�{[��
���W(��c/4�jƆ��m�h�e�PѴ�9A;��(�m���$��8̧�@`�,��6A%N��ɸ�(�9�a-��P�w"��j�,s�����)����;ǋ��QS�|�L:�4+L�1��E$���B��uB���q#}˹z�.ޝLne)l�Β�$�=:)_�K��q�Y�{��v�kh�ʶ�WX�It��J�fT�dڵf�
 J� X�9N�m:e���ܛW��FVk�a6��):�)�]�Y۶33B"��k��S2B�U�Mӄ���{�ɩ�U��n�tk�&)��Y��7R�DrI��q�
��)٧/qt�V���"�cdƦ���#��,�zS�f��ba��wBV��oŢ@+(�7+U�D��٭`���	t:@hui�Z�
�Vd���v�[X�e3IZ��嫙�Mi��CF3t#�t��j",�T�ݹn�b�ЗVS�)��e�te�Y�LT�&A�k�
{���ܢN!9u�B��	1���١d��)�&Z��cf��0�/�DS�!À�J1�����ĭ�Y�E� �d�r�JD��CSn
$'ƕ�X�X֊�y�����9ˆov3t��v�H.3/)PZ��)#�Oӭ!W� �`4��b�q�En��J�荩�'3�4^) ���p����(kıυ<1��X���kCEh� ��R�W�V8E2>��85ژD˅�t�bb×�Ke�:E��(�Ǘw���*�UB@���*�m���<I�#v�VQ8@aj4\�u)m��q��oCi\i�-;��.���OI�N]��Sc������ ��%���&�qb������R-�*�v՜�)�pS�(����S*�� v�M8�m�BR��M, �`�!%ڧyyWh	vM6ԤͱXue2����wX^�9G,V�,P)m�x�)-	˅Z�;���k0����.��XX�5�G�cq�v����� �ɎK�Pa���-�5V2��Y�� [Œ˩��"7�����U�]�	�B�i��b�^K�)�ɩG]kM#b+ܒ�,CKB�T���4��2jy0mɆ�����U�%��i5uu�1�n�omѰ�y��hE^�� #�P�X�e�¼�&Ÿڇ#v�hf�F��]m˭2��K��*���JRŧZ�q����T�شlHASW�i�]�X�ڛ���m��W����!k�����X�Iot�q�T�)�w,��UꒊA"�PL�r%�Ż�������f�Ku������JV��/,ŦyY ���ꔀ$:��6�[�2a��[�q�I%M
�a�`Hs�+1e7�� V �$X�mT��w�V�) cH���	E��fn�@��qS�o�M^������Ɲ#d� $��R��f��P�-C�����t�"�SS���W�k1�-y �`R�u^8j�#����1
	nG�݂�hT����/4f�&D���U�3QV��+ T� ���H�n�6��lWhٛx��������i��U��``	��ԭK(gH�Zܵ�8Bv:ᩏ0P�N�Ӗ�S0�@�9I�5�*���˵q[��Ӄ*mg��;�s��ֽ�o��⩙�����WQbu�k�:>R�j};h.�f�zt�̺ky�;݌����]td��1ʶ�I�n��wkB��6�� nQT���G
d�D�L�Z,ur*t�Ez�9�s'4�ZI�-8��Zɨ{@�P7F.�,��6;hi���/�g7C�<Š%��.���k�D ���4�fL� a.0����!��[f�=���3��ԍ��������Zʲv۲r�tX���ZHS���^�N�Y��`�ԕ
�Ws8pz��YF;�1�.��j�Ng!F��<�Vͬ�c۬ˈf����[Sc��'�mĢI\��f�֚�Ţ�3{��*ou�Ɓ暂��!%C-u�"<E�*�Wq:�uR��݂������ݳ���H����P��^J����]�y� Iu*�h��R����ѧ���I�Q��u��U��>ͼ�mш�ا�+��_2����
����^.�)VB����pm����؛�+��Rո:��:�>�ܺ�r�B���a�4��N�vG�ť�P�:����s�q�J͎�᫽��M�����D���OF)�VR����y��#-����L�؍*1;k�PU��=ւ��y
r�iI�m}�����gH�M�%a���nᎄ���ni���$bu�/#����eoEr�Z)�J���;8Z�uG����$�c6,¯
ba��`����7�1wegX���Ν�|-����Ɏv  '��ǖ.�|�����Z�]ܽO�w�P��烩���{��0�]��-i��U��֚ͮu�n^�_�ʈr܄5��wfuiP3v��\��%�q�O^�ݝ�XU	�q�dS(���PU�����[O8_f��b�*���v�=u��9�V��W����>�ϣ�q�����j(R�u�m����[}X(��1�WĴ��eU����e]��<� +{���a7�Tt�b���9��v�|�wCJZ�!����\� ܠ]���w��m]�6��S-�@�팚���d���{؈@���eU�Yx�v�ؘ�3r�
�rܫ�!d*_*��"�N�,6�I�;��>�fީ��CRV�H��w 4z�k�*Bs	�SF��yC��q��|ҟ*Ѣ�곝.����=>��l9]��橕�u��C:�=}]��e���ˢ�j)�Ik&X��j4�xi]by�,�3��%+CxSe��2v.�����k�䨋�%sk-S���ׇ�;�N�U�&�XĖ8bޗ��z6���'lr$K�.�[�� ����Hj��W��	mwUӝsZ�@�)���1��°���8P�zYe`6%w[�9�.��ɔ��zP�;1F��k���}=�k1�tc)��/k:��1^�B	L�₸
��ѩ��J�:pu�V�|ӌ�Yb*	R;F�*�ڿ���B]7֓�@�NP7:��ɒ��vZ��:��Z�!�*�j����5���u�\�noxEm0#��9�5B�m�a�zBW~qwj��$�z��)fM��L��C�3�@-��-�}	u��yLO.�ϻei�x�j���VR�V&{�̎���]b��t�;d}:�~�噹*���Ցu,n�OP�ӧwDRL�r;����G��Z�yҗy@Y)�S2m��vb5��M�������[�׳���X�nƷ��C/�*�뭺)�;Fܝ�G-�ǥ�yB��N�����/���bK��v6�$�,��Ʈ�&2��o�Q��t=/rT놂�_G���\/�6���v�7{W��3� Z�Nջhg�)v�HRnu�x����Q��5{#�wcӘ�C]�x+ip���$�Zq�E-ֻ��X��5t�=��D {x�;���f`��M��w[�i��ڕ-,��d��s�mD���o@ā��@�R���h�Gz��un�����,�s�� 4��gn�,+X'*9��kUB5��e7R�dͅ,��#�7=��G@$��5Ⴊ"�����N�jl6�1k	��Ӻ�%eҦ,�Iue��j�u6X��3r��|$�;��ۧ=�O�h6PJ�8��ZٟuZk�Bdp���/\9�[���1�;�@Mhk��k�88wX1f���Q&�A��p�^7�v
�8_|;LL�R9b�1۽��|���@Q�#�%F�=u���(�#99t�M�E�*{�^�ܳו؎ �<��X7��c���KT��M��4h냴�������L�*U�]�n6�`���N��n�'t�z�os�VyWnPݧzqn�Z)�ӌ�قv��$r5dT���t��)���$��S;w��FnUl�K©N�O��N'���\J���Yr�k>�-���uv�9'�v����ެ���E��VG��ox��6ԭ��a|�N�S��T�R����n�ɒ��Y���dpz��:�+�-�:���^{�u�qz�0%,� ��a��go��N���&A�n>K�
2��1���-�ʲ�*3��4��<s�נ+#�̼�/VdV�*�n�Ivr�5��͗ϙf"������nX�]�u9�Wr��4��5�0�β`��c.����.k�Mκ�e����P���G��eI*!��wWQә������g3%�u�7bAYǣxV��W
��lW6!��;^$K5�%{�K�k��XjB�:�u:W��U�sS����;:J���I�.�5���^s�}��ް������u���e�΅as��C��+-I_��Q��M.����I@��j
'݆�b�$�w8E��u���q�n���]dnU���ˬX�"Auʥ��������t��Xz�.�'��c���.�����M��|�s �H	�V*;n�ʂ>6��|�L����أ��s�����%�L2�@���ӹ[�����M�%��D9���=w˦V�����u��-���2��$�x6���q��gT��Q(��u�W0�^v��;��n.�R��_0]Ӽ��(t�{�`�cn�b&.Vɚ��׊ʨ��Eӗ�f�j"6���U��1��/r���-I(Ǳ�*��'�V�9H����F��b��h���*z��Ii�jރ�6����Gȹ�)�Y9��;��.c�mL��][rQQг0L��4<���TjuG������D���1}[w�_B��+3�����һ�ݍD�O܎W%h� �޺��l"�;�9�@�E�T/dn3F�#3�T���U��	�1w�� Ƴ��&�X�=8jkV4�u��f2�+f��S4vD��Y�bj]m3�$e���ڝi�>(]�9*oO���ҭ���	S�Y-�|�e��|��[i�!�鐟�����x��l�Di郵QB��̕Md��s���X�5)��pQ��݈�t��k��i.�qu�m'q1�h��xx9�Tܫ��nk��F�N��ܬ)!)�� aɄM�y;�DM[����ZԔ%[i��u֚0������t�!1��z�7��E����Jŕ��]֯�\����ȓ�)ۤk5�WlG�y7�8�kKl6�U�����r���1w$6�&#�n����m��.�X��S�%�
cED��U�Ǡ.Kq���/��9Q��*P�t��Tg8�=;Vi-WP7d�:����n���_aZ5R�Lަ>�@D��H�'{�G+<3��^v������9ɺxq�ǆ����0v�S:Ӑ|�gW-���6�}0K�2�@��LF�Z�<��'JxD��$�^�c����^nF
k�����f������vBfx�:J�v�{�1˽�]��i�]�u-��5R�Z��uɌ}�������=���*��}���
�6�IMG�Z��דJ|ps��e\b�����d��r��R�<ZB�sJֵ��:X��Ou�%W9iOK�9�/v��e�y��𓫃بf4-�E�|4TE�\�|��Z�F^�s��u��ԝ�@$fM ��W�:�^�� �v�gCv�	2��xv��ڐ�xVv�P�]pVJ����ɲ�*���zҾ\(����?]��+jnuvtk����!�n�Π��=�y����uL�t�7-�z1�Ү�6�U���mZ_I
2�c�]�;�����c�H"���/8=�ln���9�F��\�u�ū/��oO�ec�{]�g
}�k}۴��mD&�f��N��p.�>s�����a:�&s�e�kiE���0�s�e�i�` ��|�R[�������}W6!�!�']]����&�R�h.!

j��?gN�Qg�l���训'3(��s��b�q�OF�͸_ o{���Wk��ӛw�9��1��R�.����+�-\N@h�sh�  ��F�^���]:�wy0�]��[�sQ��tB�+���x�Λ���ٶ#���03b@��2t��{����ar0�]!+(L׭R�z;-�az6�r�t��>ƒה�*c�������J1�𺒮c�D�Ѫ�\���B�޹��\����6���\��|�&{�4�������r��np��V�$r;\�Q]b\Mn�(Q�b�'�b���J- 3[�ܤ�n��6w�(���;F��`1ͬ�5���)�Lm��������@���//���%]��X��_,�bڤ.�y�}f����4�ʁU��!N�֞�F���2��s�ya�5h��y�]y��É�ÎU��E&��;�P���b���l�{��7fol���.�g��/��e+H¡��*�ʴ�!|�e�%v�[pր#�ebX#loV�j��Ѡ�Z�;+�|K�Z�ϯf�%>���p�b�;F<��Ó�1\�b\�VX�`�xz_\��n�2pdM��s����y
��q �ft1�/:rMW.�]5�8t;�8��^���-b릻��)�,:'���']�f����mM��u�i�)U����`���*�;��zf]0gv���V[�ћǊ���"��[��ȸ;C�ft���lκHg�Z^}��	- ��-v�#U�������{��WQ�3�� Cp��;x�)Wū^R�Ep�Y�,ܜ�v�O�b�6��۷��T3�Y3��\K�Z�D�]�G�`�%��(깧��ڎ��L(�.��4��c]��/]AP� m�T�'�H��mӚ�X�1��K�{����Q�G�k�C8����<�(��,T��rv�EwSA�r�IVi͊a�5�B��:�,귋"�A�t��������r|��Vi��$�/�P]��'i9a� ھ#�]�-�,����W^�!��X�� ^���d�n�ܝ�ڝ����u����\�����r����S��>��wT3����h-�Y�����pΦm�j��5<x�PVg8��d�\�`��7��b���}�*���z�#�VNml۠�R˼wQ¸�Aܾ��gN��w[7�;�h�i��!$��ے�4U�ɽ���\o%�1-��Ҳ��to�B(#v���
�7��-�yQ�O�s�Z;F�m:�wv��'��hs	S��� ��E�b��Uҝ��k�J9�_��Y�y��!\8ѣ��E`�\�h7���ܚ�P�cbJw!]��	��oB��t�Ig��6�b�}��]0����]����m�%�1�nv���J�d�Njt�pJ��ml:����E�	�nqZM�'n���O2�n!�ٽb��ao\@vą57�	ݒof��ri��ö���u(�t�k^m���9�γʴ�Z<�^D��z��4���U��>�^��Z���N]�V���/�����]�]1�Jm7Gl�fn҃�9�+.�ie���g��	�`�p�M�W5�3;/��fe�I���-lέ���U�E[�.��i\�j�Ú$���[8,J5B�J8��'��%ܮC�9%�j�;�Ct�!8� ShaT�g;7��H�q�'B\�.�D��s#��&�{��XRڥ�G`�I�o!٣��ůU������Tt���Lǅ������d�u�V�a�X4��x-��/�ȼ��*����.��m��Y�׆��A]��6��W��]��������o�!��i����[��]8�#(S ��xk ��F�%yv�r�\g�����h2���5
�w�ث��hu���v�;�zk��̦hw�w:��?+{ںSZˬ!�h�v��v�<�^�H�o1VFw����Ɍ�F��zs�[|+�Eu6_v�*�I�Ѽ������v��q�ce]aI.�:PK�V����f���W��=Ɔ�3@ͳJp�RS�񩗂�ҫk��LR� ��̍���Sj�ڿ�|t�KG�mgj��k9ж�[�Sg��	s�"�1�R�dX����`�D��og��j[�)�Ԇ�%!�H��9 9�T��ΧNK�ݻXl԰���TG19Qvǎn���[���(7+w��Z�O��(���V�e,�U��ҕz�ɔ�I:�)�D}ڳF�CH�4�a��P�ᰈ���-� P�C�>��6�u罞�z+�CH���ۓ礁��y�3�0q!��F;�j!�]�ev#� \�3J�A�fu����ۅV���ڴ�+���v�X������k�isC��0�R���0����m=\��St*��ޭ�u�;�X�GZt*J��}�.��p`���gQ�9�*GBpؾ����.���EV��6�^t��T4� V�"�C�U�y�t)P��gl�fsiAg�b�`�ܐ�<��nv����\�����l���̗�����3hd�\��#b[�L�q�������PQ����.�)��^ �����R�"9Z���e���"]�\��r�*�l�֦W�.X'�uq��;�%�ƻ��ƞ��U�W�wA�E�-�ٹӛ�JA�/X:�	�Y�wwe�����K�@ {���������y�.�_UL�ܪ��lD�ӓ7�r��r�8�m�a�W#X�D�>�]�R��7��l�A[�"��jñ�ou�Ӈ��'���#c&9[���f�T
yԦե¶�n]]I����zsr�u�+)7�9@��3��4OzpoP�%�����^��& �[�n��Qj�� q�F�u�p�� ĩ;)�}�0j���R�	�^)w��o�f��u0�<ؗz0�]{����1�v�����;p$�S�gihm�J%ۨE/��E΀V� D.(d�8�R�U3D�N�,�|�#���Q鷛2���tw�oY4~e��E�);9���*��F��M=�}���'a�q��Z�����h1�f�]ۓCp�)�U��dKEa��W^0��>��ұ}��D�C�F���ьIв��x� �:)]tiS�/_vt��kv�0T�i�kԕ�/�	�wKwgH6�u��L8�Q��YM��;��a�)|����]�T�0�l-AS��v,r��U�ɻ��������J��Km�=�<̮�e��Z&��ղtj�4X�(;d
�v�����;C��'t�Z�Ve`�-�K�r�k�n�g`�����OV]�¾�����[钁�,�:+���������n=���u��ӂ�|�%Xi';��E#��!ʼ��sͰ�^N�|k��뛼�t�cR�7�.u�m�Uѫ(����ִs�J"��i�J�g�Ȳ]��6B���<����mXZ�Hg����'����x������H��L�aW�//��\�3�|���b��̇h�Ŭ�02�ton�e ���[X�$\�'w+*���u���sfG6E�;{Y���c�`��g��PSXh�˕�+*,�m��gG6+p��OtS�W���0N�h���-��]�,4*��o�l�6�K�vK�X�X(�H
���3������y)nȯ6��Ug�CC�Kkv��apb�ǯ��JX�����ukX"�����KM1S����W��d���\õb]h���v�껅Y��n��/*V$�ZŅ\V"�y�9���-�O"�إ[�շY2r�KްN�Ά2���,�ܡS�y(��(NN⡟0���1�����r�k���Y�eYMV��9�$�d��;Î*j�\�5�sѽ�u�J��2[��-�` �'��eݡ"�)��@ݨ`�˳^��(Î� 7t`�V\�����o_ �B�J�;�1�i�v9M�f%}q�,���i;Y��>=��Ojۮ蠕��E��G�f;�]X�G������޼/�C���u����RP���:7lVem��ͺ2�w0�I�Wa�3�E}L���YQW3�|���Fn���V��ᒊ������k�7�CWL�Gs�f	�g#EM+���zоih��F�'�x��),���h۾������b�@��#����ڶ[��Z뺦�
���f_����|��Ӭ�Ȕ��q���Pli�!��hfl�-d���@;q����=rV%��z��z�Y�4�q�᪏s�.w�I�C�t�:�tWu�
�36quiؔ��\Ы8Ƹ��5j��N�^or��h��Ejt�z�_g^rt;tlno`|�M��tyLy��=��$eo���8���Z��ޞ�aU�Đ���=�R��rpeLR�
Sk�̋8�"��������5��e��%�t�
�)�57Zf�r��h=7.O���քͣ#��� ����]����1hю5��=ܙчA�����ђ�Ŏ�ڈ]B��|p��ӗ#��$>)_>9#8�#<u�*ej�Ko��4T�^�m��;�����ͬ+d,M�*qPn㱅g6�+�2MU��=��iQA[��u�)l⵶��W��Y�qǹ��hm��Ԑ�u뜰"��@[����;�A��-�G�R��䝝��Ʈ���.�u_Ay���ǩ�/��z_֚W�W٬Ve9ܦ���ʽ�\��x9+"���A�u�opV�g)��3b�tf��+�uh�&TZ�t��m͌,u|¾w�������L��+Dy֏5�q[˕6�u+s�#��K�L�|V(�`e��D|+��[�ݨw��a].�E��]�["�陑}΄lR��y0�k&o��dP�3�J�a���jי���pd+�v\g��9�ix���}R�tBgP�z�Q	ũH��ˮ�H	��b��p��pn�^�se"6$ӽe6q�\;+�v�W[�.�KN��ӗ%\��f��XE�Vę��J��o:�{���Pݦ����w���`�r�.��u�eCϲ�U��e�1�&%�CY�t�l��0�B����0��9�;6��]�WT�����4�^�"���e��A����r��>�m���^�K�Z�Z��۠�{�G���l��`nr��c�Ŕ�����<��� r���m�!��g�D���ݏ���k����Q�Ǉ�S,�]���:)�:��V�WE#�΁F�vN\#�3�|]iv9�L��л,vmf�W��cRv5Z6a]T7�;���4��W80����WJ�]K��&j��X�JPT��o`�],��*���aV��b�;����I��;���Z�0vu� �.K%M8gpjfm��鵡�.�=1Tц🎃�,�P;=�b��6���X�Wc��1n@��Y��*t�����Efv�xl�;&��p�rP�mnr�>��=-��U�z��%m�z��F]�<���j�s�-���V�@�+�wK�/1��5'�w��W
�,}z���k�+K�e0� �8�[�E�}}]�ڻ�Ŝ�v"Z%����*0��x�E�-��u������72ּ��Όq�	�^»�q���r%zJuk�k!L�P��u�v���KJ�8����^l�K:��~�t������	@�tă�X4�m�vV��c#��ze�]�s%VZ�Ҕ��;yQܛOHu�ջ̽�I�V�F�%n���D��H�z�wЃ����NXA��3�u��;�~�5��g��ln��[���h�*ni�	�`�{�ZьA!��`�Y�_��XD���ؗh�;�Zf�⌥��je=+F͸N�F�+��)�iܫ��_`��N�Z�U�����3���r/];��/\�ʛv�W^*̾#w!��u���p3I��b��tvu��mvd���-��m�-��4Yv�T��T����=6X�e}zɽ����P6�&r���EU�h;;�8 {�����S{����K^%O ���ET9���*Z���nZ��q�	c�d�ԗf�%.v�+�n�f���׶V[m��f��V�dF�1
�/����J���SC�{�4���0�ƌa�4Lg�b"(V<�Ɏa������n��o��+g:Ek�t*�s���V(i��Eծ�նЬ��F��(d+n��V��bk�����:�)�F��3p�gT	`M��P�j�\[J���k���t��H��.�B��OEZ��T�-�CP΍��X�7���ÙYoم��](���O_oQ��`*n����Ó
#�ϸV
\�]���j w2�s79o}a��&�f�L�c{���^�w��HZ��uB����� =�+$I�����x�;+,V�.�lqR���6�Ӯ=@�`Y[}�&�����6r�#�i.�x=yCl�d��NY��f*�)����4e��nC��p �њ��<�}�%�[�iL�:eّ�F�S�Hf[�]f�ڵ�Z���{b���v�[�h��/mjZ�|�t��U+Zie���B�m�-g<��m�`Ь'��lk���G�!� #2�
7N�*�2Dn��ਰV)���sM탌3}3�p�S)v0/�]�U�����i7�="�Uڷۮ(�[vX�ܞ�xkmi�U��_n࿕��d��|1��Fs`�[�Y���	��d]��Oo�7i5}H�M�]��q�[}G�:8�l&��.�M|;w0�G)�F��)��4
�wnva.;ݱ@"b�Y��J�ӈ�Te+�e�\Z�`:�ɠ�vf<�'p���bb���V��l�6���=1�X	;�\6r��eә\i��8cc���;�}�Ѯ�,*�v�n-�+h���"5���)�^Gw#WX����=�G���rzD�D2n>�[�q^�
Ug�Z넍Гi�uKO$�#��'TۚM�O	K�*�励Q"8�LՎwT��2;l�N��ۮ���t�at�UgE��^�$5���cb�6�r�B�;}��Xd��*Ħ����W4J�+8�fL1*�+�L���sJ��7w����R��1��� �/����9�ɻok�+a:=�.@�T�8���cX:�L�}�;��s��%�!��dS�Ex���n�#�@ue ���IXC�n�p��Y��F��
-G9��Z��&�������xv��N]���z�n8�r���+��O�3,�Tt�ݬSV��iֵ����8�&rv�c���q�N��Eڻ�����4n
DN�w�k*T*��M-WN�[��-�N�
(Q��v�#`F��N2�غ*�|:Nu���A������#��S�
�
�l<�]p�+!����:cV
VQ��q�7��{\�6 �u����ڮ��5�5�D��Jq�u+�u9GDܭD���N� ����׫���@��Le����a��={;1���=n�is�>ψ;F胝c$b|�\�X����$ۙ�]�3Xwq�*��8�#P{�tnM�i�d�ߵ��(7�v�=��b5���!p��r��Ka^��Jݧ��T�[��.�����Xu���L���t��[;�}۝��w��-��MVn��9��؊��3mE��{b7D�Hm����!1SVw+�c��j��l����P�N�`+�&q��p��d��d��S�V���I[�ϩ$���踉�+�-ÑR���׎-�MX#x���$՞���nVp��B�[ha��8X��rq�G7�=��+`��m�W���x���J�n]*����Ţ8�Ѵ�]�s���h��Jw]���?VѨ����O*C����8�H���v�r�*T�Z1�2�Ɋ���f(^�$DG��}y�ڋF����Q��ب��p�1�Ԗ�{dQv\����ӗ��6#/�O%������ ���3���'��e�c�՝�źK��@r��4j�q5�@Ց����Q�ђu��]��Q��B,�MМSԩ��`�-��m�J��P)�h�a�ŇC;Mb�T����m,[�Y������4��7j��gVe�p_�6�V)�f�oG�Q�͖��n�yb��R�#��뇑[ʥ]ʼ��e4J�gSA���u�9�;�5���:��5�/R[cGaag	a��1����wݝMَ�uٙV���X�`Ċ���4;zgu>������UԜ��������yt��v�W2m:��U�9Q����R���Y�	u}�*��-���[)��^A E%�m�c�ά�+��Y8��I��)�Jw���ྫྷ�i���akf2ZB�X�-��cJ�aR=��I���#uӮ	��c��:�a�2	Z���_�mx�X�#����F0Y��`Y��^Q����*mB"gc��OS��t�r�2�����u�Ϗs��imKV��WL��+wɭ%��
�vrˠyKj��������*�8�i]LH�Ş�y�8ƫE��%mG�B�_m�	��%M�;e����$9e8gf��+c{:a�Zʴ~�ve0��)m݄�"��9�w�r�o��nA�6��mm��V|���J��Yw��K�ʱ���2�Z-�W@��L�Olڝr�ZVꢫ��1���6�-u������]��nlJt�e,���7��[�Gy��+
��vX����h�mN��hظTcUodD�����8��]��ʲ�d�����v�dP�XHo#r�������W��h�bn�K��K	��b�N#;3k�����R��}�":�60��{w�`�U�	L]6����1G��m�]L�in��j�g;�G�������;d��2#x9�����@1`�J��[Ţea�p�V��5���9��fek]U�A�����Wu�R��Z)`ڼ��ZBJ����+�
F��:�o;(��P�[�{K�\�����,���D��������hںfpJ�����O�i��=�f�l��1�r���J���j�����
�g]����A�q�ִq����Q{�e/��.��L�����<}�;H[]�=��6�J�kBG��Z����P�(Y��i�9Ppѧz��7��t~άV���b��Z���}Zo��3�u��З��2��ST�*������̩�{5N(���t��r�[���(��kw�Ht��E�t����2����R�4�_^�x��Yw��Cm�m�E�ގ|Ӭ3���嵀�+j��l&�r�4�Z̑���M��Bh�(�������&���Ioλ�͎#��wN����UԺ��ī4Ґ�����Ec����+GJ�rx��\�Z�с�u8aN�t�u!Z8Q��rѕ�M�;-��z�.I��yKD��$����ӽ��Qd}��6p�V�r�.��Y ��6��^AS;�ܮ��Y�c��e��4L��a�j���N�K8%��|THZ���#�Ɍ%6!}a�����]�X�#��W4�	��Y�r��Ee>[�0s4<��Y]���v s+�Whv���daee�7im��h�Q�7��Z�/awz��\w^�r��N�z�� 4̥W��K���-��}eoqu���(v�6���ћ�c���{� ��>��w��\F[V"ڽ�i��D����pF����;&f�n�atO��=��z���mDJ��C^h��x�����n���vT�-�T��
YP��6�x{��v"�4�e�塨�s�f��9�����}N��ˀ�7�i�z,cT@�ʛ�D�M�>	�Hlİ�Y*�Ds<��oe^�.�����(c�D��Op5���e�q�3h���k���/a/uʒ��M��t�O>kF�0�b�^���B�=��#�GA3-C����x6��T��Na�E�����H�:�lY[�!T4������K"bӏ�,u��u�(#���*5]3��Y���.v����m]���Z�RXiL��)��3��b�pv��=�	����!�!�{�kx�R����!���G�_�㼣�ӃC�I�˕�g��*��WK�z�,7������<� m> ,ٛך���6�,�[��]SF�3�v� 1ǯ�<��3i��%bɣw�%m.Aa��a�a�,�aR;3 Z��{�;0 8�ȸ�ٸTˀ5���>��a�U�2B�ug�;� X(T�2�5�2����0b�����鬲��P����֕Q^�3*#K�K�P7�A���)��n��wՈ끍 K�J��ԯ9��;eEpC!I}�����/����:�#�CÆ`��G�1�2�l���/#o�_sﷺ��.3��;�w[����=м钅�Y3�9��j�����5{��u�[���2h7Hұ�
d�@UAKV`��AQ41�D�J�PR4�)J�@R�eE+K�HU�dІBTI��SE.FYU �8N@VA@�)IJ�*dH�P�P�T�d�d��Y&@d䡐9%dP4Q�9FT�%A�VK�DfP���K��HRd��f	fdBd	���Pa5�R�BP�&I��C���5IBd�Bd�=�}����٭[ן���^�N��V7�|PU�(Áv�u���������l1v�6�������q��R�R�*���9�Ϋv�rJ�uQ��H��{��%^��V)��]�5��ٱk���+�P$tzݮ�f�����l���}!�@����g�Z�ie4�۽}�#w2�Fq���ݨ�Z����/�AH،�j���U{e�Ú�L]��:&�B�k7�q�Xg��'ZNA��!���TC�V)/�E��x�xصm1���\�3�j�Z�P
�`��i׽b.������,��G)������KF0��n���n��|�ƶ�7g5�#�=So�6"�.=��u/)rU��eړ�l�u7��MC�d�6��ۻ���V�T��Xq!���kM�ڻ���f��X�&��V28��Y=Ӌ7��T�Rㄾ��0<8"s)_�2.�P�`�a�)or�ģ&-wn�:��f�Z��{1�&��O�Gӎ��� M68iW���z{7z-HKvd�p����z��PV����*�{��yٻt��V��]sr�K�}��v9�nݨ���|Z�|�딪^s앹x�#c/ZI!��N	7-d�����&6��I\	�`;���$3�F�����-�qؕ��Q�:8g$�4V1���cT��7�w����!ݎ��ٳ����b2g�I��T�siN�r�w�ݦ��i�<���I��M�Y]��;����w=	9Â��P�,��m��-k�M5r�;��t�R=ѕ�V�e�Fa�9�,R� m�hvRuz��&��E��kh�=��;/�z�<��OD���p�X��{)uu+|jq�o����j���'���Է��M�w{6WsKsu�w��5 �N��M����R����/����\V��DPAH^����a�g-��H8�o3�4���Mߗk�TP��9�iփK���C�<oReb�c
C����R+VΥ~\:��]~MUzZ��C��5��[V���IwO�^a%��t!��r;=Z����:v5�}a�-�o��|b�0���l���)��� �����Z�3w(){uf���U����pF��k��[W��2���]v(e�[��mw|X����a��}�,>���Ejn=�e>�Mp�3"�c��`�z����P�� �++�N���r̒�m�Lη)��j���D�<3�gE���Mfm����7�M���W�f6���FS��*-p�c�a�����X'1��ݬ�tɃ+�p�wR��{�	uw+$���a7��p�:�huD��a�'2��ki����#��ow���*�a\5� ����kk�]-61ޓ^�`(&,8�f�v� ���n{w]=�\��D־����<T���	���w�ׯ#�/b8��V�tr��֣$E��d	º�¨�}b1�d��-Өy۽�nv�Noq��;�,����A��%�ʇaHl�Ѝ-��)ম��+�b��ݍԝ��\��1;}Ǭ.� ����QBE.��Ѯ�MΩ�]ת��('������u�zS��ꞯ&��>ҬF�����KD�;ڑv��r���s�p-Ml�����E�
�`>�dS��u7����y��+�а�&*;)lݠ��W��݁���u�O,�L�Aƭ�Ŝ��C���сL�1N�r�:�!M�/��`WM��@�w��,@"Uө�w�Y����������V���CL�C��~�Y��e��_2)��l̰�\��! -v4���}�#PR�h��0�u�,���ڑ��ʀ�{�ڷc��;2���eM����)�4Q.���ە�j�-��d9�M�s>�p�����Q�,V���Jn-��+�X���1�ǹTOEwh�n)wzߝY�C�z%�3��1k
�l>�D�N�r�
-]OT��=�Ձ�R9KT�{}~�b	ӉH2$��3'gz�C�.TLu�78��)��r�2���`sv���AS؏E?��<"�誗�����-#�U�@����xէ�q�ǫ��Ic�Ȱ�(�nO#"c�"��_.�J�V8?���AEW3*g
y�Zf�ֶ�e)��ΰ�6���Ȅz*��X:W����dh0���Eo%�)ז�[��h�)0Ηr�Q�T3��ݷ~��7���b�t�F���1�٭ޡq����Xv����NT=���Q��恑�N��Ȫ�N6/�зG*�穪���a�����Gkb7 �QR��L��FyJ�:k�ib��>�QR��	��Up�8�lh&�$I���7��%�-���0�m�!NR]�ؽֿ�S�8+�l�����,��/В�&�a���K�k�ŷ}Ks�c���Of�����U_|�^1Bʬ����5(��3lIɜ�]���PM�<4gn=��w�X[42�p��	'�����{ձ��b�S�W%B��+�h��"���ڶF�w���\A���N�D�SV�Ф�{����Q�>
P�L�����k��clU���
.]vQ�6)	��v�.�u[[�Ѷ��K�6���GE9V5��Ϭ(V^����S��x�Jݽ8��g�^\��\m9�z�d�ӱ44�pc��u�r8�� %A��#��S~��b�D�Zdqv����7����E�3�\"�T^B��v�}S�w�gOՁ�a�Q����]KJ����`����P�ܞ��paH!zz��)]P��TTg������`�
�5|E��b��;-!9Q����x���h����YH���;�S�pD��I}	6򂗼7�E�V��h��κ�;u|&�c�0����uk[h��7�k&�eVJ�턹�MoRR���ҸK��	ߪ��ǔ>�.j�`_2�=��k������ë6z�WZ�f��@������8���K�	�L�e��� ��B��zL�=���[��"�Cn�>ɓ3�Ɠ�D�3u�;�ٽ)�>j��}ݜ�����F�j �v�3zp�כm�a�ռ�0��λ���f:\-��Pyt�l��,+כO��5d��B�ح������V��q�'�]R��cN�FyrA�c �!d�Ѹ����f<X+�r/��bӧ1�2��1�"�2��{�e�1'ni��T��r*���FCv*��v��FS.����y{��a{97	KW����.L{�:h��s�[�L����}�Ԋ�����o�fux;�7]92go%���B���p�:�������W>J�	Co᢬�,�3�YiNJ}��}��λ��v�䒝���%!Ů"��Ԋw�o6-���њ��=~ñ'����)��t��b'��ʺ��Cvvp�L��ޓNZg��p��^u����@mz�Y�%nQi��O�\P�������dh���兩{3����ۏ(jm��Ê�����asq�y���y�lL|dO<d!��]��r�z��" ����rUm*+ubW{���E�����d;��}�h�E��}HTWM�V7:e�����kx���};�9n���RXj��������(ߓ..�_�8^���K� ���m�9�`�i�}u�W�&�\F�M�H�,)�͵�:��^Qz�C�z���UoV����}���H�ջ�6�	㫡��+��M�ɨĖ���1�0Z�o�fc�T��Z�4N�0��,�5dm�Iu�l5�Xw�`4�9ɬΠ9��f�ފ��9�t���z���0V�s�}�>?M�kI�x��x����¨�˻8��D��l�F���WR�����J���jps*���v�g֝V��� Ҫ�\^�/��mΙ��WZ<>�]wGUe3��H���dp}F!�r�B}я��tq־=�J��hdG�'
[8}e�����H��1��[<.VčE�P%�U��K��k��j;�KQ�'D�t(�!>'�|]"�k�PXc�?)1�.�\���n-�{s�ƣc���s�F�B]���h�
�/دT5KG	B���i�)��Y���9�ʓ��(��r-I�
_=���s0}n�`��d��s$`�X*D��4lV��$�n����������\�6xt�!ׯ������
�Qn�0{����R5k�͛�tK��՜��#J�x��g?�>���_ݯ�<1H/�wj=A=W�:!���9��o����\ĩ��?!%�4�g��R��nd��%���E�0��u�4Y��L�1ƏT�+�[ݖ�R
���{�-]-�ku��7MPc0)m�*�jf�ـ@��{��
���Y����(t���j˺g%�SQL�O�ݏ]�����\I���L�¨fk0�<����-S}�cۀ�%�_[)gr�5���E)���|g"�	�3a ��
�J����i�}0��շ��dh+;��[�G�aa:�ަI��r��r���eP�����^�n�MCOE�H�S|-��$b�Y�!����A��Y���,���Q���<��BuQb4�U61u�7���Ѫ�,K�p(vs�4�܎L
��FCӡ���l���W|�w0��4.ڋ�Z����%�r_�����ʁ~�t��v:+ɝ�Qoz��֑PF�J�I��Y��Uu���FDF�E'�:�aÃcg��Fy,V���Jn-�����ڥ]�dvi*�wF�F�L0��"���H@�3ʺ1�T{a��K���T;GdeU��[X���a��~T��Ԝk�S����XF�Z���`�Cɔh�܋�ޭ��qC�̕ˎr���s��s��d�ܐ&9�3|%D�h:������Vw2�8|a��?N��XfUl�ҢԱ�u1�l���fd
־*�ix7�ұ�wp>Mncc-��ub
��N�+�k���`L�Y���z�QO���U�8���ӳ�u�Sc7� 1Զޓp��%M���SClvs�:��g^������*��Eh�n%�����e���М������ʎI)�0����dw�2)O�cj/�P��5|KO�o8��h^	�Kƽu��70��,2-��ʜ����z���R��ޙ�s����Z61��V7i/v[>?ET��_�z��k��AE����r2z�=�O&k����e�W�B��d��22)X�ȫe�F��B�-�@;⢜�(_H��l�;*���v��M����8(���E 2W����8f,qoW�*�,�\�AOb-�c|�T���Z��E@���+�D,����SJpl�Ua}�g�JE��?DR8�ʑ��i)ڸH.R� �P�� KE�,��Z��f��X�yJf_�ӌ��:���N����xxXǖ����q𫡱NV�E>��
��F��dlbĞ�6+ݍ��[$����ح�/���	�2�kK�+ݖ��yM�m}H��WH쬚��/�TMn�Z�O��>��*2���5�HQ�6�ی�_��qy������?�71د�d68�S�]���콏_�5`�y���A�!z:D})kt��|�A5-'ݪ�Ǜ#�`�{�v63!&����ˀez�x�-���3�+ Iiu��U��s[/+�N�a����yB��^��E��U�.D��o�P�5]qg�.n��6J��Vk}�vřH/:*��L������t��MW�za��	������V�ȗ�(c��f:
��vV¿7݁�A��m��?����
 ��/�z�qs&��ή�"�l09�����B�X�@:���N���_��P�B!P&6uL#��B���H�zwuZً������s��]6��w�.�qa���)0pO�#t��o{l���c�O]���Sy�}{,|���L�~	�L�e����Z��ؕ�&�׆O�ԣ4YlS��2!d��q��JP�x�V �[��n��;J��TkW��zfJG���ƞ_3�x��5�(X��Jo�
Nv ����mZ�j��}3�,���܌��5Y���/Y���P���}�%��g>��x*�����C��ȕ����k������9�}�p�7Cb���w6^r�x�,%�d�a|MU�W�.�i]�m�=,/&6oӅQ~\E9y�jE;��b����3ׇbO��'hf��9Z����e���*�N	�b��i�����NEKκ�}��>Ͼ�4�B���{)��;\���;5�n�x��#7R�맏)9f��4�>���{7|����3���Ձ=r[87z�*�z��X�sO`�,'�]�U4o@�q�{-��t\^����"���|$�*Pu��{��ֹүt�-1�q5��4m^���r�8��(})���W7Ql���qQvAQ�u�ۡ{C�SN�R}~����tk�a��>��M�^S4'�\vͭ˾��x4>��e����]�:Vᕇ;���R�Wxq{I��y����<j��`漝��̭� 0�x��w.ɽ�f������YX�7��o���3�)1 �NZ�#i���X�/������[Zv;w&~�
·��r�o8�͞5�{]�~��f-��W\b�Yy��Ԭ���r��	��QX�U�VN�Wӷ,�Bڙ2��ݛ�d0�j�'��*�	f��͡A6w^�M�s�v�i�V`m���}G+��b�+�cR��`]�bo�x��閪��2���ҝ���'E�f�AGX���qLnȴ�΃/\���jKLƦ�r���Fy�mjFfn�\��� N[��ʎ_w�k��x�J*9��k6��P�A�ա�,(SF�,g��HL��U���duui��&��K��;�ݥEV����t:w�4{l��WR�U�bEOU�,݁Y�.�L+(V�N����)ۼË&��D�}��ڧ�&��(��He�Er��3ClΔ��9�4h[�3/�&H�&52�1�gi��v�R�[۬N��sW��K}��T�:��c���&t]�-]s��Wգ��3y'cO�c��T4E�S������h��1a-��nc�\�:��ޔ�ٔ>Rp�`k[�V�cT�SZ*�q�ݭ��*<+��v{Y����(l��	�3):c�r��Fͬղ�T��@ǆ�૬�&�B�A��[͕���Si�y���c1Y��>W�ӭ�Da휡k�FU���aN�U�=�BB���5�;��Z�s3�GoZ;/��	����ͫmmY�*0q�b��+_f�蕧��妑��*�gSfdL��W]$��
��ۥ}�(��whǑpTe��ۜZ�d�����=7z�N�l��k)-���ދ��	$y45���{�6G�[Yf��$����V�MԀ��,;�-AY�gdH)�7Gґӕ�ϥ�Z�/e�D���DmOo�Z�D��[װ�Ӫ��G���-v9�ޗ�ݵz�
���`V���D=Y�m���Dkyt�K�����[N�/��L��3O'P�˜��O�1Lڈ�i�A���W���p�[*2�i��i��\a���&<E��2k��G���v�i�|����[�o��,J�i�I]@T͋^r���b+LX�|n�>0G�R����K74upRk��_n:�9u��,�s�Lir�YTME �u(v\�����^���'O��X��t����Nd|�o�t�����ф��r�.���xD "h?4�&@c ��������IHPeF@ef�eT9��X�F@�2�Y��R���QMU�f!��ХVNH�T�YJd�#B��9EY�eDNI�14��E.IFC��M4E.T�fM.@d�!AT&FJ� R�!FA�QINA�Y$Q4Bd�1U4DPى�&DIA�Afd�N�5Hd��9dQEdP�fMS������4R�U��4�4U(d����@R%4%a�SU��HҔ�EBQHP�H�cKIT�@�4�T�M8_@|�r3����f;W��%M�3�S���/9�/�_?&_�nܜ�Ӳ�)�[��W�s�)}}LWL�V;sM��M����T�=��t��q;%��]�(0��8jf�z�w��ǖ��X'�v��7gDZ�|Œ��N-�V�*u��C��Q�������Ev�Ձ��ʒ��Yp���7�[Q �jtj�{�'��f�<
�G��Lo�B��n½Ιf���WEYt���"��H�B���k�ɶ�B�3�1�O]L���pJ��u{ı	]P������f��V�/\rSu���T��\q�b?k��s��}�z���A�󎌮��>��}wF���j3����tWZ��ɞDVt�P/�q���9�ͻ���ܟ>���z�U��Jo�<U�5�v��z��2��Q!�]��ʇ����Z���q��.G_���e��rT�nѹ��Bo��@����4ok�&�B� 9��+�r��+Y��(gm��>�Hgd<�HZ��): ��A����(�E��JJ����8�1L�}[7Cw;a��Vv�S����n�Ⱦ�NU�_�n������K1H��@^�si�:�_�'*�'9�mq�$V���aZ�A؁�լ��}Y	�5�`۹u&���#�����s�e�b��U�{2��G&f�j�KW9�gn�Lufu�����%�Z�	'{�S���L#�wҰ
^79�ev�S���S�H��ݗ��{z�c��xԼL �9�.[��tv�9״ɮ73��=�~���w�chz�>ɉ�����F����V����usϥwN�= �B��0hi�ci,Yl�ǭB���J6F�a�Q@�v�T�Un��#
�s˩�q�An���'����UU%8Q�ι���M��2�.$�aO�Is@�/(�R��N_��+�4�TS����S\S���B����7�F���/��t�O�!���Ӛ�a
.��Q��&﮼�].���h��C��.ӟWN���}�Y�Z��w+!�K�#�%��^�A��2Tij/�7W-�z�X�m��B7C�>z��Zt�^Z1r��_j�]C�H���q�9w���Je0`q�V��#�\]����"�L
��FC���]J��rQ���ނ$^Z̮p�=�á ��TN�W)
6�POt��Ca�veE�5� �p�mQ�������Vz������
��|���j���~w����ʞ�'8�
���b��R�8�;|�u^,��ʉ}3Kq���O� >��'o���J.�ܬ7�^�4_Q,�
�1I����W��6A�P�j�Ǡ��ğm���GhQ��8��
�wu[��DSmu�y�ڰs5ۜn�P-t9
������If���Y��1�����z�h�z3���岚�����|%v��v�:��G>Y�X��lpӫY��ň�qTu���p5N$E|��	���=�W�o�_L�9����a����>��.t����>��s��d�ܐ&3t��ehZ�R����^r:�z��'Y��)�n��n��fP�&�u8�8!�0���Se��fd
�}'�qX��*3W#�K���^߳{TBc~K>[T���m�`kl1l� �f�r�=��QQ�ko�������)���؞�|���}�n+�K�;4���/�ޫ�r�7O�)�;(��u����x槦�{�r�[�k�O�%���F�>�݇<�do�m�n�0��Ӫ��V\�z#�F2��JӐӷ}ӣ�_I���9�p�2��	��C�>Z�פ�Y{yC��i(�B�X}W�U�-S�
o{�9^�|��J����3�2����d��3D�L�����O���x�(\��١M�l�Z�,��Q�����:��T�d&6��c��X4$�2oh���t�oh%�'n��uM|��ᣵ�s$jF��ZT;��ý��=��dץ�H���j�wY�.�L\�u��ڼ.��h�ӽ{fr�0v�L��G����l��ؔT�Q�s7�X��gkI����(�Fc����}Y� ���]�]N�R�g�����([}ABEҍs���(^���w����i��'c����b�)Z\(1@vZ����㗈��֌����UyV�{$h���B0��buV�vz�|8�������y�B�m��g�����d���j��O�M������AJ���� ����t�K���D���t�>�p	}o7;[�Q.��T��g�T�Se1=
�Xy[������Y"�����4�ZD�)��=O���v$�f��<�В��9��AŮ���̅����#�'W�j/ю@(K�!��}��]yc�8�AClwV��ϋσ/yO�@��\���ǥ�.̓9���Es^Z�Gw��뇷_u����p�i�C�F6M�@�μ��Ë����љ��b6yI���c�>�E� ��a���V8_6��"b�u�3)A��x�V�܋�r��LL�1T�7<+t�ꉇ���7������J����pBŏz7��';��/{�qy�&��X��4=��k0d�9lն{�����#�V(� ]m�H��/w�(1�){p��|}\�6#g\5����fo�>���;�~�q����w�U�p�M�I��[�Ը�x��W^�쩻¸���*㬢ł��Z����b�:Ҭ�C���� ���p��{����N� ����{}}�/ܮ��%CB�0)>"��a̽��o����<gs5����]?^�0��zX�e���Kll��n���ig�CA�
����PG9������[{�`���؏-�e0Y���=m�ņ��GF{Yg�ĨUx�jޱw|9�x��H3ъdP:iH��]�\.��!��4�r�'^�`�NEKα�<�����.J�X/;�i8���}cg"�E��'<YP;$(�
"%Jc]mt��O�9�_��Jd�/�U��Q��K&�*u��h��cUԧ=mE��+�>��w4�< .���ϱ]gT��T����XM�@�!�@T!J�єuX�lRж�/JgN<I�1lG�Tkӎ��k�T�ɟs��t'*&;��e�e�ԋ�G�ӑ�	B;�����MN[���P�Gd�|z�58��Qt��g�ߺ�u��2;$�,UuG�p���۞�ybw}\<Hg�4����J��}+�P,ۻ�l���d�'�sR��;]Yc���zL�c��[�}���Ѹ��/�	���B��71(��,�����i��6⣲y]A�w��
u�|4�0	y��r"�omq�b�^h�1i'+�X ��B�I��pN�ur�T���!��k<w����tZ2�]������ӗB�U��a�F�5�����x�R!�ï�{]B!�����g~ň��������7%���y����9G���@s��x�GGt��ͺ�1�T1u���6r�
������9: �:f���FQ�.�~5�(,1���;Itf$e��q�� ���\�����LPl�"�f�jƗf�ER`����.q����(�S����m����"�L6�M�����"�:_�J�ZU�����W��9q����\U���gT�	-�\��4�i���5��yt9C��f٥嵗�R�����S �jz�=���4�*+��s�;F����(C�����s�E;�G�	��R�Tl�34oTU�1C�څyaZ�_vF��$���H�Ӆ'O�V#N^lY��WS5g���hCm	�R�Ot�Vu�L��d	��W�M)� â�.�T���� 1m��uI�͸y����-�g�=��E�$�I�X�']��d� �"ψ-�m���E��QG��4O=ݺ����5�+>����̷������'a�݉;+x��Ȏ!�[��L���:�XOR���K6��1Qz2��.���|Ue*�N����7���ڝ��]4�n7upJ8�<��S��|VyN�ۧtL��9"�|���x�R���m����Q~}μ�X�	��x*�Ky�hbP�����#\����:u-B�ttA��И�.�S�m���P��#!��ThM�T�GۋR���(�啢�9F\K�c(�zH<z&�f�R3Ѷʁ`;;�;;2�	Ί�*9�bB۩~\EA�AH�\n��;_m(Ea���GvOH��57p�>՗�yD<�blt?k9ߛ�����J�r�|e"3˥4��k������X��V5�ʞ"�hl5J2*���؃�j�H���=X�ݮ_n��G�ю���;8�������J��P{�j!��	Ӌ�P��
�*X*5mP۔s̕�����񯳫�@�ˊ� �eRl�q�p�(�ry���3�"��_,<f_cӏ=Jw@���V��Y����� ��nc�[!�>�z0��V�5CN�	ոĮ�,F�@ !.錐}6mJ�G!��V6/۶��3OU��j�T>���՜b���+�fH5޴��3(QW�8T
�$�<���d��燦j�*���jN��7}�����d��_a�ȸ�l���Wt{]S;3k�T�f��N��L�,���D�񑧋u��{t$�5.�\.��Y�c��H�����P��� f��,�7�e^,�� ���P.�8�W#�S����O�u
_p�t=�hՆ�J?����{վ�������4	���Z*���S��j�,��t�
�1�""x2.=<,����_dx0t1�cFN��wp{��XS�ʮUy�����v��Ҝ=3B=\$(�g3�oi����˪ӪX����N�p�f�6Sf�"�8�	dvȿ%��<��i�7u�nu�������gWy!��z�0s����;��p0GC�Z�v��K*1ͷ�1Zk����r�¨x��Zt��\+@�"(aq�b������q�ŕP=��W����y�c���MQ��0Q�з7-��<��1��FPS�F��!G��;��(�������=�lc��u]R���'7��� ōG�i�aH+��˄�¨VԺQq�ݫ���-�l�zМ��z��!�G9�V�O��S�x���5�ƻ圑1Cg®�d��\eֈ�͞��T?'�.Ԫ
/ˁ�js�
.ĸ�t������ME�9 �$FZ�
j�	c�n9H�Ej�hn�5"��/�T���K\�����E�%��G��:f�"##��+vq�e�5-�mF_o-�+�t�YU�$+ঊ*s���$�e-�0�ژu�)h|x��
2r��d7���L�Jι¾+��� eu�λ�Oڣ�c�:LF�޽>������]6���T8U.42p��y�|����$rɒ�Drs*�O��r(Iڸy�0�n�Y�q���qz�Ծ����})�\7�jM�޵�xE�~r2$��k�)EE@�PL��@�EзJP�x�RF��]��~N�㣆n����q�~�J&)��l&of�j�Cƛ�U�=�T����,�)uQ��۳�E3�7���n)��/oS�y����&�<-�����҇�Hp
��Rxj���i���	���W�nUr��=�7�j�Cb���lc7�QW�73���W	�RG;]����:�b:I���/Z�OQ�ಘ0���!�
4-ߩ�ؿ��GF{Yg��;`���s�����f%�r6��2+�M)d"6�8완!)�i4��N���\'"�c&z�n"�Dt��n�k���(��Ѥ�\��t�.T�!@Z]8k�0\��猲3�,n�f��.hH�ɇ֠�JvQ�x�Lm>>�-�X�"��!�ߝ!طe�c�Sn�Y���`M}��3��J5�S=��&�5��j͛����-���*�2�bNؐ▤��<�����Y�7�b�=��C'=|�,���.G��tҨ9tێ�s仪U�u�l��%��f��&�r=%���d�[qM�EM%Չi�ɺ�� �<-�PьS��6���7���w���<8C��C��(�)p0�!�9^Z�s�f�w\uU�^4�����U��i�
�Q1���(�.*�Çzr4B�����)B�q�ml�
��P���:|v�s��nEAzv1n�ɝ����&)b��0D��C7��5�:��0����JJ���<����xu��]�f$>�t� �x͌wK�
QwR����|8|�@PD{\�F�"^�<=�G�M7F�g��۫�>"��u�y�o�U6bB���h�i:��b���t0����[)���YY7֌s\{]��a�1Noɟ6�ᐬ�t�t���б�j ҳ���C�r0�n����㚹
S��5�v���X�	���ϲ(&k&�iqFhpdUy��Gg���EQ�T#1f4�3�I�����E���܋����9�.[���w[ ��^�=d�
��q�ө��e�$Z���Κ3�7��R�]˶�:w�!��yכ��~��j< U%
��*}*+}#o�����_A�Z;�<i�%p���]zF�*�]U���FL��s���W	�T�q7yVE����B�����}��ÃN�f��*s��8l�09r�����Rvo>�:�T�������_k�Y.��Ix�����p� ��#]���ˮ�۝z�4�f-���I:VButO�7���1��&B�n�g��p	��$n=H�'3y�;�*��*�K	#�1��;XRR�x٤�g_ܲ�N&^�]�NK��U@D�ZtإH���C�a��2������O.w狭��2��;a�찪Bg9\;uȋ�1E0�Y�����unO� Z�η|��&�L��ٔ�-zF
��Cз�[)�M�v��mYg���&Xڅ��֝�r����;���$��J��V�]]�u�ۮ���7�` 1�Y9T]����l��<ch�1K0��+dR[/6��g q���ܲH�>`,�)iLN��^*ztݕN���ۖ�+��2X�V-���vZ������4!P�K>��բiht�]/;Oi�s+3�q�Kp� �vdj�֥e�#n���p�KJm�\�MΧ�+z+�YN>��9��t�m}�:�Ā�4wn�r�dbrN^�Cm�t߹����x]ߞ����ʔ��xDB�[�d��5�Ӭg,$��$���]5��X�\�5�o�P�ǖ�V�:��x�ޥ2|���"�ΝT�I�R5��4pa�.87[N�����r>��]X��AEO�-jތ(������� m��+�u�:��y:щ��o�����6�b��έ%�iv�h�l��Biu_c넩���;�J�%���i:���qi�V@[W��R�w���w��Q�;��l�B��W8R��I��Wc�3��e*J�@�uMe���o2�fĻ'NI,R�vKv�|hݾU��S"�3d��H��}NGD���_1u���
K��+��O�Ez^�N[���T,��!H�3\��ϵmJ��4��F�I��J�G!�x�`�]qѢ���32'��*��e��!�+/�Y���wlW�u�G�o�4���=��2�uї��p��u�*�	x�ke�=��'meժ�V�.5t��t���~<����9fU=7��6�+M
v�9��4
�ѳ6q��$���g36��6_P\�5��7�U��]�{��X%`��*����k�IGXBc��.�YqXE�|rWc
��e����]�
u/��ޭ��X�
^oI�IQr{��t? ��'@�^V�PKV<��n�ܻG��:�=�^�e	p �`�[F�N�U���o�w`��ɮ�ҫ�T�M۩z�-�w2�B�6:����]Y۷\"�Ns�� ŷu��	�\20	۪�KJ����)��dv�uݦ���Գ��>����X�[�oGn�b=9oWW7}�E՛��]��+��'��:m�ͦ�jQ;���>�ٌ�;�gWS�M �\����7�{��(����PRU4	T���Д-D4-PPU�FI�C��JTAQRRD5C�QCd�eJT5T���AE�ATQELQM%P�BD�U!ADDUET�NNE4E@P��R4&A�HYT4�LQIF34QALENbbHUSM4��JS�E4	CKTCSP�3�CMTN@dD44ԐE5UUCH�NF5P�5MQE4�PRDP�AM�I@UDQE-,�U4UL���4�4�QRRUPQUBS��PP�A5DSUIPL�DU-UEQDTAJRETM%�4�1EIAMQ4��9L�S-D4�@DQ@�AAEPSL�A�K3��5��T~�<��W�������{�}��V�Đ|�\�6���^�����Ww+�(�D�d���M��j`X�C�ح�9��}��|îo�ջަR����UCN�gϖ3��=>{k�8��]LC�8�Sɺ8*{�¹u�j����*<ƵY����A�g"H�|pI���>F��v��8��91����!�^e�UyU)�u(�8*S�@Kν��3�zϲr/�&�ѐa���y@�������z��u{���osG��q���0�4GW%ȧ�?y�pW%�vs��C���9����$����X?�����ѹ�mC�d]��5!�N�¿A��x;�nNsQ�}�ݎ�c<.�{W�d��ۣ��"��>`C�9�.℠�~�͏W$�K߾i�x�/7��<ϵ��!>�;��rz���(}�_����_ms��4�ɗ���7=����.Z��o�Fj������y��?\���aBPP� ��8��nO������:��Sֻ�a���G���>�#�:�W�b��j(��j�pFA���t�}�P��5�=�.�2<��ہ�ȏ��|��U+�_jq? ��l{�}�p�MI�:�o�E�`��ހ������C��7�t���5?�y��9?F�*��Rr7�dS�w�ܾNA�뿹���"����I��Id���͇��_��/�˪�p~��:��b���qIԙ���+p�Ho��aK�=�#��ѫ��S�jM@Q^Kۮh�J������pL�Ǿ��';��r5��1@���/����C����G�Tj�<�F�)l�sA��	{���4�ry�&� ��4r;��u'֬�"����(u~��5F�u��/7��vc����_���r�}����Iӡ�Tc������#����Pn=����?{����L�/�a�.�&O���sx���	C�05u9����:�	�j�ˠ�
NF�)ճ�(7>I�C�`jO$����Ă����	[��9�e˽���LU���-�]�gu+�6���,8QoR����+���W�M��ү.ֆ=o�W,
)h�mS�ȽU؈��)���)1����զ�]�]���BͅPx��Q�G���ϗ`�w����.��5����?N�޾�������O$�}��&@j2������r]K�eC��=~�A��y�t~>��NI��vޟ������5UC�3���;�Z��H��*G�ǁ��Pt��ɺ]�|ݜ���
:���j����'Ѩ?A�]�:�ܿ� �t}P��zu����5����P�����~3��Mɑ����]è2^�sN��RrOɭZq��r)�9���{�f��z���5��~g�������cF�(w~��/s�`�j���yF�ì]O�|�G��7%!��������Ky߾i{���15������T�szk��Rg9��u���w����������s�=�.���s�}��o�>�dQ���X�\��~�FK��%;c���寱?u��?I�%���w	O�����y�%?��0<�#� }n��zM��~���?8�K��p<��>���5��O#P�ߚ�����2(;sC�<�#pn���.�5�)�L���W#��N�x�(?C�P�upd�_�����1���1ﾃ�2��}���UcmV�����>Oy������w(z�Z����� ��k��w'��ju���=�A�2��%.NF�p��n��cM;��������@�>�Rϰ��~���Gc�޵������w ���2/���n�d�~�o�)~�'��ߴu�e�r.��ߥ���vo�O��J��6�������ԟ��X=Gѫ�����L�D@0"�@��~c�c쿮>��u���y�{��񯤯��f^��I�15����%<��Zܗ"��5�����9��	oK����4�N�?FI�����y.@v��G��j��� \��S�1�h0H������c���~����욓-IØ_a�%<���%�XP��*r��C�`�'ן����'Q�|�OS�5<�"�g�$�O���]br9�z�>��U\*{޻�YX#�������ĺ�}]G��x��&��r�{��|�'Rl�~hL��2���E�A��}iwUC���n�'g��y'�f�L�|���}�����߰�dx} �G� W�xc5a[뎬/Zu�G�6���[ɏ1M�ݝa'3�ɘ��K9��
׼t��՝$��/0�v��b��kȊk�vAe�����zU��6QNG�֛IgR�Z���T�T��.t�4d�D�����`3o*�j�*�0c�!Y�o�3�kkr?xx{���:������(���cpj���I���}&��\��� ����$��FK�}�'R��R�jO|:�n�˒�oz)�\���߻^Gp���y��w͕e\E��r/� w>�Ǧ�{�@�����X<��s:�����ϵ�������O.�������;� �5'_`~��d?F�(��T:���7�MA�rx8˟\��G�}�{�"tt*���m�g��(��ϼ.<<���>�(����}����|��w�`���|}�A瘯�ߘ���M����<�!z<�"=�����t���b���|�������xoz��26���:�����si�S�2��4naˑ����6&������.C�<��u����$�}�Or{�z�+��W������r�����
��'�R�G� ���sMnOdϱZ�'�Ԝ��Q�u�jrO�Pm���)vyߛz���5	�>�v�&���5�{��p�������w	I��0��^�@���qK=�լ}1aT_�s|b��x�)wjx�I��-�Ӭ(��rA��_cP��bn:��s��`�L����|������߽�p��!(���/.��A�w�4;��j��H�V*�}o#������~��P:�B~�Z}�r�!�ϵ���Z�~g ����{��'�dQ�Y�~�~�'R�r_֡�x��2;�����$ܙu��6����%=^s�{�t`���>�}+�j���z���JTu�5��5�dt��j��7���i7=ϐjz����Rd�k��j�=>�I���2M�?� �\�I��%�r��y�tт���gy��@�@���:dxL�\�惩�O��'�9���rB���i9P������O$��{�=I�����������j7�:���)�9�R�W~s�����:ι��sν����ɧ��N0ѐ�����רJOoI��^Z���0�K�R�����~���.G��u�.Cל�n�_#R��py�^�:ó� Txdx �E���R�}}9U}Ѽ���7��ooow]���^)WB�6M5����wُ�{G4fNc*G;���t7�J���Ǡ�5-��nFsv>X��#���v:��;S��y��>�C�[���w�V����@�Ct�W9Y���V*�T��k��=� �0�����{��p�#�J}�حC�ȡ?��iY%}G[�5��jN����j2#P���ϵ\�#���Ġ�9r;�4��.���u�߱<� ?���|�ޘW}���hsW�'�O=�:��|]EK�P}C��٭{�d����ݒ��7	F�%չy�(?��%���{z���'�Z��T?I�j<����O#߹��D����}sNʘ�����oy��&��5	q�?t�I�S�?��i>��������@QA�h��C!��y�/7�	�t�<�sԟE���A��\�������BQ����}G�� |�i����ٓuQ5y����I��jOc��j��)�NGg9�ÐdP�tg4�Π�>�Rgؚ�&����7�d:�/N��������K�P��Z�_aK�f��G�� ���_gl�7o���R�=���/QN��8~�q^��j^��N��k�����$�Nky��j7	O���4���dR��Ӓ�����5�/��S�_�5��?�Q=1�{����oW�ՔM_����[�0<" ���?���.���W��u&C��;��y�����QG%�����Cp�G��7���`�'��1�����<����\���aGf`���7�]����O�[�o��}� ����ܝ�<���]hJz�`����&ℤ�t��`�@z{��9&���˳�i}����~;�׸
(=��惫���沟e�DxLq��2��|N���fq�|G�O�u�8s
O��s*�|�!5�hr~�'�g�vu�nN��jN���������sgP}E	�����9#�5>�_b���n�X@y	�����~�l�t���=o/�q��PW�`nM��z�kG �KXPo�kr}&@j��n�r)�\���Ey/#Pl���<�/]�pL��?����9�����P�up&G���W8�&���%v�ϼx
���#��GP�0�]����؝�C���X����'��qBPj��vI�5	k7�����L���u����=���(����n�Pds�{��x��~H�� vS�߿x��3*���"��bee�LS!��X�뭻�vݳ�W���J�]�Z%w+b�uszr���ok���c*��l���'L0�pΰ+�K�7>����d�>���Hh�f�(��Yu�Q���
�U�'�����%:*R�~����}���/��/%��n_�ӹԹu/5�|��%	G9��N���'�֓ryPd�N�採)�w�~�I��)�����}��x�|>�#� ϻ��so��pݨ�Ξ�y���{\�h亀��a�|��w!�����=O%湤>�Rd�:��k����K�s�Ӻ�A��}�;���jN����bd�N�S�{�{��#�2�ľ��|g�ܬ�)����5�dP5���r�����x�4��{'P�!����=�P��5�:�#����=��:����NZ�Rd��:��K�N���AU@P>��B���ޫj�~/Xo'o����d=A�bp9�:��:�������N��>C�{��{�.�>�M�Z��d%���u'9���|�^��!O�\�����(JG\惨q����ա�p�7O�>�8/v�a_���X�/{��L���/��y����d�?a[�����FK��ҙ��j�}��ܙ?��r�u���==����9!�1���^��A��ז����T������w��@0<)���z;�$ȡ+��h>����jɜ��x�I��w]�n�d�g��#���6�V�2�ø7<���s�<�'r}��}�<���z`E��r�����;�c���r����UPd�y�I�z��I���4u�	�w<�n��y���\���;��2(sA�}��q�w�(K�.Mi�rM�~����(5=}���|�!@}L}DW����fW���|$ͅnfs~���u�d%��֗۩=� �k�Q��r)����伏��{��9�;9�''�`�'i�~�{�#���_h�����2.�К��'^� L���">�F�q[V���y�|(�O���d?�u�BS�C�����(J;�C��u����;����9�j��O��9�]�QG'��h>�������z����0O٣I������Ƙ��?#��^O\9~���\�co
�јP�S�r�::�7'�N��I�u	N��]����L�C�kr}&G�u���Ho�'$�Q��5I�� �{{������ ">�w�����hfgk�]�76Y�z(�쳒�+����E�<hP޸�8��c���ܕ�k��%9�@]/��mNLu4�R�j�!���H�cɋSy����ȑ#By7���^�wMd�Cz�U�I���������+Se�\�l,O/�{�E3<6u���{���C�R��t���^���񘚓�2u��-��O����
����b��yjM��&��2MOI���;���j����n�ȧ���w/��r&`���߿$����c�?g���}B�������PF\y����X���05��#rx�a[��2Cf�
_-I�.�h��r)�:7��
+�vk�2�pl��:�|�����6�t�_H���o�h6�G*���?`�F��0)��C�g��p��,�sA��2���h;���MFA��r:��u'֬�"��ﰡ��O��;��c��'���;�L	��U�Wt9va\"f+���fpI(��%�
(�=��j����ǒ�׸�a�>�.K��l���\�u���(J���{��7�}��`�&��~��Jul�
�G������o:��,��n9X��&�2>����u	f'$�m�Zy&@j2�w�ǫ��]K��j��˩�އ ��ך=>��NI��kX�`�O$��n��Pf�К��1��`�ۙS�'Z�,Dx-��&�s
7'��5��ܜ�A��x���9��A�%�^�u����5��sp������9�Ȥܙ��惗p����ӿ���ԏ����9�ݿ������#�P���&�\�xs�.�(�A�q�p�;����^�>�2��Rs�G#S��S�-C�����krW�d%���4��rs�����>�y�Sʑ��gy[�.?Q*M���~������R��n�����Q߿h�����K����y��y.@Q�u�%�j����w/-}��5're�|?~�gp��.]�y�ם�BS�k���y���~�1X�;>}]����@�DG� p>OA��$�Oo��S�<�BW����5?�Ƞ�����L����q��PoyE?I��#����亓�x�(?C�P��wpd�]�{�c>�W���z�k��]���c���c�?y�ӑw��?O��h:����uߺ:���yj��}'^`��Χ�ԞO��}�Z
{����.��BR��{rB]�vki�}&��K���n^\���>QP�1����}RFp�v����R�/���8I�X֌�^��j���L�xj��h��b��dHn���Q�јc4�p5{���Y����kP^�����$!���;Xsh�֮7"�P�Wb�d貸�l������[	D/���f��5�����a��~��u�(�ܙ3�6���d����|�R{?�~��q�%ȹ查���|�}�P�h=���0S�h�O�}�����^P<`�3�H�F�cu����O� dP�<�ԕ�2B��F���MG��|��)��=�{�K�K���r�' �7�-��y�=��y'P�$�|�}�<� ;�7��e��"%�M4���vɜ
:�ˋ�[4���z�Gr�k�x}��9&Z�oX^��%>I��ݒ�XP��X���� ٜ��&I���h7>��jC��u��y��dQ{�d��#�����}_������|Amq6͹�~��3ؿ}"�����[a��亟��qA�9n��7�d�M���4&I�j)>�X<�'��.�*�tu��p�9;?o��=�7�eן�ϰ���=�|790*�YY����j3W���|��:�A����E	K���5����%���'SOq����sO#�|�'�`~3�QI�i�z2_-C�=o_aK��=�&�7r_�DDyǽ0 �j�T�_F�-���ߖ���>������b�s���ܝ��`�:�>滄��������FE	A�~�yu%n��c���Ru�j2�P�}�U�eȤ�2@�Ï?W�<�c#� �}�k�}���,K�\�i�2�����y�?K�v}����P�4d>��켵�v����O$˓��4���Jy?��.���)��kp�:��߸P�� ���L��y�gm�q[��" Q�������S�L�ք��L��~�r�.�<�i7�&@{�����9r>�_�y�7C�q޹��}�'��δ��Bd����h�{�ص��ߟu/�!��b�[!�0²o~�����,
�P�9�����L��u�ܙ?�R}<�GoX�$�5~`j(J_:�N��rB}����4�ɨ�>�CF��=��﹤��<.=����1��W��F��w�0{��3�hMw�.�O�욀�e�8�~� -/�5d��BVI�<�/s��nI�sX>w���)�=߽�p������t����A�.+O\�b	�Ŕ�Oօ������Յ
T�ʹYcEgj��)���1�f���y��T��a�ݦ��z�_��| ��6Z;u�� ܉>!+{�cw(�gij�l"�m ����&���%��zK�]K㴸�aa�v�YGz��[��r�~������/f�;��`�I��9���F�9�i�C��r)�9�-�r�\�p��ܝ��u����eј����rvoQG%�j���z�#�z���1�Q�0�1PJa���&�r͘$��N�����]q~�a)����w/��c�JT}��C��29�i���<���}4�ў�H�pDdd|���
ۆ�D�׷KK��y�{a���E�c6��x�l �#^W^����j�3�D��X�+�d)�
�ce$�x�Ujƣ/��@�`���.���Js���9�쫇��5��o�����c%y�Z¶�b^��P�O*u�4"��WJDuyep0�Bg!N\y�بe��.��D�)S���Gb�e�cÅ�J,+��0ut.��!�)v�8완!)�&��Y�5�T<��|���R�ll`�E,^�1���t�~,�;P/4l>�-� �j��p�z[1��1��*]�b��	ۏT>�S~�v�]�4��D�=~����[{�u7]���*�ՉU�D�����͹X�ޚa7y��@T"FL�ce�&�R�x��^{E�omQ02�Bh����tU��y�ߓ*�ʉ����(�	�R
�ˣȋ<b��Z*����������{�!�~?�����ZO]�m�{�r#��aK�d��Fh�^�{�*������&��|�F������-:��n�Aa�c]Ȧ�m�!��𝷒!������9R�o����F�Qk�x�x����Ecq⨞ݷOI��d׼o�_�1��󺞟k���Y�G�M<3��ݞ�@FL5�V�϶�*��:64�^�Ri��R��� �T*/U�s<�mŦ�r��uOg��V�ڗAQ�
 �1�8�ID��Ƣ��}-ˣ�Iَ�<�i�+jh�m�W6}�p2pA��zJ0�I2�P4r�2���V���+���\�Ș`R�}!�7��S�����'�Q�B}#D�o靲j��"v��SOt��7+ѽ>"�j���7/" �)�1�l����~چ�+��<�.2tGw�#�/WR�J��4�`�';�τ�S��ǜ�=���s0E���{6ꊱ.:���~��; ��iH�*7�F��VF҇+G]�}�lH+���o�牛����q���]���}��XŔ`����"�aʍ�r�b��ۿWaBok�;�p�A�mu���#�vAO���a��4�u��x�*�-Z�>�k��D�n��]蕭�Q�6�X�+Ss 7�BW��-�B��d7�kA�6G#�8<x&o�rq�\���@c5ct��ֽ�M��ÎN{�T]�3�ϑ��8\��M�[7jt��ܵ�ͬ��a��9����q�N�Z�)a{�x��y��M4�:�2!O�3�Un^y�(�9��Cά��L�Mvx�`I�W	�:�V0����(�nt���Q��;rUt9���>n�ڌrd�ZY�Z��YkR^Ͳc��g�+��/Wwop204���1���J��M�^��(��7��$���H�U����v�b��i֢A�8X�Ȓ>��!�PP�iP�nT
�5���ؼ(�Vu��B∽<{����xx�~l��8%�ꗞ�蒼z@Q�$'���ks��l�٫�b�Ӣ��Jy?aOG�R�S���>}�f��*
���06z(�p}�\(�&|}�iu�\V��ޠ��~��\}��r�������
���jak�Gb=+ӊh�enԱs�	���\'�kj!�r=A�R�p�s�:p�.U]~�:���q"+�D�'��5`�'�,vg��37�T#d���{M�>Q]k�!��y:qv	B.�$	��0�=Q�a����V2ZS5f_���,4֑�R8�J��ǚ��p�B��	��� I1�'��C&�)�v�".��/D�`�wW[S�\�����JƥL�pRRP�ya3L�tUm��)�8��ef���'��k$��Tc8;���Nr5<׼g �n[���r�ި�P����e�R̡��Kb �ιI���>*�G�8�ٺ5gF^��Rf��2�6���]�:��Jf:��{���t\������1m��ͱ�ve�m�e�5�]�+�2���s$�t�GV�Z�2�Xvdŗ� !v���5�Q����c1)�gu�:�}(����:�ͥm'@�s���&��F�`����B�9�V0V���[U�k[�sV������W��=�:��X���Ш�+��)ڹ+�#�][�evi�<�F�;�t�����]�7k����r���l������M[��6�h6Z��9��R�9o�ͦ���Z��ivX^�8�ĥ�.��*�D���Jܰ��vus���;[�*X%��R�̀��e��*�������p�H�;u#�F��5����L��o)�1l�F������_E�;���,�4�^�b��x�怚���|o.�]���|�is׉f�A�j��Cf�+]k�_L}&+�4�H�Ax��"evq��}W;�ᢓ�/��u��}�M�U�:u��T'9+&er�n�����z�C��GΑy�u��׏g��B����V����̗>w��Z�#>>=�VT��iq�%1ܺf^<g3^Ӿ��>�B�zr���&�#q�׍����g7�2:B����=���N���F$�e�ˍ�لg�,sf��Z)s�@��n!B�b��ɛ���Ճ.�;�r�#ii�ڳBf,��Յ��{�Y(�/[]�vh��
o=G�#�ܮ���5p���fv����&�@et�4{y�Ru5�z���A1푙�:�;WL�cm�@7��)oo>h�:����**Ք(w>]tޙy��ͤM��uh[�{�~��{��#n��[���.�Ǯ��3����aj�IeӼq��p9*���7geд��k��΋��n-+��=������vnj��:��*/t�MT��
\�v�wV�աd����ښ������Е��m�v�=��n ��v�N��(���voi$�Y��vPU4%�֗}����q��19��R��u��*�ԣ�{;��9uҌ�;a�ی8�6��6�+�9��ﶥoF8�Į]�w�_F��r���U�� ����}�� �7fE�O�D��f�Z�ܼkyپ!H�#e
	�+�&�gZV��ރ^���*=�+�F�}y+p'8���N&hSܘ���F��O:��i���\����)�ˊv�n�:�@��O�Z�s8�_N�8W;k��X�ӗ����T5+��v�R���hlTMj�ۖ[;����g�m\��5�F�>� ��(
))h�*��������* *��� )j(�b��&����`�������*���������	��
(�d������(J���))hh��I�Ě$"*"�� ����H���j"�����(�)�(�����"b"����������dj�b)�!&�e�ZZ*��������������(��e����
)��*��"ZI������H�����)�2
�h����i&��"�f�"�hJb���(���(��&��%������(���bh����J����f)�������(������Jh�����b*�������ȪJ*j
��r����)&(�"����"
a��B*i������3f��(�
����k�s��ߝl뽑׮dT^�ճoc�e�<,�f ��'wd��_]q�YvǺjݠ���Iv$��:&j��#{��Ή�Y������-��m�޷�!r�zfd
I
��!Exӭs��͚�>�۰��m�U��튉16K���zq��=!@>�xF�f��Ê��1���Î^
9@f)X�U���V��kq{���w����:!?5Y&^H�];����U����	nh�Ȥ�w7�F��Y�Ѷ�a�a:�ؾ�B�-�W�qnp6�����@�
0e��V��J�R��.��mR��b�t���
�")�=8PS�9UÀ�4Z��o��Z9�)�=7�V�M���r�.���@���~ěY�=AX���Cv�
l�M�@�v��^��BǪ��s��u��d�<�O���L9�(EC���%T��n\{�\�.�[����eiMjc]�
��������H��x�p�Q}H�N˅a��v8��پ�Aq�뻕�})�@������ȧ0�Ȥ'���4OE()�a��yΰ%D�}�����hTy��u;�}j/�ϥV���Z~��l9S��F!�����6��C;�;^�ÃJ��v1���p������ؖ��w��w��{Co\*��M�5����c���� �;�^��u��B�CHa�8�hx
�9u��8���.|wv736'�%`����Lε�D]�t���,��l�ؑ��{k6�������k�Z��moY��v�./��qaqM\���5o+����`܄��"8�'D���_�3�E�w��P�����ڥ�mp=N{�
,�q���^G(�$��z}n�FK�f z 8SŤqH���a�L8��uڀ��Uv��)���R��>��m���(����/y84�@؇*$�Zr@�t,���N��+ހ���2�M�ot�; ���l�K�N�f�e���$k�F�R�
��|�z�Jj�bP̖�ܮ9�=��n�+Tb�c�X�[�c��a2�cChV��������N�9\P���\C�r��Nfn�y�^pn��*.+�mZ���n�)���^s�骵@�`t#9�}����fq�]��V]#b�O�XФ����߽GF��x�m�7Cb���L���N��շ.֕�I���fڴ�j>�VE�e���G�2P���!ܵ"�����̞w���]1�i�[q�H��`j#������ױʎ�WT��j'���G����)w@p9@�G�&m��,�d�}|���T�iE�U��͌nT"jT�|�X�L*���]�Ղ^\v�Ԡ���z��ƹV��A<3�"%r�fb���ͬ�P�<�8��đ@�Wtk7^.����-��<��"՞�˭嗻F���������,���|��N�\'"���T���F�L9ȡ���HM�T4q���i�����<�iW]+P�f�z�iӀ龕(��tL}���F3~�y'�id%ҳE�����P1]�'/ �6�g��ޚi��<=�?��	���)�W]Cv�m�w\��(�B%Bkۜ�m��E=��*��c��vQ�'*)��%oM;��9��퍩���u�P��
�NeO�����qq�"���hw�Ad^��"1�;��竩宙�!\��j���!*��T+�٠[�w�;z�����Z:ʼ��u�:�,�ՙ���n�U�>��VЛ�R�HBP3��P�<y�K\'*ͨ<�uǃ�j1��s�C����X�9<)�W6�s��i:��aȓ�)E#!q���f��!��_iK@����q��Lߵ��sa�C@�=rpA�t(�!>����Rh�ecG3,o='R��>�E�%���?/��8��~���"I���ϲ�&�i��"�=p��u�u+ƥEYi��d�\W'[�p�!��]���t��<Ro:�ǫ+�B�	n�b��h6N�+E.^��B�S��ۣ:���{dj�*]�X҇n⥻`��>��R����Ow�)�t���V[V]�BO;�1G"ePMN��K+~����Zg)5R��2��?�3&��S��U�c%ũ�j�j[��U����&�~�ٿ:�jJ�~*���F���.*��u� gvn�6��t������
�_��ը�S-:E+�|�א~�Kf�+��Xǔ�WK���<||�����־�/Ca�!�唦n�P��˨t���:}4|���7�ႊ��+����.�����7^��n����ɜ5ۻ���|���\\S�*S�R�`bf�k��AصW,��j�D�x^L��җq"�}�f����E�z��aO��]��t��s��T;$u%�H�}�]��F�ח��K�� �WT�s��4�oݦ�/}�5��OU�Bݍ�!���sڹ�[
v��Ҩp���=I��ҡ5�*�Jz�=�㑍P�T�uU���H@&9�]q�^Zz-N	n���W�\^T=`!Q&�^s�"i�ȽZ�R�x1i!ʥ#Pٵ.�;
(s;2���YSkH�*���1�����W4��[�8M���B����c ��v&jp�mԻ<�f���x �훾ݵ6\�f�L	�9����έ��er���_'n��{��;'S�Z:�>�{اk��ٝp���Hέ��(>�o.Cƍ ��l�}Ҕʱ{�m�I<9V���1�/}u<���<=�KO��r��dT/�U8Q�K�;r����6��	�VTƅ���G�/N)�.��Q�,Y�7o���qшa�������V �8xȨPY����D�Ĉy�u�<\��yOOOO.��%��QH��{)�`�D�&?x��=�`y��'N.e�{}�xjލp�ы� ������ZU}��+����"q`�,WeSⲷ_����=�ߠ�6�*��ck���T��+��5�I���p9
(N��z�6k0�O�݅ Ӌ{��A�����}+�k�n��ol1a��*�YBѕ�S�<��|)}�Y�լr�F��gfs�q9'k�;ϐ��P�ߍ��B�YXN�ȿl�N��'&�͢3���Z����yw!x�"ǹ�-v�0(�b�!�̧��B�-�@;������蕾���E<(l4��C�]����'��l���O�I�X*�`�&Dd��xr����^r�do��j�3���\�8NՍ��y^("�P���!�&[�z���i������4)��M�
�U�Z�/�g� �F�T�L�	1����/��:��z���K>�*|42G&�����d�\T޸W>6����ICCy١VqL�iI�"�,��8k�B3����W)�����	*��U}�{�����F�ԙ:�э��=3->@������꯭䭜��u���;ga4z��z&��Tb��S����T�=W#���oDhݭ�����UpL��"�NÅ`�Q�`
P�[��J(^� ���mJ�"�{��Ww9������<B�q����k��L�Rķ[��:c˘:�Fƙ|�>ze�o�n{��_wY ly��WQo�}j.���S��S���{��X1^L��y�0�F�N����E���)@bf�'uB��R����Qk�jjts�^y]i�`x�VH�̺������?!�gn�yW��	}���/�] �׼qP��B���js�
,ˎ��;�B���2U�q�q���k�𚁍 �e6+��Q�"���{k뱫nE�q��L�8{bD�^K&�<�����>(�O���/y0����x����Ú�A��ͼWW��)�� �ZB��fj_`n�f�,F��#I�Q�¸0�X����IP�zu�WY�W6�7�����1c�X�[�c��a2�F{�O��S��Ec4��9=��N���5�[Z�K��A�웲60R��;�`YX���;��7Z~MV�5]N���*�[}�U��*������i��;�.�Bo��Ch�]�u+.��FcyӜ5�-yȳ�6ku4�v�IN�1%�R�.�����w3��,��}��U��Ԟ֧ZP8�
3��^�"�V@�G���G��U��2޹���[d��d��݂�b��6-2�b|H��
��
�U��M�힀Ú�~3 �Ɯ�yR�72%�V==��:�U��i`��m�4U�O�ॖ��}�4�6���i�P�G;��cZ>K�O(��L_��lX��::3Yd՜�>�ق����q��@٧�7S�1N/��qV���hD!R�&��ש�p����ccT��mz'�&�W
.(�%�ʥ:�j(���'�l�h�[��og@x�Q�s����D��ޱB݄�ǨC�8���Z���CO���GU^k-Z���'����(��������8۔�D/:H�w�,C��
�W4�4=D�7r�N����s(RR���.⁐�J���<�[dtW
U��i��[*&:kgTn�r�x!��(�bUQ~�*.���dwx�%~��T�,m����EC�=��m.��	Ƽqܴ�M����7~��L�4�F&_��St.�J�+!Y��ޅ=�fɨ��T�WZ�o��:�	��I�k�]$�j}���� �e��5nk��-΂�\�z:� o\�{�Q��mm�S�f��^-�S�v���:�&�)��X��<�Q	�v�qMG��g�ZV����k������K����\�K���x6w�z�s���j~��f��Cu[��r�l/�S�h��ﮏ	~��❘�ݘ�u�G��;�GO*�y�E��x�ˇ9�N4�H(Ñ$p�Q��Բ�f4��x�S��9�m81٪�ŗ��S��(���5b�B��ӗ�cbJ�vra$�B�2
�V+hD���"���5}�<�DD&�u1M�d7�n%Uu�2pU,�f�7�\n�
�+H%yH�Z�*�VFC�R/$�bX���W��A��p[�-$NkE/V������r-���G���ɑ�g�"<�O|���q|�ٍi�w+"D&�y��t�C���ϯ����>�\.���6m�B½�{}��B��%�����{�~�3�kަ!��N�N�y2�2w���A�g"Os�	*x:�.'���=B�R햱ɸ{���ڞ�^��珯��O�NE	yװ�٭����=Q+q�����} W>a\W�!Fu��ӵ����>n�ڌs��8�ΜR�������)814����n&br;Yv�F���yWj,�3#��2S2�+�Nmt�����i��4�JΜeښ�Wil�Sy���+Z7|gj����+�F�}�՝�/�O�wܧh�CS�5�i��m9ѝ��]J�TP�};�*�{�ʅ�.�[%�9	���F1kq��=W5�Ҧ}�2�)�u��!�ϮJ�ܚL��F�(�`��]���wt޵��ߙ�Oj��{=��^	i\��������z.�ڋ7�#KŹ�J���ro;�8�J�6��vR2+�OE��%�ꗂ'�W|�q5\6�/�p9�\�sd�}~���No*�C�|\ٽ�x݅9��Qaꬩ������P|��E.�+E-�=��Ve���_]>�k�*�K�
�MM@L�r���}w�0��!I?o,k�N'3���Z���O]&����Ң��V���w�p���_�ӭS�:�(���IW��T�������	:�e�-P�e�mȳ�f���-k�ͫl�4#A^��W����n�����i��W�2�)
V֊������=�S����/��	��Xyf�
��n�:!�d�#b:cT$��0k>�����B�,�9�C0�`��,)8 XF����Eɼ֔E�p�;�s=�Ð�h�tF�f���qP�pLd����0�C�Z��'��4�[�_A*Z ,4[���`�
6���Av1�ZΦ�[��.�����=������E0FV�#���Փ��'1c�#��ud��V6=&�[����i��.��7}��5o�Lx���.�c��=)�n���I-7�������^�V��q� �Xذ7m_���b���b����-6+*���k�U/�Xs\~aF*n��u���,�QJ�U�ՙ]�h[��� ���-�6���:ݝ�[&5NW���".�on��F̰���O��������8PS��Up�[�^vZ��Q�q��Y�ﱉǻT�.���SJs�=2hO���
=�-�z�PW�i����7�Al�m.���ٞ��A�'�BJ��E�dv��$�T�z$�clU�8�"/��v���cL���.�G=��Sq�ұ)?7a°](�9,����]Bv60�p��@�x[O�e�ҽ�{�{�/�/���9x W=�2;��no��lS�>��B\���W��c�(��q�1��{��#c�m����v��[��U?�7/�Nǹ�P1�2�iѸ���=��vm:���R|��x2�^�R��丳��M\���5a�tr}�����(�t-㯙.�t�k��������L�2�T.�ˠ���z��B�0 ���&ӗG+���&�BU��P1�3D�-��v�f�acw0��!32�>�G��Q����������k>B�1)w�;�ax&4�
��6j�pVmc�4��o�w�]�R�c�j4�MХ��@���}�P��Ɏ��/��v�����3����w��[�Y��*�W)ݰ���9�u.��[�NN�6e���A���4 +�ݛe�Ř��A���t�N+��Y��R��sP��gtU�Ȟ9e;�-%�F�P�d���f�!w�$I����]d��� v�ƪ�@s{�c֖i�7��Op�#!K��^�]u٤-
̾�����e��M��R����������5����>�t"���d��t�[���,>U�v��Rl�h�cO>%K�����ד��3�ĥ��>AP5`n��{�X���e�0 :#�<����+xu��T�]`VM)�lp����\i���{Y۬�4���T����vY7��Ǚ������m�:����lr,-'D�W��5n}5|2\�ɀ:��E\u�H�\[D@ȑ�feR3M������{���jua��oGuX�m�BH��4q\��799(�6�Ma���J�VN��ǆ��B����*;Y��Î�U܃uǞ�+�Q�Z:����ۖ������b�=��֟U�,A��*��5ܮI�!����%�dk��[� �$t��W/�n�[܌�)24��б��H�+G+2�gn�+������#�gr�9�u/q_h��e��ǝp����8�������wg�NwɅ� �E���V,��`�����Z��QXy���~�վ���+�����&��ȉH�+zR<6P����q�J�;&0�s�OI⴫��*��:%�z���/#�N�;�J[+r�'"�2FŅ���L�髮JTbB�*��P̙�K�Y�|6�]BrQ��^:���ŗN�F�S���Y��:��u�Os�ӎ����
w:����o�о�QÆ˔��ܩ�j��zd|�b��k.\�r����=���th�5�!5*�w� �y�o��.Zm�uc:NIV�z��{0���#���WVMM��v��̾j�Q�����F�HC�J3y�c�k�g2�ȳ\ŭP�Ԕ[1q=R�����wU�ci��ui�9�k��u
�j+\���Ch)���d���
����&Z3���<��v�r��4+�X�GoXz���g�X��f����c �6�Ba�\���CW�3#���Hn�0F�PX�tUt�if���
�)� �Z�ڴ��ٓ/r�z
�9t�C���ZN��Ξ��� �N�����f��.�S���d<�nd�s�r�"iI�Ƴ����y�6�lJu�(�\h��8ན�����R����w�o͏k�`g�%uEw��f��!�6�Ҡ䮙M)�vG�Y��L�1�p�B�u��&]\��=ӑ�z���~���+L�R��PQMǸdMTPST-3MI�L�USADAUITP�ITRAUDD1UQIKT�DKUT�DUMQ�.XMQ4�SQ%SULM5TEL���@Q4DM��TIT�DPLQIPEfSTEQ9%PUERQM�QE4R�$4SAC�UDC@TddCD�DL�Q5EEQME%KT51D�IUU4CDQ5T�Q�aS�dQKT��QDA0IU4�AKTUNe��If9LEU0D�4IET$�IHCSMQE4@Q@QCPTRLABENBd�Q��HQ31UTM%TETMECLDI2PQMQM,MU$L�MR@e�\�ͥ�ᕷ��w��9��h��`��͇���.q�'�t�壯��[+��*fۈ�#�r,�K��܏�x J��A��!B�:��4�hVx�@0Y^VUR*%����cV�r�ʺ��UGDM�O����b�~���ߪ�.�q~�pL��j	�?V�����t��>�Q��mw+�-�Zo�_ U�}�q�pt^�5/��ZV$����U�.���f���[/�D%��͌5]�IXG)N�ïf�A�3��J�ȱ��1A:q1A�+L�L��_~����`��=NX[�EB���A�b�lo�
Nv'����x�Q��`
M����ȼ:�dIn�*��9T��vMSй��`�4�
VFC��v���T؞��Ú�5
��')���-��p��H}��4;A��U��i`�(m����	z �9K)�ಘ27)���O_n�V���`�LOt�w�k6�668k#�����#�q�4�#[X�|(Z��^2��#�l����	�!)�i4��u�r�9�y�615J)`��I0�"��E���1uج�j�����F�V�K�"}�B|��3AB�z��;q�q�0���]�U]�1KE띲�㪒P콕�a���2����i�˯/D|;�`�-�D_|ܹ����`��f��O5s%Ռ��BmVe�d�N ��7���X6��ߑ�����u׸5�KU�!.�#.�DNwRT�jSn�0v��7 ��=:���幋� x�Z�]���~�%�S=l������6�c""��֬w�������##{�)�o�d���W�m�`ÀR��-Ξ���6)R�>�	��@�mH�;��j�'�v�oZ�ؘ���l6\]H�c�`�!"As���>���9��PX޽��k�u
��ztc��o��[���Su�)����%%A�68�aʅb�l�dU���O��ŵ-��-oo�L�^��}�=l�l;��a�nϬ'U�&B�˺�~\\Mӕ�0g��~�#}ov2yNE9�)ȿ.W�rS��m�eÜ�h'^�Q�"W�\	�N�E���v4E�\������t�B����f)�rC�nrpAs;S�G���ԩ�.t;�)A���/R���n2*���SY�O%�" �4���e�����]s|����T{�ÓY5h��]mySu԰R�T>�B
o�g�q�zjr��L,
㹭���x�Ee�3���<ϰΎf��%�p�s����n�y�����$�v{-17$��Gp��ɹ��C"�+	������n��X��:-!9����]����Է�v����
�E lRGIP�aS��*�K�y��[��ѳg!M��؊ͨU�m\('z)B�4N�7�y���2�Z��$7dm��͆0�WH��E����|aU�mDV����:B벼�y�[6!�v���<�`����*2Z>>G�љ �-��q;���dLk	и�ݮ�f�b��"�t����^���z�D�q�>���8se,����Q�.���S��jd���i�^}J-�T�"udL�Mp�&��c���[Яx�U��Ң��s^2$`����Q�z��y|���\a�y�~N�M�#�3�����6P��m�N̑`a�8��`�|�vU6;M�^�F�(5���N������7����
Y[-:4�~�ؓ���!:�(�ZT&�ە���̀�]���)����Mܰ��"��
�R2(==�%�ꗂ'�H^=
� (����c=���Ŕ�O575���Ԍ�ʁ`;7��������ʋ��YS`-"�����06zl����)��K�\g_>	@�>�;Ce�C�K�5)�.F)m���>�ژ���#dL��ꕎ�W�U�5���ޚc�v�Y.={/�E�p<�&\;DTtu�0z���_�3ԑr^;���{���.T��'��S�^�B�P;�-ԂO�]��s�������H�uӍ=��'p��K�c���Ȉ��XW�+O`G�h�o]Z�N�WN.8����Rw{k�l�^�hu���s%��)c�n~��ܽK����[5x�:���+H$�ǟ]�y2�o��X��+�u�;�l�9��u�o�r���L�6{��:�V8&U}��WJ��<)�l�����$k�<خ�K�E6�q�vz����֙��l���fd
���[K�{J���x�0��(���^O�skr���}�
^�+�Ào��9��=�Ųs�,�f��Ê�tK�GLd��a{�����u�g1.w�x�u�9�c��{����ͤ!ߚ��/����];xb�m ��W{�i�Y�{�NV>�����ddW]VB��q�}���\��4��_{ݲ����`u����]ׅ��!BL�P���dzzo��Y�U�)�z.p�����,��j*�z��3l�GU���|�B�u�iN��4'��B�nn�PW��N�d1�I7�n�'�������R/˕d�qr�흌IR�X4�M#p|D�B(C���k�K����g{��f�]\j��fԨ�D�K�X�n�݇
�t�\�6��:(���!�x��D��͂B�1
����Z^��_#mŽ���T֧��q�j�;F�HF������j�80�GFn���O*�J_pCң�X3h�Q<�,?q����R�����byvS/�tɽ�&q�|-����+Q�pe%�a�'A�y�;y"r{`ܪ9���<����kg���6n&��+ݖ���3�^@����G&E9�-��< �c�Śy<��pO;0�.4M�����*�!G���u����^[��U`�ͩ��Sް`���3wSw7=�Y�Vlf����H�@[�n�:>| ����W��|4o���z4��{{�N�J/9�$�S��"��x��k)���
Աм��|�WCS E��{}��Nn�|K��
�w,e�9�X�,U�:
�Pk���,lVO��;ة���J���v���/Y��ap./�;�P�X�,����ѣ�#�j12����R����g��t��/����ǴwA��3R� n��"�`r0D���)EBn0p�[���/x�u���p#��C����W7:ݎHӐ�30����h3��٨2���f�aa$��z:�e*��U�l	���n�.+FuZ�9 r���m��:�o�����݂{�y�-�*g4O�s1�
�����W����#������{�*ɡ�$~�z�Z93`�]�b]�A�)֝�Q�z���\����R�SB�;��˼�M+a�33�4���q�<k�����x�J����b*��Xm��cޟ^p V^et#�����[D�_ �<�l��wu�������a����dc}�u��yWaS��,9�%_h�6Ɗ�(%�>������.�봎=\Q�3RQ�.2�rԊw�k6->��уYdг�'��ق�æ����T�T�]r��{���1�k�s�0�%64�r�>-x	ȩy�X;ܴ=�����C����s��{t���C��X&�e@��GNӷ@�˽b���v��mL)�j!'����%�yZ�/z110�G�D���2�tLW�;NX�)Ȉ*_�֬qvv�9\�3��S��Ȁ��C�Pԫ��`0� 4�aX�2Ͼyn�9�����l�1�A�{����`���������(�	�R/�6'�;2�$H.x��;}|��u{�k1�*��</Z�et�������@'[2�2:�Ťh�Є�" ��	�*��s֗�j-���u��3a��f�p���_J�T6����>�'U�&��������1F�����\gtv�kڦ�Q��\o��|:�G��DJ�	}��: �}#A�b+&���O@�6�Mm$�-K��̫�|��%w�Q�m�Jk��j�#�?��sS�x�R�{k7����c��������b���Qk�{���C�c��$hW�,/�Q�ÈqDJ��*��'~�e^�J��b���{����/�q���F��IM����I��MF�H��:q@�ā���pb�5ی�!S65��s~l�-
�x���!�Å���}�"H�VA2�/��X�5iY��"���ߚ�`DD&n�%=�y�=J��[e�V�1��!_���MX��׸2*�; ̛��*rj�,d��"s{=��f�O��٪�B[[A���b��s�{L��(��>h�e�!�嘥��'�T��ĵ���U@/׷mOG@B��+'a�v���\}%FX�\q�@�X�a{�N�ߏ2�N�hw�f��vR�oS�aP)�;Q�ʬ�+f�|qX1R�QF�I�O�'޴����t�8]�`��H�Ӆ:|�oU[��}J-�xT�"�/:��)���y]�v8<���ѹ��(�r+�ӚA������Q��N>mk��;Y��j3xE�an"�ӂ���
�d�n�ps$@�"[��!6ϝvU6;M�[REQ�r�14�7֍���i��R����`(q�tN���}�`�Ԙ6�yG�����#`B��`�ӏ@�i���V=��R@�_��MX��ξ
V�o��V�6���¸-f2�M�G�+V����h�w��V-�K���a��`R���Y|�%;�b뤶����`.��m�5M����λ�a��L��@}ÓQ��݊��_W%���5��&�|3]*�5r/�*����sk������0�*���ت����LT��6�
�ܛ|;�4ʃ��40�ʀ�ke�y�
9�̨窲���PT�R�b�>�ݙ	��==^�V
�cʗ��}�kF��,��q��^5ػ��u�З��l�v�X�W|�X��ܞ1:U��������4k����\'��N�<gD\(�J�N]���;8�u�u�[�"�dI�8��D�m�79��+�.���8�����I��	��T���ή��φ���;�I��mU���"�Nte=|��M��jX� ��L���SF�{+�_p�o��Ί�{�Z��QSr���j'�.�m�o6[g�n�Ào���s�9���f���6<��|*Kۧ�^*�/9�pk}�G��Y<f�.��Cݷ~7�HCh�0�Y5�/N
����|3f�/�Q�o�D���� N$Fx.���f\:|;|ǜ-�@:�qnq�]ni�S
ޥ �����tG[0Q��A��3�L�jp�[EJ�J���\�,�w/Ga�U�۽���.m�^75r��3��K��;=E>����s���FE���Mچ���}KC�E���vq:����dԥ�<n�䗂<]�W˩�p÷v}�SJ��J��Ul���k�u��?z��F�W���=3�bHfp]q4$�'���9�C�b�S�=3B=v�6q
�i�QݧU�q��[0�V�Fai���nhW3�����8�dv���*��z$�C�mx�s��Bf��r-دK��V�z:5��ҩ��n\�t*��P�~nǇO���5a^s�U:X0S��X'v����s�hB�i��OD֕P�n�ۖ����~N����E<��˨-`����;9�7�ǈtXfx9�&B�m��c�L�ҩ����u���9�7y����� a�s]�����D1	`��%ҋ��h�>�U�.���{�m�o�[���t9�e�}���\ox��t0����4f��f�*ce�Q��d]�TlA�[oG*�y��!ś�C�e�v��ME�� %D�B�ce��T��D��w��ogl7�^{X�T��\bt��\_bw�
���K8&k��V�d-F&D�Gp�(V��-�o�q�˞�#V���QC	�J��	X�2��af�/2D��^B�zC��ߦ�A����ڷ�if/�NSU�]��}u��2lp`&�f��G�
����`�O�m7jۗG1�Z��la���=�u>��9�U�Lv��z��b�P4��#�;���Ƴ5/���!��d�'Y�u!�x���ew1!Tp:2���Y���b�+3�`��UnE�fa�	Ӊ��Zf�*5;:1���3���4���EW��n꽑v��츫�hKl���W<y��ypZ��W�t�.����*d�e�sFr+d8>�U��M���j��c��d���-����}��mK~�V��f�ZZ"�h�"�^�3�YjV��4^Vv=[��Jv���,C�����"�j�4'�::0k#�����#�q��)�xkݴ�_Y��ES{)eZ]"b�_��q�����i��'^�~.�B^u����[^�����0���ޕ�Q3��B��:i	�QP+ð�
,NӷbAr�k-�N�z��SYpD��0�{pu_������R�}�	�/���.��b��6;%�=�8��qs@�b��_�-�RB�o%;\�t�u���A�|Pԫ������!�n±��6�5�/E}�sJ�|��t|�J�s96�ew_ٚ�!��O��'��9a@c���E�r�[zF�lo\D��Ð�k^�ʳs1�שb&��,�¹�gc�۸��:�]ǧ^*;�n�IM|RN�Z�<��*n�A
�6�ԩC��O�+�R�tn��LNk�E�r���6��u5����5@�"��h�ٙ�M��F�'}�qִ���;�6K������� �P`N�Rn�Ǟ��,�Z�\�C+�����l�����+%2���8�X��6������Uxw����l�y��&�;@7�حVSHe:|�����H�@b�!�{s&a�PG4��m�:���V8Wo
@�IS��k�����������ʅA61�k�*�O�C%gsDU�G���A�ֵ���Dņ��
��^��9�E�ǗK&�iڑ��J段F�Jk�M�:ޱc���J�sa���EFJyM�Ḱ_&�7�h����R�<�\]�<Н��0d���o�*콹I��Kw�Y�0u��omF�A�g���^�N�"�5v�;���SC��s��f��Y'u�Vx�3=�[����Y���m�)�1�۠�ͺ�X�8��q/�,e�5�vi̪��v���Vj���Ἕ�)mZ��i�s��
ugX�5�%�Ep��J�\��0�x�ܔ�+k*d�,7`ak:�c�tC4���s���B�S�G8GY2��&��" �Cv�ݮ��r8�Ύ�D�uw��{��nmmoH��x��][ϫ�fwэ�C��P[�=]��5nѮ�۬yeT��H��j^��K� �����N[3�r����e-�׽CR��R��2��[(��2�wV���PT��3W�1¥�J�N}F��N��cu�ݕb}�����X��ޕ��1��^�f�th��'Gjn�靘UD;��*�����KeҨOk.>�0u��B�?�;�o����w���K�� ��)u�(��Y
-a��u%@X\6�FHru��]%{ws%"��{1��w]�O;u���U�(�{ٮ�R�*�^�7H��uɰ�k�o�n�6�ͣ�*8k\1s���z����*Q�|r�NSU7V�$�1ei}�<� u��*-A�`�`<0\���ﲧΩ�t&��]m[+�%�9T��X��+,�$��X���Ҽ3�3��Ծ�+{��4�b}O���(V��V�#MI��E>Ŏ�1�r������݀���]԰v�hn��i���wS|мͷt��4vT1�bh9X����i���tT;8�3��c�ƺs<����N�'S���P}������8j�`֧N��];ϔ��$�uܷY��2�u$0�ծk�)�Ĺq�Zh��	Їgq�Ϻ����]Q����=��tp`")F������]NY1m���J�Q�=Sg.�j���-8OoH�j;�Q54�u|U��zګ4����]_��"�$���w�ͪE�N�W��&wmR���h(* ��&�����(�����"*��"��Ƃ������J���(���
��K0Ƙ�I�
��&���*���b)(�!��(��*��+#"������
J��"&*�*�	��f*b�(��"��20"�
�b
�������������(����"����h��"i�����**b*h*��$�"	����j($�32��������h����"

�&����i��*(��"*���*"*����*���j�f����h��)�������a��j�j ��h��f��������)�������+3
j������"���b����(��"�Z�(��h�"*���"��&b��|( �
B���@��g6�K��t�mu9�YS����{�H��#k�Mt��gF|,�S�3�|�G���ܒ�t��T���9K�|v}�:��%2�\����4��-<��)�~/���T�����/���w����Ob�[g�l�|~���eB2�ҫ"l!*�68��r�&Bø��t�lޗ�g��0v��A�z>κ8�[��	�e	�.��
���<�V�v�y\���u��C�{�Y�ٿ^�QtA��1��t,?/K��1,��cݽ��j(r�^�KyG��Ȗ������������:�?)Y�E�"�OuţE*�k�ޒ�:��g����X�V������j ���[�]�5�]��]/_���F3�c��m|�D�,z�T������M^�U�����U�}k�y��*��b�'��*�rM��.�~�G1<����`��[����f�3ftC���u�`l��w�gͿb��9�S>�6x(�U�v8t�!�ey�n�͈q]���<�`��葀��1Fp�t\�������}J.����[�}C�n�_�zYP)�J=�:W�;/��Ѵ&��:í�6 �8Fi��B:�7�̞J���g�}�����R����R]�І�ol��{�E)V`'�QV��e�/s�Mt�/6���
][*�nƛH��kz36WBE����L��ecHu�p<�AyJoj�F#�\}�{,��An���%�c'�	=4r��ni�B�>Q��9i�(�8=R��1�I1�P*X������5��	���$3�\�t�=j����~g�D��p"�Y���M����kf��F��>��~>	g-k N����/��AH��`��|�vU)+ч��r�B�h�/�`C7��Ξ�P�K��H�ҍ��I��>��8��#Y�;Jj��r�x�S�U	b_K�C�Ҟ����C�t���t��6���R_Z�
�ˏm���3=bb �����sꮹt�؎���v����T�{.�
+��̨����֑PTH�U>���k(��&DF�6(&DK�򅛱���8��@Jj�F���@ZC�|�2����Szcw$��j��t��G�zqL�k+h�	�aQ��}*-p<�`N�<f�hӭZ�
���I	�	�W�iֈ5j�H����+H���~`�_&Q�7�r"t�iP��7���\w�O�~�q�K��0l͊�G��\+F��X�mh���[Yki�<e
v�ߑu���Ђ6�Բ������|"6����ʹ6�ahh�^�$'x���X4�������U�D7���/��k��1v�dcC��|#�ܾY[\~�ٻz�w'W8�tS�<9<�'D�XorѺۭ��/��.@�N�V�B�M�S�s�� ���f�)���ʢB)�g��m.h��g�R}2)t=ט���Ү]N9���"��p����d8�Έ�7�f���C������B������48W��l5j��0f�cb����(C^j�L���ٮ��%��_]�\��+ma��^��7B�8�8%��#"���!�e8ؾ�B�-� ���-�nL���:��(+��u�1���9���4�[^Un�ˊ�k�u���M��()�"e�t�]E�����޾wj��5�^v[��o��Z9�)�86zd��>�B��7����|�Q�{�kW֒�������B�)�p�T�x�ٱ����à��W���:ċض%[���`�!��Wa�S~\mˁ�%�Z�v݇
˥��6ڮ�s;��̯-��-����l?`�w� +��j��;�g���E� +`{�,z/$3V��×U~��[+��_G����g�1�k���͍��~�%�;�Ug���U�E<fP&7���:�7��/T���r�t"9m9���`yz�wD3�z6�h;�d�I	F�8xv�?:���
x;S�y9��Xz��K��oÇ���4T�ۧ��м��[��tM΢�6��Gmu+�0g9�)��}�JT#�.m�P�I�����X1^l�sLK����"���VԺQq|OB�����7�ѻ�mF���=vc���ӑ�nXQ�nC
�"��/N��0�Ex�;5㊅��VEɡк��t���T���s���!E�t:��93Z&��c�
�O�9
�1����n��8^Z������L��9tܮ�)a��^n���χJ>�]��	�|�X�۔��N^��`�k�c�Q��|�:�=c�:/Y�����券����eV*{$tA��4��o0Apٲ0�B�x�+9�%�F�gc�x�[��f�'N&=�+S];����['�Y�7�W�|d��r*�F�o�
Nv'����O��������Z��%���/��s��/v��#�<���u	_e����lS�Ǆ���y�)��!���x��w�7Y��E�8���5ٕp�#c���M�u�5|nd������3nB�F�9M̤U#O�m,G�a\�0'
���8jA}Mf�����sʵ�+h�f�Z���6X"� *S�gʟ��-����3-�r�\��}O�5�i�
�'7ċX�np9�B��+ٍ\�k30fG}'
�J���L}����H:N�jDK��<e7|����������,Ee��,�ox�HR�;6'��M���N%Y�e��g!׍�Q�HB��i���S�	ȇ{C!&�E-��P�Q���*�n�ڥQ�H�˄�æ��R�oa
F�N�.S�([��Ǹ������k���jb��5���PZ���(i�%�=tB�D�v:(v��8۔��	��n�ו�Q�ڈ��Վ�{�� �5.����*�{���<���㖥ٵ�|uh�%4a!QG�Kl
�*&9�룡2����������rT�\�rޞ�������W��Su�vյ9����\z�=>���{|�aA���x*X4�i�Cձ{I��b�]�ң�Қ��B�P�l��l�m��;���Ӫ�Fq�I�T^��6����7�߸U�_��
�s�f:n�.yȵê�X�[�]t�롞{s²�jl�iLVy��t�O�_�WQ�p˅R^|�r+iA��f�q�B����9z�냲��d�����M��Doqç��:X�V_�q��8����8���a����i��x^�� �*W�+i�#=��Yz��A1>�:,���n�[�6�wp�\�{hp��ԩ��k^�n�V�&�X��ӹo J0`�Gn� (5˻���M��3R��Z�6A��d[�tlFN�Xkͭ���+˨wܒ$�2�wuɑ�ǻ)H��'�3��aɬ��iqFk�A��7-�
������}<e���ǖ���<��r,f����=��73��`U�i�͙�⫁�3��
)7�'��,\%н�.��'�%�+�����(7Kd8=��|1�zk���$ʨ�(�b�7�R���f2\W���pT�U[�e{������; S.�{|�+ݛر�Ti&�<��d*T�K�z(�R�Xm��6�������|%}�_h�����X4��cr܂��#Z�W�/��|t傐����ʆZw���^7�	w�7�L�x��'����p������8�L�#+�B���!�>w�I�����X�{�r�u8��)�7�'�^��@�],@�FD��}�B��>�F1���۰���^��MP�j\
���Ω�!��ç�����-��y�>�t2���g+�^��լ�o�t���4��TN�Ss�z�{.۠�s;2����l�m���ʮ�ĄG�ѡ�N�K7�y��B`��M�aً��;�$�{摹��`+:�kei�����ι���wea�,l���_b;�GV{N��՞e�'j��OA��R��i�"��<+;�6����R����f��3���{*F�k�ΧIN�0�B+� ��@�
���,�����F��s�!)��L�r��j���UK{{�u����VT�D�1���4f5�~�$V�}*;ˁ�+i	�{�&���I�ӽ��tR��*���u�Z ׭S�@ Ȓ; ���+���e\k6�ju�a�����M_2�v�=�w���u=<UQ
��E�*�T��+kH��3�0]�{{����t�ڌ����^JN��q�pC�a�sS�Ce�`�@���O��s�D;���5��$�^��X�Nl�O��Pp��Ð�;gDa��oh�R��Rn�Z����'��2z(��(��ݪ��w�P���d1j\�;�&����X�z�ծ^!�Ws�\��`��`dM��fS�����Z9P�ᕊ�i�ɣ�#�F3"�^��o��a��SJR'kƦ|~\U+^���E6@!sS"�B�!��PWDf�Q��^��p-�9n�ޮ�\�Ҝ�����?bR*����8��T��I����r�-y��r��9�V.��#:��#��!�9�h!rF�I	��8��'l������*�F��Rs�:��U�8��~�����He�H���;7�	}��i�c�o+ܕ�	�;�t�K�+#-ӷA���b�C�O��b���]Ð�7~١M�M�@�T��,������R�=C���FT�ni�pR���2�kyЧ�	��(GGB��iԮ�r� :Ar�k-�v)eF9�# �9��[pC��6����KG_*�^�)ODޗ
P�n�9�r�Tz�����Q1��W�,f�ؔar�UlWe�:�Q��W��&�}�|���~���Y����������ڢ,���rޠcS.�.���b$�.�\_�����U��S#pi�W	b�p�i��s��q_�/�y���-�3@�Y��Z��H��!j�˶Ӭ>��\S�w��Qx�ce�qk��js��Qe���:���	���@(J�(�as���Քa��R񫍔��Û��{V�4�+W|�T>�/���P�����.Fq\�W_f���	���a�)�i�C�1�o�K:�=~��q�d���Al�zu^�u5�{p%�H�T�L�uz/M�������+9�%�E(x���><����{����D{\��Py��86$�!�^��]��F���:w�+����n�`��K��+sV�U�b�|8�^I�u���� ղ����F�bN�շ4���*��X�MJR�Uq�_S�}�c�KH����s���θ��p�k1.��m����Q�d���j�_%�f!T8��FCd�# �U�q�ˊ��;2��U���r��BW#�M������[�L����K�.��O��D;�B��n�R͂m�o^��|�����SB{D��fU���tP�B�7�u�6�:�SڧY�M�Og<����BI���ƃ(���.'}B<�
e�����GF{Yd׬�H�y=	�,�H�ٹ��H3��S"�tґ`�T�q���i4��u�w��9%�]`�F�ڻ�3�lu|=I6+�(������e@��B�'iۇ�D����([ȫ�,�z��7�6�_.�̕�)��3��+���w���AHxQU�1��1�����pz�94�huFR�+Vj�f�jWH�*_���֛��{P`�K8mq�LlR݄���p�O_��E9=8�Vߟ��^�gނR`�VQ1���(�L���b���c�ġ	K���5]D��V��P�Gd�Ϡ��mJ�"�}]����'[2�26'rj�P��˙:i��&Mzl�"�Ե9���)�BO�F�J�G�}Vz����_�m���F�_���4���ue݂٥=�j.��wپ~�O}a��;3}i����e޾Gq�
�+kz+9;�������VH�tޣ�<�37,:�3�4�J��r�v��by:�����BC6;�<-yл*�\o���*U����N�-�2iv)w|߼�k��t�V=�*���I��Qv&\�k�U��G���v��{d�\!���r��I��>{	��: �N� �r'���@rm(1]���B2s���l���;W���S�ɂ�ԍ�%�Y=���A3�B}'ٚr�n2s�eS���wN���`�=W6[��|�����'e�^�W�R�H��o/G?:iޥ,Լ����I�2z-�͓�^� �R$jg�H�t����ҽJ�(l������Ҭg���1`Ω��7�W=+2�9����C����l�8��Qc�����߂�桊�-ҧT����Vu�Ӷ�
���u��Bv�b�@)ӵ5���Q�՝}�Yrg�Y�M'��P��+��Z�>��>������u�O��zQ�9o�f���au�j]�Zy��W����!
��୫�<-_��O̯���T�j���^p|ۢ"/!�8l�X�df�[Ua\���*\>0��.����hf��68+{�7���zQ���I��$�b��ӳ%[X�ۦ���{�7��
T��0T�5ƕ,\��쳯9@�޽��9��؊�ق�/�V�Q�S픝]��M�󠗘�(1�f�Ʃ�p+�\7W�7��#�s�31�ƌr�g���L�m۳��<s��3��dCzGoc/���:E�
�S�X�*������˭�$�w��X�������'��Xr�񵻂�*��a,��C��ٟ�v���8f��%�f�֗bɲN4K�W6Q..S���#�rơ��V�l�4��;_CM�n͔:�PO�^��wsS��λ޺����]Zq� �vp�sЮ|%o����k����}r�^�B�u6��ۇf7�/�]MJ���A>&��s,�����Q�g̀#e%�]����I'cl��j�C���ִ�!yc�>p��j�R���G:�-���e�}�}hVkT��75#YW��(�Rnk4w(e ��/xթ2#��ޤ�ʗL�ɣf�����`ٚ��/bѢ� I���
��Wm<�`�N�;7Z��%�כ�qD���G�4��w�����qğ8�3�nj������^Y�X5�:��_�3����h+.d޴���g���y���B�0��U�OkNZ���n ƋXGm����te�{Y���;u��wR�cw��_7�kvr�9�o�&����Gi��ʵj� �U'�s���K��5w�9�5��:.��f��NȖc���P�e���%r[;r+�HY�1�K3y��?vC���ᯰ�u0Ԡ��հ��(���jm`�;����swݛ�\�z�\9gWLFj���J��`�(#�V�q�V�N�T�KS����$�_]�r9dW}��QֵcF�YW]�rV\�����tw�Xn�$t���m9�hסxK5�#P�N*Y�kq�l��;r���Y(G�8���=�ˏ[���a6��5�H�5�Y��F\3dj��k�:��Nڗ0�B�A ['3o.s.ݽZz�-}Ћ�^ht$S�E���|�ˬ--�¶d�eC�B�`bX�0��������XGA�gf��}b�٫V���E����Y&�Y7c����"x�#nZ4*־D����!���;[�����d\SE��a,]����ql�:,Q�r�Qi�v'G:߉��i���K9i�z�,�M l��͊p�Yӽ�'d�!]Wϒt��Y`_V�41��63kU�[Nu�1\�n�8$M��W`ec�F*�_t>P�����HuR�l|>�ġSB�?<���5il'z��hK�GN�3G��cG�2�܏�$���l;:��3"ŷ�(}�L�
��q��g�</�V���X���s�ε�{��}�zQ%IM5QMQ�CATST�%QMDM!TESEAQU�TTUSP��LD�A$�T4$1�Ae�Q1T�DEQ1$�D�D�AETQ5L��D4��TUK10U0QQ�5D�TPSK2U�DS4T�DTDE3IVYU4SQ3PE��TUDR�CMEQTQUL1EQUT1P1�E4QADQ4TMP�L�AMC4�E�0E%2�E1D5@|*���U *�̓m�8����9�-������i_HĮ�Ԧf)�)X͌M�Ǫ���*�5�J�e<���Xs�"7#X#�`�lv��EO�U�<�E��Nrƻ��YjT l$�QEG]��]�s�V�ucY��x�*���,)�
1��`=V�`.�K�D��(�lN{��f��r\>g�;ݦ���өhBk����BmK�C�Ҟ����`sB����^zz-NKu�/he�Wħk�W�0ķ㑓 8P%N�TM{s��#m�ó{.�
(s;2�u2nι�S�B�Aq�͂���P�]�E3M����u8QU��УX��r����9૷��9�Nb�t⛀�}w�+Yr1���4f5�b�@�XT{a�������-LZ�W�U �N�=
����&p߼��(*V�_$uc��1w1�>/^.v��{z��j�>����S��`�\;r@� r4f��TIs\!�ѧv4�ۘ+7�NL�f�R5;o�!�fЩ�����D!��71M�6^	�1�(k>�B�sл)��s-�2��;ƕj��Nl�a���a�]�r'�lA�\X�,��4��NG3���#utu7���E>��H#W,��q�b�om�t [+7eI�DU��H���K���s%B��n7|5�S�����ObO_�6���,��Z��̋�4mN�������9%GMl��1���{��*��O�+��"N;��M�Gj��x9���nR���	pLd����r71P��nۿ҄7��&nn�\�$6��Er��4�
���oU3uK�.��m��+˷�v~��_(�E������d�!�� ����,q��/uw܇�Q�!iP�3��Ux�}f]9���E�]�|�S��t�Ӭ%W�U�~-�ņ�Z���b�S����(�̊
�t]X�s{YUB�uK�!Wi��C��Ц�y7YZ.8K#�v1%J�f����5�G!�a��[��A?>3��
��iT��n\�.R�([n������XNჟj��f�&���x�AצH�v6(�±D	�z&��Pb�t��)�^_��,���Ω�|`��'��}ԇ��mE%鹆�+��\Qa��a�!G���u;�v��4|C�ʗ���,���n���L�'6�{��z��2�i�\�= ̱	XB��.�\;�%��٧�Ի
�}��m��O��\ts��u����p8�7#|��"����/�G�	�85ƽ��Z's�lubf����r���6Wb*s�Om�$�lO��;�K!�AB����%��׹[P}3<�,�����'�-:smӑv�F�Y���,wK,�){+�fY�c����N��0CFu�B;\:h�OB����	P�����u��F-�{�qr��ЈQ�.���d(�a��te�v��ME��!D웘�8n�$,}�k�k~��L)�7S&���4�<�]6���T8T%ƅ+OzZ�a�-��U�I��u����>�!�D�7Er}|�:�=����}�����$j��m��;�k�����`�l�lp� d(>2J�F�+81C3�`�	U�o�&��=|p46�Uc�.q�0���蘦��Fw���j�XǍ=�\*=侃jNv7q��%�/M���1]�{�|�sS�)���6f4[����kf���s:#�@X-�x�@�c/gq��!��F���#�I����w�.и�"��Y�$��b$�:͚��72t27e[�5���1g[�|��J+�Q3�h����Ӣ}F�����!ܵ"��k6,'�::0k#��ɭ2�2l������#z`�0�"�3����8��HB��i���z��	�P�Gk+4���7��V.;���M��F,68]Cu�l%#��<c�	��\��E��N�y�.+���,XS6`X��P'otT�g8*��8�����hgf�,�8��u���Z鑮�Z��oUڌ�2�W�.���A���Z䊙Ĭ�nW���*O��"O��t�֫0D�{.w�)������ͫ��C)N��=*��G��,ra���zq�8%�z���`���"[�D mWD�v:`ʗ�m��˩\-��$c��!�R�2")�=j�x'��b�hŧ�0a�H@r�{1*����R��}�Ѫ�/��ʋ[�:*��^}7��P��Ok���2��Q��c��w�l�~��( /��6����:y�z_��'����LsŃ����93͑�&)b��&&��d�lw%o��|3�� i�UP��Ԥ�y��"�\o���[*�w}�V��&60OK7ҍ�\�l$⑅wBXr�H#�q$"Hf�?lN�/bf�(� �uY��:��ܡ��ȵ��*�!t��m��"tA�7^�B0�I2�Q�2�ȭ�+ݚ��y���y�^���k� �/������3����b�Xa|tN)�.B�n2���iWro9���>v������KR"%��&�b�g���~چ�_	B�ZE��^��-ɸ
�.��PA�z�+�%�~��I�߽S����nfyu�+���4g�Ѹ�V<}���E�V&شE�p���f�2��2�Jc|�`�u`i�0˾Oi���ei��9��>]\xswәΒۜsH�:�e��[L�C��{��ES�I��R�|���mn�"kh��� ��d[�($���EȮ�F�\{U!"�9�@����o�(F^g�"㣐`�����Jx����y����Mu5��s���m�j��*H0[>����(a�*'gi�ت��C����z��~ S���<pƢ����cG���b_H5g"H�|}�WJס����v������_�i�_��-��{��V���^����P�7�]�>��ȯJk�A��T�@S��9q��Ec�KW���\9wp��U}&�g�;���K9kX�w+#�5�QF �]�G������l���,�D0����S}��/}����z�B�V�B$tiF�v$��6���lDJk��h|��J��bEP�m9�*d�=s�m�|�P�ϩ��Z����.;��Ԩ|����k~�V������u�@Q�%͔TMζ�`�ʁaٽ�x��n�ʚSKcWl�]ڎu�ũx�㼵�6��~"���#W���*�>�.U{g��Fy,v��Mt�)�x�F:�VGP�\F����	�VT�d�1�/N)��eXb��v��C�EwSچg#�P�Z�γbG
�/���v���r2'N.A*�d�ա�|���5[u���\��b镙}"Y��z�GZ;e��6j+3��w[�z�j֞<w�6�o�)�34ΣC�VW/�i�+�=sx)ע�h�]���9����R�|��t^�U��g+�"�v3��a:p񝋅^u����;�lJ
�b��N�aw�V���O���+>��b6T\L*E)�O�WZ�&ys���ٓ�k�]+��ee�h��+,w`9��r>�^�^�vP�&�u8�9�֙���6^L���a��ժ��=�p��|����l^`�8�Ω1y:3��]�
��v�����qꪓ�M+{YO��\"̰ٽ�~� �D��1���r�Q���C#|7mߍ��腦����LҊ6��Fwa5��������U��r||� ��挌�V*��N6�Gi��H�[n�j������5�� �_UŹ��t�����`�7X�
,}�3z�\�w\k�f������~�()�J����w�~o��Z9�)�9��&���qm��P�gj�
��ۛ�"�N��1��
l�u�%�㥑�;	#�<;��4D˽��׵J�bP��_P��T�v���>�*'�6�7a��h�55̙�(r��p��T�/9����]�t���;li�A�� ����]��^�+ѩ�(a���j�*��,)腑�8�(>��*��Vna��Ss�q��c�n5�y�j����I�Uʃ�L�v��,��s5d�%�m��qwwY�=zǄ�w���j�ӧ>�B�.�V��4w�[�s8���7��](u�gcz%���2dS�l�R~��1�z(B6�*�Q���u����ݩ�M1������Վ~���ܵ;�{�W�e����!zz,BWT+w�Xř���o�u��jon?%\CSV���5b�tu�ہ��VH���"(!*Ӫs0K�i+]���D�H��f}HV��B�e�qap=N{�
,�t::���N���2 ��{:��5k��Bw�NB�R
��-F�Z-{WէjD�Q"�>
Eo��	p�;z��lq����ݹ�G�*��K�!b:�����.�^�^�7t*
/���)�1�)l�x��W0j!�g�d�"J ���zB��+�v����ח�Eʵ�ʻHq{0��5^�.=�ʪ��3PN�LPm
�6����>2}�EP�B����>���v�Q[J*��s;ː�U;l��6�	m��Fb�mdS�:���
�̟h�������ՓA��y��Ã_Nbx���8��Il��Ԏö���fMCC�rg4��q(�%�E���:���I��ݦǝ,����Ui����7<��S�f�`����d�� 7w�gIS�<;Q{�rVq9R9�ʕt�����P�6�k�}�}ٜ�X�C�s����pn�z�*��=�4fU���<�¥���O!�\|s�������àb���/DG)e',�>\C�Z�N��f�|FF��6�F=���6�T�2X��*7f#�NE��B��q���&��ϋ�ȭ��V�&�Tl.��ⱱ��QK6����n����dw�g�m�C.��,I���ؠ�,�v��3ϴP�a�p�6���z�򮉃�|}"[�Ք{e��m��=CNkJ��<�<{Ylc!)X#��XȈ�5�hu����j�g�7I����~(�	Pe�Iq��(C	�؝�p[�:(���Ƀç�\��{mN�����V0�Wˉ3�MNG<y]Ю=*-�b�T+��>��p]1xV��/�}�I���T#,y��F��⵾�1o5~ݰ�a3^�6&�WF�h�_B*.7��ӕ�w}�j�fj��H-��o^�����|��VЛ\	
�!��r�
1�y**!�9.W ��G0X��y�h�[����y]u�4�8![��V(j��Y��]`V1��Dˮ�b��;�e��V؞��ejZzh�쫫�(po[�#��S�W%����iR ��%�V����;Gm�����9���t��+�%�fN���PV8-�G��h��v�G�-���'Dn� �D�£�2 �QP���*��^ӏ��u���Y��6�
+�Ь�����Q��a|V�ƬR���ܫ~^���N�7����GC��V����K�DAbkɺ����C��ɫ��f�2(T�t�7#��Y]�_/J���S{&.�Y2T[�y���9�h1b[��˭�Wν�]D�sY��� ���I
F�̱�'���+bGuY)y��de�{�.: ���^b����h���g�λaښ��55��D��W�×��Llg���!�`ަ!ʤ$J��㮮h��F���c��t�vtC����I�s�J����^Qإu��(ħn�K��Nv/�Lf�Q��ڷ/ }J-�z�9�yװ0y3}5�}�$��N`��xQ�;o����2y�o��.����F	���>nƻQ�r��������03�t���Rʛ��]E��%8�Dh�����N���6�{�����j��Z#�J8UH�Y���<QW���T�&nI�)��D�����8��Ecr�r�'@��[�.Of��oX�]ɨT'M�T�����9b�E�^�r�}���RIP�Z��{���7]8֬��p�V�c�� ��X��qAײ���B+��tQ����D��P��ZDNM�P+�Ҟ����c�*�Ԍ���م�ep����]f�@�_Zx\S�qyT=hW���̽�񫡓˅y���tO��(OZ|����>�\�>]� ���~��f����U}��f�j���}J���l2N!�/WG*��j]�Nn.���l�~}w�+Yr1��8�b5���@�G&s�u�fzq���t�;�%���*��+��E�:��Zu�Z�"��  v*��h/�e�荔�P�7&6���+�u�;���8��(E�q Lg�2�!�n��)w��xq��}�]e��pT��M�pvP�&���9��	���(l��Q�ф���wTB�Bcb�7��G�\'!D�q��Nl׳���P���9�%� �SG�f�t�u��䎁�R�W�P�dW�"�L�Օ�L�V��ӳM���)�G���}2OY$Bc�d1a:{#`��rrj��\�~g`R+�0���>e��F�=pMÂ3�-1& }\�n��iI&��_$����#::�jV"G�\�N��8��ejr;���_*��\1��c%���ڝ9�:=s�Y�T�<�#�`q�Q��\��܄����:��Pл`�緀k�<}ʦ.�ЧKj[�Kg:�+E���4
'��͂J��z���D�$���{fϯ:�=�	*�v����1
�f��vn-�l۴�w`n��[���:�������P�(+y�ҧ7 ���u���NU����k�<�$&DjY��UK �����r�H3ɜ*����m�(mysVb�:K�Ό��A�vsk(���2.���%7sp|�ڲ�>XⰭQ��6sj�=��u[y��w�������+���5;mѱ�i\1̂�D�6���u�m�欮A�f���M�9�.��K���������q���1��.I��Ǵ|��;M�'V}�Rb���E��v(��E�+j;!Ԅ���q�on=�݂�q�K���E��T1`;o�:�$�>�;�jd������Qs@j�ʾ�!� �![�CsF�{x9���$�	�CM��8����ލV��Ę(�'��,>�{
��I�nb���.U�m���խ�&���Qi�v��*Y�%E�󥔨�7hu���`���� ��r���7@�|F�{Gq��[��QT��O�6�DQ�j�U����=�G�RmrŒ�z�B��Ґ`�ӱҭr��v�q�����7�$l�f�䜔�4���˯v�wHj�<z+��ǃYO�@��v��5�g��}Τ��u�W�2Ł$ټx��˝�V%�Ɖ���	�D�t�̱.3���2H��d����a���|��ԋ�O����	���^n:�UWX��>�+��P��]Y8�a k8�����O��d��4�:�����k�6';�hsC&�]��LkI��&L�R���ڶ{��_r�TlEǝnK��ܔ�:�"��Mug�ڹ�6�ie������V-�(����%؞UP��I�����X"�(C1ϸj�pF�>����ƈ՚�P�Y�q:U�J]8�L��U��������2Ⱦ�‍�&n����]�,��QL<m� F�X�l����od�j��Q�bp�ff%!ʝ{`��H��߮��@��c�g�j�B�/h- ry�"G
�@����+��}Hދ�e���tv:X4z��afA���p�
����Jw��6=�)b�d�K7
I$���*	CB����;r��X��r��;P��+�ȭT�6�/e^��5�F��
q�}%5�H�h�)�)r)uQ��_�՗Y-��OO&�}7��흝��Q�舘[�����?{cZ���j� z�_�7��	]�xW��d#2��JG|��Y�2c�V.�Nk�̃fi�Ii	++��\���M���ه�����.�2�w�uϏ<�^˫j��W�����7����(
����.��$��)���J��i�&����((��������*������������(��j�(�iH� �*�b$j��$��&���*��b����*�b���"�j����32j���j*���ْaAI2PSE$EPP�DHD�QQ19dS0SIAEPE��TTD��
�)*a�1�j�$�������P��U!C���P���LQ�¢������h����*�(�j��#XI�"���
5!�
��>��gpѧ�h�֘�i�Y;�SVVt�1�9�.��:� nᰝ\�O;'@{��քuqf��&h\����3�8��vfn=��S����P�r��:ڮ���t�H��r*d����S�÷��]�E�8犵�Oj�G&W�
�F����\81���"��j�SJs�=3+��++d;Ib�9"=m@�+��\B��i����7{4)��&� _�T���:�ֈ��ǰ�un��~��FwܜI��6�L9��(EC��^�4�WM9p �V5��gY�0���Z�u�G4(���s�YmWD�
cb�
��Jj���h.�xpA�Ξ�����'Ɠ�%�S����o����[��lS�A�H�'������C�
=�D�׏��섵�ͽ���C���n/�ϥS��r�S������w4�Ap��D1	B�L��R���@��k�}���]8�S.r���旭�GXO��謑^XT�p�
��U��q����f2v(f�:{.���zN�Xt::���N���S̛X�i�ݙ�IU��9PV1�0���GS������==�\V�^"����nVS���e�M��
���wX2��u}�|�7L��v�2�R=�@֩�9I���1c2���t;/�Abw[΃{�����ˡ���B��������`[�J��+Ή�[y�gwP���S��X�[2D!O��ܱ\�!�k�Zy�q�����ϭ�k�=���`J�5k�B�Lث��X(Û�A�,���pd8�:����X;7v{�Nd�[��l�Ñ�$�t��|b�p"�g��.��Ù��RKh�.Nf��)_
c]Z�`s3Rt�a�Й���q�EPP22�&'��BM��S�9��l6�dX�e�_�jؗ�����LU��خf�j�B�tG�����y��/�Z���r+dtw���Lq��m��t��$��*E�^����n�9�d1�4�
�e�8O����bms��v�fM�]�[1�^P�Z5�'c�W���py�V��͗��[�8C�S������+�J~/�,��M"�fĂ�z_*�)8�a5C&z��of3�ߡ����ɷBv,�.����>n!���fMm��s;��^�cU����q���/��=I�w�}�A���lV<��`}�*T�\��쮂Gِ��Ei}[�]�^4� PmD�A�W8�9��V�^q���p�N�!n۬z�D�%چg���(ڱ񂷻�l����]u6ZC��Qٚ[�	^ѥr�����:��4=��zy(��J�]ue��5rl�Ԛe�9ڂ����;m��]]J�Za'�{����n��U\<�J��!��۴�V7�t�'�tJ3���V�ګ��X��A=��j�N[� ݘ�r�8�P�kz��pR���4���6v;����J��&��nN�`���%&����j� ��1H֤q�we�B��㦞�ѶRމi��Y"��N� �S���pI8ODI�R)Daw0ԣ�v�l%�^K�v�T��/�6���n�؂5��ƌN֛�����<#�-�Xu'�l������o��ݎpXMƶ�;rp뙮#5-Q�9=�ajb�Cp�7�5�J�1�63i�c�1I� <��c"��s�X�x8��'t�2�d��0�ٻYY��g��t;-��n��3�T�k��k�_oԴ߱^�^�3�̥9*�}�uz=cUw}+���P�.��;�d�0̖�NHx!�>����ռ3o���t�<̗����.i�C�RI[�gb��U���s��	��%��Wvʰ{�~���\��[<�&�L9]A��v�ݝ�:�bX��JWҡ�;/ �|:���L�m,��RnJ��ŕ#��N�k):[��w���O�%_�;
��)k��}��z�M.I�p�[����w�ӡ;w�=~� ���S�[Ѷ��fF$�6�O9k;S3��W�[y�[�kv��v���z���S1�4�����*�o9�'Թ��(�m&�:��b�Ԓ���Z�zdZ�y1N�T�q&�?FD�7#���BE%m��WWj�����:��j�b{ם��m[�Cz]�;���P]2�(ݾn��Tc�䍙���q���zU?s�C�§��yb��@R��d4��2�r��}bMU�!dd������|�z�VK��_7զ�� ��/b25��ѫ�c3���[q˺�
~O*����ϗ4�:E����.��Pq3���]WYKVm��^Z�vu�X���n�
���:��j�KBݹ�4�����f6F�ap͎5{2�g=3���71]�"�n�R�e �T�����Q�Ź�yF�2���,#�I��������7K.ݭ���h[�P���"��lej��h�i�p�)y�Ȏ�@:7���6����grǑ�6�'�������a�'��"��׶���n�8/�&c�p��Ū��oz��&�h�7��^;7�]�7nѾ�lt9.e��̇�7>Q���z��Y��x��^�²�䡼���c�F6�95J����Lh�W��i�����TH����	̤���N�\V�Y�of�L��~������9���4�6���[���lŎ�r0�WOn���*�C��n���"i���-�����`�����Zt]�W�
�z���0vwB���o	v�J�";]6�Kvv姘+�LH�q�C�z�D�Wm$�͍��Cq�]>U�Q��o�Z�q{j ^{�4��BI	���_��w�}�oˢ|܀��	�A�h��c�ǹN6�e��ΪmZv��=�M[�oK�4u�Au K����:�/�[���G��&k+mTݺ�"m����L�~�WW7N��YJn��K��t�&.�W��G�x/k���j���V+5ì��Ę+M N1��je5v���$PK�ۥ��S+��Xn�E�6�X�Y�6l�������P^N{��qs����e�m��ΡO��eow�T;|���Ub�����U�lu}�؟{�z�6IyJ�: ���������Nml>}���X���O�����7�\+=�����.��S�%{5���>�u[/���4��Ԧ�Mљ�В���P)Dm��� pq!FF�Dt�*����\:�pgn�t�B�S�
Q��2����	J¸V ����D�CG�{��\�^ڍ�KquUYf5>=��'����������	>�g��Άyq�+
G�$���y"�tjLM�
Rw)�I�8`�����k3��jR�6c�Iݛ;{�A4�x�������Vc�sJ5�P	�"�v�ZM{����ޗⲥ�z�z�p����k3����ƭ�e���k���YuS=��e��r��RIa�O���ۥ~8L�}b1�����"�����(�Lw����B`�°)s8������T�6�O9E<�X׻�)���]��R�$U�M�T��}�e"���5���wA�W�xV.�O+T��qeg�jL��|�h�"����Tw�m��%@�ŶT���]'g<&�11�.����[ƭ��m���}��O���ͪ*�Jxpgvq6_\j	y�����Tŧ�o�Ւ�ާ`��C��Mq�3bA�Y�|��լ�
�)κ���:���ꠧ������N�l<�An���"Cc�d����Gnf�G>��6�z��M�u5~}�=Sɪ|!��6��K�Ȃv��
�eA�(M%o��vZ�V�0���ޢ$�9;H�X�جI��<�d����A)�byF�wr�M�o�9�C�=��sm2�~͖�6-���x��AH^� HiQ:D�[˂����חP�����O]�(���3�֝i9�dkR:�X��\��8�T����F7|�^�5�]z���j�3��X���p�rw
7.h�Fg�u˽�֌a=�m�	N���h���#Y��A��dE6�������"싪4d,�Z��M�'84o2���T�,z4\��	Tڗ����X�	��"gvM�L�W���K����M:�����X�}����Fu9�1�W�:�V'����gX��6��[;��Z��ۃ���Q���(��$-wj³IIKL�^R���SU����8,&�Chc�'��j���v̛��2�P�Mq��W�1�63i������=cU��n��f���T~:�^�t9�p�g2��d]���o�o ��"$�����Ed\�� �1��:�7�w��TH���l�̥`�4�V���5u,U�oENjh`�����0Z�:[������pycDN:ow��4Nz��{=�#��wl���M��NZ};w<����lO�x{�s�Տv��u���w�)P�s��y�aj�Ko6Kv5�vZu;P]�s�Ƚyd�c���.�'�)�GV��Ɔ�Hi]څ*�k[T߉�|j�Nu����V��mؔ��A�w��vl[�K��a�tk��v�ȥ�$ O=}<��t7�����%��Y���g����>�@���J�F�dF����K_�4��v̑��Ja���[^^Z�e,�Ɔ��0�V�pm����9���=XV��J��|b��U
�kR��i�n�WP_m)!�@�b�y)O� �t����lv�專�4��˦6p2-�D	��6�ُ�Y��C�JULm�t�Hs�U��,TU�
B���x���U��r5��5BJ2��MX]m"Ң^&�����X� ��3�R��og8�q0�{i���5�U��ߗj��i�<�gXOD�Rq���k#��zkO>����!�P#�ՊN޷~H*�\u��PжwT*��)\6�6b�"R�~6'G3'�X#$SrG^�7���{\�A�}�9���z��`)8hk3�M��d�sY��Rnݣ>��gTM�s�m�/�j�Ja�b�pE�5ΰ��S��[9�ټ�|��Ɩ�L�.B��^�g5�V�sYX���ZMuF���Pt�_����S��wZ�����}v������á}t����5�������&#�����gt�{�FH�a�qҰ&�q�-�����S��[���6�M3x�+�ك4{�l���_-=Y�c]�c1��_F26��4m��1w�� � @�#;+6�ɜP�"���1��b�J�b<y��ګD�yҭ�����r�RE���T�
]�>s�����x]�pv�K4_`͗g�BM.��Ҝ�wU��Y6�T��pB�>�-�-�����T���Ԓ]�{~=Ib��7-�������Mq��@������� ��w�ϖR��C[�&�ĺ��<��:	��KZ�C�;~]n_� �����F��a���{ј��Vv��:�V5[MA��ޞ�����6$p��P]P�p;Y��e]��޷-A�L�����,&�{���{�kɺ.��\���X2��7���_ho�A:�$v;���j��eS�Յ��g;c���K��j��;KUW!��ٷ#�Q:D⭇ˇ�j��e�;��
��S+Wv��=�/�8�� ��1#[��X�c[�ë�����Z��U����s�����zZ�á���}��='�Y��Z���9[�.*Ч�����:����ؐ��X��g��ъ%�}S'��R##1����&���5����%�f�wη�e ;c��+ѽ��,������s쩋:�+(w0쩛zv��C{� w�C�z��-l�kN�w-p<�Y��a�PmbVvR���C���e9����Buo8t[��U]V'K�e8�M.{�-_�nwK<BZ��r3_9b@wo�;-�M`��n���Fاs�\����I��1Q9g��{2Єzh���A��`I�C`p�د�uY��[�O]��
�.eIݸ.AH��Oit[큙�[PvӤ�Z����uӫmwh}���\N���%�T�WM�c���,�A�g:�P���X�a����0Ε�zY�xTL��$��ELMouβ'f�]é�nKfk�3�tsa�����l��·�"��0C$�	�����l4v�E7{��,�twu��H��s�5�I�]��egu��Au��Cx��ٝ������Ǯڳv�uƁ��K�Aˎ�����U��Hc�f{D��Bsy݇zF�_c��ó��ϲm���rx����Ka[k.u>	��i����a2��s>��L���Lj��8+�X6�^:_p��m�7y�3^�DU�w��.�[��u�Wwͼ|�&���wv�m���z� ���0���f��nʽ�f$�fc�o��]�8@�W(v�ݳ���K7ر�p���a���Q�uۚ"��ǒ�W76��@RV.L��������Ӌ1W0]�NR{2��q�-od6w	��]��I��sIPǭޫ�5�I�)P͸�XNS�C;]i�eK�\��(೚)�����
�ݔ��q�8��B�M�3�Q�u�N[���/\o;}n��%��]������yj���J�V�[{Q\W!��P�O1Ɯ����B��U��KG�Ž�w�3N�����Ʊ.k�8�7���=��>o��L����z�^NS�fE����IaU��]�n�ҳ��m*� Et�"��{yzr=����6SNN�u�������F6'x�%LN8����l�m0�Zp�*_�+�[�_Tt��T6�����g7\��x_I�����4,c�	�gJ����[��EmLڛ��c�����zU5�6��A.��X8��4�$x�}�P2]
�K�"��<�`�{��ʅ�ή7̼�A��n�%H���ih{��P4ru�^U���"Eӏ���^^�YQy�n�%h�t�����CF�;��QPպ��@��/x	���U��F�&�c���u�8/VҥL`��$:���v&�ŜQ�ޘi�B���[ �.��̚�=e쩦������J���ͨj�FK�&B���t6��#�O��{Ur+n�s7G�N�����jp[o�+:���d7�r�	�^����Nw���rsBәӜ2��]\#���,g�m�����:k^����ny߹�o^u��kMvT4��f`4��4�EMUQDIffdR44ELADd�PP�e5%KC���R�DTIT��)0QNF@R�II3@D�@E�KCE�9 SIJD�NUI@ST�,�DL�RMT5�499��P�	IYRPSKIfB8JDTDE4�B�dERQMS�@�P��Bd�ET�A�4+���D�E%*U8Bd����N@d@�!I���`�f#�FCMU!M,�P8���IL�IM99&A��@'�rm�҇�]^�����u9qV���M��Q��/�u���'�p�]��L�T�[ ���$ �_W
�h�ޕ�9�;�����7��8`�7�<͜�gC�uw�{U�r��&�P8�ś`�]�����҃Mc��n��u��с�sfqE��4)��:_�L�̮�[�v��e6;7�u}t�%��4�/�[
������5���Qn��$	���bo˘c!L�����%!4	:�c�o`�|Mz�'�FKxq��k��~�j1�xW5�SrS�ڧ~-:�sɤVli�\d���9�S�~��Od�����k�W\im��ֱM6����ulH��C,�s���X���թ|�$-�]Ѷ��)�#��}�Ꞡ��by���B�6���.�0����z���J)(��z�m��&��z}յ���v:��`����"^j��=���a*%�<����~[mS��ZvwC�S��h��]�'��ֺ	��r�ի�T������uTaQ�vo:j�"�� �������ڴn9}/� �Yz��E]����:�L�3��F�)���a�Ie�&ޘ��U��f�ob�^�-���!�B`��rr�ܫ4���֖��|U��n@콬�V(��Ϻ=�4*"�
W���ҠN�n�l�(�2��Q6�s�@�n9T���rvm�:g3�'ZE�A(�1@ְ�����ieR+3CIE��r]�N����H�g�ۜ|ӀB$pŐ���c/VefgZ�=O�R���sש�AS���mt4-؇b�f�Y\���.����rL)��$�sY�ܛ��l�o�Kp���m�O3cR�0���ޙ�煽�m�7������m6,s�/�E_��Ӧ�����'�����*�\�t9����V�.�Ve7��V��6͖'/:c;�Wr�!0��A5��aю��Q `Xp6D�R�2�������S�ƞ�sJ.��au� �ڧ`������|M^D���
��
�N$-A��Ɩ��ھ����r�c[z���z��-:����i��\(R�e���׀Fʗ�3��c�����Mp6�| G.�Lg�U1\.ƳA>��m!Z�0e� ��\���ʹ5��j[h���05{�=��*��X35�4jC׈5S!��>o:'�-�p�*�\�;e�.�hR�C
ª��s:��=�V4�I�
�(w��C�vŜ�l���[��ۖ�yڜ��4���k��#�-gl�qF��r� ��$'�BE>u�Q��I����X�p+��C��Ѭ�3����P�~7��U�JkW��˨��=�6�k�Z"�g!���;�]���)�z�o�F�������p�v��U���NV;ی�Zټ�c]�U����s�T�Y��QWH^�2N�/;!M���,���t���n��)����D�O��+�M,r
�nC\�]�H�7��U�����k�N��sW�+X)��z���=s]Q2��k38�f-e��C4�#q�)�b��o�AW_�]i�1Y���LG�y��x�;����'���7ؤ^
nO^�6;���L$]�e���U�q�+3��nN�d��<1`��ټ7js�6�+�8}Qf�(�J!�3S} �Ms�^`�{ޚ�i��F�x��������b��MFa���!R�&��r��.=�[K4��ƍ��(�P�N�n:������hw��:(����*浣��-�E��;�2�:��VP�+����IDZ�h�~�Rn-��l�����8b Ncw$)ں'e�'����Gh/Z��ܡ�\�ky�c���߱֓^���+K�ה����!�݇�A�{x�X�0Ý^y�'}t�������k�$���ȝ9&��p�8�A�C3��bqӜ�M���E�1�vY��˭S}ϴ˄���*kcj���6$�gÁFp�g����a��o�Ƈ��&у����Г���;3|�E^lHn��>T;
5�7;Vf����h&�c:���OX/�i�ֻ��uth#p�>�P��,��3�^cV�wV��H�C�=���5�V��{��V����F����2O�m�1Kl���e��:֠�g���l�}mQu�M*���z��5q���=}9U�r�T�q-�,���t�Z���V�ګ�>�K����1T8of��8�+��Lؼ�;����[��E���I*��4<��0y���E�p#��X.v֎,R��M��_�$̺'��G}�1���[����Ev�5[y7����m�ht��lj%����w�T�tB�e�a�����Y�BVI|��[�rN��̉���w˲�zp�۬zq�S�g��.�̓j��5�1�ӔД�z��u��� ��B�S���ʃWn����J�X~<��'u��,�G_��\�=-Xw�v �Fx(�'�X!��[�U�cx���B��m__pt�\͍mv����:1��ݽi��MS��4��O���N��{�k�0Sp@o�Mu���F. ��B�:�:_���ްo��Vc�lf���pm���TnfD!�=���ͩǌ�Xu82E���R��ݬ��lv{y�}E��5�m`���u�����Q}Lk���^�]Q#À��R�`�zR��l��d.���{P��Ja�m'�{]i<�pycFp�8��L�y���5�M$�ոL%�-�MS�Өy۩�=y蔬LȤ�[�02lM�oa��
 ~ti̀U�]h�=]ԡ�T�b��zs�/:�(F>*��٨;�;�}-�Q�:�f���[y�Ehu��9������+�P���"N�:ը�@j�+%�M��ԓ-]4��Znu_p;K�t/���|��d��O�1[��&��_I�����!L��k�����;����@�h�������OT�/t���(�43˦1e���پ�~�����,H��o���k��+}i��z���V�ʮ�ij��w�4�j�y�Y�V������yT̜y�v�)��y�*֔1��7�S��M�*{�h,TE ����!�D��E\�I𪹒��eG(��|�e���沚V]s��gZu�,r4 �B���S�\Nu���9V��ִ[�yT��.]z����j�3���pI89sr�D]�������;[#k�׭�	N���� CB�ñb�u䡻",MueS&�#�8ۖc�X殛�{h߻���8,P	�-@�ˍ+1��=�J�޷G�srp�H���16ݛ�v���x�ީ]�֮v�2��vLH�x}[Hf;�Zy�{��&�^���f۳�z��K)�h%���ٯ^[4�մ�B��)2m��Xz��6����Z�]�g�.9CqGp��]O8Z4���3�m\����ݜw�'�:Xhn�/+pt���KN���[��]�f3a��+~Ơ���p�8w�N�7���Vm���E��:{嬤c��Q�^��lP��u�q��8`XF��R�F��{�qQ�4�m���̡��u�0�ڧe���-����o#��]Kl�����s�+�%�s�����ߵSv�w�ӯC��N���;e�O+Q��zUD65!.�
V�U�R�����[�kv���x�ڮ��͸�ku�ryW�:��$�����(���GSO�M~�ᢹb����y�S��k{��lpܰ%�
IAm�:s��2�q���\c:��i����O=�\7�؍���%��[�¦)��<o{)��Jj���-���;�m4�� ���D����t��v������+`���`l�v[K)�d�}����+���8P����%9eN/Q��H�$��V�Z�8۱�Rc���ĭ_[�v�F�A��R_	;�[sm�g}�f���G�����ݔ2�:�ߞ��+�3�wɲ���=6b���D���7�^��z���Re=���r��J��;� ��=��Lֹh�K͔�����8dstFϫV��k�5~敬�Pg��y�H�Rn.��
-DP���::8c�#qP:�7���AWX��ڛȺ��V�@˵l:Q�����yV�ĞFH�}��'�Y4ܞ��j���L��Ū�����d�m�}~	�mz��fOHሉ/��M
�W;X�9�HR�+�ٿwRv9�qoE�3g���xZ��a� v��z�w3�+̤��g�k3
g�j�V�sY���:�k�Qݒ�g=��s]��t�g��[�O�aA���`6���[�k�b:vUl:�N��!RIa�O�0"qҜ�M��#[~�M�Ʃͺ����,���ڌU�;u�=y�$;#�DN��=���a�)�P2�ZL���o�Ւ���vZt!�n���� �}!�'"�)����S����Q���c*3���͵˩�w�І��_D��y�����C�򀼠���$ܚ�6�0���uf5*)�g�S���ī���H���{��-�ҭ3�t��G�Y��E����*0�������-]Ys� m�O�o�s'6ȃ�U^��g$�q,c������M)k]�}�mtH#p�A��v�'4�u=Jf�z{���c/Y�vRu`:|�����w�oK���>��ۊ��	�aA\�49P%J�3]��WN��=�ퟝ�����
���xR����a�#�/k��t�j�g�X]mU�}����{��.��l�I�����)�����C�D��⭇˂��w����6��0(j���$��E���δ�A�,r(C�#[�:@�T�#f���dl��:�*�m��=V_�����Zj�KV�v ����F���ō�tW[QA��Dm��<�g-�J��B�z������-�s�u�߸"��a>���T�x8{�b��;ᚷ�"����R��<��-:���r{��؂f1��*��W(ʖJ�s��k+�1�63ic�0���/�]l� $��Ńx,�$oQ��7��n���U��V_P�Uժ���=١�Tr��i�9�0)ED�~��n�b}ҦRBg5��n�W��}�S�k��qgnJ�����mЊ�G���ݳ�N�vB��*���&j�*�ohU�y��+�oA�YI�K5e#S�[U��TO�3a���V2.�We6;=��̞lݣ�2�����s-s3e<}�5��x�I������+8L�}հ&�w��#��q�pgrQ+z�x��:�OVn:�P��FKg�6�l��ܚkx���;�1�d�~MS��C����+6$;�7q��޻��ۤ����6*_:����Q���)�M���vZ�wKx_=Lf�Fa��0�$R�;m_0E:T������:h�b��GX��=q�>�e����Pv���e���+|Yp���ی�f���;�D	�5��-�4t]��{z��]�Pv����ȺS�6��9T�T��:�O���Oz��b�( �{x�)�zzb������y{В���Sv���ҳn�י������HC���`���>�8�����S�kF��6�YHՌ�$y�3b�
˴��tU���`;�j��2��r�e��/��Gur%=��ᇳ��ͥ��_L�O�K�u�X��ʥ	��������	:6T�VKn�A���HI�^p�1p�HA˶�r�����l�5� ��LK6���������]�%,�Ǳ��$�o���:G��D��<	)j.;��W�n�n�E�W8,��Bۗ�wI�Ik��`�c&��/�@�#
VZ���&�:{z���`��5�;�{��鉲
9b�M��s*݈e��n�|9;ٔ�*莘Lt���^i�&�d�xn�7��4�]�@]zL|���S�%s�5�-����6��pt�9�3�f�}��sh�@������w����(3�SmKH;�3*����E �(D_;�a�s3�r�m5�-f�#���q�����*v� �:��;�O��0�������i�cU�o��B��Ys
�m���f�%�ݵ/��\1�]C�3��T�3����F��]է
�|gb,w �xJTTy���*�!+�:n�A���e��lF2J�[fb�ڷKL2��î������ L�]�������d�Cs�H�9�Ż�=�;�K7���r;��gZ�oD����tU<xw�"�.W��������ۺ4ƺV~X�b�s:T���h�p����g�=*<���yZ���͹�aq��Az�<��ʶ�V;�ݣ]Z;�N���i������������i�x������t:j�u��5�ΏYl��q���Z���Y�W��%��j˟7�!ϞZY�j,�^�]^0ȃ���NՊ
��
�{X�����Muܳ;�+Dm'�8�$5�0��ks��f�`�N��3��iL��;Y��}�ƚ�Wd;;J��u���^ �ZT��p��m�&��J��n��'Xu����W�� ��{��#��N��]��r�Z�GM�g�ʀ��b��jۆ�1uc�)-�����'IA�V�9gK%����4����FvvR�%�=�Cګ�ߥ�MrT�Vl��j۔���M|/�R^.l��;����3-Q�6�ꑦ��r�v��ќ��a���c�|�/�ٻ�z�aڦ���#�#��׵6�����3M�¾�Ѿv����C��dy�k^�,��唅̣,&���G��(��4�>nnU�1��Ah����>�*ל�k�c��e9��'��ջ�M��E\��V�]����L���!�V�V9�>ʚN�6Kd��^�Sm(�e<Os;���c{�'}�Vss_� ��:���k9˞��"�ծZ,�Vƅ�L���uĬ�os5'o��;��l��}���uÒ��F����귶F�{f(�M�Na�G�]ov�ͧ͗�l��p��ཾ�oH?�$��?"	F��X���L������G'$r0$��(
�����r31r"L�
(ib(	������2
F�@��h��(JZ��`��\���+ �i
�3��B���)i�
B��2B���������ɠȦ�����(i�!�JJ�(��h�)J
 �i�L���
R�����")��@�)R���Ph�h��rC*��,�2"��U�
_|��cO���_\��aز������E�xprLMv..�z�ݜ�m�[�Tj:�oaXZ�\\������J���[��g����YNk:��e�.]z��t�3��X��N�E��&q�xN�֔�;����tֹ#�[�$;�}a�U-k�ݹ��iӑjڕ7�A�:6'F#%�xm�"�m�����]��+�l�s�׎�)��C�'{Y����������~Kǲ��*���郖����쒂V�	�"�ng�u'��.��m�	j���4��^��\�Q~���7�u�lSkhc��c�5���*���.�����@��}��<�����oݔ���a�"����-����h^D�`��rLVU����
�(?���aT����Am�U7oU;-0�:�2���s�63^�c{g9�Ma�!e�,��9oaJ�Ko�o[�����asE� �&���|�W1;Vzq�b|F��
)�iM�w����T�J!a��/}�^/m���.
��}��_Wg �ƶq�/�=�.*��euu�vPWL����wV�<8�(�3]=�[�7��g�L���C�!YqM��8�K��������B�R�f:�Ey·Y���>�S�k��SW٫�U������$���؇�U�6'���QB��^�ގ:x��^>}��(���U궬s	W�)�{փxX���� ����]T��z
�OT��%��Mp[mU�w����y�Y��Q^Y1e��8�y|��<�:D�T6{��k����������i��F�*Yq�d�NO6r�<�H٤HԨ��
�U����s\ҮT�ڌ�����F�^>��o�n��� �[#qP9�b�6���(Uѝ�{2q ��I�6��X��T%�nÛy�Cpd\)*�x{9Gѷ{�'{����
�ki>p_XL�mw��ᡬ���ሉ/E�
��fUM�ַ5�ܑw���S|��;z2k�a�g=����U�Ph}�޽��*g��aYDũox�ͤV�y7��mc8LC5
b@�2[�>��V���8�n?fqs>�<��#�a��\�t��S�.��x��8U�v R�t���+�
�^��]zJ�F/��i��ܲ�p(��&�
	(7ꎷj%��]ݕ�S��d �m��3�P��Y��;�:�*�0�n^��j�XO=9���w���}�o0����kfBsP�f�E�V�o-�*jz�mi.�$pX}����J��f�~�Am�Tڛ5���mťm�o%0OJ�|�wk�;�6'�;#�D	�ݞ]�ҡ��}�g�4+S�[�nO6�4N�<�ԗY�>4�
��,�'�Ak�{�������m6�~�)�M5bZ�bi����E{Kw��{x�0zs��`ת������N�k����ޞ����ՙCc�MƈofV�M�1���}@�})A|��ګ�;���Ү�c��HX�o�j���������ל�ʅ!{x�	W��-U��au�V)�2N�U�ˌ]('m�o��Ն��QR���!�@��Ga���FVw� ���Fa�vo���9�a:�ic�B
%DH��}� ��jy�5Ee�t[� ���b	N`�teX{~ݣr��$l�9+�(خFc(��yc<��K�W�m�NP���ܛB����tg�WC�]��j�C»����̎R�lgb#W�����G*;	f�iRV��{lf�[{VSݑ)S�QM�����ypuɣ�0�C���8j}��!�+l��)�OR��EoO^�����{͉mv��6�fӳ}P�\��M(�e�;��v����m�u7|ఛ��m�����z7:�r��+q��-�x[��n��>�YY�ٿf��<cr(���ǷtVeg
릠�Z=e�U��
t�9��b�U�j-��+$�[_N���	��~Mn��۬'�TH����Tܭ׻�W����NݎAfr	�T�:����|M^G����(��������M짵}�nvjV�C���ݦ��iס�n�ic6:B��4�\zh��+��rDw	Np�Sܫ��b4��F����6�yؖ�S��-����G�lO��"G1����>�h�e&��_�W�?�>�i� ��'/���mN��<���Cʇ�2�Ǆi�W1���/f	����WT��L�xǐ^Ӵ_�'�������������Ĭ�2�r�8F���7h�O[�܉�4Q�9�e@rN�����dEY�N�y���7���Q^������U�4��w�}�\lp޿J��4��f��k�{7�(j�f�ķU��j[Ӭ=�4���F�����̥�=F,޲b�����+����������W��U�f�*"�R����Ur��0 ����7ϡޑ����1�ƻ���
iY���g&p�X� �L�U�LQv�����^\č�#o±�l�v��j�k v��=�ŉ�ȳS	Q����Q���c6��;!H�R|:���AS�>���k�kn�]`���-<T��%�FO1_��W�xm� �{�>��n$;ƍ�d�;�^����;}!m������Y&۰o�Ģ�n��d���I��j"Ֆ:�,s�(&��u�o�i�ΧC��әKp�����:IM��Ɠ�����f[��>�a��1�i�w�׺��͚�[��ȍn��(>�zK�*���8��@�T��U�e�L���-�|� r˺���X�9cm��{I�|�����ړ��2���I���훒�����i�'���Ǜ�-�,�Zk8��y�I�b�a�Tգ�h��/�w���6Ü���b�]1\u�����H>���N�k('Kw��e,��n�����u�Q+��XF��Am�T݇�������lNt=�ǻF�G��2�+�P�7fyP�)X%���-�LTt����oD�������v���z�Ă7 7�P�|�%�S��f&��i�.��X�:NƱN�ԕ�-k�C�*�lO�n!�
E�;̣}����Ѫ�Z����k�I�N���\7��lH�ꂶ����j�ź��kP\��;�F�N��Ub��6K�����ׂ�EQ�%ź�s�uQ��������t�j�;� ��E�E�&�Q]W�v�ֺW�c{4��K\��B�##Z��+P/��ϵ�W
�����P��<x�n0�s	t�&�h5i�!b�#qQ�M�����tԁ^Vb[1����^4��᝗Wj��މ[�ӂ��LA�Y}���hCz��7���;z��̊�Y�gj���2�_NU����	����"bZ�>Wq���>ԜfNǬ�.�-gM΍�R��Y	 ���q0Nv��~�S�â����2k�S�s�^c��u�URз`9�$r3�F��Ob�F[�&ݦB�޵�gW T�mic�۾p_'1���������xb��uܣx�\M��D��\��e�>�c�Mn����z2k�a�������Z#h��}�(n� )і�3z��"��fSf�i~k�&���h�:&�*f'p�^��LV�,:����l�̥~8�o(vR�o0���Ҋ�����Y�\D�L�SWdKό�9fW�*��ԯ�Sc�1�w�b��n����W�����췔�ݮ��{6$�|%FK|,��f:
��r\,�T��}4�%;V��ݦ��O��n�H��lO��Hm�Li�n�tR#g�F6��0%�Waf��o:KV�N�i�j�zi�]��R�"�瘟���qW5Ƞ�x�"�A�h�e'Z��W=����R[kh��G�U{��0����I�(v�����Ӽ�gE7S�|/18��d�ᭈ�L?-�ک�o����� {��'
X��s��R��ۙ�n�wIM��N���8ʰO������-�}���6��t@L�+s��]�v�.�O_L��!+R�Xu�C�(.�K"R��g}�[U~�q�&�5Bqn\}����Y����|V[����K	Q8�������pdtB���� x�̉��vx��S{����KH)���$4��"qQ�N]�wocj��x�ry���sJ���:�u��A�,r

%P5��[�q.mP.)Y�u��z֋�e�-�\:��\�=�j��g��������LAu��3ܗcx�Xe��Z���mX�����ؖзnpN�)�/�7loGs��a�HcJǆ��nH��F�u7c�+ɸ�3�V+�S�R��Tqu�xT�������	�n�o���v�iA�*��x����HOgr��-t?[��|�I��������R�2.�d�"��������C��4�Em�~ԃ�_]6�p�KM�c�'�^�`*-����{��0�k�!+��E��Nߝ?�Q�3ڡ.��{7��l5v��ss{Oe�I=~H�6Q�]9�<�����M�/piS:h��F[J�]�8��F�.̝�ͺ���eJ&̷�V�<2��к�'\0W���{�Xy3�j�w.�a��:H �:�܇{5�fr����[~��x�gq ���u���HA��4F���LS��\���As�m�K�l�X�A+�-�j��Өy۸�EVA�f�5J�x��]T�!��	q����C��~�-���`�ҭ�:������ٺй<���\ytH����
��m�{
li|�-]&�t]Z�[֪;cRQ�WN�Ԃ�<�c�����IE��!�	I�m��MS�b��%T�[|��=��Y����ѱ#��%2�M�Q�Ӄ�j�������V�T�ҧ�I�'�GB�DW�
|����U޷ø2y7`�ۇ��W3�	ު�|�.�k4�۾nr�Bu�,r+
�l�����$�0����L!�����X��e�.]cW;X�s��q�BlPss���"��n��#�3'qYEj��n�
������Ww$H3��.b��`/��7��M�)^�E�c�S�"������w��`�ؕ��"���w$p6Mz��2LJ�����)ӊo�j5&s�ϱ�R`wk���8SR���.\�c[\�=��'$�]f�>D.����*����u.���jlI̑�D�F#�/��nM��)��}��o��y{��{U�S�pXMƶ�;��CY�82@�&ۚ�*����^�o��R.�m����l&��u�y�;ΧC���LT����7�R�b\�r�c�v�e'�7�}�ƶ���i��w���G��L8�ac��7u��aGәJ��E'��H>��:�*V��n�ӃsF��Z���̮b���P���qӳ�Q���[z��z�������J�j��vշ��x�s����lH<<
"p�fyP�)lKn����Q&�l��9��>?g��W�+]ǯ�bA�C}E	��v�F�N���y;��k[�NQx���GSW�S��+����Wz6$��}���}<8#��P�ߦ���K�gfŽ4�3_T�\����:�������
�+��* ���* ��@TA\Q�
�+��TA_�Q�
�+�`* ��������
�`W�W TA^�W������D��* ��Q�
�+� * ��W��(+$�k>8���,�K�B,�������H��>���@ *� P��IA"� 
 $� �� �����%(�AT��UB��"T��r���Q@��(��$"*%)BTi�)J(�TH�UIP�)D��EU%J
*�P*�"CB�Z����QI$���B��J�B��$�EJ�I
$JR��$�E D�J
�	T�є IRU�@%D>F�T��   ������R�F�6��`��P4��Z�XSX[P-�0j����kemU��4m����
DTlʕ%��  n�Z���Ml4Xl�
�ʠ��04�4��Ŧ��!k`*��AYSZU,�4�h3Ue��,���%P�)�(U�  ܞ����6�(4�l���%mZhk)���@��*�BSYjT
�[KKZi��!�
(P�B�
(P�B�q;�
(�
t)%(�
��$T@p  ;v�
(P����p�$(P�B�
06(P�B��E�g
(
(ㅵB��m�
�F�@¡�m��aJ�J�L�
��Q[�%H�P�"�%��T��".   6�
�U�5QJ��
�0�Rʘ
��%J���m�U(c*�jj(�e**J��*
E  �   7\P���QT��V�T��ST5U!�EV��P
���jI �Q*+j�* �d�*�
*��  �� �5UZ���5D�T�)��A&�Y���&�a�$�5�[)��YaEY��Q�B�B��  �v�-�`P���T� &�Fm�P���Z6�ʦ�Em[f���@���d��4f����� �M5R���i�P�  �N���[F�X�c&�MZ�JP*�ƭ�m�6ڰ�hkA�b��B��&� 4l�m4)CV��&db�V�im�")*���T�� ب:(kH�kmJ��U��&Uhhղ�P
 6�����L`հ
�dm5�+(mKcJPA��(R׾�`h   ��eJH�� ��  "�)JT����z�4�& 0���� <��)�$�4j~��P�~%*�� �     *y ԦSFz�h�b Ɂ�@�*	��D2a2i�	��	� ��M��Φe�[8[�\��^�jN"f/W(���1nZ7�Ĕ{:�Q�4���_�� ���=��(���a�����?X�TAM�*,��AAQf�K����cC���;I$���*�T\`Y$��QmÝ�K��Zr��V�PTX
�J,����Z��׉Cf�a�1	N�F�I
�Vg���
JZ��(��ҤM*im�	�]ԫ�y��1JvnƔ����F�̼�nd��W��mo���-I�X�`֨ �-���EJA�F�����s&�ͺxVd�,�V+D�Xі��u{s>�y���2rV'��Ք����5y�Hb;��ˡ�[2+�vMq�i�F�<l"PA{�Bp��C�j�X�p�f��)��1k11r+0L���يKՕn��A���`ᙑV��[�Z�N��{�)cI����XN�ѡ���;�ڱ�ֱ�Y�a+��E�����%?�u��T4�U�lm�ن����,*�ʃkR9���+m�i�m�c��K�Qw���CM7{M$�����ZL�F�ڗ��������[i�����蚾�S�V���K$۠	��E��Wg��5тYJ���k���ɦ�F�"�쭖�U�nc"���,����1<iߥ�iH�T�L]�7e�aveb�m��Y23Y�&O�"b�Kke,�,�m�2�٫y�r�ǔ�+�f��t-��?�Z���j���@����R�[>�ܬ��[� �̭ʹR:Ǵ�l�#����34]���;O-d��P'� o5"�Rp�]*�@]] �4`�.�kr7t�Z����V�TpڥV�5��.�S73�i�V�' ��u���M8w�̄�/2�e��)�#�RV3�����9
8hZy5�w�#���y7�#u�k�z�3����Vu�F��nc�ZX�\�6��JE��ト�l�=��z�'��vim�k�O"M��yw@&ݿ�3�B+#��DإW�����6-H�ԖS����p`�UA�&��12���ekV�lm	�n��Vmv�f�{E�˥v1�2���`��V�7Q�NGR�S�����ͨ ������	�.�ښr������0�!��T�*S�2[���ahe*V�*+J�em
<�dsSh�\P)g���Z��-e��J��Z�7q�N�ۘN"�R(�>���\�:��Wu&��6�eX��o ��UJ7WR��N\#2nSGj+���ۚ�Tm��є��Q��n/pM�ZD�h]9�ʺT+�Y;Q�{[ 	�[g\Қ�ܗ���ݼ�V���*Ⱥ����KU�h�W�fn]t�j�2�bZ������W���v�] [X�NAYA�M�E,}D�;G)
�Vo0+oT.��J`U��7u얷#9�t��0ف�g;�1h��V`��N�L��䣲��`F�K
��zUf�˄�	#,�l�@p��׊�Y0��v��ef��&kô�	�%*�
4�I�ɯ
Ҧ��Y�d�ة�I V�����`��bU�;��M6��C�Ԏ 4f^Y/U���q�t����MfG3j�z��E�ti�꧸�]�8voM��X�-�G]�wJ��K�N��[K6�k��.�m��z] ���6�6��x��������b��6���ͧ,v�(��aT�W��8U7�j[���Y�yW�R�y�q�hh$^��j���YsG
Q�k���ec��j�y���:f�+���Z6i�H��຺Ko�+���Q����wbX`V�N�9df�mlIa.�WE
�ytowI���.K�Z3��Z�ӎ�+d�k�r�h�W��agrÏi�I���)s)��ܦ�	Ӻ�&f24;�E�4ʐJ bS�O,Ѡּ;xb� Ose�Ff7%� l������H�H�YU�Zty���2�#����w�(�cˏص+%�2��&�[�"RA���2ӗKN�G>�Z%M"�nXm
�V�ˣ��uz�� pmh��U�A<t>'V��6�$EJS���������7��،Y`�ޣE��Rϱ��b?\ڋ-�+e�H,B�f*ص�f�O�d!\�GE��0mڤe%5����ӬA�3B*D*�i�&nH����-v��o�P}�2Ξת��vCI��2�p{�hurZ��Zs3���JV��=�*�Lì�+ �&XJ�,֍�`5��u�a�(�X�Q�Wڷ��7r���:��s�K�{����4�巅�t��[���f��H�hM��Le�A�2�{�ΊA0kB�M��+��˳��H�n�J�{��DZU`�Q�nذ6�<f���t6a�4'VQ�� X7l&�j��wV�oa�W�EYy�t�<L=�m��ń�-+� �aA��ڥ��TXQ˟5�f�a�X�
v�-u�X�G7Ar�^�Ÿ�B����ה���YW1��8����Q�����r�V0^�A��xo59+Y�̠��m�W.��F�(�@Ar�O���;�i,{IeՉ0�ۚ�U�F�qd�wR��̥Ci����i�I:j,��n��1�xc�1y���wr�R!#��-3��7*mܧw�u�ZZ`=;���Ϭb��Py��V�%��e��2j��ǧ+[��*���M���7J�׹`�ꂛ�����-XXr6�=ɶhJ�7/uÖ��0c Yt�,�x�h��N��@}��sp^Ь{�����yL�GXeH-K�(ú��u�hs(�"�ݪO>�{`z���(k�z�[�W�+�ɉU�Hf#.��0t���1�wK�TzA�ɳ��&��*��m-pf��:Q�ԹeXÕR�W�,��D[�OT5#D�P&m�������R$/n��m&���K!�33P��(i�TL�/i�Z^��zo�mn}2�4��%{u���������4�3R�RK��!��ux/�\�,|
&�Cr�����͌��[e��ca�a�7���&92��WG��#n��Y�E���س�g��{\����W<EVc�kz��Ԫg=�k���l�.���j�̛p�6�Y���Ի��@�W�5�&�%;"��Sv�Z��ѡ�̥(բc�M�e�$�θe�hA�k:Z��j�ĭy�]��[ztu�*��^f��j�5���k�V�5MK{I0��z����I���E4�2�p�ڛ(c+*􅺐˫,���Y��a�	��h�ZZ���wh�9�{4
�ԍ�����0M�$�m�yh�F$vΑ[-h7B�TG�&�!c� �_�cC5��C�Mff�G�Zڵ1����Q�[C ��Z��:�x��3e��ۀ��u�[�4�K��X�����V�Yhhs[����,4��c=��V.w��L�&�Ȭi`��v�����+.�5Ym���ܽ�jLE�{XDa�ݩ�W@��cl圦M4u���4èQc4b�l��D��[��wD����r����F��/.Y$4��
Fm��H�ՙX�	dֱd������0�,��Ѭ¶��E�iwj�˭��5r�|�
ѳ48e W!G����]��-b�hЩ�wW��������vp���<jB�|��X�����d��S��r�>�9Է(�W�5�dk���9�RHd˛z� V�[u��y*Zܿ���:�``U��{���ԴX�F�^Q�V��i�D�[��%ۇX��K�����-�����/He��<l^R��ћOpy��GU��&i��Q�f����L�y��l��f�m�	\VJ�t�j$�vll����w�_J�T���o��eҩ��Da�N`̨dw�Uww�,:�`6�P4��V������7�v���S8���)n�n�fyIQ�Q�%�aէ0l4&҃b�[R�ld�-������W5��F��ZOw���{��/Q6H.m:`��EfVR�(�͛`�l	�2�[փ�a�[�81�����V�uf�"�fO&�U������S�oU��f��Tʔ�b!(n�
l�cLqaת��w���O�ֶ����Xan�f
z��ueyn��t��f��4V"Jx2�I��ٛC12�KjSI���حS�S�n����O[��ښ��i���:����v��L7Y��-.ӈ�n�	&���N�D^�r�ۂ���%��E��5�e��%n����mhح�L�;nCxbWJH�Y�sic��wma$"�^��(�`�R��P�n�#�U[�'�֕�]b���Q���+��cx��9X�.Ww�Ê�!�	wJ�oj�w�I�y���(�K�Hc-;����
x
��)��0k3�� I���,mhW�
R�':^�l��>QP���Qu)�c�hw�<ɗ���N#�e�L���s� �i*¥��t��S
�J��@�ksvUyt��@k�M�ժڼ�wN�G�e4�wv=�K1��f�g��4�Z������U�N�Լ�	aђ#[Eǒ��X\��n�5<�n�妳oF��]lݬ3-e�P�1�+e�2^VvB4�n�1Mw<J�L�*����J�YX�|�&[�1��Yr��<'7sv��m�/+���-�!,GF�`��yz�Y�N�t�gv�\
ǌ�,n�#�<p�2��8�5�&K2��e4G�w��ͽ$d��^�m ��u��4��
7���݊	&�.KN��h�[��ᣇט*�e�C,��C,GC7
Ŭ�ݡV���m��������`Y%��j�,���0��Kzs.�	�Ĭjn��6�Ŕ'�Q��i�͂�-�D�c*�n�b�Q��0��.����͠MM�pk�iPj�ލc`t�������Hq����añY$�G[@n�[��V�.f\��@$B7�D[�n����	�[��˛u"��r3e�dةGPD��L���4j��j=����IЅX�k@����I�o6��*�j�푆���7Q����H��H��eF]d�2�;�eMF�^[��#����i+��G-ʲ��}���]lN�x��ܷ��em8�v&eǹ�� �&�]8Y�%�Y��eҺ�V���{3�R�8ލ�N�e� N��7gV�4���˳�]Ք�8I6y�p�A��ݪ��;I�fb80�=%l`R" ��[bTEc�f�w,`��7+0���4�G'w�����`�����u,�2iB���ܩWcV�;X�c��>�q0r���d�
�Y��0�e�U����#�Q;��[؍n�hoYB��d���4�v� ��P��e�&�aW�����5g�0�9�L	Rbcf[����^He�J	ভ��fdx�]%m���e�@w��+ki=�w�RO\[���գ�v���r�����u��^&�20Ř7s��#Bw���'��4o�,�w,���N|&����gt]����`K���uoy�:oz�r�a�4�[�����F�[��/63m<7r\j���G�%0Z�hϋ�+l�wX�Ea,�B��VZv>=׈^��0^mޞ��*�wb�]ޅS2��v���dZ�([y�
V�� aA�%�Z�+Fe]���$	��RL�4�XWe�z�SH�Ρ��q�H�-��-]e'`�Ŵ�З�n��)+˱�\����J��k&Y��@�j�ˑdI��m���M=��f|�
c�э^l=���vp;Z++ZwGh�8	Yu�Su��(`��i��V��Ы������[�-�$ƣ�m�7+kf6����j��SF�5��o�t�y/�%�Z�kF��-'o%�U�֚t�X굔���qvYt(�h����!U�Yg^���z�ڱw���&I�3:�Z� ڛcE�2��k)�(��p��R�$�z]�$-ӓu�l^孶W0|���
�dpOw(�4���̭ln
i^2�Z-,��a�4BJ�U����l�&,��E��Il�(\wvL����*��U�N�a�hnTʕ�1x���4���@dS��ŗ	��&�wyghew	��i��z��,��Fެ��V��xok~�{M'3e��(�[MdwY-���a�ș��r�n�� ͧ�Q��n����=���N���,�є�i:�{L�c��RhU��J��k���,\�ާ�2bAe��+Ї���b�˻�j����������%��i�}��6�Vlۦ�B%72�ゝ�z-n��,�7I�̘�ұ��� Vfe\��2<�u�54����F�X�/)u�4˧E^�`aq*tJN�j�,Y�rkB�7�У�<�I�Y�s9U��~�`�u�M��V����e��5�*�]#v��Ѹ1�ؔ�y��@n8���5�¾G�FkCS��̓a����n������ep˧�leeYկn�
�cg���`�`�+&\�Ĭ�v�ۻw+q��^툱ūvɇ �"����0����>vZ��Zwwb���`koF"�L�e�Q�{�k0�b��M��=H�Uݘm��{l��$��i��+x#(����XF���,���;3}D��zi�WZ��x���<-�%�!lX+r���|�Cy�]=L�@+`0�ԩT�݈/1P �V�o;9fC\�;L�W9��u�3S��f������:x�4�V��qY-���� ��v�$&���7b�QѶ�Q�o�&���l�r:��I9�"��LT,�d܇���T��7M\<���{�&�0c9�(���`�
ɵ���]l *m0Ѭ��Fk[zeX;M���Y#�tK����;ܙ�f컘� {�pCZ��e��ȫM7�S;�>����͐S�1Q����У�X�c�$��݋n��p�.�ɹ ڕ�*�Av�(��� #Cs74e=V��^e ��%��E"�M;؉�1���L�y��Sö����K�	�0m6E�RR5H+�2��ƪZ��-��]x⣗�\:�nR�3%�o������e���ɱ��vE����#et}2�;�baW+�ܥ@B�G�UϺ�OoT{7�gl�R�:�X�]C�iJ�=r��t0a�J}D��ݝ���~�����4ү�*���[����4'��T11<��g���Y�Ni�:0S���l,�K <��^Pیn�p<��fW8�X��\겞է�Yۄ��}�o��XY�J_Lҕ��9+�ig��k��j��t!���3ږ`�݋+x��N�3��̙>��eA�S��5�O�юu��x��^\�xC�����T��fށ��(�䂁���l�
]��5���B��N��P�_lf�i��u�{���R�)�"V�v����9|�:�;i��jг�F�����o�וKws�S
Q'�TL��^�&V�Ʋa%�n�I��%X��u�2�"���_]Ig����B���tɳ�x�\eD�ݛ:�:Ae�O�������YP֞Gb�0&�fTc
A��gb��p�V��$ �s�EH9K&�xU��<4T���V���k*U�SQvq�*٧K������]9��$�F�T�B
$^��L�d���1�ESB�k���]*g��ÙgY�ѝE�zXۗ���[31ҼI5N��ʼ��v�,��75�sڛ�����Sz�r��������)	N9�@�c| ,o'�$��/�e��Q��\����U�>�y|M�w��v���,�$�i��r�r���tZ�#M�4o-�w��)2w���W9�[8ů��Vh��zڳ����^T���G4�<X�a��&7cJ�3nپ*��Lb��6�p�Q�x�#R+��U�9����������}�n�d�쭐gl\�l_g`��I�w�U���{�� |t�J�98\����Р�Ǎ��]͐\V!F����]�*z�Y+L�	V��eFNеVc�S�o2
��۷�u�	񎒙V0N�����wϻ��I��htQ�!��Ӧɒpk/�[�ٗK'5(ʑ1�_)��3�tu�ϡ=�a`��AQ(��FV=����vRs���,0Y�m�vn�@�����	�u$յQ��pV�Ӯؔ��%�yx2�R\�4SY�q��N��1EK! �2K��١K��M|�� �ag-�̩��<Mgd�4����Stj��*+o뽄���L�+4;,�he���ƨ��6�hN���}Z-黽�RT�1q�J˓l�ԡ�X�f�(�6���1d��ɉU�j�E;wT�-�PXy�T�y[j�8��Cr�,vLf\���+�a��o{�y������*�1t�m�<0���Y�gF�8�1Ww[E0&n}�f3X:�X��*u1�M:��d�(Ɨ��{Y��)�{]��8�X���3�w=���-�z�K��8�pA3WL��]�9�5�n�Ui��rE�(�Y �x��u8��8s��)�&�m��[ͻ��ʂ���T���ЋsE�F<b�J�t	�H7�U���;�"���:x��`��6�nU��<��t�˖˖���G����{Gk�TGHu�ԓ"��ڼ� ^ν�49�-�����Y#V�G�*;����"ܧ���c�&���ku*ss���y��`��e$���B�ܹ�KxZ����6X��.��n-�ˏ2S�����Bf�RZE^q�Z!�.e�ڂ��}D��<�W]a�i��8ȩ��cB�3�A��W-Z��4(�U�Ue����֮5c�p��,6�I���
���ĳ���������K����u%��@)8�eS�n����n������ۄa�s�����E��eh��	�����p*�HJ�b���Vv�����-�b��V[�z�k��z�WqϯBB��G7��\�ItP*�\����r�f���f�G���'�_n��t �N]����	��L�תP��!���f]n�˅��\2���Z0�;�`۰�\�\���[̣w��!�X����v�U+�7�e@�oYXQDv�W��]�.�&\��i[�����Ş�)��5e�.���k���,{Z�<��PxSZ����5�����~�wk.Yi��8:�ν�<����,��c*7�$B����r)��r�Y����%b��q�fF+:\���n�{���[�=����3��]㋳aX����f��%����������c�	8�Wus�����7[i悦�e���k�V����r�9�!O.=��[���@�3N�ٲ���S̫��N���+$�u���M݂���7�퉓XWI3b�g@�Q-/27����d�8�9X�	���5oZ�\� [�u%HQ���o:�lO)J�����"�5�mI�zq'S��:�*��wX"�8�q�����@_�O`V�%[6q�5�ݤWm��)�����2���9c�� �M�Rq��/��hqYL���]:�.v/�Sm�؍�*�p�Ȭ��(������B�����f�ܮ������[+6�H:��,$퓢]^}��:�4��j��>mr��$�8���#f���0�m�ZGs�3�;D�]X=�(������J����A���;G0ib�nj��|/o�o`�u����`6Ӗ�;�Wf\;6����P7N�ccY�\\8�N������Zk�5�5i�o �Ω�oY묀�x7�c$�6�����%�,�Cd+��,�gSo7
\��@T��=�*Jɲ�:n�a�&����JQ�vqd*�gS��2�n�ӵ� �:G�"��V���Н2�޸�l�v�:Ϊ'mf�g��y��E�B����x.��y�t��ͳM��u�b`��Zh�<���V�F�N���ڤjd�C�$�!P,��Ǚ�TG2,Rj��W8t8����{'�E޺��vnZ�j��}�"x��>�ƃ8l��/��gml ]��
98�u����e�3�ޝm�6�ᅙ���5��m4�zWdR�#P<
။��e�d��׶��սn�!�u��kk�����M��~Zxj�Bq��1�t�3&�|e�D����m��9�9{6.�g�Ʀ��y�L�Ǩf�{�9�Ҙ�T�}���Ԥ���bΊh�˝Zp�d�#N^Pv
iY�iӖWB`u:���n�Bnۑ��}]/4�����WJܙ�.N����Zh!��^k�0�؁4hւ���[�r�Y&#��wϦ�si	���WZyyR�.��S$������z����ed9�ӝ(�,w��@+��e��`n����7g��dw���ig|`�����u��ܼ���^�a�S���������\�hfWd�GyK�'�"��W$�>orz�v�1wV�Y׸(ލr����<����nun`�����^\�_? �׉�y�dN q�p90�SN
��6��D�/�����	ϊж�^�%K�(Ρ�����*��,�(���y���aL]:��D®���*�[�$�-�.�>�@¶at�8�1�dY�N�9:�M�hˤ�M�%��$�M�7�|o�sw��zi��=���S/Ep�e�D���B.�mc���y[����ڂ!\�u�f,��_h�U��͆w��L�(����U�F�fWn����F��V��8i��%��=[
̻A��;�����=w��]јF�p�a�խu�`��ag-��c�7����7�2�Nh��v}�wj�J��������0kk�j���9b��^�v�g�7[�vvk2���3��j�uKE��*)D���Zl�p�#�.�T{��7w 
�C"3�ވF[k���9���ڗ�yZx�H;�5����Қ�P?i�a	��Ղ�eI�9������&�cLܺYن�v�w/#�݇�(�emֱ%g^�Gh��m6��ag+�KM<�
�@F8&hͮ�A��%Z{@v�E��9�v�
s�MKv�n{t)f�޽�h-
��#a���+��*@S��\E�5p�k���籚{K}������Q��$�FA�/�R�4���b��P�vo~S�,r��eݷS��M���7�qR�A��7��3���p�5�0��}��p#uU���Nޘ��r�P���h�ve��o�����JȸQ���X��P{FɆu*���p���d��hW	3���}PQF�>�!�]���K��r*Z���5�kQnr��0Vk���>����4o>5.��q39���5|!���*��ViPyf�v).�D��<���}��]�s��͗�9�#Z�c)�TQك�c;f)a�
�ѽ����"�+NS�}��Y�'u��+̥��X��d݀K�k�!�k(���aծʩIS��ݻ�4R߻����J*{3�6���5�#b����{Y'�:У����<�n�)w%��S&G�N���]a_a�4e��������Kgd���^dq��|9�W��5ɇR�!Çx5�Z��+Y����5VM�Vr�fwE��dJ��r{�W\I�PW�z�HC�Sg�M�:7:�������9A]
����p����y�[{��x7ؐ-)�kX�p A[[z��\]�N��3�6�v�F�2�:�X�ɱ����x�)v8��4@�-�hL��S{�SK�1"o^�ɶYS`�{K�t���`S�N�۫�:�Ŵr^NK!�;w�����2�����+�m'����u��0:�2�by�ǽٟ,�<Ir��=]�H�'�l������Q��Qb5S#=u���^�*�mm�V�mv�ɩ�w]j1�Xv��W ��H�m98Ǻ.�Y�r�3vy�m�ózZx�uv��"@>�<��4��	�d#���9|������ή�.tC��5��/�`�lm���klsǼ6�gFKoja���םB`9���x��:�N��IR�g�v��:�r
c4�
եݛ3;	�II�V�	A}�Zi�}��x�d���/�1us[���KqD�7�	�ЫƯ���j��}���*7��툪S9W�VQ�xVLx2�L�5��!�s�7ss)������Gb����qԭX�ݻ��-�sq�n��GM]Z69F���+��nb�\�(�QW*�?��ڗg^B��Lc���fY��x�G�ҝv,�����_)����1"P��2��d�qbn���k��G1����4��b�wc�ڦVt�YG"�*���UXH�'Ed��v�em�H\���s�*[J��h�Qf��
u���7��S����trwj��� �]��&�{9\�te�.h:Ck!��6�WY�6�� �� @Ys�&+_�]E�q���e��n�"�4���yt��Z�����e7Qw�l��.��L9�Z�$t�/|�_<�����=ՆsƩ\)nZ/$�Z��X����}J��h�7c���/r�W	YBk�
g:��U��M; �;/�IY����e̠r��-�j����S��%�9n�\���c���Ѵ�rL�U�г�٧GFR=�b� ��6�J��lB�ZTv����� ��,@��(���:pj�)���ǅ2s�����hY�}]6\�Ѫ�v��:�+����v��堓����+��g��fh�v���[�V���o��ut��d�H�*��ro��ײ���ɥ�10ݘ�;FZ���b�^dlfB'�։$�g��}]�nWV��V �K�!�c��Ow3���B��4:�kTM�y���+/!�z�0��O.�$�Ù�v�ҹO�:D��;�e��۹Y����=m��Z�O�l��E��ɀ)���N����ތ㻹���Q<��N�;,3uk��0�����/@LcD#�Q�m=r�l3z�J��� +&\6L<�"�����<49Η��\/;��@�ͳ]�m�ngm;]�fJ��S�-P����c\�^ed���Ժ�RI��U�=�u�t[+��澥�V�p��ƸY����u'[��:�,�9Z[���<;�I'f�8U^�"��G����}��������sQ�fi�;+��L��z�eK�֒�x5�Z�j<
�X��X�i�\EDӗ���Ax����t@'C��.�V���6�3�7N�=�}��[wl�)�A44oǉkBm!$�7�d5���y���$n�����S�f���*,�B�Sˣ����%��n�w��u�G2i6U=�n�:{N��K*p���N!�k%�q_:x��ِ=z��'X}��I�xi`E P�n�^��:��V��d��&��6P
E�2bB�J�t�`9��
,�q�-!�����E�p�%�����Y�_�)w-�$�MK��%�r^N9��� ��������y��*�]�*3pʌF��p��+�C�Yr-�j%��e�]=0ɔ�J�*ֆ:%:م�c՚��-�2�$-�D�\� N��k��Ӵ��VL�{r8��R�;�f���}[�3r+��.�&t68G��S�iN���8�u7�>��t:��(��/�����-o<�o�A�%�����ź*�9]��3%^6\���@ov�>sxME��޼�}8m�p�R�C�&�Ѡ�j9���$%ں�M�Ճ;r12����^�h����٥���HJy3�w+���c��g[�����9�xͳ�Cl$sݡfY�ǡ�
����q<z��U���PQW��.j�ՍdS�K��wf,�1�C���2=�\�gv�Ww���Z���Z;n��̶˘�.�j�.��Z�A�/X�ή����-,q�/K�	c\0��ws�dV0%����QE���<j ���lf
W�.LE�L��	�T���儢�q�B����"�Ȉ]un(��.�{q���s�_�j���阌�\�VpW�`ޡ&�<�uwH {Rʝ�V�ê[2*p�y|q_8��_�b�L��a�3I�a�F��1������79���{.��RdF�wX��o��GSt���0>Z�VnA&�֥v��|F]6l�#&P�B�']�\�]]��U�f��W⢚�U�Sr�(�����cD�k���Yb��{o��R�;He�ZTe����PU��DZ�vݚ��G�MV��գ �R�	��&54r��fw��vVږ���ԭ�h܈�kV�?N�Ӭ�jv����]Je�`�
�ι݃s�*&ȾL\���r8��<l7����7�w'�����WU����ΥN�;�Č�c�I�]6g*�Eo(:P��圑�1Q�c+a�3�}[c 8v����]kQ+��ŌmkޛE��N�!H�]Xcř��7}S]q)u2�I[�6��H�5,�ݡ��Ԧ�Z�s����;^��hvs�l��S$��"i���6(���2����x1�H_�@AH��3f�c��\\%]XT��f��u��FأF��XV'���.�,+cn̓a�[,���WJc����p9R��Z�]�R̥�����6,N��2��ڷ� h��XCtD�G�Xc����ޫ���'�x�\�N���4;�5nNd2�i�{�L�0)�o�����gi��涔d�˘��GS$�7n���,�1,�Ur��t���(���%Y��(�3�e{}�N�����J�@�Ml��6�򮊟Q�.)W�ڴo+���HF��Gm�4���W9�5��ڮ�n4�b!C��!�)v�ק6%�5�.�����F�+��#[���+v�VT��2������N�U\���C͜�m���khţe�a�fao&*Ky�=�X���}yB�څ�����*}���wN�N�_�Z����'��}A��,�������htƺin]ֵ�Y�A)O�a�s9��)��՚���H��t��U�ܥ��L�
ܷS��,�����-�TA����+v�<��W�96��&�]�K`*���{�.������m�Ul��eYu�iN�h<\գh�Ιj�/2�)V���l�v��o�]\�:X���[.������s�u�ͨ$wtvh��x�т�¶�U��-ۤ�#��B�>�ܬ�yL�S'9�5�*�u%�����	*6�۾ㆲ���7LI��tL��		�Hq�<Z�t%�l��ć�W�8r�/�/x�`C�j�,���i[��5XiM?�.�ܾu2em�P�jf˼�]���X�E�W;/�vG��48t�e��U��wיo�`Uc�&���kW���e�r�DM�`!�(V��,��gb=n�:�k��Y���b!+�L���t����iR<��@CN��Yo'��	�7ZWY�]�_e���{�9P��0�oM����Z��8c��3(��|�F���(i7��՝ƓJ��]S�h\����%��won�rf8-�=9k;J��:�^B�luFSFj��zwa��֮�!K���= �죳nǯi�v�4G�sU	Ɍ�f��x�il�9v1�ƯkS��v�%���g7���S7�����P��A#^rQ�S�=kmnc�ыl�XW�o�x9��>�S����/�reL��j9v��.���T�|����˔���^b�d�I�`��\�w�`��=�ٔ�tUuL�E�F��q�fvwe�Av
Җ�Z�3:Pa��o��z��t���]�^ͱ�<�0l$Ͱgu�#@g3���A�O`���߳zN�,�|�6eۖ9�:���xT$�v�B�1�ܸ���h0�h�8du�]���閳�;�%���q��Oe�([���(iD�H/�g:)��^�<0X��y��-I	��+<%Pq�Pf�ք#.��E�D�l��]��:L��I�Λ�p'y�Ž�H�������澰���LΆѣ���r;K��$�]�@�V|�(�M����{��g�F���{��b��|�[q��P4_2[�0��ب�:�c&�x�h@{�E�E�T+O:X�f����s��eY\�;}����o����u�����aY�*u�a�ۮ�c/��V!bU��~��w,f��Jơq�u�j�����[J
�;U�j�-X�6�h��.]�Ņ�7��Wk�E�5!�����G�]�Y����-m��V��\`��ΫR����7��w9p�j������� �B�L�3��ou3��'P9���WN�fk�F�[Y��Ѯ�eY; k��rz��c2,���,u����3.���p�,��J�2�2�ᱴS���e�s�H�L7�x��
�g�0o����#���:�X��A��6H��F`�bpm�efK����
���R#G	��>��ch��@Kb|5�=#ԑ���R�
 ���ld$��J��iH݊�Y�5��1`�&wNf�'`;��JW�n�����N7����Fb�p4�<4gM�O,�6jjy��_a/5��F�;n
:�v�Խ��z��m�㕱���	�p��KZ�pŔ��1Ȟʽ;��;VnK��/��']\��&�sBw=��MT�	s���p��+���3�0�_���l��qN�E� �ܨ�+3;\䆮2���a0kW�Zifc(�4[��o�0 ��jn��1��˝��D�t�W��bqܩ����̳FE��?(��l:��
z�7����3��\�qΛM�:x�˶�+�V��_+��>k�O���-Yßq�7V��#�����)#��c�.�6�s���EL,ޙ�55Ava���dWM�ts�Z�o0��^^�����cS�=�Ձ�6���\��뼇�/�"�u�zs���te�l�[{ڡŅ���}aV3h��E��b�ݣ7Gw�ۡVqf�����{'�f�h��~l�{�i���>Q�<ael����M
5�oR���n]�G/��p��ɑ�������dת�V��U�u�@��k���D�-�L�O3]iZh�l[��z	8e����q�9�hVM�Ro��7G1�ȥ�qHr�8��sL]��R��
�јxӘ�r��'^���	�Wp�V�==e�}ǡu�X'�s��ud�����[�I�B@�/�#�WZ��T:H�i\9�q���b�x�j6��c�*�z�*�N��O��3��p��YDm]\�������$�J�<,N���C֫ù�q�.��7��|�0є ^y�Q�v]�u��(+��f1}A���렱��o�SL���Ϯ���LIb����(pspH�m8hR��:��R/��S 8��+:�gts�@.a��m��͟��l��w��F���6�.�qM���p�7]��	蔋��<�\�������㓁��j�<�d�hB���v�96t�"��l(RN�ku+镐dc�����%�֦H��^�Z��E�T�]"�oɗ��۹D�O�̣�ѽ�r�/���)�p� �-�T8�O,fN��b/$�H�#�m+]��
��D��&Lm��J"�Ӽ��5�Ac�LU�V��Ij�9�����4B͙Lq]]x,rwV�Q���Ӹ��,�%���
�Y����ȊԦ����Ů�#�# W)��*.����t>Mc'�֍$��7�\�d�F��*�u�Y���L�jD5��.�B�z��ʅ-�RW��K�v����c�J0�����eı��'�s�-�d}0}��gh�+b{�c��"�OD�e*���0�R*J>MN�Y�)���"�ϰ�=�%f��e���i��g�;�j c�N7�e���A�n9"�!sdY��E/�V��Ff�x�_@��Z�T��Z�V��62��s'|(�/&�Jwg�Z��y	����$�u�΋y�r��O���Y��7�P�ӓㆬu�cz,U��R�f���Z��ĪZ��LL,�]�<���u�p�����#��}5�Ҭrtft3B����������:�xQg:��VP%nC�R�{�`�=ux���V�H<e��!زPXt��Pk5�Mk��r��zF]����*u}v5���EY�W�YM�����Z�03�m�S.#��� jV�&�4�BЂ�P�Y�4���\���`xd�Oe�Z�D:����cY*h�4��(u.t���-=���ܜ[x���,0U�y7FZı��n�gJ�'�,2.SWԁ�U�����e���NKd��|�xkVث�2+��=�Z0
׶�
=)�!��G�ڐ�4j�̘�}�R�΋F�������;���rN7T��u�[���$�c36�帙ٓ�� �l%��/���B���&W<����@��xK.�=b�x٥����v� fp��BW�T9�[�v��M 8�' Nf��7y�WlG�Y&������=��l&sa��R� �� w��o=��=�L�2��f�u ��yT�@>�P֨m$�g\[| ����&����w�uA��N�*s�@��ڗ ��;�V�v��w�:j�fd��x�s����n��i��(;��,��:R�}��47(��йz�z�yƲ�SS2���d����G�+�#��+z�������{)�ۨ�-������ʲ�j�:W�  �I�cǕ�-b�4��[�]�*��{7	�=Ei
lҘ[�0�;]��ðb�ۻxz7Sj�16]���jl�*��ca]�(���3&�j7t�a�=��
J��gA�i���7{���d�y�K�ǥNբ��(N�݁hb��e�:B��E�/l�K��uJ��7Zp*I�:���*,��I���i����5��cA�Wv��d�%�)@V
�&�ˋN�r���Έ� ;p�`��d����k5�#���ڔf�z�ٴ�4�����q�_�����+kPo{�Ƙ.�*�,PΏ�{p -��n���:`��L�o7H7N��S����k��$p�6R�A�/7!��.����F�(sj꒚쀐g(����G֬T]d܅��'#Y.�zջ�*m�laӷ��F�%b�[�dt�覌"V��۷%����&�����Y���#��K\5/1��*��f��M��b��o����a�5�`inK!��R[�{\���"�-�·�owchGAAc]E��.���t�\�cRv�{{�+�[�.��+�tvn��t�B��K��<�i<��OC�r�%C���/pc�^T�������6����9V7�E���8�OOL�	gr����W�IZ�rk�
��5��7�Rw��'�X"��]�<�{�mH]��j��Q�6.Y�F�)��.���<���]�t�ICGʮ�O���E�N��hx(^�j7���u̩`�'MNi���i�r�o���U�J��pgw7�������H�C�Y3+Nau̘���2ow2^�ޝ�l���g*�2��Y�_R5�jԞ����67)a�����J1uj��h�D��e�ܫ���q���*d����i5��n���uŹm�u�xY\f�S̩ۨƱ�]�ݩɬ#��͒�V�����Wh���r<�cXmzs6�9�ͮ����q�&QL�m�Z�v�]������w`M��č�����,<XQL<Ʈ��_ �÷ RuZ#�˫��+��]4qA�b�Mp����Z�7��.&ʜ4+%�����/fq�甡Lt��"D�|�ø�_|7����x���h]�W�(������nҮ���;��g$H�3�����N�a��d^�Z˃b�8�R���*$�h�,L��e�ͷ��e�N��|�6�>Vi�m#��f�9\]�8��v�S.�;�Zz� <.��X��L��\+ie��PQG�u����I�jSo���Y8����<�HfAq���m�&��̖��=��R�������{q����LO�UԄ�ެI�`<u��2�i��Wg�:�Gz]Gum̩Z�a�҃����y{}e		ʄ�ێ�`-�%�:͌T0��4�d}����kfbn���l0��Y�y�q���Ä�8��<�yImkn�橨Pޚ���7.��4��+n�q���^Z�"ʳR�>��7w��C:�pǜe�V'#h ��[�SČ8T���e���]�YV���y�k�"�m[�1���Nnr���mgmm�x���f�k�f_(�Q���;%X|3]�8B���B���U�2-�WK�FҶ�=�ȳ{�\^�kS�;���lɁ�֐۾\����7o`5Ǧ�9��k8�9�In
�,�kiZ��%��^<�QX�*�R]��/��׈@	�o6�W�F�ɃW^,	�rq*�ȹg��b��M��F��5�s����\���-�x���|F����T�G�����o3KyWӑMi�Y��)�n�xp`C���ӌ*�[j.�����Z�e1Bx������g4u�;�p�ܫ���t1���tGq�����zK��wpù{y|���GX-�ݷ�h��L"a5"u��gU���Y�U`b�X��ԗ��0F�R�d�����;=�GWl�vV�+�����{J�mt.�������	5f��Ŝʸ��ٳ �0��U���<[�b��O{1�+zV�k�x�=o&јsN��ʟiաt�<�-��b���b�ΆX�P���{�K���Q�Z�\�n�'��d�<y�{�7��m��|O���d_�@�CH���?YG�8>��q��o����Dv�NP��s�ow�r���KU ��WFi���/-X���e*�E�G��=Uq���S/i��T�D0�c疴X�z5�Һ�������E��QB�G��f��*�^9I:���+8Q�+J`ʊ��p��Ԟ�2�ދ@���R��PX�r=�XQ鵻�jřC��cy�	�nW	�G d����Xk��+����j���I+$,�p:i��8�#l��w�T��e�vp�+X�����85���h��M]c���4�V^>y�]��]��<�Wm��\��Pv܁�K�j�B�����hǶ�#�eM��ڲ��s����W��^B�'X	q:v��Q�O,��g�q��Q�]G�R�gEr�z�=Y�{]ު��hV\��r��Rr�V�zB�F����a��v��Z��VPR���/F>p-�3	U}�۹���NxS5����#�q D�
{�y�yI֢�*����5�b3����mΥ+����hiJXr�|1ކqd�d��\d������ֻG^o8�<����Zd���GI//���g�ڼ��)	L�Q׵���X;AXR��%:�.��Ӄ���Yk��t�����ȶ��\�f�4�����K��O���B#)��ّ�@$��|�)�-�
�T��~���Ե���U�]L�L�Z!��+S4L�PUR��\����D�3���3��Vڢ�TR���0�m#h"
Tٴf�Da�b#s�k¥xL��ڈQ��ˬ�mV�ҥ��֢#m(��DB�!��4�Z�l���5E�U��є��V�+Z�Qb�Z-r�m�e�VZLb�m�k�֙���q����k�v[f�ȌjUZ��eθb�l���ihl����]�7�j�A�SE�h��,U��V��ĺ���U��;h��eu�m����ҫm3��L�"&�d�Z�DID(֢�neu���jZZ	��e���+Z��[TZ�F�m[3��ئE���4V�l�E5*�J�Ѷ)(���@��[J"�jQ�6�ҥ�9�ؙɵ���J�TU��.�D��Db���R�r�5*��[j(���,+Qcm�Kl��08+Zȫ)J�ֱ,�u�m*�J�m�`���A4E$P����-��E��+�6pCj��ݘ�Nm�
hmʽ:��fҊ�uC@(�;X3& �X���C�i�S��kĜ/難Q�gh���k��y�m�ks��ٍ�\��z�`!l{��FEOi�ȡ�~�KT��{!H,\��n�4�|��V���&J0c�E�u2G��vˍ���a�]<��Nh���� ��V�j���{>FBiXh���9N��$��8 �I㮍M�����aDtȵ�N�������`�E�z�A����.`���XO�9mlv�<\��1N$w�d���I�,��r]��VC���gzڶd��}9}o�-d�^5Jv�F�;gǢ����"�����$+�o:�E�q�Rě��R����6�2��ڜ$�H�/�rQ ex�R��>���7��)f7ڢ��ᓰ��D�p��d��C�3P{�O���`#��?<�.5�߰j�/^X9���V�A3�>�5�49Jq�r�mD�. Y<�ah�5�`b)tFi����۹��:%���/ْ2���KJ]E�|��] �5�9 ���-���7�H�jlJ4@}znsWIh���x����Z�H����\A�뒸@�@r�~d\�ݕ�:���[�S��gzo3P=�.�d	�Ա�*� �<J���ޚ���k� ܜ�<�:U]�8w���� ��$��wc�VH����i�.tH�y^SI��ͼ'q�{���Z�uy;����d
�!�+�1�[��.:�+7�Ox��������L]A,yyd迷���S���4���º,s�E�Ӟ<�$G�0+_XJ�iֲ��{�L!�O�쉴o�smZQ����ڲͽ�ّc�d�V�=b��;���W�#��I��΋{7:���G%|�����u����+���&��+}"�/���UVo���k:�511fT6���|�x��'Mźt����tXnYhLtD&ƚ�#/5�vuq�l���7V��I�(pK&������y��eMR/<�V�g+�Fj��Q��ݾ��k� �|X3��rfY�^�R�;�K��I���h�RCďD㳧׉hz׫d����$h2#��s�`�a�#���6%��.�IWx�y��Gs+b��k��R�nv!�rI!L�)�k����b�������`%R��w����Y�P>-�[Z�
�
ך�,������gO�yg-u�w���sN��6+p͝��J�X�:V���gI���N��ϟ��Y�VG�z`�o�iG#�p� �5��Ʀ����M�͖��0D��}��mF����#��!����2-;v&ľ�"�:��[�O^��8q�~���ve��ĝP�F���o:e"�q؇6�:�z�� s���
f
X�v�w-IDs���y�](�%�;�p�^�uɠq&��*q8Z�v�֐m�s6�E�h� "ؤ�9�O��R��B!��D+��B+�*��P����z�g��"v[C���{q�Yy��'ܬ�`��(.��]��
�Pg[�'�.��3b�w0��ukS9$�<�#�Jɧ�"�P�f8F�98c���R,�8y�V8�y�-7�ۨuR�f�3#z!�����n(�X�q�@Dxda�1n5����C�wjc�M,�F������i�`.uF'4E �V8�v=J."����\w�荽i�UZ[���#�4�èގ�l�db��WL�r3ʪ���Q�M�/����<b�DZ�Y3���k��3.X��"���הt��
�\���ջ���<ϴ�+��]��\MV����Sd�f��,����(�[��c��}�q|)�9��\�����z����AU��5�x��f [��`v�7����%�� �o�]>�b�M�2�tE��o��y���!�PLm��`(Nۨ�I+��x]��SŽ����Q�n��=����]!TĽ���GVL�h_B���[מ3:{�	������v�b��Ա���O��Ui�@�"�wM�
��&M�'*�{�s܎(}�Tp�O��eN��1�AP�L�3���^�T$�U�T�]���s��O����s��warH��#۵ܝ�!�JZ"F�gL`��S��v��f=� G0S�hGuq����5�rȊ�솬L(N�w�.�t�W9m�}�A��'�"F����'�<�r���<�(�	ݳ�+E�eՋ����N6�d2lT�&!��M��\�
��0��&^���M�zo�tn:��R�z�^,���Q�g��do�M��P:_�n?�wp�W�u՞�7
up��g�yu^r��gq��I�Ҋ�Ldj�⺼�P�ٳS��.��2��⭩���]/�n��WBo��[P�e%5DןuNE�3������4��0%�� =��>���qޑBb+Q�;��t�H_1�;t=��GfR@������T��R���J>e�yH^�ޜ�zd<�MI�v;�KH��\��ݪ�.Q�B��^M�%py���3�J�f����x���]d��N�ޜB2Ie����%���e�`oH}ֱL�{4���Ct,��qJ��yԯ�:�;��ҝ�AvH�Ί��@n[��磇$��o*|��Io:�٘z!�A��w�&m���d����A82#�QS9Q� ���&�i�����7^m��}X�ٛm�c.-O,մ�q{��y|_d��
r!�Q'H��(�#A~�6n�	�9^�SI���y��Į���!s���	��Og�#�#O���h״��4'�g�x����6qobא�GP42|�v���?{+N9��˴��A�5�yh�&��b�_�}����؂4��o��"H��s<5QP��ϑ�J���FPj#cz:"	��Ot������io �	`�d
��X��r���uG8g9����B��HdRt��(�p���m%��+��pA�`h�`q&a�8���ӖGV9��9���R-���,�;O��v�hɃ�_�s�����"c��2��	k:�U��Qе��W7kA4*�����ܨܼ�7��X���a)��9��y�K�WX�cϞ��F�
��ՙ���R:!�Cg`�8+�Ѱ9.6�2��s�� 
�&��S�gm8ӱ���TS��L��5/���eU�h�O�ͧ�ͷ�Q�1�N�p�PH\��u�w�Vl�} ���h� �r�w&H���kp�b$2v�͓���}���dX��yB؄ˡ�,��f���E�0	��Z�\W3�ĵ�q!�;�Yɣ��w/cR�#�u49Jq�ܰi�2��00�V1�20�3�nM�çݶ��`�0�Ϭ	s��#(f�ұ*w^ǔ�ר?w:���y�6)�0��i=�@�`��<{��.�d3{r��p({5��s�D��)	����M�̮'����I���K�yteÈ\c�@ݚ.U��̙o�ƫF~K�]�~�}�8�j�O������6:���>����V�-c�ʣ傝(��o�@��r�Lv�t�ǏX�<1����,�NGP[VY���Ⱦ�1�^��aƞڗQƚe�1J�w��d�F�e�F�q�T�ڎp:�w�y+
�p�8��N6E�kEՠN�}��o�\\11���Go�|��+��p��t�[�H��9�~nYH=4�߮�Ev䐉Ѷ=\8Ӷup�F�� ��m��<٣ho'�f'/,k�!h��´*W�-�ٷD���Eگ�`�J�`U �RT�f��]@jf��p=���w��9��%.���O %�iI�o��ܣ�6jot4�Cj9��Gt/�Y$�᪽҂B�?�]�3ûu:K�W��3�e	�E���˻v3:�S���GKF�(�`5�{C��G��y���Y�r^Ȯ�Bk1:�1ib��v�I���}��k�
�ù|Ue����c(W����xԱ��u����Zp��KLė��Y�*h��Qa�؆��B� l�F5�<-�(UL���v�<9��ɞ�\E�n���8B7��2-;v&U*�aB�R�$.:v��K��\��C�6ju'��!��q{�#M�0Vo+e`.G�ÛQi�����8(I�5"�L�mT�Y��,�S2 8��O����ݩ<x�49*qr��(X��]FⳞ'<T�NwW�{�ٷS����2{�J0W[���Ww8̮4�L����p\���>ת�o����}�Lt/U���Xܟ�a����C�{-WB:jB�{1�c].��]�����D�<��W{����4����X03jå�~�1P}���X�u�㰯n�yL���C�y~�-���E��C���o���{ۃn{iU����tx!UJl����x��R\s{h9��r��Q�rY;��'�)d�"�pC��^EK&�;J����w�
/�����0m�s7KrA�i����h'�;i[̇?SR�ߞ�3N8�͘*��q�B 3�Vt�D�񌬐Cm_ӷX�D�60��{ @���i(s�;��Ab��>�K>�ٝ)�\�9�l/�V���jz�*fQ
"��g�CQײ��#���/��򪦣 -E��&��#{6���g�v�{}�l�:|*
�ct�\�I�Kې�΢���s�aT���oE�>�W�����U"-E�,&���\�D!tP���LKرQ���d�f���+<ȅ��uF�5���Me=�_���v=C���xGEV|=���+A�^�*OvR����Y�����/Ip-�.ݡ�8U�cf9H=��kE'�H�aG����}����M/a��l��ށʃ=Ѯ	)�oj�srv �A)N���{�y
��m�f��u��c�94������E�gp'CM[�DT��#w.W4�(��S�i-��d(c �$�	@%qc�<�r���<��0,��:*�kV���K�4��m���w�$����ۓ�l�l�{���u͛�b�.WEM��ק5;��zu�A��	����v�N���0����w	�����ԏQ��O7A��=������Y@�[QoB��ʀ*EU�jf�j�>@9N�I��R;9�NL@�z��YC�h��꧛����Ll2�+�`a	����V!t26�rp��=�a��%�k���~���A�%^���R��t�(E��j�-�]Em<R�Dnf��6�]���o]�X,�4�I�Ҋ�Ldj�������,V,��o�����w5s��̑��l�
��ٰ�X*��()�%�L�o���1�� �[���t58eV��Li�0"�\aʋq����#��>�kX�l�J*���Q���	E�gV,�o�
���r��	��D_���e���-�qUP�|�>s���f��$���s�O#�i#3&M�����b�+�&ݙ�;�C�΀�����ڽ������i���oӳu��c�}KV[8mA�
r!Q�"��#���N��*�+�hYׇ�h�JHT����0RQ����o���cr���.Vc�5�^yG��̳3(CJ(��t$]D�P��k�'ȧa;ŇS�h���v�%3�����1�l��=������٢���E��f+�ST�BӤq���W=qH���v��z�`�@��� �VV��&������Z<���r<0�(9+
f���eJՁfml��+�\V�w�t/a�*N 3;C=�����f��6�fɭjݓ
�튉���A��A�L�6D�t��QP��|�iP|H�^��F�ʻ��:%|V�z�����j��G��P>�Q��LG���@:��3��q��E��<B�eb0��mf'.z�!�ѕ�{�$h�`q&D)�P���v �<p�6���aq2�g��qyq*���B��xJ��������eQ�t��.����3�r)�VdNvh!��m�v�܆#g3���y;v/��-���HJ<R��A:i��Ol5����]�uЕd[�Q�HFk"F�TND0�_@S��uX�)��/����(H��q=��t�T�6^\��u$P�� ��8�m��mE. Y8U��V���.�Ü��],R_#=k���7ْ2�]�XT�(ߞϔ�y9`��}�f%VN,3Yu�h�y8���U*c�Cn@��x�g���&U�pӼn���D���5�L�E,�{*z��/1`&��eћ�q
�ad�!�)���s�ܺf���#��>>�~�*�~<����U4Q9��,�1U�ZЬ;��]�6��w_,r�vVEC8�m樱<ћ?&.�-�rgN��l�dn��V�ՁL�v�<��ν�4�,�6k�2���1�BT��S�u�P!۽��R�i_@�|Os���9�����T{���_���ck�L˻���P�ph!GH;�����D���qQR$L�|]�`�ց���e�t@�6��sr�/>�sz5�9�ۈK���;�l��Hջ�=�]�N��P����E�MZ=�@m�?"7m�*	��Y��h�v�|�g���6-c�{FqwUgU�bRj����+͹���R�S�0��{��'�>�s�d�"\C���ji��E�!wj� {�aq��%b�[/��2�WB�Z㭢��w^鹘��,u���.�+@T��Y@]���	읠3%�
�.���0:�'k�nn���s��"�x*�I���}z���7���pC������9¯�S�o]�zզ�cb��Cr:�חޣ�tG��#5�g��$��:�V�Z֤i�:e3ջJF~��T�KK�:ޅ��x���ҝԽ�ka�te�gB|��'@�(*N/`���(c�h�}�V� m�3\|T���E���쫅�x�m�e��Ī*곐F�1�p�إ��:z�4��[�xs�B/G�M�n�	{Hp�p�`м5Y�k�VJ9��Ʃb6Q���J¦�t�*�<�&Vj��7֔ú��=�3�3�f�:��u����TR+���y�zj^}tt���;�v~�o6���g�x�F� 슕�r�vfM�ۋg���H�Wq\k��+9ޅIL�ҡ9eQm��FZ�g����=�W�ts��m)���}�����r���v�*sN3z���5}��.�֎t�=fM���j�պ�-YݟIвǋ[x~�6f=�W{]
S	�St���WE�Gwr�`\%�Lg<�t.t���ΣP��im��ʡl'��"faco���k���r�P=|P��η���mm��z�m�p�հ�5�Na��8��)��2r-��Z'���i�6�Pm�*��6�� ��X��U�,=�{\����\��7/�igue�H˧��K�d�qf'/�n��̱�}k+!��.�H�.�X$�3v���k�e&O���Q!u�u��є]Ʈ��Nn�K�.V:�n��\�/�M��5ي����-^�m�o�����7ƻ��N�p�޾TY��drx@@uާh��L��-��ӴU�uxo�R� *G*�ޥ�0ܶH�.T#Cj5�Z�̘�[%sޣ4ղ��-6+����|�&�y�Y�$�	U��۲�˒-)���޺Qbu���F�u0+.{��5�/"z�[�Y|ȹ�zK.XEi�N_[[O�׬�g'��0�B�KH5i��gq���W���{�g]�wX��BT�S�ɏ@��LҖ�c*R���D\�K62 ������Z�)K(6�[�ҥU�m5�k�k,�UB�Ҩ�j�m���vV�Q����J#�-�R�m�E�m��jҶ�"[+-�KB����	JZmpQX�-��4��[ZX�j#mQ�mm��J*��Z,X*e��b6��*,D�Z�X0��L�mP�CYTQ�-U����F6��R�֢��靌m��L(�(ҵ-�E-�&K�s�T��kJAKim�Xg7M�����6�f�5m.65��S;Z�mԮjVb.j��ֺ�2b�Z�+J�u+�+�eƦ֤֫6�%(փ%L]�1ef�R�J�ȋlL�e�۶�km+TV�cWc	�K�rM�Ү�5(%+V�
[Xl\�j�Z��X�KE��6�����P��D�mkE-J�X�m������[Mi��c�D��F�G��~�������]w�?ǟ��0	�����䙷)�,��]pf��zX%id���hl��Eaa�.�Y2�^9Mi���X*l~�*\����o_��(ݎ<�o}�G����VL,$�����`�J*����۩n�%�{&Om�_�&�X�U4F8���Զ��ogvd_~N�ر"�������ߗԦ.���Hb��0�y�p�o}�/�@u4C7��a|��!\M��ƩPy�⥻K9��fY�QSc��$v��9�
���36�7��"�q΁}e.��5On,���z���(�U#��CUn@���]�b���`�����|'�<�QR�Knu�fg��q�;<�哕�4��ӴTD`00�=��`q�L�<�]z72����,?_&\Nm�6ג۷�;�o���5�؅b<��������C/(�ftN<F�u�]�ڄTh~�Ϳ_9���9�Dإ��v�I
} l���\4�[��vv�]���t&*IJ(g*�.��!���9�;�ґ��+>�� wfT�����uK;5���6`f�6#L��0z���!�mBu"���p�V�Yúo��p����u�'K��۾qBsSJV��~�n>�*�әh�0;�X��c31�p�cn�%q;�R��W4����m3����ž�@S�q�:��ٻ]o�}ٵ��:�Kc�T�8ށ����BkŔ�}��T�̓q�x����V���Zd�����e�$�9�u��4q&�%N!�mW���p��ƥnh�B>O �#�n��6�#>V���K��tN���6���*e�K��םX҈��/ٔ���>��`�\F�'�C6T�9�u�@d�q+�hZ�IsW��ۮ����dZ�D����Ħ��}".�x��U�M�k�z�V{9��=�#U���P�,����R臐�K�:f�q�ق�d8ɨ��A��0bntRiFD����8�:��e�m�Ol.��Gx�s�3���M��v=oo�E����k{;[�θ�`��`d:6kb�Bq��L��W�e�e�G���)�m{��S��y�S䥻K,>j�k��%f�?6)�@{g��Ⱦ��}Nm?eI�m=zO?/�zC������e�a��ړ��H�x��b�LKغ�M�N.�L]��]�����V�$�z۠ݹW�o˲��(�GR�b$�$�����R�V��j�u㼶�V�y]X=BA{E>Asݍ�W�U�I1�rp�w�͑k
�p�{V��\&X�xn��{n���7E��%q�l'?n+��xwz����q�@�%Z�󁱆�C�˚@��@��vr�u�sd��vJ�Y���n�R���JA��j0���3p����&����m�*�nAQI�XX*�/�1��T*<Ll���rV���;9{ϵG2ԉ��V͚�Gt3��T��$���W�۵ܝ� ���U۳I�T77����A1,D�����q�����3Q�\x����'CMrȍ���f�;�u�.�;{��n
��H!N���c�<��SP�z�v3��k��k�f'�*�q���>bہ~
lT�N�
����c=��U��9���[��yq�!���{��Taَ����΂ u�7^8�%���~8�kq�9MS9��iUQ�g��֣w���6��k빋(�4��M4��yƘ�-O�o�W��f�&�8���wr�ilJ_�~H��q���q��#��>�w;�al�U@e55D���"�|�>P��VŨ�~��z[��?���6.��r}�G�eɄ^��,-b�{��@9�O1�U�s�*����3�#*,�@~>] ��!�b�Cі�*fFP���@e�&U�T�J��t��EM�ӹ�fx���)�B�~���֣:�}ZW-�cKҲ�2��2����o
RA�h�*q�[�9﷌�*t�[Vvv����1���k��$r;E�}�vs���Z�簝zz�ߦ�C��˪$��l�S]9�l�ؿ�\Kvȩ�՚�xW/�n�g|HuVt5�Mu_[TiU��u5���7J�!�j�ړ�i�e��>ڃ��"E���:��)���L����g�ggRU�=�5��W8�R�=L��������cj���è�F-���ئ[r���7��T\?��>�B�*�|�w��7�|�tm^�y�]d�/���Ny9��<���w��%���V*d�50SdA�����EC;�>FSJ�F��)�o�q	����+;�R�*#��!DA��&Lw@�	F�Ϲ߅W��p�n��t\\D��j�V�}�ώV!�Π��.`�PA�04X08�>�<��P�S�j܌}�+��"7���\��^��7ԺҶd���#~n|\W�T� �������mE����6�Gӑ/�&���C]��Q��9Ўx��'n���p�$���)$��\��Y]{�R����Y}���O�$�3}�A��'/�r-G��n�\�>K
d���vY�H�����x�R5x���B���'�2��.�i�ZY�*�w�����ğIX��J�aT�u�Є�g��TZas:ၣcX\�I,�����p�J]�X����
C�]��-���<�o!9J�.�����Ek�S���ƘL2PϿV�O�����k�!j�kܥ8�m��/a�&���OM!W�ڎ'�>��kim�s 24ɡ0�'�%�ȼ�^�w�%.����Lr��3����}�Wz�r�ܠ_���@'�셶d)��IW����*�P�n��58⦼�:f�Z�׼�%v)ڽ��@o�6V���lV�s P�!�)��C����q�39��:�H���ʮ����W�uI����o+�>&��qg
t��:ɳ�H����[TB~�`1맶��ͅYن{����߯�	ݥS��ò���̚�h9�{U���b�:��� wE����]N��SD#j9��M��cػ
���֑���i��{��l��W�f��%¿T�G���2|pG�Y�r�'N��=�;o���cb����׃���
8c:I�5��pi/i�O�ұ�K�x��m-��w�W4��z�
��̦����`]u2�(U����8��#�C�
�$#^2�U0G����V��]%��iDG�"�s}U{��rb
g)���|sI,��;�T��
р�v�9�(:�в�.�wc*.Ȩ�0j�=�c�*����t�.qb)�y=���Nα�)�����7��v8����C�W;�FA���w���$vM'��\�e��,(����1�.�>�(��xaa=(�]ʊ����ꇗqYYN��:���+���b�s�B�>V0�q����ثj��R��؇a�$�" ы�=>>Bނ�k�
�^5�}�q�1�`Ct�d9��';�~�n�ؗ�g����Y��x�ɿ-��>ۨ�P@�'DC9�hB�æ
��0\�!��h�=��"���;�X]�d�#S��B9�-Y�`l"̚-ɡ�u��%X�yĔ��Cwf�_=TpPS���-w9�j(]�SZ�FJ�s�B�p+Ҷ���N2�Y+6��O���UqS����j��c!�4�M�A�����ӊg���L���8�E�"�O"3f܉���Jy(܁��+$;���%Ӑ�1��%����p�+�cgEs��m޽۾�p�S�1Pz��i~̼��D=���`�l�LՀ�2�ق�d8ɒ8ˬ}�D��d��jT�e�<a�(�n#2 WOl,SK�g�T�c�)b�q��k���q�®*�K�92�� :sJ�G/VR$�e%�����$k���oT#o�7�:ZV�������jǊ�/F���k���T�d6y��Ҷ^�u^G��2[s�Q\{����}pp'�tk3.oY�P��Qv�И:L�����w��N����R�QØz��#��u;T|�N�\��Z+I��V�o�����n���ɘ��w���fL#��|x���B���5�|�Z���\���|��2�=Vw�.5z|�v�K�8o6V��(�=L�CQ��jN�G�.�!I�����b�$�Z��'l�w����$��'A�
��)�8
Q�
��1g���
+��E�ԉ�J{R�CL��ᨣ/���5�p2�:E&���8U�X�'u�R1���P7
��չ�%�@Od`2�Nz�pע�s��wc��bl7�n7��7�a����7&�v>�H�@��Ʉ��1�qG���S�O%H�M�Ï���;�+)���Ǵ�2�WrGk(�s}v�'�a�$��vL%ЈE�Tk����:�~���pQ�<Z����sJ#'�:1�W��g��sn�)�R�WOt����Qt�a��]��x����v���7U904�G�u�se�@���¥S�h �-:�t�_�vu��2�JȌ�ХM�����b��uw�.��(��a��f�k�՟u�zn��uB���na;���^��3*1�H����.iZ��C*��Wa�`�'\T�wndWf�dE�!�HTw��T\L]B�ך4�.L��W��x��ۤ�Q�8�˺��oEcW]�X�E8��2K]e�1pWO�>�3��w�DV�íkm����	{L�z�(ӷ�{:p�c���X[,Qe��Ңi�T��Y�&�zM���-�'��G/��!���q�8l���g��R ��=��X�P�)EK��������{������MS��&� �m�#�|(�`˫|<�.M/�u�z]x��e(ݷ�-��ѫe��4]=W�y�&��Z�j�1^�\�q�3�wćVx�/���PcSx��ʣKڪj0U^Ձ;�V[/�jN�Ȍ^1�Y��#�C:���i%���C)��~:������3��b����)�dv&�=o]b9u�������^`�Ip�yٻ���	�4�C"�P�
����S�����O�龎n_D��u!�})�c����c ���`K��i
��@IM� ����j�����<�V�WVR�^h�ܿs�k��bO��A:M a�#1	F�Ϲ�W��p�{�uǒ�S��p9��AT^ɹ�kЮ@�C42d�;��BC�,L��{gE"�&����&��n�|�%�Kl�(u\�������9��Iֶ@yi����y2.�S8{��)B�ئ3XZ��YCa����BV�bh�˝ʌ��$�����FsL���	�9�d�]w�ϩ��\�GyA*�H� �D��)D�a�"v�Y�״�M�O�{�Fv���;��7�v�m[2ncj�7>.(8 �ʡ�Q�t^mem��h�Wٚ��xڝw�4��P�9΄C6l�N��/l�L W:���L�20=�]T�R��u�0�&�1S�:�Id_lPWʃQ~�/��b����q�����+g5�L�z�au�3#C�=������B�}b�ti��)ƥ2Gj�hR�C��M�����ޮ�TS)���w����Z�#�֊�Ǒ���]/#.������QOg�`l��TٺgcS�79��(z���~�ņ��@j�bl"Ȓ�fE�T,�oa��*��k�0[���l�^�<�_��u�oS��Ղw��tj�\B�c�1�q��#*��ԥ��.j��w�1yt8��g��Q+���t}4���VL,�qt����4�eaX��[��n��X�\Ÿ����u�AoT�F,�	�[>�v<'�f%R���fpt�,���֖J�����:��V�P���L��KsWw�m�����z���ӸS�����Zy�Y0�b��v�q��+�T�*8�	W}�9|9K��!Z�t��{�E�U�aR��ǫ.u�o2j��X;�����9~{��S���N{5�,��NTt������"���1$#�9���0Z���k=�{|<�2�f��Ø��5�:a�My���
�k�)�҃����5��7
@/�n�mr�Z����n����W�/
8c:IT5Wl����^� ;�cB�MC���r����'�Q׏�yY�W	���P�"�B�(��JDH=#A�}AI��L�)m���s�����aU���������qE�e3�X��W	LH�dGu�3]�;5�%L�m�48�t?TIjyШ�a��us�v*ڡ�{���ÒI���\�%^�o �,�P4a�����X�q!�J2�a8̎�n�ؗ�dl
T�g���B�,A<�(��LB8�ЅчL���V#�f�!ͨ�y�z��|�V��j6��;5�!���`�`�:QfM�亳\<�v!ҏ�A5��qE�z�xd��I��،gd	K���sZ�F	Yna!h1�ȓ�a8�D+ }2j"�?��+7 ��l�����*������D/���N&�"�^�a���^\�ƝM#��^\�u���*Q܃.�~���+����7�XDw;]�U��H�/�Y���R�Z�mۥT�����C�b���ގ�ל7"��Aw|�嵯pb��s�K�U��s6�C�VNs�P��Ԇ��r��k6Zs��q8u��-�;���Ϋ_ �F;��I�]�&4+k3l�~<�POo�R��tj�ah۴�D��S1<Rm���]w����1IW�Vk��}��}(��r���yc&U�K��NӮ�{�X�|4NΠt�^��g2ݍ:y�U{n�y��-�	�r^_"w�ꩥgÂM�aƎ:��ǹ�ϣջ\q��ž,s�6��z�r�m�JnQӛ�IB_e��p����HS���1�&sQ�w��<�\�T�Z�b�,Ruf���яPH&�cuѠD�E[+UM�j��ۓ�n�"�L���]�XIB�����O���l�2��7��<�7���5װR��}�P�֨���4��)�6�tͫ�*E@�o�Y���Mڹ����h" ��vX���Տ.\Y���>�Ԟ�=�9j�z�4m;���Vq��GM��I����@��m���nB3�ux�m�AV�S�%����f=&]�*�>�@�l� G��5of�S�L�.}�$�-��Q���Q㲩$;Nؘ�g��4�V�wvk���Z|��\�
����2�3����+�[�)�d��QSYW�ĶO@^i��ݛ���mc���9ڷ��SJi���6��]��t��/�]E/��8��|�N�N�z�c���4�
���m�����ʷz����C7pw,;	b`(q���1w؉�Z�uԬY��I��A�N��g��Z�g2�7V�F�Z*75���ٳ�Ыy��*v����XB��a�e�8c�ꉰ�j�@z��de�'�v�ډMÁ�:W�C;8u��+6���*�i^$wˮ�\���4nc��\C���n�$��R�'�<N�x�����.���+��+���PV9ݸ�59��nt����'L.+j��%��]k0��j3yWNJ�`���D�L���5���J8Tٗ8��mh����7QSPv>6� )����6:�[p����t�Yj�����+E��ַ��mC���b]u�ʘ̴���7%��S�3b��v2�7���v�swu�J*�]!�0�{b��o�Lʓ!;�^g���wۂ.乂ӈ����Ԛu����4p]�[Ѣi<��}�Ƕ�B�Qݭ���(un;�ڲ{:W�Q��[�M��Ƕ\mY�t�<�C����J+�+�Ë_1̻�Z"���o*�wi1΍�듶6㶴��t�5i��(�bw9�^��l�ͮ�;
ʰ�t��N2���/!���c��hH��6�ұ��\�i)[�(��ըզjQeb+b��T�5�hٕ�!�XZ�E�;Ev5s+�
�n�\�梋*�Ů�T�v�Ú8F(1J�J���jj4+��8�5�7U+Y
*�Kh�ٷZ�ہcciqV�T�Z�ۚ�UMm��:͊����Y�4����DZ�%�Պ���jQ�1T�V%���e��J[R��E����ZQ\�5��8DȨ�Z�L9�T
�AkZ*"��d�Q�Vf,mˋ]�3[�ҘT�KerSWc"�e���!�j,��9EŹk.uҍֶ�J�n�5�Tm
��u%��ȹLm�6�+[q�����3���L�6�c3*Q�[����Zd��J�PU̊dc����KDEWZ�D6���QT�	�YX�j"L��"���o���ڊE]f� bnd>�yC��k&�ȍ�x��Q��3s.�EXVn�i&���{��������K�a�]u�v�z���Dq��WQj8����A�}/�2����HŖ�P_����������Z������ͪۆ�HW��vE���u~t&%5d��\�׎�\y����e���D�{K�L���,�Bq�WAlt�谶X!��,Ӎ$���513�����7$���5	�����(Z���`��%��)m����4���8��D����/q�AĜ6�سԲ��6>�s�Y
"��`�.#�e8�q�/���)��z2iÂ9�??O�f�*M����i���Llz��$+�fvK�"����w�.�/Ғ����C�P���#���U�]l�z�(���'�TT�+�ϊ�\����"���7:EsVn�'�s'Mz�TMgI(��6�ȵ=��<R��Wr�D��?Vv�c��g&�"s�_s�~���L�'`��<���f9G&���p�H�bp�z<�$�q�n�k�����L���'�jR(T�s��$��9��($:�6+n�=y=�<��瑚y�d��x��L��2�VPw�)>�d<\����K�R:]��`d�\�V�d܊�3���(s�R2n��{���ӂ���g�ԗ�U��Z&���U�8\�:�Z�z㜓Y���-fB�Ģ�᝜mw$�C����'c�,�.z�����v ��JU��0�1�qG��t�z9+Em��=u��ǻ��u�,����]+���;be�T8�8 � �:
PM��Y@��=��$-�vż��u��ۚ���ܤ��9Iݳ��&T%���C=1B�lz�G6e7�5Y(�b����B�dRn�����4`ٯ7T�)�i@�!����z��������H���LT�s*F�z�CZ��b�E8�A�d�iEa�I��A��ɪ���g�]�c���o�ic���b)�ܑ��t�
���E��
��Y`�iQ5���<����d6�-jYʂ�xܽ�[MQߏ����g��c?=���y^YN/W{�Z�,�YX8�qE��:B�o���X|O�W�».��>Q�̤^�WWlX] �˺�r}Ӹ�qcvGs���t�^�<ݙ9>�@Z�Z���5�%���#P��ޥ�LLSu֭=C#�uu�8�UT�`uU�I״�Ֆ��ړ�2#�"��#���_��Y���U���[6]NC:�Z�N��&��k��N������P����]��6-��ZQ0R�i��ca9rX�pB�n8j��Էq��v���;J��	�M�άt޻�*`�yԜ�me 뙷RhN	?P����_c��
�;C���03�k��ߔ�297��箶cp\�:b�yM<�
�Г�N�7�OX~�)dW��P!���N(g@ײ|�i�nƐ��ugE{چ�Q�FM-瓻h�� ��O�U��$+���(Q�s�*�<.���d~}wE��o&[{ˎNf�{3��)9QQt�&|��D�����/��;��뎁/;[KF����eӛck����-ۺ^�Pd_�����$p�I�r�X�ږ�����Əm�����o��ѹ�=��=��蝶��<&6�n|\S"�s*�{�_h�Kl�F�<g�.�r7#�~�#��3�i
�;J2�B!�6u;w&ľ�dQ$-���:��#C���"۔M�z���ۑ�-��{��
�*E�������.�Y��COe�Bv�n���[+T�S����}�5�eJ��{��XԪH�]BR�C��,UE��龼��;2,'1V��c��J��	�_>�*�p��w�盧qF��.���� �����ml�����\囶m2�m�(�m�!�O\^��(P0��z��U�-'��-��P�;{��x�uR�s6� uG��5 +x9�.zw{j��z��o�GB�ܳ�5U�y�J�{���zPU{�%��_}��f
�=jbf��fJ�%"�띀T{|vB�E�'q�T,�o����
�X��"J�{۬u�]X��8��"k�+�h&�A�tj�K�@���!��!�]�$E,��e���\ɞ��(n]{���c�Q+������}^��ҘX:\F�1���ݚ��Q�q=��[W�*F�J##��{ag���7�YՆ{���.7�Z��������sj��-�/}ۘ�(���>^�[:�S貁�yt��u;��SD"�8���G�����{ȯt��R�q�Ӟ����������΅�
����_M����嚑Owx]���d��-MdT��1��
�i��
6}L�%P�]�$+�'�m��-`��tb��mZ-�{}1M�*<�`�p�C-� �R/�ZQ́�qEDF���>���D�׆VuKחr��7G5�I�L��\��,c�]zGly�m��X��G�-�Nً�{�����{ݨ#� lb��!��T*9+sܧ\wh�`�P��A��)C`�>5f,�u�锋��0�����`5��yM�+&����N�
��tf_ZqDZ�7do.���f�=Ũ�����o<.P�Q͐.}w⎙^I�����qU�{�j32A�RU�;�u���n���]�ҧ�%�<�����8�86c���꯾�a^R��m�I���@э�=���C� �)B�[	�dv;v&����yo2E��=���F]����$A��8��.�`��O	p߶�׬�i�.T�;�A��׏K�gՙ6VZ��Ƭ����#��ř4[�YC;�J��!�Q1�=���'�Y�\Iy��B��	�k�����=��+���]��#�g����vS8�$�YS*�f��+���3`4����'��2h5B�϶2��t��h��e�#Y����pZ�R��{�uA���G�me�y��}�w;�-k�][��}����f���/S�����Fs������|y`t��#LTg|nܠ�:a�Z�`�m�S5nx��T	���rOc�V�0G{�U�ӢkF��5�~;mp�rb����Z}��^Y�[ok�Pf�d��r(��,wD�v3%C[(��P<1��;>��_*�]n՝�Z��u�ύV*�mUw)��
�;��<�t�Ǩ��rB�3;�̑k�������	S�'ػ��8�� �>��}�Wݎ�EC��;DJm�G�&�l�\#�l���ح|	������Uo�No�Fҧ��֗����-Z�w(��h<~��G�Do+�ѧ/[�YO����x�d��87^��O��vD-nwd��n��t�N?� < �ھyO^�;��YG���#�U(��{=F�m��� ��<B�3WT�Z|48�}��G+�psc�ͽX�Cmd��@_D�t�˰��ʿ;Y�ɋrvK��l�´��Kև���O�FO�d���E(J(��},���:BiPl���̳�U���sUo��\%�2��C��lD�ґB�{�ྜ$��9��($uvu�s��o��9Y�%�w��g��؂+�A)TN�&�F=�+���9g���U�,}@�d&g�a�1��S}J��]b��jx& ����	A4B,ʺ��u[��9�j\��m���z���<�p�����>�m��
�B2��{�T�ᨆ��'�'�d+}9��1W@�B��ɀ�.�Bnx�E�~sF���ȱ
m�ߺ$�RB3Ó<rovyb�HY�,K�f�T�9Yt�₽]w1e�7,�M(�6I���)s�
�ܻm�����^g���էpT�oے0�ӄ+�wu�X*�χ�P�KI���<rN'���U���+o`�Ha���ǲ+�Vř��F�>9S����;���iA�<2�%�&q�X06�/N�$��!�[i����4���pX�9N}G�ӻ[�0T�W3#
.ff�/�_+�ع�aa���&GF)�����U����kE]�7FX�F�qWd�}f�x����<�,T�@M⋣�5����}�L�ʇ���q��T��u����A^��h��
�.P��z��
��ΠC���ٝ]t���T4�����t�^�<^�͑Oj�흩}u�4n�i��:�Yыm4�)\A~��f�>�Ţ:����w��;:?�n�Cn�a8��P=-�K�Vfe\�=��q�9�gb�4��ѐ&w�s�򪠊��F��}����c^lFQ�p�Ji�Oo"�L8�gC"]�B�+"�VpTd����;ź�u�R�mw���<"p[��7�y�>g�|5xl	h����#^�PQ4:F�U�@@��v��H�v�!=����v����]����	��I#���<'�.�*�_o�c1@���g���Pp���rZU5Z�/u�;�����TtXPAJ�8H$Ϗ�q4k��-8���^^�vv�����H/�_�������-�fM�mB6����R��)]ɋ��N�F)`xȺ��s��n*/H�(lN�J{3ݠ��*��������Y�;h�=�o<n�u�Wu@k��8���	�/@`&�8ܻ�#i�r��@��er��/�dv]ܬQC9rbfމ儑9;��c�f������w&�ko�����`3������4�ҝ�s�͛)ө._]��"�!�4����F"VN��󴶼ze� ��
t�L>�����5�2�^S�8H,��yg�=L���i������1釨d�s��(%a}8���s����鍉��Q���D3�ޒ ��@�%|���4�
��~���')��=N?Y>fg,8L��y�����`d���!���z�/
�����ǖ2V3�w��ɘf|�}箟�{��edl��ܼ�Z�w> i�� ���t2���M�L��%@����ĝ���,�:�� �%E��I��)�_̝� �z8�z�'̝��N��p��W���c���R|���x~9��~]�����+�+aM�7�}�qg��$�����N#'�	���Lϙd�>��2r�\�����I8�C$��d�T�;L�Y�v�2)9J�G�|�=0�Ϲ�g�v�?2�~����g�a��͙�ߡ7�����|2���L��W��������
���O��+%W�ϻ��
E=I����+%O���7t�,+�<I�|�2��f{`Tx�����2AG��<�׹����*՘��"��>����{a����������7}c��"��Vy��1�S�|d�=���8B���œ���$�
��x�}�9AH�����9���3=gg�8@�6�~#��el�lլ���ߨ��G���0a����?N4:x`��VL��|��gOs���E*n������qL�}��{�ଟ2���M߿p)�A|N���x��I�'g�<�Ғ.K��.-l�U��C����>� ��t�3'N~5;d�įlP�3���Ü=�r���o)�����g����|���� �'�S甞}C$<��8�PS�*q��}�t�?�9D|����W�?2$�|����q�I�*_~����<0���C=�$ω�nH�z��3�hn,�ɐ=�pϙ9��z���8J�U��)�����AeI�~{���O��k��p�r=��ӭ�e�K�Z׻��ɽ�XЄ�M�Ϻb�����pe�V�Ťk�qR��h��K����%�;�&l�X19�q�h96�_V[�\�4��v�.�MY�h�ٻ�8+�+�*�we��F+����ђ#{�W~�����S��g�,�Ր(��y���)=OS!����9}`Tt{��T;C�������3ɓ��|a����o�p�_Xx�d�R(��q����Lι��8 A��xEtw�%��}6yrܿ�c�I��{��`d��u�N=�z�Ϟ�ؕ��Y>��8}`T�3�w�r����S����g�Xz³�3����$�"������dx�p6���qW=_a�~����o�C? �IX}Ŝ'�2��,;�S�������'֓�+;�i8k�'���� T��'!���*�_��Nӗ�C��aC��&L���@H��e��i-ϫ7q�ݷq;ݹ�0�� �26��I�Ar���O���:�����)��1�'��Ag3y��:E'iXvy��|�>0�<����������r�@�Y̿~�Mq�}�#��&`v����Ҿߖ��#��k�NIP�Y*���"��Z���TW�'�S�!���
���2w�>I�����|��2|o�ᝡX���v���È}���>�s?M���y-�ǧ>��5 �0����:N��P��aXTϬ���J�I_|��I�J�AM-�� ��@�/vO����Y2���w����I�Ϟ�礞�K>�C���s��ξ�҈�߀'�LΒ�ۼ釩�t{�\O����d�lp�I� ��㴋9Aԕ��ə3+=���R�~?S>�d��p�y��__̝�!�w�R��;qze�.�[����W��G�}� ~���d�3��'�`�_2g�v_�8AH��{���Ag,��}�<���2As��t��(fOl3����ͦO�:L�y�OS�QI�V{t%�~���9�[ͨϽ�2|���|>�䂤�v�=��O������Y9��Y2{�x��2mxI���9I�+''����AH����&{zH,��ya��'�S�'E�=0*OS��N9I����/�<���?$zg�\��P��0�sa���>a�}c���ô3�|�,��ty�!�t�"��c��aS甝O���P�+�=��`t��P��8����T�PY�9K��<Zlb����m�xFXS�B8�����wF��$xM�I�{�C�q�SG)b�B��&�u�L�`cx�Ш�e]�d"��p�-ʼv��&��7A�H,���ya�و�j\rc�]ݴ�B���#B�H�Lv�H�N��+Ԣ�{R� xx�7��������z�Y8O�[�>d�'����g��Ϭ��'hW�������giy;�3<a�frw�:gi�A}B�fL�������8~H���IO��G����~����ӻ?}�{��^}%@�R}�X8zJɭ'����A|s'oeH�|�<E�NgL�����p���g���$�
�ɓ?��"0��|�N�=C��t�'����+5��NU��rs.��>�_Y����{��gǞi8y`T����9N�|��텟���NҽOl�̓=��N�� ����8~eH�z�^�%��̙:���2m|g�# A|�Lp�s'�=V�Yٜ���x`T�q�䞾<$��w,��2y�8a�K��C=�*OS��ϸ:Cĕ�{>�៙P�~LΥ�,�
Ş3�i�p�_Xt��3�~C$�����dYG���������#w~��?~��d�°���>�(��Xq;�r߬��S��q�E�� �{��Ծ�:=��'L���x��n��W�Og߰|��p�|C�Շ,+X,|�H,������{�}�<}��u׽�������9H/i���'z�!�tsC>$YP}��� p���W���퓔
�N���Y>��u��)������"��T�{ǜI�����l9�"Oz������:�l�����u��v�!\ɓ��`T��-�S$~N]d��2|�<�z��C<�+�����>B��>L����8eO�dRv��� ���χ�{^��x��O�	�ʩ�t��={��o��O���ᝲ]g�:�^P=J�ɵ��q@�'�T�������,�)�O_^<��'��}N��<a����m�OS!�J�����r�}��'8*z�9yn�������{����X���^�����é��p3�|�`w?}�k�d�R/'�E3
§��3Rp��*���큒Vr[�R/�XR(���m���Ͼ>�z;F٨��ߧ�d��BZ�M���w�A��#��� W�w��NPX~k��|� �0�w�Xr�S$�{�)�=C!�Jԋ*����+'����}�d
�9�����A��\��{���~��MǳU��\�A�3N�ׂW�F̬�T��Vo� 8AՔ�p�t^-K\xE��R�	��&C��lk���83\�I�-��.�����}��xΒ��ƍ:�eɓ���r�k��gʖ_��L��]�z�ˍ���g��8�ӻtS�I쁝���.�\�ܦ�e�XD|4 ЬQ�&�oK�Z�١[[�)uvol�)�|�S�Pl�u[�8G���Y�/�FIc������G	ޜ�oF���d��7๗8<�1V-/ۻ.�N2��F<݄Բ�U��&�C��mJ�4l�����q%�אm\��&�,�o�Y]m��l�N�j�g�YZI��>��vU��T�sqA��/�N��
�^�5;
���[r���Y;�Blv4��N0�f�8e����m�~�e��|�Lw8�mO�Zޟ7�9)������� ��Yٰt��@R�G�y;5��ECH�k5�V]�A��a<��#u��$��r��W���f�3�V�ָ'7��!�b��쏡�aB넼��i����v��y\�6�@�kY��qj�|�e�ݜ�$GL�e�������'/J7/T[�Q#��*�Z;�9���%�+z���mwj먻��ʑ��Ed�������7 ��m5�ɸ�J߬+��ӨJ(���@e#��+h�b^i�]�jv��ٵ��K+�6��:f��u��^`�G��H�u�Nb�,�
�Y�B�lX�x��� Y�@B�8h!F*{�b�dŖE�k/���si�����:A땸9ӊ�G~������{�Q��bM�����m�Sy��Ѽ�I�ষ3cФ��R�"�P���M��w,�5{��{jW,��TњY�ٵUW�B8^�Y��O���ߵ�7m�i���ya�:�;��4es�:�f�c-��7�J:bIi`�L�6AqH�dg�޺�ܬ�Rn�}��߰rx�h�3RmwU���wsf�Ӽskrm�'�l݉n�JTB�I��D�������A�]��>0�����ց��Y�߈��yV���W�Y��S<e_<�z�v��-�oS��WZ�Z-����M�g@��7�����J�-]YuUy��:�a(�/�������;wb�D7�����g_�ZZ�u]F�w#�h`:�6��i�wϦப@c�Y	��%�Pn[��s|J��1wZ:f��J�����r�<=pЙA7Y9	�Y�S���������Vu[[C�Vm#�w,�m[�jɹ����@ �'����I{	ߣ�V3&���j�nqt!Y�_\f�Ucteu\2��/$ɂ�+�r���]�0�/+O�0��m��y5:yM�iK���#�o$��9��]�G�oY�����UX
�\V���tӄ�jv�͏��c%�����ŝ
r\}�{$�I�.-�[��Y�t���U���9�º��/ƪ��,X�jmr.\ZԅelsVУ�Ħ,U�J�(ёE��,re�]naEc�Z�j3ZR�kd����i+
Z�*�T��چj
:�K�"��D���h�2�*,��q��5�-s�D�u��%�F�E��V����
�J�*d��EV�d.��j*��*:�"��5�Y����R�m3A�Q˱iu����IY��+#i]h�梩*G%Ԣ�T`���eE�Ҳ�J�Qk����.J�ȦIYXV,
�cʅeԬ��"�
�kP�\�m�j���Q"�
��T˩�2�ə�YR�n�F� ���EY2[k�cC	U����T�TQ��lclf.ͪ�E&Հ���f�IXUj� $����V�R�,b��1+$L��fa�4��M��Jn��ϲY���i������0L���hM�����zGNn�s]��~�����F]t^��~������c� �P=Ng�s��'�g��;��Nӗ�O�?!��'hW�NO~냧�AH��ĝ?&H,�{�<�3�d��3�rO}�E�	�
��㬞�q�}�u߇��!S��&C�����2O��)����������d���oq�L�ʑC�~��r�.��;��9@�+>d�p���9B�}�r��
�����:I��� t--|��n�������>�����>�̞sN>����Y�~O��=I^XtsC�xʇhs;��z�b���|�')��~�!�:gd��+��ɒ���=J°�����>����ʧ�Q�R#��4��i�ۮ�����>%w�I^�����XC�p)R�b��fr�Xfz�qd����8I�>rO�W�VAa�Yה��*Ag���1�tær��������$A�d	'�I��ǧpYV��w�~����"ʃ�>pN*VO<���&@���H/�Y<��MC�$��:�;yAH�pk�p�2v�v�{9�z�=�|��;���OP��?we�g�� ;��vv��c~����/�q���FN�$���x��d��3>�d�(�'>M���H-@�Ϸ()�8I�g��`f|��C���*A~g��p�ô3�.}gi3�*E*�}�މ�i�D^}c�-]�:'*3��~�|���g�AD�}�,����Y�组�|�����hp�Y+�'=O�{��W����C�~N�%{N�,� ����qi�p�Y�g�;L�_^;➿�����uu�s�1�>��@���zN��2d���́�V�^q�_2�S��q�N_~�3Ϲܡ�
E�퓿~�H)���$霳�J����G�G�Q�� Q��2G������������y�}��>߾:{`T5��3=J�Y��5��៓$���J���:�yH/�T�����T�t~�O��<�ə=��$Ԭ�{ǜ�O�G�(��W���	'��<;�'��MMvk[�zH�����>d
 "��k~`d��^��l8N98��O� rZ,���O=�+��C����RXw�()�=I��ה��S�ǔ�ߧ7�o��5�2ذy9��|(1^�:$c[��{�[/N�������M�GoH�oަ+�Rx�Q�Ml�unJY
S2�u�G�^�-Ϸ�*u��V���+ecGIa�1��ܔ���7-��"ɽXgy�Բc0l���n��seF�3����9�ؗs���da�������퇈fN��N��L�ʓ�vԬ̗S�o�� |��'VÎ/�
���2fJ��
�T�|��׆{l��>�|+��>�A� o�����ט���ݏ�����A�(�z�����YP��pz��|����"��x��߷5�Hffx�O�}a�ɒ��@���Nm�>|d���I�}�38fC �_>���GN�)dTy�w��ݨC��#Ā>�<�'����^��H���<e|O�Y8IY�{�󀯌
����0Y�T��w��,3<L�G����T=O^Mg	�"�Kr���Fo�6�E�/M*������}�=�>3&H/�|qg�R|�H<�8���Ǵ�;��v�>d��~N�hr�R��9�}�O�
��+��'	�X����$FJ��'3����O_^���P�D���={��5O��Lo�G�0@3����r�Z�e��)�=a��S���S�N��?%H/���$����f����L�ʇe�����{�\ϙ:@�+:�}�u���H��__�ck��	��jy+W�A}�+�'Ӫp��J��ׇ�`fVJ�b��ӆ0�,8C$�<L��=�xk���T��~C'	����NX���d�}��<C33�;��x ��d	#�V�aߨ��S�T�u��W(�φH�x�����x�)��� v��9B���X���T���NR)7�z�~�|��XtӄS�d���������!���z�/
�����#g��I|v�+>��d�Ͼ��h��g�?&a��d��3�"���{��� ����q��=�T
���<I�+>�ɓę2A~J����i:B�d���N�R=��8O�;s;�Ɉ�O���_}�v>sy�����a�����y������,
�}�N#'�	��{�'���N~��2r�\���nRq��Z����
T*x�-�����S�,��H=F�ϒg��$�'{>f}���eMt�o|��������}e~�� z����;�6tɐ=J���|��W�gs�4�R�Uxa����"����߽㴂��^~��$�Ӧ��,��N|�2��f{`T�]~�B9;�����5�0���jZ��X�ք,��Fp����0ث��#A�Y*�u���<oJ=2ɂ���K:���d5�$$s�#�!�-�Pl�q���U{���ٮ���K�D��R){�6���x��J�Mr�ڞQ��r� xxM��Rou�����$�Hf,��I��/�:C33���� ������:NR(�g^S�'��Lã�t�9B���Y;��c���PR/�ߜ��"���|4�����O����%OGTo���������? z�Y8O����Rv��5��80*<ht��g䬜�fg�=L�3�*A}dR�g\����I���3�i*�b�|�������Dx�ݸ�O�������w�O�{�Om'�*O���8?�8xACԨ%L�Ӟ�;d��l�>N'�88{d�3�S��
Dd��2s;�fz���z��$$�>6G��H�p�:���؋�ws/k��Tm~���)�
�C���2Ag���︇H��u��p���3��nìC=�$ψ�"��Vrέş�2�S3�N5�^z�J�U��;��#ď�F)�}��7�_v�/�m|	g��ʓ�u����)��W������>L�_s����PY���P�$:��8�!X�0��8@��2�;��8H/�<N�ӄ�*EԺ�I�>(��}O���?|�~��k�<����x�'(T������N�(q:�7� �^N��)ǖOY��~��'���i�����Ow�r����S��aa�X,�+XVz�&a�J"H�'O�H���Y���|#7�u�|��O~
�!�A{O��g?RV�g	�'�Vy�gT�����~�r����
��Y3_�;xAN���*T���7�q��%@�+�>��$��?0*�@��ޒ$�=7��F��M�}sۚ�^=�
Dd���Y�#iư����!̴?<$����͙�PS�/3�~I�r�Y�o=���H�a��$������ ����ӯ��A_UHQy���m~z�~�a��_j���I���&I�����ɵ����J�J�U��h

E?"���	�Kf2y�8a���
���2xw�>I����o��9C�=L���}G�@��|χ-�rD��Guf;�Z���e�@�ﻲ��G�4|3���I�T�R��aXTϬ���J�I_}�I�T*
~�Ϭ�Ír�{�|̝�d�������A�� �3��)�]⃁���V'#V�u;P�dۙ�R��md�;�����0^jvh�ˬ4�2����s���;u�ufE�\*;)Ć�ҥ�	��u�]R�Bqn3�a���Z6��2V�)����|��3�����\fq!�$sK���{��!�?%o���e��@���~����,�*u��pΘz��G�u��:H/�NÏ�����2A��q�E���Vr{a�pəY�uhp�R�~J����I��������9�u��7���6�}�\f$�~� � �@�fϸ��z�z������
������&~gr���A>�͓���Y;��9�O�ɒ��=�v���(f�g�O2	G�"H�7���ﾬ��X���w���~x��ɘr��V|qd��|�=��Щ�ΐ�w�>�*�_}���sg,�v��M�	9��9I�+'?{�� ��?pL���YS�,8{d��p�İ������S����q��߹���r�'���'HNC�N�铙� ��׃�t'�9a���3�I�~�g�8I?y�=dY=xI�ċ%��U��$Y��R>&�_`˫�Ϻ�X�'{`fO�� v�Y<NKxg�J��y�ְ���
Ó��>yI�
�I�6p��v�����ə�}�v�$�/�d�|���{�?$YP|G���;t��;�������"��g՜���%@�Rq�8zJɭ'�����N�ư2�S���3�JɟS=�|���$�
�ɓ=���$��s����Ag�y龾��>C�����r뱮9�y�{�YG��� <$����y���Rs�~��i>L��}���~a�;J�큞ْg�si�$�v���
��Ι/~d��4����k�;߿W�߾9��L�i]��j��� A|>��$��Ox�Ԟ?<$�=�r���'�ӆ���!��'����pt��+��擶p�C���["ΐ�Y�8��8H/�:N��័���w��;�x=�//����^��Ǐ�P�8@�}����N�Y��(%B��7-���*9<�$_>�2{�'����)��|}�>�)��l}�u��F��lfw�6VL��Z��"�J��w�KnL�h_D�A,�N�v�Xf��_֕��y��W��M6���^�ЗY��� �m�˼>�YA�guQ��u�t*@��Iۢ��z�V��i[o4p�2޵FO6ڹ넛�D���oG%�G�jt�y1���2��I1�kS�֫�wo�����o -�k����i�`�y"�KY6ɏNI�}�}��U����[޷�O#��'����7Msen�L���q&o����.2�:E>�c�jT���Q3M���4㳤�Y9]
>�7�J1�g�qCJE
��s�_N��=d;2��By�6�
���B��;��"�u����Ƹ9C������s�ʷ;\a��\�e]%��f�4��Gf�(��w<�4-�"(K۵z*[�r`��J	���0��q1	r���YM�Y�s|�=+�=�);�}bہ~�b�E�ED$7�p����d����Z�����']Y0���0Û-Ę4ZJ�QȞ�W�!zW��Iy���}�Y@�u@�k�q��v�p���u���c�(�k��$���u�L�&D���N��ܻ�nym�\,a��>�_��((J�Ӹ*S�67$a�gN�w;��ĺ�ⅰ]ΊսOZ���*�ot���x��Q�]�[�|yz͋|��t�ns:k����I�)���z�ڏ(E�N��ͨ���EQ�a�O��������>�hh���hθ&��D�	\�$���Ԅ[lU�Wo�q�o��V�ֳN}�X��SK%�,L�=�~�f�ƴt��%
��{h��wR`�|�J�oT3$�C��qr9�Ҹo�p'Rw�89¹
�:�u�y*w6䒥`���{]kJ�h� �j?W���}U@I�~�a�l����N�y@z�>�.���:p�ٓ�:A9'$#�h�3����򴇧���Q^�*���*��	D�d��>�p*�N��u�,�-�}�rx��S)Yx�{�b�\�n����E�Yq���B��h g�w��򪠍�=L���I^Ee;w7���K�u��n\ᎃЍ��+��Q��.38*�|�oj��n��y�6t��pj�9�<����>=r�$ߪ����fx��#�Ҕ��6s�Su�95��o�w�}!n`wQP����3�Ұ��$gF(7��B$�0�>��SK��vCU�7)�[w�J�ϳ�^���s�î=�K�.8��k�
��t�"�s*��YP�.n�
�S�Gg�}ڂ��#�X���8Ddr]�²��	�;Bڶd�لt7>>0�y�,_�޽ޛ �_���o�6`3�@[�ν!X��(./�8p�N���q�˗�k�%{7׍S��U��$�~s���A; uƯ¥t;�$q��
�Pj,C��p5dɏ[�ؠvV^Fn:̯n��21����pM
5�#muh�����:�갬D��t�A9|WG��]\���g4�m����Z����މgS=���M��֒w�ٓDlXSЍu�fM�'�ь.;������$៪�����I��2/i���T~���YD��0|�>��u�X�]
�;=����Bi���5&�qH���t�r��Kq
0C��P��^V1��M�r}r��i{R�.uE���n7r�<޾-�uPg�b��J$F����ԂzA�l6AݼY�#&{رG޾��K�cՅ�P��҂�D�y>S���iF]�q�n%�Փ'v�޷J�a���+��,�+�̑�4n]o�2�/��_�y�����R,3�ҹ�uߩ>�@�}՘���V-'8;��8�S�EXR<�2���{agT�F�IgT'�y�{Lad�g��dJ��k���	ݬ�`�tmp��tr1ߚ���g�!��E�n{6�y���T��2bHEP3��L��U����p���^gB���l]z�)oj^�+�4"��5��7��"9�m�"6.��"|H]fd�S�9��\�n������aӒ_Xڒ&�J�U�p�C-�J�|9X��j�h|x��c�ݍOfO�c%;��s�MM�<��U�{S�G�(�̧[Wq���~�=��SJ��+�\U� }�_g	��Y�G]d�-���LF����:p�qEP]k�i�\�]fiy�����L2����C������Q���ֺEh�i�˄���� �����M[|$y!}Q#�L�)eԑ;��g\���.�>�(�s�l�3��)\s%�����甸B��#Ù������J,TI��Q�^��cj��Z��o`�tRJ27�g�V]V��4��C�$��`�^1����C؝q!�J��;Q�&͌���|���;�����X�����WB	J��#�s�1�B�����4\��z*4e�yk�J��q��|�����.Ĉ:�`� �(�'okA+��XNB̹��8'T�p��(��$����a�lH��'�4mu�#8�]I\��g.�Ə���|��L%�I��їC�ͶB))��Q��M�Ԉ>�>�� F��Ŏ����ݎִ��;(�Ah�1��U�AdY��
���Ȱ��.�:�˨���K����&�eߩ��]2^>���eX.����AVY��vG��tћ�7HUY��fg���ڤ�Z ^򀎘����-Xk���<!7g�Luݫ�gY���y읶8�&�9�>S�E�5�
f��Mh��ega -�w��=1�Xy�X�[	m'���:r ��Sl����í�}V�Ն�cZN�3Z��Iuj�pcw��b�[��آ��C:��Xe�y���R
���}����|BqyS5Q��5�
�<��(,U�1�݌6dFW�HY`�!T͚؍sz��RޮƖ�ۈ�N��G���F*�|�An0��<p>�1�`�#����K�Ȣ8�<0N=^�2"^~��e?t��[w�d�u׹H��J*�u�Ũy���K��#���^�qs�uw^����Q.�Ʌ�%2Y�
Iѝ$��:�r�̵R�&q��ȻŚ���V�_G��\	T��=�����2�~=�ę��q�\�)��w&��Y��Sz�j�x��^5윮���s��B��AFx������5�d���Dh"A{om����S��tg��"}O�ķ�N�'b`���� �����<�.�2��i�q�=�W�m��wݯ[�iXot��4<Lm6�M7�9�)��l=�ҿz��I�ˇ6��X)I����7A�i�����u���>z+b=�dH��ϋ^.�S5:��C�E�+�Ʉ�Mti�EЩj�F�;"}�-��N��s�m]��=+�����C\����k��_d�� m�|��t�}n���\��Xvm��v%ǩiá�V�]�4%ꐤ�o��g�++:e�����m/�� <=4�9*Ʃ�ZXM���pZ����/���P�p�c�rz�ߦO0�t��u/(5�PS����������<x�x�2AS��C2��������\���M�i}�b��zAմs$By�*ތ����ft&�w�����/��Xr�T�hO;�w��q��|e����B_��󧴋&1�b̆|�y��=��T�XG�n'��wUK�Ok�=jX=�Ss�'��� ��DsQ;�kV<u0uO�;���Eޔ��~&��C�횻�A�xb��|��e*���{W|q�Ӽ<���@N�L/�^X����U^)��vS|w�J4��N����~�Ui�ԩκ�Fޤ��H��c�1�S-%0g:���J��Ļ��+���7��$�|�����%Lh��G�8��u�IN'|�\��`$
��x�U�S�V� �Ix�v�z�e\BsU`G�t����f��z��E��Q7-mJ֦ /w��Y�F���e�� xosw)�ewrri׫p�����M�ش�$�f���f�b��Uw�A��omŋ㠋B�7pҥ=�ՖQ���l�n�EN5�Ҋ�@��yV��F�w�����CѺw"̸F���gn�w>O��썖@�:n�CHNz��e)PӓyG����7Gu�	VZ��-��� \��>��Bc�%]]�]�
�h��1�r���]��2�l����-�Γt�WK��t�`F�#��B��#�����x�3m1u��@���2#Cx�Lr��֬�C��u_���:����+N�.��D*=ќ��^���+���_b�mLR�Ϸp� �(�X�C-i�r����WpcwZ�K�����[{K��[���e��C�fN���i�\L��(WUǥ�-+[.�J���:�$�f��4�ti`�;f퍖�C��S�e`)oU�WND����.�B���p���К�]��n]���xt��[�hS
֒үkY���U�ݷw@Td=N�tj|h�;ݖ���IKWb�P���Z��$�:��1kxʆP�j�3��};8�ת�Ψ9���%�i��J�ѥD��w��+�7g�٬ܫ]���:��ĠEx��*`��i=��tZ��������g�*�UʗwN���k�O�QIi���2-����γ�1��f3����
�@����W��Ҫp��)@7f�,�w��y�D�]���(�O)Kօ�ZZ�(��������E���0�eSۥ�3l��RnU���#; �e�4J���XU�E�����%c�ʶ�
`�Cmp+6�N���OQ}�5=�ᬺ�m��
���65�g%�:a�C�!�1r��Z8\w=טV��\]_uX����X|� ��L�ǵ�]�hp[��y7i۹�Q�h�U�5��7�^P��U��DQ�c�W�僫�s4�=�t+vU�'/Wr��RM��3 �u��������'aUxz�y��M�x�J��Tk^v���07�$�Գ�Km��TB�]x������-�ã׹��Ҿ���v�luS��/���Ј��]��g*����Z�U4��ے�-��J��g|�T�{Di��WK�3,T��O-U��{`�K��U��m����Ǹ�]�79�e3޾{9�����"F�spb;��@����+z���OvY��ӆ�N�e�v�͚�p�����2�/"�c��Ż�&���ڧ!���WȧJ�C����h��q�u9VnR�2f�o
P��L���EY�*зǊ��7��:o
ٛ��w�,��W¹�t�Ł���f�s��I�̖�q[�}Z�&�m�="�5le�aw	ҹ�����9^��	;:��J&��R|AJ!ۙu]��[h��]r�`d��-�-��Xۆ�EQb0�f���aJ.���.��!PD*l�J�
*�j�UE��
�@��XkL�PE���SZQ�U�j�c%+���U�-���mZ#E�r���PKH)3.��V+Z��%E�[���Պ���,a(��ڙ�-C1@ȳ!XƦC[��P�eau��J�*L�3i�kDE#Z�+Y��-h�PR���J��փ�R����ڪ,U��6��*h����+��&қ�T+��vp"�Sf���TS0R*�tajX,*-H�+��V,Lږ��XQ����L���\!Wm�$Z��T*[Q3[B��fKJ)+I��Wk�RVT̨aZ�X���Z�Z��3��T��m��[H�.�d�Ńh�h�]LPS2�:�*)v��U��J,��Q3Soo7������l�r����sqAp������N#����)̮��r�L����]��^�����W{C�0qԓ{�b��� x]��Z��cN����Pw���0�o�S��}N�=K�vWw<W�1��މY�u��g(H-��%9<�vx�{�c&�8�{Ih;��i��ћwk^Og�_�H��R
{A�ۨ���]�Xy��98�-�Ś���b/�l`�RR��<�hJ�^��CY~��>�������@rK��ݿ�@%QmŰ�8@t��cV��]�DO+K�Y~֦��S�w,^vs�����5�t��^kq}�l�ˌ�H�əyu�Ҍ�N��{5kIL���lHiA}�c �zN�o�U��f]7ۍ�0fչ�{z�F]Z�s�R��SI�-(��+X0������b0�]��6�\�9@g9˭]�oy?�}l�9$4�
�ݴ�{Λ��x���u�@q�㏨���c��At�_L�~uk�g@W��*_��؃c�YCh�v��k]-�Q��즳5	�nT��b��".�Ja�|����[����"��.��� W�6��1�*��v��b��\��%%�������2���<P�]g	���0;�|�s��Kt�Pg
Z%���0�5%�#rEؔ���ꯪ��������3�(�����X�6v�W�:�j���S�q}��H��_;n�ZCrԗs��)��s�M�(�����x�Uo��G��Z�^{���ʀ����a���v�9\�(���.���[��v��ט8=��C��Q�S#��ꯇ7ct��(���0����s3,�Ugj[:I~=�Akja��iI�����lci�)� k��8�=�XQ#Bߪ������n��҂�zu�K�}�_tZ���s�l�,W۫V���뵱BҰ����"4$0��TA�z��r��=��ﺃ8���S,]r���[�i�V
�/%$l�&!�F;�٥���2{��5S���uF��h�T�<�m�VR����ˑo$NN��k�V�
"�μ����wB��97��-�k�ۋd�q;��n�`��&�+����KJ�ƶ����չ���0��;Փbf�)(6_L2��5��]�`��wbL���l��F�P�L��l�f�&�J˸�Ó:JT����ݮ�*R
����]��R��O��Zv;��nN�����S����U?r#L'x2�W�^�IT�Y���iA��eܛ5��+�1���@<�kF���$Ul�"�D߹�������f���Z�v�՞�*0g����9�<���9���^���έㄞN3����$��}�ާ�'��½g$}^9�![�Tnk��u@U1�uҵ����.��^�>���c�=݌Vo+�_!�Ŝnh������c�m�C8G���|�)��x���Qb-�,�S3���?S'j���P���/��\%IPS�lsZ�st���zck�S��
��+��k���%�!�2�si��Y�15�A�s�����N]�?d,�K!/R&o�(=ٞnver���' ߰���
�s�mu����vv<b�pH�tP=�AiR;�]�*N���B��Ѯ����J�d�C��D��یwJ��{Ӧ�w@w�]E��F3�އoӵ�"�7�3n��3ι� wm3u$�����IyR�Fvu�6:�U�V�[�S�;ȸh|Orܘ�7�˱��7zt��gn橎nbt�N?�}��|5�~�g������g<{�k4����v1�.���� � �G�p�Fo-��C�E*��M�p+>��'�^�N*Ұ��?6IN�}n*�[jUb�Ԇ��P��L-��[ɥ`����N�X�6�{��Y���u��r�Z�Uy���^���=��U˜����팢0B���{4�J9�~��ҬVA��'}k�"�����"����}�@,�r�+Wd���cJ"gp�1		(��0Pkt�ڴ.22x?���۫���~⽘My�v�.~��SA6!�1�E�Y�;rx���#�R�Զ�`���zN��oe�<�����9������f��m�קf�mĶ�jC�8�{~��NH�=؇�w����{�#<N"ױo`#0Ƌ��L�<Z�nQ�v�<QQ��z��|��g��x�;��}��uѨ!gF�\KN�����y4z{�8=�F��J��|C��� ��y�9�d�� m����=KSܫE���l]2�M��j��$�o�Nn�ܺm�ݣ�P]!ᚥ�\��wnvj˅�}��M��Y�v�؃��7S�{%e�1�c/��UW�jԧ���0��I%�~��+��.v�؆���������+�8�����otê�߆�]~��޽����y]xƪ�҇u��N�Û���}=��}����ۯ9\�GgX��b�#�Y�U1��g�=t���SFo���w~��R�M��a�Z#C�8���fi�]���ͭ ��i��D���ĳ�]�m�;�4������{�U�����'��u0���><�v�w>��8E���UQ�S�y�����n��o�lx�$���g�O��W�KFC(��t5U�{x�~�����c�B���V
����y��׾M��ɁYn��l���5ڲŤy��'1MŴU�:
U�0^܌^� �����9-+���Y�����a��b�nc5�+á��V`����h穜h,�{L��C�cל��,��+�{i�E�z�շ ��\&���Qk�e=�vE�_�=�
H��yhi���v8���r�����U�%�v���Ƴ�8hA�zki9KNv�Z�I�j��ؚ��
J��{����K֞�TE_ӯ(e�P�Z�S<��5�ؖ�}���[����&�8�f�c�y�ڝ���s�
�BF��s�-a��S�5�W�j8����:��	QL���t#5d����>�,�������O~���k�2�k��s�dD������& ��b����gV�]U��x�� ��uיTq���dM>���3��μ��*;V`�9�5ul�>�b��%b!��.m.�/DV�~R��
e��r��y�;#Y��������9����0���!����/���Q?{Mz�p��ζ��߫���t�s��1:�v�\��S��A*#����_n���Rh��5S��˜|�R����`���T�T&V*#msy�=�a����.�Ԕ�D=�㳤��8υQ��O��ϷC���T���=�ov�r$�lt>0^3b�u극g��:�(r*�$�Iܫ�sv�#;dg�6�_�He ��Xʊn���_���b���jL�!�;�s(2z�d��A��4��r���#s�7k�����]0�nͣm�@�±�F��������s�� ħG�����[bx�볬����K�T=�ز��)���Rw�HZ�"��HF����x�6��w�{��Z��ݫt��;X*��R��7L���������2B����M��*s�_�|]��T�<�sl*7�AI�+Ψޘ10�Z���cZ���x���{-:��T5s��o���k����ku���O8�^h���;=C/ϭu��x:"���	*�Y��y6�Q� ϣgv�j��SېX�q���p�|6�C��T��7�f�JOzn�P�yI��(�J>or���Q�&�'��-ɜ7P���:�����suK����ZƷ��^����k6-�*��ꪗ�3��#sV�i\*:��t��L��T��������,0X5fRϸ�0�(w����kcL����	�=C��ƺ_;�S/V&�_�=�z�6+a܌�
�6�E3��d�ǔKnnCIpv��yE�f�/�9�#�o���EG�U���k'*��Z�F
��Y�o/�����XQ]QB���(�Cp��J�g`���=ھ/	"}b��+�
.Zn�8ޏ�/����]c�0w	 Ro6�_x{��ror���r�T
�==BP}^�"�!;˜Z���y�ɵ��f�����+�)��yb��*���x�_�����!>�ܗ�;�4��
.*�g<�:7�k���X�Ȳl�5m}��y-���De\��56�.��bc�-����N�v;�1��"T� ����x���
�0߸ޗ��6�'���5��}�M�;�0�~J}&뢱E"*C,���}�-�m�o�Ԁy.�+�y�n�P����[Z��^=��p�v�S��t0G@)�/�l-�Ұ�l;�	��[���ټ�n�m��t(+�������	��
�s��g���Ppa�С���Ac��;�4�����R�����/��Z��
\�������oW.��Wia6$4��>��^kt�[�]�`Jy�cnn�;��.C��9��(S�4k����#^sw9�V�9��k�q��\�≾���G�D��HeCx�/��ŇS�=�\s��)
�f��QN9,a���J�䏺�=fwb�dj��ʖ���$���b
*/69��8Šԏ�������o��7��sk�>U5�)M��4���CY�:��bg3Q�u��y�+39z��(t�'�b/W��zoOJ~�v�X%}�˲w2T�ͦ�s^�/(bs�Z��2���h>�4�n�L���gfOgl������3+/�5ϔ���L�lA���s��U�/y%�'+��؎��2�R���WΓ�D��V��|��)ˈ�V�&�=y4w�y]�Ba�zP�Ys�BPd�9�Kg7V15n�h��s�6���j;:�oa��"`��1�f��/9��V�����gLo�L��Q�|�O,c
|�NμCW�%E��q%ۨ{6�#�e���ShL>V*��oy��cT��C}ND��r���;m���b�����Ҡ&T�'���V=��[� V	��zԮ��y}�]�zgc��|�3�E������E
����fR$[ ^%2m���*�Q��N�*�px����c~����M�V-*'gz���IW{�ދ�/�W�]�e39t(1V��kD���	;�溉Hg������~�~���~�������)	 �}!n�}��d���یa��yZ"2�:�>��4�8/e�*�U�%*l}4%k���ڳ�vо��s�.�#_�5+�o���P	�]���8���05k��Y�V�5�o��8�IgT�%�ԣ��I�`Ć�.���A�q@t>�(Qs�ɱR�1�=��b��/��[��z��Myc
h&�J>��3:+b�(���sˋ���z������*�C�G>O��^�ox�ۇ�c�d����F\�ɣ�;w�[�}d�d#`��_��Q�3�?���c{X
�����p]N�۲�u�wG3�q����nv���J+��w����w�
>h�g���צ�?Ok�?$�l��`����N\�iSkM*w�G1X��ߋ�n�<��ƇK�`)��yʾ���Ց�Vxw0��ഺ������!Y1ɻ*�͸RF=y���o��jN���/5�k��Z�H^$���+g �'��o�xm��3l�5��a>�l�\�Ky�����a�+�U%�X�*0�)vP����儾>�1���:�JQ,a�\
{,rj���volN��mh�$��ڌY9�{��2�jp'�X�ƨ΁ՓD�wұ��҂��;%C�ӆf�l�^n;S[�A��/��b�w_��f��]�g=)4���uY���sLf��Z�V+�sy2[���, �vʒv܉�	L�y7m���q����fg_l٪��m��}w�k��X����|B\v�2�CCU6 %M0�gWgG9Xo+�$Ԅ���9��֖��{h!�[���Fo�����fa��P��1���v���܅��Ѵ��1CϺ��N�ꏅ���M-�ErtOe%���}@mD)S�j�L��X<QK3sk9t��idC"�x����C��V�ʭ���L)Qf]ϥ�c�I8��,ڑ���K4ڳ!w#�V$ZMPR^�C5����̽gP�`�_�U<�6SO�m̚�+��,P(�V�ã� $��O4V D��ή�O5Q��Qm�e����M�ͥ�SFV�tC%]+^Lp�";���F-]l�s�ᖳg����IF�	�L�i�촲v�<�V��js����M�P ��ww3WX��;ˁa��=L܄�M�6���s�b|ض+Dz��S��=p։D�o�5����o���Au]&�^g�FǳRTD�X��=�e&m@5�h���co*���ހ���+�ڹ{!z�;o�Q�f���z��M����qǓ�gV��b[ ��p��<�3{(u�-�X�8��T��/�ʭHͷ�6e�^j�R����٤���czydټ��U0u�]�{b�P��h���լ�����p��wUqV�0H̴��َ�uH����u�Z��.�v��&{N_,l��!��aoc[oa�\L�i��'(j^4A���wN*m��c�`Vn�D��Hu��]+���p�p�%��PNv�ۥ���oNN�wp�M%�s�x�BwP�[$�6���*7�C,:;���;�tr�iѠ��̦��E���eo)��.��hd��܆��߸q�cSs9�k��7c"��+�>�5|��0�4U̍ y���¬�X��ݢn�}�OC�6�7�;+39��2�gf�mt�,�M7�4[�g��k��PrJu���vv���ȋv��=~�>6C��A,ЅdP��|��;�s�lձV������㣡�a(x���L��#ٔ�P{����9e���t{J�fҴ�k�5>N���*H5W\	��j�:+)�&U�NC������n�vB�O�$2ٓ��-�:7Ld7n��x[S3��­n�n�W�a�.i���6�X@�Rn�� �^t5Yp@c�j���;�Tr�͛��$�� ��Z��hͤ�ʬ2Tik�L����ҵuт�j�X��nu͙B�fe�P�QID�cQ�Y��
�j����R�fUu����jL�کQf�V�YZ���3*�+�K�Qb��#G8*.h�iRW[m�H5ɝ�n-���ډ]M���ԕ��VfWD�X#��(�V[b�)R��;UY\�E]��T-vXVLk%V+�
����*�5Ȣ"�U
���Ev�ԻTZ��کP3��TS*"���̮v��+UFV�ee�#�V[c��mKm�`[KZ�k�;"�c�Zљ\�#[2��.(�fjJ�EY�$�
&GR��P�J9+R�n؍�����s��JjB��s
��PL�Mi
�]v�T���݌ɕ3Z˩uʄ�323,p�\�Z�"�RF(� ��a�	Z[Sb�R(�(���H��HUR�fmJ�"(�Q[�q�������$�)�-�:i����5��U}�l����)���O���v�}OVs�}ɵ)��6MkV�T���?U}_ў��a��z]zt.�d���z�ss�ۧ+������h=y8�A�T����K��&P���������t�'����htr��Np�)>qy*7:�.���򩄪a�u���a��,�z�MkP�������v�G���0�/%"7�ƼZT&9;���Z��я���پ�X���݃X���(C�V���?$B꫒����y�b�V�;���M b+Ӱ$��U�iZ��{��tབྷ�X*����f�Aw�#pԴ��atAՍ���^�ҿx�ŇKBt��ͻ*ÁE����DuK���mm�!c酷�i׳�{W8M�hĆ�.[�r�l�'W��;u���Z�.2�+�
Cf�rjS��YY�U��M����K�7�rozc��{�]��v��屁�p��@�ȇِ�ʈ��ݐ��O{�˷z�ϒ��2;Ŕ�V����"`Wj��G*����ݢ��&���@M "m`&�΁
>󬆁�u�k�ۘ���I�X�d���ə��b�W��Vg�7A0�=d�:�N��ER��`�����r��	$�c��W��yQ�[��_j����D��}�Q�ӵY;Y<H�,��*N��$�+�÷k�r�ޚ���Z��9ߞ˗�47w
������9�UQ4���aE���kX�j�zv�P�.���L��ʾ珥�Z#�$���l��mf��Hv���Ox��]�`�U7;S��B/�/��x�7��̺`��&�)���:��7��sgd�`��*z}��_'ys�T��5l4i3�.#�'ɸA=��O#:��ˬƨ/�J	au����L�V�����Ls��c,|dYK���|��c�!�4��.�cb[i_v�LV��Z�������1��$Jڬ_7l9v��˩v\��S��U��X�A�g=}�5����1�.��Y�.�24W-٩؝续Ck�vzB���K�+y��;t�iW^������>_|8����/�P���"Z�;���q��Ep���Ԑ�P�M4ƩPkz5D��9טR��*�F�e��֧��V	��]��h�����C]�7�t*Y&Ew�Hj}�pރb+�ZC�,a��]��h[�k&�R`*N_���
�;��r{+P+�~� ����V:�d_l.M$]�a��{$��3tء��4��<�Xt!W�W:m��W[>������_l*�.sNI�̪�5ťV�F*{��A*����7
�WAR��Ƚ�[�{�!��O����[��ң�]W��fi�$4��>��A�qC_������m>H�	�,��o���bﲳk�:��X�lD��}�C���m�y�#pU�s/iL��V��cN1�.U��y>˫[�����R��hO5�St��(E����-o��]�ö�D�9^��.�_�em���9V�� ���R˚|�NaE�K����^(����B/�;S<�,�y�f�N9n������,B���`�cz��ڔW�!�!҃T5��-1�a
��je+
y��7��ױ�Vxr� �:G���j\�Z��׃=��Up3�Ы�Vh�	�cF�v��t�;s�0��gZO2l�y�N�7 yQ��-���w{O�[ϖ9嶍w 
�1�,�u%6+��d�{c���޸��kr���xvu���M0c�f
8&����Z�*٢T���\�UU_�9��u��
�/�h! _2��m�\�(���C�%|;zV���[��%�z�w��3���7����'��)	��Le�(�h=��ڞ���\~zn�}X��ja���l.o�y��Ú}ѓ��
���x�v.�=z��хW��;�ҩ��%��仰�uI�Ҫ
��9�[v�k���v�(B�V�]y�"6�HI����}����<��ͱ*o�;�-���[l�����y,u�IJ�#G>�Z�5��tH����z��������X-�v�I�]�Tq+��<}��ck@�5�^����~'�E��%��2�ĵ�t��A�p)e.ՇNO�<�ǌ��{��{��ਈz��/X	*�R������p�IN&�12W����ȿx����)C�p���8�^�ܡ텁9�"a���:���#���4�=���w&�M������YPvѸgU�oz�)���(��5�A<�#{���n�DU��%׽ԃ���N�z�c��۵:P\�:�ٜ��'oy��2���>iDyF�\��,�zӡ;]I6TI�?W�_W�Ob�(�����o;t�_�y�7;�'X��H��n'��c��*/4�k�wk�7xw��ox��{���v���1h���gJ���Q����Դ���jg��2�g����c{��a�8���H��2�����;c���u�"���m����{�(��[������މ�v�,�ʗ=BX"�! 8��5��{#�˲�-���7$6�'��GwY�u0���dt�WÛY�x6ɵ��������=꣌�*�rD��>Z&����k�����y
1]�Z_�ӝck��T��7=ly��}>���٫����ƌx{�S�э������z��k4��i6,�~J| hHo @����4�����p�&(%"�k��eޭ��m˂�Z*�U�䗃�S��p�q!\�@��n�$���o���2ڏ��ѕn��Jt�8��69��
ɛĈ�At�s�b���to���v�0j1>z�o����n��_&�}�σ�*l<����M2�#6Vj���ZR�GV��T�~{�z��UkY������t���T94��ŇK|�<.)�"��E�
y&(ͅ�w����*�;����	[�2Ӭ�CW8�|]�؉�~�lk�g��Q�9=H�V*�E{��6lBܘN�-eש%3�O8.tʑ��V
���53�e�1��8m� ��;s�,J�����c��Փ|��ķWjt�=ޮ��9x�jh>y�~^��j>�&�W��v��l��k��5�p���u3)H�k�]oӻg~�2�I�~+J�.���>'4�Ru�k���9^�"���+o�>x�Zz����c��/%���qi,z�nQ�v�n�7;B[=X�z�q�|�C�i�Wt#e����~Z�e>�>Qy(��*��.z}hp�N���bjz�|�{�Iv�������������ӎ�1����c��X������s7e*,�W���<���C��#}t" ����$��ڙzVE�{�J�;3�<_9��ڪ�" ��l(l�)��zk����)���j��U͉X�lҭ���X��� L�Q���v�'���=|�G'{��BB��n���(���W�H��k�8w8�kY�t�ٷ�N�d�3|�6E�O3X{�1��O����{�%O�B���?H��MMs�ڂ<Y�pw��\�I�<{���݄�S��fz�(˻��b*�j]w�,�s���)�nF���T�\=���5�P���
�)�կݸ?7�l���Al��\�Aַ�U3�˞�K���Yo/9����y��p����(){{*V�`No����<2��&���-��5ڲn�<&��nq��n8���L-sR�om��8�g�#5�ݮw���EI�m�iE�}1����������ݮw�5ߟ-h������e;��ϯ��ז0��M����7����.�4��c=��ݾ��D'��hՒ2�Ս�|��)�)��Ϋ:N�H;�O����އy��LA���gz�ՐJ�;�mF����E��k��Zx�Xٍ�[�.�2(+WAtI�qq.4Sk�O'&ʛIӴ�n8������g,!�:����U���1/� ��oYt���º�a�$���#�(�ӷ�YڱY;Y��6&yQ�{�
s��~Cx7,=��&e�$�=̎�q,,X�:�$ѫ���Q����mKb�3I6�g����쉧�ԡ��(|+�,B;Ve׌oW��Ԡ����M�q{�=��	���	ԹڙIG=�ޫ�ױ�G�*��Y 1uv\�U�|��%����M�-̈́�p����6��&�A*o�y�9�����{�(�~5��ɔ��u�j�O,c
|�N���V��c�rs5,��b��1�s�0�	��uP67��ݼa��&^�Y�sI�k��yq�̇�������F�! ���+��仔�(�*̳���h����;�M.qBҿ7����SBB�u>�N
m�MGv�˵��ņ�'_��Yw�ay��!�;*�T����Ϧ,��r�/��fgq�};��Fۘy��ЄSPG�)R؅L+�fq�J9LHݯ��K:����#{6_RJu�0���'FsU9�u�C`$�4M��@���*:Y���u���i�i���\/z�ѱF`��5�L��wvpL�$��uE��{��~���n˵I�] ��F��(8�A\�)��d���o}���ʋy9G��O_��bZ��s�2o׻�kj���w����P�W�����[�k+9�$�V15�z��9O}����F�ϐq��h��a��������''x�oH���ګzw�En�׼����~̥5�	(���zM��s&��F�9ľ�D�u%,�cJ%)���K����~[�{��c��' ��;gϾ�gV�Oã����9Y����il*)��t���j!���,X������W�k�mC=�Ϫ�[��5�ONP��1��\z5�~r��&�l=[�c���OYY4�yu���j���!ݾ�s|�|���mӕΨHבЛ��;�>*w���yb���un���'z{�:~��w�8����آ/+�:n�,��)��_�q�B��r�ܙ�U�s]=wQg�R��#b��UB�.��{jP��9�gi�J�؞Lؚ��������`���B(A��Ӛ��ɷ!9��_�y=�k!^�8��;�'<I��viH�n=��5��c,�ܗt�u�̹V��D�P|�K�Kħ=��n���O�X;�yy-��q-�;�jm\u�������u�ǻ�\�P��+�c��������e0�\�7��r3�+�l���?k-���[��׭ӊ���`��GDﺷ2�S��Sv�+��Cl�} �E�®M ��v��w�o1T�;u	�P:b
}dS��_�]Z�ۑ��,��g���s_^Wl1Y��b��I�U�Oܧ�![���^;S�[�R�e j��Ŗ{�wΫ��Wd�ӌ���cfScZPd>��ո\i�ڸ}�~�oi���R��S��g'��sy�V;�r���&����{A��s-;�k�#����vr�ixǴG�u�c���4p���X�r���������ĩ�N�9����j�����Wcvq����ɛ5���4SZ�Ѐ���v	Xn�m�M��p-�M�f�]�9��iNdj�.�eM�FPD*����39��Cy���Ի�cF@�l�Rm�����6 :��4��X�&"�>��!wC�R�ֆ	�4/� q.T�6P׊j�ek˱��iL�GueK�b!p��&+���-��$bl]49��d�kfO5u�
�|<��>�j�!9H�]B����F����iٴ��0��sA��9ᠶ�+��I��eǗ�ˀ�±[�Oo����`��S�^�/�ֲd��刯&c�/����;�����#ѹJB�n^��%ú:bƬ�Էy-��2Y�gI�Um�1a67�6�S2��R��s�.Z]�eCoiY��7����p雪Ys�0����.:���;]�O�R��e@J}S�Ox�x��Qu�6h�\��y� v��q�QǪ[���J=Ap�'��tU�p��0'�t�[EM�wH7���yVyq��{r˨�6-k�v�4�-2og.�Ц�t�ӛj5��S�#g}��SpA|�NX2|������T���%9T-�q��׋���r,�#lwk�À��V�PɄNT8z4��CN�h�bT��̟+�i%5�D+�/+к���{^�~�，^�	 ��ڻm��㩴C�qa�}�@j�f �h��K[�ld�չ�E�����bm�=`N_D+!�"1��HI{��^)�ݲ/)J��EB��
7�ӥG�gew+J��4�1����{I��d��&˷2��y����rU�+�ﲆFJ��c�lI�{n�r�K�1�ܵ$��$z@WoJu���N�����DR\쯌[Y}�!6�[���\*leby�}i�+�N�$����ړ��c��=1�ح��lܽ8�'ˡ�rj��]@�.�3
�!^�=LڏR�I��Z?M1��a��e�N�ސ(4�t�F�_eM];��0�7Rkj<��e�jC�0�kz�Wp���:[Oi�r��a�������CV�Tsk*��e)�R�s6��6���(l	4���>��%�ʽ≴3eܿ��5�DZ+�BW
���^�KFn��y�`���h4 �5����O0+s���:X��B6�O6 2ogV�Y�cf� *���E_Qۖ9��R�V��V3�wCA���;jZ�b�}�֨-u�tT�k�M:Y�vgm̹8ٽ�����-��b(L���2�/K��\�CW�������t�	����5��aw?�7/2�!ug�.�j'�`D�K/�MZ�W,+e,�)�i�s�z��v����T���Sf)���TӦI���d�r<<�)�L%u��`(2����X#�[B��-2*�d.iP6��a��`�m�m�jY�H���[�]C1UEEE-6��V��(䪑eJ�3U�a�J[f��䠱�e�4�R���kI��7h)�aP�C!Y��s
�B�UX�[X�T-�@X+�U��MB��
�r@��#H�S5��(�0V*)�PQeT��TUQH�#(��T�fE���r�������ZWjk\��*,P�VB�,6�EEP"ȤQH#̅b��B)9
��h���V,�)`���EU�X(E"��H,Ud�R(%
#h%�V(����� X���¡T`��X5�*A@F*1dQdTAm�(�Q�YTUX������˫��"��Jv�R�"���;y�c۸�M	�m�[�S����vd�Ђ�{d�Օ�{J���A�D��zE7s��{5	�����<�`�.��長�T����={�U�S'.��EO:�UϲT&a��κ��T&�hJg��e����n�Jђ�H�ޢ�~D'��/$+�,C���0w׉�o���+Ά!� �4`��3U��u<j�^��q^lу[���觗��;�q��:�<��%$��!\'��	Pz���Ҡ�O�m�I��Ĳ�L���]C�6x�IT�����*:o�y�����v���1��%$�9\:C��Y�yC7d'�_%]r$�9���c&�tW��yQ]8�\�N�켫�Mm.�xG3��V{y䅓M�K�+y�=�3ό�v���;YP������~n@#`����Al�l*�&�S�T��;:��V�Q=���e%O,C�vU��IJ� ��^��X����ݸ��h��t�H%��A�exf�4x[�jü��-����!�y;o��ŒAX�[F��q�
��G�A5��ʌX-��+ՙ�w�ʼ�g\��z�)��\�p���\%��Y��i���e����ę滄ޛ�6[r�������y˵Y���y���|Xt����78�U�O.N����y�F�)��;��r91v�zj�䙚m�iE����s�1���ٰ�!%+�g��G{쵔3���ԬaO؉i	�,_�7|���~)��^z���N�6H�<�������kPyJWEG��f�ѷ��vϜ��5���{G�Yڱ�D���lz�����V��fY�}�Ox�H���-/A}�E������a͝�0u_�E��3��Xb�G^�.��<Z�e�1�M�)=����X�6v�i簽17Ӳ��3��k&B���o>w�2�����ޫ�ױ�*�H��������]
��� �c�N4.�d��Hȷ6n��s��m���]�]�=wZ��M�|�N�Y����&T�J�:E�j�O1�ɤ��9{4$�����+��}[�-�-�:��Nx�8�VH��ށdmJu��-�KY�U��ܻ��PY�~n��	�8���އ#���='�V�����oRy6V+���>G�dg���*�9s����L�Yy�F��4Yv"rLr4j㯖��0��Z#|�\�U��3~�\�sw)��lj��1N��{y��ӊ���=��O�h���X&T�3$�MC:x���ɒ��3՞]�j���L�Ru>��`�t����s��kyN���9�iZ��PN�P���`�- ���KGe�Z\jm���E������7�
�sV[���ڠ�E�s�ѕ���j�N�J�Ʈ�w���Ưk����2���Hj��.�lHk���I����%��ԣ�G��~p��B� �����/
�v�ꚱ���X��:�R{��v�1v��层���[D���F��>P��mp�b�0=^+"��Wj�{�9y*t&�J*g �x[�9�
�X�g'5�&N�Tr2X��٨Ǵ���*�u�}?u���}���y�A��\ͪ���Y3�xx�o�E�c��j���fU֦��qEb�vU�D��Y��}W���ˑ=� ��5���ԗ��Ef����נh���}T�֏(�9����.�`���m��G�2�(Sꋝ
j�CGy���#�\*���;jH���m_2�$��wlЀRF�gK*�sP=��w����T0�y%�T6lZ��j�^P�zD}�ki7�M�԰��|���|�L��*�M�����	$�S�d��~X�L���ko�w�5P�=BP|�|����z�_���ُ�>^~ ��.��Ů�ۏ�c�L>�J	VGM�u+�d�F�FZ�Y���R*��j�������0������unI۞�Td��T94S��"߶�Wf��q������c�cR�SYm��t�}{��7І\�m�sю�O%ٜ��`�2}O�T=�a���~J�R��ji�����8��,�5�C��]�iZ��ݫt��>��֕dD��0��E*��|����}�*0�D&���~.ֺ��6y���J6�ɽ�]�����\ԭ�i�wB���o*m(k���<6:�b4��U�d�a�k�I�:3ko��z����;1j[N�D�ͦUdh��L��&�ξ���M�VIo9s���$����u�>���k4rj�63tYy�v�poB��+��8#rGؔ��q��y�͏Y��H�w���·�Z��"�ԧ���'9y/qP���.���k�g���I���z�[�ϟl`��8V��v�C�ȜcN�n�.���|�Tjw}��X��κ�ZÚx�&�튌gP:�*x�Btfdf�{��5�ؗg+��V����s������p��<���i�-k��l$����2���PU=؃���<��t6��a���x����Qy$��`������z��_.8:_:d�RR��ۧԝ�or_�L���}�+���m�����/�5���K���U�n��3��๨C�P�^��x>�$���)��U۷}x�ny�C¦������I�����|9;	�NRw��x��t��j�j�VX�l�8ߪ[9rdg'Q�|��a塌)M'~Q����ߓT=[Wv�����Nl��ٴ13g��
�j#`�}�×C�M�ކ]�j}�(p��8��V��1YnU�E^*Ofk��ɍc�%��l�R�c��5s�*�:�E!&� ��c4>�G|��q=�K�)T�/4-�(��5;6_g�Cj9ۙ�P�.�$��-,�U1����O3����2k�ો槨\XB��aE����I�7�
yԅ�M�K��X�L2oq�W1�ُ��fv�fV�[J��]?7>#`����o���1bp7���P��ھs]�l]r�^e��mߊ�R���|S�[�͗��E��[]����%:���\�|]���U�[%S�:
U㵡:ڛa�ʡ�5�rw1,H���:򽗹Y�]QC�fh6Ć�]ӆ����"-��nc��}6;}���ay��O2�糫��R��<�-!z�sjo_���0H��fJ�76�5D���$J��5d�խ�{�kT���c�A�I�P�Gn�[.z�9+�����m�x�߲1�Y�=�r��K��;����E��z7���ԧ����1�p/��Fp���.7'���{�q���YGFp�w@��n��]�|���*g� �*���n�QQ�w���+�a����@�ttZ}�eRu/,{w]�J���L�s+�Y&vP:��t�%��0�C.NZz�l��f]��ڮ7}Z'-i7.�n��$;:^�Ǔw���8�� ĊQu���g���^5<E��¡��e�1��t�4cg����D���|��%�u�"�1#y�RQ�SY�={`U�-�؃�E뉗׋,�t&7���vC�_$_"��M����vt���M������{a�x�n�y�;���A��:� ʞ'�0p��ځH&�vj�Ggb{�%H��S	T�s�U�so���!���+39o97"�3�R�o��1���y)�R�үL,~��t^>�k�O��"�.}g�G�bFPئ�������j۩�`�m��c#i���͙�#u�}��H:ԑy��8�{N�V
�%*�SA����u]���0z���H��4�[���PN��78�v����mF��9��HT�.��Z�vW�Ӭ�4I�G�ˁT�~]�loc9�u�vF�{�� �w���\-k��H'HꛁaV�L1I��{d��ӣap�&� S�z�ڬAJ��N�o��,�v�H�[i�ͳ���Jܕ�����J��g�`�%��H`�kE��\��d�^W�e�b�e���]\�]H�0vq�M�d���;���>���.�6x�	~>I;L��H�ۯ/��fn�l������:�o[^9r!<����q�]]v��%��F���*/4��	�Ҋ��g���s$B���w�1˼��,�F��q0;�����;�l�5�m��������n�q+s�Ru9S����"�꾙�aL�X���m�dce�_w*�Y{��nц݆މ�ڔV!ˍ{���o�}l�'��� ]�.:S��(����jd��;�d��_.nw��vF�檶q��v��n�2�{�X�ݛq�^9Ba�J	a�w=؍��r\�FvqkT�od.y�Z�m�I�
;;�ܑ0h��&V��\ԮZ$�{M�^�ʗ���ݿci�&z�cW���%����ϳ[��&m�EH99�8�aЫ��*�#rJѽ�x�ߌ1}�L��x0��Bb�V��韌�'���̝���c������tKBp��5�ݑ����HN]�Cd�Q$e�K�LM����v�¤.we��"�A?�����\��vg-}��c&�8�iXlaqN:���nwP����$�o�X�������-�z�}�Vvr�v��ZUM�
P�^�>�;z���u��f�󉅎�]}��>���0�<�z���$�x=D�#&�T��*�r}Ԗ��[������P�pn�sb�wyt�r�~�l�����s�؅n+��Gh�Ʉ�>�6j�5�^L��cn7k���vҩ���דb|҃/�0SX�	mZ�W~C��uH����O�~��r�~��w�ά��s���9��D�4%�E�{Y���I�U��R̸�Z�*w�R�ل�,J���}�V�z_XX�oe����۸-x�gx9Ml��*��o�d÷�*�V!�꾙[|�󦎤J���>ƌk�Ȏ^J""K�;f��*s�)��B�qXb���P�R�3��~GQOT4 h�J��<�F�tB�`�=�tۃ�iR������G\���A�7�ɅTM�LH��U($���`��7$�U{XCn��6w�^�'��3^��b4��Nb�KU��Vac/����oz:I`���cx������u)=��>����0U�@�=>�V�K���e���U����blh��s�
������=y���<��jo����p{1�f�f�[���GH�HÛ�&�);
;:�%��R'��)����c�����	���iwt7ɼ�a�X���N����+t��Y�rj�.YK�;ZJ~�{��үLw9�:������i13�xu�S<��gk�]ώVd?fu;�1�ן��F�/o<�MϏ%��͒i�.�VY�|����}۶��y)y�ן��F�HIGҢ��>�Θ=�5>7�qz�R
���+�:yp��T
PW"6O��Y'����n��r�.�;o��\�|Xt�5Qt��7
�q)`����@�	��#=C2��3�x�^�ԣ�I��bZQtL`�=�=e�����y6(�6�XF�b���6ټ���k���T�u�}�:}n5L��pS��h���h�m٩Z�����S6�3s3@�2U��:F8�3��Z��G�����YtM���"��9��u��5݊�YL�}2��Z *�?���(��wv��P��E��,�vT��ٷ�ك������Oe�B�'U�e�0�KB0S}���KzX|^�fnaW�+\:�蕱R���r\0��N�-ދ��[ 8@��F/.P��[|R�UrP�|������g}k4���I@�wE�M���Õ�^R��L��w�GZm�f��p��{����ݤ7^�W"5��í���ػʱ�G�=��,Ό�Ļ	���I��cY�?�ϯ�V�U��-��ANL+�Wg:�����=L�έW�管L���3I�2�*n�J��h��8�7V1�p_m�&��a1;����iD�g	G�*�CL_<z�iρ��%����X31]u+ݳ���x����;����Ԥ]�;�a���P�ך/"�R0�Z�Z�o.���'��;Q�F&�ivlV:נ�[<xW^%AR�镌�L���hՈ^�cq$������ˤ,��W���Ȑ=�Γ�^�Q�t�R��K�\���\�I2��%vu�XR�uc U��2��s16��%gQ��K%fY���Y��=i���
sw�F%����A�J�:��B��S�o��q�ݎ��
c�XF�� v�����:��qj���X;��kx �=٪뷢��4yZ����$���T�d�.�|]�s��Z�<�Wh���w((�T��;X%t�?[�VX�����bDDMf]B�?�V���F�� ��|������V)���mAJ�r^E�Ծ�n�^��"�W��m�[l7�-��;p������)kR�>H;3�mܨ�b_k:�Q@T�������3o��ψӹX�Hf��
�b�}�WU�M$R����#ov�/��N��
�R�:9�I��)uA�Y������0M�-�;�d�|�����)�o0�Ǖ�J̣x����*�����u�<l�~ߒ��$Q�]=�Y���,�hj98�6��f���
��PV �6�h[�Z���;�ҼZc@t�3�f7���j�#)�g0��J�ƴ3��[�m���:�y�mJo����T΍���V������*�g\��X�#�Ȫ�����	���VL��ӭ���)j���^�+�ʻ5�J��hqYx	��,��]b8�N���x����ז�Z���iه��R&P8�Ԙ����5�Q�Z��Lc}"f�7�V�x���[ݷtv0sr�f��Tәۖ�8K��[�͖�5��_-��4H3j����sb�fc�n���$K�!�D���k1�q7{ߜ��}�������8Ӕ=aR��YXTX
�",��������T� RE�`�H�� �)Z4`-VJ�$R�V�F�D�Jʔ���`��VT%dm �B��E��d�XAk"���
�(,,��Z��@�R����-P��J�R�1��Kmh���k�(�V�Ec-,��R��V,�Y
���PP���(V�EXB�AAUTPZ֡X:�(�!\$֙*H�V[@���kG6T��T���
�+����Y�UY�"�a����Ʉ�� �&B�*f���,�W"łŭPTqh�E��)�@X���b�Qa��T�����Q`�(�T�2I��`��-��5�r����Nvh綔������\��-�A-ڜf��`�u�4wk�듲^�	���MR`I�.��`"�g�y���}�~�VZ�鵣�����lEõ彽�r�����Mhא�
�ګQQ'�$UlJG)=��ymfx��n��mQ3�sot��5�OОнf��]�+}~�g(bf�S6pJq�ȩx�{u�So�3�`r���9w��̅�lZ�/M��s,NlT�c���Tm��@��ڙ�je���:�,{kT�c[Hޜ�Ϋu�sk���	��X�z�!#y�2���ɼK�^Ƹ��LOC6汦���3��{@L.�C��\�$_"ܦ�W9�����1�7�����jLհ�ԉ�y���`�i_�:}|=��t�����QvE� g��:z�r��`�6�K�j���nI�ߕwU��m����->�B���� ឪn��>�w��C}N�<���4G�^i!lȩ�ɨ��4�f��|,�ݺ��j�41)�����~t�o��I�f��m�d��xrr���{⯆�H���ǋ��\r���ݕ���9���v��d�|1�`1lJ�;X;})w8����>�)n˨r?,��}�v�;�% �iE;Go!�I;I�go�6n-����8�{J�����H���=8���Y�T���X]����{"�u�&���ޥ��Rt�i�V
����=4D���"�]Z�k��K#c�8�0�o�˚����juH�:A�۝]x��e��dX���ծjW"x����:����=~�P4OI��+�̠�ڋ�c kWCF6�P����
q{B���f��`5Xq�S����j��c!�h'L�j�K팰lt��1ep�6ra�Ȱ*[A��e8)�v-�b��y��kªzt��.�t(�4��k�H��Ca��_F�ΐ�-�[JQ�u}��F�&���da���Y�����c�s�#�~�j�5~r�_}�i��װ랞OZ�6�[��ܹ���SǦ2ctT�q`l��텚��5a/,�w�믝���u���x�[�Jf�e;�9��S��L�z�).:�Q3��]2��S2ۙWY7���b�锄Z&��O3jL��Xk�(�_4&�G-W $,u]�A��k���e]�c"\i��䬩�[�k󞞉o[��[�7>�2��oq�r���9���l��7����l�JBimJ�.�u���1vÛ�{��S��ʉ8f� SBq;��3����k�AZ�j���%��?6)�@n�lyޱ�W{IW����{���R��:9��e��g�6����H�x��^��
�D���B+y�r�4�;�;-�b�t�z:���$���ʿ3j{/�xDu(�I� H/�(��Z��!:D�ڛ�憙ʉ0�l0.$ϻ'�q�\�o‷�a`p�H�c�:¢J�aݞ�xaT���� �	~� �Ƞ*e�9}8j!(�9Pg�0k�E>t&U(�aa�ۻل��R���]�D�b	�B$��	A�c���95��x%�e����u9\��:���/��-}����M��@�x*XPAv�c�I�&f�B���r��8(��
�Cu��wk�<A�����G�x�����gOt����S=���=Iv�{j�}���|O�q��;��W1��@&�<�%�4q���*+�f��C��^�i�C�~>�3��Me��d)��df���%wQ`<�
p�:Ҋ�AƘ�-O�hU�y@�h׫<l����卶(C.�M�{�յbQU������Z.�v�[����8?-�^�A��9r�`�s4�M��_c��6H͵�^�x�R�wH=�ꮔ��p��&�~���4�wztVӇx���N�ǣms�T��v[BJW�y�e�v���T�Ѽ�����`],Qg
Jj�}�7o����at�/��מF�=����z�5�Ә��~�Dt�������O������mM��ob�f�hQ�'�}Fs"�0�%M����w�x;�gwR��j�ǉȥȞҒ~ʔ:Vm�
���%�dUM����pt+�k��7�3�$;<n��Ԭ�SP]o<y����s���U{V ��C�ι���hc0��pT��Z��->mg@��'�.�ܮN�r��c�P�p�I��\�p+����Fs�'��cp�1":QMLN\�Xu�է��G,�0�h<�}�.+8*��}ŻN�qn��\uޛ�9v�	�rSm��o=�(�y<��0`la,�G�T�k�%6����9����# &���k"��u��;%�>[6�Y�>��HD�7L�9J&#��Uz����U�q�E��w��"y^�Z�� �;�Y�}A�cʇ�R�;�"MF�8�B8)�!�r�+7]`�q�7͛�R�khK\U^�'��P�7�+�
�um��[���PjoF�/Mpܓ@�D�M������Bz�R�ާO�Ć�<�f ��up���R�Ġj^�XJշ�����n�L�'�}�rQ�ģ��%$�j8�mv��30��?z�Ǳ�Ν�c�fM�1��s��[� aT{�_V=g�q=Ѻ��/a��7�9�c���*��(�s��͛:��Ӓ�-��E�B���)�"	ܓo���
gk�aLM~��{$�f�b��!�rr�!�"�qU�s6�6Uas��0�iFڷ���Q�K3�%�U���iۅ���u$P�� ��8���ډ�tg�S.卂�a7X�8�P8�7+��.����7�|p��Lpԝ�c�~���߇1����:\^^�B
2�c�h��@7�	�d-�#���鞳�+uj�</���z�$�����n����V���$K+�h&�\��Y���mGP3 B��<�"�� ���{�c&��SgpoC����j$����硫��+�'��:v#hҲ/��H5�zH.�=��ݤ�28�1n!؟p1|���*��Q%�Q�<��|3�{�Y�7%��ӡ��|,��Jsٺi��UԺ��to�BA��\�U4B6s���&�"gw"a���<k�=�td�Y��f��,�HH#���wv臻�^v�Q�ۋ�l�ue�G"�;i��7{�i��>͵^)x P���$해��Ǫ�9���n�F�uZ63�	zi���,N��_H�I5�^��ܳ��9�,��$��tl����6g��ꁭ���SK�D��
�?z��](3�C�j��7�ƅ����b�U�-|��*Q��E�,�qb�DD�����+����H�wlhR������q��V��ݯyٹW	�J��j�x*���X���'��VPG��*�4��g蠛�������kPCٺGNs��E�����'C}v�{X��W��JciU�I�g�p�%Z�L/�7z7�zWއQ$q�r3�9+sЧn�@�+j��{���1��HP�Q;��9V�o1��@ч�/.I]����	�Q�C�!(�s���r����s��E=�]�k!j�aC��<�� % �qƆ!�a�o�u���C7mC�C�ZWEcPs^K����O�5��Q�i��5�0R&��E�5�d���;�J�G�$�]%���}(e�{���13ݱ��B].ۚ��l5��-D���2�b�67'���]BC�2�>�yoov�Z���Dqcw��,(d���tɠӢ>U��r��~Kh1۔x\(r��J�a���NhŊ����.���=���٨�:n�x�}�5lb��sI�h��RV�3��m��tVw�VP��E��=�ƣ�ɠ�.A��Eb\z>������g-�3��o�ˆ#0GC���;������WWX�6�ɀ5���&��ݷP�3�c�ҿo;�,-tK�"J3��&�R"�if�W睝�N���"��0�NQ��է���R,�5��fV�]�L}�c��������ӎ4t78`�]V�IdIh�fc��◉�1�-X�ճ������Q������:�sDR5y�hb*c���m��g�RYJ�Øz��x����*6kb�JK�����T8���B�+.Sq<���s�&v��DtQ�����ڰ?1[Zk��Kt~lQ��Hz��{HD�f�N���fݕ��݀�J*®�^z#���=���!t\Kꃳ|򏰫q��q��ê���'M����:IE��ʿ3j{/�@�Gr�bq ��'l�3E��,諭?�Xg�gި�q~��2�L�O�\:�}�y­#�1�=9\�n2�f6�)b)��L�@Ԥ`��Nr�pЈJ8�T�\�$S�b{�ވ37T��~�r�a�n���~�*�'d�Pk�=� G0z��/%�e���<2���S��~�]�¬$$�Co�M,6�Ձ��M>Z��(]�JCo0�(�o4,�BP�N�L���)X�Vs(�m�D��t�^�9���Rֶp؍
��6��Ȝʔ��O�C#��i2>���:p��&�����:�N�i(\K�~���DT��p2
����;&9Ě��,א����ǔ�rk%#��W��m���[N)Q	�Uy;�}p����/�(��AP���.��5�Ov��L�n9���yOqs���+f1�őA7\a�t�q��C!B�s7�&��g�3��� *�97��*#,��3��CH��(;�wP0�x',�҉��4#ܾ��a��~��{�K�>��az����V�o�K����@߀xjt�]E�� &��:�^���vD.ؾ�XV)�}gK���g+�9ypR��B���R ��מP������e�6,$dY�c����fUɵד,�eI�̈*�ޕ6c2Q;��6���6@2�^,{���Ҩ����Q%r�b�̙4:7>7#�x�Pu[Q�]z�Q�a�w��X��Xu� ڥI�:����w�4��p>]r{-Y<�'jj���A�0��:�8L\1P��chq���;�y���S����5���tnz�D\j�jc�=����[��-׎�R'�}7J�;cre;�e��)S�8�z���]���窥Xr�u�+�k���k4�����{�_H�p�ժ�\je�kq���a��E>��xrq7�e�]������@��!o&*��$
	�Ɯ��K��T�V�R?�EL�)Fq��
��d��v�����Q���g/Oc����9}޷�k���Ѥ��⮦H�4�H���x���Y�-�]c�������#�N;:J�o*q�D'��<I `7I|��i}����ᚡ}+Qr����<�D����iQد\q�(��"��eC��
U;�"MF�8�s���9�8JxV�����&�H~��Y�/!�js�xc�fM�cj����d�ޙ`� ŞC{2tW��)��6��
�o�,V]N�N҂��@��
t�9�e�$�AO�Sv�z�o���ː�&yLՁR�6�I���c�1A9}�CYU�7U� '}��F��C����x4|�����.S^ӂUe�Û�$w����Jq�g����V�����GfE��d��kUas:�3GM����R��2����`���X���8v͡{�WkS5혻�X�+��lt�xl�����~�Y��G� �	�-�B��S�4H9y} �+�{ϔב�_��*J�:N]�V�
������`$��]�f��oM<��] k����
���cF�`+�\�2u��·Qz�pSˢy�u�!����ة��6ѻ7���U��=�"�ѻ��s�:"�q�^�*(��:�F7i_�I�򼦓X	�s[�f�Fdo́BT��&B�����"�o9��v����#X�b��t�:$���t�=j��k����VL,�b6�iY�`htK���҉�[��⸆�`��������Y���E�%��d���9V^�O�f�L�m��]��Q�R���
��|�&+��5���V{��5�g3�y��ם\.�YV}�����������MI#��>r/��j8�r�f��e�^jf�Wjk"��!��H�
8�E�ܲ#�}L�&�׶�$+����M��
t�\�gX�W�{:Ty�	�!��ST���V�s`aQQ�$h2!�b�j\�Aβ�%�����g���+Á�=L��佑�	e�i���"Ʊ;�G�R"F��{;�5�U4w^5��l`#c:�#zZ�B9+pS�7u;bڑA{����N�S�P��¬�Ɩu�I���N{�+�����_�:J2�	Fs��������Iᮭ��נ��3oo>�o��c]�M���H)��cY Vtf_ut{�%7����m�رӲ,�8{�
�&���4����}Ճigut�d���fⓤup�KAUԲ�����kWWb��+jT�u�� r-�X_>����_�i�iJ�5e�,p�D_oH�oC�N-S��Ŋ�WX���.�vB�M1`��gsp	�S��.�Fevm��^��Ny��έ�/�]V�� �@��(���wF�vDv,6d�k5��ܭ�=4G-��GN��fb��nr@���gu�p=l�'�̻E�c�$�SD�c�	��*�p}�/P�<��҄�Ww*�;.s�Y�f�hDGXN*�V�	۩�OK M��u��^����9
z�*I�K]����nW�ԆJ.�<C��	�ȘBc:��ׁeA�^<�˶m��d[B��`<�u��)��i�P���zr_`C�_a�ĝ:���(CqӬRm�j�j�R�N�9n��ب������51b��V^�C��Ym�kC���E��n�Y��̶a�BTa
dWM�k��+�ѩgn�t��V���+�Kv����r�5�V��M9t���gCְ��j7�_ӏ7g��X
6_b�-uӺڮ�C�9u������hZ$�'*�Ht��%�qNQ��8+Fn�r����O��S�G}}����WU��U:��$�\�Z�7V��܁lw�k̚XF��f�M��/�2v^�zQ�-􋢲7_dzX�1���r8�g�S��ݾ�M�V��˃z�zzŗ\�Ŵ�a��w�힥�Q�鉸����vA�'pM��z�^�7cnv�"�MB�(�h_d��-@�����n�Kp�]x[�ɲ��j��RЭ���g��R���`1}�D��L�ˡ�� __t��*�*���J�X�WS�ʓOwjt�'��Z�#4�Z�U�t�����Q.ZB��'�b�];�WV���L�R#Kp���eA|�\���7�Y��U���\('4750BŽJ%6��U�������IZs9l���p���X���aD=�M��ʌ%#�9�O�b��]�ě�;oe��ܙ��Y��4��@����t�������LJ�+��^ނÒ��֒o��;��[w��t����+����d�ܧ�s�{*{�NE��\q��|��n�ؘ�ڇ"�A�&�ٗ�vj&�l�<9Nm9����И0�xU�Q�U�Y����n릓Y���Rޣ�;YL�;w���jn��ºD��O������*\<k��R���}�0��2��۬s�h��z���=Ͷ��t�j���v��܈��J�C������O�q�t!���U�K��Jj��4p���JĨ�i���0/L���m�F��������������TSZT�*aF]��T�T�2f)Z�s����F
)�V��ʂ�XdѩRV�ł��B�WZ%#h�a�ͭ&��QQV���\QZTm�����R,��Q��UA@XVeDeC"0ʒ�u����K5&A�P�@F�,��sb0�+KhUEF�*��TaZ�4�Zdiau6�em�rW"3[���Q�eB��
6ʮm��V����*�%J����@�X��d*((��(�,6�2ա��"��,�X.ڴH(�B԰E5
�m+��PdX"��Y�e���Ean�X�>�'�#�<O�	"��٭����J��s�gR��У�R�wk�%Y��4p��c�I�l.ЗM4���.���ƹA�n��RI��l`��B]A1��u0Z�$�#�	�G0_E�0R�[(8C3uw1hDC쩍���瞵.m��UO}��x�וӤ�Gt���#ad�!vN���+vT���=Gӝ
oW.��*�K1ӈX�'�tP��g �[na#���
��0�N.�kK�wZ�F9�3�����"����XiU�_�2TM'L�P���2��Ӎ-��pA�x,�����-so����è�7lm�F��;��"ֺ%պQ�	�&����1Ĉs�i�o\i��^k�28����t�AV,o�^^�Y��c��s�#����k��6g*a¢�t~�?s��}%%:���ýY���tj��Mh�9+Q����Q[��}��:+=�:�Q�#3܊7D==�q��X'&��t�¹����x쥲�~3��^�ۘ�W�ը��G}�v�{U\��2��&�N��Llz��=!H�]��rt��w����m��g	�:���hb����R��Zx�m�����$G��+�=ANWD݈I�!N�]�H�t��B5Q�w���)�U0�Ԏ�u`��Ϩ�<���/Q�j�p�i����B���Q�ى�
N������X�pp�!��x�VNk�%�L5�דf���،����̾����r̋��:�mԚ��satv����
B�֐�6�14���:�r���
{/�Dr�b(t���r��r�ec�\�2@~7�z�_E��p�`��#�x���:ž�	8Oz�Аe�]�57=��}���[ �:<L�D�ґB�y9�_N�BQ�3�{�\���:��ڭ��U�H�oO���)��Ί�����Q�95��y�-�,�Z�;����{�����<��CM�dF�{v�`���E� � �;&9Ě�E�]�s��`��nb��Vj�=�^V�D�*!�*����Q�5���9��>
�5�������^� ��g<���r�m�#�M�x]2\q�GuA�~����I��GUr��܆�v�b��r����H㕗A�^�{a`I]�<�',���Y"�6,������N��}��>��P:[�_�u�	��ýV+�w;��],Qg
`IW��ꙃQ3N�+j{sI}��"n<�����W�B��l�Ә��]��� �
Ok�*k�=�/}���vy�o:��7���Yc�7��̄��/��v3��a��g2��,VXύ��v���<zl-].�ةWIz�t��$w�
�3nRS��];�2�9��1 g2	������jl5���p�����*tD5��4#rGؔ��/R�#p^頖y��s�г
,��!�x�dP�Y��E�;.��fS7����M)Lt=xXڪo���sϦ�X<��̜��B�p��k����8�s��3�o��)\A`\a3�t� �S��U{V �����z��q��~s'^+�k5[c}�u>�;7=}��4F�GQB�A]{A� dI�S�'���S����g�뭘�8�v��i�*���o;7�0�I���Y�dA��8��C'�[�����J!��nm��A{��oR��s��u{J�ӀA壑"�^�H�=>�O��E��T��s������2�����,]��(��/���(Q �;�����3���5vrs����m�|�ﳡd"�w;Eo��ءqǈ��PdX�2�Ň�D���Q��*�U(�X��uþJ�pE�N�@C���y���1ݳ&�"�x�a��A؉�ۤ.o���G����׳�A�;J2�C8YÆ��zs�]e����
�;>q|�C��(�["�]���U���!�g	8��3��ub�Wn���K��NF�;�n�Op��S�����5c��x�;^�y�L��$�юo��J��q�w5ˊ��D��N����S0E�V42el͎��s.�kr?�pܜ���` �kǦX�'��5`T���l��ؐ�T�'/�r-�P,ʞ��#fcV�����mr؇;XT����T���\k�pJ�]�}��<�tC�]�Y�{�S��Oҕ����o,��2�)��=�#��W��`�R=��<}���0�A�F�?Wqǭ7(s���l0��iX4W9 �{|vB�20ҡ�7f3�|
={�v�\�|{�8t�"�0�*w�<��"i�yM�hw�2�w�����n�:8}�n��!�s�'�;+�z���=G�<�DuK��+b�]3�|���מ+��ag�t��W����]����3�-�U��1�#�����Ćx�E�N�k�߬7Dt����5��2�nר�9�uTـ�<#y�8SB1�G9>�r{=}j�%@��#og�V�l�`��a�M/�����
��<�3x�x���[��n`�|��IE�t�G��pnY��D�� 	
��In�M���KX�3M�1��v˗��>��j�v�����G�k*�nsB/ �yVF�U�Ks
���@���J�ͣ�6��l�Au�\a�~���4�.����;jQW���s��ث�sH6�wzby����,�����[�3F�Sp��q�b�Չv!d1Y'c�-�J�j�x�V�s`ah(Q�$h3�')�a� �r�W�7�6��U�$�=�@��e�佑x�BG4�p/V��+>�!�v#�37�e?T5�vzAe�躉#	N��q*-�g*!�j��%Ad"��`�k*�%����ir��I$�>�6
T cS��rJ�]\E�N���J0C��-������r8�}�U��f6+�B���;�	�9���8`��`���AC��3
o5������F�_�âd��/|�ָ,H��W/4gad�!vN��E��R���u[�ڨ�V̝b0�D���<.@��(]�5; ����4�
V���gI�S �ࢮy�n��t'C���f�Uu2TJr��>tG��1��<�mn;�ػ�N��mc��6`�s^D�!恴Eur���ȵ��un�e5D�R"�Y��z&e��y�ܻ3�`�9�v4��gpT�#�q@f^�Y��c�N~|l���y֫�?xs
!ygi�q׺x������KV�'���#����r]����N�HN%�
n��q]�4n�Tcv3	�}���E�(9�I9+�nn�H�<d�r�.���HzÕ��4q�_��7��3P̃T��G��%m��PvD�ŲŏUڰG�ܫ��D׆�j�#h�.��e-���*=�s+w�}o�]�'�N쭆;��X��23 aJ2#(���Ġxc�<vb���z���jyz��bcrВ*#;dt̤��Qg�u�Oj�p��m�U҉�]�?6(��:���w)b�\��IYs'�E�41H�©EZ��^Dta�m��=���<B��4i��!���W1�hk�X��Cȃ��uf�]�ݹW�mOe��w�����1zܿ{�e�M^�@TKQu�(ˉ2d�n3\�qȿclT(��縇�=ȯl��^j���� ��-Z)
�r��K{��	�s=ʃ=��4�9Ǧ�E���Z��0���؛���P��!�Or�I;&�@ǹ���Z����/N�0e(X��j�6_�-C;���^�/n����E� �&	�9Ě��,���͝�{��]��tɉ��$�En�C�`YT�g�m��اQ`(����9�1� �Fu�:�t��u5H��2%Y&b����oc�,81��2� ��[��՜�c�A�hR��g�m8/6X!��`!���2j6�������F�a�
~��e�kj�\��V�w��J��GH�{)��lbj��*C'uol�ĥL���Wb�W�����\wC!7<a��Nx����do�M���Z�(CN:5;x�_fY��b٩�Zj`3y�AC5텉+�0X�w���(����5F�2�c�9��u�
��>G��4%�i��J�f�7$a��8B��wы����{��c6�FF��׆�}W]�n�[�6���ض���ɾ8l�M9�c�:Du�qC/��N�g:m�Wb��+�`��U�Ft!�aE���=�>�g2*ad2.Tٌ�e
3�d[��;L�D��l��da��C�8�h���qӇwfN_��rA�׈}Iv�In6�E_Z�X���F8�����}o��q�uU�X����-����'��"�L�<�s���xĲ;%nK��,R'�c���UC�������3���N+��)�dn�vzT��'�a��klb�N�D��Ac�@�a��>�������k����㰘�!19�>^�s��(u3�����T<�r$V��k��
#UT�N���bJ#��C:����z�8�\Eb�0����L.��خ�y��[oOJ��՟_�mz��˹�m�9F�.�x�N��ҞAd�b�c ӆ]��,亙ٌ-E���fá|�Yswz*��2�n=��
*y]%��ђA�N�p�)��F�E��ϑ��V0,�7��I#(��4חqD���)哻g��ԭ�WݬA� �Fti�suǵ�p��!����c*�#D��#uQj�׶ys`'�W�竲��=��c�����N�ж��6&6�n|\PpAM�v�/66����y���16����`*��(./�͛-;v.e�8��.c+����ĞJ�I
��zX�'GF��S���HfE��`r��q�'�<���n���˵�1=�fn���/�r�63Ч��`�!��u�X�ӆ��_��I᫨A+M�t��C����12�b���ڊ~�00�V��Mx*H�Z�|�z��P���1V5�Q�m�����.E1�J⍽�)��r���Mu�@6��`-xw�����*^X�'�}��m�xA�{�B�����ΉO+�i5��j��K�Ta�b�ɜ�[\�w�Hu�@`NHf�B���	�]H��tI{9K<�>�>�y���naD�8]��J+Lq�wF���N�}��f�/-^�O�gk��&��V�;CR�"gBWy�7Ee4�]p2��/F>%�w�N�n����Iu�-��|��Єq�A,VF��9]����
V)��S6���3����mI}��3�w��vJ>X)Ҋ��M���y�֊�JF'#�����K\���G��y����GٻJ���6�1�Ƽ�ƪ�����#y�8aF�p%R�(����}�TLƑ��!(i����'#.2#h%�#�����A������hD{f�s��
�qgv��q~t�aG�n`�<vB�d�53/����a�uf�[X�Z��7�eI���|'�<FBj�x�ZQ�,�<(���5e^�X����fƤ�k�-�tHf�gO,���Y��PJbGM��:�dB���o&�"��U�7�~X�� ��q�C5-�<�{G)���9
ڡ���<�N�_(�st�\���[�v#��$�@�*q��G{9�p�%Ő�xlq�%�O���ϭI����/|�$>/�H� (Ь�H��P�i����?bؚN��t�;�5ڗ`�B7mE�t2���8��	4����#J,ɰBܜ���\�Q�;h������m	������{{�8���K,[�ژQѓZ�+�3K]g���W�iB���V:�� ~������m��u�)v*J�)�f�K���[�R����y))d��tU�r�� S�#�%Y�͎�hJA��2vn���1*랠P��\I�J�C� O��v�����Ũ�;P]V����mĮ����+��4F[��f�Uu�h�A�y�V^��j�u@�@oqL��#��xXt��ٌ�W;Uк⮕��dZ�D�s�a>�J���P|ü47W\�V��!@b�p�:sѓ���L�PU�g|]]�](�G����xX���fV`h��77�&�p���#�Պ�m2k�X�a�3�%5��������9�<x����b[Gt9��d�7^��T��H�,U�3��y���,��f�l]Cq�ɂ.M�{!�r���P��]eB�\�p
����Q�	����N��
��\��+5�F0�i������2նlܐ�.I�c(t�QPM{��p,*�R��x��<m��'��H�ޖ6�,]z�%2{sz�����U�H���GW�d�B�:��%�`'A�r��ږC��|��������=����1��P�5ΙZ+�t�B��^���S�TP�CGT����n��\��F���QZ�DC����1�Vs[�*)imd��lW*q�Ώ�e�FY��k�W'DV��J���ˢ7-R��$P��N��RFJ窍f�3�7�[�4�r&.��T�>�����/B�jN���K�7�D�0�_qӗssR�z�t�d).��8ɹ�5��ד2����*���+����d�Έ΍)2�A���O��5�����t������Y:��1]L�9���ub�J��� ���j��UEgݒ�T5�,� �;�9{�� ־yx�r}���p8N��IVF�Q���U�i�-���n���8+)�y[!	T�nh�jR]]C9��fb+��'�����D�E��뮥<���rQ���2��Xrc�B�V���od�Nk��t&�S*�h������.ܼ㪤��Gpq��I��6q�J/2����E�̗��<�G/�Bt$�u{��Vj�7��*�$^���u���Z��-��g�_���ɑ����:��;�@,n�n��t�]��jT�NZ�ѥ���w�i��{5�F�;Hob}�����L�na�N������1�F�b�>49+�����f�$T&R$vc��:���
b��o_L\ �C���qq��0��������]L�OV��摔�sكw;�t��t�����s�U�,"��4��# ���;Mf�z8�s��.���C��r��V�@�a�k�3;��4�te'%ee�>ݨ���M�E�cIM��	��z�5���
V�;Y�E����;m�Y�z��42	�obI�2�;ɘ��:�T����p�V�M�j�������t��Q7�0Lڝ)ma����ȵ탳����èe���r�
���1:�]�ж�Ԟ�0kW�+��oj��b�2j{X�ӑ�W>e���H�ݛ'&q�Mt(lj��t�a��+^D6.[y��� h�O3E�9�8\ͺd�C�z%��Ů�����:�J�L�x�KY�}��c�ъ	�(L�z�q4�2Μ"��U�G���5&�Y��H���.Xz�8��!���dm���]K��j��s�x
�����D�9\mt�(*l3�rB܂�W��c��;��C^�Ӥ�M�|�l�QowD{xԧ�r!Yy�(�Jّ����7%�eD�_`Y�'LQΘur�VR�5K;cS�;����e�5M��w8�Of.�&�V(��g6�I#4*��8��U��@���g;:)���ް�efgaRh1�ʃ��!�xZ���;�U��!�����ɕx4�<tΡ}�M�W��z�f��̴h12�V"�Wpp9�h���]tV���c#���O�rܻT">suqd��*�LF���QYj�危#�08�Wq�:%oU�l��O�l?�檪�QAk�-�����2�V�J�Tb*��E�PV���b�
	��Qb����m�b�CQJ"��78m֕b���X�B��u�QJZ-eEDPԱSYl(��AfeiQYnj�l�J7[�b,A��k+.��G�
�K��ZE���TDu"�jd�L2]�ثR
,5�n�2R+%E��b����*�&kV�h1X�P��VѦ�(�b92m�Ee�)
��+*�v����h�RjR�Ym��I3�XƲ�*)]J�s�S"�Psb�s�F,G9�n��Y��°�fQQ΍J�!PveU��¨3#���b"1�\L��~��Y������P��^�ƻu��*.�aU�$�|��m�O��H�J����2��|�3�s]F�3 ��8��2��d�F1c����g��`qiH��q��/���Y��72?X��C�Ivuг����K�F��Cpr ��JU6A���1�q@��b�U���|��]٬M),Gm2�D[�w����,���D5baB
!H0Nόs��f��cw:$���K2�1{En��{�*j.9���WzO�)�S���҉���4�M�,�ZŠK\�
��B{}{0��d&�4]Nx��M�}�b�''�-�a�����Oin+��6�&.���U�n��<�ݻ#2�q�r�92fC�QݸK�T��Sۑ!�3�W�P^g��f�N����ܑ�:,����b5H|���LL̓�(#��kϺ�"��<N�[�+�G�=�؅-w�yzש^�c���Q�y.��C���n�]k�f�U�} �y����i|>�ѐ���V�5�l�q����VY�c(n[�,�UT4��!�}4]�W��2r���HG���ă�b$�����������~7�i�w��s<��"o�=i�7��}��W�b�ʏ=�����	.�l{�������+Zz�-dw�U�U��Ut�;�aƶ��J��,�L�7(�[}(�����kN�T��vpގ%*������^N}K�_�]'f}���qZ����Y�p�?_���,�{{�/�+�
��2����H�w��3��\�Lf-��^�X!c8w�ǰ���ҟ)>�fy�9u#O���h״�]CB�� �O�m�'8�GI�����sS��Y�)Y�[_v�OU{�iB|�
��+EL�ƦJl�Wj##��M����*�����EC;��y4�<
$a��Bp�Ӥ��' @�M:^]�����[9�[)W\�\��9�T���7\{=���x��C#�1�vč����ɢ�
���jDNŨ�8�NQ�� W#;���ճ&�6�n|\Z𵁸���Y���C�t�HH[Y��NҌ�:��5�����"�#�_d�ܼJ�m�,� �~_rd������>���7�c�h'/�(��\w���[�ۘ�<R�l5�=[�ߍ�V<�}�G眳ţ���|fo�M�5���p�]�̋
�'��)�YF��Ըc}ʯ+��ɧ4��j��2AwOO���c�é�wn���>��[O1����76D��ԥ��ž}�0b�Ld�ֺ@��h��OWz�\�p�VU���Cy�\��c�$��
��Zbq�.X�w	D��i�0��d�j���!�Mr}`J����$��VB�#{��dj��
�kӼ3�yo�s�{X4Ҡh5�9 �R	�d-� Ep�����ڵ���2zY����v#���
��\
��N��rH�s�X	�k.���q
��v;cr����,"A�Ĺ�LE]���t8ߺ$����o�O�׋MXk���t��{	�� ���ҾG��T��,�QV����A�>��oT�S6�je�醴�X��v��NE����b�ԷhU<7�,�u�:z�R�:�@}P#��r�,lqiWU(�����\j�V����ێp:�w�Z�*��d��JG�:'��["�S�T�H�����z�ױ�V�hB)�3i�qn�",(�ܲ �舿����#�U�c1���?w�J�|t��}P��#/���_	����"�B�(�GP�!�(B�\�_^�A! �͠��ӓ2�,�����s���/����47�lĩ�9%��+��pΗ؊�&�̃�U5S���+F��E����*g�Z��M�8m��a�c&����&�a�v�Z��]��XԢ`�<�ҵ_:��B��:��I6�0�e�]���{y��S���7�⤙+e�Jh�y���w,�hɀ�$��:+�ye.�4�j~�� �.{��Q$3R�
�J�c���N�ظ��:��>���̮��w4r��o��_�s�ܒHR= l� Ƹ�$��g:�.�3=��]lBsӎ��w�Ӳp�V�M�_]�*�aF�%*2H��b>�+��4��{X�|���dhJ����h�.G��C�P�H��m�a�S�$Gt�
��xx /����K�iyN����M�_�p��rh:�MrT� O��E�洃me���!V~fsr��B#�^��h_D�`K��D>���f�!�J����k�:d�T �|�W��{2�ɯ)�рS�����^qZ!�9�9�%�$+� �\�cyݑ~Z�V���XI=TfI�P܌��ZUو�;$E���Pt�8k�Θ˪j�����~'���$�=���v��ɓ��s���Oh#d�aO>n`#�*�xmC�<r|֏��UW�y�MpOe�Y(��骏�v�%Ψ�戠*�����b�+�e��&l��JysCkeV�	E��n"[p�g˔�t�k 9ٞ[Qy��L���YV�G�]��̢�u`����SgS�c]Z�7�#�Q	g�M�fk�(u�-�;zPt�U���m�:�Y*�$FM�޸�?6��>��M��c̺X�V#D��p�;�H1�"�J7�&F:GD>r9USQ��z�n���Ӧ6=Dv `*bk(\C�*�]������R�"�d�ה�QPMr���EpU�͗ч������l��:똝�N�極��!l1#*b{b���GVL�j�:��%�i�nܫ�.�z�{�ї�j��Ś�GW+E��ȅA�1�@/�*��51.;�.$�ܖ[��%�� i�w�\p��H�A&��%�W��ZF1c�P*	�$�Q)��+f�;VWsbxs�C|�m=���V�wa�rH�S�M�چ��AJU4��=�P�u�k�j�s��)�V��<r"�3�����/nȱ�T(����'k�XuU�GL�R\�gvr	)�O<Y���*j�s�ʠ��>�sn��RE��&t;���%��}ilTGP�K�g�(T-�C 'B��`"�	��	�Aל�fox���\K��V�9R����d�L���8�;��ϩ��q�
uW�uӷdx>�oٗ�)���i��5.���C.�.�M��Xg8��:�h�`[����{6���a�����[feg�e��0+$���f�]�̊���[b �EϮ�6wLK@j�Z�I8i5��b��BwXƹ��[Ltk�B㑠u��ԎuĜ3 ө4���U�O�d?s�����_����z��(�7P�8A��,�r�zSIv_j�/۲�u��HMQ4uNE�|���+��R�0�-�����$�V߮5��}�6t����|�>���e�J*��-г
,l8�'Ϥ��O@;|D�9�o�;�!ԣ&���x�9j���da��C�8�h�z�Nى�ʀ�z�t�5����_r��
�X�n�g<HU�T��55y���ϱrw�+U�;�s�"��MmZ}hv*��{'"4"�:B�FL� ^߆U:�9N������7*Z��XI�o��(�A<%�J!�3N���j�n=�׺�i��h��x̭T�gMuHf/	ݻ���O��{������ڽ�jWD��5VW��Ɛ��r��=��C6��^����&Ԭ�c�P�J�_�֏�~���u����Bp�Ӥ����4��Y�k��
�{W���һ��ϟ]P���9��ٮ��<x���ȼc*( �9$4T����T��u�p��ڐi��S��Y�5��d8pޞhq����E߬5V��v×:�42�-���#$R����D�'��*w!��Ѭ��vt'�.I��\?dТ��4C��ɷ��|��eB/P�9�ۚ�kR
�
$ȇ+��P�JY�g���7t6��fL�F$Ѫ����;�\���\T�`�� �0t����`*��!�t#�,��59�H��}.��k|z��~�Y|I�HJ<WJ�'W��mnO�^�]t�u��Ut5fҫq���֑��݈�����C�������c�0�s�U���q��~̊�ذZ��_�I�׺�r[u�胪9D��Pˇ00�V1c�3'M�[��R��v�`���m��u�%��$foV�*wm��LRr��Ҡk�u�@6�zN�[�Q"1����|��]<��cO��*�P�ҍ�	��֔��"h<�)���Mk.��̾��-X�(姝��d(�fd���D]��+r�q��%�X�,��������ߺ-0�/C�����sƦ��p���ٹhq@�k�T���`Iߔ��.ّM����,;O�Uk�pxJ�س����ͪ�y`�|�o�@}�[�N7e�d���t��S[n. ���M;��sȿ�+��v�wc��N���l`�%a2�5��$���)B��V���9i�w��酰�-������<;�6�S�N]��cj�<�'��MPUꬳ�ڤ2�9̀w'�ctuņ9H+n1]��&D���U��*�!Q�&���VD�e���kD`�/�}�yukfy��Κ���Բ�)��d�
��[�e9n�H�Q�:-�dA��gd-9�5
�s�~ܜ�^r�ˣy��z���u����<��2���"�(U����8����V�^A�����4�|m��:�U�	�G�u��T�89/d^9%Ї��(]��a�s0ݚU�V�g9Sשq`.���)#A� �s��Q$3R�
�J�`r�q�5Dpؼ��T�q�ם�V������A��)E��b��$�0ǊT�u$���\}To ���9�5ڻ�l��ns"ӷbn_]�`��aE�^2H����s�e�n��M��}o�g��Q��p�9+eg�r8�nڋN�e����8(I�3+�x���޾sV�9���XF/�k��4��rh:�MJ�C��	k���sZA�5��0Y;xdSY:^���7{:�ˮ��k5�~2{�J0����EwMT/(Dד�M5B��9מ�tL�a,�e$E�$�t �6��ʹ�[vޢ�%��)M�Sc������h��t�O4��D�����dJ�����<gd|5���)�Z��][�P�����ਿ��+hʁj���Y���1/w�<+��'�^j#��o8�$͗��1��&M��Փ�n_�p�G��l�;U�֦���vE�tK�n����vTROV���0}'@r�:��u���jê[�gr�Yk��e�STE2��3Z��Eꦗew�-G�����������>nl��U�i�^ū㑭';*۰�K�`�9���t�Zu^�

g��޺K�Q��^X�23#ڢ�,\y�,����KN9+X���z�C�v6Q2*Et��#U5Z�=~M�8�`8e
���]�s�4v��Ot�ur":J�!˒Wd�}%A(r���R�����/��I!yr��1u�søz!ި�
48V�tR�4W��v�k�%���_A,���7�j���UՂ�{[]�y����Q�ۭ,r#�J18�>�����Ex���ׇ�\�<�kM�U����*76n�Er8U�X�'u�P*L� � 4�mL�!���UcK��X��."�8�t���$H��"�۵rv ��JU6A���	��F����p���ލw�ZmLc����!W��Z��9�Y\tv��%�)�Z�.��gV
��)�0�b�D	�dW�7�=γ�[M���B�q���s�ǻ�'�V��JK�=�^�^LՔq�h���)�� ��X8�M�'u�" �7�yT�~��5�ǎn�N��pȈyTGy�
,( ���!/���bY��`�#4��Ǘ)j.5Bf��S>�C�p)vX�]�+��sy8��,YD�@�Xty�
Uw�Wl�k�i�	��	�A�-�JܝأS�ǫ�n`#G��۬(�KANUL����Pt3]�2��F�onm�o���"d����K�PgL\j����b��V-��߲�X�`�=r��$*Ƶ�ӷI�w���`��(!5D�}�9 3�cd-��H�/#:�hs-椺[���T�(��z�.��zB��L�٥p���Y�6�}U��ޗ�OS�z�ZM�R7�¢��2��2��G<��i��M�V<^����=n� �).�u>ܠL0vj�
�vc=ćg@S_�֟.��[�~���USU-oWw��0T���s�Q����X8���*�
��2���OI�p���}�l���HI!E�TYďD��d�E��BW��@�֜Q�e��R
؉���	�-��!%E!;N����J���I�pK����
��H�Dg@�5|e��/�rM�<2�|�2�Z�7�Hf�x���X��_(�ā��p�0��
��.�W�����H,�!D�!n����ɺ!�������؛���B�ڳ �h��sM���T7�J8t@AQq�������	 4X�c�  
j�D �e�u�U�W�%i����RꝖ���~���a��T+� �2H*,cH�%1����i�TA{�$@A�H��DB7�ș*�,!	N|�t*9��Gb
��a�	-���[��O7�,Ӧ�"�n~p�R�Ҋ�]e|C�ڄ�˴�t
���H*/S2c!���v���q�dT����X���	���Ϩ��x��n'�9 ��^k̷N^a��� AQu'`#��\�B����$�X �3DQf�9� ���S��_T8�Iv�
\�%��.bU$#��e�� EE�c\�"c@fD�C������KS 6��@�%ˌ��PI��YB�af���Іd$��x+Ld���* ���&{�}4 nM�*->��O� ������f�f[3�\ڟv�ڳ����I1��C=g$7��<�$��5���s1Ow��
���SV��~�� AQx/�@� �	���~E�dz�G5�iyfZ�*�L���"�0@Lgeǜ�]xe{wxϻgOa��8�5�ΜZ� ��̈́�pM{6$O9p�HL`�(4�5��h� 4J�+-�
��x%@.aHAQ~l�? &wk@6ǉ��w"�*/�qD%��X8p��+R,\H�9=R�G2�{����)}E��.�p�!' 