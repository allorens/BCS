BZh91AY&SY�ߩ�߀@q���"� ����bF��    ���E�()I5�[��QimP��m%PkV�hf���+a�X�SE B�)��A�mb��*S[Z��S@2�lҾç@[`����S-�*ڵB�E-i4�--m	f����U&�يSU�i���ʴ�T��Zڢ�U�Y����B*�l�a�̐T- �/}�'�E���)�ij�٥[T�iT��ٴ�J�j�*[�cf�SlԤ6k!�J�ij���b֭�I6maQK`Զ�Vѡ�r7m�֑�Ԭx   cs�4��5\�&��c���Vv�n�U�4�`��J�����WV꺚��U]t�Uu�]��fJ��hjl+H�b�S���%��F�E�UL� �������(l��]�E�w@R�ڝ��k�uJPPή@*��` 4с� 4�@��]Ҕ�]>�{lҫh���[^ڜ`V��  t�m��v�p -��n�(9ˀwl� [��5l�.J��((�7�����@�2�t  ;���z�Z 㪻@�-�H+M�4���  ��ҁB�����  zy���@(/<�x�m����� =���և�n��+T���t ��e��h�]���C�r�6�%Rm��6�kR��x  �� Р���΂� 7*�*�������N�u�R� �ӅuN�AwmsL�U[J� ��q�4
 �`���F�5�ʂ�@
Umij�x�  {σ��Fn9��@U���*��Y�  ��u �4��\�]\� �C���)AuqÒ�.���4v�"�l��Um�6���U��  ^( QK 8à�5�΀ v���P�p4 �9u��� �tPP	�b� �ӀQ@ƪ�v��аƃ�6o   ۼt �. �8@MT ܮ�A40Pnv]@��` �  ]v��h���搵m��ٳ*��   E-T(�`4 s9��v��v8�@
m&
 ����͸ֶ�]� (��a*�5����֦Fx� z� [8� K�� �m� r��@qp���p Q�:�P����h ;n44h}�   �B��*R�i� `���1JRU�a0�h�����)�)*��h4ɠ 4  5S� IRU�a0�h�����!$�Bi�S�G��i��0���!%(�ꐧ�O�6TͩQ��dd���)�u��rū�y�k�3ұ����L��+E������w�_����~�����UU��DVEUAS�P@��3�UUE�|_�|G����T����+�z����� ���J��""��������?�s&���aO��l���C�O��>���)� ������dOY�G2�Ȟ�'�	�"z���'���"}�'��#�"z���'�	�z�>���)�"z�� L	�"z���'���"z�����!���
z�����'�)�"z���������� z��z����� z����z���������������/���!�?L� ���)2�0(?L(��*����2�>��>��>�(>� >��z�+2����>�>�>��>��>��>�*���L
�� �ʠ�
�"� �"��(�� ��
����e�W�G�D�W�TW�EW�W�AG��C�T�W���AW������'� /�"���/������*������ʉ����z������� z��'���z��2����(z�����#�
z�>�'�l�f��=dOYC�A��=eOXC���
z���	�
zȞ�'�	� |1�"z�O��?؝??_>������Fl��8�(���p�!��*�b)a��n��e��M���=��Q�M��ީxD�"j���r�uǢJY�6��:s�#� )�e�aq(^�A��
���]Y�jv����� �r�U͚@&g3'l�#�'h�p6T�˫��ܢ�r��'*N��ȩ�T�(}�ˇR����o`��rw-1wi�<��wrCs
)*��t7�v֦V�ʋ2M����[�6-�QknQ��֠�ͅ�KI��X�3su��W� �;�ܪʫy�l��-�Z�TX�X��­Q0�����j���5���)�n(ʌfM��]^E����ە�n20�{;n��ݽ�U�M>w�������{{
�[��X�R�6�r�fS��`WU�pMY�>R+���"��4ķ8���t�ٹ��;���6���Տ�n�R1�*d<����\
Ӹt`�Y�U�����!:6�pT���n��N��r�U,��Gj�ʾ�B��*>�;K\&B��+޳���EP�9��w�H�8ku��Ň�<��pt�ޢ;����~�>�xwՎm�7+��YyM�g�>O��!���
RqfX�H�n�T	JV��4V:eh�a�6Γ(�����<�9uN���+�&ɂ��9�GN�b[�0[�ڱc*�F���S(;"���'\d��n���[a�#8��e�5[�&H�]ܛ�s4�{=���E�RPR��ɔ���%��b��ѧ�����K(mCjM�s��Ȇ��K�����NsX�^�4��T�gt�����I%-8���9ic����Xx2�h�Pݟ#��^��J�={���G�^�T�h�ņ�W��mْ�ǚ/a$��&�V�j-�;h���'k_pJ�}�J�܌̋^��^����ll�A�n��]:4�����v�f�����^"�r4R�ON[�|%�Z{�����
#����}3o#�A���]:�IC���[��^O�;t!�/�f��S=ծZx�,��C;	��;w�^Ui�8%<�=nv�i���n��&�WL����ŧKyU�' D�����]Y;�L��ѫZ�V�����z�n�L�O�!���tu?v�Ʈj�u+_<��)xTZ�	�k.��L딷 9���R�붅�Y�l|첝7�Y��d��dT�vh�t�rP;���E�nB�k�s���6F�+I��0��:�h�ʆ{��n�`o�N��� ��(�p9?Y�5fgfN|^�U��WS��Olດ"��ݽ�`������a�1�A��ݳx�N�Sl�,cIx.���LP��3X)��Ftp���Ͳ�Z`Y��p�V��h걢�N�o�ꤓ3�F�p���^wr[4-�zY2�w+�n��r�&�y�����{p�ݒ�/`lbB�De`��ԨY[O(MQ�������0d=�Of��WFoq�
��KNsب��qG�}Vѐ�J��'e/t�O$"�wb=�
	O`��x��c�N��������<}�g>��Ɵ���.��(ݐ��^�oU�Q.��qv�ԭEg��[���D�;��J̖8�o�F�ֲvۮ�[�[mC/�[�Qն�0'���bۛ�R��F+G\w�n�x⭘��ɯi��hV~$)t55�ַ���h�����{C�#��륜Z�*�VE���n�\��NU��6qN���.�ܼ{z,+@���d�tt������1+w��*e�5����[�k&E�ja�IyQ�X�y&#�L��ْ�b�]���`����	�sZ(�8_:�Gd���މ�4���ל'�"�l���ُO.
����hW.L\�K����j��y���!W^ކ&a�m�r�V��}j;�sW4�nM���N�5����\Cw�F�B�W�^�o�����k/a�iu�擌�R3�K) }�w|�Tn��-��R��k4�_gm��uP�cI#�װŻ�aD�7��m�=��G��'w8R{�ӷr��M.t�gV�M�kHl�"�4uފ�Q�݅�"����hl�1�{����d2ݍ��zZv�-�8�_}|����gF�K�°�X�`ܥ��ͬ�>��Gu��^�D/_��)$v�xRFPP�IK�=s��u�zHv5N��I���I�Ӏ�p�'��ۉ���ׂ�9��V%�(h�[2�gf�\l�Y�!
���Vf�@��{O[�st�{W/Π_m��O����I�E;�D�>�M
߭�	K�[X��4�L)+�
ZQ�3D���\�:��(���$���Kr΋�Y�]B7#ͫd���d��v�s�vȈP��i�������7*�j�@0��D����@�KzE��V�H����k,�@uUc0��xKyW�!X�\�,j�	�QdO��
��ȞM=;�����c@;�B�+J��[WY��N�Y�f��(��i��,�jkb�v����vu8�r�&h�r>� �9bn��䮆��Vǧ��F����E���,{��5-�lkYl�wQ�S6��5a�.�О�v�2m��Z9iSm�f���5[Db�:��,	r�%Ƿ����\9�l�r��#��T��@9�޺� �n��Jw���t�`��Ą�ڗ���e��U�aTE��-*2.�^2���9s0�:`�x��+^�i
�̪�q�6����ؘ$'e�Ŏ���]�����UF(Id�������f��',N�nN��ђe9Q�'/`$��#^݌Uj�iJUSk}k��/�N��>[�1���U#�����y �؅���*I��[����xzµi��/���p�Ȕ@�o97������)n�����<x�����h�h����/wZf��e��oIݦE�B��v��+L{�nw1۸\DV�PVR�wCݗ��d���Z�[5z;�Zh���Vk�V�:����Vv�.��L��Z3u6�gkn��m��:1I;M�Ԯ<�>��/�DΧ�M�^A5����C�ݸr׹��d�3�++;�ʩ]�C�xL͏�N��˧a�VP�㉫�X������FyAu[̰��e�lZ��R}���&�*L��f�攺�9�"�/�9W�i��Aٵ�,u,}2yN�\8v�s���Ǧ�$lTΓWjt��3O,�Ʃ���֗	�_lT��q:��j=��	��JC�1i����/��%ܰq�r�hn��j�rJooPwg��#3:�b�x�Z���u ��^�
��M���k�[]�n��v�O�ZL2[�s8mÚ��mb5	��-�{/cMw$��rU�,��8��:��V<�=�Ǳ-�<�6Y7{&��lf��s1�9y ʣP�2d;���5M����NP�jJ�ՙj�bk��[j��u�X�2��am��w�n��/bԁ�pGmd�F�Ƥ�[�,�d�3���&�GƉ����s���w�^�N��Ϸ^"J���*Q�,Қ�U��	.a[L��(&e�r]��X��jw(�2�u�l�γf�_|��Z�����&a�b@M��L	fs-�Zk���ݼ$n�~�u�Elw$�VN�Tݛa�d��(a ��j�UI+̵�Z��H��uQDa���0q�J��a�HՈֵ���WA{7���Q8-.�M(��Iv]K)�DcWNB��f¹U��yf�����H���W�I՘+�]Af��٠iZu��>�L��(�A�Ow��c�/Ee�!��4*�h�X`��9��-&(�8�6.�VA ݷ�����:u�ݫ��,·��WZ3fjX/;�U!&a܌d��2�,7{B��)a{���O �6k�f���ah�$8�=��vbJ�S<�/t�K�����ᒱݛ���<��6-*�y�$yiQ�&/t��e�pVV���ݕ��L��iK8���n�9.y������ۭH��E7�`nf������vq��g	w��0���v�^H�{�G�i�C,��,�F�Eb��w�ߣJ�C�M�ܒ�aGP�2�.�2��HA��&��PiY6��)~ٙ�Yִ�kHʔ�f B��Z#�	���� �])Mm	��К�GjCbi�C%<�X���E]#�U���]e�f��5�Mot2��vƲ2�C�J���T���cMG�.�ڋ��_b���n�Z�K���ma�]kD�T�mw�KQj��/�_g�m�7����gcC�=4({�R�V,	έ%�Q�������F"Km]V�����//nQFC׽H���u�:��`y˯-�G&�5�+M:hnl�8>ēٺlI�h�Ҫÿ=N��3���t�:��k1ە�!ײͣCF�m�*
Y�h������[E�XBƪ7U �F��r�j��h��7�ŋ&��}�H� ©iR����Tga1��7�SZ&k+[�	Lކ�d�w��y��[���wHQh�C�X&����4hBQ퍽�4Tؘ8�e�Kj�m`�rV�8�ݦd�*U�MS+C��Y�-����0�b�u������F��;�P#of�^����{�tÛ�r:�˛E8��Hf��c��O�8����=�{F�Nѽ�'e7zԅ����P鎔���æ��Y�f�I��h ����v�r�fy������Ъ���E0Vw�zf�u��G� ]�g�:r�\�nM��z����i;��w���׻�EI��A�>ع�d��\òhbb�ܙN������iS������&��ƛ>wd�;��B5�������Zj��1Zd:�6��f�x�HУX*�zX7���͕����-ÚZ�]vl۶����(4wsގ�Ph~Pet���޽�{�;	�b���N��o4��$X^��f�赘�ۄ�$޶N�I5�FR��-=d�@�ܻBwU���B��ڬڵC���U��>�/*{d�sf�7����+9:{w���/ui<������y2YUv����p�:�%�'dY�Y�RI�y#�:)�_>�-.ˈ��T�G�a�r܋.1�+~'�f�K�;ZV�Eޒs%������_*G6�hshK�-0��\:���[�C����^	��_tZ����T�Z�u����j�a���n��k�E>V�}˻V�W7�#]x	�MY����a�0+�N)]��Ӥ�J�&Jk��;ssxw'�R�{�d��G��z��˧�Lwzm;�AxSC/�DU������!�k�1=�2"�;l%q5��{���LY���	�z-k���\i��n�.^-��UǏv�4z�hYg�t��ir��kz��/5�Ǌ���r;�بDFT$�Q�-r�\���^.d���T�ݯ����Y��ж���'�U/+s����8�5���l��fڳ&#��.�l��
����e3�t`'����Z�}\�f!� ���wQ��D;aL�'i9�r̜�f�3i��'V�� ;g�z!z��Θ�ob]|���
�=����O>��)hL\�[";��;k0��A���P]��">�^�&�tX.��h+u�NIF�v�^��)i"ͻBg4��%��"�r]�R��NIA�g3L����f�F��7*�c��)�vB�1joY�2l4)��|qe-&�;-yQ�y��NR�ea���J�j`�镹��m�9�m=V�@�����JP�
��*�kj��C%�h��sn�E��Di;B���4��|x��X��n�����+a��A�La�Q=y�1�#����lWW?�u�ݿlߓ���gq�H�%�M�Qo²�=%B����MV���Eb۪�)�G�e�7ge��^c{u훓Th�Y��;�L֝TI�_K���s�Fiz@�/4����yN�^��`"��[Ky'�{�e:C���:5hƼ���$R~��:�Kq�Q�o.a.�N���N�хn^�\����t��z��#q��/,��]����Z`���Ʒy*ң��¥� kW�dc!q����߹ZaӃa�[e
b�	CQQ����nĢ���7�wB����qb��8�dcWq��!D*�n�O0�̎�:������.���p�v.��S
��6��we�r��mmWHGf��5�e(�x%���3�|�P���Z�l�t�V��ɰ�'PB�i�j����΋t���^QYR��ͨ22m�Gqǽ�l���v�s��@�2Y�T{�ڗ�ӡ6iq�h�2޻�-	�;�Y�k�[�oR����V�hgY��oMn��-�2�`4�!�7sT���a�Q���,�;�P.�i|-�^��
����Q9J���ҵ:�WH��S�͋n���RL��X���6�������j���h�\�ۇz�)X�L�i�NM�Z�ZB��i�1�
@�5�8��1+�������Fdp�M$
ܡ5���vV[�c3��nk׏��s���	�W�V	n��M[L�^=��&����t���ɲEY�w��:)�r߸^��$8+�������Pp^�lf�*�e��û˳(���R�"6�Q�b�hMRBX .���G�}è}5]4����.���.�h�U��͐U�q
܈�X �������;���Q�������JIN&�rFYF����9�f�7��3���*H���<�pG=��u��+\�E&'ԍ��r.W9��ˡ��z��j�sM�g(y�a�� :�ˍzmOo��{=.˞�u����Y�=&�X&��S�L[���Fn���\<ȫ�M�Mlq�Q�.2�x�[�Z��zO�x�1L�:�(o�W�8_uD�vU�S}���m���"�u:�����p9w��|HGQ�+�ĂW��إ�p��������[������/M�g���������q�+�Z��$b��A/.�gfl1�zݹ��w4��/:�2`E�^�J�P۩}(�2	v��y�0R�][e�4����'N�%6��Z��d6����`ůn�!��NKg)2��]�,Rכ1��ͮ�n/����=R+��FS���&ܖ�� ]��w:�\;��W�֖�h�/�m��h�`�%r�u�9�a��դ��!c���HuM�H������&��*���ф�i:VO^�9�%�X����� :�5}5���n��Z��v��Ž/�
�M�X�-�yc
���fu���a��ؘ��M�H�ݼ��]N�Q23f�)Ю�+{���>_F�����g��}�ST^�W�c^߂��S*��R�9�mμ��/����3���{��r�F���n�u�z���Tu��r���������|0w���vm�U�9�}�nݗݕ+c��{e�o�tx^	%��\��v�����>�t��x��0�L��oGV�m�}���~P]#`�#�z�nrfQ:�׌Z�wӔ	k�/��ؓ�.o����f˛=eX�J�E7����w[D��k.�+��_P���S(�OH2t���A���3�V��/�U���f���K�Wtz ��sy��醫�z�|�y�se���sG�̘wN�R��w���l��$���>���C��U�LwC���x�r{1�Io�u ��:k.�=����/�í�G�w����� '�3���.;\���Y�ޘ.pŻ�76`����L�"8J̾!���2����z|����Y�3j�XyRF��N��7�tZ���j��p�5w`ܺޥħ�?;�'v�ߥ�x�j*d)���'A�5MJ�[՝6�ѝ�(�Q���+�M��揷�׻���,;g!�
g�����t�&!�nl�5�\mC�2��ړw5M8��f����yý�Ⱥ�[�%{%���.���e�,"y��_�$M!�^�_���ʹX���.�()��Rv��j����.�}��MA8����E��ε���ri��g_P5ѻrzE�h�)�kU�����PL\e\"�MW��[}O!��@�y�ke(�U{uz��Z���OuÖ��qܞ��S`��9i>�V_>�6)�P�]� ��s�}a��9{��fsc���([rN���a7�[��Ӊb�ܱM�26]_�N544*�9g)�|����0݂MrW�7;)%���3Ge���䵂��� #&Y�ڭņ,=�d�٣�v�(sW>|y��)^DG���>>sm�O:2<I1ts:�u>��� փ(RY[�	�df����DX����6�ڊ�&�y|-�é<�j���G3����k�9{��4\1�@ޚ��fy��C�o)J�צ^����<㜻�i�9��hG�F���m��w�BL�=ϙ��Ո���λ���2yБ������k���S�����z��4�[��b�<��=�y�U>�GΛ)�}y9�a������9�0�sC�}N�k�o$�ÝKn����"��q��iq�6�#��Մ7D��Qǌd���o]Z��@�F>�:��Zs.��{��\��x�����ވKOPw��0�!��ͼ
���=Xm���`�mVs=X��c�s7���]�>��033�8��0����冖d�Tu}G��J!ڭT+huA�d(S&���bvjE��Gv�*ֹ����阉Y�Ѩ�`�36�]q9�pP����Z&p��y뎓����L��W��h��n�c����	��$ۚ��)j���j�3pm�p�N�k�N�)ՙz0�ÏH7Kj������fh�|�[m^7�v� ��Q��3�l���v�r%|�{��˛�ko#����kd���L���J�ԙ�����<' �r������:��tDk�mW�V'&�H�*��a��L���W�����h���p�/o��J|&=x�t�5���jK/��0���'����sR>���f�@�ܓؕ���cp���܎��=�*'�w3�ΔE���:3�-�	e5�^An(5� S 炯[
��X`a�r*:1��/m'�7pi�4���{޹w/�d�}�k.O�-�nkz����F�Q���Z0��Z鸳����ʷ���q��e�|֪��ێ��f��K�l,��y���C�e-f�=v�y����p3l�v�A��ƨ�_U�Ւ���{�زq���s������J�Ftb��Ǥt���������Z�N�X��7��Ztհ��+�����yY��o�tz���%J8���:ߖ{�Clp����
����1/z���q���3wV�`���5|�"��:|����]�b)S�w}���X�6j5.�M�9��	U���-�	F�o7�kz,�ӛ.�f),��fWȀ}��2��o��[��NO���0 g�6.�ǘ�v'����t&�)
�r�w<��c��iV&�Q���3f��2�&�T�&E�c�97�Z�**;n�jK�'a����=�����{}���g2�){����V�OY�r�8�n����)<��^��{'d#����cOn�U����'�A�b�fp	d�\@>���H7��z�U)5K����5R��}-$��B�o���;�0<Āk6��({p9}�9�+�8��of��O�HU�k�ä���l�Wv')oh�ޘ�-��\}��Y�^q~�@�.X�J��:�IkIC[���-��}���h�CG�,�]ħZa����Jó�����]�T�����9��r]�7����hNU)+��	����Nϊ���omu	��໵{N�Ƹ+/,�i��q5+u�mMo���.$��ᳩ�KC0
�g�ŕ��=K�w��K�r�i�dݠ�[<���f���twEPs�J��E�xDW[q:M�nQ�ש�Q��i4(+��\1�ܘ�RY.��� ;�c�+^��=SBi>��� �n��e��
f���8�6]���7zV$��_i�ϴ���7L�b�����cȺ_A��8�j��|idV����_[6�$�u5԰WI�4�ƭη�`��<�]�f%�A���'z�So�����n���xy1�`;+���pn�i�3c��Vgj馸�-�Gic�ݙ-sTw�a��i��J����*�/�: ]�اǓ$����O�a���6�l��M�7}���l��k�3�H�_����]�m�H��^����+K�P��l�\n�����	�a�yL3Ry���Q7�
���[��wd�͸��Fز:�a����<�6kc9�I���ʪ�U�Z�t'�Hr��˻��3/5q�-]��nh(
��ۋ�������d�{���}��Mfc�N�ǉ�YS%��y�8S�u�7�n��#��=H����m!��y&�����՞岚��Z�3�p箛P�{��7Z��=��һg���e�z^Ҽ�ۓٴ��%�{U�y��6{K%/\��;�)	{t꟟;D����[�gt&���\1Kʦw2�0Xf
�nB�<��c���d�ܞԕ�\�;p�`���+{��Z+:��إ�n�}[���'��=��Ի���RΔ���a.b���������#�o}wNQW;�v�{��I�5��K�j��E�M��& �f	l���_.�V�-���V��DHl��B_oPҥ��1]R�d�W�9����:�XCk�������9����M���}�!|�y�#����{>ې����s���8bǂITkB�j��#(�J������9s�R�$�n �e���]�a<�bU�o؜��K֎"�p���q��=�^�y�kٷ��":�ǧ2��Y�8	7Ƨ��D���u�P�Uē�{��P�L�
�^�ьҳa(c'p�e�T�1���L�vE���NS��,��g��%��3l�2�t�+�U�U����N��J���^�\���d.vS\��C{�rNIp����hA�v��y��N�#�,��0iGN����j��GY5�wf:��yP'�ς�F�;W��<���:k�����ۧ��{ӾĶR\J�2�p�W��/*|P�akd�u��H��u�^��6Lk=h�Tw{�L]}~0���O{J:�X�s��]o$�&̡Lg8���S��/�wJ���W�Op�i:�nUO��,m���ӑ�2k�X|��YD��/{@4�zy�K(��]"��̓n�g��yw�q'Z4�*�n���m�fu��|v,�v�ϢfY?�w��n����L��u{�ų�ǥ��Xcb� &Ϥ	��5.�h��Iv��3�v��]	Ǘw|�>MӚk���A��ș��S�IN��̭�!�X�E<g.�R��'tG�{GQ��^z�>Ӣ�Z_z� �����_6q^��,�ƨP�Fp�3{�k���B���g�-<Ȝ7��V)�I��HE��fv�.��a}�gj�3��<���gE=���mi&,W���[�۷[�|i�ܐ�G6�j�����H���m��oޒx�4@Z{���y��-�yJ�)��.fF�;�o�gf�d��oF�gsF-��PX_]��9%%�n[� p;�����5�d˗���X���S���Nو�'n˳�!�إ�K�w��	��;����fa�(z��PE]���j��f-��}&X�u�x���m�ڴ�a��$X�Ke�8��^���9{��<\��rt3J]���<��"f*��^Qk��g,�7 )���;�P�'4>~�?4�$����<�X�;md�k�ƋGe-���Yўse�6�-r�{P}����^n�����ק{�k�k��{������G�լ�1�״F���n=�L4[���"�(k�6m�O����vM4kUJuw�.����p��1J��y�+9K4\@=<����a�V�7$���f6hi��+/~Ӟp�>�����+qҔ)�)�#��`/r�	*���6��]5�s-����	�wg)G�)Ԓ�V�W�ɬ���e�AuM�P�-{���n�*0�ޏv}BuՈ�a˛�[O<���O�ajr�������c�Qgy>�]1KW���ϝC<Y��8x��T9|�B�ٳ8�_D,��W��!��
��=�6�C��''fo?at��)�왱6w.oT�lF��4r�Dթ�nf�|�(4jH�Gp�n�4u���X�a�zܔZ5���ӆd���Q�t�R���3S���a�A���8�i��}��6����%�>�-g<���������P�/[:έ\eF���Sg
]-�{^�M�BfT�l��W���V�mf�����y�s���J6"W�P2	HÏ^��"�&G;u� �u��1-���3_T�Yˊ<nk���˾�2�vo�ٴUR�ǻ��w��7�����	�a왌"��&+�OJb��i�uԢ���ʭ���|t��)`{5f�N���a��L[�D`���qwk]hhǜ�㹋�n^�&n'u�]�Z~赕���ڛs�4�0:
m�>�l�)��΢��{6��y�#��˰��[/o+;����L��Y��h=��܀#�x�n�6��c'0�$��mj@��W�����n�M�z�@����\E�B9�Nj�j�*��rm�ځٳ&����5��z7�A��o�m|��1ꇟю�����P�ɞː	c����pȵ0�K�e:z0PP������iU�m\2]��M�z�m${�iw����g{Ȣ�v�YY��� t0��wGX�14(	�)�{.N�?I��*�{��ڶ�͐R���\�a�5tG�wh�*n���Ω�4cƛ�}��tL�k������%Y-�5ͤ���X��b���r�����iLxr�>�[2�=�rúDP���֩DE��[��MYa�U��*k�͗W����:��wc�Yu��X;r�r7��6��3\�h�H9�G�e�Oj�����t�Д�)��s��k��&.G�u.iք�؜���ݜ�V6[�0����!�S^��Qd�N�-2��,Q�ه����tF ��]���<*���!&f�+����ǃ�_G�+��ڃ�%�?n#}��=����w��Q3ZN�w5����l��B�˹vꂭ˭����|�$6���}�����s�m<��t��(bF-�wϗ��װ�#�))�V\�����O��)�/�
�v�_�_�&�.�\�例y�t��M��.���^������a��ʿ6�;vp7�t#�YI3�$g��5�\���ϖ��г�{k�	'b�5�^��o���O���w2�w;*�yQ��qw%d3�8-�ŸJ�+�y���]!�:�f��̮\,tu���\���
b'Y���^@��q�>F��Ԧ�����5����Q50Ǵ�o�ic+id�_-x"�y�K�R�ٰ�e��̾�ݢWB�{2o7���:��S�	�:�f����'[��Wl{�����R�4����_=�v�������<3��f�7�޳���\A��]�������x�SI����ك*'�V�&3xc�8VTǸ��<��}�q�5/.jI��܂a��<C���/����[svŌi�a���U�0KНiv�L#pap$�\��}�Xx7����՞�?o�*�>X�(�az��;��f;mK�^$襈di��Rމ�^V��3cL��ݻgn�JV�7�Gf]�7���=OK��S8]�d�:�9��K��M�So��`aKzەقb)��r=ɹ/$����E�-lV2�]a�,q�Jo>��&P�G� �R�M��8��Q<��z��!�IA?��E�H���F��2�KWh��g�0���@4����с�Ւ�G��h4�a_�j�#_�c�5��b� >�/��R�t�[a�l�4�)|A |�?%�(��j��>2d�s���]�"������o���{�~߷��S���HBHK�����=���t���|^��nb���Kޮ�E+������r�z�r���	�M}��ܽ}I�5e�ŝ\ E.���fW:J��;'y�>)*�ɵZ�+z{oӍ�у�j��[�gf�"�U���nj�Z\kM��o���׳`�ElyE/!*�n���ӳ�]BU�=)���9��f�8ZZT��'�R4r֞u�]�eu[�`7�CbC=a؎Z��l6(F�V	s^o+����1�s��(�]q�0�3i���F$2>�}0((1`~�������qT�p�I�˒�s�ZމXġ(R[�R?*ܣs��D�\Ǚ�G����WG�<��w{(9)==�ȅ�O�r?u�v{_�?g�28����LI�Qn�2���2V�\�^%Bc�[��w�crn%�y3O�Xgq�'�:�u�H�}R=C �ȳ7ζ^�q������ǷR���TKoh�y�o�Б���"�t�{F��N���X�`4(�ڇ�#�f]��K�N���Yn[��!Eǜ�������׏#B���t�$��WN�d�J�u�vn�e�Uz�{��۔T��d�B~|���8�u��Q�\��0�s/�)�K]�C2��G���/v��[�.�Vp�ʝ�ci
��Dz�89K;ƤG��f�����r���t�%GF�;��%��/�.�a�[���%3;������YkZ����b���@ C.�գ��r[�׷�jFN��u���dz��4jx�6�V��2��zb駜��g���ӗF[�$ۺ#�DykFV�؜�%�3 �G�g9 �Zo�JG���3���K�����j�=�C�x>|o�Ǐxb\:���c���[հ��m(�fY}�A�0��7�!r(�[č��4D{>�Q�k���ڏb]�ք2(��`��6(eY�X7f�u�kW����z��}N<�;J)
�ƷK�2��qWp�7#[ww)��f���I��T�{+�QP{�Ӈ�X3������佷�.�"�l�ۉ�]��CK�Yz�W!X�lx N�oT9]��a�U�3Hl��v+���$y�z��]n�H�cR��k�<]\��
i2(m��gw~�3D0b�rA�(P�QD@�Υ]��K�6�����n$����������~��D������Gߍ�եui�h4V�pή��M����[e+¸��;#�_"����~���>��Fx
�s�`C��v�3��o@/�$]}-Z�Ǧ+�esT�_oD� �A���-4�_���'ƞ��kd??`u��{�4֥�}���K���}���oӤV�;�T)b!6:zN�á.c/�xK퍫��RN�u���i�8�[��k�#����
d��&���sKF�� Q�Zwǫ�Y��}��=�z�4*��pv�a�3���x��EN�m��}Z,�l|P?_hàf՞j{.\�T����v��2o@�ݚF8	k:Һ��>���v���*e��4��+�MJ�o���Z�Ԗ�N��4ỏhc�
��+s��CQtp�tĈm�8F*z��7k�����+��W����3�ϵ�c��oS �	���/�d m����sī��z�=���^h���(�f�ҫ<��G�L=yH$��Wk�߶
��ڃ)��j��b�\��v��,�R<�k�fz�{�8�ٻ�ɣM����C��8��b;�uV/�x[�.'~���ON������H����@}��l�+e��7{�[����u�e�%]��5;N��T�gR荚V�]�{�\�"8�4>��ҥr�'|��A����g�p3.pn�}a	'� �{62]�ȭ�+���t)��^\���3.ȼT���@�gV<�;����4v��fr�S�yՁP�r�L��A:$�[�bEfb�R���V�0�������gK���k�6�e�V�]6d$֕�ܘTs2E�=xW��<w~)T��&�Loz[��%:v���)ǒ�.)�lZVѩ�bGhJ�dn�v,���>��:��m)����c��]v7�Ճ��xX�����!����7�������{&{�YW��6���v��ɪ+}W����bp��T��Ov���{;���`&�B����Z0�V�̀�KJ�X��W[�C��
�Չ<L�po���ݸFv�n���YBݱ�੘��ճ�q�U��T��;rA
H��H��1V��ZPf�^��q��l;w۶�9�jW�=�1y��q.-���(�~��}r�x�{x�^�n�lJS�y3��=��&_gW��s�91�9��d��OOl�u�/F0Š���s�a�;���h�#�k�=>���^Q�#�q���-N��}�n������ui0g/z����;0L���8V�1sa:�����&�t�ܚ��mH�����ō���o�Tp=Ʒ�-�������sL=�$�o;n��]-�Ms!���޽垴�wIX�@"�,mtIz���*��C�0VC�;�\��~�\[���Un�4�v�f��*��>��җ�o��_.�tL�&����k(JaM�ѓ��wk1>8r;�}�%�6�!�^w�נ5<X{�c܄r�<�t����v�ϦE8��o�NmX|8��oz�I,��V^ne�K���A�ZR:��7����ȷ�OZ�T�ӛ���ڽ�4��n�x���n�x������(-<o��:v#x]�jP�%�,6���*N|2�:(G���^w���ц{&vz��c�m���ͺ�(���1������Rp�@`}6W�V�f�xŎ͉;�+��tu�Z�랎a�Xo
x��P��hʹ��x�X�����=J TVn k�^g�ٯۏ���5U|���8�yӬ�_�a��~=��^�W����o�H�V�ï֨�p��P��yO�����7�D��̾ �}��2������{���nh~6�f(�LG���M��X�]֪e�V�U�Ի���B��+�n�H<�ݩ%����F����K�;s��L�˂N³�Qݮ�gs�y�cQ�$�6��%��1��&me@[t7GlN��1F�R�boX��ƽ�`����h��n�a�@��V�"�9Ӳ��=�V9H��ZV�n��e˸���=���GN���5�V
[xK��СcO0C{��܇�Uk5��UN����eiF�֜�dd�H�k-m�
���b�v]�5���vo�c���8����P��+P�C�.�^�ȋ���� �%fc���.���4��tD�A�Ę&ͩ,#�p��j��}Ͻ�g�%N��N_�h�%zTAH.�=�g�v$V+�xl˦U���O����[�)�.����]̹����uk�̸so`���W!7���#H��Zs�<9E�la����*�u���/gz�%�J�����a�9���Iԩz���pn\��/�� SG�X�s��T�VǠY�M<{�*�o_n���1|K�EQT���ے n�S���iu�C�0֮$������uэl8B��A`����4�z��K��OG{'�V��,�u�ݽ��
��ՈZ�[څ%Ҧ�4�|���c���&��j���{�N���X�����q�l`-Ĵ�N��͖ʼ6󓘙���/�)��t�䊾������r�(Q��s�;0K���=(���b��S�ID���55��(�oqC�:�걢$o���w2��,�����I�u��-�񖺤&�������˾�/�d<��X�qy\o��
�$^�����n];�T���/z<5��h��z!76��*2M�<Xŉ<��<����;�M�X	��u��A"v3JKʝw.�7�G���%ea֏��sg�\]�nm�\!q��3=�)'fnD�ĉ�Y�1�5�J��e��s����O%���)�1�S�ehwy�p���ȱY=�ɡow�^K���d����}��2ݣ�����Z���Pݧ�zU��yS:�ï0�����j�;*�zĽ��P�>ݤid�pһɏ^��Z\,��{'e�j��6��K]��Y�!��<�Kw�3ǻ!5�i�Ԩ�ֲZ\�;~�$��]��.af�hJ�'0#�{K��z�q��z^4W`VLݻ�a�^ޙ1�ZQ�S�{�G�����.;J�{F�ᾇ:�K9���Y�X�滍�<4E�ѵ��E�Ǳz���;�V ���f�z��xVX��VU8��s�����G�q������X�9�/m��=�:0�2�-m��j���oڗP�)@��o������j��p�\ϳ����H�|R~�ǽ��o�ٛ�W����q�Oo��A�ԅg{�}�6O00��}���� ��z�����o�WJ ��h�t�n����"A��H<�20��y�0�ŻX�/��L[��R��Qg=E���'t��|	�Z����������V�]��}��!`lg8
o��|�)����a�Ɋ�s��Jg��w���-�V�qr��n�������V�(� B���,YS�Z.�R��o%I{y��+2Û7z?�j�g,WȌ�PBZ�d³H\Q'�KV�ŵ|��.л��YT3B��n�{�D,le�B��#]֜,��i�����,1*���su�L]ܻ�7���}Up��d�ea�Z��'�r��#����f�_sd�d&3*f���챆҅�C��Wl.�Cr��f�HŐ�Y�*X�Y$�љ:�u: �xbWc)2:v�3�Z��^�xW_D.hؒ�<�{mA�g���H:ռ�����U�%�ƤYFt��KA+�k��J;����M#WwɘյS�y=�
a���֛��V���n�lM��W�r�J��P��W%^�d����fHFrb
틀6uY�f�ۆ[oU���R�o��e�
��K��]�Şƴ@��U��s��7�O��'㪛;Mc�F�o2Ա2P(���O����ZSZ�Q�g�F��輽�J�-����s2��hw\���W_oF��{�����:�Y ����[WH�չ)I�����j���ǭxE�&s�0OH�=�yN�%[�J���{oz5��ۄD����e2���\0ܭ�P��3�Bv6Uސev
�+�R��A�26cð��em1���+��9��aC�Lq�5<Ar�<�ۛ��G�M�u���eH
�v�d�eX�I��ۑ�� ��]�9ԙTq�ۉ+�QU�u�T��R�ND{8b͛�RC��˦�+�����gf�j� 0���n�ˆ��f���/�����-�j=C4�qC}5]Wt�<�źu��W�olL��Xa���"I笝��g:r�N^��u��֊D���ϋ��K���1��.�J@�+��]����`)���-ݝ3E	��-����[9�?V�ǇX<�������z�C�F�Ukt�ֱ,z�i��T�+�;��E����r4dw99�
͔u���(E���i�L��&���K.�n�f��t�;�����gN��9E]�o���2Ff\N����F`�}k"�,����h��T�yY�ܕ�>�Oi�hC��@w/|})��ǽ�h�cxA��v�{�z�4�м/��3�"�v�dFY׵;�t�t"��3��ή0�V�|��wp��h����o��I�]T˫�*U��m'�_2�����L^��,[�1o.�xAk�Xh���Ϛg�ok=|��FeV�Ra_�����]�bW�vմ�U메�d��]9"��܀�����nhi��f��J�RAU�b��N+��7Ɠ�!w�=┹����<�v��A��s|�X{��}�>�(��Y�%��>Ȝ��{a�_�fgx�#�e_?���t�s����|d��?z
&�˙���u�-��KblN�N��<�j�팱�8sq_C�M��C�s�AwU�͑yP���o@�CX�]uӭ5B�u�r�e݃�i�@��,�)t�.�TJ��[WRC��#�g^��Ǘu�mb�ζSi�ѐ{w�ؕzt�-��s�V�[W���R*}�q&�^f�o�T�M�X���}�Ľ��}w���l4S�y�i���u<�Փz(d��X1��DYT��is�m��pY`K����}]�y��̼�c&+�O�3��E*�f],;�!ن[�tH���Ҳ�eȁܰ��m����W���%��5��V`R0ESZ���S�K���Cܐ敚x���yV�\�lZv1����=�J2�,9����O5�Uc����9)Br��9}�Ys���>w���7�rX�:��ι^�&M܊!O���j�g'�JX�-N��o�zne�WZ�O�����V�]c�]Gz7�%p]�,Yy�B��~v�1?�:��W���}V����x�֍̤��1X��·��4:eg[�f�����T��AC��DX�S1�{E��oe�͗�5_2���Y��2�����;���	�{IɊF���p�<��y���wswj5�z]X����gNM!�3�O�ಜ�h����fk �bi����{V�S)5ݳ���$�̧�0t�Q��f���k�r���}���^מ_(�������('Z�S����VB�x�j���N+�E|1}��Yy�u�*-\��7nB��MC��)�M��@fV��F���k,QbV�Gl��zT���o�}W����9��wҴ��;3e��X[��<�J�]�O�<m�r�<"��D���[�71�η��`m_^Z�].gDk��Js'h��F�������۷!��X�[u�d¯8�h8 K�k���7���q�dD]��s[4���9*��f����Csǝ�҉o�h%��{V�.��Z��%�>�G.Y�oD�[��W��������Z���q�<��u�� �}lp )�k"�F��Cth�7CcI��.��5������hI$���M���oW//��K�.+�t[-�E����������h��l���ɩ}�6er�Q�$�J�*�Љi�d���L��	
k�F�W�����Wՠ��O!׌��:�:��r8:�O���ku5�"�5/����^*9x���n�vA�c�7�Eu���wv��g�l�H��OXgw;�@�3�sx��Q�x�F6�^3{�X%����/d�=A<��l��{`)r�i{C}���c�ްk('ex�m��˞���#[���ս뫊)e`�Q�ø�1�d���^�c.B�L�U�t!��|���3&�^�{U%W�ۧ�q���L���(TףhRuH�3c{+8�},GՐ�^����w��\�dV�����$g��/�{Ϋ���7o���[ן�<�C�<��b�oo[�\��1�]�]����o�V6%p��\��V��5��o)C0��-2�����V	��x�:�]4��˺��y+����+ݕ�.�O)E!Ƚ/u:��wCH�{�`KZ�u�d��see��w
3v�*&]�b��w����d�����zob�*z�Q����N�7�M[�e��mi
����VLl��Hy�7������Vx�\���]Հs��w��Qd^��C�����cn�r�.:�9^�t1�*w,�n=9��L�O6���"~��z�|�?t����Ӟ��,� ]��^n���N�yv;	:�c�!�ͩ���-��b�+�
U��J|���>"�I�"+�)�(2~!�[M�&%�#L?�SM@�-~i����d�$�aB@H��HZW���+�kF�(��+m����1�m�4Tm���E�v΂��T�(�h�`1��Z��SEkTP�Y����ca�Tl�ض���4�������6MS�F,䢝b�`,m-.�h
(#YѣAm[`�(�+X�)���m�*�*"�b1l��]b����6���A�j�(�F��c&�8�Q@lh����"*,Z
(�b�a�mSPEMl��Z�%k�m���M=��EU�F�b��+Cg%`�:z)��%�Tm�֊m�EUh�Zm�vƱP�k5��th����MF�0j�(��]���N���H�Z��Ebͦ�-kkj1�Uj\Sm���l6���j�*Ѵj3�55V��m�h�F���A�Z��؊���b5��h"&45�u�*�
j��A��1F�
�LF�-�Z�l�m1Z1�Q����(�#�}����BRS�mٚd�.>���ԋG�5ɹ^��nV��`�N�$�$�,�n�ȓӦ�ڹ��,�٦���:�յ����iiI��vո��z�U�a��S��"�}*l��\��3�4M[bW���yX,��vz24����k��ru�6t�'��5�h��-�!ݳ	}���x���_��6�C���J��a�W�1������㾽�S�O�f�'��q�3c$2*��$Vz��V�[��I�s�M��+���˽��gFۓ�}U==��ڲA�������;/�Ŧ�����%5Bq�t�#��+r/|����c�,v��*������u������
���0+{h���>�z����}�4�����?{�o�����X#�n/<��}�n)eg�2'�в?d3k��i�A������T�n��
�xμ�s��8���s��Ha����O�ӝ^��4�����=�wHǘgiɋ��܌�7�&߮<H�rC�1�˟5c���M��Di��l�6��.�N�2�Ej5�r[����q˱z��:t8��-&���d.��5)��Ξr�����͙��{,����Ev��Ei��3u!�d�b����т�oV'����,�\����N�ʞs0W�q����b�t�w7ˊn��R���\ʕuN��^�<����`7�,��ݓEM<'���^���$8띣�ȫcڸ�X��*�x-�Ꜽ&�9f�a{1Ѭj���2M��n#;2'Ē'��=�}���_d\3תg���<H��X3٫�M�:G�.1�F�s� ��"v�ddH=��*���!��)zQ�v�Z��k��T��c�ȹ����A�n�I�i���1�4C�i�;����}��T�c�Q�|fɬ���4�x2n����0���i|�{V#fFO�:D��=^쮬�z����g�����c�u׹��g{�f�^����꥗sh���Sly�׽Z8^.�Iz��ڷ����1'(�����4�~2�<j�o����k?3LH��{��{��[F���`�0��Z�|�x޼��v36��e�߉���zë��P;�o}V�˷�\���_f�����孈 �M��

u-K��,ŁjWYG��7���Y"�;�S��֙��q̎�2�~�$��6�թx�����'>�!�w5��0<w7:vc�snU�2Qy�r�є�_MO�'#���V��]��ꝑ�{S�7Ŧ��ϸ��`�t����|;�i��I	8}�3m}��ReS�#y��W?2~��6����S;˿^ �����E*U�v�=L��B�=ep^�����z�rl�iOy����^{���Aߝ�v��<�;~��1p�1��8j�y�C=�=;�^�zs���I�<Qvd����_�]�e���q�z�L{�{V���bW��q��w7Օ��&��\ֶq���$�;G�c����-�*wy��${;�j��M~�@�S�r�N�Nx�:�N\ʑ����5�du��+�:���ro�>�8r���ïu�<��3�x���t���V�/�3�O�݌�ܘ��/oi����'lu<�E����	�w[br2A�D������n��q���M8c���W�|�߲�C��c�a]�'~��v��율;C���S.S�=�1�8���1�C��j_,n�vv�%8���>}h�����x����}���l�۠�-��kR��\��Cƾ-.��\��j���mvf֡{�wo���p¯�? |��X<A�Y����^��*�
���ՆZS����r����\��r�))��vM�߻C��k�����?E1z��6����/G�os��H.A�0O2h�L��^�i��ʕ�u�a�=���%�fz;pa�<$W+{�k�hs��'h�4�z����w���SdTҽ�~�=�I �67�A�Q"��gI&�����^���ҝ5Mw���oz�x �q�����#xt��3�\Z+�ɑ�~�ON0�._���CӨ���M�}���Mv��=�.�=���N�}�35�y����|=���lAM�=^��'��l�^2=�o[پ�����~85���Q4�g��O��|���UM��n���I���|x�-����[/��rc���^roh1Ӝ{���O������}�י��^����qǲ}�H�9�b���q�Oz�=��y�&8�h������k�Q±f��1�-{2f��-BsDuѡy:w�gb�H�;���M����ղ�L7���Cy�L�Z]B-2�VL��ҵ�~1;��H�{2�9G�b�~z���}R���yri��"���ڲ�-��Ұ��yBr�7��D�D�s̽hiUcf=�ElA�m��U��U��ƭ��7b����v �ni�/oьI������ޙF��˱���H�X���w���c����/~�,�^���X�T�N��2��hG=�x.Qz�MjN�۬����?�C盂��?d�6��19c��~���я�ݯFڝ�h{�z��Y��E\�a��=[��`�3Q�i�ݞmzo;�B�{�;|�^�Owl3��{�4M������D�_�u�'I9։Ӣ6�� ��옯n����I��uY�}üZ��j�W��(^��O�2��l�:��w���p����	�s��$�鳹uB��V������ >՜�8*�z�����J�������RTv�.�,���<����������=��ߍR��c��{t=���?z����c5�y��������j����}��ۏ'��D^֏k��AT��נK�%rrʧ�z����.Vei�����r�bƣx��Tn(׍��_Q�g��.w��x&s��ߑ�Ǥ#x���I��_J(��ڽ���ƹ�7'4�pW���%?T��G�ݣܲ����m�'��k:��ǱM��ºI���q` K�����rM���m�}�;�\M���'x�w�g�8�����zq��$�}����Gn{�^�+$U���G�Ӟ�~>na����m�h{���$IQ?d5�DS�_O�?b���8|G��O��������AdM�!<���/������ �׀��r+6�?��z�ǖ�k�,�GZ�kW�f��=�F���c�8����'��m�����ʼ[�!���/_�����ړ2��4m�YCÀ@`�a?WVK��^���U����Ϋ�6���嘑��#�{M��Y��O�?g����������z����N�e]�n��6�d�"Ox�����g:^P�Ŧ�?_߯o�s���w�%��hD�H���w��� ϻ��:��Z��ν���o>,��/��8�O@���Fl�1�i ���W�R�sk����:7���uCv����>�}�y��7�%�͇���,Ʈ��v���gVZ�V���{��D�6��fO6��"��o~�{���,����/r�!㲰�Fw��p_MkGq�VH
,�n�9�:K\a�3֧ua9���k-�ں���"��rE���nO��ȩ�궲���A0����7z��=�e���S����]���&��6UX�c M3��c�ȇ$�j��~�#ewL����^��׆O{��E�����|G���F��p<���n�����޹��F�f�����6��|�g���]���3o�u�>�>:�{؜T�8_��u��e�I�|Z��铜A~���&�Z^�ۺݓ��nG��vM!�E[a&�#cϐwbcr��U��*y��U�LE1s�I�yۂ�i��������{7˟`]�B4j���<��y�d�j���z)�&����g��nW-�\��LUJs(R���mQʂ�-�y������4����^^)��v͚Q��l��+�w���7O�T�V����^Wv��\�Ǧ��Ⱦ'��I���rmy�zmYb��k�������=�h���0_(��=sۧbw����/��^�pl�J�"�a��6耩�∺�����{J�Ǖ�t�:M�y6���*�ͻ\�촥
����*ȱN�Z�c�����+g�_�
M��W.�a��ۙĆ����6�Ei�H��Z��ŭ�$2���,���~�'o+�<s%'.H���c��a��G�&�����Y�MC9Em<_k'�ٯ�����>&�=���]]�N���>�G�3~�5�x�DN��D��^FI�Dt�<q��D�qr��|�e?R\�~�+�_q�`=M��0��ɡd�f�ʼ�Ʃ�,l�VtÝ���Foӄ7�x�t�sj>��"m�x����^.��6䖺�7��]��"�F���I��I��(���oǭ��=�i�V=Kb�דlV7
"pM`�[݃\�^��L��Ʃe������f���{ݙ�Z�u��t��>p2+G��3���x�y��ͷ��]W��7��|yk��#=@q������xu���������2I��Kc#�=�["?,Y���TL-�-s�%ϻk���7Տ}C���o�w��~s(nH`��V��m����o*r��a���N"i�sN��"��p\��)ܽ����r�ls�e	�x��p��\�vFCl,-x��]�P��6r��ad����qZOAf�h�=P�I���w]ua׻]�%7]��'�s��}2y�z!>��]
��U�yt�86f[�8�%�V���u�7���D�A�x�\��;�'#���8n���RObݺ��@������N*�>3��7�E�^roh:r��UA��3��x��}���߯⭴��߻��|��j���`PЊ����q�t���=��S����3��^H7��EN��^ ��� �gl��E�&�km��{z84���ܝ�=V�n� ����կ�3s>Yc�3t��Џzu'|��-��-���X0�):��]�:�Ĉ=���Xc;�8�A���d�B^�&ݣ�J/ӓ�=S�|���R���d�5\��g��E����[O��g?k����m��9s*㹻�mvxz~�����0f�&��a�/I�3w�4����<�P�Տ(Y{�n=�ҋ��L�fK��o\K�䘃�.F�TM{Pe#KWq::x˜¬Kڳ+Ӵ�p�O��"�а��@����Z|+����Z�] {�9�ԛ����M:Cҟ�����y�d��c/ay"����H�kF��u�v�<G)��7����vx�B��V)]4[v��h��l}*�J��z����E��1����g��C�q��6�t~����;$�c�5�_�-����rE����ug�\���RX��?RW'y�����x<u���!��Z��e�.�}�����S;��:rNލ�/�_��=���A~Ӱ�Ќ@�����:[�R��o?.~rM���w���׺g�ߏ����k�w^ˡQZ|��W��̳��v$k˚󒧾��(z��[��oI�Ӟ�O��|[� �w{�>��L���ط�S^��4��dj���b���8|G��T����ܙ����m�l�ݛ�=�A�e��ͣ{�q���~�֑O}sѓF���)�*y!~�$����#Rm\�[�j���+�.ύy�Y��-�wsm�����C�c��y��wG`�������}�ޟ}��z�~�/o����{=����k��v��S����_������J��$b��t�x��j�*nyk����cѱ���"[R]��D8@����#蛽1梶j�d�Ývc��sS~n�:eT�0�V��B}><��ܞ��"G�<���e�vf�y�v�0a<�yܔ %��[ݪ�:90�Ӯ�n>jϣb��8�i$�%c��^S��]�]�|/{+"zj`nXU���P'��{�,��&��l4g+�=����_r�R�P6�\#�:��_YѼ��v{���6�*,^�p}f�=<�Ĥ�7W�|ʔ�1M8�sf�mt�fV�SU؜�:� ��/���8v�W�ǹ=��u�	G�H����~&�s���6��p�dZ�.��l���un���^�Zۤ7���Ki��ݸ�yI���ދq����Z��U��9}%^��k�|�P"�m0z����C,�S���۝)f9b�ls�L�O�8>:��K7�4��Ǵ+^�^��x<*�u��8^�o�<��;�]b�r��b�8�8�i^I�j=ð*�����͉�hn������R5ԡ�.�N *�*<�(��� �����v��M�^��q��eU	ԏX��M�;�D���4m���L�(h�=1�����u�z�fSU7Uxϼ,3#��A�}���j���x&��V�Q�;����e跩.�I�.�Gi��'������^knH���w&��@�߽=rK��L�ϱ?Oh7��*��i�ػ(�1���8��<U]7�W�&���7$�(�Nj��܃x�G=�.���;�L�+U9��\�):{�|�x��T�J��0��r�Vj1P;��zw1�{��k�	���Gr12��Kёl����,�{sx�{�k�B#l
�b��zTϴz�n7�3{�7"�	�'6�y�B���z�"�Rg�#���H轺����b��uv�舺�5r1ڮ�ur��>���0[}�mV�x�9/'T1���2�f�U1�6N���<�;�^�}�U�I@�q,�B�2���	��ɺ� ��nC��m�g�%��,K[��<�������=�yI�΅�)��j]��	���t�qdi�%Yy gGW=J��;�l�ka{��kJ�#�o��o�ӞŇ�VQG�k��`�]�
n���{�����4		dsF��!k\�r[���oP�]����p��ju��tE�&X���e��v,�z�z_@�yכ��-��uē��V��vfZ�9��e�s�����)���]ӊ���V�H5��R&�aC7,ׂVr��֞�^$�R�n��8���{��w��f��o�� �=)kA��1ୡ�4�����)����{����́��b�ѭ�8��Z��q+_y�J�k~����Z��%:�{��}"7���nZ�[�Gt�,>�<݀�N�\���2ɬ�(������8+�����}�w��v�g�:m��]�y�|^
i��yD�$ m���Ri1:#m:4i�(���Z��*�M[��cc��z1!�&���.��4��F��Z�Uj,gT��V�v��I��6���؂a-kF�`�����[1&�#TkHE[�k�Z��"v.,Dy�:��EZ4�]=.�IU�/�`�����u�cEbӫg� ��(��%�F��J�!]!�ض'Dm�m�;�ƃT�8�h�t�ٻU۶o#vծ��i��j�S��S��cZ{��:�LF��7m���P��T��R�I�URA��l�m�V��v-��S۫ͣ�(�F5�A|c���.�n��1��ty�f���͒�͂���yw=ۣ���[@I��-6I'#`��$��%��<�"<�v�[xF�+�Ts��U^ֲ��UH�5�r8�uRG#���;H�Tn:t⪨11ԑ�)��#cS�b�����{�8�7Oc��5�Q�n�9�h:�;�#[8��mwqGm����h��Mtu�TX�˸�t�c*7c�H��+-/s+T���j�ӛW��R;]a>�/)L�"oK���h͙���2+Mb��TM�/�͝or�f�t&@�o�Wbl��'�r$��z1988�s9���P����M	�G�|C���EC��goN��)f����KI����@C�|�'���編sNnf��KJ�!�0��"�� U��c��1ݨ�ս��h
��)��>0��?�F͵�,�8˒�moq�A�ȶ����F\ی�/�^mmGgO �#8�i�gO�;����,:/1q��AUcx%~ڊ��%6��~�~���~�<�)�j�>ڹ�=������瘨Z�OʭbO���20Y^�	��C{���q�IJ�<�h�W�w�YlGp��"��*Q����s�W�
V�y��?"p��ϭ�8~�6y���5��X�H"mJ/])�|1�ߵO�1�$i5��7'��|��U��'�e���m�mZ͍��ѥ����1��nC�fy�`�J�|1���<�5�U�9��.��������s��Nw0�^}A�k@��:�hN��:m�=�*]�Y��@r�O�<�A.?ngLt�,չX�]١yN��ri�H]!t �� ��|9z���Jp������E��y���1�f�}�^+��u���w��5L��Q{׊���{���z���Z$sU��ĉf67��=��AY��i��f�'%`M�.-�+8�`=�ʷ!��.£��؍�jS����z�ia��o����y^ވ�����mt}Y�҆�M�@�zn�0jp��=��Fu��-�[DCT>:�?ybC�q"�<(���t.�G�ƽ=B�Վ�ⅳ�y���8�2"_����k��O���}��uW�B4�o�9�yaQ�2�Ny@:�@��]���B�ֲ)��Q��r�?8j�mԦ@�����?V��:�X_��r �`9��|w]����eK�ڻӏֺ�)ie��u�v�hg�e'�3L��w�zҊ5xc��ME�;�*i�rz�j�����2΁����i0q����J�����u	�3Eڇv->&:�^�8�Y��"q?TgM�V\h��F�B���8�<7#�}9��m�8��WF����O�n@�j"��"~m��5�u��$f}n5��y��CdS��|a��-�{���u��k�ܦ���G;�����u��,����"��>lS-�W�T�ǘ�03����D|f��2�b�Z�!.�|'Mnn u��jJO�ga��X�E1�$k������T\9�ւ�m�;c#�E�FҌ����1<� ��-Y0y��A���):Z�JS<�YQm�����S}����k��E��RYc��;7N�x����±�N��#��n�PzGwF��+��dR������C#|��_G�	Lw�0Q�|��٨޻Ȧ�"}2T
dd+���a��&;�װ��g�Eۍ��be>1�vc�\��2>?W~<5޻v����?���KX��Y���Ov��D��}� �����$�"{�޲xh��ū��'��NJR)@
x�����1<V��m��ۗPz/��m��IN7�B�>�H8�2�},�4�v�4�2,�	�=5���^���I�����B��EP7�����O,V��(!�!�Nk��o�0%�eS�e1��y!�����ܻ:�e���9M�.��0}�����ʀK��AY>�?5���^��M�-�3K���UK#	���C�M&V�s�Z�E��*va����}�b��Xw�����2{�F��޽��O�{7��n�Rb��n�,߃�8��qTXP���fT��!��<k��q�{P��ʭ��qQUyv����kA��Ƙ
9�zzG6��4-2�n;�.��S���*	qCˬO0@��Q����Um���U!��fs8�>':Ի-Β��0�@�.�����o�̓��|i��&�.su�q��D���3�2%� �`<�x�6ߣ!�'DoK�Hr�xnN�l�zi�ӽKwOR�vZe������Dg�;>�b��P'��B�,j|��ۜd_�����ʔ�Շ�u�>p��R�٣0%�ǁʝa�Mې�g%e�d��;e<�z郌�P3E�jfe'�de���nK�����8{z��
�A3�z�Enлx̉Z�öi��n��ի�	�R"m#[�nՋ�^}��^%��X�����8�~����B�|=�}��6�2��v˰�|����?�(�A��i��ʺn%�����2�Y�o���t�i�nQ;70D�i��a{+���Z{k`�;�8�㐁r�5曌�MC�.s�;y��}�؇����Z���t"���FNe_>	�֣w�t��;���gaU�B��G���oN7��S�l��Q�/�ׇ�gf��P�΃�Ƽ����l[%�j���tG�d�|�&U劅'�f��\�ѳY{
���r���ƛ���{gh@Ű�!�0��=|����ɽ���kV@��q5�^�;�SJ2���8�����k�x�j�O�B�$�C�Q��|�x'�| ��i�C�{#�����ûM�y�{F7/!�3����;�M�Li#I�>��kT��k`�a�$D&��nz���9�y�s�����cdG�r�I�l�'L9/T�t��Ʊ_0�n/2���6�0�(;`�@�F�7����jd#����7B���*��]^����T4I��0�=P{w�#����,鮉A�����sO��1�%ց&m�W����qTa�Z��3j�H*����B'��Н�Ŏ��R�m��1��!c���zr�4J���5��ڥ\��IռV){�D)�wx��{���w7���;Ut�	kNZ�gr������ �b�jt$�Yph��갳:��*�w,��C�� |�� �]�j{x��(�E����_jW��>�s���@uM�w�^6U�U�+�J�8��6�5Y��[�9�ދ"�W?�N�;?���� �Ø_��!�\�S����3��sx�Wз"^��G{6I���Vؼ�6�֔zq�w��^ۄ�������'��PhyD����>��1��Tɪ6���f�����Ԣ�a�zHzZa/>â-�WX�}ɟ���x����H�����S��&��m��OJ���~Xdf�6y�=�>���M��� �o�w�~o���&��;��e��ޥ,�!��8(�v�)�z/�oP��ރ,ӣ�K�����މ�x�\By��Y��ᛯ���R�3�aif����X�/d�?NU{3�K��n�vPd�|�'����٭�չ��9k
b{$=�Yu�z���%��8��Ƚ������j��	g������9/x�(7}��^����ܥ-K�{�Ӭ=ہ�ޭ�|wA8���d@H8Ș�!�\���=ܽ����.��/r�d^�SL�M]����l����|BϞ~Y����;�!_�����AW72�7���;$D��6+�?ίl���/����:
�1WV��f��8�;�(���6��E�)2��ʸ�V�����R 6q�U����l��y��Q⾣��gQ
�������$`��f��&�,N�yW��������)�J��ֻ6�/	��"G	�K�'I��7�E1��&��ܞj�=9.�͋Cƻ�2���[ڼG;5��T�m;$1�a�`�̧q#M*I˼�)sυ{>�G*1c�q���e�Y���:�/�޻K��a��#��Bcc�)�^�C�a7C�(����[n�:z�V.��[�(����B��)�rsK�a�>|`|��D9�6%�=�u\כ��yʹ��n3�����k���sxv��ܱH���&�z&;�������ь�C\u���<ò~1�'�7����)���Ǳ7��l��f�!LP��mv��S�b0i�T{�Br��H��� �<��.�imn��J�)7ٺ��)Ԙt�C�UVJa���:�_���y�-��������i���5��0�5g��4*gC�c[H�-��N�Ϲ�Dwa���K�4��䢋P	�c�g7n�Ƽ@Ƃ�"����n�C�^��x��>�!9l���lN��J��x?<�Ρ48�n0�X�ZU
��U�rw_��C�����D�y3��4�)�>2�я�kN�vװoH�^Y�io_�COO*���f�w��u���1�m��Oq���z��xs-�Y�h��I^�a�	����8f���E�9=��Y�V�1�9pQ>�}�/MEse%$�TZ����`�u�O--��h����3F�[˵+O+s����#��r���+�_8g�.�����=���[=�h����h�}�g����fXo�@r�����)&0y�>#Uߍ�+�x�~��G��̅���ޱ�V�w9c-�<BZ��!�gY�ٳl� [:y��`t��=��M���2��������;��V5{zO����YX�ӌ�c��*.�ǃ0�X��=�ә������p��Bbu�tk�d���tc��9E'V�W�+
�����8�����8QS��ٷ�F���w��AB�l�t��^�7	��ŨtBd���rQ�E���`��[	�`Vjc��%�qW8�8�@YЫ��|k�H8��!�_K1|a�4Ҥɽ���[5���Gt�!z�5�W=<hӅ��-���B1�C���zA�	d�g����4�Q܋μ��.�oT漥ˌ(/�V����ٮz�� ���j��܀���n�IF��2�bw/��6�r����b�«�es�P�����RX�;P�F��vi��><�|mo=f�H63�FF.W���M.���y��$�6��|U��W1�S�T��֧�5F�M]��c�݈U��v�|j���jF�w��b���9����e^|ϗ���{9O@��Q���| ���
�m<�j�nCڌ�gdU1ҝ�K�aν�́y���U���P��ܰ�IRo��3E��<`Ů��n�#����=��C|=�}�W��}�WT��4����sH�>R�\�n�2)2�n52�Z�
�^�Ĩ%�7`h�獢�&z��X8��=�}�L$8��d5�������^ΒÛ
R	e�X�p����0�V�/wg��������5,��@��^�9�~�MO�<�v���X�?�?|��h���f������㳻��0^���C����H���g�������%���<�O�ᐹ>���B����k3��^�N�=yCΘ�� ҏLG�N�U�6��\3_�ޡ�e�pt�m>74?Vec��[��������ٱ��l$X�_�Y!L����M]1p鼣��9�-{��}����k	�|.&.���cW^UKcP<�.{:��(2�	Q�47��Mk2����Ke�r��;���]_S�b��<��5���M#��9�lc%�j���t)���Bd�D��;�.c.�e�����&�zQm��V�b�=[�M=�Ϟ|��i	ğ�`$&��CH�S�fQ�f�u>��+u������Qx��T&	���B�ɼz��xO^������%���ޔ�0�{�|g������,ɵ�l�4�r�:Z�`�F���G/Z���K_k�
R8	��ޫ<rZYI����X�K���E��X;y�p���jm��v�,��H��$Ӯ���6�)�z�x�4��XFi�6�P���|��f�j�_�x{��^����OIvނ�W��)�x�K"�=�ƂF�׮q�w0����H�]���ކO�$X�a<g6);���OB�h�w6b���t��M���ӱ�NY�6��]�6�U�hB��L���[�a;$3s(`7d�ư�
8e;���aը���T4I����7����m�����P�����:�/2mlX!<����|�3lP�r����׭Gs�1�6]��!!�h�V�dmޝ����N�04�'�`8�Ds>a��k�	٦�%��z�o��q��&��f[�K<�YY�v�N�Ծ�������N��փ|�Ga2#��6�k��m�'n�];Q�f��T��d����>�z�3�GnY�z�p�fp8Dw�8(yϪgq���ջ�f�-Г��l�m��_�1�IŜu�&+�� �-^b�<;��ݞ����q8c�9>�+�V�����k��h9���
^�(H9L��C�N=�T96u�9ogvd����q,����2O��z�x�w�kp��L�C�KJ� ����Ы�޺zjf�ث��&/��ſ~c�����v��n�;]�՝�;D������q�@��)�z�Vi�K�)�r��8�T
��|yq��h��"���@zi5mjI�.����ѝ�>��d�>���d׵Ǜ��a�F�uH٫��ށBO�������{6w���k��SAv����3��LX|c �3�ܹ�5>�z��Ư.J��=��u�!��SM��T�]�FCr͜`Z��v��ٟ,2��:
I�B��J�����X�'��F��}���j���ܮ^^�"u��R�&��i<.�a��1���o�ZĘ�|�L�/�5rl�k>��2����kz���# �𜮾k�D⊉d^�SL�MN�omÞ���=��y���iy^a�D�s���ۣ������Z ���A�K��N��1�ީƂF�Xq�<�Us1������s�C��o��e0�x�0�m>��m	��ʽ�Y��Y��'M*I��Rr���5�L�m]�*�sm+�7��CF�A�<�!�[1�tN���mE�v�0����O��Y�h������ձ��;/���E�qyAt��H~�0�`d	x<G�x�\���zW���������ݖ�jډ�Û�أ�)H��zc���,Htq#�
"��@B�Q���<L1�yy�m'�[�J��5
�(J�L�BUmv4�O�x��y��S,ٯN�ۃa��}ą?O���~_������~����~���>�}(X���[�
��W{��f�7��V�Ds].��Y��a�.�Ƕ�WяU��v�2���W#����C^��z�;,��w&)Q��hULӣ����ܡ���ԽZ2�����ښYӥ��˅��n

�sBTu}}��]�ۚ�b���Y����gb�5�Gp��Me噻���gl�%�
��㽾��k�����h��}� {b��զJ^��ب�I���3�i�ۺ�t{�=c�8BP[v/y\�=�3���iX<�����	��df�:b�]2i#4nx���R���'�4tb0{�Cü��U���{`:�9�%���-��w�6UISn�Cl9Բ��N�`�]9�+4D�Аe�f�ݽ�!8��l�ͼ����ù�R����(E�Ѳ";�t�s�77g-�7�s�s��~l�z�\�ڵ�m�,+�<`�����#ԑ�:v�v�o^ܹ8�W#՛�i�A��7�vZ�a3+k�p�*��$�[ڲV�y:%۳P���Le�ܩ5����?���j���*�"f�)�T>���i��7��D��~:U��;$����cE���	2=[��#-�2�Y؆&(�CX��E�~�/\�Nlfι�0� �Mwd�z��1�y{��\(���t
B�]qvR0ua�n\GFf:
�ڨ¬�B:@��1L��C���Z���%�|ZT�s �)e���VN���ޥ[�)8l� �y��΁Ik�ݨn!{�c��nmeсl5�:�x�2nt[s�w�d��K�Y��Z$YV�$Ĥ�w�_gS�Zq��7ƻW�j
hPF�P�kzQU.'!+�ă6bN�58b�[V�f���ot@��nX��O�z�z����<X�����0����y�M裑l��~��f�=��j�[ԺpW�ז�������חs��.���l��[�o�@M�z���zl�P�\�X�	��.���:��^���������0+Ȼ����j���B
ħ4t���Į�[+,ތ+*M)>V�]:�]�@�v�;cf޴�Z�ž�r�K��3h�I�BNk�Lg�"��7I�o�B�o9�g,m�2�[�� Rɵ̈́F|�y�ƍ��J�-��2vk���N(���6�찰�Q�;zA���W0�ޣ�ټU��$}W�,\�ڳ�ԊA��FN���z�ξ�ޕ���\�y�������ch�;�76�F.	U��{t��Z���9˭1J�lEy�=�1n�P��y�ʹ�]^B5s��\�D��������u����E�'=�L�*\f�li1n���ug'�~'�z~��-�M�ok�������i*�	���>�3#mܺ����`N)Ԭ[l`G���u���y˨�ԋ�&!���E!QJ�!a�J��i�dQ�����t����v�f<w�|�I�W�G*F�fL��e�`0=�I8���s���|���Ea�"�E��E�C��N5M�(�'����.�F�<d��ݴkIј"�١�أE��Ӡ�W:	���tb��:v݌Kvzz.�u��Wm�I3Etk�ö-V�Z
�3��n�7b�N�ŵL��Wy�ձ��S堨�n�Rh�lh5��LMUQ1EL=����AI��A��ni�a���:"6�10Z��SDT�|F��tQ��h�k���v�N`�()�kF���QN�ҶpMI5)l��5��
��Z��+4�ĺu�g��LJUQO�k��v�UWM���4A�5�=����h���;�kMj���i;���Zi���`�IWN��F�3���b��7͒�#��SCڃTP�S�v�F��̈́�6Ɗӵ�kM|vn���V�D�]��w��t>c��;a��T�ڝ@f5���6���O�ւ(���EWG�O�ؘs7nv���{���Y"ӣ�3陵5�]8��3/z���9���I|�n�UWl}�yX�5f�X$�ĒI8 �{������ݙxp�y�3�
a�=��=zv�׆r�j�u)�W�ƲǱ˧շ&+��_l?��C�&ˆ~m�ڪsݵ|��6CC�<	�O��az�����hGP�I86�
�M'�ړ�j���*c��F�$�5֤S�$��gg�#��=�Ag�X�=;#Y+��/Z�i�O� ���,ѭ�\B6"�c:3����9�z���F:HDYz�x;п8���	>���m���>V�"/����׌W����wbf�#.v�T� ��&a�ᯖR����c���XV���]���}��2�>t��>��N�Ka ��Ÿ�CP(ΰY�l� Y_)ʒbǘ�p�Qg~�1J���Ͼ���^������P&��V5�!?5�� ���Ƃ]Z�F;�2��̍���Z�jq�S��Փ��3p.)!�2�']���&��\�:!Z�9E'W��ŬTXSK��E�N���W-s�]=�/EQ�>�AX�~�������'̯��&^`p��L[����?x�J�A�Ms�=H3=�ګwoOv�v�QN.�l�	�hUӍ��gd����P��bE�j�y�?�{=ߚǈ�8����Z�dh7#=Aa������T%���s�[����`�z�%
X�8�kМHd��YN��%�Ce�[c�kP�z܊��sq+� f���Iö�c���ALt�m�W)	5�8�����8ٷ�/?�xx{�sU`�=gkb;�c����<�^�9@ߣ�Ӿ[�	F@�B1�C���zA�j�{�˵O�NOm��{
�i�R��(�Y�	z^4�o<���\�����[W�p��M7"�t��f��P� �m.����U"M�L$ٕ�V�Qy�T�(���O�����J�w��]���Ŋ�������@P�<��:�7B��̜qv8�,*�O1��Z�S�֓l��vT�ǭjԷ��NZ���`���y�sX ��h�U�u+p]��^���<O\^�J��kk3;�Qp����'��d�`�y�~j���Pl
�v]^�I�5{T'-�
�W��L��[$�������>�ۗ�(�h�W��A`p�	�R�]bdG�guM�~������F��ӱ@��0��K��]�91���<�����q����=�r�:�=�ji��)�`ާa�h<��A ��4��tg��s���`� ~90y\��&�2�VGp�&��Q�+�%�=�M�fץc؝�ɃE5��@��B��4�q���G��M���2R���#������`��p1�Iy�S����!���gNl�a����e+�o U��~�Vϣ��^T{J��٨�0z���=�|���r͞��	7mr7j�8��i<�o	��(��i,�k!x\�t�b���{�+��5��)w�O5�|y׌_b�[�,����=�{�#ݱ�V��7/0��,�!�zâ�D[��/>��j�U-�K���u�dVe
7a��ʗc��ז�]y�sW��a"�*��=�	���i��Ҷq�����:��<�E�,3����cK�F�����m�-�`�ƍtk�(��QE�vg�/�pX�����
��������Y��m�-f�m�S<��LPRU�FM�־��{lw��[�:A�Zy㔩�{��2�e���׺�"үO��Ru��YY��b����k�B��*��۶���Ĭέ�Q��4bf�}`J�ЃD�T,�w�,�'L,r�E�3�����c��$�SvP,��K��o(5�6�p��f�t7p�n�2����]i�?7x�,g��뾴���1T��Y{9�vgC�"�\<,�Ȉ����kdp�n��.�m���m�;BΩ0�p��~��
ܞq����t=�3��{p��M���G�8u�ѱ-�}2Z�UqP����e�j�j��sy[�g��(%�^�(�u	��d.�� �ØO���h�����˷�9�:3�E/W#^5��f�9J}�0���{׾�Oc����2����A�7��拊���h��|��b��"���� ���Ǥڳ�Fc�ލ��8��v:�[O8άY-������nr��)?d�򓬻�A-�d�>����6�Đ��>o{� =w9ݶc̽N�_�[6��	Rcl�����}'XE���=��n��;�p�\��5��Wj8n�)�Be�3{��؝���6C�ϯ���}D=�- �1^:��u�v!�����[s�+N��)w!��k��3e�N�k���9����׊hHG�/�V3mq��@�:����y��-~����8S��/�`���d��{I��1o�����U+"�4��f>�1w����}��"�	O�
^K�P��g�P�,>0�>_��^�S��[���� ���fK92�u�'�N���ٽ��V�A�,�`Y#������f�J��߄G^�\?ߋU|���#"zVSjW��o��Z���ϐ	!)��)A�W�)��1���Ƕ����-��
���mwt��qѾ�
�n���{; ��5���'�%�{)M2�(�kw�{njgNv	̋��2s�z/��r�tP6|bK�e	{���Z\51G'.񮋣)��T�cIMmusIM��&�����u��s��A�.�.��$(fƑ
��;<P�,�Y��4ʔ]IʯG�h*_#.�9���O��q/ʼ�Bc�=�D��{/I�K��46
͚2���s�{L%��g���ܤ;�t�m��M�3Oڽ�g����3�N�g;���p��!ryCE���Lk�V�{�����/��;�ljXF8��N��b��]a�=�)�WB��++�_}_}_|=��p��T�6߸�ލ31W𞼒��Ǣ��|�>��y#��M�;<��k���K�<wX��N��T-';*Qm�C�Z~)���Pu�Q���!��|�Ƽ952���WgD-};P�k�d.b����(�@_�i�^�w.��q"�<(��ܩ�BA&���Z�p���q��3����ؓ"�Ђj��L���16�b�� U2͔6-ݛgg��T�b�}�#[r�c3s��*aa��C�~OBz�hg�ԦA�k,{E�}[rb����7����*n,=;{�qUm�N�.��mg�幗�>���t�@g�0�N���0VSH;�/-�^n��Ί��=����[���a �&V�����W�~�[���??9�&�b��j ��Y���t�(�d4˷1/�� :"�׹���.�0v�o�D�N�ON6ۗ�8w3(M��q��'tm�^�ɖi@�<�[ ������ˋ���`���$z
��zD�c	��I���-׻k���v�MG�tV��Ppq�b�VI^(γ�l�*�i���I{��U������:�ma"p�n�;�H��X����֨���|���*){.��t���џ*�=s�ݞ$�l.���&f񡴟�7X�������|�A엛�����9eڳw���d���N�����<�Q����0#j�^Ɇn��rQ��ٞީ�=���xx{�   ���/�0�r]�:9��8���=0ۚ�^�V5xoA	���	ո��vq����7#�dL�,ݬ[z�jC�g�<�!㝬.�dՓ��D7�u�~��Xe���"��(4��5#�};v�7<��2''c�_7mu~�����Mх��5����ވL���_�6��zx��M(ʍ}�f�QN.�gv=4,8މF4�t���C+�f!��T���֦c�C'6m�/67�y;!�YZ�<�b�sȢ�\hӅ�;�0�h�d��F4�r�k\mڵ;�ѐ��{��k�]b�,m)v�0����X^2�x��m_"x�X@Y�tK�|<-����ŝ�ݠ��@C�c�CӱE��MУxi0�0��W(����`��ٚ�I��3��9��=\���/1m����О��W&�Y��.-��a�E�k����ԫXna��ݮ�T�j'"g77n��ͅg�� ���Bָ�>T�8�g�Υc��˥k������Y)���2�5��2��z4�=B9�Pw$�`��fp��4�|Njv]��I`|]��]/�[�� ���̴0�o�^�rҬd���P��^C���r	���a{q���+��ps�;����]��A7�Q^�=�
�^T�;�玚��j�VhM�)Kjlζ�S=%LH�GJ}G���n�|�:$^����V�V��3��1���t�.y�ovV3��xxxo{���Ui��V�(
}��< ��� 9Wښ2��3�[+��3+�P�s��@�g��>`e:��t(f>��R���o��߽�,������j�e+@�,+�Iv�2�q�2�t=1΁l��^]�.!�^�;�)�}�>�|���\��`Ԉw��
i�Ht���i8"�WD���٩:,�Q؎v���̈�<!c���)��Qx�ٮu� �Ku��n�|�;"����;��F��K�7nY��u^QL��Xd�l]���Ʈ���Ơ�H\�vd`|*����Ȧ��������&�������	ܩ�sc����M�8#��#^ه�j����`�YT5��^�g�{ۼ6!�BcAb�I��Wm�zw^�1��@��v@���C�	���AvZNO=#�z�C/z�X
���ħ6T�	�)*�،����xO���,�CRv����n�V��������{!�
�>ΈE�3�K�9C�)�$i0�ؾqOw0�Lsh~6*���` �kz�y�{L2��DA`����C�$J�4���Rt��ʥY�x�43�г����(���8��*?u�C��F֐+��5�ễt_g��c�z�.>�*�O:I��׃��ܤV֨cP/����v���K������Y̒;��`$8�ǖ��á��3vM� ��4/�'�*f뗆1�6�ّ�Nm�%R�*iq�!�GPV�0��ՈW���U�
�P"� P �+�����:_�eB�4�����io�B�li�&Ꞑ�װ�
7�4��P�^W�����(/�FUS���f�>e��ҭ�r���Iĸs�o����M�"�cBvi8S�MȪ��W��5Y�Mó�n�߹<:��3j�w=,���^�<v�q��A�������-�>Iț���<V���ss51Pz��]��^��ԣ�\�6���GH`�áy�BS�����3���M�p��k|e�=�.�I�O����>�z��jnY�z�p�܋)]]./OVj�=�<)@��y�����k˫6v_C�}g���]�ޏy׎��-��93P�X*��n� �;r���D��B��ĩ�{���K8�s9���-�H?x����ԭ&����D֫��~͕����Q艗��ȖxAiid�!�x�z:�i�i�ALُy<��&U�X{0�ˑ�x�0���_ʇ)i�5B��������^�ҧ����R*`���Ư�s9f�׺S7Z�A�ȶ���6q=z��]"��`qmâ���1Q
b�O�9�����9ʥؑ�jxmh�I�Yy�[˰���u���tc��g$4]p3��&>�g�;���o.�-�y������#�0vh�)3:l켓M���C���0J=!eڽ��2u�6�/��X�8sS�+7�$����� � ��� ))J�7���̩s+8wU� ׫�G�U�	���N��oܥM^X��ܮ�aG�1��U�}�=��Y놆*��=#y�P�8D�[@L�������!��%�{)M2�(�k����0��9(0N�;{�����x�'�$�6W��T/��$_I/^�N��xNH�"��(==�j��3��[��2W53��d����C5��R͵;<W��0SfS��i�I9~��0+��'zk:��wu\.��^�F��0�z,�s���a��!�n���:m�>.4k����g��V�zj����v[э���O�y���u.�a��F0>O�p�s��d���`��u�S��}�[K�j���j�ϙ�R��,oHok�z�Q�����v�ь�!��C+�X��L��s8��R�C���)�\��cB	�k�2��^#&�eG�*�f�طvm�}e�c�eQ�Wk	ά,�D=���v�I�����^�4-[�L:�Ʋǿr��mɊ�4�8�.�73�1B����S���v�
1�
"K<�Ŧ�ƻ��ʄua�pl23D|�/�Vϒ~�%�@�����œf�b+�Vp[��r��;�Y�4��J�3�7�6!�koB�h�ݏ5��)K�����b��9�H���i�[g����R�_kC���=x���5
Hٸ?����v��w� }~���@4�4	@4(Ѕ-P%)KBP- � �=�mu�t�y+q�����&�n�AVL���E������l~����Z��,iG3㯻;��\��ڊ�|`��4'�hw<�)i�Xi_����S�������Of�g������6ڠ�$Օz��9[q{C���̳Ni������ Ș��|kO^�x;]�u�D�.��,�$q���7=��=�Ԟg�(� Ũ�CP(γ׳f�V@��y�Ρ-�����������+�GB1遱5��6���oA	����zd	cA.�g
r!.��n�t_-u<_�~�\r*k��;�_��	���~ׅ1�L.z�D �^�E'IUN��/�;t�Itv�J��=\�w�[�>�f���:�4 ��(R�u/����Y�M��9�K�!�м�X͝׻�Katb%?X)P�
Jq]8�@�hUӍ�>0!�$F�����F�=EǸڟ�0����|̃}���BT�2��|�(�x%Ɓ~�/��o'�2�l��_oE����[݊��)�'���N�,Ԥ�c��"賎n[�#h�\��~g������>�_�������}��o������Q��͝�+>�u�y��Mn�ex��%M�\U5������2��;������VuK�7���W�՞ӊ���9����ṗ ;�o	�����!��f7�y�Ta�j��ϙ��+1Qf�D�ѕCԾ%ΘGrw*�I�uA�H�dh�p�f�'��)`0N!��3n�~�,X�8Zy��$�o.�K�쭩����<��,V.uD���7%â[7.��L Gh��+W��(�<V9XRtz�mkf�>�gq�0j�gZU��f�u��&AEJ˳N�zX�(\���9V�(��Zh���V3��:�}4��铟E�� ��mV3�f�(X���j���(%����غ��d�qq�gؠ��u	��܃��ضw�?������g6� ��)8vֽP�Ľ�*����"��Ӏ��[V��*M �bk)��O(�/'j�#��%o�SU�C0��v�ۿ|u�溸����Ŵ�V��U��xS���5ζa��ʔ�[�����ld+�ena�|Y)��v3eo`��$�K��w�r���Z��{��9�
�ե���ѻ��Ӫ�T�Ó�z��D��34��Rc��F�U�GUdr�d��&�e�;m\T�"#�h�߆�^��T���W3j���g(��i��XV��Ս�{�B�Y�R���������m�X�R�mGd�ovW��mzeY�Է"�.p�B-��1_�����R������Zx|�em�B�%͍a%��#[�y�P�l�pf��O�V4�(L�����yG�Efx����8uJͬ!�X\���y�[�)TY���@iޱY�����]��PQ���>Oޣu��k�V�H�,xk���ph��P����t́���/&\�����\�SW8z��'��8���"Ƌ�/������Ԓ��G8'��77��Ӟ��I��*�J�}u�7x�B�+5e��z�9��Yg?���!�z)g���������L6�$ㆲ��{��S���V��|��ڛN�l����Y~S	�D��cx�LڝYκT�HW�x.��Р�|f��D�.�$vWE���#����g�Қ�<��{��yk�U<�.���_P�[�6�^�^�f��ٻO��V�Gۦ�2m�ዃ�8jY�ia��Xt�Ӊ�4.���b�]�Mc�+9C��բ���� ��Ĕ���т��!����wqDJ���E�9_Kڸ��gZ�]]vƼXXe�����U�b&m��Hy��&��܉<�"P���4Ey��/l����;�����W[�/z�v&�+�P=C�9��
�}J��U��ݸ+x9N�}���$;&�2h;5vw�������6��7v��n˫�ðH��l�!�f�6�h�?r�~/��vs���G��r޸��Cܻ�#$-�z��j���H��9wv�@i�FP�ۜ����+QG,�o6���$���� �P���#AAM8�!-��:Mi�P�tZ4�N��uZT]b�v�QHm�7�Z�y�(�t�>]�Y�טɭ�QE����6�(����Ptn�f~#�͏)�ll�Uc�]mR�Qyg��#m:Jv�;���.��h4ht����h�CI��N�����t����&��+V�:�<�%,TPy���b�$�V�v�:^���LMm�wkN��zx�����t�h�\T��E�$���pF�-N���U٢�C1Z�sl�EQ�U6إ�GmTR�I�4�h4U���icM�F���ֺhn�h�4TMtLh�!���N"��']	TWEV��&�S)�UQ���C�AT]l����:�$�54h�[h�;n�
y��{����z�.Y��1yt`�2*5\D�W��+��sVf��ґ�/��������O��,wG�u.ђ���O����t��+H�)CB� /�����߄J��`�� ��|��K��t(�L*��熡j���RX�;P�ޱ�]k�iۃܷu믕��!9�z�F��M�"n/�δI�o�d㋾*�
���c3�2�3�����ꌞ��ԭ�߼���_�����W�q�!q񁎄ƀ��͹�E&P���
���;0�lGwod�4���*	q@.�<�<�%��!pc?~q��ϗ�lG���H�eS���7�^y?n=Wog��R��ýAXe�X�]��9�j[��z��^�9�"]�gx<!0��=Wd�k�Ǽھ��ww!V=�&]�s����v�aED�j����&e�N��-��8�r����tn���9����-i�������59Y����~��D?׎����T��J=0��[)f�N�n�ˇ�{[�ٽ�j���fp��3�"Ӊ��I�ME��_�as�l$Z��@�x�&�t)��YF�&oov��k�>dc��(z�X���~!��W��)�������s6��骥ͣ���N��R�׏���8w��Z���r������ƃ�~ׇ�_�lv�-q�������yy���5��]Ĉܪ
���h�F-�E�\U��_�����q�s���:7]d߯uEL;1*7���5���j�ָa��06�����w|�n8%K�㎱J����0N�����Q���j�
�ݻI�U7OA�a�\r��揨�P�dF���fQ
��*�h���)dff���EN�Rzҍ�%���	��JBd�H���]�.���z�o4��Ё�i	Đ��;\���J�{��t�C`Q�����j�A�Yx��L)*�ߣ&��k�<'�o���O�Q2���n�c�ٻ��Q~�A���^��}�L�N��K"�<S	L(ؾq>x�}|�-������h0]x�4H0͓�.x�!��%U�N�f):>pUD�K��L^Y��X����D�[͗G2S� c��Pw��� ��k�Ƀ�d&U��R�T��YS��ijqШ@ct�mn�v��{m�-�c����<�-�����&֨��^�E�ɛ`[���,���x~u[�jd�ޤ
���a�?s�*�w=�3��ۇ���!���0e��ї�f�y����W׹���Ʀ(BU�(r�Z�9/R�sJ��m�t[����:�8=��2��[j��u���v�z�3ln
���(�|��}�3�v����I�yk�����i���V�gA�-ï��'��'a���!�o��c�C���;+��x��t�WoQ�dR��[�&�.̎.����k����1��ݔ��/�B��x-�-9�ٙ�17&W1�\��2u�����3����W�����Z���W_k7�բ���ou��� i�}R�8�wx�ۡ�`x�5��u��|�~?���xw㏸���V*)��
& 
�b$�B���J��hF�
i0�0'�{�km��6B����b�TK� ������؝��K8�r�6��̝�:A��Ѵ_����w[�_Bۣ��HA�i	�[�]��"Y�!���d�{d�9������c1������٭����wbf�1Ja�YA
�h+�_,�-3��Vg�����^����=G��XoF���m֙�j	%L�geT<�q�j#�6-=�������c�.����_3ש�J��z����Q���q�=�N��lr�5,SI�J��Fc׭��� v��Ι���ݾ��X��HM0�O2 _l�+%W5{�N(r�d^�R�e`J4��k�-���×&�M9d�9y��x�`d�D�f�8.i0�8H"��DJt���s��-��QzQ�����B���4�����k}��T�?�(f�^���&���BG��>Hf��x�^��T_s���Y���z9itE'+��msj���y�XE�Ag�=aȄ����S�\ќ�7:r{oL7�0�jt={�Z~Y��	z����&�5l&�t��h�X(����h�w�7�R���vӓ����w~�-�Z��}�2k�*���G�m���;/nϽ�!hq���9�I���~��e�%��;X��z�Wv=��̶J<�f��.r�EΈ�:U�Sv�.��޾�*�J��\��츺��~��	�4�!ACA@L*P4�JR@�R(��0a�3a�oxd��ݖ�wp
����:%�{ ��7X�5�v0�/�R5�=x��t��;|b]�h�����y���+���f�s��j��u�ʩ�άI�Lj5mza'�#�o6)O�T�6`�k�핵�×�B&�5l��h�\;6�p���4:.���s�>vq�jéL8�V��]>�"b�X/�Ug2Vk����.��A�����^ǎ4/��W9����
�����rm������{��0+ܚA�*(��1�Q{�9�C�;V�&9���A�v* ;S�^�M�[ݖC�^ýT��)����o�����P�-?P�"O��/��|T���W�ؑ��ю4����ο�9�e#�Y����jJq�jD�4�o�i���o`D�ݽ>�v�5����oN��_�_�-�<MG��Ŷ���q^Y1jd��Q�g�ٶZd���72�o�U������r���O�@�}���_���W��CzO�~;'�����V���Ξ������%� ���VT\9������Iq�1<�+�Y5�\��A��y��ۯ!8�.�5�[V���O��կ'�J���b����KT�ɓ���ꏨN���`0]s�eG۫���o��gV��1��KvnJz%.��7�P4�
��U�\�	�Wt�t�q%[��{�p+w��e�yv{�{�Ew�Ïu�g��Ԃ��A�߇���!BP4-(�
Ѕ Pf 3 �n���:�����P�
Kw�Ɇ�����)���~~��D�����{�z\��e��o�n�[�[�Ӽ'<R�jĪ)��l�	�hTN7�H"1� ���M���Ğ]�h�^-p�7@ZR� i�I�b���(�%Ɓ�8^���h�
Ә8�7��$��;��O_f��zBuBzB�TT�Y�I��)�E�gܷ�F׎�s�Uv�iJZ�O=qi����5�
���60����w=	��H��i0���\���j��^l�,{i�����ϔ���_NI��<;�B���=y��/1n��[�О��PjEd㋿qTXK�6�q�A���`�b��B�&�C�sS��p��t[�0}ng���mZU3��o��՜ LG֫��L�|c1?޷�-�װ���*	p��si{�L����p؜���M7Ŏ�]keN�l��]�v⽪��jĕb�u^�'v�=0���e���Lw���{��;GLmLu�v�dv��`R� ��o�M.�άoK�H;�Xqx.�v8�	�v�tE��ye������ۯa����[�p�V��)���JO�z�?E[#w��A�]þ�;�Z��ʌz�z3��\���ʬ}<6��jя:�Ov��&6ޱ����^����^�����.f^Y�:�Yɝ�s��A�����L}v���}2zl��+ͭy�������j���)BJ� ?��~�������K�塲+��}��|aQ�8���� ^E��Zd���J=0�M�d	.���r��N�[O:\Y�'I��0K�g�E�S�I>5�mc:>k�[�r.w]�xݖe�ѽ�����-�M�S��z�Y�L�0Aaa�qb.��o�-��m
d��>�������j���u*<���ӌ'�1P����|��m��c���u�s������i&�5k@uT�j�%6�)�L��+�=+������z���)흐/m��`j��3{I�^��ZP��k�E�j�BS+�S��R�&��x���w��?�}ÿ~�U>��խC7q��r�w�Bk�:A��� ^��'�ƽ>�2�����g��iL���< ��b�	Y���6A�~�wn@~���1	���!�{�*�f��يN�_�T��V��s��4b�f��TԁJ�����-A�6�M(fƟGM�=!1���Q�)�N[�\U@�]�\VֶGw,���Z��气49Jw�\K���|��2ml�5����u^?���W���k�h���ϊ�y��p��V��.-��r��T+�v�j�S*�}�e�n��'t�6j���8�����8VeF�r���{,�8��u�Kv5x�����f�\���i��%����G�K�	T��k���8�Nxw ��J��T*l�.��?ʪ���x0`=��V�:ձ���l�o��P�IQ����d���s�Y9轸x��������k��au.����������]SS.�c
�ҵ����~m
�Y���?gH`��>(�w�p�78�jt����~��46�_�/q`���Cls�U �ọ���)����iܦb�������.}{ݻ�{~���S��0��B/ Cξ��t�Y��o��c�x��'�K��;:Y�=*�U�i�l�����nj
�;���\���t�4�ͬ`����O�=I��;�ς�o8O{�����J5׎��2�҆Agkd��^=��
����^r�2�I��C��f�$��B#ߨ��0�6e��-35B���������m���
x����������=������W��l�l�ʖN0-@���l�zǫxU�N���n�����{v�70d.���т��{Q^��D���(2e�%?J����w6����}N1��g3:�^�V�]'�xРd�K�	!v�#!O6�B	�xr�d^�Ji�������~�ǏZW�`��"x����Σ�r�y�=�/�i��j����7�箈Z�^𫮕��Z�u���ҕ��X��2��jQ�W����q�<�ֺf�@�.���L��[e�����@�BB���p�ޱA�;�w����{��������{�a&��ۭ�\k��Xk�e|���b1��<��]0X/��$_I/^�N��F^���-e��]�3sKJ2��[�F�[X�������W��a��D-�m���ʰ�0V�8F��F��:�cP�pL8^ޫ�/�Q���(����Fl>�a�B=D&ؼ�<�Nz���}}�kC1M��1)v�0���ܢ����A/^\^GR��?cE�2t?Lǧ�����Wo`�,�>���^�X�k&�����vE�jF�x�YPK�O���Q.�s9��f�\���P���B�`�^a�?z�s��"��j���15qT������{��q���y��7�5�n��O���na�n/��О����4-_�Ja�������r��)ꝅ=��|���9׍��#�9�Pи��|��0�xx?T񬕤 ���r~5k�vn��B��Gbe�0��e LW5�1���/��ϡ�����L,r���kP����Qs���1�5Pt�1gSy�w�y菌����qt��l�!���)��}�2\jؗ��tzf���O�'>T�e~B�sٞ~��yn2�vgê��cޫGSr��~�0hٺj�Az�����Tu^���|-���`W��씹}�*�gx��X/�}ݒ��^i�df*�M�_L��z����o%��x >o{� �� }VO[��!K}��b�i�oO����3N�<��Jq�jD�4��Zz�x!7u�7�[ѽyػz��tN�L1�1�x��I���������"��<���b�qk�ogv^��'�3t�����r�T,s0?�P5����z�~���Ҁ;']Lwh���֦S<{��k{yiC�V�Ҏ����z�>�z��'BÞC*9���O���S�	���9	w�m*󽶈l�\����D�*�
e������!�z�Pe��^v�O�Y�ޱ�/i^�z��,�!�y�PQ�r�	��V%QN.�l�G�x�ho*�L2�XxH[j�o^������7+2���_v�4�2��|�(�%Ɓ�ɫ�>5��eג��-��A��~�9��!�z�!?T�9�m�N�c��;�G�^↟f�2�N�+�W}�?4�՜�+.OB�u�;�:y󇶟�k��7cק���5"N�¨Y��C֮Qyq���lÕx�^ޞ�miP�Sâ_cX�8w�����Ǽ�s�_\�п3n+� �G�U������j꼇̷�p�9���:$������O$t/wc�EX�NQ8h�s���_�Ů�º����fɹg/ko�8����L7d��tIo��g_{�8����|��Iw������������k�9��q�z	�`�72B�����]W���U/�U"A����������?���������a���Lf�*��֯tz.θ`�Zz�1�?��tv�,���}��J=�Q�+�nc�E�6�t�{A/mbTs	����A߰t�<��#c�̪�g��^�m���nްc���˲41Qa�XR��6˪��r�i��R�ǜQ}/a��ނ%ۻ���A���	*�3�ݽ3�����Dk���HǝXޗn�9E���e۱虗iD[=3i��՗�����لC?:�xC�J��S�
�m�287��a��!憙���!r]a^"s�?�����sdF������|�}CX��=b|b�'�+S�Vo5����BQ�z��	��{������ܑ&��.2�5��u^�x���pBN&3&��j1��`́�Z����՝���c-�#�ֺ�Y�(�	Q��K���k����G�Y����c#,��]�;v���vB��{U-�C�Jm�[�%�D���"���zǫxi�=�����=u�Ci��uۛ�%k.q(>� ��|���L��)���LP�U���u��g�����x����w���}�w���߾�.���y:}g:�`3��n�j����ue_�����xՙzV�E�����C����!�ψ+r��I��r�J�!�R[����{�U���E�<U��`>�jj�eL��q���w�P�4��	LD��W�b��\`��(+��r��,�j"
9nMmx��Z��_Z�U�s����;���'��fY����0� >�t&�Ŋ��΋���g4L�D퓗��l��ή;�=��N����ey۠!��w�jT���V)&F�S��;��r�l�θ�^M�A(�]}cv����w3�麰���x��ɵ�O:%4���ݸ3�I�)#j��z��}�&{փx��{7ۡj��B�V..�R��9Om�M^`ye��|^�d&;��/,������{n[���,7Y(q~����6��`��ytq�ͅ*]A0�|j��5��׌��*o.9�q�]]ٙm���d�/67��$r_c���@�Sa��[��ǣ����X�z�ҹhu3�L�g]/W��敍��A}W�$N����Q�V
�����u�}�MA��n%�i�H�Ɣ��]~��㚕^��9a��Hk=k�L�;��/>�x]�dڡ[�R'�G����TOl�u��9E.Or��z8�P�ޓ|+�y���⹕�wJ��ԅ��o���("kU>�2٩��_m
��;���-ڨimH)СCf�|{�C'�omY;;_7 �^���4v=U�z<��e�H�ޞ��3x�)�q��K�(^L愖.U�֫Eн����8�ٷ�mu2W;m-��%�uѼ�eœ6GPP�pQ}r��q��҃&+v(��Vj�;|�=���J�e��Et�R�+��hE{G��خ���|^E6c�4&��ny�˹��E^��z�Pn/d.ګ&Kz�&��4NUr��0�ʏ���<y`�2r��F��4�K��2Һа�ANe�L���o:e&�o^�c���b,ƭgEưW*T��>�e�T��s�9V�\�^��9����>T�+�c�
Ǡ)�.�v���t�Y��ə%I�y��c��\�' �d�Z�@�y���Fennb���y�^N�|%��L�S/8|㷃��P (� �r/�+��mn!Vs]5B���Ȍ��k��`ݸy"w��NѻE��A��,\��7�+�Wwna$P:ܭ,ۚ��ԥ����7�z@n�t_صZ���M����۽J�s�k.�c��D��Q�˙���V)λ�<�RC�_.��RW�k�˦��D~�����yh��1'=>e{'�n|{&u�Mr�U��\�Xd�z�ğH�=���7ސi�w���]}�o+�L�\`�Gb�b��eoT��f��Ye���S�u�������b�G�������2��hn��a�{�<�'iY��vwQS�m����|%ʠw
�#qQ*�7φ�����K>��oe�$�6�C���Gs�|�{*Y�ꥎ(�M�>��7H6�Q$P���/����>c��h[m%�ѥ�m���i��R�8�ZN�4l`����i(:
�A�n1���n�:b�F ���4D�U~��pꨥ���+v^��������4(j�rt�t:)�f�GG]h5ѻ%�GQ7c��((mn�OU��=A�Ĕ,�F�b�֍:)�lEwm����[�ZA�M4Q�����v4�M�2U!/A�1N0�;��S���U1��MWX����Hh�cn�Q��9��ɣ��l�Ѻ���kmA@P�mlt:.5=��)��[TE�[m�SM�]ݣ�����
�u1��f�h�I��z�6Ύ�lA�u�h�ptE�<Q[�n)�A�.�*
����T\k�v�Z�ώN0���2p~��B�T{�����yf���!���n�,b�`�:��0�U�����s's���#Z��k�ӕt2��?L'A	��������:<�T�ʔ�J���>�A�:��+�M<s�|w�!Ŵ'D>W�����$_��e'X^%�u��*���r�v�su\B����ٓ�+� ��S��'���!;6;����ƽ�H�^�I�l�'L��n���$�N������(�S*�iۓ��m�mvM((fƐ#�&Ꞑ�װ�
'3�6-��W;�ʪ���E��;]V���X*�%ߚ�q^����d/����]���M������tp���*T�Չe�ßZ��3`R���@����a� \����,��"�1n���|�>�U;4Ǯz�[+�%X×B�⠗�[=�Q�>W^�H��<!x��:=�|�y�.^���:`˄�r�vN��ݷ={�ln
����:�,r�N=q��ؾ�h�ˢO�Ƽ\�xn%3j
,3����D"�!�_ƻ���l�m�_J/��=$;z�k+e��c�yFlm���!6�(�I�ū�4}8������">��bk�IgY���2�77�ջ��
���a��C�4$� ��N�T?c�=� ����'>ou4�Z���w�a��������G����W۳�����Y������������ɃGD
�jz
�^��=�=�}W]4���i"�=j��F���4�or����k/Ix-�}��L�x,9%�[�:'�.�* go��E]]3�(�K%�e�o����< �{��OYͲ!*���Y�s�ʇ6nf��Xu����p�y6��r����B�.,�ف�Og�f�³P}7��4�v	E�\�⚟N��E�w%L�`�ʂ������l�zǫxK!#��&L����XOOn!.��؆\���U�����"So(A��i=�]:®�[k�s��oNj�˨�~�9f�}\����kc������@h������N9<2�Ӽ(�t�����:۝݆Z��i5���@s�9Tm+y���<��?���1��{�6ͼƛ��y��ն]��*K�u�)��Li#I��ܞj|��\�p]��!)f����E9ؓH�mt'7G\=��
�%�HJ�$��S��<�Q���9��az|�>�a���_pB��ۚ����7�ݒ�!=(2��m���R�e�szx&i�ހK�(�M0���������V�]N�7����hP��00ZDO��lK{ʹ���:�f</Z��a��Gs�O��9͌Pm�m֫��=V����ga�����D;'�S�+�A�,w�M[]�L���#&�k���p��6�y��gF�h��Q�_����^)�jh~c4��;«�xnm^Ɇt>U,rXʫ�n�zg�{eY�.� T�E���m|b�5�f�{xL#"��Y��z	;*�s�c�{t��3���/m��J*�c��d2�ɴ����`<�o.&2Uޮ���l��v�; �A_�?�����,s\���V�Svd�ډ�my�}��1�w��n����Ⓟ����/��!ݺ�����~��ӞT&�߾}.ſ��Y����T���+�ky°�Y�_��i��>��и�x>~=�1���4m?N�ɭc�ݻ�
��	2cz���Α:8�j���c�ĝe딴�C`�f��a�sЕ��y��v__� �C�ѯq�\�m}�oO���+L�vJ-�m�&a���=�\-��.�9r�s�ޭ���n�ڪx�.�	��cqlK�~���vk�2�H8@� Ũ�Cc��+�3G:�]=��yP{eu�,��Q_.1-<�A���f*!;c�}�5.��Pڴu�j`wob�������9
˟�z`ײ �����*���`�e`�.6�$�HFu�UEV��4��*ETf4^m�Fܣ��؎���N�-T)\�,)��rq�uEê��x ���f��kS𻜨�[{x����vX�����,Z�D&I��JrR�Hʢ�]��0�v������|���w��˻l_��C���Uf��m%�7z��O5�yq��p�6�[X�uW3ҫ��D����ؖ%��'Y]R#��A}��5﹗���r�+X�h��R�t��2n`ˈ�ӝ#	f&�v3�vSd���&��qs5�kT��}��U������e�Hv��`�{��>��г,�E�i��T�ax	��y^��@ߣ���۹ق�E�Lc��]�y�I��㄁�0�'�����fFʧi����lr�d]`�s5S�6�T����˾�yN��zi;1g�`�؃��"��z�I͉7B��a�ª̮xj��\�7VC<[ܒ����M��2��;P�3��W��Xvy��6(��	ι}s�B�1卩��lh����3ً5pw�y��x�]}ZD��OA_�@���Zz~!i���E�*�f��{��o3H�+Vд����V�����Q�$�'Z�PfUԡ��;۾o���]���ese���;/�~�ڢÚ�0�@��6����8Է5�,� ^�9���P��n�΂%��& ۛ���z���^��2����;+�!ug[�-m��7 ��Ϯ�˼ �N>X�X�����z��߂��<C�\�ᧉJEQz����f�Z��=0ҴE��bm�lg��`L�\Ln���~q]4]��}�_����o~���[w{�`�o�����v�g���z��Om f����].y�ga���#�d�d\<uY�~/_忧7jf���5Q�Nq�M�OV#z���QQ�O��9�Fs����X�5�#Ge�z4�Օ$J�[Y4�̔�vN�R�2�չ�3ͣ�x��7���glu�Sk�7C�7(!�������My�\e:n��u����9aV'"�h�,=�6�b��%��	��C��vf�$�.{��A��B���󇡧Ƶ����΃��QB��k�A�]���w�J,��k����ݳ0��Є��P"*�d����ƒ2�!:o]�?��7V��G�[�����AF4���LD���"�O5t!)���)͕)�j��k�un�q���h���^~0z�he����ޡ�F��p/B�p�ޯO��N\�ķ1�0֖�S��+������=j��(�o0u���9nG���|�����*���g���w���r^#pC?S��ywvB���j�Llx��;.˅��;���=4y�� p��1�Vb�QS{�qV޺W��N�)�~���ʂƵIw��\<x��?��M����2�3��K�YG���PPԄ��s~�6��a9W�kUz��f�P�zY�KӇ���1�n鍾�s�]n�е� �ǡîsBvi��Ije�N0�]+^�A򸮾|g�P���g
�>%�̛U3�mҺ3����Pn��e��{���&����2�;K�V�7���s���M��p&,�ܘvK�fb��!�>����9h�ξ��nL�u^�&����.����������D&�'�,�Z�a�-0G��$��h�:2�F� �����;9KϪCC\<�E�C��i��mǡczm��*����G)�������)��3�cks.�u����r�iE�v2n�+D"��Gk��B�з�7��7w�E���E�ЗwGS����Ih�7e�1^�xE��Pt}��I��cB�!�K�5}�Ol�Hw.t�&���r��Z�BP�zK��g�E/ڔk�c�1�~0��~7 ڱ5�%�ꅚGN�)m�^�������T�4;7�Z|�A*��d���u��3�҃����iw�g��wN�������F�i�������K���1䥛x�ʂ����R��4Xޜ�ܦ���[�ަ��en���ј�^<��S�{C�h��<�.=<+ʫ%����Jm��Pd�Jz��#��2�����[��p@��1Y���~�'����"�c�
.�d)���'J��"�B�-J�ޢ;�z%�t7�i��F�]���Ưs�:y��xg��(���R�*��@�/J�Mm��{8���}w�|�.�_���䑤��#ry���{�� �5��,��W���k���z��E�؛7����'G��M�ši<�Ɋ�N=s/d	k��gB�7)m��@�"�n^�3��/�Y|$bWsr�\y���;���yZ���*��Z�C*f�e;�ugM\v�lba9��b�1
��:+dɁ����yȆ��B� 1����oo�?j�`fԧq:iRO�1���F���Ǟ���WY�J���B��9ޟ��9J��Ö�9$7PΛj/xT�O��n�����O ���#�D�d���)!��oOM������_A�A��YՒ�f�4����п�����Y\Q�-1�z����:T��/�c;C`)`��"���ί�dS�j��L����]��}�:���>
�?����)}X�����!9Z�"vdง�]����N������hZڼ:b5�3Wv޵����X`/m��%������j/��:��a���`6�)���k�rzo��U������ˬ��G*�?9Z���I86�5-���Z}�������e?�o���+-Q=�
s�C�d"c���ܷ�??9�&��j�.ŧ��C� �/^�x=7�v�l���[�Ԅ�zAĴ�O*z/�tö����Q2��{�PJq�jD�6�fP�6
ۉ���ʣ:_�ߗڥ����RL`�$�< ڳ�����f�kR�H8�����Kq�k�Kj���?8zRݯT%��nEw�����0��ٲ�h�&�#�oCl�AQIa^��*���ⷷkRq��:�e��L]��Ӛc�ㅎ�V���]�#�;Myi�ط-~��������,%	�&	X/M�]3��ݷ� 62����ni�ߨ7��:�Y�l� Y_)��v����o�?5����z�R�؆Ǒ)�d�Bڍ�A��{5���(@�yd	cA.�g/���/P�n2	�б\e	��j[�Ϯ�LٽyJ�E��-�����e�~���Z�R�J��}��z�k췅8���z�J�Օ�ˋW��Y՝s�<�S�.�a��t�=�'�b%9��Z�TS�}�a��и��<�̫q�/4�l+��7�#Za�'Ѱ�*��f!�,˴�I�g	�ց<��H�d3<Bc؜躇�|��7�'�V:w�xa>YB1�C���OH ��}eS��Y�I��M�.����Ǧb�љ�wJė��"uӿ3���p����x��}&�Q�)����׽�����Ǽ坓$��/r�\�a),h#�ȃ��%�����,;_W���yo�Q\볷!���v��wKu�ss!
+��q��J�
���fT�OtZ�����9�����T�/��ڬJ��\�{k;E,jRd&�UVJ�l�V���%�	Q�'�hN�{�=���[��O��q/d���	t{���B�M���cg��M��7������ǆ���q��2���c��Uˏ��s�]IUr�v�gyY.˞����q�eP�p7����(Р�8EF-��F����e*yٕ&P�ˢ���[�z%e�O���I�z�L���>�ꡔCx���ut3G���}�o�lk8e�sӲ�v�u�0�@�.�Ǳ��+�KsP=��m�n�>[��m�}�7
k�Յ�!�:�"w�~�9.�:��v�ÔXW��@q�n�|eL��@���(ke�^����s�)�8=6��[9yחt�������a������"/�)��ǅ,Ž�j�{�mJ;s�Ў����p=2��6�ƶ3�<	�PBp��F�{
�s_2fĶ��*2�mn� -�_p<�9s�Y!L���]7t�îyg���}�P4�|G.���nwNd�׉}i�UKcR�!s�;2��B��G�*ޘD5��E+�g:̃�ӿ�n�۵��s!�c��>;W��1W�R���D���!2X�J~�h]���~�m�˷����{�ͽ�t��s�<;b�S�A�0}^!��ss�	� �JseJ`�����)���Qy��.����5���������$8���ʗ�B{����5��2���O!�6�)Q�/�8���Zq�x�%L9�/�S��'���3d�!0\��ư����~�f�i�!�Er������z��3�ςe�=oRTt���7eK�e=W?o�0�����K{���]�4>�}��Ńș��[��W1H�Y�p%#}G���H� ���w��EM��d����'��W'b��H���P�C[
Jܲk�����0��գ��uf����������k���x�5�F�����-N���� ���!7\�L�y��Wm�{gw�(b�qJw�ʮ��j-?5���U~k�q.��#��r����;�b�ɽ�����i����P��Nl��Մ���Q���9�R7]�9��sU����p����5]7ݺ��%�w��yís^��M����W	V0�r�Z�T Kܽ��sl٭}�!鰛��鸴�h|셿0A�a1�}�GW�bGq`�6��Rca�u>X9
��ѕ��Ջ�N���j[r̫�,3����p�4B.��/��
{Bظ���e�*7��`SVr:��G���M������0ū�C���I��cB�!?9��-E���x�UZ��.r�Y�*�f�0�����8OT4��-ĳ��~ǆ{�Z[�_R�KdDO#}g-�4�R��s��^=���l�_��KJ�!�0��ɴ��6��-�Yy�}�y[XaWi���ء�x�֖!9l����5>�{؋l��n�vPeAd��
;A��/O�������}��o������s&*za��-,>���+��@��5�o{r���Jts++K�C!=�����*h���"����2�d�[�搕�+E8JRɨ�<��G*����U�)-��v_ d�pJգ"�w���|�����)%���P�Lޙl��I�]���G��z���3�@���]���'��n�G��)~�󨪵�sJ�0c}�k���U;R�k�w�Aҥ��1`�]�M���+mm�����������d�Β��%8Tݙ]+�u�o���'�A���~�}�6�Y��[z|�7�V�e�mZ}����a�LA��.��i6�q�w��a�U�W�n2B�H�y�����$��a'���Xs;+.ꜷ]�z�˅dt<5�7R��<�Ō
	��g�1��q���F��ڮ^�O�tL�����M3g땘���f]�9�XΛ�T�v��:�K[���9�s��ad���=�n��e��ǫ��}n2��7(�b�B��1(�J��pz�T����P/H�#�㗣׺ob�gZ2�>~쭊'���E�N�摜E+����ֳ�P������㝥�-֠��ŷ����Xn!��l�b��'n�|�S.MW�-�̱���"��Wf���,9��[ȭ�k� F�
�a4��<��ͼ��Q��n�:�w���pr��)��j�%�WQ�w`G �R�+ԉ�l<�&s��իt{�^"�t�i6dMp���e�&�,5���l�e�c��`bq�r�Om�]�Ea|V��G~�}��j;��;�`}�<]�^��K����yP����y
���C�k�T����l�t��;��g2|/�z�S`y�k:V3��Y�Gyb���f���GL�Ֆ�]�0��w��z��N���٠=�nM8z���CD�W6�Z����.�X������놽4���/�����h\���#��}F�w�h=�~��.�8�vk�D�.�چ�5��^R7�-�GM<ݹOIˬ�f>�e&�,��B��6덬�3�Yi��ѫ,I�1����+��/%�J�o�l|�]*P�V���/�@�n+�j}����1�ZSb��2E�C)�@�ǭkX3���I�G��n���x�bV���F{��j̬pS*ۧ]8�m�q������G��V��q`�j�K�WC;`�);Iౙ����re��ʹ�|	�w�OG�p�ɺ����+�U7}y�%/��}uZ�xF@��AV��:n-�{t ��&���M5i��v�b�������<���M�M֕{��XcU��(� ��9�\o�Д�c����W\�ʖ���5�)�M~�N��
&�.�ܞ�GP!f��h0,���s؆V�Ң/O��^���)ؐ�3-�`��7�4KT���j��wF�sfYu��tW;/�۽7hlg"�Xʺ�N����P��vCXz> ��yᕰ9�6�v�X�Ӈ3�m�4��%Vp?T�׎����f5Ӣb�{X5UQ4�Ѣ#�����6ŋWG��SEEGZڱ!
q�TDu!R�A�*I��)�EV7q���lS������ձ��Tm��RT\c����Ln��'v*�*���T��M&���E�"*
�&"����u�Ӌ]=A�h����V1�@F������w����+ZtTLU��X��A�u�-cY#[�htWA۷t�j-�����-��E����[gC��F�E�����=	��ƀ�UGlOv��tQ�u��uƍ.��Z"���"�qj���/v�	�&����Tm���G]��6�Ţձ�Ti*��֌lDln�;e�n���DV�Klm�SmZ������~����y�w�?{�w���u�`��y�*�j�7'k�
��\��W��o0EZ�Q��:�m�n��R���y���/���^�ސ�YJ��kռR)�j'���𠪱�W�H�"Sm�5�^jn�������u���v)�R�u�ј�oV�^�F�̅$`�ar"!�v�����E���e�V�����Dc�/u�)�W(����fՐ3���ZN1��<�X����V�V�cAi��"r)V�=����*f���D�7�E1�$i5��:�?������v�Qط߻��g�oP���TܠʱK03�2���oR��E'+<�T���5�.�q��������7�2g1o>o`3�p�G�9����v�:m�>�-�j~OI��A/@./#��tg]�z?]��U��V�	̐��1��
9������j%��3�s]��-�R5�:��0�љ8���m�t��^N]�O�K�GF3��!�:X?s�;'�"y։2)�z	�k+T����pc��͉G��xq2��T{��l�v�;?d��q��1��ʄ�~}rnO
a|���#3\w1Т���ÇӬ��\zs���j�}������:2!����S�7��AKecC5n5���ڻaOu�٩Z�)�8���6���4Sx;ƿ��b������o�+i�F�qe�ȼ^�~������Z4�lf����Xx`�w�=�
�c���i�2��4�k̃i�ڑ�oK�ya�\���$�gCᳵ���&G���UTכ[͵�ww�l��w/�aT#��i'���qh���o���-^/a�G<3�B���$CL�^�}ݽ\>�F�1�X��;#[��P~ys�M3Eی;�h�C��^>�+�[�h�s��w�N�H�T���"]���.<:N��Ӎ��=�>�� 3N�:�R�d�������־��l����/�e�E<$�`��xCV���r�~����J�H8��.̝p�����^�ް��Cw'�Q&u��l�,qL��Þ��x!'�|Ǧr	�ۓ-�79�[e�َ;�۹|��_�����A=�%�լ����e;k��O��.��<�;��ݼ#�j������n0Z��Fy��Ƀ�]C-~O)�U
W*�
j[��^Qp�1��KFSkm�[+u���
���f�/�W�e���Ib��L�ߌD�6
T-\�;�3�%�X7^Y�5����.��e-��zB�"�}2�/����M�m2�2�����E�4R{Ά�]���}�ڞ�����	e�D�bF4���Bx	�a�,�YT�f_�)?/Ǿ8>�k�ѿY$�e���]�d^{_p�9���;�g�s���k�`wXS�y&=�;g�`��Z�����י�����[wC�[����G{%U��;T%vt՗m3��|pc���Q�ܡ7�Ն�A�����5�W
3y�"�d��2��z��Wމ��V��Drc�vި�?�9�_�i��o(6��W*	q\���`�݈n��=��NrNP������sh�^�,�X�w��B/<
�����H��1�\Y�,�~.�c�y^�(�1)xS4����U�`Ԋ(:��.�E���c&�k		��W�=�x�����7�[p��Zss����{�YB�eS�m�B�(V��X�����A�Кx�K�h�}�PO�*�;7V_B�fr��sS��v��E�5)P6˦��r�L3����w�wgQN�*�l�k�7V�j�R%�04Ba <F����vI��zW�έ�Ê�N�w5�.nOL���r�Ӵۡ�e�~��g��Y^Pj�?������S�Q��0}��Gw��L�wvJf�Yg�G����H\���H��I�ʺ&�׶3��(=����3]&�L=u���(��k�����������#���PDך��^�l�.WE3����͆�v��ؼ�[�`�p�bqׄ�cV��5��!s�t+��*<��zq���C����J�q��>����O4�s��X�z�l�Ζ����*�7i�%�nP��ai��/}�Y0��:.��m�C�{Xu}칄9������|�׎�z�(�٪��vA}����W���ȵ_z�ӝ���s��CD��Wn�6>�ɻ<p����Y�"cHLsH�9��c%�U-�W}DZj�R*X�R{��B����~��QR
�=��k�Qt�xj���0���H|��Hg��x���<��%2��Nz�a�蔳�_p�-aGΦ
�w9����_@��x�������g'ɾp���k�]uyu݉�^�^�m���G\��-(�ƒ4�W�b��]D'�}iٲ�B`��OAE��͇e;+6�m�#��N-C��n�X�R���Lkغ���u9j��8zhAC64�
:���
���r�ovHZ�	2,U"M�N�H����='�⠱�5Iw��\<��w*i�������;��1�-q���9;4�_����I�qOC�}��#u���ק�i����lj�D���j����`�
=í~�٦�bz�[+��P�V���˵�.�(�2+��|oqF���E���f��`�>��tA���k��h���<z2*���X����4.�b޻��Ҏ���}8�L�5�,Ƈ�����%p�	����E��'�|����E�#ѿ�y�Ώ�{Hg*�ȑ5u|�!�VB�1H��=l�:S�Owt���$VKUp���I��L�}|�mwe-�%�@���p���K[-����y�q3A!��*<�a�*�)��C�L��.�9yA��9�׬V��X�'U;��P���לS���������t^���-��LW���������I��^?�yw#��eh7%hvL���(���J�u�=���A��6��6�$>��@"Iꆒ�-�>؊��xg�Ox�>�R��k���GOdwZY{D{g�����^=����3p�4��è%��#&<�ɴ�6p�a�irLj;����S�!O;��-- ��22����y�s��mڦn;2>Y8����w��΍F�᜻]{Pc��r�3�a���AI1�.���Z�.���>�C��=[������0�^�q�e��dl�j��M����MwG���}���<����%���C�����P���/;p����[�\$�ȿ��(FSS�[�����P�^��d��"q�S�(}�X.��wV^`p�bqH�w���<�7�R)�$i5��ܞj|��TG�����͈�����]����53s(�,ʧ�8a�-�)�N�T�ሤ�`�El�n��8!>3防��gt���#XG�"=�&ڝ���M)�aR�"�6��Qi�`O �`y��r��ҚڵJ摌d�LYn��Z�3V�Q�z�
L�E���/l�����`Z��$j�"yʘN�s���T7l��1N�e&8Ԭ�a\�`;oU��n���e��ƒ��<"N��=]�g%K���f���U�be�a�V;�U���^K�K��7����>a�O�(֟��X��˥8{s��7y���f�|WD,��;��+��j���]�q�K�GFCc��rD��Ϡ��𞂏��ۖ��VmuD���o+b�<_����u�����'+��H���+�q�w��;k���Y�g��[��d�^��8rEr�L:�ƲǱ�}���/%�1�m��Pwn����>3&�Z���H��uv-����WK��*D��pl23L+�@�LW5 _�9b�8 ���&f���o5Vgf�G�v���3�����WH㕛�}�<ҹ�0r�#���e�����\�e�כx�!< ��,h��8��}`N�vװoO�K���L�3�ڷgUwmll|ݩ���c;��Pd�h<�E�3����&s�|u���,o3�_���5�����p��3���h>͏ԩw���vq:,P�sP+$�(�5�4>͟����
�A�߭�4S�)���DGd���m䆅=�{]չ���:��x�����i�	�x��g�o�YQp��fA8����|���!�4�y��pI�[]��l���y�����y��A�k�I��H��ֆ� N�g��C�z��*7��K�.{PU<h^i:��+=�t���ӫ6,�ֲ��m�:E��w��������z��|Q��<	�%���}�ܚާ�������	��0�y;��&4��Y��v�no�L~wA�>��zm:��B��UԷ'�T]za.L֩�rg٭[lz{yS:����3]�^;U�p�})�W�!2O`�Jse*�IN(=kT�mj���x�i���}ܺ�s,����z$!��q>��W�����|e�F�T�p��mX7Y�!��`\�9�{���dU: ����/^w�xa;�A���'��/X`K*���7&�uŅ4k��4S�':�%�����m�u��s-灺vk�����\=��Ð��Bz)9ycoo]oT�u��9�w�8�4�aT-J熵P��{�������ߓH����P ���B�����!��M�C;�W[=��؅7S�1I�ɺX���O0^���f�J����MV�cP ��4�}-|1�Ӻ���಼��-�0[�#�c8е~u+u��Z�9/LeG0["5��:��I�.����;��[�}B�0p,G�� ��}�9��e�3����C.�Ǳ���=����.����?� ���g3�"]�Z!0g}�뜗d�XޑsW��׾���=��ʊ���v�C6��� =ٿ��R]�5��߯��E�eR�I��|sw��´[!$^j+k���g09�e��]u�r�CqI��t��@�+�֯,�o\��7ԨǨ��ڌr�5G:f��:�L�P�Hg��Z9O��ٷ��v��_��s�;ky��hv}_�sW����/��w���)��F2!�EX�/A�:ܭ�|�'7m;��+����TD#��hv~�j[�ځ60y� �;�y{�n�Yy��j�i�͕��ME�����y��v9��B�My��)�WL\:��L�p"aݥ뵛{5����gA-^e����̚ǹ�ƣyU-�^�R9�� Ȫ�R����8�.����*���Y����S^�C���?��4G�w�)#_t��{U-�^Jm�2!b�I��钱\5��_FպݮB�Fc��V��Ol����H|�0���j�B�K\�B©�g��
	nUoQ����}�oN#ƀ{�a��T5n'�X��h�N�|�pB|�;Q�v�q���k��u׼��������9☤e0����*|�֘<�Ā���\��m�[�$�cZ��]��C�H�V�;Ϭ�'L/�(���Ʊu;uNZ�w���M��TIt��Q+��F������������e��J��U��ʮ��j-?5�T4�.�Ԝ�����5�����n��VN�����c�|7��!�����/Cv3��i�h��z�xs,�ଷu%���1���P+)�����0��M1+�{�۝��T��a;��ᮭ��{tF�%�IU��DU
�:�
����+Fئ��-9�S�7��%c���S�ۧ�q6�fo�|���0tŤt��cs�X�����	�|Uz��f�J�s�a��l�m�$�ӧ{n��!L�zp���"5��ã�9�ꝚmW��-l�BU�+�J��u}:��j{W'�gӔ��d_W����'yQ�q X9�����k�5׏W�6���8SdU�ޔZ�gO�V؃(�|���q�q��v�׋�Q�`�AO��R��?)^��z��'���9�kvh�����xj��fԢ��}��i4	���9j��ds�0>�5���M���[����Υ�}z[�OJ׹��~X8�s>ͬa:`��Š$�CH/���툨~М�=�����9��yG���K:F���
}:��{b��=>�ǃ��S���4�5�%�%rF:<)�Ύ,�>�lGE�Ta��~_~��`�1a����d^�P~����%L�`�-�7U��D���noW-aL��3f��ǫx]]��k��?��U����57I�K0OS�
�{ۼ�!\�-kT�=�WN��=�1P���X������"�c�
�>J�O^�����m)�}oXF����睧����ǾR�]۪�]�)H\�wl�C"��^C0��;��5��Ë7=���/��}F��
���ǥ��b����6K%;�Ց^���_lO�Li��V�������[��8hbb�ܼY,)M�#����8y�&��>}힢�B	�Q,��)M2��m5�Dv>1jgO�����4]�u_4ʩ˺�J��V�6�g��唼��2��1Γ�xNq@��oJ魬ܞj|��Q}M����ss1I���G;5�T�u	�A���.�Y��3M*I��Q�+���5���J��TE0ɜ����1�Ϋ]=ǝK���G�M�;<���6�_
�jd؝Qi����X��n`�L�wæ��V�m�t�v��:�}҈��@vG��>zc^�\?r�{M�?k��W	�~0kyA��9~n&�Qׅ�Bn�I���O���v�ь��a��;�'�"yzD�'�h��,9��Sյ�RS�X��y�S�U2͕�n��#a�?�`�XJS�-@�VJj�N�gif��S�&?aR)s�L:����.���<�-��A�=9�U��x���f=����
�ֈ�ƟC���;_s���2���X!ŠvP&+�j�c�q��s�m\`�9�����{��;�=/��#Y�
O�ac��5���A����:�_���p=>�_��������}��o�������!��z�a�*��^����+[AWk�;���1��V$C�7ԱW �xGҺ�>y�)�E~�>/!��������|�6?��qe���-�7�`��sX�<+��F���0��L��oM ��y�ۚ�;��fY�uk�/a��Bno�~�#���褑�/����nq�J/���p�;(6A�Ș�+%�Ao'Fnk�r��H+oo+N������"�:��Z�Ú��x���j�������Y��S��ό�p��;+�%�$���Aʉ �w��-y���:��6�ǥ�D�m\�q9h�%����/5����VT'�ǰ�<t��i�r�[��OX�`��۶A�2�f���f4&.C*�{�b[�p�׫�[�ޕz!���q��]f��m �1�]��uYw��Ge���E"_+��ok�'s�:��ʸy�`'jؤ�l��*4��Mej���u����"���]�/�������Q�j<�����;��!�I�;Ū/]�\z���g��q�}�\�=;W��f?a;��=/����-��#l��r�5�-�p�Q�2?h�}� 9�~�Ȱ����������nl2�n��(T�[v��W���P=b��v��k06��
I��x�k�-.��~���fв�X嚘���̽��T����a=׶�}��s���9�>
"�P�k�sVt�ف=rV�%�"w��qz:<�a=r�=YN��6���^����(�F{�܉7���Yΰ�-�3�l�o�����R�`V�/8����Օ�wn�Z�������\���/y�~�{�p���v=�{ع�-5u�_m�O8�޾�_�yq{[PNP2�WKQ��2p*�}t����v֏�Գ�	�N�/ov��1��ֲ�=��f�F����o�dJyU��L3��&��{��q�C%��zK[���ut�X"���r�]ǧE�S+d�Ԅ�j״f	۲������.V1�P5�.ѭ!]�B���m�b�.G����k�u�>�釨�f��m���%鮽��_\]�9n�u;n	h�T�� ���9��7�z���\�����m)�s�`�Y����wʓ�l���`�:���Y��qa��!9狵mDQ�Z��K�Q`��M�eɏ�)��8aȖc�d�Ӻ��x�H,�.n;��A[\"q_RІu
�z�T�K�Vbv7�m^rD��7n�&d:8�ܽe�H�͋�fss��J�j����{D��{�0^1;\��腻c�8�.~�y��?_as���^�iM��;y���x2`8�IB���5�vϞ�D�,�z'oP��(�=T�G�E��Cܵk����绚Ѥ&�WV�����8�#a�����|%��L�2I�t�5��:������K�嬎�t�k���j,�)���N�m������:����j`�JD�V�ĥCL(!T"�~��(�AC����mPPD��לw�7Y��m�8��F�UOA�Mm����ntcTlVm�`�
�-j��&��F$�Gg���6� ��l��#]=uI5SEkT��DѶu���j�4���Xs.�[j�;i���wh�T6���K��&4e̴jՎ��Z�ZLm[:�i*�)�-g��)�F����9�T袂�X����S�`�ݠ���UGQ��GlPv�iv�=ۣ[[I�mEkTN�h���Tj��Z��	F��zi�f��M�m���Y�n�IOlu�t�v7c5�k:�k��F-RS��V�ͱ]'v4[Q�Ѷ�ň�Ѣ�`�ح�ݒ��U�h�m��n΃6�5;�ض�f��U��b�;hڂ1Ed�h�*-���i����gD!���~��L,K���r��j�޹	���T�`��{,��g�[X�>Ue|$N��mR�8��iT���F����ӣ��`�ؒ�l�I	?�E�#�sz���ˊ�����m�׶D��8��.��訴��m���z��3M��M�ݸÖ�[;��G; ;��{ތ��_,�-?k,A���\["�5s��y4�s�aQ���4g�o�w9c-0x8����VIE�z�l�*����x��'$穵x��B��ε��6z�X!�;�*+��!?5���z K�]Z�@�[�d�C���f�x0؍ٳl��̺��1=�;�P�8D󌩉�i]:Ųs������b��Z�R�*�
e�\[F+ˀ��V;]6I���6��T?#�x�弞ᚰK�N�/e����LZ�!2N]�9�R�j��-k���4wF�^R�s���R��`��gN7�B�>�2�_K1>�2�:iR`n�|�}�Q��c�{y?�7�PW*�w���/@;�0��B1��0B~��A~΁,�)�D��g9��/:���vCz�6�ڕc$���i��mx��=~g�
��!���=���/x�ޫ����{-n�r���J�*L*�.xn�r��PX��u�
�����a��ly�{�h�'�a��cϔ�B��*��P�{��W%f�����SY\��ʦ�;*H:��n�h�k_۬]o����ª=.��SȂ�.g�O$WoA���F�	��@��g��N��^\}��NR�1;�&Q
�}!���6��õ*���Qwq���N���n{��U�-?�'�آ�ě�f����I`@���f�V���A���ÛF�z��:ku�*;���`���,74��ʽ=#�k8���_�J�a�Jײ���������g�u��d��n0{O����5�G���i���ׄ�-ΒÛ�l�k�j��|.6�LV���Y�N�i�MAtO^/a�ɑ.�8D&#m���$����rEyC�E6�譙��xY��ǘ.Q<�^*]���c��t+�j�1��<�,#�z����b\��q�}�$ق�Y�K�ޙvo\s�wE@A����I�ʽ�6�ƶ6�g�q�p�&5W2�ޮ{���M8QFW<K�=6{65� ��; �t�5�\e:j1p���������vw�;qK:�� 踘��OsQ�]c*���R=��W�e�	Y�����u��M6�}�K�5��0���~�(������|!�s����:Y�R���D��P+=NӞ³J�����&�	Gh]��ׯcռ4�{gh�-�!�&B�|CW(�^)������}<���N��o��VE�Vj��Y�������8�~�Y����cy�ts���ǭ,M[<�Sޝw$�O6��^��X��A&���Z�^󦁽�&	�?�B���PK��5&�T�/yvi�`\MVLhFZ�%��wD?�q�|�? �)����^�����x��`�L:*c�[���z����z�#a��hN�>T�����m���k��Ё�>^Jd�X^%�u��)�FSk�B����Z���N;��[=se�����֩��SЃ*�$I�f��يN�_�T��9������K��p����;y�r�4�W�ӛ�2A7�ۚaM�= ����Q�����ʮ��Z�O�eD���R]�:l���^2+:�n�����\�p�N��W�>����n�٢��M��j��.�F���g&��F6T=���|�Wzz��t@��?c��#Xw��^p�_�N�6��-L�BU�V(���-秏3��ޙ�i}��~�\S��~���s�N���a?�S�GW����_���^�b�1IQ�f�vd*b��̭�u>_)��׸��Qۖc@ņv2n�ϴB/����B�b)����f�-Г���vݾ�_�1�IŜu�&+�tE�f�"�D��kxvwFo>�l����Ҝ��{�(��Fmci��$;z��D���>:)~����s�cF��`�;���,�|d��P��9�\�m�^!m)ou�=d�8g��z��a.�g	+5Q�ո+�ۈ�r�^pᗄF�a
��ܽW�
���Ë�:��?E�b߼�P5Ë��j]E��m협c�cR��?�yD��^?�ﾯc�9�?)��a��\K<y--(d&�l�ק���編sO�p�4��è%�t�N�q�ٟn�7���ݿSA}��C�-35B�.hj(M1������y�^��R䩛����n(�/�{z���ȶ�v���'�z��C�S�-�2/Qq��q�GyF5%ke�WW(�Ç7+���"u���5Z����gXP]�V�o	����q��,/��7dm���D?B~��\o;o���R2�3͠tA	�r�d^�J@�P�����C����=���m]���l8swE!��]�����_I/��'�D�65H�4��������&�Qix��y�|Ofv[U.K�z�kg��2��2���ڤ�W������(���6�3"��v��mu^*a,�F'e�Gha�,!�"oz�S��9���R�>�	��t[��OE<�V����|��I�./#�˦�p��0�`|�Y؎q���e��Q-���V
)>eo�$��V�q�/jF����A,Htq#�
"��X�B�Q���_���>5�6���5dx�W�\P���7��^�����; �1���Ku����dOf;�W�+��_��oX'cM��	��q�V�!u}�9����΁���
Q:�/}�#�5y}ě�O��.�������{��c����$'���˓Ca`hqW�n���������m=�J�L�G*����I��gޞ�.�����'(v�;�
���~��q:�7˕�9��T:�;k����r�^�T-Xu)�W��X�8&>���;����"���[i�ִ�Vnwj�;��9����ro��K���'�����hGVI����0�ŠvQ1\΋�I��g��=��NL�����H|12��40|�`q����4������	��;L���`�viǅ�f��(jdGC����ʇ)i���"O��^�|`?�_\��m���>�eNE�.Tc/>�wgviCإs�8�2&!�|kO��sdS�`0&P�oql�����s���h������d�+�!-@���Ft���؅����-�f��L<��zc�{�.�='�r7l��j�t!*9���qt��������z�"��n*�i�������g �����"y�PM�i=:ɫ&=tB��r�N��U
V�,)��Fŝ��O����˞��E�T\9�\c<�-�Pe��^v��n��-��~"S���b�Sc��r�3��]7A�ywF^�W�ʽ��b�V�rt�I�/�f���-Ո��mz[�����{�ywǞ�w$�n���>"�\�7���ge��C��v{\:������nQ����A��1��TG������Mz��B�3|� #[�0fח������؆Z�E8�ض�Ш�oD�#D:A�����Y��=��;Nk�l�f*�/t��/�����y���Qz	q�lGN�;�0����"��S�.�ҵ���X�8ѓO�g'��b��v�Z�I��M�.��s�,n�l�T�ȲB�_�}��h��	�^Z�s4�w*�Ԙ��H���I�W��熵P��%�#�;�0���G�ٵ۵��{���9c>�	�x�u�Q.d���Z���T�X&��]l��;:�,�a��r�}9j\<0`�51L7?��t�'�sm{8е~u+u��JװT�˩��|3:�d�c�r��ڋ,Нj	�;�8a\#��I�l�W�>�4'��m{:�j�F�~<$�NV.v�=���m֘v��MKsW�1~U�`�y����'��AKmu�����{�ȗ���o�շݖ��vN�A(��^�.ݏ^&e�N��5�l�����4=���̮��
P_�Y}��ݑj���)��z��ȴhi�HzJ!������Zgլ���}�u��%j�����w�kKq�wl[���
a-��g3��#������
��֕�7n\5��8.ޗ�|E��?{m�X8�ͫ&֖q�o�#E���'�Y��s6��P@!���9���/o2xV����e,�T[�	�$S�{xD��5�5I˟7IS�o�cB�J�zǦ��֐/ ��ݎG?x%��My��]6���O+MзM۾�u��wr��]��E1�~!�_y��yX���^UKc.P��� �fP��j�:�"�M4m]��:5���a \�C�ئx��֡�`��q�@[8ܬmT�7��m#���x�<wi	nY�B���H�=;�C�ᦞ��.���Qz�0����W���}T}�)�ܩ�[�{�f�c1ᛋ��AYZx�seJ`��O��3j�O�B�$�Y���Y�#_{��tCEн�Y�YxF��ڄ&ҡ�1	:��,��g�=�I�����g8��s	�Y���b`��k�^c��`�ͨDk^�`��
�.��\��0u���ƽ�#g�[����P=�L��s�Pmt��@�73�黽= ��a�k'q\0�0��1i��r�Q�ɫ��kej�����T�L��K�-��>a0��m����5��=4]XU6�6�+����9����q�0�B�xY;s�K%�U*��r4����[��n�3z|��k��;4ڬOQke^l�\0@�gd�tNE4J��1ݢ���~2��]vU��	�jJL�m�8�G����,~D�O˯�����SWL�,������QU�˔{o&>}�	�m��;����>^_m3�D���i�v 'Rbu������1�=�Y3St"�l�:�i�w;7��;=�a(%�^�G5�FT'w��tØ^�����G����uԳfډn�oY�yNe�v��jٶ7	Rcl���z-���5 v��1a��p�C������E��E�K1��H�jr����.���/��]g���U������z@�l[�;���t�xIC2p���i�ޥ.� ��=�ָx1e�^�D%���t��w$qb ��ˌ�0�ϝ�vrx���1r),�}��C�9��ү��7��/,���ǲv�����Z��R�iמ��=�r,Uנ�K鰡c�J<�rk�==W����sA��}<�Ir�gp,�#��:Q�͕�\ӭ^��0aj��UC��Y���]�7�Q����6a$���-�
�)N��A�ˉs4ւ�304�S�C��\��^��X�.	�-��W)F�JUzl��
�K�bR["�l6N�;lz��X����sT��@�&u�"ޱ���
�A"�������z቉6�_n���6U^a;�e	]�T���u��PcD᷽i6C���x�k3�.�o_|�`�S�f��a�}�P��b�,�z�����:.<xS͜������h��5#W/;;.b�[�3$�SntOu`ͦR���x�u�r�Ë;ЇXxM[����oW^lm�Go3S0����q<.�6cx)�M��4�J�<���7p�±��ђ񵭗����2I��a�ُ�[���>��mo?`����턵) ��:�FgvvT���*\m?t���eH<�,ǘ-�9�#ep��a��R�3��}��r�7��9U�'���n��� ���7��W!��|����1�蜧ueo�$����59�-�]�2�Wpo0�}<�[%k<e;��7�}��),�ˎ�g�6@�4�Β�u^�]հ_���G;1����ڽչ�[pП0#Y�e�r5���Q���źӰ�����JNi��˜�c�:Gp���#->�,�͈é_����DE��ͨ��O�s�k/���N��inS��\%�\2� �}	*הn�k�ʦ�m^�h�7N�n�B�pD�O��=���=9�����'�[�읓n`t��.ϋ��#�aNjy��w;�Ȓ���}B��p��`ښǃW�yHu_WNKn]��E�wah�յ/w8�H��H+�쒗qS�y�<���Ц^_Wl������{���x�wc�߹F����ƋiΘo�ě|�+5���70 ������7[}!�{����S�e^8�*�»�Vj�O�[{e Gm�]U�ǻgGq7���P���&.O��2�5�Wmy�ǯ3\*�R��Q�]��v�ӛQ/ש�Ad`�sGn#�+����8d�YG��27���?;U�1�o۴��fJ�u5m �("�HV�+Vȑ�RYs�*n��|���s8F��ݮ�<j�-H�Sّ ��H\�4�?t�R�l6}M֫����NS���z�*�ˤW4.<�]�t�rE�L	����e�K۽�s�����m���r�@e(�+��6�;<5��Vc�Y�A0���rI+���zmc�x�x�=�U+�E*F+�wI�u!C;u<�h�7	�[c�9��{:g�[�Xvåƣ��5F������q���F��u�0�[VfffwTL��ۭ7+��&A���	l�4��\�^�-Y��z���_�����}��/o�����x�/&�沧`�v]��!���^��7h����uo
�����(�����N�B3�HJ�^p{��S;Z��~�;��iX�ۗȊ6@Zz��Q�G��n.�s.ю����:����7݈�����"�`=z�1êL��Z��YW�u=Ud�ͦmx�7�3�����OM������g�].��ޒlr�'eY�4U���:�ԓ���׼����yVNvҤ���s0^� ���ѷW�{�;��S�V64l�}�zHn#}���# �ٽ|sD:A=uy\�j����Kr��N��;oj%k��,#�k�����ZI�M��%��8�+�ɠs��}w/�?h��!���s���6��A.���1��mB����hi��z�LoC�i�y��M��zh�޹�ѕy�xh�t��H��/UCľE���R��C��W]��f�a֓�1n^6�t����2��xX�K,�!�euCE^N�����.2��e�A�F��3GԻ��|��붭�bID�l��Wu��[��VW:��4����׋z�vԒ�`u�q'���,#pr��pA�n�V�:(�*-3���@)�6~�XvM=�G��h�ܫ%��-�S�p�Y��f�3(R��U�I�
U:e2���T�Ֆor�T���@�4�wH��,���nIIMQ�U�N7�g��~vp[�q{1hNf>7\%���ۂk�Ë5��v�R4l��)b�z�6�F#�X�	������N��YZp3�C�<ݛ�g\gn���Ĩ,=���+�k�L.n�s��[ۼ�*u����-�g�b�Q����Y�:�����5b�CL�س97�2�u�Bwf�P��=�/T]ȣs������>>�CC�����^�K9�.��n�*i��X*��D����OP�h*f+�k�p���wQ�M�B#%*/�H1v�����bc��vV(�>�Zct�Mb{f��q�;in�EH"�"*ڼDX��y%�s�R��<"gge�P��e��.��2#��p��k�ႫN�Z9�[�b��:�a-K/��{|�`W����-��+�Dl=�2 �e_-̷\]�vir0�N�J�bEu�ٯ&37���8�Z�N�s��bw�El2O��r�ͦY�!��J|��z!�p�2��}�,�vE뱜hT��ȉn�Ţ
�`�Y��^��L�_.��xΖ� �"�����+�N������w�Qk��fK_�>���;��梈�)�_8�. ���S3�Jf�p���ҳ�,RarB��@ǻ�R���ȓ��ރ[n��z__,Y�G�J+n{����݆ʀ��:�٢AZ�o8�\�� �s�Xw=_��7����f
���e:w6��I{���rwEq�({�I����� �6�p��ET��8��hI�����Z"}�������5m�`հ�WcE��Acv�\A�ōm���1h-�b�;f�֫T�#ZƳlZ�Z0SPl[V�c�OU�n��d��U��1�و�����3X�8��f-`֌��`�f��F���h����pu��Tl���4�e�M���m,A�Z3[M��4f����j�v�5�Umb����Zqhы���Dm��:qj+u��j�wgua�n�:s��X��S��66��؋���;F(�ūN��E�ۻ���b5�(�[���؝ݹ֝Zk��j�"����G�i��jF������c=�lZLk6#Q���Fխm;�6�"��㋢7X��g:6�����Xш�#v5\X�U@]k��v�:�.͍D֫T�|?�������8,�����S.�0͛�ھ��4M�![{����]&�*(�\�Y}�b�^������[3�1�6���k]����f7���=A�7ͣ��u@�gѬ�o��km]Q��Zl��Y�v:⏉h���l��&���[4�ƔUL�?Cϑ2"��z[��T������A0݂zƛs�������vSkb�wgns{4D3�#/;<���<�>��"t�$$�f�<�pR��Nc�c(rpma�w��w��Y�2��-��u����ؼDGY�p>=Ʌ �QJn.(�f��麮C"�ɖ{�%ow&�nz�s��84u@eL�1�3�F�ӽ�$������%��b
�9��%n%C&;e�Cb7�2���dvY��������)�]�^;�q.o�l�@�,�1��L4�k�Ғ�N�f�@���c��x]\JU��˽�u4��q9�ut�Uud[�80Ñ�\4G�yi�� ^W�<O�>��@g����-�:M�P��H�j�Q��DX�GN���������ZKpWc��9����>�J�u���BK�<!�9z1!��*��M��/�S�^��Q�-��P���'��Ħ��㒯7{�G����W��s���MQ��w^������c���ݧ�"��\bS����kx�"ȅ4SEt��J+Z:�61��m�TY��b{2`�NL��8!��Al��8j�h�z2uC٭�f@87*�ov_^��j��[d�q �l��ly�oLl��$�99�2�a�ֶT��w��D�9�.8��Mn�]���
`�e�\���_��i���������hl���ʒ�(���+��e�'���G3z�v������;����(,�}eo�[��2���{�t��d��-�F6�7>�5����\��hЌn���}�|�W���C�vH ���^}K5u�GM�E�����t����.ĎQ�1G���^��J����/,č$� �"wK�ÿ64l�Z�����|�)���1B�K#�(�v���A�h�Al�'q��kc�@v�	�%�*�Hا3����A(w&�����4n!L�����9ѓGk;�U�b���Gڽw�d�3����u묞�.��x���,�[�3��l^�y��Y9]݈v�kwtH& ���Ntz�V�9.~Y�@TJKwL}���1]��[P��d]�A��z\jP=wwC�cLEH�j������׫��4Q֑�J}sN��,�����G���IKC-��sM^�!�&�cgx���!Y�B�ْ�9�U��+�;9�`�hv�:p�����!c��]�Hg��@r�k�)�+
��٪}��Z�.h��d՞;���Asl��PE��9(�Eq�gG�<¤�VB,pQK|n񳲷%��q:a�l�k�:�@B�Hl�7��QLt�J#u��Y��mf.�ܳ���Q�zF���j�=�Cf>�p�=_���Tއ}=�-&L�ҷ2qZ�(��û�sVw�m+�V��|����;(�w���<�o��ȋKr*�&V_n�o?Lr�ri��<�Z`��]���P�l�!�{�!���^�ev�wn��K�wdr�NM��-�k��
S�Xa��ݍ��-�N��ӝQ��W�$���ziV�pQ�]y^��[�=^n�cu�uw{p�kI� e,�M�Y*��*�N�'}N�.�è�ε��|���Q������D���j�X����w�V(��HZMwh�1A��5)c1]+��J���R��=��3Q�uCz��c�(\8�׻՟aA᤬.�0$=pz�{1��qaf|�{�3��������hF���Ⱦ/VQ�����MS�6޾�5���^S�{|뽰�(����0���R�o7Z�K��鱩!qI��'H�yV�\��{�@:(��22�1 h����M�駙l�۲��:���W�Di:
VD��<K-sӜ�g�b-�u�&l�=�*�h�v����M]m�66{R��� ����Sj�#��,�f��Hy~�ٛ���G��z�ʡh�L\�.!m�A6��]����͎$��dԪ�/\M<a��ZFͿM&t:�X�n�(��{%w2
�rD����g]��ɭ��}�y��`�s'����3AA BB=[µlm�j��l����l�{�h�@�.�RR�X7/!��۲��[Br�5�!�m�!Շ�Q�Z{-��1��|�C�L��ϛ+EK�� F~ɝl�<���f+�+���Q���9]u����_{R�Uu�7��e�ä��N�ɩÙ��������KJ� �=�چ�hd�J����=�����2K7{��&L���"Z�k�ka
(�5Z�Ie��I�۶��q{��-�6�;�e�桏�'8A����a,�q�tg6�;=!�K��K'CY�������4��#��1��䪅��"�J`o�uI�te��dƲ�(��Ѿ�E�������%T�������\�-wy`�h�ؑ�p�_FJ����8�0q���a�+�3�g]�J��h��ڡ����Ov���#OV%t-����{��oR�����<��*]+�R�~�h�f�t�j��������O��5��U2��C�����N��M��vյ�+{�2D���$��]���Q��s-�Z�ݞ/$�$*J�*F�?��2��7@�bt�$$������N�ͺŻ�ݏ��p�S�bg�|�JDm]u���xH�ge!���s�k�ȁ��7��v߻e7l�E<��܂Z�r^�VE�Q\}��&]�����q�Bn_!�`��};Uϙn!��*/��Ϲ@���	ә�2�8�F���0�]�Q��� l΀����E�]�׬���R�����ަ��pL�ٹ`�=jΌi�[1�3L��`�Ó0eS�G$r�H��u�c�;�XyА:����+��)��~2+ڮ]�{J��d"��0���Ĳ���Ȥ�[݆7+��љ@���	��vUi�5l�� n�]��y�3�q����������T�{���#T.�8��:�w����]���l�p��`ý��.nC`C���Eo�)+����6�jA
�u���3���7�����8�LQܝ�	����l�%r��s�M�ѻV��1m��:[*�2d�і6�aH!!�,���:�ƻ߯(���	*n5D���dee-��Qn�eζ���~�U�'�1�̩��݉~N�G�����i���t7�0އx�L�7=�sv�c�(��ܮ�{�k��5�&����D�P���r+->׫�Cs4��������f�egb��|�
==�pn��~
�c�둜�1�dX�����_�ƺ��3s��R8��7�>��Z5k'u��%X��yFm��� �ok��>6?̉쫺�S=�1�v���a]����̽ �6ð[���7�Z���S�<�4%`Qg#qU�ڙ�y1���7��a>�tsuN5�U����by+�Ն1��%��OA�SnD�U`��?�-�?Z��&����=^c�x�����|��8��{f��Z�-��C]��=��²�}ĺ�����$���+X�m����I�n����~�)�~��A������G^Q��/�ٲ��K7���vw`�,��
�$"^*�Hا3��,t �5R9�cZ��5;F�a���o9��ZƑ�u�eg��l4�=���a���K̟���1��V��Y�T�1����H%O���@�d�0����YE^�����n{x�Ӗ
ߴh:��"�n�r��J��~�m܊�k8	ܹ5�<y[��g �g�r*a�Uz'�'���:J��v	ư]�Ot���[�z`v��QU@>�uә��@"�H@��8����]��M�3���o��#��9�Z��	��a�َ����d9�Ѽ8�?��� �AVv&�[98�3��������[P����[�x��׺���a�ot*�W}�3��f�>{K|��
�Zf��GZ���f�	w�"�s��.���%:0�۔j����250�^A��n3�h���_,��W��N�7�1�[&p˂+MK�Vn�&�����)(�+M�5�@Y*}��-�[������gY���e�v����jOP���X6�F(����0������ųz�_>�m�ú�:hG*5�&괥"��EIPHd_8����\44R�[;=�6�<A�E�#�;�E�^rWS-Y\���T��ȴ��y���{gN� �n�w���H~�hF�پ;"�=n&n2�;��nuM^��v��������o{=�e�Pc�hg9���E�$�Lu���m����5�*���5Ǜ-��9 ���Ox��F=����1/���ycbc"����-̨�=�x��ȉ������nM��~Л��Z��;�]����oA15�쉫��d�@�8��U�W�������R�7��u(~t��Au�����{%�%��A�mI�G�Z�v��f�f3���5���������|Nhm��!ׇ�xz.��{��g���3�y�j�5�z���{�9�;�-���Ǜ����'/xKO4AT�e�*�+��Z�M��i�q��os�5^��۳n�jw�ڕh��v�����e�Pة��c�c��z���T
�~�L�qb;����-��H�,T�T�[լz��X�{G�j4�̝�L�W~5�#���!� _�A"[�����N�pn��ͻ�z6�뮝.�4
JC�ÍW��N庑ّ!c$,63���
!��Yzk/��G
&����c�J\E�hT�0����P�XQݝ7�5�`��L�4���*�e4
2�j�������ͧ��>N±\���݈�V�!�?�Nyà�}M���JM��4���!�;-�Ckܳt�䞛���H�!��x����Td��N=u[˔�Ŵ�kV;�8sZ_V�v��AJ7;�Lq��o�.��^�4��y�rՌ��W�tv�oQsr��r��=M��G4�1l���y���p�s�wFq˽m���#L�n�E��l��٣a��i�y�S[3��H;*��7�[vI+/��2���Н��P��$��m���a�Y9~�{��ε��x�7�*�g�Y���ʙ�p��Z�3ϼ�*82�{+��<e�S��]��ŷ�
�&�w=}����8��Y˞Γ(^���y��z� ��pDJ�5"��q6��w*��_�\�/ V�48�ź���t��}����[܂x��n˃y��ݽP��c�#�I�����1>�HI!�t�m&�QN9���6{����"���H��s�B�RWQuћ���DO���{���<�3����[����v<��� ~��&�2R��hD�N,y�;��Gd��lj���!��vo-�$r�2�cM婹�3��T�F����S�r�t4��5y�=չ�ِ�iI,R�л$���sV��tE��W�YV)`Q������n���"o�H�AN�U�%*�S?������[�K˅m;t����q�!erC$�%VB�`�)+�xGv��*xr��+^�ѿ�l�Տ����{�H{�^� 9Kcx-B���t���"���rrL>���û�3$q�;=��a�N��Ɍ����B�l�������y{}��g�����}>���||�b9Z,+2g����>��+|�W��ȼ�����a��}�7�(6#ǉz`��5Y���0za+����6��4s������*N����/_-Ue��+���6p�a�d�7Q;9��\�ܓL�TH��d�/i6#`�Q�1i� 0WIG.��V9���T@{/��/=�ou_,��t�]\���v�I��3�W�X+{Q�s��`�[f9B��%�S<����J�r���̋�ڱ�:L����Fh�gSP��5�g�FU���ř���bӷ���zM˸v}�]\�A)s�����<�L��(�E3J�K�P���f�'{ڢ<�QI��r��U�L��+r�b���#����vX�ޫ%�Y��7%� E��Qn�1+�ۋ[��3���ХgN�.��"��RBe�j���K��%�����˾����V���p��7K]�_�Á�N�@����!����p���촋K���Tz�Cz��YVٗ��ygd�KI�k�(�|��|�7U�D��Xi_(�'�wk;��#��=Jk=_�N/�+�c̵%t!�W}鶙������!2K`!�U�y��u�o�;
O�U~���[G��5�Ɨw�F�yO��_&u>���0�#�y)[av���tt��g�����
��L[�哦���|=��~SؽI�U���ՁAl�x�+���ŕ�3�b�w7u�<ԥ�gm]�J�U�ٓ7����e���S�[�kDs�f5ܳ��W�hf(�������t���:)̊�ޝ��̻���Hײ���[�}����M!�1�a�.	��S����k	7�:��s!��c"h�w�_rr�ov�J���h�뫼�C���;UC�(��F\�B�qn�!�p�%�"WI��Ɂ�����=�T鏦���D;xd�ht;��$�w�"��@�a�Zaot]����6�#tNΧyä3S��9y|W%�	����n��zo���fJ��-��ƀ�W������-1������Тm�I���:�c�H(�[�(�h��1w7��+I��i�%�S�Z�y���_'3��#�)Y�"L���\�s��pm>��z�p��0jB�������2$��op˹�9�5تR��}�W3,Uᒷ+���c��Eۺ�5E����;#�S�{�p\p,,ɸࣸ�X�8�u�u�%�nd��yĬ����&A�םa���s$�峴�Ґ�å�m\�}tl�3���w��nr��� �G%cZyO��3ў�^��2��q'�c'[{E�9�0��W5�6w�إ��[j?���7�/Bx�9]���T�x'��~��(�Μܗ7DH�YK9��m��s��Se��3`�������Ր��@H����W��ճ�/��I�b3�)�4q��]?(ⴴ������w٢t�T@���>�9X]�.�Kn)w����:Y#3�2u��h����~URbIc��>~~5�y]߯�EU{Gtd�6�������F�i��h��[�[��椴h���4m��qv�clj5�kcu�����ص�v����v;��؊cEۛc����(�ڣ����c��F���Ѧ�Z���,h���S\Cwu�c8��j�V�hưTQLQݹ��tQ���j.ƫX�F�1��;`��2lF���ۻ&�m�mh��Zڮ狎�IۻA[��b���F�������I�1lmb��b�:���f-������b�7gvm�5[)��A��u�F�Z��j�LMU���mM)U[��ZcK�ы[F���ت���S�E�#UFe�kc;c��N�kQ[Nڴ[LE�hΝ�b�f�lm��,�#m5Mb�[8�m�-;8���d�lꭜk�ƪj6�UDX��%4�5���T��6�V�%��U1ŧh�i4cYъ�����+�ӌ(�C�Ig��>Nq�v"�Ǒ4E������έP�C��c$��!oFlٷG�n3+�-���u݋;8X8�XS&�E�s7n +v�'a��H�|�
B���kyX��E�{����a}���>׷(2�ܡs�����/��ws!3��y$^ig?��H�?c:��7m��rX��{7�VI���#����J����&��(ˉ�I�F��M=rar]�;j�g_p�D8:�5�/zN�+d7a�ҧ(T�M�3@B�7\ۧ���&���ƥ^�>Ɣ·3��c϶f1�H�/�|��e݁�j!+���'8��[�Xu�l��/�Pm�ww@��f��P�����q>��?b��5������ԥ�v���=-z~��A�
��z:�-O���J���c<wvϫr�wr��Y0D�xUґ�Ng%�t� �A�g3�m����Y�P3+p��=C��;^G Bz���h�iͥ7L�e��>��\$���onw���t.Z7�=��XUd���j�8AR��U��(�a��!7�F�h����Cl�d��9}�>��S�r�,��pηwBɸT:�.�ѷ��)�w�	�y��t]����vMlZ�:۸Mt���º��s�Q��]�;���6܌�M��!�*�TW����C=Fk���������n^��(&=ν��W*�o�a��9����2U�;��T�7]�B<R��*��)����}��3�y=�F{~�������r*D:*�z8@�GY"5^;i
]�Y75�g$^��Y�w
���?߿m>��ӪӞ�FG�!�)�U_��Ҝz��[�M��M�1�y���xƼ�:��=�Cf<{E�[��un5$��'���;Y���H�Z�%�M�\���pQg���2�����?vS��b����0^�)����ꞡ|�}\��F(��]�>�:4�X+�n�UDi����d�Bז�B���G4�,��R�ޗ��Yh-iŢ+b�;�_��t�@��}>Cz|��;�oM*J�e�6��+:n�g#�l�X�v��;Cgè7w�Ԃ�~�w�����X�d��������]�'[U@��	��k�A�;H�������E�11\�r&�3��a��"-J��`�g��Ūor�Je�Μ�HQ+L�o��t��W�M^0���v{�r���4{�:��Y��f��;�(jl]u��쫫i����C���������H�����čË�&r���7��|�y<KR��^�-�t��NC;����{�-W�����Y���b�����7�N�ǜ���FC8@��h���&!�z'wi�g�4��^���>��"Gq�!" ���-WE�=�NS���[;�p�_p�H؁�-6aZ"j���ZP4q,�8�(�P2Ӷ�Gs�Ú��:n��+�.���A(�z���M����~��E��+z��x_�l�=�mB�p�m�5׸�uSÚ��+�a߄ye�^�]����(n^��`��p�l�{�|.��zA�&�U@�d��x��:�A"q9N�������u��m�}�%�J�xD��9�Tݭ�u��B��Q��Ɣ�y�2��doV���	A�f����t�J��+�
[�͕��Nmŗh	�����շ�_7��h�����7�U��FR��5�r����;j:�"ŵlw���+g2��M���@qN�����ٖ�urRG���)R/����_33a��]S(�w���e��j��c2��e��8Re��v�Ȯ�O?0m�3o�t:U���s�7�6�V��qף�u�)6=�v�N���z��p�=�"���U E�����g%��Hо��|���v�3�o�M�r�#p{�R���0h�=�f;f^��MQ<]'aC��<�t�]oDl�@A� Y�#��Q1O�q�a���݉{�F!n��Lq�����]�3�t��T�
y�si�{7=�y��� �8�J>��!m
�n�f7�<�+�76��*��Vv��;>�*R4.���/7�G=�'���ҡ&��w�ڽ�ݽ:8[�Ty��P�c�/+W1��-�>&;��1;-�+5���e�����¦��C��YgT_*����j�yf'I"BI&���WEWm��?`֗CtTx������,���Ǥ����9��4^��:�nӯ�f�{V���ɦ򔎊}v�݈%���1�N����.4f��}�Vwr��o.����ve.Ɩ��W4�F�8B�"�A5�<�t�{5B���6�5w_�W����)���!eiI,P�m�ʢ*i�մ�}s���𪺟A���_���m�)�x�Z�ɏ8w#�֑��c�㔭Ѹ�����[Z�9�d��5�-�2���xw���:ǵ{�t���O�I��y��m
/��^m@{��$��4\�^�	wD��m&�e��Ytg�٭Q/�e��C��m���l0l��Sz���v _#<�)���I�R�T�=����DLf���ܨm u3�
���#��\��3�RV�8���kn�"+1�'��fN����*�e����*�v����P(���$�R��k�e��z�"���_n�N��C
 ��8-�׵�uɆ��7�<U8Kv�v���y�ͼy�4u_�&u�u~�]�����hJv�����-~�=��������%C��ʽ}����i��V+�19�\�����s7n�O�z'Ja���<�:�GJY��j!Y�#)>�E<B����Ψo0#����5�'׽F���݆����Ҍ�I��hf����W�M��1�Gl�c,�^�پa�z���/��&��;<��c��n\��ttY��gq�·vE�Y��K5��c6�}�j7��ɍǗ+VT_ ^5�;��u��F�g����R�:�~��V���,��2��>��C��l��Q�Aft�5��|�A2ȭ8q��Un����F�����.ȉC�vкꚳ��x�:�N��{��Ͷ8t�g�0�[Z��8��'��o�;�!�ւ�׏lG`�[�9�AЮnI3N���m�",��չ׽K�K����\������S��SǬ/�y���O1�.&��������E��U�*���ܐ�u��8�5⎶����t����MXW�"���x0ூ�{��5�VLn�7ܐS�q�N�h�{p��CD�ֺ�uݷf�gO�i�h0�K�W"�[��t
�R�1�0�)N�T]^���wdOF�*�U��Mn�
b*�:*�p�_#�u��2[��,���6����k���S�}��R6|`H"`:A���З��3�2�]y��E�EaƄ�%̸�w�ruu {�p4Vy.1��Y0�敬�;ݒ3H�/�\ZrJ+�9:�i�~L(���dݞ�f�//x��b�b
�'�GT��>�W<��b��c��KL!�ҹ�qwy�ޟ'6��:��+&l�g�{]:�<>�9�P$Nw=<DlD�8>|]%-�6e,��:����zL�m��F&vu�,w�����xr�p�����]��/�j�h���4�8�l��%t���V!����	�KU���%?�N�M��?��{�:~1����4iɺ�)M-ށW�����g_��&�d�ޞ��H�,(g�!� !��F}�7��%w�$4�yn�~���GgomwM��Bt���Ns8f�'�7�]؍�[R��s��_�D� ��>~]��S�_��3�����M;fGw�9��8Лn��5�Z�df6�.���%�H�Z��x�s!�\_V��>�m28���FGS�CNYUA�]��ĉ5�w�z��({\y�L����=ydD�'��D׎Yi!���s2O:�ٽ�2�h7bdR�=�5WUxvV�@�VD3��L"��{-m��v�>힒��������w��(���������9"����{Sݽp4��&�Ok��FA]X�a���������q4fm鍹� c���rM�6 ����駏M3����,��۵Qr������]6�&s��ۺ��w���js��^��%`�n�%��lyI�[�}]��C-��ͧ6m.|>���5�%�$�F8;S�O��ǻk9r�"���D�k���R�5r_[������U�z�[�X!(u���Ç_,�Uv���ξ˾�۳��V^���<j�ݩ��{0����iQ"5\��Zxqӛ�3�
Di7�WЉ�t��\�w�a�k��4��[	�ݹ8x���ht�\ F@t�}G_[e4Q��ڥq�tq:~�c�X�Bp�˾̖�;d�a�K���t��f�OP�U�΢U��
>�����y��8�c����B����cj�Ǎp�.�=�����n���jd��l���@U��+vU��S��#z<�_�
�����3%Y��\Pմ�Ε��{Ǻ��WBٟ6��n�Nk:�67���W��!Ӎ0�n�B��H�ˢm�\�{ϸ;��w.�w=�`h�Z.�.70��i���E��C��|n[x��q�2D��u���;��������͹�\q[��g����y�Q���w���,��$?����U_KY3�p�ճX~�g�[�k>�rG�hv,��۠��:����;��~:�G����$�����X��̼\��2Vg(�@���(��S���D������,��p7k(�(�Ĩp��|B�VF���^��Y�\0��y<��������]n���jv�V�@6����Ʌ��^_��p��B�RV#_�L.��Ͷ�������n�v��݂�vx��ܚ�V{���8�܂W结�Lݲ�Tv��_��wu����޳��$���:�����cH��>��3���
n�׭3YO}�z��u$ynwPɈ�,���fMA�-��*j ��Т�_�t^f]�3��ȃeB���Wa|�C� �T.�R�?���f�����:Z�s�e�WD��n�j���<�")�@�di��W�~�������)ޛmȷ}=<�Ϸ��ԍ`����[>��Y
(�rj���`����Kw��Z�g�w��\�ifwmt�m�HAn$Fj�����g�ͯ�ݨ��]i�r��ƸW�=3��z��Ӭ����Ϗ��۴�*���r��ϱ�C��t{N���8�G��O�0�f��Wt?<eۧ�r�q��.����Iꋉ�W�u�p�&�*X՛�h��a�߳��2����(�oh^�U��	E��2��k�1���xs�W8x��#���!3o��
�"�}�r�t�k��m^�8�k���9f3���z�5q)����ȏ�.����e�þ�8\f6t�t��GJY�(���e���q�2)�sf5�{g�r�>/W��a����{ҷ�V��n���4-J�-VYnw�]��x�5��Sh搂0l���}�nr&.�q�'�z�f��3��L��snHF:N�=!�]����<+5�?^C6��ܨ����z��ל��n$��,Ok��8����t+�5�f�շ��:���s�!�m�U�>����	���{�rZ������UH��|������}���Tv�T���y!>�C��m�6�g�~��?ޮ�p�&�E���Ǘ+�q����7�o�� �+��f���['d�V�b*&�������A���
f`U#�}��X.��@����2'��^����̌��h��UΫu"��@.���tU���{�ޏW�������{=��g������~0DE��k��ۤFq�%�*�ԥy�Ѽvn�ݳཬ�xp�N�cq�{������W�iW�%�w3�:L�Ϝ���6+5���u� �J�{�<�~�V
�OgA���w��	��q�����V[�/�<97�v��|�'�ɷ�e�o	���R�K4w[���,�+����ٳ�:B����6�X��"d!B�>�6ܢ��UL�@9�x��=�z�툹��튁Ȱ��⫚a9s*��Ϲ�u�;��ɝ�Qvrg1�C�[�.ϝ�S c�d�7uo�ղ�R��ێ%���Ìi�����kᾙRjA)�^�4Y� O�е�{0��Oޭ��R����?|}����/B|e@����Nnz�0��0�o��>��w��ӓ��6_�z����d��|�������>|�1vY�d���k��sI��pGduvrҸl����y��i\X��Znqs�m�@^v�^�}�i����́�&'L��:��λ�K�c��0������v���s�'�{���Уߋg/f�����w��B��r��#���T�{����_�!�a,܃u��wF5P��uGݨiI�
�<�v��`"�l�%��V�̺��et[���m#o���J����4Úַo"_.���ݱL�t::o�J�ҹIғ����Sd)�������w�+�_w6�V�;Ϫ����{s�j�<�QZ������L,��O�F�yyI^=뼜�Ph�`�(u^�#�-7�Ƈ)l���5�C�����2]w/!��ۄ3�7�����E(u�;穡�ߏ���!V�[����3_P�%𲢺*��n��s��ōm����o#]�lN���;J�U�s6��0-��[��͓�m�x�a���.wRK�Ȟ��Y���ˤ�x�ݡ��&[���j�}��iԹ���x���78�c63O62�vW��.�&ݓA��p具B�9�z����Jj)ׄ���_x��[g�\���# +T�>�C�s��p�xx��	�z�g�3<���J�=�=+��;�;.�荦��ka��3��!^%��^���<���w�.��i�/+�\U�.�8�qf����IeX�T9��8�՛н�ܡ%����ޮ��=�!<�b���"Ń~�戞(2�d�"�	U;���9ؽ�ɘ�P9b=�:�:����:���1�o����>+�;e֤�e	���F�%nh���s"��Sh��\λn�.+i�M��XM��\��)�T�XWƜ�˛���R��zD�	�XЗ���w��Y2�[���]��h}Ş����v�|t������K��¸��%w�,�yLm�0	@;�}uJ$(�6C�S{��M�^"��{�"���������tkl\�]���﨏����Ɲ�]Ξ�m�^��z�	z�:�J�����c�>:��� �=��jڠ(�j(��R�Ռ��D�Z*"z:�N�ŃV�ƬE�N�q�l[Dk�jf5��ѧ�a�ت��x��[V���͍h6��]�D�[b���j��1;h�ccl[TN�6�m���j1Q�[�$��rH�#m����rH�P�%͢��[4X��Ί'X���j	�3[5�ڶ*"��1��n-[Kn㋶5��m�Dc:ر��1����T�Eu����EF���#`��1Tl[1���ꦫc!��h�m��(��;;j�MAM�Ƶ�n����Y4lV�Ѧ�F%*ڶ��[n���Z�M�Q�g[qݸݩ��5cj��GZ�g$M[l�b�ݞ.64�qF
h6��AE:�l[T�����F��I�ʊ�&�����D�i�N����֭�GF�5Q`δ�m`�1ј��Q��ƱTS6�RUuݪH��kk&أm[5�����AE�lb�Q%--lV"ѭ&'O��������p����\���[�nj/�9Cݎ�v}����t��ZݙY{oO��\����f�ܕ�Zk��{*�I�ھφ�gP/���R*x>��u>� �d�����p޵����h��`��!I�2��\N����\zζcƋ��������o&�-��
o>dF��}C�8O"9%�r '���|�j[�&!r.�2�2�zw�[=k�r����<�1��8W-yR1^+���hꓶ�T�˳�Q����y;X�f�`z�2#gS�rn��R��*f���L09<�kvz�b��*=�#$m0|���7�3���>��h�3Kt�U���k����X�f�y.��N���Pn��a�`B��FFo_K�.�ne^��ʽm�0�H�OPc��ܛ�A1��zC���=x�+�Y5�����uW~�?!ߤY͵դ1�}��g�<��K͈�b,�Q����zף�.W���_����;�z�ȍ'��A�|��"���[7/-�B�ɶh��B��a�����e���c���َ]`����4*��@b��`�<�"��b����k�����qQMJ����0zr���E�cv�٪$_�w�������n�v5�q\|_�u��k����m^Rs���:mU�����#<+��Ѩ���ò� h�Z
ZԢ%�d��8�w77��A��q�o(�+}��{��꧟;ѭΩ�oᶺ��k�<����LTK�2FPt�֟��D���
}sbL;�ݜs��Lt�^�S�_,y�{����N���$g�̗:�|w3�^�����\-������N�o\������t��1(�)t�<j�ݩ��:;�!Z6XtD�u�Ӑo����;��jE�"=D�t)�/�t��sɔ�����j�rc��^D�y��N�,r�t�@�#�_Ue5��>�K�ĵ�4D�xI����Xwfa�6:�"��B��a��_�����9\٩��a2��3��EX6��d-��ɞ�#M�Ot��R;7����l�Ϙ,��[ϰS6L�Zl��.�S�׬ތ�����޺�I�^��b�n�W{#����a��a�7��/�2��U��Cw�P��z�ޫ�C�c��R��4�[�A�CQ(Cy�Εg�w�M�S�b����v�{vo�&$o<2����{�8 ��PbL�='���Z�%�o� �$�A����:�}ɻ�G����2-9	����v�t�(N�GId΁d��|m-��QH��dRVv+��s�Z��Ǻ��W@[#f��~�Ncx`�3	�x�S��֩�-kn���\aJ�m�Vrz�q��4y$�����T��Q�\t��ۀ� ��g
�����Jo"�q�2G�ʄn*�s["9I����{d��+dng��,Ǟ�e�6�y�E���`έ�nlN^�fn���_��h�T<��ט��d�YjJ�W\׼�ŧ�K'���w(�����l�ܛ@���w��
�	X)��dn>h��&q�v���11��Vw��#�Y�U�5z���ә��;�Ҍc���Ns���n֍#FlQ�B�*�bq
=��)ba~[ԝ�-��{.�rCc����;z��!��A���!!�E���:
F�]ĥ��3ɬWbn{)\�n��}��Lf��+�$FL:S\��e$��WHs�Y?=LGEt�+�.���t�����4�-L�=�~'4�w?9��A�Q��Wv�a^F���`�8��ơE6�5ew'��ٗ�9ɺ3����y\U�ʭ��U�8}ԗm[�b��L,�}&�K2����_x�8l�Z"���?%�?X)d�c�b4���S��t�{�������T7} ��:��'H6B�ȕ.tFj=�;ټ�6o��c�M�w��@>:���@x}��@e���M���f�s1\���(�y�GU�Q25���:���f��7��+�����ov�����0㶆�.��h��B�sϸ�ɵ�i�h��ث��֪U�⎨�>"��i�:�:T���KiKhME	Y����q�.�^F��\X���!y�����ܑ{Ԩ9[>n�wp��S�jfs;l��n��4�kW)t;C�6��g���A��1�^���ܞ��f�d-��,T�M׾&8裝A�]�!� hF�ymny���Qϴ�:��&����Y��I#x�����(����3�S�P�nx�<���y���x�9� ��ϵ^�Y�YHD�$�%�J%�U�0R6e�|>������
���	3=w�z��/|�DWުW��߻��F?��ƹ����nc�o��on�6"��v���oš#�J�۳G���-�ɜ���4t^��?/�ˢ�`kسZ�5%1n*��ƌ��i-�z�i�y.����̤�{0f��\-���QH��;!�"8U��~�Wg>/p	G	�C�q�h��ZT@�P*n\��/�ӕ\}�� �8��,$�pT�W��B��W���X�Ù�b�"�<~�b��y�~�#�R
�P�����Sp�#U���z��ճ7�����)\R��OL���V�E[@2�S�ж���v���J9�m��o���hx=C��^H�m��Z\X-f�`���yם�־+_��j�*K��i���u�Z;<N���g͘�_'�Yg73k�|�����9�ϼ;�)�M�IEr���}����p�^s%���v�퓳�=�)xf2��.���]�:���L�-yR1!�m��..���z��/������^ .���Z��t\dFΪ��zrn�kX�ȗ��t5͉����2T*��6�>y�͂7��
/ݓ��W9����jD�
ݷ~�k���Q�W'iV�����1�](.gE����ǜ%�Ek�Ѭ�W�j����M8�=�nI��� C��U�P��~�}!���UD���V5����\.���*��@�-ug�������D!��A9#aP��;�{�sy>�ʙj�]��%��v�����a�!tm[o��C���l�û��겶}e��eP�݄�g�ٞ��=�݀�Slmete\��oOxSX���G����7��1�u��O1�%O�*�k�C;�׻[��َ�D��B��S�Z63k�C�O	Wݼ�׺��P��l�_m�v˞]e=9�`�(��9WT/�ԁՁ�nƻ�Ų���x6��\����"�L�]>��pXJ�N��H��/���z�,�8��F�E�N6NM�:
�i �@�p��ň;RY��Vח����I�T2OH�!g$xٓ^���̞�xU��w>�K;���~���R��1� V��+V��x�#E$ǌ�v��R�*���]��[����H�@z����0���
FpB����<�%`s��g�20��u�2�����P�d����a8�K��>����'}�1�r,.��<:��އ}��e�ս��k���씩��,�'c����D�pM�POm�շIh����y�wOuFT��'���C�EW-����#޵)�l�WUD�QIrW�(f�n���sJlB�g�T�Fc����s���ʫ)��[E�e=0��"p�=�q�zu��ͧ#x0�a.d��?#Fc��U��7���q[��7���ȡ�y�#^+�|w�J�������{[o�b�AVo[���έݝ� Ѳjw��-w�[���GPn0pF�M�U�)ƛ����W�s	���^Β#P�9R��\�Ք8�R�]dl����5ou����=���= hLB4�&��Vw)o��e{�.}���Z贴�p����ֺθU�+�J�������M�d
���c�n�tMU����/v7.{����;t긂���E����S�����=����zS����8�&�p�wRd�8�%s�hk���tG�� =$�w���y��M��[�{�N+�"'�gd#dH=ɤ
�k��@�����>7�~t{c�\$����N��ݐ�(͒S6 pL]���u����N���ݳC�N�*�I�F���d�{�2,�[��!���kK�m���pG6'	�5�Ҍ���z)�\�m�8$�]Ь����n�n��![ت�;���G'V���l���z6.{y.�AHWfB]�7��%���%>�ͭ��=��O��8I�J�Lg�7�T�J�]���4U.��9�����:riԊ�t�Y'(BB �����9�S�A���v�����o_s��R������i�M3��H��C�5���L!�v^~�{�޹"|�"��}1��*�o�˫���P��>��E��`�
�+{{룷��u�2J�T�惢����[m� �j�l٭����ve���Cx�
�X�MYMEk铉L�/�?{F/]�'��⥝�>�]�q&DҊ:E0&<�sc��=ݜ��� <��ywd��uЁ���T�7^uV����-����:T��ZR�(��M�L=�k`�a��<L�9;��v�?��P}������ܟ^�*V�H�z���z`�D-����f������7�wiF���4q�kTV�}-�q�ƫ��#8\T&M��w�˞3և��^Kq�����G�7g��޲(L�_e�7ڍ;}h5ꀬ����-�v5�uuM��f�Z�����\�H���;#��U��!�[}u,ɵ|&�2t���;�A�<�\������dm)�&8�!�7���9�E���X&�p-���>���������9ʼˤ��ݒ	�����q�·t�������}��ǋ�m���OH���(�'�=����b�����ڋJu�s��t�'�;��P螨��W�⮈��<��%��t�)�3�s�G�'hk�9���޺T��C�&[��������:x�/�$C�qT#j�'⼨���@����g����c�w&��J�ɍ����aL�f0ֽ�I[�H����Gn�%��QB:�]���2����������u�}�%(�	JQ�ӡm�e:ʶx���qqr�m<�ڕs��/	�=�y���ѯ�H׋�r��h$U6��ӭ,b��,��֍���>���1���6kB7Űi���s�5�y���=�g�%���FݖU`W�O��q��0J�&�a��u�W��{L��S�h�*č-8�[�&sn�+41�ƍ�s%$�+4ijA�ɴ���{�j�h
7�R�U�ju��xu����3.go ��8T�aI�Z�\2�js�%c�(�P�5�Qՙ�]�,]苇Al�F���rl�(�+�l�E�&b�F�@�n��/�f�^Ol�����F��]@;�*��冷�Q�޵�A��&�k���Rv�T!�q�|�v6��!�`����T#��D$'�ʫ[[Fzw0��qӽGw���P2��`�<Fl��pQ���y�z���;Y�y;�2�z�狒�-Wɽ�g�߼�=�j�T��=�E��0vlqGR��C�[@F�l�_�(�sԬ��O�v̎�����.����k����Cv�g9�����9%+�n�7�_DӞ�����=�A��;�����9E�t��r`�gI�i���ȉO��jT�}����^�m�ٳ� ���
�T:-́���(���0"j���y94��	`l��Ͱ��F��|$�[+klky��fF�X�Z�el�����i}�!sIUQ]� �*/�?���_�)QE�O�8�,3�v�C�0,�ʳ�0,ʳ"̣+0,ʳ"�0�ȳ (�00,ʳ(̀L2�ȳ�"�+00,��̋0�ȳ*�0,��� L0,�3
�0�0,���*̋0�2,��*̫�0���29�f�Fd�fW�a�fA�Fd�fA�a�a�f�`Y�fA�dY�f�A�Fd�fA�Fe�fP~s��2� /� fUVvUW0��   L�0�Ƞ*�O�a@	�P& �B`	� & �` 	� ;=�<�@	� & � d@	�U� dUfUVm*���( L*�ʪ�*�� *�0�ʪ� 2���g�U� eUfVeUf  �eQ�`Y�eY�fE�VeY�fE�e�{=< L2���� L0,��Μ00,ʳ̋0,�3 �c����A�����TI�P) �h��U�����������۵�������~����D��|�������I$���<C���� *���
������?���d���K��������UTW�����?��?5{!�7�=(�;���3�wpz���v aP�A� � %Ud` 	eUd @	VVA� !V% X@XUY�U�@!Ue�U� �UZP �UX��H��DO8�A��?��S�J�*-(�P�P�P ߨ��������������G�������烥[�g�d[<n�A�
:�a3�TX�AUTW������}y���J ��
���������~�*���|�� *����������>G��>�A��o��'�<|O��8 �UU�d>||:ĒI!%�0�������#�[=�P?@������UTW�������UTW�����C��2���)�������������|���_A'���UE~����)�?�x������?�����O+� �"��>0`�~<PEu�����_��)���PVI��SV �V` �������N�����A#�Z��61HT+`Rl���R�MJ3kZJ�T2H�i�����U�)U�Be��]�ѣBƉi�I*�Zj�Qj0���e��F֙fj�CY�+cl�Y�����(F6;u�Y���6R��ƶձ��e
[Mm1�2V�b���IӜR�<�֭�٭LZ�ggm���ej�m�Em*��mYmV�Kf��M6�ZJ�ji��ٍTͤUml����jR�֕�1�f��-��d���UUٶ��F��  �/�o��r�w[ݭ�t�Jt:쌮�[j6�r�V�Z6���OWmvg��zƃ��շ{��N��4:e���Z҅�޻��wt��/o{���@��T�oZ�m�6�[a����\ͅ�  �G�
2$HhP������B�
B�!��.C�hP�CCB���_|=
(P�o_cپ[��=9�[ڽWn�Tu��N�ݵ4l�η:i��^�]��:��I��J��7�]o=Vֳ�{�卭J���k�  ����t�k��ޞv�ݍ�.I���&��lm�p^�]]�4:u@6�Z������Mzp�(6Ǧ����m^�`t��i5�5���z���a�7w�5��m���L٘�Y��  ����[���{�m�Wn��)C��m��n��R��;�ƞ�ҝfʹ�T�җ�wi�����4��q��v�Tְk�)�ũKMmWw.���զس-� Ǌ
�O{8�]m�B�>���(�t�IP�� 5��Μ���k½�@mv�4
���smC�+;���
�UF�fV�2�M� q�$����g��U/q�QB�9;�:�s��$����F뎠4ѵsp:�
���*�j��D����[5SVն�Y���fm12� w� �k_sm� �ܝ�R�]W8::m��w���Ps\�l��ۅQ!� �t�h �w�  �o{X����i�Ƭ�l5T�� ����tfV>��
=s� z<�@Vq�@�ѽ,� r��� �� �n�����zv����on3m6�-66Ŷ�ц��,�� ��  �o�� = ;ާ  (U�p@ݭp    ��� �[�@zs��  �Y��  ��g�sQ���lش���Ś��  s�M} �`4 z0  +k� � =������p 

��  ��` =�W=� ��={�  �)���R4#MhE=�	)IQ��i����2��ډ�@# a�JR�  ��J��4@��&eT� l�??�����b��Ƅ�w���P��cW�}���Ãj]R�J�U�,�_���x{�73���� �AP_��*��EA�z
�+��*��"��~�?~���,���R�io�7�p��[��+K۔���� LЋ��8��5ٺ��Yi��,���|	%-6o2İ�j��uD��
��a;�BHٔ� ��ʈ����iݭ�5H���*R@'��26[y�6�b�I�����Z�ҫ)�Nڶ+a��!�I�
IE�1)fJ#,0�MeՓymE>�3M���^M�,��,:�V�׏$�20�N'���Me:;�
t&7�p	2��JӮ�J#M+U"ô��U��`PC@��*�2�V�Jd�zl�U2h��C%� �Q��\�1�<��V, p*B�[R���,e�X��Ɗ��Z�Ҿm�DQ��\��-�����"H4�w>�	O��`\��ge�<�mL��Jb]���b��t,�J�ڭ�drY������ͨ/c��˵��\ ]��la,�N�N;�b�8�`o�ü7��O�w��	�%����k�Z��s�C}��%�=��E�#2u��iF�2Mw��4�˺�/Fj�%���
�?%�>�f�I��E��!��c7hI��52lJ�V��kc�j�K���t;4T�e�����M``V'Whe\���ɪӀ��ٵ�3a0$�BhɅo�+ ��iV���dM���u�\"����"l���J�M)��hXp��Oֳc�4�̣*�v�J�,��X54�誻�"��jlc�V����n��X���Ј�$?�e��1�U3t���6v��gu�6�ȍJm��f&ˡu�X���w#2j�FKW���j�äkhcֶ�zNU������v�O(e;&�߬elְ�*���ʹkww�e,�h
�0����+
���>��rV=U�������T$A��Y�A	�I�	3���^��\&nN����ԗYu�Kv�l��H2��*���H�f�����t�il�B$b�P��V.������3���8��4�oU�v��(E����ѣ�B������m�i0��Q;�,jY���X�Ii+2�+TJ�L^ƍU�V�,�*���3ra��g㡆d���T�4�MhJ]j���lA��W�Ww�.�l�v���,k1V�:{t
A�yY+`1��!Ч�8�,�f��wI��nԌ��"C�Ԏ�az&�Y�*��bf̑��mvP� �eJ��
�x^ m��/�e-� �"�	Jln$طg��0H*�����]�*m'�^�/��\)�$�S��Z5���eK�m�i�Wkt����WO�&î�Br�%�	-Cf�$Ѩ3�ShYq7��+��м��ͳL�L�
Ac��r��W/K�?+�W�֜YA�P�ڔ�h������&=�'q:�a���L�V�
�*.���{,޿��gf��L�9q��(i�чt-�ϐf
kKU�e.8�0,Jʸ�+�W�C�j�j�1a��ode[�w�k0\A��*�b�5�G�UŎ��x�ȳ���)O	�/Y��lʻ�6�:�J!���zl5fPW(-aS	HD�J��][���ww�f�{2ռ�*M�E]s1��'B�#{[@�b�uI�.��D,7���"�n�,e�/C�̗>t�e�δ('���IH��J�?o�%Ŭ�s-S�[w�6�ŀ:�v>X�[ ��m㉕X�)����n�J�)�����{4��Yݻ��JC�Ȧ*�#,�4�iڼ�.�RN�c�%\�G��@$�fG��d�v7y�8µI��W�/�d��|/m�	Z�7���ͅ��C/Y��T�Y�t�M�	�1]9�G5fPiK)C�����]Ez1�Y.3w�C1֔�h�4ąw+�1�������J5&�a`]mM�ф �҇DBbe�ۀ�iT����I����ڭ0n�R�U��o�A�R�w� ������8cZ���afI�2N���4)A7!�xn�	�AH�^�J�N�@QJ���#f���6f\��m Cb��Jϴ�2�Qb�������A8����JM����u�!s ,�$��ܬ64[fHĉa���Vn+rȁ��z��/N�ˡX���E�$�lD�{���l�f#l^e�+�"&%��V�^p�w�q��ϒ��ر53O$��^�Ù0m��O%Mpt%��Gu�W�����״�J��z�E4W�L�L�I�3Z�ڕ6���T��=��Z@E\�6�ʚ�$�&^�������1��oK�gM�ǐ<8�	@��KlS��b���-�jh2ˋO�����p!�� {WJ0�f� O��4�����x�!=Ȅ���y��7˝1	vjЧSrK��k&�*�)
n,�$k$u(�J!����Z��b�tmn�ɪ��IL �ඐ�U�3iݛ�&F*�A=����IZ,X�����YHm7v�2���N�3p]
:M*�aݒu�����A�C tf��jkm�Hރ�`d����
�֣e)��-;�4�LL��x�� PY8��˵z���3kzV�k� ��v�Z�;��ǖ�7(B�m�P����ܼ�˴�WZ���D;.m��QѰ�()g`�t�n'���X�l�v���(ṣ���	C���&^$��V:X:^VdL+��*�pܽt��V�<I݄�Y�R�K��D�K5�]��s���IC��G��.>BQ}�{KS�%*��8��8�3qu]��wM�����6X٨ �2m��]��WBM4d��b��Q<)KY�@WN��TD0Elv֑�m���YDb������"l��)��w{U-!�c�]��r�фVe6l+��{�5�g/U^8v��O�y�bV�7*�J�]\@R��20�D@�]̨�Ձ�
jR�<j��4m/P��ݓ��83�^���9�N��	���M�g58E�*�"��Fe�YJ���Zp�	��u$jU����k�6T�6��y�t��
;�C�.��n�Y��T��4 ���+)�K�V4�)MTnYUy` K��Q��KZF��̰�}@�r��D��T�EA(��3�NvFG�Z�Ăh��K�4i����Nma�,�����Ğ\9��?<�L6+7ocp�٭���Fԩ3kz���m'4f���5h �7��u��� @r�û�؛�!N�d�6[rT��)ӭY�
�X.�ALb�@�z���G^c��{�@^�"������3���4�p���y��V!�<�+ T5їZ#%H4�E�H���u��"h�wVf<kP�F�U�ct�D�ڕ��N�c*��Y��m%v���!2i�$La�`l-Q�wIͥ�+N�iM��Pk����*�2�i3�Cj��Չ����q�^ ���(l�PV�Us��R�dk[��3b�����#����D�n�%]��w75f�8�j��4%� ��ƆO�"� ��f5�C��X*��� *�3����(����kw�Xڼ��r5m���ZыY�Ll«Vd,�ע�c݊��j�#�c �I	Y2,*�p*j��[��!,��:(Z�{UM y�[�$v4l�-��a�V�j���l�r
V�߶m�W #mSƓ�.��i�����$hdT2�wz���kA&J�M��It�Bq�����7�lA���D�o6��^7w�^��J?�S�h�%�Htj�S;{@�.�/����)�AWS��C��F����T �û�4���������U�(�5�aun�w3uLZLQ!�ۛZ����Բ��`�
��PG��Wp��(i��2�%V��ni�lMN��e�ʻ@��n���ȩ(%+�5���¡���]�S$E��~ژ�ޟ��Ȧ����l�鹖�i�ܕ�E�vf�ɬ���1[�
�m�0�l��K��~�%��~hx��'v�^kÊa*�(���ĳ5֌���7F;����6$m٫���� )֓1=��������Oy���5,b��4̻,껙��ubL����|M�G�Jm�,� M ò�c��b�6�۩��t#w,F�Ǣ�1݇��t�S��
�������6�1k��S,ì萊��i�{�2�u�n�'VM�j5��h�6q(l,y6�L���q�񚃃rVA�,��(1��`j1���!4�jnK�ܖ��J�X��\Uuq��l������������۶�]�j�vi�z�S1���VYD��K��K;ub��-�.^����i��j�:K6̏r�T(��Z�\�����+j����ð�a�Z�6ui�9i[:��f��h�WP$)��4�IH�~r�m}*#B��&K����h�Ė+-ڔ��+f������76̦#�r��K���xc�3R�a�6g�j�{�Fd�+�HU�H��M�oAf����]m��ea*֬Y���rJC-2�I�V���M�ְ��V�ֽ���,i1#;���OiS�&��#���M�&��25���,,v��
�sn�R(LǕ���6�fJ����#4>�q�RB�6�u�Pw ��S�h���-����hڠC�(悭D����r�{,m�*��X�6S�����B�f�[��S��:%���������b����TQ8������{kR��;���@��A�T�������L���&����T/kd��Sf�[I��ab�w`;�Z�ԌBaU�K(�4iӳ��)�Z�N2Aʻ��T椝�;�gRX�ͧ�#���B���m@��l�ި	��t��gZ�s!��ZVU�ӹ�V��Wsi�4�Y9�S����Ϭ� 㘠!���2�=��ګ7�6�(��Y`0XrXXdbx$;�������֝3 $�*"��$&���f�QAO���nA�y�I�tT�d���� ��4)��J��Ut�,{�ڹ���a�2:�u틼M��ig,�B���g�Ue�X���*�,d@K�Ij����L�љ�m�Sp`Oi��8��)Р�8v�H���VY+ie+͢鳢�Pf%A�,	���aR��h��˺���a�Q���R�Z�
K#
��hT���|3w��t�o(�QE�G ��)�"�z&̧p5j�*�"��o7B�8Jf�$�� �jP����Ʒ6�d��J�[fŠ�l�{�-��7���M2�f$�V��F��hK�e�7�0[�^�S�[�Rr��m�B�G���jM%9j"��JT5	�pM�+T2�6ͩ�1V��.8�6QT`�ǖ\��n�̧!8�At��H�U�Bm���3V��oq�$�%A�b,���X*T*YU�f�B%1�@rU�6�D;WQ�\:٬���y�ٓ��p�Ӱ�4 	��%��)�ƴ*��f��
�X�W%��gJ�b7�MN���x��t���|G�%�'��R���˨6	f�6淦�i����M�aף����S��pS�S-g�d�c6�� 325��[� �����L�'5�o]0{L}�u�#�D#	���Qv36�+��۬�RNZ����(����q
Uܦ�3NՍ#ӻ�wh�Л,}�0cl7���ѻ>T����+���-�i���X��)ں8���4B����7��*�^�1��)
��tr6>۰�Sar̆
b�	�M[�X�n�
�2��"x1�%%L�R7�E.
AX!UD3K���,eA�rf	Cj�PH��\����X�H	����Pԫe�Dca�I�i�4����&sm�Ժʹyc�ԇҴ� ��c�Y�+JM����h�KNf���v���c���:fQ���sp<��SuR�wx
�u+`�Wx�=6E�@|+'��M\+�f�]
�R�e�\Ż0I�D`FKhL��n�j]��b�vh5ݼ%�F���gt�,6�E��q��ѣ*`k5K��olh��(�v5�{&��(㱴�bkLֈ����5(60�֢-�r�Sؼ�1 TL��B�̀��h�Y�V�Q;�^,۠�?���Q+��4X,�L���R	R	�ݩI�F��
�(�� ��/�����f	qU��M~������A��%�Al�@�H[�� -�7X��h��F:u`����:�r���sF���rŵ cB��8Cʓd�$����/�^7Z�H�;kR�.���F�Sc�'r��ܢn��J�R�L
̅j�l�8$�����+T���Ų��_a��%��צ^�a�����CQx�U[!���0V��B� wsr��+��"Pִj���`�k0Ù�maJJ*����e��=��9v��a�/��@[�١J�G)"�w�@t�6�1Ih�Ӻ5�Q ��M�nQ���*�]f"$�.?�r��t
��na�rXUv5���8(�{�iv������j��Fe�<��$Md��(�����2��۩uZm)z`.+ô�Z-m!�� $������埮]�D9�P��mS�� �­��[w�%�ӻ�JV���32]2����*�l-�.�[�� ��G�4�#MI�Z1����E��;�JK@�l��r�Ёp�m9�[5�a���^��RܩT1�Zu�f^f��@,&�j�N��h�-)Y�2PZMa��vw�0M��o�����cKB�Ècܥ�Nn]\�z^)Mm*�dlS"E�F�-�j��5�#�6�zwY2n�*m&���]�Q �a�&�d� ����� "zn�U�m�9NYN��V3Gw���O���QǂmA�R�wn��4>�7�YGb���y�����G���f�9�V�u���so������p��uq��[�V$�����n���nk��tPb�����V8Q v���;�w���U�6�r� ]�1Q�6�ьp��]����q���b�F���S��ţL�'5��*�/W�0�x���t�Ay�'
��ş�O�&F
��3��!K��؂T�6)�8����H�f6��F7}B_^[enL�]�j������Tյm�z�̮�V����^}�eK��]��b���������9sy2��y*����9πriX��C���Y�ZZ����%�ͱ�}�u�z�-]��p�a��mE ��NYc�aX�o�O��j����}G�{�q�Ǧ�4�[��L��8�1���=�e�y{,q,�����X5�a��Z�B���n��3�%Z��,�n
�yݙ��e� �^obWu1�m�ܡ�.E�� @S����E�w�>��I��|殧:�UNn���ˍ�c�rnS�y�� ��Va����)����u�.\���sޘ�����	�:xq�|zY�<��i뺕��B]�p����#�WF!=���,���m�٣z��1���p(1%W�W8�m���uw6jVubY�iwYq��K�Ϻv�R�����ut	����(U�@s- �u՗a�3�/�G*���$��wr�r�YyY�x��������b~��ݼ�N�uJu��ӅmJT,��:����ݭ�E+T�J}�\6�GS2�����:�ht6T\
�_I�^H��\��͘]v�XY��ʈ��]�t0�UoJ�&�ݾx�66�+On&�f�v�_]�N1;�v��V�P�`2 �.j�/U�ZwΡ��[^��x�'����}^���`ƞʽ�xܨ�ɱ����d���Ee󧇶�G"R�wf��0����x��kH1�Nթ+�tUo(Հ�!	W��닀�iq�R�F	ï�|GVv�Nrrk��v�Az��%:|�ǫn��(i՝�GQi�5���F�|ĴF:;}�1Ֆ�0ehj�����-1��E��|K)��c��5Φv���u�7��5|0��{�22�G����P@��nuk^�&��3�֢�八Ӧ>ٻԉ�����-j�{�N�7�$zh���7m�qog"�u��N��;{w��]Z8}�΀eyd	�K����K��%��6��N�AFT����E�L��;�{���]+6�q�\)=��-��Į��a��3���	Wt�R��r��w8�^Q��;0v���U�a�����P�t*�lW��J�w�:T�:�f�b�ċ{e�ݙ��	oDHGm��)��o3��uv$�s�⃘�*r/{�\\4��{+��"ڗ����b�h��z��`����uRfc'fV�|���`�JXU��_v����0Z�����ǫ�m�䊚�|ffCo�-��{���GRQ�@�p=p�d.�\X\�R��ݝ0���VH�&���R��i�y���^��e��wP��q��rX��CF�jR�j3�����md��g��ʄ�{}����h��-\��"[8Y(X�ř�u���[�	v𤳹]K	���,we~k��>�⻘�k�YW\��dt���]�r�cdw�7+G�2���9���C+�lHR����^vL�a�.��Iĩ�ō��B�V4�fѦ�k7���Y�>1+���h��,��2M��ޭ螼(*Dֶ�&�suU��F�'q��Y%�B�W�N30d���w�n�Fq$.�y]S#f�u[��;M�F4��/)#gi6�ss�w�8`�5��;�ƍ�T�>�Á���"�5l��}"rѺ��#��A�ٮ1Z�	��&�v��-���4���tK�J߇Wd;h��T�mN����W[�Ij}3$>�l�3tb���z�y�ס����x(�N��j���E��/��!�j���=`���]��i)mz��oq�����XF+�3��s�o4q��q�v9ӫ(]�Q� �������G�x\���V�[�l��c˭
|����V�|� �⮰i�Xs�7ϊ>���Y���8T;-�^��W���h�lt���m.2ŞѶW<�"҃��Y�� ĥ���	;�X�T>$��ݙ �@ͨU�B�o�ق��#�����R�w�"V�ϭ�p�>6-���C����m"e�y����(V�Ń��X��<[Q����W��E�ї�Q�Ѻ��ީ���-;o;�7ד&3����㽮N����N�nh��s�N[����SG�-�(�r�Is�f��R�`�B7X�	�*e�1e_Y�C�9i�ȞQv�
��Ս۫�.;�,�K�&,e�K�N�ςմr�e�G-�t-�7�[�>��1+����Z�{}�w ���{E��ɽ=�pK}�W��ûIz�g9|� #^��h�ɋ�#V,��/���H��!�ɋmP9L���de_1e�֑x�0'3\��u�MmN(r�} ꌇ��+����t�Ȓ��"I�2���vsT(�g�ڷ���ޢ���� ��Ln��ɢj�wSO/d]*�*��ʺ��w9Sv6�;B�ϧ�P������8&Of��CJqɴ��{�ԻS�gh[�)!�q���e�V�:���w����_�u�_e�$�	s+�$���̢�7։Z�����=a�^6�=8y-,��-|<s4g��lG98T^z�[�wouz��<4b�dfɇS����T>��/���Xcs���R�{P���P��W��^�&��4��W�hKp�m�1K��wv7�
%�glJާf��׶م�Q`"���u�K%!��̛
2���f�
J^ jF� J���A�B��w��B���p'����׺����Ϋ}u��N�ۧ�2<c�y	I.�g+���WQ#�y9�C)J������I��\F�/Vix�q�V��S/q�8^�R�
7q.��-Qrlu�k-�K!�9WU���+[6�%���s�ym��ˠ�Zpa;9�$\Y��K��+yd(�d��ƺ���E9dZHT�d�WhoVn�4���M��_��]�3rQ�k�r��޽v�Ҙ�0�x��Oz�H��F���ve�%l��X2��Ť��jh��S�f^Z+���ů�k���Z��6����v_n�۸.��	��t���F�9��_R���H�n����l;�ą����|X��������dk֙�U�T���@����P\�˹
�������;�Y�����E^�V�����8�)6&�:{�jI
�$��.��n,`��6�-�u��)�Iƻ�y�A����s��;ȳ=�t�� �{ΒhR1�^��3z�^i������v���{�n3�ʔ��p��C��z�/l�3��w�y�/>m�"5�����[,K!h#)XW-��	wI�V�sp�i�4���0�A#�vSkߺ�c�z��e�i���LΘ�]�.�dL��f ��rc�^��7`mduT;v�R��WW�)b�CUꅳ�N�2T��0�F���o1R��j��y�����.��Dy�����o-�Vݕ
0����%n]�b����xj�G7VFx|zk���r�1��v�f6��U�<5�]��@7֗�{4�֏\з��%`�Q�`����k0�^!7{/#�Ȯ=wX��"�ˍ�C��ι|*�Ľ���c�c����]v��4Efk�do���M]-�,�Fo�%ҥ��gTO��r�!d"{�mo>(��1�=��#�8q�X�఼��p���m67��J`*��>��ڧb�,�Dh��_YpG[�ؔ�i�Y8��Bx��ԧHu��3~׵g_�l��D���}��h�hw���;㼇���gw�н��F"�;L�W\,pZ��Ѯ���yը]+���*S�#ֳ�*`��Q�����
|nl۫�g���.b��2;�ra�A�p��n\9���he�F�}�濽��@G!����gϫW�:��S#7D��u$�s�n�&�^�ҳ�-���W]����wS�u���v�}�Ut�^Y�<(@��9Wb�6�s5�w�9�*�L���,Y}-���tgA=ٰXpkqW��V�.=��:�c�wo��$y>W��h�)Ce����}q�v6��u���5���������Ę��V0>����)i����Q�(��������V��ٸ��vM��h7Kwu�5Y������u�K-��w�
��9�o���9{'
퓱�޵��4(O��N{���D�B��]΅��,�G �i[�֖7Ew+�Scs����l'��^5��%Φ7v�%������%d9�n_:Au���ǳBp)��$̘2���zy�CX��yO�>�	;���J��C� �L�5����o@fc��k;�����v���T���Q߷FR�{BR�AeP����u�"_lɚH�o5N��9�)�7��4;�g+��,��]Փ��wt�V�/����(���U�xޘk��E+�ez��2���IÚ��ĪkR���X�څ��D���t��"��
n5�e��a�o�n��*�+�f��|m�
	<L�6��*�F�	d:0@�g�=�\o�I�J�ϴÏ�n��w�2F�GYW/E��A�n�{�Z�.�%�3b��(ռGx�tz�N���۴�]ͫʕ1&���w8;�v4���d9��G}��Dd�fT���9�&@e3���dlmX����Zn�6`&F(��s��:��Y=�R���/�'�Iaأ��eIS�Q��[�`T{Z��J��Vo���B�W�[H�{F���=	�[��v�c����q�ʶ��Lk�����rG��`�Vn�uJ]k���g��J�6n�	c���R��}�Fm��кh����q�\K�_�̖B2���yX��H�;�ss��9o��c
���m�s��[B��rC��8_]�ˑ�Cm��p�[J��֠ū���ݛ���1�d�9�a����mf�k��F3V>���fvӭ�T���ȕ��VWM�.de�t��x�љ[��h��tG�C��5`)h��n��
k�ts�X�`�֍�]q��Ƹ��x������f�p�	s̶ܽ�����ON�w�����f�Q��/<����q���`T'ѡ*���f�yl`��[�$'wB|-^�n>h�⮩t�鼀	��l+�MU�����JZp�b�;y)=z%-�֙:�5����"-���+����A��[H0i�%�.��Zb���	�|�L=)99�6Y�G�eFp�#�+��-�vN�+6�8�('/vf�ځ��Uq��kk���KBem�+�����6�j8;e.�[��.�ɥh�F�@P;���W j*VVY�>�v����&X꒢��ihv8��x�}���q[T;���ٴ��\��@���yi�͝(���!�e'�n6A����7n؝���TX86A�r<���iI����+溋wC��Ӵ`-����nf`'<��������$�R5]K^QK�v6F�&���Q����q֭X�3(]�V����s�F�wIT��/�;\{k5�{�Y+�֨�Ok.ڑ�c���O�8�T�˴�]0��.�ǋ*�
�Z�k������?������I��Rwn�H,L��Eܝ�;pPwi�t�u�����Ig�ܬl���zm�ӫU���*���"���C�6(�ī��=Z{X��I�P�ɗ�W��)v�x���{-1B�ohPֽ��hl���u��*�GJZ��s� �um�ZnduʷL���=i�������-��ys.��H��õ���m��cރw�p�0�ո�	mi�_9B��,&ÐNpT�B�'X�:�Q]����JrV�r/	�L>��C�6A�Z�h�_��K� �9ȡ�.��&?�E�¥�KI�XB�5�ַg
�'��b�����ܠ��X�(�V�#z����F6H؈J��J�\6Y�v��*gk^&�\�<.��Gz�2?N���,��6��G*�һGmtU�t-�e�W�nU�w.>G}��^�,�ك����mgn�;����ɦ�Uځ�g C�eH��M�o��h��g�����XM�:]ے��tjV딀�ţ�5�W*֩׬^���И��pd{AoP�����%�+٬u4-�S�ޑ+�.;4t��I����#�d]c"�HK瓚mخ��V��F�$�3O��1٢5`cK�'�����a�M鵰�.�i��h��+�44m�釵�ߴrz�險���iӮ�p�ȝ+�i�LK�l���r>n�ʦX�ʝa��v��9��_$��v i1���ᗾ�<�ߴ0�MG�$#%�i�����5@膢��98xn�Y=���v���[ۘ|I�ݍ�H̛�/�8���
\��hQs��wiJ����MHrf�\~�5��.�0aZo�ڦ�7>�n��:�� e�� ��;	n�Z�$vs(��\�L;�]8Ϣ�����X5vv*��z������ܪ��Ϫ��t��{�k���⼃��X�T����0`Y���G^�:4��]e
�-E��T"�s`�[��w���\H[�Ϟg��&<Y1z��e�qk������³�L�c��[��C���e�&]�W��3|C}�Ow
��(%��_��<�xYbG5�#�+ �z�t|�|������`�+ͻV�I�;�G=�8g$!�*|���n'l��d��I��,ձ�*،i񽧌�lʾH���,�e���+瓃�Ћ����#�U�z�q���0���h�t`���Ag�Ĭ���Q�̳������M��Y�=��-����[��:����yx����ED���XO���er�p���2d3����iO׏�x��7�u[�� �����x~<��<=�T��ܨ[5:�j�M\W���6��`��S�
����0�噖�B��5k!#�z��CJ�����H�N�ۜ+Ax.n���'5V�7�1p���aW�H�sp�}������p�������_e8lKM�{�
�@3�tp�^k�+So�����F�Z3k[���(�|��XP�Ğ�̖.���Y�+��%w���l�vr1a�r�]��~#j��w�]�豨&���I��6�X��a�""�su	�ꎱ�3;u��wmnK)��׀3w�^����vQ¢��ᛑm�\�i���� ��4���L��&h8Ы{ٯ��x�7� �7\�c��}�l9��)�S~�Z4�C�;U!!'���s=�O��rJZӼ�����r,�,y��6�!k}�D�wwB�c�mi�#)�c�%��=��1 z7]f�M'jP�߆��9����a�דBv���J��ľ���1Ʀ�A (Kb�:XR�tsfq����X|wT����I'O��ؑ��x�2��f_*���c)Q�v>�Av�vj�yWW����_��F�{Px�����L�h �NX��Q�ڶ�;z�09���Ĝ�����Yv/�7hT<��(���k�=�ϲ�bN��s�z3�ڥn'�@��G,�{�u��eE�/ke�3\���p�;�e�.CíiPI�a���Ф�W�+�.�X	YN�㺀[�F^�PV&��V�RIXQ�撈P�+-�L/WX4mZ�i1�)���_p��%Zc	헁̍՝	��9fQ���sN�?]3��g�r
����H�j��A�w�r�,�գ�����0��pq�}��W4JƜ�Nr����v�G.��U�u�G_���|sȏKc�z�n�k�}e��G�%�	ؚU��U�.��GU�ךa�ud� A�W;1Yf�Q��\�ٲ�B��ɜZn@���[�C�q�71��[rՁdu���&�Y8��8��I֯��]�R�c!����1HBײ�7�t���y;�����S%p�wPWp�KH��`Z�,M���Cp=�; �yoD����+?Sn��+�K֐y��y�/GT!�i�GC��=��a�'vv���M�B�D��͙]ݘ0�[��@���}±�J��vK�4���@�d�(� Ueo=Pp��ls���( �����ZK�dr>�Q�{=*���1��uv]j���dc]02;}�"g��;��^v�-�v�Si�v^��{���l�����]��>/oGd^�	�W\�a���y�v����#.k�K���[QpP�h3�|V�X���;J��������+%Ū���B�pfC)j�!ϻn�p9Y`�bSw��GS�	�S�Va4B�P�z�>-�c�s-D
ä6�`�t�%,�o\`2���<��U�n��jU'.�f$=�fbyiN�g��	{���j�'r=j��I���sƝ�� ��/�6��͒�6��hGՈU�l}1�Fޅ⥱'���ܞKN���l��Ǵ�ǥv1bոŃ13Yë�S*�N�Scy!�l���X&H��x�iw��>��i�,�f����/-ow0�GD�>vW<;6���va@c�k-6䥂h����d�"�o����:x�KP;&�f-����	��
y�-�� ��\�;�O��Nbi�R����>�<;*7�Y�ӵ�1B�8gݖ��v��S�7�Kf��#�[)*v3[��/N%)Qҍ���&�؀�4رQN��ź�U��=v-�.tW�do
�j�]�{{�����6�W�x&N�6v��6��s�v���dӹ8�'sVst4jU�ʁ�aǎt���B�P(̗�Kl����b9n���O#�T�-+���\�7��A�CE��{R�R;a���w�Gr���+n���9ɽ�2H��K������:��5k�\.�����eO�@14�0{[���㫩o��)��qKN��H�b���Vt�E�]��f&�LX����R�>X%e>:'�J'�Ĝ�����Ͳ�}mZ��ӸA钦��v��9s1w��cO�"�!�� �ו� .�ƕ�����	�ҞpMʲ�U�'$�;F�zu�&^�ÇN����iӞ�	j��-enc�:�ڧ����2��l=���o4���ONE��kn]��.u�r�q�js���XzHڲ9�}!k���qh��B����H��.i�b7s;9S]+^�sO�eye͚ask��@�:�ϳ�/^%K���+���R��u�e�!*�.��V3�����][��ϙ��:b����=�� �
K�U��>	A]�e�����A�F��;&f�,�u��<}|�'R�t���-�r�t4���X��OnNn� qh��ũ�4ܰr�����*�9q�����Ot\��@����|2��0�p�`w�7���F5S� n������)^�1b�J��i��P�E{w��).�$\��C��s���>��Z��>�_3D5+�-��ѥ�F�iJ\���F����Z8�'ݯW1�]�y����GJ��:��4��S|r�#:�Ţ����ѳ�*ޗ`г�Ϭ�.�'���;T.�:;�9��ęS6)�U����3^	v)i�7Ǹp\Lܖi�$��;����X�%��#�б;vz�4�� ncWY۰��`KYO���0������'g\�:,��3�����N�c����COS�A�:��
�g��ՓW�n�?lkGɡ�`��_s���� z��ޏ��]��m��ܒ
0B����x�䳡Ǵ�Ū�;a�´=�=��n�t3u@�+/���Śpp��^���I�:��J֭W|�S�$u<U�Uˢ�Ctw;g�{P;t$C-�`�`%��n��Nil9�v>��H'z�/mle5�������3Ӌ�{�lo�j�"w�Y(�,[�	r0��Ή����aÒ�<X^s�a��:�F���& �ǠdRֲtVM�uv�
os�e��)#/`%C).q
6\�&�U�H��Mcu1-(	���fn�L�P$�3�ozK��}w��-�|�-.�L���B�B�P�Y7
*�Y��e��Z�����q�\��^M��,�R�6�e�\hY�)^��W
�����SZ5v��/�'Y}�����."U �>y1�ߋ�F��\�"��tќ��(���G��zܬ�b����`�?8�n�yb*��
������ŝ��b�޲�R	R�tkf�Q+�t��0X�s����	xf���ڷ����ɋʒ�[W��6�VD��6h��(w��w z
p<��"5�'׷Vi��+��Z���]���Z�.�D�퐮���X��ԮU��Z��YEL"J֨��I9�el���Vɂ�g˛v���q�����H����Μ�:�b�������;2]<TIN�ȯR�*�BS����
�ݺ6��Ū��,��;;I�p��J��#SP«�>d�-��8{O�Fc�Ϳ`�A��M�J�{��i���1r�\շv��"�>Kh���{�|�ѝ�\s����q��q�#,;v��6zƥi�>fo`�����ђ�	�!#�kٵ�x+3��'؋�e�5ڂ�b�2��_�b�\��^���,wX&��wKFr�hݗ˦+�׸-�6���MFø�no�9�I�wy�!<�SH��AGkT����n�'��ї�vS,�<)०����d�zq��;q]ֶ�G��؇!W`LV��*=|�8gsPͺ�N�yo���t�N���i|�X�	Ƶl���e���լt�B�K@��4�o�0�Dź�{����W ���m�x����a�-Nx;*n�kA9���q-*�ůtjѬ���{�x0Zf�T�o���@�w���t�Ĭ�4���K4N��u;C�}��J|)`��۔��t)`�F��K.#���T ���iZ��7:q�w�k��mN����dTƶ���ފ��V$���ok�A�Fh�wx<�Tz^��Uʝ\�\�윧��+]�rScj�B�6���Q���y���ډF���s������
��	'_G�9X��vP '��էM��A���d��Ȧ�;/��0�Jq�wZ3�ٗ��úKtD�4f[�Ӫތ�BK.�܊�*�M��]�kzr��>���;���
�oZ��k�C�+V�v�3gj&\&;�V���v>:�!m�kTǙ
|3	��< �¡�]�41�{��u�W�}[��__��C=ۅ�p�������e������0�ohV�5V��Y����\V�'&.�~FXA 
q���k�^v�@aŖx��U���)��Sl� y�vt�n����j��Ј�>�H��ǈ��շATY|2�v���۵o>v���un.��옠�ũ% ����_;?FZ.��[�
��=Y�-R���v��X���;�xd�~����+���;���d/z��/��m�6T��Mnʮ8C.��m�^�&��TT-"'g15T�� KV7/�Щp૵�̂�v�Ŋ�����5q	n�T����ha5/����ĵV8�Q����9r�-�ņ���fa��[��i�q#`&�P�*m;�����P��F��);�i>�5�����'����_�]kU��2Co��Ca*����^(U�0���o���b�Xt{8��YtQˀ��W[��3Wu\�7��>�A�h�X�.S��.���Z�{����!����+�]@��k��[(��!�l���\h�5�Z�}tZ���[W(�n< �n�<k!#�)��V4VS1u+{��������IE���/uәk�Ң^������٘u5��y��[��)r�)MS"�����C��nb�P��M���^o%�J��(���RY�.����.(��ϻ���޹Nj×0V/V��;�������0V��ǝ�_�p={�8��Wˡ�ONf:�X<t]'G�O�fALC7-�f 9!��IH���Fg�T+�Yx�x��S/�q�8We�
�bך�4�`9|K��=�P�a^v��Hfb��t�#��T��"�-��{8��!"F����ٴ��l�[Dm�Y�S��g	ΟZvQ��,R���\���EF�&K��8�G:���nCgZ��L���9��/3��|�ܤ,\ 7���Ō�����}s�:l� P������؊�ED�[�pǋ��r��i������:���^�n�v�V,�L>۳M-HBL�Kw��gJ�_6�pǝY�[��(S�ڢ�ū\�*��OUI�'I�vet��+J����a�b=y��ȞwD��%�d�.�tᩯC�H��|� �ܜm��@ī,G`mA�n2�X�w5���uF�jφՍ�.�Z����ا��(պr#p�bf�2�.�Zb΍�z�����~0����c��n��^ {�*��i�Zج�t��lP^<��oZ��O�¡�C�*H�bfM�뻽c*ҍ+|�tRWa�VXmgcB���.��_U���v�Π��z���|��xp�����3[1�+������/7xJ4���Z"��w��\w��=o�o���3G7n+_6մ�M��������ӏ]�Ҩ.�5/x^>�&m܊n�� +��t;/��=]��l
슭�pw�����U�"�)�̻0c�U6k�1��g�秷+��w٪'�^�����K��,w�B�����Â��~�c19ݘ�B��۰���^·H�|��8O�3o5e��e"�l D��)9��uiV�*�E`�Q���<��M��8��)tb�el�땫��93diC���8��M+��]�o�t�N��IY:��K�z�9�Q_<�At����:"d��0����F���z�v���\��#�������`6�Ś
��s�DN���q��żBnW"�T^`w��S�Ť��o���=�<�v�\8�^`�o�ݩ��q1�u�	ID�⠑�wi��uޢ 5}��E���]f��h�.ŋ��)k�ww��;���S�o6�WV9.��v��s�M!r��b_{!�e��"�0�2�g��#nM\Co�Gs�a˻��/\���j����墆h3�R��ͫI�v}w	��j9+wV��y� g�3*,\�1�L�("��pf��ݔ�3�j���W�;pj�*Ĝ�%V��ƺ�7]Y�s�$^��踺Cd��"��+��逜��ƃU��U�}��W�v��*@�x�d+r�Ǐ`��.|nh
N�m��b�8p���f{^������n�� �m�I��I£�ճj	o#��ί0n�M��
#J�����u�U��/�7��C�g�*�j�E�C���؇U\���j�U���@k�叩���A3+������f`.�o7��71uk��찝ٮ�|X�b�{�)w��e��,���o���ܹwͭ�7tf
���R�߻�n�I�dL����]�I����\�6²��j���scg����T�A�{�y��f#v�ʜ����j��Ԉ:DWdד7\"MKgJ�g�0@�����3f�$��yU�sy��	�E�f`
�v�r�8�H���;�W��J�	�Y�M�jD�(:ppӋ:h�њ��=ȮX(�����0\��=��nb��a����*xW�:�=�`���_H9�X�����M�Ijܵ0ԏ�g{�R���w:���.�d�+�&�@�
N�����̮˫ ��՗]W�^��_%+�X�9��(Htآ8�1�D(*V�NL�tiQV ���a*������ã�~�H3A�B��x���7y.1ͼU��BDk�S���{������ܻ��lA1�ifnB��{�W^�l;Qb")��,v(N����p��ub˾� 跡�N���(�7r�q/���lm���+���� 1J˺���U�`=8�jNR�)ϴ��Ċ|q����qb�]iPۘ�3o�;���]W��sb����c[����V�]��[��E���`i���ʶ&gN��X�����{��Fv�t���'ƆR�|%8�[喥c��D˓�G���T�H�±y�f��I̞u��,�fhn֢��"G>�1�M�S����]�u��䃊�(��?-�46�&�Ji���K)9R-�QY;3��V�]d�@�r�&�_'��E\V�gHt�q���n�\��JAQ��L��6�R��%q�G̫F]�*��!���D��s�-��#�Y�$:��^|jި/I�������ve���-��LQ����@�[g�����y��m�i�؈4�]�7Vʊ�z��sm��t�/�j��Wg s�7M�h��6�ƀ3�A�	���43Q�GjoA�*�>Ӑ�V��e�9۔��S��Pd�v��!g���i�4ey���*k_MG�٩�mA���� /1s�`��1-8��t��2ɨ�����r������	Y�`sG��Ah�}��z+æe�h��we_]y,3O�t�����3n��Uy����w�ν�̼m�D�Q�>	R�H�b(��������RAAMDU�T�bum� �������JY���'N ��l�RD�TRDSM�QME1ATDlcY�[U-Fƨ���"*���� ���%"(Ѫ �h"��Z��hb�d�0U1SK��ZqTEQPU&�j��T[��)�4j���mP�F�4S�4�RE�KBQUh�IM:qU�i)����SKS[��m;f*"
Jij(�f��CM,l&����5��m5F�$���jj&(����u�X����
���d�:�D%ST�M.�h�EUT�"����4�%+TP�Q4Q��$ H	/��ʷ������l�=q��2�E��З��ιv��Q�G��x�Dq����Ɓ��.:�T�7u� ��-�<�y�����,[CC�ʡ�Ru�q�j]o�s1|���DA}L![pWSޙT���j��D� �/Z�W��څNNH���g:pu�#��z�z�/Z�͑6�g�6���Nr��[�����W>5�Z��υ��ҏ����p�U����W=k�9�V��֕������S��^��ՍBJ� ZԅBy�tv+��hJ��sܦ�r�2��������`W׭d1�K�p�gΧ�����K�q�®ҡav�&���Z��>����G���'d6�+�d*N�^o�r��0΋ӳ�Hqg1�[<fD����}�pW:�^Y9��@�v>��7$R���S���=��A)�Rg�5/��Ͻ\��r h��\�u�W�xk��Һ���PLm��wGN��-��n8�pقԱR��� �iI\7���g�1�r��e���Q�>�^��+��|�=j\��k�nVH�!)ղ
��@��b`��:y��|+:�g/Ef��K��U�k�����J[Î%eΫ,����2�(�w�.�����(q��F���,���
�{'g�����G��z0���|Y������"^��;;t�:��i�'q�Ux@--;�c�e� �!�Z�97$@S�����U�A*�TF]�B�����X����<�ê2X�)�!
���.�=M�d�ܕ�{=�_!	�1ȑJe��g�W�]p᎚��{,g|�wo]�����{�m�ÜI��ϗf�ҁ����� �¸B��{TۍWhI�AAn�1p�Ʌ6��P{�0���=���L��P�.C ���D�&Vӣ�R;]�W�����T2jo����P;iIl;��w�:�=I�>�$��֜z��Gy@X���`��C��7���.���-�!ɘ��|�������UZ)�'�t<�<�MBJ��\u3k�1�6��د1�z����/p�Wc��FR�:������N�c��ɨy,N�w�n8�3����C���ŕ4�P�6�8\���F	�l?��i1{��&�	S�\�q����;Q�b�sʜ<�29��]�$�������%���UHt�j<�*��րz��
\�3��s1���8��˾�s2�u�nw��ԋ�s��٘xj
U�)��a v.y#�6#�M��F��<F|�X��WF�Q�n��a��y����2y��&`�ycP��=��E�b��۠������9�$7�ފ/:�Ж`С�N���0�9,=@�vh�Z����]�ۦmPB<���Q.᤺$_#��/t��M1q�W��u^\���=��m�g�話`u1Z4��>).��u�힑�똆����@��\꣚��&�ۚ�d��e2�b_�+s�7nG	����T�I�N�:��Ɨ��U�s�;[Q{o5�:$��O����e��5�:z}d;T1YF�U���c}Ⱥ�5|FF�-��j���n��
%��w���.v�׮!�X�|ڸ}�g���Q�-g[�����f�����xK�\�Ⱦ������wM�	�*�0[[M�r0�1���E�mk��b 7g5�%h�K.n:(�.И0�AJ��s+2ߥ�.�5��o�K5ط�9�b�Wfw���X3�Wa�ĸ�0WU1(���'P�x��U����4E���yz���u �~���cc�;�pC�U�������2J����L���΁۳&j��t���77�����'0��cZ�ry9��f�/��S2��`��8��(�%7�!	�mf�s�GE	����+M�tCg�ɍ杚6��|5��})���yf&i'ʸ��N�t	��ɌV'vejS��V��(���v83/ �� 꽝vڝZ �p�0ȃ=x3�}|�qL�=�RH�k��3����{"�V�W�*)��i=X�;}X�ã�4�I�Wl�w�Ž�	֝���X!��XGWVNs��I���f+�n��S����к��uT:`9���&����y��k����O<�G�*�=�@=��!�~��9��P����k�S��f��r�<6,oOV�B�Ȱl����!R�o�`�2��:�N߸��X����7�_���ל�vӼ�z������k��7]D���ޘ"��l�B�?�����[��*�,�� ������dC[���ʫ�d�
��&��50��u�)^�`A�h��I�� ��ִ2t��:���Xچ"���,�t�슞�p�8�}���B��3K��<b���V�ţ:�9��Pp*O�������,�k���X��#���f���0�¶ch��ђ��m�3�(}�4r��x����޿+���� sw�>��a��@=�##�UC�Z��e7�Oڼ�ϡC��88o�p%Q���|aTm�Egˮ�Y�Og�T�:�����tW<O��[w��]�\=ꑷ
��P�@�d�!b/L$U�83J�$��Q{��4�X�M�k��]��|i�:�t�#����e�JH�~�r��^�tb�s��� ��a�����s0�F�K0�l�^���W܊��N�Vk�B|��]��f���4��۞՗����6f�D�U����Z��*	���̋�Ů:�����qt�6\���#k��e�>)�$�[Di��D�]��s���+�a���շ!�\=���
��c	�-�.c&��:�d"JS����|I��fA�����ms�ď|�NLc�3�)a۞b]L ����S%s5�L*U@���JR�F�捊\�!�,	��P���P&^�@̍=7�2��~�䩒�9`kp]ډ�3��J�E�U��Vנ�逈v�+���G�P���kڗ]�������8��T�,�uWFJ`;Z@���{ʱW�c�m��'$GEڑr�j�B�B��M�ot��U����ډ��ϕ��@t���?m7�b��/fpC�M����b�k�fKyP�Vb�U����)l�R����N��Ϊ���MB1`�Љ��6M�,����Y<�b��`��*z�Ag������d1����ۏ�/����`���YN�!�)�H9�~>˧���@ox��
�:*�Dt0 &#�_3#>V��-�&w!]}�kB�Nbd��N��6�9թ#X@���OeJ����}�(`�KE����}��VkU��ʹu�NSg���g�#��\|�*�qf�Ƿ;��|����Sz_��c����k�Ym�w��/��4ԥ�Tk]����VU����q;S�Ljp̝#Z=^�k��'��BpW:���u�P	gÝ���7$TB����;3]F��{�Y%��|�e�����ZTs�V���=�[C��hiZ�V���މjL����Ŷ-[񴫴���ly�����&b�Z�4���Lh@��e0T+��Fq*-����Ҝ�{;��.v���Ie��?1�:�&�W �X�'�KI)R�n���CZ����5n�M�5FP8��mV�����NX�㖻H���i��%�����T�jd���N6ci�=.�Ɓ��*���Ċٔ��Dr�\8c��!���']Ľu��/�̮ǵGK���wmM��`qZ@�aa4���f�Z=�__:"��˾�S�1�T�!��f`Ko�����]�qdϲ�C� �������-��B5P�p��������RE秸p�%�l�=v��ҳ2,��L�� h���F�kO���GyB���Q��r�W;iL��K��/�j��Kmu�6�����jw�	ΠTɜBRX��fV�q��1���~^;�ju��c���IwʆĐ�_0[���I��-c�LM�U-0�Rl�M�褺�[��93{�'�T�Y�9N�VLG�c��9o�!W�yidd�J�&�4�\��}a�"u����Ϭ�&*�t rv	I��D��C���3�>�s��H�����<+ �ziu��Ϲ;�1��~ri�;q�A��b�*�jfj��{p��#��0�Q\�L!�;���ZL^���\BT�#:ac���eX��.�鐣"[�����1v,+ ���C>�U��;������0Τ ��P��R��N��5�^�˯���zhְ��p�/�b�M�	5q9����=��XQK�O`�@	��s�;<&����(we�R�pm.'ؾ�Ž�mVŁ��h�g���8�C�?C�t�r��nR��h��N3m���^`�D��O2�b:��w�U~�\ۖ�ȝi �Xx%a]�1����e��KW6u�Y*�_P�����k���/�)�����p+Xʁ�3�����N���(���,�ift
�|���veJ7Jb�\鏹�t�d;Pڸ}��~u+0��U����!��J�2��{�ȿ�f+jb_Sy�E©c��эdY�u�Nw����<���ϼ��`��B�a ��03֡��F'�n��pD��.�ꗼ��(q����|�hU�!�{�i�[��x��Z���z�x�ƨ�t�|�j�+�l��#oq�_K.Z���x�Ƣ~��Da��M�6qq�^y��<��+�厁Q?���y��
��Ծ�L綊���u<�{z`���Q����!��9�1̡(�������
U��[��*ѻ5�fi)�I3{.mthV����gRD3�* ��7X4 �2J�$�t�<#�e�B/)�<]�L:�b�򳃟��f�oIu�7	�p�4�|`��̄ i�31ϰq��r��*(2sk�>�Z=4��!�e��/M��D6xL��i٢و�
b�l�2L�C�y�����)SJ�̒�����i��ubU�?awX��v���6ÄXf���8W�hi�x6�rq&MA�{�a�^%���
�z�:�#%���Ƌ�XX���b2�ӡY�f��Ջoh��p�������:4)՞' X�Fd��A����e3Y��;r�E���;�Ѿ�$�x�s���U0���n�TDj�6i�B?t�#4�v��J-��9���NQ8Yو��}p�!Us,�1������M���dٲP���1x��9��zS,ޝ߹�U+(d�H��HmC��,S���Y���ʳ��|G�:�B-xS=�i�M���]	�T�i"�ܻ�\�CGa�-jQpv�{jr�ӎ���5�f*f��UȮ	�,P�/f�����j�r��˜G���s�q�l���^]�Wn���{���&�iQKD7�)1>ӹԥr�z6��=�����P:p]��u���\�Hk���X���3�������lr[Σ��;����eJ7f �.3����bC�:�� �����{D�N��7�Y�W����-�N��c��>�J��-b��R[?bp�WN��x�<����1Z���<���7�.X�Hs�|)�^ۿ0|��ۿu^&���J�a����O<c{olV5�j��R{�p�+����L1�po2EǺ�Y�OS�ke��Y�b�(������<7o�ٝg�d7�-��ة�f0���ϋ����9pꙑ_)����S-�W/G[z�4r�#S��$L��4/��1�����+�K��3�ڲ�L������[���3}��R�	�PJ��-�ME�"�17�H;�֮CT��K%����k��Y�����zV�^w��dT{]J�O��
�[�K��ȫ���\"�\�ص���ʚ�cZ��A��ʒ�j'L�����Q&OR���e���&6���g��J3t���⯌���Sw�+Þu>�5ȳ��!�V!��Tcq�p�g��i[�s���f�d�s�dJ�p����<v�HW*���s�Y\��;ɀ�/��ۋ��)]Pqf*v"���]���;-KԲ�K�B��ڨKf�S�#������w�`q�lG_�;�9� ��@�?m|�]����HC���/j�1�]WШ���z?H��6�^:��gx�<~5KX�C7�r��!d�U�"
�>��
6gpֵ�_oO5]U=ō<6�(�BQ�s�P�d1��\1��{�7o]�D�~��	޽>�s����
O\·O�va|���� ���22��T��2L�bڥ��ǋ��{��s���r�FnT�(�� ��&	�K'iH�Ý���7$M�<�9����Y�)���y��b��n}7_L��j@��+H�"��Ǯ��ҵb�S8�"I�V�2l��<�)��=L|��u	�R�1��Gp6LO��N��(C��:}�����靡�%�=�hvc�<jb��T��%���c��p���*�#��ŗ.C
RGeM��]����ӈ��2���[U��Su�e�69k��󑧯%���B��;ֶՀ�&���M���9�DLI���ٞjwa���\8c���6X�N��������]��6�?f4��bZ����N��Vf�V
̒��ǖ��V)��u�­܋DB��M��&��S�4��K�
n�3cqBW��YJ�^��3p��+JWS�z���(�;�Ӭ�s�h�'GW�����0����W1Ex���%��r�`�i7�5��ZL𝺤Y�sه&E��W)�~m��.Jh^���	}W|��)q*r�R�au���)���v��+�Ϸ�=���xc�PU�T����	���ebC�{�nߕ��_;|�!ۼ�d��«o��hr�NE��ŕt|�X�c��.���Ye����i�mfͣ��m�bX���uc�Z��ٿ�6���Wi��� ��Xy���,A�H$��)řt��+��ѤČ�rVY�.3j�Xñ��IԒ�̻dh����'.����8�j������X/�1��t��W�cp��N-�ڗX��l�yYN��Q���˱_E�w������ĺ�^a.��w����۲gf6�a�H�j��n����wH��5���݌��$Ƃ�W)��ۯb�0�-�e^�w{�L�%:aq�6��y�X���w]z{Yľώ�U�n������E��u��C&n����u�L��Kd�g�VuuK+���X��[.T��ww���<��G;��}�)�t�Gк�	En�Sw[�]�1�ێ�fPO�Wl�<ުy^�K� ��"V.��e��`SX�ДU0�*󊀒�0t&��� jD="����N�}��;G^�^�!%N��P��Zj2094\���J���{9�:_trY�
�Է$
���MT��\��-�z����X ����v<����$���K�i�D�[�a�.�Z���J��6q�Ye�ܣ���A$:W�҂ C},��Y3�����y�qp���P41;��ڈ,�݈�G�j<f\���B��ÉkIQ�@���Z��F�R�[BE�'˴۲x���!j�4*]�0���4;N�c���VQ�g,���k��T*�g�{�L�t&���-�ʋ�����.�/T�S�d4w�j��g<���TC�u�y$��=4q�/�Z�)�R={�N���i�3��Q��m��û�&�����]\�+�����],�����°.j��h�{�e��ǎ,�!B_����rpUW>�.ѭ�x�l:(�@�v�_b���=����{72�D�#���6�=7+��4��)���sogmO���w�1ؓ�r�p�	t��q��Q�+X����u%s�{p�
S�R�g;����d	3�f��fP�[�(:hd�X��z'sK"���9���
���C����Y�U�f	����9y+L"�E���-���P�&ެ�lva�DvB,ݾ��1�[�dۓm���]�n�����"�c�93����n
�� ��s�T��5����t!����Y���
V���aغ4�%믿~�s��Ccd�֩)�]-��MQB�D�UT������EDMST��i)B����������"(���

)u�B
i�������)h�F��� h(�* (*������i�"�.��))QC�)�4&��������-��kAl��)�t"t��hM:"њ(hКj��i*��ֆ��.���R�LZ4% kE%�q[	��5lh�#F�Қ65)lhKcK��ѪSMF���i�ִ�AliQS�֗H�8�:4�؀��1T�-#e��"h���*�:B�R��)6��Ѥ��i�(	�jj�ul�B �UFΚ����+N�B��փIA��Gj�W<l�:�4�6�cŎ ��Za3e�=��3���.,��AU��E�5�AF}���͹	_)�5�n��k�G�i�W�}@|��b����H	T}�E��r���M>^A��W�y�����ܽ�����������p����%��%��ϝS�t��o���`���"#9t�N�1����C}j2-����8}�}�.~">��K��o�{؝��v��p^��Jz��d��ۓO�(�!C�9h�/9�����d�=���??|�u>C��#H}ܤ�I��y�4qw*ˉ�~���(�H߾�",G�4�z=�Q������=��������;��4�wݯ�s�P��F�������9=A��=@yr䔗M�K��=�Oo1�N�B�^G���wx��������V_�|+�ŋ��H��b$z7��GS���������%R|<�΃�y�����>���Լ�{��;�I����ox���~A��~�+�^G!���A�>��KV}� !�]s$N�m�̏�����:~|���ȏA�J�Z��O*B����?o���?�>�t�ےy��?#�J|��=�ܝ�`�%z��륢���O~�qz�	���|}��G�D3�+ڙ�ؽ�z����B��K_D%ӿX�ɼ��I��P�u	c������F#���'�?��8A��^G*�9�k�|9���|�i�]��;�}�G�%?�~���!�,��q���	$�G�!z-���S�D�ur�������ʐ�G��,�IC���{���rNG�>�p:��|��n_�A�K�|{�Pױ�^A��p<�?��g��߸���4�wϾ�ԅ�h�������rz���~~�F��ښ����R���b"bG����ˡ�c���'�:�
z����;��w�?�:�`���}��P�������P�O#�9�4?�:�u�`�r����i4�>�����1��60!T=�7�8�Ԫ��#�G�"4������r_=�	oe�~�����1��>OS�]'g�����<�{��|�\��7��'�~\���~�p�������N����ϰ�𼫇���_j�� }�B�"G�ϼC��M?�������{|�S�ܼ���{�ϐ�G��1����4%�g�;��.���9�����|��W%�r���y�5�����������j�{[\۩�)`כ'������t0��\MPÁ30�i�F�;������]]�ִr�V2R�ώ� T�L�;��v+a\�8R�,��]>]�Ꮄ�G�'��L1m�[�;)d���>�i�@;�����}]S#�ʅRR蕛�ЯVu?�B���<�þ��wBW�Ϝ<�����O~}��������w2�{�:=���?�������NG��x��(?��3]��Ht~���C\�׼�>�6�q�6CTA��Y��o.8{O�.�Ѥ>KC���O�\:���>K����J��o_�R::��Η��ϼMC����	A����/޺�t�`�2�����dq�����pr�]��4>A�����r9{����i4��?_�������\��|�I�ϼ�p�[�z��'���ߏ;�K����O�g�����D|,K���8�@��b��_�(G�}��?c�z�~�i�?�/ �}��)���|������������=�B^a4tsyyw�y��npt��/<��s�p���y�C��.���}�f�]/E��:Owf.���[��� ?%�z���wK���'�=��>A���9����:�A���ܝ�~a4�=������:����N�l>\����]	A�c�0w?e����8O��NG�}��ԭ�n�����}}�z�} }�4|r=|����w	A��z���9/���_phk��^sހ����]�||�����i��ܝ|�hyc��^\��9|�;��/.O�c�S���������G��c}5)vs�u�z8D����G���Ρ�G �����!����>;��G!)�g�~��>�PrC��A��{�:���9���y���4�;<�Q��=]C��8'-/�H|��1̗߄o�.g&s�?����|]�z���������/��Ժ���'�o�~�'�켇����?{�w�&�a��_��w=G!+����Oc䜻��|=���c���p�̅�x�g�2�޶�ɧ��1��}�#�?y��rW�9	O��<������ޏ��S�.���|O#��_�'��~�ġ�}���|��	C���}�R��>�����^�"����tG4�U�M|��
ڿ���>�Hz#����Е��O�0w=K�������9'#���GP����n�}���������'����N����c������Ɵ���?%�>������~?O|��]�3nr�D虌���07[�3�{p��	v�g<���ښ��C���P`ś�ҵ6��}_Z�Hf	�>����E�����#X�u�zn�/)�P���
۰t������Dq�_��&�5���y�o;#+�O����z"�sY�o\=;!y|\��)���;HP��y�A�i|��#�����@r�r�%<�A�=��:�T� ���A�O�s�O�=�GØ����/���{�g�9/�wǪ��Dh�1/��Z�
'.���U���G�:��#���ν�����:�]&�o�}����=��%^��9��·��]o�{���]�}Ǳ�/'O�;O�� ���<���9������������a8��U�:Ϋy�[g�Yg�䇩����I�9'/`���:�h�����G�>B^��;��������9�]�M?����|<���!*����N�a� ;ؽ��yS�.���#�(D���#��]�,C*���q���(|�_��c��(��;�w���}�k��|?K����u����a���{��u@v��C���e����8s�{'#�����	O�G��=��B#�T�ǫ�j�j<e�)G��`rO�rio0hk�yN@}�=��γ�^C��n�u/=�B�Ͻ���K��0��s�]�����rRS��g�8�{�욧�p򏘏����w{,0���^���ןz������O�G��A�#��w����=O�rN��&�C��y���s��:�K��������?]��ԟ��>A�J���<��=��/4�?}�>���}��M���ʛ���c��������O�xà�e�}�ʐ��~ܾd�_p�_��Ԝ���{��O�r9'/'\��Z(�c��!/2v}���|�������ǁ>�����ꅋUzغ5�r�js��A�%Q����/~a����~���ǲ���xw�G���{�������Q�HP��r�^G?d;?n�K�_o��vu���.�(����^�G��m-ގ�-�.�]��G'侞~��bi���y߼#�J{��x���}���9S�:�'���z��C_c��x��u~O��]��yQߘ�z�si
��JF����"���5��2�kqzz���1��>�C��>�]�IN����#�rO$�o8��~�A�y��C��&��y׼{��=�B^�q����}� �s��I����y��\��q�wz}�@B���:��_\IVq��F�n�6oM�A,�,�#�x�	/6,'�U�eYVV�GU��y �i��f c
�}V���鲮���]`J�^�oL[�i�׫+�6 �f;��czc����ٳ�)5�%�m�Z2=Ɠ[w��_���c"�#ȩ��D;�xw����NI�9|�����pu	Wܝ�~������K�:������������7����_����T�����w�o0�<9�=��䜟c�l~�>��xD��C	�kݘ�6N�i�N��}���h�=�w�w	u�߹z�nC���=GP���J9��9	\��.�Pr|����~��=O���pF�e�}�Ժ`��{��� � ��VB�!��5y�3v%�w�����y��y�O�v��~�;�4%?%�A����uA��������vl�&�#����Gp��u��w`�$�>��uS�:�'Q�c}��#�;7>��t_z��#-%���� ?F�_y���=K�~o�zN�{�i��`ѥ�s���8��w?%�|�=��IIN����c��?A�ܩ
#�r;c��a4���X���$}��tz�Ѕ�ܳ[�^���?g�>O'�����BuR}�Og��? ���<���~��~��Ri4{w�U���9	W�}}���!�����/Q�����@{����$����������w��y��c�~��!C���>�������\}���9?c��>��O�{���|��*��sκ(=��9	|?y�bw?oa��}?{��!)����;���@vy�Ey4=Ddw�q�Z9���վ����z���伩����h�[?�S�.����uK�r�(���9{}�+i�{�q���R�b2N�؝X�T�œ��r;�P-5����ƀ̣0Ĉ|P�3�*���=����x�s�njW/-R���H��g~lOE��yma���B��a���8�ݿ��d�ۨ�1�{eߚ���MM򻈏V��yn}�~�����Q��#B�ԕ�s�X��s\�t��ch�t9l�{���+���ɄN���Y�DN�0������4�Q�\���g:e*ܦ� ��E�]��Tp�X�n��˫COZ<p�e���[x_������o�&$r�;;����i�K��p�
S1��`��$�g:����]�r�x �w����T�>}�������&|9�ӑ��\c�L�ĵLi���(��<	8�K��oW��vX��_ow�9j-�;�F8*0Y�X�4�[��,�8>C<�/�mp�ľ�l�����)z�(	�$l�3��~��k9M�ơ�0\G-v��F���9&
�i�M��oa<Yt#�@�<j:	�$\I���'���FxE-uÆC��!�����&����[�;W(:-PW�e,0.?*�C��s���T��Y��1���T��ÌI�ԦP��� ����fV�ԉ��`d�� v�$@f5�?$F�.Vӣu�G�v����$��k���u:+��Tm��C&�u��r�9�%U)3](�� ��=?G:T
����q��7Ӫ�+�1�P{�}+�Ok��V�2d�&�p�o�b�3���wB��p�����z�R�u�!���R��YKm�ώ����ח!//�3�`�x�{ŐܓUB�o�K�l�fx��`�s�&0*�
��ZLf���l1iS��F��0���`�3���U�LԱc���N��!�(�����9�(E��ΣMq��B�Q}@�~�{B�����  �O7H�5C��,������y���pu\�U
����h�޼�m�W��4te�36���ʚЄ��Z l��ts��8��r�����ݦ��9�U�J�mT���1֡-4UMd�&&�׃EtiX�N�o^W����j[�u�f����UK��ٌ�w>	��]�械�)w��V�l4ܡΤ����F���� n��1\�d�9���U�/�t9�ѧL�>�,�u����������e�YE�u�F�ge�p�Jy�o���z��Vd�:Ъb�ؕ9h<����ֲ}
�l(o�;�\��;��JD�ߡk���t��,^�g�;w�!���v��:&R�k����ma	�S�A�|�tW��~7�mq��0is�>����;��WM���������[~��Ʃ	��:��;�Hi0�YS�Sy�E��03YP��{��ڍvF���!�yV�e��]G��C���!1*�n��F�౺�݄�e�5����9���S����v�8���c�Bs�S%Mq #��S���.Ɯ/!���wc���aO`�pmy�_WГ��As�8^Vi��.؃1��e��kL���+w���nT�x�<�Qؼ��ۮ7�|���N�"�����[] ��7y�hv�s�|�2I�.9���6aw��}q[�U敒h��l�ep�sx��A	� �5gI1u��l�w{)Wuf�/NY�j�<�]�+D�������V��5n�Ύ�<:�Q�=�F�-�xڄ�ܛNc�\�%��V ���5�N�F��!��C�&��5�SH��a��zV��Hi�
�ӳFۘ�zvE�!9H�OG^@���8�/T�iv�K ��Ǌ�B<� Q�Q�֢�!�����I�PѐAa<Ǒ�5٘e��m��s�Z��G���U�K����>��$C�u���ի�sV.���.%��T3N����Z�3KE����
�ѡN�l7�Q�u�����嬕����=X�Rv쬷~�L���ְ�x�[���5u�X'�s]F�]�� �sƬ�RT���<ۘ��ƉG ��Lv>�x���N@���j���5!ٌ��
́:�Ξ�+�H[����K��	}��p_���r�8�JP�Tr�e���3�xFf�Uwnp�A�r��v�uwUf�x��TB� ҅��,EFҠ�������*-C�]vz��0wܡo����1������4�lK�C@`��A��27��ꄇ�.�t�a��FY�5d ����3��Q5��`�
X��k[��^5���t�T��c:�ߺj�y}���J��ڕ�n�W����w"7r�k}�
����4�+���G?9Px. 39g��R��cɇw�T�\$�gm��2N��}��|6+�����Ҏ�R���ݿr���j�7�(����`>0�6�"�̑%
����3�ڬ׳��������xr9�f6��3٭�ss�Y;��X�}l��hh��K��)��!��_�j��ȅm\U��{��T��>N@�x�E��i�,]�嶨8���(��l/VMbWW�Ah��7�ޞ�*vٌ�sKG>.c&�#Dl��WMsw.:�ܔEW$wPG"��jbl�^H�Ӟe|�[dAmYd>4��]�Β��iü�l ����omd��̩�Am�#��i�>�|=3��P��[Si��_Z���e�w�S��Jσ���",����'j���s+�����[Ͳ�H��:@C��Bzc�P��!�2Urc����.�Ҽ_��Y+�j�'c�J���N�y���(	,{�=��vS�h�q�'w�!s�9��~��g�9b8#�:eι��!.��`WhEe�p�����0Lw�{7낸�s�p��h?S��nC�s�w3���t�ɼ�]c{ܽ�fDp�
�c�B�Y!�e>����;�u#��)Vs��<�/G+֚�	�7X��I�k]u(^U�'j���<BΝ2yT6�I����2\k�糞�FN$��rC����7��.��U掉���� f��Z��NLX<C8LeDA��'����|'�';e�^��ÙUC���֘����.G �d��p��ŕ:o�`�k��W��n'f�	B� ��o�yw"���n6�k���^*�Ծ3�o�نtX嵆T<O���UΫ�I��@$��,��E�ꖵ�ܮ��36�F�IO7=��p�1���}�M��z���r+_�����$�wj�eu��R_�t�؝�,�����1�&F��n��,�)-)+w��S�������j�mK��0��Z��a�s��١5��8Ԗ_�O�m��C��R�2�F���0�1�@Y��P@�$�&O#7�R?-��z���9c�K]�w��+��m�MOjU9[c���>�P�����d$k����r��U-uÆ|�����|����b�ҡ�Nt����L�g�,0/�Ui���Ҫ[�϶*��.����P�ؼ�ڱ�Ճڧ���5Z��&.5�������$s�D��tex�x2��u؈ՌC�Qku8i���G;�u�dᵙq����T�����Ɂ���s��S�y|W��vie��z�#��ż5��+���̏�լ�e�������[�9|-�m�"����,\ٛ���-�zkP=��
x����">���^l*��#)Y��+�
��Te�*�MCn�XB@jZ��\O��Gx�ۄZ:�%k�8綻�I���� ��*��\v����7	>��5DU�L�7��9��b�ŒEj�����
~:�wrF�^1X�C'��r򘮃�i]WP���ϟO�MG�pY=���n���9��	�z���Ȉ�����#�'��� (�JGR�&/
��6���E��Q�����RJ}K�"^q����9��j2�P��YԪ��iUHl�c�G��ET�Y: �����V�W����/��̫�b�+��ƻ|��7�b�OF����̅WYt}�梱R�pBzn{,�e���-fy멬�q�	� LGc�1\�d����{=��u!�e���h�=h�g �.J����ܕ6��ޝɎ��/�sѿ��
����/���j�<#v�G	�ٹ8u˰ iJ�P�č��%��`�%�%doZ���F�vy�҆y��<}Br�Y�����D���k;@�x�;��w+!b��W<%��i��ɎU�ٕ(�R��k������t�8��[S�=7ytE�p�Ԁ�i�:t�#��bXIʸۺ��{t��	�*)�y�C>Ԗ�!���߰�� ��u�{�5�ʴ"�k�h�5Q >�F��
�с��V�;�U����`X&:�sr*Cs;3����]c�N��J[���=a;��G�q�y�^��K�����ǔ��P�4���U�e[�x�H 1��U���Ҧ`�lq��%j[�\�E吳|�S��؀QJxa�]���}���O�x�5��[T�D82<��_�a���WP��4]X���r��ŇOZ;�ձ9ǰ�ɣ�l�nt������o��f,���Ag:��`�u���i�l���gܒ��sD�w�;�t��A�3���&�6]^���V��i�R��Q��ڂ�8�g�*����kw��N�8
�|*S�����Y�R�4a�TL�o k�f����j��;v;�ەX����z��!w\1`8�%C^��j�Km��A����L�r��S`h�Ä�AT���g��]��A�����H���tOv�I�4�)wVl�V/�"]2�,"Gܴv�����Ġͱ|BN���3�=�sӹ�;մp"�p���=(ҍ���o�Gnb(*H��e�r\L���=��W/�B;u���PZ`��A�4C5����mV�γ�e�ǻ.DyفdzQgnj�e���\6���&�]�i����ĒV��<�����k�?0wR9F�9M��!�0.��b�Cc�Ӵ�7�Ú��U�܍�k�� ��f�L��[K�'��T���i�A�j9��u����ʘ�R��"g��f���ړ炘�h]e��S�s+D��*Y81����ɤ�$����Mw4Y9^�	����e:��5!�#�6,\4���ՍܷP����!�rUȧOf�!�=���7�a&�Z��±�[Ն��Qnl0�N��;:��vw3y��l������\6!y[�h'2�C���+��|6\�;�,2�;����Su�0�n�( �]�I-	L�X�{:���t[���yd@��s3Ύq��If��D_.�;�1V]4����l����̬��pX���3#�M8ټ}�~#��iQQ��ռ�84C��4�L�7�#��+�n.��^*�ԩ	n�8���}�x��N-( H{ӎ�a��t��laO첩�E�W"Ͷ��=+noJ���%��f�woC}�-v{��ժ�ڳN�C"����l��Nݖ��sO{��|q�Uq�J3.C�����朳	��h��\�P���"���f�xK��	�	v����(��b��s:� j��y�cP5�j��+S��ۻ�l����l;M��E�T�ұX���n���Rr[��/.����m���Yէ��RCf�����ڑ���
�^q�u���s�|sH s��B*��\���NV�X�^f�������˨�O�� H�	 ��44�t��M:�B���#d�BS�H�"6�N��4�5HRP��T�&�)J%j���@h�)()t*�����#@Q�
����SK��*4m��&�щ�J��iѶ1�QKU#A�CE4%&�HPh4��SEl�@�ѡ�F�HP�it����ւ�BSIDH��AI@DR� D4���B$�F�"]j�()*�����N�-���J46�E4�#R�T�T%m��
����:��(��C��(�� U$JSH�	T���AAM)�>c��K=�8�^�"vDeZ؝Bb@���+��{���N)�b+Ǆ��"s6���k���#U��1E0Xه�
������c�x�[<���6��|2�~t�O�:�U�䄭J��캉wM�	L,9��!�����{X�3�n�F3\�=p�84�T+�\�j }��*�l̬�j�
v��C_n�?h�ݨ���p��9O����L���5�4�Ik�D�A���a���5�9Ǎ��Ỹ���V�ơo
��t����w6�����2J�O�Σ�ve��W����6k����*:��ѻe3�cR�ry9���sl��X����*���K�'u�i$=^4,���[�C]�T����B�i���Zms�<&LlsN��A\Xv��[��M�r�}�w�!�o�xů���h������x��:��>�g��C�G=�lkDY�6��x���wٛ]ωk�I��U�K,crK�^�Ω_\���]��0�]���ݦ����VX�j�����4��X:X�.5�MҾ ����{]�'8���;ϒ�뱇q�4F��sk��x�m���p��N�G�ޘ"륃�<{�ȾFTݭ��	�X�n9V��8!opi�(i��V&�0�\�皠�˾B����I�<֙$���v�}�����i��y+H��#�䖐�S��{��2�io�S��������kf/����b\/v`���X���"�����ﾪ���nN�i���ͯ���Ɋ��Z�KVy[���#��۳��VY�N��~��8��!�U{^)�V�o;�y�)E����ٸ�?umR�� Ҡ���`+P�r<�;�����Z^���m��	�W��b��q��PF��	�U�!��]��Գᮬ,��� ��<Vڬ�&-=���šވ����{"���[s(�� F��30g����=����r{�r��P�r)5V}��ۧ�<]��/+�Mt�=��!˳�ŇR[�?{%Y{J�����=v��tuuTO@�l���g~�r����M�ꑷ
��@�=] ӐI�<�:��E�13Y\^=��8�ل"����[V7�+j���l��;NBrmC�r2��#8�\P뎁����c�����R��,�TD�U�2�B0!�ioWϕ;l��Z8Z���&�������5��g(�}��Ȩ��)M���F���C��C�K�s��K��!N�y���b�R�ox��54��_W.T��q8�	V�U�i�"��4��+�o_�}R��#�; ��U:���>=�6������Y�پc�}3�lh]X)��diz�3�uF`��/6�����<}�캾)_
�ms���2ü����-�H8#�P��]e�Ɏ���Y���/�ED���j.�=����y�RI����}�D}��Y�u1�28Bɟ�t�W�偞�E@y���ˠP�2���]�� ݞȍ"����zz��Yk=��u��O�������Br���ʱp��T�*��%}X- v�xoTj�#��Y�qWa��tèX����ns�+�1���l?���\���U����e��U��{�*�����\��I�uY���ߧò�������Md~F��
P8{'s~�G���/��z�P�Z�8T���d����Z�c"R�w@����sJPl���%�y������Ec��@H�����q;3����`@n_p�ci��yZ1��Z�UW���T=���n��U�~l8�3��#�h�Y:!V�%Y�������A���d��w]��7$R����1	��c9G��йp�w�d�ˬ�r���k
�=-�S?z�;+�mӹᴻ��χ:zr#O�,�P���1�9Z:��~���]�$+�͚S�'��' p9�u�]R0£��K��9�RY�x~�n�d�xW>A+O�r��κo�=6�CmE�I@뮭+Z�ok1v���zvZ�>�p��d���|��o�9�P�ά�VB���y�`�
oZð'�x��l�i����.cꛗ\�/o����9kvJ�� �����ͻ��}��}�ы��v�yoU�G�GA	����fo�2�����Z̷?��0ZZ�#R8þx绀r���:3�_Z��gG�P��P*J5�@�H��I3�N�Ќ��Z������u��a=���o�I}�.ζ��nbR:�C� ��jS�݀]��u�,����#J��9ڤ�VgT��ա���&,1��Pۭ�㸚.C ��[EH���al8K.+�zu��T\;�G�"9_�>Bb�L2_ͺ�^@t�.�aU)3](��ޑ���e�*uѨV�2'K����ଃA#�o��\o�_�	��*ԦL�M�����3xn�&��J:��;΋$�su:6�S�h��5�~uV�'�������p�'w�2O�Lb���g]^�yt�O��k��������5��b����Vr����֫I���A��A����i�MlE�9��)�U�}�+�ޛ�k4��-ʻZ���?s*��CjZh�4..eH5cn��{� �uC��g�f23�O�n�E�J'tVp�ڣy��z=T�FYp�2��[�9dbQ��\]�ݛ��n�=���q3ask�,��<�t)�����/�'��&L5�zcY@�b����y�+/�)i��z����rV��G@����jh�����kh�H`A��c�^#Ⱦ�S0b0b�o1o�������W�v�!���37�� oݏ�H�s�C������p����W��b��Xȶƾ���审��{��G���aʯp!�
��Mr�e���������ۇQ�l&eTm�y�eo���O�I�'C�3��m�:����	1P�����`�ŀ��q	�e��\�e�f���ٮ�[6���4��8(�o��%�\����veJ7�)��;c��7D�ѮO`Z�&^:0 8�m\>�8���&9rK!=%��͜Hn�s��dlW�Q4�C�r��3ubC��ၬ��(�rid��©@��!-T|;�N봑r��R��y��c{Է��F���}£뉷N���w�N��m��Pꐚ�L�5@�H�5/��}{\��ak����m P=�b�"7�|��}P���|\��AyX�n���3T��/<ʺ4�a(�n-�o����& 1#�+�W�:S7x�K��L�aAsl��@�QTch*�����=��$V�QJ��v˕x �hO���[������̀���ؼ��Ǭ!N���w2�q���sv@�X~2������M�.hѱGz�"r{Qݜ~MÝ�K��bg#
����lm�S��S���C�X��1ޝ�.Qqf�C�JN��DS1I��Z;q�VoRH$�3D55 ��=N���UUU�<�'ec��񅡣�_0/$P&���ée�O�t��&,fR���f�y��s1�V�+i��ߐz��E��k��&��V�����j�WJ��{d�@6���L�8��%52#���cE�ʹbҪb/它/�Π8]x�搫L��qv�U�- ���C�E?���q�0F����}l@��Cu�F᫨��u�{�\�fmfM���w��b��.�X(�&��΍Ȋ��Z�KQ�evH���*��j�ڕ�jF���<ۍ�Ӎu�������?|�PK�u���|ǹa�`+�mC\��`��E;��%󞓃F�W��(�.���E)*� G�
`Δ.Ib*6�V@�V΅Jw,�:)on��_*̿�w��L�u;������v�\d4`��aZ�cK_�X+�����ؤ��E�|���uʇ7z1�C/ �������D���*���/.Xd�8��(��OM=9f)º�{!u�K6)��JU<9�C1����9�l��ݿX�"�oʞ�Z��/[B�����Gs\U�zn���.��Z)��φ�eO�-��Wfd��o�f#�U# l���9���S%q��z}�s���ŐXG�2����9�i,�X��Z]wM:�3GNe떺 ��ccL{uz�B�p�Tw��������̋�O)��@s�<�1�4BEt-��![Wpe�≆;' G<u"ᮮ�wx͵�B��y�8ofY�$:E�Ҩ��J��S(F7�ޞʝ� ���O�Sn)�#��T���]h�{1ҹ���\��P��?�"#��u��7>
Xwx}�C���A�9o��;��bѡ���r	�d�f��T�&����	V�U�i�8<��i��Ꝏ3�A�Oz����P�ϮB�g����K�X��",	�����B��.U��n��i*=�j��1�Nu�p�a���ۄ"�s�c!5W' 0�@aNʱa��qd�`	r]�.V�ư��.��?ok`��ps���6�wx�O0<�����MC4�7W�\�/��9N��)��$ܱ�2~u7Le���x���n3�_�vcy:�U3tY����TL7�������of&ڬf�F,P�HT4���u���T���*���$��{m�2GU�i���BmN����GVq��yS���=<-���/��g��7�w��"�C�Њ^Ĵnvo�
��J�9;��4P���p���ќl�vB����ס�B[��JdVv㝽BMui�����S�oeY�h;%�����s7���j�Q�9,����Z�Iu�����a���$��p䑼�8���<Yݘ���/��&�k�0̤��+]><��꥾�vb��ڐ%j]���&~'D%8((����b�V�o�^��$���5dwb#�:"��s�)��u\cs�ܴ~9� u3�x��=9�L����=XĢ�µG�vdm��V>a]��F��1�9Z:��aB��۱{y����d��-$]����q�6f5�Bir�ŢYz\F��ޣ���$!���]u��@�z������(���}�R?-��{�n�,��Ʈ�1Z�Z����
��v��mUr�.9�ү%����\+�h�{D�Ḡ�v%��n�d��V�Lc����3�Xm_�g\C��3���o��t�	g�F3@J�κ���	��DMf:Zܽ븵/[5����BMZ]"b�5��.;�����X#iu"��s�}n��T9��C������)��1O����P�m��t�-�'�T��ɵp�ҵ7�^j�:���Ҁ��;ga���7Ҹ��>��5PE}jS&Jn@׶ƒ3Fu�5jW�%J���~~��#¯=g�Xq(��[#l�UҮ���������&á���]��gh��3�]��R�7�I�������r�,��Y�dnnR�����q�mu�<��ݚ���x�~gΛ�E#�*�Bz�N����ܵ��pw��ꪯ�W%�jWz��W���p����1aI�?g�Km��:��]yp�d�J�d���Z����rT�<�x<���,�Py@�w2�WCyJ���P��c4�����*���{Ƥ�Yсƺ}���a>��\Б���D���~���Jj���}��J�ohY뛼�	\F����uXR��N�����������ܲfp���q���z�V�d�J9C�Wq��J��	|Ol��˧�Z�� }�/<5=�.�C����`���$e���qt2�1j��<�Xj��u��7�u�CDiaw���S̾ߞ_�uÞ�¦`I�l��EVLXof����hD����9�i�g���`�/ln��Y7{i�l��p��5_\���v�ج��=�W=%���6g���̩FQ�]O@Ķ�;���iS�X�kr�|�*C3��gi�p� �r�#��,������̏ccum���gnvq{�<�0����_`�7�%q��F�1��J�X�(�ρ�'�B�X�V�W�h�t @)d�z�>{�"�>��z͋�fY��Iuk��	b6y�z+���kw�<ȥ{0R������LR���W
�M-筨6ۜbH����m�v����1��b��]'8���R<;�\ٷ	��Z��IЫ��0���W�_}��c���,v-'�9�̆k��\Mçq���>;��!���f�uHMB�*N�����"��{/�s� I�8|`���L�/w�"7�B��BN�8\�����6�@��e��u|�+kVܨ�mP�m,�*j��$w,"FC�Vlb�,o�S���p���ھ�E�������8٬�͹�@�	�|:�W˕x ���f����G���Em��
Ȕ�ӳ�޼�ѯf�fWyUg�Q�}I��,�~� �� ���lu�N�(a٦��UhǸ\<1Bޫ��_ܝ�
g�������wRF�'�.�;��İ�f��EL��]�����p�X����2�X�J���Z�3K>u��~;�J��Y�b��B꽎�5��uu��cX�)��m�����f�n�h�WQ;q�/F�sOؽ����f���t�#}�ϊ�!.����R��%���]�:�6#9rU��Y�_��t��_��s��$�^�����V.�y7*��l%��o�࿋�=���_�6��������Gml[���w����?qa���v{��Q�;��gq���_S'+:Xo7�j�l��x�Ez�=wؖ¨g,�/�|_Nf�
X�s�L���m��36!&ЏY�U�`.���W�,��J�yK))���8\A��oqoH��Ηu�5��n#W�����7���n�Ve�.�Z��H�Z9k^��Q9�1�e�|%��7k�6�qt�+G��P�v.�u���� �NQ��h�X�\�zě�:�E��Sh�f��-��wE�6�)�3v�RAM9�����D���gN�q$�Z�\��N;9�+dr�P�x=޽��������j�>���#T"71���:u�#��.��we���)��B�M�r[%'��a�����E�ڰ�|/�j�A{�x����R�qo0W<�x6�����Yý��T�V�j`��7��sp?+Y7��3�!���1B\Q��\3B�I�}=<ۣ#m��f��ŌTk*��3v��O��%�<(^�2�ӫ#r�s�7�.nwZ�#WOk����٩�%��m��G����7;[xz��]{Kw�5� j�"V���0���6�`��������Ei�>5&�l:�;�a�ב� ���RF��[6����zc0A�[EY6����Ά����9�՗X5U�K@Ȉ���m�N�`���7��\�*غS�����'cl�:4_�4;V�Gz�9�s>�2_b�M>�B_LJ��[��m^+�|�K����Q~x]���zP��oI�~�rͅ��EmXt��b��%��E!�:d7|&�hl�՗����5���5k��%;4�W�|{n���hs���g�l�\)�	�{���Q����)�v��
�Jiun��b������?�-�Jp��gj��]��ᓣz�+1��K��8K�y`�C�}<�����Q4ē��<N^�x8{ta��!�ܪ<P+�j ��^l9�T�0g�/g[��č���R�BD	�z�h�E���h����N���ob���_sN08z3f�~���s5��|��Qv�������ڋ�fO.�WEYF��. M<s%��tM�C�[%:*|*]j�w��,��n]�V"Ҕ��������YW�kV������	��I�sq�1a���lv�&L6&am���Mbn	�7�Hfi��G$��µBr�_l��1KV��r����M���R����w^�� �V�/K�a'�a������i����{��ܦi��֞{TA�uw�&�Xϫ��wx��"�5���øI�X�qc������n|��GI;j��\��K�K��&�s =��o���G0�xU�X\j�әu;#�3E��>�Nz+�Y7ށLʍ�ź�vÙ�7��-��N���:��z85bPY���g,���A��m�-��I�{��8ֈ�2��6${F(����VC[�ؼ]Ś����~7�߿�w���}����V�)B�G@i+N�&f�����(��i
R��J(��R�hJB���)@���@��ZV���hh��hh��������MP!KT�@��	HQH%%i�+@4U4-UAH��B�R!T�M!H4�SH�URJPҔЅ�4�SHD�@�HP%P�!A2UP%-Dɡ�5@�4TB��RSJ�5J��_�tǎ��ݺ���0G=Zm^�/x_pc0ǌ>B�L��t�*��d��)��"v��E�Yދ8k�q��;��W�}��'��({M�C�*���.��!b��J�;!=3 �kHiq�A8�j�39�3���O���C��p鈸NS=��>�7�*!vT�qf ��?&f �R#-mv(��ʣx�i��$ۭ��?c���,�sw��0��t�n�zn&�G\�Ƹ�J�W"[B�M��Y��v�S�C��aW�颱u�K6)��_)T����3x���{�#mU|��}�5����9�bl �N:@���!�b.4�E-�ǡ[WfY�(�c��М���y�8�����v:W<6����N� E-�4�̄����L��Qz�r�M�.���I���1;��E�]�i��r��L`��i�W+����#ܡk�P�A�L]l�Ln}Kp�&w\;m�/WV�o+����pHO%�_�{c`<Z��lgO��+p;��ZU.��G5�	�X������W��b��~��*d��9`k�"��N�����,.�<95Ǝ�f5=܈�He���.6�8l��1�����qX�NX^@YV,;?y\���3� ";/#��T\���nu��Z�р*e�����)�,�Kx�:�,ʺ(S�:r���䳅��# Jn!dW��[��;�����K#X����ۉZ1)��ls�l��vM��)����FA�Fʜ<{Fe�6L�bff��'1�=����ﾪ���(��i�K~z�G�9;"2.���]����6!_'w�!s�)���m>ɾ�u���[�+�"z{���ٜ�8
(o�p9�*�	��T����vW����\u�� ����q
���9�����V�P��@��
�4�Gk�B���G����^�������y^�����8�p�c��{"��Y�1�Ν�2��!0!�B��kc��˱ա�{�J��01�@�u���I���Rg�������k���}���c��Fy�5�	.�ٽ�J&�W�QΨ}�1�!���ܯ[�oG�](�U�U�n�7�qfvj���j��Ib�5��'���vc��v1+�Y�=9~ae�LQ��o����vv�	�V$M��:��;�&�i�IƖ��k����5�u�Qf�f��.V���Ԗ_#�)q�G��/�ozʛ/���cƮ�i�q �X�'�:HŜ��OuzF�E���9[*R^ٽo�s�^/bV�o�F��Y�������Ƒ��j���t"����l	�������Q4銝X�#��m��;3�������h"2mwV��t�+I�G<Xx�nx������N�������^�F�^�i�y��$rġ��D
����rw����`�a�z�!�W�����L�V���:3%m^S����)�%���te��tj�^���"�Ă}{�������KU�6X܄븛�븝7%���q��XM:�4d^b�s�v�ј�-���Lb��pF����1ˤLXc%�8���M,�i��\�{��U�6�D�ϖQ�B�����{���z}���Te�d��k��8\#q��r9��Y��W;˙�-Γ�5�=?L�����v��ZW=��j��E2d�u�����>�(�O7��]�����1���W�;��s�(+;iu]B�݇{h�Mtު�s|镝�H�N~RjJ�����؎0E�誯)_h� �~�{X`��-�/�15������a��O�1s��,}_un�ڳ>���J���n�r��d(W�u��YK�t�T�xn�5Kŀ*��1aK�Fs�뙋�����ܟ�/ѡ%V�'2�6_}�������cp��}Ss(̾'�H@���w��%������p���t2�쥯A�ݳoO���W�p��hXyQC��0�W���
����/����d|t:͋���@����U��;�Z�!s���JQv|{����^A�}���9��,�>�2�R[�]��TuZ��tU�|czV��:b�mz�D�*�P��}X��,D	;�a��n�%��y�R�U��8����ӕ�9��1%3gf���</fz�Lb����go2R[�\���*�
�(����$�:PKO�7�_ �j�_+�:5X��w��Tε�I6��_>�:z}r�Zx���#Z*�>�\7���ݵ��?k;vsi�;x5ǜ�D��wm��(X`#�uB��u��`�/$��&J���ۘ����`4�u�F���bޚ"��Ÿj�}ʰ_�����}]�m�@^r���Y֭򡇕�(�,�/�sԟ\K�Q���9O%��#)�!1J���*s5{r�v�z[P�Q&�~8|�*�n#L�/v$��5���I�D3�(����z�I!��=�������t��:!?[if)���H�;��#!�-S.�1�	u�2v�"�UF4���Խy+X^���rH:�����׃�8���7�mF�.�ge�W)����Y���␞N���4�Ѷ�#Z����\Q=P6~��\J�[��\6�����&�j��SmF������
g�������7�����/�?r��˝1�� Q�k0X�.�;{G�.���U�=s|�N�7��d��E#�U~����7�����l=3��D���>��DÚ��& =�����Bî�%��د ��d|ha��n�w�]���8��_�����}{ɖS��i�������7��2�X���b-k��,u��bDƻ�s\�հ�[���� ���@~�v,�D`��l�sk��v�\7_4Z��̨�ѷbR�W�%TV]bL����0E��R�%��s����aCϒ�mc+�a�*�e�.p�p7�@���8���V{��+T��3V.��ٸ�t�^7�:0Ҡ���`+����l�"s�T�#�c�\U��Y^Q�]��b`�U�C�(\��X�Q"�u1Jq�I�Uk�U�����a`�_j���r��{)9�#r��@�l/o+1�8�%�`� ���6�q˻�:��v~u��v!gÛ���-F:�=7s������V�{Ŭk�
�`�����c�#n�+]ĳp)��Q
U<9�9��:�{�#k�7�6�<[J�ٟ����v�@	�}%0��+�Ս�
ڸ�Y�=
f�7gq��J�<��^���#\=ۑ�����L�"zӧȉK��0��[���V�n*J���>�qѿ�K�*�7��C�������6Sj�)]��]�����;�0���5�����fstG!�'hK�-owZ�������кݤ�c�%*��ң[�>yY�h�y0޻��Z�(�p�}|hҐ��ܒE�舏��I�s�ܧ{��c�N"��.c?���s����#ܡk�D����֪ߦ�r�|��{o9]�V!��<>ƺ�AՖr	�d�'��T�&�Q/~�ʞ5y��y���H(�˸��¤�w:�J�A�ꐄ-��{����^}DE������O�H>k�+q���U
�ନ���t�C'�v���=�15W&� 0�`ap�hvʃ��zi�3����ڝ�iw�g��͒��l*��{[GA�:vS���7\j9;�9�������d�ːMn+�+ʹ>>�H�<#�F�uԼ���}�笪�z��ٵLq�d���q5���Puf��֢���ܛ¢T���HT!��*;^�P� �\���ڦUr�'m�*�ؼ�U��+�)W��]�7"���+~^[��Wih����THu7'�Fˮ�Ș�vk8�]@h���=���������b��t���c���j]ו�GM�Fu�{� !�R�I������}@�䊵<����#�W7"n�'���ָ�b��"���r���N'3~��9�8.2���Nht�p��y�>i�����rC��7�h�If����������R�;MHT6�|s�����=��$��.l2o/����������P^s��#,�i_5���ږ/���gn�d��/"����KT��U�N�2j4��J�s��F��Yt�k�(4�;� K��Z׫�W1��Ӝ��d��@����L,��F�W0Y�١5��'k��ܾq����d��&6�mb�T}��Od�2�[%IX�`D�ii,y������n"�e*�\�~du;�[�w����,6��K9Y+����i�9��E�HSh�&��b�]]pL�θFxE|�����͖7��n���p%��
z
��L:
�g��V��w�-J�圎�\sa&�������o"�v��e�����U�w8�	<�r8\�k��]�{ɾB��\�o���q���J�R�9���6K�6`��-�gg�9��<���H!9��ߜ��5�P��[���Dg!���g�ٕ����jؚͼF���Z}��*h���Z����sP�A��s]��c��g�3}/.�W]�ǃ{K���7��{H���i.�V�8|���:w�q�=9�*�m	j-�4����P�m[�>�nQ�d��X�l}�U�Z�;t_W���L��W+�;�7�I.8��93��р맠>�`w'�.������2F�H�	�8x����G��R�x��)��^�=�/n�������uu��'�7l�Q��
�N�{��8��9�X��r��|�
�����V�n��1OC=mzӪy^�tj�u�~�}
�܇�Q79BSxTv.g�T�����q��ۓ]<�%mb�yu�h��z�i��m(j5�ፊ��놆a�a{wK�8=�E��[>0�	V���<�U�Թ��R�JF�NlQsqP�^b�۽����4��t������Uu�������T@���݃�G�k|�s�F�s{o�Y�7����C���GCG6t<w50�m�x2�y�����oMB���ֻ#�q�_<㔥*�PP��^�.���O�'hi��	B��p�),�w��N_u���=��Ź�r�]#p�z��;ճ0�ڎ?g�Y҂գB�hf�[�ji\���"�si���x�ez{�4m�xI	9���B�.m��Y�X�2]�\�0Խ��Ξ���}3/䒭@fܗb�M���*������_��ä%{7aבy��^�w4%����0gjslC<`�I�=���M8�ݢUw]ߪ���:�㸸p�C/��U)D.��JU��J}5Իw'_=ᔮየ����;�L�I�\����k��ω_oT���=�N�����2���[��u�R�ϊ�����b[q��J�"%oBv:���(+^�*� �伞ӫ��c�M��Fk��UZ�IԬp�5�eTk�'�c����ꗪv�T�֞���Z�7���[�J_\-q��^d?h�|��/N�ͭhL���p-:�c6�e`ʎ��#r��R��m���ʜ
�Z���a�+і��et�s�]ǱdM�W�{ï�'���z_�U_Mj):��=ԆNv��]�׳��6������u��%P]^��$���վ@Of�7�5jA���U۷fQd-޿Mr��'�?P��Bsp{Z�Au����5X�J�cb�����{>��d��_nC�����[�v��,	ɞ��ji���K�Jl� ��:�:#xk2鳔xl�&�+V��݁�S�B|�j�Z��ʗ�5�����W�u9�4��3r�\l:�n]`�QmŸP9��in ���>�k36�����ե�J��)�Gk��>�彩��޽2�3��uT*��ꢶ%*W9�����������V�ә}��ľ/;��$�k A�@�uR��t]:{4�<��n8x�Q�2��b
ԬՔ����N!��A����+�В_-��O��s�7[�{L�|��~��wb^}Jyxr��!w������Bj�-�휪��!�3O�s��K畗�O%��wa��2�"P���Ϧ$���W���\�X�lZ��T��R\��o��L.f�U#?qGht�/�yb��N*n�P秥�{��d�su�u�}S\���;�n&�:�t:�ݼ�� ' �T@ۘ=������s�q	�5�Zp�D&�^���0y��`c�Ȏ����7�.Q��y%���������g6�vb��Z��Ǯ��YU���-u�_M��Z3c55�������hȮ�|�h��۶�h���V�I�.�V�މ²�V��V�l���8�����M�x=l�%:��@y�����\#|���$c
v�j�G`]d0U�2�H���.����t.x=b����
�X���^�ʉ�@�&�Q)��=�{�J.�*���YӮ]Um�Io`0o��H���Ѷ�H7����yNl���M�s�p`fѺ�M=�Nl��c��n%ws˕/[���2���
�'Ǚb4�:����:�^��/�Ȭ���w��*��"��\Q�7��w^u��1G	qf��*�]pJ���2�[���j��9*��kQW���\ON��1KK��s+�niv���[=�e0�/��kv�G���" �R�^���������[�׃�
��qW���o��nhӗWY��u(^��!\�'@I6$��l�N����ñq�3�o�_C�/0�ڄ�@�2����$z���g�����nE����9��K}-�G�Ru�쒁�HI�KJ�I-Ҷ�\ǫ��rp���J�q�}w����/��z�^���;XуsM���6�m��}���t�|�k��Ź�{6�|T�Z(��Ůp���.��X?
�G���w:�σ=�w�,�p�m�Βa����1�����V܄o��Y��hͭ���i��S�4���}��s7qj=︜[�bb�#��]\����V��ved��O+,	M�M�kp�\�ENR�-:

_�L�nvg��_N�rx9��^��ݒ�<�8=�k
8y���^��"�R@BP����]\��=�`6[����\���;u'=�5;������[����[���?^�Ҷ�Q��f��Y��ռ1�҈��QK]�!��v�Ù��-�X�ӗL�F�Z����I9�P�%(W$c8�����1��nI�J\���'��0\3�n+�bլ,	PW����o���w��+�Z�G����R������M�ɸF����{PS�������8����H�:\���s[�6�3���/b�ܪ��6�yK<#ruO���V��W���\����/x�y���ݧ�"��E�@Vc��������BZ6Z�R�]�'�3�zZ媰���V:��.�V�<�� ��o\�h}u�7�h�'��f�{ֻ7�Y��_j�������)�����iU�J�_M&C�`Ԋ"H��PA�����*�1�Е�!�9�6AM����7�WQ�Pz��8�:s��m��^��eTV5a�s��S2��[3��-��Ӕ{�����n�L͡�hhz�ζ
���	�b���P��35BYGHɯP����w�2��U�+�Q�;^���[��b���=��߬`�� >�h��[jќ��+�w+�,a�,��	�}���-z�j���e6�v`�*�r�lށ�`[�T�؛'���nN��.iz�N���t@� )
hbR�Z ���R�����������(B��( ��(����J�*��((i�hh)Z��(J"/��R��DP�T�ERRSQSM	IZ����ER5E4�CTUPPRP4�KIH҄HSKE4�%5H5@UICKQ@S�4QEL��E�PPE5T�PUHUJ�UQKC2�DD��!@D���4R�QJQ@D�QE5KIE ևE@44Q�҅RR���RPKA@U	BU Uu���|�����Ys�^H����h��q
���f���|r�efMua;/�Y�)C`�#�f�Yy�>!ml�N�}_}���킣T/�aW��n5���v���tj�P�	��4l�T�qIrSƊ9�۾�u�7wa�>w
g�����n����|Bڝim6�(��5�^���g��J�;��T���j6ֲ�sb�'�{3U����M����֫iC���N61���\��_muNʄ��V1�k�����s�%�w`9����C�!{y��ۇ�\�4%���g6�X�+���8j�#�:���'=�%��'/c�2�܀�*��ڔ�B�.�[�t�5���ش��y�e&�E�~>�����>���.Oc��ֺ��d����7V��q�Ɣ��KZ�q�m�؇)D��wwň!��r��r�Oq�,nXl��ϙިZ���-+5�B{���9P�����`,���u�����	[�_m>{�#��I�p����)��K��˺�Ϯ2����Z��mwtٰ�vC��d[�ir�;���,\0зj��/!P�m[�:�ڢ�/& gIPl'�ᵣ�mTS�z�:�~⭞��c�SZڊwm�v�Z��n���c"�x��uxc`S��Kf�)�n\w��>�9�Τ�&�	�3g+�uF���}Իf��M��G.e�����] l�����3ُw���3q.�<���uY[�W\�w�t.z��tȷ�g:��S��s��;���MƸU9쉏��ka�����Z�oL֩�/�7�d�5mu_\ru��Úx��'�Q�ޱ�-u|3���lU�h�.���w�9]��bq��QoO�N�3_s�Ow�̩�
�$�ˎ9ϲ�V]-�zs7���k�_Dn�J���:���E<\ڭݭ��r�b{#iBl�:�g_͌�.��ܪ&�+�)��*'�s6�6-�=ouu"T\�)��o0�Os2��+s�휔�r�m:����{���Z���1B���߈D,*C6&8���os�{cf�az�뷔'��{�ͧ�C�ý�gYtO�3�z.�������M>��'��{l�Rf
��U���.Ct��L�	(j=�F�̜���,��M�T��`�8�ɤ��ث�aV����YQȈ��r:]�T�,�+���#Ac��˳�3Gpb�=��|m�M�'�f?Ir��2�����Cbs+ν����؞\�5J�
&�*v�M���DG�]��p���s�vv�:4���|��i��͵:��ʤ�>Iof����|^S΂��;�E��K�oMB���k�5�uD<㈥,Q���HL�y�X"�wا��kE����Gz�1>4��_�>�����&�*��^��@�������0`����y��R�I4�7O	��/:�js6�3�v�1�Y��y�����
}5K�prl�d"��SǰOs걏�Q�M�v����H	�Չ�hs�o�}���N7`�<$a���>�L�o�k�bjq�FF�!Uo_	�L��L�|��^��=o�XY��o5n�����X�OBn�YU��Y10��f�^�s������Qٕu=}��w&�E�Z�ʸ{j�)���/j�s�T��v��Qj{�Ҧ>|2`ZT3D��+\v�[���z�碯��K%)�Xw�m+�R�����6t�������M·С���/�P�^����x����s�$���S����ȅOVй�/�<��OG�{nE񻽩���ê×4Έu��`�\J�ى�"����2s���a�M}c3o�PK�����p��Z�>����Gj?^O$n������Q79P'�:�b��8ڀn�,�7�U�O��F�Toq�̦Ü{К��݋vr��̢�`��u�۾0�3��E��U:&;�6lr��t��ʻv�_L^��W��7I�W�g��R-���)<)znzzz�s�mj�M>��\��l�m�H�i�͹޴�U\�:�@�t�/�jz]��U)R��7�CYx��6��ZaǍ���㝅E7��.9w�C��mJK�n^��)O/�5�]5r���q/�uXR3�mGcz�R��G\wϤ��b����wB��Yږ�lٝ��]{8�s-�Kq8Χ��(�w�����������V�;�w<������d����$�����Z�0Sl�9fa���@�W��Ͷ^o5ʫ�ˇZ�s�ۨ{�*桾l&*2!R3�Ͼ- I��y��d#�dy�mq�:嶹c�V�j��6� ��ݞ�+0g���w��o��x%�՟aA`�R-��'��c���>^��V��o+�:��tK6�\�F��#��=�gu∳}���)��'B��Z]
=�q3ܷo)�	���PJ���S{�A��Գ_���ux��QO�n;��h�o�y&�7Ш�LLܫ�j�Υ�e�s��7�g�{c�����+����\��&��pȂ�×u��qQ�K�,����G�~;�^�_t��G`�=T����9�Zyc��cC]	�>�X�ef��'
z���o+����:E����"m�u-_|����^2��q�Svh��s���Υ�WM~EeN ��Khp������sz�_v.��v͌��ތ���+>S<��Z��:�4�>Д�I^�Z�.�
˯����^A�ڛ��;�b���s7+����v�½��yn%�N�j�m8V�m�tƺ�� ��u5J��X�Ůo�����pᵝ�y٪VV���Jam����d���'e��PU%*�cY��OEI��:.���@_^������Y�(t�B��ݩI�-��3��0,oK������1�e�U
�m
t���6a����z,n�M������(>=e�}��zQ%Rh���Û=�^1�����}���I{@[�bw'.��]|�	R�{�;wun�g+Ou�f,L���E�]�%����6<^�+VGF�Ü�I���>mㇵ�m���P��;��W�̅<��}a��U�	Ub�8�V�ħơ�쿡-k�\gU�2��P(.���H�<S�n�:u*��ծ�s��_,C9c�nZVk܄�E|񜨇,�P�5��7,��"��v`p0Z��\�Ջ�$��2�;���\Ӻ�؞��?���s:j=��F�z�*����k�v��'P��\��j꼾���u�Ơ��ь>���D�!��Q���b���+���[��7��bKo8z��֓�q�º�Dgܮe�{~=�dI����>�.� �a�.��
3�ޭ��j�'[-p�x��|�Uo�:�r�M�	!��������.{�$����eGSѷ���[��/V�����ÙS���cH�w�ݬ����s�B�`f:����fr��|���)��Vc�dOrϽOb-��,:+6���k�ܸ,%���x��M �w(J憄�7g�גa�X3����g�Z�M]2[|3�����:.n-����$�=���x}w��Q����΅P��t��a:�;$�{�7�Aǫw++�
pJ�����nJ�vN,����6�]�sr������
���s7
�b����p(y�Y����O����^Qd-����8�7����P��p���4pm��$N�e6���yɽ�i���ۇ}7�r��'�����{ �ua�V躾���2�~O�̞q[�O��I����H�+�bv�3�8�a�;�ޭ9t�K���.����o;�|��i����T(t�o�sJ��O.y-i��<?�A�k�_iI_�h�ޝ�R�\CZ�dk��,�����d~@7|}��z�nd������Ti�ެO�C��ac�35�s��Q��..ZqS��0ޔ_ȅ�%�-+�d#�P���h+@NƼUx�v�u+�̍��v6�)�3�]BR�}7K�x��Z�`br�o3���,p��k�M�h;a�7
�3�l���(֋s9(�GB&�9<=j��]�sU���Y�����#,F�[�e{B�K�#�Ct�2s�:=��DJ[ǲ�e�GT��V�jj�mŗ�N�r�{ǵ������ۆ�R�]ԛ�����\t���,=U�s�	���s����(����߾�D�nڮ�}�ٸַS/�Ꚏi���k��+��tD�!��6n�n_fj�x�ĝaO?�;��e�S[7�kUZ��u5)������D�A3��#}/�	⸋�Z���.��s�y��i��/��s���^���#a�����w!���Wd1�_	��]�S���5�����ǜv��}�o�3�W4̜>Ԯ���3���1�P]�b������u5uƈsF�b�=k�d8[��y��־�Mw\u�Ż9\�es��=H��r<5��������_�?�c�����͇)��J�~���H>��R��E�ۻY��3�������%�5ұ�����i���w�+�u�ս� ��qX� U�=.��)J�����5������v:s�.a�q��i��f��B���Wϖ�I(WE�:{4�<L �u�g־�ͮ�љS!+�"�P3���s���l�����Jް^:ٝP#���p�j��|v\��R�N��vn�I*5VP+,�^�	,3�Q�6o��1�	�;ʇ�I==s��
{,�#�F.@һ)�ݸ���IyL��;���*���ˊ�����W��j^]�m�1GmD<㔥*;�}�$�}�$�s�T��A�z��Ux��h��=�sw.��q��q�O�r�\w��X%-��3=�d��}M��+�����g���6�<�P�9P�D.��ȕy��f�[tD!ջ6��E���;jk��l&�h��5a���W�J�a��C�<b�s���hZ�`���+Tܮ���N�Z.����I�Ż	�ݰ���o0����Ș�6`��[�y]��t���v�z	��ާ��f��eL\�����oXwZ�cxZڈ}Q�o�y�*s���]=�#n�Q7���H�5b����i����Y�Cz�����鷂+����s��v�9�#�g�D/.98ֱ����F�P̨��7م��c0�ۧ;Yc8l7�W9���e�v�������61־�N�v�bݜ�dV�6����fU�G��T�>������}Cs%;�ym�w���M�|1/]ۤ^������>���|e;4��X��\�b)9_���0!�WN���"�Q����Gn�4�V�Ӫ�>�RSҳI����ﰸV��;ڄ�_�Ò���׾#nu��zhߢ�}cLv.d�l9�;�X\��p]ڼرO+������~*�ڹ~��ʋX�1c��o<>��%�2�Z>=3�����ꥳ�������s�<��r6�X�&*�N��_�ڸy4����W�����.o׷2�u�ς��I�me�n'�u�%��o5���=�is{>n8y�o��ƒ��C�;��Cհ�mC뫦�,�Uΰ]Qpξ����%�4��_�k]��3��NR�A>2�u���ϧb�wy���Q�U���d#������y�S���r���p��<�ܕ	�a�.eO�e�s�{��B:�q�I�q�9�@�](G&2���,�����Ȩ�E{ ��k���s���k��d
��Ma��u�`�학�_w0� 7��'�(��5�c`�q�z�d(����`�j�碹leu}�,����,Z�0������gBQ�:v��d���J�ے�%����{��uRǼs��.. {U̳�I�uT�3�]��Q})�� ���Rܾ�]��V@o��Q�a�'F�\�L;/�ƾO�t��s�[ݷږ\K-2O
}z�ŏ�n�ՠ��fe��+���j6���e�����zk�Q+ec���Y��%q�1a�[���=	䓇j�Kxe�^��X*���|�u�^�h��eo�Z�nl�*����Y�_ �h��wa�e RQª\'�s�m�|壴��*��B.Rt���wZ<L��o��kص�Q�����������i]B
E��r�|m��v��uXgЃ��໥�*����� TN��A1ץ�	X���Vq֕\���7n�
B<�;��H�&
�V�'I������ܦ��/Xi*b�YN-s(���|
N���@�nQ�fofS���P��K�E�H=�n��������3��tc��=�<�o_.E|jT����f�w*�������+�c9X�Uۭ��8�ˡ���|�CL&�F 6������se;�!��R�IT�����*�&�[�Z����bw �&5<�cHN����h���etq�Cwn����Σ`ӷw�����"i�s��gOJZ����n�U�ܔ溹|]019�Ln�Ov���61���^<|Dl��u��w ��v�ŗ`�})�5�_r�H�z��38ݑ:��Ʊ�� �B�A]R��v�LO���1�׳��S�M�x�o�`ј"�ʜ���U�i�).;@,�v"M ��o�cH6&�:��]]��ʧcw�@��8�hS���i�>�0]�|��^��+�`8�;�ƅ�����2ѳ|�����[�,�^cy�D�R���6q�}4��_Y�fˠ�;##x���>n�q�]��	�ar�]��0��Ӣ�Z�gB�����#�ڱ�q�g���{W�����ؼ��@�f����L��#iK�ww1ea�c��՝���ɮ���6��9���υ�DvU�vf�R�M�ݽ�	ʙt`�ؘ9�3��n&2cI��r�ȧ��"�H�s��;X���u�BN��W��k���Y��$�}��M��w�WS��7�'�oc�s�b��8Bx�6�_|{�i��0[��	�[�}Ş�V��d7.�6�n����X���qy�B�U_-`��w*Z�br;���f��^ �_�Vj�A�Y���բm�]֨�z	ٲ��5�3Z>��x���v�e����-{,Vw��K��+𥍁8Nْ�R��qt�8�a�Msr��M�[5](�������� m �������V\��s̎ն����g�	���zmZͥ�˞�>��b<����߹�uDKT�Alh
��i
@�J���(b�)h
h��������)�iR��JV�"P�JC�h��
��(��h�(t��(Z������h����("h)B�H��i
��E�@�h)h�
(�T�(�i�i�B�Eк*�)
9#����JB�����4��B �(�bӈW�U_<�2�.=���<-H�����"yb�D�4|p��a\�+�E�Z`�t��D����J5���n�/�ۇ��i�FL'5�c�{�W^��^�|}�Qi0i7��\��dWgDkFov%q��"�ݕ�Q�9X��jo5�.�V�����r�Ä́�#]���;x�׆��_j�$u~,p�~���k"[S|�O��^��g����{�zhz�m�K� �9���Eg)�g\<�<�f:�&��	X2�3�LEc�/O
۱��٣]ТM)��0���-�����8��;�
YQt�{����帗���\�զ�u�-{��!��Ő����hqϪÛ��l�҆�uBY1{mr��Fr5��+�?5^=�sѳ�2�!n���=�a�Ss:����^N�n5nYR���-t� kb��yq	���=��g��������95M��S�����Nξ�(�'>\����c�����%:�7x5��87 F0�m�6H��%��+w_�躖��B���ֻ#\g,��,üy��VL����g2�G`{.�Z��o:d��EZ�;zJ����.�VU̒g�T�)g�A��^�Y]k^E������=(C�����37��N��U�Ꮑa�2܆<,��\P���F��ӷtsG8�c["0];�Pe��e���"����J�M8r�$.�wD�Z/O5��7�ރk��3||��ھ���f.�]��V觌�C�g�B��
Z+OO%\�.*���B��<}A�-V��wC�mD�*y���JUA)��!	Ȫ���뵚���I=�z�3I�0ШJ��66�]i0�Q5V�T��z��SWK�w�tje�}SQ�15�͸�a\N� �.�#;�_:�5�2�7� ���ﭜ�"F���
|��i��fN^����-�mC�����KӅŉ]��ohfuK��Z�5�ʷp���V�^z�<�.4�.лG�v1�Άb���AX/>�N�4Z.s��Iצ+C��ܺ��K��~����o��8�䰭�����}�D�N:�c�=����ld:�֚��ًvr���ϲ���P^R]�9r�(.�ڶ�j=j���,F�Q���-��oC=k��7*�<��i��lǫ�5�}�,����Xxv�Q�Y�;ޑ<[�kA���x�T-�b�<�����I:��Ys\QX���C-�Tz��|E�pq�}>6�c�P�̕ٶ;��AN�J��w�R�bz��8ꁍ�\�s�v��}�ad+8E��{_��:{k�l�9M�U��[S�QJ�r�6+�妟9睱\�k��|%��n���=��H��W����mQ��=�yoCX9H3��ȒI�w� ��q�y���.h�܀�b�[R��t[���x���Mk��Ǔ���΄�<�r�JU(t��>��I��JK.q�9U�Y��M־��/�}���x�W�Q�Bﻰ�����M'0��(��%�o��/������RҸ5���l��9f~D&�1J�ؽ��|3Y�čN�	]�Q���|u��%�(�v����ە;���i��[6r�\m\�j.�l�&��������a������7�YHF�Y�q���іٸ}D_1�
��H��煾{]<��_Ѣ�=���b��]^�ӁI1��[�Vh0�r��+sd�(c�G��P�ʦ�怩��#D�	���s��yz�Cxr���M����`�	�܌
�	�(q��@��ѽ��nV�����{H*��k���5�se�v�aT9Q�Y܋�P�Bn5�WU�ȟ����kc+��y���~�y�|֥���}��8�g!���__ܝu�\9��r�ʯ�a�C��k�-.��d�ٙ^DC�؜��+Z��]l��/'�ó��;��ʽ4=�T��/�){�-�O�29k!G���K�.�^�9�%p��Q1X��B���:���u�{z x���"6�z�~��CA�}C�\��&�(J��1D�b�J�I�Ney��^v{s<���fyۛ�9QH.�*�9α�����|1k�N�:�L�Mn�j��f�z.q
��\�N�m����'��ʧe��V�d�Xў�Z��,;:�n���e��>-<�{��O 4(����1�ܝ�ϣ��������S�P�=����:-��)h���|�
�e7���^���>�\��|Z-%���[�P��_�k]��3��NR8��zM��57ڨ{ϋ�p�3�����*���F�3��*jв��j�Suj[S�f
��5�^��i0l�!\w![�C�oD3*��Z]�lV[0+]�V	}'�a\8����l:h�Tt��un�.��ӊ�{ph�Sp������.�f[}S���[�,A��2NK��}�b�0!���4�Y��R��nZW�O0`���2�(O�A}M�}�E78t���y����b���jk�1���ҫ��y��]����L���*9��t��|
T4�o��7���O��od���q9W��jlc�f�P���7�+��(����:snM�����ڮ1oL�ʼ�u8�frmn7�]�ک���5	��qLƺ"c���Ne�Ŕh��������ۗ9�Q���5g.�V�������O*�]���v�n��q��_���}eM��k"[7���x��NQu>��$�.��y�|�o�I�&ңO��2��03D��+�r����"��uk�5T�v"�Xj����|gq�?kg�^Aک�KG�NuJ+aw�Ϫ�V�s-Ӥ�{5c�XD~��vD�Uv�fwHj���z����9����Cx)���W�<xRƟ�u��NOݚ��p�䫮�iL�$-f���=ߢJ;2hs��l̎��P��gT^P��� �ZGj�$��G4��/�p9gr�q�M<� �����J�o��b�PX�s�g�Cq�眹k�}h�������Z�����9T������0`�)�*�Z>Ϋ��*_WAu�ҍlu�oOWΓ�;��g�Os���ݓٰ9l��A	�F����+bR�P�������چ�ТUs!�]�V���ղ�fS��p`�#�La��t]D���~kZ��*�J�&b��F(ػ|����r��_

~�O�A	h��_ ����
K�W{���fi褍b�N�-�䯏�
r��e�܎�1'-ҭ��9��t
�[�/�Y7���6�&�;��y��y�e�
Q��7�o�����GUX2�j݄��ݨ�M�w�vøF�aR���U�d�u�熧V�a\�R騺]�q���S.��i���k��%��Ó��U�X��s��v�f=��χ�F���O���<k�ۛ��
YV�����t�����29��KUD��f�9���/kNЗU�3�VZ�喰+i%��r�zn�U"�j�d>�d˗�K�B��|5�{��T���N�}��ݍJ$�5�'w��{�S�q������֎��."��P
�M�W=WCwM���p��m�ǲZ���yn��E����{��6��l�~��<��>ۍz�*�/)���Z.v��y�
U��;P�g]����|�1{�%`^M)��kxn#�!�7��wxvy٨�u����Ɏh�s�]�bB�i�5(��^k��L���&1�c��<��X��]�{?[���fS���I���:��0�z�a�Elo�N���Ռq�1�\���<�]�p��cp=��YCv9񾳲��z�uR�iBW]+�cb��7��i���}c���S�Զoz�_/�!����=�T�kS�Ν���6�e7�]&��.0n�p������P���ࢾ��VԤ�!]C���ਯمw�뻘�1��)�kF8{P�R��P���La����HÛ %O���tEM��V��}5��!o�8�q��QȄB����͉��-���q��U�E
��)���uR�b�s[�\Q}�ՍL��Tg]i\{~������|t�
�+��v���L鏂�{AW3YO�6�u׎�W�s�?w ��(����ËݐD��_p�|��b���1d����:��B��nQhjF����v�w�tz�����oW�{��R҇z҈06��9d
�� mQ��΋�����-t��K���6�����o���Tu��ڞؕ�U��fz���:Yڈ�sk��]�w'�������U��nj��Ķ�W���l^�f�a;#��m@w09��ydo�xy�ju�!�����Z>j�o8���Zp�|��p�r5��t� �ڴf�7����'�m�ayXO�N�{�/mF�Z��Վ��m��Ն��V�M�,�	�u/K[9S��W������n����//��k!����f�0D�'��ZQ��7ҥB��ɛ遙�s�S�v��|�L�a�=�y�eեO(d�R�+��)��ݞ�|3*���Ss�T>��(���s%sc����S�S�(tR%�/x�,���F����s;*!�ٷŇ�̌��DerrS~�/��i4��u��Vg9�Տ/Hʇ@��š��7W�j�k��L��=�(*��J��e�;�r�u۰QRV^�^�;��ЭĴ{��ZE�� �J�z���K��4Y�HV+�i�^��#�:,˺���Z�X:�y���ҙ���4���?oy����F���T��<�r��d2��Y������
�j�`��O8�^8k.1��-=���O 6J�'o)-���Z�v��X��ӅSϱ]Q-ѯ�'��Yn8�|���T��x��n,�����s����>�k�ZRW���q-�r�--k�\gU�2P�2�S����=��Yu�#w�O�!%�G5}�;Ե�2�A�p���D�Ͳ���J_�����î�ϻ����������itVU���]!ۧuw�.��w���9�lT&�+�L�̫�ps�mTޏ+H�W�3�����B���X���3I��7�Tb�L� ����8�|U��|��b=����gvKֶ�s�m����`�&�]�3��1E�=g8����z�Ȝ��|=.�VeG�K\��]V�'[k\9���y�ʐs��M���ڎ��=��*w���1L�:���hr1b���,'xxlSz�U�w�x>��ݏ�F�
�37n��
���9u��l�G�!����fq�smY�yz��Y�)Y��g3�3�D�krrN>A���=��(î>���Q�9�����Y�m.EM�l��ߋ��;<�?T�e_M�T<������d�4E�L�}BvZJ���	X2�LV>u_T�oa��8�$�{��i�8z��q�ke��|A�֖�9~�J�s�z��1n��`��m�O�Uz7�ڙ;��ڹ������*�QWz�I����L�}��mb��#2_�[�k�P1�Q˛܇i�}��:m��z��˸znaʶ_��aC~zǕC�魮���Q���妟\:On ֻɵK��[���v8S=F�Հ)����Q�=.���R�P������p�Ә��"�<�z���(���yV���0;���t]G�ޚ�)�N`��Df�O�ܭ���j��y�*!JT()����Z*4�Y�#��$S�USTS�݃��Mݔs����<���r���S�S?�?�!.\���ˊJw��vv`�X%�D�fM�{���Tx�XF�/�xic��Q�bL/��EK�n��(�&d\5z����,�u��h$?������6Yb����4	Xֺ6Į��w�A�`�����6�뜳�w:R�0�X��lU��ohKlps�R�D��3:^Wf7�;K�;�L�y�E]l�����!"����^1n�q6����띎dK-�|lꡙ�wD�ڛv������w{�Xv
�[�Z�����5s\�;>��f�k]I�4�߁�6b5����;��`���:O��ֶ�V��[��bwh 虿(��)�d���%lЌ�I��r�D�*+��N8s	���2����)8��R��D��>��f���8r�wX$'9ޅh8۾��w�=�AN����*'���ڻ�E�ՠ:���r�<�Lu��ѱ!�u�N��M�+>�CS�T�*����P�#i`U�d1�ɻ݇�q��;�EHE0�f�N'9�ȼ�{�X�������]�4�WHb��@%6*�]B��ѐۙ3��ᆃ�oh&A��e������]�G��c�,�-8�[�N��C�M����XV��j��bi�p���x�u��Zƪ7����9�,.�+G��e��FR�O,�r�[�[N�Zgk�w`m�.��V�m;���t��cZɦ$�}��g���Xע�*�����T7���~���[�u�1ri���T�ۍ�\��$\l�Bb�m��Vu�Ɉ5,0j����G"�$�q{�����h�k���)�"��H�����7����(������C���؇�q��ش��\]��**]�:��$^'js(R��s:��bᐿkpe��Y���ua/��pL��9K��罼�1�j_��V�RY:�$B��5��Q���}ف�>d/LÎ6���j��P��l�`ެ���Y�1+�K�X�F����s�*0)�����c��[�3S�rK��g=���p�8����&�bי���*-#��yA,��k7V�}�����ꈼfV���2<�k����
��1�D�f��ZX{����q�U�p�jt؇x��	햷$E�D5�-��س�3wc4�:��� ��+`���E�L��G�*����r�,�m^Ed.3hTė,#_u�֚�N�ͦnb�f�=<&("&�x��z.��uξt�vh�Ap͖f[�!�q��=y�D���'���*^�����Q�[�F);t3�:�_	Z/���#EpݻX��*$�Ŷ+�ƫ�i�rU2�r�2��[+h>*b�6�Z-`Gw@ۙ��CX�	����NF��̖sY��"X#ħ���A�7Y*�à
�Rs�-K�f�z�k50���,ԛ�^+�-�wH`��p��C��;OI���*i��K��¹���o�ު���=}�`�P���v�)F�$?�MPQC2��Ҕ!A�JiC�y�\I@4:��%Q�Th4��CLAM#l��X�@����[m���"$��Ӧ�l����1)J��BP�q1�M�����(iNA�((�$�SB�.�C�A�J($�N��ta�[Al����ƪ����i6���:@к��qP���1	C�Z]Ph



@AGďA> �=����n�5�f"qJق	k��wcf�gprwp��p��4�J;�s���hʼO��]B&/��
`gqU�W��=�qK3D3�_=�	4� <����Ȩt�t��^ԗ|���J�ҷR�BZ��������s4���;a�7
P��FFc�w�� � �����M]>ٽ���[}3��Pۍj�����I��^&[P���l[��+��2���YѪ�_�:��]�WD�Z���p�Z�ٵ�q�sʯ�]�:�H��3�<��7���s�)^��:/�u�(��p�__�\9Oh��;��f�1��󡘪m�ێ�NU18�;�WH��Wѹ\�/��u��9_z�c�7�]�w7�l蔸Z�hr��|�ms������cv>ah)��]�׳n��ܷ�9u��ܩ<�jz7��誁�c�ہ.��:1��˛�=�Uۯzj���ꐆg��p����w�G��d�ͥ	\t�6-Cw$<�sﺰgd٫���Y�sLʉ��"�m1�|�`!��+1��fyQs.m��0_r��N��x�1_{��	v/�5��sl�-�V�:xa�id�-
R�}�rOr�rt��3�	L�S7a�EE��d�;��l@YH�iYٖ5�
�՗:�jx��.׎/|�y���ț[�o*�z�q��1��$�w��B�n�ڷo73gBY�7��oz����A��l���y];Gx��[yY�gM���f�����,<�
R�C�;��Ejr�'V�vnt�rĦ�e���{[�_K/u����ڶ�2�B!)��m�'6�k��/9�ۃC+�TiifD�P��Qi �Z��6�^fWR<֨��:�ꝅv��/�Dt�t����]K��mF>9IsW�oI��9W1�aS��������F��y��+\�E���N�֋���V�sy�fW�R�7��ž�n�z�� {��.��[�e���i���mJO��1K}��Tjӆju��C��2.��P���sI��|�� B@���Z�q���]����7*��uֵÚ��r����Xn�P��CS����Yz��%�͙lwe!�e5Գ(����8Vz���~Q��-�`�f��,m��f�F[yg.8��`Ss�&�.�4�0�r���:�\�0��W=�w�h�&|��p.���7�cq)�����
,�xE�+;�y�r�.�C��ɹ�,(Q)�㻰)hEV��Zn�V����������z��W���H�g~���*/v,"q�}C��iv�T9���X�ڙ��C�}$��0§�3�K�I�7�a
u��kӕa�AC�ع�"j�n޷���Q}�k$~����E�����hqʰ�i�vT%���
�ɫU�N��s��г�n!V�-�i�î{f�c��TRg��~���ΣK�2�N��G��~]�끭�8j�cO�%�����C�9���&дOon���a�X���+��rqrz�5�#=�|���L��ۧ���77K��$K��qP;��)+�mk�o�9}���υ�]ب�>b�κu�a�YdSr��PS�}�?	-9��Gz�k�-+�v�P��T^�k*W_%N��N��ܷ�tT[c)�3"�|�[�'�kޞj�>X�V�X�.^�f���Gp!��Fh��fbgưm��X1T�����]�^o5��s	R�z;SQo�<��yQu۵�^�z�V��F���v+*�}�`Xʯ�4�NDv��=s��w<Ǩ{�v��C&]n��0�Xw��ٸ����^V��S�so{�o��ؤ�E|陈E����+\�;�'g���]�d�l��_$���g.g�|�n1�W�o�Cg�Sꮾ6���u���p{�].ٽ紹��M����k��c]�j*	�ݾ+o�"G{�c8�Ȟ9�յ��������sO/�qN��UE��̦���6�v�}�b^e}Դnju�Ox�yC!uʫz�4��^ǍH�`^����֖О�K��>ڈ�e�r��
�o1��%�w*7���G"֮>�[��n�\G!�E\�������S�j��{�+V=j��z;Az�u�z\��j�jwHaxY~޿-���q)�jv����y+������
�J����Q����7��>��۶���8w�o��;N�,��\��%���&�mOMm(*�Z�X��[���O��{�QT;���Y��d��
�7G���ԁB�P��@1D�������V��o�D�5�Eܖ�9�i�p ��Y��m^,I���@ U�O��ں�}���&t}�\��P�b�6�|M�ɲ���k�����8�oBO�ja�հh����N�����T�p��WԀك�.['��]�Q)Q�\޾^)f�Wu��]�O=�V�v
\���O�A��'�=�|��[�׮y�Ս��u�Z^x�>��t~��y@���HW�>���-y��[Z.1�SBuLe߽}���I/���%r��|���ŹJ���yu{ϟO�b�q�-�	4��o <�I��t̢T�n^� 2\�Xnrބ���p8�����3~����3P�������Z6�Q)�6��z������m��뚺]�q���S-���kםG�j��*�_��O��PN�!�r�pĮ�'�cb�í��3%<��[Q����Z�Z#v`��+9F��T�ٗ��M&��|�Uk�'X�khgLw[K_]��OQ8��>H���Oc�V����{gj�ț��_:�������Bk�f����q�@�j�%Oj�����c-��n�@����-���ɡ72:];Eu(�*��]o��N������s�QS�Jw�ޡ���P9�eMp"�gq���
2m~��3mY�v�W}W��N�K\�@����hᄜ�u��nAò�s�K��������_'��Ӟ��=��BK3�y�0ʘ{�n�����z����ꝏ�G�	�>��kk34�S���XV��8h��3���S�%CW�����̈́�=���SqcC�5۔��f�K;3;5�n�����g%9�P�c�C���
��&��ǡ��|��=�O��[���Z;�k���'�h�q�1�a��<��?L�/U��W�܊���6�ٽ�:c����ޝ�$fηU���uߤ���
����'�4��=�y�P�*�C�;��:�0�kU��"WdT�u��l�= ����w
�M9}Q�n'���2����Y�瑏Vl��5��QF;����.�1�]� �mv��ZH<�'�.*�T�j�ֺ���i�àu�R4{7��簕,5���c ��e��n���{Y0Q�[Cd��*W;��P�#"��ke�Vɥ���A�(ɃC:���u�8m[����s^\�6f2�������o�1��a�p]S��WЋ�.��Ơ�'$.�q���lVeԹFS��Ldu���˳�2��k;xd(�x4�Z�vN�'R����!g0h�]�;��e��5�0�7���@��9�|��2�;ܧ��E$�řɵ��V*��k���Bn5�WU�Ș�c�غ�9��I�Ś�:gn����b���w��b�W�u��Ú�x2a���3�;&ɞ�ۚ��7}�.z�;�����Ȏ��wSQ{N������kY��:�i܄!���TZ�3m�&�j�SјE�yBy�������[�M�t)=[+���m&K���]Oԇ��gϬ��o�%y�~�)�9K��UhK7��ƪ�p��M�/9�bW��r��sT��_e:�9�{	N�o{��1��oH��ojZ�=N�+�[9]�H��3���jů��YӔ4������+���g{�{�����8^{	�e��P��Rإ�|h��Uץ�C��շ��i��8�e�}*�������p��5�I$�+K�S��;1��6�����Ž�(����˼Uޟu�mv�9ٽ"DQ��S�]t4[#����lq���d̓ͅ�"o�Ѣv]]Ԋ�qW���TmO;��*�R�Q�����E�x�,�%sYnuо��+^��N1��J�;��)%��xx��]�0�:r�tJ3��y��v�z-��o˳�!�����b�_l9]:J�{���|��K|ZK�qw5�y�߭���p_F���}$Oҽ\.:����܆�����)s}�O����h�u�߭�����#�>�Հz=7�,�xa�H��d��C�3I���{ת��
�z��̿�B�nW�6�>D��O��>�
sNfE|�=%HΨ�rج����V�2�͂��Cr�>5���k��������4n��;�G��ɞ���Y=\]��*�-2O���2au�Xb�{+�Z��Y�Lu���2��\=�T��V��o!���N֨{���ۚ,_�Ԋ��U�A�0�"�[��Ώv�1��:��*xW��1uތ�7��;;��7ԏ���+ژVv�Za�߭�x|M�P5ߋ7n�)��%i8L�x9�ԯ �c���]X�1v����1���1����t,��>�=�48r1p��;�!�l�6�tK�:oz�\��sS��+JZ=���Ǳ����b� W}�����=�1���~��[���G
R��W7��k��$�FM��곫J��oG�}޿�U�s:�Q�s��uq�Z*#�9'`�͉����a���AJ�H���v�쑞�}�8��f}��\\)��'>w:�gɻ��Vq�D��O�;`n��غ��3�̥����G�g�n!�z�\u*s�g�+���6�/���"�CR*���7�$��{7�CCظd��q��OY�A����>�U�7��3o�Vo����=^���Qwv�땱������lߡ��#�*Y�(�����.:�zs�Q.��q{ףOo��ڭBb}�4wr�+�wѾ�\{�Ǹ��¡Rx�qd��0�)���J��|v�����Ǟ�����E�f��>����>�3���W�T�s,>�l�� t��P�J�oY��S��9�w�U�H�s��G#k��z�8\��ӣ��둷�f��,�|���_��]��i��=:��p̴X����_)�oԑ�o_����&���}�zF��}7Nr/�;ދ@�ڟA���RFD��EGZ�g�)c��dm���-��ώ|}9�\� ?���1�H��`�e�S��%'�^;�:������o_܎43,�04�����Hî�jX5�u'�������x��9E�(�9��*�,m`��U�k��V
|zM��.�X{9βu]L�cEW%օ;]s2�/e�v�㭱��r�l�$����K#ű� ��c��T�����A�?\����UG��v�j72���}o��o�� z� ~��Qd��A��W���N}r�z��0e�1��/vr�K�'9(��!�'W&���up�~����eH5
|J��qfD�����Tܜ�~�+`=�5颸�#�}��o.."�y}���>�eD��ۖ/�p���X<jJ`N�����v�Ѫ�{z����O��9�����ڸ�f}�99�V>�����Vi���3��=~���f�WP�ς/�3c� ztu��i׉���[�q���x���������
�]������_��g�F?{�R��x�wn��|P���_�N�����)o���Mz�`�v��*}ꐣ#�G3܎�O���LO׷S����u�f�=QQ����:� �w��:pO)��|�;�����犤����ţ���c�#�hxvM��22�$�!x�Z�V��2����������cv�~��<w����{N}����7���9��s�7�J[��J��px]gZ��D���E_�Bv��OQ,�Vd���$2����Dͼ��j�3�)��A�PM�޺X��}��'(�z�9��i�GS5�����2��J�s:5���oW�.�6�-NY�6��-[�l���>O7	�8K����^v�n�r�8�>���i�㖉����������pr��y���"0������.Ѻ*�}t�ǘ�-�����=kEP�|滸�~퇰���4��:��8w�;�n�|;��)1B�5n=���"fd���ʊR�t`N�˄�6����z�.vk��5ʈ�֪��(�:�'���+��l�*�uc`��B�AY0��]���uZ���M�yki!��Hb�xf�WxM�K+���[��m�!�s6�B��̱�t�u�8�^"�����=��ԛaWk&㕦x#�7}��Ctt�ԍ�]nu"J�R�K������M�S�6�w���J�1ס����$�/8r��.�W�8o_[���XC�ŕ�Z��7B����um^ݬ���w��6%E�C�<9SOU����K����3p��(���^�+�g���f�z��͢�ĭ)݈ss�O]�g�-%�ծk��>�H�\��4�i�-��eֻ8r9�$����7��gVs���P@8u�������2�Bw#�s�0��Bh6<}���0�S.����z������Fhhvu�-<oh*�G���SXhq���&Q`M7t�БM����j5V[���W|H�C���Xk�a=���c��m�X�y��MVN�]�.�\��%���
�m@�m���+h��/�$vjj;ރ��񓰡�?E��i�����J
����wY��5H�����&;N��{���;�V;��6�#�~PhÙx��m2x�SCA�\��=Y�)(iu���G *�t�jv��ڔ8�NMuI�w4�4�m��k�qT���&�
tӼ�7X)�|�����q6]}Z������4#�W�fۑ�� �M}ݢ=�RWu6}6����F;��#��t�X^@t�F����x�$���2VGs��Lz�E���4�}��4�z�I;�I�IJ�v�.�B#�\0;����+�{u�u����Q�⺓�E�"�&`��s��OS�&4�m;���V# ӂ��b͍���jF��_M���nIr��Z�	�ζ@�H�J��oB�Ô	�cHV>zI�\�QX�ia��jrT��G��R���$��^���V�Kt��voh��*׽M�N:s3��A��;I̱͛Zi�v�f�����C�-���C�QJQ�VZjw��RY��^ϻ�Ȯ�� �@�p\ǳy��g��c#=×=ǖ˺�{������m�ǎ;c��^V�܁��V�μv�2��67br��5r����u�'3���9*g�Ķ[�v�e/6Ȉ�{Qy&��>�bs���b�z�P�v��j�lZ�$|�IxCTP���G'S@UhօĚ*�IN�e4��*ҺM%:JB�J�i��Z-�CIV�vαABklRM���Ө�Z
6΀�Z]ss�bti6�&�(:t�.��ZҔ�lRr�rt�4$LN١�!U��N��P�]����btSA��N��4q:Ӫ��Ԏ��m��j�h�1i�ESC����+E��6ZҔ�.C�J�v�h��&���Z�Z�ѣIbƍm���\��<�LA��lh(h�Q��%�S���:*���@�MP�
������׻fb�k{�%�T�S�˧1�n	�L+W�-!����J������,��!��箍�M�UJWK7y��2�E�wT�(l<��W�'a�~Ӟr|_�:���m�2�P(��#_��vՖ/���_H��q�x�GOQ�R(b�g!ߩ
�W���ָ�?H�����غ�t�lߜa�	Z�e��;��B��DLIo���#���]�C�C�;c"���HЏ7"sط�ܸ��}��O�=�q:mS��	g��O�]F�Z>��:�X��`s�}^xb��*۫������g�z
T�yӃ�߽8;wJe���2����/��o�r����s�l�L���o]�qT}O�y�>�I�Mׁ�W��k �l��W����+�K�8�@ru߷�뛶w��Xr[9G��|m�uǟ�T��9���~�����_dɥ08���b�9��]�͜s�z5�w��%���o��#z^��yp�]���7ك��w�z_�$�q���ʵ�2��t	�k*m�W�[��f��`}&��	���ۑ����u��qp�^W�_T���o��u�T��̓0��7>�U�uu0���]��2�3�H:Cd�{���򳻼T�2X�:�}��9 ��#�oj�[���9,�3h͉�<��;�
�7�'��um)��>|�ᢔHs��u�=�q�̵j��i/�X�1���׺��gW��U��Y����og%�	މL��t���w�{���s�xTg��T"�̳0��t�߫*��>K�@�%��z�u��ɧ��� zw��2"��zO�c�{~�Ý/z��W���	t��w\�с�"8|rvג�F^���>�s�9��L*�r�e��.�Ͻj�n=u¡t��מ󧆥г.���ۧ�|�~��s���*�d�)�w�����+�#�����>u��9|z|!M��{��mE�ůw��H4V����X���W����ĥ��У�!�b��H��z3�CT�k����vϮ�eO�`4�tQ,��/L�%�-��z�'޾.?^����b�����O<ٺ��U��|�*��PpӥP��rQ���@�Q�뉿�ex��j99�,o���f}��-ǜ�2�����\8������UA���S\@	MA��1+��Wg���ʻ]ⷮ��Ӝ����F��o��p}<=��^߽0	_��S�D�e.�*�Q���?s����Z�[��G����\G]$xg��}�{��ۆ��M�O�>8}>�� ��ә���M�w>�������"�F2�G��y�:�81v���	���W�D�8vĬ��{6n���*�Rg4�G��#v��m�!��Xqc�'Z��E&P�?'t�Zdq%k��.fD�l���I�����M�ḇJ5�h�}����8!�a���Qީ�����N��.}��f6�6*%ΣB�/��5���Q�y]ы^~�F��}���=s�W�0j��1�x~Y|>�L&�\���>�/i�622�{Ƴz�檬1����������/���xuN3�N�x(z#��"���Q�X��
�[���s�ݑ�lx��m��;j{؉��#c9*����{�>���:}fF/eH�,�߁��_ʇqY^���a ��ھ�X�yk�W����P��.���_�7�Z��n��߻Ӓr�KN���.�E�nb��c:9��p�*�'�O%@_-�'�D�+��d&��U�k��`�׋�v�o��4�/�D�P&PWt���z���� �}^���ឹ~=/�7p�K���tК����R;r����V{s(�� >�,:�g�u^�}n�6��a��xq��ᵃtN��f�_�}�p�[>�W���S�B2�(:��L|X_lq��T�Ӌ2�]�yb%����r�Ϸkf���z;AH�����c�r'&
�Ƹ�OT�O�EFԤW{v�������_kL;5�=R��`�v��%Ks+a�&^9	�-�j�fRGfr�t��0A)&R�%_omg_*��B��-�s���p�qt��<�RQUtcEK�}�n�O.؈�U��^�U"�{;v�vx/��9�^x�����)�/98x�7�?Ռ~�����?��^�3پ�=����k�a���< �Ȓ�4�*mUt�9�kڦ�g�x��Y�F��\M��i�x�*!�tu�}r7�Y��2%��qcٮI�w�y^�J��Ʀ<8��"~�ՠޙ�>���7��Q�߭�}�~g~>��m��[`�ç�Ҽ�.v�S�#�d�7����D�I|dWZ��퀥�_�Ypڿ�~�#�_��,ƐJ��>HÍ������g�j2+u���&�N��}Gc.{L��ԃ�~�;���W��Z�����G%^&��|� ;�����R��>���w�����z�`ޙj���hΆ/у�'�hd7�6���~��z��{jA�>%P8��}S���5i���S|o���l�>�S�7��>o�h��P�>똝���8G�3�|
4�!W(�=��7�{B+�;�=,u�Rp������~7��<Y�i��:����O~�ӭ�?ԵEُ]L�8y�sӆQbͫ����1`�j��*��������3�#�"]/g�������~�b7�3k"��Ѕ��ۗ�H�S��i[ޑ����泒ˏ��XJ�MϘ���[h�����VC��z���]~ک*ֺ�C<٫l�^��s�/T���^|���X�SU��#��;�� �h���7<٫���!㨾F%�޲��H���C��ŕ:mN���yP'ȱj���A�@y�π徵�"�5���3�������ª¿0}��=���9�W��P���>*�e���+g����}�=~���os f��>yU�lfz�w�w;"�=+ޞ��SY�Cò&���r�<j"J�2���A�k���SIi��䑞�>�r����hw��r7�<^��\W�xvNWp��K�խT:��ǎ��[%K�<�;��y��g�G��b�!�~�R|_�}#ǯ�j�}�A�e�����������(} ����π��37�l����}^�)}>���!=��v;�4�7�0�C͵G;�:R�.�=U�
�%� � �"bK}$_L�9��9�z�ឯ;a�9�2~Z�4���$�����Ol���`��Q5�3%��D��<LLJ�u떏�`:�w�Bl:W��P�ް^�������J'����{ՠ_��Ng�*@)��>X�`>��q��AҮ5���Ӊ<�cvz�\6{��j}^�H`�x�blwNL��Y<+�3/��z�K�a{x��gJ��z��֛,�ݷ@�ԲE�p-�D'��� m,C7�qb�̱���K���V�]���(�)���n��SW)�o+�����}+�|uK"�*;S�at�W[�(]>p�e�3��Z��x��l*
�$��J䈵Hg�z^��)���}���\y��I�W���~���.����2n�|A�#�o�M-�S��d�$����N%i���
_oS�|�.~��}��=��=��6�D�p�2�"'�i��;�p�G�%T��Z��N��n���<��xd7^쌛�MW{ Oc�V�#֯�)�B�X����B��t��%w!1�v�9Z�U׷'�-�_U��;ܬ��G�'�׬���]�צ�����Q�ʑ��s4�<4|��ΜǞ�0;�yR����N�W )o��F}NW�'=u��y�"W
���;qr��ۙxkT{���K�䇟^��z�ۻ�;���|z|��x������\?��qݟ}�+:rN��(��qJ|v�Fjʾ�䮝�%ze�P&P��3n������x�=�|^���_����lU��9O(gM���s�>��(����e0E��u�,ʖn��pׯÆDySZ���Bj�e�;�+�O'�׃9�T-��q�H����AK�#�m�ژ�z+��2���W�W���/J�Ron�rG2����R�
��#b��B1�W�V������&�:;�������&��n,f��5��8S��Z�m��Gv��Tɇ��h��4.|�jiY�q�=����(1U$'�Kt5}�Q��"�]���G1Q]wK$�p8������%����7�|��W�Bt�s��e�`�10[�&�ex��k��}�m-����d�+�wuE{�^X���{_��q�����G����ȍ�#�|կ�m)����u�>��[�x�r7��j:�o��9��/����נ_��f�s$�v����#����
��q�W|\�2�!W
�����)~7��
�mW����'� �s��"�+���|�k�{s���f{ffCr}f�M��Oxи�t��r�������Wtb�y��8�H���K7��z�+�*̓H������TK[z26�{�f�1�UXc�|���kf�i��Y�>����*�~�=p��,_{jA������W��*���k�"y>��t�R��a�g�4z!�����q�}�4��x'�����T������C��c��7i�[�i�u��k>59���t��U�\ϱ�������������䜾����)�{y>�d�_�]��n�(u�UiZ%%�K|�=�}2�Y7��=���%7�~��>�5s�މٮ��,*Y�cL~[(��[��q����v�hK�]Z����}P>�ŗ�O~h�w��:Wq�]h�VO�ҧ^�rb�6�tש�����y�>𮹖��:��+\ͬ�뭻�C��D�/�o6����x�|�҄������K���.�
�Q'�{Oa��1_��9)-�Z:V��t�?yu_��3��7�t�|z���Ïc�n�5��V^s	,^��C�f*3��M�e����2��,\u�z�S�ˍ��N>�� ��f�>콮��Gh�h��������C�q��vT�vX?�2�����W�!fTKا�Œf�@����Tw�#cu�G�O�܍��c�M�
(�x2O30�L*�2�yG^dl��#eU��룾�F⟺�mӿi��s������j�n���Y���bO}��!^+��>[�.|��ަ�3�^>����<�^��As�+���=~�\���4���ib�eL��۹�$ ��4��tDϝp7�_��/zxku�l��uy��g�e�$P{�GO䨭�?��tE�q%��M��M�/�gɘ���T�=�#m%l0?v�z+��|��ڙ{��:}�s���x�d
v�&�R��0���D��Q�˖�k9S��Vo����w ���=kμO���o��'��eW�����L�)_T�.��x��L��n*sm�=�.y��M�2� ��^o��Qiw�5rs��=��fz�tT���iٕ�y�>�}'د��|N*�+6��3.�)�u��v��x�X��/{o�ށ��wގ.��smn.�]��X�P�[6/��_�����Yr�����Uo�ƋsG�������1��ɷ��?W����U���mH4�Ī�p>.S�ͭ��U�'5�n�ޱS��}s�|����o.7�_z@�)�������fp�$K(��{~�\�/�G�rp+�:�e!���:{z_��m��d��q�O��/~�]����~�S�g;7]��������g�����L�������9GE�U�����������t�����D��gK��3bU�ez-�y����V;�:��b��_������T���}�q8��:	��׀I��˛���A�8�U����N�.�3���!�rO�ӶY>Wa�tV����FJwW�?N����Z��3�>o�w]�y��zȷ����e1瞻Còn�T.ʑ�r�<jJ�Y��x����-���7mt��/��k�U'Ǿ�n��{N���}p��"��òr�+�l��~���p��,̫U�� I^��B�B��n|�ϊ����U�N��<���;�<uG�\>��/�Y�e���[Ԗ���`�� ~�,	����7�[,dC���_�
��z�ё	ﭣ�M�z�T�
��� `?l�ֲ���|RH�焺�\u���>�{��AW���3�α��(���O���\��j��&�����V�ɻQu�:����o����������[��m�2��c'q��%�"X���)y,HG=��J6��h���]~���pv�u^0�\�iA*>�&K}$\t���fx+�޴�
��i{�wٙ����J�3�<V�c���H����H�>��ܚ���^$��WQ��h��i���T�������'�{��F�o����|ǧ����Z���g�*�=$t���;����q���T}�g�!����fcS���C�����}�3XD;�&iK'�t{�c�[S���;�.����Q-֊�˦�Q�^�{�=�?;�7�9~&M�����`���#Ҕ��ׇz��&O���(v�S��Jӣi�xVl�.9�\<O�h�C�Ez��d�TP3���º������=�r��-��O�r[ c�A���}j��e���Ǯ3��xQ�>�f�L�~i����z=��9��*�=�bF|��8oK'v���	�0�++�n:�u��	�ɫ�W7��V�{C� ����dK�^����w�ϡz�w���Y�jY;�a��P�z2�\����N�{���"$ޒ�k�
�[�쑑NW�'>��g�qy�!ep�ΛG$^'��U_���2	�̂�V�\�c��#*a��G'){\\��\�P:�����n��Ȭ�0�]�=���T�����8��xz[���(�����w#�2#+�.�v�ʼ�͇��;!F�8�Gegk[7#\��Z4.)�T-[-�A�k�h������!]�e�;���)����=s���#87�F�4J<ϑ�`|�D㸝�V8g3kGOYH�>\���̆!"�T�-TH`eа�|��eջ�;͇GOF���nn";X�g�7�F��}u����J=
<�wG�YC�}ֵV��+/�(�d�[{�LEdo7u�
�$��헵�OQ���|��#X70�$�ϰ�y�إG���&uQ���՜�&��4��5�\�����'2p"T�|M[��n�������2��a��)�#�	S/0���ҷ=O�b��^0��On��3j���#	�fZ|��U[�*�ej]JZ�u�e�=Qs͢������s9��Q�1GXWm}�'��`��:��O���W
j����/A���3(�r�j��Iff�tJPF�H����A3��G��u8�A`��pc/:щP�LOa3�t�د����W������ңa�8���4{�^zC�2�������3z�r��;�&Di s:����.�V^�uΑ��
��6�O���YWs\߃��hP����u-�^m��=��QkH��3�ˉڴ.E�g�f�7���b�<{�v�^zK]nɢ��URˋ$����5��K�z������d�j>�.bᆩ !gJ�K�K�NHVܼ���ˤ��w�_r�L���^X{�u�w��o�_?Llw[4�jX��O�� �����ϴ:�q�{��[`��(q����0��r�W6�)����i�2��]ɑ��Wl6�+5�m��;��rX��c�\��ΚY/�#���o`{�.���,��<	e��p�E���	��Ř�GHXƱ����M��P��
�X��;a�,�"�>m�w�Xp�K�%��s^M���[�u�G\��ilA�����)�Q,p��}�!Ǎ�.$�"�%�>��{&3}t�Xvĩ�Z�<��>����G�=8�0U�e���uK�=石޲��p~c�#&�uZ��,Pw�v�gp�����=6�q��Ʊ�x҇��9�0����M��(����R�F�1��v��˅;�Mt�l@Aٔt�֣lu�7�7�a�j�a�O��7�/'�_l��ƃ5;;��ѥ��S�Y��A*�{i�<�X�t1�a|�Y_���D���Lsۇ�U��5q��x8<@ڌ��M�uY,�t��W;E�6�n!J��`a�����l/)q��]f���V�ap���h�&�|�WY�P]��u&�]�����y�IDR�|y��-w��(�,ƵҾ\Q����z���}mC�{�h���X���*�'7S�� '8M�ز��9��F������E�֩bӈ�փ�tQT5���Br1�4�.-iIثj��%;cE�:
�ZX�AAAE	�hkZZ6�M�P6�:ZC������N�N�G8b�-T�T�ӈ����ѭ�rE0E4���h"�T5I�EU&�6ƃEj�-6�\�A3͍�Ecj��$��DM�\�%DMF�QM5T��D�ƒ�f�8��b��Q�v�1T-Q�DQ�5E-s�6ƚ���m�F��k���"֍�KZ5���+lQPE5�����_�,��a��~�oM%��R��#ᜭ��on�K��u��[�˲�jr�ؖ��Ϗ4�{n�41u����5:͋X���g�w�7r�6p��8�O���x��=���޵qݑ�w�K�
6sd]-]�!\�O_I%���g��+��3�[�.n5��<�ޯ����$�\���l��l.�{U.z ͣH�f�ܐz��A�,uJ���R��MՉ��~7V�MgR�T>�[;h�QR���p�}���_���ݑo�Q(�>$�2��/L����먟w�g��FF3}~�+#y�;��{�����>�2�#ʎ�{i	���>%� a���,�nǺ����v�ֶ�����1�}�����d��{a��q7�{�F�z���s%�B ��/��]G���l��j���G���`�3)��G#����m����>���߽z�x�\<P	���I���=�-$�>���*H���B��G�hR�n#|�F�6��m�|��������ҝ��5�w�AE]opg����[3"��=5�����n���O��^�=�*�1}�Ӭ�W���"w�
�o�
�`7�x��Ji@��`�;,���Z�џm����c�~j�����d��6"�ù졂�U�d�qy��Jv_1�N��]�J��)���T����-�2ٛ��.�۾�u��Snحnh��e��ˏ[�2��j�ڦeK��k���|�ybsX=y�Y|�1����&�+]����������J�#=��y;�}C�6�>z׳E��mH<|J߆L>��;�׫t�����I��G{9a�55���_��3�/�!��qϡ��x��u��7������w;!�L�w}�:n����j���}]M'�N��7����u^�L��Gy�/]A�ܽ�rmd&z=�zz6��o�·��)����&���G\VUi��E��ʣ�uK���wǟ�Gp�9��E�Mۊ�sg��̰��8J�<�׬��y�;>X�_�NW��U�So��_���{S�) ���#���W��^����W�}��b�C&#�Y!��w�ð7Tѹ���5mV��G�C�7!����J�o�R�F��$�|f�A�LuL������r���=��Zo�==�B���FG�O���P�z������F�ITf������wk�z��r��t�V|��'���{�&�ӿi��s������j�q��q �)�#�0�1���G�Of��d�"JCT����e�Ϫ�#/ʢTz�i�x�/�a׎�d�]z�ns�\o�c-�:1!�؏�X�3*�|F�k��~�������Sv�P
�ʓܰ0�=G�q�R�#�8�'u��r�]q��w�H>�ʔ���V���{�3����P�֧Nħ��7��l�{j\J������޵ghaX����Z��uX��Y��dT ϋ�:%��o��7C�F�*C��^��dA����h�}~�.$����Ø;���"q�A�D*�d2KS�A���u?D��4-[����z����C��sN��μ�;�ٙ�=�K�Y7�Z���D��Y=Qf�Oa��_W��\��Q��:g�Յ^�{�j���7���1o�:�>����Q`k�܃Q
Y=P��z�q5'},϶y�!�N;���ϼz�;��~��ϟ�\���(���}��U��L��|J��¸Q56�O]�|�=��������7�+��߹K��WP��]���@z���쨞�{r�A�Pc�}����+;Ӟ[2���A�G'�F��6�WO����n#��ǲ%�{�d'����wP�R�c;3}�U9:��n�~�����g
�Nlχꁳ���9G@�?���u0/|�~�ڻ\��'�J���^bM��qAއ�ݟug���S��d�����"�½�㆝�NrQZwJ��Vj��˺��#>v�~�/�]O����ι�4>�fza��zO�Ŋ��c4U��������R�I�W3��n��B�7��-�ܱs�To9��spF��Uٽjs�5D��o����[O��݇G%V�	�h[�O;bv/�e�����wy%Q�*o��C���[B��b[~��v�=�T�6f��(�ˉ+FCՁl+{'gr�v��3t�������h��}@s��P��Q{+ޞ߽�ǞG����S�WeH�,��"n(�����'�g�#䏌�C�sJ��\�,޷wz��7�<^�o���yׇd�pZ3ܙ�quT��V�^�yq��&��I�Dπ��C�����^]O���B����}�'��Ϸ�<yx�r�z���1|��7+����C�m��6�B�Te�1J��-�1��x�z�HU�>���z��G��]�o�Z��l�w�N�0��z��Ǫ��K8�����C}$i+�q����e��(�ޡ��7n������'la���v��wq����W�&��,� 7Bx��^���/�,ϯ�q�o]E��:����$h����J'������Z�=q,�L�6Jz�3�P��ꛮ���S��#�+i��)�J��7�j:�W�6��@�>� 7�� �\���F̯G���{I3�x�ǌ�ild��e׼z�G)|m�uǟ�T��9~&M�����ѷ�ec��69���G��ɧ0ʚ�������w�JӢ�m��VoS�~�(וw���û��sX��XO�:��v��ا��u�i��u�U(gw)��r<ֱӷ9+��{md�]L��J�vPuy3�[����wM�Yy�(���f	�'��vq�|jO��-�0Y��=��g�Bĺ�k���=��>�p�(�Ej}������Į�oaB�p���҄���{f���3�㏉T2a������t*s����U�]���zM_AQ�����ǡ��w��X����B����Nf����N�u��"3���.�w�r����@��+@
��+�.}Y�*��^D/U���<3�2/�wl�<5����&p�c���V���/}N��O�+>LP��d��)���箣=Ҽ�/�W
Μ��0��>u]�;y�`�<�+>�P~�XAS>�Wtn:��<�����x���^>��\?�U�|o�fѽ�7���^G�rO�ےOTL���q]U阸�t%�ƿU���^��G��%x�ۀ��U�UvO�W����*���3|j!�(�[�T`L�X��u��Y���¼^�Q$L�t�Ni뽿u�-����\1��:���{��}�H���� %鑑�-��g����u�k�|�^�zk�=�Y�Eïz�g�W�^Rp�m!:mӨv.K4���Fa���r}dwS1~�Ӌڵ!cq�>���[�1��}�qW�����:�:4�nH�z���s%�{F{w��x��L��!�m�ûx?'�ל�#*3�3u��U�dO�͈��>���5p�t�:�F�u���vW�x�
�;�"�<'@a��q���e�+��+]z���.���/�tM ���sB�ֻ,!#�S�,��AebR���+��5�O���*H�}\�#��j9�Z5m��8};��#�8C��@�Ϝ�!kӯ��o`*���&}�R6jS#�>�!W�h���)~;�f3��~��|��_u��ǽ����}��}h��VNi�Ȥ|zA0�
lo��h^[�Ʋ9S�mz��䬪���7U�WX8�u�nz���:4}����:�����&�d�a��}f:Z�Ѵ��iğow�e�D@�靎���/O�g����G���E��T����'�{4X���R}��U@ɇ�'t¿/{�S2����[����h������Å�^_�7U�9�CƞG��O�dЮ�T���ŗ��JNt]���(��|�q��Σ���6j}���]/��_�K���g~����z��։r�K4kLY�7�3c<�>�<�z&}��
��*���J<r\
�o�ǲR��9����1�P�������G>��Fo��x��:.��Ib��3�_]z��4�y�A��
�����79�Ym=��;�٥�=,|���dE5qݐ�Q���ʝ4>\e��x��3�;��2�ٿ��=ѻ7�Y���
:�=��+qA͛�C��gVL|Y���/gm�U�������U(=�yP��c`l-�G����#����0�9)I(N�0����F���V=NӣE쮡�b7�0����}[l#�&�VYyh����aM�t5ۗK��C�vX#ў�W��?S�^�Cڠ���2�ŖI���?2��X�XH:�˫�z��H뭟B̨�����X{�����P�z����
�%�Y%a��T���!V�fe%���t�0��̼}w�>�TK�^���s���oڪF�Ω��K:)�������$ߔ�5�I��>8�e���������?àu^���~�%��O�h��̟)���Mx�$qA��]2�p7�~,n��6�R���ُ;�G�{�P)_��o�O���&׽pv��Uxȧ2Z�&߇Q%yMV�x��>[�l�7Cن=�� �.�do������}9�^x�d
�v�&��z�L����0_O���d>�ʬ�Ů]�r1��yS���x\{�������z|�"��+����z������V���@vGUx<|E�C/����ӴR;J;�=�����!��ɸ{���x>L�X�d�/ǌ���}�</:��kuzD�	p(b>;8ҭ�mϸ�E�}��!�]���@z��lT�����-��z^]�+�Ը~���d�/][�]��7��;q�����ˣ����2�/�������`����}��h�$,b;{]��!�n>@��Z1��yz�7�
b=�-�*o�9[���5��k��x���2V�D%�u;+����5ۈq^Pz��f�$D����#�vg.=(jK
�l�w�᪥�:sK񽮨�F^ݟO�.�P�{��#֯�����՚X�3e�_L�~�:���M*�N�B�`M\�T��>���m��F����F�OS�x�]o���7"��
_�c��l������֬�0���	iU{ˡ�U*'�-���*!�x��k��r#�OǱ�!�rO
���qe��pf��;}��â���$��f���;wtmڠ<�z�C������^���X�q�<;"n�R�Wx�ݻw\�N)�Q!q��B���F���Y�ꡨ����}#������םxs����k94�T۪�����|T�ѯ�K�CS�����؇�S�~�U��i߸�G������M�lx{vn݇"�-�w�{���3�.��Aʠ�B��7e��C���_�
��k�i��E�-�}{8��,z5k��x�:�=냷�z��w�_( %P}DL��H�W��@���Xu&C=~�{f_f�}�{��pR�!�������'������D�C2Y��@n( ��6y�/�X�ʲ(�A|�̩�q���`��B��F�O,���q������`5��/k����=�����V
Z��V���`ҟu=�x/E����?+wԑx��E�L9���vZ�ᚏկK/�� ߦe���fu�kr#K�-���̎|��n�o��+��]�x�s�ֲG���>�"}�Ӄ�����@������3�n���xt��b�U���WD$LKt��B����~*#�f��5~���@��W�����0ۨ��$��b^�ɳ��r�2gޞ'E|f{�ʜ>��W�]/�����ƪ�q��d��n���չ�G��rHtm,�����+&MB��SG%���JӃcm��VF�>-U�?\/>����T6�����c��)ѿl�O{Քw���%t�j6t9>Ã�Γ�hn�C�L�ٺ�������uޏ�:�ddC�P�K؏*�=m`�P��8t1�/A�0̥����|�t���f����|k+���_�{�~�K�^�:�]�צ�����ʑ�
Y;��N�9�(xoɰ�v�}��_�:�*��>D��`��d��r��9��t�9��s��B���c�y���Yc��o�G=-��`Gk��32.��0�s�iJgr�&V���A5�m�u���*����ߩ���^�Jb���EI'�A�����}S�[�.o_���ޯv3���ѵE��w<Yt�����

�;zw>�B������F�;���,r�	��'�s!��Y2if�2�pTx��tH��\
n/x�T]�&�uə�'G��Uz�Zs{�wN�m-z�I[�f�:�x>�J�qY=��{e\cT�/��J�O�\�ZC:x���1\g������z�G��4�a�n-���,	�|�R��yfT��U���-��݀��y��O���c�yS��<��=�׌&.J5���`X)zd��{��}��]�U#�[>�+��t��$\:~�{>g�yQҽ���r�%�D@���|���p|�$؜�9��Z���C�w��p�|��&5���n=^X�A{^G������{�F�e���Y�Mߧ ����	C�n}�;���'��㌴}��r:јކ�m����>���b�m�z�NQ?�<�~�����}�3]2JF���f�I��+�G�hR�w��c}^�O
>޿^��V���w���g��ӈ��=X9�3"�zA0��X*%�xм�K�gܩ����8|:�^՜B��3�/}��1p��f��}}b�������0���W��މ���1�¥Ef:�yJ}\k��c����~����=R���O\B�h��ɐw�Ī���*<I�Y�X|yF�.1^����Eq�(�~.3�/����}�4��u��7���|L��`#��.��$�vee�U�/��E�3f���#����:s�$�n�`�����u<믬�;�������%����A}�o���mt�d-���Q�4�4�3o�*C&E�w��-���<w"��_!2z)!��ͼ} �#~P�FE�DVÈ�Hu�Hj�sw/�,XB���Se!�l�|A��h���۫2�䩄��Y;B�������}l���~�YP�mm��Vo,��D�D2�0�ɶ��F����4]uwv�
;l郫�t��U�w�En�~�-������W|"� o;����kv=S1���¯�ū�b/��{]�PD:;׻DS�
�w�a:O<�����u��N��_q�?X;:\&�5�#��5˷ܷ�4��G,�k�h���EM39��fS�f${��0a���U���p�Uf@��C��W�7��{pA�ru6
�'�1�H�,j�<%^2�`=���M������^�桮��<���'=�K�\�E�<��0��cJ�u�W>q��s�|��3:S�Z�ZI!(��,�ːw%w�ݣ��5�7�9���-��7�<���R���3�ö��R;�u��8[�>���8S{�����T�.v��9�l�c�j;F��<BpH(;mۇ�L9�����u2ys�o]�o<�s�ݓ�F�Z��K|���+~��л�L:]�R�]���TM����xV�>��9�+6l�I�>M{n�oq�D_-J�jY�F(K�&�E��:7�I݀����׺���� {zv�ǁ�ur�����]�J�	� QhYh]Xμ��}�̳�W%_`h�$�eC7	=1FcE��!���ʚ���@�
K�
J�O-`Q�͎��r�ܼ�E��4��8=�b�vg�헜����@���U�)���S�raU��G2�=w���7�~���}:x����Z:����w�&�yh�V��P��W�n�X��W)�q&s7&L�'��A��qhy���}�!w��j�[u�r��;KN�E��ȯyd�K���ͳU3�B��`�EM=��亝ϷtYj+�6�nW4� 1A%$�	�%In��Qk�c�\0.��9�T�e/�'�-8B�o��b�y���͗�Gk�f����ђ�Ԗ�8bd�+;���C��u��z�._$�յ�P�}�SE��ZI�ϭ`�r����s0F֊f&T�+��B`傘ٜ���v���X�k8#�8��*o
)!���D\h\6<	r6�0ـc}ݱ7�N�u���ͽk� ���bT�O�K]J2��#��%��sN�F����泃ӯ�v�xǙ�{���j;���T�J���P��$p���-���>��B#�RV`���֌�gyW��(�R�e'%�;	0?�G��=��t�����W�����)�W������#MMɍ���� ���
���$���nj*��+��j؃&�ͶgMMKE[:h����;b"I(�(��U0DIQ%QlF�PDZ6�&bv5UEQQ5m�4b"&��a���h��E�&
(�Mm��D�!E1AS1��:�c`��DD[i�F�
"b��EEQ0V�"�"'Z�6�cZX&�&��������l�٨��IQ[5U���b���m���H�*���6������j��)�j�U5Q��TEPE%EUU�li*�
��QTZ�U46�KF�DTEAUIP�M��*�(��ƍT�6؊	"�j(�4�4ECQE�%�Q[e�b(#f �2�5Llj&�*f�b*���� �L���T(��@QhǪ��2��)��qN;��\�nÓc+V^���x���i�/�%Q��;����͸4���+v6r|OY+��ScFW�p�ш�هՔ��5/IӐ�_�u*�Q.��靈~��9��;�&�/D19s�[u���ϐ��9'.#���ۏ���:�Uq�5+Ģ4�|�=�ꗏ����e��0gLgwH�K��Gu�����.��+�#�%%�o�����tY~c���� �Fz������^�"�Ϊ���5S��>�~;/�7T�y�S���'�/> ���w��3����W�G�V�L��� �;��a��}^\c�W���?�=�'8�䷪�rK &;�pǪ�n���ڼ6�i���C��WN|�*'��X��{ף������SҾ��
��Fn-w�n�珆��l����>D�:�z�_�t�x��'���{�&�ӿi��s���������6\=�4�,��'tW����l��� ?MD�7>�l�����S��z�!��Zzs��/nǶ��F��F����G����F�9��s �P��UO���끾2�X���F�Z�8��:y����=���W���+]�t�wI��\�Uxȧ2Z��S��"~�����+�z��E�וQwQ�l��9�ka����B�k3'�������#9��ְCbWY����Kk��P��N����.�~�I|!�c/E�wb�Z �n�zzົ��}�ό�p�S6�Hp{wY�Jɔ�䏴uX�b$[�/���pfoʱ,���G+�
���VFߚ�0��ώNx���Q�*���,��0�������{��m�Q5۹�����]GV�z!�c��r</�Wt-7^'�����q�W��rD)d�
��8߷�gq'|
��/*+�n�Nm�g�#�������W&�{���x>Q-7o?^O�q{�2�ck�*e��8;�����n�ۗ���)|{j�C~�G"z��9>�����fn�m���q�ݿD�{�bᕳ9ł�����+�UK�t�����W�]=�޺\j�r�y@���#����^�������P��g�#㳷>�N��9GE�U���Sm����j�v��[c��wz]/g��Nx�~��Y�*3�S�Nf���'Ȱ0J�}g��N�Vm��9I^���q�7�6��R����������!�s�£;*tݖO��m���;oEK��yj3�3�H�Ϫ6���7j�n;�B�YJ��}r�^����7\�(���
�p�|�3��u$���4eTz��F�:�f�[����^ӛ�/s��������֞R��k�h�5b�f^��.X�g
�4[5�[O�R��u3��Sy�)w���/!��zc�
6UvLEH�V��:�4� ����kBb�+��`
(^��w���v��#Ǌ�gb�ނ���+�y�%D�=ю,e��B���g&oe>�C��sW0s�g�)`�-	=�L�&�C��ꛟ�yu>7�U������l��uT��ij�,ns�|(���G��#\�{ڪ��8˸�F�<��,Ex��a���}�W���\��wk�9��k�+�J�cF}��h�zF���޸;q�a���J	Q�?Io��SckK����s�uu��^O{�fx+}�A�W���}�~���MǷ����z�i�,�z<��z�|�z6���&=;��ڹH��j9޵�87�L8>�"}�Nq�z��z�k޺~yk;�����2�n-L̯#���I���r���J������M_���ޤ����JDP{m/o�����ɚ��O
�3�B63�}Z*��x��/����|����C�ua�b�\u? �=�L�Do��=uCx�&M)�T��c���ةZtm>�
[���>�p�fK��_u��4Fo�����މ��	�z������||J�0�l�}>ӡ��>�盻*3/o;�4�D�a{:�G�Cu��ϟz�z_�Н[X(R�T���ݿ��� ���W��"/P"4GؿiF��1]3߻I�)R#�AY��i�.2��Ξ�B��{�}�����FU��n����zb�����1gv>Whwd')����6�p�;,���Ջ�}�Tىox��]�-F�hzh3����w��^�ќ�v�o�o��+C֢�	s�,Vb�eq��h;��������V3*��^/U�㝳³�R2�o���w�cѻYA*Q��>�S��4|��eV�5/ĬL ��\�NW�'=u�^t������x��
9^Ey<��w^A�+�s��m�2���:�wF����9z|o�Ķ{�����bd3U�j�Ւ�|�O���}��;���Z�9'E2I��eW�g����T��[�.o_�Ä�����6�٥GU�,�zd�VC����q��NqG����H�h��'Ĳ���!�G�k�t���yl�u�Mf�����>���p�!�cw�<u{��ݐg<a���#�J�2���p�{��>��=���s+�q��O�+���V=�#ޏ*:U�i	�q�C�rYI����i7�`��{*�3U�@Y�3L�Ķ^11�^�+���^X���{a��q7���7�g�m�#��s.)�U~�(���@	�}���x���Q��F�j:�[g �w��A��_��p���]m��^�jm��2KF�Kf���2�HUºh��E���5ܖ��dyɬ���G�VWw^�|�qm-�G�:��ym9���%��uyZ�otv�6���F�`l����Y%dٱP���^i5�.tط�F���m���_&L�>]b����03�DCт:�^�9+�p�y(��Z��� ���
��)d�r���%K�t,��>�R�K9�����������e*����yo�Ĺ��k���7��j�Uj�
���I�������*=���|FWO��5�z�0���,ط�ryK��~�sq��NW�{����ޯ�j����[�P�M�O��^�;�2
���[;>0�z^T���m����ވ�c��n�W/����u��73�)��x���^	�~ɠ���}���>=���Gz#Ӥ�|�gv��Y^DIzN���o:��dK���g_�;�z���C�{�fMy�������ǻ]5X��Uk�0�vzDTF)
��9e���W�����.$�Uד�3�_Qd�㾄��Y
��}��3�פ��X�'���Y�t<��e�j^���:��+9T� ��`��/�����F�C�F+���vY>Ve��g�漴V���>�����P�s�eB�C�ȁޫ>��"�1ǫ�q����J�kL%�R��d��<�� �Y已�
.>3���;�T�!fTK�o,C���ё�>gs}@{�=�c�s�'�viz�߰/Gfn�f��t���/,���s����[(��	b����a��u���T�L�
W+�,5�S������8���8=<y�v���r��S�޺s\}޷h��S��J�n(&�s�wnJJ��Voj�-r�܆��h�^��@��G���/"]��Ͻ��װ���s���vvrI\_��l۹O�R�Jr}"��`�>� ��K`7^㌶[顨�~Wq���G�g[�^�ʹ͟L�����u�}����fv�,҂G�E�u��~,n�sȢ�r���ӷ쫽�ؕ�s�m����l���o޸;~��_9����n:HȒ���������#�ر��]����zA{ܬ��m_�}�g� �sļ�����ND)d�	�^�#�!R��z���B��*1�[N��\��Y	W��Τx/y]д�x�`���:�b���l(�N?+H\�.:Y%���eED��ӑ�>���zu�i�?:�6������{j���k�U�]V.dgO�z=�R|���+��<W�k`����;=�2�y�Uq3�!��E�T��i/	����[>����{��L���jK
4�}Y^p���7���f�.�Y�W�'5��:7ލ�OM{L/zw�8�]��՚i���G�gI��p97'#:6�q�Nn���o�����[x�6��I�[�r��ѝ��q08�R�;t�y�&R!6N�ǒ���׺��ߎ�T=^�3fy���d.��wß�gc�)���OX�7�Gf��'��,�坌�����z��d�.J��:��G���Iv�q;|�Wo����R����D�^������c����F{*t����3=�9��z��b���Y\�{��℣<}����L
Z�x��k��|׿��|7M��Z�8狙����*4�e�d�+'�J^��,5UB�UTw����]�x7޲-�z{}�ǞG����G{��<ka�^4����R=qs�O�Kf�2��\ר�\�,�kwp�w��s}#���~����7'l�w���N��B{3�X�D�pW �*��Iꉖ�*�}uMφ�˩����WNx�u�y��f-�����.���#�T{U����2�P@򯌰&��7e��\?3����rW��f�|}
�!V�ֆ�������V{�o�LñrY��������zD���CG�rH��W���x�p�ւ�����S�w��D��^��fK5
�u�^��F�����$|��������o��>�j9޵�8_���}�D�>�'����i�����qsx�9H�ڇ���_�c5bGx���}G�G��~7�j:�5~�oޤ����=�׃wWT��K�~��]�����i$�a[�x \����3���0DA]rg�F��6���t�\�m���~�uLG����5��u;�dGe�M��䷹+��eb��V�y`��������� f�	��N�Y0����=|o�f� ��G�`�&k�>'�������VT����.�\y�>9~�Gcs����s�'�Jdɷ�P�wT8z�JS����_�Ӂ�Jӣi�xQW�މ�TϣTg�v���͙X}x}^\,o�|cz+�o�>��^���3g~��Ta��ᵡ�c�P:��^K�oϵ�a����^�'�#����]���n����;����ꍬ*���Ney)���N꧴3�΂��{���7�h;�j� ����u��g_��^/U���<953��a�܉{����ߤs,��|f=�%0���H��J��Z�H�r��>�����*�Q����ӽ��r�/۹��o�exTgNI�,�3be�+���f�%�?r���z|o��&�(�9�S�ajp��nVz�4����Һ���z��vG�ШΜ����'�&P���L��;�B\�&��P2tߴ�ºH�mwW��tn��V?K�^�Q�P�Q�)=S<�XW>+�\w�JmWė�b�!��ٽ-���mi�����^���1��������~0�����'�qQ�S��?Ry���ڈ�-���Pk#�ތ������!жz1]Y�V��N�$g1O��`֓cUs"���0Z�֜�rU�����)>�dd}��r��R�
*�m��c�ïK�E+��y3 �ejH>��*T���r84]��a)��!�=(󏽺�h*|���̋�3���LO�{��Eç�ё���V�yQҮ=���r����=8U��m�^�廜��q5�:�x���3Q�޿+��W�!�9��=��Hq3��K؝{Ҷ����|E��^�.r!����Anx�-k��h�s~��A�=\���r�`^�/�]��>/kA^�`��s$�n ԶnI�HU���<;Q����Tdꥧ�3}��.y�gѾ��nM�O�>#��O�̀�sNfE|�=5��^�
�TK��S+&�/��=�W|�l�8�gզ������G�{��_м�f�����s�>�$�,��0�xa�J↹�N��Z�{H{��z���T��oS�U�9�]�{��P�>z�{4X�d�=8�iSs�'{��S��i/�2c]����V鿡\���U��^߆7U�9��P�{��~����"sJ~;P'z��^�D�`���#/�R�*�r�w�?�`P�ҵ^�}򬍏.���8���Fgf��g�h�T=}�o'�޺��ܽ�rN_O�Ӷ^��TF)P��R������""|����|�9�a���q��4Y"�S���H�R_�_��e�}c���wd"�&S�$36[=#��9Z�=�Cr�vw�k��N��7�x<>�Ol��d�t������6��φ֌n�����M݆s(�e�é^���K$�^��U����z�|{��Y
�K����;�8r%�o�������C��?TPw�އ�����al��;<���7	���9���M\wc�F+���Yd�\c*��Q���� �{�>�:=
�ER���}4���.1ǫ�r!����J�o�.��r��я�f輌�^��T�"��$���D�p���^�Y��)����G�3�}@{��c�R��n&J�A­Z�v�Ϸg�Q(��I��O�C�B�q>3�uD�u�<�ju��/��]����.�-���s��||��H�j$�$7^��e����?+�؟:��+�(zwVj���W��ӌ�;�4��}r7�Y�s ��V���-��e����:�X�����-M̮�`�4�9*C�!׭����9�����z��EC�-M�ja��"��zc�F�^�s�Uc��4=��#�=>�r�6�~g��V|p�sļ���P��J,t�����ň���~�=��nN,>���	Vb�*�7r�Md%P�5��ŷU"���KȀ偶�,��}��G�?�APE�"��APEr
�+�PT_�PE􂠊��W��*��PT_���"��"�������W₠�����+�DT_�PE�EA�"*��PT_�W���e5�䙉��u�!�?���}�������@ $�R B�HU � PP@
>�0#�BTH��ITAU%IQ
-�)UEUIT"� �4��u��B��")I%EDOc%BU��ު�< ݶjٵ�,cZ��d��j�ֲj�I���2kj��J88�)V��f6��M�  9�  n�  ���,ݙŵ�$=UJ4�(n�#�)����mٌ��Le�F�V���mEPR���X�DFD�V���4mTXV �f؇mAٺX
!)��álM��:�`EP��)���Gs� cn��7L 2 ��i���p��9�����V]����l t��-PK �iRE��7 Z **�Y���U�)A@uFv@�v)��]�L�F��%%Sp ;]�j�X�e)5&L�ff�U�ͨҶj5�5cZj*TIT�. �8���Ŷ�4jcԲkT�՛,�f�	(4dK[d��m$8 wv$�0ږؖBZ����l�����h��-ml�
(�� ��R��d�&#��0�@�LE=��)J(�&A�A��d A<�4z�      E<�i)RHF� �hi�&# ��@h�#=MG���d�4<!� �I#!RB1&�(� !���JODGр�ͦflF�uM[�S��)`  "�`�J�Qw��("( �0��-A.�C�JB���T�gc��ɟ#������ h)
� DE�B�&TTE�*�����Q�&���SE������� �m��P�[�P��6P��P��d�7l������u�P��E�����?ԹO-�����T5�Xq8.�8�4.dU%]��۩�G-�>�� ޛ9sZ̲*fُ<��֬�Sq�X{j�úu�0f-�ehcvΐ/��Z�nƅ�!�����^yAѳA,[��j�cc(i�@���e^�y�i��d�0�e]l���k)^��R9*h,5V1Q���-^���E�Z� w�ܫ`���5���l�8�� o� :�� ˼ !��4ѱ��b��N�bw�t��h	v�,nM�fnU�L!�w
7�k
2XR�$LH�1���Cӷ@c��R��u�:ڑn����*�
�S�^+9F�AvX:�D]����ڼY�M��-��d���
��r�	� ��
����]��U����^<z/sn�m�z��������/ �M�
��s3�e� f�X!F��jͱdCPi7sX�f�7m�Jf:�C&̽ڛ��,[ѳS���!V/o�sF�s�_�� c�id 5��þ����vz���:n��NX4e�&ܒ�8g�+]�n�L�B���+�:t¶�r*��&��/��$N�0����(�5-wa9W$h�2��R�){��XF�VY�ڵ1�/t^�jƝ�]�Xi�pX{������ �� +( �[-�������+6��.W��Mce+�,� �l+Pۢ��F���tfU�u�˛/�X㵹J��)��hG�kzޝ,�0�	��XvM�ބ��#Lkjͣ�d�UۺLt��(L̑i�W1n-�\���Ca��yf�u�sN�,�K�qi��w{�����H�M�yYQ�z�m�ҭ�������1�(�8� �%c0���*�U�����e=��tlZ��+�3��.u���p���-���^�ȝ�����2�G7)�Z�em
�ǬR� A�{��V6F*a���@'��4�-�6��c�qe�GhT�%����/B��)ƄTN�Ȯ�<˺֙�n�<��WWؗ���:��@��CJ��9NT����6
������h�aR���d��'�^��P��Vsc4M�6=�6���uc� ���o~`;0 䛪eK�6&��Em�/sp�Ж�PЙe��]cu+Y3r�Š7Z�n�r��N<���
�b�)Q[�ܿ����kq4cQ���K�*ԃm�+hT����7I�o-����v���)�KcEYIJ�.��$��&��"ހ7w.����'nL2ġ0�Ϭm���I�K��m̍��A���ؼ��!��.�E�U��p���A�{�n�;}Q*�F�`���:�]I-�x����⻣x�_<-��Sl��QD]j�Rڻ�)ջ��k0�T,�w�S�e�i[Uwk��V�5��1����N�6�Ysw,��Qy��ނM�.���[H�6�=�jS{J'�5d"�`�7�t�wmZ�F�KY�Q�i�7��ڭ����W�n9H�ʹj,en��a��I �ãQ��V��]x��Μuy[�T�q���7��#��ۭ���l\@���c"i�Tl��WjJshfh�s!����#%j�r��,CLժY�AS�����W� 9RΓWbE.C��)z�5�0��L൥���.m��V�YW�VNSz�	OQH��4+oQJ�o�]�3�+h��{�-X���!�5�r@�I��HQ� `,VӒ�f5A���.��6������%`+ �z�eY�x�nԬ�N���� ,���kT�wB���s��I��.�is�nz����@�5���Yh]j�eޫ:@q770���n:iau)]i�6ʌ���e�i�V�k����IǊ*̭�Z�m�"j��yL� !�7)ő���ݡl!�r�k@�iC	Z���������� pn�4�.�d�� ���+�`+�ѕ`�,8��(W5�,�^ث�D��5�$;�m[�[MVe�&�1��CQ�$X{@m���x��h�[yr�؆����6!��e[���̳A��9Eiv�<yj܋�v��ۺf�Q*�SvP��k/,IYYt�����z�K6�ܶ�l56����iG-a�o Vr�ϱhTvҹupM�V@XJN�.��t(]�k-L��)�@�J��������#y�4Yј�ۛ��k��b7n��SVn]feN]X/л[G��%gH���� �QZ.�h����kv�[�Wf�G�w-$4�f�ܶ�V�ʉ
ǭ�Q@S�7.�&�5$]��o	/L}�7c���eФ��a�r����WwlX��a��$�F�,^L�^7s�l�E�y��j`(�P^�4L����\��ȓ�Y�����%`vd� ���ٵd��3�h��)Kr��m
�d����V���n�Tv8�(�T�z+��),U�M��	.����h?K�f��U��'�(��L[li�F�ɔ~U�E�{�٫��u�	6��,)�qr���J���=�d�ص�˟J�GQ��5l<2����St�חejy�gz��QPX�cy��9h��F�4���Mf
�Ȋ��YI��!Eփ��b!�>K8u��� ��J�T��ٻ!���W+K�e��.��h*�3(8��eJb�h6M���(j�b����t��!�n��z�sY�P�蝭S�7�+V��X�;B�A���K�[/h�����齴̕uYe�65n@�[�� �B`�����e�1���Bmn8���A2�6��X�v�әy��Zx%]���=O
�pY�%ø�"�!�15yCL��~;j7w�h-�����Uܨ�Ve-.YX�I�Ewf�oJdX�����lFٺ6�[Z���ψWi#J��#aV�z�(�ufX�`8֒�������;WD0f�/h�@�YLm	n�b%eR̭��p����sQ1�7>�.���y�]P�n�$�D��ͦ]f��Ţ0�>���.»A�i�d��n�j�4�؀Vdj`�C4J�QV�C�@(��6�ܭo�gc��
�6��E=u�9OV�a�Y6�d.�rѳ0� 
Yz\�u�#ǂ� `��p����+/]�$.�t�ml�j��C\OSW@��`m+Tw�[�\ްhe�������ȥ�p�/,[�^0�	[m�	��[��o%µ*�>#s NA��AY�&�>گ}�U}�_Ք(��)a[�Gj3��L����~��}�$���y̔�3'�C��f~=Q7l?;Eh���c�?�T��~f�a�U��)ʱ��9V3x�*�o�X�✫��JT���HwwI�I$�I$�I$�I$�I"I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�e$�I4�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$��I$�I$�|�t�A����p�*�z��,Q�ja�{Ϻ��f��4��<Z�A��[����ν���#G(4�Ю�e�8|��L�
,�\��;�9����ٷ&��TouݎH����=��v;[��Ml���N�3,&�!�+C4�� �o���j��c�xn����^�c&?L@Y�c(�;e���de�n|������[��[0��
)����WN[V<V�V����<ޚrFn��m_(���dݤmJ����S�!�YwXм�7;fm]ծ<-�\�+��������݆�V�R�m�9����
�+q�( $���X@ӍW*�V��Z���7h:߸��S9�K���c��stv��\Y]Y���,P�T-�F���nCn�O�ͭ�e���b�i���v�8t���`;k$��
�U�k�yjf��@Me�H�u:Ļ�{�pK�u�Qm�FcΫ��wá�t��k�ٮ���v�����GXj��_e��E,Enq�Q/�����ʻ�*>]�v�ÿ_o+� �>�rrҗ�܆@�*5h$P2�P�xI�yE��������q�x^2j&�<y�9ćX�[�b�{�:�2�"ؽA�(������TtM�^�V�����e���\��1t����6���n�j��-��<� �X�o��q�aRc�К6�T���.�Q�x���]�Q�u|�oR���0��[S�4�S�c�Q����D� ��2�t¸��-o[a.{�j߃�a����ݾ��Q�T�8�R���Zt��YXH<lt����]�2�e����G�;7.����x���r�����r`����,��7DH7f�>k���N��E��[�y3sX�7r����r�m���,Q�W>�������3�۫PY]���ۥ)�.S��C��lyә� �;(�.�V`���E��ѭ����%�u�rf�<����B:*�x3�jv"�wJ���j�:���7l���t�	�W�F7�;(m�HVc���'Q�+D�}Yt�������4����<�>ri�y��O[f� ��Cx,oh5a��}��`�����s��"���:�ʴ��O���1A��3G��Y�a����n�̑�����9A��t(��Y��nekx)@�`{�x�v��*Ġ
=ό9w�.d��%���,u1O��'�G����
i���n1�����c��fq�!�w�n+W+a�Zp^ݠ�<ak�*l���}薅�/<�ܫ����dڳf���8"���S+7z��ڊS G��7�LL+&�YᲛ}n��;������f�ڲ�l�8f�
�ͥ��w�C�o%����-�;T����\Ƥ��*޺Ω���S&�C§����\�@���SChu*wQc]DQպ`�N�*
[о�z ���.����c50�CV�ol��IK0�;OP<p�]�(�֬��C/��R�cI��������j&c�T�]�tYv�ޖ�'qݢr�����'WL�.
�wa��!m�E~�D��p�i�-��d�`=�����X]��S*�i�z��Rm=�B�����a�ua�R��ٔ
~<�Ӣ��]	3�+:���̧����L�B���������1Lk�C�-�8�'�� ���PY�B���Gpͨ8a�a��f���c���X���ٗ�o�fԎ��W���U�!�W/�9�5u�Ud-'Ҧ��=�pPw|)
tR���Ǯ\�J�wy����9s��nQ�A1�|Ľu]�E������mY=�J�����ܵt���fĖ%�s�AX�~Vh&AY�ժrD�����:n�b���ѻkn��`��f�ڱ]��Z���J_��{L�a���v�iE�9V�Ȟ꫰7��!@����3MP��i3�����
�԰pd;��X�.���Ñ��܊U�`����]�ɟ7mGti���*�s����v��ʗy���㭛kV�l����Q���suɔ��t��;�	y}K2��/v�m˩W�1j�����v�ժ3��5w�͈��CH,�z��8�M{۳o��Uȴ2���yz���u�.� �Z3	t���a&���jWL0��B�.U�Yc�N�+y �\6�X��z�
�d�W�� ��q��2����a^�����=E|���n0a�^�ֵ6��8VV��ʹ��^�x���1�A�b{L�1�&P���	#is{�\\��˘�!�[��:��D�'Q��e-�5�t�R�0��</5�g]��m>͡��j��^����^ˁ	Y�nڝP�Wb
|�p�u�P�BCc�^'�vV��r(�����_Ibm��l%W�������İ�Z���l,��	5U�&��[.�,q빕1Y��(`�8��`TN�<0\���p�o1e�茋p�3cԭ���U�]���o����Н'D��n��%ȟ�6��v�Y�d�+]ܰ�
A��[�3�1�t���.����ຼ[�C��jk�k�C�b�{��_��!��wXF����"xt�z��9�v�NP����v�Pj��C�"Lof9�������}���5-�^�w�)W�*pU#zsC�|�ݺ�T���YV��}շ�t	�z�K���b>@X��3 �X���Z�G�3�HlL(����_.�T޸N�r�_j�w0t��^ͽ��d��U8/s��
u�/xmM�6�\բ�Nӳ���̤��m^�л53��YX��2����o �\�#9�}\�.�X�%p�L9�_ݺdV&7c ��bj��]W�I�%�-��1�:朾��=�B����;6��`O���ӢGV�sB�գlf�aIk+:p�X��)�	�3���x��>�ZG]�t��@��.eE���&E�0��qC�I�]��xӗz��n$dm�]��������2YZq�QGCȋ�˦�;�jV���JQ�ĭmby%���Ԩ1JuM�Ů�>�)X�B���z��a���}�W��G��I@`Ĥ��J�D�RI$��$�I$�I$�$�I$�I$�I$�I$�I$�I%$�I$�I$�) ܊Pnڔ��:'�7�l��ӵ�,��s�KrE$�L��,�˻wfӫ7=yWV��8j�<�DZ�HZ���*��U�3�A
G�K�!I���3�����/է��u�_���u�^o<�gW+4�ѫ�+��ӄ�Q�b�]T7��<��2`��6�493x��V�}^vf
������qPJ�����_�X.R��f�'�S�:�s�f��&�0���(#�����}(����4a'{�e�!Wb�eA�A�=UN�+�&ݤs�����<L�W����n��
Ԩ탔p!Q�z��w=�x͌�[.��a�L�{C`�`u����7��mV8��4ˤ3_]�E�:��76�o_m�0;���R���!��ٺ%�5���ݕ�qn"��n��x�h�X��i;�컺WK&�~l�;���3��֎κ�!'-
��|�52��h԰E��];�^_�v�t�N�n4Y*a�ϲ�`��g�Q���1�
��j�n ��눻�%�� ��	�]q˘p���]
�)-(ܻ�b�Ycˬ���ϯ��B&�]Y�ٝb�	hBAL����g]K�%����X1�fds���о��(�7aT3f��k���E��O�s3W(ޔ�hj+W}Υq}�p�K�-���7��uD	�K*�9Q�[u�)����Ņ�;CV�2��*���EKQk*��2l��c��Db�f]��9x�8��� �ΐ��Id�����f�ׯOE�h��E!]L��,L`P���g�r�&�ݕ���4(K�2�
4O��t���t
��M|kz�mVN�M-�Ν���)|�N�����̐i���L���Y���eV��s�]����.��7zv��N\ � ��Q�k��	<�X�X���ӉZ��*�K�B�mhl4�w2F��vB=B�_EG ��\h+��cx�+�ne��%y�.�H��s����ơ��k�bԑ]2�iJIg�S//�ّ=����Z��e���qV�����cW�\i���#�F,�2;�c��gR���'�}�kWF�ð��jX�V]ä�$�η*C�P���{��6<���pʘ\7:��]�2�!�Ҕ�3[m�,�6�$��o�E����)����Ť0�nY��vWkͺ���u݀["z.����OM-���S�4�Uc�4*%kH��gΖ��&��\B���0`��Q��|ռÂ�ZF�K�wBs�b[��h%j�\ss�����eZ��
�⋊ (ƅY�;+F�M�1�
H^�����{N<�7��~�7U�ĀI�%��F��U����}^��r�����8,)K{�ʆu��Ju�pX�2�8�+ɺK�������J&�Zڶ[�a|�9� �l^��}���*��������vgw\�+qU�j�s��:�p���0��O:�]8Ǜ�a"��47#�TF�묾�l���]�t)��ٗ�#LR��mQ/�i1WN^�H����kOC��k�d*lN���X��W�-|C��I l�9
��ʑf4�5&��
����-F��R�Nt����mAx��.��Z��\��qP=:e�|�ۨ�WP�\V��b��tb�gq�kJ"�ΜY�]u�Q����g.��������s#�A	�Ӈ,S��K�T��'��Ҋ�k��f�;N �� ;��Z���*6��-M�m��ݗ����(	BYot*v��L$�g7��J�Y��[��Z7�,�)]�Վ�l)s,���j'&q���y9�����B��h391a��=�XE��O,�=�H#�iTJ۾�R%�C�4���RBsuor7.f �|��&�{!�]f;�)�X��K(�\�n���@ƙh�<0����%�|��)U�������.�v�%��t�T:!/F���=K5ݝ��k�p6�`_U���f�l��\4��>|2�R \9���}��k������2�w��NJ�Ga(��n�\�AV���/k��]JO��Q�� �o)L�.��0=f�gv��_j�_<R�&�U�5A��b�d����'l��Z�Q{�*����Z7W;٭���ia�QQc�js�Խ\���ǭes��]5Bk�'=6�e�F/��<�w[��<�Q��6�J0ec�it��N�SBB��w� }Z��XydN���mޛ�j�[6q�v�Ϻp+V�V��ܧ]-�D��Qh�<&��֌�K�Q�L%7I�������TʆZ0>D��59u��뛮�I�B$�Ф�T��0n�;EfZ���1u�Ʃ����SQl����B������7qW
5��J�mj�����0����>�>��9��o���i�f�"�F��䎆J��Ӯ�B�oiB�"��m�\[/"M�v���K�B����������j�Wq�̣uз�i���e������"�6�ռ�v.����\A��k5�
6Y"�w�f�V �R݊�w(�ŷ��+��ݪ62{f��� �iU����-W�F�ě	�˵�S�%���xṂYd빛��I�(<��ʾ�x�z̣[��X�}��Bj��5�֤���:s2�L��%e�f�a޶.�9#νYw�9�Jܣ�U'ˀsFIAhn���Y[6���r�u[dn�anT��iO/��YY+�x��1wF�ACWQ�h.�OL�Sn� Ff�:Nf]wjKWa��4_�!��C3N�Z]��+�K�����4f�o�[l�V'�t�l��U����[��av����� ���X�^��eʃ+p��*׳�4�Ʌ&���b��댏�"ʦ>uyf�N�vV(�I�J���0��M4�X�tG���z�Z}�����ֈ�1m[����0�.�&ɪ^Y#*a���]���$R����L�t��;�Ϥ���2����؉J��X=X70>yn�D���b�30	�l�X�x:��9/o��naw-kXYp���e×Eb�)u��l�؁�˹GkL]J�������M,ێ¬�65���Un����C![�����c�iX�l�-0�G���am��%oJ�4F�5!u���.����wW�/uq�VX-�5�Y��z��R�v�#>����ʩ*��a
ʗ8\O�5�t�:�4"$�OS��e�
�@�/2,��QN��9+L�y�ݺzv1B�Aae��ɀ��]t�]�Sv��U�|u�C3��C��9�g����O���BDd�hd%�-�L�TK��#��$'_�J�i�I$�I$�I$�I$�T���g�.���t7�JX�9���7�S��p�ǁ�󂷧U���ʽV��A�����v��ી�Y+����:���7�E�}���,�u�|oez/� �&GB��X�u��p� ����f�ٽ�Ko��롢�M�\"M+�v���&�0͡�{��mʍ>ܩ�r��0�ߧ�#]�&3���L�۳�u�@I[݄��ղ�aID��)�)a��.5u(:QU�\�"&�;vzX�W�,�2\ʜ�[se����z��T36����� .v�-I�Βֳ�i\���������6cy�OP=�I'��s�<���P���b�Ɍ*I��5��X�KV,��3(VE�e�1�kAH(��Щ4�a����R�I�Ǭ�bAH��I��jH��0d��H�S��l��me��(bUJ�r�� ���GB�L.#�d��2�f*�T���J�[l��b�ܵ�j��S��. ����hJƴ�Z��\���T*Q*,���]Q5��SQ�3N��wM"�!X6��F�J�P���VJ�eKl����ޞ5�7�^��[��Ԅ��q��Jbx�{\�_v߀��{�������|�I��W_*Z1j��:~T=������ͺ�J�ә<�xk^�,k=Dt�*<��X9Е��yr������t��*{b�H=�W��+oPp�̓�Ү��J���^g=H�H&���M��{!6X��Ϣy7�(Ժv�4�,���b%�޵�^���T����gW��K}�X3*��{������{��b�2��W��K���BGޭډ��7tߋ��g���il��'N�X&g\�j`�Q<�s�X;Dl�ރ[u".\lۜ��ws�a���~9^^��<6�Pݦ��}m:;�E�"A��t��O���j�-�3����I�4x�s�W�����+��U�aJ��EsUj��Xŉ�y��8U��nU	������z�.�9t�M�gA|1�0�pw �7��s�7�9W�
��O=�:ۂؘ��ƒ�=�䷒6�B�;f��y�玭�;D§����T%~��&{�"Ś�$p�y�&�:��Qr�Z+���p�`ȵR����;�n�0�B\�\�r��w��Ql�}��%7_�<�
2���Mi^Qr�s����r1Ma�x��縚��Ik{-�T^��y��N)yKYћk�wU�4\�Q�2ȅ��U���U.�t:{^$�F����*n;;԰�'��o"�+��5zhA�J��۽lw+�լ��{��G���r.�=yFxA�O=Bw!����IJ�nM',�^Z�^�W���	��j��LE���ò��}C��1b��N�tw�9�#.��e�����]9�\�_��Jy�l��4��T�o������&��6�;6v{�"�-����Ub_��j^~G���� ���v�)o����5���<�,�&��^Y�<��<0�7�V�cu�t�t�`3f�I�	�C��K�W5z������~*w�<4�9������?C��bQp퓙�\�k72��s�N0h��VH�+=�߆{Sg�Ԯ`�{:0��{�G�ӛf�ECZ�����R�b_;=�ê�x�F.�B��[̀V�}�f�v.��m-�p�VH ��F	�3n��%�ct�˘��\c��n)ꝑ�7M4���S7E�QF��溶ڻ�S��c��������%&7���|+����v��E�����\��\��聻��ءj���s�]��dX���E�؎�y؂�6Cq��U���4�yF�$�9��ƪ�=6��mY99��[Ę�a4k 76&\��{�d����;o���m�Z���\�i^[}��ui�7Do�����+�%�怚y�xwË6zS��/c7,��$i�W�7��٧�[)��ŹkL��!-M��)�Ƽ%F�W�yI-�R�L�Ͱ�û��ߍ=��Y˗�#q$�PS��7�ZD������H��GFx[��Z�釣�8��z�p�3+H{�D����e-�˽z�7,v\�@���w��!��*sm�ٍ��
Ӵ��&�WxW�'�dʮ�y�-��
�-j<��pO�_�h�5O�{onem�I���B�st�5��HB��:1�[�ֳ�����tn����l�����p�q�6{&EԵCs��,��6W���e(Z�1�QU��u�9X	��}^�+T�Nh,I��$�f��s5f�՗�dh7qzOy*���݃9y�n�~�2�B��(�]c;�na��ҟ+�֌�S�}R��̕������t��~!w�ʣ�;oY�7�'��^�=���y'Y���^{y1�_*zf	�G��)�8����$c�SʎQ����:��u�|bK�ﶧb�d��A�Iq��ΉCƁ������7���З�^J��c�M-~.�>/��w�O%�3Eb�	 ��)�t�j7�ʮ�T��(lA���MñfjIH�B��H:)�.�<~#�=�u а��>��][�����^>�+]:ޗ^�M��"��I���ϡ�B���l���R����Ӵ!��	��E�ݳ��9k����cx��T�xR�b�
�iݘ��>��"7q�ڵ��[&{A����'��᫻it5�:�kX�<uѬ�Z~>u�� =�I:�x|ȥ%;��b��-�3����ۤ�b����/�I��
�F�EƓv��؝���J@��B��]a�!��r��,[�&�u���;�X�ư��[��)�ug2$�yrً��ia��e=n�3��x�[�:��N�-h�LX}攢�(��`�j�sW}����o(p6 �����)��Z/�ǩ�K����ш:��9lIئ��1��C'NS]�sB}^j��yy�aժ��G�\���En�����YÓn�Z<�/�؏����߱���k�u� ��ۃ̘��b�9�{��ht½Զ	]�Ngp��(�j�N�:��x)td\���ݛ�n8Y�Mu��b�wP^��T	�.�'!��x���@��!VO8Uu�e��ا�/+Ր�6�2�1�}N7]ֵ�;�����`���������T�xJ���<���H�2��g{[L���ܻ��ko.b:�b1��u*/�	z�oRa8��;�qOZ�]��a�d�����\�g�2���X�.8�f��0MB��w�7���M�?W�dA��g�g~~w�wp���ҋk�]ma-�;�9��F���;xՈ�)>��O_$Ѿ��َ\�яGLV5p�`�H�i�n�U\�c��eX�P!OjL�0��i�B+j��j�ֳ{�T�kF���p�ۓ/,� @}�)mm�����,�"ޢ83񀫼�R���'@(^�������E��h\�*�/]d�����ue��R}s���YR��vM�K�H��ZB���r�7�`�J�<u_�G�5�2>����ٛ�g;܊��uЅ���aw�h��):D�oj�]�+D�kw����n�l�����fV�ng�8�	]��CTA,|��\g�M�E$�I$�I$�I$�3��Vn1SL��]%R��g�݌���1�g/�nıF����R:{u{ېZ}|���/����.K7��7�Y�JJT�.(���V��=�j��i�֊ξ��y����B�ږP�<ʹ�LMM�BY���Q�ad�3P�e*wg��ʸ���	�; ��?��;y3�`\��՚
����-=���ˢb�=s]��)ٚz��R���Ȃ��m�+p�n���{\�S�Y�+�72dF�u��'*�R8��d7�!��:��]���8ʛ3=d*˛�W�^NqR�m"h�$�(Ӓz�|B�]R���ȩ�+�MVm�j�����ءl�Z�ܰ��B�ƧHq>IFb^�f �(�PX�UB�ëI;zH,�* uAfe
�<�Rf��e6�0��&�T�4�13(V�X�d�l�t�GV�=�N%EU�(
*��D1
"�QV#P&e��Y�]��I��w���6��������k����9�7����V����ʿ�
��x����+��ߔ�ߨ���s/ݩ��G�_�~�����93�K�:�����Ω�����j�G�l}m����&��%�(�{l'':tD�בP͝����u\~���wzj>�n�y�]��P�p���ͪ�z�:&�v����+E=��u�ʖ*W$�/_���G���?g]���BR��Y��m[g�ux&�ք�=���]5�BGvW�v�9��\�SVι��5tb����Tkޫj�cWq�q�u�������L�Yc�2�.�5���k���]�/��J�7�ٕ�x�y/6}�-�D�gm�]�L��_/�y����cl\O�~�۴+e�ǽv�R�S���&����b�_k����*ϡ����~��ݝ0L)?�G���nY�)��[*���������
���V*�8+]-ʓIf���_F|������#�܍�@f��K�_3;����-u+���<wz�M�b� 8!y�|�A�C���'�~��"��[�����U�:ѽ@���{`Y~�;}隮.�iA��,�H�ӊ���lk��!6��R'�������Ēy����Z{W�&�@��3�>Z����(3�����.�ŅK�����"�d�؄��t{4�|afI��*��8x��=��yY�y�����$D�[^؀����Z�8eW[N[x^�!i�k��l�x�}�
�o5��5��~׹�E=Tk׾����6�CWk�^��=�q���qH���B�{yOu�Zق��"�赩B�\����啤ĲR���Sl�wjl�H�����ع@<���GT��ѯ7��"3�(��Yв���'��5'��)���5�YyUdW��Ʀ��.�u�Z��Su���PJ�*ݾ��{/ض?`�Y� �[��o�?Q
��k<s(#o&;�^��1Ȩ>)F��V�
�H�줱8������T:�r�ݸa^s�8��Vǽ�޳&����Мd3T4��9�{�|���;������ ��T���ԇ�'g)'���(2Nk�$���t�k�g��ι羒N�>Bx����uH!�OXi�l��$�:d�I;@2���ϼ����Кt�Xv�=g�!�S�z�5ݐ����I�>C��$6�`(Mr���yy�
S�<I�r��`މB��WD�̫��qK����eHG��)b��]���zL�,Ս�)���֕�s�k��y�\�E$g}{�}�$�&'�I�`e���v���Xb@���=Bw:���
�1�:��!�˿u��=���2v��H=RM�O��N�I<`,�@S_Y!s�Y2z�����������n�;�礇I���r���d�|�$�!;C���I���=O8�:���@Ξzf��Ͼ��o��ğ0� q����a݁ēl�ǶM2v�6�M3��XOXi�I�<O>�}}���!�t>`,<�=d3VC�O�z�i�L�q��C���'id���w�^��{�7���P�a�,��=j�G�C�O�=I6ɳ�MO��ON����g��Ϸ���C�}i'�����'!�P��CE�ē�5Ւ���V�N<�>��7����~s�M�I$�ChOFN� v�l�P��!�tj�|�Ϭ�hh�C�'>��}�|��{�>:a���a5�l�����<I2v�Y=I=`,&�<N$X̡4�y�z��������L=����q��^��a�!�<d�$8�Y'l;@5�$�%L�'����fp���g�Ԋ��r�;
���!�Q:i�ړ��ضϗ$zQ;>��6�
y2S)l|����%�? "��[��9��!��hv�.��uHa�'���T!�
23hx0����� _y�k�{��$�I���ā��C�^2J���!���!Ć��=I8�Rx�P��u�y���^s����'Li�����!�=H01��H0��<d�;OP�_X0vo���y�{���d��t�u@��gԓ�Z@>O�!�S����N��d4�b0��$5�J?}�z믽��l��t4�i&��K�$+'i&�,'�
�;Hq�ެ1 g�N������gں�����@�>��Ha�mz��̓N$��q��I�f�&��s�$;+�߽��}��>@��ިN�q��������I�	8�I�I�Yg������������'����@�Ր�f��u� vô��'�L'H��!����~������IXK@=C��Ԑ�`,Rm��M$P����$�ݒm�N�wu����Yι���{Bm ,�����OY�іۦ$���x�L���S�!�t�g!��cE�ک:��5=c-�<+)�-��a���&�jw>�$� �:�9aE�GR:`X�ؠ����?����I$�\�[�����r�~1�������N��XO�-�t������8�2}C�'�=������y�=�v�$�'��RL>����MD�yd6�8��XN0�<NP�����z��λ���6��Ad!��OS�!�'i�	�
��8�!��0K��0:��Ӟ��}��|�ІӦ
@�,����2O����>Bx���XO7Bq4����H^�����+w�_{��|�t�x�S�,'0� q �Bb@�P<d�x�C���(��N�}�w�uמ� �O�	���~��I�5�HY�1�I�:��|��,���B�S�Cć}���_u�s�<�
0��@>`,!�HyԲt��=��I�Y2��{`i>Bju|`
����������)��}��d�0�$�d���'���&?'^�!L��	Ğ�gW~��:�x�C��&����8�w�>B�|�t2OP=d�I6�z���>Mk>}���o�|�{�8�H�=Hq�@��́��`(��ۼ��_�uߟo�9�=�]:��
�(U�E �D�J�d��U��"�l����`>����ߢ�
���3�3n�ߞo�oκ�� �!`M�Ӄ�\���yN�F���82l掇�K���}a]Mވ��?�y�%u�b��L�A�<�����YF ���YC��B���/{�M�H����R�ʷ)�x�����kޏ�XZ��Ҟ�"�m'҈nT$nȮ�tm��)֬G����R�ٞ�qza=sv�x�����CZ*5��.:3v'�7i��(�2�5<�ۯ�lz�km���S�{w!�b����ggX�S� #�W�0�o��Д�vލ����e��cR�A\#���Ժ��@ ���#���@"��R�g;��u���{�'K��W�����)�CJ�k$���w���$Q��nk��x:.�L%���N�'�r�❽�\�h���tޫ��3��+�*\��D���ײ$�T���n��>��E��}6�$�yt�T8o�k��^k>鯗"�̮��Ao�Z�	�D�{]U�
tG�Y|�L��Ս�h�\�O[��#�K��>��K u�-��[��%u�1��c�?��Α�g����H|�+��]�O�o`����8-L�p���Q���$�E�DRAdPdA���X$� ��B(�,XE ������QUUDb)�u��ߜ����t[W����t�jW���n�?<�y����%=�ypys����O鏠w@�a���o�T��7�ڑ��s{F�wz\f�ē�fz�9s�e��wofm!Ǥ���m���*�j'IR+�CZ:J͌��ގ��pG�exx�9yK��P<�|�ޗ�}�j��l�:�&�~�V�-���;ܘC*ȫ%���#�X�m��ѻ9�����O�byP�����[#�}(:vL5{88n�t��__!��N�ڹV1��+���Zo��<��
�]�%;���c;x�d\��P��n�VS05�2;1woU�5��W+Wa͋r�hx4P6����g��~�1�%���M��N����Y#N�S2Ԣ��bؕ�D�rk�;���|����T6^c���t�4ڹ�~�W5�\��g�/��`h���a�1,U���H���a���ގ�)CC��SF�o
U���\�9�DCis�6/��ʄ� '(�0%��"�;1�}��h��LƷ�8k��W �� �'��=u}��ʺUgwn�֥�<s��SzS�^�D'�h�K�upi�$�E��ѫz���
����Κ�U�����Mko�ԒI)$�I$�I$vg���e\�Usv��:�n-z�vDoO����r�n����Zr�]Xre�+M9W�u�n���Zq;7
��ܮ�Z�^֙��\�:���\���IB����=���6��s��K�t�{���Ԓ��C^�8�֎6��y��;�<��,2�r9nNr�����7ur�Z�'tVXĽo����ȷ���}%��4C���uk�l顑�\.���M�Y�E�Nɨ7��T���N�ϐɜ�hG���,EՐp]�����<��f���T��#�%_K�zg8`��QT�w�������Ȋ��\���$�Z�y%��������A �b ��L�C�c�
֬ثU6���i�4�1X)(Ԭ�B�Ta�c26?&e�YhVbfRLaի�AR*¡P�X.��Z���vɎ0��	�t���c&�*V��dDX(Q��:e`b�3Xc1�M[;d��P��
K�{�	�!���o�U�ݗ'L=�Jx&��&�BV��F31��Z�����m�߿�~Y�W�y���(9?gS�s���*�r�խww��4�ɾŊ��؀_O��]&��sγ��j����'x�s]9�D,k;T�gb�1V6|j�p8��WXs����1�P���sr�ǈ�S��!nxz�*����1eZ�d��r?wT�����x��va<��n������}�c��H|oqjM����SXs΍{+�A�a�ų~ �r�=�w���T.����GP�՛��G�z|8|<��C<�e������p����s�J�������%?���hZ:f3�������J�w�6lW@9.�q{&	�.*+�{v\�HN3�$�LZ��x'�����|������Nvl|���l˨{ְ�2+��� tuY�Ou��D�!ŵ�+�z��v��8���[/����1�a��h�{�ȝ9����z��'��<��9o'�wy=zM�Ck�#�R|�E;��ѫ�a�gz����>�[�Y��}O�v�Q�z��m�U�o4$
����d�N�=|5�.��ii[��ˈX�R��A싴�W+���<<=5����*���Ϯb�a}u���SiiIq�e��f��%�^[J)EmH�C%-S��f��r+�Lp"��:ň<��=:��_}+��|(��{
	噉gUCat���=KGo���wS&ڗ����r�-�SMvڀ�eKN-���|��!'�+��U)g4ɎEMc����8��)[8���aC�?���/ӛd{��4���b�R�ڔW6�,����� �o֭���T�Z�-���:�1�ߦ��jD�wx���:��"s�}\�_w����v�����G��v����^C��w��˰N�}�x�D�	!C�ri�=��И���6�^\��<��Pd��{DV1�l�K��,���|�4�%02lh��Ϊ�ƕ���jW&�j.ݕy���Z]�6⧵������b�-��;8O��537�ܽ���{���y�c�v�ez��'_*m>�����9X��N�Is]�Q��U,��F� O,�Z4q��Ω�_��+uua��	*��K��ػ������ޝc'�QK:����Un��0G|8�s!d�?��O^ߖbF%uk���,̃|��{��P��CmT��SS/Öׁ�3г��\�����.��~�"�m\�@�v��x��+C��L�m��1�|�����k�Pfp�����j|9��:�I�63v�i[��L/i�s��� ������{��z��әeV����Ru��^�]	���ϩ��"%��z�kp֋���B��꾵��䣜ɝsu�h�k9S�Ҭ۹\w2f���伡��e�v)Y����]�����{�Q�X��ɩ57�
�Ƅ�A��ڲ�f�o0��
��j[]��KET���n��ݼ����ϐ��	��!���E�_8�zcs+vÃy&����Ч/Fmا%��du�9�^Q0Ҷ�$��w��V�s�	򚄷i�s�Ǭ��7�{5�����\wi�Q�Dӣ}x#<M�F�	ȸ������|y�m>neА��I���S��~:Mw�VF��Su��	��zYG��n_�e�E��5)���z�擶��� ���]�Φ�����Á�t"�U���M��"/�_a�X���y�ǯ��ӉĨ_\�鮁yOt(lEݾ��)�l5�4�ܧ4�fK��>��xu�ho/��#(s�yq���׆W"�C�˰?!^�4�{{��[�B�D�U�h����B�g�ʤ�S��b���ߞ�ܝ�K+iy�L��:}+��܅��C1g��tk[�ԨH4�޴�A��N�=f�9��Tu����:�Q��AH[în:�aiT�g�Z��3�g�&����oqƌ�5��{�j��NGՀ�������-8����n��R����T�g�S���ss�+�=-�pՏ_E��_tO��t*V�_;��s����̓�	b��E��V�����?`ܠ�
;S+�&���-���F��LM�}s�]�7��`�'�B���fY�������qm��Vb�\�Vf�Y�5j���tcD��S��q=8��^C��^ �m{�6��,�ux;��x�y|�]��BE�^��X�-���=��+wO�s�|@n;�;������ꪭ]~���;߄>�6�6�ْ6��C2������*��,X�*�އtګ
����+�	s${�1h�w� 9��}��UAܤܼ�p:]1�!�n�ٛc��w6]h�ѮwN��=N种�
_u��i�s{���K-�Sol�#g�K��	�flqh�
��{ ����|j���<,z�?az�9��)Qk[�Y1�&�,q��w5���5��S������!��)�/��q�w*n��̨r��_٫��o_s��������81~@U��*�fV�?l������h��w�N��˧�=�����8��.�[Aw\8���~���W6�j5A�_�4h��K�dyBAg���"b6��^�uܖ�@��7A���]�4�[��7\�b�dF# 7EK�����"��U����c�'E@x���t�L�xR�^t'3=L��t��ѭ�|�������C��Ṕ�M��	���G�C�-�=��=z�c���Z��9K��t�u�˫N�[N^$���VU��Le�N���SJVu_r��9�BH�F�������V���2Q�N�^�B��\��������4�d�uq���Q@��l�WN��]�������w��펺�a�r���j�t�����+b�R��b��V�y)N̮�q~zfX�x��t�
�ϡ�m^ʀ��� P-������t�Z�9�'Hr��i���;�t5|�+�;w+Ab�v� �r|p�1S�Pa���,ӥ۸��ԑ��r�\�*�3�J�+(�4�º����]5��ە�����p�v'j���Ն�g]���p��Ȏ"1�ʶ�s�c7�Or�Im�ܒI$�;K�R{x�� ��;50w��V�-(;�Y���/�9���3V���]��,u;�����}�@݉��f+���g-WO�I�F��&nn�،���i_6Q����-p�D��(��x�Is��X�J �c=[��lpy5�+#�f�.��Bo݉�)qV�N�29Ӧ��ي��/AwK�o��hs]=dOw[Fc�W���� ����. hi�+�A�헊�U�}Ǔg#�Ec�W�7�Ԗ9z9F2��A���g�H�ݣ�M�㬑H.$d�ph��s�*��ZӬdh��r�1��:S�qGR�Y��I$Q�$�Zݿ��QD>f��P`T(�T��b���1�˓���+
�IRWHi����_i�>ՎQaP��L��ȸ�����6��CT��ZAe`c�Tr� Y��*C`ɗ2��6�Y���Y^&.֥ո6!hl�~e_39Z��wװPqr��r)�����4�����5�Ǒ���H��xu{�-�=,���B��ќ��F+����nzC�N�˵{� ���yR�J�s��Y�B�i��_n���V3����fϳ��Y/4q]ȅ��k�go�cm_�����l�����j!���l�s������i�}�֪8tgDy9C|~��k*v���刪x����aYr��=�ʧ�����A��b�H�t^t��BMD�@�G�u��!��㦐H����NLY\yVŚ�aK�Ә����ӝ�� xNU��4����i�݅�q���r���1���[Q�����(AL?8���C^�:Y�=���z�6c����\�	���ҭk��K��!�jr^��z��k��c�sͦ�{Ӄ;Fw����۳;+�~^P�����g�F%�o_�����T�e[�K4xȘz��|O�@��zyt�R@��gN=~Θ;t|��藰jR��b�b�t�k����M쨞(F�������!֝OD���R�~D�����{#��WQS<ܮ��f<k�=f���}�}��<���S�Ϻ�45�v^U��	�$�r��I�Rq����Ó�5�YX�µ���,4����]S���}�A%è����ҷC^���3a�������0õv~�y�V5G:�U�(���7b�be�{�Zɬ[�Kj��1��[�����ZL'����qnv��RE�۴D��dy�gxT��
cz�$=*z!�~�U����� �7o�D�g;���qٗ���N���Χ*��yI���[��'��4�Ǜ���C;=N���������W���m?Z�y��W���![7�X��OMK.x�3�Z��$�uqn���Y�TZ�ˇ��
�eL�)�K)�ak���=w\�f��+	��[S��|���W~p1����%����^߰���3�O���<��|�����zi9eV�G�ic�f��}^��К��~jb�u�9��c1�ν�^������F����}���4p]�в����7G���5}R�U�G�Ԯ�;o!���s�����YPs��@�]���B�>���9������9<?Q��!��F7Z*�����R1���h�c�1�"�_9]֟;
��=�ە��`6����f��o�Q��
��@�0����R���6�dL:]�$G*�rb��P��*7f��٤�E��<��{r�NЉ�.@�)]�Z�VĊ۵wӧ5���W�ԫl�~�Ȕ�G�S�zg���|�&�\|Zg|�{�gϰ�*���,$X�+��u{N��-��w�y�W����ƅ�M�l�͜��)N���pڇ4U�Kh�����yH�O�~����$���\��Iϼ�fɘ_z-���Sw��o;P��E��r-�uv��t����6��Z;o��_9P����\�s�+ݘ�杻��n�V�ݡp�S�W���*���b�f���x�J��Gf����8�[�D.Q��5���p�:�xbݫ12��B��o���[��7�t�U+��pK�>^�T9Quv�f�&.!UvClF�XQ�L̕ƋT�{L}�u^0�U�$u|�����(j�9Z��&�.N>M����1��F�y�S���o�2����G���j��r(����69o�"��T�V���ˡ�ar�휱�/nw�tϹ�}B{b��>�sa�Z��K����Z1���s���D\���.:pɂ�5�0�`pʁEMռ�ė
<h�9�G��l3�b�:�Kq�z�ۚ%��6��{:p���#�慢����K�jx�g�x���T��Ǐ���P����x��T�"&(��E�R�g`r�R&]UҘ�U|�MGe�:�-���$>��[i�l��-���M�.Ȧ9��;�*�[.�.Ռ�J76�J��=�w��"O�>�1���M�,��3:m�ƚ�D�.�Q����b`zv`�˥�_2�:Qd�����id���Hڏa	��-�pϔ)��qğ43dq�q]�wY��V�JQ&}P)��7�%�-���в�#ۤ��"r�{r�L�l�ː̇�2�$-�\n�//d���)�
<�3FΡ�4`�`�x?F�]��Dnu�Wa��
�u���n}�H,�2?:XP�f͛���vs)�>CE�⍮�'�=~y\�$d#[�At3�(�^��z{��V>)f�6�-�g��V�K
�6��t�����q���u�k�'t��e���+�m[��R儮�%��U_}������GW�<Dӑ�d2G31�9�sVP���ϰP!�IФJ�(��]��O����7��>s|x�]�#��t(��o�K�P��ީ����}>'��(���y�9V��ǿmG�Ξ��W{�u�K�u�|H�n�
ԆD���Ok��%�z|bH��OlE+uu�(@��U]�m�}�I"�����^��!�>g"uX��X�8t���-@'6�j��hF2D���6��iWA�;�p;"�$=�}8�v�r�ӓf�����i��(�v�$�TV%��V��{n��Sk��W��mh�|�mڢ뙓I�9ـ�ÈC�u�T��&�]ea�홱qg��Hl��T�����j��Y�Q����ȃ�Ӌ%w^��n���c���߷�Soi������C�H�{K�g���a����*z}�j�1����%��<D�رp8�Jx��3pT��YV��}���ĸ-��2DI��} ^m'm�c���S8�H�I�-�>1R2�;E�[ӎ�x�!8d,�%ƒ��IEC̩A���6YޏC��A�6 a.9�~�=$�1=ʼ�����sƝ>��Mjv���)��}x��:۽�;i�6�q5�}*=a���B1������(��ۧ����>d\}�J��zGdcjý��n�=66��9h��BlSUf���{Ҷ�=6��E�gP�K˰9�۔���c��D6ʸs�zEz�ї�����U�5�Cכ��Ũ�ޥ̃PID�\����F�]o8^ꃸ-��-�w�cm�ReGZ�u"��b��Kx9.{2�B��Z'�q�����f���FՁ�b� �~�����רe����V��Ȳ���M+�E�v��GXϞ֐����3ru�=�Q�7($�(sJ�l\yH<�P$p�%gE7D�w
|\��c$4]*�VqJ/�7�ǝnT�kEYՇ-˽��W
�i1�Ev�y�P�9؍�BͪM����9V=���RI$�I$�I$�H�!���[�q�S�k���W �S&�gn\�y%��BH0S�n+�ò.r��d9��h�\���	�]ӐI��x��]h����*.��s5� �^ʹ�-8��P"��j�@w�E��mRD�#g��DyYeoǫV1�z�=4���6B������̫�`��q	�B�W+����j�!���v̚�=�ѫ���� �Uo"J͎�r�O$����Wr�ʅ0���l5�8!���N�缵��.�� �8����(���"a�!�Q��Ӛ�u�>깺��o��J�wo�wk��ۼwz�K�T?�" *B��f#|���$�jں���JR*&[�ӎ%Ʊ.���ְ�f[J���+4�Z�Y���i�4�a+4�ȫ��8� T:I���-cl4��<�z�X'H^�V)-�5�H)��RIYY+3W��!P�㈤�L����GT�ՅE�P+Un[kL��11�^��VVZe�%Ld�jeՏ�"�����8#����fJ����ɿt݁^�G;g������ɹ�zc�L\�NY�p�nFD
�*4�%���w���Pq�p��'L���A�"�	��\�<ja]֮}�Y.<�iY��Q�YÁ\ѲQ�,dfr�Nl���2�=>4M����껳��״�9�u�ܭ��8�l�)��'����P���"�֔���ս�C�L�J,T��p0(ER�el����S�rxD"L����� [�"�iw��#��{�������/N*swǚ�9�۱����gO��y�링]|4TB]�����G�1ep}�M��kV�D\Y`���@��9FD�2xЗ"��]u!����$}
���=���U4�报GՉ#�����ٓ��)<��dt`ܛhښ��|Ը��r�k�sy�����Bߌ���n޹�?��.�ڼT�k����~�o���5#n=��AGxt����0�d��z�Y�����S���1�nG��08���M�Uӫţ�D� ���8H�E,끒T��|R����˸WG��8p�(�@捒�Yf�#�/����f�Py�x�FlzΗ�t�1P(�y����mFA��#�J,�����>X=`
;1]a2�m�<S_u��2�}$��s`q�|2��9��l�Ǣ�p��3P+��� �1����k�r�;{�+e�v�#M�]L�l�ː��>�-�7������o�З�k�P�4lWof�݆��z:O�
�G�!�B�R���(b�gSý.�;��
����4��F��H"N죉�!������WY��~�6b��%��!�8{L�έ}����,�P�D����6�V;��vOm��z�ۃ�,}4RA1R�ҽ��
��]�?~L9�=����M���0�b�yE��a����s�(�j󷤍0ENHJ4��"E)VF8
c���*��Kz�4� �� ���.4�d[�2}�WG%=�붯�hAĚ:YH>�H}(�F�1K5�of�{�n���}d�Y,�:�I���\X�i��%�����}#2F1s:Yd2�:#F�ٶ��*,�p�"�`�F���gK��iks}���h�z���<6�
{���	��a�A^�!�͖3���0qdL�����*M�u�#�/h	<�3!��}�gsm��B�?tz�?R�@,���8���vNP��7i�Q��M(�U���-P�F�p�w.�z��թ�0����炂�L����ˮ�<���0)��y�w#Ƚ�F�6b��:dU�C=Pf{4�{HL��-���-��>}N�T�:vi��gfn�̿\Q�������i��&�\d��V��W<`uR��'*p�����yS�ɶ�>�D�DnG��1�(\Z�:Q뀰|ND��5��p�o�Y����e
��D8�����J����MP����Ƿ�v���C��9x2��O��9G�u�>g3�&+�����#�h`�7,���(Q��+�P�t\(-�0fۧش�E��\�q>��D�EG&��>��j�qs�᳤J�讁�.4�p��Ȓ�?���e�����e�?�zeH�6F�"�g:	�M�}Ӽ4ۮvOq�vʉqǍ2f`i�4�EB�X�Qb Q܀ɨ����2��TǤ{wB9�=͈'A�:Q$MԋՎ�\PP�J�c��З�}J��ng��,�3*E�dWA<A���	�n�,p�NCi��2B$���,��sEȾ���"��p��((�%Ԣ����Z;��a�Iy��Щf�jt�9���{��Et2���<����v$���&��p�>Er��o�����t�x�J�+�����⬥\h��<cI����[[�^���4Ί��@��c����ݻ�����n�����{~-�_�Y�x������ Z�4�B�׉LЋ]I��%>Ӕ���\���a�l���x��Y�Z�U�#Y�����(d�i��,�1���֍Z�(����y8d"Ƹ$m���"i�̜���g
B�IgM�t(�0"=�a'�cD��y���w^��J��g�����<7��|��ȹ�-�cJp6jx�;q}��(�8ڃ��}S�y�����X�o�;}�J���s�w%J#.)�*�z���K���D�32 �vF�p,�"sy_>��̎$�,��ѳ�:W@}L�H�<��$Jq- 
z���ǀ�ܹ˵y6n�Uڑ^��,n�8���kNr��xw����'%�5�)�����WF��r��y�������pi�m��ӽs����7dY��G�!6�3��xi͏l�inw3�)�>�&�#{h�pd�8�K���no&j󱸯A����p�~qdm��"hB#a�ir���p�B ��!��0�_������Ds���p,�L� ˊ�@]n�x��/!��[&��(7/�R�2>��8D��L�>%G;�Q�PN�qw�dagkg�YF�.���_u��0}�q�9ҡ*�#)VF8
Dq�"�+���)���*0,�D�%F�h\}��O�(�Nb�e��k����v�_oc�Z��ͧ���Os2�OU� *��[i�X)r0@�a��.��r�/�W�U��1�����Wnr�Ô㒖x�O9TǳW�b���X��0��Q'�C��I���D*�u�zSylveԚ+O����)�w���; +�#��n��E�Dm�nbH��Ƕd<��L���q��ˬ����7�|x�����̵;a!���4�O��Q# Y�f��QN*Ԃg`R(�'5#���W(j�\�iŸ�u��QD>�eԼ���M=��+`Q��#M�}�"��M\I���o�z&�N�Ǡ��j0���S��K��4�f�4��ӳ&�
�p�h�xE
��������&�c���0H`}���1oP�!����jm��1�k+jj���6�����Dv^��uZH�s�~���3JI����ö�:NT��S�P��=�*z}b�e嶤\�4��̌��8�j4��6B�&f�\��>�t�dq�R	����I�MH9҇<ܕ�R܆;$	�
}g+�0�H�r ��-�'s��b�]�mƑ� A�!F��y�ѳ�nS1��{M�G:�2yǡ��8F�".Ф��kx��%��,���x�8d��ٍ#H#]��{��p�#r�$�mt�]�!�QS��)WY}�ݞaA0|\YɈ"���Y��T7"<�mY�����Q��!�:@u��G�u��Lh_`������ca�q@�V��I� Pz���p��t)`,�Tu~���Si��9\$�(6�qJw7����ګ���U���A��t�Gĸ��q��D	��Ag	� �z\���Y(�y�u((�n0�
*�g�C�-J�����ǋ���f�?�A���/�Yk���.U%DԲ2�@�P1DX�2�}}�UŲ��Y7z�fK��E�Ҋ Z�"�4��=k#�>�X�ةl��F�8�u�à�D�kj�f4�n���+ An��v4�T�<I[$tC��gmj���0�"r4�����z,D�&{
���h�

W��C9P�I���O`�m�n�^�	��˖hGHwj�l�=цH��h�{��g��Q��u�UƑ�t�vDW�M�3m�����Z(=�{f0ὕt��<�Vڈ;d��\�׊B�e����ޢ,e�yW�0ُ)q��!k76\���M��'cGe����,���Z �
��GB��M콈v��i��ML@���+�W���ﶶu�̤֠�U�T*���ɍDo+pLyJ�V�V�on�7��:���c��i-0�*8%Y��v���8N�]^��܁��z����=t���S�h���bŚ:�C7P��0?�J��(���ݷnN��)�������&
?>�Aȍ���@q����h�j����I^��eI�ZM���dX��wN�!5=Հ®K�9$�I$�I$�I$he�5�,����'f���Y�n�X���E5��M]��=w�qRw�� V˚�&%u�������v�d(�uѢ@GU�v��B�#>V��$�
�Y��fo`�i�YJ�:M�U���=�@�Zu�/��0�=�Cv\/F�4�{s��;Ic#˙LU�w�	_�E�V]H�mM{]a���M6�kC�g}f�qЮ�z�ߵsݸ��ھ!,�T5�	���.��y�������Ӿ+b�v\��:�@n �mͼ��)��@ڼ�	�(����U�'�J枞7:	3��p��k�p���NٌE���k(�e�I,I$�} �$ނI*
)�z�L�S@��1���,���V��b6�)1P<�hA���a�[,�=�ƶ�YR��-�:)Q��z��a4������8cE�&$r¶�%ḏ@Q�:zzg�sZFbI�P4�J�铉j�5m2�SY1��j�T1��+��\��&��R�M'�o}o�gw�{o���m�Q5�)tD\��֬��n9����^���qW7����Y����G@��E�6c���o�#v�j�Z,���ټ
'o3f.�����;y��=8���|�cS6VD�!ta��8F1� 3���[Wʟ#��"T��2FlzΕ��l��U��;�#LN��"�6##����r� Q��v�N��z�i���.��w�z��x�,Snl��_�5)c�����>���[����P��&]O
�����BK�t�Q����X W�]i���e�a��>/v"F2Gl��F͘P ��7w�������Ȓ/#���t��$>�t�Zl+�
��d�OZ|�g`{\�n���+4�3�h��a�y.�[��q��
�Z3Q5��g�Ņ�f.�;>���.�np��4����]�lQ�,ؤ>�����c����CQſyw�8.p����r�!�0���/�>�HE���r8��.x�P0��B�X&j�Z<`�JfY�H�r܄l�w�œsT������t�p8�|�ۀ�	g���2�{M�R�]D�#�=d�y(�@�`̣��l�E�T2�xW�x��u.�L����^x3omٲ�G�(�p�`�x���4�"j�s9�':>��E�e@-Ϩ��xB:Gr�$�ZI��õ	��#�MtqN*Ԃdl�b63�4�u��lm��$�z����g�h�he�H��׷�֍�P�$��Am03�G$+�u�kƑ��nV���!���;�\��~�?8'ޓ�۞]�L���y���"��g%��{"|��y�x����3Q&��!.����B6�H��9,��965k�z���V�{��(����F�@s�&n ��WE�j�!n�Us}������
Q�ȩ��O�b�i�sR�lEq�\�'�`)2f 25�����(�q��ۛ�ɫV��u,�=9��wO�Ö������L{�{�K+:�n`Q�������c�32�
�7�SGٞ�U�K{�0Xw\̊ځ]՛l^>ދ�R�Kw�R��J=
�L�#bd=���:wY�Ǧ��j��5���]�@e�7�[�N-�K_�{��I�-Rr5�K���oj���r�L�W�H�S�*�f������U�֯��O����۴�����c#�͈��('"EA���3�
�Ef��3b��1'X�Q$
:zb�r3���ķ"nr�kJ�a9(f#�Y�\aڧB�3썼�8�W7qy��<s���u���<�*\�v>Y5����g*$�p6T�9�u(�����j3.6u<���?l"��/.l�>��&G@���eH�u��j���H��DL@dR��*dѫ���{\:��׎��3��8�C$ˁr4��b��V��ms����C>�Q�d�T�h��\�#�՛���zTus{_0m<N�3)ok�b�f'K=�����z0:��MN��;Niշѱ��β��kd����:x�o{ϟ�:��J�Ω�ע�6�,v��^���zev���4`�%3�ۤ����ҵ���φS&c�I�|��Ǖ�w*p�r�D"8�@�B����(��I�ק���
���Q�8jZ��qyYmw���#�!�p6�Y���O��*��R�y�.�\�r �^G}���� P��ΖM��z�]b��:`��'��p���$L�Τ�ț�]�\���g"$�:x��=G����[�C����. �"�:h(G�*�`q���謤��$�m�G��@rx��Z�.8��������bP��U��0E����n>�(�nZ��f��[�L��Q(t�ϧCԖ:��R6���l�Y�]a%k� k*��^@����2�z)�ؓ5�Q��%��W5��0�������3P�7 #EB�n����#H��d2v(�"K=�{Qٛ΃4t���
����S���pHk�a�R��o��2�&EO�W/`3�Y�騳~gL�͋u| �����v᝸
B�YG�ys.�W<]� �0�p�302�E�G�8��aY2����������6`��p�����G3�C˨��힦d���w�w{swn{N(�Si�)M�]�7��v�4Q݀�tqu}�͒^B$�o<�'�}9�J�V\E8�#xDѭ������}�6�J����)C4L��L�VTsZ�_+Jځ�K{�/�C��������|��S\�<�;v�OYfd�÷oƮ�DIÄ2�&�ql#��YN�\xX�@����k��h�oѱɚ�6��*r�x�E�gP4�H�$�|�lW@�*4�)��U��mm����<k,"0���#����½�]
mf]N�"x�`�q��J)G��F�6`��a�޼����v�kr*FO5G�#O�b�r��ֵz6�)�:i���l�n�tX �5��u;׭�;�rp[�AF�"�R�F)F��1nb�-����F��b i�|ȃ�0\Z�5^�\͒��÷:���K��ѽa,�ՐYjދ���w_�i��tNbW|02����.L఻���?U�O�{�ܧ��S��f�C'`t@���E��{+{���(̩|A�ʬ�����)x
�(�7�`/[�qg��R2���6(B��
����\x�Z-3���_�槌��L�]2}�a�iĔ�Vjv�(�:\��jdv.�G��u��>�z$�G. nE%"j�ty�PPY5�}�\ɥ����@��.b�r2�K2.q�y6��:�Q	p�E�a�(����2�[�(=Y\�;R!�e�1r4���z4��b�wu�GI�"�;'��{q o�W�K7멂UӹWK��17�]'���sE�$�Π�cz'|]�:��bK *p*������vh�3�{�4�����O�9ՠI�F��wOՙ�˹:��6|ȠE(Q�6[�Xޒx�����}Y-�c�}�9(�@���L@�H�d�Ǵbi��]l���2�D�q'I,��QDP&���Ǽ�htЖc�>��|���vK��Ƈ>պ���@���M�\xA��#!��s�Ѻ�kiv貉<}�audFF�"�'��Q��S]�"`��v�~����7��S�W��=£��d�$�׵螞'�:�5r:a��9M�v���j=gL�>��#J#v��",Ɛ�������>��`a���=�ʐ �=�8̮�&��՝s܌IBF$�̓�R-�ʰ�{:���Yx�]^i�s����9Ad��pl�OP�k�{&�L�r�����c��훧��;��/�����u�; U�gE*�y�VxY�nW��;��e>�
߷�y���+h�6����vJ3�Z��w���H�"�V�5��P��0m@�8�zU�"��S�>a�F�6R�Et�{f�S�>]`lUv�}٤��FD�:��܎3S"\Y5�Վ�;{ T�
4�UO�c�g Y�6e9�>�SC5�	�S��ޡ�s�I���@�\>pؤ��5(�,Ҏ#�Q�
ȹ[�a��6 ��fv�}�4������+a�!k�FlV�(��%��gT�OF�ɓ[���M$TER���[�蝫���ug�d��9��.cY��ftzbXWS'�՟bv�/�����ww��E��4oM`}�27hE5pC��:�]�Ɋ�|�KXql��h��Nt8�Z�v�Ar�!\R+p�zy8��h��J�,u+�f�M��l�-����9R���Tr��7-+�)�����d�����@��r�eө��m�0�+�}]�VD8�[}8�uIH]�i�˰q����^���rTbˠ���,�����/�'*J�{�)_ �$���ZL��N@kVL+_�&�f�b�[:RȬ�lY�v�,��&�˫BH9h���^�{�����$�I$�I$�e�)��A<ҟv�S/{kY�&�j�|dSŐ]r����us�K��ej���V�1����4�eY����D�f���z�d�t����#��	8�����&��M�n��5��oE���yc�4��C�ܺ�&s�g�6VR�L�
�u31[�H�;�5DҾ1o.��u�J.�L⩋9.V�������R�6��N�#&�ӳr�䨣�ʩ
�C�R�C��U��j��ж#)۵C�	�vp��s�d�9[�D�;T��f�1l�6�Ej��=��w�	��[X�K�rL'����Ht��:�'Nff��ĒI,��||I$�0�2�F�z�b�8��$R�J�VhVc%DAb�������)]�@DģL�-b�kFԵ��̑�o*�6meee�*��m�34�,�آ�5v�SE��2�ݠ�FV
9Jέ����֭˂V������T*Ԣɦ��eD`�Q2��*$X�+���	 �NFL���b*�U"��.�f���������{;)jf���(�^���p4�>:|�f��B\#�s�M)v")\9�o��0��31�8v`Y�H�!��Y��_uKz�V�ٓ�Et{�8Z��`G�8�=�m�q�-�GqB�O���Iw�idF5ipۂ\��'O8�0-��d�<E�>�گ9vtQə��"�A�����D����,w<��s؝
-D��O�L���
s�(�u%Ż\�Y�@>P"�0�,��r$�H&�]�޽�f�0B&2̐r4���PVxS�F����|���F�4+�9��yQ�A��Q1�M�kX�^|�(1v9�^��ȋ�����TJUk����N���of�cf���&�d,΂�l�c3~���o�_�SF�z�}�ENO5G�#�Ŝ����j9<>���M��֮�DS@_X�tz�*���w I^�1N*6A�/dR�&�b�F)F�Y�y;����F����I#H}
"N(�
"l�Ҭ�]��:l�lO�ٚ�2gѲ: dƂ�����c��=�a����������֐�$<�ž�wu]Q���롹Gk�]c�b��dS�]%?�O��I�aH��$�1�O(�(}2d��<mK[�@d*�����#mD�(�`Ⴎ��,�#���7!�s�_O�Ǭ8Zb;�����]o��X�6���ʩy�CW��^w�Y�������c�����7�Z�3V�5ʋ	�ָ�Z�ڜ������x:v�!>�O���Y�!TΖope�$߽^���9�ystㅽ��:v��w�n���Ä���Ƒ"�ID���D�l}�;dW�=u�si��{E� �߶$��x�B!� B8F���j�Ǻbn*2|��QGj(�s�ޒdt{�;��g�d�c����h�3)st�B���b�7�U�/������v��������t�J�(��4\��S-c�.���6rT٣B 9Sŭa�D�ts�ڳn�ۺ�ɚ(,++�p(d3��n�2k3�)�yԉ<Ig�1wCB���6��Kw�׹^�߰hG�6�ggc�l��h��1|��<�oVL���9�`���3�����j6d�p(N�G�qV<����6��Q���3w�x�>���FX�d�K��+.DL3�9H�����O�@fb4�@�����	\��r�gbt������.4���9D@�*�eD[�26k۲,���N*`3=g��L� A{D�cLM�����,��fx�e�7�9�wv(�u�C�-I���eK�^�l�er gA#���>���唣*�.�>{E�Hn�؃
8y�2:	����3IX)��Ǖ롯��Gް�c'��"n6��J��O�V@�D�+\�&�q�H�cp�7n�z*	ɆP!"Aî9��̌�3S!��v�aziӚ��9q�'��	�n�����k/���|iي�~��RԒR���[�N���,���ڮo��ߧ/�SPE�.F�"k����#H�v��d�Q��~����j�$���/Lp\ vg������/uk�q�Fvq��O�W+`3��z{��,w�/��Q�5WW�`�{(�	�"�7w��5w.W�a$q�,�`�����BlQ�������<l����N	�ڣ�w�x�w�[���4�f��>�}Ӈ64�P8�|�#ex��)�.Zi�ǣ��.��8פ�,�^�{�
՝�;`�04�GTA�v�ځSD��[ښ��y�;�&J=3<x�/��Mt�B9�đ.C&+��/�����A��]%��VU�sd��G�cTu�3w�\,9J��=Ƙ�7��KI_|������xޞ��1�d=�7�8�ҏ��.�	����Y�`�C�i'HkaF��#�[�$���Zӆ	y ��>�N�>��k$)1Ʈvb��j�kd[ɺ�WCp/����Q���j$8�����h�:xȬ�5�4����9���Q�D2.�mf����3G�VM�2*$��9/h�yK2�k���F�ͳ<�5 ϱH���.�-�x��Ҷ=#N2�k^�5�oHgJ��dqs�!t(��̓״�si�"
�<x�D+�#v0ك�3���L����Kn�gN�"�rR4�ElN���8Y��WU4�0�+���B��2eAy��]S�A���R0n��q#��7y
��t�46ԫ�͒��Ͷ�A	��L��v���R�s,�U��G7��

��ۯ6�)�W� �V�IE���(������q�]e�B���������h��xS:1�.Z�/e&/MO]=��v>>�s��8eup��<�M�n�]s^�P���}Ĝ>���6`C���u57!�[�C�Bp2 "\-���<}g�����&��&ݦym��j�����wT��7�x^�����|$��.��2Q�n捐�8��D��nWfd���s�#7ǰAB�`vlZѷ<>i��;P#��5�y>GN�$s��& 	q�\�C���x'�����_f,�v#W�� ZT�2���ٙύ����ɦ��P���^��ʎ��U�X�ZM�_�ٝ����K<d��#*�Qf�4�B"2�YY��]�8�}��D�r�=��G�T�0튛4IbQ}{Y��Z{2Y�q�W����C�Y��n0ʼ�M4����e:���=u[R�����E8أ��s�,�!DA�r�K�U�,��[C ��q;�RP8���v�5�~k���j�}˓5����u�#'7:j�ǣO6òD	b�*̴��7�t��Cs��>��T�3�Ǐ��|0�X����;oX���Z��%J,����)@D�:D��N:չf"$��nMǤ\q�����;V��y�)�䄂�9��v,�|���[1�x�n�S+�U�)���<fĉ�VF�mr�lu�ks�
Q宓F�<�'8�;��`�l�����u@ߠl��q�C5�
(��Q5��N���JI�D�uF"k�HUFQD��^D\����20��Q��"͒p��^�8�.\]S���P0��$�U(��Ǝ���dP��GʋQ#/�rŝ#j�"P�$�G��c�1^�j����,��OlE�0+~����`v)�8爘��xjɶZ�Z���7`�㎊�dP��j0�
d.�͞z��y�"a9��q�D���"�	��F�p��bʖ�Z�+�uǑY��o��Lh�������n@T��_@]�O�2�>��cJ�Ј!��u7�JO �`�[n�]��EVy��N�j�T�e��fj�U�p�
�t(on--r�y��r!�w\P5�5F��W�?1������gG�¹�uvmY�F���������#����F�F�\�A�訓����*�Y���$��F�@N	��G�*`Z��6`A�;���U�S��wA#K���2'��Mt�B8U[�*l����0e\�u��D��53�:Q��[������tC,�I����ȑ�P�E�_j��!��ΓuI��Rf=1�[�T�����VȰ�JP8Q�Ly�������=�{EA0;��|<LbnoJǩ`YS�R�xd��`�1\��~�A{C�zͩ����y�s*W�h���o�XZƘ���.�eX:�j����q�b�v��5��L�¢�"���b�
��U���U����KY8����19g@���qŻK��b�e�d��!w�@T���cw�4��b.�ӗ��_��L	�p����=&��wu�f��/�=�Bt"ȧ1��� ��MRj�aVx�� �!R��a���u0�D��5��đ�	��mV|�D��BU�8�{Y�s��iPN	��*�]wtM$��0�=�U����6][�wW�'y���1ϐD�`[Ưe3�N^�<ov�c�ot��@u[�Y��j�s�B�I$�I$�I$���Z�.Q����P��|��� �N�"��)7�$=����/����o��LQ�,^�5���Y��.D~B�p�OkI�3��M^��༓�v9��囸o�x4�3r�rS�j�3OE�JV
��6�,K��}�oac��\�ʫƃd˹��<�Q8�y�1*(��n�kU�&���n�Ya��Rap'%tof��F�m�l��ݐ&����S�Wʘ<F���4�����ά�ǀ�eh#wiB!�:Ț�:�����Vkmo>8p�fG���nj��8sؚ�fō)���"�t��DɜC�B�I�b�s�$Y$�X�I$�� �H'ē���$�j5J(���RҪ(�2ӻA����mb��Յ�i3,PQ�c�����-c)A���+5l�kUJR�jѭ�J�,���c��D�K�Lm��*7Y0T�1�n\�(�[�g���(�*�i[eEEDSM2���z���[e���fd+0�h���ޮ[��ڈ�����
彴QǬ��Z+����Q�EV+[�c�8c2�Eam4��:��C���8�)����2��r(�U(�4�Rvˍ���Z�;��i�9q];3�J���(�K���1k������f��ӑ�Mu��t�_^���w�L���x�o�g~�kދ�I\�"/��m�I�#5p�f��5�8��&��r��ҩ�d=<{���{�I[fGR<�7(s�����x��v�zZ�g^��ee��{�HS��ܜZ^o��G�o]�Rm��V+�+�D{�9�Z^��̧G��w^y��͓�r�^ੴՐ�S2䩙�a5B�u��\�">˵�υwQp�����&�ˎ��
���v���jE"���f���k�I�&��vv��_�6�^K�#��<��K���+eT��:-C�!�e�<��DOg�[���������hI�s�-y_L+.g������b���^����;x�C[C��6|Vr�9����@�P"�E�3wWdН���b,�\kq<z�Hk\�б�&�\������Gf�=Ձ=���0�ul-^����f��Z�����:{����f�.�5�wr��'�*)68�f�H�f��/8�.aa�|�f�l�si�o)T�t��1�E�K�:['-��*t�㯷?<�s��e����a���d;�Ͷ��zc���/�q����*�k4��z{��_cy�ш����U��1j��H��Q��/���w`:]�4t<��p�nͰ���KP����=����k޺l[۝ɬm���H��=��+c����k�^%�i^1n����'vs�.�!b��E�!�W����y�#S�ܞ���^�W3rA3�GJ�����C�u��V���q��[�t��7�IT���ro^!!5�:��?^�#9��~���8v�8��
/������y�Ui�3f��F���I��Z�P�ϫe�����
iM~�'�5�l�Zfܤ��5��I~�_��}C4����ޣhm�f��?g�z��:�r�!g.?n�)����]���y/���|֩��0b&�7��^5���t�}�ҳ>�d^\H�k9�m]�;�P���OSN�RC�ҫ.Up����Y���e�*��Zg���#���v4:<p��<�\4
���J��r׏\�1--�����[6y���Uz��&��׃Ғ��I���[C*jz�F'PKlm���>�ͳ��ݖ���̧(ѽi�![Y�shD��4��N�y��1�Cm���'��&���ü�{��������Y�旂��q�is	Gݪ"���ko�l��Y�Jl�J>���/A�C��͜uڛ�k�g|�(��ޗ�+����<|��tv��S�^\ȼQ���([��VV9���&]� $8J`�,�s^�x*�uM�%��zrܧ*�'Gf���6!�2�.�/�� ���;s#^�Ǜ���N�Aj��n�O9/�f�֎��D�c�હ��r�Nt{��,���Ǌ�W�<8M�Y͡���z绛�Z�l�Pj'��ע�vr���\��x�,d]�E�[��h�㻃"�ֽ��!Y5'2�Y�컼��'�:�����{��W�~�r���-�����l#�ٱAo\%��yH���Ss|�F��������&1d���aډe�w�
��]eQ��^A��UَD�gw��WV�$���;��~KL����ᚒO�^�Q�Ug�N+>�vu+`���u��t|Г!�V&��
>��.筤�<>���l��k�v`����s�ͨOO����������w���n��|��$x���V]>Y6d���7�,n��1�� U����s�7�>�	��U����=1]������(��]���`*o��ok>��(�:FcK*V�� b��v�������1����H�0kG=��h�價c/�YU0�E�M��q���t��aU�w�S8]��{�1�nw"fZ�R��9%��L�\�|�齵�Y���z��PO�.�޵.(�s }�s�W��Q�{.^�\԰g��������شՓ��^��|�Ѣ���^n��Y�P�Ef=��Ӂ�'C���|���͑ElcW��Z��2��xR�Ɏ��{�+̔��%9ו�9zc$@�d�8��bi�謃�g�<����,����j�۪��a��.�s�F׷.a�њ�Nzd��y�bŘ�f:��4���w���ʍ��8q9 ��|4�G
: X�X�ܣ�8[���o�5(��XșF��4��rTˣ�)E��`IZu��MN��z8lz[]��k�)î��:��fg#!�S�J�F�ުF k��xW^\g6w��ˣ^�~��R�Se.F���)�	sty��
��c���5]��=�||�=.��ʚ��ӎs���R�z�A���)��ժ�-ݭN˧藨t�^��-����O	~�Hף�d_G�4�
���OS����(�R�Ntz� �~�Z�^F���ezBݤv��ź]�[��(��ۅ�K*�Q+54k:��M� �j3���Q46:�,%r�߻������o���Z�:�i��5��=�v�+����2�Ef�v�$���N�\�{,�:r����S{զ�^�i�E�����V�/z�{kȹ;/�S�ĖQ��YWL:C&�b����� �%�81M�vMzm�S�0�j�����M˅8�����r{ԅm1'Z��&*�+���Oz5BxÞb�i;�&4WkNQ�5�y�F[��&^�S���T�@;���G�y�,KiKk+�Z��y�y�MkB�f�2�N���n��I�^�z�ʽk{� �o���C�Oaf<Ε��ӡX���D�WϬ��:j]ɳ��tS(s[�R������\�ޜm���ؤ4z�[��՚����d��s\�s�'y�N:��\pr�wטq���ۤ����њ:a�Om�*�n�oH:����D����P�L�Z�xΕ��M�.f�ְ��GK�RZ�i[��	���E�z�j�E)d��]rn����P��*}t{s��!:�r�eJ�ӽ�E���O���7�aݻ�8��,�>��!�f�ʯ`&e͂���OB{m]�m`YS�� Srp��mϫ��3WU�Q9�I$�I$�I$�F��
�t����\�A)WcD�.�$Wr&������wH�2���YK3j)�Z4Qh������\�dg)�lm�6K�BcB��2�/f\��`仮ͨ$�Ν�d�~W�<�;Pa�CY�9P�/r�X��՘���{V7�L�}RH%ա�_;��!(�Xq,.Ժ͕�'!��ei��II��Jb��ao ;���v�v,딿������b�w5�H� ���$tM!�z6���)���o�.�
�K[����+a��Q=]sr��yjޥ����J�L)[��C٪�P2PN�vovFF��SK+T�}WNU�i%�.iCX���V��W)b���\T�Ԩ��̨��2�UW���Ab�T���*�q���F*�EC��f"�e�6�"�KX�S�pJ,�,QFE��1%Tju��K���B�3dU1��ZYZ�6�eJ�m��`�U6ܲ�"V�C�ň`�2��aN��Z�TkKjPEcQ`��n7-0��[h�j[J��n�EWM頢��j����T���`��VF��r���EAE�b���Y��׽�����~��N���C��9s��[�jB��8����x���/?3D*�Tea>H�#L ���}�(V�}���S�<3+�1����8��{�Yp���sd�<c�2g��ұe�1��Up��Ζ�A+�v5)����ہ	b�V&��bI�����M�g�+\��p�\3\�ˤ�v��1����f�\7�.��[{t�M^ܾ���jә��~�y��������-��O_{ג��p�2�'�f��W���W!y���	��ks�����-:�w��в�+�����Ä�%7Ĝ��t���{މ'X�3մ3�B8\~����Qt�t>x�Rey�H�vOM���8y�ܘ���B����DN�����55w�ҁ{^�{oYk����u��1���Vt���ÿ���zN�B�c��=�Kn�C���o�q���d7�j)Zڷ)F�L�X.>�k~��Һɼ��w���Y����x���]��u�Q���6z�������{��|��%*�p�l�P��;6��HhԘ]	t�2�ف�8s�
R�Q�3LI�ƭI�����R��@�������@Λw��{�oem��v);���2��a�tG�<晉���*^Z�%��K��%X�\���5�~����|n�F$�y�1��hf������j�ϑt����dЭ�u�Tޅe��4]���o��$q����v}ǆY�-�3H������Oj�K��}��%��f/b�J���I��8E�sxFpȖ�l�MK}k��o�O9����ueg�%�����L�<Y����t�Y���EJCccb���۷.��|5r�$�wL��q3.B�U�r1���(�;[ϦPA~�;���O�`k�z����=Y4�zZ�l)��0���9��Q���l�K�۳��׋��ғ�70�*a�O����#��iݯ�1�\+��k^��}S�'Bu9��=�sY�w�����[��9
2}%fp�:��z�^fsl�{G={L�t�[����-�|�;����>+�贇�a���zs�{���L���p+��0�R�V�Dr�{�o�<ˀq�g�b�֮ �(���P��B����A!���Vnr��fd?��m�OUЇߧW��D�tw�ݼ�j�7�oB�N�8�ڳ�������>���t�yLO�1ݪ֬yr�q:�+������/e��3�q��$8�Y�g�:�tָ�8�E>�VA�y��v/3�Ş����]��Z��������(H!�J�XC�znWK�c��㲺>�t�3�<�|�{����iU��T<WT-<��yF��;��I�
�34��u~����nSˌ�MD8b�V��mV$L`7���*ny5$s�x���!���S�52�[����q^�7`��))�T�?U�zl���9�|�E)��T�΁�?�ۣ�������O�8��٧�d�z*m%㼷$���E#vGk��n%������)��M�t����:�tw��:���^��<=Q�t�9�B��'��qNW�g����mՋLv�à��դ��ww4�o��}�� h�9jj{C]��X����ϴЯz��t)6�Wn*+/My�N1�+9�$*���*E�+��.���\��+H���/��R��.U�������=�F`��wrRz3Ow���8T2aو.Z&�|r�#{�xw��
�D�s��jU��N&�b�PK��U�*4�뵗����@��vު��1��T٤��T��K�kK��X�s��b��LL���2r�Z��
���������9�gA�q�{���,�m���|粵�R��^e�P�!s��~ܪ�sϵ���.�	hUN�[)u����[s4�E�1�7=*�tSj<�(-E�Mawg�uw�!��͋��O��b���r���:9d�a]�]z�P�z+]���n��PA9,��/�Ȧ7����~���?�,OD�U��/6.��J�����Ou�N�LU������.�Ȅ�O��-��-N��)_�l�MJ�>�T.k
;}=5׽o�Яxz`A{Y=��R��G���t�r/bcH��+�eN.���:<V�y�K&8�Sk����HΊ��u��I=�F��9��O���x���m�(����'��TOA�+8=5����KpՑ�����^�ZK��:�8�w#�8�{Y�t��>D��b��B�}�*��E,��7{����]���N@q��rU�#q|���ϔ'���p��@���{]�/%{��S��v��7
��f?��{w��f�;��-�l2i��봝3+�^����R�S塑E�~�r�T���੽�e����6��n&O,wj��y1����t�^��J9�g���*"��F3o���p���f1��[��e���U ��"����h����2��}Y ��Dp�J�W��Nt���z�ݵ�b]쮽�7��+=Kl9�w?�ՙ�$��H��~ԠΆ0���y(�����z�ym9��=��	���43s/�Q�+4Msǭ`�1&�q�}.���\A�qQ�*��w5�Ni�E�;ܒ{\�Y@j���Iӏ�`�,0�w�lR�o����y=ѫS�/m�n����a<��{�U�����#����.�Dt��s�D��f�蠦nw6�Ws�/��C36���~��V�GDɷ_�G����f����P�>��_��[�g�^3&�U�K�[uP�!�hҲ�$,�շ�'��^���`���$�ͪ��1ON�l��z�߫6S��Xb�7
��Z����.H�f��������pX�4�[�J�V�}r�e,6*S�`�P�����R&�!sNդ{v���w6s�r��[�Q|(�k��_]�@��ȷ/�u�K����*5��u��ͨ���Xݘ�*7!���]n���,�MK��ӱ��ǿ]��Oh��X�T��nH{�hz4�(f�9��i�]�Ap�fGi���4��
V�����u��6�u�8gM��)5gp�(��-^�n���}M��ՌMI�I$�I$�I$�G���*�wj��f����/:,f��޴t�)Yba���z�,En=��U�6k�x����7��X]\*æZ���Lø7e�&����tB�\f�[�%�T8�]:�lK��о+8se��2��I��<����0u:���-̢��0��ח�I&�W����L핎"`,���́3�+O��f��#G6�-�@�çU�+=h��㙊����gvm�A��4C� ����Vr��v�F�����v�pjKcp1'I��7��ʾ�é"}Cs��,�\#�@dS���r�>;u�)�Ι'<A�aqڳ�\�CrO�u;����ua��W,�3��c�+W�1�"��`�PU�Q�w�bGT
5驊�FU���HP�J�Y�\n%�%T��aX)����Qb���%b��k([EF,+"�VEJ�[* �R6��LA���V��R/�XY�
�B��TP�S���k"����@R��P�T
,դS(Ъ�T�C
�-�"� �8��őH
�U���1 � �M��1��O%|�����;ڹ�8�u��{6��������������V��P�D{ǡ��枻�/8,2ج�9�0�([[x�Z�=4�#m��}�W�9J�]Ў˧֜�r�hp�ż.����jk]�*/f���\�Us�/{d��p���p�gN*J�����R����vkX��J�Mu��:ޕ��K��W�h�maw{ٹ�؉�4��[[�CnJ�f�c.���d��E\�ɗ�J�h�Ӣ��fXY�2��X"U��Cc���{�����w�s8=K7���QB���=	1{s�أ�RM���O/<���Ԯ�\����H��^�;�k}[uh2�Ś�d�W����]����%Ph�`H�U��اK'P^,�bȱ"�u�ex��h� �λ������:�E�y��"p�W\7��X��<�G�����jN���kh�b��_>�{^�r���Ew>�s�����y�b���ت��T�S|��{8$���'�d��-�-�:�X���X5��w!�ͮ�T��;>�_���]3�h7yvֻ]�������Qj��OPV4��;!r�V���;]vC8�X^6b���_YnH�O�>�@Fk������g3е](4��:v�uת�[:�''�[�;2{e�q�2�5���ǽ��u	��./�b�Ra>y�ٸ�{�-�mҫ��8�3��+�G�ǫ�vv�x���9^ϞM[����9�M�{�ߛ�RXo�wL�N�)����f�E�.$7��M�_���uj`�z��-��u���͋��v�mON�w��'Y�gth�8�M����7#��ā/��3Uq�^z���ˋ��֮�U�[�Cn��(�����6������.l�{�3I��7q�����0�SI��d��[/]�0A�`�׺C���
�:z�g�6���tc��~��Q?���  �^mr���HN��eq�Z��.}v�� |�^3����5�H4��:5pb�����������=�©k���M��p�C��q��Ū.zG��z?{�Ht�OzѡMJk�q�wHa|�6A�S�5�*�c�!̽N���N�Spoʅ��h�ך՟R���y�/YVu�]�w�9�W�D:����Q�te'���ԗo�w+F+U~��K�o]��{�&�wzC|~)R����:�=�w��g��}�R1�ة�<\v�A�1q|���M1v � �O�����9�I����ն3'8�O������Ǯ6^7Z�1��{�VE䵻Z�jn���M=ws�<u*b�:�8Gԋ�?S�&=�]���Z�U<���KNu޽d����U�)���͊�����P��' ��z�s�}b��v�W!�l�Э�D�s�wr$�Bh��PT;ZV5^�G%fvpC\�*E��������]����_R�R���;w�'''����?X���>����3�Vi%ނw�+�C�9{���Jr���{��ޓ���JD}���1�~�{��ןc����TC�=~Qf�ޖ�O}V��
�q^�eѫ׻���h[ =�u>�HU�!6O���ۃZw"�yømn�s��)$�R���i���hӽ�� �Vry�n�X{��H�4����?(�uA�J[�騸����;UzNtUՠR��i�wԂ� �8�wk:*�'�.1���'a��rћ�)���ʽ��ԓ��Ak�g��o�M+��S��ԔW��I<��^��]V޼�S��2�������c�����<b�n�tv������k�b�q��Ψ���O��*v�i�]�}�>SM�f>)�~�z�����:#̍��5�e-d�q��B>�t=�~�o��e$�차T������O�7�
�C5�R�W��`<v7�.WX�.���.����r��}��L�ԇc��\�"�D[+5g�,t�1����Wr
�3L�0�aԜ�4�ee@yݑ&��h^��[�q~�ԛ<;h��oy\ը
og~8/�F���w�Fbk�k�KI5f�+6��|�P�;�X�;�������mZ�:�]��`|)�W��%5Ko��]Ej�P=kǉ�m��\�y�LU��V��Pb�����X��_zʙ�Y���_��$~V5#�|hW�����ʭz����2��Zq6�v�]�{u�����=�]P����<U��7r�K\������h�;�J����Ҿ��2�͉�g�>��Y�H�\�NT���/U ʍp���l+�:�s����<V����xߦ�ࣴwZ�ٹj'�2��<�[�~03��=���"�Ǳ�Oiu|,J3/�H^+وy<Փ���[|�&3joZS%�Ui�x�yL�ұ������z7.aB��"Ҏ?L���L$A'9;����C\�օ*�{w!����+6z�~��%��7mN�U1�ؘu�����'�7�tT<sG
[1�5%�]����{N�}�M�
�z��9��U�f噠W��~ �hZ���]xf���fN�n�r&&|cI�JAf���iX�Cl��vÛ�{��"u{&V�k^yQO�����R}���ˠ�-����1f�N�L�^<�gZ����̩啳!�x��OhT���>�Y�W��L���B��j�<��+}S�a�0�x�U4���G�z(v�2��[������,�T��o�z#1�Dd'�˅3yo�Eh�.�J���\u�����X�t��䃈e8+WU�	;��G��������~�z�7{�C���?hC�����AT���@DE��>(����(9 ""����HF���,�0�\iyrK��������ِ�B�P@TP%h��"*�G�Z؋zٽ���vXX=а?&��Ho�K�i5QB�d��E��`"/yMSW�_ޛ���<�І�f0�(Bo[�*�n(�	����(o�ɟp)I��廓�	R��4�al������t���\�����(���� 
"��oD�(�8&��.�&���?�?;�������?�U:���:Pq�:}H����O}����@4YJ��E**X�z�q��4/�M����A&B{
+)��rR�EoV�n9@�<c	��ơ�xB����A��Q��Q̓l�J��g���B�U���d�$��t�@�Y���Sl��nG�87	��Z�.4������/#$�CsxqCh=7�6�ø��R���:��6�쉽֥���`�4<C�� P����8�*�h��n#E�eP�Jj/8	��$5��^\?k�Ш��`	��S���7Pt�Xv��� ׈��ү&����=���� ����,	��_8���Y�É�X1
���
�htb%Ҋ]�AQ*h�� ������d����vO��4�.>AK%ME�<���TD[��6V$Hs�I�������Lh�lQl87������'�w��(�����Uo��ڄ����X�ŨI������""��:�c��hާ0",�'��/�V׎�v��ixi3�i�9��?�k�T���Iu|Nx@�6� ��|�x'��{�b�|wiLR��P����l� ���( q��D�'`"-��PLZ��z!�A�4��3biv���'ov���b��5Hz�P�� TΚQ ���ݑ���L��ÚM=�f5L#0�i5]�� DE�G@�ĵ�n	]��T5S��1!ۀP���5mY�D�B���v%����6�Л 0Q�+����w�(
sO'�����p�(���y��ڐo�H^�=4��e�Aqb½�C���z��F '�Ġ�-�\�.�p�!��