BZh91AY&SY��U,�.߀`p���"� ����bM��     �    7�$�R�"�ڕ	UD�����$ �*�IH�%D�a��"�)P44	R���TH��T������B��}��)�*�T�m�QR��U)J��RJ(R�	!$ ��AJ�%HB���D�
�#�@j��̔(D�� u@�ڥ�m�p #v��Ud�-�U�m)L��[֡"R�"��H*P��҈��HJ���)%Ki�k*���'�G��   y篮6ڦ�Qlm�V�5�\�ִ�pwv�*�I����j�۱�p��ێ�uukVtu��T�j�ꣳ�Ӫ�mE�닰��
���%)E���  �{��U&�H�n�@�*��Ω4�TS�n��R�q��u�J��ʊ!$����4�[�}�ԉ*]�{á�UV<�ޮ�IJ��¨���R��I�$*��@ ���%UU)�ʽ�J
��K�u��U+������*�V<ô4�PwS9T��)7K�����֪W�)E��j��M�:j�l��/��$*T�	AR��"�UT����  n]�j�WM_wg�Ҕ%@�Яsԧ��ҕws�N�QT[��z U)]�;Ӯ��Lu_{�UR��{'W�z��SΕ�yD�:i^�=ޯfP��츀�RR]d��� ��o�� �޾R�������n�R�[�w���ڔ-�vox=*B�8�{ﾔ���TV�^��)J�/�+�m��u�U��JM�n˝-����u�u	%@T�J�Wlo}�@ �}�@�Vƹ�wt�!�7N^�P�W���T����jR����Y�V�Wm\:�<
US�F��:�F�6;�B�ݱ\��M��ZR�]R�*P "��+Xǟ) ��i� �u;�%Z.�pU)]!�����x=���8����c��UP�p tM�u ���j��풍�)!$�TJ��{  ������:\� Qw-��9�qJ�껊
c�� 
��m�t ��wN�w$h1J�H ��JO�4  w��AJ��;� ή����:UFj.� 9� ��:� �rY�֌����%H%5lH� �y�H  � 64 ���*� s����:�е��r�� Ѻ���wTr1J�� �       50T�J00` &LS���% M    SɐRUO�@ &�&   �1MJT2����d�d	��$�J"* 2     ���ԢD�&�5=D�O(2=FG�����?����_��
K��Z?�sʻ���w(����ͼ�����|���*�9����>U!~�*������K��K������B��UPj��m��/��������D|O���������58ٓ��a�Uƕ�e\h�S��c�,�Ƨ8�\h�'�jq���n53G�2q��N4q���h�f�8��G8��S�N1q��8՘���S�.2q��N58��.2q��j�.4�4q���jq�Ǝ2q���K58�Ƨ�h�'���b�Vj����h�S�N4���K�N4���Y��N1q�Ɨ�iq��N1q��N4���j�N2�2q��\d��d�1ƙ��N4q��\jq��+��5fN2q��N2q���d�G�N4q�8�Ǝ4q���i�W�.5.4q���q��Ǝ4q��d�*�5\j�e\h�4q�8Í8�f�2�2q��+�8��h�&n0�'8�Ƨ�aƧ8��58�f�j��4q��8�Ǝ2q���h�S��b�ƪ�G8��d�'8�f8��S��jq��N1q�Ƨq��Ƨ�d��jq�Ɨ�N58�Ǝ58��N58�Ƨ�U�8�Ƨ���8ÍN58�b�N58��N0��\jq�Ƨ����N2�2q�Ƨ�d�*�2�W8�Ƨ8��'8��'�k4���8��'�h�����Uq���jq��S�d�S�'�d�'W8�Ǝ0�3���8��N4q�8�a�8��N0�5W8�4�Íd�G�d�Uq��f�8��N58��N4p�d8�CYd5�8�G�k�Y��N2q��N2q��N5q���jq��\jq�Ƨ�jq�c�N2q��\b���.1q����jq�Ƨ��Ƨ1q��N0�S�\b�\k58��S�iq��.58��S�\ig�iq���1q�Ɨ����,����ƪ�'�b�K���b�'q��\d�G�՘�S���+�+�e\ef�4q�ƪ�G8Ì���2�8��a�N5W�Vj�E�G.0�G8��L��N0�'q�8��W�UƎ2q��8��N0�5Y�q��j�2q��8Ì8ҸÍl�ƪ�G8Ś�ʸÍa�fN2q�8�\h�2�4rh�4q����Qdɵ��a����q�8��3'q��U�K����ef�j�0��U�+�Uq�ȫ�J�0eGG��K�UW4Uq�W��4G���ƈ� �T���Ҫ��q�8�eGI��%W�)Ʃ8ԧ��K4+���R8�')�	Ɗq��h�2��q����.2��b�'�j�58�Ƨ8��S�N6d�*�Uq��b�'�h�G���j�4q���j�2q���2̫�8�q��%�j�5Y�8�Ǝ4q��8�\d�'8�̸ÍaƎ4q�8��e\h��+���2xР�B�
a?���U��T���9m_�U�J�u
s�n�{���Zt�� �dȲ���Qٕn&KDTwX�
�@��r�ؼ"n`����+kn��O����4@JP�sL+8�cf���ִ���-JW)Im'�V��5��I�P�j*�jCd(��ӂ �/	��je�R�Ӧj1�76oRZ[ۀi�-^ى�Kf"w���r�=�Ce��M���3I˧�ϳQ/Z�Z��#�z��x-[�az�n쑷r����t��-/ڶ��
z�(�%F�b�1���!�4��G�.n6�։rX֫/f-���*����iK!Rm7wA�-:�對WH�V^�&�m�^V�e�;�<-��D �R��F�Hj=R�S	�u���H�%kz�P�T%ѱ7m�؎�t"�7�0eX�n������u��z���GB�pc�
�ei��3!R���6�P8��bB����m
Ӯ�`�E���"�q����B7�Tʺ�,n�*����N��"��٭��b7�kp�h"���SQdf�P��V������F-��C�Kk��+�Y�YZ��s%��N�2]+��3)k׳�2�MV&��ʻ%H� �H�ڗhc�7�-c&�Cr�Ջ���wA�yP<t.��6�1��ؘefm݂+F�i�\���;"�Sh`�
��w���D�S;��\��-*�6�+�b^�Y.���˷tm�OC�F N�Iv���Q�.S��j�����I̒y�,��&U̓�[Vm��$�mӻr�J��і��v�bu�9Jh���u�0����r�z���x�A�(��Nm�xۆ��Vnǆ0wcYN�6��
у)�KD��\7�:[���F�RǴL�XC��깆�fWlHU�/00��7�h$h�ݺNҺ��&�e���	Z����kIׯFR.Յ��q�r�.U͠R�+.�`�.�ɉ�&��uvܡf\seT�mIp��F��U)d�����e�uJh)Lљ�yA]��EpJӣr)QJ�[K��a�LK.ҿ�m�P�]6�)-�Ka��%)L�Wr'�v�<���F6襶�f��Yd, DV�ւ�Tk���� �	g���6K�e�RVQ�U(���ƶڽ���1�&�h�-6A��.�����sn9���r� ���	��3]e`���1"ƠV�	�yOf+U�[W�0�«I�����F�>��L��n�B��!�)�����'�/%�.�wr]�*��wɋ(�o6
ǀ��x���6R:���`�w��ض��(��H�r��`V�i��L�ڭ�0�Ѹ��m�]IOk(�j��k4����ԭL��*Җ����Z�T�i6��L�'2�7��
��t
�_��5�x#q7�vn�@M��P��Q���_ � R�ԋwE��B�;*�w�*solݫtpH�n�CXṸ�I�����W {Oe	+����Z��j�Q�j�d�`k��5���^ʎ&#������ͭNY�Vݒ�Dm���ˏT�[��`v�U��L��*!���.:4�H��u�k#�
�"jhW��qL{�1�f������/]]�j��٬ʡO��q� ��h�35=9e����z-L�n�5����fy[���)Ѩ/]�O$6R���WO<�	Niˣ/�e;B�v2j����j*��+Mm��z�y��R�Tܔ�sL-�8
�5��k^�$T�0�$�F���P�	��b��7WA\��E�pa*���JX2����w�N��|�V\a�FЬ�x�8����J�-OhXP����6�3�2i3wd��(Uwm�xfV}i�J<�^�f@� d��%r�	P�f��.kQ�u�۫�w�5�!�����[�u�C���Y�N1o�e��7!;ᤫ!��0fJ��^R7KMI���H�:ΔCد��=Z�Ջwv�ֳ�j �͹��3�G���ad���pB�U��2�V6nneŬ6����),6I3}�YXs-(�a
��6v�Xn�S���ě��d�.7iV�ؒ��6H*��e�ȱ�ݬ�Wu�lU&�t�0bsuMHsa5�T���bjU+m�[�o��%*G�q��2R�_;�H'CD[X�\Se]�T�N�f�EiR�KP�w�kiȋ����	i۴33C��sVi2��0�ꄁޒqk�mU�2��i��9�B4�{��$9�2��2�ވF+�n��P��,^�-�v���h%.��55i�4��6�u�BT�Y����n�E���r�QP�ܽImgΰ��ˇv�=YZ-�r�s]?@�I�F�ڴ!�U�[v.2��t욺�eͺ�J3���Aj\����36��2:с�E�����P뻲�kb�Jݵ�)Z�ҽk�D�5֌g�B���f�]�0�1(M�Eۧ���]��E�.uz�2�'���d�UO�����9��ٕ�q�iݝ6���YV��)d.T��2�kh�#R<h&��9Gk�y��AR=�@��Bn8m��3Uj1�Ya�Udܱ�ܬp�4��Yb�.십y-V�aj�ʊ������a�a�-Pݘ0<M�J��֥rT[����)�(�P8�aU#�3tE��n��z�hp;���Q��x�B��Nk2�)Du� Z��w>N�L;���A��]�)�MUP��%1=��n[�.y�zUu7$�ۨ3j�&�ͬ�m<�Z�*ꮹt�v�Ն&d�3��V,U:�-��MV��uZ++q��-D�;�,l�p��-�J���fT,`T��Ceme�--C�C#�XY���	�
&�	1A� ���qK��;Z�U1�۶yf�$B�*֏�
z�5�P=q�S����D�`��B�-��k(<-�z�ކ�įql��Y{�������e�F��f�X&�.-����l#R%�kҶ#�mkW��0+��E�ڼ���/[J
����sE�����a�uz�՘��Q9�jXA+2��Y��:���c��wEfi��)^����7� Nf��#=��X&��#������Cj�B�H)eX3.��������J�6F,�wS����d9gQ[�F�5�U�2�BY�[��eC�+C�#,���ɂݸ��t�ܬU����o�4��kxuU����A����B�����Fݺ������[V�hŧ���ר���t�ӌ�#.��[r��b��U�);�ͽ�y`�0HyV1	�+�H�יaF!�Dn��p[���QaV��l��w�6�A��Yۢc�ۘ��,�O��`ݦ��ވιC@b�����Q����Z����I���2�Qa�QC�?K����R�å���M�Y�֖,�h�B�ʼ��\q���iY����V�tF\(k2ָ@V�t^��Q�Wy���ֳBYɸ�EL�j�t63wq��Y��.ֶ�b�c�KY��	,�N�	��Y|��S�_D���wIW�b��y�^
�]�1��$�ިs.�:W� ���y�'��6Ya�m�	)R���krk`bɏ4B1Xa��u���F<�0��.����b����U1JS6�r�1;��aY��Q[pM��d�����溭b������(�Si��n��;�U�܇fE�,�eL5"�UW0I�CM���33F����i���iїK�i_�ǅCwh�2��6��"I1���Q�S�H�$/dd�X�^�k�H�onD����5b�X�	D�[��(�^Jf�Q�Yt����ѵ\z�;�*��ku����1Q�*�h��P S�������ٛ����B����潊b�4LSmض��l�U-�`be���L�0���T��8|in�hG*�ۣtˬA�[��ܥ6ҙ����Vl�a�M�u�Zȭ'��
ֆVՆ�d�մ��n�\�N�aݚK2c9��,�5ZՖ�Q��V��0T�k���ɮ����f��7�=�Lmi��:�(�41GU(T����ɶ��S�;�N�	VvSv�t.�Ȃ��l��6i^�o&�to�"��#/;o/R:Q�x��v*�y#�GiضY2�
UQԱ#V����Y�q��R)���(���xB��`��!�����rIM�F�U�1���ɕoX��P[��Ln�c{*��X�ص�[U�6�7NVU�ih���]�s�b�Y[f�a�qZ_h�V�C�h�nl�ܚ�H�5$k[�}z�Y�T�Ƀ ڳL����R�&᧵TK�x��TM�i�$=e�����X�����L��5��������x^�uZ��׆�	{ ��VI�B�/7�(ނ��@e�--��ilU�('�C�x���y�m9r)Ú]�8�-�t̽AҼ����Y2��]kd���M%���b�T�YhŖ���8�{.�ҤS�k&�ÉD&���V�6�������%�yc3'en��=X��Á�ۍ�]J�[sF�Z�ösk(�Ww���DF�۵)}�9ć.�փ��Q)FyF5��Lt�1T,���5Z�U��f$d	Ce�ؖ�h�x�K:�H�,�(#5=ȯ/n�k˱���+1+6E���a�ū��m��Y�I{�oK��^ʢpFőt�P�����CE�J��V(�w&�T���쭢�2�&�	��Hi�,���^�8l�L��-���1WA��Ui�	(ͨU2�����C���/��R�]�xi=�ӆ��rT��U,
T�8��9j���D��/�NȰh�4߅"19���������&fQ�wBM
��v�7����0M��.�6X5��HJH�PyvfE0-̀��j�9{�m]�eLv�c�-�F��OC�*u�r��R�ˤ�4\�sr\l�v�K��e�D�������m]�`���XF��Y5u��mM8Z+)�.i�y���8�Znb�A�Mڎנ��d�${r��6�q�=)��Kl�i�s0̔�dSe���*,��2��J�;,��F^ꆈ.�b�
�⬬�M�{����
��m�-���Q�r�=;�hP��4�[Wd�rbc���p�t���7t�8�@�i^�V��f)J��.���1y�B.����b���l,��0n�Zhж��Z͌�zۧi���2,��(�NG�������x�O�~q���'z`�zp�5xӥ�@ļkH���C��l�M���:i�c2Z��]��6�kڇ�ךE`�083(�J���O��r�}�[$MG��u�l�3�P��˳K�I��j�"���t�n��$���RN��
�.�(,C&-���,�w$��ob���D�MOt+

�Ri݊;��%���wV�i�D"F�6ol�v�V�Ǡ��khڏf��{��x$�*B�#)I��f�-�`�ǋviW�Qv�c��1�Z
2l~׈JR㠓�j�^�&��q�R�ʍ91�Z[�e��^�����tZ�l6�I9If�j��苍�*n��i�c(�@����Gm ]e^\�g .�N�����!#F���Wj裨l����y>t����:���vp��������F�KN�ݰ�M�f�����񚌸�iR�i��/�wT7 ̻u�[Ʋ����2�0�����j.�D�hi;V%/{��H**��1�V�Z��0G��nV�{�+y{HZ;#)Ϭ%E���5w�Ƣ�N=�+g��J��8�;{W���f�6,�6Z��"�ƱіO�@��;"��-T�����]^��LAeK6�~#	�)�=+�z�}yJ�ѻo*;�E�:i���oHP`�L�5�z]��;ƥj�*6��8'�.���؅�^�Mw��e�t��y�ƣvأ�Ov0�ה�.^�wِ7�������ne")�]���ע�L��Zb/2M6NX�]�f�Ǌ�h��9��[��S�3��o�l&��uV�8�fc�`s*P�2�d��k	���AF-2���a��3UCCj���Q�Iy~޻�Ǯ�]��-�fN8��h�4.�h��q�nE�N�6���b�
}��CJ3��jX*k�9�Ò�W�`�&���H�����R�����o�U��U��b�JJ��r���%�_e�6��N'eX=6��k"�ߙ{j�L��v���Ћ�!��j���o,���`ͫwk��ĝ�oy�A���]�6�@֣f�E�>`c�T���$H��r!u�Z/*���QɁkŐ�`��8�q���"j݇��E����
�0��F�zb�|	�����$6�ދ�W�]u}(���y#ޕ����b"u�1g5I���N�ҥT����;�s����@�a�7��(�&���m���ya<�8��$�.-3L6�ٓ����܊��XHԮ��/Ux�q�u���yf�p;���V{�<SU�3��ғP;Z&QL�9"Y��T��-|a���tq������˄Թ:�BXw��!ѱƔ�}�`,T���g�ܾ«�6��ȳ�R�̛�0�Zy�.}(�tN��p�{}̶��@8�t2'��1��t����
�%6#��֠N�D]ͽ�u�S�9��8�*ޓ��C\�PH�*���d�d�+�8��K�����ge\�-����qA�wT�Ŭ�*�|�M5x �q
�J��9.���+��3y�ب�y��wB�T�idDnE6F�Z(�c�*�^�j|o:���a�ϝI�Vtt'r��:��ե��=�Cq=���YY�H�9H�z�=���M�t�^���]�j	4ҭ�W���Ӝ�������� 1��,ǫ�if ��h�Ij��$6��j��0!����tκY�9>����nL�k'�$�JwB84a<y˹��)I��f�,�?��R���#Xj��}ki!b�X����Skc��c�J#t�����o+�j��\�&��J��[M<����˭�C���tsh�:��!qj놳�
g;ɸ0M��3n:Y���`�MJ�5U���������w��/�{м8�����_^f�������9�ÆMoN��)*VXK������%�邻�m�i���q�9��.�%�|���'Tע�&�m����
�#�{Ϩƶ������Gq���NI1�'��f��7���]K޼
e��QS�m$;�U�:�+Oh8���[��6T��*q�OT�:k��pfͮ':��wL�ݥ7�WWI���l�ó/�o�"�(�`���v�p�;xo��I����K��R�G�n8��7��r��-��T��-���nou�oN�fI����Wz�Fų� 5ꨒ���Gj&�i����ѕv�[���$f���b���hV1�v8>d�ރJn
u8�Gs��#=�_$t)�Ş�yH���f���gswü�ӟ7t͹ܝ��nl�)w 8���3���I�>C����B+���ȍ�y�Β�)̦;u�����.��k9۵Se��$7�r�@�%�ֶ��%���K����V=5��R�7��m7F!�����@���3���j	�9V�+BK�]�T���O��9:�㜨p#.7����uD��N���p^�JZ�9��Ջi�I��ʬ�d�z�Z0��z8 �����'�-���
���9����5�����T�'p0r	�1[ݎ�fcxվU0⥴uҹǚ�.h@�Wq	��W�*�_2��gg��.�w��uo�M��ֲé��/� F>����w;v��ʻy�{���jJl=?0q�k��,��g3�r�H��w���+S�@D��ZV[������=���e�C�yC�j��:�]��*@s;x���ln6���g�/>,��.��G���{�9]t��g7c�N�G�ٖr�UM�������q��Q��H�rUt�ǲ�4����Q��o_)6�Bk��9��i�����9ͧ�-�o��Љ[�Oi��C�N����l���I'jP���ٵ[��2-I�����J�N�a��3 ҋ�[�%E1��U�5^d�3�w)ڰ�v��ꍭ{��� �7�.wTv��gn�F�n�r���k����[���\����w;5bb���zp�5\k3��;��]B�
�Mk7u�35h�R�+�n�B�*Xv�"��8�<{:WX\�z�e�7��89`52+�T_rr�v%x�T{B�Q���{����Ui�k2�V�\GEM������6�ޘ�×s�򂺡�V��}�)����wiv�5�ٷ�����x<j��P����v%i�2���&��Y��7	r����?k�N-��sS�f6�`k-���F�ѳ���!�=�KΉ��)�
,`��׹�o����[��m=�AegU�W8��]�*'a����7�x��r�9wru]`�Lb�(�Ŧvm��9R��qSӞġ������r[�8Nu�G�:����[�R<y�/޽�v�w��j�a��;��s��ǡ��Ԣ�J��on>���*1b�q�4�Fu�g�O��締q�QB�ލcK��U�s�)$���<�N��of����[�s���`� ��;�M51��#L�u,[k>�+j|Wn�S��#}\u���TZ�Nn�I�|lC�X����o6�̇k�U���]���Os�q�NV��\�5ô\7ة`���*,�wRZ�ї�ӕv&U��-�N�ǙyƻeJ���Ĝ;����QU�;t�{!o�vcW��.ʚC�8��ŧG_ln�ؓ^�&�fN�MnU˥j]`0�f;E�&f�D6���eV.�Jܬ}�ٟX��g1,����t�}��� ��cg)���od|:t3)��'�)�p����Js��s[��f�`u����,ɖ'։7q�9��v9�Y���a�j��z�Ӻ����g�r�޴�d��u=k�X��ا�U�;�
|1`��30�5��o$�䭹�n�,/�֫�"�8&=�[/Zg�8(M෷�d�vNML2_}����@��W���F��θ�Q�̷#�5P�(=�r����j��}��Wj9Ö ��ok�tR�#�nVu��Ƕ4�}6��#�hC�9��$��S��fV�Y*�=Eԏ�y�[�a��Ļ����!"�7(K�؎͓����˱B�����Ū��aҝ�+��U:#�u�m!<�⥚���c
"��RYw:ԫh��gp���\/w�Ӽ�gu�	=%wi����
�}#�kU�ws1]s	/U�7o��Lx�>��<���K:`N����Kmp����U�E�����CR�y�]ݢ����	Ι}�:����a�<�UUv��'d��U��P��\��xo�dp�6cs�r:�;�-S���a>�6a�L��֐�A�3�*�H6��/n*�Ug���oE�4�6VU(�m�dnq�k�YU�D�hL�;���7������y�����L1�/4���v���i�ү;:q�lf���{K��۫�(1S�8�P��!��#	�M
0m��(���ȼ�fޜs
�e�C�X���+����q��ŗ��(i���ʽ�GYQ$�f�;�ꪧ�=���%4�Њ�C+����ʠm�p��p�OX���v즲�J��>�n�k+�cz��Y>tjS�>���\����u�x�9���Kfk��q�i������\���mR��0M��Ǽ�*�"+Eۊ���O9��էT���K�en���Ƌ�p�گ�bAcE�#��Y�]�}�8d]*ۅ���z[�S�̗�uZ�]��N�ˈ^�K���nƫ�+9Է085k���\�_p9�Ɨ�y-Mb�$�ݡ��5��%�q�fQ�=OZb�
FT�Y[%�����n�U6ڲ&��:�5��mف��Ʈf��r�삮�*AȤ;m�
xE�M��Շ��;[�I�i���%��E�����f�ۦ�q�u����T�4�M|�I��-mNʺX�!���r&��a��3���;���<z�0�B��y��֫�\۲v�G�G��H�m*s\�,�푘C�Ө�Z�hJ%`�YR؛M���y��v�R7��8z��ӅЋ����aj���c	ʬ�d�2wdt3�b颲��Y��iTC��t0l������]��їAZǖ�Y�bv=ǫ�p����n��Ƴi
����޸Y���;��Vk��:Lލ�صE,����v�����{Xu��ޣ�k�^����P�協�-�"t���2�Zy7m����y/*eu�U�{�a�&�<S*7���-�9ZSe�^T{�ں#0�C��s�L����5�:s�8	�u�p���@wxA������4%�xEe�+o��μW�7B��A[|7'
oK��Н���L����IZW	����n򴥏yT{~�_&�^X��w�#Rߐg
��.�5vom�f��ih��I�G
y������j�P�W�(S�k��ƎHet��4��Y̫e֭򖊷�<��O��N�
=��Km�H�{ YuO��P�W7��A�7�վw������p�f+ܙ|�xsxc�͠���!K9b�V�7�t���;J_u�N��1���<�}u�����Gyw�Q��^�w&��_[Ӷ���(iP�x��&b(%%��a��)u�L�+��_S����r3Rm8�����moFL�|+8��A�$���Ή����В̸���s�_
;�'cͮ�-#����&_U�17�%e�Sr����{���;��:��6�m�v���"&K;�&���W`0x�vu������Yk��l1lR�}�C_M!�.�{I�w։s��-Ǻ�`���iwG}�ɦ'a��(7���9��c�R����۹���N�	%&��M�u"U-��!}�ێ�c�h2XU]=c��z�r����aT�K�"��jP����<�oB�V,�6�MN�N�ʶee3V�KR��s��(��w{����ʯח~�eC�p�ސ�-I��z2DBZ�� �Wyۚ������b��&����Q��V�K�F��Ae��`��W|z2:
t�}diէ�f$N��&��ʆ:�0k��)�A�r�#���q\ۘ���
:���f5r�R����yA�=2�R��[�W��R��j��]*r�x��7�B�n�9c.�R{kۖ��Y*T��4���O�+����9���MA2����Hk���T�C��0�WgǷR��#%Z8s�}�^�0N�j>���2�`J�sqe���Zæ���ov�k��*U�V�n]�3ix�˩%�4���]t&�]f�Ġ�4�; ܀Ip�-W�H����7�&a|��)��wT��6n
��23�
�����͝����ƎU���b%�ׇ�����-n�]�|l͙(��6�h����`��Zr�c����1ݽ(���gh�MT�kz2�ά�/�K��2�˺!����d7��wDs2]���Yқ�,�zĴ�HW\e�lѳ�ub쫯�/�4�A�YrQ��[/�#�:y�r�UU�6�N!��t���6ｫ_uz���vt��{���7f�nU�<�2;8foh�4�j��˟ad�$se�κЏn�XG��T{z�d���"���6$��z^b��I�M������h��Y�d�(UM����G�S!�pڐ����T��HR�͡��u�͆��ڵ�z�9-�Y��*U۵W;�>��ð:k������m�a��Y�+s�V�"2��Y��Zx��#�Ci��ZFV؛�zԼ��!��fY�e��c4��Lv5F�����)�u步��w����6�ҕJ��t@'[�`�޷�͖*e)d�����q�z��]��<�W���N��|���'D�y�����N�*8+����b8�RoQ��n����6�e3Ŋ6��K�K�{c:�WH���ʕ�꬙Ժ�z�s
ki:{x���7_�Y�%E�0W��H��c���6�t�Vs��t��\��ogv\��d�:��/��L�n�Q3�j��>�G��:��֬��eX�秳V�ݮ�XKv�΢�Ͷ�%SI��ӎ�5۴7�;5�N�K7��ӯs���@�$Q��ㇲ��f��A%��ܾd�bj�Rö�,����F���en2�V݆ΊL�t�%��I��7�@��2e���;�c[��$.��� Ʈ_s��W��
���o�E�v3K�����o��Ɠ�շ�7���<�o�*��̳'N
�n�Tս��`1Z��m>i�j�)xc�r�ŧ%I�뼹���Pغ�J����C1�f�MY�͡�m��zp;�w�����B��z��4��.�oR��4=U{��N�ڜ�� `=z�q3@�Zkx��z ���,%�9t�Kt/���kH���x���w))�]%Zxo�4�	�4#[o:������7%�V�p��N���9Y��!v^���S�gzc��윗�f�j H�ѱV[DASVn�'غ4*N���l�%Z������]98����/~�k��� ��EM����n�8�O��*�P��*��B {e���r��@[���;��<`}� ����v��w���k���(�6�Vɉ�1���Q�7/��u\�T1��6��!�Z��tP��(���*��f��*�ϯ�N��ؾ4+f4���60'"��s�A�Y�=�iB!@�]�g�6]��"�d���X��iWm��]�������=<a9���v�J�M��.˹�OV��$Y��P3n\�:��)Ζ��r��6��}�����uL�e�Ɔ�g�:����)��D��z�+�g[����.�	�N�	\�Jo�0�;9�\8D��}��z��̮���ƞތ1ۛ��_Iڝ���3㒜]Cyg��xIYrN�9�c�J�(#��֊4�o:�3Dޜ^]@of���wbóx-=�5�*Y�β�v�")_��C2�;4�JRQ+��Db`��˹H:���r�u�4.U(��\<w�k�\�=m���:��:����{�wwwwwwwt�6�I;��y��Y��Iu��<]����5p�������[���)�fJNlbO�Ӽ�ӑ���]k��&���&��țy�u^��wJ�����f�b��l�]������'wwww7��ُ�����{�Ք�)�Zʻ�Y���T�*�QfI�2R5d�H�F��1�N�.�� T��'	���F���{�s��^뇴ߧ�����2��ɉ
A$A�Q���R��G0H�ԧQ%�%ʲ�K��,�Ax�vb�ᩊ�� �0Q,�pEP�@��}L�!P�f?/:J&�J1HK���
�e �L���Dx��6ܛrM-�a�H����V�%�M�%�'I��4E��uJU�&6�b��`���Y��ꛤ�#��Ȣ*:~~4��p&�\�]�)���^m�FN$���m��)6��eGT�R��7N�>^@�B�R�EJi��$Sf�․�RHȤT,'T>a�T��}We�[��*�*I���MB3�)AH*S�:.��!�u��#lq��d�]:��S�(�fJ��
QUb�J��b��gד������	=�����e�A�)4S�9(2��R�, MR")HDK(�(� ��i�J�N��&��,���mۋ-�.T�U7SAY>0���W�M��\�D����B�t�.��T�W��IL�>\��)!(DRf�u�J/��;]�r���g�T#(R4E2�z-�˨�T���롵G06�j��6O���xzI�_����z��W㿣~O��]��@����?���w�����?�O���sm@��ó�gN�T2�J�L��Qk���z*��+��);rj�Y`�4
�FBU�C�˧�۾�t�*�M[zZ�yB�Z;���}]FN�wѐ�vx�u<���~W�e�U�lPe��p��W[��]̔C{�ۦZ9�oU|�d�zэPp�*Vn�`��[�[y�oE����9�V��1
�U�Xx]7Q	�4(B�oKn�p�Yϫ-F����]pN��`S�5q��Ꜻw^�=��A\���\+�]ْ�*��,S���n�'6g4s'���V�*�Y�����=�+LW�M́��V���WE�y+�2�)�|��:me'��5I]��\hw�P���ghD��S\�̻ɕS���k,?B(>���B�J���pn�>���.��J�z9!�ꮻ����=����s��4
��l(=:�s�~(7mP�Q���#]4õ�/��;F��r���fq�7�J<�,��9l�+�#w<��l��p"����j$�W�S&��&Qu3r��(��M]6G�L�wX.U�ƱK�mV����*��x�i�z��mJ����]c��Z���8��w�sJ]����>�v�H��VfU�Y(;�^��-���Ew���\���kR�����o&��T�C�XͰ���LtLt8��������]x뮺믇]uק]u�]u�뮼u�]u�]}:뎺뮺뮾�g]u�]u�Ӯ�뮺��]u�_.�κ뮺믷]u���u�]}:�:뮺믧g]u�]u�]vu�]u�]u�g]u�]u�]vu�]u�]u��:뮺���]u��]q�]u�]};:뮺뮺�u�u�]u�ˮ���_n����u�^:뮺���]u��Y�]u�]u�Y�]u�]u��:뮺뮾�u�]u�^�u�]|:�:�O>��u㮺뮺믷Y�]u�]u�]�u�]u�]}�κ뮺믧]q�]w����i���6�=�撆���=7�LU_��l=�}iZ�Y�i��U"��I��@5y%�O�AZ�b�+�Ʀ,����{Y
��'�:����ز�wYY�a���/�RI[?oiĪ�������*j8�B���]G�i9/Dk�x%n�B�m��݄xY���C�j��ۢ�";�eW���Hw8��*{��}d�F���%wg�D#�!D����2�\� ;��6ni�����Θ�vtI��ߢUy���|���� �=�s.U`=��c"۶v���õg���9Α�Js�[���tR�-Eur��!�+���˥+7S�5��k�I�[*�œ.]���	R��α�NL��I/��i7UZ[$�.��7[��$�$S��'�\1=��qU��R�
�P����]���Ĺ?�{F.�S�rtb���"���+�q�*
k�;'&imk��)*!����r�T:`=g�%.#��
:s�u[�v�tF�a�C�wV
BL�Z��r���u+�+c���of.�EJ��$4�.�6PR��jL.�7,ۥY� �QK��o˱���i�� .\D�,.��s�M�bŠ��S��S)��r��nʕU�
!<�v�:�+|�GmglF��\'�
�`����>�,\os6�u eŎ�d8����wR��y�i�t��,U�;ȸqQq��c#c������c�ts��뮺뮺㮺뮺�u�u�]u�]}�뮼u�]u�ˮ�㮺뮺�vu�]u�]}:뎺뮺���]x뮺뮺���u�]u�_.���]u�]|:뮽:뮺믗]u㮺뮾u�^�u׎��u�]}>u�u�]u�_nκ뮺���]x뮺믇]uק]u׎�뮺�u�u�]u�]}�:뮺뮺�u�u�]u�뮺�뮸뮺뮾�u�^:���]x�vu�]u�]}:뎺뮽====:뮳��뮺���]uק]u�_�뮽:뮺�u�\u�]u�_N�돷�����f���6�a�@0w��os�9R5��W���f�(	J�.����tF�S�)�og����*0�ѷw�q@���T���9Rܠ��%(�k��T�4�t병����q5�IQF����*���ge�=� *��
��{i�J��o� .���n�"/���ݪ�BU�jө��|m��t�ws�j�M���9��S.K�w%<(*�ޫ ��ˊ@�'@P۫j]
&̮�&�Zރ!� E�C37v�.�/����X5�Ǌ�eU�HT��\c�}N#������(H;P�b�n&�wP}�qmvm�=��-��8o9� ]V�xG�I��x��[t�5-�k�JGԑ�X�5H��2��a�61J.Z�Tlώ���gV��
a��B�U/��E:�u�j�
�b�0B�s�i���ho��D���n�C_TR�n�]��YhX�58�cv^�]�#gS�R�p	!�B�l��]���,�E�v^P�-)��VNf_X2��\����lV{�S7��dZ2�k)n-�VE�G����!�1���f<7)���ܧ�&x�b�P"��Y�����9�;F1}F��l�}t�qQk&���� �M�X��U��_v봤�.d:�����у6 @[��E�|� ��5`��Z�2��Z���$ڞ����"زvJ������,GS�3߂�JU�f���{����cf�WX~��WtN(�xy�1��� ����\����E���Kӫp�9G&��x�x��W'���Q+˨�Z����/�I��Õ�W	�yk����WL涭�(s�>H��勚\{�[���~9~�!���Q�;&h����F�|�&�F�;�-�`N��+/o�F�:� ����NZ9��9�(��zuLE�޼��L�ҏ
.q=�1���n��5:��`����h/CS�Яԅ�e�κs��dY�W^�R��̾��z<�Y��}�ĕ�+�8~�nX����!c)��9}��g����I��n�\�㵹P6�]�kdY����!�Oi(ܖ�֛��;6u	>F��HK������ٴg�0݃x�|5�9u�٭u\�A�$�Ⴒv������6X�]\�=f�B+��f)��gk^2�7�4�ũ�r�ޅ��OM�Kh�<�b���jVU���FR�d(�T�Y&�Wq+�	�z��-ڹO:'	bf,��uOG4NW.;ZEA㾊;�%��Μ�#�XC�+;n�9�I#x�-M��]FJ���r�n�U�:�z�(K��������4�>�{�yI�).�-j��j7\
�z�iXh�`q$v���n�� �oA��{H=�JOh�p��#c[.�^;���CD;"��[ѹiqj�a�(+` ^��t�kxm'B+�6�b�$������Xs
r,���5��ę�w!�4��4��}�L��:�
�,-�o��s˵�+�NL!Û�%^�6��c� _S�4�r,Һ]����vf��&���W��ɐ謆���t{Q>�������p�vwa;vZ�A&�ɺ��w8˷�V�1�W0�0a�V��0EMI���ď��(T�1WVfU�1J7�nvk�
秓�rp�j��1F��ة+�j��;1X c��&{H�7V�$72���`��E5g�����K"sa�A֠���O�M���W@���j����[�a�XaV<�"��60�E��{�5��
�U��|��qX�H��MGk�������s��%֕N��#x8nR�E�:�P��}��h����-ō�)��ܨKv}wy��,�ʽ,��t__ p���ӖfA�x� ���x������|�
���>�,Q�;����]x����0��9�9��[����t��+�	Y�!�In�m�԰�U�a�Ti�
F��6�QZ�ۡ�'L���.�>#m����M��ix�(h����ڹ��v�_vQE��Aу���������y��Tb�1�2�첵w](�%�^a���A���oR��fZ��(Q��qkQ&�4R�]Mf���}���8��9�M����R�}�1��z�4�����f�yQ.E��t,P���o[s+�ka.����D`�C�WTs��pNм��^^�G�L���K�!�z8xmۭ�p'L�D�7��.�o*���b��b�����Xv攟>�JwU����yO^�{c1�E�T�*ѕ��*�Vc2��yl؎���sB���I�*}#�Y�;�ܻ>ԥب��+�M�V���8�u��h�ٗ��k�y�:�Vx4�m��w.��,�h�iΘ��|�n;W;�8@��2q��*6�U˨�y��'����8Zr�%e��a�nB�X��y<N�2�ʁ��+���6��m�\�3�܇/��ҹ��%R�m���A ��F�"�KV�W0.�S�*��#��ڙJ��[��������j^�Uu��n�0;�08�yx*�sa����G���)���3��s��v@u]9��.ү��O��g���`�@�:�q���
T�f�jv�۷B�\8>�2!��{Y�́�m��*v.AT7E����9պÅ��r�;6\]�j�}��D����2��Ee_t��z�%�7��Ya���s��fBp�=նL欣�G1
D㽖9m}��w3���s���1u;.��gX�n�c/��qnVG7�oY�Z���Ÿ;�YW�(`˕��¶��ز�]�[y��1$��]��qX�"�,����޽�e�m�4)1�.����T;7l�[�LM��L�D���:^�$����cP�]����K]mЭ6��(�6f�w�{$�R�Z���v�d�v����\}��fŋ�p�0d��t��V�+9G�X��H`UNX��;H2���D,�d����kcIM9-MG/C��n��tCj�g06�Y�!P1�����t��%*T�r*����4�^���ǉ��V�:�O����p���<6$g��f�{A��+�"�L��vl��^�n뜪�[�U�{AS[�hLҁ9�[�r��![^����2�`�|�����E#&�޴;1i�y�2�7�]���
��c���u$���=	
.�˷�fU��e�V��vv(	6����f�͚���lTȋ2��Qj���v�s�=��d�Y;��1�u睛O�|����x�,��o_#n�]��Q!ݯ��٦�v(#���Y�};+)���<e��ݹ���3NtWF���绢�����#N��1w7i��9�tb��z�˼5��mN|{�����y�V�a��!�Xr
 +Y�u��"�(�G{��ټt�,/<�9Vk��͟L`tq4��۝y4h��9Np;����j�nZo9iw�a�WR���JIm�|�*��ˊ��=[]�	��N��qP��Nf=1�cj�&�sqw1�o7�4���rn��hn�76�:F�ě�l��ƜsYh�����a����l؃RX���:^R���K�j���Ҡ�f8vS4y�[,vR���VwH���^�d�H�'��Zn�VT�Ց���)����2��KC{h��LA�"��V�r��j4V��e,Һ�i-��U�w|GGiI��W�Z�GMl1!Eͮ
xKQ��[I0�=�v�f 藽����Z:./.�f�1����֬��X�t�]wJ�͊.WWC�5{ݍ��5V:��hz��!X����-�*v/���w@����,t��#�1Z@K=:�ԓE���n��^g`�Фqٜ��ڹ:(?p��J��ʝH�}�k�:=��᥮����`�Ky����鵕x�Ir��%���M���̾Ű�e01;�f|�j��ȫ���m�w�fѷ��\�c���@�r�W��q]�W��=���k��u|�i�)(� v��S��۵��+y4u:�*��N��ۻ����"�Lmܼ�G���;fU��u��EɻA:b����ì;u�*������WjQ��m<79��q�N�{s:�FvM��m>�։ݨ��Wi�3U��}&X��V��|/t��7J�Ŕ#�'U+�Wc���Cv��ef.c�D�n�ʳ�9�zk�3Xӕ*������Iu�W
��6����顋�\*�ޱ`��ƔGT��3-���ȃέ"���ձAV^X�^�ZS]��bξ3�Z4hn��bB\�{C�Ωz����o�K���h2[L�`����z�78%��r���w-5V�z���6+��vޣ�̃1e�c.��r����)fѫ�=��y}��eJ��Y(�+:mщ)�t>�n7��5Bͽ�"�:#k-iZ�c���O��*�I���<�]��+q���!t��ivk�gG���`.����LRl�(G�s�ֽn����;W+WrR�jȌP�%ʪ�&��M�G��ی�,b׺F��v�c8Ue�̅-�٘���mN���v��oJ����i7�aU�B+�,͒��F`���4c}$�{fU.˪,������Ӵ��K�a��/���ݰz��çB��{���UΧ�������m��^8�cD�]�u�.�+BwF ��R՜�F��	wcg8cv��ɂ>z�[Mr<��dY���u�B�_$:a��/�$`�ȃ;_V�ҕw	�5,��yWv'�㋷,A&������+�Y�)��	�֮��X��N�e����s�)W<[&f�F=�4i�)�uwc�6�&��:��پ��� ��ebʔ��e¦�9x��tjm};^��ku,�_c46H{�D᡻���[jܕw�Qt��ʰ�H���*ب�I'{�z�U����uͱ��<�
|�k]F�{�lS+�x��Kd�t&h�!�]e[���L�53��t�4v����M��{��uϫ�;,0�ཱ���m�:S�o%�����sK��{qunE"0�@*�fq�JЬ}X1	4�G/0˧	�k��{T�@I$���������$u8��Kh?����nZ��R�
�yr;���w{��ن��#�g0�Y�^�fe�yA[�/�����n����oTX�ܺXW�V�{�1���k�u�F"�[�O/v�w��D�k:ڳ0͒��g[��S���.��lý�
��8r�jU:�֍���������  DG�$����\��#����G��ԛA���������v�4���4h��j�!��t�M��f���
K��2�	I���:5������T��*��^V�C*M��ַqn=��X�؟Y�״�g#Jܡ���ܫ
�y���ԙV��E��Î���b��^I�$��'����x8��U��oJݑ�&k���L���vֳwq���p�>���/�"2.M��*��V��,�R^��J�w���mF����s��S��}�7��!����v���ɷ֨�`&U����u���ʡ�iG7�4ŋ����s�l��uM�FM�RW+9�.���9qy�{�$��27{��j�X�;v�*z0|��:E|��s�%��l[u׵�gCF
��Ly|�(Ά�f���ì��ζ�bՙ���3�moN�Xz�'wmlל�M���O����!%�S�|eǗj��3�s �봪���:�m�ab�+q_u�G"`����[�9V���7�1N�ZyNgBۻ=�Ս��J4ss���b;�K[B�Y[�CR'F�Fm�Л�>�/�ඝ���������W�_����)����`������3*o*�1�bj呮�F�S����'�W�F1y�ܧ>�������-�p�c�/��-k%w'O�̧y˦f���9��H�_v��c;{����6��4�z��ǻ���y�Fi{���y��M"�ԠA'H�aD��~�E����.ϓ�:�RP=�<L����I�1)* �i��]SOČW Ӧ�� �F�U�ZS�b�FH>eV�FK#��2FA�YC��U���-����W�䎈�Y�J+�v^<z|>�n��u�u�]u�]}�:룣�bbbbc�#�A�@�e4��mT��g�O��A>��"+�T���+�QɔJhMy�/-[z�׎8���}>�u��뮺뮺�vu�]u������|پ+Q]+0�ȲH����'�}|�9U�MR�ihY�$��Uȃ�{���r�e?hr��(���W"�TE��eʺ��s_^z�\슊-I�s�uB���UD^e:5΁r���8���U"�" ��*"?%���{#�Z%�wA"
���NTUL� �D8N�
t�UQTr�d�h��"��G(��9DQTARt��(���H�(�b�0�*8U�\9P�,�@��`Q�,)Z
�Y����Dr�E	+�%�)3R�E�Ģ����M*		
(�]+i`OĲ
%��"��>Ǻ��(��p�?)|�<Q�̢��ܧ�U�,���.a:�;l�PuM٭G���.���p*KL�[�w���[��W��޻�u� �k������uIM��o�L�N�HXǽHwkpL��d��.L����6[Aj*�����e��%S�̕�����F#+�%�f��	E�fW�ۏ�P!��Y5���F��U�<�y�G��U;uq�#h�v=����H޸���Mq4H�U;�[��C��l�}[��ӼC��=��x5�nw�z��Uq��f��=��޿�Ϟ>��zP|�nq���y��L�8=�P�o���-�uz�_]T<~�0�n��OslŎl��jn�ngv�CT�����<�~������y}��������i�{��7t�Kӗk)c���������/�mY�ʎ��S��s�������G�����=�m��d�s�vs���W��t�˝���H��^�m�D�%�
:��%�߇��9\�Y�{Թ���]ޞ���*>�=�����3|!]�jA�[��h���}8�Z��|��m��P�����z	3���i�y˧��5@՚���zȋ�=y���]�:���4� �Y�7����\��K�b���`�p����6��`W�Ǵ���x8i	����Ӛٓ��P:��]�� ���,�wV0�dd�~�6��ESy-�أ*k%u�����W�LT�\��viZ�Զ2sT�2��'�vD�K;[�`�-��;gX|_,N6{|||vs�ۙ�5�<+'���[K�`m�ܖ˪{���CkVK�;~���q��(U��=tg|�
v����\���R����Y�s�޺��q{<�����M$��w��>����{�"�I����Ƀ �_ۯ��=�Y�N?	��¢tu��ř�禧R���\8ٙB���v�ڟwb�{ݘ�Q�������5~�� ��/���W�*�� �������G�hOk���˹�7�W@t�b��:���|��������q��W�)YMvw>���X*����{Y�׼.��n�����Njh��|dc337��vt�m!�*�������������[�484o�x=�v{v�ތu��i��׾���# ��A��I�>��q>�x����zi���>��q�]>�tq�]��x��w@�]ʁ�=�o�'홾O+�7�M��)z��=k���K�;��n����_��j���d�Ͷ�?�.F��FzA�i���b�{:T묞Ͻ�V��6q/��A�4$"���e����]���ֹPu+��u>6jY:/�]�L�u���bN��Ӏ%�R7J��u	d(��,)S�^>>*�wggv�;�h�v�Nn;Fqѽ�:��j�l���/M{�[���1�\_�f_���z_��z����$
�xI�U�<�y��흂ץ�ܬ4�F�~�9���!�y������ޣ&��쭏��o��7��{�)��s�z%��|�-� \���XPz�_�L7�����`Q�o���=C�-���w p`��I�}�o+��@��&�<�<��^���s6��Y~��z�L���v�u�R:�����:1�g �N���a{�������z�:|��>]����u>�|��R��v�C��H��C����>�B��Ⱦ��ǽC�q���jݨΚ�Xg����lŷa�$,F�P���M��B>�|}����b@ܗAfR˼����<FT��^��}r|�T����.��?^o��5��AG��]�I��|m�Lq�O�T��^��2�i8�M�72�s�+s�};���s�N�̠�9Dzgg�У�D�l�{�Ys��z)L1��`����y+=f`��\�\/'Dk��X�Y�^ʄ�Ei��}�K�c3��[�n�[�[�L-���ΦwZϟ�=��j���;�e�kf��A������'0c�&�D���u6%�Y�$H��3�zv]dGzl�d��v�c�=���'i��	$�f����O?��	���B�`���� UD��YϞ�t�F4��ng}_u�������*M�6�݂r�I��筤Q�h�0�B�]	Uc�O����z��N���{��`
;Խ�s�]�� M~�Ȩ�m<o�����2��{��P(����zu'��i��Z�JY���0wV>�u�M!���i��&�μ>M��s�0)=�;������Vԓ%�����ϰ���=�Kv���f�7{:d=u�=~��0�a�9������������d�K�.�Ot��l�`9e�5���jȈ�g��(�=�n��"LFǞ�c�	��H�=p;�����3;;���4�D���۲G���9�� 99���H8�u*�g[�lu��cuu����#�gq���m"�W��%��2���w{%�u���o*Z����j���J�»�:��e��z�`����z$��>}�a�i�egp��L�WJ)��3J!�1�`���0_;���7i�MhRӂ�ČFr=	ig;�I2�����J��+z{���}E�y�ک^�-9qwIϱo�sh��j�����Y똈T����AE���?]<���{��*������N�Ck�V��>����w����f/{"2*��N���m�p$t8�g"����#~k���G(tf���t'0X�Z;x���T���V�W4�i��m.c�ٸ���O�h�������cq���/�}��8;�w���0˼A��m^�K�i���:�o���N�7��|l6��s;z;k��q��;�dk�9C�{o���Oz�-W�2��=��zvC�96�|`14u�sެp9������#Y��4El�kI��l����j�KHΚ���<�(���,��U�����-)<WV�� 3Vq��^='vɭ�
7��븞�f�Z�I����ܡ�ӎj���$����&*�S��2�f	Y3� ���� 9Y�����9uw�qi��h��?b�@����e����k��^oR:q8���OX�@�Y1�7[��v����qZ9֌��Ghν�f��鲯ڨ÷g�����ƙ�E@�恇tookt��wg�͡�ݳ�}�ԟ{$����^ս��Y�ݨ:C���V���:AÄ?fO���mxa���z�5�Lvs���]�}G�iu�y߲�\ʋ��}�S�q�ڣ�.RNY�!�f.М���;�.��<��쫷��S2���&|���a�<���'G�O���R��7`���*��c=��m�-����d�n�g�._VN��jc���'�}B����ˬГ�F[d[~<�ӂ����������}=$ߟU���/����ij1-\&�:4<V��9rkf��:3�V�.�+#(%ܹi��}|���ڌ�_�	����~jw����S��\l XqW<x�:8�1��{S]���M���Bx���"�b�9lVc��+��z�(��oc�������Nr��7�+'�{`�H�؆���F�孝��C�M��&<�Y�Ҡy�ˋ�&)0�v�GU���IKN��L�)6������B�T#�����[�������l���T�����j��;��fj��?�%�y���}��b�q� c����^�ig<��D���wt�	6c6��K�P�sf��`�������-q��&�.�]�0��l���'(����n������&��L�)�i�h��3���c�-�}�cn�w`��{�Y�^Psp�F�8ʫ揷�k��:�}��������mV��G��:s�g�^���r?7��-�h.�7���Ѩ������_T����k�Kiޏh~$�i��-���'���=�7��IPn�$�3v�`}����U�����t��ng��ݗ�������ڈ���]�
QaA��[�0ﺠN�D����1�^?�o�W�'��:,��uZ�x���$_���k�dF���ȫ�܋���)��~�h�{㵆���aS��݃�.�Dk�;|����7r�����\㚕CK�v���	�rٜ/[�Lo��7�U��^�Y3#����n��[M#�\j�n��Go�F7�^�b��u,�jd��|��\R��w*Pܓ��ar]�͑��Ux3d��t۹�X�{q�!�\t0Q}��N}�<�^՚�` :19�wot\s��꿾'�lof��|��s��p���M�o������~�{��"8��1ޙ� hwO�G┰W�P����^�����S�x�bۄ��	ϻ�{��3��g�eT��<¿�����t@��ܚ'+[�pQ�4�%����q�_�=���w�6��h���ˏAգ�߁H>��_L�)�5��oy��z��/i2��@��^3���wN5�Q���&{z+�̌�|z��m�u�5�R�="5�	X�'Jzg`W��q]~�g� Qؿf6τ��'���>a�>�5E�v�=ݦ{V���77�Z���O�U���w���:f{�c�D�}�=�\׸	ͷꮗ���^u� ������U�����<�v��f�r<#5¹���G^�h�u-v�=�lq���яL�5Ԭ�0���Ϧ�{�`,[�\��tv_ �=I��R�N��1ffvv6�ӡ���c4��8�2�	Io&O�T}w���#+�Z�QoQ	H����*�+iKR�i4��Q���nbQrSIJc��o0y|/���7���5:l4��k�;٣�g����<�?��OxTQs��]������6u����un��9ݧ��nl��jR#h�=�(� 	��{Sޔ��r˾R�ޭ3~�1��s �ۡ�y����-GA�c%g����������"��~��?g��ʗ����W!����mdL�^��g��]�����E����H05���Ա]t�����h�*fp��|h�S��&��`�Hs:,�q��&���7�m������ϕmOǰ�o|)fOm��z���L����97����𡫍
�x�����B�:�}�6�����ʺ�{j��%�AV͐�G�5&�}��gR�"���%���g�0 x�0�4{M>;_]�D?fw�*{���;�C2�2��2{�[̚�y��gӆ�~@���zcB�*���ʔ�*���ޝl]0ySͥ�b�`,�Z��ۓ�/x�JW���)�^�ܖ6�=|�^����:�}ݩ�f�wg�ލ\��X��yvJg9�z*���;�7�+\e��T�yηN�9�YQn��\�	� ���k�o>�9��%�<�P�K���S�`(���:y蓪�ޯ/]�[�5+�ةZ~�պ�&��@�Eß8>�zO���U�+�ږ\���6��zdT�Οg4XdY3���=b�����>�g'L�1����݌6�{8��q��=�`����on�M�h��X#E����g����zߘfw�-5�Gf��\n�'6�J������c�2�����8�p��1"ݞ����<�����%�^V�rJJ��wN�l���MQ�P�Ѥ���	���K_4�r6^��/�pg�����N?���w���._t��f�vwd������N�V�]�+�`��t����:<��n�j�"�Ow��|�2�?uf�ϓ�8h8,w�eR�����P�6�/Ot^��{���<��[{����x����Qc��� ��f|~:�J*��T�s�𧀙O4���],����Z�=&�"nm[����tj�{�к�x��sY�Y���;}]w���+#��R͹ĸ�齘c,�+��`�7z̷�;=]�d����5�ppY]W�,-Q�9U�1�F�ق�먢G�]�Vef5����:�8�Hk� &n�R�X���:�[��Q�疠���F�oIl�LXU��v/1Y����n�Wm���`-��L��x��4�/%�M�p.�����7K��׈\��۳+Wl�k\�Us�ӻ�u���[�����#��38;{7��Q�'��e��t���z8w�1�4��|b퍽z�-H�+ka�i1�L�&�/f���K��XVC٭��j�<Td�%P�����	uaۇ�+�w��rxn���y���R�/p��L��u�4������s�*�X�T�Wf�)m�H��`�R��OZ�ƥU^���m�v�l�CX����j�&N����g6�8JD���+۫Ѫ���+�뛼�!ޜÝY3�d���QIƞT4���뫻ڪ��M�K0�bP*zޓ�7#�M-b�oWNW��8���Z��V]!����k�VZ���jG �<,-��ƮsejM7��6���m�FC��ou(�섒�έ0�\�AU���Umi,1�����ǲ���v���un��j8��Z���VE��u�@�8r'�_#}�A,���|5�Ʌ���YxY�x��l���lίSͪt���	�B���]���X~��O����c���Y���D��}�*`��i�E�偻��y�r���u�U��Q��+�2a0�4V���v�^ʇ��]Y��#��&%__���Z��V���>ڱz�>;�WQ��
�O]�W�gpQpp\ĵ1%��W��ʅbg3�����ucT���R�ۈu�S	�6\:V�cz��`~t�ZԈ��9�e5��,�d�8�ڎD� L]PE;��)�����lV��U�NL��[6PyQ�vA��\��4y����设6Ű�,�X��2�c%.%��㘭�����֐sSΰN>2�.��b��²��x`|8kgtUgn��+^a�_Bj;5���=|g,��}P>����|T�e��⇠ci���3�;*��ڏR�کX��.s�n����eI��CL]�B`;
]t 5�����74��1f��3zfdd�#0^= �ݫP2�#�N���/�m�����ZX�u�F��5�|r�S��q�u,ޗz���\G2�X쥇��[��np�Q_�[���]p�Rf�]ۼƙ��pl��9Vm'#���d�F>��*>���{�Z�tZ���q�u6�Z�y��p:�̧�r�z�ovs��w���6_>u>�H�W���0�& �qL�Y,�N�\s�x)9���{�p�pp���3�b�����uہW'�!���� �J�N��(e��n:ػ��z|>^�u׷���ۏoooon��vu�]x���^پ~����j��-��׹{r@�O���S���C�Jq�Q����pt�����t�Z+m2����w�(i�Y���G���O>�/������]q׷�����������<x�����s�9��3+��w.]G)�F;�v�{�1k��z1Pw~��X�ʯD�(\q�
rC���������1���v��p�goD9Þ-l�:�+��ۄ����o\]sl��9;��m�*��''P<�s�/B�	�K��9�8C׼x.�xi)������$�8�O������ˑBH�Hjz��E��s�:#����/f��rB����Dtԓe��s���{���������3D,�r�G$<�Q���RHr��s��o{��
�T�����\�����t*"��)�=����s��@Y�	�,���xC��z];
���9��^�����(�g_�pG>��Ң;*;#�UA�Ȉ��)m�T�\=~Y��z�dQ�4�8�[r|�p�!u��I�"�"|��פg۳��.����\Ӻ���P��\�~ށ����J�{��x����m�)T�:�k�A�D�B�A�ݎ�u�����\Z������lA.O@�%��o�瀢&qzF[�Q+'Ӄ��D,ٿ���_��G������=���	��ݯj��^eD�%)��o
*a:���T�A��2��=�P���ޛ���'Y�̏��G�c&;af$lg��c^�,���(u[k�Vq����T���;�A�P�$�;`w�M'*��o�=�Ά/�o���8�ON�����@������ @�'W�1F{�G~T�����s򖬸_~�A�Q��ʉc�ɤ�q�NUL[]�և���/��MB�>�����l\�a
�Nb�2�����f��� �s��'#�gc�gj���=��1����U�x6��	����yl�m��-� *@�u��xy��=�=�#b���[�{�)}s	�:���J�a9�w8���
Z��&'�Vh�X�[��˾c�+���ե�Ky�_��!�ޘ�^`�зĸ��K����q�� �6����в�5Up~��ehjΖ��};���$�߀���4�a���.?ܨJ��8Eǖ�;%�10��r� _�/��~%,�كK��\q:�����6��ߎ����g��?&�_>���[�m�<��ɓ�G���~�
Wp�[c
a΂ع�y�#;�K�����Tx8������-�yC/^���^�m:��|ٰ��rj�xD�������uu�����W�'�])���m	,�LL��4�����T���D��z S�����~�땣GwWO�Y�p.�fXOO18<��D�����Ba���=�@J�_�&���t��`�SE�u��OG�~������"��L)���l���O$}�Z��-��Hk��d���6��|�=�?[����.��^�S�P����=�t�9�aBM��i;�Z��C���7��[e*~�q}.�:�����C۷���_��u s��
�=ߋ����U8�_b�;W�-FRy}Zi}u�_����t�E�d 9R�� 8�����d��>��-���� kf2�3��U�,�������?���<�S󲼫�)a���:B��Ho��,9n-w����$�1j��6;����iw�%�^���L֚��c�q�g����+�f?T�7�u�����/fD����J�E�ݟf���W��o{�����x�����Y��s/?�����Z��,���F4�}������_eu���,�^&����o{@^��y
קYsoMa�?Y�my+�O�,j�am^�S�����ޙ�G4/���S�j�㣖�H���m�i�����vK�AziT��5
UX��T����:O畬긳b�P�A��T׬��]I+;"���xմ�l����qk��E�3*+��MR��Mk\������M�t)��J�ʖ��܉$xB��P���Ū���zu�>���A]�%?�Uk�S�s��J`,��L�����0�5(�qN8O�,�����֬���s03R=�.��ӷ�K�O���=l'X�vɡF!s��q��=C��҅F��o�s��;Cq�}���r�d%��3�;�����2A�4b����ؚ���Е9\Ֆ�k!�ڌoc TS~Ē`��(x2|[C���'���1���P�ܦ c�i�s5Y�Wm;�8C����� ML��v3	�H�^*V��Q�!�ʹ��W�:w��b!9�7��-2�ͼ���	�\��2Y,��'�b�j��x��s�e����T��Q7�{K�r��_�)�i�I��Q�F�����U�Ŝ��R]�nq�䤰Z�ƻ:�v�t)���g1��#ȚO���������+��[��ؒ�]ѱPN@�ʍ�A��k�C؊�s}����4l�A&�����|����o�A�4�]�j�Xah��h��~xec�(���x�ʀ3�H�"t�{ئ��gןu@oG*�`� $:��H^����~SQ��&.��>��$'�������G��g%͜x��}��Ӄ���!Ε�3c�\�n���;���Uư bg/����>���ۓ_q�$-�1�=�D�ȋ�?k�Aǜo�e�qb������=R�hm����g�k2�����B�y�37m�V���zX����q�����~�R�ɕ��p�fA��=)�8wL�T,>ɺ��!RR�Γ�y0��2a��섟��#�׸�'�M�i�4П�Z���, 3}�?WP�޵A��n����#>_�_0��������k�N��$2(@��Ĵ�v��Ւ0Q�����$C���P�[�O/<K�?54���/�����z�>�"D�2*&�±򶨫P0����=��r��}iwQj�+6}��~�����z�x�?M5�,�-�RB�25�#h��v�#�_ݏ$}մ����_�[TI|���@jkgc�I9���Ƶ��ZZ�r _M����`x#ͮ7���l��d^ǵC������r�ƽn��1vۂ�7��k�j�M��G^�݃�z�u�Lw=�酥�Mܔ�oRe����ݹ(�|mN+��^g[�uf1c�ѫ�'g��GG���&�����զ��1�b�[R�n�T�~k�כc�ugy�R�����8��qy��;��5Qt��7<ہ�Jy�>�ЂT�r���9���)�gH�<Ϣ�0L�KӘ�v��k���gywg���w��@ࣝϲ(��S�3T�ͻ����=i��薍Gmꑇ*`
�����r^�5ma�B�c��d��]Z�$�8᰺���ɵ��Mm�a�"���,+$ŕ9�.FA�ɵ=3�V���� {��v���e:x}`%����ņ8��)��4���X�RyD���
26�"{�Z�`(P�%�{y������ͮt<��������e`�҆�A�iϾJ*[�cɖt�y�F�6�C������,��_:�����/өO����|.`H�p�0�[����P��9��.IK�W7U�lM�&�#�Ǣ��_=��W����9�~���.0w�8����x3���)ih��]�`����@�(��)!b�=#��Ň8���O�<-��b8���m�MVC�{��/f]��xe��iKmOi�^�1M0[�G��d���2����Ljp>&�'͢�͗2��9<�{�c��G�������� �p��>t'+ �U�"8�˔d��G�>����>FB]�\�i���z<ÙB���(댰'�q��^�%f������8�茘� F`r�NL";\�qv���	F��E)��N0��9��{/^���9R)��\ǆ�FV64.S%��v6-�δ=����ː�<�0�0	��v,�m���P�N4̌���@YN�26�����<F"�'9�dҩ����R�zS���rcsU�黻[)�/�z~9�u�Kں�n�������L[�V��EAm��|�l9�i���K�g��3]�|f�y�D�/���,�7*uժ�A졅���/�֚�Uh��GDÆ!Æ"#n�Pu�A�� �3�y��绣��E�mE'��1�¢��cC!y����nؚg�c��{ݿ�Ǥ4��D�k�LT�&�w?�?L*Z�&&����V4�`6�o��{.s�.�$�o�����FQE	i�D�CeJ�>#&�y(�\|I���ַ�N��8ǾV���ޡ�j�ߚ�%�ZF���ܷ((�`gs�^��ҹC�G�I�bf��t�|���>��|�mϳ��"�m+,�b�O��>�VP�Τ�>0�vY ��SJ/A����y���+��^;�ͨu���ۈ�:J��\e;&����$�<��Z���#����H��V2�i�)����B���<[e�)!d|�~p$vO��:gK��oTe|����V�oH,���2#���ը^��Q���t�=7��@;��cJ|�F�����xc���5Z�L[9~�Yݾ���� ��s���"A�耐�f$O�0��]J>��#1*�ut���b�/��s�l���w���E���!��H�>LX���,�y����}r5��J}���>e�x�8��@�j���X��b�F��tN"�IwWlH�_��y�L���ՖY�'v�9W(8Z�WVh�e�e�:$ I�2n��.y+��;��U���e̮��\�ok��v��Ԙ���s��`яN�fG���:��;jʧ��ە,�ܙ����)�W��18 D��3��w���x��}|��_��yFB�߶@��Y���J[Ԙ��+~��O�L	�.ˏ��oF7K�ҋ��؋Vvu!�f�:	D���{ผ��@����D���7y��$LdAQ��˫ZhD��خ�݄x�ۊe�q��v�~c��y�@�"NP�N$�Ό2,t����g�z��Ҟ;��2`0lQT�0�Y�n��L#���ql'�`o^�!�=L�+�YcUkxG��b��p��g_DmưR�0�T�FZF�W�����Q+����ʌ¼e��&<���<�~��7"�;=?t���(�z��M�n@�����vޯ4Y��z���X�%N6x��@��T�[�NZ+��<mTl.��E������V/T�̂w��3~j�>+�YߞK�.�My�g.�0�N���;6�f�w�Hz���L�����b�k�y)�vr�l�9���*V%fO��`���y�=�F
?_f&�������ӜY ��B�<��L��GLo��{jQ{����Z���C�ל{w�b����b�`ز'�M�:����� *<Zzǒ�dφ�q �U�,Q� �d�ఌȦotJkfc�z��-�? e��3�^�Q�q
��1��:f奆���E�,�>�t3~�\��ʩ���Tt�$@@�O$^��t�l^v'#�d;w ӧLVM��s+C������;���
��]&�.�`�,�x�n����U�1tȮ��yn~J�3���O<J�$m��x�N�-ک� s7Þ��C�8��=�.=�VM�O�� �	��O@�2�RX4K8�̢�i�ۙ�!���C�-��|������P��w�beߕ	@I�<�����j&v2ofI���p^԰̊����r~�L���1�I*��
��"
�cd������$���K��E5
)�/a��S����1ٺ:�y.F9��1�ƠG�������Δ�H��7�vO,''u�h��Q�G���/�>��>T���51�*��&F�]�4��2ڽ`IM}X\%H����'7����1���ݡ��M�ӑe�`��h�)�GL{ޔ�BF	�6��Ĵ'�wǁ�J4�e��1�Ş��f`�y�H��q���1�N�l�'��g�a�j�P%8jC�m�;�t5�iL��U��g�+����kaw�/e�w���H���C�M\M����p?";�e���x���le(��?!�Ɂ��Ɓ{P��9RV@��ٕ�9�18�(�x8�.]�g�T�u(ܨ}ktN��u�	է��醧Y�l�ʱ��UЬŵ�H�f�)��+dᓿ,��="��l2b��}����p���O��O��ֲ�YU�ˬ�9k��O�RS� �,�U��4.�mI��|���gguر[<��;���\���;U(l�vf^��w�C�4;k�9E�29��Kf�N����:��[���{{�
#~ޣ�_���ĞO<����E[^���	�;�ɦ�_!�}��<s	L�[��qTȾ �ͷZ��
�/�㺨f4ԋ:ǧt�<e��{���u� CWd����]0�-WI��1�~�Slo�������H��c��5/���u�!�kA�gO���&pTh�!�T�q^~3���ͧ����n��ぬԁ���a��̭�(y��]��^h�O�@OCk�>��S�S��|���	�&)�y��z׷�f�wT��s4���oe>��x ����z/��� �l9���}�}BS�@%㽕2v��6<mF�z>�����3�-�r'�P�㍋�5Ab� .���r6��'zS��Q�.'��*�y�CCkj���d�"��=���h�;�U�P�l�؇�6|�L��ǅ5�ȃ�d6$��)��K.�ĕFd=��;,��Sͺ����G���u}1d	����b��ʕ�}�K��wf������x%D�/�zP������-��Q#�9V,?NzF�:ř��OH�i�Yw�A�03�b��u���x�����~�H�p��B�G��T�.4���͇2Ey��xf��,I,(��	�� �r�UۺKô{�qJ�/:�>�ۣ
��km;#xK��4����bm]��}If�ҵ@ɸ}�d*��n`��Q���#s���o��#U�o��w�n��u?S�J)���1�ʾݩ��O��`d�w��|������������q�<yDQ������{�ϱ����#�Z���'���,�d_O�/��&8���_}>�4�j,�x>�D�����3d��B�T�,�;�N�9�W�d럕!50��S��_��F�G܏:_��˜T�a�τ)�HQ��{
�����~��d�h�	̤D�y�nc�%*j�T�{� 55��$p������[Q;�������t�>��{�����1,�X+*����Q��i���s��Ŝ��{��<س��d�\`3q<��Άgu�uo=�d���s�[d���`ʭic�j��~��h����}_F�j<P��M6��I���U��*<��	]?W�p�]4��X�i�0[��oo1�,��z���ab���@Wk��*���Ņ�>[V��W� �d�|�N�;��*���UQ�ɪ�e�V��#��t�*�M�6�;�ؓ�g�W!�	��P+��_��5��9�[e�tQ#!��}��{��CӘd,L*ML&�;������$�[�v�|��ȲL{A8%?r�^=��'���b*_�'p�Ƒ�a2��*���\���~�FIu��z�)��$wv2�b� 1��t���Ѿ��e��(ar�DN��'4�o
�(.�C���h��f�nٓ����{Xۧ�V~��7���>�7�ZN��1�m$eԺ�� ,\�e�Rݘ�8z� wM����7x��j�7;6L:�Ϛc���H�ko3)�=m(��H���vDC���N��k���`��q;����kF�ڹ-�%v�ήz��G���K,<�!t	r�����G_][�u�j�6�Z��Ձ��ݭ�x�
�Nn���i�޺��mwm쫘��:����;���v����+FK[�w�5y�6C���w��Ч\.�ݢ	P���[CK��$]t�t�SF�3s�>)c��0�D,�xQ�٠��U]b5[�n�uwE��5n�o2��ے=�qڙ�H
�bS�5������h���ݔ ��F�&��cg]g1��\�Hk��Yx�nⱙ�*�^��fr�� tq%�v��ܴV��l�������(5e����1�2�RѶ��t�taN�e�	3��P����^�o��tx��o��;g��/m/\�T�[y�G�[�JD�]�މ�i0����Jh�坻zSCu}��n޾w]1�;}Ķmf�0��GhU�����(�yuO`��R�`���Y	 뿕ܑ�|z�u��rV���<��O��Jc��i�����Ys\"�$�E-:�%�Y�����h9u�5�m��%;N���vI����x�8��	��TEVd�Ƣ�t{�:�Z���oyt-{Ҏ]
et�4�R�MnR��O.8<�"ǃClaz�ql�U�9�`��xz�B �0f�R�7��'�G�� ���w��׸�>�wW�q�)T��nu*Bc�'k��6�Z�Mo^A*qJ��Ɲ쥨K	��qs���6�wSO�T��wW>�ݒ�䝽}	�)Ț��y�L��f(�^�1<�vvi�o�	k�/��v=�v�D�Lˡ��X*X��$ݪ��4�k�����W`�s�2Y�SNp�`���+z�Y�ӌ���i�=k�����>]e[2DQ��J�LI���:�hT�@i,�WA�Cz1��`�b��PJZx8�m�.��z����n�_+�2�ø�'5l�xiP��OL��\�uɬ��x��S#��>SX&��?��Kgy�Q���N�5�(��SڸR �g{B]m��Ƴoy�2̫�H�A��+��g7����j��dW�gk������>Xw��O�f��X,U%\u��a7��P���G����A�G�O�����u�#�͘%�W�:�8\�#�w\Y��Q���ZrZ�;̖�JpwB�g ���g9��7�����t��r���m,6��v�gs�ӳ�0��uQyc
�Jp�Ns��m�Bxګ�N��`ݡ�@rQ�/�郎��f���9	˟��X��� lI�u4tOW(�j��+It���R96E�(�ڌ�	U �'L���(��! M*�>���k��珟��+�=�׏7؟�{�a���/��N箵����2���rGP=�~w��5o�?���'�w$���Y9�@�W�+.�οߡ�c�Bq;ֲ|�3��������u���u�\u�]u׷�������������w���N�B4)i����
���ע�U�h��EDD�
�e�~�o���{{|:뮼u�]u�ˮ��ooo��n���~��H���0��~D/�/D� �f�@���Ӝ��L���]�.�s3.vQA	�ZPJ4�I�*Fbe�B��TP�g�����<�?#J�DaHg()�Ger.��p�#��8#�����}B+���dS=M��#�SH�r(��9GU��+��QpT�*��._��=yQ_��v�y\"��UQ�2�.Q�e��a'� ��aUUEs�]B��'6��ܜ���\�lI�%T�Tp��*���U���G�}@��s���C���._2#�����\#�U[��Ⱛ�U�9Pr�?�A�J-�EE��Zi��T�	���䖫i���I�k5������*&j���ܮ�����Ft��v������3���`��j��F �2�[原'H��x<��%����������ϗ�3ǒ�aT��~>���]��^����|��T��U� >,^�EV��evN�'�se����,z6���l}Kk#��f]d��؇���4�hgI�pR����xБ�ä��lx=C�3|j����s�Ŵn�7}7����j�Ș')�3��`0#��� ���S�CY�!��xP�o�6�a"0n켝�ͭN��ܰ(�U�xt�vϖ�!�ޠ����&��z�B���6{/�z�	ރmϨ֮�#�ަ�*�7\�W%��[:~f��1��Hry�۳�_o��lij��U��U�G�7�7�h��c������p�	:�x��B�>�pj;��<��l_w+uN�uj:�	z��Wle�G�5�����'����Β\5MÉa��;���[ޢ�A��hy�}�v�U7�+���c��Z����֨c�e�� W���X��̢��A|/od�oǪ��@ �/�&exm5q?� PvJ�(����k��m@�ׄ�SP܄Ǟ��'�w��SQE&&��}>���w�1���dLƈ�Y��vq����h�f��5��[�s/�W�S�!ӆ^%�����Յ��I�
���c#��'�7�^h�*��s����:�k�;1�u��v����h��W��ݫc��38N�E�Sz.�S[V�ފـ�޻�:cޅ��^��R����h�:�ܭ�Lf��_����g��W3ǔ"����������"o�׫Y�^��H*��HQ6����YGػq����+�Kv�c��At�fJ��9�%���2����H���3�1^���V\�j�5ʟ�V�B��ɜ_wZ��ia��t�4le!�i��A%�ӷ��7Z�@�
8�	�����0�V��r+M���"O!�a�<��0�1��3�6c��iO7� ��,,g�.znhX�t�T�C����Yv��B�,�X�T��%���]8�~��V����!oL|���K�6�\���F*�o�Y�҄^�F�i��܉�L'��|(�BT�<C�덠Y=�7�^ 
�����L�[@�!�ӷ��ʱ�I�ҁ}q��hkN�8���m�x�և�A�o�KM�\�����.�~�[�O��9]]��z��6��Z��F��;�%���B9�w�T/zd��u �;�x``�/6�j�e[Y�h~`�t�d�3�̼�٬㓀I���WE��nJR jeb���>'���|��O������?r腓�S��6��k�V��c~7#���x4�q�hO�����x��ď�9\ћYӹv���_7U�$屳
���uW �����*.��S��r�8�s�UHP��7�h�F;�yԋ���u[�x;z���1�ܕ�uͮ�����ƈK��ӌC��,�)����M��s���X۱����||_�O��zy*q�<y ��2r���aaw�d|�|��D:*<(M;��8�M�Eտ�/FE;�(��� �K���y���h{�;��+8���޺dm	l樦�䂾4e��z\sR�� ���2i�h�/�"��.��(�C�.)wѿe
�q�@��RK�ԁ0��ÇW��j���J4�{>Qx�3|�VX��<���g��b�K;uf��3�޼�v3�M��D��R�ژJ�����J�1�
����"��7��`����W�KI(_O
bB�z>�.{$"z ����ڹ�-�m����u��b��pjn�q�o[*�˫�<���� [sM��E�Ȥ�C�I�Ba�&6�w`I^7^F6��/U��z٢�n�_���'��>�p[p~2/�B��Q�]��x�:	G7HS�{0�_X�k\�5]��ԇ�_���^ϔ��N<�>Zg�Z�&@��ן����&�*�{����e�nr����:�Yd<���Pu!k����`�w�G@�˜,�, 	�-�~��g֤Kt]�Am�I����!�΋j.66Q��a��jƩ�6k�m�l������D�&ЭC�Ϸ�!d�Ƞ���r����ZRp��Ýw3-����>ף)W:!��y~z��t8���e�2m� \���d=ܗl�ǫF^u#'kFek=���E� �0���Ceeah��v��'3�sh�
2�~����D�1p�@C��	������5}��d��i����(vN���T9/̈́��>��0�G��:J�L��+��{��3�R����שt%�àײ�ZC�{��["ã�zw�Ws��Z��fy���H�7=V}�u����F� �C�	���7�q���%Cf<�}O�)��H��� ���>34\�D�h��5�y�/�=�����`�=6�ʆ�'e�!\�P���͍�9��73^hÆ^@5�hk�=}{�G�����(Υ�R��	3�U�e�x����r|�^s!ϟ�N�+��.�v-Wvw=��t�#��P�?@FY�4��i>a�];�7�$g�@x�,b��9?x±4�g/��zn�{�'R֦���h��nw1�O����V=�P���Q\�)/^���9R*t�MV�ϙ�ND-({9�6��7ͩ��p qٶ��A�P�ɶ�Kln�,�2-M��H����؞�Sxֺ�;�uCS�ב>w�qU�9�m�Ĭp;����(��`-�M�T�=��1	�f��O>N���{z��o�����A�@p zm��K�~�K_ *d�n5Z�*��X�c��p��f��.P��ٝh��ղ@y���~[/�a�/Y�؆��%�"؞�a�*?e��U��J�����;��;����Z��Di�pu�#p�b�Н��*�����N�MK���|i�Nl;tܸ(�T�E�r��2ٔ��u"Ye�q_�@�d�q (paÁ  G��<}~�g��< ��ɐ�n������^���������>Z��ĸ��QY~�3w�·�[r`��e�y��{d�/9�Oڌ�?�����d_u�䈯��G����k�~~lgdۨ�yym�Q���=.��-��oU��k�4C�.��EoZ�no;;kf��7w��s�n)�pk�6���oDzZe"S�"��H���z�,�/���x�����s��0���ܜ�Q���"qx�8�u/ޗ��z��/L�UO<��h�hOG6o���,�<O��k�Y��;���B��Qyt�^����)J�!$�����~��%^k~�W�)8� �M&�|�ࢶ[��a�}jg�϶������EZ����8�� ��Ϥd0���1Ƕo=a�߲`[��[�A1'_71zsOe�͈r�v��~���r ��&��Xx���f��_��s90�1v����z�2�B>�ܙ?EG���v�!��0��?Z�������*`鵟Hr'Ӧ�{���c�����뿄v,�J������QQ+�y�Ę��pxL��.��5��y��F���R�Ƨ�h-t�L��*UfWąԯ�y��|2��S��ˇQ������̥=���O(�]��E�:��.[�W�c�c�����jp�W-�ٴ�3�����srփ7�P���K.=VX�uQT۳3o�a��VՇ]����1  ��� 1 ����_h��@�3��TJ�B�	���b�����yB��dKeS���TC��鯆���3$��g�v���7�#ŉ�n�n=*�Q�Qk�y�X�&�²r�R�ϝ��:�A��vF���mN��Jʿ?��)50���q�5ݙ�45�L瓏g�����[잉���A?>S�9e7n/=��dH�Q�f/iِ��!#��\DW�b�6�q?p�}ؐ���4��/�!b�%�(��#�ok1�Q2�0i����|w�2 ��Z �C&[�]MI�����Mz����Ӽ��$����9�u�b8���[�������&r29�B��������.�5>��^q�\�O�	����e�az�-d�y��L$��`8��ڶ7����[/xB�hnyc�-���^�T�.�=T�G:�"�N!1�X��y���m)�z98�N*�2Y&1��m�u�kRmw�Y�{����$:�"b����@��	m������=hЭQ��ل�I��������W·��-�/ $�i֡�ͽ)���+��P�{�R��c�,��$��$oO�}8�a��e��#vw e��R�ێ����1��+Z�	�=?��3��l��O�|ZT1�[�aJ؇��<��j��>�F'~K_�{��E�pЮ���t�U�N(ΖT��m�F���>�ښh�PwD���?�ʋ���*��������R��+�W�O�c"��S�hkH�m���w��i=�
��@�x�a|v�tۿl3u�XKQ��=LZYB�9���û�_���Z����`U�w N��R<�������=ڭ��z�����/Z�J:���d_ӄ�F�11�B=�0;۞N��r��gx0%~س��ے���gs��oT���E�z_���E�:�aP�J���c�%�����M�W�|�=�|Λ��}���$|"��`��{�թI��6� �������c�S���K�ˌ��оNI���	��F߸��Wo��A@��i1�r��5�;��L�|ak�(����|�����Ʈ�M�z�z��?�g�!jBn�	��z��O�\��W=�z1��5ы�C?EX��8=ퟳlj���*��C���J:i���.ar}���m{ז.�{i�"�>�)v�*kh"�:,�\`�TG����ʻd����L�t�.u�-�����Q�8�)ꪜ����yFa,�h+���߃C��x$矟�K��M݃ޫ=q`�p����姙��Q�ʟ*<�h�Q�j�7b�%�v�]v�ކOC̝F+��\���6*��˨E���c' ܜ��_�'h�bc˲�@�X(���Hzs���9e�9��!J�]�/C���δ� ��N�S�*Ø��ݾ��m���^���a�ݱ�i�����o�U�u�%.<g�(�y����ut���� .��������2��g"�v��E�O��m�F_���)>��en;��T�om�4�跖�1��|�}>�/jq����@3�̤�s�J�����Y6(VՓn}�ut�Q�o{Z�]�xzb����?LK?���}�gO|�CyP�
���D���ߎ�u2��t���Ojy��iN�h=�<z�[/q��zYaEc���z 3�R2�0����84:�^��4���ջ׊�����;JH�'�EOz�Z?/�lua_��F}�����` Qց'��{�T���3wdxˇ-�z�ꥮ�(��X�10+�a`,��]�?Y|/X�Q]Nީ-u/��;��ߦ�{}����GV�!q+�=�(H���1���ڲ0�����w՟}�v�f��.GV�zu띵�3�B�˴vD3���=��	b���N}#2��\��[ڵ4�����qd<��Y����:*_ʡ��GI(�AWə��=A�x~��'�__��f�j��ԇ��f@*��47W�f��=�nsУ�`5�0����)��;�x/�W<�r!]�w7�t.�M���:WTj�j�/����~�>�{,�/{�s���lS��1��J����!�=k-wg��d��J
Ė��T[aq�%/㙜;���Nۗ�T˲�8��g�|�}-�*�6q�ܼx�R��^;��T�/���}��f�2��m6�e�N�=��x�{z��� �;��7��p�  ٭�ޱ~��W��A�9�m��Ft~�������'��?�~����@�{��|e+�`YV�<^R쬋pAn�~�O�����	`)	�ܤ0i���*ޱ�b��0ɀ�+*�l��U�r�5��Y\5��f�������-��a�hF?P���ƪ��v�{������P�c��x�k��<�ot���@��`�dC%�}1MmPT����?<0&y� �C��of�~��Uܹ�����ͯ��dVMu[j�NJ��������tzb�6|��� L���_O�3֔쉨�]{���M2u �}3i��)�0����\��lKP5��F5���.p/��1gp��Pm���xI޷~���N�6K�&��~~�eѲUG��{D<���لN�K�)E��ݻ8�݌��5H�Y��M��t�����e�d֑��1���;�6�}�N�.;�� �������܂!+#�0|��K��L���[K��ߦU�;F�zQ��G��.���^ݻ�2+�����}���Gug�xK�}�-B\ky���);遛�S���-�!�Zsb��F����p=5E3�ʙh�tr��,���-�x�|�P�L�HS�/�3j�&|S��_��UwLʲko�TB+b��C��Z��u}ݚ����އ���:����V�u������S�JJ�z�r�C��S�� x��g�ȫ���檭��0��:�^���^��i��]��=����	�� ���!��]B�z���	g[)�Z_#H��J&�W��(�zF9���?~��-$��4��טG���rezw��RqqU�}:ݵۼ���vY��%#�ղ2���,CH�r����WT:k|b�w��L���F9o�^�%�G��Zo�����lлu�<@�b��;�9����b���y�F>Ռ�}i�ec�s��g�����/V�-�G���nx��1EB�#�O��8y��(�lWMT�u���3��k+�e����E(�	YV�D��"�A>RhZ��
�,F�����X�i�_)���L�RD]A�~�դQ��d���.YA�Ĳ �C�(��}D,�9��|
h^}������)jj��Zծ��y��j��
��ۢ0��d��6�1b�0)��4�Y�����9p��ͳ°������L��e�)�&��b���d�cƠ��ȈZ�������/�t<K�j�C����A�'ֈ�=~��
6ޞ �ye�`���_�ߧMn�9V@/F���+W���2yP�\=�1�,�>#�޼��w}���
:o^�=Ů��f��r�����B���xr�
��N]E��j�Tͨ���.��"��s(4
�:rz;�4ˬ�l83*^�M��1�㵋�%	3�2����|��!���Ћ�L�'r�p��Y��E�k���0�*=F믵�p=�z0p�����l�tք%e�^^��e`�cN�lQ�; Ɉc�5f���L�z[��6����tH��K�܊�aڹ�Z�0J�s�;��Gs�.q�H��rmЅp��9��8�Ju�#��<f�ٵ*�8ֆ9��S���#3�$g���h�u�����!pQ�ֳ9���,�Y���w���F�c�6/�qt�Z�������f�=�+3c��/qݦ�wJ�Si=�0��
}T;�b>~��-��B:�`��U�7v�f3|7.�u�(����]h�6;J�d~̤4b��
�3gf❮u��fT*�6E�P6&=�V��`UZ�od����dQ���Mkky��h+��R����F�Y��;�ĭ3kj�� Sb*�V�=��.��٪��ƨ��HU�m�dw�ֺz�v��B{EeF�v];�~�M��ym콷���^��܁*��p>�e���S��\Kס`�qn�uU'˫%�d#7/5��Sz�/4oZ"��z��PaNmS��}J�'�5JS&�U�[��a��U{
-��]�Ҧ�w��(�=:���V�8]���GgEZ�0K� ��r�T`�ct���#5���b���V����=��,탋����wL]�{�o��\8tD���'o��N��(I��R�wr_:!EyC�ˀ��G�]��MT$�@%�,���/�iνw۬�萓���̞���.��L�N�ٮ{��Zq�2J�o�
�%d����|{�T"�D�(V�֤ŪË�ՋgV�.7�vE�9�7�,��R������v%��nG���	�+*��}�9_,gw7�iЖ�wl��S��TV����3{##/FoTN�o]z���I՟���i^k��w�s�ѩs����x5�ﮦ����/�v������l�eѓcFtWV���B���}]՜�Qm�)�Wu� Ou��)7l<Y�gs�Ć�ټ��$o`���S��lmu���:A��J�r�Q�g��I�;]W譬4x�y��n�Wo){Z���\��ogź�Rtݜͮ	[��*��J5ג�]\X/l�\9t��#��D)�����Z��:N�s&Ю��TMK�d�U@�}�(,�����|�Mp#Q�+�	h���T�r�=E�D+�
���Q��Q>��s��e�N�Mo�����6Aݓ;efU�� b�ԿdQ���L�*)�p����&K���L�gIy��}��O��������뮺��]u�_.�κ�������������͜�0)�@��%��QUr�b� ��`�&�Q 1�FÇoooN�뮽:뮺�u�\uק�������̫��$?��T_���T\H��""��,8r-��Qs�H�6Pa��*�b���_i\�DD�����>�9��p�|{��eA}b�PD�:I�
�� ���Q�vUU&�C�(�
(B
K�r9QEj���r�S�P��a�+�4�<*����>q��P���0��y2��Dʩ�D��GiO�ۑ���������H~��er!���Hs�~ā՗"���.TTQ�+�2w)�ԓ���9dL(�ʫ�d�D@0�2i"0J1�&u�V��\7��W�~�g=��L%|2�9<`�G�xr�V�w���T�U [�M�T����4x-m���3������pc��Uq�<xW5H��/��|}{�[v6[���M"���y�ɐ�i0�0[�ۚ��hs	��y)X�i�ߩ�m�Yv��E�2&��= -���iفR�hLm�p%<�ёvc����
K��L�3���x��77�{��`�E��Q�i'*%G1������X��hЭP�n�ZCY������mE/gϺ<��z��${M�k��[��f�Q��#����T+B�ձR�f�9pr�����0���6E����G��25�zbĻH�>�>�f�<��mݪ���1g�%+k�2�H�2i���`$>A.+�]<ѯA+q �1�`3jwe���î�f1w���W��:�a;���>��|���
ϯ�������@Wtf����w�[;�x5^��Tr�Wb��K���:���&g��o�,�H���VE��,B|=ޫ�Or�q���^\ۻ���}F��Mʽ-jQ!�pZ�0l5��b�����9՘����G7ܳ��O	��8�v�j6�cz�跘�tȑ���)���@�0���Ю���źk=�5NػՕ�U��w��& _���p�.�8�8T�.p�,rϲ��Һ���k��g<5אZ{3]�A0�	٨�/�r �D��(�s��Z�x�Z�ݤ7��d$��C��㧫gҮM|F<�o��uռ)R��v�t{^|��~��\x�<x��V�mJ�x�:,�[ޤ=��E�"d��9���|��7� 6�1RVd%f���M�%���j߷�R���}�6W���F�6�Cu��m�X��^X����6�Sja/r��k����}WW�Mo�K�%�����ӹ��	�L�UM>�1lU��+�a�*1���^�b��2�/5ze|�#��"�6> a�Z
9"N7��z��)*����n�ܷZ���[iwt�Aִ
�l����>g��O��M�q���H}Q~] ~3��p�g<��t�b�':��M�ˏJg�~A�P�����{�c���u�`?-4�:�Zg���Ͼ�>���t;�*ϋ{B�r{�s.��F��>xx��I��d���s
����j�oEa�-��V5uB8Y�
�����H5�)��'I�|�f�`e������d!e�H�K�77{���u���)y.j����4Ԇj�m��mO�9v�@�f��t'������-�qץ�UjB���"윈��9fQ�&,S�g�F +�,a8��0 ]}P'nI���<��U[�
iZ.{J�%�3/�ǜ���v�9b]�w�cܢ(�ǣ�9�R�K�(Md�D��f��̮����Tϵ�|\�o�	 MRa��y��\�Ȍ�ݺ��V,=��f�B�n:�5ީ���W�)��{Je��3�+9�-�v��Sٷ��q� Q�
w �����5^-4�-�*�=y�����q�L��$�`O�A�x��{jH �a"��x���8��0|��HK>��<�帰�9遲`[ck��jc�y�x2[gc��,��o�ޤ2�����(�I�Bd�����\�������N���e���N1�٥���ק�r�!5����Z3��FM��|�.$��-L����j���1�]v&m���V-�=�S�P,7dA���i�V�!��W0���ͪ^Å]h7W�=�8�@��{�5_�6���sL33�Н��R5Jf/A�}W��P�Xb`��S�%��qb���|>��U��Nʳ�����~�ĕ�q��L+�So���R���1nb ������ے�'B�`Yԡ��3:��t�Y��0�����䜹�!.�*��.��6׶bN=�<�-EJ�74ٚV[cX�337�:۪��a�tXr������yР;��������zذ-p,O�#w?��M�bd7�z�W-/y.0v��Yn��LN%B��2q����p(느U�!1�zbU3�o����c�8�Q8�h��:Kdӷ��L[�����P&9P~�(m�g�2�I��2u�<Au_�����Mì�Ş�����Yh�1��5;^�}�P"w�t���O&sȶ�fL%������7hS�2�"����������x���-�4��QO���;i���;�Wg�x�o��f�+�]=MW���L83s{ 9�eݤ�]�6
� �G�C � �=@ 3{����%X�>���yd�r�_t�H�\��]�ѭ�
;bGR�K)12`���ܸu�$��$f�oy�YbV�51W9�Z�-\�Ͻ�)�ZM�%�Kϟ��2�UGK�5���|�[�P)�����M��d���:N+�a=32��G�̊��y�P�hOG6}~ ���i��m��3�&�~��ը�q0�Y�=˾����)��]H{Ƒ���_�a�x[��wrU��9�-Q��=2=�i|kȃ��a"u���'�kֺ����N�~/�������ǘ�t\�)X�_��-�E��J�[�&��<�/8�[���S��S��}�C���vbؼ/g��Qm�6 ���`Xi�W%��x�t��yw�jh�k��m	�82��6d��!I�Bjϴ��0/��-���9���w�[1U!�Ì�0�Q�m}�Ș�f5aV��u�}y��yfL�~Y*�5v��0�r�}�P�2%�'�t�vέ�Q�:�c���nN�>>�o�{GK���(K�y��F(��o��0�+��[�>����x����[9s�ORۧ�~���:d3�7�K��vq1km�-n��+��&��:����e�+> ��nv���o(�S�ۣ�H�٥�]��y>w��vLԏ:�3Y�Y�mu��2%���-�0l#��,���<�^_�?/��x�ǁMe_6g,+�[_ܷ,^�3�%��D=�z�򠕐.J�(��H�>!��X�=?z����:�{Et"g��6��Z��+{b����^*s7�3=��H͇dh�-�Q�ǀ��puEV�t3��(f��- tt�� ��M��'5X�z��[�&q��>�}w��*���J����m:� !�#C$�f6Z��1��˟�%>��#r7d�d�w�t�uP����_�[�����
�N�Kc&v� �Br�v��+|��O�-�c0k����Չ�(�C-4���o���~�C��2��#zJ��K;��P��1�� M����1T�툷ٻ�*��O�{|�>"G����R��1h�>xz�b5��̔�@� A�(��Q�L�N����Iͦu����a��oGs���O�H���5���]�����ןrm�:�~��//�q���\�I�%��˕���)'"�@���`zb���L��I@���U! �+GWu��S��~�8i�X4{�ˬd�9h�Y��<�r\1�_����=���B����"�P~��^$e�_��;���ސ�r]�SOM�x¹�f����{�+�X+�cjc�#1:q�� ޜ����x��M7%ʹZ��W����s��w����FVmX6�`�Y��o:=�z�����92:ik�D�Q0��m,���ʶ��Ǟ��;ޝ^_�����U(�dtq�I!��5yH�D�x��[�a2#�u�����ﲙJ��[����n����e?�\w��M����a��a��wP�s����d��2��R��Ư�{�{۾E(���o��.���`�{�����gKMf) 'o�a���5M����rˡ
�5���t�T�5'��wZ�Z��Z���)�?��1���'d���o��P�^5z�?����edm�+`1%>�DsD񐏫ﮠV-��H+#����e����,�=��y&�iz�B��V?t<�k)�x��3l+���H׊�z�J}���U]
�[Q���S���z�k<�4��S�]�0��t��O�G���<;�S-�%TȽ�{=6�a,�oZ'^�i�r����03]��{b	M�8-mm��i;<�z�%��J�7u�=Ì�fq9�&�*lZ�^�3��Ņ��/��Ӑn�8�X7��ꅮ0�6O��E�6`�t�M�tEs�XF ��*V���������la��
��6<�Z��[m���t�{�/9$Tv���	*c�7��u �zۼ�Ep�2uӓqq��5wz[�L�upLT3�P�D�A�,��y��ߌ쭮�];�go�L�t�nGn���6�셁�z�:}:��n��r�O}{x2Kb\垵X*2z�V�΄|�ר�'���F��o��[�(p 	� ,Q�޻��{���36��m�_���x�k�P�\�_z�r�,<d|�&�W��.9�⧽��cȧ睬�Yvr��^��W�!��g��d
+�G0�2z�@j%ke���Ѿ43/041�k�p��TP�{���x>y��T�|h	Rt�y�F�|�s�5�q�v�c["�e�ܶ�0�[�_��׈6_�X�`n�^��U+�|����#`k6�.�Kw��FI~pt������7�>�7�͖Z��4#��H��9�/��,xPS�ϥgf�aClx6��X��8��z�Qk������o�F��:�`C�@�5$s�Lq�0��y��*7�(��v�U�C�󞶌r��8����g�GP��}H���:.c�k�	�ϰ���χ�7}��e�����j�[�=�9�^����7i�0��5r�00
��0Ƒ��C��O�N�Bbu�Bo���"U�y�PA���Nn0qJDo���>NTO��N�a��~L�������Gn}���*m����h�!��;5��J�"'O1?6�7B`i{�o�[�:Ϝيd�`��>�;�����OX�	٭��nbC�W\U�B	[ՠ�<j�;�)�-�_UU�8���ǞD��7���'�αc$��-��Y�7�TEi5X���p�L�ׁ����f·�f��u]��}ϳӻ�T�rl��w{g�mtX^��1os�ߟ?�o���>^�x�3ǎ<F� �(�)V�Z�.�μ�����+����S��������<�i6�暡�5�;��{9p��R)��Ql��Zt_�Y�K�kb��٠��-pjO��`�����2�h��۬=N��k�0��R+4Z�a�\�r^����P�
���d��3�;)����l��΍�Y��!��a�������(��H��H��9P�{�_?����l��e��߷[�E���C��E��!Y�.��G��[WO�1�[g�vX��]	�����@�>�������:��Ϟ�-��"]�@����#��2���c�N�^qصc]�s�(Zm0	J�� �ϒ������K�t^�?4U�v(�]�gO��y�3����k��)b�_�ӦG��Q#p���@ͯ^g,�ӹha����cT��_Zn�sjYw3�v�M�{��Y��gH��j��}�>v>Dl"@i���#+="DV�Y���x��]Z��Z��ۥ�o�����IX-����7����,3@3;k�|�~�	\ƿ��U�?(����T'z�?ߡ��wO՜L��({Y�����������&�V5���n��L�(eR�ǽ�cf�:�.`Q���6���C��G���]��:�3���Aw6*޶;�a���N��삋�b[��U����{��{~y��ǎ<Kd���X��6�h���������d����F(��g�丰�rZ��Ƅ���-�S�R�M�K�3*�3|���!�ȉ����՝�`��g!Yz��/��Q���G,7`fš��V��_f3I}�e.�a��*�� �y�� �����q���0Y>�i�My̽r��6�3�6޿l��s7�ʏ	�[�=IxG�m�?KF0���`��M��Ɖ]K-Q�>OM�)㕪.km�"7 �v�ݒ�x�;4C�R��TUЬ�U�3��"=��,��|oR�0��^Z��#V�F���5T��vy-Me�~�����k�C�ǞbYY��qQ����h�h����7�k�,���R��י���Ϝ�!]4�ձ�'�U&����Ьy�}���8�!�όwҗ�p�oi���ƞ�^�7}Iy�A퐃@��:�S��'Ι�Eˀ��Ժ�d޶�3~i "![��յ�a�e��*� [*r�Ҧ41�tf:hÒt�o	
I�Ԙ���9�̕��۬�WUt[�M��^����C��\�����?���HM��O%�Z2$Y�.?E&T	<j
Ψ��^�2�h{�IQ�)e�=�o�L�7p(Y�\{M�r�%dt���̇mT�M7�\�<�Z��A#ܝZk���3z�'wKg�u��w��4}; �7��lna�Ň��Ì�
�Ԗ�{2T0ܝ;;/�Px���{��^���%�l�Dٴ�[m߯�ӥ.��|@c;��~x�a!l[kP\C֥�d�燪[�&`}���n;Z�y�Q�Փ����yl��*)��fƧ�y�!�����i��Qȝ�LhqI����b�v��:��N�)���4W	G�]��g�v�^YHe7����nd�E�RM�mj&1��`���[��DsŞ�r.�oV�5x�!㕱`eY�/�L�y
o�0k���O�}N�DCu�,��qAFGj�j�0�^��>WL�������alV�HY�zБ}��.cI�}��~���f�oh�_|j=��)N�V�:�q�ޑq5_U|�����8�u�����- �B�o��k��:r-[^p���ܫ[щ���t��BL�o��k����7/�z5�� ���cumF_Y���nV��<H���	��hkH��Q�.��b��ZK)e�D�u6f�j	��s�1�����
>����j���2H�e�ᄠ�%%m�s��ޘv�cƌ�-��ٺͪ�m�Ny�@ꕕ��D������.4�2���*͋�YS��4Kb��v���\�����Ku����T�z���anOe�1�8��"��͈�g�M�/:�NU�}b���ފ�_h�γR[N��At��Q�X#���n����Ү���56�Z�GG��&曉%}�I\�ݳx�&�6�.B��(b�.YD�[��f�U��R��u嫻��D(�u�
������2�@�|�e8;2p��T\��õU������̽�VA,G%��v1v/�"h㭞Vm-�:v�)]�uҥPS�O_q��/�S���v�j� rkm�Z�U�v����*%�u��t���xk�R����/:�;��mڋa�d�;�w^@rڒ�q�����[5:+���ˤ�N��&p��Ǳ>y��ɺQ}Np�Zԫ�i̻֝��h��u��*�Z ���:-�ALI�76uF�5w�����������۾��"��z�E��u������\�U������ҷ�qӢx��K��z�_r3���Q]WOVұ�A�] ӶG:2�fҲVMo+���o	"[h-��PZ5�����C�ym�_]��w��Df����(��N6�2V�\o�Cg�S�ײ不{T&�	.���5RZ���]��ə���9{��I8�i���\CȽS[�U�b��8v��V�k�5�����*א�vʶ�=�=�$��Pݱ!�o���]ǻ���)s�fӢ����ix�MY���hӏ��w�B����׍�O*�WA�;����
nU��3u<�Ȇ:�	�2�U�PŸ�.���H�HVؚ�a����+bp��E���������r�b�:�"�
��U��hk̼���<�a>'�Z�Y	�L�#���`=:X�iA�e3�bT�3��x�t( Toqpb����Ҕ:�t��M�YQ[��Ȉt.�,
o@u�S0u3��'Yx��-�t�c�#��h&�Kۛ�3���a���VRy�8o2���9�k�F�>�� �;��t㜡����uv�	�
q���Ȳ�Ǚ"���oh��M���fVRPp�\�vY���f�RN�ۨ��"rGy�^�� 
�����;�2�p|�P��gf#�M��V����q��P�Օy�A�Q�l�-��c����f,.�7���� ����e,�Y�K�F�	���\�����N��x_\E���\9�T��ݡ\ � ��_-t3�F{�U���3F���o�Ԣ��wV$fgM�Co%<gMv��no�$W/E���n��:$��G&36��Ww*M�f����'K�TT1�k�Q�pW$�u��KZo{h�z���]ֱ]�{.�hGv������2;�O�,�Ţ��g
��f�u��wd�M��������'wpyے�^�	��Q�2�u|���r�����Y��N������s7��A�5%P�Hd�
-�Q�K���l�H"�th��IU
Y#E�"c
�I�h��^8�y}%�f�{�q��<�UD��P*y�ܫ!�X��B�2d�$I"[���Sa�,U�;I�8\y=ǎ�����Y�ks��՞�����O�����{{zu�]u��]u�î�㮽=����S�@���$Gy	?�A'U���C�~�ʂ���ʿ�淏�����}���u�]u��]u�î��q�11�TL|F3��
!4/J�����)�&$�o0 � �W,��)��)�*��\Uy�ʟR虄$�'�?#��J�z�|BUw�G_Rw~��?>h�e��n{�
ލ (�Л����<�)��d�t9TU��3���A���%��	C��SJ�"/�T\��O�ޔ�J�>	W'�
.��r�+��8�n��>g�.��"(�OF�y��˿Wg��	�^����=\�L�B�����֙��EO�{�r?>��ϐ~%�h"@"J�3@.S���#��q,��F\�;z���R���ԎnvV661�w�\oa�o=���f0˝4j��dX`�{Eb*^|��D�Hê�*���>��3ǎ<M�e�[I�����|�߽6��D�I�m��! �S��ٸk������}{�Z�fSbĪ��'�N�6�����^?]5�P��Fd��K�D=h-�u���.�z��FE�=x'ИZ�B;�ndLQ7k4˾¶��*��5���Z�Ob5<5G��bB��v��}�`��H>OC�n�g��p��L;sD �._%��J�� ���ڂ��J�Cӂ��(���/i��c��'�z��`��0��%X�	OyR�Ӟ��7U{�sI1�a��u*ξ�w���8�OVZ�֭���d����3��<hv1���.=��FX��1����?��x�?{˳:�Á�)���L�_�Rt�Κ5�~9]�cSU^�9~v�&�����;�K���u}ײ���� �ه�	~a?�)<s�"�yK�0�=�W��)�ufl���g��굛���T��>�U��]�󂎬	\%�~|D����Y�g��0qfh[(L��~�ٯ���!���vT�������Cmx�j����h;G��sH�����;�x1�Ϡ_t�=��ݦ���#Y�j�L�뢮ڸ�)3����G]Eͼ8^dkN�w^7oBA!������ЭYR9|��9��`E]�ꡕ�RH3��7xHm�
S�6r�j�š�r�IoTL�`�]��=
n�� zL(`D(`�-��Z�k��M����Ǿ���z�5��J��{�6��4�D�
��Yhr�s+�G*KI(� U�0��B/ݬx�����/�{G�ˁ�O>�Ҳ.���6�!�y���ӊ�C��O^�f�j�	̓q#��ne�K�מ�SK���V"i��:;��X�g��;}^'����(%,���F��ϴi�~+n�};���6�9R[��\-��E�,o����+z���z�K&�6`�9�Gd@y��OvNv�үi�}�Y��g9�5o�i���G�c`%��^CNV1�WԼ�����kM��-���{�us_:�(��gdQ�(}�VjÃ�Z5ivAp�|�٠���ؖb�����g��v�0���=Д5*`�d�qAI��|��f&����{��Wb��
qhg�q��%�ǳ���-|��k�0��P����Y��@�74ͮ9��)>�J�������P)�v���Ō�`K�؊�s�=,	�Z�.C�i���]ҍ����;�z<Vd�{�5�NiGl2S�����7s4�t�jwv��}%ދ�?r�_��D� ͊缪;.Vy�`J��DՇͥ��3F;J�u[�}/��0T�`�p2�� �n,������hn3�<[�t�3�e�F6��J�h��V)�U-)1����R�I�7s�qm�k�8�y�eT��H!�wHl��y�{B_���E���2Wd����٦eV�=� bb��۵� �l��Ȋ!���>�'����G����B�̠�Xk�$>���%�^���ߘ���#j��4���j�����Z׎�.�] ��w���G�xK:��/����U�ٕFz�SS�{Ɇe*���m˫�#=�3\bH�ƥ�"6���v��Z�Lc9z��ڇ�@w@��t+�:��U�9^�z=[ gP�_NP��6�	�a� �oeY����48�y���ڸ"��߭���ȔY�|��*���.��$}C�zm�ƾ͗,,6�KPsΞ0q{|�p��w꺕�ֻ�Ŗ�d0$	�p��ۋ��pG�}��m�2;\PNYy�P(Af\�͝8��ޜ�YӴ�q���G�y����>v�$(����I"�54��m���ō��F�~��m>���������1�h�`�]ފ��T�:�?��`d����j�Ύ-���Fv�.82����A7B��V���q�$xqh�f��D�rig��_pA}��^�Ȯq���a�S�v�@�=�՜�Zr��n+2Vܶ���1���7��R�_�C�2-���G���Iag]�賸0���+��E$�L;�9�b�(hE`��������ȶ��M�t$�M�����a%뮩E��ޛx{ns�5G��+����B����z*9�V�fn]AaFxr �zF�F���{�>>�u���ݕr8S���f�`�u�8Um�.gc.>ߙ�vq�W�7���@��O��ȜJ����1��(r��z�W`�0q٠�i���2��s5�W�q���V@!��o��S�v��P�1L���py�w���f�w4s�硵��Nld�<�"A�ý/����sRմ������^S��l/A�zS	Ԗ�>��љ��C�������J�׆�����Ayqg��Mr��Ա㼪1O��`D�6�$���smMZ8�b�E�F{����wP���"0�����Q��3�=P�/-�̷�>��/C�{�B��y8�l�zJ;�҂�Bֹ��f�g�6���&[]s��TPw�������Щ�O�%�9�P^�J*Ml�p�J�͌�F-���������nنS�㎇;!H>�C_�� �ʥak��;�Ke��}z5���"5�LVX8ط������e����j.�p�[ڝ�GbޑX���$VB�i��w��H7TG+v|�Tn�HW��r�֠�r�:�������0��>��L����GPb.�* ���s�.�Y�VK��6e]���uU.��)�h_�n�Y8p��wmRou��u��;�0B���T�����G1��I<��.@U�C���Ec?��5㘯�_-ڽU���f�!���*Y�G�{�;f��1Wp;l=6�އH�k$%Y;d��ǩ��ڧ��Ǜ���{�q����8��8�6lխ�e�[��L�9��Εj��p�����;�wÈ���n�Ba��򮖵HI��..x��tT
�����ӻ*����-���^�/�y���u���o	�)�=���#e�5�rp(Sе�料?�5q��O\V#��ƵO�)�z=x�&��!2)]xV>��U~��w�gT��?AO<�[<r5��_~���Sv�Z��in�.}��V�/e�iU��(���πkC�;+�g��Z6�C�����M�M!�Z{���A>P�Ҹ���%����A�S�����Vf�(�6�;�aDz��K�d�$7�I9o���H�iI���r�]х4����=�_<��O6��F-��\o��i�3��3�px/�cǞ��=w3&�{ۻ�&w�?��S��&x���O�iG7T}����"��(q ���/�ķ�)����^�Y0i��oZ�û����>�X��F{�J�X$�]��g�G26dn��Ն �w��i�OMt������$���^��o���	NȐ����~�m�2%�R�֮p�D�(�ӱ�c��?O�/�w
ݷ��2����zlDq����O��ÄM���NK&�a*ѕ��;&Xc���[�k�t�c�ڠWږ9�h�K�#�29���Y��4��%5:�Ԋ:����Lehhѵ)F�9ɩ{��&�[�bx��az���~ή���ٞ<q��mjֶ$ �b	`��5oI�J����*�~�!�w�����:e�M���m��mTW��l�I�Pd��	9{�X��D\�`��D@Ə>�"]JOr��^�#��b�C��~Or��r ����W����w�p���k*�zYk�YG�����
�^�G�+Ghμ̚�Y<��u�����|��������DH�9��� ��p�O�a�n���8K���<�%g!Y1��:��^_�g�C�-��Bl�vl��b��s����J����d^��ͯY���ܰ�L��l>O��]C��"@�2��Y�4�q�=�Nr��\��8PmuV�Doľ�bmJ�d;n;�i��=0�1�Ά/�S2z�1-�YZ'�T�~]�_>��Y�>Dxw���(nN4�P�f�.n5ȓ��>P $����bݳYkyޤrp'���!�c[Z=�4��d���ȭ�'�5火�T�`H	ส
4��[�*��D�P�:5g[
���P���Z�M��ֶE6�k�~O5in�4|���L_}����g[��!�)�"��2q�`�\.��E�"[���"3����{7�i��k.d����s^��jR��V��SU��:�Y��%���\�̧����-��[�ث����>�C��w�b�n�ۛ���v�<����z�8��݇g
�L��`���g%��[JW�Lw8����¡1 �*�؜^��+"1�O&p�^����k��g4�k��_�f���䭟.�|K�	c>��KX�|�μ�sÕi�r�ͷ�2-���q.�{I�kp�̑=�BP��� ��m�K&�aڻ 7�wU.s�c�~Q͸���\�p㽧w��Y�_�U����r�BW�}C$O �j����z�e�d�]W�`B�OJj����.tX���Ѣj�λ����>���%ؘ�f0&�/�yT���{�?4z�Ȯl���&�o̥P{Kp�Z�F9�]�>� ��8�Q�o0�4;c��E�[t��LZ�ڌg+Fc-��s�E�u�/^R�D�z9w�nx�P��쩛��3޴���]�g��8�ͪWY��
Dt>�ǹNͧ$gtz&9��3%���/Ϭͅ�+�n������Z�E����UH_Z%x�=�>���$x�-�g�w��-W�z�BfQ7��'�7:3�-��<h��Hu>��C"i��,�*0]�X������\�p�(S��я�v�B����ռ*[�Xܔ���b��P���������[Δ���m]H�Ir�U=���/m6nU�n�*�H��u�����θhaͷڍ�ˆ��o���a��s�z�	J�Ԫ�-��rn�߁&L(�`8p��0H0 �`� ��Oo���FG���z��m��|��~��M���<�%U�f��|�.�s���}�f����U��w��D���Ĕ���BzZx�J1į�B��ء���ZU��)���~[���s��P����W���L���(�c@��Y�q���Ɉ~�v��=�C���+��q�u�1�O}�?+<O0yv��y	�=灊O����Eۊ��jH��mT��oS>���ceS{���:.$�f�S���	��=����oؕyu�+�;����L�n��ЌT�9�j��~.]�3�����N3�eےh��Z�[1����2.yZ�{b�Պe[rͼ0ҽ��v�y�
�|�a���{f%|p�����Ǉ�Ƃ�x��S�mV��G�T�qꚷZٮ���nOͥG[�?zQfcUb�lt�'�%���T1O�G'n�>u�g&�����A6�XY&K%�ฮaAtcsP��x���4�A�"�/V��o='ݝ�^�u|l]��/�c�����~FKg��5ηjEv��G�������������K8�sW�wL�	��`�������縚�y>վf�y�<+;�����j��v�v�q^����f
" ���E$�3����k,�:��S{��dq�\d'����q+v���Y����BƢ�ټW�__
�bCܤ@
mȩ
i��i��l�sI��4W�!�@��I��A�[���>�{��l�TH;|A?�Ǽ�e���J���y���{�J�v	�>���9�MiŶx�ʠ��K�:B{=��N�5A�<������aq��sG�)�I�Zmo�0�L&�����9{�w�U�]ѽ5�w�%���	_--*��gN|�`�d\XVzE�p�$�6����9ɦ��ն�g��4����	�^��Y?��PsrR������8>�N���;�8��G���Zm��S�}�����r=w�ƽyDs�$.5����<'�w��xh6������o-"3nbl��zՀ���!tBt�_P��N{4s��ƺG>�S9=�����Γ�����7��Mz�z\[U��ͱ����!�E�y	�x��X���k��q�f��S�q/��^y[���kb���N��T	RϹ���P�2�Y�e�U��I��J̰�c�7�o%�v���lh����[_G�/�0�ڐ�(�y�-�y�����VnKMv�g)��Y�ysf:/-�ԖT/nԌ�y��q��[��UA�n����<w�R�aV������{]wƣ����m��}N˺_`��T�!X�Ϸ�=������8=���I嫯���ӳ�y�)>��G $�>W��m��)u��[U|^���kS:��(P3���O]�A>R�W�I��#����N����=5)�UH�O���@
�b ��o�'U��b�Ϭ>Zn����4�k�IxrVǗA�tV>�����l����ɭ�k�J�2z}=��x�󴼀�y(��c�t��zv���ɿW`5)�)#�8��M0~���95���ˏ"��6�����]~�.(k�xAN'�˯���7�]8�i�M�ʞUy��ܸP�X\DޱS 6͙�.��5�-Y�%ܶ3��>�����R�w�������
�[�cAa{dH�$��L�^9*N���qVn3��h���3���Z��2{x�n�Cb�.S�#x\��Aò��^�<����n*�a۳KE�}ޟ\��9g`� l]�=��#|>�;z������RZ�\���m�.�LXL=���F�&�H�4M��݅���֡�%#��[mw)��6��/��~;I��p~A���ɿǟ�a]W*�z\/w}65ٷ'2��(m�>=�ޛ�9S.-,+>������NM���~�ނ�/|Źv}����q��L4���
� ƀ=,�J���= ������z<�uVHa����3%�cz�N��Z�"��uUٝV94��}�E�Y�PF��1�i�id^��(�R��PM�^������[�P�9.H�"u��[x����s�k&��+�Cr��*J'�J���PVz�k���DJ�1�efP@pՒ~]�pw���j�3����}��֮�.{to�0a����4SWZFؾMfʢ�Nf
�3hI��Z������o�Nv�
s�csc��Z��\x2�h�B�&�QYr�'����"�Z��;��!v��^]O6@޻�XѨ]ܚ;[�o��P~���g�N7���Nl������>Z`�+��؄��=wV)Z�R�F==5�fu��'!"%�c`���9N�F&�}$�kwO�/S��Z�yF��Pd���P�Ž�*�\�!���6�EL��=׷~X���nH�b��@.py�}nT�EH�����6;�̯	t.�#k���j���KǾ�1m!zT|%�]@���j����V�j���LٽŴR�Mo�r�*�[��W�z�|M�Ý�0:���sU�H�Xݝt��c5�Қ97K%$���ݥ����5��k���F�Vq����&n|�i��0O6�:u����l��Ɩ��ʻ�����t�W7�j��8���`��΍w]o�V㓫���-�[K��
YU���CHr��}�Sނ���YY)%{�����(WM�I�L�#�t�I��������&��X��*μ�=�:VP��^�#��<��c�p�&�����m�im�� ���K�^%p��\����p�����Τw{�Q�K��j��̔,�.V��u��Nd����2�X��dϣZHV�u�>*��	��Zp�>�R�����Ю;��̶�:J�z:Rw��a��v.��tU���w��]�s%�v��dY/�T�gdB�3��5wҩ	�p�0��*ή9��+�+�θi����\
*��6����E��6o-�!���9ބE�]D{�fl2���u�]���� �}��vv�J]63��غ��9�{*�\ ��94�΂3W���U�U��/j\���h H-@�%:�����ºާk��٭GNf�;�>y�;<A�LY-�L�e��]���*�q�k*H[���ᮻ��'D[�i½���S�yN�PK����L/K&�w�tP�xջ���:�l��yF
�����odo���^�Q�5�l�����3Jp��%ծ�5�ۋM�r��QN/�Ob�˗��F�|)�tmX��b��86N�����]�*�fN�,�]���։ ih�k�7�+36tz'd�Y��$���X��LV�6�s';����KL�'#���t��,�2HY�sZwj���LHC�!4�O�2)�HY�#�p5�\y]��Ǐ�����}����]u�_��N����D�ё�,��0�F ����L���Nw���~���Z���sV��x�����}�_ooou�]u�뮺�뮺�ק��������Z�rI!�#|��M��N�w��y��w��������q���p("
��Wt.��AE�S���~6]ԧ�>��>�r��~��[͗"(��{������O�|xz�A����O��
�
'׽4�\��	�q�/؝�/D�*��WG��'��C���Ukd��?�I䄝��Z�r��y�^S�����A?���{�S.?Y���Rt�~�-���HL��#�y��[�g
��ܿ"�k������9��d\"N$}b�R����+��ӊ�9>������=e�]���7�v�h�H�iR��k���S��x���� �o'uܛj�/��'�����U�FY���3N*i�[����9ؼX� &d���q�FA�y9��k�=ｔ��=��r7�v��y�kY�@���Mu0'�b�\�.���;���CIw�Zi�;{�q�(�y�4��i�ץe
�Xb�e�0��.��,nC7C��(	�Kޗ�1+j�棽ݺ�L�O>*"�1E'����m�V�k�(�{�ۻ��h���S[7�k`�p��z�0����̎�`�S�"���+��k�e��ē�b}ꥏ�F7+�^ժ��ܶ���#c�K��jE��z��m�ySd�_a����\�?��fkT�5y�.��}Wʇ4�9Ccx�}����9h���F���ی^��A�2���	_��>7]�$���T(t��6�<�Ef�I�ػ9;zo_l����{��)���Z�c�A3~���Ǿ���/�\��R��K�X�%�u\WtźֶCQ��1�hX�M��������5�/@峆�N�觶36���Ϫ냿H�+D��B�	OW�a���\=�C�2ǽ?�5j'�8�^MBFcDp���X��{6h����{���|�ú� C����G�W^-b�rO����0�~������GL�=�Q噺�L"�i�C瀊y"�-0W�;;��W�l�ʊ�F�fuA7u���R��u1�y�ؖu��X��Tu3xoH�v�8�bQ�C{���}B��D�}��}'���O����ȝ�%�Y=C�@��j��zg/��6�	�?ǉiW}3��;>� ��k�2CוF���c�F�>�P�sO��0�Xg�З�2���}��y�U�^r�����f��+�,"ǖy0|zŲl���}�]#+^8�.+�^{s�șW-z�j���ލ�Y��?:�}4�5��*q���6{�,(UMl)�O���܎����,Z�os�P[~�iz���=�@�󦽑���S�U�"C��\;�P�B��7���Kk�������L������`I��l]�ۻ��P�¿T�9��?H�{�{����o&���g8�r��{LSO�?0�]	���b�V^����<�=���gj���A�w�
���8\�oR��^u�@��[��xMMCr{���-�E*�q���v�nc���{*�$��<lçei�7�*-�����),���[�͞�C�|����[b��t�k.u�Ι�MtOF�d��VNKз�qM/p#4�5C�G��А���3X�j��=p��5}�|�}~��R��&��ٮ��gp�+U���c����&�#$z�JQ|�=�wr���KdPd�̖t1E؁�`�$�:�N�������}S��s�:Y6\[�����J��\�E���4q�N���6�N3�om캕T��r���m�_织�%��p��6��j�0VRǺ��w���IrH�3����;��lu�udl��[V\�2փ���ŋ���.r��
י>�2�C�ξ�g�,U8ܟԦ�]<�EJ��f ?���g9������K{���\p�Y�{��zˤL���N	�<ü�6X�e%���mj����[0O��<�G�kx�@�-����DF�R�5�ʅW�Uqqy������ZRXw�v<W4�f�+5Yi���<�fb轉��� <�Н�ob*o��OTc����,�ͪ��O����\9��,A�2���~"DCM�E���<i�98��-}o��C��W]����h�F�@=Ba�tl/"���CT��>�w���0�<9^xP�|��&|�^�j��S�s�ʷ��~.1� �TZ���w��|sB#��*p���)���w�,Au�׳ef�X	kB��z<����}k��½�W�T�3��`4%]-j��B2�?A���Ϸ�9~BNW��m�K#�$M>����m���-��SiZ���|���Ԃu�!�GF�^w={����3fX�4��&	\z�v����y4:o^b���@���}yܝ;[w�)l6��.�<#Rך+cF���>Rsk�۝F��7MrEr��o<��9HV]� �H��т#�́U���p�� ֯)e���� (P��!�U����e}���I���h`Z4TSAezt�<d&U��V>�h	��4a�����O���آT���Vl�󳡡&�<��Y1E�T���P��Q�e�b1��[���py��W�������勷����G��W,��kj��jzNe-��+/ºOJ�ܲ�L�]�n��ӂ��r ��E��L�c�q�5l_L�uQ��ƚ�n�66[�b����q��k�ӯ����@:�N�XJ�7rSM�k�[��\���hw���=�V3e6�]UOe=�ۗ��CbBh�q����<����4<��IO������Ҡ;A�p��`��Fc^��UY��}x�AAI^���ή6'Y�YG뮞oM�4"�L�7'�Q̺��F����~|lS���J��s�5��[|�E���r�B�	|w��k,_�I�^��]�%�h�%�~�����]��[�ʾ����&�C�y������D�1�z�U��:lL��
��ƴ�����.�j�d�C�.i����4B��oy�*"��,�[�įya�)�j��H|�^~:��޳�.� �,��N�H�u�|��g3�ͳ��Q@X�Y'Z�Ue����rf�4lP�9ڹ�J�U�e�5Z����Eoj�5��$���
؇j8|klc�P�=c���]ۇG$��wQˮŇqNW(�f\d��\L(�@p�@ ���O����q<��~��tb�z�Ɏ���e� X��"Kd�`�o�\�Q��-�r��Okb�o���9�O�n���-���x���8�M��T�6*E�Ѱ�u�z}?]?%��r��d#zu�K��c3b��ezF��� ��w'��8΋�/F]GH]^��U_����J��f��beă�⚳����N�ɑ j����a�ۼ�ϋ�$�畛y���iY@��q@��]�O����N�)��K�!��*N*`TSg�i�i�ǎ�s�l���;&�vw���Q4�y�.�Q�v۞T���5e�d�B��������ߋ���#.wcU�os,�(1k�xd�U̿��{(U��L����VnO�"� �҅����뇧ۦšF�Ȩ!x�So��[��(�� ��M�T�=�N���?vп�xv��ߍ��5~fH�{����V�'�<�����B���/K17����$i��cƻ�A����L��}��ף��1~�ba|��mW	Gt�h��W�`L������;b�&'���[�Ϻ��ֻC[~#�>7WD�i��ͫ	㼦}k��ܟX�����nIJ�{
[�p��h{�c���hY�\�Tya}ZU��J;�0N�oc�ӣ�g�c̬����*U;��o�\�������ۮ���^���!FB���B�!ݍ��_��?�C?�~b��1�u0�f��tS�Ze�}|�wK�/�͞��쪣{�a�^��.�s��En?C������u&�fB�0�(��.���<�-@�m�_8\�쪩�J�鼠�1���Z�S&�FK/b�a���5�CYA>ZF?>�P�][[���De;�[Hv��e�|*�����L���5���>/��:��_�편�N3Hn�ǟ�W;=i;WW��.��R�V�z�.tЭr�]�1�:a��c���w-Y�჏-�Y2e��Ӥ� 3�;��&D���<M�k΁��/{Ѭ7�<��빇K�U��ʴ�}����"~�L^!x�!|}"�6�>�U�/m��^Dol<qr�f��O����\�UΒTl�s���lѳT�~-������Ng��I5�{_��zu��H{f� U�i��u]mNCS���[���Ī�,۔y���\��Q�r�T�@pst==�A��M��8����B{*[_P�{�E��Z��-=��,��6{�����Ll��Vp�6<%����W�:��w��V���)G24ݴ]UnC1	Ȅ.���(�X`���+tި�����I�9@Wmѡ�کN���i#�ԃ)�.Г����vv��7�t��u����4��#��9��u�w��H�":(�
�]п7����k!���}�~D}j̑c1ј��y�И�R�i�S�%�\D9P�톜�9t��Mx��3���g�Hx�>k�^q�F�&����qޤ�_=���-���*o[��0ӛi�wP�0��v'Z1�����*
�ȹ����7t�O�������)�<F(�cn�-D��3k��(P�\mN�
1�A�V��ݱD�5��2Ge�6'8퍕X�U�n)�f�蝳��o�찘�J|dRYclJ�ɉ�t��g�y���A�~�sּ|�Y�^��ec�	�v��έ�!Ɍ`�5%����}�ʋQ��/ϋ+�8���|0|��{��jwn޶��%�]�E�e��&��z��|}�O�~�Gj�B�s�����uf���{��6�7��8�DB.�T{�)~�<\Q͘O��)���I`�m���*��VpO~�/Kj����� Ǌ���ܨL��2ϭ����"���8�b�⎛W��<�����N����k���>�7�z��,ސ�~"@�@�7�.h�e��BIw��~Kk��}�K�ʱL���Sv<T��s�h���k/�7F��~6���m�I�2�$��s}�P����gmf��1�����)�;]��p���DۗYS[Co.p����p�.�YoUZ�]L;芕}�,F�v��I{�i5��T^��ã�D(P�D~���}���5�5z�[)���X�z�7�P���L�^|�%�>0�l���V�Y���ع)9�P�R7�8��O��6�mƦL)����Fk��=]��pV�c]��s��Z�����x|��wm���Q���B8�
�`��m�=���*c���Il�9/�mN�j��|�I��6`D���a���k<��� df��,-��Y/84�<hGS���Ӻb擷$�-a���E�sM��n*y�H��%H�Dԉ��&��;��F��؎J�!�kӽ���-w���1����'�߸��_�3s�~Z�__���fs���(�l�V�xRG���yT��~׎=��6��^X��Kj�q�1�h�	Q���*���ʃ�W�¹��R��A)���Z�Z�-ہ�[���)��]c��``{a�
�^��n�66*b��D��4.�����;yD�\`!ze��(s�t���ݼ�n�X�����c´Z�Q��0�K=���g��y�	����W�A��>��8��?�����J���bR�P4�.-%l5��p�&*��4d�Z+f��̖����݌t��n���X�5�u�v����t.�#kej�(���z-���(-�I"�;�ep&�a��� {�;�c(�Gj+T��e�6qs �T.dD�{<��� $ӛ���3$9A��]˦�J�׏H��R.Msz���hMz��;��s-�9���YssYh�|�Ǟ�1Z���#�� %��*��T��c�2���%�dsk�9�!��yY�[e۔5v;�f�ݹ���Uu^(���ƙ��g0!o�s�L��ޞe��a��F��w��+��!֒���`�ۑ�GxK!�z_��7�Mb��UW����^�[��3PӨP2}��SH{#&t����\`��U���.#��}V����ng&�lb;5	����Co@�it���{��yW����4a��+:��7�v0�ޢ&ĜN�n��&3��}:��>�:�NW�#���r6�ʆ��W�C�tćá?>#�p��jj.]'�>�ie��N;K�_������3b����,e�"w��Txݿeg�w&�=[�PgĎ>��g �7O�w�	��m	4��4����#�{�	�Y8�T�w���M/
��79/x5e"$w���9RW򦬿?)V��,o�ߟ��,��g��L��0��;75kޗj/]�}i�ީ�q,��݋�[74���,M�p���� {�-�➷��*���8D����wJt�Ϯ`���].p�9��i�_�րCT�"n+������
_KL-܄��5�!�*�{'o��$=C�p�G�(�+���,�[�G�(5�`�-^�ɶ�R۶��"oΚg�>��%1j��Ǿ�D�5�;��s7cD�ۿ���Y �׎��7a1��6����!�P+�|gmva����-k}�g΅�&n23ܭ��&��h2=ׇƝ�"E�׶'H�Q���a�Uw�C{}��2X4	��Ul1���ՙ��o2L^V�7Y�u���K+#t�z`�|���&����zx�.��ł��&�%������*�P~#X�{nAB{)����t��E��&.����vM$ö�ʑ�g�&Ul>T�.�s����=���F��GlSCk�B�,�Cl~U��k�隣��_�}E�:&l��]�'��˕I[�`ܒɩi��{�aǰ�9P5�A���N=8E?=�X."ۮ��Y��j#�����<ӡN�/���^��m��u�= l�Ɏm��{h'����6&���������O3s7�ï4�G4�IGk�y�F���qn��G:DmU� ��w��дk�ll�<���8| �EL�Hʯ�LZ����*���23��&������).���Xn��Q��#��~��V����g�_[��Ep�s��vx.����R7�+�x.�0�W���zԵ
D���r�ʮy[1uel�;~����)O.0tp�7�-�;9B�
"웩Bʳ�(�;�˅��:�H6�q��	9v;��LPm�S;�9��;8'�����ú�eF�n�F��[,��(!v�j���/t��g�e�OF�Fк�܊j;�U�R=4�[$�S��$���;љQM.�.!{��2�f�޸,�b���v�e�;\�V��m�E�����84�c�����O3��d�n�!�d�A'z.L�UZ�@��j�E�%�g�tz툪��6��S*�6�.8�.�[^�K��K/����g6WmRN����#�#2�W\M,8ͻ9�^s���ƶ�����,݂򽊷G�s�4z����pX�0�wL�38�-�q]�F�H�,���^�7�Ia��r��`��AeZ�
�j�i|Z�����з'�����u��s��ڰPJ�W���j߰\�A����7���5��X��u��]�w1���͛�#��u���H�8��/&���n�c����\�X^M;u�V��2�v��h�6�͉cG�Du��;79����+�)�<*5�ܳF�{n�+�NR+����T���a^p$��bbT�9�=�_���Rt4�y
�UH!"�w`�PRI�N߭!I���u���Ѓõ[TȚ�آluEN�%q�hIj��~Ԫ<�%`��:�	�B�+������E[ˆ��0XOY(:гt=��;���\�bʜ��*QV��QdCN9/��_ט�	ˀ����|���;gt|ۓ��flY��_mܽ��֩M���7��jS9:�D�NeȆ���V�K%ڷӯ��Q{�׻yz%������c|�֜�ꀫm�3�s�@�q�n�9$X����{[C$S)-�{.�i=8�{1!��&���	9��_N�3�J�Ll_W�I��9q kN*�S��������}��8B[��gb���#j�U�ۛ�>.Uu<t֌�n���%@j6�p���5�l�scY�_Bn���i>�b	�S��A8����:�����9�����k��ηY��.��{R���M'^c$��$�R�vfKY~��[ق@�X�v��&��#,k"]����N�,�{�gC��6��d���t���Nq):7U�w_VW��,u7 � �m�L��m�X� � v���z� ���]<u�lK��Q;,^�g]:�u������)"55���4�.��E؉dRV�J��j�]Mޞ}������]�<�7r�����'a烧3o�e4�4+z���u�hw-�ӳ&�r�)v6Y&�$�b	��)Ⱦi��ܜ��9��$|-�}j�J�dm9���I �䰤K*
`̶�jAnY��� �i�A��]**U:���<X.�APB:(8�4b��T4��H(�l!M���J�*GR�-�S�5���������^o[1�݃ȧT�d�ĵ�<��(.�������ǧï��ӯn:뮺믗]u㮺�OOOOo����6�6yˋ�~�NqM��y</~�$��UM���͵̜�Ox��}��o���u�]u�ˮ���]uק���������坿z�w}�¸P���<�ğR����BA8�e@�u�(3����Ξr�)��w���*�Y����i�{��#��O��
��ݗp�����|���p�|���jwT�S\B�N�M��^vU�v�w^�A�Ӷ<�O��C���8�\�������2������}bz��΁�eQC)�k�z8=w/!��Θ��%�����gM���H$�G�^j�w�Uy;s��<�)��_�W��J��9�|�z<����� ���wc�4H>;<�UPm�ﴫý�Lܫ�,K���X�5��,S�X��ک�:9}r�c���g&�`�k�:Ğ�M3mj��
*�L�4��e�ZrRR��! (B?�!�ُ���}Uu�3�_�j`� ��X��#Q;����E�wʤ/���6zE�b������ŏ��x�$�{Q~=�_u�=덥���K�c�IuRcK>��}8Bj�y\N��{�\]�4�/};�LŦ�0[���8�U2�Sb獆���Fqf�Fա_N�::���/�����\�� ��9^��*x�9�>��h�wch�d)��wy�]t�p�S��jMڐ2o�z\x���qJ��P6bY�Z�ʝ��Z�_\Đ�F���~+t�eh�`q�jYy���;:i�nư�q���}V�EڴY�f�Fg��Xjߣ]#6�{1}|�U�xHnWV����ƪ;�#1��iX����C�ƽe��3}JiM�sC��{;�����ᙠ<d?ag��d�Y+�R9���5��d����H�g��Wl�����5��v�@��]�y������,���,��wۗnmz	�������lN�M<�G:��ۆ�آ���8�/D�2`{�&�Z,f�3����L��w%��X�0�����Q��_�|�ZM�������U���/";��<�}��pcI���t����0gQ�ۢv��Qp�(Q�5�?f�����=ZX��Ǝ���)1��^�kk�[��dMsy�s�jc�P� �j}����g���n�<,���=�5���Yimn �57����kҁ��ބ5�i��jwo*}عY:��׃Zn�]Wo>v�CcZӠG�U���}ۋF�o��ë�R_r���z$=��鬝Hb�y�L�^/8��M�\�sz��F�0_��\�v��R��Y��f��wX�$�>���ޞ���޷�~�^�J�p}�8�5�Y	7kʏ���w-]�.����X��X��X�v�-�<�c!�M�>i*��wֽ<�F��zO�ND���'3�����oʄ�/�w�
�����^��V��a�&�ʫ��ANy߻{>7�)�=#^��㕖b�y�{w�P��vw�P��s�ӱߙ�c{���K���3�/wn;�W#�1W���EAuӖ�R��Uϫ��zس�9�Q2��˫>�t�5�h�Y�k��-�Hf��*����^���
�zv7�j��]-u���3���I�֕��S�e]�N��i/�LbI��j��%��ٚk�bH�C��!B� suXo�t�p���ZmiJ�q�=W�[-w�mƭ�ܛ�[���h�Ί�-G{��s�Qrm�*Y9$ՠ(�ȿPleR��S�9�1��Y�kK�n*��?�r���>��W%�����/szu��[5S�����;�|�Ǐ;n�����?��q}�J�m;��+]�܅:j��y㙙����g]�m0N+&<�W|/�������S+zo�y�T�8p��~6s��o\͵7>���+8��ې�B�(Ƿ����@���xw�<��͗�I�=6��
%d�:}XՔ57@�0Zޠǋ�.����tU�oGguUv�TR�1=h`�{�������2Ȟ�֔v��lR��^�����B�y��wt<�t�}Y�}��g./;vP��?�׼����a��w���:R��a��+,�W^��4z��f�\�)M�g���#�)�M�٩l�^�����;�_���4�I.���V���y���������k7T��e�,ןd }�$�M����s���'>tdu� ����w�]T��Xc�]EUw���*:�Y��w�}0"�!�2��B���!=�m�}><L���@����hϡO����cOh�m(eS�����4�d����ر���z
�<W*�=5w�/��7�w�y��/5�n�ik���]ŋ0Dyb��2� �y�A��a߶\��8����j�иm��U{bFXgz�`�Kv��^W�ht�)�V��)������z�[x�qE��=1[�9�t���ʯ[h�"�����)+���f+Vdo�X˵`��[��mܭ������#C&�]T�#��ᲫPW�%[�9n���D�y;���.�G���p�K�ߧ��z)i�=���]��7S�fP'�|���'sF�+����t��V�fD��؜�Z�[\;ա�,�6p,�68<�M������wg����u߲���Hv6T%>>��@�!�뭜0q��sڎ��P�f��qvej��Y�7$�vϰ��c��.���S���}9*�@�i�����ڪ�n�4;$�5O%� �,ƅ�]_^�7M��}Z:��4�F`W�7���n��o[�|k'���I�������'r��1ٽѾ;�{�E��])==���>�%�S��{�R���9�T��SV����0?���Y�k��>"D��T��B����^�{��;���kZ#�D�kO�}�����BA$����2+uu�In��Ɯ��a�+פl�̲��B�e]ýǷUs��3�VP��T[۴N�5d�}��u��H��j1m��.��-q\��4>n�wJ��1ݖy���8�F=l�҉�.Kv��;ܢ!���Y&��l��r5����{M���wx̟b��Y��{}����E����F�8+)�Wmzѣ���/x�VrΜ�V�ǭ��ƺ[���mM��^=
��&�0&^$�]{���+���	�s.�Ӟ�k8�m��)}�jmR4Y�`��hο�%�׏�ߒwJ�~�{������ޤ��+��^ԛR4^3x}�{("`���D�}�f���|�L�2/�x��&=�Sx�M!M���O��h�Y��s��N�d5T5���E`�7��F����2�}SK�l`l�`�מ^�v<����E�`!��^��T0A�i���7y#��DNc�� z��,[u�:_�gQ6Fz�Ï�3ע���SVc�f���m�[s*nB��iYJ�9�d~�o�r�7��u����3/4�6����^�6��5z<Å�B���};]4�����>�x{����l� ���)+v��s
���ܔ՚�G^��?�"�N*W|���Vƅ�+d��oϛ-��5�uvc��k������ ���S{xR9��'jEw�]d�{�{�x0�:����|���&+�E�S�G��q>e�s;��B<>�mSҟ�e��;;�����d�H�G=0�����#:��K�Y+s�!m�E7t��K����-|�{�����B]?��z:�љ�\j����H��lL�@v.��?[N[�U�	`�Zh琿��7��y���L��R"��`E_jpϷ"�t��L����W��A�f�x|����?����T��ꂪ̖v����Kp tڕ��7.^����9H~�rlL6�+��p�ڙ�E4&:j��p�]�,��gfc�q���l`�fX�h��k�/�xU�=�_���g6#O3l��4��7-�BSݪ��[W�c��lN ���F5׫��=Q��l�]W>�
�f}r�b_gh���N��	C�=���-GK.*co��5�E�����j��״�d|�G+&���z�������oR�D�e�ۯ��E����_-�ӹ27�,G*MƝ^�[���)�ok3w��W�<��p�O�l������8�/����ߢr�v�˺;(⭶>tU�H���IQ�|�H�\_���QS��y_>�������fj{p�j�X�v��=�w�l�wnT}Q�r��U׍car�t=޲Ɵ���酾���G�ùP6�
��@�9@q�� �˱k��Ľ8<�o�+8�i�;&N�8�x�{_Wtpo*�Rz''EA2&]���*���Q�k�dm�S[a��-9�u�άȳ�+7��
1��M�aY���o���霱�bU5Wo����6�����c�`�62qh�\4�?��+K�!�Ԗ���ic�n��v�'{�l��e��U�o��!�"�J�ԥ�i�<�v�l�i�_kE�;��6�����ڱ�1oT�q^|o����vs�c>TT�e���e�EL����z��Z��3Y�x�l���+�<�N�}�⌿b��5���*�^_�wN�XX�V����=�Y���#�S�Nv+B��r�w�������!�<����q?z�(���*B���8�Q�Ç
�s4-���W���Ar%n8���ooh�a�}]�|O���y��F�C�l�x�<���f냷�;x�z�D��H��^�v��-=�V~��=סguP�Bc^��z��l*���u��m k`���������`��7�J}��ôF�.Ԉ+�a�J�-�a���x�.�X����=;[7���[�}����b.<�g�G��x���;�y��a����O�X̊�sB�P�w�z/�P0+��w�۹u�T\�S�P���r4����<P*٣�iԎ��F5�!��Uu�.����������hqG�=�A�x��*w����-v�It+dKK�P��ۼ��v�f�I���ӎJ�+����
+d��@����w���^�P���mr���מ>��,�]}W�5�N�;Bԝ�Q�s@��*��1
�jow�v⋩�5ia`C;{&ѸA�ןO����|v��/����"B���Tm���c�+�!�q���N�'*L�M�X����'\[۫WG�t�7dԷ��r��N���\��5bpKS(XV�ޞ����
ᘦ��Ģ�dh����J��T)שR���˔�Ӑ��UJ�����B(P�Ua/s��k�]�/� QMI�_Ȟ?}'��WaʁM�?��{�d.y�BYE.���t<Q��r�77�O��H���O_����*�a�^eפ8�"1d�CVMn��9z��6��6*��j�;�OO`p�X�7��oa���{�O۽�0���s���jI��Gl��ր�k*�o���5��!s��r�^�m�6��DAV���	%���X՛���۾�h2󏏭�����2B6�}��w�]x�v̵.����egwO�k��:����]m�t��nøЅ�k%W�O�br��k�v�S�n�0�՘�;}{�k/�O[f�Y�h�xa8U���ű��d��λ�9�S �KO�x�'� U]�ç׸��J���E��pȻ��{= ��k3E��wB����
�'����l@�����H�mR6,�*7]<����of�-�ռ�d�?z�����^����V��n�yWّSQ���j��/MVc�~*��	�:Pq���/��VN�������u6��(��]gUw7�o_�E�rI�јq,�!�t����34IEWz6>��8p����۾S��Us�#�m���Ȅ�B��@e��|w�o�;�\��掕}z�{�,���,ߥ�*��:��֋�ԁ�*sU�`�N����%�K�X-��k&�.r�flGLL�P/As@��c��+:�ڝ��������8o*��7~���@j�Q��i��C�u����T�cv����	���c��vGVGq��c(m�C���~$Dg�j�r�j�f�P����5|	�ܿa�͜�%WO+��c-�{�X}�boʸT���@ւ�6�fw����fx�`��n&Z{F�г;��)�+�W�C2*�	��B�����V�ۆ��Z3��P�r�c*=��jG#�����W�f]�\�Ә�춷�({��)�:z3ʼ뒮)��J�bV���<�5� ���%���P�7*̲|���� N�2oz2��h;;n�Y���ǵ�4���=�����V̧cU�iɚ�J���ے<7OMŽ|�-@mn�5%���(�1L]��Oj�K#!�4��%�J��X��[��E�V���,��j�]Xԩ�L��O��p��8]�]F]Y5���5��v�Ě�幯�q�F�k��Ȧ��Aƹ-�<N�	���HQ�R*�SY8p�:A��l���$�w�7	�}Z~on���� ��:Vu�	ښ�P�)od�s6��� ����b(y�4͢��n�d˶ϳ�gnə�S�x�f^�U�Hc��
]�b����Y�S�{5s�S���zsj�\���Ln�&�^���ˇk<�V
����Q9���:��ޣ��/^�LV�m���V��%ٖ�E՟t�H��v.�B,ײ3�]����,.2w5��r�mv�b[}��=����7[xn��k�zUɽ�H�tMhi�繑꠺�J��k�v;���������:��>��[ݳ�=��P�]���6y�n`��0���w���&���\����ewn�h��u"fC�K�B��5ؗK�SZ�Z��W5��e>�w]̢Kb�d:���s�'
8�w&�ΔJU�(��ϲ��/oK���:��ؘ�Q���gP�v���3i����M����C������k����uP��Yn�a�X�P�-
e�oP�C�'	4E$�4Ÿz���z)K�k�F�ݷ����)�ڬ� Ace��ڸ��?��-�t'�f�SVJi�Vsk%^Z����Rz�f�B�w'[��7�'w�`�F)�̗��;el3%�G.��)c[�-(ڒ��K,(���²ݑ)ndpӻ{��1�].e<!�I�%e�f�9�k���7��m�oQ��ó^a[5�5*L*U�N7�_RW�21�Iԍp���*]��U����G�.*�������M;�;�y���V��vN���[�)��R}b��b�{;��h�mp�Z��/�o��s��5��_f���2�S x��4��kq�����7ʔzv�e��%�(�u;I�O�f)�'ڦe�T�.����=}�����[���Ώ T�--h�� +u�a��묷Ke��K���εN�K�ȵ1W�T��l����z��"t	��7 �Sdx�d��{O ��Uk�����]/q<}WW�NCy��ŀ`yD���q��ն�3���0+YO�i$P9���s��%�q�z�gN�����`]�.�XW�涖�:�/�sq��&�`#����Ff���͡y;+�X�-D�NSs���.�7��M��Z�a����8l���,������R�����k���V��:N��{�8�L�wqZ���WڦCo��X��[kjn�8��]N�)wi+;����s�}',xl-b����ܧ�b]�]��-F9�#�\��e��#�Q�� �ms��Ǐ�ïn��{g]u�]u�룡�GGGGD�������nj6� �ZA1�A�=4���Ja�).De�p��
�ɖ�~�Ӕw�,I~kv����������{g]u�]u�Ӯ�뮺�����ӯ���w�J��Fd��E�fPV��U"dR�u�"e����H}x�*/�ÅC�8o���:!���n�w!<Ð��']O0�-�9TAx�q�Ĳ�z�;���h��@#$�^�XN�j�rs�\�=���Q�H>%��_���\�H'$)2I��{�ǕT^�F���AG�\��N�����\.zXOAe�ED�(̪�F���W��.\��E~2��߼}}�Q'B"��Qs�,��Q�J#�S��4M�
=Yr�rĹfG*� V/c]�19�
|ar��#P����q^�d,*�^����G	��(�<��p��"�
���	e����b��#z�bν�ͩ��ԧu����o�����WCc��3� ��T�y��8����x���r�m��d(�p�C��T��6������>M[�����3�����	R��u7=fMR�����M\�g���L��TO�����g�fw`�P��jK�����.z���5/��36I�����-���d
h����(�ʋ2*�ȁEY�v�`c���ݝ�mufC��l��#��Wë)o�{�ak6�`{�@0����Z�+�����u��(j��ϖ��:�X�P$��V�j���5j�BJbl�5��t���/Cr·˫����d4�hܬ�*-~�A�c�f�LwT�]��{���w7��K���iMw9[Ӛ!�Q[�^�S֪�14d=�x7*�=�H\MA!�m��ܡS�Gr�3Oj+��IK��r������ߢ7�@j��u^6�n~U�}�U�f8O��ޙ��mK�$�,�rr|�\yP2�%�
u�v�y�֌ا>��Nd�8*��fXŰ��(s6Vs�:)�o*�MN}�daa�ko���:���ꬴ�"ښ#
�
�����H˳+yQ�1��}[���a�C�M�o���e�P��&n�Ԓq�u3f��{g�n�՗�T�ؾ���p�G�(`K������M}1�C���1z�xg��^�G�3�ԕ-6�?�iNR�v�w���ܪ��wPq]O��]j�}��K��w��Ωh�~�R��OoM����,���n���B4��3��|��0�k�_8�造�|����A���z�[+Q�ʲ�N�~:}��Y�y��0Z����`�A��+�=���Kz�gw6�wU�|mT�r�X���6���q���|֖썕�7����P��i����sî|a�I:HM߯ >����gG(gj�ڿ8̍�5j��6,�9]xwm�^�`�p3�5a�y�/f�޵v#7|#��#�J	=&�[%~l���{��s�;�,�yn')���p���l�q���*h���N�Ϡ��^m]����T�/a����[ͣ��
�6��$����s����C&y*��b�s��]�� �Wb��WkO�.>�7CS�I� 3����J�E�.�4:�wc�j�{z�U�4$^P��6Omg_J�۩��ڨ`�u˩Wʊ�B+���*�0	s$�d!�'�ԃ�5�ׯ_�|�b���5��.*���Z����.� $�Ȕ�_�FC�p�C�*�༚;����9"Jg��H/�Nf^���c��X�S��6����k5",��0��v�v�C�;�W i� g�9o�U=^��Ң l�~��e������;�y/)�n����4��~���X.s+k�\���e������v���)����p���� ^���riI4�[ܟ�k^j�hk;���Q�YY�q�U�l���oO����
�F.���)�f��ى�}n혝�kɭ9XE��5ч[�R�aW.BٲW�|�#ވU<#�M�U�߈Q((�ħ�yc޸8�Q��6\��Grޠ�=�p��p�wm#5�~�&y����z�k��ͩr��rL������+i�[Ԝyp�̽��^�N"�LN/��߾��ξ��W��z��W��Q[RX՛�zjU�Ȩ�������=�9��|�%���<��3��j��tM��/�PuQr�9M:������gj����:g0��a�AL����BPܼ�o���������h�#��F�A$�C*�!�4!YϺ�|{����:/�y�f�tm̼��ꄆgMh�mmF��\��voi�g��4�U�EU��EÅ�=@9���*u��}����v$��y*�穛M{0���c��S�OQ�/��͆�|=96��{>.1hp���ɼdb�6��Ͱ�5,3Y;]yD��Ih��`a�<⽰ȼ\��.9(:��y�r�q��X��?��r�r@�&(�b�\�|��k/=�\���
�\�\�"v��}�Wp��r.{��� ���X4ٚ��1{K0���6��9y���X4���t�-�1�HT��?0<}�p�S��!��Y6�vOG2��mL����~�܅��~�͹���d�5'�N�ݻ���}9�ѡ��OU���٧�n=����W8�S~�|�q�S��=a�Ǧq�1ڀ8�hyŮ6�7ǯ.�̏md�=��]Q��Y�}���j�]��K�w��������SW��%��Č�E�ɺw�,����4x��O[��A��E:�ץ\��T�X�Û��z�b�Ce{����4u���Q���
�<qq�k΂jG�ѵ�w T4�Q���Oe��ڄ��X�;�������/����ʃS���K�@�
0� �-�>�������|�{��ݸc���`��)�m	3q�*�6��k�VNa/��$�ݗ ���&���kx�[An�Gt��R�x^d����F�|�l�PG��{���y�)����7R�~H��OS=2ыD�Ce�?mr����z����l�玿�K�����/�L���!��
̩ϥ�wb�6:����`�ֽ\z�yx-j����>G~�a_�7�����i��G^�\_U�Hr������Eu�����|���M��r�5.�]�����xC��I��`w��L��zL�0h�6��!��N0;qň�9hR�\�tEl��,+�Ψa�j����W#{�lr�:Clt?A�]Z� O�������u^��n�{)��u�ś��㏮��sx`�����z���r�����@�mr)�ˤA)�f�g8L⬯Ae�4��B�*kh���A:�
�is��[��v^��v��vr�e�+R��B��/T�U�*%](�4��8�	 *��(+�$靷���7�/��[�˦pxu�@��l.�Z�Փ�+�s��=G�C8P�D�[?|�HO�|.�f�/���Q�k��4�`=#1�3�TN�=Pݑc{�K$N��n�<t[������]��;� �l=��S繯�����R�=S������̘)���u�hv���+�6��\���(-�b�6�!֒׽��15Y���K���\I�z�tt%�'����j����UJ��6�9�3T����m��]5>t��_�d$vClrV�.�䯘��6��y�,���k'�P�뫩�>g�ɭQ}�\4�f78|�|��ѹ�u���v���{W$����E�u׳ѕ�߆�6�%oq�6���Xz�jj��=ƃ;A�2G�^<�r e�l	��t����۟;�(�,�����{��n��8n�An[Kz�ڛct8e��G5�&��,�_mn[5�$DaU2�g�:��Y[V�m���'`�Q}�����)?�QV-��LOؾ�i�����%���!��]_���|����!�MF�T[ެ�C�/Z�=4��C�AĤ!M�"�M:f��D=�&�y�xN�p���8�Nحa�r�:�u�>U<��v�d��{�^
̦q�F��|�����pcb�N�UW*i�E �$�%R�)0[�S����(`Ç
b�yD�G���;�.�4�C#��8��Z�|�mT��_t}�_(^}��8�o��j�B�umT�l�_�2U>���|q�4
��o0k񎗻��U��Xc�oP���Z6|V�K�h�g.�u]1Ȫ�1w3���b�4j�3��m���zā��}oNgYϊ�7ɇ��&���7��u�N?�k��a�{"��wJx+%[4r��*��{%���٠R�q�odg:ۈ<6+���J��ܱ�W�O.�
��3r�g�[�������稚��f�>�ʖ�UbOB�	Oz��vaf�����nm;�1�M�k�Fc�;�Ѷ���s�c�sS�~��_������gW�k;]�y�����&��;���G3 ��<U��c��-v�Epq
�pN�F���Lۛ�+�4�'���z����2�.��w�����A��h[�Q����ro_�Y�{>+���+�u��{�Z�B�_^��wV����#��l^f�����"�[57ޅV��N;O8G�S%R�d�.}�ΠR��"l.��ϥ�a��e�n�۝vY7�ޤ�,�u���{=�q������{3�㭵�>'8wĞc+u���#hĭ��6<%�*f�F�C�<3N�Dw)/���P�
��EyH�ް���>�]\���s��^N.�s7b9��>�Z������g"⊙��딵J�'.(�Ƭ�|�)5��wc�#��Y���(Eh�)T���*�T��5��,������j0�f������ԤO�d>�;�}9��]�zV>�n�wz���E�vk�Wc32*u����lg�ې:��1^q��O`�IH+v�L�h��ک��d���h�oW����3��&<^C���'̋�_G�����j�1�_dCm�e��U5s�};�a��q�ݖ�p|�D{�f���v1i�����.��3�{G���U����b��.�0�����^w99��3���C���IO�jKƤ�`f��iٛ�1�dgQ<�N	��5-�{p���Uv��5�7ss���*���gGq\-ŷ4�xej8Ϲ�>t��,������~y�s�+���;#�`
��
��zdk*Ww^9RT�Y���΂��l��=�򠎪Ǔ;7J�P�(p��?{�j�JxK:���L��@�i��������Ԉ鉝�A��\������]��i�ٻ<:d���n��_,w+��|�aa��� ��F��	�ʜ��]W�>!�K���X	�
����ux����q���l�b��,��������%��qq轍�~7\RF����畷�������:�얋_��j��ˑ�.e-4n�oO}����>�ikJ����ݛ[��v�Q��s&�G[˶��;Z���#L.6.�^h�|��j�l7J�[��un�jb�P9�)뷟{Y�S�tNB�ս^�1�h��ұuWq焈��W�e۞v˒��^�Hg�,����<�Q��nzљ�7��;��:�X{��a�n�'!a'��o���o0Z]�;1ۜ�j�"���e��_?Cu�7ݯ(�P=��6h��8��|l��1s\]�&j��v��vlY:�T'qr�Ar���+�ڭ���ie4���&=�y��L|n(E�����ԁ��i"��oUlڪ; ��[��2���׷��޾���]ԕ$���i�8v�*g����N��_~���C�0�3[��}������3�"�X[����ӝƤ�|�3�h>�������ܝm�I%���;�ą.�b�_�b���=�[ۢ{V9\v�U�����~����k6Y{L�zXb(�/� iO8/½�KI��ռ�����t��`�4��=��#��5�WuCV�+�㊦�<4U���{k�:�����*fޗ7�͡�i���'i��2M.��&a��(���9�;�4ILvm47���eoNdT�e��ݷ.��6U�<����FX����� QV`s�����0�M,)Z�^؆{ckޥ^g��r�L�aӯ:YZ��s�3�"V�g�Җ�\����&4�V	ua�a=lM�J�u�Ҁf�56!�GrA�h�J�����x��n��Lb�m���;�}��7�;i��~���)���g��ށ�����sD_%�3L�d�$'�,�.����L�)q'n��5��Z���д��_d\�eK��;}����E�x�5i�����Ci�5�B�:�|MU����%Z�ژ붦�*����mG��n�#��3�A[{3q�AZw�%���=w��{B���ژ5��.:7�������CmZ�f�g�>�5��M����yHm��-W0��	m�I�}�m�c�h���ƚ�.��t����Jt-#�ޗNnǕ��7�x�(�f�k����
c8g-uj���vY�uA�yN3�Ku9�-��7*�$pFs���V��wR����]��Î�����iv�����i��̄����K�v�:l��.�ʛ��4Kf�y\���4�+�>���kw�k�N���Y�;U��낪�'��w+���ۣv���K�w]'\��x�&팦�����".Ng�l��B�h�yV�y�j���l�QR��r�Pƪ�r�e%]ڥ����oE���"�.6�oT>��U��՗�oP�����{;J��l�Q����v�e��1�ց�Ôz��}�к�f��9�fJ;�83�ع5�+���x�˒�lʎ�����sa4�c׻h�$1O���ըoϪ�sOf!`TЯ�:���Ѿc\A]��9L[�]x����+�� ��bj���SGR��l�h3���$�>#0UF盡�X.*�u�*veKZNeUv�mG����fAs?����THEbu̗��*��u�eɆ`�I��gV�Q���5����V�/�7�]]q�>e���-٠�Xv�Ǉ�+E<�0v�)��7sR�Żq��_C��p���m�6"ᙓu��Q��Ψ*��]Ŵ�T����6##i�8EԱB���]���L��e.Q�;�-�əf�����/x�_E���{���r��Z�2Ӗ�;tij�q��ÙӬ��p�����9�R��+][;N�����=�o$ar���s��� �"b�͵z{e�����:�6�n�:x�gNWG9��M��UԔ�����}cU��fݻ`�듼��|ի62�&����&�YW8T��w�;s��ĸ���E|�%r����JT�j��W3w;t��]�Eq��T�a,ÇWYF뫍�J��q�����]c��-7@1S��8�weˆQ�d]^���Wӛ��+w|t�ގy}o�q�ok��vm_C�$���U����Z���Yo�M����ɽt]��U��
�]�|ŋt��3V��ݮs��4=ˮ}YP:��b(�ui;Vvr$����5wl_h�I*�%�ȝw�;k#j�1�g˥*�^�T���g9����rҝ�3G!4J+V���O��O)��q����U�oi�V��HF�t�یw�/�Y޳̩��q���b:�S��R�l�{���f��ٻ��׷�D����T%���æ�3"QJ[EL9ne����a�!9P\9�]
��Z��D�:��M�@`D�&��h�Ei�k-KFb�*�&��m��P-4	�4�HL�����wr���;x��]��x|���������'R3���YG���2�QT�e�Q�Uq+
44�r��<}�_/n�/ó��뮺���\u����11111�c,�!q � �KJ�"�H_>=}�8zR�\_.���E�$��O�������}>��ݝu�]u�]}�κ��ooooo��?/�NQE_��TTQ�PSD%BOtC*.TEpΝցQ����"kR�,���"
.W
r}�r(��k4L�E�C̪R��D���F�˓�/�^�Q%)*�Q��;�U��[�r�B�0�A+��9׻Y�J�! �Q}h�$}� ��(�q�{�O$��QDz.��ʂe
��B�D�TG;��3iTG,�VU�e\�3�ϒ��*���Z�W*��('�.�r"��#�D�U�$���云r�Ũ�:#���PE���G�ªE/�!�9�gu��Z���-D�A8���C�	U�A6B}�Î��5}��Bt��@���󊈯=�
���'��ʈ��H>�,�K� ���\3���-��n붮�x�R������m���|r5]��T��O:�/Q��s���#�˚"j��V96_��j�A�&�l��@�`��2(�1���Oe��TRFm�O������{�{8
�_='���T.r;=���ԉt��z��Ge�ܨ�=�
���S׭r��8�~�3��:�������}�I��iɃN��-��3(	����͝�aPK�e��<��㻡�:Ü��^�����t6�;�o���یJ��x�}�^��Dߜ;�t�Zx�of>y�?��W��$�KnTÒ؍�����}��"N�sc��ս[ɯ�f���d��v��K���Ff�=o�6n�*z;'�j����fj�×�x��(H��p�m���2��4U��=5<��r��T���<A�^�ϸ4�9W_��}��}!<a"/�������ؒ-���O����0w{|�
붴�ڈR7�©���/�p�ԩb�������x�󖺺��)B:�}�t��3��VGZ���l�Īe#������B��C7v4��;ln��L�Ӊ�]w��ǭ��,��G�u���4��)W��%֗�M�U�!��W[ Ш:�^���4�{C#%1ص̅BRI[�B�9�.�kM��Ҽv6���:�a�Jwg
"D�&��S���}Pc�]�{���jߜ��2���	�h1/hq�al�rKm�w���]y����n���ͻǫX']M�7��H�͑NjF��2M<�uD̨�������*��9�@��3)�3t'ַp��.����	�vn�͢�r�㦎VMK�`̃�8ףT\�\\u��SȪ��Z�v�螇��*�(;�$&L���y,�+�:�gS��ʉ*���C����n������*�o<��yG��7��sj�H��h����{�ҳ7���n�ǩoy�����W�
�Q�z�N��O��$�<_�>�����.g!xγ�����������2��{�^)��zf�v��<�+�-Zck����nu��@�Y;����C�Fc�(�Dt8zʞ���99k��;;&�,Ů2Y�u?=i�G{8�f;�4&Vl7n60[�4\��{m���F��]����vdZ�f�8,��Z�:u<|�Щup�����eoe��Rq�����lf����9u:��{�-�q���4�"�;�]��*���a�yh�q��%� �MQ��t�7��y���֗ �ߣ�1�9��>)u�(����4�v���v̘/!�tYw�R��}��]�?\�MK�̽s깥
W�Y��5�=����pr�I���Z�u��I~�]���=<����7��d���w_��j�!*-��K팖Lcp�{Z%�����`�iLMu�nYg���<�ʷ;�&�KM�,r6�`0�f�Q���w&����.��#��^}��]	P��2:�fiڲ��'�o-�銿a�U����T9G�c��N�r��ܘ�٫�u��k1�^�Nل��/'�U����u��u�ٝVٝ��vE�1��ݖԐHG�]0��n��K,��D�U��wV�մ�
���X��e�Q��w���+����[߆� n���ʼzV��%�xb<LR��L�n�P�=�wPFT�j�q��9�+�yH�/��Kum����#�9�bons��a�\�r���]������[wtU\�|2�鉡H���#	�%[�'mK�Ya�?�:7F ��az���V����@��,{ˌ�;�����2L�����r���y��i���R5�ld��nUo����
(����>���fm�$������^&��
G$F����vt�C�v��J)�Tnn��_z��\�.�[{���b,��w+�^��L���_�g\�4'��"{��\��X}GL���ZӶ8f�~����ic�����H�ao���q͘1��)Y'���Lwgq�>���8�=0��������3�;:���R +�= :�k�k�N+���r���Y5V*�аv+N�[��N)�n��`@6dE�����/V�����k\=�[������N�gp�@�k��+@���f)t�+/A��{//a�^��H��,t��a��S5���i�Qan�aރ놮�K���o۶���
�ܠ���m~�:�+[���ut���O�ןM����g����ʠ=r\2��f�����Ռ93Hm(�g���l}x�EM:�f/H�z�}�6wKTq�g`�ȸfv�6!)j�*���I^��`�	s&eGz9o'0L}�Q3a_��ׇ�,��z��N�g�}G;�����Ha:U�e!�6e��)�t6��
�WY}�vo&ͮ^����/t7�a��oC�-lt@�Ŗ�0��e�X�
��IR���B�j hQn�:��uT���S���dFQS����d�zH#�(?���ݕ}	�H�@�uy���
��]��,w^����/Y9�zu�fq���X�Um��X[X?җZR��NT4K]��ʇ}�7�zzf�i����ֈ��j�3�F�$vi�y)F�p5�6>�γ��,�wVt�ϫ�'��'��]AW��/}�FO3����m� �M�m����,kݥ�~~�����JY�!�ղ���2��9b.ȫa���f�׎����=AyM�'�W (2>�q�y�gP#��j����K�{dsQ{���j�?�h����苁L����P�匕4V�M~�A�mJ�	��E�R��MT`-�ݍ��L�=����>ی�\Zc����V�c���ۇ"�lF�D@�ᧅ�r�	09�f���ԧ����7t������*��l�|ױ��ͦf�C���ݑ��e3���nEٵ�*����yS�n�?^$ŕ��9y�����u��`���}��/�^�?d��]Vӣd�m�*n�����=ә�JJ�J����ӆau@��-��E�W����ʗm�U�ԇ=�ڦZ�؜c��0�巶6O[��_[�I=�b�|�1����4@��W7�9з��˕'n�Zsz��r��^2Y���r�>�����6|��3����̷FN�9��!�(׭l]��P5�o�S5��X���c��yh�̫�&[zZWzО$��XS{Zn�,�y�<��>���hvc*���f���aԩ��Ce�kd������6����u:��a%SX�0��������[�j��ľǳw�.�܍LzC]�j�g��5�1���Xf���ጌ�`����)�vp��;7�V�;׫=M��ʢ��U��b�M\�*sy�-�3W�#u#;�w�����L�,��u��en���n�ꖷuY�i(�ZV�����xE�@�F�d=pz��6�F�[�f�U��飜b�$�n���k�]���\����.����פ�K]r݈���Ⓑ W�R#(-1wgi�ӻ�S�E�mw`����N:��=h��5��^U�ni�Ht�����4��&��^��ܞ��YI��H@zA�e�'$�^��X�ݪ��wqo>�e&PH���:<� Ah�zVQ�m�G�ۦ|�&��Q!�t/W�y���3�g����}繹nQκD H��J*�{���R���$6�<�۬��g����k[;0�-����^�x���zK�kR�c{`��}k����+w�"��<��=�D�8p�2͡ط���j��B�bm��x�|�]ב��pߺ�yR{P����[�t�y��8�i-l@�R�Kc\̳;�u��ݓ���$�)�	L�۾>���t������D��9?\��2o��k�r�����=BR1���\��8I�R�>����`��1H�i�~i�����m<_��37H����q
x���/V�8k��K2�{Z�;j��/��9�2�4:Y����U�b�c�y��p�ww������0��Q�ޜ����ʟ<Ƴ�5�����[��U��|�γ�"�����v��]��7龃��b�x-��K��������G&���ۚA���"�F3��u�.�V]x7ˡ�=�T�m��Hn���Qun�͡J����
�*<K�Mf�&�ᾗ9�9�D6��5s�(��󵻽)V��t��g��a:LҚB�[��`}oe�+@j�G� �0c�'o������5��5d�㏸���7PYxT�ѷZ�y��fL�g�4F;F�y��c�w��{O�ҙ�WB���{�Ւ��0nd��dR��r���،SBoʉ��u0%�34:�J�n��1��!�G�v�lr�ҷlQM��6KF��ۭ��0k��)����[9�ݙN*h��]�n��B$nF�N�md��ڞ�~g����$��� �;nM?8�X����u�TQ�}֜���}�	 �3D>f���>wTV��K�B�����(�k�"
=6���'.3l?\\a����|�%S=܍�s)/$akV�y��>�o7O��ª��7[-U�m֫*Hxl-�m���%Y3�"�/Q9�T��B�ʹ����걯9\60.�ù_�N��0g��%��:8��lG`�P��M	���ל����7�?b����,� �{r��.��=&�/V2.��7�?{r,S�R4oԧb8s����M���ȥv�Gw@��r��!�5È���;�Q��I�����u0��A�/9Bj�VK�	c�E��L��Ϛy�ݚ�γ�X��]��Z%�tU��������^o��ʣ�h<P�XvJfe�v�K�ԣD�0��Y2�KI�*)P.�~���0c�k6~��[��o�Tߴ~���^�})EGe^,ɋ*l_E�H�B��oU�m��OF�5���2��ƝH�;8�����{�:�������x<5�sW�/<Gq˞5hS�.0�[��6�>�l22 e4���M�OX �Vv[U9���A<�JA�����;�g�8+଼\�ovWgSG �T�&��@ U��^ f�,�.->�yY�+�t\$n[�#1܌`5T2��?u�J+7 ͎:-��*Rٱ���˦�#r�n��Κ#��>�b�;�3P�s.V͟}-k��P^w��7F������y�����[����oNd�5"�AS��<����[�'=�˸�Wl��ͻ[��e�B{�'óݛA�mP'w���%�ǫd5�Q�2��:'����b���#�9�9!d�������2IY�x3��XbN����9q��tU�7jS��&����X�κ��D�Ǔ��{�s�����'m�)�41��[��a�WӞ���u�C�s랻zӓ��7}�%��kC�[��mɖ4`8e�Uo#�[����&FD�^�0�y��@�J�k���D9P��c=5j���	n�c�[M�8�r{���&�3�����<5,'R�3M��V��Q�j$f3*�w��O�{�M��>0+����HI@�o=+H!��2�
�S5sMF�f��*�����!u��{��q���dݥ}�����"ڠ�;�nY��=˭H��3���������z$=]��L��:���g��d���ګ�}O��p��\2X뵝D)Oz'�j��S���$���f��Ϡ�;����U�ލ$)�$l�ʝdI��Ŗ3ov]��&-�Tޘ������'8�Z^�����ck�b��yض��>���H���aZ�fe��NT�J��xq�L��4ԭ'b�rߛ�r�Qr;��)��mLݱ��?L�w����_�>�uKk���R��e3�0�Op��rG4�i
����Zͷ�{ʙ1Q�o��^ҋ����xqF�g��s}P������pUo!��Fd�l*E.�䲐���%�Y�zؔb��4�nU���������E�+���ᾏ��=޽�:�ոb��o�%�s����'���J79p����t929eWk��Xɧ�+�{j[AG��e�l넁�yU�����E���N�������}�,���sP�;��2�T��ʽÆٜ��I�
�C�K�B����ML��:塻f�ⲫT���ݝ���q�d��N�Y0bw�p��o�?���(,cqU����J�i�P�p�sB����6�b_f���v�w�/�Z�Vf����h+������s�D�v K���h��n[[S�}8݅T�
���;*q�ȑq�ҩy;]���q���\���j�'��K]���	���'3-��Miث:����hw�Sp�=����k��D�Ga�6�˵]nu�0�sq]�wJJࢗ6ګ�ʾ�����lmr�I}:J���C��0�fj�\�>���l���h"'l
�p�x�.I�;u8I�|���aɳ
���Mk�WHP�WP�0�Pڮ��Wl�'j���A{2:*��K�aL���o��R�~ˣt�x:�^��=Նr�PTb�	uQ�i�g��UN[��L1��hS�����ɝ!�K��Y*d�E�L�[O����^$��[D`�5�U��7��lͻ�5��қ�R'F��~vk�{���oF���(��WZ��R����fIبK�ӯuf�v�8�;�G'�y��`��yJژ��z�-�����	d]�!᦯�
���`ۇ�iy3)�N�l���;ˮ%�ڜ�8�t.���Oӽ����x�Hvf� ���_�M[��T�}�.E[�:]I}7�����'-$�k���Њ���u�gLY����:kHX�M�>f������N�"�s�\ui�z���UO�huc�ŵ-�g��*�i��R͔�PҪU^1����]���IC]�١鵼pm�_j_vE�7D��l�t��ҳ�s:���3�۾��]*�.�¹V�O�;�RF��3N��B�̾F�dt���8�34��hk�)�V�:D���º�4�rRq7vz��7�P�k���c�Jֺ�v+$e���LpR�w
�^��!`X�H3��y`�ه]䮾��_G�f��wbR���°m9��{���?e������w@�#l��;b��_ޝL�OuSo���m;��u!� �0`O�[Q����s���u�z�!����/g��(�ܒ���{]��*V��UЫ��f�ٷܸ>���s��r�ϻ��L��l]J#��kI3��~^�z��NEZ#����ҋ��EDQQ�Z�8ͷ�qǏ�ۮ����뮺뮺���u�]u���������.V�6Y�*z�;@��p�n����,�DN�"�ȉ�Owj�6�o9q��������}���κ뮺뮺�뮺�����ӯ���^���Mk�e�n�Q=��O'dUn����V��y�|}�R�iD}^�Ez%4˨V�QT�4*������.~!
��8Z%z��Ңt(��r����4�>�eˑU���¾R�`H!D��5$��ZbDY�TQ�*��R�{�ER�A���q�oW$����閵6r�J�p�0P �aT�DWtS*��$�Y�FVJ԰Y�]�I�8��|��ʹBa��򯈊>�"(��A��'eT\9��(��J8��
B�f���QQʦU�D��e�u��!+Ԣ�*T���
s3�����+�+6�ӝP��*.Z�����ZS�*���1��!F9�F�fUuB�"�s�EF�f`��#�JNN�k���5:T��{	2��Ds�/^v��C�k���&��9z��u]�U&����R�-G����y��p&da������}��XkoI���8AU�˰V�
��n���5��� (���Q���u�6�AT��s�AYeo�ux�e[��>I�����ơ�&ᐦ���z����rܓ�]!��vL�zl<��Y�a��j*�C<ϳ�Gr�{��;6*�lqK���*��y�&���E��Ҭ�ڗ�cmd�n�u�e㮽��N/�d(Z��^�9��ȸ��%3]���i<Se��8�7�3��o/4�6�e�*5d�q��8cz�{ ��n���(��3q�Փcl�I��i�Y�䳯ݖ�AƬ�f��G�_�~��1Z����!�`Æ�:�wXoY�<��ñ*t�n�Ya{��mr�3g���Ǚ5Ssd�wNI����fq�ix�i��v�C��s$GV�;��?^�-y�q�a*&遊
&���nKx��ʹ��s��~�nn��*�4�Sǖ��\NdZ�%cg&�+Eu t����Սb���j7,7�Mغ��n���ݟJ���t�u�L���n�AYM+�K��Dn���%e�~\L	����ub�3��5�I?��>>Cߟ�Y�$f�×n���|�S[5�+8�g�s����ˢ���֦�|�[Tt�H�OP��}�jm���l�מ*��y�Q�{w7��C~͝��P�a�o�B��j�h��x0�d9�T�{4��'��LLmonF�v��%N�Ü�0k�3��*�n����UM˥a%E5M��sh�{xc�s"��]�\bW��a7��.��U͹�]���eNFs�>;���Ӯ�T�����K$��q�5�,%.[�U�)]��C����ޭZ�u��kı��C��є��CC�9W�zV�]�rs_-����dlİyZ�,�B7��vڙ������J�@�Jy��pc!K�ؔ��K�.�ꚺ��;����M��\���b��foP�F��T��a܈��ѝ�pI�0ĝU�F��V���b��)>��QEϚ�9���۹��#���uIeF�88���:B���h1)�ף�M�r�X�/�Ӗ��8G�b�<o䇭^9�i����N�%*�e5K�*������S:wnci�369�Wj���y2ڡ�Z5tT����E�YwG���a�%M�ڨ�R;<3r���"#��FL� ź�����[h~��P`�5C	�o�o���ìe�đfb�G,���ŝ�'yx�����)�Ɯ#��[��뫘�m�j��e�{9?�m��Be'���<�|�:��%�E�8�۲:��8�%V��3��=��R�R��g�z���ܖW@5�h�R�;�!V�v�����{�ސ��\8��-}AG�0���������z�5<�u��r�J��?�M����n�Ś�u��ǡa�,1�ع�5�cMf%��{5M}/=`��k�cN�ү={�����t���5�L"���O��/!�kjۈ�޺�'��R��������,]�����<��+.�&g����9�,/���@��"��ʇ������`"�;�;�~�4_�����h3$��!��3@��`ޖğ2 b��&��
��P�� {�a"�0Ҷq�k:������P"u���A�E�}W!Ta�k���x0�BH;ώ�I�:T�E�*r�:�i켿*�{iAτʖ͙:�xfe��һP-�^>r�fj�Gi,V乢�3z��8P���6es�\�.^�k!���=*�u;8vV�JŴ��^���O�1�����is24�$y����~o7�Y�n&�����ݭ3_aS���>�Є�t�{&/B������G0�'ra���Jܑϸ���rS�)^Ou�8`ح�x��lB�d��:���7�[[A��{&�/x- i�W�N�5����(���E�1aմ�uk��U2��˸��\��)�n����u��'�W/�t?fO�����, �vZ�z��;ͺ�'O�l����*`ޜ�V(�+7�ï�$����p��-,��77�;\rl���κ�R���S:}1��ڲ��z�$�wLϛ�V�iwq����:���Q̎"�������O�Mʀ�s�\�N�>�	~[Ow۝5��E�V��Mǻ�6�>�t���zDb2 ,%����(GL�����ݛoKk�)&�ɗ��t�a��&fL#���u�y0�7��T��lҏ�~��p���,��[?��h��i�u1�>��D�Q�X��̮n�%��K��0X��Q��|�Ljd_>���0�~�o[��k�����qn�m�F�`� r���>�[����X|�9]R._��#zh�; ���O��f�-�Ҿ��R��hR�t��+�D������ৗ�fw���]��]�<l���m��X�q}D)B�[6�.�����H���a�߈"�<`�5���5�7V��=�H,MQc$: |��ƞ�ه��e=���.��x7������~�N�Vh��ڛ�d��s��Kp�f3�Y[adR�}L���5i�M.Tl�޽+�7��_���LA�^s�i�7��fh��h���ߊ���Q�#�<��X{S����='�焟Fr�����	.� ��3M���Օ�g��&�$��v���d�t�vSyx�)���\��l/�F�ʽ��%u�L{k�	Ή��7��{Z�Bܽ��e�y4��g�ץ����S�xrZ�A��T+��&���:��w}آ_��950ncdr�/Y�ݫffd����Si8gu56J�o}���'�wx���������������{��7�����M�Ѫ4��} �]��쁁���螗�q*�9M�4�A|#1]�|���9���>f�=��A��}��M��K�]I�.�e
[+lT#�"0ۭ��#'r9�/�+\�#Tn.�����'(����v*�>�7�&�ᇃw/?��+(湓z{:�ύY"63ZQ�4���������o���"�+����
��R~P3��NP9ϲ�M��8f.P����|g\�yo}��_�3s�alCu�L}vV��m7#��?���������ǵ-��d���.�Ny0���9|hW84Ex��]x}6��g����9�Z/���f9m�t�����j9�=��~���x�ȩ*��ع]���\�=r����2$��b����Sjg��֕��U��3�e穞b�P�F,�;�o'tt��I�X��^�:����i�x�^�ix�#��V��Y�:W��/��LU��M�V�����>�����̽����ʷ��1�����,n��̥K/ �WU�8�SPhΞ�:X8G������9_��*�Ӓ�p%b���J��D�*��q�r�ϿJa�4��܃�e^H9���|�9���n���F�m�u��ń����NnF��ޑ�j���)j�h3�AZ#uXCɎƩ2mWuo	,Zy"81s;�;_aTe)~�{}�����'m��q7gfզ���{`��p<*wfr�r�E.)9$2�%�
i�QI�!ɄG��0c�6M/=���g��Y��I�1��)L�)����_㕳o�+�_��I���0E�?�����{Y�����Һ���A��zr|�r�k��[#����K=����e�,dma7բ����<��ߖ���[��_�l���X��������F��壼bz";4��iz�R�H.�[w�8C�X�Y۬Yc���µ;�3�������U�i5n�wn���[>v�����h�����Eda&���&F���&/�Z<N��g@����#��ޤdʖv��K����d��[����Y&�0��`6�=ra�4_##���kT���d���wӝ�}��4ľd�3��l2R�d��,�� ��N�%���*�9y��pka����3�P�ݐspr��h6���O�"�!i{ű4�������nټ1qd;u��ᮌ���qqp�zY�����>���WҺ��3s22o0#�hn�R�*�77�M0��Iqn֎���L[�н�Sr��TD�$���#�v��ə��]�Y=��2�`ݮx֨��c(9�2�R�D7���u8ܑ�B?#�;ܛY��7P�=��;����(0c�K��o������]^*����0�3�/�V�9���_pE��w�:�]�#A�m�@0�{�(��T�̈́'�)*�r���Vt�>vU�n�Q\u�϶[=��kTz�.Tް:ӫ�ndQ��L�/"G��7k����z�����w*�ٹ^���1�A��_J�S��J�:�vNV�oR���6Ոv��_��<}��Kz�W�L/oT�얟]��=� :ԅ�3�L�v��]�w����S��wZJ���y�]��C[�*5cD;�+�0�U�b�v;�I&�["g�u�6q�N�Ε���w��Ћ���n��-���Nsq=j�=��)�$�H�E����)gi��qU���&�f�wyʽ���M/�Q+�-�j�usw���(�Y�|�pK�O0��t[���]X������Z�G&���v�zMxLjU3�6g�]{y34���[��,]���L6i!dڏ_/Y���cwt*���e���o���.��[����Mene���e-(Э�>]3��T�,+ں�S�Rn�u�mpQ����A�����zB�o��\�<	��������]V��hsu^�~���mg���jqW�����v�DWz�߰o5)MKc7.�==U��nDp�臚�Y�-^	�vY����׽��k�½�����hiI��{�x����c�C��_c6}y�^�ʉ;9��1����"w��ki�j'���_3^[�y���^6���r��S��s�f��<8����+�L��扚��;cB%)�^�v��L=�뾨��ݕ}�[�^uAwn�9R�/mgN�1i�tf�� k�!�|��Uk���9GB�u�vGb�gOj`���m�5�1��V�-fC�ӕMqՓ��Wے�䭎ޫ6����^���N�Y3gq�F��22fCes�O����Օڈ��Qǐ����Y"��Bʭ��}l��50�Z�n�1��!X���]��ݥ��$^���T�``Ƙ�%cuw���&�P�[��U��D<��W�ͦ!Y~�D�E��Y��A����\�ʽ&�vl:	�[�;�}�.���U}���3��m3YV������\�]�扎�ޔ�y8.����	����X��v�naph�t�<����Z��k,28�]i��{<�oO5�#%?K��!��D��gj���+u,|i����<0e�T�̓��`څ�/|2�	l�f�6�/}�3{���t�:�ae2]}�u��{�&��0��ə�g9�w�QU�B4��1����@֙<k�Iw���2�L��Y`�C�}9~Y&{�{���W�5�`��D~P��v̕v���To*�cZ�ɓW�����;���>���.����d�u�t36�.
���-���Y�j\Dybˮ��e�;�� ��O{�E��3�	���s��Er�"�w�S�{wx��a;�~�dRIn�m5=��Xa|���8����l���f�q���Go��fy��;�:D������6kqS��0 n�u��9�d�ƹٮ�g�Ʈ|ܭ���d>�YwVn&�P������8�D�Ř�Gk��ot3X`M��-�����"�>�y������.q?x�����I'��������� ��D���r��r�3���ɤ-2)iZiV���Q�5`���M+CL`�i�M5U�����J��j�LiV�U�Ui�M1V��+i����������M�����Q�`�J�ҭ5U�0i���i�ZhiX4�Z`�J��V�4�V�4���iZ��CMUi�Zbi�����b�+#M0i��0i��Q�1V��+CMUi�L`�UZhi��*�CJ��F�4���L��*���d �|7ow�4� 82*�#L`����*��V��MF�4�Z`��4ʭ5+LV������i��0i�LU�5U�`�UZhi����5j�M4�J�V����4ԭ44��0i��M��i�����V�U��MUi�M*�UZVUi�MUi�MF�4������&����V�j4�Zj�M0i��UiZ�̅Z��_S�V��-MJ��L"�4%i����+M�!Zm5B�5(�
���Ȝ�ɫLR�6�J�5%Ze�B�6�i�1%i�M�2i��i�1R��妴����jjEi��
��i%i�i�J�i��M����i��jhUy���-6�-L���Zm2V�M%���4��)�j`�p50jb�L�5155U���150z�ʞ#SQ��SJ�0j`������S9S������5b�5hi�MU����������W�̪�m��֯�}�=��������쯫���<�����__�������\������_��������W��O�_�U(���d��֫���v��������~���UA�?ƿ?��ޞ6��������/��K��\�5���ܶ��r"�0�SB6���f�������Rֈ�j%i��"�(V�*+++�U�iUYV��%�UjYO޵H�V�U�jUY&��²UZ��Uh�VE�Uh�*��UiVR�IiUZ��Udd���*�SJ��ib�,�L���*��C���rܟ��j�H�I����*��U�Io�������~��ڻ���^����9���+�9_�������^�����W����?ؽ~��*�>������?_�}�*���UA�����_��ҥ�+��|֒���\~��_�����pA�����n����p�UPo�����O��ޒ���~��گ���
������_���^�/��]��I�UA�����iUA�U�w¼���?z��r�W�����/���w��qo��T�[i�����U���_�����_���������M\��Ǫ�Ds������������e5���W W�� ?�s2}p$e��ު�CT��+*�AF����� P� h�����R�-	� J ( �(�
)�SDl͵����M�����mQ�V�2*�j��-��4��m��B�����Vf�Ղ���im�j����F�#f(Sjk[m�6Vj�Qie��ٚ�ւo��ml���Y���4�2�D%�Z�kU��Mj�k5,�l�+)d��4�&¡�KkL�T�YTZڭM�Z�dfm�m�-���lYm�J�ۜƑf-m�x   A��b�it�3kj�4�'M'ZةQ��Ԩ�a�[KUZ�+��:��ʵ��[��ZXͷu�Z�Y�V��qw3kl�m�qi\���IM�kX�ͬ�ml[m��'�   Y�44(P�-�an{^�:(P���hP�B�
��������k��jkc*��������X�����K��۪�������jV�Ev5�l��ګm�h5%[�k�X���   ��k#6�m��nwSU�i��]�ZUi��a��[U�Uit���VQI��Ui��ӝmje �1ә�[h����գ*�ӛ�̪�CNkmcK-Z�mM�mem��   m@���h�)e�
Ut]]�U]tt��#j��إU(U3���
���T�J��$���̩���YZԫF٭�1�  vx�
Q�QJ�5F@	.۪UQ%k��vQm�WTj�*�ԁB��n�U([9����(Y��@R����5MP�6�b�V��  ��)�Ssu%u�F7f�B�@�Z��]��]j�j���U�aQ@�;��v�7i�Y)(�v��cl�T*�,h�ѩ�   ۯD: lu�  �� ��@��n  
�� LӜ�O�{�� @Nr� ��� h`t���ɳmU�2[%��em��-�   m� ���  3�  ���  �Ӏ  ƙ�(l  �+ [��4 :\�  9�@����hmLfUi6g�  ݼ  wm����� �s@ g�  g��۶k�  ���
 v�  ZV)� 3�5k-l��jV��5J�   !��4 m{ P۶q� X  �`�c�� Qj� �Æ�(ܸ  �cM�x&�)J@ �)႔�! A�������jz�4h)� ��   ���<��L�  �Q"b���C59�Ʒ��o��{��-d�V6!b�-P��ld<+�Ԇ
}kCҁ��P��W��}_o\����1�co[m��cc���co��1�m����1�v�m�����m�f�5�2�P�uSUP��5Hܩe/`:JYܳ��U.�Տ��0n�.�\�$�ޑư�4J�R�vPw�_VKʹ����;$m��:ܼ���G��K��{a'�z���V��ɤ�,f� X��J��S汥��mӼMj�[H����v�o`/%�� )P'r�������tp������}���l�>L�.��:�7*D�ki�u3[�)V���ZJL���#���3>*�ǧh�R��&��Gf��lՉd:�B�\�5F�8j�	E 1�ظ�#tBrK��"ӸfTQt*�X6.����0�ǘ7YM��J�91� �.	vb�,c�����*�n�^F�CY�wo�"q��πّ�_ۛ������n�sf\N��2D�!1��a駃m.{K-�.�ʟR=E�ͤК.��;2���t1*d@�i�G7�|iu��u��=��ۼ��ۣ��İ7hE���_"Q�J�n����8ڗL3{�5IOv�e1���[C�+L-\�᫲>lXo��1�5��[&�v �oV�x��t�:{�쵹Xpr`�(��Um�ј���
�Bip�Ye���Bݘ,F`M7XM�W�Qw>��4����$C�ɞ͓�~�ؑ0+m`7LY�X�@�5��VĞ޸�)�Te�Uk)r�mM�i�%I�Z��k2�ӱ��mm�c/n��xD����X�ndb��n���V0M�&Tas��˸vO��~pd����;�S�L9��T���fΜՁ]^\y��M����}΃�0���YP�"龜��ۼ�B�@�!�vX�a�i5��WE�j��i��mfP��Xʛ�J4��4��Y��W|��ֲ�C���V�<T(̫�v1f�/)f�Om2Y%$��h9�q���N[�z��ǹt)�[z�[h���b6�H��[�LrY�2Ń��v���**���t&#�Q,峠�ei����#��1�:�f�j�1V#E��ʵ� 2�;cS�F���+L���)>]W�M6�gܬX|>�F�e����){�y�x��>�e�cl3LLکDK.fd2����
�Ɇ��*��^:Ԏ]n�Q����ߛUg6��t�i !�3m���� �r�چ� ��܂%SqL��H���si�M�Y���N����`f[4��5��XAb�15��cN���]V��㨢�5X�~�����{�։Gq��,R���-ͻ�@Q�rb��IV�{��G?}ݛL��1ZZ���ff�S�i�,�,�D�s4N�6������3�n��0 8�N�ɽ[�����'q�L���"��ȭ9 =ܔ�5�A�]<�jAL�h�pbZ�Ŧ�V��$�x�p^�������ϝ��u N�_�Gn�m��M�,0&��UX������gsN��]0%�q-�I��{ Į��5�t��6���l:�u"�;���d����0�qLԠ �8����7�`P�Dk�0�&�x�!c�)���PƁefX�A�c7U���1�(�J'yo��/#x��1��K�(�b5��ؓTK,�ӎ�;��PTP<�j�uЫF�ȼj�5A��]��{�2��$7�V�@���3q)����E�j܇k,ܴ�@��T{�3N�;(��H�W��t.��Q^%pdHI��'4*ںY��L�S���(PD�b�@8��"!%fM�okNkq�k)�_��Z��[��]&�/�i�H|+�4,�����Z)��յ�R�SU�(ojݬ��r#J���7]�@3�V�[�#yD捭��݆�iP:������uc�JH����hӺ����<y1E��
 +��u	�n�N�f-�.��#!��9��ы����
�m����<1֊��W�5�I_Q����G����癋(�|SJ��z�q� ����k7�a�%�2���u��/^��G6�gV���k�t�z���i\fq����`J�B���x�J�
���H����7��`��񛺻RŭӨ��K�nͷ��ݣYOͲ^l��i�����������Z�/V��M�%�+�j�ސ���
C��x��֜u���'���`t������� V����Ŭ�vr ^*)ƣ���;vso7��n�:&R�p��N�"���Ǹ��4�ĞD��ff��׊h�Y�V�>Ƌ9��Fh����"��S�KU5�{E�2�z�Ou_�$Ƿ�Д�H�{ui6]?%���b\ơ](���԰L�,<�X�AM�MYC6��W�DacZ���Z6!y`��\�.[���%��Gsn�˻TԦ*�TX�ݡ�n,����;3$[�+�hZ
{�J�b��r=;�ҍH�(6�_h���vl��E�b�m��MQ�&��I�>N�^�nK�e�s�{ F�,�*h��F�6��E�u��u�x�yM�sFd�RV�,��D�-|��T��Ŋ��:KX`lk�I[-[�wc�t!wz�LÞ���0Bc�T���̠T	
qkJ!��M���:��n��v��&n�ݒ���ŷP�6�op\2" �!�x�0�ׂ�e�0�V�L�Y�-��r�N�#�f#�YY���AV"��[�� �If�8��f�n!z�t]�b�`�S�jF��Tu�вU��~5�S���ej�1TП�,#"�*үm�ӏ6���@ Sz���z��N�/sH[��y���v������
ݦ-��Z�6��Y�Z!	�,��5�PUn���3��"�*�͔8Ml�C,B����%.j��^��]��GHݑ{2�wF��{!�w�<�(lt�K�&L�9��sY�P�Fe��ֱb��PC�)0�IM�0�k[�8d�oZGi�F�Yw�F�A]jyO�rIk/Q{h���Y%sTs��V��6�ٝ��av��o�7�WIVе���i�i�զ9iCr��G��lg<��ػcUz���n]ԡ���;�M�c0�'6�[�HS������k.ff����:�n�J�dݢ������oPj�]�r�!��[n����>u�Ei��B��՚�N��d�J�$�ipi@9Z% j���@ˇ)mK�J2ރ�d���7l�u5y`�� �mk�Z�����4f�ykv��F�G�4s�Ƞy�!���
f�qʺT��+�W���nVRz�9��(�v�t�ϐQ�5�4INKÍ�"�6`i=z�M�,�XÌ1�nμ�`͆����f����b��zy�hw���LS4��Fn�B���vw�5�+K'���������,�g��°|��Ѳ+y�
ѻ�n�����^����3t�1;�u��`\v��Mnd)fF�^-z偦�)J�X0}!t)�mѫL$,�m�Z�ʒ�� Ɲa�j��9{��n�jX���DBu����PP�O1ȎG���[9��!��Rᦰoʭ�&��ǩq\�Z{���Iɥ0Le�vFD�� ��Zrڬ	#��r����b�`2���cv��ō�0B��`�,�2�nP�ĭ�j�Y�z.�\0$joUj���7��7_�@�+cj�j���ь���M:��j%`fZ�mm������:�|�ս��QF��mڱ"�q^�<���B"kUm5��JY��	7h��5l�ܛ4���0�Y��Xi*�"�`V���p���2�Yߌ�-m7v>�M�.�̨��rc����ZӋb��FL�!��ǽ4�x|�����X��S�Z/0�A+�i���I��yW5�"�����p�%n��hł���(<��k��%5�u5�=��u��5&���a���H�g]l�_\���0�̹�u�ŵ�Fƨ�J�E�3R��l�1IwR�:ʌ[�Jʫ�Z��(L��CN8N�f��|4�Q���d����p̂H򊬬���eCY[���Yq�W�\3%M�+~���w`DS:>G1e���4�\�Z��neK�f�C�1A�ʐZ)]�&��r�ق�`��L��(C�����\�еȧ����+�]C�I#�֡�Ջ���0�.���B�[�P[��.ʚ��,|Hf��U�����:� �씪]رt��w�C3&7E�yݙ�9��Y�>ť��n$çz�Khm�+.jl]n$'!��G2.����$Y����e�D*�T�Dϥc���'���bǪb����dnP��g��٢P�4%ތ��[{�;�\*j��	��ҝ4.�+|���\���xxA�;���y��a�����f��)Z������F���V��+sN^����A�!ɇu��F�I.���o:��y�ewP4����DBΌw�h5334=SY�r-+MƱ���2���Y��I��j��[ �N�b˴�fۢrf=��m7/Ry�Mj�������$յ�˧E��m`�A^৮�VRC�Ц�+����ݏ--�(�ȴ�Oj+�OX�e�Y�V<Ҷ[a<���l=mf�ݙr�����iTwMK�[Hr�������/(4��LR�ǻ��`,��$i�x,<�b��c���6(�h�Ei��Q�I��7Xi�tmhInL��]��Uo%�P�3	H�.�S�G6i56<�֫pۀ�h֬����nmآ�
e�8�iy�P��t�7	G[�gQ�j��̼osU��R�Me%j�4Tӊ��2���:�#ͅ���G�;�}�����ı�ct}�8_�K�5�S�`sD#b��>�h�̒�UF͍�H֗.�3Mk�&(Ӻ������xkQI�V����F=N�d��c�R�ޕ�t\�F��̭ҽAi:(�~�mME��JP0rsdǴ�j݄��˼l�xk ��0�Nn�w �z-�w�n@�&+uհ��V����:U���k"�0V���W�Vp^�yh��O��Xt�}ۥ;|Ckǖ�XF���,��m3h��f�l*����a�ݝe*�Ǣ�hb��Ȍ!�rf��KP@� �(���&p�gr��z���)�գ����E"Ʌ��B��bXl�V��t�	�ũ��3�i֫�d:�\�7���c#v��V�r�5Oq0�EO�I!�tJ���9x��-w�N�Dcf�ٹ���ͭW{���ʘ�W�
�Z��c�A	13v��ͺSSJ�7D�mef3����sMZ)K�J��&7	��)�1�M�u�m�N,,O���Z��cĪ�V�R6l;�S�"'.fEWx����ʻ�+5PS_){3k&9h�$��0m%w�h�Lb�U�T��*D9w�a߷*��7t��)RAl'1	ɔ��n�`�Be������Lw����qƍab����;�kr���g7M(�F�����k-��%��KF�34����^��9�ֵ`�\-jj����U}��WY�D*68����m^�"뚳� �Qx�3 ��8���"QB�
U{f�;-6jUټw�kn��Ji�Y�����!wHs�zwh��f�+ͪ¶�XH@*b��c�U2�~��}4��kC.�,�k�"�TyD�Hi���ɑ��Ӭ�f�l��Z�v���6�����b��ݱ��,��^SҀ7HC��Z.�5�)�E�M� ùWm��m:�g�m�pLC	��0ؠ��5,�T�x
z7*��I���X�mcoR��ݺ��iԇ�wrڡ�Qg4]���;����k^�F�0��Z�.�i1�j�8�ɨ�m�S�q��FT/Xԑ�W[$�'�:#�.T���f��\J={�{WU���gv��S��ʲ,��
�M`Ь� �I����6��:����%9�N�-fԱW�㑣�$�d��JQ�u�,��1�X�0ÛvU��^޵ ĕ�.���ehZ�;m�	���@챁ZʬWW��$��a1m��{��X�i��R+M��J���9�!�.�zA3idV�6��	!e����{�YCu�h]�ل�piʖrд�F�=��l#3-�8�.�(�hfj����� ��tB�OmP�7���(p�2�84��&9c���Yø���}T��U�m�)�U��;qu��m�� �3j�MV���־�`��3b�^��ݠS�Z(C[r`54%#�9v����v�n�Ơ�-��٧B�
��kg�Lx��4�M�T��bF�c$Bm���^0����q3��3kj�Է5���wg͏ �r����Rԟk�K]�p���M,��y,7N�ز��E���yF`�7�)ۦ"D��E&�TN�a�wT5)w��3��f�&Àޛr#F��zV^����DM<�f'�txF@`�&�e� �O����\��3}|�NۭGem[����P9ue^�R�C g�^�6�]fnm�A�i��(���Ƕ�4�!pQ��q:5	�K�ʶ��Xq*����/C��j��cZ�	��(��CJ6�h�� cʂ&~l}�o9ѷ�M]��IB�0co*�f��.�`���-Y���.��q҄QP7y{�(�V��c��G���I�Y��_Z���IxCA�F�l�v�m���1!Z,��$���[��7Y{��D��5�-F� Љ\���K=8���Znd}�qS�p�Z2n���7룒�ֱ�m��sP y5c�y0��;��(F�.>���ќ��r{"Ƙձf�~%d�0eh�QzN=m0�c��h%�(Q�f�'ח���ȅ���FQu�5m��#A�z�S6�akrt8� [x�*���Ե�U�<$g7�;�W�+M.k�
���h�š��ށ���)!҅eաj�V]��0��,�v��6S��y�*���`�!E�5�fn.���R��'KUf�bc�� \��_=anP rҤw���zy�'7�bM�5�0���Q�ݛԥ�ZJ�x���*Xp( ����� �԰h�7�P쿕ӫט��XڕJQ��mh���e��z=��vSLa��bC��sDn��-G�Cg�w��6�-��zﺳ׉f鲂8�Z�}�fi8�؄{s ߉ͤ
ͼ��\̖NUŴ��l�W�0Fk+��r���[�v�u�ײ,j�9��XpӦ]�k2�RΤ)J��wQSY��qݝP�z�[;@S����YlX/��4�0�Ʊ?�sk\C����9b�i.�����(l̡Ri�v�Y���(q(]=�y��rMn���ط��Q\��&�낞q�zs��I͍�20�塭Z���vn�1�J5��Te�^�$߇��>��[\�|�&q<���F{ ˂�/T��� �m�l����!+�;DN8�3���}/k"�䃉h���hM�����G*�Dۇ8����5+ �J=����J�x��2f\@�� :�%�wn�!�j����r���n�GV�w6��7MR9������ov,Kk�ҏTín)cyٱ�d�Y��v�7�m�@A��+�@'�@h�xW��#�L�VP9���RGk{͑{�z��W�^��z����Q
�dc^��F�NP�#p5{P��D�坺���aX�A�Z9���z�R�o��F�Î\���@H�h�νJS*m˛��Z���p�c4�,v�2-FI��6�3����ˋ�F��vFGY� �gV��Û��_^��>DA�T6%���w�+&.�녋�nX{����Do%r6��ğƴ��bj*֣��e�tkP�����n!ע�������q��j�H��t ���<zI)��y!�V�s��K�қ�����-m
�|þH	Ƈ=p�7��w��L���nv_.�松j������Y�����Zr(�>����I���EO^��N9��/bJV^�h��ʜ�.��@�����on����e���h'|�X������CpJTȩ+N�ͮ ~��^ޗ�|M��8�Ճv<��C����v��ۺU�W֯:V�5�/,L��[�ڄƹ!��Ia�t�������fs(]'�R�P�
��Ә�7�����U3�O.q�Ƹ�*�f�̀x�t����t���z)�,ց�l^�2�4� K�.^Η��[�K�6r�w�͂'L�����6d��+�=$hQ+\�\ST3�v�5�M9��B���-���<�� =����/:���v��u��oeg���Z���׸����
��S}8S�=�݊��[ꀾ�i�|�Gg2��13���4��+m���:����͊�ĭ'I8�!�t��m���A��,�[��f�F�z0�8$R00$u���Цn�"1�z��;%��e�t�or�Ӯ�2��ڔ�%����2�JS#�U}�iܬH��-���=Tm\�@�υXR.K�}�BF�1l�L_VX�=�� ����L�G��*tJ�)�ulO�&Fg.zma�����p��nzH�!�6���
 �<��4W��v�o�4+����j��Q�v�Xl�x��$��(n�qޣ6K�����i�f��^�taR�C�:I)�`X��r�+��θ/gv�ѯh˘�BaL������W<2Y�O7{�
$�`wW��:�z��PS�r-��M��E���7X��3}0U�Φ�(���}a��W���
&�^��ZPP%��M�%�g_\6WtX.�s뼵9E�1C�d#/iѾ��41�w��s��%%҃u�S��y�齁Fr�؉�j�>�|�=�j^7�sG,@<�ҷC��"�l����e�����iC!&B���2/��s�����������Ki�Cl��;͋|3R��[�T��8�^����[=��u��H�I���V�|�d����r�]�qf<
]������Åj���X�9�Y������v'l��� �Q
��5]�XY��޹��w9��v;Z�E�F��Q���@u�߇��d�1�ؒ���\�M �b�M���R.Wz^��%�t�8���#>쓢mw�Ĉ��-3��{����\�c���;&�Ӂ���?e���\O�,Q�^x��썲/Mm��1�gL]Pc��҈�6)&�wH��s.�:V��}F�n�bhʕ:�ϺW-e
	S:��2���j\(�ȺI�1nwg��jC�w����$�j\ǁ��uxn�����i��H�w����f%V�����Q�{�4�h�>W��Q�C��He/[���W�a�^�������J5��7�k{}D��&�Q� !�l�2v��r�#NI����JPiG�f � ٜ�^*�f�7��H;P�G���ĞF��wo&VM �Fr������I�9d��qcC��$�ZoI�!�l�Go��
2�}�qR��Dظ�xj�\y�:�fn�2Z���հ�c���˥�s��u��0���ϱi-��������}�2�k��؃������$Q��01㣥>����|�?-�AS9�.ܩ2O�9| Ε#}9����Z�y]�#�rژob���c97�oe�;�g1׈!��]9|0	-S��O�Q�p�aY�\1S�v/7n��kmy���p��t��Ⱦ�Ze��� �r�=,t�^eǻ��<�X��K��[��3j2Aqz�5*40�t/!%��ҙ���Ac�4�8����V���V���}���Ң��j�j���`wnVK�4цxeN���,�F�C ��#����ǥ;�#x(E��ܦ��5$/�}�����onn�Ь�Ѽ�m`�q��a�]SVt�K.�n�ٽJ.��b�c0��*)˼y(Y��x��'%�kسW$��\�1+��&a���6-T�����zU<����y&p�:�;ܻ*�s%fb��h�|��a]�7��M@��l20`;r�Y��qp��������cNw!��F�b��N���o6G�-����<�gP��'s�
�	�Q��82�փ�Ƚ$z��+�צ�
��B����Ojb�r��t���ܭO�0:Y]tg}4c�4�9i׾T����D�Ļ�M>���C�Fl�n�:)�E�#�b�E���P�^j�����o`�sҥ�rOv7e��l�"�����s+r�"j��^�ɧ�R,sU����Vyf���8B5����Q�젧N���q�'�Op��u�:����y�ݚ��n,���^��w�{lKtr��Kҳ�=��Sb
y�Q
��s$>���y��za�ځY����[��`�m;qQ��|�7�Zw7S��G#u��_PX ��#ޒ�G'a�wZ�+�\�d�V�]+m�5ʲ&TY�X[h��E(��@Ӝ:�u�s�>��^�@�*DP5��לּ����,Q{>a$�[j농�&(X��+b���f��[�v*TDPݚ׸���z+(L����Eu#���=)���<7m�ao	�)2������挟aꏚ�Q���*�4zr#�Eo#�X���2rΫ�Y���B"�!�����D������@�6Ҍ)j����P��8�0�����uq�1�7���s倭�lp&%u��9v��vo��
��I�����#�A�(i_l���VCa�7��m�_b�����w�h�e��Y��΀�3�Z��3O�ܹY	�')(մ챹���P�ᏄT�K�OpTxt+rRw2�Wd'	�9��wAm �]�=��4A+y[�������ION�2�k6®�t�%�m��xY{�u�>�</ps��[���/�cu�i9Q�s��$A�aC����Ed��Тq%LgR9{n��Ν�.�h�����Y�wuHI�ξ]܎�˲qN�<��W������M��a@yڤ����r<\1����=�-4		��(�R�r�M�F��d�:s��������|�'{����p��y6�7���(��/w嘀M�VY�m�0�2ɡ�Og�M�%���3c�&�
h�4����b�MGR���J��9Jv
�od��aҳ�ԍ�{�[ۘa�5
�(���XBjxz��oQ���$��m�E��w͒,�4끥[ʘJ�z�|�-:C�;3M�;�vu;5��u�ꓴV�QB�کEV�_���fOr��낑|K[WC�+�+���r:W���-o5Zڙ�W��t6�V��V��ɝ��MpT]�>(��D⎊�i�P��t��՗V񗝕��j@��k��%}O�X��+��yq��lFhoP	k$\�k
B����x2[�:��(�!��=(�ā��ĭ���,]�0p*)(�b����s���\�2kft�����\���vf��b�C����ʏn�i"�≈���H&-Q}o6,rv�b���4��C�Zt��Cb
�!R����cs(Yp�S[�J��������ɢ^
�;�Y�V�C�s��g�\��N8��)�[���Ԋ�]R�c��x���6@��O�T�|������AY����q_ayrG�B�7��Ô�z��zkS�,�NѺ� �K��W��[M�yc	ṽEh�ZxE1ӝ�~9����x���	����e;�媩jڽ�M땊;f����=cT\F���x? ǖ��P��~4$�V�k�/6���:�
���G0;�� �W+�u8_4{K��:ou��өk)ҍ\莛�,���;��7g�B��5��"�Pl���VpK�&�f�����u$d��T�q,��r�@����Y��.�Q�̷���:�J�i��]N��K����{�l̥�Pt���E�٭�|��ZIS�)����K�D�\�+)��t��\�f>��`��<����\{rKO.�c5�	��d̷����09R�,���^MŢ44�gX �Wk����9�LANE0UG(�͵w{q"aY0ä"u76f�*�t�c�Ԯ�P�b��>d�/c��v㏲��m)��D
��h�i>�=͋�4a[���&r���hMe�B8cY%��x�_ELhgL�N�,�D�Ģ<�r��7P���f\9�JM��_SC�oT�\��r���l�FTAa�v��`L��/E��;��:�{:�GY�d�]2-�J7��r���K��Kɲ����v:E�]����IOT�B�i��X>v{���J�s5I}�@��\�s��{y�,��31=�4�P�s6�[H�E�f:;��:;}v�i�Y�t�S��[��z*mɴg<�h�j��D��A��(�z���Z�{�/ke�u��	ɗ�mp�{����9��>��"�j�%:;�ukj�a��-���\x�y�f,�Iݻ�4�i��}�^�}&)˿��c���eTD��R���(��8u.ޔ�on��0��
������#\�YO��{F�"� sW�U���-����#���s�J~�\!4��Jͅϡ���K���S0f5��]Xl伱Gh'��H�^�l^�X�x6���xo����|�@�U��C�A�w�U�� ��Q\���L����o�
K@�r���:�����.����C!�C}�uc�E�J��qU�H��]qтl�Z��}��m��+��ͱ+/���&Z�wn��˚A�V��C�4�v�Zqy�6|s~�[�g�z�����6-�wD4�iED���|Ȏ�Q]��F̙wd�5�z.��V�Mv/MZ9���.":���v�%k>�.
���@����o82CVɰ����=�G� �xج2H�s�X
⸭N]չF�c �S]nvδ,�P�6����ܠ�S�2�o��!V;#.�l��i���NeY<���ܥy0��3��Kq��2�A�jc)�;�����t�A{F?Q�N��+]7�ށ�sk�w�ʺ�����^�ART��C��_��^ʪ�$�F�tU�}��O������u7í���+tJՉ��!�8^l�����*��55���x]�ԯ��� l����ɢ;;7t�	�ĸ��+5�Ka�6�j?�ZM�#���Y�Q���f>��7��2�fU��;,��҂3R�F��sr�Q�A�fQ:�m�C����l��@h�}�D�����tv��řI�%bnwp�$^w!�W�|�.���<�e��(����!��7�چT�{���/��R�&����v��}�i�mu�\�+�.�ʘ��g#�6R��˩r��4o*�JͰR�W�����]�����kv��%i�VQ:_/&!�)V�zT������������E]�d���v�̬|�T���h>ʺ�_Y��|�[+�b�z�V�dUۦ�`�מuoM���p�=���] ��n��^jc��%�L�.���Q�V�[��_>���dS:���6��c������3��xۘ�#���1�A��Bnt^D��=!crs��
܏��4K�ۣ��j<R�)e��|Rg��뻦�O>z�ʢך�v�y��(OhA���"*d-)�ݮ�Ǧ�PM�Y�N�"�4礖����ԕ��f4U
S�+R�Xo�N�5�o�9���tk95ch�L^��7Zo����n蕈@�t���+M�gfm4�;�&+����k]b�n��.�5�E�P]�(`쳦T��l�
^ym|e�DP��;���G1h�֮�;�gv�fD@��I90�2F�W�v��rRZ���a"W��P�skz�6�Qں��*;�)Ý}{�B9&]خ�H<ߎ�k�������Qoe�;7��\��}H�QY}�O�K�ʜ/R*������p8��[6'�.C�X������dM��������ȟe`ፗ���kUv�3+dC
�!^=�n�CL��}!���#��PqH�9hi�(�4R(�P�	6�G]w�S��h���w���κ&�Qm�ɓ&+�ShB[<�u������y�Rv��H�����Ͽ��m����1�m�������Ϟ����d�o�����RYw�i2�=m�:9��S4�o�k`�X��H)�������p:C.����]���$�6�E�� ��:���ne��x֌��"��ի��Βs踺�{�S�_&��;���{(�3���c.�[ت��[������u�׼ʛ�0��{B���j�J���t��ŀ����U�ޜx_:vhJ�C���li��u�W|��ԁ�m�+;�Z�_--q����]C��j�����!s� e��p!oS�7Ts��=��|8�*���5�m��^�:��A� ��� �����V����Я�R��)"me�W�yPWy}���mmw��aEF��g{���iA<��)�Zu�|*󮄂@��c1���::�s�؄YK�<�/R=/+���
p{��/"g�l�g%<���G3	�r�tvY�Ն�Jf+&��6�K8��٤�3�pρ�D�,c���Vѵ�6�����̺���I�BV�R�#��d�H�>e�,�Z���4tn^�ĥ���l��\���X������	Q�֦��0�S������𮧕 �
�U'ݸÔk���p�ץ��tu#��z�R���w��VV�Т��\^~k<VՉ�[^ ���Z�l�����{�ic$b̽/)�1�������'v��C`Wi2�d�.���S'D��|ٗ�k�]̚º�d,#�������b�����j���i)�ln]�;�ܽ�.��ʮU�C�	��J��mS69�=I�����qu��F,�+�ʆ5J�j)CX�B��ol�{�|��WT�h�q�%{Y6�НkV�7�%�4�� ��a�*Ҷ��`G�em����l/���S@�){�/7��ͦ���Xb�G2�<�Zѕ	b;��j]������EL]���^�J�ɺtV��5m�)���0,ZE�}ۀ*-f�9���(�u�)PҌ�j�[�i�C����Dv�fD(Cju�^��ͺ
�� �K�����$�<�����%%����g;�mE�{^˭:���ۦ�Ӝk'e]��Q�1�<�^P��|�	6�p}���^
�Y�E�7�ΤQn�o�I#���n��M!:��k�\��^�pչ�f����'��{(��8L��[�Zk7�w�'r�㜻���L�6캡Z�X�Ӈ��r�p�E�����;�#�eЦQ����.��;2�Rr���޼5��Ж1�9���Nd�}B)>K�HY�C%paT�V<����KA����1���ߍͩ�)��S�q8,lpr��DG%�+�,�Q��bP��dO��Lu��_W�w\�'U�ڙ�U��W�H>ۯ^��'�o_��m;�u�{ETk]>�$YJ�4�p�iq��&����R'm��GR�s%*�%��q��9�[���Yt�=���
�2nG���(o�[.������|���A�6�ov��Ν�7lid}o�x��y�����b\�բ�ٞ/E�֨C��_���ax��T�enK8l�L��[�2��oOe<�P1�ܝM���_X��D�TU۔����r�.e�e{��ڦ)�ntƆ���ul�1Z<oK����gNs郴�X�}٥�}h,�
���!����/_���bHtox�=g���Io��qmޭv_
�:t;�YB��v����O*af���ht�%�۔���C��R�|0��W��=�-��TyW5%�7;7F�����b��{���m��d�x�R(ٸ��J�Zs/X`+��-�4�=F:u��s)y׏(g�زuG����78���h���L��ycN7[Jal�к���<����ۇca2�t�Z&�b�F�_ۧ��T�'&&�k�SB���a;��P�t��1��fp�6SC˒�ْ6�[��S u�m�ѯ�צ��Q�w�D/3F%��<Wh�'$뇴�*��kS�8��t&�9��NF��R�ݜ�O�{'��ƫ����Ŏ��\�$��_1\��i����H�E�A\��:x�W0:�A;O%�p�&;�wQ3K�6���L�t��ԅ�Z� �=�:�fVf凰ٵ���6���F����U��K���y)Z�b�hh<�U�!�-5�Q͈a��oV�W�tD�r�uӾ#&��k��d����wZ�8r�� �٥.e%�ڀ&�]3��YV��WX�u`��-i)g*u+��bY�k'^*]�c�'Rسw, O�Od`U��F�&�tئ9�.:\�P��;�n7r�e'�6�ް�,����cW�{Kܺ��ǩY�Uu�V|���#���ܖ*:ü��!��锒�[��++s:��ø���7��!��릂���(Kf�'>l�
Õ�H�I�y��p(f�G_U�U��nZ`�˻�y��(d�Qӵ�{[H�+�m�(�.�H��Ve�A����1C���w�w}�
d�]�D��N�ª�#5U�]1�e�w��^���2F}�V5�×Gz�2<(��7��Y��w�Ⱳ�[헕z�'�����ڐ.�\�)�n���Xt=萿�+y^�A��a�y������na�̈́#���LZ=�.����U�R�Q��B�n����K	��}Y�^�t�9ڰ�y��;&L~>�u9v5�`D��5ЏL��gG��Ky�ː��A܆�NHl�n�Q�y�om0���l��&��=P���\��=��_m<Y��:2�nR<�/7��.���9+rr�ok�;�y�5�*��i��p�U�b<��Xu��-��bmӤ�6�YH���վP��aڗ��$nv"Gה��goz�҂����.����2[`�i��Pu_2:��9}zC��T�;-��;�[O�:r�WVԬ7`g�6c��7�dwhͲ�-KYU�����(m����F����V���I����.�ޛ�+((%7�[�5\�v.i���vN���j��uT���WJ�z�����N}4V����Cte�a�9��ұ�1����j��qK�L#���j-ߵɷ}�gg��OpkɃxP�4kJ�-��U�Z�M���F��*٭1V���N�ծHV ��Ǯ�:�⥈ʹ���c�g;yP7l�m!j���].$��1�
�ڍ�$�%������4@��Z��ٴ/��7q�ɵ�٫5�s��mn�p��y�q=��<f���9F��dXU����y����4��:�E�x}��O��k-�Օ7K��@S��y�Ɩ�o�ʎ���p�U�w���K㎘u�������KJ�H�n���7*a��x�X"�������ւOp�����i����{+^ξ����1�o�Eon�G��.]5�tɄB÷vEb���%� �0�{ȕQ
=�'^H���
�%��p��Ta7h�@꣟Nl�7ij����0�Ыy��gmՕ����� �.�k3E����6�dZ��2���`��ы{��O�1�i-oJq[����ʼ�K4��]�Q��T�۸�6L
��("��8.�{&K����q4_���qml�+���6��b����˽�ZY8�`�����hU�'�fc1Wr�!�J��VgJ�]�i�mC�[�ذ�{Kc�\d�r��gU�!CX��#�J�Wh��&s���tC���&�|`lWժ��.-sN*����F����(؂�n��/zOF�U�C������(v�[3���4ڢKۥ4�gj����v�*L���h��l �/�ayX5��`c�t��^֎c����[f���TZ�nK�-�����訾�7D8��Aw��I��y{v~jgr�s'k�=���	�o%�J�u�"Css��o3���x]LΫ��l�˭��e-��W7�wp��Km����#̖����ԏv)�0d��(��δ�L�I��/�JؑЩ��e�/��)��ruQ���{+E��Yf�Nr���e�4�L���f�"����^*��>
��S:���ږ ��/S�g��cdoJ�b���ތ7t��b5��z�{�u�s��L�r�}:�]�,�=�ULS1P���[qKa�z��b��4�axfF�My�a{2�����yl�畹��̓���$�RAl�`�~��oe8v�f�=�w�)%�z�$���)+�±i�%�q���b��̽T	�=P�o�Awi8�,T���R˅[���q�]ݎ��u�(���?Gg[¬٣H�o�&`���n*��3Y�a�7Sx�k��sX]S�M�����.�^)�����lb�\���<���Wk���&J�-�d�e'"Hw{�V���.���A�q4�(9t���,�Z�Ӿ���g^�w)���N��3�,f�L{��7���ʯÒ�̧�e�n���)Cp{^ C�;��o�Y�U��@파媊)K�����{ʯ�k,�Z)5ۤ-�G0ݗ�Lxr��xEm�8����`/F��t������d {�k�}�tCn��/���E�n��1:�-ڔ����C2|\�H�֋��-�����s�M�ډG�>��c���-p��t��_��	��"l�O=0�^]�n��ﺷ�>�ǰ+2VC���ٮ��S�a�}�p��魘GUń�(Gðs90���o;
|[��xq����K/Nmơj�X&��T7�i=+�Ye�/�U���$���A��Ġ;*�����$�v�鱇M>��V!X�ni����+E�,rȏjR�u'��.3�'�	&���'4��� i�ᙎ]J�ua�z �8��uǞU��(�X�6�ϝ,���e��:2t���=�%�v��	J歸uF�۸����ќ��Ig:&e�����C5ĸ�ybTX�k7Ӝ�Ai�ވ@V,PC����j�-�o,�V��A4�g���(5�k7fc�8ud�y�䀩��ހ�8p��u3Ҟ�����ޛ��3>8�tI$�t8�e��!6��,���K�I��{���\����-H�wp]t&�x&�f�N!����7h��J��,�Xa��j6E3t��L��ٌKk�������1���Q�WZs����P+���j8k�b�e6V^.tl��	W��
˽G���q���*Ȃ��Vo=�gdٯt���Mt���2օHD��c�e~{^��mq��@�c�Z>b����`R���6��p8G�w.�G�mGLX��2"�u�Xo�d+7%`�8zW�]#���vY���A��*��b�γ�M���H�� ��<�z�X�We�ź��e,g^P�k��,��v.�X�ᆚ����`�����ؽ����Q�j,ɇ����qO�Ȝȝ���x2���Ћ���U���*-]H���}��c9;�:�{s�;zi!&�P�w3p��p��#|�X�δ�n��}�6�hs{4����t�Z�#���{0�5J}E��'��Ӏ�g���`\OpM�z�ãt��)�A9V@�`�Blo+Uܼ��+^D�!�r�d���x����\�1��z�]V��<+����r�@�GH��J{;���G��h[鏘q�� �iTX����άof�E�U�l�Wd,�tjC���m[�x���2v��lJ<l�s�;��uf����y�Sy��X�#[y@U޹o�l��skD��;��2Um��uf�s�vo�{+�D�!5)�����9ݕU5\�
�@=��SexWx�Wo
G1E���B]-=�e%��ܚq��s�i�j�f,�2�ݹg��!�oq��&��JYU��3���*�Y�JĚ�L�U�W�k��Cj!�[��K�2ڎ+��!Ք��m�J���6�fJ&|Fh.Ф	7{�uh�gkUE��\Ŗ�G�3V����X�Z�a�X�]���[�
ޛ���[���#*��6P�uj�C�]f������u��#n��"�x�c��3���wB�>�3�o4�^ݳ�J=�BD]���Y*K$Vj92T��jih�6���3���'Vէ
�j�k�ػ]��F��!wvHr^ܜ�?"�;��E�}W���X�Y�w|v�d5�M=�(5�v�&s������Gu���Sx�N{�"_r#�, �	�Fc���T{:)vF
W�(�ޥ�vM^JסMR���&�P��贫*j�ښ�A`��Ifb�1���o;�D.>��`��f�E k~�LC��o?>�	���CKH�F��hR�g�l�tʾ��,Kn�7]��d�1�lс3i�u����g6�u�sN��<��^�ُ[]�P�� Ι�'q�����M`�{7
�U�ʽ�$���[�y����s������M�j�f.��X�{�T����.��@齘�����v���n�C*��b���X�N�0Ke7.4A����{/�0Ӕ��Kk�[���4�P��/a�j��a�D�ӲQ�̫�wyj��
�>&5�A^N���5J.�4�nf �|9�}-Ӷ�F��� }�I}�_g����b�|�&���3k=����,�n3o_V֛�Aj�BtV>��� ����#)��j�N�f��������jOU�"q��Ym�9ۜ�+�+�O��ћZ�&���U�4�Q�0��j�q"=�.9�H�M՘:���D�a̫]A6�Ք��:��:-v��ft�;P�m$�+l1;�[{tx�u����5)��z��(�'���!�.]vk��{J����.kǛ;��d��I���37�oaON�J��n�Z@`�u��;:Q�
���v��D,�󊮖�U�sU�µ}u-Z�_U�ҽwj��J�Yk�E�ҳ	#hn��X��C�Ϥ��z	ғu��,�RG��V�
�׈K��}����`�Q�k�0�1r0�C�2���5�
Fkc/���cz�����o7���o{�ƱS�,�%��S�n��x/k��(*�g��s�=�Lx�� �͠n�^N�RL���.X&�<��d���vz�&�b�m��XZ3v+�U�u+��1��÷��N��Q��w>V�[Caw��	��t�@��G��{�����Z�5�.���T)Ðh~�l�w.���
'~�/I�2�nL�r����r�"(ljL 9Ƕ�ݎ��Y斍N��g�g%��ß�=�%[�T�b�W�W�!�h�|���!��4G�k8���L�*�3����Jщ!����ۜ�1b�u�)�������z�H��g���PÛ�*`�]�()�5�a�e� �d�[���Y�zH�cK3�oa�0�zw��m��WB�+#��Ϸc��\�_t�0�0��1,�o�4�T].�n.��v��=�E>�*�>DR��ÓT�w���(��)��6���i��e4��ǡ�UJ՝u}�_Յ�IL�MI�}aF�zm��"h\��s�}<�NP2�E��m�Ԭ�Dڐo,�H���z&�<�Fj���T𡽔e��>�6�Z�>��0m'���������ۓ2G;"d����[��!2�hsyn��!QT��1��(�\ǩ D⼩����i_d�	؇��)H��41�7`b!�.�v慵ҹc�\��u�J7�5jN=�>���	zBM�mK_̇Y�b���,�
�V#Y�� �憑P�x�N�(*����2AR<V�"�s�4Y\�۝�(��Ȩ��%�G���Xyw�ĕQ^�8Qq�X*\9���d��8���ͅ�#*(2X��zʋ�%UaPabd�v���W(��ĸPT�(��h�[rc�� ��Ur)6UΜI���h���I�]�(\��i	٣�.30��H*���TQ�<q$�ʄ�%j����
��+�.p���G�<F�ĚN$�^VR�Er#��.r�-�B��p��$:M&�N]$�n$ȓ��!���;���'H"�H��A{h��\֑�[�(�Up�L�䊒a	�I�=Bpq�GUJ���Y\��Ok�:EU)�V��[9���h�AW4OR^AP4���B�dB�5N��CPQ�":��E*ĔK8\�PU0����hr*��&d��r#@(�2�MP
��|P �6�����f����Ln�Ife��w�Jؖ�����WB.�5��kujV����ɸ6j����L�qe|�+��H����Q��1 ;w���wF�U��'=�3�������˗�ޔ �U�0=���Vc������#�O<E����M5� Wa�B���na^w�.L�P3�L�@n�R��N�� *�G�u��?
�(1Q���E��p��c( �K�HV�m�75g������}�V��EV�*��g}�`d��>��3!���Xz{��7W�^�]��wm��ᕾn�ߗS�L'U޸��� �:��v�[�Ux���4O���]~�d��V7g�y�b�����}s�m{��u|���{��Vq�a�����:aY��l�K�3k��4~c�
���l�E!�iV��8S�����Y[�*�̓��v��J�b����� �M��$5!4>;k���Sڑ�RToI��U��W�
�3�^&j:]�����+��C��+�h;�MҶ�ŧ����2ju�y�rE#��[�>�C]j�<v}~d>2����%5�BZ��n��z�:o�<���nSn�Z�\��^�BЗ�>q��L���sG���/ww����M�Ũԯ^XZŦ_CQ.8'G�\�c�i{�ՋPf��ɸ��u���zn��΀�J��������C�M)(���F�S��(�`ȗ-�X�Cc�Σ�-꘩�%|�qB�_����3g�խ�*���;��b�c�lU¯��=^Z��ۜ��he]�!�_�Z�7�Խ0���vQ6��=*-�|t�xㅂ�gz%R�OcpO���R�ThL�S���J��`L�"��\�=��R^��k�>��Gé\���b�K��;���ʇ=��5e&c~�t�ۿ4�T]�wW𪽴�AU��;��/�nc��st��P-C	J!\K&������OG5Ū핢�Oё��D_���/��c�Z��	���İ�d8H�� �M�ݓR<���c�ٜ!@��w��J�\�C���Ň�;�^�w/j��/8�<���J�>��;YR53�{��ye,L�P�ô�]x4�{��ҭ*�u֎���VNG}*��[�S�7R��}ss�����	ԶĀ^Y�CN�.�>��>�o2���]�4ZQ�$���p�bɻ����i�|�֩�d�]��,5���I��{"(����C���sF�=d���"N���^��24ez2YX�Z������mec������ ���z�JΧ�Lom�_�YҴ���q��Nڻ�P�ǲ����w��T4���!��>~�g�ٝՏ���#�:����z{}O���g97�'LGI]��x8r9:Fu��[���J+�7ST-��PҪYk�+�����g�Ŕ�f�	T���U�۹1�3�Kq��qɣ&����i��ąW�a���O��b��引�י�T�n�P�d]Z�Ea�\1��^��!�Uv3��^�^@��T}f�:���3��c�G�q;=d�r�������{�f����Ӷ��ؽ�ŕ�_O>��^	�n���<o����z�2|o{�<jB����o.�B"� �:���Hy{B"��:���Q��kϟ�VԷP��Vu�Y��.��}�+l��pTװ�iW��p�]gC��c�Y�^O�2�{|�}8�`�*���aiL�5��#!�Z���*��R�P+���yoľѿ,�J��r�l��҂�xz�u���go6H�껷X!�x�ju^K�q��?E��AS����$����	ly���u)g�[�e�}�����z�NG���e�3�� ;c0�Z�ؾ�Uv�Ǜ �h�*X򎣪L@j���rN��]��	�,�ף *�\�<
�f��ݒ�ն"hF�ԭ�D�&������N�����og/�>:��U\礣�W�>[K��o�&hV�6��axS�m2�;�X�ͬTk�����	U�Q�x����ԉǲV���)��Ыn���C�Yp�օ�Z6���9|L+5Z;�vZN=齓.׮���f;���/��|���P�yrކz�%�1T��:���}=�љ[�um��ɬ�VW��fG�c��z*�]��x}CkŚ:b����;�<��-W^[�~O��uVxW���Ơx]a�oy��=��-��h)f�Ҭ�x�BqA�P.l�����P{��]/�xj�V��_�#�y��,cjm�0��դ"±�;��Q�vE	K��|���V*s��ڢ�"����D��v�����n܋[�UWk%�2؜!��)6TG��\Ŋ[ ��@�f�	Z�Z<�+a�X�|w,罎��﷐�R�����/�W�ʅ��y�.������q,�4En��uhѾ�	�V�\��)J����+k���n�[����M�=��~!�4�����/dF�U	RXI��/)��cQ�%�By��B�j��dC��b5R��C��6�ݰ4��$�����1�#mƾ&c�*��N����κU7����������q���|���Z(ge�/tp\���������`��օl��!��O��V̀��L�y|��k�r��B�Z��Ou,߹*ɕyq��޵Q����;�/�T��r��:�u�`� +���
����턽ʕ0�֦1a�q�G��2���9���ǜ3��ؐ��r��/����*H��� ZY!��v�d��
ZΙ�sw� ���'��b�E�	�*�ߘ�5�s����6��-���eu஗�V�+�b�
E���R;-�r1	̰On�Ȫ$5�.d�>;[�P��y��H/u��q���Y9+�~Οy��bw��;N;�^�S!ÏjXv[~��מ;=�O+�� k��S����t��x���׈�Mx�o�R����V��=�ي����P<=77���N�`�w�v]#�_m*��0���.Mq�]�ʭ�6��}V��6¥O�����\+<�brh�ZU:i|Ҳ�QVS��X�5��:���\�`D��<��*��S^"��i�j�\rq�w�ד���y�9HOM�0Ͻ�xϗ��OK *�G�u�O°Jp����C�(���X����<�{N��K��ƺ���P�����3�sx=t=l�Ɗa//i��}f��jp���dHe9��-�.��p]�r��u�St̐Q���=⩄)z]�9�Οp3z���Zύ�Z�o�`p�,+/������*:7}o�o����s�5��4�r��s�3�4L{�~ZW�`�Rd]q�+{-c�����[j�)SG*7��/������F�H�'Vܨ[>ݬ5����]Q8qg��o�C��w��v<]����]��gA���'�7�� ��	�v+��K3:���oqxi���&�D2<c�t�C}��+����<���?�Cb����gÀ�l����]��4�CgS8L���[lO���fyx�^�v���|����.��:������W���=Cx�G��*����v00=�;��>Ѭ�{�6��~���u]����cZevc#����`�b��*
;�>g6����d���>�<=`�����2C[֨��8\_>|(Ġ/̒NXOo�zvz�����1� �\Ck�l3�,�t�X+"�V�­��t�{��9�-������=Y������7`*j� �����$�G�E�|Mx���-C؆��['�X�������H嗼��dx� ��F���s�lV�M��v�X8g���M�S�r�CQRww�8�h�.�K����R�k~�5[أ(*=�o�b+~��K�&��~��k �
��fU��V��<*}�U�&<���x'���.^_��1�[:�v!f�˶0��o�Q�׺-���t�Gט�~X��rW��m{>����W�@��y��Uv��<����Z��K:S�T ��\�.��1���0�_e�����s��J�����)�}xw��]LXLJ��
٩��-���ޭt#9�vʔ�	��E�+%��yܔ}���z;�w;���r���XwiC7�,bv�{|��`�]��V�w+U�SwK�$7>�#�f_��zï>���W���Z��X�`K� �S0��8Cjl�U��R��~=�O�V�Ƹ�b,p��������ZG�^���G�X��V޵��{f���k�z�ݭ�5��#ʃ+�˖�*����V�x�xx���ӗ1��j�T�D��n���	�� ����9)c��>�c��Ua��X��P�j�	�@#I����u9K!M��6K�2���A�w�=��5�H��)Z�r�
c���G�;�+�s��������.�NUy��W��S��k�"2�Uy�cG�u��3�.�F���9��Z}��Y���>g�(j���CP�g��Vϱ�dƊ�nĊe76�K�պ����Vu�ġ���"�S\F�7�vð����(��*���M[��ŧ�%[`�ޤ�)�9c}�ͬ����Q���O	V�puᾺP�o=bד�L�]���6�iI�{��h�I�^$ƙ��
��:���1�f씾�˹��yo�o��U�|��b�wiN����U�C��y5�:A������1~x%��=��1Y���J�S��A���[�����B��:{�#��,[�%�%fͱCv�ŏ`"� r���04W	��PG����B3J�w��QT��V�h�j�r/�˱@H�4�}��{�E�x�H�*L��1z����N��)����c�:�\��Ǹ�UMw��wu$�ct&3s��n#�>�-|�z���'��
ï\��t}������9)�(hZi��`�D"h�Na�GZ��S������Y炧��԰}���2�� ��hb�k�'-9�塓YVf���\,C�l���d{�b�Zb���j�?IE��@����׹��&����z'A<>]]��3+~�k�o�>�ZE�ۧ�{brh��.�_�5��$��aκ*˦GI�A�gu�V��<�l���[�~_?+E�Y�^OX\�wũΑ�t����b���3]�ș|�C ���x����eA�2�1�K��^e�ӵ=�y��0�ݸ�oI;���kL�"��wlyJf�[��As�/Z�3��o�k��V���#��0�?e�+��:��Ј^��ۓ����1zf�	�������x�(�}�vp�{���b��.	�L�7�$N�<W�<f�zK�
�����՟��<�+�Դ�dC�XHF�aA2�!Ó��3�y�n�g=���bl��ya�����m��~&��|;!��%��Un����Le���M
�{��P��6YZ���"A�LC���
�?;�h2�wn%���΋���QnV䍄�H�]<�R�g��^�b��;*���vp��:���[���]I�+�V�\�+W>�$9Ӛ@�ɘ��n����1�~}�o�n�a�]�t�nY�ya��uKXV�#��n���T����o�"+
,�n붛�q؟�^y�O��ļ7���}a��-ǳj�h��E�J��m��~�+��W��{��3W3`=U[~s}XƘ��Vo:J4�o7����B�k�,��L�ώ��	�XT�����fs�~Z��мN��Y�vyHp��S�q����*��jY��G�Ǜ"��֋�:-ΆǕp��hP�Դ�FZ l=Kk/�]^wb� ��$���f�~
=U�}���c�k�q����Z��̛m��u&S4A�XM^���v�4tvm7l�'���j��?�7��g^�뽒��Cw�au�0���u��K��*��X"'��4���^a�&�.�Ug��QCZ�lw�|�Ɗ��#R�R����7v���g�sрO�6�W��v���X{����ˠ_�i@��	�{zT�:��HL&��7�Qh�M^�W����FÃ�u:0�ޞ�[p��D�x��M�y����o������E�7�f%ĭ��թ�ޕa�9n���mn,���j���{�IMO��v��Vl��-oQK�+^�ׂ��W\��*<�&1��Mppr�~��t4y3�����2�{�
uŀ
�?�u�����Ӷ��L�م����`��\�����}��1��E�3���SH�H��fur �g�g}�Z�mb�j�j�4G@�~z:粼q��n�SU���z]����0��~��U��Uo�.4]S����^����DTԭׄ��а��
9X�t> :��O�T����7gJUl�d�ڃ��Þ�Lrñ����F�E��Cb��=� _�d�wh�2�K�iGvKLZGU'�e?�]�E3�&�.�x���%b�-g�:��C(�ʷ0�%���r�ݾu�krNV�9LqR�2ut�}�%���&{�+��dp��X�v�n�_T�J��S<���(�'&۝Ղ��m�b�>˄�
�PP:2�6����k*!�~d>3��jgQ�� ���ɓn��{�0=Z��qo�	V�h����Wxغg8�t'V��k���slB�M��E�D]v}������X�ݶ�MW վ<��O��	��������.��}_ii�K�Z�C;�m�&���p�̲�`n�Y�#1Px�8�b5�uL(r�^t�H�e8�X�"y6i�ѭ�<��u�[Z N�[F�g�A��'��i�VY;��5��±�2�V�}xQzz�K�v�,ZGn�QҺ�%�d���d���'M-!n��x+��kL]ǖmx���ǧE	y{�9��R��	{E]k�����*���7�q\�9:F�j�Fې͌Y[���l.;�s`��OwV`�e���'kx
K�k3��K6����n���������L�uYZ�o���Zm�Y��(�b�uJ�m�heֽ�[��.���_0��ݦ^�U�y��zog��+�z�:˝짱I��î��(.��w�sٳ}x\a"λ� �E�ŷ�Q����6�kX��V�r���f�+�o(�ށF�(Q�XI��6�1�م��Y_B��]G�6�u��3 K3��,�b�Vm��, $)�c_>l#�7��an��|8S;�(�n�hl�ȳ�w#�]>R�k�pVx�H�{E� J�;E�:�/�-f���1�%N����d�����6pF��n��-���4Ǉ�c3z��v��߶�58A��#���y�֩�0s�GeYN�PN���>];E�A�/Z037T���f���)gv��W��:J����A˹Wu]���yy�-5ҫ�Dp`4�@8��i?<Y�D�s�^�T�%6�׵���IZ�XÄ.gj�=��i�+U���uB�"<դ7Vw�֦�
N1u�_��3Ld�I5Ep��c"fc�P�}�]�J7q�i��4ky�yΔo�ُ�!�f��;��&K��v;��_kH�:�.�*�H�ո-�V��H������I;���$x�"���2BiVb�� q�y�=g*�f����\[\����V���jW�ਖ਼�u�ԘzP�������t�oZ_,ֱ��\'!�"�j��H�1@C&�ݜ�|N\��rM�@9�&[nv*��矎h��	���v��;8�i��4�Kγ0�O��z�������ڏ�W��r$��tqZ��uB�p����vI�N�l;F�!T#��O'7��8�0Ns�9K���XW7C�5*�Ӎ�i�kUq��h�b��ֲ���:U��u}$����_�X6C��}x��{�̐;�\��|/����x��,3V��[-���J�mm��8��{�S7����*�v��T�W-JKED.��V�j��נ��|G�]�"���|{�A�у�W�x��J�+d� 멍%[�4P��j�/�-���-���mvr�A�00P93�e�	p�88[�Fl��1k�ź���m����3��p�0q��Q���R������f�Wy�Y�A;�Ӻ*☗1e>w7�4i�z;���՝Ԑ��
 ���ج�#%�����ӷ��^�̦%v�2�?u9[0�=�b��5�)\����(�uYS��nѧ$�ss�=�o1��1 ����3a�������/6��]��.���9��p�Ȩ�$��	��rU*Q��.TT�Q�9%��6AE��#������i���e$���Ehӝ��V��U&t����y0.AGDN�[�P�
ŋ9\�0��\��K	*M������d\�Am�*^	-Ee��8(�
��� ���NTY�(Գ�T�*��Z��L�/"x)"%f��5�+���*#"�R�K�J�Nj�(�S�����S*�8D�d�U\��@�2͡E˕ErMR*"�`�h����"��TG8E�	�K"�uidY�YPA\<BUr"��:AUՄq
�F��*��T�Adӗ�U�*�VlԹ�QDym.\�)˼����!EPg$�ҹ\�R��t�E�r"**��"V���ZPTDETAUU28Es���Et˜�*�Z\*Ι���
+�QFdEÞ��^P��5-�fTʩG^����9^2 ͑R�j%����~ ��޸<�f1��8^ِw,+��zpG�̢��ݗŲQ���Tb�w����1�Z)��($>n֝�3�������kv���ϼ���*��͑7�븛�~�����������8=�����x�Sq8��ҡ�ğ���{�x�~������w�i�I��x~M��>�q�ߞ�s���z[6��g\]�"Ù����2v�woqsI��;۵����px�N��������aw�����u$�^*���W�q�?��\��G/�~O|w��og 㾡��C�o���0�oΞ��շ=�{�S�lS�s��7T�����P]��&��^����'�߷���$�Ҿo_�tq	Ǉ�w����q	���x������s�v�
R�o�G��~���oϡ��hao�z����d���kxM�|N3�w�ޞ;���o�'��\}O��o�N�|��?'��>�~���iӾ�����x��'oA���Wq4�wN}䄚~��n|�G�9����`���s��B���"m�6�l��1{q�v�W���׊�|=�������ޭ�����>[�<L.��Ͽxy����:�_g���7���]�ͺ�@Y���=t<@�py������Y;z��LJ���t�hÙW�p��3qP��OI���&��ۺ���@�O�����:����$=��R�8�����n88��װ���>��sn����M����x��0}PW�LR��)OfG�����oϧ���	�|���BO}w�qa��w�>��'�Ǥ�0�o������L/���������C�q7�q��l�}I��C�8��&��S���T��*��y[h:�F���QYc��K�y��f�ht��x�5?���?��~�6�W�?|�� �����P㏏{O��p�0��oon?'��aWx���oHI�!?\~C�{z�����;N��ￏ�o�_s����k�oC�1v��o����w�v��}�sx������Y������O�w�u���q�ޓ��oo����:��O�oiǞ�C�i����y��Pp�R�~����Y�����R�45���gh�9����ggok�����7�!��z|C�����p�����q?�q������U�$���]�zL/�z9��q�w�i���y�<C���?�����@��{MRzݶ�o�N�����amM6^��N`��V�Nw���Ϩ�ǫ3G�O�f�:��-�r��*R�ٳX��S��l8���BX���U󵧪Ԝ�i�W>��f�\������#��l�6���$M����`�B�VN���o��TA��ɶ������������~Tݮ��OE����_׷��#����z�_G�~v�I��+����L/��p��� �s�>!�8�~N?�z��w��=t>�������C��8>c��~0vgs�����59��R�P�1��y篟=�7���I������c����X�o_`�z�����!�@q�{�������z��|C��{w�ϼ���/�SECk�޷o8�ne���p�+���Y��uǴ�a~�͔�o�H~�/��S���O��x��'i�r����@��{��u��oWP�o�O��������qľ�8q��;۴����ũ۟�Oް��m�k-�%۰�Q��:cS5;zݘ9{���b��.��2}�?GS�>��)�n�S���&7��vS�d����P�I=X����}���x�&^�?%h����<����+�c��oyO����&�ZN!���ۏ�~p��$>&�c���c�ߐ��=�o;��8���s�	ӏ�ר�w�i$�^+�v����wyS�q0��㾿������΄�<e�j����	;��Mv&x�]��|ᾧ���?s~w�~O�q�����H.��M�X���$�ohI��~����ԝ�=���<N I���8�q?~�8����!�8�'���������,�ÄQb;f�sLi'�?���w�S![|w^�C��z���<L.���w���ߓ�q����u�I��'��goi�>�1�����v���w���@����{���fN��Yo2��5�6�:	�^wf�ohO�}N��8����è�}g{v�F���|v��ފ�M�	����O��ɽ|��o_c���_;��ۿ���N��4������9�L/fr�w��h3Q�<]���١I?����~w�8���S��Ǵ��n���8�|�����=���C�i�O��X�Ԑ�����bM�	�}�����W����~M�����î"��{&��e��&g������{��aL/O?y�|N'����w�����q�=���&}C�޷�8�q8�S�X���:�x{�������@��oH_#����Y*~��ϗ���e��d�<��U�ӏ�,��������(�����_P�G��S��7sf9�����Q��T���
��+�0�/�$�����Z�aw�#(�Ӆ��6�"��K޿zu9V�!<���t1*����U�S-��UJġ���w�f`��f���?-�ϼ8�SH{C�q�s�0uӴ�w��~K��]�q�A�ߐ�[{O�_N	�?�'�p'�x�]������{������w{���ٶx��F�:J�j�p6�G��������J���E��_Ǥ�8��:���7?��'iһ�k���u7�'�?=suI�~�8���w��@��}v���`S~B}��=���������~�_|��7��u�t�3�����73!���#����x@q\��8x�w���M���ï�'�8�%�>~�ώ㾡��{�N�CϿ��'P��=�p�,q*�_�	$>&�I�/�5T�u={'.�5l��]���;2v���?�����W]��������]�@?����n;봓�������S
�z��9��i�:�Y���=��8����o��aw��}�Hqi���������.�VG=�"t��t�x?��k��4?�<���i�߯��P>���zN'_n�@�����u_'y��P����c�A�M!�����=?\�i�����zK���������_-��8ח.�r�Vˍ$��޷/�`�����ߝ����8�Q�zM<M�=�~�+���?۩����q�N�z��뽿�qǯv��v�+����u7P�}B}�>�������|v����Kt	/w����a6�y��]����;��}������˪�S{Bo��n'��C��Λ�v��u��x�}�����®O� �;���C�r2�@����;�!ϟ�sw$��6[r�ع�"ob�y���ػy�G�>8�|C�M�������q]�~~�����}wﾟ� $�߿�'U�������x�;^_P=o��}M:q���=��{v�N���O3��x�/�у-�Vѻ$�{__�]�Φ?q�!������7�}OI��QO��P��@}}��M�����?�t�^8�]��_����{�����>z�x��W�	��y��x�`�`�G�YLPa{ B��̸��=���C�4��������:M���
��c�+�{��o�_ �9oΟi��r�H5�s'E�;[�1�,�j��%o��y�rΡ���j�WjG(�'u�׃et�o��.��>"	e/���h�r7��%6�9��
L�o$I��{&o�6�D��3�:�2���ǽr�=�t"�o
�d�B\n������|bȒ�/�(r����"g(�n�޼�n�J�Ĭ�z�������]H��k��v��DC�	���'�k��;{^4�� �%=�w��q8��N��j��2<ϷbX�a�Xa�N��f���@�5(p��f���VE���.ߓ7s�-^RA]�|Me�<��܇�J���]aR}�0�^eR��u�\B�W�_�I"vv�_7�|(�ܸ��}p	�� ����W�-���n<#԰e'�h�1���}��4\�����cQ��B�6�.��,�����#�"~�Pc��Z����z����s VƜ�Ĩ����x�/�"ps�c/>���tN&���Tμב�3 ^��*x$0��'wj�_<���0o�]�qX�X
v�[��^[�S���ID�c�c�L��W{�,ݸ��ˀ]fPB�[�n�T>�¬n���pp
�> n�߀��h�ŵ�iv�t���4�X�v���G�@xڪ����6z,@��S�a� Oec��'f}�'s��uKs9+�[x.~�u�ڃ����u��.��:��xe�1Sƙ��4�ٷ������wX��Nٷ���(\3����tqi���uƎ+�)r3����B��[�ҍ#���U�u-	�('��h*�5l�AIF�EW��]v,��7܉s8N61�&=��W֝E�3��6���U�x��2B�9iR�:f!4Ьm�����k$�N#��l�G38t�,�#Hd����w��=�i�۰��0@vWr�+9R�kW�0��^G�Trs4=SuKPc�+>Ϝ'(W����(6>���"{�=�Q�e��ʱ�{�8���k71�.�a`zBz��l3�,�u�!��wg���&��Yh�:������8*z�������n�MW �P3p]�J�r��Nש���щc�C�z���8q�<�ʻ�DR�cY'Ҭ��_�����,5���f�z�[�ث Ug�t�� K^�M���\>���	�kC0_y�J�q���V�)�����#/,�J�NUFnީ;#�ת�Km(b���Tۍ�J���iF@�\H�!㣾�J�`c�궖ur�	���f�:M����/��>ճ�X�O�+��7K�����p�^�� ���x��k���5}�ף x�6��m�v/�=vT��9z�ͧ�$�O�B\�O����|Ӿ��Z��o�'[F��j�dM�ܷV9�ሺ,x?��^�O��yS��4��':�V��'��}N��`�]�Er1�Uϼ�]>h{v��
w�G����qQ�hq���K�`�+�\�9�E��uM eL��@�����ӛ�Mo��	3����|�܈�Qh�K�t��y}Ժ�KK��ڤ*#��$�t�-S�'l�c�37�����y8�Ux�!T���N��{�ڏ�Evk������W[�W�<e�oEa�c��Vo�����������B�~��<�Ӓ�c�p��ʨ7�'�n�s��5�B�/��B��/N�^�뀙�����&ź��ŕ���gi�dB���������*էt��M���Ng��.�հ��ь���>J��k����1�u�~����V]�a[����"O��m#��\Fl53b��Ӄ���ϫgPՊŕ���ʗ�k�k;�S�*Ί��*����v�]7�Z�<J��K�z��lV�x�0���^��n���Lى;���N��l�B溜�)�z�d��e7��`O���J�Bxo��������*��)Eh/M����V���S�c��L<�=�-檻"�P+����[Ǐ˻�c�z-6���ލ��G�<��2׆_��z:������#ܡ>�K@�CC<4�1��q��V(����44դkEX�[,����x�$��;acŏ[��z�!�VP�Cx��+}�:������qtu32��[��W�o��(�+.��Z�OM�������fηc��3�６ܒ�."V��,Ƭ�W�<�m��PH�ܬ��.$Ĵwl>�9(�3H�{�I�j�8�N�q�-\Y�l�gR��fM�G���p^e�����y��FZ�V\�s�!���􊫅�}[�ƘF��R���0ȼ�ʤ<y+�R���PL�/�d���?{�e@�/|ݒ��!��b���~gئJ��y��a�'�b��չw��<3k~=��Z�3Y����^�2vONM���u�]����*Ll͛�n�g}[Q{:��>�N�ԣ��XO��#�xW����44^i������t2��= �=U�~�`{l�c<n�@U�^�JixnYPy`��T+}��J����Rr�aQLq�@}Uʦ�Sn�ԏ��> W�7c�C��g��\.R^fR5�0���+��ct�/T>��	�I��,w3w�SnʦV�bq{mJA�˘�UB�lfe�Ip�Pw�|�r�!�i0?1`1�����l(n����d�*�ll�Pό��J©��̼x,-n���l�lק 3戫�J�EU���i����h{%^� :���~�e������K�o�6G��ٔ>`�^j�l�J����W�v8IO<my�g�CU�m��j�蚖�3tţ���Qȧ< ��'Q��&�G�C�&�aKN�Y+2�LX�z^�.7��3��&Um�=佚��e��qí�E�~�K�;9�p6ys�c���U/6NJ͑:��4�܈�� $e���O��^S�_}��}O�6N�k�Ǆ��'�����[1w�����}�>P!�I�F�y�O�į��ȋH�XA7;o�%3�g�����~~%.��'r"�j��}+��;Q����!T*���a�I��S�}nt&�Rƙ�L���pQP��UO��oLg�:��r��z�~i��a��=�=?,������b�,{�Zq�"ɩ��THkd�=�[�a��:�d�����S��m�	�Vr�<8�R����<��J��_��ƽ�Gz����{F-9
�:�]�$���r���#]*�/q�GGf�v�2pzOi��/��ܗ�@2�W�́:��61�y��b��W�Χ�芇UU��{����U�>Ֆr������f�ۯ���9l��N�+�x�^�s��?
2�U�7ތ}~��_p۟y?�2U]��ac3��Zm�km"���@M��n��ЯJ��Y�u���o�
��
����q�
�~��Xxa9~��^{}�)���Tn���@�`.��^}��t}�4��[�U �-C��u��*(�ў�M^���X�\Fְd�'-;ޛ�!��A��ep��{Bվ�;�ŷц"-��6��C`�2l5w�y��u{�Fu�MOM$���ЕjTD�Gb��To2B9̆/�M���㘓4z�(�`��!���\ ��(��ɵ�e�!�zv�9��oy��i���R9n�>%��_�/�ŏ:�ǅ?��Y���ݥl����5�
224������Z�xB�f��a���2��z�V];�OWP�
�a��^_ظ�q��߲���9��L�xr���%��}U��|�z���;^h��K�:��g��� _���<� ��L-μ�L�y�"喩�6T[��n���{=�*5n�8�Wd��C�^��#�&u{yܵ��,����p/8r�>:�h2|��^�{|lY1���H!���o)3�{Դx�!O�6>��``z�d��ia�������
Z� tcj�/,Ϻ���R�����uOnb����F��^
3��Hqv�Mh��s����6-�t71P�_�Y\ed	���/�³5_���³}K���gSvj� ���d�T�]w�ܵ�1��0{|
'4�Py�ܺ�ĉ}�52�g|�*�>�s>�W�D���6�T��>�Z=r�v�(csmm��Wk�Mx�n�b����a�x.'�a��(w����uf�{J��{����4��;�Ec}V��Y����u�h){jZ)p��)bcZ-�7�ȓ��f+����M��]]Z`�<��s~�m��{ÕwK!�	�Q�zm+��`��{t�V�8Ҝ�0K�v3�ҥD�F�[%M��ǡ)��$�]�8X�(!�?UW�UUpEI�g�Ag�T��S��v���.x�W� �N��!��&<��\��Tv���+/��FQB�7C�aqf�,S�_�.	�t]�X�ճ�1�^�E��]R�06W�p����@�oկ��.�,��𐻻O�.��{W-������lO�^�Y4�C;�Xփ�)�����St������\�^�k�t�ڭu�-Վu�"�,x:�>���j�ǽ3�ֶ��"�eI�KY^�[�T�S;��6�a��]���#j�j_���1�t_j��%y�-\�S���O���wĊ�Ϲi?hGL�GM�,u�g��?��]��s�KѻݹǻY�׾��P�<'��׀�g���B��P�QxYD�즄-�K���9�(�Ϳ1#f��N���T�U�;�����?�h��t�`�DE��3u�Ϙα�S<`q#d[�nCx�ig*���U�s3�Qg�x�7�}�z݇���+Ox�lɯ�z}^v��o�U�c���_i{Ohׇe!�kFQY�+C��'kr���fT�K�c�7O�jdK�����mb�)]�oX���XЭc�˾�Jp�C��&���-��2�[�&��rR�WY���/h��'0U����Q�6� dV��ع�*��w��7}���a�j�L9�"�%jSG���[��������;y���4�bxƥ��wgؐ�X�_ ��ٮU�m[���l֊�B(渨a�%�>u��Җ�>��2�L�ι��&z�n���X�J��G�6Lf���K�'it]�'���v*�:��N�9�vtol8��:��,�|BPv@�w�²qWd��(r���5�ٵ����WL��0�Z!�,Q9p-\�j�3�R;�4ޏ�w��:�<��+
�hZ�PO�*k��Dk#:��,J�L��m���Wtms��ART��w���i�蚄<�A��bG����3H`�Q�H(��w/�Q�[�IB�D'x�=z48��"��h�&E��bX	*���-e��9C�X�r�)j#%�H`p�b@���k�������k,�w�M�9z�=B���y!��ң+��G#]2^��o�Zէ�j��^M���M�(_e���m|e�eHa.MjZZ���,��SnI2���7��(+���I������|n���52��ʵws1*�R�ej-u�b=�PK��{�m,��R�j�5��)�Z+��
4�ͺ2J-i��e�<��w'AY����{z�Sϲ�t{�9�-�����CП*�G�HE��z�	uڢ#nq�ݲ�GC����K���rj��E�:S�m'xz��������f�AQ�r`�ܼ��.�bZ�����e�Yz�������M��c�&�-�5w�L�,�k��G-���y1�ů&��1�}}0X
��^s%�y� 졭?�C ��m��m:ySb����P��,��U�T=�[S�+Z��	h��d�]��s>`;�s��cSo"��.�{���g�����w�O�R�@vvR�r�����{�9�M!Z�ݛ�:�`_A ݘnF�Y��p�*1Ji#u*��:)vt��G(��כ�(���o��F�3u�.n庴�d��Q������ �
��v�E����צn�]�����R�.`�f�a�LGVmy����ʽ_Vmp�V޾�K���kTWع����t$��	�����e���O�Yk���a�s��H���x��T�ue��w[����[��NX22L�����R{� ���$��f]=����P�m�p\�*>T�8�j�cx,F�pd��.�ܘ�]��!�ϗf�����7$�	lF��m\3��4�'9m��-��C�[�"e��hO�M�*��Ƀ��L�v��P�%�����;��V�k,,�ڈ��]i�i�/��X�@�S�}���m�귇Ԧ	�u����N��)z��C�pyf��F�.�4q��uQ T`�4B�"�B�Q(4K���hWr7e\�DEU��(�Be� ��U�d9bE�VtÜ�r�r���r���XHY$�&�
�T)�Z!ʠ�������%E�U	&�$�k5$�W#�
��Liʪ(���)�E�.E�	* �U~$r�$!Z�#�s��	8�y��rYP�x�$�F-	3�9�Ȫ���(��p8�Y���Ï_�Qx���Q+Y*W�N%�P��)�Pr���!��8
��"���<�r"d]�\�uVz��GC� �\<�QȪ�"��0Ȋeʹ���v�9E��d��U)dE�(��"
O8K�ED�UPQr�9*�W9�I�ڙȊ�aBD�	�����*#B��B�q.�"�W�"(����^�OϜ������pL����=]��T�3�<�*��"-c*��=moT�l��&��X�b�\Nq��ܐ�s	��O}�W�UU����cf��_19Q��1}b�*7 T�x�pq.���x{�﫮�!=�3ݧ<r����y�u�L gU^{�>S�j��R�P?.��yo������DA��a(f�w�~�2uxU��D��/���"���qk<z|H�҈�r?�n��C���jN,D�^�9c16K"'չ>�eQ! ���m�l'ߏ��>�(�I��neYS�n�onz�ݻC0��B�Śj
��>��.�뮔Vi��Z+���==���y�yf?�.�ܞ�3ج�e+�|v��Z;,�����Yʩ~T�~5��4�j�
�ӊ�ɼ�u�	��K�Ux���z���ם?��	�ة�^Ô8L�^����9I�.��2z��<	-���c�Z5`k��ԩ���i�nJ�xO��~V��¼��|�o�}�Acy�c�iyb��*e
��;�iB~>�Y���QK�W
���=���Ƶ�L����Y�UZ�ӭ����< �
��S�g7"������6:f&�z�їޟݡc�`;�5\���a�nj��˕t�{n7�'c�@�{���\5�\$q����i��rvӤ\���s	r��,��t�E�z�#kf�\��Y�9���Xq:7B���vX�U/�`涟�F%���̸n�#�~o333z�u�M�I\6���=��NE{ @�f�ݕL�(�b�Ӎ���Y���Y��Vy�Q��W���^�F��W�f��[�s���?�����3�V�N���mY��O2������(���~	�]�V��2�}�W�W����*�ʘw��Dz������y�9xٸ����N�R^*��c����Qsm�A(Zs�7H��䫴���D��_��Q��O��{hd�[[��k˔ȪX1(m���d�vO�J�az7�˨!+������W�@�ʔ�<q:��-�8�s��Lǧ�aX�J
�*S��6��{j�����{;���ͣ$���9�_�~����)w�R�5lW��
�rƙ���cxn]��C���Ƹ�A�P&{,�Ŋn��PI�wmuꋗ|Ȁ�~�%�}P�膷/��۩�U��:��_�����=�G[^�t����rX�������2%�;f�*�p����uM�<v~{����rY��u�I^�`���TI��B�ƚ�B"�!�\�Q��'�����W�q1��a�5]�eV�Xjұ��M�e��f�{�ؘ�O]][�Ѷ�˻��D���a�8Fm_14c�lôs+�'.s'�'_�g�P6"��n��ޣ�ا+�C},P���r*�7Evu,a%:��)��ξ���u��N�ri��o7���o)>^�Ќ��O͓����V�� �=�D:r�~�=�Z@o�]q�����[e���e2���{��l���)��
�R�мwc�n�c�+�X}�������%��^O��W�w�-�֛̕GC�u2�$r������m��%H, V�����`v��]�
a��fb�����/:���'y8�On��c��_fT]�Y�,�=����S����c��OP��j��FQ�ۨ5f��H�P�@d-j�5>8�.�=�
���S��*ݞ��������)w��F��2�^��w��x�,�=��GNP����V�j�pu���²���vՙOT����=eq���]��pU��s�eϐu]�.įv�|���c�Pح�Zɱ�s��/.k��ס]ݙϖ@�s�*��7���~��O��%_�������V,�ߩ���l���i4��g�����9*��y~��wU�/��,pk _Y�\�
�̐��y7==̍^E�:ߒN������j�m1�0{=A���`�:u#((cܨ�l�V0y���]{x$��i��H8��at`ݴŞ幋2p��v<�Q+k��V/o�ö�����{���ʆ��X�pc���V���7�!(u9dS7���3�M�P��ݫ��r1�ͥ��޹JkT��J�Ir��7Uie]j��ܠz�Ɩ�V�n��Ϣ�������j/���-�,,Q�>Sr]��S��^��UZU�Ҳt��=��Ǐ�霥z�3�z�'�A���.�Y��W^��ާ�t�ٿ7`*j� ���rwX�V�{M˭U��LW�{�L������hw�*��{�׫�<H�Q�e��ټ�fb9N�jzu��(�і|S��bdi���BRH��]<�n�F�;�BH]u�#�(j��O�� 4�6���9��:�HT.����I�~��^�{�;��EO4E��D?s<^�ok���-��p�N%]B窰_ٯ}0�ǆ��=e�����g�F{��}p�� �e�-*7�����7$0w^da���)��B6���{]P<-���*�5�(�-A�e�fjY9S{�=�fP����>G�H֋�M�]����v��X|-�d�<O������Y�-�V�NC_�G�K;�1Jɜ�������+�]*�{��X
֬uih��%E�,ݫF�a�Cn�������:D>'��b�'(_ν� U{�!���p.�F^����}3����Nu�{�߫��4��(l+}�Ƙwyp
��Ry�v���F�J���׻��Ja�Y#\y�x���մv�;;r�&����r�� ��&�����$��j��U=u�Y秺%޲�y('6�����hC�R�"�Vb����8�Ƕ?7���y��E�J|Zv���3N(q��\|w7^g��Ӿ7e�6m�Õ�̴2b��w!����"O����u/|vr�K*���J��\n��8}����6S�Y�:���j5~�]qs���ZF��0�`�R<#������ʧ��a���[�:�i���z�G�6��\�+s0�@�9gO�2ܘB�U���j(�o�]�c��_i{O]j�l����ҭ�˫��ҥ���#�<�������������p�O�,n ���^@/��¨��Y��/nF���|uh�=�q����\���tL<�{�{5��>�[']�=�ʥ�R�>�%z���`����Լ���S�ب�xn_���D^�^�ǯ�@�O�pkw�:74�������%?#�XyW��m����;��}'�L�^{�N`�w���.�6����v�*�q�ʕ"3�D���@о9)�)Q����
�2Z��H�����R��϶�M>��ܤ�r��a�j�.�ӹ/�kj_|v�\G���*�-�R�p��x=9���3D 5`�v�ٯP�k��܈
R�5�n�YN�PP���r��1��\���;�Z���,�~��D+f�rW$^����C#��t��[���[XԒ��E]�5�P�s��PS��rWVt���7W�[�&ٜ7�`�U�Iࢇݕoa{������}_}���db����=���!�ϩU0��R��]�oΟ���4��:A�|�3,.�rF�[ư����g�{��)��>�r��_�>����(E�{V�7%v]c�=��i�7L�%k@1qwb6u֒uX���Ň�0�a�L:���g��`��r�<j4�7/�*a����!x�sme�Ii:e�5���݄\1Bw.��J�g +�%���7^�^�q�n-R�:�����gg>hP&������>)`���ҽu��x�u��ɂ�ڮg��N�>����OH�:L�I�=�4Y��!�ج;7�_��t�Os_�ʅ�W�k��I }��n���DD$����y"�w|�����4W�vxK���cC�/��Y��ߨ�>�G& =�ڃp����6��l\j�{��U���U�X�xp�>��?T�VA�,�e�NWt���~�k�,?)��#���w�|��������v����l.�{yo�][��tj0Ml�&��_H��|!X����m>�[������n�>쾞��yum���D�p���pE�%���]�1XI�Y8��x����]�vm��b��P`����V��V�m�ܰu�Y���}�n��	�M9�Cz�3���U��Y����-�����k"��[���u�S�R��Ӽ+�ҽ��Ch��kr����}��}Ti�7�b�����-�%K4H:�����rƼ�8/�a���v�j��{z�V��܀�,���鞭̀T����s�U��jSX/����K"��֋�:mf�r�g�~�.�Y�.����d���Lg]����;f�*�xk��m��}z5\+��"_V��򑉞ՏU�Y�*�
����$&�����i`1�
 �k���lrg��3�h�	^/�.}zV�w��jd-�ƥ6�v��yaD3B0�ŀ�")�;[�j�������j�L��m��5��PUg����8��Gw�`�x���@?7��s�
���U�5�F/wNg��֤9���̀�Z,�}�
��a��`{���0+� >�s��˽ف�W9���d�я�<�4[�o��VZ�'Xxzs�<kk{����.Z.5ޞ��B{;�G��^6�.��Pf#�4�6�6|j���+�<����n�J�[�VZ󆬱(����yY�J��t���c��Z�^�ÿ+E������߅�e�|�(�ɯ���o���r�7�Ŋ�k��F��+8�moqK����(
��ڭ}+aj��w��y��Q�{������l{�ɰ6y�WD1��<��
J�!#�p��䐷��h�)�a��j�F��9E[�3x��qG���ҡ�X��F�}��5�t�ۓV^�n9���^��o{��f��ʦ��3�
n]��<�w�*#.׶������T��6=�x}ۇ�]𾡆���gg���etQ�^7��,�}C@�����`:�x�zh�sZ����_���a�k��[���s.���ʯKPk�-a3��3Z�O�jK�h�@�<�ٍ�3�Ps��OB����6o<~��v3e�c��i��M<'T)((Jڝ�1�����T[6I��/�籊�d>3��I`Jk4���V�h���N���m��nOo�y�.�ѬP��/`�X�h��G��n�bM
F��`v� ��� '�|y��V(S2�=���M�q-}}~} �W�<������xI^Gp��U����]C�m�a�.����;�ŅG�8��4�o�ʰ�����:�����7�x.'�a׋��?)P�ۙ]G*�Z�����)��5柡+ęr/'h& ��y>OX%��H!Q�{~��?4D�J���;o�@���PO"z)�����V}���תa?^{Na�����,u�}�_����`oA�������IZ��^n�I�(���H�`aR�X��'oi�<xp�1d���X�=�����P8�[�e���<��ʷ�����Iq������ڶ�L9�F��`*m��Ti_�&pkV�1�y��y��[��J�A4��K {M�w<*�"���^×�<-���t��N��$+ޛ�����Wy[��8�2��W�������m�ѓ��uڨ;*���X�c����wK���(�O�=Fo]�'��D1S�o1�C�@��T��4l�S��h��кq�`m���I���P�O?9��h[����ħ��x����lW��>�Yh��<CWT9���]��z='싙g� ��禠�Y�8�p*��;��>�>E7����@{yE�`d���Pe�ʘ����I��z�J����U~/P�Vw��>�M���^���Mf���&����zo
����#t��Ռ���x�u{hR�k)_��(j��=���x]o�`\Nz.�s�||>��x*e��+�݃�M�e�C�į��K�{Ik>5�DJ�j�mp�ژ"9���}�W�{��U.�}����+�
�:�����Y̩~`5~y�~u��?�C�,�机	��l�O��n�̀�C^$����u�/��l�S<]'���<=�'�oݲ�&0�(�-`�P*��x�L砜����X��U�ng�k(B&s@}�|����ɚ���*]�6�R�m��WX�L�_�3ewn8b��h#�y�G3%�Fw�MϞb:W7գ��ͩ�;Y*n�xU�}c����3z����\��]�WA�������TW�x�?A����z�b܀�P(�bF$�I����n`ζpӽ�M�`g��Ԡ��"}[��%>�~�Eo`0eW�t�N�|�|��Ru�P�{�gJC=���С�o)�)Q���R߰
;�ڏWy���wR���n�K=̛lח5� ��ԡ}N <φ5�8;��%>U�bU[f�����~y�y���Uy�e�y���D��	����>R�����IE���@;G�6��y��3�s�,������2aa9t�H��{�[��2�f��Tϵ��[^�XȬ�x�>�R��5����~����ޤ�����~��s��2i𩂷�A웹�^�g{�������G7 ٭Uz"ո�*fL��:���K �Gz^�eAW�,�W�r/�Cߪ���/˨�I���S{�)��|���&��[���S�}�䜡�}���h̶:�yNOQ�|��ҟ�s�w��b�?w^�򛻜PՋF`J��;���ݛ�6ʴp��."��,���oA�x�K8h�Xo�h�8��Ak\��Y�uܺ�渹[�q�LS��K�ńg�����g Z�b1k^�˧�*���R�@$��m�l�ze��Dw<&H�#w��Z:�]>+�.���ʊ�P+���on^}y:�Z�q�
�n:sB�(���Ǹk'y�ê-VD<����U�a?H�����COS�w�H���V �h���	����e
w���j�`]؟B�:��e��QX:8b�J���t����)Ownpےw&_�*�[H,S*�����Uz6K.�ȨD7fv���>�yu(k�3S�gT�Y�㕋�ݻf�6��'ֈެ�c�oZ�x8X>#��/������O�f����V���P\��ub��Ϗ��RV���`�U��3w�>���-���=�s�9�6��J��t�KT[	0��ki�&�e�[��_�G�@��s�Bcޘ�|����P�lۗS"����w���Y�vLM|��(��'�W���w�][���]8�ŷ��PR���ԋ:�D3��7td	�ǆfM�o-h�<ȥGV�F2���]��Ř�n����>�Yf�5- F�+���-���k)�����\v
�=B��Rgu��lM���\�V�
]O9XjX���9FM�t5ku�2�����0�"qC^#`��xe5��9,r*Y���)��l�e<
�K�)w˗aa�2C-�=!���Һj�`LaW"E�ǯ3�X&�I�u����&�3���1SL��Z�(��p��/�
ۋ&��j �̱�FBù݋Pz�*%lx�/Pc�u�k��v-d����l��8]%J�3L��.�o�F��x��x���GI�]\/q]�W�w��}2V����Mb��ghp�\�%�w���\���R�kE���5�x3��s}sR���f�a�:c�V�ܫ�#�s'v̐q6�@�/o-(���{6X����f.�!s�v���\1>��(���GmrR隕���k'�G�ttUp�X�S3v�H�kUɷs�"���7KǾ{��%�3z�lݬ���k�� z�`��:~㤇�wc��Xm[�[��q��l6�:�甩�)�<8_:q_2�j%MͰqݚ},!b]Nj�\V�mS�BX��#����r��tU���q�Ϥ|v:y�w���u�s�טQ)�[B�ky��:[�N�ċ�%��f����CqT�Z�Җ�kUB^�(Y�Q���ma5�G�~���M�Ae���
@�+D�+.>t\CN^eE��+:���&�e����������{�4`�8�uy��'�t�{y΄FF�T��*#�TEQ,��D�5#��p"	Z%Qp�B �Ap�����E��]�$QiHTPU�MZs�\��ESG9/i ���9PQ*��4U���PADs��*
�q��EJV��PEBB\9\�Ps�d�VU${�<�TQU&�8U�rIyiA��*9TDr�^<y�iEPz&�S1��tDTN�8�" ��G
��r�Q8Q�M.U\� ���g*"�d	p���)��7[*�Rr"�����ŔL��EyB��"�׎w���<x�"����N3����^D�EyGmdE@W(����aG�!�ϔ*�7Q�b�i����s�UDȮʹQ2�&.P,�J�����YW.N2��xʢ .
.�s�孵��!�6�]t|B�f�ˆ������a1�Z�T���S����E�(�vdbX�(��wO���������^�<�z�E2���4t}^����{l���LB�O}��׼^�e7�tA��յ]��h�����B��>��C�i6�V�Ƅ���w�s��s��g[�>J�6ǣ����2��uz�/,lE[:�h�ߒ6�(�-����u��������ҳ�?��G����O\�#9?����#Y�ڒ5iz��Hh��N���2O
PN�öq�^��!�M��P�96^Jq�����Ce�P��y,	hf��b��J�(�&���ǋ'KF�7���}��R�u{g���k)�n�_n��*?s��b��X�ؾ^{����a8��W���6CJ�$�Pm�k�)��<�qQ��2�P����z%91G��O���7�+YM	�mdf��!F+���4���8'���V��������0��&�~�Pw�����7)/&�e��g�Z�l\H�F֝��n���k�W4��X!�.|� �撯��+�x��2�K&��) �w��	T�z7(��:Ҏ���7?�6�
�c�Ygl�V #4,��|K�謨��f	z5F��"��#�mu�r7�*|�y�,��*��۾��ꪪ���Rr�����P=�����Mͪ�p�����}s�M<�L���m'h<n��x�K�-"�_�<�(��;ρ0yb��y�g��6���y�թT�J��jG=�j�8�`�ڎ������8x�^W�V	��k>�{g���œq7x������}d�}� nO
��:���a����t��.�Y��;�u�/d���T��ӝsp�����D�T���-e�;ƌݍ�����t���#6Z�%��:�s�uU{�1S�gkj{޶���m�_����>��hi\0�2�W�~�޾���x�O���\��H���l�]��m�薩�g�,�PZwA�ĩ"���2��X�N���צ��5����U�jl����WyΡ��R�(o��������0��*h�\�S$�Y��4�`�L�H��Q]Ԟ�!�6?¯	�	�K�M�O��H�ںȿٝ��^kq�v6��	�[�h4#V�VR�A�c�һ��z�Ѐ9B�A��U���t�6ba!���~rguF��{'��z+�����GfX���T��D�T��B�f�a�����]Mv��	���W�}��V�%�N���$��揨/)K듬�*��+���Fs;u`��ѩ�K;p�<|���7͏���<���7���ʒ��Wa�@}�����n�����Y�� U�Jt��zaw'��T</�Dב{]��g�k7
~�õ�3t�Z/6/~d��K����]��y=��0wY��֕j�P{GF��≼�c;�y*�^�>�8���޾��p���^�8��453#�k�Bܡ&嚮�����P���_�&R0@]�&և��<�b��~�{������m�V�ٻ�bF�������_����T��L����yr���1���>��7^�6?��۽��B�X�gޝ��K�u��q|�a{�`�_�硫u��/K�#�?���=�rvW���OaC����&�2�������~V}���c({ ��3F����j+G��r�1Q��TUt�)B��n���8�V������ű�ٴ��3`5��19�y��KR�'��\����� P4����0�f��+�����7V�r.��E]qRn�Q�-�����o6#���%Xv8�%[� �[�j���a�"Y����_8������]J:����3r�7���}#\|qt&��&�xs���<���Y��P�q�'�wD��)�#t�J9m)l���f*��1ƃ>1D�-^�E�ଝƉq&d֣sr�E��i�*�r3�AyT��f�o%C����y���`���+�۩��QVڽ,�wN:�W�TRT��@��{Z�-/R�; ��ܩ��u����W9�Ǭ5/ͺ�F>�l�#��b-Yc�r�f#�f�DfN�E���+k��>{U�N������݇s��J~�\/1��^*�x56�26��4�Q��x�;��A���!y܃���{�����I����40)�6dN8h9p/�w�Շ���M��Z��1ک�W=��i�L�����J�L�Ϭ��"M��;}��=��~��r������n����ޑ���]&�r=hL�͑���GN[�R����Ѹ���~�o��f�K&;�����D����TP�>�[%.���ZZ�qX��U��[��T��\7�;(����L��1]�W�[�u
n���p��Y&�G6��rD�V<�VA�{�o{�Jm1��5N��Y�(�T�yp����W�V�U�S��Y����"��'��(��Ҽ	]@��m�5�2f�M�ω
K��]X�(%f���z�tm�FvM]����׊�)[��{���%��9��p�G���^�X�=���^�&-�{�0u)����>�R��U�����/.Q�y�����)HS��>ކ�{l���4�J�i��X�I�X����^i����������K�W�����F3��
ΐ6|z�2)�M}���BS�K!�������C�半��f^#6�3�z��5���W�	�>����j���X`��V�:�,��;��ZZ�U���52c�naIc��1��+�L>��k��P�<�GV�"+�Z<��7�┓$�����]1�*��޹P���I[\ߦ�x��K9|Q�G��������p�Lq�n��mf�Q��݆����IZ����g�h�����-��b�ST���+'ש�W��;��L���r�J�����1/�u&e����**P�9Rk9KN�4�:c��&l^bp�ﾪ����������;�Rv�#�����k�*Cn�U�6���q��=^��ݦc���);PU��dwd��6��T���6젺0�J�w<�>7�چ��!�wI�lʤΌ6�c�2���cR�A�zW���@�F86h��R����zѫ��M��N�; �CLSl�V����K��X���<�$��ݯa�$���kl��3{cu<ϴ�ZB5�[�UY�lR!({�Խ���|Ъ·�3��o��3��dȵ?r�Q���/2qz�Y�|ARE�X�jT-����5Z��,p�*�{�̆�"�Z�kaHe�;��a�KZ/��\j�6�]�C��5-K	ݼK�{��,�> G!8��^X�}+����4�&*y�;^����-*����^hW��$��x�S�K}FQ�/Q
Q���y?Nz<0�S}ٝ=^n$0o������$'KX7[�3�Tv����)1���_ٯ�o6�SD^3��4���B�]�cjf�Z��L�#vu�{�i��r:�/f�j�\�M^+"U�\t!��'��R��H��8f�[�w�CMk�k��W��[��{�fh��M�D����&�g~}�0��q��B��������i/�K[�f���p5a��K��$St�ό}��ӈ�2�Ai�'|��#�{w۞�Nk�hrJK�S�w�쁘�,��tN�>�h�hZv��I���}�!'ysk��{��?G�Y P՛yI2�t��A-#)3��H��-;x�e����n6"�4>>����g$*N��J�y�����
q�z��r�[���Na�[�S�I�2� �Zٷ��^��ڏ���Dd�:+��A��6���@3ܔSW�=�[W�Jm�@�@we�cگ�秃��.�M�R�:�R�:�����$\��j�"�l�6�\*���A4b�'OG,%���3=���^��ygc;�y!p[8,f�
�ǥ���^�9^@��c�Y�4}���cw�^�h8yfw~�"�e{0���K25�yR;Ə��B�v�P�ҚM�<ܮ�kr���GMkQW��<@��M�H+�:-F�(.���b����2�,��oX�����
�\� T�3����޵p��9������կR恖Wg�����$�3̲:v�#��NK��uS$�R�"�%h��o���;�t[�aj�����y��L��r[8�J6eK^Ö���Le�ם�ۢ��>��c#���a\<�-KU��5��p���^2f�["�����c��{<p�K�����]��Sm�� �����(���������×�y�8z�����䇷�,���6���`��l40��2��Y�k뮨2��G|�L�^m���Lx5��T&��o<Өa���<1�д\o�y���FK�-*��G-�-���}ӕ�}49��Wރ�m�;�bS��r3�� �s�p�l*��j;	f���)�lBz�>��Vb��i��]�zC��Z�n@v>o�z�lnW�u�{D���L�:9�z0f'���%D+p\�9�Mc�d�o��m�8z�:y�"�,�x}&�V�hAb�II|�(����|z�S�!��r�e���V���y����~�Ow3�X�s�2���\�{{M�#��zgZ2u<>T@��E����*ăWd._^�X)zq��&�30Љ�:;@�Ȏ�b�� pe�����3�6�A�d���&�3��T���q�oύ��|�#|���r�xv����A3�����&�x^��`�W���y[���xm+�h����B�ÎNH
��Td���u�,i���`�U��{+ŁpK��@��W��W����k2��G��$�8�Qlg�XA�|1��2�n6�l�����M��M��bo������}�J���S-���HumJN�
+_w5��l��jH}�������x'��`�s�xT���^sa�;�%)mъ�j�j~���r�a���v��.Z�8��۲��Z=�Ղ^��D�6yz[�oO=���>�`ც���(����|��¢ؖ)݅0��v�R�i��l�[��B���m� ��3�<�{�A5�cmd�n$���J�!J�pyi�M��>8�Bn!���g)[��CD��gr�偹0W 5@�CKΝWJ�C���قS*�G[��D��"��R��VCYo`�{y�[��*b��WZ�C}��Cw�5g�50Qq��4k��C���2_K��[ճ-;��J��k�����)��j,��dޠ��������	Rȵ�/;�'&��m8n	�A~�D~�O��&�q�o|�O��ga3��ZN�ژ�uQL'5M3�U6-�Vy"��J[T�� 'c�m�[(��Q�[-e���o"�y�5��i�'��w֣)��S9o��F�X�ݦDK��q�v�y��J�ʩ��U�W7鮌b�5Ζ��=7b7�m�p�o����Ъ�=��1�r�T�TsX�4
��h�VQ1iMQV�vQ;W�0�[��ݖ)k�f�����*VϽP�Ri�o�x}��-�1'�Ǭ��m�^�iN����*؞U8x�������iچ�E��Gf�Pk�/5�EU������1Y����a�ӻ���i�%��Y�2f��Gg��ms9�|�q���o���9��vugZ�W�P�k)�[d�,����r�I�j&p��0�m�W�߃���ne��|��Pc�,ҥXxk���jw)�	���ڝԹ�b���G��y��.��4����rjC}������㝂�2;�!P�7�NQ� ��n�}3L����s�R�Ԩ�`��]�RZУ����9����t�L-3)�.�݇@I�t_�Xl���	=�[SMށV�o*�n��p0�<��ݓ
���i�c�Ez��)V�֬ռ*��c+s;lK:�#tͦ��/����Q��g	��[�z���K�V`�$��1��R��V�[�)	��΁[���K83�w�8�V�H[%�mٹ��,XО�����Y��ep��i����۱ȴ�OH\��1^fv<�����Tth~cd�g���=�śW����/��).S��Yz�Ա
��0�w���v;��|5�I`�i�K&��B�(٬���|iE��rݣ�y��ܚ���#͞hӐ���[V�ջ|Pn�6v���P��F��^���
|9ڭ~wR�����	��W�Ok,X�}�n'ٱ���(:bd�xs*`��M�Qgs�i�7b+�F�RX�/"�Q5���DWZ���N!�3^���Ӹg��Rs"nY��
��ZȒxGp��%[���DO�<��I�Y�,e��8���U�xrn����IQ�l����<⥾彇�0i��n[ϱ齮����ʏ5Q�.'��{\ԆP�Х,�]����ӻ����l�8� ֕����EY;��]�˕l���v��
������3�wI��E��h�gb.�9�F��7�i�g@"¯6r�{�,=�I��A]Ӕ��H��R�cu�M�`S\��P����.H�ݥ��`D9|^h��$�X�/�f٪][���)�V��N�l�.a-�F������+0f]�]��i�d�v���c�8�9���_=���?�*�y ��l~Zsz�i�vAp��V1�c%��s:�����`yȮf,|����:jĹՖ�Yo6��M�p;#r�Ц��se������WY=���Nv�|�^�',j�Ԟ�"1;]��ȠTZs����ФQ8T�U���j��d��+�)���ރ�`
�Z]��$�$�އ����iVU��߭�tb��<���:fNu�;����/��T�S2��Mw����K�ؖd9n�{|C/�������z�.�ba��nVh�pˎ�-s`kv8�kC�ro�[kx��oU�L�wF��@�L�J6o7y�L�r�r��x�{:�4
���z�7n��h�&��F�fygHG-���6E˻Щ7���\R��]�z�n��Ky<\��giuR��!U�e�+MnU�}7�b+d����I}5��k]��q�:��؊��y�N��.��gV�yv�+\)w4̭��R��]���ǹX2v��V|����Y�¢��r���Y��#jvsg;��Z������VeK1l�yk�{cQE:��\3'S�l��޷�Sz�u�u%��^cVht�*��M"�BlN�d��ό�q,�(]�PE
�S(��DJ%��".r�\�JH.2
��U\�R���*|��dD\���/+�D���q���L�z�\���YTEC���㣉*��ed�EQ�TTE�	�)��.�v�U���^�\�W�A��Qʢ"x���'��+ȅr��*�$��H]��*��%r��ѧJ8R�x��P�"���B��.p:�p����$����9V��RE��#QȜ�P���)�*��q#��ܱ�PD�$��q�w�8-�A�h�Z3��x��{˗;�Ǯ:�G!g#��@um|��E�$(�(u\��<�TUDS���E\(u	I�����~�<wm��x�	�x@eM��N�S��h�4�O)���쀥~��w�q�v������V��u�9���33>o��O5zu�ӟ�6V�a��"4<-w�Am����j�C���K@l��� %��:��`L���Z�|���[U���C���V)ڴ.ֵ�}��%C}��#k�&���JVUs�\ߏ�zZ^D��fF�2�BA�kޅN���x�����
ꅬ�n̵��#\��4�$sY{���(���lTױ�r11����+�M�U��0�>��������G��.2�m�x�aN��|ߪ�&q�-��Z�++��P�:�y���#�Z5j>-�����3"��)�^��-����D�4V�C��^�{���,��C.9���(=֧��+�B���� s�;�Re2�k��M��bj�Ɇ[ V�ڲ��^��������V�6d�D+�.��S�|r�\��7z���/��wS�m9���=[�kw�<�E����M�c��nO���z>U�EG����[��³�<��^����l����z)9�WIYzX�b
�����wu|3-!zb��ǜ`�U��穧�o�s���T;��c�9�/:���N����aͷ�d��*��*]�l�*�;zvɐ�јf�b��XP�i�����i'=<��?�W�|r�Y|+'�q�g�	Ēo�)1�"�;!��	��ޣ�%���^��B�^V��^`+�W��j��/3�B��2{ԙ~���>�����8�4=��y��3��'��VX���w*���&[/s�Ȓ�)d����s��v~�3�gE�@��z�Vݮd�=�q�3=L��gi�͢���L���E孙a�e�f������^������5���]K����S띗-^ҟS�����5� ����t�~�Kg�
����Oa����<g�u)Y\�ޓ��Ka��'��2}�5�9E����~�G��6gX�er�w��eAm ��|�u�"/w�@.� LT��Z����l���hi������3�)=���Vdn�����s����ms���p*��B��8E�����:5��׷�zVA�7���AdCx�jT�5u��k��z���Nޮ��1y8*�+ݷF��	Ap����2�`W��d��}Ky{E�#+�n�n�S���KՀԩk��r�p{���UoC�������tWc��)䛶��v{ȉ��0r)�+"����oH՘�es���{�5n�9�J��e�R�����ͫ4«$�&w��|��О�?A^b>��}C#�PN�S�y?F{�}U48*���z���d�M�Oh�����T4�B�Eeo�mWy�*����w��"����-v��Z�;�F]�l?=s���_��m{­�Yj�U�zh��{�#;�="}��j+�:���
��o����I�G)�+pmc���?E��Ą3t��?��pZ�zy��T��l�=��n�+E�����V"h-��:H����nb# �i���4���(g�;h2�J'T�z[����qy���R2oүq����"�/���{A�ؽ�z��5nR�m�S�V1��z���i��>^=�z��M>����[��4�l;��NM���n�WkhVw�" }�����t����ċ+J��!��ƫ3�7{�	ҩ��³3Wi�$< p��z\4��"6h�R=�����&ŖA2���XQ|n���FWd�!��Vi0Y;z���x�t�(wiPT+�s��ו3����+��oh��X���y�ޑ�)��}U�U�Ǚ��s�\�֔/��Y|��{��Sxgd�ګG�o��9qZ4^N���)����LԦ�I��7g��s��h>�ќ��j��̆���1O�gI�"}K}JVs�]�p��/Dǚ;�|p�zHW��b�
跬���y���[�SS-i�㪶���զ�Ť��Ƹ���M�!f��[�љ|9-�1��2�_RjS��-O�6�sGR��E�
�1�J����mf���3zz��(��M�qjf�Մ�>t����M�,	���e���-p��Qߘ��y)���S����P�<�OX���7r�]���"���S�ƽ��{­��Fe��*G�-;���l
���ru4V��d��%J)�V�,*
��~�*�͡����A����Qƻ���$�vz�&�|����<��y;���mr�'�B�Vo9yj���[r0&�ٚ��9��n��[�Iw'sx�t��_��P�b�`f����!�Y��Qm�(�ؠœ]�ya�̐1v�zs��(�JzU�ӽ�͒��_=�dP�]�uқ��)��b�~.hw�w7���7u��|&��J����J�ۤ?��搜xE��}SѺ*~ѻq@>�2E\��<�v5#�3\�2LbB�ׇ��)��`ѡj2h2f��9N�`ǯA˺�9Wt桱:�rMx�H4s���Y���K9�r�w��V���k��k�‿s8h��.��#��u�~���"���ר9*Q� �)T�[x$������f�ky*֒���������V�е؂�����/c�b�������/?N�&�q��{#��m^z�u�g����w�޵��墧�!�C���R�y�.��t�B$��힓Ϩ'�8���қ��kb/��YwU�H>�T����7����e�X�UGܽG~��W|�yh��AX��2x�8�ב�@��}��I���R�����2�-KYm2���Qx�w՞%�
�QN�H"^8�&�I�4V}�Өa�C<���c�}@C�>	F'u��tٱ�9ia�2���y�䕌��9��}�牧:����mz>��>K/|�v�0vȣ݈^�w�ܚ2]�M�`��qT��=���΋-�&Nj���3�w�9b踽8���2��oq���s�m̒��W�W�x�a��>t����/�y�dl������)�b�VmJ;�DB�ּ-k�J�rm�2Ǧ�(%)���О����탔�)�blYU��N�1[oΌ�A�"�JW���{E���w���8�sq5ꄥ�t��J�k��If��a��������A�HY:����c�+7��㊢M�.$��)��v�'��I����sύ\d=��N����s�3
�*v���2����'h��T���j�]�^��Ýkb�~d��WL�)�>�e9}�y��=�K~7̺��%���J�<j4�c���ƻx;p��*R�K�s����6I��VB�U�d��i�S#5����n�n2�$��Ң�R+3f�׶c^�-��Ja��>"�a%l�8{����N�}�f�Ug2J��Ey�T{fU�r�S�d��k!�d8{̛����XsA��ǗSEc���ʇ&S�1+�9�ү��G��?Q8���&���;k��E`�^���iH��J8��b��>�"�f؃%�7N�Q i};/�-m�!N��[K.��4���Vb7m�?��jU}�$��
�BG�$�iڶ�iY�����am{�H�/U��P�g.��;��ݼ3��f��&Z�ըsofm���Z�\�kXZ�(�1-�e���j�,����|�W�{Q���-e�O��6��,�A7nɚ+��M�.A3}�H��VM�}����xz1�
~)�.N��lo�c���n8O:���N}鞝C#�dQ���OD~���}�2'�7d��t�k���)��y��h��'�1�\~hі}Ұ�G#N���
�!�Zœ,ժX���z���Y�V��s�cGގ�lTW��kG܈{��Z�<���p^��3��:����j�J�s�E��=@���tW���ջ�zN�f����@J�g̹�dJ6ݴ�Pl&�T[T���Z=�����Y��Ǻ1��)>��狸=E�x]A1��W���w*ꖟ���DݗS�}�¥�Ֆv��K���$:�a;MYs%NdYyb�!Sz�\��O���-5����ۛ#^(��ؖ0!D��R���*����ӷfV�+�E����yn�\�l�l53{܏���Wm�Ҏ��=�%�[���������z/zt�TP�izLd�"��"��X�.�XE�β,�B~�=`�r:�"����֎��B�~�Cpu�^�R���/��J��b6��BnW��K3X?sk�p��T��}q��Ӟ�x�N�Oo��R�y��+����R~;�o̬�0D��ta��=���?̻���u��'�6�Y��:��b�3�y��u��)�vM]�j����	�ꞈ�w��X�'���R\ߵ��}�W5PR��.YC��5>��P�+Ҳ���폼}j+-�-���N��J��}B��~dj>8{��C�`���3��de�'3-j6Q�r�Y�-i�c����ms��O��?s(�㙞�`�jp���	e�'
�G�&�6��0�z�,��?x�>���w��V2�W��AV=�$������QV��hv�h����-����l=�O(�Dff,��d�B"oo옙�`w���9������gP���\�����٭��=�s#I["c���o��-���	�����BםO������{C��+ĿlUq+��sd�f)s�����q�)�Ò��`R����+��<<�z�T{"���2�׳�鲢QM�M+L�%1W7�E�;A<�i�
`]9rx<���kdW�3�Oyuc­��Q�;����7쒯ޮ�M�j�5�[��m��i�4R(���z���^�o˥��vv�	i�pX���y/�����}m�(ǴB���W�T��$N�0��Tؘ'h�K�U���Gq��C(�72ڎ�U�4����XV�O*�<�q`��@+mz �ޅt��R���)y
��S�;�iz��$c6;�ҵ�z�(n6z�>��\�w�|t�e2����BU���zv�5�YL�2�Q��	������^r��d5�{B�����C��x�W�-g>=y�Y�O[q��z�{Mv>X=�7=V���+�>���x�L��˺$���uV��ݴ�q�5�݄��a�KZ/�
��o��� �\�{j]z�C*�;�d�>=ٿ0��i�`���b�H$�J��wD�0��4�%���C��O�SbƔ�x�Y��v�+#[֜���#n�;�%��vsZe����|o�!1VW�L�G���v���U�Q�ݟij5�ϰ���{�kJm m^��6���P:x��:�J�,J	���(��'h�}�C�����G,{��� �a����<�����z��+���b)Y@&�.S|1�RC�Ŝ]^��{I�*����e9�R��mr��S�|&q�������{9Rn�~�O�"k�����l6�h�^�a���jK���g�wqrke T��H��)l�ے�f�����έ����������^�� U�d�G�uZ�>W�]9�P�(�&�eQXb4Å�]��ȭl�nZ�f�VjU�ɮ�}�)ĤW������9N�����d�-%��f��H,���+z/x�������OZ�U��pq�U��r�Q���&����L3Pe ��sϪ1��o%�p��kۤ�zU,�OQx��^�)��R��5Qde�3�V�͋Ƽ��՛��;U�xK�m��B-a��*��R<�`2�[J��[]��ڔ�:��|�C0�/S_n}��D�=6K�+��ڐ�]<�{9���c{�r>��
�<F����H�)W^�^���jڿ; U���4��bh����*�Vte!�oؒf��6��AX!6��W�5,��9���:,��@�&d6��rCJT�e��V����s>��L��ѕ �}\Բ��0u��-��㾛S �,v�JsxS���
>��J��g9b����߬Y�Bm�����f�3@P6��u:Q�.�$�<�;���C4�rcz�X{h�-Ö�Y�����z�]�5S�ib-76��ׁ�0�!l�����P�)��R+0�4e3�
 pa�WR+1m'ȹ��<l[	QϘ��ŵY�aw���e�r�寽2Qf�{��s���z��۞�(�I�]\��eY��s6�U����Qsɍw_x�6�L��dV�b�DChq�$a *R܏��@���l����J#q����,�/�Ƕ��v.�껍��E�	����yD*}���Q��=���F���,i���F�E�ԯ.��Ґ�4c�|��I��d!�P����ñ�rI���
{���G��1��4�o2�S�I��d�+GݳZw��`��M��8A��ŧظ��.'gd����#n�6d<�*�?d�\��׫$�k���ب��mJ�����X�|V�M����CKr�iGf�^��K�6_cP��겘T�۱Lve�����@�]�3�8���]�,+��(V��.�D�*΄*�mI���j����8��r����;�Q��bu�{sP��|��,iʛGe��B�����]��߀pѥ��s-���������#�/Wb�V��/0��6ELm:�7Q��8E�����Y�;�wYj�l�${��7��z�F䒮�{2_����Ɩ�(��T\b濒�ľ1�93��)�0y�RAMk}M�\�R��k�W�;�f.(n܇���:2����Y�(�3�R˥zx�m���Ox^^H|�E��������}�5�������3Ӌ	��c�X:S����o R�h�T���gxc���,���7pk{B��tZPV+�Sx�a����7�]C(3A
�7]Vj�$4�je��̹���ྫ���*�TE����>y��wjTda#1qp\{��h��[����;�Fmw#Pު��J�$�u�!Fkj\�n����j�h��Uj�#�R�t���S=�Yޭ �h{�孾 "\�6�`g\�[�l'�P��I��\;�){A�f:9��%��_^��k�U3��˭�]u|��	���2��hq1	�L(�Ҡ��G�f;��`�1H���b���mC��b�q�꽰nf���W�7�]pd���q�AL���f�_j�oE}''�4{���P�
��r�5#���|�fvS((�S�^����rg$�(����U<��(kU�&fW*�M*��Њ	��)�D$�v{�Qp����]�Ǘ��2�eE9H���<�W���I/r��x@�.EE�I�
��0"���L�C�l"�K5�$BQI+^'E8���r����	��'+�FU�E^$��9fm0��N�94���O��p]"�e��)�7<�:�4�L	LN�k,&x�"�<�Ǐ1	�s�Pγ0�kv��8s�����.+y��\����.�K�M5V&yq�Rdz�\�!ȥ�\����bi+!:IJr"�d�ʄ�Sۜ�rʊ�<�3�\�E7)M<�
/9'!(���N$�4�F��x��ﯞ���_>o8w0��������W��Ǉ�o�F��I���-�hbr� ~�`ˢaӓ��^V�j*-�iW�p��[��Y���d���oiE�*v�H3���½�|�r23F�@A-�E��N���-!�[����~�&z���M{��+kӽ���ג��ԶA�Q�2�6&��O}G��k7��x�4��8�^q��_r�R�h;<��Z�� T/TfcǇ��(�6����w���3�j�&+��0|��� ���}O�lt�g�/���u-[��ay�^�y��D�&�E�<X����
��r�8���O}�v�W���0-P���2����.%�>5/�5�lC�z��ӥz"�ު>8���C�`��lCL��<�y��>�}7D�mF�%@��3�J��'�����B��>�܃�M�����լ�#IH@�3�Rߕªc������T03����X����I�#p̌�/|4�Egڜ�u���_2�Gm�-�l$�ey�z��lbd�÷�ċAVY�fJe�q</>����w�*����ݩ�/O5�h�(����de�r藟j��M �uφ;�@j|R���]Q��W��)f��jo�$R������F���� �9�\���R�.I�b�k�������&�VT+�^�x$kƊa�%�lUC�>��[2+��5.VmJq�lë1d�iR�@�3Xm)�8	h�(ŝ.�ik���yLaQɫI�ط|+�۞Vxt�����8�8���Ɨ�ή!��t�Ol�zF�}$!a6��
�͔ک�u�dkN%���D�^x���ԋ��}~����M�Ҹ߆����y�輩Z`�g��vD�i��3�:O�)��>�h�Uy!pi~�$�b�)�l`8h���z5�@���?)#��Ŝ�t�;�����9�a�O��6Û��pA;r�*���ĊƲ�*����*an<*���-V��qS��.��5�z��x��}����.i�L���A[�7���Xgd�Uږ��gޱ���\������'^�&:���5�-56"���T6|�]���n[����w�8��P��9���E��T�\��e&(�J�qnr��I���R7�y�gZ�[, ����&�q��i�X.K�YwV�oj�20]�b��/"
7 Tf�6oo�e��W�'s�c8sxu������c��;pkK�geqX�����W�Ja�$�c{SS{.�]����?���ҽ�y�1#i���ԣ\�W7������o���m����%��������4��5�FQ��R��Zg��~��Z�9=����C��q�1tO���lVÿӆwԛL�vV�RԵ,�b���6H�eG|�8�?}���H���d�%��h��H�P�>��W�k���iF��`�y���d�UE3��iKdۦ;��5��Acx�L=�+K��&ж.���������M����r�1nS�|%4�\�,L�����@Ƚ ���MZћ"mn�$��J�lU��V��D�2���X�T�L�}��I�S���U����xVO6�)����0/����JL�nO9~(��tν�(��-�K����H�k�)�+s*��"�QM^��o���=��������H��ZhӥP��dw�R/b ��"����&���~�"V�u��V��o��B.e�Y������	@�V6�9��^�H��{dZˈ�<�����$i�(wÆ�hC��"~W2�]曻%@?O�c�{r뼕���
8"º��N��J7r����ԞQg��ꥅ��*��S���:�
��!D߷��0�b1b[�Ӟ���k���.������?z��
��uf�z��j�����c�D�ޮ���F�Ž{s~/o��]T�Z�M]����O
�5�'+�U�̹G�P��Z��y�V�������������G���YXAA��9�ז���M�q���t��g�u)Y�>��ߏ��}�V 8я3�`���.
��v�������0�<��2���r2����F6���XJ��vedE�^�&[Nݪ	T���mVô4�|e9,.��\�;O{�N��{յ���^w�� ���Л�M&ح��3��t,�oD���x����M�Vװ>|J��"��*}�*�W���^5OD�GYSX��e� #�/y�z��ms���-O^W槼]d�{u�����L��Y�Ehű>��OS�^@@��wWX�մ��S��U�6wy�̭��5K��&������]8ѻ*�h:YZk5�҈q�h���F-��<��&ĭk8�����%&pbL۱x��4��
��='z��)��͑�g�qE��1��>��fJ`eH��3P����4�1�[�cb�W��}I�#Zf��GkJ�V��
"�*vJ�F��Ty����{|����dou9$+��gIt�px�;��z�{}��:�S�n���@3ū�½ٻ����{m=�3T��m��sI��
�thhP�gn�t���|D���v<���vȵ9�m�Dd�����R��P���X�W����Ѹ��;������}���ɽE��f���=����L����X1J�2t��/õq�;�yGo��g9�	\"����W���u�S-r)����H�YK6M���wk����gx�gP>\��3��x��Vw��R�ZX&�W&s���3^����c�l0uP��:x�,R�K޵/CO����}���嘣x�{��'zx����G���V���V�îV��>J�D���h��y�@u�טtz������k�n�m&��V�텭�L:`�쬹aݬһR!֭�r��������W���E�wB��^	叺�Y,,���]$��x���9�
��NQ�sM
��=O���5?/l�Q��(�����w�^�,�֬d�%��~W�ʩ��x�w��ף�#\�?Q����*�'���x4�q��7'K�u����{Џb�w���^�t{�P���g�"���>:���ݻ��d�6��p�KH��2�Zh�$���1}8��2u�,�G8��ԯ��oOZ3�)5�s������>0X�3E4д��kH�1��[,��jׅ=;�ݶ�8�wI��6V�������GoӽD�l%��K=�Km���(�ow��=�*�e�}a���+�*f,�&ݘ:��IY��I{�dW�\�����wR��f��u�#]c�����R)�բ�_�~f�ʆ��T��:�e��2ԩ�N���ԟC	�@f��[�Ps���5��O+�s���YY�f�S��9&���`�hO�F��~�9��s���D}�wV�xs	��U����ɣ'�#���zP��h����1��6e�[���r�k��I��t�1`��D�w$g���OY�"^+�we�@�`�e��V������oAeG�պEt���x�w�!�O��X�ٜ��7?W��1����U��{V�"���H���s~0�yBփ.��FM�,O39YKH��v�u�3Xar��hF�1M0�)�J��Uٚ�!�f�</�@Y*���J�,�i�L��}�I�%��T�i�|�����P��j�X��l5��w9���gcj���|�O�3��`�׊������s�P��ҩzU�f-���힓�P��J��ҹ�R�)���T|p�50�!��C݋id��
�K�v���hi�C˸�&FB����4���Q����UYR��'(�*
"�{�ͱ����>ΪYT~�+�V;����<������uH"���QVΩ�[Z++��P�8g����5�_���0�yF�su��"�OmdC�O�[��V�ϵ:�t�e� ����)�y�#,z�0�����^c��+�,�i*}�r����4-*Fߗ�֝*��)��ZA��s}�B8L#��m<�����0{*	d��څO2�� kߩw�������{�Zx�~�B(~/h�������M��cܦ���%.us]t���&��}v���=B�V<�)o�l����Z	��v�T��G��+�֖�\ݢ�'ᥡ�QQMgbU�EL���6���]����v�_ӫZ(�^/H��i�[T�US5����B�ҳ\�{��Ŭ�m�wtJ��!��jk���Õ 9ŵ�;wNT{s��J-h��nz{ܱFt��X�ǫ�:�"�X��G�^F8���*팝gl�AP(�+7t�zՠ��
��S!e
�6�,�1�P��5��2�YMv�'l0�t/T@�6�'H�ژ��W����iL��l��h)\�rY���d�����3l�|����2�m�_(�s��Jg����
�+���_V�g�Nu�NӥF��^�<�P%���u/+ͪ2����y��OZ��k�N�O|+~�����!0z��c�m��|:��3�;�+*�����}E����c��y<�%�@؆zH}�{�0u,y�2����ׁz�)�֡�u쬅i�/iھ��E�3U	�[��	��{w�^�c�	�N�C.������ ��h���9���<�c�Pr�B�]^1+W�z��M�}��m�}�l�4=�����Q.�Os���u�#!��������-�9W�m���ǃ�X���i6�l;CLu����d ǝ����<����%r�
�-�i:q_�^K1Tr�`�7nM�v+E+ެ�=��To��ps��=G�P:q��>%T�G-�-�l9j�m5��`�9�����9�++f�a	4I�?����l�z��T��S�����?=}�:�ơnd*�t�QgP�+y�MF=�����ب��.��#�:�fE
*ͣ���M�4ְ���T
�KD�J���*��f�P"U�s�K/')3�f$ӌ�LKj�
�16���3�����Z;�rca^�6QH�%���0��l{ԧ|<.���^��.�.�Z�8����fd���_��� <� =pj�vA�H/(�+^��(i���NC&D��9uOF�O|���ޣ<�N4��{uI�1	�ыe,�F�B��D��͵[C \N����/*q6��+}��xy�H%���ZD��+3q���������`z�����
+�HkI����wu'w^�$vR�f7�t�$�STRT�ݲ`�f�e֥9.�cU�R��V&�W�,nt(I9���aI���T�.Z��ǚ�	����^����y�ݱ	@ҷ(�n�
Hg3����6�>�^;MvN�`�SsՏ�^��Ã�6�03S��R0!��[G((�r����2�k'8���fU���{�_��<�\|)��f�T��T���v�W�ٳ8���:x�,��lL���)����A�c�;�̌Zj��>+s!K��$2��5B��b�/��U�V=n��+�Z�5�t��uRjJ�d�ƵazE{lၚ��=�M���?B��B�Z�Z�
�Ni!+Ď�ެ��3_�]�]Y��r,�}CY�gh>��dQ�����G���m^�7��2'h���v[�	�dS�N�P���OW�ݮ��q�k ���uE�����qw�'���P�j������k ��F���IA�ck4�י��:ܦXrTRTϴ	�L�Z![�rJ?}�J�@��ȫ��z���&��s�6$,�U�ς[0�4n(VC�(aݚq�l�v}IT��4u���t-v�ʜ�Ul��MX��R#6�
i\)�̣Zk�}4eeqq�]J�`���$xX�C��kJʃC�{����B�U�X�ӽ@2�wx�u����ǯ�� }Vԅ!Ք(�%'��53	@3�y��<�h�i֞���6�U�#����°j-�� n�2�ct�^��P^���mE�AXSC��Πk�U�uطN����_aWo�:�.z�OM	 pee���e�9N���G�w�C�axNþ�8�l�������=S��Ho�^�r�=�i�g�������3]��As�;z�<����V9r��>_'�D0�)[U�w*t��&a�5�z"�ac������G_�v�;QZ���Y}�GrcRM]h����啜ARiW|�x������v}��m>B�A��� r�}�"\�X��ɑ��oA3�]�ohf�5�����X��(XG0�D��oi�{�Ct#7�����|&0������\�¯��X����յL�*v�fu�&*z�(g$�7|�G��&b�m��ךȭ�=s ѷ���|�VOɇ��1��;��xthL�J��ցu�1�ņ�ѡmF^L"�:��M��Q��l����V1�@oa8�666^.-��]oh���u-���1q�9B�K6����X����Fu6��/qMv��f�2.���ݧ���i��՛�:o��DF�ٯz�jnĄA��h�DJU	cV}��� egѴ�:�YF�j����@�=����0qg}��L-Vc����8u�t��EΆ���S��'�e'�x���6��ơM��^��<�eX^�I��,�𭽯|�s���LA��l4g�I^��
�2�;"�ToLԜ�:��t+�mY�[W4y�(���z��g(����m�S5�o4���5�Nq�n:��o�������-�j��fM\�͖�j��5j>�:�KE��DRY)tA>�t�Zͮ@u��� O��ٷWyh,���9C��B��x�����I�X�-�r�OX���a��!���V�M"���;U3N�. V텉v�j��n(��s"䋋L�	�O��yuʚ:����D㬀/��8M�Y)��ec�Gw�E�����j+�g8��g���ɜ��֋�R���*�&��;�VF���6!����^^���470y�F:�b{��z1ƄY��ظ��MK+�����M��SK�x�>��d��x)-�H�q\ 7a�'n�^(Ô�QI��Dy��_uG[�c;�y�G�p�m��k�������
$P�w�ol�=ܮ����.XO2�<|OeЧ�5F]��;bՎ��a/�A��|�F8 ծ��s
9���X^��Y֍c�+,_�w]ƍ���6h[%��֬�3;�v����^���1����u���5e(��|���Fa'����s�T��pQEN!�-:;C�P����U�U"+R�(�����#/.'%�����r�mnS�\,T��+��;D�w)N0���G4����9ǃs�<�;3ۈ�[���$Ve�w�ySCv��rȪ�#�&ʼ�ïx�r
$l���dUP��W$D�8H�x�*㎐jc�8�9N�U�V��D^C*�np�^G���2��w�v�宼8!D��pX���*<�p��8s�
��Nw�x��(�E�U��K"�BZJ�L�F�XJk�\ꪨl� ��jX-y�<�������<�dQ|�r���U�KY�����Q�9�i�r�l��Q	��UA�s��Ѳ�XyKZV��*B3J��R'�T�)�%|���9�[�|  ���9��Ggh�sW:j�
u0� ��:�z�ũ�����Oy$Y܉���L
76���ί�;������u��������5��O�>#K�I4��ؚv�fEc��bs���N������z�H����S��1<��}Jw���ɬ�]w��uVpS�^�W5��E�e��w�����,Fe�������F�Z�#��wQ��ץ�㧶���$`�`��[��Ʃ~Q�;�	c��rE`\7m�X<�٤7rPy�YD���]e�i�}��һ�@޹�0%.c��E1�y�c��r�X:EhX-*	2i\U
��sT髛P�M�U;����CeߕG@S��t	�W�}q�"[N���h�]E��=*���w�؈�B���cM�dt5b摢��q����P��  �_�鏸m�l���Ջ�����Y.ZF0�=9�LPθ/8+ٰ\D��3]mϪ/��:�Lx�<t��]�X�9��=�csڭµD�}-�W=�=z�'3gC�u0�N��&�w�=������96��:����c�/�<���y_��|��ۇ]7^���K��Y�zV�?�W��9�w��_�\^ɋ�5x���gU�wL2||f��n���YO\i�0�6���7������I���h��=T��i+����v���yYm:�m9[�=^��2����4��i,�76ң�|4�P��cojU��sHE-��b�g��c�SL��-P�iX�k���#wvb3K���{+�/��5����\��ڴIz�f<���|-�'�f�Tʮ#:+�9��M�	��x������땆�/;P�	�Hsr�I���0A�-�yT�mӃm3n�[�ʮ �m��t�
x��nn��V������+��B��Ʈ�"��l�dh k��P�&]��L۸R�P͈�Wg&GI����/^��ïڦ�W�fQ�ȿJ�m���
��g70�,M
D�w[�qk��7�bSf��\a�}��ߛ%9��~}�ʓߛ��#oݲ0K.���y�M�;.^��na[ě�Qͽ��b���m�f�`���":��,��.�z]�Q�Z�]<pFh;��BZ��/�q�w׻��~0��SX����l_�Cǂ���z��ˇF��FL��M��/c�@mb0w�C�;�F��p�����z�(<�+�R�?����܇���-�.����/�ձ�r3��+5=9�K�m1�U����+�=���.����Ί�s���]��U'a�6�����O\~��5��a���c��a]/�/У��
�ynW= Ⱥ��7\�mǴ��E�םq�5��x���l�َu����۩ud��A���N��6f���D��B{.�6ƨ�G)m�eLי����D:��ܞf���떲��)��T����~��WY���IN���re�q/?3z�f�E�չ�B�V���:1�d'�c|�/��WK�	���)���_^�KuE�X�{�f�X�Hu�n��F�v׮su5���m��>�N��=<��fBX���������:���3}n����̦AQ���_l��^L���l�w�4�ކ	�ga���h�����5I���ܨ~.)��c#!=��S���f���'�d:�S?\�,�l�GOK:�ES�֩�6s��H�Fi�~�4J����n�<x]7����b��7}��V�9�����M��EI�~e�S<J�Apθ��[n�(_�X	
e*q���;1-��p;�M^՝'�܋#��3E\A![lC�L�=�߹G��x�hVi���j81��INy���woY����o���LFY����MoO"�\Bsڦ�>�]X�۱�m���ܜ���S{��U�7�a�}��ѯ��M������Ck=�R�yj0x)��dD�vK*r��U5�5-����˫�\%�P�n�w��=<�L ��:Q^n�N��~�a)g��w/d� Tq{c����Up8;1��x��sw�1ީ�ܺO�ZeqF� �,��3x�_0o9q�4�씻s���B�ԻFQ��Skf:m�[�ŝ�T���θ&op��J��Q[����ndSW��Yu�η�8BHAx��p*
������T��<)}�x��M��U�1�E=�\1�cz�T�.��;�,0�2 z;EGb��m�b��؇���'��E��$&�e�3)����}
���<��R�G!M��]oLG3�Da�흡ѓ(�*w�;�{f
�q�{ѯڦv�5��=:�e�<��zC�o�;C��G��"�kS�ׂ��n��N ��&rFp���<'�95=�B�GK��"�Էe���e���-�r��[w�îb�3�Y��ޅ$����쫜�ʯ�`N���g�|e�<�3�Vv��-B�lጽӛ�*Ӻ\�����Dh���<�lE?`�̖U����h-�˂�[��E�ٲ�5�f�9?{vd����wL�����C��Ekt�s���!=�_N:��q��!�ӿp��[Y��'��N]���J'8;�(;.���X�@e�n���M)�Ov���hh2��4j��v��'���
��5ӽ���zk���g�wJ"����VvThnV�Kݝ�*(����IHq��#�G�l~��,v*������l��U�'w�)W9�8�^]t_glj��[�x~�f�v���+�
>=�!4�.���a��`{���9x/���.�*��t���e���ݨ��D��lfY�m���+{��:��)����]�B���Y���[T~�}�6����<��q��6�fТ�lp�� ׋�,n�<������u2K^��?F���u���e�����q�\G9W�t�L�W`��U�	����wa�k���by�{2�]=�/�ƈ#LźQq-n�ӽL��)�!9�m�W,�}�B_6����nh�J�$$�WW9ze6i=����6�t��^Q)�l_�[�y�*g����e����"���q�Y�L�=H���i��D�A�˶x�n�ꗚ�4��8w(Ktl��s0�V�>��~��Ց'8�$��wB�f��ds���uIu$ۋ�(v�cz�S+~��	�!�!ǟ]f�=�	��ܱ�w[��t�=�F�6��E�9�lk�dj����$(��W
������p�	��k�.��I�#���N��`�m4΀�+g�X��xO�cts�2��B��'���Q��*�e��;�'+��sg]�~�1,��ZQ�����43J����xebO<s�n��!"H��3�h�Uv���*����wuM�]��&���C��Ϛpxm�2=?,G+��gŗ0�r�u�ㄞ�����Om�m����4(Q�~"�L���r�ܧ�WmQ<�p��ց\��{t��}�|�!g���XN6�5����LguD9�������5�����4�Pu��Wm�p��{8�
�C3<%�5�I��m����.�x-���f�e��PS��/mЗ[�M�z��͸�`���l���*�f\�9�f6|�q��l⒫4���_���gr�miNI߮}��DK`.L̲�:�ع�h��~<.v��A`��0t������/�I;�*��V�K�m���q�81�7%;ǉ����9��m�(�vļ.��
9���wDw)�>�H79�s��Tb��%�׮N���Ȝ���6Y�A����;׳��FZ�:\����A��������-�8����3�.����][�^���+<��Mh~/} �Brbv�����Muv/׊'�N������`���2B~�|.B|�5L��3��c��ȵ�T#Q��[��U:EJ��¤p[��-�'�U����e��>�Nǁ���}7��-˹]$��H~�w$1��8�n�b5��|�g�[wB������-x�� m��<�L�T����
�x�P�<��9�f�joH�u�0��/^���[j�uL��{���:-����J�[��vaӯ}x��&�w�y�2]�o�0� �t`�S�����~{n�)��tm���'���̫�S��ULk-ڳ\�C��n�`���ζ�f�ZI�l#�!�-S��)�$}�
�ޢt�:6���~���+h�B�n�[�.�>6�&��bۃ ���h�)�1%@���XM;�G�,W��TI��b�\{w^����hLW�E��i{"�.i��@}�aS��X��ONsF�c�u�]�#D,U�.�`�,�hz��wm�=�E6�������|��^Z��C�.��e��ȇr�-�C���1�Df[�.��̵4�<�\�ף������;��5��Վ���A��)��u��xm��x��)o�X����탷���$�b^��L�^1�@�Y.��t�*�zC�A�tF�t�s���Dh���ڂ��en���U�����͛F�3��rD���=�l�K��fA?O�
�y�s���y���~�S��W���"�*Ye\���`kb�q	�H	���51].6)�D�w'�"jFU;��csVi0S;�����0HѰݕa�\v�Ѯ#!;���O=f����{�����{��{��n�Hb8��Ѝ�x�V�������xfx��G���R?umf�L�M�}"�'~'�{�)�ۙR���'��њ��!� ����r�׮8�]這�K��UЍ���[�Lw�B|�-4�4��)����-zǲ����8�pve=����5�߲�ve]g5��l�<tW2����>��L�[<Ғ����ul[�PE2��2�E��@C?3KG#,*Nߋ�lbo�<��0�lJ�kqX�ƺ��gQ������ki�tV��7D��sOM��E����v����o��1 ��+�mO������Y<�{z�ꥎ(B-&l�ϧu��y)f-y���2ѥq�OmnV�����T���~A?�x�E���^��>��q
�b*�]����ʅ�}��p�g���҆��l��l�xXj��D_�W�3���!�Z�
����	�j�Ǿ׎#B�k�����n��L�1�ny�n��uC��}���)�Bw[q-l�Ҕ�Ϩ���Y5�,���׌�2�O35s�"��e]b����q������,�T����!�a*g��Z;����̮9O�����&���Coy�U-�@ ���ߪT˺]=c�t��4jm1q�S���&#z�yfI�����x9	̆K�v����3@"ۗK���6��!@w��M<�(�Ή�֡��Q���VmL��(G��sL��cPǰ���t��m�����P֣'�"��k���㣦"�233Ţ2�!a���!ߚ1��m����d���C�3|��� ���5GK�Fߓe�lF�c�(���������[7�3ю#b�����{o��p{��V���t�:�M�V�N��4_�&]ɰ�_8!PL5��:�_�c^d��k��3O���Џz�/�K�m��bI.������K9]�X����
�鯯�R�".Ѹ���dUt35�����<_�j��/u�w��J�5޶�T�Z6��v�G����YqM��(e8t;ݭu㌩�л0Sw���q�	�<�X�q鎒��9����i��#�ꊛ�_�TN���S�w�#��U��vh�9Ɖ�O���i鸼.��C�挄�Wӎ�c�-�T��j���m˛ӫ%G2��k�y2��y������^�ne4חeF
�61��5	ʈ�b��F���fu�3��q<6��������ʶyf�=}��7�}���7�Q��`�>�e�2�n�I:] P��%��`�ˈ������?e5�'w�5����\����:J��{�������푑�k���1�!}1��n��jS���\G9W�t�L�W`����7�ߪ���c��"�A}�+->�vl�6�^T(�F�K[��K*pP7��X��OC�VPV��N�ݨYS�Q��;�
n�����l�;��C5�HyU����=;�Rϱ�wt�Uvrx��՝{q���],�T���t_l-���AɄ��t�7B�u���I�g����V\\�&��6K����d'3��������ṵ�g�{�Tź�H缫���k)�N�t
'5�H놌u��0�-��`����2ճ��L����$(��wղ�(��v�j�M=��6�y}�����7jt�����[��t���慎4f��Y]oaT�0r�bV݋t�~�Ѽ)�C;�5h�@�]J�+R냱@�a��V��Vk�d�V"�&Wd�dС�Ӗ4@9C;��b�2�+�mD	̴�����y��F����,Cv���Ѯ��f�h����l#1�~�����W����|�G	�ȻZ�����g��u^n4���S�L�捗J8~���%l�l��T M_2XЬWu�j']��~��Z8(w�>Q8�滲��]uK�4~�M8<3-ퟞ"Z���Ǹ
��F�v a����29���B[��NP������3�����V�@SMQ<�@��u͘ �Oaמ���w^j�����Ҟ'!>����ƪ�W�̎����#EwL����;�b0���L���N_��fs^�,��΍�ӯ�q�:��pW���FBw�&���ζ{�:����<)e������H>d�'O
�E���ZM-�Mo��	x��@g��)�x�>����@I�m�n���{�P����N�<�{	Ǧ�;���0�2�Qp�Z�v�b�|[�����rk�"4e+�_H��~<�bu�uk���>���E�.^��C���Tʼ��8ue5kr�U=��s��H��|��]�8.7]6h�Jq�|��4�]�S(�r�ߦmܳ6o5�K-�˘�@D E��a�K���a�]_�M<�뺧;e�_J�[����<	Fm�j/eQ<�9��_�lǨ=6��v5�A*gv�
�`oϒ�]�a��*�|en.�>�n>�x$}rM�w���اJ�'Q�m>;���2*��O�V���y༮_=�`�[x(gAClc|���=ql�Rw�1!<�NVȽ��#IV��E\��v��o���t�C�b���0еt(N�<ۀR1�n�9��n����!&o�П������3��{�e6f�מyIki�&T˃޷ �J}ڷܒ!��EJ�UƉ����z��>S0+��V��R;�CK0�t��gk���:��H`TS~�˽^���B
	�T-�Y!g�ܵ��I-|�94��C��}��@T����f�����g�fo*7��3K;�yr=���7���M��ی���\7�b����޻���溺�QT�5q{^_)�n+��5�4��R�EV�^$9�k�9�^v�n�a�%k��5{+KW�,��fP�s11AոL�!
2L���y��7�3�5��N�ް�p�*���:l=\
X��%�ݵ���"NCj��\چi Ӥ��1	9Д������᷎������Q�,�[hl�#k������Ġ�.]C��\���-����-�H�_^�/ 6.�{7�w�J���K��u�Hep�������送}��V��A|�FTYq�>T"����5�6y-[�yN�$�(ր��4U������ųxh��y�*�8�&��0�x��D����ܫV^���H�������!�1���<>�v�E�3�m������[�Fi��[v93�Eh�4�H[�m�B��}&JF��Ev�gs7x*Z��?Ӎ�G�����`��(m�J-�/�]�{<e�X+OK�?]��{�R�+�%r�]]�hԝK�+}/a�*�tLQ�U�ڈ�
l�hx�7������ء�gezݨ�b��h�;�(�p[�[GY�¬n�˦�v��������3V�����N��"N��걎�%�c��i�{Q�6�}H�����=Be�|+�eFJ�W�^r�[İQ��ڑb�@�qk*���w�:����,�2c�[���*��[�̥}�$ ��%쵽�6�@*�B�]7���U������o
Cwћ�ﴆf[�*$O�ցt8 �z�W֬ힾ��OOj��p(��j�	ػvۑ�J�r��+>�+t��@&�-�:�������
5��Z�0:Vf�B���/5X^�z�J�ң����h�#��*3�rD�mv�\l��hvQy7qZ�������4`��9� �*T��;��Sb%�vH��P{wdQ�l���]lA�|�V���,�I4*��Z��Cz
��zٷR�^��bQm�,η+#��h@(�xb�=��]O턲��]�[�d�!Q`��{ژ��cwI�j��^��M�Ay��+�GY�V�5�Y:���f��T�"����m�R�PزM�.EZ�:[9��#-�!
av�f������AV�8�Ĳ��`�uS�ZG.#�p�ӖFi�EpԚn�^2.PY�Uw���F��S�8s����c)�F৔���*�f\11��ZWeJ;��Fr����)#�i+X�fjʪ,� CL�.��,�"KUi��fq���J��-*
��Ҡ�FJ��\��L�r�m��g1q�N�󋗃D4htU2)F�V��f��Y&DWe(�̩R�QE2�E��Iz�.
)+㸮㨌��q9�Nr�I+��FN���JT�\N˲��NP��21���2�$$��u�=�!�*RL���q+*(BW�.U�h�*�3�tX4*��f�۔��Τ�&�9]Q����Pݏ�7f��p�۵���B�����a>\���/�f��7��wM@k\=���-��,�w��BP����p��pH�W�S,�M��CNgPz"��������f��݌�ry��Aw��?T"9��z��S3�"1��_��]��
����+�X��|}�kz�F���i������{������
r���~~\�?k��pe������{�<nM�胝�<��!`k:[�{yh=&��G^C"}S�ͪ�DL�p%����p�����ͧd��n��]*a�˧��c��"�ع��x�tE�,9��`��"�ꓓ�;7e�q�k�0��t�}����@y�T�ߘ0�LӲl�vK�u|89��ݎA�v?�x�%��:���mR��B�w5�t�,���=4wDlVtF�5�)��K^�"�^�iFn�:�fHu-PpC����t�X��)&xT5�O�1�c?K2.�)Y��7Tfnq�<�\���3�*Yez��\p�^y`)�c���'��1�T��~`�U�����n�ɪ��ܐktv���,��m�h��l�mz�02�^Oh���-�����-�_�!
<��:�!��&b��M��>k���7k�ٜ8�3��5�zQ�<ļ+�}*ވ,�6��!�/��ܱ���'�؊͛���7��ӹ*թ�'�|egKU��$.���bU�
ٵ�6��,0wI�g%>�ЈW�zo�1�E�X�&w:�."�ܾenӐG�Ҁ�ª�du\S縼]2�h�eb��YS^L�l���_D�K)~�s��uCmaS��n�]ߛ.�;�q�A鳧�h�|��8�ܲF���x+ѐ���)���Z �H��ufk6������T��57�g;���Te�}��)��5�rq�j��bfy��NzT��R���{H�3�#6�:�V�~�d[=b���-	e�i��L���V�ܛB{Z#u�N:�o:@����:"��H�1
�$��S>�p��Q�b�t�O��-�Q�fg0�m�:	'h�2�[C�Z�(W�Ő��m�F��m]9㲬'�����2S��>���m���!���ϵK��l*e~��Q	�m��Z��)w�0x)�dB�`����w��{ϦJ���v�h><�uus�90����StBw��{�������qsM3wV3{�4]�Gz�NsnC/D2�2�$R��Ѩ.ank�� �u8wD&l����`�
�K3.M:�y�z\��2J�\ث�5n�*e;]�ۢ3@"ۺB���̮eHwL�TݴM�B�y�0�1{]�jƎ�g�{á��p��|�-�y�t\��Ζt�ٺ1��gc���[�֢��pқM�3�Εl�Z��7u,.U¥L�V��.�r���}���q�{E��W!���n��(�U���z�+�C,��E+���j���6I�C�:�
������)5Ȏ��o:9�ة��.q���I�ֲ���a�e)�n7�����9�m�=όH	���ؔT4��ux����
�|Q����L�<��3��6�*Yez�02����Ml����pR`������Z��^Ы��UO��)�G7.�x4�a�
���w�w0D�L�O�+י,��{G^Z���{s��.8���`A��j��a����3����P�qx]{�C�ѐ��0ވJ�3��{�N�s�T�
l�b5ӾQ����Q9��`�h>]�M�dX��toB��ѱ�Vr�:r����Zv��GN=������y��=�n���*���g���ۺsEy�o��]�e�3u�ry����A՛g�Cs_c�辘0��{���	�#8S6(w�Cf_��e;�4�k�NO6�ښ`mM^�����.z7n��=�h�ז��
�1�Y�OMq�5�s�~هO���I�V�㉬��t��}��U��̗O!�]<��|{]�K�[/*)�źQ'V�ν�ew��"i�eZ���`��p�?�$�v�)�Ώ�[�c�����3�W�آ�Su�\u�*|��jk�[t;.���&Ii{���=J'�;n����LsdG?	�����c�����0/L�Iev2h�{�;��r�dq4D�].��pѧ�)��h7Y�A7=o�9���s��h<�u'�Sf����6�PzW��dT�w��9P�Y�Of�q�S�'c]F������h���)���ʟT�-���t[v��Q���`��
�C�A�Ylh<b��6�B��~$f�s�.�����w�j�Ð�f�Nf�q�2]I�AI�ͣpKuҦW��,�0�:���{�#����VCAu����!A�w�s[�T��.� �3*ZЧy�������g��vm���;!3d4[@5�J���#������φ@dlȭ�V�gQѣ�Gx�Iq֗Yw�ʦ��+��g�2��tC�`�o���+���Mw��U��xFS	�y׮؞t;�i��w4˲���_T;�4~/�N�/2C�沘4�)�ꋉh<0� su�͢��	c/Ӈ�P+�ߴ�3���\�ϛ��B����s��U������ʌ�çs��oN:���"}��	������+�������B��g�ήE�u�9�fa<�f��p�|?��w���6^<�ְ<3<�����.��������oJ!Elȃ%�n}j��d��#j��{��Պ���0n,���{��G�ݚ����5�;���]]�CD@߽�����OWM{V��RMyV��.��k9�J�}�E�4*q_AN�K����\V!�ҧ��^.ݛׄZt��[jw#�Ô��wX����g3vDi&o����pj<����#*2Y]z�'�c�C�u6�w��H;�wn�&]�������R\U-w�����6�����\��t_LoޙebnrYU��
�������8���3E�[;�g�Ӯ���4zo��2��4Ǯ���oh���2B��C���j�����̦LsLYxZ��;�#t�i��@��{�#��3z�]M�R�UϤ4��w�F&�8.��YS�\UX���W�yĬw4e���8�U��C�g�=���pDetq
�6[#��`,�R6��k�N�'s��wݶ��x���!>�\BC�Īǚ�̢1�ɺ]�Q��NƜJ-�vΣ�g�'�9U���GH���t��a�}�w�0x)�d�3]8���\�=F1z�WB�s�d���HK�C{͝!�yW[s�9�L�:Q^Ȃζ =8=��m������OC'���H�-�^�j����z�.���wO	R�r�]u����,�i��O {.��S��!�$��'�� �a�����~���t㻪���^�/�=d4;]����P�)翪N�)K�P��ekǸ8i�1���X�IB��es�6���@�h�xң;���'�SL�̘&7�{qp�S:�K��!y�\�6O\T�,���<�w֑�gY�͋�ö,�J��5c�MԹ���:�X���tA�Nj�ۄ�[�F`w���ܖ̡�[3�:t컪nR��bC��yOΫYw�+5i�a�`��0~<D��9�pC�gFp�p�I��RL�j�]/�-�F3����j�� uFk�����w�0@4:�	qRݕs�\s�CF6J~�yl2�M#����z3ZltEld]��+ynFi���w�OE7Lqm-�Ms�^G`������b���!?8�pM�:�{��L@!��6��e�E1�o\^���`�eC/�YS5��	�dv�9�p��]n>qXA;��A���f���������N��ʗ�]�q뻶�7M��V���6ϼ�{��f��n��dg�S6w���yz��Z����-��Y���ʍ�d���ɜ�ZW�@z)-�/�����(�m��GG��kU7�p�����]�E�c����rʌ��l�98��Lۼ5F�OW�U�q
�!ү>�p��Q�b{j�i��52��`�;e���tm�l����n֙A@�lͻ�Li�]
k�Nz�U��Ǻ"_y����<;Hۗ̕'�jn��t�U�;�w�hA���i�?j�U�ij��fn�P��Q��G5�����.І�p�0r�g{�LH��:�qZwl���-��r��/��K��5 �W���iŖ3hV�u��4�+����v��.���l�̚יo3I���Ǟg����\�O@�T����D'u�薶xiJ]�
s�^�b/w.�ZnX����ىSu��$,qϙ����ϻ������>��WD~ض�koT�]�ӱ0��K�3�(��Kqջ,��OQ"�t
ݯ��t�^��g�+�wHh�~e9�Qv�T�m'u�h]1s
u�q�p]�B�,l�ep�t
��M��U��sI��C�Z��鼾�sډ�=r��Z�����J��c���t��ӯ��giCZ����i�X�	P:*"TZ�s���w�λa,�q&C�4�F�T�f��(�H�Q�6�'�95>��e>��N�tV��*��G6F��E ]�_��ߔ�p��a��YW9��_N����t��x�9Ve�N���2����e�^{fA��.�l)���.]��"q�g�����̖IT6��r罭���yΝ��9�D�d�x�O=f���ޙ��-tμ�F7�E�@sb�4y���wl�ن�kj��uͽ8�W9����Ϩ�[u�Q9����8��̦�]�3�&@��i��Q�֢���1`_pA5�VX��$�3ka&�6#3�9�PgL�2i�	�3��c:�3[a���v&�J{�X�����rR�RN��H3u��[r��K]I+��AV��d����W4O��[�://SW��=;�3RrYق@c�Uj��D��;�KT����l����Z�1�{�~���m���s�(�,���C�Ez6�Q�l��}�ܕ"#]��-��tr�T�g3.@�I�9�{��jm��+��o�)�n'zf��བྷg�r�E�]��fS&��hע��ia=�qJx��By��i�+��{�PCW�c�Bۦ1��l�`�0���7�q�Uq(�KFȎm(�'kvL���.���G!��UV�~�x.in�ыo@�J)�[]�z�17�5����zQ�1�-�[\lq��Dj�dY�O`���j��.���sQb]!�R�N�a� �O���q�Ww7k�t��g��)��9�X�YW�T�)�3�;E4.�pL i��y��H�B��>u>i;����.]�\�=���mPP�&����uL�RA�������Z����y���Ӥ�k%����|y�>�R��R��t�N��g��W�'��<�g׍�e���h��vϣ�4�P����z�U6=yBƽ�<����b4�J���"3'����om�w�mwK�ɮ���f�_FJpo���W��탫��glp�c���V�H����7�\�n#{u���ou
��YU�U�T#G*����Ҩ䕷�E�Rxu��ͩV.��˿a��ɻ�����
}k{��"�H%Ҧ�bmN�9�61r`���{��򺹣i�
�����fzyYu����o�I'z�N�<2���s�-�B�GK�u�D㻚n�~쨙w�~i�&�>��Ut��&�\�m<o����ؤ���ȭ�xe��H+�ߴsB����!r�<�z����*U�*���q��n?�<?�\2�Xݵ�)�/):����ƪYd���˘	��S���}��.꯷t��9���Lw�����X��cY�G�"rS�3���ڧ:���.��9��u��#VT�܀��(�;�<n��������^��Wq��Ȝ���Bw�O�ZdxDH�Ϋ�Q��w�唝�ͪ�h8ݳo7�'��wE���1�cz�%�5��=Z��b�mႱUƻ,���|�هO��&�訮:���7+������%��2B}3��Ŵ��Q��LXH�u}��|ulg5s�3XL�
؄�H�vl�\�u�f��r�z���AOn�Ԩz�T�զ
�t^��1�W����tͻ�l�ˈ=Mqz,����a��θ,�`[-a��q���O��u��6q��т�@x���R��m�=1�<�q	�����6�"-���I���P���B�j���<��h���G��e��f�Ƈ��u���yZ;�^�j�4�[��X�-�7#ZÆ��=���t%���د�����~�͔)䦂�W�R�G
����,x;��	�b��#ŕH��
��ˈ��/�$a7S��1�p����Gz2�[9Ɏ��M*�7B�u��0�A����y	̵gV�=K�&�^/dE�2+z�o������P�p���=��QM��!ҊȂζ ==��a�Ԧ��#[���Fj[&N�4�6mk��t�$Z��[v�}yf��P�L��2���)�!�V�ȇ-�G�i�/���4�$��h�	��܄���*e(�@�\$�ӎ��S*C�~�ݺ!Ue����y�钯�ݘ4܇�1�2�3��N��t�-�B�Fp�\;��uӹ�V9������0o@H����ђ��6���}ˀ���<���	�|r�2��^)u81ӏtf��Z�Qᥣs��L��*]�dl�U1��*Ye3\�c�`kb�q���Ā�lW=�k�mM99�5��-�צ\l!��]3��w����8������ʯ'�oq���Ft��X~�6�N��S���ݴh�����3����{��� �/2YX�k�]�}��z�o�$�aӶ�CH��.�&T��zs����W�s*]u���Y#F�t�{�fj,�a�5�9����q��f
�<�(n�Cn0�Y��ޱ��̜�&�b��o��e� ���*�g�o}�����.��{����__{U�!�o���'�8'K�+4��j��K�/sⅭa�f`�{�niP:�I\���:[����(�*�P�|�wѮ{8�������vi���+�],N5�S�q9]����'0�Y R�����ܝY���i��m_��݋��Vx`A|�,D�]�{ʕ^"�AQY�ݨ<�.�.]�*��c��I�V[�v���M;�a�V[ˮ:�r���m�S�VV�	��]o��"ܤD"{��OJ_t�.�gv=�KZ��4x�C.����X���c�a�j�R�\c��>D����U��ٝ��B���"W�%�1z���we������B��a{��A�dv����+w�]r�V�,�f���H�QP���O�p閵�h۴@A��X![;���"�x�U�C���T��й��i�+p�'�?\�z<p��Gg�R�qӊqA�59#��D�:�W?���z�H�o�vk�Q�=�?]��r�a�ӗO"�P��f��Xh�	��I��U�ћ�xѵ+E�OV혘T�\ܕԻ��$�j��`K#�7�p!f��P������n��M�:�&&��<ۮ����z1�Ҷ旈g��OnE�-�VL��E��q[mVkO�AU�qv���.K�3/���"3���7t��I�u�釐���_%{2�e���R�������RM/h(����S>MN�����y��k-��t)���wƈ��������ra�ͽ�@@mXmU�.z�0��ȏ�k9q�4��&]��':��B�㏡:�F�I!�C֬3N�!{���G�*�z�;��59Y�m�V]��+2� �W"����*�4j��Z��v:G��.;$��_q��#K/�-yA�,�
Fm�΅b ���2�\9�n��*]+�Fr��e�\�΋�E}J��<��6N7����)��~�<��G[9�|rʐ��}xl=�R7�ԖtĘ3��-7:�
�F1J�=�)U�_m9�r��/p*�G�o$�|;8��t�S�wd�
H}'��դ�ӷr�*�	�ʺ*�����ˍt�,��z�}L6e�8�d?i�{��˧K1r��7Ҋ��٩�Q���Õ�����!��CtKd�V�LYC�$�o	#��*YD�b�������A|rn��XۓV:W��7��H$�ʡ"����@m�]ɂ�e���l�@����;2�q�d>�Q9lҙxo���I�:���o�N[��+�v�r�Q3�P���1K{e;m���o��P/��sAY��vU�V��W��gcǘ;N٣���}�(�7Fd5�XN�U��뻻��U$u(�E�*j�$Q�'�f����M3�J��2�r)V�H��$�UDEQI!F�PXr�$0�t���rB"�\��<���%JH�Y���ࢋ,�C�Q�t�BB�Z�� �f�E�9T��P)��f-���t��I"�����Oy�p���ˉ�ej]%G����l�"� .a���4نW��%D�A<N'YSĹaDR�
#9��5B�ʕD�@HN��AV�w��Ԥ��N��D�.AÅ�qҢ��&hX���PH��"=�/(�T�3�E>s��D�"+)B��J2��B�ر�E���J IUDR(R�-0�̍�!�D��ШU��pfF�W:AIhb��QE�EQQG)et��f��C!O�S<��2��Y�EUQ�<��1$�
KD �U�f�2�./���%G9g��<
�eH:ӗ`s��%DH�{o�KW.V^3�Gr4-Ƣ�^=DwKǪ�Â��i�T22D��$��n�5zθ�1ɿ��7�K��=V�`�ϒת��ՅVp3��M�a�|�{n��h���qQj��=�B88>X�3���|�����Ά�P�F�~�dz��Ԥ��3�3E�K��w �c����(��]�j8Wd`	e98��S���x'�\F!MqB�؇J�g�[�n�Y��G;��"����C{����]��o��k;Z���H(�i�w��!޸7����6:��\f!�+pj���4�Ƕ�xDj���ܗO`�T�}��QJ!;����x��.�����T�ʚ}cI�Wl�,�U棷�I�Ds�����>�7m�]=<��@�8t�z ��D�b�Ǯ�<sF�;�3�]�z޺1S<�n��Y�vYS)�$Z�-�^1箕K�.��

��o�QˍQ�3�x�s��A����{��m��O�vY#&��`3@"����0u�+�]u��s7��oN@w��M<���i�g@�4���:gOY�:�JgiCM�1fB�QLg���}z=�ё��z턫������tݹcJ3�1|�g���U��������ǖl�� �/bϑ +pښ��X$Zu]�c(��"�I��݃�"�Hݙ���9d/�y�94q��r�c(�ܐ=�mrH]	!C�U�#�]\�;o�b�a��XDC��*�>����M<Fr��ٹ�;r���#�D-�O́a�R���W�!�5�о��Dĸ9?οԿ~���}���=���gynU��#7�,���02���f�7?v�6�9�(L�����l��a�
�w�,��Qr�>�b`��s�%��z9��.���z�N��W{T��u�E�wj��@A�G8��;���<�C��E.�ѳ�Sĵ�t,���Kl�_��M{8�W9����<m���B3��y��F��̦������]���cZ��A��$�(���/�|��\����g3�g�+O��}��>��z�����@ge^��V(4#��}M4�r�CW,y� P��)�Z�p'�3��|U��X �1�(	�ѐ�\g>��w~k%RBr��J�u��2�x$/t�`!��Y�OMq��{AӥŻf�]H�17�''��wL?>�qU�/9O!����!T���๥�򢼦-ʋ�kw�j���GPm����0b���h��Fw毙HS\Br��eO���cq��~Ξr��L��70�]�v�q����dȧV{ݙ���/��
�����e�Y�,�ϪI��۶����x5�}"�0� ݄���>��c��sjw�Y��6��5Xr��h#G1-<�t������7.�&��V�#�#��Ѹ@;��U�+��{�{*�M��{)�Q�g�]��K��v�T"��3Q>�kn�+%2auc�x��O;b�X���[�s��e��:���j�F��!߈AC��i�{��)�j
��NN^ֺ�Ґjf�ѵ�bը��/�V���w�MO>�̬�-�@��a�s��a�Z �6,(</9-[:�T��$��5�Yt�zpS�i�#�������ʹQLm�4r���L����,Fc�*{m���˶���R�ݦ��b`o��p[�m�oU0w��)�v(��w���Qk2%�k�g~U+�1�����b0���<2�%<s�[4���E����y��zh2���V�"��ح����E��\3�p9�,#]X�2��oX��C���/ܺ2���*p�9\����*&�I����'���/��~)�/):����I+��ʵ�4��OY�'#E5�M�=�2n��3�ȡL���X/�>�?>�5�`�k�y�X��9)�	���S�����[�z"�9��MR���[�A>�A�t�/#%��v���' �}$���G���լ�3gA�N�۳D;�v���m�+A�㵏/Y�'��<�n�0�L��q�˥�?6�a�`l�S��tCl����H�A˸��ޙ�I۬:�΁�Ù�
�ʾf�Kv�3��L�������v#uu;.�{��O禶��R�S�Ϻ���5��`¯!9j�@��Tq�j�Q����M����49w�}�r����J��Ӌ�\�UE��^�{��t�|����u�`D�9���Kqy[�_��bz�9*�S���==`�:��t٣�)��� ��eR��-Zt�
Ȝ2w1;���&�u�f��L�PC\G�m�L�s���
�ú)�(k���J���5Ǩp4۪���Tλ���8��渄�^��T���}�rX5?m�?OK��fdd6)����_Su�ɄoJ�MХ�m��=�BA�Z�
o%9	�u�<�}���=�����Ms�w!)��t��>����C���m����4�`lP�R��3�{��ǔ�V�h�޼|�[��N�OL�zI˶K�m�A�溕CחOE2���0r�"�E�\EJU\����ͲN*~a{<����g��we�3)��.5�>+���[e�<�\ʐ��$§�� �	���{u�p��/���@{��-�p���nL�ep� �;���2��5{��-�6��H'��2��;��n���2C����p�t�|Xu����{�C#l�ą��hjr�@_L�jSz7-���=�N�4��:���:���C7D։�Hqf)���L1�+<�shG�Ԣܤ	�����GqE�;�+8�~��n�3i�S{ǀynG>C���]Iw�1�&wiY\���VK>�,�#J��F��hݿ�>W{�e�*�Ö83+"���Wϊ>��g�n.����1�m�T�ˌ��s�B�B�J~��젖���u����~��>��D=��r����\���w���c�ۍ�����'�!�iK��f�[`�#N�[��%����z�28>(�3�!�B=�m雋��u� ���ea�-$�Y��V����I���5�m����9j�������)��=w`�~WF7Q�˹��t�U��e��;�яus��^�&��wΊmϒת���T��n�m#�i�|��9R�i�[Op1�N�_��C�n��pb�z�p*��gCbTc��^G��Z�Q@��k�a�"_7g:7�-��טi��ep�H[)���f��x'���B��8�{�5*AP!_?���5�	����EvXO�t�����FZ�mG=��S����xf���
�w&�dI�/��a����W.�Ǘ��Տl�È�]<�c��Ċ�*�n����5�+�kg�*��SF<� �v�:K�;��d�-]�ʜ�$Z׎#oݲ|�������
�C�`;m�x+E�w�l��V�=M�d6,��ă�n{U�Z���u��f�1��y�xs)�7n���ԟK���e�*V#ԅ"����<� u]���M����-��Q�2,:l�Gbꎻ��]`��9����������l�۾�7��([[��-Q�;��Y-[�ʔ���� ����=]T�<Sa�u��5)=P2�C����!��}�S�[:sb����n�*e;]��#46nLħ��ƹ]-��w8+p�6�����s*C�L9��]m�f�����A���=�oN�r����ܺ%�Q[��^�71S��Ftƻ��L#��C�{X$6�n���N �(�H�Qϻ�q��O�n9[@�;�Zj{��$y�i��j:_�-ߵ���	n\��0g��Z:��ǒ���L^����c�����^5���e�<�)��w�m���xc{���Y�"i�g��8�lkt��g��*v/������z�N���d2�j���̄s��3�̪�[,�P�;ȸ��a��yo�B���c�#���:�������!���ޞ��fB/��r����n��13(>�uaF�m4�ʌ�D�V�d�c�+m����3�|3¯m\�xt�o�����7������{ؼ�mSMgeF��rǝ�}0,a��-�x|%�����<�nR�Wf���=��QLՌ�M�ە}c;_'Fܰ���^���=��2w��:9ئI�݌Q�v�:u�[աN'ᖏ�-����Ą��Es'�.KKe,�z��q�w�f�mnO�vq�U�stV|���<j�\�>Y�����i0T�{�.-�zY��ʹ���"q�1�Yr��{�PCR�yH_�c0l�-�%�ԧ<�:��׋;�[�d��}Ӷ�1��6�:}G��_�2T'ޅt_�h��ִ�
:P��3�����(���8���oi��B"�Nx�rʼ���_l⾸r��̧s�`�fr�l�kn��u�#���y�'�b��3�5G�b���el�	̲�~[��ۅ��j]疚����nɞ׮�l�X!ߐ�7A�u�3rХ;�T9	�����T�u$��-��e�.��컛�DK�+�	�L���=!=�!�!^�h.��f�b��#���[����h�Vnz��7����2I	훺Q^���i���<�\��6�9
�CAu�[J��	t������U��z��������;4���n��u^��`��碙�hDktC�`�O�iC+����_F����*E`$n��u�<�ϋbPL���2��w2ˮ��]uK�>�X�o2�;d�e�{� �LM9|�fH}�R��8;H����XzD���G4)�~<����;����l�hW�}��O�����^W7���u�� %�����k�fi֫��Y�(l*t��؃�r�Z>ۇ��y�<>#"�QG���m�9�!2s"�6�d��l�HV VȺ�<냓����i��Lw���6��K��Qϕ���Uq�#|��Y�dt0��8J���+�[���b�g^x���� �[}1��F�ϵ���q�8)�G�"rS�ht܎��u��oVD������2~�S���T�b�ݱ/��j�����Q����'���N$M65w'�=F!����<�JwYC�x��w��]�c4�|{]�Z���pSt��M��+���7[�n�a��;D�sg#=C8;��ه��k�N�TWdJ���5:����^�d�7��լ��&��d3_�Y����=�6�Tq�V9��[�)��3zن�ܻ����}�l�7+�sH��_��u;ҿ��#]�սL�� �j��=��>��p:޿LgP���AEK!وf�;B̙��;�oi��ڎ:���w[~��xf����n!!ڢ�����G��U����R#���SB�n��n�I��z��m3s�H;Ϩ�৺�̔'2]�f�+������lR�=7w*O|^	}�%uu�P�<%�`�J&%�=�M�c>�����?�Ӑi�������mc=�N��n �����,�q^'ҁL}8�Ui�h��Ǥ��oN�k3g���1�nGH��à01K9���
�Fu��PO��1��-�%h�K�ebߟ[K�u<2��_���{���+eJ�γj�hIs�c���6�Ni �^�P�����-�}S�Ҟ�E���[w�/W�կÄ2��cK�� Ʈ^�sr���w�Q����绦g�\7:k2���l�:�ߗV������[������lvN�T���ײ��d4sr%F��u��k �Kf��u2ٔ)�<:��i�U[�s�9����t�;�u2�;�7����$?O�yf��m�'�2�˺������ڻjn1�gV<nT��X�e���b�c?R.��W= ȶ��#D�+��Z�`K6(��r
P-T�c�S��g���ٴ��ۺlO(�]l��;�qw���s��n�s�+�
9j����q�ӳ�����C��q��.�*y��A�ا��n��ǰM�qx/���.��:��U�2#�J�7�1�w�m����4�މ��{�I����|e�N:�4���{�D��q�v3j��!�Ĵ\`u����i՞��K�`'���]{�٠T����K�<Ma�i�P�3.��/�'��B,-��gCbT��������9_\�a�����%�)���=���o�rX�:�z�7�|*U�<3�Y~�=�񵨩�b��*�����{K��Xc���9�5�桙�L�S�`EoR:��N�,�`u�ñ���ϭ��Xͤ�����F���¬R+$��Kk����h���_�x}����4�Sg\f��# H[)��"��7�z��B��8����f:������v�g������?!�\�,�6_v�pc�Ix�W��+n�UMo/F����\�&���qn����2��F�eXOCWV=����]<�^St]=�66�4t��=w�$�u�ɌP�<qz���m��9��D]vKB����>f�w��G]��1#���z�����k��u��;��Y���D��d���Y�@ �lݯ��Oa�~���V��g�߼vv���
l��Cnb�Ol�͊��\&�e�)F�A�I��]4T�븻��w�(w�l^��|�R鸴w
�CAu�3`G�Tow�l[:z8���g�huuln�����<�̚�kn����{�Xg���z�Ј��M�v�X���L��k���,��%�Gt�u<�3�=Ϸ&�s������C������Yg	g�S�0��5y]s�O[�h�l�7�gx���Ҡc�
wg�Ä�͆dp����|�~Qr�ʄA~f��=������d~qoQ��+kk�6J��
��e�b�u�#�E�V	C	ǈ�Y�nў�\�x9kgh���h�x�"p]GW}I��s�����/�OyO����� �7��F����N?��o���d"�P����d7��{2徭)o�����C���"^4n�����V��qe���YKg���`aA���7�&亂��Q�yJ)�t[��{g:R�L&^u�);��͕�_3u�5^�.�-t
�^Ĳ�wQ��&�������L���̗٥��y�z��?N.ܹyo*�Z�^p���uwk�D�1�֗u\y����J;x;cLM�@�ԛ��Y�.�h�����T�5�o� �2�熞nuq��x�����&h�fأ4P͘���B�r�����,�T8;��mξ]�W=�K=���[R���J@�.fܻ�awDoe��iJ�[J�z [�W�z��3.�K�� ����L-�/�w�#5|׌��p��S�"�eh�a��+��*i�Ch��z��v��靴I=]9�U��ÜC/z�rU�k�t�\s�L�#4'eh��Ӷ{9f=K�1鷸�_1.�M��ݧ��p�|��r=����Q�N,;�if?*o��]��fd�z���7g
��5��WV�e.��(�1+aB���+S͕x5].��������&\�$N(,<^�\TvO��9w(S�F���m��4�&��^���w\+��;3�]]$ �<C��u{^�TKX��H�fY�u��k���R��Wv��Mo��dm�v�����ǋ��k����Wb�uf%+3hK��'e��pa|$�9y®��f�Y�*��8-���0�w���Aк7�y�5�S�\E�Q�mwQ۾N�Z�^D�}�U�<�Q��ps*Z7�S�0ш����x-� �
���8��4:C09�H��j��+���[_]��&��>qn���<%�l�F�$��w&f}��lut!k\Շ[�gC��^���_NѮ�h�`Rk�b�+p��q�;�y��zO�G	���uq�U�e�]S�гٯ�	�"�����[�q��N�΁^/�T�I�'n����Rg��_Zn�������X���s��M��Ԭ�}}�CY�{t����]�p8�;��M��շY��Y�����خyb�;IO�t�=G� N���o�q�1!2��^'�jMK�'-���\Zڃ{��eqT�T�Vi1Fd0j�c9վ�7<�}���f�q�_-���9�:�#eH�szΪ����;[�;*9G� �7hV� DI�l�gP�y3���ĢbU�Μ�@m���5�v6�����q����Ckv��h�[A#g.�Y��&���.�L�-�
ı����(���VvhJ��u?���<t���1v]c�&�$���:}cy��,zS����@w{7�M��-+�yjh��Y�V��ըR1^Bt1�w>z=�ϝ�y��Β��*�(l�
�ybEQR�Pr#�����q-T��̓gd�Q¹�32I����
�O8Yp�E��D!Q"��eUP�W4���yhp��>Q�rM�Rd�JY){���.��-١��B��g"�B�N�$��H��rJ�t"����<)�^T3�3��*���3=�M�w�x"�(��԰�)eu	̌��%�Wyh���G-фs�)"�+,(�jΦ��T��ל$��J,�fr+0�>W��"��aD��g,������ʉ��b�f�BdQ�Ђ�Jq!�\�Y�:U*Å	)�J�GS�*�����a�Uv�H�E���U�x�R�i�V�fT$!A�2��I�D��I�$%R�����@�ʂ��N��3�6\�����r���5"��:�!M���84q��p��`�z�_��cKf�ZF�]j��e]�|�_@)d��Z�a;���ێ��/��%h�@��\2��sޙ���ds�{���cQxN�����wA�:t�S���!�Xƌ�{��u5;�?lEhN�g��(���9�{;)�]xu�A�E7n����"ߛ��Td��+mZ��y��i�=��hr���(WrՆ+9���,Pκ/A��ط���T�,tCw�2��F��×����U�nNW;��)�YV����J����}�]t_o��PCW�c�C�]�b�?���SF����Q��y�����B�!9V�0����������.�̻)>����n�ы�7�����)Wjz���5�^�:%��Om1���\Bs��\��}S�-��r���қ4���WTGS��E���/ۆ�H�{�ݐ�k�S�ض�n��Gb���i��$�e�8�x�u��e�%�fVi5��s6�f�=��Ac�t��o�a�aJw��(rm���l����GdI�1V�\Uԃ��Bud�vXn:�On�:�K-g자��l���o�0��h:�vK�_���m2��n�k��Q�R��vy� �֜5�z�}������:$'�^VE�.�)������uC����8ed]�-])�(%���w;�`��ͭugKr�y^
]�f]�n�lӆ,u�!�]F�Y�_] �
��s/2_CFXl�L2a���_~�l��TPO��B�k�w�W�l��Ж5�<��a���t�gmk�Ü�/�N��ڳ���W�c�$f0�Zcts�)٤���V����碙��eэ��a������we��o+�$S`(n��+Ǟ9�-�B��S�,a��Y��;�t�5���,p���vp~��ѻsN_/ْMt�	���V��L�2�a�)��w�2_$6��-ݚ+1�ZN�\�;�.]�T(
u�'�越�|�k��W���	�DO�'�f5T�8L
����$�����'6��Ŵ�ş�O ����w�X/鏸m��ϴ�����G�")q�K�Lʧ'!�
�ߛn��{��L��<6+�%�{����qw��L�0�h�et�=�:��Z��O�L��f��|D�t!�þ��Fiz'���ی���+^��N=rǝ�m��أ��j��r���j��wkQ��;�=-�޽��M����0��^���鰩�z-�n7Z��{����+y���m���B7��Fsd�>�t���T�W���P;�)��yи-ꖼc��4�a��Y�O���J���ɮ�(�c��ߊ�i}+��#�.��J��͋�����7LHC��m/WM�����ؾRKD�V&󺅮��Ps�F��P �V��V�с@/9��Y	�
|�wneX��L黜8<�����X�����-x�F9?2ݘ@��w��S�Zf�ᚷ��\AP��ǣ\9k�=��-;�\���ް5�sg�s�Dvt"*	��dr�y���y�J���/�|'֗�1۔��#%,�������{�u'B��+�n�s�6�biT+�
]���=�BA�᜘�VK�6ͷn�64��'o�
�	�z��_�۹Jzn��7�K�Muu�w�!���Л":�M�:��)	��ڻ�sU��T�?z1J�~ ��!�-S�Ҟ�E��.�����WR�z]=ɵ�(�R{�����w&����	#��f:���\�x�;(�`�p�m$�+hF�r�pi�uc����Ge_u0˭��;kQ��ߩed�P���Fp1P�Tn�8\3�
Ķ��t�-�@']��M���_]�vwp�f2+���2�ܕR���zC�wDm��n���$?P8!�زy���{6�T�5��j�5.�x�{��A�	���Eӽ2��
E5Lv�qR�)�+X����8,X�靭�ibt�����s� /xe�����Q/�h]3��qw���q����n�`�1��Ɋ�{v��zo+��:��67p'�AP�9�V�+{K����&���Ƀ�թ�zU��`ⷪ#�e�E����u��i�9H=T�s�A�Ѳ�!���tkߴ�1�gMb����)������Ԃ�0h""m�'cX�&�MPj�{Tk��N�m��φ  ���@6˦_`S"�O-܄�^0��B)�k���㮎��챡Cekݖ�kɜ��b�����*w�Ӝz�ݹ�/Q\u�2�ع�8�8�4I��;��d�7�Ռh�Ow,v�E`N��MϚ��$��
q���n�m��՚�9�Gm���s�*�n�8��'�k����kA�Bf�ٜ��Yė�����n4dξ*��g��F��^��T�~�ڂ)d`	�pm�m�*7�z��@LO�5�t��Z�u�������Ꮮ��]t��Vi��ukx�R�QS:�ٝ�4�nq5L��GyX;D��א����'+aPN��m��^8��]<�Jn���l*m�wK�Gb,r@.������rb�V�7}N�y�Z��s��|�`���Y5�,�ʒE�D󣱏o����F[.�j'*��Y���Ѡ��C�fQ	߶/�!�%,��Gu�d�"kvY(�$] ����v
���,��n#%������3=!^wH``P�i�{�hS�]�Np^���5X�i��j�O	��~���mCف���V�j4��&A���ռ���)�$	��te�А��j�H�t
������n�]1�37W��#���Wf5O�8�3��ާ2��ij��2��wA������Xb���1�[�~9�w}����O��z��}��ǘXs%��u�M���R�G!Y��Pңxc�0�81mv�Lރ2���b$f-�6jz$vf�}���TwDttc���`Үz���F[7M�v�N �}c�R�`����cI�鑶5�9�όH��J����w��w�<%���#V����캜���s�°��fv�X:k�<��F�S�131C�u0S/|,���W��@�~�_�d�!3��ẟ3�S�
��n��������-�d ���`PU��cpdWU�P]��=�B�<.��s��ѐ��S��������N_cp�l�Q����zS}��
����T�CZ꘠x�pWK�|��������pW�C�G�=w�ls�`��gr�w㦙�U�g���M�}M5��
u��a����j��o�O���{�P���8�O����~�?zm�a��B��yj«��f�8�˲���CO����N�N��~Q�WdgRɳ�9�G7mN���7��[0��W`��S�n5t��r�/�l�D�*��VҮɱ�׶��m�����yQ�kB���x�&GYI��:P��o�{}�VJ�<ߣ���tsd�*q,�'i�q��`��~rQ��d7�s�8��מ+^S|�S�L�)^��XaZ'1�w�{4��j�(2=�����=�l��n̺�+O�v9qȟ�o}G����A�se�8��!9�~%KD���l���}|��,m�˙;��D���m�ݒMi��ٓ��t;Q:�\�w�2�=Fz�>���dڠ��>.%�Y�18ZIۼdb'���z;E4u�s���6�;�)�����{
���"�� �cX�lx/���|܊���4^�=e�}l��n��!~:���>Ϣa������q��ж��Ƹ{���vH��1���4�fW�Q|󚺩����x4r솂�bc-���:��|ʬ�㨻snV,r2�s���&2yc'�&��sܩ��7uЦ{��xm�y�4��h_Fj;ϛQ��m�4��{~�vYᕉm�y�[4�����j'ܱ�N5W5����݇:�b�1g��6�w�B�}����e�f2<�~x���?��O���a2�z�4�Nk�P��"����ο_�`?j��6��w�[�n�O�~�S���@�`O���t�C Q�_^�޶�k���\��A���F�n�~�:�=��h�>CF��{y8��-���������2�,��.,����R�u�Hc��Z��A�˱F�g�vR>�*VK�C��:/'*܀@��j��a"���E=���3ܳ؈?\����S�7� �U�1���}@�2���vbc��O���eʝ�+���+���ܣA�2��<L�芆A��o��.����2|Q��7�B��x]S63w �^�0L#OW���ע����x�'���-��O��{��|;	�(� �D�W;���SO.z�[�,y�U��R�D�	�I�g��l���c{#[;⭖���.�ՅVp3�ӎg���A99�2z��V�^��ջDqzWw�g���>��Sꈾ�tϤ`���W=5�.�� �^E~z��<O����~��;.6���!��^nǁ�n�U7��J��i�]:������[�dL�*��ξt�d��'�U�l5�5l�(R�N���6�CϪ8���s����(]��)&�[�3u*��r�>��������e86A��M*�7A�u�閰S>c��Y�Fy���(`w�n�Z�d󙮜v�E/k^8��v�|�.�����k��\�vNxn��nc2�9޶}\�0���ݒ��8��l�Dܒ�])�~U�A�箍K��+A}t%��G$�a������w�q�"<
�"�Df\4��*S��/�'\K�XV̸����I���p�����$:��L0@e��߻oկ�6����O냠�{tD�n�B�mb5�9^Y$򩻏T��k;��<�F���b��O��R#,��8,_jA
;�F�%I!8�>�$Dз.�����\��Sѽ/���O]����3������!��TT��i1�2�.��V%�:[�(�c�[}bN`�ֻ7��]�l'�GdFh��F̷u�K+��P����7\�y��L����췹�ރ_��o���kMOm��]�&�S�~1p���T��� �4�q~��Yq�-륱J]�:}�WE'$�[���'�%̘��C��oK��C��1�gx\��t��\�q��Sw�Pf���h\�=a�5��������g���̄�O��2��D�s�"��,�O�_�9�湑�*2[�SY�Uq)����.�'+���g��\�E�"e	i�G�M��/�Nl�u��6�͑�b��r�J���l;>�+�>M�x�ܑ�uZ��Y��gŪr���P���_y)m"��i���\�C��|6�)�}q8z�3��:9?j	����*8�I�K=�j�P�%���ۑ�[�J!�qnL��To�]P��Lu�F����C���!ԭ��o}�y����-x�j��4�`���i�K�l��s)�PS����̹�2F1	JY8<����޸G��:V��.OPYO4�dW�e�u̧�����m�����K��r�*�̼�A�}�L��³��(������zη��=���bSpt�ʓǈK���HӤX`C�)�w��m�i�E\Bs��*�z��Տ|L�z9�1�]7B��ܑ�Mhz�=3��ME�%�σ�"��jg��2�-]���DO�{%�3�$��׎s��M��U�gM/bl�KDVfL�1ͫ4��A��ktAw�<�4L�Pxw^K"&�J]D��c��MUkl�$_c��<��Z���q�����%�!~S�,���������Nٱ�ٵ����44�љ����5�l�/\�4;��E�����R94r솂�m��<zTo{͕�X似Cڗ��ӽ�3��[	��m�����+�ю曺��d��w�,^��|���	����e�q�$��Q�@n�N)����Q��O,����:_�[B�w��gy�\)���=�1ff�����]-�L�8쥩N@��;����^=w�C���~5�]p3e��S9}����N��`�N���c2\�~�Wp�o'�[�"Z�	کOXfG�����]o}�H�\!�;3����B���"雦X��O��n�\lc6�<��jy}�=�z�'MZ�ԭө}��d2��}���[Z�S��Ζ�'j�]GOv�wj��ƞ��W �=*zu#YdM����!�f�S��2x��᫫W@^ŕ�D�eM���Ƌ��ԕ��fV$�LhX�ߊ}�8����,����1��[1�CE6�w�N��T����_���vCeƢ� ����_*2Z��ӎi��pU�!��
|��ꨌ'�ϓ̂w�R4�$ʾ�{f��]���Y����Xy���F�m�|,ܱ��&Z�l���:Ol";:�S6�?e5�'w�*{D[.�}�h]v_q�'HjY�)�+����%�I��O�s��?�K�+�c��&�����-�w��l��t_)�Ct�������8���|���c�S����ӝLmƾ5�<5E��OX��<�a2[�E>p&g��Q����~��MId��.���%;���n�&Y�c�Ÿ}�ӝ�ɯ���
w��s��bi�׉���ذp��^ȳ��U�cr`���;�)��������)N�P_���#�X��э=����x��)�wu$�����P�ԩ�?G@N[!�!Y���a�Wq/t�{]Q'&{q I<0J�4Wd6�NN9�2k�'��2�E��|�t���QM��9��ԫNmZi�ɀ��*k��[�S4���l_�Df0e����!L�.S���]�U0��o7���{�x�1���Lc�����1���c��c�����co�c�6���1���cm��c����1���m���6��8�1���c�z��1�����6���1��\c�����co�lc��1�cm��1����
�2����"�� ���9�>�H��EUR���CTT�J��RB���fR��P�*��B%R����(DPPE
�$%UP�
�$�UUR�J�����B�I*��}ػ$l�
�R��bUP �AUI*�(J�%JDځK��IR�����$�;wem���E"J�QT� 
��͵�D�
�B��&�J��m��J�H**�U�*��T*���bّ-eR��˪�Ul�    A���p�*��R�(UQ�T4�(�V��4�ъ [3LT��6CUPdV+CEC�6�J�T �^    ��A\�eT+Z�F�T:��E@��$[���QE
$w�wQEQ@R�ۊ(��(��9׭�I(����;�(��(���n(���-#��(�)�h���  =�����pj�)Zʤ�`�
5b�	���j��PK5���Z`IKmB6ڠ��T�4��4IQO   ��jԚof��1�����VP��E�bֹ���j�(j�6��43j�n��d֨���ݵ7r�Pl�hwgKf�Ҕ��C�qj�"P�*��;5j�  w��m�SOn��Y-Q�fƊ��ֶ�5�lJ�[�ձ�MU`�N��]ʖ�&�PM��v��v��L��7SMF�Ed��.U�v�"�UN�"�  ���Ь�6��AT6�������,�nçu�Z�[cE����:�R�C-n�N��ֻSU��Tʥ��L֍P�m4�n�4-"��R�ڝP�� �x  �q�4޻��L�SJ
����if�+(��;��������+B�mm��k.�����5��J�u�㮀jk]��W].���J��(�*���x  {`mb1jհV�P@kL�3�0���)������]w-m���[�(;��Xmk4	f�Ց�Wj���F��ԫ�FR�@�P��   ۵c�N��v��Մ�)ݫ�m۸Uݕ�l798Mm���M(U3MV�EFY��nխ-kVV��N���n��v�r��T��(��
�'�  �{յa�n�r�CXZ����(�Ω�Z �Ԭ�N��Z�P�cl���7D�*2�UKVQ+	� i�5�����T�� �S�0���C"�F����  O��T�C "����Tb�C	4�eTH ��ÿm x���`����2�A ��`�*���w���}�|��H@��	!H�B!!���$����$��$�	#!���}O��h�����=�o����1!nfɻRB۲n� mMt�	�R\�[7�[@�Xl�-��,�D쫒�l�n1yV�z4�5",�� �kܐ�U�0�z��9v.��6)l��E���۴�B��I�)�u-9v�J�S��ۚ��4�b%��DF�%xw/iʽ��W��y#`��&U�z�����{��B,���	��yE�AY�Q�B�kX�4��:��l(�Yݦ�.=j�0m�IS�n��
aY5A�!l�v��`S�̬�{#r�'{pҩ{�pb֫V���3V�j�*ʳJa.�X�}kE �^��8+E�F�r�j��TIKQ��r=�	N�b��5��櫀��y3�q���x�TqL��bU���bF���ʁ[�X\�gqĮٗx�$�]�v@W�M$hʶ�	n�[��
N�F��V�z.��i��c6��*�m��J��>��{�e��F�6��r��$��n6N�Y�uSa*��kc��`K3o1]Ez�F^1�R�"$1�w0�i�_FҴ��Wn��u�h���N켔c۰�*N,�b���.�����J���^e���pl���h��ن�����j2����8^*��.k�v�t��fS7�R��X�i��ܷhJ:�5{��7(B��*��K�	xȹ�U�p�{b��3��t�`m�654.ܗJ�EL����XF�xF(~M�36��b²L��[��
��x�l߈���9Q��]K4&���� "1��%i9�Co+6�U������;��`����ҕ"ؔMmâ����E��ET��ls�Q��@@�%��[30��2��R嫓p��z��m뻜�^ĪL҉Ù�Ru���y���Y���Z�Z�G-�Q^|n�db����0����������=Ux�e5�Jl:�9�B�c��Wkhb�������ٴ�b��ofKkH�Hj�J�2lǵ�F�JDQ�Ὥ�t+Y4�e�;Ƅ�-ƞ�ZQ7�>��)���x~�k0�w�)d��*�5�
�;H=��;jR5LY��(�YUq]�v:��mj��L2�6$�S��d�ǅ-��ۨ�]n[�ꭡ��n�Lb
6��ޢY�
�v�W@1Y��q�{�M�a�3oO�y�(�]+��:a����lǅc���(�Up�"��6n�`)����o��]��ӚE�5�-X���i�ї5;�1 n���n�sqj���V2�{�h���>9,�&��M����ٽ4��0��vśgdn�X�^��^5�!��X4��7�L�t�\�����Y6\.[t��9p�m�6)R�(bO ͺƍ��mڗ6�L�~BC��z��L�KP�@R��P,ōP���k��H�����q-��5�ͽc.��5�TV;�f)�ac\z���e�M�^��-С��SR����M݈VV}���8�ځͤ1�9��oN��=�7C�w��N�)�V�;u�^�VF�̠7&弰�D.��+a���Jb�-Kj�q�[f<+흌�\��t)�4�-�(}��ŷ��)H�+"1��x�V��d�c[�VŻ����1h
��wu�H�t�"$��JE�nf�Q-�r�aǮ��2V��M8�h#@vR�G0ckP��4az-���5�
�Q^��j��/)��B槈�8ơF���I��u�]�ב]@[W,��i�0���[�E�������Ь�B��.� ��t��!-�,br���-Y���`K���.�`�MM���G5GXSH�{Ff+4-[���cyF]=n�۔�)n��韴�إ��QܷQ��D�����׵��VK��(<��#�OQ��HV�:�����Se��nj;��UM�RD*�ڨ��Z�����EJs6ӄ�ءQ��� p�pX�;��q��p��i���ִ+n6h�z2����.-QnVei���r��fY��� ��[.������wI=[D۸e=��7t��xFZ���3v˫b���b��@��]�aTr�vV�2���v.mJ["Q9���q��v�m؋u6M�r�L͓Su���f��@L�����&���Z�ˣ�.�H@�S�Z�~�pEVg��,8ܻX��7.���L��-йN�ꡘ"P�,}�ygc����-Î�M�
gl��9,�5b!ʂ�$<�����I8�͛N]�<��37V�EzF+���	T &L�޽"�:�H�b�:(��z��B�B��iѻOtR1&��/�F�� "-��չ��qZ(QnZ��Y��Mh���2ه$�j�i2����o2�z��������L
�[v����
�.ҕ��� ���ϝ=u�d�r�%��:��35L-�wM����hɹ����Z{YT����d8��h&���f�4\:�m#f���+uî��O,�AxS�m8Y�\����n���U�n���,m��u��1D�B�w(;u�1y�P$PXhe�)��[���m�G.	%�S!��c�n�Чf}�N}��L��'!+�s�@����٬��mn$�5���YW�bv�Ks`,�:��,e'>�sCL��<�+knͶ��I8jf�&���NL3�ɋ	��U����*ׯ.�E1��7�������i�a�H�EhhƤ)@)�I������Zd�l`��n��[�w�jմQ��j܄ 3"B�{�a.Y..��3fv���gɴ	C>�M�m<Ҁ���uf1+s�t��ƌ�0�%kی��P5�ѼV�`�EӬ�f3mi,��Nة.�,!��3��5BR2��VG^M�BNecZ�˷i5W��;ڐ�*�%��Z�Lǌ���Ȩ`�2���T���e�b�5m#�S�b��d�y�┝D��-���4�)��2O.b�SP�9��͔�AX�l1��a�K[)@�8 �{� ��yJ�u�+U��I=�V[�b��P���U��2��L],biZҗ/�˸h�;J��Sc�-�G��	�o4�T�w[I�����4lS�+`Q�Sf�<t-��R�L&��P*ն�>&X�%+T֍;iVnV%@��됣`^M��5*zLf��;����!Gl�0����Uq�ݒ�Ҋ����؞�r�hV
�{0ݩ����J���[,�d��Խx%`,*���.�LK �
��PfU��N�G	�-��TQOb/l���G��ۖ�u���y�jc��+���8���ͨPV�ee����kf�v�B�
Sh����rb�j��*�e�IV�R�k6)Kd�@��`���4�ը��]"�%�vc˼�0�����ɂ+D���e�-,��{��jI���V^�6���.�4�0Jo4�r�Υu5����t-�(�@�D%Ӭ0���ܫ��ʎۻqڤ�hCS��	�Kj���#U�����'�+R���y�]03�z^��(fi�����;��gjiL�F7�V�
�hQ�����L �S'�z[�it ��J�f޽���p	:ɼ�Id��'op����A�޹�f� �c��6�[�j\��Y�X�/v(�;uc.�n윺�[��D )�����v�/f)�Y�oq�;Ԡ!�sP{�ݭeIJeĬ+�"��X�ɺ��u�w{�Y�֮#��r[�1����m|�.��ML�bUKj� f=emVq���V�k3J��J�ʻ�#@Rz:��Y�&��^\���V��Ju���Ă�x!��Yh퍇��5���TU�Ƀr�D��A���1&�(��{��.�m5%�:V9Wr�����f�R�e�X�gғ���& ���XN)&��[����h��T��@��2�Э�<���d�vٌe+	j��+R��Kէ�hHZR9gbV�����ul��t��V���)[�����B-x�^˕�q��Z�hB0;��K1��+K��E%=OL��A��!�yn���1�6�V��%:�R�݁i�c��۰�e���C�/�/V�0)�(:�n�	E�R�!
�����aYJ���@E�QW�{��fw~E�/*Q�P�rY	�j��j�sX�;�N����q�&fS�z����l��i:2:�5��[Z.�o�Jd�%�����x����z][�dld%�-��1����w4��7	L�����<.]�NV�X#c7-�Z-;$6hD�S��T˴EJ!��e]�Ԙ��\�)Q��Ʀ���ʂ�f�b�W���U�/$��}���w���:�soqĂ�HG���n�t�[��M�1m��X�f\��Ǖ+w8�a���[�1����n�$��$�.�h���U%G6���q�����a����Pù0L7���ل��6�r�Z�0���Ա�L�Ef��0�Z�e����P�q'�۩Ihʁ���۴H�q�F�fbn���.��k2ڤ��wQ�h�Wi�y�Zm
E]�e,�!�B�,-Z�[A�,�(�U��ӊ�;��8�&oPn��17�54%W�I�ya����l*���nTѥ.U���2q��E y��rfԭɳ7�3fŐ��uc6�7����U;L�n&����V2v�(�Ķ�LwDZ˼DK���U��*C���ӌn�T�-]�̔A���91|����8m̂Pw�^#�-F��U�J�e�2U��-�Dn�8�S��JHTP�F����`�Ƒ��B�*)�7*�β��E쑐�֛4]�&VMl%�,գCR�<���RY�x�X�̉�v�D ՔV��4r����.q��Րe�����t�+�1�f�:���p�(6[��CC,i�V%blwy[��6@�՝�Y`���7fV�Nԟ DLƒ�eCl�#QT	�j�jO(-��W�d��X��d�3k�t�Ʈ��'#j
�kfn��Q�3M�
�2k/u?�)X��Ê�Q������.;���UlI�ᵄ�y��EQw�}�ڴb��.�E@$��$ ���7R����@��^��d�f��{W�ec�3h��Y�������-�rAY[�]��Z���Z �Gk-e�霫j��dMͫ��Ż���#����8�n��ݟ<�T�P�\j��-;����ۦY�T۳�2�;%�@���M�blQ:�I�p�����7-ۣ�eY��d�����i��?�Q
�Ѽ4��0v�	�y	l�FP�H�X��J,ʰ��ؔ�����3k	eiM�#@�v��$vT9�\�0Qi�R���.E���C�=_&h��(�s�Z˅�tn�dǃc
��c36�*}t*$N���[-R�Te�e��;-o�`*��u��,<N�u�n�	��T�~�)R����/�wJS�����q����"�0�ib�v��S-��5n���w����tіS�)��u!Y��홺��n���O ��̆bH�(�o61���	[��1�4��`VBm���[wP<���GX���[5�F���V�U��#,����A�]�EJ�f0���tQ �E�5��.(*�8�K^e�&V�B�K9A�r��L�iH<��%��ˀ�˺EٲU�0�A�I�� f�m6�!����Y���[c�]l�&�.<-꼤�		� 
���F�p���"�ѭV�&O�FLOL7u+�f���j�
��l����*
�n�YF�r�2�F��ۦ�^�*�4bʺ�D�3E6�\jnTĄ��X�˦A�%T��B�g-�S�Q�ݷ���@T��tE�[i8�xt�r���d�Š��t�j����4����A-С��D���%l@�4d
�7m�����6���LKU��p Q�� wN�Df:;$�"�c6��y�˨�/6POb�6�}�U��,�zv�
({*��J�i!�f��y>қt��wL���fL��U��ȝ훣&��Xw\�c�YV�%Ҷ�։�̻@��!��K��"v@�d��Z���Ԃ�TZ�ڰ�ӈ�z,G�,��	��Q���~���Z��Tu��X1̐���*�ݎH��P�����J�����3�4��LAW��ܠL�6���,�y���v�V[�hf��h�%1�iloRݗgQ��6�W�-"�|��K������.��Jق�<C�q�D��/$��NnE+!S��;���D����uC�%�ީWu+�K�b�6��v0�iJ��l��d���!��b��vݢ��jtn�-� ٔfmӢ���1�Y4j�����$�l�7i��,ˀ������ͩn��2ap��.4*��ɕ��9�{,L��(��e=_L�R�t1��EQ�Dۇ��)��S�w+++��ګ��jƥ�����ǩK���J,2���hݽǅ��m�0`��o^S��wjR�/��b�٬�kvY.���d��5-�i{kCq��η�طƵ.Ǖ�Xy��a�+$0*�4@b����Ғ鉦��GT�mU����V�4%�8�Q�cTU�	ZB� �kN�1����5����+ݍV<Klub� ��`��f�B�.$���%��cKb[�l; 2� "a"�VZ�*��8kq�[�N�G(�J���m�z��۰͔dwp;�$ֆN�OZ���e���t���z��Y��+����d�I�t�2)�չ��>�� �,���(����z�"ن�
e'@e�x��";�񵡼v��SӔT.��0�ф�9Scv��r����D;��R�e�s1��	?�Q�������[�tuT
^�V��Bgk0;���m�� ���)�n�WLK�у-]h��;��6�l���/.�h����Un�$}�ʕ)�a;�\���C��W[�+]��U�c:�,���r7"��X���4�)���+��j�߭�|�
�˙�,s��:�EՑ��՘��b�]��}���Z�{պ���B<�m/h,�"������]2���Օ�_SH	u�(��īw+��;R��9_�N�ioe��ϱ-4�1��@��6�82��X��juλmE�귯^�Ml7�28��t������[���\	�������%0x*5tHY�3e,D���ͩ�z�\zW;��Fet��O��0��O�����D�5mn@���^Θ� �]�.NOO:���
���ɵ���JpZv�n�Z�á�Λk�\^.�o;��Ao��W����'��Q�Uq���OcmŦ�\-�^8� ^SR��֥��G+Vk��خ�v�Љ�HՊ5�T�?%].��Lv����/SX�cz8l�خ�쩙�ʙ��4��&(6��(L/&��N�4^�]����d�fu��
��5w��É�V�\��<�A�n�Ő�߼VY���4�C{dOjH8�=�w�g��*C�aں���ݧ)�����(�	@��9es~���O�x����Q�wR�=�,)V����oJD��1Cm���d��ѥ�x��+D+�������T���n�:��3�f���'g^!��o����E��^�� %:�w;(�}�����(2#bm*B+�9Z��ۋ����2Eێ��r�]z�YK3n�"uΚ�xu�=ܚ[o�c���`����ݯF�hn�f
M����*
���$�e�q �<R�h�;7+�t1Ђ �N��GE>l�R!׶��`����ou.}�*�f#n1./5>M�ī���+Z����.j�Σ�r��%�����S��k�`#����9F���m&��U#t]��[�b촤c/j��Ⱦ�7]�}����q���0[<6�Cs{H����RN��ف�%��7M2��oݽ�T̔^�����}��iLm꫇�=���f<����ﲂ���g}�]iq���]v�ܐ�����d::ͺ
��[σ�W^��]�E�ƌ����َ���Bcn�����8�ge�4�*աbr�Z�Y�I�&�-�޶�_d��G���U�N�Υ��:�ԁ$�yR�wT��A��kX/����[����zD��U�5��k|�򓔫�����dn�9�,g�7^�֡�Q`ro
�����o�d]���ie݅2���B���XŒe��4�;�>S�l-�E������b�{�<�9Fbv��74�u��F�TV���9Ѯ��:�sH��׶�T�;�����|As:}��n�2��)L55�\�B�EA_L�8"��r/l�Α�opS���J��	vhڻ�x'J�GuԔ�W+�%fJ���2��:����`�3]B&#��/����y���b�ISb��t��E�Xgi�����W�M(m�A�S��2����8-31P��>Z�,g.�:��5�}�k�h��o
�d�1�uq�,��mᚁ�V�ml�-��g�Y�]������+$�GMX:�Wm,y]����Z�.JE��JJI��hZ��<%6�f�-�U��)��\���y|0/����S�)�2�*��w ��˳d��v��C04���/E>�W�dcm
���X򐥳]B[�+y6���u��*�ﯷh��z�bt����)$����c�>-l�֛IlP��C���F�],�s��@&�tN�qH���v��ɔ�3��2��Y|�e]A}N�^
ɍ�H�a��:un*�[(g3�Mm�v�:�Pw\����ly���Ո_y%�)k�W�.���`��.R�W�5$��5���->���Okw���+%�s���R��.����vc��1d��YS��Gu�<h.0�s�J��t9�H����>YV5�[$w8ӻ(e엏/��m9'SA�JfYh�Zγ;7:
r��S��^Bre�9��.l �E� ��RﳬtY�G�e��%8��]��˼F�'o�N���934�F��D-��[��䴁�R4�^mi*S$�f`؝Ǥ�ٜ�]��B���Ha�,F� ��Vِ�IL( ��a{�V���ǃi7�����{����C+Z����:���9��&.��,�m�E�&��H]>�hn��4�m�7��d�օOU���f����>�k��F��2�&�^�a[Z������R�Ǩ����r�0��<�>i�\^+�C�&�[۾��� k��bt.�`�t.Gz��T6�ɞ��Uԧ\�lZݗ�fvKhI׮�F;�[����+;��t�ˊ��o���RG�@�����������qq6Qŏ��c�C��g[O��d�g��GP*L�:���]���-0"����|�	�=��>�/ǘ��"wý�X��Δb�}���
v����W��ش��|hnNV�}�];
�2+G���W4�����[�4.���3�5�oڨ��$���P��9dØ����kI��yʽR�.�f��;[W��Д���`���O��5 p�+��)�1u*Nh\��J���`��9��us9]�$�Q]W[��b�4��\�)\t�>/:�S���^�kc
.�5���8�*���)9���(�*�����N0,�uyu�a�&�v<t�aZ{����<�8u����l�\xu��E�T�U�|�aZ�r�;
�d.|]�T��Y�Ī�f���ͽ�b��'z����h͗�aH]�A������Mj��؝�/3�7��;;:��]I�6���參KdU�WG��e�2R�
��L��tn�)���k0,��_rN�ʋ||��Y����~�8J3�VF����8�CD3�[���Ty�M��ݍ�u�o���v�*�N�%�HC�I�9����1���D����הw�lZ��Օ��3��b"�B2����߅u�s�mc5l�*�M��R:ļ�Xm�����S�A�@p�Ѽ�}�6�*�Z���W�P4���b@�s��� 3�r��o)F���,2�@U�r{���eU�+�_҂dhS.0ƣ3��p��u=d����9 ry�P7��]�G�8�����n>��7�k�%һFL�*i��O$�F���3%��a��-79+�Y��M^ǣ ��+���N�A1B�ݞ�o�f�
��T����M����m�2���X��bT8A9Z����t͊A��J�ykv���3;.�<Y�Q�F�r.)Vs!��M8��0�m���V�F��a���-m� x���V�뱵�d��̉�U)��YW\P"���A��KSi݋/�+*����.�˜5s��'�Os7��F
�P%�<%��,L�qu�"�ҙ'2����6.G7�����V����άT��ZvZ�d�ͧҷ����1,�m�!�ըqT��j�K���9��5��iT?7��g�wob�N�)Cӹ4����O5�cj�[l#��Mu,Ad�Vs),���7���%ĩ^�A�qp��-�'�T>��&��:�e�!x�N��{�I�*p}�F�)�d�!����B�H��]u�'it�	���U�Z]٪]���9A�����Oy��A�ǏE+��͵�ȂUj�w����!o����g�Ƴu%A���ɑ��UԻ�X�v��]K���]��l�h;:s��]4�j���(z++)v^��M2R��7Ƚ�Yڹ
1IQ��:bs^��򤑤�ϳ;e^����N�'}����3����V�ʺ�qs�f-r��ݧ1q���c�(�Ac����3��*й���%+bˑ-w�y��4����oe�gc}c��lq��Vq�:��9W�FV'92v��˾���	w��!�[��D+�������1SgN+�|y㸛w�̚��b]=��<{6��wʤ;�)�D��b�(���ލ���9d�7.wJ�ذf8q���NK���]�,��[Z�U7��h
��3�����W��t��[��Őr��;o�Uy�rhʭE����V5{�f
iWХ�ܳm�\��o���bJ1Al��ÕbsB̹��^��u�=r)V�lZ�oMe���܄�|U>�Q�<�[������	��Z{�'x�N�S[�veq�܋!y��E�.�Y���_��o1]�Օ�4^�]0r�e�\��T�͠�1o�*x�> 廦׏�2�z�Q��#��'���HV�oj�J�X�ݵ��e�6i�7^1y�����yJ�B��h='�I�u{v�y�g4���-��\�wz�J�j��d"zk7B�����oɚ.>$�m8�tᩝ�6�Q�%w���a��1�O(j����n���qsu�>��
�{Ӆ�VU�L����|�P\�� �f����ǧ��a�����Eu�xn�-#��
�Lݦ��F���Rc��ma�=�FA3�4�٠����(.��٦�pޑbܭd'I���.ق�C�W:�4e��E�z�@8t�q�el���r���O*!!�,ź�����ln��L%��5+zeiz�T�e�Zm�_,�9��
N�ಸ��8.��*���<�nP��LV�ܤnըo0QC��k�uz��N��e<���w)��
��O�g(���@.��lG�%&���|;@�(�yȋ��F��m��9O�c�g%��C�kl��{5�w@�8gn8h�,�{~�O^yVҽ�`[d�`�{���I=��(��
�m�UƲJΪ"効Q�T\u�yg�[�"r��/)��u�k��Ric�4Ԭ��9g���;h�w�N�F�3�FU��;�1Lj�rs��c�`q���� �=%M�"��}��=׵&�=�t�����om�5�5גBtC]�.=���N;]��1�����BK�U��A��܋����,/]n"�,h��Х���u�6v��Q���i�E��7��}OE�Fؑ
����g5"�3��Y������<{x(������ 3��Ѹ�b�p�f�Q��g�[0N�\#%�zk�bwh���q�[��+"]�y�x�8��ɏY+Qr�f�c6'{aoN�u�J�d�ہY��j���B��ʴ\+1t�
X4�W�l��w���Ϋ}�RH�R�]�hfoSKwWV-��4ƕ�8��`�|-*LJ4�����6�g:��%�D�*X�yċ<�η(��.*�UB6� �u�9����N���E�w@n�"6qm��X�:�����֐\���r�jb��L�o*c�k���+][;X�0R����0�-�Y��S&�O(}�gp42pwA��7FqYKL�{ӓ���G1���e#�䚳[O6�8bxq�4R�}· �M�u�F�*�	�����*�֙��{E��̮���F�kE��EVp���N�)��Ŗ%*A�ٳ���n��k�)�6�#���)�Јy҉�K�T��m)����;�5�w����9���dnu���#T�ٶ�:㥂	f�f��������׈�n��niTh%/`I���@��9�X�&W������O*+x���ǚ�Ʀ�^�^Fa�yZ�ՋZ�<���]b�[�s�R��M��S����u����fIᡷ��@COT��^o1@<��U������YG�7eq���P�6:���+������p���؎on���kj�s�MU��x�� ��G��-���ZYd�&�J�ճ�q`�b�}vT�����WS�j��*h�
��uFl�V�Rm��NO�|p�pg[WX��`4�a�`�V���{ʳG"3[�m��z�D��Tq����Y]�6������@7ǣ������{j�c�`F�����r�>S7�/v�yJ�|�n���2�d�����/�}���&E5v5��mk���ĸV�-v�o8��n��[�6���i��W\������J���|)�C}���Y �+�.`]��&����ݓ�+�'�3�(�l�v�]�AD2�q[��䆷��W�Ժ��z��z`���5;N���9�Mg�;�
Uy|o��� n�DGO]#�㽔���mՕ�Y5Z��r�#-�����!��9���l��0���3{�l=��i�={}[�v0n�Ά�R�c쓛����Bv�R���G2 �Qa��wϻ������&��S��!3Cz��Nb�b�ڱ�\1Ps���]�{*�픬(óL��T��"�27��_�ϤN���s��J8�>m�9vz陏RBmO
ȴ�{T�*�c1�N���_S���Gt��˃�E��Nm=:��ٜÒ���u>��[s�o�F�0U��c{ޥ�îU�Z�y�c�E�fĸY'�T���-�6'v@iS���y6�T=��$�s9:����/����b�_)�z�\ZN��@��,v@}��[3��_�+��;�iN k�vuN������HJ�=�u	��o��5��5<8�e�8�F�Bj�o��'��݇�It� ��N��հ�uaL����.����o�����Wڦ��z��}ȅ���x�+�Gh䩝�sw�X�\�Ɉ�X�α�"����(n�Ō٪���m���%y�~2�Q�-�j�2�d8��kD�6�-����tkU.6��r���2�/Wf��];]��&��uy�����|j���m\v�u�벵����Uu,ٖ�^����p��]��D,:�xAA����-E�oP]��yB�o`O�9�d[x�-7�����L�e��:�I��A�Ȕ�����ۄ���IiIHRKU�R���)OJ�!"��J�̅�mūT�%�qb�K��*V�[�iy�8+)I�	JT��jի���ԑ����ң!v�7���P�I!�+Z�17y���� �	!I�}���o����WK����xR
�r��;�؟S�N��`;SUc̛�C������5]`0
��<�J��$�*k��]w�Ɏ��q_�A5!�۹�d����\�E�ei8wqY�B���]�xrv3/z`ɸ7�W���cp^�Z�ߺW���d�p]Jt#|#����(���cC��;��=b����Iv7(��ٸ�՛=Z�5�oS\�L�m|wa�1V�m�g�m�h%f�2���I�%zib"u���PW5�6��Y :�3F��*^/9�H�"�E&8�"�i"`�1Xz�nV�[wn����\����H36m B[f��{Cw]Յ���=��X.LC�MHeB�q��1�
�uLu6qs l�`����R:������Z7Fl���ʫ�I�o��sy��ʖ��&��[���U�%ݫ�1u�9�賡�5>����n��)��Cis�{�ץ�hb�H-nf&^����ţheZT�M��z���d�b�
K2s�[,dF��;��{�gN�Mm��lu4t���<�mr�U�*��J�u]ZK�/��5��l�\�s%��˾�(V�KQЕm��3��8�v�tؕm��iΰ89���8cMrxpˬRSǼ�u�̬[��v��A
�B[yρ��`.3yw>��WN �3��]S��k��&�L��.�lR�_ ��?w��S��%��ّ;ܫ�S] �J�EG:Tx���`��ë����Ԩ�U�J��J��ݸ/U�7V;!]O�=�)嗼 D�8�w]5�m�d��K ��G�	��n�9v�U��YY�q�V�18]��9��Y����C{<tf��ޕ��0�l��E�y��s�RE���:ʘz����O���_>�171f֢\EL%�ߞ��Yb��
I��s�`�������O8J��\֗�`m���\��]2�9�/�W���(SݮSъ�ʢ�o��,�VE�T�UJAg��C#�V�m��qY�� ,�|�jH@�/;Z,����yV[Ȉk���N���=�i`�˵l�AT0Sժu/�ĩ29�]�;=ɬ�3*K!�"��뀛��s��s�����a!���ăC��m�{�
�ɣ�L�b2���[�>'�w����%�B��I����Y0�P�S:�o+W��̈��D��
t�1W,6��jg�m��1��Xuꣶ������fr�+`Bu��#�.w[�]7:#,���Ǵ�U��I_p:��7HSj�E
��Â]��+wi��KΛ-pD���JOl;�rl��&3AmK��U�X�;,M�2T�V���<{m�s͛B�����#�|�2^QTqm^+�#�Ek���m�qWW[oB��\�T�
�>[�s��z���;G;U�w��֍h����Kkn����ƲdԀ�d!]�m!�$���A���b��Xl�tѤ�\��U)�5ʭ	;�厰�tۼA<[�\�Ђ�-5ǫm�\P�nV)�`G�T�2��0u��Z���7dV>8�V�MɈ�<A�]cx����Me�-bL�nWge:�
-���` ���X�Id���nd��&D1�"�JX�b�+~��k�ۘ�5�"�e���FC�Y�؝ �s�{Vּ��z���cW��Ⱥ��xw��ʥM������K�Qr�����%��:�KT��2�{���Z_9�˃����<�ΐ��lMU.������up�'8,����B��Y��`����sa����_EC��P��[=�Q����e�@�!v��sWP-��MZ�ur0���|1̒���: T���Qu���@��:��ـ�d�4�Ylm;�$�F�Fk7���i[��p�JŞ�����'׉��ȝ�r�����-=�\D;�q���1�9Y�]:��o����Fq�vNa��@Eo79��f�.�Xҡ(�����Y	�0 ]�K�������+��<{ftv�.m٠2�
�LG�4�I�J�Y7��n����V:k[Ps��wl��m�J�����;}R�v������/z�T�0���ʒ���Ǩg`K��/�.��pvH�'�L�Ǜ*n)Q�Q����,}����V�Q����ƶ��׎,�_g���RŸ_)Ë̍�J��K޵-J���+�S\s-r�z�vE�]��w� �}�ݷp��Wڭ���UK�",�m�X��IP�?5g���{ �^*݋Xp�;��^Dyc�*�]����9�:��N;�:�ʛy���As�T�ltlALܾ�j�9� a��
��t��L�^TꏲS)�إ`�H�[43���˿�Ŵyuɕ)��2a�;unk���vZ�U��{��� :��tS��1I�=�/�3@�S�1��}�]v�����Z��qVB�����Z]�ur�#5���(��cU�*/q�ED�3/�+��(;�Cl�X�	q��=o��4��5���.!����U<�9�CY��+*uG�2����U�'�`Q�52�]���X;�5]�Y�l��d�=}�7�B�5.P{6��Ři�E2����j[]W�p��*�y�o��� �8*4��l���yn���:�ճeNKQ�� ���D�n�qG����4�V�W�Vpn��їZwCX+���[S�㜻��"�ͬw,>���ެ��6
��}z'��u��W`f�Nd�
��p�P��N��c+q5���I[��fWe�ۂ��:�Z�7^�o(5�-A@���`�� l�nX�e������ˢ��1
��۹ū���J�չ%��QI�j��vu[��qo`��%ee�IK�&ct���Q�{�����R�)���f�$�nC�R�2dy	��`�����[ٽ��*Bzؙmn�n�="���������e��k.J	�K��q7ô� �ʻr��m�b�*�m\�|U�kB��Mܦ-�EF�p�څ���.��:A5�RR[�z%X4P�Y[��Ab�-r+jvՋ�����`n�3pV�d5P��k���(#�:�L�V 鯴�qX''w�3�K� �GN�R�ラ��%��0&�%LpY9m�U���m��T6��Q�)) =�YM��]d���.��M��u�r��F��[���uL�01��ڹ8V����0�cr��u*�&�m���yХ]3�ih=ձ����苤�F��^Wen>��[#o��ע�2p���{��fT��\p�·1�,�w�^�I��N�H#ꅳ���}�֣�
్�<�nP`��.���cE����AZ,�'Z2Gγ�(L���YA�Ѽ[
�V컄�P/�-P�o;s0=��3�"��8h����I��XN"3����eV36�1@��Gp�:�G,�q�z��.�ق�s�M�.��7M��m9����P�4[�ׯ��s���lr�(%\e͑�� 
�m��I�z ��TD]�����+Y����Pi�gt�������T�^sC��`����o�[7^`x>�Ll�Bu0�ڐT�Vt�sA�@|�8���J��j�.zgP�R�6������<)O�����ƪ��nΓ!���VD�`F�̫�s{'hzb��(�Y�	�)d�n�;�Q�Ŏ�6z-u��z�[ ���s� ����Sp[F�C��ڻl���gk�8/��`t1%����<�\�+�֫��M���
�݊��d���b5l^'t���{J�\�cn�qÅmJ:���u�:�"�L�9�]n�uu.V9ŊG����͜Ҩ��] ]��!��+��Ɋ�u:���B��mK�
��A�S��!��ٔ4R���1�&5�F-gLѼ��l(ք�]0 4,)�:@�R7�]�Z�9����& jR���d^.�F�֑U�1��V�Ε�/��ss�;:�Y_�׭���r���'���Yj��`�[Ĝ�v�#�E�te^���0f�R*&%
i��]�ը�c �%c�']+�-]��\TH�ީ2Y����nEz�9 �6���sUEV�]���yԐ����G6����[��k�!�-H�}�U�{���]�=yS�����o6�ͼI�豉��N�b.Q�W�Ʒqr�'+��r�_,�c�k�x�d�+Ai������ȫ��r=W���^*Y91�κ�L�0iD]��#��D������؝�Q5�=|'b�Vf�����a�O��i��n�]�cBM��I�Fy�����W}������j�]+D�r��3���:�$.Ҋea�쏣}�>\�Y���Ӹ�O��J���5���uh�]��W��,JoNcA���)�n-wK���s1�զ���q��I��/l[��馮���5&_`dM�}Ykh�7��rՒ��f�\K��1�{SI���y�ap�*ā�x����{|��OGVn��fþ�e���3
u�nC�t�yYD%]} �в��ڶ��?�E��/�\����ІfJ�iD�.�Vl����Kr�e��N��	�M��զ�6�yqc��9�ӑw������-��v"��ѡ�KE`�.�2���F�j�	}�޴��or�H˛�uS�&
khf#pl�9�Z��]�̓(J<�I[����l
²�Q�"CVjY܋�ʽAS3�&�a���?��Y]���>��X��E��.WN�]öR�3XVEʆ�`L�.={�����+f�v�)G�{̷�[榬h�9���ܮ�%bĩJP,�q��r���3�G�u�J=���2�"���	��Ѯ��Z|wN�n�򻖉����Z
��;r|ѭVZ��+Zp��8�>�1b���n�:�;t����i�k�e�X�L�01+�m�I�Öt��Ӿ���k7�EZ^i�V�Mu�Z�5��zc���P��k4w-ĳt��eomUf����~�^RXy	.T�2��[uҢHh��{A�[��V�&w-���m�p�*�����c)e��z���5�8�r�"�A��X5|�r�z�Tּ��򭗊�pf����:H �u�2��qӺ+� �;��(T*���g\�&���'>El��W.̇������j�W�#�27u*wh�!9�.���N���`V���؛�]B�n���B4����6��|�M���Έ�P�Qe�zʉ�xt�w5��Z�T#|��ծ��Ք���B5[�/�%+�y˴'.����V�c0�^r�=��e�0����9��.�o����O�h��ܚh����]\��^�to5Z��
�l;�t�&�q��2�0a�ͣ؊/{kY�#��q��wb���1b�+5A������]�e�����é�
7|'1�����:u	��]C����x�w-[*a����A�L�U���ED3\ླྀ����vѬ�v�k�B�Z�8kz�(P�q'�Vi���b�RTG���3�6����{��4ԏ\7��%
��*;�n�A;k��9E�=bh��{�bze�i3A9Zj��3q�lb\��gZ���\T���[p:whr�{�87Ѹ ��a�G|��dmq��9E��wue���F]������̈�'�C�,<E�<���P}�]ui}��'F�ZM�3�9����yT� ;��'-v]��of����t�t�3�N4�c�(���wt�ϖ	ن�l�)��b�}�oX��îK�(|�(�ݝԪ�o
���մ��EJ
q��PJ�ؠX�j� u��B�!�5�������+�:��b1�pt�H�^*��H� �j��|��շَ����ݹcV!�N_(IF@h^J7�Eݩs7�]A伢;�Z\֗U���W�c�p�[l���[�l�Ü��o�c�Ҩ��Q ��
�fw��3�<���g�p�!�`�u�9&jR
�N@�Z�[E^ט����ݍj-K�U�f2��s�Z�,ޱmKz:�T��!ky�G[�2��ݹ��J<f��Y:�nS �����ei�h�%���NI�G��]�1[}R�}y����Գ�:�r��:*4_P�y�%�7md.��w;�y�s������Q��cJ�t�(���fa��l�b�]ԻM%4r��F �V�Tό�O,�k�탶Ԩ����R	CҟA9�\��� �l)�5ْ�S�h��i�vwk@��++:�������\
/�R�	���
2��_oD���àQ|�������	nh"@�:�&��� �%�a���|�h���'_+��~�\	##�]��j����za3y���R��jL��tw,嬓Ҹ	�m�n�ӂd����7�ɯk'vE��(jx8��Cw�j�M�#׷s@�ܝ�:���������*n)6��Z9��D��y��
�[���ָ����^�.����;����i��pZ�e���,� �/Y�r��oi!D`����}[vf�v�5�+��K#�\�G��/O'Qv&�s,t�Lc��x�E�.�u{s6��N�{D�XT��]q@u�S�/jm�b�-�5MS"���jOn�MU��]��jVS�ԯ%��U��V�i�C-�i�ĐO+[(v���Y�>�����X�]�u�;M.�B�"�g5�Ȉ��Ζ�+"J6N���͙4����i�iWj��Ԇ�ښ�na";�������O(���hm�>�F�rי�����چr˸����_IR��r��4f�Ǐ�ẺJjy��ھ��N���M�1ڙF:������;�ԙ]MS�ϯh�5h2md���d�S�b��4�,-H'���H�4�>8�Μ��K�Y��7� \���k�Dlkx�X��i�H�����b���yϲ�;�J�r[�j��d�Wem�s+�+�X����Z�t���$�C�Z��lڦ(V=B
�4B�VUoeA���ɿ�������^�K#1<���VhV����QZ~<�H��K����R�1��U#�L>y&�Fsr��LNln�[��ql!�,8+V��K��Wk��%J�㾭�J����.�Ӑ ��q�#�����%F����ח6�*c�$�a�JX#��u^�=CڕچO�}�U9^���sS:��.8�
/Q���ĩ؛�����S���k��D
�2k�4���>���ddȕI�%.s-��u�����ZO(�e�&�.�չY�o����;Ƙ[����e[�P1\������Yta�u�4�[��(
�(�R�FF��z1S�Y��z�\_�&@�����5a�N���/%Cur��Y��]�U,\ٔ�A��zw��|�!�ͩۋ���|W���}j0Km�Q�%w�vfJ�x��2����e�]�\CTW�i_,��r��n�)C���gfq�5غ3�ח�+�`	I�s�%L�ެb���Ƴ��N*[h��]ܪ�����S��w�O ��t�i���vN��Jh<�Kze����f[p��n��[D��<g�i@�U�*��VC��f���b
Yy\oUuМǥJ��+)/rba�������tPܮm=x��os�ه9���{P�5�`_<
�ׯ�<"+�3;�V Q�;C��V�ו�^�ԍe�uy����R�3��������p�¨P˺,J�V1�|PT���pJ�k�at��k��ޤYHg�O(��̺���f�Q��@�g�G�[9Ӷ�V�
�U:/z��P�m�~>>����5�ڪ��E�Z��Z���*��P�iU偋QL�F`����X�DF0Tb�0X�e�Ub(�mX��0F"�
ZQr�q*0EJ���*(�",+R���X�1P��Т
�DU�QE�e��Z�$Dj��"�LlQ+bTiX�QEJQ-+�*UUEի�T�T5J
��X6�1�@TQ+)Z*�)YSv�X�UUB��iiZ4TU��F6��*�T���n�"�i�+TPT���F��aAQ�E���Čm*�k��A�%++-�
1#e��X%��V[X�����,J�E���֊���j2��V6���6���-��e�`�PUf�j�\�U�+���D[iVňcFұDD�"���QUr؈��QEE��4�em��Ķ�\e���2�*Ŵ�Ub�j���TEm��X�[EE���#YE�(�v�c���ŕ��Q�V�QUKj*Ŋ�l\*�J�PU�#lZ4e*Rm�h��U�[UdU�mE�clR����")��aZ�1&
�UQ[j(,+U��UПU�n�M1�m��-`�,���'3���Lj�v���ۏ�+��΍O^+ǝ���+q�spWu�oV�����Ϩ��%h�S�x��:����v�a�|��z�e��"�9ʰ��|L;�IQ�In�¶2�D'yz��N�}MT
��Zf���:Z1�����(�y�R�'`9��k�g�'9�~�N�u�`Sf�W�0ؖ��s�@='�n��{{W5�Ԭ���5�{,:�<0#[w���&�vt˘�3{�w%�V�}y��	u�^��&_D�)�Ҽ�����8��N�\��4����A��pw��B���m��6���N��;՜�t�;��j������[G���g�u�|n
`���Ǆ��ȵy�t��/s!�,�0���u��c��s<��^����n�PC5Њ��$��
�3W��Ǵ���;S,z���V��r+��;�im͆��ɰ��
�륣�d����}O�淮���hVjf�[�~�|�g�o;��m�\�-��M��ՊCtɮAw0�Ui!z�q�w�֙IԼ�
5"��7���p'y�3;����,�mc�����mO=�׶�2}iD-?�Y��j�5r뎳d���w:e�i���d�v8Fa" k��3�}7^%N�w�G�踘��1�,f�B@��͍H�Uζuj�S�uȗk⍝O{2h+�جq�u��>�6E&z�Č�z�Kq��Q�2%6V*�ی�aGv�o"��-��;+��Tj�E��3���BR�\O�����D��m����~Qݲ��J,>�#F�q�C���}��Kg���gD�G���+t%��>���=�c���^R��#�g��wjr'eR�IA�Z���Y5U*�9i���BBN�_Lv�(g���Լ��!$���k���8ӟCN���!܎][M؞��
�V�)�1���@P9w�����O�H=c�����g�+c,JʢԊ��V�T�:�w�Pw���H��m��޼�G9�i���fa	��liv'�ȕ�>�������v�>U�m��}X�h�x���N�y��hN'Є��b�ӓ�����L1��X�=j���P���ZQQ�G)��&r�l]�Ǚ�d��q�9ug�o�'��^gHmojy�_��lqT�5�
k��]�ގ�B���q#����l�9y��;DnV������x�n��:X|d�we�ƻ9>��
���� �+�ԏ3T��D�z�r�zav�H�ṛw�:�M��k|�܃��3ê���g�Y�jaW�vZqrwɘSp��u��d�<OI�yw��-��Xo2[�o.\�"BOF�sX8��SU����7ӭ�ި���(M��or�
�lP��@k���K�b�(6ԍ���N�L��y8�G�I�L��GTz��Yi�珯���12V[�p�s�^�^S�Y��ܷ��ρ��S��"��(M�ft�j�Uhb*��+z�f����U��k9VW�-����7���:7z�x..��.�1fs\���y�)�j�s�J��{c�]o^��HX��wW���4Y�ZjL�ړ|v��->���=���n��t�Né��Ĕ9���l�D3'kuw:U�*�[2_��.��)����|��y����\�:����;wT?z�r���@�}��Y5���\�<j���su�B�c/fv����s�$����\�q�#�E���8!I	����Im^A>�ĉU[�oFn��>�=}]���}xc�+K�h���m��PW6�����9�d�����l��\�;�1��Ӗ��S=��Ơ>�����VpD,��V�W��ܺIun��ġ���:�$ص���a�zl
�M�~t���x�E�-����I����j����U
��`�O T�g�ا`!��V���T&��}��}|�j����Rʽx��{���6w T�a	K&�*Cz���H�ȴ6��9>��X�ÕB�9	���	��Ѹ4����[�Diȁ~��umu�'�T\q�ʝV#o(Jq>���Rދ�'��LDY������N]kL�2�]���c�C�ԟ��<��|�u$}���S�c#��;��o�[)T��;�2l>&=����������w0a��M�hS��;3�f��
��](���<��vN-7>zZ�s~�2��{*V'��ݎ�汹�4�����W��2���|*�~� V�	�a�9
+�x��l=(X�CS�:n�����ߣ�<C�^�c�A�	�|G�����>sxW=��o���#���ю��Hg`qD>w{+��9�w�\9VS���nd��-nfq"�\�D6`�6u}��R�)�Μ�Ut����\�F���t�L�4ue�����2OPFn.�F��nPJ��~�9>�U���)�X��N�i��V6&��<go���uk/'y>��my����",�d�2��IKcg�xCq��>b޻��]^6��.2%�N���Ev
��]3~�ݛ)��6-�K��k�����&-�d�n��G�/)lp���l���(��[g&�Ơ���6��:�n����;������xB��AQ���Q�^����$���⯵���<]Z�>Jnv���z�s͈j�\Ⱥ���̮�ୁz��ѐ�p�"���s��pdkl8��l��e�l���G�����P��eR��q�2�+S9\iP�|���/A�qjNqҼP��Z�|n7
><+����q[K2�:f#�_�P��`;��ϵ�����	�'G3f�0ܡ�Y�1�����Pg���Q�3�o�MO�q�u���- �����4f�u9�6K�K�K��I���F]�|6���墢��Ϲ��C�B�C�8��o#S5�v��j�dݡ�Jw$iLV�u�m%�*�����pg�0�ؚ�:�ѷ��`�IHK�5�;�޵[�w=O��6P�
;JO�n��`r�����4�*�y59�n���i!�ل�9?jy��}��}���s�s�٠�6�a��Nͧ�SV�=��ՉɟV��`մ12¤��Ǜy �fQ�~��C_��rL�&�IZ�b���~�U/�^w]��r'-���bf�v�һ!e<N���˺f�[�9�ʹ��Cf�=���m�K��Gm��^�ĺj���gN��\{�5p��-�x��b;'��+��,TcԞ�s\��3/�9�ƚy;;�V�3����J9W��k�O<�}��u<֡~�w g[�b���A�޴��}�3��#������I������Ն��],��9؞u�)'sb�TpL,qY=)-N���P���c��O}���ګ���R9��c�oҔz(G-�� ��0[˛�uF;4�w{�f��!�)�Y읡=ؖv����'-Vm':��%��ˀ��ݐ<,��k<�foyt1w	ʬ����;���]_:C�Y_T�P�ĳ2Aܦ�[l�s�s�&���:�һ	�d�"�@�ͺ3^�|4�]f�ڣ�b��ҥ�j�
'/jRx$�kw��ә�3����9R�2�+*�U�q�Z�ʎ���⹪$��ρ7��y�S�)��%W�]�9
��9-�B(��~3�ϓ<��'�?^�T��aP<�P	��i2P�G�r�Ӓ�Xy;����Pa�i�z���fR&50�tp4n�q!NC��wp�Wx��s�r�;��*��f}��[��(P�/�	<4ѻ�1g{ɇ'���mB���1(�:/꼛yW-�B[b��k�*N��N%5N�u�.9��j��X�&�1�m��ٻyBn���	��pF��ay��7�pc~-���)�`���U�'�k���Q�OT�;��3��V��Q��_�[�|��+��ջ6�Sb��M�zzt�G'��ʵ9�](0�5ۢR�q�^��������\'�)������g�jB�� �E����>[��Y����y�Z��n$��V�Z��V��l���U����x��$�ا���f�ҥz�t��&��y��v�HY�Wgv�i'ҤJ!mև�Z�g�2-+w�ӧ<���ٽIBk9���G�wAS�vp�r���:�bEDE>�=P���TbW�p�Q�Y3�'
�3aO��k/x/V��j��xS��r�T-�e|=����ڻ�p������Gt����w7�T+�C3��m��߁YT*�jd(1[�MskV���p����c����5P(6��?:i�9��q�̝L�w݊b��å{�m��c;6�ҵסSM͍�@�)�<Ճ���n�߯9S܁Q��5�W�γ�K���}\qװ9�xf5�j`���p���áT��U��ؽ���/�kܗJ��s�ɍ�N��S(����Z�W��w�*r��F�Bq����rݍ����ܳ"-�7<���G�t�bqc� �k��޹F��K���"��Q|j��*��뾚/���R�xA-nq�����x�����zv%���UF���N��o����J���
��r�2�:Yfج��V�_S}v1E��W�Lr�0����_i����<[��C�(���yg�9հg�Z��3L�4��b���W��5�y�Ω��w��������*�X�)�5ՕnS�.�8R�)�C-�C��j���6�sg=�aID�{�}����pq�$���[���!b�����ʶ�kz�b��gZ�;|-��������V��Ldeh����&df�h*�^�׶�\�]t�1t�<dt����&��`�n�l���\ؽ���^�٤6DRg�#��MԽ���ʌ�Kp��o)��@*k�ǲ��u��ˎ+Nۮ�6,p���J�Rբ���]j�9	�v�r�ؐ�N��л���ɼ���F�PR�IY��=
f���o˫��|}�<��zה��t>�t�Go�&;k��s]E;�f�
�<&��^��g+�=�9��k+��^�\Z�zW[���.�p�^N�9k�'a�VlL�ŏB�u�6VD�`�F�llK�Ԇ��+��]�2JՖn�v��˚�rD�.�%��O%'��R�盆��{�����BU�ɽ�z�;M�Y�y�޴gw�6���;�թ-	s��u�!$�˙�B+�����0�-j7���/�
����/���VM�I���0/.u�D�u6�.��T]�s�Hi���������8��P��~�����g)Nye�խ�A��J�нwretLV*�w��8��ì�:�ao��N|d�.�e/����7F��
�v�'�O�m,�,�R�X��[�-�ڞ�z!�jaW�vi�pds ���Gj�ѽ57ѐ�%ڄ��ӯ�e*�k2�
�Osz{����]� k�7�����(�{�䔎�l����3e��S��Ǜ~kv�u��˵��i6Ԩ��'.�{�6��94����ƅ{3S7�6�Û�u,������_%��z���I����:#�*ާ"�/9�*']��F��]�&X��c�<|�N�ϟ7��~�a^ɫMd�ާ�޹�ӳ�\3δ�8�6�����j�%K��\8Mm��F����]d�ar;S�O���gfU��d�2웃3[�-�jA\,����"�8�ډՏ�8����\8�pm]��`���&:��������BkR�D{�0YDMٜ�o����
e�]mG��=֧�N���K��[�"�5M;(��{W�#���3�m�����q39�)��k��WP'�ƾ�����w�ib��M�v:�fR!i�؇��2^��j�Լɴ1>���}*sF�Wk*Ȩ��1Z����o�wI����
�)et\dG*j3*^\PپX��O���uzҜ讐��iEV�p��n��V��k�[���K��ޚW^{R��\{�r�s1���q-�	್QM��8U��!֌�v��`L�6goe�Ê�.v% n�� QV�J���31XE���twM΅��.3N��E]�H��0��vwP.c�v-I��.��9Ї����ӀJܫ�$֮�lB�)'M�k��^*�]$s� ��jJ���f�l���}�cSv���8N}�KW]���6�s0eͱX�ky�w�D�s\j���&�;BQݡ� �>;=r�5,��Mz37JsO.58Q���0e)����N���e���e���j�k�l�]�;=҈��A5�`��o����^L��N�]e�d�G�!2��;>��73/���7�C���q]�)�:hb�8���Z�8#-��x�����Ɋm�h�=ʂW�K"�u.����2k̎#��on�6>33���P�|����J����t�K�q�����*Xp�!�+uh��tlv]$�`
�&'�!�h�,���R�F�1�w1`i8� �lYUW
c,Y�<tAL�˨[)"@R6
������n@�a<���B
��wD��>��na#A`��f�%�,42*���j�$���]���;M;�N[�U�q��v�����;r�*S�DJfV������M���Ncuv�{X��
a�'!êf��HXk]�p�J�,��uvKK��\��Ӓ�P��~�I��f�{��V�OE�Z�����`��X�tw/�]�r�|?���$/�r8!�ۦ �nT��ޙ���3k6.C�b�V:99)������)��^,L����9��3c4(�T'f��L��>��aV�,�z
W)^��IG��I85�3����7�t��+0�^lJnb˻c]�Ow�}*%��mAf.D
�k���nT��5c����0��O��̑inv���3���F��EҚԞ7�G
Q�B����C|w��O[�YV�f�46*�%='B��c7��7����.�ڀ�V���{ܹ���Ϻ�sx+d��*F媖_E�ٗ�w��>A����D��4ƪӾ��Wh/9; ��C;��:A�vnU�r!i�9�e�c�!�T	�@%���ނdg%����u_h�+�
��_��h��U*%,��ZT�mb�E""�iE�"�(�X(�-�Z��ȬEc��*�ģ��(*��h�D��"�
֊1X�F�QUr�Fb
VZ�-
��ł��h0�Eb*�QfR����Z�����mE�Z��F1�&]0�t�5J�1�QEQ��kj�(�UTb�",�k���km �FEF,�D�,P�lPDQU�D-(�m%DQETb�ƪ�9leJ(�AE�D*�Tb(��e�
Ŋ�1��
ł
�l-)eeUUUF1����V����DE�ih�ct���+b���]P��&	E"�� �c�����,A�,+UUm��B�*DjU���R0D����e���b���aR��(��Ơ�"��,QKB��.�\bQI��DZʢ���F* �0TF++EU�,��V2(�iAE�*�Z���c"����e�Q���Q�Q�*��T��
DV,�QE"*��Tb��$D�Q/�1��]�]��Fs�6�wB��)6�Na*��Ϭ�&��&�;����kEv.��k*��JԉE�/Mb�+P��	ū.T��ښ������k�g#\^��I����ƈ%f��=\��J�V���I�r�}����(���� ��E����"!��d��[�0��vJ����÷��b�w�:y;qݲ��d6R���3y��C���{Uy���U]�\�el<��Vu�J����֟-{���;c��0�}uY�����E��J�	����O7P�I���*�Fr\�kf���Fm�ǐ���hip��W:yMm7bz��S��a�U<���oG>J�KF�Q�~��ɺh�
	�9�3ꕱ�+*�Z�8�$�
��˪�kx�#��vr#,�y�����U~��	Lϡ	T���]q��,`m�UJ6�&�w��/`s#V�� �i�T�H��±ڐ�l���M!�i�ng:�퓌���t���2
Jvkύ��p(2��6Vr�M��T��h5�+k%����t�uJ��%'�@dw[���	����ʻ���;2�|4����9q޺�m���])�{j[����B뵇��IV����� pe=�>Z�fp�~�X��,��[��N�������N����,���D�ʰ����E����c0mdMy�B:�6����B/�`v�@�{�l,Ӌ���!9�yݜR�q[�D�"V��,e��A��!�{+}1���OoV��~�R7Ue�y��v��ޜ�9V(�,��z,9F�0o;hs�ފ;X��の�/Z*S�k�ͧz��ɠ���XUMX��)>���Yz���\���hWʂ�{�-A�ݛvLë}yr�	t�竛jc{鸠�5\:[;ؑ�ı�iϜ�;Gv��g�S���ٷͱ��3�C7���k�;&��B◷�.톗W�5����;�'8�kT��ڬ�*�Xv$gn��X�ѯ�y�~��nc�%~<!OoGt�
tOb��ڨV:�F?*�{.����sΠ�f��O�J]Cy���/�Bw���7Y6)��M�8����5)�����c#\��=Hl7Rx�>L�o��ֱ���f�q�wE��O J�-�d3(�o�tA�d������*˧��;�LWWGo9������7�Թk�(�O&��-���^8uiiˎ�,D­,�uwM�ȭ���Ys��Tl�R�2��,�%����z�M��J�^��I3X,��H�!F)�J5����]$]�P�m0�KDKq��jÄ<'[z\�i�{���.�w���l%ו�E	u��z��]X�ÕW�]f�	'k##�x�������]^2��S����Y8�enw�V�YPލ�n:�HV2�U�T��U4�����e��pgX09�:<3U�^T�-���Sг�.�!���sJ������?m�(g�*�zi�̛|�'l������B�͠V��z=zN�^�����N}y,VZg�v)�X�m-ۛkNP|�U��Їz)��wdZzØ}�i����́[�^�bE�c5#�Un���\����v�Y�+75<�8�t�qq,f���Zf=xѮ��5��}/��M��w�m��+�̞�y�&��紂|2`x|���I�'��I�d�;=�q���(d π��a���cp�*Of}�5uC	�kee���F������$���6��ҦP�*����݉�]�˧:���j7�������-�)ׂ������J�*��qޤ��P�N����u��E�}\��C����G(�=��X�,j���:U��Q��Y�;+68{���3nD�N1U~�|�j}�3�}�kA�8ϙ�a8�����I�_Ԭ�g����ì�I�,<�C䞲U�U�yˑ�`�y�bA����6�;�E�}�r��k>�Gޢ0��|�?3g��!��}�>x�u'�s ��Y1�O/����,Y��w(�~E	��ğ�x�@�����M��_|E��w�l�������{̉>�I����d�OY�?r�Y��w����i��u2bu�2�*Nr�Y'�h�~E	��ߍ���^zW������~�s߿w4���t��>@���!>Hk?d6�a8�j�����Y�!�<g��6°�7�jd�@�o�'�m�f�;�:��ӿ�s���of��o���U��� ��"`� ���T� ���dRq��M>߰�����z�q�$�g�쳌'�K�C���sL�3Hq-x�[g~�W�u����?wO�������LE���+s�Y'w�)?5��ֳ�0����Rq�����!�}Cl����Ha��"�>>���AE}�&��[�m����	���d��}��ORb,ٮa�V�r�8���"���I�3 |���h�'3�hN2��q�����ov�*�k�s7t�s쵶���P�&ӧ�u$��M�!�N����<E����xɖ����d�氺��d�_�,6����L��}�޿Tx#��}�F�'��r�����k�}��>a�C����Y<gR{!��E��$Rq3�2VI�����{hO9g�2e����Jɟw=q��޸R	�8���v;�;�_՟}!n'/3s{�x	 q��$�Y���
��!:v��'YԞ~�zɤ�E�ԑI�Ͻ�wvI�l�2I����y��x������+��p���Zo�ֽ� ~f]��<��T���g^
;�����\U�2��v��>����
�Mb*P:�r)�4��~�o���]̅(�%.ΝB��;s(bOc"*̡#f(���P��
����'$��3iɏS.vVLr�r�8����^��:N�/���<픙����d��>�=�8���&��O�2u�z�g��:Ρ7����E�g����N��� u>�Ú�M3������|�����T��Wd|6���G����xA�>�J��!�`��?2xͳ�T'�i�}�ԓ��5�qY&��	�N"��O�8��5a6��y��s?9fſ���\Wd03c��|>���g�H����`~C�4ý�z�T<�w�E'�1����>d�Cɫ!�dѼ慒~I��8�I���q���������|����]�urV��>�տI Y�� |�{Ì3ɖ~x�~C}�O�<Ȯ�wR���0��}ԟ�O���C��!�d��Cɫ�M$����?$������wop��WlG����������(drXx�O�d��3|�O^�:��fC�>g�C��I<f0�I�s�dY>g��Y:�l���<���S���</���μ���UY�>��>� �"�7����'ό�a��yC�$�����!ԇS���3�N�rZ!�=d�8�~�$��a����3_��9�w�9��������Q$�#���A>2���MM��I>d�s$��N3�>@�u����C�|���C��o���8����u��Lg\��g?o��{�<����{�$�����$�~���C�fN����dP8��'��Z��y�&ߒN'��I�����<>DX�#��vK+���8z��1_u;��~��w�u{�� t�ߵ'P���hN�Y2y�Y'ל�d尚;�:��OZ���8�����!8��}#�~ {�z��D>��/Ъ0��.����®^.?y�I��|;d>��z�����=f�<7̇Rm�f�s$8�P�h��u'�p��$ѽg?0��Ld�Ě}/r��k�o3��������mf�kq	|4aވܣ��X�-�1�\.�<M����,n�Q_v��m�+G5$R�gV�*f�z��w��}��[�X�[|�;��t.����4�6V����#��.=RQ
�_Î��u�βpૢ��W���{�>�ָKksh��(�y�0��@�>d���2J�f��C�&�w���=T���C�=d�Y�o�!�NX�q�������vy���
���\��K��v�P������}�#�}�� �d7��g�4��<`,����I�
�L���N;��u��X�!Ԟ�e�����b�9a:���>C�����΋����U�G��$��aSĝ5a�C�1�߸����6é6�x{H(c'S�XJ�S�sA�Y&��������G�� ���_M�~_c�	 	>n�1��&���M?��M�,�x�Y1�J�!���<gO6�:Τ����&�8���"�����uoq�2�D.�������`i��G�/� 6�n�v~� ,��>�x�	�G�,����O���X5�N2OP��N��&�i�2qP=d�N�ui�ڑT�;ࣺ�ۺ�_t}�� #��>��Hl���d��'���iN��+���)P����=g�0�zj�~a��^y����7�N"�w^����h��Qcy����^l��@G�a��2x��N�|�|�����n�zß�u'��O����<M!�{�~d*�;�
�3�`|��!�y��4��g�荸�����|<����	�di�'m���O�8��S��6����?'XO�9߰8����������$�n��$��;�M��C��W����o����9Ϝ�6���guH|�L���I�&���,'���'9l������g��08��<z�q�ݧq������C���=׽��]y޷}�z��g(A+������#�e	�@�<,u`q��=VL�>I�&����|��Y;l��,�d�9�$8���s�A����|�dy�atݎ���5v����8�C�>���]Ϋ��iڳ��mͼ�W�jV♴��MU[R�� 1ޢѷEP�U)[�A�|��@h��7�]�8���kk�q�1!q*S)�z��������X��HTxw�������
^��:���kQ��nщDN���� �Y\R��s�� _e�3�4����5	��}��:�8�O�B{�'|�����󮤟 o�O���=Iԛx����� ����B���~���u?x}����޳�N��u��1���$��0��pY�	�6wY�"���2q'̞�'��qԚ7�i$�y܆�������0����gk泖�� 	;`v{ġ�=gS���	��z���4��{�q��1�|>�	ԕ����$�=��R|�e�@���dݠq q�X3���9��J�N���nO��G��s�&>��g�����Y�Rx�S��2�����p4��@�;I�d�g{Bu
��h��q'ǝ�d����O5��C���ԭ�j;��'޳�tD���Hz�i���O���
�P�Cs�'P���x�N0��u>�Cl�$�{��OHg,:��LE9�`N$��>�C���C�����"��ǽ�#�����a;������z�q����!�!�Я�'זé4χ���*a��gXN���!��"���7�2~��x�?&�FQ߼ �3�L@�P*�r�8�gy����	�3 |���jjÌ�c5�p' ����$��LHu4r���*t�9���K�~�����u����O��?GO�"x�Cs��*��l5�p�P1Nk=q$�#���a8���<g����q��͟��gMyOP�'P���׿|"��k��wg����Y������f��"�x�w�:�����d�-��� �C���+	�G�(x�P�O�`|��&�y��	�9�n�;7��gr��ߡn��}�#�>�l�'��l=�x���G�H��=�{���&���d:�����z��'��y߲d�3�g���0;�(z��N��[Yyn�0.���G"�r4��H"NW�o����f��A�l�Q��畭R��W���{]�ߐ�9�Ӵ���*g�wT��\Faԭ�z_u	���䭌�h����u�L-1s���$Owrz�)����<��#u3aX��80�?�������{�������N�=�di��>���7���q�����O���d�Ϭ'�M~��M3�l:������a��:a�Y=d*?���/<�W?���|��ׇ�~�zT& w�N���g�xj�z�L�7�'XO�o�d�E$מ�u��P6{a���������ݳ�'�w�$���9��������wd�r֣cw~�|���|7���� i_Qd�<H{��|��=CL�VC�dѾb�?$���q�f��8��d��>>�Q�#��5&�6����:?��(����y����|>ʀ�@���xoG����,>a?3s�l�!��!�d�L�>I�&����~I�Y;�y�>��}Pnghv�_˺�����=I���s�	�Sgu���!�O9�|��~d<��u��C���Y'��3� |�Y��d�Oa锇�{O�L��D]�"�//�[�ç~�ُ��RO���=a�|��{���<z�{`,�S';��|��O9��zɌ�xw>�'�1�Ŝa:�����(=]3�G��	�-�f��#�
R�K���׺�|��N�I>@џd6��u<Փ�M�`n{C�3�|�'�d��h�~g̞�H퓨i����N>@z�ē�y�%-��d}�ǯGM������kZϼ�m'M�|��Om'�h zɭ��Bu!����u��c�m����2C�~O��XVg9���H7ܓ�m�e���yT�~�����z��VW��G��PO֒s/?2}l�N�<I�����8���a�����Ru�fY�q������{ѝe}d�����fO�{��z��i���6�f}Bq
����$�s"��XMM�8��OY<�'�۲�q���+=d8�Ć��M#�5���}��k�y����{��p��yd�Ʃ�5 ���Y6U�-e'^�F�۶C3���I}.���k�������������3�-X��|r/o��l���΃f�vw
��xҀq���|:�����y��[r]t�K��6��:!w]Su!2�*v�tu�$g�=�{��o�
*�ޏ�{�|T�ṡ���~O/y��'��8��6�g�su����I���m�$��2�+�&$�C�c<��q�����=��tGV�W�w��:����=I��c'S_�ē�
�ϲVI��^`u��X;�
��&Z��!�La�9��	�M߲,6����&|0�O���}Z��*��䟅@����<a�Ca�<a��l�'��L`qGԑI����uY'w�d�Н�rb���?NX0+	��${�z�?�Զ����O݉9���a���t��x�Y7���0ѿ��C�M�g�i���O?~�?2m'Q|I6����Ւi��`~k!�YP�"����ik<�-ݬ���7��+�y������
����a6�5�:�=a��d�gP����4��Y=@�N��/�M�u8}�!����>��+����D�;b�|)�?|z���'g�������Hy9��2bO]���<`d�0P���<fوOS���:�z�̲qY&o�'Y8�'�y>��n�U?np����s>i�}��d��~��XO�7���z���������i���I���{��j)<a��0��l��x�2zo�,��Mo�<�${�yf�s�syw����jg���`~I��NZw��0:ϲ��ROP�w�0�?2w�5!���'<�=a?&��O���,>CL���<����G�`��O>כ�>���`�{�I�����d�>2|����ORu�i���2C�3s�oS��'R{l>C�z�nw�ē�79�u�~M���'��!�3�:>���w걗�v��j�o�Dzϼ�a�)$�&�����̓�d�>�u��$<C�$���C���|�!:��O�|�Y4�<�f|�`���8̍U�WQ����jȭ�q�ɻ�t�N��2�έ�[B��q��%9I�����?e�����Q7���Ȭ�aR[�xvDx���viѻ�)�P�p�Y�>�ÿ�JT�{��:�}+N���%�Ř�#�F�Sm\,�j���_��x+�׭�P�{�	������F@��M~̟$���Xy2��Y5��RO�73�'��q���N��`q��s�a��y���xì�h�2�b_>߹����Y�gޓ�?DN!Xg��E�q�'Qd4}�8��Om��@�OX��Z��s;���I��Փ�O��N2C�|��}����u��ܭΎ����Z��<	����ʇx��<��'�m���su���h��8��s�����u�5'�3 ��4�0�`k�&��:��ױ�6�-���������>�NO��3��r���I�9�Hz� y�d:�l��6�u!�J���E��L7�O֒o/>a�������6럼���y�����;�����ȏ��}�q��O����<O5z�?!Y~��:�zs��6��<��C�=d�Y��a��4g2:�N0�(�~����ߓ�o;�k����.��߻l*~I�VN�<C����!��3�M����i4~�d���џ��uI�u�h�=;̇RzɖÚ�:��o����3N_���y�n${�w?��}� ����?0��OMXu���o�	�C^Si���=�1������T����,���Y7l�{�۝�-}�����5�`A i��d� 	>�׺1��&��)4�Bu+�g���É%fk�&��p�xx�l�gRz2z�08��H��_y��p�������εm\�0O׼����߁�w�����<�����uf�h�|S�>����Ȝ\�z���馳2_[���m8̪v�7A��"�%�9wT,�=�3,ғ�
+-��MCuP��D.���L��m\U�d�Xt�)6i0:sޔ0��I���p�>�%��ت���ʍ��Sj�|��4fU��kr��й��Er�a�s�M��|�yy��W]_,ӊ"ay��E]��	��K��z�핂�U.�e��5}������Q�U,�6�_P�.�B&�L��wV�	)X����U����� ���*�r�c�	�m�c3AJޭ*'fL�Q1e�����C�-�hpKc���i��0�/�{z��<����g��%��#4N���u�Fg4j��A���C����Q�v��M�:m���?c��QӵÚO�#�O5/f��:M�fc��n!۷>Ƞ�Kq�ՊH�[W��;L�hޮb��c��c��f`�|��lv�W��V݊���aL���K���]J������N�ݻ�2��|q̫�PƓ�'��f����+i��ofV�i��\�L��w���닾��ք�{H���ʇGQ��3*NT�*'R���WZd�.=���Y��c�Sx.�{�KMGq������M�^QEO�h��d������%0�Ck)[�A䈫�G�"�BAٻ�^�[{.� ���m&��uNO)v���ܽe�[�U+��c$:��ZXX�v���ь�P�sV��[�ݏ����b�^=k�n�m.��M*|v��uQ�`.1���N��TZ¼����^)��
�B�X�|^�R��<����N�ޕz��3�en���47@��hݰ��n�&�ۺmK0
�u*"(F3%dB��U�n3�*YbEDV�Pf6Qʸ�wy����˦�h�>ܕwf[o'�nV�
���MPQAv���nY��T`��a�fc� ���R2H��"�\!e���d�I�N�h}(�1�SC2^$��M]�)� �ڃpϛ�'�ۼ^�Kx[G]h*������$t�ԥQ���St���n���Y���6f�i�qq���Z]$GSr�NA�.��r��*�Gj<�ݫ��œ[BD놷w�',��*��j�`}
��}i�jV��>9�"�U�C�/&*�T[xR��2:�)�tCz!u��X�;:��rt&,Q�jD֪�	�U�*%j�ծ�l)΃I�{�f�q��r5C�s!wn8�˽&�m4���g.���]b�]�(KY�%�Zh�nMǝ�;��v���*;UdK>j6_Bd�7�S��7u<����@T��J��-P���(�Z��,�����ɂK��K4$�
���*�eP�6F	&.`����<Ў-R���٣���_^��J�V ���#�Q�D��u�ct¥.kwmL��:Nx���^�y)M �h���$Ɍv�r:ج��qqm��i�6N�[�.NG�r�N�����ݳkӳ���PRPC&dI	���(��>��Q�c������QTATE
�[t�AA1*��+�(�PV(�X���X��&%Eb#�KQeJ�U�klTiDQEAb#t�W)Ub*����b[V
1EUV��b�����U\d���J��a���"��1�F
��Db�����QDDV+4¨�q��eA��ŌdQU�"
1T�1�1��eB�b���������EYZ �TV,]0Z��[(��Ȏ2̴uJ���)�-J0kTDQb�Q��Q��E�ՠ��Z��E1b���b���EQ�TF
�b��*�őT���Z�V(	R��%�J��(�eAf[�+�QE��А�I�p�G�U�pu}u�{�/"#{ύu�)c����{~�������'6\����0+x�nduJ�=rVq"8�*�g�������k}�y�Е�K������o�으Wy�s���<�rx k�Tz���}�^�F_;����jF�[�|��+�z�f��2U��!���ֆ�h�x�'�OCɹr�k�υ6:����+�c�����&��l�f���ɻ��i䡻�"c��#�R�3֑�/�ݦ�t��U�E�8˾���ճY�d%�z��tPR8q]`��=^��P�j��ޛ�4��xaE�ٞ.}#��/N��R�=�hp�Wa�V�Gd�+�#@��r���J�4���wf;����oP�K͆�B����CC/��8ʛ��Փ�{�05���_����={P���Ǎ�̦��~s1�:�;��������ʣ�Ei�Yl��\�T�5X!����]ۍ^Q��v�v������u`�u�(K��L⡁��� F���땘b~p�a�\9;zn�,��lñ��M_ؓ_7cr�ٵpm��g\]C��s7�'�J�2붻*�6�T�w�.��]���U�)�b\�aܻ�`"�T�v$֥ܣ��K��V#�kι\�`M�����������X�f�JS�[�� zRV�N�&y�;+:q
ݸ?u!�!O���I��X�8V�pg��&�-�u�Y(R>+�>5q*r��y^��km<�T=}����k͊��4C�b$$�ך7@���)>�!]|r�;9S(y>]��n�\�P��&+���w)�֖d��`. �lpW���Ou����,�~-�l�C-3��v����|���b�v���rpyf윬��ۛ���]��	����FU'Ϟ�Pʱ0�1�F�"d���q�����wu�J҇��5�3���hubfFkF<�5�N�oyodK�(�܌�c�\��K�x�
�z�X�ɤ6i3�wj.:Nqv�]j�dt�K;��g8$e���r��e9��e�kL���U����Wf�e�gη^ĩ�0�����+��-�ìC���"�r��ن�#�.N�q%eC�������:Gd�Y#�L�ܚ�P�I�'m3��c8;;}[MB�>��քm��38��9m-�Sߌ4.��鶡�I�?,)�s]�%�]#�GR��ӵ��<�2�r1;�o����ꪯ���OV�w2�ir��vMF�AW(�x(�^�yÞ��z}��7��Q�&Ӓn�o4U^�Dlv��tm5c!{C�Y������z�{X:M��m�� �|z+�ke+ϻ:+�9S��@KM��.65V�e��z��1{�Y69�H�bP�4��.�%mP-O�q�5�v���u��ի���un^���칰Ӹ�LȄ%4+_㐺<�a��%m�wqkw"X�r��	�I��v)7&�0!	t��L��r�+��]׍��l�6�Em��t�8<�8r��F��J�.�rڴn���yl�RR��	[~����R�^��nK�[�����J자a��[��<�Ȯ,ꢘ���T"��W����P��خ�G�l��ń\(�жxrۋ�{�6�[�-[��Hf�_�&}M�\� ^4=���9C�����u�Gʆ9N��L�w�X�e�P3X�PUF	��{�q��CR�n���㝕�TU53}$�5t�W�	H0�p��j�k[;c{k���cn��w4w�OOvs�c��g��oGr�c��y$k���mP혹_NTfP2'BK��u���꯫�����6_:�?uZ֝nm_ygn͆��>g&�Ֆ'&}Hm��vz��b]�I���,�x��M���m^�z�eU���YA�VV��aQ��L@�6\�����v0����FE봫�8��9K���Aa��kv�H�i��`{k��&���3��)v��մ�)����YYc�cr6n�r�ȱX7�t�_X�Y S����g[į�ڃ�{C��`Q&V�W���>Q{�^��V+��/(�cD�%��y�"r�;[���T�,�6g��k���<���ڇaC3�~Shi�/��eSrkĿDyK=�n�sxw�.V{��Jne9���#._�!�&V��Eފ*�_>U��c��MY+r�X�n�鑓ͷ4	O W���Jh�A�k}0`�M7;���S��>�ީᏯ�ν3�	�i�cj��{��"eD4�ǽ�rv��������xA�6N�[כ�n�����Iqt9�]M�N 
{b��TSc��ˮ�{Eu���ZL)]ɢ�A��&�����k8�=��4.7E�f�� �Os��71n�ۮ��=�mۇ��<��+c���mǲ�| ���M&�k�+b>Br�pVu�ӑ�,V)��j�L�50�b'n6�s�ͻ�k7���4�q}wy� �!׏	�q��%]*r��rPu�%Wۚ��R��)���O�v��`�x
��+�k.a!*���hy��l�P۾A�[��R��Г���v�M��m���D���l�
&U6�Y�[{�QO��G�{P�*>�y�3�6�y���ѩ����5����|L�	s"�{���xV&s�*��խ�^�׻'��B�F=M��=X�NH�U�s�"��lv�H�Z�T���;{�����L�'z�����t�\W�j��oT���	���o+3�F�N۬�Ɯb��c2�c���l'A�)4��@GlӞ*_k��ӣ��"�=�G�o�7�^�r|��!�;�9Ýy��=��X+4�3'5�n^�[��0�s��M7;5�>�I�U��v�Q��&�pPF�����wTY{�����IK�ipj���)�,�!κ8�x���j��a�v��m��pC�8=�ج��H�L�a+�1h��1J��jIUX�����f�˔ļ[��T�D�%տ{���<�������>�3��C1l �kiݾj�\������������_V�,u��M�SU�l����wLws���}���9lT^�li�ܲ�{*�J���y�s��-77�����QKt9�]�
��h1i.���W4t
g��z��wd�b����x����E7�A�*q0���q�&WD�)��+^�6D�G�볩[�[�i�d�{�M'bCF��7��c���;�{���J�b/�5S��eԡ����F��BF���	<47F�`s�txf�9����ͷ�s�fU�:˔(e�+�c�\����i�:�d�gS�.]3�[��W�[)�"=�T�3���ݪ��<ڶDr7y�"�_w��\o=I�RU�>L�AV��h�VW���w���9�z�9��%�@3~��#a{���ӻ�/�������:���,*��s˶��B+]0�S�%���3D�Y�Wc��(�k�L�Pv�sX�λ��+v��O��z2ƚdٻ���}:wT� ���.n�vY\sx�7L�P}_}UUQ�\�̮~���r�˼Y��I���:ٞ�Փbri�hv&ENh�!v��,ٽ(N��K[K��^�۱�^�++�z������jV�ۏt�~�3�Ө(�y�#"Ӷ�n/���m�C���GK�gEh=��d�<U���nv�w-��z�q��V.���O���ױ�Ca<��V�b;���O`��5`�Gd��z�*�s��α�9��[sz��l�YT����=���Y�#qWa�VϪgnc���(��sR�)�Ͻ��z�-�q]6����t���._a�Zڜ�׫����]��Y��;���^]o:ɱI�
��ĺ���jWFB��ZE􇘷r���D'��d��,,1۰���	��%SB�<o���3'T�<|1Nf�����[��zO0�t84n�q"�25J��0/Ps6�N5�Wg�>��ݭ[�A]�7s��ɸq��Q�Ӊ�ŪgxsXL��Y���9���n�3=���f��%��'��7w�iĸf,0n��c�$��\�Y� 5����@�טX;���y	�D4��о�2^��s��]C���gP[c�`�ݨ�/kb�2��Vz��@���Lu�����d��E�š�z��ћJE㧠���9L))�|j@WYۡ
.r��mnjp�r�;gF�Ǟ���*�
t�u�v73�+�T^܆Őhɋ��3J�}]yŋ�w4;��w!�������rށ���b�i�%K:��b]���7�m��6�7 cQf���Syp��l�k���k�v�*ݙ�w&T��su�z�W6�y��J#>��@��b��9��9�w����M�~��(�o�����)7��VdҾ�lV5� >ד]��{o������s�>�5��H��~WȬm�M������R�z�_fc���[}��܍͎�#�E1Ը��J1+m5�;��a3�`��y�v[�݄_�|�h���_�,g�\Vm=Ƴ�����2k\�7q�0z�
M]P5����=�}db���#�vet,�Y^��R/���O	��}$�FnlJ�f��5��#O|i�Z��xV״ rHT}��Ӄ:)9צ}Omv;���Jf%�rnJ��/V�cv�#���E%�9K���j�n�ĭC>����O�;�7��o�~ێ�X��M
}Q֡���\=�e-���:a�q�*���7ܽٮa�:�����ī&�:�	�9��)N�*{co-e>}ļ�;��㎆<۹zdG7C���a<�2�\��>�kB�K3Y�{�[���X%lMgH�q��c�zpG0�t.VkZ����+^��kX��GP�՞ە�_�NL��b��J�C��=��ZMx�(-1!��.�Ck=V�o\�Y}�_vt�<���.U��[}d�M��p*���v�
��-<4ѻ��s�����?
�<���[ >��$�>s��dL:yumT=��syy߸��ӀT4\ �ͷq�2, �C{���m����x�H�B�{�~G�{�}�k��������4���.v�T�*�uC��fV���$^&sR<��k������u$D����F*�n���a�p����2��STXv��~��r]���߲�82c���.���r����R�+4���/ss(��%���ك��*�,���/����T�ܩ�"��4�o �&<���s�w��꯫�+��������?����&$k&eoS��T4��x�X�J�HB�B3�&(�<]ܣ�ee���y�ݛV(
�9��b;&������V�z����;|�uӽYZ��M�'�qݳz���}JG	�]����Wx�,F;�k��a˾��Z�9����Լ��L�Μ�'áv;�9����Qo�w$�M<W��=^��v'���u�6��Tc��7�q�gL��:%B�g��O^6�rV�X���	�����Ϧ�+�[Y��lױ��5������jsE�܎��U����6(�~��
Tt��u�{��:n˖h_Ll3�^�m*��J�pJvEs����1f�F���"�]H�"Huj�^�q��+�x\�N>=x�'�@���{�XWej�8x���3��q�9B���|��>)�t���j��{�j�EL"�H̔=�ڝ�L@cT���bB�S��fp�PT#���tv���YϾ�XBZ^���r�̝7�����(�l��XW:��ﮌA^��1|2��q�p�Ejvd]h�+۳8�/�(�(j���-��s΢9qM��8#DU�&��6�m��GO�{9v[f�❇��k�n,����x0�MN��}��bG�0Q\��ذQ�N�6��*
�#��������'������v>hR��+��t��IA֛r��Q¦;b\u4��,�����I]�1x�)�)u��	Pa�FS�ݗ*�wY����ュ��Ş�k���]�o,�9Z{|�A����H[���wB��]������8�:&��[)�&e���(��]�Z���84����-ˇe���Z� \��v�*٨�`
�*��H��E��;��Q��f�\�k��'e��`�o;��Z��@I�����]���Yq�*�e�;-RD����2�]�������ޝ�n �lc��$��[w�V�a��C!����ѡY&s�[Ά4��L�JAuY�.�J\�>�6�1�dt������3�WSt�u��j�Dv��T�ض�	rILWu�jΥ��ñ��5��)�z�(�gl�h9�ܷXY�W\�_N�GT2�[Bnp��r� �WL�T��ӡnH�vW�USLL�E�x]����c����vgf�5s�t�5M�[����E�;�<Y�P˺��v_w8��ȷ{t�E�[�os>�J�>͢U*7u��p)��`ns_��v%q��e�vح��i��&F�)�'1���5�P�C*--Gr��[ʧN
}�F'9U�%�v��J�-�2������u �xfxM:a�W�b��1%Y}�:��o�N�b����K*×����n����yCc�lAlp�<�BۺIaP̸���[�r�$^���8cj�����\Gj>.=δ`��
�F�Dʋj�(�'��z��w/+T���f�R�a��1U���0]2$��s�bJ�j��)Q�*�M�@8)�1�"���S#��,3Aݷ&Y���u�񹺻�2�$�n`jp$�j 4^Z������˷��d�o��OX7���]>���E;6$9ܬF���mEY�(���[�VoV��k�÷f2ej�z��Ple���޵ʐ�S����N���T��J�IX�o4s��"zhf[�/u�&��<�Q��3��Y7�Re��t\�7r��Mi�Mmr �[8egV��̜�A�,)z�v�]�mV���e-�A*P�U�|Or�W��y��3w}�%��CJ�ivȶ�����_l�
�.�pu��ӥ���(�	kct�pu]�K����yq_es�V[W`_�0
Dp%,ʍ.Vw1�Xvģ:�^��%�� �$�7X�������WG�Y��T�T�ъ�(�*��+[-�amV#kJ��&+
�5�*���W-���(�(���k��QE20E��-
-J��b*��EE"��mPc"�"�j���G(]P�QQ*��j�*(��4�Q��X"��+X���[~k6�X�r�J���X��[DX��ŨTUE6�wKDc��E#-
��نDr�ֈ*��V"��m�V)YU�i�*DPT�����Z"�[Db�UU"���������DE�YV �DQ�Er�
�e
"�̙���GmA�J�bH���������ݩ+F"0YZ�"��Pc7je�*���",V*��"��U��X�DWU�I��0A�Z�Q`��""����*	��|���;u"z�^����yj��s����c����doGm<#qS5W{�t*�R�s�oWax�O������Vs�Ra���ُÖV��ʷc&4��S&�+|c<�2&#��W�{��1�1e=[� �Õ�},���a�S����T�c���u��u����ڜ�mvE��ՌX�ǜ���+˲zZ��x�%#��VO:��-��4P7�ݤ\d�rӸ��&�|mOj|�;�1�ho��X[�n��=w�Q�p�꺤�p���EF�~�D7։��&����>�ߞT�/�a���[UN�a��A��f������q���Ξ���M2r��ڞڈ��(}��Y��\l{��d��9R[�8:��bsn��>�hЦ���opI���;"h�����g�9�(���c8�R���EA���Wlf�Rꦲl�����8�wj�@KW�۾���tn)r���z�җ�-�N^�e���gR�].�N,ı�r�V�]
�_�;�A�s���;�T�T<�h��dn�w�^������<ج��wIԵ���1��F(j�N}����a�!l_L��zm�9Js��ϯO�����&��^¦�Y˴$+�5�8����b���U��F�J�c�� ڻ���\Gq���i�7��3�9M��;�\|���	j���C9����k' Ӕ������#2��7�8��m�1��A��ힻ��Bm�㻰8�o>���A\.�9��Ĥ(�j���x��ɘ/z*]B>��N͊��V�(�s៪����SC����t՛�����g*2�8�"�r�KڀQ��I"\3�`�n�����i��)���'F!M8��n���p*^^x|;�԰��|�!��6��>��{�ˋ�܌��3:z��8�����d;.��jD�N���,�@�Ø�&�fn�V�V���r��g�0��+S�:��Oѹ�PLPu��X4�7&)9s��t�R�TPW;u6���m�t\h�P�8�D��umZ�6Y��$��K�t�

$V�yw�{(�䆱���L1�$���с�A���%�R��u8�x��S�@ux&�^�5�jP5w��מx"��Ǉ%WpUw�^� �ՏG�w7ɐ��ڤ`=bd�ۅ��V=�����|jU��'��4�X��{���f���d\ƙ�,�/X2M�r,a��ouB����!��CA���v�-��k�oB�;NB>�|*�*_l��=&V�����������jP��p7��/#JFB/�s�ŕY<��8m8��M߫���v��VH���{R�¡����]`�;�s|z��Fd
�=*
�"j�ķ� h�c��=~ӝ���]=C�r����.g�~Ϳj\����E�"E���w�z��M&%v�_{����ޝ�ܞ��V�LeE�}Nh��xչq
��."���0��OR���X�Ɲ���8��ރ#�4<LS�4��:���dP�'��Q�q���9E���&7/6m���ii���n���
 0Q�Q��H�|��f�Z��F�N8\�]�|�!�z.���\{h�0�Z�t��<aF� �A��g�WIF�GLb�QN�2KZmK��Fq5��c������d�mй�q�=���}�ʺ|��Vt��⹯��0�:�l{.��	~� ��D�~���q�Gk��&�:�J��oЎvFO:�*���]凯��d.���n�:$�Ьt�^���债[��<|�ѺRȀc3A�Q��g��&�`���l��1�	tUw���<%�g�~V���:�C���o�_-~�׼c��f;-���<�G����O�
���MU��%�|��c𬸩�d#�Ѕ�ӌܵ�?gjvAe=�ɟ{���^�[C���q;�\�~5=�B���|�*����*��Nn�ڭ�<q�E+ ��31݀����/SG�!�;�+PX�1�n���k)J|�V��9��ao\��]�H˼珠S�;Yȯ��y�����v���56w
ytpJo����;�t��c쨑�^��d-9�� ��.'[�پ���!�":>��8h�")�8r���'���!�.#�1�㼶;�Q����^�>��K�w�3}Aٺ�:����)ϻ=4�:͋fU{B"�gD�y��==>D7�-_�����U�ٲ��,�]]{{����Y�~{,�V��K�A�w�*T�-�e��XEc�y�(�Wj�ˍ��b/�yb����H����fz'+6t�������aW�/�ěP#pS��\Ni�v��$�Ц���r����='�Uqlm�GG9݊v%��T\i�6#�4��4
f3�f���ͼ���{�qc��
�,ҮVˈ�<5+Fl;��t%��84L��+0�1& -���L���aP��V +s�(��P���yC6�Y�llŎ,�h)��g
j�;���s��%og&4��%p�5/�9g�IW2V�����p:�3`tˈ�9�b���Q�a������`�/Ep5�H�Ftݕ,ׯ��W3�l	R�;,�q���畳e��-���^�D�06�����uTq!�5��\�T�p2�=�^��ӶI��~�%�FY)�˚�Kܚ	�4t��
x�x�ǁ��]�ae'Ź;+h��
W�iK�_��-W�� <�>��n�+S�oC��@�z�k�{&0p���L_/���������{T9Q�Uf�)�N�9�}�I�<�H��6Fl3~��r�K|�DƛS"�VY[�_�&��11t'�|�*����
��0���)�%P������+-V=n��v��^��EZ�p�k�1t|�Ѓ�l#��#�#�|j�i6�J=1���<�O5W����r*�G*�`90'��;�PC���N�!�/����b�8�u�!nz����9�;�l���L�ܚp�	�#�51"ly*zbژȘ�b �L�C,�'�Ym��u2�S�3�:�$�%����P6�sn6�J���Yr�)K���M�����:���L۝&�c���E�,�Ƒ#mPˉ-�lI@�%j�.G�ߨ�,=JgT�"&7�Nuc�ǖ]׹�9=��6[6�2��,��@�0n�JUv�W5Վ�V���}��V@�h=����Eo�v�rF�55�K§MP�(q�n.w^�����7˻f8��'8�5W|Q��Z{�]��ͻ����	��t�΋\s������5DV߮R��/�;�5P6(�ţ8L;���3��}\ڜᢨns�ݙX�����brD��ނ���qS.!i�����gow�Г;u5�Zy���_W��+�WƐ(�(���d=�NT��}�q�3�jH�e��Ӗ.��{��N�rc��Owmr�״M����'w8��nA�ŧW�������}ϝUn�8~�%��Q#�1>�E� �ˡ��k;��(�#�׶��|�5YV�Ұ����TLɚpX�g�UHؗ*!X�Q�R�k�]|�;q;�*9�a	�1ݹ��S�'ټ�#�Ԣ��D�8L��%N����a�(}�G�
��p:�������c�&�Dz��U_|���ޡKW��6Oau5������>�����k'd���^�'�=U̠6�:g*2۫2,�ɀQ�H^p�a�=h���׋ ��=���3T�2g'�������'](ˁ�����Vd]O��1��]�p*�u��Fy�IG{�W=�M*pK��x�x�Z�lE	�d;�X-Cȑ3���Cj�*��L�=Irv)̣H�=1G
3l��,�&\P�<b��cۑ`�jlo$�&9������}�ك�O]��N���\TQ�>2�3Z^}!��D<[���;��'evn��C��@��	U�����-^d�����EO�躆�<p�c:�T�*�\d!�c.���p@��:��X��L� _=M=�e�v���,מO�J��a�SՂL �Cʲ�
`�:�R�=�� o6+�Ղ���ϻ���0'N]r\R�l=���?}U��_5KƐ��H���~��%o�&}�T	�y�9eɓA��������#4ePd*�o�����N�X"�b�*��-z�U��ٿp4:^��O!�;�Q��;�}ï�\->�Z�-\�Y^��5�P�»��n�M��V�&���/H�뗢�b�������v;��jGt��߃m-�/P^/ ���FT"���謄��62��ZV�_G��9��a{�B# �t}Y,��2�(�R��J�e��<�x�Z�"]Z�_��X9��(Q�^�����q��D#X�^�F�'�7%�&f�SyN����,�j�ΰ%�,ߜ�_T-
%,{B�< t)x�ri�5Y� �}3������C����xG�t�׃��鷽x�|��h�1�H,�@�,B�$�B;;�,�a
�wmrs�n����e�T��s_��"V8�suD��(�`��(��'�6,�^�
R���w�;�K|�a�š��|=)���.�W�N���2�r�%�{��Bj3h�w���sHz4l�Z�h��5I���+9/��kr#ۢ�ӹ$��r�����6����D�l��:����u-�*��l�9�����r���F�6��zf[7�3Y	$2�R�W�$��6eY�z���7�/�����<=�+u{�S+�;��K�G�B�o�	�
��c�'$��o}^U��\2d�Yq�E�zhdmPD�q�$JAXhR�f�_3�?+	�|�_t|���p'�M�ʾJ�����~=?�iR��u'^�Bb����t_:��*a���3#u�LHӞ��6g�e����=��'zl+��'i������yO�%n��x:��^������罯v�z�>ʠΛ�C����@�A�8r�]�;��BZY����ڄ5%���gix�[́Z�j0��������=U<���wY焱�l[2��p �3�2GIY��Rק����۪æ�i�eK��,�cg$���T�Ų�dVJʙu��I���]!���h��2.��ED`�E?y��P7����ˆ���\14�Ú�EY���[���;�wjl<�v�0k P��bM�uE P#f�0xީQ�,�z%u�7Y.��*��Z.�V���U�y��2�:Λ���"}HH���1b���_T֖��X&���T�Y�n�:��,P�tz�8�'P����+wh/�����L�F���&.�j�FY�a:�逤w��:
�S4�v.[���*��}]��$cb�|�Z����1�*�n��Y��_}��R�9:P�^�	b�䷀O��h	�!����dO.o�����4:]3�c	CUȳ}Ό�ʺ���4*qf��+B��t�^���|:j� 7Ћe�l�����Ό>��I&��_�z���GMUHߦ(�WS��2�:�Ҳik����*���q��#j��a�v����=��QM�$#���up\x��O��SQ��R���j�<��1�0�߹.%�����r�]zƀ��Q���]{��M�ﯦ6��3b����ƶ�O�.�3�񈟫7F�/ԭ�3����;��O��A1T�t�G��Dn�P:8�f�9P^���'���m7��	T;��/��Ms��P`�KI�&�r/��Y^=Ȯk�h䞋8�R���������e:�m���b��`�U�L�k�/ZR\k�,�v��s�h><k�ۦ�52߄�O�׺�~�S&����j"�bo3�{ �ib�Sɴ�p�r�DC��Q�sa����P6�sn/rh��e��ڢ&b3��/����|���0� hWk~]|^��fl��g��6���V�cSLܱ�R6�;y�b�|�4wA4����{&ֲ�h<3mJxO'�����-V�!���B]�|gq���-���J<���d9&��U�Lܛ��Z.�&��W�W��;��[nX��c�j��"��
���
C'*�I{��x��-p��#�G&���~�xB�A����ghQ�V��=hj�v�=�_�e�uL�.
�Q��W�v�ր���-���D������}�Xv�s�6*���Eh�\cm�������w��篼�h�AӬI��lW.T�!\s1$c��h�`%i�:Q�/���\؇����T;ko��G<�z;�2���2���vԒ:�R1C!�p��s���*�C,�En��#g*'K���+eOR����͵N�:����6%ʈ[2(��C�tK�C�E���j�hv�v����;��zC�d"�,�L����@Z�F��6��#Dh�+#��G4A�1��֮7���1��U�x�{Q���:|��P��v�m�����߲a��ӽ�T��j4�iN����5�}o���8J���ٺ��C��,H(ȴ$�.X`�n�3ݛ9�S0:y�ab���ŧ{l�tܹJ�p0rW{Q���̋�:f*3д'b'�aeo>�.��i ���;}�$D��CNs��;i܉#z4'Љ��7f�Į}}@�n'[�M��]7I��Ւ��r��K�z�P��J�"l�(<U�+^�__^�r�i��T�)q�|�BU���O�`�a�[��z�y��qn�GxH�fIl]����q��6��10X�:X.�r������a>��
���1b��
U�7��O�(�ѺĒ�ݗ��yӄ�jM�<��*ֽ���SSV��gV�=P'{��ig�*P�'�N�"���'C���
S� ���x���D��h�pl:)����܃`�2WCMɋ������	.6���h�&\�V-w��T��W.��+��H�\��N��Z�-=`�X�j�D�7�a__Svr<�k�P��\�r�_]D�uW �p�T�S�ؽYB��*���aP�Y�ݙ�ԥʊ��wOF�:ۓ�WK�� 7:4��=���T�����.�aa`����V�����]^!�T�t(sr����=+��[I[ɩ�\~.��eb����a	���[�W^R�_�&���e�u��n��O�J��:٤#�>��-镋#-|�^L����.�fðQz�,|��*iv��@��忡�s��Jr�9�q��"���ʱ�7k�*������r�vMjX�l�|(-�\f�k2vM:�6��St�7;mL<fJ�ٺ�V�X�st������h@);��LJ���a�[B��+v��ڂ�e�O���zg3V���q��=��n=��&�;��&4�ǃ{u���0����,�X:�_SȦ�q�=�z�ֻ��귆�7�+�[3B�-E�`+;�Q�۫H�[m�q�jy`K��iӟ[9[�WQ8g=���4��]AwN�	۬�@E4ڬ�8Lo)dhʌ�V%���(![8�P+#���t7���9ܐ���[�둶���J�����C��o]������7���%��|�ew�6��'{�6�g7�M.\�j�p-�1�,����=��J�˙�(*}԰�٫��^�Xǵx�;0v�Q��۝��Q!��<v�g,��.���'�oi��q�Ō}}�+��R��#\��i��T��O9��R��A�8*�*�������o��m_h��s�`��
��9�c'&���\�ɴ:͜�H�ո����RZ݌X�q&efG8&��+=��Yܧ�n�;�]��E3�ޫ��^:��k��S.�P&�:w#y�n�=3��b����t���e-˨v� )�;�&Iǲ�*��[�IǓT
�>�o�R�%[��uO��[\�a�J�Q]��N���̱8N%�v���eʗ��P������B\����8^e����/�M�;'\Xy�9v�n�p"{5�n�NR��kM��I�o|;�v�{
#8�|So,�S��%����Ȏ�.���􋁡�E�tE�:�]ʎ��5�	(K�� ���* *�Fe��~�5J"��%�b�TV
*,B�(�`���V%��V�X��0m*ͥb(��f%TV:�E�UTQm(1X��V
�*�b*�e��*�*�ы��U��*)����DEf�X�Q���b���J�"��,m�ff�UQ��D��aX���U�EAb��*(��*�UH�F)uqX�U`ɻEUAX�F"��*���i)�,\�X�(��h�F1QV�`����V+��"6�ET�Qv�Fڪ�P���,
�,1Ld��m�DAfY����$Q�*�DR*1�TݱTQ����kX(�U����ib��,U��R
�*ĭUEb-V��w��~��oy�S��X���i�G�25��z���%�fs՗�*K�'�na���(�À�Q�olB��R7�t��k��<<�8�r�]�e_�+ִ �TX�ƞ'.F�h���6���H�J��6�����rM�ι9]��N���%����(�F@�v��$ˊ��LPz�`��u^nk0�ژ�K�J�6� ��X���߄��)���r�/����p�O�(uiڱ�[ق���spԡ<��IQRc�9�Xw��K9鈞��H��
�:=�C<i�db�os�,�%{P��į%׸*�c�c9eɓM�/&o#q������U}���ڵ��ݸ�$?b��p�p���'�(��ތ�sǎQ�.(c3R]��ޏkλ��O�G�Y!��f����?N�9<$^@@�a]�p���g6�v���N�V7��BY�N7T8;�/z�M�xз,�d��ґ��,�^zy�ۆz�]o`ʙa�̜XU�i���{[�{���]g�
�5��7OS��z,(q
�Yq�E�a]q]g�,r�#v��L.qѪ���[�Cqs�H��*-yG�P��ez�ブ���b���]mNr��h�,���^�)�h��>B{�k� �&X�Vv`�/3T�>�z�j�3H�"���K-��A�	h����_f+Hmd0��Xy�3F|��:���=�ܤ��ݢ�rו��9�G;�?W��ԇc�ثC-3�u}�Y���J.���E��%[P�tO�!��W�X���p��cr��}�;�`��ƺ{,�8p�C�,�g+'����w���/�F5������Uě�.Jqz-�P����:kr�!�0�=}a�O_N��$1mй���Ȕ!�<1�Y*�n�gbS�~յ~���uф�â��^c>�=G'Ǆ�u�xӫ풐���e@+��S̬����-�\�ʢ�������a^6\Ьt5썸�Nt�	�lţq�A���k셯�1
�� �U1�&B�Ю�f��8B�a�/���^5��Й�0�;�>)�K��超��-C�� 0R�Д&�"�鞍��9�^�"R���󃗼�=���'��%F=L^o*�"�F�:ȋh���Y�Ԛ2�+�U�}�j���i)~�s,x�Pa����`T@�P���|{X�4���"��k�`�p��'�9\#_y��+y(q��-a�闑�++���t͌��G��U=�9Nvzi5����<���Q�%V����y��F��h�^�s)����MޤS{�wM�9j��R�C�����Z]�;:MV��H�jY�C]t�7���ݖTk���j���A�Y�z�X*<)�u֗M��z:��/un�>�MmBz����I����5�u������7�kNWNn���Pt�6)h�Ӧ�b�7�(��e��,�ǋ�;UX݉=#y��A�=ۯ���]�-��ċu�B�Z*#ɉ��62�C6Qq7��
��I�sc�1��-�FwH`v�#˥\iO�wE`+N�0k C�&Li@��
t�hX���������=k['�[z���t�s8B;�+�Ӵ��C)̞�}AiwFR:*�t%{��ZR�/<��0a~/Η��(��A\�y̎؝J���p��BP1B'���ض��T�Me�q$�h.2@v��B=}87���9C5�2ȇghl�7���,9���wt4U�Z���ҫ�� φ9��X�Қ�|+á��`*����f��?fQ,�u5��ꓩ^��g
E��q�h�+�p��.0�����p�pg˗���;K��S�c�:�a��"k"��Q�N"C�$!nN��]X��,ׇ�`z�ۼ�+h句vt]|2��g
r��X-����^�H��ʐ�s�`5�kM�8F%f&��{Xw��6�������G�{}�����1�09���rEYQ�1���:��v������CM��r8]J��pVO�97�����2����69|hn������nv���(W��Z�&�jvX��y����wJ�YS�̰�dYL�{A��e�d���*��5�xyfn�	q}���Gɝ�7��$UyHȘ�n�UX��a��L�ʣP���.b�i��Э�� ��|�=�s ��'cQ�L\.�e���)Ȉ�����`6ٜ3!xJ�r�"��=��^.���]T��+׹H��S/I2�P�$�LH���c
	�^�3t3�?S/B�Ą�?%�^���W;^O�}x�tdYe���eL���{Z�G�t-��"^u-0--�ڜ��5�\�(��f�1�m��%��٢�	��Gj=0������*���*�C�«�+y�l�8h$�r)���i�kw��2�j(\2:���2�2�Б'�o)Lp!���͖T_��aH�m�"��kv+��}B��aq��_/e�e[�=���ǁd_h�#^Kf=�*�(��w��Z���4��F�DH� ���÷s��_�׷W0�޸2��:��<��v�q��Eۛ,��V,g�K���XF+�wLs��djm�]x�=�j����i:3�(�uHߥʈW�,�X�\<��'��G�K9y��i(���ذ��S���iny�!'kr��%ei�@>\��ؼ�z_tѨ̮���%�'ld�O<�keG�w\���|qej�WH-R�(f���{9�+��䷰wa78�)��yI���wyլݺ���L�*w1����G�_�[���
��C#�%D"ȝ�̥�ZTB:%ͨ�ܖn�cO�>����Dw	=���e���:J*a߇D���
�s�H�Ȭ9�7z��d�Κ�x־�{�=�}�x$��V�\�����ݾ���̋�2�Hu� �a$G�3��Fj6�a��%Y��&�l\c�A���S>�Gƴe�sƯ��nٟN�T��F(C&a���廎�Ě�����'��tC�V�
��V6V+�'ϝa�L���6�k�rI�y4�0�ӊ�|��כU&�L߁@�¿L�&\��(ܸ��Zi��x�&(6�)�f,֎���jVV����`ta�1Cz\�K��	G�L>'D���w�q�������;R���Х9!�\v�Wv��i�dp;^OCF"�9&'�ņ��g�;6o��e\�P٬r3;Ρ��Z���Y�7�}2X<Wd��<�v"�qC����.L����o!�BN���[���y�]#Z�Ef�0ldb�'Ơ��q�,N�<�u�܈0��F�����(����^|�T�o�^�BCO��Cs��6{�k�Q5�dP�^Ġx�������M����Y���X�h���9��X�ǉb�)���&cѲa�G�bWZ�9�u��#]]�?6�W�����}�mtk��%f�i�/2j����öT�k4vg~���3g������T�T.:�Ӟ�$^�@���SD[�n�Kޜ���\z�j���ӎ�$PKh��z&�(N��3�N�ƭ�6&�� �Qvs��
�L�P�.��f�uGf�#�(Ʃy�C����[*���e����ZPʝKC�9���>%LUN�ʜ��t��oj�y	��e�%���#P����.�p��C�5σ����N�u�jv�6�ol���f��.î�Yp�mCaD��`��d���*�`�q�DX ��_x���Ή�����k������6��d�}oz�ùu�[2�c�8X,�p�ͣ��v]Ng� �^wY%�#�0�W��WOR�vH��T���縟!u\�R(ڂ)���ۼ��談�)��<��5�yz���=���υex��H[�r��	Ģ\�F�ܨ����"��3>�'�.\�8d��*9=E.�=x�?�Ϙp)�=�-�Q;ג���c#M`���D@J��u']=���	W9�1�XS(Y\8H��r���mMյ}��r*D��6��]�+@Dw]�*{�=�;ۢT��j�7�����F+�sׇʂeiw��@��٦�*U����[�4ْ����3���k��+�C��W^��'w`�����.�l�vE���8�M�U�.�GbV�,���<�m�!��F�_v��gC�`�,]��`\ׂy���5	��%�|��6���|s;R�fz�&+��^.��U'Ћ����ᘆY�*K'�Ε4�)��o���+^+����������5���xng�}�����4���g�jŹY��w���ʫxI�n�F����#�q�YL�e:fv�:l�'�qU���XZ�
�o6&ʱ(n��^�\ޏ'x-k���>N-�V�5��M�*P9���,�C��w�����縭��B��Ozs�8��j������!}|�TF|*�T��}mu�E�G[sJp�#)�ܫf���=ªȝ�Vy�,�8:�Ǖ�6İn�5풐����B��bd�"��B}��6�n�o��ʈ�oK8���ΫH�c�W��]�X�l���q���W=��%��IM�mn���6��8@��q�Վ�ER�=tf7��݉�o+Fm���'�1f�2!o7�r��U�k�K�HV����O������:�{�4�����c��`���*e�o(���\�����`6M)�����s7p{����ZFی�%����:�]N9���(vaq�WFs���o���3���cYG��mwI�+���f�h��v�t7[}֥��)#xgt���+Ter����M�1��aL}z:�]BP=Qس,�2��L(������TN�g �vG@�����uצ�3�<��q��{Aח�&ϖ	(r�X�'Y���1 �3�j���gP觽D�.��-���ج���2%�Z�����T;����k`��J��ϝ3�4��:~̐z.��J�Un/Ũ���ftȥ(Á+�E�]tl�g���y�5Mf�\c�"���7�H��:M�8:��N0�PWl�J�P����ńW9��w�������%���5�����V�6��/]��9	
�u���1�,���S)�N�^�&���?��&+����5��̋�VZ~>��� {S'u4Ȩ����t����ewN,�79�e�7��a�1Gi^�K�e�	��s��n:�Z���{l���͎��w�'�r슰����w<Ʈ�Ȃ�z�A�Q�>�pVNU-Ĩ;\�,}�U����n�fs���%ak��V��:R�ˊ֫�m��ؼ��p�2�(rk{&���9���s�'l�N�r�����l�Kz����7F,q��ᆘ�!5�L�a::#�י��7��n�$4��m����qC������	e�	��R��W�\��U�s=`=�:_4�na
u�{��Na������C������q~�I��N;���;��D�`�EGUq}Ti];U�@���v��}��v�n�2u^_�%oq^�p0769����m:���Ւ��k����}\� ��o]y�VA�@+��a�謇qJ���͵O�tձ<k���	�p���(��2��5�DL�Wu_>�B�򫔿wJ!�����:�Yцe6�0�Dv�<qB�c78�y@;	rb�넪$�6����Q���:��B��vT�2��.mC<:4�ꊝ�n�<���{S�Ȟ�O�N�v�^6_�g�4z�����>�Pk��ð�����c/5onQ�_�^�7Nsb�ϯoܯ"(bT�TSsFAe�ojF�	'��羒�p�_�z$��ػ�;귵/L�<-�^���C�<��J��&3�(*�~�X�$0����lZ��K��Be>$��ጳ��-8붎_��ΰ�KW�t���
����䘘�pkHdmoJ�����b��{��4�r�X��}<C�X�>㠠�Bzb����:�k{���O}�[���񬨂Ĳ��#�r��m���ig[�7�*�Y�k!Y�w�Wi�N����b,J��!ǩ	�WvP;��v��*�L�(��̭�.E�E�8r�3�#+��]�Mt����V3��m�������*�w;��y��(�yԜ�\|J�u7�6���^O��|��0B�8���A�����Q�����[�f����d�M�1�	��a�zY�&;6e��9P����i=oU���֣�1��a��_n?B�����SFE��j���46��G�)�=�r����-�ܗ3�?��7&G�H�L6�#
�6UF�sa�8h��1Q�i���W�3y�y��r�g���T/��6S(f�@�F�ʪ�An�ٯ9�����R��`���Zܞ�se���w��=eh?d�e���{g�C傽��2.1B���E���b�_u�кV��2�E�.�V��<�hu�ϫ	�=/h��OA�b��:������MX.�>}�r]�ذ��u���e��ł�n��x��P�^pF`#�\�-�ێ�X5ףeI�\�{p��997��3F��-OR,��Ψ|	�Q�ԇ����WB�K�ٶ7;�CڼI���q�dk���gT[���gVs�}"���]q����tAgG�b:#��t^˒�a����*�!�l4����;��3jKg`�B�qj*�C�<���r)����*z�����r�c��N{(w��kd��O���'zm�q�U0�{�h�8Z���+�����Y��D�X�(<z*f���eq��{�2�K����co�$�����ԗW-�,�|L�7��[�H���-�Uf�n� ��/B�D�ة��Y�;4K�メ���D��+��Lo���ع�YM<[bo݁B{�����ӨNK��/Qc
�.������3t��U��K����Y���(-t�:Cz"z<�:�����Aγv�@b�{v��s�pgY�i��>�F���5�7q`U��V'��G��sQz�`7��:%�Z�}�G��Y��j����*w�ϜE�9��sD��\n��3����|]�KQ��@]Yug7�eI�,���w�ًd���G4�;v+M�.��k��xL�M�ׯj�x��zr�Ǵ2��7j�ɘ�{[�ol.���2+H�ш�UY���v�8C��RV��J;�����.ƻd��t���n�)��jmJ�YQl;�8�/\��ú��de�j��y1��,�*YL�o+���1;lZ��W �/y��C�n�.���;fvYdԍmEz��]�s�$L�mqܑ̹[�u���k(��:�쮶���}��Êe�W�ZB�c�aͼ��8������ueXT�l�.�J�K��s��->8����yMf�9�MՑ(�1��>:e�ڜ%F�̮��?�י�Vws-11͚�t�d/�s7�;�M�z(WV�=:i�X�K�3x�r5�a��0�u�za@wҕ��ʱ6�1��,�s;���Z9�:�1N�d|�4�ҷ��(���������Aj�1S�6O;֖tZ��1q��2�WV�|\�@�4 ��nL�O ��ј��6[r��r �����@}1*@��Bң�/�C�lh����V^6�8����5��vp&A�$���BG5T"�Zc�K�|3t;�)`��b@U]p͖"A%ޑ�����ަ�VCP/3���]ė=�fK��d֍�@�Î��}����]ۺ�g��V�u����F ^N0��`M_!+���Z-q�u����v�IMlJ��^���9e`؂0���sW��\��)���P;�e>�/�<|y��S�+GmB�v�tk{y^և�V9L]�M}���Cĸ��V%n�\|I��LT�;@���n�4Ռ4���{�5���R�ڃz�'Ë���Sĭ��F�l˱Z�h�S|(p��$=�\.�5�T1�u����B�N���a�5�+�ie(^쮕�6���ܐ��,�7��:�x�Dw�<'	��i�es��U�Ι`�QؕӺ�-"��9��aס���qhrIu�x�2z�)r�M}(�K���V7��v�2v��s��ӹ/o�e5��S��pG��E��n>ض���]N�8�x��t	��N�"�۪p�����8�V�Ɏ'���V#�W⢂%=��]�ugp���j�F,bm�1�<j"�q)s0�V"�T���E�T�EU&�N�X�-EZ�hQ)J�@Ct��YJ��,�[i**�ՋR�ۧb�Mf8"��Q,�b�D�Ŋ��Qb�K[`�(Z-�m7�G�D�KkP�R��QA+JŰ�V���Dr��kT+B�Q��ˑJ��X1�іЭQR�TDF-��ET�Q�X�6�Z�1UTĮ�M���kV�1�����ږ�Fʕ%Xٻ1�u�D�e�Z,����"�TEkF�V�D���f5�
��-.�m�Z6��
�X���V���i�-n9�֭�k-��V(Ŷ�5��*�b(��V�T�U�U�[Z�-��EjR�6�FZM�d�� �"Ĭ)-
*�[c�� ��A������5�{<:�mD^��[y.R����Tf��5����堹]�Rm�Ǌ�$�������M&pػ����ۼ��J�h§il���!��}aOMtp�T��Mй��;q/lG�"�#	�X��͸Vd��#hF�te|
a�\g���kl���Q�s�1�np����n�^��fbKR�Έ�$��THu�E ߥ��1=^��a���k��V:Q�Y�c�3o�G��j�"�R�0�)u�A��z�U�)f�4�=�w�
,S�3W��3;�
�w_T�r}������*��GLO�����lp�h*�f��.�>��\N�T��2l	�}���K�e�tȯe]��naP	���Q�#���œ�b��ȕ9RYxeV���b��!�T���MF`Y�ߦ^F�3���x�^�Pf��T!} ��v�Rk���#�]�^�_wx����M��#C�X�4eiy����t�S�lnM1�:G��7��^�Z�P���o�s�����
k ��kG��ki��^W�Ƀ���k��2����g$�Fwi��HӐ�c�=����.�MI��/L�� ��A�8����#&)��eJb�T4ٲ�~)@Z�s��X�B�7W�V���0JIU��a���6wj6���cb��ܺ��C92f�X�ڱ�j'2Қw�e��Cv�]�%��c��{��^i���i�¨�NU ���!k�0ym�rr��+Xh��q����fj�[�H��\+g+���6�0i�Qp�"������������"��Y���؄����A��b�a��iB�=	��U��*t�tnC��O�rD~
pk���+T���"Ӫ�4�J��>u�S���:��L��;z*E�X�m0�(��� ��Hf�fP�J"��Qǁ�E�o�2H��J��թتn�m.�M�Q�7�:=�d��%Q���%�\HV�=�����U��s��nH���F'|�W-�C+oU��PS�C�t%J]#�!�:-U#bb�b�����*n�	3[3G��]�޺8N���j3�$;��D8��!W�
@�r���s��r�sT˭�/0�������y��h�(܇~���j�M`�H܈d27�M*��O��f8�c)�I"zU��v��7"��'1���{�N�R���M���i�b��b�AE*:`7h+���3���o
�ؙ͗����b*YʱԈ�vY�6	9n�Em7؇U�����7�\͐{u��N��r�b
cG��S^���?��񿰅\���( ��6s�Õ��J���la����CT��1����k�{1x�H��CX@�eܠ5�:��EZ��:.Y��9���3��x%n��Or�͘1i��e ���K���Wk�s�|��λ=Y��R��}��+]�_v���]�q����}�]��S;��4wT��������Ze�����1�ck�e��=�����W�1���3���]�X�tk!�xy�>
����������S<VF����A�Y�����c���ߍ�xu�U��*���yۋܚ(Y��t��y��W��&��I*GmQ^i���s*t50bF���9��#���b*z��[˭��Q]���9���=0�Y�s���*EחS��u�<s�g.*�T�m���3��EڳckA�����i�����s�
�U�p>�͔T_���s�/zl��)�ӶXe.����U��{�8z�Ţ�z�t���N�8z�k����p5��N�G��ѕ}���잖�(=�:��,U�49	�T�����nIY)�d'�e����z�s�۪SX��C�+emi~ٖ�q�!�9���.h�ٔt׮Y�mU�e��Ӛ�i�F�槉.�R.�OwM(�2�5�d8��L��3�ޞ����xW3���tz�{�6EgK���D��ֶ(�-�L;�xƯHZ������/��'o8��$��ܫ�74�](�f�y��VM�)�0Z{y����M��1�΋����r��z\�Z+�ƺ��g��.��l�͒��F����0N,S�Ԍܨ���b�|���돵�#b�T�g<�:!ǫ5U�p�j�g*3�����<�5��q��>��WN=�������`�k�����)�tX��kЦ�J�*8ZufE38��Mn�xՏ>�7�d�k,�'C�6OTz�WDy\�y�F.�˜<���A�~Q���p�9�gf+{�_n����j�*����2%��l���3��*zb�8Q�l��,d�qr�FP�s26*�1��0
�`�S��8s�T쎬,y}�-1�>^�
�=�/^��<LI���ړƲ�X��D���AC$���7&)7Pei��&�YɎ�[����Ǽ�LL�ׇkz�L��Z�ףD�m�I[�X�ⓜ� �� ��Yo�w�[{I����f��6�Vl�t�����H6���Ԯ(���鲗e0��{���M���&�Xa3/�)�!��w�}��wYlX�6E�́�cX-��ݬ��~�����ROK�7����i��}��.���t��ZO/Pw��T���*�[0�z�VF���z=Tqd�!C�Z��c7:̕pF�xhܯ:��{J�ПI��*��E��q�[�R6��ߍ�r�g_e�h%J�%_�5�[֔�y�;{����C׳�i��lN��Z��J�:�_Buw%�i��8(��,E�CiZ�>��3q�̡m≉;�kV�!�yӪc[�ζW����[´���hu9x��Y@<��즲�6���u���q�dR�E��.�=��f�!�̩V:F��P�@8���ȵKn*9��kj�n��fV������q�ㆹf��]�]8xx�<g�<���|5�chա�Y)��FBj+�K��9��=������ՠ:'�O6�\��/T��|zeS���_[}y�AE�A�jנ	D�[���箻٪Vr�go���}�r�r�{�I�	���?1���|�%z���/`\)�D���b��f�&�s� �� �A�}�_�hֺ�ހ�ݪhWK��*GD7�e�=KIu���ߖ	�	�V:���8C�����9�.��Y��y[6<��`6)K"�*Y���VB�!�������Y,�@�������z�(�)r~�� ��]������I.c��!�rod+����H0��7Il���s���qW��8S���B>w��B,Jsq<ќ3%�E-���=��o��򰽸SW���M�M��v�w�����َ"F�¢����b�ƴ��W^;���s�7�0ҽH�*$�uI�8v�P�{�-��m�s�gS94��/�f,w����o;3�\Ǹ��]�շZ��u���_;}}����*M�*�앶r5��z_�dJ�%�g�M_���4�$X�O���(��g+=��9�̄n���0X�5eiy3�b���c)�;p�ѱd1]"�����y��SU5j���|C.��7�I����B"�j5C�fż�V�5��w�&2/%�#r����inI�J�.��46޻�7^գm���j��i�W�ED`�E?y��
��.ʼ���;�~l�*�
���eŻ�#_K:�z�J|�+��`K�(Vצ�e���>�_�/[L���Q(S��Z�ݮ�Y��}���ٮ�U��]�YbQ�R��\�)�p�Q5�	���dWp��b�@b�q�tf�r�p9��V��mڕ��!����ֳ(e��EH��t���G]D�h.��QCӔ��ԫ�%c�:@����ݯ�c�W��U�ͭ�w�Ж.���,�j���*Ƿ!+��Bx��g3=Z��T��z��;Yܳj`2�e�c���p4�C	��A���6��a��Jy��
n��=Z!i��Y��/��I�2�r�ۯ;\�"�tx���n>с�W�&��E.�r{ݳ[�Cl��
�K�3q-�h�m;�5�P�	�x��`��Q4�[�ɪ��Ӌ�����F��]+/��ݳ����Cְ�>��ڥh��$mv��՜z�qS�]�F(̝��9�j���,���g�9q�̨y�)����+-�7"@dk�4��WK�b]�EH��*���?9�7����j4��V��j(�2�ᑢ���
^������A��~��ԍi��x\�
O~����Hm�2׷^�x+�v| �l�"\���՞�r�^����|�ߒ�u�5�XV>Y~��q�d8�8�o�c�E5��t��m;+ss-�ᘯu`ϕY~�&+����5�Ⱥ�o����}jz��<w׺�F���Z���&z��&�{�ڋ��.���.VWü=t����N6O)��#q��
��栱�ج�8�(�AI.{j���:zJ�c�j�Ȃ��bp��#��3��{���%�9V�Ky%;P�y���"�M����U��:l&��b�i��]ؿW����]	���}*N��Z;u��8���`�0j�iUe�R5�6�Va���PQ�/V��F*��]׻��׵,`;��y�X��u�Y)���W��o���
�hL(�wS(je� ��#�ܖq��n�*P��UN�'�r�"�@��UFv6Y*Գ���X9�vGh)
�S���8�4�3�P�9���%k-f�S[R�ԃ��ēU�8jFw~�k��d�s����䭉k�j^��|0L���ŒF�)��/�݈�y	A.��'9��SQG_�U�jg���B!�r7z�v��:��!;n��(����M�=�^9ǜy(^_�<d<�D���Cf;�iB
eDW�C��/���t��d�=����F�X�oE�:��Y�4b���5Q.�K�[q����:#uzB���.�2�J����>�����}D�5�����o�锼��+zY.���[/�L*���z�e�R������Ί��x�^�$O��1q\�]p���L���ƴ#�����1�4v�<���o�ZGM#!��Υ��ʈ�F�[,�pMO�fy]�?:�}p9\������7���+bq�;U`������;,U3~(�y3�Q��ɋ98�'�v{�I�0+�^�%A׋wI����W!A�.E�^j`܂��y�z��ԦZZ/���o�����+�M⭹�͐��ͫ��e��Jΐ�TT�H�ћ�91�$<��=^��~x/p�8���g���/�����Ϟ'�#���lv�#s��p�u�J�����3;�^�$I�l�#Tӹ�w;��)���:h\&G˒GB��x�{ّ�u!�mWwKŔ�ú���(ZfnQ{@������G��w���9
�V�������LCq���A+ ��yp��2,�tL'�H�B��<�!��7��מK�*X�l!������%�FnUEf� o#1b�>�qEk��\�~媤#��rw�w��X#j��� 46�"�T��3����
sh lP��N7��;Ӊ�����E�7���t��r��
�����9X*�0�u-��2�xY�B���C�cu��V�7����*烲��z�n����[<�v_��n��a�:����S�H��GF�{��47�g��j��:t�Eޡ�Lq\%e��(���uNaH�T(#A�u	��Lؙ!��yos!!�)Qo\��7�Qvu��9J���F+��g����7"Qi&��Og�z�`�9"�hu�U���8���,����W��Z�t���0	�����F����X�r��z]q&�B8O��	T��ީgVvH�G}����f'V�r��w�:a�Y.�yf~�hbz C�7�(�	�t�z��r ���KO#@]j}���{�3B}�A�vV"��r�z�Z��t^~���;�mr�a���6f���@k�}��7�c������r�N����I�T�}��u��w���[#�T��[|����}]�U��p�sv	�w^~����r��=]:o`|��l8u+Ԩ(����p�=&/-
̧�@k�Gx��j�bKfr���mn�T��uC�LW���n�~�,��*Y��&�hODz���>��k��:J�O�������b�/#U��`�����Qf!��{8�d��]q�g2�[�M��2�_�/N��W'2xS���z�=Q�hpr�.Szl=Ȥ�{�c��瘚�����n`"�ԅ���z��9)�vj��~�A���T!} ����Iؾ�]���v7�7ж��V+Z\���l�dBX^L�l؊�GN	r�tK�C'��[4a�[|��Nr�8�Ɲ\����Y�l���E���#��������Zra-� �z"��үs�n�fR6���5�*�j��^l�>�=�8^�����Cc����0��jd��ؤ}=V�Sb)~�㮭ܿ�[�
���ղ�F���,�1�%�y/ ݭJr=��ID��%�1��6�P<qB�@oK8��-U�i��+���f��t�/���c�چ[[[U��tѢ�ˠ�zd�{�<WS��t��u��c-�㔨R�P,-T��o&�\#��W}{������jYW�W^@�9��)[5!��uȤ�P�3��z�V�Yq\@����ss�j�M��0��ۛ�<�X\�u����0�9eY���'J�߲?�N�jU�iI����5�ęݬ���F[K��)�C��R���qAr�����q�e���(�+ݗz����Y��e�d��Z���2��}������k%;ԑiu��:���o����佼&��ʂ��m���/9-6N���un7��1�atBcwQ�7��������۽��1�p��9X�삮�p[��Hsc"�2��{m@��}8*]X	��ot%��}B����]H�-aNW���8����֠7�;�z���h*cD\�1�C۩u�;�S1��.�
����<���i��c��*=r��h���y�Z�w��{m؛�O�	"A��A�\i]��ɵ����z����j �
� �7;u�~�!f��۲�ӄ��ݏ\GG��-�BŶ�kOU��sW�f�Vзx����#E���%E�b�ʱ�hqg�φ��x�7��tq�I�W*�֬Χ\��Oj�����Nmź�|�8�MV�]նG�+H.c�K�Pׄ�]��������٘�������U�X���1����uU��KAҲkt�=���*ئw���t/d�i&����m޶����_wG�2*n{q���1k[������}B�N�N�ơ-0cU��S}iȮ4Th�h,��X�Nɠ�h���Qf\:�㪹�9�p�0'���.�L��aA#XU#E�,I�ȓ���	�(�$I�s�Xa[T0�ZVrVh��&G�v�P�:L2�XJ��4-��,�Ɩ"r���	Ϟ��F��Fj�%�Ғ
1'QD��%'��2���$g�e[��r�y��S1}��dֽ�ʰ�M[��+H�,��OXY0Q4:ڸ���M��+(]�t��cj�h;�d ��%����X+��yJؕ�I(�;]�g
����J���hh�<�p��آ'+[{�|��+X��\�]�r��=�����.�-��)ԭ�t2<�'pY�y�vksŴ�:!�Mu����]�Wn>�egҲ�B�lN���y�q*��y���X�k��l��)[���I��a����>�ˈ.��0lH�bg�n%&�'�9ӥGoM��ɓ�v���Ɩ�)묭�ޜ�߅b �T��#��|K�4�}�c9�ݼ�a�u'4yU��(8m+�|��.�:jNT���u��U���s��$�;���۫����v2���<-�f�V�fC�]��I��,+I��e���t\�\������u�����]�t5d�H[���_Rۗm�4�*Юq�tt\,��w�tM\0��d��!g���(jGbPL��UTG��`�6���qeFƌ��ډ[J����%����iB�Z�+~������iR���JR֕H�r�5��(ZZ���R�mvT�֩B��aich֍+mcDZ�w�\1m�Tmk�im��J�u�WZ�%KZ��qb�)�⺸�cF�8�Kmj�֙pqS32�M�LDkQV�jYijڍ����-��0�Tj�h-
Ѷ�j�,R�V�Dh�F�n��UmQe�4��ִ�5����ekUiPkZ-PPl[liTFY[F��R�4Y[V([UXʭ�4���l�际,���F������R���sa���cE�(:��Z�j�J�p��G[c�b�m���ҴD(��j�-na��jX��-mvܲ��bі+*-��,kM�2��b��h��V�j���e�Ym�Ҹ�:��"�kE,j�-�����wos�!s�J�]�՛��5���f��-[�Fs(u�-c���`|@��+Th_����o:��Y����;����TD9j��U�2_D�n�� 1k�\��h�+����/ϼ=]׼&���P�:lQX"�1�S8�L���V�-B6��E�<������U�=��1��;#�K���6�K��GF|�D�hu���U�����+���F����u(9�7;P$k�n�2ȇghl�g�mД.���DK:o�e���m_oy�En���Nb����r}k^mF �*���U8��~��	�q˦v#9�e��=�Ъq�{e����QD&&Uƛ�/#�B�f�1����t�ȋ"C�$;Rt�K^tm\�*���G��D�j`z���97�`,z�6.�)V�b%E���8�N�ȕ(�fՉ�9���/*q��=٨����u�����G�T�� ����+��,�'�<����U��}����jG�K	�a��j�i6�����~��x�V�V?e z�����9�㼊)��;�qdᘥA�*r%��F��m�\<��o����}1f����}k��%��մ��&�F�C�(M��EG��0��18���M�xp}4Z�-5���2�<9{�.�7�o�����;���)1Ԡ	3j�Si��h��f�����ʞ�,�oGw���s�<|!�b�ƃ��e���ț8��n�%ֳ�䁫�rWh<�����T��滩7ҧ�ݸި�ݓG������ж�������ݩ�(؉����E�z�OJ7e�.LU�W��u�S��42��f��"ガ-t���=��M����錜��p�O]�q�c�z`�b�yq�QW��]SW�8`�͔TX]�����8�ެ!�=)�N8�,r������}]8���l�cݛ�]n;ݪ#�C���7)��G8Q^W|Qy�Gb�dH�ճ:n+�����:���X��?pY��E����U������<��ZH�,Wu��
�)7F��}u.�nY���⋡��k%B�NEA���}���u�p��y�:c^�u��׏oå^�L��k�
:g֥�<�D��Ћ���J4)�N!�t+��:eth/	ي5[�-mD�Z�C��;p�Ω���J6Eb��٪�t1���"���h��!T�U��^u���]�����k���.���)j�>Ns:ex�1֫Ȋ�.�r�-��>�.iQ3}�9��>����{H
U��l<#�U��EP�ĹhB�p+6��4��<��:P2GLDF]�7��쬻G��;�?r�����Vo*<K��0�d��Ƣ���2�us�⣝���z�/�}�ޚ��Q��$�=!��
�ֹE�����F�\]Y8���d���@������ݡ��IMw�%wM��}RM�=�K94��ɦ�ۜ<� ���K	q�.|p�]x�U8Εcgu���fٚ}��ڴ�Rz���D1��mx�U�mKؑ~�L��b��{&x�*nb�w[�ý��]�U׼
y��OU{$ˊ��Bb���X5�Ɋ��Pt��E�;��Lp՞�'k�/�,qN�����5q��/DIB��%�ޠ��R�"Z3rb��I��aޠ��7�i�Qs{�Ж�:(=T��~Up������xt�����v"�2,�v5q�7�0o�0�y��LE���'�//d����lجt6�2*sn�8m�qx;i\QMGZ�(��q/vE�J���ݫ���A���"o�و�9U<�0K~�M<��V�x�0��W �"*�e�Im6=o�����sUW�����JqK��[�o�R��������d2�nwY�����Ib�x�cB.��xeVOk�a*��GS�R�u=q�];m��{����=AqM��~����8���RW\U�+m��ĥ�-��M�<
�Z�C��F��c1�Yޭ9V�.�������I��;_:�ȕ��ժ� �ǎ�>/���"�T{��@[h�;�D&�u�e;�y�`+��a'6q�J�V6��ES�\�P�n�_k�ҳ��_n��`������E��3X32�	[�.�_.��>�����
oJ��ɩ���8�E�ͅ
!�P��t���E�{��;��s��y�԰1����w��δ�q�uȝH����q#�J��F�N8�rά�;'����w.����Ov��v��rAd0t�J�$ߢE��M�쮺:�:�U�׽r���B�L�Q��zܲ�n]׫RG�h�|5�:��8�tEK�9�EЎ��Vo/J����ӝ�o(gM}	�}3Ǳ�6�w���&\:�J���ߥ��'�(]:�;)ΛtIe�h�ܥj1\&�vl�b,���GLl�l8F�E���"E�g�
�����QJ��k��u�{1��9�4/i �S��,���V
�p�MR��bJ�3�[ٛ����
�3�m@y3ѭ��;��(���X�郼�йYޛ%y�_���h]��gU�
�%�l$p��o���9>p�<�:�n�&g�V�>��C��5Osj=���ᔐ�г�	��v�j3Ԑ�/QK��/Qz���*���d+�SP�H��6�l���3UK�GHQm��98;��c��0�m�t�
�.�f�x��Y0!�X
ab���*��Mx�J�د�M���Gn��QS�����U��v�.�&��KS_^FU湜�M�EH���q��H����|�n��ɒ,}����ޗN�<���6-���y�Ef�;�V9�p�K���m[�p�wg&�i�C'�$�]v������罫F�W��-�i���Z*#��:xB���(Ov���.[�V�����ϥ��w�k�g{ͫ{���U���l�i����n'&R�\���k`17�bM�:�<��:`�Z�Dqf��ũ�#��W�&-��ǻ���۝ItS��s%��3�X"�8��!#�x�`u{(��(��AvW�k��T��G>�����d-��>o�%�.Dl-<����}�Gjq�=:�̯�лt�}�WR�꺳����ބt)�D;;Cf3�K.Dp)K�v0�:hZ�����b�W�=}s�����64Dc9����$�w�8�3}2�(	��	�t.����{��V���M��賌ˤx�D�\a�*^GdJ�fۚȫ�H܈�8�zD��H/U�_�Cƺ��\�Պ��ŀ��c�k��`z���r�K�J�q`�pNp�Y7N[��y{Azo&+)�a]�R��h��a��]��e	8�ݕ������oFܫ�.�Il�C�n� Ga0Y����p��?/��@�ۂ����7��� 4q+�o%�P��i7[JI0n�u8��]W�&�3�k��bxpJ]ӕkE-�����$Ԥ�}W�4c�r$�@ڣ�ʞ���C=v�"���g<U�b�����{#�����f-}<������c�p�uS3��F��.�-&�5�QL\^9�xB5�w�?�6��1�y�a�a�ERӽ5�"2�H�
U�ߛ3�aHf
��g���
�n-�\<����u�����Y�כ��~�4�Y�#S&���s9�&��~�1ʳ>(5��fe�H�Ǽ�}ܟ���������rh��e�[TD�	S���ݩƦN�����_�
��rr����q9sE��D�}#/�-�lI@���ua|:]F[�t�[Z�������O�K5����+G&�г�e:��Fl�o�q�
�U���`�͔T_��aH�abv����3o���E,HoWv������{����1��5�)E�+a��_�k;S�T���ؖ-,Q9GK���Q[�WH,��ާzO.�.OR�꧐1���܀sFa�=Բo�`�
��e^u��2�N�E �:���~pe]%���z�;~�O��x0�K銕�oo��+7G�ޢ��v²7Fp�ݖ��Q���� p���]J���5��)c27�r�V7��v"-⭲��}81��יc�c�Eu9�]f�sX�������ɗ1����x4	��L����҇7u����i�UͰ�E,���1ё�ڡe�P�9%���ݚ��"D��d*T)�!,�9���ӝܟ+{Ӧ�U3r��<�J6ER�;a�1���8[��|c�hN�6�\��ǜ᢯�&.}��*�`�{/���OM�g%zf??�o�p�;���d���P�����{���{2��u��
2-	$HpʰeRK�\�U�k��LZ��AN�=�ݐ<�Y��k;��m�zHKШ���Q~~���?�R�_��.�l������SU[���In��I޺��ۓ�S���Y����5/bD�f�b��B&J��G�G��\���]d����wmGGK��$azZ6�TO0�k0^r�I<!�V:�x���o�����=�G���ڵ��8�%�^��C��HЮnLW9&:Bp^�EF�̝9��qޣ��1>:/�v�J|���S�C�]Cq�X�%`�qEr#�?Y��:m���2�R��[v2�#����;�6+�2�2(f� o#0E1#��-��;��= .�r}W����큺-��P��z�=k �_T-�KR�}�>�k8��AK/��L2�*ːx�!��T����m�$��V�m@����.�������ӭ9A�Y���d�:���[����br�?}UL��zg���
e�L~����U���߂!Wuc�1*���	��S�V��V!�΢�Oڹ�Ƀe�el��yT�a�V�b�=NF^�®b��KZ�]힡,�f�9�Mf�Ӽ��>��S����ы
�j�����}����P��nB!Y�lj�������Oa]n�a~�B�ED.�e�W�)U���N�.É�!�̩�<	��c٤Fɏ}��f�{t���,	��^�x׭ʈF��q��l�9E�u֋8��������Y�{���΄a���g]�.��GdS�2��8�{=n)�����;�wE�^�Uu����s�]��3Z肈`��\�(���5����kf�&�e�+3�d�X��_��ގ���v'֝��S���FY����f���\qȿDQ=�܉z2�n�Ğ��ڌ�[���ᓖ���i����#�3
�\���7�f��q.�q���8{#�_e�Ht�qVq��֙���6lا:b���W���1��A�^���|��jX�ռ�z�0�^��\��ւ���ˣY*�����r"�F�C�l�N��kFi��OgU�]m)qֆ;��'0&��O9m�5#;�j��Q�9d;��[�X��Y����Nkqwp�t�Ҿ!nf�Z�ow쎓�6�W4Y]����s�~�W�G�#{U���3pE(���� Ď�
�
�p�p���{aT(7�a�)Z�wt�X�!1W_�i��*�u2xU�K��=�b.^���=�����Z���̻zL�`G�h�\����x:�Km�o4�Zz�GSGm�u�zg�Owڕ}C'RA��%����s=�=d5=�z����V�����:����]N	�gU� �j�����aP�_k��]�E�VF���`�j5�f�=�ӥ���b���f����{l6�lR��^�ײ�H+���A-��Ucq%o��G��-@��>A<�g0����;ۭ��~�Vb��	g��czYqn��k�g�ϩdq�ku�.�W�M�[��"�Y�c��N��&�:��m9`��R�+7��z.�u�U�3��q5(����ص�1�{ȿ��Q[bYTQP���E`�<FR8�L���J"��Q�K�wy|�/bW%���,e7l����R�f�\�@�H�ɔv�.d�5+���ea�)ŧ��S6��͹��i�Ji���d����iebĈ�V��]���YJ;y�+��1�1���ks��*�����Z|s�zۮ]��H��T�L�+Q�-wt
�T�s��o^�#��6�k̶s�&G;�p�x�IE�֡� 5�f��o{���G��Ӷ����әdC��6b�k
ـP;�)u�F e�2�աp���
�y}�LKŻ�Vh�UR���G^�'hb�Q��u��q?HT1
�F�Lr��#�5�3n���?�'eD}t��,нPWD��/�v�Y�}�.aw^\�A�dp�̨�-��ۙ�Z6���)��"x"���6�S�Ȝe�^���j��i�7��V7m���9��.k=�Vq�
�_;~�+�sz\zq@*E�;(�ge�$��t2+��}7���	�3��^>��@��=����l"��_.a��jZM���j.�bG4��R�"�^�s��7v��^ٸ��~��A�)�m��1^T�*�)�Gi1\+��"f�8�km�s�ێ�,vMl<$�AA"�(M �<E{�c𐺑�
����Pѽ��iѽ���3'�qyXȲ�U��=��b�{�����wꑟ$����$�uoTL��q��"v��[��l�@��.8*��u;�{"�#�]x^���[���}�uvQpֵ�R��S�N�i�(��[��[�zE��q,r�mv=����f�P�ȭ���܄^�{�����t�B�ewur.[�׻Q�����]@�nN�]k�J��ά*�un�m��}CF�'4��/��.cf9S��y���7v�Y��s�u8̻�E��.FG��&��wGy����ap,��u�á��>xucE����X��nl�=����@�S�r��m�CS��f��>Κq�h��W4({�~\�6S���{L}�G�?�9��!�M])5�-Ol�|t����Wk�ˆ�����B���1)�ô�L�Y��n��#���J�'Ř]�O��|�z����a%a��*ӳng�ukU�ř��D�-�Z���`z��o`#�Y��f�E�Ek>���j�K�_,C#p\���0�TVy�H�oWZ��
a=0�>m`��v���[E�7�r#ȥyw��k�����L�ѥ�2�ܵ}Ö���Eg��Ҋ��N��eb`]K˫��ɭ8��=y]��9m��C�tÈW|ONe�Q�`"�P:�X/j��] ����3��f7�ѦE*�üܮ\ۇl-���[{�;���<*�I��/KDgC�u�r��� )��J��iγ�E�L�T�u�������a�1���a\49�s�|�G˰rOhr���v���lWMt8�.c^�K&���@6��f�4oks,���搙�xU�$vqt!Wd�9�Z�{�T����=�]-�r�;����Gp���IځۧhWJ��L�9Y�I��Ŗ�X+����W��ю'��	V>5,�+ 
U�$1&n��qBs�]:;�0�ƠU�NKlC.�h�XAR�	����df8�)P�/�P�NXd���Vԗ�����b�f]0ѻ6R�fIB�<x�j�M�7�&FJ� �s����] ��^�c��X4��.�IV�cS�q��r5vj;٪�kv��Ҥ����Z�>ڷ��љG�ږ����W1a�c|m�5}���Yvj�:�R����eV�z� &���:��5�R@f���<�
��^��"�VWV�] �5�GmJ�p�r�uf��t�uc{���ѫ�Z�Qث����*t���ê5L�������7R=���w�ɹK5զE��w}-�'^b36�C��h*���`J�����u�5\�.u}����;�uO��T��\�18���`Զ����K�K���9A�uO�\]��7k�0�dÑ�9���M�<���5�T�VF9Ӝh��b��g^:�ޥ+�!�ba��I�y$�Իn\�����G�;�yb���Tl�3�%��|�Y�^	�5>�'=�X/���> �P�2�5}��^��B�pxuZ#�#�D��Y+x,��mnn!ܫ�YG+#�J=�W���0�t�Xhw���3�ۋZ�+IY�}�*;�������ѝ�BR�� 
 D�F$��j4����R�4,̢���ʸ�V#��*+�6�r���(UT��R���3+�mr��D�h�j�֨ѭ��F��Q�X�����q�m��Lq��k*-M�Q�I��(�̣����%�FV\�q
V���j�k[k+
&\r�̸։D(�TKB��kq1*E.��-ER��C+H��b[-IP�Z�Z�F�E�Z��V���PZSneĸ�ҨҢ[cj�YZʂ��f-JU[l+R��`�]�pTFD�X���Rږ�)F1*�ʕ(�m)R�)D��"�2��[KV,�4��iWaV���\�a�6V%�R�b�
�Эj�E�
%R�P�U+�v����UR`%�P�Z�P��Ѡ�m�Qd*�U�jU*���l��j	[u�_�7��
���:�7�0�fA5���[l�웤�����.�]g#�xvdɂ�����QR��\w�,�s�����R����=L�#�Nl��N����Niahڊ��P�1��͔TXWx[��4�1Ցo]b���ɐ�,�#�g0�o='�8%/s�]��=J�eC�*m,�X���`m,�P�A�"���21�w��U��"�-�lߝ���c���r����:m�⢻�e���͆H�Y�/�nl����3�'Tڝ,�D�A��B���:��^+1�k�C��{�ʪ��8Xꑅ
!p�Q��U��$�!�"�8��Q�eDS��}W�Q���GN�m�S�=�P,\�8�L)¢�П�O"�c����$����h�)EL;�rD\=�Ob7GB�\�s�7���h"vU,0J���lOa����P�|Y�����fKNh��T]�P��2
,�ɀQ�He��|.@u�	Z��C�R�9�X�=ɴ#�)+N��qR�Qť�U=���{M�O�>����p��:#e�l�>�wr��Tjݤ%���OpOgu�e:^�,���Kؑb�3��T���oa�Uq�4�+f�˕�TY����@��Q���zWv��-�n"�Z����oK�����\I���h�:��[b!�f0���o�R�(�"%�����'�<���YH�>�<�ʅ[Xeي�D]v�Y1�-��P�Ga�����V}�h��*,���k��t6��j��z�s�rѴ}C��XVC�G���DP�ņ��`�7&+���P�*��6Y��'�7��,�9.�S����9ƙf\h�P��\���TT�H�ћ� �)Į~����n�y����Y�1ٳb���\�QƦ�v(�~�7��m���t|3'�nx�Bڸ�iuaJ�`��\A^�ǣ��Yx�S�Cl��ͪ@�F8b�����v]���;����{t�(��[ўq�M�j`�����Ck�.cL��:o�LPu������ϱ+����ٞ�Gͪ�1ŷU��ޭ���\z�����&�*_=����_��ke�}���y��qaƃ{I���B�E�U�`�U���78��>�}�g��o4��;�6��Yq�R�5|'�Z���\E�U�����]���-F�L[ބ�6Z|��x]�̡CtŃS�B؞4&�(�p8�1�6o��:�E�s2��ûms�b��{F��,�`�Ԫ��C�D��P�Upo��O��|���,���Z��7Uh�[�'$�t��׼S�ت�������͊��ӷhۀ�����v8����wB��s�ʝW��D�П3�^�\"���qrho��j�#��>��]r�[�YZ޽�|1Ez��Bl��1�m"k]8M�}�έ���7G��H�ne`�\muF��3�q�)�{�(��4X,�J�$�����Ի�	�m��R�i�>՜��m�ed>����#m�1t�'�E3��K/LtF�.8�X2������mv.���[��B���q�L���c�^��ě�.�E����,�fE�=*���-mr���W3����X|_�hz�]���V:�Ι�3X"�K"���ݰ������Rq�_B�s��=e�ĸ�9{H�@;����Θ�=L3`�Sb©V��sk���Õ�x�����'N�P���Ӌ/���R����!w���{�}#�o�~��/ά�I�g;�Re�����my\8�ὸلviոs!�;2�J�99��n�ME�T��v��`c�;P�!8���'U��ɂ�g!�/�dm��GNU-^��ӣ%z11���1�yne�A]KUh�[�r��:L��bٕ��u�pdz�Lo�Ao�>�h���n������k6Yb�p�M{�ˮ�V5t��A���j�{��w3�YιB[�sԻ���2뫢��N�D�g��Sd6�9p�\]���Z[r�@����A�ƸT9�%��ʧ:��]�%�0�)�%`N>Sr歮[s]�9��U��]v5�����}�L�J���Ӽ�NSd�/��(�V�y�D�k�^'j�5�x���K^�+�Y`R�e{v�����f[fT��f<���N��JBR:�@l�t��GxoK8���U��D^^]*�sl�,g7|sϝwT��s%F�g��E�c��p&duT�;ջ�z�oW#r�V��\�XE�ʙ�27bw�#)����@ʗH��e��#�J���'[5wAn�u�|��/i��R2k#�����^s���"����:��:����;��u%I��q}}�1��񿭄d]�3��u\lUL.�uC��������rOz�A`3[2�1�kM%&����b;=]�.�U\,���A��ib��pO�/Y�=g����`o˃Tky{�Zd�TA�8�����w�����E�E��>X$^I��rȥ[��m����{`�.K��ś�P/՜kL��c\�!ڒ��ˮ��(�g��"���ΒDٌb�Mp2�3{�����7;���UX��a��R����0z%�ۦ�j/鋄�[���ib�S�����ڹ��+NPF��9mHr��!ԵǤ�i;�KM\���؊��Mc�Oe	���4�Dy���G��qO�-�����]Ҟ�V� �D uoF��_wݚ�5�p�+^���'\��;h�N!WE{���ܜ���E6�v��/�@=Y]E:�m�8f(L�B�,ף��
�q���#<�v�����c����Ww�͚p�C��DLP��T�ņ�2$&7���'у�o����)�8�*$i��^���k6���~�Q����UX�d@��n��v��eTC�z3ǳ�w��yt"I���F
��S1C��t2bKq�bJ�l�������*��d����@�RMS�~�޴5}ݰ��A��9L�/�|+_Ѿ�L_����EBа��,.��������L�)�����wI�Hi��a�q��vj/>ks��C��V���T�x;Dּ��U���Qǔ8�:�7����"�-�l��q�}�M�9SG̣���E�{,�F��&am��ӽ�c'��)Ÿ�lX��S)t�9d2,Hr6�P��v���5m�%���U+{,�f_,U��O�σp�Z���{�iy��WW�f�?��8��b�z����;\�!?]
�k�3�K�5�UH���<�Fȯb��٪�u�}kb��Y�^Guu�n:=V/f��Q@[L�u��9�V���XѼ��X����n��qS<d�]�.J�T�!�\�ahVS���-�� �4�褧��F��cz����BE�v���@>�d����H=F��WS����@1�kecN�p-ՋW!���
cȔb�?Xw�D^y���r-��<|#�xe//�@߳�vv���]�y3�O��e�ɅXx���BI3�`�n��j���ԕ�L�`�k��]��{_"9�!އ�\?J���M8�VTu�Vd_�:f*�:3��3�ʈ��p�}��l����ֺ0v��xk��{	�}��ܙ�aC��s�CȑB�3��T���oa�"a��`������$f�׫��V�3|gnxl�.9���ˑ`�j`ܘ�9˘v�CuM=�����9���
�z�R�|N�g���|lA��f`LuJ�.GH`��R�!Gte�+f�C�%N���|���
�AX������ٞ�H��^5/��u�3���VV�9p�["`g��.�:�~Ę��:�U�yF�&9eI���������3��h��deQ[�V�^�������O>�%��y���
����a����N�6N��E�6uc�1>�~.�͠'�j���n6����)����x�^���g�9��l���W�zV���-m;%�߅b�b�����&s�9v9e�Spܦ�� J�b웗Fb�9��m*Dw4w"��:ZaW�"�5�����[˯+���[�uቜ��K��(44��qͺ�W˚��l�by�v��f�NV��P�$X9�c�O��9�g#ݖ��6�F���~�%}H�d���r���9����>ړqW'� {V��e�P����O��ݛ~L:�KC�^'�b�q�"ʰ��������R�F��Tk��
ܚ���D��TvԼ��+�T(ad9�=1�-��jB<Ӭq�p��(���4�i^,�ڕ��ii����
�Cł��U P�T0 �r@�.�.zO	���2��L=Uu�s�S����\�Y>��V����aJ3�]Y�X<��\I%�GLtoNRB������-�2���ՃN�MΪV�d���sJv�^(�fM�C/tFx˄r:��upg��Y�����魭�"Kp�k5s6��9e���/ޙ���H�����W���7���Ԩ8�:������J��c�׬�1�`/�{�d8�T2 �Y��Q�=-������9^��ZO&��S�)���"�)E��j�鉞�
���)�=�.�em�^p�C�\�!2�.�v����'2xS���B>5�g��Ys2����s|9���5Сάx8���M��Z�=D�����׉#V:S�	�c��ͦ�owV�{�0q�A*����m��	��+�\�NK�N�!��n�0#���5�5qӳy��gMsL���c-�瓐�jVoru)�W_&�4�b�8Sl����.[j��:�yW<w���o{AcD7�ϛ��ic��pݏ�i/-ի�����/�XE�
U\���6��ږ��T�V��쑘��]ڭ�'��l�u�(���
���$7�s�+]Awގ�����"��N�������g&���j���ı��1C�YU���XZ�y8r�}�0r��Ph�48��!"�	#s���G�Zo*X5�,�y���l.{&���v�0>�=�1V�n&��y��Ve�n
�Ɂ��3�Q1dd�7<w�R���(��ޖ\[�"C��[�xv�f�[
�v�ߚ�\�:�'l��b�a�V�(zn�Z��4m��M���@j�q��0�������⋮��g��\����;�Nģ�Ψ��fz+X��'Ԅ�!3�xF;��@��^�U�Z&�͍�!,�ʗ�>�h�
hm)6^;|%�|kz���-���kF:��5Ow����\�r���BC����ȇ^(d�p�g��.��{1���^�{��n�}����с�o�U"Ǝ��������9����h�xW�W�����貆�mX�WMf�?H^�P����;Kx40�e.��#��Fs���'+j��C�ձ���A��p���9r�Ϧ��ֻx�AB��p3�V��պiV��h�7E���d󵳞����u�S�S�T�{A֮|0���A���PWJM�:l(yp���U�S�Z�[[dV�P��XȌ�7TzD0C"�$:�H�E�윣��<��p�J�W�.X<�u{Z�7N�9����0�t%=���S���*B�9��q��\-ϱ�S�i���';;��Z���]�H�[��������SxLP
L�,�:^�3�^�G���5�U]�k�.���EQ�riF�""'y�
�S��3�b���9��4Bs���Tk�6���y׊�si��5"fG�B�z�O�jJ*/;�P럭ࡅ�z3���f�Qu�W�����p��4��Ź�7&�6p�^��DM�遽s�e4b���#Fޡ=̾��5���k٨��e�\�ᴎ
Y9��({�U�VP8.qAR.�T��v��SÛ"&7�T�iܵ�}���x����͗�8˪�µ�F��:��xۣ�j�A�?j�o�f�����2�	f���T�c�.������,`�����YN�D�����n[�<�Z��#��H��{JuL\Z���9E*aL����0>���Xih��E]u����8J��#Dr���7�S�\X��r͘�����Px�s0�I��v��q8i�޳����� k"�z�^K'����2e�ŧ�7ft�D���X�B���/�~��z��+��:��F�M{��Q~t�΅.�aKA�e�ĩ����k�U[���(о�GVKF+!�p��s��Q�)�!N����ܸ�̦��w�Nck�\�&.�Ix`No������Ppu|����$�|�;'�����I�z�h;w���ڭ�R�R��.X\)-C�F��b����D���m�w>2��a7V��+�n�:(��*aq��ѫ�9�$t��1�b��R7���,PxZ���"&obq��pI�O}̠��n���!�f��cH�Y�1B!���]6�彇�2��uam]�w�v�c�w:h	r4Ѕ4�sUYQ֝@�U??πG���XK�����E��$p���:V�3�Y���b�B�Ξ��S|:BT������
���*���s�7�d�܅m��c;q=�[|�ţV8d�Y]�����W�S��X4<���1
���[�1j���9m�䏩]7�|r����r�/��ڵ�2���t��0S�9��b�ʲ�f����v�Iv�%y�7�B��fr��)��,�nL��w-1�i\1Zōh�%<��	@w��.��n��᭷L�}�}h���/E�{e�]�Iw()�5�	1�i
��Tv ,ң���}�M�W{ڲ�X�f�P<�Aܒ:
���Y��T��G8��d		p`DL�Rvu�*�{�(�W̰ypJ����������GHG�oe���g8d���/e��2��w��1ֱ���9��4��o%w\�I��Gj��ږs��H0�i��S���q�+���w2[t��k%���������#�����wu�q�
i��U;j�����P��Eg�N]�_7�8����J��t�x�u&��u�`��J�6/��ab8�3mK��Z.�gn4�W�̧���=q�T*.�z��Le�[ͅ��ׅ��7�P�]��� �R�:�+�9�jiv��d
!�U�.7
:k���k}��������c���pNLzN]�T-�*W]���K�nLO<���.v�H�vӪh�Q��6���˻Q�>�wnK�+���Tϭ�*S>�ɲ���yu���Yuo��[������B�k��L��H��4�;�Mza�ԍ����}�dWwq7�bObY�Є$W3���5�R�K���zT�#{ٚ��h��s�M��n͡w�Ǎ��}qZ���R<���1-�0w]�]�Qm҃C�M,�{]q���C�CU�>(�3R����0�����0�١�J_6�B��90�"
�K�VR��l0�� ���A�7�������o�B�F�:���N�B��Nɦ��PIM/�An`IR�F�rfKS��2�YR�M�	���c��Ff2�S��$�fT-`��-3�K��y�(;O6�n�*u��u�7��d��j�joh뮵\Mn�P���9w~�$��d��m�j�.���{k_S��ۚ�ѧFe*�ق�"q>���f��0��uI��9�n��<7���NH�(H�u=G*�-ͱn)7eNndD{)m��
c��v��5t���-���,�j�ZZ噸z��S��MS��10Uѕc8R햌��栵���C����i׹\o�n�X4��b���oe?��z���I:X�|�-#7,��)2%��(�01����Q���Ϟ�$�-A����Q��&>��r饔�s��.��1�
�;nM gGRCyY�T�=�������F��Yϻ��9ǧ�i�����b��B����J�\	�v�qf���yb���V�N�[���"r��G��?4��>��(�h���(n�X���ӳ��{g�&�=��[f���1&xP��0-��F��dP( �n�Þ��~HV���ah�)YU�Km�R�Z,�m�������Q4%(
EU
���,**�*��VҖ��ZZ�Xa5t�cV��.4��Q��\j��"���B��b2�j�E�5�6���`��J�����p�Ԣ"�-�ѫ[jVUc6�v�[!TQ�*��h�U"E��������TV�ADKJ���Df2���-�DQ��e,�V�J"֍h�lj�V���ո���,V	���ib���Am�[kAX��Z%�D�Z�V��Tr��UYkT�V��aV�mj6��Eb�A+k+F���*"���"��U)Z�U�M҈̲��t��E��֊�*#D�Z2�"�ҕ��TTQX��Z[mkTEZ؊"[TDd��(ֲR�Ar�UAUA��rʵ* ��U��AAM�Q*�U�jb��PV��a[lJ�D�[jFm�W,U�4���v��R����ɢ���tj��(���c:��Ur*O�H+�pb���Lkd\�vݺ�l�gqZNk��o�j;��v7,~~�\�+���<^�^)�~up�⪴�>񿅅~�^EP���MxT�q�ޞ�]��\���G����3�I��\�^hmqx�͛�c��29��j���oXBw)^l�H/��"���WV����T��kD߼H�0�2k2ʀ�U*�YS��%�3����w����t�nk�;9�{���d9b%�z�y7�y��W�z�Q����5�R���d�R1a\�^��`���-��SS������	f�X��`eJ�ˌ�lѡlOp��V�."�J�J��d'Q�0����r7�q�Vݖ��Y�J�u��T�HJ�r��XT��xLr�c�l��<ݍ���2�:�:����)_Tg9F(C�S'���T0�G�|2����2'n�z|�M��XC�����>��o:4*���.�.	g@,FʤI��pTH�#V�ظ˦��u�vv<�:�*z�ߵK:�s�D�r*"�������,�1��a�<ԏ�+}J�p��E�V��tZ�X�%,�U,݉�
X��Y�s5�[%�������ț��ɡ<p���%�W�R��`5ʌ����[\�*��&���p��"�T�*��:��Z�_�t����WTaܜ���j0�7]]�:7��	�9�
�k���Z�e�B����E����< ަnq�6zS��#
�+�¯`e����L:'�G���nU%���u�_�J����`׹V�rM�k�/M�v6����`��<J����.X$�k���V:z�ۋ���y�7��ܕ����X���;�Z����3�M~hWDxJ�����L<25F��ug����FU�7r��k5]�?�3��G�'���>nM셂g�f�)j��2��n$E��k4�U5�վ��L�1����4�,�'Xl4g�	e�*r��xL�t!�~�.�.����g���{y�3���E�6h�b����	��w6kM_N2w��ZTV��uCu���ym���V�JF��S67&��6C�������w� � �h5�x/
p������-���7���E�UiӘ��K5�,�cg$׻g��hPY/6D�1�I� .�鴕������e�m�z�ɕ�}��+����DY���v��b��������\��4�h{=�vB�6Ƨ�:/���k�l>��^�)	�(*Dd�t�ӽ!t]W����*7ko���9�fvY�8�vlM�NE���t�qǻ�s����ۉ�HV�Q���s�h�HYSK��<6+8��uJ!h��u���v���m�SǙ�w^����^�����\U�;�#�Jp���ł�PR�gM�zkA�0R��{n=]�����P\�<̖* �:�z�Pe�t��6�t��6�p���^|2�����L�i
�YK���y����8О�@9��qǭ�BC�9�ۺ�`�ȉ|:�s�ª��-��[:�����V��%E��Z\0?�7�"ƕu#��q�3��X���c��0Z6�f�l�V��=b{w8�Y�P�[������?*�Tpl�����gY��>[J!�p>���r-����k�C"�����0(:]{�*�ӆk��b����Z�s}��Ӽ�/f^S{8���'Zd]:F(9C�hV����>컣��K|���e7��Bؾ��{}��*e�d��x�|����|�o�a;C�gSxGC6��;��������Wy�s�jl'X6g�*��FY�پά����xyY�OEOQ�Cn���\�t����\kI�	���;�⻽6�X­� C���a�ulRQ�U���9�7��Ym^�6;��回X*���6ց��j��%�y�R�>��M��oʶ
]o���>#I�����J�IM�,���Y<Eom֖����ʞY~�M7V��^]���B��=l��]'�>������8t�]�G�w��;������a��fKpz����?��إ��8.��yN��6J��6W)���M����U7�w���y+��L��U�[�͚<�2�0��#�9�Ө5�F����>�^�O�,Z���Q
�CѴG�����f��BO�3�XG�]�u�3�@�}ԋ����He�{Մ�Hd�%��E/����U��V��Y�U�i�����7`p�����Q���]�f�W;��:h<U�Wg#M�&�#�L^j��y��I�Ng5q4���-V��x��Q�w"�V��|iQ��Q��8g��ͅc0%W��;ԩm�U��W�\09���.'�*���*���u��=���W��1[{s��}��'��#�<���\,�����Joχ�+'.���.F�F���F�TA:�1���L5��5z������vLX�슽��b\ۆq���k�]���m�Qx�����"+ؕ3�-��7�� ��A#3�b�@���� ������<�:���Gisu�����3*�v2G�¹��n�+w:�:��+s��̫��>�6�:"+Ljf�pJ՟,�k���������t9T�h��{z�j�G|Ӿ������Z�VՂ�R����y������ڍ��C�N�+�&��~��]��r祟g�M8ˮ��-�Vd8f4C$�6��������v�=��5��"8�E�Zg�2^�̧C�*T�):��y;ԩ�/��;Ww;b���jeu�6X:
.��q�+Ҧ�(��l��̂[��k�0���"�ޭ��]a߹rh���v�fm�"(Ed><t�J�FD��p�J,%��%���}e��U���r�٩AU� W��
 ^�QU��+��-^H��ʓ4���Lp�(���i<�u:��USo�w�����a���u#$3QёfhtLO�'�&�u<��!�z����ej��K1��E���{�N������dTc�/���-�/��D��ň'��A��_B��X��H+�kg���O>G����Ǘ�۳�-��{6BL��c���6�|�{�LӐ��\�s���<�1���17����!�V�S������_E^�\�qeVN5ܪ��oT��w�o9�{*M�SOj_�A�n2�[���{nY[���ޑe_���&����gm��t�e�?k��)u���t�)���٫�{^W���7�Y:e�w���ݛ�>�R_1~X(�E�V�-� ���s͛�J-���[]1�aZ��%�2����KDܠfl�/��ġn���s�f�������V�6�u�)������G���6�..ͦl�Z�ܾ퐞�X�I)��p�!+�;�tj�/���#�<��T��R$"�!��G!s�`sW��+<�+Ů��62����ihWN���4���n����*څ�Q��g�P�W�U��ˉ�Up�G���eg�ur���96� ���t^�eX�D�B{׊5ˮ2�FhF�%�b8�<Im͖8�˾�J�Ǥmm~��Sz�=Y��^p&"[����(�`��20�c��ͮC�	՛�f��X�P:xY�h�^��:G!�����yF8�P���.�B� ek�m3�{x.!����F!]~�<p���'��
x��>���ly��O�e;�[��e�����7	օq�Ӥ@?	�&BB�sbz!�2�Fĸ����{� �R�!�v��<n�r�v͘��g�6�g	4K3D�|&�Ĵ�>U��O
5��ڏo״}����v���ł�Nl��qZj.C�$<RZ2��n��ڮ�jn��w��+�PvX�y�/r�q����b��)�DW���:�8��^su֗�N��²O��au�3RJ&˥��!�g��z�kG�4ϼdq ���:����o����vЋP�.�< S��lk�x��Xxj�b�w!��bw]���N|��2U��*=�����5�0�9f�t�~������m�� ?_ �h|=C�b��F�v"�^E=�Ӧ�b�62��l����]ۀ߶>��J��c��|�I��z�V���v-�i���|����GseY��_�S�_��c��>T�M`�P�m=Q9�?��EoJ��~�;�Wδ��d�4u*��6�u
�T���x�D̃�9'��3y�Z�>�\=:>���m���y����C�'EƑb0Lq)��!�O^T��ou��<��.v�F��v�"�J���P�ĩ��c�D\�(�۩z��K���o�Mq��!��Тt���85	��m����2bV�!���'��4Uo
�_���=
Q�,�UHߦ(������O��S�׌�5�qO��;�J�K_!����/ՕD��Н+�/?$�+��=PWJK!�)j����q�nu�|-��Z��fRج�F���p�H�+���udF63�_N�T@��Y�N9Ew��=�uj�^U��V�q�=���F��٢zxן�����i��2��F�u����w>�QW���V-���-u��}��Ψ��7�`���}Yte=yJ��M�9a�q�8���l�K�Im��;`}i�|��A�xg(.Q�:Y��C��:GA�l�~#8�cyXU���/����`4���gN[&�6��6����w6z�U����N)#i�g:��q�hR�b��5~��w�\��r�+�x��a���
"���][�`�	���1!qN��p�PT�x��Wt�M���oxbQB�Tf#�Q��t�����az�($G�1B���v'�8�pJ�!�9%�*����6/SM�-P��Xܚ.�p�ũ%��u�sRLof�������u-0s�3�Q�$'�rX�/����u%=���1�3c���5��^Q.ȼˉ�6�A_eG�F�m:m=�Ȭ�j��͈)�껍Q�z�'�����u=ZO��w	E嶂���0�,��w�ڐΚ{ՄX[��]�]�Nn��iQ�=�͵V�ŝx�n.Gn;���<�Pي#Ttv]�fVOl��-��{~Xx�Aܢ�FǴ��vm��}�I��{euY�,�-	�Bܒ:�R������J��8�R�ߪ�Z;�~���5����P��@Fc��yI  \eN���� � �_��8/zkc6���=��<ITUID�fre�Q"�ѹ9��ǁ$72e[F�8�,Z�Վ�μ���]��Ei�M�윥r�3�ѽ�S��t��l�ǃ��l�殓�^F��W�ܦ�'��St�%��.�<���4�	�*����9�ǒ.�|c�]5�*�58q��[4�L�E��F�z���KV<�	����X�AJ�I0-��1N��ۧ����u�Բ<�d���2ƿV�x}*� �à"^�#~���Qo3.��Fq5��0�W����մ9^DV.�r�=p�Y���
41	$O�z�e_�� ����Q^�T͍�U �ٳ������y?�[�&3T�8�t�W��Yf<n���&��w��s�u��>���D\�Z:*<
��]�V�Ј�P�Nf�jD���읗����`�hꔗ
�;*7��t��,XЪx��^A-��x�Jv��4r�����X���0 k`Tcz\�!2�B{�Պa��d�\J�|dd{>�0�Op��+77ǹ��� �Ut��	�_

N�V���+@ea��ۡ ��Ň�8j^&���~La���y~��w��&��r!����D�<�#\^	�x����ן������OmH١瞳�/��kM����_e�bg@8}w��\/(
�V��v2כ�2;�tC[����� 8;�i
<�8e��J罏�T6e��V���oV;5�,uA�d�ɺ�5wV����#̶̑>�P>������R��KxlJ����#br��%CJ��vJ���r���R���/��ś>��i0��$ѱ/�|�Oh�·0���#��C6BL�X�u:l�[ы���3���C�Y����G�X&��9YU��[�6ჹ��7��#T�]�j�Uհ����ܷP��3�_��W]�8k<~Z]y��῞&&�ѕS�ç�Yq�"ʩ�"���jʍW��w�,Q*�1;���9J��nԻ
Gr�C"sq^�'Mz�\B5BY�+�_<x�^c�TXg��9�/'�l9��Q��kʹ����*�~>�{fo��o)I��+�s$з�;��qƸE-tO���^(���xU#5��f�`�1���G`m�9OS��Z��,�r��}�k50=�>���S����h�j)�)S��>�ʽ�y��E^����1k�s�e|��JZr�\��ޯ_���K�&�� ۄ���|�w�	���b򃈮^�hc�t뎘q���FEi�*��͛�F �C��Nnk܉2j�d��h�|�a�R��Lo�7���-�֨�N�ڝ5_E]4|O��Ui6M���d\�'�q�d�GLgFK��8J�U��=�U%݄3Fi97p e��Z&iA�T���|�<��ݹn�"R�R��L
��:Q�PT�6 u�yEm�k�Vw:���U���9�M�A�����a�mU��iݿ��־0��5b���ǳ�媵Vĉ^��jb�i��skd��{�qPlNw��+��ܷACwM�f\����te1�ج���ޅ��c6�-�ܚwW\��*�̔ ��9P;���`�1�u����P��/m�"�'G5��qY����&�/��N�VPL^��4l-E��/��睬��f@�f#�����������.I}'L�����f�&����bM�����$�ɔJ���K��чT�]I�v�/U$ *��b�-�HG���Fvv�Ә}��su�$�H㗝����i"�Z���{���teN�k�ݺ�P��X㥳zp�٫#��]n���,�HT�]����[��l�ͣV�Xe��,yV�Q=��Я@=R)᭜cFf�md� rNIP&t�
t;��e�-k��[��ۍ��dgL�����A�b�f��n��`�e��<ë�o��fs����K�^��%�����1U�ىoHݍ+9�#��.��2���Y�\o%i��P�������`}A���1�[n�g{N�URկ1��nueX��M��ۘH�~�6�4əqhn��.m�:qN��]�d�Y��L9x����Y$˽{k%d�D�%�19X�G.f+�ݖ�rX�۬������s2s�r!��@8�-�{��43g�����Hĭ������g��
`�OO�����¸�.��ec����&73�S��,��g9\�c����ef7�i}����+*s�q'N��9"�G�q�n��B����j�',kzvڻG���1��V�	/��
5lq�Λ\2pK��(�}�(�{!�%ڧ�[��;�;E>��;���aUf⫑wa�WS5�/���˽4�\:L���T{���.Ѧ�_Y��ᗻJ �m�w;�Vx��L�As���4i=7J�a=�Ʀ�}u�h��<�Z�늞�����8 tL���h�t�G�a��͑SÃ�����Q{Jۧhk�(,�p���մI��s�S9�,rӔ����t�
�r,Q�gm\L�Y�4y����i`Q��z^P�Aw1r��nШ��6�3KD��\���Yq]jtU5)��5��R����:��<ҟ4sJ�\om��^�}�����\噋o�\i�����Y���;}��. ,���1�v����b*�,u��n�	��yd�qeǖ�Xz�jBiw^�G\��}��vaW�.�r��[N��?eY[b���ͺ�|||}��Ð�Tj(X�}j
�EAEDX�Rc,X�J�)R�ecl�%J��d[m�X�DUѶ��(��
��#R�"�mEPKeb�Z�Z�ՌQTU��ZՂʔb�mF�DTQZւ(�"*,J��V ��Z���k�Qb(��Ŋ�(*��UX�"(�JV���*��e�e��EPTb���e�b%���ij1TH�ZTV��6�!�Qc��F��A�F"+b��Abn�QAU�[��I��ZѴ(�+mQEDcR�DEF�����i����e�E`�ETU��1Kj�h�J�ZF,EF"��U���q���6��-b��h���%UDB�f҂�UQrьD��խ��A��)hEX�X���+V�IVm1��Em�Q�EQ�,����DEE�Kh "(����we���Z��"*��($Qb���V#���m���j�a�ECP}�I(_Ie�{�Fl��ܗz���ۨ��펩N�f՜��@��e��k瘺�[ke�:�kF8M����Q��:���ct�X΄.�G�3b>�5PD^Py�4��J!���g��XsPв��"�3�m缺��V�Fۜ1(�*Y�o��M*�]I���1W]%�|���Gʝvv��i�|i�����lu�+8�"�T<X(�'Xm�8f(KpH��`�Q�u۫��5���&4��~�4�Uڠ́�%
��\&"��dEs�k].�;8�Jt�Τ����$�S�\�dm��h[t��r��{CO���V*�w��j����8��\���e����w�߸`�U7ƷU�ԻX���|=N�h���N�6�jW�4�[���KQ
.o80��M��ʐ�[�P{ا�@���n�߲��͆Ym��^8�w���
��7���Ү4��wb��1�,�%�ؓbbL�B{����s��į+1�0���[��/��A�qw�ZF�	6��9݊v$n��M��]1�37
I-�S˹UV�aj�;�պ�Δq㠋.T��dnD�iZ3a��
�[ᵽ{HKog5KVF#�cn3��ͥ�l�|V���8k�\���~�w�;�|�H�#���e���6)�
:-�}E����`�hXUϙe�˔TŹ�:gGs�E�vH�y��\�vXKR���&��ܮ�ĳ�糲Ԗ����I3[�m��%�x4`�}�&sޢo�9S�2�И�X�eXK�#�K�B�5�^��{�C^s����+i��f���Qx��ъØ��ŅBv���ᖗ�S��)4t�ka�?l/TۿX�|.�1��Y�M��YԦ�xlP��&mzGW�B�]#�t:�����q:͉��o��V$�fT6�q��bgry9yv��C��#������D`�:n�.Y�-�a^��赜�ݧ�8��V�J�<��V��qG�Ru�EҤb��$:�0(�а����<{��WL��!z����<v���n��xFSp��Q��s�eK�\�<)gG+���X��[���άO%��j���hw��<n��ig���U�C��������[@mż�Of{�-��A�+�&+gƮt֏#2!�r�<�������[�2s"(8ԓӸ�D�>��ݸƀk��^��:U������[�Q�^�g/���|���������{#b��{�ԯr�J{�w���x|"?�Τ(�"b��w{Gt��~dY���FN��?"�V���:/ ��F�>�-��Qeuv]���&"��F��Zb�;�*�C�;Hª��q���aY��:���w�wE}��}�=]��@	��۝�X��M���+K[�����C�K|��+��+�ZŜ�./���v�����q�5ե��uoha�~kkr+ i؍��vo;��D-E+>A�5�}���Z��ݞ!�`��8l�q`+�-@g��XE��݊jt�w����N���E:`�*��wpŝ���^��u���E�f=�:4��̈́�<G|Q�!�W�A�\GkaVTk�K{�K	f��,f�w��rc'�p��h3�
ܣ�
���Q\�2��>��*����If1[yU�_�B��e�
݋�VtD#�m�.��ұT��|]�bZ�9�:��y*�F�F8eڹ��Q��
"\D��%�[3�ON�ꑇ�7�Nݭ���Z��v��!���w��t1��#f3գ�Nw�1l(q��"�l�^�%E���,?_.�Dn��-�r�Y�,KB��s���y�K7QM�*�`9 �6����h�W�:7Y�i�2�'n�)����^������O{��nӫ2,
t�v����q���֊��$����i.�=tEύh�]T�u�׳�2���RȠ�U�����92�ʤ`��F�gv�����l)�d�m7a�c�����dr��ښ�ՙlh�oNWI�ҎwG�y}�����&"�6-ch��!R!��ӍM�]grmh�g�S8ŋ���=�t]�Np�i�
;*�w|2D&[���ں���ܔ�;���<��W���C�ׄ�8<�7��~�71Sx�w;qc �f��lc�8��r�m�����{Y���X.���T��UB�|��]M����j�р���v� �|k	޲�r-������QBv ^��^ T�H�ћ��r"}�{�&�Y�1ٳt����ܺ�v�K]*�ځ�l���(WI*|;i�4�v"�ȳ5����<�"�Ck���4��nn}��|�r~�ݙY#>T>"��,��]���b��D�b	�DL����k�[VwuzG��+��+�C�G�K8w�LP��!B�Bf�qE��O����V&����zZ{����Yt�/��z-�xu<�?���:����� ~��s@U۔{�9O���!��9��g:�j�������5��7O-��W��?�xx�)z56�K��Y��u���೯�w�A-_��??:�\h��He�B�R���+��"��.،�/�vQ�R͛NQvu�˄�j�(�z,�yU(t��6���Y$��n���%Y��B�+{��{����Yǌ��dY�� �s\F�Al58�*��y�P���6�.�פ9bu�K���9��F�d=SJ�S8�n�R�G;�<�V���+���"�bӰ^�͚�aT)��!�'h���K�܂t)v�s�f�[v�F:���E�q���5Q>I�p�Ιvz����E�.��Nl
���g%�az ��)Y&���ӕ�ϋ�={�xH�b,7=q=�5C]�[��]&wKQw�jg����eup;"����	��;P�
�ٌ����6�JG��tũf)��o1VnE�%��Y�}!DK~�q��9U��K��P5�<
�O�z�B�l�3:z�QW��17O��q_�C5�/ԥ� ץH2Bh+
�le������FmMq�.�>��oWk;:�=��j�b�1#��@�g��$׃�D�!��Hy2�g���d��1-7�m�!0�/bp�rȰDtQ19�<P(����ќ3,�%NT�x�*�B�-1ֻQs�h,ÌL���Rʚ׎�ʠ���(t��jbd�s�3�cL��{���e��\�8�W1 G��A�YV�zR[g%S���t��b(diP���c�����'6z�Md�mkA�K�x�����=��Ui�C1V�ʖ�������F"�����	|ѱ��^���Ls��8�
��Sw�$��cwq�i���n�e��K�w�x3C2$nڂT�Zx1��]m2��Um9+G)�$�����8��d��s�j�iK�ׁ&�T��R+�5�G]ԩ�>{°�V-Ո�R6���ƕڞL!N��~������j���ѷ�B�傢2�Z+��=����{��&���z'���X^��meU��_�B.)ݲ(s�g�y�,��׺gy`7�hK4׶JBU#l����1��;�KP����E;U��`oK���,�uH���4�i_�4�*��y95�6�2���e��qZ"��\$i�y�^�J"�U3�}!d:��pt�퉴ݣ;n5�m�DeU���i�]��T�U���'���*��=2��̑���5���85���3vˬ��E⚩��oc[z���)�10���@�R�2Κ(�6h�[��#ƅu�$\������;��ڪ�'X��E��:����z"�?HTؤyK�v#!Κ����!�r�G�,M{$^����hy|9x{�U���C� ,x��bZ���s�份\��^�}�����`r��46_���B��;�����ų*�ɅM��_�!\��i�#Q������wtȭ!�ߨk�N�p��*�ئםdW�m7��U��)�)S1�f4Ȯ�n�Q�,k&�G���j��07��Ϭf,!�P�I��{qLˋ���p�!Z���������ʾ��e�]��0��Q���%<(lX�8+TY:���{DU���MS�øoF��@�ęx�J��3������kE����Q���m��|ޅ̾Z�Ö_��x�##�`7�PVy�6�}B���Y�Y�@[�B�a�v�Ҩ�Cn��E̷�e�Q�֙�S�	B��/g&���lc�r��M�Z��_o2��q�h�=�},�g�_x�����k�3E=��~��̶�� 6��y�4�Fs*l4�L��XhNl�sFZ�r}t5nOz��.M���B�Z���K,XS��]N��:m��Ȭj��V��[ח:��ٛY��ֆ�r{��nN��a�-���c��6Qq~Wx]�v׈���u���5}�l�ߔ��ۭ�4D��~��6!~ǜC��[R��@��T�,5B�
�l�w��ocK��8�=�w�7+u8=�վ�c.�G[Ԧ.L\K�SԴ9�m��P��Q��n:��U���r��[Z_���S��dK��e��KbçVt`�GM[��Q QF]�Z�EX�{j��P�>��������+OO�V��9.%��2:��\D.�a�n�;��F��r��Ay��e�I�;k�Cq�=�a�U�B�;�t{������^�.���_L��Ztՙ�>���\�q�Tμ�M����:SC�����v��f��l��N�AOO9&垺�XcΨ�s�P���� �sn::G�@�c�ujg���.܏[��AQ��1k��ϴ��@v�7��o�1�M�������>��p<_z��Y��ٝ,�W��-��&���Ds%N���bM�J
��q1��^�GX2��rP�^l��\f��yT�*��Ī����2����0l���kC\�X>*C���p�޺#xDn��F�d�V�ޜ�S����f� f���y��!nnFjҕ�"�S0k�X�d 0�mH�G�F�Y^ <�^-�Թ����01y��87M�b�i�:��>�/"��~����뤴[���է���>>_gb�1��.��ͪ��{"K�U$t�
�
�I�1�噯*ذ=,����Fv<-�5U��Z��~�g&�`�0V��p�p�B�I/�X2Qf�Q"̾�1>�%�V�����ޒ�oT�Ɔ+8��͙Α�22�8E�`�HvӸ�ak��ٳ{Coՙ�.��K�L�I�&&�Xc�I^��B=�ەIo�٥����� p�L�+���S���ܢ���w�)��v�#��;T�WV�t��~|K��#:zc��a	w|B��!��/:��l��]��I4�~t����m�͡�;r�5��[��=�����.�.3N�G
����W),�!Y��g�B0���@J=�ce�b���$��<�zKf�i�!�X�4{���bf��&8	З(UeT����CO�d����:ms���,�R��
�MZg�}Hm6:F�F�ė�w����lu�BǶ9���ݗArr�;F���d�y�ϙ�[��-�ׇo��I[�ɺ{\���EA�#�n��yfw%�V>Q�K�pb;'ղ�^�j�*�r�,l��7`D���%�Ufb�N�F�tRb�h�lwa��k���[鮷m_P�"�;�/�Xʣ{6���FX��6����s����Qջ�N��m�fs�.7wO9�γZ��?n�d�)���g��dT��b!d�P+N'��Ё4V�S�X��]}�qzS�T�&��O R��}�>}V=�趺3�=JZJ�G
/]�j��w"X�V�3�L������Ӹ:�ĈBU4/]{�ñ��E�6�b�Gc;N�9l
�W�9�f�pN�H�]:��m�Դ��\�'Ky���u���:����t1j+�t�ݙҶ�6��dӒ�
�y��g�����72#����Q�
3���g5 ˺I�ѻ�N������:�S�[{���N14��t�]b�ɀ3y���Y�/'�;�'��F��l�K{JdK���Q���N��-�(h��jb'�<*ևs3ʜ����(�6��vynC�xf����WN_N]!`Sbx(���6/w�`�AXS����W����Eo�6OG=�O:�f�M�˞O?d^e��õ��uTמ<�	n��kNW��mf�,Y��M=n��o�zM7۩y�o͑��Vp��hߦ�����{{����r���nm�9hUn��f�٬��~�5�:����iW*�N���]o^��v�=�.+'��	j�W��&�Z�q���"�=^Č�N݅�;�btn����q�G6�͍��T�����NWK�#�j�\zq����c���ӫU���ie��^j\�BlJ����d��٣��3��R��ng�}�B��`IO��$ I?�H@��	!I�$�	'��$ I?�B��`IO�H@��B�� IO�H@�XB��$�	%�$ I<�IO�H@�hB����$��	!I��IO�H@�{H@���
�2���/> 4������9�>�V�Ǽ}T��*P��R�J
T��PJR�QQ*��UEIJR� !T�BJJ�JDJ�RR%%)UJUAPA�j�U
�)$�P��B�6�JJJ�H�� (P�UR*)TQAP� BT�֑UP��f�^�RIR%TB�J�QH�QBIEADUBU*����U�PJ�U$Q*�UUT("��!�mQT*(�  h�ֶV��� l�ƭhU"�LRBR�0�h4����J�_n��QD��Y�ҡAVʘiR��ڋ��D���RJ�J ���<  �@f���dU+l�j��͡��X,�U��H6�֕	��$%U�����)fKP) 5�KaEU	��+Mh��A�B�(T�*QDB�.�� v �B� h���@ �C@�w
  hP
�w
(P�С��q�     C�'p
  448��
 Ӷ��j��,4Х��d��Z`���T��P)\  �P�kjTX��m�4���mMT@�W��5+��B�U4i��B�h�
5�,���I�U��j�m[P�֚Ԡ��Z
*��$R�x  �@�K0!U���AKa�Ui�m�VK�km�2��Gl�S��kCR���kT�h�a@f��Z�F�,�QR�$*T!(*J�^   p�mmV�j��ڑjUR�[U�e��X`f�El��T����ű��QM�5@5aKR�f����6�U��JH�$��
�*)$�   l�IR�5iK*S[l�[U�T�ʕ��QU6++*kl����[@��XcR�6��m
[�Jd&����T�BJR�	Q*	(\   9 :Y`(R�h�%�mk@�LkJ�4����B��6
�M�(�`h*с��[R����}�EQBB�<   L�) mK 
j�P����ִ� ��h�Y�����@��!��e��(�V���J%@IP�H"����  ��h4��`��h��+�b��`-�� 6��(hUj�̂�5JVh��%R�i�ʒ�i�h�B)�IJ�h  UO�5T4 d ���R�   S�G�*4<�dh I��3*��@`)���8��w�����d,�{Ci���J[���m����Z����@�$��9������$�B		��$ I?���$��$�	#!����}�?�U��'C�Ӕ��D��®�d.$(�3p�"�шE.���Xj�˨6��5�2���z)"��Ĉ2�D�"��;���1Zb�U���(&T��
��k�g",U����Vj"��ۡ{��(#̴Kc$c�"X�-��uښ����]�7�Q��1�p���Ul�zV�0s��;x���)���7��9m�D�C4�#c,�V3n��j��A"�`���&�0z�K���FkQ��9�8���v�HD��[��q�-��
�m���-ydⳮ��צ�JKsn���T��
��.70Ls������a2j8�M!�A�7�ș9wD�-���	�W�ن@���R��a��l�@��KH�ҕ����o��%���$산mņ�,`���E�4m�N载yM���j�	GE_J;n�V1k��ػx��Q��8d;�Ѐ�è0껕�"�"�x��&-iz��j����5b{cuN�X����9��T�Q���J���k�۽ӺU����.���P�I	�0+*Xf|�8e�����{[��̂�cu��oA����)�4Nn���8ʏVZe̓F�5(�Q�V˅]$��y�w�A�5(*���ݷF�VXN]�U+ܙ}1= h�jU�mY� )�X�y��3���ql6�LJ%/r�HF����QҬ�]9Z���U�n�4b�����W ��*&��|�<yf�ٻët]'�ƑL�����+t�A=�b�ӸǙYMV Dt�$^^,Ǥ
J�"�[R�5p��:ǚL�V#Eg�Jc0�B�F\�c���%��0Q܆���*�3A�+J��V��^e:��KfK[��|�@��@5鰐ܨc[��@MIZ�Џ���ZMJAt�(NAz �;�a|I �D9���8�����dL�g��7[u�5C�1&�aZ��Ŕ&[ڙ��4�Y���e�1�"����e����I�)WZ�*��&f2�fp5J�I��4��r�}��j[b�on�',�ƥJ����%���.�m�9k[KA�m�Y�+*@/,CZ�1<���$�3
�!V��)��U��UjA"�/H!�[,S�J��4Xw��vTi#اTȤ�ŗmk[��Z����ݸ���޴� +an�6Fށ�����;��;��6�"6�F����m<6���(|��1DF�
+P��YU� ��{�;c/vVR���w>����6��	m�V�7` �V�6'A6j�(
@i4��%AͼF04����M�f�ܫ1���X�Hd�Ć�0�T���h���$�R�ݼ�EM�K�U�*	<{YM�e�w�
��4�h*'�)n�-��Ø�6U˽5zmJR��h�HnԻ	J�	����U�ȆϠ�4
��t7(��0�;̇b���!-BLPHb�&��z�3m@�6��0�d�z3f��E�	e�F5T�b��#�ȷ-��lf�Y�ل;ܥ�Mf�]�� d95D��٭B���խ��tٍ"����<��L���'R�X)f�Iaf�f0�P�I*�ٹ1�M4�m����0i��j��r�Ru@}����ڠ�fam��lq(Z̙�6�ݹ���'n��M����t���u�H�K�07.�ę9t�ݻ{��u�\9aB��2�䵊Gq�2�.�!bV3w��ofmc�D��1S]��Cai��D�UjJl��۵p�("1���Mɬ��k��3]�WwSh�.��m+ɖ�!ZT�X���4%��5�^$�\��Y��7Z��f��wLQ��iyl=
�f:մM�HIs������ע���R�|�����SI�.��7y��F́:�[ԅ�݂�X=�\�p]���V�;��i����+ 7�UX��Q�m'q�6#�ʺI,7M޴�{vM��(d�V SS �a)@��o�N��n�Bd�1�34��mk�PLdf���-�&V㿍�]�j�%2ѱ��[0e�ʜz��[gD�
�<Pi�����c"��r����	��`���WY�n�֪���M������C���@~��O+F.��itJ�صZ���L��B�{�K��:ƫFV�L��L�%7t�l׭do/H��-PtC��lf)Z�w2�h�JP�Q!+�q���[`����D��GK.ƹ�����7�@�qk"�W����~F�Jz���b�@��4�h����ެ׈�+u�U�1�����ɡCXȫn�**��i�1�x��SH�ͫܩ�^dor������`�^]�%e2%:�$$��YZ��k�ǲ�T9F�)�u�⤍ӻJT�(��=ykQw���_ʰ���^���Ӂ�e�P�a�U.����(7L[�	-XgL#��S�ٌ!�����{oU�t����2Am�
Ŵ�Y��!�̭�5�4��l��7N
�Ŗ��	��J��,�)\,�ހ�#�;[��+�Uw���b*��SI��	��Q�C^cT��ۼa2S�	K���8�Y��d�"�Q���'�,�dʕ�Txc*���&�V�d�	R,V¯d{t�U�+�Ó2�\̟#Վ���L�sl�1կ��V"7��.�ifD�e
�ӟc��Q�	bQ��R�kb�ǩV��[��9���*5��hX
n�$���(���)�V-�HM��3j�in�wIwRyvU�dd��I"��̼�ʉ]єaEz� ��ҕ�q�+@��--<x�S�/2�q��MЙ�p�r���+\(�a]����FE��*�.��L��	v���:ʚ٩�ed�u#oV�V�)�Px*nXr�0/�"p૘�Ў�8�(p뺿�6����.-Ԇ��0���^��-c���J|�VhT)��&۱ut4y����[�߬^l��!Yi�ݕ��?1qaNap̬��hZ��e�IP�I;{ .R��f]mѭ:�7!�U��/5ly�OV��11j�Y܈؎�P�C,|0�`�ed���7j=ooa80���j�`W� ¢*����rl�Y!�q��Q2����0�hL���eR�����U�od6��c��7�U�H�6�^��h'(T��Lɇtޒ�[�l��`n�Ô[4�5-��&��IK͒i�1��\n�7w�VE��E��I����E*�1n)�)b�r�1P�k�E��e%�K��J�-;	C��D`×YPᴃq�M[N���-Vc�H@�  ��7%f���	8����TY':����0��0^e�WO.m�*^�SUڊ�=�4L�lQ{�.P�D<P<��=rE6�yY�n�=B�e��k2ҡX)�;��TR���A\+�V��؉W�4H�d4��`2� J���ac���ޫh��5VX���܌m@�TaM�y&��(:�ܠ^��Z)�^��k1nT�X�Y�BْڏM"���ȥ�#R�@�v:+u��V��u[6I;R��&�<X�J,�[���.ıZ&��/dx�����{+a[�ʆ��rŊNƅ����C^7o%�J�C9M����b��A�Bmi=F�t�<�4�'Yh�ɢ���{yWZK��"�����z��A���11�j֙R<��鏉�;G�][���i�E��[VsN�	ܣKK
�Y���D�AM��P�7�(� l�!*��m�-�׳i��֝� �&j�	F]'EJ�5Q�����%��R�V�V�NK����jL���Цε�f��0�Y���һ�����L0^�۵(e�{Z5�D��^��[vZs���r����I����>/m�#Ɋ*	JLڢQ�<��F]�MƩ4&c��7CZ͸�JT��aDU��)aM�D�D�F\�oD�������B.��.4)cr\%�E����[`��-���!��׻o^�a�ZM�6����cf�[�+c5z�Q fNg�;�ic�J�e�EC�YLZ��@dA:�]�6q:H5���ej��f�i���n;k,]�ܧe,�B���jdd��^Zzc�(0I��L���#SQ��b��t/>��=$Y�2�ZKb�nkO6Y�����&n�ݗ���l:w�;2<�b�8M��K&���r\��0l9t[*HV�bX�����;{�J� �1�kNQ�ܫk7K���BP=ګ)r��9SvV�al0R而Y�C�$�f^���v]ф���㴌��t�(���)Ŵ^\�u��im�Y��Z��M@0����0Lw[�E�,��Rތñ$/f�Yt��[��b33M�����TiVR��%s57Yi��P�9-���:-*��xB�h'[m�F<���4��ne;�Y'Dn�]	X�@�J��س+J�Rڎ�:�+74]����ʻ��)��
�X��j��K��śf��E	w>�n�!��R��=2�{����0c)q�֕":J�k";�!C2CC� o)��JW�n�M�wdu��hTo6G&�"hX���(���J�Y.��Y�7r3��Z.�� �1�Z�ܼךN �,��Y��,�SQ�T���G4-�r�x�1*�rk�MܔF�h0�L�sw��RZ(z�룗B����1FHLF����I!z
�	{h�T�#�yFM�z�mȪ޽��6v�j�o���Z�&�5H�J@��1Oql��֬Ɗņ	�C�KN� LE���dw`�
�'�S���dwJ��.�v6X��eK���D�+z��M�LN�)ZD�T���(V;��w �j-�wTe�i�ot]n���j���`͙I)�3Sd���͸���U�k�Ww����J�5q9�ܧ*2F#pjv�A����U��H�B*�	u&4�b3.�^]���[�GX˚۶*Rk#rُhV�(�Ǐ�J�h��mK�[��ٷX6�+ĴU�*
ZEعZ�c��b����:�D�4�� 7,bF�����{��t��Csj�v(��pےΝn?�-&�K2;ʍFt�V
j�n}��0M��T7Pl+]к˭���QK�F�aY��Vm�D۫X������`Ԇl�*aۥ�X��Եd"���2TM��1��'��Y*7G^-r�s9B��v�K{v�j�4n��t3G2�Ԡ�n�vm(�϶D(�E��|m�.;w)4]�y�Fb���Ǯ;�pC-��M��f����cMLWF^�D�Q{��H�L[,�F=˭b\���ǋ�q4Oѻ3E3
�+tL�b�n�i����,;{�F��β����#���"k{7	�3^ؙf��>���̫��K�+vn�ԫC7TP�قe�5�n��2Z�%��H�����y9$X�ub��^-�3����xdd ��M�vl؄ct���Lض�Lb�����X��k%��U�EƷ-�Z��э��+p�M4��kO�9v@���%���fe9waA�r^֠B��9Y�ӱg��<T"��I�[,��t`%��ӷy�R�H�p���63vF�����wF}*��71f"� �D���h����([�}7dC4��-�S,Jש�	&��k���5<`��kQ]���lѭ�o�c��gfb��"��)'0�8JY��4����K!��!������7S��c�2�Ku�l2H���	�� j��[�aP��=NV�Q�z*��iV��1ʼ�U��j,�I/�KN5K7%݁/F�m �f���>cI�3U���oLM�']�
��g+0�C6S6��ҷ�����5@|���D��t)v��u� ��[�Hܩ�YwJ�J�	�2�M�qn�������Y�JɊ�xMB��,2mZ�fyV�
�̰ɷAj���Mf���`0&İp,[�d�q���=U�蛍[�d�T�ڰv�.�Z8\��a��x������5-;Wq*l���c�[`�W�W6��˰CBO!Ҏ�] (�W�Y��3��`zpG2�V
ur^n[k*5oY���*�:������Cae�{P���Fl�lR����K���!�����	��YcqTl�"�%\w�lPPQӔ�c�IL�����8��isKâ
n�C���&����NiXi��p��9Y��ZgJ�VI�cJ3�6�3Zi��t�

��NƑ-�jG(ң�"˱�{�*�ܸ� ��T8��*�'uU�  ��5�U],��j�����+2JB �G4��[YknX�A�����#5j��a��:u�����ۭn$/j#�����@��]kJ��eZM�D���,�Ҳ�YrGVu�S`u�Z�K�:q,������E92�-��k�+�{S/3n��-
B؂��D���u��ZHIR���5�6����]�W�6;ǗT� ��H�uh�j&����,������s>& ��oj%Zޙ�)3v.H�o2��J�ц�dQ8�M�P<:ڡIcMi�.�g�{7�����_e�U2-��Y��Z1̧(�D�ƍf!�,�W�`�mt���kWښ�3B��ܑ��x����Q
�r�nV�vh�j8r9���wLhR&�];i�l�U �c���r@�YQ��WD^�4�e<��70]���R�r0E�jV#CjK`�`j�к�u`,����KW��ú[���)��5q��i��a-ʷڰ(Y��c��Nr�՚��ƾ� �3-N�
��0Z�S�J�F����Uj�q��i���á��Ա�fd"�	Y��5�r���:�m�Oi��>֎�� �'C ���(Y[���̼����iL�t�լ�^�9p���C��OF"&�y��i��SE��1��������N�k��1G�]:�̼V�[��g�ս]6��K��uM�M5���V-�f�Т����d�(�V�a��6�а�N�:7��u���S1����̕c��{ysn���'^rٜօ4�ӝ�����'%�c
ZT�`"k�n'WY[�]��QGbgm+�Dq��TZ]]S�F-��^�ت�n�d;/w;�9�.�E%My�/���7�f�����o|cޤ�CչnV��Z/�xՓ
wvp��b�u��M]���y�j��:2:e1d
��FvL�*��K�}s�k�S�p
�^�Zq�`F�\�-*D�υ��wnV�,��6�M�rK�S�T#�v{�k������_H�P�e��Э�*[���
��@��ϱ��0�ʕ����ur�}��|��{])�Z��)m�:�7r����h��t0}�8f���D��j���)4��|��D}�E�������9vݹr�����n�Zy�>�ᕖ����TF�YoI��4;x�gn��6E_h�쥑j�|eu�N��dZ��*�+����
�s#FS�B�;��u��ث.������Mh�;y?�A�vѸiǷOeʘ�����Ny��ӕ�.?�\��У΅ʛ:����S3N�<��;F���Ճk�I1�K�r>�u������~^s%qKS^������2�lV���
���X<A��X���rUdm+�e�2Uv2J͓+% �n)&*�7�u:�������'Pu|�ۖ�^-��`���ۛ�H�Ӧ5*���A����®M��ej� U�.�S��)c��PA%0�|*; ���Yڗ8j�[	��дSk:�32�)�\jcY:�,�E�P_f���Ν��ˉ�y�D���w�8�^`Ȧ�EWs�
��ݎ^�X��]�t �墀���8��v�_lR�ڒ����y{]GWM��!��"��uӎA����F�ii����q���6#�+�V��0�'-�coo��u5`l��<�Ĺ��̓�ģY���k����UnC�շMn��� ���<K\���ٝe����\�Xh��b�uᤶ2t����-Qu�9�y���p리P@��8
�ڽ[&R�j�[2S(1X���i�����D5����śq'b��S��(9kNP�%�U1R�k��*���u�ݻ&y!�;������wr�cN���<砺��W� V^��8&��eJ��ah+�F��{(�t.�ɾ�jVV�s�Y\�9�Dc�t�!�q���#͎|ɡ}�G�j�C���q�;����8���9��`� ����}k&E������T�et��k��мJ��g#�}A�CyR齺��˼ܬ�F��ͷ�uJ���^<Ep��ƾ���b�d��.�7ZZ��^ꬪ�W������zS���}������\�������un����%m��MWYW��-����?�+��L�يf�>���)yG���Q�q��qS=f�����u�O�,[_�Ҝ>e��N3Ȋ�6�'x�c]�y|��ڿ��О�!*����Q��B]���;���x!6d0�����@E��C��OUo]��.��3����� 9V2�߈��}b�����%�ᝧE��d86���uc�EW�>�tQ��n��"��Zݶ䮝}ը�R�v,�|�Xʘ�gMZ��8X����8�i�`7�SOA����V��}o�iYCV޼}c\�ݧan\��).��`��4%�Y`�lʎ��*�	���sջb��9�l����U�]���Oc���:�mռ��[t�Mڋ���tU^v��j��� ̰�%͖+(#ګ�*c���[a ��ԩnPY&�
)��D�v�Tˏps�̎7�c�^l\��/���;�v�kI���H��ٲ!2��Փ��֊�v��j�O�'fR�{��Uݵ/�D��5�b����7�{j���UZ�k��C;����>J��X��+aDͩ&�E��%0|����'V��_* ���0Eszl��	��P:
Gj��YF�M�)��3�>�wK+�"��n�¶�z�M�����}\�YP���<m��ܼzV.7fr3.r�JD�N�Gٹ��4�5:܈p��ԫ�h���v��40<��ܜ�ד��ݶ�:����|��u���ٜv�`f�fJ�c�t;�����]u�rKV7_kX^)*#�r���� ��h�M�.�p�dH-��ZɏFK�1\��̂��9O��ٌi̡�Y�i�u�uR�h��*�]����� q���>]}��Pg�՝��خv4cX����5_u!X!�5Ԋ�2�E4�4WJ��KK4u�g:�� *�p�w\W;�@�����;[o(�|��Wu�������W*�M�fk4�K���ͮݏ\f҂�����8��\��A���	���z���YW�
�s�H]f�������u�k�S4�ro9�ں<�F�	�h�y��Fn�u�ѵהz��΢�T�P(Mp��0���N��|F)�y��g�9-N�w,����N��o.�[���4[j��ʵ�[�Ȝ��t۸�4D�%3/�pt-(cy��S{5����iZw�[Z�J�mޞ��^:{�1���ɢ]�1�5[��������U}"��s�qΦ�����K�Mɯ�V��Q��X|��H��LsV{ 5�or��J(�v�*����%-�}'׊��7����T��i��7�+ľ�1]�]�ϲ��M#�o�3��P!�d����
ݭm�zj�Ywt[]+�[2�m�\�qO���<��,���[w��]���M�N�i�Q&6����#5T��əB�R�eF�ol�f�u�4S�k�Ӊ����w
{��7��k�;l�AR�i��%\��8����7kE�p?�@�jЬ�
ɗ�+��Һ��
��qD��f��͏Nұ
�K�A�Lk�[}{v�x�d�
.��FRi�,��Å�t�����vB�-'��/k�Չ���2ת�ti�0����X���U�lFT�������&wnE-[��,��`�yP�U=�p����1J0�y][sz�I���N�ѹls����$>��9��۬�y,�l�I�P�+G8[̽��n�UҲ��$�)a����sTBк���$ی���ge9p�Z�M��Dޮݲ��mt��kD7 �m���\k�O*�mC/k�u���Y��aW�Ó�ږ/%Nn��gg�gT�[��+�p!L�f��k#w�J�l��<��F���S�6�^t�1SR����,Z�__a�ay�_N���6w^q�g�4�+��`\W-Xz���a��\���⭇]��.��M�����mC�՚_�Ʋ����ὐ�K��V�jg�ڴ%����%!�<��G�ۼ�跛�bR���Nh��[Ó����W���yL���@�+ޮ�o��&�p�"��R}���#�]���j�C��z$c��.[��8c�)��am��n�����t��]@���d��d�6�V�t�t�"S0PllZ6�73����q�K\tPt�y�e������.�t�La�t
�V��c�
��JU�Ʀy1i��Ť�F�=�O�����i��@Z�O�[�#�������q,$����B�v����s{E(�gI�T#�8T�.�O�ͫF]ʻʘ�]�����L�WsY�G���6P�)e�fc|�έ�u�]�_e
}���z��Њ�v�+��rn���u�bҽO9):+��l�L����qW�Sb[nV�L��,���
�`��8����P�J8�'"3u�X�iҹR�llm�n���
%fhVnq5)��2�l��Nev�=�n�\1�}��
,l���b_�x��V_5���X��e���P���QR�;�8ch:]#�H�Q��ꆄ��KR�-����S�j��-��'�{�gH�7�Y�� �;�Yn�%��s���" �g]�'E:�U�áVE�)���v��VZV6�$0�¨����Y��ݳe��]ɑ<+��~.����1�0[�z�;e�O*��v���W��K�r�v���H�ۥR����[q�lRG��:v)u��
�Mٸ�N�@���c�ւ�9b��M|�+�6�^����i��0��_H5u[�ޚ�}WR�Q�w��o��|gu�a0�7��A��x0N��ֶV���:T�Ok�5�9}���������qU�B�grޡPvZ�ƕIY=��}�#%�/3M1���|,11�N�"�8�.���&�%�*U�s�gN�����D�X�f��K�\��ܜӉ��9^�K�a:��s5/#��g�+�*��u2�l���|��I�|����]�9���O��n�3�Op�{S8�>v�t�2�����yX�<M�t�=�K��3�Ŏ;靥��Uh^*���Wv��/���{mv-��A���`6駈E�/�8�iJ�E��xVP����v��������C�ю�>�Ie=���Q�����'-�e�hW�d.�NN�gB܈YEv7�c�Uuj2�^�RV!}X�N�L;�n�@������ѽZ)��Q|�t'�r����v�Q)����+�0��g��b,�].U�Y�ݎ�]�f�9r��93��m���eL�8e�#�VҏK�|���\�0��2��$@+�O7c��B�V��m6�q i���.�!y�tx�{�?!j_���+��i��Cw�8�����m�l���4�h�fg�u;s^.���r��us��K��O�/3K}N���ki�ui�����S�����d����{��Ŝ���g*wGΗr�Y��\�\;�OC�k#�䬮8����߹�]�k�̷6.j<�Yo-��� 
�ɻr�q=d���G��v$��aW/Gt��
�z ��?���m	}�,U*ܼ���
ۍ9�r;�>�^{ ��2Koi�n���9ۖUs��q��řb+7۝@�32.K��D"�ﰵ��5F���LW���|+�|'�K0��~̛�|�7�sX���h5���]957]�fm���`�Ac�s����p���7'z�4Ӗ��R.�Rp7���*\݂��uQ.��ȴE�����Z���:`��u�N�=V�Vf;H�ut��X�0�]ڎ�P�66�5Ô�9D�p����e��g\�c�*c��̺�e��(1u&@�J5�b;u��3�7�Nn�&�$:���D���{մ7h�V(�t��3J�#X:�W�L�pL"���N��Z�Klm�w(,΄��\b��dWw�d���a�1�G�|��m�]JKpMqWewƀ[��Ԑ���m�԰�t��yMo��Ve�K���,��M�ƃ�-�D��7���	�;v�֜����q����&�K�օ�\u{Օ�/Nb*�Y��m*W{}��gNbS�J��en�݆gCw��.7��.����9uO�
C9��q����r�z�mneZ*I��Im�S4���⻻��fuv�LƄţ�Z�sfi��X\o�9Iq��q�ii�gU���:gGס^^���y��J�����aERot:���;z.˩�d\W�#Y8r���A��	��t�v�i�:{�{>l�m�6o9;ҲQI�����t�8�ȱ���-V��I�:�bF��S��gr�A]l`�*E�h���¾�O�nO!���5^Kg	��K]W� w�w)��t*R�a�xts�ר��k�0^�^���nY������k��@A4^q�cg>�kZ�KI�mm�SK=r�5Y5��d�cP�c9v�R���z�6�
���VM����B�=z�p�̐�@o�] ��n�䆠/��T�jP�K/�$t��$5l�J;�!vI�E�C�w@]�٪t	�NL��M�Gi,A)ݷײ�0��*$s!�3}l���ng���C�fn.��+�����ZU�������y�+�3n���)�K����v��p��95FxKd�0�kZs2��2#���R���Bg &�V��wewm��!�G�4�Wv���lN��uySr	V��W�������+��F1}�*|��7�uξՓ����u����f�o�b:st�uu���f��U�b������W�RU�Cb�e�
�Oe�Ӹ�c]W7�V�v��.�nU��j�`�4и�
����ĀA$ ˵��a;//6��#�oX�������L����֞�.)��k��g*�E���-�>��S`�qY��Z����P�Z�[�����U�	L٧/Ty>�rA��Vʇr�7���"'��>���7+��f�v�wy�(��8@�ۚ
��VR��������틵��.��rq��
	��\Y�)��QRYw+�z_��������hT�'$I ��
�K�����̺�4\��Y	���<�t��5�*�b+��Q/[�ɣ�Ŝ���}��R~��3�?fn �'���ۧ���%��k:���
���ev^G�{]�����v����y�&[��t�nh.���[f,K��ӆ;�G�NOy^��y�L���J��\�O����*=�D[8�<v6�I@�s�AѼ ���t�6�K��6������Gsw�����Е8i�\��^���9��CrN��.z��=��J�E��@���1/��k^=g'�.��n�T-
��h������������v^-�t�[��@�٭��?�,|Ew(�1c�@��J�?A��M�^�$�
:�5�sA�Nx��Ah�F��fĦw
K��NV�Aa�������%�]���:��M<L�.}��+�o�;��+CL�����
cȰ�nupK��g`�7@ea;���.JG�g���]�R�,��۫��z��o��)"j�������vX�I9�5:��K|�����s^}���!���$ O�zk�0zx:K���m�����GG2k\�Eux��7.��`e��к���i��U���n��!��\���vgA�we[P���E�%J��6���M�w�)�@�Y��m��ݭ<�a�U�CRG.Ѧ2�;����ϲ�o]�Ə	i]۝Mvc�F�ɎP޳(r�c�:���N�k9})O�^R���1[vh5|(�������2��5s�	����'��g/� �m�o�e����V�]VHZ��p� _
������2]�nHw�ȸSr�2}�ݞ�޴`��EW��E
��:s$w��o�N�k�{��X�
v�0rάY;IP�%NS�9BmH��z�4s�p��:��h�>J��%���}n+��>�* ]��X_J9�_Sm���P7���)}�4&�"J�AHQ�5{��%��&p�-�\{��S�(e��u��HRؒj�3�Kr�i�,��vW+��m����Ʈ=�V��e��w.0�7�<h��C
�Z\��ͣ��Y����:
o�j�_-�CR����sZ/V�BY�tp��n�0�y'q'Ϩ�ۧ���ȩ-����Vr�*�lF��`��D�L>z�0A�Z����R�A�iS���omot��u��ʻ�gl��Պr���:ҍC.��R�E�\�)Θn�<���`��j�����}�,o0ʋ7���0��r�<�Ӎ̮����;�UΙ3s�8��gd]()g:�4g]��f�H�˥c9�	&�Qe(H9+�]W{.�܃[bޛ�V�t���fQ���#�q#kn�ǌ�T���ec f�t�铰E��D�V�'a8j;����;˕��Sw|qb*�P��:tY�yn��L�#�ŋY�3��R�����
�9�����8@���T4p����8�	4f��W:��Y&�����5=n�2��J!_d�Օ��w8tu�X�W#��W�ut�^���>�uOT9�nܝ��*T�V��m]���ӥZ)��q�6�I��۽�2M�CN:�/v�[,f����CvK�bv>��ю��|Mf�j�_V��TN-�l.�3�*�j��e�ơ]�t�8�[��[���-������A���sw�=Ӎܥ��5P�t�:e[Q�ӤY9�NPrx�	��E�wNEC�`�uV��ú�u��6�Y��hy��M;[x�v�*
�+r����yZ���;9>����TX��P��ΤUY�{R����`������u,��f��u�o2q��F��[bwY�o�k,���N���L#-�"�]����Tz���s�@��Ԣ޶޴q�M�3�uv���/���e+`�-(aP���vR���Rz�WF�{[RY/
\���|	/�s����lTݻ���9v5��{�i]eDo�h�Se>�.��%�P�����P���n��:x���v�$`�F�^��I���x��������v+-��cS��ɵ+�f�IT�K=|J m�x�gV$�l�(VŇ2�Ω����p�|��4ܗB����,F���cl����]����ī&��Z��p�+)q4z�C��gb!z��]�̜j�ۀ_h.z.��W���&=����B_���� -ځwj|Ү�X(�0�ynq;�6Z�@[ǯ9]6�nZ�L:�wg&-i�ɑ��&6��k�;��:�B���U^d����4񜑍�S�!n*[iL��yXf�i�S�3��!t+D����ɂ_
��Q=b��1�յ��EWՌu�"0��V��)�txn��u�vڀZ�/��g[������UjHˉ��Yn�X��q+:6��6���M຅osX#B��{���tj�L��#΂������Ə1&iN�Do $��C�C�lɑa�r�[ݣ,2���]1L.��BJܛu%*�Rb�L՛I�.��Y�Bwud0o5
�4�]k�c_ea���`(� ��!Il3fgS<oz�NӼpTŅ�} ��nҔ��R¾ZӒ(}��+T�6��-"�򺗔),�h�
)RIX�:���V�6���h�f�ʰi�u��(�
3tЋ���]=�ڥ���z-t�u�ul�]ա�i\�ctѫ��w���{��
�1��)إ�y����^��C�;���ۈ�J\¹�)�(n_���Yg�9f��O�:��qڭ��3�jAm��f��/S�Ү�6�RYhPG�v�C��% F��*/n��^^Kie �Q*�-u�,T�2��J9]�� j����q�ْ��whM3i��r$6])|��v�ʕm���VV�!��)�M�bZ���5�4ް�Fp�X��A�.R�Yܶ%f�b�k6�+�9�V�xd�-���Ь��o^�=l�AI��ÚbQ�W��u"gT�׌�=v3δ�F_t�>�Ls]�3'9#"���'Π�������erUsGw\uvp�w;�aw�E:�l6A	�oDT���vNN)����V9Ю��Qpn�������"���Z��}:��
ix��V��V˫��k��mS�y�>����(sy��Ep⦘�k/`9��Smְ/���۰�W3L�.�*J��J���5��Z'f�"ܡ ��.��4��=G�}0M���q.��ڲ�el�9��0S,b��k;L5���y�P��V�|!̽�M�1��7Y����L���-y:��VR�n?�2(S4�O�K����p3�y�]���0_P�,M�f�����TB`��(vxF���}YO�8)�n8c�1+}:�3#��� 9˝8�nm�	�=��ŏ DӾ���1 03�ȕbYٮ�V�tj��<�HV�t6��A4w��1Qz�*�HS��z�j���@|�[��%9�X���xmϵ��AV�#Zo:�ǯV�-�\6U�Bg ���bg�n�SV���#.w2jK��s�����m]b��MUŃ��幢��:���S�����\���:��i!]X��.W)O�є]I�N��F��!��[o�Z�o2��
�j�\B}���Z�I��Ɲ�,V�s�bbUz�\���q۬����%Xð�]nj�m�/�1��Wц�G�6����;;��dL#b3;�*�*�k"#\�d!v��o@lN0��x����\�J�Q��'>b��p���^
�Y4Tp��iE#�/�ar��~a�_EG�����tﮢ�劺�=��1���i� �o�zx-�M��h�3,Yv�JF�����*ǐ����9��}V1�^mq�4�]6�gG�%;3Y�J��������I�Xv��|m�%�(�����ѯ5Eb���`��*��ʙ�ξ�O33)�ꓨ����%�yp\'h�w\QcC���D��۩�:����|��S��G�t�W��q��fJ.�m�)`f��lM�n}{�m$�`G�s*ƥbc�i���sz���Ҝ0ͻ1��:h�a���wl���.�7�Ҵ��c������wQѮ(�3VF7$�`�4g9�t�M�T�t95�2��,U�Ӓ����|��}��i�-|8q>	��{|8�b'��74���-���m]��e�ۛ6�%��˹[ӛI(�Z�N<&�ʼ2nr�;n0�i�Lj�3"i��y�.���%�"�g��]xj9�qnƊ�m�s���i�j���w^su�]َ�[yL�Ƌ[҅�ݵ�/:d����D�V���0�Wo)R�k���{��VV����=����{ݙvƸ�-v9Mɗ+ydi%�	�8�&�f�t�l��p���gX$]��S�o]G �:b���kt����:�/��GfK��b�f�XD��4i:�zL�b�N�Q�����탙K�jI(�1=�[m�k�j\�vJ�������´�_0�U�c�V:�E���+��C]/5�b��#�)��m��*J�Nh}��e��[�a�� *�ѓ$���֗9DŇv���+:1pp���n�z�YӜ���$ԭl�����޶����y����l�W�y���S���n�S �R�Ķu�l�9wTqG��1�ڶ.����W��ښ�q���G����f�8��[nK�O�I��l�#q��}��
7)>��򴟗P���!����똠���|�Kq��j%����['��a���k�;��>qPbT�%*�7
*������C�յ��Lb��y1l�!��6Q���Wg%���4'
�z�u`\�C��}�,Ôn+�R�u���hT%s�w�f+Z�1&n�t����6:=FN���Jt�cpH{i��'���y5 ��J��: ��/Y�D���v��r)A:
gm�{�>�z��C�v]��W\����#�J�M���cH����g^Z�8*�}E�N�mi�^��"|�#H��p�e�֪����d퇼 K���|��p�xF�N����K��\+^R�\N�X�:6��lj�#) �Z�D�n�dVQ��%D6���C�O���tV�ͪ⻺�I|�ᎄО*� �%�]��r݌�`�`GYQ
f��ϦlGEg.�g+A�:)<L����ڵ	Z.�蓫)c�Z(ܫ}&�̃.���G�[�}��_i��ᛏk��2o`HZkH6Y��A�*;u4�Νtђf�꺁f�K��6r��J60�1:�m�h��k(t�f޹p^G��7�ҙ���`�V 7a����M�2ս��A�I���s�z�5*Y��z�9�)�6�b2]�+b�|�.�t��Ȏ+��̤�ekю���j�%_}���ҮC>թ���%�HԪ�X��6��K	<2�-	�W���tZ�j�
]YP�*�/78�(�s�B7�*|�]��R��v]��޾W���.����b�eNXn�w�0v�l�!��(������ N'o��Gӥ&���v3LwS�*�-%�����p���S����t붞�v-�ʝ�[��eL����{z���m�#>�]ާ��}Q��X�i�++����n�"�;�O6h.�.Vڌ<J��p䬻�k�|vf���@�"�6i��:��$�¶��"5�Uv ���/�k�o9��J�1�-���PY(]�h�c�Թ�\V>�0*���Fͧ�VXͲӡNM�{�&g��CfMrmohq`wV���^��O�H�\�"狢�m:�̛�5:Z����}��I�j�Dq٬`���V�t���=J�GS���u�K�6����TO�r�i����7V���f��h��Q�j��',.jU�U��Ռ�x6�f�gy�)1y�r�wa.�*���b�w�����B�M�]M޼lR�V*7��"�u"7�c�Et.�we�N��,es7�=abf&2��&Ы&���ҭv��:1%�n�(I;�_,9�v�.�v:!�Q˜4	VS!f�sG��{�Sr�,k3ܺ[\�h��ӈ��kk]�e'��d�w[r�?�t���v�/�cV.@q�M����*I��R2�^֔���/��(���8%\%쵴��U.#��%�dۼ�L
�cb��ҥ�� z����"ubp:��`���7���dpe$�:tT��|;�����un�.=
\�=�x�=�L�%�>}9]��b7wJ۾���TM-�ګ7C�ҰQdg�[�ծ���ψ�.��b�es��WV��cr�����;� !'`ڶ��W@�֧] S^7��*y�`*���Ua���n�%<�ɽ6�+ m,�[o����^ڶ٥S�H{��V�*�ly��j*:�$�W�e`�6�Sicp�������S~l8� x�d����?B��4|��5�k=���@C�� g⹩\6k)J��gMc�J�[r	Ql���TV��<�[��݆�jX� �#����"f�����f�/�ZV�j�V�<&�tz/5��{R�R��:��(n۷���B�<�v������+0Ĝ�ԗqw�����
O���`u�q�-�(��̐���,X�W���`(�J ����;�&��V�0�+-��7��PWR�4e���vyPA����ʅ��%Y�;7+\z���tg�p.b�j��������L�+C��r"½7��H����e��z4�{�����Ȳ����P��ն߸��e7N�*�>����)��r��T���s"�܎ݬU���	cl�ۍ��o\�M�D=Y�*_L��8v�-t'������3lu.c�."�l�k���ި�/���f�v���C���k�>D��R����/�qu�0�1W,`IC�se3��q���(<�j������ig�Si�O6��.f��V�5lb����i�4�l�G��1=ZJ֝u1�������:��4�9�wW']�m�uκ�ߝF�׻���_
�.����D�5�4���s��/c���^RM�[Q��V��]i�����m�C`��HOvl�E�c�I�aj��uZr����B]C��toe
,Ƈl�/z_t���νզm��h���+Gf���3

U�M�ӬJ�9]�u����D�Y�Cy�O0�K4�{˷��W�[[�l+Mcm��Un�{0��V�S�}�	u�Z�ô��A�����ז��'��]�ob�Z�#X��F�Π���
�y2���0��Ь��+`��^Y-m����桌-{W�����=�v���Üp�
]V�ua�b�:���k��q�U�,hj��R�`��&�z�oi	;����tSo-A (vc<�q��۶�B�V.%,DD�7��YsbcGk +r[:��,��v�)�]�<�S櫺�طNݪ�㹹���ß4�E�&����	:� �š�9+�$����j���gu�gnf�l��}�
+n(MN*m�C��!.�.�yGc�[���fM���w��{>]8bH*ݧ�&u=����oc��vsܺ����o��G���G�ꈄUV��dڎ�Z��-�wvԀ��[�[�;]c����^V@7�Zr��X��Z3�fd��35rНJ"].���>�oW^��k��(o[�J�DQѤ��,՛�n��]��.����i�����v|��-��iv�:6N���|y�Z6�>��ۥX$�I3W׆�.�D!�qj�ܸL�f�0�؅�vJ�G F�O}v&x�w/)� ��OLc�D�=�P��`��j��x�:�ԟ�ⷜ� -8�l�3��-��2lǹ�oq�������-�]´VS��[���Jr�^_��N���v�Ň#��|ɾ��vĜ��9�u��ȓ��e^���]�����}�uu�j�@lV����䮑����|yr-C��њ��Y[��>sx����l��1j*�kw˦�
��u����2�r�^Z�A�[�%FM�4A�JĮ����յ&yf�ec]��U���̚%XNS�@�j�\7Xx��7a�L)�e`��s+�lV�S�h}���c��E�J�PwB�rEۯ8s��=��u�I=��|m֕H$p�N]��p�WZc����kW�rQfc�Z�����M�җQX���+�u�I�zG=��Wr�Wo�_e��l�o��k���9[�;�0[t��qε9{/y�v�hBN0�{7lU�@P���vꆮ��6Ԃ�R�N��|V�r��=M�2�.W��GTf�Q
Ň��#Uʺ����q ��ŷ���X�^�X�'�)�KlH��u��qDQQb�
"��"��R����*��AF
"�,���Db�1F(����(��+UUX"�1X��eEV(�Ԋ �+UU�TF"�,UT��D�EX���ATQb�b�+mDUTE�Dc[U�(�UUEX������m�ATETU*UB�VF5*����(���F"+"���E�(1�Db�T#X���Z0U�������j*((�EUb("���QED�KIAUET�Ab$EUDQ`�#Z,�*��J*�1Qb�QDQ��,PDb����""**EJ����Q�EZ�P�F"
�UE�QETe�PEU
�"��U+AQڈ��Q����E��b¥Q�Q��"ʔ�b�,ciU���QETb�VV*"0Q�DV,E���Z�W��"��hs�gks:��4i]�m�5��kr��%ӌ,ui�:�B�}{*�K��뛲Ɓx���x���2�v��Ek�8.�ƷM>�kR�mn5�`C��;��Afwh��l���f��v��0H��	��i�����Gʦs���Gg�W-��rй�'D%ʶT���z�F���f�'�i|��C�Uk���Ӂ�u8O����=����X�{��!ɹ�Qo�zE� ��s�C�Z+�::��1�&����(�1w�)>�����DN�uXn�PK�b�ǵ�K���p{�o�C��/߼�ꠗ�6�493m�z,Z+��3��4f8:����NR0�W4\�<|�WPr�&8(4��r���aMD�CcF�s��r����b_��F$9���M������
x��֜������bӨI�*cx�"�,M���|���=o�K.�R�p�o���墽){��2���4'
򔜘��{}�&B���x�|z�2){��W�QA�5X3�'D%x�����K�1	�K�{s�����gJ'l�����b��x���%�1d�ˌ9.L��4�7P�k��\���y� jtP[|b��s�BȐf�<����5�J��@�=ƥ�����7��-�S�l����dZ����z�5��n�/���B{�Xva2^�r��	�ݓ+�+��u��)C��,�:�VS؝�'���G.L��������ʛ��ӹr��U^}�#@����|���ʎDV�!�'��bac�u8)ͣ!��e��T���O��E���.1LR�}&9;��؊���}u4m�mD��.���U�:�����g��
�z�z�@�*LFS�t�Cs�RЊT�ϓw��g���O6�JG��睚8�e��~�&��٦���X����1�u\��Z����x�mi�Z˧�i�۫*��P�{%�"W���*�M#�N��j�M(��P3��#ܻ�9��i��[\R2���༗�p��RdOJ�|�-���	�cp��0��}"Eછfi�����y��:G��pg�1�Z5��(����*��Eʑ4�ۣ=-����B:�{;��F�6@��K�����L'qS�#Z<�M-�%Ł<�8+f��9�p�\#�{���́]E2��.u:�ni�]���N���9���<�q��R��2�bp�5�	����c��9�C&�2��\���tܚL�M�WB��.t�m�/1�-�j[H�IKB1��3�����m(���K$�����8]-�k]�"p��u��q��,��5�E�E�
z� ւwr�v8� �Ic�y��X��ϲ���)U�頠���gR�����;y��x�˧ycP�v,�V���.��-|���
��ʁN(X<}&�la�ʙɨ�όNʱ�;N^�*m�����7�S]��=g�{+�q�F�+��J�<�9I�S�D>�����}f�{l����0N�µ�ʼ.�MP� �4��D�z}C��K��{�ķ���֐bn����/c�b�o�{u���Y�W.�	�c�t[A�6��긨��S
�A����1Z�᭗�F)�i>�5�)+Ni�����=�r�
/�]B����Q{�����6>~�q3�0���H��F
��dQ.P�2�o��Raݘnj$�3�k�r�	�y}�iC�[ޘ��=����ɍ�,	��t��s��֪����1���Y�ծ��!ފ���v�xVi�o�����ؠ9�P���K����.l�����Z��A:<�uy��
�=,uܡ[�az{A�j4)�|o�ն:�*���f8�G4n��G<ʝ�����6�U&*vZ�}i07%��:���:������S�cPj��^a�Z�ƴ�X�w���>�t����r���yʳ(�i&2tԂJ�0I�0��b�P���2��p*�s���!`���iZ�f��I�m��p����髓��GI�̜�w�Ri݋i>9�]{;_�5��Zٯts��:����u8{yR=L�`��9�'J�])vp�v��!�=��Xm�lu���hY.�W�0�)�����gR�D&�:�N��7Z���85s�yբ��B���7Չӗ)�0�6�ڛ6ꫵ�M��7s��j�Z���ФD;[��F��x^�>�c�199)ݻ��	��;I^i��x�L��o��`e�̩���ى���^�en��FVk�O�S7�Q��#�M���G�J)�Ʉ�S]W=*i�ׂP�n0=u���T\��^:��+s��0p)3��S7{N껃��E֍"�����&��Xn���
������r��>��-Zd�b��4��SS�u/{bM }��Z�$=�"���5r�:>1�Ćui�)�3��!��lu0�=�XP1������\&z�\��c�B��oa:�"8jca�5�(Ξ�ɹ��7�C��7���0m���A�j+���.@+�����h�}��Zɶo:{���U���gem� ��ex�TmF�,xuʷ�
w���E��6<5��Ե�j\~���h�r�귊��_�ʔei3�#fـ6��fH� N��fxԶ�Ip8o@P�<����sNJ��/�y�kT]s��̋�K���V�6�����z`�i��cK����m@�!�끃'%����E=�֊u�;dx2m=覼mć����.o;	j��FϨ�VҾ4E��T���$z�
�n޲�W6�S����N⨬-��n�x\>��<�8��zz�<�=5&c=YP�v�YО(��qT�Á4u_)�ℾ�Ø����E���֍��e{U ey`����\�W�x��	���!�8�[ ���ߨ&�IcSg��3�Y� ����Bȁ���j&�j:���~�G�POp�]B�TZeM�].=
����M�����ؑ�ZЖ��~a�ǒ�M��`%+���wr���U�==)j�	��d��X��]��)nEx����#�I�ԥ\1�q� �Stj�PL[0�XӶy�	�˽�9����9�S�/��׈�&l	��RNV�Y�Fm������K��ٵ�1ڣo'$zߚ:���X,�V�7���گp�#�x��Uf���3��LK�S)C� ���r�a�lu�n�R&�
x���ND�ẘ�` n��A��^*�]�|�r�*f���e���4��X�ߒ���}��"�gd���gbUWGqF,Bo�U��5Q3��g�uE������CT)�w\H�k#Z�e$G�t!��+�[Zt93�+5%YN)cv�F���E�y��<��iYc�ƯK��f0���N�r9=R�yWL;������N�ew�p4"��G<��AVi�黕�Yc�����пY��^H�sf��!5y��!�����FT�D��Q�� �B�돁d<70Q�9.a`��L����gk�c|:�m��\1�	�ъ��Ɛ�A���1����RX t��V Y�CVc�8��v�Z��8��sR�ah���x`���Pw��H��3��V�<���gBJ���凛u����6wp��ub�NRP5[>���rlEN�o�NW�� r���ix����nH4�6z<S�KX8X�b>�}��tf�j.����n��0��
*2{z٫Ĩ'�]p�^>|0x��)t2��:����
�ʂ�ÍL7��.=j�C�Ib_��j4�gwo �<++��7gdI��A���鳄MJ�������ᰮ��`�����#�Xk�S}��n�
�C��*�Ҩt� ��7oa?|�{���P�/G�vZ�WЎ<����<x��DF>�����1Rc[���/���_/����s8s4����4���.�Zjki]9n�e�t' "���^�=}������F��λ6nu��R=��Pg#ӈ��G}{��/�d�e:�6\���v�3r%J�]@�Dt���W���|q����g�i<C�j��yUAҨ���t�A��	!�T^NM8kn/)��p&2�0����=�Y��q`O 4^�x��=7�����s�=��B-b�����j���;8F���w�&5���t"j�wr�\z}d����O���Cb�D�1��W^`l��f�x��}�U��δ�:�d|UD�5vj��bc4p@W�J�g��^cM��NX&rJu��(m�r�w������]���=9a��S+k�Ztf����#����'��J�D=�>���֠� 2Wv�Y��ᯰ,k3�{�U=��SW-1X�ȓ0㇧B�ٹY'a�9Ig�Jg�+Z�v ������] �[��V�rb}�z�>��iD.�ྱ����o�?#��JFj��9c��ŗ���Y������1���.��5X5�'o�F����M��WFry�]NeNB
��-vx��ҷ��^A���.Ŕ��D�+�V����&@rv�:u{�z��sJc�\�{��Q�� �<(^���\x� ��¤Y�to(���Q�� L�T���f�s��� *t��^!������:Yt0�W.��%T��pNvV=�6l����������.��*:�n�\S����{'Wg���u!\+�CΰS�8R��g�����t����+Z�j��͇�veż�Rڜ��R���S�k-V0h!�TyX�C����/D�pu��0w/Of�W0���u�ޫ��|2�#s���
����zU1�H����/�-�*t)P�����d;���s��E�Fl��!AuU��*]u6 1s�(�H���K*n�t̠9����e�W'I���~�A�0u:�鋎t+��_�0�)�/"���Y��ڲϓ�y��`yC9۰��bq��j�v[*n�.
O�龬��˛��L)�1�Zck�Ŵ��C/��UOЎ�=�*"�lC8�71P�㮹���N��OP���1cێ��M��y!�w%��������7NC�}[�Fa�x*W��}>���G�qw������x_-.+q`�Sv�٦^�L7����>��3�W��0��+�E��@�SР=�.^�����i������t���Xʸ������s�ZT����s4���td���r�R��l����B�]ډ����tTÖ�@9���V�l�s/�{��3z{2DM�ֲ~��<�s</Z��m/I�r)����ǳkF.�{J��
�=�:Tcq��5�� V��-F/��e�F����:���7U*߻F�$�&;�O:S�&�ւC�2B���;yG���2\�K7JnnVp�b�yt�%Ted�H�sq"��R��yĹt��X�*{���|�vg�����E(%��؀Ϳ<:ȼ+ 5�v�m�]l�]IL۰ p�U���j�tt�� ��qu���>f��˼�q��>�Ff�m9�r��2��Hz�_pL�����vI�ݝ�Wʰ�����R�*�]�[�S��L��Qy�we��
�{���L\�����"�}�v����V*ZWƈ���:oD���S�xښ��6��lNΞ���=�c׵U����!l�l�/#��u���<�����bWW��u�-���(K@�Ø��HIT]�q��{Ļ�=tlc��k���K�d�O9{�$��G�8�:|>��u�����`�Ϯ�)Z#qY�k��*�k�ޥ�襖FOQ��cS���.�g�U,�B�U�T���A��������5h��)P.��Xvm���~q��T�e�7&Ez� q)_<p�.n0t�>�·Q}J��C7o�n���Z���X��{�Iݪ��^�Q�̮���ߤZR�����]��r���Qn�F,G��mt�Њ�d�%v���L�̘�Y��ev�����N�6Y]�\�%Y�ѵ0�Mv����ճ�geOغN�d6rD�#�IJU�Ȃ7Y�[�X�w6�бs��fIЩPe�m)k-ߺ]��Mľʩ��l	�����%Hܭ��ћn�eF�\�n�s�^*庢�WRɋ�XqW^%"��مb�ӚpZY�{W��C"%�V�W�C�(Ig��O�[��c�eb��5pvM�TnSb,�麲�9cj�}��Įm���@Ƣ�6��0lš?I;e�������v}lU~~�1�@���WL;�F�=�i[�0�ܤ��Evm]E��Jó��s
�ƒV�e���$:���6�q�*#�r�[]6tg�n�W�yX�+�q���[�.9N�����5s2�\Ԭ�i����j1r�f��
�v$�4��A�yU��|��Ϭ7�j�&�!�1<zl<�����fUْ�����c�R�U�z�����_$o��3Е� �r��"��;Ϩ��-�=S�O�ڱ](��]�=��/���c���^�6���dz: ͪ�O��*�t/�sTӾt����AG&Y4��=�����ʖe�������΢*����;���}���ַ*Z�6&�z[��v�$��c�VK#73)�Z��
�����K0�iV�|X�-��3���mH�T⣱�v�:�����j�wKZ���Lz��;��B���r�d�Mw�7��%o,w�T���|+4d�-�9*�U���Ԃ3h����Խ"�m�������]"OH]F�
��h	
t;����+r�p�]׎rΧ	]H$�NvZ���3���"��Z�M��0��0hY�c��H��n��7�;��A�w�J�u�8�[Sz�Q�{V��l���ZA��۵���EJEv�D��W9$�C����G�I�* iv��C��±�U�=�2���q���9:��[�m�x�4��`�,|�v9Qܾ�*��'h�1ݬ�iM-���C��s|�G,�m�ڟ5�J5rY��"��8A�E�#cX��v�f��1�� (r�]%<��di�K,�!�u�u�)
r��<�Z���oC��F���rdT�ݧ`\��G`���L���X� k�{e���Ӆ��z�i���,���aB=J+�u!�M�k'�@�
�t�'q>����z�i���S��wl��T��\w�%�L�rM²��3�ǰ���N�#�.����9���}{SP��(ҏ��T��ui�ڙ}��r�f���׮T�K;..N�˨s,\t9�)|�[x�[#[)�Ux;���-�y�y��rBhȏ;cel�J�k�HFJ/Nf���clΆ��3�sH��:�7����f�.�ڛG2IOSޚ��}U}(��a�촲�Б��g]+kh,'��J�SZ��G�7@���E�6T:o2aB��6���n>Wi���[�7�ef��wA��.T~tV��MM�#�s ���+X4��v�r�5S/J�T;t�tl���J��N��0��Е��wG�F��腕%��(�u#x�qYk���Kɢ��Ǔv�{qB6�9�B<n������f��OLK�Tڲ&�P`��L9S�[�`�w�ѸХ5���k'̴A�-��B'�m��.8l�)���>�PH��4�:�G6�c&>��M�*]�7m�.���h	���]����;� ���^Y w�6,�����<#n��i֮w�u�gWR@�8e)8�Z�+)R&�r	���R1�n�f��G�kjV��o~ŽSG&�7yۮ�q+�F�z���W]�����Z(��F3�yJ�R
�.V33��T	R�4m�˂��A�r^铏N�h�y�u6��ų��5n_k���6���(�*D�(*Ec-��Q0b�EEQ��X�X���0 �����c��E��EVDED���*Ԩ*,DU�h����EDJ�##VAZ��c�QV"�FF �"��V"��P[aF)Z��)PU�PLeF1TF**��F��\QDb�ȶ֦&�µ�)*�Up��Ah���ms+���7�֪���Z��G.&*��EX� ��X��QPUX��b"��ETQb��\��#Dr�ɍiX����1b�b�H�
!hPDb��c%�1R(�Ŋ"�"�Ab#ZE��UDQU�TAFT�0\�)EDQ�:?\�������w��s�u���5�"����u��D}�?j�}�����T�rs`�j���6�-"�����f�|�oy[�(�륎�T�S{7���!g�V�̧�q��Ni���uF󚋿&v}06aD8u��3��q��Mp�<%L�J����z�T_��&3�>Lf�\���A����
0�J�\���+:�h�=�LN��#�\MP��`Š4Kn�u�+Z��w�8`�d�9+S��c�l�0�zB,t�lJ*��%�fm��78������eW��S��<��U��>Ʃ`L�J�@�.z��c�RUYG\7�fgb�f�C���� �R�֝��b=0}`�Ld'Ja�U��顏�˹��~�M�M�2��#�ޭ>q1�N�h�58��Lj����m6�3�M�j��N�ǜ-̮�Ot�r�W�z),�6"\5^Pa
� X3�U�����P|�y�L�Qʖn��d�13V�z�����0e�Yq�
�i�. �zj�ld8!`�V�{~ڷ|C*�>�U�l	�r�W]�ڜcD9���i��Y4�J�I�t�'��JDC�2���z�6�Q�����}O{�]:��FA����U�m�A�CzrE7�}�L���{-�
���Ky��!
ǁ;xM��9Ѝ�� w�Ҽݔ��&�!pz�oT����Gd/�i�bS]Ruif�=XoL�
){�8��ӣfƭ�
�KF��G:��F���h�6�*����_}L�I�{4况�S��%�� �Q	�ۜ�*na���r�N�r@וq�u��U�t/f�ۇ�fe�QKt+�a����ʧ?��O�6�`�r�l��7LĪU#������N;�o{��n�S�RB�VOhf�܍��1��mB��^�n�[p.1���.��s�����.�uwM�@�sh��|H���!�����lxzo��N�аuה��u|��sǆ�[y���=M]6�W����׮�nW:�Hz��v�e���*�#���of ��ms��Yk�\<97=���Y��N�H���������K�2���.�v*��`K]o'�P3I;���T+J�j�[�;��C� h�	t�ٕ�u	K�ZW�;����)�,c�2Q�U�.`�
C��UV�n�T����:����'r9/70��U���uJdNJ�:X��<x�����z*i���C1��<
T��`Psȍ��UD��S�m��3��\�>���:��*�T݈�
M�7Չӗ7�Lt顡�wa��q�>)y�pU�R\�V_��P��ڏ�u2��=�Z[>���^e�7'oʣ�Kf�[�����-���a=�Ȳ�ηr4��Nr��{���ۢ4ҩg��z*��e���Kz�"�X	b��j嘙��UPM�9�]� o>ߏ;�l�п_�G��Ћ"\\J���[�����T�{_R����������'������ub����z�"�~�t(*�yxQ��ҎV+
F�KĎfi�p/b�����i�Z:�S��4|^�M�}�p��P��j��=������Z�v�j�xr��G촺�X�+����9z3Є�K�9VD'w50}�D֕&2�WBI���J�)��j� �L�1�Ȑ�s�e�N��K�1Thg[�� �n߫�nP��Z<�cե�^�w2�	���c޿�������k²U]A}��z��v�FmĶbhd�-��w�0��]�
��j�������YxrY�/�M�QQ�#iσg���z��}���R'�a2㝝�M��h���}�:�_�P���>��
w��W���;��yr��N7���d����8;�]v�]�~�0��v�)yh�@Պ��Wƈ���m1�T�L�[w��Rw.(XW�R�C�AD�_���c�m��7U�e{UX(���hsѰz<Neu$����U 7t+����b��\Pv�9�;se�¹P�9Һ�ո���T�=KJ�)ns2��q��O_[w���v�o��1���D�y )'p��w
�v�*=�����7t�s�w�us�Ӝ��9��۳�����m�����G�=���p��w#3���PFJwBR5�s!����d���x���e�|��OL�o�=��$z6��.(ٙ�"�l�l�Sq5)�H[����)�#n��a�c����Q�8����,��tx)ȣW�(�ܼ�
|<S=:GpJ>s���{j��}�Y�M�k>����b^SجU�c�u���;sr`5��TJ]Q]t�2�r^ȩ��Y²d����ѣ@�Z=�n��l�>B:aD��ԥ\1�q� ��5��V6:������/zZ]����T982[�w��Oz_���&Kl���������TX;+�)���]:r�X�*�>�Ҙ�لGz
�款�o�hs�gbQ�����*%,����9�b��S�Zn�E�4#0)���ﶬy��J�@肞Z��J|�Ez�'�;��.��JT!O#��3�:�8�'��������؇�un����M�g'�A�&9WL=�UP;gf�8��訲���֟W��˟y|��g�+n�p�)-�Dl�Vjq����-�T;��I�8�!���*���N%נ��;�n2�fǽ����,:&
��x]`榼6忭�˳��=�.����,��A��վ*N���LJl�=J���vɜ���Y��B��}�̿���Y��S���5/D���S�`]���y���,�p��W�_UW�\�W,+}��'�u3�����:&�y�B��< ��+�_��V}fQj
뺥��C�_��8�f6H�<=�_�\�I�4�ΐ}�V��}�@���jp)^�u�,z8r����L4�+�`������(�k�q��s����uY��ѕ���/��3���7�lW��/�J�lG��j�t���{�{������f�Bb�EN��ǽ�@9�ޚU�
�Zʞ,3�bo���~��V���Z������q���:3ܪfoU�Cj1^�O1>S��J�)_ޯj�ª�R��僀���K�Ǫ�=�����a1������bּQ��^�76��M(�[����-��6:l��.����[��]4��5m��>O���H7u�w���iZ�em���R��-p�-�m�I\���~��yq1��_t� s�mצ��Hwb*zWJ�����'g@s~��!&z��C���t
G�;y�Uxw�6�"�����˴�T�6,�aL6�7�|F���|�rc���/�ݽr�r:+��ze)7�C��T5��#���Q��y)b�JF�e�>�-��J���I��᥆���ް��R�X/$���I���|��L��~�^u6L
��H�n�)�f5�Tv���L�<;�nanoxI� \*V��ވ��X���t��g�К���
�[0�LcN.b��T��h����u��������7tzk�'�D�u��� L�4��#|�.�P�>�NLwW1��fo��ͪXy������/԰���%Y�����V|��`�s�2!�uh
w��-$��cFB'�`X�:w��ZV��!��mz�'Fiv�J����ߨ����	��s��x�}�#���U�33�S�,�)��i��70�ҫ����ʊ�r\p#�� (l�/�o˨��gqxApӨ@�_Mi���Ⱥ�>�қ0w�!4=�no��]/kg,e���(U���+p�K�L��`����u
+���Q�`��h`����䟥�>�ܬ��H���!��g���{��Q�5=:ǔ�
��vN�5�c�f��飺����/�E;��8�\)!O�]�����8��P�;�Xc��A	�)-���(8Λ|������b͝���S�/�F�H"8*�W.϶�E8�=Pu
e��t<G��Ű�=9Q�(5z�#��]�"D�O�}3LJ�	]�v� ������)��N��� 4�٘-;|�=�Q��]�Һ�����_v/��Y\�Ct��g61uE�ᯝ$��Wf�r�!��X��;oUL�,�o;��}��}�ěsĸ�՝���=��X�ϫ�ҿZ�sF��/�ס�5@`�7�]8{�kW�t�ٝ�S�(���r���q�0xR� ��ӕ7ۺ��N�H��g���o�&=���~�f� L`�WQ�p�l��)1�A����L�0�g�4nh��u�:�ż�C�5@_�˃�b'�`�m}���	o&��Ȅ�˘��
� ����ї0e��|�7yUV�qr�"����0���E��W��<u� � Z�7t��8��g�)�vz{�j��p�Ɏ�F&&��!�����vb�*��YPX̉�#l	�4�/����m��R¬B���������[�3-��)7�X������n���$�H/�V�e���7 P�����g:�@���|=��u`�>�(���8�P�}�|��JU��Gs��>y�E����)����}������sW.ӣ�.LHb6��-S�����H�֣X���8*d�N	�S�c�z�����²]AV�#�}G9_� P�=�v��i3l��
r��w\[%���g}�{��X
�������_�U
�:޼�@��~�{�:
WB�ћC^�Q����Rcoom�kh�Q�?��K�w#hjgr�Ρ�Iܖ��nM�]�!�{�'�[[��b}׮����]�uVB�c 5�nڱ�����)�iw�����{���kA�̱3�f/ЄP� �{���=e
a�[��x���gb���k�g�_��bv|�<5"SXL�7gh����:lVƘ���V_��ϧ
�M3x���(��r�(�.2��u�����v��us��pt�Ȍ��X�s�[A��i��(=���q=&Y�^�
'�j+��b���mVi������d-�Z7�����n�ʅb��18l�R�Q��0+8���g�%p:
c�!����E�l�6vz���U��ߦ�SU���^��^����Y�S@]-\>s����x@�{˸����9��(�Cvm_N��^Vc@0�"waת�
U��q��~�aO�t���Ѓ�];<����[v�)n:�_�͜nxß�����|"���CQ,���j+� TJW`����p��"��[�)�7�����a���Jk��L�۷��B:aD��*��A�28:��C�H�y��ʁ���Z=�D��7�e5n���*n_��#�6�h���>_���&V;s����>�`��eH�P��WX��ծzv��#k�ilVm�
r$t�H�r�H�+���JT{��y��j���>}Z
�ŗw�+[ܓ�qeE������D{ވ9�kg�pa�2D��2x}��I���.�5�/�����T�L7���<߂��Qw�ܭ$\��S�WL�
���-����b�f?x��:�)㓦�{�U���W]o</��yc.'��TĢ8�9��1���~���e&:n[��R��h�#^��ܤ����CmL[�F�{�t�$M�mש0�<in�Zj�����`�t�8	�Qf�K|􂄮F��tC.L:=f^z�5� 0P�:��`V�ȹ���28l�:�֔�S�:��K�^�k�7�P�đ}�t���GҸ�]R�nj��lu{B�����j�g�zL�����n�l��X+�O�z�Z�!��@�`�[θ@P]����K�O0o�QÑ,�bS�	VlW;���n���Du��1��h�32��Yj*�0�闥�S�*�����3l�7v�	���&0B���,�܎�)��au��2+�ub�;P�3׳��v���E��	����)z�����Hu~U�}CP�f�u������f��u�q�Vt����ݎh�Kub�<�$�YB��
���s��=O"x��y��U!{j�;2�NK#[��f�yu�Mͷ9�u�D�K�;{�b'�5��^7x#j;�$1�V�=��H̭���U�K����#��G�k6N1&�m�����p�t�g5`����3��
�����R�uƜ��8�zr�׆������.@�ɌiZ��2������ԉ��1��.�:�s�w'uX�{���jd�'�����_
�G���lB����'�{��k���P�p������9?t:6�ύ�RXW��7QER�Vc<�)�p�7�����} !Y����c*���y��	�8�V�W�?�i�_,|$�M�����ɤ6]Rȶwd7nqcΌ}/%�+���2�p�}յ����2Q��:��B�Ƅę����Rۦ��.+m��DY�ˊh�Kb�a۫9D`f]^��6��pB>ʙ���3A�p���<��~�<mZ�z���꾗{���EK����%g��~�\�ԷΞRy,T`�"�-B�v�p�7��'�{����@���O_�m�����|�g��1|�@Ĭ�u�;�22x����M�����30�Y�
�:�����+'�M��/��U^m�����o�_�s���5��C�ߩ
�i�o&��'=�H~��S�J�d��R<d��{��m��&����8�f�k����Vq���d*)�f���g�����>'���gb�M�U�+�gsܷ�O�>F��S%�Y�GE�!�t�A�J���CU�n<�V|uӗ��S0,<�@i����=�{Y"�=PWTB�3mu���ks�0�s�\�_Y��WG�J�۶�V]	�t�.����� Uȼ�ҭ��o�z'J��Z\�j�H>�N��wmF9X	/�ҷl�6�,����i1��
j��Z�}ASs�Sl<yH���&(����Whf��W�W#}yQ�J!1�wzHO���x�`���-Wh`!|�k�*��7�@���U��C[[2��Ҷt�����%Hw/i#���B!5��9|�Y(��Ǣ,d��l���-�\�E��+n�\7������ek��L;�P.-�:�����6��LHS4(��5a��V��r,|�g��*�l1������C���3��'�X[����ʵɮܬ�����Z#��k��>�c��A���:�Cp��'x��X1CnVKv�Yr�f�"d(Pj�F�l��2&n���}آ�z�ݤ��w>Ê�u�Ȭ)u�u�;�U�c�.��������A�u����z�Ӭ|uMUu��b���VE(� �s;G� ��-��6Z*�t¸P�Z:�q988$���(]����]^C�]<��7sEj��E˶T�P��u����B�!R�l9y�,զ�EV5׵��p�&%�,L��X�n[+�z��،jV��yo��J�ήAh��۾��刌Ju�:�<���_^�-9ie��o��<쎠R���Tyxp%���񬨆�"��R��9�m�3�Kb�k�'M�A)���rXc5h[/J�{��K���9#���k�9������zQ�nV��w�M`�Y�:����X�z�9lQ�6�yvUˣ��r��醃%�G�����z��pG�n�u�y�+2���u�2GF�šu-6�M��e��b�du��Z*X5��s=q���r�j��4Y���L���:n�p�|��uN|z\�Ÿ�;^�j(M筳%��Y�������U5�	�n����5���x
&#�pve�Ƌ淖��� Nb��Bƚ�\5P�e˨4c�u�T=9�1sb�e&ۺ�3��䦛VU��EJ����=CscF�݁��6��5�����+�4�*H�L;FuHۆfI�ya ��"�qb#~���ʝ+.H�7�Ar�~���g���V��QY\볫4b�9`�����Cz�v��\��8� ���ٔ�[ic�Y>R��[:�7��kԨV'�A�X"�e��S ������j��r�����\Cpʉ�}G�[�z�� �a�.`o3�+�}A��`���K�x�m��7���4[�8��438S�; �t5&T6��2�P�vs�y�F�x�q*(�iq.�n����P�E�"w I�]���DZEo
Lv��Y�\YђL�˷��S�V�e�t��"��G{��6�9}*5�{r닩�t�a��[ϢS��3y��ۗ��q4y"�qյ&�V>��}��1���,���"��lDQAJ�īDQ�#�,`��h��#"�"0(,U�Z�
�cEb���,X�"�A�2fY����J�Q�X�1�TE��b(��
�eƨ*�aT��j%�[Q2�DA�W(�F0E��QƢ��E)DD�X)l�q�*(�+��*EQS)A�fQd�`���QT�0�TUDQC,���R�֢�1X�X��
e(���-��.61Ī�
�ŋ�������)m�n6V ��U�e�*#R��1�iS-C,�Ub*���1X[La�0P Q#�[��lx����Vl+���5��K�E@[�:ۓ$Y��L�٠����Z��I�l�Ӛ�=�FoG$�	���G��F^⥩E��G,��'�q!�g%@Qa�����O��&$�������~�1?M��!�����톙�%g�7�ö�Y��u��� ����i:Π����2z� �}������&��ϼ��o�1��QH/�����v�!��p�$�b���
������sL�Y1E7�?!�s�&!���$���'���l=aXx�Ʃ��2T��γH���`O�ƨ�j����-���p�+�E��
퓼�<}`V��>�w'��� ��y'��i���1�I�$״���Ă��U�h/�4���oT?&����x�"����u?]���d�K���9��w��)�O82�4�b9Ci�q���3Y�ONy�y=d�=B���C�m����ߵ�R|����Y�%q��Ky�1��+�{f�H������2|g����yS=]�}q��Ψ#�1��l�+��1�ϝy�Cl��!�,�����v��>���&�Xzs]�6�OY1'���2m�c��;��aP����+=d��z��}דK6�����Ί=����=>S�QCLZ�^�܁S���ߖq�v�Y���N��q�Ϯ3L8���c̰1�N��s8°>k'g{�w<f��b��<B���LN^��Y�ڳ|#/D��j_�*�W�Uj�!�Xi��+�K�|Ԩ�d٭d?2���J��}�i&ЯP����3��k�N�]$����Ne��E�d��O\IϏotH/�����s�;���_w7��yz���`xצ��~M���C����T��8���I�+'���i��J�C�13VJ�6�Fq��(��Mӻ���'�Q8��c�f�l1:��n�ys��d\�Wo	<C��{�B�)�������h��d��w�B��H/��{�ߖ�f�q�q!�gS��iE ����CL�8�!��1��bu�M�HJ�����1E5������}x{߯�}��;+_S�Laз�*I^���y���Ì*a�;�!��%gs���QH,���CH�X�ӽ�OX1�Aq��Y��Ă�|�0>M����j�3L<La��7��޿>����Ck��6�vG_^����*zc�������[�Mb�g��ҫ���?B�Ǚ�v�c����j��6B���gV��wt/��Rz����0��:��$����܉�2�w ��!y{��L'��ڷ&��n�Q�=�W�D{ވ����t�>���Lzd�1?�_�+�Y�c;�&2~=��OP���'���
��WN�����VN����P+:���X~eU@�]��os��$�+����\�>��Pg�4��.�{5sj�G�~�:�ɴ��f錬������`c6��oT�(m ����a��1����gS����&�@�+16g>�ᤝB�y3�M?����8��s�j�f�(��s^i�w�y��;~��o�IPY��]d>ݟ�*M��a�����+�t�2w�L����W����G��i&�Ǭ:��A},8�f��}̅t����<�b"f&}I��8������X�f�c5���fءY����;a�1>g�3���5����11�& )�����|N2c<ݟ���W���0�*!��_�
�2W�m�uE ��FɈ��-I����;ݕ޼��:_�~�s'���������DTAU���
��A{�0�<f�TP�Y�?&0��ᙓI�O����
��*zk2����1���I���C��m'�*N���g_�1��Ve���~�<���׹���}o]4�Β�Vi��0��d���L�%I�W�������t�Cý�o�&�n�x����2��VڤbO�'�;��Ci�&k!U��M��:��O�=�����)J�M�n-c��U@PT���8�I<B���x�<b��Cl�9M�6�u���O̕E�9�u'�,�%I�|��~dӎ�=����*m�[�|큌���3w0ԩ��sO�y��ʸ�����Nۦ�T��� ,��������O��=jCV�;�f3H
,��f3�P������ވ.�|�'�s'�6��;�N>�b�ߵ�a��q4ɛ���6�$���f����*]��yϣ��	�S���HVq��T�6§��]��ɴP���J�`T�8�Rq�8�����0�*)��3L8��r��H/�<��u<E���_�����~�w����o��i���d�t�2E%B�<�����
���i��|¸��ۤ��k�L:ʊ���8�g��&3s˧��Lx������N�M!�)1�2w,����|��m���)����;�f;�I��.���.NYBA�voQ��-�H��-3)��M���svpY��Ѝ�<�%$5�R��X��mv_q�T�ǵ���3�6:�7kY���U���`>/�eK���L��q��˥�=��V��	��銅T��{�����������&=�$�w��N�C���&Օ=a�;�t��Y�<OKܛH(M����|�q
�ڡ�i�8��d4��Y����q��bq�����}�螵j����<������
}�4�:Z�l*z��=�׉�2W���Rz�$z��W�LE��ɧ��{C�w<`u�-<��J6�Xm�f��Y�q��H.�|�HO}�������z����g!���;��M�|��|��}���}��	=`k�y��_XO��rɶO�P����4_r̇ɹ��PY<g7���g��7��~�/�?o���z�ٌ����6û�Y�LM�g��������mq�@ߗ�L�����~�h���+;�oړi8�I��A�?�1�����6���T
�w�u�l1�Vo}�߽���e�u�[�����޵��V~d�3�y���'�ǈ���a|�q:� �L���ϙ��͡������hbC���Ua��15�'��:��N��ڇ���'��1'P�hw�_N�~���v�T��O`\��YC}��>A����C��~'�@�Vq�Nf�u��~�Y�'�g+�n�C�O�<g���a�
�Cf�׏��$�[�̞&$���&ް�b(~7I��������a�p���	y�O�����+����}��	R<;̓L�����3:�$��6]��Ϙcm|�r���Lg�Ȱ���3s��I�T?0��/X�����]yHVz���{�y������t�o�פ��2k,��ri�d���<5�ki����u? �$�:���CL�&0�}�ɤ���I�=z�$i����Ax°�4�&�YΟ�
��+�DfwC�����^~N?�oO̞$���Ρ���0���1���Y79�5�4�Xu�{l6�gY*�Xm�2m1�O�̚a�VO������Ͳs)�u���H,�ٚ�6jc�h�������#l���h_Ѻ�	]�.g޹ٷ�
�?;C��@��%c�0���
%N=dĞ'��M2�b���9���Ƴ�w$��2T��wL��I��O9���!SL����i*�c��"�W��.����ǔl���r ��k�� �F˾���v9����VGD�;w���V��}M�R'_�����::��@�f�Mښ'V�U&e�����8��h%_oԝ�X����\j��}:��ax�	N$���Y��oS��VEx�dr��{!	
�V?z"=�*���[r��$m�f>�_)Rl�a�b)�|`]X~�u�0=j���Ae@S�H,�+=��<Ci�湠��a�y��
~tɓ����P����f}�T�Ϣ�#���{5�M$�
�����ӟX��<5t��8��B����i�0��C��&3�%E;?S$��k��.$�>q?��L:��G<��H,�&(�}�K�9�b[h��.�2vb*c�.w�x�At³���z�L���x^`mE'���4��ɉ=B�k�ACO_�������'��3�Jì�������Sg�6���q1����;��]�;a]v��C�@�Vq��<�~awd�w��]$x�������QH)�s��'�I=�a�;a��Xc�l��lZ�į�w� (����u6�~��L�2�b���>��DT��즪;��W�$n�2��>d�vv�"β{�z����I<B�Y9˧�
�l*}u��㴂�S���}d�J��ٌ�����bzw �0.���'��ư��6��LDsk��f��vL�t.�Z\LǢfm��q�CI��:�����$��<t�S�<�f�Xu�w?w�8��N!P��la�szȡ�x遳�޶�2Vc
���g̕�>�w��^����^lߺ��s���B�ĝ5f��x��:é�R4é���N3H�Tזq6��b�]��1�
��d�&�>eg?O�;�<@QI���g=�bN3��3i8�z���Z�����3�gKrz���C����4βV'���U�Ĭ�'�Ri
퓉����0����~��̜�'�CV�$ۉ9��Ϲ�k�Vy~���@��))��:c�%6DA��~�����՗UV���$�6ϓL1'7�P�&2�b����C�1���٦z�Fq���I��l��8�2�I�*|��O��y��3��
y��ɧ�K�+!����V�p��Ͻ>�����4��<Ф��߹����?0:�zY<՞�����R8�=�s3�uH.y�!������-H)��='�@Qa�5�}N2bOR���º�;�v�-wwJk�*DP��++L��;ގ��{ۡ6���v�KV�}õf*N٤�~�L�L����w��B=r�B�[�:�6n��vt��S�v9���Tۨ{I5 b�=�˳���A��,��Ҳ��`O��e�\pL�nd�����}��_W�o~��W���3�T�u���9~a�8Î{d�y��>d��M�s���2T��u�����O��m?3\gy?fu�Af0�g��C�m�˾�u6�ǨbAt��b�<���}����;��{��<���|`V�c+���&�P���LI��u
�����3�aX~C�'��gY+�ﺛEY1+8�>�M��qi��gX��^Y���SĂͦs���=�w�o�z��y�ض�{���9��m��bVT�q��1�Z�U��|Cl5&��q4Χ�1_֠i+8�a��,1�l�Y��O�d�fa���J3�</3H
,��e)����{���}��f}���?2u'�T�P��)
�i�[ɴ����$?L޵<d��K����+?2W�k�g��Oɚ��u�`m����Y�V?XTR8���Z�0������gu:U�k7����������14�0Ƿ0��S珓>։��9f�S����xky�=a^��1?M��!�������L������;i�ɯu��� ���d�u�Aq'��>ϵ^o��|���k��7�=~H,��
��*)���6���4���<�0�$�b��3�=k'��{�e�Ɉ
)���3�Y1'�1'P�_�>7�Oz°���T�
�*}���o9��o�}�6{���[�f��*��+4�0ĚB�2t������������$>�$�VM5����x�C��xgp�A}@��y��.!�Z������i*(J�'P�9�x}�?g�w��������*OP��e~{�bM=C��P�c:�F~C��� (�������
����w'��
�Ӿd4������}³�J�%��c?2W���Oh���xw�?{_;k}�����������٦w��C�gU%|�d�R8���4�ߘ|�2~����N��<;v��5>��q��s]�6�OY1'�ܳHz��t��~�P�
�0��l����ޟv�O*��NMocT����)���L}��x���>a�`��ص ������Aq�3�㤂�g���m�YQ`o��&0���k i�'Y�xs��XV����So��& /�~~ŜB���U�!�ml���&�um���XV8��c:���'u�0_p�IEl�}����gr���p��j^=5��A���wФ�Ò!��n5Ո<Eeŵ;j^rz�(&���M��j�N%0{4�9�%5����@b��Њ1�[�f���9�-�16ѶK���c&
���!'o�u�i�/Z�r�12���z=�DD�֍5	��5V\���O����v�P�OP�Ϭ����
��m>jT
�2zkY̨�'�a��M$��g�`V�O)�Y:�t�_>�<d�Y8�Y�J�$�Ĝ��3�\��y|�f��x�]�w�ޖ>��5�l�&���1��"�R��q��N!Y6���i��J�C�1?nɷL�E�O5���Y��ug*M��
q�SR��|�lU�Ӯr�}��&Tvo]?0�>d���N�;��u��d�r���|�]���P��R�<�p��é�i'�皝|He�J��] (���g�P�<g�4��a��g`��Dd���5��?}�z2��@��|�d�
)�|����ö��Cԕ�l�y���Ì*a�?�i�d�߹�P���|�?sh�X�A�᧬
�Π���3��1��2!L\�:|&&c�wڀǘj�1|!�}������ǝ���m���v�|�q��?o=aXjg�ǉ�Ld����
�n��8O��:�t�}�@x������A��T
ΰ�Ұ�d�_�5��M��+��|����5�������߮~��>����ǽ��l�� y�c+'�d���?Xͤ��5Nv���OLV|C�@�Vu<a���0�EĬ�ٜ����u
��g�*!��}}����g��~���N�o�/���Y�w����
,�7u��vu���k��z��Ǭ
��O;˦z�YY+�S_�R?$�n=a��R���u�C�XW�us���|��������[�����k�z��E��^efءY��M�X���1=g��wP�Ʋx]d���L@R��+
�8Ɍ��C���=��
¡�����+4�]���N�Ag���wO/���(��w�����C;�~��(
�> �s�1�O��u�z�LH/��0�<a�TP�ZE���c^�fd�Av���Az z�<5�YY�l���و��
�~���I�'�F��C��_OW�>�϶}'�g�'�Shu�T
�3g?`m�QVM���c%I�W\���y�B���s��ɤۤ��g���O��T��I���}�������Ұ����.}f	�#b��PY��v��J�ض��޾w+����Ç*<w�J��QV�nN�RM�\���xʐ��f��P�f�?�R�k�'��7g�]�8�.Y���Kc��[j6J���G��G�Y��}��3��w�8�����@Q@ĩ���:�i>B��{O���^!�xr�`m��%�nO*�?s��O�Y�J����A������<����*m�[�|;`c>d�����)�k;�k�]�~�n�o[�A�� ��wT4�a��X�������4���֤7l���f�Y?2��P���!��������ﹹ��Zì*~}d�����x}D!L}����k��f����{��q��>q�t�rM��
���y��~��0�5M3l*yi٪~d�(q�P��	_�
�g]$�8�s���0�*)��f�q��E�6\��D�L{RLN�Z�ou�c�6��°>{��Rz�ϵd�y߲E%B�<��~�<I�&'�)���a�
�j����T
���L:ʪ�g��i��T���t�0ǌ9 D�=��1P�)|S��w��]�Z�+<d�Y;�����Y�O��7Rg�1 ����M+_�c�� bV~O��{�h
(M��jm>a�8�f!�c�)+�=7�Cl��a�0g*�w�:��e<�Xw������/�:c'?Y�Jγhbu��;H�Xi�N�s����>d���uS�R=L���q1M�Y4���a�8�n�jCv�gy��@Qa��f��Y�q�:�~��7ϛ���Ͼ��}��~�N����_�6�{�8ΰ��g����xɌ<eE�XW��Zi'�T=I_�܁�=�s�?>���妧æIJW��R�d����8r��F���a�p9�")��Pm�)^��ҙ�t�ƞ������2����]���St�����Yg�"yo��_-_;�L\�±]��A}~�5g4�­��洫�6�,l�!r"Q��v&�C��B�gh9��:�q�j�B>ֳ�s�ܪ��b�ڻ��XF�Y�bkэ/c�d��8�&_YW4T�
5��A��i�<����w�P�~�x��2V_�;�i^�=W:u<|���9�����n�3��^�"� :���es�㙷�@��] ��mU�:�bT5�ވ�DDc�Yؕ�8{R����0�D�۩�F b�s���u�_��u���1�ۋڻ�܈G�w,h"�kMe���;)�a��,=ȺaT1^�}5�,E�0�`2�7!�����/��d*Р�L��ԞT�vzAbL$D���;.pU]��Q��������.�1��L�ҫs6�o�Ȃ��v41{��x���:�đ��HbuA�sZn�������n�Y@����V6D����6���u
_F�Q;��������p��kq�{��_%,5�3v�>�Ҩ�� �rRY�ħ�	��ά��}�=�E/�v#��/ϊ������W�,�� �hy������}J׬���"�P��.8���Ω����?Wf��{��E�ϛ6p��l�WD#���w��N��Uʆ�⩇�rTP7ظ�{g6D��:K�ێr��&{�M#�VvD�n�F�>魉W֦�屷Ov�X�w9\K�8����l�1
�5\p>rq�j]*z5x�b|���&��ӄ���q���p܇�p�I/�䞌
�oQp�\���F�".doV�r<� l��f��?	Z+�=��{�U�VL�v����>j�w����N�8P4*�NR�msޛ٨[Ý%���C��䡚;��YSt;7�1�Rk�rugp�Swt�=��gvu8p]�`ُ�EC[f��-B��؅6��J�pN��-�8dT�}S�
-N#=A�&�I��R����*�T��ў8���b*`Ń�1�Ҙa�6@���f��=]�gF������9�"\\@���\ ��΍1�[�0�ܪ7����n*�/�ogaA���;L�[=W���LF���s�u�'�j���� h1����xF�g�-F�c��_+���cXHt��u�ri36�dL;�3����.��>�4�v�ek�l=7��uuv4,�񃂩��c㒁���Ӆ��EK��	W��q�ɕ{��(��c��ֶŒ{��70�Bl$.0L���58��銔�\��nE��T��0�Y=]:�GL�ԯ���(]zt8���)g�e3����ڴ�����(��������q��R�f�	�Cn�E!� ��~��|�cn(���*�W|�XYk�]B�̗��{�pƓ�ɹ�d?��C����=���?�j�}؉� 0f!��F�C*��f+�sE[~��a^���ڮ4����#gN�&M��<2�z#X���,
dLq �kѺB�H���ƾ�e��G��\���G�{)s:ࠝ���U԰���|�w^m��Oy�u�w�#`���Y��ջm��<� ��u+��=G�n!�<`����(��W�z=�Dz���#�O8�?yt�FQ������uce�)��%l��X)�>�p:��u/.��ׯu{���n�����[�zn]觢�Ә���n�ry==,u���1Ӳd�Y)��h�\r���.�V��[����MꃨX��ø^��&++���>R��o=�)�<:-�Toڧ����yh���΅`�u;�����R�B��-:r�����Os0t����5��c��dc���: �꬟)5�X�R�W��uh���v<��ׁoE��[���'ه�M;�GG5@_J�I����"�qK��.{7b�C�=�=K25�\ED�e�]s���˛�:c�P��l۪�E�./��9�E �k��]C:���5��ۆM�S3�=�;�����==C��.o��c�1��Ð�lus���'�)����Ϩ����{�T=�UN.����=��M`�.<�~ɢW�� ��>�=�y�����ۇ(�z��e�&5�V��.��� 5��|=fo*�L9��V�]�L�70�'�D)Hۆ♸i�c-���|����̓+L�{qJF���4;��I}A]+�Z.�������!�+i�9�7�V��y�|.^w[�8�B]��$� ]�D8S���\]�.h��,��u�P��7��a*ɍ>HU�\�D�+0�CjoVl'��\����hw���01�՝ܺ�̗R+�u6�T���k��Fh�h=q0��ih����Vq��N�6���yε'P��In��`�N��:��sjY[����s����,�s��7�L�b�b���ƗW*�g���Í]��YILl!��m��D�w��˞l�����>a������5SX� ��t��r�9]ˍ<�d�O�]�F]v�L�O�N����]U��]:M�kg��$1۳ϭr.fw[��p_\���1|���M��a�p ˫��a�]�� ���\s�������9�n�S���TmP�gV3����ҩ;�A�)q�ZkBK��Gwٴ�� 4mVj+3V���zٜ;�4�Z{�w@YZ.�!��v "ux��r� �X.�9Aev��%a��w��t���3��ă}�5ӝ�ծ�ӳKJwt* �7�� � �p::�R\�R<'x*9�<���f��u��C�v���4�!�
��^Qτ���ci����ʎk6A�ZM�#x.\��d F6���|E�������ᅑX��[SZ$�r�#g�4/6�$xSH���.�r
F�i*�az��y��ks*����m�6n#N\���i��8բ����;����E��S\n��M(]4�s�A�5���\$u��A�h��O=���!��A��č��3+on+��V���6�^L�	{pA��`�ǥ\!l���\+v=v�6T�rUtFv����ʟk`1�U]�
y0�8���Ն���dj�vԶ����;��T���?\�O�X� �2.�k�t�Vu�ů�7�j&,iVB����ݡ|����|)��1���[%>Z�a�K��:�(:�������ܺ��^�I�7�gQ��,�f��֐�8�|�&��q��MVy#!H&pa���ݪ����~�÷���\6����ug �w�-�//<�RtMAZ]�LpU+/1�k��	�0l2A��'-:�w���u���n.��`j@�whm[��ݛd�]�����B��:v��R0 �c6I��/�C�CT��F`Ր%����ܪ�_R��e�1��s%���t4�B�ﲘ��2	w�:޵@,��8�Ţ`��#P+M�2C��T��Vj�b�m�J1�[tq�b�i�D[,p�{P4�+��7�Yt%q�~G�xv1E�u`3�5��Nѭ7�Q ��P�/8��]WzlY�S���E��G\Л;�\�Eb'M�D�Z���m)���m����Ϗ�*���#\AVV�)�&8�m���+��1�����4q��
6�ĕ#ip���0D�Q3.��J��P�Th[U���b�r�-2�YDAU�*�aXҕ�V%�+b�+K1�aU���U
V�Ĳ��H���FثB����V���bU����Q1
�kFةR��[J(ZZȖUYZ"�ZB�[F�h�RUFEX ����Ad-�֕DD��m��U��婕aR��R�D�B��PkFШ�j&8��aX��VԱ�V����#,ER�[UQ���UKAkYm���Җ$�H1"0�s)�5�¨����Q�V�J�X�V*0PR�,�XQ[lQk�����e�fk�ԗj'��	)oWjz��o��@wnh�s��� ՋYՁ�C	��56_ʏ3{f�HPO��G���)l6݌�7v)�ӛ{��<)�<>�>S��>��r�@�j�[���mȤ��f�v�UW]\�N6���T���I���pT��q�E,�MA��X5}|�!��a����û�
Ƨ
�({�ޝ�1��w�F*}|������׆�aB��SԽ��p�G�ޙ��K�l���.|yP�4������jw����ϫ_�^Kj�\�����qT��_���O�VN��Q�&\��b�����?y�x6{�L�'N�����&_M��?|j�Z��4l?r��9�򾫅S��6)�;~��Ć߯�v̊܊�q�6k����I�==q�����Z�]A�6=ҕ��`^>��U���&�gS
c�v�?3�;���:g�P��e�h�
���堺��x?S��8�����%�oPȎȦkU)84Ϯ�#DnB���D��o��rzxZjP����7"��W�g)^�3/���|㵜�Յ ?|���S}�ٍ����U�1dK�72�W�M��gi��Ҍ��FTttv��Բՠ���d����\�{b��Y<fm�6��|����԰�t��p��\�I�8s��:��Nk�5��ʈX&i��k'!y��o�V.˧̯�G��ζ�gV��ښ6c�����U�}U�<Q'����VVvQ��m[�&a�r�OJ�c��I���.D�0�z�����6z�o�y�����
;Ep7���S�{[)姞SO�OK�pV`.v4���Y���J�� L��\D�OJ�2¡R[��t>���)��0�\��J��>4ȣ{�^tE>ݴa��0����yW�+5��
~�����5*��Х��<���<����m""�Ri�k\΃�n�'��G]�K��>1�h�{�Lj�\�|�Y��]&�Oh]&\=��~�eI�*�t�Ûr.��Th+b�(ĬƓ�[�f���x��OfWx�˝��R"/�ԜX\�D�BL$D���˝�n����S�� 0PrN@r=[5*'�]ާKh�;����" t�K�K���i�����b8 �.f*St��I�u��u���pbEN�bx��kd@��N��L1�)}���oGEgt���0�vt��779,��Gz/�/uQ|��1,�b<Sƥ�ά�({�9��ޭ�ue�)�V؈:�+*V�&�<t#� �,<��إ4p�-�o��~|�e��n���;�ѱ�:��5����6n��a�{�����p�W���1Du��P�8�QF��o'�/�FA4�۰nc���XVr��D{�wٚ�v�׶���W������2{`��+�Y�a�;�x�t6\�{ĉ��wfdָ�PfܸF�B�tj��!{>l��6��byMJ���)z��
��'-}�4�����trn��I�U
Lp���u\���	��K[Q�
���H�q.c���'�Eb��U��d��iNC��E��#�D�����]{U��8�*S(��r�S�������dl�R̰�xr�Lf�5�ܣ��/�_	�x�~5��M�ʠ��o�K�wZ������8��g���j��y}CH>=>��u~��|�S
�hv��/��e���=]/�؍*�"\X�V
�>G��б��yf��a7��%�ʮ�T�&˭�V��N��\����BY����!�s�G�Е�.Q��s-v=d�q��LB��`*l_�cr���&c�۬��x�
�0����Wc��7ot�jemgq��D��8H������dK�{���T�>O��L��q�G�{�=�j��{�m$`��*�w�yh�Yf�FXc��h���\�V��/��y�U����f����YYfYs�٬��mS�n6���E��A�a������i���-�&���Ogs��7����'����oj����1�Z�ٔ�on��H��fI�v8�`�-���ncm]*�m���iu���O�+:���U�U}۞�����E���
�Z"q�@���5'������Jarr�)�wL+��Yg��B�]`�0�O���Q[NORo=��f%Y�s��^�+��;����&G��߱�������eVyLI�zA߬
�=�2^��hb�ٳ��Wկx���:|-���.��y�0f*-m���퉊q�R�Q�1P$,[��[�k�ʵ ;=��ن������1����
��ˑ;��FD³.��������U��w#�tZ|%n�a�f��c�9M����U>�{Ss�H�ϻ+���jw��U��\�uu/f彮��%U�{���Љ
�<�.ϕ���1��D�����7>IW�ʟ^�����i�nё��e�&r�<����9h��S�H��=ƎO70}��r���F��
3�����`��ǫ�>�\��j�k�����4�}���ǡ������W�Ʌ�.������$���.�p�x#	:��M��~fsTd������j
�M}�sdhZwW|�+~�^Py}�[
�r���\������씹a�:�rʠ8�:�G��Ԇ��qV�d��۷S��e��\b��HZD��ʎ,��\ܫ��R0u�Q�5$��h�ƫ�DDz#���yK�����A͐�RaJ��Lt���}��uW�%��b�b�!�D���c�D�	�����n��L��j��;;)߭�OPMS���f{j2&��!��g�<�t�Gi�z��Ub��i^�p����cz�[��΄���|�g\�^o��e����^w���|6C�N�a�]V+dd�|�J��Cb�˲�y�J�����`��M���y��Oju}GKU�"N�"������,|~y���tf�O����PU�����x;�ڤR��c�%,+�!�9�5:�:>1.LHC���A�	�#|*�N6�v;������QT���c�}��q��-S
�DtMGu	n�:�"-;�3
`���ŗP�'hl� ��}��s�'!E.�b�G%h\*w�A�;N}Q݊̉���ԘnʣV�e�Ձv�ѡg&J�-f�H�[)�����p�،���n�N�8�o�L�)�O�.yfm��rd�rjK�8��]� �̩Xשr���j��to�*F��+���Y_+=Cnc��o��;�^m�FZ�}�vT��+)#��k�ʣϻV����4S�+d�ak�}[�\�Ύ	��$b��ήc�<�VZؕ�-;���qf��t%�[3�e(�v�v����̽�*m����2�<��@�ȫO����Ս�T���궶��u��Nӛ�.�v����}���Uv�Q�S�UBu ��� ����`�`�x6�& �J�I����PH\M0��#a��s-gc�-w������P��"̳����t�ř��ϫ�V�4/���X�]5`ΩSVu8b�0�>��8�n'ҵ�V3<�)���I�C��4�*�!0���ܧ��}5��6��AH��H��~����}��f7<�0��F,�nni�&N蓏���k�Z���~`TKu��H6#�6!λ@����%��z�{�l\�X���v��G�9}y1Q-�<X�8�x��M����1w�)>����֞yM_�:$�"�=��0�G �G �IПo� ���z�'��ū������]J�tK�AK��k���4�
��KH��!���XDJ�+�`����N�����Vi{��s���r��r�K�9�D�3˩p�����Χ�pm\O�u1(��G]�K���ga6�����X �������ǃ������:0�^�c�U
����E�V`�x0]���g	��E�E�����b�^E:Q!�е��i��<���n�ǧ\}Փ�cJf�����d+�>�ʛ[��Ky�ȷ8�r��LuӃ�3�(�gVN��e��,B��0{14^�qp�嵌9]W��7���ҹٸGB��;V8������R�[g����nP ���U`�=�{�/�).`���7�f�q"s�ԩ��������y�
�=��!V�uȧc����Ļ��=C+x"v��	ǸKo��)mb妋�t�f�s�gxUyI`������	�����P��+�� ��x��,����E{G����m�:����83�ӓ䳍��xo�PW]�e�y1�o��o�75k;G,�R¾�	]�0���i��45�ϴ�]N��e<v�	�
�O:�=�[L�SibS��&\3M��emT]�.�}m�^��b:`Y��}56�O��#���9ޛ��'w�!�ur��)p�B����V�V�'"x��7#ʶrKu�p���&m�`e��	ln���g���*E⇔MA�0
�m
�r� |��c�jq��禘�q���-+�L�="zo��LN����	]�,U��6p���;&��%]ؔ���������r�c.��Ҵ6Y�*"zi	�
Vϗ�t4��̡�W�J���V �R��Ϊ���>��t�3뭱�Rĳ�����h��8�2�8j�
�A��\C,)�Y�y�kn�Z#7^�����h�
fu�#7���²FQ'k.�$�h�c���,����DpN�X ��݁�oZ�	��K�Z���l�o{��ݹ�3ʬч��ܯ���S�ĩRr��>aL3᧦������ʡm����#x�e`���J,kQi�8���U��Tu�`56��r��ή��*�]Zw�'^�[��xDI��>bs-qx.�o,+�HN5FE��ʄs$j.n;��̋F��:���D���p@W��@�tX�`[]�&���0�"pC8H��ǲvU���^\G;S�g��rC��*�1/�of�R*� ��}����t�)c�M�x� Q����X"�;�n�x�Yr��tm���ι�
��ۗ^��[c�E,����Y�s��]�`�x�;�MU��ھq0�ܴQ!�W���{Q>�����H�@�����}u�g�X�����7>T���Δ6�O3�s>1��r�rpC�'gLK���2�ޗ��wu׈KZu��w����3�n�MNI�U�4c��1��țI�dd���U�P����X(r/���^v�[䫆8�w:E�a�PgX٩}��Ɯ�ߺ��Э�NNr}jZ��5]�ht����nͧJ���"��6<3jt�B��n����=Ʀ����5P�idOg&��+p=٫ה�1� ��jZ��g���fnS�	Nh�^gP���	�zyo_RR�:�Ű��<�iړ��e�����3�
Xgn��l.u��ы;@A���-���P���"�}9�C��iic�mY��+t�/Oo�c�Iw+FD�9��MQź�Y��F�6�S�89thlr�XM*ut������s(J��� t[>~2�^��9Ya���sp�/Dg����|�ۀy�c@Lp�Z��<8̫z<�sWh�&�m�wÂK1r�UǶ]�-��%�Ql)�h�.���q<T�1�6�W0�������FY�O�m)* CAI�����.n!��1����6Z�D�!����輺�9Z�y;]f�NPW�Ң��7����3�zUOM�����];0��Q�#j0�է�0�V�2���6$�v���e�^
 �|�?�:��Py�L�|�T�[�=�(�+K��n*/*�|��-�fvT����By����·<��B�
���Uw@��<;A]�@�'n^��Kˡ>թѱ� ��V�*ssSǖ�MiRn;��V�>�4��Ŋ�V����;y�i��7)��K�+��s�!�TkT�.p|Fq�)`�m�c�� �|���`�1ŗ�+id&9B.yoZ�[�4�r�>'���єrU�]�m�f�ngM�=�t����wY�	b>�s{�:A��I�)u7V��o�p�Zx�{�ϋYd-�����z�+sX�D�����}������{���*��&���s��S�"MDwP�������f7ЄP�ܓ����������]��;�x�Y�l�L<�[��w
�����w�v��^�op�{	i�<:7���V�i��O�uZ�Mc5���
���g"��]h�r|�d��yf`��T�[x�;�ݎH���a-C���j��uF��yV�;~�+�Ce�:zMJ���<��x#�ر�W{)�{&�lמ;�hsѲ������_��u�6=ґ�g�1Ӛk9�+x�����&���ԟs��u�<����'����r�zr�Y�1����7 �g�^��N��^ٽ��6�Զ�Icbg�n�����r�ޝ���χ'����|Up�wt�Y�츛�U)�s��t�F�w�����1������q*��b�h]�1K���.��vwk%K�{� ��Vz���nc���]�zzV@t�}��kxr�.��e�V�q��s�dJ�S
�y�R��N�PL�B���Τ�:�0䦢����D.qӬ�Q�F�u�*��ˈ�=[����ܢ��qD�j�2�U���j[b���:C+u⣻|1�{�ۣa���4����ۘr��Ϋ�QJ�;$�U�:��o_c�:�F�-���c�ӭ��[5f��ğ��\�Of��t9[��뗹V�&�L��Ā�;T�Uً[1�0JSN�|8	�ϳ^� {-[ˉd��j֔�Z��H2�ܦR�'<�o�Ze�w�h����#�.�GxK����4��ڦk�b1�e�]δF�Y�q����;kuh�vF��9\�Tw&��L"�PŇq�&���vN4�!t���[iF�B�5�U�5�Q� L���$(y�����ꛕ?!W�]����]w�԰�Q;�1X6u������[R��3\�u�X��ގ9b}n����=�mO�&�A���A�D�gCM��=3�kTRQ�*�����|{�g7¡���n�Ǜ@]�;�ZȷA�/�C�z[�`W���J��a�gl�Tte��[}I�W.
��r�k�r!��扵�Od�K_!6 cae�(�i�}q���s{/{g>bs1�z�[����mA����p�b�-�7èbt�����'�P�4&�i�L';.-�|B�u&�捠���tmV�μ�+�cymc�*����0������.#\�q��K8ɾ���e.s����w�o\/u����s�/�g6�������٤{�v�MH�[\��*�h	��bv_.��;��x�EX�X�:���d:ܼ�Wb���ʃ&�䲱6�d��$Δ(u���7rm��{������M�2�P��� ͒��S�Y7b�1��m�[K�<غ�T��!ˍ���oi��=�D�.��]���q��nn�P�ʡ���k�"�'w��4�T윗ki^8��ۛy���~�C��O4�t@�ILv׸.+J$Ft�P!l�ySt3�e[(CKMmJ����,���C��ֆ����Q��n�V�)z;�|y*--/�����t��Ɣ��y��W)�Ѻ��+"}��p��*�h�+�]-��唂�B��J�r��NխZ.��I���\����\�e,���(w���J�G/+����S@��)ي�!ӨިTn�}0�٭�e�m]�h��ڧc3vS#_%w0�<��Yl��y��FT���*��G�B2�3 ���Viv�[SD+�h�2����Q����r	��^\I���m���SB2E1⥮�������K�Ii�:b�r�����QK�v�i����6�ˌA���|(�V���qm�3A�`;�#u��3t�!�������ig3�>v��:��;:�_ ��nu�*�A�������Q[l��m
�+h]Xc�T��E)mTX-Kl�Z���b`�,�*Q(��E�+�e���kQ�0+Ym��[T��-��J��մl-�Q�
�P��[aXj�b-j6YQj���X�b�R�E��-h)Zԕ+U����V��Fڅ`�V-�
��h����YX(�aZ��R9�b������X
c*L��ihUKl�h�-�6�J�1(�Z�X�*R�F���E��*V�l�k[Q�VڡX����"1mE��
�(��*0D�ȪV���m����D�jQALr"eD���X�V�U��ƩX�2��Ym������J��V)R��AV6�*���XRڒ�F�VZ�5)YY�P�Q-i��H4|E}��t�5{��_ulX�v�ӓsw�0�h���^gc!�mZ3�S5�]�fөQ�l����7�nP�K�`Q�:LSs����S]�q�,�زOM�W�}�'�=*F�'+p*%������m&+���.��;J�f5
J�i������=�ȉPr#�xW^*xFe���U�wW����6q�L�frp�D���Y\�YU�ue<r��>�.%�Y��1��y�� F��V%*���rԍ���Q��[`��귖���y:��Mx�)���� B�_�͹tyK�o�ۭ�K��V L��~��S��~>���/��DxVw��	��c�ȥ��2�ō�s�v�e�{J�}�_ŕg�e3u�v<P�?b=���U�oB�Y�{�-��+j�\��UtQRӨ�|T_Ȧ7�j�İ@�cÅ���wY}WE�X[k3r�&�{���YC�޻�gظZ.����TFzZO�B����Z�߬�����}���wi�-����ڥ�#=�x�}��)��4���!lcB�	��3_�6��a���w�ǄKU���eB���:S��en��{>�n��F10*�S��{Ay/����>����RV/u��?�9�������D
F�a�1I9�d4�*Ž���&�nK���rhd���2�ݑq�z�Xf�fC����n����V��^��N��-�M#;�rZY���of.)NT.z����5t��mY�(��eE��'�u
za1�W(�V�''�csʶriZ:��y�D����*�����<�Ou@ƋA+�*�#�5�=oF�Fg��������!��G�vVȞ���J���	mE1hzn��%�u�1Z��_�wA���}GȔw%8a\V����H�s�P�ԥ\@���A�����Po��U�U���{�Ѫ��*iL4�!&\�Z����=x�T.dK����l����Lc���E�]��Ӌbf�\ӅI�R�V��,S�>���.xg�46����9�蕔�fdS��5hOeg���܍g�.񕺷��b\���< *�x4�QF'��%�"M��������9�2,�Y�6��~�������0��7�*^�&��\�b��m{����GV��O;hI	��3������)���n��50qNqӷERÓ�K�*:��]C�O���q�(��bA� � y}9�G����E\b�޶����P���Q� Z�����Q>�H����r�'�G�Z��ڥ�L�T^]noa
�ݵ*�ZU9��Y5gS�2Psi2�ݧ0��;�N��Xe�ţ2<��j�R��N= ���̦�f�	�{�7��q�已e@�[Q��CrWܗi.��Ʉv�#lL|r�����z,Z�A��+Tg�ؘ���N3>�S
�t5��"���7��A/�X�2�%=Kat�oH�\٪����8�0��2��c�m��@�2|^��"�Z;������Sb�i�/�ޢ�#��Xe���kd��59&5ה��q�w��a&�=��6U�]dg&x�2�]\��M?F��W����m��j����(अ�s}^Jٹ������4M��XJ,%Є�S���8�᠈����G�
>iic�eY��+t�6����Ѻ���>��b��3�]U�W�;��f��&P
��R8fD��&UtƁ;-@1e+�n���
����V� �H)�p�/Dc5��/ܑ;=L���32�d�Mz����qETh�V���۝��m�=��ޜ�T�OB��\4��.����L⸞*n��88]�y*����3���z������Sw'�t�V'N\ߐ鎓����6�<�"\b�G���ݻ���W�z��7M�g��q��s���w��/ɢ���p{����s��Qۼ�'}�49Lw�3V���Mt�}d��e�Z`���;f���^���9Bl�|���8�})�^�/W��U����'V��ݲt�osl�ݨW�{���VÆ^�i����:��[�Faׂ�*뎧��x`tqw���Z;-V��L���&���3j���j+����}�j��GJ���ea[�Vȳ���в�ʱ�]�k��y{�%6z(��$�B���ì9����
u5x|_�	)��A���i}��u�ZUY-����Z�*����c0y\�j�����W�\�H`�Q���0|Fq��%�q#rUO
����ܶzM@r��!�~_c�k�*�D{����N����@k�\q�i��]V[J���O~�c���3Puʷc�b��l�3GiϪ#��%w>˜�5�h���Z�f�6�N��T���t��h~
4���r���=i����8�m.Ju��=��H�� j'�y�z>�u��o��-�_y@���(T9[~�}���}�!�qr��@q�9�6��ON�ۃ�ʳO������Xχ=>�'�����r�K[g�=Ks�p�e �,t��H$���6w;=A��Ϩy��9L:/��j�=W[=��F�Wp��nC���[+�����䕜��+�k=��4 �t=�0#;4]�V�%��(;JΧ�^,3�^QÉ�r�O%���wX�>��+r ����-�'��$3wu��rLo���Ҍ���dt9J��o�׬z_�U�'t�����Os��K	���6Ex�C��jy��B�0�>��JV�܈Vbt7H���|][xo�����gy���@�eѩ^1�c�U�����V��z��T�h�p���f2�9� h�J�MV=��7�k�`es�̳yR;v���%�"%,�z�ק+x�^�Z^���˰c�rU�7�Ŷ��b{�z�kEus_+�N�c.�iiuS9Կ*����!��m�����r|��J���gn�L >�UK�84è��r��>/�Ǡd�v�%����T�!��
��|\������9��@�"%[ki<�C�ւ�i�IĄ����3���G����ߤ9���M�������y�*����{��υ-��K=��%�ax&o��KecY"��g�K#����ra�f�s-�c�U
�T���[�&oxb�)�ý�U�in��-dE{dZ�6ñ�
�	s��%�V��qk�����l�X6�r�f�@$k��"�<E�,�Ò��J��=�xi��~�Rw�J��Z�EWQê����/d+��ǧ�v��Ŵ���lJ�N��(������a�]��:H�F�:�!ړVw@�a�Yݽ86Թ�5뵜���W��P�6��e�ea0<�sxbv)6�������b�)W��UW�읩p����U�����*!WyV�Ҹ�Z)��#]d�,:E�q���bN�vpOU�}nY��m٫��
UyM�hKP�w��F�AgVS5H����H2�T�UP�l�z�$P��T�lTY���.�+g�y9�1��y�&���i�S�eD�p���Sh��r���Un��9������2�n��{>�n���10/8�3Me�������h�9���q�V�:�E�HuW�
Lp��ߺ�QX�NNz&�#�B"F��`&�.2l���5-���s�&�h�ğE(���`h�.��J��j����.ے��E�~�ٽ{��'\��8���q6��c����?Q�*�V���y�!���p�-�=/�׭�vQ�ˡp�@T���:Q�e�<6�k��'p���6�g8���\y�s5���2�*�qRq�=q�ʡp�"\L� 60V�)��2��#1y|E���uV��dΠ�����[.��ߔ�{9ns^}i}����fL��n:ض���:�4-�n��j�t���*{���ETS9�>��ׂMiiWeb��j��g]�ƧF�P�U���`#6�nf<LMe�7�Щ�wl%�
���n�g��/Jƹ���zvp.��A˓�Muʗe��w"}\�`��M����_��*'���@�Cd��L_us�T�{�t�^
��0����f:�u!,��9��K���L؅ѕ3�Q���Nʱ�!��EM�V<�/4q�t%���fzxez�;�������t�$2�@���� T萿Y��'+Vn3E�o����jp���&h�^���ig�pr��o=� ���h�]�z��Q#v�s7��Q��§91;-�	��ұ��r�W�Y�:Q�گ~f;�`F	9�v�M&����^�/E�U�(�^�.�{.�c'�j��H���͋���{����|���l�?m�S��r�	�g���={���Gz�֌���92v���E�ۗg׃k�]���>u곁�]f}L���`��Yu�z�L���>*��|0Z�NՆlW8��^��A�ez?��iz&�A�%U��(��6�ﯩ_����$�Qx/=8o�W���ԛ��'c���z�U�����:�u��tQĶ�
�}չ��So���%K%�t�����oب�fѮ��.�Zy��8)Pk�葤b�;S}��Cut;�J��K�;�T�f���IjlW8��k���y�5Í��2��l�:�q����5�m�Y�wha�������JP��� ���uP��1+%+����!�B�U�|��	��;�%c��F^��� � �ϔ����]|�s²�M�
\��m�_Z*b��
����l�Ч ��h\B4���M�2`�1,ޝ[�ꜥ��È&�aٯ:�T݈\�_amV�\��8�׹�*�*7:+r{U�F��^$�k���'�˨���m�&�Yf �S㎵���qn�z��h��ֈC���{z��sl��0[F&&�r.E@�w3g���-��PS�:����-�Ӧ���B�^�.:D��^3�d�5��^��)��J�D�.E�Ư�E�h�=�VI�k9�V�H�!GĹ��EȔÖ.�$�	��L\�������a�����S[��e���k���Uu2�1�$$=�!:� �i�~��X1�F��Tg�qG`dr%�w����z���|�_�@j��xVe]AVb#ޕ�S�Uޙ�\i��h.�(������\�>*T�
�X�,@nB�����u���ۼ�#�}��S^� ��dhJ=����U��n]�PAP���,^" ���)�?u��lfм��\�9���]mn��Wp����4�!wF-�Y�Ykcl)�+�X�u���2s��f �+�V0Ԃ�w!6j�<\8��3��l���GS�N�5$��A�L�NT@C�9on�O���Qz�f |l�ǫ\J����Yq��j�9:C�EUK����-\��l�]����+�Ӛ;q�X5�v����X�i_a����^[s8�'�m���+e7�RQ;m�:ŷ���F�}Q�(k� �ʺx�]��ʣ700B�yo,���3����-��1̉���N�%�,�L6F-W�X���x5��P:x6��:&(�������C�]*���[#|9�'�R���h&�Ņ=�1B�m;�`RWH���x�f�ɪ�n(����&]�B�U�T�].=
�������f�d�9QRt�9�}
-`���9�]������TJW�e4�`�@�X�:�==)A�J�o<F�v�.����W��v*];�WlK���j�G[��m�D����)\X��:�>\�m{�L\%����;�W
��Vw�L ?6ȟ�
A����T���@wb�*ۧ�W��:�y9#��:��ut�ѐz����ޑ��C"%\����0c4:��V}���C}=KNj&��d^tޮj��יG0,��	��,�����&��wR�)9G�����gk�;�:�hp<ս���pN�ό79ϧ:Ĳ��9�V��ACX�0���
D����i���y(f�o;彽[�Z�����oB���q��{l4"�l�^)㛇Zr'��"$]d��
��«]�IZ�\���9�!��UFp��ױ�g+�I���Og�r}܊�yB�̼�4�Hڌ��dKF'��Q۷e����*�4�w+�M@�TFʰg�����H(IH�s`�C5�*��ʞ��ty
3\�U\Y��L@��s�0�2�z�M&��n]Nu��xun[	MD�c P�+�6�]�p,,>�E1��F�ȖC�j��I�ut�c����z�Q���������\kh,�\�5u�/��#{�Dg�+J�|@:����V�>*�z�ɥ�Wt�~c&�Qx��tLS
���N�Dg�^��{[5�϶�9��]NL 9�	ֺ��n	~�y��>V;�W]79i���emT]�.�}p���99�
�53�+�A���SN*vn��O� �����砇~U��i�����)b*nkQ�Y8ӻ�6��.z��Cلݝ�%�=#E�$ʾ�9F�$�(yD�� �N��+�r�C������C*+/�f	S w��K��SYJB�I�W�&�ҶMz9�]}IsuYt�"������ت��z���R��z�tQ�d���8�����wJ﹗F�
���6��X"y]Q�@�c�u�1�)�|qR�èt��x5���/�l\��5��`���)o;�t�s�Lf�#�|���d�#���&�����f�zF��^��iZ_�M��Bܨ-��\}j�om&�Ӌ�kВ�^�9 �8�E+���a�3�ě�v��s���մw1��!A���XB|�󎭶7����	�e��H4��\��o���6=�u=G���gY��E�/����j��*���5b ̈
�����U�j�1�3a��2��z��oy�&u	.Q�`PE
�K�qk�55��]z���h�(�v�;���R�-��ef�jؾ�?J��)m�:��"�,χ"�'Y���������ӳjȊ�]�w٦�D����)}�K��;\��4@�e��o[�j�bP��9L���P%[�+�l�Y�i���P\ɴ�4n��pz�vc�m/'gw:Zq�m��/�JZI�5����u��iX��kW{����rz7)t�s(�	wl�Wm�/^7\�E!����q"�ٸ���k�%`Q�
k&ͼ���gfrW �Kl�e�Ʈ ���O��j�s���w�\������e�λ볢+2�:��2Pv��ٓ�wM�Tg�*�#��(��ۮ�Q��f=�I0��#��:�h�(�2_�]�#CV��(��磚��9ع��o����i� d�R�ty��Y�>`�F�
�/��u�v�;ٛ&|�,F��V�L"����A�6��hpi��-�j��9)*���$�����-f&#E$��p��Q���]n=�Zq�6��XٖNC��&��3:��>�כ\�\�ύ-��i�L�2�N���j�G��8��.����WH���2��tnmQ�B�K[S�B��j��Vk����pbem�qb��&����SK��!�Nl[�]��c��Ҵr�VX��Y}�x���A�-�җ�HO�R'#�5VVb�2!w����P3j����x��L�{�̩�7M=`=t��C���w�Uғ������&��m�f����ҋ�J�v����g<�43�2TEmܱc�X�'��i���+�r�Ls��O�;�f:��oz��ϋ����3gE%|��J�t��S�=V�$��~�Pĺ���������:�=����+u��Lr��J�'o�V���.��	T�%k��N�/+W7��5զ�e�mE-|)���nK���a��ZK9�/lP-e<ku2�摝5=!�=�lI�5N�*���I�zGJk�y(�qA�Vs��J���ñ܆)�5u�z�K~|��VI�X��ɽ�-�ړ8kcB�w�t.�	#�'5Б�O�JPf����ǭδ�щ�bD7I��
�nN,��fы���|���>T(��݌9R�^Vwv�*ȥ�En�(�$�����Ԩ��Qe�V
ѩ[FV��AJ�ܖ[C��T�I[KP*EQ�(6�m+�H�آ�F"µ�EU�P�m�JU��J1B���*V��ij� �J��TJʶʍim"��E��*R�lmj5+UF�Tm��Q�Q�R5l+1�R6�V�����Z�@R����2ڋ%JҖ�1AUeE�؍eKZ��TR�E�X-�
U�X�l�U�eJ��)QUUdX �@Ym)B��UjT
�+*X�)�Q�1b�U+BV��aR)R6�ڰq��cl�KEEF-�#j1R�DA�UU[mB�ڊ[EYQj���b��PQE�ˑQb5����e��J���["²���P�D��+m"�*�FZ�Z��R�X
(�ieE��QV�����R��B�V�"ԕ��(���e�֨�(��k
��B�,J��*��6U���AQYR��U�|� >@�gt�si�i�T�G]�|�7�J���s���g�=���D��Vh�����dȶ�YUO1��<�G�١�A����23��Q�cU�<��.��6����1v��n��G7�ʸ2�֗��4�$����_�H~WًG,]�=T�_�h#�-vѮĮ�%��-��=%�3�wb�2
�۬�f��)�Uǥt��c�-�Nˡs\�Ԥ�:��"*J
1RN��g;&JYNh{J/'&�]qw���`�Lg��0��ҷ9�[����t%�x	���B�����M�]`ً�"�w ˨��s��ڨ�7;�e��w�'^�[�ׄD���[,t1N�ζ����t6+�@��#�=��:���d����W1�u7&�1�]g\oe�h����2��h�)B���w�g�!j�xZ~(k��W���m[���X���&�����y�Mݣ�;�,?R����i��W�ȕ�Jr��b��=�g[B��MD��[�O;����7½��\cj���i��&D���#�[��disWu��ի��i�2	�VY#��J䮀�����O91+2ߨ}]uڞiU�2A�~���cn_p��5ü�s������X$�訫z�V��c�m���d��ӗD\CU�C���s%M���~Ahj:v3�]^����>���n��G�P=A'w�4�PК�<���E��"Z��}�����G]�+�Ev�Cs�u�ĭ*,��躙�(�,��;�Gޠ�kVK�UO]�:d�u�5¥��{"TB{�����egd^<���;j�u`R��cf�]Y�ծ��;ҭ���
�;H�U�����םL#Ã�[W������5���`�C���J'�}��Dި:��Ǖ��Cv�Vw#9(��I���ϩZW����xw*�I�R/k�GI>�]0����V��Cɾy,j��H�ǳ�q��eL]EFB���ʛ�,������F�>P: �k�p������wI���\ό�9R�T]6�/�1p�
�����=
r ��� �)�$����=u��T8�wus�UlN1T��^�T��ऐ�ӄ�sp���P��:Q6�7�_n�kN���O����AYP� �j���=Q�u�_�ge;�}=A�s*[[�ik��}> ��_�

��~Q�n����
�EC|�?G����9�M�A�/ �;�𨭵�aMۧ.zh�k�N>�2�d��I�������ٗd;�Hj���jv�w�b�x-ȟ��_x���6�z�vu�Zw�+����i�hřۣ$�E��@b[|9�E�4혭�|�X���U�;(� 6h�����;�y8�����3"'�{�p�ƴ3c���.N�v��Fn���ܮ�'�U���v����h���*ۇ�J3�Om����v���ʠ#�|<b�uw�S���Ƃ
�n�C����':����m���}�і׾�Y�Wt�
�@��� ����c$1�X�*�Ë�b��Р&�7|s�.�sd�� 2l3���F�5_�E�Y���Q��)�Ԯ��3�%���N�޵\�];��7�
��.�`���2�A��c������ͧ>��jD�f�E���ު��i��z<MK�x���=X��*�_�ǅ��T׭3�{t�QN+�ml��֘�����u��2e���Tsj�ߞ�����Z�����U�J��E��YXX�]ޤ��U4��&Ne邇c�s���M׵U����!m_=k��ؓQ�K�fvMk������;�Q.�nℴ�����"-:���ʑ��TL��v�|����K�l���T���� ps�d���SSu��hM�]�R�S]���>܎�˻^�=7'�?q&����h�eo[�����|%T9�r�0�����~���{PT��^tz�̶�J��Н�1�����xs^c�<A�}��NI)C0l�Cj]�d����)F:VgR��+���Q�{�v9˔�g�uu��ڏ��b���4A�3u��
n��;F􅽂`ʼ��3-C� ��]%�u���-%�=f�nй�n��0�F,�v��Z�����8���-��Ҧ���u(�x!_���#�Gȕ���Z�x�y�ȗ�#�I�ԥ\1�q�&�����GQ�� ��L���3aQ[��A���Zȋw�~c���K쪞�J�ͷY1�H�D�n�4fۣl��a��Ƙx�z(�u(ɼ@��W^'���WL-��ߋ���zF9��l"%_��w[�'N-��H�4������@��_��螓1y�؋*�n�;s��Zr'��;���Fx�ʁ*o�{�\u�ʊJ�c��U��1������4J;��R�{�S"(T9�.�7K��&�8�JzYt�}�4vW��g�&���)5x�`�S�!+�xl�W7�OW��3���=�$7� ��~�Y;67Abf��
tW��d�Ʌ�r\�c� �|��g���~���0o��۩>A &�s�3lF`jA���"��`k���X !q��k�}s�� ]�-c�t�?Wo�	A��Kz��޹FV�������TFz�d��4�Ah��"�)�����W��t��j�T�Kvj�tp�]�sY��fn���I���OĪ��;y��Lש^������]`2s���U�L���WP7�፻�>�n�.Z�F�(�(�b}�qd�5��ގ%�%og'�voY�����rԱ�7�v�6�7��b�L#���e'p�ca[>��N�DdW�*m�l�F�IEȩ��Ӣi�9�p<�������"Vk���{�]i�*�4 �g�ɈZe���/�[����[��)���Y�S,�����ʌ��	�[��1�9���XzE9J�80ھ�wEk��4���vtr�`�b:I�6p�MJ������s��e��`������F����}���*�èG!\��E�u�W@�j��%�`�|��O<�x�[r�{1�n��!M�q�].����|Y�d_��$��ۯ\�����l�|Z/sE҅c��/�FQ��.�S,	��t��T�4��{4��q�%Ōۉ���Q�^uP������Pm���Z<�N=>�Lj��*n�i�Q�:nx��t��{��啝��6d����.8���+��!\���#�#؏����6O��b�;����*���� �R߳:��={Q*��YkU�X�)�x�O��la�;V]�=��U��|��?X��u/mf����͹R��g���z�lg�4�v�Ũ��՗l��m�xQYS�}���Fu3A�gu��V�A�9a�� �Ѥ:z�˧L��x��ᆘ�pI]�W�\Y��%S�6�.^�5{կ*=�!w���0�}{kد7hbKgaA���L�6\�"\�3ꔝ�р��O;�pN�LHA1���,���oV<�u.��R�}�A��Y< !��_8}��x�!K=kv��w����r�����a�V�9UNi������:�.�U�R��G��^�i��C]މh�ND�ܵ�^A'���V7�W�1�>>�P�`VSp���	�.|���������U#�@GL�θ\@���^ˬx'LhXg���Ly���3�z��p5ּ/28{/R��K��f�8Y8����B�ST�t�Hk���d�1�GN��b�њ�V�p���r�sc3�����kV0h"G���5�g��jTI�-�nz�d�`Ŝ⻡�i ��vy��R�>>�wy/c��J9�T��kCc���iP�o=��Vn����4uB�er�(�^N�3���`c�1��PDd!l�ʛe��2����"'�pt��b�]��kx �J�Q҇��I���Z*aLV����6a�S���E��0���rT�WSΥX�6��⥛�o*�D��9V܌��:��)wl`}�����[�x
����(�w��{:T�q�X�íb^z[>���9l�ם��� ͡h�3h�̙�N��˶0�V#�xm-����@�Y�b��
� AU�ۣQ�v�&h�\�.�'�al�[�'.
l���.\ߗTt�Y�mB��ݕ��|[FjS����U�;)�((}��Ŝ~��{j�����)�5�}�W��mt�᳓��bw�Ӑ�\o���ك�Db5��
vJ�����uٮ��K;�St�Lt�~�9�sGŮ�9��������GO���XVߕ�,��y\�1W�����TV#
�C����.A��rbaȕ�����s徚ү_t��[�z�>FL�kg^�y{ڽ�Uj
�Tx���]�+x(=>�'�����ý^����-<��q��b�A�N�X'��{�]��1݉ʅ}&[L",��W���Etk%���e�9X� w8������a�Z�:��^>�J�x|�G7F�+"�z�ʑ.[fn��j�;@����T@q�0DE˕}|f�3�����wn(��O$�Mp��p���_z�z�2�o���O����Պ��WƝ#a����K�i�ެ�[�ݍ���Z)(����T�Ǹ��Q�Z��%[eL�e1]ݗJ�/T	��{���Ŝ���K��J�Nhh��D�����<S7|9AӰ�ޫ|���.9���e�Ғ=����ێ��˵	[2��zaJ\Τ`����y��I<��a_p2��Ov�W������^�d-�/��=���"v��Ҟ����յ����¿.U��H��|��
@���U��gzl�}Q2,���&t�is�D;�=<���S�F�ɮ�>>�[ �aJ��	��B�0�>��Jq�A��T�_M�l'=�����P����1:�PS�\Mz���ʅ>���T�G].>s��}��H;����RWH�W#�t�|;��{�^�U~�76�� TJW`��ah\�`�@֥��	]���ę�z��s�m��V�? �N55���Ȟ�َ�c�J�}�jl)���A��ޭ�l㩤��등i�7�e2϶R����q�2b[t'Ǻ��蜭���Kڠ
Qݶo�F���t�(?R��1q�f�䋚��&��a�"t�D��$�j2��Ÿ�B�7T��B��I����}Q�GM�f�t]7VS�6�ND��X���}</�9k���.�|g����Lt߇#���1ʺa�Z���֙���o+��+\�L��f
2�eÍ�e�X�tRd��R�N$��j�h*I��,��s���x�җ�G˟�����,�]"{2��r�
fIE/[�Ύ�b\ �LiK���F��WP���[L��5֟��]�,b�XxoX�u-��Փb�Wf���u=��i�E.Zm����i6�3�64H�p���/�h&��SsO@`���&�=Y�����K�q�:�A[��g�'Iܮ�P{�J��:��j�t�箲v�M孇�xUR�/Й���2����y�.q�5F�>���v<�y�|U���/��R��j��7
�z$�z%�B�b��6c	������)�����-�W����HJ�ZY>�*.�z��ngL�B�WP���(���Ѿ��C|h��|;a���B���^�Z�f/g�ܩ�M�+�yM�\3�·^���4C�b*wW:p�/�j�ᒯ5uMr�j�6zx�>���՚�a�^Cs�W�RK�^+"�-Z��̛7ު�K���c�p��'��3oTR��%W�p�]��c�@U��Y��=1*j��æϪ��e��ܶ��:�^׼�0y�]WM�"jP#U�fܨ��4��.q ��{U���'5�jr��*�����*n��.�j��%��S-ឮ=c�K����7^��R��)��\zVG|}��д��܎'�t5p�=�`/;mAR��^W]}�/K�1�gN���*�u9t�{"���˰}Y��n=�ƺ%�J��s�H�>wz�ӛV�,��|�ҭ��,D��uH�N�p�X���嗼�����kT<�^ֆ��O��µ�e�|2���te���.����`�L&����xҺ����Z8�p"n�zi�=d݋�%C\���aȘ(-�z�J��m6�/щ;8F�ۄ��zZ�w����`e�̩��p�b�yA��@�F#):__O�}�Y���ߟ��[����䶲�W/��i��b�������/����cM��"pB9S95i�NeWFR��(�N��4�9�S�h�S�a�r�תRtf�D`.D����߉��D{�b���س��f��N��]�t W����a�)�w�y?GM�;�^�6����.m�͋�vs�}���$�ת���W���&7�ۥ}��K��X�@��"h{Q�Q�(��|���0�:�A{��w _i����g�`B�����[p,s>ar�n��F�n�+[[TQ�wD6� �p������=v�=���DAu�_)��e�ب{:�=n
WWG$N����;-!R����P���8��Y��1ޖ�A��0�pyP,oȝ�z�OUIvw+[X������	[	˭�1�Y��W��J�W-��L��E>���vb�/6�󕶄[��29�+h�ו ���t�`�C�R�-gs�)���,w9B;tK;�2	DBm�X��Q�r�ԝ���	��լǲ����S��[�
Z��&���g[0�9T�}w�y-˔���j��t��;;���ck��s��Ts�Ys$�9�io9�"��:���g�ֲ]�U&�Ko+��7�m`5�A[y�ٸ�ەݣ3D~W��o���� �-���F!�
�9\8�7x�2Dd�N���t��_�N��G�J�
����Ji�N͝W@���%���Pu8/�3��K׀W	��Ԍ̧��gW��ʷ���ҏDs��fR�V��VZ[#6vo����w]G�R؛ݗ�R�fnuͤ�]^���{���Ж�V�A*z%�Qv^efW[�v����g;IuX���O5�o_
�S��	C�n9��������Ld���\@�*x*x8v��ܭ�E�.4���ӵ�9��
\���t��*,�v�����tYz�1u#o��I�Q ot��	Fɓr*\_�" ����ۃfj3��o/u��cY��"� �=��Io"�ij�k�'ٙg�;�`�w�;!��P��Lav1�*.��%]X��7}*���ك��y�)���Vx�����G�D6��O�,��	�ֶ���!5ٻm^�70�"��3!�C;f�jSv�6�e���u�O#)��uv*��G˷�^�P:x7��uݓ�ս6�K�}����-��t����!L�u����.먁�*��k8&PrKט�J(�[PEA�����1W-e]tB��u�AmW�����i�&=2�B�����쩂���_Ƚ�ڵ�� �;�2&QڈuΌ�[�ju��
��L�hV�̍i�f�Z�^J�J�w�C8���Y2KW��eh����4��c�2�mέӋ�7{�Ϸ)tY,�:Jb��J������sĉy��Ѧ�AgFFҭUw�ZM���{!��ޘ�ikߒ�{n^��Ѣ���o,�I��F֨����N��S�L�᪶�m�@��I:͠5�"��L�ҭv|��(ݗ�uf�U�C�H��F�E_��ڼ=I�)7��޴����׹�ɉS�Es	b���6"�$��:��;1��2�0�1X/w��m"t�fa5;�>}.�9f�*�@�/s�\M!@Z���u~��1ْBǎc
a]M6	��@�t���pv.��DѱR�5e;�kr�Ҧ>�5�ӄ[��[��颈�V�e^��� ���Һ��g@%�^$	zվQ�/�͟NtԳ/]4WJTh�r��-Q�YZ�Te�@X#*)X6�YYm�J����)J�֕�jT
�kb,PZ�X�����V"m��ёJ��եQ-*�m@X�-��X�m-[YPR��RԱeB��*�H�UD��B��b�QV5�"#[J�PTa
ʑUaQm������(֖�Ő�iQTV�Ң�b�%K(���R,kDX5im�mF*��U�Ҋ���1�YU�e�E�UUk-(�ѵ��mkh�DDFإTU��Z���)R�J��#[V�ڂ(�e�lkj[Em-e��0Ab��" �����FX�dEbV�[JZUQb�b�QU�[KKVUbѪ֢[Z�j1�e�EV��Qm�mV)R�EDb�#h�AV,`�X�Z+l���b
ڶ�E�KjZ)Z��6��[-�XQTJ�ڥh�%�U�UU*V�)QJ�Ebȫ-�VzkϾ��3.��>�	�/5t[|$�s��\^��]��{��㹚$������jd�[5af�H�8{�L��;���w'�w$儴�R�*�r�N�,]o{g�u�֮�g���������,u nmR�����R��
���TB��֩�ћ����g�٭����^O�Fm�-Eރ%�8�@�c.`�9�����,�lFC5��/ܑ�="�k��!w�v�����|�<�J����N\
�.��M��W
XzǕj��c
n�Y��v`��KZ<։͍��+u�W��/�>�hpՊ
��ڢ�Sv!pRn龬�N���.�e�i�[	���1r�n;L�uq
���%UR�������b�?O���c,�M�"�7yV��geN[�w��.E�ӂ�l��t(/yxQ�j�J3��R��cًb�2�i�^=.�z�����*\X����)�s]���n[�3/#k'�M�"T>�#���"o�e�����yA��n\�
� � �?p,�F6&)�r�\�.A	�%��Y��ML~��83hSc�r��t:�^�okbX�*��ڌ��ȖǷdRuq�j�*!�U���d�6�W����˹*E����h�Ƞ�q����h�㵺Gs�e�9Wb=�$�5�����Ԍ��z�e����9��ݖ��v���fu����Վv7ݡ؅< ��sZ�yA�/��-��ܮ���D��eP�$�pqY}�#B�|��o�����ib��C8�IX�n������;5'n��ߧ*I�2�ހU�KB6Z�`M�S������!�{fb��5Xg����'J��ǥa��g9����z�)��[�������IMdbW�&�yZ:'��̗^�Ud�3><:�[��I|<��(�y�����޹lӉ��˒���\BxjL[äusKV��ѳ��U�J�׻�g�m�[�>�.�����pދÃu-?��c��̫^�S��^�H��z/%vK�f��s/7�m��sc�8 �yZ�PC�]���GØ�p� ���#�#��;�{y(%�%f?!�i]Ws<=�n��:7���\>u9`/�Ǆw��66g�q�=��9�Lu�F$���pMgMeO`�~vc@0�"wr>0��TC0��|�w�	���{rvI��.�ن�~:g���\}?|�&3�C@��I��3��>>�R�q��B�������W{����#�6s���R��s�X�E�d6nD�#�IJU��8�A;*8���i��>ꝒMg�|@��"26�V�޼e�_o9��m�GBG�kR��rI�w�}��з:]�Ǧk ��\�����ק���C�V��Mo����G��q@�%#sv9,Vb���aWY��w]�t���޺n�>��L��^�<J���f�镻��
oF�5��.��7/��ت��mПwR�[&U����k.�7�c�Fmu(mux�n���`م����ť���x�%X�"�vS����z�T���X*�d<n(<�ﮘЅ]e�x�|�E>}��D�'�~;Yh���&��q>mTĢ�u�ͳW�������-Z���[`��h�.d3�׮]֐S��-�8v`�Tc���le!��+b�*kY�9p��\��eS�yn^fG�ǅ��|Λ��V�E(�إ��tI���0S��7��x��x�����F��+91.2��ȴ�vuSR�%1��I�ˉ�OD��\�T��0~�G&�q5=�Oܧ+��M7J��;��3D�0`�f�s6`�=B�1WPu�n���Q}��(uu��E�M�^�<u'��ʺ;�k��~�K4؅ヅ�+�*�����1LR�}'����6/V[�4�:'8���-�"i�`w�.�ɬ��a|FZ��b�Au�φ_ژ�w"�0�
�}tsgcm��I�F�b�0{@ּ���]�b1�;K����t���7笭~�L?I^�l<��-�x5�����cz�Oh�3�ͭ-1�C=K�Kc���"����%��T����˨s@d����Z)�I1�fE�`+S�f�7�g��﮴d10	�vT����)z���V�p�x��!2���'��$�1�-��ұZ�������txu^��FC�Z��֧fPH��0lL�5m�i���R��f����j�ܭ�&1�jq�w\;Dba�%M�:��(ʊ���N�8�ݻ�S�9!b4Z�(��.3O��N{�C�q`ݗ^~��hT�%���&n�!B =��7댱z5}�%@?�P��:wW�DX8�)�hqSx������=j�y��z���G��P�g�V
�E?����L^�*���`�g�+Z��vD^���R�|o��і���Vx}���b�1�2QʈuP�06�PM�u]
{����q[��"�]C���GKb�a�����C���cM���hW!v���w7�MB���3Om�]Ӕ9��y|T��0�9ck�):3\�,�:P{�NSy,U�g��h`;��)s�����8ϸ�EL���<iТ9��W-1NfvL�R�������������������0B|�vU�v��aEY��K\�N4�轒��{R,���\��\�}Dt��(w�س&F7�IՅ��c��ˡ\EFx�¢�
�e��(fhS"��l�������f�����m���v �;y��o�5�f�䯱FpX�,�����{(�Ft��=>T���5���X�̓��72y�TK�&�i��qY�.�7��*Ӌ�a^��WU�Cޠ����Ć�u�<��ɵ�"s�{7E�3���������#1�4����>���`}>ƅ��_pYZ�sz��T&�L���o�dM�'��3��68+�%�ك곁��u�)�V邚�`s�fk��w>��h���~B����9ɫR�+ƴ`�D��z?�|iz.����u�ڃX��
5º;7��ѓZ�3s�V���3�7�h�/����t�@qfV���z���諻
c�T���n��˘<)C<��|�3*m�z"ٮ��F��41FU��uI���cD�.z$@ұ�KS��{�T��鋎t-�Q�;3��qj/��W_��畚�`���fW5@_J_<���A])��T��v�"��9wto�]�����,���L98�压ڸE�..UDZآ��Yf�(C��S<��]�O=�����7ƅJ�����T�b�`�gm-�f�Uy�����2���tE�!=��u"ɶgu��qk��FN �އ]��wY�멇��vv�ΉI��W���=��B�w,n���ړу���G[۸(����!�;}n�z�j���=��LM7NC�~��p[����л�WJ��"��@�j|#eeҞ�4|^�M��s/���&�P����Q=�5��;�k�S/k+���"p)����ؘDn��9z13�aɈu�"VD&zj}^}h��yZsVm�-�)F�Z�'5�$�;�Ȩ�蜝��>�!��	��v�/�\h�k/^��,:���7S�G<i���8۵c�ko�/'�����{o���[Y{d7��*n� r�JՑS�4�� im׋�`��f�����쀹���� �Orc�˼�.UR'=�-��	�CexW̺�F�B�:J��h9�L�s�nr��t]A:�U�X�V��.�,��V��Za�Ѵ+EA����MK�^CD��]4{��'��Ga�R:j��Q���C�:|^_d�^��+ت��a�5�Z�����ed�`�h*
�fǸ���0�:=ƞ��6v<�ؗ��^���&bNlHBő�k�
V��Ӽ��tF�ݘT��j�m=��FI�?$����[n��u��G�����d� {}��\�z�U���
��m��3��'R}%��$����H6*䢝��{RN�<���N�>|�S���F���Ir���\��>��:��ά�x��xT�k����a�&�G>ȵ["�AOMJ`����5&/q�t�(��ئ�|�yӗ�7!Y��a��˶�p::E���GO�4�HWU��F��
����k("s{�~�*�[�Sq�����9�!*�"�|�*etW� 
��0^ې�Iq���<�\�eq�~�!0���ԩ2秱����gdK��Z+�3��A�a8n]��睸��{6:��E l�q�B��)�w�lk�^�aݾv{�d|̉�EF���{/�Zy��L�}M18ʦ^��x��z0l���ס5���>���������:�r��]�9���!(r��T���Y���R=��dwvו�o���8.q��ش����s����Pū����F�OL��X���\�6WA�����K�ڷ~�L�}�.�0Ôbk]HO�23zj�����oQ��'�yj2�c���8`�����c����KĪ��.���wj?�����d�Nu�����yU�v�w��m����_>u{�F��4X�۽�ǅ�8#D)�5rP�c1�Zt�v�G�!}���7۹�ɴur�rw +xnwΚ���-k�Uf�NK᥄��7&+�e�[���]���N��yp���a�]l�UDN0�.���9��X�_aI��m������и����U�F�=r���T+���4��5�$��ggm0�G�N[�+����y<���f+59N��[D�yc�D<�7��ң���B�w�9j�p�hu���a��]���Y٬�' �m��K"{|B�>q�^��x�F�i�"��`�8�OQ��y6�^ӄ�y�U�M��>��aG�!�*���/�j�3coa	J���V�S��LyQ���<ˏr����K�cB��
d3YE�Eޛ����6��#a4�ä�s̭˯���p�Oc��.�aP��A�9{&�:
�t��]Ū腪�C��Z�)���S�j��mG1�՘n��oL��V*JW�������N����!"��|P+w^t�s��5|
EȎEa]�j�����k��q+~�ٰ��%l�Wm
Kj�f��fmg,7��-u�{��U��h�]�P��.E��_�P��s:m�����Mİ�1c���!���K��d��z:�,�ήWW�oe�.兾������j�œ֪c!������⸥/�U��v�
����O�n�瘔�~\����i>onD=���uD��%����Hо�	��}R�]U�=������Y�\���Z�L�l9GҰ��3)Y�y߽{�Ft��.ב���I��-0��̳�:� ��{�7Ү�}5�,��\3��UZ�<]K���yE�>+{L� ���+�kq9ȁ\PǷ�Z��ݘ�ui��*F7B{�yyi���Õ꜎>�1Wq��^����A{���|�⥬�oat�y\ӻ)g��N6���Ǟ�Ϯ�l=�qw6��Ow(H$@���u$Ruŉ�zy�u	vh�1�	�Mu������X�K9�n�bڣ�� h�J�%��Aѹ��o��R�)J�s��^���'���{�nv�:uq��r ֝��-{�~v��5anf[�T~��Z�])�tZ�b�fC��maF�Bn�Ꮞƻ�X��ք�G��-��|v�L[�T+0n��篷;u�V�`���CwKњc;�rd��ۥ�c�����S�. ��ӝ������8*�p(����h�t�rb��1�v9���Kogc\��X4�r�/��Ȍ0��iML���%�=����A���;l������x��ɽr�1/��Y��m��S&c������7�6��Ci+���1(e�P��mlZ ��<�\�V�&3ۮۭRuF`���suܞm�7��Sn\�@�&+�>ܝ.�u�Sv��:�'ݺ��`��0�㷫j�Jf&:/J��➹U��+��3Q�p�:����'q=��.���"�^�Φa�/_����ti�+�;WSu�!��4��s/*ﺘ�\��oww9�-�EE�q(��70s�Q5Wj�Wm�lh��m=ΛJ���%.��Z��^\!�9���$��(s��Ƴ1������f/��(���X�+WC�a�ղm��=��,��q�M�i޻sq���5۔�5��݌p���ӵp���5t�;7H�n��}LSWYs|i�׋>�f64�8,@�va���J�u���§�3���˼Z'��n���<�i�5\�z�u������lJ�N�B��[�:�(^�m@n�����B�(��aw9��"(��E������63#�S��u.��R{݁ݕGO]����[����$�/Eg)�����Z���g[�2���@��RT�P�2,� �� s0��ι��[�\���"�B�Os��n��MXn��(E�>}���\�j5�{7���u�o�T��%,)���gvl�҄i��f��δ:��f��&,3�u��ӄ�f�v
��H�dG���q[R�`B��	.
��]��W:�š|t�(-vC��jy3�4��I�l�=
���Ȭs���w�n�S�� ��Y�h�֪V2��%��w�{e,�H�v�,�P�,���v�Yʫ�Y+����|E��l�9��&:�ÛUy�y.eu�ͭPM�ŻfȒ�`���*]� }����o-����~U�v��;�ށ�!	]�/�gjn������Sh�\Ɩ{�v�]AiWӍjҸ�uu4���g�Cm\A*b��ޮ�1�=Ҵ:D#뭥���p����-��P��Z���}�v�k�M�B�\m�C�К��tF�P���ky2�B��K3kC�@#�����'
s�]�"���P��-���y�:�a[6��4't*���ٔ�π�����|��1k�MӢ��t�e��d/���[Ǖ�9�.����} (1t6+|��/��Q��N��̻�ݝ��岻rDnB���'����.���=,_ ������T�
N���y��wY �|%�ax��饖NNc���]Ѡ�|emF{-�]ma�Q%��o��;}n-�����VǊ�����Ҧ.;���Z��{(L�9\I^sT�˷jT���o*q�� ��pe=v6Zz���1�N�\�l/�;͝kL�������x:,e���v�s��⽋�ڈv�6
V�P󀍔3.�w�r�q&�
��՛������7ҭhj��ebG]e=N��5��	�&�&�z��H�e��;%�������Z���l���Q�w��3���w �vQA�]ݦ�� �#y����R�"���+�E:���W�S���
���Y������`�o�:В�s�p�^�V�׈��a��R����g^�ZIr�k*�|`}R�2�N�۫�W�"�f�p$��m>O&�����L����]F�wB˟"0gu��%�Rz�L�c�ۏi�w&-��7g�����8X�n�1%�'I��1	[��<�R�2S4��A��/�n]2��;����t�֊~;YA
�Ad���SQ�h8�(Z������d�7�u�����0���Nk뇍���ޗ+�@� ��c�$�c;�x���]�0�*S��
Ҭd@�I���/�hv��S�y��X}�~���߿}X�T��+)`��ab����K�R���AjJ*,U����D-
T�Z��6�j�K,�E�h4��Jы�-����R�(���+(�U�(���X�Ԣ�kb���Q��DH���U��(�"�V�Vڢ!Pm�����E�V[B����DKT�FJ0�DZ�R�
����E��*�*6Ȉ��Z�2��X#b ����!R�++-�V�UmE+(�Dh��
���B�Pm��U`���jU���X��U�TmJ�Ԭ�(����	R�DTmj-� ����H��QX�Ee��
"�m ��Z*���Ȍ[j*E�UV ��h�iR�j�[kԶ�`����*E�m���(-m-E��ƵaiEQaiD`#ѕ�`((�*#���E�"�������(ƍ����
(��b5Q`U�Q��j"���%�R�Q(�mTT
T*V��Qڪ(�����<��a�u���/�m�����;Yۈ�t>��3fgNfw-�t���b.�e��&��a0�*3+��5���0�e�Ѽ�@0~�r�J��W;��9���q�{3��S=�3ce���Q�j/ViP+P��sڮ�uc�5�N��g���1o�-�m�MN�Q�jP^;U�_!̍����^��緂�LY��o����TUꞦ�=�`d+9J* �F0*���^�W[V�E�|D�^�Iwy�d�k4�dQ���dT�P�l�[K�{S$ng6����^Q�t�u$����,i1={���U�Olhf�	�����]�\��z��v֨mg�.�r��W�[��K�T�5`h1�&��y�R����Owlqz��q�5~��0ږP�Pby%Z-�c����N\(��F�̓�S!&i�]s��ʠ�|��c��}9،��\���Oޢr�������ۚY[P/�4�o�����yȲ���T�`m�$��B�t	��{G#K����>uA�Iɝ�����T�,�%��REw5��pV���.��n���B�-O�v,�����,Z������D���6lƊ�r���g��uN(�x(�;*�vŌȒ��A7�#�*��I�#��mڛ��Ex�����B-�Cr�>�n�|2�
�`�޷�.����eBYp���QQ����Pq\^��n�n9�*�-����]�%v�%��3���f���"k]Yj�=��u�[�Fq�o�=*�ĸv�rY�8Y���:�q.�;B��\�X��Ί�5z��QL���Ȇn�}Kd8V��iꊍ����#�t��f�2�q����n���,�����+��f��Q�@��3o�yX�6�j	"[�a����ː㝎S;��o�a�m;�³盅\���C�צD�>�zɳP�(����Ϻ�QY�/0Ňq����Gʽ78c��VK�j���[���.mGZ;U:y�aI�y�9}����;X�R렱o8__rD�����0�-�2�ZWj�e�r����\K�bQ�J�9� h2/�ڹU.<LrŒ��Xz.�|��Y馇*�ˮ���f@%K�g���Q���qý�4t��%L�uY���R�w@�E�1��֓�.]�׶:�i^���W&\�:=��gR���^I`��w���3]l�����1�ų�(��J'4�\�r���V�=�eh+�=i�3�Hm�����Y�1ƃ��5�揸�V�p:���J-�9�p4��P�i-�%�qkm?C�.[/�������޺|�ɤ���z[��*˭��gF	d۴�Q�T�A�=km_����z�j'_f�ݪ�am�{�e�qGU�Wt�Cm�q�xm��IA����⸫�}������;s��3l�;�ͽ�ES�ķNWkԟ�!����ꗰ���m:��rUݧ/x��_-�Ҷ�ZT@M�}]�VC�F"Õ�����hX\�KlY'��
�.*
YUﱻۉ�ϹIg��1,���.'&�fr��-�̞���1�<�5�y���ά�����S�wQpQ�}G:Z�`�i�gbMu1�nkۣvnݦ3J�ġ�xJ��U��t�M�Z���p��]�{Hl���\�OU*�H�F����q�]�c(�W�R3��;�v��o�b���:aݑǥ�د���3{n���X�0��%WUs�w\L �R��N%�f���j��O�5Ҧ�d�dw"ų��
���)���j��� &��|�
hι��P�f�u����-���Y[��z��@�Q�GQT�;�����y�l=��km%�X�J����9��Hб$-ndC{���dwJ�n󺖂�5W�*s��E�VE�[�+ПTjy�ŋݳ懑J�ʞn�5�0��OZ��z�Uܽ�����cEE�֢�a}�k��]&�p*k64�+��-U͵����-?<�)�ܿK�bW)ʅ���ZS^6������)Ú�ڽ����]�Zls-���1ճ�T=�b���-�/�og"���:[����E�=�����1����|�EDN�D5�j�*����I-j�B�͉K��?5��.H���<��O{q�μW0ۗ:3M^]U&j�4�x�0�X��ʭB7S1��,�`=�oq���3�1(�W2��mm�<�7�����u�W�n��Jk[�C�_`
�s��\���N/��v�t��y���KTa�r�.`esv�3��b�{�^e����Y�ݸǦ�<�{�α�jl��)���ˡ�ִ���I:�2�*sb�53������58��
���GyH3�+Lߨ��j�����rX.�{�<�Zjf��w��Y`�j�d)�Y�i�+�Aۋε��Bv���3�f�.�=J5r��֎��ۮt<�s�:�u�B>�W;�+H*C�2�x+�\e끱�<�h��l���2o��Յ�3x�#G*�`��a���v��C���&�<���y����>bw�K#{�}7���3������.O}A�8���5�O3�^�:,m��IwG9�\f�c)��R�X5�p�c�W�kz�Ɋ���;��8�7���\�`��e�F;�����XU��_��pݸU�G�-=Z6c�:��͸瓦^l�>���dV@֠�٨��	P�|�q3�'��b�G��V.�'S[����0�Lq��
1P5*�+�m-9�w%������e98#"n�u�3�� �p߄���6��B�d۩l��D謜���°��6 {�'upE$�;d�U�����p`�m8��Sy܅��npo�����☮C�Zw)��[��WI��,�`�����0g��ܸHI1�qmZɪNl�Vk��r�w�$j8&��=�6Td�gJ�����Z��~1�.0��w)�:mo�b�ls�]{��ܞu�؊��ګ\�qz��%�c���_Sr�5�3��M5�J�"��^q&��VE�[�km*ȷ��&S�wr1��wv��,*d\.R�T�5��ĮRj��=y�Y���K���[޳Yޢ�rX�{���~R��d"�G�+�zͣVQS~���R����>���@�^=��w#t��5Q�¿7�e�Ț�a�:��W���u���SYN.�i�k��F"u����:f%��1·t�?m��%�u�T���~M��N���X*�B{����ć]��b�1��!C��Q�:��{�m{�N��6wOAcY���=P���ƕ��դp!��OnH���������<��k/0�Zu:�R�Nm�yqif���YUd�W�1VeE������<
UT������u]X�v�<��E�rvFst��i&�e+�Lp�;���Y��vg�G�j�j\;�'睘a�,	�fz����eO%��`�����J�+t�%�ah[n�,�K�{��ӂ�d�p�qt���O��I��o�<��y�\f�
�<�ƜW*���&5���wD�*�B�ڂ�l��O6�y���\%��W����d�lpN5T�ʅl�q��-t�8���N��l��MՉ��W�ђJMN�7c�H����7dz|c{��>M%n���r^�V�$�m����OnԂ��D�B>a	w�j����yvA���;�xy�{Q똣y�wj��<�C�G.Q�-]QJ�ud��ו��Wp���^�w+f��8��=�ֶN�V�\ou#��Qj�ځ�a.y��J��<�#�^3�"�����KmT�CIAc��X�@���zcv�d��坊�:�1S8�Sf#�l�v����{����M{sa���b�V�<(�\��yZw�[P.�%��Ft�aRT��� Wv��8���5y��ђGgW�|q;��s��r���d�|!�E'��v<���Z�w&9d.��X�0ý�f�Y�clk��C��=;�/{�ky�S\Q]��Q��HOG/[�x���[�g�S��]�����,߼gMt;��L�����i��>�9obًR�h~�b20]�n�2�P��Bt��M�5�ެR���y�Uxe8b�0�=~��[fEv����4(I�R曄q�V���Ӳ>�N���>ϯP?���o�
�d��uRy};�F�7j]J����1'�*�t�"�b���l覌뙾�dZ�X��lN=*Qz�G�!�d����=*{���ym{)�:��'^�͔<Xf��w��M/f��X��Tu�����9��ӱ�|�Ҟ�bП��1ۢ���W��gVi�N7}�Է�3�a�ߟW���t��y��tW���>��m ���dx���"��(��s׭q�l��/ ������=ɓ�_��_N�����=ׇ�JA�D���	�W�&FmcG)����u������p�w�(V;raڸ\e$M�e
y6|(�Wu5b�䤹]�v��b����]�K �nx�فIms��� �v�\m��E9���o��x8��ܨ��{�&�	�Ved���ԳJ�X�����%j�l��]��{,�ޭ�ۀ�1/������.�Mq*�u�r��`�p�f��˹\p|cNse��`EF�kb֭���sw���]9�E�B���\�^�w�O�[��W1Pۗqz��^]5y:�5D�4���<�"���B7S>�ՖW0b����M���Q7Q4!�C:et)1�t"���A=1:��kw:h��G�>sS�|8�/g�ѧ���!�@ά���V�,z�:0��}��`3z�jK���e!N:S�bY�g�8ǻ]��RR�O��][62��5cҔ �v֮�d�Q�.#��q5�^��i�Ӊ�n �1k��s*B˺�Ȯ��se�S�xZ�Q�F��TGrP�����pt��}R�7�**��q� (�S�q�M�iP+V�3}�Ӿ���xM2���O8+t���%b3hP���r�:\�7xŻ�0�_fQgZU:M.�W�,j~C/@���z���0թ����� w��ko:�Ը#���}��>�t4����;x��i{M�S�b���h��ЕuĊy�{O^������Q�"����_fb+o\��>����q��,���1)G,@ʚV�fP��O��9M�n�QY�:���>��Vx�%��4!�_s������h�Vqغ~o6�<��y���ȳ+�]fȩơz-l��N5�:Yxf�4'˔��<[j�A�q�b�n,gȳK\уjݎ�A���Y��r��ޥ������k���.C�ˢ�]#@���D�os��9{�u׶��FNپ|~�'=6��>U^>iC�Y�.u�o����E���~��J�TH~��j����N��3�󗵓;5O,��7u��)�G�᫚I˃9I��#/}�ڙ����[��9zh8���Wd�	g%�o��bү1�M��r����e�N��]�ϵkS����c�.]�y,�w���!�3Y�m�U/�U�+-`�U�y *�'@vVXd+����JR�hmk8���¥�.��ᯏ"@�_.�m���[�Jy���ݺ�|�q�M�K��#f��m���jK܊蹽�wV)`U�et�[C�V0k�J|����[ڲ�Y4�;)���GR�6��i�(����P��@�Q�`���r '�[K�v�s��d�޺ZG_g)yf�� ����;�Ƙ��nN�7���C>tx�zS�ZUٚ��O/�[�Or%�x���	����Sxmh��:s6�ww^(���6���gi�����z�[�D��s9`�Q`�g&�+����Έ����+#ڴ�
x�v��%M���fѨz>��,��[�����d�3M�Q�iͮ���,�v��	�&LU�HХ�K��՝�WM�"������o��������/�oV�wv�堪�
/�'�-Վ�%�yҺU�K�qj�G�IY��#.vքE:{xu�)jeo̀0��z//29���:�B^io���t9 �5�b�l]V��A^m�fٗ�D��+��[��E��;���w)V,����|{�έ���BT��cx>���8�'C��ʺ��7�5�乫�%w^X���,�B#}f�-�k�W	B�����2"�^�wEH��%��ѡ��X���G�
�'uv�[X�CT�4o$Ѯ�^�\�gm�5�!���J�,�zc
���9ٽۣn��Y�8�.4o
Q�g�g7�����s;'tks�r��s[�;5�b���	��`��C���5�r��Xv4�wV�9��J�d+�i��[PpH+v���t�_%������T�����i!������0������|��4�ĮKD����J�|r�H�*��*q��
�3��kP���ɓ�ZKi;su�3����jj���r��H�y��f��`q�|��:��$}i�r�ARI�28�@$:q˷�u��;y=�r9/���aoSW,;�A-8%��#��*��B���n�M��Cq��"5BR�W�wd�fX�Q��C�Y6.β�V�"��l[�P=�uu�3w�m�����-e[5S�бZ��˿���q�� �Ț� �̵W�˵t��`P�dR�7c��Wf���)�=��[�פwgL�}��U�'�,�C�{����2M#������_<�b-����gy�5خ�	��O+W�(
�(KQ�z���wYRgKq�.4�U��*�!B�V�+^6�a�
J?�e�� �غ��X�3���3L=\�-9r��|1�!���]m3j��ܶս$@-��u̫���E�� ���+�S�9�Z \2�j����h+V�@��[f!��n�[�2�E��s�Rܬ��s-��,�=y%�m�v)t��lQ��(Wu�J�VuV9m*C1�d
A���e�����6aY4�:��J�f�r �4(
<j�!ӲT��C�Zů�Nn`��U�8�4L�Ք2<��m;��6��t�����6Ŕ�*�,�Z+ֈ,D�+DQ��X0���lc
�5�@E�6��Ѷ���"F�k@U�PR�(�

��K�ʰDUEc�1��X�R��6ڔekKBģ(,D!i*�EB�-���D��J�֨6Ѷ�R�e"�YX���QDUej�Ҫ������VT�lX���"0Q���**�X��ETKm�խb�Ȫ�� �Jm��EAb(4��TQEJѪ�m(��"�aFDAVDF#(��F6�DF��kU"�[�B�b����5*��l�)iA���F�jQ�TQb��R%j1��DF**6�b
"����(�E��b-�(�UU-� ��DV"0Ab��j�X,E--��Tc-�QAUE-(
(���"�"+`���b�X��eX�iI |I� ��q�oL��7�r�W���%fv�����ڭ1�����[���tה�(Ֆ������A��K��;��ݸ�T�Q������:u���y^�lĤ�>�p���t;XsC=�*�oF%Dꣴ�E�1��-ب�o6�i2����}.ڐ:�s�~o7�J��=��{cF(�٧��^:{�-��NW*�+��v�CmQ2{�z5��r�\�K������Y~��V�y�
���{ʳN��V��{�+��\��5]��� �z�Aq�^�)om ]HM�o�{��]�'��є�V.W+��}x)ឭ�{�\f�
�Rjy�� i�{�4�c�t�j��C����B��|�������{�)b�W�K�W��<��A�0��ąJ��6���$��*}��4sޝ�Q5%mV�t���qđ�L��x�U��5A�ܮ,�ڸt���H��m;ݢ��w. ]GˡP��WS1iM��8�W�/;5���Oh\t��c���*଼4�^iT����2�q_�[���0���eC�ˮ0 E� o<��Z�ܚ����vwuqx~�%ɓ�����-Mͼ���Kt�S2�>�]��wB�v�ǽ|���dkF��'VNp�
�\��6��{���a����)�LK�%�k��9��ѧ� +���D�����K���s�_�I��#Nse�T���ŭ�'�"�Z�3��:�0m&ou�/�'˽ϧViȦۃ���X�G���u鳘$wF��ʺ�c���ϻu].`<���;��!��xrU���b�Ў���I�+%������ǧ�4yi
=I��\Rc���i������]U��5NW��F�㸨/�FF��b[��N��E>�G����EL�������N��(�>{�,��)9�J�ct����a"�S�:���ũl�'lZW Cnz�:�-
�P�c���L
חF�Kޕ��L����VD�z�UIՕ"u'��l��λ�ˍ�����%�d����՞w����I�O:�mL�G'�W<��{x(����^�V�H�
.l�����A�h]=1Z�P}��{T.K�:p*�����˹�d{.ƨ�r�r%}��5.v�4�Md�1o-���oG)�Z�f����Y�+��PukVͮ�*U�Z�'AY����n�9y���yeN���Z�vVbIw��H�����a�D�8.��*�K�1k��)����]Q1&��^���jY<\�i#�ౚ�5wz���7�%ہJ�aPo:�w���*V��pu#Ы�ޞ׼J̜�|��������G6�T֢�Ik���yN���.�����t./	��ݾ	f*��Mf�ľ&Q�p)�>��	�z΃'�Q�{g���E�M��᪷W�]^mk�v��t��c���I�Q�2�c�̰��F�g�̃I`3���㪈-#e�Sܗ�Nu�r�G*SPyf�����1<󹃑G�V��u��|�z�S�/��i��μW0��z�w�)yQ|���3y=�&sq�U�	ꋭWz�ŗ����{�]k�jwX��lͣ�N>v!��z_C��h�A�}���K7��25�F9��b�p��t�][������Şk�ek�T��P�,��*Vmo:��,��A��R^�j�fI���8�vuqۀ����#��t�xihL�n� 3�S7X5���\I���b�f����[���'&����ݥ�Ô��'5�-	[��BH�Sr����{�Wa�1�,�J� ��(m�d|�d]'�\��Sq��iw�{���St��r�\o��wZk;�n8K���Y�e
bZUdRWS��w�n��,�5FY^��<��:h8�%�q4⻥��c�*��)��S�}����=�����f�
SCi:��pyL�}Y��#\c��w0�#[�G4<�l�oԜ�W��toc�'��g�|v�
�P#y\�Օ��
׵%w#vj�7c]�*��(�Vk
w�R�~y�O��Y0\=�J��b��2��6�;o����мw�h)�G�b��2s�I�ڌ�t{1�څi]�y���ս�>Q��n)��Q�յ�|���7����;.||��[�i]����yf�o�r���Wȋ�ol	���/2�SqGs�0��<��~����~>��[���S�EWN'��*��ֺ�,�Jwy�Ҳ
�R��5����V�r����bU}0�x�FA٨ѳ��A`g5ArvZ4%��X=������u
k�3����\��=�V�8��8Ն�����&X�,����\[&���љ�GN�E�ÏF���h�W`�(j⮧�(�9�Cl�4�%�Z�؃]Qm�k���O!��.�GUz�B��J7�Ό7ݓi�Fr���&sqMlQ��.5��Uq;����F6�v�8�#�u����c^�;�w1Er�|��+(�ߖ��/6��.,ڨ�OO���\�[��%����·~��^!�3Y�X�U�!;�<�;��إGjj,z�V��l���)�1/n�L�rﳳ�������RG�2�73��1PR1��ְV5�sI�4����]����J�ʱs�{���G<;�JG8����Q���"�
��ƕ��vo��ݤ��N��U�MRUczhg0+��׷�2�������iPUv$�۸ղ'8����oitY�>��>��h�.;V1��§X��=sX�$��k{�k����P���}x(��}/tˌ��S�n��GW=�
��p⏜��H;���ަ�^���9R���%�PK��߼�=��^t�=�󹺦��Su����u�6��w���z�h&b	1��{�9sP�WV����ʶ|����r���3b���g$�(�;��3W?��.�)�+K��e��$�㣽k�ww郭���%�YyS�k=��ߺ��g9=�������RŔ ˓;��B�[���7�W�&���׷���6�nߣ�ᕏ�t��Xl�r;�5˻�<\@h��=�(��))���c�e6����5�֝�M��wv��*�ɩܰQ��T0�1]Lť5�1W)sѵu��:����2�c�i��<��6�y�-]QJ��W���Vj�=oF�f�Ka:/��G�V��ww��:�,N\pUx�1IjV����wut�������T�,%$�^�t��D'�ƽ��K�t�%�R[P�uԵ�RS++:�����,���}��z}Ox����T�_2�Yڗ���N'�r�"Q��o����Ъ�ҕ�z���U��΄o�����[c�ݓ�b=eTW7C_e)������*�"�]y{(w�*�t�O`�,�=,�!A��[Y]t�j��v� �ꀂ�{A�-g�zR�R=G�;��x�7j���\���cs@Q]�sG'!��K�j�H�܏��^Q�ܕ��,��W �^��b�ΥX,�;2Ԡn�-Ra����Fo�ٗ���{��]�<�P��=t5�[j⍧�;�����>�P�r��u�<�Xj�8�ȥ��ܪ��#�\p���
�^o��U��]j4� ��w�:�57A�aR�q��w!5��u�M����\nOc{�qT�y�L�=�ɾΆ�̢g3��[3���\���\��s$̩¨�X�<Ѿ;�WQ>���=�������ד>���y�@,ü���ЫT�����f^鈖sn;5�A�ι�Ж(t�>M Q�4c�gSZ����j�y��oH&^�G6����E�-��J�ALv��"4�ުڮQ;t;.��8�u�κKw�Κ����ҏ)+��z$uQ�ُ'%�s��rH]��O�;UЫ�ǥ�e�*18�s�=E�p�ngI���ZV�q/;��(����sw��GW<Q��4�G"��+��^MK7
�n�n��E���*����ȁ���Z�2th�NLT���[�������Z�Y�������<�lpv��>b�cL�c��,k�(�H���� 
��	j��ǻ�1f�f�]9�B^�xwI)M"��1�	ʹ;�;M��6�u_i0�k'�3{�n2�7ӵ)�[��ӽ��UN�(��H4&k�V��+ae�Er��~����ݘn��ߋ|���d���IK��J8}]��5\Ȅbb_9�V���.��Gwr��FAu���qGmV�Yn�i�>��Y!W�s�&����WQ��Ʋe���Vk��W7ځ�Q���aW�����49�G�,��+��g�fY�b�=�NUFA$i��~�"�b��Wt����UӸ�DS���&�&�8s�#U�U���6�/�1�ҝm8�R�<	�SS!N:��)�N��q�!;�c�E�ʲ��iP*#jW#�J��+L��^H7;<�Siz���u�t���}Q`\v��ƒ��|��L�6��_w�ۣ��~O2O����g2�<�b%�c���"񩈊��r�X�{tӷZ�������;�/9�xb��T��	�])��᩽�̸�=��F/�0�Өj9����r���%�&*�d�^
�ݸk+�n��F�[�gu�ܵ��/�vګ�gݪK\�\W)��z;{�ڮ�8�Ք�B����j�{�v�)�E:V�蔤�X�.�
�G[wp���y�ͫ��"̭Fúۊv$t�[�,��OD�q�*�?7�i-�Oo���}��w8�p�6�)�M��7wZC�F���Q=F�u�b�7��tךh��ҫ��X�W�t��Ȋx�tL�ő��l=�J]Q�ؔ_��g�
��=ׇ�ڛ�ƸI��
ų}eO4l�ٱ�p�p<ʚ��W��Z�U�vz�&�#g3sR�:�Ԕ��ȭδY��ҡ����~���N��+@�ӗ�9I��W��ў�9ܖWr����p��!>�y~+X0�-{a۩�%��ؽ�j.�	�� 6�wWMک���1[+���_��3���<b&��DFۛ���7�}��,!L�Q��P������iR1(���G-=������[��i��R�nT���\�0D]�X���i3䤴ŲI�MD(���^���V��b[N�qg����x��`��'=�)ޱJ?	j���ʕ��a��WC�;O�*d�h���9�E�.�m�$Z8��r�q=[9Fһ�Y�x\������Y|_L��A�vd`T���>n)7��93z1|��������%qڰ�o��P�c`V<�6�!���m(f����/\g2��Z�O.�oY�c�5�ō{qZ���ńaL(�n�`(�8��N�EVp"Wo\�הai�F�ɧ~�ڗ�+5����T1�赍��]@_�v:�7��j�{��B�myo��_�6G��+��d�-V=W!|�_}�W��.�U��-�R�|���ޅ<�6���]m��j���I��&����Fu����TX�1�ɟ����u��H{9���!��N�H��Ξ��}��W��T�m������-��9�ܜ��ٍ�<���K�b'T�8aW���S���m�B�O[�}ы���s�6���65dC�[売�ꇶ�JI�F����z�<��G�s[�I�_Zk<�f8n�s}�ݰ���U��C�o���1۱o.�I���1��®O���.C�;T��t2T׌gU�d,P�(,*a�SU�:u 2U���*�=�7FYE�x0|���eH����;�x5�Z��RT*7w��u�ùÕ�y�HJ�Y��v�}6� Bx��"�;R�i+8Srrn�o{�<�݋�7��N�f�7��Ż�~��UAi��:�W:k�����v��;V�gj�8����\(�|t�^�S��b����Z���ԙ	U��)Ƕ�9�cn�닅���`���WZnf��$ ��V��㻷B�"#f��w���0=�k��GEҰ�zؾ�NC{hEvU5@��N��c�<v�v����SĖ�Zh���}�������d���ER��.j�rQ9(���i�ȉf��W��R�U�VtT[M�	�H�Ŏ�ʝ�5i�e��(#��H*Σ�,��XݼU�E��,�Ah�S>�ô�1��]�����G
f��v=* s�^"�t�E�i�Z����K{t��C�a�hT�&�3�ɻ�L@F]qi)��}�y]S%��g����NI�l�P���]�o9��ug]3�����破Xt9h������x�tz���3�<� �w�;�kL��%�u�ϰw5�PJ�����݂��SO>�Gu&K ����I6�R�-���ϰ��p�t���]0]����T��-��yhgeI�����	�.k��β��ֵC��5�eD
�FV�x�hP��[:9S*R@Ngo\U���)Na��S��vw�c�
�*r/>�1�)l�J�5���-K�N>crUξ��>�J�咕u�<-^�������cul70bssf9׋���.��h������V^3ViH��^{9e��U7\��h�-T��E�YTU@�U�e����V��8�J	k�/Y�)q��M!>Ղ�V`�k�3ܝD̮��;<�B�"Hm�4���R):�D�7yW��'V�:���&w[v�$wjc���ln���ۥمEͭ(�b+�&s&1�.Ѽ�q�L��&�p(hA�d�.gn����
GW���a�g�-#�/������J�J��є�M��\��ӈ��aa�:��#R@��+M�ۭw��+6��B�J�Er�*h�p�p�Х�N���k)�[vK�� (�T�mg[����L����C��h���cb���(���[���P��e�=S���������<��n��7����<8:p�s�]�����PH��6��:!�<Gm�Z�j����9J+K��|̘�Jsg�D �E�r�]ЗP��+���wn�𦐝'q�R"M`VT1Ƴu��ѹن�D4՛{�[kBT:�x�I�.3S���WX[�NPNg1�i��ӛ-�Etxg�������AU�b"��EEDQA��
*"*����"*��DE�m��DcF*�U�b*�(��*ʒ�AcƵDQb����b�YA-�ĭUV(##(�1�E"��
Ȃ�
0DQUUPAE�%�U"���DPUEQTb�UUF1D�TUX�EDQ��T����Ŋ��V0`�$b�1����ȱUYm�2* ��*(���#������QPDQU����F#"�Ԩ����b��U�0�k
�*����DF*�TVҢ� �� �m�EUb�X1PUb�EAUPb1Db"DQEUb�X����Q��*���*�AR*��b���*�(���V���"��(�Db��Q��F1V1��TcTPX�QF(�DEUR�UTTZ�@ �B�
�
}{z����vv,<���V9��)w9�M+��F�pd�m���_)���<�fO�6gY�6�oB砮�7S�;�;d���L��N0td<�D/�2c�{���	�={9��`���<�WQ"Eݷ�yҢ�WUx�CV��ϣ�V\I����y��7W��Ԯ���=��$��t�+��n��1���N�ˈ����Xy�q�R3���v�V��g�q[i�Ge9�����X�!����ԯ'�q�<�,/�^U�UN��E�I��p��G�"��|+m\EN�cw!=��܈M-�d�q�8I�eTr��	�] W{R���]P��-v=��)��xZ�^�Z*4���r���cgo��w�*݋ѝ�W�G^�VN�٧ܼ�n�z�m���q�j�ͧ
��N���0�����q�X�iS��5U����ʒ+ؐ&z����q�Y��/y^��cɐ�ӭz\���:���NF��c^�>[��7;J����[�`M�"^Ux]ͧ�(�w$�u�Q�/hf�h�gSZ�U���q=�dlrӯWe�ݩ3�*�m��{�\���f��x>���.���ɯ�����4k�^q�[��Gy�z���ơ�n��q;�@����gmip^lK�G+/�2T@ެ�zy�0.zd>����蓪���H��{�%ہGӭB�ɬM�1�3:�^&씬\����t�h�t�j�����R�Z(�&2PW�+U�;���U�9��R�馞�$ӻ�|�8�%�v���ض�j-Q͂�l6v�z�k�A/:�ù\p|q��[v�<�d*J�����.�OC�Kt�z��H��W�>����S����ɦ�&��@�J�lb�=j��ݩ�l�$����&sq]Qn���W���E��O3�t8���)�Gw��!�,��7�B2���R�W!�3Y~F�4{�-�}Y��(̀\�/�u��sfmLM-t�k�})S�Dx]����x��u�2��m'ˋ<�bQ�p��Ґ�5��R�.���2o��yr٧�OB��W����niEGt�|�cr5 k��3MkX��:9�]˔;�q�o^:$�۸���4ԓ$�qמFU�^a5��0�� ���wڳ�U�mv_j,��v��]'�.[E۹���d���G3�9�H�;8+F�i������@12��EVt�g�Q�oqrf��y��h��%��u��b�V��R�om&iW\��v�W ����xb��i�R�\����"��@f.ݩ��N������I�G+��	�4��#Ini�3�K>}O5�M�:\�l�}[�8q[��P�͜C�����[K�}�{ƒ��	���m 6ž-��Z9]\*�W�'����e<��0��;J�)�՝�q*������魸�U
ڻ�ټ�{�,�V���S�]k{c�����O|cR��[�(elդ�����ZWp����+z��hd�����=�z\+�e[�{%��θ�W���$a�/�����������W+*���9�r���Џ�BC��<Wv�O}<k��0<O[��Ǟ���R��vv'�rY�Jj�*�}���q���&-r�{�����ġ��N�%�x��I�i�޼��ht�����sq_���7�S����yK�Ϫ燚"Y�r5�c*T��L�ג<%t�t�mZ㙩�i!Wѩ���C+S������OB�ceʐ���%evN\��XWu+�x�NW���;��8T35r����G1]v0��f�c����}R�����2���V����"�|Uxs����n���}��l<��UC���Q3n�4W����t��pF
��E���}{r�����3/n�j���%AO��É�nb��೓����N����� W��������XO|Id�>��Vʩ�L��Čv(�p��j�z0�Q3T��D⍣�kW��a*��G��������pq����
�y���g[9:�+�z��(���(���u���^�3ҍ�/ն��O���L���=�ڏ���2�����9ޤ.P���J�w�O
ח#�K��b��:m�a�����:�m�9��R�+yw�������&�U	U��+rs.x���x{�~��3�s&���$ߞr�eW��tˋ��p.w�s=�I	��t�'uoCL�n��w)yMv!���8N��S��<�ڜ��U��m�9`�ޝv��B�=w/l�W#kH�l
�i-�NM��i�-�\�A����z��YupԢ� bwu����G�GM���:��Qo�M���?��9���7�w����9m��n����V}�];m_��jx�m���(_hE�t.���[�}��'���h1�N���et)ȨY�׊R��C���}�oA8��32�Ip��hW������o&�W<���h
I��k(�Q2򷴚��d�H����L���ns���}9px)# l��˷��9;]f�[��N⌺ט�8���6=]���̋��s}6naH�Z��6w��bn
���꒗�z�:�Φc�V_�$�����+��U�S�f�E���j��ÔX�&0n;��GT]'GJ�-���֪a�7��]��6����C.)�Bd#a�1T}q��d��A��̡�x[y㯰,j�}5�R��T⢚��CK�C|+m\Q���3�wV��Z���\�f�Wt�@դp+�CU��שŪ=^�!�M������Oy�\*��.�LN\!7�3�m��܆���L���In�W�۞���b'�	�>�X6�����']��d�
��ϓ���.6˄�6�}rT3���B����Ċ��>95��w+;
�]X��y�NYmɜ��嶕��.�k��/r+��l���Tg`�ip+���&�<�l�W�V�9cR��}��8��ң0�ͳ�e�0�w�N�,�'�P���ܺ��vF�������M;{�\fN#�x���v3����i��N���=CSX�&��˯kޑG�v����V/:�w^֔4�V��E���4{1­�W�n����k���7D=�(�߅��Ee�-�}Sz a��G����}.�{�T&�ۤ�q�a�;� >��(��U����7��\��s�N���5m�W+� [��lft<XaWN,��t֞���]��9�u�9�ꈶ������hw+��`�zd�T����$\�f�q5Ztl�pp�˃�7޷p-#��6��N��yuZ/b��+WY���o	��ڜxՈ�n�������z��<���Ţ����/�mX�{�FQ���$�セ���
���u�14�xp������̡^Ӛ+׵��k(�n0�h��ZX�5��X��h ���
������ 2S�5��Z�4U<�+3)��/6
wpi��ND��l<Ȍ��:7�Q�|�q&I��BNK�[�������xי5�p���ug'J��_E鑠"�y������V�frs��i+9����i6X˄ߕ`rVq4����ՅU��s�)`��/V����!3ܖ1/b^ĵ nC
x�����]j���Œ{�Ғ⓺c���z�ԫt{���+��b���:�4�Q�gz����WT7�\|����Ֆ�-�-�:>��	���1�:���p�͜KUWA�%ìο F���;���k,g����2
�����v�w�
r�^��7��f��;�����위s)3xTN� \	�Ό�#)�+V	��@*ə�	GaT�:�I��m���OpwD���q�F;��Q{�T�<*�B��U�k4rVՠ�61=��Ռ9�%���-�=}����a�K�"�k����<Z��n8��=��g��ژY�~�5��i,�u�Vm�u��#���Z��yv���[F�]
�U��^�P�6�����ݺ���\Z��{s	�����2���C.ɏ�'�9j�n!#�7���=�Wsi���B�s5������2mvumbX�2���㛴��Nk��h$��uH���<��Q]����+��ܧ�Y�ΐ�H��h�߳;�<���O]8�%�2��P��ut����^��|�l�n���}����-e�]�:��\�c8��]*�T_E�TR�]^�l��[�n���Q�Ei(�B<�4��w����E�N\��LNn+��֘��z+j��7g5�*}9��XL$ٽՖV�S�}�g㹊�IAc�䪹xj��+�u�Ņ��=AO)���cS��זWX1�>}��nB�e��F�]^O@˖�ڸ��G�m�N��:�\B�Ϣ�=�nz��ǜ���>d#�
Tu�+-\
�L�V7��L�#�PVyڢ��ɪ|�:�UXW���15��c�E^�1k9ٴ���Q�S�(u���Xj�8�r)vP��h�Ph}v"��~f���H� k!Z�*)z&N!��T9l��\���R�3�W���r2�E���Y<�ۭcƇ�Q��V�?IK���p���/".�(�#b�kV�z�s&$����:��뒣\��2�r=(XǦ�Q��7�$�D��	�6EIj����\�M:r�ԝ�k��梥�������3s��G�u]=Vꛈ�!�W���QL�r�k��8�!��<:���v�,x���V���g�kd��S�}����uf#���7	[���82`�ʰ+��[���������N��"_�D�2�VɕѻEp�cL{�ʺ����zzNv����%�ۭ��ѷNV_ն�p�C���_d��D���.������f���gT	�M�ti�_Q}��Y�����\3M�č�Z+'�S����=�t�*��Fp��(c̓���cF�����r��e�f�v��#m/>��;)[������爕5��K-t��̩�4�-�*b�:�f:�B�/"�Y��7�M�u�8��%
���ݲ6�<%Ҽ�.�(��s��Z*napS�t�V �˕�:{I�_�6�dK�Ĥ�'�y�����{����q� �A��'ڇ�3�x��z}=4j2���4d?h��U�W.�%ժQ���ʉ�~j�TM�2��ׂ�)���:�.�ၜ]�+M`�R��5��5��ovy��L�5U-�tZ�6@z����+-�9�':y7ސ<�x<��͹�����B�X��a��Ҡ_n�����zیA ��C��YY�^�=�����H��]Ɩ���u�9�`O��N�軣�w������g6�.��Qz���`t64}��\��^:�·<��E���w��Ю!�m��
���+5ڬRH� ȕ�K�Uq4�&jcl9���.M�v49�-��;Z��|ymA|�<�x��՜v϶����+ܥV�P{�UT�t�����
��4�X'����]�:6ٸ������������J���Ds��횕�2!Z(������ך*�V�gϝ���~A'��U#cpϋUYc��^�'0�^*�\u��J������{P����t){%�%�|>ZU�uq*�,X��o�5i������%w.o�d����T:�$�������
�$��o�6�ɪ����Պ��WƟ��~���eD�e��v'�]���ų���iݻ]ʳL����Q~�d-�/��=�Tf�eB�62{
rP��ܑȶ�ڊ}	P3)4�L6)�)v����l��eW�P:x6S��}���e��}v�N�[$�/.��{�M�J�!�J���O`�γ��H��Ț�}�{�I��$�	'��$�	'�@�$���$��$�	'��$ I?���$��$�	'���$��H@��	!I��IN@�$���$��$ I?�	!I��IO�H@�hB����	!I�$�	'�$�	'��PVI��k�~ 5.` ��������_/�ڀ�Mj� � �-� �R)T�T
��`�(P�A@ �
eR����Z
-�h0hh��N���)ED"j���[�IUMjR�����	"�`J����ک���z�����6-�PK��v�uc�6���X��1$/�i�HG�P'eaT�g$"魬Q��j�͕P��WjŖ�m*kSf%tҔ))�
Vm)ED+mR��ڮ���UP�4�  �U�J��6��2�����0�-h�psm]ή덬�3�-�:�K�\���v��n�Z�P�n�m�e܃�gj��J��:˘ӷt�w��Ί��j���  >  ��}tʵ��n��ӥ���Ԙ���v떭�]���im���Q�75�fہ�.�J�fq��TnwW7(9mժ��n�vU6�39;��a+g^��(�!An�(�Y
ў�  s�vj6�ۻ�0�m�N��뭳��56��m�u�m5��0-�v�r�]݆����]����s���܀(ov�
4�C��קx� �B�����	
(P�B���J��`   <  1�(P�B�
({v[� (P�B�(ZE�
(Pp�	\��Ֆ�5����8�u�ڙ�VB]�m �V�����jV�]�9J!&����  � ϼ�EI�ݙ;5l�$�v�mZ�gKn�u����m���e���µ�R�c����n�qT��Ն�*��eMh�j�QIJ�{U=k۾  Ύ7ں
MU��v:��;U5v1�UgC�v���e��f�Е�k\����δ�dS��-]3ZP�5�����   �   �{o��H����۪�gU�A��q�V���֚�����p
�DջU7A���ݶ�S5պw1�l��n����ʺ敻����e)�^M�B��ʉ+X����   s��+�۝�n/m��ݗsȝMX۹w��z��ۭڻ��v�gI�6����vʥv���֓J]I+]ݗm�Ms�����ts
Z��]]�%b@�/Z)�  �   n{�u�vn���Vk�
�v�仭���@�Ү�Q��N#���vӭYW�k]�v�]��[��ݚ츢�]��3�]˵�w6�N-ݜ�ܮ��� kTa�V   �   ��_Uu�v��wnݖ�ѣw���&���we��ڥ���Muu��5pZ�e��v�u�)��4.�Ɵs���P��.u���r֥s7k[wn�7�O@2��  h��$�* �S��T�� �JUOF�  E?
a��M `�M$D�T����������_��>�
�W�6l��͜�:�X��PX�	�Iq�و2QD���q�&?�H@�f��R��B��! ����IO�$ I7���$�@=��Ͽ?�����tk*,�E���Y��C��&{ޏK-e�b��=|��D^�
��b��Z��zN�p�{x�h�O��װ=���7�)нQϔԎ��e'pmd��%�OE{z����V�+�Z#����ub?a|��K^�%�1�%#>�;f�5Hm6��Y��[C^ՍA幦ѻ�̗�1�@�Yw��Zv�:2Wx�8�_��c �����U���+�q;����X����E�����m�������=z!Ǳ���5���]�O(�%�r�~:��8/;�}���*>������]4�K� ���઎{,�{༝��o��K�ߵ;�[�s=��V����'0�z��"��ȴ_ad�/"2������@V�Ay�VMc��6�!��:ú�Y��J�kq��������˅g�e�9�??2�>ew#�K͙ǎ��%��0u�x�zK/&���F~��z��wA5_A�j�������H=���i��5�f��4\U�H��@5�.�&�<z��X�P�n�s8��x��z{��!��k�j�D��@ꔡp+nk��l�5�8��f���`\4tּ�\���xw�Ep`����H��� ����e�t7*Q��L���F��W|)yڻ�ȝ��DJ��h3�]E���v"�˒c��{��x�_��ț0��$�W=c�՞q�U'<]X��ރzڹ�Ǹ�x�y�{b�|�:k�����4ؚ� zk���uv���3jT-R�N8M��t�]m���@���gY<!�;PXI@JFee���C�WRJ�(PD��W+n������
Hâ2L7�SB�fz����Ml��5G-�2>p�3� A��"��.�����(�<�VJ{X��VL<ŌM�O#���<�ρh�T���=|�Ng�ߓ? �w��{�H���M���C���q�P7�l��p�� skcl�DA�g���^ݭ=�	�Y���##)�?:��%]��d�:%��胰�p|�ہ�,i����s�y^���B�R��v
���7��oo9Z	�&�ý���Xz�F^6M6��)�gǽyB#�/�"�{zZ=����,�w�ʤ���z��/8]i%A� dŗ��߷M�^f?��#9��~<�E�*>��[��ѤTe� �/ �z8~�@o���Q���/��C@���'�:*�o�g	�yܺi�=����9����~�: ��e�����x��v��*������n���=�1ǲ����ǆ��'��>=~��s
��
�(ֻ�FsЈr�!`섡DJ�i��2`�C[t�`YZ��KI�nh�z`L��kΦ{t�!s�^nm.(��6t��s�_x�r$������\P��|�*���ʽ*G7[�aU�g֋�mlGV�-�o�EǤ��u���+1g(�d{��0۠X�Z�CN��QQ��f��4�Z��3�@/VS��ˍ�>�z|��SYP��V���xw%-��J��t} �Z��
���4�����t�L�CN���>��Z��[��1�{�;���.�;t�m��3�X"<�Z���Hûow%:�&�����
fx���v����˸'���ן� �ard	�MҴ'��o2ܫr.N�|up,e�9,���k3���7���i(�����s~�����=}�Vw�\��(�}Ob�[�s�97�{��<�N<�P���Z��1�ȓ1����|z�/o�htɢ�!���`�s��c��5�k�^�v�*�%q�۪�ԛn�$�����8^+YM,=�]�8�<�1��_Ȼ�y�h=���v��Tǂ��C�U�z��`s;�:�m���N<�VHj���-�g�򞻒�K��Q��=����D�'�Ʃ}X�v�/JJP��DG�>��'��Q�w�&�Ө��s+z�6��;Q8{w�sR�{�'� r��Jl�������/!����1��j8�/��L����-RE@�,��n$Q�!N��8�l�Ȯ���R)�5S�)���3̉�"���7<����-זu�z �V9��|��[���g��a���.�\o1Ȯ���#y�@��_1��������`�%��J�Ŵ݉pf��zu�cpI:돝U�m� ��*=�T������Op�t^�E����aY=XϽe!x2���y���ܐ`�����I8K��^~�J�G�Qy]4H�q�C*�V�[P�hG�a��m��b�� �S������ާ��z�O��L_;���^�U��:����w���1�ǈ�$��r=}�5{i�d�_{�<"�Fjӧ����Ry)�2�F=:y�5���W(�I=�J�E��;N�6�K���%`c#]���ü', Ʉ��xz��^�?s��۪��(��ش2�5�Λ>+��
V ��T?��d�A^���ox�yt�^��r��pG�v7�:������Iޤ�G������H�%凔k���O��z�9n���!<lޞ3��.F�͜�h0�C@�3U���.C�v��}-��g�E_ �#���,ͮ<���l���i��{6T�d�{Q�g�և׷o���a�&~� ��gѧ�O�8��KT���͚z��t�S��9g��e O�{N۳��9��3{��P����^���	�=��m= ��`r�hP˦���6D��5�w��žZ_�1L���aS&j�j�aQ��Zzm<��B ���6�.����y�m��e�z���H3(يJB�7N�.�&���|���ذ�C�[*1��X�?F�,m�5�����Q�V2d����=�"���\R�OaXr�n���^w��^!���B������V��2�����O���`}�3�t�w�3��*x��/�G����I�	~r��=������:�?w�,���S�PN��v���p7\�׫��Ѕ��|o\y��~ܦ��t�:x\�H�V�h�7��Qq�.V�L,
h�1L��3fm\�e]]WA&�^���~�j!����$ó������3�1dI>�-������#K�D`�f��;�k�PvInFQM�?Du��MG/&+�v��^���u1�9��p=M��"xɡ�:ű�z��p��'�gK�{���o4*s�������#�ٓý=��^�d5�LW�m�u/�7�)�c�w�����SG�+=�����2f��>�����TuP�d
�z�\��.켩�r�L�\ۧ����g^i�{�p�(�P�4�����J�DӁ�em�F�w�*���ӒG����	�Fg�k1����d�ãǓn���*�A�m�Ե���h�b�^���1�n8�~�N��^�}����0B����{®�N�z2z�W�x`�见��ӯW��Ø���(���¡��myO(M��K�a��#���I���!�8�"f�?V�{�����QgZP��.�����4~�R���=��OQ����0�Ix�v<{��ly5�>Z��\��'Gzc�y��_H��K��o<Y�մ��F�&�4�lB!4n$�Vf��(4�+L0��0�.̙��ڣ)1� <]�����M����cR���\��r�%��"^����S�ϑ�y�7/��.�|�bB<�P������� �}�Ν�,��P�'gK�p(�c��{��R㤧?����"u�}��e_sa���o��[#��<
���r��|N��3*�����r�B0Gy�L��x'�4 (�ڟ=7��O��r��c'�|�?9����g
�MA���q^:>��vF8��79煡ι��mֿ1p�ؕ�� [-N��+ۘ:���k�p�����7m�W#,�@�L�q��	�R�%C��;s7�"�������<N;ooZ��}��0ʓ���\�ǯX7E�Ǐ����31U� 8��mO�>��lQ��±�y�`���{���|�Q9yuu��<��
�G�+��咰�%�����=�8�,{2��K][��i���d�sg��q]�8��Z�:ޜ*Z���b�S/o�k����;>��b%,| e��T,��5/ky��@�zQ
b�Thq<�S�
�uz���n:g�{�ш�/�2n��z'\���Oݶ��](����0�����"u�מ3��-���d�
r��u�]8�v�J�Ig��Y�W��S�������g(�;f܎�)�'AMk*���N9Q��^�z-�=���ov�����PE��-��T�{�K�z�oƀ��w�y$���;��,_N�j�}�%\Ú{�:��<���[P+�_�����炖��"шg�H�� �PD޼���~V��~���8��|9�&����^���oO[jjE ����X���R�V+Vem߯�<|ϻj�C�b��7�	[��5�|L����_�@���>`�7���n�-�Ǒt\����c���7*̜F���s�6u��#Y�w=�� �P�B`
�՛�z��YR�*,i�l�(�fޓP��)>�><p3T�\n>��=T8�^��F�ӸY�-�`9���s��fawq�t��TpX�c�Q�s��5�_���{d7j��0ن��i	��4�k1TX)�Y�)S�[a�j�á�k�$�v�z�����^��Le���A��iSp%nO�Ү�@�]��e�NQ>��z����%}���7���/��E�@Bݭ��K�3�,V>���'�Z��q)�q�q^P�r���SP��e2�3te5q���s��RhL���Ѿ��*t�\�0�"#;ɸ��iMn�0ݚ`V�=�Ù��KB����$^��X�P�6k<��O?,M{u��^���5��y�����Q���gY�{ohb8B��l���
�J�hJ7*��۟An<�@Hmy��Q9x>���#;��ڋ���N�8U�^<�J���S�[��	�ĝ�}F	B�����k�%"��nZ2���)=<3��3{����F���8{,�s�WLi*9��كSVְ��*�c����wz����m��)e���=����!|KɻW�3�=Q�����	�d�{JC�,���*�� ��0J�4�`5�K��m�r�Ⱥ�Y7*��*͛�֕C��/�� ���Xz!Le��0�in/)p�z@�=�᐀A��VL�x/z��Oy��fC��0�r��kP�f*9� I��m�	�~���~|C�<x+�̵e�Io���s{mi愮�
���4�O�ka��.�wG����v���<�SôQy�}���[��pٵ,Ս/`���H���{�^�w��g�Hk���^~%N�)�ό$�Ի���k�,�A��z�����C�ƌ2�2}�9r�:�(�'����
$ӗ��f%}7�!<NI�D�(�^\5�ܩD��b"��z"��
H�زP��;7�������;O*݌�)Kr"��R���L:��?)�<_e��8s�ޕz��v��HJzjҙ�SThaߣ�������40W\[Bӡt�
�c+r����8�W.�h"ͪN�W�*L�kD4V-�}�wi=�_g�K��Ay���D��%)�*�I:XR$;�U{�����Ax��#7�l9�ѹ��%5�8 ϕ�/I��,��Os:L�x\��֩�a!K9��_O��� �o����r>\Tc�>���܆�$�k��2�+��?y�_�v`([`�P�R�-���a=�'�aة��ǳ�u�_�}�{{~'�j7�ry��q>�������	�_{����&U��2����H^��U���Qԫ�,�����O���9�H�vM�n� Y��@�n�09\�ДZumkhfCX)Rk�p�s�ڳ�5�z��x/N
�2��}�֖}r�,�2Mw�!,=�G�]+��j=t���������τ5�oK�����uN�Z�����S �IQ����I١�n�aT��@�'��/�ُu�X[�x` ß:6�3<=ާ�ÞД=�Ol5×&<�{E�������/�Υ_#��y�������fG�H���5��"��d�GP=H��K9�m���Eg�HR�Lw����b��&ZV��^� E�i�R|ۄ֯��,��_|�O��x��Y�Qst{�O{!�$�p���ѥ⍘-N]�{�Y�xoY�w>"�:p�����Gt{棇t��Ţ �~�1Y���7�ND4��+<x�t�MH�n]7D��ԫkl,W�5W���Q��D� ����$r{�ğN]�}�
��݅�*lB=��`��U][�8	� JK�!�$R򛌅�������HՋ:�(օu��|jI{e�
��揷�4hw94�g�`97|����Y!V"˴]f79�g�܄�
����'0'5�[sjl���Z^*�4��cU�Zvf��fj.�~�WǮ��yW�k�Ώ����J��:�g��i=8ySz7�s�ԕ�}%���x^�`2���8okM�j{!�}�����o�HRWy?f��R��h����|�+��xŘ��m���x^����O��N\$�2їo�3!x3���G�X��J���ز�"�e+�:Y��Æ&��Fwmq�̢�;��i�Xem��)�i4�\�U�7E��y��M�ԙ$ɜn��=�����;1���zd�F����|�s��L�����=IfȺ�Q
&��./{�U�}��ѷ�Ww�Qҥ�2n�㻭� ����dY���ۭ�K�P�w����چ�B�oe*5�M�b�ħG��X�2�u�V�y�Y�����w�A��jn�=�ՓX�}�N�\�k���-�wl��
��� ��O���Qݙ���|'ڎ!�w@v�Ϯ���Gt�Ь�&�jĝ�t}��^�F
�O�A���s���B�IQ�\�cW˱M��%�k7}��J��v���mp������#�5DAbi�K�<�Rԥ�<	��q�N�e���W�Ӯ�_Gq7��:5�7�T� �˩�����t"X,��Q?(���j���d��*��{txv�S����}����BU��X,��M�e����<ڃ��ф����[�S&��F꒰��� ATk�t���g-�|��LPoX�5�.���i�1b�X6n:n�:�W��Ʋ���'�(��N�]J���"O3����l��Y�����&m�H
i6*¬7�l��L��K�7M3�v�6�WF\��2�MM.�ͳ���U��f^�E��8�r=욤ᷖ��D�\��J\��Μ�m\���"G�3��eL��VJ��p�Xw�F"���}�:.�bdc�˯���PU�N����/l9��f�gh@���:C�'AK��m_`��^��:��z�L�P)=k^<n����z�)Q�o^�V�F��0h�e�\Wי�q�H
�R)F�L�6�h�)_q�+��8z%��,�|Ԑ�ݫ\��[k����7I(!��i�N��屪��Ƿ��iW�s9�v�kZNUꥈn�m������GL�B�3x�`,rX�']m�lH2�O�l-��h����*;��-����u���-��:؝����Ջ�)���D�mZ�յ���c�V�b��)d�M�r��;�Pp�n�T��u�J���yP��n��H�Ej.n�o]�W]Z�9N���<�'b�5�S��wS�q���q��ICO-âZE��QL���f��3�u9sԯ��</s;�%�55��4���]���	�^�?*y�U74\�5��3a��3\�GQᇦw`�E��[�i9X�;�vZ�8^�L�&t����ʲ񣖨@�b:�����0�v2ؗ��Քslr4N�}�F�wR�F܁d���Ero�OP����:\��&en%L_9})�;j<UY�Q�l'�Ԭ;����Th�e�\J(�f�A���
�m�)|6��s� \��GZ�9y\�L�)\�粸e�n�າ��0���s�Bvj�Bx�c��BZ��+[�����$1f�f�}*��W���E�tn![���"�e��H�4.����Q��V3if���;�L��ʟ�P��g�����w�sqJ0�+.�J��X�θ�n���Ę!���-�@��bv�ZKu5-Ӕ΋N��U��"�����U�T�Z���܆TL��	��y�G��[���f}|i��ok�	� ���L���oT��m�����[yᎬEȌ��Y��+LVt_�w_u&�\��^����Lć>�r��v�΄;����9�Bt��2�Ma�CUvh1�?�m��
T�Zn���⍱<#�}�= ���D�6�W���R�ny�ɧ��!;��y�L@�$�o�jd��"���6�B�+��7�QJ�`ّcC��S��J�Ȫ,c��yBã�;��n!ԫ%	+ivZjx�2�AV�� V4N ���;�^����� vwf��pQ�-����h��'i8n��ǆ;��Y�96��ٍ1�_k�G�2km������|���}�B�Y��U�.�I*=t��a�#�>�k�h��*@b��7We��w:��4h�S���w�.]���zwZ���_4������:Kj�\۳Q9�b��Χ�b����S52�.����޸��;�A��	�k�릵��T���)�	cH-��\��L} �}}X�����L�o�kz�N^��������K
�6�q��"����h
wW7�fq�6�E׻oXu"�������ui-)��VO��U�.U�9��YGi�x��$�w����r���(/6n\��yH3
�����Lh
E5�{�T�������Wmb�%z�؆j�y�M�\-%��%��k�9�[j��p�d�!_d���NA��Q�qm�]_Z�Qb�O�a��&s���3��롭��R�b��}���*��z�g(��eBf��.�$�wY	�5�!%A��m5i��^���eJ��,X2:u���92���(��8�5v�Х]������߸�|�͋m��}}ot)ލu�ƺ���"��ۃ�U���,s���t�ZcB���G�tǴ�h�Rތ̓�չñ���H�@�ɮ�ڼ!�|s(>��nS��Bdܶ��n�
b���ۦW���q�m�y�U��TIH����v�Eb᷸+��7�	:�N���5I�m�qx��L����z�j��O;H���K(�������+���j0 ��+U�@����V.��>�.˶���*>L!�.��ξb�#��l�:�^e<��l�xy������E�ū��Q�9J�X���N����v9�{�� ���ծ�bu1���h�D�9�D�kF�N��W����;���sZTۼ�SZ���B���h�џ"�7�&]zj�=�!R�]ས��po��w
Əf��Zr�"�=t�<�/�k�5�M?y���Z�x�"��+t�de��.����̈�-E�-���X�gbT�fɛQXKT={�+2相��<�5,Q��>�|HP�o����,����^�D���A�rHu@1���o>��0���[xs#�-�5�B�ewL�:�PL�W�y,�b�w

r�#�8W^D`��F�W'*t�y�D4���MX���۔��S���[�(�w1V�̋�7zx�dꋹ\ee�+�;G8X1�X��ɰ�t3����y����+��:h��yt�V���'arܹ�I�wsgb6���ok9�]��u�K����"���!�ڨ-��\��Ƌ��/���K쬥����WH.����z7f�P⮏*x�Uic{K��^@�V�dB������"ѱ9V����K��|�ihv�u/�P��{mɹdX�S3!�����BC�l�I�{���$t�]s�auE�ԯs��i����s�7X��,��k^/�u6ee�3���Z��w:0Խ�#��oo@�y��F�����Ak��",;���	���Pڃ]��3�Ԧ�ϗ� ��c{��՘��o��)>��v�gߖ�;Z�NJ�����:���⵩�Y#���Mm���ݤ�@r�]i����E�5/,�>�OP�����h���ز��³���H���Ǔ�kl�72��H���N eF��H
����c�J�+7u�1k=���`ʔ�#�C��,f��ˁ��A�)�n���s8No�o%L�Q�LɏF��w.
�x�E��y;g�	����v����0d���sm=�[S7��P홸sX�k4�}G{8-��W�Āׯ���yP���T�2�x���mF��)���X#���Tj�;���p���E���E˾��Ab���e��Ҳ���d��ׯCy\����A���k8ܐ��ֽ��M�Z���WL
�OdT2I�q�]�V+��˚�jZ�]֥R�ʍ�P�Ӵ���\�₧�PP��4ŉ��ٿ��'	1LǦou��ڭ%m�sST���#08�V�Ʊ�5R��8lTz�/GAtZwז��.�z�n���ük���᧤�����
kt��^M����u�e�l,����V��px�:�Y���@S�+��*�%>�x�#:�d�� h�h."�
w�A�u���D9��۳�w�[�BC����x�v�N�c�A�j�
��N���p�I��ۭ)��8�	��c��]]�;x9��t�,U�]�A~����2��i*ʨ������Y�{����nU��;P�+�ǭ9�m�ά#y�K�j�땗f|�*.7N�Fdؙ�	]2A�V�
���,*����.� ��N�)nιPP�c�&˸��v�, @�5��H���g&�lǯ;��uM�&�n՗��R�p�:��|��̋�����Аd�+�5�θ�kF�t�)Tk&�+����ic�Z�v��=\����QN�"�0�QP�1��(kq��e�{Sg\}���A�5Y�y�f#�k���J��Jz�s�3����ɋ�}q��s�P5F�=\p
���$��8��Ωق=��=zyF�0�h�`�a�N#2LT��c,])P:���[�^U��T��Y��hط��VY�N�k�*����*ő;���R
��[�M���:�|;_�s�E�F�3�A[��gG��N�p�!F�3�*]�$8^Ԙ_j���ք;�6�U��.&�����3�m���f�n�f�H�������ޮ9R+��;(��T��{�aD�����Q8���Vi�S�B��|c˫��;��::�I��9���k�Y/��Q7��Z�tWq\��"�k��6>��y��ܽ�2�I��n��p�0`�YO�?qZiԫ���}ڑ� ��\�+���qF$���]�[���{����E�z@k��;�јC���/L�Q�u��a���wU�!�\��٣�e&�p��ɰ�\��	�d�u|8��w���R��C���v[a�0��b��+7�X�[ݨY�]b��æ<8�����9�q>_k}�'��#�J9��x@-y�1�>3�>��tܡe�:��&T޴v��G5es��KkS��F4Vѻ��&D:u\�0>�Yr)\'y<��]?��5+\0[�~[Pۍ�S)mE����6�poq�7���f��ؾ#+|��҂�2E�ף"��[����.�S@��V��q�٨��e%�h�L��hr�6H�pd��0=6�.���:��!�$�'��f2��d�l���N�l�j���,�P-^�8����f�;��"��4��Q�X�b�K`0i���n�9���v�*�{h��"td��t��\;M�dV�N�k�V�h��تU�`o�j�}��x#U���W��݅5L�W�ɛ����J�F�u��"˃z��w��TP줍��l���2�U�ʯf���4G�pӼM����w��;�`̲j��f����I��tv��=�J�m�����ߥ�vb�{��,���R��=����x�dg[]n��p�G�d�q=W�I갨��#0חW�;ls[+�vF��+�ui� �V\kV�GJ�0�۸�u���ޝ�SOU����Dd�<�KԦ�dS�v��N�l溽Rw͉f,k++/�g��>��0Z��S�" %Ў���C����jK������S�$ړ����k�|i�	V/2����Y��)�h���h�u)`�"����o�E,5+J���R�4��}33�H��>&�L~�ݒ4�(����"H�]��V�=���-^�;�p�����j76������o�%�}���g�c�^��i��K�f�<�����1:ةT�E�Wc\�esf�v�짷r<�CY'[�������B+q����8/w�f��F.P�޻v��d3{��xv�040�+��<T�qJ}�7EF���n�TX�꙯��Ru,��g3f^@�{��W86ˏ��h)I�se��p�T�ǹ��ԨT��<�»z��v�M���фYz7/X�����2����
����#�r���v�����,�!L�;�wуÚ��3!��vD�8
GE>�C��������R�C4�@�Mn�7F���N��;�;xl��j��WM[k�{F�T��	x��� �;[��f��Iw:�r�u;Ó�t�Ċ֫2Ò�\&'�o��r�%��3E�=c!d�]7�*�T�;h�P��Z�*�Z%��&��=�W��y&���C�<��!X����y+��γ,��R�.�vv@�/���@����XGzU8�ԏ��#��gSh��uu�b:��C�2��m4��G:}j�]��N/,�eh��s�e��ѩ��sY�Zm��ji:ӊ��o{�ΑW\Gp
��Ur�
=�-%�ُ{�6e��3�u<v/�+�:�9��{��K�ʴٰoM,����ʴ5|O:K�Y{�]��T�;�odc�`.��K8Ṵmգ���*1�3��4�W3.	�wWɥ�aӢ��Y���%B��Nk锳o����p䕡2N����uw*�f����$��Hh�$�*ΔP~�p슛����{%H^����n�A����iV7�����j7���OxmR{)Nyf�P�@�ku|�k�n�Uu�w-Г#1s�9u��Iaۢ�]N��{��h�6�!k�;�ED��,+ނ��T���w��u�)���\��� ݾ���n^U�}};�Ss���	N�uǘ�º"o7�u�J}�u�.���'Q�ɫ �Qr�mԫ�E0�����3�G��ݹ]�o�Z��m=�Q��pm���W�A�8�z��#o,n�،������F�K�3�]G谍���w��ufX�mw��q:�㕏�NBfw=�G�n�J�
O�o^f)��rr�Gٴ��
�p���gM]�~\����������(v�Ө/����N뽬�S�3����7���?� �	!I�L��D�ܜR��/��&���tuom*�zT|�߅��MGt��u	{Ϲ��c]�:G5��Z����d���o�n_FQ��pW'�`�8+�Z;
����lĸ���_0xE1t�Z�W�eٽ�sD�Y\�f���]���F�IYM�{yi����^��p�07��V�QS�Cm�˦;[�N:���jo&��]�޼�[�:���h��]pn��$�p�MR]:��wf�ȁ=����;�Y��ں��|Z�-%[�i�:0��e {+���WS�^�ck��1i��������{�W���oA޾q��;�k��m�+IH+�������PL��.�O��Fp{���a��J����[3��5�n��}��.$��:���oOȣ��3�t2���d�\�=��a���-t��u~^}5�)��3egs��r�ksx��.t��ܵٵ��lժ���FQ��(�Ի��]Уit�k��&�JDis������"k�%�
���;i����.�u�Q���I\h�Û�_ݙ�iF��T����R�;�M�D�i_G����F!t)��R�-Nu�͉lEr�OF�#ɇ��A�n�3��!����M�*$��±����+����T�-T�n���`ۡ���_F�ǵl+,�Z��Cj�ZK"`B�Q��|.���orՌB,i���3�]����Wj�3�nv;m*�Gh�=�	x2x��"��8�&���[mU�8"�u:��j�������c���s�
�U����v��/���8����,Y��S
&��SF�_�hk똶�������m� m�JR��*k<� [Zb�1*��Ʈ���Fn�̪t0
:�ce�.Y�f�yVVl�A���M�b���V6�M�xU��7����^j��x�s�4�,�.�9KiB*��HZ���+�G'+��	��R=C��2yN��̜���G�-�e��\]��X�Pwƞ]" ����.p�T��[�3Q!	��Y0��s�zS�/����+ml�|�q�r*�a��ژ�#Emܼh��(q=��<�����v��� 
��o�S�g�����%ձ��h�י��*?��._B+iR�����wMÒ�����څ�x>��
�W�{%�غ��-7ս�WEn�4a�bK�B�k��B�<Ѻ*"�5H���y5� ������˷F���_J��n����4����v�CB�f��M���.�717t��c�⡜@��+�쵻��@��r4�z</�-��nDfm�J�3�]�^�����2���[) ���֐�Q�䫬�n���yW*�c�(�ck����oyr�z�>�O�u.d��K?{��ɺ��Y"��� M�]|\I�t�7���a!й���Yf�`����7��`.�Wu�N���1V`���׽Z�\�f�Ӓ���|hiT8�	4-\&dy�P3wV�/��{yL5S{:��/�Vm.T��ƶ�n����1�36��0 LN�-�ث�]hZh�Ņ�twu�����{Q�
٢,��[Q�4O]ct%�*,���u�}-�y���/���loe];5,D�4Dwrl��ޮ���֚��Z�o�ɣ�����6�h�er���Y��JW8ޕ0���:yt��ђʠ�B_
�[�����BQY�V()�x��J1.鋅Рx.�uIB9q����ݣ�<M^G%�U�@0�QŨ�ɅĤ2{2�d��S���X6��.�C��!�k$�u�wR���a����Y���,��/^^rXq� �0v��Tv����Q�	o�n��5��7f�^gT�[x똢v�uԛ��yj��+z`׈�&�0V5(Pw� ����4=��c���x%�O:�mAt�їJ&��G�.Zu0���q�Fs�!����ڻiy���5�����HA�X�a�Dzm���+nÝLϵ^#�\��Z/���wWb[V)L��:=`�W�-W˓�v�z1C6��F�tl�Z�jhjj�_m�m���Zj��5,u
�'^t�y:A�b���'|cu��L�oL�Z���uj�r*��с ".��z)�b�E��ӵ��Y糉EB;t/S;�8HF�՛�, o��Z������k�������nƭ�oAS]7a%f�ǵl���"�ت����C�	���w���s�Cg-m�i�*�]g-E���KBަfdEKv\��t��滑��+}/��+j�f��kT���?f�	rԪ�����u�������� ��[Ե!W0	�KMk�����	:��
��-jh[��N����ż�����/l��}TC~\�{��כ�����)�Y���yr��u�*e���Z� �Ɇ�^�Z�]t_0i�*�����G/����&�Vek�����#����+�����U��g?���]�e��-lK�fVV��ICy��hR�x�3%���e-�f���;��D��%Ֆ�&����S�p��y@r��-F�/T�l�����
���
�p�f�eoNb���j�>}lN���
#X�byd+��X��5��&�xR�.ݽ��.o{]�B��+n.�c���@��ktpGQB+k��/m�)�V��U&7�]���t�.<bJD��x�Ԧ�5n������ʒ��6]|̶�Ns�)@ wO86R��ܳ6&-��wrT��=�*���^uL�=����:�O/k���z{�$�f�x?5o����p��zv����=?�����kvQ��.�߱�X&|T�ʁ/��RZ��\�'ԃ�U������6��:��\�˕��"���P��5�AH+�8�-We���'T�M;O6%N�"��\Eश#g"�ŝ/��pb(Po7����rυ�*�;�T`B��GU���ŷz@X)���*�0�в��ѭ���X�v��k��!XT�j�!��3v��f�\Ɗ����>��{�n7�Oj�ż�5��ؚ�� ��4;#�w���Փ�� G�b�����E麍U���Ps���6��'s��S|j�t���\�j�L���ź�o��oB��/����+� 
݄��v-ce�Ƞ�nΛ&�?5�!ʸN0V�od�6������,�b�|��֪y�m�i"6�fu��ה7_]���sh%}h��[���r�a�[�w��9�:ٹC;�x��`/߰�_{5����	��UG�H`u�LazPlQ�S�����A�1�5����T�kp1�H�oe�Q�\�F�:udv�ђ�"wB�*����{��ާ�p�J�-/[Ŋnm֫���U��ή��Sc�B��k��;��ʖt�]�����,��A)���%���yt����li�(��]�cd�6� �����9鿚��eJ�j"����Ybwth��\�2��4�]�(er���,�B��%�������s5�e�A��r�)7�`��/�ɦ��0�p��Y����|-T�oS[v���� ��=�#��lHd�%�7�w>9G!W���T���6ŴL mlSt��w<�g2��!\�m��i�\�T��|;1)��;���!�u6�kq������_z�`��#a
fe�ɮ�;.<F�Gk{�R
��4wMcb'�f���*�t��4]$�ו�8�䝞+S�f) �)bwnWPP@����t��!�1��E*1�r��Ru���7��Y�^%�O�.�[D:=���@�x[F�&7��*c)�TB�34��Xo:�amG�t�*��	pKzI�����X�R�C�Mbv����GXָmCt7�
淂��]A;v���Rl�!�/B u�3�nx��v�fq��1u�P:�(j+����-���=x�r���Еq�OJ��w�6R�K{W��yv���7/���짖���U1�@��_̀���r� ���#��0�ݧ�%��n�K���{��@]q���� ͆j`K9�9�/�����u���rY�,�+Ae��JQTء	���]��R67� 6��Խ�O�l|�5�!��3Mg;e�%�v*-�*U��̫�èlj��s�Y�{�Z�X`����B���-�~�iiz��v��l钎0h�g颍'�`h+��M�=��
�+4Ӓѻ�G4��������q0�̗Ԋ�7[��vh��L�6j	4bx1�ܳճ��B}8�ch^�j���f
�Ŝ�.�Xy&mn "�M����D�O���E�y���P<�n�o�r�<(X˨$�+��)�r���o�o����I�hcC�-���B�gX�Ж󲯮�:�9G]�-=��W�m&��jK�	"ٗs�9����̝09(�.����hW'g�8�Y1"���v�q�97��2i{x���[�YUш$��ʽa�t���:F���g�<�(#��w�u����;��-�+]�c����²}uhm���N:��9w}�V0)-JTu'VܘF��$:�9%v���i�Rb�S[:����#5�ov�S�f\�����W�=O��V5�E�z���4��C����%����љh@wh�w�R9V���8���J.Q�iChc]#{ldS�\����� (d���g��������)/j�UF��+6̛�0�������N�j�ΨwG@�m�9��Ki��#�kLZYXp]����r����)�%f�����ג0���5���u
hq]4vN3e�5�2[Ϯ]��q��9��|7y#Ó�ݨf�O%�UR;�=�R�֊�9jo��8��Vk�n:��;^7�:MS�;3 ��2��9K����X�LT�Ĝ�Ewyr�et���@�V�e�z��;���{*�J���'�ic|�Ъ������<�ԍ��T�{�����\��:��*z��._�fBy2���5���R���Y�e�a���L�W�Q+����<`�( ��X%ژ�������WHF��HTWVWV�Q��O9񦯠�Y]HA��ϲ���Ѳ��lT�М�DE�`̣֑������� ��}wǠ�ξ�b���̞�����P섄6��Q(���0��cYS4�)_(��,Hձ�Jvp�oE�)Vj����M��YǄ�'G:��l�b���M�,۽���Ry���W|��V8"SҐ�Cc�^�ЋJ*��[|,�u�3!g]��9��^cۺ���]z�7".�+�����mXb���us�ZڈT�/7�Z�i��t�V�q�٤편Z�����[UP�߂?��-n?�&�7���b��l�vvg����6�+]�]���-��u�r�2�r��8Wi�����f�g��R�x�� �Wb�E>]ݿ) s'.�"�$՝x�*��]��������i��bWΒ�tc��^�\��z\���Q"8�k�7�fħ�F�_��.
XUk��6|���#�U㓹c�W�`������t(IS��h�rN�f�t{�U�n����V�q�9\j���-�v�B�d�|�*\Wq��ru���E�E��}��"��0A��-;xɴ��r�<���e���Ry˘�W�d�6�F��֌mao�������lʈ��c�����妓���R>x��"�O�@V���c��v�����C*VH��r�Ԕrre�M	��ӧ�ܘ��+�%�� B��ަ��k�l��a�\�m�6�"�1���z_#W֩�ʴW��f����D�(�X{J��T܎-�ԯ��r��V*�8i_K�s^���bɨ]�/�u�b�@R�#y.>�0�̩dꅹt�� p��� ������D��wM�cv���Zxy����#�n�����E�:�PKc��m�6�E�����oj�O&��݅��ܡ+���J��O�u8�ïT�YBX���K�:U��;$�lZ�� sCzf[�)Ϧ��e)�3v�l�Z��v��U��о�M�Fb���w*��SR�ë��F��2�4m�xj��UNkT�&^�U�A,�T���V8�;��-<�.n�����a�F�����e5P ����%j�1��Wn֎Ł�����˴P�pͫ9�v8زPݬ�n� ���%4[Rٺ��k�+^�A����v��
X*
����$5�W���гu|�f�>������΂;n���i�X�z�\�轺�J��E���b,�V��0��@�ȴ�&�(u�s�Ѐ�l� �����+�3��;т+g75o5w�e��O���S \�����oP�-�/���\7v�|ֶ��q]2�ɗ�&N���b��V�ȩ���t��r��I�kw���7��o���r�V6�����KVc}|���[�~s�s�ܻ���qb��+�:�>�Z��]�O���K�J�=�4Ś��;��/��Gr|j�b�m�'�5wX�x�ś�Y$�@9�w;AE�d�)�x5Q�(*�_ ��ݣo{M��	o������*\P�����yfw:�<"����䚭���� �q��,l��Y��8�l�]Ä}��1c^.4@�����9����С[N��Uc�Ͳ3����DV;Z�L^.ytD�8_K�����E���N��WY{)�].Q�Q��(����y�L�)�Ioj�u��b�D��׏Q7�f�<=w��ֶn=�9s$�oPP�:�7wP�Y\ݠI��H�z��k�)�k%DsK[�k�s-��Bo������avs��_3�
K���e[���[���%pڌ��)��f�w]u�V.R�����0B�˚N���I�Oe�N	S�du���־�[��'e��+j���|Z������f�[��tQ���|���n�Ytkϼ?���$eT����\�q�ܡ�Q��ȩ��j�����*=J`u�;{I�Hh33��]���6lz��"�N�LQ+�\�Ն��9(3Y�ce�P���W���mM���h�Z�-=2��HB����f�_�8�:���v�-}6)Ny�5�q�+@Ef*���\��E�"����D������b�V�Զ!s(T��y��P['[�6;o�к�n�wE�.Y<3�u����n�&tgZ�9I����K~}ՠ*��$�]�cz]\���+-+����O-�����;�lֽ`e�T���"�Q�yl�<C<Q�X��T���zD�lJ�Z�y��k��f{�����4o�i�x[�@�l���7Z�8�7�/��]�w=�aRN�ኈ�nb=+r��rx%�>{�9p�X�����B�HUe����(��J�C�F�nv���݃{c=צ5s����뇍>|"�zŰ_�4��N����U��h����,��"\,Sx�TA���8w0������� ��Ш96m�IM�YIo��8���8���銭Z΢0�xu�]����x���!ypǳ�DK��l�� ]�r�W(� �$��]t<*d��u�y|sQ��Q����V� �� ���OxW^%ͷ§'����ݹ*hU�ԛH1���x���"�j��R�N�k����d�Q`�ՀG�ԙ�\�w�Ѽt>6��+kB��;���WTɳ<"��F)� ޝS�ʴ��KX_����#��%ai�m��}�B���W�:��M7BI�q�5������q�b<+2-s��'Ǻ����Db�ъ6£�qQU�J�+Ke�ԫ�Q�V0U�hQ��ETAPLJ#X�+X`�����ml`�R�%b�E�TG���A��U\s(�DAU������G�2�A*V*�T��*�U�QZ�c(����R�m+��1�R�V��,�3%`�*B��EP��b*�b
* �E-�[eA�,D,����B���"�+UjX�"���V�EfZ��Ls()�D�+R,EEJ̵�W-���)A��R����EQAR�%�UKh�H-l��il`����TF�Em�YTE��"# Pm*2�UUF1+PQ`�V+Z��*�!U
"�E%j#�"b1DR"�0Em���"(1EERZUUY�
�c"1�b(*1���UjUH�Tb�J�A7����oq���>A�����@a�Kk��|���J%n�u���X�O�l}��F�VcZ� *¹��s��{[�g|�=�iIs��ޫz�5�;n�[��ʝ��;'���)����p�"���#.fn�[�v �=�r��&��s�J�%�}���P��[�����ζ�e�u�a��t�Eb���a�@z����Ȏ���si�[8t� ��!�yAW*�"�_,G��+â5���C�(���fx��л��:�_�Q���<j�ҹK5��BO��:$>\��)j�5��q����;W{]�-�6=�2��}O��.��.q
�G�Bjf�1��y�D��K%o��o�'hCx�Q��w�'����,g	Gw T�uV�2n���op���Vf�V�5AQ����4#)X��E�R�T(�Cv�s�9�ͻ��?��;��ɓr�F	���|e�f����ܢI8#Y���J^�,�2�PJ)W\#��^���䭳":>�{�x>���*b�ηK���)�v~_�<]��p�2Ɩ�g�f�	�i�{ue�9��P�}-`�M��f�b��
tt�*����D�ԭ�kgN\�#�Q�h��߳Eq��:�_t>�k�:Kt2��QQ��J<�;��8�U�h�e�C
��Iq\��M״*�3�v�˛�&.⸻��+j&8��� [��V�H�j��d����96�Hݷ��p�Y;+.��v�TY!�(�D�#��1QA'D�`.w~���Mۊ⃵4y���.:�Q9y�,h�/|V�*#bY��W�vz�M}�*�T'���� �-5�l�~��_���r�$n�O��^�����.�W�=\Yƌv+(Aa}x��WP#<k�T V�Ew{gz5�R����ly�	����_�Y��@`ffzk���sՊ�ᳲ7�ꝗ%\��α��W@ר�9|�� u��\����r+G0ڈ!��н�����<�W�\�f���ٚ-p�6 �*�ܯ\��0!�_-ٍ�����`VH�QO|l�֗.�-j;;R�ˡ.�
:lT�豊I�c��!�{B�r�tK��n�=GG�nl.�3kix"XC�Ы��d�4S=N�`���.$#Bn���
=�i����G&mhZ ���,ui�x����x��U�Z��[r�k��Y\k�cU���A|�?
=��93��A�4n߻�.�
�v82%E(�M�U�UR����mn�KPwryIz�m����TAdݭ��̚��!����1����;|rb��ˊ��Ch�����G�gX D�p��������2���	����զJ�b:���UϤ[��o��<��*��
<8�g]�R�
�tc�T���ٙ����ú��eJ*�Ԓ�15d<�QBܒŅ��a��$�%(����Mx�P5cR,\�J�xU�j�g+��c��z�uqW2�9��Sك���
������k�>Gd�`��f�،�����	F.@����Qf:�DF';��U���F���5:�F���/v�����Q�Ч�۔���wJ��*��[i���pDH�s�,�-�V���Fr��(�TK�יN,�Lz�5�E��Q�*�@�])	S@�<e��x��~W���z�3�}� milTa��w�?��]8�K�<X!��1��Xʙe,A�*�����Bx�E}����S�ԇ��6��_�V$>� ��,m�S�}F�J���\�{�H���q]d��8_�(,�JT�� �&c��m���3���mE��k�S�@����T͜(|p�0z�[���EcW��G��"#0�w�ou��=�q�$?�Ț�٪��ȓ>�$��d����P-��!w�>�3S5r~{��|u�ܶ�f�x��8\<We�4�p�����u[���U+�)-V�sv~�(,��;��G�3]�j����f<J�d�����w7V ɜ��JkA�̨$0*.���/h�z�ᔮu޲��3�9g�3�
,���H#��PF��y��32��o�/?��$D�$+��qca�r�]�j P�4��M�<nv訢�t��O�sL����*�[���})��j�N��}*F���}⎗���yn�L���w��ײ��������RLhRKG�Ǉ�3k���)U�'�m�Il���6{v_�,�{[�sy�g��"=��ûS�a9sJ�G$*��m��)-�����7S�_�ّ�WG�%�q�,�r�c��H���;���dsukFEf��ޥ�zM�
�����j�%7b���\�X'Z�R���{o$��k��r�b5��o��F���J a@�D�j�	�e�@W�ϓ�1�'.iD�Z���\�q��T۞�����}�!��LQs�jMj�f�o0HDk���g0{,W/]���]�Lë4�ꆼ W�V[O��TP������g����|���M u�c�{LoZ՝<�΍4�Y#��eN
qAԠk�,�dwN���,�񉀫��y�A�&��u�w��x��q|�3o(�А��Xv��m^%ӯo[�R��/i ���#�*�k���CT�9�\� ֗�n�g�-	��ݭ�9v>1F�@�s��t����퍯bظ���gt��Z�ۚ�yj�p\!#�#0$
��U^�BcQˏ�0�_R;AUA:p9)�yT�E����p`@�MRj:�=��^?]�^M�&�U�a��7�
�Ȭ����z	�$E*�ݕ�}������3�����5�B��7�nz�W�O�\�l2~�2��y�R�z������H� �	�_��o���u��Nn�տ�9�T6�ӞKa �X>J[�]my��q���I
�q��va����Ҩkj�h�]�b����o���g�Ƿ��zE�q�j{G��$�����#�$�(�{��:m��6ƽ�豊vO|�X�W�D%ZZ:��7=���m�ob��Q����VƖj�ҹK5��A�_H���*�؅*y@��"�u��c>���{.>�٘��h�{�?eO����S�9��6���VZ"�(�u�S'P�<�^E�r֟^��Z����Z���Ig�TB(��"E�V��#�)�]l�w\7���i�Lh��)�a�'�'� ���
%Lv�&�r�av�Q]�B�T9�t:*T3e`:%��wJ7B��(T���{E�_x��)^�V�̼����tɺ�[J�<����kC�|W�F�����|�՜k����VVe�RK˻Z�����[ú\%u(9�S�e�W�{�Ml!W��(�*)ru(���wM��IqY�� U���Y|'� 8?��������a]"��@�hž
�a�(z��RU�w��zc�fUz/qC�{���D�K�F�狷G��x�Rq�=,�V���(uͯM�Z�zup�U�.��1U��N��DC
��rٛ���U�� �GTY�w4K8]�jv��>n-L�4{��UKەe����fS��zY�|��j�@`����2���]��Y�u���L���1QA'D�~S>��{1��*p,�MF�]����z3�R��DlK5+�ʼ���Y)�/���'Љշ���ܰM��ڣ�K���g~��t}A�2��Y���xo�G�9�ʦ�%6�uc4Ҭ~�4�i�zfv
�b���v^�_\G}x?���e�|<0*33�]SX�G:8�:<ϼ�V^�p��4��pXB�(~��eS�hD�,s�0Qf�sι{�,׃���L#�(��#%׎��r�{M�X6O9���k-��]p̸�����O@F�Y�T)u��˖-�u�V�)!���y�U]=��3l���o�����bɒc�4�D4���hh��{5Q
�Qg]��r�N��s�3��*����vin�����9$��� :�iP\k�.�8�����1�}ɸ.�^c���|���p:�u�Ω�k]7��<��}9�k1b�V�.�Y��ڈ��9η�������#�k"=R�$i�5�Jz�I��H�Ƌ6UJ�I���q#�Vg�r���Y�Yr��A��U��r��^�y����s�z[�=L;U��(��b*�ToOT�u-)�%s�\��=�Z��u�OR�����l��c;�K�g�D�G�!�$�z��mEU=���n�gc���q��~��"��V�h6Cȯ<�Ȥ�Xx[BJ��c��@K�'f�ˤ�;:gz���.�
���,�óe����{�6�c"��V*�[��t@G.���Q���2��d<�� ���lV���+���t)eD6 �vw��&�|쵝:�w��GEVk=�(�#�3o��=�6*�u�*���j�^�'û�1AU�������E��y40����^t+�L�]�^�����Jb]�r�d@�"S�`o_��p ��[DkQ0�|88]?nMT��K�b��@��+�T$N1��:�,r�ʨ6:{���"��ˋS�8�y'f���s���Ż��Ӭ]�H�IS헜�+�!�!��
�n�hu^L}9�F��q6{qۅ�
N:��hwy����������U�A=�/��u8�ͷX���ǈ�)AjM;���f��&����u
��7c�02�$Q[N�.�ě.p�f�J[4,�rWg�b��V�;��=����M� l���'�:�n8�Xi׶M��j�τM�$��G-;�7�����q��T����[��W���#0:���̋���<4b��#�Rk}�}Re��_��f|���T�	x��*C�@�j��x��^�{_#J�uֆI�K�-���G.��c�tJ�y�lퟡ��Q�vB�V�\�!̌
F����l����x�ugR]��9D�Q"�z��]Զ��}iű��})��r���Px4]��T��������JU*	��α��*ک0�t�h��M�feK��#t���-5�pU�î���͕�S7�!�ؿv�tE��
�=�(O`�w�.�e�{F[��檞�!.��&gn�S�p,���Q^�+���cTi�HN����R���U�β�d���l�I�ËhS3i��i�P�Tg��u.���
�9�m�l�[&�I���{��Y���=�|�/%�M�H�62�;�u�4��չ*�el�)��&���$�] ���V�}�%.[�m��Vx�<e��
X{r����F��+!t�<C6�n��8N�U���x�eY���Y,�ׁ�w��g���Ƕ`�_�:��ywz��Mu�X��&ɹ���,)9S�P�<w5��B�O
}�j�w����+-kx��o�N�Q�|>�C�ү@�r�ҏ�P㉂	��.�&�+/b��ȣ�2�اN�,��t�E�Oˮ��yl��DW�،=VH�'ؐ7]��kE��\*�հ���o�v��7���z��p"Ñd��o.M���EA�G�>�9�tlW-w���_P�d�}����)��4+dt�p�G�T��ݷ�!�� J�W�
�y�F�D��]�r�Ώ�TZ�9�S�x#0{9�)V�ތH��g,&6��"�4��n�o+qYiwɭ5��r�&�ٌ�+9X)���Z�>�"��]y�q"\^�������]��66��ۀ������T@���଻=W��uEC�K!����.6߹�띯��2�7���gK.Ǿ�`��$������!P��ٲ8�k�#�S�
���L�Y�s�� ���2%����o�V)lֆe���G��Yպ���wXI]h!>g�T�xH�M��bެ�bT���Np��{�W��<`����B�!���u�rۜ��e�P~j���,V��oX]��[��^�w�0��j���9ST�'�����υ8��-�����S�o��d���;�'>xz�.B��|��h���ٓ�K3еK4��f�W�2�)���`pu/�J��ux�������z�'�w���[�$�`�%���/�{ܯ�Cb�f��v��o�|��g�PȻ��[ї&-z�ٝ�j5�t�f����E�*�)� �-�����7��8J;�W�Hn�U��UĳǟO�E��S�	<���E����eز��*�Qx�,�K#*{0�	�<�ptf�ϫ� 8?�����M`:�|��RJ��`4=��,O�Y��#bdg�����@[�iD�0�`@N bK�ϱ}�i�zl^�ޞ���i��HUjؠt�CD2�.�"�"0�tup�WCt7nJۥ`ء���!�7���F(����6�
���� �MϷ����0�6a�>N/�Sd���)�\�B��R��'��V�QWk�~UPY&�pℑ�w9�`���r�MD#C�,�D�QF�;���������2��̓E�+�s�:��}H���\j#�Д~�hU`1ԩ���+AQ�[X�ގ���de��Q�D��\e���8{$�R��L*QO�#�������}��d�(��0K�h�V��et�a
f�m[��wmS*Q�+2�v�-�tQh�5E �\��N����a�Nj�M����A�,:���SVGS��j��YsW��L=�5`���{�
{��3�,�`w>���}R>�#+��蛣�K�^'�Gf�ZЧ�qۦ��;Y���A�,��4�.�%r�+�<����E�=�]>�9X�MZ�����z�r�G��0$�������I���.�2�C������U��v���{;��%�n�=σD��#T��ۓ!E]-�-�u|���:�<#y����V�� �K�s	��Ep�q洫T�{9n�t���Js��[\������ZB�f�]��Ol��A�-�2g<6���k*-��u"�Иc�Z�J�J;Wկ�s�ll�W[�둷)�*{��i�묬�Vf�wjn�opw�mi}��uP�N�ԮNX6殰;�ʰ#t���J|&j�5����u;��=�W��w��sC��Z�m��c8姶��gղ�NT��/-��wE��e��&��X���G�-74%��l��eڻ��Y:ũ;{�%�*Xs���v��Ǜ���r�<���q�jZ�!Vcu��~�V�s�:_��du��`X�17+Opk�=`*�]�'��OM��9�,��§/���w��K73�^僛3�m�$_�M�3`��5�[���Ƙ�r^ ar4$�O�W�
g�ۑ
'
nƜ+@��8�]Sq�����g�J�&�!��8�N���%�LJ�<	kk��L��qH����L��p^`$ʳ]�wf���Z�Ok��e:��r��ĝ�W�m�X�AM�ŐD��6��X��]Z�%�.�A���nkD�Y��m�7TcC���Anܳ8��[��M��a�}K��8��'�=q��C�촙NF���b����EŊ#�`7=���	�A�݇jl;Mt$��U�0�M-��/�$�<Q�L���U7���9Mz� ��ڳ�&����(�d�!<ܵ�V�p�A�^�iOV	��+8?�;�����0}�Վj����<4�9�ؚ|�+[l��_]��8:��)�k�vT�7�2���x>aѲ�؜�Ԛ+�Kk],���w�<fx��Ng�8�ȷ�&8ϔx�9�Jn(�y��MV���*%���А;�8s,V�TkU(���j
�b�F,�Ҩ��T��QUbʊV1b
�Pe�UF1��թdV)�F[b���dQb�UTPQ��,m�X�R,UPD�"-�Q`�B�E�AA��hPQE����*�R(�����E
�FDb֢�jT"�c-�
�+)QV(�U�*,PQ�eB�X��)mUUU�mTVE(�c�ERȶ��`**Q��*
�"�`�Ȗ�P`���V`�EQU��(�d�Q�2�U�PU"�H�U-���إ�Q"�l�UZʈ����QUD`�ZQF*[Q�*�(E"�"��Ym�U�ţb��%E��J�Yl_A �>#Tm�%|N��e�_��-n-]�2�ќ��HZ�T�8�¸�S��gi�մqΙ�e��Ú����HR�N)�T���7': �MeA�YW ���>wg���xjz*����g��H�c(p��x˹2ʭ>���hX"*^D�{fQ��a���Y�� No� Bf/�����1F����c}N�I]Ǻ@͊��@�nhN�^Y�g;��)��nD87��Ԟ>�֗���w'wDO�Nu��������}�o�x��
��kf<����Ɓ���[#3��nyʛ(��sә���Z� D�7Wު��/��?:��N+�ҵ�V*1ou��;ˊ�����á�*#Ehc�˝M�Vٮ��WQK<��袈�s����ėnzv�����ޥ�G����;ӂ��Ӓ'�s��i�(l�!������&m�ac��(��y�B��3���,K�Ú�>:,r���:���r����i����s_�6��\���ݓt҃c��54��ޞV�h6CȠ�c"�������@�:�;�z��������&��u@��8ߏo&i������A�t�R�sN�w��hQ���M�bJ���>� �ԌB��˵��6���QC/)�=�:Ym�o��W��+�����u���O�tʜ8��ܦ74@��ь��Rs�	���в��٫t��qӪ.�E�SNtJ��[�;��)�����W��S�oo$�u�2�W|ƌ�V tQ��%�yzwa\Ζ���Tʈz �s��J"�ǯ;DmR�,&�{��)��E*v�_�R��r�Э��|k"���N�XKY�̈́w[��j$,#���&g��[<vP��a�5؁�8-���YJ��WR� ��A�2n�nz�BS��
C����6 �? lU�Zч}�,pz���O+�e�ˈ��Y��v9�o#�`�q�+���QG���N��1��Ċ+���i�X�k�.�O;:yr7KT�J�av"hl�.��H��c~�W^4�	��K𹊐`�f�`�b{6n��C}�h������k���n��A�W���b�,�xΫ�_ep��t�8���Lñy�(�SA���!異=�-@R��T�8ݚ�nŔI��L�<��P-��:\r�Β��C���|��<��4|�rDA�Ӳ�K豰�Qf�;t�%�f�Y��)��&�8�~�y�V�fmsXz��Ub��|>#Y��Fq�������8�}ѩ��4E>��^ۣٔ��3�-:^,�%��%������topn��x5tCJ�lZz��Rܦ���>@�\�X��Ω1�,i����M���7J� �5�
��NF����)�=U�Jd� ���X�-\R�=��5r���vr�?'�d�F��jDʐ�p��cq>�"�-��
�U�4V
�*gX����yu������&3�H'�l�Z�3y��A9dTr�Z/}�*)9s	�c36i�\�.�������[�}�]T5�vZ�i�8/h�Ӄ�_tpT��^f!�ёM��w�?wa'0��9u����z���6�Ć�p���Mح�0���Xcv�M�_�����;pu�T#��:s����=�ѴFt>���2w�U�]5��\��)����p
x�>��ez�t�b�h;$�-O04x|�#��Z#x�W����V�.�"��"��!K�8ɗ-��E�d7=�Ϳ2!�E���_o�R�o������:�ꄄJȧ�Ǻ,p�\���Q��^=��������>�l����xD1�25���;��p;��H�S{oՊ���K9 *�"F�.���Np*�8��E�\fQP_(�c8���_�D�u(�Z���Y����k�ʭ^�"��QKz�*���Ôrmm�/w4�ܛ����c�fx��pj�zG�)q]ncW*M#�+�s([V�e��bU��W��ї6�)���X��t]�g];��u�-b��k�LwA7ہ�lJ��Y�v��i�W��Z�9|��kP�H���ݰr�$V����Ŋ��h�]d��������%��}�+�ʩf��>
˫=��e����xz�'HO�[�]��g�o�w��~� 3#]�μ�x+�����
�
��ݾlh9y;��V��C�C uN3��3�5͑��m�w.��%sx��f�t�!�U<d��fr��z�ф�͑��tB,ĩ�]6��>�dZe��xC�b�Y�J^>�=NU��]U���VL�^�,�B�,��3@��a:�Zpm�Ie�5�/��׋M����N4���%��w��wR��6mK��K���-���m���r���M�#�L�K��JV.|�� t����m��a
{��I�Y�C۴����'go�㍋�U����9�H��䠵����[@ةE�r�@b��2�>��9�����i:`�Ab��W`@pb���Қ����|������'���\�S�q��4�bBR�!c��W�����@{�8�8�,MCլ�s��-)Aӻ�!���w� Kn�b�j7�u`n�ĭar:���o_sȄ����z��AW�qپ���h���G���
��,�7�Yͳo��\ugbk�6�X:�p�� �(hbt|//��m<RAC�ό��]��l�h�*3���Ő�z'y_� <2*�6�v��Ǿix'�9�Ǿ��s^�Ƌ���:���k���' 00���..�N�ͷ�g�n�C�q�U��d�Er��%���T�(����1����ۺ'��!P�s�S�D�t赵���[�j��dh �ο��%!O�}�Y�u�������|�5��ǒf�[����b��ڞ�X�1�1�D\ƛ�Q�"���JuK��m`$so7_C�ږNou�Td��c"�s���f��O����/�ep3�Ŝ�nV�b�F��{@����E��8�J��b����`#����n���:�y'�}<���i�% �S龱6�N���e���V�LUW����_k�AѯO'z����KU����Q�8u��@�9���3rnG����T����.�z��4����D��]ʀ�O{�֐l�ɕ1J\���]�ܮ=P���{^WfQ󮔥ZB�6�x���kB��r�������	�T�f��֋jp�ѭ��"�t�B<VJ�eD�@YP�	���hpþ��~�\�J�֫��`��X,!&!���p���|{6��yV+:���u�R���{TSYT��)���	Qb�\�Ӣ��92�����$�eJ�vd��s�n=�Io0U��{��cN6�Aݮ�K�e����zV�M�o�,�ʪ���{q�y���TU���yCO�+��|�z-w����N�.u\���	_yo]	�f�L����\���P�N3;�;��/(3`GeJ��I��%GH.�;�IT������ר��%�⍿d�MN[�"��{��j��F��}]��^���Ч��u��L>���Ǔ�, 3�`J&��:�tcv�l��N����8J�"-��]0��j3'b*��^jJn���1ȉ�N�*� 	�d��x}��Y���8���niW
);�ܽ���]T��u<�4�4�X��(Ћڒ*qe�$��0������E�4������Z�� �#���'<�����xt��4E��d"u�Yp��k{U��}\��#��pR���rv u�L(�!�	�TÍ�fh�a>��5:�m�E�
V>���C���� ����=��+:��1n(�`�hs��~�6��]�Ulu4�uwNڼ�����J?Y���ޝ�0Y8��U�*��R<����q\4����h Uk�@��k�c���|8.wY%��c0$�1qJ�T���15�4�kD��%	��wh�xe3�7���-:�H��El]�45w�q9��f����su�=��r� ��;�q��Z���\���9X��++���|d��}�}��,��^��qY��3HS�����;ax��|�;���L|�c�`�e����v�w���8y�<�;x9�� )P��ID����Θ7�	��0�=���ab�&��Jq�B�d��s�1��� 8o�_�ªZ�����bZ��Sӓ��wR]�h��%�w.szJ���@�v��_cC�誱l:�}zI�a���z�Jپ����/�tՀ���7��g*R���K�lj{RG[U&�U��i,E�X��u��研_�E�O�3��K�v6l�J��!��N#���z6eB"���j���wz�zͻF��=��$�����]�[b�(d��s�-"I��
D�i���?wL��kX���oj��(���^�L�At J�j�,UaP݁��]3X��c��W]χ���/�����1�(�ҀP�O.��e�LEY��+�2+/a%j�����Vjϕ���H��,<���h����z���v��A���e-�'�%��d��ol�ˑN7�z�Z�=���q�3f�jJ��x�[3�U�/�̈J�A�G��z1&���2��#-��C ķ�"8���|���tA�­j����ٳ����u�[[�c�4�i�t�1�[����ج=�y��H�{l�x���,�r�L�j�iӻ�5x���bt2r�]|�꺈I�h�2��p6��FV쭨�����<:Յ�\�����_\�D���ʮ����E�ȲL��\�WU�C�Ͻ��>�f���t/Mc��|�K.ywh�4�]1y�uz��s�]��Ls�ug5{��O*�������a�*�f�;�.^Ϯ,�u��3DO@.�%9�SG.p�͐|�l�{���Ǩ��^!3VQ*
2�K(u�
��`�V�y��NH�=[~��f`U��E����if�7&63�xM;/)/�*>̕�8k����=<����,����%*�ڦT�| B�D�� ߾1��������}�%o�7�\~/u�D���B�zGC$�q����Ȋ�#�[U�F�x�^P��/��+��ܧq��w���Z����cn<KẬ�mY�t�B�k۞��)ل]j��T�Y;�k�{�KQב�z�CET��V��GD�������q�KDe/r��YĎI�ȶ��9��t���M��$���㵉}�������6̀�>7��nb�G�+Rk�G���u�uH�}=�@��'�ᗜ���hVZ�D���Z���aU]Yf��ʫI,��8~ �OM'I��V�ڣ��"K8Q�n*B�
�)X��Ċ$ԹJ'*QDA-�qݫ���kWMʢ�7<�#�U�g=�H��䢡�%X��`�U �*�oX������{�
~�M�Q�Q4n���s���G�����ٌ����V|�h�����Ʀb�����[�D�h]��!f���w�y��kӚh+��&���zk�e�����8�)�l�X&���z=�Tћ��`<S��;�"Ɓ��:���\�S9`u�k�}oN8��Y�(���$�GT0!���$A�B��(j��z!���$�dQ8�10�΁��NC�����5~����_e�A��g	���S�����Y��=(��r
9�$���~MO2�<dۺ��[)�g�agl�i�U����^|� ��ǒ�~.^w#Ң��ή߀�⍚���_��?9��_#^�g�jL����z��v��A��8'�Nb��wk8xL80��WPT�����nЈ�O���p34V[VAYMoyu�!�6�g������Sٚ�맽���xj���;u�f:���dڸ���f�v��o,(}j���h�넫��|x����hC��U+�t�����۾�:�[I�Z��:�Ή��c�U�O�iw���߬�S��}�xxW�1��Z�FY���p�2c��d�������^�8Axd�\����lt����I�]�W`�,�M�`�C���컦��M3�f�Y�:�S�����3�<��-�f�$]�}���r��z�1�3���vK��\�e����S��Z��� �#1o�:�y��2�*���j��iFJ<UJ�g�'���gR�<Y���]�K:`�BW�Ss��h�s�:.��<]zsD��s��i����):��@(=�ۇw���
Ĕ���T���Q�2���vE��؎ʕ�ԙ.lJ$�Y���a2�L��S�޷e �آhT�9��e�9np���8b�Cؾm\�g��uܩү�𾦭ǯ6��ab��|�5���Q5�i��:8ᕇ��elks�(�=�81��N��\8�z�\-���^�����J�:Ռ�:b ѵd�x���Y���	�b�ͼ�#�]��A]9�����1�,�R#�:���0Y���"��YbI)��HX=�9ޮ�х��ǚ����i�飻{Yb������f�Ba��3#'�M�ꤩ��m�1�B9"��oLmj}�v@�/7��ZKh]��f1bJ���b�����l�g���ҭ]F� �iW���w(��f�\n��m�e��c;���5�v�'aDzi$����k6�EY����z������.� �{��p�)s���5� }*�!^kި����&�3f��)�OT���s�ywQٓfjfP���`�v^G:�D+�.�0H��'tA�E�T�Z��u�1��гvO�u�ѝ*v.��{dv��d�V�!�qT�z��x��y�S��t7�Q��{c��yO�lR�*b�Y*e&���jN�[`ʝ�F����tg6�t�;&Q���7�;�����j���	���I=��[\�	���q�,��ˤ1��;h*7K�l�6X�@⢣Y��u{9�ԮU�5��Ab�΃ܒ��V�Z��]��P��&��q�w�)ʾ}ܴ��v���ۧ�erˆ�j|oz���΃utq|]h�kz���n��O�<�{(�[��r斓����K	m���r�=Y{}!��q�N1�+��sI֮LKp�3�9��i�����U[a]�9��H���a�8��t!�u�̛gӊ�V�G�L�ܦ�\a�mEF�iM;W�_`�~:Q�W���/l:Lu�xyF���Y��L��)t�媝X�����\�2��sT�bL�d!D��3��-�$<ٰ˴Ch|����UI��
�L�ܐAg�[��;B�B����f���u{'1��Y=@�2�S$�ч������+�uD
ƽP���~�-��[QdUND�[
\"ݗ]B�����Tw��'�2�n�7cF!CT@*� ��"��T���껕�0��E˷~:�ot��z�|�5��w=�X��}�`�����_gFGw+�sT�'����Z���R!]�\��G��A���T��-(^�����h�Ĉ��VA�̩�Q�[y�c��[�V������ �(�g��Q�f���հ;��oBD�A��c=2�Q����7bڄ���:�K�x=ChQ���6�f�g ��c��1�����P�n��H1�/���a��˓������qA��:���3��F����B�{�'EY�*oVeՎ|�C�l>KcS��52����XJ�q38��֩�����%c/#��i��5�w��t
��R[�;;F�46�Qpۧ�d�׵r
쨦�,�H�]����o�`��c3HY�kVa�z_5m,1t6�؈��pRbY����#(���{�ё�좎j=қ���n��5�7W��s{&��X{}4f���>7�x�о5�DEgR���V�Y�@
1F��%��lf�۪b�vU0̺V^��jݝF��iq4RGNwTô��p�]�.�ŪMT�qѪQ�rݑ�*�i��[�2<��Lފ�CԲj��$�cV:�&�+h���K*�4�c�j+�J���ڔ�o΄��	�Ny�r����p��2m����V�� �P"*�Z�h�@TQPZŪ"�D@F,U-��Um�D������Q��,����0X(���1(�UPUd�E(�,F,mV
(AVEPQb""����"�bʕU�AATe`��b���"$PX�*5�X�Q�%�TQ�X�����TU�QX�AUb�AV
��(�� ����,+PU �0E5�l�D�V��6�V��(��*�,A��U �PPQ`�`�*���H�J�
"E�YiPr�V�DE��
*��Ɩ�UT�X���#�PP�X��FDV��R,�FV�TU�+��,AS���e�0� �s:�Z�ڮ�4�8����v��v(�JU�*�.�g^<��{���؞+{����\ ���0Y3�_ =�W��(o]�뾪��Äa�,�0��#�o�O��`jG��ýj�01L\4���[�Tr�t/�aWD�s�S�5���b����v��n:����9�o�/���xcZ5n��۾K{xJ|�K�*�D*��=a�i�T4�d!Ω��4��#�Y�J%���}z�v�}Y�QQ����ͷ���PY8��TqGS�jG�:�n8��i
�n��_�?)ۧ�'ݫ
T���E�b�!kvSP;2�xj������>��ˆf{=�N'sk[»�],��&�H�"3^@R��7�[u<اJ���R�AQ�Ա9��K+Ŀ�]Po��(�[�����U?j������?g��Å�U��+<V!��/�QT�js��˹	��}p�ޢhR��
�{4�]����}��*�[�g9̣8m���&���:�������K�F�jp�;�sS�O��(��x�]{+;�Э���0��OW]M��.�&!0aC<��f�W�+g0l�wa3�C�:�wv&�2ZH�'5��=Kp��y�ɪX0Y��7B����n�Hr��Jdk}n;��e<�)��4�o{�6�ѕ%���0����C:k0�5�w����P���r��r�����z��b<�jV�P��w�8xu���ir�	�#3�������Z5ؓP��������!se,�`������TEw	u�ib�A.!�?^V�Op��)�����6}l�D;�ˑkH����/P�Gu�!�@�/_
��n6�׮RFqL&m�Ν}�(���òk#�����v�PtT��l��w:
7��\�~��`f����xGX���
a���}�/I<�:>w���B��+ք�KQ|��*�;���R�4���+��PdR������E^ I<п�ͨH#�џj�K|�ݓgw//o�L���xxL=���I!H�u�q��N3Ν�l�w�W/<N�o�p�c�s0_]z�
��v+^��^�3�"�S��ݱ��~gRr�����f����0Olx0�3ە���*��7��N��J���`�=u���Y��0�֧vxW\1�-+ vT��;�پ8P��F�L����5�Z2�ʁ�A_xPK��Z��Y�>{~){:���pؕ[:L�D�<���͜�&:2�.�������򴄼=��-(���Z@��r�i_���Kt ����q;r���9��z�:�w�#�:v f�r��Kn����d�u)��0�=aeJ2e��r7��:S��,�E�jX���0a:�/:6��9;	�R��=d��5v�}+����yepQ[��< r�^S�f��`�}�3��2�PުE��6DW���#��ݛ��c��M��}�R�ʹ,S�dX�P�C'�_j�pt��P�W��t�"�\�g����R�WO�cUPA+�Ϣ
��!������<d�8Q��ҍp�AO�5"!,c}�:9j�mQ��\�}���0$�����;V���X��U|�A�:�J�����c���^a��3}��7��8QU1�bzP*�+s(�B\�'�g(�+�)kd���&��Rջ�B�Hk%Bܣ��uu�ӆtGdR6p�(.(��ܩ;Q�q&UX��H�nu�PW=��9�i���"���?�k�:b��|��Ç���Eg��&o���tUk�@wy{��3$%=���}
�P�������3 Ǵ�	v�IL�6om���ןM�Y�Z�������.���\$t�	΃O��<k������ʫ�r4� ��=HF}D莩y��\υo/2��	�m���|M�j�u��hj���.�N��V����4��.7<zr]���u�2��=�5k9��ʔ#�-ۢ����_�M����Bc����P�Ȯ7òY|����K�.�QMԾ̒	.�������뜺N���C���:� a��r�� BS����yp�pylVߧc�<�V
K�*1"0 E_u��)�����k��`�z#r{Cz{e�$�v���E��1QA5D�~
g�\�a&��3j�����dXȼ�*��9�B1��:�b�J����dH(�C�aB�}$��?������凌�3�ś��S<J��K�{}{��w�nN�`���IMX����UեW����gu](Y�#K�y�=U!X�/j���.�r�̻�0�8��U��=Ak�A����^�8Ay<�Uh}����K<��;�^e���=��������N�]T^�@`a�e��2�Y�[~+3�m%���Y]4+�X[��^���Y��˜Ȱ!>���LpI/iϼ@�cB����a�͉߼ݩ/�)���z~v6r��'���,�C�r}+m��k��U��Ӓ��2��[�I�v̴�۷��nc:p]P����0h�8=���\���5D'�o�o�t͇�׽7�^�����Y4�3�L"ұf�9�� ݇�~�7�*�M.�d��9u;�gpE�!���F���#��W����SΛɂ9����ى�Ļ-v�4�u�N�{�����8]o��vV�W���2�����P���n.���X��Ln�$3���ˤ@a�p�����m�k�n����ω.�r�\������⺵s�͂N~5C�0��OO��ܮyX���L�@T�ꭓ���(�X�6���n��{�sw{��i�@�>�t��{`���[WS��G%��9r�	=���^d�
���9�ʮ��󍎥�R]��2���oe>ҹ���R�����,` ���B��#�}�{e[�U�-Z/�z������SnV]z��T�d^���^�ܺ�\�e�;�Oyk��	�m#n-*h��C��,�=���48e�L�&[�Ϩ4�P��6S�޽4sz��X;�~4��n�N9�:�u���#�+h�T!�&@�TJx��M.	�|݉�m�ù
�)��_�xusQ����_m��s�{>�FB.�Q��qFU�e
��l�`v�t?IX�D�ە8k��_�f�8�J߬��bj����
ˎ��#ʟcq��[K�w�����ȃe�̫6��L�#;�#����f�
�jfU_/S_�_��]c��J�آ-�$�KK�8m����j�::�����u��|���T�J��Hm_ /�,`����W����`���<�;�e��f��hgõ��U�{�(	�f����CѴ}(�7��Yy�Ҧ���V�zAvW1Pمs��B~u2|�ؑ��Ef��4�Hύ��b<�j��TtF`���{Ht��ძNG����㍃�-���������$/�mh�b�	Vz�� f�Ч����e.c�P��k��-@f_��:�;�)�Q�O� <=U�M����Z��㫶 � ~k4��b�z�|�~��	Zl9>^[�
!�l(���;n�g#B�:ْ��yG	U��xF��m҄24�b$#��*s5����拧} |��gE/
����N�*�i�!�=J�qb{:���^ɍL�J�]�L�'f=>�@�Tq�ᶓ2����x:w�J�����w�݋	�"����b�kԎU�`�5�s��4Gq�ܚ"K���|]C]��)L�;ܭ�̝��M����%Fݘ��p,Ǜ�C��s�/�H�����'\��lEu",L�'`H֭$��iFrx�Q�"��Y��iiy�����<>�b5�a�cA�����,X��ʊ�2���#b�X�݁�X����w{��4Dl`h���FVH�._�z���s�{O:�D���w=�x�kE��Ө*a�ZZE���P�$�m�ɿ+�u��ޟb^=^�J��2�����v�1i�V/=R��U���n*�jְ�	��wz�&�(�a�7�$���L�!5����������)(kM�cZ�'�71�q��\�9~�5���	��C�M�[��%\�꠲(�
���\����t���v����E8�M��y�֭�P�z}��8%�y�fw�ʠ �[�}�QI����2̦�Y���o��aU�[����1�λ�e��J���g����l���6,)0��փFfz��9E
��G|��)��(�����L��8f�_]��O/�1I�a�bD{.��y���s�>њ�E�:�Lb�-���&�@�q\�I��m�S,��D+y��'vܭ���Ue��:`w�p]� BWb�ݷ���3Y�����6D8��@��E���~|�Mx�O^�e>�un�y���W�3�b0 �>}�;oG_�!���P�W�Uu��<K��Y��'�?&�HWh��>DQ�|}��ms\c.�ܟ��:��(�Z�T�]&;k>�@'� }������Ag�w�iRb|�����0��!�湀i����/�k����d�,�|��8��̓L��X�=�hi"���O�4��I��u��������5�λ�_����%g+��>J�0�����I>B�a�ֹ�g���Aa�k�%xԂ�s�q�z�c�i5�O����O����
m
��M�ì�>g���7ys)_3��;4���J��q@�<D�i
�{<ֺ�Xx�eH�����:�����X(J��~�����I�+�}�����g�ܩ)9ˉ73�g*T�o�f�X��{�2�����&v����ۘ�W0�b����摐��Ns:8@B]�w��e��)�)gͅS=��UD�q���g���[��.8Cl���ӫ���{��؉��U�7U��8���g��w-۾+��e̋%���Q�.���Xy�g���{�;�Ӵ/^���È�z�Z����z���7M�@�+:��oT6� �~a�i��a���i�>C֡�;�01������2b��~�v~a�oX'��1�>\G�+Gĩ}eLvf�7v�� �R(~a����m������o�B�a塌�:�5d�{����PX|������ ����4�:��?s����N&0ǨwT����15���|�>�꯫�'!b䦮߄q�L@��Ld����L��*�A~N������K�u�B�L<��4��T���c�$�
���o�
��2�>�W�7�f��K�&?&��&��{�~���o����߀�� ��?��Av���0Ӵ��]Ͽw�ri��f���&& |��5��&!P4Z/�|eH���I�
�OœHJ������'�>�>ﲮ�_���}Β���Q��bπ���M$X��q�<����x�̕*N��H-@殟�:�M$�9�n2�Ĭ-���qL��OP�T���6�!�mbȼa�ζ���~��o�?@<n�k�?3�wz[����8��Vz�S�b�^���8���'P�
½�sXAH��ϻ�1���w'�u<�!]3���1�C��}�owr�0*Z��x�AL������?k�]��ξ��'�I��c�a��OSc�z�H/>L��;aXk7�3Lǩ1���2l���?�y��$�"��������
E�3�x��B�L����u*��'�_J�����ǣ5�Q�6|z�{7��OS����o	��T=k&���K�&:w�� �`6�/�z�$�x!\AN!P4s�۶Zͳ�g�� �b䮓g{��(� ��������$��B͹䢱�&��eB�L`V�ĕ�w��̞ q*��wD߷�$�����_����b�S���3��*|��;H-I�X�a�u4����`W��_�C��ٟ�+��<���������4���=f ��T������'��<O��ԅ0�f��ki5&yCO�L@���4ì+��>~��J�_���*
E�������AA?��SM�2��uǉ�95[����q�.Z�rY����m�޴��M�w]<R�_�sjǔ1*��X�2n*����c��R�+������g8�a�Buf������tu��ϗG�o��
��z��Y˚��pBMҒ�y!<Q�B��B���}��}T�9�I�;؍�ādD�4�#�#��?w'��������4�ɉ��$����b~�p>�z������<H.�<߸m�
��|7�I�m����z0�c%e~g�s��}��t��>�_~��bO��(m+��R/~���;g+4�o�M�z�>a̧�~`T���������0*{�bE�J�>�s��������i����!$�Y�w�����l?��{[������̲!� �"�>~g��4��P8����`����ɏ�>a��������񁶡ĕ�|Ɉ%yl�%��!�;�Pۦe�L�AH�I������l���[{̙���,`����bs'>�<	�>�3z��Aja��=�2k�1��eC�{`iă�<�3h(m+W�f>��>��$�>C5�=v�`u��g�=Ci����Ϲ�߳~���9���Xc
��'��m'�+
¿xk\wAH���:v���i����glǷO�
�3���{�Y��Av}C��|Ϝd��d�*J���'>�d��D�>`�q�uZzx[����W�y�����"������WL���x�%̓�����7���x��Ro3x�d�
��8�ϙ*~�_4��T�����L
G�^>�ϼ�����G�����SY�������ߝ"��:s�L��0��p��x�]�s��P�uH?w���8�f��%t����<5��
�R�{�1������0��<O�F�Ց��3�GVo|��Z��߷���i�& z������X�f`q
�̙��y��6��b��|þ�6������}��$��1�é���8��P�y�`i����#O�	����W����ߎ���=�>�볲qĜf;a��$�=M�:ԋ�u����=tɈJì+�HsZ��>B��j�m��nsXm�_�+*y��ی�L���{�O�
�3�k��o�W�����33�\���3�6||ğ5'�ӌ5�3�+�O�SI�'���������7�J��I���:풲�^��@�+%e�Ę��P�}�4��4Ɉ,�N7V��t{��m��D��>@�*$��k�O�7*OZ�~�$�����O��e����վ#�rۮ��h���s��jz��4�D9�}��A�+�u����]�J�t�`�b�1r�|��"�f��-���ʒ�-G��0E�]��x{�S�z�[k�#3���Q�q�d��%@�*~��I����X�!��O����f�R/�����c8é����ښH/���Lz�@��~�f=@Z��B��q�����~W'�F����w�7(��q ĩ:_�x������6�^��|��ڛH�u*Mk�C��z�Y=7x�Cԗ��O��u
�̙�N���m"�4�v� ��o�4�I��D'�QK�c�*mj�|�&vU��-M��w�gO���Q������ s�)��0�6��~��f&�i%w/rjO��h�{۳�=H.�~C�R,|o4��.��ɉ�����a_�'�4��V߽��^8��{��~���H���|0���!<f�6�P�g,=����/�g��	�잲�0/���ԟ���5ܓL�*��y�G��Atɹ�0������2Ch.�T;�5�?~���=0'w�Tֺ���$}��z��(�� Z䬕5�ٷ�u&$�T�B��'Y1G��4�����ܛg����4���S��`z�q��c�톐R/����k�H,�K��y������';�ň���g�<	�>��'�Ğ�_�,�)��1��`u������6�R��Lx�`��ӛ�m �?�<>�x�ʑ`~jy3�9��}g+��1�//o��=��`�W�݇k_}qx�� A�x�Uc��Y�f�\H,�y2�LI���)�������� q�~jJ���=�~�o�i3H(i�Ă�'Y�����~CĂ����ݴb�����c>ߚ���{��'��rΦ�i
���ɝ͠z��W�f�
�hV�XW�Af��:��0/��Ɉq�;g��&��M��C�Y:������Aa֤���<�>�s�uϾ�+���G���x����op��a��cϹ�w�C\a_8�%egk��'�%d̳3i1%g��H��偉��1"����<�Y�J��}ѷ������ﻳ�Yˡ�E�z̖|}��4��c�{���_�����a���d���A~��R|�&w	��PSa�}������4�3�1�O	�!��V
=�t�Uq&K?(&������d枈Hu�R�u��	�費5��4���iX��֡�F�|A�Ef�L�2�u�5eL��y����DJ���*�Kӛ�r����e_�_�@�1q���˦ʋ��r�b����N���oe��V�5jʱM� ����B��q��"���κ\n+��$��U�&�Kk��t)ؙW�Y�H#OX��H^Ƿ�BS2�[�ݨ�������_��bn�9^�bJ��GG;M�y��ΓȽ��)p��!��#�U�
��\]s�dx3�.���˧�Mmk=ID�o�2-b���]�4	YͶ�/Z�|�{���^ةČ`T��Rv��\�^��.�������D�,�R��E����;Q�dS��"*�-*y�����s��6x]rp(�<%gNn�jr,��j���
ԉx8���\u�^�Sf�#SE:,�Y-܉N@m�6�&5����g+U�v2�Iu�AvC��ѡ��&�Wv�k-(�(��{35fh@�E�r,,�9�mȺ*AE��]�5��v����|cOU���� +Y�Z��5�F��+ug_�9@�ŜlZ�gJ���s����kF9K{GL��8���_KN�R��@�B��9p�@T�k	;���(n.SF��?�m,��滙y8�9۹Fm>���D����n�jD�{}�}��[�$�U���Fu��A�����O8bąT�����Ϥ�Mԕ�C�F�}k��.u�d�rE�i�u���������}?0�x~�������J��ů5ϲ=�H1��do�����CBr?b���T!�$
�VQ�mx�:;z��F�V$�ϝ#�:_��v��k����5�/�8U�덚D�K��lG�  ub W@����4|���5̾�ѵ� �x��.�(�dv��:;�" �)\�Bb�m�0�u�L�ǲE���N4����.�V�>���%@G4�=���������U&�6i:I�4�����<Jdf�Y�h�&�WQ��$ �
�x��|xb�Rtd]����iA-��,��T@���KoNzp�;>9��A��^
^e؛C�1s� A��+'ʰp����Z� l��u�^q	�D� �\�@@�E�Ed$��*�2Ѝ=ia�i�R[vw� �ðyl�Q0x�:^����b"�h��X���
����ȃS$F�E�v#0W���@�L8@�*����ˀY^H�\�\� ��0��,V����U�d�hdn���	RHa��@�{���r�r� 9:��I>��P &#I�]B�8���z�����L�������;tI�d'4c^3�n gF�.�(>pwqGo�N��7�f����lkH��4�.�p�(�3�"��y��UEAdQdF,UTdb�G(UV ����P�b�#UF��E�[[AZ¤cq&�T��,��UZ�*Q���T�@X���,�Q��(
��T�UDDQZ�m+�����b��)"�X���1�`UT��V��Lˎ�`�U���(�R�A��EĪ��#�"�X���c1X(1��U���(,��0X� �AH�TV
�*��,��b�-"�(6ª����EA�������6ʋRTDKJ�%�P�VA@X1H�
�EIQ#h���`UeaZ���2%���e����	��IFe����ker��k8�n�n��-/d���3��yP��[Aq���x���E\+�=����Sj��Lλ�UJ�z��T=H.�A�}eH�?:0��J���bns�E4�䗷�{;�CĘ�g�3��ǌ
���;����Ă��z�J��$�>�n������<	�� ���O��_D�os!zHJ�ơ��L�C��Oi�i �I��7v����$������H��̇\I�
�������%g�M�}�n��bM�XT*�`T����D	>,���}�uQ�����gk�N����W�3*��Κ��!�L
͚���=�Wl=�1��I�z&$q%W��J�H/Y<La��1'�O:����,�YQ����=dDAu��)��#�߫��|��[�I���I�+�5��P_���u��R|θ����6�2T&���������N!^��|��1"��>��Z�Y�h�C]�m�4��g٧����~>�:��f��)R�ϻ���x>�-C��0�
��d����Ϭ�m@��$�
�
�MK�C�>�����Y?j�t��+�6ɞ{�q4�`^ݧ�Y6��V~M�XovO�� g]f8u���Y��I��Y�"kw?2T�=~M3�d�L
�aߺa�<H-@��b�ʆ%`c]}܁���|�!���m �I�g�������{�<a�ε"��Rm
D�"f��O#4p��2~kw{詴���=@�Vi�٧��I��솘i�`,�s��E0ӏP�l4�2T=C����� �0+��p�ʆn��Wi���H��Ƥ����Yԟ�ig��H�<	g~��7<�k)�ۻ?|w���V>!�t��̟�\M����d���ɷ�1�S���L��:�x}���P�"��u��AH���5��q�l���ϻ�R�����'��� ��c���b_V)�Z����}�����:`T��^wRo���>�^Xm���j�^0I���� �@Z�%N!X�n~��xΡ���m6�ԯ�V��O�2o>�i��G�G��sO&��%<�kO�i%'�?gp�J��.�>��X$���f_�
��������=J�2T�>}M?���`W���~N'��7�<eC�X��Ґz~�U��+`��|����[6�z q���+9b�>�1ә����.W��W_��]�,��^��G7oz��S��I���f��mT�� �2+�&��9�w�o����q�v���P3��ˎ�ܰ�����:��Wķ�S�
���D�ýB&���߀��=퉬���|�����<OR���C�|�2l<�M?0��5'�wZ��Rz�O&wz�'�J��~�4����8��SL4¿[|eH�Y>q�}��J�2T8E��W�< � R���7	S�n{�9������g�oVO�]��@�?2��g�I�!���f0�1���3O4��!���c�'_���P�Ʋy5�&���L@�_l��~gc6Y�4�A~N�������~Y�i������}���� �Y��_���J�+�z�>d����<�I��!^���0�<x��,<����izԂ����ɏHo\�i���O�5�5<H/�Mfi�E�Z��{��k[9�_�>�Ƙ[{Om�>����|�|9����W�T��f$� ��k�>a���"�X|��W��<��
���xo��$�����f����F9q'��3��*N?��C�Uu�Y;o_kn�z����Ls���x�Z�.�2��VOӉ�q��`%H/�:�!�|�0�~�CMa�����01�<B���o1�Y�����v��;_r�U\F:{r��w�R�:��'�(�A��Ԩ)>a��ځ�VJ���S[�+�����8�5d�~q�PY�*}5C�?;H,��4�:��?s����N&0Ǩvj�_�?&������b~޽��;iÖ�3���<�1�9i����& w�p�%ez�$��	PĊ��g��& �Rk=��l�L<L@�*~d����2�q
��&��5����Q��!g�[�]�P�Ν����X���f�޻�|�}�c�i:s�O�E*�u����N�����H�+�k8ϐ�����ɤ�i^�X)1
��^!�:AH��8�I_Sѓ8��g���7��l�ླྀ�Ğ�}�gY7���g�4�b�����9�vO���a���� ���6���Ă�߷�m�T8���2i*A�g�gjx���f���&��6@��C߻>y��ܜU�����{��!��^�,1�=M�{���1�_:�]�c79̝Cl+
��y�`i"��6}�6���������O7HWL�s�&�a�9�'�iW���@'�_���I�����.�]JW�U���u����s�&�Z��P�8|��J����Ѝ!��)tQyyU��r��Lra�+u���2�G��ӥ�)��{/�E��V�U08��'C�E˥�v'2��9�cv(�!�q+Z�S�º]��Z���%��?ϫﾯ{*h�ma������|̑�H�Q�I?'��7�=a��8� �d�g�+��Ƴ��f=I�>gS++�Y:s�x��*E��������O��%f������=�~�;�n|e[�Ғ�5�@D���E:�����W�����<0*�xL|d��d߶c8�{d�O���E*zZz�H/P����6���B�z�����g�� �b�]#����g�i���Vl\��Q�O�$z�G�J@�	>���w0+P����������C�z���<~`T�����O2�`T��v�~��1�d�S_�m��AjJ���I9������;��p�J~m�]5�Y�p�D�S����I����1Ĩ9�;���x��>C?!_�=C�9���`cRo^`i6�d�{�a�����8��V�l���R(u�@Q�U+��fWg�D��,��}{࢈z����
��ẁ�����3�<�;I�����rz��N'����1����7�!�At��p��������i����{�
u�F�����2���-ޛ0�T{^���%e{a�4�HT�|���d����3���J�>o�M�z�>a��%~`T��������I��
�{�4�q��k�wP�=d��~5x�H/���9�ׅ�������_Si+�)�
ÞPӦN���u?&�1*����
M�Y����|�YSɿ�4����O!�����q�>J�g�?&�0*;��4əx�G�MolK��#Nm�%��?y	'ĉ����o<d��k	�||H-C�n�OX|�M2y��^2�Ծo��x��Y�(q�@�V<�ǉ:�C�~OC���Az��1�5�=v�`u���~x<������N�G}���w&$�iĬ1�~t�нͤ��a^y�|���CG���Af!�b!�glv���8�ڧ<��4���/�qğ3�>=�M2�����'�LB~;��U�Gnu}�=:�>q���w�p��$�=���g���
���+
�<I��d��++�l�{�x��R[Ax�d�
��8��!Sn�1�T�>��?;0G��x����֬��jw.����ٞK,�2��Z��4kZ�[��o�.��d�g6�E�h3Em��c_�������_#R�����"�=S;���\�ޙ}\�b��m��/�ڸ77�����-�p5lt�.��w���Wt�u����n�>�g�nb&�)�K��h�4P�lp�P�u:_n�7fQOm�����79�u������G{j&<  {����M,�c{<Lx��R��J�;��c%��}��Ԃ�ý�[��bA���T�N!Y�3�%t����3?`T
��tᧈV
LB�(���Nk�A�s���C�̿���ԭޑ`m��:}CO��L@��j��/׌O3�V~d̿3���6�X���掾$m�Ûލ��I��}�v��u<M0�+�
�W~г�(��/��QA��-S�xqs�����!�=@�Vw,����1S�JH/Xz�5E�d�����bi���/ﷰ�m�XW�H��*VO{���`)79�6�;|H,�3����@dJ�z<=���4z[칚��2�)9U?�q����{�@��5I�0Ě5�Hg��|ɦh�CMd�&�q���'�<a���083HE�~�r���w���{�I�Ld�ɤ��\g�</��~3�J�ĩ�����a������~�f��n��!�����Ϩm����Ϭ3T�����~½@L�w~r�F�0VM�9�N�^��o7�6������t��j\'��߮±���,��c��V�%^/���{�O�8r�s��z;�<�T�,ȸR���=Y���33�1��80|wܠճ�fTg��#����o�j�:������tz���F^GcVG0�ck�9e����T��n�mX8aօ�2M����*���Nm��������}�Z���X^Áۨ٬����fI~�dA`�R:��@`�ɒ��D�@}�E��[���@��;vwv{][Y�8��Z(�?f]eGx�H�>]s<
�R��N�$q_<P��(9j�K��]����Ǽ�<���i^��P��� 
�h����Ί5	Ò]S>���P�r�P���K�@���$+��"L���'s1���/���.�,sݱ
uS��<9Aõ& $�|G���P�>t�~���.�c�]-�X�읲�]!��r�Y�T �%,��}aa�k��/#D:�ؠu��Iv*��|_�(����7&C䄡�T��8=�K���t���2��Ԩ�G(P�(F��'ďLyr
�x�ڻ�8��0;X�8B���B4��냵P�����i��]�DoF��U����$x:b�7�_I�K�0dDn���!����゘�p�O��.!e�|O�*֍0*w]�޻ً�e���J��M�@�y�H�W�HDk�D�veFx�$9I������#��v���#9W�[���}۔#�a7�W�����]e�����]4r�Vۋ-�"�D�˸��S�����p�d��*b20��s��o�W�^�ǯ��Ad���z-g��s��:�D��A�W��>T�t��\�(��f�R�u�6}e#�^��Q"��H��.X6�c~Y�3��u�	އ�gP[��X�zޤ/��ܤ����>��
NT��-a���F���'zN/���g ��N�J9�f��rV=�bF�v��{|1^iRQ(^p��:��˛����sjr���5�&��1v]t%��{�x�8��2#%��ޜ^6�10�~O\#jf�,���:���b�ٿs��_�x�/j���c�1܊����X�{�ğdo��Kt:-�Δ��>z�.cX7y����"�ty��^Q�T�X�V���:��Bu�׹K՚옚��J�!���z߭�{��������/��QW��]{Π6��9s��]����q�oWw���أ��C�{�N��A��R�*P�|�a�-���yjv֪֪��/w��M*�u�7���Ih�� u+��C!WDn<k/Q��@�e��dj�6�{Q��^=��˵Ğ5�W�FVԕ{���ľ��;��3��DOG�����<�#�#�d���'��w��ζ�jP},k6��j�ti��l�g��%.��>ǻXƷa��wIsW�$�F.�x�9q���-{O�1 #�O�q}��W��Bo�˱\J��U�c;�Il6��)�Yҳ8���q�S��d��ե�O\��$�V|�ܶ�h�L�@���𘣤}��§��J��f�KMt""�)�f\�uM�/�il�3'N���*�E���m�;=r3~����[U���Ml�æ�:���n�T"�*��Ϊ]tu���wO�1߮��������=~o�;y4�\���K<������a�^�w*�ΡP�aY��9�)��<����@�/��'���*�v9܍��m4boZ�@��3�gz�gQt�g˘N��n��`�P�����{Y���ݱ�g�H�_�-�q�]�UZڡ�Z`�	��.c�7��md���L��z\�������	��+��8��������W+��S�Ϲ)V��س��Ʒ���`ne�`����{���^����Bޠ{P���a�[�#V	c�(�ƺ?b-��&]����j��ϲ�;�ˊ�"�\�M�+��؆-˵<,��oV�	Z�����GN@�ɏ%\8*Ó��|�2�e��G���R��r�6��~�B������[B҂���f��`�{$��z��� N\�'�}M\����w��d9k;�8o���3Vv���D�#aO�8b�a���WfFf+�ف�c��U�7�`P����]��	��Jb,��h�9<���M�,ar��>̮��2�ƌ�t1Λ�t߁]]�f���^��3e�{w�~���T�|�^�,���=�=�)�ʥݱ�^��Bs}7ނۣ#8��y���y�6���B#�W�r�\$�iH�J������@�.^5��45��ɵ��GS΅��T#�M�T(w9Im����ݸ�0W����m��VTX��;�'-�����
�� ⨣˨]v�n4��������Yf.��ż�߷ :�4r��q��ތ8�:v������t��������R��ken����v+��R�W�i˫��b�`��g!�m׬+L��{�e�I���
uȂ����K�ˬ�ݞ}�h�?��m�*��x�B��S���0��6�9�z�gJ�N6�g�1	�f9n���&�a��}�T�2U�B�dE�T�9�����r�6x_��Ďo��v�~�>e�X�Ԯ&^��3.�to�Zt���V�µq���]R��|P�����ϰe 6۹4��\�V��Db��E�Ӝ����p����|PwX���;��O:U�.ƞV6��oU�k&�f��v�mf�9W+h֊�04���Y?}_U}Kq���Y�f���5��zU�;�.��1�c�7�T�|��Z3,zǑ�/�o�N!`nW���
c��O"�v'�QR"����a�Fߟ��2/Qg�.�u��{�F�;5k�T�n�0.Ùf�{�
�S�ܥ�M�43�~�b ��'��Xq3��uN�HyOR��8oݥ�ӌb�����I��{�NP�y��1|�Tj��aK؝P��#�U8ȗX�T=)�珞�<�sq{Qϫ��i󂊤�MpB��+�	\]l=�9���X���}�jٹ�~�۶{B���	58����=ϳ9���l�,}���R�9ٯ�P�ݿg�~Zs[�w�\)
�J�l:�ᣋ����UJ��`�۞>�����z�7�w�N�6��<�5a��r�s���Ƴu��7~��f=����+#Yt�.�JOOZg'��ˣzWv���#��������[��-/�Z��.Ű)���w�S����Q�OE�MA:��7��=���ŷ����e���1�f��L���;�����z��)U�;X��w�\YAoKyu�A�P�F6�NrӦx�ݣU����)l��{����D������mն�����5~�Uuφ�twu��7��ЯI꺷�n$�w�������u��6
��i=;�*e�]��I�'��h��^Js�{f��ep]aŉ�b��"�k��K��3%/LW���	�i؞��;@򹲔��٠-���m=�i�Y�ܽ�$�	�v��湍@����1>�j�J*�;��$7�*۬�����݌(�����|�L��?x�w��6��Jg��}���߰o�{*�a��k'���vX�C�٩YZ��r�1�5څNy�K���0��!{�5��t�$n��ˌ��7lC���8��7�����'�\~W㼻�s>, �z���{���;h{�xp_a�ƴ5e�ȶ�'����:l�J��zX��]�Ǣ�fm�î��G}�c�%o�Qh���o�ɵwi�Ԭэ�3ų]V�q.�ޮ�5��*%��Z��\�e�.�;9��1���^��\G���EZ6�KŚ��o�׀�9�&�({���J�.�`�����ȏ���#o
��<�5�=d���1;����v�]sm��].[S���W^�[E��*�2+%���p"<��ūRt�{�A�z�4q�����y�.���[��!I
��mIM�Z/���gV>�[��bE�V���ۙ�ܘ�:Z�*��W�7sRS���Y�8�uG�b7����v�\�Lou��� ��J���j�%7�[n�02�MK)d{�{������S��p��(�0��na@LXn�rWFT��0��]�V��}�¬̖-�]��̙Y��z�\o1�z�5�����YXL.�SOڋ�a���tq���
��ʎvu��Z��SAr�'vv!�=+s�0�0j{'9&۹;4(�tQ�CnT�|k=��o��ێ�H�H�^gSN�e�v�L�d�k��Q�"萓����bU�|�ڼ}|�����|�P��g2�"�{k絥���*�u��������ܚ��r�{N��ګ���k��V��p[�7�u�#@��;����x�*��S*J��]+t��u��:"3��b�哚@��m �U�c�����S��
��Ї��ca�Tg|M�>���P�߷�u�]���0h~��am�w�<�t=���gy*hQ9x�'o\jb���6|�3�i��j/�!Xq��W1{Rs�LO	�2  j���*=N�x��N�rɅϵFm�k�C��&�H(t�ʰy��ˠg���y�®�d�qp��>��ڷV��v�(J2><{}�I���`�ǁR��Nq��������r9� Y�ɵ�m����:�Uva�x$�a9�f�m{���Ng����/Ȕ�Ê%ޘ����Q	U&A���h+
�*�21"ǜn�x8`!j�Z2ۺ�X��h+�X�ǞF$*#��N�`j-:b�7WQ�����V:U>Q����M7&�(�/:����<�1�Qe�v&u��AةKv�{Q���K�"d!��E*"�suS��e���3mۚr��5�$��Ba�x����4(B�`��&�^l0���ЙˣQn����Բ�ׯP��	l�q���B��mjݥj�)��	Mסة���of�� ��1�/���g2c|0�&\# b����P�{��]o�K��{�?EX,,��`�*-��B*2�E�(,����֣,j��RՂ���(��VUJ���.%F�m���F6��D(Ԉ�V�*
(�1F*E-�ʕ-mQ�\LdXV�"�[���B�EEdRUeFѴPPX"5,TXVm*сm�mE��,�`�F,���T���X��)h[J �T���X�Z��eYb�kE*\�0�R�m+(�,+�j6�rܠ�R��W� T̢2�q�� ��h��J��r��1F�ܤ����Ҷ#1��"(UEZ��[K[�l-���XT��T�(�[a�T�U����JڬQjJ$1�#�
�h�q��.ZZP�Lj�KkK!X�DQ�U�������h��ξ'�!y�ۭœ�	v�Ĵ�뽭�+!댬G�'�_gs/��m�<�h��͢�!ܮ�sc�Ev���3���;�<Ho���§��Rj�g˦�5�v�3��;z?����~\����EЩ|��ځ}۷��l4�u�c��U�Ð�sk��z�,���Bz܋��u鲗l���CZzo2x����k����wGf�~=�^��q.��@8�-|2�Tz�jҍ�Ɯɫݷ�әe0���m��)d�׺��0X��ی����6���J�t�]Ѻ4�����A�ɥR�P�+�����*�ыj�a+}���/��y<�,��\���ݓØO��M������>�V1�=�-�����,�Z]̏b��,zv�s�N+��0�Q=Z�	�x�{|0p�`��+�OH�k�c��ꅵ����v�XF�!�5���)T�t /���>��~W��tOq[��"|;>b+ۮf31ME�31�n�-sf��(����Cpno���N��͖�LݑQ�F���Vf���7RS�!���n�Bݓ�78�����[$ɒg�xvNܖ���{S_7b���vfqM
/J�qj�]�f�u:ؤ����m���6�>�s\��^�s<�P�n�VCB���� u�[��cR�����7�������/uؘ�|�N-�Լk�hCf�ͮY�vgez��^���5Wy����\�9��U��0��vPsێ���J����O�ۄ�.�O��ޤ�f�y�R�uf����o21�9���1hs��[ྜ�	��ir�p���f��?[�L�or���N]��v���o��HĪ�Ď���	<E��+�^p�s�Rwf��Y&_��9�+CSy��Oc�V���'�*�K:�FvR������+q�|켇^YТ�h*��Z�s��]B���IDQy���^*�9����Ḭ�K�;�ޜ��7`�4��B��C�r��yv'��flĎ}sk�;wR��cr uJS�.�|���ކ�$�����7��w�J̺p5@n�m`<����Hv�h*�F���N������%M��R����_I�t(^�M�%B亽 �D���/U�M�ݱ�ǂ`��S�{;S���+�+��J��,�_�P�z��V���cr�u��vV@�T���u��2R�rt"_l�·�tֹ�3{z���{�{X��ʉ��ѥ�1�J�y��p�=:ҵ��L�41ᦳy�o��I�j�M��c��z��;ۓ�v��ֱ�9'�O!k�6�N�{�������g?[G��ɹ�Q��bܑ��`W:˞���7w��pLu3��Y�i(����O: ��q��B]��ŏB��
�w3����5�RD�v�4�����b�ۘ���W���������t�dً��. v3Ϗ�L�c�%<���l^��5GI�6���F�g���`ޠb
�z�-��z�T�!�C5u䮡m8�C�^��x��^o�/�[���^ޠԥ��u�u���@����c�����JgC�w�I�]����e��,»��nwIvuE{�qk���%Υ��_�7�ǈV����ZW�����i����xC�ٔ\����'^� ��n1�(�W�������6qy3�N��:WD���|�q�Of�
��,��B��6�u77��1�ބ܂�Ǟ���x�Ŋ<��Ι7<7�Pz��+�u]�*_*���+l.k:��T�]ʛ(kt�p���>�=[��&]%���3�����B�-�6�r�u�HXS�]���S{kՍ�vĎ,�4o9b_{��:��s���&��vmW���|�ס_+=��P�H#����j�%���Ȱ��y�s��r}Z�f�3�w8,�ZrCtݝ��V���[2"D�R�*TU�[��w�\ �{�koU޳�;�N�b疫��Qy޲P)D��6^(��:��֭��w	�*��˲�Zq��эW�zz�9	����i���N�-T����>�����(`W#��ׄd��c$e����O;�wB;p��f|�T���h���#��xG//c鋟�嬃�����g���r�c.U�;�SbBb��"��_U���^}Y汱4!�=�ٽBn��b��/��vAr0��w{40|I[�@㛵��,g]��Ǯ�Yr�.I��ݿk�3��#��d�V���eP׆:]@��R�-��P��4.|7�6C�c���iyզOi�w������F(zٰǱ�Z�#Q�� ��gG�������;�tq�#0[|�qnc��j�0i�P��K2������|C8�-�N���7W�pL�y�8jPAvwS�0<����`�[L��Z���X���:�u��3�Vxz�soFE�;�4�q��귨�3{��6���챯2!��Us��c��@����^���b>�G���$�����������9�
�V����bj_XB�4{���é��N�=�S�S�V��[8z�yC��=Y0�ۓS��T<]-�ަsX���y�5x��"9{OO�#{�Ǣ�fm����B�\�x)M��SQ}w�v�)h�4-�uY�tȑ�dϮk����و/+��`5�U�y6x�W7����Μnt�=dlҜ���������WW-O�,�՗ƭ�%7u���Ah��&���ut�_�mPv}|1���;�˷��c�5����^�S�_�);�XBTp�C�N*�<��[��J��� �d�~����[fc��O,7��c +�d5^8R����W�cg,�G7OoRLҩ-Zڅ�sm�����׹(�֡��A��}�/�uۗIՍڈ����D>'�b���ނ��O��Q�!�ju�4P:%�����2�7F.�+(��t�uI�{�;�k�K>�]���SR��pYN����N�f�O.|�\�r��|V��8.�]��c������uևL;��gq����
≝r��Ӄ�9�����`����fy��3�ѸW]����Qy����&��Mॴ�����<�j<��;~g%g���r�k���W�%);+j�7s�wz]a�;��Ɇ:�`�ybU��'O;iq/�����\�	/�n�W:�#u�.~oD���P�ps1m\�bf'���>���$H�<w����L}���d��J�|,���g˩zi�x�wy��N6f������SJm.�~T�`ߩ{"���n؆.|V�q�646��"���(Ȼ�3ܩ=c��VN>]�|jy�X�M�Er߇�7�t�m��n1� �qe������?�&wM��7�H�Fgc�F%��w��{~��v32e��ry�5z@��V�S>U.�ڎ$kd���z��7�>�lM�=����QB[p����uDMD=L�K���W��nK�o4�K|+EEB�qÒ��.ƕ�3^��|�����9�ϑR�u)��6};zZzK!\ߖ��sc�
�v��n��΁�Y\�{8��>T���n����,��l��]ݑ����^�d:��0=�����wW�������ў��a�-��/��w#�<�QE��Gp�mP���R�\v�7ޏ�c��J|�N[cO�'یkצ�:n�{�!.��;9j9dP;�a�I\�eB�}K�Ә�Cݠ����N�,�'.h��p�9/��_>�q��5����-TQ�t;{�|}:�`ݒ�T����_l�"#�$�3-�[-v����F��u�׋yC���Pw�b����7���e���7��-�V�a.�v�3�s��f�������w�qQQ��Y�7�
���2�c�	�9�8�����U�q���zx��]�K��b��G`��<g�}S�+�%�:ly�O҇:�ſOR��obb���j�U�(٬�8�#Ji��@��5�w5�3�.?�..�_��,E���^����K;adZ��S�3�특��Kb�v!>�n��9�w�I�[�g1��Q��Y4�QY�ݘ���X���X���̘(dʸ�.թ[��ڠ,s%��P�h����3{Xt�=ux.��x����g<�cm��meʾ#*N�F�۬��V�Zo���²g#6���s��<6����wK��76ޘ���ˤ���_}�{.1��{b>N�ns��ﱌu�cu���'+g���'.�~�x�{��.}"dy*��4z�T��{j��T����;^~��L�{=����n��e�{V��2��UߏZ��=rҰ6�2�)�v�Z�z�Nν���)<{�q�5��֕�WQB(��������e�u�w�ߕl��	����`�T��H*�w\M�υ-�F
i�*�]_��W'P~��=��G�F�)\��k=�����x�rk=a\����Wmo���5��v0��I?dkL��)��,�{Z���ɴ�Sw{,Ds���z	EDr���z�oO5��7�-���:��\өR+:�:�yȸ�nC��`W:��hg#U�xm������WI��㹥[n�[˕R�<C��#��xU~Y��a4K����!�����-�4��;�8��ި�`#5.��z�\��i����ݠt	�:�+Zn�Y|Xr�v8��(�-͚�7�����^@��W �t�<��p!]OI��	�ʴ�q�Dy�+g/R��D�0�R9�DҸ+<{[�	K�\+���&t�VT�[bd���*� ���!;&yۑ^�/��y�����N��j��:z�U��|�x��AnB���n�kg��uq<��Ȑ�mٍ׹I�?H���k�`�F�7�`����ݛRK�a9��ʺ��IS�ٕAZ�3���i#��b��c�^�9$�m�{�6�P��lˇK�(��ML-y���1�W�~�-����шc�j��-,�*O=�ы+*'6�`X�z�nk���6��Ẏ�!�ũ��۸�k�s�t;Cip%�����|��ԑ��b��Q��rwy�#xY	_��ٰ!\\r3Kn��;J�7��FqW���~�R3]W.Nl-�.�]r��𴠪�&M�u<�Rhn����O/�.�������*�U�k�,Wr�!_+���툫�9r��r�ݮ��2oFF���2�P�K�j=}۷��o�V��w����ݧ�QT�:ыW_s������Y�a'�o�}V���E�Ѐ$�=�n�<��b�&��rsf\FFq�/sYHl�y�t� ̽o���a�lB�On@2;��$�[D=f�QciT�u$z��u�'�+��ɼ�Y�C�Uq�׿��̨�)�h��⿲9�	il*�$ڡ@O'B�.��\t���8b�'K�)\��X�Mq��wIX�y���<�	�AU9s��Ùn��b�{�˥�؛�$#z^���{�➛�n▼�x05>6uP�Q>�W��̢���ơ�z{u�wu��3ҧR��i�QS�C��6Mj����U�ੂ���=�ڹP�u\Ӥ��N�����0ݨ�!7���r2ݼ���Mrʚ뙞RgY��*-�{15޴����ε�w3����Cw0��6��K�6�.����_щ�s�߬�/����K�t�w�75"_��`]+P�5���k���m����{�<���k���__Q��=B�����|���ٞ����Εx�G?U��=S>�7�־�q45��ӻ�8�[Y�-_!!	����NE�\�k��Ǒt��,V� yؼ��\���H��vc�i���,���+^��.\�������Y��mD���x��n��*_�H=��N�{�h����՛�	��!P�o�Y�IZ�BDn�B���:w%�:�*l���	Pr9l(�WiGZڗ%��^�K���}]@�&ŗZ�P6p�8a;F�I�͌uiC6�.	aރ��GqN�դ���`t�{���OS�2�ejѰ��T�e�]af���I����.4=�\�6���T���X$�U�g,�9��u5V��fI\Gt�K�g�V�zGP�`�q���v��t'���t�w��Vw��@~5V��Cg�KR�2�p�&���}�' 7�E�MM�u�VJ�#.��0dɛ��E۝�2!�V�vv<�z0K�פ�ͩ��;��߷	�rܴB�rp}��;�\��WgB��Y�6����¹���Au٣i�'Em�V�p���
|PE��֋�0SJ�n^l� ܓ��R�^�Qg]Y*��v�y R��pQ��$�"�������%�u��/@z�}����zQ`Q�m��jJ5��R��k���3���3U��	�+�g\y��쯸�Nl��%8����ð��:r�ٔ�::P7�V$L��H��Q%�*�l�D_^7�;vr�ȓ���ϵ]l��9Y�a%�6��Æ,�,U�Â۷�����+�Յ2�h���5�P��۵Vwk�S�q*�ݚ�B���%��o8�I�(�a��Er��Cuᑥ�VL��vۜS*�b�,|��U|wkU��9�c��M/���}��̓A�0!�8Q
�K�%��2�f\��CE�Ov��9]�� 2���-&��𧡍O8�7��Hڵ1Iw4���8���c��O���ȯ���Wq
äQ�6]ҝ�E�ێ�^Xr[�gG��#i�Nb.��æ��uۦ��Y��}�s���&q}���Z��X�ؗ�z��1�Ѯ�\kn��pGh;�� �-}+H�v; �C+q���%[��n�(Daмi,x���;���އ�!�%�@�۰�rlb����&XtPB�l���#>4y��l�^�X���2V�p嶬��BA(+���ú����\v������n1&��Օ���[hp\�I%X��K��
�Ȣ3���}R��Q��g%`�L��M���y�o�RLd�����gۻ���Y+��s|*��9g��C;����"��Z�uYL�ub�6م�#��+q�D�>=o����,��C9\�w�hVX�gemEpS����&�k�\�u�1r��7�:����-r/[���Y�[`�x/V�䡸Ψ&���M� �_U���ӛۇ���נ'�#g��Ck��\��X����PR%�W[[M�Z�Q3�Q��F+������]o�u8��G^R�!��d������f9��U=^>�C<���b���f�H�$ã�y��Ҧ<���da>7'F�^*��Z'+I�}!y�G�\HB��盻�P{n�Lo(了��y�4�	�jJ�b9v�E�r��3]S��?V�����b�K_3��9&w�#G'��T���ł� �Lf`�G�5i�P.�u�*��V��� � �'ĀE�qZ��j[Z#lA��)lQ�Q,�ZUU`�UVTlm�T�h��W,1T2���2f.d-*+m��jT�*
U���ԭ�EUJ%*YmQ�UX�X���Z����UD���QU`eZ�+kE��R�km��B嘊�
����YPkV�X[Damԡej���mk**����(-�JY��T1R#Z1+b����9E��DUե�jV�-���,J�P��A�-�UmFT�V�����ն��R���"��l�Tm�LA\��j6ԬE*#*E)R�����h[B�VUV�Z�ikEZ����J��eeՊ��[m�����U�DQETTmjҗ0�E���(XŬ-��h(�X�B��P��J��1Ʊ�[b�����V�]�}��6�]pƝ���t�S�I�����v���ys�hbڸW;Ϛ�6wn��^�#k�{X�)�����Q�PΖ�j)TJ�KP��{�0��ھn<��묗K��}�0�����lmlC�_E���{�Ru۸Vm��ѱ=����+k��d_z^�9[��.�6εҪՊ�=�P��%����T�Tk�c���u��G���k�3M$Z���(zH^��w=����X���E�$w�M�Vy_k{�w9$��3s;���$���7Wo��*٥�����']57�{���wz�̘}���KV����.ݿ��Sc�:+ҧ�VY��<A0ZP��#�G5W�{u�����b�ޜN[����vː�w�(<P�bw/��R���z���ں{S��!�����v�[AY(��&��7W÷+��;LF/gLX/n�-��*�4��x%��hƴ�����j��Z�FN��ð�7�1����1��BwaR���ò{�n"�-9�����c|��KL������q�x�����T���N݄��9�%I�"��b�`���,�p-m@�,�Μ�a�%{G<u��7gQ����H������AA+���_H��o{��9[[����J��E�]���3Y�/Mq��MT9�>�33�'T�ș�y}�goT϶/=������(k���L_����<h�:9�cP+m���6[�V{u�z�jlc�L��՜S��yK��sM���mz#=<�n��ؾv=t�CX�b�ȱ1.Fyנ�c;�y��;,F���7�)�j�����f��/d΁]B�d��֙��avE�`U䆺7lC�+TT��Tk���H�}������<�;ў, �yi[���{F!%�*���\�[���Ѻ/���V�b�{�5�o��z�(q�̧���A�*�s�mτr���+@\���
X,ymW	�^�|��ت�ܓ�#����T��>=Å��똗׊_��E����@=��x��KG�6�8-շ��vz�v%:a�v�*�Ţ���{qN��z/�WZ-��i�}(E�M�%0{6�q�c�tzqb�u���W����n���LPT7vG�̴jG�K�	J�J��e@SJ=۲�����0����[�ۙ;k�98���5�G�^�h�)�ݛ�u.89�=��A��ׯʲ߶��s�����L�����uލ���1"Q7ul�;��96��SOHa��I�2���)�꘶��t^m<nh�VSJ
�̲����u�{�6�]�F��E��l�:FT�݉A�s�һUћ�*�h�I=��*�"��H>{轉�W=S����qT�lv��\l�=��څN:@<�v:lKv$s�"�K��As�n�oe��Q��#�'�C���RBx�;E��}��cYk�o�Q7����f-94v�������F�œ]�N����ƽ>�\_t]��--gEn=��S��6��I{��x�U]e�3�{%�5��܉���<h�9�K�F��w�ߩ�x���ǜnЇ��j/1u�A��aSwP�_vJՉL�cj��S�τ�
j'��e���-Emvx��)o�F���.���o'�N��'Z��6�q�z �׌�!K�]���h��� ��\պ���*��E��mOr�F�3_3ӏZ��}�L��Z�GQO.�(4���8j�w���M���f���sՐY���nX:�����1\�-è��'
�21#[3��Zy�c^�P<�oד��D�Voo|{a�'Լ�����s���u�{�'7�jZO_e�
J��u8쩞�S���Q��x��CS(�C�=<u�wfC�:P�,�ޭ劷�A�iO��V�J��O|߅��{��9g~���8nO,�Fg���A�]</�F�vޭ��bS����I�B���T�m���hC�=�%�׼�$��Rb�����s����%@�*��E�̽�Hz�)޲��8�|t���Gv�	>*ޜ��@�*k���:�yH�í�oIs8��I�c��
���}�y2�?9jiT�����[cGd�f.k����-;\<;N����ϟ��2z�y�jlJo=��0	�:��N/%�m�{�i/)����x�;��q��`�5��w0����]�ӯz���������ه}R�4ZQ/��:���ld˦ZJ*rl��=1пw��������`��O�O�����9��]{tk4�2�i���+���^��{sbVhr*9{K6��r��om����B�`r�s���ňs��;m[�v��l!�N���׮/T��bk�b[���W��x�\sb�`�8��S�jw����h��}�|��~�=��7]�NI��y Zf-zh�\%��2ej	��V���j�&sh�Y
^��b���rsC~/1ؘ���Ҍ�K�+�y����B�9ҝ�lSyI�nߡ�iH�
f+5���Ԣ0�r��um�-�8�By[����kW�e����k���$�����vjn��-P��kskY�o8q�d����J軾�P�|�����ݎ�R�B�Eʄk���E�f�3|�&��&,T�ou��&�KE�]Q���g��8�u��8�B ��=;H��5�u����Nr���h�V�U����:�J<v�Z�Z�`�2��U�]��,�7tԴ�JI��}��@���7��%�n��dwPq�!�����Zv6OQ]Q)p����Jo��RF1�+,���7׆�,A��2Dv? ���r��Po��8;�E��S��c��f�&��<�խ�]�e�bk����BE�V&p���qLz��Ft��u���zy�\����7]��a�����ױ�vÝG3I_{�s�Gc	F<���~��k+^<u��ہ�Y$^��"�a�P;j�mL�z�c�������Zν���	�8�I��c�g�&Zw�dH�nm<�
�����z8����si��e�Q}�G�*��y.�,�L��Z�٤a���0cǈj5�K�3��巗�Fg.��
�;sJK�a_=ͿK��jAٚg��l*�>���n<�hc=�d%N��A`�7Z�	�f"}؁��Z��p��$O!�G)�䜫ݱ�H�l�Ĭ%����Tpk�&z6�@���FBXcm%��]ƅ�y7)說:�L.�6��%�z��}s�|�Ծ��m����Vd�Q���d��D3M���T�O6�S<	�>�R�|ܬ���6��x��wX�ڳ>�l�^nVRQSs������"�QU(��c`RM�U�r׻*�k��&�B���	c���^7=�)�c�ו�}�n�f����	ɮ^�S
��r�M4�}��%L��>�;��������v���d���r�fU��uj�e�q�(����5���T�Y.a�d}ٻ6�G��l{U8���=1	K~.U�֬SP\F���Y-�R�a�jN���d��_l*��f��.����p�n��c�b]\���Z��I���wx��H����2'z�iV^D��<����y(�8n�Q�ӏtY�cl�]�~[��욕�:ȷo-�a���M�ű�G:���h>5\hN󫦺�+T�m�[�m��H�|*s�o�q��)�S]�r���C� � �k�V�۫V/�������vw��3癃}�H-9<_��'�l��傪��V:���<v�c"�R�n������5R;y�㟏6h'b^��,���WQ|��a�q�=�n�_�u���g=�:�P�IߺlKv'���:K�%��iq}9/ϝ�;�yO�~[��O=��ϦX���.a5X9�1�v�����q��`-��8������~�k�9K�f*��6.�EP�{7kztٶfdY�M,���!��a_;rw�?L����J�����[�����7c������>ŉ�|<�ٷ��}�;��qW6������@[�8_ ����'{�q�b����;.R����N�����k��_����'�����Fd˫n�X:���2oݔ���Aչr)j����gzO7z)]kuz�`A;��ۨZ�����\�Cȹv��m.ջ�;Z�X�%R��7���j��{���ܣꊇf���>ږ�����m޼Q�U�X3j�Uk93#y�7w��7�d �Wc��gf"^�j�Ow�f���塴uR�Ǻ$���_1������RO_n�`7W��x�*w���M�8�S9��L��1���e�NeF����&�x�]��PUH*�t��w=��b]`îx�tœ��s�T�8�Ľ'=���s^���C�5zԋ�sSݳ�e�۽���_$�e�y��\�h�	�V�4���r�}�8�7�λ�	\p��5df�*���:ʒ�����o2�+������Jr���o%b;��֭��C@�Q{����[�Mk��Ұj*��S8��Է�_m!&*q*L:[�z��g"�����z	2�ۚ�}��*P���qɈj{OR�	4N���-֥��OA�jj�`�<7>|�]Jp�/��MY�Vu
q`&t�(�Z�%��Y׼�.��se���4s�>xO�����M0{'�U�r^�j?U\�h����ژRxu?9+�[�7/v|m���pJ^��̟*�aN��'U�O�.G������}�XAB���^���=^<ӵ6$fb�R��D��V\������̶'ؽ����G�y�R%�Mb�CU�IZ�4�<��d o*t둙�7#gE�������9�b���G�5=�&���k�eT���!�h_ߨ�w�A�jrM�fj���nFp9�Ճ�����]�C�J�r�';���ۍ�UX�����N5�YL](�sy�\�S<��\����Q�]J�\�c��M�����s}�Mʌ�'���o�a���W����+��W�F8�C�8�OU�܌u�����s�)"�[ӻѾ�3C}����k��oP�r7\��(��P�����	�V3h��t�^�!>��m^ͧ�]�-0l�v��=�|Q�ͦiJۚ��l �X�2�M�7xi�ۡ��q�[�ns��d��>��{o�������r�����y��eM��[W����ܽ�~�*��'��[PUBJ�x��"_%�6�s̠��W��j�'wbm��7*1�m^'�ɽ���T{>���U���7B�t�S(2��|bR�e{��9!�lu��;�a��nP�U������<)��0���}"���3����zVW��LΝ���B#� \��J74�V]�Г��5�i��G���;2���Ws}��9;��ɧR�s-;�5�"/�̓)�W��sD�IdS����+��K�Xq�BoS���w.�O{><߾�#(�z�uM��(�u��S��aP�c���́X�	y@�����)/����6�W`�ɉZ:��m.cP*匼�������s��c�vb'�} x�>�J���Z���C�qLv�������Y9�9G����IF�u=�e6]
`e.1���w�
��]x��[�֒T�NZlA��\u%)�عb��g-��0(EI��i�`�oeٻ����s��jmR�[Z�u�O�0m�,bS��͔Ƕe�&n������U�1yz��9(�NC��ڧ�ݛ�w,�K
��\D�ٝN֤������-�v-�j� ���{��Z��C�:�
t�S���>�ŻJ
�yr�Nql�����Mp��]��F��u�i<��|Sw�YS�[�n ���m�C��`���gZ�v��(�er7K�����F�	�w��ޛB��V�k�$��Z�;-�eoj�s3�����I.#��8��z���t�-�ϸ��tօ�Vd�����Sb��בOS�;��n[�GW�ܕi[.$�#���V+��D�ˢ��V%q���r���ؤ8[�:8)�
X��a=�g�Jk�	]G*I�Gb��;H��w�҄�%N�f8#Ọwv���Z;�mn}aS����y������"8L}�ջ�Ӿv�R�s�*x0�W���n�Yݖ
}GGY��,r�j�'�cUc���5ݹ�j�7�@��C�R8�TYfof�st�����[f�]��-��6-���ld��,��P�6U3/��Y��^�y�A6��)<,�A��%Ev�"�]o r��ٳ��A\�p�eѰpvX9���[Ι[�]f-י�'�k�U��s�úL{�Vi��в���oS��\^u��|����Z�E�ݑ�Z�q�`�P�B�
�v�S�T�"�[)J�;����]_j���3����hы�����GV�{
k[�0n�wWv��K9�8}�E������CfE؋8���p��XS�.2�q(
X T<������[�m;�q��ی>��,R-
D�GI���b��>�1�p!J!@Vam�Ur�d�Z�;�3���Cą�XlI�d>�7�|�x�Wr+��z"^0��R����?q6*3���/e��鉥BR�9ͪ#[��Dx7;|zm�Nm��v���,P�F0w]�Q���/���rC�b��9ҹم�[��pe���B��-�Ӝ�Y:�����N�S������;S��DL��ZYt��뜱W���p0ޝ�Ł&�-x�xv��[�ݱ��|�����24AIV��X���[���k�ʼ��2���������b~�=\- �A�A���;���}���c�jX��E��M��2�0*\�⢲��KAEeF�"T�Qb���[kh�4m�+
��*(�Ң��*V�X�V��,J��e�h�mX�+1�j-����--hR��cU���3r7*� �P�J�Rңh�nf���Z��Q�6���"�R�DE+V�EQ�ª*�V��U��T��*)iIh���E\e[j��Ym* �m��m���kFҪX���m���W�[`Զ��e��֋m��ň���4�D�[0Q�UJ+Q���%��J��[�0E�cTT�)QFڶ�ITC�䵩B�AjVVڵ�[B�֪�J�EPb* µ��Dc[nU�(��+RР�UYm-*�,A[q\V*"+m��QKm�F�ѭDUYi�QA�VV"�j�b�"Rт����j"�*��TR��X"���U��T�J����kf�{����ePW@����a�ы��	{(-g��/�r �*��uwhxC��ڥ�{Ss#����n�1󝙰NG(Fm�N��8�$��9��_+�<������M�ˌ��T]B#;'d�c��gDnzWɨ�xc��55���9q�l�ɰ����~G�@������2�7�@��B_U�W�s6�1�N��8��mOb�.���{�=(���_w
��V*5� ��=����T���gʲ�r���w�/��$���gm��E:'�������s;�!HǙN9�;��b� 굮s$p������<��:ܞDԱ9����HbN�]���.��{!Q3y<��W3ɋ�j�=��@��U�N��|��=<t��H��sV6�l�܇�i�n���ԗu)˚[��ێ����=��Mu���Z�\�ee쉶��Ԓ�#��;���J�����I�3㽯)<���윙�)Op��k�Tm6V�Xȳ�.a��
�1��,�yof`�^TZY��<�+�.ܒS~�!;��s�W�v����f�.�;��RЍخu�++�i��d�t��J�4	���\@V�����|R����Ҵ��*�_K#�M��TP͓��9g�EOr���-9<y[ޡcy��o�QF�9U=޹K����d���'��f�v%��^�n̊\���ui�F�zgJҭ\�1W4��cQ[��u��G	;�v�ow�SUQUmj7�VE���[����;{Z�GI�k-s	�S6v�F)���~[������>������_#ws��ί�*�yc|�H��4/�P�{�,5�f�tKLuV<0���^�Zy֜[�.��Q���2���3�&���*e����;��N�y���T߷��7}�{LY-K���=*�4���	�R�.��=��t���Mߌ�!٦F���w�����{V�ײ����~�m�{B�B�oϑ˿�)%c��� �eט�z�r�7�a�ȯ{z/|�/�{o�+� ƔǓ�PfR�Vj���+�yܤ���ť�&�B�L\�!z/F����c�����E� 3[�T��T�]�sU�Zɻ�f��H��i,ԥ�c3*ir������Ó�6E�#-k}�76�g!w�N�7p�N�V)��Nh��;���)0j�7��&Ͷs]��;.��zކ�aԪ�U*|�S[�2�y
����C�����zB$��W���N�ZO���z����v�2�MmC���U��:Ah��R/�ϒZFJ{���/��sUg�u��Ի��Q�*���S^xBTr�C����c���ڵ=�w���c0sw�V���<ğ~zrC���'�V�S���'5�R�	36n�,��K��]�\�4|qlP/.�s{�m�ɞ���wm��J����:�Y�ocb��RyX��p�dt��8�1���*�������wf�Q*C�; ��x�m:��w��j&�~<�(�W�%}�`î��Ë�g6tK����S��)t򾀑������s��7���ss��J��}!9�����f"G7�7�kN��������^;x�yN�,s1�#���������������χ;b�>N²e��e��ʂ�k�\j�/t
&P�Z�&9gF�y
K�j�p,��[Oz�L\+�͸����<��er�S����^�o�S�f�����3���9�%rB	p���]�T��+y�K���ӓ�6�������y��7e���ϫoI}<��#&���W9Cر׵�Bu�;�I��e�D���W]޵���c0^�S}~��Bs���!#U���޿_��k{���Ų,�G>�gte9q�dm��S[%NMʯLc�Z�^n�r�Nm�Pձ�����.�ޚEu�����F�C����Ե�`&�}%�^���g���{�f�'P�r��V�ބ��,�ג��ӋQ��A��w]��C��Į�f��z8��Z~{�p�Jj6jD��V�9ZL�K�����h9�G}�����ww����%:N��7���vɆ��X�,�"��~��FAuC�H]�9�P�i�jޜ�;"[��mN�$r�h�җ�ҥ������5נbr7s��tɷ���H�$p�ذې��Vjn�)�,��>��T���eX�m��HkӰ�dk�_����1����@L����<=u��X�奁����@��g�NȬ�tR^�y��b\�tK)�	O���tNj��|7�	���{����(�"M��ۏX��QN\��}걷T��qX]�w��*&�I�H�����{�����뗢�U�v�����W���V��J�`2)��z�{ໍ��wf@�������3��J^�9�������<���	����j\�Y��J���˘t9��9ш�{A�uNs��줝��q������3w�ֱ���s�V)δ�]j)�,����1�
�N��H��Tʫ�~?`G�j?�{��55���n�fS���w%1�9S���[{	�V{�ܨc��F�j[κ���S��B��2�cչ��%��zG�m�{�տQ�[����}5�(��Q�Tk��O�n�<�P�o�s�:.B������'ʀǑ�k#���P.Vm�͙�fN�X��ň�+ujnW<* �21.st��B��Obits�K۞+6U�;�F�C5#5��.C���m���d��E����B�C=}��;�l=مP�V�[�s)ڢ�S3��[�O�,��f�]\��G9����7�򴅲1:=	ֺ�Bш��Czr�XÌi��:�	+�YN��o���1KR��G��ϛ���E�n�h����I�=��-���Dw;JF$��,���.��2��{jZNϯ�M�6t�==�Ϫ�9�\�V㬎�c#5;Μ|��QV�Zv�t�����}]B7�]5Ӫg�9Mp��[y�Z��X�����zq�;}�{>VBU�"�`9&A��̯#���>��'�mE��{w�ރU8���r{�,o:>��;2Z��,�9$ý��,������Q����y;o"�+w0lZ�]K96l���M>{�����k��W5��4+�e�GV�1-�)��=ƺ������Ž���تj:gx̴c�j���v�d	}�+���b�ʍ	�r^y��oa���d�י�?K��S}}��X��w~]�_X*�*׼�8ϔ�]�}�ju3iN����3}�1��c/
�����U:��V��U͝-��g���+۞cy�@����r+�J��)�F�]�燧��`���*�~�p��$n��4�oi�7�̻��_;�y��\��~��)�T�`��x6XY�2"���r ����y��F!��ׯ��><D�T����>�4W���M��C��v)<���v�����1��f���ӒJ�>�]�mI�1����m���:�5�텏�ٞ��^z�r�\fYo3�ykԢ2�r�Ҟ�cl9��n'�J�<Ϳk��=��<êɼ�K�Q}o�فÌG��:�S	V�N�\��S�)u�e��1|wlY;�'��ҜH=k�\���t7�V��_.�S�J�j7W��"�m�@qun�����7�u����}����u鞻�Q/�ႋ+����vTn�d�ƫ�9^mqk~�#�I}8�@~�9\�r5�}Zh�@��Uֶ���E?/3�⡷ϲe�Plm��
o-�|@�gvN��t���s�6�x��m^ř��F/h��f�
�<������D=��7^�؃{疰U��o�P�m՟k-ii<�&F�u+�b[�� X�DBw�~���zRX=��a:6xjnüݞ7�J��
o��
��"�����{5�>1�v��.-�Ş=S��p���ԫu'K��}�k c�e��pm���� �n*�ZR���� w���QG�on�mu�3ct^���`�����ЭO~������Y4�n�t(���޾::>�Ш�X�>�z�w^e��[iͩX���l>�m��=x����c��[�Z��9��gy�B=Ŕ+�	�9#����Dv�4�Cs`F�k�{REy_\�%�7*�W[�c¼�����d��gB7��X�EU�fz����`�tsf#jf�t����ж�����ܖ��+��H-���|�h�pL�7`��Fv�����w���SQ���|wj�^}�z����r���p>|P�U�w�h��A s��/�;A�����aYs�Ѻ{�l�+L�{<0�P�/ν5#ʝv7'����e�}�aJ��ln\3�5���Px�wO�~Y���Ϻ*�ͼ���d_�)g���O�a�3bw{1L>��9���;)���F��عrH��"hU�d�t(��$��d�PN �k4�9�m����-�Wq'~��oX�N��v���y�:8Bp^R����\(�m��_E�al�eh����E��^���ٓ6��g]�n�g���Kl8D�w|UX���|>��5҉�qtϹ$^������vJ�%�z��#f�|�M
T���u�ojH�j�±
���f�en�z�Q��_;Y@侤yӐ��o���+�"��{+K|�h�ݞ�o�:�V�h WLw�: cv�6o!0�ư�F�)[{�e#�.-N.����AX@��/�t;f�Pԭ���݅9��;:�9�h���^з�	��Jk��K��qVk3!ks���w	��:�tq�uQ���վN�w�N�}}���9~�r�%^
9ǉ�3��ď��{�kq/
�\.̔lM�G���f]���G���ˢ]}N���[71��>�0)u�W �\!��hSF	<�E��s uv�8�.A��}�E��`=�Ztc8)��}Y�xZ#x�z�t��x:�zL�0�qL�=�3��k��k§�V5���2;x����òGݸ3�|�r-��S�pz�\}Ӈu�7�%���Ϧ]�1옪�R�CuQ����`'u� �6S�Ý3���N��L8����"�M�Q�]p�ghj�����Np*�9i��vL\�vv�ef}8���n�"���ɘ��
ᑾ�Me"��w�䈥֪#8ʽ���d����<B��Xb���~5���d�]2�Y��;<��ǆ�����ck��j�^Ѧn5F�� ��|�\)��wi��F�˵P��W�S�I���L��4�NK�q�����@�2@t�֥\)v�P睵�q�PRsjM����xz�i���ں8.kT������r[1M�����ٮI�KՓ��HR�N(��,s��-�.C��[G���e��JGN��'���W]<�X(h��a9Ȇ�n.�굎� q ���7���
.�z����̳9a2lS��YU�Mn<���j�����4�����3�.��� vn��]�{uX5�Y��W��t�"�\�^)لa�b����G���>|�2Ehʥ$>��Laf��))f�[��}#,'T 4���VMS׾Mg���,G��5
�pBv�[�U���Uc���x�[��'�����9��2Cv|C��|�#�W��0p��T�M�J\�c,IT�yoip�>x��U��R^�ѕ�m�wCw;ۚ�xqtػ�k��7�Y�GdR#���(�{�pUP<!dUHKH�8�����y��eE<��>���&<2�|x{�s�>�T,�TCrNFR�,��~=�Kl��	#cW)Ƨ�@N�s�a��yb:*��!�
��@�E��{k��:��xD[͆5Z�������+D�9��]<A6x���\t�s�շ�&��	&��s��u�u��EV4���W�=�&�o�TiVէ%�}��+���PK'~ڕ7�Nz;Uv>����܂��q�����Ü�_-Qܫ��K;���;9��O�F�dI�_Q�f|�����ӟ<�Cϧ�I���	ʝ�n�n�L�T��/��2��F��}�G(IW�n��Sж�/�U��-���&��7���#�RξX/����T�w�4�2�+{Vj�W� �Ϸs�- �d�[u������m<T�k)��9u��Xzn
�K28��i�^�R���6�t6m/�3�[Hҳ�b�[����/bH�)֪�"]���g6�Y1h:B�E)�����n�i��
ϫ̨Ă���q]���Y��E���a�:�l����8>���iT(��auZ�[��&�7����^�;�;y����]+Ἄ�w$*b��	�G~�8�	*R��� ��͚�[���@��/r�-���F���1��]�Zc��phh mj�rf��K}`ť��.��sQ����[�__n!{��+�F�E����f����`�,�;J�)��s�Ǐ�p��kwi�cʽ�>��!�UV��I��l9N����λL�׭�*hN�;���6:�J�ř��������,�!ƢJS*������z�t��ψʒv��T8�3 �1*iε�{��	^�nc��S
T-�L�=}m�n��RQ7�D/3L�y��6Ś)�á�8��{�a�X{��,ͷ\�ջu���r�ǷXW���g{JUv ��ztޖi��q]88����5�&�$0cu.`UqI���8!��N�������u�۴򅼘3i�&�r��2җ��۬��pX��(�_v���%�3?�o�8[�d��v���S�C;�)�l�+t�<�"�1U�(�k��n��=���r@�t@O;"�	otةq7�����E.���º`dM1]�W�\��Ij;B�
5-m����� �.���F�����7�p\x9H�4�0���#	��V"�[�*ع��餞U�J�=�=��iPL�ܱ���]�B-�N��.���c����e[y��(&�i��=�p�٩	�h���yԕh�(�[���0�faU����6�up.��L5'lw}8�B��dY�*R�&�v�+5Z��k���z�g{��E��?��AK_���6�+�"5���_:_m=�}�:3�o}�+�9!Ww�q&̈́���;��;���?�4V�0��G���i�΢r�E�W[��S����%��q��������ֻ�v-dL�)���彅[|�[}ϔ�{0_����C~G�y>�Z)l���m-W�hV,p�������-�3t���!Ϝv]p'K��~���۲ɣ�'"�V��[�c�x)�ӂY��D���]0�$��;�nL�����Ό���~ϧ��� *����<a;�2�],�.�6=w��z�=[�p�"�;'7�q�eq��X��N�����sP\.��7�jf>�/�cƹ���"�PZ��nX�\-�$��!�7�Ĳ�;rG�XX��%QZ��\�JU�^.)t�d��<�+��A�	*���YR���ڊF1�6�QEAX����Z�(��UD���S,�̤�Q�KFV��Q�)m��DDJԶZш�)j��Kj�mQA�-��������"�Z��+R���Qm*�Eҥ�)L�+ն�b��ƴT��UDX�U������*�DjRTR�Qh��
*�)Q�X��65�b*���Af2�-j�-�)D�ZYV�QE�B���V6������X�Fj,-(�Dc-�Ԫ�*,Hڥej��V#R�j�m��J�UkTTkV2�Z1��ZR���,��UZ6�j����Z�X�ZXU��J֢E*Q��ŬU�ja�QX�F�J��#h�1m%+օb���PADX2�1�G�Q���eq�6�����h�&fdKIX�E�UTQZ65�R�[�������QG,��r�*"1e�E-*�R���aU)V�6�j5
""�F�F��DV(��J#J��>�ߍ}u�׮.;�nGS����ݼ�k��i�F�i\��9ͣ}}zv�&��k&���}�#w.��q^����7�Ic�����}��έW�[�A���xq�����)��e�P��c<=���|���d�*{�d���Q���T=����(VO�����(WY�w��O����|�<���;K��I���	���}t��$��fz���3�Ԉb�Ϭ�|�"�������W��y��;���O��t c�Ιc�v�ɡ-/pw�ע�������X��Fs<\��Nv�/rS�c��m�A�r��2U3N3��i��n�0Bpe�����	Dwܫ��2_�����񞣽9��/|�*�}g=Ԭ�nk:h��k�=-�=�y_���ơ�5r^�S��C��н�D����a���������a�W�=S@kU�+�|�R���s�-��.�xφ�0�}�tc�RV��M��� o:ƅ+;η��/�_oBN<��G��*>�����k޾�ڴ�,�H?+�r�y���em��p��޺Ɗ5,=�������Txa��"���t]�����T��'�*�ʣ�j��BS��6;����ޣ##t(~0�2/rB���y�V�/
��΍ۧ`��&8h^����%BĮ�V�u��g�V�b�������(N�z�h��wn3��;2�+Se�ܴ2�wir�-?���o)����<0�6�5( �Ou.���\�Q͕��A;�/�f۱f�9��7a�\����eJ�
8�ɉ�d��e��2�;��^��">��]�0"6�L��}��gd���ŀ�c"�����ْ'�̒�X�;��Y�s���SI���}� �F�q�2��޸*��u7^ҋ؃n�X�YωKV]�$����i57w{P�!�F��� Aω܊�r��0��'~�@��'A���.@�w�juv5Uo#�:t�b����#���hQ�����N2�	 2Ngw�M�r����d�܂��g҉�GS�Ny�����;�G6`b6��e�{���c�f���������G�¬g �y���; T`���F���~h�V/��2�ܻÊR ^*0�l��3f��1qY��i]&B�tL8�/g���ȏ��)'�����%Mt��*F哕�+~�>W�n��ᄯ|j���H���q_���-��o��]l�����(�h��܇n��Q����	�Uj�&>����dv��?��kT\Us�u�[����]�ݩ΅�#�Q�M�<{r
B���7�l&
w���H���;v/��y����
�qo�9��T��v�wx�L�V4y��ͩ0)[>�ze
�o�n�w'%5Z�n���jŕ�,F�S���.:�׭؁׼��1yHvb��n�m�SΘw�����w�%9Bf6]M��)�g`�0Y=�׾فO�<��6>_K�Q��܄Uqʅp+m_Xxӥ�9ƋǴJP��U���u-�P���q�eu��g_��]��Yܽ�UZ���ǽ�-����9�<`���3d>R&T�p��u���\�Bک0�B�(����qk��dN.+�^��<Q~��>�03��/��ٲ�ڕ���݋9dW�_XYUq�pw�^="�Sń�1Y}�_lYnf4h�x�����^�F��P�q�C�ogA.�e�|>3\nÞg�h���'�XZD��X"����*����E	�#���#�G21��t�ER�;�i\tX�:�WhE�#�Na���JJV��A������U.*�?�?uv�����v�!HW^�pv!����c8)��}�g��7��^�w��W��M�]�3�n[�`�3b�x�c&z(GJp"�r,�!7�ET��}٢?�5~EZ=��o�?,�XV�[�:~�C{f���|�)l���A�0�v����S�Ǚ�5"�E#r��i�f��<4(��	XBک��L�Зۨ�=����N�V�[��luj@�(^X���[�R���ojl�M��#\�;�F��G9��`�Vµ}E]7�������z�	aέ�:�	Į�Ƞ��l�9��B�/��iv�8C&�-�"�*l�>��G�pc�ȥ���5 趹�5�x����u�H��Ǩ��^�Fj�&+�Yp�z
߸�q�o�����H��_In���t�3�{���N�r*�s�v�2}	�f��I�h4}�+�ʩf��0+67ƍ������Edl2�����Ȕ�V�&:6�����ְWk��'s�����B�bp��0&u͸ne�8���S��[C2�ް��ÿ1�M�Sj�VRƫ##j��*���ۍ"�T�Y�S�7�Mޑ�6w����~�P礞�^�L�o\�7��߾r!�C먐�N��i����:�^����GP:�Ua�WZ|��Y9������^D锼��O��pJ%��>��8���Ϲ���j��}���EQ�1k��|uM.:��^�~�n8�A㫗PӼ�e"����2���ab��RF�P��3��M햤nl���+>C_q7�j86<s`4͆]�sf=�Ǘ���1#
i p˅��fDM��J�As郾<�sT=|�vKKd`�]i[����7:\jq�(��������9�fY���l���E}x��w����]�Բ-j����ȏ+�Qi�Gh:�P�GdR6%Q*�wX&��*�R�S}�Ts��3�]�̞�xV:�{�ݨ�� \xa��3�Ā�U�s��`BqH�oFT�����&�C�)5�����8G��ML9����f�J�
�qx��t��w������w�$`SO��\B!�>ע�cC:�C��,��&z���s��Wэ��m������$�t�y�z5��D!dY�^��r��q��g���x���Q]���ݻ;���a/��s:�A���F���5X��$��Y�͔v�n� V!��=yֽ7P0�ꛬ
�⾏}N�����)Ek��5|k�lt%Q8S[�{�䛰��+�ę�ǃ�Ԏ�\x gG��>��Gk=��Bd�\�h���TZ���11�ض��N)������k����6"8�׃�	�!ݕ�Ę�q;Ɇ�d�m?	�Q�>�Öj����,}(?�zr^�8x_��ja��lq�8���'~2��_%q��t�ƾ:�9����,{�Ǹ��Ц.ߕx\G}\�����.F�����#n��o\��sj�w[��K�<� `����}�z��3�r���
\7s=���gY��W/'�wMv�e���o{0CS�-�t,%��9nkx3�ebsD���vonD��O;M��ħ�-c��Vom�Z���$qطH�
w#�s���0�oNu�uq��W�$��s�L�a��,�������|}���u�� �Ճ�����W$ *hؽ�n�w����]s��#�:Y�Lp�4��}s��]a����cl��'g;Ďk��+�>���+GF��81���έ�k�\(\�<�'#��<���'KFrK:`�ﲶ��f�P��U���p>�`:�twM@�'��	�v�khQ�l��ƔXĔ�K�ҡF��N7s��>������;*TXQ�
�.�%d7���Wn̺��}&k��z���冋JP��%=�x���-��E.}�jeb�6	e�=�������~��X�%�t����b :�Dr�q���t�W�Jۇ�=��w0zx����R:�u�v\���J~������)Wl-����>��wa_�t�=Z/[��g#���{��:�]�~�=K���OK������QϨ缙�Gg4)�딄0�e�i�d��r�49�BT�ʛ&t�Ӻ&�T(�.l�Y͘�3�v%��4���"�;���CrW�:�{��O�q(����{�7��kMsg�=��*�O�"%��\n���H뷯��V7�9��W]r�tzH�.G\90C"L�:%5
 +���U�i��4\�����Mʶ�R�{{<S<�轊cdag!�d,�DÁ������>5pN��Ds9r��Ns�z?wn�ո|W�xD��7��bmָ0��R1T�O*����ȃ�dh�q�m�X6r��Ԧ��Z�K�7�J�XR��iUF�;t��X�G�a���k�rc���M�g����dw��v���������ziC�e���$��&�WU�;=n���)'�2U�;�������ٗo�NK���RE8�����Z:6��8s�?��\(������Ƹ]�����Ҽ	w1"8/�p�ޢk��"���,�i��jx���X}jš��}kRxt�N̬�7g��xŔ�𚌮��٣��+a�9۴�H���H�lr{RGj��s8��;(����| ܪI��-?���+��͕�S7���ŀ��+Я�"khA��z���%��g6�2�n�������XI+�g������:G����K]C�?��1�od�k���'�:4�K��9hK��E�G�|���c�r�PQ�}�k�.bZ�.���f)�Wr��r�v��9d'��`Z��T�������[Z��oU>O)�N\�B'�Ŭ�8�i/�'�`鉢ڃ�t��t��9��ퟱ��ǋ^���CU��B]vU�&{(�u���^���mt J���:P*�6+{�9�>i<�Y��a���=ǧ]<z�@�>�;B.�PN\����JlF�V#�f�����gAZ=SR{�M28��6��Ɨ�֛Z*|:}]<F	s̆2����#��Z#x�z���8R���.m�HUv��NP�!�;��v2g���h�E^ .���4�'(��m��<;z���w�&��G~�'�B7���Y��6I
v]t؎�
q��8I#1�w�g�VlJ��9F?A�x�!G8�!���Msپ�F1��吿V�1וTݲ%���3ۗs; ��+����PB�����Rb�>&̳)���V'Ua��%#��C�4�\Fp4\��;g< |l�ƻ��N�a��F��f�Uvkn�
͎��^gҟEij���%瞬P��6%jW�|�z����D�C������%���%�i
E/U����8��X�Wq��,����G@��d>��nY��~B��hfZ�p��S�6Y���P�ǭ��Әs�nÍ`SvI�\�י�R����tή��r���]�BPFH�*�`�>>��.�{���b�r�َ�$8��Ά���y�|�����xn�*�NL�P_J'��u�x�Ij��.�9�.κ�N�|�|!��,�r���隚]���	�Ά��u��z���.�?�8�t}�}��Rg<�D�:�XF�S��2����ܽXX�ֈ\���t}�����-��˳�r�o�].yr'��r�4<�E�@Ns>�4��;���87Z�P�>���ǟ�֫;fwK�8�Y�
kҥ�<�e��I��rebй������D�ݾ�r]W8g#�)��Gz�U��Mz2��R�J�T^�T��5Ȥg��������O�j:`��E���O(�W�$�gܣ���؃o��.;�fk�^�wyK��X��Y���T����z�}�OM� \P�uwmY�N|樤��RfXc �0�_k���޿qv�yG��Ӣ���㋄:�E����{g{*ܭ�wpV���i��@v�����~T+/�@���n�Y��z�^eKy3�Q�p����~�=Spծ�[5p�깲42P��}�����v̡]g���gƳEr=<:��g7[���Oo�n�n�D��h�i|�:�3SX�V=@��-��g)�n�s�xyw�]�]�~�};�e��D���k���wp%�4ej�O3��m ���'�����ֽ��\.{z��>uxv��k��C���d����'�U�g�  �~}���6z6w���d�tin(Q��y-[�;| �����+�����z�#Ǆ ѡ�z��_v�~���,x<���U�E�i���pǺ�pI&=�Uh6�i��n��������K=B3�>��a�83�R@^����� 0a��y�y���Â���Y�
���5��ަ8Ay<�V���!װu�w|����!�b=d�����¬��^�9����D�J�f{9�ś=e�����k
�	��P�J���2����3��ve}blVP����}��X&�A�<��0^�f�)�>��4}����}+د�L��tK�Dpt8A�|9԰v�t�W\�����el/�$�fZS2���+ot����y��kqs��=>\�o@�����1���SoJ�r��N���3;R��Q��fh�a�\����c\gre���V;SL׽��s@�Z�P��uڮ���u[�t��$=�{1�I۰�z-)���He��?'����V3 }�[�죵�Gm0p(�Ԛ�/3�R%oy2�z��N�9X'���9����,.�v���'K�'��Idd��7X���b=�cM��s���n_t֚�C�v�3WK����kas@u�}|�Y��V��Y�;;]qm����S1�˪"����
w�*k�e��W.��g$N*[x�Vڼ�2��tit����K�V.Ȗ�KFu9fj}N���j��e�sOL���#{�<�{X9[�A�*��15R��y@�2�����b�X���R�H�]w=��yWM̺��f��e��ﰕ�b�#�_�\�
@�|��y���@'f�<-�q��T!m���\��eoR��Ee([�t	��3�u���Sw����x�V�vt;�u�ɠ�to2d �_mb�dKg�%`��7����Q�����\�V�f����m�'h��S��Ւ��np�:��<L��p`��H*�����U7���w:�C�x�X��
R�LCb�f�1[�9̙�n�r�}|�n��+-����k�]t���'0�V�f_`\]%�2�F;�Ã�h�!��g��¸�y���4¸��a��|p�M9ԭ${�"����+���po$ �sV|��͘k�Fj1��ٟ
7�3�C��>c���NwO��[�cn�u]ɺ$�{�ۼ;�.0�`u�b�ik�!���c�[���f��`?�<Uv����N9L]C��QW����������yWw�huBjtt��Y�h����l�;y��Qn�8�F����P��xcັ77ȁ8s�2s=�B
�$f���B��u�VL�`����?�B���a;s��iVʘ���WH�����.}*Y^�^Ϛ�Bs�oc]�PWs��-8�5`��7�}]E|�S�EHs��:��F���G�sa��PDٙQ���I�,��#a�UwU�Ư��I/9��I�7���b�+�o�ק�\tM�<A<�1s�r����H��}3C�(�5��9�a�"��e���T�XCn�U8���0���y�MEZc����� p���hH�7�	���x�H�����a���-�Q�������}�
�Jj�J�ax��,^C���$�h@�R uNe)Ua�s�������W���!�4��F��gY�|�<m~����v4$�i�5�EAC7�>x#��9�5(%4!mk/KK�$�V�nX)[�rH�Ò���-V6��O^qa��o�a�dqOt�Σ��ٝí萵eٌr��1�ԓm*���z&-H֏=����S(`��C��𘯃�S{n<냘�`'�:��
hu&zH��iX�Op[!5����C��+U�	�����[�y����=|�8�
1-�e�£J6��EQcZ5��
����eAml-([JT�QkV�Z���3%ULe�AE�l�,bʈ5�ƴUKkb"�h��F8�q��!h��-�j�V[T�� ��+J��eZ���AJ�,m*�F�ڪA-�)B�R"��-�Z�Eb��U�&[��[H**�Q�k�T�D+��6�X���1Dƨ�b�V�Eb��J6��6�EUh�DTEeeF!�LK%j,Z�QEDQ�(�1�QV,e�A9��������"
�1T*UQ!mUUQPUX8�A2�ii(Z�X)mTAB��%aEVT�X�[jڡZ�[b"��"�mUUR���m�F#mQQ-*1�j�c
�V�Q��l
����f`�[�Rը��-
+AJ�e��nZ*$Xe�m-��Qee�YQk�D�����U�-U�+X�մ���+[DV*���(����l��*ZH?�Þ��b��kY݄[�ʗ6�]ҭQF��ͷ>��ˠ����2�:�9��(����Pd�Qh��|�����n(����5�+��H�%j%v?aauD����iq��;�Yk���qV%+n�=���;5�5��Tt��k[SN�="=g��3���d� �0{b�!�� sjkh�+t��SZ�K:�њ�l�F�� ��
��*�o�zߢ�GT]�)�ιHB{����+^]�,T�*�C��
"��dҋg���ꗀ�TqQ�2���j:�a�ܾB{(�t� �w!�rbΑ�fӭ�Y�� �v0:q^ T�@�h�O�3;�JgL^���{�J.n3��Ʃ�ث>�FG]F������#��;�~�"�o���yڒ�����"��u!�QX�}I[��|�M�pa)�?e��>U�v7Ng��\�e�Ɔ;�4��nD/ۙVl�bdI�OD�fJ��D]����/S���*���J��㤫*�WTژ��s��Gv�;Z�ؕ�܍]dV5z禔0X��](��;�RuO�٭��t���rۚWU�92x�%�\��z�j�<�����!�x�8r/?��\(����v���z�7632M��C�7Lf'�=�oby�Uꏮ�Gc=�ouV�����<{+�7϶�����c]����f*>�+�<��{�U�0l�ེ\�BB���W*H��e�N[e�L��G�h�G����^�%C����uI�����z5lg�८*U[���������._7S&��X&v5�}z�K�X�Ui�lU�7�+5q<�G������b>�2W)�d3%�>R&�ۋ8�}#�6\D�.�rӕ�v�/��j䘁����{O��V�}��`�wbۖC(=]8�����1�$�k�� �kO����������b�}<S�5C�ogA,T��pd���J��QCkcN�e�j{l��*E,"R��`��wQ5�*���Qu#���ɰ��S�n���eT"�Y���N�����s��0)O�8�'��ޱ�/�7BfT]"�eq���m@Z�`+��2(�c������X�g��=�"7��f'�[����c"Y�9�<��4;�[��L������ʌ8� 8IM�Q����3F��M�0|o�#��b��Ħ������X@�X��㫨t7Q�����r��8����֔eQ�=�u��x��4k������3�6#��DT�ǱȔ4Z+�.k����ˡT��H��Q��i�)��|��W�}&�D���� \�*�w)vj$V���v�*�a����B���d�M���]�o�i�@�^�+�s�d����en�C�:�7��70�_5�6�)�]]��^�1�q����߬<Pҹ�|���65aI��'"�$��F�uV�E��S�ʊ�����u�H�,MH��kQ�ѱ��O��ـ�%��>��K(Գ\ 8J�i���̧��P�Q��T"�g^��C�3��)��d��"63e�*�����oE���׌]jS��u7Y>�mo�l h@;C��.(�ޖ}��e�3/G|�a�"]k�Gx������5��]ѱ��N������J,;��'*�H���e���F-M���(I���x}�>�.%>�+KGmD��C >��lf�7p�K48S���ڎ�2��Ur�����Ȟ;K��|��3�箪���^��v;#T[u���l�UFx��ݺEºDi��\UB��R%u�~��D��({���dS�ųj���N�<d��n���D�ݢQ�=L�z�Q}�
�U�u�L��	�u,H�Y�[�Q�X:tЛ3�i�+��<���GL���.<3�,�mi�Q��\�ʻɝ&,r��������9�b���!u����R4Glm�wX�G�6��4f���h]�s0Y�or�ɫ��G��H ��%��
)`ȧr��9��__�╎;k{DظM����k)�s�H��_p\��w�^���Φd���W�i��B�K��a�κ��u�K��an%]�Jr�V'��]=���z�nPU�Onj�vΕl={�z{G�pQ�/�*N����C��@����z�X�f:�k�{��v}맦���A'uC��9?Yه��)��Z"�= F*�
=���xG]��)б�\!Ԙ�ʥ��K���ID�h,g-�6�	&�H%tc��3�A�UE�CT��4J9C��0���v��r_hw0�+P�zΚ��~��_���)��9�'gpod
�`�X!�"�����B�g/sM�(��&��j�u��,�S>��؂ݺ�:��R��pTFĳA������x�n�k{���ݽYԏU�(_����zX��#� ?�y��ʷ��4��wF=gFKK̾�{W���ޱbSR���c�������2���!;�,����t,���c(\V��3Jj+ �ib6If�s�h�l�BB�*6�m �,�`v��;s�$�ˆX�.jZ�뺵
��o*׾Yf���Yk|�=��T�vz���a�������� cF�%�v�{R�����ߺ���7cz(Qb��dX�J�߫(QF�L��E���u�(�Q6�9M�34�Z�g��$����}w����e6�����as�_���g�=_��|�(�3h�R�,�!oZZs��鉞!����I�R�+��Go����R �^(�U�,��/�.��θJ�N4�,w����E�L���cB�����)����s�8.�G�Cj6!P��K�If%Ҧ��b<4K�}{v���{�=MfEa �k�),s�8̰���
�3�;*Tep�Η�A����)s�P���}ڷ�X�[�t��S�b6d�{�=.T�}g�����kB`��&�N��/�r�^�&��t+x��V�O��L��=6�y�z^������8{�Wޓ�9�Mq�`�\4��q8 �6�Q��q�hT�>+��0[YƜ�9v������~�î,D3�a:|�势+�LЕ�g�R�l�10�J��JAf��dКJ͵&�W.e*��AP-����ʙs��Γb�'faB�6S�&�z�U���f���Ӣ���S0Z,�!P�E��
��&{��3d�,\#��0&��S��ۏ��]�� B�^M7-3��k�
��ŪC�6m�U�0���GƼ9�|d���k#��OƠw����ן;���t�{#���a@B�[x�r��LYu�pv�V�L����[��6��
y?w3�u��K��
l�Fa�%�n��ɾ��.���egu�[�w,'��11S�u}/i�7�������bfv L7�����WM��n�5�ڹ�Z�d��6ݥ��
>�^Ӆc���aq�ٺ��S�Tr��K'ܪJ�O)<�cx�Q�][-�z�,)R@4�3=R�v+�L?��������:��Z�e�ڙ�9#���	Uq�F^GcW��D��ч�Ŋ4;1Rn7���R a%ӝ��Y�{��
ɾj������C!��0����+GF�6�(��9p�xn�z�`�N7��{�ˬ��>�%lmGDw\��T�"�P�����'��l��2���R�7��o\�B�n�ج|��j{�G9?&�Ҹ���3yV��*���{G��`^@vL�'��-�+پhPp��& i*�N����Gi��v;��z�A�f�c	��{��j��!���{R�ӗ0 Є��af�bQ=m}�.�;(�@H�=}[�맔>	�eK�vH-� ��o�?Vt�쑩�2/d���J,2�#��tmt G��!H��^�Ѿ��xw,M�3�c>gGΤQ�w-��#zQ�J��v;�g���0�����T�C\ʦ�9�2"Ň�kݛ��D���_�����<=����d���=���u|���LL����G��ވ�}uGi7�w��݅�:;$e5���@�$(���}u��g���\ՎL]���l�ՖՕs��� .Qˑ�JI�`���+.CW�Un�Q�����;ёyRܲǾ���P}�y�s̨vZQ�whր{2��8�^�-mUҮ�c��m�����e�:Nlec��έ����]�5w�PX�>�@^��yq��`yOi�?E�
�>Z�������Pf&k��f��{��t,S v�̌<�W�F�o�`�K�f_,w���UPF�P�d���rd#���s�&��':_�ӻ����B���9>�
LW�6e�T�Y��W�EEI���_qk�W'l8[64�+�j�"B�s�b�<1(�L�NCs�'}�َ�p�MP]��z,��s|��G���Ck �8`�}Vs꫞�	w�j��Z3ԣ�|���_�Z`&�=�4<�GE��s�[|�6��Su���A5�� �B�y�8]d^}<Х�bVO�s�������a��D%;��T�Y�"WO���@�J,�)�Ξ�\I�W��g%6���!5�s�c�;UE9��ȏV��Q!��C^�ҫ���h�M�AԶP��'�榚ƕ������e���x��g��I[��@@J��'YW�5Wu��
�eo`A�u�*��
�9�O��v��Fa��E�r�R�Y�G#�5U��v����ꭊ�
���	��o��*e��s0�5+��{I]_dv�����;S�g���.���{ʎ�ˑ<e|�_���)%��S3�;��t).neutv�+c%�b�,_Vla{#8T��+-g�"�j���]t
��d�	f�[0v�ʺT����x��P�?tΖt�}դ^p�wq��_��2{bQ�p��P�(�oGvSU ��r���j7�l)�ʠ]N�56d%�
!H�[�k�:��`X~/��ΎWJ��9yx��ac�xA�����`:��{��V+A�Uγ+�ovz���c(�|�"��'������yp��ιܽ"	=p�2KQ~8����7�x����fQ���dV-$rǤ>y����SО鞥��Р�P����[����ӏ�����4l@`�	۝6v-�e��/�j��!ϓ�U6My7��� �a�1F��đB]�T-�X����\5_[C�(O�t[������ q?g}���T�<���Ek�h��O��C�t�_%���z��MWB�K4���t��ζU��d�֗�ʃ�O���6��� �z�����p�gNiC+���mҡK�5m��Fcn��-�}��f͂��8c���6i�]�~՜8���{W1L�^WebH}nv�o��v�5��Z����oPlzZ�SD���qb�WOd��w�kKMΜX"�;��y���wn�{��K,�N��h��2q5�2f�����f5�	��yn\���Ik��>�8�BV��!7n��/�ۜ�� c��Dʐ{�9�}jz�F�Dq�y_Lٶmߺ��y
7�D�<v�m:!׊���tg���o<�kNY��vT�k�X�����cL�{:X�O��ѱ��!lX�8k�J|��#K<z_7y��>��[dH��<��B�2�YG4u�oؤAD#Eat�`��*� -.g�l� ﬋�5t*Ħ����ѹʘzsM�Sܗ�;T�����S�@�;� /n�l2Z4����U۵x==�D�Y��(�ĨY�ޤ�.��&Z���uA�Ź��n�Μ����Lrt#�O�����>��w)U<�S�պo�ďN|�њo*����aΜ�,l{+�v:Ct� !`=l�kY�+F(��ء����&%1?}��u�n�;ኽ���Q��m'4��"C5g��N;��:�^�`��������Li����ü��{	J�u'әy�l�S���kmi�|���y�>�lZ��*��J�&gu8��,r���k$*���L�G�&����=���Zɣ�W33n.�`9�}v�ow.X�%��fV������wVtG��)A���8������Y����=�u�})�m�T&��yC�#L(S?|<����|�BB��Ib#�2�	*B"�m���y�!�w$�*����x�]~Y��<wo�8Bx�d���t]E�����t4HW��N�tJy�5����mm[v_9���S�jccg�c����G��{��+<<�Xu�J>,~�W�wK;V	H�~��=b}�X�xdą|ji_�Pz���6��)�lוC���3ܡk����N��͎*���}�Lp{�pO��
T�x�z$Cݰ�kX*���`P�OB�<��R��jUb1�*h�v2㍌UI^y��+��:�"3�w�
y��r� t�$������|�;w���c��@^{ �l :�^����M3ŋڸ��� ��o�������|�xx��FY_��#��_E��X!Y��D���n�o8*�gcZL�>��1#��y[{C��m���U�a@��ja#8�7�֖9⁇�o*K�t7_*�WnPa�*^,�i��%�z�<�7���c�f���X���v�R)�М��:�u���ri�L�@��8�4��gĮQ��Z��g�r��}�[���30?�!�o'(�C*�bb���+Ab�]c����1H����)�^�;#�Qַ�����Sl�+
i�c�
������[L)$Y]��˭�ڈkӠ���I�o6���
Z�PM�'�풟uc�)NS�2�2���e��Sʼ4��R��3sH��g�{:)���{)�5�����v)�x����V�7o�*81�yw���,r���ƏU����2\���HP2�7��5j��s�,CJ��	�Xo{tTƸ��+�%��wTj�v���Z��/�lԖ�
�F�cT�rf��K�mb�y�#WR�m�+����km�J��/�M֍��E0(a� 7i�d\�M*��]�.�n`��geM%�J�i��.��D�+��/�D��Ko��,��\�`(�D3w,��m���g��y��`.L������un@�m���e%Kq��-���\�����h|��[�3����80�^V�Vyv�����/8�q����\�!��Y�w@�VB.�ǫ
(�|e_�S���e��}|���6˹Ԫ�=�*.���W���g���Sw� �Nmn���.X�WN��p茌p�'�ً���|4;wq_e�kl��1я����I�3�+�
X����fp����iӹV萌k:�yWv�
�,rul��i(�|�S������R�;� �jnf�(�iօ��\�u�4Ku<Y�tN/ ޮ��S$��O�Fq�S�����[H$	NU�(i�T]]�<��� .R��nn ;fgItS��E��G5n��< 7��b��t0����WFmǜ"Z��L�wegS0Ǒw�IZr]j�섹JuA�E�-�ڇ6�`�k��\���<��Pb�7*�n-<�`r�4�^QcCb��g�,�,�&cԍק���J<oF��t�
���S<�g��쌇I�`�z��Fz�dMh��Y�	��D9'��M(6I"�y�C[&�K.���)l�ԱUƂ��q�P$5%!�!��t$�8c6G
�C��m���t����6�8��ˬ����-���[��x�Փ��RDI�Y���׬<��6����47�Z�6PFM��u��'.I>�˶�tӜ���)WLO�׍T��%KH��ST��j��L��\�NAB��v  (�>�A�َ8+"�,��"�h�$P�������R�h�"��QF"+�b-�APQU�1& ��ek-,�Q�5�Z��
���AQR*�������Qh�X�ibԨ6�TJ�[*�)J���-���EX��Q���Lb�Z�H�T�DX,X
��
���[J%�[A���UAUUbţR�T�U��ʔk(��#����VZ,Z�"Q�X��#R��V�b�������Q`��H�����EU�
��Z����P���-[Q��Qc�JƖ+҅�����-j��R�Y��*�-��6�D�-�DU�L�#TQEAU���Ebe�Uh#�Tj-�Dj
��m�6�AUD�ʔUAR�d�-J±QQb��1QB�m*�kE�E"���R����E++"��LKDU
�5E\�����mZV�Z��1U��U�IQZYQ�T�TR�icU1AJ�F1Q�U�Z��1�ƥ�@�
(W��i�g�̠[���<����[�<�C����mc0�Ӎ7��gz1
ru���:�b�Sp�_r� �ׇAsE���7�B�y\v_;�v��Y�]��h�O��:5Aõ& $�����F�`��~ܬ*Ҧm��q�^�*�}��)�鲺��\gyy!��E�,B��D����]��Q.��������.�s��%�vF�d����ۖ����qq.�C" x�$P�:Dp|��:���eB�#fl͑Ƕ�.4�s<F3�t|��Di�u�]��q��8dq�}5,���`�3;�FP$J��PVА�;���2Z�,ePh�����~�ny�sj�Sx~�X^�kz��kE��W�O+oO�
���ȢM^èq�˭��Q�/P�-�r����ی�QC��B?�+�����<&G�>ʊ!l9�k�r�����S�ά��Gx�z��ʍ]x��	��Ȃ���u��*Qe�=W�~��2��+�+;+���}�������F8� a�=}E�Ğ^��|���y�>P��zQ6e��=g»��J;��X��]cѯ��v`���U����l���ճ|���&c��52��zݡYL��s2�/�l��lv�*���^��P��D��F�ʃ���-�����g>�zD��_]��ӘiP��l7v�v f�s�Q��Z��q��(�tYb��]�r�-;w����{\x+]2�s��V����\�n�登9��q�Nͣ����g�9k�jJ�VlHhـmjp����������g��[!��Y[u�>�����/�q
�K��
���0q��@�D��Gp�Q0h~��=򫴀"���{��Яn�C�<��>>ވGm��j�ŔN)� ��r�k�c�7[1��v7�ժ��U^��at�z���rv�,�]>�G�a먐���i�X����a� ��h��?^Od�!���_�xJz�>��\��+�P��%$��<<���vWq�מǓ8g������lt�a�Y퍿Z�]��D_�(���)��� �
FQ��jv�r/<�̮��DCԳ%��1�YFMwF���A�w��0�L�Fϒ�J�Kqʦ���1%��{�G.�q<㝂k�1]�0�:.�%�v,���tW��l3+�a׋��fF�cݾ�2Ml����>N�Bh��N�7d-!�RR�!_C�I�m�{��s�H�����ق��q�d�1�-G�ъ����
�__��t+��;�7�Lf1g�fS��_����Ɛ���ͭG'�P�s�J�X8���2l�ʋI�x���A+��3Nn<l��}q�����]��>�Rf�k�t(���
�ws9�M �)�$�.VȲ����ư�Z���SěӦ�X�Q�YxY�*�3�.Wj�l� ���ǀdS~Ȗ��B��W��qHM��a��IS�2qZ^����^�7:��aq�n$�x��nv�t�L�~8v:k�nP4��%�H�s� ��P��v'(A�*�E�g�	�S�Y��o��R�xm����g�sP\���3n���&M05P�đ�g���6�UW�w�@���Gdi���$�7툲����b�3U����3Խۣݚ��$
4_8��� �u���6k�UDj��*�UЪ�,pu�]W 1��=�o堸�fۊ�OW�G��_�X\Z�J�������S��X�xB�u��ҫ��n
�ķbz�ٽS��̸�\��bQ�Q�j������d��)��譜�U<s1p���t�[W8dj�m)f�tV�a����k��N�_�e��A��zO#�YD�n�k��\����ڮ��D���:�p�u��Q��"�.{ �T'EeQ仯f��\����Y�(�+s��l���I��=�])�]�e[�(�u�lb�!)�1.��̰�^�����_
�܁�������~ʒ�o*a�͵KN��\�N��8�:� �t1�U��,l�
��u��;]���<��kG��Q;�W�[OE�YнL1\��N7� �u_7vУFض�ƂY���	��T���T�T�J;"J,��Z1+lf�'	p�,�R�)�Cw����{8Z�Wv��>�rcπ)k�_P�X��>��
Jqő#���!���ci�^�VT\�3!��1�^N݇���"��$�9/"�� ��O�[�<nk3c��n���}�ۦձ�Xޤ�y�KV@,OWy����[��gB�5�v
U������I'!ы7v��J� >Gg�+b�4�"Ȏ��>v��XWT�A�a��Dp��	���8^va��N��B��t��w���T�J��m=>��. �3��$�	\˰����:��9;l4t�acv�`c��Z6 ����\PFB;�EpJt�J<������6����{�ߘ$J������p,~�x6�����?xXVxMAWh&���8UG�h$��@�?{�F��h����ؐ�>5�(���RX�|��t�V�U>�~�q{���ZM��gl���+~�3|�ŀ���=�LeA�B�L�^�g�릠vR��3��A��x�Պ��7��7f��\ �<��u��� \9N�[���e�_;\e�z�T�%�<̾�:J�n1�U�Y���YÔj��ue��g��g�r�KS��8i������n;-��d���l�B�wV���2���Fm��}ԤggdhK�Z�����Ov+���<G�r\����j�G`�[��� S��G��¶+}L9����^]E��!G�У�	����t�i@��){�>�9i}ì0�m���S�Xg[�zt�¤�e_{��� ׍�H�1��*����>�Z(�n�N�b�[�4VQɅ����'��VԖ�D�9@�4���\���N��_�P�U�i�ʗ�̼2����˥\���j��F^P�
O�����<�>:�& $��#��R���|���^8�-�G����߄9�I� �u;&T/'.`A)I+};��(.�C������R�`]o�W����:;#M�/����C��}��C���"�JE���`��v�%��؂}$�|�����PK�d��lUaF��/'x{D���h�x|�<i�,!�/S)U�����\�ݦ�E��~�VL�%�U]3]�5�T��N���]�Fzסb�s�?90Z-�n�}��p}��G���7$a���Y�<�Zr�HDN���NUtX���DK�}ȎP,z핻��{��Mr=ǘ�fm7�=U���׌�oQR%YP%,�XG���Yi��66Y�ju�6V:. ��U�E�V��xϳ9���E�sr��\�x��v��A�����l���7�U.�B3cN�:m��]F��cb��ͤ�ηJ\��\����i�N����:�`� ���	�ˣb���_�S��~�X��*܇V�\"�c���Fւ�c��h8I�wN��U���_C��|2Ϫ�`�Fy}��G�J�V�*���K���=}G�m�<�1��^  Pj�bn�q��ލo��*in���S*�ufC8",������1Zl��)��q�Q�3]X=�vaS֟�p:��e+ʆ��χq�g������8�g7�����	},�=~M�Si<˩�kg�c[>6S}'�\*�,�{^��B$�g;�"�K���%��!S\ѶX��4+�$.�|���=����p�qE�.wU��)���^�ܞ�ϋ��|��{��'��9�u��運���l=uQ!��5�=�U��>ݎ��d�ޮ��D���z����tr�=OUy�tp��.D�<g�>n	_$���K�0Z;o4�|xǱ�m�Ҕ�͜+cn�"�VZ"�(����K�P�ڑޓ��ӎ�1k��Vlh�uj�x[%�Ԩ_���s�	@=S����&��u,ЬU�+Լaê�]�1E��Z�������l
�r�B��o�啵aC����e�۸_u]��t�9"��u�0��u.2��g�\����u��&��;�<��H�ޯ�� T�o����)��2c�jVsWeu�����V�g^C*�&x�Y=)%�&��7��h;�}�	b1݃*C:Ԅ�.Ő��x�h�0:����WMb�n�fhͽ����ȵ�}��c��׵�����y)w��q�'v����9eGrk�)FL>ޜw|�j�vO{�Q��>�8���Pf|����V���D"�I��80�����SSݮ���"�5�g��-�����'HQP����NP� �QdA⒡f�L�4�vnJ\lTW\Q�l.!ҝ�F�
|�XU6M��7઱ԃau\��B`j}u;ȼv��]�)�BHbv�*,��F��'�؋.��
��?� 6�f�0���+�ud3���:�<Χ��@k@�b���^������S��x�%j�q@(d�t���ܦ�P���G=n̯uxgP�C81�ج�`����M�P#!���
}<�`��)%꒯�=������b���1�L��X�O3�	
��)��6�SK�}'���l�z�Q7��]����(�'W����{w�>�^�h��w)fK���C/��]�_������
V�9��
�om�ޭ���J�B+��-e�_z��L,5�+��L�*�rV�X{<+��U�~ߺ%������y��6���j�>��q1��V-R�x>���&ㇵ���vz����i�'MS|�q��$*$s�d��M{��36!�o�֑~׵=�㈮��
�C&�B����$� ��Ү�~���
��}�
_a�~��/�b�ʇF��G���_*#����H���;�Q���#A��Z�׶�N�J'�z�39SNi�*��*�;ӂ��y��o漴�����f��vR^�UҵT��2�|��D�Y��!P��62��~��1]�9t��b�bl��KA��5�+��F�����[B> w���=ŀ�����ܯ�
xN��ɔ�[�K���`[1�A;vY"N�,2JQ~1�J�|,�f�·���⑍:C����GJ��VK=betu���Q��+����`����8a�gI:���/+hZ]y6��w���.#2.�̩Y[�ѥ���r#��5��`+��",s��,����3���F_�s8Fr4E	��ě��C��$2��5�Х�1�@7L�b;�J}ѻ.�l��B��r�=^�$zW�i�+����;��"��m7��s�����3I�J�}�ͺ��-Z��gqR}�Iك!��D���wT���Y�t�V;c\�[<�R��c^���Yx�]��d��b&\�*��t� ��m���r�`z���Pw�s�������:D�q]FB;�E	NgL�TWu��ùG5������%����R0�Lp�7=��W��U�DX�k�2���c	:��%n{����?H���+�V0��$QU�߮�3xj���e�u3��t�\��@��P���aɪ73�U��UH�W�H��ع�`"ª֪�띉�&�d�L=�N͐�E�
n�Bq��.�l�C�X}g�}z�#���j���/b#0��@W�s�lE�,-�y��w;��J���P�z���@\?=뼙8]��(�T��:M�s��6%����C=�6jع{����AC���\N�ҁG�Ėj�]�j*�v�LI�<�g������p�⮯<�[����4;��%��|>���U��>;�kJ�x1IAҡ�2\����;ĭmH�+h>��n�YDg�i�^�H���Lx4����x`#��Y������ۧw�eY�1m����)F�D�+�f5�w����`t[�Ĥ��~�Y��/S��-�kCJ,�Vb�Ve,�{'Uk.���V,�W����ŝI�������w q�r���i�Ĳ3�a){�V8T8���ju�X�ե�:�⽴�P�'W� S9��Dsۊ)��MU�_Qz#���<�ӮNКbܐ,7�_l�9{�w�t�:�ٜS�pj�8��C�zrT�	�"�@`���
�s�)��p��8� y��N5[���Z�5�_��C�bԆz���#F��A���]�4��ͽ�:ыڜ4o%�ق�J�:#S::�S�૧��\ո)��p��f���ˮ��b�G��ڏ�7$a�,�p<��o�\+&*�J��	���I���)����P!��d����.���,��k�y��3�yq��^>�����@0Lg�J�������z���G�А�sWA�^ lj25" ��Q�u7�`�2��x«�3�>����X;�q���$t�H\�8�b�U�Y���IB�=J�y!0�����e�rZ{��b�E`�\&}]7p�WUDo��V��́�LR-׵�g'$�^���7�r��t��]�P�h��0�`�J��%���}��}1A�����t��3(�7)-Z��\�V�Z�B��+U�a�q�נIO�$ I?�$ I?���$�IO���$��$�	'��$ I?�B���$�	'�$ I?���$��IN$ I(B����$��IO���$��IO�H@��$�	'�H@�z��$���
�2��E�;h�6� ���9�>� ��zT�	D)D%$*)J*�
�
�QU
��H!R
B��)UR��@!HTH��"TRP
�AW���i)U�Z��]gL7wB;(c��(Vwt���R����������v�����M������m����^���[m�¨��n���ݯv����樛���6i�u���K��;�n�H�muM$Mk���5���TEA�m���f�K4:�2U��M֥n��L�J�5f�M��>���蹊��;� �S
_`|ݜwmt��i�v�4t�̫Q��z�����{R� J�^��+Gj��Ѣ�j�烧������K�(�v0��u�Mњ[k;aRkm�{� �x������ �t�+SA�/�m�z�6z������@gzjMh3���� #���PSݹG@9璴�u�����m��;d�π  7x� �� ��{p���wqp:��^������sU{9Y@��5�[����z䭬j=���ֵ���1;1)�؊��U����  y�W�5���G*)Ż

������(QE��QEQG��]�
 �B�	
��<P���
Ͼ�((P�}�o�����P�B�������
(P���n���j��q꽻�r��ݛ�  ]�x�� t)�{��Kֻ�K�U&��;��P�uW�����f�Ӈ���UC�
sK۸�T��ۺkTS�t��"WllU��<�A^�����B+��[ݽ��W6��˭���  �>x�֘;B�A��( j�n��2��t�r��v�Y��M)��@�Z�����AwV��V�N��=z4��U�=iV�+cM��K�v�   ���aM46+n�4�e���G��mC�uރ�^����hR��N���]*@S����zP�n��r{�z����f���u���K6�m�u�@��E��V�ժ�N�|  {悋��un�u΀5T�Qelͭ�tþ����Wf*���P+�(�v�T�P�X ��[��oi{68u���c骭��G:�lѽ{�/w� ����mZj��5���5�uv��&����Tޕ`ʀ]m��ԡ���Z��{�z�R����z�ѻ\�����S{�{�T�B���{^��)��û��Wcl8��>  {��� �����lz��%CM],k�,뺕 )I�nP�����y���IG�,unN��WW u��i0ү���eIJ� )�IIUC#���`���ښh  "��	JT @���U @�HS�D��#�?�ߍ������fx5�s�w���w3	bu��ȕ�&*�_up�Y�  =�=�w� �L � $	'� �$�� I �!!��{�����M���b!F��q�G#B"�(m<�7V��I�<��>ô�bD&��{W�kS��b
�E�P��a��ʽ�c������mT��x��u��{
qU�XoN�U�/v��1D�&���� D��I�i��cĩ;�����ʽ��֢�t��	�bf�-�0��[b�p���vڳ��퐅ڨ��l7(�v���S��i��A���״;MC��]O�|I)lӢ��,�I:ID�y(�Iʻ�%i���W"��mMAuax)���r�ǟF6��p��&»W!��*��P�0�!���G���C���r�5EV���(�X��-�++M�o5eD�Vw0SX*0g�>S@�H|`�J�ڎ<�G���wA� �wM�qh(��=�-�źk-U1cp���46�k���Z�2��cv��v晲�����v#Im*T�����j�r���:R�BR��*��`��E�n������\x��rZ
���U X,K����fmW1[�ZH9��wi@�pSoZ��B�Z�n��ACV�1�n9i�Vi.�T]!��DLl�: ()\&�i�浑�B�*��83 �1���<������i;{��Ԣ�Qx2ռ��Y���%�u�$�7�*�L�
.LҐ����c�v�T�#3h���,t��4��sF�Oq���`�2����X�Ӯ�4����B�����r9�PpVP7��mC$k%�M�lL'�t*:��9��ַ0غ6X�[A�Z)�<�����ۊ�Y���uRܕ*�)4ħ�Z�q���5��*fC���#6�(�rť�J߁v#�`R���)�cVRVt�D6���ZBN��&�e�sa���Bj®��Ҵm&i�{�l� .)tժ�&�wG�$XU��k6衖��u�*� � �v�Zfi'��WB�^4�t��C&R�D!D���-����t�vQ�"�.�Gn��x��v^沚�P��C륲�-�Mք�FϮ]i'�Z1���j�"x�-� 3���X�e�J�6Tc^<�;If�n�OXښ6�^V��Ɯ������Yՠ��yVȣ)�2�����)�[SF)��*]��m�.��؈m���/SW)��e�xinX#[n�hV�Q�zA��Au�����߶�6ޅ�[�i�.:,]a7��
�`��0H����
ͬ����pG ��x$�Z�l�1۹�q�N�U�_K��Z�]xh��������3FHH��a�uk+'�Pܷ`�򞳏N�&!��V��w+,!����� ���a�y�H`{1L�xަ�!
��U;�w ��Z�BZ� �ݔǏ��sni����(M����3t�ոɢ/Q�a�1�,���Z�<�Q��b��'�H"��b5g%JqC����`ޤ���$�i�4��1(&��۴�L;�j�f�U#Y�EÛm"�l7jŃ.�kB.ʶ�RY��6��Ϝm=е=�05���h���A��Z���4��р�����4���^�9�hg��(e��%��U݊K$��[/2�l����� ъ˼��#��i �����*p��+678h3D@֔c��`�x"ZvL����yY��+� �Fw��;]�M<̕1ˠ �bov�^D��nҠ��"��1�(���3sP��0��B�	H�92�;N|�f�H���Q�&�1� ����iyKdh-R�jR�ЫhU��˴޲l�7v@�۩z��Hpxh=Y7v�O%��"��̳�J�)U�%��@�v��CI����2^��oUG�� tӦ]�����)q�5���VC����`T2hhN%��s+2k�v�3 ��V4qB]�Qvw
���0��1Q��oF�[!��Pי�
��
� ��f�[rҩu{��۪��`��C"�{@G�5L��2=�Ш�4���(��7vjvي5-M��۫L U.:���5�3l	b���0:�s/(�Z��Mag]��(���j�q�aˍm0�Z��Q��Sie-*��W�#U�<�9r-X5����5��+q!�-�X���`��b�4�=n�&�`j�t֋[��Ŋ-m)���à�hQ
����I�|5Bs3�@*kM���#D��#/6�e��R�$e��1u��NXX�5KYln^S͇tF�M7Yf�q���.��pZN@��4hEì�H�[�$���V���2wP �M���n�G39�M����D�wN��B:S�B�Y!��n2��EB��`��U��e���'7-)�xYf����ӘNZ�eԣ{V��ܴ&�0�Y�A���^�fӥ2	
�.y���ѡѧO7L�(U�8��؏�D����*�J��ؼ�]Z�E�Tz����IX��N��f4��W�'�@e94�VU�5%@]��T&D���f]ڇ-���r�k��d%+r��)m��.�9����Ɋ�R���H��qLo^�T2��Y5Vs@����-:q��\�v�Yr����D�sG%�l[���Z�ZS��F�Y��{�j�h�Yb�4oiƵcTH1}��P[Uq��$k&�{F���[{Bi�ð��N��޽y� )R�ws^�t�4���٠̏kY �e4��A��
��,)�	q�	m]����5�]��D�t)��.��$7m�u[X�c,����ѧ�V�E�u��{��"��[��ކ�gV�y!�x+ ׆V�E]IZ~�a�J|�GB[&
V���B"�l��ӿ�F�A!m�V7wί�Fj��&Ґ%�ӗ&�Z���M�e��AE��bq�6~�-�ۀ�^#h��ì� F��ݚ	����w;RڂI�2M�BC/tS��'e�:�[e�Bի����������ʋ�ߌ{�E�s�]@��׃Yʙj�P9�����:�(�x���oe۫�H�4�֬Gf�
���4�J7��m�-�#%�h-бSK�eBf��&��VZ���5�e��ڳZ�IEh��t��7��h=-f���t�Tb
�oUh���j۩):��)+w#�+��b�S^����c݄l:�Ok���[m���r��Vn��M^
i�*tO$��x����f���'�C��~�%l,�o����g����	v*�W$1t�YOn��U��o7,(^�Yjԣ-�h��U�l��蹖c�B���[����G^&��(��mZ9)m����8��[yn[y�Z�2��d�6�:9v�hM����$�-pj:ư��#����n�����ϯ�h]1���� W0���۫4�$�I��!c�V���NŹ���d���V��Z��\�]%j,�r�K�x��J�wN��K
ե*z�ׁT����^7��`�9wT���46���$mfThҁ)mV�Zٺ�3%[���v-A��Ұ��$x������8n�e�wUr�7y�D ͠N�6�ڔ(G�Z�CK�qw�#���,� 7�
�&��v������T�+�7E�Zj`Tl�e�̔5ޜ�6��ϵ���ժsN0^+16qʏv[R��X�;�M|N��yL��9j��ؙ4,����C^5�I��N��VY�lY�r����YgX��Ae�[�.<ʁTJ��b���H"��ud86�C��XZMa��1Z�y*�m����(�;��Nn,5�];�gd���t.�Y R�dl��~���0��3J��hT+
�!ޕo~�X١FTz��I�@�v`�"��)xVպ`0e�2V�q���Z�J��-W�b+x7kf��w�a��{JG�0�:\����n�*�V�Zf,�.�CVrM1�R���k%*ik��*{*��FH�5��U6�b�����Y%i��a̩h�JD��Eڒ���/�Ћ�4.Y��a�
�
�hѳ��Z��M4i�n@��S+��N�-R���䶳)FpR�E���*��6�&ॉ^ݭ��귴�HS��X�M`�`��e<jt�Ϧ\5���3��^���f�e�Hd���w\׮JI W�9` �;��åf��M]4�ĳYvI�1�L�j�R8�M�hVn6�^� �Uy�6c0����P�aa�j� GB�t�@f\��Rz��*�*ջm}6��5tj�ۦ�&�h+M�"�D+RC2�Fkk�[X��v���a�n��5Yh�Jr�X��B��S[�Ki�J�h:����0e
 �
kM]al.|m�Y!4��twk7�J�)da��b�[b�-X�qַ�4[(��1��zn��,�  !S^6&� �����z�X�W��S9�W$���uf�+l�,�
��ϲ
���x���owo5Q��JF&�DH ʛJ$�����&^-�M�OuPơbf�B�G�� �[�]yX�Ƕ��� �u�c���c�Yxj
�&Q�
�Q�^�����J%�+��-�e��Yq �,c@�谄Ưfl��[����J��tNVKT�IH-�.���3�i�0`��/1����
Z�*�h��:Bݤ踄Y�	�ꂷ&�i2��E���1b�u�^�+n�N�:��oi��+�;t�%J��|���9��{e��m5w���@�;�r	�R�9n��$�e��
�V01/���J�¶�m���jZ���˦������vE1V6&b	��+yVTx(1�@��[��	�6U�l��$#M9�%��5m -٣�EQ,zu檒���@��t�9)c�r�z�t��h�a��6����WRT��M���D-�1/�"t��Ձfcn�����ҏ)Yq�ܽ0K����pD�d,��80cH^]��IMK#4��uRi�re]ڢ��=HJ�/H��Aڭ&��8��¥��e4��J�U�"��Lm^��$P4�5����P��E�0V�2�K^ތ1=1���w�u[���SnH�K�&�5��7*�yR���wH��jA��� �E^��k�Z�7�OC-�����2�ش(�v��YO~j�'dAG2V�2�qK�l\� M�h[�LEz�~{������\��Ɛ���Y�i�4kif	�jL�SE�G�i^��)V���J��ܓ��̀[yW���a�X�9��Ik���'I�j��Y��u�� $�s(iIl�z7eKŅe�[P��	2dN�kN֔��]�2-g9rN��J����įU��7� ͻ��F,�����"�%#R��gB�M6��];�������pbv�he$N�\Ոj֥��P�զaо���i�ě�c���ߵ��*���w1�������9��B�6�<Wiݦ�T.<��#��h!c��|�A!h�G7���JGm"r�h̵F�̳(	����ʆ�Y��v���1JKTF��*�}a�tl��ݕob��!/~9�W�>V*f	bM�YH�#�U�j�0r^�y�`�٘�F��.��v�tUM^32�hmC�S�.�7�����{����3(?�	ɚ��A�VB��YmQѴd�N�â��{)X%�h�@�e��!+�VY�x�괂
��݂2�b����-E/Q��.�!%H�C�t�`�X�k^�y�Ga�ГVB�� 7+t�N�Q�����&�z�7R�!�o2=*�Ǹ�2u�=��%�G�	w$5R�f��HGd��Bΰ�Lf*em�j�C�SFmmM�Ǉ2i�a���Ze�Z�r��ϒ�������Բ�M���ǖ `h�@�����srD�n݁u�Z��t��;a|�Z���ć�R�탔�ɛ �VZ�,ndɻ�#m0�[�9��Z��o.`Tn��X�����n��ݰ�a�hB����FT)�N�޶T[�i�m�i:{�o�̰�m�%k#u	-	�����ia��A[5�d�ܧP�Ӄb�^��(;X���l��2�����n�����[J�����»i���͡��Û\ȣ��Z2�"�ؑ%$2�!�)���P7��4�b��y&�%Q�H�(�8�:q7L��LlP�^�n�T�e@�`V]ɐۦ(�ѽ�6�wDT�"&T��ą#+MYh��+#$т�8��v�+u�!SWL��k�N�4��.�ާk� �����������ɰ����\!�V7-v�w�����l�º�RKB�Ti��˸��*��_fa�K7�TU�YsJD�N
KbO����kyPVR�.fL�jr��YB\���Y"���QN7��-�h�m�F8H�m��:�QVK��K%�$��ڊ��s)YJ�+�toum-�&ҕmZy�H ���O������9%F���j-�
��wM��v��hڸ"Z2�Sr��nV��6e�S4�(+s%Hw5��1�}>T�eͷ��h< �Va��n�wNk�2BXVK�8���O̫�X�	\�1LdT���� aD�;�i���w{��"�Ou�j�n�&��d��Ԕ�5D"v,];[AcQBf��X��� �y��T��5�����V�+V���	AH݀d�(m�$*�iX���
Ga4������VR!iǒ�y��.��V��̬^�ŕ�<[p0H�ȋ�-n1v/Z�]���3m�@lzum�T��))���JI@Hm�]��գW���E�PXb�t֙��E{�k5b�DL��عx�d�r�QÚ�OBm���Z�S�ɤ�
I}� +Neކ�+���[�}_������          �m��m��m��m��m��m��m��m��m��m��m��m��m��m�� ��)o����Ӎ�m�F�T�˽N�;�*�����"�7����I��\�d^8�on�,wFM�������7�[S��*�sf������%��u�b,�v�ú�⊶!7W�㑗�����	�R�Bg]��j���v
�:�jэ���Ðe���P���u�K���{�?N%o��c�n<f�t���\�;��X"d��|Ԣ7n
rWu����T/h�M���%H�
�Kx��@�y$��#��d%k��$�5n��V�H0�lÇK�O�Yǹև�2в�uڥ���.���N�zE�����#%�o9����m��ݛ.��t+��-�/;i��iK�����؄�ܣ�L<&�2����������:k�
d%��n����= b�:�Yx�l��<�j%,�v�:���u�Y����S)��oSO����{"eު�|���&��z�C�%c�*Ӳ���Z��]��,�O��A
TdE�Ȗ2����׬]5*���pt;�G�
�db���m:����ݽ�$�~�]�[�c�7��t.�@� �{]�D�8����,qL;�#`q��9��|ė��u�P���j&����W�P��aЍd8,nh9n^H�WQ���š�	�EP��t�r��V�)�о�찢�'� "���e�P�<�]Xwx��_
V��"��f�tC�m�Os2�yQ�n���H��1��XJf���ME�G�
��@���4�����܉y�j]�V�K�x�V�Ƨ�p�{a�+�?72-x����5��UM}�y}fͲ����mIM�	�g^ mU��ȽW� ╜�d*������ޜ,�]K>K.q��Mjo7���Y�و�p)�*8/��wZc6�v�+�U��1U�=Fl31�]���@�p7&F��3:���5�'Ƅ�]���8P0o?3�%��}�sc�`*����wZ&��<)l���+��B��6?���������C�]Z��o���}B�~G�g-Vb��J�k\�c�$(E[5��%��e5��Jٗt��F�6�;�m]κ�\+�F�Xd}�u�RO��N�].�a��_^��78.W0�k� �Mڨ��Ace��k2�yk�>6�۞���'DOOv�iZ�M�y�7e����+j�>�U�i�M'*tf����B��9��K��46Lt�e;?H�:�S��8z�Z��&>W�"i�Z�V��۰�Q8"�1U��o��d����=J����C���Y�<��R���W����d���b���沓s\��6�w�SZM�YT�K,�-�Z���Wm���e�B�l�.8��mūީB�9���0�<T(�X�����|qXK�^,p��I��YΥ��_f	/����a������4������JW5u>�YR�V�	�f����ʂ�W4z��wr6nR{L�ٲyk��L�U�ح���A�{F.v(��YE*;a��ʛo��Y��yή:�n���.�C��z�<r��u.�hf��s]�2�l&�͘�B���7D8��;ɭ�|l�bW�o��Ssk,r]]+II�mʓ�����o&Z5 .�eRX�p]�DA1$5V�}|Cيd[��X
i��ᕩ�Z�Z�f%�[�~2�e�Otj[Y��$�j�Tj��3���gW%B��Ȇ�g4aޫ&�dN��F����}/"�riXdXCע���_^�1�['��p�<�έ�h8�����Y�Χ�Ԝ�Gux%����ɜub���Uv�<�ң���z�(i�����v]��:ip&�Z.�/ Ԅ;��+{^,	�y0��o*��k�#3���w�c��To7y�홯���q+� �ɜ��Eu^�3ZU�2Y�jPH�Ԯφ�+)mu�Ux@�+�ݠ�	X���8=��rA���$3 W����6��|.��o`�r4��[O6fgt .���/�l}�u�<|��\8��j�`M�Z�N��Y�6g3C����Wc�nX��'n��E�ꉅqjKC}՚O=�]k�]��D6n�vy)����.vf�E��2�P��Q�Pg ��\�ͼ����m��:Z����У���v4��J��l��u�;t�`�Wo�.�s�9���o�	{+)�����]vZD+�q+���L��d�5yYa�ec�@�+��R��_upo<�*�Rkߞ���x����w{�mܹ��[��aHb�{�����Ա[��c��n5X���(�1�����1�)u��|�"��f�|�8�n��k�����h��n�H�����9�c�{,ղxr��.�[MR��X�L.��ɔ��J�R��b,1J�L-̄�v��ǆ-�;YIr���n�@Wa�Pn[�K)�@�5ǽq�lR��3]����B��vU��7¯�[q#ɜ
54��]��� ��枹�89��f�}1n`*T�Y���1�ó��M<ۣ:[��II`@��.��3�n�}3����zjI*W� �`�79h�T�}�
�%4/��<�i�c�Z����1e�j�2���T0Ӗ�N#8+/�l�'D�vL�3Ec�R��lux�̍��Uu9חv�a�t�<��7��4n�0ެ����<D�C]&ˏ�*i�4��Ĝ{;'���w>�4�N��s{��wGoRXL�����J��@��mf��LQJ�;]x^��]&3^MOwsi���������j��|N��2^�j�r�+H�'r�Y�
<!����:�O���BM�)�G�f+H���[#8��q�T���9�X� u'��Ӷ�U.WD�3P�J�<���]�M����Tk���8[k�]`�cBP�n(72!e߅GVS��R���c%I&P����i]�z(���R�--M�/.�@�Pi�`]eV�яmn���x�.=��.>Л���<WaF��]c����QA��c�RԊ�&ڟ^(Tz�vU��!U	f���)�S�Mٳ���Qˎ`��"�%M^$��Q�rnч�r��OJ��6�`z;7D�N�*՘���7Q�X�̞/�!�5�r���~���Y Tim���O�,��V���m6�=�[U�nK�v�g*���4t�&�	[�QD��}���ۆ�+uԬr�,����k��3y��8˥f�ts����J�ؐ�+��7lO�\U�Xs��r�n}mL��<F��{���}�cC1�OYP��{�t���%0%��+��s����j�5�7R-H��9�Ļ�{�B�+��G^OVGiufT�De�1§�ҍ9�#av��):�K9��f)�s*��?Y��h�;�4�n*^��Ԭ/-SN��tWپ�9"���ǯ7"��=���Y�f���Q�Ў.�uqzξ!��YfV�N�|���e
a��]��.s\ճ�p.�w�|�V�E�F2�⽂u�]��*�l���b�޾u��j�C�ʼf�)�a	���l��K�wN�"w�{��L_+� ��F��s�tWc�3v�ȟ@o,�#�ٺ}N��7���^���5�:8��i=[���6;��V�d�gg,�wa��8Q�G]]ed�|rI�,)� �M���W]r5deF��3j��߱%gT�a׵�C�HAy^4L2�*��X�Ѧ��_'7lR��eu�M�.
�2��E [b*ݼV�C�i�=C�89��CJ�I�d��{+'uZ0��Njm@9��bdBݧ�'`�W�t�H����1ox؃U��/z�h���t�q��.�X��)n�i��A�1]F͡J�����eH�i_ n Q�h'%�&sYܩ��8�v*��'4�9��uc.)R���7W� �ܩ{��*(.�m7��NS�bܾ
��p�9�I���g%�V۷&ԩ��[�{.�݀rd��N��op6��8��X/+��J]O���Шi��d �R`۩5���^MF0|L8�ٙM�"�I['Һ����9*8�����b�c��_,�s�%�h�\�v�w�2���265r���[�����y�i9ʒ�b�M�X&J������_5Q��w�����/h��b[�Jٻ���T�q5����n<�Iz�ӫ�����drGn�L�OO��Zh*�WY��.Ɏ����'r��GH���\x1����l��V����D���SX�Ghc��h�wg�God�_G�+tLZWv���B�F���߆����B�x�يzWWwP�;��fW�-�׏�P�X��&V�s���Yxƌb�C�.������I�_TB�Io�Rq�0:i���3�ϭ�S�Vxm�F���x�u�N����K�\�*��a��r�j��W�:=����h�!<H�*�e��+r���.S�R�V-B�vݍ�@��a/D{���'B���k�A�w���2M��#n-��c��;���Oϫ��2���^NdJ�y�ݎ���[w6�<*/2u-YZ�!��M��X�e����8^�W>2���r�R��|��&���s-13���%�TV.em�9A�@�B�"�hj���u�KQ��`֢6^G��_P�nX��:�p iB�����ފ+^�LY3����E3,O�)���ZU
C�5y��}s����]3m�7w�Jv��r˞��}S���y΍C�f�vv)���)���ڂ�}3��Od�n��)�Q�і�8��=#��Rh��Ja3
B�9�E.��qe�;��X�'Lʖ�dɛS����ʔ�='5�ُl��Kf�]��4��fnb��j�c����jˍμ���7��Ÿ����:��t��(&�i���.[8r��l�������f�h�VVQ�ϫm�wb�Iq�kO	��慌���Xt*_-u���7o���F�p��xv�㻀�q�r�u� �r��JRcK�O�����!���5��<�;Ws�R���Vb�MA\����Vq/s�jWD-���%^dw�ܝ��F�j�Ԧ�ko�j��Grl�݄�¼�Y}.K%��eι'�fW�/,�nԈ�3��^�������V�71*Ge
ϨmI�̠�A�1dq��N�M�����2�VC�PIoT=|����쭝z݀婗e��]予�&�u�Ģ܊q�eX�Օ���T@�b���fooA�j��B�d�4��0�^�?q��V��o��Vz#�h�d���N�(Fl��t7[�K^�Ŝ8�L4�jaf�B��]�2��J������^6X�ÜuS�9�D�׎]��s�@!�pz�hX�J�Á�).����$D*�;Bm`�e���P �f�36ꉽj��Hj)ع_9Uq�vY9yĝ˛��q����S�E&�ghi��M�s:�w�P��jz(��D��ñ��Yݘ�#rEVA��fئ��g��Ŵ�l���*�IN�ܥy�'�3�N�&.v�f���޷� $�9�@]��1�\�!R������S�9�R�a׻��X%S��]>`�Oќ2v���e�X��v}�!���f����V�Rz�S���������ne<��0�sA�J��r[��p�(u+P\V��(�	�����-��ϸ�6^��vE=k������n{6��%C�����&e1��Z��h�N�r��v�Ӭ��HM+9.��Dt{+o8��5���_�CZ��Me�0�$Ì�O��:����]��78�m��W��˜�d�D}�լ���LX}+L�m��J�B^�٦h?jY�ӧV�L̝�Χ\�zB�ŵ��%=��G%�:�q����yG^����N'@K�B|Sʱ�DX�q����%�69,�}�z,B��ov�k���УY/���B&]c�2 {Ն6��{L�Ot�lu;�oW���I��c�T�t�+�j������\����ӓ3P�Joc��n��$; Yr�S6y�Yˆ�<����`�wv�����_r�Nn*}v�<N��Cm�O>�5��>��Y7��=F�̢q�ܾ�� �i�W����gZ��tV&�͓�-;t駽թ��4 x�k�W��Pz	�T�/���ŋ)w6�z������s�Wd��1C3������mmC8��^�6#�]��i�w����1^�+�G���]0y����������^�沧�̾Z�[����zfր@N��&���U��3:�.F�+f����n_gkǁޥ*��Ȉ��J��V,��èӵA�����j��`]gg\RJx�	{y��&bl�[���v9K�b�J��c=A��#VU���;:�Ǝl�No��x��|���\SR8�7eΝS|��5u�+����.���N)�}p+[��	4q>Ž�V����t���p+���>w�ɦ��ݛK�M.�9�kZ�J��J�YC孉��"�$V�Yx%���g!&շz^��u�ʡ��ZՌ��d����(=��6(hw�b��� 	)<�33ywCQq��%�FY{�aL������5������+��:2�`s7K���7���̔�WfS��AwXhu��N����}z���-�?%��FI�P��6�#z�q33Y�f� ��d�a����|�nҪ����o,�H�p�i�ΐ���4Pw{Sr�u����]L�$ԓ{/(ٹ��='��eG�����=ǥۆ����\&�﫧a=�ӥ%Y:�����R�::磝6�۾�0��`�d:��,�әo'���k�Av�J����\������r�۸k|mH5�{��NKQ��Z�%�o�� I�N�ͥ:�rI$�I$�_�  xx{�� �
��M_��	<m���ur˅�P�uykz5��3:)��FgABU0�of^tr�5��l#�������Og<�Y�3nf���5��s�h���b�ݙn��nƶ�k@#4>��j\�/���E�y�w�g��^��[�,��i�r��=+*�GRK���f��U��sI�&`J�p�h�m!�t�v��`�6b�#tR���l���|%��������	ε��6=Q:ݗ�%[�M���ӪC��胶���"w�ʛ�ٲ�a�e�[MQ�B7Ae��rƊ�Ė�, L���{8�yAQϸ1��cU��>��d�h���X����w<��;�/�M9YCq�i�vyNx1��8^\Cn��@,�bm�֬���&��m�۲����4u��իAa��Mt����Z�PS���D�1��l[8�tYݳ��!2�qL�*�y��2<��HHdʂ&.ovtZ����ۏc.���k�����K�:��t8�t�]���D�%Z���%Ћ�4��5��)��>�Ŋ���0�*�.�<��6��
O=ZY�jz�u���j�e>9�Gs���
��̮�	�gH�Zp�2:�M\��u@�S�Ņ�.�ydZ�6vd�I�iV���`��91��r-U;�A�G��Ś����.=E�[p/�T�]���L̳�˃��J�I�0�+�����ddi��ŧYJ�t��x�+��x8��/zz.����J���Wq'ME(�bR7����+v���;g�V��^ez��JY�;u�@���@l����^oٔ�,��Si*@V-h}҃�qf]l!���AYG~Iգ[�|˽���w���&�^6z�臩������)�vԢ�ɦ�)�J�S�)����5���<-u�m8�o�O���=]���u�/�Z�U��`D�|2S<#�w_���[��qYen�Ė+�	=m��Y�v�qx񍏹d�r֠6*"�Գ&�hӍ��y��P��m�����BK���<�\|~��n��:��c��d3�ۮ��' �C[S�
�NS��gwO���PYZ�U��#î��i���tjc������G��2�-��2��g���Y�	�g<ʈ�.TӜ]	zR�N���;�o���WMj����F�gT��J�F\�tй�lѮbPJW���)Ҳ��:F�����*o��V�9�<7c4LƊ��&�-�A!��N��s�l)U�;J6�8�Z�,\Is�vRzV�O֦`�z�n��.λ��*��m�J�I��+gb�r�oy��g@��5+*��A`�vpf�*�\%۽�uu2k��3���([���-sO����j��D�*�W|h[\�쾕|�-��S���ݐ�jTt�KV�Zf�Q�b�)vK�P�+Yބ��M����U�����]��Ոu1�w5��v�o�=":y��;r�Ϸ5q41M�F��p��r��Vő�@\��EU�wd,٘I�#w6![��~
�7ĩ�r�@����}3O�b[o���M�X�}OU���L�6���a�t[;6��;S�0�=uz�:�$zU����ٷf��
On�;k��j\�t�����v���Qv�����M�j��V$F7M�(0��C�U"ĕ,���#'u�f�r�Ȍ.w*t�+����/s�<D�дt;i]հ��ō��~��0Vd�G��փa��v�R��$]�@�EQĬ����-����'��<�h&^�uǳ�<��m��b�;��љx�<jFesf�	LM��v��v�I��3�_u�P_�y�lx)���W��x0�&�����8�bx��Z�m�{+4�Zjŉ�����[�$���E۹�ԩ�#ˢ��a燍]�TB�9�ؓ�-���WG1��ܻ��S�)���9e���U;1Y��雗9Qņ���^�`*b΃��]Z�;R�:��N�¡Wc2� 	y�k�4�wQu5�4�\�ٔ$l|֝s����N�<�!n����Z�nX��<�4ee��٭�o$�.k���I-gqfv|H�%�@�
�]l��W|f+�f��\6��qm�SW[
�[x�������h��E�EB����2ɀ��q�9�+Tw�&%����c_V��]����|��TH6����n�@�1er�l�"��kZr���MP�;���؟��2���#t��z���P���N�70�N�������}�E\�1Ų�YM�ޙ;r^��2Mݭ��K��J�Y�];!�E��Y�}���p��7�����]ژ�;4�bG���i������Չ��:7}A��9>j���F\�y���<#3YE^�O�)I�F��=�t�N�CnGC稒�u� ��u�Qlsc����G�Py�^@�mE�A�#/�u�0bĆ^�\vc�pfZ�A媂�������C�i�p�P�Rq�������Yr��O���+!�սz'\��T�̥(���ݎټ�E�U
{V�*�㚧Q�S����PJ��� �\���QKA�Fn#9VJ�����7kn%u�;6���>���ݥ*{�VŸE��:��e#KOM5��U�oP��M��X��,r-��[�/���R�``��%�wY`�t�0��n���}Ç|��V˘��Z$wL<ΧP��ˆ�h/B���<���t�E���!�,`ƖV,̈́�J��4�0=r]�ζ���|x�2��j`�Β�4��7D5�'��w׳������%q�\ӏoG1pN��áS.މ;����͠��*��e
4N�9�]Lӯ*�QݽUa����|�n�Sł6l���-�ak.�hn��V�/\��W;:���9[u�Ѳ4�2�(�QFf�b*W7F�=�̀V����E�8i	�+m_`�Zhr����^�"� ���Sb�^+1VP։��(	/
�����]�X0�7AC���u����Nܽ�sФ�爻��p��g�"�h��y�ϻ2����7��ghaEy��ab�]�O9Ȼ�^.c6`�(���l��e|�-���ƪﵺ�+�B�ZVSk8�7���(!t.A�E�Ţ������e��ɑ��SYռRM}���1X�ʼ��F�wSǡ��H���VQ����k��HM[��IS�ګ��B���(^Rg;D�u&WeM�f��n!Ei��>�#��ؾO��ˑ�1�Ĥ�7g��N�x�7�!�b�md�f;��	u���5�N���NG�C�_yC¥y"�0�	��+�
|)��[/	�t�U-�d=t ��Le�2�ʏZ����,V�|�,�[R]3e����*I�w)R�ܺ���)|c�D�����l2� 9�r����b4ՂU��Y���"��֜j��]6^�ѺY st.�/ǭܳ�i�>l��'vݣxr�� �|�,��V��R�hhZ��2c�{ѱ!�*��j�I����d����*xۙB������ev#�$U��gn����y�J^���_c��&�T��[F+�z��7L֭{�U���[]ԛt	B������uuk�K���U�no2�'V�|�K�펌:�ݕ7..���ۮȐU�q�q�!
�Z�U�pG�KW��
�\�p�;���m%3��ܭNW.*)�J]�FJ��U�5�݂����J����/��;����r�[�� �_;�m���-�D��(e���"��'s��ﵬju���8o��R�V�a��Fo'qۥ�:mwwU�W &��£��� �΀�Ƞ��4Uց�4/A���������&[Dws��Q��q�6���o0�j�;�J)�v��L�F@z ���=T�܂�;0�?���!��P=N�܀iU��׻������B���PqWf�P��J*Λ�a�,hZ�id�"k4u��!J0�6o0ݴ�f���(
��`�ZI���Ow���å���}����]�Ex��P�I5t���۠/Rl�;�a�)d���i6جI�z�3N�پաy.�.�a���+��� ��y��l;]t,L@� ң]r��Tt,\A����V7`��P˽(Q�M
��� ��V�-(�n���)�af!�b5N�\8�@/���f�"�z����G%x^mH�v��C�J������h��T�BօQ��m�����C��u�����n� �w%mXw���uJ�O����o�S�j1��@WS���P`^��W���ERł��T*6����j�[��*�KU�/���yVj(KGS�Z��$.�����fs�C�(^T�ۼ4��߹�3��J�#/���,=A"m��u��R���1�)�n��+g,�9V�N��`,÷D��K�9���ۡ5ͷ�(�T�_T�j ���D��K�s�(��c��dG^Kx�..7�v������$
P��7
�1�b�����o�jn���Ё�q���F:���/gb�($.���A��գ��|W#
��/��W�p�L��G�mŲ�+4���b�51\3�������sYV��,sZ^P������6�H��X`�DJyܝ�	�~3�VE{��4Q�c���T)��-A��&��Vn�-���<�̥8�1 �gը�di�m��]2b��m��j��U,�K��o�wK�ݷ�F�ۄ�٢�b���Η���;Uy#� ).�9_8�RΩN�2�㫷3͈�˔��hO���n��Rl��x�C۝�0˾�jb���������ST.��}��
�`�u�/lCm!��j�&G�ȫ�8��cs1a���a-�,>��:n�fi�O*�&�;c�8��_/F��H{B�P��'o'y��.u
��v��EB���B�.��]j����-s�cz/��o����Y�e8"�f�w>���i��8%�Zn#�WEG�/�c[V�v�l\Ys��#۫��U��4m�Q����9�Kݵv��)�2��Awm��+W���t�ؙ�t�U�S��ś�}�*Ύ�-�9���Whq�ސ�S@v.��{J���%b"��:X�v�yD�<c��w��O
��v^�n�nĠ��L1�;~ǻz�	��wғ�^�yހ�	�� ��ֱJ���v��p
��Å��t�e�7�1�+���]�9.�+�-ô��iQ`&�u0Y,���J06��B`�"w��X��Ցl<,����T���Ӯ$<X�c{`Nq��'#J4���r����;$��:E�C��V�g�\~��h��J&?�[,$�Ռ���:A,�t�=���a�81f�!Ӯ��zS7�Vtc���[��{] ��Y�'Z���ujMr�e�)����1�ՃO�Gח���KB!�6�Ui(_tcd�*�%��Z$�r�̂H��L)�����-�T�����
R{F`"]���oV囡�t��!��Y�a�mU�����X�a��rh�p
�Da��^ֻS�V�����;ܣ�4Ls�ƒ�2�ߖ>T�O-�r_V��F��V�b���2Xr�PaRI��ӫ�k���J�zNG�̯���U���gT�4
3������݇�#�ʶ��w�5d��������J�(�˳�%��n<Q!Ƹ���]�W��hEMڋ��;��Xj-�"`M�n�^Ae���������E��X��y˳}	�qT�NqŲ����ts����^7\Ű:_oAγ!����P7��<��p�n����}]�t�N�K�r%�cr��DӂL�B2 ���#f݅K-�͓B�f���P�=�u�3;��Oo�k��җ-k���f65�]�}��]7��S�	NN�A�UmG��pPY�˂S��\͸j5��/%6N���t�"7òv\��C�*:��%tm$rFnv�y7%�]�퉽��Pⷶ,�t�$���jf���9M(��ޮ�s��h�h�!o��<G8�Ed� E��ӝ0R
.FIV�K�"h�~����)��ݨ�q���p�{Bc37�,����wk&��nVk廃���ᄁ�`3������KGS5��w �s��٪�j�X\ f�;�xv��j�a{��Gl�ZΰPض�5�gM��p��v�H'��3�8�ΖN�d��w����I]a��!���jQ��� >���d�m.�#e��u��ݹu�8yI��5.R8�טu�P��u�����#$]�omWA;�� ���xE=�Ҕ��m�)ޚ������ZZ�[�¹Ӥ�%]e�(�L	�'�SIB­�|;/��X2���o)q��'eV�%��CE;�2(���4q�(]w�,��F�fr&����e�=Vx���Ю�+�Lg*�Bȅ�B��j�7�&�n���K#,�^�v�蚏�n��	n<'�T� �0s��˰z��w��[u�	�n�T�;Y���ڤz�=N�������J���|�0*X�8������cw8�ǡ�gv%55%�\Wn8�&ud��T8q��͎k 9}Ɲ��aa���	j�[-9�N�Y�5��hU6�Pd��o��.#�4!֨͆��	�(�Irg��=�86�蓚�n�3-C�Q<���T�蚋��G�v䩼��CIu�U�
�]-����ɶN*���˛�x���3j�INd����շʓM�{,�{�3/��ؕvk� ��KD�܊���� �{���*�/:0��V�X�1u���αl���r���ʴ�!��ٺ��;_HFgc��۩�X�eJ1�s�et�w�kD3 �)A�1���y��oe3:��1�l�mui?V�G-��M�t�nI(M�v|��GP#W7�gS7�t<߾�^7��� 	I�j&s�w��� ^�����r��4����vMdr��4���r24�ʭ��>fQ؜㝂�R���j��"t6ulp�LA&�N�jV��w�s��I*�� R���ŕ{w|��:�9�u|��#���C�i�M�8w��SdU�qɶ�
oUA������P2��aU���_�H�-�2?��|����>���}ͺ)Y�^?u�=F�r�t�>��/�s����M����^4�v�f5k Ŝ�"*4kV@������6x��6�R��ĦnN�]ګfu �����ي�v��o{�Ǖgh�<���Խ����E�gg�h���������B��cO>2�U}�Z� �w�J���-!�Z�E�和�o�i|�VT���K�����MB�U|��sm�OC��"0�й��u2�rQ����P��.R����\�"b ���>����D�Q�=��*!GD�}\J�d�ۦ@��V��Z�}���<��;��"(S��Fa�Q�uwl���^�.zVP��T@]oW/�A�v�w%�:�j��X��?Y��6�m�Y�n�-����=�Ț.�u�sلR�Ku'��2P�͆!��z���]H
\5t�ʔ�B�o�;��ġ�c8��U%�k��]�Ug6)����Jzʯ�<�V��g%}J�f�IN��zI>��Qb�`�`��!V1V�F �ZDA��2�*��Gv��EPDĩ�TTEX,�=KR(z�v6UU�J��,\k��Pݲ��T��&$G��`PPS�($�H�,h�BQE�F@R���"�*�������Hm�mX�	��c�M��*9BT*f5Y"��ME4�3�Y7h�¡2���4�����C��g+�UT��_ւ��ID"�J0DC�6�!�yM�0F
Y;���q��d�s+(
((��J�a�8�X:h�ʐ�
ȱH�J���8ʁP�"!8�@GL'5M'PQq&���IRqn�R��c
��&�欆�,b�U�,�SI��T�
 >��S�`g]fU�ꀕ�"k����;�y����nL�I3��Ѩu��0f$k��/I��ɹ�_x��i�z}�^�o+�؞L#[�
�H*��D*�UEn� v�¾�A�Eh�-Q����:��k�]�<�t'Rċ˚/���P5�n+X�<��N���E��c��^ź������ݵ&K��I�lb��}sJ p�"�2��v5҈�k]i�G2����wV��,R�V���ß��8�t\"L�Jf,�*yMX�]�<���n�T�7����![�]{f�W,�ȋ��l9-���KC��UJ�-����u���K�螒h5tȰ5��9����P��WkcH���P[B8��C�ŷ�&�{��F�#{Hv��t���X
%�q�Jr�BU*/�Q��Q�.�s�r���0�yh�ê����h�,��R��/e�;Ўx���~�'�W���6j5���-I{{�B$�=O��O��]"��=ns���Y��^He����Q9�0&��dۤ�\�\�L6���=
�G��n��*�X�����JF�b�����><+d��l��w1֫�;F��-��:��8\�V�yEV��[�ļOn!�l��#>M�n:�5�ۚ�K�xif��m���]G6�n:�!�ܝ���B?g��'�/�KP��l@.5[9���0"쭷��&ô�H#���(�;��k�{���`PN�������R��u�gMX�F�zgJ���:皤�G�B�koc���t�IM1)�="�ߠ�LӯN@a)�=T�o��*���Iw&������W��e9��Ux��5䩝��Y��Tf��"�v 1�|����c૷�t�9݋�����8�̈��cu'�)d3�b�����2/֒H����%�}��"A��#�g<h�ɫ���eܷ ����t��C�^hϠ�՝թN�s��X�^�}[���c�9�r���yi��P�]CѪ\@�`��Q��ݹ�ԟ��5f͛p�`�s���3N�td`uQ�
{��V��t����&�{5��ڎY\c�p���=�!�{F���Bё�k���`w�\o�R�9�(��8ռ��,�W'�t�iUa�r��iW�׷fl5:f��5��2;Eeג���~�S��iJ���@�����."�ޟO)�q��>�pq�~y^)*�{C�2WMZ:� ,�g�"�wi�BG��3��i�MJ�]�/Q\��NB������Z��9�fmv>Ŕ��z��"�i�N(Ewb�ut����Cw�#�6L�W^�k@����j/���6.r���Z�]F`��jcٯ탇[��!�{d�9%�e�ީX�V�eP���������|�DZ�m�!�#�7��:0�s����-b� �����1q��ẒȾ�CI��v��X�\`W��7����J7��S؞F�N�s����[Bp�n��(L���\|v�*c�:�9*z��|�+֪	��+��3�wmP���h3a9�Z���~��3\.8�dr�~�PN�M�a>78�u��`�z��k�G�,.�Vt���M1�b�^��v"��}�i�D"��Y���x�°�t�=bةS��:R�,�~\(�yx��һ�kCtD9�d�H�w�N�AEˮ�;~�t�pC5�!���R�XHM��>��Y�R����X�=ȧ/<�tCA�{�!�j�>GnG��RJ���pvl���u@xc��`�;;#k'Q�k�j�+U.�� G�K�x�+D�PN�>��;�T��)n��\~��U}N��:��K�j���kS�������I�dLPNɃ%�z9�Λ�����F��?{�h�{P�����(�;ٴ���h���=�qΈ��.6��ŭ-�5V���bUf�\��7���
!�Kj��A��Wb�㗪�i�;�������R��ѧ|*��s�f����B:��ŵ���)�3��RvN�&
H���-�����F:';�tA˦�ؿ|�A*lł���i���	a�4Y�B�#�Fl�K$�"�2�V�+-�����B������p�'S�x�q�D�\S�Z�7]/����<�9��NU����X4.3�~ޔk��a��A�N�l�j�����M���Q�Q���e-��͞�j��u\�0��7#TP�T��s�i�۠��9}�h[1rv�t�c��f�R��4�N��:�)r�N4;���j�U��V�n��q�[��Ҝ�wh��F8�&�H��5)E-��Y�`��.@�"��@��2�fq�����6�F>�=���)���=�����@�2�4`�L񼺠����k4 C�S��~�ዸ�O�|�?ps͎=�~�	�_Y�(C���*��i�t����t#�ׄ.�����Y������^c��6'/)��w�j:j3SZ��aEEe���BŹ��un�]{[�z��Su1�:�3+z+��s�R{i�>WVj%V�hW;_��W���G�R�f�p �~N�H����<h糨p�kq]JSQ�i�@�\R{!���k�x�U��Sy�n�|_:�Q$���P|j���zJ���W��ݺU0�Q�5k���)*��	Ҳ��{D���N�RX�æ�l^K{V7��Z����{W������͔��(Kk/�J%I�^�tϪ_F_��&[���=�������~��Z������	<�ç
;�A���NؚY4,�g��i-=�}����$����q�Un�D�/�f�G �Mą9���P�S�L���$��߆v��3�x·uOfF�c[)6Z5R��YyOoV�8�r�DS�Ւ^�����gQG'G|��r53
�:�fN��s�T)�94�y�J���%-�k�mx���trjP�n4+�{���[d!��]����^��Ğ���j�y���\W�c�x���=7�y��V|���)&�x��~�q���n޽ٿ+�>O�1���R����ll�U��'3�rԬ��-Y�e�J�%�]絽O^d��(Ynz����N=&b7���5�vweN�Y��ZG�UŃ-u�Ǭ>�HOuj��E
�bw9 4m�{��SA�ɶ�J��O�9՝����c��[''��GIVv-ݜj��Q��4*�[���}z'L �7���mw";������o+�E�C�1cs��&�2߆s��;����H#��ʵ����J���J����Ԣ��;V%Uz���y��8�V`���s���)��ZT�e	�]�j�S�!�T.��_f�����r�.x���˲��]�;Y,>db�,:{g����Z�[L���	ۜ{ݩT��Wf�O;v��Z����E�3R�������b�X�a��*��yiu��!oP��%L\��+ʜHL˥�L���e�,�t6��:w���Ŋ�OJ�e�Ǻ��{^�0��,PI���U�f��R����dJ�mSܨ�W�ni�лW����3����[�����5n�`�Y�ϭs��$�\�)�W�w�i=����U�������L�ȇ.�WU�{=&��`Ƿ����^_��ܧ��P�v�Ø (:�eMN9��Iv��w֡ν�2ē*�b��a�|�b�3"V��8���u�v���ם�p�)�~AM�� _uy�'{�>����\�X�㔡��WH�ϰi��^�r��KVp���Z��r�g-�G��LwE������T\�`�j��;��fX�w��O3%�:1\D�9����G'¥��9��36a�jY�L��۱Mr1![^5<��S�eS� �����&��Fw�V�U]mo��R��i�	9�ޞSu���Z�����������z���� ��Ơnnԫ�K�R�<
�؛��f��+U<���o^�ۼ9M��WR���31s��K�-�'���J������|��ˇ��k��>��}�l�K�T%���`t�>����b5��<�3)��s"�ڱ�Un�{���w5EL����%58�q��XΊ	������,F��OW���Ǆ��V�5Oe�j�{C�^ދ�֓�K5�o���X�8��<$t>�w��Ns�y�'a�G�yt������]xv��݉�b�ⴇ����7�.�L7�fښ��g-��-ȥX�U�Y�[IK��5P(Je3D,�G�b]8��E��˝ʈ)P�O��uh*U��1M�[���>���<h�ᚚr����i�w�1�m-�+���+{ f�2V�ñ��r�us�t#G_f��`����i�X8�3-rAZ�V��V����5�LK�:���tn`E5�w�����,#����S\qW�f:�<����o U��E�C:�y�1�b�gCrf�i��\>9�.N���_����'���w2a.��S��4�A��(0����j�E�7�ނۃ���]�5\�fP-v��f�9S�C�c46�ç���=���BN��Tj�y"��瑖dy�1��I���w4��J�H�sh���4�<�����y�:�\#��f����δbU�v{�69��b��W���'q�ޥ��g�p��J��R}<7�֎�X���ݝ�
�0&�qq9�M#؆OnC���tBڧ�:�П^&k٪yJ�v�zx�h��y1�ɽ�|����IfK��	����lJUWCdRfo�7��3�=��^a�	j[	���m�;�m�ٰ���e�u�Õ�.�H��������:�5b\3C&VKǘ�ev���n��K�\Bх���S�G�v��:5�.��Z��Sv6L�oO�9Z������8�ݦ9u�+x��Ձ�)����YeҾf
��on�:8�������k���%K���{s;��)�k�"����z�޵���lc7����9��}�Ɯ{��D9�/{�9�Qh��v�ɱ�����H͵j��e{5S����z�����r��j��Q������R��sv�.�T:�wF'���9������2��I�w	=��M�Z��h��������R+i�z��,����U;�f��8�vJ�XL�8�7���(#~�.����R�2ķ�%`�8�cͯC��٥���͇�m���������������.{�5�6�Crj���1s�+EI�޷�8�i8��O�!;��@$�yӉ�/����N���yr�ɸʼ��J��2�_m���,>)�h�=�PV�[S]��X���/��q���r���yw�/.���2�c[)6Z5S�>&\(��*aS���
��y���AA��B�=t��B��s�\�S1![d:T���i���H���;�ۈ�ǔ4�z7��,0K��=������.ˁ<Z��Y9�T��,1P��7�(��S��gm+�:��wm;�v`�[
��1իn��+�0��Y����Oӽ�d��i�o5f<9��]4�S��N�b�]��vv�;]Wy-�c�r9�X���H(g�{�o/����f�=e�|�u�V�Mc���7��'_DH�{����O�:�����P{pS��H<�1�<��k��ԳB�n޽ٰ���2����Jv�l��4�+�E��ú�x�����bSʞkx�׻6�"���D���#(��qVZZ��îg�F��u�H��u����>�o�����s�My�=w��C��y댺ws���.�8��8�ps�YDh1[/oU�M�M�7�� �e:�<$t.�~:����u�!u;Ʋ�S�͇kcfns�N�-:JjW?sJ�ư�?v�D��߶бj�^B��P��K��W�ܞ0���\_��^mHr��R�/6ŪJ�nK���9n��-�15��hOTŉk`PT�33�ё�T^a�w������Y�I1��hH�.�\v���� �r����T&�Q%��HvX�J�d�����\�ӈ�+q�]w&L;طd�_9����/����t�y9���^,�XJ�jq<��%C&:���n�f��p��V]ڋ&�e ����SIp�����ӆ�+��޼�5�)RF���]*QKW�r��f	�u�۴�w�M�ו�0���c���-큍aj�r�'b�2��Auc3�AK�u����1{p��_cJE�bɓwM�ht�sec�g6�u�c�٦3��0��Q�<{-<����rJޱ��'M��a;p�A��˄�J�<�&���-jz���v�è��/!�����ژ̭�ť���>�b�WW�5h(pC�;�=e�A��{VnV��
��8<ǁ>�Y�Rd�-2�G!��'Ku���:��^tO%���MuM˚�:);�e�]R�F��#Q���oTV7_C¦�:ݬ�{�������H�'Zghe���gU��Tk�A�u�*N=˨����t��bw�����y0�NٽQw`�*��f��V��t��
����,�>�/�}F��ծ䕧)Zv���$�I[Ok��c��,p{�ud+HܓK�1�Y�8�jl�Wc@^*�j��B(Z�S�K�[R�E���r�M>?v<\1:�N����b�V��b��@��6�` �uz&�J�E˳��!�ȇfҊ,]�|ɲ1�}4m9o�X+t�y�:�.�L$�����kM���,��������Pȕ�r�v�$sp����]�t�ؕ܎���v���K �K��sɛ��r	)�X�%5�wᮨ�cz7��D��nk���;<~<79Պn��.ҴgGsmdG�u5hL�x�E|Yk�������&=#.�ǲ��:]��� c�1�|k8lc��������3~��/��s���qS�3l���M�	*9���7t2���r��;3`�h�P�D�6N.��+�r#w��b4���ʄ�}w�:-���-;��R�vWO����i9{aY��F�&�l����Kb����V:�T�{Fr	Eg��t y�I{�7Ճ�H�v���8[�4��{�ҮLU�u�f��§q&	P�oa�P�����_BD��<r8/�1�/b����'i�rVa�Q���/�F�oU������3�-���dt��%1�_p���=t��2��7Vu}��w'����H��$��ւ�����[ӈM�պ'Nr���k3#�v_e�vsF7$|�5*"�w6R��tSo��d�sD:��¢WϞ��AMDƔ���ζ�B)<�T���ӫ�g�����+������^M%�=�p�\�� dmC��k��\h*��+C[o�Ө�O�(����u7L�Ҍ]�vn{��o�K`�,9����<<�S(��,�������]_�{�9
�c1�䒰Y �,�
�RJ��P��C	R�d ]3lċ�T1����\��P"�RLaPU�fTH�f�TRHT��BV���
�ł�Ơ�)*B�8׉��V2�x�`m�I8�1��duV)��svV�&9���X,1X�ٌ
����K"�N8�#[��T+|J��(M���x°�!�x͠Er�3v���P�����:LqYRO�Bm��VV�LP�'�3i��0*B��WyE��)&$�4�R�_��r��i4��T����R� bm1H��A@����dXCm%CI�M"�r�������~���NR�p�N=��Yf]��Nm��wyŉ��h�Ke�o]�ز��Ԛ{���E��Q���r�L_����1[>�s����� �u�%�	=�^t�A���1�S�3�ɓ,<����;�j���f�n$l�#��(4r6N5�zB���WՏ�v�����]��g�<V���Au^���f�G%�v���)}]�~�������]5�./z�߳��T~���"�����m�[�����s��3&����q��:�̜Ŧ��K�jA ��9_{_[���jG�����c�{�7�b@���l�<��z�w �S���9+�s	�^$(�<���֭T�wvm���Y6�mt�o}[���eߺ��{tu]�>�L��j���ޫ�׻2v�D�φ�g��D�+:��|��~��-�~�D9[B�m/�|��i��r�OS�LWV8��ĝ�_.�Ͼo~���Jt)��r��8�5��bT�*�pmҪ���۹l�KL҄/NoM)�Ȱ�i�w��b�>W��q�&�TT��� :ٖ��⣾��% �۾C)�ꨧ%q��*wXߕЫ�m��h[}�N�z��м��;��))�Ʋ�qF7H#��A��ۙ�����3��e��2��.�q�j�z��]�x/L��*��uݿl�k沀�sW��[�7�q�^�h����Gg�8�̪��sME��H/���G���ﮀ�U��z_T
o���9��gi���T�td��w敟�F�^�jkk>�?^��Ij�r���|nsY��Z�s�3h_����(�}�y�mz�)�8�fc�6����"M�7W�vJy�Z�m|����$93�d��?@�� w���J�^�ឳ�����\�RI�-�<A2�L��_8�)2�t����T�*�H��ߦ�M��HE+;ڙ���}��-q��@4r�s�t:�Cj�O4N�RsR�xJ�ٴ������wf�ϵ o���f�BD���|Uo��k<{̩��}m����c{>��믕f�쿤k kF%[�a�ۛ�$%�q˘�Z2�B� �e����t�h�^�}lZE��S�S���P�������.�*��.�n�pV�W�Kg����WЉ��xhӺ�W�*KC�L�<@g5��S�3��1u�����/��6p����٠5��lqת��B�|GE��.���_W׼�~��d`w[���fݪ��(^4/s��kGib�#�ǫ(xOi���T�3�S�c��[U��:��L��R9J��%[u�&9�����Ӝ�ˌ�]I��vlxd&���x�.��_>�S{���|u mt�`�;�#oo�]�=��[�>j����a��6��,�9u�����s�d�L���6'��n�G���~ƪ��#���_����rJ�t.�B�!I�BZ��ԩ���e�S�Y�]n��e�;��[��ꗇ�=�x4��ׯ=�����->��(7��Kk�R�C�+�m;Y����/z榠�<������HIa�9xt�>��lR�V�qջ�Yz�)�ź��,�:/�z������5P!���r��R�2����R�8��`�]���Qsfm�F�,W���3�I*b��ą&Us:dT�����^��=3����3Mn_u�Μ�e+n�Ѵ�����_D,��3c��Am��nfJ޽W�v�-��]
�ƥ��R����ŝW�;�lz;)[�f7�����o�0��;�_*k���u�oو�]�x��D pNr�dS}ۋg��ϧ���u*��=϶%z+t�yC��u�k}9�f�j������~������XQ��w����♦�A�&�T�1���_'Y+�$N���\�P��z���>؆��(Ｋvgځ�lD�٦����oDs����H�k��%�ӼNn��z���M�˔(� k>����\l���Ǹ�,�+gr�o3'�:-����׋�n�O�:���V�٢�ԫ�֜O��z���.^5ͳ���?@7�<�ɓ�"iά�P���4$g���4�d���W��:��n��ٵxS��ڿJT8�h��:X���J:0� [H�k���r��5�O^d���g���r�P�=��g:�T�d,b�)���F���H弯�u�kT����oAE^n`Й��L�P�}��	m���.3�N�ƅ�g��G����d�J:�N:6��[[��7ӊ�E���H$um��x��ܜ�q��~�kU�GL�C���N7�`�?�g{ڛt��ݻG�`.,��s�)�"�
��n�$�v8a[3)>��=�p矏-�]����3���$F���u���t���ՐtVj�3�_�A�|W�u��1�,�_�w�1��ھ����sz�3��+�a����b���͘�L�̚n����x�m�kW�����@��2��ʕ�l8z�ulu)�w=E�O
�aiݽ�p�h���!���8�̺���nN���չ�r��5-�[7֞�f:�k�[��K��.\8��Ў�?A�m�a��iq�f��lM<������dcq;,H�-��\ʬ��ǯgl��T���PXǱ"�cp�7*�E]��M戁��<!nlP��;py�[�Q��|!�̦j�y�.�A�D�^Ky����Pn�����J�,��;��dw1�yr0�gZ�ɷ���q9��,f�Sy�Q�yS�q� $=�����*��хnގ{�7�bu�D��͕!����SΕu$W'*�d�������o�o���YW%t���if�e}걽Tj
j��[OSɢ��2Q|U�e��mD&��&iਮ��nr�޳zMv`�lw+Z�D$�V2�"E�V��������t:�|�i����{)��X��U��^��=�G)��ko�U�{��`5�"�Ȥ�\��]�4�FRݍH��5[T�]!��3Y�yJ�V��z�r���j./t��g�o���-8ǽ85J��I��H�u���`)v+0�ǣ�ռf-=��ǽ� ;fD%,�Z-�ۨ��.2/��sНYU,�	�KĞOe^Ob]��(�v��	��B}л�5m��rw��]	�)�qڢ���v%w�
y��U+X� c�Jg�����S��FN�;��L�r�K�]{~���R+9���W��!i�iE`�pS�ubb*.դ���E���jŹ��W.��f��-V�)��y<�ڡx��O�D���3���R�2�)H��̷���!�C�b.��F���Cpdy��X�(���C�9>o��9O���L-ٷW�<�<{�U#\_��e�\��NS�0��t+�!~�֩�����ʅj�Õ�Ig=05e���i�%���*̞�kR�P�ZH�R}u<��\����60贎��-�{[x�c��[�I]M.=0w
.���9+��`ƍE1���>Mą&]�k+��&�w�;��1���+�R��'yt�gg��^����h�A�&<��t!�q���S�w�+��.wο<Syu�r7X1�L�M��T�������Y&�Bͧx���ս�
�4��Co,J�<�ٲ��:��F;i�ۘ��?s�����:��K�9ޫ�=��^-�\�"�Y��U�Z:��i�����v�g"�s7��m�H���l�M[T���z����'�	Y	�J�7��o���;��v�V���a�ݛ
��MFV3�ւ����z�+��92��}�Lz�����+���Tݎ��a��.��J8s�D5�.�t���R��Ȋ`4��K|1*�mH弑wݬgCa�J�w�:���d����<����)Tf�]O���c��j�)����w�qHEoo�w�Ӆ���w�b� v(9-���)��ת�q���`H�V�Q�,��)�B���*odźU���%쨅7Q������<�~LC��c���B`t��IW
���x�@Z���i&��]�8�\����w���w�":����!����^^v�l��Y�w��}���mO����Q�{��ۇ�ӵr��q���,:e��66�Əek�x�B��"���-�%/yF���u��n�W��&C�,:j�祽�X�5�"���]���Z�����Z]fq�/6��A%LCyC��*�3�}R�2�R�(�f�9��s��e���f׸1�[��48��ˮ�Y3{�Hy��[<�>�tu+�&�Mz�����8�g�X�)������06V
�Kζ��3;�9�Uyc��W�ԋ˦�vdj[~I��gx��14�����{=&�W��ʥ5��x�yrތ�B����r&A�L��_a>f�y�6�H�mx�����'�{��JS�U����
{�0�N����~������ z��<��h�`�������W��h���,���������<���>�P33�tHUd�tx���-�]x�@/+��>ܾO'6�$9c��������J�..��caO'u�]����(F��<:E�����<�h7cY
��)�u-<�y[�I,ؔ�~$x�O9������i�ٽ#��c��U4׻6���2����-uv�~�վƌ�fW��w�E}�&�]�䧕<�kz����;F%�ف���gx�ᔝX�7ޮ������d:�=5�ZWC���y"��G���t������԰��!]�_�������3B�8�S^'���#�ϫ�B��~Q��XΊ�ҕC(H�]�έ���C�+��[�׵��n��9y�qz��υf7m򹱬##�aўp����,ZF]�ȗ�ϋ�cuS��,Gu�j�ݮ@W���>���2��a�5+pѽ��{\>ʂ����g,��"��X�hB͢܄�1r���*q!3.�^�y�Sj��Nn�LNaEF�[K*�)�#�0�כ@�u�K���Y��E]Sʵ�>B>�>�
?���Ւ�?Zu'/���0�7��DcU3b4sdr�]2�iǼ��7&=<*�9��M�򌩎� r�d�����ѹ����FP7����̈�Aʅ�4C�{�'�]�U�(r+;2�n-�dz��u1�{� ǵ7��S��V�bhr�R	�7�g7ݛ��nj߼�$A$�|	���u9��%:v�ɜ����<􅎇���߬���.?z���L*��g��2�~]�$I�h�����5�y-���c`�ӕw�.��������y6�4�a��j���=�@ϧ�:�&�6Y�I/^�o=ƘJ����uf�
ju�ִa[���no��'_DN�G]Q۩٬�{Y�Z�jX�޻U�U����Ô�v���n��ݕU��)�E����ې�j38���[T`��Bo�9�G)Z��|���2X!�Z��0��&�kvUYĔe=��aJ�cdRfE�F��p�NMjy�T<+�:����v��Xm�N{��t_F}�;-=C�+�j�{}���}rs��;��]���!�́v�;Ѯ+�2�C(OB�V"h"f�ka[C��E[�P��^%���S�v�+���ҙ�|�
;2z77(e�N�v�POn�`O6���k�-�9M6��u�YؚS,*���t�_I��5�����cwюڹBB�fs��3���q�[�<�" �}�I$l�}!����!Gv���C39Ի��À����$�ɔ��Fͻ����>2,aƺ���f�ꁜߍcZ�Kb�WkEk�/B��������1I36�J��N��� %=���[&y�[�f[����>O�~��خ�:W;eN��C�5ԧQ�H���c,���ǽmm\�Z���S��Mev<!	�����s/PE|ʁaW7�ݐ���r�N��:D5{}�"_g�����ƒ�^9�s���uŽ�4\��Rf_��򰞥�f��!�@+�*�٥�.���t��BOU��m��t�'����FscӺ���Ί�O�1��	g�����a���^����h��1=qu�^#|L?Y���`Hj���-��媽qP��͍����x>룀�
��(�;����2U�n�(��J�ށ�6��/25&�i��#���G�wK����t)d6\G��lBP��WP%�Q�%��3Na��f�٦�i+LN����[ķ��b����87�uШ-TI@��<*��	3"�A�Ҥ���U�3xѲк��'k/*�Ɛ��K��c��3%�w��ݺ-��h�2��]r ��ʓ����`�ec�*;	���xhU�ӄ���� ƽK�Y�Z
�H�oݓ75ZN,���P^���j��"�kweX쒺�:�\��C���E���mE&�sRӺS�a���}�N;�v9�/	��v���'0'*�ov�EZ|2����4�^nP�g-5+����i����N�ܨ�V�!\*��@	T�ݡ��m�U��9���[W�:�jY���̈́wz~:ֈ�YH\IP�Τ�M�v��u��7@n0������z΍�%o���u���֍ظ�P����/�W(eJ��p|kCk:�U��z�XD6ڳ�Ǘ��ٹ���u�������7�l;�nbᰄ���kQ$��[��]77�N���R��8S�[}�S�����ѧ�6��Foz�`���R�Og���ɧ(���ɞ��/�[W��/��֦�"q%�I.C�v�̡SE>�Hvؠ�5�w��q�B���r�����}NN6���Rg�b�l�]��s�/�������*�/�/�S�����f��?3��guME���ݑ/8cW7iF@U�.�ī�`˾�ik�4�{�+{�hi�f�����е��
ә�*#w�rʸ
��#�+�]��.1uwE�6�s�Y��$�罵��ﾏ��K��wNh/�+���&��g�">z���'Ԁ�4�l:�-<�-���JJL�1{x�w��_(3N�Ӗ�#Ԯ�m�p����p��^u-�#$l�J*3��$�W��9����ᇲd���&��̰�6 �P�+�+4�R���@]ǌ�l��R(iY+$2��4�W2�k&ٌ��HbE+��m6�1�((T�
��
�&$�
�YMd�!X��+�I8��4!D`��c&�I�۽j�RT+�8�$4ȵ�����q14��U8�Vm�ڳYd�+�۫�d�E��a����0��cRT*c1���5J�c=L@X�m��E-���.~ȱC-1&30�6[tœ������4歵EIKIXU�r�X�����Y4��bJ�e�-�D�X6��ۊ���(�f�`T�bՋ1��)���j�QG
bJ���!�
�(����LN3a�L�&��%ChT���r�U�R��&&�Q%�\��P���VV�*����*cZɴ���Y,��°+XV��m3)9���FE*�V��"��3v�c=�	�7�~�&.8���s�o���]`�ǳ��7۷��<݋Y�j�WG�*��`P֕L��@�e1X�5)-�Ml�꯫Q���G��:v���9�{j�B����+T���
~��}��eAq$�]���&ص�B�am�6إ���\�څ�^-�KU�7�SA��][�}n��J�w��-aӵ+�,K{V)O��*��k�U6�Dz��ݻ��-��~lJ��\`
L��ol��ڥ�WjE��tR�֡u=��k���N<��0���[��A���Re׺ex�7*�AB�Sq�w0�Lj2����_ؗ�2Ѹ8`���Έ���,���U;\�e���o3�^]7��#X1����5�ܾ't�ǌN�\���>�f�H�0
yU�M�l���k#Z1*�=��3M��V�\'Ԋx����`s=�b9��6�:���	�hP�S�mU84�Rz�4��bqk�w�x�����Oc_De��4-��u]�"�2��{�����vԒg�u�1�\|�oǁ�N��7��w:r�ufA������\�w�:�z��ٳ�%�}e����~S�h����-~�Ǿ^�r�uu3�F2�%��`��0�z�J������ݣ~��D�(�)����{���r��c��{~mڰ����+�)���V��R�Cmt��h|6���w���H񴴻޺䧕7c��_�{�n�)B�]hc:���;�t�Y{�i�]��Xt�3"�ZĦ�.[��cXΆ��f�mM�aX�}��+ͼY��b�S������P�SO7��qR9*͝;>Mgk����,5���(:+6�����T:k+��>-�K����8������)�I�k�m0��~�N9}�J��jEm7sׯ���LH���t󵵱��R�yM�
��d9�æ}R�2�)T܉�n�`��C���ރ�{�{7L���:[��N\��K��K����iިjgl藹=ʦ�l�U�_y�1>�-�	=���5{�7a��HƵ̘�:�-���k�k�j|/-��dcq#e��)���	q�q�9�e�������ͨ�%��i����U�p������ܵqj�m�j�8,U���X�f_y,�xhve��Py,�]I"�.M�#�h�9[f4�d 7�d��(�Θ�+��Y� ��4X�Б���:e�$�<^n�J�^���竴t�_}U�>x�Jq��폜�mt�<6��t�+��^T���#P1���nh�FHy:����k��r�l��"py+.����pz���/.[ܹC)�;ԗuz�*��j��.�Ga�������(��+*��F�mf��� �2_;u�Z�y�}3��W ���[�����6���e?@0�ɚ<�Df����"X�˪m��Q�
��y��~��q~=�6O5��ku�w��vs�XqU9�O(v�v���k��ܩ��[�~z�g�ϖK�:�_5�(9�E���
pW�yW��Rg�F��t9��eJ�?t��3�����O���4�͇nAJ�t.�bۘ��ϭ;W�V�[yI��I����;�ʾ��`ps��`�8z���;zw&���W	�SoB��}��.ȉǽ�C5O�f6�*��##�@XtO�>�{zWN	��:��R��y&�1O��\i����q��ݾ��Ʌ]<]p�%u�v86�����|���+�w�Ir�ey֘�qJcq�(����\!o��i����VӳGN��!�Y�7b�8ud�R�)��T�dv�I�)��W/����c)�s��������ỡ��z�ܾ��ѐ�>Xt����.'��Ƴl��w�VX�ݠ,_H�8�mY�[��1bZ��N$i�2�\�3�O7Z��i��i���W��]"��Y�μ��!,;��d�F��������صt#Տ
�Ay�������Z��xZ��3��7�v�꺵���R�|L�)3�gɸ���;@�ٹT�+�jo.�g#�ڦ�B1Q��;,s�����F���k�:m(=y~��i�ʣX/cj�FҦ9n��|�fl�k3&��c�H�sm�},��SV���/������lmʺ}Y��xe���Z1>V��=ۛ�=�d�C������x�~�]c�x�y���{�*3[3T�v���n�U��7.�T���-�<>�A3'!��-]s^�׾F��h_&wٮyJ�W���T;L�T�a�߳٤z�fu��h=+'K�B��m���[=7���v`@���2�%G\��y��x�'�i��pM1��K:���I�%���ex*K���ϫZ4���K-�'����O2�$��uT���w�n�N�յ���b�S�����0^�\�����&��׻6�2���ӁB�v6i3|��4�'�ݰ��瞆{#�Y��P��y��zi7ё�;-1l+�f�)�iR	/Z��cUV���Vn;�tRe��2���v	�4E�����2�yL�S�N���%���
y���sz���sq�[t�jy�����,|��ʨ��_ջ	�v��n�ׂ����-��$�l�%�!�xt��}��ՋR+k˽�Y�s�myri�K]㦩.�Ŷ�5P!�L��8f;bׄ��b�qŹ�������>Q׮���1?ޠ��(6�N$)2����\>��T�ڢz�Շ��YԌt��<�2<�|�����c��)��e7�ˡ�k(�����TWX�А]���=�s���YEע-�^�ľ)�h���yo����,�yW�k�½�uKT-�q�pt�����Ј�I��.İ�p�����jM��ם۔VǙ�}�w�2�(�]����[R�2�wQ�{��Υ[;׽�\
Ǚp�ֽ�$*�������Xp Z<�^7s���ة��նR�� �+:����PC*��Ϳ� ^]7�vg�������f�ѻ�{1��}�K��M��e˿?;Zu(钅�]7^͔(e�b��U�����.�vs�Z�{͜=���i��<�5�#*�	�^�Qh�)�#"`�V>��-��ת.^?sm��� ��7�uߞC�����W�kSA�^�"��R��]��۵o^쪳�	���z��ҕ����d����W�����2��^��JySw��ͽ�t�I<��� 6�Ӟ2���|Qq�]S�"�ڿbUV�-��u��gF-}�]�#7L�������n���E�Oh]OT.2-u�Ĳ���S����35ڞe�}�;X��́o�)�:a����E�d.��1<L.�;/�NV=��m_nj��R���?t�:e��:VeJ��?xV{˞B���05"�k�)_ܷ���\�s�ze�5��	��|�o{*V�ԨRPǾ�@8=���F�*��:15w:��)T��vV�YKs\�,�ܐ�s�E�7�	�prVL��h`ב%����{�y;����;����i˽k�Dr_{��͵<�9k��k>�-��^�w����|S!��[�����y�^婲!&��^�Qm<;`��u�ڇ�^2�y%LCyC��&W3���Twq�O�o籩gM���V�l�f�AcwKb�O`ӧ�Ω�G�����[��wܸ������b]��yMh�3 cq#e��3���΍�����ʝ���g��K�pB*���_��k��4��(Ｉ���*66MʻZ�f�_~O�������a�.�������z�˔w^s�fL�E��-vGs�+��
�4�ɷ��-��g6��a��W��d�b���;�H��k�C/�T�h�^>��8{�e?@2�\�3!�S�o^)���3����^"��zox�ee뵶�[���ͅxmu���5<v&�Q��cl�ھ����Z��f�;�g��P¥����R� �I��S �	Q:zI�*Uۗ�%Ʈ�Т�����6+���Q�xp���~r��~���Q��������74�v��f��s��o�'d�&R��O��O>�W^e�Fx�%�po�����5�;x�f8���諭��������g�o��;fa8Ynz�Z����M���'�m�f�{"��ԡ�+���v;ֵM�ے�!]�\5�I���Na�*�Z�vmx�{{��9�[�潬gEy�J��8���V�e��T�'�PSpg��b|+�|��_����>����\ް���Jâ|���%�]��ȵ�0���b�ĦXb��S�]{b��k�+�n���o����Ѱ��&ov��fnWo838Qnop��[b����k�m܏$��������2�
�X�ϋ��[0�3�3R�2%^�L��/F��2ڣ�R5x"zh��sE-��?'���D�2����ڲ'֜���c�����EJ��|��}Fm�nS�yY�tO���A����,.�A���f�SȺA���*q��a�JkO\���bb;�:Ѹ3��X]xt�Pz����ڳJ�Y������g�a������N`͆�F�
�*��_d�7��i���ǻ7ff�C��a-�'4oUؗj��]�JЇ
C � �����5;G��-�F�Aw
�4��}��x�n�j޽�}|��Jǐ�q��ށB�Ag�ß�0���%7�)/��Vs�zٗ:�gx;R.���>�{S0�gZ�ɸ�Q�%5�F+�Sz{�����1cto+�I�l�^�Z�Z1![�c�����u^$r�g͞�!�y"�{�2��T"d״��:����}����Ǜݬ5YiI�Y=�S���owf�ؑ��1���U�A���/�;��;k7J��s���ŶD��1��Ϗ���U�;�*�բ��e]��Rd��3��[zD���[���yt����l���k����]�+靮����AjF�׮Z���d���f��3�Og�w�Z���B#�7
�R�Jwgm)�R��~���U���Ĳ�j�O5�|�oXゲ����;Z౵���e	�}�Jͻ�A��в;�>uZ��]&���� ��g[V���t�@ot�i
Bæ\��~:������Y���]?WMDL�dW�Zzglכ�2����ǝr)�l�&���w"?I?��ފ�ۺC��{;�?*h6l���q��5(���l��&(D.�&D[�
f�=o�U�;�i�0np��|��}e��T��¶�4�*��������R䘴�n�6����	|e3-aӠT���%��Ʒ�e�����źw�4r�zj��1�!4�0�o`9p���������K sn����[�8�!�e����1�9�H�-���M��Re��5�B��͚��r�P��q�z�w�i=�-;�hlX|S4��3��7ΦJ�$dK�NK����`y��4�"������I�c��Q��W)V�l���a�c���st����yC�M�l�����yYͻ	���o
�|���0��v��͆��c؉�l��Nj/�����znR[�.`��n�~z���X|��X���ݛObu�D�l�I[8��n����=f�Z���t�^S�ӎt�t�Cn���ݛW�SQ�1���(�=T�y�7�e0l��z�ղj#Nw���>�M��y����۴k�[���r������ܖ|�̮3Mq�F�Y�6�¹��.��w�s�ydqD�kD���:bv�=��{O%w.����+}�����p��5�Nd)��*�(f�R�1;�]�ARg���5�Z�M��q�)�g	x`�7��v7�X\��jk���jGΖ[����nZ�����/�����ڽ@��i#Fov�� c*�}�9.Q����_>�Z�{���n�OA�z���[rL�:��5z���<�CǹOκ�m;��D���o{��I^�5I����6xL�N+ma蘋Xf�@��3���u�I�q\a\.���v�k�5g2oa�y�F��h7V�a�mbڕ�y'��yFź�ͱ�������d���,[e$#���LZ���1m�P��W��4��;�w5rvE4r�X ����o��R��șj�b"��S����( �]ڹ����}�5W P�����mrPf��#C@΂��	���l�b��z��Eh5��ͭ�]*	OWr����;�eخ���P�:wv�2�ް�6� �^�#K��<�����<���ֳ��R�e����9�^k���[��q���2�i l���]�w>�䛡V{�f���Vڽ䬕�˓�R�ɷ{`�wq�u*cc���q۽��eu[9Սx�����7i!��5�KA	�4�rÇ�Y���<�b��x����J>�r�T�qh.���^W8���x�R�q��U�G+Ov��[����Eu�0=���|���[m����ԫ�j�FA���X�Ĉ͗��hoj<Z��L=F��P�ջ�m�A	�f���(3&7��\�*�)�g�ֵҎd�F8x!Ɂ���M/�t8�iz�jY��4	s��f��8�FY陔�]�'V������t���|L�����|Mb�l�y!��Qv/��Jl�Ź�;�+^`�Q�ӻ�� >tr����մ�U��� �b��4aTWV%���ӗ.���G����ڱ��|�1i�́�l��I:��f=ˬ��l{�q��8/5�80f��n��8ݬ�b����Wl��vr/�5"dF�g�[u-�[���Ӛ%ne����e��N���ѺĠ����>�E�)������/&�ڐ���W��v/�9�S�:���{���6eG���k=���N���x���+7�a�����
�FtǕ�q"�
�K���ᎎ��Gw7$"~���۳Y\x��B��c-�V�M�Z-������ȴ,Et�{k�Pf\�}}�1Vt�+o�H]\��+
l2h�j�(M��i���N�hC��{D�t2Fk���\��T�í�VU��Qb
�m\����s�4�c��/R�Q��KV���4��h&�i��B��c�Y7�Eq�C������+�:���ݶ�|J�i�L6V�]dd��	FfF�Yh��g����KV��]�rW`��A��#�T*��CJ��Q����M3m3)+!�o{�����&��1ģ
�VM9�����m1%H��
�(��f0�P�)m��a��-�SH�i��͔4�Sl�E0� �/7�6��,]��
_[:��%TI*�9ea4�+��+*���Kf�� q�Ět��+�&%d�4ʩXQ��q�ԊTY�����P16�P���Tt�(TAdR,1%Tr�T8��\��m�1���	uL��&	5h)1�4�y`�M��ۦ
���W2�Lf �b	�SfՓ2�(�[b5.�Xm�b���I�[k<J�m�������a�Y�-E*C�1��G(K���u�1�dEb�P�+!Y��k0���"��m�HUo7]sO�k���vy>��{ك�xnW�x"�{}�.�nUΣ���6oγ��t�}���U���*��Up��Y6��� ����W���t�ȅ����Sͺ4��:V����3�����֭>o9dY�{N�`��
|yBлE�oj�z�.3�{"46�����#e��١W\���w�q�[��xgC�#Vh��P��~#Ry{H��+;�Ύg�'��<�^��a~޳���,l-�,Z���![�G/c���j�-詨��.�9�W���7P+���C�,:f�la*^i�܅鉨%��MD_,����qױf��!����!���t�T�N7�/tc��p��"cp����XK"�����Y��נ�Ct�($���HNQÜ�ݶ����ׇ�3��;t3ڲU'�NNR�{t��cq;,I�t���uʬ�|�b��NY�nID�NC�t�(m�q�h��y�x��@f�	��q�\��ƪ�-���jˠ��ל��B���>� J�S<Fzޙq����O��/w�;63����
'�F.]kR�-�/��k#:֑�8ƌ;U�3!�E�s҃�X;w`A�ܵJ[򵔸Q��;[hWe�q�(Z;y�n �^ V�.�.c�l_8�^W\�:R���������I���F���F�L�m��y�7�ű�g6��:����S3|��	Q�Gpy�+Q�����ܼ�k�m�5�a� �IG7����{��c�/u�w;=A�}�#�����{5H�7��o��v��˽zܷ
��F�fv�ԆNvڌ��i�u�,tֱ>�H׆k���,tظ�T�߬�AY�Xv������}y����c	�s�-�5e9'���gv��Y��<�ֵM�rR�(t.�Zͺ���+����ԋ1��� jW��;���7��F�c:+�JT!�'�v�զ�4kq�Y�7x��9n"ԭƲ�T�cw��\ް�?r��a(n\��\��/���c����E�}e�v#�p��g�_L���N���wU���3lZ�)�xϪ^ᾇ�b�֜U�6�,��mw/V�s��H�F�3�|��;%X�-���w��MbRk�@6��T��u#��f���U�L�����V�R�Z�ح(�(�ٱ0&�&�^C�侃ȝ�:&5��^˗�WI�u�Fc"�'��y��8a�T�dFjH�Wsh�U�e�Ξ�qLb����WI���W�mdO����L�ظ�t'P�*���f�Bn��\�<����	R�}m�(Ro`ӧ�T3{F�N��ɽ�U��;�ǽ8��(�����#�^m	���[��2����v�o�f]�
��c�88դ��vƣm������q�=ܙh�� �]6e�蜑m�Y��h�q�]��e�כ��0�]�`ߵ3�e���|LX� ��I�h�Β�[2 ;�ʔR�ݶV��{~[(P�R5��F5[��Df��a\k�H$}:�M&g��ϟ@2����T<��h����f�������550��}ܝ9N"���>>m�>�3���\ק�׻O0ux]�7ɒ�s̠c�6&E^u�Se�R��ST�CoU��vm�	(��աB����oڔTm�E�=<�]��j뚐9W..����7�l��,�S�����j{�mDS3�0Vb*�A��ٸh�~�y�v����i^읶�לElܺt0>�O�΍)|�S#�]����g�6�[�Ç2#&:�U<Q�ܥs�0Zr�}_��Ƶ�T/n�N�����ѩ������,ZH_��ݸ���W�8v��s��� M�|�/�,��ܪ�ϯ��Ī�m�弬(�v5�蠙lT�Ț��3�6�4�6�aA�o�[B�z�W��+@f��]��\�' �ڢl��.��ss� �ל�Ǆ���o�j�Q�x!u�N�;��o=^@��������1�&N�碷/�\�`��v؟�J|�_e'hl��.���e�vr���_��n�T�2��K��J������X��h�-C8��]�����>F�{�& D	�<a�����望:�'��Ԟ2b;��	�LM}��Ւ|��܅aǈ�d���G��;�P�(��U��nn�UW�����Q~r0��>D>�!���P�&��p:�<Ce̓���=��u���l�p��&ZhO��>��9� �������v�vv�k�η�<�|�aXx�2����g���I�!��2q	��6�RC�� ���s�IRd�rN��h�X|�֠l;��~d�O��������^�ݫ��c��{���{�>�${�A��2&���R!�~aϷ�u���'?Y�!�C\��q�u����&�jy�IRg�d��I������Y�������]��R]��t�����0@�䕓�8�=��T�O�}��BbMOl8�̃�Ra�����8��|�l�gR?Y�M2|���8����p%���K��SJ�+et��ˉ�{T=z�J���D Y�񭽫�8Ẹ��8*M-۬��+�S+�*�Ё/%b85:��l{g.�T�e�+f�{b�*�wZ�p՗uG ]D�EFޡy�@�.��h`���ښ1dLA}Ы l"{z/#5i�V�a/�������<o�>��s�(�{�k�'�g�^�8w�0<I�I���E�S!��x���M{�C�<Hi���O��aûÈc$��SL�"�wz��W�o�&�|�]�o���2='�D����O}̒m��w$��'����'�?'X��!�4���C�C���b~9�
�P�!�f}��!��=��oZ�>��u\���_	 �{ȁ��0��L��P���OZ�g��2h��j����RO���:���w̝Hx���p��C�!S_w�C�7�����:Pf/�K-�-�*{�[�}�}� o��P�I�7�mI��:�������$��8��6����!����Bu�I�?3�;ܝHx���=����?wΨ�jq�:����=t��P�N��u��M�x�8g��!��m�O�=�����Xq����'��m�s�I�ߨx���x������K�������
>�����|�3�wC�&��>C>E���d>I�'���;�:���Ւz§̞���ϲ�8�I�����i�����i��q���:�wm|���t��t�2O�`yڲOP��h(�O��w!Y=E���0�a�'��H|��Y�XO�*u&�RO���B���w��,��w���#�$z��;�'�P�͟���2����:��L�z��4�����%M~��$�4}��yl�r�P=Iơ�y� Ͻ��cb�����j�X��XɃ	��>��}Bz�Ձ�g���a�C�'��By�<��2u�I�}�:�l����I=ISA�r��߰��'��#��~O�;^�_�Fw�_��>@��<a���0��^$���n�P��	����~g���a?'�yu�u�>�ϐ�'Qd�k�'RxɈ���	�K���sӯ�S0������b���o�kq]Yo�(ޱ�J���5��k����Vɽ*�=�Ž�3�3��
�JfX��8���D���ֵ9�{��c킞�/��^-�n�ݫ��9tv���]hڴ�����Tt���vR������.���x	�O��]}Ǟ���Ւm����Y=jB��X��qj����1���NY�+<B|�`~eC��Y�I�.d�D�{� �|}�'ޭ��GdO�R�UoU����8ɍN�7�<I��nwy����0�ٓN$��i!���WԚ|M'� �t�!���i��P?��8ì�O�y�I�4����y�f���{C-�j�Ub����;Oq��}��)*g����*6�]��%f�~a]8���N2u�&Ϸ��.����Ci�i
�� �=C�<����P*~a��a�H}is0��a�I:θ��t����|�zy�]~�~���/@SĞ�0�`�I1&���m�Ȳ�5v}u'YP�Rc6w�%tȱN:g���Jʓ�~�i��Ld�+��d*n��T9�8M0����� Y@|4�#wMN��������O=�2TS�
����4��r�'�LC�K�y�R
qS��Rw,Ă������ĝq�öÖ��P�T�y�4��@Į����1��4}����AG#�${c�\Nd^��{�k�{�{�Y��3���s6�$���&�E��<f1d�Ұ��f�8ʟ2ny����*r�$��H)�7�d6�'�SL�{f'��'"���G�L��y�=���v������gk���OX|�d��w�<jz��1�;�?!��C�g?Y�4�E%I���:a�d����V0���6��Ǫy�Nj���x����Y���F����P$)�v�.X�������<@����ީӿ�'�1��z��['���4���㤞3�~��!��'þa�,�AO�����l:�*�S�Y:ʇr�P=t�O�o�Ͻg�g�G���ӕ!�~���v_�<�w�����ޓ�i?��� )�����:�x��&ӓ���O�+M��8钢��8N��=ev��9N}�H|��a��?"� ��79O�d�Y�a��:�'\f3Y������dl�){}������x0@�>����}LO�d����d�M����!���:Ͳz������u%`_��3L��(=���,��*{�aO�S���n�P�'�y�w�c� � YY2�/Pz��Di�2�{��U�H�Q��81�Y����R��i���U<-���y��p�e�;�e����.�ww�z�����6��r�#w�������_PB�r��T{�,�Uƍ��I,ؔ�{�  *���u�c��$��"H�$w@J#�Q|?0��~I����8���p<g���g��y�zìğ��Ś`x��'���u���l*>E% j��fς>A�U��s���A�]�����[���6��htʻt������SԜ����_a4��8�l�3��C�>��h��@��y��6��C��i=O�~t�i�j� ��13��ui �������CO���j~ֹ������u�Ns�
�0�,�C�d��e���Ͱ>k"��*�L��T7-<B���&2l��4��?e<d��%a�8�}���{��g̕��}ɶOY^2i�}�m���r^�4�q�ge&<��L{��� �l�S�o�d.�嘁�S�������\��Ƴs�LA`|ԛO��2|�P:�8��1�j��i��<���4�RVGz�����fk\����7��k�|�O�3�K��'M�6��+L��;��N������W[�:�}�M�2{n$�ގ�m�&�L�옝@��<�E�m!��nr�!Y������X�La�c>��y����z�:�|�=���+�S�P�~C�c�k��B�Ȥ�{�Z��M��	�N���o��ێ�1���͡�?e��S�~é6��6�݆���Hp����7Ә�w*���W/}���g���
��[:~�bx��n�~�ϝ$�O3XVE� ��jN��uT<;����*�l�p+�dSY�i?8Ɍ�eN{�
��o���3�:ͤ�2���7���.��~�X�ww�[��Q�� Q�}r4�!=@����'�m�%E=g�1��������PėD��I�]�Ӽ�$�,��1&ÿ`i1��4���ą�5�{��b�C�g�����_�禷꽎�:Ўπ�8�>g�H�����ԩ��!����O�Y<g�O�S�M!ԕ�6�4�{E���eb����E@��ʚ�쓭� ��g�d6�d��~§�
�I��k�:��Q��>�����R]v�����H� �$}�Ć�&�C�<f l3�]$?Zx��c���Vi����s�9�3�u����>�&Щ�Xr{t������,�ea��?8����߽���>� ~�[�����#�eLq��� k�!�p��6i^{����)-۶��Őz��Z�W��>��k�%�Y�f=�1o[������N@�D��#_�1y�m�
��D�k{Us�]]�A�޶]��ٻۣ]�;8���mœ��F�����S��O\+��� i�0?�{��*�����Y�ʞ~�39H)����6����Hj׶O���g��d��v�Ro��i�Ȳ�7ˉ�'S|�+��2��.	���|i�f��ݸc�|>��gŞ�VOs�ٴ�!S��LO��r�i=Cܦ��l4��+'����� ��*z;�TSo{��l���CٖqH(z��<�|������c F�}������Y����LzO������>q&Ͼͳi���{�C�T�{�'SL>aP��d�6��T�O���N2x�ɉ���yCI*$����=k6�|����d������fs���n���w�s��~��T
��/Zu���Af���4�2}n$��CԜv��
|�_~����C����XM~g�ĝ�t��l�OC�Ͳ|��$�܁$
>d>�����
��C�[�����w�k��&�I�8�.YX5����
��*kvu��\@�����Ԝ��'?SH|���9���$k߰<g�����`i:���@�r�S��:o�}����y��輶Pn{_�2��$p'��L�;=���=La�)�]$;l�2���st�`|�1��=d����I�6��OYRz�2��@�=IXo��#�{+&1s�n�2ݔ�<υ���c���Ӿ�P4��W��Q� ��}��'ȸ���Xi!�~�1�,O�?8���~vͤ>��5g]!Ĩ,�٤R��N~�3� ��4��^un��;�߭-�~����+'Y:}�O7Cԕ��u�>k6�ug���OYX���2T����߰�c'��Avwy:�i�'��/�LH/����AO�6r��'��<>�ٓ��F�*��TW\�������
!�~f!�X|�!�l�ܚd�+g���C�8�Oӝ�;�N!SH���Cl��yܕ���~�V��3���|͡�Me���Ad��/r�P���pD�3�����s)
�^���V{�AO^O�M'�<LT��C����0��m'Y���M&�uT=��T�Oi���Hv�4�j��&0>j~��W����� �_:�s�Ƅv��}ⲯ��kWQ(�^&n6�`L��R�pn�q5���ţ�5��NSUh��}������rZ����O��Z;�6�mxrٓ7Œh�;�7�s�ڔܧ���B�,���H7\���d5S�nZ5����g�����xw���G����2}����#�@�s���C䕟��W�
���a�1���̢�@��2�f�N��ACs�\&�d�.$�{����əN�:Ɏ'�O{����'7|����<�΅t�$=�:wY
�%Ad�}��=J��7��N��~J��쟘m��V?S�~���|��i�k4�t~�i�Y�ْvҠT���bx}��Q���ySj�F7]�{�����bJ�dո��r����Y?8��S�6{�q&�Lgq� �q�����I֤?Z�f�>ed��?:O�qgP�=�!��<��L`e����O|��*�x;���c�7�Q@Y1��i��+���u%f����]�;�I�1%C]�O�2���0YP��5H.�i=a�1Pϩ��q?�mI�u��bA�d�#/�4�����h�쏀>I�c��4��l���4�r�v��H�gY+;�f�q
�v��;��%eI��>��SH$�ݡP��z�Y�fH���3r�E$� ��A�v��㚧�ԫ�}OK�2}>G)�x����.!��&$=�My��6�S���w6���m9��']��T���x�����ɶOP4�g���1��4����`V}�#�@�F�	R�`�Ϯ��۴�r���5�a����d����1����\���O�:ܤ堡�J�2{�f�
Ax~���Ă�'﵄_�q�i���'wH"3I���jC-8_���c`�O�-��#)o�}����>}�t�!�1�!��jq!�I�/�q�`z�nr�a�P�=f�|¿8��i��T:��_�
��*O~�q�i
���p4Ρ�>Ձ�f�[����ԫ����H� �0�"$��� ��17���cğ3�?wy4���<E�5��AO�x��?Y�Y����g)�4�r�??8ȱg̗�d�3I>B���6��*O��8e��O���WCĮ����Ez��'P+���0�>f:gr��u��g��6��r���Y�>I}�z����p$<�6�{�i=a�T��O\f$7��jZ��)������*�:>9�|��%	ܽ���|��c߶��6�B
�"�iY5m�����|��Nܼ0�W���ÞУ�0���r�5e"�N[�ѕ�U:�ª��B�&E]]�,w���8m��w�ӨSwJ�+l�X�^�[S
�������菢"6�M79���2@D����|}c熓�z�>e��I�=����y�Ri��Y����n������'�������z���C�g�M!�J��a�ق��>�׮�?' �y�W�O߆�W�h�Y�(�Gº@Q����C�7�̛`|Ԇ�~֤�+'YYý�z�>C�ͧ��*C�I��~�J�J�����0+"��]�����8��������͟��s���{s����&�P��/�W���w�B���&3�8�5d�1>@������m ����G�??�u��a�;��Ұ�w;�M��&&nv�*,��k����_~���~��^{߫�΅f��)1�{���,�Þ���T�!]�4��Vl�!uO*'<��C��Nj� ���3�&"�@�~�}��m�'Q���_�� |G�G�D��v+��E�{�?y����;� �2ӧ{���i?3�Z�����;�ơ��>�z���X��VOYX~ݝM&3�d���4��3(u%w=��4����ʟz���{�VX]0.���}��W���k>b��J�߻�d��<d�r��0!�J�O�ar� �s��Ӊ8��Hs0è�&�Iɾ`n�D4�6�0>j����u���]���I$ I��r�_C���Γ��,Y��?3䆭'{�'�����u�E|�~�Vi��Ӊ�i6��T4�j���0*a��f��s�B���g�P�]�*u���s��<*�d"�Q�9�m����^8�7��Om�O㈠(+���f�
bO�SL:�*CW��ԟ2�ܤ�w�J�"Ř��wl��&'~�����Wܰ�~�<@�{��&�@�$q�y4���>�n~��^&]g�|�x�Xi<N�n�2TS�
��a�i�'���*I~�y3�-H)<�Z��f$�Ͼԝx��3rw2����~J��w0+P1+���
>��A�Vgk��}Zշ����=N3����,�'��(z���f�ĕ��]���5�B���<f��}iX~f2m�>d�w5�AC�J�/rO�Ă�G��i�O�SL���ɤ��6EO�ʙ�#�u�o�: �SF���k	R��h��ѝ��NV_\���x�|����\�8L����������֭��P�7��p������[�v(�R�ݤD�ׅ����}��V��vfa3'g-xq�l��+���e��å�.����h��:�0�u]:��Ӧ&,eveouXe��toh�O���M�5��r���wF�7A�o�:�Uot<n�T�R��XtܻǧN_��R�t.� ]�bc�9��s����imb��U�V|^�Ҿ)�5v�8�K��=�y�x����?
>h�xi��	Q�V	�xoB������>����)7�"h�tn���Z,]�\�]���[A&d�=�5��Uۭ����Sm�£Y�Q��!�޼��ڏ8mӪ�n�'{��⥭���'+N����)��u��n ֑�QS�}_�P2|��d������fA�v��ܹe�7 ��Z�oR5����U���sv�Gd�m�ǈLp�(ꭕ7u�)���y�(�@��wx(�O�]]-�~2�Ö]�+"�ׇh�rI�����X0���[�>�ϫU�y���B��e@ êC{���-�eQ�k+9Kx�����KE�$����G�P�{�eH��<�ר
���&�<VԮV^��"_EO���9cK`�����	w��\��x$��/6���Y�.�4{�&5��s���hQ�AV�J�bI��ov�=�� A�5K\j%X�܍!�u�]fX����Tu�T�`��u]��wM/i^��'�:g��8��crv2�8E�.��MRN��j+����d'
�oz���^䷢]%t��8_�V��M�h$�wYF��T��6p�j�g�f<+Oe:� .ٸ��^������l�c�c{b��2�u�c��abm���t�����@S��Y�h�N��凓,{���q�����CaU���ϓ_Xtƫr�*K
�9ְN�mg1Z��A*g����$�H�l�� ��`�1f��,t�ë����ɜOf\sm�rӽ
W/����}k�����+�@cJ�]1%τB��y�M�4�b�n�PrI�->�.2���NTr�o��wF����YvE��ź�XڅA�����5��v���r�un�F�o%���.�N�=z���T�g�����V4�Mt/(ڷ��e�Hҭ"o64\��[@�9�x/��P���h�;��qw�7�u'�߼���-6"�sD[۴+s+��ͼa*�4��É)�vxJ��.;���s��c��E�q'G�9��lD�[��֔q��f��}�a&�k&���F�d��ރ͒�b[����t}݋#X�#�wv�ۜ"�Wt�u�yvW������As�x�]��'��=U��Wu^�N�9E]��[��Q�1�ò���^;Î�\7+�gW�7�/t��T.��{�n_K��y�[ۼ�_F���|��!����)^wqo�}l` *q��L��"��U�������i1]R��jV)���)�±GT���#n鈖��X�UդX�"�դP`���-��,+�X��h�Z)��E(T�h_(WJ±u(�5X�YTeJ2���E�0XE��bX�5��((�c��ډmQt����0�'�!^'��N2�QETA�
�m��H���j�x�X�5�y�*��&0���[�1�~t���$���j��$�`��ذ��S�̲"9lB��5Pՠ�\��KSl��T�m��*.��QA�vk,X[)��3)Km��m`�m*y�#�7����UY"�:k4���I�[��E,?!Q�H�S �1SV�����F�U�.�pbe�'�Ĩ~���aL)"������_������l"uľH|�wݣ�r�����"9rC��Ʋ���N�(Қ�G�F_C��9)�^�D�at��������z��cg��<6`x}���K>��>�0�,�2�i�i������a�f��9�͡���&�Y�aQd�댞2���w�ٴ�~eC;�ۆ|���i?l�¯��uf�ȵ�)���@���v<qDx� i�T>����3fwS!��6~�M&'�8�'�㟾�iiY���~E�H)�8���a�,�?S�Y>eC�I�'�]2,Y���)~;�n��.l�_o�-������y�A��
#
>��<Oǽͤ��:�W�:�~C�����H,*}��6钢�@�ђz���r�>��>I|�����v�P5�}�'r�H:������xf��s9{����y��Lt����N����~O�����O~�L=aY>ey�N���=a�~��N�l���Ci��`T>#�|	n�`)t4����j�ޡ��Xu<�r+9��*��B*��#���F��i�b,����p͉�P0w���3z�%
ڨ_����2�7s�1Ƅ��7*z���+6�5oh3m�,���P%��*b����y��CkW�K�P>:,���|��C�<vʤ�<��+�L��p��MYe�}o=���r!����HVc"5Ծ���aƚ���_�3{�6$�=�тr��v�,�G��" ��L�f$=Rth��uO��%]G��4,�fqS���Q�7��k��l��5)Ť&��3�Pu,�*��WΣ#��*�{�t2k��`h�xe]5�Q��hCR3(Xс��#Nt�Y�yEJ�gwW���^����<��%����B��+���Oθ��.+�5�2��ԛ�]�n�9O������R�7+����N�ۏ���)@Qz��1��%M]����rY�I��z��&�r�3M�+L?ddT�s�@�`����3�b��ȑ
If�L�E"��c���F�y��靛��&���l�3�P�#(��E���1��A���ə"5��3;��&Q�t��y�W[;ћ�����,��$��LКJ�0�E�s&�N���Ed�j`�Y'
#6��*3g,e�qczh��e��P732a|�a7�wS;�w,&���B���߰�Oy�4���y�L�.eW�ƜɼK�DT۝VR�(�.��n:�Q�vwb�Ιc��>�WV�ㆁM���Qy9��2�.+�4@c\�E��ʩ�8F�m�7箴�`Yzb���:oc���8��F��vnl_S\�aܓ�r02�R1�:�C��:E�L��m��t��:pnP8~��[�:�}g���ڲ��8������W�����D�����<�S��g������<;=�����U� s�2�6�y�h�\o��kB��OZ�f��ua�f>�KRY�yҏ�՝t���V)K����kM�W�u�;�g�߱��U�e��ɰub�e-���ӌ��c�����R�t.�mӥ�r��m<����̩܅M	�d���V�w��=�:��ʑw	S*t���m��ڷ�d;�;�tj�  ���0Ӥ��#�n�#�O���:��B()�9�#FeWX�۫�-ZD�e��<M�^1�y8��<x����e�:F����-0K���L
�-1�:F�*����@��U'�øo�(�<��g�x;�=��
���.���
���_���q��B�z\��3[���Mp�!�G(;�[��Ͱj��iU0l��$P陯*��Fn�_N�&}S�\!���k�1�B,9ׁ]�I8b2�p_�ٲ|�W� }R,wlE�:b2aUD:P�Y�)��lA(=�()��~�������&N8���K��gk�%��]�,�;ċ@����ɯ=(�R�R�Y�����"��Z�}�X������u�{���-���D�\E���E_��1!��4��!��@�ɢ�B��Gno5�R͒l��&!n���\�W��\D���4�V�}pbF��2i3����w�՜g�纛���P���op������TF��p�̜3�p�`k�8$68Fcܽ�qc�d�xj�dt޻����`�+qP6,[X�����P�c����9$��s������*;�3箅p�.vw똷M�;1��wU�Y�0���m̜*3/�[�Y��LΫ��A*��2,穀��Tӷ8[s����D}g3�s�Z{������g��I��L���*yM{*�B�7箽�&jv��Wn�Zf��μ0R1e�Wx)Z6le��B��}}(����8���g3��Cx�ZΥ�)�ݬ����P����1Ա�*���3�ZN^%�/�9˄^[7�5�1���/�*��-�:�W�K��8�9�~s�JS(GD#�"aB�p�x"�L��'�IJ]�}���K�/ײ�s��GoK7�O������Gg��a����(b�1���m�-�J�ON�~�*����C6��y,�m�,��`��tA�^��>"��L�*���OS8�a$��r�{6+d�wD�Ryԥ{��z�F��сA�
 �;�Njs1�6�� �m芺u���b��t����聛C4��b)���G/�Q�֔�t��a���A\fC��%'硊��;����X��[���/����yT�9�jmb���fC&�y�bz/�����V����QÅ�W�=u��хz�ox����w������חTkyԩ�
����S��S���ۼ�7�%��)�*6h��Ҕ���4�,�������N���ӎi�zv��]݉�A���b��r^�t���<E���Wv6�rŤWFX$�t}��f��Kd�&w~�����5�s��r:>�ړ�	g�3�a���sȇ�Y�(�K5��%��޻UY{o��.����;cQ[�w;��o�᎘2k�^hϢ}���j�!�����Y��N':��t��$�[ﯨf߲��42搋����"�qi/ k�Z�e�.�桩U�p�#}�HÃ��r��N�vy]A�WR�lN��Z�E��\;r|��
��)jSq�V�L2����>ϔcr���i�v2�g}�R�
t,h_Vktj��y����Ns{.;N�e\;���9��!�hc�띸��0P�2�^��~�̆3ʼݚ�]�{ӄ����2�mC���3�\n�;�p$�H�^*�:��*ڷ�Oz`���#2o����@`kT�/���# r�(�K����s�Ȳ��U%�#	�o�\�Z���/u���j��Ĩ��
��I��AF�#jv���N�	�8g��k儓��5���J�ʦEv�T�K��)r�}x�*��C��x�Dֱx}ME8�ŭ�kº�{����<��UO�9�H���v�2;a�Pϳ�z_U�CL�瓐� O�������s�:r\���nեP+��Ҩ��ϡ�����7xУg�p����voҳ�*�tV)����҅�3\}�*�]� u�ZL6�\�	��zC�>5����0�Fx_��.[g.����R����dz*0����5��G;�i�0���v"��}�Í4,@��¼�{5=I��cm���}�S�����v8��QwN�MzU3	������XuG�ᒮ���8���W0\�X}غ{��5��i��a(i	���>+��+���=�Fkϑ�MX[�+29Q�x�]���a�v0��d#�"g1����]0l6gL�	e�0��B����nv�N�Ga�P�[���#��de��!��&db ����b�W▪W%y��#�p̞�ֹ��x<7`z����Z��xw-pw&���#�S2'�p��s�f<��-��t�un`�.�hr�1<�.M�͊�8l*3g2���颅��e���J&ӽ��׷��ݡ����&�e-����^���j��R{��+��8UlK�5t��s0٩�n�ήSjYnf�����G`]�����t�$fl��ۮϻ��p�t٥� +��������jJ5X���p�w��!٥�T�Z��$Rݙ��DѮ��q�7[��Eت�·Z�����m�v�l��I�t��ON���뫦\�b�X�+W�<����r�!�7�w#���)
۫Vp�K6+�� )�*��'Ej�G}�6�
���Q^�T��#M��z�N�ye�	������wԷ$�z�^v>�8?c~����q�"�R1c ;�V��ݳ�dgCnp�w)^��ݫ���C�F-*P*5{�~pmYC�:��	��X��zZ��ϯʲs���u�]�agy��=.u�{��s7�ˡ^�e]2�4d�g����lL3jx��HEd9�ON�9�����[��%��#zk�1�GhN��\��&V%�e�|"��H�q�{�%ivD�ÝmƔg՝L�r�p4��ItTi�Aӥ�2:F�ځ�n��)�[�Y=MHz�U�g�!�-h���b�p��(Ү�[ufE�N��ϙ��t�U�"����߭�Ls���ٲ��	�'¸�c%�
�9��T��X<Y{)�3&2+�K7Y��(���Q���Wu$�ʻZ_����>x��M�(Wq����LR;��V����>�a<�Z&�������Ip�H�e��@!~$ua��Ёz^\�<����c��c�lRڴ���eٮ�-�{�y�K;�Ԕ�x��,_9�Ɏw_�G�jQ#�:�l^�����Jt����o%ڣ��A���n�T��9Ȧ�|�7h�R��k����A�n���Z��T<�����{���ی���O#�|�;&(�6M{A*����+����E�Եp��d��]���՘��5�	.Ȟ<X�|�D�L���]�kU%��4���!��(�k�f�hb�}�S����Ot#c"�+��p�;��k��X�~�AU��xc�<}�,��9���Mú淐���9W4�
8y����7RVy�:;<�V�c��y�C�G�z�����i����%�z��
8�E<.&o%3F�<��^�j�甅nFΌ�K-���*���.�����J���U�U|Ò�NJ�KC���q���=�����+v[��NsU�^r��x8���j�P����:�:,J��3r)��^J���N26���ڸ�,��OeV��Ԉ[R0�4�s�&ß3>��P��{�g�ΚUC���T@g���|+����f4D��&�~�h��czY��O�c�x�8���.���!����`S+x��}��[{��߀��\��s�\�(f�5y,�m�,�,c����A��OD�"���\�q���vn�a��V��;z��aR��u-�^s5��65R�z//�V�}��c؇R�{K�&*%I�̌�L9�*'�ƙ��5+���l�3���ҺE��=ב�1�v�}"X����h	�5��B�e��۱Z�=��[w��U�-vr��#G�â�큂p�^��fV��"��PdJ�Y�#m��L3Fd�7Qڵ�������A����b�������x_�����J�"�C6g�8'v���ʸM�Kk1h�+ˆ��tE��u��%'硊��;��2)�d-��f�v��6��U���?<��/��&t֣!�A*gd��ܳ5�FhW���P��Պ|�?����cF�bw>�~�f�o���;V��׈��9��������a]���<�{�(��>[x�I4����UojR�2�u3,:d\e��F�1"$c��(���z�&��>����=�����k���s)PͰ2��r�P�6^�`��. M ���?x+V��o��֜o;����{5�G��B�
��;K4�ף#�׃ݐ��d�U�ha`�
�+�Ȏ�&%�o:�ʹ���m�ʐ�=��*M�g}.��C���s3e�C#J#+��k��M=~��#��l����#��=��M��G����W���wN�]���n�Y�v��i8@>�]��`��Y����*0���{q�+��۾3�Z�u��]���cb/���E�>����Yj:����Ѿv56!�'4��E���{[7�w�BT�M4tS�b+z�seLm�te�]ӭ�΅;�����E�Ԙ~~��w�MѾ��v�ȍ���)F������g<u��U�<�d$�H�G��Q�mɼŝӝ��������(�K���,‎���F�K��mθ���Jd�<Χ��WwiFwf*r���R��Hgj�h+/�
�߲Wc�)F�#~S���R��b>T������!k�O<�AV.z*Q��%h�/G�|�l/6B��跴t�ؘ5�&V꽲�gOu���B�3�~����p4a��_�H�:���-����9���7Kb���8b{۷a�����q�m��{E:_u����^ӄ�>8�\�´�RCh�"�-wgv[]`��~�;�b:Y�
QEߩ�"	�*���Hj�*�c�\3�)��$T�X����(�Ɩ3'�p�n1!4X7���R�Ҫ��c�FG.˞U�kp5=ҫ7��cj��I+C�^��j��Y�!�'����3�bd6z���3QS��&_�}C�'�w/����c�N��rl��L��d���P�>��
<��_�P��^�Wm��'kҭ\�y����Am��sm`/Z4cX�p�GH�hbԏ����,[��X��4k����'��-�u�l�5�.���:e1r-�}G�#}�	fCF�nRkr�sa��9�of�]�z�vd��<��dܴ�����^�YY䝃y�tsV�9��
�r�+��/^�`�����1�$țʮ�8��&G�(��&��,J�G���0d9��#����]E�� �У%f1٪r:��׵M>[�;x��*Zs���LX�A�YY8���:�p�{���j�1g�'�3ڦm��[��*�)��5��c�oP�6�=����u���y�w�ZP9��I��Q�0U����f8M�u�W�ka]Jv�eK|��*|�s� o��$�j�m�����q�]l���G�S�jQ�|4�M�%y�gL��m�;�����[ۂ4��ǣ5b��I�.�����nw<�q��p$���l/+\he�ꥊZ��*7b�eG<Yz�����-S�Ȣ����\V�nLD�c7Gs�R��bV		�|�D5��#�u���װ�g����)���۹}o��:WNu�b�'R%e�T�+}q��f�Ge��m]����wE�%h1��aX�q&���.V�4vZ!�X��I��2�'h��61]u#䗥��nE]l�&,�/<��u�_@��2dMRy�!�̑��,3��d��C���e�ܩN�$dӶ�Hެ'���e�m�Լ��5p��!��ο%��H��]N�}���J�w�������zJx�A���ɦ�W�1Kͷ2P�5�n��\��ܕNu�N�덇���h�`�Co
s2��d���Vomr�ʃ�x@�k�h�k��X��uyV+�)O��Y5{wQw7�p�J�����ᔖoJ�V���{cgMU����nf��h�NŪ3�Y���͹��֩ch��ymJ��u�� ���:��q��?>k��fwu�*�� �Qz)k������_0�}�>�S�w̺���M%�Z��H����g�)��S�O^,ݣ`ы��뫩��x�k�䩞t�w���]`�/2�G*»� iTaU��.�#8�e.���:����b|��uq����M�x��� �n��
"�ӻ�L9t�o�*�d�Մ7wI�0��Y��7ٸq(j.`�%Q�m��Ɗ)\>�k�׋k���*��u��nu�g+�Z���{n�w���:U��T�&�rήnr���9�5�[5�6�f+���D���ñ�a�f�+'	.ɖ��ɃNPt��"�O�^���{�1Pm��<[��-�X�z�� t{����=ĉZ�P�����Flk/��sl�7c�-����&�)=*��1d.�ڶ�'�|�yz��"�ﶮ�jG#�f�.cXL%�N���[u���<�gc5���jI%LD�QD
$�P�"L̢����\�4�H�Җ�fYDv�ңY����EY��S��(�0UbͥaX�V��ADV˻UA�U4�e.R�J,\J��kJ9]f(-J�J�c��L���5V̸̈�Q��ʬATV&�A.S�m�QLB���
Ud1U�+����\Ɋ9eMsY��!�����L��b8�[D\M97ab
�E�f;J$ZѬ4�V�!��8�.\�UX��;��)�TAjV�V���UDUb)Y�f��QX��Tdb�������[`���3l��?Rň!�TW�U�Eq,\�X+#MR� ����b�+��Q�o��X��yl�MZ��
[DEJ�?P�)bb*)��Z�,PTc�(�Q�Ң
�6�~��a�{8_����Ȫ[��q���Oj�xї��
�XP�ԩȜ�I�E[�a��j�i�T7�{�H�I)�=�t����������Z����Zڂ����.ߧ�i��\��o�Ǧ}0�+:��gum�<�Q��Ȼ���`��ȹ4Y�P���aQ�9�-�{zh�|8�d�����ZZ��Ł�,ϗJ����7\{"�O�{&�*��&�Y͹uq ܻj(dHu@�,ʹ+�H���p,oJ)�������G`]���N��t�'��W[e��g�_H}:��v��cg
�ͱ�)q��+�R<���۞-�;Y嗦1u�� ��gw����N�c��/խ��p�`O��#C��#\��* _B������v�l��Kk�����2úf'�矜VP�/�*|��T4z��u�8Ծ�ʫ�^1s�iX���É[X�}2�R�e��˦x�]WY�R�d��Q%:��3�
�Ւ{��Ռ9���Z��~P7��z��~��g���Y3㋰�K��Z<����(w�%ԡj��l��c��#J5�,��3a���%�ʍ0�Xb���N��a��*T�98]�-g��U���X�>�w�:��^
�[sm10��3�tÛ/��)�@�%���>8n�Ԟj�d���=���]\Ak,�&�f��ׅVv_l�L�r�j�υ����IO����H���+�;˶����V$�U�g9H�&B��R���!F�t��q��Y�t��g��b���,{�U�TCu�������l�����*:Fm�T�Jh�l�ؑ� ����!���0�^�e�ܬ�3�`��X)�-
_�$��:'��[��D:!�4"X�]�\�|gV�E)�*�0��"��(�Tj��t����əF���)�L�$��5
)�.���\�.��fV/�4�#Q��5rLhN|Ur�k�	X��R�Y���b�����u�s���ⶮ_s��]Q��q�\���r%,���]�&�7�b�sdW���z�:"�ܩ3X����5pBu���(d	<{"�W���C������Ey��֯B,c�r�ΏE=������Lው�/�ލ����\��-�dů�t�8��ZE���'^,��Ug9���؆On��n*Mb.��.8�EƊ$��b�ҧܦ���ՍƳnf��^%-�
knK�^ٷw���VÒ����KC�UJj��}o������qyx�N�',p�^��PB��ö���mK���dۦUz��s�P��B�PZ�u��W44��e�ëc����Eb7[�Uꫭ.��M�l�z�����AH���a	��v��Ssqv��zV������+�}�l�^�.���K�ሥɽ��wl��n눾r�K!���P�J)dk�t^v�0Q���{< �X�r/fD�=�z-Y��!�n��#ElqH���Ü�Q.<��U(E��2�p�\�;�p^J�*��
�L��������#"8^�<�zF7������!�ē1��I��u��Js��F�ʉ�D:�%O[��>��GE�Y�7Բ+!��_>�B�����	�ӛτ<5��2_�2�3�#L��"�5�,�Y*a�!��W�1�| �@RI;��}}Oo�E���Ag<���PJ���tՋ�h^�Ҭ���3��RI��TCZ�G*��z,�����_K="û���x�����1R��v%
�C�6{��~|�,�ϱ�ĻDiy���"e�]�C&��@Ͻ�s	���#1^�e9��Q��g����Q<uh�hgŃ�q�C2b���I��`�	d
�Fp�Rv��=��4KȽ�`y]%����C�c�%�E���l�T� ����2k�яA�ð�3V�a��C8�A<S�3��n��Ї��jh��Ck�%�-y�ˠ�6=�c<�=�p�{��&��`D���n:5�V
�ϕ�aK聚N㏍[�r���z\:��K�B��Y���	Vt�Ǖ��o{���	,]?���y�O�fonDq��J�\W��ٷ�!�sHE�dat!��T��4��WrgiJ^޼����U�8X�$��S�Fs`�Ѽ�70����6U�ha:�ӝ$�������e�r��/��Ʈ������Z��Vם��zYz%[]B��|���m��w��T�i��;�PG�l͖�):UCA�{vf��t�}^��q���m��J����K������W���HƂ��,�E�O���hj�q��>�F�̊�⒩"���Z!\뭄�]yVb92_�ٿ}���Дc(��R�XR�r���7��6�VE�Mc�ժ�l������d\�C
]&��v��D.04djo!w���z��}P9>ݮ��N�ó�&�N��<<�CO-]\2Q���K��.[!�y_{6�%���A\���RSSË���Z�������L8�`lR>u"�`~-r�9�o=���u��3b_=[͍Rwa�>�+�l��u��Cp�p|Ez@Xgb)Ծ����LV��v-�AaP%R\�V��jG�� x{��a�}�H��Ƨx͝su��*��bz�r���[��(hݗ��f�V���aP:���K�맇^�ŝ�n�Y���^�.��b�6�ݨwW|��Y�Ѣ�ߗ%�7бj�RK�_xx=��n�P�_z�ء.sb�
Y�R�,ۄD2��Lą�j8���1lMb��7�"��G6�-+�\*p���!�,��5-Ť&���>��Y�UQP�l�`J�.�6�2c��a�Ҙ컯d]Pg1��ș��ר,#��`�cņ)
��䡳Yi��6�����#t���5�lv��;62��E��!��3>�(A�Ă��Yzf��9���+�)N�7���D�%d�����di�&t�g��;уrQ���͌�#���5f��'jU�kn�nI�������~�A]�"23b�18FTf�^]7�n8�E��}�-��U'��N5��3�TD��{uǲ)@}�b���wŜۚ��X�����f�������Dg����q��NG:&�]��PLu�d��ݶ�O[�ߦK�_�C� es�ؗy�w3�Sj�ۋv��B�\E{#TW*�ls�#M��#`=u�je�<`�;����ئ2��6���ca:l*�E�'M��"�R1�η��kܭ�7��;�lR,/(�4�ei�=����rѶJE0�p�wz::YJ`z�-nn#�;x�F��ii"9	�7b�d76|
�d h��}ʋ�q>��J�ݭh��;2�'(y��6�O���o3SN5��Y�N�yw�6\��;S��{�K�֯�U��n>*�&ºF)E-��Vxg�J;@\�ƔtF>�dmb�����.��r�t����}�l,%�b��ˡB�@�B�����4[K����
�L�bup�|/4-�ivEɬ���03e����
�2,bx�c�Na�(r"�edocEV\��7���tX��"�9�4߆9g.4� Vu2�#fmϸ��	x9hv(R�����|/�q�r=�=��*���R�z�^�J�"��5�Uø�挎��xE��/�ג#.����SB��7�є�p�E��R�l���*���C�B7��R���D�c�4�=���$eN~UQP�Di*]pWrN����߂�N��>u��0n��.SуN��a�׳[Y�e-W�CL�b-9b)לD�F��&l���6fQ���vɽ�I�W.:uó�ዟb����2�g��f-����'�r :�D�l؄'בn��qU!l���fm텙�ԇ#x_������Ɗ�JYqќȫ��˂( ��I+>H��?Avp
�*M�8�,.�{�*n�wz���XR<~k�ǩ;W��!@3�h�����b�y�l���W��r��I�*u�y�aj�ǎ^lJ�f.�P���=��U���#���kэM�-(wX�;s�Zn<�%�\���Yõ,۞_��.��UP���NlӢE剢�0�(4�F�8hR�&���"�o+V�#���%���^���2Xl�#b#ٱ�����B����uB�](�7宴��5����m!�婼G]�::�p�|�L���-|9�qy�肴8x ���2�`�ٵD��s���U�����'��![���^ٰ�4�8hc3�yJѳybx׭�/���.�=u��\�[S�\�T3��WL���z�w`Xv�EJQkcH��Īb�X�#�/:we�(C�%a�j�F�!�qnQ�r�Yy(��� �#TM�>d�2�`uD�{�,�8]s�9i|z����>�UAX��^�,��Q���s��0�z��ՒǞ�4u�k{
�ux���!Xs���P����^�U�.T�����m#W�e��q]ڢ�z�$��N��l��@Ɇ�4�������#��p�}RΉ�׳ba��ȘF�ή�:�h�UΒ��W�[�F'ADPpAea��˥^�~p�B��4/L�[#��A��I�.'#bb�������D��.����ús����q���9���h�Wp�u��'�]����sŽΣL]r֨w�9<��^���T��\r��͏��k\�8�ۣz�WLΫ��<����1{4�[ð��h|py���E1N]i��ּ �G�k���x���5�N����K�vG;�AL̇�RN�LӮ4E�*�~"�9\K�꧇j��ک�珧�z&)���kܧ��dWq��JY�1�ׂu�'��#1^�D��7{`����UZ[>����ǍɊ��4T�h��y�8f�eNT�8J����zq8b;26p�vl��&�3�w-ƟA� F9`�⋈\c�\Lu��S�ڍ��&Iv==�	f�-��r�7:�m��!�.i�dae����	�;�D�j
�neN�<�+gs�!��b�q ���A|�ԳN�td`F�)����v��w��^��̶sכyܛz%K��|�C���qnW��y��ޱVs���r�ǢU���v��?���X�\�1��J��^R=�4��okۉM��Y������Y�T�Vy���nx+�P��f�R�΁c��`�9e�_���9HF�M����2θ݊���!%rF;�����[a�U�.w��(��Գ�b}.@�S�b�r�R�R8�~�u�ۮqGh�3����Vљ	�����"]��A���f�vC, �iu�h�4|�Ы��do�s�s���x��G-X/4xS�=�ƨ�d���N�/7r2�`q�pQ����Qt�"h���w��]C%�3]�%چ�`�9��3)�K��-�|����ﵨ��7��ԖGC��ꐎ��������NUp�AF�#ux���wa�q<�]5���dYm	���w�P�\�|0�H���K���?tIn�;����ע�r���ѿt{^�A9�Z���~��&k��a����]�F��q����A���5[�X�#f�_�Q�]>W��.tԈA�F(>"����9��� ��.
Іƞ�ķ��nrxV ��8��ob�NlX�)El8DA3*���HZ���{z ٗ�VK֫s#�t�$\�R�;�� �3C2C4YôKq~HM��>�R̹��;������5�BË�*-t�:=V��;H����W�5�R���Q,�\�E�Ү�|�T���vf����"�=A;2���䏆)n����7�y�.��q��Y�C�,z=�8xpe�."���D�'d��^@f�:L�.��]����7��[(x5ʶʽ8�^�������?wI0er4&���}U3����	a�!����,�6q���W=�:{DDN�#���d����R�Y U��z�8|�Օyk�|;�X�$�\ë�ffK��)Z�ϮqI��O.႘�Ԯ}�F�_�%>]��
���������&9� _Z{R��sʮ�rY�I}�N�^ �[	J>Jh�{8Q���3�TD�YOa�n��E( �=�l��*g�t�<�=���eף�b�^��\gBz��V�%q��c{���S�S=��'��݋���EZ��v�#��ЁY����*�ls�#KnB$v�6b���Vru���o/LSN����N�DP��tԞ��:	Y��e�2	��Y�ok�:X�vӜ�wh��F8�&�H��5)E-��Yញ(�r�=@�w
��`B������,�鵣��>ϻ�5�K�5��6eШS��9gJ˪GyWS�a�V&��T�@������͔k����@ކE�bx�?*����Qu�V�%zb!?u,�������B��\��
�#N�R�X�(�gS/)�6eǸ�i�[���t��Ȏ���h]NT#��V���b�:��ۖr�^�J�#\3�F�p�2۫2�w�{�j���<U��`�Pl�kg&1Ӧz��l�k�PVK�Fh�n*US�^�bum�� ޭܞ�v��&��0��P�ʨ�����i����� Ɨ��g�����`M��rwued=z��ќ+l-��Y�\��	�
��Am)���9�+���\�!Y�i�{��B�j�[ܨ,�aV�"��zV�?5��{�p���X~E�|2Ӄi5'�8�e&��5d��Z��\��#�{���oXԇ+��Pzs�E�����s&R�wo{7������1C�R�hL�:�i�!)�n�H2��VA�a��/FN	>��W�]RQ 8T��۝!d�eυ{ڕ�GL{�V2�Lk��ME�Y
��-y�Q�J��`�6�Ǆ�X�h<�p5:��\�#��P�.7���fR��Dݤ!�w�;o]�42��V��+��+�F�Yl䛽�� ����-�o�%w���|e�!ͦ�%���1f7j�&��؁�N�������0^Fz�)Hnv�S!v�r���W�.�7�A�Z���^W��[�����9m	���\Ǿ�Hs r���s��n^^�L���_;��B�±�䓺��p���(+kz���u���fA&�1\E9�h��y���jP�_R�gu=� �8ۭ��U���j�[D>&ue%MR�����n��^N��L�e�+n�<H�|������Sl!��F���L�?��\+�`R��U�ۂ�f�.��di_U���s������i����I�1�ܙ%��oznVp"c0�MP�v�[U�P�$2����]wLR���z�_w[m�����ڊ����I��)�GW��U�B���wY� 4�}k����n��ͷJ�z��ld9���i��w5���5�tcf����S�横�V�Ӕ�u}��o��_}�fsy��gM�<���_�W�6���X�;{�溋2���@�o�ݬ��w8figa��+|�G���7w�-��gM� ���yz��2��MX-۱��V�aWi|�ʡye��̡L:k2��J�$w�kvo��e롡�/v\�����9�VE��R�K ,I� eL0#�/w���c�d+�ގQ�l��%JU��L�JI�:�icOH�洮u�f�Xuu�o�=��W!w7{x��*\uf^P�d�K���$�ܾ�"��c��V��a��0ª+���Dec�ӛvmR�2���ن�1[��지��[�']1ĳ*��=>[��fv�y
m4�+�g@��=4��{}FJQ��K���i���a-Nf��#�]�mA�b�|luv��U�T=�ͳzզ�婓.LU�Xm�iǽa;���rł�}��m�P���Ǐ^��娱A���ywV��PN�M�h��F�N������R�W�H��!D���#{$�\Z�7���8í�X�7���Dl���W�V��N��-΢���(�Goϭ�n���$��"�}SC�}�{���k��ds1U5)�̹���5�R�D�6�E����:d+8�f8�3v_wx�1*���*֠�?���:�PPF��k,�T�0uj�T@Qb*-�%��j��-F�"���R҃�QX:�X�AX��"��H���tʬ�UFEA�*��Dx�+啂�����X�lE�%�iī�*�b��b,`���&Z"�x�UDX�b�j*e��#Ti�1��b��6�WV����DQ�1��UQ2��b��Q�5�PUQb�?S2�DE",-*i���Q]�J���b<j�+��VX�@ݤX�`�EUY*U�UDSi���1��q̲8��V���EH �YaXr�X���b0R�`�S�R�,Q7J��A�#�1����Ő6TV��"EL��ٸ�l�*�d�,�v��S���):��]�)�jjn���[-��yٽ�ܷ:cW��3q[�)mb8Gl��W��"���X)5�]�$�˵�߂�O�6O�Ŵ�,Tǽ��q!e���^X����CQ��[r4�S�8*���'ڂ��x���
]���)��s�s�}�b�c=Z�A^�!Y�{B�=Ȍ@���땓^zQx�Q�_K8�E�:Cjڈj����c.�U���F7�����3�rO��\E���E[Uʂs��SX���Wdr߱
���xF\�	�&�(� �lӍ��R�&�W��V���ۥ�������G�a�x�=�C����K�|�f�v��搁@�hE���z�Dq䦨#�v3H��igV$U�e���i~n��y�-|9�qy��
�� )k�"�Ғ�7�\��y1��խ���h5}cz�(=u�
�	�41�����Y��%�>ʨx���{7��|��T�-Ɩ�ړ���+"�(�d`��;�)	EvBu"��R@�mb�CM^FT��b�c��DM��<��R��x��*��^��j��?x#��QYݗ���p =ss�2vP��mږ#�?{�񋟎"W�hڛ�a��7S6�`2E�c�����0UӄTX�R��Gy��;�%�O?t������m+�Yy�%؜�)�,�=L��bz��r�����B="r:�Z�㼳2�~���;��m�}�t�lՏ�m�E��*q�]1t�.h�%s�Nw����6�f9"Y���e�+T%Ė6Uv��G�e�z�t��=ns\�+6��y!�`-z�v��n�v3y;V[���{��1Q� ���9e�`�(���6&^��"�wW�Tڭ�S���1���B]�}��nEtE8 �+�E]*�p�b���*0S��t�؊�X�-.�����l8��J���r�H�w�+��q	ϓ���%�	�_��y�x���<�\w2X}1���\iQ2Ƞ;��M����fkʌ׹�V���3�3�ffԾTu!g����צ�Q�p�,�d�Ecu&�T�R0�ќ3��&�D�n���s������&O#1ň��8h��^����]�q�A�����z�-A�� �J����K��<=�P�� ��5�:&��D����?�-1^q>�,���5mb�YWv[Q��;�n� K�j�C6l���I���-�W�R�;�c*5�[���7_�YC�o������c#&�������4v���j���/��p����jJl���ԎR��F`����K���%�2��U`nDdޱJ�]6*�����-C{,s�'ALZZ���_X$�?�$dP�W�nL��4MX���a�ӭ[�|�%|�u|������՛�4��4��SC�c���9�x�T���{KBp5�r�z�Ǣ��G���7ݬ$g�c:Y�di�\���Gz�5�7�g����)^�`�'�Wf䙰�n�;��$��V$s2�43�{���#Z��ny�}���V�j�<�7n�.Q4���9kDX�wr+�����zq��2��8�׬�ALN��=ܼSֽٹ7�b�θXcG��48T�ΰ	��p�R'[���v��B*��!��dJۛ�H%�MNB,=A��'M�p��d�\}(�႑:�ѫ�����T�^�Wf��ZV�����ɭb|Oc����|tY�_���l��qc�^�ȧfƞ���/WS��*�&��u�_�/�:�r"�ܣ^����9�ё+%�~�Ozn�뱒���H�'�eFϮ7�AFlP吺$���(�&�S1I���(�}�$;RU��ɛȄ`7R62n�Q��t�\��dtp�n1!4X,���!�IȋN��.њ�f�=��g�׀4���L,Ȫ��BZ��^r7Н%*띲·a��ػ6��؍���Ǘ�I�;y֙�*w��<]�w^I�6�_�J�C�5z���O���))څf�$�ي)� ��bY.���>Um%V��Y�;�*�]�������rn�W�Ϊ*1t�:6�y�;u#���I\�*��͖�U�^��e���0k��U��n�)N���阡(�%L�׺L�An{#j��2��o.�`��]�M�w>}�(.XR��fP��v�
(��jc"b�vL�k���JL��N�ތrQ�M9�O
%�����y�e��~��}[�LS4&�Tً(��f�L�%���,�ءN��%7Tv�V�fe�fT���F�='_��Qczh�~���Q�
J�c���q�Un��5�f��r��ŵ��\� I`�޹��"�W2���K�tM���Ơ��h��p7m�5kR�3i>�팞��*8����U�U�Ui�s����B{!Y���;�p�5��*j���Fmnr�]�)��[n��c��_{�4!c9��D;�Қ��a�s�5��qf��y�y^�݄WWR* ^���&úFJQKc:��(��EU�S夀�����xҳ�����.Y�.5��UŌS���$a���#:f�.�z�@��ѣ=.��r����0}������7m�8��n.��[�`Kt�8��5��T�#�}	'���s�|EZ�WZV����F�C	�r�&���`�����S{�i�KZ�6/�xw�E�l<^�P�R�۬n�Te��ur������"Մ������zpIY�y,ؤ� 
�j)�FX�Wi�`"'��PW3e���Z����'�W���PN�j�3v*Ϟd�i��ُ|�������)yAL��4�)g�tVu2��4g���G\g�A���jM	�)q�e��G.Vޙ�׬]B�m�9P/b�N@k�QҪ�ٝ��v^�v��}n��J�2��4Ux_XXK�>x�]??�,|�E]�/`T9�&����녛��T��v�0��@�,���3J�*�YDԺЮ�I��kC�������j���+{��#�t�(P�wlE��`%�y��W0߄�AAN��tV$�@��h����1���R=��&L��3��3��S1a���b��D�ȁ�)WQJ�������v`���'�aQ�=y9p�N�=�B`�9%*e��^$4׻E�wpN-��F��:�qt��EB���$^_��n(�%Y�X�9�R�%����ɭ���N�E{�vw�=slk��� 絠��xc�	�lm�t �\�(-����uB���ef�8[]]�X/�zj���}z���AB�yr�V2��;�;�q켵kvA�P������<_���+>�kN�+��0aUk	�]u��A�܆��u1��K6{N���[w���,�7���n���YVӕ3�~�/5.N�n�^�F��n��v���'Zd��;�ER5b]q�ƈ㾸D��L�ze)����k�hO�B:��+����*r���ͫ�0h'0pױ��͋0��܊s��ǎ�#�ɺ��@bܳѓ��8���WL��/T����Q�]�v#H]+�e��9c��К�R.����8��>DP�(�9D,�<�K���#TM�>gk6����p�m���޹�muW���ѵ�Xm��=�b�p��*�Q�s���,�{9f5�$�.����9Ȋ�Q�Z ��`7G�q?���꨹l������c��tGd1dL���8N^��IMHG������`�1��-2��ȱ�H���(���70:�tVȷ�SۗP�|�)Z�ܓ��8��VcȧLn���8 ����`�U�6tՋ�m*܎�u7�e�1��z
�L���>͂�3�$�،�,�w~�����Nt1Qw��0QK7���٬|�	��2!�s��2/��C&��vLXw,�Fk����.c�rB!z���#�9V�X.l�92�2Jky���oS:s�)��m�#n{��2�B�N����H4q�ce�d0w���M>O� �=N�}?��L��H'�~�`���U'M�����˧��j ��d9s:yM=���[���WQ[��1�����N͊��VJ8�5�1Q^��M�`ג2�3�b�:�'SYG��[��m��G��K�R����͑%����\eܷ��1�H��:`ɽ���H�⦧[��)NḎF=�܀+��>�C��.��O���n
f��C"˖ʝ���4yҭ+[���؁5�[��8Ç�rLQ3�|}K4��]F�(/a�P	���������@�X6z���яhW/��<{*p��O��T���3R��k�1y�8�l���A�+TD�Sl��diF�Ua�r��iW������0\l�P�1��=�>Iwj�S�Z`�
�T��b��)��'"N9���_:�vN���W��݊YE���W��{L�Y����L5��l:.J_-<M<դ��x#�eu�/�����>��rȣO|��G�W�\�E�JS%��P�m�Gh^U�Ȫ��Q�+>�I���W}��o�֯�/0��:�;A�b,��w�J:Uq���Gl1�O-q2P޺P�G%LU	�1b��r�nS� �ִd�)��O/�eb���l��T��,r�AЋ!�M��Ę���X&�/H�s)Ö���6�.�K.I�Ie#���mSͮAi�n�.�|�	p�n�<P����� �xTٱ�����M�0��U��:���dzh{A�nydֱ>&ߠj	��hÎ96)Z�&*;�/���gu������^[g-/Y�ھ_tΞ-�芍����W���Ed�fsB׆��q�Xa��F�K�)_�
��7�qB�D�v�� ���f:z�t��]��C�S�-��y����6�>^;~�t�z��k2C48v�j[�		��mk:��p첡Wen�5Og�>z���ϥo3gE�.G6G��RJ�~�g�f�O���ύ��wԼA��ޜ��-Vx���Zft�T��QC7�f�s��t���+�^]2�(v��8&R)���I�(A�7xP�ŗ@51�1^Nɂ@g:L�4��y.�͌U⬺�]��k-�Uԇ#[����0���&�f�ׂTـ���_D���^,��nҋ�b����.C0T�*�������������S�[�<���q]�Wi[�%��"px��������B�&�G6���W��P4.1���	�a����YH�t��Z�N�N퍋UzfB!`q�9�|�jp.�vK�x��F�V$��=��,
��7���յ%�x�T(��X5wm9�ŉ�1��_XZν3��L��:��13�ۛB���(�,��n;j�f@��Y�^�|WiQ�� ��u�::�N����Z=Nbʮ��V���d(�D�+�¸�]�*�P�-fp%����媔��^IXMPf��Zv�,�1A7rt���GJ�Dm�ݻ߯�b��!
�^B��SJy�gdt�����N��Ft6��S�
�������G* �9�TS�(��uB^\�o�e\u�%�qx���z����X��3i�@�����+�D�|����.<͙�R������oDF�)NZ'�B+#6�{\E�z5��1��_N�鈟LD��}������?�q�2Ή�l��<F����ҍgK.\�:gj����+t$�l��!���]<��֯.�sR�%5]qd��jak��u�Y��[�:�1A��St�V�Q�ګ2%�0Y�؊�U���3ׂl�k�PW연J�wJ��	��<�^�O�5[�-)����ؐ�Y�3�d;��xUz��K)pC�Þ;��Q̽:�WOt����ml�:L1"��e���i�s��Q�f�L�n8��M�>�t_�W��G%h��u�u��Qt�_���ں p5w4Mg:�t�0�z�Qu�GyH�t��˨�|�2�z�r�I)�`�Z��o�t��-o;�����uvY�#+$����@nV�O����v���1,�ږ(��U��Sje�r�4g畧6��L�"��I��S1~j`오��+�^����O��$U�}��"����������z{Ԉ_o�!*e�[Fs"��%Ef��O(4�������:͐xG\��"���n�C�;3��z����U�Q$�?-�KI�K5=�+go�BW6n��pcWT�8���b#ٱ��A�4�
8Z�"��ޓ�x�|_���uN�;����WK+�� ��Z�s�ϖ�41X6 J����.;2嶱Z��������Ս�![���^ٿ+�0S�6m�ꌾ�=�{�
�W���,.#8�܁6�2����E�+�E�r�Ny�gv�"!(�țj���yL\�{Zw�P���AӴ�P�vܸ��)�"�J7c�#^+c���8��#TH�F���Q���\���\7R�_L��#%HӕU�zW�f3J&/��&����_"AqT5��O�C��ڛ,>�Sڂ:�����y�0����h�=U)r��?J��t��	��@`ʼ�`PU�4�j�;`|�UEς�n���ی�1��b�dY�nW[J�*��"�88�|��
�;d.=�ꖪ�gX���=����5*�sx���'Mh�Xڵ��6����v�|em'���$kVƷA1���B��
��#���n2-��a]�k�mq��*\v5��C%GGZFRDQdn��B�->mH�6���7A�ʲ,*T쥆���27�M�FQ���*�(Zlg���'+|[;�0�-�ڳ/��4���ks/�4�O*fV��s�����֫���]m�ٺ��y��v�l����twF��9�yR�/��)Էw[�\�U�c5�)N�����S��s:�T"�"��!�;�3e�m.Y�I���I����S!5ϝ��R{�>�;)�{�e��\'�J��A��p��&���k
ޣق�XXle��	�:���T ���H
��'�WK��P=]����E�N+������գ;8���B)*����;1���ג�JwR�>C F����	9��_\�T���t^�:h-9P��d�[�G�d�Jc|��x=�Ľ�km��֩Ò.��Kٓ V�y�V{��`����Lzg�.ZEYN���;����mf�[ Ʃ�[A�j�%J1���c��``�2�5�&��x<�VGN�r��v(�][�Ū��xf����^^�� zC��8�̰[;�9м��.M11t��;���h�%��iO_��(��%��G�T�v���m�8�&z�t�uܳ�q�]~�Ӎ��/�ffs�RQ�J ;m'��KT�Ν���:v��R��;��1�uЪ75��>�DD'OtP��T�oM�W/��f�)V�1s��f8�a��5wQRɭ�]�L�V7��:sf�&2 U7
��h�ɹ��\÷�J�Y嗓q�VM��(�@�i�Jt��z��ɶ��^��E�<������=��%iPu���ݒHM5�@cX��cd�k�rQ`�Wε���K%�5��E�*���<��"��3aC�Ʈf/�7v�{b���#a'7�ͥp�i9�/�M����)��q��a32�K�ƣ������NȽ&:�m���T��0�GU��u�3ol�m*]q]�g|ʇ�Q`ώd܆�g�������u�Vֻuqs�����׸Ө�@��4�o$�]��������A�O�w˷����[������U@��d�:���fJ�o�ۂ� bK:�Z3�w�۸ $d�QcW�*O�u��5��JQeT�Mt�ݛ	
��^:W��bW�[��n��7wN��<j�K&�����<����Ҝ�s�H��̬ΊPg�j���F����)R�d]�'j�v��h"�)�z��7�9޳�9v�!ۃw�̲���l� �ܚy�Wٯ�;�N+;�w����=��)�1X�Җ2*�{LEY�-��"���EX���m��
��Y
:�dX�R�T�(��D(QX�.2VV��b�mA`�l�4°R
E�a�"�SH(5-����H�
��X,QE�1�E_YMY8ȸ��9j[e�b,���J�(赋a�R�J��J�1D-ĕ�� ����(���b�P�m���3iY�Fˈb,2�q
�`�(��3�1�Sb�J�Ū�ݡEj?�UTQI1�ª���R�(��ee�`���P��� �v�(�kQR�+Q����u��:paFJ$FEU��`�s11
ł��C�E_-��U��*,�+�R�咼J0RAU�.����$�)��Y�P��C_:
�ތ͝�:���w��+01��}�R를Z =�;�[|�Ρ��*����x`]ܓ��mE��]#�)���B(��Zd	p����R���6?(v��FZ���g_m�.�r����Y�#mȣ��� ��,3�*}e��Z A�Z��=��^�xz��,4e~�[~��lT9f�J����U�+ɚ��I;Q��j.��ոu��[[�W"f��"��1��b�|�he/
{�W�u��1=�й�g�n+q�a��k͹�RH�ӓ��u麔p!�kٓ�n���$e�.�ΰ���w.�J��9fa�3J����tC�[x�1�i�u�}P܋�9���F�P��/�{!E��g�-m�DԷ\E ��A�rLKU��I��~Re`j���k6�n���23�\ұ�(.�)�R���8B�QRt��f��$�UWȂo��0��iۮ����U:+�谆n�ɏ���{�\l�����|pdk�����ih9�V��\��eW�8y�s1ɋ�<�d��z&�e�aҎ��c^R<t���׷fls�a:�㱟g��vn�]�׊tw�gضwhÏ�߼�g/ ;�{�>��!�γ����rr�4; �r*|z	k[�it����p�w�h��(�t�I��v����.�CO�mwX���6��f���	h�TlVi�v��.�!Tks�.�&5.���r�]ϡ絽ֲmw� '�fo6b2��?y��s�ȣK0P�̤t"�8oO�@G����1�BE'VGJ=}3��Ș0o���iԛ��q�������
�T�/���#1� �q���O:�9��Tlچn��`�,��J#:U&��#�w4:�����9I=ݓ<&{��YS��FvTY�au�(Ѝ�;A�����3b`����㰎l
��h2Qn��ޥ�+��=*�ly_f�F��l7<�k�^&F?H�L��7w��n��,���oV%|ùh~'�Ø�Y����L��-�芏�#��W�N�d���9�38mD?5zp��x�uPׂx��J5�0����r�J$���� �M(����e:{ϡBkz0}��;�k~��i���J���\��fHd3�D�p��3Ҫ��7�s��R��Î:}N��*��\�!ѵkϑ���ܒ�:�\�-+�vK��I=��s��g N�L��Xt�<)rDW��U�>��;�>�-WU�^������i9���i��Ҥo*����L��%��
kyt�d�U�ٔ�^�-<�;�T��a�����˶��u������]u�X�^;9w�'�/߻S.�e�b�:o�}����8��U}���w�>��ݣ�xt�23�3��\CQ�`ϋ���24ה��/���7�\�p\���x}�\�/�G8&�f��-��Q����%%g.��<ǁ��<K��V�������[��z�
��$kx�:��Z~�}�\Ju�����=e��C��-�3=��=��E���M�6����̠h\c��zQNf�tF����2��N�kx#s9O_n ���zl�}�w�d�>S�^�9�Uy]
��4���ĺ��J
�H^wu��=���?�l���݈�7���s�)]a�j��{h�R�H���w��4[Ą�y��[.�|�é�Z�zx�
<����r�l�
dgCmX��z>��}����8e�d<�՚V�覸)C���R�*�h�E\^9�-��Q/`k/�{ɗB�)���p.�
�5�[�`Vi�,�W[�9��R6&j8��!�^͔h[��-@ކoX�0V�C�����m8,mj��~�=GI���8���7�R�Z+���p��޿h[V���޵x.�~�|�R
tۢ�<�P�WQJ70���|�k#WY�һ8�] �|�	�b���]:�#�};t�t`�Dَ�]�����+*p���JdĜð:���Ru�Ecyfz۽ijZ�U6���{�[�ʜ�`}?���)�ε�gMѳ?>�$v�%W�ʍ0(:t��D{(T�޹�r�
�{*p��������Ư�o��8G�7S�p*�ρt|*�u�����#����
���ʂ|�R��\��ƈ8�n�����fߍRp�,�Ȑ��3AUEB6#H�s�o.���ЈvY�����{`lv����x`tW���-����"�y�J�T���͑���3�a�|�Ov�����t8*$�@�Z=W���$ɜr ϲ%��o��;&+�9������k}�0����):�ɖ����6t8c=�ס���"��T{���l��7鶣ν]4��]��uA���W��"�1=�!x&�q�A@٧5�´�;yI��h��;��]-:�!;�7X\�]rd�L�q��Þh�u�4ŏu�털�ܪn8r���8��T.�R��ak�"��^
R���=����s�ϖ��D�>>}#bn��c�X��ł4�(�/��
B�7箽�`+�0h�
��B'qv4Y�Ԧ��'��smf�j�:���[Eė!�Y��u�ܳ*9pH�X�#ډ fy�/�|�:l���'�����)LJܹt+$XKj=�j��њe�R��:�u�xO^j��S9Z���m��k�!�Q&�.��ĮڮL:ʙ]�s�)Q�&s����O�9�mw-�G�;�Z�&�QQc+K������r�N8���j�>��=��Ǜ�c���J�SN��n�¼���b�M��L��U�Nj�f�tk6�.X�7�[�xv{4]D��pGy��+R�Fꗕ`�*��I�| �(^�6)���Uhk���D�E��)�AYI�t��0v��Z:�|�T\�y{snA=W~f<�A(�]/62/��(�y!�m���X!��N: �@��96)��p�����}\�:D���J�V�b`u��e^��
�]��p$�A�
"�Y����P�U�!�_t�q����|�/�\�^�gK���:�}��8��b2���W��fC�ε�xj]#ݯ&s	Q�z��;�A�>F�LXO��-�^�x��h���lr�!m������-���y��u،�xj��N:��J"�e��ԚR���#ke�84"D����}��BS����3�b���?��D=8�Ή��W�c��U���˹n7��	���3/�vA�λ�gN\�d�ޟ�K1���[i�G��N�i.Gz���̡!���+n�̷�~�N��'�|y�%7$pK@��gg/���[G��m���ܸn��v��\]�_;/F��G�ۃ>�k�}�Zm�� �����9]@m�(��nZ��	|=�v��-�x�(h���p2x��5�>�>�$Ć�"��v��Redn
u��*�5j;�NF��y���L�:0��}T��4��a�8lk�E�Ś��L�pN����X&O@���a�=���n�[�8�ɲ�\��1�\�s������=��d��.}Y|��č�8�;Z{#�WR��f�>��(��U�]�;�4��`=�n̙��V���}�ä2s��b������g�ȣO0P�@�t��,oO�r��Sn��ׯu��6?Wa\�+�_�64�߯J��kD_�J;c0W���WʔE�qxt�)ؖag!����[R8�aK����s��Y)L�F{�P�m�Gk�sC�L�06��z���O�Y�+e�t2��+dR��F�αzx�3s�g�*���l���5S�P�Tɩºj6�LrE��WHܹW6|��l#V��6�Y5�O����5��؍Yx��u���t#P�+��]�E����<=��]��~z"���w6��}�s����w��:qe���k�́.��.��ˮp�e���.�Ηq�C���a�z�Ϝ:� �$4�F�yݞ��NDS~Z�yʹ�<H�Gc�{���\Yz�{z6-yx���*a�y�D_.b��b�b���U8�����X���b��4g���8M���\�V:�Z�xg���J$��2���)�ek�Yu���M" ,v�Нzv3���5ZmG�ᒮ�F��9�̐�g�fX�	��f�7%m6���bh�l8gO��3�UEGo��F���v���\��:��U����3D\v���{ݳ�y��`�D�L�l#��rDW��U���=ù#�W���!�����՜�����3�(A�Č�.!����NɃ ����`���^ ���d�-};�f�}[-����(�˚,�F�	�cS4&���_�>�����y�1ݴ�
��$"7���a��͜��n/��E���tz̍r�&�S�u""�4���ER��_bGk�aΊaH�	�UM�m���Ez�e@\c��J4uXHT��n���t�7���'H��;�IΙ��|���sx$����Pp�'6�þ�Q,dut�C�t��~}T�qda�۠��u�k����:llq���J!Ԉ�U�q�[���v�..�q<�ne�n�&�,J/�'Im���w��jK���+"C����CY2#�V$��bT���ڒ����V���WC�[�`H�H��痗��35��ۃo�<>ɣ��E��ٱQ��KT���ě���bR� =M�{���i��G�땄hr�l�S#:s�K��)E-�ӫ<9j9�v�f]͊1{��E��pʀ���p��U�8���
�D��~��s)�"E�3z	u[��soDs-ƌU#��]R7��M��o=!�Y��{\E�z)C�b9]�L��Wڡ�9=���z�ja����/�Q�sdP�<F��,�ƔF��9ק�7u������)Ӯ6f���D�BIt��L.Vߦg�M�ߎ3���X�<�n�c�%ٺx�ݹ��mXvr���9�t�����28S�b��Xcb*T��h�L�c�y�m�[��.����i��e�tvFu���%X!��!�t�Ҫ��C#H�R���h9���c����5Q�k�hX* :eQ]N��/�U�_?��*��<�E���-<��a+y��y+�`�F��q�W�H���etF9g!�g���Xj`옍���7=�4�R��hfwg�����ul؎�f��
ʑpu-\>�k��ޤB�*�9�4_\�\��b�;h�<d�����!�a�.�O<�c�o�q�1�E�3]+fhYf6�4��u�ὺ����u��s$<�(ĖgQ�t�m-n����_=������`�8��n&��[f�[Ħmd"8/;�dM��28>���=�-���;��h�fs"�:��A�sd#�	BFj���L)"\j�.W	�z6�l��V�(^�������E7��+\��&Nx&v�ߢ=�~wPr�P�x���C���^��/
����w�K���x*vc�Jw���-�˃��$�tdmT�y譛Uj군����[�I�y=�=�o)�+��B�6<�׶l,͕7��S�+����7�y\��������=r���Uu5p�*�Y���tȿk��Y�@�Z�A;ݮ��|:P�ĬC[�{H��Īb���R�+�BԣwΑc�u9�e��&T���z�Om�Fԍq6�2R��oR�D�Ն����Iu|�,T�\(�לPΕXR����weM��.��D�ek�)�A^�Gdt��1�6Q�˚�D:�eː����afG6�.ȩ���>��Go$2�}*␆
1#xז�T���E���(]�G��zӻә[z����m]#b`u��e��D�z�E8`w���+�,�1��b5u"6��{u�Q�p_끼z�xK���Yp���	���\;���w�Og^�����G�^���O4��V��Җ=H�&��L�q5��^.����9A��d�ˆrٜ*��/,'�`�D�$Z��h�3.���ut��8�����8z�B�㼳r�}�+-�[}9�/Y�0���.xн3�����>͊�,�IU��NY����Ь��W:�W���/�,���IT޽To����t�������х/
{�W�w�O`�T��.��-[��>��Bu���#1O��X�S��O�,W�Wh���ԑJv����T��\����e;����zx'�<�z}�tJ>U���0�Mt�q�r��N]<���E�&���Ł�$D�v�5�ˈ�4g�dk�bCU��I��`)2�7=N���̼7yy���ٽS��~��t �����	�v�,8Ç�rLQ�fsT�{���ݒ�Y��U�{FB�g��:na���42l�q"�hǕC�:�N�K/c�;�}|\h�X�H��]�r[fC	����7���*���x|����y�e�o\T��/�X����)�uC�>����������ز詇U�C�2�5��E�X����]��c��ʵ�O)�빜��=��\n�Xy^2W'-��Z"��Q�0W�C��TE��}��۬�șiA�����^�hAxs1�M��!���B�u��g�ʐ�Uۂ� ���-��s��v��w{Ҭ�ǏP�r���j*3^�ص��bQ[Я��֎���{A�fH�$�_�0m�
�Y�bZ�4���bہ����L��R#(L��IW>��9�<ɳ+Q@�w,��0P��s0e��bçZ{�ܥ�Հ���{v� F�3r�>�Ш�YM��tu��N:Ə�˝�R��4{϶�J�V;��=���Ԉ�b��|�!�i}�pZ2j�wk���R?6Įۨ�=Vu8k����k �|k@�a橞y����g��0h�'rZU�(���0D��fR���Q3n������S|w�B��	$�=�1���V�I*t&-ۧ7�i��6�Ћ*��fX�/6�Җ��7�v��P���[k2�������.�븻1כ�]���}+�Қ�����T7C|�Mv21�$�u���p�k�K�z�z+f�<^Z}3�#ɬ��udj����z�Wr)d�8�W�����d h��m���BA��+�:��u� ���8����$	�j��Ij�/�x&���Jī�];�;2D']kl���U29��'T��Ѓ/�톬�+iUD��Z�a\��I�ۅ|,Fw.���oD>�q:��lq����6m�)�a2��<)��Vכ��#�O��c,����#�h��#����/`jOc���#̨�P5Y�T�NK���*3��+��RpiT�c߳*�w���[ye��]�a�6u���ؕ4zڹ�Kmꎶmm]xUsNkxj��w����O�*K���2�w�#���z&O�f�~�}+V%J�)��v���`k�h�9�1�E��9�r�K]E�m'h!��赼�K���s���n�34R�cVs2��`�DNZ�↸oE��F��Ӑ�[2��b���j�t�e�Ⱥ�7ym��l]�����?S�%^�%����3��'���<�w���F����B�*����å�u�ٰ��oe鑻@�� t��r0t`�M�2U�_�����Λ{I�"���\�I�Z�i�y+��7��+Sf�@�
_z���˜>��6f��[����NDm�=�{�G�V'�p���u@=��z�2fP�����D�wh���4���9��V� �8�;��حcn	�M��v�'��S�b��U7Y��{&��J�Oh,Z��D�Q��_+;�{���zkt�})����P�6~�i�N���b�j(��^h3���*&�y�;��ǡ�D����}EP�wNԻ��C��.�p�XR�t���x�!�|�����|���rb�����؍��E�3�|�Suٷ5�8���F�1ԧ�cVU�uĻ6'v3�k�&^afߦ�=�W��y�};+s:���3����"R��0g7Z���}9�[kz1%��U`
10<4�H�b=�}�AR,��QAV)�P��œcU��).Y1��,@r��!�dQ@��?�������
VC�0`�
*�E� ��$�QdTQ�ؠ�!�9d("�,X1?&�a�mV,�1��m���`��!���B��*�*őd��+AEDPU`�R�Y(��Z�H�
�"�D4�c%C�fPհ�TQdE'�Q�²(m��AV
(T��)+*.�Vb��`�IP�����X�Im�U�C������_d}�E��Ɔ�I�Rv�v^�v>�^��n�0[�Ebzk�2�_o@T�E�X❰��͵"��:e/��I)�m�mUa���BR8����86�VE�f�(��#	p8[eVj.�j8Y����Vn�������e^:dr��F��u����;��%�t����S��UE��utʽ��*c�mK0��G��(qB��f۞Y5�X�8�#��K�f{�u����p�.��<}�񣦾���7 �E�X]>�z���
u��EV�ͩ��
(KNK�y��c�޺ߏ�M�@�q�l@FkdaW�؅���D`��7Fm�M�]W�D��1I���v3�Ө�i���J��������z���ٍ,����Ĵ<'.-Z���p��,pΟ9�g���~�Q���])Q;�D���Ws�Q�Vu���e�e����ޟi��;��f0�h�Y�"����}�v���i��:�Ok�U��MKu������L� ߆6(W�\E�2&);&y��q�p����i�}B+u��½>���p4<xe�o�D�`ΦhM%M��Q���獺AgW�VQix�fh�u-��9ֿ�T�uQ�
N��w!T\�ȄA�u 
K������6��j�^:���-�I���ej�<��s/�A��s9o��89��d\��F9�G�dԅ	p�,��k2�����s���y�j�+��zZ��b!߽� ^��"��{�N��J�t��m�i���3o���~��>7����t�]¤^�Qp���ˈj�UX�y�Y���H?���^p��=C*������$�h,�v�zB�l��];��z׆ywWtV'\f�O>�[=\iL�p�2��2��U�����^ŚѠq���{	E���s�im�E=u�k^����ӧ��:J#jr��re�^�ڂ�(�X��$cFG���a�nx_%W���Kk��!�����S�^U��u	�uZ�Ѱ�K;W #>�=^��Y��q��z��(��/�Č阍�5gק'+{�N�i\���}2U3��]R0G������Ȭ�F���>�w{�7��&�ڲ�gHڌ-�+}�C�=h�%q)�j{�d�+��9�g�����Ҏ:Sv��=Ի��ٿtu��:F�۟q=�I.�Ti�Aӥ�8��*�G]?/U�\m��)����k��EdGF���t��qM����!��,3�t�f6\�����GED��6Z�:3S6�	sʊ)�],'�M�����h���<}�޺Y��\L�n����8��ÀT��Tr�vam�x����ܟ�����l�v|�\��:=�Y-�g;v��N��L'lT�"Q�=n�f"^_��:�4����8�ŮO؈>ZvF�n@���f٪n�4X6/bEt�וTT#e��A\�G�gpK%zW{�s���7U����{�"�FD:�gI�$_q��[r4����bM�f�w٠I��W{y�W�k�)��AAN���Y>M�Xr��yoï��21ȃ��_L�(�#��b��;�j�-H���U�|Ur�k^�^)P���,���r�r���F��&��1���n���̪�����^$6�U$7�"l�rg�!�&�q�A@�K�{�4w�PW<�>�IC�Bp�R�&���"��Ô���]rd�gk�?^�FE�oGv%ɪn���M���z�0t�Y����]�](�+\�2p�]����u|9�u���s5�y���0����H�͐��I�^Jf,4����P�S��׶lw�ۈ�j7�L�~���&>�"�p:��S����<h[�$_J*/+K����tȽr�NXj"�g2.���7�v�D'�r��1�yWY������?h��C�Z;`W���*Ҷ������P�FI5m����s�uq3��̶���,�i����y�<��fm����뚩و��bYIX����/���/;��xF���ر'�o�T���ƹ�S��e9"�]�����#M`�tl�|'!H����~��:t��yN;�
��'���F��C2%R�_L�����n���g+�]�T���A�p�Z�k��켌#�a�ބpޖu�����$Ϻ]v;��5�u���q�
iِ���J�������ϲ��H��Y��RȬ�
18�Ƃ� O�3�!Mӎ��Πck_R��UB,�ﮙ�L���E�Hdj�Y�#E�`StE ����@Y;k/�Ij+�����ì�a������5zgJ����3�بr�y%V�K�vCȘ�6\J�P���*f�l�l��)'b&�ք*|�;�A�?#g�V,'�|te�D��Fp�#(NNJ��Kh!d���2����|K�xb��s�?�G����C2b���s�ć��W�,W��Ku<s2�Fp�PNٕ;R^����Q�V��*O�*�]֞�{�(�݀	�!���2x��5�>!Vy W��>PǢW ��9��-�������eN��N���5칮���C��R��N�E�Ç�`�)�r.4�~�ͨ������7M�uEM����g�u�����ש(���.�����9�P��>�*��D��ZK)�PX���y)]�Q�+���׫#I߃:&�%�%t��Sn�P��vV��@��iugYi:����ȋ_ݽR�f����m�3wl?G���8�F�v�}'�v;�:h]K"��!^6UsChǵ\�s���쩾��r7����*������j*M_f���c���c*P5�,��4��fλ�um��z���bv�^�T����{vf��銇�2׀����-�eʛ�{�{Jg_�.g�-�����;�\�}��"����U=������VW���N_��ƴB�G7o���x
I�L��2�/8s�N|���|��)���K��mθ�YfD%RQ:U&܄tS�Uo�0�\���9��H������^Q�ڝ�����Ӹp�P0*;�8Í��c���2Ͼ�d���
��R���#��Ͱ�{A���-b�M�\k�b��X�ACkW�Kh��0�E�b��z�B4�qBT�F�"�ǐW��g��my紳�c�9C�zd��S�NXO���'>��F�<5c�׬�8&*��5�3^V��Ώ�cg��ȓ��r��aK0���`PR:-G��Mpϡ�g�Uk�r}V�}���/���w��ׯyh���Lu�n@6�)	�17x�!�]���Q�]�7r�T%gK<��O)m���1ۉ�[����uj������,��Q7í��(GBA���H����Z7�?�4*�?3�0�S�M����YY��%��9������v/t7����ӴJqi	��e�>s�
�*��F	eg��E�;�▧C6�U��:��ctآ������SYνFH�.�6ٝ3,�'�ff�I���6�4M�������C�*0�N�����(�_�9&q	q�#�\E�2&('d�����g3���Ac3��qnL�k�Λ�v��f죕Y���s�`ަhM%M�,��÷'D��j���'o���>��a� ��T8U�gԬU�@�.���i��{g4:=f�e,�ΨZԎ�]�DK�u�9ӷ�) �ء7�UM�y��������
��<��T���"����s�(&8�'<�ݶ�O^��h#��C�o�+{�e���ZW�_?WD
��z�H86�v�\�$a�6�#o]i�����y7rt߶8��tOhZ�lNE7����{�.��Ǒ�"�R1c#��PG}�ݳ�dgCnpR߽=�mX̛�K5�w�=S���ӫ<2$���8ȥ=^<]¼�U�W���͕��{�kLA�ϯ����ר��D��*�^5��J��3�gx2��JOa�]H�]+:������\Lۮ~G���&�y��z+�si�Y�Yw�P�h�
	�R-��ֳiJ4ll�"ASx�oEwP���u��.fs菮�j�'�Z�:Q1Tb&��'�g�X������P9�]0K�x߲ꑱ08��<m�����$�a��{j]��K:,*�&=�;�����C�'P�PS#�D���g\�a�߇d�v��}sӌ��4�n�ldv�~�,�t���#fo�}�bO��������Ծ�MW�^[�k�Wj�P��n�̑Y\��R�Uø�挎���̬3�t�f5���`��na��Ԥ�--�L!6}H䇹+`T9�j���I`�^D�R��*��G����En���ɍ�9��9�$�Ϯ�W�h�f�����^�O��-�n�"l�����-��؇�F�
�}�4��ge�;�ܦWA0tc�r'K��s(�9|��S���]�F _r���VMy�ZQx���Ȱ[�"�w(������Gf�:]��B3�w���fX�/ˤ���q���s �z���N���5R�qQn5��[�xZX������A�[o	�^�."i�y�M�a���'ں�ɤ�컿�
�=�W��u6W7�I[0��� UTa_�Ӄ�q����p�R�P�αZ��N%�Q;��v̕,GI�es����gv��E\�X��\�b�p�=�ȴpIOF����U�m8H�K���1c��ƹ�Z���Y�y,�_
�j��	��QO=�+ # k�c](�6��-n֑6�������"�l�JK~���CwY8��#Nz���l�4.&E�b�F��$�;V5@T�=u힛Q,�wqw���U��`�{ȋ�.�%��p�}r��V��EF�iyw��"಺�Q�b�}�}�+7���POr�0�W@��Ԋ:,	T���BԸ�Q�Fڔn��i���`�e�y���x������~Q/c�s��&��30�J����r4�F]�4SI�f�(���(�+k�605d�!�"�e�q���,��ڂ8�8��t��1�����:P��꛾�鄊�8�JE˕juǯ��H��e��qH`���� ,|����j��5O;��G�ce�J�_^�w��`�\����
�]���"�
�
"ʘ�N+W<Su�ٛb�h���E˟Y�::j��5zgJ���:#ٰ\2����&#���)Ju���2ηH��ۿ���7^����B���(T�6zd�C<�
4^�c31���-�������Ԣg��._n)�YK�H�����\��g(�z�**��bK��D����1�b����g��2���LC�b����si�8����ڏJ��������%�yY�Y�ޘq��#��G�S/��=[�fw�Rq`��N-b��?7!�A:gdŇr�וMz�y�(��Չ>_+��t,W�%� �۾Ɏ���̊�c�F�/j��U�FY�3�b��f�m�v�b���r;+���Z������se)u���n4�01��X2s���hϠι&'�VD3}'k��k����gS�*�En�NϯU�5�4�^FB>� JN�BaZ�f���^z�I�̊ƙ�NW��&A��fyE�Bw������d`퐉�d�U�ha�X>���&n�ܗ�=�����wNa��#ٻ%�24�9÷p��׋��Vppu�݈�ߨ�O��.Z����\v�~�Uð׷fZ�{A�_�زf�U��u���z�8����i��՘�SE�R�?>��56�p7O��\n�;��I��5�-T��U�u}R�x��,�6��w5���'�;�:�1q�g,ɬW$�n�\�鑄̅� ��^[�ZQҡ�0�w4��"��rW~�l�Q�ߔ�oX�=)�8d�b7iI����ƴ�kt$3K�k��`�Z��⽘�����N���].����.�X�V�"i\���V���:Ƶ%�h�b�հeN@A��\�\\.�V���}�ֲ�aPd=]�d᷑󦇙�!�����H�
{�ul;߯��w^�ۍ�դ�~r�����5�W\lJ��y�,��з����ɨ���V���Vb���E��%w�&��@Îg�_�5���x�9�Ip��ھ�p̶�%���#�Ӗ�.��F��ȋ�.�E?�儿�״�6�R�pxk
���u �$�TU�ljv��7zt�@�Y��'}*��	����q�S�����f��_=L���#�����)ސb$�@�4��0�4��`ߜ3����l��|͝|�+���B^fו�R؊([Ŵ�Vr�L?+�����hddT������$wLlΙ�e��L���u�툛����:�j������#�~����L���3>�(A�Č8x�^�l�ɪ��*�x�IR��}g�!�܉��l5�di��gM�v��_ً����ٱJ��w���o\dnѬٷr�Y��έ�ş]��1�%���df�z�#�Fl���q�P�.��n���|;\W����܁������dV) �ء69Tl	!�ڝw����UQ��C�ǎjD�V{2�X6	���v����4g��L�,&�u���D��A��T��cpY�8.Оۮ^L��S�)��&��;�m�%��� qd��=��lRͯK�ͪ��(=]���Ke~�IؕDk.3��Df�}o:+v���b�-�����3-�Le�S-U��Cy;X���3jz]�9�����]�a�!\�҅�4v��W:�K���Uc2�A��-+�s�μ��ə�5jRޫ�䮏7᲌�ZyT��<qN��,3nD������1� �[Y�ws8+#3�U�[K�38�Ƣ�XJkR�ΰ�fD�h�gܚ�U.��&Qo�˙�â��t�uq"������#�}X�@vi,Ϲҫs�f��c����LwRD`%s�}�#@�Gm�b��Kg�d�%s&��p���#*΋��gάp�'!��u)�:�	�r�چc����eX;��Vړi��V���.��1�v�O��棃���Ob��lMN����^�Sep=�R�:�@4�ܹFX{yr��p�7�
���4mJ�G�ޅ�����<��g{�pYR�`�`���}�4(5�B5zv�ě.���Sn�H�fH�9D��}4�k�3�D�mSξ���痍ju������>Wt(�_q��D��NN�M�``'ZT�=���<�u��x�=7Q�y_c�cx�͢�����b�j;�s��:u�L��t:�ꑉ�{i2��/l�{꩜ĕ��j���j���wl���*RܹP}�e��im��{ C|+اz�����gKさa�&m�Փ�'�Y�3�MRM����9�9DW:�e�0݅�Z�-�\�Æ��eY�h����į��cR��ӷڪ���7�oV�6Ø�q��e�U�;�`Z�-J��dݾ��MZQ�W!���H]h�<�B\z�ѓ��R8��\~3�Z4e��v�#>�S<�w�y��,�:��,�bܱ望P�Fn?4J�%8I}	�.��ʘ���5�e�ҹ�y��s1w.W��5��Ԝ���R�����(��N�kP�eLwe�w6w�'�w.�}��u��x���/�[�밠���)�L��xˎ��F%R��\�ׁD�ˠ�Y0�q,u��3�#.���rZ���6�1h�Pzk^���Nz$LteD�����S�V8�;D�#���yA-��ѫ�G+#㉾�3C�����n�\iKTdB��/���p�����)-1E��d޾h�MZq=���[c�K�תq��,�f�L��T+��
#.^��H�J��w6��No��R�r�0uD^CL\�-�V�N4�0��V��lAL�1gu}�|ȭ�"���˜|��ϡ�%�6�ݭ8GG��V!�����L���m��6���rJv���ʠ��FW�de�2	D҉�Y��;��fYsݜv����O�I�>���欘����,�j�" �2�L�"�bȧ��ݚf*�"�Y���(M2C9f�3yG���'Ԭ,UD�aRAH��(�V"*�Uy�3IR"��U(�X� (�+
��
Ȋ�����ȱ@��M�*m��b�dv�
�E��ێ�P_V)Dt��"ŋ�)AA�)!X���<��������@�CN&+),
�V�X��cĨ(�q�BQ�t�A�^XP
(M+�5!��PRq�J�t�b�׶2)���UTa/���+"�b�T��(���&5�U�T�,%��Q�h�����P�̴��-[J���IpI�w���{��2^��7���ǔ����u_f ��$ݺ �����G0FL��R����ߊ7|�/E�Y�~��-��gO)��K4�V����uwE':gcLS;:iU��@P�J����ܕ���(dq�:���qdaIH���Zv���&�N���B'K���-[*{�[e/jYw$�Z0$_JF,dy�{��yS�xyL���i�#pm��,���и����VC�ug�����dR��]Bђ���s�����5��byN[�ij}��p�jg�Rr#�=K��Z���.7�R5���J�5.xqk�5��)������-��@ކlk�+�rsF��G����Gw�xmי^��U�~��yGʧ�y7ivD�^��ˍ(ϫ:�yN��6�q1	%���C�KL`�m��AΫ���f������Ȗ���ʁ{%N@k�iF�p�2۫2,
t�T2+l@��<;]#W�g�k�9+S;:u��>�9!�^��C��f��䦋�e�H��3�X �L�F7��n�+.QQe�G5=\g0]�;1y���#FFD:�gMD�B�q��#��{�hŭX7�z���9���"$������D:.�gPF��K����W��<�o<��k��iܒCt�rso6�	��@��f�t��Xs��c��V�Ϋ���*y�BAju#��.2f��޴��	i�ڹ�S�0w1��nd�������.�ƛ�*��sЅ�������a�PP}�e.=�|ז�:�P_�n�6)-���=����q'��F	���D�9���B}y[�"�����oqPԓ�����tw>Ȟ<sDAiH>J�qќȫT����A͑�ɞ��BE��;�*�8�u�U�c�=�����d^��8hr�&���"�yXr�Tŵ&J���
��*޾�e�џ1f�)�}�L@����!]P��J#���֑kv��Np�AGC��?�jV�h��]�2R=(ӕ\n�q�8׮&�1��*yM���)
�˓��m˞xӪ^�;y>���G�܈�|�sNJ�KC��T�j��[��5Ç�MV4j�{S�o<ś0���`���ap��a�]H��Īb��'�Z��<���Mc��q�� �T$���4�R4V�aD��9�F�����U(E��=�!�à��M�Ř�q������p��t`�0/e�;Ўޖlk�(=�#�#�|��1i�{���
�i�z_wE4������͗��S���>ߑ��\Ϲ{�q��;�˝�a�ݖ����XXg-�T�+{��X��8#m`2n���w����6c{~ٚ�,��w��ѩ,ǚ����.�d8v�taJj}\,�ږ(�_�
M��ӫ�YF�y�׉�r!GS��}��Hм��6�RȬ(���SȁsC�O^�J�n�6��Y�}�l`�,ׯ���L��(��uD�^�Ǒ��Q�=�o.��k�O#;)h����6#.�{��gMX�F�ƕ��{s>͊�N�u[�����.Pu�
��=����ק 0���!WM�A���=�;�v���>��2�z�[ϯr��L��N�L�u΅Fk��+g|"+�V(�?���p�z�ֲ���tL���ձ
"}x�/��h:ֽA��4g�'l�	[pZ1v�͓%ӓ��#���k��K�g	{�:о��[Ѿ>��$D���2x��5�>�>�$���Ȇiw��5�[��F_,b;J-ɝ���ٶ2��C.i�dat!����qRt�;�0��2"Ĭ�]Q�]75@�f��̩�x�*j s[��枻�:na��퐉��+\H��-����؊�yث*�/7e��eN ^ǧ_��`N�y��7�e��P^/��(�'W�qx�z8�5)72��ag�:��ޯB�yuf��v�Ij�K)�	}O*�"K��N��̻cm��Y$������Sw��<�����Jb��3�]��t�\��e�uu$
�<�Ȉ�v�����}S�B��Pݺ̍�&ծ�K��y��jw��������#J�ogٓ:����:�n0+�E����;y��}
!UK�Y�j��9�)�P�j�q���db�Ȧ�e%rrÑƴE��v�1��Ü�\+�,$Gy�ܸ�iJ��Y��(Q�s{)���,Ȅ�J �t>ZN�oINҚjP�^Hgh�����M�"��;dPQ�ڝ���X�33�74y���4��|��r88m��X�=J8�d��4t5��\�]b������>{^���ڝqߗ [K��3���i��x���I��Aq��6)P�����T�썈E�N⫅�n41-�ۿ?6�Ѽ��LE���>"����_{s�0*��4+�5�+㈱�ǉ���%�����Dtf���x�Y�r��hJ�b�fh;[Q�z�GFL�g�<���v�C^T�������hi�Y�8�p�R�$"K��>�R�Ҫ,��t'�lN�f_��s��Y�VoE�-�w^ȡwcMc2�22*k�Q����]0l6gL�K,�=PﺜT���isK&���x+��A��f&�j�U��F8�YOy0�gd�L� i��f"\
_!���"g���غ��Ю]�����j�Qc$-�lܣ=z�D�����/����
���"�t������s��=kq��w�ȭ� ��Gu�mxZ���q���cF!B6$a⋈��ՓQ5��w~򽜻�0���#�6�hj
�? �K�I�r��f�-� �}]����`�!�5}X�Gw��Ж�s1e�\I�Q��B�*Y�A��(.����M"��Tq�nwO>ȭ<X���]*"k�)�<n��E( �=�\�6��ۛw�^T��)u�%�;a��;��ls��J4�V���R8�v��W��O>�l�q�o8��R�Q���Wm���~�)�N�
.#r5EUH��8F�܄S�Zv�e����+���Yϟ(��['
:d�bzQ.��5♁"�R1c#��r��r�l���o2��^�9$��=�����a�wL��x�����V�8c���/�-%�4z`d��/��� �dzd�KqX0^�WvJbUS�%lb��aH~�0P5�v����j�|���~W��?K�2�ĩ\Ӭܱ�6;�-mq��ebx�c����
dqȋ�l��˪E>��R�Ţ��SX����weڭ�LX LB��λ�e���:�T?f]w��~G�+�V�V4y��h:X�<�'8lW'�w�,��\���7r�8�L���wj�Qd^����#���_k3�f�n� �]�(��O\Q�\)%���:э�N��#���8�l�EVu2�#fmϸ��$�]l�5������tS�?<���
�O��.�4.zܳ��^�(�0k�iF�p�2۫2%�0Y�r� t��=�G%{Ț�:��et��*g��&Ϥ
�C�!�ͳT�Jh�oŗ�"n�w���o��9&��B�y�͊�X+)�=
1v�;�Z*œ���R�0��r�+���2��"��br4�9�&���%j

t=㢲&�Xr��ð�E�r��;�w�'�7/B��sOe`��i&}��f-���b��D�Ȁ��N�B=W����f�V�YS�]�{�Ǧ,���M�����7,��_�JTˈ���E50cCypE ���&{ ������ˋ���	�&��� �6iF1xr�4�Ȧ��`�O�uɒ�ܒ�֫On��ݢ�=�j�W��!��V@G\ȫ�J#��z�sz��:��fH��a~�qu,��%����]#V%�<h�;p�2/%zW�#D�2;԰�8�ɒ�����❤�cə��	
�����"B�#��c���*�U�x2ol�dgr�b�o�
9R�Ad��O�������Z��łQ�r����@�}X;��l.�}5�]���f�l�Sv���ď���s�G������-�Q��Ky��0�pf��ۯlߜ�w��-�%�� �)hO*�6�}���L,�b����i<3_W���e��9��(���P�J)d9�B�is��.R��r�/F�����Ú�-Y��!�m)D,�<��^��#TM�!��Jc�Q���i�N��*���h9[ê%�Ф�C�R2:z!�p��B�Q�Ј9���'�Sڂ:��$���С)zћo4+x��r����Ѳ�'�Z��-�Y��ڼ|�^��}e�P�fa���e��n%�!i�VA��2�3�"�)�0Nh_]3b`u�ߦyc�2$z�Ai4�׬�q��L�>ɩS��Y>� ea����^�n:h(н3�^����ϳa&���l쥮�:��{g���lF
�Y���q3T�$�D��\d��Z��ѹy���g��v���Q����آ#K̝5�dV�ɤ����2���{�f(Mxj���dqW��l	�ֆr�3����M�1Q^Τ��#��Fp�Rv�ҭ�.��9q�J��g�`��\+E��b�ώ��	3ӡȕz:w��/�q��a�i�'�q��٤���<���r,~WĿk4n�o1q*�rҩ���}�"��.���=DOGM,UA*��q󼕜�!��]m��L�f�.;H$�=S1k�6Iu��\>�~b.��{��t��_��u�Cr.�/�QW���^�E�SF}@�$��9��0inn��37�"8��e��q�N���E�˚B/#�`�5K�I;q�%e�-��X��ܻ���l����0db�0doxa�,ӷё��F�)���j~�40���8���&wz�y�9�r�pdkG����ZpU�5�c,�´m�@�l��uE΍g,���z������H�F�p��k۳7�L��,�n"'�r����U���۔����k�#�,�F�{yHF�����}���N��J���pE��b��jj����b~n�����%��zo����R8�~�u�ۮqYY:��1-]�͠�/O��굑rQ)t4���.�\����7����l�
7�
v�5#_9��k���4jX�p���CO-Y��!���K�苖�������O^�H�0���ԩ)���Tw\�!>%�􎠙��a��2��E\��t�m�����3n���΃i�,,��V-��5`B��G_=7������s���æ�nq+t!S�nD���Cҗ.�uw�i���ݕ��Zm7C�\+w�3@� ��J������b`G0�R�_?���m,�j��mK�GD��wϮ����t����l񮇛��G����Vu2�T�"۔b�^�,3��R�6#�j�m�R9��z�c#k�n�-�&��Y\��h��6)�"	�*��L�kj8��u#�'*^4:�9�Thfl4�E�zk�N.�f��!� ��D�q�HM�gO�Υ��U
������r�uRؗ��c��a�Ҙ���{"�݆k����S���G{��`�lΙ�5<��ٳQʷ�iͱ��t�����f�.5�lv��;62��򥗻$�� �6(@�ŷ�x�w��s����݊Ր' F�`���00�y���܄{.h�`da0��7��S�\FV[�m_e����<��|8}"O�j �Xh�E�"ȳ�Q�9yt�"��m��V����^�3�.W���^����b�Z� �q�� {&�*��$3�R�� �Zϲ���ݞ��ۏ�_{�fu^��q<�.]��PLu�d����������ض{5�6�]6�^bYOJ4�;\m�:�������F��ʩ��ې���Zv��voj���ܰ\�7�n�ft,�֪^ �E�јR�D:T3���%lێ�N۝���)��	x�n�U�^�c���R	�o��d�ɨ��mQ|"�t>x&�D�L��zZ���ts���&dX����R����Jtx���7��к~����V���N����ca:lJ�Ez�I�@�`M��b�<�+�L��!A]�k��)��7�ZD�WH��)E-�t��%��8�)����䢮���c�8E�����-y��a�Q/`^�#:e��p�)����+�F	t�.�#������`���&���&���Ef�4�x�
l3cP�1�H�	� ���:��5Ff_.�M}���z���cb�p�ӎ��(Ȭ�e�Hٛ}�H���,����{_��s�we�y\��0�g�b�,��R�TدJ�"��f�iW⛚28S�c�v��d�m�ʘ�[����-q�h�DP�u����X�6}\rB�2^��r3D�p5)���͚�p��v;k�6�i�{Z�B��dx���>°V5�[o�����X��22!�,�d�ذ�QJg�ضou�t��H~	�LBp0�k�8�L7�>����Y|,9Wo���~ 	����>�q�7;�pO�V� /�B����E�^����d�:�(�R������� �$�� ��� �$�� ���$�  I?� HO� 	I� @�� $	'���$�` �$�� $	'� I( HN  I?� HO� �� �$�� I?� HO� �� HO�����)��a
����),����������0��=�A9��fz��`�)�P�I����S@   h�#�*���  ��@ `20110�L�L�4�MS�2(    RD����LA�@ @z��jcT��y&�����P2��y�H����\j|��@�8�+�YX�xH�-�xi�a���J�}�U��D�b�
��8��eZ�c������z+|��L��&6�Ԭ�k��jYB�6В�[�:&�Sۉ.12f�؜��3qrGkp����I$�I$�I$�I$�I$�I$�a���N���O.���<R	�w�V�h��bbbrj �8�Ơ�	��jG�d��
�%,j�m�p�US������<��� e &�沣3M��歓�����k�f���F3 da���"$ۇQc�$ޫKWi������WX^P"#&˝��ɽ��bZvŤzz�b��H��Ԁ*#�"T�,��fJ�4"M�:���̌A��Rv�}�S�6����ecPчv��j�CNM"!��Ʀ�$e�lvt�;5/FY�o/K�c~w2t���T6lf�R����I��P�=�_0S5�X�Njq]��t�.1�qAm���i)"�D�Y�]�i&�+u�E�DP�"Q$(�k�	���M�^�њ��������� KA݆���թ��#P�%�2'\3�W����.��5��ۅ����2��r���v
�J3E�t�}��ւ�c�ȃ�Zy�a\dXt��i(Ԙ���M��� @\;��6ph�BIfp2�❉��@����<��RG�T��L+�\H��Z�g2^��� �}X�d��ԐP�^3��d�,�q�:��<IVp,�*`|��RS�����fS4�-�׊b/FW|I���c
a9k�띈"o|p��@�V"!L,2&J���YN}��ҩ�A����-KB݉���iMOx} �$yq�zP3��2��W�ħG�����|�z�~�5u�2Em`d�&&ZÁ4h���U�1A<�X(�O����P[�=��GU�f�% *�D��<0���k/7��%���V02i�o�2ϸj�_{V��Ғ1�s!��boW����ON2%]�^F3���B@��Q�$pY�Ƙ�����`���($�$5. ]��`��ف<qH�C�B�x]h� ����DB6`��_0�}e\��C��v���S���EN�Ԅ��=Jk/�Ri�mCZL	ˆ��I1��dl7��<r�O��5��1a%��Kr�JJ��	��;���k�&H�d�Z
01m��bX\�����JT�����s��-T����$�&A5�o�,�k�\��+n@`C������/�s�!��~�:��:�A�a�.�D��-�,��s�$AՃ��1}k!�"�Km�B��=iQ}9����h;c����nӯ1 ���֐
j�n�!�Z�fKyV��M�9ԲfA��̐�rԎ[��]��B@��