BZh91AY&SY2��gi ߔpyg����ߺ����  `���հ  A� 4W��2ց  �r�    �tА        �t:F��ǁ�@�m>��     }   � _W}��WA����)�[�0u��㷟M�+W�zxh� ��5��O��x;�ފkTS}���pz�{�� � �����H6·S �����w=:�ij�-��u��:P���<6ګ���^Z&����z^9ӷZ7����ػ8�H� 9�  ��v`�ݛ]n��pn��Ng`�p�:.�;���� ;�}��o����k�K��'pv���;3W�'� K�^�Zۻ���m�l���F�mwD3�����u��w.����kk[���=Ηvm��c5�k�
� z1�  y�Ǧ�}u귃���9�F��pF�ρO��m��z�*���sQ���6��      yY )	!BH�DH`    P*��h~�T�&#��	�##j��D)*�bbddF��i�	�i��Ԁ��Tb FL�h�24�LI�@���` �10  �#IL�4
f�T��M0�=OPiA�M�z�(
��OJ�D�Hd4�`���#&!���yI�
^w���� 6���PA���oA�!����*��(�Z�_W����Cg��~T`e.O�b��;�*�����I(%I)7>lU@q>4��s�Mb�.	$�I$��3�
	�Cl~���O��]��t��� �1&$�1��2��26b;/�h��/���>�Gy�RĽ�i9���l��G簞��~�N��'�i~'>��5�W��hq��wˍ��,�$O����7��w�U��zI��%�#��$�C���!�a�yl�j�7��Y�uvx]���~VZ��>0Mx<c��G�k4u�,I��Ci�C�Z�Y6h��ɯ�2hMi"y!����='D�~��$D=�$+��C�'<��d��8�GY"{�i�O�~����D�'�O}ߓ�'��O#��[�8=,����IO����{�����Yq"'��:=�(K�O<�pf�C��"s�:�_Ή�R'v�4<�O�<Yn��2k�MxNP��Ot�����e�9���p���Z',O'J/Љ�:'�ؑ!��"x�H�~I�0�!�5@�t�:s�'�p�|Nu�>Fx�h�$D�$D�'�4'�e�A/B&��8=�(~K�Ν7��ȑ/�>OD�hw	�"pH��&�'�<$M�D�RpvB�}'ւu�%�f��8�;b2��k��"o�:D�����Y�pA<ԏ��4Q>��!>M�si��OxIӂsI<s��t�H?.D�AD}ʉ�D��N�p/��؝��rr�S�o�5<W>e�v�;�cȝ�~�O�ӛ�ml}�}��lN�Gĉ�C������|�����H>!w��'�8+8k�ND��񇭬�k�ߌ����w�+z;i\Dz�����4{�:T���]ҽ�8(��&�Q�i��Du:{��O�dK�T�L�9���R�ӧ8lvԻ�|jY��9ƧI��|��9%�YZ����s�D��h�y5~f�����=�ʱp5j�㈏f�|�5���b_��>������'�#9QgK4Ϡ�����"�m	;S�uU]DFD���'ȋ���{��=Q�����R�u'
d�Q�*"mjP�ڛ4?j",�Aʛߪ'
�S�a'��"<$DROV�#�TD^�O}�֥9ƥ�}>NuR�e�Duꈛ�R�2|��U�(Fz�&��jY��FUO;���yQ�*Yj|��U9ឨ��jP��R�>�'��mԢ�]D���7��d�֪"/jP��DNm�dO��%���6h����j"����[jq���:3���9g�Sq5B{2����h젦}O�䣔#�G�O}�}sDѢ�F��{ʏ�W�ƥ�/[��F�H�T�Du�<y|x����g���^gh��V�b$%�>{;�Bx��|r��!��=���N�v9�ܲ�J�%t�<�D��E�)�J��rx�Nת3�p���%���X��U�x�<l�ޛ/�\񇖇O&�L�Y��;3bt�UPS�cŪ?1s�\�}I�RwT��5v��3)��z����g�Vv�4F�8�eg�Y����{ڝSя�Cu���FV��dg�3݌�^�3p����=O}c�7Q�j=���$������j>�H>�v�z�SS�:]%m9�'NĮ�wR�;��=��k;K
�`yf�������}�;�y975bq}o����C��}8Ml�Uja������zl�]J��#����Կ���F�Գ̺U7�\=���q��Q��{+��{On��l���y��y��M�t��9ԣ�|�a�p�F{��5���3Yկ��i��=�<��y��.��l�F^/n'���.�~3�f��d��_�����/.|�ODu�(~FD�D�N���͓��W�'����^M��I/��ӄ/�t�Y�����U���J#�ODN������lK�c{�d��vR'jX�y)<:����ʳC���H��I��&�y6��h���c�J�D�O҄��D{�_'�D�5)�N�"�W���+biܤN;�����En"G��/���:��U�FQ����H�bP����jR&��D��D]J�c�J���MwR�M��������S+��ܤM=���2�h���c����eY�O��JD�^4:�}��r�8�R�n�ԯ���D�u*���H�YI�ze}_;�����9�WM~�/�C������+D��\��d��A-�V�	�2�~�T���Nz'����S�d����U�D�'�p�Y]:o��T*�*���,1]<����������B�������eMW�nI�<�o�xY�=�WnxD��<k��<�ӛ��Z�n#����?t�5,N<��'����H:�Rh|H�US�I:q�~�l�Rˑ����e��z���QӬ��/��ڪO�G�d4��s��s�} ��������vޯ3����j�4��6�8�5ӵ��F���V����o��+����:��6��[~���1_q��;վ�&����U:�ܭ�Q��3ݮ���x|S���t�9��=�8`P�����9��5g�=��6ϽOa}��[��:s�o�5s|����(yS�y�0{�t~Ny�:6�PVO6�Ǫ��Κ�w+=�ړP�6��f�H������p_w�t���Nx�ɭǾ�go�%�Nh��d��-�5�=�:N��$�'4D�}V컪����?�
1MeOL�*z1M�5�m�V(Y�K	%����R!�DK?�\�f�0���,�����,���rx��MѤ��g2Iy�A�F#�y���vn��4'y	%���'��=�{6 ��xCftO2)�vx���&���D�`L���u�Q2Y	�m�br�>P yrގ��o$ �Jw;>N�[�==���8�GC�,��:?I����l끗`\ȓg��9����tg��;�)i�$�=w�����Y��w:t����;�vnㆽǎ�<m���I���yػ&Kw���>���f�m��.���ո�`�6���O��z��w�
pKt��K�������e-$i/��Ň��R���}�H�-�s$$���ɛ�xKc��c��rv^�s��@K���#k6�m�$�����&U�>db��37
�/��DO��߷���ƍ�9V^�����rtO���M6|��<�N˘X\1tZl����x2���nOl8R |�o�u�!�I#s[RT�)GM��@��F]��]�k �cT��ٰK8gn��ɰ���gF̳l���wa�?�.�_y�c9aeh�l�gy!� <0 �FG���m�|�|��=6rp ��]|�!��2��+@>@ �:�!:��a|0�G���\9qvҘ`ϐQ�� '�O���o'	���>A�aݓ��!����  aE,4��)d9`�W7o  �|��P � ��$��{� �D�p3ǈQ�!��7�� _#7�( t��m���^����  (����` i�]U\��@c ǧʀ�#�6�8��v�*��c�!uV���X;���0��3}l��մ���/W̅��&�%9�_�L�_�,����.�^���o�跻ʔ�ϓ��)�G��&O�
%��ch�kv�|�v�Y(�j���k95gf������`�����yO�ۊ}ܛ�>��+9��VX����>�,���ӧɐHzO�V���=p�z��{+<�� �nX���>�$>P��,�X�����/�֥ȰW,�K"B3�>�"CWjXh���s����̈́^�igs�xW����֦Y����K/��[���ZT�X[�Z�k=�1�櫌+��i�n������L�>A�ˤ>W�O���jin::�~�X�%����t�����Z�8掌��]�����4��3	{ B˒Q�d��:%���w�179&웲wl^�Ve���M�E�;�p��x�F^���� ,�$
9�����%^jk�d���g ���^��'�0���U��P1r��fY����g� �(����H1�%:�Y�R�Ly'{'=0� �C�(��;}�Ffl &Ηb\��� �%ٗ!�s��p>A�� 1�1�2<� �`��NL\�z�x�>�%���3 5_��� �"���vw{�X?�e�·%�h�Anf,�il �1�ay�+x�'
�lrp�>����|�Ʉ ����ѳ�	N0��ۋޛ�f=��}�FM��Z᩾r@ 
0 %<��^i�zCl	$6�og<�{���� Ng��O�x��H$ �0~�-�ќ䏳�Ζrt���S~�� �|�`ɒy�  �!��    � ѭl3����ã �  �f��L������7�!�	�&ޝ�щV�*l��H�x��y6|���0 ��2�l  �6@ h�0�{���7Ѯ�9%���fd�py�m0{���@>A�NN� <?d�`�  0i���d����w������Ӥ���|I$��0 }\�f��� H80�2���� �|z�i   ��!����L�S17�� c>� { 2��Q�9ǜs�[���H2�z��q�8:>��'|�{�� rɻ&� .R��vM>�@�ܰ��`ǿ�0K�8%_�`?d������y�{^� ���@!v0M�U�2vE�4`  p` %�# ��`����`�$&��P)N�?Va����Xc��dׄV���� ��L�EN�T�N�>#�/9bu�G� �={��S��txw�=����Hs�>���2OLR{��-ˇ6d7G-�烞�n{���[ds5\8|�Ɠ����{ �y���#|�P��̲�:9��5���ȓ����9��{|���M�#����+N�:���&|<c!m�@�@ =n�0���|粒�)�.7Hh�}{��쓌`��Yi�'�A��3r� ��*O�' �d���c����>�9`v��I]����ن���O���#��y#��� �?�I�e�����k����x�����f�s<p�}:xy�����0�ܒ	V�0{1w��z\|�0�|y(�:��̐|��$������[�[S!;�"�r6{���ˎ���4�M<s,-��w��>V��9��d ���ž����%���������|���Xuv�����ٸҦy�	s�0�0mbO��^b����[�Ӭ��Z�5�n;ơ8���ϰ�ur,s�˕�q����G֮�6�+�#�Г>���aOf��hX+���̪60��ӂ�!���Yh}2�4�gb���>F5�Ⱦ�
���@���Hڊ@����b���9��>K���S�]���q�e�9Z��n��B�-�b��2:՜abZm����2�v�
[U�Е��Y�v-F�cۭ�b>�*���J����=���	B�B�qɅ��+f�*5(E�U]o�j��1�L��)*(�'R���uۋL<É�Y�Ͱ�W	1 ���aLl���$:�kL4���0mГ���r����`�F���s��+h��c��Uh�����v��O3݅i�R�e
\�.����+�U�9��2�*d��^dq/%�k��:*c��Kr��r8�r%ĸ�wE�(�K�2��r�J��FL[0B��b+f8YE�Z�e"fae�.�[�oFkF���b�VGg�^�Y�RA,r��PE[fjB����Z�wwB�anJoEi�DC��GuRS����S9ec m-ZI3MHL�ꤝM�V�Մ�eoY� J��2Hy��'=RI���m$��ݠKI���,`�����:k���z���hI��	u¯�䀞tXД{v#�̨ʁ��3t�o�Hq��L��LXy�u�5�x@�0-��ɦK�S8���%'̓�;��N��T/��'�RN!1�$�B�I>g{R����$Ć�o���a�P��R��c���<��Uk��8�	���V ���i�BZշ ؿ���b7��k���ξ�OC�`�0茪dF�KJ ~o�k[����~z�X�Uz���������Ҫڮ�Uz���Ҫڮ�V�v��U⴪��*��b��WJ�U^,]U**��*�����Ut��V�U괪�U�U�_Q
�*��d XB��I"�
�  �"����TTdQ���T��[Uګ�V�t��V�U�"��|�U^�*��*��b��V�Uz���ҫ�VեUz�����U�]�N�J�*��]*�V�v����Wj�����Um_��@XHu �$� � X�Jm$"� ��XQ@���g�H|}��{[ګեUx��V�v��U�]*�UUQz��������������V�U�UҪ�b���UW�J����j�j�UW��UU�Uz���եU^�*����� �$)X(�RAc�Rg�7�ff*������եUx��V�v��U⮕W��U^+J��R�U��U_"���*��t��U��U_"���m�U^�*��*��*��*��*��*����ﾐ�>�$ 	YT@E��)$� ��6�- �/�B@��$dTׁÐ�*�������WG����@6���y��9/�i��6��-��V��[�ukX�:pK ��"lDD��GH"A(DЈ� ����bhM��Bh��$,DD�(A(DK�,�<��F�؛blК���h���$8"%����b4&�x:C����<�� ��"%��<"xN�%�(J ��AN�DК4"lM	���?�u~�����Ֆ4O�tD�5�q�>����H�m�qF����+ZtG�QC���YZ�6Y'^a�#�둲�B�d�i�lVR�h;*��h�6Vݰ����X�PUJӮ2)#����f0��,j±�1Ҩ���UUq���+l��1�,���M��N��?�\�l�����(��::�
�]�G�
��L�v�#q_������Ls��@�V��aT
۪)?��eEt���Kei�V ����ڃR
C�K%q����N��񄨉�WK+�V؂I\�����U�FS�dc���S�7�i��@��*?c���Ye+k�J	��!�q@�*B�pn�k����c�J�E�6JȞ:@j�'aX�
۵��?ek1�ʛ��J7H�uTA�?س0�NI~pv�1��r�SJ�	*���Sn)�� D	�<�ʲ�[������ �"�F��#�D�I��ǎ8Q:��"D}kM�	ba�dbn� Ӡ�G���X�+v��+>m@"�_�����X|���+	Pu�E�Ϩ|H����2<rH(�+(Z�>s�"��J�RY(ڕ(�*��x�E�����Zܖ)eBj��	]v8�"�r6��lX�>�[�:(�B�-V��%�j;Ɔ�ݖ�\��1 �(�Li9�J�1�/��d���E	]E��k����k���nF��Dթ�T��N�����ۑ�Ȁ�q��]��+R���c�R'�q|K�9~��,�8⮳�Y̊����ڶEm���&UD@���>�y�bm�ƖET>�PڲϜ,�N��b��i�UDv�~�ʬD��~jʯ�W!�n��n�R�n�D6�R~nb&X씊�0uʢp$�Е�Z�j([r��*Z�e�J�P�d��e�b+�w*yaD�u[%�����H�m���#-�.��by�,�M�ٱҴ*RT�e��lu��$��x\h��ّ:A�Yh�Q��j��QbrV�U�m�����i��n��~u"�`�(#��X8BA���D�r�v�>R�A+]��AK��-U?�����Ԭ��R�K�Ue���L��'�<L`�GF	�D�'�WJ��RѺ8�*���	*���E���-��j���Wh�d!+��D����E$RUH�� �mT����H�WUt &�>�U؜���qH��##�U�V2&|WTl��g�7n���l3?U���}~��8���T���}#E����Z(傑��R6ӑؠX�'没��C���3�U��ײƲdR�Fm<�e1('1�?��8%]�Z������MF�C�c�� ��'��Ѧ0Er�h�����B�)d$p����Tn"Ƭ#m�A�+Y]�r6���h�|ʸ�!��m)��v1��5C	18������n�� �l�6�Z�-NJ�L��q�Z8�'��ǃ@+��j�����V�T��u�ƈ��(� ���T���[mh�����V������[%�A۩���U���&��~���_�f(��wwk��|a�����*�����ffffb��wwv�|}�ffff(��wwk���*���㍶�1պ���Qqj��^~�H�!�m�rإPjWP7%j�����)*t��M���G]r:(�-M����M�E!S��2 �F��G$��~��X
Pq�厊�l�Q�D�#d�VҺ�}V�2�X��i��EYX }���YJ �PRY],�JY%a**��U�WK~�+ce�φB��Qʥ�lb`�n
�b��Q�5# Q���Z�m(�en�7"n��C�)#�ZGA�9(ҒGY�	�K���-QX�ɶ����IpN���F�QEjV���Wj�E���i�ڔ��#�&�T��t "��?��~���}��[�fY�r���;����V���ǯW&�fq������Θ��s)7{��b�oc';{���gȿ�Z��74Ťŧa��o������2K���UU0�����[��;g���|���p�jT�}7����Ubhf
�'��3��1<�ی��[�j�pF�R���ϧ�TG����e*~���۫c�un-Ӯ���yr?uԒIR���a�o,�n����U� �>�"��2������Os�gf��*�����5�P߇��t�F�L*����*N��ku�J.r''MNo(�zl٬[��aӮ:㭶�un�źu�q��+ն�UY�^�Z�V��+!ۚ�~��;��껨|l��
0O�d.M(��C�u�L2��F5�>6nm��֩s+I�c��\�8v`�X��.�Ro�[���á�_!�p��NN�^��P����R��ӥ×yR�^��k*ۦ�cL~q����[�q�Ӣp�f���F��m�|UYѭ��w�.n|�溱=� �h���x�@��]Ça�]�p�h��P��0���pW�g�t6p����K�쫻�p�2a�-�]��76a���P��J�d.T��h��6x�㧎�8x�t�6X�zU�0�̤�m>=7#.�f�"���zX�qr�$�1Z���O�n��"-��J������cu��Y�=����ջ�c�{:}�ƥ�r��j��-�C���'gQ���sof�ܯ�R.�}�{{�Ӝ�M�M���C&*九�bϐ�sʩ�ή}�j����sYt0�3��5��&�|d�~U�Ȓ�t�F���(�ў��ʁ�%���v&C��Y7\�%�	�H*r�C�6s��&h�Л��?S����6��V��[�WP��E�Á���u�9�q��u��~�-���{����Uտ�TK�˫9�«,�cD�D�kf!S��p�0ЙĽX��6�%�;XS�;��k���O�������텼�WyI|,mu
�IR����iǫc��[�un�źu�\Z��r͹n+��wfY���5e��C�qw20��0�Ӿށ5�xa������.d�a���ī)ʁ?ollMG�AX�#j�~\�w�|���}���݊/��%�hvh�����ܣ"�-J4\��+�(V��	'��oŸ�n:�V��[�]G�X�����Bϓ���P٨m4�8��v���P�٩މ���r5CP��¦�a��̢�y��Po=�IE��<��ǟ7��|��<<ha�'L�>�S%������Z�m�X��[�t��oO��6�����}�D�& ����>5��2��U����6ڍDҜU��K>i�  ��({�=��8���s������vY˼��ARƷ�����wu�s�"�\o�b>��OX���$�����y�֛w]��Q(�����EC�Wé�\Y*P��=�K���I�C-ƞ�����}�æP��g�p���f���˄�7>,���R`l=�)߅��}q�x�ʃ�T2�,p�ç�u��un�ո�N��6�i+)UY7(�d�(��g�5<r\ó�f���;�][iE4�,�0��p;��O�ŧ$����]�ϔM,HB�C�xF)ݵ|ےB������ﺨ�CP�L�;Ԟ�<jU�OvOiEV�e��ɣ��|ƝLJ�V�-��x�&���������%��GS�~y���Ǎc���b�����Z�>G�4�>k��112M���b�����c��vO�~N�|�����)'�x��;������N��kkI���5������jKL&L�G�J�d�L,������Xר���:��1*1�ORI1�'�1�N&#�6����bW�cm4���jOR��wS�cƱ11�y:ǘ����mjcQ�bcƱ�����'Y�1�������?'�cH�J�H�M���bD�#&IQ�m+I���������2O�`�{�U2���p��9�|{,�iә�{���O�ʵ��i"{w�ۡ7���f/ܗ���,R'5�o��_��&/���-s9W��q3x���?jW(�>����(�����}�}�Js���]�{ڵ�d����c�f.���\ ̙����p����{ڸ|fL����s&fg�}����m�q�1��ո�O��!�͘0�$�%ޱj��%�g+���-�R�!�980+���50
'�0�a��mb��"� �M�͖D0Cs�������ΓŢ�.Gg��fA���hNQ��.p���(�UW/�������3,�
;2�`�l�2C�&�_�橦��Гƾ����n� ���5%v?��(�C�."`��U�&��`�
4|p����e�q�m՘���zӟw�.{�/]ǳ�\u�;�UU�X�JQ�,�'ǮKD��`Jd��}S�0�m޵�&ɫAeCh�Cp��&�0�&�F"!i!���BZ`��D��O����|:2xd�0<!ힲd��5W$�������8Xw0J�u&-n,n_��Q�d��s%CC�d*%2v'�j�J�m��!�+�4�4~uE*n2����
`�&�!)��*�+�m�_�c���έ�tO��Ǆ��~7��toTd֙���4�ʾ��~9��C�����7�~x��d�J�T�G�1���8����!���4٘K����uX��Λ���wf�.��Rmw8p�qkP��I��5{���n�k��fY����_{I�U��4_a�%7u'��*�E2`���D��P6wVu(a;:]��Ji>��p@�`�Ё��*C"D��*���O+$|J0e�P��0�F��؆��z�|
W��������BlH�l�i=;
�B��HS��Eva�dR�;��hH#'�I�I�I� 1��]��N����A�ah�HX2j \`P�� � z,�GܽO���q��>[o�>un��Ӂ��p�fsڻ���d\�y���UTj�R5A�%V�T��ċ	�ϊ�5F ���' �.	ibT&	�І 	P`r%��P`�'(�3pd����11��K�_'�	�Z�@��؆��Y!GD/I"�ި)�z��I��a�g�l��O|*�(0I�v��=J�o��&�T*MP�H@�F	!qu{.L�j$� ��",��Q�2"%:����ͺ��Z�[�]a8l�2Jߥ��qL����`<AJ�]~V�'Sq�2�Lȓ�2	'��R��%X�g:�A�&&����a;,�hC"K,1�d~�0DJOB�.��d�%<�
AE�TK&.��V�b�Q�)�Ub�X�WIU��h�V��:��IQK-E[��F�\O�Ϛ��L�~C��m�n��O�Z���ǭS�

�T!�Щ�2'D��!p�lԩ4&2hB�щD��8�UlT�-KO�&�VjP��]4_�UZKdR\L�C'�of�?����Z���:�uǯk���a����:} ~��.�t[>>t����'5��s;psT�������l����4QbdL� DC'��q�`�XrlA���U+�O2�-W��᎜��l�\��$��T�߫���M���S7�&��CB`��A��
�R)���c��J,�2Hj���"˪̒j��U\
�CC!� pC�{��Wm5i��6�s���Q��.2\B�C&2�@���ţ�I���*!�=:!�@��1����9YZ8���cn��Z�[�Ç�pك�� ��/�CZ�)`��]U�!uMi��S�ש�R��p#�ӆ�V�m��J����n*��n����m�e����/&s3�x;:���9�Ƿ���3����W{3׾�ꍧ8�5����y	ݿ�߷��^]U7f8Y����U�Ã�@��2t
2 c5Ԅż.��G>&����(��'���CBCl,a����F0�p�K�B��:�KX����p�W(�*�:!t�U��h�6}
dd�+-��4!Q�da���j\bpds�}�Q��>6;ҵ�Y4	L��l�����a˪�O[Y�GL��ȫW?� ���v}
?J?q�rS%�p�
2F><T�c��׏��o��խn-Ӯ�t���:pZ2�8��S��̎/E�����UTJ�49��	�T�A��S���Y�59�Q[��0� �(n��k٘D]���a��SR���&�ʑ��0�2zQA����(�/ղD�R0a�O�P�}���S*��#.+��!ᐐ���^����4'��Q���!��ц0(e�CFE:\�`�%0���>{YR��Z�RU[�θ���c�H��<<C6_g/S*J�t�I��UUTC�vm�ca��T�@�;(n�`���J��
4��OC��rR~��)A����!�R,�eI�B�Pևe����:!}���֯[ػ�,�Uam-X�z��['�,a�9��l���eE%�r��n�s���T\���6!����%0��%!ʕ\��5�{o��e�6V��1.�K��2hC�Ct�u��E�RRtd�j�;��\4 �i���`����İD�=[��c��c�Z�[�]F:�������ڪ��Q���%Q�H��X"��<JVRQ�2U4ރHeϺ�a��lϖ�F����I.!~�0?A	�Ý=0�`j	%0�*()����	FJC�[���` ���RCB~i��V��d�iU݀lN�\���04 l��MB�K�Vk

���%��ap�4!-
 SիXh�KDt�(��bǅ�|덢�MV���q�N�䴮�����L[X��LKLLG�Ķ5�ljӮ4��D��ǌy������bZc�i#��bW�k'�Mbb1Ʊ+���lj�7&1��4�d�$�>&	d�!�<Od���:��1�Lm�#	�k�5���+�d�Q�
8aVL4^��%V$�~2%�	�,��,�0"O�ت�g�D���hF�ƫ��N&%q֫m4���#���+�:��S�jc]b�bz���&�ĉ����Ʊ6Ʊ1z���c�6ƶ���bD�VT�"��z��0J�|8'�0��������(�n�k��O�k�uǯ��,�	��)�ԫ�A�]���%���mߦɋ�st�sK�*_����M�p������zϯ�����`na��Q0m����M�e¯��[�����{s����ֱu�}�Fr'�{�5���=�˼_��}��߱~W�%�r��	�{�*8Ny�ՙUh�J�<l�˗nV��9�I+?nFSfi2n�o�-��غ����>�f�Ԉ@�d�?�LP�7P������B�D�����K[�:�����ՙ-w"�V��Zƈ��D"�(���kHq�N)��~B^��+rJ���}z���Ϲw333~�﹙ڬ��fffub�����g�32�333�s�wy��̬�����\���fx,�N:u��:��źu�q�=~n#� c+l`J���"���� ���B���6";>w�q�,��ב$d�,���݂�;\��pd���ǖ<���T��CR�J|�bv9�Zɗ%������JZ�m�C��Y
�n4�%�U��:ꐬ(W+���e�Q�Y~�"eʬȨ����XYT�X���b�F�i�A[Su�Wie�W�ES��;o�J��*i1ʇH:dx��D|F��QO��0��(T3SY.:�t>�$�&�T��0���1xl�7�Ub�>~�m����������u���ys������Y�r���\T����}q��ÑrsWÛ޻�x�tx�i��{Z���ڿ�V���am�e�Zo3Z4n|	��.l�P����|"�X��A!I�!_���,�����0��a��F�RP͈Y�R���P�3�T���O"Pg_R��Z�d�9%OD,aߧ��)P8!u���в�%=�M�u��m�2�U�S��pBxO؆�Y>��.'�yF/~6�O;�kf.Yd�̏7�L�'�>Qg��\?���'�B��E�9
.Y��<Q�����1o�b���:�8����<��$Ǯ� �n��ͪ���TJ?D�����d�X�H���� �gbr0؇�~���fWܼ	���.	4\(�\�>�%�X2"&m�Q_����6Y�L�y�wE�!����ȝR\`�Q����Y�W�V�-��F����	�aA�Ag�d�a{Nk���j�=�O�F�� �մx�՘h��*�4x����-n-Ӯ��q��ߒɋ�8�UUH�`K�G�CF�/�ʺ�5
���f�h:$6aPRr�N60��ߗ�vB�|����۱J���:�9�B��t4d�h�������ݪb\�nϲ�ܻi�[pp��X��������'=��_�i{����r��¡�\0CH(Da�0�l�?Mhd(B�U(��h20C���d1��P!�"��n���Z�nj*��������V�SQ5Hi�jߛz�����lZ�[��l�كգCS�UUT�r����yх����Ða�Aa�*\���a٢��_�u��:o6̿�d?�f�3�*�x�9E�~Z}��uUF�ǥ��x�� ĝ8�P�`x�1�ɅA��r�,B�ڡ4&��ܹ��-�3�������v��a��C&��n&�_�q����ZW�jڪ��˟���~��;?B�Ü�W�UC]<���_��z�X�|�lZ�[�]G�׾�vz�{���'���P��pT�ǖV�0 Q������Q	m�g3/�m��hJ-8��v�T�3�s9��Ӽ�ٝ�1`�fɵZ�8�dx�*�l��]9�n^헙��p�7oX�꺲�_n��g��
�>aҪ'�t/&���C���Q>1R��y�pCpd�Y*P������㇅��ٸ0�~°��U4XdB�ͦ�4*w�h�jX�z��Ӂ�]M��ˆ��d�Sb�}i7�MCs!H�e��;��r��������K���O��0����K�a�,������\�)���ۏ���qվ[����0�]�Go�{��޳ޱ�ꮾ��rS�����ٲ� s�3��r?a��-\���{��M�'�l^�os�^]<��\/����/{ͨ�Y��~��t�p�JF�z.*.��Ms�}�o;7�ӳ��0�l|�\�<7�M�NC��ڪ@�Vi��*�pyM��!�Uk�H�����]=���	b���3��Z�"�K8���E7MuZ�
��0�IA�����5J���B�
������0��J��/�T��U̬��t>Q�x����na0��MR�pف�0>�����,٨T7B>��
��75�%Cb�5�p�0��z�����~[[-�c�t��E�3���3��/:ڪ��`��F���b�c4�WCD�XĠ��djYXX�6`P���T>=K���p��aA����K�O������a��Ï͈�:aR��F&�+�W�B�ϡg־6K|���$��Ĭ0*!���@����V�̿F�ud����9�5��z�ƴ>�Ǐ����)A6(��!�:fdg�\4��:�;qk|�1�1Ӯ������y��$��UUT�sRn�I�]ݹ��"���8ьOL{�o���;<Pn�o��f���E�"��8��ѳ{+5���Y���!|q��E���e����7������:�A��G!�)����w)�O��#��9Q���Pt�.:]��q9wP�?N��u�i���έŭ���8�N���>+,��3I�&q�E-?2�|�S����u&U�~y�1&�ا��!���3z�m��o8<Oן���:'�˳V�;��g���k�t�~��z�{gJ�f�wݹ�ۘ���8[��׳��*��s$�ư��|�����!��T�����IA���8�??7hx~���.�M���]h�\��w���,�&7�(�ؿ�\W�q�#�ʗU������E����ҡ�:���ϊ(6Ұ����i�#����reRI�YrA�0_�_���Oi��?x���i����|��ű�q��um����Rk_J�������UU 4J�Z�j�<w������2&B�����=�2A��ga��;=>�`X����Ew�tl����hș�L�n	��a��MT,�^v5R�����ٙ-�u�Y���]��e��5(�}�h�&��2c�r�ɰ��_�O�����n��oi��G��=b=O�i�Ԯ�i�|��[LKH���-�ƭ�-�-�b[����D�c�bcmbbbbZgH���LOS��bm11�V�$�4�&��cL~i����c�H�bf��1�S�k��%�?5���bx��>O�|���1>O���f4�J�rO�	�C�#�ğ	�l�O��M�Lj�x�I���H��b:��������bV�	�ŉ�h�!�g��I��澓��Z���c��&'����b8�cX��LԖ�����4�bm��ʓ��2I��bD�1���#H�b1=JǭW�i�d��w���=/�{����M�lfy�sa��L���r��T�t�������w�ƴ���g2z�.���ϭ��o���N;��_��U���hlOxq��w�g=�\+ը���k�ݷ�&����y�+J��r��33*��o9wy����W�ҷ������J��i[�]�fv�t��~q�1�c�:�8��Ԛ�b��UUH.�E��IfCghCz� ~jLh��%7F��'��(��s�K�e�'���֨�Z՚�9���0�)`��t�����Z���f�Z��GC��j�p����?�YuYbe�V��æ�6p(����{E�kЬ0��_>[�͸��[���Q��o˛�{.|���j=FJ�}���4|(�.aaA��J|�s�EV��R&��e3���l;��w�����E��Ջ�>�O݇"p>�Z�J�������F��D��1�~Bs���u�yX�.�s�aA�υ=�٧9N7O�+u���8�V��[屆0�x��4w��9���Ww�ޏ:�w33ǟe�b����x�������>�L���j1�9���5�D�h�p��UUR�3��Bޝ����1�7Z�"~7,��z�p����[�X��.��]��)�
�VG�;�7[is�u�>0o9K>���8f�������zh?�X�h�Eeʈ!EH~�8�>��������vdXd��L5H�Y�+*۸�r#7~�4p�e�u���]>ϵt�g��6��[|Ÿ�1�1�u�-h�oNMa7��C9|��\��e�UUH��醡���Xg��Xl�<\��T����(�T���_��4c�l���#Gi X�?��Vh���0�^����XX{��cٯ�3/0������NCG����4XvQp�L���ʜ��,D2����ƚ[|��:�1��e�!�E��v�9���:���T�)�V0���,��ܣ�w�n3���0��<o!�D3��2���*�^[m
�h�;-�ϕ�w��d���90����UZ�S����X{{�_���O�:��C��ύ�k���!�C~��Wv-���c��>q��#Ǧ%4���??:��-�a�0A8h�]�W}���ݹ���w[�˙�+Y̻���͏�I7is;oXwx�9�9>UURFg�}=��Hz6"��Q�(��5�w ���˄�ݷC\����+t_ؒ�E���:噳tl�h�X!���*>7A2l4�⒪��cu�!3�x�������[k���l�"SB��_?>z��\qվ[�:Ŗ�u��Z�U�nS��wV���%W0�3��K��ߖ��鎚s2�&��lQ���j�uW:򪪐3}Ύo�X�ݝ�.���cQ�������NN���~.��'�9:���k��{S�}��;�'����&.��W�q�lϾ��[�44�C��*CSի+G�cr�uY��l5PN����W����4�%^�5��v�t�9FHK�U�ZY'�BI���+B�F�x�4e��Dk��(ƌ]Y ��ćء9O����J8z�r�5CGwFh��&�}~�.^����=�]������g��h�5]/*�x���۳�&�M����V��0��"C��e\�J��UU��M��}�0n�$>,h�t`�!��6cПd�<h���FOC!��b]C�a���,��9�����|5����=��o�,M�~��o�ғ4NQ],�Z�羂��_֕7<]�"T�<Y��틳�%k++o�V߹N��z����l����m-m��:�-�cb�Z4Yf=���ꪫI�e�v5UW�jl��&��y�h�r�O�ڃ�=k���s�X��ȧ��43���Q^˼�f���8j~�u0F��Sz	���U����;C�fº������GE�OO�Y.:Q�(Ҩ���x���u������^#�q����8���[�:��Q��{_�L��<��K�I�I!uZ��nG�+:4A?D�j|qS�ѡ,���6Q_
uh���'N��XT0���NLEZ2�e���l�2 �%R#�W�ϙт�=Fˣe]]`,�������ۿ��{7�ͻ��"ۻ�>�w�~�q���(��H\<aB�"��P�g�a�ك6wj���ޚ*~�-������b�u�1<[X��KcV�LcKLL[X��Zu?&lk�&�1��1�bu6���i�LOS����b��b-�Z6ƌMɍ=cOɉ�=F=j����bzƱ1ƺƣ��ʣ
ʒ��L�(�a3�V$J�Ʊ֫rc_�����<c~I�{'�d��J�cO�$'�"|?"BI1"1"VI��5�|���q-����'��!��O%�ćG��~����>8?3������<��?5���3���1���|�[��W��0�#ʒV$F�%�%i��&�d���~M*�&�!b?"��w�N��ع&��g��+�?7����t���k��>� �E��)�T��d'Lr���ڮW�Z �\`�n�q�8�ΑsnsA8<Z��}���-�>�,::�}����<5��}E��ӝ�w�0�f,�f8|_�Ӛ���v�{��Z�{S��T���:�y�E�mq�˵k�*���՘֔�C�UZ�]��՜����̞pߵI��s@b�0XY�&�U-l�%��%F�Q��c>ꪎ�$�ҹ(�eS i��UJH�y-\t-mI� e�W$,N�Tr��x\�������I�e�pi�k3<��n���331ګjҷywy����U�]-�r�333�����ٿ߳3�m��8�c�1��u�.,Qg�o���}$r��V�j�$M����,��EE>tj�
��������?�
�b�TX����Ҧ�IZ��A�~�Q�Q
��������m!���i�$M��R+��r,����T�Q�HݎKh�jT�n��QEZ���mߝE��W�򉯚��!$-�Ws0�Y&8�+�8�j�h�L�.$9`8╊4�T�cu�:�N�hPu�����냒3��C�V$*��)KA�$�S�U�(hd�`�KU����X����6�lJ������5km�ۉ��5	j���|dH��T	؛p�l��J��d�Y#+����m��B%�ו��y����unOVN���Y��̽.{�Sy���79�X.󓯱Aa�[���X�ȹ��]���W�ĸ��*K���Bi���~�X���CxhI�+ۅ�<ks�h��v�B����嵪�f�����n�BL���q^���NV�Կ�*�wf�
0F\�l��h�;�L4��&9w�6C%�bp�e��S��Y�E�6t��O��b��X�]G�<{�i��y{UUi �`�w��!���	F~'MQ�ר��@��ȭ�F�4�%v�_�����K�d(D�Ҍ?l��粽y`%��\�r>�`�{7o�+0�;p���@��}߾���3�=Ŝ.&C�(��a���9zQNF�{��G[un�q�|�lc�uӮ���)�}�ɩ�>�r�;���	P}�+�q�YꪫIQ���[$����X%��A���Yr�vX�(�j|����P��/~Xc�yVB(���=�m�]��WW URh^`p��IU���uQpr�V�K0&M�9��~�K���a&ψ����?uEY�%�c�TA!��K��z�8�ž|�1�:��Q�%��x��#x�UZH]�$�ѓ�u�]R���E��;�{+�@��Ϲ�X����kqQ�	8v�#��f\��t�?���ĸx�T=�Y��B�C!�B'\?a�p�Y4�~�m蔚�Z4h�U��!�V*���p�0�?_⪌���ֱ]��ɼ�2$����'k'
��F�2�{ߞ����X��la�Ӈ�l�fk�BFQ�3V�������V&k���R�����Qp&G\��
�]Q3�+ζ�m������~�����չwc�K�����	���!�'��l�ڶ�?y��rnV�={�|P̌��pܾi�T�;U1�}�Y�a�(����u4Si_b?�H�ͣ�i�m=l���n
�TC^\8eP�dO�'k�U�r6p�V'K���Q���<�Raɽ�0Dn���_��UC�:l��;0�8%�}*�b�*�٫��Z����r��n�!b�0�5�5��x��	꘬�F��^4�>r�|��|��>[ź�p��,ˆ�=�9��w�O7��������o-|���0V�����w3��dוUZHz��f(�v�A�fh�4��'�0����I0j�>�v�o�G]�~m}M6�)��i�>�rLѬס ��)��a���bn�G/�0��y,��cѝqxqm�>��ڊ�tY�?�?BϏ����?HNB����A�G�����\��~���{!>x�~F;R�W�����c=|�n-���1�]:�8�ǿ�'��h����j���CUo[m���O�O�0��{kjɣ!�2r%	���WC{3�y�h�pO�T�̇��/G߮�n��E,E)�lÇ5>���S$�O�a`jxE�"Zl��G��f�g���˙?{���)���Mӓe]u��SOk��s�q�n|��c屋u��l�e��.�UZHg�B]{Z����t��g�Н!��Yth��;��ؼ.!����K���dɖ�r)G7�����*�+�p�4k��}��g8n^"0��WqUW�/
����EPwYf����Mp�6"&�ea����(F��/�	��L,�����|���ȶ������J����]|��q��[�]t��o���<v5�������^;�^?�����vh��ύ��9�\�Y��ӈVuw���(�'��T(kZ���UV����s��q�s�y3�8u>a���|��g��=_�۾�A;Ǚ���o,��������]���6l������7�k����|����{�o���D�I�\w���%db��|}SO�'�&	�p�svh�e�0K��F�:�##>�F��|Y�>�eO����M�˷�M�6Y\=�8#��`�\4hd��$��4\(�;w�*�r���m�10��2�?yw������Iʿ�}���"�-�qk|�0鳇��4Y.w�.��UZH@:��hL����HJ:m�Q�㡒_~�����ˇ�w�O���SƄ�����M�����,Н)���	V��p���âgؘ�촿�3�K[b���1�6��jp�s��'ŕ>�����,K�D�w�S!�pD9j�!��W�|��ߖ㎸�V��[�u���'��NA4"'"tЂ$4"l���6"���M��6&�	��DM���:hM�D�"l����xN2X�blM�6�e��(�Dd�!�|��BxK(�GE����Qg]cz�1���<``�DM����pDO�%�(AAD�d�6&�ؙ����uK�9¹�����7���yM� yy�۰O�ͯ�Y���[�o���L�\�q��6�9�r�7��NG��o��_.�'\���͝[,��!ׯ��k�]�^~��z�7��k3c}�<�;+�t�xZ���@�����T��;��8��z�w�n3OnR��E��
uU����xS01�E#����QO�}�;G���� ��׷�Ϋ�Ã��tm]��9���t��~��Uߺrn��z��D��(�8Si���KW+��GV{=��ǯJ�ld^�j�g�
�^�w��S�v�'q�'x������d\�f�9��G��gy��9�]�7,�k��p�.����&\Rxۼ��=c3�b>$J͑y]~�k8�M��L}w6p�`�?��.\g�3��}�[�7�QŖ��y�>57��ƀ��]Fl�����ؾ��*����s��f̯�G�'s2���g�ﳏ�^�灢��<��������9ҙ�Ungz����������3o�{y��t�;�כ�.�׿F�ੵ�M��^Yf��^���Q��s�2c|��fn.��k��7�{ͼ��V���ust�޷��9��u���U���]�fffmU�]-���fffcj�U���]�fff6��Wm��^fnΜ8p�Ӈ�-�[���:Ӎ�Ni	���iUZHk8v�۶�&��rJ,IDJ�/���ͩF��2b0��.��&�.���%M��U����mG,Z�/nZ����ѓ$&�JH�p�������-�P�B�6kƃP�sF	��+
4N(��'��n���~;��Z;�zO�?>cn-��-�]ui��=���2��x��������/T,�ԩ�rp��3���&\���T��Qw����CF����.n}�`�%빠Љ���}k���v<�e��<>F���O�蝛8tJ(�X��,M�й����=���B�׏+�=cc�ֵ�[��u�t���;���ZB���жb\F7m�F+7���{wZ�	�j2�͊��Z
�q8���B(!g��m��B���6q�G��{}�t��]�q����s��w�r�]|h�3�g�-]<��=;��ĩ�l��;�{/��a'��WńQ�ـ0��˩)��q?"h~�W~�.nT�V���'0}B�MK��>;&���[8r?	�:Qΐ���L���X��V7�K�MMM�,{��DOߖ����	ºh藞�E���uM�]�a�ʓ!E	���x�_E��><�6����>[��u�u�x��3:�K�s�`�,�6���A��>�?7.7e�g�A��4`��}�T�a)��,M�GC%��+C��C�d��>�&ˇ!�`��{ß����9=54A$���_�#e������y3�v}N���a��N��r��`�5��p���ʽ�ܟV���۬[�-��]GJ8l���6g����o6k�S�1��Vq�';f�G����m�Ј`Uu�IB_����/	Ȕ"W����2���5
7""��v?	�7��K��L`e��ב���%�K�G(a�ݞ,MP�W>���2_f����vlON#B������П�j������A�!��5c��խ�|�ͭo��1oκ�:ӋTQƹ����r���ٿg9>��X���ݛ��՗W��|n=�<n�{��V����UV�X5U����'�Gk��0L�EN~=�Â'��ڿ�j�4�U{�����أ���f�XlNyTF�bL��ɚ�����;FF�h�ŉ��P�h�CT|&�H��=�v�j���OM�|3P��J3��'!�໛��B�U\�c=[n:��ul[�[u�u�x�ފ3���*,LQ��Y�>�v}��0��j1[��X�?6�m���[�O�M��uo��-�[�����5�a��]圕��3y�/�&�W��߿j,r�ϽY&v��s*l��Gy^r�|T�C�����F���Y�y��̨�VDr������i�?S+O+����i�T��'�d8^͖%������K3��~����'x����գ�\�6hJ�
����e	fO���~�E����F�M"gEQM�����3+2��Ӑ�&	���}��Tkf���ض���[�_�ui��wǫ��K�Gƫ:�5kf��UV�(�C��,K�,�p���N�������"jP�p�}�,Ќ�:&4b)�:u��!�C�2v����qv�*���T�Rn{x(X�����*jJ��\DNLֵ�*�W�z��?>m�[�-��]��-Q?غ��Z2T둑���bT��UU���VH�Q.�Gj�X�l����j&�	�:Tl��$>Ѯt��n��:l��_`Ho�-�ob�ee���r��e���h�D��}s�T}9\>��Ƅ捪���ҏj#��l���P��^6ݴ]��
2j\:aن��.~���=F���mo�ű�u��Q֛4Yx"����UV�Q�,�D�j�z�!Q��I��=�))Fkw�(��32����C��vD��J��YsAE�x������h�|z~�OT4������q�ǎ/I����w������S[�$착�C'�Θ}�mI�8��:�|�qkun��tO"'���� ��(D�f� ��b"tA<X��4&�١4A""lDD��B����lD���<��,M��6&�	�e��(����(�|��Bx���'D�ǫz��z�:��b������c��[k[�[�[�6��f�AA�6hK,N�C�����R{n���/w�����Bo.d�."f�O���V�`��hTx��q��Nn��,i���:�����N�O�<���L�ȘV�r|#[_{Mˤ�py�q���*}-s�(�lɓ\fnw!�e]�9����mnd��v�< L�ae�[��T�n�\֮�x����n�ty���9�q��ssY�d��G�d��u4�V�f8W+*h�=�n@ev����Б��#���~#\��C(Ԁ�'O��(ӕ*A���t�*V����M�A��l9lwb�E�*��/wS�׈kW���mU�ww��������Wm��^ffff<WJ�ۻ������x��]�w{�̳�,�Æa�a�x�ǈx��S�j��o�ILu2"J�%��]nJ�rIB�:5e���#*���T��",>�X�e����!�����	%��I"�z02�%�ȝ>�AU���(���5�Ved�pBQW�%jl�u���W�w���`(�arrW��� Ki�Wc�҂�cVY,�p�����݄��4x%��̉�i���X�R�ITcr7h�aJ���AW
+$��X��v�D'ֻ�S��쥑�
)-�$#��=Y�X���27i�6��:\B"	-v1�&}��$M��PVV�gűB�q��*���UT��B|q�q/xonH続���5�{��>��fd:-3�vN��ҹ3��$�#��5ns�x����]i�V_�B�eъ3[<	��7H`�3"��Fw����=G��=,��%����M���2�B��>�u�ƏFYR����9��,,׻<d�(���d%s%%����\��vѝ�j*RS.�fN��9:jT�f�M%zj�m��_:�$��c���:ӆ�0���UV��I�����u���ѹ��ઢ���S�3@�:`a�M˽h���������Q��φ�تxɀ�n���]}���_��}6e�}��¤���Tnh����>%=Gݮ��+�э��]d�k~m�8ź�1n=u�u�x�I��2�t��Й�NI��deSWe}60��!�7&�/��?|����O�Wlӕ�t�����<.���enYD�l��z�?�^U!s;��B�8���2�#��⇒��4h��'����a�8vM<[g�!��vLDQ?L�7�60��G�I�8����[k[�-�\|�V��l��pM�<��d�%�oUUhO;Pٚ3����2|�4�9�7s�\��l�qxŨ�Z��ưz��h����Wț�}�쒺6�������n~��d�;��`���Mv�.��	��^��vM�ӟ7<n
;j��C��Sd��_����C��8~>[���V��q㮣�8�2�i��cn����ׄo'�!��T�?��"�Y@�Uc��m��Mg�~h�9���=���/9�t�כ���fv;=�����l�7���Gάa��-�ߟ^s�߃��1��&\Ⱥ���n�r��Ow�>t�3�O5�䜇#	i���V�G0x�de'+�g8f�Y�Y�h�Y��N����*B��o�cB!!m�����������}�c.��F�GS�,8k�揻���.}��a�S!�&	�Q�H���/���9̓����f\�~_��l�8d��l��o�b��:x��㯜c�1n��[�ui�תֵ=6��}�Q3�������U���s�������e��1ͷf/ʪ�	�<%�CB�tf�m>������۵����}N��)նWϕ� �^�&�CIf	^L�썶~B�k-r�dc���������}��Р��؟��h�~��::�5�;59U�|���1��V�-ǎ���٣�L�ɥUV�h�����kQ�_�P4d�D�W��v�*�����h��>�痻�bg�����T&�3	�bXQì��]�!�$�Q��驩�ƌ7|�}�Φ���G�l��R,~����jl�8\?l���f-�-ձ�q㮣�8ۼ�F�]�P$!m�^*��&ɳ�Y�P׾h�`q��c��������2r�Yn>�?�hҲ�i��S��fɟ��)3ŕ3�8s��=F�!cq��[����G+m�{	���:�	�v�P�;��C����.}���W��[|돖��Ÿ��Q�73��ݵ\|c����\�5U}�ϋ��cQ�J��N�Gv�ꪫBbg�l�񿹲��������ϯ��܊�ncƩt����;3�ؽ��ޞ��Iǭg<��5j��>��'��fm��'q�N��i�똜����l��ɜ�&Z���%T=��H��f���,:w�*��l�!�� ��ή�V�Z���t��W>��`���`�؄>�4��'MU&���n�?|}<0�
����fb�4^.���ʤ[��-�(�)��}k[��>�[U꽨�qx�žu��uo��e�8C�l��C��ȹ�1����&��_'�xVG�$�E��V t��p�\*0�6Y������~�)���J?>�P�?'����̇nY�|���}��̫��Wwb*�ݫ.{G��Yg!qy�d�̅LN�둿]��ƍ:{rl����xO	�<'�DO�N!�b"'DN���Љb"tDD�8%��6p١4A���'M"A6 ���y��X�blM�Bx��6l�2|��	�"%	�b�\[׎?-��0���c�1�[�q���Z���cc�0D�� � �"%&�BY�:^�˱��.�뚽��������ښi�_s;�f��㢥��1m�L]8��4��ޯ�H�z ��ә�/.qANo;�]x���s�*����5"��^�ߤyT���/ϻQ�V_8�Ҫ����ffffgҪ����fh�����e*����fa����V�V�����gN,�0O	�6YÄ8;�G+8Ҫ�Gu�H+� �45\7�I"�G�=�eq��i*/�YM��Rν>�y+�����Z5�w� 1���͟W�������2P��~�Pt�Ӭ٩=�'?c�W���}n0�}�u��;^W�z��q�-n����]GZ�}~��߸�AXм����
��m��[������r���:h.��_\�ں�.�ӲUO߾j�����=wA�5������N�ݐ��H��)�gS�~��7OC)�W�T�l�IS�)>�gڦߗ�ҽe[�1��[Z�<|t�g��M�Ƕ��0����O�z���j���5��s3:����s���L��gM�ۍǪ]իfLo���nmٱA�T� ��,*u��iV���M����0]��ٳu�=���3E�ғ�<��ܖC,=ߖ�r
��a�}=�x;(���{e�L��������p��`���0�juP�~�}�~��}QSh�,DG:67��� �����3w7���]6�Žc�:����6YÄ8;�E��zc�s���p�3F�х�[��|f*/�4p=��.nM����Cb�a����p��ʹ]7˕tl=�����5��:L�^#��n�PY�&~~�8����J2-�ؘ����5���~��~����>u�|�����1n<8p�rhkxF��UU���we�W{J9ڞ��MvX}�>�s���͢���6}V�=w��o���������(��<}�0��p�C����6l>�Tx�#��ܚ��.�KZ�{�t:4����ja����G�[���[�[�N����6�;t�$���i���&N,�'��磎��Xٞym�>b疦��3����`|-�;��+�s8֬�7�g�{V�*NM��*9ٿs�t@�l�N���վ�E׺��_����]��*J��w��㹸7�Q흢��5�=B�U�{�(�@�\w��Ɵ���+�r�5�=�^�����T|c�k`��vl԰s�]S�FY���V����C��T�5�7�����`���O�:�o���qkuku�#���p5)���FWZ����g�����'��4Q^nfk���՟18.�ΌՏUUZ0�M���;y��el.vk���|٘�o)/NI}�7;�=��oo	Ǉ��uX�\�f.��l�y�1�)�_ћď�b��<���kG!�@����ϿB�aӵ�m#פ�	�IQ��I4�M����%��VB{��5�����Q�њ8І����E�s�^7�X�,��\�P�|o�?L>0���8��V�X�:�:�$�ۓ�kLs�UV��D���6v�8�m����A��������E���5
�)��v����M��2��H���;F��ϞK<��8r���B� r��uC�x;8	F�*"��NOͳT�R׉����q��YӇ��p��юbA��UUh�Rp���4 �&{�2�4g�?IEѐ��[�V��n]�cw��ZU���=�Ϧ�V�'��p��w�p��}��u^����*��٨�R4��Nm%/�[Z�1kqkt�����:Wg��t��5Xڗ1�*��r��,=��6	g��s�����[o����un��*?3#��>�L��x���8��nl�a�dɳ�+�]p��Y8rI�nV�����"��=�J�V�'�e��O|w�?V�ڧ^״�0u��1��N-�έ��V��[�ukZ�qn?(DJ ��<'JM	B&�D��tDD�blD�4P�$�<'
D�"lDN	�<'����؛4"l�4%	C�}�!�A7D�E���kmkz�?=[�4�֎��a�'��B�DM���V�1�6��4��0�,��D�4hDؚ,MM����(پ�g3>��{9��6� �R����-F�jʹ h����e�k�e.\�����˖�w��B��
�ҙ�Hsro��֟��~�g�S��yy���?ë���qNjL�jֿns�~��
x�],̧��|7��}��pQ󊫨S��rˎ��O�ʳ-�q^c=�q�җ����M��x��O���g �Y�{{�Όu���b:]��-�&1�w�c�ɗ"�Q7����zيG+�9�o���EEj�4��I�y-R)Zl�Wci��کV���Q�n�u}���O�Q�G���/��4��wwo�fffffuiUn��������|�U���s33331�V���s��8pیc�[�[�quq�o�̿�H��V��	"�[	,#�PR(����ڪ(P��v��v�|�$�R�e���B�,U�W`�=�WZ!1FɮfA
��m7��7 ��*�H�U��P�k�P�%V%A�T�����ptUY�[.M�w�2J[*�M��0LE*j�SiEb"eee$����D)�V�,����d�¤������<Ȋ�c-a ۖ�b'ֲ&}B�GX�Q@�[~�Im���R|2���b�L�:(�b����"�~�q1�_��
R���mG)%j��@�5H�(*Z9�̍W�8�ֈ��~��5�i�ˣW�����[�?6�m�������5�VO��r�[��L�5��힫Q�8s�2��ag0Γ����]|;ռ�s�ݻ�s,�nڟDva���{��R��q{9�;��֩G��¡Ð�2x���;K�A��=1���Q�O����}Z�/��.H�~�:��&p�y^�u�S�N9LȈ��m���.=ԊDӎI$�X� ��?(��?����i��%W���Zc۫qkuku��:tN�,��Wj��"gn�V9Xq*��?oÓ��p�ΨJv%�ι�������0��N:.���mh3~~c����j���=;8|mUp��4�sF��N�Њj	�nb�G�SG�-�Z�Z�Z�c���{�{�H�� �c���!��k~AQ���>�Ϊd�afC
k��TE��p�r�(��,<Q�R�s�9{�L�&A���U��ݻ�oU�Hj�tp4Z).�	}@�3.b�t+�58rd����v	r�4p��qkuku�#���<n���/�$Uc�T�z�Ð�����4{�(�9�Gkm2�Z�To�!Ӂ�?wo�Θ\,24C�}�t8��d+]xɺ�W(�Ē<%V8�M�7�K��a�`�*!����7,�����c�1n�n��u�uǍ�~Cy��1�w/�߳�X	�ڕ֊��ʭ��sL�1�e�e? ˍuh���ǋww��̈́��M���u_��'�0���g5�e*�o�s�N��3����ҡ��n�p�3�\�|o��獙�g4���&�g;�+"�3B}U*��Rύ�Sv�O
��2!���V��^�0N�W)Z�_��/A��T�-V��F����ɺ8l��f�=�mm`[r�ķ����*�5
�������J0���[�[�quq�n���g|U�h\9]��������n���c�ʲ{���ڜ�zns��q�����t�7e�N_*�h������揌4��U��B��QUuc�cB��ǯ�f�X5j���V楗=,���#WJ�+�;�L^sh���]��U`�t�ÂsI<{��������r���z�c��c�-n�n�quq�i'��I$�j���G5�����Q��VCF�����79%oY�CA����9���5sY}�����7����b��ɪ>K���ce6x<l�3����J�n��cĔ�*=��Z�7OZ��Ca�I���"DxE�q�1kqkuku���:p�f϶~t�O�P�j����ð`ѣ�5O��}h._�uW��,�n�**����+S��>�͋(��,J����T�ۣ�R��4�'*��
r���f�ݑ��m�TC�'�I��]iʬ`����[zr�ӒH��z}Vٶin/�t���lu���m�\|�V�XpN��657���ne4e�c�d�-��HW����a%R�Y�r8�jm� �h.�m��f�m��NG��u����_B�ן��V��Ů�
��z���Ԅ���W�͖:�>km�M7��.�y�*婝��$v|�f���n���*B�gn'���81�!��G�*Yن��U�[R�����8�[)��(��Ҧ��=MӔ�O)�eD}]䧕�X,�]�ddn"�K��3O$$���~�c�ۯ8��-��V�[`t�8Y���<�7U�--�Ua�����>�!���D��T�UTtp���fC�§�r̳�?&�!�Fh�5�X��5�x2�Ͼ�=ތ��inj��G!��*�.�+L[������o��|��״�u���=w�z���n�պ�V��[�"'������6"""x� ��b"p��"tKblM�d�DD�"%����"5"#r">�<'�	�E��6&�١4%NQ� ��I�����lК!�:�1�c�ź��Yk[K"X���'��ba�
000000D�&�ѦDؚ�)�}�ߝo��ӯ���wzi���;��_{�;w�ޟ��L�?j��ٟ��ng2�C��;1��g;zu����k������}_�o];ؗ|�Oh���n���|�U���\������V���s33333�U[���̙�������wwk�g~~mkqkuku�uq�o;*@u�U�����]��U��a�v>�&�%Ϡ��E�I���Q�h�l>��>9X2hٲ�'����#�n�����V����چ��_K����*>.z�CL��ߧ�I$t`��߮.Mꁣf͞,���u��uku�uq�o{�V	�w9��0�r������Ϳ��;$S0�:Q���9��p�kZ��0��������t��l�@�g��>xu
���{���w�h�y��G��-��^�w�7Y��\~�1II_��������S�[�-��Ϙ��q��Z�m�]G\x�7oc�9���̟U���밥࿶�P�P�ܲ�,�1���7��a�uʛ��~ ���w����w|.�rk�d�[ݿ;�M���]{}�β�^[�w�f}���Χ�ʸ��;�^��������绱�Ŏ������z�+�j�FK��̃����tn���RQa��_}��.w�������k��+ݜ>�7,�r�e�>��t�j�%4'�<;�"ԕA���vpN����nt5K$�$���+����۫q��Y�σ�D����?]�we;��*�if@�:��8a�S��Ml��+��r76�j��B�ݼ��.���V���~��:zCBn����v���*����4��y�m������7$��&x�m��mm���V�[a�Q�.{����2`�@�~@����v��0�,�/K�2���`r�L��!�<T�!��;RύO��Ϩ��_י���^e�~�B���p0��{�~=#��v��Y�U�`��U�H���&���UM���MB�f�SK�$I1㏞�[���\Z�Z�Z�%��.�(���x�W;�d��[��?e��3�s���:}�!��c�q��|�n���U&.n,��q,�^S����g_	b�K��q1A�����=0C�.�N��gj~��EW0�k��8pf��S�;5����5f�d՟�����;�ԩ�.��O���m-�����[�r��]\B��~�S�������|�������P��&�p���7���/�Mmf�jx�Lb`�l�"[!cM�&�@CS�� }�b������Յ��������S��n�1��9�XX��ʵ�k��ZVݞo����}}�s�;���u`�����}�=Z�<�Z�1��b�7�F��w����hJ��Ht��cfd*vx����g|�#�gvD��BNl�1F(Dֻ�QZ��v\0����������~4h�.��9��k�����\�ǐÓp��?|�=
�J����Žu�6�-n�Ű��o�t�7w�U'&�&�?|4t���P����z�����f'�w�_?��G)�	����e�p�:֎�M���¥����L���V���60�4a�EA0a�ˆ�g5�5K�Vr;8h�f�>mn�ź�î#��wٮy䧗k{UY��e*#*����:np���U^�|^�*.	���?J0����0���Ջm\���Z5V�O�	k�>���z�.{��m���r0��!� ՙ�gb�����M�����~[���n�Ű��e�3���̕[��Ϊ��?M�>��;�J��>�����s�y�Z�Zӟ�$������^<f�~�[����	�՚+�c_Q��Th��A�1�G���Y7��ܑ훹4RRfiy�>�)�ϗ��EFn�ՌdR�̘G3P=�w��I$�$�I$�"�Eǩ��{��?Xz�~ձbl�� ���""�"�A
L'�K�)��,��0 P �;��. �#`��I ĝ�P�ă�E"##`��`�bF�#�b �bF"� �#��DbQ$�A�DFtIq1 �"DA�A����$`�b"0A"b"���bbF ���#Db�D�"A��1F�0D�0B1��DF"�"#�"0DF0���`�#Db �`�#A��DB0A���D@DF!�#Db"1 �����D� �`��"1F"#�`��1 �F""DA"#�DDF0D`��b"1�����t�X�`�#DD`�$"�F��Ȉ�	� �""2"#""A�""2"#""0FDbAb"2"#""0DDH0DFDDdDF"�D�`���"� �""#""2"#H�@DFDDDdDFDA$F�0DFDDdDDaHH��1"#�#`�dDFDD�b2"#`���B0D� ��F�0D�0F�0H"0DF �(�� �F"#b0A���D"#F $DF!"#A��.��K�"1F"D`��F��A�#b"(��A�"D`�b"0DA��"1F" � ��Db�DA�F�1F"#�������`�����) �"#�1"$�#Db"0DF$F"#��DF"#��1�Db�DF�" "#�F#�1$�A�1##`�`��H"���!B�D � F F`DA*�B����	J���!D�A*�! ��(���@?�AZ�H"��R��RB 2 ��FF녔Pв,A d�	  0���	J �UPB�J*R�JQ�TJ�PAUR��D�)*�J�AAH%U ���PAP@��
�%*�	UH"� A
A*�ET	B	UPJ�B�ET�D � J@�UEJRB�� ��!HD��A�%<���	H%AT�F�R�"	H"	P"RR	P�U�D*T"B��`� �]� �D#�1�1BD �"�"�T!)BT"	U���`�DdAdAdA`�A �2 �"��JB�P�%!�P�J�D"B���%!JB!��B��J�C����JB!)
�D0A� �A�ai)Ȃ �2 �1`�BRJB��!)BB����"� �AdA��"�"�"�"�"�A�2 �2 Ȃ ȄDDDA �T!)BR��!	H ���0A�A�A�A�� �"�2 �"�"�DA��"AbA�t�D�BR	HD%B�P�BR	P�JA)�RT" �J�B�B��BT"�J�B)BR���"B"A�B!*	P���J�!)�!	HD*R�R��!!%!�� �A��AȂ �#�B��� ��
�J�HD%B!*BT"�JB���B)BR�R��" � �1@b���D%B!*BR�"	P�J� ��D� �D� 1� ����D�Q	P�% F (QX���B
��FF��#"����HD*R	HT�*���JA)
JA)
��RR	H%!R��P% ��R)�<B��D�{Z����R�� 1�! 1�F! �!��1A�� �1�!�"�`��"!U
�FB�� �%�5HB��JB�!��*	HT�% J�T�D�0B1A��F1 �b�0H� �� Č�A�"0A�A� �#�R!ъ@���8�[X�:4�	�Hl������T$�@R0P�!a��'¾Y��3�~��_$ٿ���!���#g7�NE�?����2����!xn�nBL��r�И9J��ok�hڵ���ټ�����'����M����F�z�t���*�?��������A���Q�4^����?�4@����h��Ѿ��?�="�iF@��%
n����Q���Ʀ���!����� ����*��t*~�4~>HI�!��i���p����Bbu&K��蔔����xM]8�n&]x�������˂^B�"���;1�F��6�@ XA�AS�D�u
QIQ$E�b�TE@# Kd]��
hi�kY�*�۳�w\�+ ۢa�x���hT@U@�P$AT02��@�d@A��{�/(t�`�&"f��w�x�r���i����.
(?�a��x����-1y���4T���Բ�|����=>���D�u�j��.����\}����9���K��H�y�!��ᾷ����d��s�QT���ؿ����W���������p�7'A֨���t>�b��/[�Qk�p�M�r����ML�d�R�D��PD�Da�م�k�u��A@A�'�'0�p�y��e%������`渶�F6��\��/K�^	��l�9"��Ҹ��1��ǳ�r���s�QT���Oq�����C��a��>?s�A�X��>9�-�5�9Z�P������ˠ�z�
u�s����C�x�%ܢ���u�����A��WȨ��<�I�G����x�M�����C6x��׎h�"l�b���I� �0UpO��43h�6����/_�Q;w h��oـ�<ئ;V�x���MzC#EP�=G����w�^��Nt�v�~���$C�=������g�E:�HVX�
�R�᱑����d)�jq�DO݊z-��Ȃ�p?��8���	�8%Ҵ������,�e'.�=!�^��yҨB���nL�����ܑN$����