BZh91AY&SY�fq��ߔpy����߰����  a9�Ϣ�@  
�    M  �ݪu��  X����@%
@*(�P@(
��(�@�P�f�T(�H�����@"l �P@    � �
z΂���l��o���(���;���v�͋�����{u�:W�޸���x7={�C��b�o��x6�l{�z	z^����.��hb�����+O{�*�.�}�f4��w�_Z (� �7�� =*��z�Z�e���yW�{hQ��@�KC�v��W�
�}����zz(g��{���
 W���{�Z�4R��ϣ�%|�݇Yh�ۦ��:��������(}�o}�>�E� y���  �}�Tև����E��^��P=[9�1�nG�t�(��o�[۶9(�w�qq�sS��l
�础��kT�)�( �p�S����)�w4^C�A�&�L�� �ҝi�P��civi�{�w�����n�s�O�z}�9^����P�� ����  <�@�5��rtq�<���ƶ�^�G�z�k�� <҂�{�0�CCJt��:�ȣ��((                    P   ���47����4�@1  h a����"4� �i��M0 & 0i�R�e*4h�  @  ��@��DɀƓC# A� �B�hL�1OM4�4b��i<SG����!e)R��'��h �A�2ܟ��/ݴ���Y`M�4ڛ\�.��h���~���n��^�`��ʠ(��`��#�?��1��{��j	$ ~�y$���o�?{������>��2x-�S�	h��!v�* Bh��T5�5�eU�~݀*��Ո����T�i�x��X
"�R�H��%�@����~������_~�=g�������=��XW5�4�âzΥsV�M�Xv�����iĴ�{'�����Bʡ#D�P�	�FzMt��,��6$l�:x�����l�u�I�&�ٲ��r2j�0���FZ��K8هVSxt�0��(u	�}6u�g�zWB�"q���0H��jn�zy��DGmW���-�a²%�L.���})0D�5,K�VA�H%>����e&�V�y��fۈ���YB#؉ŕ�g�D��r��D�n�`�D{�ZGH��w)�D}����*��r�:ܤE�]6U�H�R'<��񕨛d�F(��%�DG�(}��� �D���:�".�aö<��:y+�oە�-�KYI����i�H�})���L8;��:YUg
-�D�^���z��5)m�D먈���}��O�"oە�-���r��핪׮R&�JD�2�l�S拏�ӑ<S6o]I�2J���ʮ��2�t�UK��'r'��u<vN7r��sPw8#���Z�8q�9&ƥ���o�=�Sų����5��!�AU}4�j�z�U��j$��᳏�"�1��w69���M��o��&���u���d��N�{(CnW�;*�|H�URxrI㬃�d��5"5:rDr&�U]j��� �JS��I�3�a���;���g�2ӻr˾��\_OC�����h�9��%�9��L�f{�+*��PL�
�'ԓ�I���z���֥wI*�.�.�.��NħjO�'��BJ�K�K�'�Wa�į�+|R�t�<�Q�9�����D�KF��s���b���m2�$W����o���+�}�o|��m���D<(��Ɗ�{t�	�M�H=�_$�2�萇��5�<��'a���M��R&�'SɈ�9�k<IZ���'p����}�8�؞l�Gh��Y0H��Y�*�l�7$N�O&bOJzMټ�	�u�=(�h�kd&�ӛI����:�Ӑ��גy2�bX��;�\!����D�;��C��;�g7�7�Y��	znN���10s$��䓆�x���$ć�'���݉ݲwg:��&�Gü�!����2j!�Hz�;�&ĩ�5Ӓ���Bд:��������&�%����⇰����5�DJ�A"&$=�Ći:��be�RBi:�O2D�,�✑�pJ��	:Ɍ&k�O_�L&�X��`����u�%���='����zC��Ζ�N�-"x}�P�Ęt�ɮ��P��U$D��DO=%Ӳi)֑6=���LH�9�&����}"_D�K<�$�%�[H��҄p�F�DN�DE:P�q/ۑ�����4��cp���Ĉ��L:S	�	�D�I��DLĞ:G	����͓H�'�m"%u"%):l�m.Y-=�
mD��'��%�C�8"{�&^�H�ĚL�8l���tH��K ��"%M��H�ԝ!�m�4q�"�'zK/�:�L3���u�l��R%��M���&�t�	��K�cRQBQ5�<I��N�DF)��ȝ9�0�	�!�u ���P�b:�TN�N�u:WgJ��ODh�0��N��D��ì����n#��O焼�L9��8rN �HW$;��%�C��&23\7����y9e��d�u�tG�:fO�x�U,�n�5¥���Vq:�<��G�H>����
�W|#䮎�%�fj� �����#�IExN�fQ�	���#�r�g���k��Û�|'�ڇ�q�I������9�u��}�=֧���idܔvNt�����Q7��"P'��F�::ʴ�0a(X�����,�t��#�K�"���@A���TC��������PFUDF�Q=�jA9=SH�"=�O�"tv���H�����"r�#���\��n�Q����"t�AUv�%�J��d7�A2r��o*'J�SI��L66H���I0�[��4���D_TL-jP��S\ ��tۺ�#9Q�TD��(�X�i��'G=R�fTD�8aC���T��po�v�%�g52K/sIc��D_TL-jP�w�N�y4�6��TDw�/m@��Dw����#2�'m��f��d�&͜7"<�2i��"�݉�v��;�Nd�c�N�^�.�m=Sg(�{4��E�m���M'�(�%Bf��6Q�C�H�e���y�<7<p_TOo�8t{ҨM���.��{H�50��t�x�m��3�]��Bz�n^�E�D�G&l��E���q�8,�Xư9�PC5&ǻ�����*&{�:���g�������N��bRa�jt��t��JN9S�qʜ/^6rJ$��SOf�MmQ�eu�B�����8��gj���L����2C"�l�����"48wR7ԏY�j�2��$:�^"��6a8lu���r;��G�R�����{����r�T	������G�Q��Z��jv�������[����㷨���H�i,Jૅp[���3l&%�BCc��!��S7G�Vu�����v�.����5�wo��贆���Dƌ%�N�����yҹ�N�*rJ7Q�'���\������Q�iQ�e�|�aH��w�+���h��m�9q�޻G��s���B�#s�3g��6�F��w��R�]"��@MQ�SG��Z=g���:-r81��5�f�;
ȉ�H"��ؙ�Y���p��Ox�r5�R�F���#�E{}�U�e��H���:�N,��<�'{��r%u�#���{#�(�w)�D}����*��r�:ܤE�]6U�H�R'<��2DK�̕�Å����R#�=��i�H�nR']DEܬ8;�:})��+b[�H����핪�r�(��H��W����~��K+�ͺ��w)���ܬ6;�ӯT�M�)��"�V}��O�"oە�-�KYI���תoO%%�{)���L8wc�"v�[&��I8S$N<�N��蕓:ʢ�U^rVd�'��u<vN7r��#؝eRt�Lƫ/ݕӒXԳdGr�؎N�1<q�7�	�p�J���C&��橪�k5�N�R,�et��G2S��dzONQ9 �G��ڎD޼rNN2t{{+;T�'�*�0rHvx� �vA�Ò"WNH�D�x�S<Q����q(y���L3qa�A�w#3͝Xg�%e�v����q�;�mal�9���З�,N�7�:��{/z��Q �P.��RO�'�Wq�䮵$��I8����J��Jv��R}㡇�%i%�&���Ev�+�q��!�B���a����
:g�m�l���z�tN�L{�M����^��pV�@�{�eaa ?8��T�Q�ݑg������lRR���*Ð\L9~�B�&!&G����Y���C��?�����ݚ�����>�h�}�����!���*�Y��v�A���4�>!��բ�p�K(�C�1��P婴ae�H�2IՏ3��[���B�{L�aM{�l�U2�w��a��*�`m#���4\�K�h�$m��8a��\<p�vX�+��8鳵�v|�4r�'utM���(�$֥{�4h ͋���1k��}$�msW�Vݟ(bCe�*��)�ׅ�t���V6���*���5t��=�z@�9S�Ѻ4�F�(C��h��o�-�z�Z�W\�g�g7�e��T���J�Q��[����&�k�!�C�������R�@��DCDV|�Oة�n�4p�Ξ�$�L�.�����L�(�����oٷu��d�yV#]��2�Ff�E,��q��Nd�L(�
����p;\�M��ո��z\�j%G*a�=4p��~Vޚ)��D�ɵw������Ǌ����$��E,�U��zc�'M�Y���
#��Q�O_6rsL��=PF/r���6b@��.:eѺ�G(�2�Lh|�����l���"�W��GI>��3w���Ζ��@K��W�D�PK.����۷��!u]��Z���'��g�-R�x�������˟:v��m�)  ?¼�Ud]W�M�Ff>���N�Y�faGw���4�4|��:t�,,5���91���R���ߏ����f�Պ�V�C�XVI�UQ7����l�m�3m�)�/�H
��OUa��������l��7�r��җ#�ꝺ3ǝ��tm�Ç�Xf�HٷNΚ4d
z�ꖊQ��2���rN	>�Mk��ٌl�M&�=���%+��M��	/�Z���Gn��l�6t٢�Gw�$� �ӧ����=rt�Ji��g��v{��1h�:hC����b_rr�:6��������P8�t�G���<�㧷��4C�����B�ַn�-��4p� :CZߥ�3Gh���K�L\:gO�o=>h�E!u�#ݪ�����T�������M�5Y�T�EM�*���e;H+:E}u){ m[AqVt�q;���M^OHpr�@n9�޴@̹��tʷ��`ѥס�� ]�����>���y�'�b��in�d ��Yύ�,Ѣ3//
��\��@�م��G�
�Š m���N��T����<Qj��{����f�@D:3ᥘ1'�JtJ���LT���b��c3�[� v�c:C�܂��}7���Wu֗G�ٍny��+_���Z4P��	�����%α̘�*�4��gՔ�ڻ��G`P�)�J�Ʃ��Hͽ�~c-]��,ͅ�:TI�0xä�}|Ee�+,|Y���W�DT��!гĖ��Dg�'-�f������7Ȕ��n4|7;]J�߾p�ݬP�����g0&NBB!�\Mi�'Ⳑj�끈��Fʶh�"6���T��l��ҹ�ڏ)�3�N�� ڏk+�J:a��U����x�l��w@,M�џ��~'�&ƍz��������G���$3�`p�DQ���>h�������T�J7��OO��тt�ԍ :[*��&�r�{qU�ς*r�=�ՖO��,Ѹ����g0��(Q�ɫc!��`��Vvk�4��8��f�yJ�l�Nݸإ�:�7�v��h����n�����|}d�ZV?SD�:,��<ET�+�(႖��s�+M�a�D�ه�V04Ѹ���Kת���]p�oS��G+���
�c�F�Qf8i��ި\�1"����Z^�x�:{��b�Ub؋,ô��e��a�o�-��
-kWM�`�}<�xh��>�C|����3�wf������8YG���0��[[N8�)�e0�,��w{���,GNFN3Nh����mHd9V�Ֆx������|M_		�*i��&��{v�J��C���h����>YN�8p�F�~�^6hj�R0��#Q�3��Q�<¨Q�n��h���l�HO���S�~6Pj� j��7R�S:oq��u�
����l���L����gf�;M����;.f�Q���P��W�������ɧ˾���<K�IS���k�A$ތWm������X�Ǖ��0�
�k�vh���>��#�y�<z�����9m�zY��>�W9��~��,Y��O/�Ƌ�oM?�����ٌC�QGo/9r�������
�n�zx��Y���gO�;�Qf�˶I��%�D��\6a��Id��-෰'�5y�=�N�C��.�ڵB��p�u�"ʹ6��6x��>8��}:i}�]��d�гB������sw�͝��8le4A���%<t��TI�z]��H3� ��w	`CG
�6S�p���gw&���}A`te60<s{��lѢ�l�e(ѣ�H��,�w�el��G��8C�p�}�kd8��Sc�ｯ����?rh����|�Z65#eh�7gS���L�Cn���2���K*F�8p�f��yL�π#�<o3��Ц^7�e�o���U��7d<h��&�C�|��'�^��x�!��x�M;�=| p-��;u�i���o�m�:Xx��8vh��o�62��x�F�,���S�(�@(��ZO�TAN�٣rN ��Ma(��京���ʏ?�0�~��G6�'�,����A ���Q��Fѽ���n�ּ	%Z��	���Y�ļnS��6Q��c�o�tnS��(d�ep٣�D�V�v]i�2��U#xF���N�����Q^�D�,�$���;apŹ�wZ5�Z͝����l�K2���ŧm��8I��w�C��x�1;�#�a<�PP���D�Z���ei(}B���8�3k��{B�8I��2��UX�s�O�=v�&(��Ng��/�,�7ok��Y³+f�%[Ӧ�:�
Wyxh�Q|��4hŎ�7�b�a5��l��dz���.��S=v	���WU:p��O[^��z��}����1�ꦤ8QS*� �wzm���7(�Bz������x �a��$�wn���Re�wv�ٳ����%��M�}yl�ԍ]�f;��i�Q���1�b�[=��|���$u�8�G��[v��
Y��_<���wΘ�A9m�~��5z9T#l���W&��;�+N<@�7�|�L�S�L��q�
���*׸�J6I|TeY�@C��OC<f?I���k^���(�9�~�wP�^��-���pѠ��[�/��~�]4-��ɢl{���t���7����  ��8h�N;�aG��,�F�vM�>���x�N���'�D��iGf�<x���ۗo�aS�ᅲ��
)���]����B�9y}��9������f����އ��㦍nn��Fx��N��),6t��,�[�N�1��h�ϭG��$���V�}��j�t̪�|�O�6۱�뚭}{t�A���U\r��u��$���0񆲳^V�0r��
i�u��Lj���P�����(P��1�������O����<�����{�������������l��p��}���\q��nZ�p�R8�J	��U\q@��ih֓	A�&V���)�� ����f�R-F�J���]�$�Ji��;��9���-��ڂA��b�Y����)��B����u\�A�R�d��FϷ�c}f�:��oB�i�A�IbrCX�iUD�4�wR�kvJ9v��F�q���A\���)��<{��F�+d�}��_C��)��4�n3s.j=Fd��iX�BmB
�T	�B-�F��5q��˪6`���d���oI܄,1��M�b���4\E�3���LbE��Mz��U5-�/5�F���(��Bf�u��-���h�ԢH���
۶w7YB7�m��2 �����on�{hӵ�<� `+U�6KTL���"$xă7\WQ*-�IJ&��CZ1 ���!-��Wǥ�}d�h�l� ݉~&���O�6`��ާ��6���!��*P-y�.K1�7?��p*0��c)�q���Py�XQiZ-���1(8Q׵��#C"_�|==4�ThC���s �f��4��ij�լ��ND6�F��	�g&�^�R{h�y=���[se��-�c���+��o�{��J�&�a�^XHOz-�8�VP�8)�cGi��c�b�M���l�5Ċ�&�+c7^��!j���m1�v&�;l�+[c%�r���[����fV6�B��Z]�̱&HЉ!/t��i�F�s�83eȎ�d@ܒ��H���
��'w��Z5
Y��g>H=ڌ�Is5�b�q�IH��+K����H!S�L�� �{�ztâA��8������R�dR'C-���vA�!}���d�B�F@0�DDS�6u�,��\��e:�#��$�b|��A����x�]��)ćP�"Xy��\}f��q��S�����Pw��!�'=����y�P%u=�d9&@e�gp�OR�I�<�]�J�q-!�{�7܆�):��)O�w�5#Ľ�{�﷜��_փ��~-��s� �����������*��y�ʲ�?p�<�����~���_���~���rC0�%/���?G���}��v��Uڪ�Wj��V�^*�Uz�J�WUUQUUQUU�*���UW���Uz��[Ux���/V*��*��*���Uz��[Ux�UWUW�J���X���^�����^=Wj��[UmU�j�h�굢BkPԚ�Ԅ	�!�P) �
PHu���$2�R*PA(D���(�"P9*㓈j	�5�k�[U^*ڪ�V�U�UW��Ux�j�U^��Uz�+|��UŊ���UWUUQUU�*��v��U�]��U�U|���W*��U^*ڮ�W�UV*��v�;�u]���iUUQUU�*��ZUW��Y��@$��Z���B�d���$��A�F���V�ZfQ�*�!�*�|ͪ��U\b���UUTUUq���[U^*ګj�[Ux��U�1v��V�U��U\EUW���Uz��W����U괪��U^>Z�W����U�*���]�{UUUUUb��"������V��kR�!!� %�0�J(�F�CD!�m/������ٹ�����*���U^�Uqb��"���UU�Ҫ���U�UW��Ux�j��[b�^,UU�UUTUUq���ZUW��U�W�Ҫ�EUW��U-ZUWȫ��j�J��Wj��]��U�U|�UW.�db9d�H �!u:���d9 �(jhT�3R�hA� �@�@\%EԀd�d�ى��
���T�z��
���2�8��054�JO��>����3R����?��o� }>�~c����8?1�:~�����<$�"bNA(DN�0DÂx�,��!b �	�6Cb&�؉��tO	��&	�xL0��8YB`��Έ��'�"A(A6"tN��`��D��ĳ�l�"'DL�"p� ��:"`�"a�0��0���e�&�d2iCH��%��"Y��:x���8AD�8"xD��	� � � �	��GRD����16oM���u#o����^�КZ꼥���+5#�6q����D��F)�����ġ���t����qu���a�f�B�d�E&v1e���x��vK�4��i]��;b��4J
(e�k�sI�k]��82U�6[,�k�/fٖ���b�eԛ���c�^"7dn��asZK�XFm����Ժ��º��u�������x�h�}���&�Eѕ�dm���LRB[���JXJjX�j����s�26�9��d���p�Sj�u�*���V�2�WBSGLݎy)�ա��!����j�/u���;�Mҕ�VZ!4+iT�{�H�Hh�I���Ek(�	,��A��7n��`�"C�]�u%�s��J�]
�5�Pl���j��WjndZ����Z@�nkķP5F����L�J�L��������J�K�"�ٵ�n�q�im�5��t�����)3��-�L�ieim�l���J�+0F�e��0l��4@f2 ���%G3��F�H�Yet"X��1�ͩ�P��V���X�-@�f�Y�鴔)�vl�km�ev�ZM-��j����� �[0�h�d��b4x!�������uu�V��8\�LS��ĚMa���\	iq�k���Bl�e���e�	uX]r�l6�HhԈ��)�ҩ[Y�YucpL9�-Тk`���l��b�[Ͳx�g�ײ]7�ն�ձ��^T��4�#`cl��	n�vcF�Mu�5�\&��q��]]D�.�-��İR�-u�,�ް�'׼�g�`�K6B'7S�ĸJ�]tP˶ŕ�����q�V���r�n$l�B�@�N��#�}�WmV2�(�՚�T0mm�k2����ص	��,#�.�� q��]K��@-�5 �4�٫��[,fml�6���]��6��Ț�mԺ��p�Ck#ue�S�+[Ym�W>Ry��6��.��Eq&.�%���P��@lŖ�^�ff39 �`�i�ͷS��-�i�\(��5-v>]�z���흺2��-�(�%%�ٛ1l����u)&MV�Q@QU]�*�U���ܣ���	B%QnZ�r�]��UV��VPǔwn�ZQ��H��hvyUĒ�h�{�	�J�RAV�j&Ƕ�9w�/hkt�m�͆&L�:�@`�K�e6���]O�{oVek3,�6�Q̮u�lAsa���sR8)�XݪhSF�kk��u10\6����l%,˵���Ơ�b����Z])�p�[,K�6�[�F��b�v΁��ǘ�lʼg�]f��~��}�)�A�f7L�]̠�r�ٓ4�����8��<���k(�&��`���ta���1�3[7X�r�L��B��8m��iJ��*�:ia�����A�M��k*�6�i�a��0�A��m�]4�WD���d.6p��e���c^l��f����2��s-]tWG�TMVZ��g2���-��ٲ�õ���P2ݙ u�X��4L-Z�C#ұ8�V*"��Nu	G�m�6b�ÕtV6�c)��ú�]���xN5-�h���JK�Ypj��EB]JSE^���%�8ªme���Z]�eҮۭ5��v�2e��բ�N�-b۱�Lw:-\馤���ZKm�e�$�^ZB�K��l@�8ٚ\�:ڹ[m]6-�͵!�i�.��]<�Q�%0�bQ�SKt���UZ�,�c����(Zf��9aUmpʲ�jk��z_A��fJ�M���v�n�ҥ�mX�n�3�n�-Η��8�˫��4�V��a5�*jl�2h���g�(���[��s�kZ5�QUW�UU[��s�kZ���(������۟� Ҫ�b*��*�wv�ƴ$�ԑ���I4�J4��a�����a�<t���\jnf���|����o[H�v�����)�i���PeQ]�k[�챕����2�dJ���h+.P��r��.J�a[2����{�Q!j��kb$�RgJ�^x�&��cZ߿q�Y=�:�r���֒��df�U5�̖[�Ԙ��jg��֭&�:�U

��\@R ��D脋�Ү�Mxm)M��-śmn�	q�t��C��ٻJKlKE�m�\]]6��R��{|�a�.\]i�i�덣+����]�Y��Ă��ԣ{+-n�޾��`j�2�*�j�GJ��n�`��u�Ԛ��]�1�]4ֺµ��ڰ�L2�X[q��fՓl]���kq�ͦ����2��3�Ԫǖ��m�k4�� �f&����2H�����Ŕ�;�Zm��B��L%Z��.�f���m���6�S/CE^%��f޺i����6�V�I�t�����X�m�Md,�TN��C�����Ä0bd�8�b�������v���]vg�'�W10�LG�$���x�^�������0d�H%������1HS}�Ap"S1CRt�B�-IJOt�D:���&�\���Љ�˫:�揇���Ä�I�r}t��GߣK�I0ؖ'��tDL��	���e�E�\먭zի�aI$���=~�hë�#����)��h���Ȩ��'�v[k�A<F{V�x4��y��r��:�+�$A��"��12��W���~�( Ŋ�%�<`��I&Ƙ7��%���ȋ[�KX����j��7
�'I��YcNQ2_:uJ��R���H�8I�K(�D舘&!���D�X�I�J�	b�4���� ϼCM6�x�$�s��gs܎\����b��і�gU��F�Mp�����ZR��R�8�a|vK-E��Z�F�Ø�.5&*$��R�XS:{�\/�*/˥���J ��^q�3����66�~(p�7��]�6��D�Guf��`�!ӆΛ0��舘&8���`�����5@�$b��j���97��bva�i���	�&xx3���iQyqTo���̒�b��5�=�A��ѧ���M�]pɚJI���A��u(@��:�l��1��0��;R��q|�%��(��8AGm�!A���oW@�Xۓ��i��I��0�舘&	��a6L�KIL5f_c>�~j�̹KЦ��c0�o�I�v6h!L����ͶM�QA��`����o[ fDo�����N�*VO:V�eUN���ݙ2��ULծ'uDuos��O��q����ŝ��C�)ř�]�e����a�Cڻ�A�}���۔�Ʒ��|~���Ώ,(5�:�z+VV	(�*&j �n
�Y��l�^.͢�c�*H�,ͻ	"��оn�O8O�%�j���h��s�O[ѣ
R�'��L�6��imT��CL�Z �!�TI�<�<�zM��A����O-�R|���-���7�$k�Z;�I�J��!+y(�FƘ� ��J;I�a�i�/�%�N�^+�캪�RI��Hx�g�Y�舘&	��!��RL�+r���R�J�t� �w<������b �����:R:g dZ�n�-x�B-�
ԜF�i��j8xV�z��3޺�J����Z�=�Z�.�غ�}9X
��+�4�AQ4�^H$�)��HXS�hc���ϗz��W��L�&\(q��G�h������!�9����e^���GI	:CgK<"tDL��	�!qmL�ބ��	.��<Ի�LО�ݚ w�`��&�b��w�p	6H���2�s+V���������x~8p�U�f�S��1��
G�t/W�Y4FDD��K"`H��'�A�da{�Po���#���&�ޫm��˧bm6�A'42�o�����*9�y&E�ε9�a���%G�Iц����\^t��i'	4�ƚt�<a��pѠ�ε�y!i��)��x�� 2#n�Y�{�&�{*zŴ�HW~�y˂06�D6�2D[a��LW7�V\�����1c<�����ӥ�g�Q����<�!�r�"
�"�K�!�GK[a `���s��C�%b���ç��;��v�F."N��.�8x8�O��È���:Ce�0��ό�"`�8X�G�a�/:?%ٕ�^0aU�%L�B+S\zSMs�^npX*W�TUH+r�N�5P�Q�f>		w2��rx3�CR������$�Hb
��Q�)Ǧ��%�=ѓ,�n�b�û�^Ã-�;����U�Y��c{��*���Y�X�츊V�A��T�h�
{���(Um����\C� 82Z�XD興	P�4`�K0xۈ�G�^%����<j$:�q��ueJ#��o8ǖ�h�� �%i����jѹ�Ϻ����В6��s��Uv�*��t�5�E"Fx��h�C��>�@��K���llzJ��K-puK�J����G,�Oh@����UYd��R�F�Xм��a���Ϗ�����`�<A0�:l�\ʤ�t��5D�I����<5pc4#��-4�55�g8�Cq)W�Z��yA���0"d�J��:�X��SD�,�F3��ԩFx@�Õ2�9��A�� G]�L�
<����o-:�t�f���^ˋJ��c�� ���ظ�1I����ogX~^����GЏNH_�,�����>��2�6r��H����vi:=GH��l�4zIl=#����ޏ�4�=��:_��0�2c2�
#��M!�[Lѭ��҈
4�MєiFw[�����4����� �	=���h�=0�G����z<4��f�&��hQ=N�����x=,��ih�4�F�Fk~:N�FQ�h��@hη�P�kFP�4���=�%���h��4z=4�:DA��4�4�:=,�����p�����pz|�P��m��t>N��&����a�U�^va�D�QxUG�Z/	����0���4��ä�����:=GH��3H��$l=#����٣����=�4����0�l9�f�l�
#��0􈽦=#�9	�1$#�WĂ�y5�㯾��v��.���9�Ɵ�HP9���F�l.Z�a"�R2�2���|����u����͖in�]�wy����+�����FYl�J����؈'hm��5�.�\�^�-� �� �yH�L>�cS��]7��1X����|��4�0Wf���Zm���le�Uo0v�/d��6Wr�p��f��q��3O��ك��_�v���e��#�� \��g����EUUE]�뿷�Z5���ff}�,UU�U�����4�Vffg�b�U\E]�{~�37��������Uqw���!� a�0�f0������	��$n��*��^/�<B��G�O��"�Ғ&Ԫ�pr�!����N14�$�:�,��htA�Jw���C�O$6Aߐ�ͬ�mJ*&<�JK[Onù��)�&`������B[ �[�2�0���-QDCO�P��EtHe�c|/���͌�"�� �TW�
�O��s3$��f�M$nX�����6�ti�TX$�t`BxG�����{���>8�K�g5�D%����鹪�k�P�M�q�)L�о���	)+aч��AL9*��4.���Yc4�O|Q��O,�g�,�Fa�<t���9Q�"&�x����@ ����C������/'�0^M�m���d��]a�O��A�h��k��L䴮#b������qH���7w�G9�ra�I�aa���@�1�9�u�: ���GI�/b�šw�~kY��]v������Qg:M)�d��=���;d<�^aG	�A�aC�� �F��[�Kl�E2���s�g�,�����<e��N���TF������0�IĞ��y�vA��4N�a�����:ꪽM' K�p�:%xc�]$�#A�JB鄚I�F�|t�<a�4���Ç���T�r�l�����Y~4�}o�<���n�~�1*����+�z��9HQg\��S͔J[6{&f�V4�3�I�I������+DJ��P4������*��a��H�/�f�*��>T+r�YfЋ0/]^E��YZ%gg>y�XScFuk��d�P�Wu��AL]u���+�x��et�V�����ѡ]������+��v��1��dO�s$c!1�|p�=w>�Gg�m|�B�iM0�0i����_"v�b���#͖#�F#�!��9 �5#�.�tK�C����!��$a(�J�����r��j�E�p�UPrX����H[�=��ѲNH;>m�d�A�&�NMa��w�=��AGɅ�J���P�b:@�a�u��r��,/�l���d��$Zd���>&�sX'�:�30�&	��Z9�UP��4�ۆ�ܮp�-ii�
C �H����tadT�P0����Pbe����(M�<40��|a'ĖQ��DD�0O��g�����;	eI��� �HK:n�N���	u�0Y6G$�d��*�DH���짧���)h:_��B!UN���ѯ_�w������:I;$Oz���i�l%yH4`I�/Dw�UUӣ�Ӌ�ǷG�-Y=O\G�����H�F|���R��a�L����`��ԏ2�Jr��% W��3K"��^��Uv.QfL��S�U�P$�c���x
 !� �LC�!�18(��8�фη�R
*����!��6Ȟ�4'$$������cF#�	��XX���h�K!�(:P�<I��|p���xDO|%l��+��{��Ա�i��i��Bź�
��'���jM����e5|7��6�_�/,��������ӓu�H�	۬B��z�8�86�'.s�5�� f���@�iH4u#CbE�C=K�5����	0���ə2I�FEV~��=n�)u�IGxWk��'I�$�Hm���b��A�W<�˄�rNXo/l��E������.��1`�Bf����
G $a�1|4����Q
G$����vƉz!8Þ�Y���,�S��QHi6�|��60�N�Ǝ��e$�`�D��nӀ蒂����N����'p�O~>?�`�"'�	>�6x�L�p�p������\�:qe��'׈s.�b�yH~�K��Q��pb�:H4Ƥ�0$����)K���.��*HA�JG�Ӵ�D编Y˜Dk8�/�z~�� UYU�"�I���!��XcL�!�Gy��f$�Pㆼ�8Ht�Cgʍi	���p�=;��DE&����iJ\!4�F�O�v����G2r��IهYM6[�IjH��"��|�e�s8%Nc��6Y���NP�d�H�)4���8D�Hd�&�{#�O���v�i�	Y�6Aك�>�1�Ӌ��|$����A���rh�LO\C�LH�m�R�H1D%���p�O�0����0DO|%x�Ts/|����8qS���6y�ȇ$M��R�O���l��r���2��q�D�n�5R�'������C��P���BEg1d
A$A$ڗ-:���bB�څ�I�꘴�Z���Y[ƌh�:]�lY}�f���uv�W�*�S����t���*���Ż���ۻ��0����"���ԛkAi��
ۭ|���u}۾\{h��%|=�Í��F���U�RT� ���u3��G�J f8�Tb4����7{La0�\TtX4zۀ�$�R�PG}�fd�oBT�Baц&/1�4&��#�^0�	~�pA�F�ZX������Ga�u��-I�;M���Xd�,�l�_77y�O""*91\x�:��KH8j0m�`E��MG|����������2�A�$=�%�Ũ�2N�)P�]$��1���4���f�Hc!g�Ѣ	-����ln�;���q��x�e\x��&�M�8<���1vG�N%$HQ��E�qs��&�'I��h���f>>8|~D��!���01�W8	M?2�n��
 ����h�ʔQZ�(>C���D-�K��{|yO>�L| ���%�����������F&n�y���	�FgH�5K�AѬ>d�A��pN��4@x��"v����Ih�1���a�
Ppa�M��.u�ѽ�;�C8� �g�Y7�"�Si&�FhU:�>���^"��q
�ãI�a��Fӡ7�s�t�i����A�3�I�ُ|CDn�'c�8u�,�4Q��IBi`x�	�g��8|~D��!���gF����y�f-y9���:�u�\@ 		d��Wꅶ��ȩZZL���\{�2b��;���s��'/g��n�q4�)�4b:L!>T�
�$A��i�G���ys^i�29�,L�o6%P��8��
�e3�9Y��Q)=�nʉ,�ͯh</�\P(��I��)9_���~�ᘎ�H�D�Q������a���A!��Ӈ�7KȚ�M,%|�VJn1���6p�u��gσ��K�t�(0a&���|��9pM�<-e������%J��6:��v�p�pa��O���3��p��!�C�g��N�DD�<xHa��x�5�D�����e�*P�$��BY'�zS�ghq|T_����<�� 4`�E�11�d��a��0l��ge�k��%+SX��LrDȘ��x7�1!�g�i�#N�+M2Q�Αӈa
�:ID�T���`�D�QX�d�-�&{�t{w`��5�|���u& t>��1�� y��� r�Q�K�L�FR0�,1�HcRs,�a�EF�M:���$�҇��i>���I�%/�D��=}ؘ��:UM�!�$�I��D�-��\:��H(�������G�.c�t�:8?!�1���9o�>>��i�4z<4�#F�#Fi&��4}4��A������A�H��}�E�O�^5z^�O��^�3�H>��χC>(�G�-1��4�F�������4��Z<�H4�	4�M0�����G������~,�4�=�I4�p� �3G���� z=ђi=|�=����xi���g[�)� ��|C���r84��i2i3Gf����ä@��A��H4�4�$�4x=��a�����4| ���4� �zD�I��$��n�*�0찼(�
#����pi�ѭ��G�p=�����=���=r\�f���M��h�i�L��x=�A�H:xg$�Z/
/<6Y^5�Q�D��E�D�G$z��Pza�Q����W��*��6�/P��N�<XV-������ղ2��ِ�u'`�mM�}��a}r��U�9=!R���6�6�׌1�5��t�9������撫S
S*a�i�-v�g�eLְn�\4�;=%!�y�6e{9����Xa۞��P�����ś5UCF�#la��RĔCy[k6Unᮥ�c�PP�i�>�Y���\�V�m\/�A�\ߞ��ER�A��ʙ�*໴���ν������Le��j�˜�]����ƹ��T�e݋t��Kv�R��-�@�L�4�F��ˤV���`���ښ��-u1w��q����aA�*���W��H�-m����n�.��q-jS̅���v��˵V�>)N�u@�؄"��1\�U�A�@Y#CLԴ�Z��U�bͲ�[dmTJʙt������v���28T]u�omB�v���t7g�.4�lt9��#��n����k��RQ�5!���N�V>�GFh���\��g=��$������~���������39�a�O��{w}�������fd��o��>�����ݝ��ݼ33&fs|׽������df����M�ə��0<3ǉ<I�D��!����M}�O�b�\�qK"�!��X���L�l���lB�]�Sq(�6����ۜ�`�69X�4q���]A�2c#3K0;V[G��X4"�[3�`�q�]^G �f`a���+)��Dь�S�	\뮸�X�%*��n��i�4͖���5���2� :&�t�+Fab�0�Y�J��ZU��9��٭�awZ�	M贁���\�6(��-*�H-7t��hQUV3pjM6Q�R��[�V���U%��l����CZ�-�Dm�U�N��laP"��Wh^�Mv�Zá,#4�܍�)n��lh��U��]GM�̮@��:��`��ue�ݑ��F�Gk�AQEQ�n����&�%��Q�U�yDlT:�A޳��ۻ۸���
YS�M��0um�dڄ�4�����l�,�k�Kܳ`���{�WɅmz{E(�]��}ᛤ��6�~!����H��%�HHc
C
��m��4?u�j)T�o�E�����a��!Q]�a��2W�R4Jh�T�t�o��v�㣇�la�h�>!̇��ZM�o��,���x7a��bS��7�yU(e��8�ux��ACB�����X�!�þ%q:F$���9��ꩵ�n�i�/�C�W�:�щ�a��': �{qo�pm�/�\�͵#�ح����.�z��npw�X�GL��A��#\E(S0I���)1A�aR:AУd6xقp�?���"x����ic^m��l�%�d�#��wvYe�Y${	:>:v�aC:�'1H0����)h՘]=1'0���h;��gpA�����-�� $�آk��a�[K`*x]��l���i��Ȣ�G/�d�����veE�2va��u���L] :0�$��`���݇3?���XB�@����i�^�HI�Ӥ�pq��3��Z;91ye�%3a����D}�m�F��"0��Y
�c$mi�ID���A��E,aEU�M�J)��ڀ��&GN��7�]VI!�&F�q�����	$�r�p�'��w�tt)h>D�%�Q�)@�
6C�M��������DD�<xHuu���%�b݀��`@ڲT��d��0�#"��n�u�lc� <�E��QɄc�ˣn�|�4a�tH�n�l窨�x`��֓�0)4m��$��dB�%��Ox6>.M!�*�A,R0"]$	:>tKl4ɐ[[��}�q�bfZp�Q##h៿Kf�әm�-L7�>c/�;MH�E��ݪp�����("C���pA$���F��ыG_32�ĝ��F'!cr:���Sw�{�6�N�<�Ds8�p�����cɎ/\bD|!��������a2x�`� h��"(�h��4m��}�Lqz:L\��kɐ�plGFY��I��>:i�"'�	0���GT���V̕*�,�!4I�=b���h��Ѩ�4����ւ�Q�8A�$4GH�;�O�\/"(g��I�h�t��BW�8�`~mB��7t�P(��!ӳ������ܽ�g�<#㪛�)G8F��T�K�~̚�t�m#�Mt��u��r�3K�����ߥ�i������r6C�L����r��,f{qr�6�ve�e���8M$sݤ�TQ��������b�J8p��,b,�1ч��Ԕ�f���Ӥ� �9c�<����̸H��S	O���4�[�/XǓI���:Qbl�6"p��:|"`��<$<xe�X�<�c�v�aƾ���4�Ր���6�PUqЧQ��;��Cm��ۮ�TT�75 �����UP
�Ѕ�c�$Ж�y �)/ە9��UM�^��8��~�W`�	��{l�}|�Ga����v���`�};���w�6���-�su�ţ�}����;��ܙvU�ҰT�y�{,0�>sa�T$N�W����vѭ��mh47`-���nm|tki�5���;8Þ���Szm>G):M	�0�|�m��V�+ZT�(]�j#��_	:P�$ai�B�#�N�5V� 4!rH҄0��k�ہ��Ltx����.<�a�Dp��죁Ĺ0̓��P���gBQ2��0�r�:��|K�"
h�0���I@�<�}dV��x��l6i#�&�5.0r@pa�'2a���]���`�(4N������ ��0�
�D@�w���T�ăq���~5'�i��1Er]v����]��\�|4b*P3�c	�@P��TFᴸ�A��L
QL$�O�8||t�<a�Y�<xe�X��,݂��|��[V�4���1�bMqLO?'�ivl��vs���<�;4�����P����R��$�% ����#v����6��n�K�y�s|g���:#�ܯO��2|>UǮ�=y4�
L�T�#Y�I)P�Z( (aw��
DB"�-���
;1#]��f	���h��;�DD�I��XrI�_�F̝��!-��M�J��m�����x� ���=ϝ����$Ժ 27���)Q6�a�*,h���Ic��*L]�%�"��w�qZ�G5�R]�vA�=��ђiB��
BS��� ��G�0Ç����D��!���}����\���81�c�BK�I$���p�R�p� ;(
�>\��(	�
^�t�#G��paHa���ꓤB6�%Ģ�)}ѷ�R(h<0�p�T0�j� �(G�U
T�
S(���	T��?\��(��_sO|8���$��GH5yB!��@ȅӊ	R�	�J|�!0�3-΋�Ж�>�r"D�22%n��{̏���͹��� �%u�F���u2�b%Dm6b޼���0�4A��Ǔ=����u]��5&�x�
�w��6>��G�:E�(a���6D?��,"����z��L�o�|M:����ģ����B�	pjd�qP��p!�~�@�a'	 Å$�N>0DOa���ٽ�J�v��#G&�}=}ZR��,����0��%t5���4�	G�bz��l��×4�DdO����'�m�d�<[�D�PO��G�U�f�-q���b�~[]YFI�̋)'�@t���Ƃ�D2mB��}��ceR<��@���=qt��g�u���eɤ�����",a�P�$�F�SP��D%��$��"P409��DD3$�$�]CJ����(��b�)6�8�M(A�O^0�	tH�u�:&�tm��ѹh�=qDW'L��8ǝ|�1�KsD�{��8T�P�4�g��'�ç��`��<$0�>u.X溮�p�o��V-�n��,�%�*�ZN��nJf�OYh�a+�)��uq�LRj�Ë���1�bH>�ԾpM]jk��<O=O\��;��7�^�P���F�x��Lu8�o�oWfJ�Vn����O��'L�{Aô��'Pm&	Bv�����.����13��1�@JV[�>kz��oG+�xq��(�3���$�G��GT�K�<5��ZV�gM/�I�D�ߙ��p����Ra�9cLv�u��^�M:�dbG���A�xq[t�޽�3C.M}]�֋%u2�FW$ta�֪*��F���1::7����;<u�"0��I�\$$�f�"$8I{NO�p���LD<��wa�`pA�pЦ	�HG	��.LL�8<t�%$��i�$f/&/'i�̟A���ƛo�b�[Zi���'�K-Vr��8��LS���ތ1�0K%+piB&#З���G���0q):�h�(��H����,K>>8~>>D��!����*�H�%:��oHˡ4ãZ���͌c�$З1��Ф��ҕ��D8��qJgZ��RA�N;!tq�GG	��lrvc��=d'·FY,��ؿJ�����4��;���8�i�+8�Ar0i4�!�:8���^��ME�M^����q�Y��0�@hra�w,��x��XPu*�@� �IR����嘪�HB]����j;,
$c!6Ҏ.qs2b���Ǌ&��.���%&0��ڛ�R'l�j0f+F�J�lwH��쐡�#��M!���zw�M�l��,`vi�RG	PÚ�:P`�Q�B}4���W�Jh�H!Qѣ� �� �E�����pzL=6^�����=9N#�l������?�>#�������������xי$x�QG�>�F�h�ѭ҈Ti�pzAh�њ;��z3Ɛxf���<= �L#G����A�3������L'ñ�iz=4�4�4�:F�F�Fh�y���G��Q�G���f�#Fjm�c}!�B���!i�G��zT6�� {ƚEF�N��ƒh�vp�����ɤh��G�����#�H����"�Ђ���n	DI!h�A�VxUxa��
#E���Gђi���H8=�k���'ja��R%`��8FO���٤i���tz>�F�L������m��H����oa�h=m��׆GFxQxQ��=(�LK��(C~���օ��U���v��Rg�/G��T(J��R/Q�	��ذ�7D9;u��ۺч�&��+q�v�vس[��YXxv��w-��4������-j�vS��CW=���Vw���C�n����W��WrN+��lZ�L�k�3$�3�l�ѥ�0�S�dGgT�)��B�*vw0��.��0��*�^/�}}��7ﻙ���n��u��L�}�S37����V�W���}{������f}�Uv��~�������s32�3︫�W;��wyS;ļ<3�(�G�4ӧ��`��<$0�>��ʕ*T�P9�� �j�_�j/�x@ \����!�A��3i'�$��e�GZx��P�J|���+��j�8L��;u�/��L%��đ��QR�#�
�g�8�@X�|�_f>� �I]�>�5'�^��4��C{��ͷ}�4jT�����{��Ƞ����㣽�9��4G�u��tk��H��@��(�"�uY��m��"�Ms����zGH�ll�J`P�ζ6�J9E0jO	��()��R�I pa긇�8`i^)�q29"�}��1}�6gku��:3�V}���Q�.�1�_[�Bk��R
,gJ8Q�4�馘x�,�x�./�8�� X��!Cѡ�m���CG�O�1�
�!z�!OP��;Ѿ�$��"Wa�:�8��"ض�t��"���q�D�nVUE��E���B9"�#x˫T�2Z�x�H�
G��1��u㤠��p���KR�%g�"�qH@H��d"�mdJ)����+%|�P��m#���!��6�0p�BS#-J�J(�m{��JE��Y6� g˄#�Q�j�p�4�D�����;�k������b�A���<Q�(�N|t�L<a�a���i�^� ����lmKR�(��5�느�7Gw#L��Wb-`\��e�9i����i�xr|���݇Ș�o�7���ؗq=y�	��Qm`��R	 �	/Ke�Z�,���J���_�zt�{&_��tm��r�ά�Sz�3�����Գ�T�^X�9���g�W�ں���S\���ަ(�U�]P��U�X�Z��㷜��{����n�j��F��	D����L�Rh�T�J)b�Ao*&g�:�aј�~q��$�E��R-|�����<Ӿ�SL�����N��"=(���xd���tp����"[\E�GxAGQ��7ôp�>��c)UdD."��Ǝ�ꐡ��[H�^���#Z��/��X��r5dr�hd#�)Г�x�>P3J�J8q\s3ki)3I��B;����mr���8�e�DP�U�y��\���+��:gN�F���DGf��'�F���8��Z����A!��FY����N�������D�aL���fC!���^m��m��&3��D}I�b��%�&G#�����ewt�$(0��|�!8�H�Q��G�F��E.��<���#�ԯ|��*C@Z��"�>�w���N�b�����������2��,V�( g���Q�HZ�Q�g���3ض�!
����"����e��(�Z��K6>}ȃa�QB��	P4I(��"%�ff�vu�c��%�	هǱ٤q��U�
J�zY*���=�bdB�K��|q(�I:I��:||Y��x�,����,��7'ò�z�Qny�X�N��Dͺ�S{�@ ��ߓ��Tq�4��.�U�G#�Z>k�!-0!e�3�V�=LN0,zw�G)���Qo��P���H�"��m���HMD ���2�ίÈ�[Ȳ���(g~�K������ٿ1��6��	G��!yI$��dJ�|G]8�]1z���ʔj!@@Φ������x��x��zb���y��z�'<2P��(���la�)Z$���Ɂ��&�'ZnSF���;��tTZN#�٣I���h�%	D83$�N�x�Śi��0��<<2�3�6C���N:�%��l��h.=~	D"Z��M���SJO.�.�6Fê��ON9.=���Я�|u4�-���R��UPJ��y`΄(F�jQa�C>R�>C�]��b�}���2�����")��(���#��e��]/@�������S�ӥOw���:�]CE�J�M����#���8��,��%AP�(e�!�z�qޢ�CGǈI�k�r��uE���C3���L$�f�0��4�Ƙaff�Ǿ#����ޙcNX��E$#[��n��{O�<�k�L-�VDt,(�!��'��z\�?Є=Ӽt��4�Z��DMv7V�������Lɶů��c1Y�7]1�+��WsBƳ����30Ѧ2�`��O*l�B����y|F�.���Q�]J
�J�BA|/ߍ~��;����1i�>#N8Hpe�G<���(���s��{�*��$�P����n���:-�M8���<,g����<Y����K�#gN����Ȅyd#�9h�qy�3�!���q�H�c�&Έ���p>�	F���G=�WVZ�k��K0)��]�i>8|��Y��S ���/ʏ��*�q�Y|I��N�|Y��a�Y��ǆY~�,h��}�{�Ү!�5����� �q ������F�p��nh靓�t�M�H�C�!?+2�wv�-���2-1<Z^�� �h*�+:�D"�M�Ԭ�a���>m�gǑ��P���7�s⎮~��������놬���H���F�r'ʈ)p a��Rߡ�5b�]\��~�]GW�%P1�h�'e?����X�
�� �ƒx�����O��4�0��0f�`B]:���Q6�R]���Z	!D"G�����X�MdD3�:2��9
\-�&+,�
�fp(d2��|�vp�����M�k�>�
�d"��  da��>rC���8c�	r����SҔJ:a+N���oz�w�̃ςP�����!J�i������T����/IP�#.4̰=�Vgi�!�OnF��gش�ixm<BBr.�5��:a�HHYd�aei����f�|'�'����������L��,�c:Kgѽ}<����@ ��T�(���p>,֏��V��˘�+�J�v��?m��[ XO��&�ǼZ��Ȅ,IU�p�B��·�j�\<?"h�єq�pgLs���8J���8�Ը4�h�O�u����~���!NZ<q�С���m�6�W�J:�D��>Ez��ĔÞ<��pG�ЛL;yN���A�.��8?�C~�HѳH����N�G����~"��d�����i�4z?l��0�6��n�k�9'e��#��0��|(��63F�h����5��G����>,��A���xf�i�/A���a�0kG��0�4�4�<;A��z9�Ǝ�:N�M �`�g�ǣ4�,z:���z=���������1��Ϋ�K�6^�˂���҇�����4z=4�F�M"A�l7=��H�n4zۣјia[�8x��Q�1��	4��So�F>�0��/
�"�~��S�>�Ã9/�<h�;�q�|?����Ѥ1�= ��:F���͖�xi��x�m��zGFpr=���Urc�Gg�E�Dh���Dh!����`޵���S
��.��d҅f�e:P��@�Cn�0R@CF�ILi�18��#H��?;�T�+%,��/`w�������,+w�20C�?]��mE�}E�G.�U�sv�˼L��nXC���[#L�����gF��	�۬�v��:�Ò���%-a;�l��力L���*躍�^��'҃00ڳ��eZ�lmΫ���Y������w�0V):�TN�����+��쭶LY\����)b�j��I�f�ߛ3�icS�p�Qc5N�뺵@�NS�'VM�:ڗ6�U��6�$��?+&V�Z�ґ�X���p����{����C+���v+����vI�.l�I�վ��\�Ѵ��f6�n��ԢA �:��8�W�D�R�r(`!�6���B:1Y(��\
��cm�ꖑ�3F��3H��~�_MUn���{����� ��7�?qWj��i9˿������}�]��U��������y���UmUⴿs�s333��}j���V�����k6Q�a��O4��4�0��,gN�=U3��5�Q6��V&�.vGà2h7I�l��B�j���
�ަcq"�ֶDKk1f��m��D%�mbhJ�,�(2݈���W4%Gio8�f-�C��^�,X�q���lY6��3����:&��\R�)�����Y��ny�s%�q7i�e7;�.�m�XM��6����l�v����-��F%�J�b�v��k4q[�&iyҭ�l���z�nuq�
�_�k�S���3c��6]�]^�],�6֥Y�����3BSK\# C8]^kKk�o^4e�γ2��0�l�����#�<=s/bͬ�k+x��-�RG:ѷ�����g7�D��M��]%1�[�;b�2Ʋ�3:2���1-4��.$��@ ���ޟ)�딻	�,�z�	����^_�;$����0�c,AA�����G�u�&B¥�mлV�$�g6l��f�ʡR�UH��
�������p2QD%f£�%�s+Un�@m���21�[u�-�D#1�6�K�n&z`�;��4�7��!�3Q��T��td�1�'c#�FY�3|�E"�g�83s��2��:�AL��X��y�]#z�ӓ��|mS)�W����$�Y�9J)k�
ֽ=��0�8���D�
V��W�ш�!�Đt�GI><Y�M,�M0�L,���t�3��l�YJv�@Z�ZG��6�l��@��d�bb�۳QjW���;�h_�w7�+�J�^��&1Es��><��G��>���((d���/!���F�E��!�����%�^����(�h>G
sP���Jh�nR�/�JU4�	Y�����jJ��/|i�[��]U����'����8  g�1O�J8skx�%e�T��1QH�H�Է!����ͱQ^xZ�t����A�H,���a�Θ|Y��a��Yae��W=g����	J��{�� �D���"˴�b{���={M�yPϨ(e�Q����p�f�c+�6:,�\u��bb1J��Py��a��Z�_��u�YA!2��0�7t���!n���v� �dzR>_t��t0i3�6��1b-�j<�B%@xdB�ґ���Oæ�⣝
�#�u��N���G�S$�RJ�pS0J��zx~���^%p�6`,K�~�,��0%�)zW�Ԭ�PIC$��F�|iӦi��i�XYc:J���ʩT����3K8X�~! �@:��v�j���mH�\-���K���S�o��&���e��N5kS��+�,�M!x����.����a�'+��1q5
]��oHϑ}��%:a�H���D�x>�+�g*B��{�%v"+R0] �G�ܝ���PUV�a�0�A��I0�� ��pgN�@p�|J*d���@��Y����F�|p�c>�CBN����aF�t��i������$�m��Q�t��䮽��fU�nB��jUs�z���b�V��C�v&�]�] Dw��@ ��ϯ�Ӄ�O��U�t�XJ��PZju���X�*��G����y���ݘ2�Yx��@���]��0�k�����6]�v9s�Pѥ�ʗ��:Gay�P|�>��2�cp2d��7L�!���"BFu�T/��V���	����r���>SR�qtΒ���U��Ҳ�h�j!i���ř�~V�Y�	Y�ⅿK#�=�>�
��p�����vn��96�n��:s6�UP�!���N�)Ch�tgNĳ�9U�:�auS�`����Q�y4��$ $��((��>4�M4�M0�����?K�%�%�z�bF��X�$-���H ��@�M~QҔ�!u� c�m�����S5]cc<�oN�P�����u'+��h�P�g&�AC�ꡛ��8�D�ـf��=m�(�Jh����:ˌm��4�[>^�_��B������.����(&LĒb(�\FaO����!ĕ#��2#q��x�('!�׭_��ktPpa��	Y���a�1WJC��F�iG���4��M4�M0���Ҹ]����d̪���4���i��i���\O����3OaǕZ�������Ã=��|_`������(d.�Ih>��F��41uCX���uÃ0����$l��?7�찖_�b�c_&�>�����π<���8�P�I�D.HP�D�������	*�����}�ψ���-�F^��D���t�G��d#���$g����̓|ɦB���Z"C�'QE�iG�:wG�f�i��x����8���+N�?Y��R4ͩ�b	 �	B e%��-���tV�`���pg��B����EK	q�`�
��DPnQ��u�����U�L9�b��r�"�΢���ۋ�A�ii���:���4�>��I��@Pϒ�"!7#�;*��z�ܯ2|2�D���f8�UWQñ��O�N���ZYJ��C��ѥ�CD�)(g�0�J0�N�|Y��a��Yae�,lf�a�>6"XS�n��	|�墥�vM��V�Չ
p��5�y������������A$^e̷�Gh�o����ᒃ.L����`�d����ܘg��ض3ZWUh[�R�TֲL�f<��jEXVV�Q�N�QeZ4##)��3d�nۢ�~�լq�$(�A��y��uq������j6}Sh����|�ӣ�Gab:p�3ſ����b:�#�!��QMq+�k�����TZ�EV��x��ؗ>�{�1;O,;#�(�*�#B��Ie����(--�c�����P#?�MSlӉ���HJ��R��t��	�A������IjN���]"��y�I�b1�r�L��J׉X@� �F�YGƘt�K4�L4�,��A������	:[����������� �D"��IGʺ�8�zR>+�h�FXH��Hy.�$�HT2��f��s�w���X�"	1��oå�y� �r��#�t��k�(�������(!C3��ǈ����2��F-a�GGd^�Q��GI����w�t!P�,dY&"�D� �Hpdȯ�8pF�Ѵ�F�eLQ��,�,�,��l���M���<lA�b"0DD�8'(A�A(�H�&ı�X��`�a�`�&	�`�0؉f�6 ��&aø=4�
<Xi�$�M0�O�%pH'�,K6a��DK:"`�xK "A,DN��'̝ΖlCi(I0�0�H4��4t4�ؐHpH"x:x�㧄OD�'����&����e �pA�࢈|~`��ܻ���(Υ��%-p�����3M-+6����`|s�*��t52+���kj�����@�PT��=s��:�<V#eip�Ĩ��%,����J�BG�U5r$'��om�u�d�A�zr��i�>��������5�am��Y%UG�Qm�=�ti��%�$��7��V㳏�'C���U̹f#kHh�f�^�Wv6�6�Κ3��u�Ӂ]N�}��9�������q��[Ux�-�˿�333��}j���V����י���Ͼ�V�^*�����333���U^*ڮۿ�l�C
0Å�Y�Y��i�i��X� ���s�Krۏ׍6�m6�4#^ ��I�W�s�4�ccm��@�RJ<�¥���àx�����4�sUU�	G�Όa�C��iࡘ�2Q���i����/�	y����U �bu{�Ԏ�!�Xr��u�~� ��@�{�"q��PȂ
�����P���~�j��&���neM�;=N06G;=N͞�����|�����u��Q9�|\EZ�!%X�!O�:��A�Ӌ�(r��AӇ
0�O�,���4�4��,e�t�����>5������c�ܕr ��4��m��m�h_{2/n5�a�1 Ii���#�|I����u;~a�ֶh��u�[���j547T�J�q�T�q�.b��y��G�fk��>F������y�Ç�M�XpgʒF_<4Q�:2�u��ȇ0�Z9�0�c/�cy�����UV��<~'�{/��(�+�)�}��I�\Ga7N��, f���GO1�!HP��6�c(��� cG�!�0�F�i�|Y��a��Ye����l��N��j���TE2�KNYv�/�$�`��P��Wg2Uhm7� ���I�Ix B�ƄXC�*�z]�*�4��oQ�=�,��J��1v6ؾ=x:�ͪ��������ê�a�5�}	�&K�i˱F��IH=��]�h�Q�=l*���L�$��(|ъ=���N^CDi$���4�W��{fa��__Dl�b����"��ݾ�h9#�'�4�l����R5��D+�� ��-�˻�ٟ�יI"�9��}�a��e�G�?(
{�r�F%ђuP�P�Q��k7L�'${������m�@��-Ia�s�m�IU&���A��m���o�-��|{��ɖ�G (��3(�����p��A��p��Ǎ,饚i�i��X.&���|�!�do��&(���30��3�}��tD�q�iF�8e�Ev�|5��t�P1^%4��GǂO6�|��S��x�=�_*Č��\�|g=4�O��gKX�A<����0x�LY��m=Y�Z�%ui�qHp�7���1�]rTL��*�xH}��^�J��e5��v��4��/���h��^;e#x>!x:2|�m=ll�V*MXx�� ���,�ƚY�e�i�i��X� ��Xҗ,����Oj'rP3%_ۭ6�m6�4�L��./#�d�23����	�t�
$�>oܰb�-J/Qj>��yb9Hp`y�����Ѓ��/�j�M��!eu��H�Li�3��o.��D��)5�p�Qhv�*�OGW�X�����p�]<�ȲQ�[�7�Ir�I���!�W��f%��8�%�\Jk�Z3���Ȇ�<|Y�Qk�Yp�{P����0��pigŖi��i�Yc,��[v�b�/�ب����b5dwݍ6�m7��PqqWF��3B��4fvh���^����^�;�*�3��܌sWU��qoU�&����Y������;\�J1?���haB��#������H���+8q!�#���}G��<��R�Q��i��	8�G�xZ���$�s�8�:�q��Z:��mq���{��:pe�p�'(��>,�M4�M0��dY�eF]@�D���Ǌ,�m�pYx�\��E��n��)0��H�	 ���!��3:X���@ ����|�m?����Y�x�K��oi2��;[w��r�l˃�W�9T6����9�zj@o�83i��A����_��i� l��Ȃ���y �oJw`���c������%GO+*N#��:��7⎝F��oJ
-M�>��|lMZ��i*�ߊ
F��.�O�e٤����>�n�U52I������)����!`Q����e2
)wA��_�[n��Q�F�Җ�&˖3���#bb%Đ����[�z�̫]O9���>O��xclv�sㆫ$ޣU+a$���I�J0�K>,�M4�M0��d3|�L$c%�F�j[�Enz�" ��A�-%q����8h'�o���9���}/�F���Ԕ%�>K�,0�=7h�q3Hs�1����7������*E�|����>T3���<53��g��(wK�\@��ʐ����/xƥ�i(ֵ�U�"Wn7եV{@&�����Yг�p�J-]m����|	/��0L�>�7��C)�����0�����$4���a��gŖi��i�Yc,����%�y�
��I�Ix ��F��0�$��s�(뢅�
E�#�0�%�Ȁ��ce�$�T��{?#u�L�=o�AÊJM+8$ ��)?(�,�L��g1~x��B�3���p��3j%��+���TuQ��%J,���F������>��Qą�k �>�͒`�9$�q��y?��&��%!A�����L��Y��<Q��K4��4�4��,e�t�N��/m��6�3Q��[B��C܊�"����M���׶��/�w?>��a�t�@2~�Sf/�����c:Ѣ�n%�>!�N���^�q쁹u�9n-�L���a��2�*��cz�uqR[m��R|.��]�tE��"�RT�&�A,����� ���J�x8`<뉙�����ͤ���4|g������^SM���0�i�(�R�׎">F�(��g��i���T�"%x�>/�Y�e��� ���0�"A,DN��'D�<p���A؂"%tKbX���D�&0�0L�x���D��x�B$�DO���!BlD���4�M<pӐ<8a�
0�N�3H��""xD<lA�'D�0N��p�bY��ؔ%	DA<"B%	� �N�'��:x����><P�$�	�DOI�8l�AA�B�|p���'�=��I0��:�0�ݪ�P����\!YE�t(�:ޖ��Vᶫ,f���D��U�ְ�W�O.�%��&6��!��xɁt%D@j��,	�L��/dkN�Ge�^W���ݕvr��?)Xe6��oi�1SA�F���xHjx� �5��ه-dk�ASj4'F��dݡrU"�$�L�� ���)�*�գ*�AaS��ͫ-��g���O�먅��U�H�._�(/3ϐI$�J�k8�o/�̪E�{L�D��x��((�̢v�B�7 �Z��]��,d�Ԥ5d�#��Ty�[t�t�}�M#AE�Jεh��#(��	!@e��ke��`���r�V�u��	�]��P�+Hm�U��m~�-e���k�6�%�=c������)f&�f����kX�e*���PPD�9����-���$�z{~�wҹ*o:��;U^*ڮۿ�r��fffw>�j��[U�w�/��ffgsﶪ�U�]�w��Ffffw>�j��[U�w_գ!�a��a�ŚYf�i��ae�2�:o��\��U��^�/�
\B�J�+��hP�����n[�ⶳ@���ʤ �t���h%�Mճ8�|gͽ�5.�B���rB���k���LR��	��.�ny�D�(�ҘW\��w�����1>y�/Y�<��	+f���JK&�vζgCa�6�-���g�T|5�n��c��.kxٓ[[fh�5.��(�;U:aiF�jK
:�  Ul8���)�.�]+��W�Z��/��Yti�M��ȚTA�&�@�̵qr�2���LVˉs�tε3�ݖ�X��>�nt85�n"ĺ�-I	�[a�b$��`qn�Y��`�T��1��F^+��>�z� �u�TNzճ�R���� Bk����q���SV8�tᰱ��{�:�ob5ܹU;��fq7�uj�������վ�Mcux�u�V.�n����r��F�/D�t��.�f�͞"�Nf��Tk9��غ�)Rp���Gpy�b8wF��S�����-䮶ׇ�8��/���(YM�胡GϢ.f꺵Y��|D��%�EK ��{�F�3��|�3/����4u$�ۇG�F3���l|Wɀ�-pV@t�k�]K�C�"�00��.�A3�d�SSPp�!�����h��g��ȉ���!�L$<Iӥ4�ώ����4å�2�:�+܂��!��l6��Z�������2�VZw����"�"!B-b"@�7���h���d��I#�x��Y�|��|�_������l8=9HF"o�G��vY1D<P2��?��������.���I��MR�m��ͲfY����җ-0��k�t:�h�I�((��}�?Ӧ&�e�>m�7�1���	"��d�$å|ag�M<i�i�K,e�X9y۵Qm]�W�
�� �	 �"dZ�s1UFj�%f,G����lp׍\RY��1HJ\8w��|q<7��>��'��C3��~�^*���<�-�,�&S����A+F��Η�
_#W�y]��
"�uZj�yA��Ͳ	�Ԛ|�Pa:6���߸K��U\�U)Sb����*��$�>p��ĵ|(X�t�$��t�� �ĝ:Q�Ɩ|t�ƚa��t�Ƹ�����#�`	���^#M��M�My	�^��A��bx����* N�&��@�׼7ܹ��. F��\iԎ�>G�#hH�47ݿ�(����"���\n'����(�|�q�_h�1:}���s�QH�:�q��?p:U#�]�7���_|M@���ʪ�.���uT��ｨ�(:t^0:��j�)��Hp�v,����y��C%��2Ft�$ӥ0�ύ,�i�<`#�ӽ�D:�Fˡ*7�]��zz��|g�{���h,�A�8]���DA$^Vg�i=_C�ە�W�c\k;s��Xy3����A��8/4_,��u��7ݤ��ͪ���N��n��rWT�e�un�{r�Lw蹈x9���9ʖq=��gV�u��x�=s�M�J�;Tم�RW��
��7����#,p�C|^G�GCF5⏔�E���\, ;��c�C)4�P��G�5��$��S��V/�LN��	qYa�]�(:��1fy�y����@p���C��g�!�0L8)�p�e��wc��h��ń\|�����F�|���Ic,��	4���Y��,�L4�<X� ��㈮�b��%d��K��'�s�" ��A��kpg�8�\���$`{��zM'@o���q�f99�v�/SI�v���4iG��)�	}�qRK��U�5aŖ�2Q`Ϻ2IG͍��:���6���X��f|ν�x�ڋ������
�g��m73�#-x
F�2δ����n*`�$u����
�T� �4f��0��Y��c�eE�t��A��:I�OY�4�4��2�>�^_c��<A$A%����G&b&H�%�rt�iQ=E���T����\5e��笓ڛ0�H�3iUbx�/�q}�Ys�~�	�I@�kt�^�%v9E�\�{K�4��(Vj።[��A���T#��?������4$��dO��+�V�+�7��j��x�?�������R�0�4qZ9�xc8A��K$����gƞ4�i���쎌97Z��PY�\8e]�i��i�����ť��_��5

)yԮ�D:Wh�§&`����d�A���>>���l���{va��6I�e�fD�B�Ň1�)p�,�p�ꈂ�6Σ��G�G�в��2�2����� �&�|yq|P|8Gɯ/�̇#��'�A� l���J���Q��KNCį,��F��AG	0��igƞ4�i��<�����+FƑ;5�Aj��j�5V�fU��ܨ��X���E8�7kb�W�h���$�H$�b������|7h����pmf&���e+z��9ۈ�r��;]�.��Aq�J�c&���1-�������V8��9O��,0tUW����z������7
-IN�Q"Qg��~lt���-B:I��&�p �[ccoʋ�����Q鰣�M��ӈ�T�@j�A��1�v���Q�8��c��yfd���_"p����l����������v���E�O�:��8uD��k��fg"92��3m���Y���EG�{iE��E��Y'���x�� �I0�Śigƞ4�L4�<xe�ur����8��W��m��m�k��U�Ff�_� ���:�4����Q������ϑ�s�T�Ó��F%�P|mQҾ|�I�Z�;��쯜�CV`̅]'aL�ㅣ��ͱ�>]�sƥq9��!n�%�͈�$�l_w��1��'�߹�>�Q�epӊ�$6��z|�H:�`ϓ2�����
FY�b����x��g��,K,�� ��""&	� �"pDODO:C��AA"%Y�D؛8"tOd�0�`�&	�`�&pDM��
 ��""xD�4�`�0�8a�i��i��iF�Y��t��d!�%���H�!B�DK�`����tN,�&�(���� �$�%	� ��d<<p�Ӧx�Ohi�4�J4�æxDD��8'� � �&�4c����L�6,�q����q��C~m�q�F�!�!z�#|깇�#�ܽI�U�\C����Ӥ���*��1nܾ�2�:gg=惮����'Z�w��v����VO��::i�+�Z��)�-[uͅ��!��m�x�Ź8��LZ�{khLV�`�[[٤Y����S;U�b�����۾�/��Y�}�7����J��]��ws�������R��Wj������333=�Ԫ�Uګww}3333=�Ԫ�UګwU[�/�<߉<I��Y��4�N�4�Y#�	 �	/��)�q*�S[���"fH/�Ѽ^8�E�0j׃�X��8�<s!��D�_x����L��F��ucA��"jX���M�7������� �ί�	]]+��E�7$�a���T`���J(:����>m��Øg=@?	��/ө5i��N}�FO/�JaH����8qg��3H��ĘY�Śi�K4�M0�ǆYo��&ǽ�3��1 ��(m/���	�۞��DA�p��|����#�O��^:��
��>�g�0�?~7³DE�m�D/<��.w��t�ZqPy����x2�|Q���#�r��~��5�;�����ӽ�g/{|3�����m���ҷr��z��~3|�GV�$(�v|�#�tTNC�x$>T�[��g�/,,�����U�d�t#:G��'ĚY�şx��>4h#�y�d�R��T�n�U��޷�V�4䁦ɠMA�����~3'�O���[��ZM��k6�����$ �E����V��6�3���a�d�_>��q��r�4�����2�I�9xo/+��m�]��Y�e{^vEF"
���ʆ0��c,�l�����<�깍�p�0�(v�qB�dC<�K �z�X�.aag��W׃h�%��bv�~"��hjL���%�"bZ6Q�J;�XHb^�G\|���a���q,<���GQaFXƘ�h��RŻ��diyØ��D�1�U#i��ӈ�A�HuJ9��^äm*X$e�M��I,��|i�N�a��Y��,��f�CM���ؘ�^z�i �����6�m6�{1z|©���.vG�{檫��:<6E��Ĩ,��$��#�g�lpb*�{�.#��/�Qtj.>ӊ�km�G+�V�������_�o13&M�*�`HC����Z>��G�����W�s�BE�I� �h�`v=���*�
(�:����@�(�W�߆cm�|z(,:N����+�GM(�}��te�M�%�i���4�ƚY��ag��o�Ɉ��z"���M��M�Z�@�RW=�ee��k�L�&t���B�?Kv��
N�7y����t�|(��6�B<<�	�tg��_<#�P7"%%B�Ee�$���>|�qP��o!�ނ�b<A0q|����QextT*Gh��(*BHcm��ۢV�#ǎ��� ��nN�y��#��0��<G��'I>0��f�x�K0�L,��#����;�D�Tƞb�Ϗ�� �g�~�>�0�;�$�1=9:'<;͙QI<+��y��ǌy��iD�F�.^^y1#�{ǾF��K�P�l�!�aש��vU���p4��Z��Q�h�q���a�}��Ç����(I�ծ�����uR�<ώ��D,$:��x�}�3��zZ�"��5HI#:G�'Ěi�>4�a��Y��<G[������Sb�4!nZ�i�fM5�bh�(�L1���*"���x%䞮�!/�+�{�џ-�K7`-�h��t3�]>�ߢ	 ��ו�����ƫ	�����Wo8.�u�{�V9���9�}oc^.�i��m^Y�r��헪���le�� �58�¯v��$5K���,亖�<�y�LAN�Γ�j53�/�ŃO��m� ��%��uE�m��|r �-E�#����V|��G��vWv��uam����h��W��B���7�}�i��ח����$��BgBMVt�_˄�dv\7؈J�F6>-�����T٫c�x1�)�>�P�4Qg!t:$gH���K4��gƞ4��4�<xg��x~_[���6s5�?��.+8a�ш�P��Q�SI�:l(�u%��/bx��y"k��ثLHKd>3�h)#\6������yG�Y0�����x'����P4��;�X�t'G����珕����N�Y�ia��L%~&��=l����1ᝧ/�]�	�8rHm�J�E�E�_[�Ce#�e,Fx$�ψ��$�L><|Y�4�4���:�]�ʈ���O92m�Wo4Qm�쩅x
1ץ����M���͚���q��g�%��Ɋ������r�H�
�.�B�K�ibk�� -���6����Ί6�?#���_�m�ի�i�P���߇c��<7�>M�|�FY�����J,��Ih��|T�����`�����16��"8#Qb��DP�}:x��g�GK��X��J4��Śi�M,�M0�ǆx��FE��=��)b�R��~�(�QC_i(�uuO� ����'��Um-��vDV�`�D�n5��8�
ݕ�tcC<|F�#FN/��n7�x:�O�qG��FuQ���f��ʮn=�k�J&�řTY�G����+��~0��:�!y*GQ#H��g\����l��Fx!�ƍc(��:9�~8p���|�DD����t�H"%��������6P � �"`�(ٱ�؉��tL0L6`�xD�0L�`���$<'��"x��DDD�B��e	b"pD�0��4�NI�L:i҈(4�"<��Bl�$��0LǄ��:t�7�(��2�AA4�D�6$:<<x�Ӣ&	҄ �i�4�Oa�L0�Ν8a�H0AA�!�B�'���Q�{J3㏦n�@��+UK�n�[l4cQ�Ds�9l2c�$����*�!n��K.��:7V�ͧ������G�W��, �jHiQ��v��#>A�Μ���UR��n���N���*�E'Q�6��:�ԩ�n5O���vح�Owm�myO1�6?���e���D��m�8Һp1�ʋ"���\�M�2]q�eV�ۗga������[��s�r�X�##��VT�G]1^Wq�e��ל�-�]طzR�D�����'�n(S8�[gNn�ֲdީ�Az2:Im;5*����	I,��.�P~���cA���8���͛k-��5f�hU�4E�,h�&��/�����l�
���X����*p�u��t�ް1�IKn�lɋ4�F�YxA=6�∈�j@�QI�M(�Bhh������ �<\��{�~��_�G=;�x�J�3��Q;��f߱�Ϣ����[���/�fffg��UU�ҫww}3333>Ϣ����[����ffff}�EU_-*�wv��a0ن�,��L,�Oi�4��㤟�I�L,�<�r#[�N�5�j�[�]T��b�t&][R:\1���x�i�%�u	�u�C(����V��I�k�f��kt	]4H��g.�n�����0q[e!�ꥍ֫mu�\�Rc4�6��3�a��K�X�+,̸�æt!�M�����U��.oE�.�����0Y���I�m�R�3�c��ٺ�L^f�WjL���U)��و�T�ݦ٥�5�ل6`Ɩn̥�̭���V5�Lv-�6&���v#Z��t�%Ֆ�`1���M/9�	�f������ay�Dcwg[�u�F.�!�Z�3�:�m�h]�+�����Fk3�D�f�.��-]��ߐI�Ixj~_�;Dm����]����s��1{Q�jĩ���뫢���]p��ޓM��	S7I;�÷�[o�KS*�L�ѭ�J۸$Ҥ(�̼�{%.��I�1�eaEX�P����uyqo\Mq}�P��p$��[l�t"Σ�Qh�&b�
�ߏHthk��_%��
b^��3���8�s�{���z�ݬ]F�RQ�0��&�Ü/��GaB��hW�,
�����h8HP1{l�b�bT6�B�j�N����xp��!Z$.Qh��1'��C>^D�t��p��K(��i��4醚ag��ڋs����%4��5t)У �/�1�//<jj֟|�B)�lZ�˪�ãP�����jfH!�B%&�u 83[
5�"
#"�y�� �8R��U"�	KLC�WC��{p��lM���O�z�d��*\N�u[ײ�l �ʖn\1�4t��ή�C�QwU�������Y��9���y����Av���I�z��E�p��(�ĚQ�t�M<i�4�<xg��e��sd$���-�d(�ldx��666�����M��]5�;�}����q鳳��S���57n&�Ǎ4�p�2��-R��9|/�UEU=������ +��(�O)8�z��>Tp�Q�[_Io�u^_B+�nWPRS��M6l��gA�o�,��,����'��A�|�\D"V��$����`�Q,�'	:Q��L>4�t�L,��F�nURP�UT!���������B���h��(��08�+��/-%�h����/�A9hMDZ5�4�:*ʾT_�}�� B8��QJ��"���o#�ٍ6a&�kĒi�����ӳ����tQ���m�K|�gۛ�a�A�R��	65H�%C��4�OF�r�;���=��V�3�ğ|Qft�M<i�4|8`Ѡ�O��X��:YD�ʊBP7Et1��M6���C!�ET5�Yu��#,wFD�)�J��ժZGZ���35�]M�}o-l1���0�k2w��};̉���R)C7���L&5[��Ra䕻.ܺ~j�v�B�i;�D����[Z7�6�؂5w7m.�0J�e��nf�yװ�,�k��i(�
O�w��((;���D���Ǣb^"_Ͳs��)M)X�{�I���cztţȮzQ����2"G�R%|YGWFR�q�1Z1w'����Z�����}zƞ��(�-]�ed�)�q@p��x�w3����˙��m��R�$��$�ύ$�N�|x���4�i��<1��	PU�|��Xsɦ�wT _q����{̦�:Ng!�lǿ�������u���GxZ8�3�#�E�usNI�ˈa�!�i�;vXJ8B��GCo���C��z�o�jfE(��~cm�l�1L\�6�\]�r{�DF'�U����,��S�0ȹ���N��3��,~��z)I�H�J鋇�fD9q0yO��s*�}PΞ$�'J<|a��M<i�4�<xg��kI�dq �M���S�A�P1����q��Q���>�ͱ��7��=~'I�;�0t��+uQ�gI����J�a���K��ju��Z��}$��y�9���hӑ�(��ԟ6y���:
2+���p�z��h��B��a�6{6 b>���a��DDZ�{ŋ����ㄞ$��>4��4�i��<3�H��>��uȻ��1���mM5�"l(�j{h�e.�WC��>��6���w ��Hb�l^��F�O"��-E#�#�jHV������X�z��93����殐k]�Ȃd|��Ω��&sZ�.g��ǯ�~���T�A�K�T<�&G�^S���%<��"ɶ6T�R�(d.���*4��,���pD3�$g�$�'J4�M4�ƚa�M0�ǆx�GM�M�UU$"�@����.�4�p�!�N�H0��nU).%*��v�.��.�W;8��d`P}�~�-��|%�T?,���� �<Q�X,iH�P#�L���N�՝m��q�ά#OC�cH:�Evvƾ�ۥۻ�Ec�N�,A��E��r<H��<I5cu�Y���Wٓ&+Ѝ�ڊ=�ǓoA	�7v��!�⫀���/I~K=�d�IFEŝκ�u14x�g���:����7�8�PRh���?R$��#���F�0�m�����R��.�>�O�Utt[��8��:��\6�h��Z�KA�2�$�N�x�N�i�M0Ӧ�Y��<Y&�|�"11&6666�M}�((/�Q���8�0�Z'Ф��q��CDj����͋�	V!Q��K���ۯ�Ď�C��W��V��^8�3 ����i�*a9�#ćN�ϑ��W�x>������eãnκ��pa:�Ɍ�͉�
	DA&�8*�i�;�y�ĵ��(1A'���kC��E�x��,����"'DL�"%���	�&	�pN(A
AD��؆Ͳ%���'D�'�L!�`�&	�`�&��x�x��b%�"Y�"&	�"%M���'�pK�Å�x�����>>0N� �#�I��0O	�0�t��������L�AA4�Dw&�jD�"Y��<x���t�D�8"xD�O���:Y���>�AH||B]��'=}>�kĭ$}�]^�Ax�������7�����5kY�lQ��j�G�c,�x�U�meN(��:���r̤u���^Wb)�B�e�2�������yL����z��������SY�Ƭ�@��O�b'DsD�<�C1t��A�Ij+�t�G�uV����EL�"��a��Aд��FͥkZ��5�a&}���ٝ�1��(����f�P���-��~�����ʾ��i����>���ZUn���������UUq���ݿ����|���1U����3333�UU�*�wv�k!�0م�a�M4�ƚa�M0�ǆx�JW�6^�ӫ��n��9��*�w4��\�aH�:R:v%5!@D�Dj��2�ˣ:��/#��A��m�[q1���9<�^X��qK?�uE�ZQ5Ѷ,\_��g5Pw��^Pp�B�|V,Z��^^
'z�`��ș�%�F�<��<�,�
��#���n�*<�4Z��at�'�0���4�Oi��4����+۷3��S�kO4-y%��  ��!-�����P�N���3�������	�UN�<�m��y&��\1~S�I��Ce�3�]'��q��	8��}�*��x����_��q\8���ث��m��r��/.�m!�����r��M�Sc�����o�P�ה��G��Z�%������N�x��4�x�L4�x��I駰�M��bT )�����O{�J��-��߄>��`��#��ي�Y��T�&�W�;�2�cL�"4�6x .c5p?�WG���>4�v�U�ժ�S��}��gwu��.��f$PɻJ�:��:�µ�5��FR�紵]J����T�$s��Ӕ3k�9�P]T��T��UUr+�j�:9�a��~~G�XB�h�G|�co�J,]�]�+��x2L+���Δ�23��d�aǕ�t<���*G�R�c�"�t#�0]�f��R��/q-�N�	���m�Þ rQJ�5��G��0RDv`j��3M$�%�x���L4�i�L,��,�G�}iKR��P�hT�hL�=E��� $fh�<2�h����x���4ʪ!��Lcm��3�g���L;��t��~E*_��;܈N�و��{`����hIHu�S:�]
���@�D$Ca����*�WUt4w-��,�8���ů�_�"��JU��u��{0��s�D�Р���2�^Tt:P�0��K(���O�4�i�L,��,��E��"�Z���1�)f>� Z�퍳U�ןFlS]]:�x�#��X��-1���J��#�b��R��MvK+��k^$j�x���x2�q/cE�M�7H���<�^�H��娞��8��|{�LN�i�p��x�<w�eMf`�tLu�X�:H��4Pt��I�L(�4�Oi��4����"w���H69ɮ9mg5UQ��;�-񏉇�l[F��Ө�d��l|Z29����[��0��o���������"K8�1�8�����3���i��k��r��q�P�a�A���t�A*Ϲ��$s.bG�|G�ʇe��qp�u��p��nͨ8<��L�����Yl��qH�i'�4�Ӧ�Y��a����X�:I��h-TiD�ueQDC7hYG�,�+���K�Z"�JUR�QR9�OM��s$�˒�+d$V�x ���C�ߍPB���}h�!��ہ"w�-E���s���`y���Yl.������E����`�i�n��D�U�K	��9}�X0�^Vj�i*&!$��r���?{��"�*AS�S��C�����ui���k����������-yZ �x�)}ߣ�	�q.""\��($�aH��'O�����|qUɲ�}kzzy�NLL� ��i���h��ǃi���A����CDQGB��i�N�Tqp�8�c�c�����=82�Y&�||i��0�L4�ƞ,e�$r̉�2Kr9j��o� mT7�Yn��ٴ.�����-f}�ػ�[~Z��\���d��.j&|1���H]��gF:4B��Q y�B��-�63��ky�xm��P�Wd#��Q�kR�]m]lP�3�9��1ua��<Zß�XL��"N�0�Y+��
��K�|��jP�l<�������Z-�|��L�.)0$��p��:X�|t��'�|Q��!��ΐ��LYݦ�-�-����Bi4��U��DR��� Qv�,�!�K;w�6�[V��ϝ/E\�	H�2���0�#�kZQ�j:��o��"������"�1����y�o�}�l>�U����l��ᐰ�� �թ������kB�M;��-+��*ۥ�);�(��'�?7O"����!B�'���(Q#���Q�K$�E�|t��xi��x�ǆY�F�&v�\MDӞD3�n�m�0���t�p��`������h�2ϩ�Q�ˈT�*;_I�.g��\^Z�f�5<���qq>X�Q^]Zl)Ջ�����o�D�j1B:b ��+���ӅI�Y;c��E�]8����s�GN���? ���P�W�QE%P0�����g����H���$ƿ��"I�������I�����La�N� I"b�@���
i�bH�f �&"	��p&���	�Ba�f��&	��&	�bb`�B`�f	�&	!�$����$�H�$����$�"H��D�DIĐI LDL���LDI�DDđ$B�DLDI�$,1$DIDL,D�D�ID�0�D$ PL3L2�D�$A��KDD�	$@D�ID���D�$ADDD��D�I�DB�D$DKDB�KD�$I$DDLDDI��ID�,DLA$ADD�,DK��KDD�,I�)�DD�,D,$DK�D�,D,�$AD,DK$AIDD���D�,DK��DK�D�,BB�DK�D�,D,�IDD��I1K�B�DI�L��1LDLAD�0�D�ID�0�D�DĐ��1I IDD�,D�D$DLK�0�D�1I�A10DL,D�111��`0ID�ID��A$DLDA0��1LD1IA$A LDLADA$K1LDLDB�LD��0�L!$0�$�$LA$�Hd�HHd�Hd��  � � ��!�	!	�!	!�	!� �"	!�	!	"X$�HBH$�Hf�	!��``````dB@�� aBE�� eP�� aHBE�� a�1��<�`H�� eHR��:6h0�DD�,�N4#��2$�@�0�@Ȱ0$�L@ aB����`e�� `��`dQ a ` eQ eS�P&�HP��``  aXVE�� d�0RA��``A��`eE��5�jҌ)��#*�ʐ0��:aqB��*@Ȱ0��(�Ȱ2��@��)
@���@�$�@�$�@�&
��(��(��
�# 0) ʰ) �H���B0	 �� Y��1 �@B0��@B0, @J�B�0�� C"CC �"C#�)
J0��C"CC+��0$2$)+�,2�Ȑ��"C(C B��0�2�2�Ȑ��
CCCB�$2�2���
C#	�00���`�1����I��
D1��2C��B���C�C$1��C$2C�C�0B�X��8!q!�e�!�e�!�!��b!�d�d�d�!HHba�ba�d�f�!�e�!�d�!�e�"ba�e�!��!��a�d�d�d�!��!�e�!��Xb�$�!�a�e�!��XR!��Ha�Xb!�!H!�!�!�a�!�CR�
A��2��1��)�C0�2C�pNC,2C$2CA$0�L�D	$�DA0A�KIIA0DA0D	0DA0D�IDA0II@�A�AAL	AIA0A���)@L��A040D	0D�PI��L�AA$�D�A�A$@�L�@�D�DA�@A�$�DALL0DA0!��@�A0A$00�,�0�$�2@I �@I$�,�@DA0L	$�2A�`�2@�0��L@�@I$��:���H d�H	 a��
�`$���`f�	�`&`Y����`f`�`f
	�� �`&`Y��"�H"d!\`�&`f����`I� &	�`f���	�& ��a��&�&	�"Hf ��&a	����`� ��&�_R��N�L`|c־�:���yLS��>�?&U �Q�TVaM���ԗ������'}}���_z|�����h���/�6���o?�?����6D���������80p�``��y��L�����SoG�a�Y���9���óG�`��o�����;�`}������ ?���w� �������C�"���Ch���@��*X�O�#��?��}��!�`c��0S��hO��!��������~A�~�S��P ;�/������@r&�t���9�����`ߡ���^4��'`������ C?y��C�����Mo��~��q��D��oo�:>��18z0e@@s#-(�b��"��A� �9���	@��U�aPH �*,J*A"��C�Q�A���`��t?-�D�)
����@}����������#��	@=�� �P"��@L
��  �a��!@D�@�6�����?X��>	�v�A����R	�]�ڇ����c�0����O���7����������@'�;4'���q�������/�?X��O����	���}�3���_���@�#�����?�C�a���~�x}a�Z��P��_�t�/�J������B���K�L�����:�������t#��ټQ @ ���P ?W��?�T��������֔���=>��:�v���݆���`D?��b

;v�}���cO������@P��H~�@��H� �<����`a����0d��b�r���|huÏ��x4�?�x�v�Bv�\�>	�G�P�>��?�����>�����*���f�?� �O��_h��Ǎ��?�y����@}��C�I���O����O��~����>����)
��O�C�����G����xz�@���_���?o��J?�@T ������g�����`~����~���q����h������G��9��`Cq\	��A�.��@k�!�H~��~ϩ<�d��Y��u�E
N�No�EĀ���9}�Xӗ�#$��~�~���@�^����p}���^ô��b��86��~��ȼ�������!I��+������������o�����?�<EG��N��?W���?G<��~A���������1����:XW��!��߷��w$S�	
�gp