BZh91AY&SY_�uV_�py����������`ڞ[�
� =�  R����D n�  4  
�     P �j��� �  P  	}�  ,�6�Q�B�1�(m��U3}I�w����#�I�L�R��;aZ�R�`�km��m�F�n�<�  >�;�L�mM�l��̀�2[��[F�co�/1�5�T�e�6��8j�5��Kf�H>�|�  ]�
�J}�Z�����ʕf0-Z�͏�S�Ƃ7����4m�����ٕlʶ��Mo#� >��`}j�,U��fHKZ�A��6n����v�55�w̍Vl3&Zm6�kOH8 �v�jֶ33im�V���M6�V�Q��@#f��mf��0����݅  @ �   @` )                j����U*�F�����C��J����M4d��h�`�&��&�1��Q�ꪪb` �0 � 	�# I�A7�*�        D�	�D���4'�0�d�hz�4zd��DJ�F��L M2=^�d(��$����I�(}��i��o��@@K^��P�( �z�D=��� )��J�����/���������)���C�!	$"*��mo�%-U�'��`UU�����׼���6倁�j�	y�����n	��w����__�=���f��k?��Z��ׯ��(�.=>�)�E���+�H��zA���RU���7]/��Ձ/�;�B�.C�fA߳�ኸ���&yw����zzQ[+��oH�R�Y{��嚜�}�o����,�ܪ�<�\R��>մ�V�o����n-�
�b��[bg���T��mZ�i��DаBq���}4�-�){KЖ��(�l�����m��G��Qm�(�Ojq:���z`��	*o(�.��Qh����T4�'w�hV�]7��S�S���E�����Y8{�B����j<��Z���h�7ąȹ�rTH�߻�=�;gl�&����h�� n,�\'r)����W(�A*�`�&ŗ�2B��!E�㏅���0ڝ�D�O+<���}V�ju�
�V�ݗ��%��ك!��Ƹ-��e�RV�*ʐ�%z�Nb8���&�ɀ\�[tuř��'0j�U� @�)�B�\�'�$	�����F�PT�x����J��y[�p��3M(��]����Y�	A����G���(+�Tў9pr�wC0okR�� hp x4,�]mB�T��[國9��=t�A�{�h<QXQg�E@&��;l�0�^�^�\�_O�a����D�6�Y�1kG�ЛZ�Z�Z4�ySI�a�$=-}�F%z��h�6�ON�H+���ȏ�j�،��Փ�7��0
Ҍ��oGQ	�{��	��`����߶�3��'қ<�����w;�.h�
�E7�#*q:Q"wV'/���f�<��2�*�5J��/B�U:B����7�
����z�]۪s5Qs��Nh�Т}<$�jW������%mȹ�}��^�(����&qf:7��5&r/{����U��A,����M�/�d��<}tS�t��l���l���'�yV{��1���P��\*�ݗü��Yك!�Ƹ/H�\;+J�⥕ �<��1N�I��I�x��_���9�VJ§B8�t�W9������@����	ASI�AN����0�=0f�7��(�a��ٸK6! ��`]�A(*iS�!˃��o�}��ó�dѐ�&��k�7<��=Yȳ�Y���C6�=�4
Ҋ���M9<2�T�a탘f�\��<����=_W8��,���V�+�J�J�J
�hg,x�"3I���!���Vp�'b>L��6u}8� H���I��H��v#:zud����7��.��gG
x�J�O{����/3�˾��g�d8@�����_�naݹ��a�ᕞV�pʙ�ܱ�F�6?O�|�����(p��cC��
�7gĭ��FW�,����,��U����U�0~�B�P�U0�L���e��<Z<Y{��K<���-z6�SJ&�t�f��j:�`�**﷫WѺe�%��}sW+�J����VV�TI^��T�Բ��v��y�n��y�Z7R�%rƧ�>�U��P�+�!����kݠ���خ�ezbɃu+�Jl*U�Ї�*>X���
�B���-3�4�ڐ��d�F�)�J��lZ4��6,nЪ�x␣Z�))CG�߲bK�����d��^�ȭ2׆ό����֤�YD�.�����G�(�s�hV֥���t�-��(�54��8eK=��-�Y<�<2��ޣu/�.ǵX��̢��T�}(V��x")xmR>�|+D<D1V����wrũt���c��+�
��Z`��\�b2�"ߠ��b���[yf1�pL�a�(���
~��N�į�*}�}���5�|q��7�`�ԷS��M��&*�DϬmX��ɦ��1j�
�F��O>�m��oǓ�D�ء�6���m@��F���M�%b�cn�)���D�T��E���Nn ���+)�R�R�^�z�}�Z�Y�[�[#�<ޯ[�DV[�Y��b���YЫ�WN����q���}
+�m5�J�u�u>��JȮ�eph��������,Z�A;�ʏ�0~�B�P�|���-3�ɣ+�-��Va�8����1��F��3�У_����凛�%�S�T��I��5R�����>m��	��T�/*n~��W�&}cj�ŋ��"���b��֞}��%?(<ߏ'���Cmߵ2Z~�%��&)���:FSfJp�b1�/h�
�9U)��G�	1!k�y�|!:��
��W�{�}�OR��$)bb�	�(LR-U���B�B�P�R��W�1h��R�&��b�6Н�Bh������ܓ�p��4]_���:�O��7Lʉ����)x>��c�YJ���
�̰�4v�/���d~�����<$��A��D��g���x�9É&ص��ΦFΓ��U<�K�5��^��|����J��U����lS�As���v�u�n�Y�"�m�w�����MZ?h�b�8{��ӽ���k�8���ѷG��~���ë>Gݣ���.��ӏ�:?C��9����B��#�A�3��t�ƨ�����e���7H���f��������{/���z�>���h����o�Gα���0�b7�q�{�>G�=��gۏDt���F�8�R��o�}Iœ��pG�r�+����5�x��1'Ȯ��K�M�X��Ӎ��}��UV89�t|E�V?�/zN�|#�qi�B�5���ߩ#D�sۛ��E���r��n)�h��/��Jl�LE#c�\�}̼:,�i�#�<�9�;�6��ҽ;��7���rr�)�o�9�%���>Q&)�u�y��#eWu!����Ǣ|�l��_��:��.<X#�"6=f��#Ք܋���O�u���8��4�9���[�#c9�IJ��ƶ���7�֪�Vb�G޵��7Y��5s':��xe^�MT����=�����i�9�o��i���/���}Ü�/#_#����G/E��d�o��M��^��?���Vr�"���D�>yru����Mߎ�(�XiZ����+��t5�,^�]�b��t�{����2���9y(�-�K�����|S���yTO������Q�gЧ�9�;d9����(��7:�<s��7=o
N��U�����p�Í-��ݰ�WR8I�Ӈ<��7[�N�4�u_rtӃ������қ1��4|s�T��sݺw=ˈ�~��Th�k�<�i��>��p�{���!j�}��DD$˞��J"��NR���if���(���\�Ԋ|��ߣ	�hs��8I�^@B�?w�8O�d�>i}���s�ћ\�M^F�9�
}�3��/o�p���̘�D_C�d�;Ƕ��R�(�x�l��/iNs_A��6Ti�|��>Qo�Ͼ�{�t���N�T�e�
\�^y���/U�o)Z�VR��p�Ĺ��j�l6,s�_C�Kr�jT�<�M6!z�$Lf�<��	�]8s�zw�=�w�bmqog��ݖn��g~�^d�g�L�!�������e��l�pځ�}W���ř}*�_�|֞�`�y���O���!ƾ���5"_�3]��bsאJ�3��.q\�\���i$�G�1הG~؈-N�:S�\���u��%�5�Cwې������A�1�y'�<�,5}JH�G��1����w�3�82�i�����%��ٳe���mu�&��>���ș�~RJ�WW�9��p}]�_.x����d;�2Գs���	+����{�}��w/�?�x������'��ݟ��蹧3Y��p�R�	xi��M�gM��oY*�s�ܫۯ�Ú�.��Y���A��/��)8����4�x�(hx�"��8F�p��h�xG�
p��!þE��/�]Fx��e
p�CJ>�˦��:�υ3J|S�8R��F3s��ִ�0@�@gN�Q�����4]@�BΌA"�^����1'�Kȷ���bçO(�#�� %N-=�~Z�y��!���)��C�H��5q��tP�hQcd�v.���%oe4��!H2(0e��V���GAA��Q���N鴿st��!e4F1(��x_��VvF!�3J0Gi��8L�ͣ��?Oч�HA�4�!F!�65��p�8pУ�Q�FR�xn�)������#�)��V)��J�7s�})��!f�
���p*��uu�c�xӆ�&w��M��5�^��b4f��:�17mݚA�c!D�V�A��Cᔡ��c�o�Dq��C:i8>���X�R�(�E�Į�9��C8p�(�C��7�O�I�#D@�_iyG�T㤐CB8�������7V-z�#�/���{��+��b��hN��
��Fڹ�c�N[��R�\뗄,+���f�r�<}�>C�f�5'Q9G�;5��+�����:L�����Rk}�w�����WG��;��w����-�dP-k���?3�?{�"l�"�g[��`�S���GYɢ�Zi�������=���fw��T.sb뷆g5E��ӟ{��kϾe^4�v����Z9��|q�Ep���qk{̾y-�ov�*�Ǜ6�7X�8�k�q��kdU�I=��I]+�����?�����^�t��^�)q��ҟ�߲{��2�v���̝��B�e^���j��4�=�c=������P�K}��7̨��KX�{�{��V��;�r^���MO�Q�s8y+ޝ��y�y~��۶�wb����w���;�Z���U^L\�u���b�[m�ȏ�ֻ����N����s�n�<�N�����I�cNo-��<��I�$M)�sw��.�����*���1F!��^��W1�����'.q���\�rY�VX���jB|^m˞�(�Z��ێ{�C_��BU��N��Փ�.���/�;3����j��|�k�`�g���JqE���O^sxj���z���������>o$�E�Hﻼ3�w�̙��E��d�o�j��Ҝ��̙�cz���-������ms�YÔ��t�^Ӝ��Gw���w��Tw����Q��C�;˵���|�z�vO{�r��]:z-5����!9ͻ{�.���=�t2�ۚ.�׭\֯n����\��v�z���U���Sv��S7��tFb6��5kr�ާ;>��Zm��#�/M_�yqn`�ɫ��W����dBsz��͆�w�ν�Ω��>�s���Y���������6��q٪6�}��;���cq��1����3{�X��؜�>��퐿�dwf3�(��_��V��[l�[l�*��9[Ԕ#�-e[�vp����4���$j�g��ă~d��Ơ�$�8�ݛ�Q��\�Q7�P��������U�3�����r��nF�P��K�˔T�FImn*%����&��m>�պ9ɱk��U5���qHJ�SGW�����F��������B�#q)#�H���`��$����-z{�T����j��O�v��N��o1q&9E!�'RnR�ⰭG-�K�49��FcXޓL�hNc��G<}�躙��[ߴ���Y"�T8����["QH�U��+wv-M����Y;����m�����L��V���I1"��}!�w{����N���8�_R�lu���IG[��G��6H������黿,�O{�D���}ޞӛüw��������b���J*�Ү�i6A�D+j�j3�����k�����s�2_x�>���FDw����5�er6�r7QZ���'��]}/
s�uw�4�;V�q+�*�ي�s����:���:�(��o���ġ����/�Hq�5�	�-��� ڎ��<�7$��"-�"5l"M�m\j����5�HZF��3z�o ��|�>p"��q[J^��;��y4��2(�M	���D�$H��UL���X�W|�q�!�s�vH�#���ɍ��BM4�����:,�P��9���M�E�tO�%I>C���gy�ɳݝ�i�GXৗy���Ԛn֝�+�������60���[�����I&T5d�wﻗ9ĜoKà��7Ⱦc��C���7�J�:�t�Wj ��#��ai�mj״�Lٹy�Յgisw�Ϻs����ٻ��������FD�Dl�rZ_v�k9��X�c�P=����^�T m�V�</܂��kp�~>>������������|(�Q�>���~o���9�r�� X P� H   P���J � �x ,�`   @ `@ P��wwv�	 
 ����H��(� �4G1/���V`   4`  X �<  �UR��$ (@	 ( ��� 0  р `@ ln���  X
���/����/���_/���U0     р 0   UU@`@   `@ � �<� �L D    �{���0 F������~(����w`@  D      0T��   р 0 F � @� 0@    ջ���  �����'wwa  x , � h0  � &\̀         h� �<	 (  � �ݍ����A��ﾖ�K���K_|���� �� 
 �@
 � X��� 0�g� X   `0  �  4`�(@	 (�n����P�����D��}^����EUH����/���uJ}� {�>���!!!,BP�)B$!b��G�+������������^�-MB�!R�,P�-Bŋ�4$%I	M^B�*B�*V��Z�
�/)B���T�P�K�R/!y
BBBBX�
կ+B�k!R���4$*M		MR�>|��!��]O����CxҖu�ƭ���M��٣ȳKjcv4�k$bY A!�Bg�(��6����sxP�t�#M��S�sn��×� �Sj���. �$���H,Z>(3\%c��yGX��5��j��MʂZ��,'�5��i�-�%(!h�l"��!Rs$�&��Ph�ct��iHA+i���%� �Ŕnd��c&0�UX�Ru�#P�CJ,�H]?6�U�<cD/P�9��eD�n�
0b�4��� R�p��2H���<D1(�"c
2�S-��2���t���E�%4�z<��A2J��y";\5KIJ�B�,^������T\Qʤq8�E��K�2^슽�H[h��ԉB��\�ڪHj1X52"��}��-|g8S����=�(�����m�'sK1U���ɵ*�V���
"A��(��Բ��R�%H�F�)m�!ىب�PV䐊dL��jZ���l�el�׉T�Y9��|:�Sj��V�*TX�QC�n��jRfa�>o�_�wo��~w8���9�u�]o�{̹ȒH/9�s}UU<�zw�$����ꪩ��DG}��$�wwuUUW.�#���/�ϻ������q��#$aÌ0�U�r�f[��~BH_�Dr���DZ�B!IJR�E�CC���%ơQ)F�!2%y���a���6�`����X�x2���*�*��lID�|r%�!q�m���[2ޏ`�\ʜ%����ZkK#���l5cF�1�pdQ9$�$8�=H$��g���=�nY��:��u���o*˩�S��8�?�P�w< 8�}3�Y��9X�cCp��e��C�W�,(pX*��ǈ��Kb?��˞2`}���a��F�����q�6ߨ�f�:u&MG	Ƞg�2�Ό�����R|u�Y3.1�j�����J47��\��Y��GDt��4<e:����&.��aN3?g�i�=O�2$&Li��<�e:;a�;UW��c�Ճ�$;���e��ˆ|U��r��e�KX�eM�w3�����s�Ko��x�2�A��BO9�7�n!� ��'D�LόС�CK��_�� �B	�t�B�hi���=��o8��<Nl�H��3w���g�0Ǫ�ۦ��:kN*���J��@`��:g*��fg��	H��ȥ��	h��i����n�OS�挞%>Ob�ֵz�%Ɍ��:�ٻKn���,��3g;�l��K:=d�h�t�_O}���w�e�����L0�J!8A�f��_:<I#��ZS�����*H�b$;A���QP��n�B4E&Bc��W�vD+�T��IO�B.�v��!����;M��C��!+i]�K��LC$�i����it����nt����y:2,j_�̄��m��>�Ądd$#�����̹��'\|Zϗc��ᆋ�C��81���B�	�$���ӟ���W��)jםYu&��a�*�n4�1�_/�Y��Y��@//G,�0��h�n�p6�˔J�dht��8�V$�66t&�q�l��QR�#����x��x8c3�+�$~{�����Gi�I����1���L�mZZf���28��ٶc�Um�Lc&���'��=�m{�Z��x4�'�����L�����F!4�m�9�3��P�t�j��vM�zOOM�ew'��&2h�}����3�F��!ko�-}Ɯ�|�I���$؛�3��'�,�4CoqZ�bg�������K�C4Lf}�P�h�L�nI$�%y8'�<4;<�n�ǉ��>;N�����o
���!_���5���3T�y�xFU"˛�!\�mӻ$��`LLC�!d��œ!r��
+���x�ܼ$��(�bN�+m86��K!'��G��g�q�N�ޢ��R���g��#�#��l��"M\r����dL"�����Ǧ۳������'S����z��qy�k���q���"jA����eY�%3��|���)���x��Sv�-�^�!B/>�� Њ<�dE�|{�x�ב�;̗���,��a�z>�:!Mｔ��3�g��k_s�,��ڃ���jg��lC챧P*�C��[�0��+#M���]��Ý�2�̖�n���EI!=��گ�j��_����*��{Ȝ�\��Ԝ��O.�W#���\x�1�/��q_/�v�������97'S�w��.��9$�.��S��u�q�/KŜxϕ��x�q����^/c3�W⴪�Z�Wrk�����J9
3��,��7��7��r�؈�T�Ӿn9<B���rb|��s���r{���v���ۙv�f/ū¸^.wnv�:x�=����;^wn6�]�ƙ���j�����~^�`�I�`�]'I�"6�9����ww��2��>k�F��t��</-]q��w���}ǵ�x}]Xs�8�K�r�w��:p���6c4�߾!����.�o����Z���]G�?�3�yN,����2��0����Rϟ�S������f���=���%���~�ER�M/�Y��P�-䬟}�;�����˪��]���'����wU\��";���]�wu\��";����Yww|��C����]ϡ�>���˻�����ir\�-4��xWi��iӯfZ�Z�jѴ�W�R��nl��%���v�G
�K'�2KG�o4KOR���'��4�|bq=1y��ؠn�n�Ն�����oHH/sڨ�6Թ���$(��n��q�=(1*r�Kҭ�&Y<���t0
���F�!���{�	��L���hV�4�i2��(�ŠgZ����Ju?[��Uվ�i��w/:u����>�ͻwٕjիV��*bYʝI��4�>,���Ĥ������ ,��_�~D,,�8�L�&�:�CA��Ћk�vF)��W�Ia�2��!����1'*eG��R�Y��I���IC`&��X��8]0\n������I(,�4�`堤�F��:�CP���;J}<�'���Y�Y#rQ�Q�0YS���0��]x�!Bs��� �׹�'�Iqٍ��A�!�<����T!�\sSDM���	A
A�Bo$��������7nE-ԛ�mD)&EY��i��"T�(8�ɵ�^���P�����kL�q�B��&�A�kh��3=��ũTy:0�B��p�|�}<qJəl�m̳D<�^�&b������D��X@�iKD|��<h��ʒ�Dd˪�r5:�(���<�ԩ�Q�޸})��sL܌K�s0�"�%G����%��x��e�=�g�겫H�u٠�50~j���R{Rm8a�t��.,k�Z��Q�U���b@�	{Lf@�2��ԝT~J�T��փ��X��Rä�dh�v�i��_�!C�>��[�p�����[�I�KSR��vU|�:�3l8T�'��x\J��?&!�F�)i�����N�aFu���)6�]ظ��[ׄ�.����zKk��&�zQ���k�c�v�5+[n�T��rH����.6f��'�&#�<*4�:9]�N�����}�I����a�w?]��шy�Ã���-��DA��<��B�9��WO謃.���㺵jիF�L�^w5#t�*k�ú�)ra4Q�T�ҝJ�JeN���M2'�>����2Q�S�S�ěRm*g����!��\�Q�%"bi-]�6�V[jtOS��p���e�c8 �YM�`,���hh�>�&����2����c1#^�B6ذ�3A��Z��,�u�،L0�:��fI�RtS�d��]���Y˧Fݫ�3A���B��_�  ���n �[Bi��Mӓ�Jy	�&����׺|z��fg�-�'���e�S�~��~Ri
!��T��E2�!���X��!̅Ɋ���c���Y�NKV���;���)���1��<LJ�`�ً�ݵ��[���Χ�c�LN���GGO*;=a��J}1<:0��a�4�lӧ!C��:5^xD�q�!ʱ�.���<S�K�yi�����h����L��Mr����e�!����S#\�\�qC��B$�:���W/���[���O<���-���h6���d����mq�J^����м��q��r�:O����\�9�`5f�.;��fE�G
m㝐�q���E��(�6Ї`2L*,Et�L��mk-�e%l¡
��J��I�헊ht6�j����цݫ
�Lc�O�4�D!�-|V�� Ԙ�ȱ�<�;t�LN� Xz�B>31�=O��?Z��}>�-�m>5>��i����e[�)r�����;v�����l+\�LN��� ��BC�rY
�)V�A�Ǧt·���0Ў��� ��hv@(� �=�|s�rnM'�GN+
�Lc�O��4_���?c!
��˜ݯ+&�3���V�ɐ5C��'6�-�)�<��Ӿ���x�i�>L�=\�x�d���B ���Q��3������^���:J?}O=�4|tu��fL��=Զ\�C����5��4�L��qXV�c4���cIVvT����PTŊa ���j�f�[��x�I$�$�Ⱦt�2d:8v��KPjO%f�!E��A%$�M(؈�y	�6�R�k����3�.1������ك�+�Nt�ə����ܸ?��fi��3h�>2��<�]�x9�bB`4:3��������֋E���j�:�����N̝�6����Kӣ�u=�MȞ"x�_�f,�L�~Z��W���'�����^+���q�8��Y��{WK���ӌ��\Z�Z�7%�Ļ�����Ԝ���强g���������+���q]>g՝�c�W��j���g�ӌo�s8�^���ܼg�8���B�-��R�N�8���B���>��O���E�Qi�'
S���m��/�¸���k�l�̹��gkΗ6�4�f/ū��^1�^/�����l��4����\��sM8��s�\Tk�45�=F����G�Ţ�ԥ���7�9ۼ4��T�Q	�W�NB�Fmw��5j�i�I��>[��3���XA�f�h��Q�s������:]����7ɾ�M76��Jm.��g�YJ��\g���|ᮋW7&��=m`ź�n��n�l�Nij*��l�t���6�2{t�
�w�)�4�)d�2�D��j!��*F@(���4r<��n�Qf�!JA�!`!�)�]����wD7k&`X-"�RX����4\�������Nj@�LжEDv��OZ�!J��#c�\��zF*���W�׈��V�+!_�~7���{�ȸ���~�p��C��B��Q����_x3��K��S��ϣ3}s;W��BV亢ǲ������x�_���A#j�r7�J��Q�F�kC�Z�u<q�)�1}����mmA�[<�9�Ƹ=��e����Z�ݍ;r� �I�A~8��'�� $!��e{(�F�q��œxY��d+��6T�SE������o#�G���(�J�E�NSƕ�E�?٩~�M/��e���.�}O�������w>�'���Yww|��Cwwue����o��������s|�����U�w|���S�+
�Lc��q�cM{��5y�D0���Q&'l����ܭ�<�m��JQA��+R�!b�H1h��j�I�Y.�2���8�񳊉���vl4Yj�E|�u�$�&T�4%�pZq�Q3�?�)�AI =��Y`ֽ#lX�kH�T�OW�Yx;4�8�:�ߓF&�om���,ȩ�z쭀¸Cw|�!04��29�F��-��6�q4��'C�����0����~O�-[��zxS��P?o��eY���Z4(�:A��Qʦ7�UUE"Qb��w�߇:�%N$x8�ܚOħ��+
�Lc��?1�i�>�i���k�վ��?8~7��\x��ߖZ��Wg==L�ߦf�w��:vB��� i.y�h�p{�t��N6E�"�e�a�z8�&2˄PuM��1���(�I4%�ɥ���3��y5���MLJ_׎p��{�X�g3t�1���IV-Ko�e�§]?�K<1�aZi�p���4ԥ��eHTAdJ�mQkT�&C��q��Cg��&#cq9&��L]G3�&��qF�����}U�e�Kj�ۊ��z�*^��Fk���ƕ�r��*-#+H�ز3M�5M����:&�CzF9QB�q��j�C�ް�4.��x;^��3���~<;�\�}�"g͸�cI���8i:ON͘l��&�2ݣa�]���S������|�颛x�+M1�J��QE��yyE�1{T�n_2�SC��*׾���_���'�]N���|��>0W*!+$N,��hci�w��Ƈ���͹�{}�'�i�R�+��_63�ֵ����=��<�
�<d�L�t�z����KJ��[!1��x�\U��kx ��i�ô˾G� ���6�+�j�<q�cN����L�ؐ,@�2"l��"Y�?#jb��>�5 Z�b,XŐH�&:F" yB��+$�6�f5�cD���5�b�!clHq�;H9���z��i���F\Y�S�����j����D�Rd�r!\�";H�m��'���߸ĭ�T�J��dĿ���g�=L/N;L�W%�1��UZ0=tde�� ��X%�c!�4@���b��^I�~�L�����O;U�ںM�'�wJ7�x�2�L�K����Ϊ8� ���X�d�]
���c��!$#������%���v�R���xV�'�:ק��+
�i�N*�i������Ԝ?���Z�Og�Yȗ1XS�B������0��[t6ϏGLMͧ����_v�<�)�`�}^ʝ�s�i�特;4�ђ���$�����S����5��^��V��]�ե��\M�����ǭ������M����Ř<ϒ�'�:���c'�1�M��U�Ooh�f�V���V��_��M(,�0��i���o��@x�G��vt�ԋ����~��>�Kz��g���h�t��]3n(|	�y�g |����և��I�G{�3:@t��i��O���|Mlu�U�����X)
nij�L76���]m?&�q�ժ�-�O��ޓ��ٿ�&�I	��Z@^
��C��G�?���HD�?G.��a��O4�(�u=7�n|k�J9?y?k4����1��\��1懌x�
4�2<t̅��uC�ަ���J�=�I�.�E�Z���o���M��i5�X�����5����<�V�X��~q��w��~O�'ɉ��ӵaX�?�\)���8rcY�J��D1�U�D�l9N��?�C����]:R�4�c�ɏ��a�h�*����+]W[lZ���H�PSD�m���I�m%�z�q/Yz1�^I���&$��'i1<y1#�8g��.�k(�Ω˨��/���:�l�^>]��G�!j�"w�|�O�Tꞧ�g�bm���^��/&���{N�O�|��:)F?O�YY�~���y�S�QȆL'U�!���(,^�<ᓣ��ѯr[^�1�vh�aX�8V�U|�:��Je.�Y�X�*��ɖj���X�z��·b|qƩ*I*����a�'];AN�g�:O��4�i3I>N�i�ɡ�a4����n|���-��T�QbE���:gs Vc��Pƿ��2UB;X�lϿ�=<pp�,� � m,6��:8��>6�t�]-V�Wj��ɹ�'$���;�]I�<B�b��U���ڿ.�����/q�8�+����~WJ�Zs-��^w\��ND�ܗ��%�K����ˋ�W8�qg�l�/��+��z����q_/��{V��j�'�.Q9�ܗ'�ˮ^�-G'�r�|���Qɉ�!R�d;Q����z����\��@�-Q������v�6�.���:i�/
�x^+�����;y���gk���3J��^�p�/f8�+��������˽�O�%{�m;YZӈ�(�5I���ܫT��̅��d<W�-WT�{qh�r/�J�{zo;�"��me�Ӿn輵<�i5r">���yj&���M伫E/"H�[Q�x��o��I�W~wUe�����o����ꬻ����-}���Yww˹�Z�������s|��wwUV]�.��c����]��Ě\�6��j�8��n��Vf\̽����m�Ӥ��>M�S�޳<U��T�`�kӤ�N�'�M�'�gϻ��٠}��(F�\x�-P:Ǆ��rto
�J<���a��8���txP�2�Yˈ�^��� zu�O>'��|�+��HtB:RoM���V���a�9�ms���6��OӾ�C���2��l��+��+I�Є!<;�����z:����MN��=4�����:��V�q�[I��nh�v5EJ������,�,�I�tkUKe��h=���;���<t�+�jӍ1�͹��55A3���4��i�O;{Ӓi �ì��
Q(J�C&��H)�ѢP�FR�Y;$\�x�d��%�pԤq��!�oY�<C�����0�E�l�4ǲd�[Zۉ�U�|gLFw������§KJ�/Gb��p��IU*y_ņ����~��	�I�z�q*_zN����^��δ�>:0plw'��z=84>N��� g922!J���l�#5?'N~��6rz��G��ٍ?6!��Q�3���:4��߆��M��O�sO���;�<=��N'�,��60�:�������a��wd���`�0q�����+1d �	r�*�ETJo���[]�Z��|���ğNT�9�O���É��C�<��Y.e�M��v�0��+
�tڴ��SR����
@���P?+�Ec?6�C�f��c���MqzM'N���m.�L�U��5XZˋ,4�S�b�ٳ���<O��m`8ݘ!OeZ���J��"�%d1��V��d$
�l��q�t��0�i�`,���a�STQ*�,�[s�TBB`*ν��cw PS�!��R�1���v*�2	ѵÁpu��pɍy������w����J*B�%�K7t�]v�q9SC�d;)���'���I�9ǳ3Yrt�����r�>�������N��w�m��ʫj�N�~>4��;�i+G��&ӣi�[�SE4ڰ�W��<1���H���	���p�p�p����Q��i�����F̊B]6]/ �SKR�9�YDmw(��}�蹽��lH�1"&$��1�����u��H'M{����h�YZ�\mR���D�E�\m�6>>20��dq�	`�P������V*�94�����U*��t�s�
�wwڭ��&LOzs~xW-۹������s:g�u{4Θ����LcchC<���q��4����fͶ�+������
U%
���Fp���CWX$���:Ko�����77:t�mhxT�{�R)��R�m��Ԯ�������yT�hhI �%�=��$�bt0�%N�X�8���xhy>�Y+�I�vm;�=;4t�X!���1�M9��HiZER�cĩ2	�]��R<8Հ�-�٤��ڻO�|t1;0׆��NҟO/^�N�1'�rd�ƊJ��(��R��A�nAxp���c]Ϧt�)��/R�Yk,ؿ�{4m546<��d�gg��y4};N�)�t���zV��?+
�~1�1��^3-e�761�$'A8�Q����Gdb713g��'����ҭ�<j�}��F�DYF"�bmV�,D�UR�i��k����n�p읧gR��j��j�6������H��y��~t�����h��5[�;N��i�E�=�VΆ��߾'�����]�^�U⪺Z�V��W��j��ʳ�LÝ	�.tn]]z˓�r�u�z���S�Y1�_�������2ޗ�j�'1�u�'"rnK�w�%��K��$��r���/9�x������r��q�^1�s-�q̷㫮D�Ñ.���.O+�\�!�;P�>X������V�j�n���-Q�B���(��|��	���;���v�6�]+��1xv���z�[c���<{���gk����y�q��j�
�x^8�z�/�~��,[�q��\����$�ˉ��iŧ?(u�Ӭo��ڈ�=��Du*���G�e�wg>9�����w���u��d/мd�&1dST�s��u�G�WQ��f>�B�#ygje�v�:��3Ij/q!aHQ�MM�)������J\~��i���h��G�&�q��]Z����A'G
Rא���ψUF�^�-llQ��2T|v�]�O8h��˧�v�B��hɷ�xx�Dr�b2�1Z� A���4�|�Ռd��"6M��\�8�F�Cd��5��"3	�G�b:q��b�243r�/Y�#��S�H!')d>���}mw����3^�FS��4*oy�Y,[�ÂZכ���HA�J�O(�j���o���x��Ț'��f�=�y��W�{\ˬ6��mz�i:�7~�F#��'������95Z��ڻ#.��q4���#.��//<N]�{y���o�k�+k�oCkCDv��rD�+�"X��*�1:��#V��,V�A�ȭq�*ti��4k��V�Lv��p����#$8*�iҷbX�٪�$B�kD�B+Z�"�+$�WH�E�{��QŬ���'DR��ଵ�&;eϗ��y�IeUe���o�>���˻���c]���U�w˹�ƻ����.�s}�wwwUUe�.�����˾]���N8�+�t�1�P�����C*��!c�cP�@h�*r�b��2�b,d�B�����)H"*XQǈE�d�Ul��Q�81J�B
J�d��"A(�b��J�0si^me$��n�����e�r�8�ۆL��&���S��y�ϓC���UV���m˴߲���{'c�T�<�}�C/\<�[�Ό;�����|ya���M'Z�'}�z�rv|Ӡ|:�'�1~n�w��[t�xw�ΒY=�j�ٳ��°G�g��t��^�'տq�ı�U���֓}�:K'N��O�i����Ѥ��I���3i����y��Hǈn5��.b�F�?�~Y�4��#$�,�q�E�b���D:k!����4;���Zj�����=��N'��%���M'>U������4l��c�3Dh��{xS�wZbB_��06u�N��I��j�NMxtw�Mr�]�-���f�UX���<N�����Ɔ�@9��E�E��*V�
!�?Vn����������C�2v���C�7*�R����j̐��p6��a��O3�=C�l1���];W��/��]���c`z���PˉA�L�LgH1YcB���ȼbԩ�İ�4;:��%;��J�ZY��SO����'�����Zc31{3�O����c�v��?*�G�S�I�4���$1/OJtM�M'���~�t�tl��b�c�WN�?��q13uV*�$ACq��d~�T�������G4gGcD!��1��"ֵD.Iw]��:V�(�^��JW�.E��A$.�j!�[kL�M��\��B��IRA�#����emº��J�!�1�`xd�*Jև�!8$��g#��d��Z���t����$���9d��i<�J��1<O�m*S����b���{5N�UM����@����?�H2ѫHQ���pc�eH��N$��V�5r�����F���âh�1B����i���������`J��r�s����;�L	��r7��i�a� ��Q�/y�3����#�<[P�2Wac�܂.$7f���s�Xp���Pvu�����*O�>Y�H�㒺�&�q14t�����ҫ��=���*6���3'���0�5W��l��UU���t�T���Ng����+\��M�4��WKsM��Z�(�9������Y��:y+�Z3��cUY]�ҧ�'gS�M'^�%M�3�PϿA�R&������p��?KmS���z�y�������b�Uc�W��{��5�\ˤ�u�]���:�\�gt9񞦏Ƨ�߾��h��UUZZ���gA�G�f,Y`����3�t0�zG	�)��`.�X<�Ǧ�l8���R퉚��n~Z���4�:>N�vx们��6�Br���٧o1.��Ji�b�Uc��n����-j���Em��%�+���B?�w.Hh� !LUD1���R����"b�Q2(�Rي!-�6�5$��$�y���*)HF!��e$��yT] f�!af"�YǊ�F%��Lw��l�p�j���x�H�ö��Ύ�T巾_���m��r|�~�U��#b�˙���G�c���',&��48.��ڝ�K���fC:D_��D+u�M�X|��N���d*�eٜ�S�n�c�V;Ux���_�Xֻ�;��ՄX��G�$��!8���Q���;:<�%N��<Nҙ��O|���#����E.�V����OYf'BWV:F@(.�L���g�X�~Ǚ���+�陖�W���&�}������7���S����ޱ�������Ϥ~��*�U�>c;YU���j�e~u'"\��/uuȜ�r\�/J��x�WN3����\W��^/�cNjڼZ�Z��ʮ	�^/K�I.�]Ļ�w=ӥ�_1���v���]?3��}i�+����ܽӓ�us�.D���Z�],⸻q�u���̷���^3����ݽk�L��8�-q�;z�!G�(��O�����pܮQ���x��*�8ʼ/��L�x����㼷n3k���c���{q��8�.:g���ͯ�w���m|�;3WM�t�M��Y��p욢&p�)kU���>��}�{~��Z���Wx�v%Ҫ��M��Z�VN<w�bT��L�U�CmJ�?J��>{>���ߧ;�בV�ֶ����ŧMunٕ:�͵P_�Y�.Uq1�Uw���|��#/��'޳��W��wU<��������-��_���in��[�������zy�O��������^ǩR��f�QR�>��eUV]�����������s}mwwwUUe�.�����˾]������UU�|���]��s���;㜷p��c�V8������FPy��UB�=���(U-=�.7��%�7�g�'!$�X�� ���F�b
F�����[�$�������z��';�m7��Ovc��5f�=��w�i�����0톛�~M�����u���4|��1^��⫅~����<� ���HG[����������81�L$v�1�7*�^u�g|�$��=���A�e�q�����~���)�ͱ���R46��sr���a=��,YP�r��|��S��ff[������~=��F%�v��UX�U�3ry�L�bJ�d�hC$-K��!H	� �~���<��[(���AX�Ő���Z�z�n�֚.E�*J�a\����%�EQ��b���$Z���h�,�X��,"i���A�\��]��GG�²kfG�����i��f��<Z��ڲ�m��o뷧w�ݖ��~MN�v�}^�:�Ø���qd&d�t,�9�1*���Ǉ���Ѵ�m4Jz�b���J�=d�uu�������V2:����/�&�~�/I��׺>0j����m2x�;��C!��z��!�BM�����]*�̟���N�I�y�ӹj�'F�km�i�s�Sͪ�M&�Óѱ��1��*�ow�8�D���K�����^�~ �9����Z�#�����|�.�o�Og3N�C��$��yą�v�A�E!	rRA�핔cCRY����(��\&����tS�s_�'{�d��:QUR�#���t6i�[k������O��)^��V:Uq�>���kM5�t���O��U*��jp�]�{�j6�;��Ԯ���j�j�#&e�M&)yTi�V�霦tɕ�L��>y�j�G�`:6n� #f�ƞ�\t6	�88�l��a�ˠ��ݝ�p:�[��A��z6
[���?R�WJ�x������{k�:����s�U-q�� u�j!�2C\\�HA��D�qJQY.�_A=Kx>�8�K4%�󵵸�ZPt��TLz�����X�l�R���"����/��b1��w&i�m6��Fp�hh.0 ��\n�����h:�N��H�^��p��M��k�G��k:�xy�Y|4�ό����GIHL���ѦP�~2�$�ܙ�/����r�D�,Pϳ�i��aҕ�Uc�W�>�k\c{�֕����&�l�s�>�x���b�m/m�۞ɹ.*ո�+������Xf���`9v���^�
���CO���$IF2��̙o�i���%e�7�ŉ4�3��c���щ���������l�ǉ�S��LN�*�J����G����o֤�^�0F&����N�N-V�}�y���~��2��f��������x�)E�j�rѦ%F�
d�9�h,ܷ]�%N��'[=?&���gH�5���&��;J�si���?;6�*�jW����J��]�V%��4��NYjU^�\�^�u���\���}rS��뇥`+���B�e��n��M�ʋ��6۵U�=�p�A�m{�d�����'��3'i���&��Ϻ[V�4��b�O�g%?Q��޽��7
��$$���9�j���-���J�Z��x�y$�x��z�t\����u9.Y�l�]����8�8�W���]��rzK��	Ȝ��W\���.���KĹK�;����̓��t���:N��Ҏ�+et���˭ܽӓ�us�9�ND��f^2q�Z���q�8�����>{���
91�Z���Z|��o��R�G'�Qɍ��r�>B��!ڎW���.��3b�ůY���4��Y�ܽ��yn�f׋��+��¸�xq�^5W8�^/y׽5���x�"��/�����3\��"ee �GA�!�b�!��b!����gx�Tj�TL�Ụs�4f��w���
!w��rk���#UB1�S�r�^��1�6p�NA�8h�2dc*����#P�B}���㨈@�&�*򚋳B
�?�N�����'HBg���(�]��E*�nB"(Tr��4zR�Pb�F�ɉADJP��
Re���&�A��$cHR�n�b)v(��&1aaԔ�F$,����ې�r �dZ�n�r��e拪�9��5hn>H�O�9�9S��+��˷��jt_O|��ߦ�vֹ�%�
����ýw�;y����yѺ@������zwb��kD��+Ʋ�)l�62�Ez��I�5E�L���*�u�D�.���u��{T"��#Ȗ�G!bV؄��2GK
+qV���V�-HR���˳�Ӛ�NFݐRҸ��Զ8��^��������ͪ���������]��.��ꪪ�����>�ꙙ���ߧ��wT���.���wT���.rݧ
�
⸪�\p�^c!9�d��.9��,d
�(\�D��Ѕl�d�*.3�!E��ۊZU%'�Ee-n6��򬤩��uZ&G�V�!b� �h���9!r`��!�m�A2��5"�,��7q��0���p�8�N�����а�X��ϱ@�;����>�<�\��&�N~0l��[��xgLa������;�]#e Ȉ�[�/��xmL���һa]��V>�MIj�4�.�qO�H��Ig�`.�z�$�It������s��Еv4W*ŇEhlOΎ%N�{�ڷ&2)ULſ��U��v~gIѴ�N���;75)��Ԧ��S�t�MO0Ҫ��F�C>���?��Yi�
�����#2�-�4��B�D���,{%ǁ��-�`NZ��r��t�!r��DUvɺ��T�%x7�ΪxV�ۇ���e})޲i3���J0i:�mU����v��U�,�g�M��YkG����Q`��h�3����6��ǳ���o����/3}kw��q�̬GǨ��Uc�n��vխ��� �$�g���nZ���ph�J��rhsCa�|�duCv����u6i>V��YF���T��Ǉ��m	<t0غ��
M��Ta�Ç)U[cv��v�1Ɨ�2u��B���֮ܑ��T�娸���R�1!
�r��m��.�����y��X;f$4!B���n���f1��X��0И�m�K?�X��
	'F͊��̙�����I���l�t�f�Ȳ�����1�2�{��5=J�������=N�ۅMύ&�u�{���Rj��5-�V��WI��~�:dL�&��OOSrqU�cJ|Ǭc=�uY�wrh���|f@Fi�~r$�Ppm��CR��s���c)���}{�6����vm����3�v����Ɗ("��bd"I
"֐����f|d
'��AL���{�z��a��jc���c��i������^�x��v�1ڹ�w��O��E�Σ[��$�r}2z����zw)���}O}�c2��7%)g����G�D�<���\�RE��*h�HrA���n�o��]I�O�0�a_J}���f\yUF�%Z����`��чF���:�$�Oɩ���a�xSD0dhΌc>�?���k9yK���ͺ뿒ge����z�mv9�3�rtΐ�����iS��� �4��#��ZI�Z)�=U�Rڹ0�x>O��ےڶ�u;V*z�ע�\���_;u�uV��c�m4�z�s,˚|��ʲ��\�k�٦-�'��Mz�Mrl�ZV���<c�7�yJݫ�SM14?�w�1���sv$B$�"�?��k>�}�w��n�YяUϭ�r���\�}�#�p�S^�"WO��I^4��%������z���̒�m�X��x�<�q��
��RBB��G�����)K:������v��u�4���4�>(P��n��d�>dq���|oG�L���l�FL�TTlm������0����=�4SP�t|��$!��X�1ڛc�1�Kk�3���-~�Rݮ-f7����6x}��Ͼ��˩����O��G�nt�o��3.]�q:K7���b���nh�.��q�3�����A�����%�5�QXeʄ�q�Ƕ|��B����P���۩��x��NO#g���OO�HV���B��(B�14-���+������ON>>>==z�<q�t���c�~_]�i_Z�����(R�*B�-V�b�
�^R�!Z�!j�j�b+�Κ|��+�����t��o��J�*^B�&������!B|S����r��|�\�Qiӧ}c�b�5��V�Aogw2���fΥ^o��o�k��J[)���|?�����w��d�Žl7}�Ot�{�N�>�ILo�{�y��ml�K̾͗s%ܤ�Y�+fVy��{�k*7p�BC/֟�:�W���o4��^��[��m����߾�}��33�˹�w>�ꙙ���߻�;��f{9w7����]�������{�s���\V�c�cZ��;!�]�Ɍ�2}�L�v�j��z�'�r�zp�q���,�I���<|�������ƕq�c,�m�\kX�njf����w5*xx;����B�K�vɒIA��b��ۗ�)����n:���P��!g���%�JK2'������G��C���psM�9	q�����BP��GZ��j�ӣĔIB%��/����J�MJ��b������"�:�����#)��c�O�G�w�{[ǯ�w�('���,���F��	��L�.�2;p~a�a�UU�1�|�m�l��m����4����e�JLA��-�.1�V�S�ThH�XEJ���N�D��[B#��x2�Cf��J�D*�����KU?�n)���b�w+��.6�䠠ˁ��G���α�g��GSIُg��U[j�;n�q��_O��|T�C>�? ��1:تC8<�tc펂�Y�4��˟�L�ό3�4�IgE>;a�>UWLz�1���.�嬙պ�u�z�i��C'ѓ���S���>:��I�Oxal-�|����5��:Z�5�&4�˙�cb�Y���+���m��z�:*g�d�+)�������c����Lc����Z�)x�[[9zq���ɉ$C(��������r��C�i��b�SDB?����'�,���M���GcF��њb����=���}6�ƓIM�x��bmO͛��|�N����c�!�:1��=�N� ��BA$����5C���3��ιwP���U�P������p�t�ϐ$���[�q�R$<%��۸�9e�t=L��oa��vMJ�k���#��A��-U�)�<6�;OyUm��}���4�mU]���n9��)lI�a1cc�QEX��3`��ќdPcc
h�",�td��Ƈ�x�1�c��iMQb�*����V��`6�6�bۊ'j.��]��Ȳ�x��*W�,��`�6�x�6щB�)A����tˁ��HgƺB�QF�$���:u�r�m��0�LӸ���`�&�R�n|\ҟ�Æ~�s�?��w�<�Mra��rNUW˓�5Zֱִ�q�8�,|��[Oܟ��ɳ�2�B>�g�V�t�����W�{�ըƵ�u��F���k�6aD5�4*f���~�%�Ly%�S����a�����L�3�����cݧ��K�3��e�V-���I���z&��0'��2�j���\2V��7�t�*y��k�)�Sa�UU�c��Z�>�VFB)qK�IO���.���8B��.<�����r�LO:ju�v�EnR�(��bpY�,\�[�2(�Q��ӔZv�3#Ac#�ѢIf�A{a1��:v����ͣa�*�lv�1������Z�<&�q�Ǔi�m1g�0]�}��>HYV"�ZY%Q5���[jv~O�zno�'M^1l���Q;���PѢI��<��
#��nm0�9«�w���Ul���n|��d�ͦ'��;ON�Թ!.HJА�ג��(B!�>z������|�^���||zx�\q�[�ΜqǮ8㎞�r�А��$!5�!R�!R�j����P�R�!
б
�P�Z�Z!R�B�&������*^T�jЩ4*P��(M					�^B�K�2\&�Q�B{��'ɚ�[O[�+{���GcM[,B6�"��a�-"}�>���8w��o�~�Ӌ}{Rf�ܞ��R���U!)&y�i�Q�L�P_*��%ݫ81�c�����pB�c�r{�8}E���z2�ϐ��b=�n���p�4��"	 _y��:�t��H���F��r��:p��G8l���wnN2o�9�Y��!I�O3��B�p:	у����H���O��S���$�2�D@D�(� �0k18C���1�:b,�"7����3FMe�����gQV��_S��Ʃ�ʠ�6M7ao{i�I��"������&�O��k6�OI�c�DcT�����y3u}+�k�iX��3y�����r�n����Eߧ���nի������"�EZc�j��4�@�8Q�U�n�D��X-�\u-Mk��f�2���^�����9�U���kj��;].h�w=j����cE��w�}͜m�uH���"��G�6�,߶[�/��7y�sV���1iQx��듂ĭ�<Ed��Bk�������m�����߻�;��f{��7����}������U3ݯ��ww{���{��7���wUT������c���c��������b%�e��E*oU%ȫ"C�X�72�TFZ򲔂��=��,�!rAK�NJ�NW���I����I��8B
dMW!ZM2�#�1ih�I\���N�(k�jպ�
0��$O�.M����a�S��/�Ǟ����r�^�n7�e��3�S*�0�,x�.�����gi���=�g�[�(��*JYe�Ad�0Bc24>6e�[�tpr���A��A@�B4g�gOO�˼�`���k4Պ�3�u�1�l�'��bk�'C�<N��S��bi�����#Hٌ���$0�d2¯��2clO��L��HJgA<$!7y�1Ǎ�AT�x���Y<8�z��X��c��x��,6j�Tl�i,�t��g�f~3��9��	��w�p!�|�b��Ć�i���O� ��ϟR2B�#!D��T�#:��a�Jޏ\|�	)�1���m2;��~��gI�v���R�j��'}}}6vc1�c�1�5���#S��5�t3�,|�lco��8�!$����#���f�pX��u��n>0�
ll��<�c��v��D���Pt0�HCC�Ӯ�$6kK���l6�ǜ�q�x-�&F��:!џc<{'ϿYpvEa�4���6q'��6p�Gh}<TS�#HM�Q�LZ"���"�c���i�dq�unxF�(M^���[1�>,z'�'�[v�Kkے
�d��6|!�U�FAD�&�pX�Y��>�,͌�07<Ι!!,vln7u���i֪>�h��q��+%�p��|y��I���'�L5+������?�C5J��C-,�n�{9'���'|�ө��ã�c�Um�X�>x�jn��D	$j�"|c��,8���C>�|&T�wL��-�l��I����{<���S�c�ti��M�R��Q:Ʊ�bi4�"b�Ǜ�^
x�'�f�ݪ�����u9��'LM'��y5&Θa�*��:c|6]�DW"��F7�|`}��TǸd�S�Ŷ4��%?t���S�|�ʉ%���Ŀp�{���|D%��S�'�L*a�|m��md�hl���F�^�q��e�#��cj��1�|�~��Z��7m�	��S��g�~��1%�T#*2�4<qC���dv<��|B�+*��*3���b=8Z�N�Yj�§�طkGq��p!��C���q�u�k`����j��/<=O*}?u��ь0d�hφ1�?n'썈G2^����G3v	<l��h�B�b#,��(��EgD�9g"mT�S*,*N�B����)u��b�e��S�$R�6R�$�sVx�rh�'M[q;�V��k��O��M��o�ȿ���Us3.)]��4t7Ё����p8u���#������k5���p�6o�ux��ӧ5g&|�)��cJ����p�{�c6F�nbfgc1ΰ�cA���a��vI	b4ܔ� �c���z"F)#��+�e2˫ߺ�п!IJBp�!q�+�M+*\x�$�#Pt��m���%J��l��o��{�����*ۚgS������J��f��Ӈ>>x��+O��~n|�>x���ͼW�+����珘�����||x�\q�/���Ǯ8�ǯ�ڸp������o�6���V)X�-B�j���V��B��-B�!b�hT�K�^B�А�4$$*��N�;v���M>i��j����&��B����[�|��������r�t�]o�v�^��9��Gy7n��F��{�B�./4:N�ӷz.��][���;��y�pm}>�c7k��=�7+��x�9�T���}���ӷnT]Œ�z#}PM�OF38�iڕ1T�\��߻7l�}�Y[�Og���:�X���F�9�y}���;��m}=\}�J�ު]u{����9s0��~q�˂<�yS��6*�j��j\1��7��D��W��ʟ�׺�-���j]���7�8�����M;���UL�������uUL�=�]���wUT�s������uUL�7��;��z��{��]��=UU=��.��.P�%�U�8�1�2���̾iߒi,�1�1d<o�F|S���t: MĄy,Cb|#ND�VkX�2[3���{��%��=W���d�6�����ے��ln��I�Oe�'o<˘�����1ڪ�1�3�~�cg�!?*$� �{2�?3�L4ɿ���ő�d$ʉAcdQ��*� $ۨ��ہp�ņ�
x\y�L�C����K@�Y��$�gs=�3I��ܦy���˔�O�w-����>��}L7!����I��4f{hh��8!�g�1����Z6φ\Y�\ٚ'��G��a1��w�}Ι�A	銦V�ɔgB��9)E��Ia�Qj!Q�w�Z4�:����L�k8�U��M�Y��D�dRb��m�H���,S��&3vYJ�$qC$DQ�UU2Q��U[�-�-J���9ɴ��5/����=OV�μ��Oi�Ð��ə���1>��V�'�)lZs�8ų*d���y]�zKkL$]1�>��.}�;���ZR���e�J�jĚ������3�o�2��ӎ��~4�t�����c���Aeߍ۪���)N|�C٣���[9�����յ��M<�x:۱����PXR�f��7ƶ}��[Lh�kU\d�dd*M7�˧��ǲy=��s٬Nph����^{t:g�4Ǧ~���0`�!��c�w���7O`�l7�;��ø<�����{:M'��dۉ��e6�昪��q4Q��"I2�����HbY��Ϙ��c��7;�q�f�16}ɛO
y��NMY�i:K3f��f�|����9GU���VDfU���FV�o�9��>y��BV[|x�<��&�p�7�uLcY<�%yWYf$e�$P_�L��s���1���P�8���K'����9r����95�\sK����ԝ�0��U�:�I��u%���45�O�t�ß�`��8����>�3N'}��8sA���aFG�U{�^���5h��9�~�j�|���hZ�CdT_�pǣO��dD(�c�5,ĥ����Mb���3�M@�/��+i�bi:�p�186|8I�tx%��n'���ne� )�3hm7;����3�:d���? ���M +f�#[���WC���)��3�Ça�*��<cכ��m��i4�����i6M'ɣ��9Ue��[�Gɓ����!��j~��N�yԫ�SZ�9Zf*��<?S
%[TX�e�q6��q2���P�R%���s����3q�����e�O#i8q�N�a�;UW�z�1���rsV�Է7�L���ݖ�mo"i;Nm9��:d|�������l4����ɪ5��C�	�eF�	�Tښu�{�N����ph2�����������Yb�Ɠ^�����1��U[c�1���+k���{vN&����t��[U��eFF��BI�s�UR��a���k��0��4h:9F�&̢E�!��q�P�3��<M��Y�ތ����U��'G�^���U|��Ț> b*�$�9��+�����O����[,�R ��X1Q"��:����+~55���UUU���ν�6�R,��TE"��Q�)$�X��`Qb�B��H, �P����"��(�7a0X�!EHQ��5����
*H��(�"�$�*�j�#����(��*D��(�(�J*�$�)"�"�R1$QR%	E�%	EBQBQI%D���R2�"��SJ�*Qe(SJ�J2��(�(�T���BъF%��R��R��Z*QR���*Qh�E���R���Z*QJ(�T�і����l�R�6�`��R�QJ��Z*RJQJ*QR�(T��T��J��0T����YEeL�el�Rʔ�eEK*R�+S*YS,��T���eEjYRʖTʖTʖ�)T��J-
QJ)EE(�$�E(�E(�E(�B�R�Y(�E(�E(�E(�E)
�R��)EE
�R��R��$F%����Y(�E(�E)
�R��R��TQJ)EJI�0T�R��R��QEJ)I)E(�E(�EJ(���T�J)EE�����J�Rʔ�eJYK)e�R�Ye����Ye,���R�ZT�L�dR�QJ*QJ*RJQR�QIE(�E(�E(�I)B�QJ)E(���w�	��EJ-(�E(�)"ʖT��*YR�K,��-e,��Ye�VYe,��Z��)e�R�)e,�����-)��R�YJR���U�T��R�ZR�R�R�e*R�L������,�)K)J�R�e2�RҬ������T�,��ԫ)K)J*)e)KJSWKn���)J)eR�l��YEE6R�e��JTQSe)JU�)J���S)el������YMJ����ԥ�ԥ�Ԧ�5)e,��Ye5)e5)e6ʚ����e�ԥ�����������f�YMJYK)�K)�R�jU�S)e5)e5)e5���V�R��YMJJR�K*�)E,�Rʚ���U��Ԧ�,���RZM%��d�m�ɩ,�MIdԶ�MI�2Y5%�RY5-��RY5%d�l�&J��RRjK&��jMIdԶ�MId�d�%�EY�,�L�REYd�d���ϫi�"��"� R,����RIRQ
���Q��4�R,I)I����!H��"ȅ"��$�XIH�Xj�� �Q
E��E�))�YR)�P@H xS���S��z1r�Ҕ�ZC�������! ("���,! �½I��?u~���o>�?.}��z��t?�%��>?��c��aD����u�{�?V? ����>+N����������t�OYG��I�-�ѫ��>��<�lYN�~_w�y�=B*��쾿Ѻ���� ?m��B~dA@?�"q}� @Q���E�����'�$��_ޟ/�!���A�%.���V?���E2�����}G�!�~o���@>cg�UD��?����$��a-�(}/B��)��ؖF'bfʚ����%%'�&����F������Or��������`0��%���}:�Î�?m� ���"^(삪]�҉(���*j�!l�$����(CL����\��������°��(��L/���G��TZ�B���T"��'�$�b�*""Z*���"Z@De���M~�|��-tM)��[X}����!D��K��z	��a^��d�~�?�Hz�~?����{�QUD�������~�>�k��o����ܓ����
����y��?����0̞��C	����BD�ϢC����|��>����q���?P��'�~X!�_��,��t���}	�:x~�a~�=C��g���UQ=��+�O���b}���l9Cǵ����[��C���q? ��Q@2�k�$!���%�v>�,�@E �II��{�ȘGP�ޒ\l2��~�����t�m '.�G���m������By� ��t  )@{ΒHO�����F{��TO���	�0��O�����'�?��������z��`���J����O}�|���������}^����
|�I��!�!�z��n����)_�z�=j�D�ߙ~��"H2b�F�X���ب���1�QF66�1�QQ�ccFѴX��EE�*ōcF�TTlX�hъ�EF�F�j(э�э�ŋ�1�,bƋ1bƌh�b����شQF,X�X�F6*4QFƊ�QcEcQEQ��(�(��Q�(���(�b�(���EQ�EQF1EhѢ�(��b�Q�EQF��(��1�(��1�(��b��(�(��1�4QEQEQF�QF1�c�Ŋ1F�4h��(�4hƊ(��(�4h�hѣc(�F�QE��Z4h��QF�6��E4QF�Q��ch��E��E�4c1cbōэ�,X��,bƌlQDc�b�Z*(�b�cb��5(��EQ�cF���1E��1b�(��(��Qb�(��(��cEQEQEcF�(��(�F1�QF�QF(���4h��1E�QF1�EcQF�1�(��b�6(�(��(��QEQEc�1�h���Q�F�(��4Q�4h�EQ��(�4h�XѢ�Q�F�(�EQ�Z4QEQEh�4QEh�E4lQE�1Eh�Q���"�11�b��F4Q�h�(Ɗ1��Xƍ1��h�1�(ŌcE�EQ�h�,c(Ɗ1��h�F4Q�cE�DQcآ�ƍcE�F*(�F1cQE1E(Ɗ1��h���b�h�(Ɗ1cQF4X�X�1F�QETc1�Q�Ѣ�lQ�b��h�(ƍcEh�1F�Q��h�(Ɗ1��h��4Q���1ch�1F�1��h�(Ɗ1��h��F4Q���hƍ(�b�Q�ƈ�F�DQ�hы�F(ѣ4E1F�Q�X�F�Q�h�(�b��EcF(Ɗ1E�cE�F4QF�Q�F1��X�,b���1b�h��(ŌQ��Eh�(Ɗ1��h�(Ɗ1��h�(�ъ6�Q�X�F(�b�Q��"���h��4cF���h�1F�Q�hъ(�h�1��(��b(ъ(���4b�(�1��b�Q�E�b(�F"�b1�F"��#�b��4Q�c�����ۻ��,z��(���=>*}YO����=���/�p�� �(�>�|�r�bF�cr��r+a�G�6���,���x����J�/�a`J~̦}������UD�}�X�q$�������������ꞻ�}���z;x��~O<HD���͙ �:�'�T~�c�O��?��!�������(�'�?p���@�~��zD؞�.�������3M'�������?�?"U``0S�֜����)���+�