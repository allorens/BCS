BZh91AY&SY��E���_�@q���#� ����bG�婢     |    �  P @             ��   (  @
 %IB���*�P�D@)AI P�
��E@�B@ �U	 �  IEP(x� (*�@�UP� P P  R���((� @  �"���(
 R��(P(��Q@�I    �� =e )�) �J�@5� �  
��P�
5T�[ (&Ͱ ��PQ@(}��A*�   �@`��@-%������@�,h�m�h6�:9)��N2� �f�F�ES4Y@k )y��h��� Т��*�� �)�  �;л(��@m�h=Τ (�1��m 6.]��ṷ� �j�\z�t+�iUB�a�j�P��p�p: ��RB�$X  kzJ��G� :QC�\ۍR��v�㆝=]�Ҽ�t���4ꀡj.n�����^� ��j
�T�wi@
{�(�UI@*T �)  ��iB�l�H��r]] �L�I�����]�C�ES���Pli�jm��a��
��$�`PӮʲ��H)�  U@�P(�  7 $6��Z�=��2�M ;Df� 	mF*�Q�����S2�Ӯ��T�*�5eIZ�kB�`ݪ��  ���JQBU*��  cExEP�Z�@Si7�hJ������p(Q cSPR������
6���UQ�j
=�J   ��UI� �����U-&�J�VҬQB�5`16a�Z��� YLҒHf�P���lr�D��J((P�P�(X �UU(��TU�`UR��4B�������W11� ƭT(�1URRb��QUKԕ�Р%D��
)J	Q<  ��R���M@��mB�R��EU+{�u
*U�)���Ҷ� Z+
 R�Ѭ(*eU��     	
L�)T� M0� Ɉ5ORUHd ����"�h4���b&��Sɩ�4d�4Ѳjzj<RR�&� ��` �b41z�U�P@    JH�j�U1� �  ���'���|>�o�D�bfbU��S-�Y�kYt�K���"�����))�N�W�@U�AT��D_�(�
��3&	`y�����^�B�� 
�2���OP_������za�$� D�v����$�@��'[ ����"�
~���2��2'XS��u�:�=d^��YS��`��X�A�"��:a��z�`N��Y����:�e�YC������D�u�:�C�	�P�
u�zd��aN��X���z�=d�z�X��� ��zʟ��XY�:`^��XG���"u���"u�8�=eN�'XS�)�T���:ʝd=ez�9�:ʝeN�Y�)�P�"u�:��e���Y�	��
u�:��`��XS�u�&�(u�:��d�YC�����
u�8dN��X�	�����)�D�(u�>2'Y�)�T�'��G�ʟ�T�0����`C���3 ��=a��X�#���+��"q�:�`�Y���P�"u�rX���D�(u�:��dN��YC���/Y����:aN��XS��������u�<e��XC���@�u����P�u�:��)��(u�:��e>��e�'YS�	�:��`N�'XS�C�)�T�"��zȿXG��1�A���z�=eN��XG���Y��G��A� ��:ʝaN�?�'X����:ʝaN�XG���T�~3��*f�*x`��XG� u�>0�eC�
'�����2���/�DW�  u�� #�P� u��(��DS���YQN���`Q:�"zu��
)�ES���Y ��*u��(��A��X���Y^� �ez�����"���C��/X^���eO��E�"��zʝ`�'��YS�)�T��=d�/XG�u�>2d�XW�#�Q��Y��� ��:��e�u�:���{��`?K�����K��̴�<�Z�tY,h�R��^a�9t�mCJ�020d�G^9cm噻X%�˽�4������n�Pc��[�&�yt���{5���´,ua;z�jJ7w�N��(��lS��s6����z�X���F��� ��0f=��ɺ�!˘N*��/$ř���Ӹ��W=y.���`�H��M�ZV�n��5 �0�r����2\oF#x������r�i]�Ŋ3��L��f��xeKe��pm��$ܫD�7lm��f^jYxm����V���J�!顑����t�FU�,CJ
�0fL.�m�j^V億�cb�O^�mF³�,��	-�p{�XDi��mf^a�]��[��c�{jD��)�B��e��r]��fX0��l�H�7W�r�-y�`�Ik�Zn�d�!�`���xhK{n��ipF�\�IS� �̒̄�5�+��m���4�Xo!�҈���M�Ɠs {[x7�F��#7�oAt��e��݅���o/M
z)+���uemf^�L���i��7��Y$��^�̻�z�TtP��L�ot���d�V����V�LՉj˺�{x)�L��Ѵ,��j�XA����,y��Z�[ܫF��K��7�1����Q�T�=�5\Kv�ܡf��d�`6��̭Oe<�z]�� �j�\��M����ZH��J��J��I4]�ʖ@�/rB/E'��!��y+,���F�� ,ѕ)���	q9v&��� Y/v��Z3(f�&�l�s2�j�n� �uթ4��9hf����EY[��J�$�26�J7W�V=��f��h���㥘�iV���u����Cv(J�ʼ��V����i�т��ƛW&�̛��면v�˳�*ՇrB�	ChK�w��I�EM��Y�U���^��ۺ���/rVD��k�X���R��e֬��mT�,�F)���@�Ua5���`,�F�ne�[ dJ��a�-�Lڲ�V�LmkW5��$/)�m�qe�l2�d˷�G-g��;GK��(`�L2v��.�3,;��Ɏj�c�� -̔1ۉ�4̼h��?�d�[:�D���W���"P!-�`֡�N j�f�kup�/(#�)[�����T�/n�[bG'b�2�b�T�������AV���/@Rm-Ӎ�ÔʸX���X�;zR�F��Befm&�[���yBP{WW5�͗L]!�h��/&ի�y%ƭI+X&]������Z�؁Wg+Cn�vͫr�4f�-��uئq���˵i4��j�p��%�� ��*��w�b��d8�`�ZV�P�CkC�P�����a��ǂ��l"�[z���1X�Ĝ��4�t�40	���u��T"�c%�%zA�����Z4K��[[	Q��L�Kud��%��f*X�``e;�*V�Ff������Waӛ{�&i�x�YG�2�CfZ�&]�i���ܰ�Ġ��{@�\V��S�\��+�S�n��`�Hj�S��V�]��,ʡ`�N8�:j* �m��W��Mfj9��Sp��B,���RfJ�ё�˦�Y�y%;���Edu��۵z���U��ǘ �.��*QیaA(nJs60�:��av),pZ��l��饛+6�q�5ff$�Hf�y�EiS��
�ybZذNm�ʣ�n���m����U`*�M�ѳQŗ��Y3(�����sS��ٷZ�t-e`ڲ�ݸQXKVh���fI@�C��C3U,��6k+�ݬ��>(U�Ѷq	l��f�c�j"�E(6p*W@Ƭ����f���ՙ#�-m�"��Ш�ebWZ�)2�b��٢�Љk��i{M`C:l���G5�W)!�d���7Mc��b�e৚��1޻ҍز4����E��l{6D�V&���a��7uܗ[y{�����Va&�ƛvH�[�u�ɸڕ����DKw+'a)�wD�9�un^�6◊)~$��e�*���;����i�V���ܡ�n�[wbڊIG�cW�/�K�/w4�L���P(�7X5CYf�(�H�:I�͙�V���������y�ǌJ7CE����]����C(�L]dW
��3QY��UM�1�KÎ�$Tv��Í1W��;1�l���pK�ѻ�c�'e�L��Nާy[���٘��ƕb��M	�Օ�B�weݳwdʎi�9�cV�t/B�:U�����P�ҺW�cgJ�t�m��j�0��*V�Fj�$CqVG�1��� ǖU췇%j�+ۋ]��ֹ�z��C�m�jd�ܫj`I���i�iʗ�wM�
��N��86��^���[X�H���V�,�tPz��\��Q���z��ԱQ����hH*ȭV��.�nU��T���n��m�!V���rV��$�����X,�6��!����5��]���*��6��Y���^ܠr�ecKb-��L͔F�B���b͠@ĉJ�bY��+<��J2�+�M]�t�8kJ�FEbY(R���r��n�����\Kwv�'��P˽Y�b�ZeЎ��t���5�*�nՠ�R�ݺX�]$�nb��˥S@��*T�,�O(J�k����)3�Dۣ�G))�ݚnG
h`9�t�siM����1�u��b�bF����9�-�i;[�'㈬0(F��Y�] 2��X�Hs���	D$��7}v��s5vY8rP�!�%�be�0���n�ve�QVn��al���4n��+E�lx6��u��Q�fД�ݗH�;N�ܔR�\W.GN�dT���Gj���I'1�sd��{a�N��`�e��V*m���:q�G}�h�mh�r�C �ra�P�&c�r@M��lO#�2nc9K��P0C�H�UKoj���z��6�b7-�{���v��B��s0̽ɡ���u���v���tQ�s֤ŉ�@g)�ڄ�(-���ܽ��1��l�mx]���щ]�0;���^��/&Y�d�ӂ�ۧc	�׶��X��rVn[ Va;G�^ŕrcU�A�@F�x�6)2�z3*�7Ri�[��P�gr�Y:�	gEi�b��{va�����<�)Rݼ�X5�`���Y�b�H�-�����HQ��S˽RÞ���`���(���1zm�X"�6�@�Z�G�"Z��s-�m�ݻĲ�Wq�� � W2Y�E�hc�������^�2��qT�z��W�	S䴳���̴�
ݐ��b��*��2��mQd�-�ۨ�Ɔ��2��~Đ�Fw���hYA�W�f�v�1ش0�o5�WW��Ҏ�ʏwZcd�O1��6v�MB�A�8�攰����&�,L�@mB��dږQ��r�
f��z�e�a�Fm��n)��M�O|��3�C��yu+^2A�kD��yg/M�f��U�.\V�m�B�[f�)�� K��d h�7V�l�3�t�6������ݝn�drȭ��R�V�R���%� �:�&Ɯ#SҜ�׵���졶)�h]K�!�Ĝ�u�)��#���)`�q���Qn�%�`RɺI�G��j!䛺䲫]Y8eQ�����ӧYv//�$��\W����CU�v�x�VF&��-��n�8-�)�[����o&aw&�g/.cXNTJ�nʲtǒ�l�
k"�6�F�Y� #.�[�xJ�.���ݩcr�nք��U�&/��:�v-�җP��%�:�r�^\ٲ�/��6�x�86,�0֘�OO8q��Δ�+��c5�b�����)�^�.�0�kJ�6�Z�=IA�.�um��3����U�nk���V59+o�g�ffݫ`D���D�eVeա%=6q�ܭ	H�ڀ�U�[y��*�ܫ�Z2Q��s^8ޚ1��uzeZOј@�W'��Wy�sK)˼��0K���b:��e��wV(ne����)�������n�P�u��,��:���Uy�t%[QA�wn������	
��Y�]�M�[�9f��وۙt�h`�Ԡ��
B�c2�#d14�
x�T�F��QP�o�+�t���=�{R�+h͏��v�4I�H^�A�!����F�a47$��oӢ�w��ɷkqd�W��M�e����H�R�򳡥%�j'���"e��]YZHH�5x��D�\��d�ue�����1��ZbͷpQ��.��Ù.3t��}Y��J�NTOb���w�Mn+R�l��ȤN�.� sR�hm�o[ܫƍ@1�nۦ�6���eDh4�Ec	�2��+�4h���K���E
�Q��x���7�U�H�a�w=�6ּ"�7$�n��!�	V����[r�a֊�5I���1TW(�,KbeE�!pp�ù0H��ù-�0�K�4J��^�V��'6c� ީr��{CFA.�䠑[vPĮe�Z��ugXb���2Q�q\�����l��k�7l�K2������Y�u��d�[ܫfi��sb��Ͳ��$�Xvd*��YB��ojG�X�&
v,���<E�v�N�%�=>�Q�x��֭2�"t$��F
�Aͅ�Cnj����#q �+��(d ��YXt���V���x�v/׶c������z�1�mL��b�&��Ë)�D�[�Ă4���1b�j�0@�+^��J	Y�[��j!�)�M�ZC6��l̳��VtJ��L�B���,����B�ؑv�
WV�x�:V)%J���J�-*�n��*e��3�e����N�,l$&m�� ��-�ڹ�n!AǛx��t���U�-V�I+2����Pk.d�����"���M�R��n����{;jN&����˴�gRͫז�W�Y~��Y����Mʅ�V`��.�H�@z�`*(ZU�@*X����;�2�á`��N�A3��1Rocz\Ѵ���Z]M;�̱B�{d�#��mE����fyf�ڷ=�q1��st^a��6M���"bF�KL�%��O�U��f�^�햵k�$�7��*ե���K1�d�����Dn�N�к�(\U�&:L��"!X�^�#�q��54�ԍh�JfeG��Ѷ}�[�-[<fe6��H�V��M�i����t�c��4r�mZ`sn���S[[���`Gwf*��0c�u��p\jv�9A���_`�DM�=X7�v2ؽH���lD�7]�,�.8�[�Y��o6��b9=<&T4cɵL�$,������/%d	5n^aL9���B�4���7�b�9���M��!�9��E��Xv֩�8���7^]&�w�C]2ZR����$��sX��֐��2�XyZh�E����Z�2B��c�,�P���n�Ձ
D^�Ƚ�tUx0�-�e�1e�ת#f��$R��}H�f��n��p�U#���*�����z}`Z�败ݜن�������8�أ��(a�f\N���H�U�dDB���B�AT�;*����k1��4ͻʔpn�,���eM�ּ˫�Q�-�,��� �����4.�ǧ	�T�Ŭ�U�l�)�Y�t�ݶ�X�'1`ne�R��#L
2!���v��I݁r�]��F�4msd)Xk&���i�]D��j���9cY�;�dɗw[r��s37t�]����ٸ�O״joE��/�w�6	��A�dlb�P�j�*�I=C\�.�iY[OSr�ՆS��)�˰A�N�[�j��%�:�LÎ���bVC�XY��im]7P܂�6�LU#9�e�ޛ4H[Bf�w���~�Me�*ִ^\7�lH����+r��C�.�]���
�9��ַ~�z�'r���);�4��z.���+j�u,w��c�^k,�6#�ȶ嫌�Z�+�K���3G��`#1����ۿTv£W��t�J[��ݛv����R���f�x�����Z��;GiM�+p�ƂcE�6�K�LE:�Kq�O� A9��k	�[W��m]Ah=��8�а��7SN�h�KR!,���5���a�kTаWu��%���a1+u�ևM�lȆ^,䰪El�˥�4ɦ�M�V����+&�JJ$!Vlɽ��èL
�U��jY����zY�4�*z
%�� � 2+��u`�b��#%���ͽ�챱��u �J+u�1�/ئdpұ6�OA���f\1Jݽѳ-�m^����;oJ�m ��xqe�e��\�ij(n�̳a꩸7ʳ4h�P���c���K��1L�����n�L�2��hͺb���IW�*J���.�	<Mł�d�J�+ �n�k@D5��Æ#F�0�AejX.d��L�@J�Q�!��թ�7п �W+&E�བ�)d�(�wq�4�2jܛy�ud��8�V�]�k`��VF�l�L���jީl��[e3�Xy���K6�X��Ѭ!,6�o �m'>f�7��%���{"��²c���p��P=��Zh���A�!��^P��ŌD�Qh��݋~�S�b��UV���r�U�Ӣ�㢍-�f��u��\�hA[Se�E޽۽�`�ZV�2���V�j�-���E��J�K���h,ſ@�.����»Jӈ�=���tR��.b�Z�X���,�ܕ%Hȱ��ac���"�m�Y-�K,��qL���d�V�7j��,���2ʠ���2�G�;œн6�^eEٌD� ����`�[V�zZκ�b�P�aF3�����.�e�Y��pE�*J,�"ʂ`�&�"��@-�ǈ"
�pK���6���K���mG!�p���((MHD��W�ɚ�������ǹ
�E�J�܊�\��w%}��iXoO3�B.�.���nP�6��{sC׶f�$��l�9�a�T=�a��"׽$#i��7C���tb�NoI�fq�v�Wt	>��0{#.�/A�n*aAtfH��!�Kfh] ���,�{}sMi-l�[��ޑ�qh�N#l�NR�}�Bt�1�̎6M��*]�	z�ݝA�	��Ȍ��X�03��ȱ��a�,S�������Qf����aY�?[�ϣ����آ�x���^��{�	L��~y�/�6�m��m��m�y�J8�gC+�us�N^���Q�h5���5B轭�̓����v[U��M���Z�jFe�T�'�+��orsIT�a�SS1C�'e�ј)�"-��t*[Ӡ\z'@v8`�:��m����9c�i*��
N�eDP;J1�)�b�)	�e<��f(���P��"LR|)�Q;ջ`h�ґ�^2cb�5[�R4���6\^`�1��x'g`����\��	�)�RoRz���ȃ�Y�b��B���L;�U)�r��ON����ˆ���!;(�o��{+r���D�Vg7{{��g>5�N\C�Kg,�㸤g]n0�nb�%]�u¦l�n�Zt���%��`g�����v�ne�{�\Ytu�R�&��8謝s�d�?v�$F����Z�-�������ЙnȫWzf�. &�Ct��.�G�n!���OTb���b}5�DDE�b�u��Mr׳�R�N�56Y�z/;�`����dA!\9��"�+,c��1\`�bwf�m�$��O2��2�R�-*�{�p�Q����\r�T�Kͮn�m��:t�fc�v�6���G�Z�-뤅�h�J1��󚴯d�1�m�ӥ[��˟�w�'�ޗ�C�x�yt�]��ZjK�ʺ��0�Ᏻu��;׭�ż�m�ḕ��F�)	�b��9�v'P[�P�8���%wǕ�ݑ��{�˜�y��jܠ����ų�\�^\����ͳ���f� ��*m��B��Z�h�ʪ��nS5�J\�X�MӁ�)������y4���F���ݖgb���OJ�*���"��������#A�F�r��9wm���K����<���+g"���6p9_K��gF(I��Z��-!F�(u���"����j*��w����Q�v���*���!�����Ի�L�Pc��.XX�F�w6�a횲��6M6�I�U�%��[�ц���	[��ѐe�lY{��3qYT�v����b�%�)��i3����,�����Ds��<]��͓B�H-�����%6��s�˴�F_v �+(�ec��؄ɺ�<u���-��`s�4`�L��RLy/.��o��5}���t���{�ε��I��=��So�	�rj*u�m�Gd�9t4���R�$�]�I����B/	���
W+nx<���]n^\����	u��n���bhZPƺS�
�uȪ\��!��mk`�9de,�5�l�j�tg�C�\�����M*�B��/B�g(XUOM�[nœOe��v7�7��V��0��ǥ>�S-nꎄ��o���a�qo�D�+���ק�����Ơ���C��X��o���_k<��s�ᆠw'B��yn0ڻ�gN���˄uIej�Lir�@�P�Ɉ�];mj9�^����w�a7N���Sx�fYƬtT�2�/X&�l���wU����}U�d]^T�͉U?V[�34��0��[P�tK�zww�.4s̻(ot>�/h�G6�aKl��u���Mv��iV�N��|h_0�x[W�!������S�b�lΊ��8�eX6��<����3��3�I|��̜G��\��!�/��L_�Ȍ�P}���Q)]���c}y���[ia�0�x)]-n�F�
}cjsC����v<��L��Y�'p+Ί���o1�E���+�Ծ��k������"X�8a&��Ю�#���� :#o-1����2R]��� �j:k���ݪ���m��h��
�����xZ�ا��KB��b
�3�Qz�Z�=���a�`p�7rub�K$���6�a�wf,k)	v������zm@,����Ģ���ϱ�27�[�\��o.jr�����L�,ۛ9�+��A؝xe)ǶL͠�G�^`�&웂�z�a�̻ȳ��Q��j��LDm�k	nY��e�3Jz��4�>���[� ɽۖ;�����݅{$��/�Ut��hɂ��rm���v·�ܹե�զ�α�
]LxQ�.�/�7N����k#~�K�:Rƙ�ȋ�1���j{� �pU���I�ޘ�=�M�\���QJK��ȑ��U6,�(։j+v�
D=�,��<��<�ոP�s��	������{������*J��c��70�{���`Uzp�[G!`9OMЫ��t�w�2�H1�IJ�wD4�b�h�u����7V��}3&`T�6>��xtz��q:���m���9���ԥmr��b�����/{zm�
�1^n
�~����]�2�}�I����U;��{w���*�;�ѫ�N�����f��V\����4<`�XZt��֩;�����9�����L�*@�z��R�x[:�;��f�̲�>9��W�s���p��Y��юv��5a��n�&�uٰ��HNk&���F�X�cK�zz'ЎZ�����G6+��������a�LP���`]�1Y�<�ug`w��U�\�Ŏc/Ul��ٻX,��g����5�vԼ
��*�0r�&+�|�#��vT"ࣻW�y���V�ܹ�.��Ԇ��H10å��uUUfI
��D�Z��+I�$;Ҏ�0i6����z���j�6nAɬ��t\�gy�����w�e�Ւ`|�CbvT!WM{��a�C�Vk%r4Ӽ���ɛq�`'J�����+1�Sh]�����>z��Vcܩ�k:q����{�%{z�Xդ���*cTV�-C/u��:�jS��0��ł�����ɩ��5Tڱ3�>"eĻm�����^�d�.e]tb��Z!f��c�{���w���aZ���<���`y���fTX/I��<�)Թ���M��˽�t5�����ɳs*��u:(�����GF,�%�Ȅ���v�*�oe�9庱�C���+�fB>;� >�ms����{�� l�9owWu\k�9�N�6"�5[$�e��\1v+�R��D��V��,i-F#ulLå�Q�5����sr��H��jMf�h�,��s�zP�}��3`φ�|H�x9�p^���U���Ǵ��d=�s.����-о	��^��fǹ����^�o��2du�����w�/�w(�Kx�vgK�R�[�d����<�g�&e�<�=���꽸om���Q��,�g��-�g���&�t�+ -S�#8lkks:��0�z�s��]on�ZR��Κ�ѷaW^�b^J�y�]TW���u�rw�&6�Z���&!=0f���hL����U+b�&]u��^]]M����n`0gM]��n�h��]wy�Q�<������U�=e�}���7&��8߲�͗/�P�ж�f���ڠ�&�oI�V�^����gR�N�gYf�a���>|l7m���b��*�*t+S/%��DnΥ�d�����0�j����I�Ύ�n��cp�gj!r��,�O��Y�v��d,��՗�nh¡�utrm�K����j�r�M\L����5��n�f,j���ͩ��^�i�sZ�EĬv�)��S�F�J�Ѐ!+6��t��@7n��¶n����	�p)c�U��ם�D���4�uŬ!��m��n[dC08	��w-w����T�:v5�]�pU�u�_sK�)RR�3L]��|�-wVL��A���H��F��и�H����n�}�M��qe��R����ΰdĽܾt�Z9B��.u^\=4�X+�ʻ
i��x�I��¹��tS^��3ݰ�Z��W��>�th��(=��W�4���z����H�w��*�q�d:)��tQT2����;�J30��Mcj1��gu����YdjQ��2����X�R\]�ʾ��ůz���d��pM3N^��;ʮ�����9'�Jw0���1�
�D\���d2{gi�D1�Pns�}����*T��@Y)����-c�4VpTM���z���{w�7ͧ�gX ur�wu7��\R�w�T�E�rJ�Vw�)�X��q����|�u%��J�9�w-�PQ�����v�/.������r��z}R�k"��'f����K�=�Od}����8Jy{���ʫ�kq�t$=�ѸP��;�ottX,�YH���4w���81�kkVU-�3��k\�BVD�����4T� �X��M�éɸ]v�z�=.gd�Ѽ����hi��ݭ<�V��I��6��p����rf^+��{�D�V���D�
�Ṽz�J�e���*�w�W��M�[`[�㹍�����V��Oj�ٺ��`-Ǖ�4А�k����k��2���a�i�:
6I��v�ꆭY�Q��\�X��7�^'�MIط1�����K�ӗ21n!�<oF��[{jb��z0���bFc��w(�-�P�4n ��k�d@5W�[F�Ӳ�M;�:H�!���Vv�j�bՎ _�sm��{up�v��%i��@W]�lR�b�3�Nۭ������9A[�[����J����]γ�"�Z昧x-(�˧�]Q��|N[|8�X޳X��F����2��=���j�D`�2��2��Ќlk�T�b�qH�F�
S��@ü;$��#��8�%'\r��4�̛�hG����{2�8t����'����VPM�>q ��w���$mK���£�*�eL����A��˫�����+�h�h��ydv��]akx|������m�;	��ft�=iP�}�L�@^��4`�ܵf�]�&��� ��7�z�]���+��CT�OXp�n���=j*���gl�LCK,*�k���ӽ]Q2mJѢ��3J�ͫRA�,wcݕ2Ԍ��e���s"�F�Ȱr���Nb̩)���3mwm�%.#Wx�R�U%����B�n����fS��� ����{o��mv�dۡ��Q�`�un����
��iW�2\��ޥ�u�n�łB���T�y��m.W\຿��;�2�A�W�6#�`�{B�$b�z�^-�wnI��p�� uf���]�C��u�^��kr#/��m8��E��W0*=ξ�T@�x�Y���+��Ʋ��u�C�trʀ��ed�Z��=�Z�5G�{����a4z��B�v��M���qj�:2�dn�6���5����=`#�����P�<�	m��ͺ�W
o���;1+GO�s��qɔMn�UGqwmnl.��8��s����6�K�zmT�s�-��M���"���ȉB�v�,�$�ι�d���i�5���d��'`��-����&�AX�Ӽٸ��"���V��qe�¸�������r*`�H����\��|���8��7���G�<�H��g�p�cGm��.�n���ۭ}��	�P��,V��tŬIٽ�a�&�̜v6�:6A�38���{J��EX�����M�sj��7/�n�����e�ɘ����Q�P��s��p�{��Ջ�9�4�c+8زo���ǝ�p_&�ge';f��,z��CK%�f)�^��q�XVSgTD���v�mʥݑ�^j�ј1����6�3���v�9�����e�	�w���23nM�{f���F�W
�`�xi�Әu���W����)���Ⱦw���Ji^Ub;�N�х,m��ŗ:Y�����7�f�n��h2�]Jf�r�z�WH��T�e�5�ڰ�P��+Ms�[�H�n�۝�Jk�f����^]j�N٫�Mu��n�[����9Y�6e�����;�)�	��+[�v�����T���4^���:&t�b�N+�F�Ѧ�(T�Ø�{������9+/��dW����V��b�i^ZG�:����|���o2q�Z����A��\ރ���,wh���K������☧�[n���r��w�f6.��Zw���R�#0�f�N��wl#6��k������a�k�vkf�pn���Ȕd��������]�|�ו��{VV$�)�b�f���x�j�R��Ԕ]��/W=T���_LU���A�j���.�����c0�=�wm��4C�6����;"E�zzn��vm�Շ��©�a�'��&a
��N\w.0����sp��2�f��7�{bR�G���[���D�o�B�+�1�� w��d�|�!!�ӳ�A4��v˛����b��*��cѺ�ó�x�.��=�N3�^e՚�X�4�^�Ҥ�lW�Emͥ�Ɣ�^aӛ}N��B����5�h�+�ww�A v�㮜ࣔ�;f�t���oRF�I Tu+6ԛ2�;��L�ز�ЉRE�p��*0(E�%�v�޺�{z�Zԋ.H]�v����wǑƞ�lܣ�5Rq��Z�j�m���M�c��bf*�J5ַoZt�zݶ"�Jm�Ž)�l˳	 ��㛊`�e[sU�����<��ԘQW9{��L]mE�����sN�+�M�a�2�����|/���f۽9�\5f�{�9d����wZ���"�������U��Xּ;���Ŧۓx����)�.�n1[v��t����%6��b���o�m����l��{��s�xRm6�i��m��m��m��m��~���+H~_ �ϸm�8���.�4�?=��?�a<���=��lG�������Q�%=�C�+�%���"�t�����^K�~�K�>F�/��G�~��|��������y�'���_����o��'���`$9/���{�s����~�>y������=����K�Aq��옂
 t݄Ӆ�"|r5*����}u���י�US�Z��ad���qe#:Yeէ gy�_���%8u��W�5Z�"iO6��w1)U]��]�3]��ۙJ�Y�־{�Ӻ|�7u!}w��� �+h_)%�9��B4��9br6�c��}&A��R�jlt���d��Y;�c1��E�6p��Q�Zu�w&w��]�k�`eoi�캫�(��{�&�g8
�"�v��j��2ѱ�������X�]��SV���8%7�L�bT��ZA�;iQ������o���65�Ce��yR:��;�wJ���ۓb ���� ����rmu�v2���n�
|�Px'K5���[u����b�n��9ًfR��=}ZLݬ����[�D�w
l7y��� 	jA��1�����P�rls�_3���f�tV��Se]�m�e��w�u�Df�v�t��L�p;��<���(��j�_V�!s����T���	@tG9M7o�Sm�䢫jG�զXx
d>�xC��ʬ��"gN�w�$�VA�T�U1�#����ZS�:q�;]#w�y���Mn�ʠ��d�&��-C ��C��1�'����pa {x\�.��4V�:�f�6�[RnӝIM�.�/Lٲ�q��N�O�u�tuY=�ǰT�y��Vgu+�F-�e{���u�p��6٩o������"]4.��ZE�����!x�������x��蹈B/r5*n�o�u��z��8���IV��^��f��.��|3r�p�e��GAf-,M[ُ�P��4\&�.�N�n�p�&̕�pVu���H�f��K]��P�K%�̭�0��*��v�z���qۃU�4rغX��ۦ;h�.�rXOdֱ=;FE	�ˍ!�nҔK�*���i��j�ݳ]~|��^���aW'u�۬�/�l���|+//տ���K���)�;�x�+�,�6�"���`�_i�J�����ڳ{A����f�����8E�7�c�ڦ}�9�w���b���{*U"a�Q�JŢ�ͷ�Xp��Fv�s�����:nR��n	�m�$\�h1���=(D�H�j&,�U�:�|`ݢ���Wg�PJI��&����c��V�N������F̩#_,W������=���9Y��,3Og;��v����i��%��R�o�O�����-��jU���خm,WH����2��\{\vh��pJ�zP���U�v���J�ے���;6�e�i��;8����A�H�V�rS��^[������;8�wf:�E�W�3lvIEY����r��
�d����I�F�%
O�GA���H:%[,�c9��:p&\�	�xF��1�\핽���!b�m\\���Odv����n���zU�=��81̾�s����Y[3�&^���`����N��W��yaQP�A���t/N�sX/&-�Ѫ�Cj���;"0n��P���}�^vjû-�vx�s6�ee��e�i�틽�{�e�ۇ�r��P��!�7X�tL���!�Ub%B�Z�����N'��H� �l���*�44�T0ƩҫS�r��*�1�b�*���D�Ԭʽ�:h�̹&a�v��q^`.�q޶��bD^t̮p���v�uh�8���`۷��2��:
�j^ɘ�1�{e�켰�*:Fҋ�K�]����)H#'{MR�o<,�k�/!�,V�z<�ט�İM]����hv�\k����l��5�&1��kM<]A;d��e�-��]��,�e���h�]m�MgY�sy��n�VLT�N�jRn��+��Z�}S�����1i�-��X�1�p'&ٌ�p���n�eK�q�R�M|ly�tZ��a`$�"�N6��ѳ<��͋�[�6��,@���>EE	��e�pY�XXB�NHV�ǛG˸#�B�8�P�'�CV)�z�t���	�tR�N:��p�JʈُiR�t���=����(�l]EN����W\D���2�Γ�מe�G8oN�J$�3U͸��5n޽�F�&v��ø[n��:)���9���n�a�ԹQ(W}v���:`�I[�*�������E��<���q��|s����/�͙b��os�T��wZ�� fޥh��ѡ���%���gqA��wSN���V�-��T�ݬ�/;1Su��2�yZ����ǽ�s^�Բ-}W{I���'].C���ڀ4�nbm���j�ޮd3�������q�pT�<�J�나�3�5sǱ��|%�.B���9����\�72�wt^黵7/mQ�]�;�Z�lE�T��:�\Uuex1Lۍ�;mB9J#+;��/��-t���<p^G31�\zr�+�{��@��0P꼨2���̳M&�i[�C�؜
F�3K���V1գY�ܶ3��Mf5\5 p��P���HY}���sݹŃJL�]~�-]�СV�ةư�4!�V=�ma4g�	�ލWM�1M_%
���9�Qp�m�Mm�T�Z[wZ�Fn�w�
�	)'B�؎���ŗ۩�{3:��N��XJ���Iǫ7be��KÕ��*q��"����~K����DQ�F��ۍ��M^�vF�{�xqA����{"��ԑ�SE+�O*�����9C�c/yԡ$y�]j��\L����^�evR�q���gq�K�kL꺻�/�^�@����jl����9ю(ɸlcu�̉a'�`�5̛a��q�r��{d��JHb�Q�4��Ĩ�;]�[iU�]��E�xh���`���z�XcuL�Cܨݸ ����
I�܋xee��<��d��I�Jc����k�X`1�-����(��B�۬�WɜAPf\Z�-Ỷ�3癁M�ztIR�{2ښ�Z�L_"�|���7,�%ӡU��W��S���{Q"�.FAJ�X��Kh-�k��df��̩{F�66�]������P�R�[w��
��L�&��˽�3��zh͓z/`��w�Y������뎆r´�w��\�yc6T�v�l����7E���S�Kk\�0Cvn)^NF�[�4���8�l��k9-����:�D��4q۰XNЧ�5�{w�2a+X7���܌J����k�8C� Nf�IM��"ң�f�'Q��sL�o��p8��;�3���R.*{��l�SI@�U�ֺS<@�G$��~7�;l6ske��ݜ�z;�Χ~:�\�ti!o�"]�a�VWv��{t�5�e$"�am�� k2���)�.1�~�Ee�Al�M��٪K��C:�={�������h���թY��>���;�]���.]����ٗ�BJ�C�,(�5l�u�Є�j�fQmf7|�Z$� uwdͅD��;���G}�=�u��s����ɵs�g5,�E�i�DfI5�w$J����f��"�����ʽ��WWl���yƊU7*n���
n���s�r���}�;F��&"��k��,!����������jQۙ�-L���"��ڛR��r��zv�c��%�ew[۷��Z㕌�iք4����Ƌ=32շ�*�ӎ6�{)a�����J uVwB�D��:{�o5�6��7���d��~���ݹ�{o�j��*
��x�P$�x5>���[�O���z����'�JT}gs�x�:�gen���
�=1��E�c�w+�V/�q�V�S���=h�agCG<X�uZ0��@<""i#x�=��df1Y�������gq{�hu��r��7*�W����0��p}R�x��Ȉ-{k%c���@ze�se9ܤV�����u|H��WSzд�\Oz;��8]�7��kjX9؀��b�ӥN��3����&�Igx�<�b���!�ؘ^]��u§d�!�0n�� ��������7�1�Y�����G��MM;h=YLp>{pc[k���ƪ�����{m�0�NM�,*����{�3��]\Z�nc���к�I�͝�f�wV�BI3Z��VK�g�������q-�d×e��3s�b%B�)��[1��\&6oM[�+G�7l��j��
������y9M�}��wY/u���.ˇ��}�+���i"����h��[�Öo�V��;��VŹ�w[4�����giR�H�T��s��{��	`bL���Q�ql�Na�W�,�W���M���FJ2������Vٽ�����.�����e�w���L��ۡ��fd:�2N�M��y]���Ɍ��cW�VunBY+�銴P|�7lqT��뒯q�Tr�.#`���i�;�R�`P�BM!��u�ja�q�##�F��j�����bs�3��]�$"�����{�+����l:��R�����VT�h6��q$4��(%-]����]g+V)�<-���b�{1/H�<0�*��Xn�gTd�y\r*����]�xUއ���:S;b���
��f�<��eI�u�0����S�����H��vɫR� ��c0��;�`���4�n��:khL��3����f�x��1�)N�.6u�]'8q#��=�������
�Qr�9��I���}zI�7e�B��$V�,ڲ�	Nk1�/vU��,�3/۸l�Ö��8k��sp�c����3-ji<V�pL5�sn1G��# �p=N���f�]̝�چp�WA��ͼ���Mp]%f�t&�{V#�^���H�N��(i��ج��w��CTJ1/T)�G�U�m�uj�ѩ"1�r����J���7<�p��H]Z�#u�u���U�\�u'g�����β2�eq�R�o�]G6��̀/e�q�޷���e �%̊�����oI�GY�Q�����}o��� �x�WGǻsLt*�+
k:�'P����K�-&����?��#d������lR����o�z!/WS]��2�Cf��JZ������ԗ��.�t��i����^�X�m�*�:�X!��\�C���k90؎�W9T//�.��h�8�{��>	�p&
�t�����v�#kI|E>sU��I�	��OP�AeQ勧+�#�b��J�k6nFAt0�֫	ָyN�<��`4�,Y�ty$�����t��T�b��a 騪K5��;N��0WFQ������J�0u)W�7w���x�W�Y8F�:,�5b��*�t_ �]O���S�9& :�ݞ�[���4WwgaX�]�[�2��;�c��[���^�}WWR'��U.�ؤ�3���3�a���56%�1#oZ�
Z��RK����h�,�.Qt������,a�ݤi���qa�W���8��^�a4�eɻ���q�(ҡ��7�x��JF��Z�p��=��VW\�buƦ����dG��F,YB	B)iZ"�p�CC���5�B�{y��kǂ(��'A�A���[��GdV���1�*.���b�S�mю��37�hC]V Y��H�i�V�J��Th�.���x�Sմ	�%����y}g�^�,�˄D�5�z�Go!�3[Q��m!G*g@�-d,��;i�ˑ�n�Z7���,+�0��Zw�=�ɃAA쫓�BCy`��丗V��j���t`%9Xfr1�R���pdbg"�[�%�<,rnL��CV�O+���$�U	�u�)ʄ
���ً���oC�\մ�y��-�i��y�ۮ+��ޣ�1'�����`�Wkh's7��lM�m%<��8�T��nX�1Z7	�F��V4`�ňe����A�M�gm��3�3F7d�8b})f,WP����X��ӌ^]�B�@5�U��t��V�e���;��8в��2㬹�3��ߋ��vt�EJW�f��(e��4�ғC�*�V�w�z���]q n��0��4��|}�ME���W������q�FXJ���6�!�fn�s�����̧��f��l����hW��ʗ�C�/3X-�T�G^uA~��6����r�}N�W;g3pe	�󱣂.�U���	��
��:��]}s����	��UPx'��엶}N�6p��e'@�@���-�Nt܆�yz���v��I�y��Fi݂�g*�k,�B�X�\�&���ir����WB�hM�[X� ��I��� 5>ngS�dP��N�x�V�1 )��+����2Dr�W74b�&�#A��y�|U�%Yy(��'݂��G�׾�3 ��6���0e���3�|�-o\��O9�Rڗ�p��Y�Q{��Ⱥ���E��V[6n-9�E�=
�t��痼h٩Aq=F��>��2"��#@A�كV`�{(]Xٴ)M�Wil�� Y�����u
rQw��S�R�8�O#�/Y`>����ob7��l�J댿�i��Y�s WXxڔ7Uc#�!�nˎ�-������o���rXosJ�Z�F�bl����b��I5���2�OTGH�+� eCj�Xe�n�^^���r�
��d�׵�ι�;�TP�[[Ө�8�u��waY�k����b�T6�^9���YGN�y0
t��`8��3l�Ǯ��Tj�;�f�/�K���a����q��
|�wf�8i�,zZ��݉��DS�u�����
�Z�R�zԂ�;�p�vTWb٦Q�ю�D���B�h|��M\�r�n��N�;X�C�S�ͫg( ��"R�7q�����E+I�gctɫ���wR+�;N����߁��YV��fuY���,ʜ��y�d/��[�RC/�h`�,w,M����P�)����Z�r+��"��֪�hd�Y�j��t6��Zȩ�͡t���˞	Od�v�4b���[�m
Qͭ��n�pOz��{ʝQqj���Yf�]m��l�V�]u+��4�4J|��Tt��:�����a@f�������^���������˗ob�nn.N�G7GkFƍ2hѣF�6�h�F�5�f͛F��1*�W���*�!�0�(Rd���EUAbn�!4ZF�i0)2�%� *���,�a�`�D�"|!�����DhQidB��cpF�m����
� �m�A(����(�B��J�K��$��G���n(E{�̆ck�j�\f8����r�.�t�<�t�9ْ2��»�:��v:�B�������@\�GO�u���ӚzY�����!�LMl��Iwۛ�Q!��9����l�N�qa�ۗ��T������kU����)����gi㲀Nѫw9�+JU��i
�fPO���T�(g�B��MW��O�z������,՘�8��Z��{��s1c킠͓_;]�f��o<�@��m�9=�{�X�ۈu���7M��V���з�t1qXb(s=Z��f�R�X�vk�D���\�J@h�+evQ؞st���1`�үD�YKAY�i2e��U�Tˢ$�o������stv=�zdą������rl��O.�A4#^�.a���{�Tӂ�R�Ϗ4@*v��g���Iے�a���<gndt���=��Wk�LU����gew1.=�S�z43x�
�g��������땵�����k��{3�/�rZ\H�om�nZF����g�E�H��3n���Xon�d@��^��#ne@�1}�9ۭR]֍L�,�8`��HB�^�y�H�ZsguN�1���W*DuL��Ǌ�S0�[Y�����WMVX��ʳ/�<UH�d�xj��6f�ae=�m�۔[m�i��)��M�u�Qr�DFM���M�t�"�A�LQ~$
h��<�M��^�2��(�I�i�	�ʠ��I�K@�ӣI��N�mI+���&%ҥM��F��I��.�6��@G��)�.���H�  �Zi�`x�TM/D'A�4��D�i�AI�4���	�N�m�A��4)�tP��4)1N��Z�R~ti�i�i~t�&���$KA �PTBi� ����H- 	x"�y#&�tJ��F�)�Hsnm�ۗ����I���<��D�t�6ö��K�����|��i+cQ�����4Rh��Y+N��О^Ej�E�El�t&�&���gITb*�-Y(Ӡ��\����4SN�tMV���U�cd�}�.Nf�K��X���+Mll@m�4߷9K�y����TV�T�9M�T����\�m�E&�mX(�ý�1-�>Z��4��F�Z>A��$���D�Қ�6ɉ �,i�l�@r䜚��jkm���MP�:�'KA�5�i�+��,Ese���g�d����EEQJ�W�����b���G61�Ph5BDTR��%DU�w�Q��'�<�'l��֨(%$����SLE�ê*���j�G+�����U��CAE�"���Tz��]����|�<��-�Ȁ§J�l0B.�HݛY�ź9[��y�˚#l-��G`�/Q4W��gt���v�%��7y��P�9�� ��̽��_Cb�U�N�=)���CA�(0i���AxA/H*j�(����C��VY�7�V�-PC�H��ҡ)��'��_��s��of/�V�����
!��o�p�H���9Զ�X;���p�q��|~�޺����m��X��7n�D����������I��o�ƀ���������vWc��h�=�������7�����6(e��lS�1������w�5�
�R[R��h޻z�3³�>�[�.Y�bܥ��b���"vB[�x�Ѻ\�-:Em6��W���Xn��?]6�S˕TDo:�4���_f�F=v_|;�/��'��;��Sԫ�'�`���m34����S�<QS�?��T��a��;�����ם�_ju �=/��F�A���/ޔ��\��O��g�y�[;��g`�mu��w<����[��"v���f��v��"o��3�F�5. ��:�:U��|;��͹7��6��Nn�FĎNN�u�����+%��][�8��;h�Wk��(�ZL�p�q�.L�u ���c-؋�9H�q��s��$��浛� ��hf��z���-^1��7����@a�{m�]��$�ݘh�](���s3Bm�n���oA���bq �u4u��64�3ם��^�����ebﱄl7@S#��Tpdk3]�>7������R�����������\nM|�a��L���Jn]�����C��U=a�:k�8���3o�w���w��i����>�����!IWr���bnI�b�m��-t���w]�oOw�_�Α��w3��l�ƧI%�sw��;��fƘ.z�d�L_�ۼ׉�g9�u!5}Q��Wv>O�c��l����}SO�^�n��;��a��x6�aڎuU^B}[��L릛�}}���2V퀲:��������������a�p�7�=��J�=���|����=ϕ���v��˸9&!����^t�5Ž]�Sk�6��C��h%o�a�>�W�Ŧ��5�e���8VFȬ�Ѯ��d<|V���Z����X�e�	� 䛳y����Jp�]_kp�c$|Š����Rk��I�ʝ��|Z��^�CSH�kտ��(d�P����"TV�qq��8���XU�5,p��.�c{i5��T��1�8v���-�l�{�Qi�A3	�4{��F釅�  _E��\�K�t��:#a�f���8�wU���a�?q�AP<o�j�\��t����;����`��#uor�z��W�3�x�P95TzU-��0%ܲ�Sv(,�E�l�R�9w����ƛ�t�)�y����^wB�xN�5�R��NS����E���k>�4
X�@�HQA�ꕼ��Ŧ;6n,��Yz�cg����|�t���6�+w��3
bHP���K�ut־�UI!D��Z_���� Xnضà��E�U��TN����;�og'{�d��;�+�a�����M������8�t3;��;V�2�.j`f<���M����-��G�&6��Y$O���s��ewԍ�f��o��h^��ӫn;@W]s�_|.�2w+jU_����ϩ�;��������ȯ+h�&� ��ӺT�S5oZ�Smv�B��� ����_P�E��bsy�fU,?�bؖJĞʸ�@�26sZHTk�V�����*���OP����]�hac���Ub�t����~���*�VRl�W]�M-7�C���x��4{�w�z�{n�z柧�j(C۪C���*��)$�;��<h�t��1���3y�Ou[��'�bCC*&{��3#T�K�{.�����2�p8=k�	��t�4��.;}E�j�}�"/'�M�HѰ4&U�G%oÂq�d��㐅aQ_%}ݰ��B����L��y�v����l��-����7$�p[�EOWW�
�5ך�[_[���U�f���X�̛�v�;�e�޾R��W
!�4%���U�·o5����O��X_OS����٧�;��4c��v6�i� r����]J-�o�k��8I�o���.�c�'xa��md	?C|T>��'F
���4��9]I��d:e`r�/�������b���F�.]ɳ��q�xo�����Ϡ�9�N����n��`5m}�N	ȧs�o9[8`TqyՂy������7$�gr�3��N�t���u�]v�:@
g�淚��³���b��"�"xj�4ب�Պl�_v���8�]bް�|;,�`�����R!���h�$�^0��x����n���[ٚ����+P�آ�9�n=����*��'wM:�З���Hj3�����S{k�8���s(Un��C�b�5]� '�>Ͼ����)N}�r�>�/�W~�W�Ш�����r��ѭ��������Be$;����Sr�� hu_p�S�݂�7�-�!�G���^=�k��a'���1Cu���Q�C���qW�Bə�K)u��u[G*l-��|:�>��_}�VmL`6���#�˟v�hD���2Ez��W�&8�}ל�W=���V�&#j!�6)��16�ՙ��O~��f눥�V.Ap��>�����E�d���K��n��ؚ?>�)���+�����Tov�B"ps�����-���gP�݋���u�X�̞'EF��+ �*��7���q�'^.����N.�W|���¾�*U�����ᰇ�>=������w�(��KO�$!Y<��]%�pT�J-�C-�&��j��ү$�6oS9�-�v[�9a�Zu��$���	n2	�2�(�&$���ˈ�X������,s��ŀV�N'y��ɕ܍����3$�P��z�D��;U���M���֚���2���m����L^$����}��]��V�9g����ҬuD���m��;;sM�$�6x	�_w`��)5`^�����ןOb\Rw;���[?E�L:�U���D᪠t� "�w�Qy��6{xw7�ֶb#"c�t�B�,�}��h��h������{����?oo�]�:U���b���]�>����r���F�h����ŀ����u4u��8�͍UR�v$J�-����M��9���V���dcV!�U�F��k�����0������qY��Zk2nO�M�l1?Rn� \��ϸ:�f��ܸ	]VKD����VW��/7;AD��'�M���#��Y1x������\o_'g�ᔂ[;��wJ��X/�,�ìggX�{�s�l�Nu������M>y&�č#u9J��݀�$�io�G��kn��lb���mR�+&Bn'�5޽X8)P�����^�޴��HP�E�U����6��ɜ�rv��r�Zs��;9��Kvw�r��f�h�8v3�J�+�Q��
Sff�[^�T���Ϟ_8�}7Q�;92�-7n&���4쿫
L�=ܫ���7çD�	lQ���t|�Q�y�w���R�*�'3��u�>�������r6��M3�\-ɳ�(�X�(G
}��m����������ݹ�7'��C����]Ƣ;�Mcerv��¸u�������|�a_qi|޻�6n�73�B�u�t��vq�c{�� Cl
@�U��}��_�Q�~c�>:_x�NP��&�m��&��w�(5�� ��L��jή9�'\봺
]��3���0�t�5�3aӨv$|�Ngy�J�%w�{]	]�b��p�"NY�+���[��e����p4��0��� �N�7�c�Q=��=��j@Mr�v:J8ڵ�;MX�b|~�B�9ⳡ}�3X�]�&v�d�N�
>kz	I�Ηz�e`Rhc/(h��|;�0*�7׹���ќ�6�tzM�<0j������v��B��F��p�#jS�Y�U��2�h4!\5���9B)b�Z�$WK|�i���eV�*�_-��=4�-�=v
}��6fn�� ᳵo�u�YF���m��;����q�P�#

�u���e�@3��`���U�� �3�o���A7�#]�G9۪��eV��j��tf��O�L��i����Xw��n�$з��ۼ�i�HG}������.5g�+��C��|]}VhI�JN=�w�`�p�����WnF\��5e�Av,A��C{s��=!\N�����s8�r�ڷ3��od�J��9�2����l�h��	�i�m܁sO�(�QB:�
�"�$��)���NP�Z햗����&���hA3 �܍�s>�`k,��jvMI/9:tSR�DLl x
��
ޏn�M �����|M6\k�a�+�rRI7H��P�-��8�!�a@E%}ݡK��9
�7��Q
R�:���ue.�w�$죟p��O��a�{]x�P[o~�.5��5v�bL�N��}	W̹6ՠ�h���jXJg��L�}ikǲ��}G�j����km`Y2�'NuW]�Af�.<���K1�v�����4��ղ��v�c��f�Xŕ��^U�ĩ�����;�9�LT�.7��N�`�Րf�i޼[v��u�cC6��R��ܝ�MNB�لu��z4ƚ0cS,b���2�]S"D�Ϡ[��۫:�8� �9��N�CH]��&'��I=ݧ h�v춿^P`v�u�+)�:�_Vp���|z�Mk�Y��v	L���;Rw�xl���� J�>�Y�zr�S�����-ֆ��7zF�X�ӽm��Õ˹�`u��X!^l�ݣ��y-�w����#�$�����׶>D�*�6(���G$����h'��ldL�K�i�!��"N,��צ ���؃"7r���tUi�J.X;{1���adu�H�؁��eF���
s���Wӭ��m�|I�<�;ا�U�����&��y�̥��:��M�:�>�����L%�|�lZ�+u���Q��;�b��b��%8n(ҁ	�e��X6�,�Y����om�o3V�W,��
(��r*�l��Oc�
�)P��Z��ԣ	�-�03���ˏ��ٕdJ�$z�F�ƨ�WY�BMIm4#���֦b^{(|
�rl�ׅ���+N�s+����s\Q������+9c&iJs����)H!��g\ɨh�^ա�5��Q��skhRĲ����K�3`֞��{wX��*���	E����h.�M<�W�'��"	|.���o���r�d�Rb+>�N���9W�O	I�Hb"p$�T�i����rb����Ӿ{
`������3�b���ӠoHZ����2	$l�z�5���ru�*��U�*��9����b�8+�>�{o�u��}|T�n��?]p�u�Ma����0�k�::)�����.�{�r��狫��Ml��`��"&vl��ʍ4�}�83�
M�e�ۭ�S��.���j�B��R���fᴳ[�3"��	.���ʭ�.��\pw7�4�v=㥂٤�>���;#���Ég@��)d��7v ���1wύt.L��*�����S��mhvlZ$�t&��8��Q57��)�bGOtǻT/_��tӶ�6�S#�Ѱ�t���?P`���w����x�x��ϯ��______������o_������_s��\�^Ϫ�C�J�|�ju�o[,LV�oQ`J��֠�E������j�,c�d�A��Ȫ�^��}���KZ����aVk,�.�ٺ�n� ��U��<a���n��cv_^e+F�n�i�'a��Dv�nTi^"k�rp����T/�]��A�T�JpU��뽰���?����p�/�f�ېeT~�^��R��l���q��-�@]��=��l�:�#XN�)M�}��M�a��_J�8
����	�+[�bI�	'�Ɲ1)5�裎��	��_q|j:#6���=���]79 �Z2�B�Vņ�&�����@`�ͽ�]ӺŽ���� ���m����9�,NQ��e�6lDΒ�a�4	;z6������a	�9�ڃ����t,9;%��wm�լ@<.�v�v��}���Ӂ�Qs�YE�iC0��j�P��g���Q�US��$���5�.��E
R�r����§WP��"�qi��v{q�NYўqُw)��CU�z��Q_��CaϜ۱����*.znm`��3o!V�v��SD�t�� �4*Q���|��S�s�M��H8µ����}��#�����p-cˏ^��j���J�����跐D�{pM.�mnt]!Ԗ�nV'�pќ٤��.r�#�r�c@�;h?�u�Lx��b@��G�6r�;.�Z����N�`od���9͝P�[7����P��Wp�¤��*�B��,��Y�J���]���$S�݈�o͞�O�Td0���6R�2����f�Q©,�8�u���ˤ(����I]P�g�X֔ٵ��O��.��69�H�xZ�M_qΙ�d�H����<N� ��B�ph��ke;�cp�Ԫ������1�L�L�Dd���@K�5:]��SK�Zy��EP�N�=c��W�W�m�����@�*kѳ6�u��`�8������({.ďM��I�)]L����Amcj͝R���y���R�B�������}���;����tF2��n]�e�[�;�0�Ëwr�fe!m�ELӡ�Ѣ��ȶ��8�=��f0J4��e�4��p��|�e�DX��;�H��6��$���A	,vf4�]
2\�q���&�T�,S�Ɍ����xoi:�d�4S2�TE�i�*��aT7:c� +i��Wk��7ۈ���͹]�)�Y�N��!Yb��u��C
f��ٳ{��%d�V�ݞ�}z���kum�<*�[�"��Swy�5��7P���mƫ�������<�2D$�Z?0
���+D�-\��X�	��l%h�#rȨ`�Y��Ց5�_�k�qh��5%�j��H(��l�^S�ǂ;���&�3��RCK�5ff�#��%9�n;����dB{.Q�2�����m�۔Sm�-��6�m��8Kۙ���|� �\���C�ܔ�X��8��a�y)�$)*�<��|ؘj9����ADE��llS��lU�D�lUUG�J�]͹�EU��550�t|�|�J*1�G�h(�b�4r5��T�r4{:
(��fJ�*�͓��';8�����"�3����I�Y��ȡ)��7,��)(��|��kX�4��X
71�h9/.DO-4�<�\/�כPLE�d������r���<*	��LIN�s��s�D���m����E��s�9���[g�c�:�1�����c������ڷ��ˮ\b��0Gft��r/�����I��k� #�~s~^s����>����ט#m�X-���/.p���m|�9�I�lh�:��[����.Y�Ob���UI��tr�3Û1�C[%lA�b0U�x����f�.���G�^[�ߛMx��78ьj	��bkm�-lK�ѭ��D��A����g\�f��X�N�^7�܋����^9�������Co�;5Kd�y�1�v��0��Jb���Y�6cp2d㵔]BZ���7��V�;�Ff�Jg���-�����}��}eקK���Pm��X�Gt�$@"x�v��;��p*ldK;{��W-�)�+��˼����R>���!�Z}l���ǵ�oP֑������,8�RC��p��ٴ��g�K^)�E��?{	�;�Ě}fj<:n&�b�ǃ�� e9�*���W�6�5%L�c�ʽjm�`�,���KR�޶!����+T��s�J�Q~.��R��ҟ��y�w)��J|�W%����OcoN��E�ż�[�Mc����v��O�[��P3���K��ul���a`�N�.��U32j�A��إ�u����+�5؈�|j�t�)�� ��
$�67���YY�.kWonN��Co/	�h�3���1%�|��t	`�&�~���"����݊^�(*9q�i��GU�ۍ?3&�3�f51�o�vK�S��0�;�����b����)R�,gu�!�Rko�Eݵ;�ͥ�$0���%��B=����"�w*y���R�'!7K�F-?,��,�;Wp�qI^A����t9z���&E�R�Fߞ�.G8�xe�C�f��9W5�0���������5I��Èy�#/�аؾ�R��ZF[��KW�T��a�Ӗ ��o�%�-*!n?m'�6�`�7��}�L�Ȭh8J^9*�;��1Q�I%��i�������YEؘ���Vp�������wj�q�1�L�Gvp�V�����]p_'��������~1!���0�����Pv Kr���{���OO�ʘ�U\� ��|F˳�Z��K�;z��9�ɾ��^e��Ϥ��F@�%9�S
z �M�ˉ��xb�w5����o��)eVO�:�Ʒ���z}]`�� �XO��;t����h~goh1]3��p�UR�����s[;[��o�$n*����		��
$@:�&#�A~�Pw�Q{���O����쫦����l�=���:�xD��V6��s}�A���aq�f��x�f-<k�~&�I�p"�ַjO��G���6ݼm"]�|C@ۇ�<C��t�Ψ��rB��w;"+V�b>��}sHv�{�AJ{�4���2����^���>���-C�A�W�M�K#iY��ng�z�6抢�OD7�-�O%<�1��'���|7�P�jFq��Y���ђ-�=zw�NI����M஬��S����������ʢ��wЅ����� A=z����c=�|j�T\9�p� �[z�6�e:���I�b��'��x�'��!�� [!�?>G�����b2%B��X��!������M����oC���i����ɤ�;�֖np�l;]�;F���$�F-��F%���z6�`ɑ[:Lv�s�>=�;z>�������w�4�9�9aѣ�9��SL��hλ����s��syv[wv[TM����ҼX�$��3�S�S8�/��/�2oLɛS~��%��l�U8��vww8А��
Y���E�F�p�����	�(p�%9��W*�qm�|�n��y���ǝ�3���S	����zq����!�(8v!��˷�ޗi wQ��	�Z��Aw�8�8{r���;���� u���� ����MP���~dr��}	�L9�v/H�zƝ���-m��d˴5q�W=Ċ�ޯKyv��2��Y��4�����zk�����\=�-y�0�R�Ȏ���R�]wIѲRjV40���{s�3<o�n8�"��H�r�v��f�wǿ8|m��}>2�ۗk-_���Ns<u�ax�u�y�T�P�^�����<�=��Dt�ʌs�&�R @�{qLv3�&bWnu��<W�����p\�d����4-X1'\qn���(%�ʣ�����h=k�5eA�u��U���+�����4G���t[L������,5��*�������4���k;�&�����x��;�q�<��V8�t�go ����������m�X�fI�{6]��$�sڠ{��˃a��&���l�1��n��w�ѥw�4��[��hՠサEc���������=߹]F�Ґ1�>�j��n�I,�&�/��td0Ͱ/����]+�
�fu�CJ�j�#*SW۳��6�M8sM��R����[�3�ki�atQ����o$�A|N�ګO�{��iX�����Y��\�����(>���~�@x�zA4���A�r2� �eC���K��d!_���:����i�x�����fV��h=F,O�j7��~*�!\�y��n���u���5-DL�q���|^[m������r���sLe�sߪ������ԣ�k��2�R%hJ��zޜoK/f��!�3�k��p�tS<��Y��`K&�q�1�K��R���D��`&DZ4)8�&@�I�j�0���tv�U��:w^�=EĴS�;@A@�q%�$3��CH�y��	L[�f��������ǋ��)�Cwt$�[�e��J�VB��R�(SCy6� ��#w�nuY3�i��]�5z�F���%�t9�D	,�|��r'����T۳�1�v��B`����ӞO*鵞\�IO�7�>�b��3vEM��aH7E2��P�@��,�^�=0�!��QS*�[i�h����&ژ�,dvo'qTqWK�ȴ��9n ��J����Z�/�;Ml-�[���S���Ƙ���RX���w�Up)dw:�
���o?�֋4�`��*\r�8%b�ҕ��@�5crvK��-54l�	8�0bn5Y�h"&����-]�����:ϲ�]M!0 ʱ��d�s�S��UE���˭C&V��n�"iM���"Ɍ�U��8^;�<�՜�%��}u�>
�Ǝmf��/D�ݝ&:�*H�B����#g���g�.=k�<6,�XepMc
'�k�C�s�$Taz��+z�>�9��&;2����.ñ%�BhxS.ö�g`����m�z3�*t[��V\�{���;�{����>#�} ��j�Y� /`xeX�3@( �8�&�*Ԟ�:��R�ѵ�u�sɱ��C�܎O�^=%��H�v�����ų�C���.�[�sY0ƢC�V��<���!��Ow}�<�3���>Q�=ƃ�ͬa>�C�$@"x�v+��ϳ���~,�;
?~�cυ�}��`�xVEŠ����b�~�{D��	�QILѠgIj�+(!@b�������Z�H����2���4�H�"2�@�4�&��a4�FS�S�罈�Ԕ�j�(2o;�jqnw�\[X����WX�E����0'
���?�hv2bi	��������)��ڊ����D��2����4�>�Ot@nhXeMBњM�(�0�z3���x/m��N�" 
�3���W5�sB�:a��W��d�j��≉d]#ȉJ�[�A���JS��A��̔�=={��>���]hKK�15��S�]���<�}�r�a��g��,���e@tE�LC�Y�k�}D�����a���l�/��72V�8gGU�=6�w*Y�j���^��;��mMd���Yׅj�t�v36U������開si�z'2�OI���K�ZD&
@�i�"}}'���:O��Jr��H�je��O�p齂mg@�n1бv�>����74��f0�1��v
Gd��0�;��m'�1I��)d�`)U{�������p���WEQ:���1եQ�1�㑓m	������aR�>9	�]�����J�U�I�s��u�\��@�`y��y�[W����aἥ[����8���g��[��
fW��w3I��&k���s�����������TY���!��;�'�"u�{^;դ*�\��Q*󻛺�,P���y�	>�
̛z�s����-ݛg�a�9�+����|d��*�N{=�q1(���/϶��]���*�ĖE�Yk����5@u�ד���;d�0`7	P�6��d��,gN�޽�ౝ"��ۛ������M���s4¼H�v�����6z i�u �K=G�FΥ����	�0G3��&{���H���>;��P&h�Q2�X�)�%A�FĵE��&c��#�%�@��n���P��<15���}��o?*̿�z��|o�}�-^0�,�t5�T��LVd�&�_p��FX6t.$�u0N��2����M<*c�Pwjq��ضؤ�� (i]]�W���rvmd`lF��U�)7�b3���b�Qa]0�-e��J���
7l�[�����EF�_^��n� ����k9�Ie��:����DK�wN��r���}���6��2���Zz�x5�N���� ��E��W>�7	�vx����]Ð��Xʌr(_A�EG���=�%;�'f��>�2�udW� r��f}�ܲ��+ɻ�{����c���F�!8���PO��2Y�l��c�P�5=�Ј]J�b�@�x�<x��DO8�bzD:��s&�� azs2װL�i:�F�.�z���/�q��������bm����ake���3Ĉ�2�,�@L$�;��	��M�o0�'��%9HȤ��86��4�+
�1=�\�\#�/Q�Ɗ�Ӎ�� c;$:�ϕ��{��#��&M�z�;�a�Gk��ӹ�9���h1�E���[�0�;�z�H܁AƟFzO��}�,���:���Cf_b���;����^�s��'�L��fqls� zk�����8{hA�א!�n��Qw/��ٚү	w��[�PJ�+�I�R�\��˔^�%%�r�vû4�|v���ӛX���S�pXЄ@�I�^S��4,ى8������<ʭ]k�O�vD�~����u6=rϤ�Pm��h���z���:��T�����-�)��	^��:vn�4#oh��#X.F�=w-�=ޜ�e��+{Vͮ@Ūp�H-)`�y���^;��pN' ^��ݣ�����B�h�4J++�q�,��=y&�u�:���p>���oU��d���0d��t�rɤ@1�ή�sl����N����~���(I�Tt|�|�6��ރ��o4{#�:&U�B��y��m�g�����7$���ڽ�����}��}�����̳�rwL�]��D�g2��5,Z�����g&;��`���̓�͗moJ�A�+:/���Qڑ>�^��֚���[�ϼe��������l��^]�g�Das�b��7�9>�q��s�^w{�<��T� fE�+��@��F �W�2}��~�����@g�
�S'�M<Z��7Uou(n(��H�ջo��U�my�4��H<5_A�T4r5���t���|oEj{�9!p�VK`�'~1<&�����"�v�ӣ2�g^UK[V�!s�A���+R�����F�DF_��z��u���-�0��g�#�pLa�s��d�f���M��
=g���'V?zFMx���.���i+�]����ᩭ��b�0��s�#�@e?c�.W�߲��Q�6<���ħ6��	�BJ�����5�z-��$8�L�|�1�b�k�3����7{mi����c�Y��^��,r.���¸e�[�W��C+m�.wF�8JH;�e;5���,�M'Ȑn/6�ڌ]^�zdЭ�fguE-���;ۡ��G<rnw49P֌C;��ݵ���2��K��u"�/�B������Cd�շ6���="g��P}��tC�fi�ȱ���^�1L�u�bYXuzY� ���_8k���5��� �67���/ȯM#��'nߌs�s��b���y�dQt��T��s�.[��<`���P��R�(:ͅUo�ƭ����ɦ�cv�B��=�I�UU��r-?2Nc~+�C�6)6�����S-��Ѕ;�د4g������"�kt<Y�%�W�˰^������ק"�d�7"f1�CM��u�@d���G�?�^�Z+��Q�^F��=c?G��-���MkxJV;�����=�3�K��-�L��gǩ�w'}���ۈX�`K��@�:�_N�E��-�=jCͨ�lvOܫ	,�ݺ��F�,m<u>_��N����,Ƽb�;���ǃ�����$��u��V���ث_-ץ�\ȼ������Y�� �='D[Iwb�<;��lA�J�-ي��o�x-`�E���O�ڌ�������6��4�A!� �M;H/��yINB�U���#�7�K71Z�.�^U4�,��ZP�-"�'�zǣ�ޡ�;�i�*�K�U�A���>���q
�,E�W5��
�k��j{hB��Eƞ����읤wqƥ�c����L�r�y��F�Q�x0�B��{n�]��.�t�qU��,XȒ6AȘ߻sR�o-�0�vm���^��Q�7pnD?�ӓḙ34��* �ϡ@P�%%14��h���?���?}��~}���l��Y6����Z�9hb�1������^��`$jJ���W6Vv���5-|'s9����!⬀���pIU���ɯ*2ȑma�E�Eǧ�Uc���v�=u���8#M��ؽ}BjJHe�{�ԫ)�p�0��c׭��վ;Ϥ ���V"��O�eP�C�y��KM��LO�]��d,m���"_Ƀ�bYHĲ2�%�f�)a0�8t�A�/�j쳳�7*67M��@t6���,�iO���<'I�9�Nl.�L��*Mmq�<�T�{]�WT�Җ����p弁@N-���,�^���}�.�H�;��O�b����`Fz~�f=Fn��;�nR�����r����[ ��"mLpm�/g���P��!0.͇+<�,{-�Rw�P϶�t�^���:���8�z���`X��o�y���4�ȡ���Mr��@��E�[K�o�'5�@ùC��8A�3�� K�GF�����2?s�;'��~DE�u��Pr3�gy�(	��Ry��-��pK������fX8��j����n�ؔ�����?���������������������>��=~>>=|XeM���@����Պ���f\+�x�<�c5]��uފ��1��y��N�EB������4kL��9Jn͌m��Ȭ�F�v�x*Yvmw�ۻ:W��P�2ut�	j�Ӷ �ێ�O{��r�`AP���Hޭ.�r��7v�V;`G�K��*&��'_\C+Nm��9��']��ֶ��CiҊ���lӲ�Z|��p��.mhL�Yǎ���x3쪪4=,d-l7+e�u<r��o��ܜR�b�r`컪؉1���]^%�&ˆ��DypM,�r+�p�ۮ��s����v�t�R�� T\tu��*��^�(�؆R0���DdQ��kv����º�cX!S-otf�ޥt�f��]����8uߞ&Y��R���0gM�(�g[�ysu�o#ˇK�ξ�j�: ۆ巍C�#/TN���V��Ӷ:�㔢ޔ:\���;�u�HW��[A+�s{��k���u�*�V{f�!wl�,U�[���A��׉���:��Kk][�Yt�pܠ��t7�X�'�o��D�۾�V�_�d�Ԫ&~-f�uK"0��ջWE���v��/%v��U��ay�ú�f�R�����=��	ٕպ�b������Hp�w�4�Ž��[&�h'��=��<�,����k+����!*1��;J�;b��i�qU��f]�\���)&r�8�̮�Ή]�4;*\�z��Ă��s=YF��fX�����N)��ڼ�N��27�":��!����j��u���u����k�+�bf��[�5\����68�&�gVe�9�YI͙��6�q�#�ok���.��׋[ٵ*ʖ��zs,m�V��9]0Z�vv�;&$wl�d��影[Ƶ<��^�F�%8_S�,�[7�Z]S4�df��VΧg"�emX�q����NL�hT��M�g9�3�`ZG$���z�3��Ѩ���t7e��6��\�Ӯ�'l6����S�1�T�m�@�1B�(�)�n*�M�`��	Ю���Ƞ�zŌ�����������)Z�[�2 ���V��ui�Uw�N�-1YW�*���[��=�R��p���K�[��n�����|l�͛uKnn�������֙��̼�vR�����vV"�)]�]�w�}b��5����7��{e^��6��������h-&���Į��W���x�}�K�l���a�%��,���&hˢ��dHw��5٦���dd��b���im͙�Dm�C"��Z��"ƹU[��f���N�I�Y��jһ#L�ũځ�"�ʻD����˰��T�ٙmV�ܫ�R�rV7�.�*�,�p����F1�o��4ACX*��#[�g�|�q�v��2�X2`_p�E�3f7��-jwP��!��vjXYS���2���KAV��U7�����mi-�M4ڶ�m��l���M�~�H��j��5�4U�+�bv ��j�Z4Q�F{q�"(��U`.O�~s��pc^`�I��ci#6"��3�5uc��v(61M6����h�5QF��".�����O"q.�7˕����1N,�|����n:�6"8�&ygZ��(�T�[�	#Fi�Bi�F.ss��ȏ7ͦ ��(�$Ǆj��#j��^s5qھl�btj$1�T��$Q�yj���q�����)�3�\���j���g���mE|��b���I���+��j�A�*j~�rt��TO�8PD�D�݈�y�q3m���Ey�5��p����*�e�M;�b(�����wy>X�Z�'q��7��V����Mb(��ST�~Yy�LU�-RR^s�*h���(#���nq9�[;X"��J*�
H���r��M�b&�N
"#G�g�衘h��������Q�l���%*���ADy�Ir�Q@TPPU%�x����y��~���qy��H�߅2�t���`���w��n�L�qfdj:�I䣶$5[�&,e�����9ٛ0�Z�8v�0'X��t�gg��d������Ur���tP,�D��i4Z%�H�	`�6�4�W��[i��4��P &���=�y��g��y����BΘ��ս��BDCdH(kh�*�T|�G
nu6Ia�^5��=�3:ĿXq���ޔ�:�@�[��X���x��IY4�}l/��7��I�!9�aD��:K�0N��jV9���Ճ��u�)e�$����2��(�V�����g[�
��_D����Vw^t�|d�aѽwr(�r�~L��o�����y���!��!�h[sO�a'W���s�zG���<�_A�˅?no��Eۢ�8{�i���S �ęv�[�i�sͼ>��3�#@{�d\����V��f2�o��^8��i��⅘A�梮PjH�3�uj��g��z�����2����X���3�⡡�ޘD\xv�TU�P�~k�'�U�����3��fL`+jz>�oY�@Ԇ���&��=k��2Έ�q��N����M@d�����s�����Ф��鄰���1)U0��YYz�5���c .����g���*Y�3H���N�7%ۄ��S�OЙ'�1)�z⫅�y�f6�Z�j�g��]��h�b7�Z§"�{����p�C)����׽.�W�����𨵾��u�m�E�$MT��ˇ��j\��ǹnwXF������7O�Ҝ��1ط�;y��ێ��0=���u�1w|��׿{��r����=�i�aM������+�2����ۦ�.�S)��`W솳��H>_\����������u�{�xx{������8r4�R���Z��g�`&Y~n�I��^���;�0�7  ��;��	�G8��V�Լ���k�ur܀IS�T��~&m�u�c�V���zk���3��p��<�Zg=^�g�6������5���/%��S��I�W�J疯�E��J@,yl�	��·!���g�gg��J���Zx,b��Srz��sBxв^��T��=�̪º�ݾ�-8�::K��zv�w����`:N3����l����LW��c�MͳB�s=���s?s�}	=�����l���L���N��n�^Oa�OG��y����9�&�k
�Ú�<��od���N�>�R�N���&}���we�j=��3�2%�=ś�7���s�8	�/b�T�E	5�f�Y����zu�ė�	�c�@��i:"��@���L���S{K>>��w�́5%P�Lq��9�;<��L�YJ�����Mo����C�* 2�'D[*޶�:��Z�G�eL�>Y�m����E�D�/b�/��cFd�/��z�W>J��O�Z=c��z�����lY����]KX�&Aڣ�.]l�H�썛�w)(�ɀBݒ�g�RV���7���X�MIWV�+m�ឡd�y׻�$<͓bX�AU���@�XムD����(�YӅ-LV$r�z���f�۝˯�6iλ���W��{��x�@��$ �Ͽ?���9���k�x�9�E3�"5�������Ȫ�`+�eT��jR=���ز�c�]�Q�;uy`�xW.�o��8k`x��}�6)���cH�0Za�s�|d�neÌ�������]a�O���/u�^�\.	ط8�pn���r&(\ש�:-��̘���
�>
����J{��ǎ���e�|Xטė�&Sx&�	*~��ǭ}Ǆ��|w�ý��H|�?�u+��^$�k
�ܝq�-�C�W��=�%:oc��K"����L��L+��|��`�xk� �&6o.Em��W�Rf*"�.z~�7�Y�3���]0�0����-���/�8�w��Уetd��'ϰ��4x���h�n�0t��B��4��P8����E��%�x���ֽWq=MvV���^��'��<c����8F�P���T��.Y����u�m�by�J''z
�x�����?�뀵�8�M.� 8�#Zs���M�n�LKb�L��M�ˆt1��i<�Z�೻�ck��ߒ�^����Ŏݸ�����;"Xu��t;�r��z|�;U�{*a��\H:���q���	�ʷd!S�*`8��]e"���4��6y_�u����(ju��I�#Μ���ӓ4�;К�&�:R�54��h�ɰ��J�[�tE�٦�Nte��7��f����ͽ���-���e�u��z2���m��A)hV�����F%�@)H�������w���~�~.�ñ,~�i1��:�,����1�z���[��gcn�����T4vD�ЦFb��V�G���"%9ǅ�w}��ٹ�G9&|��&�=��#�������[�Ǚ�h	���\������{aK��OM��{�H�A�l�l�	@>iW��v�7�&����]�g�W2�O�Qt6%�<�wy�Sq1��J�͜�O��\@���>�*6����\]��r�=��dM����{�����������~b�~�y�j� ~�*k��Y3P;3w+JSm�D$0��֦�&��Pz͜O�4�t�w���t?|mZ��^����k�3�T��GM�y���H�Jm&d�Z3I�J3��@�f=zޢ�K��硝��ɰy������Uם���k
B "�`�$�w��!�LK"���(JSW��Ưs�8	��qI]�����O��.�W� vg���$���%9O�bS��%� ����T���h���';e�38�E)d��k�Tc��[O��fژ��Gd�=�o������(�O��z}[۩78��,���&�q3�[ju��\H��
򤭤U9̣[М��䙜ӎ�8���Yw��M��C�R���{U���)V�!B��,t����ʻg����GDr��_>ŗ�r�u;Ո��MF^ǇWN4�K�Y����	�����+kB50�����=���S�
-
ҬH�4(
!O=�����߽��Q����/S��F�t�N�L'5����,P&0�dz=��G�9�hL�l��5�*]�9�CoT7Uڥʛ{y�u�1i��G����;��a ��a��8�!����L"�(e�sMa9�����<�}����3�H�K�,��e����2�q��ݵ�v���-���A��G@{ۺ�J�gn�R~BvE1��mv;�'�֙6�`+�A̰qV���+@�7N�y�V�y"�ϴv
��~B�zQ�9���}
Nf�j�Ia�^5�����WX5޶e�w
N�ez݀[5ݪTz�b��Ҽ��`mg��s&����K�|��A���I?���i�x� ��,/�B���!�'۱�{-X��ޒҋX�q(ɀ�Z�"�o&-�&9���X�����tV;��ٸu5Q�\��ռ�f[���L	:"���o�D����t\sH���tŶӖ���#��63b2V� ��z��
Zk�	��n ��A�r2�m�I�m��ȧx	oHA�)ns\tY{�~^��Ӹ��k�e�(ΟͿ��x`��m�A�������g���M���΋�	������ O��n7�B���'wmLm��i"]����lN�E
K!��To��5N���co��IW�Em��$�3W�(2`4�Cdqܽ�����۟]l��"h�ޭG���bqHkѥJ��ʨ6X;�osu�"/��T�u�7��4��r�Y���7�=�РңB�P�Ĉ�*4�2�L**L	?<�����MJ��O������"�jܨ�e����xa�j�,�$k��|`ɽ�*���.^d���ώ�&�θf^C�<�X#}j\�N�8βj0��t7�Z��b��FD��>������*#�gosWd����
<R� c�ڟg�h�ߢB�����0����v�"�Ss7:oc*�"zz$`�Wb�!u����r�����U$��:q�c�N7�A�g`.<C��Y���j	T��(/og�de����*�,���[t�OIC<s�kK�A�mᄎ�"1�C����m���+�Z�ӈ��:���>�.;W\���~&m�u�`sJ��@��=~g�8{`/�Z2"j�Z]���o���P�kץ乮�B��4�U��9P��
J�[.�Bxw��d��w=WjUއo&.����g��^�����f��q��QaK:y�_����Y��{o���l�]���{p�G��tX�`��� �cB`kd���������p�ڸ�1uu�_�7`��/ٲ�������4L�t Hb����8��9�1~wQ#r�xk�oG���*ȕ}WF���<���2R�����ө�:������L2��*�DI�a��tڙ�/��^p�n��բM���p��업�)�E+m��������/�㾀>笅[�E�]{������ҧ�.�hW�խ�d=i�s�����9��� 	���R�ZZX�~|����w���_�6x=�Vg��Q�;���u|���HC̙����i��c}B�`�Rڃ��~L�^��.�{_)0�	����a���&e�A�ǜS ��^]�	oVM�!,k?VT�v^'m���ʑO/M�z]�ȴ�C�A!�p�r�v �����,[ڣ�-?D���;9������#a{�T�Χ�U�my��#25������F���y8	�!�*�n�.��̦��������x!0�a�	w4^�TcW_��Zچ��A�� ɽyv�+����y963Vtg����5{�
u��+D�]��~��`yM~�8�|/��L�k{��ID����s}�������0�L�ѡI�J9B�Fc�=[�O�흀�1m '_*_�ꍒ��t����X{���{"L�dD&<�%9����j��}���}ǅ���<;�����0�1r/��Vv�[v����O�����|k��2��xd]&�I)L8?E��S�0��mK��e*�sYZ���a���6�D^��h�Ƒ
��y�o@]0�0���-�yoT77������6���@�Qe��`�Lf�؉����c}�;� oG64�>�Y��5f3Qjꑍ�+��B�b>���"i�H�K��u=:-�e�9cX����O&qLc��6X��s5�F�Xjj����CVE��KR�֊*Kˍ��@?ԀR+2�R�B1
%J�0�D"�1 �H��~w�o�>���n���TX���!�63��&����I�«�����K�2j]u��N�x��m��+���)�|j��@�y����Z}#[�L%�L�;B��YkE�jl�K�s��'��~��oR��o�s�09�ס�87"|�%�!�G�2��W���Ok�U�%�7�1�Һ���s-t���r�9���6�E�~�t����MO�z�4�}v����k#�z�vf�t6���)�OO�	�N�/;=r�h���}��ьPv|��Qѕg7n�_>����y/��]����C�nFx����^��1^�v<�lXM;cS?��}�E1�U�}������xu\�|D���3e�j3], ��c�8�;���H�Cx��,Hc�W^[��n��N�S��g�*]fĳ�� 饥�>xkd�>yZgx��(H��T}Zn�g>�N{�~
U��a�z��~��|;���X5YM��zxk������҂����,�܏Ip*{f�Grz�+_+VE�vykWq�mXeT-M�L$r��l�z�o
�E;����~oo�HDoE�*���d�@𣻻�HUZu��>�P�֮��T��26&�#�p�3�w��}U[
����D��ƶ���L�ҕ����Za�z�ޑ4�d;P���a�t�Bh=�ek5��I�wR	rfu3C���-�m���,��*�=����D�����Fd
�h �fY�R�")(�Ef(x  � 3y��姷:iV+
o'5���4��hq�����^��L�O~tX%cj+��Bl�eMV��I�Q�a������7�a_�@FPE��/�Q���D�xa>�&A���; ��d����1,��	�W(�[�����`W��F�vv)�n�t-g/͎�1Š�	�f�r�gcH"E��z~�N��x[�'�F�Ɖi����$���8�:<)ױ��>y�ฦ�BR͵1��d;�����g��`����Hf���)Z\�Go��C�dQ���d^��#ϲ-� �y�p7��@y�{<�]�����D�$����Nʔsz�Qi�g�H%�.O#��%�x����q��~l���MhӲ�$�{K^���(�>�0�1����v�/-����^�Q��cHw�s0����Ra���e�G�M>!ס��*��ꀞ�
n��mvt���ӷ�G�+�@5R2�-ݛwV��P}n1T�I�=��'�>7�S�;)�_0n��a�^/����N�pҴf�_�8��#|�?]��>Ud�!LY�[���>w�nP}�;i'�x�jo�y��v��
y�q�h}�zZ/d�J�f��9�SL�ݬ��"�R�5�ӷt2��<�����κ����j�ܫ�@ی��笿U}�jlr|�;;�EY_ř�Ϲd�q�K�pZt�L	��QR�I���F��0��L��{e�����ʘ�Y��E?�!�eB�Q) �P�dB�Z@�A�E�(� (J<�����Y����حjO�5��s�<���D��;05��^��2V�Z���}���!S\�3�8�wC�|�m�׶D��!��.9�'T��w��E<d��޽$k��DT�h%>�Yq��<�^*m�nEza�c�e��6�kdS���w�h�Ԧ�-e�����s��zw3k.�qE�mb
�A�1l����T2���n�����q5w����;�*N��y��M�S9젎mEcr~	��a�դY�P�{
�c=q�#K���Š�������+��;@B`[z�A���iQ�����ntc��6r�yU5�n^��'�N����{'�Pp�.1�����A�p�;`ܗn})��fq�ѩ�S���x��tħ64-X�S�C�[��N7��i �؆Y��Ko�$Ut��-ߝ��3`e��q���,`&*�t�N����3����o$n@���uvz
��	U���Ձ�0U@A<�����N�;*JzoY1l��c�B��6��zw�~} g�����{=�>^�w���������������׏���_��^?���o/���k��t��u��MAl�Z�:�ڻ�v��z������˴��t�U��]�%�^c&�8��8z��+klӥE��+
@n���G����z��넺�����m�;��!Gt��]sq��e�K�Mw<;��{�_�L�6�.�U�"	�3rB�F��%f�fIwvD4�U&��B��������fV}�|g��]��޸���B�t�T�̔o2+�U���en#�m
�M�W+����O�YƎ��4���h�x�J�P�����2��L+��&���٬�Vm�\�7%�TMܤh�/�B���Ӷ���1��9N�e�l�p�ΰz�*!z2����0M]}�]r���9�r�� �l�9��Lm�d�M��,6�W"++7X@��˾+�CJ/�v;������0��]�xol���kVٚNY׽тl�.����R���E���{������6h\�@��F����3�=D��f񥖙�zz�&��]tID��b�ۧ�{j⏱�ft7V��lI{��v�(vb �scn��qn� 巰���:M�F;ssnd��r]�e��@�&�:u�
�n�"��4D���A�:���6�-�5[r�!kvti^��ȑw��*7LB�3cG+}�l���D�[yɝ4����{���c
�εC��w59J��`���B���Ku̦54�I��sX����'���@�i�ݙ3F�@�Ժ����Y�o���àxi��N�Es��<33R�Z�ú+ɽ�
���X̓�"n��i�S��n'�ƹ�9���͈���&c�v�s��zCZ^c�4W+))$�lܼJY�y�V
$*vmQ)`{�FN��X$�C��^3[-���Z__P����c�l �SwWF�
���%ê�t,��F���ZԆ��S-#h�Vоٖ"����t���� �mȲC\I�}Re�U2���(��laW���L�{[��zL��v��9��],�I,�G*Y�ő�lv7���n,�ڂ5�V�(5����+�ȱVC_�����FΪ�6;A��8+��an�x#���x_<pޔ�O��v����Y"����e^�{�PL�a������tnK#�u���H*�F>5*`⃡��o��R��lR�oqaf$�N���ZR"��n�i��G&<�l�7|V���׹6�wdڊ��V�J��w��'[�F�O$����R�R놺^�\a��n�`WDj��� �����eX�8�-Q�(�J���ۉ:I��9���؁/EZ�Vm#�������
�����{��n_1N�^�P�������|��os��q��n'i����/��4m9�XӢ!	�Ylb]nٲ��w��q�N�KX��\���#4��]�L���ڥ�6�wwv�wwv�t
�� A �AD4EA1DM������
)�(��$������!�b9i�*��MEUD���fIg�W݉��9:K�1RDEEED\��i֪�
j��&�&�������5�������&"Jj*�h�؂ngTDU$��i��*j�Z���"��~lTTQ-5EDTTEEARAMQK�SUT�UP���TE_�1DT}�Z"�G�>�S��E3��$����f*�
&���(��[cQ��LEMܴg�$��2LCDUMQ7�k�1QE3EE��4�EE��K,�PSQQCPQDDTSRU��4�T�APLT�EPS�h"�(�����7ͨ�����(&"�
�&�"���b�(���$��PS1$�TCDQ0� w��Ƽ�����_i���o�䍙M�袧lgT"��l��Yk����3U�yiqaV�y%�/q�O�}������|���_���F�B� V�R�
P!i ��)F�B�e�( =�oo  �Y=�6V3fd��qiݐm/��_���dQ�a�¨��,r��	Ib�{e�Bӏʠ�EOm��۾�4�rZ����̚��#�gB>j
l��.�TXRΞe];��T[ҥ�8��V$)ÏS�b���_��8E�G1����8O�s*F��a�j��N��TCmV ���n'{;��a�Ol�� 8�R�迪�x��'��(I��u�q�B�{��v_���q�r�se�exO�Z�	�i��5-�yŗ����ȗx��`<h��F.n,�; ���߳VC{
����"K�
��4h��bK�&��w�P�xF1�`[?<��������63޸�2�.��V�LBe�K�l6*1��7��a2,�w@$?� �#.���t���tI��i�ŗ�m�O_Z���_�*hE�fJOb�/��lcNd����r{��=�k,�6h����ڼ�#����C�9��!0���w4^�T�n�2
��yϝۣ;���}M�:�v]\�?|N�����"p'f�6�)�{b��M�8&O��s�|d��������|u�h~J#�UŲ��h�Ú>��Z�]��fNF�r�~�hma�X;2�K�l%��ey��/\%�������z�AUU|�����m`"[����=��\��|���K$Q+y��Ob�Y�m�J����»2���?}��������~�s�؇�J�(P)H�D �H��
��K!@ L�)Jϟ?��w�o��ykS����)	�Z4)=�9B���cռ4��;G�7�f�'�5i.���ˋ�.��$�u�r�oW�k����%1��%9���	�T-�.�<5���	�[㼨�g��8�c4�y���YS����,ǟ����5��):��%�u�n�)�$�0nz�;J圅W8�g���6�E�D�0R͔"�R�18ўiZ3��W� ��,�0���X��N�<�,��������{���_�y�6�zhfƟ�	�&��a�
7���T��0�έQ�����v2}�e4�F���^݄Ɨ/SC�Rq.���C�C&a��Lp�n�1%�L�Ҽ;e�R<K�E.�sB�'���x�s��X|���#��\p���y�C�0c�ܲ�FJzN�5?N�f푱���|W�+��ߣ��݅ OJװ��k��+�i�b:��;"Xt&~>.��~5�w��-�;[�L;1���d���)�'���cя�&9�T3,3�o��e�]F/���b�f��"�<#��"u��]���Hv�ܔ_��zKy�D�LJ��>>�R��|a�#�r�ffZ���\{ic[��,+�c�-����1�_�w��R⩭�>�Z�$+'#d�м�����Z�oI�鸢�ⱄ.R�L���^�zw�:����n�f��QhTQ��J)M�٘J(8ְ�����EtZ�![��ʜ0����JU
Q��f
Q�D���I�E���1/%�f��!�i�.�h�WtՇu$v���1c��H���_�eh|.$D�����t��df�0���$9�pl6{Uڜ��[����!�V�;Iz8c���g� �xBKI�{d��r�5����D*~�p��Yi;t[f�4!fSA+��(.�Y�P|^��9���Q��9<=�A�¡­��՗
�;�E���\b�	�U3k^A�Sl$nC�������ȕ�%��7�æZuF�I:|�Υk#ϦL��S��^�W����L ŕ�4��������o������;g�Yg�s�!�:G� DA��v[�Ed��nt�^s���+��0X3a򡰑��m�y�IK�J�?��gKd��Z�H��Zaq���3��<��'��Jr�0��j�`�٫�}=}:�mVM&�������y\�U|��_�06S]C��f>���H�\k�[N�]N����5�W<�g�\����V�X�"�-�Ú�1��>G�e��BG�Ȅ�mLpm��k��P穢*ժ��]ة����HY���N��?"�A/K����3L$��4�Z�x{�������͇+ �/�t��߰AvZdf����.����@�>�N�੽�A�XdB�W&�jP^S&���׸0��m� :<�9-����r�:�[�N��v���Z���]兖�"�oTԆY�a
B�B�v�ڛ��l�5￿�>\�ny����ݾ{����V� �F��B�)P$��biQ��i��Ϟ�;�{���b�N>����=�s�s]��^V@�2��w=X�8�a��Ƴ��b�b�L��Z����)��wfN15�E�c~Mc]�g��Z�&ެ+�@�F7�3h�4�}�n�̘�m�e^��@���AC���|���L;k��ͯ���B�0Ɖ,:�Ʋײz}� �KSC���.7�9�p>�,�>})?"�dP���E��]{���}A�^�.�ճ�H�x��y��cܱ�D16'����XM%Q�oIͪ���l�H�Jxp`�(�Uy�Fuq�'�D"f4]�U��0)�}����m����FZm8�^��^ךּ�;�Hw��o�>���s�mΘ�{)H�����6�5E���gC�g��+�Z�n��3����j����-�=ŷ'�Us�C6m��$U�A���Pd�[>�f�2����$����׳N��]'�x# d��y=���"�%�QW�{�Br�����@�Zl�p̡�;���]q�]k΅ďnF5���}�ւ�sb$��x�m
1�vL.v�A�8�����?k<�'��>����Y�c�O��]���]*Ѣ<�w���J����b&©ɏ+11�j�v��t�������m�_n��Y%�P�*Ɋ�0�{,��]��2nqU���$���j�5�Pgrjd��X�n
L�4w�䎰n����aҴFiv���C�JA 4)M-(R�R�R#@J��y�������^sO8\\�4���X(�aM^��ơ����9oP
�\:Nٹ.�6����͎�X�v��A�n��|uNm#B�ʤ�]�N0�9{gf�Ӎ�cO��(e4�����jý����6#��CK�v��4�`c1V�Rz	@؃'��ٱr%t�&+����,Uͬ�=���YD�,'�p�}�d	cWƝ�ݕ%=X&m�u��w��V���zk�72=o@Ȅ��t��uK�u��C�b<C�=K�~�uo&@�yj ��/V��9}�2,��wy��MvnZv����1�NX���"7�y�T'�7�q��%Qaq���-�/b����V�K.�	=��W���Ƹ`�D�v J�:}@�
ׄ�E�וMIf>v�4^�df���N8(~������\�`�s�eۡC�D�
�X�'���W�F��`q��"I��-bVl�C�y�<i���X��~�ײa�v�5-�5�0�x��s>2%�85�/�4���7��wq؈��gx/Ja�k���f��nQa@���L3z̻O��� ׺���~U�T��m��T�����{�\Xvffٲؖ�*m,�Z��0w�wh�y�inZ�=����uN�+Tf��{�ꙡѻ�z�&6��9ȵwtr�A{�@Ӕ��G's�or��Q^1jƬ�3u��TO(۾���I�L��C~Կ�\�DY����}��I�
T�Y�"

 0�D�/���j��r-�~�ݣ�_�nq���f�e����@A���l�V�,�x�Ә��XH[�����e �DH:����H�&��љZg`���rC�V�}0�r�V���qޞ�or�4�m�5t�ê���Xt�=���`�u�1c}ve
"v�l}������܆k�0�*�t)ZTu��ޜap��X9����5�~F�vu���ܾF:�:�6�L�c/:"Sm�!2�hФ��ȭ�u��=��y�)3v/7\;�X������0���"��5?!)�/	�Q�(IP���ǭ}Ǆ����n�wu��{�<���tC�	�Ex�GM�W���):�t�tS*�J��^[7��B�ˇ��u�\�Tn��g
�r_
��yߗ�:{�:��k��EL-�]Z��]u- ��1+4nBάE�F����;�ׇzh(f�~����7w�M
o�N�$=���FwV�4��ܶ]Y�OE�r�t(}d)�j��>�B���u-����~�Q��U=2��"6b
��Nj���u�o`7�e��g��ݏ�����թ���$����ssn0����'�F���I���yZqw�,JV���#�E#�k�eDXrn���^jTeظ(B�'=�Mōf�Dͺj���P��<�_�<�{�@���B���H�iD�Dh�JTbPf@��������t��^nV;��s]�����C����d��F^�Y�iU��v���8���ȑ�g�� :��>f��uǗ��<8p[o(LKq��֛`��%б����{W��j9��Ցl�t�kC�f�kVKUFb���<)DE��;-"�m���W�1�y<u>�}&9���1�[�&���WT��j��҂��F��:F�����8�[�Ӡ���~�5O6���PhC�ܕTwˣJ�&�h��o���Dck*�Ļ�XF���G�T�{Q��19�N�sjGB��vi�l�F�(a��1>����1}(l�*���xg�Y��KJ���z�u�Sٍ{�3��L��[�sgW!��q�h��Ê�.R\7�i�y�V<�43�Ɩ����7��.�
�|�w���߬�9@UMy�s��m v0��ٻ7e5jo|�5�%��7�9���W�|)��uܛ���k����{y���}P���8^b��jUc�^}�w)��L�ɞњO��z3lf��!�.O8�xa��%^<^.]�N2=�%�`����d���C� �P&%�t�K&��y��7�,[3�'��p���f�D�s�sb+;���[]���`���^����%���31�x��=A��l�"Ś� l�J"���-��3�#z�;�Cr��Dk����ݺ����!5ہ�N\ oP=���[u;:���8���O�	J��PRR-(ħ��~�v�M]�\ޕ,~o�C���ȧ�x�%D�f�	�̧��#:O=�P�ɁQ�B�C��PkKv�m�r���Ȧ4����������\[P���k�O�d��]�>,Y�Y�vr�p�V�'��)9X�R��n�3�__#ϡ���	���Bm����s�<ՙ��]�6����SR{Ο������.�O�(���(Ey�z������c�����C�����3���xb^��i����������I��·�c8�1.�zh�,�7�ɝ��	��$2����s��:�:-��wU��BO�V�6�j���"tcm�e�����jХqn��;����;k��ͯ��hZ�bK,����[Rh��޺�nӼ�({v�q�({rR�QD�1NC�VX��!^�#�%r��;���,�vp�К~�!�tK�D������׶��� s�<h�gh�L4��k��2��&;Sљ����sEPt��hA1%�I�b�\����h�/~��x5�%�<q������L׺&�-[����M�Y��gf�3�F-8����E-�]�[����MA�EB���M��&FjhP[��Ւ�j��aֱ�ѓs��.���N�iơ-���ue��Q�̃QY��Qd�Ha�9+��ro*fh.�"�T��;_H��&����IO��~Q���Ohyfϓ��'{`n��W��d�v�-��?4S��0��Ѥ��k�;҅���@������S�Uϫ�ٵ�>�	]��U�I�rsiQR�I[���
��,�����@�S���zap	�y�ѪOׂͅv��On�9!�'��I�g�B������{lʋ�Up��I|mq1%�G+p���Ϭ�f��fٜ9�Q�M߹�����ۮ��}6�,b4)B��[T{����2U�3Ĉ-�
����P	�j��c	����;�Curv���Ũ:��=��Nl$iy��U$��:q�c�BΜo@�c"6�_c�q9��7��;~6${�S��P����v@R��p[�n��2z	@���zP�;5����<&վ�[&-g�x1a�����5�G<�@�U��N�;*Jz�f�XAa �.O#��ƳC5��z�ɨ��FTG��I�@�$TYZEL��A����?WQ�G�n��]A�[���ڑ��q7]vub���N�|^��痥� p����	��/:��f��8��@?�����N֞­���
�f<�ze��!w�e��&7�=�E¶�D"{�tü˘�.�Ho�WGMC2�N������E'u����jO;�Y-��w٬ܺ���6�9�1���!�t�۹o�o���4{��0��3M^pz�7�78�Ve�l	���{��o ��M^#E,���q˘}��2���(ӻ*�v���<%���@��Ŭ@Q�j`cc��ǖi�z�6���?vZ���\u��J׿%���Ts�Z�tL�t 1?DW�8��o]���u�`�q��;nKe�Ua?Mk߉�i� ���@��3�D�A����TaIm��;r��� ��E0��6���fE�l;n�����^��v��=8���>[ꃇ++)mmCY�����e���y/�+�%��28;��FdYx��	E@A��k�-�f�Y��I�
�ƺ&�P�ρ@�B,��̔����^�s ���6-��J|l<��p�Ϋ�pwB�$p�k�7n��b��<����z�璁Jwj��ˋ��9�<W��v}���C/�ct��ބU��JҢ��^ӌ&� �s[�M�83�%��G�~����na�������ӳ0�����~%z�2�F�'�J9B��׏Pȋxjkgb��j�Tܘ{��^�<��M	�ǁ�nV]F�׈mT�bD&<�����	�T.�g1������|��>�/G����{����������������ǯǮ[�?;y��!�¢�V0XʚU囵�/�9��opS8��(���m��.�e��V��E�r<Ǡuk����+t%������죪���r�q��C�.�-��p��ZN!�q��L� �y�3�(R(��s�H�B-˂���4tc�����Q���Χ6ynw�RΰU%]�ǽ��m8���]+r�k��+��YT���V�5wIu�$v�ꁹs@�8Ĩ������)��Q�f���v.Ԙ{ƑSCsJ��&�î�yj���|kpʈ,O�#M��p�UJyzbq�n;,-!+��oed��gG��W@���t��6"�©s�shM���-Ѥ3 �T��V��v�����E;r.�M�J����[*�M����n�	e�ͩ�J�W]��7�@�^*D� �87y&��]�:UXr�H�gz:��-��&&#`�j�q�;�7�����n�8�1N�H-S�k�s,J	��ui1�V��s�j��\2k���O���ٿ8;�]����l��)V����"o��:�b���{R��|q���]�a�3�><��F�8W
�t�zA���6������ܧY�{7P;ˑ�5gw��N�¡73m�H��}�6{nP���q��.��s�t�4�ϓ��c��r�wo�U̹P��tQ���)p(���9�Y�ûɧy��[�hz���u�];*H7W&�k�kI�rs�Ւ�5�d\3(W[����=��)3]�}]�]�˭��p@��/N�"��4;ߓb�W�US���dJ�A�V�k��ȧs%{�P}BR��P��w>����4���W՛St��ux	c��!ט��]�y��t�-%�t
�_�D��
Z�p���r�rT�;�.���.�ܖ��3��#�QL餂������U�
Ҟ�5WI�Gv+4�H5��ʷc��LT�G�#]xӺ*���bN��ԧfi�B�K��p1�QF�ՈJ�P3D�"΁����zs7+���*W��Բ���Vʸ5���d�˾�0���r룵z���C};1���ة�K��Q�݃�Z�
JWt���=�eOk�`���۸&�����(�:MyY�BW^�f�E_��ǜ� ���;W������%P�o+ ڱrd��ݗ�NJ����"�XE����T�h�]sfr�H�2P��P��	�{8�0��o1eY��;�7ͬ��mҳ+Bj^�+ҲI�opJ�n��6����� ѩ�n�^�vpn3��ɖo+�E9�y+;�M�g/g7B��ZĦ����1&d7N�w91�BMu���1b�&�u=S"g7��a;������K��dMTɝ�3o/i��`aSa����2<9|j�e��wxh�2v�F�ެ���a�HoE��߀ �}}|��hf�B0��D)�.��MWs�u��	�;��11!8�БD��XӖq�S���v�km�M6���w)LM]���A��1ET�Q4��5MSMEEO-Q'3����d�h�������1�h���Y��#�gA%%REUQMEUUDD�L�_-E5Ash<Ʀ��P�T�TD܍EUPDUQQ$LQ���`�[��*(hh���&"
�* �lU^\��W��E�����((&��j&��41�Υ��6�����"�)�j!�`�i���gY�J*��,S͊	�b�*��4晠��d�����(���	����/�*�F���֨���֪"��)����*
����/,��T$UALy����&����+�*���0�"**��I(fb�&���DS4M���$�"&j���&�b"j�">�J�j�"(��O�z|9�(Q� $2�@����Y i*a3\z�e����-��b�y�[Q�K�)���U:��tT���H��Wr
��G���c�ɂ4�veh�+�K�h�B�EG�S�)��0�@�)��d2ˤ���$�A!L�F�N�$? W����z����8፱=��ӵ�T�&*�V����;ć�_�|��B~�pEq�p�I� �%�u�%9�Ş��qs~�l�\3�G��[\f�ι�Ϳ�~���:����]�ݑE�
�3���ʙQ�;��۝���tSq�0��4�9���m\3c?M�0t��B�K+����]�Fr�����׭uu��d�ܔ4�TK��.e��|��QS�����&��5D��k���p����8�������sW�t;��Y�ϝ�=�BG��7����L{�~i����8{N�	�d�e51��0'�c���T��\sH7r͵�l���J�L��>Ze��CA����D;s�O�;6�����؎T��	��ɟN�x��s5ۂ��>�J���a���腓�&��A@x�����c���>��އ��e�O�Ӳ~�6����W/
S��sB�W	�M`؇e>1.�����ĩ��6�5��h1�PjG��W���n�g����e�J��&����N�T?PȖxBKHC ���N���ee�x���F�qi�Iv>ӓ&ByQB�=�F���{�ӱ��󪮅�vٞ�8������F��[�0��w|`vʉ]wΊ;R��1�x�GW$��zep��G��l�g�g!{`�i����ٝ���WY���v���7j���Q��2#�﮶ճ��S?��g�J����������Ê�h�%�=�g������M�֊qq-�~�t�G}��n(�AwG�9=v}NN��^�\AD�hZ�`������F=W�%yL#T�<e*�ׯ��V���;�5�6머��k%cj+��Bl�L�ɨFi=�Fq��L��5��v5[�Χ]z��z��8���1 ��d^�U���'�2�˻�˅?a�gb��Ş�u-��̍Y�f�)c	SGH$4J��}jT��G�fW;e��B*b�l�{b�yC_o)��t�%9\ށ,�%Q���S�^|��T:<�i��mLpd-��zo���V�LKY8]^`����٩�Uԓ�yNR�)-�Û��9�DG�d4[A�Fʦ��T��Ĝ���=>�
X��O���'�*]��&�uE�`O�)�*GW��a'�?s�;����M���Ƀ�pr*;!����OD����s]���Ad�c/A(�ze�������Gzd�_���v}N������ʿ�U�wؤ~+�M���\��=�	��Ů�6A������Af���zC�������vvu��*���Us 7p�th���{a&�w"�H�0��X��H}���u�C��l�m×�KȪha�5:v�\���v��.�Yۂ�+�Ϗ �GV\Nd�o_+���q�v���dH�n�EI](��������rc7�	��f�S�����d��s�ML)�N�Rm����}�3Z����×u����E�=>���b�zr���p�.������Vy�N0����,�;��۸��H�6���D�LW1n����� s�>��v�`PYS]U8�����i��if=����͐����@���D�1i`��DYz�m�׶D����8=����<���x!L�EG4��=1m����n�P��t�v*)�m��iZ��EB�l��1{��;��|�^)1槆�\JL0=Ų/uW>���X�1BAŗA��y�A��r,����.7[.j��Ým�]k�"ج�l��=;Ń'$�!��o��(~ڊ���Oͧ�3��|�yk�PNӵ�9�7�\/���\d���sN��(6"K��&'��j�d��Ű��l����[����t�k״���G=B��*L)�;'�@����X.5�$G���Ơ�ˮ��\����%�om4�췥�	�[���I��Jsi�Q��qo�l0vE�.�a��y�ص�����V u���kDxq�.Q�J=�/7�/��z�t(T�z/ ��&��nP㝩S�U8p�>9�#�7Z�ƒ� N;����Q3P��@/����n̰{R�A���#��C^���5vJ��ܶ�q��W�뛺��;a�Wɾ��H�A��K1o3M�K���4�`�2�n�I�"h�C8_���]��5k��汦������� !8�!�/t&���Z0�v��)=Y7����R����s卜[<:�(;�~vmAk0���C�Ľ	y���8��������Rw��ńV΢��SNUs3�k��?,�驑A�6�0�0t�"/�q{��󪓴,�-�O�.1�)�;;yqkQaAgO2�S�4���+��:(Pu���t(��������N�0�Wg�O�/Sg����g��d뎿�Z�9/LUG0=B5��ÿs�O�
��{)
��s(�Ʃ^�|c�-�0̳rKm�J���5�K�Fo��\X�d�!4�Syp�yc�M�jV�pB��T!����~����u�ٽ�E�^��`�2�=�e�k���������/l�8��k��.�b��D<��Ϳ��aܯM��= �i��zE��ْ�8o�G�®ZN����D����f|��\dfJOu�~�ՂUP��<}��K�d�g�Jh��f�BJ�u�f�ĸ�L]Z�1;�%X�Q��lB)`�t�����|)��lY��ā{7R�f�s��8�O������n�vVrr�]��X֜z3�YӺ*�9�v>ûN��c88R���'���;���X�%G�����ۜ�W�7�Id֞T�;���)B\�4�C�<�T�	� ��+[M�d�˧�S��t���u^�x�,"ä�D]�.�O�"y�]�8��u��!�|���P5R���!s�A�WB�Rq��{b�p1lkbY�!	��Y�=/�b���CqI��
�]M��(�3wP�K��L�y{Ф�(��Ӻ�1�ϢY���r�SFh_Rì�8-#�O>T��;'�6x_)���� �'<��5BJ��^v�ʈ�S���=����x�9������]_�5ԽSzy���.p1�nbfگ�U:�pb��Vd�N�j�i0��qA��־�zA�l�D(s��;f,_��L����j�}�u4׫�uŧ�r�k���
�;�{ 0i�S�mvji(f�~��L��`;uP����q�o�U���Ԇ�J���X����Z~k	AcK�C�&�}�d��Q�t*�UN-��>>Jxdڊ��p��LO:������ZMyY���;\���������rD�F����6��3 0oFR���}��c�\z��a��%��v�[+ ��	^5>���/tꜶ�\����Ǐml�?qՑk.A*qVaM+�<*�(�0.�_6ի���Ơ�mTrƭT`fB��2BkgNΉm�'s��ˌv��^�Z�|���H���3\����R�T�m�A�q
f^��o �����"Җ�#��Azi�a&�6�Rӥf;��r> <4u��&,�������	����^�wvmt�!ٶ�F_M���1�����dϧ^��i]�w|�j�q�<�!Yr͉뙃�ᛁ�:1�*a�����v�W���������:p٧yTOY�>�p�3\/7:c�ö�1^�lZ�_�;�D��X@��\LR�O���䟺Y���{�<����gu�܂�,!��C����k�1�N��2%� BKHC �G�JֲA��]�l�I��EѨ����B�w�F�ƒèt�R]�Ƚ�OC�m�^Y�d1{�@�|W�f#T��'��ƶ\.Lde?Lǡ>ض�jJ����Pc^�6�2F�>��'W����Fwt���Uo�K��-���y�\zz��^|}��b&Pd�h�'���E�
�ExԻ/�c�����J̲���S̢�W�W�P��'�_}FW ��U�^~���5�)�D�[�^�c.����1.���W)Rk���Ʈ{gO4���Ivl���OcH>��m�[=��ڳރ\�O��:h�鎚�|�[�IJkk���ȸu@ty��a)f���<�}I����w^sdds��EWEEKvw���yx����[M���GΌZ���B�cW���u��v�g�X�Pٍ��ݜ����-�X�4���@�2��Ln�SQ&H$f�n��\Xt�y�Z��ZT��`��i�� �`٫nQ)���$2씮m�����r&ӟ�@l�T�#�L8��I>9�NV7H�^K:��z`�ҌV�}�$｢b,��!n>���Є�B`�2/d�¡ہ�M���bӯ
/��i��b��Z0���3��Ι����9L#w��\?q1މe�}Fi�:��[(�זH�2���M͉�-tt��}Aǟ;OY�ؑ(TK�G��	���0~睘d�bk�t.�yۿz\r͞�T�4�S�	�ދ�O٦�/sj��r�@�Z���hA���v�E�]��@�-��\�����iE��}�'��ͨ�>>���PB�@�`ϡ���ŝ�������]���Z��u��ɭ���Ph��s4�t��m�~���#�Зg]Jw����&��0��®��\���w�?9�2#A3Eؘf-�`��DY~h��{IHMKK�ޫ��t��C	� ��jS���-�)��	��M�9�
�d��jԞxr���uW�K_����5@[ͼet�w�`0&BBu���Ʋ�5���Ɵb��������y�Ιr��+�q�����%xśINݎ��0���6p�%Q9�+�C��ygZ�vj�����p�����n祐sJ��F�P�]�u��Q�m�ԦFC"nZ�TE��2�@FQ��Ά[�CYooK�Z�8��f[Y/gg&\%��-��>Y��p}��1����Y�����m�L��H�zn���
7 �QV�(~dF4���-���ʃ����Ȍ}e�N��Z��[$�m�@1���2��͸f� �\��Iq��1<�
Z*Z0�\�^�������@�QvNGyֿ&):�1�U&�d�PꋇT*�ϬC��5�n}E��svWS�[�p}���v!�"�wy��2�����F���I8�ӌ$vE�)�mb���ԟ�{�1��eysy!�Z}�q0�2��f���ޗn�2�w��LU�M���9@�Wз�k�#r���hW.�F[�Я(��������f�ǆ����9%=Y3l��$6�[5o7ӕdvOgV����G�0��0J�*u�Ƣ�����Уc&�I*�L��.j2��>��:��Y�E��RX�-�a!<;���~4po��֕~�?�;;���f�
�w��A�<qK��t�*�=��X�ݕ�dM|�@�%C�T8�&#��K{��u��x }�~A�X�T,�s'\qn���A/l��������z�?��Kc?2�4���W��;r�B�����bG �P��b^@u;PH4���kf��	�:�.E��V��i)��s䭇�fU�'m�
M�ͮ�+�W]�ʘ�����3kw]]V-�b�8���3q��r4[��K��f�%��K�q�X�#�����3�e	 �ۻ)v�/�m��*j�[:� ��5K0�UhXp��?�f��6)��1�������ԨO�Z�	�i�f��.��`�XE?��ꓫC<�"]�7�4!�#m���uY���ܢ1%��\�=>YM���\-m�6��ԝ���Z0-���^]� `L���S�
ٹ�Gp�([�T�+ޏ�12��g�2���pi$˴��eC�m����cU!\O�vR{��Ƕ�<>�P��ۻ�gb͜��2���^9�T�k�7n��b���L�0Aaa�p���V�r����Ž6�v����j왆��`-u�eB�Ф��s�=����|�L��2�ʮ�'wu]oh.�u���@��6c�����?)��	�.�%ԣ�.���x��Y�.�	���h��B�xd>��!���_*`$$_W�i�y�?!)���%9���	�ak�m.�u�Nv�eۑ�ȱ��vG������$8����pB~�pG|k��锟���*�t���+����Gc�k�b��J��y_�n��thU����+���B��!���D��x��C�V.�:��s�v����O�Bʕ�y&'�<ì�
l�ν"��r��i�-+U�vڬH.�3��}����lϔ9����;_Y ww����Tm&�5OjA�ʹn7u3L�Yٶ��o�v<�FM� �=�RnDa�u���d4�3_]�T/6�����j��c/��Ϲ��J+\�JaH7E2�����0i��؇��l��A�b}Nv��3z){�I1KS�1��{+΢�*�*�z9���PX�]*���\�|�	_O���=ʞT�_�q���2�^�m�ħU�,P�v��+:�<i��������p�rD꡻*�ոVdN��q���c�(�8>��b[N�kepMc
��t���r�2
/��S�=��غ�"�3R�������$Gٵ�X�f�|��e��Y�����>��R�������8�^N_��u{���,ʀ1a�����぀�4B麛Rzj#ҐlL�G{�QU�V�瓂�S����Oԧ��ϻ�>�����-4��D��Ņh|.&%M��2+EIG�U�}R�{��*�gCgt����N�_E���P�C#=O���yL�b$L�����YsFpլ�=2/[Qx���z���⦟<о�è���%�N��K�ɨ��^��X�����[q���U��"�ZF��g��u�UO���b�uW��m�2�mZ�`��H�py�}�~?������������������������}>>>oo������D�x���$G3ݝUw��rݖ��5����Z�wq��W�W�}-e���ۨ1T(��B��5ۭq*&c,�u
�ꉓTP�Z�r:���\(ݑYa��o�\)*U��EF٪�n0��q��u���4r��5x9��9	��\c[VF��n��E�gr� ����,=^��5�Vn�YP���鎚��.=΀c̰�Mz8!���Y�&�ޛz�g�f�3�a���WL�D�kk������m�o�b��#�\$"�n�J�䳗�6��6�V��Y�Ė+�OE��R�nu��3F��C��C����]�{ږ��̹�(�9ة�K^�!fi:K�|*������n�9��������y��7D��_�6��l��s��[�sU�&�z˺�b���S�%�\�q���::�eݠ.KW%f���J�F�U���Er��!fN�kw��P�Ą�˾�.���|ƺY�����P�ꃞ����m�D�jk+h��/&���z�pc���m+95�kAq]9kyP�Ӷs��.�8Ú�Lm9�,;%��A�3����4M�N�����/��"AǸd��,5b�(L9�fs*�آ��7�)�	��]m��4��,�mkIꙭ��v,F��4���I+K6].ku��0�B=qw��llfU%�ǰ40�N!�o��qZ]��9R;ʺ����	�J�	�H�K�8�g-���-b�9L��FK�y�5j
����3��L�Ly-0���fNε�F��g����æʴ�	��9M�Y�;�B��6�\j��?d��H���=�nb\%��q�����"�ch㨦ƫ,�U·"�������Z�U��Ƨ"T��S�#���q�&����rV�W�J7݃y��$�ݦ���;�����o�mF����t�a����4�4�퍕@�(��ɻ]
�S2�ݵ�}��#(-T�n_�vs탱ݫ/Y�ur���Pb����
)�z����Sol�+I�R��^����=Sa��˷:"��w�e�;�W�/P8#�aL��%b�h)�ML����p�4�a�-�����薷���&Nr�oWT�v���ى±-�c�ݱNN_�RWʝ؝K$�!�諸5a2�/�ne�Ֆ�����cJ�����sn�n�V�h��8&fSso����Ǧ��w̠��pO�e�<̂��i��0^f�
���'Cé�v�������Jdw�6�;#����V���3l�%N��D0��0W<`�ĭ^&���з65�s��Yxo9#���7�<����[e�V�JĔ[�1o^R��#�yc5���i�['Q�ڻ�iI�M��؆ȡN��kZ�P�5�LTV	{L�m8YT/�Rl�s �Z�Z���9ì79d��C{�[�E]��t�[�/���F,�b�oE9�&ff�rul�Qu'[&�M�`oQ#r�4喋)�[e�J�����I�m����;3DAU$TAT��TW�)�($�����h'��TPDDCD��_��X�:��(嘩����A�(��F��EU�LQ���ILR�S<�h
�j�Q''䜘�����(����Ѣ`��x��B���譵QEm���&����h����m����mP�AIT�STAQMD�4�PEMiЖƂ�A���ڴb�lSUTV�)UQ�HW#,Z5yb"��(�����/5���4ET1-5Xh�(�b����MPL���7�d����'AQSQIDBL�U!UHV���IDRRN��&)�fbH�� %�J5�lE-%1\�QUT\ƨ���	��ETE��DE7�i� �"*J��/�UT4<��w��9��oo�?3�3��i�+`W�gK\pLWkXəԦ�8�v��/13��7�u��q�ꕻx���52�/�����ݕ�$gJ��֝����3L��,~�]��%V�*��W���Jm�`&�jjٺ,�UV�f���_f�=�8���N0�z3������( d�	f�pH{<��휮g�!�i���|譝�N��čq\�ǝ$f�\�I��Gc�Ww����#e�]�(L&jGuV2s���9�۴�S7_2&Iz���u/�s��]"�PIRkk����S�\:��♟Zb�ڡ�1�u��=�==p�N�.C;%��0�;��O�9�NV7H��z�9}ֺvU}.<nصV��W�Smc<c;����E}S<�b���g�A*]��6��Z1��`e ���<��Q�����u{]��u���"�)��i�:���k����9W5��E�dc/1��i��l�Ъ�ub�t׬��2E��@�U��W1G��G��%Kg���l<��ck!��񈞀C����ƙ�����_lz@+�A���6-ݛga�?�~a ������K��8ͲS�{:���7wn N<��o3�u����j���XOP�n�^p�,�lX����g�j��ף��#f�ݖ.��P�Bk�,��{l��ҙc;�t�3X�.��7��W���]u@znʭL.Y�2�&v^}����5��Ǔ���	���ªb�NƘN�nC���u۴��<Ν�;&2�-��g:�{�v���<�?�aOX�l��Oo�! ��0� %�|_�9b�����{C��;|T�-z��ǔL1r��u����kcz���i�4�ba��s!�8深��j�b0��ӹ�m,���ĠdK��Z|��i�&
u~�m�87����4#�;p�Sl�jX������s�;���*|k/��y[r)�0((F0k{d@|���u�6��:A��v�(s��-���3�x��r�0��!��)�"��z)�T�����T�q�U��;��9��̛��}���C(�r�L|��OV�g�Մ����c��(�sB�3:
͈��6^r���J�t�v�v�"���=50����8%��&):�dJ�%��vN5{�.[�=��R��(`�|vV"�z��zc�@��`�ir]�M����2O~s�ߒ4-\�I�؎�a��Y��5V��G��5kA@����Hp�C+�l�pi�#��\�b�7H��b,�F�n��Nk�/fO�z�|�޶�7`C�;r~�0��q��ӷd�N{<��Yw
�Գ`�"<Lg�a��o����.n>�R��=Y7�M�Y[�"����_]�v~̜������')^b���Tn�ޚ�R��ه��-P[�m�Z�o�չ�	-_Y�i�
���P�� ��-���!�l����QW�b�VF>�W�(}��jj�Ϧ�nt&'CA�9.��2B���]6w�pM}BT�&�8X�?\�&}	��Q�DsN�Ŧ��h�Q�ɵ�y��[3q�;~�Д5�S��'�u枏l�����S�M��z�-�R]n���������6�*�q��%Qa@,��Ua]k����N0i!�JK�PWM����{��<0^qp�T�L�qP�nd��=*��m�VzrQ�c�H`�(S?4w�4%���0d!<������^Do�������*�����`N�9p⫶w�.]�v����x��^x%>f�?H�Hfp���0��o�&�.�>k�n�*,+�ėn��~��L0Ggb�bs��6�ّ'D[*��64'�{C@a��yOl+&��f���EG�J��{���`��x�v��-�k�<7P��@��B,�v��Nr���1Q)WmJ�y3�{�9�s�*/��i�d�}���O�܍��d]�n��{זx�����CkN�+���4..��k�꡼ӵ齺ij���x[Ѓ*��K�4v�^
umD~^�o|A���s��
Ɯ9=���Y��^ \V��ջV���#A���3��w`,�]i;��w�u{Z�V�����{���Ps�����3N�㜆<��f\�]֋�xcf��Mٶ����Ӹ�K�RE����h�X��v��m���L �0���38�3ֻ|b}�A�\_��'��}8�f�K/5~c�U�_��L�ѡI�J9A:/��U�����\G9����z̲���
�V��
B�*����4�)��%5#��s�KR��q�9��©��]P�d��`�엠9휼�ۼHqlY��`$�;/�{ W�������-}���s�u��L�%I�s�8j���� f�t�k�pe|)�;��a�|�1�W�H��d5.��<����jQu���T�F9f`�����q�!P�:�S\�ln�.�>���sޑ%4�ă�z]���?7����KGl��m�Fyi}�WU�{��51e#Za�?PS�9��H�T��dk��w=,��b��T,(S�ʫ�ڳر�Ƹu��Ͼg�ã�9�51-��hSuGu[
�r��a(%�!�7s
��,�{#zv-�1wܼb�>�H`�sݛ]3�6S�:���d�r���nVm_�K�=~�'ǯ�S�.Þ�E���T"'�qȂ�C�az��'��z<�ː�o�N����i��@e1�o�������D���A�)�ҳ.J�[��yY:v��)���yn2n��b�qx󹈜����ũ;��a�hT�4��C��U�X*eˆ�,ƫ� �*\^D��lYoD'6��f�;�KB���ڗ�����f{v��7��;w��<�&Cgp��D��P�[�lC�����^%��M��.BT�&�.�P�8�V��uG17�A�p�0�����H�g�����l��n��5q$񑯏�`SW�cm����\wK��9���������<*�!\����i�^{�]�S��,���{��u�O,���@k{Nsª}<�/b�u%L�fn���&���1�&��}~�5��0$A>���ؖ�\�-�����6���g�3Q��9Ʌ��j�-��Է�u�k�C�Oꏭפ�����ޢ�K�3R
/��b%���s��c˙�X�j�mf0���޸���$�ȿ$f�\�B�Gc�W=���On�$��^�A�K����i���-o4�$_I��,�ۘ�����eI*Mmq�#��`����޺��I��a��O-Ĉ����^�����`-��ک̆��.��:�J�b^��e���:�FHw����v�G/:9� �z<�#�a�6��/B�K��r�=b���2���T<�<}��d�Մ|MvG�O�^N��<Ѳ��ww+�pk�m�*6�1X��I�wׁ��E�$��n��|��X-:T���ﳝ��Lʳ:�%b��� �����ó$��Σ��_����{7��{��C�/o+,�{?(;*v��N!乻1��X�Ct�.F�}�¯p����[o��8~��-�ɔ]O<�[���~��k�nϪ$��8��*���r�(7>�^�ϣ�$WM;�dZ��	�����!sס�q�γ�ld6�DDH����m�ߦ=�����:x�*���n�ݮ����y�C�t]d�чɺہf�/2sP�����F�嘒Ë>���z}F#[=϶ҰT�W�H� CA�C�����3������c[({c�^�d�;���G��a?M0$89���j/���8qc�0�w��Gk>���dL d`�����2Î¬J�]�[���!Ň.5ѯ3RX�e�܈]��mz���>�A�E6�MOzu]lO��D�`��7|�A�R�2�J�RH�3��heY��>O�|��O6C3�0&P�aql�ߪ�}T/&��vÞڌP�ktow.��0Va-I\��䌆�ٶU�-�?4��.2å6*wg ���{�w[^5{+R\��;z^i��AO�xa�Q��$f�����*�.�k�
������0̵��e������1_: ਞL���V��1;�*z�y� Ul��;Jj��Ԛ�Q�x�!mEl�r�uf|�l��1n7X(�TFDk���kv)K���I���/9n�w����aW�Cg^6#ғb�U�E�m�1����>�L�	�5�G{�=��t`�S�h�@��r5��W�<��r�.y��e�`#	�F�+�F�ᚼ{'�T\;ưM��գ��V����?7�FȺ�ې8WBmn~�Ƚ�1)ͤh'P��z{�s������(����~�R�hTg�$=��(8�rMt��zdO���i2�1����ݽh��:��yI�7ըuh���zw�xa#2Dc8��	�G<�@�U��NِƘ���7�s�[�л]a�d�g��&�����ǌ!laV� �C�!���/.ck5`�װ�؉꽣�믳ԃ�d���ٙ������PXױr�a@'�q�&lH���Y���NeW{�>*X^.^/�:�O]@�8�T�gO2�W6�W�ƌ�t(;tpP�|���]|��,%�I�}�౏�� ��a��������d�'�k�PK�XU���6ʗ��	t���U�۞�ffe�����g��� >�C�+���	�v�@�~������.�d:���s/py'�]���qx�=�r`3W��C�e�C�/Jj`����w���LY��S��RF��j��RT�LDؕ�β�vb�A�$����e��jN�)�ݠ>��� T)U�;��E3�oa�!�r�-�� WB��|��[lc{�)�VL��8��ӎ��~��v����jZy�U
0�?ӷe�����1��DƋ��z�*�����=IGpl��s��QNw]�1��Ӄ�[9y�x@���^��=���1Pz���V��B`����y����(4�LvJ����x��5��p0&P�./-F��)m��ݴ��?b���/mxc}���U�z*�!�ϳ�q�t���ז|���I��Fe�ݼ��m��Ä�X���5���Sн�kj�d.|.�*U>%'>f^mk��}�̝a���j{β&��9�\8�y��_��XO�q�I��F�'$Q:���<�d+�Ŧ�;k��W������iϱ�
�i ���pH���o��y�G!)�	ʑ&#���f+/�y�x�~�����dR����l��Sۼ����ʘ	?c8#hkne�Ea�U�͗�;�W�)�.�Q,���I)L8?E����� f�t�k��;�����Z���2w��:���f�K�s�t�Q�E�y�)�������-^w��ϔŌE���dZ��ڤhb�z�k� ��2$�N�A�=/Hŧ洠��ҡ��'�O���5���0	�{W�\���s�R��!9gh��:��v({B���"d�
���<�7~�X6tT�����r����w��`œ�9~&�j*���U�9�[-p����V<�"&�¦�,U�h�-��g&��m��9�k� ���_GQ;�t�3���#�73��^{>��4.��sW��л�38<iG^{rR5�u����K��5(K/SӇ���}`���k�1-����o4��ez�u�*Uw��2�9~�+'��
̸��V��`+"~c�@A���k�vf�|��Q{l�{Wj��f�b{���-�K�z��zu��=P͡��v�H��	�½�T�=-�?o%�wכdtrlr�t�e>ܞO�^y�~�]���y�ұ�W]"�D��"c���u;���"7�<������ܸ7�+0&u�'p�Ϻ�J?)���Z�J���Q�S���t��t�ht_�*�V��)��;�M�A��,W).�T=;�
)B��_��sJ��pR�X�X9G�Bm|�Q������/VK����ˠݺ�XɁh�1�F�U�F�/t����l��gb}5�������{q�Su�ļ�7Al��+gj�y7�����,m^�(2j�S�H�0�z3���ջ3��\�,.D@<�y�B�O`^�w/v�77U��������ڄv��+��ʹ�4�m��C2����m%�����W�Շ;&�tԽ��Jг��>;�YtUp"��M���X�Ig��Pͨ�Wp�Tf&����"'p�ss��N�^]u�؞Vl��q�����hm
�̽Ͷ_=��N®���چ��-A��Q0��E�$f�\�B�(�|j�=���3[��A��P"M�J{���K�Z��`�v4�&�O;s�I�9�NR�,�%I��T�m�Vܫe��30y������uk9�^P6K��fa�7Hr���;��I;LR�t�IIa��Y�g�J;��.օ��>G�E��!�= :�hLpm܉�I|�]�ܲOD��r:�i��@��ubʗ<���L'����"�@!F��r9���-z�����U-Yo|�d:��w}��u�Y����J;����`V��9(K�T;ysY��퀙.�=����'6��]�0��\���ב�ޒ�,���|�} �H��l�4�g!�p��w�dr�qLy����N ��)ۘmn[���$���Yk�=>�gZy�D��L���u&�u;�vb}~�=�[1A���{b���g��n*^픜O�L+�� �x��j�~�-<��9&P��L�SםS�t;�����������Rj���'p�%�i2�X�q�����������������>�����w�����}>����<��h�<��0�i�\�O��9�Gc���ut��wYE��_�Dѩ����]c�t]sn����?m�K_b��,���'�����jsK���gx���M��s.�.XɜZ���k�]�TԨ&�p� ��%��wq����sE�n,p˦!�F֬��m݋0`�g��ʐCٲ=ȱ�E5�R�a.�I�-�zl��֑9�3�&�5�6�P�W6*v�/�5��.�Q�)<=�ݗ#��Fs�k���ui?��w���2�Bt�ܡ����=�q�Z@A��Ү�c)��X8ޡ6�m'��s�;�2w�*5�u��t�Jµ��1��oOq#�I{�f����˻��:V��Dz��ků����:���j�j�� v��=ֹ^��������cy�_7]җ]a�,|M�}w��<i�Z�V�zHػf�vZ��Dɂ��~�`���g7.�h�v�{�7����[�oE��%:i`�q`ڹ��[Idf��ԉb�Prݹ5�u�Cm������3TY�+wW+���n��)���%�#��b������ƼecR���J�@C����*LťlI��}U��e������җf.�mɍ5�R��o62�o"�au��AQ{1��9CF�B�"/Z�P���׆�sn��N���=����J��zM�{���|5h+��P\��O�G4f)�U�W�L�
=�&T̵��7��B��d�2.Q��a'�xd��c�A�Y8T����s-\�Q����ŕ�P<H��u�:���㗳����W٤���SN��_Xy�nyV�K���M,�\��I���:�]�h��e�A�/V�������4�Jeh�pr>�Z��h+/5�nřU�裳/G�����x5��F�U�3n�\`%Iåf��S9����.tl�(�+}�-cf�����)P��ޫ��}i@&���Rɋ�܍s2ˣ\�3���)�K�Rpsu0�5[�g���5��N��ڠ�J�?����%�Z������Us�U�m����}�����˔���ܬ�R� C���o�qھ��;(�7���u�c�.������]7����|iNfa���BU��}ՂX�v���4E$�ȵ�f�8�6��Yu���V�Q�r\\��N�mn����7wSy��(�K<%�t���wU�.W&���pB�7P�s�Bp/h�c�����Cecqb�7+^�n��K�"��e����!;:���)��y�vY�eNN�e�/�*d��۲��o	�ؠ�l���%�vNu�^���/�[ ��5�3h:fETiwf���SR.�C��j��.hޝ���|�ŕg�i�k��v2�����X��!�r��6�M4����σ��?\��FY�V�嚍��Y��щ��z�N�79�,�$nV�]6�e;ն�ĳZh�i���ۚ3��{r�+�so�IISZTTQ�T�D))#d�5M4	{)����TQ^Fj*����&ؠ*e���r����r�|���
δ�j��PSr�CE5@SMU�,O$�M��TAT8��rփIO��54DPLE�7>sp(h")#͠����*�$����31U>j΍�o�8���jMFΈ�)�5��f������e�bj���5UE.�)h���UkQ�rM,��DUE3)���~\�Q��3DEMM ̔T��,�L~�<�8AC��PTW��G Ѕ�H�C\�*�LM%i�J]5LF��AL�$ZMA���72iB#��� �����{<|}�)�VX��ָ��H�(y��MҧA�
u�'ݦ/�#1�췱wb����<�r�'նGc�{NKIi�����y�"�F,�5��9����-b5f�6�AN3A2&P	��LE4�i�H$� :D�)*i��&t��"	_ҫ� 9��3�[�MV\�7z��U��U��륜g��R&}F�U�k�M~�ekV19���fG������ej������4�vj�vB�G�L�I}kO��v6��(=����E�U\��:�gCe:|�4��包�P�����BFC�Z`Y�ƽ����&ä��:�j{Z�4��n�~W�L�H]~ʊ��0S�X�'��%�l��c����:ᚯk#K'5�Q5ռլ�BP"y��9�A��-��_��Z�dE�B���
j��Pni{h��MFxy$���PbH}o��v��&�SsS�&E��Jsa#A�a�����*�8t�v�r�p_b�.ȶ�C��!�$;�ke��N�bۿg���T!�&�tߺZMk�à�c"���牱a�/�����	�ݑ(!�����١q�x\M��Kۄ�ݩ�7�������:�s��ˢ�C��ɸ-/#h��=;�׀���8X��s��Z�&����[�@v2L�+��Qij��-G.Q{Juy\���� �T������?1�0��>������Gశ[*�-X3��ט���TJj�j􍛋�L�4b/ �u�P��5�ѫ{c���m;v.�"����uy׻v�ԃSn�v4�d���1���~��\�ͱt]l#�0ۺ��N�0� ��K/n'�P��9�m�j����-[�[$��?@�I�:�'�@�qvJ�ΞeV��k�m�\���Oɢ3��Q��˙�{����������01��pд�8�{�K�K���Ts�8^�Rq��|*����f�G�<6vN�������� �W/�TwK�@�n���kޱޅVf�vCk��V���ޖ�?�6!{R��@��z04 �fX04Ba����~�fI������\�g����p�gor�^5�F��fD��:���9��046�yOl;5���i�T��13Ո��_:�8�T�#2-�Ұ؜�8E��s��o�k&��ƄD���!b6�Ѡ[ݽ��h�,�v�^��^��}�����z���_B碮B����ע6�7C�;i}�ֈƝGm�{T�g!��p�����*�7��^ܵ�5)���ں	(6���Ű����h����?��꘨|��g� [E���8�y�(�J��XH�"Sm��	�Z7�5ުRm�6��}i�Ή�9�Q"��؂�֜K\� %ux���<�/?�.2u��cn�l��ن�ʼ[�6^������뵜�`}�/J4��b��7Y��b#F�F��6���atS>�ۤ-��/B�+g��v��h��1���q��ӻ�9F�ꈮ��,��ml��q
�_��P�p9U�.'cy��3t2#������k^�)�������b��6��	�BJ�ߡ�s}d�ä�A%Y8�B��;��-��»1�7u�o;u�!c���2S�cȽ�tS*	*L���y��ָ�]��b,l���G����0�u.�)��)�]���E�F�X��-2;���Y�6�]���"e�R�X׷؝�[�x �F�P��{�%h�I�H����b1�����T��W�]W���Q�ub�4�$2���Du��-�Q�9���ڞa�Y�hY*L�dk�F^����b����M�ubn� �����0e���֏�hS*���,�0�k��n'�)����ә>��f\A�l	V�@���W	}.����F[L�)��~̮ZCwv�-�5P�	�S�1��&Tp�a��jDF �Mp�tՌ�OiG1��7ٖ��O��W�̌?_P�%+}/zk�����}a�[1詊SS2ss�������Z�<i���N�5	�_X��M�c�^}�`�=�Hz$@28�v��-Ƿ����I�	wQ���Vd^�	o� Rї��mh5]{WV������t=\�$�Z����@x�]�[}a���r�u��]`M��h<[1��e��k���!����mH�Bhr�5!��Jx�Ui�
ʡ�,.�Nj�R��'^��n�v���"���ݙY&N����z��!����r�=��;�'�Q;�M�@}���.;�r�k��Ej���d{o��d�h3q44WD���������z�����
4C�EvDv&�q�n�ϧ���j���V�P���U�N o�دc��4D�2�P�4�#}��S�c�㦹U'��wv��ݛ���xJm��MV�S�H�0<�o�ޭ�zݙ��,/�a\g�%uދֱ���O�.@X�f����O�b���H�2��N��|j���'�c'fi�hȗ���{�q�WT�a�C9ٶ�;m�_J�?Bd��ħ �JE2��&�~�m>tLbh�b�V�vK���((������0�O������q7վV��zb���X��n-���:oY��Ǉ��\��T��¾��^�R�"����~�������H'l]7���'/���T2���y�n���`xzT/�x9S��3�c��Spp�v�(�wm�P��{id��^�J3�Q+FjiQQ�)��P��\������]�5���c��X��Ty��`��Ÿ���B������Ti���,��%�5^t�Fj���2���<�0V]J謇7um;T�)]^�t�ww��w��6}Ւo&ggAg�]��1�R�g��W��*�F�AM��儻W�\n��%+�� m���$^�;�"�&��%���禚�a',���j�Ʀ^Ż�G��3���V�6B�L�2Op���z��xdٶ�Q Ė^/�\��O����_�?��C��)��M�aOx38���Y4��o=�b�۔6��)86���P�,�����y)��W���@����֏!qa�@׆x����![��H,���� ��B��.�Kֱ�-v��lͱY����������wtE��u�"]�`�8./��5	=tŶ'�	��ٞ�B0O)�'w�����
��Qp(7.�b_{ω�x����k&Bl��a�n���&�����p�p�tS/Z�!�z�nb�m�FCH�{��lO������N6WM�Mn�Zai�>z�7X���S�9�h4��͊�'�0�z�YPH�3�^��(d�í������0���9�kz&n"�	d�"�N�vt�@v�2j0���!���	�b4)T�H�p�4�aVfY�S[��+z�.}v���oP.�0����&�SsW��2/nbS�����ǌ�h������lc�M̡&����E{�5��~��_��B���}��o>����<4Gٷ�N�_
���/y��O_N�@�hӥ]Hؓ�3����V��Bn�
���}\��d��cV��Nm=J����2��e�����Of.��k>��J�r3�+0,kb�Ӎ���L9~U{L�;`ul�\w��A;J��;�i���uG{D;�"ds�_=y��ᄌ�F4å��é��m^��l���#�_8	��r��*��\oͩHZ_gǧ��8a.�Y�f�]Okl>Mɳ۽�b9��3;;�u��U��A�F�]�t�Nո���4u1F�FF��K �L:Zj!�p����a+v�w)��{��v��[s6��e��5}ٌ���,j�Ϙq��v-�)��{VP'�����MC���Ԡ�N,��}��du ��=��]^Y+�t��<�U ���mdw�y��EҶ�{h���F���K�U]�T���ͻ�N��ͦOj�L����b`�����gϢɫP��!S��<;x���y޾z�'b�M��D�- ��y��C���y���{]�����B�K��.^���� �f�*�� �y�s�6�.��X�7�{��Uz���pf+Չ���X���{ڕ�v�'���<5j��ݷM�.b�ʬ��	�����#�cP��F����8�`�����Oz�	]\/���L�#�fF�ҵ�7�8�����ڼ��U��"&��U0y4��@��:����E�Q=�`t���g5Ba��Й�W�"�[|A�&�L�if�����q�es]��=��}�r�+�����.����g���_{oс�fu�!��H�o�]���	4�tw2EI���^6H7d�/˰�4�n�i��\����X� H&_��ɨz/|��]���M3����T�v̚���[��m��T1����RѰ�I$�~���N��0\+t.�0;w�&��NIXПӾ��-	#>x�)�歧�C��F�H
�����c8@���=�ɷ^��~�~��K�S��e4���I���'������:���$�NF)iv�ߡ�o��%��4����̛�14I�pW��v��wo��L^�����8[�"3���O����ot��<���.��;�3&�V+���ֶ��Z�yv	̢��t��i�x�Wha����pJ��%�G!.Rd�)j�
����v����n��[��0���8a����uEm)�{�s&YF�`:����,���Mn�l���i5���w�U��-����ϖ@&��t������ �p�͈��l�
�7_�<�:��1)�z;�������Z�|�7b|\J uE�����~ӉlF��SC<3�;@����O���Qwva������bܽ��4\���y'W8g� �%�j�Cޛ	��/�ﻇP\��+�%Gc/n�e�7:-!ꊯE׶�*���*�M���{�"m'�)Ez5����7���m\f}���u#e�k���������g�a���%d��O������q2��q�6ԋ�P6Z���T+n&��oENl�+Y�t�n�酨���PSJ�z�̐.i��2���zGnń���;��].[R��ӂ���)(��$e:1�n�ڭ��ű���ޮ���H�kp�6�-�v����]-��{IT�$�g���ߟlV�������^�Q� �eK����ׂ�-mlr8F\J��O&\�'r�(;X�%�8u�)����e���v6`�O��,KGt�G�)֭R�o��We�Ί�X��fՁL5����  f#�&+Y[8�[W���f�7�5�ΌX�+����˩�b/�0-y�j4��`M��F��-P�C�?������
2�Tzoy��@Kl7.3�f�ξ�z	���9&���{W/#�Cf<m�/K�r��T ���z�%���a�M?r��$��c�9�{ew7`an��F��!/W\Л��C��͹X��>��c��Xv��.�ՌY��ǐ����Y;hT��p<h���gt�a�WU.�>��%���J@V���i@5Y m0q�Om�h��{|}��TM��wI��y��,Ү�/>�^Y��u"�5�9����V����',0�7�a�XM@Y�s �K�������8���eo���������
C8���vu]W<���� ��[�]�R�����jx6V�h{���
3��2�ၯ��)_Eb��p���}�p����Ay<xF��=#�b�b�'C`�!D���ђ��U�T�E̢ʛ0�u��[]�I�
�P&J���Y���V$��B	vC��S�{���n��5��P���7�o]��#)N���̱��-�z�k�.8�^�bY�6��D��h�P�q�i�%:�Owrb�ĕN2�~�^+�Qs�_�'�������!���8�C<��e-T�u:r2����G�4�-��E����	��C&*u�/� Ȣ�PH��37���y��N�n��4�@��p,B�~㖎B�n!b3�h�s��"���;[�w��v�U{Vn����5��А������]�v��O��5�9}��=��&q7��;^�v}a�V6F{�xx�3Z��EfS�+n]WzK��ݦLgb�V�JDϛkd�뇜��t���uGM���\g_4G3�o>��P�-rUҸ�K������頥�]}|��ip�m:CH8��3�|�P8�$�#Is���=Q?'���㖤�y[���a�p��y�騂�8��S��\�O�V����lvo<k�uq�쪂�, R`�!�7�s�-p�bl�+����=>�g�������������������������矟�߫�O�/�ޔr��3Y���x��#uJ�Lg+wj�tn�#&���[��Yz�yP&"U�tޓ�^]��E���ke�BV�F�b7\F��|`ԧطf%A&	0-�·�r��5�xq�g������j��[�k;��%���B���M	8"�=�M^�xh�E����R�i��:��Jm��b���UYk�`utN:�L��z�;������Z,��W�.�Y�3g	�V-�ra�S3gLY[nc��*i���K��L�ً����yQ�mn�u�eŹl���Z��/���[�t*�]u�5ԫ6��f���ؗ����Io�Ѿ��W*۷�i��2 ���̵n�ۛ��$(*��hi�ƚZ������+��﫭��nMX�a�%vq[�V;��r���ve��9Gs\�7���Qf�d]�2/�;�8�&+7�1E���h�����k�J��}(�X��F�䶶���y��M��b��K�ۛX��C����6T���$l����W],�M
�@����#�Q]Ӑ�itd��i�;[�i�Z�X�7���բp���7hU̗��{T����co�:C.�8���I1[���'�Hѽ�k)]�RcT-�@^���z�����P&]��Wun��=����n�ɵ3��B�L�As�dn���uy-��uo����Z-Τ�pV�Xɀ�`��x�,&�[��lX��Ɣ�����E��v��T�v�H��V�k��<`�71;_Z�]k]���W�T|�oZUJ�ȯ��"�[}ۙ�;���0���.�O��*2f�n�.LƎ������h�=��ޘ�.�V�<��i���k��a4����Nūzխ�̋�D`�X�����d1՗�Kؖm����M�&`;\�^��ܕ���L&.Gږ�d�t��wV���uzj�v��3�kDH�W����rr&^��Hi����9��˳q��	Ab�d���K����Z*���ˮu�.��T	N�)6\7Q��'(݅�*S�ڙ�Nd(���m݊U�s���ˡL�']	h�`�TW��L�0����6Y�̅_��;x�-����œ��|i`��.�ܸ�3]h��uf8;�yMdUv����������6��A�{k(�ea�QJ�E����������j6�S�mi�k7A�h��WP��n�d��;d���@�����{��t$'f�G�C�Vێ�l���QH��g2n�$Y�u@��8Ϫ�#]�&��#K�0m��"m�b�%�̚9�ٱui��G��1[��3�6������L��"[�Q�"���/dřD��)�gN�+� zàkRś�r�$ؒ�`4!�cb��<�O�jh�4��rzOe�ݠ�x�t�
SN�c��U��^M����	��M�a<IV��v�錺e�m�L���x�km�6�-6�T���_�<�}�)i*���Bb(?mS������A�A�F���IED�2�KD4�T4~^����%|��������J������r�9:*�("R���Q�)X����PPR�gEm���_p����)�H��J������(la���
h�C@{:iO��m�CCB�}�TQ�t��E'݈�
���	B�!(�	�6�����Jh��&�#��<��~A�D���4�HSMJ|�u�s���۝�[�z�D�*�[�-
�(��o�� �wmO"�*�[���M�P��-3����k3^i�5Z�3��Ufl��/���"��,��C�� �~�N�P�����AK�^mVU�{�4�^.�t[�Ϸ�}��B��sh��b;��z j�W؞/0
x%j�Lq$�L@�a����'����B��s����%�R����~5���àN�$�}w����2�ܾ�h�L�B_�f5_.�G���z1yU�
:}­��ʈ�i���sݻC�qw}���sL��E:�k+^�Q�Uk^)Ʈ+��
����"[�.�۶��-w�]lΝ���u#e��S�F<��0`��b�R���6�E=I�:[�;����*�eP�nN��K�^�``nL�߼X^չ�-����o&a�r������!�t.�y*��P}�����8���m��<S,g����==p(�̱������%��#Kd�J�?_�Y��y�n�Ln<KU�i���/h,�-W@��\�M:�/�Y�u[�Q�J��G/p�ݳ]�S�5�ٲm]W'������v��R]X�õ�:TI�du�xk�?j���1M��C8��u!��;��f��{DJ�ۗ���7�W�q�(�	A/SmCY��}�"6��cWY��#G����_y���4��imҤ��.�qsfۙ��r�4=ђ<�7K�Ʈ�^����,y�[+�%��5=Ɗɷ��Ͳ�L��.������U����xЖG{>6���������u�W��M6k���J�o��; #<�	��z*��i�����=RO�L:�I�7u�w�iP�m	t36���;v6|.��}�`G8#��u/�� ���̺5Æ���06������uܧk��H=�(Bϋ��Ш�{}��,lb��h��Q�o�݆�6��Ǭ��;3Ɛ�{"g���Ee�Dp��C�4מ�Ĩѱ��/#�� �D3����O��l`���_k���p��u���!����J�鼣y�.臻�ʹ�E�[��ץIz��,C��SiN�9����!2�xD����N�6Mw����`�y�z�f]�;C����v�>�˾A�B�Υ�>��;���h�#�
Fh�%L����mR��y>+�;�m�N���zU���M��
0�"ktE�����ـ�����ٝ���\�:�̙zbͽ]�s͖7c+������E�n�����Q�t�J���6���&����W�GFm��V6Y���w�������oׅ�ݚy��b까�B�%4��=j��ɹ�2(V�B�ؙ��wQ����!\��4��>y���=䌪�d�U呱����f�+�JMה��8�,9����;E�_.�R4���H�;6T}��&��(�ܻ�+����~�K�3���,z�@ש����Wv�<�Nɢ�G���r20�ڸ�;��x��$�ǜ��)�_-���m��X�ouQ\��������-г�;aw6��S0[.D׻��;6ǵI��Y�ln�k�������FR�^Ս �������sE�؄�7n�E�.v����A3����;�Z�����ށ���Y���*Rɡu�v�r�1p*�Sp2�.~=����{�|�x�x���_�2c��1���7_*mu
՚�E���k`;�;b��D�X�ѵ[�a�NN�	�Om�[�-��.���*���6H�+��=�x0�g% ��e�,������2���T斓�����3�v=n�#��uh�1^��n��Ä+�݇�-������qi��nMX_U�����2�R�@́�s���/����̶��K���}���6�A>�y����h�s�T�u�IN��V�g�.�d�Kiz5�r���ޠ1�)$������2�#�����8k��l�S]h�׾}���$7W��(�5"�"�kݸ���3X��9��7��( =|���n`ӵ����qR��!��u�,T�Vø�����dkzm�����z�T&mu��Ԗׯ�2=EJH�0n�L�YF6A7[��ü=L�� ǝ�,�td���B�]�=79&m����]%au�ٚ<)/g=��\U��'�t�W�[��w]�k3_y��''w��y��y$T�&�o����vdH���!��B�rb!�����z�y�m����۹�r~'[�EXn��:�[^��@9�32���?�g3B�7��l���:��q�p7I�fi�^���<ݬ��N��9�+Gf�eĤ7u�s�X�ǚH���U��1]�$��}{8L#4�J9;�S���y`�w�LT��;J��n��/^�������]�,eb�3�8Z`�S��I�u�(�5��w����K� Ƕ��B��{�J=��jR�����3D��S�ס�Νƺく�|�i�=��P�Y�w�ā�H�]�t�p�7wd���Q[M{[k�M4c_�������B���κ�\!gr��h��0j9{�t��d ����e0�3a��?�.��S�i16�e��N��z���|a2��Z���s���:�pO~�{=Y{��s6�T�TD#y�K�iyx���=.�s�a�V�5�a�Ág��f����֚�Ǝ6�7t`g@�k�����2H9 ��׿Y��8��z?|PB0�#���}��{�-ļ���n���_$ط��o�(r7��墠C��N�cy֭'��q7ܙ��Bɘ�26j�7(^"��wyY���Ɯ����U�'/����L�e�yz��8�x������uc��$P�>�?�&�g|)��/��a��h�'��i�²*�Elf�>��jkM��{n� !Tmۮ�̷v,�/�-��)ʮ��r�7�F��C�~��Zx�W���gF��:�U_=�
���m�#Y�tr�S���0R�=���E�ދi�(��Z�EP7�Q�U�[#�z�g�����[[=�m>����ung�,�S���~��|}炳UN��\�w�J�jd:	���"ѕB�;w@D��
�p��&�FN�/vv���={�#�@/	�=-�)��]D�N��ʭ����n�wٷ�F�l�ٓ����"+�H�b"��JJ����L��SusE��s�L�#\{n�K�G�%y�c�=�V2۱�hF}H�жÿu4�wz�y��u�{+oM��M��vC���p^���B�Th�m\�n�%=�.�r�x�!rx�g��?�9�,��6<�T���-r�������wv�z��I��R��;� #��@N��&��𞲣o5y,aRh}Yn
�����y���C�`���K�����̄�Ԭ���;���Lt�,�����<ڳZ�.�;@��� t���y���Hí�a��˭�BX=���f�3vֽa3(G�Ծ�Y��f��2���)Bŕ���{����G���\3�S�--1�=2r�\�X1��IVN�ًt�mەyq����4.��������R�Բ7d;�� La􉚥i�V+�C~ԙr�q���\�,�r�2��ܳ�3Qyu���#B��=��Cۇ�J=ϡ��m�[����g-���ڻ^�a���Q���Y���%ct\�/#y��X���{kU�/��9��XU��j$p����u�|˱~���"���.���6�����0�@�� lS����H�<¯���L������H��G�E	�F���Zt���.��(,⁾a;�Zz;��&��sF��iP�ﶮc$jAmx�҃$���y�sNw$8cF�.]�����B�f��
�E{P����E����T�R0�tiټ�U�5��Zy��ҷSV�\�T�EO�������^n�,�Y�[�&�Џs�w{1�ǁ�u:^���?M�oy�dq�Z�ԼF�#�Z�z7(�4�&A<��8d6c��pB؅�4�o����s$�C͜��Ӭo���d�Ѯ��6�ڊ�4��K���*��o��u7l�vm����价�g--j� ���޽��p��q�nj�T �(hS8ˬAem�3�.��>#��zU������k2�1�vӤ��]Rp1݌�0���^Ͷg������'��W�-5�^�������['=�}~��0�B�����[Lj��T΋��S�N�S{�W/}��������[_^HdK����)�s������!��9�"3�5W7uOrI^�M iWfqY%c[��qF�;/7�`w}`>���pQ���qM����_o�lMn�ü(����7|ۧ�w��d1��{|Âu,���5�[�g�jn��\8�[Z��L����u;�<�LDD\R$	�:��s�)�(
���}��y�΋�9��}�9I%��E�c�C��k��3��U]��xo3��ae�e�O��鿓B�0X��;l�A�c�ۊ/�U�=�8]�4Z��&��]P�^�6P<�%.YJ�m�nCDa�ٍӼ���r1�jj��7>�y�T\�Ko�2T�z���na�L�;b��w�Ϥ_e�={v��v-��X0Ms�����z�.��y^�48�Y�w��6	���b�jL̓l<�S[M3b�Vn�La�P��@�1]LG��څ�np܋6���H�M_�����f\T�+^f䉰���f����P��عp��ΰ��r�?�$������hA1�*�5C~g@����nZ9��EoD��.�j̫Z�'��jʥ奔f}̛4�M^���J��!!�k�l�n��:�����H���	A�"�@w��U��R��̑n��L����:�.�;�;�,���+g�#v8�b��д�oJ��Ϫ��OF�3�(�u�\��`�
C�� �ڕ^�-�`=+���)t���e<FLҙ{��۵�y�A}�����>��:��_%T.�r����m͉�ճO{�:K��[>�ʉ>�P������UG'6�ܹd1pۜ���A�ӗ{��ޱ�N�Y��W���;��J�h�j�*��k����b9{���so=�|��>���	���
��^�G����y�Ħ1�aԎ��%?VP= oF��&�a�!�&��x��m=V�N��V<��|�v7�������֕�X2���A��Mj��œp��t^�襆��B3�[!`�R��b#~�7zl&�n�s[2���n���;u��+�c��h2�("��wr,ý(t£���h䥪�ǡ�����NcQ�VZ\�*�L?ߦ��#�lU����&$�$u�b`��NK�Org3ss-N�&�B��4�$�t<m,����/�6�1?w�
d{){=��Ɨ���}��n�
"���S8�� �1礭^n=��*��ԡ\�מndn���}n[C��Ռ��S�����v�~��a�y\�*��QZ��S��~+_�JR�i��q.v���r�%�}}�_��un��}����0�9Cy���hʡܝ���pj׵�W�*�>s�53`_#:�g�����2zN��݄M��܂�и�H�ISmU�2��CZ��n7xN5���Dc�}lDV��I_��4ɒIO9ݮ�N�x�=�5S���q�[��x(l�¸��rZ�"��g�i+��T6��O�0��/=��<d2m�5G����#S�oz��6x����^�����������������}{���y�������SnW̥�������:5�v�̼�����GtKVv�Aj��v�u<�{y��WZmk!c;�����(eƬ�b4)�T0�D���jض୩oPu���5)�8u}���g�,Öѳ]e��Uh5Y���F��˭����D�Cd�7���3r���I��#���]{��lܨ�15/���P�t����x����]�f9�f�a�e �	y0)�1���p�����\���S��ZD�H<z3C����R��,�ܾ9�յkn��悝�[7^粞�!��ٺ�������ZV%��"�-u+�����ҒW�|���+ݿ�7��;s����f�0��Wùj�˱�qy5Ł!��W��x�0۶��>����KL��5F���=��tO{��X�-B�F����V�`���F5�\�;Z��\�-���+e�5�%�k$��4ڼ�@m��Ϋ<0�����*�F����ws=P�y,�F4�n*J��V�N]�=PG��0s�2�ӌt;]�k�M��nYƯ�j��)iY����Qt�݌#<^Z��[|o./2�f`��Ғ^CМ��nvԤ�5
4Ӻ�2���2�Q��_*��ϴ��L��7����\Ȫcf:V˃%Ҋ�8�hͫi�y��K�+�Ի�(8R�[�fl�2o-�t�����G�|8mĸ�jΔ�/�U�7H��`;���^L�O*G/TyŻ�//}[�V�eଡ଼wkQ��	M©!�Y/*�Q�Aӵ�C��3$�S�#}H���T1��I�Y�2�Y�vˀӱpkF`Ee�Y	-.&K����dCQ�S���o#eݮ�O�(��!��uF��l����R܃�G$\H�ն[�(�%f�wK{Fmu�'�8���h],:����<75=���y�x�@e�GU/ww��ޡ��#�b�i���!+]n@�N�wg�����2�<��b�T��f\� �S�t����Ei�0�S�\��'kle_α�1�u��س&_Mr���[� �������X��u(,��&*N"r/2�㲆�9�D�}����S��T��"Tݠ�ҷ�-�C/@,ȳ^��YyV2h�iĭ̇b�I4�ȉ@m�p4�N�B�#C����X�Yu�!�W�**%��X�'^c�8�<��5Ti_�\3���ou��*w�0�I��G:;�ԙb�I��u�;r��i��M�M����֖���z*cp�ȣ�*X��KZ�c��h"�p�z�}���K��J��!s8N9Ƴ�x"5T�j�t;-�rM;P�T$۫�t$e�x��0s7f�1H���'�h�];t7r��9�t��}"��G*F�����owmwB��߅�:p�֙��4�e�=�ؕ��J�;��
�Сґ;y�,_De%����8l4�XnR�E����p�Нg	�YЃ{�l�Ͳ�x���w[oN2�Mf�wv��pV�J!����G��W���W�(p��l�P�ҕ��:]E]=��ӥ��кОHj�RiB�/��
hi�)�
h.a%'mS�q)�IJi�kɠ�� ��h)��#�9+�)�N��J|����ihӠ
4[--�2P�5TDh+M(D�ۛؠ(9b�
j/�$��4i(��CAA����M��2A4����ti9 h�<�4}���	@W��k��1+M	IER�?��9��~�:^]
�A$4UPe�5�($J4@�@�=l%��+�Ͱ�
+,d��hXį��z��5��"d���}�xb�y\J/%�͝ۥS�r�6�|׍��Ѧ-IRi��H�0
!Q!MQL��QF����Tn�t*�TQ�L�M� �&���Bp����g'�����3�r�jf��'*�"�/�q~y"W'��{����%�������bϣ��ܮc-O5Xw���1zېEmW�Hąy�>'t���$#<�:�A�]>2������Y�y���6ܻ�FOH}�T;���DԫuC	�J��	P=��oT��7�c2���02�,Ҡ��G>+�P�UD��:�ǷH6w�N���c)8�-�����M!Da)��g����`+�X�'s�W�wv���X��J.�!�����V� �g��C���'}��V���9[�":cjws��%K�P�0�6��)k��;b�
�~IP�Q�U�NvQyW�y�������]EZ�ȴVRSs�n$hu^�3=�|]��7��{{��ݷ��n<D����%
�7}ƒ��4�ڛ�󭖙�k���jYS�tԝ�
�F<�s0oU\�N�׉� �.�֫�9�}����367�gڬ���A�F�TK]�`�,7y��W��da8h����3&r�K�e�@�ɋ���pD�FΎ� R ��nn�swQ�5r��Mǳ��b`���_k��*8 ]V!F��Be���c��N&�7�jԖHQ���X|����G��ߡp��T�-�P*�L�IC*���.��Q�<y��k�g*��u"��LE;{������2ڑ�����m�D�������"�Q��S��8��t�F�ä!�(M����7�w�v�-�$wn�g4�Om�d�&�l�ۯ �ÀB���T2-���0�{�4��t�sm��@&�+e���;ag�x��^��H\�K��l7g��M��ܼ��D;==|�GZ��H���jƂ�#�֫��`�>Y����u�G��U�z���zN ��Uؒ�ޞ4�N�M#*.zoV���0_��ͻ�5���y0.3q�is��ر���V_�ǝ>���z6ǎ���V�3�<��_��nO������ڶ�,���t�gQ2�WYfs���ip�w�p���rް�G9����Ϋ������}��]��Ŝ$�h8�@���i��O�65k�r�.��5�xf���gH��-!ǩ-l\���ۖj��ը$�bk*Nƕ�u�+��q�r����W3��@I��'Y���h�U��p�V��75n�~M-%����E�u�}���G��,�=$w8n0Ic�M����r�!�F��[�7�a�ěy�:3T�O=Ǆ�����)wE�- �'��gr�umjwzA"",Z��x�&��.�#������S��4]���-�;���
+��_�66
�窓^���옩Җ��o��L��B2 b>�{�ܝ�b��i�*%ԁ��Wa�y߄��F�ϝ.l��V��VooJ�N����k�=&�U^=��/SL��hPn}	"���9v��
�����Ϙs���)rMP|�;��}ّ"�M�]p*�^����뀐�h"w�v6rE_��HH�����<���]��ٜ��Y�0%?D6�#�Ƕԫ��S�+�bm)K�8����T?��N;����Y�8$��n�ot����U]n��G��)�������1ҏ9��7��vIZ��%b������JU�Zy눲Í�"E�}�˴���
]	n�v2c�vNįT`Q��
=ۋ��J�m��3��`K_R�DY��4�/\�oz�6xMb�ТX��Sn-��&ZO0�zj2��3V���/o������`���	^O*��O���nfx��ѷ|p�1��ڕ�Fh*�6�|y����!��0R {��^qD�0�s��mӧ��Љ-�K(Mq�n����o!�_@8����\�ٖ.��4wp��;��h��Q)��ZK�t��a�jK�0�����w]�ĉP��
����h��A��&#݂�kO�p��6*j��<��g9,�Nd�#}ã3b�l[�p����1��|�[���n�����m6zS҆�=�����>�Οv�f��Ի�7<'���u.9X_�E�K�b��^���TN��ޯ�v��=�2�(�i�t�B��dy��gfN�:���ԩH	p�z��>ɧ=�v;�&L#7~/�����˥�~���F�b;HX{�%BѕP��n�+aW
�����33�����y��a�3f�2��C\#x,�$�s�H]���p�W4 �gd�W�/�p��{�rh=ʷ�����Ct�.v��$B������gq��T -p�A��[!�Y��`H;4���Yq�Y�)<����>�l"�w;������q?�~uk��[��Y�6%0���;Y�4BϠ@��~�r�@Ո_.�G�ux�J�$���v�)���Ѧ��%v�oq�s|��C8���h�K����Gt���a[%�������������V���k$1�=�Ylz�Ǩ=�J��a�`�5I��'�.�=��;=�����;ㆧ �n&Vŧ|�}�x0����>�ږ���Ӊ�4uXH���>�m�w�`����7&�H���Ɋ��%�#u5�韽�]�~�%W�;�mt�Lی��[�fQ�m$nFon��<-/��%>���ݮ�ܖ�H��
��E��O�B�hI=��f�}��"-��x���wS������x[@9>���}��ҙ�5�k6�����ő�Q��a�&t8A}��]�Γh��C�s8I#6a]{�1�~L�a�Ih��C׵؎���gc�ѧ����Wc��]|'�t71ݰ��?0��}+/����x�f�{���!J
��%uA�{�nn�ӣ:Wa�̊j�ht�s$`��.V��f����4V�̤��lDF�T�ZM�.�ʷ��a<���tt��ۻQ��ӭ�����(m�x������E3&�iw򊾼ɫ�_og�����!`i��Fv)�FC ��+��$��eAșF�#^����\]����
�9�YJv)�䵎~m�"����i���\s�(!T�U�֭!w�,c�m{����hʹ�)�~�X#o2�5W�s[�g�������s":ѫ����B���
Pd֎OQ4#�)U��u����4�B�F�c0��do�j���P+|L�"#�٩�i�{�*/�q�n�mU�_��Ц�q �NE:+�p�|�&��B,m�OQ���|��7(�A�%R�����Z4�p<�g
��ؖo��o\��~�e�}��T��Y�(�а%ǉ���۠��(����nwwON؎^����h��M.Aj�{��S���q�<B��-�';rb�`c#������/�Ϻ��ZFy.�Ռ�o7��m�5L��_�t+�V��r&�Ǒ�7��誄x�[���%P�U��/�8:m����7�:����ܶ��f���^��"#ꝥT��J��y.u�܂p1��N���;fE���iI�i�X�7s� � ل7E���K���X��e������8���l)���~`��;���].ǟK{�͈�{ޫ{`�:Z��;���i��x}��_@ �C����J���g�:|�9���Nb-g��1����e��5�gR!�X��}}y�>�C�Z���R�Na�׻��Ci�����J���t��#������8$�g�d������ص6s��.x
�������A%��7�8����Yx݀�g'�y�=�Ꭶ�Z���+�����" i�[j�ܳ��T:�J3��o_F<氯96�~{�؉��^\Z$O7��T��O]��u<vɶD���zZ��	CǪ��L��0HԖ���nr����Yv�V}I����k쫓8Y�S�@�~嶺���e,������7U7w\��A$��^�ʨ�gD�4΁������}|��t��l��(�����z�urE��g8����g����+�Da���6f��:S���;(R�V���!�5�Ƚ���egEw�*y��'e��L(U�rMBǚ!2�nc&�\���9ڽ?hcX�Cp.�5i�JM��{�*��[�����k�����DE.(9&�)fϲ�W�v�Q�X��ӻ���Q��K��v�O�]h���v
#�)�B]�ZHzR�Cy��a�q��d��7>�&��m�U|Z\�@��7�Ժ*�m1n֬K6���3�ep���<�z��*�u����O�8�6��e��l�gJ�^iʤxi�|�}~�F�V����8��һo���gj��(�Ŧ�8���߯��_j`T�7�UL�Q0��o�S����\!p=��]R\�W��Y@�J�q�Kv��uH�S��#i�V����t\V�pj�9k��C?Y�b����Xq��]7U����ah	�χ�����8j����E[^Z'A2gă�L5ZnyDc°�4���Og�M��_�oC������^�;�Q;\�|����b}J��Ù��n���h��E�{Qa����.e�^��l�M)��m7���Vn5�J����C���6�}�~�ω�y6��#��Q��Q�WV	�2�t&��u@�Go;�󰙏m�ͮ���++�:l]f�'����@
�S^7!���ӷz���oM���>�M�ח2,��y,��V��zQ~R3j�cw[��i7��-���q�&��<���{��6;�a��	C��~XcӃځ�*�kl:����<������J��.���SsNge�
��b�������zxo:�;�z�c�|�=&>�|��3r�{0�d�믧��<���Rგ7�Eߟ��XD��h1���.'�0����6��Y�NOb��^$��z�T�i�@VJ��9z�_:RVE��b%,�X�8���ȴ�}����z�6��U��Ty�[!��h�\\!��b�W��Zt���׼��Zo��B*� �-����1[�Y�V�[5�gv���Pz�7g˹��t��u�j@���k�7u+ckV��#,I��N�^Ó=ˢ|oO�ݯW���Lۗ�o?��#�aUY𚮫��A��#V�ˆ*Y`Fa��mVQ�Z�-f
�;�����g
� �H�P]��d�� �!��<t��p}2�o���b\4�G/_i6ૼySP�?�d�ۈaC�U��m�Hd�b.����"�4[6�.]k�-È��5k9�r�0�1��	��QwJ��X�������k�����^]�������魜سv��̓\!ɆW���u�_��>���s��9��_����D���&�ZHFlȀ��^Q�;l����A��ͨ���٪����Xhk��+�B�SC���^�πV}�#�zj���[k��uZ�wtp-���N�x�$�y��`��/װ�2���9�su��P���u�b<�ۤ}�ǨhO"�+)k˛^��~$E3[M��[s��.�IU��S��#RB��ƒHm�͵s��opK�kq#;k/%�V�7,��`t�p�D�c'QIAJ~����D<z�k33yٚXEd��m�5�w��N�����ق^�0�^^���p�;���k^��^h�f%�����ODt �ϵ[��^/<PO.�O�
��������_����������{���w���������{��~~~~~�}�3��^�mc����O.���q$a�eˮBewi��//.�(���C�9q���L���"l��xq�Ŵ5��&� ����$�5�v��gt���#�*���X��;q-�7j�S9.�b�����J�j��o^�˨v����W�+�#+i,Ȑ�ܔ��a;�Y�[̹U�(�A=D�Ó[0�ڻ�3r����75H��l�Y��ܻ͗���AO@Bny �{�mmĨ���3�_t۲G[�;��˥lF���ۦ�B1Q*��o�ٓ0
���1��D��|zn���̦����h�79���h��e,l���a	W;,����������\�se^��"~��-[�v��WR��2�9R"`�dQiiٵ{�����M�/r~��C$XiWa�t:�$���U��-�w5T�2�7!ih���*�UL��D���j'v� ����{9l[�������*�=���9���qv�ﴄl����I�Z���a�i�H��%�Ӛ�����B�bY
be75!i�S*ֆr�	J������9��;�u[f�^��-#O��.mLN�yW�p�oI��-Y�����Dݕ������ͮ�S.پCnGj��e���W��ۻ5�r�FT8dYE_I/�Z��Y2��q�u�+ ��Q�Ҭ�Kl!�"�ʠ\d}*e������s�ڽ���z���-v�]0*�
���T}�x���7�����W.�2ٖ^�[���4xJȐ[:�@~ Wغ�v�w)�B�b)�����r���|_L�:���e�va������M��!�-�Jԉ%V14�w$��s���O7y�j���p�ݾ�uen����^gZ�p2)vq�m�켏��q;OA:��dNct�&�U�VSf�x�kA�j*�$l��}
��]���/s�i���z�,�I��ӭ2>���B��_m\��j-�jv�V�+��yy�'tnd�6�c-��·l��vp�-����T��vA�wY4$�f�<sr]ގ��pV`���K�^y���zM���4&�I-��i�u�-T��Q�wh�s�V��78Ph[��w�9t��.�i�a
�ˋ+��3
����:����cz���v524�f�Pa��o5��޵�t�Ώ�ܒ�cUn��\����,��B��2��p�g�{D��h� �	P��Y�zD^m�ΖT)��$hnd	���Pf��p�/8�dk9�Q��u�/k��B]�H#F���R�&�d�5"��*�^�ToX ����b�JQ�V���pe��_1׊f�̗�i�81.�9Qͅ�jL�5PF����{�y!�ܽ�S�-��v��u\�Mi����`�]$�k;���yhY�.�se���gb��p�=�S'�`��^��rjqC��
.-��b��e�x�m�h��֓m��m��n���3U3b����_�9<�htۗ��#G�����i)

>������J&J���Ѥt�AA�>`�C��sA�] h���������MV�̀8AD\���`<�КkȠ�ʂ�?`9��<���b��Yk�����4�4�آ�����S��[g�:�|�ȉ��槗%�s	�ej����E y�>lP�5Jh@��!䚤9h
ym'6R�4�Miit%(�:O�c�Ei4�T�SZq�J44{	��Pi����ڍ�V���#E�ŉ1h�b�kDT��7�1�������{￝��Z5��{���۝t��˜/z�� 3S
K&��w[:�3�ʸ�cx�df�eӣ��QP[���K��eM?�Gp�4�t���$s��)$����S��p/2 d�º�q����ag�̌����)\Kl�����xۮ��@���)��/���a���z����*N��C-��x��鳙�۵�Eh��޻���!p�������]W�����~��c�.���g5�fTT^n�)�]���+�0�M�$gG�c���|#Mvm9��M�qwԲ:��=��'.�$���'i��=�6@Cz����d���i1�%^5�t�<94߻�+�{������HA�}#|Â���3�NmT��A��>ŬJ}�k��_<�W�×�;f}��ӣ�S�":��������&�g�~eBg|y��wtP:(χ?�ήv�7�U�v�{�i�
4ig�ǚF�̲��xID@O2���o	�|ce/��Gj'���}�Қ���9�]���y�\�$! �1�im.��q�+:*�]�R�5Q�pD�[�cz�bE�ff��OF�ΔcqE�Y�X���u�g�Ṷ��������ugjͩ�rS���ݓ�a�G2�%����e�����~���ml�� �Aa�ѩ��^\f�Z������#��]�5;��+і�/��;ᅊ�+��u#���K0I��,���G[��s;�2�������w8�}�A�EJH�o�\TK�Y�W����*A~���-6�d���H<��y�Q�ޓPyUx�d���5=�O��Uv��� ����-|z��ؑ���EPrMW��#��`�q�Y���i<c����戹1Z8G�z<7a#~nH�n�>H�����s��	'ʏk��|�5#Npm�S���r�}lm�Wŷ�J�Ҹ����'
ỗǃ5������.�۸�K�VK�]0�:��_%U�������HxW��SM��y�;��˦��/SϏ7C�@s��=�RM��ҳ4��u�i��u\O%��T�uf�2�9��m���|h�����CjpZ�u-�[W
/"�d�,"��m����ڻ�i�)��Ś4�X�x�)&C"m��҄4)J�Qy	*v޻�.�����Y���;�h��܍O13��z�C�*P�I1U�'X�Z��X(���fh�\�^�Jg��`�DmO�2uw��l�ˁ=�@[?���]�=F���{��)N��6z��o��U���f�^�nF�����pLy���<�v���vs���i�j6g�P��4��[���@!�g �P2��SMWJ�I%�5 �n084o�;���Tjk��|��>b��9Άt�E�uF�o��p��:�3��1ә�����^�����A%����|�1B�=%#f����!^�W�NI��:�Ϥ�[^�v��'&��S�}v��$E:�u�<�gK|Rw��m��t�M�o�z{���*��u��Z��7햁�"g�r!�\�]kL�����y�t�8U{& �w$��~��q�+v���s*��ICMs֗p�А�gu�Y7!�ȉ��Q�7����Pʅck��Z�k-]�]1͕Dm1��q\a��!(��"E���t�<��|�R@;��ު���ʪ�0�vy6�����qV�"�rO��Q��}�j�{x�o=�q��޵*���6�9cv5݃��
Ow9�4� ��ov��2f�"2�RSN"�4�<q"��k��Oei�R�r��Y�p)�B����g��-t�?�k�}���/@�k�R5�P�����ʳ'�'4u�'p�f��jx_Y~��g���~-_��2�:�.���r2��S���"6����U��ml��.�������v}֗{K#)�r})��@y;{�D�j����u�F;����@���6�|i���s������mL��f$^x�q�f#�ʐ��#�ܖ�Y�n����@v�@��Xu�OYC4���K��oyp� 8�\e���UжG>,�T��TF�3��6�ӑ��쨁�#c��ށ����홀�+�K��q�����Ӌ�M��>�0��,45���:��Ǟ��.�r�3~}y��v����։��|�$H$<�bN��~x�g��%�Mq�����ҵ6����=��ؠ2U�]��a��UzЮE�V�|��U�C{��u����,�����=5dn�H�l�LZ0�--���,����.�a��Q1[�2D��4P���PNG����HF��ܴ�3f��:���n�3u5TDU<ѳFٻn�~<F�7��XD���b�`ű9������Q[� ��r���D�,N4�L�~��F�Uix�;/r4�$W!��4�%�<��D�TD{��Z��&��d��ȑ\z����²n5����wݽ�Z�f��������fڠ{2E�:�^AT
�[��}�޸[��ֵ�7]��o;�wpĬ�)]�ڨ��U���@�w�/b
^��o�:��	Na���d;�I3���0��cʒII�ǘ�:�0{��5�E����;�wl���r�]7����I\O�d�<��*	��XD�<�p�=��g�4z��w\7l��/��n��+�V�`,���j�o,�N%���p��p��l�&j���}}�_���U���^ �[Ol8mo2�9�X�
ex˝���C6<�t/�O�_ݍ�g��+Kx)�x�>f���>���F�����0�3�Fi��>����ߑ��?����~"��/�J�����Z$ͧ��%ꡦn*��ږʌJ������'y���I��O�J{̹X�oj����L�ؗ�'TƓJԇn�	����c���"��ՙ(�'\8����L�]YV�o!�ew�3�>�uJ˛�V�'˦gw��*����z[Y��`�TX����/����z�7�5�,�9u���R�؁�Z�¸�B��-�k����4��,���O5�o��M�k)�?U�$Mf��e���p㤖�C:q������ѧ2mY���x��f(��`Qha�<r��V��̴�;�ǅw�D��x�˸*��jU����u��c�u:XPy
0�hצj���#�7n�*�q�/_�f�QJ��b�s�Y&u[�,�X/�	5Tu�3g�����2H]��r����op�����ǌO�z���@���W�O���i�`�Ӽ������زo��XJ<(��+ŧ|{2zi����T��Fi�f��鄇YZv[JF�c�W$�y�ӈT+H��O!xF�e�t�^?n%�=y�����e��� ��݂��䊰�^���. ����*��E�}k�L��D �6�z�i-�yvl�gs���
/��·KM�S��R���3T���egK�2�8P����
ct}�`�wkǳ�3Wk5�J�ᨥ�acZ�7FxǏr�gL�
��ad�O�|zu�X��4��;����8К�36��N�U��v��Ԏ�
�*�>�C鎄��9��&�H�66̪ţ�J�Y��F�|��M��>���9W�;W �a.�Y/�t��!e�95p�χj�0��v�;Е�5仧�K�Pϸ�a�F�y?/6�蕲��ڿ�־����ſ^�J�Rw�qU��q��P��*=�/c��3L�S��F���j�'���W7�H��nS]A�yv����z|}d&�T�\�[�"�Oӕ�ѝϾ�:�a��E]��ƻf�����	�`F�_P��
���N�d�V�q��OS9+b��n$U�߰Wg�\.:��:�qV���<��K����Y��|7�c�A^\)#�l ���"��/#�Y���M=[f(˻��9{�k�>�Id�!�<v��Ȝ<�E���ɯ�D���؇��Ck���ц���|ו׷�MN���.���B��Me\��w��M�rݿ3�4��]�7,]�\{��ف��˅F���Q2R���r�L�.o�7;��U^o{������n�IF-����H�^^�s�N����8��~��UR�5����𠦕)K�������G�)��on˩�V�2�c'+�q*Ɉ�i(䕣��vkn���6��[����M�S�[:pɹH�XD�����}����l�bf�)�}��'L�R��҃�޷����@뤈�J���G�x���4v��B�L5��nQ�Uq\h������pEC�����l�4?�����|����fÇ�=�x��4��7J�?k���	[EO�A��e�E��,=�==�0K�EM�x���A�� ���'�OZ��ki���2�[mQ�s۱��p 9|� l;������b|�:$��6�L�k���e�nu՞�`cY�i��T���ȊO��>�ux��~�Ͻ�vM3�E��(�U�����t\��P�Nf��pG�{D�F�v�Y���:}0�p�ĂM�D>n�uc��g�#0�{*�4��n�}��lܮ��Nu��h�Ц��Ih��7b��.����<�x�Ltw;Y�
:��o6��l޼�:lGh�I�/��|8��ʶ��
�Ӄ�,�V$zku���:6FkՑVȚ�ܶm���9����k��x�="�����9��`>ّ\lm����p����~��=�����m�W�C[���|G���ˋJ�/2���3�af�r��|
��M��p��˜h��P�C��(~د>� J�n_cm��-G�qw�;K���6@>��r�$"�-��[n*^2Z{���*WI�ޱ�#!/)m��T����z� jHW/�(ڬv]�Qp_
��������{�>��>϶��qaw3
ɡs#Q	�]y��۵�;���i�&�y���Ӛ)��[�<5j�h����V8}�zۦ賑\r{A1÷�S�	U�Fd��N�� 	���M�h��}Ǝ�yǴ���7���b��-�n��J�A$��q���Gta��ʬ�t�����׽<+�z!�4S.�^�@�R��Ƽ�&@'�Q8P�{}:��D�dUz�X`�̏�U
l��m��z7U��B��3d��,\�gH�R�lsVi�V�V;��}A�����t�s��.t2�l�J�M*�F�t.��Z�o�Y�o6��ޕu��r�� ])Tجb��ju�d���n!DVMZs��.t�-w�,5b��3ƭ4�T�4���;�l��oK��vV���t���������g�==Bߪ��Q�+3N�El��JԞi��6�QՌY���[܄3a��\n#��\װ�{+�Ď�K^{���%_dwrw�jN�҃U���7�$��#�8�ba��(C��;��v�\���ἳ���Ε僺��vg`"o�t�n��0�@�k\ �6g+[ݑ<.��9B�f1��K���Q;�+�reu���}z���׉>�ʂK۸�^��6�Iş
�{�
�R��B�]m��6���=�UR��,�&��5Mq�pB��}N�Z7�c2�z)�1�a�N�m�~�,��1�X˭��,B���F��]W�/�� s�˚*U�V��f��S�5DI��rpӜ������U�;�:~y.R�2@e܊�������P?��A�����F���?No�B�̋0,ʳ̫0,ȳ(�H��̋0,³"̋2���,ȳ̫0�³*̣00,��0�ȳ*�2�ȳ(� L!̫0,ȳ�2�³̣!*̋0,��"�2,ʳ�!"̣2,��(̋00,³"�"̣0,ȳ�0,ʳ"̫2�ȳ�2,��
̋2,°�*̋0,��̣22���"���������3̋2���� L�2,4��� L�2x�9�fU�FaY�a�`Y�f�F`Y�f�eY�a��dY�fE�eY�fE�aX`fE�`Y�f� �`Y�fE��e�	�	�f�`Y�f !��F`Y�	�f�V`Y�fU�FF``e�f� �F`Y�	�a�I�f �P���9BBUB0�*a�!�@!�!�@!�U�y*���x��0�0 2 2�0�2 0 2��ʪå� ª� C
�  ��2��ʪ�*�9�� � � ª�*������Ȱ���p,0,2,2�0,2�2,0���<�������ʰ��Ȱ�������0�p,ȳ�0,���(�2��������}����*0� ��	�pJ�ᖫy���$|��>����
j��O)^�II��R��0�*���r��`� �w1
�
��`�D����@�ևj� ����/��kjHj;������%������V+�l 
����*� R�@�J�!��+*�@Ȃ�! B2��H�� �H�
��, !"�  +
�"J��@ *��(	�B��m"C����bz(��("P 
	�C�*��_HD�;`�=��p@ddwVO���~���i�M�k;nJ�S� U�lC�m�խ-�TWR� ����pa�ZL�PD� �j�@���@d�'�Ƀ��������0������i�> ��V0:̍f�=2�j����Ȫ@SuŅ0�S#"wP1`t'�pw��-�* 
�.Б���T@u�]�2���"Ky^�Q� �9�:��[������	??��Q U������*I�Lm��=u.�IK�AW� �k� �+(���o���$�i�����)��� �����8(���1"]�OS�U	"*R���T$D�T���U$JB���T�R�TH�P���֠IQ>�R�$��UT�$�R�\�[���X�1�U���ڥ[5���3dٴ�f�lY��Z�W�v*��-�Xm&�CfҬ�Z�l�m�d5��M�w\ųm)����i��=��z�a��a+*V̦�m�)[m�(�*��*�*ֶ*��m��4BəmehҶ��cT�-��)k*�H�5���ʦf٭,Y��%��ݶ�YKm�M��  \��������ףm�]�MT��N�th�z���M��[W�ޣA��S������\���Q�y��N�[=��U���b�{ս��KNn�s��N�W{�mj	���b�,m�֫f�  	�>�
JC�Z[���D�CveJ$nW���U(P�B�
��^��HP���Ω��n ��gN���{�9N�O{nkͽm��n�nJJ��v��]��ݞ��ݩ��\-��n�n�mog9��V��+e[&�����   l��}�Y���b�rd�w�S�5����;c�ܧ5��=+k�ޞ����c��uz�{�ӣZ�ӇOZ�@{��%^�/]���^��l]ts=x�[@�+2U���Б��|   Z���e}��;=�N�]�v�{޴�VӮJ�=���{r��ݷ���m��[��o��׻y�Z5�y�꧲aM�8i�{w7^/S�٨��k6٨M�"Qe{�-��   7;����:����Ͳ��ٹ��+ն;�=�֭�//=�a��Q���:o]֛��햭1o{;ҽ��������^^�3�ƶ4=ƇV�m�%�5�[[o�   �{�����q��R�j���4{��Wf�z��YU���ޜ-k�0�Zog�[d&{�o�<�x�U:�FY����{k��m�ki����ub&R>   ���O�fe�7�mY���F��hky�����y�(S��<w�  �{.4 -v�  ��  ����E���Zڦ�-�5��6[V�  �� q�@  �����g. � �@ �+@ ��  �J��@ 9�� \� F�md�[SMjj�D���  �� Z�p����r� Q:�  ��  hwW8: 
6v�  v�  �� ��ޮ� :�mb�Z-f�m�f�&��w�  ��  �  ϸ��h6��� �]�
��y� :.�A�� �o  k�� �X O_ E? 2��#@4d �{FRT�� S�6LUR7�  �~%*H �� �7����R � Iꔉ3*�  �~w�~߻?�����/ţf��wL��^��!Eu��C�!]<�#�K���UW��}�Ѣ{��j�km�mV�kk��Uk[o��U�m��j�kl��m�������y����� q��G��rhGq����ܷV����N��d��l�_2݄(SH�l-�e���X�.��z���Yn�]�.4�%\o6�V�.���k���I�Ֆ�j�{�2� �kP��υ^�yovI;1ô�#,��gg�0濎pq6q�R���0ܨp��!�q��z�5�^=8�l�Z��y��\�^�t�����I	�"�1�(�ސ"NC�����ҳ6)S��ދ���u�k/Z)n��i����u�r��R(0$&A�t$盖�m�g-B�X�n�͢�ZK/oD�%
�(Kd�V&Vk&��bW:��g�p@�
@����
�b�A(�Q6��7�)Y������	t��Y�^,6A1�HG���޷�v������ć�i�Y%��8�X���"�#(��8�gkt�LcHͥ�ҥ/5�A�&�(;qk�n,O(����Ih; j�IY��$�u!��Y�WF��e҇1Zb�n
����4X*3
���A����+v��x4ʈ�h�2jY`�K˃>�,Z�;r�5K3�J	՝NX���6Z2<"<�[�����W���C#&��{V`��z���
5���sM����{�jDŻʵ���V�b�g�{fGH*6�Vn�>��F��،�q��c˺�����Wm2C%��
!n�MF�%�o�%��qV3N�IS��\�w��ۘ��ǻj��)������G�k �6J��QE��bţ,S2��K��#2�����hK�d�N3t�	�e-N����w@��mnc���CX��u}�mG&Xd�tsV�֠!(��V�h�����\aX�7�14.�a^���4�f�Xp�E�eޣ�KҼÚ"08�ڝ#t�FLlK���Eڕ`�����ƶށ�]��T����@�F����.���S݅�� ��)�.=L#uik��བ�YLȦ��ɒ��`���.ܷOZ�~���'E��)57U]��q�M���f�[�Y���Xa쌜�zZTf43�$Yv.H�O2Y��)�f����U�B6+�;jMu.�KnI�%k���]B��������.5U�i鵗v�f�6ѡ��d�4J��ډ(ܠ����n|�D��Z��d����\z����&Z90ִ��m钛��},��ֿ�˧�%�b2���Xb��GS#U�@ڊԤ�/���
��]Ԗ� n�cvZVU�SA�v�ѩp�N쐋�mh)�"��d]=�Pe�nmղ0��3����1���H�9�2V���ǥ] /\�Q0KI�B�"P�]آ�1@���b��s楪)��ۄJ���`��3+b6�;1�כ-���e����*��Ҭ���̛oCX�ݳ���f*9a��n�q���T��h��6r�.��v�e� XI��,�2��h�[SW+vjN�ڒ^���L�pRb��܏^���Q]������3�jeDȥ���(MsY�n��ܧ���*��Gl��_ؓ/p��7��j��`M�u�`Ҵ�V�	�횹,/S"� �7i�M+�qk�U�.�cFn�OCV�0�b�6�Ba���l�tP��5`�Jj�0X��Nlw(��)��������DZO-�N�%�c*ّjE^d�#S��
�6�ei.��}S�iѷ;���L����X��;�wE�� p-MՖ�;n�#!s*�L����{�N%[@Z�|��F,�pm��M#R��OD���Ŏ�4^Ѥ��HoPɂ���fd�X2�B��YI����&�z�k�X4�:�`�٪:ԭ���֞�Ų�JB���i��Iz�K�c�1���t�����Y�d9�Z*ə��42ŕ��.��2n�7Y��C+���%nK%�%%z5-Ү�Y�nF�1ol�Z��]ފD4�uuH^PE�e�7�Gx²�f� ���x�L��n6��,-�Q����t��f|)�Q��V�S�ˆZ
����ɖ�
Waq�j�c9������)i7�5vh�+Y��y*	3%�S[�N����vj��з-��)K
df����VI+fhQ�	Q���7���ь%Z�qT�N��PôBYkv5�C�)��e�"M���(� 4��a�kp'g ��M]��Y ��q�)(�׏Z(��^�*�m��.��/+�(�cqJ��k�kSݣWb��j={l�k6g��[�Z+uq4A��iջq�I�B�Q�bM'T�E��k����m��#Y���/���M����޸�A�^����A�7޴ʂ���7R:��
yOu��f���+3v����S��S��m�{�/2�+�ma�䒶(��ϋSk'D�8���gA4I	�<;T�'�0S�]GXUT>ُ�k�7�Q�R��*�|�ՙE�fVBK4�?�PB�����#S+-��Q�H�5-N��m�b�C@�3�Tp�V+������*i\��6v�8Y�U�Yf�ݩF7�fl��EBQ0�
Uut��)��bm-|�X��S�Le��=5x�rZ�,�Ic�V@�k�u���Vm�,&����K�o!^Uo� .���X�S 	{(n��#N���@����pЬʍ��3R4J֨��^�+V�?
*��T�ix���j
Ķ��2��r�A��w�6�R�pf �� \�Cu̈S�1�-3�p���2��Ǜ�f-�<xw2�%(rñQ��e)v�&ƞ'�-@�$}E�%��%����o`�j/1�{v��>�4�jA*I�,jn�\ŪS�i��Z�+`2!bCv �n��c_
��@YˑT�Jh5/^���������AMC��c����@V���n���Ł��U%N��!t��8�l�5&$��ˠZ�1��F�:��w�֌s4�OI2�y667>I@3K�����o6��k��Q,�Ԋ��fe�C%�c�H��.�ME �&�����ɗ���bD��Lu�2&tQ���zcv-���{�R���"�䪵m,0R$��v��N���Vr���#�*�4P�Mi�5�>O2ؚ�ZHh!i^�㵄 ���.���q�)��wGqϜE�l�Ð̔Uј��ifLɬSq���G@��b�Δ!��wYcd�����
��Ѡq�'+i&��""\m;����4��g>���/^Z���e^�wP	4nF�]i���х�ۋ�v4�����P�ZlJZjfD��͗�kJ]JQ�ҝ��<DkUxq�eDor��q�R��TP�E�gZK���!qah`7��S-QR����Q(��%a�u�,!SY��X�R�M3p��qS�S4���PL�+>�նB���C�#�L��se����@�8cSF0��7Q�"@�mf��!�2��c��S�š+����t�Nf�E��q۔�r7�-��P[X ���kJZt ��dy��Be7C�h��T�����Ұ��t�Y�6�s^^�c(��<L8s��d�%�,̻N5N1Y�M˛Ni[B�=����]�4�eR�Lx,;b��2��E
���2�$CHC�ښ�)At�����M�e�	�t�l�V2�wo5�u�p�d2�t�S�0\Y6�(�X~�Ga�]=ڲ�L��V�*�T$�o~B�`��j�Z��- �I��Xu�K���V��.���-i	���[7i�V�SS_,�I7��QJ	R�$ܗ��v�kV��+b)c{��@�tK�`� �swP�1U� &�"�Z��^�3f�1�`����)x$˭�<X��4�ç�!@2�.\MU����e���C�����2D_@�`Q�ߡS 3]�:�٠�:c+R�"��T-�{PNZ�m��+���XOה�R:r�(5n�Qf�os.2nEÑ�Z6�=����T��B�N,��w��h�	�)�Q&�u`�m&��]J"�ղV����A<�ϩ�6�R�ڞ����K��u!��-�a��b�V!Ǖ�`.���j�46���b/�h]m��Z���^jʉ�[�<Ă�P��5���.�:��@�ؖ�i�ճ�J@���Q�#Ыe�i�ˆ���*Q�I�e�D*��:�Z��!b���#���F��b�W�����/"t�s��`܉5�x�5a��8�vFf��^�2��wh8,�����U����׀ԥb7���zwt�ɺs5�����Ҥ�m��GU��$&>Q�2S��ֱfй�n�5v��M:��=̺f�����<���j�&�)�
�`��2��ƶ���koB�q<�2	�0��X�cp����	JV��2�DM5#�L�oJh�4�t<Xի,��K�{k
[�ؖ�*��m����fM�*�ɻV�S2`I�̠o.�{��`D���H���Lڵ���oh��Q�G�J�n��P���h 0,��1����1�0ku�Zw�M���؍%��o36��nk��J(mm�L�1G�5q��ʴ-F��ۈ�����ll�h2�c�Z3(���6����]�J�J9v�A��n���A����7^�� T�n�x�fM8�m�1Y̵ P��6U4$(����d�"s�7z�6K�<�p�޲���o-�Q�N�%2��i��~��cFfiz�$��0Y�gl�LP^Z�J����m�.'��*�OC�[I�믬�d�\ְBmؾo"���N�,0m�Bdݽ�>���1r�X�����O"�/U��R�\
k�حJݨuRłS5��s/B�i �ҕ��֫+cF���H �����'r�S��'>��h�'k� �\�LZ�PbX�^ϳ��ש5nG*��Uv��Č[�[�X-Ǔ)+w.V��٦��l�\���L.T�wj�3l��ѣ�cc�C�+�0ѥ�[&�!Y�ںDar$P�f؈��a��&c�#��>R�;.�Mnm5@��͙(5�y��H���VN��aD]Ke�0���qJaL�jHM��[�h��B���(Df]���3w��S�t������������n�w`gKf�K���p�Uz񗑥+.�}�E`ZM*v��Ǵi']���޷��	�pmX����k4CH��vAq� "�E�n֪;RQ�hTVSج�Hc��Wj���-�n=㢶*�+�#֭w���]bjZB�0@�.a&U��jD�z����a��LҚm��aM#%J��f-�T�Vju2�������SIF�Vfۢ�m݆�ҕ�ycU��fc]٫Ij�PtV�:�y�)ud�y�,�V̵i:D^���6/ _6Љ�|��0�Z8�
Q�0<cop��Ιz��(���Ձ#�sskVe��6KL�ܫ����
E��:M�	�e�< =)ո���N��F�TvR۷��+H��%wW)�rA�y@L�f�<��5vYl��Ɛ��"��b��ȴ
:������+%^1��Yn�Fd��`tRV!
%���!uF�"�'�����-Uɐ�e�;y�������Ȍ���̌\�CYV�2����z�e�nV��0��fn`��[� Y�Xp�u�iD��۶�`/#��dA"��ME����S,C��B�t���$Hh���u�>xׅӤI�������<�1��6�*��RԬ�{�b�Y�,Z2B1#l�f੡P4��wN,�Y�FPǴF�j2*��n�1^A��iRƨn�܁*�6�z�iP���-;F�1.�Xi'��îH���[����oP�2Vؕ��1���^J�Z,hS���%Ӆ8�<���t'�块!֛�v�KE�52Y4�)�{)��H����8�ڥX쩘��9s6]d�.��hS�Ab�)V��X�q����sE�p���ܦ\����;�� �0ɠ74
�kne�BՋ���ܳz#fR'+�m��1(��i_�#��t�VsѡY@�����f%�%��lhT�T�	�Y��NQԱpt�l0�S���.^��b;zrd30S�HY�P�ǐ���ə���lx۬ڟ`��Y���2�\i�Y���R�┰)y�sD)N�ᠵ��汰
��Z�CV�n� ���s	�Ɂ:H�շ���^��e(-�WZ^��ћq����~�[Z�AB ��V�˵R�j�{���Q��hHH�&���6�/f��e6��T')��݁�S�m��5���jϠ0N���+�A��
�T�+�l�)Q�hݙ��]Zs�Aܺ�&�5���e]�hc�z��h+x�`�BP���E�pLĲX$YQZ(b�3c�.��(�7�X�)]�8��2�LE��y�J�(Y���f�������,l#t�m����O5�y����&QV)���\���
�%Rh-UҸ��4��Y;k���u7slvX5$�5�^\kLg���5r�[X�R ���hK�^��X2��-�ڷ�J�a�MIB�b�h��Uj�f��ַ��銶Aϥ]�Ւ��0m�4&
�Y���4���W!�{�dn�mD)�����2 4�m��:IP�`*�vhL�Yu���A�1M.��(*�&�b��+^F��n� �F-?xs���ӎ��@�u%���rV�y*:��8�N�6�/>�HoC�(���kq��/,f��&]�j���إ���dGn<t2˶'��eMe�gUN�jR�o^Rce�a�Y�$D�.��;X]cp�@bY���1��y	�Єa���H�2N���3F�KZ
�#4�i2�5ô�?���d��0�ESc�c٘���ea�%m���X.�t�3"ծP���$�kq�Ba�-6��	�4�ePn��`�=ɫ5	������C�W����kcwk'{�q�m�����{�k΀��8�cB�Ly!X�#���S�ȫ�F�Wz���s��W,+阧!��qS�r�f���Y��>���;]�]:�T��q��M�\UMy���µ�[d.��k1���tf��u����_��tb�F��.���j�B8q������;�޶�aA�m��\w�}�{�Fخ�۫Aw�N���R����o=k6�>Z������oT�g��gw��kk��� �$�кC�s:VfP�ݱ{�'���d<����W� в��:������X�n��Տ&Ԯ�@,>�'s��u��:�T��%����v�6��Y�B^��>s�a�(�B.���YO��}�TW�@��:�5��:��;��9��ʹ%�!�}5�J{Z�Mi�m4Wu�v�(���.�ޡ��>V�  I�����f��K�WgS������䫡�u�`k;��Vr�8	�8YS��P�~k��@�H���e���:ﳁ�{}ٱe��#jҘ ����Ԕ�)e�ˤ���4kW<,��AG���h�*=pr���˧���3�۬��cs/燡�L�u+���-'�r��|�훣�%K���pc-�)
ғ}�2vv�\�� �`K���W�ϝ�Ov뮽[{��&�r�z=���mM��AP��6��)q��b�0n�J�Gt�euʭ9�hq�Kl� �K�u���lM�G���SG�a��A��O�;MP���bG��]x���n<-��V�2tEc�?_��n;کTwN�딗R?���V����Ŷ��7�]����c��UV��q1r���e#2��wl՗J�� ջQE.�ߣ�*��>si�8m]��w�h�����ݱ��9�S�Eq˰�[�K|Ӛ���a�Ƅ�\{0�a.���	/Uz�ݳ������N�+�pZTrk�3Y�ͫ�5ԝڗP��攒p�LS:9���iF]N��{����o���
�Z���aѣ�w����/cZ|tX�,��oZ��'�BK|�>���w��Y紸8��p�)	^�셒 �r��u�no(W|�Zř�kO.��e=�8]5`N�d��c�s��(x�g�� ��"���#�g[	o�Nv��]�]�H�M|��\RШ�����o;-α���<)�I��d'R�NLל�+�^͚�����Q���wf�(A�)Td�X��~��廢]�zVzi9�]���Xm��U�aܫ�}��ݭV�\9�u޾���=�ɝ�6�}4��,��a�CLi�x8��z�Ƃ���T����2��Jȳs���i	Z(L�]�cWOm�+^Н,튇B2�-�b�i����ݷs��ܮ{]���&D/ʂ+�(oȎB�wm�r��tUN��2u���h�����;�FE��/0�V�q�B�8+|���Zs�,+'��8�Xo�V�刅���X�8e줷���F�s��k�e���HJ�66MN=틇)|-�#Tk|k��Ǭk�wk/q�3U�I9��8N��=�2񧧎f۹1&�%]L�Ц�u�Q|�`j*����\\�Z���%]P���i�`�[�|]۱$�C!��m�hC��Zk8i c{��)q�Jɸ�]T]^���|�������$K\��~�$��R/}��R�)7���R��)gV���	Ե�v���dJ"�&���B�̫�u�����7���K]O�ne������O�e'Y\J��E$�+�S�-u�^�ذ@;�^�-�����Y�S��cil˘�Y;qf�`������K
)q�wF��Hv�Ըm��X��
�"a� "ʋ�3u���}��dI�޽o�q�r��*k��p.�)6�:�bK�}e�$7hԷ͜�-�dr�c)�\��N��\�Յ��i��Y� r7����Xk�_)w���̙A���hU��֟k[]��t�aq�W���R���JS�DZ���xV֕�j%��_oB-������f��N�v��o�4$���Iޏ�P�}�7Z�O�֏2 �6�[FX�&��P�n_�X��ҭ��M�V�Kk���M�U�;=���+le9������OW�V�}��/7����Uէ���d["�-w!��h�p���v���n��_ Mvkx��'2�(�>gp`�Lg[�y3�}�͚ R�]�hE�@e�ʘ6��(o�k�؃�#K+8N�M��oz�qe��<�ď��WQ�q*m�FeX�C�.J�t��O�5�G�%+W�u�x�����q������QT��ݐ祧pCB�|�|T����Z5��(��3���n[��Ȧ��p.�=O��]j�8A˭�Ge��t��+$]Ccy�Gtfd�S����v�U�ҹrІ7z�{RK���
OeJ�3&j�KA�X#]b�v��i���t�� p��p�q��v(BW�u�CVJ!��|z�f٬ÃUqH���9M�Pߧ.Uu/&^N��a���=�=V����rI��c/4n������3��d�v>�������$g;���G��%��c��4�:�'��m�*m�w �˹�7M\�dL��%� ��C���(�x�V��S1]t�X�����Woh%!b���qks�Oq���	X-I$of|�pw۫�&M�N�I:�{4ގ��TX5��qrA�62�wnZ��e�2b�*X��p؋1��9��u��*�l�Ҝu�e!����zqA���b��k)���]v�Xn��W��@�-45�,Z�詐�h��;r��Z�s}�f�qYM��H�p4Yޮ�E�1d6�\U��b��ހ� rX�"v���"d�1ݱ��k�꼜~�W�Uf
�^�N��1t��u�1g��]1��%�g�yY��ni(S����j�=t���J�]�cRحGFP�Q�;�N����:<7�Du�;��{wۨ�	�n����sjsx9�<#��H��C��jw�
c���:�'n��U��[K���f��^+9"}�]2�ݞ�#���s�"���o���=K1�ؽ	e�x���E�N��<�q!vj�t��6��!^K��e�՞�ݸp��E�P�7���yV@��=�4���ԡ�4du�U�km��Ά,��32�2^r|S[`mǇc|�ڊ*&M4�.��v��~�D�u�5��t�E�%t:]N�qT��_i{3z�ڻLe^d�N���p�sl�ȸ�a�pͧ�5@���sb�l�']��k`Xy�q^�+��X�
�dN�V\�9�{���f9L��كִ�s�G)z[Ct�9s����Ճ_LZ�0+�����V]�;3zV�
��yǠm�l���C�ҭ�jh��5G}_�N0g�A3�9�u��Z@B�N�,�]��5�pNaՅ��ܱa�ͧZ;�8�c��Gm�H5_l�HΝB��.����9��P��2Z�9�Csr����t�����F�;%t�OT�{r-���=��6�W3�i�K�>���d�Yӝ��֧G�EL	�%��\��`�2��O���h`v���G��6���;b�p�4�ԍ�8E�F��=Siyc)�Ng۹p9�
�d�6g_MX�(�9B0�R�Q}t�i�dN����%�9/��L����{<������+�5v�J
=���y��E	)��x�����5��,xz�f}�{39J��x�{x��f�����H��zA3�!V�E.f�)��G+3G��]���n�˂	�����] [�S3bT��|�o7���+��ZLJ�̈́Wm�W-P�K���-QWm�|�T��o\��_�ӷ��4�8�v_I\��.��ۆ�G�$��k����],��=)I�,dX�50%�еΰ]�56�ۑB������_55�+��5tw�;rwnu�J<�~s���aVf�왽�up����7y�n�.�s3�0J^}�jL\酵�.�L�}{��ʹ�Z�����p�w��S&)@5B�\��p�*�t�
�� -��g�H��f���5J3J�+��2�;N����M.���(�
�W�Odܣa����ش������}-��u"�|��7�M�޲��F�p�F��;vke�x��������j(bq�3I�	tK�J���7���p����:�!�J����S-���=K�|�c��n��^������n��ݶ`�^�L�{o,��G�j�ޮ�U�<`�$��n�+(�o܇Tp��4�8��*�e�շy��B�i��ȇxT���G.�3�d����˂�I��2Rw_�25�S9}͞���`�~G��I�7��;��Xbs��md�(WL �C���}�z'�T]��c���ݡ�/ �~�FLD��/�}2И��VDgo���	�p��O�3�8�T�}�V{%�pW�Uh��!5�kF�g@�[��	Iʹvu�;���z�1��-�L+��DY�c��TaWR��A\��������D�w׈R��B�lM�o�a�H�U�t5�6ļ�R�^�4�x��I���`V�\p]Ñ:�+6�.�5++0<"G�Z��}82M9�qbޚ����W($��<����,���L�j"e�ѫ,V��T���J�\ދVS9n��,k����������qV�,[�v�� q��������ԇ5Nu��+NJM't�A���J=WAٞ7	��2�f༻<��b�%yN���`~# ����)�dx�w��]���i��F7޵.��t1»��U:�<Ŷ��[Ԉ8�ѣ����H^S?oB��Ի�'��מ���36��+������M�-�2/g*��� �ohq��0=���عw3Z)Gkp����ܜs)*r��'Uo1W��,��%h��!Ȫ �`o���N�v鲣
� �!�3��tK���;��5�Ue�/^
ª��.���JR�
����f���2�Iy��Jtg����{f�ܗ"��g�:��;�(/S���;r�MPTa�J�I}52koR�XSrC}α��V�뙠tKi(M�ֳ&�z��C�ɀ�Z���^�k��e�o(0*��ܬ�P=L��!K*v	���t�eu�M;틩č�ċ�>����S�V�f�o��Y�N�4�g�~�q�oGE������f��o5Ph�E�t�l�ź->��(l�hf�N��R��1ŒP�C�H7�o*��u�=W�P�`׀�Ǧo���n 2;�7�Owr�r!3r����M'ū��V��Ҡ&�^���ݻ��]�������i\�V��R���'S�=��a����?n;|bi��#1�V���T0�#cg+ű�U�)b,�r��i�Z���+���o�u�eK�b�5�nt�bm!��>wuv�D�;�-U�œ��J����篇$����Fi�4�ü4��d�jS��*���R�[�`=RqQلw�9���SU�����ժ�w��l}>օ�%r����a�X��Γ`w��B�y�7sn�� L�����k����-�T��f�S��ߩ*/m�<\�4�$<�_��M�\����Hn��B�>���g��6��֗����]��~�N��i��$2N�����՝��s�A1Y�<9�u3���0Z%jG-��M���.F�����N������T(�����ǳ]�x易6S |�	Q7Qk7u�j����4�h`	��v_>ޘ&��>���+�h+o�Ue��A�K���S�G��f�:����� ۖ�0{�{�3yu�d�7gu,5p�����J���}��b�}K�y��k��H�u �zk�κ�
�LF[Xk'��p��n1C��7�h�c`�l;{]֨ px[���٥�\�yK���l�'(�kL����췢�9-��*ܧwq�]4vYg��������&�4:m�rg.a����z�uJb�!&�f�aW�s��O�V���Zŵb����N]-�r�o��v����B�a�9Vi����."�Y��׌�����8���3�A�U��l{vm�H�� CS\�.�U�S��e��9\����DG ]wSfwM��<�۴e�J�!������f�D���Slr��3Upm!\))Z�o�fn6�a$7Ԑ39v'�`x��2p]�:6��n�d�ڋ��b �{X��_>�qs逋�!�;����t\�C�&�Ou�}�q���h��[F�K�~��-������e�E����ɤ�>T�
�9ܧ��� �e���",��5�q�f�m&%\�����q�|⫕�np���|:��6�W{�����t���o���&�&�^T�
�Z�C�����2�;� x�����[���4.�êhZ�u�%��I�p��<*��4>7��.�0�1E�/soֶ�K��նi�TS7�㼭鱡�@��7��oT]����~�=]��+0?bd��nznupFm����k���w¯���8^��f+[V7�U�:*uX�����4�O@^����=aG���+Q-Y�Xq]wXx,�R�N֓�ˁMu8v���+WHW.6�8��ɐ۱�:sJ�ǸM<�n�h(F���ȃ�W	��ҭ+����c���l�^�f�`�ދ0�E��_vU�;:w�Ҝ7�u�	���X��Z��`�!܋�,	�rĹϔ�غ�]�)V�k+nIn��m+�p���t0Z�u���:�I'�:חY���dT�Z����G+Us���Sy��Vd�σ�
)��(u(�/�>�`Q��Y9��s(>x^���-㻰�\Q�����}�B|�}�ۂ�tW��P(G{�m.��t��f��7=�z@��z��H$�.�ro��8��w��n�����i�#M�l[M�m�;��jڍrױ6 ���=܊��ҫG�"��W�G�DG�}���� ����]~�4}��~�^�n��,`���?��,M����vٝ��Kjd�#lg˥}.yFI{m�:IEh`��5;�PjwZl����]ٍ�$5tPÜ�v��W�����צ���/�+�&uqv�W��������֑��c�4���\�ۖΩ����t�_�Ax-Xb�q��4i]����|�_�&��������8� vqe��b��J�C7�aU�Z�{J�}��S0j�a͑��7��by�h�4S��JK�ғ�|B�@�n�J�]xsB��:J#�H�K�fk�K�uY(��o��[)�!PoC����һsyW�]�p�<i� /������c+y�1ىt�ү�"ԎA�[/z\�[��1��������B�N䌊���tlp�͐p����Jd�g1�aΆ��m�{
�d�jqɃnme.5*��*38���)ͮm "�$�l.Y�w�XZef�z/�wx��隟2ب�&��Հ��/�xu׻Z��6��*�N/�#(��� r{�d
�%:œD+;A�B�[҆A>D��RUtca�2�gEaa���d���}e�\Z����3R��n-�&K�zd�D�9���ݾ8ﰀ;��]�ٗ�G��6��H*Pu�i���i*hs�עyb���q^ޢ�g�71QB:��Y��R�F���d�#@�Be�Xh�#�Ƿ[�۪����թ&�o�ɼZJl`�j����F� ���X�.��!��8�(_A�����Y7WGW*ۻAT��]�?<��
�,��ͫr&��V�5 rfc(L����M�������-�(�:&ڼ�i	}ٴh+K^���y��z�a��D�۩%��ՑZC���e�7*o�$6�[��^�P"�o)�V�M����x933o���VU��u���C��B$p�������R�^��<�6�=�3L�����3�/2:VG$��/�g[��V;�t�lB�˲��Yz��Ɋ���SR^k�K��2��tb\��F�6�ˎ��]G��W�k��|V�v�N�������Bvr��-�j���Vf�XK�1���kG�����ߜ�-�^tkcɅ�eS!}q�*v�C�֟=����w���K�v�Cӷ�<�+	�{h��h��ch[�)��͸X�xOd��s�>�k 6�e�#������1q/֝�$t�Ȩ�,e�t`�=s�)�l��&�M�{�@���ǽ��L"�:�(Y�4'Sj�iyB�|�.�+LV����µ_qpz[ǋ���c��	�+7­:Y�Ƙf��#���� &::���B��[��C��Q��BƓ����11i\�If�.8��ՠ�n�J�o�Tp�g�"R��ýԶs�&�1f\*F;���]���;����t%�Z;�WK�E�Rt/x慹��Y<2�4�ûx�+��]�z���FL��ʶ6,�Q����|v+2�p��>͆�r��m.5��
B ]v@-�DN㇦t��,�4�ѣz�;;�k:�CX-�Zx{�vq�~�����uZIT�^q�C�)^��j�`�\�(�:8l��E��VA	/u+���9��^o^ovW:��;S�Po��4���	��یt�;��,݈���+r�&���k�����Ԋ
J(W5G�d@�{�Z.i���d�P���C��\3r0]X�W�nE��JZU�3 �B-TӾͼ�`�Q�L�-TʚHξA�"ӫʰgD�T;�Q������=���r��EC@{�S�T�K!n0g��Zt�mͧW&�7�6g-�$J�N�rk����r�1�����^��O`u,���BJ�D��oVNHc�^r���"�;�K�Ѭ�ݴ��2�h��'�{� %�Y�M̸��Ml����蔫mQ,��������Τ4S����ޛ���JT��u��А.�>swr�u:Է�>��v�d]ePc��b�u���P��v���U�ͨm��U1��������eu���@���5;�&��Z#&��6�ɕ0]:߷��N�e˖�=\0j��w<9�kd=�#��,e��:��^'% ����vֳ�_�֍�����U}شݢg�s��` �\��m\v���4��P��fb4#��Wu�����T��mk�k%AէO88Z>�������	�ةs��L�7`1+I���>W�V�;J�
w���(�WJ�<�`ǅ��5kn��<������>y�dؖ�u*u:`��@Q\P��e�p�x�p	�_�M��ӽ���8m�M�dG�֞�`��Մ|���μ��]�+۬)��}��6���I|�n�[���:��1ܼ;�<.�g<�Z�8�^#F��}�$�,fAN�,Z��Pӌ�6�̺�g��%{OG$���br���BK7��c^g'ʭN��W,�n��bu7��TE�l���,z�]}�,���u��KH�ϷhU���� ���*>4�V*���C�Zٞ!�2[F:7@��̍�Z'�4�D��.\,� �pL5�P�̝��; ȨV�+�I�/8u;����D!���N���O��T[����2	=#|��/n7/9I`��U���W�v�:9W@�@�d�B����^U�L�͇�a5��+P��f%�j��'Y��Er�6|����|r�`p�\��I�g	�3�b��0��~�;r�:Ջ�ʼ�R/U:���yvd��9��T�5����c^nFHUs�+e]��|b��t {��ٯ�}��{����ؐ��R2w^��f�������*�wU�GL��ƄM���A[������{� ���ں�QZz����f�2Gb��q���6� ��;�-�5Q�ݭ�
���dы���':X��Y��c"��VR�=Iv& �NL�4��)\�3��U� ��%��Z�ō��\z�U v�IFR�-��T*d���p�)���n�����T�9�]t܋�*U:��!EԷ�����:i�ʚN�����̊����q�'�Bo��
˩�0XYQL�����j-�^N4#���6މ��z��
h�6��4��2kD"�<8�H
���-n�uZ��9A�<��s�6l�ǝ�v�n��ƫ���'���+�ox'��ZC�k��ң�l�g2�.�	1�|iڿ���l�Ǹ�D�t����E�;j��akYf��2V;i��cUgu.>{BBڊ+u���.��'d;�s{��]͟f7\�3����L)��oxұ��̀��b�qWԫ+^\���
<v�^qN�K�+HB���r"�R��������R��h����m��n�1X	W3x&�T�GoE*V�[]w�^�]��n�\�s��d]�(G���@��y�����Ź��դ裨�[��o�g����=��lb����s�[׮ڢ�H��Ɠ4]^$�b� ;�ؗ����p�V�hH˝I��PR�ж�'�׊��<+{�Պ�`�_�ENKe�4�C0-uNA?
�p�:N�q8��^����h��FoJ���½�$,�oI�}�7���� Oq�5k;�SK�ha��9-%A�m�9#��n��r��jH���1{�k�e��cV���6� K����6X�Mg�3 �X/���pK��!;�WWY�`�#=�^w+�Q���i�L��Z��/�vj�I�9r7������ͻ/v�hͥ"5`Gx��Q/����������QR>���2fVf��c4��@X�U��*h#z�Y�G�yX�ΰc���Y�=�]�f�䕵k��[E��R^>���68�:Vv@��iA�9�Z��mM�e��o�[kb(K栂��pSuǯ�ǋs��.�N���1�9T��L��L�����s^+@�d�'EkX��
u,\1���iE��ح������TZ�f�Qd�d��.���&L�y�s��?Yv���Oy'��M6{5��{^øV?$��j������1�u��������\<@�w�fH!��W�S,����0����(0�}mi̖ѿ�A\{Q��#�0�ԡݵ&�
z{��Z�wIf1i�8T�6:��m�{P�F����N����ѳ�;�Cz��dU��@W�+Op�$��a���à<	�N�ٞ��2�&�Cr2��̫pꜭYU�۶�[��q�r���T��p��X�5�m�}R݌3,֍�N�W]Ӿ�/�{���V���j��河)|��f���z�*�#�Y�y��ՈqSm���e� uGy]8�|�reR����,kκ�O+��:#O�ttU���{p�i#�n�z�M��:�(�L|�nM�Y �����[�Z��̤7���s��+4y�(��{�8��Y�c�#.�h�R���G'u��o����t]�f��_o\��S4������T���˩t��:-��?hБб���Yy7A�Pޥfs�4���S�1��_]m͚��"P���/��#a�P�~'�H9Hs�~��%>��Ar��v�Ղ�W6z�Wvl��|[���;�F�	�-S�	�V���}�.\����׀��:D����0^V1�b�O]K�� ��n�&�
�g�����6]�ǁ�;0y�eL�&��M�i(U�P²���ݪ�vw	��k���g��wK4ħo�
��҅��b'��	��X�)��T��F-%b�WJ�Nޜ�K��q�zeKRly�6��p�k�쿓�\�4�]�`�_>˙e�_#��]S���=Íu>��$\߬v����f�EûRV������E$�vL
��l/*+�'y*�D�'����@f!���dc�)�}6�3�Ǘ�6�6��p{�̦x��*�S�e�ڲ�\�E�Z��0h&��G3�h'7Z{;��p��Z�b[�gn��ұ��̐���H�����ʷ����O��W�s�c)w�B�d��DN�n�[�1\r�`�-����Ό�����S�ʙ.����\s TyO���úxQW��d[u�����g�KrP��\�?`��=[���:'�dKn������o@��O+�462�㍞Gu�Y�K�@���D0w�3����؈�N�����_�6����������<����gl�ڔG�c����:����`��f	�W���t�����.n̡�2�B�)��;����U�Z����Z��š�U�4_#W�	O���ػ
ͱ;*��hKS����"�ܻ����D�x�έ`��\�˯�&��"�ֺ졬p�c"dk����4B�E�ύ��|e��y�̽�+tciЖf0Ч��e��{�9H'��i�b.[3��)GR���
M����m��3. r�i�\5���}'u].5>�-�'�2.tW0.�ﻴ�A���$,�̙�Ūt�ܔ����>��A0P����v_��=0ջ�UA��ݼo%��d[%�"���L�p�Lṝ�x�߉9%��<�ɠ�����.����Ǒ E�թ�_�u�W]�U����&%k�_�KN���5�W+4�vm�ht�.�Fru�Q��ܵYɅ�mR�\EI�-^Fw�z����M��5���R���k��!��w+Z�J.�${�4�q'p����#�&�Kܱ�t�lM���9>�oag��=�<N.9I�2�uZ�Loe�Q��医]
�`缻V��y1�9�vV�,��&�A�/f��)<�Gz����,;��n��e,�mkX�l����{I��&)�p:�F�Ļ�V��1�� t�Z4��x����z��a���sX�IH�3����.�`�)��\�K,���m[.�]�hX�3a��B�c�|�4QG��S��S�٥
��3�W�̺;V�d�Ү��Vu\�Ȼ5Lf*�/>��R�7:ER�����h��Jڨ��L\���9e5��;96����}:�X�Lּ���m�{d;�?r:���pq7{i��i^+^z�i�	�-(N�z��E��L��7��w°�g���v]AS��<ոL�U��.��1Z��1m@z�y�ScǗpN$	�)�[�[��=�$�K�e=����:�����jp���y�/S	4)`lp��K����Z�:Ӓf<�k��˱:?��e�X�j��(��Ņᥧg\�u��r;(Z���L�љ�G��B�_�2Z{UA{4��+NK츼������b}�cn�u�d����t֪�T�� 	ܫB*-�c4������m���]7.��f-sf�nP�`�A��U�b;��ӭ���JP�G�6��W;�sW[1byC�����������؝d���XL9ji��U�����ܬ'�OK���d�{�<T_U+J����-�����	�.����^�;A��;��K�^M���Qޅ��]��m��Lܞ����@��Fh�.ߋ�]y�_��!U#яC=6���gmd���/��Fd\�q�P�.��7�Co�8�NYn��:�e� )+jr��K�[�8��ٮ��l<q���7{���ĝ�J�����K�˷�]���r�v�lN�t���:�Պ���eYǌϻ-c)n��c�9:��-����4,���3}t�0LJ&4��B�t��gn�يo����x���=tX�6��8���
<�(�gp<���
j�V��O^j�����{x�D�X�U>�	{գ�Q�C׫��,C���F\I�۝���</4�%���_"x��S�ηJt�W+�c�q���z�i�,���-����v�M5�mgM����7T}��}�h��S@r�^g�Vui��k���Y4��|Q�Q�\k�E�����F�-Q��]�ωg7f�D��a#����G���?�A�ɐx��v4պ�uzfc��ͺ�n�j6��Ã:�S�g�]&�aQ�������gWIʎ D0�W�(zRuj|3C�yq��4�/i����+�r�;�>��!��~PY|�:�	��y�fu���S��x;c�i���=��۵��Ҭ;ũ�]K���1|�:�g`Y�ML�����u�W[P�|wP��e�ɝ���y\]�:���%3 ][2j�(����b٢��~Փ�B�v�f�5%�/ m>���۱�`tM6��69�Nf�����o��MJ�s*T7�%���^�9=��)=f���t�{�i/�T4,��hQ�L@	r�q�ۛ|�)����x'�s�1�-m�|1�ǃ���6�����J}ˁW��*�^ޫ��t$�ċ�e��0A��L���y	u��Cq{���Y�|��\hz�
hb����[�̕>�O2h:�ߞ���҃/���nխ���v�;�.4|�o_�2���b��E�_m) ,qo0
(�Y�ӥ[JLX0����\�"�6	�8��yf�c�^n���/`uv�eX�|+w']
S�������i9������).����Z4�i�x8�`��zaֈ��f2�' �*�pO�O1��s�;�d�<��4��t	��T/mn�o/0/IP�=��y���*|>P ;�s�n����h��.^wy�W5��E&�F���-':�f1N�Q!��wv蘓h�%�)wW#���j�;�� �Cn&st���� �PPN:�D���Y���"4m�N�7��.Gs��#���dc&��qIFS�:�E%K�����;�4Iir�\�:�sS���&4':��3r.g��0b�����.��#^.�v���h�q�s��t��W#<��y�;�����+��wqݼ^M��.���ˮ�]��s�y�y3���nnkƼO�����[��r��F��c�zW��oi<��8-p�e�obj������\��t3�5V_^nv�;5�Ҹ&�3�u�����kg]�����t�v��+����(HhyW"��Y�Q�u'�:h�! ��u9f^��qιI��Q��b���Ub�q���X��vs"�>�)^��Qе}�$�m���s�%��h1p�ݎ&oL1�;"O�ܱ}R��.:�KA�U+�uon�^�s����F����ޖX�/��@a��Գ\<�Z���D�_����R�mv#������K!��t���\�=��X��Z�-���p��:{�	�91@�P��}u�4x7��0X�
��h"-ޟ	K���{~L��}[ӎ�ԆC3��,�.,�-��~�$�_Abx�FڠχU"�crE}�y��t�u`�輾���cz�YcE����>ʑ�s��$s>=_h�#(i<}A����BVmu�=6k{1n��$F
��r�H�jX�[Z:P8M*〓���k��4�ׄ�e�TZ}�g�ñ;o{\Ǫ��ꁧk�5%�� h�5�T!�As��F�A��J8�'J���A���S�b@Ҙ
�3�F��c�����*z�v�
DN���O3��e뭗���|�칈dWٜ����4���������ڔۡ�,�U�ٰ�:��ݚ�t��i�u��Ν"}读7'^}]�J�DN��t�q�ۛt2��Rޘ�v�2��uSg��k�,p�ik���H����כ��Dx��m�/6dbVr��v�u� �ZH�[S��W��??dS��4�n}"l�e�f�L�5���aB}�[�iX����jz�����%k� �I5h2�	��ɥ=���G_�7��%Wy�Gz�N�9�񣦵���#	v?��{N9�>�c�y��!	��i�YݯW�������l� pb,UH��D� ���<���T6��jL�&W2K�6����l����8�)�%� kL���VIZ������6��ǳ���]%�ݾU��%��Ac���˅��ݲ3e}	�`�͒�͆f��a��:���d�]��Z0�Ww{�wݸ`b�=�֓�,1�h1���FDjt�������Y��n!��oޕ�X5<}�͂�3�su�SMA,`9}���a������1ڦ�i_l�}Sr�:�����j��yƄ�r�s%[e�s������0�����u����:U�)����1mb9����ASy�S{Ճ�ܭ��V���K�W�MaU�u3�ͤi��k}a�Z�M����Y��ΞB�s���]���W�Kw��H�,�&�uV{.)w��}��$�;oQx��%�:�,��8��u��ʘ�V_��s��Aډq������=͵�˾��ӎ�j��E��t�+���>1���pw����j���A,)��U����88��I�8��aV$�\��cU0m�^��2����!|uQ�$�g]�ai��O��$��!EC���3ԅ»���bD�t���t�c��|ڸ}�Uk1!O�n�Ei�8��Xf���B���:��f��zWN�\*�0\5�ч���s��"�����\'WD֨NI�C��()�t�f�|��c��D��M9n�Mv��q�r�a/��5L�(������1�Jt�iy�$B�KxW�
<�j�ٔ���q��kx�8#Q9��ns@��b���'��k��@O�x��=�^�Nd����Y��n�,j5>�%�!g/!�*�$R�����Ճ'�`w�_6�,[�r���� �SM��Y��!���(�J�^�����,�Ab�LB=����Q����(�$5Bn�?@g����f>�w�1e����Q���7Wrs[c�i�2檸*���z�T�0pở���"Ǐ$ι�����<,x�C!x�L�Z�-ٛ��+hӾ�ν�-VT��l�'��K�mmnG���w]Sk�XS�������c�J�vy�CWU|��wr,&C���Ms�(�%�n/u�I��s�Cq�a>b�IA���b@�9�^��p�ݚCH����b/�N�2:'6F�����4�P�l�4���B�Y�m�0o�9��;~�Ub�v��;�
�V2E�Y�Z5���\G*B9�;�=q�np�s]Dt�1C�eد�ڷX��*g�H�fdOy7�����r�'&�.ru��Ŭ����a���D�)���{~��Bmƺ�R4���EBS̰e��.�=��Q��a���ԙ��{5�Է'��,m��B�Y�u2�l����������"�NS=�N�4_՚8٣�QZҜ�JlЀ!�K�3Ԅ��bd�	B�v!F�X�[�����#-�i���_hj�o�E�Ne �d�P�J�1��
⌤{��%��>��� �J��i�3��)9��F�腦��Hۄ��v��Hzj$�
�*�B������:5��N���c62��G��J�<�k.
.�
�]<���F����":�����ͯ[�����=.�G.�D8N�}n%���#�U8��.^;��ZL{�w�����(�O��~��_Oj���í�';�Ӣ�Tz��@je����1�aC\zH�x_�J>dT/a�Z4�Ft��d���NWL����Ov���q�Z~x)r��-�3"�u�e��J4�H�U�"F0c�i�I\��������,+�S���C�e�c%_��о�ΓӸh7���E�N���Aq�	F��b��rj�W��A���bឣ�JY-3,hu�E���8�V�R1ѡ�t��Bӟ�t����6n#6���-��ԛ1��Ź"p��]QdҼ��Ձ�����4����A��N�{c�š��[�΃��{��:��kE��X��ű�Ue�\�]��n�rn##m��^��b8L�p�Zϻp�{�Y��wyR�|��p��)L�u��ੇ�q8�(�w^�f�"��iD�Q���ȳ��F+���sq$��Х���^A F�޻�:�Cʨb��y������e\��5@�iC�������3��c�#��P�vB��A�mm��D[�>�s�;o�ׄ2�P0��(y^�Y�1R���,RW�s��˷9�k��J��g{^�eM�wL���kUg����H�7=q{=�#�N��2�p�n�� ����n�X_Ce.!�p9��3e4�9˰M��7�F���%���#��X7qX�]h,����'����f�%.3�����0x�)rT��(��rS�����
��y{\`�m`��X�p�^��lHc6I�������D>:!@(�uTp�:��>K)67�\�9��B.�&`�,oD��"�i}�'%�*��u��iq���Sw3KU��u���%���Ƥ��ƈc9�\ �_|�( p�PAj3p_}���E=��Z�T�,���T�ϝ��j!�0_Ж�H��I҆3�u���5g蹖��>�S���\X��A��EG���̎2�W�]p�N���L�9d��e�g��]�z��]И�T~�������׫I>�F�4;�5	Z�4WГV�.Q1G��8����eK�����՞��gX�A�4�#Gd�����\r�k�;xLf����^*+j^�6ɽ3K���ؖ �ЌX�o�u���P#�]_*=�Å����� 4��x��5�G���z>g���!}]	�I��
^���M}���f�
uC�o�E��qԳ�W�:x�p�&�E�P��!uI�-��lm��g���^�W����>��s��f!�K�nBWk��v�8�̎�Z7*�v��u+n�%�8�����r�0�U�{�j��P��T�gM�WӲ�>Fj,��ޒt�]�6��5hV|t-4���ruZc���\�<v���̀��Xl2=����ܶo������P�E�#�瓾ZH��eqh�b�>����##]|:��M5R�Ov�S����w{(�x��~P.�=��zh�0��@
���1p���[��(��=IR@����X�Ny�}ͯ��j�v��`��(���2�x���� *��g���J���	����`:l�E��{�]�{,�1��#	~�����Z���n�	ǧ�q��'P�jfq,�o+2n`k%��D��{��ݹ�;��u�w�{D��x:�3�r] s4J��W)>/�w�]0��	1KU|��`�|�/�7=���f��z_x����C�V$n��������J�]+�Vgk��܂h��rv���:C2�gk�������~�u�՜1ZNoM�1�Lzy��P�$YS�ULK�V���R�ki��N9��x�_�U=�xN� �h�C��E�>��a@�)V�d�+3�k���ӕ��Z/�,�į
���+�<��P�j�!O���<0��n�}�w��D���
C��T_�lRԾ0�k��)��v.�_u��{�4qRaX�Vé�K��x6RY��09�U^�if����S����F�L�S�6��Y�Yx����eIK:�8��mRM�ق6��!4�J�� b~|JU���� B�s����^��G:����fuI�oO"�s:!��v���|��T�(TuJF�& !3�m*��3��	�k����2Q�o��77����ܛnc�19�d�F�
�6�
�8Pp�}�J�l�9ݶ�����})�`�cB���K���Rb�N̛����B�mL4MR�\�T	��U�߻���������eJ�SC���뿐��;�!��7,@Η��n�(/r���UeB�{�&b�:�,a��'t�Q.sQB��,MULA���kK��-3��ף-�X#�O*a�
vt�u@��a�u�׸�j
���S/����=�6���:���Ad���!����{�|:�u��p}��~�|kV�������6������L�bg�Ԝ0�Dd.����aŬ߂�3�9G_«����=�zWt:�39fO}n&]��P0�8J�3ƥt/���}/x�Ӟ:[6
�`�K���S���yQ�m��!ۺ�nh�D�i�+���%��/�\kw��p��S-*�t�Z��^��O"͟�q��ʋ�^̯��v�.Y����8�in5�3�)s��f����ۻ*�-�p	�㳚-L��a���W�L�up����1Γ�u�^���U��>c�]Ll���c�
�Ϊu���3��h��x���N�M��i�4b���*����s���U\5�я����<�9B\�&��9=�{m���3�`��[/�����F�ё��-�B�yv��=��-���]c��l�\'%�ײC��fF$��w�6J� 騉(F��	xw3T��,3j��=�y��e�
԰��-�����ӟIG��2]{/�j���)}[Da֐�)9�Ǌ�:�z�r�wރ�������烔��ڜrU�BH�l���Ğ41f���U}��>��Ò&J�4.)�1��XW�m|�[c����1�����`��S����1���@��/�BK��*;�E}w\ȫ�ޗY�����}�S%�ٙ�{��9��ͺKC�S5��dU���DR�>'(v}n��y��na��ڄ#�<�1T�zv�ƺ�[��$��h=�\"�+�健�3B��π{c���Xng���s�?kWk���ZmQ�Gj������p�j�MM�d�j]_W<t��C&��u�!`�_L�`��%YO��%4X�2�C<P��S��+QWιөe:�ƙL@5v#�2=r�+�ot▶����`f>�}�d��Ԁ0�V�1������uyuo4������<7L�x�sS���4��on��7������L�|q�%o�K���{��5�C�r��D� �l<�@��3JF,5��
�*�7��ң)�6:|ճ��,:M���9����Ҽ*זB�H���9o���=��|r�̾��
���+>���l���i�t�va|��m��D[�>�=�_�A��tnK��z�U|���p������d�f~�$�E�㴤���A��ܐ�&�5�E�����y�cgw'�)����ᖻ'϶�*,$�h�����P
:ú����k������]J�Q�VD0���&b�c�%m�X�:	;Q2����m�f��b[����sۛ�,����"�	�\��h�^�D1�:����^D�����l\U���T;.M�{��L|9h4g��T��v��,p�ik���Rp�����x�N����7r�T\t��u�:`zH���ә�P��xh�5\3�X�n��}JՇr_@���v/��۶���H�7ۖ�F�.����֯3MA�siL�G-k��� ��z����TC��[�Q�3#UKaa��������|�U�و.y��K�,�����)p&V®gL��=��v��qn4�S��L�
�E��x�Vh�4�Ыid+�bT�XK9p�u�	r��L
r��!��ƧU�^��X����ᠯ��/�]�j���]���^o`����!|�Q�l����y�#��
�w�I��)R��p����	v��X-��[��0Y�0���x�Mb]�^�F�����T�V�*Lł��J��P9�F��
��<.Fi�s�9n3�F��`)� 3k^��k�;��H.�=���w��=���.�ہ�9�_k�N�Յ�ݾ&eL�cP��}ӹ��ƮKn���Z�e<`l!T%��Ի��τh_B����%4�[����� �91s�����Dؼ�}P�����}чI�MW>ΧApy��E��.:�|V�G��f�ic2��>jf��2�Ա�2F���aB�L�Bl�έߔ�)=����k�Ų���c'TU��Ʀ=έ�Z�
�Z���e�K�Ŧ���ڈwuݒϽ:7s�r�T���i�3�!|~1�tqp5Џ����������`T������V���_N[mY�{nl�yf�{#��3T�Ù5e���P�3��R�t,��}�^PR�\u8'Y��<Җ*]bhʇE^I��O�M���M�z�����ۆm�:�m.�d��39<q���WJ�vR���dධnY���"��S3K��)����mӔ1�z�+�g:pۣG�@�y.;:>�־Tt��F��޵n��b��H�QR�v�5�F���ݵC��iO�YE��>T��7ԣr���U�,�M�g#$mWNx�!��K*�]��g	�y�ݳD'�DTjlC(�������C']x�.{�����5L'{~�aGG4*޽	������]��*3�Ք����@�h�sV�.�pi5�E��(�I���=���/�v[̼�3}[E��UpWx�L`&��q^gr}�t����hq5gg�� �M�{m��W}Y�$�gC�Ɋ��;.���6h��)�&��uf���]��h+����aޢRT�{;Lɳ7��I\�g} �Ԩ#����3��1��&ޝm*
�	KV�.��,m~���y>�������J?s&�c��Xh���E�N�K��=0�ɩ��R�Ke&�N;�F��5���t۔���vQ���ܙZ�^�aɐB��w
�Ν��s��6 �11�P�u-s��Ȓ�Ԭ��/v�T=t���Ww5V�:��\�.�*4;�`���꬛�x۽fē�Sc/�.���v��z��.���)<�eԻǴ١A�mx	
�c���ё�O��u>��S��ڻ�ؾ�RX	Z�G+�Yb$��\�v�v��v=�ڰ@��h�#�9��r�nUr�wk�E㤧�˛�wXۖ�(�s��r�x׏�;�s��^yˎۦ�gv�p��E����s���7
��v����Ƽ��].U����8G+��7s�s0���\M���t�wa��[�C]κ�H����sW7]ܹ�I��x��ws�72C�ċ�$s�wtk��D\��u�wu�wT�u�x���u-�y�C��t���^(ӻ9ۙH�Wv�\���u�.w1�[�7;�W����9��#^0��+���;����2�����K�K��t�w���t�m.��r�� �K����㝐wݹ;��*9t;+�s�x���:;��/urH�����8N�;��D��%�.�s\qĪ F�4QI$H�w-j�,��2��L�W����֑��9G���1���8���U�T1�wwLM{E��&����;c�[2�8��������գzk��k��Z����\��Žo�;�77��{������ţ�z���m����^+��[�~��o����+���_~o�ߞ�͹W���|~��c�}�u�}�s�~���U��Ԏ��+�������[�\�m�����V�7��wo��|^֍�sN�|x��k��x5��ǿ:�m�ε����/ֽ��{^-�\��^/������@��秱��f�����J�K��姾����~�/x�����7�n�վ}��k}W76������*-�W.oWίo:�7����ү�4i�v�-�}^7/ּ�~y�������#]G���2�'X����׶�������x�}��M�_��~}����W��k��ߞ���+���|��η�x�zm����6����r�}��yok{W+��?�z?ݷ�żo_��i�m��/~w����@�����5T��mwoG���ۖ�>����m�o������~����~<~�����H�Y_h���F��_��x����^�"���{���޾������/�|���o��W��x�{o=u�ȉtW�W��f�}Xg��c��D`�����w^��i�~]ס�͹W�����o���6�������o��/~�|ץ�+�[w�/=��o����[}~�ţ��y���<c7����{�w�_��=|��?]�yY��{�ԣ��P}�5�Ϸ޿��k����/�o���{�Š�9���Z|���c��6�]�_7�n��_߾ož+��w����߶��U��m���ֹ�QM.�o�x�7���zs�װ��]U+��}���/M�-�_�����ֿ��5���������������7�x�+�_���/KF���x��_[⽭�^��W����ί>u�����g�U�AAAφy<1��S��ǟR��^���+���Ϟ����|^-����������^�>���6���t�/�k����nj�<*���c� ��!_~ �}¨�gW�����{�:�߫�ѿ������DH�!����/P��R�_u�-���������j���77��y�չ�����>v���}�~�������_[wο7�|��x�����/�<���6����/K�����mߗ��W���^ם����<"�G���5���W��n�yp�;]Y�+|�U������C��=ɴ��+0�����.�;��v*.�g��Z�Њ>>��.��'*S��>kE�ٵ7���
,^َiyr|�/�A}����^koW�_�8�o�M=����$��8��gǏ(��m*���=��c�#�>�Y����<"�} c�����u�<c{�?~����o����꽷���j���ּ_V�^>��^7��׋�}������o�Ϟn��W�^ٔb���}�}zs��4�߷�������Z��������o;���SF���WҲG��!���U1�|�o�������r������|�E|m�^���!��1�+3���H���ظu�����o�x�_{��\��r�}�y���^/U��_5�z��/��o�\���ս>6�^5�~y��kO]���<���*����o���ۛ����^���c��Êo��WN�>�M��>��K~<[�}��^O޵����w��+�ţ}�u���}W�{+�7<Z|����||[�����~o:�G��菱�F���G��}�}돐��@������&WY�=oo:��p��6濼���/�߯���ν-��~��y����ץ�W?W���k�ε��������zU�������o��w_[r�^y�ϝ^���y�+���k��eoԁûW�y��ħ�y�}We��׋��ߞ���h�wϿ}[��_�o��^o_�\��}m���U~�m�m�u�}���ߋ+�������ֹo��z^�x��Z���m�*���<�ƍ͹n����}�"}���x�$��%���1��G�B��Z)
��Ú��L}«��*��:�x�o�{�����o��^5}��-��[�}����^/�v�*�.k�y��F>�D}" ۘ��	}�$}����ɜ��Y�u�������DP��"�_{���͹W�z���6�noM����5�Q��H����1�	�D5ꈹ1����y��׍{oKţ���ƾ�ƼzW���}�ޕ_���v������z�u|<���37���y�X��P��"=��x�<���?��hߪ�wo?�ߊ�i�}�6�7��7��ߚ�����^7���h��s����/kE��ϗ�Ͼ���c�#�/���O�xP��)��w����#z�1~����$��$G���}�������W��ۼ��[���k����w�zZ7�����^_��W�E���ս?���_�ߞk�ήX����~�y~*���G��1�c�
�>g(�^ڵ���� �:֫X�0�s^e��~��-��]fS���u��R��_��֕�=KQI��èԶȕ|���+�&P��C)A/=GJd�fQ�CG�C��np雝���K#!y��e�n��Ȟ`���i;<w��9I�ݒZ��(��dz���]H��H8��c��k�������so瞺���|����^?��ϞW���+��^���צ�k����o���_���~u�o�|o/�~�KF���}����x۽v�k�"��D�}�e��T�{ۯ}����4c��_~�����⯫��o^z��__��-���>y{Wո��|^}����i�~��~/m�m�|�:�^��77�^�޽-�]�m�o{�5x���x�~u�^��k�����0��A/1{o��{�>�>b$}_|������^>+�����Cb*�k�B#}�ﶝW�>C�>����"z��7��m��_~�|W���W����{��+�_�t���o�6�{�ʾ�K��䏶�y}vvE.�+7���}��#�"�����K��[�x������ֹ��ߗ������^�����zo��������7��*�|�祿��x�[w�z��zo��^/���o��F�_����7��W�x���ы��:�.eQ}�.;��}b>"G��"F�wl�ur���{��W���׽�y��o��~{��o_{����ߛ⽮m��η��|�M�*�~]����F�͹�_��5����Ƹo�������x�>�}��u�=o���Vr�Պ��f>�>���8��~�������om�+ƿ?;^r�oׯ;�:�U�y����گ�����K���ƞ�ҼWո��~����W�ߊ���w��[}_��؏���r8]_�{�SY�wup]���#`m����W��W~������?��[��ϝ��z��\��5�|^6�noּ^5���yޖ�b/;���^->v�׾�oM��oͿ������Z7��������i�#g�9�u�,�G�")h/�=|�����^-��W�u�����}�������o׏��������+���������^?x��ڽ��Mͻ�o����U��wW�u������g�6�	�8��]�ǻh{�#�f"G��}����=�����������������ּ_��W��5�ח�����U��}��ׯ:�c�{��}m�����7��������o��/���sQ��ݢ�\���C���s��vg�3uzoxz>��}�}��^��4n[���o��x�Ƃ ϔ�D1D��|�>�c�#�"6���⾫��i��<��~������_}yW���w߾}W�������׵����""�X&)O���]���]�a��Sܡ�`66����۲��cpf»�F�P;��"h؝�1d����B��4�6l�	{��;��Z�љ�ѯ���\�x���/]κ�v�Aq|�#c�#���K����k2\��Kj񇡪�A�89����{��\����m�}�{{W�x�{^����oʼ]��6�^��nzm�y6��ߏ��x��w�m������|j�G�����O�|��G�#�ߌ��G�>���H`C��	���[NG/]���h6'߾W��^֞�{��xޛ��o������h�>v�.���[���w�<�[w޷�xߞ�o>u����7BSb"�#�����}���A�U��"@D��׹�u߶k������������^�o��<ޛ�n���������m���}zcxۅ~_ݯ��W���wv��Z���Z���/����{�����k�_���~�y�C}[��z_���0G��">V��鎯d�fnW��M��|U����>����oM�[��y��ssn�ܫ�߾z[�soן{�v��nW��__�4nW����o���_��wx5�_��������7��k�__X���$}��I�ᨯ-�^�����޼�^�H����}����� �DA~Ο�DX��3c~����N���7hxF��T68�fpC�~7,t��]І�'=��3�;���=Ng��߯�;0�qZ�ߣ��q���h���:��+|���6Ւ2|FzW����b a7�W{���'����>�Y��䣠�-qIWoFZtU��F���mi�ƀ�tUpB���q;!r �7��w��y�4���kt��|�W��Y3⇻�e�����F|nٮ��iu��թ
���B�pڃsr�s�E��(�,ꝝ;#��}u{`������hd�,$�h���:F��᡾)C�תRy�C��j�R{$�Jٍ�<AQ�tp̡(5%_�
^����%ZY�2��EA��R��V������᪋��~�4��sp.A80K�����{Agv̮D�;{X�=�n�,;��YI��aXY� v�+�M�'�Q�Pfnk�L���=�ӊ�fP�����Ϡh�_�n1q-S���,�p������@D�6��>:�*�w�/���N"�Y��`�_"�	������,�9D1��θB�.q���(�\Қ��&)��K�����,	,Y��U&qۯ���0_�k���Rt�����u�̋����\'WDֈ�.N��U��I�<�s�B:���!�W���h��R��K�AV��(iȊ�8vbuTN�<~���"U�&9�2#C���P��0R�6��:��%����3�����p��%I����a����������w^덪��\��p�L5ۙ)����>�*59�OCn��3L�ьL�o��5�و63��"|�t˜@ν���h�L�	<��5DZ)�'�t<f�o�NGL#�9�dۖ��%eq�ۮ6�3D8�_�U�~X����wݥs����]�6�;��az���u��'����Ӛ�Ic,��,�v@��� �Ã�N���Ѱ����a?����5{#3s=�i�P�JWST�
�@��ţQ��:�V�p;�80UϢμ�R����Vi�/M��}�>}
�9ue���ׯ�VT��]�Gn��-�.n�<��5������tU۹�U���O;z��O�@J�.��J�{�����p�_Y��Vl׊�@� l�Ͻ�a#]�ad�nnN L�!(*ȷ}�!��Y���cӵ�E�6�
��ߵlhI������:QXe.�;��]�!C�D.M��IG;"�B���s�"�g������9?j~����AO��Xk�;Q�ٶ�ǵ�SǙ������CF��
�)eꇗ�
��M�q��Sf�� T�y��{^Sr����I�([�L��S/�:��1����ƺ`ۘ�6ܦT�_o3�{�LWs �|��^�+�Y�?"�XEpt���$kLة��ޞOh��~0�߳98���l�����J�j��v�O��p\p����C��Wi��:^�t����,e5
k8
tz�����>�}�D�u.Ġ�p��剃�F���QU��xL�wǯ��Gl�� ,�1in����铙�+�.�>;��M��`��uHM)�������
U���w�ŠZ����{���k�p��}I:H���s���n�lAϔ�(WT�Z�0n�B�F�g2�:*���T���K�b�/4��	��9q"���1��Z':v0�X�X���=;s�{%�cxQ��Xo�s�l�n�:`���=s�ֵ�a�uQ�+N]���Aԉk y���Z҅�w̋�:�����6�]sZ^=�es�Tb辡�]��*U�6 cY�u��T�ci.�&ۘ����q�МyN$yςV�����}�d
�>��V�m`�SH����b�V��:!���TB��f�����U����ߧ%�%�� �Va�{̖,������hg����x��?�d���{�!ƗVi��x�����[��-6D̷��P�����M�y�&���A���$9�^�o�^�;N�;��ok�%Ug��UHE�7A����T�&��Lʠ`�2�c���}�'m^{̭��r�i�W�֭�<��m���d<&Ҧ!����Ш��,0����z@��u�4����捿\
%�ʮ�x�HGbeu''Q�:�v��ldg��c�ټ[@�h��F��%�O}�-m�}��ӂ�*�i@$6�����`���2���f��qwR���DID�ԷY��+j�6p58Gub�(eL���"�L��*�
��*Bh�IN�-��e��\��mw��d/�<U��{k��B�+_	M-�*�gºWN�Wi�)���^�9y��Y�`���l��x1�Vl	��oc0����fU��G*D�C&��rV����4�w�y��o��:i��fs��p���NX�����-�)Yq������A�� ��)�W/h������둺���S�6���!�׌o���S���h�ɉ�2��n!��鿥epY$��2Oh5�#ё��.��)	*�olU�<]��3=�V<�W�J�0�&���!鿞�H��;���d�� �!�'*��7uc��X���j�P�?��:�<�A@j�'�$����r2�գH�Dn�k�q4���z���#��@/��
g�_\j�p�U.B3�6��C<��V��^;�m�m�G�hק�Tp��T|�||��� �e�p��ڗS/��VYK��y(��EW��s�v�ʗIx�7+�C�B�i\�J	V��i����{M-������k����f�0��̬S�����>[\K�e��"(��'�������;�>�O����U�_�2�#�e\U��x��o}axn;[��NWF������;?	��N�����8��n5����H���$q���p�>�1��n�_Г�Ӛ� ��a��m��b�ٜ�p�V(ܮ$mMa]���,O|<�������Wx����Ty	�wAY���=cP�>�\�q}��痯�%6�
Y/v�`�f��/�v��['��vj�ur�4�u��L��]3��������8O��
Xo*`�G�����vs䁿�r~�Z����=�uc�XӖ�{��	/����<q�c�=5�K;�����p�otr��}���/�y6���0���aL�
�r��x�s�P��q.���ʕ���B���k}Y�*�+�ݐ�|jd���$��������q;0�`x\	��|�(�����υ��߃�Iȧ_f��=��Sƃ%.���0<��X�3�w���*��Y\�ru�sRF3�ί�S�.�1��|�m���'|�����g��tiy�ڮصm�}}��B�������s��@�<��	�-K�+o��	��`,r�S���{K��d5wﯻj�f�0Y�E
�S��Ԗ_��םP�8˫���qW� �ѹI-���h��N�#���%?_]Rg>v�騇,p�%��;IҢhos�v�Y�{�v��h��U�دJ/�k��<���\u���C�'��N��:�O"�֩�7֧FY�˧t���t��K?P�=ƀg���z��B�M���e����ٜ����f̘C��[�D�a�Z��q51����ؼ�ъ�i*=�+�p�d�uZҴd�{֯x�R���X�on��f��4�k- [.Yeԡ�<��=^i�u�0`Vo��м.y�D����ʤ�[�ۻY�هN�#b�ge!B�N�+To����3]8�X#/H�:�-�����;1����Y��}�Gܯ4�5�޹��V�|��r�a�ڝ8f���1�)�S1 &z�TR��)뜼��.��2�`��CQ�7���Oo��5DTZ�ɓp۠9�3T6�R j��*4�\*�9���'^^+�^�����6��?;}�����{\u�[޻d`+�M��L9N�܇Z�}Ϊ�5Յ���7�"�_�c��ε�
)�_���7�5S��R���3�Y�)e�����c\%_�w�����@�g�{*�B��W�߀�V�3�vk�����l�=/�+P��Ÿ�߇�:�裔1�^�sc_e*�+�;��U�Y�?��+6n�EĶ����e�n���D�/�.'�Cd�"��}''�a�O��Q�F��U�m{w_%7]U_3��2ve:J�@wi��<�%�S̾ط0����WVt�oB��b�Y�g[�ֻ�;�,� XN��_Llu�b�Z��p5���^�J�{>R_�a`�R�-���}�#���ϼ|(�<DtV������ۺt�!d�	���c���t�?�,�d%��V�Y�CM�}O�T�N�PѵK�B`��[
��˂e��l�OQ��R�\�	o�uA�\�5���x�N1{����#��{�c��u�yF,�n������B���)jB��oh������5� ɶ��˻��@�P�[�xU��0Yy�yZ�ږ:*m�xaݼ/�[�j	�Y�3OI�@�����Έu�J����W�,��x�B�Im~����i��b$/W�������+�w.��j������YU,��N������C������R\g�ڥ`Y��v����Ww��v!8��.y1�U���a<�W0��L���{"�^�`���T>���紃\�ܿW��h<�䒭��u|{Y��J���;C�<4FR�K��0�6��E�J�:��yj��Z�޼�m��Pa0���YN�Ų`�؊B�����4Գe<�(�\T��e"��j��Č�/�%f��N��)<��NzZ0�3��ʻa��<�#�w�-]���H�b��G���h(�$!���#�Os��M�ξ����w��2�J�a,���;nn�C���j�R����嚜q^TwJ����7��kY���v�t[`��f9|�t��\�fZf΂`��W$_��'�z冀z��H�ğo7�	r�,�^���2�mB,��{f��{2�u͜ޒZ"u��[�B���k"i�"��$2��ti�9�����aG,B�<m����3p�n�S�X��j��0пx�v��B��uqqdy�����S$�m��G��T˧��������oS%.�@v�X9iڱ|��b-��*'h��FGX����a��Me�rs�vZ����,�^,9�4���X^�2�vED�����x�����*\l��2c�4,�nK���^��/GlwYԑ�Gd�Wv��]�te�\(�}B�����wc�k)�{5�.�fr�C-4A��w�0d�CHS6��_%���h���	�%�T��09�h�:е�)Q�9N�9���V�=*H������H�����@[���h��[a��=
ӹ^��v����_�i˓�0��u��ں��N��php5����[|뙱����yp[�Y꽵]ahl^���Hޫ����rЗ��!Ílђ�*�:�0cbTgID���z��YF�ez�Yë���R�HZB��fE��ܞO���0�3���'��~�u�/��=�n&��E���e�t6 [M�9�ݔ@���m�������M�	sea%��8���*��,/:�q��@�Sj�M�Q,����}k�G�%�$��i��|1�֤�#�X������Ks�b�\9�h�iy]��b�����[�D�h%�rm6˻������h�4��,\���.��'����l��t�w:f�9����fKAs£P��y�B2�4�K���<�#��l�k�%+𧫞�����+�1��H�N����%��"9�F5�;��:	�v�`�ܘuԑ��N]/<����wu"A��.�ٹ���ǎ#�pԝ�L�i���u㗍7]�r��ˀWws]#8��.r��L��RF.ww7)�Ɲ��us��.]u��r�,y痊�y�D�ˎ���SH��c�[������y�x��)����S�y�'�����%;����1˦�p��Q�K��M ������u���wF�.t�t����R&h1$+�.��9���v��JR�;��p�Msww���d��ʺ\��uB���x��)9��wD��n�7�x�(��&���<^D��sG$wrL�t�F9��M�1\�n���.M)9vF���Ƽ6!���:�NE�w\����L���ww8��n묚�r��ߝ��׵��j���A�=����J�%��u���L�|�F.Y�um�t���Ʒm�;��6��O�~'���G��d}�-K�ܜ��feF���Y�ňA$��Ep
��$:>U�el���N�c��B�ꋺ�ɼh>���A�{M��p���84����$�C��
��U��'�/n��{9�uyOj�Q�W�e��R����Q�ߤ]�L��b]�]2T�q #�L�N��i�Y��qP�@���=�$C�KxW�	:H�pCeC���w�[�g�2J�\_v��ѕ�o]�Z:�E) ct�������)���m%��c�0��2^#Z3s��^�o�Ɵ���~�9C�hfW�ܬ��Qe���aZ���Ra$��/��Z����o�����U�J(`�Y�q�K@{+�^2�<�_�)�'���n�ר߱ ҭ�Ȭ����]��?�Dt�D',j9��^T�Q�����N����s�P�ϣ�w@��+'<{ڳ�O��Ӫb19�bB���!��+�x�t�c��9n�e���ۛ��煥�w|�51�0v�f�P�1�wPz�����.�|���z�&��ދ����|�����!���5�m:3Eq�g5YyYՋy]��3BMO]B��On�n�4��&�:Bi����k���u�u4.���mݧ��v:K�d���kq�.jK�G��kض�l;B���oi�qNK­�e�A@�:�	�JY� ���+�諭���%��ޯw3$?������[��ô�Ў����"2'/���rz��9�ķ���������`A��n�_kK���=��8��U�Y]�|X2�3�	��[1*���ㆬUO-ޚ�a�p�^��+�t
��|�𧴨"���]| N`F] �����n�hޑ�b)H�E:��A��0��Q� F�*�!u3�o�TX��ĉ��L#
x�S����u2�'5z1�c�9���*��d�k�x���?A�>0�t�);�o'��s���6�.�WU��ȩvv��k�!��{�#n���6J���7�Ì�,}�ͥ��w�
je߽>��	<��e�ΰ���}T'�����@L�^ȩqK���2�N�v��Fm;�b�A��!�Ha��W��xE�\j�p��S��`9��ƕX��qO�$�f>�MwY�s4�{�jR~�����G��DW?�"#����_�%<>�K��7	��h�N�(��VM�v��H�`�D�f��T�&�ʓ�A*�O��4F#r.�JV�������E���ޙ���ie�~�2mo�ef-^
����}<$�a�8���>R�|N��]�2�t__�}z2y&%�:�մn���W��
��z��׽ó7 ����:3���u���u�ng��3�wZ�]׀���z
7����?o�}UU�UQ���=�,ܹ���MS%�X��PDpD�D!i9K:j�@j�����-��[<�g����p�>wL'�R\a`+�健�3Co���&#����J�"~2����cݼ��+�.*�;u��U�w��y���*_�͇���P��z����zy�_^T���_c�G�sc���u��;���=Ba�ta��1�{N��yAgj��h�!X`�_���L`�|2p+����|'�'/���d?eE�'����/;Q���Y&Jɐ�#=����<�V��h	QU�P�i����4�#-�sK�\m�S�K�����
o�>�о
/�Mɩ���S7e�����!�Cs��\S�Ag�ժv�9�UA��������yN��������e�q���f!%�o�+��_91���;��w s���a彸L��-S���(L%�k��d�YW��>��4m̰&:�T�0��\�E$J�OK��!�Z��[\��q��_��O����ly�Ə:Z$Vj�L4i�8b7�#�����
�egS�U��/��G-�ҹEZ��(4�Y��]���Ш0ಞΡt��?<�Ug}�<5�tOb��I�5:v>���٫Z5đn]8R��un��qʋ�g_���}_U(���=l��������%0:x�?_�uI�N~��,p�ik���8՚�Vu`!��׉��s�8:��_*�b���}�@�q ��EA<�s>�2�R�\8v�J�U���ɩ[K/Z�t�����wq]�񿄳���"Ut���]F�hy��.���u$�V5���0tM8�� hM�A9t�����ɯ��}�d�Ha�� �L�����(��z)%�=�@�ԇ���^��r�d�Cn��� p�F0	UH�3�회�c9K9j�s�o�d��_�����6�U�	��q�+�O+��`��2Q����w�c	%`Qhos���{���C�I����ͬ�h���?E�����y�C���df�� �̫��i�6��.���gX>��Y��b����Vr�X���<8:��1���&��ە=S��Dd�"�v��j4�\?�*�T��\�^*����1�6j�}쪰�������CȔ��
�,�Յ��{�2�r�B�9s��T��g9��s�}_?�Ƅ�j�9�⫬�>��-�j�鞋|�� �FU���lj�}}Y�1Q�K��u��jGv �]�ǎЎ���Co��l�P��Umǈ����_����3�'���Չ���-�(ޥ��a�v<$�g+�3�O��`Bip�K_��ʲ�M[�?*W�3��d�Rg�z""#�N�|��]�6�L�D�|&81ؕ�q<�'���U�Fy첦<�<�n�e��՗��E��e��񨄰�&m��l�A���%#̽V��|b�Z�AL��j���r�V�Q�|\w�����  ��b�_L\u�b�Z��c]0o�0x[)���0e�u�ͫ���5b�~�pb5㢏��A�����p�k�+$~|��E	��k�>�M,����a�Ks_�"�ŵ08�Bj��S����!(�'�
��HgʻL�/P��eh���73�s�jY�3;���T��p��F2!��.Ġ�p��,L��F�P��,) �Q��jg^s�s�'��2�⾞Blv����X�;%?i3>�!(��>� c��nm��3i-�Z��p��2��y�$Bⷄ��:H�9���s���6s���_�bz�6{4��w��$�$��0�$xEIZpfDi���7���K�ɸnc�1ng.�m�qc��Vָ��J��%\'�]����|5�k�x ��R�uv��},ʢ52ax���;���]�Ԟ�*�H�noYD��sr�Ⱥ֒8wr#x�?]��I�3�̢��߰�8�XC몌/��Om��o��N΢��>������:��X8��'$��&y˶q�Ț�����[*KТ��;��z�^�D}}�\�%�z�i��:e�0�)�%�쯵f*WT`��T�֘C3>�:!�t:ƭ��R�y6s�;�܋��[,y�,�����B�v��Η�٨��ͻ�i��	�J�`xj�	L���P��+]Ɛ�k�
��ˠ`�(Vݫ���{�it��Q���|ܥt�0�Q�}l`!�)K�\�����F�>�^�O�<�.�%��btF��@�-6
�	��O#�2������9}�%�c9��x!g��t�ܴ�~|
p��F͓�K����/3bQ|��ò�Wj�Jy�3e�,9sѐ]n��R�nNm�T����1zp5��#���p�$�#~��Ad5q��}{�����������;�w��]J~������<U��xm|~�hk�j���֗Q��d�n���,M��wق���� jw�	�2�{D=n�xJ����QC�+`��L���nX��/��0�Q��b˸�bV��
U<8Ԗc^�͙Ϋ���ɣХ^��=��p����VĖ>��66�ER�8=��	V�Y/r+o�o�>��yq�3�����O z�Y��^ݪ�==�Ty�ܭΙH���T7�.t�WE�؏��{��m�������9Ϻ���j�Rs�������������f�14���	 m��#������ι����`uP�zrJ"�ׯ�K� �Aw{so�v�O�A��TL����|*L����.4���d*vٌ�se��c.W�wv��|�w7F,C��Q:�Q��(�RD*��A�hgԦˎ2¿���j;���V-�i�'�܁͙��VY�c%_��ХLM�k��UvF|(���s"�;!�3�-�yM��T1�vB�Q��T�y�2��D`	�Q; ��;�V�4o��jR�ٵ�����D?eL����&���a`*������/�*g����J�lF�����B�m�LX\Fܾ-��Ɗ��lBI�a�:ɸ�A����5/�9�ꩍ�k�����Y�X+�Q��`���(�.V��N��y֯�*aᄜN3�1yc�.�;�t�5]̓)D����3�#�����`d�W�NQ���d��v��Z�wW��'v�{Z��!����'N�՝��N�os�Fm�N��`ʃ0��|Pt�ve�Y=[��vxE'j���k@�5(5ڻo�\je	дv#�R��+���0e�Ȯ����!��nI�:�$Ӣ`)s�����g����E�Z��W:UFÏ�v���!��.x�f|iS��n����2�����vp	ͭ��NΪ��㧻���PD��}���ї}�M-nz���V����|3�t�Y�:�4��÷���J\g��p	�ܐvMv��y�Ņ����鐄p��G��P򘎹u��ȕ��B쩷��C��~ɁRէ���o�����}_I���L(Z��`�ON@�<�{p�����ȕ��V^F���/��{�s1TH�a�$�*�ޡ��C�Uq�/�`�P�&�r��>�!��4CةF�-����q��o^S���/�`(�( p�Pǁ��iO�uI�N~�[�b�"̨�<���s�V�P{��¸8���aQD��t7���ZH�M�(B��æ�FNvj}ijk�:d��_6sK��wp��O�,����{�z��_S���a���{����N�kQ�ێ5�>�E$ա�]"a���m� �;����~H�G
 σ%�=����o���."�3�}���
��0��m���i�8Z1�J�@�l4�'���v�m^]sF�L���~f�oƃgh�t�6����UU�L�6۠9��3M.��B ��n���Q��/�u}�0w̃p;t	Ғ8x��Mz���h���4Te"8�[����AFep���q�6vk�����j
��E�왻�R3J2�	k�Ó8���Uq�ݬ.��^J3YCv�^C��7���#菾����M�3��M��c	2�8���"�XuS�~��[lVAд���[��񊺵�ƱZ�U���_Z����K���V��d������Y��B��^A^�=�
)�_�<*��P�Q�8����UY<88�K�5�c���^;�`�[�c�n��VƷ+�^���L�t��޾��ۚ�4��*/UCT��;�r� �/k8>������Ρ���U�zj�/��Eڊ]�C?z%�!S3�Od	� ��Jȹ�P�9�b2:�''�nj~�u�F�j-9ζ��ݧ�_��r��F�	.K�D	Ń��+�JG�z���¸���mD��S<���;����=��Z:'�&�t)%��u�b�Z��t�f.�L����u���`�լN��d/l��>��zxh��>x�8�+�T�pikѕR�J�$���"X�mu򽆵t�h����n!�v�W��g�b�ㄝep
��C>U�j!ypmԇ�{e���ֺn�����B��R���h�>�������p�If�Ѽ(y��qy]|��1RQ9�ʹ�z¼�Ruٍ[��]����>]�� F��@���K�Y��ʛhm�C�m�JwvaG�����iu/���em9|��ܕ`��E��-���g�Bog�9���3{J�꼓.cT��°d��W>��z���+�}�}�}�ov]Ǐb��'�2�8���lv���|�)��熒�{0F��'�S�`��l}�+q���{��8À��ⶐ0�}���D-�_RN�9gD6s�;X���{{�i�Tvim�|��4 �(��=�Q4㢈�0K�
���j�w(ؒ��(�vUU3Y�k\�]v���ix��G3F��}�r�$U�;L_t�7��o��n��``κ����U���Q��4z2?����0�)�%�=���DE��z�r�WK��{aq�HL�w��rso��'m��-7w"�d9�� ��8>���H:Y=W9x��ԥ�PgplJ�l���l捫-ܱ���CE�,\%T�\bt���ǖ)����M!V8����*��aOCJ��vBɎVSDI�c#�S7���P�1�u�{/�tǭ@�����ŝT��}�T��W��(��VUiҩ�x���Gb4�ׅ���8V���͏9��U8R\�Y�
pՇ�F�ϒ�tO�>K���������CxR����X�&�_7�5���U�l���xSKk*��ޣ8.�E��[B�	Rl×ֶRo��R�2ݮO7�B��V��� g+��k����K�K��ͲE!3���+)��:����(�_O!#z�v�&E���ۯ;\w\���BJb�4Vb���|]�	9�w�Jڡ��`�s�jو,����pC������7��Rp����*m��X�*�k�z��Q�.e-{h,�fz���c�oI)�$��$V펣I�t��Ք��k<��J�W��J��������W���)���B�+���j�c�Bu�N�����Ck�����@��X���mj?oX��Hr9d�"`kxA���t7��^�{��7��M��UU�.�n0@��8���C자{"�dz�pyT��V	t����Y'�疺�����WV�[��B��ۘ��V9�wo����l�.�K��&��\����5�����ɓ҂\7Ԋ|k�'hڵH
�֖�\��WR���Dqb�`b*ߞ_r�Ygu
�	W$�+�kU^���ž8�vk��+L�ә���Eg8.�j�4���Vnk�<JD�'+�������l�|k�E#Y	�;>��h}VV1G�#^�奈��+z������ ��U-ٺ��u qU�V���k(�\o$��щ��0�s��"�7��{6��O���T0cj�ܮt���`�їD}6{w��D�&���;�>)5v�c��ݓ��,bwvf�Wog�S�n�/&u�wg�"�T��C�B�ʾr��#�\�
g�c)�	�:yd��Q�nK�s��D�bV8lg*���}+Tf�b8��{\��1]���w{� ܾ5�	���1M�e�����a� !���+࡮���ʰU�&�'R���K;j��\|v���'q7a<�]���3c�¾h�W�4���Y������
�ٜ���`���7��C�&��cĭ��)Ł��](�b�����������+(@�g/�U�	�h��t(�w�=����m��謕��fJ[�c�԰�]:���{��x�5��I)��ì���p�֯�Mb��vK�}t�WP!%�:�K��d_[��j�Z{���W	l9�Hn�XP�b�<�\e)�}�b�F��by�����=�w�d������!��_N��ݾV��ĕD��U�h�*�H��#�_f�,�R��t���_ 7E�hk��4¹����Q�K��7ŷ]C������7����={��S����}���fj���#y`�LA��܇{0�����f��.qH��NJ�ڀ��$õ��²(���zV"�A�CWL���|i��y�z� �W�]��e��S𕼎n%�V��,e>}������w-Lv)�X��.���f'id*%6�2#u���iv��/�3�[\[��:m�����T�"H��E��Q�k�8wu#�����Gv���y�yܹvo�:���.o<�������Q����D��Np�b�wW-�-x�RJb�'�<��d̛d���Aå�1N��u<b��<�A�����H�;��q�ݺ��@ɮ\�r�W
'�睉�1�sy�&)1@�ι��R�o;���LE��8&�5#s�w�1Iuvfa� ��H��	�L���xs�ɼ�N�.8󮉼��J��B#x�5�.]0��]Qwv�p���%��GQ!s�n�G�ux�P&RA).�H� ��#�\�݁�+����t�d]ԙ�t��w;�w]'3�B���tܺ
,c+��Gq���K�(�מw����Ɍa�]����̷w&	΂��(|(
 TA�AE�t2>j=�:��Kc��M���p]Y����#�:[��냢og}WE�^I4_�_'v��{nTT������a�m榬�]�A�)�S�3m;�b��:~b;�� �C>��"��TGb�>�����K����HZa;�
����L�u��3�*eJ7��4|��\���).9�ۨ_.12pBj�؅�5�ѐ�L1�h������J���Q�G�)�0J����U� ������Te���˸�lR��.��RY��{D=3٭�ޓ�fЀk��F��w<22i�H���<�0�BG��ʰ��B�����}T'��Q�oI�5�]σ�˦��{�k~��Ă*�h�:���������B�-�̡�����\�pL.y<ա��G������j
�{ΖJ�S2%U$B�$Ϧ��[�,.��v�f좚ŋy�y�$}-r�e�,���z}���\��u�r9U��m�I��ц�ƽ}��7��ּWZ�fQ�k�p�Y1�~�IS%��̰9�sGNo��ZT��NJ����.oۈA]��G{)��bx/�̹������X���`iy��/�1d��ԓ 1ruL�����v�.,�] el	ݚ�ZM���W�i��9�tާڸ�l�٧8 ���y:���~}��>v��U嵸�v3H{qI'�<�լ|b�X�������SOzu����{���}K�e�y���pQ��,
JNu�M�ۋ	�cd�0MާR�}U_W����^^*�����h,7�lr��v9Lh�����I�����&��ǅ`\�An'�(_.��g%�Ǽs�^�(��g����Q�\��I�f��ƹ|��Y�͂�Ա��Wx�<�����ΥU��f�"����a/��)�g�Ai�77 ��ooo�.����)�uݢv�C�z�����m���yƺ�[Xeq�.�\>���ٵ|�8{�����֋W�un�`p80'��q<�φD�L��u�io'�on��<q���8;���n�B�����n �,�;�(��p�䊌S��k�b:�]pcs�[.����C��^D܊N�;#��k��'��5����G~Z��gÝ=9��<��	���g)��Y�����T��ݞK/�>��iW�N4�
�����\k�lTx�����\���C/Mmln����g��9M&�s��vㅗ8��pj!A����<ҟ���3���ҕx��c��}6�/��#=v�֤�Vq����U\+��#���5�@y|v;�V쐲���cS7�fUiw�c;�q�ܢ��(�j�͔�E��u(_4�X5k�T�2 ��L�lAg�M� d�h�!�����vWN�&��ʬ	�}�W>=�o@�}�9 i͵F�8ï�\����JӃ�\#�������'��  �ɻ��ɪfg���;�1��U�g4���q/]D��,�(��]_v����67E�c�!��H�������7/�CW���V�C�H�b���$[�\�b��:ͣa}A[}7��֭@}�B$��/�/����1_.B�yL2zu��%�4r1�_"+�z;+>Ŏc�����:�U|�f����=�ÕE���en��>��O��9���t&�NZӤ�Ufwr��I���2`z��2UyU�V������N��� ���b����a|�,vD׵�"z^q園�Z�|��M��ߛ��|}�Y�i�5��PUc��k�l=���}P���9}M�����I��)[p�:��?�w�«�����pg�V���/�ǉ��.�3��ڜ=@K`���lW���
\�7�T��ds�� ���V��:���)᫫W'=��&���û�b��d_!�]�	`� �Ĭ���P�8X�}7�6��s���164uorɜ�K��p��1#	B��aF�ar\l;�'i��ǌ�%}�N�n�ag����|\��va�y�Q�D]X�l��/k,�0�h����:��D�x�=j��stYM��m]�:�بk7�j�m6�>'z"��	�錦]	(v�<����k3 6��|��m�0�Rt�����
#9)^�᫂6�{6�����_i���������Z8'�&�:<�X:SR�b�P���_(�,h�C�s�3��5��_L���#�R0>������8�#�
3����4!zxf�ӥ;T�XE<�3N�o�w:ܹ�B[N���Hf|�;_6�dZ���O��'��w�$��J<��KL�G�Sr���H�őN����)���Vo�7q�#Q��$G׮��o"eUwk%[��=>+���H_>+��;c��D�V(�싼ɱ6����z��6G�n�fuK�bԝ���$h���A�ix@�ǡwWԓ��9���;X��V��i��K�U]�O�*;@yN3d�:I�& 0<"��83#L�loIu� :.�����]�i�޴t��g-���HJ���3��X
0ą��0�v�v��e�^�)�^�ݧ�ٲϲ�U�t�G�#P��ژ}���']_c�}5��×f�%˰:ח�E�;���{*[ބ��j�x܋��f��`���5�H:Y=�&WI�}��s����[�`fp��;��&��A��T���G��'��r5���n�M�jL�M�����'eP��I*��mH�K��Y�`=�\j�J�9�����]'�h�W�6�RmZ�.��_y(������	��ԯ�Zo����W�_W�s����D�5��V{�{ѽlh��VXJe����36X��fĔ�*�BK���|��K'�M��r}`��4ژ��%h�t�c��?&a���^�M�)�8��Z��AxnW1��*���/��h�z�����(�dx�[���*��x�;@<��u'$t�y
�&�+p}'��('�ZD`��3(���s�%�T	P��(��5�����$I�ɵ�ߐz�}>��خy�3�l�
y���㼨�8Nv�pL���eު�Wo
������B��[i����g.���	��T1Rskl=��v�q9<�ʕ�
�+�[��[���Ol�8՛��y�Ͱ۞�(�����>���\v�ܻi��,N���My����漬yo9
��5�����PB_wnF�]j�M9}֎>���Ɏ�� ڻz��W^��w�!�J\}�>k�!����ބ��k��V��+���Kyk�v6�b��f-�� ���Ş���i��%OG6��m��%@���;G��j��9Pf�]92h����wW�-��n��,��Venm?�<6oa<ʵz�=�ܭO3CgK�mT���o�{^:����f|�ԭ�}_W�}��r[V��t��B9������D)�	W�A�Ϧ���6��.�V�If5��*�8c��|gL\)G�8��'���ꉌ�J֑��y)���K���"ǵ`7�Gދ�G���C�ょK��61��P1+2E���l�Ƹu�ݞ�_���b�c7�s%��o�����x�I�@��~秜��~�+��_�r��Do-��I9��'����w�o\���a�7R����:�ЫK��_M�l�}�/g��v�0�B���ι�����ݛ��&j�f��x]�ޫ��Q[�-�񫵽��"�ĝ��n�}�?�Z���YV��*ͽ[��+8��f z��G��x��T̓m弞���b1�hy�����*t��nMkJy��Y�>�/r�X��yOʝj�u�jp�<�s�r_Fc��c���Z:�rp�KZC9&P5z�w2ޥ¦d=�
�V��`�&p����5�q��zz�FȾ�����ؽ�<� 4�:��8謏[q5�ˍ
}n�Kn�e}��6+�9���^"�ٚ�֋��:L7�.�mF\��>�&@�Y��n^t�;]C���������(#��tw��rR����PV�T�[��z�z�|�sY�+�ŧ���j�nӃ���,5�nA_>WR��=��9�٥5��nm���܍�g��I�ُ��2K�a/����CK��866r��Y�[rw(�1d�ˣ�zZ�^�w�پﷲ8KF��V���[�뵻hJ���z���-+��׭����C�f
{�&6����oy�g���y,���ڇtӄ9<��B\+V"y�j�(œ;-�)�v(�8�᠕�j�r�닟{P|�RG�=Mz��������(�ɩ͕��Q��&u}�9;�۔���W�o�s�/�#���->�Ib�=���h��]�9���C� {���DW�y��]7�=��g��[�ug. �-�2A
��I��ml��=).%���YPZ%��.��6�r��}<,�ք|����rw��Ң�Ձ��\�/ V �u/g���q�%�v�;���i.BA��woZ91^�|
7v�R��]��X��c�x���sL�tL~܆L�;=q��g-�/{���b� �XZ��}�U}]	݆��k��y.u{V����<df��٤R���N�wʲ���0�.Iy-鞗�T	�qڢk;�
��'�����򒖐}}|����_.>�k�u�g.`v���!��Lv$+�ϛ�����MU	���xfJ�H��*u���O��C�Z)�\'�����s�{��b)-jiN^ܕ�c�윙�>�{Z��|'����~��Oz�o<���s��.�K�S�u~/��חӣ�S����k�xy-����}!E���"�VWVM�;�w���s����������y�6��X݋
V��TY�V���걊��۹�	v���U
��)޵�vC��-8�	P�B�&��cw��n��m�y��o���J���s��d9f���u��v��N����Dd����	-k��o��&���	�"�5Ѐ�h�ڞ�j�i�ob��V|V��o�1�/�K�m?p*�d3Ē9Kؑ����-X�yF���t�Z	�K��ls�U��Z��\&�:'�s����I�|�����5*�`��ȯ :�K�L��ؙ7r��2��d��-;ѓ�U�����#�;m�w�stl{�ױQ�f!��%P4)�ԭ̽)�-ὣ�%�������f&�͙�����0и�T��R;P:��%kͣ��=�4
4N�F�\>1osn��p��}F�I0i7���]�1�l����7C�����Yig3��vV�5�f���_X}B�W�A�@9T6Y�A�n��2;�)k\:�7�㨕�_u=�>�z�_uM��(\P�5�����n-Uҫ��we,��[U��Q6��V���g�}K�q	=k.+2�(M��,cs��2��fs�k;�2�x��ʰ�?\v���<�v���`�LKUү{�iZNn�}]��N�nkC�u�c��s_���]^ޥ�rI�0�T���ƕ�~�՝��g:t9�3�}�(��c��*��u7�l����sY�{o7ų蘜4�1�ݾ�ؓ��Q�g���%���}����ע#%!�xh��b�M�c�S�ٸ�7�7���U{Iz�&��ng���Ma%��wK����\��̪�G}sjPY��q�������z)}���:s_��b���ҕI�v�X���8q������ �Y�����|�b^���͜����S���n�T�]W�UW�q+�����s���{�JR�*1�X���������z��F:���O{А,�z���U�ۃ�\u�u�l�)O/�[=k$rX��[��1.�҄�V}���XR�ޘ*\+�7�b�`r��ңf���5~��/A���mݵ�gF]���u|�uJi�����	�o�WwR4@���Kz��7�����p���礇4J���}��О�D��~kw���wT�Z�
q�ǒ��sW����f8���<ʼ7]J��Q�����xvY/�O��7"��:::;�zX��8���s�¶�O+E���u��<�)��m_�nfT�O7�}�d�������l�[l{ʓؖ����U��Z�L���t�뚇��
��b�>�U�N�Ɇ�E(�/Vs����ؒ�t�Oj�9�c�[ꁘ�鷕�Rѷ���
��'����Y۷��NY�r�v��7���=`j��PD�('���6�˔]��I����a�=��"*�,�i����'I&l�����>�}��������0t�,k��+����o6�m]*�B��l�Km�کظF��7R���SekX&r�����7e*�\����Z˂���{<FnHՑ
�h�,�}3����O{E�����6�V;ϝ>pO)�b ��]2��P"}�V�Cj�ը��m�r�����V��������>-��q�u�����e����so��xn�+�IB��P��ᜬü��R�b��'r;]QL�{Y@��&�U�Mft+�W
{�ÀcT�������ۨA�i����X�p��{�V�Y��e�������5��'}�\ň�ϑs�_u�E�m
z�kV.��Y���b�L������&�$������X�p-�W/m]�+��75�?��,��(�7&4i}�q�^&/A��շ(����▱�g ߔY+�QR=���|p U���Һ����QJ��1]�y�9NnM����d�i�'�I�z�J���a� ��3a�A����-�[,�[j`�節��.�����e��'Vd9lr#�L�Ǽ5ہȯhV����t��f�G�PO3��֜�SB�e�\S�s.���A5��l��.<��R�z�t���M�ʨ�VN�%�Or�����oH!">�k�%J�\����S�s\�K���_ǁ3��vj��;z�(U��ܩ�ɼ����Zg@M�+9c(�Oew�3��
�r�EҌc�Cq�19ax�wl�:֖��@�_b3"�E��l7
`V}Ϭ��#z�r�JE�z]���Y�7NT}a7��C@�'T*l�Փz�)�`]��d�C��|J����u;Fw"4����˄��ղ���;�qrӥ�����U�J���J���T/�6��{Zao��R�C+X��]ȯqC�P�yЙ��~2%]�Y��+��JH�j�Bt��#��v���ۡƸ����~/o4�
��a��m�Q�}
���.�`�$n�P�q���9��_Iµ 1Q�B�m��
�l8\ʱt�qT�)��m���[��R�fBzoU�C3/V1��F݄��}(�����F�{[�$��ҰF�X/�'��oO�JL���0�>�,�[��qA|��G�:f�83'+[ff�(��Lh�����vR�",��Y,����-*�]o
=��q�No	S�^�1O)x��6!����ov����������r��3w���*C)����]�����ǂI;���7�7����[YA.�:���'���u!N�8��yb����ӽ��O
��ss�y���Y��Z�d��g��F���x.XR��meX��z���N�V���Q��Z���g)��.��kƩX[�t�N۽j���9zDMr��4+z�X�䒀�  >� DB3\����]�$��ݻ.p�J9p�4�wW0єRD��$�i��˴2"�$��L&bI��Q2�2Le!�����������B�ᐅ2w]ʹ�d���Rf	�Iws���q*�Buܠ�Zc+���ˡ�ě��0�+��ɤfa(��ۺ�E&1�I��F4s���s���H.��I�ҙ)λ�$RX�u��H�w8lc��5%.�u�� "�\�@�e��)`.cr�1���#(	7v3��d�J���0N��7;�G.�$)Nr"d1CH�% 2!K$�R��%��a(
�}@V���<�u&6��Y��,b�{@SZ��w[i���wvt�%����z�`� z��[�FY��B���P����G�E�^p��[�9�gu>���sW��� �>���{*��˜�ej�ɼB57���n���8I�.��;'��8�=ڙ��j�δ��q�T��wqa�{QJs8ϳ����)pw��.9<gFf�A&�vvǫ���]�@�		��ժs��gn~G��	F��cb�7�����X�6��o��gbRsP�����45p*�/�T�U+����> �[\0�emiLn�s������6J��ʢ�cG_������[8{�>��{�L����5�C��rۂ��XR��
�伫�t��;���;�"fN�*<���s��̆�%���]�8���\P�\�Wo��P��-�t-}����k�o�TC�v��,�!���;,T����i�w8�n%����Uxm$ҿ�|��1M�����}�4GM8-Δh;=aLÂ���{;���gI�Jt������˾۰���*��X��^��Qo7bw
�.��|r���&Խ�������%�`}nor3+����Ҏ�t�6��˕sAR�,Rw:7���r��s����n^˒�l*?�<hC9��3e!]�Ku�Ͻ��	#���ʲ�g}uǢ�O����+q��|�@x�Y�ʺ镭������J�{lv �u[������r��q��ʍxG!� �߯��Yڥ����Y�;.��p�ǳf��o)d��t�rjb_l�u�E����(���j�y�O1n��ַ-W��pی�w�O~�/o�w�F�ֳviiKJQ�or�i����������_U���O=���#��3��#�[ׯy���*�<Ea��
]�Q]��r*��������!��6���gL�y�)�TN��u�);��hga����*���g�J��lB�P;)E]�u2��y��:7r�$���۝������_+�y
1�\Ay.�q� �V޾�������%���'��G)Ўz��P�_�*�&����j���l�oV����8j+vJc1h����Wl$�1v�����CM�T:�{��(�J�.2p�~_�`ݵ�C#���}�H[Li�o��$�b�k��.���s�%"楻)��Sn�ױl��i�v��t��l�����}�n�m��1kT�J�C�R������{P�{pV7bZk�;RUjC�τ�$���xexv�7�����:T�QN�!�k�!�ί�q�崚kEi�-��3+��ۑ�3�|ލ��.X����z��${��e��R�.��וQӆQ
c�JD��Z�x����ڏ�i\�������,�U��Ό�����ær!��%_
}5+s.4�fyY�\��ʺ��$�6d�oW���a���L*C���@뒵̾��5����ykε����	�W��DF���
n1�9��6-m�`YK^{�ݭ4�I%�s�8��R|��i�;�7�3Pہ��k�.�T�NF�z��_�l����ZSr%3���s̼�?������B�(u�p�Y����i͕V����ͦ.).���}P%`��N���g���w|�F��Ҟ�ǜN��Tmsӷʱ���Ǘj�riyc�Br0�7���ǻ'e�g�(����[IT����jru;m�W��\S'0a����
�v��Vo��{�5����w�y��ì��'���:�5��X�����綥��^�u��7��ٵ���������TM�P��끊�8�\$�7]�^IOS����=) ]������ה�`sٞ�=�EJǋ�P.�kesg��3�U�W��uH��}�:隞.��;T�u���a�Y�X{W����#UЕ��j�cb����O�g����D8 ��s}�Ν= N[��i��DI}Q�ʥ�������o.�BN�*������Y;'#��%�{d�x����t[��b����,	ޝ���X�h�v{���1,��m����Uf�;�(�?y�=��dNuGVl�N��t����Ok��q��jb��3��R���xD���ձ'��ܝ�3��>[=���e���������X���Y�D.��;��V�^=1���hM��s��_`�����o���.�BL\l3�s��G����������k)��ݰ�׻� �u²��;b��9c���yt��곕�~^p��J��Va��	���<�����o�:k�l��r;
�6Σ���<�4��f�;ָNj2�	n?g)�^v#/���%v��V�)�_�}_U�Mk�4Gw�3��騕�5�ξ\���RL6b#���oE�ُ����q��t{r˗[���9̗�NE}}!^��/ǁult�e>���l�{��Tu���۞KV��O�����L�g|_g#k9�����B5m�����vk5���7����v��ky��{s\�D�Q;Z�/Wv����T�no˖Wf�ߗ^g����#ʎ���qŝ����G��垨u��rͽ�yH��O�|��ǝ�.���k�U�!���<��\r{H�w�&�'��֔�چ̺d����!�#6��j���X��yX֨cb�9s{����K��˅�;y)d��<��ߖ��E���zm�L��*1�ݨj��-��Ǭ��K����C�߸�g���P���ᥘP�,��7���P&7U:@�0an2���h�\7Ϥ������9��1r�:5�^�x���Z�]gT��J�n�4�ꙺ��̅���;�����Ж��-���B��t�]Ŵ��aF�_S\�4�c]�'�}�"�{��닮	2 �}Y}�-{�;jeO�km�i�v��i1aJ�邠��C�S���C��oe��t�úT�lҔ��ֻ!�����軂�`kAތ�u$�l��\�OG*��J�_��q]K_0������)�;ND;����+�.���r��dcϵ��~����k�⺖�ԚK�u�g�Hn�[����ˏ*3v��#G��Ǘ��V�F�:��5.e�כօZ�F��V[֎�B�C+]��*���G>T1����>�)��`ӣ�ݛ���fv-�Ϻl���Q���е�ȞCg�kh;���ܢ�lJ��-�e���{��PH�F����$�� ��&-�S�̽�"��YW�}]��=�g���&�l�^�����΂\>���|՛�QQ̭x���j{����%>�)�t�����|�x.z�9�Y���[sܭ�[(^�I�cWbu���M[ywd��mJh;ھ�ԶL�}���^�%;�>�.��M]�/4�M��
U�����N�9�+J���^�/}�44��]h���\V�Bx�y�iVCB =���:�ݲc�y�ճ�v,-]o5ٝWҠ�hi�mr���_��UR��I���59�Vn�h�W�57Ry�����h�͇�C�]))ɲ�nq��K7q?O9����5n�g�:�Z������N�zk~�zK�~��N�S����6�o/���ݠ\�<w��eCm�`�f�����*�XT[]*��E}��{�{�済��ݻ���#Y^�d��(�yb�}�v�۽�x�TB��ކ��x�,AX��C��n���76L�~�z���_�v�b�Kf�Jy4ֽy�̊�R��w�'��)k���u��!�9��O�g�?W���W�r��b�\���z�a�:����O�|<#y�<��]�C��O/�q��\W�v��8�s;���٘D)�	T�=��(f��!|�����wy�%��*�8c���o�b�L\t�v��_@�/fw�c!@���֞ө�(`�%T��zL�?/n7#�V=IL�T�'Mg}zN6�dg�F�҇ �
u�Rی��O:c1��5L��ޝT[�	:�)��$�R�0�j3E�	X�8�S����V������= �Pb�'%8�C���J�? >��:�fs�ί�</z09�EϨ��MF.�9�h���!��`y[�� ss,bsk6���_>�X�� ���y��OR>�Q�ڮk�D8X����gLw���j�ɥ���p����i[J����r�;�	]�f�1�@�����B_j�7;Φ=�vJe�Y����r�kA�|�����W�f�:F��`�L@�#g0Oxnge:��k�Z��;weG��<o`2��2�3wŜ�WY0h��d��zo���=��Cg��Pu��jVE՟H���t�s�g����c3`YZP#�xu�;�kSl�p�:���p���j�cb��������ܺ��+.�"�ʴs��1hʞ`��:�$��ej�J�����ݧ�R�'����R�xoZz�[���'~Z(�z�Os��.�R2�<�
�2���ͫ�-�{a�*t)y��}�)�J�j��0��j�ě��uڮelW\�*�UaY���?��T�;��s���CuÓ��`�V���"�c;VT�����lWF�������"g7x���"�I��@�k���5ڎJ1��>ŗɽǼ簊��l-��vW��w�_o��ܬuϨp��&mK��i,활�
R����c:��9_:��,��ޓ�KE��M�bLV.�����$��_�ZW�opSl�C�P
�����[�r�U��%u�082�ju,����3���|��1M�J�g��z忧Ve��h݊4��c��Jܝ�|�	���&��ZU� p�s'U,]#0�u��u|��G���Ĺ㿓T^GJzg{5,k��:�a�Tdll�b0���<��Lŋ�_ٽ����ƨ����Ue���-��H!W'�I�l�kg�z�]�%�bJ��3�ڮ�c{���w��ת'�3���/<�ƍh��b�	>ڈA%[��33��.3���e��K#��ry�ڛ�%-#o;��8iS�R�=����:,���~��i^���/�G�	C�F3b�Ӄi�����K���r��j~��UɾV�Ĥ�Oy�����o��:�{����SV}(X�G���J�2�Y�K��q5�7D{ﯲ�U�/_3�.Gk�WXF/��? \r{*F��7-��Y�촲[�R�69<�'Ӱ�p���:���}��Սj1��G.oA�BÇlf$u[�t�Ӛ�V�/�c_séo��r��Q3r�/Cػ��B{BX9+ک[�k�s@��7��O�"Z|�°�h?>U���㚡1n�h�;V������k0a��T�i��҇��|�;i���og�Tp�+pз�)��/+����t�Jٯ���cZ�|3��N��������e�cX��v�N��,'���C�]��_0�xZX��o��YR{*�f� �YK�:�(?��]��.j�]��>�����;#�F�bNP��s�LD���à�\����+����j���mg5����9mT��L9h���\������v��q�)C�����s�t���Z���jqjg4Ҋ^��նX;��b)�w�	]��U��q�a#k�˗}��2f\,�����ޠ��kNPp�'w5'��5�||�L7�ב�t1�r��;�v��pV�@C^3��Y\��;�i,
y�p\t�5v�>�X�M���0o\�����9E�Ւ��.�1;wkr�.�p�.�!f�*ug
�������l�n���;}����Y��k+�"���w�W�[����q��X���	���8������'l:���cj;{Y�ܨu��k<����K}��jt[�����:^�Js��h����]B�kZ�8bi�sb�է�M�d�+ՍV#a���C�����J��i�҈�,<�+r�΢�.���w��|w�*Y�;�MMI�f����]<{c.V���ī��a�׼kfQE���e�L��7��c�}�r���âGueK_[V�
�$]Er����g��*�Bՙ��=��>�H��u�+�;��75V����9`�a�J��)�J�1��M��D�!�d�8�*��z�h�v���w^��-��`��J|ګG-:]���89���Y�G�I4����V����c�WfRj*�o���5���Q��";�퟇��VA �n����\�Q�P�֞XH���\Xw[%��R���S>�wə��e�v�*͢�l+Rd�b	�Y���Gs$�X��!/z d�ꓶ_pw,��6��"�����dr4�y�v�D�t����ŝ�o�v^��iۋg�Na�h�)L5�vT�[H�quqj�wTo���Ϛ�ω�a����(ذl뱉m�Z�g��.D��B2�#�{�Tu��a7l"t��kg+��)l�W�J*ѻ~BC�Ί�=�Z�� �S��u�%�}�Le8�u\6nR�7:M��fptm}����V��i��0eϐ�)u�r�:!o9-'���a'6ٴ 묳��Z�;���8��k+CǕ-��cs���j-а��S�b$-J ��i��jop<̛Ȧo�Ϭb�Y����w�5'ٕ�sshhU��A+�v`�61U�D��͈u��� "W��Cg�zLB�swj˩���5o���"$:�K6���ܥJ��F��p����]wk��&��*-��c2m��ڙ�"V[Ut!�q	8���@G-se�r��Ѵ{5�	�
u��N��t1>fF�9�n��,�T�N��pQ:�cQf��4*-�$x�/�FP����Ҵ��>�`��q��7U\��`�olA�4���\�n��0]���a�Z��z;A3&*^g����ۖG1�dpfi�<�r�`�yKr��AV�r���V����ַ���*�:F�v�[1���r{œ�]���\Pn)M����9A�D�q�C����뱻�p��5Z5a��[1�r��}.���y�c0����������A���e4zp��A�\He� JI$�$�0�R&E�LQ&�l2�\�s�4�BIb"h��K���&D�P��$Q19�2��d(i������$P�MݮD)�w#2�E#��)�i&K��b�J�1Fh4̆C�D;��]�(�]�ā���%��2H)� #I(�41�wt6)�!��Д�b�a�;��H�1
C�w]@Rcw\E6JBE(�@�H�)�&�b��$��솂F6)1E��&3$�  ���$m�BF�F��&�ɉi�����	�1�d��3l�5����%���~_��������t��%cym6�w���y%`�t��;�{�y��qB��'��a��73���s0��7N�mՋ��_3
�2b������4F����A��㕮ȞCdZ��=���)Q�W˒8�v��ȧuX��@sW�E}.H=�	2�^�X�-^M�����jY�����Y�c7��(�̷à�^��H1�
����tgzK�;���[�7��"�jk���ʗ��z�WF�D	�U�N��_���}�{ɗ+|.���Z����ؠ�r��
N;�b��;J�ww�
�!��8g��F�}=qh���bίGs5I��5N�bĦ�	������i��nm���cé��;ӏ���B���~�����&��^�W܏ɧ������=U�l�\U���k*��nm�mI[Q�JU���R���n��r���+tt�q��jO'����W S�`!�Q�`��㮋�Kf�Jx��龏�#وUfqJ�t���u�cK=h�K�o'o��u��� Sө<�W;�J/3k{�@�?_�����%��ui��R��+{{Ou�n6�����l�i�p�r��C�-�y�rf�Oo7�u��V�Fಧq8�f�'V��DT�����p�UT�ox�j�i�vV��X=�l�����s���ˇ/�8��U���O.��Z2�^��3����]�\C��C�����8r�#�j������ٍQ�9�Kֲ!��_6��9�!O�!*	zrfP��p���ǋa�Uϙq��]�!$~�OuÂ�u|�@x�}����{��ҽ���=��XwZ��:O��BI��/u���|�LF����f�$/=}쪷�f�X�ڱ�����(_A
��֞�a�`<���J5j��C�-�Z���;Oy�*�9�zv�Oy��$�V����Vg_Xz�<;\>�u<��1�<�=�.ʦr�c�s}+5e�3Ӓb�m��vsY��޵�F�~�k�k#�̢�#1TM�d�F�����>ǻ�p.�N�s��9=�2;�f��f��� �]�=0$Q�ob�Q����Ie#�PR��\x9�/q��6_�#%�ܱSU�"�^
˞�g=�\�m 8��s#|��-5�*
4����xM#� ��;B�}��N[ݽ��
�Wcq���-�v��9T�T"āQI�ս��*�Yg�]f����?-�ԇ*;j�������R^�X���v�:���ʋ��P���Ns���9� �CG��S���GљӜ�%u�kj�z��o�z���{-X��-��)��%���S$Y�w�lն�J;�������3���Q�_m()j��5�����]�f�z�z���j�N�u�y�ń� �*���lg�>iy�O��ݙ�l�7õ�0���Cڈy�l�n��a/�����$wm���1Cgi'�i^a˦�9����ݳ���}2_D���`k�"�WA�.�vNrz��]ݎ���%�h����ʝ�l�=�!��h>��ﵱ�G�^�CI���ϰy��;����4�|��TCocK�̇�,�]�m�/�*K⋨��7+rkw�|�A�I�Y^þ���	k����䜤���-���:��Q���}'=��^�
���sp7�V�JP<���v�>#� �_E������D�l]�=��pM�j��cx1eR<�W��n�
ȵӈ{����ﮁճKx ��3f)\�����P���)^>�*����t�ou/q��
�ۛ5ZQ�+;"��8at��ꪪ���x�GkD��-@�n5�3����:`Z��;u=�YK\�Z���ݳ״��oc~v�oud΂rj�fCg��]C1hl�����8ޤ1,[���߶��q}z�>3΁�͋�dĹY��w�+�����eY�!��U�\�N�R�X��[P'�e����;��റu�j��Ϝ>WR�Gk��!\ϫ:K���iTAw?ʾ���)���{
<���񼌻��y�"��7��p���ۯ�ߔ��z��Z)����s�I��:P`F��o��Sm�?}����B������;�Q�j�y���_n��/#n�r�R�\������z�aUZ�PC�Qj��׭��&����=��Ů:�5H>�l�;.o����d�{�hJ��o�-|��B[Zk���sr�v� 9v�]2vNޏ���qtRg�z�S�QBw�Xx�yJ�Y�kzo��I�3vHm�S,��J�CgmAӠL�"�W�$�L�d�Υ��\aUɇ��X��~�/5������keZ��hk@��M�љ;]Ǧ��oS�Ҧ�pͮ��l�R�"Lރ��_��Sר��v@]|w�\��g���7����.寥�������GZ��GL����ZeCT*L��p�|�Z/����xjM&�Wvj��|�-]���e���y�hR�8����0���v]��pd���-��7s��ْ%��q�M�l[�ȘT��ԃګ�p�?d\W ��6e��akx�mi�r�{_>a�'�i$�M�>G"c]�1�l�Z�=7fA
�������]�[�V3{P毬>��}(	 ���Ųϰns�	��U��t�W7�%���E������5ͽ�;���t���L~!����.,|�qUpEf�Od�J�����e�ڝ����
�ޖ<�r1�ë�ݷ6���ѥ��W�\�x��ʉ<�_�¶��H�{�6��au��ʙ���9�)�=����x�������ú�����P�[:�9Ԙ ���n5�W8^�ს�j�GwNτE��N��zǡ���c7X#f��C�^�D-Z��ɲ�89�C�T�5�i�������c;��;3ue���P�q2�������>Fva	�ݴc4��~�:o^+�XT_1�@��\�/��]��.��;QLwC�R�rT�c�c^���ܞNN��]	X�����	e��\K��VuB�*U�d�'kV���� ���=������9J���kx�7o��{Q1=<��n�)�Ǹ��[�1c���⠇ʤ���]P�lҔ��h5��&�c{D��[���ˑu����'�
W��E��	wd��O��=:�;����l1w���l���)�\F��ϸ�[�\?�υ_�#��5����DLuY��U�`3��_�ZL^��XIqY��
zBU4U�$�F����o�_%}�z���e��o�������d���AV�Rt�kŶ�p���;��oM].��M��O��I�pˍw�9U`0^�M,�WOxM�0��+s.#+���jڈ\��j���u<'3#�7����]�ux$1=�,nV͟[άqu�����9�R�if'��+5�s�O?:S�����?k��� ��qܕ���֤�H3@��w��Z�g��X��5(Jp{Y��Y�2R�+`�J�+Uꅢcoc�o+�s�b*��j�7/UrB%�����yO�ю�ǞKio?D�=��='���'���'�-��7*�+�s��·�1��Kmv�Z�� 4Ef�����ۼ6�B�J�.^\BN5��]��w�H�s��b�4l֊����=�smmZN KC.;TLV.al)x���ǛsF��̛ ��|�ѩ�d������U�=�(<��B>�9ϳ�f��u]�N�ݘqFO�����7_s��\�m(J�l�c$��M��N[�����%����ڮ'&�u�-Pƣéo��r��|���J
���������ꪙ�/0�|�w�-�T�I.�i��g(����PC�Q%'�%2m˨&�p�m]��o,�/�ۇ������9m��ذ�}��<߹�e�a�R�;%تj�X�nz�N�%�)Q�vN���(�um��J�T�@���s��G�~C��/;��Z��9b�i��[ٕ.V�k�ϭ��v�g��1QU存��/ŵ�_W�����*����Y!�GbT��!��_)�c����	���R >�r�5�8N&�N;���մ�]�m��vgB3d+�Gn�/�	X(6��⺾Z���J��z���xβ��,��U0X:t̉�z�W;F?��r4�[5��y|R�[�Ri/����8���"T0�n]f7#����g�P)T�rV��s_.Ck�\�(�f��֪�7������h[��Q���r�|���@ے�&�N�ܴs�ڢ*f��d�����^�Ξ2A���ddr"�ç�يUJ�;��`}�ߵ��f���Ͼ��jU������ᚋn��Ć�6��:��>���X��d�̛�kT��c���͒������tvl^z���F�}M遯�n�\�Ѳ���)�|���+F>�^������5�WDt��!�i9�pS��n��BљG�,��ʁ)���;�ϛ̵��F&2R囇�s�y��D�����*ÈT����u�lʭ����H�NO7���#l�"�Mh���9��V��b`�SK��.=u6��Gƃ���B`G�����5u�j[�.s�=U���<qs=|�Y��Rb�h>�3��o3X)YqݾLt�.�����q|(f9͈���rx���W:�&�X�ws^#;'���a�\��z^�6�Vv��d�|/�u�U�/C��c[+0�1By+�6���灼��O�OB�_.ª"���þ�z��]3#c�ނ2���.�;��.97��5��=k��Э��aQ18{�[�k����@�_������.�_ut˝����Lg"��&.���(fkY�N����,l��L�Z#�L3�v�K�Q��︾7�w�11����ɹ6�;_9fa��JC
Z(-wq\��uc�yG��ö�[�i�ݙ�h�sȆw6�*�(�=)T@��j��Wb����M7����/o�W��Ci>f����3�4.3�HLu#��<�uՌ��4����ęk�R��[7��.a�}E$��Mƴ.3]�<��F�	���w��{0Λ��n�S�2�.�V3{y���7�B�ھs�=�{��D�Uyӓv8v����p�iQ�;PY>&�2�8(����y{}�TS_I)� "uq������)�2Ө��w�
���N���s��^uv������+��@��V�˙E���wj�e"<�tFF��v��{��>�Μ��/4_�_����ZSk<���~��5z�_uM΂Y"e^}]���8J�����~p�W��	�t.�����]b�n�W��j����_F�㽚��[��>�����&j���@l�b�����U�/�<��ur�d���������s�'���k7^jʳ���s�t� �=���$J#={���^��R��i1Isb����͸��gY݊c�ȸ2��N���I�Wc���e�]6z�ZC�%i�ҵk�
�C/���"���7S����^�TOzP-�/����p�R������\C����Zz��y���oV+v��1;�a��:`�?ʢJ]}t]*[4�<'vVAWqp�ժ�51�ERp�[Q8�}	�v,)_oLAP`$�%��K�	�&
�0kr�Ift��p�'p�>�lg<f��2�]�p����>�$���@oFl:ԙ�Ӵ��y�Vu\+��PΨp5����� �ge�p�Ďg�R���cye�_V7��\ձ�����d��o�q�+p�Mx�w�:
���W._���&)o�邸I�t��JtҲ�����1b�X�9on��:jdi���x��r�_:��A�2����@ւ�|#�@��K��n+{E�V$�qR\�D}��sXH| vz�W�eڴ����9�2���Dݭ]W�ݶ�V[Gc3�ex��PNƗw�]���
f����-���)_<��a�e���m^�)Bַ��W&�P������*=r���'�Ol��KVr�èՉz-�+o��C�j�����GFWmv���Jn|e���%��Jm�S�T����o��/��� {��&v[G�W�~(w�H2��*�5�����s�I^c5L�%t�b�
]@��nSu���Z>�	64X����CV�C��q���`H\��h��H��1��ڼ���.�ѻ�Lc\U���iqXC�l+K���Gan�V_-�Cs�[x�mi9W��a��J펦�}?wk����\�O�Ps4)��w�*%��cd��fwF�%sin6{2��ꡛ�^�JA��̗L�� :�Ǆg���(C g'�����+��VdvaqBؕ����|����̲%^T��noE�YQ%QS������ͩY(�]0P�}���>c*�0ż����&�`�c��me�z�����|�WZ��ȇvX:>R�@�K�(*�_Pp!(9/�3�Z�Z;W�v�UGf��|�ITw���q]4x	J�;���d���3S�J��v�`��4A)f�أ�9�O��nحGQ��8L�C��!�)&�<K�w���r�h��|6��$PM�B��=�ۭ�l;ѥK:T[�]��;��|Gma�epvrG6<(�v�,�[��嫱z�t�ή�sM5T�3�I,�9�E�:Z&�wZ����B�i_pt�yj�؛�2�ԊV�8��9g��!�`����v�٨7'^Y�}1�F���(E3"�d���,�n�ĳ�+�]ڳ����D�R�8G"w��:u��C�Ŝ���8�{w��P�����+	,Y+�gt��������	�Q �L ��n֓�cE,�8�#v��2��y�L�hW9iCl~`�g.�I	�4H5k��<��d1��OyE<�[wL��WX�(���}���g+u(�)�c9Vve�1�U2�\�@���:�W;<\v�4/1��L�L�t��-H��t�a�T�9�a�0����b�v��u�]�ѣT4�p�]ٳ�n:��JK�p�ŉ�6��$n���*�7"�"�����m��O1�eXk����qmwPcl��"�K�2��ݻNnV�B<�Op�ӭ��hqb�e��2>6���Յ=6��(]��S�`P.�}΋л�܋�߾������������%㠀B�,�P&@!ˣ���Ɛ�H�F2�@i6LW:$$�!����I�2Y�"[��J(��NsY(1�4-�ͤ"�3�`���
%�b#JfX��2L�BF��B0���	,�.nA�]�e�� ���P�1�)���M���S��`C$e!�C\�3bR1�J0���w]	�v�S��� �����4.m��L0 �awr��Q  �w)�Iw]#NvP"����d�`MBF�҉�0s���&Ca)�EL1�.dэ#$�&	2!%�ѓcb(#)��"���JBe���0�"�1=����?�ߗ�X�'j ����y�h�O��}ֳ�jV�ۆ�K�db߶��7��&�t޴��sc:�픝��8�M�5t�m ��"�C��R�b����m��,�!Lt�����,4�wjJ�4hpe\��Y|Z[�7书��a[9	q]�i�T����ܗ�/���������[}��F������+繷D��Ӫ�֜�Thª!��l��,��s+���C��`t�w�kqm'l����kfziB���x��>��	�%g��[���Y�������ۤC��&H!B�lI��+6y���3;j�ޞk�fIN(��W�jG�/g�ñ��N5��]�{5�5�]��Ңj�K'O�J�9y���-.|=M��,�Y�r{*drU�L׊���PHU����.Y��֧�#�W�-�ίCV��.��>�9�etݛ�я7��mn��2q
�maU\;���\�}��+-X���o+4�ZJQ�&/oM�]�v�}y��i�U6^�Ǻ�8��ԃ`y�(Z�R{w�/��d�TI��*�M�"]#�{6��Nr-�m�t�O��^�cn�6[xUh�4lΗʞ2�g�s�Uo��V�{��}�����]|�wq[W5�O�t4<���o��q���Q�j�yv����F�ݾCZ�L%�S�->
�p��!h?�QRp�څCe���}�K0a��T��=������-۟Y�ϻ�0u�5�ez�fGd~:ny�A�$��Q��l�G�jd8��w��{M�&��U�����x����>"=~_y��C�7r�uÛ7$z)�:l�xv^�r��.������E�?�H�~<�jV��)-��M+e�t/p�Xaݛ���39tM�=��NєY�R���V����5��5�e�-
��X7[��bH��8\r��eƴ.��r?�}n`�ɯ���]G�aMj�ܾ���{NE�+� �p��}��C��kh;x��f9�־��<���}r)�V3{P����lgA
 ��&%��6��;�e_PǞ�v�N���5��Y�u�B\^ت�\�Q��8�~B��8�n{{�9�Y^�37:QWFOHܠ���%K,f ����]�i�����d�j)uc�g��:fՈ���]�߉��;	͸�ٽi�E��pC������Dm%e���܎��zd_Wf&�}���ڷq�^�'ֹ�c�SWbP,-{�<�Z�m�E8��̢Ԍ�_M��+_j���󿠩x.��D������ݴ��+��3�2���v�D=��V�޸mueE��H��1V�6�3����b�����=�\[����d�\'���P�k.;ʭo7:Z̢63�?����z�_n��֪�3���9�:���ZFt �swOu�����-j��[�7���Z}qgT.ª+@��/4�o[�4g'���9�k����9���Sɼ���z7�X�ps��]����z����&����`$��KR�R���ֻ"�-N�&�`,ɫ|\%B�������,9_oLZ(s�+�펐������o8�n,���-�Zn!��O�r���S�%1��KE���,�vz����|ҺCK�I�uC���r�zk��Xs�j�hbZ��8ܴ4�,JW�W������R�n�IUއڡ�b�ǒ߮�z	�u��]YM:������/�s�,��T�ɹ�C�Gv{�3������� n��..@g��3��#��͙"_˒w淐��m�:eB!OJU@O�v�-�����r��7�B�qǝD-�	s5���a�p��Gk�y�J��-��|�v�oFゞM]jپ��t�Q���q���r5�N��q����ض��):a�^}��͌���_[��B��ۖXe'���5�VT*�	�}]<��5f5S1�c�緳O~J^쬚�N9c�ڽ�ak���`�}������v���fu%�|�q��un*N�YD�ĸ<{|���u���������w��\��%�臯�(�b@ }r��+��{Hs�s��x������������
z�T8��l��r�ZǋYȳ3�e;��r�hn��Ξ���->+��_Fv�I�Xm�����������A����EOz��[�G��Eie��|_=.�.&�#c�ߺ���h,xS
d���a<��{��%43�i��b�S.��t��5V=�L�(������yE�R���s��C;�1:�J�q��,�gt�̣���.}�Sg[x�T��k�*+ò껐��9�	�x=�P�Z�;�n�MVy�h0Z�yTI�ٗ+~V�\o-�Ś�DQ���:�M����Q1��,)��t���TIK����T�@��)g����oW�pNm�^q��:n�XR��
($�@K��9�E��k[Ǫ^a�S�JBTn��잽s!�Q�B���~0��A��gJEP�+��ם݊�!�O��[�֥���I��_6�Ӗf
�uU{tխx��Z:���SR���!o���e�w�
�*�U���%�g�
�g�^3��/\�����:|���>�I&�)+��2f��-yɫ���7D_������G��"�y�O����ԙ���,���WNbMlփ�{�KMƻFg]�:���_{-���l~��kqʵ4��d�f7�pv��r-��!W;bMNYY�΅Y���G�v���%���C(�TWZӉ9�k�5�x�<)��y�7��P�\ h|-�:�Y���ǉ\XnZ#���<�IK�[HP)�,'�xc�s����}��{�ͱd�RoNmeqv�̈́@ݪz{�2 aE�
�W����ys��<j�+(J�a0��x[7[�wgn[PD߶�k�^�=�^�A��]�{6��7\�b��E#T��7��w"����}WX��_������짏���[���cM?lw���T �vU�+TJ�
�<}�wl�<�-/�ɭ6i�Q����"�s�DS��Q�8����h��׾S�:�^���u!z��������C��R7���U������f�;��]�v�4oO��s���hx,����[R:�x�ƢJ�L<�3�z��,��^��ٲ��ǳ=[N�κv�wKܺ��p��>�I������9^u��{h<�	uxz��`H�ns�Ay��_���ם�߳s��W���G�;ub�!�~�R|_�I���ڮdV���Y�p@�c��f�Y�����.�.��r�����޺��G�ԅ\z�hho}O��\{}q;~��a߷L��<����e(���:2L�t�d�)̄e�o�h!���3�N��v�Ը������me_q��R�h��N�k�O�" yО&&W���|}��Co����*@��I^P�H{��X�T�������^��1�k���x=���ne�����u��W2�Z�������,�ٓaPc���ˍl�y�lN�>��a��ucT+)h�����x�^ ��nt�Q9L\ӻ���(�8��s�rv�7������@_�w�~�p���ә�ʿ��ٸ=$LK���WmB��\4����Ǚ��o�HqKt�C�������h�_)d���êå�x�ڮ)��_�x��c����r�E��<�i��=�}�d߽�������̚S��9,s��;�W��8�W�[�����=S�:.6��·��P�����w�3_��'<|��{f㏴��\ẙS���"����y��s���օT�:-_���ަ=q�w��9��(����;�`�VCN�G�[Ν�A�T�#7,ר`��*p��s6�u'tø��q��:�w[ ^�W��u��O�e���T#�uٟ�����BY�g��n4�&�]e�k���!�� ;2���ڼg�b���JWW��Wx�DJTۓ�����pY�h\j���s�P�]���B��U"+{�~����x�/�|�b>*|=p5׉�NW��~�\?��qݑ}�Z9ǅ�I'�&P�����C��w1�g���<� ��L��.�����C�^������x�q^wX]j6��,���W{��a঳�R���A��Oh�M�����x�7��^�
�J��J���vv�1�,'�,*����2v~!�N�z�)��X��Ce�ӫ �wRs�RP�񖖾�Jj���k �*����f���PĊ�RZ��$�ZF�wd �ц+N��.\;7���~�>x��>�.:�V��_�޿�=Ln}�>=~��w�Q��lc����{s9��}|azIf���O��`�}-�WS�o8Pr�X:<��ʌi�y��f�{;,ur����>8o��\'M�����d�� jPf	-��Vd#PѸ}�qS{;;b8z܈������A�!�s���~�8�o�F�e�nd��@�A��2�p7�/��k���3{�X9���f'y�=Gй����[g#�;��;����h��s$�J���*XJ�/�evow�vw\�b�9�F�)��
�mW��z|���L��|�h�$b�sӸ�9������ռ�9p��K�V
��f�����J���Dz��]Ɇߨ�~.�|�F������� �����U�'Ћ'�2c��J���m��s�4���j��	��E��L�˺2��瀞����RV�+��`<�4X�{jA��d���N�W�tڹ||��W��:���w��}��m�;F��}	���z�-��޼�����ݨwY^F�K�t��G�0w�/D�mcS"x�qRO:�9�ZԻ9�Rр��]Y�[2�� ��m�\�Ӝ��J̾��e�JK8�X�޷J+�^�\��*�-#��W��a���j|�9�Vɨ�vw��j�SA�U��^���諛�I�h-��w�TrEF�$��Ë�V���>��ld���N7^�;�PU��s�ù�9}>N�L�4}:�y'�2���f����ߛ>��2Yò�R��<Y���g��}�;�X�x�d΋��:w��)k����ÙI:z᮳�/�&XwR���H��:1ׁ�t�|G��~+)���������\��繥?2��]zx�Γ�\c* ��qS>F��e�頮:`�Z1��O�w�ʵ�2�����hJ�z�ߠ�j1~[R���O��b�e#u�xSǏ,C����W�GYU���>�.�ջ��vH{fҒ;S���x/��3ĕ_�`�T9���D��_�z�sO.�����K;fgW�ӵ����d{��q�j�p�w���%Ӑ)�,	�7^Z���ݨg�u}Y�����D>�����\U����Y9⴯��:U����ۏ�4̲Ag��θ����d�U�����N��2�d#-�ʐX��ٌ�N�����=�߽���W��3��w,a�5�缢�x��ԑޱ�Dğ54/�s�;�σ�|����W��}�������/��^�]UE�?��ʅ�����w�]�����b�H��	�|ׄ^�A5��;��Lf��"�h��f�u���
nu�t�<=3�Y��G��=�2�q�_.��.0u��Ev�Oi;��+��"��٦X.�z��¾���Qy��;c�^�uX����ע`:s�Rz��7b{TK�����t%Lz����o��D�)�>��2�3<�Ӧ�z��}d����;�Х������**_V��+�io\>>䞌�a��k���_�NxB����8g�@z}��|����eH5��z�`��W^���ք/�"H�uw��;�w�ɜ��Z}�yp��V�����Fz��{#��}��%sW�x�6�H�M(Bk84�����^�3������f���
��߁�\{%�{Ld7��{�*��?^��f���~�ޜ�5�ܻԻǷ�9:N�ΏI�:7�^�����W
]/g�߫վ+=걼8C�wYK��֖sԌ~�ו,�x�wA�y"��VMi�.����Z�
�L��j�^f}3#2�*�r}�s�J��/�((յ<n,�����Pg�ת���ty�����+�k���ownkͰs�r+��9A��և�Z�N����Qi'KG�W:�e~���_8&�n��b��`n��yz�=��{N{���s�p��"�����@�-��ٖ���w���s*��'$�;�*5���wY0>𔎹V��s2� ����3,�=G.$�����>��b
�0�$H�v�����U�h�ڴ��z����ܐ�~���y��k�|��,����w[��8NF�R�Ч4[��3�7`H�0�QW��c����Q�^�^�����1m��[w����Р���ɳIK�\�.�)׏��m�s�q$v�d�jՅe�P�8�P�����(h����NuEn1KQ�4k���,�6��|j[� 8R��&(T.�n��i�L�ڡ�=�{[�wl���� ���f�x�Th�W-N��5��i����|��Z����+���a氳�=�RF��57��~�SbU�2�F7���{Q�E^#��η�ׯ��B>zu�M�_*}\���ڞ7y����:��|;I:��^��)=��fx��*�Hv8y�hI���}w]o^Ir���9n$z��� �@��>��͜_�{h+6S6�|�_g2������+i��ٷuu��%�S���DgU��Fs��4ꪔ�/�ima�ڹ�ż˧v&�
��sh���I] 3.o+����oM���m��y�n�'�%t:�6��yV�4�r\����F`�|D��xn�;P�r�v:��
2�����A���+���+{y��uqrh���w��V��-�m�2��j����t�r)������:��W�<n�w����\|z���j&R�f��U���;�C�f�>s���.qA���{F�[�Л������b������#+1��mZ����؏�Z]��z�#��i�C�X��B�IkIh]>�I�j�񧷤���.��@0�X����S��^��
Z�����Yp�;��bw�V7��P�1�
��Z�k#فX�����N�`f"�a��M�ƴ�,U��Y�x[�V�W4/-X�b����ޭ��Ӑ��0�D���\��hs�I^Փ�tC���ǵ�e=mrT�ˀ�t��ǮI�w`9��K�+.���䣜8)�+;׸�sCжL��f1v�n��[�9�<=�����XT�W�\��}�4!�{�1��h��o(Yxq	Rf[O�ͼ��G.�
�*
C���-�� �.3#�h=@�Ό<-���^��'�sRw��y�Az���b���z�}�W;۴��СG-퓝qX�]Pƈ�/��R��Y�M�λ��F��Pq�G<�]�Hn�x���	͝r��6/R��X��n�P�:5����n�̐�<A*�oY[",��ջ�����X.=�iR�Ov�&����
��-f⣜K��حӟd���X�����+Zm���d{OYwiJ��m��@�-���Jm�xa@^���EjY2sf=ȑ�N�*S�Ͻ�`�8֌o,
���Ǚ6����� ��Q������ا�{��$�M�R1I��H�`2L�1!���R�	�t�F��%�ˠd�ɢ��"���I�a(�FJ	�46���S2���2�;����"C$����LL��M���@$X�Np�nu�Q�"&	�Ԍ��� �d(�͒�ą;����K�3&Q��;�!#d���@�L 67w	�H��&f,�"����B� �!�IIdB��$�a0*s�426I40h�2$ɀ.�2���$����"%w\��B�U��}R�����Z:
F�o�.�?"�*�����һ�wR�aW��7�	�+�'d8V��gLj�Kk�LY�ZV�^+Y9�詟9A�L��;ub�w�9R|_q>:�ڮa�o���Y R��{<EǸoWw7�wxG���A�#����</����_�
�W��z�;�'J����v�g`v�c��,���'_D�����<k�@�F@s ��E���1a\>����Θzw�ën.9S�6�S!OVܥk}��ӄ�#�����'Y��{x���^��t_n#PݾXG
����uW����{-$l�4<������������Y>���!�q�����z���hfG.U��އ���廣�X}��*:��_��{ޤ�<k��C5�:�
,�e��6	�_�Q59*�f���{��u-���n>k�q����ɸ�/���� o����2j�*n�C��Fz��Ů6�=�}����Խ:/�u�V��*��y�~����o�~��bߋ!�)�r�_��sY`g{۵�=VgJK��2a+�Z�O��T�ލ�cםw��!:�df�P^���$x.!�2�K-D�A�G��X�\͜�J'v���	�0��ӭqu�E��$@#���uyS,Kޛ����@������V��f�oi�|��bu^��E�r��\3^(`h�1��Dj���=�'G�@�$ߩ��x�Ѝ���̡��Wz7]}b���<Y:����h����[!!�ˠz��y�M�}e�Y�J>qp��V{:�������3k{�,ԖL�9��֢��C4�=|&Kh\�^'2|Uzˣ��z;o-{�**���/u�������9��� -J��O�Kޓ>��t���pY�h^��=qs�Pۙxh�T+׳�����q/0߶���Y�h_�E@h�*�r��r�}�ˇ�+��<��S�xWOj/�e8�O�{S���ٹ��>u3�B\����a��W����|}�>�����;�,���Tfxz�ǭ	��zo{(�{(͟E�H>�<�
E��T�UL��+Ub��~3�z�܏u��1�h�{�"w�׵_BV+\u����$�L�%���H�_Kjs�Q>�o8Pr�X<n�Uo�����-8-�Ԝ=�m!:n����|i��0�_ź�o�W��&5X�\��>��QƮ���ٝ2s�^�M�Dzv��o�Hq7��H�L�:�K�D ����1-��y j��$W�z�m{kQ�f��#Q�r���9�����h7����.=9�4�IaIl���'����Ow�V����V����gF��6�
���W�>��'����>bp�6��{9x��P=x6T
�mn��Z��wU�k�t��]�z:�A�;��Ć�̋^$nS�ӗ���V�ںG^�}�c>᫅M�u����R��&�_!�[�9�p��#:�3����@�S;Z`�;��|0M�4�R^wPzqZ���+7�K��&��9>�9o�����f7��`��4�~�Ʊ*|n���U&:~�&��}�pw���i��<ŭc��J���J�~We�t�b�{eP�a����fۯq�ަ:�j�	��E��'F!xL��곭`Zq���yJ ����V�Ɓu��<���(,�])�y�t���c��p�^�:����m[7���UY�S+O�ޡ�7��M�{V/�*F^�'k�p&F�����/9(5�u�&���n-��`��t���x�u��ȗU�'����~;C�?�K5^8�(?XA<� n .6�x��~���k����W���5)���r�+�{œ,���G��9dB��:*�t��F9�ٗsO{8�7��ҽ(d��.��.G���`+���t�|Ez���j�z�f����Z�k�|jq
�Y�G�ԣqQ)\A����,I>G~�ty����:`�Z1�oz��~��Yu���Bܟu��WSa�j1qmK7x��f�T���F��)�ǖ!��n'�nh���^_G�.�@�c��[;��#��SҾ����%�4�����we�������e��*�J�Oshy���5�¿j�i����4p��w�T`N��Gz�gR���=9W������0��pT�0wR���#�E�ʞi�Qlfc*�I��'s�2crY�����;��t ·k�O��^G�0��k���}�t"�.�`o��za<��XGo{k}��C�y���u�7�R6������� RC �1*��|������w��n�gj�~`��_�jǑ�~W~�ZG!�����+�ꑝ�fî��s��sp��E�f�>�|{�xq�L�c˩`�3���(r�׭���z�����o����De��c�~9v�zK�]�2pתHj�Q%yM	g�q��>VG\6���*>+����Uu���Q����.�ӄ縺��9�|W����>l�^���W%��ĩ�\y;#�)����ط�����cH���'ԉ�}�>��3q�S�\�_)d�D!����պr6�x�n����+����޽�[m�p�^.{h?9�+�~�=7�_�����;�Rt����pvp)oT���+*T��}�qW-���W}�_μ�y��k��7����{�ţ�ˎ��ߣ`�C}����Tw�3�N�VW������/��u��d��i���Ew���]�_�Vq��cT���4윶�~X-w;2ϡ�;;s>�l�wS�tY�^'WKE�G�K���;�z��w"[멛}0�t�˲
��a]�I�{ Eʡ0=6�Ê�����<7~��9l�gz���c�)%�+�&�ث˳\m��דwb�Jc<���Z���9ܐ�yk|d����E[G#�d9M���s����!G�����j�*;����JsTT��=��5>�ma��(����q�N��>-�Q���Z�;�iouU��N;Ś�����A�:l���R����յ<hx���0���z�ϦQߺ� ��u��b�yu����q���lX~��ȸ�J�����1�>�<9}/m���u��x�I^5�P�u	�7��{�����}�����CP;��>�|}�=��r+μyH5����s����:%=d=���#ե���GI>��+��[�V*�w�9�yI�|s�'ǽ����狘Pv{�}y+r�c��o��^��!J�H��t�}^�)z�hho}O���N�9�}^��nW�gي��vrmk.�S��]ޘ�@�,�B�*� zAo��%yNdB2¸}�A��y�
15��2�/^n8��u��[�~����.'�����ĸfK5�О&
�����s�j��Lo�ٞ�$�6d������O���&���p�TN��L�Cf�I/��k�������մv�؍�j���x��1Qɪ��y�ؖ ք���0j�x_�_�QtQ���V��'[� hD�$v�Ց3i�����:�&3?y�lM�旴�-{D@'%eX�3(���Yc�4 �&TY�2�|�\�kP�oM�P�*n
΍E���Y���B���֪b�X�E�����b5}Ǎ,�����s����ۡio�wI-�v;ق��\�QH�K�eC�?;�7�_��q�z��123c��2r����q��QJ�ܦqt{�MϾ7,z��ꕧE�����zSW���ϵ�+�s���EU��?E�F�����L�3^�>��t��|J�1�6�9>ӃU��{7��^u��:�d:�t��WUu���85��䦁�o��g����<dew���[���n����6��s�WW�6d����_o-�ٝ�J�zC�k+#�X�9ϩ���'3���Gʡ�eV�3��Z���*�<�Y�x�^���W�
� ���d�^����>�{θ%�3�I�s�P�]�gcr=�����Vf'�=��Ez����*gO�;��7	���o�ˇ�ʣw����;'�_��q��Zs]��q���s�L��	�
I�ߺ�	so�Vw�����|}�"=�~+>�;�.��J^�nw�f�;�����e���TA���X��U!}wR��4){���yS��
���W��g0�ٿGw\.�>��d��3Ĕ�H�_Kjr]D������o�}K��̦���`�e�`]���(!��,n:��s�(���Ek�iơ.������_d��w%��ۢ��'nE���<����ƞ�F�(��V3�qM�*����=�������:�[8Y�0��XK9����#�2�M��]'�ǟ�����_���7�~�������`�8��o�W��P&�!Lي��]g�v׳0z.���+ޯ,C!�ב���&���q�&��sP���>�'Z�s�;v@�|��;�]���=��G��|�G_�߭����>��OV�q�z��Nx�9�X�Z{�ޯ}j����Q��!�==ԅ]O���x��Tu�j�'�>D������d3Z�>�s6�*�yo�:��G��W.}6fc��>=�AF_�q����Dz�~Wrb�~�'���� �	�T8g�v[�U�M� U�1�������큓���1R�ތ�u�5���5Ua���G�u�^r��ә�-��s�=	�
f��|���C~�mH5>%F}���
};�a\�>P�=h�
���yVf�o��y�ז�C�W����M�,���nZ4�{V���x!j�m_����݇�ݺ�dI�'�t��U�]W������9��*�}����Iˎ��xL;��.FH�^��r��]�NVUi��O2Q��������d��>�Y�;�Y����v�q����<.������Z�1�Zz�T�� �p!^\��p �T��r`U[Z�Щ��3�pSs6�u�ؔ0�7v!�v��e������' n���8� "ua�tl��</�E� =��9�Gl��%=v0߽���t��]�i�6���D�~��p䤸[	h�י���,���<��^��u�]*6�(�U�w�]|�\jڞ7|JW�2��EL���A��:h(�,Ҙ���z=�EO���n�3zFz���ʟJ��o8��ݍx�ttU{�es��.�>���S���B�
!�m���[�R؇���FG�O�w=�G���c�r^�"If�g�*��8�a�#.����e��/ҷvп[8�%;}qV�ߴ真9���D{��UHۇ�d��r �:Z+<����e�5���J���]�ڰ�ȯuG�#��H�s�i^��*����,�Oa���EyP�Nӱ~�t� �$G{���/�Ȅe�p�R!׭��޿3�t��ė�~̜���.�S�&�g���H��#��'��Q*u��,*[�F�BJ�c�
P���+wNVj��t��:��}�Q�9�@�;�&azY�����7r�MbTǽ^���̑S3�[}�<�즷���j����^'��>���h�R
,��d>6}�����옢D�Ss�xm.�D,洪΃�T��aTHi[{4k�a�K�U��C��_�Ր��r�Oo����܄V�<�R�w}p����n��jN��4��gP㚒���j1�mY���ش�rm����ү�(:����M���;������ٓ��e�>L�z>��=���^�jO�������4�34;�2}��z��r��V`D��Ifyvp�h�s�}�=���)|n#:������F�P�q������,\#��T�y�F^��\}^�]��6;o�>������qY^�}���/������\״�|ߢ���z�
�k8� S�J\���3r�_����3���'��6t99'@�?�ĺ��W�z�'Bw^�Z�E�����&m��~3�m\ΝE��fa�@�"��Mi��:�6XՎ;9���e*]Z��4�J}h��&VE:Cx��R�jxݟ�0�ឨw^�G��w�O(��N���¼(�����#Y^���1�^�<yHs[R:�x�ą�y��z��q���H%yyֲq��}FS.��,�uP�}/�Yy�u���_K�A�8Kź��h��{�KK��Nop$�|w���>	eԳn�X������>/K�t������>7<%Y��Ǟ�µtK�+��,נ�ޣ,E@)�����K��CF7޶��pk7s A�~�VR���y5�R}G����g��M�|�i1�[u3t��.�Ի	ЧS���J�i(v,�H���Ko@���U3�܏��{�8wI��Ӯ0� ����;�e���������̫���<�p�F8��hX[���Sv���p׾�w����Y,�|���=�I�+�s!a\>�����}s�{+���r�����C�9�hs�����D��z�Q4̖j!��O�]F�>׀Ƅ.<(��t�ͼ�w���5��s�8[�����R'�3���{ޮ����s>�V�����~,g��}���[��9�G�Q�;W�w\&Zbc{���O��@���^ w��԰x�tj!Ls��Afߥg���>���Q;բ�.��QH�+潷��w&���2n=�P�&F_�Ou>݌n�9{�ս�빓��>��9<:�)��*V����+>ާ��j���0���I�C�ݯ;^�1~�=ol�x�L���Qf(����O��V���cםw���^G���z�R�}k�h�i��y7A9}�yo�E�W3g>����N�qY^�%΃��{���ER�{���s��ԩ}>�^���k+#�]��޳L��F�<v+�/��kŤ�m���,��=�������O�+� R֬��W�{�g��yN��/u�q�vO\\��6�"���=N��G���,
����!�E�_vnVN˹ۇ�J+G6�߉OnἬ�V�ӪWP��KV�|l-٭H�A�z���c��b�|+���V귙�m1:E�{N5��Y�ф6���M��s�u��y�c�W&��J�T}�ۉ-Tc� L`�ޞ� }=�����b�b$oX�W��t+@Mb*�S�����	�CA��Q=Y���"�ؕ��e��q_t�/=L�ޢ)K9�) M�p�Mu7S(��Crd�ݤ!�[qS�N
��K�8%ӵc�#�]�o�G|�����l�E�����m�׌/�+�6�kWؗF�� �{v��拮ʚX�f*�E8f[�^l��VPך���;_�ķ"�]Z��s�2��..mk�N(b�Mm�V�Vc�U�I��)k�������#k�@�$v%�ۖ������ʡ��T6��{���˖��㙋�ށF���d�F�m˗ׂ�@4uj纋n���s�mS�{�o��59Af$j�Y�n��v��X��vӧ�8� ��qS�d��nN(u^I����qB���Vf�f*\�B��ȹ&|��$9�OO)_�;H�ǳ����dKU3^4MG�1���q�-޺ߢ�1`E=��I1[޵�>�Fr���yV4�[HK\�v�4�/%Yo����Z�aY��Җn�b��{��Q��,@\j+�����r9��5�V�����;-�oa��~ջS/l�	���[7b?P}Y�����p����b*�;���閝 ��2@�I+�p����[�GZ��zkF�V鸇Vi�ۮ.h�;#���x7Lг��՛R�����}��qց�1\�$33(�6����F*ER�iJ��T+x>8����{-0��m+Ds[�o�#��hڤ��[�D'��LA��fdT�%ձX�ʂ�W�Z\2�p��*fW)�P����Y9e��w�s;c0��i���b��X�����דt+Zq�m���y㛎���8����2d$Lku�؋��9�U�`�8������xܸ��
s���#)�:>�,�sGv�r��9Wج����-�E�;��1�`��\L���p\�ڰT��wR�Eu�8�q�V��yJ�r�rɕ�M��m��+�wt;W7/����WՆ���j�Q�,��[v�K8�Ȯ���Bfq �)��B�,uw5NC����T��a����u5���'�S�qsTS�fa�p=���С͔0�uZy���\�[�V-n�-�r|(Q|N%{g��*��C�[�*�7Ɯ�/l�ORĝ���ЭX �\�V*Ώ��C��(M��������;��UwʏZX&Ј�A]�=��G{U�=�E��3���[?z���sҌ�5ms��]��	̭X��&F��$��.0 ���F�w!ϨV�ܴ ��zWe��	���
���f^擑��;DK붊ρ':]]�Ҍ�
3"�Bb)�L�+�A1L�Ƅƀ�dr��L 3�#$�4�
(� 9�D�D���M f$20FbH�4"Dl�1ݸc#K�H�Xb�*S(�&�b����wWL�2�&"(�,P�a$�#32h�CA�DJI"����J�4�$�dę�cd幒��"12��I��Qe0�B
m��� Kr��@ZD�D��x�x��39(wvD4c)�)9�^.�#$d��R���/�$��
2F�<]���$�@�(C�*���Ɉeo�*���c;�M	v(�nh��-Y2�G>��t�vLuه�ea5]\��D;�w"�0S�1�ܮ�G�����a�*�7�>��}���p��v�.�����>�3x�}���S�+*�V{���n��I/�,:�L���L�L\u������χz��O�������ܝ����߫&.v��=�{CV+}c'�x�+�QA����>�F�Μ�v�����R�X��]��.��q}�/�/��G��G�[���Y���J�2���"��[S�,����<�.�z1�K�kY�3>�CΚ����W��<��HN������'ƙ9T�`�\H��گM�U"�5��[v�o���癨�����+��h/��ב���&���~�bi̗( ��8:�M�����w�����~ ʛ��^d#Pѷ�Tu��l�}����==Z�޾�9�;7���y[�#]�<���'G�*{����?Kt�\T�:7"8���Tu�j�'�>D������G���t�"�O�+��F�5��zoĊ�\��3�U���47/Ը�%O�^�<��]Ɍ3~���7�5��=��k�O���w�&26:}�I�Y=P2a���a��koE��������?���0�F��;ܩ��22�|]5�z/��E��Vv��t1��s�ӫ2�i#A��=��.k�����c��d)�|҆�;�/	ɋ�vK�{^vwg��Un�dHrG���{����G)��X�[͘ �|�`��։p�d�{��V��t� �*�m_Z�l�=	;���L߽> ��ࡿw�����d���aO�p׸��EN�m�z�;Ց���ט<����lpΫ�n��s�~��7�z�7�Ջ���{(��f�ێ;����[��wqwL����q����!t���_�DK�����xw����PV�/�C��8�����W�hl�y�B�{>`�^��!��ÿ���%���wȗ4�|N�zw�d{�����R�ɕ\v�o8�z����.�r8r%�[�	h��_����Y�`(�^�n���3o�����<�J��>�9�;����b�mO%.��Q �.�|����4`r/�r#G�]{[�s`�<��C_���RX[�X�T7��Ih�_\��Ur>οn���0{f��ܯ�]����+{=�#�s�`_{���s�D{��c�T��|2K4�P0�5���X���f,پ��Vb��~� �y]TJ>�o�*�ӿi�9>s��#�o�j��U�� �.c�$I��@t���筬�����!��	RetBڰ��w�qW�ZG���;��+���f�n�ʥ�P������]ɣ�ӲLU�T8eFe3��ުQ}������y	��gb�[����)����fBv�b�@I�:oX��z	�B+��Y���/w�\�/��U��og���@��,;�]F�/{ݯ�z˒STl�azupӶ�	��һfe��|m�u��B���Z�������s �A���ͺ�`?/�FZ/���}I�zw��B�^Ȏ�w~k.K�p��@7��T̊s%��U$7c������Ӟ�܈F|����9xeeED�OǕ-��`���Bs�Ϗ���&2�1-rz��/X��/��n2定��n�9��9��owG�gj�8'�R=�n�O�<g�w���+����z������QՑx���-�n�;�[�o���>g�7�=���߃󚒱������4�C3B��eH5��y۱ީ��2�v�۟h�>����s�wn}���)|o:������k��7������,m_�.��j1�z��]��s=�<�A��V6tzr|3a]>'��~.3�\{>�5�1�ߢ����.���X�z9w
��be�����F�f�g
99�3��4�{�NQ�f�~'WK^�dxd�Hd�Y�_�m�5��s}���j+���T�g
4��`����W��~��5�5��@y]W�`��!��8fn���s׃�j��O��"�&V}N��/�((�[SƇ�HvT�e�����uϢ����e뿺��9�J�:�{{+a�9�S{��K!�ʰN��i������kI��=�߸��(YA��3n�6;�-.�k�Fs�m��[ŁX��֖-�O��ݚ��Y!/y�����k�f�p��淳olen)���m������T��<�o�d_��{���c�}Hxqy\5�#��<M{D�y'��YW��N����7�E|o�\	e󪆾����t�nD{���yׂ/)�ͦEP==�(���y�uI5��K��!*�u2��b˩f�۫m;��)>/�G�O�ޑ��ȼ���:�j�o���v�����@�.�|
G�z���_�
��^�4��n�(��>ؽSV��o.82�#�9:U�}q;~��aŒʀ�@��H��|
��~Wu�Gz���3�O�X���#ӽ~��.&����7�TM3%��D��J�~zȊ�)ė�i��+�k�U��kY�f���{��XG���J'��tx���\�����9�L����%_���eigr�ww��V���^��qG�ڿ��<��LTu���I��(8����ր�X;���:�ru�j�����zI��2�o�ӂ��Z*���=G!)|n��{�ܛ��/�ɿ{�x_?@�~���L�O�=;�&��"��KNIZplm��
�ާ�ڼ�y�~���^h�an�ۍeE��n���4��'})8	.�	
=���6p���vְ�֪@Pٴ�.L\z�\�z�r��u���V�A�S�&8B��V�-m�2�6��u���Z�=<���֪���{�g:�÷�G��(��a��Y�v�j̫T�,;��#�T�׶n#����>%FkFև'�pl+u��}�LyR����&tk]=�6�������t�##}����V
���n��d�٘^���w��;;^u}ޑ����b�ט+��7~ U�W��נ�8�k��V�yR2��,��a٥m��>�����ue�r�:�=^�f�JD�L �� �Oyɗ1����!{��S�z64�l9��G����9�<����>3��uH�G\�g>=>��}>'�9^>�]C���Tn���ߣ��}������
�Xh���OTDσ�x<��)���З/�4��7���&[����xt�4r�iHn�s�]�	g�ը����,���A�2��ȱu*����F�Z�kw�8��wʷ��g.&A��P�G���_��=�]o�{If�g�*�� $H�>��=�����L���v���	��a�V�z��FG�W�[Tt������~�\{I�9Q�p����,����T-�}�-�����#>����d9��=��RMǷ�#�=T�ә.zq,�Q�U ˾6�4����������/������ѻ�9W� }'������+W���j���F�q���;�%�|;[.��&͕'�ؒ��|����%�1W�E�W��)�ҳ���۶�9�b�5C�o�6�S�Dȁk;fb�n�R��{��	O����X8��3�j/��ކ�m���;��;���n#�������/������:+�=tg�&ǣ�-=$LK�!R_��^6�
�mW��z|��.���$QC뫭�gz4���������E���W(2%�x����5�S�mz���f��ȱ�����g.Su�}�cП+2n��;�Ldo�>�$�Ћ'�>�>�-m�ͷ^�V���k����|�7q.�[UcG���r1�G�T{��\/f��{jA���d���an�8�o?i�]����/���>e��lp�μ��n��u�G���X:m��ו#4�q޾�^��C6����t4���a���;���"K�p��~7�j�2%�{IȆ�ü�az�
����<�Lj�4޻��
}�z�9@�ۙ����*��į������{"\���3�=-X�^�;��^�\�Dסg�}|�ƛ��N��'�]�t��3�Q~c�+8�����&�iB����z��,�՝�:��6VEy\od?_3����Cĥ�X�x�qS>F��e���ꗕq�17�D�g�;�>�t63Uf#��(�1n�W*hG8�Y؊ܭ\�Ņ�ĳ��X�}C����йI���'��E��ek�L���||�^&X��|M�����O#��"�j�����:������=��Q�483n"0� �����]K3+�?@~���,b��~+"�Hyau���[R���OW�a��T��y��w�������b����u¼��j{ף#�'�;��#�{�Ǹ佤@�,���%+$<��w���m�rkO� x�P�(ϼ|��%��o�*�;�����=��#�oڪF�?]�x�S�S�d�ѝ]ޭ6��d�<�<���l�a������W�#�g|W�zN��:pe�7*&��=M��*>�^�uzj�s ��+f@>n������m�:��`� �����VUm{]#�-ޖN�>������Nd�_B�!�DO�W�Ж{�9�o�=J,ܣ�v��ǽ�^l����v��G��ώG�wĿ	����JF\��a{`Oa��}Fc8�OU���r�4z������]�z�=qN��~UR;��x�g���3q�S�\�JY=@�|K��阧Z��Y]W�狻�nz=��V��۞g�#z��m�m�d?:�7���ޯ��;�R�\l�A)�����=�;簜���~#M���t��r���/��u����w�5�����]xOr�u\ܓ�Q7
���8���)CW�B��wڟnR��j���J���b��=�)�.�������`���B����)�..5�;^L�	Hh���p��wy�i�~9͋��Aй��u,��E�v��^�`^��{���#j�RZ�n����;�9n|
5%�t9����|O��~7�u��g���a��������2�K9���{?,�*�����Ǎ�8P��͉�ѧCة�:��Noк��-VND���3�9y'7yWw	�=*���sǗ�V7�ը�ʝ(2s7�0�O�b�kO`�3�ŵ^������Ǻ����U�+�k�����9N�+>�Ho�3�gM��3�4�23�s���Or{ђ�Y�z� �� o�d_��{��~�<�������C���5gpp.��A�Y�{�����p��;�Q]C�|���>�,�>wp�z��=�|}��~S>s���z:�I��9�}˱:;�Uz����*�����(�yS-φB˩fݺ�W;���O��s>�ʨrg�٢�V?$g2|p���v�8��@84��ʌ�$)@�)޺~9��ԅ!/ʄv"l�;���E�����z�;�'J����v��v�<��Y��U�= ��E�J�{�5[����s�O3�W��~dG����ίQ�.&����7�TM3%�D@n��1��/��s�y~ۏht2�����D.Ȥ���}�/�2>U�ɲ�nz�y:��ļ�]ݡl;RЫu�S������9�z���eE�W��x qM�eѭ����Wl��췱�h�=�҆�[t�Z�\��sr �����W0���^����Ek����"�"�	�5���o��ȏO����tx����p����9�L�mG��k̓��[}���<BG�I�J����v�x�ɱQ��j�&��R���x��f�
��K�3$�Q��X�WtW�B�O�|fy�Ӏ���e���9	K�5��5U�c��d���3z��c��8��1V�M߀�~5Cn#��(Ǌ����Ӄ�+N�����Y�O��W�7�-�F����,5���M�97�z} �ǽ{g��͝�>%PɆ�mhr}��u���*��=9�Է{Vo�=��!��W�#5������X*�ע�ü��icv����tЛ|��ګ��=��r�X�kɟT��]~ ^�^
%ׯA�n���=��
����enZ��NeIt��g�v?CJ�����YU��5+Ĩ���kVE��/zL�c=ң�u�g��hz"���������x�4���~� <-�Z+�\�:�O1�r�E	����T;�L��ޅ��Z���%b����C��/���SQ'_�p��Z=_�T����M�w���˪/����ݷhvn��y��i]�85y�S೹���T�ۺ�.��ۧ�@$��l��J&�))����ܽ�"��g;��v�I닪�BTɷ�)-��'����{}�tY7�����\�/�<�R�U�ɜ-���^���w����#�ݗ�����岲��<���XXe��� �|W�T�>�k�	�l�q۹��?�\{���^b]�7.g�W��lpϼ����I���;�v[��%��x��`X)�_��TR>{��ۻh_���#�u���B�?^��>�2�#ʎ��'C����$��2 r��U�����j�o����%[��p��|O�^b5��Wq���1�ב�z��o�o�G\z���j���7�S��/�v}�zG.|끿�|}��4n!Q�߭����>����h8�����7�m���*�S�����L��J��6zH�~�*�_��W��>B��W�5��ߛ�}@�Y��kz���p��:��xցNm�+�r���/B�j��?�H�ރWv���Ugf��ηۏe��l���URc���d�@�&j6+�a�k�Y=P2a���a����O�A��=5G�׫5ގ��^�����B~��q��=3~���ׂ��{jA���L>�e+���ܯI����Y���/�W�t���q���~3��á��q��3~L?��pJ�mϾ�f~���P����ЬC��/�$���sMVʷB��|��h�C�tB�\����A»{�'v���0vL�3��j�(��ޚݪ]�,��Qp��SR�]o�CI���y��Ր�~�-��=��mo�}�{mF�؅e��ѳ(�v�"�m���i<�����u_LD�Iv%�Լc��
�Ivw(q �c�l�z	�(�ନ���]�c7Bҵg�[yxvH"��[�����b��q��,�sN'L�s�����rQwi�R��O�=��$�$i����A�}�r�3|�8�������գy�5wN\E���-��C$~m �� �[�a����"��l�����C�z:L�um��P&�٫,w�բ�VL���	9z�ġ�o�z�Z�k%��3%��Y�˯O�Ѵ��ͰLeA�Q@��%l��:Ң���,WU�Y�l}ET@E�0_>k���ci.R��je�s2��vȸ8k���0R�`�j���Uwد�"����[�K�Z����kMk�PP��Y�*$��2����c�:�M7�_q��c�N�5̋���u䭳�We�㱼�g��ݳk.���!�6� �f�9-"��V݀-�ť�ɕ�ˠv��Ə�l���s{;������y���������pd�"�)��n�Rn�?IQ�@��:q>�r�v1V��<V�-[����U2ųƈ�N{�1�oL0�s	N긟/��w�O�յ�Ws$.�B��R�Q�)��[��̀�X���4nl �(%.��7�`"���_�����rYZ�T/d������5��}Z�A����w���s�6�Bh�!޶jg�W	�q��Lf�-��5�g<Q���ˁ���������(v�w.m7 ��[9t�W9M���Y�w��mXo*�>���6"�����6�,��LW��S����j����b{M�C�tE\�`��6�rͷ+tp�a�k,hX�;Y�S-�Ɗ(�U�6���%����6���7��pJn���$Ӕ�ůػ<�S�%�ͮ�S�p�&M\G���ѓg4B��K��@����/.��g���y+vNv�f��G��bN�a�j���(X��� hvC�<O��tϫ g�_IW$�饚�.�����!` �Aձ�[�wwe��.��K�8E�Q��`#]�s�N �&08ǣ8_C�;��&�LtЋ�8N�e��yB���l�\c�v�F	�$M;ݴ�=��f��o������c�ހ��i���O�!y��Vt��-v>54Y�n58���<�1�J���;6�9Mbq�X���ْIRn�ܧxu��PL�������N��;�wx�h���+��ڠ��I�C�d�m�	��բ`v/�}x�m�q�
��#�'v7wu}*RlѸ������sQͩڬ�̰#�ٌĄ�Jl���� �   �6���X���y�2ZH�$E;����w1�C�ӭЉ Д`4PD `��-�1��$�E�F��1�:�s\�;�w#��M����.��+�i!!0�
&�B��λY��@h�v��nc]$��Jwgq�1F(�l3$�"#+�H���S)�`���$I<t��LQwt������&�V5�1��cZ6�I�$3�vL�K���r;�1cx��E�Wc��t�nD�y��#$�#@ıw+���#r�wq%ݮ�C���n�Q�� ��@� 9�Gr�ř��Y1=����#"y���3K�H�w��a��73���K�oaWxF�%' �V�[Z����&oTwX�G5���� ��k�!��kV��F��
�g�򇏁s>�[�j}�PW�lf�~��M��ht�f��=뜓�x;pV�����jW�G>;.-��DK�^>&���<���F{ٜiŬ�]�N�B��7��gE�Iӷ,e@���N�4�yN���4���ԭx�����+����+��VSW�լ[S�����b��g�S>D�1�-ߜ⫵�1�G
/�;�3��O�ez����Q��e���z����ݙ*����yy��s�I<���)+WB��^��	�����j�z���Pj d�\T^�E�jr������$�0�zz�]^)]TO�;}qV�ߴ�y���u�>�22bu�[rpm �;5
��4�/@8K� w�d�$7^erڰ��w�qW���Y9ⴏ�'#N������Mώ�u#<�Ư�25
�d�끀�P��e�p�R	����$<۝y}��{k�A�}��9���=3�O���L��D�\B�!�DL��4."����x��z�1`�3����,c��6�8�
k��h~T�n�OT�N��1o�`����r��f�ss׃p�)��*W��V�*	���uYʒ��5���Ya�����-�;�֖9}��-���7f+B�C� ���k] �v�CB���g7���]L8@ͭ���1+����\�~U�ǋ�,��;�^x�l
�ۨ���f�����5����{�Z�]��t]��BTǯ�����\Cn�O�<g�w�����,�����\y:Ӝ{v��wݯ��.A�~[[�kaS9߄�N��ߙ��~uro�~�=7��~�����Ι'�F�oR[W��U��t�T�������[�����<���3�.C~�����}���egR.���_�&���h�����Ǐ�g8�z ��+:��exm����Ϸ���u��\��u�{^R鞥��+F��cЛ��^�z�
�������3�����|?o�6t99'F�U����{2nȷ5ힳ��������|�B������W�|VD{�c{>�_#��:mN�0��<j,�@�0=iJ[��_Z�ύ*���k��\탑�2�������V���R��������}�ަY�<>3�*g����n:dx8�z���^���~�<�ԇ�){hI����p�{&�3�|[l�^�ދ�|k�-2�=Q�#q�.�p��Î��
�t�o����Th����H��g�rGw���L�ߤ�^���UˍF�}�^��5�uu�% v���C��ws*�	����S0Ug���wnn�����.O0�1r۵�K���ڹ��:�d��X+�8�	
{�����8qz���I[��`�b���pi��jЕ��p��H?|�s��İ,yT;�����!eԳ;ub�����c�%0�g��TH�]�}����6ϣޒ�_��p��|}�ˀ-�,	�
P0<6#�t�jE���3�.��ܷ��홟h�C�hhϟ����):U�}q;�f|2K5
���"�`�f�\�RS~��ݻ[���s����_��Zdz�팏N��v�Ը����x�ޯTMC2Y�D�^�ȃ�F�g;���8=&=4�(��E2��n�|��ߝ���D��Ώ{ޮ����Z-��aE�ʬ�s�F����C?���v�3*���r�ew�)�*95^���� }�x׀�Zh��s��N{+5�F*5�԰Y�tx�����K��W�]/��%/��5��D?;�#uN߇�Vz���{K�&O�ܨ�}�T6�}�%eN��:�zpz��Zt\F������������ű��{����~��N�g��EzM��\{׶x{����U�j�ևq>ӣ(x���z�d��ޱڲ1b�՘)�w�7Hz��xbu���~��/~�U��7ע�ü��q���fa{ئx5C	�"+����� j��=]M�P޲�-OaU�bU4H�`��
�O���[E��j��h����,�H��6�
&�KԶQ��}�9����e��T:5����:�p]�&���5�Ž<�a]�u�3�:�z<�����z�m�T0�jNwtu��#�V�%N��i�^�_�D���-����83M����HL���n�����y�뤯�ۋ�̜^��n�c�YU����ĬLP�� �J����F�O��G9;txƩ���2^gq��T���r�Co�a���B��U#q�.�}����'+��6�Ś��5o1���q�s�E'q���S�x]��z�P�	��g�c�ȗ=�VeN8�;������=���hBtx�9��VW�ǖAu��2��7}$�,	ȱ%J��=�dN*ܧ�o���3ӅR���~3�z�܏u���ǻ ���@�,�<IUX��+ݺxl��m��b�XH����Ϟ]D�v�t�z<�|�?*:U�{i	�o��d�㴑T��s}��,�u��< n��H�%2��h��+���yb�k��ǽHq7��H���գ\���[���E{��NO����H-���>�����>B���[g#�;��9>6�/z�z����5~�kPW7E�>���6��C�%�U-���DĿRu/����+��!�{��Wc0�����$��d��Q�V�yY�]��I����ֳEmb����4>&f.d�y�zȞnѕޝGE��N�=�1; ��z*rn�f�I�\C�g �ޠ�}C�n��nh�|
	N��l�,���v�`��/B�]�X�͉_���}�L��#5sȀǙ]Ӌ3�6g�'М�'�=3�'�N��<Hu�yj���A��^[��*���Z��G���W��r���ܦ�tz���#���L[o�d���{"�د�}�I�E��&A���(����EZ]�+iwa��:r�׷��j�����\c�L�{��eW~�M���~'�mKQr^�׭Nea]����/9S�z���ܯÅ�u��d7U�9�C�n3�`�oj��Ԯ��˛�f���n�pW����v�f��G����6j^��K񿳭_�D��i8�xw�쀽�4g�FyW�&����(����jg�3C�`����2TjW�GˁK|�=��ǩ�����8�>Ԫ�rZkI���}�QY���Z��L��w�l�>h%��_��(�1���D;�/ݕ=盜����U������ϫ��V}M\od?_3�jx�Y�)\c*�,
{A[#�'ٙoJ��������/Mc=L�9c?S�Y^�<�żE�;UCb�$�͉2l�>�����W撝��<>2�����q�t�<��,C��^��p�x�D{��u��Ǹ�K�A�m@�?����o������Y�9G��R�����k	��6:��1E�9Y|��kz�K)����툱yX�d�p��m����b��sٗ�����V"�疈��OPp��M��
�������`��eb��S�ǧz��L�{%e{�y�}��p�0����t	��PV|��'���늷N��̟9������W�w6	��}���J�g�WeV��p����7>l�[V8�����H��@��$�*f�ԝ���u�ۆ��y�ҽ���f��diAU}2�� �b2�'��+���n�������t���G�z�����}�TN���dT9��*��DLI^SB�=�V����S[�r��G|���|��mW�=>V|r=3�%�F���ۨ��e��&�s�#i�.���x5�=�]F�2�>�J|<����p���[n�O��|{>f�@~��^ZԔ�M@���W�y��o�!�����un�����Vo\>7{o�>~urn1����{��8�Vi�0Ukޙ��`�G�*A�s�z��4�[^��q�=�vz�F����L��R�{��(��a�R}�b{�,!왾>����N��VW��+����/�:j�ґ@��>�bF����9��J�Zc!��]���w\~�{��;�#㳤�~�:��Z�D�~{�;�-��݇F��[t���Y�v��7��ߐZ���~��OW�j���PM��AN���V���ǖ�����	õ��7����S���}3�eO;o���gz�iF��|��bJ�>�r�`ɂ)y�j�L:�qwx���x��˛|^��:��=�dxdK���;����U���>̭��<deyA��|+0��گ3�o����L��.L��#�W;`�S�ʗ(f�~�B�mO�mA�n�^��Yo9��9�d�x�v�;Q�T������C�����e{Ӯ/�ǖW���Ͻ^��8�3�Nj^����+�d�UУ\���~�у��9v&�����'��pT���n�=f��R=�}y3�<8����.�s���2��)�m/y~��p?�Ϯ�K�e;Y묽���@�YL�V�{�����W��<|��p@�FXJG���I��m��u~�{7k{0��n�*�^�4c}�h*������ݳ d�T 9l�;9ȋ|�m]O�Ϯ���׎9#ķәς�޴��y���z�;cޥ�߷�����`�eÏv�O�i8��^���{�������P�m>XGo������>���o��p�"}���7o-��wEO�})�3�G�H��W���j�����G\&��}�J��kr���]�8�B���N���f�HN9��q�/���p�.�B��ŏ�M��i�����]rZ��q��B�"b��yl*��.�WS�U\E���1uw�Q,�]<���Na��|����{}z�^h��*S��%�������<վ}/`����p �����] k�,��~6zpT��e���9�R��^ۏLm�-�;b�6mg����/d���2n�@w��j��O�d��a�5%������ݷ��F}�js*����opk�}yq�޻���7�z} ��׶o�>�8n8��C&�Z��s�W��繌K籛�Z�Of�!���u���~��/c�V
�V
�f�}Y;�ۓ$���&7��o��%G�w��1Ӓ��S��]lQ{�~�נ�u���V7�s�C������K��>�\�j����H~r�ݸ3�PZ�wYU���R�J����֬���^����{�Ϛ`	�����~��������!�Z�I�JL�5z�]z������@w��W�;\'�=O=5om,�J·�w<��������aF��</��$�L��3��L�L_�n����c�t��l�廛}�}+s*|���`߶����{��V}^wY�u��2��7}$�,E�7�C+������sۻ�Zh{�u>7�Ub�!?_���7"=�|{�u���ǲIf��$�7d���+��N��.z ��u��,�/����o�O����ɀ��gfڍ�oS�&�h��H��|�'y�ʙ�x4Y�&�m+[�8P0�W�/����zݝt���g�����Y�+�:8^���%C��ͅu�|H�^��m-�)6��j�����=ٙw������G�*}�N|��%۷�(\C��ё���V�Qҽ����~�\y�!�vh��Wf�t�}s�Ѥ@�3
�z��%x��j7��+��W�!��k����ROj;d>��2��Wf�vi�5B��+Ъ�MG�K�D ����2�p7 �>̄j7����m��5}�G�����5�Ue{]#�ۆ���ՠ��޾���ә%�U-��=$L�R�5���c���/e"��o�{���W�=�ԛ���'�=3�'�N���"�˞������U���=�AsQ�}��4�N/��^���xk��^���#��]Ɇߨ�O���&27��d�E��2a�g��(�F��>��x����Lz_��mt�5�,j�r�T�}��=3~�����h�}��wzR~��N������د}��Q����
�V�T_r�~3�����i��P��X:K��! ��{���x=��p�����7fVW��R��9���R��}��B=���[*�����>�S��e����_F����:r|}e��S����~'��qz��R`�/�Ix ?k��u�61H�D�n�>6�k����1�vh���!0"�9Ou������v�S�tlN.���]t��La#p�@g��xh�7�ݗ[y�v�mv�ӾL)�h�I�^�i�c��j�gr]�3|��$�3�ɜ&������qoJ��[��J�a3>9���w��QQ��gB�8p�/�L�W>����#�����t��o:���|T�\w�m�^>+��VE5q���|�\jڞ7gĥfX��u�N����=��YW^[[��X�u�]!�M�9htƿK��^�<���b�ږ}���T�M?*處ؓ�ټ=ě��񯌺bI�;w^�<� w�z2=�}��=���l{���Qb�D�7ݞƅjؚv�IGÉ/LÁ'ʡ�c��q>7�\U�w�9�'�z���M�R�����lN\���ﻺ�m�w~Ȁp�N@��K`7^e,���uE^Qӆ�:ʾ�R���>s8��?Iҽ���z�٫�25�8�� ���`?/v���u������v-�f`�Q�4��g��ٌ��_�ߣ�=�߽��L��d�R�!�sE�#�έ�m7��S��3ٷ��%#���������x1���>�L�y5����e���^�.���o��YĚy��?�pz���54o.��,�E�}d1p�Q	*d��e�֪0��DG��m���V����V�����Z�ۭU�m���Z���-U�m���V����Uk[o��U�m���V�����Z���-U�m�Z�Z�u�����j�km�KUk[o��V���������Z�Z�ͪ������ֶ��Uk[o��PVI��]�" ���` �������N��E*�TU�B!TE��
�IR�PQ(�I	T�*���*J
QITJB�PJ��EU�T�U�U ��D@��EU+�T�
H�хkI+�URJ�@�EJ��A�tȕ�J$QR�RIJ %��E!J�**QB)T�OcIJ�-)*R�RU���RI$�[ �)J��B�IAEEPUB RH(�(�d�D$��  T����a����Z�j½t�S����+�. P��h�eL *M�m 5`� �fC@����j����$�P�x   �⍱T@�R���QF`� �F�Ԙ�ѣF�4P"�EQGF�(��th�:4`�� �9�(Ѡ(Ѣ��0(��ѣ��Е{eQR$��OX*�<    �N�gQE
&��QUD2�*�i��)��EmU�
&�e
�K�*�*���A*�J�-i*JHB�/   ��@$3+ 55L( KcU@�l(U۪r��h]� ���PnEj�5C]�n�:h���hu�uEP�����
�*))/   ��5v��wIwl*�5l%e��SB�kl����w4���M�5]���ҳ)�3s@�J�	���[4ʖ��5�t�vȢ��"�#l��  ��%SJ�d�`�5i�����T3v� 3H˰�ܢ�i��,�٥��F��Mi�뫸�5]��WS5�Ӱ〺n��Uf(�BB�l�I)
�<   !����j��v�UX�iTF��u�J�a���4v���kJ���ݻ�cl;`t���7e5�Z��إFD֪vĒ�!Q(B�W� ��Z2��w����4�VЩeV���ѩ�� 鵳`�٧w�렠�h����F��1A�kU�ݓ���J�R�*#���U*P<  	ܭ��uFt�ۮ�ݬ����K�J�� �]�j�:
�S�l
�5��U��)U�'U�]�@��k�t�V����!D��Uk�H�*�(�  L�l[S��� �L�[���p� �md[V�F�P*J�j�]�*tVي�������t�����2&��6�)�4��JT @��a%)*z�d�L�z��L� )� ��@h  �~�&iUS@22 I���b� 4<R�b���A%��"�#޴�	����,�y����k[�����{濠$�	'5�P$�	&�����$��	!I� IFB		���?����2�z��g�詭�n���%O�鹨Jdk"BP�3*���0�ݦNb�t��AIݥifaI�#eGYY��;�d�]��0]Ku��>��km@����w����2��t�],��e�uZ35$�fd��+8�yt�m(y�G�t���M�x+(͕qi\Zh��,�u�`0ȣ�k)�&]:[yf�wjmh[f<���ښs1��9a����A��N7^U����zV�ILŦd���x�.�B�f+U��:kr��!F�J���X��t��u��C�2x��@8���*�D�f�1�xc2���e�m�]�ӵ	���l�R���v��0��\�X���s1��h��bn�ݬ�vuO�ו�iWd�2�=�J�)�����r�ÁmE��m"���b(����K��*܂�jB±�Orn���u\j��թ��T׋�4m�N'��e�B�L���t�%]elw���֝ dhH4����D�iM~��m��rm�;�0�@�P<��Vbyu����f��L[k],����X�ec^�:G�
�{�1���z�n\1����b�� ������[���JTͥ�*�pH�R��"�WY�.h�2a���k{�Rm8���Ҙ�E^֧��D�-L8@�u]�x�$̗n��1:�����չ�]�IM�YREG^����������A��;���*��x��i��U�V;y�0��	̬�5�����u�F�84�6��7D�٠A͘�Nm=�ڵbFb(��"`ǂD��\T��KP?�q��`�w�wq諽�亼N��Da9m�I,$�n�utZZ�^�$�q���n��A\R�k�<����k2����2��5�1�'u��_-������۱��ae�	��'�H15�`�#u�j*2}yA��{q�9%��^]i��/��6�jwMe7k�R�n)�WV����k߀j�s �/FZk-�&U担�̔ �ER�r��Y�Jt5�ѝ-U�p��
7��'t�5��-WH�$�Ȭ��2��k�ͅ!o.��1<8��W_m�Rh��
�p;QeX��-IAo��9����_�&û��;�d�T؈�V�D\���4Jڗ[X9�dȈr*@���V�`l%�Y��6mß<yP��@��=��؅�#�4�6n}Z"Қ�v��h�8k*�wv�&��-�ba!����5���no�L�id�U&	̙�#�z
�d����V!xґ���D��2R �ẩ�kL�$��ŻKoi�h��@�]�V�ڙ"����ԛ|ݘ�1,��b�fXwj��wz�n��^iӖ��2�57�&򠼦"�^��wִ�v����ÑF�d�h�WSLfY�(�����@�(��ܹr& ��г�i,�okv����H����BB�X�1SS+6H!�nXWn�P:iS�Ccktahǂ�[��	n[ٺ������*�:`J C�T@�	��;ԕf#$��
Q�nLy����շrU��-��sT
�]�J�/N��n�JKt!�&(U����w`L-b�*�{(n��w�pTP^	y60�@�hbf(�'W���;����k��Y)]�G��YNmH�km��]X)�ifLL�\D��.�AT�c�Gq�5mji��
�a���+(=��:�	�a�W*,�m	��A�X�[�%zḴB�i�-U���ۥ�o �����e��q����9
�!�{�.�ͧ�~45�P*�FfZ�1Z���M�AS�kc���{�,��e���;I6������VV[��xh�Zë�C��(R�f���a�-&��;��ܗ�����Y6Ֆ-�ĭna޺M,��)�y�IAYB=��v�����0^=��)����1n�Z����rҹL5p� յf�¶��֣(ѡs]J����2���a��MV9�S�ԣ�7�Y���0�4Q���(��M켺���j���[$��[$���� q���upd#���yd�mE{��ZM�N��'�VE�����Nb���`e�*Z�#��h��m�Kۆ�ɓ�\�X�>����l��V��-<U#�se�ջ�Wi���vh�6��$�ׂ˘Zn�%� �u�U�B@��"��dk��ywn�VT˸1Z�zF�m�fE�������Ӹ*��J�i���x��d�6L�{��P�œ ��m:W�����!�#��� x�n���2�5��0ЅYڊ�3	E����2Ĩ����J���6�F��Je�.�Q�2Ǉ �7)�6�U��R�ٔ�2e%9���a�Zwcte�&0�LgעI�-������9�����4��w��t�<��<h����R�A���t���+I���Ԩ�ۂ$���r�
W���շ��׃a7�B��z�[1�e,��ujC	@�B���h�t|�+:@e�!��XX�[n�:�;����e�QV)��B,����(L������:i�YPW��YE!�U����C�EJ�$N�w� �^X܈@鼘��M5m��0㩳M� t��8�Q ��6�`o;�� �z�3Ph�+w�ԹA��+�q\S&{EVē���4��#I�������ӗǸN!�o>�f�2�r8�����zf�e�%�����w����4ȸ]��nɫ����R�f���Ԭ��.��n�[@-úhn��x�a�򙼘�L�B��kso�7dj8���VT�D�a�m:n��U��v,�e�!���d�&cW�t6�x�K��r�k������ �rɰ2��x�I�e�/0Y4����7�2.VVf!Jc��h�t����&��e4R��x	��]���	0ث�R����܎�p��ܕ�(R���2r��fn7xR�WG*J*�[U6��a|�,K��N��*�Lm8��fl3�;D��
4,$�ӥr�hX�(��*�o��B3 �NH�7�8��j�̎"�)e7KL� �i��h�R:���J�Zcv6��Ӱ��lԷw�]1.����/��QU���0����a�r�1}��i,
�P�m�/*�ok7j�i:)�)��n��dH+wZv�s1X֨�j���v��V�۬�Svݷ��o%Ee\CC�I�P��>F�5�V���u�	�am ���S�aY&��݅��.�e��V�K�����J"��4v��Q!��1)f+�@ڴ�e�M]�t1Z�PXAYzFc��靌���P�2̷�靂���Cp�n�Ҁ6qQ��ײ]kwr�����s[30�G�ul�R�����X­��v���԰�=�ͥ!���XȓC[3eX�v�Ù�!����^������R*�	"�i��IX��8sn����,�c-���c�"mB�8u�srh��b��� e�ߕ��9��r�J�J9�ú�L&(�3����n��|U2�+0oJ�J�h���N��r�%���R�T��s(VPM��6l*�"�$�et��3Z�N���6:z����V7%Yѱ�X���vv���`���Ŗj�V�+]8s5X���ř���1�������v�%��,?�j����`p����I�\�
��v�>)�yxr�O#Tݚ��5V���28Q��KnR��l,|r��eT"�[X�,Gui&kT�mnác�V��GrD��w��Y/U���ջ�%Z,�:��G�73+r3{!B��s43�ZW�A$��r�����9�Fd�5�Kvh@��cvPY�#���������Y!�p��m��*ʆ�I`�a4R�ܽ�����	Λ��ڡpe`բ�e�j����k�z�O��"��5Y8Feʎ��[����q
�nP����dSj��h� yp+ u�Zɘ�Km�O0�9ô�Y��DMˢrބ4��uok �/���w@d�1����^3�u-m����Q�E��H���خCZ{1Yw���1�hc��ѣf��jʓ&a
G�4����)��m�b��V~PVҫ�k�%2�bE6�H�.cw[��9��e���L��; ��i�QX�e��ԅ��5�F}(�d�X��CU/�35�x�6������	*1�s3 �yj����Eڠ�2�.Pc]!���^�"�ה`��e��c���z��c��Э��\��T�o�$լ�v�f��j�P٫��5��`�wG^1�&�h�-fkf��Fh��2�Tn��6�v�dF��<F��V�Zrll�T �6(�1Wv�7�#��LÂPGQ�v�4�0G(���\	��1tc�O7�{r��$�m�1�6�F��Su��Q�{-�U�r������ַ��y��70\!eG��Ř�E}���(���+uG0�3*����՝-��%�(��VJ��f��Y��Fl�kb�ii�JLˬ�Z-Йu*12�ɶT`�)��PU�j�[t����%��b2�bj�b,�J�]�r��5f�TT؎��Gp���t̙6��D^'PZk/0��i�NL��(K�ͻ3)ћhPf�;T�j�]����O"2���-㗘v�[E�� i[:�1[�|Q��6�F�F&4��fe��P�YYu+VUĨeb�i8�����k^� ���M\�wښ�F=nZNDcR�Vn+U�,#B�^��4�٬6�]�b̷f��L^��s7�Hk�n�ɧw�0hT� f��ӥ�����o-B\�Ih�d�8+QE,W�l�I�P6�;Tm`{��j�@��)5i���m�j��X��:.-j����u0�![[��U��7d�&Xʁ�PF��
�`h��t��2�&�"�q�c�V��Tku<��6"݋8�
9���)�Yu�r^;�5��h�.-�Qm��NS�F� f�����86sA���{xR)�K�a�8`T�[1����4/2	H'�MJesX�H���N�������Ďkx14�^��բ�uwF
��ո%���t��le[,e֚�I���)9t�@n1���t%
$2ʻU��ܖ�0��c�m�F��p��ܶ�x]���[�:�1i�������6��X�[�i^%[�,ʰ5�F�X1���t\�tA+/w4Ϯ��R�C�j���̳F�L�
A؎^,كvh�r�&��-���8Y�/�F�8b@Un��[�9��p<WG^��M�2�e�P�e��Y�����ƍ�_�-��`r��IQV��e
�Um�B�!��˳!-�bҡu�����7���{7n�c%}��ݶ)�8lj֖m���ҖH���T!
�.��^�o �A�0�S9
5(��6�w0=p���v�Uuw� ��#3$�톮+��͂+h�8�AP2$��o�5�n[��U���9f#��k��C/$��,���a�#\���SfmV�[@fA
����Ct�0c�J��:B�M{0˚�э��j��GkvȖ�V�:����Vln�kh��=��^�+b����l͋V��x�JF�]� =��uD.��t�խxBQ1�%��Mef����i�Z9y�\�M֦+ �Aō*Ǻ6�:� ���ϥ�t���J�n0V�m�3sar��%�A$��qc2�!Br�w�=Z�ڛ��#	��f�Y׎��Sj������/2�^�@��)y�����Y��2�X�e
m'�Y��dXj�9P$@Y�n�nn勍Lu����%����mb�c�RRR�8쩭��,�a@�Kn:�7Z��G���E�NR��o���j��!���I�5i��Alaϛ&�>�+M�q]!{�&����&eKn w5ԣn�n�YW�p5id���k[jc�ˣ�4��d�.�5��AGp� �N�S�ǡ�z�+�1���Ur�jj�yHۡ���������R%2̦)k�mZ����,���y�--׌��"��̥�V��,�mj�WV���miU�&м�7��Q�aC0�X�`jD��A����]�Y�+ʻrdn!t��DlT]4��~���T z����rջ
�^�Q�6Q�I�rkJ�� ��f���غj*ࣗ��-�]��Z� �T0���	��ӊ �l#JDtJu��͑�K������[w$����w����]�:)`ۤCtqխ������@�'y 2ېZŏ�+-4��U��$��B����*�!x�l��X��nPP��Ys6�x�ܗ�P�v�I%�ӹ6����KN�6�K�#@+�UWyj.��ʴ,V��4���0��Yj�A�j�&K��˔p$��+@�;ԁ-���F�5.R�ѱ�S"SO7`/-݈���L�6�d͕dV`��F�N�3Th�*�D+u�o&�HU�WY�+L�TK7�����4�(M��$١T�BZՠ8�Tv�
��R����`�5�c�~+�R@̇
r��2�r��n��@���*%���)^f.#�AM"@P������O�i�/�Z��b�=�ʍh	�@۵��]��)�v��,x�n�m��j�Q��Vɀͭ�F�B���V�Ⱦ-�����7E(����u7V��9@C׷:��֭�o(h4�IVnD���p���T��[_h�aie-�b
���8Ie���5�kw^�7��d*X�3�`K2$�i��с����UK�)(S���e]���0�#�K�9y{aD�"�mh��;KU��N�o*L��X�/@'e�,֦��4�C-*n]fڈ�p����um��Ɯ�ۺ��{���A��v�C�뢺��ʢR�;2<0��Y1	(��n�g���c�ۮ���P���\�ƩV:��x�`��񦂹�t�3r�A+)rV�����ff�\���Ui̊ ��Չ<�O9�G�5�w-�W���v�0^J��ݟ1�F��h�N�;�� �����,ި�b=��D5�)]r��k��q����8��UړzI�7�Y1I��;cxL�}�:�"s0�۲���h��HÕ˒�ҧ88W��ys,Q�Z��R^ZUm���a]�7X��/:�r]�8�ue�!c��Zۤm�+m���5N���R���r��V�j��~VŌA�ǋ�B�wX��T5��9Q�Kd�����8�s.*N��X�s|{lu�3��HU��E"���]�F��mm�W0v9*�}U� �7����˕d��ʥ���v�F�� ���=�~�����)��=@h��+�VL�MS�왹���l��-��Y6���WY��˔�r�rӾV����7y���p׆�
�����l*��ƕ�\ۚ1�˳���W�k�����6�R�p�N]��&�6��Q�
����_��+~>t<��5�ӷL]�	�FVGۥ�d��u"���yӎ\4��%y�Λ�ņW5�M:N�y|���<x��̕�2_n��jk{���ѡ.���ugV��0�8�U��E=�5l^�R\+ۖT�(,��iQ %�U��zY��87EYl]�y���7|r�b׍p۝0']�]�oҳq9S&^����7�4zW'!�a�v/��X.����,�y��j:gك5ku�6|�Kd�K��[2n��m��Mط�db�t[��	N�$�J�����X�u���{X KїY@F��|8�4"��1��m��2�P�o�N�N�cwCBw��q�= �p`u^t�8�7'Ҷ��2=/R�
R��-q�r�k;M�L@�-��&-vq��������R�OE(�]�w�{,���42>��K�˹��*ܸu�6��w%��*;�k�!��!̶o��
�ܳ���oo��!ԯd%|,\W��Ow2��z�\:f�����aj{x��������2��c�Z���"���i�*�+��sɸr��	Z8��8�A�<���)��T�=2���nS�4e\���1𷴆Pպ3H���b����r�U:_\�<`zm��<\!�����+��"�F��(Zh�Z��]�⦪ݼ����ݤ�;t:K�N�;�C����R�m�2� �݋z��p�o��1�����S�����,��Ai�/G=��S�`Z�&{\�p�	�\�t�n����K�[������n޷�ヒ�I �eq[V�일2�'%3��;o��g��a��p<���C��tM��+j�+�Vz��t�&B���b�5��B�s8����`�G�]��Ԣ��$�/3\;��� �<����PgU��:Wc��HT3 ք��pTj�gVJW�����u�����=1NN�燊�̧n�)۽l�����7�(�$b������tr�i3,P��z����\����Z��7p�V�E����ӱ�X��p��mz����n�5B�D���8���xo�ge�D$-�@�U�1$Ҕ��l�p��8HEߡ���F����E�%/E�{ƨI�l3kf+*p4r�Ov�b�8cC�����l�Y�3xq�n��&���pZ�������t;�Z�����r�����՝���D��q���}x�&��׈�+h���*W)���)��m�vjn\����[���\w7IO�]ʑ�i�YO9��u�MahL�d1�xvf�2�A�[7�G3�V�%�m�,+N�1��*
4���,��]j���rTzHp�$t֛[Q�j��[��=�R�;��S.#�ڭq���9�sTɈ\�u�g���fV6uR��yC�G�̛�we��9��i3O}�d�g�)ݛ���,��xq<��y)�����yA�l��qV]qeT����kPIv�F���\����"��S+(u�뵗|Ŧ��K��ܩ����ݛ�RD'�,���0ٙ��Fon�q�t�}Wh�[�8=�)�X�uZӎ<Z`��;�xe����ME�ɫ:��v�X2}�a��Q�Y�q��jcT�kX�л ��C���5���k]u���v�t٦ǚ��Lh����鱱�!���d��S�E��*�;����Vd�������cj���f�1�8��t9��g'%%ڪV7��J�Љ�Z�_�_^b����R�c_p#YNq(*RB87.�\���#x���|�'�r�M[��E�̩Q>���r����3�9�7��ȸ�2�T	-=��<��Cs�ɔ�)��.f,�49MKpߢ���u�����C&\�R9���9;m�����"]ʕr��XD;h��}��j�X���v�+�զ��']���.>�㛓��`X�P?\��Q2:Z�fY�Ԧ�=����Vs3���nF����:��D[�7���v�g�h�5�)TDK�m��)r��*Qځワ�vkH*�R9��K�D57p��/uT��fZcsvf���=bu!r.��Y��l�+et���A�H�)^��z^�u<��s�׹��v 9�Jm�}XF���`ou�f�hmuL����v���]����;U��3��v*uo7��׏��c��T��RW�����[�eC� �D���b�ʽ�}�0<@�$:�L�f���
��m]X��������"�����(����T*o@dH�sOqd��$]��&� Q�����5C��M�،���&����[.z��	S{9a�"sxn#�w;�~�ml�r�1�)$-l����؛j�Ԥ�ၶ���ۏ��}|��2�[����m������0]�"#�]���vQ�]�1�̮���z�&"�û�$�_Z*��	��+ɟt���c��W���=>C��Ә�w5��H�� �/-.ӱ�"�$�a�B�.���	>�Ί�
��ZXN���z96w�g:Ĳ�˾F�A.�#O�o�._Xǌa���[��r,k��f�'�����;%�0�S.�s��ocxo;��H��}��U��Rq��ovm�{�7�tQe��9V޳�^	�J)޿Y�᳢�zU/׎)r�t/��J"���o�|��.Ǐ�y�Qm����1�Ɲ����-,�ܡ�kn�R�����Ww��*IY�%wPlҹ�ܜ2>aNWqr>3.�4.�����,�;b�g#�l�Ūup��ӣ�T-dݘŕ�Z���gu�����*��H�Y�n^<���S�������aP!��-ci��S�Tp�h�u�2�Lr�R�Y���ws���'�X��"X	�X��6�� 9g��c�kg÷�y��L�x@9U�zs�i�L���!��b�S�β����q^ku�V��j�.�/�Jt�۴��ŌV�Q4���D�yY�mYtv^���`���j�"4Pj�S;���ݝ�:�/�&�*_H��;�<�<6I�`REs'�����)X�n�u�5-�2Ա�5XKݧ�)��ZQ]�M�-e���P�NkƐ�1Ҿbgk�i:��v�]嬐>��u�-�Qt;�ɹX^0�M��l����3F2ۉh��p��t������|���Yk�.�޴
�[��S��6�f�F��uP�������'Lv��e��גa��H�D��3�p'or�`�>��N�r0�7o5,Oy��!��x�e��`����6��/"X��Ě�;�ް:���:�i��#p4� ���*"mbP|�6.��G�C�����MT���mY��+���9��8����)F���QғuՁY�Vh�nT�֞�|lI�#��i�Nڋ��^���J�ɰ���٭�Y��l��L��PNŋ�7j̅��	���S1i���mWV�����}�y�����"���lB'����˝6��Ei��$�r�:d"��>���-�yH�eS՜���Y��{�q�|q;�TV'��b�k ǰ�zp���v����
��v��0��	��uqӻ�'���X��jt�x��IѼ���7xQ�VԌBh����(t�P�z��k�Y�|ÆR���l��:�m�wi#٩>�[�:�X-�;�+�3�L/��
�K�M-����v��6�GˎPb�v�"�f޼�j����"��ڠ,�[¶�1�ӊ�t沏=�V嬮1Iww�t{}A��^�i�mi��6i�ƥ���,�`.�����r�a��N�vU�m�&�Z3�z���v���lc���u��?C�]�5q"ɞ��X�H��u{�mtZ%-G"�yZU}�%[�׳f%��
��
4��s#t�.b-@�R�o)\z�H�6"�N�8��gp�d�vgӲz�]��s6�m�\�Ҏ���V�v-�io^Nջ��i*���R��\3�:Y��X�y9'5�:y�w;6b�����kUe���	�0r�H:ω���8�c�^���[ʭ ��d�I�e����_:	�,��k��⮮��C�������nf�Վ�Ǐ�r��oQz�¤�_Bƍ|j�Bu���z��<��9�ص�[�Q�>E�� ��C��5�eVsM^���������-oK0�d;��
������c�8تM�S�[���q���4���[�Q*P���8�	��a�ha��0��!9�w3��;���rʔA�U�wr�e�s�Iɭ�J�I���%�
�B�W+��=g���,R=�]�������xn�}о\+��.������S8h��om���m� '���AI^�U:�(.n.X��E���c��
˹9+�{M�K�-o\�v�Jy6��ڽ�����v�#ҏ|�^\�t�nc��|ì���ϊ�x���o���u��@��{:���]j�9Vc\h���ɩ��{���*U�P�su���oҳ@G�h��^t�BuWf��]�v���}��d�x�)��-��v�`��m.N����`�]�
}X�[�hӲ��=��ON���q8Į��J�!�6h�lp�Y?pM���'���e�.}˂�L�]ʏ�2�Z��u�Rj�s��֫Os����sm�-��TV��kR=Nk^P�tc�����F\�+��!m���s�	}���9���)ON�cN���AR�C��(k:a�ˆR]C/��Ġ���e�<���8�*Om�u����N�[uv)�+;���4cht���h:���+�7��vvJ���;�^c�&��F�|�Jgd�8ї�A�)U�70Cg,9Ba�X���\��!�L*��uMѹ�:逻��D珻s#m҈�=��//��(T���%.�����k��N�X����.m��;O{���{Mޒ�z�6ooNteG����K���]�����m�h.����"��jv.v"|����5y��ۤy���.�`�X�R���Mv�Kn$�N���u���c(�	�Z�d65-�s=%ۻ�2�;�WB���U
�on�vS�NN��f��w���}��:����F�,k�렎=T+���4,�sz�ˢ
���^���'o��@B!�J�!G@��op��]���n�X.��6V�z\��Z��52(�����pl�Sʽ�9�u�]����P����U+��̤�yu�Tw�y���0T��P��guAe����J�|�U����9nL(p�%�TVDI%��;.T���@�c�@Db�q�H����U��^�+�mg 2f��є��gTF �c��ur�Q���kq]A�+5����o(��&fƉl`U�]4�}���C6%q�5lƛ�{��8a{{�Z�vō]%|jR��p��Jx�L�e���U�SJ㽘�bG9�^�Шt1u՝�CTpC-ݞ�i 2�CTwԺxhؾ�e.\�'1�ԅk��]J�9��WoJv0J<��,@���!��m�|e�vh<��*6��)4b�#���n����zbA�c
g<1�qi��Ǧ���]z%��{��L�#�s����;�[Yy�BqvQ˂�쬔�Sc.�������M[���]���g\�q�G��r�;��]n�oB�;w�����oe��c�T[	�9ڦ�a��Aچs� "�R^���Y�s�SRz�etX���Pl8���A7vқ���"�]8Ѕ�5:�+��E�l)Z�7CkfwȈV��ky�ٴ�����4��G>������.��u6E���5`���|t�K���p��\��M���=���z�fbP��6�����=qMЮ�r�X�ݻ˨�,�0,�C-��Y�%����t�<�h���7ٌ7�����\�v��%6*=�(��;��I1v��b���|tݢ95f����SŠT8�%R�q���l�ҭ���H��ڼ;��gc:�!���`|���0��k��x2�UK-�.z-��1�C����Ki��뾳NSx���G4Tp��<��Λ���?+�=yس����\���hN���E,�Q7"���ٔZ���bo,ʕX��Ÿ�=���Ay��V�u��[Q���r]޷:���jmG��H�P����}7&�滧+��,�]fv"T|[�]R�e����Fuc�iV��c;x_<�!95Cf6��n�c]Y�A�|/�e�m��jʹ/��9c%m4�#�����5F�I3�M�9�ԧ�X=݃ø�T�b�V�� ���JW��հ��;y�C�������-�{ύ�����[�-�'J��n7i����90�%t�g��b�Z�ǽ�6gS��ufm4�J�k���,�;���}_W�U�����}D��$��v��O<��{���._w�߫����{�m�h5��"��=�rJ�i�JP/x�����ed�t��7R^��Υ\c[ܹn�f�{�E�L�g�w.��B�%ʝؤ</v�X�.�sv���P��d:�-qW+����>(Yi��u^�M�2vZ��r�on)�ԭ���V�K��@\��kwKv��JN�[P����&u:�����X�n���Z��
�w&"�˷b*�3��r��v�uiݨ��/���>��&3[��\<��<o_,��A�Wx����� x����Ӏ�p�@��|6�]���e�7��8���E���vU��i�ļ���s��ˇ�K�� 9���Y�5�8��YN��+%E�S�$G�"�)�lً.d	aDM�����sy�֧V��goc�u_n��-ZE��+k[�!�&�45����L��W�8�[)�'8�'-.˙k�_7�*����!lw�lv�rѵT6��櫠΂�E2��zl8�T�|�=�]eU��R�9�l�t��� 9����!SH���I���>i�]�`��Cz�a�.�gB��.���'��7;pU��K6v�}9w>=|[ftzr�Pd�5;�s�D��ԣ�,��L)�Ը��ұ���W ��=V���7�MCqMi�KT�1�1,�XX=�vEAoL�V���sU^�ޜ�(Rj>���[s:��5')�RO�1:깉e�p�ڶ��u,a��̢3"L�]����V�{/�X���|!ǻ�{#X�`���%83�Z�j.���(|�2�S�D�/��(���������y*�]s��kl]�l���'ҵ�e��׬P�6͓�:�o��f�
�;�֘��7Z{�S���J�ծ4�G,
h��Ai�8���9og?�Ir�b4�r鯏v�b�<ޕ�l^�D�W]V���&pf'sC�^�m1\�S[�fWh8k#��˔SD��::�׶�q;�w'�nY���5Wb�&4��AJ8n��wWf���*% 2�Ku� ,t�'%��Mj�>���ܻΡ�һ:�3���$�ڤ����\�`�%�f�S�Y8��y�˂8;9��ս��pi�l=7�4�����R��0r�U������,�ʹ.N	��Y4v���%٨f ���L��L.����E��iXQ�Y��	c���T���LMw�E��	P�e�\���υ ��r��%�3/6U�-�-Z�dQ�7���ܥ#2���(^+R�7�If��ls�w�U�8q
�W��˙�m���B�ir-Qv��<��'f)�a�IC,r��㭵������U�|'t;{�1�l���Ƶ�=���cKn^��i*�'�6a�7Y���r\�v,Jɼ�[��>�R��"�ܸ���YA���9a��'|�u�p�@�����t�Ã�{�����D�ǧ5r�h�����u�����(\�G+bG+��Sc�ɥ�&)�!��2f1\qTͷ��JXkrk���73_k[8���S��y���1-�/�c�m!vc©�}Qiˤ�����)��y*��A��ٖ.�/*��}ksr.��9v�5�	�o6��ף8�s9<��s�[�Os����|p&eM*un9|9,_)��PB=�{G��@�%��Y%��C��tT�k�l:��sb�v�,sW)w�(n��ՖL����w��:��RЫu�	������bjUhwWN�e�۠9������ip͹.��Yhj	!lQ�+>ˬ�撕��X���ɻM�m�����;�5�Pa>�,�΢��x�ُ�x�j��5��������u<�5�"��x9ဲ������Cbs�H��-��޽[D*�\9��֫�$��#�^�����=��@�XX.�ۛ�V��WP�]}�C���x�'�{�$8=zh0y�I񮮄�W�Y/5]�����kDU���K�R��,ηe�5�ジ�۹z*�z�n[s�.ؔ:SI�qhNΙ���A3G���V���%��+�u�FvR:��b�xWL1�:�AӺ�U��%+gpY����*��=f�Y���޾X�F��X/X�u!Z
 �G����騬_nf�����N��Khs�M ���A�n=�����Zs������v]�5g�1�,�`�=�K�ɩM�KI��d�I�f&]�w~˔�#zR2�`����@9�i��U�� ��\i���v'�݌��u�ãP�]���i,��yu���_�j�U���*�j��Qa�e����B!�
���gbs�7w �sK~�Z4�
�&�����(㻫�iQQ�tü��-�n&�y!Y,̔��G�w���b���1�F8�����}�"�ڋ���h���d�}��'ӡXb��R3����.�ř��p[�u��&�"}��.ݧ�d�2�%�6����f�Ov0����k�=3�lp�4fj�*Q�tzڗ���]�P�R�,��R���n��;�Օ;`��.��E�L�����&�7{y�@#�՜��( �P��u��.h�l;�ǜeb�j���WX�X���7l�Ūuu*���9|AU�O4�̬]\�n���Y�%nym\�F�Q`7��}�u��Aޣ|<+^�����YCRK�f	�®�3+T]V[�Eڐ��nE����������kkB";����V��U+E�w����I�jb���@���V�od�g3�EqU8�	�R_[��{Sf���u�-����x��ų�n�a�ٷ}�(&,1ևk��(�5c��*�W ��=wF
��Hl:jλ���@>mB�騃�w�8r�.�N��=cQ����YJ�B3[s����Ғ�:��殆�)1\�:Tq�Z�EN��['���f���W[o"��U�ջ,i��h�t���k0X]k9엀��Veb+g��[��%��,��Il]v�[|pʕy��R�T�e�Zз�l�f��wL��E��d��s�J��]���N��v��]ӆ�s7]:}���!۽��`{j�I9���:وJ	V�J�j�:b�+�<v�N��\M1�f:����ӹreR3 �����w��T�X��,[8�1�$�Ws~�a<�c4�\X�n������ur����BT�h>�ŀb�
�7r���}��u��Qp{��� 9<ښ��|:(Q�-r�n�����uoZ��@sk��jl�'�1��W��B�l�0��R�sS��n="܊K͙k۵b�V�FY�x�ǻdn�h"@ε�[�(Cdi&�[>m�k�,�:��*����n�Q�� �N,��OcL3���l�|<��y�*�`�~Rl����n�c�8���6UiZ��CKuǚB���֗3�.�s���̿�+骯���Pj�n����ȱua����i_N{x�mou�ԈGt�GS�����4,ˠ�P$�*YQ��n>��rC�>,��X(�b�J<l�;)pu�S=V��-�4Lȃ�}������i��;̜��Z�KY��+:��"2�}�T��cZ&Yqkr�8�]�g<_-A�a�ܭ��ݓ�Ǿ7��t��;W"`_:a1Iݽ%�s����@�v�4!�^?�kI�:�,�;��u�ڗ^�gb�q`|��.f��YO�wEv�����w�$�,׸Y"�\��s]��v��`SûQܢ�[��eic	l��i!C)R�;!}��GBc�b���L�yuر^Y� '�Yn�H3I|�ISw�^U��]���ζȾ趐̫�&}*o ����:�gP��!or�A�
��k�}V��%ipO�Ԏ��!j�%6��TVvE�L󶺶�^���ܹ&����ls�2����������u�/{	�9�5Ԝ��Y��%腜�8�f�<v0��f���Z`�+*��`����`���a] �xqJ=���^>0���	Aҡ�H�^���Tn�dގ�'KF��o�'�h@0���In�n��B��9Y���y�ljq��ʇ^�V��9;�z.l�E����T�~M`u�-Ώ(�Ǧh�vɛ�@�l�� ������,���㙻ͤE���F1�t�y||�9�ƻ�(��l��*��4[
��tMQ@�d�gn^QJ�gىTu�1T��;��oG���u��:��|ݺŘc�e���p�]h��⸋�EѢ{�
%w�^[�jA�u=ܧn�S�H��O���;�eMQ3b��r�لR�e�'�v��*#L�ONS��B���wU,Z{8q_+iv�֎F�bՑy�I��y��F��3D�W�!:���9J��-X�k��`��w�5�A��]T��ֻ�,ڽ53���Bl���ݥpLȳ(��L�\H���ֶ��B������;�x�&�������gC�7J����Y�P��$��+Enj����ܻZ�7 Ί�v���5{n]��Z��.�{}B�Sk�D�>["��et{k��p�.?�̱4�4l�j:�����wO*Y��j]Z�7.��lf��p���]Ltv��AX�к�y[�]X/\�K(5%a�����/VbXCE>���aIQ�^e��*�m4����0��Z��zhwݓ�mӻfe�x��@(��H擦�e���ָ�]hѸ
%�r=5�m���H`�v\�FP���X��hD�\g�&�k ���\�)���aW}L{3��֑����5��V����ެns�1������7�z}�q�Ls�&6��Y����G�ouչ�6�]�X����x����R���FF�>3P�.�y����ڱc(Y��Z���˵��qn$r���s$һ��4�Fa��%���:�ii�yڻ���A��R��ʽ��ﬄ��tj���0��0cήH�ܘ	=�����t�g���k{\���K��@R����c�X������ݬ�7����2����Ҡ���&�{�/�\�*ɫn��6�G���[�km�Q[D`�p�돂��O���^A���u˻��2����R��Ul����M��V9��@q*�7U��&�=P'[��cw|y��85��������2v�3,Н����Y�Lsɵcjm��]��Z���h70����N���[좰Ӿ�WJ����!�����ܳ��];
�����8�uu$���7�qv>��d�j�m7�Ud���[��LP{����C�A]��{��d��{y�,�}�
��������$���cC*�A�N���t��b����7$�Z���8*{ǭ棝�en�T�C&.y��%-<��oG�ݻD�޺Q;EרE�5�i8��� 8".�$��pk�Yr��֯�:���z��8�i��F%oz�olɁ5d�2��v(vL��Ы�"�j�	�RI+��&h�9b7���l�d�h�i]WL�%z�i�\�<�j�m��ǔ���,U�{tr;U�ޔ�9��0���.�-��nk�w��o+8�6�ll���''v2Do�6���M���՜�ޠ������:�����Vx�M��}�G���"=���lTܢ�.<���;3i���!�`�n�Q��K��}kwb��ֶ gZ�j��E`�@�w�a�J��+�����wtbR�U�.Q43����)Y�r����E���i.�1,����]Ƹ�fyD*|w�E��7ё,'yG�������-n7���i]��Q�lpW�%,x���-���)ˇq^>��%;�&���>�@���R�ގ�Z��\~J��ͱ̸
��.ذ�EJ��?
�Y�3;`˴�|a�ީDo�JU��x����µ��� �Ju4��Tѽn��g��LK&u�YX�R3Ij����tţnA��;C��{���K9�)G�����o��{$�[Z@m̢�;P��˝�v���,�6m!;�{oWIWbq������)��u��gܪ��s�	�fM�3��܋��E��q����
�@%p!�8\�l�������se��Z� ���.�{�F������<�+�3� �ۦju��ruׂe֤��R��3�qWp`�Ƹ0qY��C�	���g=ŮB4���h��l\�<1h��e�_F�V�@:eb�)�.�UͺyB��=sBaPYm�f[f�0tœ��
_1��ww:��E�77*u� �&�X�k��c���fn��J���m^	Q@�=��A�Q��lS��*cܑ�v;JO�H��g�N��@*��5p�b�ͼ�7�uܥI���u�F&��꽽W(;g�3U�
�Q�������;�e�*��Z7��\��]A�hus�V�:�u�w����R�����6��ܭJ��"����G>�LAY$#a�٬��ZzU$j
�v2�m^�v��c�T�o���Iz�B,	qړNM���"������r�K"�h
��� ��T@\��b�YWEp
�`ۆ]i�C�V��T:�pn<o����IT�=�h�=�^�c#uնKqV�,΂�oq��ܴ���^Mˢ,��J�F��ܥa�!��7�e��v���֚�-��uN�"볓��Z��(��b�e�B��+��fa��X.�
K���i���8%�'U���^M�V n@�[�.V(u��Ԇ�و�X�F�V������D�b1ՖtU���W^�x����n*\(��^���繡vL����q�3�U���$D���u�]�J�������θ�\�C�cUj�Ay��B���N*�(�ٵ !�-�q���5cT�@��b��I����;�Bz�S�=`m��*L��KU��C=��ugsV+nu�L-�b�i�r�to�鮕��+:�F�NG�`Qeu�NW�m�坡|��v}�ۢ&�?}���~y���_�͟�$ I5���~��׌�0�j�&>�%!�Xflw��� q�H�Y=�n��uݵfȜP=��q�t��؆u��7�����ӴԠ:�`f�7�C���W{Ջ_#N�徭�v����y6(��x^�^�5/�G%yX��^D�&�p���FY�2v�N;�㭻���U��.:qI!��9l��)>�{.�T�[��W���΂%�āj-],��3���޾Ccj!yiM��'N\]��#rk.�V�Z�Ѭ1o(nm��b��4;�)�koeh��;6bwJ�s�`l���X��K��d��w�<6@K[�g�/�)��GJ�՝��#z�wf"����2m⵶M��S���W�3�L
���x��$H�R���eh����wK���Ui�K|uG�b��~�ζk�=*>Vg��ٻJ�έ����i�Y������+w�'D�n��n7�i��)�N�s\��k�xRg�����Ҫ�xa�u����
%��n�x��2�nwe�p�Ԭ����|���;RoE��	�������E�.=�G�k��1�����n�*J�I䦋x�Wusj����^<��ݎ�.�-N��N�^�v���ժ��hm�ȳ�T��T96f`)Ր�ؼ��.��R$P��X�pEc{p�e�W��#{�IwbΦ7洸R��>����[;)�\#G�NJ?
���ۯgH�ﺇB���1(�E��Ym[FĶX��mQ-VX����*�R�-J5mF%J�eKv�P�UkVƍJ�e[C�mjV����R�m��[m-��lV(0mU-��������e��j�Z��VU)nYqAF�6�*��32�iE��s#ZR���i*Z[j6�m���e�T�hյ��j�Z�mj������q�0��e��QQC�[Z�PFEYZ���Qf`�PFF�is%0K"��"�m���E�őUm,̵-h��ck���r�UJQ��[e���V��E�[E�T)V��q��9�b%+JѪԶ����QaYZ���J�Qh��j*��F�j*8�\[B���[\�Lm*�F��h7���33"�-��VѴJZ[lD�hh���@ �����l��[�yY%���CTY�WX����;6�.�/�6��wȞo�=��������*oV����V:�]���Nwʹ�z�Z0O�o)���CL.(_:U�c4j Zxk��f����e�|c�.[����^�{OZ�9��*���)pR����VI��b�������;kP�����������P?������e�ۭ!B��@r��!�=%ب-W��o�A{��;�� ��a�Y�ue%e��;�]]�(�^y!��
��ʷ��Y[/tՇ��L��o6��R�<i�<C�4|%�U����z_�}ܶ��I�r����r�V����}z���9M��2�
��u�>��^�}qpwy'���!��!]�ۺ�fq �N����YG�x����fŻ^���~��\�z\|6E����k����f���ֈ��R��3�����`�W����T;�G�FV�%����3����g��� ��&*��3j���2�Z��nfz5OMeG������Vnѽ�/��\MS]�v�{��La�=f���qWN��"�3�[��bs�\Uវ��n�{�����u����_jX]�ޡw�������dI��������e����Y^�=�o��9w�]���K��Tr�r�ɭ�WRc{�T��c��������H������hd�
iM�V�i��=�;k���ġk�&�7��������m��2u����-��t-�c> �
�[��_u�	T��0��p�:����n��'�΄��w�)CT��_��Σ�0t{�RKG��!Z�[� ���1����.�|}[�)�p1���)���:Uk����x�.��@�p�]"�i�٢��'<R�u��~��Rb�U1o��];��¬�������Ga��442}A���&|���8�풳w6�Ra��	�[o°NV��kS�y�==38g�'�>
�;wB�w�9(��Y�K���/���0=��yupr˄����Ʋ����^f��70��0.#Pl}��t��[�1[��fwtc���zY�H�򻧧���Uޱ�3���P��'�_���ƕ���!$�Ӟocj�¨Xѫ�!?"��Hcb�E����Z�}�2�$/E#W�����m��>'�}�|{�-ip�u�g�P��a���c��[C�^�h��krN[a�� }��R*t)���+q(3��>3+�i�yT�]˲CB���7`˄v�Y����j��o v �($p��q�\�c��s)�o�f�R�I<(��)YEc����ռlޡ�������zx[���ݭ�A)r\�/���3#���M�X+&p�um�}O�0#|�7׍+��֫c�|���Z4t9�)�v�����������~Oǆ�v�d'Uk�U��9��>����vr���|`�b�z�ɻ8�]���u������Z�WƵ
޴%:\�&
^q�T���
���ň1�¶����F���hv]�9�i_b�*�u$�_�Fq�9-v����B|<4�[�/W)�p������F�~HS�<Z7O��,�c��c>�xa3�j�]A��,Ô���)��Գ}l-���=��k�C�}k�OeAZlZ��}Wz3䖏O��
��j��MW��6^��D�p2�Ye38���z}[*��`L�����Jb58�T�sȟv�C�����z:j]	�]O����;Բ:c4�q��^��C�Tj���B�U�Eжf�YjzϠ���4vY�;�XƢ�}/T��DOnt8=��<��W���-8,�f<���7柧+B��pW�Y24k���X�i���/T��j�R�N~�T�Sٮ�E��w��)�=-)��m�(�,��Ti�\�]��4��U��f� 	g�^�k��!�Aq��	}a�+Au��+_,چ�[��O��OZ�*�\M>��x�WϦ�X�=�MI�(�Id�ĭWn%�^�ճ6 �_N@bF�L�!f�
ԩ��36��G'V�h�.���l2:%�dY�Ж�+�Yt��XjJ\��4浯��;�*�r唤J*wT���8]�j��d�+��t���nwlgs�Nϙ���^ԓ�UK��:�b���j����m�'��F<�����O:�}� �nG�ۥT�=�z������]�3�f>W�q��L�[��ߎw@/�P�n:r���=t������H�	��c�G[�GV;���L~��S)�е��0��z*�黿S9��Eϛ���[��l�ϧ�G�K~�y��}{��YYr�|~��+-��v�ըJ����t�5�QA��+v�+�r�^�Oޣ6�����z����ϮL>鈿|<����j���q��^v�^��kz�O^��=�{ݛ�x��J���U눸���9�uS'�
�t[2}=��|���@����'W��=�x6���L�9=�K�9��>�rE��=��z�ee>*�s��N���j��������i�w�W���2���OsV�L��ד"A��	���z��������W�*yPK��A�.^q:�]��W2:�c.�`��v�W}*�y]��.��_�^�f�┭�SY�A5��vE��v�\��e���h۞���^�{&��l��7��0zn_�y����6�m`����0���q�uN�oD�oyך[C�X��q�۵+�>U�'b����~���u��gϽ.��r
3ySĮ;�ݚ�t���gcx���*h;v(�� �<�|k���Y"~;���Ֆ�r�Sg7�}���ʧkʻ�Ί^�R%�EN�~�8_ǧ_)�o���_܆Q璧L*T��Ӻ{�ڏ*{�EՕrj��;Ӕ���6�ϊ���}����9��Q��?M�Ku�"��t��{ROU�0�[�2�0����"�`��_�^��YW��ٙ�����*�N���[�pfN��wk}�lO�W��\_v���Ykrw�fC����'��[K��+1#�}K�˜��J�{)|�=Q�]W����ug���n>U%�p��Jnw>��3�?/u�.��m����=�8��%�V;E���c����B� g!G�N 1^�-�dI�f�E��Mp�>�V��y�"W�k1d��֣�`��rY��hp�u�I���ڔ��/�n� ���t�9}X��9��s��k�f���Ǟ�w<G]O�y�r����z2Mթ�i^�UC��%su��;gf��'�����z�؜�G����F�{�h������[�W�f� |����@���ϸ�=��=��Q��+��pe늋�G����0:x��9>䷷�g��ҏp�(֡%w�c����N<�4s8�RS������l�_d��y�:ƍj���'b�]u��T�H'������ݜ��y���>�߶������1�c�CF����:��/�[avg�����0�Ҽ�u����U8%��M�f}^uݭڧc����k���:[�R5�VHWs�i��o�g��m���wӺ���&�K�iUl���ch�X����l����~����u�&;����?w���9��r�9&����}y#}�{�oM�т��ѧ��w�g�T�ןK^������p廾�]cO���s[�.�3�v���'�h�o(j��9<
n�	/�Ea��Z��mj g]s!ݍTGb�ծG�lmMQ�;��=ظ�h���b�k���޻%$/�s:�r�L���֌{ʟ`��8uK0��Sy�X��l(W9�5�R&��[>�4�8]:�[�����_n�i̍A����WՉ9�]�����U�&毢���X�UE��^'�R��z�©:r���z��v�}�y�1��|�=��c���ڭ��_g��A�Z�p��9�}&���ty�0,�[5vw0/�P��Ncѕ��5���k3���8d�����`�j��f{�z�o������(]c�*�1�ϣ����xVN'}Js�kxA���H��[�vj���S��"n/g�q��dɻ5>w�z����o���5{��;�y�q��J��%s��-���Wr)��I�������x�ύ��w�>���N�P��w��eMNs���
T'�t����s܏��y��^dm���;h,��u'��7����"�i�<E�J��O�]G:g���J�U7�:�k�ǭ������=��6����P�K#�k.zj�kH4<�2�����+��gk��?�38�M���qM}��� �o�S��tu:K��gC]O�u�&�ToY�+N,nu��e1q0�r�%�F�+tI-�����ᜅӔ0�x��꼚�9X���<�s�n@��=�SD��M�U�g�N؇k����Y[����pd��{r�ܟ�5U}|��?c>sޜ$�����F�z��H�sH�[�M��,~m�aͱZ����t�������?w���Rs�!pC�ҫ��k�	nto=׊U'��]4(�� �Ɯ�����k&W`x�;�5
�s�K'�����T<�:E�)H�};h�kN�[۬��%2o�w/3��r����^s��KQ���ܧ*���W�Tv��K�}Rl��C���e*Hd�ut�n��+��*݀]7#���r�Ґy�y]�1=\�7��K0��j�Oc�۟��%�[�ݙ�]���Pn:�r���yf�Z��'2���t��g�+�L��t�P�����W�-k|k����r��8�Z�b��1?e����hI�n��ʻE]�A����<��-��R��Q�7�P�b�]<�]�f4�����Ix���Qt�3.m��G���b�ۜ��BJ�ˬ���0|@��{V��N� H��&���Ǵܬ�e8�.����v�!��Ȩv����V���8G��������
WO5���X6l��Z�ǜ�MI��#ͯzM������V�|9^R������J�'=+���n��u*��qf|�ads���۹O������~/׍���Ai�5���w��R����iγ�������T�}2yU
�E�;]�^��gݾw��/z�(֠�]��~s��3���W�fƜ��W��o�.�ճz026_��j�u�ca={*h��ɳ>ssx�omGs����J��l��)�},u�WCcD�0���l=�=ӄ�d�9����&j{�/��;�ڥn7���bȮ�cj�k��s\_���"�3l�Q=�r���=Ϻs��)κy��>x�,��/��أ� �<�Q�� �^���ն��;��J���ge;^U]�gzd\�H�EN�hV��4�Y���»�zjXT�yf�����R���=�N�y��r.����um/{V_hx�)��<�C-E�JAyy�P��R>���-ml�|��y�y�ِ�����?1 }p���f�����@^qI �����C�m������GZi3z�s��2�r�]1�[{E�[�9�yՓ�n��;UN8�O.����ۛW{�=�ws����ty�V��z<�����2<��/���|��� ��wzn����Ʊ��9V��{-5���U�=%n�
���159ь4�����wy�ީ�ʚW:��V�`ƶ�y���ٙ1��T��0��Q^r��#k���!�'��ԉ�F1�z.��ug�3<��<�S���6�/�,�5�MX��E�G����R�����V���?4P|h��Ls�{;1|�ď�\��j�;����Q�5���S��|��<�eh�=ۗX]����׻��k�4��N.���]�pe����}�s���Y�<���:d�ߚs�a^𶏭�3��'Z�����z�.t^�X�u�M�|a��3���NNS���ۙn�Zv�-�v86�� L��']�Vy-tw���;{�߫e{�l��գk(l`k������=�g�D���u[r�;-���4<YJI�f 7�]ڥ2�F��$�J������0_D���;�1�:��hLZ��ѭ���ַb�6�&��<�i�T�\���85���:��x�,icf����9�Ɲ)����\�?:���Z�W��%^����r�v���@ue"܌Q�{g�f`�l��=r�JH7���O[�%���.�{����y]��i�:\:���Tk����K'=�Nө<Uz�.�Gٵg�j������'T�.S[�o]�=��?f�r�!^�*m��6|l+{y��u�����V�{���LS��
�uش!s��z٫�+�PS1]ir��U�>�T��76�h�X��3�IJ�]6����8�'SWrsaв`70�z�Ҳ����K&v�kJ2���y�֋ӝm�WS��3Zy�;����*��F��N�Z�֎tjoq}Z��u���SV$�(vWb����DSDau�$����0��z�CGuNeAm��X%��7/'������V����Ķjm��a�ܶ�����Љ2�\Q���"�����w�
�: tRޮ=�r�����<e0��Զ�}׏��U�'R��ٲ�+�\�ilC�y��w��2�Ts&o�S���S�v��C�3��{�(q����EZ����Pm���ŷ2��6����[���__>61�5rB%4�v�V<�E�\�E)��7C�wME���}e6����këJ��}�r���c�eopf�""��ԫ�ˬ�|�%��5�Z�⫩�;m,{���s�w�����С׭B�s7�1r�����:��ׂ���&'˪�+�q�np	��� `'&�#��u_"���c�z���)mV���`u׏:�����]Ƕ�h�}�s(٭��t��$�Ks	}lc;�r=ao-t@� �
i�=����:�\"MY5��'L�$�/&AP�*�u���(snS����C�ZD�*nR7�ъ��A%���i=�`��-�9��a�('�����6�m��B.��ٙJ�3�y��[;�O���^���C�!v�� uap��x��b��
�^�@[ژ�t�gT���1(���N�����ީ׹pC	�C�f�z�%(2���s�}�e�;\&p!�e��Jޭ���%�*�u�؁Ԅxv!��4NeofTp�����Xl�+�J:��N����t���t`܀:��s�c�Ƌ(Z����3����m����69�d�I�x�+����ޮ]{P�\�ԍ��ЩP����Q�N��(Ոk�c�G�SwDo+gn��2*��G�]<Yp:�Yf��5��e0Rj�� ��t��)�"கe�3����gP�`�>����	-�#i�,U��z�g&�vBΘ	��d}k��^To�?oZ���q�i[DRؔ*YF�hղ�UhR��(ԩij�,iEJ���-Fڶ�Ume�V"�J��U�mkl+��6��X6ж�V�QTm��F-�Q�����kh���B�[X֪Z�V�����--aX����Eb����e�RکQ��F�Z(�V�)��K+F�Ո�h��V�mb4��Z�±�#R�Z5��؂�lE"�-[��+kb�mR���2���KmƢ�0��m�5�PjZ*��[A��l�X��
YQQb��U1�U��Z%-�e���Ю!F9JV��Q-�m�����[liek*�mmAPVұJ��(���m(ֵ-D���T�[ZV%Ue�QV-�
(��J��kF�d�)A���#cZ8�\���\h�3%��kJX�"ʣX"bQq(�fi�����r�4Uf5q,DZ�PmJQ�j�Je���?  �bջ��4�]u�J�FO�u<���q4N������ӯd��"�WL]58#}R���ʝSk8E�ZƻP��K٪E]��}��_�Q{��r�vگ�����Z�r�c�1�k���V����yd�P�ܝ|����uN�y��G�>���U,V�C&��:��z�%��2�z����6_C<��q����󢗫���X�k��ϼY�����o�T��p�S���g��s\7�Ŀ�L��f5���}Ѿ�^T�َ��.`�Q�jt�K��e��^A�d̑.�;ə�a���<�*~�UEqS��؋�e�L�W��پ������^���^z�܅H�')�(ǭ�k���j/|_g����	��b3j�Ѯ�Ov���IU'��w���qҪs���ߕ�A3ϼjn�b��&/#���G�um���9�D�>_k[�z(��X�	�z2�?l���鲰Q�{m��ϳ�P^��Bl�N�T����g׹q{+�1�Py�k$ۥ��;tkkH�K��~V�ܫ�b�����ޝ^�����bt#r�ހ~�I���=TN0$�3p�
Ch���*o�]�Eｗ��~�*��h����6��2�f.�5�[�ӹCo��V��y��:����``7�7�n�	�wa����-�x\Tv �=��U�_w�Jϯ\_V%z�e>V�{������S�UŶt�&��߄W�(S��"�^9� �W���'����p׽(��ty�9��L��(e��-���Z�m�3�"�p���~�M�-����G:u�)'����2���Ҕ���Q�O,
�.�����0��/��xG���o&�~��ΧlC���T�=��nM��=Z=R�G��6g�����<\���p�9 ��-��[�rg�a�)��X��me�������<����CcRīt�~��6�wM��x��sf,�S�������G�#N].볷v<n��/�g����x�eM��l�oM�;��r.Y�(��4�8]�j��͚�3];�w��[�y��V:�n�3�j<�m�9W�$���`=c�ǥT��
��/:֪�{��M�.B����J���d�zШ�_h���ҍZ�
��~Ww�@v�ӊy�d���}�WAH�I.�w�Z�֖խq���U�H�D+Q�w'1��4�Y˔���8c%2����71g��j  ��v����dُk�{�ەW���\�n���T6�9OiT��հ���U۞�\~�Л���.S�ˣ�=�[��^O;vfw@/�Pn:r��tT�k:���[���������ǰNyW8��T���O-�Wo�k�'�ͪ��kh�ս������fM����'?�[tzy��Z�k�}]W��z�ϐ֠����Z��)m)�-䜝ʹl����s�?��z[����қ��%���d�k�{ϪU�D\Y��ad�G�R|mbW��{p����ϸ��9���`���}K�����E�����)��d�"ɜʳ{�������{�ۼ�F��k��'[a��΃������R���7躑�{��b���?QC�h�8�U�U�������=�SDy6w�x��>ǃ?����]�?sKU9^�*v:�hڱ��y��|��
��͠��b��3;py��;�ٗ=Wihϱ����1�8ӍV<�,���j��Ʋ1���*3�ĩ^!�&��o|��L�u�h5sl�n��������U���_A�'B:���%Qul9w�`A�������a}�����{mrWt��ėv�~�����}�RS����v(��mX��v��9x���.ˁ����󰟪�J�N.n�����/��Kx@9����j�Xg(�H���p�J���#��3����:)z���};hW��N�=�sg�7�/c�!|�}sr	��ᱹ���{��]FOh�'���Q{�%��1Y*�����|���'>OO,��'Y8����l�CG�d�	S�;�i'RN;�a���R:k�;W��ߵ�~k����AC? ���`O���A�a��u���IR��nȲo��Rq��O_Χ�l���ğ�6���=gY4��^2J��7Ͼ���x\�z��{��yۮ�I����'X傆�=Jæ����~���8�S~d��sG�"��,�C��O��vd�!�4�&�}}s�Җty��TGq���������;��O�T5>�Ad�?O9�Y8���{��N$��;�!Rz���rI�OC~d��svE&�Y:�L��H����g~�V���w��YS�����z�2q��{5�@�4�����!�7>�Aa=C^��q*]�'�8��T<�r̟2j}��$�����O��A\���X?����opg~/}����<��Va<M��P�N!5�|�̝b��Y=C��Ax��O��2u4�=g��a�N%Bh<�q�����s!N��_�n?JGt~���)���.���ۆ|��k&��v�ޚ�T`y�)Vu9���N�"؈�F,�޷��wY��S��?uvG��Tv]���%Y�yfʜ�ޏ��ռt�:o��j���>�]����5T�0�|e�Ѭj��m��J��G%�*
��l���O�w��v�x���6ԟ�>J�z�2~OfY�I�V~5C�8�����N �k~�!�N�g��'ug2u4�<>�����h�����!�q���t����l��5�N�̓���Y�$��`~���R~I�k(OS�'SFY�l*~5C�,���u��,���	Rq'n��U}믿_�鿸\�԰�ͣ�?D�w?���I����o�'}�d�O�2{�=�'RO�3Y%a�AC�VO�qr�z��8�+$����Aa6�����D}Td�1���~��!�h�V=o����M��M�$+'s�봓�6K̝a���d���I=vɣ���N0�O�IRm!��>ed��OŰ>C��M+/ﾗU멗���AF����^���d�z}���J�����������HVN���0��	�&�9�>v��O=ᐛf�5>矡Y&әd�6�Y�+��*�����Iy��3<���G��UAU�OS�IěM0�c$㼡�N>2�`z��N�C�� m$�9�|��M2sT�I��vw�I��&������)�_��?�2��{}���%|EP_~���
��ցԝI�jaI6����I�{�06���C�f��I�=��d�	��6��`{�0�f�6�OsZu`5�����k*w�_|n����ʫ�'�~氕	�^���J�P6��6�L,'>Oڰ�RN3�2a_�:�Üì��y��4��	��>�;���O鹉 �i����z���]}�U_�����3L�b�?wu�4��8���d�+	�q�d�VO2��d��h�a8��x�ְ�C߼��&�s�ѧ�<fg�y��s����w��a+6ç���d��̜I��;�P���;�!�=d����$�Ms̒�I3���o�2��O�;��?Y!?s9�nk�ny���m�J<��RBfQ�Wh�v�n�D�t�vq�|s��b�Cq�k�H��E7Ӗ;�&^Ҍ`�j^H�r�Vj9�O/����]�s�=Z������tZ����-A�Gι��c5�w�1hJ�>�b��x���{Q��N��ڛ�yk����3z~��>���AG��d��&�j}�u�T�?s�u�XLMw�4��)s�2|���<I��d��q&���_,����Y:���V�9��g�d���}�}�_!¿+Y6�~՚}d��������7��Y%J��=�Ad���d�N �4s�<I�O����'�?{���N�y������d��wޞJ�ݏ���b���Y?2q+�M>��~d�!��a�u�Ĝa鯲��'�7����r�Ad�>�u��Y��8��>�^����	 �g��rm���UZ*�Gӳ�{�I�MO|�+�	��n�x��Lє:�|Φ�冘q�ߔ�?2u'Rl5�I�4��'�x�Xs��~d�
��^2X�g,e���˲kz�W�B�������Y>~I�X�|ɳz��'�{I�Y?2q4e���M3FY�I�T����	�[2�q[�$��u~+��NQ���8̏�߾��W�*�)�?$�C���Y9���w�8��N?$�ẃ�'�>|;�IY=@��'�d�Èh�!�?2u5�q�z�?MXq'���v����l_������uWuT�aRq�iY�}�8��k9�Y��<.��'XO;��X|�Ӿ{�N�O�3Y%d��t>J��'�,�����]�k��7��]���l�^u{[���Q�;��RL��*d�V����'����|w�;�$���'M��$�?$��<�'N2��Vd.�m޹�}�u<�׼��SG�1_h��8�2q*T��8������6��d�V�}��:���<����~��'~���5�`;d����u�M������т�v���/�ލ�_��>�߲J��C��T� ��i��'R�a6���~��~I6�,:��,��������}C��$+'X~��>vϿ���hd�Fu ۯ���/iPu�#��$���#��[���aYpWR�7w�V��FX�^�t4�mw'.�C��鸁r�����y��r���;k��N�2�+a�b�t���^�;�z��J&������Ǻ��,K�9�/܁I9����7;��r��P�����UU%s��=�9�������L4�Ѿd'�Ms�Ь�i���%ABm�B��"ɴ�d�o$�N'�P�?0�f��l�}Hxs0=@�]��;���{���.���ϽϽ�����t��i'y���O4���u:ɤ�w��&٦M5�d�C��J����6�d�VO����&Ҍ'U~�~�O�}��=Fkv7���)���/C=~H}l�$����4��	�N2~a��;�u4ɴ�|wu2h���~9���I2}x��m(��H�W����asެ�2���W ���﷮c&��l=�l?O���&����d�z�����u�s����'|���X~I�5;�	�>d��	Ԟ�k	YXN�{Ogo���u���{���J���
��OY>'XN2m?O(i����CR�O�6}�?I+*�s'Xu�s����'R킇z�ϫ�쯨]|��_����{f�f��4�wt����~I�|�VV���N> ~�N |���y��Y8�~�>�i��y����Oy��RJʇ��d�IS��a���]U�}[�X���8s�_�^���(c'�t��B����ް��m[�$�Y'u�H�z���,6�4��;CL�d?O<��u��I�����'Xsg����TEW���W랓�B�n���s�'RJ�>�d�T&�ܞ$�'�Xy;�!X|����$�'�~d��	�kt'���Me�'�SS�I���a�i����z���'c#�T��~?���~���_ǩ8��~�x��h�0�	�4{̝I�VC]�'�8���O{�l�d���2N�{�O\d����(OY4��8�=eNl��~_߹�y�<�sϹ�!�0�<���8����p��N ��	��a��é�I�9�:����<�d�&ߒsT=a��<�+'�Ǵ���m�����_�_��=M?Z���JWW�:0����*D�{�*�=}t�ՎXr�f�����aee�
��e;��,i����L�t-5ǝM�V�L�	��w3`�ˮ�;p�ES���w�ui4�Y��{�����΃)S��.M��B�{��������|��ݻ��~�$?'����Ci'̩�ՇX�L�N:�ɭ��|�:�<?}��a��a��	�K��d���:ɷԝՓ��ǿ����~�{�>���ߵ�����7�������>ed�C�d=O̟2�l&Щ����>Ӂ�N�Hh߹
���J��=�N0��:�u���u���K��/��WZ�k�_�����g�I�L��s��q�m��*M�=�%d���e���q��q�|��5�è,&��aĜe`s�
�����~�3�_�~��|��{ϫa��+O~�;�����4��>I�M�������d��|�
�6�e���C��|���
C�:���ˌ&�q4~��~d�to�J����>��5~����,�)��w6�Q�'̜|gNw$*P�w���'Y4��P>vɤ��{�	��&����T�l��쒱a2n�B�|��H|�:(������ҭ����;[1Z>V^���k��m����̜��vo0=d�&�P����NyO���&�>9���'�4��a6��>9�%a8���쒠�3�m
�Ԭ�t殜�=��}��Ϯ�ߟ~��>���z�L��&�|Κ�ƲM��~d6�߬���:�<v�ß��'�&���^��&�=�'SL�a���rC�4���,��y�n�[�����a�g��~޼����	ӗ�'��?@�N�s�5��q��~�Z�8���!�����xs�:�|����u�s�ܟ�8��w$�i�h,�;n�������{��{�7���4���a>I�޲J�$���J�l������2u�������?>�u��>7�]�i}��%N�V~�u�_~���k6?~xv���������z|ɶ)�܂�Y>Ag9BuY;���:Ü�$�XN�dY7��)8��'��_�M���i�l<=���G߇�X��+��y�5qq�%�ԃ�m�I�����}���Q��ǳa��ckWR�B�]��Zz��@�oS|�u\B�t��\��0���I[1�8^(wUwf���XM쏣��oh�c�0�Z�������nj÷Y��N�3�Lo��������{]wr��n���$�X���u���)���,�܂�>J�}��2{9�?2N0���+�$��N�`~�d�|M�X>���5i6^�^^�{�?,I��s�@�I=I����@�4��<7��	�
���Ad�?O9�Y8���{��N$���<d���$�&��I_'4��4}��G�e�k�`��oP�v�s�)&>���a���a�4����k��i��/7I<C�o�a��5=�d�T&��Oq'̨xw��O��%��~����=��6�� ����"��ڽ�d�'�a<vɤ�������u	��'�y�ܓ�:�����$����d�i�z�=�d�V��~�*����ƾ���7�W-��|?>M����=d����g�'��zԟ�>Me���d�k,�$�+?MP�N!?kx����,����d�Vp���N�ygS�$�>�wÏ����/{�����}���:q���	�s2u��Rzw̓���S?d��Lۤ�R~I�je	�~d�k,�	�?��I�i��'PY5�p�W�W�|Em�]腿ߋ�g-�Q��>Y�'�>a�;���N0yN�u����m��>x��y�u$�����̆��Y>a�+!�c'�)���:��C�]�_u�&�S���W��؃&��?2z���{��8����{���9�u�I�/2u��2q���L�z�_w��q��y3Y%I��������)�Up��>�
2~=��y��'o3��Q�|���6��6�}���J��>��������HVN���0��	�&�s |�'��{�!6Ͳ}�d+$�s,�>�_W�W�Pl�tH*���3[�w>B����,;l��&�XY&�q?��~d�u7���}d<��Y8��h{�����y�;d�L�Ny�u�Oi���toc�~$���H$�[&����:�pS�Vq�9�`����v<�?!���G�gQ�4}�qr�Re1v�Kr$
�7Md�܀2��׫5���A[}�H���>��oUԣὸo�b�R��+Om���1��m%���B�VS߻���꯾��G��ֿ}�o7��V����J�����B�|����m'm�I6�����q�ߘd��!�3�N$���:��	��6��`~>��c��7������﻽��I�~d�ۤ�O̜�Ad�C�*
�׉+'R�~��q&٩���'��VjI�~ߙ��̝a��e~���_��Nև���[�V;mS�͸�W'6�s�>d����I�~d��;���|ɮ�d�C��J��ϩ��iY?e':ɿ����q���凨���:`�]�/�7��c/��?}�'w|ì%gk���d��Ld�OP9�d���{�C�M��'Rh�%J�g׌+&�4~���}��i�\�� �}����3������N����4��<�y �I����$�X~�0����;ܚI���;�P�'�,�)
�Ğ�Y?$�O��������%���y�/%�������d����,�2|����d�!�5f�Y4é<7�@��d���$�Xy�u�W��N��
CS���N2|���_���������J�)_�0���A�G�>�g�'����]$�}dXi��8�4���Xi�����0�:��N0����?2q����OP�s��J���_��AD}�?���p3�D������C�&���sx�2h�_~�m��Y+���O�?3���u5冘q��M��ɦN��Ou�I�4��?}��X��>����v�/�S.�,�כ�z�+�$��s2u+!�;���|���� |ɶMo_~����i=k'�N&��|�&�Y�I�T�ՇXq�����8�]�T����w������'�~��uN���=����CY�:�$�!�S����w�m���}I��2̟$���%d�������!����'SFY�I�B���O�~����~��n��5��9x��>{Ql.T]C�r ��+k�އT���
��vVj�i0�U�]R��G&Xq�25��'o^o>{�Ro����|`�/T��m�ʳ*����w-���uj�g�c=J���G:P��]�B!A�q8��+Pビ��ڽ���[��G��~I�2���"'2�qb����{!Gw�DT����!��c�R,���rb�����O�cJ����cx��gY�z��y~��y��ۘ�ڿ$V���]�K�@Pj�>��`�鹼z��<r,��Iv뭩���+��	?�sǬz��7[kt�רN c�`��wM�|/	g;�c���8��'�k������r�
�kI��u�>#��Y֞�q-�u��O���n�uQb��W�[u��x��vi�')y��9J���3�h�)a�^˄�v�:&��v3Pʲ�5-wY��Jۧǆ)K�M��]L׽+�#�=�Wi����Jjμ��֋�����8��+��wWr}�F}�����>�Gև&��s�\��L�� �E�X(��0��]_�O���=�v�*�·���"�3 �<�m%HkQ�vf��.m�A��wwf�v�oj����9Hd�9͜�J_a�L.6.��+6A�*;�'e�^{0ce o'((�k�s�C�uxsƻU�s��rwu5w�����pEvʚ��;O*��S�f
�G�Q�[��*���ה�j����b��G;#���տwىS�7{�x�O��W:[���Q�k�V�bF+q�)��4�isr�Pd�b�F�R�����݋��/�mn�:��sO�)��F.�Y�m�i�����d�Ԯ�pL�E�α &�A��������pVnS�� ��f
f�g������;x�tn��J�ǅ�k���+�.��&&��%���L�R1ۺ��ķ$e_U�N���Ç[KL�����v�~�C�Ԕ�V��>�⽠�Sd�ȃ}��:/d����hZ��k���qWY�uYB饠�`���*l؋-^�+U��\�b�e�.������Գzǟe:��ʗp�QǍx���fH_�k�ܞ�9�@�j�7[V��,k�Wz5�X��ڦ��\�m��mZ5V�1��,ż��7)5���\@)����ٽ�8����:�|;���o&������ݢ���pnu��՗���Y�[��᫸���w�[ٖ�Ba��q�|Q���K�=`�]���J�R���4����Mlh�c_+2�[9X�HO*��R�`&�9(��p��+�g���5�J�EJI�2b��5���gt�n�<{M�ฮ�#E^���`}�|1�,:.��Ų��)�c�"� XGE*�tR��B���MS�2
�̶�+��׵�˝�u�m�b\E�yڊf�����c.��g��R�R��(.�/TK�l&�����R��U�Th�Rآ*�Q-*6�Z�6�#R��U���km��TV֪�B�R��-���Pڢ��)l�U+J�UkEb�h5k*�KJ��F����cKb���m��F�kTQ�m�YRUJ��i��R�R�EZ�0���*DX*U*���Q"´KE(�s%+Z���[F�Ŗ�ѵ-��km�-�E�E��J���1��)EJ��A��*	s�J��DJ�VQUKT���5.S�B����Z�5�[X��h�V֍Z5-V,�eX�m�+jV�*���j�mU,��ږ�m��EV�UJ�����-��5��A-�JYAm-��.S�Z�UV�kJ�F#[F�j�ڥ�iU��1��KhVX%eV(T�մ+QYmP��b�Tq�5�kU#*T��İѶ�%EkU(�A�1�V�[J�F�Ң�r�R�Kq��j5[#QL�"e�Q��e(��hYm��%�X�U��F�`�(5Z"V��h��q�R��l���E��p~���n|��p��癹�}t���t�t�aM��x�W8^CK2�0��2l�<4�s6q���JB��������ފ�3�s���������ʇ�8����r&�8�����:���u�a:�˼:�����@�]�s�{�N�O�&k$��0?��VO�8Ͼ8xR��/>�y�wϼ����Hx�Y=N��I�f��8��d�YP�'R�4o�%a�N%f���C��d�쓬</0�'XO=�O�k����a8�=����:�u���;������{%a�!�hq+'�:�)!�����ē�8�C���n�Ì�J�ߴ��Y8��{�HVN���d����
�+���?-���H����u�7�/�X�mX� ����]q�)�9�N�������X���M��j���,q�����5�mX�s�R�j��{�N���4�z\�wwNc7[��/��)�9;���x@9��9�����Yj[1�5��Ϧ���;^����rϔ�TT����*��-l{�n���M�����	nW��u����ܧ*���M_ER?y"���~��A�{���%=�����~�{k����܏>��/����׊νfo��#�ޏ^����9VWEG�\^�ݾ����6ܡ�APd3s}�S�/����^?���a�S;GjY��}��}� ӰGw+x��yͤ��H6�hm��8�n(=uh�{�(�n�n�d-a�X�{�|�
֩!&0����\�vh��0e�9V�^���S�_�����N�h���ꯪ���z7ށ��Vʚꦮ.��}�쿏,Q;��L~�k}h�	��������v�j~�So�?uΌ'1�{|�vk��$^EX�y2�(,w�s��s'og>X�✝e�E�r���
�����;�rت��;0��Gֱcl{k/<�n�.}�M�����
���^�Eř�q��o��{u��q�R:������=�۽<Ƹ|Ң�-::�u�����彡��*�q�[��u�~j��8���9˶X��W��M���u��l'�:T��hw��u��;��Y�ӝE��X��D�_\��lk�'���:R�d�R�c���l���>���[0r�c���W/��U�y��~�S5���¿R����/���z,������V���5�m_�\ӷ�x�C�s�M�k�f���k���>���_�7�c��b|�A۱O�y��Z >�Y��L��l��/���Jz�� y+�֮�B���9�ް^�����ص�b�}�s;g5b��qJ�X�}Z�y���j��'`[a���-�Or�x�E2l�S3�;1ћ��:��Mo+�j;�<���̎��͟�着��1YE���fZ�Ü�Z�pw�gM�fge;^]�g{�r�R$���L��J��Y��ъ��Q�A��>��������gu;O��o�}��c�C��q���]�g�+�]�)n�G�9��kT�R�κ�{S���}-=�"�Ε��9Oյ$��O �U��uC�����H��Mxs'C��qG�t`_�r"t�r����c[S.�X��ޱD8�-����JUo���0��r�Uݩ�tе�㭩1�ϣ���M�����yѽ̰���*�k~�W�ً��<��-�u���Uk����aOvk�o9����p�
?v5�OC'����Tg��Mx��מ�������_y�;;�ͰS���\��E�{�o{�����|�����~/��wT��Ү��2���\����߈n�Cq����[>����\{�d�"���ڣ늨��jV�zTү�bE���8��=�5˛��E�<'J�����y�T�[6���3��2��[�zv��@Nvs*o^�cJ�a��f��K�Ld)ھ����t�DMvI9�}[�q޲T��kb���WI+�/[�:ӺySK�c��՝@��?������!�vz%���?t樹�>Og�=~���xh֏����{��S[�u��Ζ��%Sӧ��S�[s�9ϟ�+ܫf7�����5�����;=+^����*�|��
��M�#���k�o{3λ�k��}��"�R�-��zxO����;]}��_�y/I�qp���;�Q�kۤ�RtV�<�-)���أ\��ϽTk����k��8y�S��j}�{7����nvr�s�Z�m
:�G�*�OW�Õlў��&BQnp9�n�����gs�{s�[�E՟\���4�X����C�IN�������7�`�X�%[�G}U��*���ڊ�x����l��ە��o{nU�9oΥ���̩��=��c�M[�{/Ck�j�{���}^R���e�t����S��r��qҪs�OL���gAhǲ�� U��qy9������8�����3;�.�oK��!3Y��:k4v��=n��^>�wK���ޠ�r�.I`�7��Αa��tKH#}׌o3Wѵ �^u�y������ӻ�(ܼOl��1��es����諭L�~s��r����=��:��x�;įoJ�kz�E�����3����_��x�"ry�7�������������z셩=KyJ��C*J��G���^P��|�t�Z��5=ק�ͪ��6�k[I^v�~��k��En���(�>:g�}땪����늋�3�n=ɮ=�L�؆{������ce�%�۾�VJ��	�� ��w��S�qJ��N~�3�E���])��I�F�>��֭֠�����ΝA�����s׬����<��~����:�l�ǭ�'Y��U��U���~�q����W�.�4zNj�[�m�uߥs���9S���cj�"��j�d��]p]彾�vQ��_Y�.�#u�5obϤkb��Q��ں���v����^@�#���������ާs�T��d�1e)�ST�GxAs/2M�@髠�%��������x��ͩ�yQF����r@cގ��SF6�r��󭿂�U��N�����\6?<�y�{ږ���|e��꾍,��"��c4d�S[�}/���L�rL�|{�-�s��n	��iv��cAoci��ugsI�Oz����u��W�U_=3!-I���ѿ��w�����s���-n|�\�H��Sv��f�5v��{c�!|�Uͺ���y-��KQ�6�)ʽ�$�G5r�¯y���sb��� נ�e��U��ev�-��r<�u�=��<�����c��ko(�O�1��q}�ڋ>/s���%���F�L����׶�]��]���\�5�)�lc���]���Y�'���a�����n���|����r�8���=���ӐOݞJ��^����ݒ���7�a�����R�N��ܬ�q�SǛ^��5�QA�jc��eb5fM�A���kz3�pJQ�m�߯�%e�E�qf|�c#���zw��ȭ�no^��|���T|ң�
V؎����ʫ�q3sܮ���"<�XY��q��}ǖ�����[T}q|_N����d��}�(��yX���䳺��޾��j�-�p��Q�d�J��U��/Uh��wZ�V�9�SZt�{�Z�GC��]v��!7Kj=���9vX醡����0�(�l\����p�mt��O;�P��7v��A�zJʘ��:�����f����bk��W�UU|�k����;�����/mG�g���h�8�6u����t�e�<*v\��q�r��@��ٟ9�V��/�`���CFՍ�:wn��M���Z�^�$�����F�o�p�����ْS�2+9��>���Y���ۏR{��~kҨ��q�>}�S��,x�,��&�;���u�dBf�ns���o�=颧��_d3�����ղ{�/���6 �/f�}K�:o�~�����j���vTzu����@�s�����*���a��Բ%�Q���{�tѽ����ɪ�*��X���[۬^�+��2�s~)���~���[8�Jٓ���J�����,�<]uC�9���kioa�ji���}s��oJ��3����!U"t��zc��V�vkjf:�����a^��c�}+V�fgd�wj�]�B�r�㎕I�FTc�U�^^>x�O�5�,�J�]�R}�7�3f�U
ͤ��t�h�R�n�V07ԭ��լ-Eѷ�f����"��ti>���y���X:�,z=-�IL����|3jd��/]�K�%$�n��A�6��.A����Z�k�H����}�}�Ė�~���X�Z�����%o�k[�z/m>�%��yw�w^�"�.�{�(����V���ξ���l�uM�/N>A>�g�=��mz)�����f��}I�U<�/x[_D���d��"}�8��T����\����Z���}5Ǿ�<��wj��"�_��g{=�V��I�{v?~�^b0��.tσ����_�znQC�h�<]�^
����)�?z[�� עA<&�:e_zw*~�7���~s9��*������9��þ{Н��ʫ���{�7�8K�<�sOSs�~Tu��+�r4��=��T�m�6���+��_/���|Ϝ��꧛�Ŕ��_88�m��)����$߾��-x"�b����ϑ�������|��kkg�n+�ۻ�b�w7�g�"�rMSv+X�O>F��(>p�/,��ɜ�6�Y��=��&�\}�s�ො����h��_��7�%ջl�Wf�͊W
}IM���r5�� ��t�t��n�u'�Z�]��n���Jđ�`�:�s@��GQk`Ɛ�=1�Rr��u�ү���uZ�)����������ꪘ�;��gG�G���~���K���Uɲ�u�\�=�E��6K���3i�¥O���_n�ȉ!���{J��,�<'U����J[<����Ϟ1���\?+���:�n���}N�����z@DU�np�y��]ʯ`ƶ�]�쫑_����S��r��m�ׯ��E9u�׽��"c�ъ��uZl�~tW��#��J�����G�ɠ�N32���r��ޖ�	Z�&=�}����1��%�{bw]��B�ϣTm�=~��!�����<�\�\���a�L���ɭjW�o؇+U�*��϶�kg;��O��n��y��8��������-�^6��;t���,�wo�{�7v=Y�{E�)G�A�]��T���͡��G=�鞚�p�7���;��V��`^p.^�w��:���$�9ҟ�YV�� W$�K�d`g<xC�al���	�m�q;����t��
:�qGlb�;{'A3,W�b����U���m��hWtz^�V=띁c�_f��bS��� O-aZt����rV�g���F�R�d�r��璟:�?vCw�c�}�+�?}_}_UR�W�g��.�~��6�h��'b�ݍ�z$�M&X{�;:�o�tm�m��ϲ�ҧ-�9;��F���W/�\w����*���-ŚS��͜�y�oE�V��v(�V�5��`��L���;K{G0Ot�����~F����jNx��d��NJ�vУ� ��:U�~��5rw%��{���j3�����9,�"QS� �{6o���s��%SѢꌎ�����yVE���j8�ӗ����-��_�a�>~]��v?w���UluA�����{]��V�F�~X}��wS6bž���|�]�Ms�r�W*�w.���l���ۧy�����i���u9繻��Wtt����p�U�,a��Tu���pL�j�|��֔����M������V�B�Ɯǣ*1�U��m�Rº��2��^��}�������n9���kF�Տ+�3[��6���_p1�Ǔ�:�u^�9�ٱ�Cd+�-��;o�^d�F�/I}��
�
·
��B��ۋm"��aR�`T˓B��7�kc�@���q�ް.��kM�v�k��z��z�,˩s3(i�S�OgK2���Z+��VV���X�_TpQ,���n�۹Ga����ݡM����w7[�³�2���S�YOV
�2�&�h.�XoN����[�#���wJ�o��c���{r[ƣ�e4���[j)��I,R��Z>��)L�*P��u�5�ȡ�r� Y�ʅՉѳ�H��YA���fT������^0V)�H݅�D��,�}�j`��.���D���[;#Je�B�);u� C��7Rmڼ��t|*��{�\�A���v;�_�t7}W����Ƨ�^:���V8NZWC�rmr�{#'{��*#�I��6��CohXB��1j�wwv7�,��*������I�5�HzLI=ՠ�����4[�K��"�*�\OD��G����4���͹[Sf��s���Z1e��y��3�G]�1z�^�3���B����u-�r�(u��!$�F��YE�}p�#[�>��)�V�0Σ�/wu�ؼ���qd���@�ء�c�M�|��^����	�,�7ݏ�Y��^Ol��m,x�������N�-u*Գټl5u�a�JN�'����D��Z���ŷ�hc	��{�k:7	���E)6�u��'t�e�zT�fܫ���Zl�SIf�[C�?f���x��,�cԒ�pf4
7���b�j�}O�5����Ԅ\_q�E0W[��v�kC/F,��bge�*��7P1��*I�0>���M�mo.�t��m��JY���[���z��`��O��kFn�T��F[�ʅ*��	lȭ�]���'�f�R�\qVՁܯOSߞZ��kFTS-X��<�ٲvS�9�n��c���TVj��Lz;�բh(Ͳ�r�E{+i�͸惸2L�a�MՅ�LX���u{�}�h$��c�b���G�^*�7qT�Ն���L�k�ŉ^ĳ����VK�fn�t�jKA��u2��~γ�tyt��;t��i�ݰWv��.k����/e�i����2��ή�x�$�c�7O($ے�k��"ڢ���5�oy��y��4�r��,�
�K��uމH�<�^`\���9���
� ޞ��z�͒��wtQq+˺y���i���i#S,��\�-��f�4׍#	L�WW ;�V]��3r��U�Ք��b��B�c�>�=���12���.���92�z��h����N�,��%e�`���̶�:�J��L�[�:��K�(qtI���u�VM�d,�T�v���V��.\v��q��hۼ;�@on�%��2�R఍�y���!X�G3N��jgyP"5�3��d�֗V;oP݀�0�0^3�/�.�9DW� چZ�[Ki���i[j5���+8�-L�DEaD���ʴ��R�յ�ZT���TUX6�e�ER�5��crڔUH���ԥ1��kFV0�-h�Lʪe�.`ո�b5+[J��0mrܥ��*ѵ���TKJ��mQ�f���T�m�VTX�mTk��2�
1�ƥcm�E*PU�l�Ҕ��1QJ���c)��FҢ��*U�e�֔�X���R���+J�b5�
؉Z�c���(Уl�T*�UX�E��%J���F��UkJ�(TRV��b֍�*#Z�r�J��(�AE��alU��V��V11Xe���ldU�[kj0��ZJ5�l�`Q���9j""�PE*ZX�VґU�����+Dkle�b҂�����ثT�*��XV�mb-J+�
�h��
�ʅ�ʢ$��s0�c[�cq++TX��j�Rڈ�+��۔�p�E�
"�KeD��kT��Q��-�(��B�"�H��Q�I ���Nn˪�~9����:�6���)�ka_w9�ӧ����9ĝ�J�T�wr�PlQS���d�����/�_}��UV���!�{%���^g��-�I�Dܯ/8�>�{����4]ח�9�IEqz�rTq�=]��e�d����^n0�#��$��^��	/g����q^��p�Ǵ=�?�Z�t���ʽqQq^F=�A�{^�=3��}�~����'������<��=�x6=S����S/6Q��r�hy�\�J��U9�P�5�X����S�lW�KӃ$�,�)�w���O0�~����߶W�b�hu�V69�_�<Z�;���]�xGR��^�®�9��$Η'�:��lC��骰a!��mx�μ��-W����*v�i�B`S�WI��ç���7u���ݞ����}#Ҷ�1�9�\���r����ywI��� o�r�7���ͽ޼S��y\��,���ԠwU��f75�c�n@ԩXo�,�~"^W�7q�嬙Bĭޡ��,��ǴC�u�bn΁���pp�H��vñ�h6*�t5Վ�Ӗ&R+����f���=��o��U����_N��[������Z�pg�en`gw6��MX۩�B7s�UW��S�r���|�����t��>�5EG��,�����z:���5�y������kxk�t��2<�۔�ROJ�⧀��Y�KB���ƺ����O�;��]3e;i绒݀[r"t����ǭ�k�c��o�U�mfzxƷ˵�Vܣ~�=��'��T��W�(_��JLz21�t��0�VΜm�ޝ����/n��˻R>��N����\�q��aP�z�������o�e�+�uV����bT_��]uK�C풝^�X���L�@��ۼ��{9�I�ϣ���n���|����yKkd�ה��F�Eɭ�=y�>��Qqf7�Mqﾙ�Rº����]uE/%J���A~���ݏީ�<�V�s�"䮍o�s��y�c���_7�C7,dw�v{���w�-�[�����~۝3����ҳW�{���j2�S���U��<5�q���Ζɕ�QH�v½���~e?�m�E�Ӕ�B@���nD𓶍ǚ*�2DF�Ǭ1C{�U�
�ovX��T8��&V��kmN;Ν���c�U���^[j&�+��S},���(�4�� ���2�*�E�����嗀3fv�ޜ����U�\�U��{&w�Dy6����7Ꞹ�Z���ur�!��C���5�y�.��k>sӻ�*��Y.�R��>����R�Ŏ4�f^p�9j���h���gd3�.ۚ��^���z���l��r��Rs̨�唧$�;������gOD�vt����������:}-{��f-�r.˓W�S�� ֱß�QW�qoyZ}/��gt��/g��ܯ-�|���S�j�(s������9!�;�������ڱVTy^u��`]7"�-�r���uJ�=���׮nk{��1jϥv{MY{����W���zL����
����=�Ý�9��T��B�ǭ���c���-f[K"�[�3&��rgY������߯fΡyф�=�z�9�e���P�ؼ�tR�wG|����B����O��7|�S���5h�n�y��&�v����;�C<Jڙ��t�V���!���}}�$�`j�Yd�.��-N^-��&t�k��J����:c��Rms�z�z��	N�y����5+����rV�3qN��ﾯ���E�7�v���^���*�"����L{��G6k�mu�e��(�?y׭{3|�n������Z��]풲��Eř�q�9��Ŷ~�iy�t����g�����.��~�tu�Wy�����������S�޼�;wm�ؖ�u�8�O�m���,�VJ�u�r[���>����㾮�9W9�gw9ؽ:��Ǩ[?Z�4<�o�g�C�}^���G:�y��[�)�m�z=��CK��i���q}t�}kݠ8<"�ᕙ�}���k^n�,�'<o�g�G�_�3z(��H�l��أ�mXsG,{��Ed�ɮ�����n?1���oy&�JR���;��^���׌�m$�u�\�>��Wq;�ū���8a_H��9,�H���j�r��K���1[9^���}e� >U�u�����u�W�Q(��۸�+T�ɿ"	S
Z}\թ[{��y�)n��73k��B^5�׉�O-�_H��v�W2^3/%�Lԓ/�`^[y�En�J���*�Y�I$���@HP�]Zf� �[�f��e�s�y.��3��Pu"cǵp�9?�}�U}�ÛK��s�MR%�m{>h�u�{-[۬^�;k��ڋ�h�� ���^�&c��/;:}\nS��RcwmW`j,/|�w�X��l�W�f̾O{�y9с~p[q���z#��=����M;Qwu�5{�ȼ�>")/go�ϟM
���+�d�8ӑ��3ႰB	B��jy�&�v�zA>�n3����u���'�M�U�8�.m��4�Љo��׹�<��:l�p����|V�|���j��b��!�r��D�fU6��H��zny��T""z{�#�ܱ�~��
�,�8W������`��	ũ��}7{��`�S�&����c�<��i��G׳��ZD`T��*ϑ�G�����Z�P9���aY�����N�3Ì�82�q�����+�ߏzM�;׈��|&]؊�֊tg`Ć�d��m���W�g�z*���3*j"A͸2�����FtL{o;ލN��A�h�m�Xv�������}@�>��U��]�����pW�z��V)��s� �#'Y�����ܺ�J��*��}5�c] ��wz���;�!�ާu������jQ^rc��pe=��j�W-�W�;v�v��A�i�N�
;��&��߾�ﾪ���fِc���g�w\��W*ԟ�W�3O�Y�y�F������1J�`ڞX��H罍w��x��̓�� �^�ɠ�߱�u�v����L���eW-�tq�^��;��|W��UQ���TB����2��\����hd�y�Z�F��mm{g��2KOg�G��Xbw�3�{���hP��	Vz˶9e�`O�49}���t�Ky9ݱ�^��;̮`�tt0.#>QA�X�`
���Y�bϒ��)]�6/L�,����o<[�>�]�Q�����I�r������$ x���2wb~�'Иj���0;��O+��W*���A���IR\UT���9a�ʑ�W��g�E���7���D�n�k~8l����X.�SG.P{�4z���V�J��N�ԗ��;��3���W��6�x��r���{�8�Z��4�>U.Rb�q�ǆT�s� ��`��w��fe���wMK@�[����@a�^4֋��@�e;uDl�l����	Z3IK�ppb�a����x�u��]�K�\�'7��љ�#�T��<���G���P�zki�ݘ�>v��z���o-#v��WXi���!u<�x`��.l��Ϋ��c�5�}u�@K/	:d��>�A�L�L'}WZ��k���Õ��cz��y�'.����������6��p>������VT�f����ح��CN�<	��x6���U��e-�u3c�s�7z��4���婉������&��Yu�����
��	�'�~����:��W����w]"=��iź��Qn(Kxzk��
�}h*��Cv��9�Q"�d5�7<_ 
�2_��}� 
��C`�=��Jr�l�J�����G�ď�����B��*ػ`1����viHH��S�i"<����
��mWn�U�~�3�{���nPBV�]��'h�����5��c�i�K�{@�c��=׭^��Ƿwͬ��]8pz{�x`���D*wf�_Åz���f]]tX�0g����t�Kwd~'���ި6l�\*Ny��2(�{"c2b�+� ��S��o�:��<옶A�P�e�5��9������}P�-9N\���E�W�,��\+����&�yy/�fDL���/_�l*�CNe_S�2��J�c���{k�#'����	*k���c0��k�����޷̝�=� [(���r�a���BWu^uS_c�7��:)ђ.�p�.nם��c�2���3 ͬ.�"�-ᝄ8vo=Ω�evN�9�3_J�.�e��[r���h[��!
mk�G��h���G]�s��}��}UK�p�����8 �����K��>�c!yU��82��$ӆ	.���^��Z��ឯ�[??w�.�*�~�mLJ�Wy�3	��m�1ȯe�i��I�+�g{K�����Z=�.�QcaIl ��<�Z���GƟQ��^u.U��N����H0߀��F���x����֥<�Dp�^������Pew��>9�m]�*I`��G�n������1nӼA��{K��Z��8�9����QV�
�諬X�Ŝc�#��`]�}�ْ�í���Y{|*V^�p幙^�_O5i�~�ö�uwM��[��8
BV�*���zOr /�\�g��T =,N�qe?|SO�EeԢ/����te�����emҌ�b�R�ѶzRX=P��w���K���R��t���I����9�m�d��^LgAxo���ARayLj�}$�q���ߪ�t�x���G���X�%9�E<�E(�cg~�W��O"�U	����(v
3M���/�=������]5cԍY�mV(>��e)|!�Ɲ�T�oS7|���1����ͥ�e��)�u��Z�#ҵ8%#մ�:�k^��:y4���6p0��Z��ʺ�O�V:Vrl�!�G/T���5b냦�Ai)ܓV���������-�,���]w�O φ��=Ꝅ@�{�R쾩-����C�-�<G���[�г%�xu���F�j�.�j���i��X���J���Ꞹ+W�el3��Y���+o��f{�!���l����C�\���ٷı�z�ţ(s+NS�0������}�'�5��͸�n�[���2�w�鄏�S��=ō�>�,P9�R˥p^x��%���z7�:|`��9�+j*����$���Q��7�^ᛈlS9��Q}�߫{��3�+����dr����wb���ﶮx���:L���exة������?a���Vew<�W�@BfA|�[�r�Dj��b���k�D˻�sݒM~���yxۥ�/��3��/������u�ek���9�g��cNUG�h[���}K�82�Y�Oz2���c�(�L�|�ќv��l*�{s �Y�	Bq�Zܥ^���Ϧߡ��N��2������{g�r�+�̭��x*A�[��}�&|3Jdb��!\�/�HV%w�{P���u�;;�ݷ�lf�)�-�ڬ�ҷ�Z�7W�i�x얾�:_�������Co���9o�0D^��cqop��`U�;�$�;�ݼ;Dl����Q�i%�vy�$6��لu�*4��%2��Hݾ��������ZOC휽��{b����Y�zѲ�͒�b8)�:*ʦ�ۂ�t0{K��w.) {d̏�;GK��4��H�}sZD`T��$z�)���W[�ݜ���U�D�>;q4�Ow�+�\�ס����xez[��<����!�G��wbFa�:~�;Q�xH�U�G��O����&�Q ��\\�{�u�ٙ\��G�{�45�{z.G�������Uwb�j]���3O�Y�y�G���$��*���V����G;����yO��E�V�#�|	U�b,i&��_�M�)ܮ.d(6� ��?`�A�ޝػ/hj����TB��C�-;����:�[�N�ݙ�G�+Rf+��x&�����ↈ�38b�ch]
��B��\%UY�{*��	�`��շ:���w��{��,�\�~�y����xA�.I�
��X�{��*��12�MF�䱼
��%tͫF}6�9��s)��!Iy?B�NU�Ք`�b�z�^uTB��(���GyNP��;8������� �9��t�2�z�3�̝����Cˎ]Y@��)(�*g��է�!�5x�$K��J����[ѽ	��G��0rv��*���wu�bwҕյ¶}V*roe����MګrA�Gw1�-�IP1���{Pfmh㢁�լ��:���rL��i�������P����w�\�ٶ��˻��bH9�:���a'�5ZN�Vf���$�@��ܠ�۸��]����.l�N��X�����1m̄T���+�ɬ]���J��`���핪���|�^�g��4vNx�:�6������1
u��<���4]�Q��E�xP�Ò��o��V7lRO�.�x�W�os���Rv�mӭZT�hVv$�9�:x���T�\�����L���V��������٧w�2P;I��ٕd�#��\b�,�]��+�1#��,1����0q��Rc5�'u��lXm��)��	#���B��#O"z��O�>uT�N��)�31�j=����oq���*7`w{���m�z3��=*L��v�f����5�VܰzphӸ��3/���֫�U��Y�R�j�4�嬫��V�7�|R�@�Kr�Ǐ;�+^�N����	k{�3{���	�!YA\�����E� �w��9���o�8˙uyK&��i�I�����'q�i�>��|�˺c�	aqr����]�)�׵m��J@�I�C��;ʸ��]6�m�?<�B7E.��ژ�*�xP��ȳ�YQ��x>ˡjp�49gT�x��׸��r��c�W6%){,v����U&D2�Q�WJ�2�L�"��j�]1Rv�z&5e�M�`�Q⮡L���o+��X�Ցn�R]�����}'@����nQ�޾�-��I[p��2������h++)����nkQm������ek�u���]��v�v::wP�a���r[�i�+ax�4l������A�]h��E���Dtz��J�RdB>�`8�*O#�^��v��s��\�u\5����� ĊhəG�V�	�Àw�e�{1���k!��F�y�^F5����6-�0nN�Q�[�|���'��&V<�s����;\�ys�!�k���z��p�O�n�:�U2@�{�&���T&�R�O���[�J��ܻ@�NN�1Ѭ%��;g�������B��k6����끄</ =�r�V�
�_R���p�5�����i�J&�!�Jd)���0N^���*�z��J��F�j�5����}����+��U�άu��ޞ%M&�	���us+����<����+_U�^ge���us�=Gm̧-̙��߄Ten"\��HD��P���N-X����L=/�V�ܬ,HA��"]��D[�s:gN�h�J�E���g([t�5� �6����QQL�ġJP�+��R�"�b1Ɖ�kDX�1k%E�Q���ڪ´DUU�Yidb��1DQ��J[Db��±��(��Պ�F"��cU�R��Z�D��UZ�UD�j�DQQq��R�AUT�����
��,T�� �QV+bŊ,`�Z�*$TX�m"-�mUTX��"�TV�U�V"�T��T�EjU�mX�R-�������U��UQ��*1*TDh�T���
Ƞ�2#[QEQ��B�X��V�*Z��khT���b%�cU�UEAb������b���(�H�VQQb�ETQTX��*���Um��EDc���PF
��1E-(���TTX��eeV(���X�UeJ(����UQEDEb�UU������X�,H����D�1XŊF"(���*�֌b�)+
�UU����֑QX����UETVڰb(���������c��v���*Jض*�]��N��1�Wb'����Wod&��Y�%��2iCr_p����!^u�ۤU�^�݉�+꯾��4��}�ӏ�@����E��Z���D��IpQ�'Ci��}"#D�9�d����q��{���e�g��*+�˅���X�:1�;����**�T�e�9��v���/t�t��XtG90��;�θ�K�E@���g�b���ڱ����eDTZ�X�������5� Sj��Ϥ���]{"#|Hp�^u���h�|*d�����>�[�0��:�/����G}~U�f�X��e`��*��my������!]ct��%Yuꎷz��5�^-LL������ӕ5�+}_LUvg�V�Lsm��+U9��i���O�U� /�*��p]J�x��|�.\G�~>���ƿT�T�I��w��Cm{�-}с�V�<fUޅ�*��<Qu�p ��Y��l�je/$zof�g>��0+{ͱ�FY�����'IЎ�>�|(�y�JBFT��l��0�+�j���D�F��t��iK��D��j�o�Tb��A�����g���B;R 湗�<�.�B�h�0�zj9 �r��~�7�[[Qf_;&�8;��=N>�|5é)�R��q�[�<�x�_�<X�z4e�5�m=.߲���ɻ���7-�ލPC�$�>{2�h�ۋ�J���ހ޵-��H�<�m�fpZ0%����9������M�j�>���
��⨧�:�����ɹޡS�!}�=
�ӈ=�������-h�5e�$�ݻ�ϹM>w�{R�p�U'?z�2(�)l(�%L� ѻ��'�qk�ۯNoՁzQ���}�]r��tL���Z�-f�p�r��(��*�̗��Ts����\y�wl\`0=U���h��ښ���ώ�'2e?B�h�,#�-g����Ŀ{wJ���)(���{� ���s�­U�h#!{����U��)��[߹�������[A�a�v�8=��Z��yt�pL���a��FG���{s'��ʑf�[�A�; (�����`��yj�Wyy�{~߳�E,�
�H�C���^n�s�?<̯q�_��S���Z�_yǄe	�����+־�����ٜgOu>�h8�c;7�B�����e���>�x��r���W�L��O&;�*��W��f��J�*k3���r�޽��]ޗ.��g�li+��R��¥;�N�s2��w#Pv��w�����r���un�^��o����Y�/�F>�F�`����+U?9��k��\~[�OŤ:ОY������F�y3u��b�o��6sǊ�[;��A�kwW�9d �Zse�6=�	8;�y��Y�n���AVq���g9������iz�_����X��`�
͖�0wK�����w���x9V��z2P~��^�LM���i�p��=2�׈����U�#2�DYn��vp��	�g�˭�z�ײQ�N�������M��G4�xXTU�4��]p�I�Y�ן%����V���ݏ�ω�{����"9�Z*9��uүYΞD<��
C	�O/�u(�o�.�$�z�W.�X�g��~�+p�2j"�ʐ�/{��-��=�1,&���k�J�!kj�'el�J#�ցB�p�k��<�}N�Yb�m�}'<�O\�>S+����[�vZS�fs�������#Ĵ�{�����V��Y�SU��>��Z+���ѷ`��z�'.����i��yQ����U������YWkCx?��~�!ZM�{Ut0�y�;�ӊPw�6���tjy�$�ֱ||"Ġ�^��L�9=�xt�vχ����o�~�<�WK�p@�Zd(�������0���.����+�/����!:��IK��ԃ�V���-l�y*��:r^1�Y>�a}���R��O���j��]�2޳Eq��Z�����[�^x�^x�K��b{1�[]��f�W�zn܎k�{�OՂ}���c��I��`�l��cK'5r�_RW(k�vH�9Կ�}��_.�Y˓��x��_�x�q�w_
���e�� !S0:	ʷ��h���#]�1ow�ޥW݌�����n�3N<���C�}{���U��k����T8ӟG�h[��2Voe����^���͘< ����|2�e���̂o՜��'ܫ��s�g�62;���H&�=����9�0z�n��J�X�z|~��F9��P�)���D�yr��P[���d<_U����G�y�[9���s�y�W�Z�0�/�#����
�׼n��aл��z����E3V��x|Ɋ.��͍S�Y5������H�
���:�"���r���P�-���sG�\�z�O�����]U�b*��<\U����s<��W��Q�|%��Bh=���jH�z���a�R*�S]J����U=�9��"
s� ���Y��{�1��Jf�u�Ӧ�S�&��7D.�A��w|&R�˒lf����aSϲa�9��.��7��u���qo����
�B�ȑ⨻#�;WE���=��;59[�b�
����|�*�����-����c.�[����� k�������K}���\�������N����Ϊ���&^����9�E*��TJ��.eҪ���S�]��Xr�C]�1��b�P��L�^��mM'��wT���Sb��혀��m���G�Yn��X�J'��U_}E�y���h�:������Q��D-L2���]�,1|����|V�qޕ�����ͽeȦ1�C���罹g��Ô
w�WA����?eg\X[O|�I{���(t��a�X�|�5��Z�Kù��x{�`\FR���c~G�w�i��ܦY�6�ܭ}�Ox�%Q���Ϟ��T��"B���it�ZYF5TĄ��7������g�vv�1b�T0n�8F�oP��9�'+�|vʹ��T#R�z
�wo��ԝǐ��"�	[h��U�
�|8l7>~~s�xj0g��Uk��� ���1��r��]�co�Lt����pFw}g�}>��G�K��
�K~��&�A=���+~z2n�w���!�g`{� R�\��f׍5�	�`��mK�ݤ�E�w}�vN�l��G��ʹ:�j�ap����^���z;*�6V	�*�����n��o,�b��{d�u�V��V���+a�֦&[S��8^���A[�{�jx^�~p�E�hR�
�qO'���Ip��]���2��$�6�k��Q9�5����+3�;5z�No6A��*t;m렗N˘7�p�+�rs�m>�Y�c���d�.�J��c��%E��k��\��xb�`���U���gdE����D�6����. �w����7�>��lWU���Y��ª�̃�G�z}�,A�V{Nom-��icL��ӗ*WO՛zoj����ބ�U��J ;��C`��a_xz
�H�չǣ����������Z��O��ʸ�٘ZO���\N�'q$�w�A�JBFT�u<]���k6%�ˠ�Υ��F�����e;��Όӳ֡F&2q�5<��t4��f����דi�ۯ��^�>��{�O�T�������<9�[#y#B��
��fWx��W;�{7�~~�P׫��:����{��\)T�����x�&3*b� ՞����O����3[�� ALo/�]Hs���s���8mx�O��Z\1������T�$��{�U<E��,�v�u������s�9L��*���S������9���/*�6���ʸ�,�А�墓��k����n1�	[��.fVMt�ʚ��(L�l�7a�n{�7}V\�+h),��x�<��$�����n�&]��n0��'hT�x�j���u�$�S�r��D�����;J��P#Z*��w�%XvËc*nNeV��1�5��SbXT�|����PN
al}�mY���P���;:U�D����a��V.�;�.����Lu3���.��=��Y_ʪ39�1v���G��Ѣ��:X�����`Q��^�΂#�[���T0f�]���T����x�b�9��Dr����P#�C�L/I������*|��hHm�HmH<��8�u���O
�I�^����uc�>��W��������ߢ�'��N��FG0�Ώ2�{����_��N��*]����>JPꥷ¥e�[���S�>�#'Y"5��I���q����b�+6Z�6<�.Z
�h�!OW ʽ�'
������'���*��NSO��g����|P�l�>Fe����t.��H��f��M<�t����};^�gD�/���ބ�&3��5;��=)��l�~������׭8��]w�-���U˩��>���Ȉ�h������U�9�ȇ�!�G��	ջɡ�:]y;&�Y�����l$S�rLd��b{�a*�甆T�����J�WOa3�Vf��Q��-�]������"�* �N�6H{=O�3|Fv�w��w�=ޞQu<�~=�Z�y�wck\�,]c���N���w�)���3�7��/x��h]8�*��[����.�>3a&X��;�����g��*��\6���~�Û���2rݫ3��j�(�lv�Hi�;�y���2���e�J��j�Mu�x��+��^q<��Y��[��(�оva*��U�b��p�j�V����<����R��O�{���l�F��)sTi��h_;!���]��^��V��vomn���ޗ���>�l����Rc�`��R�]E��I��/�,��R���e��Ź��-����0�3�j��DL����� *r��.��.�@�xW�VDG�WK������W5�Ǟ�R��i{5d>���VwED��y!��
��_�ڍ��^P��c~���u��[���� �~�C-4pK2�/�zg��n�gtU��k���9��C��9��$��=~ܧ&9���G���yh�
��j�J+��ʸ�:�����U9nC����J�w��mM��r��by�$�H������S/}e�x+��[Mr��W�_��Ȃ��u�7Ǻ��Z6$+�^�5���/%���W�4�*�b�}IHV��0��6{��׶�#��zBC� zc'>Z��V�`��5OMg�5�����7d1+�'�F#Y��9���R�.�s�89 �3�,��e�����6=s)���BEK�T1��(
�:�g�����C.��m-�`��pȗns��{M�N{�v�T��k�-wu�K{�\��h.�\��R��vI32dj�z8�=C@�]5��?�W�k��&��?ˮ�G�!Pϫ�[�ס����QqW��[��Sېw��w��0J�g�\]����/���,_��v"��+�u˭�J��aϦ� �\\S�*~��{���6yp��<c�~��u!�:=�)%�Ѥ+_��p2�ס�}S��<�L.ʎ�^��XWz�ߣ����:T�-xv4�]���s�+���S���%�QJ�A˖/��\�~�R�=Ы*-�B�ѻ,
�$hpd�ņ���"���2��<p{�ey'�����h�~Sǵ��d<�.�~�D�����W.T(Q����-g� �k���?{X����W�)R��;����p�����<=�0.#>��1 �J.k�koi�w��Mq�����eY��X�N*��.C���ϛ�D/�K�i��I��hue �L�w}�A:ax��o���nDS�C�ȱx��=v!N��Q&C�1ЍsF���ct�*���؅�O��ip�L=�
c��~~��X��z�Oh �O,[�O7�����({)��˲�{7����o�h��0/8W�`{�ՈZ�w����FV�X�|�F�ר���Ey��|5v���NVv�*���B;����83L��cۮCD�v̌�V���rS�Pz.���#�C�����S{�����N~T����z��R��3�v;:u]��~��3�i�Ɲ�&8/���<.���W��7�{�v�s�s̈`�k\���o��.v=�1!�^4ք'��ƺ��Ծ�Gő�֪*���^�^�5Gp��������}�m��qiym6�;�����b�딭�7k*o=[���������mV�X���]IJ+a��婉�mL>��zr��o���n�vo������k��ޗ�'f���=��Lt�����%Ud����t�w�f�k�
�3 -�痪�����K�&��9^\>�F�V�g�%��-���/ w���Ƕa{��4��{ϻ�>�No�f���==�)V���U]��d�;U�����J$4�$���ӷў�)�n��ǩ���ҟ�z�}R�x�8������*5H0�Ig�N�{���r*�+2N��xJ����z��{�ȉ=���꧹�z���";F��V�}풟)�x�I2�~��J���U��÷sǥ�^�U�s��z���9쉌Ɉ'�^勇���~qz9�t���E.Q։�I΍	t$���XꙂ���CVj����w������Ǣ� �f���f��7+�f�{��}���Gԫ�6NҐ}��"�Z��r2u��R�w�pWBtB��R�j�I$q��R̭X�wmɊ�8/����/�DU}�>t�����!�w��m�t﷯kjc��W�#��c�C8csǋ�op��̱�H&�u�i�ʚ�uu���C[����E>�0^۰�G0�kp������#pgc;/��Ǌֺ'M�9�V�̽Iu�P���fIkC����=�mX#�/ �����jv��.��v?צXݙD뫮���i%��`�}cn��1��u��u��L�K�Ӻ)<�������As��
��4Lkk3���ҬP`�s���Մ�M�2	)��2l����ֹ	�q�į�;����uM��fm�$F�"mRZ;�4�\�Ģ<˳��:M5˓vɾ+�^�p��Ui@�9�J�l�2�W�v)ڂ
p:in�S��rN�>w����9�o���A��eq��7m$��I�J_=��������{�P�m�U�L��,@��%��J�+ �֭�l>�i�X�m�Ƒ.�͆�KY��QGc��<�9N��S�Rf��m�8�Wgi� M�3*�R��z�"�F��5�S�Ǻ���*z��|������Q��K2�.Yàށ������@�+�{�fˤ�St=+Z+�yF�R�` Wd
_v�j'hj�Y�{�<��T%X,�4&��W���r������bE�cFwa������;�95�GvT:��o�M�:59e�X���k���`b"�p�uߊ�ө��܅g��L*�V�t%h���(	]5�Yo,��em�(��f�X�Sd�]Y��S��Oۺ]�r�w&�9���hY�Ke��b�k��8�=�&]!p�L�Z�8]���KZl�
Ty�D��/]Hv��x߱e��k�K�̆~��s�9�{p�}�p�sC9��i`��������]�6���tt��l��{9	e��"�\	�l9'�RF$��tOv�g-stl�\��2�1T�Cv��)��w;��������1��.��v�)�T�%֙��p�K��4�=�S,o(�E.���J�7�FYX`�7[���wM�a+Up%oa�63E�gu61��r���;�u�Y�d۫u}��m���fሎW�w-�;�8���Fu�O�-�}�)_J����M&��݂ť���]W]v+n+�C��&���*uz�$5QW}з�Gl��L=�
֣ Z�.iQ�}ʾ�u��>�����dv����][��.�F8�\�=���|<v*�s�܎�2{ԝa�q"6���_���H**�#��3��.�X댖�Wd%�l4x��z�L,+ Q�s	�f	������c���*0V�X �"�l����E���E����TX��*�UQUD`�e�*++A"�UDUF+�*�m��(�,��B�Ŋ�����"�TDUF�Z�#���T�(���J1U`"�F1AQb�EF"��X�*0E"�,X�[jT`����� �"��UVVQ��
�EQX�[,b��b#R�UH��,Z�bEV1X,UH���DVTX��"ȣR1cF1�`�b���HX��UU���"EU���TAQDb֊��VEX�*�Ĉ���(��X�"1Q*QEF2(�URڃPQEX�X�YPQkD��*�U��,,EQ*�X�������",Q`�X��Z��Z�b�"(�����b(��PQ#J(�X�X���*,PDADDUw�sk�7�%蕣0�^q�[DW��f��tW-���V�w���/䞾��u��L�W���hHƮ���WF_����yN��k��]�@A��ӅVp�h��=T����}U�Ӕ��=�ۅWu宅�7��X�Ւ��"o��Z\+Qb�b�x:��00�uL�B������j������7��2,��ͪ�s�pDI9��~9W�O�k,_��یi����(��"�olg��M=,l���������}��l������K�E�U��O-F��F9n�+��ޘ�z�xx4gsDU�`U# *r����O-T�Z�2����&����:fJ�KW�kƧ���ӈ�w��Z�^q�~&;"�yyT�]�3��ťO�����ϸ�S��?fK\ii�I�\<���-U�r��<�q2s�O&;����]a�\]��9�V��0�^�H��"J�ȗ%�/S�OP�x�W�R�]�3�M/?w���eo'N�"V��]�^ �����m�aU�-tJǡ�.X��2޽ ��,��k؟�>���<6\Ք�˞.�@�z}S�2��^#��h�������/=��V�����}��zD��L�����iNPs��k.F���+5�Р�{��YjĬ`et��b�5���J�w�.�����P�Ӆ���ZO^h�ܵ��j=���N�\SU\��l]΀�/VYwҞ>y�N���;��孀]��� 6.������=�=��s�j�G��'*j��;*x;�n�[*�ƚ,N��4��aP���^e���+u��a��D�+!���pM��"O]h�������U�9�O"}!�q�/�ޛ�mfy��\3hB`���]
���i��7ŉ��v�甆T����E�[�r� =���7ʹ׈�+��/��!�B�rv�7ǘUُ�0�{���)�e�٨��)���uw7p�F��Eb��TßLj�d�}WlFr��.M}2��p���h�H{�̀�87���{���#��a�1K�b�Oi�49�>�p5�RPr��] ɒ��zE�-|��u���E��&;��P�.
�F���$��ĖxE��1p���X�/wҹ�XR^q�8o+�ֈ�U/!���[�2���]��S�.������
o��R��/4�<�j2ϸ��/Z�t襺���$62�A�r��;#e�	�M�P>�����l1�"�U�m��>̭����OC����^'�\�Ey̔,|�l�����r����_��w��m�kE�Mz�4��'_`���pv5����>N���m�^���ˎTuc}T3���5�ON�<f���\w��Y��[�����V��e�X*�[Q:����@��B��j�P����fgVS:��G�i��]�������O�U\�~Ǫ.���U;ѫo�����o�nh5H�^�������U����Ƨ��Sv���nd��z���}����� U~c�&?	�Z�k��[O��ǥ\|�_�~}�/��P�_-��w�Y�^HW��Fg����d��ܯNV�#|`�[}t�����q�N���Ӟ�=��t+�y�~�U��=�S�Y5���z����#lZ���oޘg��{��g�C�^*��P��5(eWh�ʽEmN0{���NOK������~�N�&1��e�Ǜ���58�2�o�n�R��W\���J{fr��S��\�)Y���y�pP�
�05�kc�.�n�4R5w�ɢ��������H��rM��d3ǧY���m��7�\�M�����2����J����Ƒ�#�&���tiS�؀A��7�lGd���k�����m?(ϰ�����`TQ#B��v����4X��-���2f ��O�n�>�s��°I�y�|z�xN�/,����5{B�}ʅ
9�x�3UAD?�z�Dw(��%�j�,�)u������kQU�i�A�xcxp�Yd�w*{n�W��ATԖ.��Ǐdl�Jn#�i���s8�p��Uz���Wɍ�q;�VҒ�fw|�n���&Y�Y�B�W�S���\C�w2w"�����} O��W��l�J��=هM;��	�?4x�7k�/�na��`\F}J(6z087�2֍�
9[��� 
�#��X����w�V��T��WJ�'��9V�U�i?e]���jY'w��pAJ�$4vG��U�6+�E�����Z�Wt�$�`���K�a��y����O+��ݓ�}�'K�eT��ѿ	�Z6}5P*��a����uV�*��oG�ʓק�N-��K�T�a�::TU6��_9xΓ:{�Ġ�~���˴�h좎m���C<�tnU4���{3�����dՌ���s *�� R��OA�G{�;9Tܳ���>ӆ��4��|!��h/=nϫҸ�5�ټ�J��8l`����U�z����*杽Z�d��Y�{v?0�9Wz�e[U�b�*�u$�eq��V-LB�#��=��kPV��)p<�PK�d��3����7E���LJ�kP4�:�Yfk�
��̂�V�^���jn�N7��i���t�ʂ�*�X;IG�,�Ih�����m����8.��~�<��5����5�̺-��,&o�y4h	��<)��;+}6�Yg9����el��ޥõ���b��RM�h"c�1.�/3j�gr�w�{�Й��:H:�c$���+T�V ����0�;��T��t�w��T�����?�W��zJ�����ZB�N����)V��CS.�qI�}}h<�|(�~��l��16�7�z�N��w��LR�B=\�_�z�����P����4(��
�3��[f�4���ބ�Y�S��2R���(��K�{ӑUOnt8==�<3�`h��#��hWxk��<$�Of9X�6+�!/Og�WZ�.E�n�>�=ҥ��JN~�OE<e�>�J,/��5ܽ�\��I�n��Ke�Jc�)���!���0��0yWo�>_{4�\��+X�ђ���'�V�	��ou�}�&p��*�US�u],�U��P�6�MV�9�t0᭘�1���+E��v�z��7iٞ����*�b�D��,��r�U��z��5wX�fϲҙ�{5�V<X�$�B���9`VА�>��S��"K
�!�얞�)s����9}vV�T�y|=�Gaϻ� �s !��� �܈��:���ٳ]�諏��~�G�����ҋ7ROh�*׈����'�xF	��9"��J��if��
������ʻ�� �XzwyI��h��^T'K���զT���6W]�Ɛ��Un{{#N�����v)�K������y�y[�!��gHN6��3����r�vïN�e}����n��G\�0p�v���;1󓡆������3Y�K!��ne1��au媽S2����L6���ʳ��#������u�W:�ma�����a/���׫�6�-�5��<[1|{>3��1�G�T�R	|�>�����
�^Rnq��W�.X��U�/x���յ��1�'��j�}��_xh}W/�ʷS�qM>����Ol��U^#�p�d�Y������j��G�kI7y�Z~�����ד�Y����r��);*z��6��*�ƚ,N�\+C������z��z�Z-`2�|j�#����+�B�qK^��'Q��K^Wi�q_k�#�'��H��>]Q�sq�OF�F_P�~�Es7.������_��"�~S���8��#����߼�Wy�f��C!`[�x��< Th����k�ǧ�����htw��˝/e�}r}'�G�{�];�P�Դ�!\k���"e�e���V��jy�䝛�CHh��Sޑw�}�ܱh���O\�H\1�WMS�hs$2}V�����\��~gk�S����F:�&���ktܶM5<�cx�M��p������Ӣ�;��"Z\X��suc-.+��EB�Z��{�c�5-ޥ<�U��.��aꙁ���VYN� ��q�}*N&�f�V���5��yg\VF�o����G	]}�}I�������@l�\Lg�S0k9(�I���.�a\WO(�;���jt$�����o�I����owM��RP5^��Pg��h��/l���[�2]A��ب*?�`B����C�'l~ �WV47���n��m"��)2]'y��}
��_�su�Y~�o:'�۽�̇�,!c@f�����f���ߦzn�gtU��J��2�|���e;��}z���-�<6�5A���e��Fz�G[��>�:3Y�Z҇�f3=r��n
�ں���c&i�t���8L~#]��m:\�z\|�~;G�坘���Jc�������Z##ԹxL�!^��Q�Y��>;Y/x�����5E*��Ɓ���N}��ҋ3��|���=��qjbg��`��T���s�����i���V㱭�̧�ow�0����Ң�t(֡�����V�� r�}���~VO�7ޞ��Ʒ��]9r���/�	y/ƫ1��������/�؄��a�>��@�����Aoѥ6_]�R�^�L-��W�嚫"�3�RO]*�:t�Fi�2}�d�C�7[C�6�:�y��;�I���fAE-�w��h��f���J�.V�R�[�ػ!�Yg��V�4�f�,�c{z�΢u�j0P����b���_p�E(^վ�O�[ODN8��s~�*�ݕ��a�^aQ�4P�w3��o�6��[#�vB�ұ�r�\�.����:uP��̭���[0*�i(�#�P<9WE��2���-���gpl�C԰���b�:����k������?(ϰ�h� T~�y ���������sR�2I8;�AIzKU�PV��~OǷ�1�C�`�~�I�]O>��
��B�I@>�4}~��^r�[=Ƕ;�t�V_h���`S�G�cqV�K����� �"R��]�m��sR��͎�|���g�_Y��ϒ��U{E�q�9�Ss(�
��T)>.\ͣ�~��|���I���aT�ƍ]�2���t��C���UQۃ���<d���M�н��q7�nf�;�B�י(c��ϤDh���Fϴ�L]�/	%�;w�6�/Wu)��F)��y�Į�uʺ;U:�¯�M��s�L��^~��h��el���������!���O����Ռ�\@��@*�1={��a�^g��v���!MD��j��Xc�{º���l󗩍a��X����DN{/CΚ���b����d�B�c�vxQëFԶ�S턍�+̙�=&�n���<��cu��kJ��R��m]�D�{�V�4��M�39K}H�[]�)S�9�sg�nHa��F�sA��m;߈�-����;��|�xL.<2��<#+�ʷOC᫹�e�n��q��&�t�ߪ��4q=
ڸ�N]1^]I:\ka���12ژ|</O*�ʇ-�K���ݻ��~HS����~�V�]�3*�'%�:޲�8��|����n�R�.fݸ���k�O�ji�б�OeAXPLO�g�XT���O��� =d����֟L��؉�g�,���jg������Z�C��˺n��v��|,K峃�x�FdY��<��9,w=�I�FS�u<r���vR�����\�t�T�خ 2v��K���4�旽r��"���>�f��q2��i��gNDE=�����<��Q���g���|�W�eA`�$9�o�i��Ы�\���d<h�=�\��SO��^Ե\)I���梨�9j�ܛq޿)����d�t[ȀP��Ү�s��G8��V�mx��k�E�Z�{��^{#ӵ�eWK�=����W��H�zF �l���5�ʡ���X[QK�=�����-�����ƪp{�9j��A���;l\�_L��X����l�ex���`��ڟ>�[JG-cg91���Ǩ���bE��Me���2nl�ew[ݏ��}�pv����:��ۻ:֎p�i�z_�r��p
�S�tVV-�.��ϭNO�W9#�l�Y2�̥Z3�,#��"��*�U��e�zU\�j���<$~x�C�b�5���>�4!��,�N9���>r����K>*�%O>�"K���I,�IrO;�չ��x�ֈ��[�a���� ��d�[ (�'��z���e�EJ��sG�^�~>(�q�����[I=��:=;<��
�ϝ��X�W�a�tu�Qogwr�]yiږj+[P���?fz׊��[I2k�}�!K�{K��U�ǉM5Һ�Yī���ǭ�ԉ��cv7X4:Ӄ�ݥ��I^ᄺ�^zܡ�o�J86Z&^�c}9�=����1��2i)��O�}ry츾
�Z��Jǡ<p��7����ɋ�)?Lݏ�b�������qe?�^���~5�!]K�ᵁh��W{���z�gV���W��f��P���$=B]MPR�.vT�w&�{e_��E�J�: �繹}�;uq�^���n���Y��8!��^��N�"�U��hw��z��ʯ�4�yy:�f�7F��s�Fι�.��F��z�,��r�p�k���:ȱ)�{�9��@����`�]Ʈ��B1��_n����9Wq���t�)�%��Ω����[m#w�n��|�[���[k�d�X���s��[wB����7KrSgko��ˎ.Ӓ�Tb>�-��)Qr��h	[˶f*�=����a�����m>��|�oj/�rs��f�5��fѺ�)�W/2�v�]|�(kEn���lX�V��@�r�XQo	d�v�/A,SY��^����'M��l���fU����S����-4��hʟ���0�>ي��'n�+H�E���^���f����T<��b�_�r���dЄX�Kf��(M�[\�<$X��}��&�k���Z��b���:fҕ��9_U��.{��$mof���9:q���ڤ���w3wLt�KS�C4�oEٱ�����ZQ�F���q[�!�`�e\�o.��!<��"�����ԹM�p�5�;���ۖ_��WFd�ː��ظ�ԛ���r��eo5�3zS�g[F�毴���L�t�ч3L�.�Ij�Cv �jŎ�}�) ����`Mt:��-pݹwoM�g78�JM�s�ʙf%�w1K�v�ͦ�'*�*9�a��X|���m�;�/�Xq�D�iu��ʲF�i�[~=̿^�$��Q���^н9K^|�2�o�ƫg
N~m[���`P�Ш
�m�<`����غ=�Gu;��c�-�M%&�vM��ԼA��J�j²��j�����k�Do���]�2<jk
�3o=�H�W���Ϋ�}Y���$v"d��;��:o�+��뱮��5��q9�dP}y�.�V�Ԟ�i����S�z�vT����k���ͣ�� <tr���ӱ[��9�yh�rV�t���I�8хst�B�{fi=<ݨ���866�η���w%��NL�*]pHh7o6��D.����_)ܮ� ���Y��[�0)�b�56���$����bg]҄j}D:s�;��a��E��vۅr��1u��.Z-�͇�ls�Q�������Wz�%)o
 �ѧ�6�/y�E�EC/�֣Ok��`��v��]#�F,��i����_>��!1g*��d�}j�X[�\�N����O;@�W|0ȟs9�f�`xI�_Aւ�jT��]Y��`���]oVf�m��ی�K��u�c(�L�ɖZ9�Dw� �r�X�A51��"]�]ȝM�t�k��%��9)�76�p�F�(ut1�1	�n��vu���\ݥ[��8�cYV6�m=�֖����P��e�β*r@:��Q�Ȝ��Z��ҷl�e�]zbس*8$����IӋb�8'r�ڑE��j�F�l#R�$�e���4�lXw7�ڋ�]���ks�Тo��&L���#m,��|�ҙ�{z�ܓ�w��6v�����	3�]��&� }_
 | �V�F,��"�Eb�E�((�UEQc
1UUb���1���(���c�TQQ`�(�UEb� ��"��EV"(1F1b,E��D`�c�b,X�$UPE�AQQQ��-�UDDUb�ŭTc*#FD�"� �0TU��Ab"�V*,T�Qd*(��#dX�"��
X�ňȢ��1����"��"����R+Xը�V1���EU%J0UH��X"�*-E*�#f9�AQU�*�Q`��(��)��0VV�H�c�(�)V1R
��E1��F""���A���TX*��*���������PV#�QAU�5QUA�\B��DTb�UEETTb*��

�Ŋ
)1(�XȌX�`�(�)�Q`�Q�(�EDEER*�*�Sϻ{�5����j���=�|��䐁�ڝ�:�Vˤ)�s����Eu�[�C�K�}�iD�x�
�ZO~�Y�۝��wN|F����΅� �]d��R�Wgܞ2r�o�};�Os�C�F!k�׹�b_��ִ��p<��!��!`[�x� �5���Y��Lz|�b��[�ѷ��~�1���Nez��=���pV+��x-��5f��	WlFr���f´﫽��Ĕ�u�|ߍmλc�}Mb�]%�3F��\ÕS*���4/���V��n��T' ^^�T{ٵ:e�R���qBv �.���)1������J�����$�M�_�w��z<g�D�����|L�����z�M1��c��]�!A��Ci�3�*�A㴮���
֭���s�EX���U�o�Y|ubR^�s��V���蝾��C��ya$&$o��zv��Yh�9��a����=kYBh�t��^�!d��'�˫���,+���go��t���:�p1�4E�v�4APs�!�B�/���;���Ώ�2�	��}ۓ�bW�Е��V�WE��ǀ5�� ��;�^��t��[����3;�o'X��ޙ%Z+ K#/�'B *�ޟ�!��m�5�5�<1'J����a
����'o�YOכzk��x�m����/M��N��,Sn�2;����v^|�.�]oJ��z����d�3:<��1%�).��6�{Gj4ѓT�g�i�����Y�@�S#��d{���d�
�y����G��:>���A���Z��B&}�s!�8w����xV���*��Д0{K�������:��G�0����[�׻�M�Z���'�Zg*ΣK��\UԡF����9��b+jq��\U��Y�8�B�Ga��{×o�ɟ\_a�5F����$��6\Ln�pc�8㞋��Q�z3+M�xg�N��6�5�k��U{3�|8Z�pN�t�xĖ�d��UrM����Ů��/T7;=�<U�^NY�O>ɇ� �se]1][-Tk�4��b���s]��81p�v��Gn�'��Tݯ!P�,��<���?(ϰ��i��e�QTH���:����r~����L����%�߾ʶ��KT����'�����g^^&YG���j�6�s�V0"��rZ�*|�^��^Uձʲ�0*~h�n*��y�9������v��s%�={u��ѓq  �~�g�UV\<��*|W�\���M̢$*a�<�'�-��=�~.Sw�pW�wT^��w;��c:�U���
Er�KǴ��(mh��<�|��ڼ�/ϖ}�P3+n5�؜��]�'��wܮ���ʾ�lg:���	��/C���"�#��nE˘��ջ��5�k��]?�7�B���Il�I\ъ;��79��ZYE�5LHA�O�Ȱ�ve���1�����hC�@BS~��i�{����$͗�c���uT��
�%�p� R�>�QAJi�yf$���-��s�s������*�\�E}"�AU9xΓ���[�@�3~��j*D�n-b���J�I�
�yw�U��!�	ծ`}������ݎ���{ޥ�{���ɭ��~�� �Ձ@Mdږo8K���\�~��o�w�ڲ��E����b�-�Mn!{�Z7�=���s��Y�f��ۆ�'j�+1V��t3�5��ϖ�&[S��EX����N�<�=����3~3�m�+.��W�,0&8�Gؗ��R��t�.��a�e�t�5c����>���-�D��� ��ʂ�ش;	G�,�Ih�~`N]�[�z3}���y 1�;��l��S�����8ʯ�^�� a9�t�1���wuL��l�����oB�FD�9)	8]O�dG��K�]o^us�t�T�خ���bml���n�:��==G����[j�a��Q �]{he����"�m�����z����oWk�z�3�LӖ�ʚ0F�5���ܭ�{y�����P�m_۽�Q_s����ʝ�(�hKT�vU��]�N�wW��:�Sij�\��0�7w�y�T��pvrN�u.�����=0VIȈ��:��y���ђ��~�����V;�RGn�jF�]+hY=ʺ���Ȱ���ꗪp�h�����E>/=x��zNm�,9>Ơ̘��L�����F��+8]5G8��V�~y!�[%r���ؽo�9�ӕ���VL�L��LGBY>�b������^�I��� f�+f>��E��̵8.��Ӗڒ�i�e\�V��g��E Q�5�����#,����i�R����8�ʮ�(8`yP��e9`V�_Ig�Sĩ�yX�u�!�V���r���Z���U�G�d�=ITH�e���#��}�`# '*�Gd{)I��Ƚ�o�oN����-W�V4;=�Y��VV��x��|�}�J/8���;�YR��Kٽ���d���EZ�Z6�۪�ȗ��>�2k�k�GV<��WJs���/��C�����t4MmBr�<��ڊ�pU�����]%xdK�痃��=CAq�iE�Z�Nn�d��v�[�%�'H��k��A�jB�rwb�}[�#�C7J��s�L�v�f���`K�u�5�]�=�YM�}A�d�w�	4�$�����euN����W՘��d"r��C�*�X��.�;���n�os��J��Yʷ3+�����~�>��F���XUf�])+�|������aU�{�+�S������ e�2�Ŕ�SO���/O�{fWZ��t+E.9I5�
�1��7��,���+�B�[�����'>���E�ʞ��M��ʿqʠ�<�-�Z����y�v�o>����u�Vn��R�Cd����o�az�D\�l�]�����/���~�˥�eS~DL�$C𾠉�MQ"���Wgo �C���E��T2Rh>Y9���-����o��9�OaK9g�@��|h�8�~�S���\o1ײYS��������0H���S�b��h�jZ�RB�rpTL�̿�`k�3�4�	G�[y�<:9�7)��O<�z��h�%�}=s!�\Õ2����к�d2d��4�����������z��I@�޺���v �.,P?T)1�	ghu)pT�5&)u�3��	��w=�R��X�f�*��c+��e��DHP��o�(��k��+3x�pH8i�I�xp`�gp�Z�>�sr��U
T�����m�.������!��"�-�z��FT+&p$���e^�7���C:��H"0*R����A����JGv��
%�,P�ԥ̳'�p��
�ǹ��r����w[o�ZB�:��u���G��߼i��rw_
��yD��� �#��n����u�::���U�'Dj����Fk��X:��νIx�ݐ�q�Ƚ��z�,v�s^��ݵ����Q^s%�8a�2,ed��:�!�J+��ʯe���)%B��]iN�k��[��~EЕ�U�R�g��NM�C��M:�	�Z�k���<�Ḗ�Y+����k�d�P�[���q��HG����d�
�W��ʯG1�P�O}=����֥%z=�����fY�I|X��'x����	ũ��nfz5OMeMj>�{���y9�M[�s�k~v���7��vΣJ����ЭB\����9z�ڜ`���}&r9Sf�8���ښ^����*</�˽Fe��t:�E3��mW<������V1�Q��Ց=�w��y,��l�J��U�zN;����:C�������MX�S��[�b��L�ٵ���c�ՠ��^��|L/�}���f�T�*��v4�]��U�h������̽�5^*h�Y��J��r�6N6���z쁷��EC_nP��^��@��SZ)��rudLu����s�x�;���0_7�mV�BŶ4b�L���z�6u+k^��&�����.8:X܂�Y��i�h��Z�îuv֬�J�Pw��w��˹+'Vw:f�#H<���S�'6����m��9���el�*K�B���n�}Sy�����FZ'hC/�4xM�-��b�eQ��;��2�f�oڞ}
�87���k\�wȫ��jgd{��TI���>����~h��ל)xl�na�:U���#-�y�6��>�DD֍j�cB Q�g�!��~J�^�r{c�eSs(��!�\���o�v��b��9V�V|`�ULHA��,���vدi.�Zh^��>U��g&��ޏ/F�)ɔIU%�FD�r�=RYS����}�
�P��U}<�MM>OA}�ض\����;Z%��� >�J��ʕ{��0=Xx�ۑ;��w��Uz��[l]�ׯ�pf��y�T��φ}72=�������S������[���ך��{�'��~����#�\7
eW�d+zД�/60myǄw�;��A8�^�;��F���fs�˕xn�2��.��*b��RN�W�egԵ1��2���U��{r�z���~�2�D�[�<�\(�����	�c���ij���W�4��&��vl�6a=�XDt�K�� X�7d����jVq'<�'��b�}`T-TӀ���z�f���:v\�y����vm��v=��}��+;�&�Hc���(6f������n���mn�A��f����^��t�I��T�%�[���}�w��,ƾ�U�� �o��g_�W�dL87	G����Ė�z��)Td`�W�v��%�~�y.�Z�s�va�q��OOoJU�����t8�:N»,I��΢{S|���^��h�f�R��)	S���Ϧ�?N�,�u�pyњz�x*{\�q�w͡�}�9��_��$�=	,f�Ųl��\�ӕʒ�M�'���W�⬨5�|�������z+�=͆1�]���,�fe��5X�1���K���Z��iL��>�
��V�ӷ�E����x羬��ʘ��UT�`_; ��p|��]8s���85Yw��r��ݭ�[Mʧk4�z��Zq˘{=� ��2���d/���-.��\37륕��'�i{����]����}�s>:p�TY2��J�c�ڒ�i�e\OBC������I��d��^־齺*�]��C����83�"J���Ф�g�X�Ig�<J��T�wO��u���{+o�����jX�m:�+���WO�mV �Y�¹���Ӵ���[6��me$�2І�����to5s�[Yn��S�_�'w�j�t�sm���,�,�!���h�EL�h\��F_<�t���Rp�����Ō��*��=�DÕ�k�E��
��`�	�kղej��~�N{�y�si��!\jV48��i2�����N+g�|,���J�r�`��KcS�^n�VK#�C�&w2)[�^�QZ�����?fu���
I��\�y	t����z�����:�b|םg\%Z��Oo W������\�~�H��<�^).K�^��2ђ��a�~s<�[�i�	T��Yz��ʷ3+ާp2_���7K�X3~6*³e��%cг�<����ND�Sy�~M@^���z�@���qe:r狆�/L�E[�x��8�������<��L��e�"�V[�vp��E�NT�/���=T�<�OՊ��=x|,�(ꇗ�.A[�MѤ,Dr�Уdu$�u�t-Ql`���Q}<�D�B����0��`��o��f��^��t�!�D�a�Q<)�(�W��Q�N�_�<5�/E���Nl"������H����)������U�򫧰�2!`_�Y�< Th���\�y�=�,�F�X�Pm#�Wkfvķݮc'���%[w�}e;�z�8}��m�j��fx�� G�/��u�u�a3|P�S�u��Z���^�s-�Ur�S����e�h��M�z��ԮFx����4��N��Z�WKʗ�l)���c�>�ޅ�]����L0�����:��K��ּ*9OҶ�.�hоva*�Ϫe!I^��ߺ�x���V�R�����]��W%�zy5c>�)��z�B��ʺk��خ�Y;��}�{8͎���w�����^�]n.'a�����W�Rc�F�P�`�~���ʫ�i�5k;��F���j}�/�U�<'�(9z�M1�G+��h���@�L��6������.��A�����DIu�W]��S�.���V_Wrh�>
��td�'A���N�KD�<���3��6'%NU�'*4F�(!�֑s�C֚<%��p]ߥ��JW��k��NrN[��z{���ҕ8��cDxn�)
A��a�ύ��/x{eٜ�t�c�ݏ�+f�@����=�r��\K�~������{�d<�T(�|ҋV����y�c߆m�pt�&ҡ���!�r�]���Q�Y��>;���>��|;�O^��.���m�:\���p�.�����%!U����ip����\Hfƫ�����2箱*�t����VS��Κ��ogYe*\�cYf�����b#s�l�_0{{"�֤�W�R�56��3[��� ����tp��꾨�_�[���;������meM��7�Q����oj�����#ɕ��P9&3��Kr�{��l]�89��wZ��,56�( z
�w;*�v���K3��q�y�v��r/�,e[�i'��+��M��T׼{M���r��4��>����]cH��#�&;y��%��P�� &վ[v��ېu�\�gN˹��F2��K)[�'e���x����
��ѝ`���	�G>Br��:Ѽ&t-鑉'D����Er�;읍���ɵt�7�6����u���؉�
��V$����-n�]G4��]@�]]�Zj��������e"=�XT�Y�N�\OC�F4�<��t�r�wx֟7��_εwvk��m�ab�}�r���|T�Bgo�n>��`�U�DgR�ا%�U�]����>�����G9���w2D�Hl��6Օx��-2A>
͇]�����c��X���A� ��2j;8��F�h�+(�4�T�o�)��pM[Y�A�Q�l��O��ۭ|�w�)K�өf6�(u�Wv%zݫ��Ovk�� ��~M�.pu� ���&Qk*g���co
:��F��Q.�l��G&A���ͲZ�])���촠�ǛY-���X�/��w])�71�I`rY���/8ƻT[�C�j���E��GF��h��0BF��7�����J�X1d��L^�N�Y�YG��9m*�Z\]�5{��T.�Vu��^=@���;-��n�ݳ*��mp"��}�r�Y�t�9! �%�u��\�#9��\�A]��n[SS�n����*�s�/udty]�M���e��O�k��9o
)#�xF�/����voNě�0	۬V�HM�C�Q���*�v]�T\����T�O+a��@�V�֚��Z�/�G�σ�}�j�>�,��~g:Z�T���sɽ�<�F���zr�v�añ��WbŒ���Rl�}Ko���RP����#Eu9N�mX�.�53��g�p��]�����0���0�^J�������*7���\p�>�R���t�_��#��YW����Ij���v_u���}���퇛qNHx��L����d
�5\���Ɔ4�Z����դ$̼�,�
��P�q5eb}J�~
�aH��1�i!{YIT*�G8����l+�<w��=�h��d#z��պ��x޴�t��5�uѵ�hnA��p�	����n_��v��X��A(��x���C㷖$KiR��7D�0Z�n��)�V�pn������Aqv+W �S[&�W<��B��,lY����h��)�Ҵ��-��w\�ĵΨ�8ٶ�v���vnn�UE/}.;����g���X�T%QZёV)QD$DD��`�D>lUU`�1���-��1��*2"��"�#1���
���PV1AeU��EQb
�Ab����� �����*X�b����X�Q��X�Q�VfXT����TTR"��lb��`�EdQ�"���dX�(��TX�����
T��@b�QU���DAr�V��c���[UdF""""�
�AD�(T�"�X��j�l�b�D��bZUF�	�)c�Q����Z����g�,|8���`��5 ��x�m9�Z��ӆ����S2j�Y���EP���2�TVL��g7MU�gs���o�:n������׮r�^��6D����Ҫ.늫�B������C\	{�Jק�KKso;���Ջ�oǦy1���C�*�Q�Vn�R��ʐu���],�&��0���}��xΘC9�Qqs5��W^���0ǯ�Σ�0t{�$�x���*�����}�=��Rp����>�}���el�LR��s�<v��:�0����y���}��i48tȐ��J�����?
��\*ʪ���^�6������h;�]v��m�������p3E��&7��h�w��y�\��nZ��2��:���ъS��qS���0ς�]t�
5�\%U�g�����	�_�<k�����h�E�_S�U1��-]��h|��ʥ�2�j�!RJ1�����3K�;���\r�A����ʖ�����.�<�f�2���*�������)�YA��$1�^����{;ɷ4����{�&�!���ed0Q�3r�=YU"#B��O�|fWX�`/T3�#�oX�ܙN;M�Юn`��w�;q�>�r�:ľ@�r�Ϸc�!1�C�:��FU��:��,n�?j��)�,$�����`<�,ĉz���5ݽ���f�T�nw{�ʶ����{apZ��(幛��(X]��E^�=Yyݡ��f��c��·�[/~I2�΄����TW�*t���>���[�A��r��W��~:l�v�ң�Y��Ђ�3�x��֙F	�h>�PK�1=��yoZ��/<�<9��o�ۦT/k�5�	�V�5�ڗ�o���x_�5��z�z�b�+!b�������x��z�|r����p�0ӳT���'�F]x�b�*�u$�eW�e�kw�}O��tq��_��Ϯ-���ӟMj
�ULZ7L�|7tZ.��]����u	�Nr�>��=����.�BW��YϚ�­��<z'�б����u��*�E��%��Or�㢚�.?U��s����+p\ *�Y���z��j`q==�])V��CS*��ɬ:Ǌ�ft�ޞ<OxʹhB	��A��	U8]O�dE���Rʗ[�W�\�w��U۽����6�Ҹ΂Tb�a��2�o��챭E4��^�+ީȈ����pnEld�k�hf�_�썭���:1����Q?Bj2���鉍w;#�>~�u��;m+�Lp����[`>0�>�o��n���P�A�L��Al��;qmoSЗ݇��9ϮR�`R��b�Tv���N�U�	���6�*���6�K�	)����]��;��㋫�:Ӵ��齭Ў���������ֻV�����i���������:�#n>��]N�I�Ur���dLfL@@��,�dt+��j�«8]2M��J-��1��1\�����.SS+_���O��-9�0�z�d"���|���V�ѹ}��kU�Ω�(�>�
�o�әGG	UE�)��J�g�XGk$U8�L��T�$�_yȶx"=���W�~^�yhz����3���C;�4����&�0>�'C)����ώ��u�ɹ�=�8�+t��`U[G�]/-��u�2�.Zpz[�dq t�s�,~�NT�uNO+o�&wl���j"�lN�Um�f��r/*���
ߒ{G�0tzWg���_<^�W-1wVjy��9��TE���4Ee-[^�QZ���:׏�O�jL���ba���ާ<F�:��������˽��ζ綝�����Ǖf&	�ζk]���6��Ô�tߩFOU�weꮇ>�3+ާp2UVF��;�W\TҼA������>�9�>�yg�}}z
����n�=\ >��&U������}8^�T�̮�X����O�i��va�P�@K/U�nu��)�.�{ɍ'��k����!�:ͧ��沴WDyG�{5�������%�og#�A�U�jKRWm�9�pf�/�_r�۶��-�D�"Z[]��;׹��}���ƥ*�K%�{GR��mgbǗ��!g¸R�"�ëAؽAnp���\��T�*.vT�Pw&�o�{�x�Sb�N���]wa��c���J���>�_��lĥc,��\};�Y��|$��vz���m�j������t��s�D<��*</���\ʥ�Ϲ<d�cs�k���|oYO_w6sN���� S��ʙ{޿IV�鈆:����x@�4k���Ͻ��B�%d�����W�/���1 \��twJ����z�X�Wa�x-�d��L%� |��g^���y���o��,�Q�K��V��[�S��7�8�A��f�!�\�}�^���Щ�׹�o�zt��C���e˂+�;k�@;����,A�\X�~�&;�"=C�-��zo��$��&���u���M VS��$��-J^��LeWm��ϷZ"eK���ו�F_����[�;�	�ʹ�c��T���Q}�}⾲��ϒ�үc�ྒྷ%�"͙z4�o��ό}�L�|ֳb|���*ޓ�#W�P�®"�#�]#�Y�l\J��e�� ����ǆ��L�:��u%��C@a4;m������{�Ƀ�b����*�}���d�oG���Rb��K������Ƭ��^R.Š���ݘ���=I�ilvS������hRQ�y�|������:�	výѩ���{!~��LT�Ԩ��(t8ӑ�nj�
��X½�9U�ԗoR�
��h��a��<�p^��p������)W��d��~���t*���jN�J�}���f���G�N��V;�X��{͊�V�`�}��>=E/e��n�>��}��to��X��D��5&*����N��x{��x�zR�H/��#�J�tc���وof�6�ίƣmG�0��vB���:�"t++P�Pϫ�[��~�So�v�����|�xl�������������8�!�</�˽FeY��J���2�:K&i��g7۱�X�2���}Op�:����kղ��ٳ�a�U�Ǭ�
���n�yxx�U��ї�=ئ�Ԥ)��3O��Y�T��}Bg2�R�+b]��<{Y���r9����s��6�P0s&�q�U4���;�soa��{<1}�}�����$v\06�ֻ	�;���Z��zY;A�UձV[&/���)ߓ��1�3���_�5�wVZu�d_4�c�bϽ�}�XB�[�$/���D��9�pFm<��z�ƕB-�߯��sLͱ�>\m�f��W�4x:��3�I��c�m>dri">�Ӥ�w�x޺庺�`�ā����뫑F=���Y���xhe<�A�3��a�}�ݙ�,O�9�T*{�t(Q�b�+�<�eUձʲ�0'���w�}Pz�8��%yM�ol^{��y�r���1  ���,�y]���r���+'.M����og^���>�2�R^CO�P���ʴ:������)�Y��C����N�4�2�ZVwy�<Z%4��h3�]�(��K���L�C*���VT��]���>2\'(Jw=�]���hb�r�P*�{۞OF���$�tvEN����gI�Gg�/^}��[C}���nol�Ǿ�F�J�@^t|�\LpS<���v�d'�@�y� �ֵ�4jy4�'Ѹ��dn֬|����ɵ��!<�ʖ��=�T\�~���W����=�������I���-ߟw��K�i��{��0ӳ�v���ȼ��:�I�7�5��e�C�n.��T[��u�.��-*��������wy�1h�>��z7A�����U߭��C������5S�R�}�VW���t��r���\J������S�PV�ւ��l����t�U�4�w}��9����H�&.\(F��=0n��wPpGVa;�5��H�`��WI��A��gc�,-�'v��/F�W$:�NK*!Vs{k��eq�C�����>�%�=���$�f���p�Ծ��/y�]�s;��3�<"�3�Ŷ�dםϬn�+�
���Dw�lª��jS��w�R�g*��j����t�ӭ3�=.��� ˞��R���$M��C�ӽK%����(�n�8�}�Z~�í�T߂��TjI�B��:�N��t4秼o�z��z�"#
���n�(ͼ��6��W�V_t��#��dl��4)|8VPTO32��_Yc~i��z$=�d�YOf����������ܩj�R����`��S�=Y�)����d
��Q�����^�Zۛszf^���jek�T��i�����꬙�W��"�&˲����e�b҈o��˗����!^����s|���:p�Y2���F|�v���ze\��:9/l܇�ި�����E�eS�#|r���������fWjpg��Pp�������^�?L���o(�cu���'��������yt�pL������"
�0����f6�y�Gql��M�T��L��>4�P���ei��'�x*׈�
�������e�g�V����u�Z�Ϸ�N���]2�G%H�,��=�o���Ĥ)����d��u���+F,�urS�z��W[�M\��prB��"sw�7�85�,M� ���y|-J�;r>��]�o�Z�\���cc���g4X3�5�^���z�e{��ۯ	[b�t�xd��zz�5���Ev]O/5s9��x�LE/����^�)�C�y����cw���G ߽�W��Pñᙳ[�i+��-�x��m��ݘ�z��
�����	�����}��o,v�PWJ��Rr��RG����X㋽IX�b债��U�.B1�� �^�*�ڮʡ�8`���zⳒ�,��s�"�{�:ںwVʫ>E������#<�Brj��;*VGW�g��os]N��{�׮��+�C��Ft��k�ЭG�Ԋ����C��%=�ý~����K�o���"6tU��;=(�����*$C𾠉�MQ"��J%\k��r���/mE꙱9���m7���y��P�8�[x�b��	y�?#\�q~O�!;y����C��]z�9�c�7�a�=�=��=pV,�2�<���4%\�ʖ��'�=���>��oT��OB�j��)\����Ռ���oֽ1��w�%�[�.��ߌ�� �'�e�L���+w:�"�1���ut��F�:���|�ø�&�w@ÙVɂ��YdY��D��#��":_w��e�i���T�
Ü���5���O�>�sr�.Ud��������Z��բ7g\5ܷrE:�����ut��н�C$�[IA�4�|O�3��b����j�(�@�qT���4�k��ì�;�F�L��$Ҫ�I.Z<�~�L5�n!�O�9�7l��	w�9��~�mg+��@�r��R�U.�@�uu_x���ڤ�4�٫!ܬ���^yy���������)���^y!��P��'*ޓ��5QB�4��؞�^;��oP��>U���z�����p�E7��)QU�2P�p1�#�4/�5AHRh3μ�x������c�	��7��	n�d����dz�{��m>�m#�� ͿC����wƥO\��{ӗ_	Uֹ�~���yX���:�%S���#˗����Q�N�tf�
��&��i������{��7,07���H1^>��*��-C({K�����0\7��"@S�>減~���~���LO\n�C)�j�ΣH��*�У�G�6���	=]�å=���]���%�2����[S��������܃�x���:�JK��Wh��o�j{Y�r*u��k��l8�?��.z�7��&�҅Qƿ/y��c6.Y���jF��yyi�W9nd�=,.X]{�QZ�k��|�^-7�V���z��B�^�x�w6�,�@�Yy08���N���u��EKrvHw[�P�f�hXUd�9�م"�sVΣ���-t��:��8BWݶY�*n�9� r��{*�ݳ1���<C�+�5��ۉ��2��Ǹ˻�yJ�W.I�q��3O�Y�T��}Bg6U�ճ�Ȳ_I{�P�]oa�E;q�O:avGR��]"�Ɛn�ߝ�9�h�og�<��a3��#��C;�����H���摡|Y;A�][e�b��1Z2��?�jc��=��^ўQ+Qɽ�����fp�dOPT)�B�*�.��qةp���}|Κ���gA�"��Ss�c8�M�K�g���<=P���QA�XU�+~�g�!��i*|A>Y��X�}^�o����ޘ���bϛ�D)/!����P�����)�Y�b�
]"��o�&m�N����p���#��y`~�hC��2�2(왎�9a����LJl*X�f�[C�����E��P/�:�>~껼�;�g�wDI�*�슝��:I��վ[����1�o݇�b\;	����4!���b�3�x�����<<"�0>�kE{p�Z}=�,�W������GQ�:��L2�
��^@���Ԧu�7�6�V��hR	`�`�Д���N��Xr!M�ƥ��f=���Q�1W{x�*���i˺7�먲���i�O�N�#�d�Tlm޾l���^�����q�� �%�ޑ����MB4�d�F�Ŭ��&��7�E��6�=.�*��ult��~�gE�nV�+{rX��U�I��`U��l�SX��R��X�z��i9�wlͺF��S�V�W�EY\�hӗ��n��}�":����7On�.~խSϊ��/�(��'�f�w��:5є�무�G2�:���Y�8�jr�'U���S�H�6R��}�"����r�u��E���Ļ�G�T�����܍��0^�VcY�d�eFZ�㶱�k�f�奪�s[�i��*0��em^�ejX��s��쮓����M��\��!��K�R���Q��e��v����.�R�gy������#:���%�,Z��̥
���孕lit�f{t��Ѝ�ԃ��M��3��P�.�:Y�YYK�e�h��:�Y·�p08N�1�����|��_�a��_PMY��59��GgoS6���"�Wq���.����um�F���]ii/���p�A&����B��v-5(��U�a�!��hY]Z�L^��;#J<=ףDq&��
ꎹ3,!��5�n�9�qAXUr��WM�uKӇS�f��f��A[-�M�L4MX�C���� �W�m1S����Q�k���pB�{6ȴ��[��z��q�[���ܷ���ڒ��Z�'p�NG A��\�4���ǳ��e�"��̊�n��Q�gr�J��@T��,���7���R\�&�.ҹ�5��7���&��z��<ھ�X8�ik�kCp������B}��=��V�(���^i������{�!���k1񠻻v�S�S�X�\r�ȞҾ�F+TWe\׳s���\>3Y�v�!�;c��uǣ�}���"����|���b�����}˅j�N�]#��*���%|�����M���cE����l^��v�X}m^�x�R]�,�]���-*	0ͮ��秅�J�ci狧4(|�n�w]��ǒ�2A��n��W)����VK�Ob��.+UY�҈�;�Z]��Wl���Cb��5�6Q��z#f�x��.�pP�ZWmJP�OJ�n��&�&Zޔ�+�oR'�� �9K�Y��k
Vp�����S��a�;N:.MO4e���Bugf17�9�X��VE��Z� �.�V)U�ͳm�pԑ(ց�n�˙�nYE���ɲ��`�[��ɅDj�]�1�`a&
v/Ul
�nr��SXu�_�Z��k������TiJJ+�t!�<�J�j������eE��=��d�[�z݊�̨���ZM��
����B��B�5���hZZ��QQ!R��TY+Q[XңB�*�"�X�iTE�E�"�-wr*
2(�7J ��imX��)QEU1[���V�
�kE[T���*6�b�ыh҂�"�V��*�F�U)TQ+R-K-��S��Y%����K�V��R�-���ڌUT[J�j���V�"�T�Ė�-J�c[�(*+��j�X�+Z
[jT���j��2�bmV�UDڨ�[Z������m��me���+YclV�ZX�l��V�*aATn\W��W-���\��+TeB�ؠ�iVյ��V��jX����V��F�#JŶьkTm�-U�iQYR��� �Ee��J��h�F�9Qc�2�1�wg>���I	�y(��g:��֤w�w���!̀�b�H��r�S�V��]7np,��8��s�ww_�~;�a}ݎ��!<�5綥��
�֣!�f��(b�{�{E�������v"m�1�oԧ��+�i����p���f�JK|d^u�*�S*p�W^��F��?n,�7dW�BV��]^�������/NT֠��LZ7L�|6�tZ*��jr��Y8��6z����`{ή�p]u]�,ÕM|�V�d=�ꅈ5�Uxش�z��D�R�7훽3Y�Ҫ�B���j���p�$6�0�g�OOt��q����y/s�k�3���$*z�*�ʠ��;5��<�D�Ɣ���.��M�#��cl���K��lw��y�vpNus�W?N�	Q�~
�8�'S��t5p�i��PW��g���rxd�yŖF���Âg5�fl�#��F�Xb���O32�����r,<�<�s�&��Ξ.ݑ���2��f�U�����x�"c2b0X�; �\<��{�׻^DO-}]
6d�j��;�y�����i��n���˘{=�L�IK�נDV+�٣�j*/3J��U���J�q;[�u��{�|�]]5����YDȍ\���k�[(X�Y�-����/T.�9��ޟe7Y�r�d�P���뭫��[�y����ټ��R����ً,j0��M��h����е�y��Þ�{��G.b��]�O
�?�Td
���s(�aÕL��*юXGjK����ʽ���v�^\�y�j2���-�f(��e�����ڇ]�Pp��Iн���ҽSi���<����@����⾮ĪJ�d���o�����e�\4X�;'�X)^���m�S��������ą��K\��r/T;����Q���}����}nxӪ��S��MbV��5�|F���]z\vƂ�Z���axL�s"�[�^�n�j�2U%���y�k���U��O.?s����̚���y�]{媽3(x*󉓞�Lwo�V��: U��3��g:_<�j���w�׾���J�ᤪ�l/��2P�<*S��]}nfW�N�d�w��ǫ�9��w���5�7�HM:U�.��A�Ȁ���r��p���\�](8���u�=_q�~<�ﻹTE��W^t�����P�TK*$�t�(p�mK�W�NMPV�4��A���4�n��֫#L�Ly�xw���_�ti)��l���=*��N<M��F�_-��TJ�S��ҝ��b���:�� <���b�P̵�LNa�$z�מ}�\߷��+m=X�=��5�i��޶�^%;rjH8�V��7`M�.����d]\;�w [�O3��m����V����Ȅ�s�
���r��η�q�n�yct<�ryV����}�]ȵ̋W�aW���f��f�s�{���5�m�Ϣy	����T�"=�)�e�z�%[�"��<G���[���/D�j���{��1�4�#,�.S�;�e����/����z������<��K���ӄ�{&f>�d/`XtL��\��LEj�zF��>�w���Z2�Iy�a��؋fٚ�K��ӱ�[\|�ܫ������Hd����RPw� �U��������W��VH]Z2�r�KW���{8hc�]��H��*x�5kĪ�|"�JUV��7ؼ�YD����Ԭ���g!�A���dr��R�R�T ju��_Wr�	���r�3��oL	���³;�Q>jCbC��2�4F������2�oT����ȷ�D��V�}��C������wEZN�WG��J4�xF�[pf��*RY3�p���c�(��#���Z:�L�_����Z�c��}��Ew��a|`+z.�͵�҉��Rڿa�����l2V.K��+2[�T'N*����d�@���;�]^ WU�v'����v�g>%eb���8���ܝ.����'����I#u;E��!���1��"�޺JGu�J=��/�ѣ�.͗���� �̭�~k
���nn{��)�3Jd_�D�^�	$HW���"">�^�rx�=^�J��>;Y/x��ܯ��g���
���x��	���p�~�����^�����ݣ���n��Ӫ��}sui�6-C�ug�ij��i���r����)��7Є�By������V�����2�ӓ���{r��!�Tx_Nٞ��#e_�x�ž@�xT�WOL�{frnu����׶U׻6{�1��lS��7�vx<��3�� 0s9w|&R���I�r���3O���aUSϲa�9�͔����u�4d�R��ӷ/��ƅ��Ԏ��^���!4��cH<��?g-Œ�*^qp�2�0
�M0�U�<�x5'7|��*����%١�œ��i�ĵ�0��j1[�S������G2JBf{/�{����!����%�;"p��r��
s��.��;)R���z�X�-n��ωs�ۜ�=�W�w���^f��3s �"��� �GA#�u�����X�)��}j9v��]ղ���uW3��<��r�:�giif� 	���R��׵��]+��V�q��n�v��h�g��Q�dS+��x����+)��z'(V�u_K�v\76�r��;� ����Ʃ��:V'V��̒+�:��Vm\g��f��SE�r����DuIy?B���*���0A��$ x	��hn��:�Ha����Ӟ1[�U��x����b�eW�\W�f:�z��Dh|����{\�~���-C�N�`Vvb��{���{G��t�O���*EN��w��烻�(����gy'��>���u�g��@^g�K��
���<�|G|tX�ս(q�gW�͹��g{y��]��I��>��x�ݜ�f���g�s*�
eq�FB����r�������/��Qxv
K��Y���S��a�e�;9�����Ot��ض9�:����*�J�RN�V��.���!w�N�Mj
�LZ7w�⯳�nx ���:txٙ��jϥ�%VJ���R��Yf���­��=G�z`bs�ʂ�O8ww<��c"�J�y�[7��&�(̫��'��Qu�. w����{f�S(8��Ux�5���{�^�H˭���q�.�i?qN�&#Sϫ��s=��#�MO�dJ۠8�:�xV6��S��W��Z��65����u������)��Y�Qlo�8e��(Q�)�+W�,��p.��㔫7�.��#���i�3(q>�HWS��/J��eM'�2w�V�#6M�L��������s�4�B�ܰ��'�jȻx�����|�-_�'�޵0��TjI�B��8��h��ME4�Y�����=��V�wtg5��"/��:��yឣF���m��a5
bY�11�~���#oD8�qn	~���8,����RN~�T�S�=Y��0XU��8ng���m3����:?W��5u8��b��s��jek�KY����\����2�ʸ����Az�Ͻq�ǽ4"S�<J��)�B��� T�o�Әt0�Ȳe?T)V���	��=���؜��)(����q�T��g��Z�c�=���h�N��-���2F�y�_���^�`C�2��m�xmCk�E�\.��u��g�fS��Ӽ�Rчf����G~�A���G�dNU����<Ѻ��#�O��=7�I���h;z�#�̓'����^��a~w��֥yǄTE���s"�[�^�n�L����.s�ȢǶ�~�f^#��z�d׭k�G�W��zfP�U�'*o���F���h�v䶠ܿj�0�����[SF��[h��&�a4p1e�3��
`'~e.&� X�|3J��ͥۊ�^S8&=N�eL�*ug��v��d��;��ٜ�ۓo�82 J<��J�2��8k��[�`(8>d�cI����Z�z��Ito���c��b�Mfu�/����잡t�h�T�c���U�(9��]h�^�ך��M��6�ܖ8APz͖����w���/x�ظ@}{lL�SxF�G�
	zL��|��i�����]�G�|+�[+�=G\D�j,p�������z
*��cS������r��R���~�ۭ�^�v5�ti)��!F��Fw����5+nF�|-w�\��g�[}O����U�.v6zQ��ȇ�"Pj��P��d��<�L���娚%.J�n&M{�v�甆L��_�����t��D,�ݕ��$;[�׵�w���l��r�_F�F����x2|��u>���0�Ir�]��dLi򲢽��ٻ�m�<Y!�4:&Z�]]*�\.����Ƀ8��bџ���X{�>Y�[R�ޝ������d5���h]s�*������}[���}���/���S��0���nz�3�p�є1K��EWQ<D�����U��|��y���a�@��j����.��8�d�:f zQ٨�PZ�=̠���R9�'�6
X#��.^	iřw���V�ud- Gz�3 ڈ�ܐV74����z��V4�]����#�+U]4�I���Ê�iwFA{����$�I�'`�b]X=�iE~�x��)c�V���6���r'�t���m���D4Ǥ�x�U]W�*��:����+���`V7w�s�zk�Z�+��Vgt�%W�Hld(:Q~&;#̡a�����P���L��<��M��mܳi�ˁ{�y�w���}�i9Z�*>qJ4�xF���kj�vS�����΅�~��Ѿ�yd(hg�i�,o���A7��eGz)k���q2N�)�����55���h z�0�i��J�X�zQ�[O��ǭ�Ba|D���!���P�=���>��>��v+g4�5���>;���T�+ӣI�z�
J��iHUw���y�p~5`>�����?^2e(�<��3������^�����1�j�:�k�������f�o���X��~�WI��W���3�z���QqW�zrz^�nA޼D08�K�T�巷=}��n��n�)U�����%=�97�:��..f�[*�ݟl��`js��r�^Ԛ��ɱ��g�@�!$�H��I�X��x��0�>SA�UU+M��V���NCI-��c6*>�8�b�n�fR,�g� Bn�yi#��]Kr�C�/Im��q��k3a�8�p�N��gZ�vhe��f;�EÀ
ڞ��
J����v����Z�S��{�q���hW_l��8�!\�cG���]!R��S>�!�:��<9tX�������ߓ�pV�U��S�g��wv���62w���}P�El�*K�C+�'h/�[.���-��b�U���W�NK>��S����m�.T��P�84z��g�D��)���P��/��R��o�M��v��zc�6��Ä�O>F��~����1���*F���G�*VC0K˂��r�ow==�RUU���{c�e72���i�w�zQ��j���i�8����������"P�¾���yH�x��?kB=%�C}�z��w��J�P;��C8�����iX��6zV�*C��q��;��c����߰���&�nG?
�<C�f����]�t���]W'agdl��4�<�\LpR[��[�����ʑ�~�]��{mG�c�mVT�ج.���2�;� P��N�@U\0!G+r�9�����X{���e
^~�,���lOm��W���<�� c��	�S�P����t�5{�Q���0U����j,���Dog!F�l��Z\RDxqa05!؁ﳛ�|�M;�W]/+X@s�We�g6D����d���oDw���I՝E�l��n����F��l���ÉH�7��Lp�k�\�}S[����n�����V���+a��jbe�0�{��zrkPV��-�`>Z9�f��Ǹy_�q���%�Vc��=l��eB:��e�q��*���=�螘��b�a�e����>>^��R�~���{��,�K�)%�����`^ :�Dw�=�
�q�[���9�o՟�K�q�<^/�Y�CS��q�t��*��yUf�<Q �!"p50�YnZ�efoZ�S��o�T�E[r�Vz	��*5$�!XgrN�#�����R�����=�ܜ�jc�1ﮒ��/�S۝Os��+g���4*�1[@fc��h��ɚ�7��kԔ��3�SL>�<ܵ\)T����觎{"c"� �8��ݸ1�!?mvw��ng�K�^Έ"c���1��h�/w�:X���V�~�g��||}f�Y�w�R��~��Y��دxJ�E��Uv�u�)����SU�CN8\Y2�uᾕj)�;�����5^�UwmH�ix?DIU�Du�K�E'IpЅ��m.䝠�����mQ���B���[Ȁ��w׽�A���<���F��E������r�"�t�I�)��n��Q�¬v9u|��>wj=���wf�6�:�2>u�,�k�9Q=ʵ�o��c�&�X���:�yx�}l�r^�L�(��4�́�:�-�9v%���ATǼ��T�k�|�M�R�шm��A�����P5��6��B�NP0����^�[�/�{�:�����;tZJ�p��LCۡ�=��+��P����+4ݸ��vwm⚱(���V�MYlQ��~�=�g�][c���dޱ<2�gv��MS����Xy�W�yw��N���6�JH�T錛�^�R��*�sTaޜ;iUM�\�N�[�L��^8�:�2��^�P>���s>���Q��\KM�:��؋�$�:ɗ#���w�h�/n�Sa]�.�=H27�M��9/�zE[2��̣֞YC�+�I�^�	t��
�X憉Y����k�QΖw��y��T �I�㺵�%}ysN�����*]m��rjܒ���͐���1��Y�q���58�*�K��ŗ�7F���ZŖ��%�4�J�ck��kc�O!��f�bv��cÝ��5��]�0�e���8�3p4�%ؓ:�1M�N�!(�G���𔺵zq��K�WGR��.88t4qN�Ft�5v�iU�7d���1�4ݚ$ͺ	U���[��:�1���� �uA��w�ˌ6�?r+�w��ZB����Z�Κ`��r�^c`��ٮ7XvZ��Gy���,OhJ8=f�n���	��M��f���U�b�dv��Iᕻ��37�XR�Md����b�/;Nt�)Ct�Z5����������43nG��� �w�g�bάT�T�|4P��w;U2���}�(����s���kY���E��o,���1at'Q�rw�i��G'~9�}�4�����p�W�-Bl�[w�٨��5��v���he���G1�03�x�-/]u'a�˭��N���9O(�:����9��>�uo**��m��&�s)i��c	��hA;����`taPJ�j[ۨ�e�Z�N�����Iekj�fn	L]\�p���t�qڤ��6fI�d�:]�x�ќ�4WM������Z,v@lFy���TT��Y�����ӕ�ׇb�^�d��u��C���(i�\]_:bK��xI;���9k���r�s��1�Vs���������z ���b멖x�����ξ+0�h�놬8Cj�RVlS�Cv��x z�C���n��T�-�՝�u`���Wt8�Ilө7|�ч�HF�/�]��WD���t��a�Ρ*�V�[�]�ʹ:'��[�P(`�M�t,R�}vx���x��.�m֬�l���X�ǒJ�'�O�҅J��{hct}�(:�f�_�9���V�f�}�7ݢ�B�L�[$}v,KɃeof�ۡ	�}@O�is0�+�,kTTIkJ�R�kldh�b�\�PA�Zն�R�,T-��Ĵ*��ek\��Ե�J���(�ƈ�Q�-mEm�nY��ܡ�UJ�J�,e����V���eF�Qm�E+(��%R�U��h�JZ5l+mm*��R���E��l,��+����*6�C2�drV9B���q�XұZ�e2ܠ��[�*�֊���F��kKV�6���&Ze�qZ�UQ+X�T��1)eEb�V�ڲ��[c*	R���-��F��cq̭�Ҕ-f7�V�+Dm�4�e+emmme�miA��q��aKZ�U+J��Q��ʣ�`�6�[V���(2��X��[F���PiV ܤ �P9,E�X�۩�{����>���3�H�t�����o�љ���-�va��hie�A�`Ŷ�2�>�M�Vɍ��0m����9`V�U%�������,u	��/���S�+�luJ^u��:a=��Ogt�#��� �s *�,F@UNU��;#��ץm�f�h�8�T�$���N��TsFN��Y^����|V1^���
�^"0x���@���azLvEo��A�2靊F�,�T� ��v�{�O�9����2��<����^�+�e^q0y���j\���Oqb]��q�4����hשa�|��.K�yxu�~���N�WC��e{�;��o��ӼQёG�nOww,�N>��F�Q�V�l�蕏aʫw��ƀ�B6�� t�1왾�|�rxq����ZU�Br�}�4�z}�ˉ�,����QW.� � z�cyg�b����^�gD�*.vT�w&�z�e_����bg�x�a|+��f�b_yQ
Cܦ�y÷��z�Oh,Ot�")�Z ��cgj�U�9�ȇ.�ch��?{B��я�g`���ح�)�wO��c'>��,M�N� _Os�C*�^���IV�Ξ��r�����꽮�J	o�zeבR٭\u+�ʣKy�U;(��+�����c/�i��EX稛]{b�cc�>�ojgc$.��C��ꚸP�-�����oaj�
�bw�}�G��q<�S6��Z�m>�F�rPJ���]%��@�ૢ/o5�\̓�ػ���5rP�S�������3�xg�t�w��8�����X�X����Ǌ��wQ#��к�f��b3�tX�\.���鷟;�=��bя9�
ϧ�Z�9�/m�*���iR���j��d2UU����J����>��y݈w>�l����e&;��P�R��Uu�&�X�$��-J��W��jp���p�����vDr�@�6�NU�#%��]��S�.����n��c$7�M�N=�M�n��Z|=��Vg��(��P��/��zNF��`�2�~����ӹqt����i���N��,΋��y�����Y>r����(g��cN,��q���n&��c�߻�`����HR��0��ih�^�L�_�Q���_�+�O�[KT��}�2��b��I�^�9���Q~e�e�F�W��m5�ǥU��И_)��!̼Kڒ��7t��m�|�ֆ͉
EM�X���x���k����1Xu(��������=G�����'�����8v�5���T0��\���ܗ��F!�P%��4{�絧phLū��5;�.(;���L{ŧ�e��+�VN\�,1Ʈ��hʆ�v�]��o#1̡̞�!S��zc�vE\�a�cN��Xitc�f����L'�nu�ݵWQ�b�|'n��Ѫzjk��n�z�ܫH�
��ʳ��b�b�[�#�~���	դ�Ш�,�>��l3������<\U����{<Ϯ,:/�޽��4��zRj.s����oI1�n�p8y'vP�oП�zｓ�s�e(��
���0���>��ph�(�u!���2�%�ҚB���6|�z�q0��؂!V���W���f�q��vT�t��Z�*즑⋲:�<&�kA��*~5�;�sn��s'z�3C٩(VC���+����{��s=g�8�Fp�wL��4a���i��5lL,�	��}V:�y�TJn��}b�O����wP�88zzfp�}�<8
wN�P�Z��UY�z�eA�S)�G��9���ω�;�5��Z�/3G{�na��u(�ܘ�a|�}�����3�X.M�4m�j�nݝU�i唕N*���]�s*��Q8.�K�r��������P=�9^O6ٻvD�A]�U�6+�Ǳy`~�Z�wL�L�
;U&c�L,�M�]����_�F�7� ����.��o���V�R�%��k$�cƅ���Z�Ά��X�<��:����c:�f,��e��	-�G�	4�g^q�-�l]m���VV��+
4Y8p��S��q�[��ݵ)�xԽ�wա���{�Lp�9E��U���׻v�u����"�c\=]h���@�����uwy,vρ�� H�>�z��&�zE�z���mz��K�t�Gg����)�ό���iQ�R�c��� ,Sh;t33ݧ��on�����h�l\�����3k��!�<綥��$Աv�w��O��~�)h�5���X���P�<<�Dd˯xΗ��r�x"FI+6C��lzώ��񕊘��w(z��l2���&}mL>��zrkPV��-�gK��p��Q�f�5�s���M	�'ܤ�a.z�/�]A���_8z���=�螚�����Y�3og�����q�l��E_��Q�l.;I-�Q}��}޲ل�ן=����:��^�$�ܞ
ڏ"�~���,�L��`01����M�U'n��z���u��g#+�7[yc�ѝ,���z*�3KW�y����U
5xd*�e����isF���掫3�s��<'&��S�PW�Yg���}=�<3�񁢾��GcHЫV����*i�دv�DY���Zx)]o��;f�\��K.�0hѸ��wM�p.����cu�R�ǫ�|C��3H��1�A˶uG�{7���ѻ�5L�M
����²:p�-v��np��������\�Z���zt�I�7�(�=ZnZب78�K&l�o��D/VVT�w�u��54��z�ײ�p�'?{�z)㞬������[�۷Tw��$���\��� j��ӅVp�c8���J*���E��`�{<D:�/�':[��ݹ=��^&�[	�/��J���*�1��*k|��á�E�)��4mu�|o��r��ӹ�ޮ���g��N9�ʸ�2�7],��r�U����EC3�8�K�T�g<ԭ�{[>�i�cg̤�g��[AIg�Sĩ�w�%����YSv��̽�Q>W�?a�99ǎz�J�:&��*�� �# k�l]����2�>�B��X��ുY���rd�u�>�[�~��X�I�Z��N��uܠFלxFU	��9U"��/*�A�W�n5�⻧���]%��gג��·�I�]j��#�V���xz�Z󉓟M�c�w�n?�d,�5����R�jͻ�+q�c@�@C��򛾫��%ר�ڞ��K 0�\{�L]����=�龹<�\TҼ��Cs�g�Ö�AU�}��#�~5�g��:Ӟ����s�v'S��N�l��#P��z41	�.	M���'��hi�W���n@���{)*�z��{�}O8`
��y9��9^�ry7�w?�3g))����Ք6q�j�X�{\mn�]Xs���o��c���.:���|�r�W!�J���YO��ꆜ/O����ϭ#��Y#,ͫk���6�ʆ�/5u&������O�I`�L�j����pw&�l��i��O��K�鏸��ݮ�����ٹz��Y+dײRN���U=�N�"�U� �'����s��*$C�k�($��(���fg�k��!,W"EHR�Wg'���,OuT�"	�j���r��U��f_�j`����}�ʹ׈�9��g�T5��=f����Wf>ùg
#W�l��-���m��tw㢒�JeL8�\�НrpTL�̸����L:ٍ��D���O��p�m��Q��_��`\��V�)sTi��h_;!�Y��J^������n���-��N���i�b����U"=C�)TUu�I��/�Un�DB�����f�sΰ���1��c��]�!A���d�*��T��UK�P'�]O���=)W��ϟq��,=̗^��OO�.��8�+�$6 ��mS�oIϺ 7Z��|_���IdK�3���1w��zb��Uw)�ot���խ�I�[�W���hp�ga6N�/(�f�r����1�i��0�E]q�^+3�����d��+���UՑ��evv�9�����s�֨��� �cA�EZd�r_ǘѹ��)]�s�p�׻�@���.,������%�wd"��{i�~�r�8�	~�{�W�E̵����{a1��LS�jߡ^�U���L�_���U��c�ȏ�_���5l%���';OVSRo�U��z��['l���yZ��~��њS#rT�A�������Ȕ���B��j0k+��|v�^���Z3N��ʳ��,W�Y�h=��ي�uGX�M�r���GY��t��KZ��ĆoѪzk&�^�\n�V{�7�=�<�M�xV�^�{��ܑ�z��ԡY�5(gݢ�g*�C[S��P�m+^��N�g�%Ü�[�q��7;w��Z����h���1�-p=&g�Ju��\\���I^������n{�u���r�M�ihh��!Ϯ��v+�rM��3^�i�L4�x��Y������"�푷{i	������\)Uk����G�.��	��]v9�J��r��Ӱ5���_v�s_?\���T�{<3��3�0S��l�*(��|Y;A�][+e����4k�����;W{.���Rn�[�f��H��ݗ0�Ղ4�u�����Q�G�V��r�ɽi��X3d2}:��b<@��f��DLᝤW%� �L[�AcV>�](L��n�>=؃�����V4-O�u��a%���'ԟccf\�'`?|��t��D�v�������dKFw�ÁP�t�
?k�4�%,�7����}JI�"��=�L
���ƛ�^n��h�S70��0."����b�kv�DֹY��=��x�Q��L@���*���CY�X]���p�i�w�zQ���^"�ᣗn槭���pAObCF}�E� �¬��^"������s;�Q&C^ˉ���+��n����!���ژ��g�M@T�Y����:�1��Tpc>ܩ�N{�ml��n�>��QTڧA|��8M��GN4�.�ѳ���/?�*�)m��q;c]�};O���|��=�@�w�� Uy� ���G{�;9W�[6|%q�0}���~	��=ˊع��ϫ�i\V��z}���.^8l`k��Z��HOo��wR��=��{�S��Mٻ�Z��p��;X�
��RN�
�e:����mL>��zs�AZ��Fmɼ������<���3�0偑}h�l�u��_I�܂��y#�QS�Ζ%^��	�X�@��n�Q�|M�h�m�k��`�\fQ3��ۋ��7�Il�1�üq���Z�l�vkW�͑��]�]G���Ve�ɁҺ����Ӭ�(9�6�ܺUU�9ג"[3�W'M.(վ������ãGގ�U�0�{����\s䖏/ /`^ :��Gp"��_S�Wg���[4�g�����Ή�iqŲB��2�f���u;���7���yDd��z����[�変�]?��?{n��ʳL��^�7�t��Z<NPuD�1}����S���Z�>2�`�=g��QM>��
��r"*���pL�c���U[<�즑�L9�͋�_e�c��1�)�^�	zxѭj���ji�K���Z����`��S���(LH�ߓ�l{��I۽���Ր Vrw���B��y]�����Qvib�ᕬ(<R^ͬ�Inl���v�||e�ɕp*�,���Y$�]g܂����0M}}��;��Ѿ��_�)�{T=O��xN��ʑT�*���s���r�_
�Wlr(z���z�ť1��q��x�>��W��ϡI��r����K>-]��yX�	��xQ��*$�'�u���zeֈ�y|=Ztv�� �,F@r� lvG��U2������K��{40.}��xX�|�soy�{^��W��U��Ȩg�:��/5�wG�#=Σ��f��!���nl��C�&�Kϔ��o8뫙.�J���q/�ټkJ��I^��q����b�A��P6L���+U�f
T�t2�1����Dk�(��c���E���׽�J��g<֥yǄTE���4E=8��啓6�U/��w��i�6r��>y��d�Z�^B:�V�����mw���a:��9��ި��Vٞ�ڗ/j}{H��<�10r�%d��)C�[|*V}z���y9��Z1w����y����NGpn�ǏF�*�͖�RV=��u9��`R����r���ޕ1���o�@���yn,�N\񂹞��V�U�p�Z*��y}���g�q�i�yu�Ej8b�ﷅ�H��n���~�u��^��~�i���
�i�����w�3'���f��zvY��ϩ)C�c,������aO*�Qs���t��r�y�.�o2X�wo�;���z'���)��Es7.���'>���};�T�<�2�^��J�w��|��0�0d��� ʈX�!�Th����j���
�1��\���X�޹�%=c
��j�a�Z��\�u[���CGO������~�����}�s���$�	'��IO� IO���$���$�P$�	'��$ I?�H@��B���$�	'� IO��$ I?�	!I�B���$�$�	'��$ I?�	!I� IO�H@��B���$ I=�$ I?�b��L���lL =� � ���fO� Ĉw�$�R��*��*��J���(*�R��@"�R�D�UTJT��D�TJJJRIE
JRA�JT%$��U�ʢ��!��B�*-0�UER��֪�D
�)ta*�����H���P�jU*CYUI*
UR�cU)����R����
�m�A AT���D�@������4A@�T(�	R�ETU(!J�"@	�E"�I�;j�hԢ/  ǩ� =]`4�V

����Wc����ڴ�;Y�@ta�.�(�+��lhtV��f���`�4�.�i�%JE&��(���H�^ ��"��u�U��]֚V���¨�rT�Ӫ�6��w v��vv�t�ݚt��gWc��ܗ4�WGv�m5�()�T;j�T�JJZ`*^  �懅
(P�c� P��B��a@P�@(P���n(P�@(P�m�n(P�B�
q�p�B�
�:n(�
B�÷
N����Y�"�5��W+��WpI(TUPPD��  .�zh�=sX M�qՇ\Tt:Gf�@km�wgr���Ő;��]����ڡZ�.���Fh�MuÐ����JJ�iR�   �z���]�fm7gWw �p� )�:��w:R��۔u;��k�i�(֙wTƭ��B�һ�����`˲�'[7�(!���kB�4���R�   6<���nM�� 5�\pE5m�هA�R��V��wUݔ;Z�mU��f�.v���e��:�n�@�Lv�8��JR֤R���5I)�  &�N�:�Ҭ�ڀ�H���Әa�҂�vť7`����Wgv4��gG:]��r��B�`UҘӮ�t)Ͳ�t��H�QPET�̓� � j�B��X
 6�l����h mmk���  �U�P�� #  ZK P�%�%%HT���]�  f� �  ZV ����@ w8� ��@eIQ@gG  ��P�Q�P5�0QP�]��TQ �� �� 
�E P�  mF *�	� ��� �V� Pm*� x��T�(��Oh�JT��  �����  O��T�   j����U@ R"cU*	�##�&�[*�^.��M\`��3z>(H�$q@Fs" �ywj:�?g_��}^�+����TA_�}��_ꂢ
�* (�������Q���+
�
)��������Ґ��?��ʔ� �%�y�q:Ӹ�/���q�Zqwr�v��P+%��2	o�ji��2n��X�m��榤��k*T�w�E
ݗE֥7Q�<�K[��8n�u�3��؜�X��YA�(d��K]����<A��N�Z�M|���"�l��c��j/c�U �j���-4�[b�Ct)b����m@�][O�Z�H]���{�vӓ2�F��0�9��r�$����H�ȝW7>/B�̼2G)�,j %�U�>L��K�{.Luwa�w����+
:�'�D^��Kt�u<��1��������k����P�̕��~���ج
 �N��%浔�[�a���a\�v�� g��u,˴�.4��3�zR@��ulll+$����x�P��z�-Aƃ�x��"�;J�R��̐����U���M){��l�{Y	,�*Sr��G4�!�y`�t�N�#3C�A^��m`�0����P��"C�`!���pԭ#r������KaNe<� T�V B��	܏f^#l�:u�N��#Uk�A3K)�:�im`b��WX\�R�4�-+S%�n0�/r�9�. ��pM���3]�J�!��!�Ck[����n�w�� ~x��÷1����N�@`^Z�(boqd��tݬ�� �Tf��#B�*⧇u�Z�w����?!#f��R��q 1��#t�Z��wa���8a1HV���62�e�es��bI���g3S��I��`�u�ЁP X%m�&�m�{�V��+TW�-R��r�xޭ)�z�}0��Ի��WN�ik�X�˽L�̎���߲�+�;��TYS^Q����J�YMөEm��6��a���+{�Sױb��U�b�k*��JI��U��)*�h̥�l�}���mVEOp
9��P�)��L��;ȶ������GXw��6��`T(�9v���=�$�x���ԙ���$/)0�j�8-�5�Z��m%X�u<���Ďf����i��<nԫmb� 彗�2��*����9��qNSX��%��4r��iY!���DRvRƂ�42fc6�V�ɕ)�K-�[.��-���gV�OU���T�q:׹eQbLf��Ȳ��b�y��y
1��E{>WV�Fg��um�/��JC� <@��^Gu�)V��YY��u�"�
��ӊ���ly�ԳCU����Z�&��(��+d	�U�c'�,2�.�l�P��s	�73�*��D���9B]�-=Z�#�5��و�r�V�~5v��Ō����]9�p3����(%4��51X#cn�۠in*�s,i�n-�w�2h�
�ء5���36�N�{z)� ��Z�� с��`�PSW�M�ʍ�bv�D 9E1���N�K
�j�\ڻZ�
rbbj��j[C�Ξ䝵��[˵Xګ�r�]\�wF���5bV�3�ð���2�N�%(RDSS+i��v��aI���0"KB���n?�F���5�֌6e��~��S)R%��������%��bƨR)��f)v
y��J�Z�)�{��%�[sic?�����{wkF6Ȱ�O�@���t��W�^
�f3/v��،�ۂK�m�6��d���[q��Т7d��WD��3V�����۲��܍�yC��$xo��`�k�IYu/tH�Ϭ���'��̢�u&n��U�q�j ��<�٪�4��'J�Y8F-5��0V��fi�"�4��2PNXj��qJ�RQ\v�^Ӭ�]�7��+s����:�Hڦ/O�t����'�L/���h�bh��ܫW���)��Y��;�����%f���Ǧ��.��V&Ҳ�M�2IwUTP����YVH�?�Y�Q���,Z�����P�˼Zk3ZSݙ�����M�b��+ ���K�(�9��6X�����Ɋ=OQU �ͽ��Q;��϶%�p�܆Ų
;�0�ғ]�h� 4�j^ݛ�e��G ˔q޴eeK�bI	�Z���m&^ˠ�ӿb�%g�v�n836��h��"6ڗ��Z�3 I�ʌ:݂��@:�ݺ�Hv�������h̢i2�%-�IZn�fm٭	�	Y���E[QIP-ڰ����Q����P�= �������wt����.��Mי���%$�ٽ�S�qQ�*�[��u6��W��.�����0f"��^�#"B��8vn�ʔin�[�|��"�[z�IL���$���X�ק~L����fP#Ͱ�j�C&��N e�(f���M�#N��Q�����(����2�.�^:Ь��(Z-;t����"����;�)����kZm%f�t�`Ҋ�+�9N��N�yQ`����;;.V��Cae]�Ձ�B�%��r�f9���Kee� �Rb�%+W͸�Kblݤa�����,7W�V�5���L�0S�x�m��؟73f�۔)��A
�f�aq=��B�jDE<��8��;[L5�#�:`�CS�`,x4�
��1m�KY�KS���̩�1��
{vJ��Vͼ��r��m]�U����AW���4 ղ�L�V��n7WZ��ׅ�j�Rm�S#ܷ�%��U��ҽHCSpfi�(���i�� � o �X�(j���{���WbnٙW6���q���nͳ�� �j���3�^��Vc�;&��hQ�M��[������&S���J�`�4�� �uyyP
����>+Q���	�m�,[wx�ܕ�,�k(����^��:x]-��ܧ"A-סM�kt� WB�yt�,�F�L6]&sJ6��K���mIn�[�'�/cU�V��,P
�K���^��skEjG��h��;��I�()�z.Zb����LSN���%ҭ�ƢŖ�����Q���N�iK���P����!�ᐳ��� "n�=F��4/Ft*n���r�&�l$F^,']ަ��F�ZCz���ˬ7��3�eYͻ��%6�Qi�u�6�V#S 0�a�7r�鬤l[�jG�m�RU�dEʁ�/�MmJ#&:�[x��J����nj�Q�l3�hz�je���a�ł�l^FX"�5pDV+���w����0[Гyc���#�>̏dʈ�JJPO�U�d�2�c��Gfًr�+���3�A^*�*�T(�,�t֗*|$�9��D���j,�-$��ji��ٚ�])�Ԉ�t�8�w�����k�Wj�޶6�v�恄��y����N�vե���u�Һ"�?.�)�XӲ�K�A�QFm*Ô�N-�\A�ͣ��
� �1eL ��v:wKF�u{�c�������@KJ�e�{����MJ4���;o#��n��haw�2'RZ��e�8^ -�I=Uw`��ƙ�\h�b��f�Aki��l����4m�gaX.:2�%��#IӉ�el�D���͒����Y>�+qT8nPe�!��=�E����TĒ��e��0țB���f�Y��&=��Z�F�L+�n�&��4�Le�J�%�ݑrԽ	ۛ�v���BD�Yq8U�%YEԔܤ@f�:��7��.&�T(��y����6��
��wm��)h��l��9y��)2wa�����J�,���V� �j�j����bZ���ὤ��qQAG)n�,DUH�Dl���5b6SN�����1�Ce'9F���Ya�K�aݭLʐ(�G��p�@n
�bڨ�0��#��;&\z�Ւ���m#X�-;����⪖"����ܱW�-ͧ7MTh���D��[PM�Ƨo\��8��F�j��Z�A,���(i%�y#�/t�%56�
NM���Woh%�i\�Z�U��2�T)wp� �nZ�kMT�3q�XǢ� ��.Sʔ�rͬE�k]#ӭlb
^��-�N�hW��U�$*ޅ�VZ�u�y"S�,ݧR����g$��	{�)zrR�3jT�I1m���V@1�Z�ĥo��M�[kVPDe$q�ʽ�E5z�X�/f����3L̽�!�T&��H�kn�գC%Ȧ�� � �AOj[�;�+@���)Q�4��ٷXDJ!r�֩�i��]^�w"M�P�q�v�+ܰ�4MFcE����3����c/q�D�`��ա�*��B��7����y4l��A5Y�4�$'V�e�3/f�4Ś�T�m ^Մ�%������i=��͟�i�mfQ�WfV;�wr��c�&t�6��������B�8a��bZ*�jS���,
v�f�d ��9�݉c
S2��]��-؝�=y�"�af�4�m�5�B�9����N:'߭\�VX%�q$ŧ�T�34��1Vm�{�B�A���i�&���W2�[��q V��| ��ݺB��I��ʌ�9dʵNY�I	�ow7znc� 7���f;�r�k+@2ݻ8Pr�$�Ѣ͈7ʗgk�Lt��Vnnj��)0#�DV����94j����:"�g ��T�<��e�9*��w��A�sa�P]�$[j�4n��a:η�8�oP����ꐺCL��vp}�M
ծ�7j�7jK�Xǖ	6]�=�E ��m�ġ�4d*e��R���ҝ\�S,m`u�L^�m�`ݻn����͂@e p�Xע`�T��Z(Fce�̘(��vԭ�7Jo��Ԉ�Hݔ��S#@轖���fLI�mn �;Ô����,���$��d�	��a�O6���.<�e�A��6n2j��J�Xg��m� ��7D겣h��UP�[�
�̨�U�s]HXll$�-Z�:�<�j�`)f��/[�@ՍS���;+ ��rԈ��;�㥱$��f�^�Zt���R:�T��F�֋?���ΠAʠ�ve���"�ڊ���m�n1���u
���%2K��m4b��)a��F6Ցn�ʶ
�kpMQ᚞����O%�f��%��a�m@�t�j	�vM����(��ࣩ3���%��n,�&�j��@�3xn[���LB��E=щ����ƌ�:��F,�����mC$��d�lޘ�]�1/�i�!��%�F9i5hކ� ����3T�� 1�@��T��/�ؑ#Lz���ok(l��6����%1�	(ǲ�OEUX.H�ý&��Ot��`m ��K��	��e: �ۻQ�'�l*9��U�"b�Y5���V[��RZe�%e/I��V&�Ĳ�2��J6�Z��.��[nnb�J����%,=����)Z��� !��6PŊL���B\��c�V&de���okj���EN���o6���u����TY�
)�2�� ��:�i���R�P�a���u���im1��ૈT��PVR��fK�n֭9�ˢ��\ʑ��*@���{/]����r5�YLeb�
���W��+�yu����r�H���HS�l������H��q蠲��e0
M�Gl#sCڃ1����1ձ��s�Eȉtt��c"�a��ű�ռR�oqr�p��=m-�x5�*j��Z%�0(+M!���R�wwXq�P�n������u��̻�v�,V3��cNc��ūoF<EVV�MpXi�x�5����5��IE��M�,q8*��oeb�`�P�p��bM2���/5��XI��p�k��J&e�/^�l�t�i���ݗO�O2�Ӵ,mnj���@]l����*�ܭ�N (�"��#�Gҷ&�Il�wR���kp��(�C6��hn����*�7
�jmc�zeІ�:xt�cUc�ؒ�R�h)���nj�-`O,��Ѧw4�Y�6���[Ƿ��-�f�
5��F;RD�pC
�J��P|��E\t��!ŵ��>|�r�w:7 �5Y��[��X"(�Wj�f�r�:��j�	U�)���UށM=	jT���h[��];�Wmm���,�!��6��fE�l\)��U�l�kD�Ъ�U��5�ۧx�d\�(�p&A�����,My*��q�$��c��\8����eT[�a�BHob%�s4�tۻ��{ ��".�V9YX��e�Gt�yH�y�8��u����"u�J��݉I�`��Vf��B�N��bY��9*bՉ+M'XD�3��kV���5ܗ��(�]���l��}s��K�1]Y�@���#։�Bs�w�U��N���V/71݁�f�u1�`<$��7�V�b���pl�,����X7E3@ت�쑇L]`ˬLKe=I��SBT�ɰw�"��ӛQV$J�Em�آT�����Lf�n8*����9p20�C-ղ��Xә���\�1]h&��*Im�[7+]/��nPJ�H�m�6'�l��H�ae�[49�I�L�ݲ)S`A���� ��P�T¡�\�D�`BT��ĴnVhN��hi{t-;�NQ	2��ie��
��R��
Z(b#vG�Ɍ6�'`���x~u1���:#��^�λ��m�\z�w+jp/+��V�2[��|U
q�J�ۺ�S��i��mk�Ĉ��& ���8���i��tI/��{P`��bv~j�2U�uEq��Op�V��8����*޻�X\�U�-���v���c�2$�-�u��찖�&��:� ��*�:����b�Zd���7]�),���U�f�`yL�]$ĩm�WY���LE�:�5�M�ݣ-Y�,�1�Xi���-�m�֢4�[����e�,�Ʊa{�`5���u��r|�f�c.?ս�H�Q�Y4��2�&�������������-��R�i��9Y�	u#9_5��T��9};�tk!XQ痜�\�lU�&tԒ+���ڜ�yf�S�@�_V�ܯkxu[G�.��z&op4�f�-*�k�9��ε^-Q\�V�Ƌ�a<Y]��}Z�5��frU�֧�e���RfAyB�Z�g���j�ww�Í���[��v��0S�QQ���\�0�x�u�\7�4�����0䖥)�N�������|%6�i�GkWʎ�`�&е'l�k�p�����s� 4�V����K��k���+��Z�����k0^,R^���FL�ɷӠz��A�v��[Mz�8�U˛c��s�pl��[��Kɗ�zbO,^�N䲊쮃J���R.,	�Wۚ
��b����}˾�ӵ�<�Ǘ.��6��s���� *NG�V�ZZ0����͓�Y�Le�"��,���2+��M�M�]�iuݷřz�${)�7�d<Z֍��;��Ϛj� Ǭ$zpc ����-��R�uo����Sf���<jҏsGlf+��C�����c� !��:a���7e�00�	�v�儝qo<��_�z4�S��
wDT*�V��b�����{��(M�L�����1�M�p��hV��4NeFyY��K�J����F�@;��l�*�K�R�{�>��c��j�m�K�9� ���":����c��$�/���.�st�K>�ϵb��O`f��ju��-�Ӻ�S��l5.}{N̰�ov������l��!O6���V<qw"��]���PT�xv��e>9��Ӿ6�N�ӭ�G;	9/��J�,C�k�f�ѽZB�r�6�+���!u5��+׷�[$<��Z��05=-8Y�R��z&1�̭ťroK��k�%�"�z3�f߆�Q��n̻�#Nm��c��'�p���)��+e��i5������b,�l�|덜c��{]���F�3k�_���]�v�n\����9&j��m-� �T�K�8Ʋ�3 �}���,�T��Z�Qz3��R,�Lǻ��hִ��ɜ�7��H���G6�K+��1�G&�9[�������w�KB2!-<��s_o�iN�Z8���˱�w�C��)��'E��A[93�vkW,[�L֓�q����k�72�[�v��E`�T�Lw7�:s}�dO�����=dV�Ҧo�b�����󮗔r.�
 �:x�V���t�8t��umۣ%�Syg�zdҰL7�u]����ٷ ���6�dؒ�gp
w"����OX� ����0�
Q��!YWg��u��or�ï�4+i�Q$��K^�%m�*&[U=B�9Rs�gEAlm%:��s/31�ф�;��Y�!݈�W}uѫ�՝��u݇��r�U	's��"*+e�6K!���f<��S3�ζ���:U��-��r�:����s)����M_*Z���;`��y�b����y\�8D��M�z6�r��}���c��i;���,�`�C9�iխ��{�ooY}�b�:�8C�^[V9ڷ�Z\���Z�JH��`���yWI\P)����V'W�B��]'C�ש��X���8�Rq=��d�((��E�}ԠZ4�n���(�9��E��R�;����^�1���x�ݗf��3v��n��tEj��ʇ{�v�������I�=�������E���V`�p,m��"ɫ�΄w�΍ٕo$Q�-a�fP5������K�b��2�b�+nkݱG��"�c�*�G���3�6�O���oK\h�}x�r�6Nqފ��ݾk�19��ÓF�[š�/�y���d�Λ;B�B�1G� 84�$L��v�n�g�jF�o$)a�hr�q������ ����o{�'���٘�b�;��c��v!�n����z��Ӕ�	QG�iu�Ƕ�%��s�'����a����&
��@���Er�v���Wn�miK�D�'6.v���T��7�o����I#wAU�����FB>'̵���P\x�u�,Ts�V���������z{'Mhm8�jU�b�����Y���hZ�a.��t��!ov��0q _F,�����J�#ɛt�0MV�d�o.���2��h�ݶ:԰�Ԡt	(Ia��8�=I�=v�
���ա�'�vs}�Ya��gU֙��ȧU���p����<��D�,�/�$�G�Г�.(u1F��cm\��wnܸ�X:��:�+((�72:�iX��c��i��]��}���P�Z �ƻ�Ѣ��]rdf��Rڼ���[�����^�J#O��̲�r��̎�b����y�}'I�w�ZB��06�h�pe���t�B�=���4��w��ҵ�hq��x(��M��BC�?R����d�tg�LG@T��^������C�Lz��4����n�7x�`b8/fW)W1r΁����rݾ	=�W.r ͳ"�}ljc���ݚٗpIr��ˇ�t�Sf[�Dt�uoq-�]B��ފ�	�l�L�;�@!:�vs����4���ȹ�Y�����{6��1�b�=~����)
a7���DU�n?5�r�/e��D�m�옠n`�g���+9*��]�F�r:<6�&�)Z�x��oea�j�� �`ju�+�q�+Jovt���e5�z\Z��κW(����^��ϥ���v(Ϻ��T�^K�k�e�[ F���811QU����P|����VN]چj(�Ar�5�ΰ�s���5���:S�[�jsz� ���J7Y�����g�-g`W����\O>�a�=���)k�[�� h�s�L�-V���[p�R���6�ѱE�������v�o��	e�ͽ�0��Nkʺ|s�P��wǒ���X�uo�Z�g��B��������3C���Q��������q�c�$��8�|E'�s�F�6��Y����4�K�LXrlr�;��o�.����|�7�7 �N�3nO�c��tn���w	@�6�T����B��)K�Eޅ���ù��ɅLi����a��]@1�/�$Q���v�d��������ϬK�k�;r����ù{�s�)C�J��;�4�0�6��&+���n�(�<�h��2"��_e��o�bJ��wpm�;�w^)�f�.;wpL�Q���:/L�ӭj����� ��ˮ�I���!Q�㎸��f��Q#h�}XZ���* _*�W^	+P��JK1n�w%�˺��W���ádt|ND��[�j�6,hLLʶ�y��^v߆p׹�V������,)����9�\ٮsk�fG��s�JlCE��v�D&Ca��J�=�t�c-Ż�E�%�%վ��p��*Mc03���Fg:�d��e�L�0�u�Hڴ���Sh d��lkÃ�PI���|_j�N�R�]#�,�лf]�k.�F�IR�f�]
߳"��DJ��l-Ҏ%o�m��ق�)+�9K4t��nu@ɵ��2�v>�ݷ�C��d�O^�H�tr��� uI�dnq�����J�o5Y���>p�͍;�����u2��.,���G���Ҏ,����_\K#�W>�%2JL�H�i��}kh��u6�̵E]��*�Xԯ>���1�[��s�.ZGl��&ȷ)�BtT���_eN]ڷM�.iv)4 "f݆Tk��N�W�%�^���ڹK�L,��u�@\k�pڊuJ�fvP��s�2H"-����*Qđ�=Y�X'�!*�۳=�m���9�u�&h������u���}���h!3�%cOU����=����֊Z8	��>�/�!h&�6�fnMP8�� ՗JGHe�t���3�����e���Ŷ�t���J�uʺr��]���̾�pv)��#�QF|�R�Q ����WEx�e���޼�pv>}|��X�.���诼�?���S�>�Y�R�+�����WI�WN��T�''>:�5�Lb@�,��;�)ZC)-ԛ;�.ZuZq`<+1r�BJt׍)�z+V�gJ���g ������N'��+ǧm<��=u˪�D�����_ׯ�䶅���e�TyEeb�Q��çzX�2��1qtM'�l���ήwu����{��1����Ӣ-��Wj}��!]�<�H9��T��]�L �������\4�P*F^]r�$/�D�7P��Y�LBb�Q"a`�^<�L4:���4�����w|�!�Si��*嵻�n��T(9Q��y^q�	_���e'����&����e����X�,�ew._-�5m
 ���Mr)o#��yc���ДS�#�n j�%��v�����PgY�G,�B�L�Ѥc�K$���P\/>/�e�,�\�v�0�@!��jᕪ\�ʹ�2�qKյ��]ԝstق���f#�	�X5�WP�	2�m+-i�\«s��5�dGk-��J��p� �JV�8�2_e�̙���;�:��%��S��ܺDش�/��������O�.⻵��֡��ì7�hVb���5�N�f5����e9r�F{9�r뚍V){��ɺ��$B�:Z�x�[�*4�)u�e�tS%v��o��5Z���Ԯ�s*��Fev�l�_S�lR1��|�����ʦ�ߋ�r��<V��eD1�����*﷓�\����=p�0J�*�s�x<ދ��+_u�oxM�V*Ď�4�3����z��;���6*�Cmf%����붾6X��8t���YS-�s�d�4V-��x2�)�s+HYes�ݻ����h��ֲ�t��l>����vЎ�����l���S�\�k!@\��i[K<T+�����҂���bN���e������&������sݑ��.(�OsAiJ/f�w��V�f�b�kjcouG� dJ`��뫗���ZBo&�ȡ����s"�*�tf|e�};��	���e�%DQ*��@���+4�a67!��`��Lu��N�^��s�'�.���%+���e���'��Ɠ��R�*S�5�N�77����6A�g��;Y�,:K��Y`�;�A��5�j��0: (����v��S]+pK�q�6���U;u���2ŉ�4F��x,᮴ս��V�v)E������ܽ��r>���On�q�s�b�,9�ɱ���-�=��ܼ�:��Ji�\���m��th	\έ��-����wd�נq�J�f��l��G�21g��e�+ �j��7`���bf��3z������-P���ݢ��pnX�]�+�T�r�f9�a$�O���kǵt.�@����uu9�7�Ěܮ×v���kPr��*���4I�*-.�r�K���S;�c��&m8�ǻ�50ܾq��7��B�r+/���wK�{��1K�^�{�t�-��u�������٭v5�T����;i�;�#�W1��'ű�1��gp0�7������.L\��6��(r#��F�=7D�W`;f��`��Ԩ���������ܘ�\(X��p7d�c��	�8�=��d\�}�v_�q�- I�َ�C�"L�]4z�r�VZ�x�[}LN�#h>���$ᵐt�O:�'Ho1��M�8��H�N���]֠��
Y�[b\�p2ڛc�`��Y��JYD�<�@�Z�o��Em�a.�7G��+\͝�m(D��!�wM��!�t)k������ ���Y��鹇+	֌�yǶe�N��li��Pu5�)u�rb�a͟eg+s�S��H�-��tq����L�tmL�՜�J�ig�J}�T��I,\(f7��:�8�\� U{��l�f�fH[&��h7)�d'w��ĵ�z��5�}yN���po��Ϋ����<���4���`�4b�}]BG�x��]eo�Ws9��M�t3������Ed,�p�t���K�y�f_Kۈ� w[+��2RݴTk��N�, ٮ|z�#v�/XW�j�j�[��3�@nd��]��e�R��Uk]M�a����{���b{��_e��ez�Fjd ��z���e�N�k�856;���HR�<�I�:9��9�����P�B���iM,9�U�K�6�2�*�;"륮V���Lm;�[��e�)����4�ui�ج��!��/�^��ȧ�>d�0���)a[cO[ T�|�2�X�0���Z+��9*+�1j����x�P㵂�w^��B*eR�;�Y���4L4�D�/�+��͕b�(f>ީ95(XKe�}��ݫ�iYDm�B��Z]�ƪS���eM�Mb���cWX�N���`e��]���8b4Vjo�wAہ`���G���E0�&;��u�o`(9�FV�1�0��:~�A-�뙧����1���D����of��I"��MN�F�`�-y�򞂾ϔ�������70
�r��b�p�jH��wN��j[�s����]+�V�r�Όͮo+��px��[X×ƍ��kRC���샯m����<z[]]��xf����EL�*�pu�0n	�h�;�R�ᨵUq嶚1]z��;3P�-#��z{IXbz{���,u���{����Qύe,�=P������s�׷kl�4���wh8댍u��Y��;���֮�۹�H�9wH�Qײ�y������g.�Qg��z>s,쥪�e��ࡤEm��WzR�� q���ϏW'�ޡBm o
���sy�NU��"����f�s'H�}������(`v��m��-�@L�T���f*����X��M�K�@�vaN�+1r�us2�o�*�xй��<��\)���dRo6��@K^�(¹�vR��X�F��oAW��Rg#3��j�٢&��r�Q�xx�x~������������TƜ檄M��!KJt �(>��X�j�@�����.a����N5���諓ke�8����:����_u߲��3�=|1q7��ZO�!V��}ui�R�k��p��i՞���]��qjv.��]LL�3k��GbM�PYYjH�)���Y�r�n>�e�d��)��¦��Yy}�%�n��RJ�7V��X�V�-���M�,�ZN�x�5o6�q4����ϟ.�.��]�O��
���g]/�o	�� ��5��mL5�'QT�ֶz�4e@w>�u�RV�&�i� )�l�t��Q*��M�/�N�;��]��r�r���ה�:�\�NP%�i.XWW"�ýܩ�FT�V[�Z��<�@�����ԝ��O��ޑ��|#�}'Y�GumZ������F]�|�\�ד�[�re�����]t����2�든>5:����3���3��)������:<�`hmS�6�gC/^p|����4���jr#Ҁ�3h�N.;��m+�`"-e;x�9w9�!β^��������j��q9�1T�Gz�A�fm�2�n����٣J�wys���J�`u�@�Xי��n�Ɩ@2��� wro:�X=�N^.�f�Ú�6�ͬ=B(:�����Ŗ%�B�[ݎ-IӰ벗ac�]�C�l�(�@kO�,�qq7`�6������t�<��P&�!�c�(�-�"�m���Y�qg4�����tm�4(�R���l٧�\��ZŦ�Y���%�vը��-Һ����D_T\�E���q�ޡ��Q���ٺ�������Y�W�Jn��a5[���$Y�y,�����h؁+r*RV�����҆��&b\~[K��|�a�����Ӯ���޺>h�Q]f�s5ҷ���H�TE�S�:sB�.��R�����ӵ5����JW	��b����>R��u�ˮ�q�4V���&�4+�
Z4�Aڟ<.�4��!��̙��9#B��e���ĭvȦV��\����:uJ)3�d�hj��V�,�Z�7$��A��e�U�`\!�.���s�� ��wȧOWqsxsHp�`n6�A:�l]N��f㸻.c�-�_Tڼ:Hn�^CĺrՕ"��!��}5`�\y>��[(�%򅝤�U��n1A��e�GiN09ԭ\�� ,n���q�U��)�+%R�M�L��htrŊ�K�]��A��g]+W#���gMR5�jW�d�ÉZ�6�]��-���r�K�gi�}�-jV�LCz���XC�\:
�Z�n���*�B_CA���l;C�]���AC�쮸	|���8�=���ҋ�8s�(n_P)��D�%4ؗ]v��	mb��"4bvR�El�ބ%���.Qެ�h��O)���9��޷A�!;�U�E�nح��d>�αֺ7�`:`��)��(Ͱ���Mjfv�#�%��iVj���nB%����ֹ�����nl�� ]�ҎE��m�����֌�ĵ�]Pڃ,-�ա��d*�!ʛ�+�� ���[�;U��㷅�3W3Fe��YM�V�î�a�����Iʚ��{��j��n��;tA��F]�{��sV��;A 7�"+&t����t�����EX���-v[�Bc2�Q�9jQ�N��n>z����^ա@�(o1m[[ :�kO�- �.�i��L�r�u"�4c�mZ���of$�m��\�d��[>�����2�1�ֶ�}�kp�V�JC�u;/�;KaeX����Ӭ#w�f4�2Z4=�5wE)�e�-�x�/�V�P-�z�J�Y@�|�Y��t�n���,�﷐�Gu1��f���y���۪-ޠ��d٠��-Y������-9����Ie�M1�w��M�k�I�e\�;��������Q��\��b��:��7�5�-�	KNXÝ�!B�v�(�X��H\�>�`����u�V�	��:�ԭ������Pp��$a}�L�o;�d'�+�܂�vG ���u��{�Vn�ٓc�ҋS.a�CPt)����Wg;��d�Y��u�C����{��m;2��|��*iv��У�z1Tntc�IX���L�/�k$�l�ѭe��dz�V�j�5�6�o9S���6�·�ɥL�r���vi(�,�ywlV���^���0�]�<,��S��*$�e��&���"�+,k.*B������\���MH��)`����XRT�����f�Js,����ԁ�]^� �EՔU56���|�)[g6TK�n��"p*��{� �����1p�P,B��.��k5��(��k��5�7Jup�εd��NGf;Ղ�毟c���F�c�2�+�*�ja�4��C�/W%q�]Kk)��o>\�ׯ��n���.�7���Y'.T�R���l���(�-Si]� �]����ܺ٤]��z��:��]h����p�1�%�i�ΰ��9F��3���1���_+��ms=����f�g$ 9��Ĩ-z��e��3��<`��`].�	+�X��!�s*̳m��ǀ�3��'��=2�\ͦ��}F��8�bWbYv3ƍv���_b��Z']\6�:-=)�>�xFU��������*ݹ��M����j�ۏ����H��Sgo*�t7�V�D��پ��T``��l$r�8gL���OGr{:�6�����k��ì:��F��
�G��"�Yo�Jt9M[��v唨9���9��#�ۗ�n����G���L5��j��h@���o(nb ݉��VE��}��	2�l��-h�N"vt�;wG.�*P2�b�����s	}{��Pz�V;�6�7[�} ��J���+��eͬ�8��%�����]����.��n�+f��3Q�B�f�kK��g3
��AxP\��,�鮽��郰�s{U�����-�]��AB��5\W���Pk)��\�(-�Vkc17C-���gc�vG�NF(َ^�T�5�q�MD�������=X)V���Һ*���6L_a�O�����Qաq)ˮA��+�^W ��7���:�i�9ϑ�Q���W�KF�Wz��*O�uc�q�K��ʝoKs4��uco]<�D��V
9�$���x��v�ZW��U�r��Z�Ok{_X�+v��FRۛ�1�g,�i�JJ
�5A�����P�r���j��\"0�ܡQ�T�]�fcdu�5|V���m0;`6��̹���r6�#os�c|tq�T��@ h������	�C:[�O��%)Im8;-^)g��/��1$ؖ5X]��7h�MKkN^c�ǭ.]�`>� �����:�O�6�_U�8j}�|C�ƧgLo;�B�%�khj�v!���'�-� �e6���}���;+��X�=��]z^�P�����T�C�����)��i���ֲ&�[������-���
�[B�C��ĝ��rr�gX�t���d��%�W�u���ս���P��^`����9�� +���Ƶ�cY�Ʈ�;��dr�a�'T�8�[X�j�q�k�)�Xs�~���Ut���=���������_�,��u;)g.8�psث)�y��v�����k�i�&�#��)�������b��9��r�˨ü�f�e�t�|�qC4�^��4��i���*#S�OK2��"��)26���L�8�֕ ��Q}������%\2+�D���3q���!��	&�1;�u���+ �j5J���Ƙng_Z���32�Y\�.�Z�y��&�r��2cu�	�j�r�vd湍��@]�ïnF"�q@�{PϮ봁N��f�l��Ǻ�@����9*�F�d��79���V��Q��/��ۮ�{�a�Z��F��qD	�1�2�/*�Op�:����i�c@a�vt��C�! �V��%OQ�k,}�A������� �w���e-���2�;vj�郳�vS��-���R)+�pS�%4.�Sj���"��
qBu_K,b�t�fwa�Ӷ��GwA�+v*�W�#�;̜���#���6�eƊX.s�u�R��阹�H���5 �v7D��[���;�
�ɢ�LB��W��z�궃ይ%��u�_ BY�D���d8�vhd9j��'f��_[�F�%ηl��y����}`�Y�J�c5m�l �pc0f<[�Lq�Q:�0^)�h�]DBS�f�������.��'A�yԃt��[{���e_z6��G�C��w]{vV��u)�^���C���a�[�l�86��P�4^��Q->�"e�s�͇�)?��M�;݁���أ���t�c��JT˔���*/����uu7�}R�-�vw�
`���h�s�q�ͅJ�{h�M���tsXm]pl.s��Dn�>�|u�K�k7�m�GֳC�(J�_F6�����ތ��4�(w/��V�y&-��BY�h�iԂ�k�8bf^�8��·I�s�|��؀�p���鼬����Z5-I�h� �3�3R�9�\�a�!�A��r�:{�)=��0��e���(��P��k@��/khh)<W'շ-�F�&�n�m]�:+�e_m:�����j��ep�.�ͱ�Z^��/Uo�=Gu�
��k�5�l��ܜ:���p�o闗s�Q��k�s�֭�=�:v۽����2����ڃ�"�W��P�]ګ��Yksli�'���!2��c:ҦL��+�:�M��k*;�2k������ʕ�hVP��#٣�8��\�?va9����n�BhA��2�сt��!���ƙ��+p�0f��0������s���ld��� ��-�����;t�X�ݲ��V�������R'��mՌj�AjMr�n�z�ewXӵ.LEEs��em-�<�5)�gO)�/2��%LJ�g������ǋke�s��u>I�1m�9�(2.p�[�y`�O�`���֭p�w������z���ۜu�;Q�����kw�Se6�e=EU�G��.�
��㙶�v��
`l��|CP	�A�1�0P��7��t��RH�EV#9�Cpѥ���>� \w-�n�q�x�fh@��5=}'�Ow��\��9kjG����
�����v��}�|��ZK�C�3��\���γX�°!�����]cH�z
9�AC���W��1%���w8�G��t����ڻrU�$C�C��T�U�6����ZR�m�86�u��h޽�x̃ �}�P�'J5����E����̦��Il����̀K�qN���"�{��DEu��Nz�=�`s���`=��鹮R��Tydp�:�q*v9�TYΨm��tp����ٽ���ܴ^��f���k�� 	��Ʋ
���#*`ѻ���y�l��9�W��G>=Y���R�`u�r�/��T���A�M��ؼ��q��ج�Έ�Bf��/:���Ԍ���/xS� 2:�^�Xr�$�eev��zݥ���j�x�t�.#�*ag26�'^�Z�/X7'u��*���èv�6�d̀�xc�}��T\�uJ�\��v�gS{# ��ͅ�M�*���|]DEX�H�1
f+Q�>��˼n���[�_�n�;A�gTܢ��@r��u�:p��N4o���A��CF��]
{�A4��i�˼�2^8GN��؝ �6�ɳr�Y�t��\�h��*��q�y�q�,�U/m`w��4u�B�*�|��ߙ�GZ�.o�Z��˗х#�f�l�G��'+�rp���M��b�[��>��Ϟ�j��\uv�ڜ9�F�`��]]�bEI� ��`�eJOnE�mw]�ufPA'�)�h�죠��9��j�f��Oh�b���+�AӶ��2�m_.�{���M3��X��-���V�Ӈ���eX"F-Q�RIB���Hvo]ǹ�)�e��VRD��u�Q�'���w+9}e���g]���Z�t"8w1�9�i9������)>fD�:z�ӪѡY��MsW}�3���'5���;u!�l���S:����v� X[������ǓthفS�±V�>�6�S�n�}KIK�ߑ�z6U��ѐ��y]�6�8�v釰,�3�gV�6����IҸ9���]�����e�F1���O^�1�����.�t��6��}�u���ňr@*����޽���n�E��4㩁��%>��T���)@��\"���Sgn+�X�T��Q͡��h���%^/�:L-�z���V�[u����[C}د��˥�;�$o����j�k;�kbu������;�Y�e@e7Ypaڵ�-��y]�ӃKo��ǽA��� E�U���R�'�Y�}e���B�Cw�0&�T����v����V^պEXc�M�ف�m��~�d%\ֱ�/�[ma�\9���oV����ٙp��.M�ɥ�O*f�R�cZ^tg1�9�wIM�V�%�n��%�T�*uQĕ^Ԣ�ة��v؁Nk��2�m�ʥxn�G�юV��D:6�0[.n�8S�2�*V���؄�̎�JwV�bՕ5V�+v鼦��p܉�(�l���Xi=ƩP	���y�@�]�g.±�Q]Է�q:����l�Zp\�,���b�Q��/U�eDd&�]���,v��&�1/��y�]�8S���J�u�f�zhe�%
H5�7�$�b�����bs��wݧ�#bTNq�R{���!��H�玅���j̜^�
��f�b��3eb���4��/	��P�/ ��:���-奻D�,!V+]�����-�%M��#��b��qWhU�8����V��0U�X����hSmo"q �9}��X+GMj���0�.��F�F�L��\��ׁ��=��z@���t�ٷZ�G��]�'g��#st<��A�YK7�p�4>�ɒ��jغ�c��\� �E����:ѩi������ׯp,�t�rS!�����f�uom�
h�(��PUnרg��Uz�4�X�t;��[���.J��1w<�h�@��8�tz�Tƛ��t	:!��L��H��y[� ;I�_v@F����[K'gR��p��TQ4��d7�mY4ݾp�������:��V����+�z�*���p`���Fr��OCؗqZ��*b�V���#t/+�I1Qч*0J;�gh�B>0۝t�̫P\�剪'��v�2��Å(���gt��u��je0�Vz�@��{~M?{Z��^�Uv�s�<w��*vt�x=���A7�a�c�6�R�:Y���]odK������f��l_F��XV
k�I�-X��V�q��n�sU�&�����=.Eĺ�q����Q���Dgs�ev�[`m��^����l��u==r�D�'�S���6�4fS�Ή,�8��y��W%�]�	Y���n`]������B�V���6]���Ԧ��d�TL�(jT��I����{n�Au�m�#1�i�.�]�y](�>��)Ϫۺ��l��7�F�ns����FwQ�nd�1Dd[>���R��#��ܫ��қR:�/�����������o<��u�BҔ4�!AJ���r��B���*�h�Ȥ��2D���ZZZ�(�\�Ȥ��J\�
�
s02)�2V�h)��$��*�B�JJi���������,���%D��!ʐ�2B�
��\���,�$�(ZZh�������!0��2C*J�����2
Z�ɳ�*����i����f�L�ɤ��r2JZ(#!��))
��������JB�%�"���CG�w�>n����|��
�vS��ع+f�b۬[�wˑM,����г�9Xh�\}�kҬ�\Z7�-��r��uۆ��_%��c�p\A:et��j�V��bs��0w�҂���R���ɛ�����oHiW��h���V[K�ut�핯st�}���篘��~j�ж� �{΂����j������̺�.�cc�Om���l���۪�u�:�ic�B�bF������}��8Q�b��R�w����cT:���2�;pI�d�Q:>{T��ؘ�=���kRD[
�r�3��v���Nc@Mv�:�s�/�J#�&�1�ִ,`IƬ�.ܛ�h�u7a�a7-�ɦm]�jJPb�1��]��)����8��N�o�Y�[7���)7��MFCf�tj��q&�щ�2��%��/�"s)N=o+��}����C]Z�f��۾Y�q�������z�8<��J���<�w �t�k9�ь��Ƹ��7(h��Xn�ޠ�[����a�3�0�=�3�Q�u�x4�\��V���y�鋟x�ƺ�����MrY�+;{�6��:K�����-�"���nR\�О<���fJ/�������'<���ݺ ���n"H8��n��N�[A�]�5�͉�JBp�ꮖ�_s��S��=��#��w���66[�6��m�<[�.<�l�a(�e���-��h�(1-��[M��Ij��tM\���>Ӭ�-t"1���֫��c���l���E	�6�=e:[]==[5{�2FQ�AlcG��ݝ<��;wiw4t0��%�J��kݖ��
V�諙F\M��R����ձ��E$e?C�/oC	a;��J�!�Ĭ�7���C���ڧX�6)�7��>�5iT�%�W!�D��V�h�dnV�B���w�C/��K��sM%T��s:ӭ��!�6g* G=P㭩5y��hK�Es����;�\u��T�U�Y�����Ҳҏ�K���OnR�x.>���B��={K@������M
�w����I1�z"�}wM|����2R��N�I�7n��Yɽ��#��w��7Bs���͡Nn��m�5,wŎ�1qaʦ�u��<�9��j��)���@l�"�ޤ�9Z|w�#�*����`��Ȩ�����niei�diP7�u����#��R�݉m�!'�3�V,�6ܛ��o�������%�t�t�Gvjj	*70\�,k2@���DNcvo�YY����i\�\/�Υ�X��tos�-W����u�o�i5�b닕�#v�R���qLx�Gr2e�K�}O��X��s�fS��P�i�XN�D�xF�����<wӼ��n�s镉��"i��#{~\ç�����OWv{]�4/"�U6ET~�YQ��k�h"�*6u�ʚ���W�[M�N���~G�<q���%�=<��OsPC�3�
�WaJ�Ko=�[��s���.��F����� �$�d6:�)t��vRlN2��i�p�n�EJ�vi!Xup=�Ӭ&���Wn�Js(uzQ�{�&�ҽ�ixb��M��{�{�������W9h�a��^}:�!	��-`r^Z�qO�Ť+��$)Bʢk���#2�z�ˠz�t���}b.
���)�W�	��	�k0�-����$^E�P�ڮ못�kc�^bDb�r��k}��|�i���V�c��]2p������{��K�N���M�/�����c��ia|m\L���̊f���o��#��ft�'p���gX�K��)U[,��t�A历�L�y��R�*�
;�-��h��=خ�z��!�0PL��}�\8����Q�,V��\%7)��gŊ��q�Rx]=j#��^wT=wH0�G����Uш+
�W�_K��z�{ܩC�v.P��.uo*{��Q�]����{rpAL�"7�2$�����:�b�L�_vmȼ���:/4���t=���cs1��s'�N�]�Br���h,����j-#Գ��Ib�K�z�s~��^�+���?i��3��e�N|a�M��r�K�&`�@�>�����(�YMȷ�j���sz���G��O����y�m�`kl1~d8��t�7[�5�<��|+�lw#�����3�|��u���!��sR�N�g�誜ޫ�U��{��(��^��=�ϭ�s�O2�=R�����	�pR��[���q��օ�Z� �vS�r_��J��o��d��Zw�L��FC�P�(x������z��M�z.p���%W�r��[bI��@أ�����6�d�����@���˽��)U����ݐ3��Re�����Ʃ!��:��Y<H�Ǟ��[���3��V/۝r%�Eq�)��cH�b�<��a��*���h��W�Y�����U�̆gd��L�d��1s�.E��}mҷ��#S7�]92�O��!A0�s~����J�*���� ��|�`�յ4)�����`���#�Td�z��-:�XH��m.�^#4���
++���Ls�kjm�.�)ʿk-޻
����F�Bv'8���mՍ�&H�5������i�3�5�,�F�{v.k"�����ٍ!����Ku�O��齩��]y�M=�
㵩F}3N�x���5
d(�����}n//�Ο�>��rϕ����-������@���a�G�K�0�/O@30�+��ʊ��Т������\�iؾ��[#S�J;�j�Mt&[�����h��f��Z�G�7� u_��(3��֑�m���s/�:�W��
������y�QU�]y��Qю@(K�>+�s��dx�/��,9�:�M������i�9�ш�cT�����.\D�R�άկ�LP�nD2�ڝ��W�Wf�[[һa��Ò-*�μ��v_35/�;����ԜdPj�Q�o��1$l����jg���T��71V��,�i�$�b���; �k���.uRw�ۢ�X�c�ַ�?B�SA'z�N͜1�9.�wN���HN�^v�	i�����*�r�H�;M�^\{B�,o.�&��&��g����F�ۚ��W�8PL����P���f<X+UnE�r�'N&(cB��U���[�p �M�d�g�+�q���pBŏy/�\��J���ǌ)�/H���.]�X���9�X���ջ6hy��ok�BUe�]/x�l
W�FC�v��=�T��Ǚ0&t1�0��ؾQ;�LzF�e\,�J�E���T���C@R����m���X��y;pl����OU�O�8����qz��/<ʁN�ؿ7�::0dr;-`)��U�>U���%ɳ�/v��z�
���u�i����6K��׭ˆ�t�V61%J)fס��G!bP���+J�J�g!��\W��2�@���-�n��r���mӏ%-N��Xs��ŋ�٩u*���i�q0}CO�C
x�C}j�&;7݄'5o�����r�I��١��h��cb�,ڸf�05*�y_�B�>��+��m��L�	�ȡ��N���N��vN��1/fc��ie�� 8�����,BD�Ӆ�T$ͱc ���7�(��q�%�0�jI�(�h�k�я�Pt?9q���L����?�??p"j�k�+���-���ڰe�Y��pý�U��-q���Vvo�����]��&���E�RBnf��E�n��Ĵ����q�d�Ν&�;jԴ�)�}]������� ��J��Bxd.&�S����]�����2���N��4�͖s�]�P,.1���*ջ��a�nϬ'U��Ը
D�V_
��>@{G�s�����~����ں<�g�ĵH�>xF>���Œ��9�: ��^�<�o^�!o����Eec�i�����x����hڇL޳1N[�n7Ew#7P���[�@�cN4�
3^O��qM�!Y0Xc�?)1�.�\��5�v��O���n��b[n�)�쉤��j���5��T�����N@7j�ݏL�;�yY��{�Vk�f�*�=F��-a!-���襾_Z+K'~�<�^�h�> ��$�,���2�3u����˶�:tGC�vW��n�M�qKME��(48�'q�,[ofk���Rmt\c�D��q1�f���$�7 ]LC�N9�����t�9C�i���*G�Ny�@w�Y�ty~U�V�==m`}��F:|�lIr�=��T� �� �`�D��2�R�m��J��IE���V��T�/ʄ�δ����VLSL4Ȇ����	�Br�"�lt`���h��r[θ��lk���#�2;Km�*�Lrg5�,Fh�wrt����s��D'V�T����v��Jig���ȯp�s@�0��+�*�d�S��l�6��PUpdH��/����9Qr�T�#9y��:�VF5�QG�R#�A��c��3��4��eY@7�Y����'��c��n�b|�u�g�S#�J73�'��C�2�*ƌTc��1���Ps�B���t�����z��"��
�R�&�7k\����\U�q}�Wwy;�F�x2���Z�� J���bwr��m��3�.�厊�2��z�*V�0}������X�Z΅I8V�`)�'`:�'�eC���У�X���E�Sqt�o�^PV�:)Ԯ�dgn�=7j35`�f#Є�cYWF O�
�P�}.,���`�J3�#Y�w���]���~u���6 ��N�2%WR�K�V���*��Bُ�!Ѡ�^�\N�X�չ��1ܑ�tm��)�n��T���T=R��2�EkWJ��,��Wֶ-�wCإ�<�Bܕ�Źq�9*�a��ˈ����}=�����Pv����B�7��T��9x�v�="ur�%U�.C����D��^^D]�ތ˷������d�콒�{S�K�[���b��[���s}�J��z��� M�xI�96h�4�Ul�Q�6�ވG�v�T���n��^��T��!6@zt�#"ӳ���[��N9���f;ͪna5��C�m��ʜ�3}F��@�7��=�1��5����PW�+W#���=>�Ԅ>�p�����t����k�-Rz���5f�R�}��F	jfAYU�Un�lXδ-�Ԩ�\S���k"��}����o����C9Q�C�WFP�$�ql�L-e���()��Zf�t�����1(�m�ފ����eӈy���'X�����(O��("me�Xa�L���O*����]����'���K`��\�d�qbY��%us;u�A_:�X�?n��51�;F�G�۰��!� \\'�i��q�.�NU�-�}aB���%��U�;J*����Jr2tr���n�螌�@�V=D	�TM.��W�89r�J�%^�jdu��R���:6����EJθ��D遲������C�
=�Μ//�����gO����aqkb��E�Ǒ8��+g���`�g뒰A� �O@���"AݗJ.,'�E��5(@��'2�Y���jw�*Ώ4`�]K���^S��,�����-RV�R1},YN�G�����l��|n��Ƕ=����U"_,�X���	��b�o�6�9�ir�k;o�CN�ϳm�v7�-��W����cZ6��Uю(L��Ŷ����rkY9�G-�Q�AS__S�~O��yq�B�:��e�|�R<�DU�E����RaRBn��w[AC� z��QkN��;<�_	��� '���c�Cq:r^,�,�Dg����ө#Q��a��2է)L@;8�\V�����.\9�xr5�>Q�`�qs����s�O��7}�c�'o�m��O:���#��s��ɗ�����b6�5'uv�[1۬XkWn�aH%���c�-�>�5����N��������a2�`�Aq�͝C/8Z�6�8�/L����Xg�$�r*�����n�U��9؂ߗ���uq�{p�L���x�-N-;���ڬ�e���L���"tG���c ���]��ƹ������^gk�ܱs�0��Cl��r;%z��TzV%xSt2逼+�f3��2��Kk��f�Q�`�l�M�p�/ڈ�/P)��!�#cak#���ğ:^��}͋������	����٧"̸T;(Y���:i�����nD<T25%J)o��T�����(���Y�q�ngʻ��:�u�N15��K���Em��ˊu-��ٽCC�!�hK��۱�p��w�l��y�wjr�6���rKswsq��)�}˨s;+��Q���Wj�]-�*���;� ��R�r鼟�ћ�yC)��2c��-�kx5��VS�м��-���*Q�\�/�u0J#R���1��
E�4�S5���uh�	���껧�ji�.`[�-	@���&�u�u�Z��3�ɏ��}|ƺ�ۗy�PV�Ʃ�PM�En��P��ou��Oy_���TFuC���(�^9e�ueَIut��P��s�b�56ۣ��KJ�3�Oa˃2ZG��̂�t��T�C��]�6гY�a.¹�R[���kuܴ��ܳ��<�p��g�;|c�Z��w���Xs���ev�EvY��L���JEY��k��uh�ܭufZh������㻛���m����9A��CNLM�8^Ώ�O;�> ��ŽZ��Z���������r��fm�	ԕ���t��:�ı$�Ū㆑�Բ�Y�}���!�;�E)3QRތLm�հ�W�P��zZ4:�\���K��jݡi4��Ҳ��X)i{�rk͌}�on���|�P�I�x��S�^e����7eک�_]��ve�&��X���z��#�������s�FG�;�]b�Oxo�j��Nwc��0�r̋fm�`['��͒�[|~|�1Da�	M��,�Wu�+�x��2�\m]L�	n��X�r���6WZ2�}��pN��6�b�m��=�rس ������Bo-�����c?��m�O�9���w
W9���E]f�>�d�s3V���� أ���ܻ%mZ���[X6\3�D(i%2W)9v�Kŝ��v�e�����a�u���+^Ro,��ʲn� {x5�x�S��o����c3���	��]>}���fNs���JHՊ+���]���������L$ב��l[�Ӈ�����bu�Z������s�w�!�����ljCB9˶�����IvI)�{`9��z�
i������Q���x� ����$esS�����u�$�g=rY��^�ݐ��V{�~'�eX����+v�v
P�x�o�&�S�� "��J��*�f�������(6�U�ޏ�n��h�]������*;aސkQt%){`��X�S�^�n����o2���oy�b=q�� ��,�k�u3M��sw3���a<&
�Ν���\��&$hۄ7G
���1/����tvb���j���-�{#V#ܧZ��Ulz��;�H��u��θ����p֏	Z�|����˻�Vo�.+#��wն\3M��=�`u��̧ϗ6��+A�ߋk�+s�^d�Y�w	"��Kj�
��w�� iY���l���5�����7z�Tk��7�-7n�����&����ʈ��)J �*)��%,��&����h2���$�(���2rrH�JC'"�rr@�"�&
B��$�i�j�L�2���)+ 2 �2�%�(r!2� �2V�2���@��ƀ�rL���2"G	b2C#$���'#"��c#	L!�r�!�,�3���&��p���#02
\�rJ\�)³2ZZG�3��r!�2ik r2�i�2����rZ22h�����C$�Z2B?#���Z�2�q�~~���5
*��������1�6R;gC�'D�ʵζ3)���p�k�y�f]�'	���#�{�^�)��x-��o��f��Cզ�m[	D��A�=�ˉ����vݸ��R��U�;W�ȳy4�2r��`���"Xs�D E�蘡���v�վ�r�d9}�C�uq��̢Nr��$�#��j�p�<�`�D(��݅c}��dv����܉D��8���K�Y�����V-��MH��6�Q��qu"�8^���K� ��ܝ-��Y'T��b�_���]��mȨ/N§n���nJ�ȭ���'B��	GL�crk]��[���D)�(Ӛ]��J鎗Ҽ�P.�;��a�n��>r�E���BW'<�����ެ��>������4�k�����N��v�9��W,��r��ʨ
㖫}���5v ���i�)xm8�h��b@s[NP���#�:g\�"�@��f=%FJ��ђ�C�VCΓ�2	�B|N��h�!Y7��]�Z�Sx��l�n�޺��1÷����M�P��n�+��쉤��j����pdU v9���9x����iZ���bۼ�������5X���ʹ]���Դ��K%PEY�p=~q�/EE��gn�c�ȼ}��h���a�%��NS7���;;AW��X��F�lՔ���������\�VgT����T�:y+�g^h�&0��N��#��Lzπ��PÜkh1b[��tz�u�2hq��0J��`-��rDX{��9yMn��ZlWU#|\<*��rp�C��o��ϰ�
[j����|%����M���t�$+������[&6�w�d�!���b��"��v���}�7y4�q�ja/��w�n&�*'���IS^8i��;�dӅ��{&��ʊrh]F���a�v�1�"�+ k]��
�HT%x��+�(��qGnq�T&﮼/7���.��P�#��;;}]xN4�X	{��Z�VG5�}�e�[���PB�輄 {]�o��w����_3|��F�(�5��A�i��bFb2'�q���d�����������B��Bmˁ]����Z8�7�=<d?�Q�5WR�D��gf{�_].\�⮖kY{�QL@��\�L��vsC��L�+�K�c���==U�!@$n��gOE	+�=lZv,�����L��wU�҆�]}
0%�۝������E���=�~uY�k�y���M[sy���<��
,e\8xiC:N����T�Zj�^��)�/�q���v�K��}}�za��z�Q�������2i^΂mo|�q�i[:�9��3��и΂�7��'P��:}ۦN�}ٜ򘷪Q��oK�X�ރo��[��d{��J� >1^j��vS�tHW�g��9C�>ع m0*�Dpr}�˙�Ӝ����u��~rpA�t���dI@�&N�,ݫ��:Ż��|�s��֩G��Kg�����빊s��rP��nH��_�G�U���E�ॴ�����._�twy��s��3([�`wS�s�|a��L7<2[0c V��<���ڈ���d9{ra�O�߾͛��1��|�:
�۶�05��C�nOM�繛�:��W7f��$�Oئ:��FC�~ň�/�q_���N�6|~���v�Ct�E�Z�Z�"�T��k�g���.�~�ΡK�]x�j���EP�N63�
q�%@>�F��C��|��3��C9�{��@�^�H���|T�p���^0��e���Gnb�hl��v�7�qUe
�|�������ӷ��i���V׆�J�����h�QȌ�'�J*���-�{���&ps�(#`�o=�B�<ٸ�N,K#�Td�z��r�]j��,�V��'�ו��\�K,7)e���|��a�+���*V�+b7I	j�\E
�<B��nJ�6�3ni�<��)e�t˭���(h��:݌��M_W ���V�E�B�7�B�:(j}i��38<�+��]K.e�3�pAm�}n$w*٣4��R�c���b8p�vu=�J\:E9W�P����,�b�%��U�ٷ�3�'��؜��X�;�ʉa���4�d���4�Pc��u�G���P~<F��b{����W�{Y�����1��g��e�=b�C�
=co���/�������l!��S;����<U�e���\�;��ǙY�_OT��A� ���LÔ�U
��EŁ��(s�l�J�{<��9r3êu�HP�j���o��k���(a3O�"yC�@��������ی�he���C��Ҽ9���!A�:����h���@>B\I�@�*4���ˑ2^_i����\)J]L96���om9���Ӫ%�o��A����e#o&��sy�WK{<�������q��O]�Da}�K��X�M�a��3R�����b6����RŭZ��OV7$�A,1J*+�2!����߯���s�5=�Ǩz��wF"�9���(�k�V�����X}R��k��=侱rs�>��͎���S�`]X�{L>�#$�(2��I���w��qXcJ��t%>p}�Ϸ97tS�2�])Y��WcW�oOvvJ\�����W`c���Wt�vvL��h�T��ky��(g|��pͶt]�m�pU~��A�����Z�9Ժ:taAp��Em	_u�y�Y/�f�g����P���Ϯ��Z6)����qjn`8u�r����B����hs�0��C��tk��sF�Κ����xxSt2��u׭�B�u<4�G~�w�Q1fX2��M�p�
,j"��e@�t�v}�.Z~ʘ!X��ӻj�wz�Ohr�a��E5�/�zd�@`Ơ�m\Q����Z��kyZ�X��WoV±�ژ���%�UQ��L����e@��B�۷D�*ƱB�P��i��o�g5�=|~��[���W�;�_R	�ԃ�;��Qew��<��*N�t��ou�-�H��SC����އ3cF٠���t�x'�����ϥ�2_<�0;��ܬ�UF+#���W�M�ʅL�s�V��/�A�ߍ�'�n���j�^�N�è�sS�zX:}��S�\qȨ�}]����7[
���iU�6�&�q�(q��krU]f�{�(bf:\u��l�-л.������h�V��'r~ϻ��(��
"��cy׬azn^-��M2\�P$�Wʥ��b��6$"��܃I��1�SV���������iZwN��ޛ���������\�����{}ß%���3h;�S�n�����m�:��p�v�Q�Wb$f���ۢ��V���3�Zk�s�D ��Pz���Z�GU^Wϒ�D1�����
�5�ˀ�S���%�Z�ڸ�l�i:���"xYQ���P��m�#�:f���z�R7j��x��WL�S�\�nN5�t(�'�4N)�.B�q�B�=۶Dp��mE1t���U}��r�Ȉ���n��\bf�jƗf���T���7�\���_EuŨC�rH��n�d^J�r,f����\�3��@<ϰ��d���������½��x_�mtЛR��aI��#/}�"<�ňu�^u��l�8��QcP0j��gW_%Wۚq��~`�>�=p���;@ۿU�Bn.�!�9�j ;1&p,�s9�5b��#Ij���D��|F	0D�n^
;��ۅ:|��#N\\7a*R��ڌ~�ꑞ�:��¯��a�3�z}�0�r+DҚA�@��
�J�B-О��k�i�r�ʦ�,�9'�W��ك"��-/rּ�w+!�|E���/x���m�oU0�Eh����dVm@����Xci��6���9t%�`n�j>��oV���Y�-��qF\5��p����'Y���m�WJ2����U�6ܭ�iG�|��D�ݪ���rihr�[z���ƹ����sVb����/�O"�Z陋4K����ɉ�w)\�H�H�KM�^�F�(�`��z�u�K���Q�3�${��Z�v�O����f����tc��-�	�6�@�vScQ�"�n
�o�����֢��>	����li�F[�Q� lX'��Ǣk3m���*s��T6�2�^�Yg6�oa����|��L�fZ��j�$yq@�9/��^��o�n/x:�}��{Ty\L�N�Y\�Yd�����;������b<��X��y��!_���j���+��'o��}�T�o�h��� ��y���g��H2$�v���+��MDib���̮��2&'\��EW�Z2.��`T�� �T����Z���"�^D��s�j��g�Ε;�e�$A�"���u8�9�>0�&�b�(l�0c V����0.F��@����"[(�:Nl׳�n��l۶�� �p-�E���u�8�r��Ǝ�6�(�*�_Ld���+E�C1XؿnۿX�(C�5�C�઼�BQ���oDǗ��_J��)vg%��=��k_P��D��a��OR�t�)�K'>I�����t;u�{AK- �zX,nݾb�f˫ϕ,����T���Cv�����!6��_�O,Λ��X���8�j$f$�7�xZ^�WA:�����a,�u
���4ddUn[�ԅ8�e-�x����=#�t+s�(�ض�������9��� �&וA���	���/w�F��"�;���aȅ8:u�W��6]oz�;@N�M)���'�C�(WZ��r����8�^�?N�`0{�;A߇i��l8n�hSg M�@��84=���6h��X�&��y+���=M���'�å�u�ՑB=�8Z�ۡ���ҍsU�z�ϙ�����Ҹ�
����!��X��"2\t���w<�ܸ���L���ǬV�F&W�c��yy�^��Pá�=\v4âB������v��֫᳓�6���7���J��N��a����h�.=r^A� �O@>.��[B](�DUI�P�✲3;ۯz8Əo*��Z7������Vȡh�xOGz3�×�^c��uuu�J{RF��ޑLl�
-p=Ns!E�#�Ӯ�����5��/'`�?>��g`����c��͗)�=�Z�]×��Zu#�:�Qh"��.�a�'Ʋ�,��I[KE�4�q���ն�c��P��TˡR�uY�H�9컰�����ط�����k�N�A�	-�z���2ƿ�� ��8�j�A��np��w�eY�<�R5�������KS~�L)��min{f ����ߪ��Y.̓$��t���2�qmG+����|>�C�-ȉ�p��)6�K:�=c��qz�Ծ��kmM��˺�Zlv�fi�9���)[O�X�EzE�꧟ߗ*�ݧ�ۃ�@�GQg��s�
4��(��Э2��MoD�L9�B����5��'���i��t;赸ߍm��4����`
MСn��+9���`v1*��X��[�ض�QZY{Zl���H��^�ʦ�q�k�*��t:+Yg�MEo� pdi���3�<�P�B��;��WR��3�:+��]#�F��%g*����O��o�M�r�?eLʝ~ѣ���c5lQ��桨_D�5�1\E4�X2�4�!)^�4�瓯:�϶�׫b;q���-�����T��mz$�����t�~,���
[N�8��,����Q{Ԝ�$|Jg�z�����;�N��hi�nx�CmWD�c ��vԮcr�+}W�Ø�]ce�r����z�?R	]��Y�h��R�5�G�����3���7)��Yj��ՙM=o)�-dC�au���Om4���:r_S���`:�b��y)^�����A"s7�'t6���m��	�+��Er?��f;q��u�u:.��1r�2")�g�:�]�K���Y+*�����C�Z�ko5�Vm�7��V��]u=�t�Ϧ�eB�jf:���(�e�ԋ����[x.�{n��/V�ֽP�W��P�4x���\��EA|zS�kr���yQ�n�e���\���i�Y@
""�aߨ�Mt.��t�_���*Հ���U�>F�.;}�0Sܹ�Ů��bʖ�`���@Pc��1�EY�e�r-p����,�Z�����ŉ:3T-K�n�D�Iפ��9}�)E#!@+hL6��07�����]9)��i�i��g�&�d<�s�Fk�	��h�!Y7I���p��tT�WX�m%+����upo۴��DD&�u1^l�"�5�V�g��q�M��V����z��([.��wՑ�✎�5����H��+å�������յOt��n�1R�K\3"���n�@�e��p/r����Є>��7Kf�8��Q��}5����-x�wPe���<U��*��:vގ7EY8�Q:[��[G���78�	[�ꇻ�i�Yk��Cz�Q2v�C^ưk�$�P8%�r�L�\m��X^��]'�ܩOz!��u�hZ�����#����q��f]w4�i�ݦ��=��Yf���.]|(Zۜ����?��<��q�؈�߀`���\u���6y��	�e�1hM��n��-f� F�A1a}f�)���B��o�e�����R/i� �}�Ib直�+�Ei��ie��"�c躘7]{$�|5�I�r\�F���6)_���7�d�r�U���n+/_��z��E�K&bO8v�J��j۾4�*�,��M�}S�v;�Qh�`��Q�ɷ��M�m��vtś4_i<�z(ih��
���V!�cvi����w.c�
�xoU���+����PeX��*�vX���#>B(��opfCq�D��3���1���Mũ�����[rL�~&������Ma;�B�q��3%�S�T�<�J]sjn��ν�X���ܼuk&�۲qe��ǐY�r3Y#cF��^�Ў�V�ED
ٴ޶�u(�}^��'��z�i��m�!��{[2�P��Ӻ[�g]�Ǳ;�w=�֓��^�y�]%Z�;��+];�uϥ�\��3t ��>��q��t��^vn�I%]��W�fa�)��쒣?K&1w؆�2LU�veڎ7 ��F��i�c�Tt�:�@�|��7x��ff�.��맔�1�U�-�M�苒S��l�u>F����E�{����sT��]��94De��_b�:佣�d��Og6�*������7Yz4!"S��j2	}�8�;˜�`RMȜ��dC������<���բ�lG��nͭ�8�X�pܡHMJ�S}N���A�5����"܃�ʱ�h] �U���κ�Ρ�Ն�e\����|
Tѹ�5;\���*�#�����J>�����z�Y�{�}�������S���ν����z�sZ)\�ǔ���G���c���6ĝ�tu�shl5d4���������2�^���Wu�mc]��{�Q�ܭ��WՄN�y9���v���[�TRe#�]N�)�]�
]R�TpB+r!*�qb�W���l��F����������c�/��vH�V�Os$�RvD�d5{l	N�����ͽ�7��V"j�[H�PD�;�@ŝ�������W]v:x3!�d�uwȕ�u��T�[���r�����2�ݨ�-1l�W�Q��+I髬b'�`�֡�3��|�ry��T.{p���.(q���z+3KO��t�y�q�d��[G	��zb3�r���[�$����؜veŝQ��r����4��]�ܷ �%i}���[cy��V�R�t�w�枋YC,�0j�c�+6��n˱��hV��;�8dn�R=�p�z�U�ֳ~��f������Kf
����|�kYך��{�I�E&�,�rI��3�lĤ*�2
V�2��r�$���)�irJ�ʖ�3�r���r���$ɣ	2
��&���%ɣ ��Jr�"��$

����
���@�H�
��$i�&��%�� )�� (h(������2)
��R����2�
�L��(B���Zl�)(��h�)L��P����1��*�3)("�����22*\�Z�j���2ʔ

*&��"����2\��)�L � )i���*
�����2��I�hJR����j�JB���#3� 
Z�����"����gv��������ݜ��$��ܢ�8��Ǌ��٬��2�t�|UJ��cZs�-ܰ�ky���]�w]K{����o۱U��+WP3��"�0�Ex�V����6��/��s�u11�.!J�qHP}1��c/[=\����sa�f�TV����!n^���+�6�F	����Y����4�s�<ۥ�*S�R�`bg���d	!���4���a�����y@��f�ꯖ���h��Ժa���xo�z�G��d�4GW��S��5�pW%�w�;ؔ=��a�9��z�	�vk_�����5���7>��z����	��u�W�2�f�rs���0=Ы5gNd|�kk�[�r�C����(J?��ǫ�u����;�K��r>��;���0���rzy��Jn��i�>��\�?f�'�e���i�]O���g����)�/ksU�߽D@�꜃����!�?T;�Oc�Ju=k���I�Hu��nO�����ߟi��䚊;�5�n��>��{���ܺ��y���r��UXF�]��J��2=��k�'�Ԝ�'P{Qk�2~��oz���2w��:�Z�n��o�$���掤���������A�O}sK�|�����sa�%�.Bs�סꎿ��5B�d�m��t
� =����I�O�u|�A���L���V�������=�#�x4j������2�Pt~םt�N{�d�����x<�F���^#�R�N�uEVl}��g�Ly��A��3�{�p���_}���2��`uI�X�����4r;��u'֬�"�������O����c��'��X�#!4u�{~� (����q�Y!_UN��ך��]o�������{�ǒ�k���h�O�˒���.�&O���ts�'��BP�����S�n�y��`�&���NF�)���
ϒdP�u��<�#�G������G�/�z�=��qj3�#��+ ���kh�Ŵ�`�1�WkW�f:��U]�ӽ]:�8U��w��V��ND�.�Ȳ۰6��s�� %���,�wM4
��z�]
�p�jl�XÂ�Uܦ</~�3;����%�n�mn����]����Q��x{	i���z��/�Жb~�Q�=֟$�FA������9.��kTP}]H~�zA��y�4{�h��=�zޟ���2y'3@UP��{�5�V��:DG�R<&<|���<� �ڗ{���﷟��⎤�F�5;��j�ȮoԿ� ���9P��}��4��P�}�]C�2sQ����I�29=?sA˸uK��i��R�j��<4x� 
�1��L���0����}G}o�{����=����y����l�x��~�2��R{�����:�����P�����	Hw�5�+�2�x���;����ds���%<�����%Ȥ3g<����O|�>��n����y��{��웃Q�{�7�>K��;ϴ��d�1��%�
=�2_֡)��=���^Z���&��&\����w	O��ߞw��xP����^�@�L���L�B������{ל���0L�ʞ<溞I�j�O5���O�dPw�����w^��%�&�ټ����ё����G%ԝoE�r��x����=�>��xLxtxLz� ������_\��`��q\m��N��p!��@��R@UP�=���J��W9����=~滞Gr{>ơ��Z
{����.��BR��i�
9�.�:u�4�>�R��~���2{�y��;c�*z _ڶ�ӽZ/3u���#�#�E��_��������0��=���h��˒�\�O����sx�GP�<9�6�������ԟ��X=Gѫ�����uj�����{Α<������1#)m�j��z!G�G@p̺�7����voC���^���ȥ�<Ӑr�' �<�b]c�y�>�<�p�I����X�\��\��=��P�}����z��>��y����ӺG`��h�c�xǇG������S����_5�	Y!��S�t�49�	�}u���:�d�5!߾�s��O$ȣ��'$��z|�:����s���&@}��Y�V�_6j0��a��O�lL\�|x�TPy[������2u&�p���<�.��'"� ����.�*�z�P�9=~�7�{&o˧�����NOq�?>�������98+���Nڟ�o�y���z<�e�!i;	j61��9pȅ�H1<�9*;��d@������FdlՉ�E���D�<h�S{X��	�s����ŰEȳ�ˬ1"%b�}�����컽d��Ҳy���s�@�<��Yo)���<=�)���as�����(��]A�jB^a��i:�{��ԝ�ޞGP�N����w	I�k���|��d�\�
_�I�ZM�ur^���.BV�;�k����s����=�]�~/W3���>�Ǧ�{�@�������_�滄����ٟi<�P���'�RV��zy����w�`~37ѨJ7�U�d2M����/�����.��]
�x�����9漺�]y�|7��G�;�_����4�K�G���/���B�����~�~�$Խ�~�� U&�0��A�U>����X�+~�G's"��ډ������r~�S���%'$��^h>��K�N�5ͧQO�dޘjaˑ����p}]�o7����O\�A��&I����:���-`�]��G%1�"" j3>�]���Λ��j�*�DP�9��5�>�<�:7��'�jOg��n'$�5�4;����~m�G �'��wmri�=�Qߟhr7 ���?擸JN�����?@�|�,3����>��xnH���<9��n��rdQO��g�j�y�����u�����w&I��w�4r:��p���upd%{RW �;�� �5'=���;�-�w��w�y��k���:�Bp��������s��r�\�p��ܞE�O���_b����oQ�Z�Pd;�#�{���$ܙn�}�r2�G�>�������"6���}����z�K�9�p�?Tu�k�9k���4�Pu>I�ԝ�sI��|�S����)2O5�A�5	ob�QO�d����d�ˑ�7������ݥP��f�-��߀�Pd�9ͯ���:��惩�NE�O�s]O��WG��r�(:�:�n��L����ԝϱ�:���Ρ)�MF�ȡ�JN✃��5.��.
����wz��}�D{`(����� ���|��	I׿��uK�P�{�%�)yj��rn�ˑ��i:�}�!��h7}/����C�����Xx{�nN�ְ<���-~?{�F~�끻�[Z�؇���jv�o���e|���n�W+�K1��P�v��Q�s���W�}��$�n(s���Iى�p�h���C�Z�FG%ӷm.���:)��ć*��f�$�}ԥ�H�+-L�t���g	��ʚ^�ײe~��=�製�ڷ-�� (�w�Z�q�Bfb�%}G�x��:�Iѽs�&�!�5޿h��P��r;���JC�#���2�<����?I�����1�\��תּb��(>So�0"ǽP`��<a��A��k|�2O�{j�w������wu/5���J��w��A�s��h�}Pd�'Ѩ�u���<�S���4�%''����y߾k������^�p�!��� �<�ã�"�$���4�GP}]G����� ���C!����/7�	�j�MN��-`��4���
���C�	G��h:�]��3���9޿g>�:�G�Uq�y{7]񏇦<z��P>�����)�O���w��%�'��?G�jL�^b�Ӹ�>��<��Pe�X^b��vk
MG%�}�:�n�
^������5��G��}e�r�ϟF�{�#���w�
�^K�Խ�{�p�5��~9�Y�d�I�a��FF�)�>��P����vI^���hK�����/؛���ԝ���P��s\�����# ��r�������zc��(�-c���my��2��4~��=�z����PQ�}�v��!�~�#��\�}kX&I�ts�=^���7!�3S�r�^����P���u����}ٽ��5�{�y�}~�S�}o��ܟT<��﮴%=O�jz�4���o����=��5��to�'$�Sԙw�4��P{\��wͯpP{<惫�	����G�{�h�	�Wq8�C����~߿��u��M�Rn-`}?��j���	�Z���jOd�p�ru?�Rto�~��)�N�u͝A�'{����r>�S��iw�.M=��� \ 	��}v�/����Q�u��p�|���
+�>�u'Q�Z��kG �KXPo�kr}&@j�ٻ%ȧ�r(h�%�j���r5���ӿpL��39�G#P�{����7_+�uw�[��Ne~���aMe/����CvI^ǿa�K���u���N�!�jޗs�C�����:��Pl��' �%�߸R���2��u����=����K���P<"�0��n�B�֍�[;��_�t�}l��8oiitJ�d��kFU��gƷE<t�)�7t��{2��62C�ٵ�[��%\��%ؤ��n�)I��]���J��U���2��˂�`h�2�B%�O�&*%t�#V o����n���8�*�4C�Rz����{�{�T��qim�w{��q�G��3�Re�s�ߜӹԹu/5�a�obP�o�h>����1?sZM����ܝ{�BS��u��ME	N�0��~��5N�5�'$�S���$�	����~Ŧor?( T	�w\��>�PPl�v=]�d;�����\��z��2w'"�}� �u.I�9�uP��%��i�=O�Ru'g����:�Ƨ�p���Jz�K~��!��h٫����6�� \ �	�����9A���w��N��G$��d=��͆Ob��y��rdr^Z���O ��vk�NZ�Rd��:��ˑN���5�仍Ef���P�����٤> l8 ����Ju�	�u�����j�z��>Z��ȧR�,��ֵ�	w�ty�����bj2cW��HS�C�#�i:����`n�O�jC>���a~��y�EUoӰ���%�W�g�=����?4���M�;�`��2M~·	C�;ތ���Jdto�n������&��r�^����(J����꜃����.��A�ɺ�����q�{��]��ܟgwV�߂�`xDz���_�dyI�BWA�h>��� �0s�O�j)����2I登#���6�V�2����%湥��O$�ܟG�~�} ��\�y�;�z|>w����VX��D@�@>>�O-I��~掾�2N瑯�ZO���Jzu��Oc�<�"��`j_' �y�
���Z7��p� ��(5=}��zw���rdr^�~�]���>QP!����[ݝ�'��&�)s{_����^�:��K�O �y�;���/#�u�(z����sI���$�Z���X>GѨξѹ�mC�d]�hMHe��¿A��x<���25�3��;c��+T��D������gP��˾b�(J���I���|Ӿ��^o�y�kp�B}�vy�R��9<��Jo����|��	�4i=�/%��n{�g�כ�}�w�{ݿǟ�Ӌ��.Z�鵅	@q�({��?C��GX������~�=��)��k���I�Ht{�[��2=��5vy����NI����5�n �=�#���0 ����K�f��UEf5J3�sn���:�=�p9�ps��]g+vĸ��G����MK�˝n�����V⭮��� �o���>���X��k%�X7�M+��&GX��B�gJ ��L5�+�]��\lMJ,����r��Ε^�~������ӷ��:�� lLlx	������}��sI��MI�:�o�E�`��^��@UP�N�1hu<�&��~��&����͝���5	_�����A�O}sK�|�����ɉ�>�p}�L%��'�6�)��>�5>F��їy����X���05��#rxa[��2C�3
_-I����.E?G�����4d%���y�K��&O~~��£=R(��4����AaG��� �y��2~����3|ѨJC�/����	{����w���MFA���9�S����vK�BQ�����O���u��/7��v���22?{}��J�o�wu��_!���=�@���m}�	I�����y/-{�~��I��r_��~]�L��˨��=�
��`j�r����0L�u_E'#P���}���2(z��3OԻ�c���M�.���<&�{�Y�%��I��z��2Q�yߚ܎K�}��(>�.�:}��Pd�^k��s@u'$��;����A��9�j��Pg��	�w:�?{����r���(�ϟ_�	�>H�ܜ�F�:����5�dW{�5/��6����Kx�>��m=��jw~����?����sZ)7&G'�`r�A���i��R�jNI���}�����s>b���Uq��Ll{�#�ϼ`(�A�cF�(w<��/s���u����G#S��]O�|�_�h�P��}�[���!-翱z���159�����T���{w�o/<��s/wq��Ȥ9�������Qߟh�����N�L��2]�ckK�o�h�Z��zǸ7��_b~:�ܟ�˒�����)�._�u��XP�{�}�ZΔN<��:���������9�_�L��<�ny'��J��n|�S�L�O���O$���}ǨK�MA�yE?I��#g�(ur9.���:����=��=���������U`�
+㘢�3�$+7��w&O9�{Ob��d�>}���
�GA��BP�?Z�y��u�	�w�5��;���5��ORy�peՐ��9��Q�7	w�Ѭi��ǁ�{��7�-Yk�#O˱Tfq�~Q�����ٚvwn7�q,�)nw�D�j��p]b��dH�Z�V�VV��F�A�1�֞
u�M���$��¢gF8�2/�^���YD�Ԯs�(F��(���0�1j��ʄ�
�Xf�,����=��ճ�����ơ�����u�(�ܙι��}�$�_����Z���}���;��.E�<���@Q\���'#�J���a�x��{�y�4u'�>�Q�j�t�P<`��p�P��1�z�;��>��٬���$8�^`�I�������%?^{��=\�"���4��.I�;�:ؗX�^osI��$��4��K��h��Z��" W�3_=�S:3���c� \�z�^c����2Ԝ��:���:w�엚���5�9���>��Zϲu����n{�A��~=ր��O^sTB]�r3�y����s���s��W�"���c�������{.�9����[�ϱ7�d�M��o�	�y&Z�O�� ��δ��������P����o$�L�	���:�c�9=Ơֹ��p����ɢ
����p�u?l{c�����(J_���P{�P��w�4�M=��jN��<������c�
)2M{�/����������Ԟ�P��/��E?K�W�ח;���~�3��p�Z�{���޸
�G�
}p\��s����u'�9�GW��p��Z�C>�y��a��On������u��jM���f�!�5	F�ʡ���&A�r�O��ߞg��ϰ�+m�Ι���8����=u��xdq��~�?K�{��wr_�@s0���e害�b���}<9��a��O�^�2�_5�!�kp�9S���
{�d�p��f�s��}���;�=���A��'��xoNO�jy&GF��)=�#���p�X���6�E?I��zh�×#�u���qA�9w�-�d�}9փ��hL�����P ���}�n����~���y���uUA�aA�J�ޚܝɟbo7&O�ԟO#Q����9��05%/o����9�P���ݵɧ��MG~}���<�'�#G��@���v�K��_gI��G��j�g�؛��.�O_a����2ܝ~� /0�%�j��&��^�=�����9���G#�Jw_~�}��2(J;}�K˩@ o��?I�Q�����;{��J�������@\Oz�C6Rb��x-�̗�α���X�/j:����wS���jY���UZ��E�Σ�y�]������ �����ʅp�fI�dK�+�f�5ݽr�<1!fOlp�ӻ|�{����^w7�y����X�Rw���i�:�Q�N������r)���wZ�~g ���׸]b}&@ut��~�~�'{��Q�Z��x��2;���k������*b#�~�������ͷ������!)�����XR���w	Cʏ�����L�sO�S�}���o�}�1���FFGί#4Ms���V�:s��K�ϮMC|ˊ�fձ/<��U:�y��y����in}Ρ+(�v]�)�)��rTuίK��g`wZ�ed("�W�vU7=���̫��n�F�E~Vl���n�9��ٷ�f��H=C�
�(��lR�W�)Ձz�uHp�e@�_^F񞍲��*�/��p�����k�6
�^�P|��OƠ2�4�$!	Ll�,n�Cw�
Z�e���]j�?K��P��cc5J)i�L�To�2�vJ���Pn�c8�����&��1�3ʿb�������kH�o�|Q�ck�AH�.�
�*�8eVb��e��mF&�@���٧<�汨��w�/�� *�2ta��Qyx�]+��<7M[O��!�{ao��=��_�n���L�9#���qu"Q/u:n��{xY8�5���(��3����,8ɴ�M��ܓT�@�w�B~�8u�S��8/�bo7b�llqJ6q ��<�W�7�+��g�NE�ܟ�o ���.Y|��Ρtm��\�Fn#���/�]jQ�N��:�I���ų$뫆p��J/�wע��{������
|�#���ɚ��T)M|v��N�����:V��M��I�#�)���|��˺ra��&���bfa�GX�Y5���e@��58�P.��.V�b�k��nF��}j]��|�!
�1L�tHd�������	[Խ�^��ݠ�.Ꭳh�w�e���W,��s̝i:���9}�)E9
���4�:_Ff�\2�����`��s0\�g�&�d7`����Ҷ�h^i�S���C��sש����O��HO��8�	O�����-��@�����_X}�칋���&ɩ�9׼�n��ל�`���37��@�F�K�R,f���[A�nf)��#���.�B�/�Ӟ�Ar��Y��52X\n��R+������#/}�"<��!u�^{{���������<�{?�����	֯��UC��6,�p;��g�u0a�i�����M
c$+r4]�'�[�|~��|a�B�x�m���5W�b��M�j5b%�MM�U�S�n�Δk&/)e���s�� ��+7��(.����d؛�?*yy����'+�V�u�D�m�k���k����k���u��7}/:�Dr��Q��[�m�3����v�(����G{�:H$C}�*e����}�������1������=ԴE��u����K>Q��Un^Ԣ��RdT���7�\��u��ԡ�3��Րߒ�4����C����rUt9��O�C]��8Gp�^�y:�VF5�{vM��
��VB�Y���2D�1Ψp��g·a�Sc��e�n_���@=V�K+e�Ɲu��͡�/q�w<6	E̸�4�A=I����dL��U�ؽ��j%B�����7�Ց���C
�k�)/�O��������
�4ʽζ�`�ʀ��T�@y*��s\�n�W9u;Ls��:eE�ꬩ��TbP��Fx�p�
5���v˷zܞ��k��]]�t0�+nv.���j�L�a��T��@�1Kӊh�k+3],5����3i�jH�C�=�d�*/�p<�g���E�]~�	ֈ5ಜ9E�u�m�ѩԚS�5@a#�7�<�be�ۑ3�5�v���7N.�9ܐ&*.bn��:��j#�t�aqZk��e#�W%����h�u8�8��XL�ƀ#9Ø٭;۽��U~<���2]��J%�8a���d��P&�U����&�r,�swY`��{�jvTN�Ǣ��A��-��c����9 X�v��ݹ����|��pS`�2�d��iمV�T"�۳�YJ8�[Cl��A+H��v5c�]�@%�����L�4�N�%m�m�k ���5��^B���
�Ի�N�P]�L�T�P��6��l$֨`ɬ6�%T4�t��^��_6�e�J
�vI����&1g52��%iy&����F�q�1�I�hޕg�Txr��)sj��3�doT;2��Q��!fˊ���Ϲ��ZC��6�Zׯ3dcfSѼ�몽

:�ӫ�9�ǻ����q�Z�MM�ОR1���aᏎ�v�L��B]GLq��Ow��0�+�p��m�kK]�(fU��>�9��Gh��E�4�]�Ӫ�2l]f�g˚�)j�L��}�{H��is,CyR�ƨ�tҞ��xx�����ywJ��)�S�C*���Yژ�L=�G���\D�f��Տ�ȲW0��[l���3OV�9tl�wz�\�����1Y����㕿LW��BE�DYzn�)��:����&��7���R���)��E�UE`�/��gk�y� &���ܵp���}K-�� Ci�\�<�;۽n��@�=���vi�bwE'��Q첟\��WRl�٫�.�������z�^��\���@[��1�Pf*�[v.��Q�OU9�[���v М�)���h};$�n�vR�l���XAvgwn�9}��=N��nJ��X�=yƦ�sE�N�݋p��7	��s�j��4p�Py����(*���\����`X]�s�X_L:!�:��MV��[6��e4��C��k���u�Z���6=<���OMn����i��f��wy�,J�gI<P�N�\���۱�n
{:����h �t�u�l�{�DgU����.��[�W{@s��"�I�V;f�� 1����#]ُ�3��ή/+�C}I��3x���b�lzpm��F�h��qT]��.����4V���gb*���8�vwP��
R�%�8Q'jJ5A}��&����c90�[�9���6>o��EǏL����L9Xo7�;��U�(�\p�d�W(�"0����fQ�vi)�
ou�}ێlA�<W�.�T�E�e��t$� ��Nw��<�qgz��%T����n���rS��0).�D�Ș#�0޳�;�@��K;_^Z��1����g mZ����Y`��G�SEe�G��ᗕ9V[����i�m�`		O��ﯦٳ攘:�t3j����V��܂�,�'���І����{%��)}����dp��)���J�{�m��E��\��2�Hkw�M�MS[\/���V�}{�w��b?����z:�w;�C�6*Яo;D56<o�k�P�~�>����A�*b���((Z��F�i
�2�
F�����!*�
� ri(�(��" ���ZX�j�i��)i
(Z���!���(B�� ����@�J"�X�"
(��"$�%)2���(����(��� ���B�J*B���
J*��(2�3*���Z�(
"&R���"���
�)j����R��$�)����������)�i�Y���J�bJ(��)�%h)i�*���f
j�*���&����(h**
ir"��j��j&(j�hH��&
T�f�r"�h�*	�h""�(*r�b ��&�* ���i�I������*�*� �*����- jɬ\ȟ4(;hg��JA��͸��Ef�Mo4�-w)�u�Yq�<�wk����N`�؝�ŵ�yV���=� RΎw2�8�C'?	�1�)��<
��!E iֹʜٯfIn{�������T�+�Y�{��xpa��-��y�e�h��.Th9x��T21������ͩ���z�Y����(B|�!�r�!�U��3�J�Wy�Xľg��ȸ#"��d&rnDܣB��\2�31����:طBT�7�@mR��n�NV��Pu2UmyU��w�y!ORz��Իܥ����U�+���aN�*�p-�;-^���V�o��)�/.-�u�'N��5�r�b:e�?�00�)�(�}��{a�mFЦ��d�qs��e�f��=G9L򫡹;�*U+=��hq�ß}�iZ�ՑB8�E�++�r
�g��V+�t�\���;aWD�cb�!�X��=Z\(1�7���u��s��:�����㗁+����N���2�`�}1�z,�
z&�A�re�+I��
v�]E��>���Y������kz��˹/ Ð��kn)�ӿF�O`�b���Mp�n���Φ�j�
��ƻ����6{+Ɣ�Goww����]ruB ܉]4j'����.��YK��WV:�x*n&_>�Z��jZ�O�U��E����0��	�*,�]�XgV��NF�:]3
]�:�r[7C�ݙs_�<� D�©�
�_�$���鞅�Շ�.xi>�p�Ѫ��K�+h�u��r��vz�oR	�T�vC~��^3*(�;4qл�t_�����B�6�A�^GGOaF���nU�R�5ۂj���e0�_��:�TKW��ߵmȽ��$_N���̽WK��QTcj���?"2��MJ���a3�
�<xJO]������t����C���g���gw6�/���$�Jܨ��!���b�pB�U��k�y/��G׈��Ƴ�v.��t�f?cx�V%V�[F!�N�LShV����Ձ��Hڇ"��
F�c��#������#0�u��87}Y#�~ͫB^�`٘�n��+9���Z�s2��u��<a]4���M��h��d8�]��vU6'�|Ö;2�7C����Li��9�pޕ��йMa�f���W	Ct* �h2�R�JDyg�
�T�!�T
w]U�d�+�����ڥa�;z�GFk#����'����)GM9�*6i�`�BS�O���E%��Ut�����gf����;O�ҶޕK���VF(�E���sqG/$��V8����ڹv�ODi%��*�PضQ�ʘn����]��3��o)u9k;���{�N�^2��N툔�2��u�{�E�cʂN�y�IU#��()�ص��S�w�/��=�	�:��l�=�שˆ�p��ca4z+���I0�"�� �&�e@v�ګ�3�X���=�
��%�ۅ�f�~�([�� <�aN�:�tL|dKb{2�,��jq6���4Xkkbb��Cr�8ە���s�A�M�@�;d!fb���78���֯Bȹ~2�8�dp�h���yQkr�EX�^})�P��4�_�o�u}�wa�l�����)<��x���--&uB��u��t��[f��e�Q��p�ǐ���y�[���*��)Ra�j���%A ��L9P��l��Њ��ke�����]�:/.3vۍ�V�l&
����겄ߔ�
D��
������γ�Nu�E^��|����<K>C��_���BtB��:[p�<���N�!L9�ʍ��G�4��2���;ůl�J@��[(f%n3Є*g\�<�l�
�kzX�W��'����iJ���b��f`�~�dT'>7{V泺�K���,Jl�hl�!��sLU0_L�;�x�������	�P� ޞ�@,�ʝ�m�/��L,��z�4�;S:�ɰ�^ޫ���N²��{��zCYPD�V�\�����A�jO���B뫹]ٮO���p�ّ�7�9=ӓ�����B��5�(i��B�m�)1�'E���� �����b�1������� L��rb�`j�,d��"�MCbq���[���L���������܆N��� ����~sFs�7`p���n�!��bdz����rC1^�tO�6���[�/=���zg���&/�RO�Q�:���t�d�l�n����UF�m����Ξ*�;qu�GE.o����ݛ�0QT�i�>8$�׎r�]�9�0nvJ�����-	���4p�~�|�_k�7�ȯKν��	���� �r(�ɕ�k2Тt��ӎ緥��~A���4�;��_����)>n���c�����P>
�d�n��l�66�ݵ<����-�~H9�Hb2��쒪w��e�n�X>oU(U�q'_j��c!�P�yӽL�e�?D��,��đ���!�W����mʁ]����G�Ĺ���z��Oe���ƶQXz�E���祺ꗞ���B�@Q�$$��ks��{�"U�S�;8b�}��a��ەX��N�P�Ԡ�����
��6z+�K���n�ښ�(��i3���ٶ�'�8���_o\f*Np�����{��=!�Xfކ7"�Zz�Sh�"���-��g9��\1k�aY��yoS]��]\���f s�f�%k���I	��E˾
pϹݖ��mE�z�qcU�'�#{��*�"����<< �u��5\�&�FF��룣9��}	MŊdj���.}w�D��JT����r�����=�i��糡#o�bl����Ң��V'N2*v��:�apDQ��멅�x�#��t2p�"�1{��Z�L�[�r/5�7��kxIp�|����֪��oX��X��2m]+อ
5�J��c$�t{���6;��9�>0�gɸ
j"��H�(�1�tl������O��ri�Z�=S�5�}$]�
q�#֮6Ş��6�Lb�!�"��f���!���%�茕p㗔r73m�e~S��U7����q���^m1��C���ٮ��c����'��]x���DY��#љ��R,�k�]2g:��C2�lXδ-�Ԩ]��H��w��!���؅��{a�Ss�M�L.��ٕ��ަ>,����TߌE&E��Up�Xz��Z����\�[�7"١���Sٹ)��f�T)�	����nlQ�
�M8��ڍ�M����\�ch�i�t`]���t�u�"��Z�K�r�R��n�@s���NN䝁�:�{�8瓪ָ�L{oJ�a튼{��]kN�FV,\�Z��!�'p�k�O���#�ҡ��Q�Q�w�9�Z�v�Q�������[�$��]q�x{�� �'�F�G�x���Ύݧ����<��㋁`x��U�XVE���-[n�T6�ge[�G�-XNÅeҍs���;aWDН:}A�������,߫E�3q���{����k��s�m�h�]X�GXN���]l�}1�z,()�R����r�A�4u���#q�:=v�Tj��Z��[��Ug���s~���=VPl����U����J�i�����*{����X��%ҋ��Т��Հ���5`[������䉋Z�vpm��v��-�Y@���֮�i��+Uו�d(���59�̅m��j'sөw�ϡ������sn���r�R�c�$0������o?x�v�)�<m^�IF(��ڍ��όQ���U	p�K��yI��|�O�aʊ񮬅��9�d{�Zj��:ڦ��-���W���jAōfj_7Fg�,F���X�#]
4
QQ@@�PL������:\t���S���2�{���~yJW�;
��[�m�('N&(6�i��k}��tÐm��b"��uw���ԙYn����I�FH����\�9W��y��yq��'����/H��}���'���z�)`Σ�ta��U�1��,��>��z��G�u��]YK�n��J�b�]l
;�-�������՘�!�u�_�YKǷrl�����gs"�z�SІG��U{"훌�v\U�ա/��+ɺ��-�^�g:������K3i��B׽�HPS(G��-M�쌇h�=�T؞���9�ٕp�7C��9��f9R�nk��m�HY%��٨��72F�F֊�+� �>����8�0�t 2Î�ؼΗ���8�L\_]b�o�v}�u�E�yV���n���a�+ƶ���D�7�u2�[�'�z5���t#���z��ȇ�C#|���mz$�s�^�E� t���G\�y5��tVD+���)v��q.Z��B݆�ǨC�:�=(�֫�b�ϐՆ.�v��-�UA��^�X'�M�Qn�Lv2oa	��m��Ȉ�41��֛��p�B�rd�Ԕc�qV1��X���1���P���
��:.���Į�u�������mF��6�yT��Tkc���X���Qu"���ލ��b�Nh._����ݪ�i�O��y��ާ`=����Y;���q��uI��YhJ� i�L��Ԥ�|]2d�ku��=��9��z�q-��Ds@]W�*��x���*���'%:(/������pɡ�u�
?����
�# ��H7:��ϫZ,]��Fc���.cW�ˮ�|��8�tO�SGzn�O��μu�0�_WnR���;}�u������{�z'�l�C�0������V�C�[���uYBT84 TIF (1�r�Q��X�M5`���m�A��8z|�]�8u�������1w�: �u�
aț2�-N^s�#�=5O5C�:�T��vk�B�u��s͐���Y<���\�Q��Jj�1���o�u;�BWL��ɸȡψ�ڵ5���Z�,Oy7S��C;ۘ�zt���[y���qFh0��@�&M�s�9 �v�#!�)3MCbq���S�]�)��� �$��#��E�PR�s�{�yG���Y��G0�Q��륿$O�.
�){o\kZ��冽�"9�����p�MF; ��q�H�P�hx�:X�r�p>&�{����Ó }������
7t�
/��)�G�']3|<&�N�+V���+��`5��y9�Ys��j�*�J~��N�a�
3ӧ�7Q�-Ԣ���L�����7�]�� �l��3v�T�6��h*�lM)�����%WDi.ȟ%��-K�~�ӜJ�xh�s�����v�����<m�={Y#�A�����t��9V��D���ڝ`5�YcU����h�^�b$7�Q��W���*���9��Ci[ruwv�8nn�#黋�dU�b���x���M%��kr�E"̝��吸�մ�`\I��{����tF���m�M@Q�? �1�*�m�:��M��L��#p_��|��UĄRkt�,�\E����z�ы��p��_z�z�41�
�D��*k�T�t�z�����y�ʦ�w*C�v'[�,	���
K�S�qT��- �G�.kT{{�T�2����;����p/�����(�:eE��VT��`���T��Ex�p5��43�۽T��%�s����Jr�MKp��]25M��@V]�LZ�`�1�p�k��K�[����>=����+�U�ǫ�/�B�<�N�<gD\(�z�ڝh� ��0]������j2Wl�D����o�M��P�!d�����:w=��qupW
��7��S���KQ|�H�[UK8&U"�V֑����C���7��q�d�� �_V�ig3���L^���7(d�0c P�}'�
����(�N�ɋ����j�K��Q��n�vk�� �Wm�c[a�� �<#��oh؇ ��\��Q�9t�⫴s�#8��|�(�gK�c��}y��J��Zq>ݨ㔮�6�m�%�mU�I0��82dպ�\쎏{M{su2���yd��
�)6��[i.�]0�WC�խ��읁��R�3M����w[9_>5u�Vs-�D*����{J�Q�y3�����/^�1�&�n5^��̥^?f��d0�{# ���l�q3�
�%���O8>�Z)`�ح�U��
��ζ-��%@:�edZ����V�zn��SJf������ F�js{e2�ȶ'Ǥ�=�Ux�M��s�=��\8��Z���=\*�)�~/ڷwUG~���������mO��p!A�2�ߨ�~�4��Ck�6�6b��҈9�k�z�wk« 2�8�!d�o�T�V{OD�Ch|D�B(_�_D3�F%�rVB~ܩ������3.n
Ar�k-�nÅ`�Q�a��8�����^ \+�:�[Fѷ�����
F&�� �Yn��{��-H�����N���˭��A�tƉ��)��H��[Ñ�+^i��r�P?P��6<F�wQ`/��E�Y���������z��6]�{5YT�m�n�]Z6��6!��h�%�7O| ���������sJ�tu�ہ�
d�^Q���}�؝`�!>�\P0|�Z��12������(���繐���Ra�ܻ{�}��7�C�Ǵ�"o���$�d���qeɖsn�gj�[�Ţ��J����ǒ��Q��M妴؃>.M�/7�R5�؊��.���C�������9���o9��p���k�#���X^����v�_DY��SeSWd�wF�2]]L�u�]]].5��mqiS�|J�]L��T�_fnV�V��@Q��j���W��r����W<��OĚ���{�Ď[s��}ݎ��U�tU�J����.ǎk���#(��),}�Ʋ	�v�CN���Җ���@�=�����	7��#+t1d�{D�RR�"-�dKg4��ٝ/F�y����-��m��U֭��>Dv���%{ۊ��ʼ�+C�����+�b�����m4@<���u�������0^u�����Se.���0r|��kWݦp�8���%��oMȥ&���B��"�q4��uj��7���KnL�J�=��d�r��MQ���dL`���Cq��P�}gj�l�n&�U�J]�F!N�E������R�κ�Ԟ�X��v�kf�Z�8�U�vX}�:+�e�j�@At�[����N�T/���h���g����S���ﻹ&���s@�Qۛ��17%�]L�
FW"��=�X����Nr�D�4:�&����C�h�/A�7o6�[�rz�a�w�(Ц�-݀i����R_!�p��6�*[q�P��Us;�-6�������v�^�}X��E�\�P^m+2.۩���)��#i#��V32�+�R)u^^r�K�%���Il���1��͢2�T����RgMr�~��/ұ��ہ�^Ӭ���|W��v�Z�����i�����A��6q:��,Uݽ��$�\��a�������\����u;2S���K'�[���
����5���:���]ҝ�V��E�͍�#�MEoR�[s0w��VD�]�,�MΧ>�8�2>ƆmgVSR_m5�P�x`$W��|�����zũ�.�hr�n�ܡV����$��2�bUr����/z�p��ƾj�}��m;�����N��7�����T}�+۝D7]������`n�I	nTJ�+�.J��`r`%{w�pauRa�N�܂��buϤ���������Yã>�d����b��[�Y͑�XBmU�ܴ�����M�҂�A��(-�����2�r�q^�C!��>@X��7xi���Ի;���|�b꩒��̦"]A�<���i��&���
y�ܥɀ�@�2�6�ۛ�[�\t��C�vfi�f�=P��x\����JH�]�R��&����,f\v���g�o]C��6�v�X�������.X/��$"e%�����k��x+a��.�P�_ak��q���?2�P]�j.�gb���v�ھ�t�͍��  �*��
 �J&��J�� ���"b�!�����*�����hb�*
��*��)"������i)�
)�J&��J"���""��2�
JC#
�*�)((���������`*�h�i�*��b��h�$���*���h� ���i�hH�"h�"`i(h(*�� "
Jb
"���h������
h����"�F$**j�*��)�Ƃ�(�(*�h����)�(�� �Ȥj ����� � �����b*���
�h���+02)�����))��"���� "(�� ���
�j��)("�����H*��)�*
h�*�����"������"���h��%��*���3%�`�"H���(2�
*����̦�$����b*���������&	������")���)�s��kγ?u��v����d�z���n�I(��]<)���<��kR�S�"��ԡ9ZAh�B]m=+�j$�yE���DӐ��}��V~���2�������:�P1����$���Z����V܈�ý��S�U�t�sS�Aq|�x���WH��~�F������G����	�!42���-p��s�\y�pt_���}��Lד,F���:�&�R������1V���8I�&s~�M��;&�_�fv<�U��Ct�a����������誱ӷ�Sތ�L0B����j��@�U�~�v\U�ա/u��LW��^�/���]y�m��]n+�,bL����W��-��q�j�]�M�����Y�s�FB�Lj"�Ep�C�nɿu�5|nd��ފ�+� �|)z�2#��`�Y�j�L�ȻaX�M��Dj��y�K����Ѣ�<�QP�7��1��?�'�B���М\��'���Vץ���4BSs���N�Nˆ�P��ca4z+�^��0�#��lB����w�q����Ġt�;p��iۇ塬P�a�p�8����y���&u�P��������%��%_��ާL�X@U=����w^*�@���?3�{�/�$�ca�]���ح�Zzڬ�A�gQ���o^>�{���)���g!(mF�a�V�8U�����C��ˌbb��ce�����!v���"�B��{�:n������"[���蘡�������ܬ�旺��{�n�.�����e�q"^�"Z5^��� 4-�
��=p��讥^}6BÆ����U$';��l�<�(�e�ԋ���N�Q(B�M��<~�l�=�x�W�%��6�b��+��?Z�:	֙Vrb�*���<«�Hx����}�N�C����˺㫍ӃX�=�tt��fT���YakP�)�e4Hg�buO"�^�f�iS=�#���=s*S�ap�5ry�sn�n�d�Iפ#D�F�q9��7�ky8�*�f�q�$"���ٮ�`�!S7��S��(�2�d<rtAx�dOP��;�;x<������'͚iHVM�EϮ�Қ��O%�DD&�u0
!��qBB-�Q+�ܚɫeE������P����lR�Nv,x>5�x����N^:k*��Ϋ�Wڇ-�ź= �>�=Ҳ��P��h�V��ቑ諾{u�Ԏ�_�3`�^4nѾ���%�v$����TL�W|h��X���f˻ާ���aV9eMv�Skk�E���|w�v❓���eԓ��W5L8�Rڑ,�\�n`���z���.-F���t۽�V�X��5��b;ȥ+�Q��+[�� �5�쯳��빌���C�>c|��~��j,c�>�
��0���mÊQ�v��Ӻ2�;�&2{k��i�q���b�qH�~��t�vtC����Iaϥ�ǳ�i�֝_!��p�R͕r�
;�VP�'O�m����|TS��ȇ�Y9����uB{wI�aJ��õ��b��Mlѐa3�-��*�`��p�����c�����Gvr��J���k�9,��0�Z,�P�j�/x��Sa�>x;*��i��
j�.�8sȘWN�w0�r��|ոX]-� taG�ZW��=I����,��G^��b���ˑ�wKY�Y���e2��FEy��9�n����蒼z�� �v񲳕m_�����4�fD�Jҟm2�'f�]�vSGL�z����*
���06z�Zu�-�YyT���3�磢��*�`�۝�\%7�dj�	���>�ʘ�-v��NFs�Gz���]�y�Jɯ1�]ш����B��y�����EB�κ�̙�\U���PZ24W��to_uYշ��6�ް��X�����.���� ���S6G�*.��
ˠ3����}��K@�̙���XM��1�Y�����p���ǩDk��"ۭ+K�ݽ��v�����p������Δ��h"	��4$uy��1P��5������|E��t���F�=���~�-+�h^3 �@#@s��|*��[�3Jv���M�5������9���W4-mLwE)}>0����l���	�1�5ϧ=��������Z�Nl�mmH0�{Y8SwCj/��p���1����05���p���o����6E�B8�&sh��-�P]��]���<��xӳ�g��)�U��m�T�����^�*���S#u�G}����o��aW,�ȥuY�e8�Τ)� � 벲-N6�G:u�=qWW{ѯh]ov�%vb��FD-*%X�3���
�")�z#%;ܪ����W���sVq�g�h�J�1�p�%���~j���P?_��H�uö�Ƕ���V�36��w�f�0huq`sU�,�N,zYga$z��z&���8�<a��^�4DU��Q�[��Ա��K�� �V5�۠�/J5�K#`��@�lW�@�^�oR����=�C��Ί�033�2��+4R��&M�n��^Zj���oo�>�{��Gx-�*E�h*�Ӎ��N�����{�1��PA�6�R���l���<�̍ۙ�.���կ+��\�Ƕŉo-c��y'Q]��u6�N.3��p�dY���j�.�{ϐ�>Dװ�pb��n��g� �w�#���S�W��������׸��Q�K7�^�!5A˺5
�HQ�6��E����]3J��XnlB��W��2a^�'�>}Ƿ[���� G|��	0[�.������>�,�}B5V���5v룢�Gr�d_8�.��A0�,d�P6>a2�:ׅ#7HV��c0j��¸ƈ���oc,�ֶ�G�bVX�L�}�ME[S��t��궎��iA� ;�;_1=���(5Q>�ļ���u�}y�1W���K��\['�R`����r��ud*��!k鐛�ۮ��su��"�%�Tn;��pd8Z�Ծn��&X���P��t(�
QQ9������bC��Q�̌s�(�eb�(gZ�ؕ[�a��e����+L�L��V�,�Lf�9"����\;�_��dU{ё�̟de�p-�qWƐ�����b�Gv�U�����ov`{��o�u	�G�8��}Xp@�U��lOt��:�LDH�F�K1%vطbs��so2�M��mMЉ�U[5��4��-���B.�=�[c'+!����1��٭k3^`��α��{2���ME�枴�J��O�c�N�ժ��<c9P�u�Z��#���6]��?(lgD�������]��𗷍-[�|�v�3��tV�U`��j�x:�-���+� �Rʚ��:C�����3�^2jآ��ɺP�ZC�̨�f�|F��dj*�ixf�U���~H[�-�7�5�7qe>�c��5��"B�؝4��u�r�%�X�����k�>&�J�x#u��^�4��\i��/G_DԔ%�ˁ]�(Q~��n��0\��vݸ�C�:�%�z���5�A���܆�L6�'4OX�6��b�����x����߸*�V䷤��-'���r��1����'�4�P2�8�E�T&��<���C��ԫϥ\�]-�w�v23#\����-��6..�>�T�oظ�_��k5k(TSys�8�B���V*p�{�����	ܚ���x!U�W�{/����^���͡�F��]��jt<*Շw��ݟXN�(J�F��ePtHf�[�Ǵ�5=��{U^N�v�ڹtb��g1(�!��^�]tA��g��s'D	פn�'6t��EaHG���J��9�<����A��\F�]�p8t�뒗j����L���U�X�+�=��4̀�.т�(+��	�oC��Wv'����۝OaF���Vgf�+R3�:��o �nj십����{���eV1�����gQ�{�=���Rj��H��*�Ddu�
Em(1]���B��s0\�l��P��N�ڙУm�J��`�A6 �ۦ�P�J�W����])(,1��I�q��u<�����۵��r����}*#��.de���V��X�/�*}GXG��u���(z�
��z�<����7cW1�HKOh1b[��n��^�.��"�{K<Z9�
�#<r��2�1l���{��@.A�F]o����-���+�Pn��p{F��(=>��Te,�^��u5ݴwYx�&���s�����w��bwqb�R)������l:�Y���cӔ~����Bk\�6$��®^Gb���ۅ:|�l�n^ ��[��l���{z%I5r���7��nk���C9 ��dn�Mt~�*�d�S��l�7��[��%9k;9�:��w=V̻��c�=���;2`l ����!6ϟd�S���e�����T���x����4����|��
YY-z$tiF�&v$�>�!q�(�֕	�m��1�����.�f�{+[$���Yݔ�59:����z���x��AX�L��Q���R��e��Q�h|.��1��7wJ#��wm���gE������ںf�s����h���!8��ZfQ�r_p�����ݺy�,0���-�=r�s�������'.�=�$��6���٬qZ�Df�x'[�&�6�%���
�$�Ш��T2�tq�om�]]�HΖp���c��g�m�ó{.���QA��T[�YSaizTe�|�u+��^M�߽9���{o����x�K�B�P=]
3�;nEBSP�25M��@O�N�V��AD����?4�G%Y\.��{��R:���萯�����ɗ�t]=�|{+n^)J΁.Q�㽝Q�����'^��uxѿ��
_0�F�x�������(��L嶱���;���f>}X�ytr��T��"����Ҿ	�Z*Et��#)*%�Z�h;��֟��]_
R{Nũaό=���Pl���fd
��}$p**��:�0R��2��ji�ߣ��a��>L5�5!>�ƶ�!�6��<沎Ê�@�.W Ƶ;����z�����[��<粎F�b��cv���!�s��,'O�;�ӥ��7r��bc�}�$H�Z�8)`�"���׌��v*�fS���B�rJ�u��Y�T�����|j-wF��)�S|�*f�NtW��Ĭ�`R�A�X�X%t�ǝ\�XA(��v=�HL1��'V�Q� �a�픭}�Y�˸*N���BN�:(������q��4�@�tt���t9�|[]���O���o4IS�ɬ�r���u*�ZSL^���U�?"�L\3`pde>*H8\Z�*�`Sc%����S�߮�7�=�[��)�7�.��u�'��$猽/�[Zy.�_p!A�2��q
�M8Fl�a��.��_,��؅B�9��d�qbYV�6��~�k��c�jF/�z�<������Et&��{g��[ܠ��?[5�6�ڗ ������p�J5�94s�]8�3�=[
:�S�'�����0(�NTM�p���V�s��/�t��N���u�]*�m(ˍ�G��a	أ86xɅ��;|[���}*�����-�t��
i�S���YY@��\��T��&X���B�f�%Ŗ���(q����U�7��fc\��آ���o�'���_����f�-j���B�X�;�T���y��̽�Ujh�͊�[!E�^u��ɚ�5#�|���9
�����h�7�cs7��#Z㤏�JK��s��@�������R�`�8
��:�V̅��:�F�e`²҇O`�t/��N~��xn���C��Ӽ��a1�9�,ŤXsOFkb����(�=�
[#a�����{6b�ke����[L�v�w���=;�>�x�9�O;z����ҭ*��(��1����.L�@
<"�L>�%nb��/%�I�S[���ۃ���48���u�\{}��L�n�L�܋$k�G�o���u�@��n�,�Q�̅��F�+������X+�r��9:q0���x���a����޸W�o�f�>2]B�U��ё������VE��e�X�hK��l��n����b9v��v�ٓ��sKr��%e����g R�2�^��T؞���Gtb�1���51�+��wqYd甲��ɺ���"g�p�#l�AǦ���';�Y��o'!�gD8���!�P�}��5��M�D��\m1H���wZ�pT������Y"b�?f�p��%*tӗ�שˆ�p��ccj�R���;���N�q]�q�T)�~QqE�2�@됣�zv��{�3˱�P�mۀq�-��&e��#9�>u= ��P��"Z�(��砇��H=�]����{���ߣ�F��WҰ��1�F7�y�8퐄����BW�� �T&���*-nP��UZ��xa��kp1��xcXtD��]v�x���n�4
�U�2k��|8.��vLj�:e؎�8U�\X�ky�%�\�����[���Ph�5>�G���-,1�q��w���{̩Y{Z��d�걼�<��o:�^�&��m讼�1�1��Ȗ419�V�h'��s�n��-X��D���Ֆ_q�e�cB)d����.p��V2�QQ�M��5J S�U�q��nv�i�U�LK8�Y�2�_SS��fdIN���	C��`�t묦�f�ݠ[��<��p��rK$K:5�z�'���5֎[�U��YI��-T�|wA�-|�W����a����;�Ce��P�w�'�ނ�9��"9K��N�6ՙ�w�����k���	��@
�3���;8!Oy_]К��R�un@U�ElҖ�q�V�9&搹�|���:�-�t�+��S���H��z���K��aӗ�H���E�K4lY����!ޥ�҄�vF��c��F�Q��X�z=AC���L/��w`�7Hv���݊Ob�NNd��z�\:��,�+W]F�����!�-U���tr�a���e���M ��ssg�����d�oPXVM�UrH&��l�$�U^Ơ�T}��n�1yjo:�ȋ���q�.]iK� ����_�(k"�d��kvFhđ�:|\诣g��\�N��S:<���x��>u����0ę�z=l,�R�힮7Soif�|a\L�N�K��د����rȤ+AV'�z�7mUJ4h���/[}[�Dk0��í����]87�K(�y��;�.�ҵ&n-�o�4ǹ�yKZ��
����~�7��&�����7�wJу,��1=�@����L�7Y���2D���D)Ձ�,� �=����>�u�]#yA��(�U��շ���rU�VK��I[�^E�t�G���zһ̬�[+���g[�[Ӳě����ە��W]��Q�to��R�Bm^��(�8a�79�=v��t���n&d�j'yKgJct�X��Fe���v����<�(S���G������;��.���i�g��җ����v��ٽc�
�X�7��N�*��6��M9�iQ����u2�Th6�memLj8���;���YN�/m��*hv���7�2��������ʷn����(�����;�U�{�o����v�	}o-4���V�sC��*p}���#ہ����y�~�$[O�}�<o�)
��!���ڮU�?��Gn��x`���^�\�R����`��*ue3lf}�������<�T�����c3�m� s_b{�t���`���w^��u7�K���0R)�ޭ�q���=��yp1�|f�FE�B��X�|�D��Yl��Ї$�kC��Q��,u����8䵻� ��̍�7�z�Բ�=�	Kw�V]��D�EM5�QQ$IETSSMSUMARD�QUSP���1�i�"
h�***� �*j��&�b(�bH�b�����
(������)*!��+,)�Z(�"��h����**��
*���"j�j�����(�����0���j`&*���3 Ȫ�!������������b�&� "*�������Ȉ*��,����H�""���)i�*"����������i2ª)"j���h��)(���i�a"
&*�b��r&f)�b*&)�����*�#()�)�"�������&��ib�*!�b
����"� ������,)�b��# ���`�j"j)�������
j��f���" ����"�(��¢�&��bJ����Bj��"(**HC�� �M�/Vs�<�ƭ�j�5oeÃ�=)Q2\+9����&TO�WL�{��b�1u��N��o:�fR�w�AmF�#x�.��S�-�����B�߼��(ߓ..�X��=����	X��>�1u^C���������uj�Zg����e��Pn�ʿ2:�Ťh�Bxdj&�Q�R�ƨ��]��ܒ'6X:�߶](���Z�� ]X�}˭��d�	�.�<�Q8_s}�<J��?1�z���~���C��J.�c�ׄk]�2�ł_m�s8 ��/(=�Me�A��w��Y�����4FC�ȭ�;5ӄ!
��fb��d(p,�gD�#�c��_Q����	�#ѣA�5�4�+�77>7{V�����\���A�le�����9�y���/ͺ����C�<S��/���*}GY*x�6)}���U�Τ��^�[�1��ng)��W�a!-���73n��:����ٚC׻+����٫�ϟ�D��^�ڼ�����v��oHBvW���l�8��l�����>���]�t�ll���NC���P��֎xT�Tگ^�bvwS�����z��{����A{2�Yɳ�R�R޾�/�m>X=b�Y8.�e:6�V*��R66��^�L�튒�ICiǇ�OR��4�<��M�\�ـ����]�ls�X��T&���G�;�����ėa3t�88�^sy]3_:�@MƳ��+;f�.�
t��}�l/o�q�7���4m}
��V�G�����2Wk�>�k�<i{ʞF�7{�6�G����]��~>�C98M)�dn�k�+�iV�==T�<�>nRLSθx���X���[֐�3��(;$u��ut� Anx�B2��쒪cM���&�l����vY�������CZ����x"GF�b6'=���!�W��D�a;
xZۃ��t%�S�(,4�pj8�Xj
�o�g������#�ux� ��Z:�ގ�W�N,�:5������#m�ݛ�w��P���VTߖ�PR�_��z���8T��
z(;�>�%B���У�c��T%5
��9�[��;��[/qk�UXn���+��zW�ј�U�1EaQ�/�E���Ӈ�����ۻ�g8,T\k����h�Ae8")D�;�cg:St<W��!d��߳O>�{s��jd���0���6ڹ�s����ؒ��7}ή���2�EH����
G����wi�\眘"��j�&�wT�1��j�g�5��X�B�O^�z;C��Y�Ev[cn����#e���k�(@�pv��	B�,k8VQ���DiL`�홓d��ޠQ!fq1�V�LWi�G2�-;�(lz�v�-(� �������E�SmV�Q���[�cU8�8����f�(6P�x&`�@���xJ�`p9
/wg���Feth*�����].�U�.���>�v�8��ۜm/̇ �g�a�����a�]4����)�7D)�gl�7��v67i׏�BG!���l�NǪo���R�{5A�9�ܚ�EK>��>�-���{��q�}���Z� �vVE��V�8u���B�ަBWú���+MM(8i�����ǌV�'_���ޥ�Q���x � �W i:�ъ{�͊�������Xo��[αM)�鞡>�\2���!���-v�Q��%1����\�q�Al�m�@��85�lg����à�u�!������ES�M���օ��q���vu6�ۗ:Ar�X�n�v+.�k�Yml�~�<����]>]�y���Ж��@�V(�Nz'e�j��g�F�f���P�����pIAF����Q�k �=N�=��^�����bGA\w>i�@���o��X�;Qt��*���S>q��z�}(�*5�����w��۶�*��U�ё9��vC��a�lkSue{xȊņz���O^A|DY�X�e'%ߕ�#I��W������8��*�LqgY���|i�x]ƫ�h��q�}��� �TÝ��#��YH�M�Dh���*�QY��V5.�![>�������%�p7����b��[�����(���/���ʣ'T�쇧�L(*kl�M>�=�^��2���f��kWH�́HV��;3�W��Df�z'/9���
�CS��Qfá��:���N���\c�����,&6[���q8/��q.w�RF�'n|X�T����vxj���<�����`�8׹�^�(v��d��܎�4��}�:
��y��o�+�������K��w|�b2��X�p3�W DF@�]��p{
A,1[�ؘ
�p�q�1Ӄ�j�rUnE�������<�iW
H�X&ާ��ڦ��7�x��5�ŋ����)9؟F;.*�jЖ滑^t����,���}x*��ꞛ0;�9��Ρ+(����,R�V<��rn؛~�I�cW.>�Z�.��O�R�fU��7C����M�{U��ih�{�U�IdA���x����ӥԅ�gr(��nNÜ,C��b��S/�#S��8ɫ9@�\n��N�\m9��18Qk��c�Z����#N��V��W�=���$Գݩ2�� �������}8�n�0(�`U���ދr��b�xt�t<{�\�{r��|�V+�fQL�}��Af���D|'j eh�7��'`��wk���$��k�v�k��{�q��l;%�p�7S6iȰg#�5�����M9x�S��/:���(��6y�U�q.���c27�BF*\Pb������e@��(�Nӷ@���ޱBݷn=�U��ײ��o/O.rZ�}�բ�ϼ��a�%�=tB֫�b������:i�A�����W3������� 	�;`�a�yq�!w�F̞z&��!��젾jym�r�}f��oGw�8'v|���l�t��P�Z���=��7�ˋ��ޝ��P��ș�oOF�Uw]���HU���������g�ߺ�u�S��&4,Ut%Q��lm���tL�Ocj�pKr!OF1F��<�]��J�7�����;�r���3Ya0�/���1+=�$���wҠtH�_��]��P߾J.�c��p/Q�!:!T�u�n)�; ���j엢��c�5v �}!�
D�N$��Y 9���vk�B�oY��,��GP�pe��[��L�.GEd>��G:�P�L�|H^5ı�x��Ls���]��O{�����c�ݬ)��/y��,� V[\����4�v�&�B�� �CX���@eMy6�T����e�w}�,Q�;�c��7������u�K�Z�DĦ��Y��n�����]lo7h��	N�P���)h��l�q\/:��y�;�n�SΗj�.�\�p���dD&�u1A��nMd�˂g@�Ȥ'`dɹnL\{$�Z��"!���u�|vf�r!�Td	Ƕ ς����J}�b/|�9C�]m,�^�0��5s���-�<�t���7�e�sѣ�!����ٸq]���N��Ξ�M���?f��y��m;��c�:v�ʝ��}y}HC���LC�r�N�<�U�""�h9�a�[HҸ�Sq5 ��|aψ$��p�����#�Nt��.�r�ϩE���C1g�`�+�R��o+��WG��X�C�t+���E�"��e��-l�g�]j�a��9pH�����=U�2�[��Y@�!(�M@���6Anz� �g̢��1˗V�>N��,,��Oa��o���W���V��x�[/H�ҍ��I��C�g��Y!=<բ����iD`��hMM�p+�Ӟ��G�AP���
�<�x!�l��bX8���s���:M]<I��E2@p�A� ��w:��e3���{.�
�2���YR��W&	�'k�y1�eu�tmz���]����j�36e�ѤꝤ/WIVѸ����-:��;��˳|٘j�[��r�wח��s��H�z�q���;�믂��5��^}�֤NAu1��{#����nf:�s��[*�A� �6`l��*��
������;	M��#T��7�'�/�u��QC]�Į3 s]�K�A��/5b��O�"���5NL��]��׏<1��M���r�3{M�{��
�]~��u������"H@�39қ���G�J-��o�Փ}���31�9}��>׈�]�.�L/�*�WJ�&V�"�mi���OU��os��i���P;�S��\[����L��6P�x&`�@�k>�����BZ�"&k�e<���j鵣Tl0u78*sf����P�]�8��b�!�"��f��oh���X����}��)
O@(Z��b�席��J�g��-�U�׻v���;i��jE&��ZCN*T����U�B�|�"�Ks@�
��C2�lX�-���I�Y5��V���{�����q�n�T���TlBҮ�T�� �qh�L`�l�FCʋ�	<Z���f⣔*w��(=U�e�ذ$猽�~j����U��P(3���kw������y,Yo��k��@������%��:.9EL�"�8[oxL�^�n#'n+o�Q�+s��l�w��*��M*��`���y搘�Wj���dȭ��gSe\�G=���N]�燨d�S�ĸ�LJUȲ�+V%�����`竮ْuک��޺7!n�hSe�n�q~�B��I��O%����s{b�2޳L��7�����Ç]��M�q�.t��kSn��eҍs���:Js��o�N�م�eİ.H�=��H�N˅7�ջ��q��"uek��3J��O,�U��)�خ�ǫ`����8Ɖ�aO0�����|���v����>�S�1��̞
�Gl|ࡽ.O��Z�n]I| ���"��:](��'�@Wh��*��̕l7v�7Η�g�����'w��+�h�L�l5��kH���`�a��>*��Ng�<��纑5��.�E���59�d(�~t::�����Vx� )�ʠ�S���"T�Χ�*�5Ȼ���@-���NӉ��E�ߵAq}���T�X%�����F��e��V��E��A��]u��<6��jO��K:�=}��q�d���A	�#�]�����9S��/���ձz�Ƌ�k�������� �����'�H4bš��7/y(ȹY$ݚ�$�N�nؠ��gH��y���k���k5��U{�LN��J�ӕ3�39/y꿗��_�LJ��FF�umf���e	t���Ud�{`�U)��Z�W4��,j쾗�����@�r�U����N1ґΈ�����1]�����:�0��i��of��|d�C�TFFCv*��n�dt\Wv���1gK9�ѽ�Em	O��`
�n�([����kf��� h�`�4��JFC�����ܺ��NR��1�k���9�P�7C��yWaW�,��BVW�fQB�w�kH;�����m��h3/Z�R.8�PC��C�̨���6/����YJE`�1
sX^>�cL{^����Ȟ��0�B�lӎȐ�%7:i�L����T���-R�
<�q��Rt�r�n�V���>&�W
.(�&�YP(v�Ditᩘ.]�k-�j,��ӵan��B@�se�= �=CO��Kbz�D mWD��@���A4)���Z�Z�y3�flRʞ~���ٱ�����5*�����̆"�"G�lX�]eg	�E�EgwOr�uU���~�^})�P��3A�vQ�ˋ� lOzv:�(BNGH��ъ���G����ΟA�[���EE���u�y~�Ι\�W&(,Ut&Е$���z�g�Z>˂%��'C2EL��ު�5���9����[dt/)BIV�yK9Zm;i�9�>�V徼��6uY#�F�er�C��zi���R�l���r����E�s�݈�+�7���U��Wu�f+�bv���,|[i��a�:VՆm�|.r�یo�<���3Օܥn ��1��
5�^-о�T�[/���@��w������Ӫ���ĩJ���&+w�jb�d	��'�b��i���@g��ϒ���U��k��u����nŶ�dkwg��	�X�Z[�����U!���+�f�{�]��B3�7�V)V�iS�y���9/ɐ��(VCq8 � �����i�W�M�En|cR��s�h㵪���֣�)�"I���ϲ�5�W�����T; ��rܾ��WOg
�sK��}��������܋�i�lN5��	nf-��9״�s6f�K�?5.���;��o��Nt;����{�p�^xf]�=o����l�8��QcP0U����.Z�ow+��l�v��'+�p7������<6�_�zQ�~^z>�qo'"}їu=�����>&�N+j?/����Z�>��R�Vp�6|�;˪ܺН�Sڮ6KoQc�����qI�:��o��<}�	^7�[V)
2`�|C�N�C�:q�'\۸Aɣ1�oEN&b<ƻiT�-�j�k��b�P����r�c�	���7�:_Pα�j+Je�qU����G��)mt��a�e��96	����9Ҹ�G�Qݧj�8P�4�V:�PD�L�ޗc�m�;��N��@I�v�N�ҳ��Z�n���9֯���]�&*|����tK���r�M�ٗ�u���♮��z!�jh�;q��I;f7ί��N�Tg���z��=ǟZu���+X��F�W��/GY���'��-���x$��4V��CRX�j�O�,��.��Ĵ�m�u`���/��.A@UƘ*�ͷNѶ��[$^�nl�ۤ��t�K�f6�9\ٝ�����a�;#���o4���8%nкp<,p�vV�5\|��#ٕ����cu�d��X�۱ī�G�g؞��u�|.��ۉݼ�-�q�Ih�#6!5�^Ro�t�TM�*��+�TV���q8����ˬhd�U��1{�YJ������u�&r.�� ���hM�5uk�p�"�7V�v8�E�Nݵ��V�v����sB)���7tU=�U����o<em������HH�Ē���/b��<{b$�S6����/�W!U(������軲VW/�/z���hI���$'U�`�)�\u�,Ȏ��.�Dt��� ���hވ볪�Y��u[ڈ)�N��R�u�&;qq`um�fG�5Ǉ^u��J<�Z��1��l�9�V���w�ئ9%�q|�җrc��%#&��Ԋ-:6��ɴ�Yh9��[���G�_p'���:���^·Z�#�d�@�՝i��Q���%v��i죒�ٖx$`�}��(s�:C��
�Vk�����ge�)�Wz{���Kb���:v)�r�7�+���T=uɚV�4	�h	��Qޮ�в���s���p�kUL�]AL�LR���KF�� �J�~�*^�Lv�b��noF��%��:
�t�T�ar�T�j�q+2͉]M���rK&6����\H�꣥fW�a0J�O��8+�����Y!!t�ݶ@���b�PIt���!-J��'�t�g�;��^�w�dA5v�|5�6oiF�����(0����C�JDnX��\����JD��8��S�V!O/qBSq�k�k�ˎ��b[�M��5B����&Gg��QU�^�W]�0U�ۛ�
i�.ZeU��o�dX/r��Ⱔ�.�͆��-.9+$�	Y��Õ�����u��u�)R�;�s�t]��Ǵ9#�@������}���;��6�me.�nS�[�:��N���^e�.�u��i?�?��뙘,Yil8L2�+�N4�oq?k����ꖩMk�x*r�:���1�phm
�CT��+(rqE�n,��<y�;=�v��[c�0�9UT���b �������rf� ���j���Bb*bh&����j��&���i�*b�hfb	�"��� ��j
(����b&������`��b�)"&�**&��j�i����������)��J��"J�*
���j��&*
H���"��(��j"�j(�)����b(�*�������)�J(*J*��J(**j����"�*J��Jj& ���&bh�**��*�*����h��������*�)�����Z�d��$���*j*�����d�""
�"��*����j����)",���I�"���*�"h&������f*��*�&b"�������h�Veo	"Y�B��\��&z���Uʹ/���mźW:]��rt��Ф��raΓ��}l�k�|���Î=B��`��3jU��' _�R|Սv�穪��-h�ڬ�jTF��R.�"Wo	}���i[�KR@Ϲ�5�6��ep^�|�}j��Z��Q�vJϔ�ח�Q+�7�Rd�9��X�p��tX�-�	�r�h�4��sQ�"ڂ�[�FEy��8�]R��~�ո�,_jR�LK~*6� l*
�QQ5��}�)�-_���q|�K�K� ���H���章����iP]�*
�=�%�T	��K�Cg��G+tԸ������p�_g�p�/$�x�M�M��Tߖ�PF#����4Ʋ��
.��i�X|���I�H�{�����ЭQ�Q����h���"4 ȓ�`�D�7қ��=
��K��)����p̉��N��>Q]~�s籺qq(M��9 L93^�*'D�/]�p���O*�{Q]�*v3O�%@��jM�S�r����m�6^32gҤ�ɾ��dNv��+��P[4�\�����n݅ �u�s���ņ�T�����z���>���е<���Rɀ@��S^��r[R%n_a��L�ǣ��8LTqj��w9p��昳Sf�-�Z)�,�*���.�h|��n�sRoG;M����
�:���j��K{.IO��2fԓQ(���ۙٽ���MS1�s�Rt!ܦ�e*����QG9yG#hf+7mߎ�B�U�����r�ݯ@3=����5����|�溅(�#�4��V*�fS�����Y=��4����-����b@��dZ�IW	[��sMM(8i������q_+^�n���>��ލ�����˞ ��w�:�UÁ~z���W�~o��[�u�iNS���ל�J3S�8�l��ju�\�]7��i�i��Cv#hSgn���N/��[;��R�i��9���"����+�l�7��aψ�DW��C��J���n\�ʿk-�v+.�k�.��Y�N����J�x4�8�@�lP!��]'ԏD֗
W��79�㗁+�lvuv�щ�kp�ҙ�ّ���˭���}1�z&S�F��$(���;�����ݯ�q���j~b��'�m�'Rj�i�v��}�����r^z�|�= �L�	]P��t��-S>���N<�p��I��Nܿ};*xm���+bz��I��=�P�Ce���?��t���ow=*�md�ߎl=}M����%�1
e4S�z��3��W2S㓷
w��{�p���S��^�g��s���	B���iaTQ�;'����Fvwd�;�8ϟ\
�E �{�_gm-"M���o����Js*;ʛ2af��X!Im�ֲ�N�ͤ�:E=�AE���59̅o·Cg*�'W�j.1�	Q#5�#A�=I����(��c���Tz}[[���+�����Uz\,���2������\3��#:������r�k�!�s|�8μ�X����Ծn����Rz����8��q�#6�\�X�l�o�(��
&�X(�et���ł��܃�����'1]f%xVo*و���(��Э2��Mo;P�Up!A�����7�����u�z� ϻ:�gfrx����u�y7Sn��+:���EL�N�-�x�@�y��fW;S�e^kD�k��@vU6'���sC�*��n�Ek!1�{Szf2�{)�=���;�ef8�.��� 	o �}K֬Rmq��PC��C�̨�fŧ�::3Yd�u��6:.c��fL�cP��~`�b�<F4�Y��7%�h�BS~�4�|Z�q�
��Js�¼=��tkwv-�����(��Ѡ�s�C��Bl��vHP��;N�=0\��q�2�싾��J�$g+�"R]1�{��#�rC���J��c[6�[�� ���nc��ng]l�&������j�G�����s/�4�77e�JlxwO[��*������tڴ��ՠ,yʛ,eA���"뛎���Y�؞�(�Ov���m*Q�!�S�J= ��WD��>"D�'�QZ����A�d�P��sP�;W:.�؄mʇ;�5 ���8쐻�#fxl�g��+�C����m�N�3���Q�����hsy��n
�r��s��G@L���~��ލ��eoP�=;9V�+y#���S�<}m�)������`y~�֙NB�1�]	p�+��!�Ȼŵ�N^���Z]*򂜱�9;dc��Q���P.�S��e���'4���)��뗹��V,�-ʁ ���HF ( G�ʫ�ʳ��bQtC�#>�]g�n'�k�#8<��1T/e�]��: ��u��Ñ$J(�
Ā涔��v�����lNv��$`F�/͙�S~l�P7\�hs�FP�E�8��f��d�d
s#Gs�|l`����|�5�]���P9-�f����>P�.��
�X��]�p�n����J��1p�VE���^i�lN5���c|-�t|��f��2Pn^2\GU��De��5w%>I�H^,�sV��β�<q�r�ӳP��+�x͠ҷ�6@�kr�}O(_`�W�.��&ˮ-ka�;��\E-DY�q��Dt�Ê�����gc'1����St5���ŗ���9v�;C+�_(�SOU�EúRVz�!���7G��=t�"}�ѽ!}��6{%q]����Y��S���ˤ�ѱ!tyb��*�{*����X���uٻ��a����L*���۵��:8��nr's�Wg��)��;SÀ��Lߢ�(��ݱ�������(�9�ȇ�Y|7�]>�g"�M)� �f@KV�VE�[�Cψ�o��X�;�nˮ_1�zl�r*�LĽ�Z�N����j_iAG<\FQ̊�9ƞ���.��H"��N���6�z���:��)ed�"GF�lL�M������%�Y��h^�$!Q���nT
����G��T$���A��9��6�+���O�����N�T;�����R*'s��
6�P,;7��
5g��ܱ��Nu�*t�C��YSoH�*�L��"\@�l8Pog��F��Z�ۇ9��#�����9%-�����T�Z�^F#�ъl�k*S@Q����Ё�T�7������k՝�]N���i��m#ي��Lc������}cN\����D�ڴ�Pb��տn! ���!�k����Wh���vj=�!�G�u7�h�h����R˝��������mnL�
C=�m�����m��HnJ=;�_+��Q�'T�	Ӈ��\(��_�×�Տ������RGW��4��*��}ݏ�N��#g�=e�NyO�Wk�e��.�L/
ut�pL��*�):�� 7�!O��o!���z����I�4;([�c����z��������32��0;m��+{���#�Tl/}t�`i��f��_I�\)n�蘏lA�� ��P�I��(�1-.pW��B8��|oh�(�!��t�J���/��m{1Xر�n�ln��2*����r�)5x�f;��{{n���=9q�����_R�����F�>�ݏ:�~]j�-mPBp���^v);A\cj�ted[��j�s�[��"�LUȩ������╯	�+ǘ���V�D�Ի�w�����=��\8�W���bǽ8����x*b�C�����t� >
�;�Դp�~�FZ��-�4��Cj6�6q�Y�[��,����=S�2�ΕO�S��1;�����\�B����4�mq�.�\���B݆�8^�Syz��v�rκ�q@�9{�fU�\'���{oסP�Y.(bs
�0�wB䕶�k��n��}�P����b������N��7�O� ������W}�
v�6���u�ZZ�J���q�g�3�P����ֺ�"씦& �;�����+�t����N�cb�C¿
 R����.�7<�ܾ.��':m���5�.e��z��$��E+Ƨ����q�LF�*x�o��^��i,iA�O����/�^�}.��a�g��z��˹/ ���BX*�ov��Ոe���_i���$)dtd���|CSV%�G9�y]m�`x8��h��B����B�H�5�K�U�#��9ܘS�̂�uP�.��p=Ns!E�GC�Yy�N���\c�*��͘3WW�u�n�"_��y#����j�k�ӵ"�����P��n�U.	pǦkC=%C{ל��V�m�<~�V<v6��MDl���vϼ�Z}j�xup�VJm��VDk[ܨ��3���6E���=��1�2!����t��{3�`�Mo
۾�yB9;y)��C���y�q1M�<Fw����M�4�Ү�bǽ)��Rے�l������W�17t��1�J��y�lK��l@&�b�udV�s��ܮu	_e����Ao��E���wlt[���nX�j�8�A�&oU��@�=��=0c��*Z�-����-�.jy
Yy,j��m*�;�<�a�����#�����r���*
*!�PG����r�0�H�����uK���؛"p������f��d](�Αp���^��T�����9�̫��n�Ek!l��Y�QV8����!q[���ګ�m�B����,hC���#"��8���!�*2��4��GC�wV���Vq/9i��i��^\
���|��OƢ69҉�m�]C�Ê��ϋ��B����b!�9�cc5J)g��L9Ȯ\PM!6YP+݄(Qbv��r��mՑ��b�+-��F#���Es	ۏP��uNzQ��*�B�X�=�;t�u)�A%�u'�cܭ��u�8����~�F�Xq�+%�7�3c�93�a���J��6)u_�wU��@�#���X[Q36{�����ޡ5��T-�:+�W�M��W-L�Pk���&\]H�@ء,_e>�;z���O5,��(,�>��]5�ϣo����EA|z ���u�U�ɉ��У��/;��S*�P��D��0�B�5�@�B�P�l���W�2��<'�OZ��8�h}�0Ж��*$���Fc���*.�	�]*f�$�/O����u]�ץ�nsT^z7��4xW��n��a=U�|5���[7�j�{[�ġ����=�q����/l��\��U� �IΜR����w���O���쓭���9J�d0\���\���7����wY�@ͷ)TX���bQ�⋝�ާtͺ�: �}#�"xaQ���V$>��V�n%�qJ/wms�ڵ��o���9�!EP���N�4y�G�|'�J��_�tt����Vv2線=1p�b��V滋�l""^	�����C���Ml�&tpdU���f=K���s�u�MȀ%Z�^�E�Y��Ԍ�0ؔ�\�3���Oo��}�?�|�KxΨ�?1�������[�[��Y�dz���!u�^a��y�3�b��*iGW��ED�5nP0h3�FVr�:v�ʝ��}x�!;=�LC9vvS�r���,�m��_,ސp���ҽ��!����x��tW�z[X+/Ç�cghPZ{TF��Vk�5�r���)�!�V@����`�|C98M)��j��;�9|�X�Y\�5gs������OU86O��v���5N/�9Ӫp[����	UB�U�s\sӷp�v��e��/�N1D1��;:��6�z����������l��H�Ҏ�!9�5S��D�c���hɅV3�]�2�.�ݜ�P+�s�3R�cp�����58���c(_��N��^f���;��fA���I�x���Ll��)3�7喻 ����bW#v/����ӾZT����76�=�2A�-�����;7���Q0�0�W(ArQ?0|ςO_��X݅adL�궻����[�FA�����p�sv㙮��.�r/��U�/OD��z���(����[r0�e@�f�]�,�����\�86h�窲������Rૈ�:ʏ�sK�GÃ��G�S���'�u��r��w��\'7�L�Sa3���yS~��H�b=>^�SFcYV�sQ�T
wr���I�<���o��+t��;
*���u�Z �YN�2$�vyQF����]<�җ{�wX���n�<�1����=����$�sʘ^3>��F���]ccng�z"���Uϥ�����N��f2O�:�(Z�{���{a3s(l��}ٷ���Rڎ.�62S�~`����@4�\�sf����a@=�M��[A���oo'�(�؊�|ª��>Ӣ0��7�C��p:#%Zŋ��q[K���Ϗ؄�tP�$ՃϠ��ƾQDsN����5Ӱ/<�溅/�X��"�]���U pa��3�Y�>n� 9�W&G�mT�|��ӭ�p���ʷ�&��K�E]�&�{GnD�h{�%�t�NVo
p��"��H
Y@�f%� �6��t0�vB�gF�;5��F-���sxT�hZ�ү�˥rP`̺w]�P��\x�{�m�����q��㿠*�fwN�ܤ5f�v������+�$a��lS{I�\���#�r3���[�iB�WF9vf��;�tR�v��.�F�׎�0N������uC�%�g���yS9�]<�M�M1Lyu���ȍm�e��zi�˝��eed��E�f�X�\OX�/������<S���o1C��xǔ.���nV��9&QX�ĝ�����H'4��{��}gT�Q�S�0�ϻ{��Z�u�]vn�]�:+�[7��u��F@�z�ft��hH�P�MQ��]�<�#D�-j�f�L٦j��	�<���.�}}�-�ۘ��c�$u]E�� �d�s�cik.vEw�����閞�S��3�8��Y1Md`+=��%��Y���-Ƕ�`naY�JM�w��诬r�Hlj�h5�0K��e��V��V�Ӣ\)�綞aP�aX֕׮��z�<S���Tg��݋B��l����v��<���c��zum2�wRX�`�V�-�+&X��K������2��y ��gCkN�l����ڶ&[��q��,n�q�ӎh��5�!d@�����fn�ǃD��a�� �ُ&�K�Me�� �D첻z�>ʸ㇅m�����_mǪx(�.Z9eG��c��;�hs�hvc2��%k�I�(��&϶C��m�ו�"s/cT>��.�bl>̫����$�o�Q	{5�#t�=�*�.Ί͙�YGxFF���ϭ���
mb�xY�\Z2fL�悵+[b]���]-���|��u+y��ܫ��O�a�u���L*5t#�0�p�+L�-_�S�\��w���7E������vR��L`,�g۴��qgn4��]E�b�q֮w�ƃ��h���7K��s��׶zGT�¨�o9��\��r��'mP��h�L�hZ�vV�d$E�7M��v��r�p�Zi�ܗĎuJ&�M̾�ى���.U�[�7ws7Mp�ձ|��@�����w���=��������W;@[Ac:3��KK�K�Eb�9�L�����W^(g�\z�ՠ9�ڥ������!�J�GCU�g+�4�{�n6*��o����&p|0�+FM�p1����
�b���Ӥ��A�Oc�\�Y�U)UB������F�;���}v:��F����|8,�{��+��M�u�,[�:�����1��YN�a�ٕ�klp
[�y
QU݆%�I O<<�_-yX��wS����ս�����jː���]�&���i*�͛�*s`�o'��vV�2�7��[��Y�+AY�ik�@��k�Ll����0��*�� �B�"��
��f*���ib����� ����fb*��(�j�����J ��3&*Y���`�̂��&�(b ���"�*���j�(�H���"(�`���j
����������B����"��"�(��(�&�(����j�����j*((c3*�f**��(*Ij��������!��h����$��i(����$���*�-�MTALUM4�P�ɦ��fADTSEPRE0�DMF�2h&NfePQUC%F�
���I�6��ppt
���o�9��9wROjdRK���<.'ZX�0��7Ӎ��"WaRWYf�9�x��{2�g�Gr�
+�u�V�F�k��eW~��"���Q~�n��}�/��\��>����(����u��qܜ��m(2���M�ѳ��=��8	�;��o�tv�}5���L���yb�Ҙ�oj9 �Z( @�:��q
��4�\t1��)����t��,���S1*2�K�S�[	k1�US�z$�#0��p�:{�ҩ]4��] �V5��u��ڣ���Z�S���B4(�z�7�<%��u,����檟V/:۝=r����(i���k�VeN��b�Ml���x�/<���GCG�����B�*��"K��q�{��p�z�{����}�u���Y�������U�.�.�O@�b��
�T0�I��ݹ]��cz-�p�L��	��P����:��v��+dU��DR�c�k�O6snz��Enz�KaK�2M��߆ˠ�����2Y�:�e�v �_	��xV��E�_Pԡ�ku������W�x���q`�Z��k�[q�� WM�����/'1q����c��mv�����uYo�I
/�b��Ԉ;Z��M.���J�)j=گ.�f_�İհ�#�w!"��o�hP���Pɻl�#3�r��p�ky#co���ټqN%ý��ϖu-�kI鮒x�GS���3�+Z9h[j-�<�sY�٥o	X�����G����L9Q@�VB3w���5�y��X�7��UU�ټ[Ϩɛ֝�',E���X�:�Q�T�!D�y+(�ec��4MU����o+g�����LUnE��C�8��Э3a3{5`q�0�P}��"D��W{��pow>F}P÷Y��e�_��[񷢩���s�f{�4�+�BVQ�;�8r�k�Z����ލC��Jf2��W�ò��=�C�2���V�Zo�'�>���O�m��{m�����x�o�X8H�o�1��n���WR��U]���i\v�F볘j����pxpgs�D�}b5��q��b3��_')㮵e�P�sɤU�ؒ�8P��{
I�H��s�Cv��<�ʷ�%���N�N�;V]Ǭ.�n@lv)^��3��m�u��i0�+mGSV�N�5@&�߄>Ү6$��6jKKz;9�b��mƳ=O��6��6r��۾|��y߂��v�3�P� ��ѕ�7cI�al�޳K�z�ةw�\�8%\�d��C˪�o�>#²��zl�����F��]3�� �6�9П�b�F 5���ٽ�l��+����8��M�Uۉh�b���Y+8v}�Ċ[m�]���R���HkQ��f�t^����1S���,V�$L0������(�(>��W��X���;�7���h|a��Z֮�.�,���a`^�2S;r�W�{����dݧ���������w���������
%DH֫�t��T6_:�Tc��f�йhz�NaO�D:�5�~�S=������A���D��d2�����౸����2X�6�-p_[h�([�8'\��K �5��.=�^��z�셉�fҒ.�Ѿ�n���?���X8�j�	O˖3έ���*8�a�&��7��k3#�6��1^M�Q�ŉ�8}��ַ������zp,�Ԑ�'�39���ۻW�2���>�a�Sײ�\B�]���=�oV鱎��1�����Ne+	�����F6���7h��![
'eFq�fJZ�g��Z��xl�j��H9���7RȨh2�5�۩aŦ�̢�#�2�9��S�j��KlR�qp�Z{?'�`.���;�oL������Wk�o!��҈B��ޙa�q侻�Fo�%�,r�Ep:����$o�5Ԭ���t�s]�4/"G�%X�t��
��6��On���y\��X;�n��N���s��ȝ�񒳮�gP�2�"��q�����ڹ
�ٌO��q���%�ջ-:�α۫g`q�P�G�{w��}�rU�<��]���t�V�N��W-c���" ʕt/ؼ��W��!ƍ�a�&���Ѡ;)uX���P�tP��Z�Eӹ�^í��ٶ�__��.�lO���P]^%�J���m�4�v�­-�M
[ME��zۦ�U=Vh,TU�K���*'a�w�u�[�1"L�)�Ļ����>W�g��ut�ד�VV��k؏��jr�u�y���<�Ӯ�֑���C%$�s��+X�U{:���![�B/�<$��n�:�^5���$k�t�9>����]cT:���n׳�{�hC�t5��ͦ�X��.���ѹ<��Nn�-ywk!j����U����|��d���f��fs�iy��I�Ղ�3&���W㏪��"%�6^�����������(u�v�0vuf�[H�[g�"�ث<��ܽ��^������(�ܦ��V^K��&���k�tHD�,d�rz�ѱ���8/SE�v�c�f�Jޅ1y>W�D�9�izK�~7�jp]�F���C9�p�7aq����W��C�"���Xk]�g�<�{�`����v��^Q[MM��{ۨ���5�W5���M�&��F�`l�s)[=�Ҙ���Ú2�92q�ve�a�w0�̧a���[������=�p�>�j�h����Ըrs]]gWp��-�j��=T�~��?�n�W�{+`*W[$k�aOF��ث,"p�G݅��66[�ջ-���"dBf������<���	�N }O�-��{��ǒ���G��!ja-`�k�O�&�Z�bi����>�'Ժ�h�l�l��ؽ�
a[�S�T��m_1]C��հ�2;��2���g+��$���hy@{O0�q�;
����������6@�O�٫�vⴃ�X�GZf�;��[�[��-��3�Ѧ�d���p	׺�>5'9�������Jm� ��u��u_Z!QƄ�'��.�e
d�{��y� m�=Id�3;dH�I@�B��a���W��K��U�����m*�:��4۩a���ZM,�G+1o8vL����\�ST��3a�u�U��5�i@�a��b=���h�p���X���Fk�t��U��_�j��+6� �g]�#$f�)��-���k,R
�[�:Eb��o���������de3��mњ����pO)���2{��>�O^�w���*x��Flo%04�栮�Ā��͉>�g��ш�/��J6�;�j���\��R�\�ݣ~��A�M��|2k��k2F�O�b��[y��D�e�ѷ��FWd�bﲽ��҃Mk��u�y�'�:͗�z!��qZ��xg2�������M��a�̧m��k���X�R��3�Z�k�Upw5j����h��O�j�4�\bu0��Mpx�nf�jq��U���j����5�_Y���eʒ�l�g+���;قGYq�����NQ�H�!�=����7+8���Eٺ�v�u�I�l&q���5�V�I�X0=w�Ժ�nZ��G#�z��[pk��C਩���;�}���l�&�p���li�܎������"���j�8<�`(���"l�����}.�@մ\V1�	tm�@���vn�<��	�Vli8K�8P�/�p�Yy�M7��VL4�{��pε�-�b�6�zv��N��@#p�luE��}T�Y�l-��Pk2[f��M��ְ]���Ԃ�<�!N]l�<q��y]�۽
����
j6���e�����-j;����f�u'�\k��#��_(��ȞPF�r��ګ��ͻ�Xn��d���(DKϦq[B�yoQWĆR��}!�@�"[����.�k����2-\�襹��b*��1+/�'XE,rQhb>��W��UGU��G���f��[���k�!�ڹ�'j�3���pI��O�b"N�*�j�"�ܬqұgwn�H�׳��䂧z྿6�r��'�$
�;/M��yf\�2;�v�x�3�vd��s��T�}�l�$��%�2d��ُ����Ԝ��T� �G:鍐���Q�=7�̊�;6�o��\׵�/�f�`{H���P��f�T"\�b펡����FU��9�%�UcNp�p���ʌ�Rz�.�šcN>�̴䋽�{�4�76�;�����l��҂!�J�1�#,1�nI�v�YC1�7�M��X�n��ec����3_��?���g42xc3�Ji�����`�A�L�丢im;o3�o���a���a�w��TN����$Sy��*�A�i�b���6��,fD�b�*v��n��h^G��8鎽�����p'5��
����o%Nk1�SoQh:n��f�N���ؒWFe��A�7nFw#�r��h�bh�`�u��m��[�jܴý�@B�=��ǖ��N�fq�}z+o���FFoQBEj m�5�w7�}[�Iɗ���xh�6�g��E��ᙅ�8na��%�Ѯ�]W�V�7}�E�Z�*gk%���W7�=A�Z��w{z]��%(#o��\$CB���ub26�w\a�V�-5P�ٕ�~�7ƹ�:��zq��3Ղn�0S��؜��}k4-�F%#�J�H�˰�s|m��C%7Hr��b��
�5]��V��I����c�{�^�Y�*�l˭-��]�\w�e@�a�lN�\�XBGA�Yb����eU�.�J�[*��f�X��,���CJ�	�q��{f���7.�$2���}m,Һ/Zy|��~���^��p�mu�Q��n{�`�"�U{e�Ú�s�-�δ�IV�NZ}��B�
)c���ڡp�\}#3��ՊN޶�Gxj�]`6���"��םW�}qw�#T%��H��:2{�FH�䎽�{�=q+]>�Ά(�E��Ē�%C�ъ�I�^�g��1/��v���h㼃�Xꧮ�X�jj#J`k�q����Xk�]N�7�f7��wj�'L��jouK�}X�"��à�1C����]��֓]Q807ƃ���\�Ɗ[��镜��}v�e �;�uٔ�6�YY��I�1�Ty.�t�I���������gSc�1��T�kϷƫ���|��{�a㼖�ˁ��H{�++\�h���A��-j<^�F��Ucl�-���.J�R��c�(INV�_ź|��4;Hi���gJ���{�t}S��˛�iwv��v����/���7S;ŕ���3�u��#=�u���,E<ܔ�Y�6ډ!�
"p�~<�%��4�in�ڷY�e(��J
�y �1�F����W�F���|�݅��4�{ZM�C�H1��Ne��s1ǘ�B��P�0�v�nHA�&�FR�
��ھ�o�yY�,k�uk���ucQ�V�����p��҂詾]*#�sv�5\Ҍ轇�ٮ��Ut��6�U��c��^m԰�7�s�޹�8{�S����o<��1�k�4og�Z�j��e;������]��\,}z��jl��3!�Kp/;��s��tx:7��:B{����&(�hj�q!y|ڭ�9�#�%������d�ï��ԟY9
���˅w���暪�+�8$�FO���=�C�Z幧�K	���q�/s�s��OP�w��l&�<�F�$�h��O�����D_f:S�kD@;��u8��a6Y���X�[��\�\�8������;�JjT'`B�;����#(�(��/���5�y[P�HXtdee����#�Sk&��c��I������Ǟ�/.AY���y⨯��v�+��5��1Qo6	e�d[5���W@�{�D����vl�k��L�O��Վ�t��q�˽���}��+��y��ʱcnO��.��x����Z�-��r[�o1u�W��IY�����7��Ae��)�4�(�k�h1P�bFu�l�B��l�μ썇ܴ�}��Z5m�����7�ʎ9ܨ�&TT�m:���HHj��s�X���hgv)�vL5�)	͍��C��+�
�i���Mユ��8b�e�;��8�M���ƭ�,n�a�Q��xvb��s��MS�x�咑 �����r|��N[il��ꙡ�5/{�i:_��B��;�BC��3B�m�7���vgs�\ࣔ)�8�:�	R�Ow�A�����)�`d*�Ehg,P\��*�d���&v��y��
��k�۔/{Z5`c��~�I����&Q�i�]c��tQ�#%�T�f��R�U�o�$K��:p:k)��\5C��a��%jKȣ+ Ʀ�5��ib���*Wֶ�-呃�2��lN��qV�t�Lfr+��r�YC��r�g����	��"�n���w*X��a�zl[.2����n�f&��[�wv�[�2��W	�2=�gtSq3�X�t�7����Y�e4�ba}����R=o1�Xw�
T��wSt\H�8���7:�k����ʐr�}Aӱ��#���F�+��(�ӎ�n,��Dtv�@��MҳpWn,;G]జ��#�;�R�g7*ޑ��%��s�=#�7����=��yOq0� R&@% �v�V﫣���VzZt#��{y%��6��#��ţÇ@�)Hc����_^L4"C�N���)��K�ѱ׵�ŭ��$/�mN��}�TǊ[�OU��$�������+��\�]�N.G�ާ��86�6�k"�c���oJ��\�g��b뤇_�X���Z����K_jαZ����2��]3�� �wۓ�֦��=Yk��+�1�ToL=�%f���.I*�γRP��Rڴ�꼜a�BY�֧�d�;-�B��ֻb���n��"M&�h{;):�/�r���7 ���x����0��NKN�\���?�]�!���՗�Ev����� �qW��N�ʲ�`����2ćr�����ħ}ƹ�n���z{0��
�؞]��kO��F1��_�ݫ��׆�UK����]5/Y�yR��,ݜn*�BwB�h[�r� ���[��9��a�K�=���b�C�+�[�5�-�W@��/��:;.GԶ������x��wM���l\�ˮ���'�ˤ���j#�0r��˔���K�����&�j%"j�c	hH��
��������#�&QIAUDMLBU4�T�SEE���EE%UM5L�PZ�)����������� ʃPc	M�*���j���*����`5`DCHUT���E%%4�dAQIT�P�LP�M-1CEDTE�TDQIE9C4���SCK0��1d4�f$E%SSAUJL�feY���R�QT�CE�#KT��d�R�fIB�PP�Y!Y�C��+�vmء��2�9�VUc�T�Ĭ��E�,268���{���2����oi��^t���{�!{Gp�n�ز.yg#=�܌��x����~��rn|2k�a�k2t3� �[To%��}��OB�&����]��t��A��1A7�v�:�`_X�w]�\�"�k�L(li>����>�Y^��gs�fS���du�7LwI1g��n-�Ԭ,=�&�D�xF�ۥgS|-��)͗�7����:�5��Պ�`�����k�&�#��
 N��l�e\F�<�j'��S͈ޫ�s@�RZ��;�-:�<���Y� ���dN:��c0�����#^w(��1�WS{�0Sm:���.Ӽ�'�nf�U�C��P����J��-�'��m�w��yMk�5I�w���&#���(&�ئ3Cj!�3YB}IA|��]V)[��,}���H�%<X�>�z�e�iuq�;��K	Q,��m�%��*}��oQ��̈��L����1V�[�\:�YW��ު�RL��kM�q��4�ٚ[��e�{��\��Q�x=�B��+Rm#ԯt��7_w3!]�J�_pV���%�^�)�X���z��n�̩�è��&��1w	�ɭ^C��pΊզsBޕ'yv�Y�_�*"�����d4��2�P��Nɜ]
�/Y�A�F;�_�Ӻ/�	y}i�K�
$!��#Z�8Xݪ��PC��ݗ5.}p�-u�\�`v��[���r18b�t^Unc7����t�<��&B�NO^�~H*w�p_[h�Bۋ�̻�w��U4u��V*'�o���ۓw���;w�b�p[Cܽ}[�]�Rq����~l�
o�"$�sY�k3#�ͦŵ�u��"�M��-��5w�n#56�B��Y�Qþ�RF�xc�9����ڼ̦��p�;���N�B$s�V���:�8�	��a�ٜ�W�7-:\b�䑼�����+)��_k��Ӱ_m'Kw]i=�y8<#C��]�2�S���PU��L/�1���i�n��;7�=y���N* �u�]�5�����:3�]$�O{'l�H;Q��y�77f�D �}����Vv�Me�Ua�G�m��F�{�t:7Ws��Ѯ=ձ������:v������]�g�tWe��c٠�2�N�E�(P�[�k�q�NZ���n�[��0rvvҸI���^�]�+�-��-޵n�i�<�K�7T��p#bN�|5-S���}F��P�|�ð�^��t�W�SM�cqJ����O3����Ů{��C�*ǣb}�r}��4���a]SW�����݌ӎ��e7�i��;�~֣�=�W�cc;�Ђ�	CY�i*�=�������t�;7KUj�޺m$[*��eb%p��/o@ia�
�3�ES��swKk��^ؼ�����ig��ut��{��V�Rqq|p��ٹu}����t\�GMc�/���4��ql�rx%Mr�d�Z"��j2VHa���	��rb����H*�P��mT�V�����]1��Jq|+����x(��'�X#$Ss״��;w�x1�V���wx���{Ϫ&��`��;rlֳ'�<1Ix�˵=}�=��[6�S��
�\�ǲ��\[-�t��S_�����;9\>�%��[�c��^�T	(Ob�ܬJ���Kz�&��kLN�u��b��������yp�YKrP�E�G��2:T�}L�E2���تG��������j.�=��f��ε�����M�kM�ߥ!�Oj�~����]�/y�NW��N�5��Ό����*ۻ)7Xm[�k*��<4��3f�Uʵ��Z�;�M�Sv�S����Nskl�W�����a���v]Z�n��|I�x�\�X�s���l���S�z3�Ä���AgTݽT�:Z���d�a:$��j�}	���]Zu��vxgw���v���7`F��c��9fTD��ָt�����I��3RH��lI�Hn1�ʻ
"���GVU��cY�ܲs*�%s��N�m5bZ�bi���7�J�N�f\�U)�k+Mh8�B�5��������+���	�v7��lp��9�����q�����Ŝ;fS��F�f��j����J�펯=Vi�R�*ۋŧ.�}�<���q'
����ps�N�F��r]MR���
}��*v&�������*��6�u��9<]t���tƱ�կxG`l�ԥ�"��.:��lVL~gG���6e%�����>�3V`�ٛ��;o�+��݉6��:V��N�'j������ �U��gz�H����}�z��;�6X��L�rBU�Y`r�0��\�ʁ:@�U��p\9�iQ�k9C܌��Ut1Y��*���ę�t,rAB�k|GMb��m�G�F���UnL���mL6ư뭵T���X��#'�N����d:{�fM:��b�\0���N��}~l&�7'u�<>ъ纹#�rS�]�f�}p�?l�Sw���Sm97��ΰֳ0�8�Dw颙�'4)��t�Ya����vo���v����k��n�ךb�ޘo$ճ��5�K�!��l�s)N=�������:�)�wCF���S�/Ds�Ņp����8�	ި���0��p�4�\b[Xz�mu>���ѻѦۘ�������OWvw��FpxF�%���r"c!Ϸ�Xd���w,��p�%�-�j���C����*�bHy�YF*+���û7��uBfG�HsW}m�[��{����I��q䂳��[A0��t:[�2U�7��-=f��Cr�ەf�%#��Xش����FC#�C$.r��%�ԹJ��[*�z�P4uZ�}}}e�lu�0K�"�]el��~�+�|'~��~]~o6Kz�|�t#�>��;�}���/�Z�K�,�.���	~<)�^�F�)7��ְ_j:���c���P�r�cw7������ƍ�P,O�(;|�e.��o��JK���/��D劾ȌV�F�?��l�ލ�w����@�P}�ܖ�Uv��@EMѮ�Oi;�x���=��QՊ�� ��z����RZV��y,W�t���Ӻ��]s��X�+����<�a�A�
$!��֕�H�].��6��I��}Y	5�N�\�`�S=�ŉ�nA8��:�D��f�mJ��id�u�H���$;�ms�-ۜj_�Q��FTe`<�=������J�`�[rE��6s�a�XM�"����]��R�K6�ُ�c��s��씹>�²�䗷�'��eJ��2�t@RJ�$���D�V&�]rf�a�f�h����O[MnD>�Ё��B��yx9o�#���p�Mj泊RV�v����5M����]b3zН@�\n!�W����aw+�S����4�Ωu�]��oj���dK���K�{����=�gU�+���pm�a�s�5Τ����R�8}�O!%Ү���V]�<������9�e�A���a�c�'�X���n3
�WwZ�c�6핃/14Nv�|���x�����n��|Mȟpyu�j̬��?M���6 ��׫���݇����u;7<���hFK����;OTb�ൎ�!8�
w�<�݅+�im�%�j���1�$���b�YʮމJ���ǭlO��"C}@&�>�G����i�:���:w���{�P�|�W-c�}�X��rĠ��B}IAmryɇVӠ�nTµʧn���������𡑾�r����Q�b
�H_j�UUm$*⻷X[mU�w��Ҡ�ʠ�Y��QV )����xR̝=��gib	��d�'��er]MrҺ�OZ{k����q�V�Z�ʋ����4��~�=�&�h�z� �tژ��F���LuC��:�Re��N��MʏF���W�̱�ѽt5��][wp4�Gi��Gu�1r����z�뽺W�}B��LJ����W��J�Gܙ ���0��n_U�5�:�M]]./��z�=��h��Fs�6Ec��|�.ՎiZt�{8Q���Y3�B٧9}�(#T%��A�
$p�D��D9�b�6�� ��T:��@k��{}�Z|�Lզ:1�N	�3~N�Ϥ�+e7=[H�6#������ʱw{�LiKb{[fBۉ��k2x"}����e%S���������/�̿cv��Sm[��-�ɠ9�]I<1n,w&�aYW��Vk6ȻyC2�;�4�+��P��:�k�$��0�m����5]|
�җ,0��e+۾����á}�����Y���ll�\M �MM�F��%h���'�M����-�=T�=o�����Ƞ�P�BU>������כvG��n�#�Z�ǽe�Uӌ�hM�6�P��&O}=�x�5$��ؒ7�6g"�)�u����pS�fv�Bt�m��j���
��ؗʖ�e��_] �S��A;�����k�Kj`�y��Víh�dΊ|W=�8%2���h��Õ��D�W�JR��t�9���Zp�E����co��q����p�'5=�Q�qvĮz�:m5cp�]4hWW��9�߅NP��jg�c���چጶ��n����+qts}I���ƃ��&'���Z��K���Ǝ�	��J����}mU���Ŵ�}���0� �b��k���b���b:F�Q����ѱ�ܬ��X�����9���a_B�vج�~j�յ ���X��P'O�P/���sDJ�WW\�W�=q����(�i�G3�'Z,r

�`H�莬G-�9��w��-_n�����_�\�<X��	#��8+�ݟ���h'BK�����v���"�}4���;��lhMv�đ�����=���v�c)����Ǥ��U�)���JT5B܄�-5���bʚ�Rɨ��rؤ�Ɠ�4�g+7��k(�l�ͤ����n;����l��ܟA�dˤ<�7hSv9��Y��1�p��#ide���hZ�rhd�C6yX�����k��$�o�c��&��,pJC�Mڼ|�e�^��[�Gd8'$ś�8L�˯I�1l������[�|���ew�irpǘENow2C�Y	��;#;�Z{�?`D�l�̥g�Y@vSc���
���^�e^'o1kݻ继�]Z�i�XO���Qn���)�LUk�26/�5gTub�$�L�*�`���n�%^D���T�:����|�Ly�f��'X��?U���[M�i�<���C6$��lc�U�d�5��5�뗣����z[u�R�[y�[�o����.��[�Us+���wvO�T0�dH�@�4�6�;��M�u5cX�C���M�Kt�es��.�lp޹a�x�IF�3ݓ�ϩ�����L�U��:��f�"st�ޣ�7Eߣb{���PJeؔ���9k��zh�-�׽L�:���T����bl�����OU����A{x�iQ;UG�!u�g
�]��J�42�������Һ�O�<�����A(�u_��a&�tz�^y��@ZCK7�hn��7��p��J�^�7�i�t5|&�;�݁'���V��SSO}�6l�6��sGVjǃ��T�]�pp�E����i�v���Mj�N�oAT/+,7�e�_q�p�|/�+i�,}�X�.XOu#X<8:�`9Еf��~刪�w�	���ljs�j�%��<��B�]����C<$�ͬ�ܾ\���B�Q�r���3|ؐ��%ܖʫ�+�Nj�a
������s�^����t>S�\��G"������ҝV9�cVI픰]
р��愠���g����N�k5�j!��o�V�bF���=���a�F}�n[}|��7�!�X���tę���$()�+`�+wu)Z�����w�"�U�q�2[�{us��qU+	����U�<��1징����Q����o��=�m��^h6�%)���p	]��5n�v�x�����H�[��ս!{�@���-w�Uq��j�Yt��s,��$�D+����Gp*}PE��r*�]^�%�#]�p��o,�W~�O<[�ɌR��J9`�	��u6�e���\��^�a�Ui��	��}]+0*�, �^��n��փ�Pr\Q
][�\����j�1o	0��ōE%�N�N�΅�7+�����z^���~[é���fj�g���͜�%�֣S&C81�-)#��t-%X��Ȍ�(K�� ��i��'P�@Ma;�,���}t�Ln�Q�,|�y����X#��:Pf�sl	��[�i��V�S_k��En�{)�����u������
��g_7�R�����wyDڜ���&ʸ�޻2]��L��S�1]��]0L��"�z��E�A�[��PV8�Ұw@7*�9ʹ�����Q`�yM��b����]
dw�����Wt%t��*%6�H@s�H}/��!7x��t�g�z��c�b��)�I��8@y^��GfM�`��a2G�>[���\N
�mؾ��(�9=ET�����P����>�yѕ�o����U�gbޫ����!��]����3��+�����5;A
/o�T���zqG��ܲY�ܞ5՘�ym6����W��~��%rXy�����u���׮�u�\n%�^��=]Z�e���U�].��e�,��6�1J��Eb��|.��M@��:Wu{Y�;I4e[�ĝ�¥nm��)i�:�*�Aϴ�߮���^K<<M�@��U��˜�U|.��}Q�q�mf�7b�t��3�f���/e�F���U�SVn�s�Z�))[�@R���n���f���������Il��F���d�fq���b����c�#K{U�)v3�Un�̒3Q[���%f�|�x�1�] J�.�yL_Z̾����m�Èt�N��3���@�Ա�G��nL�^��#q.'��4��\�p��z�L���&�˫W}�zAO.�-�o�:rՄEU%5�MR�!�R�PSTIMM	AM-#AMddP4dЕQSRQKT41	E%5M4�9�QE���AE%DSE0�ddSQ#���T�Q+AME4��4�NK�LLE%DP�R��dC�RfIC�Pd���CC�@fcMP9�e�f-R�V`SHU"QKHR�D�&B�BY�DT�19!��R)M P��Df9U@ę%5E9���d�R%%HД�~�����|��[[�*;���sS����V��U�Ѳ2�!AU�y:k�㌭��b�q(��a�[J�Awq�Euɾ�V�S���kUP�|�p����<�{w�d^��
{zB��Dv�U󶪆C.2w:�SZ��[�$=q/x6��C�� �uf�B5T�Wb���fJ4g%b�xE�7{H�s�a�X�%G-TVB6�'���4J�n�W�pֳ$pd��D�n��YC1�2��m�ޢ�a����#J���n�]���Zk�I<1�9���o1�<�tf��\/�ů�y�]�����]��ޓ]Q8���z���G�L�L�4�_��:�t����Vf�w�м�����CXZ&��&����^x�Tl����-����:l<�ͦ��n�T�M�J��Z4m��C��Td��yW�
W�[x6Kw�[��n����V��s����ܯG�}��SWM����]����ޛ�+�]d�ɋ�N<��m\��ZgXYW�>a����;�c�b�:Ѫq�g,kc"�i�)_;X�K��è��zP�|˴F���Ћ����O%r�Y���9�բ�L�:V��n�����]F��J�۳g�9S���Q�,Q�{r;��ʣ�Х^��CV�C�(l`�D�J)(�.У�Px�Q:���Y�/��U_��jڄ�kQ���ޗ~����AtX�wT�9��Qk�oWsS|����m�V��ՆҦ�S�Gm*�`@UW��o]��u����,	���h��r���N��/�{��V
�F]�/\S�y��#�c�=���mb66_+���X敧H��}�Rk+�wp��{nq!y|��h4� ��"��D9�H������Ź�\�2�j]�r�䔞�aO&��C��gB�46d�+#$
nBy��i	��E�u�U{H����{ɘ>Mv�١��7���Ξ��y\�Ԉ˳�;��N��xz���ɾ��cn�d�:�C]I��Z�S9�$ԣmE<ݗ��+bo�X��]�l�m ڶ97�1�i�u���|��'&C�lҘ����Ut��hf�f�}�~���u�u�v��aj�;Z���˚�嵏I��N����>~1�Z��Ӌ�G2�f�Sy��y��M6t���I�G�r���H{�v%N�+yP�/�BxN.�疵5��q��^�qL�9�����uN��T���#DNe;�y]����aо�m�wc4誋��Tf�r��x��R��}|M����
"qҳ��6:����M��y�oa��y���֝.�8�Q���[ջ���͉;>
3��<�ak/�B�U�1��-��M�lB-Xm[�ۨx�p$�Y����!�8P���Y��t^�m��=Jt���x:KW�S�6��KZ�G�N�Ue� ��L4}t�ך�u���X�M��l�e'V�ڱ�WcQ�V���Qǲ�K�Η�Lb	�0��g�ʹJ6��ﭪ��w���lu��[�����Kf���tw��~�{zw �v�q�}۞���l�Xu:�\%zg4v��u6���i�ZU"�Kψ�woُ��=;#�P���Ca�q�N?=Nͻ�L�rgб�!b�H��x�C�*HˁB%��DL:q�G=ىT:�Re!���C
�*� �\�����:�Վ�Md��v��T���Ė����˙VV�!�79Bv�v$5w�:�ge��Ƒ�^ޚ��]ܷ]X�a���]Q�[[������nM�&��E���$\�Y��_;���ָ:���2�;�	�3|N��4��d��6������{z_t.L�4����}�ӱ��Ʀ��'=��;1ӕ#n*�vU�P6��v,��Y��ܑ뽴{�hs��n5�2D�em5[�����;��ol�̰���s��뵔3�~ͤV�`I�(�Q6��$�9�P�0ݖ5V��/&�dNe)Ǿk(vSc��·�!�v�å�h�+\N�s9���a%�5��x�I���
"mҿ=�v��f�]��+3z9\�c�=�.a�x��Y�	����������0SU�qU`���κ�؇k�)Zg����\�Kv��~-:v�y4���2"��ŧ�5�=wKnAb��:(K�C��q����-ߵ�m���Jt���;1tk�˄f�}���8�Q>��CC�&�Am�e&�GSV5�v(e ��������ݼ샲�'��͆��>�'u�重LHpk���8�N���'��<'f��\�%���;�ٛ��J~�+�V���WxP�/^D��{�Z�2�a	�c�޻l��GY�nq��� gm:�Q��9��Ld��-���2�t�����A�)(��f�-u>���AR���}2�t�4fξp��<�h�D�#c��%Ĳ%(�]0TK5��+W�f�_;�E�2������f�*"�Sོd4�z�oeZbZO)wS��͊�p���_5�Һ�|�K��	���AD�6smw>���i�K��9�#�V:�����uu��i�<=�ŉ��s��r�9���u8�Y!��>����vC�Sc�[���~���ڠ��e�Q֖��V78$�̑�D��@��Mfx���'��y�q�(�.M3�y��a�������Z̞��M���ywq���-��*�35H�a���}���1I�6��8ts�#C<1��G9&�@{�����ܪ��fe{2���A�S[���I��*����#	S���eaU���%Z�R��].�Z���R[ẇ�/u�;�r�ss��ֶT��vk���x�Z�4��r������N�v�%aO���@雒�����V���w÷��w[����*��V*�o�.�� �A�ͨv��ދi���(�ܻF��PNu:���Y��(_S�w0�v:v�L���|L��%R��Ԗ���
y�T�}�'%d�3�¨/�F ��Sv�v�wz_</_�K*�pѺ���=y�$<<
�����)p���-�w,�i��G'0[]ݪqe��C�Ր��_������&�:�]ZO)�)&�5V#\Z�s�VjƱN��|��X�}�X��7  �W�F�S�=�=#ae�\m�W��@,��z��BZ�wx=�A�/�b{���55:q`|j��ǜ;_�dJ�#m�am�V���i>���Y�J�vgP'ڶn)�&c��p�[ˏ�g:'a#�ܗ�[K�������)y���C�ڠ��vb]r������jF�b��|�}����dcW*�JӧޅP���^��bL�*܅�J�n,9�Iz�FTyOJ�L������N:��r�(��ov�Ż)tZ�[/��J�P�gi�������vx��6�헫P���'b.ܬx���E\6G�뫪��M��d��[������zC ��%���TR���� 	v�Z�����Gu�J�Д�c9)���B:�T�z<��Fxu�����e,�{NV�c��(�~��\��8/�341�rl��d�D���L�-Cv���Kw�uB�fѻ�7nپ�m�c�n��&��Xhk��F�Nɘ�mĻ�-�l4}9�����e6sJ5�&�q�i{�:�Ľ���a�as��%�Q(v`n.ʛuN�e �=�á}�Í���k���Z(+�Y�3��f8;�`(�:W�p��z�.�^���;��ҥ*Go𹓻J����ݞ�|z�bHv}��'v#�GF
���;�NV��d��V��-�$��fĂ7��wl��\�nWn���օu�;��Yմ�Β�����Z�p�N�];��b�!ў������$ �x�O��h�N�SK����GRj�NDAF'�vő�4�W��������bk�d����վ�S�5��-4UuI��K7�N�#;"��p��{��Yz˩ndw���M�K=mι֋V�|�k7yf���ur/�a����� �I�+{N��-$G6��GAp����9���V:�in��h�\�����68v�K JPF�3�ST]}��6��C|��qቡ9�c��,=�5���wB���TN�F��r��ڣn��G�;���s�Md�Ł\�y=�a�i�J�W�Kڠ4����⥹SP4�X�r��Mu��LC��J��77z��c��(��"$ky�5�[���'�қ��]Z�#_���%'k�WX\u���+���n�Yn-�)�c(.�ܫzj���.������{j���c\�B���lLĖ�9���Y�9���=�B2��pf�+��m��m�ݎpX����r�^��#j�v����P�~{Xi�:�Fs�o�YY�ټ�A�s!���Z`�,�v�<cu����b�S��6m�H��f��Wy��[Vb˖Ty�O1�ڡms�ٔ�[��;�kݶ)W���o]zG������w����l\�YO��6���������j�Rul�:Ƣ�-�`��R[}�P���9�.�˘�̃͡mW�䀓iPw��mZ)�^��_T4BZ���Z�궱�ӱ�3;�������b�Y�\�0�
`�_*P!Ͷ� wM[)���=5k�����; ���ݚy8<�z��ċ���-c��o�[�/�=^6{�ь%{%�5NZ};wH��,��f���̥��eE��P�`1H����B��T;
V#Kob[^�)��q9�/Bْ��eWyi�w��$�����P��{m���jE�����Xc���	9�����Ҟ�ջiW��A��b������ƃ;\Kq�5�^�3=uLV[W��%@>S�����}��A.�/�}��6Y�g��ZB��]ֶګ�>�m�u7��=Vh,TEWW��:�/=���{yZ݋�9���Y�u^�|�.�k�u~�Υ���:�)c�=6'��͛�\N������Dt��T6_;\:�W:��U3��b��i�n�֋��w��5BX	��	;��!֩��n�
��p_G�ᒻՇF�Vܹis�hm�xNW|�o��#X	V$��]�Je�:'Jw�'u���BYVןz���C<Gk�,^��[a���5����>U�9o���e�JU��Q�9��&��u��*�2��<J����y���I��CXi���Zz�>��+��m����e��q\�w>�m4tc�89���b2^+�>���n:�q�{ٸ�C���G�����R�iD�z̞��m��ی����b�/;��/�ݳ~ͦŵ�PM��v�Zk�I��H᎝�8���Zr��{w�>�Y���ۼ��f��-��kkv��zM{�3��\ȕJ�7��φ��vp�o/�xk��JWf�Kt_E�=3�pk��k�;���/�D�xF��`�Tl��F ��Sv�b/����=0�౨a!�F���;��3`����'vg�v��o����R1By�u��]�̴����q�bA�C}E	��T�F��̸U�*�v�wto<7E����馯X�X�(j�}�X�#��B��EZ�SUd����Ѿ������{�~�zi|f��.E���ߞ���.�����Q�Q�D�W�����ED�؊�+��TA_�����"�
�Ȋ�+�DTA_�TA\Q{TA_�"�
�aW�����ED��* �������TA_�����)����x�)���9,����������1$}�| �TH��U ��R��H��
	�J(@)UD� E	
��
(
T  lФ�%JED�@�E*�"U
IE) ��b��IJ�J�V�J@k*���"@PP�T���$$����mUR�%Ih4�I)E ��J�PT�ԔB%*TH�#f��*D���UR�UR"�*�PP�E(���Uݺ�PB@+�  �����a���!�-VV�j��@*B`�m�4��B�jS`T6���kjd�ڠ �TP�"�-��RT���   �CMjFeE(эM@m���VUV��`��b�3Z� AV�5@Ͱ�&����P���S@���UR�JAJ��7   c͚3#�&�la���jTe��&VR�5��Kk5�E�4��KQ�(P�B�
,�
(P�СB��n(P�B�� w)U@�K�	AH��[�  3��
(P�B�	���
 	(P��P�B� P�8� �E
�a�@h
a+l(���L�aJ���m�����JV�eR��J�PIRPN   X�T��4��5�����0ƃj�h��$�a�Sf�YJ�)��Pd5��6��!$�*TQ)D�ظ  B��R�b�UT6��-h(�H@T���р�h,KB�6B"��5PV�RT�EIUD 8  �J
��UTN� U@�@��5P�j�UU*ئR�TU)�`UU �(l�%�dD��*��8  Zr���6[T(Ц��#@���ҊU1��U�2VP�$1�iU���b�3#kb0� R�,U�)ZB�1P�R�D����  ��4�Sm�h 6�٪�m��Y@6ڵ�� ڲ�m��D�0f�������@(б,�@5f`-6�A��P�R��R
P  �PCZa�(� ����U5���h��*��b�j���*��fJ5F��T
UP�kCmA�dSZ]�    ��*REM   a   O�*B� 4`4�L"Q4 L��L�SM�56��эO�`��J�� �`  1T�J��� �F@FF�$�PLT�F�i�� m&�`�@3-2U�f3e"�[hJ�	X�I0��r��pH�<N�yO������8j~w���2BI$$��s����ڊ*���nUPS�� +T|�"���VS�����%��Y @[�TXR�,UQq�� U"��UQo�ǝ�)����:����"
��]�Jڍ>�0,򔞘��s�1�((BJ��R��C�~a��ۋ�BoM�]@$wQ��a5�0��lS�� IM,��b�b�OJ��iGyp̡�H�Q+*�#2[//
�c@g6�*�@�beP�D|����jλ�
��JVɬ�.N��;.E �bZ��1�J��v�X5�ʹa
&vE�)�\�[��~:�v�@���VV�-� ȍ-$�7	�k1лW���r\�E�߶SٹD}� 	�hǩ�7�h=�����+36	f���Ŧ� �G2�Ľi�S/#h]5Kvd��-�;f<z07Xme����6ˬrBJ6�[Vl�5�/�wtޤA@U�cp噁�Ҭ�/3�4\x��Wz�"��|͠D��{��ۡL�%�����8��4���k���dP�[��<��q��Vg�%��%�wJ)�9a��� e2sv����Q�i�ü�j�t]�w�P���LU�d���3q����Cm�$��(��������f�ƍ���i���V)�Ö��Ua�������ȵLh�!;\Lչ����p8f
Ѹ�G6ܸna�{%k�=��6��L�znInf_����$؋{ �]J�6��0�)T��v*ԡ�/�bj�F�R�׆bg3Jcv�Q3Pj���㭘�)6Cw���hh���% �ٴ�Tdr��ݛK%���֣�dOK�T���m�X��y��m,��+tB��Tԡ�r�@-�,]�4��T�Z)v�Z˒&�x����y=��(�}��$�Z����Z��~�V]�d�H�y�^Y�d+@��[�*Uٕ�&��V�@�Y׋ut(Yo)i�pa
<v���Uo��C���Ɨn2kwy|j�QXOgҽ�"ѕ��Q�f�e�Vo)ڲ�,��6�j�rr���XD�Y�J��ā�4�����[Pm֜��l�h�E�f��'�麐*��R�ZT���3s7)�[��J�a��tlY�
	�������=�| �݆�K3N�ڄ�ef�޺t]Z��4U�74r��I��U����
n���f�b-�e8DyDe*�xr�a�b��1�,5�iz�`���nD��ͷ[u��҆詪^�t�=.[!��eĮU�ś�=�7#=6�;����v]7Sq�xFm��%S��4b���r��8��8od�WnF0�٪�
���Y]]I�μ�M�$�7ZKTo{�M���.�B&��Y��R�kU�����v;����H)X�i���;m%KB�њ�Ƃ�s^R�*�1����@@e���#��k��Y��S�Y�*Ȅ��_j]K��k� �ҧ�$@*���Q"�^�ÍF��&�v�m]�v��2�eeЎ��j}��ǣ>���XX��h9mm�nn�����f����(�6]lhU���HH��˳�Ĝ� ,��)Bf<4[�/�ڠ�h=�W۹�
ޡ�Z]M�$n�5���xC"���En�8��ܐ,"��+��1Q�e!BŸw2�E
��rk
�#
T�(͸- �^�V��2{.]+$5�J:��K�ތI��4n����R��aɎ핚�˥z�ɒ�*���t�P� -ةi�ԕ��ڬaѭ��٪��(\M֊P�	5^�i�5���$�t;5�$����T����/0�w>��uX!���#09E���W�#r�}$�p��]3����R�,�ք�$�O2�h6��yY,Twl5t�`�N��@sD).)s`�)ˠ�ٽ߮�C2�25aa�Y��R,�N�a70K�����v�Uk$K,��u�`:m!�b�c��!Z���u{��+(�u�kI��R �y���a���)*�����*���H-�Z70Zf���[�%�i/��)=xμ����~V9�,�#�nv�v�Zܔ�7F(odg+N�1�/rA�ur͒�w[dm�2Y7]FޜZoAw���O3�y-u>]�I��(��lV\��`��浖��j�n�e|��kp�,�bOsL���p�W�������˦��5��9��H����ժ��c�ۧ��� 2�ف��������/��G+h�˙��N�YX0�T�u$y���ㄕ˹Z�3Es#���V=��S����dTF��Ʈ�Z;��v�
�46�1+{D՝���	Yj-��t(;	#e�Y5V�K,nj�d]�Ac�7m���t��ʺ�,-8rnI@M�#i$�B��A�ty���٥��J�e��\I�<wI��v��gh�I�jɰ�]�qc�Y����E��ܨ�qV����7i���裚3,kֺ�	��f�j.�'V�m���&�c��S0[Pzws2��v��G@ޝ�C�^��[�e�Y�F�r�,�#3mXD/Q9xw�EՅJ^Pĉ3e�Zi];�y��Z)!�n�=р�����`ޗ�&��Q��n�$���wPͧ1\�kMebx�,��j��j���ph��i��
��xMb��1��F���:�U�i%[b�D5��9e�1��Cz�D�a&�K9�e1��7hm�JF����Ӫ�e9��J@�����
�\0��kA���$Xx4G,�w�'���ýl!��zv����5؆�T1��U�r��h��Zp�v�%u7T�,lޔiҪ��w��kstF�j���3*4^ٷR˂�qVы.@�M�ic�G��t�遬W��:��X���[�lj�9r�
�Wϻ�^�K���q��ѭ�o^=vn�6��
Ҭ�Kl���m�-$2�E���[���kp�P�� � ˭����^R��-��
��e���顱��g0�8�nA@�l���utAZ�*��@��r��N�Uo��+�[3U;�,>4���(}�:�-�4��*�k��k7f�M�g+fadkڵ�,�x�v���7h)5ֹ7D�(<�\���wh��l��*�����0i�^cYY���0h�� Y9���2۹�X�e4\�R�Q@��e.�yŊ���g^�������Q���n�-wS`��[�ڰ��D����Z���ݽJ��@퐤;�D��*��fɟ*B4�Լ������2we���)��KX1qk�(*Ӥ��M*v�;���L�����+Br$�x�$I� ��&��ұ��¯m�;���[��{z�U؉f���U�E������	.�E��tp�z+u]nŹv�U�I���Y��LX����b�N��WtJCL��f����ڴ/�ݍc�	�RN�6^�5V]@�?m��bx)������(�ϻA�}������W#f���/^�1�@v�Mn��aA�4αG>�v����ͧ�5�;H&��h׸k&<�a�9m��lV�S�pb���m�Wɯ�'�8��6+1X�kMn<�M۰�<�j�"��!0�ا��0Ƕ2���*"1	o*�_�8	��3l=4v�4�q���g���j�Ei����/)eC�q^`x�"]�5
n�@Fj�p3v.a��NY�e�^Q����v7�M�pTCa�6U��֞�k�v�-�-�[�m-eM��d�PT�,T��t�n�]�K���T,5�ʹ/�c_en�Q������GQ�tq��JE��XԳ��F�ݺ��R��yXl%���D��z��/��'�;��oMj���kͻ$�v_�Uv��DV�ۆ������՛x�:���n�l�����`WWB��$;�)@lm�;�eC�ׅ��1L�	��[�]z�.�E2m>YWF�i7��/[�������
�j��Ũ�	4�ސ*��MZ����� �@��5�b(0�zsm;�ǩ�8�*ZN^�)!��D�R��E�k//����iq�i*z���b��ض�u2	�y����bI⚌�m:υ���0��������i���nX�B臆lH-�����N����"�e�ZT����&4i�
7{K+o���7�fF^���u�Z��Yj E7��)V7f�r'Q�M�������(	��ޣ�5b�P���(J���ӗ�5c��kzI��
ŭ���n�r�6�tn l}(���#tF<7朶֦W�6^lt�VL ����N��K!��Q�4�B�2�ح�Y!���'۬���d*.͹F,k�q�̛���n�t��6@��*;!M�SI�ɋT�ȥ6�۠ͷL���e�W��&�&19��m-�X�:j�����,X��ź�=]y���h����{yx�+U�T�w*=�p{�ٯe�	�;K.�+���Ǳ]��Mb�H4�P��u�# Q��h�{e$nT�V�n�Q���1�SR;a�i��_I;1��u��%:l��r��%�(�.����7kI�W�6�Q��I��̼Pi�-�ɅV]�j�2������g�%��Z�N�^��aS #&�/L�5�Ϧ%�Y;leAK7��I�M�H��PAX����Ƚ��$@�Mv��m���@���Ŕp]GF��Zj���6�rW��mp6�mi2��^"S�z�[TB=��kr�BƗ@^Ln�"DZN#��M�	[b�q�j�ܗ��@���#M־�ki��]tn��p�l������XU�k��*{X����Ɓ�M����.5:��6�fL���Upź��L��-h�q֙ 4�Qyw�u�����n0n�n<�(+���e'n�4��A	�͇��[C*�-JXM]XӐ��[w���p}z7Ml��,Y8�M��Du��,a�
ͼʳy��7p��w�c��C6~��;�\�!r��OA9 �Tl�2��s3n��
:��jדKt������G+e�C�̸n^��"�Ml#����K{���>�m�&
���Ոsp�/P�t�%�wj�5w�V,�k5U2��.�]���1��kU\q�kb�j�*Ջi�'v�tcd���P8ƍ.W��oKSl��DB�Hv�37�r��,e��*Z��9/����j���2��V��gɼ�5���bå�:^a:n)��cm`��@�bJ;�f�NGMՑyL4�%I�]G��^�HQ��J�ӣK	ϲ�sE��pQt�[NG����Uڻ����f=Dnk�Y�1 ��@k2M�V�6ٙV8]�]�t8,��D����5��4��n�Ƭ�5��*Kp:X��	˫���F�eL�����������3mb&�X�Z]���u�V����u�}YE��m�q��8�=���� Ҋ��Xf5B!�2Ӽ�4�t�/6�L6��l�T�}+�J�&�0�F���z(;�"�V��P�L��䲍��֩[�T[�h�HU�4q� =	��׋(�X�]���#o�U�w:�a�,�F����h��J�r
�1��a5 b׷�(�c!f�Ԯ�.�F��xȴ�ݖq\Ѵ���x6Fu����*��i=H��6ZH[�z���b�b����wfb���݀�GW۴��Z������諵�2��PU�2�Y� �zUX�.�Hi�ү8��G��]̝w[���Ę٠�����m��e:�^��-Ċ��捐N�m�ļgh+:�]�uJż�,R�72�F�!Z��m@��ڠ���m��S_h�4�������6ZT4˒D�`�Q��.<�DDů�ӂ��N�8��w/E@��v$��E;x;�`��RT�����\�44Z�N�N#�Z� ��2�9[��CK�T�ͬ���V*�v&�۽��ӈ̗Ur�;���.fڤ5���VŃV��@��H����A�1]i�HiW����՜M1x�����Ӻ����=�&�Ζon�v�;J�J��N��C�R�N]K�S)iͺ-��t����wXl���km�\�����WO*�@�1Ձd̰$�,�U�����-Q����%b��ۺJ:�s�<�u;x[
�������ݥ�N�wN�mcwl4%� :{qm�{_�i����f���6��8%�ǂC�Y߈yd�+.�*������)�wb�h��$����r�q@V��2���`B�#0h���z�����^��M�̤�L�B�7��.�n������EP9W����!��+�Z���i,!ദ�?c;�B`O���+�V��(Ғ:�i"Q�`�gi�&�9S:2-Y��$�q
�I[2\d�Eeg�յ�*%J�kp���a/8)�4�'J�J���K4Rx���#MTKA�{w�B*t5f���!�����Qm�8����״�LvY�"C*�c�6v	�/&Z��øQtVH`�)Q�'W��p� :v��e����x�lk���Cp�F��O`o*iћV�>�B�h�c�ˢ�`;��|���U�R��ڼ��']e���P`)^�Z�n� 𼧻�wYMQH�7Z�+2-{�V3��2��
p6�vaEbMoڌ������n���4�D�ā��-k�?��ya#K^��h��g#0��n0%
��=�����iyBa�Ol!D�Zt�D�l9Yaḓ���Ex7`���^ܰSa£߶F�Y35Zv�5�%t�J-Q���*�ː���:�����=݈�ss/Xuz�Vڬ.F�m�5{w���	_�5	n,:�
�{��i\W�K$�4��&EE�$�w`J��B�ܧ{9Rb���"���V�5��ƽ�)kӧUU�'��@��d�(�����iM�͍�>1Q7f��b�O�r��iՑ��u�V��������*��!�`�С!�*7��p}�12n�^Q� �f#�Ur�,�/@Ų<����A̭�5�V�Xz�-eX��V+f����rJf�a��G�~�珷za��5�/ �y�_��P٬��T��m�Ԏ4��D�B�G Ylʜ�cp�d��.��}s9M16��ޮ�ʲ�{;����p����mph��w�чw5��1�Uc�()Nɸ����Ev�*f<o�wrZwZ�aL�53�՝�5|�M��p���AH���T�3O���^�įL��=��IZ��7PۻI�}�g�*c����W(�Z+k69�
+�s��v��K����s-cwM�MyR� L���tfF�����Or�-��F��TpU�7wC�Y|n��x�k�s���E��{B]��eB�-�k��m�:�m('f�QGs艟^�]״"��"8�K�w.��چf*��ݒ���К�;5y��s�׻�Ƹ��u�N��h���t����oS��pO��E󈼝�_iy��%�أkrT�Z���]u�l�J��d.`���\=���s*^�,Cy��L%g1v�ޮ�#s�ee�h���2�Jh�=d�����$�
ٸ��\�3b�[-�W}Ջ����ޫ̸l2P;��!�Vb��f��j���T�Hr�-R���I|�}�;�0�0e�{�*�]��z�E�*��%{��3�Y��=��e�Q��}{LE�q���Uv��7}�zѹ�%��͝�A�<5Y�N}}-=��Z�0i��'������;4r+d�;@�	-�3Z�G���뒭|q�ö���@��w�3�sPk�Ɩ2��bf�[�>5�Z�~�r�;A�
�R�����Q�,�Ʋ������}��z���T����2h
�A�3d�˻�(�i�y`����*��V��˦Wp�r�2@S�E%�^ź��V\M!�Owf��7WA��a��1�nb7�c�ͥ��[)���u��z!�zV�ѽD�je�H4��<��������{�1��J�Ȁ�WT��`��tI;6�۔G)`�];Rz'QnA%�O̓6vbaa�����!���8+�����7����Z���ճ+[��r�X��Wz�.���E�f&t���ogy��d͈̚��K�T��l�.}�L�ɥQ|�>&�m�>{V�M��f�vRZ��+H����2V����Yw�����j>�՝8f8�-�/!��G��m���LSzBu�a��F)lW*�#t���c��4�iEմ%�T���-�T7��u�qWL;������8��f�N��{g1nS�k��[t���Sl���ʕ��D�9�:�3@�j!O{��Vk� P�ֻ��Eǲ[�8<8t�pq����S�4$s`��am�-EwPq�mP:zT�J˶�[n��K�R�w'7V��v#�-;���"Z��w�+>DQ��v��8�[+�^r�b�ܸb;��v�536F�C9w/qq�pu_mo�
�q�%,Vp
���4�L���yk3pQl�Y�D�T2ED;d>�uȪ{N�ww��]�)��0
5w��0�:urŦ.��=w<m�VE�\l���6i�ކg9[���%NL�%�]�ӯ�X3��Q=� bfAIV�y݂��U���T�J�	Eeu���}Ehcf������CGtz�4���﷈�Q/U���+Ǵ�)��q�,f�k{����օ
V���k�f�L�9C��a����]�)�Z��/���ۉ�:���:�\�!�\/9:O-��Ǫ�� U�E��!=��߱Еb��P�{/z����pP�ʮ�1]Z$�֝�u�vW	#@�x�4�=��u��������v�<�䣶Mk����<���]�bf�m�O��xw����ѫ<,��J0Je<ja���-K��Q�݇��~ȼfؗ��ۼ�>�O4��}����>�y@���<����<�c$�y�v��.�蕜��1������me��,e��ָ��j�I�-���H�ά������& �Yy��t*HÐ�e_1S{h�s)�W�	7�Y�4�|�T��l[5�j�5��p���h�F���;���b� v��ȼ���He�������qf���$�z*̡���`�"ɸ����(*K>����K�X2Y�FC5�����L���K9_C�@c����;�LY���L�Y�sv7{e�Q�&X�SJT�_��ۤ�
:�[v )N��,���w�Ҏj3c�80DP<�;��.c�E���R�.%�o,�u�w�WYT7Zj�i��;�\�2���OW\����
��b���|��MPR����o�k@��N��,[Hu$6�.o�Ю�1�X3�k��h;���)�>�ZJO�}����v4�;��f0�)e)1Mʵ���\��Rԃ/5���MH[�F�̝4���U��f�lKP}z��~�5��N�p�Y̥���a���=Qm��Ʀ�ݓ��*[�Q���Z�HVV5�ժ��,��]��ø�'�Z���=��v���m��|H�k/0�Y�J��Q��Jc
sCv0�s!�Y��mNә��w+uؕ�	����t�}�I�]|��}�a.�U3�8���̲*�r�&�$�=�7>EƬ V
�����iݺkA�|�_�0��#ݪ��K5ʳF���H�̒�Q]JL�g�&85�d��g�Jֲ��ct4V3L�*f^h�� I��ܩ#]=�!)$w��3�����v�P;kk�(֫���1�Ai[|�r�B��g���xf�X�5�WfV�6�CQ�I��W���"��k�z�qɿu�c1��*��W����yL�7D��Zk���e8x��f�A��T��y�\,�����Vы��PV�����W0ꜫp^[�WaS��؀WW�ǩ�	7S�ňG;n8x��ghW���ܰN�&T�F��J@*U�M��i<ɡ���y��a�Z챒���z7
��CU$S��Mee77�N3z�]�n���z;��˩��w-R}&��ޭ��l`w��ݞ [��CCāpՈ0И��3c)<��Q_¬�Ok/��j�c!�4�/ 3����ǜ��Z���D90�r�;��f�S
�K
�}��݄;��h]
%��XMl �D�5���f	�
����r��Z	��7���]x
��}���N'����K-���0�n͈Tu6���; C�Q�#�s��W ��[s,_8������Z�}Ң���>'�2W8���{�<U�d�l���+��O��C����<�-�՗�H��T�I����4�
�2�'�e��t��6�(�p��h;+НmZ�J�t�\2f �uo2��U���4A�;�[��*ӏ1��>�ג�=����(��U$Tb�I�E�4v�J�����+�l�_��QZF:��)�j6�Rŭ�n�&��ȭ��Y7��3���Z!�V�7���]]Yǁ��^v�Q$��F��h���e�*빸���d�.9�Li�i+n�郰�=n>�w�����o�Aq+�lU�.���L4��]g	���L��s�����6=y��1��vz+D�]W�D��=�ZVfKTZǋ�[%����VVaM1�����ӛ���U�"s���{���r�����;m���$��YL���^
#���7J�.��sl<Z_�R��nf\}�s�u2o/�)��+3K<b�h���4�2�CHJ��V�*��;Q�(�ȩ7]c�k�n�P��$M��ᬃ�>��A���r�t�7u:��D��;<�ٛ;�kx4���\�~�JVR����e
��2�ʀ�1����ZXSX9pvaJ���:���,n[Y����=�dr)"���eK�B��W�Z�D��W+�û�F�۰�����hHU(�@M���8�'~Z3���T�ٽ׽��'sw������V-_$�;�u��6-z��4B�)#Ϳ��
�a�- �$�\R���opu.�BPC��*�efG�e5cvk���y�ڎ�ՠ	�("�S��lٚ��0Q	@:��s1<��]%u���ui��K;�t	�Q���|󰱺s`�y����+a(^Y

M<}#A ��Zv:�gd�]�����;hW�X�QZ�룾f2����X)W\��2��2��<jM�ev=���&�R�b�Cdy8k�s1A�N�Ѽ��o��c�먻�2�;-��qx��[�o�Ƀ�6�X-���Srp�z����y�]�5(�bl�I�.���'��ѐ%�G��'����Vs�xDw�S�{0��-Z�#NL�g֖�<n.����������WgmU��1�26��6��ܴC�&b��P�k��܌+�tf��b�Q��;כ���iǄҺ���{Q�l���^���j��os���6�1}q�d)Gj��
�<��ս���7*�˭�q���NM�b���is"�B�1���g:�5�Kc��']�#��kQif�gM탂s�Tc�W��[�����u�D���
=�Gn�P����s�[���k���4�r'x݋;�,�fh�;dr�,{��;�DZ�R��_3��u��`���JUck��$rd���]9�E3�ym�(��q|�Gr��er�k�S<��qb���FΎ\��eP�P���g�W�#��aE|kke�Rf]݅t���d��[�E��R��L������2`��ѭfn��+��4o����$����R
�A���3K{8��&*H yG(Eϝ�<��)���c��t�j Igxa"�wt�jL�Ŷ棴)f��o�O[u�v�]�m���ᓬ�o#lU��3&�(�{ʝ�s^^�`V��WV��⣝���FB2�k�YBpޛ���|xT�4'A��b��35!ë�FP��[���@�L���6�ɛ��2�^ޝle *�o���@���G{'\���l'ʎJ5S���"�t�����g�B����oT(����7�>�kc�/7�P�\.���v!;w,�D0+4����[�|%� X����P��l9�*<��uu��F��.��O�s�6��M��.n_u�YH�-4Vz��/%k��-cM���4��|�Ԥy9H۱ō&�mcɒ�,v��6�r�\�&��:�jN�!>9��Zo<.�X��Y��b����{l�˝.G|�mZ�Z�5+	�:-O(^	���ٔ��C�m*;��S��R�	G'
�hGutPvhV��3�-|EAJ��g�=���wݧ� +4f��B�1]���>̜;�r�\��"��r�а���bU[l''M'τ�KXΫ���SRڠ�!V9��t[�1��u.��%.�W�,X�P�¶s�'N���ָ�\��Fl�yn�N�y������Ȣ���(ռ\�0�vG"�v�����dcieK��B.�-�:���$�|�C"��qeo�\ɥ�v���Y �m2%������ʭ~��cd�;4����f�h.�Yq�R��Ed/�>&y#|NT.�r�u��9�ͻ���(��ʘ_��Җ_vX3k�r��=Ji�SU���b��Θ�~K��)���t��LU�c�}2q�,�:�o#�Z�u��m^i�N�9X�Q�׀	>�d�J���s���2�jN�x� {:�4��������֢��N�r�R��:��}�і&��
���Y*b�̓�#�d�-.��b��҅��}c��=��L��w��[�T.�G,k;�&^�M"[�:�UIuZ����/�2B���ǭ�7m��FS���
�_lF�+�J���P�BCהR��n��t���]43�
�M7w�9i2��]ms��:(�JC:��F�ӂ�[���<�)v�Yj�*yS)2D�I�vFK��s�7UZ^.�rp�,6��߉�wO�ĩ�_�u�n,b�T�	u	�+˥}h��j�H�^)d]�yJ�C��uej¸_s8�=kFGrM+9�q����Z7q@�ٹ�nX�^dGO�PT6�\���;e�H.�mwhj��SX��[�P��ۡ��K��2��Ȋ�-x�Z����u�-�}n����˷��t��`V T�xwJ�[�D�0Y�Ğ�� ��Xg.��{��!'`�w.;eB�WB]������T�зy�*�V�;so �%��p�@=I�dQɍi�Ϯ��;�t�]���|���dF�����a��Pu���Zs��y�����>��|��5�[WX��� �8��įbCEܚ�7�.jK#�w	��2�,ڎ}c�^glr�u����eʻ][ԫ��ٗ���[C����N\G�&]l
C]���T�^U��ʉ�4��T.A׽�k�-Q](LY-���E8�mD�%6��1�+�U Q�y㏟n��M]B9����Ʈ��{��+yY]�j�Iū!6��>�O����G�E��Lr�=�mQ��֚k��i�E��:N1�
���)\���w�kԇZ�
9���evi���jV�#ۼ��KV���ǯ]�t6��PS�)V`��n)1=4-�k�蔠�mw={.1[����uv��inW8���O彴8l��B�>9�S��`��&uD��1b{���)�5d��x�dc(�Wi�۰49(�U��������Ъȇ"KL�S����X͘��RB�oc�v;s�:��v��U=#sO%�Evp�����0��U������;`��Wvt�q��Z���z��r�*�wR�R句����ɼ͎6�eC���d��V��!�i,ju진@%`�Q�vn�_\�]uf��vy��BS�Ֆޭ2����.���<��Cˋ���,�R���l�2�N�����k��y���(���5$5Z��P���
W�2**�����3�!H����k�f�H�݁�9;Jun��X7V��I*G����(-,MԌ�E�o5�ǹ�J�:��:�jc�%�*��l���^ʸd`-�gd)	n�����f�ft��z�F
�:=�dW(����"o�!����GO����Rj��<�M��8;K�˫����|���M�,n�m^�.�<�B!F<�	$"�+H=�͒�,��-W<����Z��4�v����8�]]���o�"��vO��kX(�������[w�_5v��x$P啷�{q��,Tx�"�\�a�c��9�,I`si%�v��κ���Oh�r1ǁ�tx��2�.�؀9L��+����h�g=��$KY�R9��,�a�(���h��'���� ��9J���ƒ9/�ا�T��Vމ�Cz���;�g#��3�v��eҧ�\�Z`W�3/Z�[��k���j�$��H������|肺��̎��
j�b����u���9����Lvf�X5���n�l;�=�6�&$;�5WEg�P/@�$�i��%��d��-�R]�
V+�sm�q��[-�p�v_rr�rյ	��We��f�9�0[|��8%b�f�n]5���z�ɮ5���:�#��,�oe��N�0�rK\�z�A劻NJ�r�l�=�޳Y�*duc���	����Y��Du��E"�����N}׽�9�j.Y/lg<x���T;/&�D1�:�_;�L�5�����S!fӸ��j�M^���v�9����V�A�;z��i�V�T�;c��Hi9vlӣ���\�"���
�X0�{�ӣP�4�ӥt�E��p�"zZr��cN�[��-�.r�vŎ��U!��1�|d�P,��ЦbÜ�D���5؟L�^ǅ	��%,6��R��;�Xs.�wS8������;/s��b�sGZ|��8��Yڝ��V8Nn��3(1�y暊gJkq��&m���.�]�����0�jt�-AB�7 kO����� :��d�}i@�!�4��כ�9s�ћ��|n*�lg>��`��s��{�RU�(.�{%t�����D�7��l�L=×�`=-q.ޥD����5��8v>6�	�x��alq�xK��u�1������	���
zY/c����A����z����k�)*�\�b�ȡ[��.���9�X:e��Pv��]��1������C��g�H�1B�ͻ���u\��b|�C������QQ�"�lܧ9�WPc1�	 c[�՚O���T��n�Eӥ����BރM�i��_LNe���{� Y"�S<yýƭ>�՘�a�м�z�ل�y]�����&�����X�j鞳���׌���_=o P�0��L��H�v��ɑ��幔3V�.9ך���c�x�q8�kOm������Z�(��޵3 a�)X�|���Lu����e���ލ�&�����02�h�f���a�N`2�J8[��n���4��X=�@���&�X��8�n���f�Ϩ�8^�Z�Ea��]�A���������wGQզ��d��6��*3'vZg�d5)�nSoiN૛�xMh�`����7\��k�oy�Řk��ʮo�._�Ӡp|�2�f�Ժ���N�$_"f&��h��$!348B���k�+hXo6��g2�G�_Lf�9�Zި�T`XۺTb<j���)E(��+\ز �}� �[�D�
��<�dR+��3(�v���2=�S
݂d�z��&�#	�*C��2��.�CV�D����:��:��Wh*h�;�������̻6���p�{.:�|f�5sVm�"�K8w�c����[ŝ��[��nmj�����-��̣n��*dS^.c���*lo�
��8�*X2��#R��ej�ㆬ�u�/	���������d.GM�����/����{qP�zԆ��j=cLB%`@�+pU��,����N��NC�t��n�J�VrQ�#c.�^��1�_`�]�P�㜮����&�/r��3r�3�
g��X�2-|��ȝ����ƚB��٤�)����q1��X�B�rv������`�m��������n)�]]��o�j�ҋ�}%e��5�����4��ҘϺ�`$������7����]�Y����]�2$E��BR�z�JWi/��ʶ��Vq�MV�X(�U�Κ=9Ρk��18_b���OkeJ`�����Iw��`�莹F���ә�6����`�u�`�,��.�W;�\;����-�ވ)�vn�8r��_*�0��7v>T�-�|�`7�l�0	�����C��B;ӏqR}�W-���,�I�+.��D�L�y�Fr�eq��$���L�9��ӝox��Y�
RF;o���'�[�k#n��Q����E�[�HZ����[��;�P<Ӯ<t�Z���ժରܔv��$������cƻ����ھ��%�W}C˧�.�ݔÍ[���Y ! y��T����k#E�6v��L�Y���1�(�2�t���CLT��0� %�dRۇ���#Vkd���<j�rmL4�F��K�FV.��7JT���V��gc" ���Kz*F�{wr"�im.�RMmPᵝ��b���=ï���J�0c�y�) 8R����r���*����,�y�S0��[��h���T��U[�}|�9���R�{�q'��8)MUɤ��F�$��A���gl��ݥ�ymC�e1ԅ:���{B�C�M6E �f4 �%Ū籔i����+��e�=���[�8��4���e\}�;�.�MK�*P���6����R������	d�p���5պ]ɓ�T��T�Ĝ쩯m!vh��"�L��kLT���Ta���ֹ��j΢-�k+��R����&B,çe6r�e��V),0��9l�3]�e^*-S�S�g cj6�Y�2�'����s�i��E9]t��<�E3����U�dˢ(� z�
�.A/Ȼ�nuZ	��wsrj��n��`��լ=mdl�T)<G+B�����]]q���C��R>�N��x��G�o����H�|x����eI��ϙ����4��I_'Yu���l�&��x8S5��y�n�!�H��ږ0eo]ȇ�ؤA��Í��]Z�t���%c42Tǹ+�X|����r�Z����L�֙�Ib�;}s:����+� M�-�g%vV.tc�M���V�F���4(��ri6��D�kCIt�p�9��|򺬡g��u��W5���/;3�p�۝M]�cam�c[��ݏ��)
]n��Y�G-u��a��3�z�Q�Ee�'��K9%�f�a"]��>]�f�I�*��{C��֦@�4
n��r%��z[�c��s/mf��A`T�w�j�I��2�N�Ȗ75<�F�ƒdÏ��<7��.��UݽO�ݧ���]<�������ܣ-�ب,<�Ϲ�<k�:(�9Wo�8t�)!��
&:�VprW��⸕���8oOW9���*�5�̪�؋�b�s���0V��a/����4�J�a��g��hMN�n�gN�R�p/�*e�sQ�}n�kMŖ���\r�)GY
�1X_=`՘�nQ����9K�l,���"�R�,5�۵��$�/�7v�%�;FV@ӫ|v���N<M	7:X/���@[�^'��X }�P<F�� Uh�;���r�2���ą&�7�i�̬�
�s�����l���V�,���)!��U,I����Ncr�ڨ0ܑB��j���	B�Q㖻f�]����;"tTU�9��(<�����@MyBr��J�%t	�j����	˞��̦��G33��[���38j͏���푫;3(]*�N	bۜK}Պ�ь���<�N��6��(�i������𙨔�r�ۓޮ��j�|�r��]�����y��a���q*��naf���M@Eۆ�}Y]K/A<u�e�v��Tï��@�KË��� ҄3��cl��k껏+���\�.�"��Hc�
dh�t�OAB�%��\�]iD��;Ӄ�X�{W�@�����:ʕZ�Ȑw�B��1}����wy��ѹ���*��:�!�E�f�Q��v:`꬚l�������&�Wn�4�W���"j�]L�ۣ�c��ɔ>f��Ӽ��M�P��v�q��p���M��U�Y�[Z�Ű?�����A�b򰥨^f���\�m8N1��(��5�ep�P��ioz�@H]�*iN����޴�i���fK��t����x;� Lx�ZRP�Ae�)���9Q<v����i�d��cS֧p,�|F�{����3��;�����np��Y!�S����r��d�a��Ld@I�]'֎��g>�� ��Ϡ�pttR�O{oJ�e`��dP����s��޴̼�V��%)���ȵe#�R䈇�Lw�L�n;�u�[Y��f�J�+,��k�ڴ�e�{�oI�}N�]��®�h'�����f`i^��nR+jgT��4��+d�u�Ϭ�'�͍L�Ni�4�� �sea��m�)���iV���e�4��m��X?!v��r��ZR�\0<'���e���-�u�$��{b�í�Z��p�PȰ�@�$�p���N���7+��+�eN`�l�7��v��f*�K�8�E��Gfh:_VkU��zN;��Z�p���~_v�d^Q�f��[��pd����o����c�r�E-;{�h�s�P�E��#ozڛ
Ʊ^�жqZ�fs���Ȳ0Ec�߰��N�z/��*�hv�[��)��h��V�j��D��/\,�y��[2 �sm2�Y|L=��SIOD\���|�N����^X]�|\*��o�5���2:I#��
e4�>J,�I�HgwL=��k�Nat�!Ť����A=,к���#1��R�t�.��:���\��;�%������2�%����<�)�:�.dq㖗f�D���r��LKwj�[�f8��F-��lp���k�[����`*��)rQ�C�*v�,��]F���t���^H�˅�����a�7H����:������H�@�ۍv�W�W�2���E�/��u�k
�F�xXPJЫxJ�б�?�`�A�k���1����U����.B��h��e�Ŝ�3�gh1�:�FQ�`��uEigZR���e�B˶{&�4s�,W{\Ш6��k~n\��4G����Wgӯ"�����Ct�����c�Ɏ����Yűj;�Z@r]��K5
���Wt�}%�k�#�D��Y0D�-�(�z�$����Mm�b�]÷��C�=��"��!��CJ�j��[��`�s,a��Q�W�!k$ҷn�Z��9��k1�26�.(n��ƕg�",�9��*��^��6�+�-vf�
�i)��g-����L7N���-֒(ޞ��c����wz�+7��y�m�8e��"՝�Wsj�wP-j��;�[�h��HwS�nݨ�f�n�!�Hܥy%�y�s.e��W���[���w*b�-�wU�u��i�z�+���oF�7���J���^�lSG)�]&U��xgN��/�.��\���r<[L��e�jb�í��:ι��Ҷ�iW	�0R��-�&�L]k�-���$7�d�������C��de0K&����ܵ�7��s1e�&�:�߲�{2�Xz����B�4wdU�Aq�{��)��y���4Ȭ毕�1'�-,۴Ly��b�y&��:l���v�N�&鞷x���Bl�X����]�E[��բ+����=ƗC�
��6k-�׺�~�K�4'�Fj��[
��<�4*{9���� ��Qʾ�klb�'��������3��T�ʆ�/��v��{����R��肁�/�u�L\M�[�* ���*5n����*��-͑hv++P�6��kx���b�}4J싴�Y�Wo���<�������D�	�ʂu7؄�y��GB�T:�R��c�#�--V�a�������B�g}�8��U�Qf���+I�A.e��`�3/-�`�}-.{�ج@9��;�w%ѥ�����XA�)��lc�S�Ӄ)��D�����ub@.n���c�L�c;l�nc���馯������ih��&��tSU���l���t*Q�]֌�;"s)�zkK(G�F9'��A�հ�f��`��03f�xeX�(� j^�D�/��5="����!yõto6b/����2��Q�j��A��L�E�{����q�FQ{�B�KYF孆#Z��f�`���3�vp�5��ڸ�z��)��ۇ[ձ��|D[w��e�_���m��M)(���Q�y��\SF���]A%O���x�$+��z�N�F�ή�D��k��?u<6m�
�')�R�C �//`�U��{�uy4�Mh���h�~T�̢r�cz��j��[m|�*A˖� -��8�t�r��m�ɌF*������tV՚�'�<﹧t1�[��`)��#^ǘ&�lyF�sk�K���<�$�ܼ��7##:V^����]at��j��"��W)�E��C�7�,�72�,v/NO��٘�\�·1|�|�=@�:pIZ+w��f��F�:6
� �3�;��r��������'D�6!�#s���D�����
�,ۣn�[�54�7vM�Z�5ᖍ�,�o*��N�`�%X�����e�O`�p��6VLZ0뫪�cW�Xʼh�Dd �K�,�����<�]� a��K4y����p�S��-����K�31�UE�$Y<��J��#������?����W�ژ��"�n��Gndvŝ�m�"�:�90k�)[L殩|��ۊt�(�.���ԙ����~|���,�ı`�������e��l7yQStM굌f%���-=�I*s���Aõڮ����n����t�H	�R�.S�O�#�,"Cږ��ݷ��#V��]�At�9�xCY���o��:��A�b�V��f�]`�M�Y�-�]��fu%6��>�X�B1�%
��:�k%��雌.ϔ�}��ӔB�*�#{o��\��E��KU�4A��\��@1u1���j��x�<t��RY�V�p�� /Y�<t��y�#���m�9,1W���-�0��J�3[̩E�RX߆Aôm%ʵ��2�z��{����n��ө�K"�c�i\��XԠ�a��� J�(�Yؗ�ul���m�(`
��}]a%CJc]��\5�j�� e=X��Ytk:\��_\��;U�e�:����kb��d ��[��r]��C{7��G{��oT퇸m��6Gsǆ���)�W2C��TOѭ�����L�P�E����B���z4�2�������ZH�E�\��o0�s��O�0;)s���/r�.��d�Ht�H�N�Gy|c���o"x���T*F
"p���	C���-ќx�ڌV>л�S|J�]$�x�8����5!���T�[�d��řX�ű��%b�b�*[EU6()���D�]������L+[r(*�,K1rL�)qfaR� �u���'�+؜m���m1��QVM�)�+--s%�̙�����@Mj���H����m�QPH�EUY��\�3\�Af�6i+XT*T5�#��Q+PeJ+*e�delp�����4F+F0��沠�k+,Y���L�
�VХcK��EPQAr6�v��L�2ʈ�&U[d2XŖ��2�dK��nҪ)�ժ�[�0�)�n�X:�R�1Fֹ3�jV���QZ�X�lԮJɚ�������j�lK�Ԣ)+�j[��&���h�Uk]h(d*(-r\5hZV��[�乲1.��m*���k[l�c+Rڨ���C4{!��Mz뮾y|�����I6:�� Y�+J�1AƏ5���Qu�H�Y�Pj��\��*�'��2f�!Lt�q�L���l7�H�������1�D~�9n"6���=�V�c|G�n%GiH���t����ܤ� �.}�u��3Jgʆ�U�ƥtI�P�l�⮦H���=}4�p�%��y�-Y�Q9,$[V�j����b��{�׸����'�:I�!1�d�n�q��^��r���~�]3�WX�8����=�K�.8��G{ʂ]T�,�[M�N����b�H��5<�HGk�AT���������m[V̛�9G2�ƕ����yL��Զ�҄X��� �9��BB��o;�!�t"ӈ[0!�[g9����_ڧ��w���VT��D|I
��ɒ*Xkp�b�T�.�ً�.x���o0�r��3<~�u���@כ��!N1`>Hl����:p��t@���rzDSiJ}#�Jݺ�Ϻ���)���j(e�s	jl��!��L(��#�C���_sى��FB�c2FP�w�璧qE�yL'� ��\�jA=�.g빍RyagBAgOLk}���;�uԆ��wc�'%�
�t&fz�AT����ڈ�+M���j顯���iŝ"��A�3���IY[hm������{���m�����],��1c�>mX�M�:�"�ic�����ѥ�*�EW� �qb�d3���E\
����D����)��N�Ȋ�I.sr�%ڳ�,d�G�p7p2\�|�"�G8˩w韶N~+��Z#7>*.�[�t�l�>^��_�֭�j�c��傝+���8��z���*-Ki�y�c�V�Wo5QS�0�dI�19Kj�6����f.��.t�Ø� >���s��_Y�t��.��@�j�]\�LIPQ�_�w�%dNFq�@��tN��r�4�U�ҹ�s=��f? +�~믧`Ў)�2��	ӤE���t[rȂ��L�S��q�K�����պ���!����T2���"o��>�!8��T�ENTR%ӄ.n�bkk���C��ܲ! ����DD���dF�b�G�g��z�Y��K�9%&�^=H�i���XXn�H�f��Vd�%1#A= �.{��$�kӭر
����Z�-�K�ٝ���� ���H*�w��!�J���;I$"�J��o�
�k�t���t��
nn�ə����w�N�ɻ#��i�j֛�9f�Zٺ�b���`6�G+D�+6YE��+]gq���7��3M�ӕ�̒.˸�%up7e˰��ɶk�Y&�W�;yD������R�cp���WoLo�.�ܴ=��=�բ6�P�ܝԶ��+#���d9����E���r��
,�
(�FI�G=��ƧvaIO���jsdꇂ8Ϯ0����X\�!��6�Ӻ�M�ؑ)�);�ff�D�T�9<�vr
�Y�^#7&�@e���C�k�49*q<\�>k���nkH;��_T
Sj1Uc}��ɆD��p*^׫��؋!e�d#`$��-@j%9d�8����AH=Z	y�V1+/�|���6����^>e�Uп����~��?�������QM�o 6�w�����?j��p(0:6�5�~�{h]6���]!��ʴw��B_�����O�{q��c��C/fY�B͘*�6C�������-ƾKn�+z�0�s�����I;Y��v�>��
y�4Ȳ�Ψ�戠*��nǨ(���E]z�rd�=���#~�}�p�@�3��7���(�R8��z�%UMFx�0l���E��X�@E��+t��i����lp�!��uFg`)�0OI+�(9΢���#���iҾ)�%�z�M��eoS����A�����lT�����:�8�9;Q�j�Q=��^[����}���K+�(]j#D=�@;R�9�Ƨf�N��v���x�ם�pQoD���;-��m�;��R�F��W�|x<J��2���r<y��æ�,����$��}�wF��i��+�c;B�դ<��W��b���5ڮ�nf5ˎb�%ߘ�[sE��d���W�h�UC�k�:"+�t�(7��m:���kHf]�3|y�67`�-�*+��XL��;���R
��g��D�Ґ��c���Z��U��IYp�ua��p�r���!�I)�oj�7"lA)P�W��^�L��c��0Y�k��vo��)J(��p��t4չdD=�# 炥Gv�J<y�72*�1��	D1��6�X�e�@[S�IKP��<��S I���}�/{�7C^7)��
'�@��9��[�u��ـ�к��q���O۳�ft����� y�ׅJ<���P:Y���^�q�
^y�K�t#_7���&�EJ��gq�r�-(��4�A��y�Y�3�͚��9~����vr����YO*��抽���d���vl-�
��Y@��j�}�7�05��-�d}���.=>n%>S�s&�q�ᒹ!	�Nնc�|���Z%_mf
�������Y�aУ[���$�J��G�S�ċrt:y���s%+2�x9s�����l��wjn�J��h�n˷\�̎����c��(qԧl ��\;x�q�;Q����7a�ۗxE��!�Z�2�%Et>�d7B�(�l8�h� ��1Xda$/&�G鞽g2��t��/=P�s�Ť;��~}4]�����62R�Ï--ouu���$�Hf�G�MUdFwćVtS_�ԭ^}�u���� �_�^+�_�nA?��伂��-	�!P4�4"4��fL�a�$p;�8�[ �����>�r�O�{��^�������[�[1� �lt���"��}@�Ц�p��Ƭ�T�{���ꇘ:���2݄�7cώMdsR�$�B0`t�犪����7c�2`�?0t�"_:F�j���͟#!4�<Q#ZB�i�HG"le��;Ef��ݹոIf7 P�+��S>�b�� ��n��k��8��E��lk7j�{bc-]�'��fAb��ʢF�f��tȸV�=�d=���i�K
���Jw�Ӎ��2\è�a��8�� �9�A�`2�!!mgX���u��Txe��ڀ�9�jt^AsK��rcf�I�#,[F��N˛�KF��,`�=*��p�"ku]:(rt��a�{�w��uwG1�Uo�NDw5�$��8��2�o<Ü����7�J�*i�@z��KGG�q���ة�q���Q����2(t�f0���n���r"�!P
|R��'C�3u=��l��M�J.�"��c��/�E��h3I�臅��]@�M�c��8\Ř>J���S�)tvV[��N/���=���hS��H=��$�r���P�������,tjb��8���&����A����>�
�@̑����J��g�b��x4��]s�0��cʇPqE����Q����f��g��L:-ڧ;�zh�����y^S)Q��Q��;7g7����Ǘ%M\O0lVл5.U��W2c�����:������1��&N7��ٝ���C,�^�v1�}{�����7z����<pQf�i�|�OXf+{0���w>��R�=���qC�8�yV����س����ͪ��=~�u��4��]�}�;X�nƃ'���pU4B(����S�VU��l�th����=�`]��3݇j.�8f�t�:�|���r8��r�9S�5s��dA��λ��j��^������xFYs�d	�.wP��tT�ꎶ �f�4��WK_N�竗*�2ٷ��֙�-r�I���"i�:d�����#*
T]FR�j���q��C ��nem]��*]9Y�6�Ξma�sT2���eВL�3&�d�J�舆
��ǌ�jf_E�"��]�����2F|��]3=��\F��wK��ƞ�˔t�6�(Q>00��:�Q#�zfY瞺�^�e�佐w��=1�:�*�0���{��I���O���bv!\x%"$h3 �s�D��N�~�#�OuQ�]�^+{�u�=��3���h��Q`7;�H[ l�1�6�M�R'n��`�=	�bގ�2d�ػ��7IFz�ߓ��;�Ҕ��T� �� w0����W\�3.)����:��#��e�������+ .G�qN5;���ہ�Dχ�����ʹ��v��r��!S��2h��8B/Fw\��k�<����r��B����X�Yod)��[��-�D˥1���p+Ҷ�Q	�؋!e�d#i*��P�0���;<�{����#՗�Ƭ����.��ܟ�`����V��c\U�h�#JO��'Hk�;��˻������D����Ā��i􈹑Ca��t���|�/�*�x�D��`�s�0l�i���%��@�ҟ�>r���w{��+�S�fm�bb:�
�m��#/z��{3_0�eȸ) ��N��}�N�(i��y��f?H��m��n���r��ۮ����vQ㚫�5���;{x�#�;3�#����ؾR��ڦi��nl�W�dע/�Λ�y�^S���^�.G�h�﫵ײ�m�SH�*\�Nh�X�g���yE�\��|.r!ڽ��C'B�e�gbJq����1P�+�_9����Z�=~M�"�t4�r���9J֮[���dY
L��:T�=$����'�p�E�f4R˾��+^o;���"�Y��}r{=r	��.�2zb^Ŋ�ud�f���ة��v��:3{�U��=��U�x)�!��_r�J��U*��5ΙZ+�t�ӟN��n�-������ݛ����8�R\
� �O��Ni�N�T
�^��g���;Ʊ[_���b�����*�:�])��~���s��wc��"�۵�Ȃ9�%#WtVf���k���0a�<�(#����	R(�N�:k�����UGS+��S<�-�<Գ�`�P�#��;&�Q�^Bڞ��5�9�.J��sea���f9=:��N`�5ˆgp�Uc�e�v�	e����̜t��p%kT�T�S&�|�fK�ͪ�GU���y�Ė��+.[���Xp��Ry��S�c,�諠��ƶj(>�� �����z,�]�F^-U.;{B�WB;N�K��Y�q�i3vj|z'�Ho�}�C�t��҉ݟ@`��g��uf��^#\;�l���>T���e�M���K����T�0l��Es7�1ŜL5������\u���[9z���W�i�2���`v���}S��&�QA�1ps�W�P��=@�5;8p6۶�R������vP��]?>wf��`��,�BjI��S�~>g���[�8s���J�Jk��|x�8��r��6�x�ܻ�/zC��L�{4��C��aEՊ�D�[WX��T@���-��R�(ʷ^Us�G���c���sϦ��}z)ͅ�]U���ob(�̙6�A9'$#@�B�5U�'�AG��}�)�{�ʺ������i@�?3�l|�(;���e��ә:��$�Y���8]�up'�B�v���Vj�$�w��1T�k�z����Xz�f6��Ҋ��"��1N���S���g-�,P8d����T{'�S��7�|�j���&O06��6�m������%�S�a�&|�]#�;�^�m�]��2�k����5.Ɨ����&gM^~�^�=��i���k~X��)]�ɡ�CA�So��4��y���h��>�W9���i���n���Ճ��7lv�	Z�8�-×�g)$vnu�v�ׯ,jS�A������gpl�Ҡсc���'�=�r���!�oc���q$�L��s�Bvy���}��W�Q���֍�!��P��Mt����ȭ'���������2��A��F��$�)�*5�Y!Z�\<�SR7�mlJ
*RyϞ(�CX�V�����#iϡ�9�x�e�BB����aA��Y��e.��NOfd8���,��A;v,}��z"�!PS�ע	��Lة�Pڋ��5��b]��V4�w�Co�S��9���۪�E�1���>HT�W�u�����T�6Xr�_��I��I�r����A�2�`a-M�0����E\�[��m���(�"̗1�'���72FVk�+ J��{>S��ZRN�\wV�F�
�o-�ط*T�A; ��|���T,�llq́55�җ:$M:�/��E<���o_[���K�<�ԙޗ����@�*C4B�����7*G���3�������O��ܡ����ʣo�Y��ì��{u�����F�`�p��rK�F�y4�:��%t��p�o��B�f�{P��z%l�m�7W�������f�����썏���n�S����L�P�1;3z������ˮ�dsQ,3o{.� �]�!�5sWC:@x.�L��̲U+�,:���ܱ���ώj�HʠU��sd]iN�]�yb�,���	�8��:��M�7۔T��|�sW5��D���k=��$j)>�e�z[e[r�H���MZ.���&����z6V�uш�E���5�L1k�g�L���Xd^P@�ӊ��WdqNY�ط�ݯ��_$T�B�l�Ñ�Y�)g��A�N��1�cm������o%!����MG��2�So��R�L� +w\�����WH�vJL����5���2�sm�4���K@��^_$��z5����(��&T�M�C�18Dj2f�қ��q�ʇS4��+x����%j��O�x��r9���ZJ�j�Yw���#��!��Ni�K�-���o)M7^�rnJf!���v$���xC3��Ws�aP|�Ӽ��U���h��q�v��%�.�/@�v�<��*}x��4��n�W���'kw|�c	<*��Ԃ�^���\2�f�.Bv���e<#�eE%-ǈ�|-�,Lʒ�xӬ�N���{s@瀾�D�=/�z�,oPPr��Z�7������-��v�4�Q:�(�1���@��3-���V+c��v��`���3����[�O�n�c��!�|+0�WMӣW�׹wF���wV��I���+L��w%#1k�>�/Z��\���7�r7�d����t�X���hK\�|0��⣸��;�+�^bpkc,m8ŝ�!�����L��s���y,%Sovm|����6 ,�����v�����'��ie��^;��q�Ě���^�̈́��$`�p�G-D���'���+0���f����Zr�굮��@��rU��)ޘ�(8����.�mm��`�E|Mf
WzW-HVi������{�hV<�)^�U�������y�t�Mv�FE8�׌�_u�\V=aiB=�Gi�Ma�'k+�;��(��\�#��q9�UdO�B�wE�g!7nU��n����Ea�vv�=`��p�z�T��C���'���H݊	��ʾ�P�X��eq����S�P9-�m���zWq���S���RE�N��µE�c���K?��k�Nݠ%�-��&���I��̛���US#%@s���@%)�kU)����TjrN��P��[�"U#�5�mEƺ�Ê�!����e�QV��^	H���oJ)�}KK��Z�Q�'K���I�.�140M��F��(�K2>�u%�WU�o6���d>;D�G�N�;�(c2��ze��7��
��_����>�s3�P�icۜ��[nJ���ivع66��̪9���Fks�����ܔr�j���J�Z��l��n�kn���Ѭ�`⩶՚�[�Q��m��cl��Du�m\�Z[m�\����3PiM��P֨�Vڪ�]K��L�2ۭ`�!���(담Q�h֢�����[e6D���9(*�
ƛ3mk[L�f�Z�AJ�Mem��G&s����5��q��iV�*kR"�#R۵-6m��DK���mUֱX���ڢkB�-E���U*�M���(�E*Q��%�����\�1�J��)Z9���sm3Z&�V(j�X���uًm���i��֮kQYQ����Z�kJ�]����[�W5SP�cG1�[�#�%�mTE-������X���[iu�lLҥR�fhً�V(fA�n��[u���ArT3���2�l+���i��v�DP�lr�*���iR���F3b�iv]X�-5�15J۬m��*�Q��X�2��V��+���5D*R��m��F���[X*�-�����Q�?��O��Ǡ��
l+Y�^���ܜ�T�J.�Vc{n�Q��J
�YY*F���e�!���]���۔��[W�w�?n�e}�}�G�����ފ#٨F�i8*�U��:�:��xjS�X�� fk�gLHE��K:���Ֆl=�ّ`w�靋��t��:�b�FG��K�m�gw;���P<�����_F��!�p���O�x��:�a=(؞�,�������bTA{˂F�O��`�)�3�:n�DpQ�:&2 ^��[ع�\�ֻy
#��%U�B�?�]��PG�.=|#�2�1
���:�N��3՛��í(�GP�"A����:L:&e�x.�z��YX�`=<zݷ{�o.�d���%P���7�L��'I�G��TUeuPC�tʦP����ާ�R^�^�bs�a}&a.��Z�jD�R�nv!ߜ�HR ��f��<�\{[�29�3�����ī��N���8B7��2�Ba�Qh�(%#���M��8���:-��7`�w;e`.G�qN7�����`{�v�|��Q���x{��s���Z�r�nӇ���vw�t�[0�
u4L[�DuL�^�'���7=��>��=d}����<��[�8�Cuo"�>��2�v1��f�ﾁ�+o�nS�3�̋T���g��Q)��m�0(˛�7bQ�P�v�X��"6fMx��5�y�Rx�q%J�C `z滳E�WZ�-�3�9�5���|��"���uGm���!���^N:�օ>(����ʓ�N�s}��Y�$K2�4��5����4=����]�L�:�]��|��0����ot��ڢ;����1)�&��p+a��t�9pO:gr�������T��67��ŋ�QC2�;��{���X隷<){�:}��m?�����q�wL�3SՋ�F�#�'�TF߶@���uM",.uBq$r�X�<�nǢ�Z7;^��t���V�J�5'��4�xeT'`l�gبq:e�e�E���o`�U�0�ȍ���=�H���1��#�t���)�BzI}yA�΢��ͧ��,&��zG�����3~+���=����] (0�7���,�;:;".��Í�or�TV��%NCh9W�mvW(�GR�b&���{Mu�+B9�z�'�#��_��ĸ�	un*|��3�W�f�hF��p�@m�n��.���:�֪���'�@����SV�Һ������ew���eθ�L�����<�	{���,�D{�ms?�LmFj��,��}�[u.��c=�K`���b
4�r�"�(��R���.�F��ac�ZhV��6�du[���mv�@qvz�R����CH������u�XlDWC9��3�5�"}O�Ey��Q��;E6;�#�&��j��b؉>1�>� #s��B�Q&�#���i�nY�GE3B�N����imj!��=B����B,�B��U䩨G!�8qx0�j���D�U��o)�u��0}����L���(* �"�E��*x>[�%e��¨V���=3��.ԣ��L,7T
m��r�&-���5^���dn�-�A�o1��C�p��A���8�A9d��J(Pq�2y���W��;6S�u�z�K{�[���Y��~�8��0�Μ#��wf��TP#STM>꜋��[ӝf�Y��Δɘ�k��*�U�0#��aʋq������czC��S-f��yV�{�	6��/�Q�\c�C+���^{PR���TZ�7>�^W<�3��Xsk��b��yy�xN��|�ա� ;P��������{v�(�RH��[zd5o��݆�����ωi&��ok;M�n�% �hX��J�I]g\��Xyȝ�o��9���f<���P*gvS�eޖ��2go�J�a�Vd�uv���>`D���{)$�]ڱ��-�։�l]2wl~��vh�A(W�rM�3�g|HvtS_��w_���.�vv��<���'��p�޿}��FJ�d�@��Zς
���|L��������kSǮ+H@�T$�.�p�<������g��]l��Ѣ:QV�Z�cR��XK���=ъP��,z�B�*�O�nӰ�_�O����5+�8X�/V�y��{n��~��K�ՏX��8�)�=������gsg�ϓ]+��U�nD�z���*zo�ֻ�q7z"	8K���(��sU@j�p�����^��_[5�2����
}�aY�6�i��$�f�!��z�VA���=��,���s(�.E�1���6Ҧd�ڄm9�8� "c����������O��{U؀Lfm��s���8S�Ca�[$�$,���L�1,���/��-z�^�{6����O$��E��
�Pe8}�t1E���f��V8�B�.b���6��X]�k"�d�8��s3�<�NWuhǣpZ���FepKF>t0"-��W�I���S�7���-W	w�+8�"a�W�܋����1*(t��7�ԮQ�bS����Ť����.�[ڛ��*����T�1��u�E�(�*�78jMMޱ���ߵj�p�vo��{~�"��'�'x7,�j(aq�/����-�9�]�J���&,�Y�Ff��;��35��]E��1I�{/�I��w�-ŀ��q�
�O��@S���P���9�&�f�ZI�\���ù}��]mݒ%�2���X	��q>��y�@ح�vj�*�b��u������`ߵ6T������o19����>�:�@7��:I��a]!ΑSr4��.::���\���前=�G����Ω�̀�K:�9��&Ǉ��,Īq�l�<&�-�\�Ci�刮����~�=�v�7���WN9���8��h�mG8i�l��'`>�npB��鞺[��̈�`3tOB�R�8ʂG\y�
�<W9f��Sy��ˡ�Ö�ʷ�=��",��<����)�$�������:��>ƅM!ǫ�s�B�n�81��=�.��Y����1���S/�ZQ́�q�
"$�4T}��S*�:Ixw\hW�;��mgN���e4����HN���qB-�Sj���t���r�w�z��F�3���״8��u�<o#�݁�O.='���E���~�<aa�'�Y\2��QLr��՛ؗv�Hm��\�y�e�+ʜ���9bΐ���,;{ׇ~�fw	Q�r+:�����bR]�Pڿ���Z/���C�⍹�sX��W�	LH�uQ�.���+^�nu+"�s��.�pr�q�΁�^��A��J,6'b�$�� ��:��6DtdݪƔtĂ�-s�.I]��p�%p���9݋�;v&ľ�"�Qd�P���=1�T�t�)����hp�T�$���H�g WE�0RI�+��3bۄ�����j�����;�i�-�Y���fB	���2k�-��w�RR��$�n�!�$�ě����k��v�^ �Z��'�J�s�Lm���$�N/��YC6��:�йWc1Ǻ���Q*r��=/�:d�"�kӖ��䶃���H�2��^���(�iQz�7W0��
P�VHv;�-k�[��\ *�� ~�F��w��aŃ��Ĭ��m9�N�r�QTm��da�d7����C�����f��x�-͘*��q���A��U{6��W{o�kA`�鎌���g"6��t���uM.���s�0>�!b�q�J(TB1)x�,px�vL _'�(�� �t]�����hsT����
��{5���#9�r�SK��D���H��[f�G��[��ѣʞK�Oo��-�G�-����̔�fK	����·�%�ewP
��V��]]
)%����H1H�t&T��p��2Y�!T͚غR�:��D��g�e󑊪�)�z���{����ow����<���]:cb�"�����:�*T���R&s��%���޼{X骼������.a®�{5Q�=}r{.h
44Wiu�����P�R#��ӎQ��zz��Ofw���xv���Ieߓ�݇*�ʎ��FLr(���Q�e>{����<p�	��=���0p_K)Ƹ.�1�*J�^p�H�u��͗���U�uR�@;s0x�ٔ���dH!�ȡS+��ZlDR�s=΃=њ�>��bm��p�%59 ��0��v*y��#�P$�1��5�{�W����k�n�E�N�t4��QW0��J�����ol�bm���L�d��vA���Qg B���ǒR�ᮑ�v�Ag�I�ny�z��Ш'�zO�)�S�ҙ�8�{��PO���E�Ʋ��TO�N��nzqr#�lܨ�f�!7<a�X]���7T!M��i@�)GT�x=���ǖ$F߶
f�X��!��5��4���Jz� &�@�滱�8=*�f,�(���H�GW[��e��ڳGM�߯x�����8o{�z��y2�J��xqQ��Im��s9)���#�-�֔�YݮU�(T��y�n�N�*5"�d�rs�s��uz���םF��QN �nY&�iEa�8���y�uy���[@ӓ{�tË���5ڂ3��wi��J0��$a΋!h�wu�TX#CJ���S�es�8#��#{�z�!ھާ�`�!�9^;�g)��(�n]�7�>�kX�Qof�T�Vu�N�y�\��ᷦ��:���<M!vѻ7H��
��@nU�u�&��6��}[v�ط���Kku���C;e���ެ�<^��΀M���!�^��ؿV?f_Q�v:e�j#pz���!~��*Taə]Ϊ���q��-����ا`�pT�pV�����l9���^8}�w��P��w��9do:���#aOS#�&�=~z�f6��th��r8jX[<�y���wܶ4͐�0�h=ѣ"�VpT�2���7O�GVt7bI�A�V�z�K��R ��zY�ʘ�8��IO���;G0j���͟# &��'E��9��{32���I�Ŷ�d�QǢ ��$Ўz�R�3�s>�Q��a��fwk���y%�QN���ސuN�_oW5�w4K/�c3�yC�J�`��K��5�i��f��J�.ܛ�b䭼�c(Hf���CI>.���lbg&Bɝ��&:ҙ;�j�����R�l���X	ǐ�u��M��d����/�bYϟteA��\qdW���b�:;�),�D��(ʙƹdt`����vb=d�Ғ�r�����j{��jٓsP�����R�D��>�����j�R�l�Ԣ�[��)�J;T7X�8���(P�:�p᠝�����d��O�SB �sd��`����xq>���Wێd�-��zΨ��X�/��b��4��(�1�ƺu�M�����\)f}�����iۄ�ԪH]�$��)�8�X4QC6*�;7�z+u�jkin@D��X\�:lȘ[����^d����n]Eϔ���l]��˞v���v���P�u��6�zA�lȲ$�2�|3�I���;rqr�^OE��W+yޒD�򼦓X	�Ҍ�5cW��@ح`ݚ<k�خ�ܽ�Mdтhv�����q� �4J�e��i��9?���{�>�y��o+&t�����W�e]bB���h�zqoE<d�/h^_L�b}���[ag��4�Y��P�[XY{�#Ta��Ś���U��7�$���{L�X��17�ãF+3��q��/Y8�u�o�qʰV����%$Wu�5��'S�o��(j/5�eA2�X���v>��F;��V+�x���%�Y�)
�mC-g�
5!�7invKZ��֤�Xn>����7m���N#Cc��S�~ >�! ]":]s�1$q^Q�ZnƜ�ü�VOxmM넏(�Q���:�d��;y;
�]G��:�O��`�+��N�(���l����ҧ��S��u�">q~�/
8P�M�U�($+�I{L���#��{�����[��b��ʺ�	�4�T��(U�"���B��=#A�}AX���D2�o���I�\�'���/�Hb�+�9�K�1�*��qF���85�؅b<04�����QK�N�ue��j��ȓibRv
�B�����tE>����Qa�;��I$*!X�q�LNjo���x�/��:�,Ct�d9���v/�b_]��yĬ�Q��<|��a&1b	ޠd�%DB8�ЅчL��<�r8���`Kt
�W��~{�|m���ʙ��B)�)_��ad�rhd^wT��k�.s	Κg3��{L�w�j���Ȍ`�>��B�75�d��0��ہ^��$ИN2�Y=�MV)a��a9��C���s9����]����,�7Y�=�+�p��i���U5K/J�����4kb��x.O��S�u�[-RU�;!��=[�lʼ��F�Awc0�vxLojU�J� �Z��S]���q�u�Q�7�-���$g![�t�j��;i�)h�Y������;����%W�uiP�n��Fۧu��P�Гo3Ptrh�ˊ�mMs��QX���3p�ځª
����ǻUp��>W�K	���͈R1�`e*)w�WU�N���A.�4���4�
u_�i7|w^���� �raK�I6�M��z5�^�r��Y�\X���������d8N>��=V�2����k���:~/�/F��Qd[t@��]�W��+.�Wan;�[��	�{��X��NQ�s
s��sݶgw]���"K:Fhћ�dH�ϐ]�w���g,ef��>�Ѻ���@3��e����[�`[ǌtr8��_F;B�o+�������q���ïRj�h�Ĉ�����[�^L�q�ٴbwe�b%۝H��9i�؄��P�{��J\4s{%�1��m��!�zj�E5+���[�樳X�*�Mn.
�m���As>L
X��݅ga�4���JS�A��tA�r�O�e�ͱ�8h�Y2�f����am�kit��TQ�Ҏ˜�V��y��Cw{#6t��id9���Y��r.˗{t#K"��3�4�.mQ�!���l�hZ��:+�/X0�0$��l����滙Y/�
���g�Y�ה|�G(�;Zpօ�L[��cd�dk�;X���5�)�,��J���2K��"XÂqk�ڙS��$�q��-Vt�M��/M��W����"ו&����o����:�vk�3�Sh��g`�����P8��@u��E<���t��.��w���9х�Xu���0RN��7���ō41ɟv�a�˝��L�X_R�E�Of����#�� ��~����Y ��� �������k����f&�=���4�T#7t��{��!p�W���8Ku������K��X_�(a+4��2�=5h�JL��sk7��.���r�>�lv�=�Z3@ܾ�6�Ǹ󢞈�+�xY�D���[�{f�^�1�̹
�8���|N�����3�GL�բ����&�R��u�-��Ki���$�"��KS"����۫�v�*�z�e�j�
����cEM[�7ܰn^˦�L��� +#z��v��a�z��+��.n��"��An���V���s؋�2��h�D;poj"���'q��t[�����h�>^�C<8��zK�K�.��X$u
z>R�qӚ�^q�+3�&rF���]�(le��<aA���;��܆��}(���rv�O;w�}`sM�E,Ζd� ���W�eӜ�Vfj�6`���[��+*խ9��8(��+>����l���T�\���Ց�r݊�U,��FԶ�т ��%ڣ��(�Wl�5Z�Jݖ╕kb�52�Զ���R#mnVa6��ʬF�nؚ�R���:ĨҷR�]nb6�YS2�JV��T�(���6���Kc1LW:%(S6�%�C%5��M�mb&�f֖�ѻj�j�mJ��+R�h�Z��]f�ֵ
�n�sv�2�%U�i�+V��DE��f�\�Z�(�6��6K�m)eV��v�[�Q�沱m�D�ծ��bW]����\�2�ڶ��(�K��K����!��
���Q�S9M��m�[��b�V������b"�dɮ�Kr
�X�5�[���1͋�(��,���;S-m]����GYqT-��#hЬEED)maQc�7a�)h[u�Gm����)�2�3�w�?�����]YM ".�X�7+��r(��L/���.��θ�eA���;�@�h�#���|�ƺLj��������uã�u'�}��㙳U�8���'L��A�{^��{�8�R1e�0x��[���[r>ӕ��U�s;�GUHˇ�$+�wdXZ�VI�	�%��6��t��P�3��FVUgwrGM����gfg=��3*�-����X!��ڦj��3���靽�G!�<Q�o��\R�5c��a�W�ׅ��T~�]�kO�����7�LQ���	oh֥Ln[��{���涶L�L����xs����B��5�*Gw�Q3��������g��Yx�k���ޮ���O��h��6�j��	a�^HU�D��D�HBBڳS�,�_>��F���^d��,*�R��w�5Q���=P	�(D�b�_B�Q����f�r�s'vD׳��ZrNU��
z���W�h�ܤUz3��ƳS�0��	C����ę��S���AQ�&���i1����3��Nu�i���H-�D�D�7�����4��&T3o�{�5�"{͊�~���!yx`��8=ٲ�\>�Ë���t��o㛫k8�/X�*�����,)��?/z��dr&�兼혷Ō��X*�02G ���fƪD���.�����	+�=���m��\P���۬M;�IT
=*�[��&�^b�t�9mrq�G�_}@d��w|��[V�}�'b���D�2a(4c�⏑��L�+V�;�4�]���������TmhӗD1/n�OEK�pAA�vA����E�[������v�$[���K5"c3�0�F�'|`a�N�X�6�\+
/�ED%fA1O=os��"ʻPl.�K}y
eF���c5��ف���A7\a�u��sF��n�2.ۙ��:l��RЩIF�T$�V�ySƘ!���C����뺋(�k��$��l�1�i��h7=�[6��D�~�?m�����Ѯ��M�H�Yӄ+����`���5�LD�0�vP��̶�bܙP\{��M
��o�7�����S�k��y^YP��vk>μ����~����</��h-�P3��B
��
캤z�bTٌ�E���Su-��S;��_jJ��hE��!s������g8^bB��U������xe3�$<�S�{[{��|�#ŗ�%߾��f�U'�ڱ;�Z�����'�;�� �[���#n�[���{P�!�K�50�X����q����z���4�ϏoO7�K�4=���:G@�V�q���p�x��;�.�����ã�����09�)���x�f�o��J�K��SU�Z�;L��v��mµoE]E�ͮ��;4@KR~�����8�~e)��y���8�h d�I���\`��S��m������ѽ��ҞPg�2OQZt릻{X�ZhD"��@�tP�8)}��S�����O�GVtP��d���Z�d).��ź� ��b��J���`h�n�(�O+���4�G��L�7z�����g/f��-y:��
��*����B��U�<%4���i{��z<uG8d\T��O���������n�ݓ���"�}A�cʎ��
U8I��2=R�����WE�H��65�U]�l�|��VC��N��j���cjN=9�# �\%@��k'�i�s{����g��ՊƐ�:J����YÆ��rlK�EBQ�En�U{и��U�����a���]Ot;��#��lPVT���0�[���3)��h>�z�aұ�'�P����*�F��u+�M�JqcR�"��&�)N!�r�u��Q�ݚvKsj�w]8�Qa�K�
����6fae����7ϳ}4{�^e�y~$�I/���f]>��AY���@U����� ���6*�/v�jU�=YR��N#���֫WC�+7�Y�Ñ�%z?{ҥ���rN��mq#����/c9�z)��o�+&>��}��%'@����ڣ�7;A,�_N����Q�ߪ��滋ؾ�m�q;���fJ%#y���6���ߌ�"@)�dIW��G3��q*j�?rwZ��jy�j��~I���~�D��)�X	�Ҍ�5}.!�p7p2exb���DxCy�zw<})SY��]QCr�3}��}щ�D��}�G��}���0�Fp1��jv��u�.�R��M<�����]���.��Y��|3��y����xOb�J��5v6���;~��7{z�@Q`��z��vUH��Br���\ �h�Q�I\��:���8'4eK�5�f�40�p!�6�T��6)I#�'�o��j8����B�����x�M$�	zs�iW~Q�:/��"6$�D`=!u�̐�$��>@wb"���x,{=�b��;7y5�G���e���R-8QC`ak�DI�C�
LL�}����m�vj�B�٬b�H�mS,��E�'���qF���:�dB^��$h3�(���U�W����ú!�)ŁQ$q�=�ňV�a��u�v�v-�t��Qcޥ���m�~^L��jju9+Nu���>�e �]+#�Cx�xV� �̱n�V�� �W�T�砛�\�g)Բ�u��e��l��bl���^��ri絋ळ�R�U�����#��E���9u[YV^�N#J��O��t���_�xx��Z��aI���T;�{��+����p�%r�,��p{�յ�徺����7-�DY�Ldh$�$29���qŀ�.�`�I�+<\�!��wy�n��.H���Y�Rɚ=��ƺ����\� J���+�Պ����3b��}E�ܡ�t'U����bK�c���|�E��ָ���Ũ�p*VГS	�Dv���nm�`�u����Z#y����ҫ������N�4���9`���3��b��ٻ��p��C����=o��?˦X���t|GW��h}����%���D�MQ8�D\
��'p8�^�ƥ�}���{������xw=R,�4G8�3/,,��}a�y2�?9�I�c\wvY/�Y��<�o�j�^H��$3�N�v
�r#od���M.��S�q[z4�ꗫ��@��p�D��^��q�.�����Y^,�Bf�l])q��ъ���|�Dc�}'>��2��j�U���X=�e[�|x���E��rB��;i���M��J�I��~�f����񃓷b�]��]r�R�:�����L��)!oC�yS���M�ӣ���dʃ�i�q;��Ǧrv�s�9���L�>�Y���k��e�u)K�T�6+�뒳�L�٘Րl2ub}���ٷK�������5}M�-q;(��wG ��R9��R������j4�o_\�ːH�+����ai�� ���ܙ��P���vD�A,�	�nÕ~f��C���&-����A[^xm�|}��Mv1ǈ�LoFTS��.$�C)�xk��e�t
�M+ p�H��{�r��#�X�^$'�]Θ��%���iH�T�s���M�"�3�9�g�3\�*���my� };��*��׀���s.��%*��d�PA�8��r��;�V�j \FX�.�V5�k3�0��u5�RȈ{T�hOEK�H!�Nh�IE����dm`��� �ϧ���k<��0E�Н�>.)��
�B�ED%`��g���ܶ%ma����iƩ�[���t2)7\a��~s@�=��J�E�/ݚF+�]��;���j�B9�!��5����8S�5��ZQ6w�$�Ar��P����Vn�t�=p�˯�f�/�N�Kq�n�:p�}���[,Q`��%t��\)T��tu��̎U��m�����[�x�+`���h���c�T����a��vܬ ,M��3&�-drCQgR��:v�^�!#�12���|��ف�ثxD�=J	g�����E�e��%`{3L�fv]��̾D���:Er=�ػ��{�
ʎ��n[;	�n:��b<����d�!K�Â���t���VF��67��,ݚ����j�뱘��z_��
�Π<ea�?A^۠��P�*l�^R.,��2��Bv�N,Zڹ�YG��P���(>�.�=Y�N�2r��䜐����ءM��,�����6{"��dZ��ʙ��U^ԝ{O-Yl�}�r{���4�<K���U�Bwo9��6Bb0ʊ��{�Br$��q���7�=L�M��✘ȋ�4����&��r����c�Y��`.�!��N3��w�>e4�7Rn�˔��C=����<��7�������g��~��8И)�=��1,�:�z� LW��&��fߢ19��UI���SN��N�ǉ!�/���6*e(�S>�2�:��:፶�Z��M�B�Ӻ:t�踡qǈ���"�gL�"�s*��\ g˸�faͼ�1{�]}�A��7'Hp��{
�{�:'m�fL�E��P�R0�[��"tD�.�o�;�����⼜�
����k¤�Wt-��˭*y2���fP�ӨT��˕���[�e-/6�}N��˅u��1��t��Z�f}�Z�r.K���YO(���8�,G����,�8aAN�Ă����UUKN	]՜�lƂG>H{@gX��S��9΄C6l�	۹7/��&�!`�hd��9V^)������S,D�q��}��/�Qg���ט��NR=z����|��̝M��?0��ϐ�_������2t_����������m	#>y���]�em?!�>����G(T���tF�!PR/�ӛd�"��z����fró�p��y���^���$��9����^9��<y`���=����3ϓ'�o5�&U���y�gj��n�[���t��*��C�������=RT
���<I�+>�ɓę2A~J��'(T�S>��;xAH�N0�	�'ng]���ԯ�O�c���R|�����M_�?A�o0ָ�\����Y���6�����p�>xL�'�bpϙd���x��Ar'�y�I7� �����
T*x�-�����S�,Ȥ�*AY�L�ä3?Nl�����̂������ͬ"2�~��%o�IY����͝2d��y�>d����|��9J�U�3��r��ORp�{��v�YY+���7T�,+�?yI�O�&C�,�l
���r��b<	�蓢�:'�S��vr]-�$����0X/L9C33���� �0����:NR(�gG�юXr���Lÿ~����RW�哰�y��r�AH�s>���Y��ht��dᙞ��2�Lǽ�s�ٌ����S�.��oj���T���5��3���q������rY��S0���qT��ȥM�8�?!�A}C�9���J�׻�
��+?{d����8H/�����'v�������?Hu����纻�0�l�< ���2iS2v�S�N=J�έ��I�S�=�r���o)�����t�YC������ArN|�=$��!���8�P̘1��kG��u]���-Ԭ����2Ag����q�I�*���Y�L�ô7�X�{fI�jEԬ�Y�� {��3�Nu�^����U|gi2
E>C������'�G���.�5Ѷ�¬��r���癤����e���{:�)R�L�ÙȽ�Z����jΧ��.z;[a���vL��kI���d�;ަ�z�"��͢c�>/5l�h|��X�w�TLD��7��EM��V�=�c���w��k)�٩��MwܝL�Ɩjލ^F�JZuob�{��۴�m-Md��AGޮ���W���$�=L���~����*:=�q*��d��m>B�fa�d�恟d32/�d�����Zp�%H�z��48a�|�ə�S �=��v�u���vӝ�=�߀d�!PP��p����y��)��O���پĨ'����>�9}`T�3���'hW�Ol,;k�%a���3�3��d��dR�" Q�*��͙��eS�Գ|�z��32fOY����(%H/_����I����I�_�?< �]���
�=d��y�g��ԯG�yğ���C���(p�dɟRt��}�Yq����q�D�E��ݟ���26�÷�� �e���O<��8es���]�<I�r�Y�7�pzäRv����g�|�?�~O|�$��L�}���J�o߸�sc>��鷺��K����Z�X�#���ӯ�9%B�d��l"��š���AeAe2y�8a�uxk��<L��~�䜾0*��c�r��z���}��
Ş����~����wU����tǂ}�;��|n�]}K������*E��낰�*g�L��L�I_}��I�J�ALZ��Aa��@�/vO���ڲdS�C�g�W0*O_}��)<B�>>�3yf�*��vm�|�T�W��`������8gL=Lï=��t�_̝�}�(v�!��t�g:����	�&eg���hp�R�c�3�VO�'W�l������E�|@2�O���	̋�Ϛ���i�2T_�|e���g�N}��r�ɓ?3����
Dd��|�')�2}��;~L�\�l�<����Ƕ�PS���'�&H<���(��"�]��/�������g�M�
�_����:|eH�|���q�'=Y�&C�CĬ��k�O=�NR|�J������AH����+��AeN�����)���g�I�Z���w�n�K�}�(�	#�t��N.g�T=C��:��fz�b�Xrw�9H/�;C=_1�;C����yg�r��H����>NXV>yI�@�*%w�~��$�T9>����$�O��CD�A&�NBT�ަ����yfz��z�a!�+0w�0�!��N���o%�05�6Ż���� i�Һ+|�<$��8ꕲ�30�!qq����]1��I�QDe�����-��8�gss�eNã#$���Cp�[ؒQIvr����
��￹��{'h��N�o��P>O�+���a���NЯi=��Xt�;K�x�g�>L�{�3�� ��|�&C���@�����"ʃ�AϺ}�"Ͻ��]�NZ�_C٩���������I��X8zJɭ'���� ������fH�z�<Nm�o풲rq}N�>L���7���^�2g�����
Da������ ��;�*��e$x����;�^Gӭv��}�z���O;����NX9��xS��&@��gi��N����3�2L��KN�� ��������"�����Ι/6~d��4����k�:�z�� A|>��{�W�fNn<{��9U�PR}�pv��Ǆ����哗�O=�?��!��'����pt��+�����ʆC�ft["ΐ�Y�8-;N���ӆp��d��Q���� �X����^�7��μ���9�:OXV?=��8@��
���ܷ�$�T��d���A��x'����i�>d���}��O̯�
�~��<zI��ά8AaZ�O��x�|�(I��R�u�����{��}���+:O��8aS!�z�I���ωThs�8@�+'̯>w�퓔
�C�18jVO�'�{��A~~d�>��:AH�|�:=��$���>��̉<}�"K#�|[�T��";���]�s�������L�s&G_�
������d���͆����d�i�P=rO}����3�����'�T�'ɒw��2��2);z;�r�̏I��@�<	���9Z�H_ʭ[��]qg�G���`�'�}��"}��Ԭ̛_^N($�
��KC+�����)�O_^fL����ៃ�q�_�
ãm�z���t�ھ�d}��%uh�ҏ�:�����k5���A���1W��t�^t{��L�!���p��ɒ�^O��f�O_^f���T+8�g�l���r
E��'2�H�z��9����>d���������w�~|=q���'l�l�����$��'g�i9Aa��:�i�T����~��L�2A{���H�(p�!���Lԋ*����+'�Z�}�d
�:�����A��{=��8��z'�.�n��=Y�k^}�Mq`�=M�UX��j�Ʌ�5�m��m��t.ۖ���UaL��]�L1��a6m���_k�pH��U�w�ʙb�lyYe&��Ӻ�n�P�gUN��\4�ͫt �ʬ��w�^Q�ޒ���pb�Z52p��̌�~�4ޥۿ7]�,L���6��Saֱ}XU&�uQ��`C2��%����l�,�n�;4fT�/�Ќ;���ώ�-/���E$s6vf��_J�9B�T�b���	�2
:�c�4�u�O5�j��o�)����)�={�w4�D���S�<�ҭ�r�Y��c	Ԅ�-�{���F�<��a�L�PJ����Ew+��֭ ^V� �۾�y�p�`mٝ�p&r�0u��������5)�0�Z�V�s��Y�u�{yB�;}�Ql�,��&�e*Ya:\Wu8��9�G���6�Qt��q���� |�e�4�SB]�\�ٶ��n�c��g`LpAF.J�s����Lꗯ���"k���9��B��R�"�3y�NX@p�o*X�	\���;v齘o�n>΢4��S�ht��)7ь�r9A���+��Amх�'c�S�I��QyJ��;�2�ہ���˖B�C =M�("���&�Q��e]�.��U�],CD囒��]�.8P��wQ�6���]���[����`��6��H;��.�:(kEL܉X�zN�AD	�%)
��|�_%D�w*��{W�ZÝځ��9���+i�E��~T�Ԩ�;g�^���7��^�䷣+b�[��u�e���ҽy4:n&w3+�uݫ�Q�ז���U�;HLfn�������VD�8y�v���9�[+>�	k7��o&�[*c�a'�/�q��"��c2��˕e��+�ҭ��{���,So�����
z������Ϸ�e��p���(���
cc':i�7ݯ�V�-c�w%vM|ƈ݀z�ow��Ǉ$��N�5��p�Z5��bs�3lBz��8��}�4�BIcP�Փ��A��Y"����n��Zc%�;���i�C�!u�d�j�5F�zi��G)�t�3z��]�ń����\i��Yr7en�s��r4�FN�ȭ9զ�Y�t ��{C�@&m\�zoV�3]���TM�\�y��/h�����~���(��(�wԪG�T2����X�&_u���;(�f;C	���qn[�����};�eeo�;;�Kh�"�:.�D�`%����շ�n �:f�i�mF�^C��C+,��&iZ,��W�����E��6:��VǴ%�Bb�"o��q�k_TWY�F��L�]q�eay�:J�2���S�Q�H0����)�ح�/��x�S�1�������Փ(��N�K7NGy������dj���\��I[�gu�3�,��75���Bt�^��-<:vT�9�`PQ�d���\���ډ\�rU,�%�Q�զ�ً��nr��ե�X�*d�[]b��mF�6j[FV%��[Z�ch�KX�\�A�76����ب�آ\\YRg+���u�h#���ŤYVʚ��&j*�ۆ�]j5Z�e���S0�%Ȇ�M��*X��7����le���b�][K���U�R݁C$]D�n�-̭B���ح�DT2mVTMm�b���7k��r�+h�\�T
���L�к֨�s�5֒��k�W&I���a�m0��l�k��k`VWjUKvD\"%d��TQrZZ���XQ+[mJ���+�F�Q�k�%�f���5]��-d�E�1p�f��Z*��̨��QB�#Z,\4a�R���q�+
��V�k�`��j8�i��6-��j��*6�-��a�����L>*� Tx�ה+��o9'!� ��n-�w	V	�j�Mh
�v��o+��'F�v^g3i]��z��x�Nn����K�<��ʮ��㵍�� I����~r
E�s���|���%N��'������~�AI�퓓ߺ����PR=o�t�� ��{�<�3�d��3�rO}�E�	�� �{8��c��U��ݩV?Y@�����|sI��|�$������כ�������ę��"�'�`�9g��Y���NP;Jϙ:��^3��
��}�r��
���a�Ѣ �2�N}5�.ʗ��ƅ|,�+�=�[�g�gӋ<O��=I^Xu�Y�*��4� ��+��c�9H/��{�<C�t�P�:�௬>C&JÐ����XV/�7R}� "��k��*�h�޺����}zJ�l��N�Ӕ���9��
EԾY�h~g钰��<�������8I�>rO�W��z,;k;�%H,��~���Y�f��~>�"� I���sͣV�Һ�w_�~���"ʃ�;��I�J���4�ud����_��yiơ����Z���Y+�d���3�K���p���g��$�
����zt�=�@���v&�kҮ~�M\\�>�����~dx�z�}�I���I�[�y�Z������
�'���X�&a�P�*A~g�Y��t�`f������"�Rz�3�K���Ã⣈���g�yϚ=�x" �+=C��:����=B��<�r��gS�w	�'��;���%~d����v�����e�C�~N�%{N��p��ʇi�i�p�Y�9�g�D��K'E����U��]���-�~
��坡��%za�2Vtʁ�V��^s���&@�*v{�9I���a��;�9AH���w=� �P<KϿ��N��>d������'��@�
#�}&H��or*��1�]��v��y`T5�P��*Ago&��V3�d�!_Y�|�3���A}H�����%@�P���3�y��2w�;�� ��d�{ǜ�O����߾�Dt�H�>yw�������QYW�Z�]���z�Ù���S�ҹ���;`p��+�t[��ANN(a�����,���O=�+��C��0�C�����>B��>zӄx���I_0��9��NQ:��κQ���l���q�4T\�ɝ��Bi�}�'6�_�G	����ۻw��:z���o�� 5>v��Қ�{�Ye�Y� ���8]Ea��,R��v�������=�:��y��ސ�@��ޥa��X�9i&c���_U}@ss��S���D"<	��͟�zΟ@��o�i��<I�Rts��fd��[�'%g��l8����=N�i�p�U�^x�$S䞾�3��fJ�½�A�| � ot?��/]>���;L�i+�߸���YP�{����Ag�w�㈳�&`w��a���!��h��C&J�2�*qfO�2�x��g�l}��	%} ��L|���m���������q��d�׎x7vO������dS�,��_����')+>rNN��|`T�}��Y�T��w��,3<L��+Y�z��Mg	�"�Kr���N/�g���~ׯ/_q�;����}
Ι�vLÆd����qI� �ox���Ǵ�l:L�2v�v�O~���2s���t���8B�o�I�g�g_}�H���2N~��Yd��������x����պ���?~���P3��a����IPS�*zù�S���S�{� �� ���|�����{&�C��x�>����������s>d��A�
�W��{��b�2���|����߹���u�T��_Y>� �R�����X������ᇌ+��=O!���Ag�T��1���z��1g�=L�~�>���f|�G�C��>$��7��L��mem-T�)1$x�"��O����$���P�+��i2"��9���
E&���q���39a�9�������Ձ�zϜ���Ǩr���	��>����._��]U���3���:a�f��O��̊T9��x2����8��J�S�x�t�ϸ�d�&L�_�����i:B�pqL��d��#���p�2v�w՞� dA��5�M��Wo{c軜�����2z���<g�y�}d�3��~ӄ����d=��3�F�?}�d� ��>�o�2Ak�AJ�O�[?'	����p��T���Y�L���	>�f��H��ڤ�����q��#���� ~JΘu��g,�į߼�̝u|`Vw=�O��+%W���PR)�NO~���+%y>��$�Ӧ��,�<��'ɓ!�W�A~�_���u6b���$6�~(әU��%�+����uǁ����ݗ1v�"Ш�n���fD���ue�8��_��I�z*�J~f2���	��%ϥ�V\��Să�g�N�YKۘɒɴI]�����J�v�`f�����׈VJ�W9ݫ� =�uy����G?,���2AO������a�l�!����ݜ������I�EԬ��pÄ��ɘt{���%|�����'T�ǁ�~s��9>�|4�����O��њ��qzWFv�ͫ��~��{���<@�6�p�_X'l��a��P~8�����Y98�3��a����R�"�7\����I���3�i*G��
��+?8��|���dx��Ͼ[�ɫ���}�������z�I���p�2p���S�dҦd��:��p��W�u-���I�3�'	�?�R#'ω���3�F��_4��8H.Iϕ���_@G��y0�l�T}x�o�Y���AN������x� ����9@�*�~����<0�����l�3�r[�(�gL�7~d���|�ξ0+�6��VJ���=$G�:_/��_o�a����tf�ה�ʓ�֯l�{N|¼�����'ɐ��~����*:=�q*��d�S��|�b���d��0�fd��� ���:��8J�@�-��
>G�zO��w�x����#�Y��|������C��
���a��Rp�AC�u�8o�AH�ydSyd���>��J��}��Ϲ���������㔟���
��텇m`�Ĭ9=����L�'�'	�ȥ�������Gt~w?~��?��{���:C����!Y�~��?�Y�p����{a�T������r����!Y�ﴜ5����
u��8@�S�Nw�q��%@�+��q'����@��A Q��IY�qbY�n:���zy�PR#%y~ׄ��YN5����Ar��焞}C2u9�<0*
|��8�ğ'I�޸=a�iXv{����$ό<O�ϱ�Ak?$�!���9H�d��׎~~w�^y���\��y�w��ol��$�)��&����T*VJ����~LZ���T9-�����ᇈw��
���2rw�>I����o��9C�=L���i�;B�g�?&������y�~�_ϕ���F���|O����G��î>��:J�@�{��+
���<���T���9-'	*1h/�X��R�d��:�Փ z�j�?2��Rz�I�㓞������&^�Lޜ�g�;g�;Z�����n��Q���gi�-�t�����ʿvz̥h�`Kk���FF#vU64ܧ���j�Cu��d�E[�N$]�ҳ:���&���8�	vK�]�;�"������-9��k��xE��?��#?,�i�������z�:�`8gL>Lãߺ�|�$�'gq����d�����,�����	�&eg��ա�J��+�VO�'W�`/��N���i�~�ߝ7�z�����~����~J�!�Vv��*���2���g�Ng�`�_2g�w~�� ��{���Ag,����'��������O���y�x`T���8�YG�v�l��}�9��.-�}�u��&a�	Y�œ=���[� �3�;�N_�䯇���Nz��L�^�%g̛^r{����
������
�S�߱+��AeN�,8t�ΠQ�DG���~$�pm'Fv�n����$�8Om̝!85Y:C�NgԞ�qa<a�ə�$�?�i�NRNg���E�ׄ��<H�_=�đ@6�f3�8���ǛY�]�3��eǀ�'�Y�;K����xg�J��y�Ѭ?3���Ϭ��'�+�O�6p��v���C3�&g}Ӗt���/�d�|����c��*$��|���5t���ʻ�Ͻ�"����}y.��@�R}�8zJɭ'��~�$�2v����%Oaۙ�%d��p���g�Û�OP�l�3�����0�|�NR=Co��^w��{믺���^��*~�\{�YG���� 3D{Ϩf}�<0*O=����'ɐ>�Y�v� t��{`g�d���v�	���V��
�����Ι/6~d��9��8g̛_�\{�Wu��s��=s�<��_������'�T�>:����9x�Ğ?<$���'̟��=�}�3���:>����%|`^ϼ�O������["ΐ�Y�8���	��$I��qH�%lq���ݽ��m}�_�㏡P�9@�|qC��aS��:�(�B�����~�2J�O=�H�}`d<=��R�d��|�tϙ*�~��;e}`T���>g�I8B� Y�� ��'ݵ���/VEO����;�G�>�ReHTO(�T|�d����Q43��]�A�r�3`)�0�d!�vM��umu��a�Y�[�;��4���ym]��#֍,�W�Vz+"f�{7|UX�u�vi�� V�R��'<�7^^F��ڏ2^+�F�Vj�����/��D��Ĩ��ժ���'��;#�����f�`ut:ƞJ�uf����=�̍���<��
b�.Q%©P�5͕�c/Ǹ�C���>�<���t
����ӄ��U׷�����ᎿH�B�3�� �����sIN")C8�1�ؾIEVSW�m��ӻ�$M.�a��q�\��!�JZ"t�0�1�p9+����V4E5�Wb�.2��G}�4�'CM[�DW��ځ�=.,8 �	:
PON�fP��ŀ��{H����lY��}2Yy:�0`a���Ûp,V*#1	T,ݣ1��5]��w7��A,Las�Q��wճw�t2+ɺ�u�ۚ0l�n�2:�l�<�t�,uo�,Yy�,�1�OE���#�W��"+ٮ(+���QN �r�95���pOM�;�t�iD��Ę�5�u�>g��=��{g�X�Gh����g�,��{���\^N����6�0p�BJI}�7��*6B�9^�
^F�8��(�I=AQ��V�L�[I%�=���7dw@���u�mE_��Z�f^È�l���ȩ���u�4�[��;D�lΛf���R�)�XD�u���x�*GI���n�=C(L�عn�=�B�W�&���4@f���g�kI��w���M,�"O��|!(U۔z:��3 �����H���G&P`X�q��ʷ[T :aj�9��wiW J7ꯇ������Jݶ7��w���r�8U69H|�MV�g8^��� ��rB*�!�H�&^<뫞-I@Ss*B�Y����UIÙ�b��qvu�ncC:J2��$�wn�oY+�I�Gت��A9gy�8�*���dn��P��7U6�r�t�}<�'g�x��V�up��N��i` {��)����)�;��D��{�����Zs�]R[�����c�
�6�t���W��P�5_�A��l�{����	a�;��gpl�M+�ъ�t#�P��d}�2�)6�V�[��>�=��I�M0*�-Cp�a�����<x�o�2/�ų�q;�����N�1S�����z6X�\X���N�d\+]�²��tN׭�fM���F۟^��h���Z�s�ZA�0C�����ؠ�����`K�Ҍ�9Јf͝	۹5��0�	|�o]�oam*��E�F׺|R��θ���}�H�7���5��}�=X:h�w��yf���.�	[GwB���1N�.��c����V3Hn;���qSpl�2Nv�Oھ�r/F��S��*V1�|s���g% u}�z��N�ɽ@�4k�����*�eG�*�u��8�ʾ0��)'u9��(�%��+1�?��}U�U��(�+���kUV8�YD����g����]��H��'m�Z�����s��Z���Z$�fKq
3��M����'�.b�:d24ѹ��>�	R��=Q#z�[ט�sEZ�<�z����QA��LPNX4Ҋ\��`�OI�l6}���ɜ�-�z��Qp�P�4�f�$U�67���&�W��k*��a|)�"���[�#�Z��\D�al
�#�,�#+(s��A�y��<�>�>��^�T��kqj7z&H�@M�qf�q�7Y�F��ȷ>@��{agT�F�IgT<�Ym+΀Y�ޛ�n����Lo�v���3&B6b�%���X�ʎ��Ed d]"1�a��dlLp��ޝ��r�.޺���?el�z`���V�����V�y���G%<��̍x�ՙo����;��G��5�)�r��8�E��Q�J���pt�B�kg�������VC��RD�IQ���p�n(:T��(U�`aiB����;n9�	���Wm�cw{د~ò�[t�ǟ�k��q�F�g�r�;�u��YBm%W٢��4�`�%���[�dC��^��"�N��e�+p�s���F/���7�gV�:��zľ�󥾖F������M1j�:����+ԣ���~x��5����c�D�������Ƅ̲�L���g\�-�<Vƞ-�m�9�=��D��؋��z��B2"߄xr04��%Q$3^��b�A�󚽍��V��9,�o��2�x��u�,ۊؾbv!�rI!H�6
T�s�rJ�N��ܥ��˾���Dg���Y�oR�`��>�Y&PA)W�� �p'��
�[Uv�p�ܝ��}��UyH�.G��ۋNݍ�nx(A�)�)X2Ll"̑�,��>��t��Rj4F)w����JP9Ğ	�臀�Z�vsZ�F	Ynb�I	���ZJ#2Fh�Ge_s�a(�OuI�0�a���!AG)�%�|��NX-��fw���g�߽�\�Ɠ����(/fUB!�]�~=Y!X�wd-rK�I�Y����<����N9�[{�d4Y�i�u���eX�<mTa��Wr�u����cY��ٰ�X�,I��e�6m-ܴ ��1W��D׆��5��v�Na��&�g�H�f<�+�yc�A�N�Y��K�q⚩f�Q�(;�x�h�sWpy1�YB����M�kmTs/V$et��5*ִ�G�x��#Cd�NL�#��P��K\.H�>ڽj����敖��W���L���7��U%Emr�������� �nRO[쎵:3�5�t�c�+�c���6'&ص]r�¹��]�_G�ܱ�vUqOwD�^���>:�����+�2�������n0���㏧LlYGI�
�n�t�lU;y�lgF@N�����{��H��T�8J*®�x�QO_\��)��R���eN��c�$3�>�#�����YY�¨�ΒYv��*�;��\�;ؚ�۝0xf�GҪ.��U!�5͕�c4�(�.$���q�\��RޘU�d���{��Vp:����J�x������4��R*�{�ഫNV��F5#�^�);�ց��wvB;���$��>�m�ی��AJT"t�0�=�5�Im�����B=��v��n�D�q�8'CMrȊ��j �����^@���g7�
����)����o� x�:h =��*J��r�8z9^N�X���+
:M;.�5O��Wt��hfLB��L�zb�P�0��^�~��Ƞ��0�����9���,즚��Vث
�Z�+��w���w�u�v�Ï�p�]���,�O	Qdt��f��Emܤ;�U�5��DG����y���>W�ح���c�n����K^t����PK�ݯY����B)˺�t���dܬ���1�{[�~x  ��������[hY����M��BWS5b�q�.�"�\*��35��uDէk%���n;01��w�n���Ϫ�܌�[<x�x�1�
��o�TK�Tk��&el������IG�஥�t�5d�d�"�-x���]y��Zԡmʌ���
s|�^�My�)�Ж��^�o�e�rY��:ƇGϹ�B�&���"�Q���9@�bw����>�䰆l�zWnvz~���Q������K}���T�~7|������M!����H���fb�6w�(u�y1d�&e`u+i??	�&�'�v�ظ�o�+�Z�ߩ//'��*�H�эT&W���K�|��@wZ�5��r39���9�]{i-�~�L|,��u	����q��y��0�}�H"���{�W�ET��<&3؅���*Dh��</�ܛ�1ub�BZ>y��՝0��
�!�;{�e��ewX-S [$�%�З��:�ux�)"o�]Q�=I����D�wV�L�3"펎�Z0�$��w#�;�>�p�"��][�>���三:���{kC�K�<oh��aB�>��J��ҡlʹ\�p�]2<��2�����Y���ptCd�M�x+��N�;�
�p��"ܤXc,S��SK��|�;B��#�If���y�1S��U�fݳ��˜)�X�mue(�xl��Ь
�r�f��e�'-�C¹#$ҨvPfV��w�����z�7��[�f�����8;ZYx@;� Z�[t6��V+yމ����)�si5.�M�ۑ�Y�i�X�<.�l�X�B�Q�Dh�A�M�87��{�PuɁ�V���[�%�7�u>���ϱ�NZa��4oz�b�&ō�ݠ��n�Ҭ!��7��*1+0�J���nm�|��$�^��z��Uq�\�ST5������:�äw\��k�h%}�u���0�Em;�M�����	*� ^��[h֬�z�h�Os�YU�ud�&G �4ɔ����Tvm%a�:�wLVY�bmnIć��u��=�5j@o�e_yQ�i^J�е�&����z^��J�O�C��ݸC�*�t)���iƚ"��[A؃v��������qԛ���A%[� �Lx���ӈ �I8���J���/xd��b�M�lU�~kS��m��+�������RP��Z�U����Z�ccEۡ����hP���t�L\v�:J�P�%��avAm�:��@Q�����8�6�e%n�N�*!��kc�U����l����q�]�G����K���o!����* �]������k����B�'gL7�l}F��3 9��d9d^�y@
�
K�ͼ�"���B��Y+�&ڼ{k��Ų��+�@�
�N���9��B�}�h��J�ڱ��^���t`�Y\���α��3gX��<�>Ysk�W��^�݄����0��Q���ͼ�.ZT҂����E�Y,���/,���4�+����"#mp�O�Z���]����G�W�w�c�seD�����z�ehՆ9D�`�\y��,[z���gLW��"�GIOs0���c�@����f��\:�{)��v��W�
�o mX�� ��CG�pT4v�[
��_�;�v����	��+�fû����SF��4�u�����M��\�]]$X̿�r�p[���,Uۇ���$�:?�5���IT���:�()���dm���e��Q�{�;;N���t�I[`�dF̭�)�'a��1!�b��J'�;V�w"������řB��wf�iC��@F���,�w\*������SU�z;��\Z���.uDԾN1]xE��� �K�>@�B��B�k��T��a2f)��\�̶̪�.�֣Z)T�ZZ�����h�9k�r��(S%Bڪ ��B����Pɶ�Z*��5�T6��(Kl��P�8�Qr]�
��W`���ڊ�l�.�T���#hfB�-V�F0��Ts�ЭD��s]��[iR��%����m2bլˮE��[��%j�d�R.n��bȍj�*)Z�J;Z�(�Qu��uLʆZS[.��#kk-�Z��53$�+3P�Ƶ�䴠�h�\-��"�E��L料��]Mhkj�L�v�$��֪��b���
�33��R#fQ&�ɵ�̙
�4KnE��s5��iF��QJ��"�iJ�v��[l��aRL9����mZR��[V6U��m���B�TX��봨cPu��L�δȲ�&n�*�%[k#j�j�ѴKFإb���2QEUi
�(��wk�N����O�l�R�N�d���C�<�[!�CųHoh;�@2���nf�b�)�K�t���'�������
,#�y��ag_���o}�=�S��;�0�/%�N��I��w�Gg���A�W	-m	��:�K�
ǻ�	��|��.�7���=�α��'�&:����
z���uX�ҿz�x����gDs��k��/�jሷ]c��.����>�Z�=�}��%�B}q�R����}Φ��-W*�n-�A�*uk�����O��;;�\>�7�w8����6��e�[�Eכ��A��u<��ȉ�g��=�����e{�a%SAc
i6%�u�������C.��vcWF��g���D>Ւ]Z��]kXsA�)�Ж�\�c�����]�',�E��}n9g1P9��C�'X̎PU?��b��S�+����)Mi�Zʜ�A��gs3!�6-��գW}��L�;�<�=�Tm
�[X�{|!��W4�f�t�Ku;�@"�O.=\cJ�q�]Xme)�6�m�Cȴb���������>Ʒ���}�mu�"�\(�&��'�IҖj�K'eh�&(x����JR�宴N���-��}��"��댛�)�f��j!+�_W�}_SVx��/!y���ݍ�,9'�/�znv��2�[Y^}[A{,�O6�7�6�^�� ���T���-�f��׊uo��ڑ�)D��vcY�]�ʌ���78�^W;Q����ۮ&.ì����݆h��$��8���=��8����A�n���	>Q�׈a��jv��c�躗ؒ�6��)��a�u���4�T�7.ex+v����j��#�tb'�хח��� ��iT�u=΀*�aqy��՟<=�!���L��a�>�A[+|��ߒ�BB�;ϬP[>�z�q�F��>����`�u�-����[�!�;Qb/%$lq0��ˊ��F����z{X��Y��J�o��r�ÛaPq�
TF@��.�uW-�5��us���r�P�j�3�.�5���E����]�/H6T��G`�����ܝZ׌BͲ��y���+����}G�+��wulL	A��C���ﻋ��o�t�o��-��ٹ��c�O_��~����(�b�B`ٯ1��7m�EKޙf���q���_�/Q&����'��]v9�{�ب���9dОy@e��ת�IT��g���`����Q�b)�����aC��u�]W�#`��Q|`o��^�kz�����6� ����k=���G�:���Z������ru�_�ޙ�iI�L��Sn^$�����xs��\מpn�"��V|蓐y��,��C�Dr�Kݚǋ^�ٕ��L��y���$�������Gn��'1�i�s[&i�m�X�_>4:_5�ro��ݷ�cn��=W ��K�0yoia8ܣ�}x�V�_l�3(�R�����'M~B���-=kgzCUk{k�G?R& /���t&B	Y|;
���&�0��;��bb�n�C�G<Y��.���m�4�D
�ӄ�	�����M����0s�i;
;���D��q�Z�7}���dkHׂ�
�?3�P離�F�D뱏�"�c�L�wc����7`x�<W�O���D���-�>�1�O�2Wn�b@NnMq��Bu�������\�V��i��&�p� �������X�7���}�4"�*�D�$��s��}�����E���uv� ����2i�E7��c�����/`���v�W�FEU�u��ΰ�r;�
I�*�vx�{���q�����C��ݭ��dZ�N)�i��8
�fs:�aPI�e�ާO,C�f��*�[�*2�v%K�X*�޿���V���\��&��.ڕ�:9����R�K�}4��Fw9�oֺ����=��מ<��֏J�Ul�+�cKH����s9�fn�?rQtL`�5�+���>�ٖ%<�e�0���{��$���������Tז0�6#|�tX�g��VՓs�P(e׍uZ�w��Ґ-���r���K�9O)MА��+�I��WuQy�j���h�L�n�Y����u��L��ʟ<��<[�݌��݉�j����:�0{.��^���-��G��;��.	�O��@���wk�FS��؟X�as��g*�l�*�)X��s?�^�����F9}�V`�#M?o��T^�ջg��]��ǚe�M{��N7]X-��f;�u(T8�)����{���m6KW�.�2�酇��l{Je��4q�y�+n�ҋ��}�}�^��kJO�%�v��U�~�jP}�`��BF����r��zi��^v��H��8��1���^X�{�ތ援�n�Z�[��[�4���ݽʌ�B�ok	�NW4z��{��H��r�Lw[��ynԙۼǫ9�58�2E�����apM'~Q�׈a�Z#C���<� �N��{r�gA��i�JTIJ[Αte~>cW��U�\����V� �iň�w�	��'[
WpV�9��	��p��>��.�'���cw��L�R
z���n+�m�����Ko���d_8�q����5��nWEG�_YV
PR�FǏ>����>��5�pLaM�&f.{7Q��l�.�'Qt�㲬8�t��j�4%v;�}7�k9���n�Է�fï>��$˿ĵ�u��0W�����׈@���^����\v*�����f������"�Fn������ �ӫ^7��KY�F���3�<�&���ra���,sx��r6�k�R-�ӭ}��l��@�T�JW\�vJ*�`BD!u٤7��â�'Vh���u)�!'?�����8O�����u�e�Vs�a%R��<�҃:����d\�7����9�e����.�d�#��R��蟵3���=+ 9|s\�k;բ3���'&�[cΉ?g��*7��F]j�;�~���}���d@����kV�h�����ܳ!_������Z5uk����χyI�c��Y�i@��)��ڴ���3������,PX6`��Ps����Oy��ʾ�^�<�K��Uhה�;S-�U���l=[b����W�&�����0ꇼ���z=�����*o�/�78�W;Q�ͼ���W]앷D����1ݒ��u���2:o��Û�m�r��(��ل{�E����{�! ��D��r�L%^�i]Ej��kw^�S9+b�hC���K�={���μc/%����d�zc������aO��ځS>~�3V��K��tn�}n��i0bj�#o��<��)i'�窗�b���gSO.Ɯ��6Ý����na:d�w�N9��s6���8��Hlp:j�g\tq���Փ��b�.���j��1��Ͼ���V�@��A��7G~����lao�l�������T�on���%�]Y ������ﰯz��<�r�a�4hB�䤍��k�fӵ�������⡻]���4���.�r�aͻXqJ
Ina���*v�Y� ��zsr�[u�Щw9M�a���nq��txt�	
ec�rd��P����v�ܚ�VZ��z��*�9�M���K��^��xɋ=S�K$z�X�
���ꇢ>۸�y��^���,�"l�<;�n��٠���7�+7�%o������읬�$l{���M��*ߦ0\��{m�.����CSe�<�!��W�g>x![��8+�d����֘�ìZt��L��ʟ<��^����e��$�V��P6�i�B�0�9��Y�#���rUOq����/���^�M�|�9���GJFMh�T;LL]��� �Ml�+Ԗ;}���BOP�E�KG�j0��|RLw=�/�cl왊�mNc��R
��w������v	��ӏ$�� �:=���.�r�ɲ��l�f�F�v�0�A����6cݍQ�ٌ����K�tm���"j�s֒P�vr���¯rg�����׌s�==^�P�����
{�S�j��ZQټ���W��"/$�!U��*��W�&T����P�|9���0_p\��;G�O����s�ߜvu�[
Q8{}�2�{��}���8��药$�~��՚���0�&�����a�Z#Dz۽�H�3O���]p<ן&�m��W4h�o3���X��>��S�c����0�Ǝ8���MGLZ�HY5��+�+y�'�V��{);�c^��+���
饸�^P����Am���$ҿ���I�θ����,���C봚��l�WIK�~)�ԭ�	�d-�r�|^����Jw�P��n�p��#�:�����\�V�r/oo�=���t���gJQ���MD\���ٚM��J-�E��X⺟Qۘ]�r�q��z"�W�,����{��/b���#�Z��8�;��n�:�f*fewl��Һg���ͅi�G�=L۶��#>�TLh��[:_����D��" �8���wi�-+˾˛I1)"+%!�ư�n�ݎ-�&�z�Jb��ku���\��O+�5��H�}_}��XQy�U�wٕ�s��)�&�KHK�5�C;�.׉����	�4�켙��|U�*�o��r�Ս�}~ZÚ)Jho�D��9����H�#�f������Ϫ�\�9C�2�WD,�/S��s@<[�ʙ��_ɓ]��N�����L@]����*����z��G��;S<�L�EԳ�ہ��޽|����37�����W@��K��%���'����{c����_u�k"�g2ڎ{�7�޽�����`��0���݆�SY�F�[KV)��T0V�JZmӕ��vu���H� ��yoi�H�����8���3�ze�X����h�y`c
SI�Q�׈a��D�35NX�eDm���c�f�И킹誏\�a��0��tS}N9u�uV�/)Gs��眸a����HQiP܇�{�W:6j��Gꞣ��{��qh�~�S^߳�:�4!�jj�T���`D-�e_<V�E�dU�K�;���������$s������VgܵED�6:^pֶ,���ScE��
���ۘdAkC3�G�X���)o"�;%�����7��V�H1�X�9m.�ߞ�� ��S�x�8�ۏ�"�m��]��YK>�+mO1�iGY= %��K���1#y��=y9���̡ʜW�=�~*�J
[�6��R��ۓU�qLWj[�$U��m��b���`���vӘ����VWAJ��ծZ�f�EP������ح����}��2�ű 5�t��Mc��}����d���{�$��K>�K�$����$݃���t�N
�Y��EL�N;���uY�o�������#k$lB�C�p��W-a�y�)��*�N%a%r�9gW1���ǰn���G�N�#`���~#�����W����b�r&6/������nʚ�κ�B�9��q���nv�<�P�A�{���i�/��]����dO2淋�C��X�Cf���F���l��aZ|���b�Hx*��r�ڙm�}`&�l�cf�`<����܌׫�m�7�T��qR�@�3"��-�iw]EС� Q�ۣ�DY�*�K�06�
�&wt��i�`��!V���l�S�޼um^�[�_ύ���Z�Sd�cIG��7v�!W�9]� ��<�0k.N�\��U
�Gw����)+�C�|i3�d屯tVr�1Ь}bx.j�t��R�Ov�v��
�l�]O��x�+��:i���s��:q� ��3G�ۧvR�wSos	�ۗ�ƐEGK)�X�,�ڕ��*ѾT�g�զ��;���:�Y8��Ƶզq���e�]��5���NL���p�,8�t:���g-�rg)I۪=B�d�W^d���$U�u��3no=�e�F]A��P��t�W[�ǣ��Ѵ]�h�!sF���M�i��kn�5��7�cɡ4��B]Fh
��Gm��tm��:���V�:{&Ʀ\ͧ�l)�arTÜL��m�=z�lgNL�%��,<��5��"�ޔ�Q�*u���N�P-�{�'��YKM@U̡�NxhF8	�l�>�%�َ
i�q/����b��Q�|�#�"���/+9��Z�&nE�2��ˈ�2���$�:Ee���yE�|$�)5�y��ȯ
��v�5u�nB�Z�n��K�nظ��`?,�ܔ��~�,*6���AG���mc�(���[�}�r�ɥ�r�ɹ���9��]6�رyѽ߷(�$1ΘOU��u�F�^�P��b7B������5�ΰ:e*�B�V�n]^���*�6���V�@� �J:��wa��Sݣ�;M� 9$֡���(^K��:����\0k�Os\��#�.����P�<�� �?m��&0�ލ��|�w"�����<;He��K�e��Hp����N_\�4�K4��Ҝ���oV2^n� L^����Y��Ri�Ua̕�®!��cv"b*��x�]"�<��YU�Lk.U�ܮ�\��P���i)���W8�����:�ܣ#�"(ɛc3l���K��̣%�̪�s�>ոS�]:Qu'k�è�3lQ�Ѹ�W���3�	�ep�dz��	�����ը|�����uK�%�N)�HJ��H�]L�Bn&Եv]M�mpC��wH��mb�k[�讀���69R���#�]H������b���u���u�gme��P�nV^U��W� v�P��>��Zl0�
�صvV�:���k%�twr�����,M���w���=���W	m�&��N�Z���\��m�u�.�=v�wt��7h�nU��*�Ӑ���jFa5����+�>ں�8'M:�qj����w:��痜�<U��08Q���H�����(�V�8�����i�>���!�e��nK�l��t���rM�B��,;;�BG.��F�p�2fڛlm�Ef��sMg��1ܔBH��XU��7sl�w��k�������؉B���X�+9�� �g�1�UͩD-�*lmQ�ґB��.j�SV��L�ّ��)�!S4J��-�v�TX�V)6*��KV�����
$�E�J+�5�eʭ�"£j��]k��)����\�F#rQ"ɭL��
V�Q���R��ԣZ,�A`��-�**�P�1E��֭n��J��2�K�EI��U�PDUX���Kr[T�1UAEj5����rIX�+#n��R�b�-%TYd��VU�����ݩ�.�I�(��(ȉm�d5�dJ(�
�Ajd�ւ0��kB�`���R�b�Րm����6�#���m��6�����
"T*��*�Yn�d1j*(�
"(��PY3+V
1jR�ے�mL�H[U"�S2��A ���\���1_a���#{lZ�2
���&�����c
���3vo6P�Y���xɲͫ4�u	w�`5.lEi3�ᥧ?�U_}T6�<����bJ�˯N���J����.n]6�q�ԖFʓ����УCZ�T�z��HՌ��}BPKg��u@_n�6��Rs>���e�E�\{	�#��Q�t�t�w��Ba*++W7���Q�{��%�0�s5s�]�l����䎊=�KJ�9;�%�''yE@���Z��ά�;��`�2E>qBҰ�����L˒��󕮯&�;���Z�v���m+ �թ�S�d���%��i9כ���
�Y�]ͮN2b�}^at��aPI�e�.�]��t��9�~*Ç�C\�Jz�\�c��.
�1��j^���;�W�s�	�,6ؠ���J��u��1�tF��G��yru�߲#����⼠�I�п^����G��oֆ�B�ǵ�^�=��E����.�� ���"��3L�ܛ�\2�żR}~�
E�D�kĚ��}�F;�Ս�E𭋻��y��g�%�+�=�zF�=����t��J.	 �l�xe<.�;Q[��� �����ӬWPPfe�u=FX�6��Tj��4z+Ok�nV[���I��]}
��Cp�.?}��UL�إ'��̭_n��!	��b�������S˅F�nL�B�UL�x� �!;���yk�Þ���B�k9'W�c�7Uf,��y�)QX�����#�Oc̅9�~5羞^!�%�T6ye�N��8C^jQپ�quh՞���v��臜�x��v�TmqǶ�m�-_7�ut(�*�Iͺ1�BT�	A��_	I��S���`j���ْ�E���������^��q0���ɇ�%�!��([�UX��:�u��e]��I�S��lȲl�6��p��}[��Ta��,͘&մ��^�wy����/R�N�Q������R#D�FU���\��8�v��kw�[�Y��k+�Ry���`�2i�Ey���Y|��Ss���J\�r�]�$,�+S
Ww�u<ηN�>B�=�Z��n-�5��1x��%�����ֈ�U�����̩��{��xR�xVq��_ U���v�s�I��D8*Fe��Yқ�'����sP1͈����8�YB�P7ҝi�]�l̮]�
Ȧq��J�ܔ^��_ =�Y�Okq��j�/�~ޟ6�B|
�H-��I>�^kxy���v=�4�em-t�)Z~����.����l�hJܬ	ϯ�r�;y�Y��u����3yVm���.���d�q�'U�܋�վg���mױ�z܌�����5�34�QtL`�5�+���Cr2As�,V��vd]�ܟ��/r�V+��u4�ׂlD���tX����Z^D�g]^��ی����ڶ%���.ioC��9�򔦆���;0潄�t���f3!p{�����V��Y���.�tB�����\���bKn�ئ��m���=XC6v��W�:nv����_>v�y�����[��P��p!O4�B|�}>y%�Cgjʺ ��K��(>�*Pɬ4&�����v�5Aw��B\��&�<Y�Y���1�����B�X�췶��<��T�q����[�Wv��n/��a��6��1��A*;��/j�}R�.���ط�L��H.5;�q��:���_s��a����N���H�dv��i(��X�T-^�NV�w}b1[M)���>�&[F���}�}D�|��b�f|.v}|��[�M��;z���v)�q�v7i��Ԣ�6��s�Υ'�_�� �X�N�vu�y�md���)�ԧ��D�2)�1ʄ�s��W7��ݿc
}O�#�6uR���}���m-�ԓ����y)�
BKJ��Y^�l)]�
Ǻ5�nY�v��8�o���#��d]�j��螺`��u>�P[>��Nrd݉�ι�{+ww�9J��妃����{N�V
���Dl}4%k�V}q�^�1q4�wvjC5��cZ�-�v�I�]78�+��@�u��C��b����y1��<���gt5�3��.�bZ��,cX���i�4�$�@��+��r3/���ṟ<�)^g=vU4��5�ؐPM�6"0�ކ�T�}}ϯ*�1�j��x��y��'�N��{c�s�܊Xg9��C24s낅�v�M�f�=����k���¡�͍��1U�! K��1�5��!ݡ���*uѽ�Zsdsir�"wy�S�j�͓���ɮ>L-�
V�U�_:q6��R�`{�:_t�v�V��"�Jn=���/��}U�zЎ1�h�H����7z����6N�"�=T_��P�*o<�.�H�ʞS�������u�����z�X��ȩ��՟>�gh���eU���rfy�R�v��Wp�UM��7|������"p����Y����jY7����Ǒ}�d�1,c�b/��K�`)�� �_X	��z�6�Y����,qL>�w}Ϲ��ae.UKՒ�_/�7)�t�ss5�K��3w���T���d�WK����8/�J	VG_5Û~��8.���n�s��˦2u��ԑ0h�[��nI۞�Wf}�?{��d��s�w���Q'�T���{������I���2iA��Y�up�˹
�b�w���S7Z�Z����|ཕ����~JD�RZ���#dټ���j��LPJ}m�m+�w�s��պq^���`���%|���ޓօ��uu���u���ä])�Dս8��X�'������9c�u��mRǑ�<p�����ɤǐC�):�@���RBo})�؇a������GȌ��\1Y"����Q;�5S
�eX-��S����ռ�^�O���\9�K�H��Ti��]��t�*� �?;��{�W�(E밽WJ/h؏{-:��T�����׹�K�p�d��e(vڧMu9�P�ܜ�p�Et������"����v׌b�(^��ᾴ{��k�ͫ2��$��קy�j�>���2El行_����u�r=�y�iv�n�r���M}�q�����9�ĺ������t���F��'�G>OW|̥[7�u�S�f��f�^K�!���o7[F�qV��U���E��}2��ʟ<}-[׹a��fܖKb&l�ή�v�Sf���7;R���/��|�)��x�`_h���z��"i����d�Mb\-������l�>2�:��~�ۻ���i���yap�G��\��KU��co��Ǐ.�cTЂU��R�`c,u��hO"���q����Q�85���݈U����B,�+�{79(ݴ���oF���NU�h��[+�ͷp�}��ÓE�A��!�������Ǌv�XS[|�X�Cy�GT��j"�m�aJ�e-1�ܾ��)5����(U��&�);
;:�%��
D���Bc�8�����)��O��{9
56�2}o������v����0�D��h�Ru�D��ܾ�k��-�CN�
���I`R��=}٬d�O��vŗ�N2�ƌ��e�n�s��_�
yԅ���+u�H�<�P�{!��#c�I���-4S˖�Lf����߶�BAX��-�_l*�NAW��E��׉Z^��^G��E=X*�����O��{w�
�;p��U;��(����ceX.�S��1OZGub�Z��55ǀ=��#$���]��R�c3a����fxؐҋ��cV�}����ި��uӇZ��-������P��+�՟X�u4��4�-!>}�b��z��y�N�MM^=��Ṵw&̱*��Ւ2���K�Xs^)'��#�,4��W����iV����98��v��Q������LU���{��
Plk|��g���O�n�r:f����?�O@}OD��TĽV�k�����u��n�-G��1��^庆���Ř4��G�d�Y�nt���
�k��(.RO�^���&n�����Q̟C��%Y���.�X镼�딉�{=3}��e��ន���>��վ'ȇ��FuxL�+�~��VP~~�������P\����Z|wZ�������,B;f���}�%y�NV�aԒ��erx�EjU˹���<��z�����y]xƬ*�8S�⢶�V�UFn�q�_'�ȷ6�n>�ο�úD�Aܾp�k��B�"!rm�)��������} �{AנT�Tک�<&2�xX\�nM�0��p?r�H#u��{�L%Bc�ت�usy���@��w�3{���1��a�>��1�=Ay)�HH�S#[
V�:�U������-%�n����:��&��ܽ`��O��׎r� hyn��c%���ڮ�I�kv�K<^e'N*Ӳ�JJTF���a�����FW
;�a�֟_L�QB�L8ܣKgp놂U�8ӂ�);�7�&G	��=�W�Y���S��{���C���rn�gM�{�S�$��F"��JX�n�aV5��vk�Y��/%�R�;g)fғ�'bis�p�~���IsV[�ç�N���~*Î��";V$�^��Leʃڗ��2{�ѝЩwT׹&]�����n"���q"����EmW6�Rܸ����/r�[�k(g=vJ����4��h���&�5J����֠�X�
Z��]d'�
�j�H��������J�n	��mxr���}����`���t<͓px���4�X��e�>��3����5�S߇}~�g駝m���mx�ᘢ�2\85�F]�*r�]m'i��<�� ]-w�<�L�X�X��{�aa����&�v�Vc�5.���<6~�M�F���﹨�ێ�`&�^���r��Ul��U�y�v,����vC�|����=����|� 8n.�jez"Ȉ�p���ˬ�S�������sf��=���Ӣ	>UR���)�
�u"޺�j�y ^�Cc���%	��7���NC�s�]e��1���2+���Z23b�.i�1��XB)�l�8�lpbc��J�W:wnm�ZOQ\�Ƀ)d�T�<��������P�9m��Q�d����z�bP��� ���L%Ba�u
��PC�;qz�e�%��
�7Q!T}S{��U�g������4@=�|ZC*�E�K����׹5+l�l����%�����7=�m�.���e# ��G0�a1J�M���Q��Z�Am��ކҲ�V�{��p^�F�)u�z^��n��if��0EA� �o�M$[��n�t����GLk�i�=��]��Dj�5+r���gt%��|Z�	y$r1L�Q�9���W��e��Ql�+qC��6n�Д�Z��z�t��>�y[.*��%R�^cfi6$4�ν8+�� ��>����''z+��i������%{)�V;\�-a�y�)�����[ڵ�}��hM�?-��J.y�	�9X�����{�X�a칧�%��[�|���Dy�H��i�t���0�q����o<��}�@(���d)���}9��v���0�+U��7g0/�u��5.]����ؗkQ��Ī��F�[���D�Yk���ų%�w$jV0/��c��SGܶΗ�L�\���̙�MP�Ķ���s`j���[��ǲ�=n@�j�,�:�uE 2���M��*;�j��VQq��`�M��]g�ԕ[ώ�7��0�([yĨ�:N���T��������Hz���o�՛��j�v�Xb�v�=��I�Rw���]_h*�D�J��-�Jn�\�1$
ܕ�x�=ۙj�)�H#n�9��ь�i"�1�(�fx�+���Zz�wsկ�N̴����2I��Jw(a���X��\���e}���<�9,�Q�s@�x���m/�Z9irA8�MS���'�v�W�Zw��n'�a�Ϟ^���[��+�Z6a�^"k󽛲�A�ݛ;��&�Pt|6�;]Hs�Z�-_,we�{��[�.,�D��@yyƶ.���f�]w�\���e*Ί�9J�]hA��>�Qp䙸�Cp�y�T<�wJ�j�6���A�L����-ɱh.�nNw�uoZ4�rau>�\�@J}*t���8-n��9M}"�C���7+k[yb�a�Ls�ԓv�#�l��%I�G�o�h�I\hCAP�v���ņ֫���,��YW�� ��w�a��;<����Oq��U�\��䕦�@��w��D�ht��44+fPUT�A��v7���q�/�=��"�$vU�U��|Iv��x�4��bU.�0C������m�<ת���{ MԮ��]��Z5�JQU�/������h9�:�y�!ե��^m�&�<A�����٪�c�3�D7/;WBƶbb�j�*��m>B�m�.R�h6#�6�b'���rf�2h�r�����M�F��h�/��wN�MG&���WmМ�a��U�i�e���L���X��n�f\�|z�F��(�n�����f%��B{Q�{�ȃ6�ަ�
m:x�t�D��K12i4�h�Y�_w-T��&��e�0<̭�5<FM��sfy�	[XӰ)ӱ��Z�]c.���';�7�ѭ���zƹn�=C���wt���8�u��z�\������F�Dr��QX#�v�rR7��ө[q֧�1�����i�O�;�t/uS�>�<���;uى�Spf`��XD���]Z4J���2.���
��0���-3NG��fw��V�W=nF^�]�I��0��qM6�{Odeu��Uvh�p�zT�Y�՜�r�+�e��V���b����[u TNB�Y��s�:�r�[��Ve�\�w�R��tz;QN�`�r	͌7pm%y" �d�'3oWj�]��9�ԡg�f��ek�	�4<�Jۓyl���Cf�sAdNY[C7f}���k%f�w�����j�ER�kf[H�J2T�H�2kUւ�Z�Z�f�"%MJ��C�i2a*V�+
�Zf������kL�WZT`�-�Q��De���(-H�#
�����eE���dR*�"�+mR(,�U+�X+iD
�ȱE"ԕ�IR1���YF���Z�a��¤��-�P�Y3	�$��g1`�Eu(�!P��"ZU"KlX���f �m�2AMKR"A`�X�Z�E*(VҢ"�-Z(��R��hJ�*g!ABVQ�B�P�U��m��P��L�
��-����*([`��AE��dZ�Td*�XʕU%�m*����AX�EV,DJ�X�"��bϮ�賛V�l��n:�f�L�X5&�����bC�]��r<r�:��0�OM�2 �jh�5[b�jI���r�HqE(��[[�0�{�+>�V:em���>A���0����B�8�!y8��������z���Ϩ8���M�( ��꽚wm1^i8-ߩ/$>�,B�[ڳ}W��V�^J�TeeR���
z��C�~�;V���n���kő�¸�<��cUL>�A%�7��D�W)%�;�hح	'�ۯl�1��&˳mVߜ���b�ˆ]T;���O0�1闝b��_&�=�=���4�=nس���9�X�%��N�S]�ݬq��}�W=���;�z��X�����fͬ���iECݧ����w�'B8@/���HY"��Tn��.y+�݌�)��>�f��{���u�X!��r�!%c�ȶ�w�zC�=/S.zM�P9 �3��Fvf0w2�ʞ\9�`�W������L-��=��ز��'/E\(k�tɊ�w�:�WTΏ(��z�᮸Z�mZ�3�si=}bw{*����9�X��Ǵ���qCss#��*!	@]\f�u)qU�0�hJ��:f�}/2�Al�&Ц�����^��	ɵ�z�Ƹɺ��!���'�d'��h&���jb���J����Uix# ��*f˴�b�8��T��}�I��ؖ�[��/��"�>�JܿiG�.T��K�V�O@~/�w9�XM����>�w�r�Rt�U��Q���q��[�ý����Y#.�^���-a� ������Ի-4{8>��3�����2}
�_�Y������o��{'7Y�5f�M˚x�,�c/�䃊�Qq�'����ș��1�=-����q��w|�I��wԵc��v6�Xr|q]ޯK�)���OVnZq��Z�Hx*��mRo��L�aO>�ޫ^��Y���ٝ��.����X�v\��M����[A���m�W;
;:�{��~�C�왞�խ$��k�T��)+��]�	�aHM'J���kC텆��,�2�껷�n�Nq�31�����˄�Q%ev���ri:Q��9ۙ:�T+7�[��Hd.I͠8a���uJ��ڀ�5"u}X��W���� ��b�׹9�=�����>�<v8JTɏ)S��*D��{�;�[\�����qD_��~�.��*ʿ9ےe�����a��90YTig�X�>��U�9l�B����h���ҡ0��'[�J���w[�Vc;�wc)��R�.��� �$O��\k��~NM7�޷���d��w���m+�w�g�y��8/e�*�T���d�e!]�hvD��x�VLl�Jj�>��^K���=	�]���8��ګ�n���RǸ��*_�Ƿ�MK졖�wB໪y&Z-�t\Ne8�;9��$�뵽��?�>Χ��ֆ�DH��z_��I;a�)r۞��%>���o�Z��-���pS��}}dnO>�<��h��G��j��Ѥ�^T���r�2�=���:�Qs:�h�̅o.U�	U���1fw)f5�.�N�_���XO��X�g�<��d+�3�㏨�%�S}s1~��Sz���1�߷=�݆ŀ�d��� ƫ�t'h��Lb�����tks�x��+��L]�oX<�'B��$�J���T�'&<[��=m�\:=ku���ڻP���Z&�9m�"�l��[�����u-z`%)�J3$yz=��K�C������{_T0�Ȝ*��Yy��}ǥ�zg<HO�J;7֦����J�؄�ƽ��ڙm�U�{�^m�#��#�v�s�]
1�VT����=^�;��.E�Bo�7.��޴�r6�5����+�b���<d��\���*�����T�q�7����i���<1�xu	���<&2�F�T�ymV��P�J�X;�:�Ӻ���/u���z�̶9�}��v;�0�/%"4G�q��5T6�����ΰ�s	+�7�J��r�݀k>��(C�V���?$�Z��kr��Ľƻ�@���Z�=�x�]�z�ݫt��79	A%��Q���9N'ޅ�k'�|�ˮL܇ңA��4�-�v]�p�vn��F]]:�t�)Z7�P�aAKի\ԭ̤�;�W�s��8�<�lӔ��ʸ<k�dpWn����H^c��y)X<o��m���:%�x?M�2�&GQViۗ+��`f�4�C7�+�����I ��l�= �0��P�c�N����]Ǎ[�`<9h�%k�E�H[d�u��%��������L⛠�겄�]^nq��n+��GjD-ɩO(�l�î0v���\G���!���u4���6%�u��^c�f�Q۟G�=°=���������/�@"f��:�����"BhH}�qZ�]�[1n�)������qҜV<��9^�s�V�oK���9��<p�7wL.��Yܪ!;Xݸ�a�V*2cm��vr��Q|�b�y��<��8��̓݋wW�i�mI����`�9�h��=o��ƽ��ڰZ�l[�}�w{�;>wؾ��1z���W@��K��(>�1��ID{˄L˃i��v�5A
�[*IG<�kU��cn�� ��u`�|��L���+k3^kBq��$v&�rvm�O���Ĳ���'�YcFw5��q�6��q��Q�ɻ�a�^0�&�����0���h�}4K,^5��Z�˄�Ty��VF��ow��Ґ��bד�y?�B�l4�E	�}�m:$u�k=17�}"�L�j��e]�`�r��e�t0S�Ͱ$s��̐:;47{�2wr�cS����f�b*[��˭�G��?�l't�4&~��# �8=�@���T�`篻��)�FW�W�D��|���I�=@/$tP!'yԅ���T������
�'�i2��qg.k�+u���{J�������x�u���q��o�ؑ������r��L��Bt��ͻ �P
J^�)��ۺ��y�sZ|=��W�^��Wp��������v�5Qt�f�[��AJ��feZ���;G1��/?�{�>=D3�Q^�to��$��m��J.�L`��8�U�4�@s��ҏ��w�ho��9<@���XX؍�H.����z�J}���[�+�km5�d�O>�<���8D���Qz���̣��A�� *s���H��&d��8-�x�O�[�g(bs�Z��^g�v�CLOӳ�)�K����oW�DT�Q�fŪ��P����{|1�NFGtɃi�Ķ�K��u�M��z�X�7DwM�TMjg]_;�h�֬SF�о̪j=�"{7V��S�ɛ�-�V!��,�V�G�y�g��� ��Rgݣ�9b�t�X�3\<�X��P=���N�`��v��c�f'�z[���$}�3�ѕ���^T�^�	�W��v���Xr|q] cz��3z!
��Ȍ�Z�{�ъr�:�z�1���S)Z�}~M���l��V�D�AUnj�{W!��������c��\����-�i?9\��XDV�7�ដ�֞J�QlW+��c�	�膔��|��ycJ&��f����>S=Yt�C��,��y#��zc�ت�������N��#��q�H�I�-
E.�o��1��y)�◚Y0��F�~���s��V�HVB��`�6�T�&}(f�3��.b
�>o~�9V�Jnx;�T��I��t;���M+.� �ӗӿ�^RR��G����������Y�s�p>�}���sV|]�n�����6ۮ���#���P�f�&���Z��]���{;�R��kű��g)�ǳ��X�@�Jh峫��⚞}Iq&�vvhn�`�Gw�YxU��/e��i<�>Q�V=�e�$����?o]}X������H^o*��y�3k��-��{�ݏ����ģ�lE�(��S�Iޘ7'���{~u�T�9��:w�S1��L����!��?�T�ϭȉ<x�z���vΫ�W�g��Ly�3R7�L�&Y��dP�q��im�̅O7VXܓ���ԫ���'�v�n�u��9y*u4$4�n���f�܃�c��4��5{=��-�!��������~��������y���?Y�>z�_a�, ��\:{�>R#e'9.��9X��վ�J!��'=K;wcLP�&�s3y{��u�~*�|��a�!ˍt�v�[nl^���T/�a�N��9�'�k�������cU.z��ݐ��!"�srz(桘�y���~���8=CZ��2�{�X�w<�X&P�������(9����2d���ԉ�+X���m�r�����nK���[W�;rA<W�w�G�O���sfm�S��kv��)�ܬ��=Ay)��f.8�P�C��;3#��P�����U�\}���+q3&vК���S��#(�y*�F�Y�ؤ��:7kS�/�H���?���BǴs�+.�Eɯ����N��N�v�;��/�Ֆ�J{��
�6�l'SD�x�^�� �j�\~�ܞWIex�]�-}٬d��!�+�,ܷB�h=�Q�[�{P^6��pq	y�|��6��z�ݡn�7�J�/t�A�w{�l��vhF1�JH� 󉅎����	&��,Sv��b�E]��O{yʾݹ�*)2�8����\ԭ<D�o'����1���<�{��&aض�#�ĵ�u���V��-P;Ss{g��>���#O*3���lD��);*����l4��}���X�X4�����{�8ûXJ?�y��z��G� ����]kXsO�M	}�qCY�U�e94S��~�[��w��{��F���}kX�a�y�|^>�suۅX{V�k}�-F��rA��s&��J���G���2��S�S�#��S؝8�{��,j^����,0X�9_����zٕ�+�^ix��+]��b���e�o���*X�@�fZ������C\��3����+�����m�70kʱ�\��� ��}��*��ӭ�h�|��XVĨ���6�˛��=9-�]�/-L!�zZy�dꦆ�@�V:r�-�į�Y��r)J&b'[��vv�>;�C�����/�,C���0w�oP�J�)�:*{7d�������'�s�
��<��5�޽��$ո����W�,�镳��SA8��/GOaBo�6�k��N�vu�[
Q3Qn*����x����z!��Q�|�����,c
SIڎǘ������Ė&�1����$�c�w7��_����b��Ry�篻=�e-7��Ds]1�/5R���{���1��%��HH;ν!dַ^R�A���.���ծ�c[Y����v�S��V��o��V:AkR����X�-���n�'y�X/5�/2����sn�U����S�EZ��N��x��q���}6�r�4���t���2U8�W!��"���#<\�c�b^ޭ��=����3A�$4��>������ȳ"e����9�j��g�7Z�wG[��Gx(
�fS|��Y���v^mm5�^Tu��݄�f#3r]�6.�-��=���f7}�4a�Ϋ<��<BZ�Yޘ�3ZVG�ET���l��̗x!����	��(�ol7a�v�^t9u-�$�����l����X�a��ѝ�:��,8N�s�ͤ���k�omn ���75`���u�*��q��fhSi�"*�ӗo(�A�k�1u�A`8\ݺD�v��R`���x�{��pdt����c��պ0_X�N*sZ���\
)ӗ��d�ƌ�Z7\��)��v
�Ch�XVU�m�Jې�`��Ya'e�rҨ�^��'��GQ����;`�N�>;�T��m[�.!�G��Z��7���i��U�$ujǟ#���kr�R�h,�xkO�n�������h`�ᓋ�WCDi��u��{W��B `Z([�b�hݳԒ�킶�{���#�=\��FH�:��d��
��I�|x߭������8c#T��B�v�@�WK[�w����5��g[H�zJdE[�	���T�/ ���f�Ae�57����� 
+��y8F��Uj̐�=�b�a�8��������'���@tgX�����G)�v�bT��8���4��:v�,R_Hdw��,R.�|)��iB�g4;��ځY�ns�ef�4j�Wj����:��ˏN�|5�y��x�"�5��]@�I�j!��<���9���{K@e+�E]����2���j ���z�T���V�{i!Y 鏃+tj9o�m|^`l��N�]Z��B�l�X˫`s�ҙ�׫_-*v�A�V�O�IαN����aU*t�b�M�Ƴ:BQu��tO:��j9�Ś,��
W{mނ�/��.��i<��U	M�f_P� ac]_J��X��ݕ�c�{4����[���T�ԩ�m�0���6mq��-ma�h���0(�d������X�Ra��
�s��ջ�a-`?^ ��fj��$�:�b��� Y����/b����*��-�!��jc�V����1ҫPK��cw���+3;�]��P���;֬��>Ž�hp�#�h_^��R#�z:,T)�p�fg�����H{^E�>Q�S��D���n� �s
U�;m�z����f-|��z�1҉{;���J�P
��2��!�z�o	��E+Y� �pG���]q�mB�[[�-6c]������MTkv�#$����r�Wm|�h*�6Q�b��[�l���Z�*��a�e�Ɛ`�O�j�(�˘T|��͙t�m�=�vT��8�=�����BksV�Q���z8w1��)5֚�5R����Y6��v��$/u)}o4)��ŝ��{¤kq��$�XdV�1X�3�޴��c��܊�n�f2�쟯�~�zߋ�����F�B,@U�
���*�Jʂ���TdQAV�F"��"
���
 %�*�Y
�6��F����V!ka�+(ZЭb2JԅJ�BV(6�,�X��T`�h(����ZфP�!m�T��KmlEQ�RV�i(�ԍ�P�hJ�Y�*��X҄QImQ`TP+�QVv�AE�kH�X�XT"�T�)XTX0a
B)b"!*B�UB,�H�d�X�Z��U��mZ�R"²X,��d�+P
��iѴ+�*Q����PP�Q*B��$+"$Omo���#V�w/-c,�!4g8�Yu�l�w��bt�����z{h)|�P�� }j�,�\�F�1���Ѳ���;��gDF(w��hny�7�=_}�X�w:���דbYF:�+c5���Vܶ ��X�G��^��J���2�����
]z��Ŝ��P��e)�HO�Y�:������*�P���$��	m��rvr󵾹�Sld�A�����G�����`��5c>��7��;�#��!������:�#j#�2�'[�:��cU���z�	��a�<	~��b{N��U7�V|J�ϝ�L�jy��ޫz�4OB3�k#m걓ۭ�I�b��kê���)��7�	��-ͦ�9\�ulIDO(r�7dE���yV����m�n�A�ïN_S�OK�z�@E/l��K��	��w�ێ��,� �(�_*	A�z*�������%�v8¼�D���6��Ey��c���lh�����!��2�`8an��ˍ����Sr��f����:�����.#b��k��HR���b�4m��8�<O�`�4s�Y^]��Sή������Z1+ƶ�����ݜ��j�r��x�S���J*�]�F��N���4zF�ǣ��
Q�ZZs�R������� �{�4��C�M�/���k����	\��R���|c��+�'����4�Bi_�w�`/2��8�{NʰVi�7Y;7M��T���:ʖ1�ܽu����З5e�.�vӘ�h�P�we��;N�[i[9a�{��Fuk�]}��{��NO_������/pb%���@k�e��Q1�q^�}@�Р%m7�0�a��S!��.�Y�»1u��SR�512�*,�*%�L�j�k�t{��X0v��Xt��ٟS<+�r
�w��{w���k����ur�n�]��
(�ՓMH��Y��6_E����(�2��q� �}qN^�yܺTUu"��@d7�{a`�ɏ�/�������_�疈{��>�^6����U�L��/^�����ӷS�b���� ��LO(�:��"��X��F�~5n:��6"R%	���p��;Kqfl�Ĩ.;!�P�:!��UU�yS��򡔪a��$,�XF��m�a�H�<�����/�F@lݬ��w�d2�R��x�����,��%��|@����+�!N|��S��I�������[�0��jS>�{7r�8�թ�w�p���(WR�/��iA�r�MGݩh-)���{�����t�ődt�zB�3;K�"&]�7oҨ���aL�,��8rFZ�io%�S�wd?m�.�+��Dta�m���V4Wiek���i�3�+�ߏ�<�n�|�u�,�˳�����K��|�e߱�nܫ�6�����w)F"A� H�g-9�"��dck0�ȓ
3��I��-�{\�q�*8[�i���]�ɫ��3J9���3�c.�`Y�l�2��Jp��)G�T���$�����ڥ	B��/9M?C��Ɩr�r �b	L�;f�F=Ϧϑپw��t�,D^�;�:hv�����$�ƻ���N2�ȇ6�� �K�H!i�v|c�I��Y�����<�%MB4U�}�X�<~`?5;A���yB�S�x}*���zS�2��{��P���.��+�ڞ���S���-���lܨ���d&�4]2i�6h7T!M�)ZP>��.ׁ�o�FOu��w2�'c
b�"���x������A��h4����.5^p�����]Uo�����ٷl�-\�v9�(J�xq���b�3W����4��˩a�7��з�9�S{P���XK�<�Y�ʋH9ٚ��z@�Nl�
F�%�
Dڭ��7Չ�O�wK�N�o��������q��/���
�	��v*<��&U�jp֚��`qN5*^�����T��v�Y���s���X.����O��"\������TE>�}N7�k��-��-�bߕ���<�,Vt�;�X�q���R�]/)����4�M΀X�fiQN���Ezad3G�E�G烇sn�|g�s�򖖭�օ����Y��8��2oT�pd|������d"{T'��˩8��>ק3UD���g�U{V�y{�.���ۨ��`���I)ˌ�"ɮs�S��-b��yC���'y�8�
�#Jz��s]�z�&3�-�up���ۧYn���~�݇�9��P#Aj(dK�Ҥ�O��`'a��5½8�7�r�(f�=_\�s�:'�7w�Y0zt��rʺ�#�L�������t\q�>FSJ���s�9�������7����~�r!�*"�i2c� �	F�Ϲ�u�A�	��>v�_���cN���Wn�(��x{,��A>�ȿc*XpAJ�G	�'c�H!�k�B�i�NQ�lĺ���Kg33!W���ݡ[z}�Y>�耮�����<����w����;���1p�
��D;f���7��.����{%��׬A�����[˘4g\�R�n���]}%�D�=k��M���t�Z�\����NK��8��g�'�Z9��s�(�^�Z�GBs�p��2�JAa}��5}@��S�v��2E���F��(^�;��p᠝��n���$�AO�SQ��J�4Ef�۹שVTf�u)�߶I���|�9���C^.�8
`Q��V8�Se�>k1��&�Z�ǻ��A���c�^��]�C�r�|Ю�T���P���P�V��H��99C-���O��[�/2���
�#@�vO�T��̔v��ޔ���)��L�d��1-MEK�Ժ�v��/q�<�M�= ��ّ�H)�dX!�a�Q/&2��Y�z{T�[�6'-'�u��yM&��̺5�t���1�<WPf�κyef��R+X�G%���<ˡ�/b�]3�Z�>����3M�{�8:�>X){0��X'��>.����]&E�1n!ǐ5�h4�h36��:��{6QY&F����� �Ts����v���i�3�lT����h�@�<#y�8�M��������z]���{�6�jpg	 cd0Yk{���Q���ŤĳX�%���+���@j/U@�6���e`���0r�t�0:�F���ڄe��B�h���x������e�=i%��">zuX(��z�"�Wb:v[�W�U��f�5�*�J��0�w{��}���>���|���+�>:7Ԥ�Փ�"�+�qP嚴鸺�P�{�+"�/'u�Q���<�qE�,�q3ĕCU{`HWI-�)���q�J��j}]��_ofZ�n-�7��UМ�G	�a5H�T�El#�yB��@D�a�&1ǟ>-��sBjzW'�f��"�����9%P���M �]����=�ܨ�����2$.m�Ӻ0�ˎ���7Xqd?TIhJN���r��	�;�j��R���nI$+�4���U3�\N8���܂ ���{��	]����	�Q��J����ؘ}TB��w}$���u���,�&;��� �`��Ezaq~���F�*��e�esn�S�$�bw�g\N�W=�|m�uެ��MY�Ӣڑ�&a���ݱ]���{��ʵ�%'G;�%��f�����������.�a�����1�D���p*V��8�D+Y��e��-s��Di�٪�(��i�%�}���`t���1eu�:pМ������X���[KU��X�R�� �ܤJ�I�.!$�އ�"��P���}/�wz؝����R�Q������+��4������ꓤ�j�+�szQ�����A�K�9Ѭ�� e����Zi(�:v\ e�:k@�9�}�ʉ�ʗts5�1�	F� ����H�p���W���Z�HB�3A5 �-*���u�P{H��y�x�6�Ϲ���s{L���,����{ad}1�E�?>?l�ƹ�4�0U8�8�p�g�~�z��W��6���ճ��'0���텝S\�a�s��!����r�$�f.廋���f�4�6Ū��*6kb�Iq��&|1P�:!�]�Y~ȣMy�gw�^��S�ݟ���(T�j��N����G��V�a�f�+9����ܷ�њ����!�# w,���y莌<m��'�\�}�.���
L>�;�u:��̈�{�ky�󘨠F?\��C���`gI(�rNU���S�|B�9G�@.U��g*�΂K澮���@�'��1��8\I�_O�g��p6�:Ez�u��8U�c��Q����ǜy��Wh � `"'���"�*g��Jp���s9Pg�0k�E>t'��7��Z��f��Yw���ڴ���N�HA)'lJ��g���;��e�k#� 3�٬�ެ��6� �]\�Un�a�����eVM+FQ�)��xMf\ד(�Z�2�c�=�s}�n���@n�GXSn��:"#(Hf���V 	>t��G�	��sZ�-}��4P��J���$;EX7���`]�,�Л�ɝ��G�ʕ���=�@{(�5�0L�$�x�8�q���X¸=����ڌ���pc3�0���<0,�	ݳ����S�F"� �:\���lV���҉;��>l���E{�ܯ #�	���^s��n�2,B��R��}�Pd��m�G�bfx�����1\iԆr�]"��c�����h�Tq�25^p��V`Q�5�Ó�]������gf�':ra\2��$a��8B����0.��Q	��Ag6���ҕyx���Gvf�>6�qm6,�ۓ|p��1
����"�O+�)���{�����!̞���q�/�񠷝@x��5��{]v]#�|*R� ���#�ܱ����&r�X�~}��}	�jl���TPѱd���U��N��)��d���5/e���D�~��Q�T�8s3�\��#o�ޜ�ZuQY<�@��[9�k����]U��u��f�P�ײ�'��q9�:��{뢩�3�{K�hk���Q��b�%C&!ћ�.�*�+��6���y��n�m��NVt�wY�'��l�͛������smZ���Dm=V1��T4t-��dg#p�ŉΩ�>;����W�3�Y�eZ2�Db�zv��]��}�A+����qgru���Mwj�ؼ�KV�����dT�ފ!��VD���U��-�v�0�|��:/�*��.�xHy��t�Z�]R�K��N�:8��#�L��"H��;��E�V�/��������FOr�~�|���*�M��N��Đ�' @���1���}Ogʆ����م,l��ܙ�oo���J�Ş<F���eC�pAJ�G	�3�<��@F,��2v1Cw�9�u]�l�#/� �F':u�fM�LmB6�C�-�2���{r���y�]ƭN�E��v���$�(�w���8h'n���Yl�D��x��S�u=ݼ�5iD�i� ��`��5b��6�IȾؠ��1A9}����L
8��[�f��{�8���dU뛜z�͈�����c�Q�.|״��[7�I��I�R�EE��*bi�w"�Z�J��Q���q�	�s�<�����	�_>�*�p�Y�`듼3����7Uⵛ�3P)����nz�Jh$��s�@'����daxݙ�3�|&�I�͐r�99�����d0��o<BN)9�im�p�K�룖hv;Ɋ�bS �n�PZ���n�\{o�.�����]i"�]�R�;�<3.�>&uY��͵H	eY)����(Px�pS�v����v�8�L��q�����[]&EzTsgj\��U�%�;5�~�ޯ�o�k�-ܣX:\F��v�(J��=�5
 E��;�L!�R��m'���A���,r�g����駋s�������]Ux�y%��Fr�)�bܺ�i��L.��0b������6�K:��|�_���ݦ͉P�+��wB�+T���pw�k��MU{K�=AP���p�$�((���i���z#k{��ܝX2�YVX�灮���'�B�ۏ4�Vz8�r�D��9W��w6_ume�n�]�9e*��}���g�*����"�ZKt�mxw_ѡYwa���>yǯ{wR&�
���yFg���ST���V�t�#�
"���>��ʮ"��<��&��n�A��G"�2��K�1�*����My��g�ՙ/��[��It�4�Lk�9-d`,��*$�5���J��8�wG��v([T �/b�Xoh�1��F\"�D�.[�I$[�**�js��WE]\E�t�g���d9̋N݉�s�?6�4�"����������i��:�Q�(��A�F��Vwxd)��b�u�n�Tl?�������S�(a}�����h���J��A5�j����'H_e^>�@�]�Z;]�-�&�Ծ���)���49uib	�n�ns1��⡦�ʰΰ2��ck--��������q��v����B��XB;Y��'@��op c�j�ϸ�Aҧo`w�EP��N9��z�����!�����nrøދ����(2���$�Dǝy���͍����me�4)̣��3\�,q� ��
�I�'3	��8V�N�n_P��c������\N�	ڵ�֛�0c�hd=�d�]B�lj�6+��q8������|a|��J"v�f� �+v=�LЅ[�:f���\)N��K���� '9�rYYA�a&@�(w"�Tdzd.�"9Ou�S�:\���C!6x0�WN�֐)�I�2�)AM�ǚ��vst���V�z����
����Pۉ\�΂����rgh�	�y���lCdB��� Es8�u��:��+��DU���6���o�::����e^m��h7�7B��Nŵ���5mW�5X��?J%�/
��	��,�r�=��&̘��[�Kcy&%\���;��e�X�Cm�]U�f
�4桓�nL���{na8�h>�Q)�W`�2��&e��N��7�����o��♰!�L�/ u���Wviр��!�R�a�6�9�έDrv���oL�Iq�f<��k�y�h���4�)�wVJ�yҵXjۦ�w���yV�r��Ei%�Y>┮<�V�aZ��u��iރ�pAԽ�^6���îK�r�:���t\��OW,�+����[	ʸ���o���9�;K*&�;��H#��r��	�#�]���.cZ����4��u;�R+�yg������/���c��P�i(�D�WW�1��׸3,�<�b鍉zX�l�պI�ʏxmf 6􇯾�ok�4\kp�3�ʖ���qrM�e��wb��1m*K���o�6�e�̠.��mw���F���S$��Xf�񮗙W����g#MR�퀡�X�WG/ol\Æ�t]o����1��I�Uw���Ǒv�om�Y���K傔�6B��u�l㬾�� &�P-�Ы���+3�4n] Y��ȥ��&���r��%	�]�k{����̟]�ȋ*�V�Ŵ7l��Z����CFGm_L;K����.Ј��<� t�*ֵ9�Y� �nr_"��8T7r2mn6��ֻ�5�^pT1,���Τ�Q�t4���V�Uv�l͸�b$��=�:���rĭD)��s�,|wy�Ff��qvvͭևoE���*Ӹ���6�a�4�N��r�]E��>���eӹI��z�����fV#�̻n<�9޺Yl�<wߞ? ��P�+AeBX(�%�X"� �V�Q�+l
*,("����,*TPb�
T���)iRa%Ar�ks�+��Aih)��ڈ��EE���ejUdu�"��\*��*����`�M`��*��`�QB�aZ�6��Æq�`X���&L��**ŕ�#l�����QAB��TYZ�-�-�����T�AE+�c�&@��ۙ\�`VJȫ�eTUH�jZ�R���-�V�Q(²�B�U��*�jJR�Kh"�5����C0�r����DօV��"fE
�]n��%Im�m�U+F���U"�����e�T+Z����V��UPPD�J��̣�TB""H�Aj��o.�t%èlOu	%Wh�Ч2o2�!�(r`f�X�Yѕ����8�H !��9�`b[��w����S\�c�рI"Ȼ���#.�g:�)Y�D9��!�VF�*�Q�\�e;�]�=�v��qR�[~M���~�2�Mk��
z"
Zf���|t+�ӫ5���b����NM�h̪Zڈ�bMڕ�@��a����[nb�I@��
��0ߦ�4 ���r���Q�lK��D�u��8v	�A:d�T �u���q��4Wi�8_q���K,��na�[���҃wx��6�ȯ���yݑak�][�E���i�s"��1���*�ݭ;'5���WqU�yH�
�da��.�(.��>�'?>?l�Ɯi�|^�p�S�[o3��Z��ג62hDz�rp�9G��o*�U��+��k�^Y����捜`<e����Q>�0̤���6M����\ҁᏐ�ً�Wδ}0z��~n�P(l�1�o���;U�m�s�TY��n��}c#��8tVfv/$(�q�t��=JW ��=��X����;��#���ܲ�Ҿ/":0�m�I��#ǈ]�����F˞[f�v�	Se���9�Ze�Hv�a!0���7i锑�J�����O���3W׬�Y����b�����f��s��҂^�o�D7{�t��R>bS3g��MU�u�3s���S�Z��t�cD�o$Ӄ�1�Tݭ=gf�	jG�9(PRp�ў��].;�﫰��y�K.�:ߜ��*:�x�r#�#j��bnS�q\��c�̀�TJ�TK����Ÿ��K����QV��&T�G\f_]��V���q.�yޤ'L[D��Ă8�4�LG':-*�q��`�3��I�xl�R�`�q�w�/��ٓ){�~�M���Pb	J�I�R�f=Ϧ�|���/%�z�~���@aӻ�����Y�k�����,��{v�b�*,( �	:8���@!rB�W9{�X`!sW�im�b�'�����D7�ˠ��>.)��B�Nb��b��x�s�-��6l3�Z��+��S�������`+��	��9d�0l�uA�p���0Ԉ� ���z�JM���/��L��F�e�dVk�	%UP,�,',�҉��4�A�B���d�X� B����˥��`יtٳӧ6�d3��gN����g�K�Y��u��kgg-�Lvu��ND�#���W�Х�a�Jr#v8���#��>�R�����9����h2��\z�Ө$�e��.�vS;J�N�+[#�}��<}LC��wWa��stz!������ǩ>�q>2SCR�cf>�E�:RʹAdt��Ő?Yk%9�N�qFuX�Ƚ%N>�w�5��z�r���ѳ:-E�q��[QBRĳ^w�ʿ{i�����_�vn��>(�|�8{��D�kZYk(�{UCM�r9��E�|�;�2q@&����T��/�U�ܗ��6�R���}xK��]o��q����7~��ea`>\6�`̊�]�^̸�2�Ӊ�~Xn�N0ˉ:vH@������O+��)�dnk��\��]Sظ�������{���GK=`���]��D��*A���v�ԢPwxNL���s��[�2x�5�~엗�V�Y�犘�8��iM� ��v�w��q�I�A����LqQ<Z�Z����.��l��3�Bp��H�' @���1���s<`���S,j�\��*Ɯ���\y�tv*�^o�2,cP��W2�iP5�qo���k_=�p���Ȅ�a�VWQ�}�s���~7yb5=��:�d�ڄm9�8d�؀r7�%觷Q	7k"���^�o(ٍ��$=��bI:J���3���y;w��1� ޫ�y]�9��JS�A:ɼ�^%��.g�s� ��-�C�u oqL�;"��0uq�܄�L��<Ģ��u1�[��ՌWy�:Y��Iι��[�/p��h�d��:�u��u*�q�N�;F����;0�MU��:��]xm�!�8�uw��4F\�P�^wnuc�r^$_���^ӓ�ᠯ�0�>�hCYU˘,і��Kem�Ȇ'k���k�F���K�VZ�9�HV�n�A�.�,����*���kw]����2�L&��.b��3GM�+�}
�fJ;~޻қ�n�N,�]ܤ��آ�g�b�����s�@'�@Y���'�8̉*ᛝ�a��@Yyr���0��E\i�T�Ή@<�)MX'CKw(�t���G���1�8Scjjiw<�T
�`������r�#}V�*�u������}<t��0�J��1u��9����Ͼ:�SQV����/�����EW��(�	܍ະ�E��k�^㛷��J0f�x�9�uY������ݵ^qY��do;�������s�>��)�$��~K½~Y�q�9��5�:a���� +]���mt��C�6�^���=!Ѷ�j�'dɳ]צ3��D8���>�fHF";�=U,��Z�x\r=�j�f���a�;tY!�d9ٛ{�G�.��6����@��d�/{��SUh�tnB�uV�=��V욲j� ��	�i$Ge�h��:ɳqw@��gc�%Է�.h�����i
]L�!�����F��C�\w^���+~[�a,�	��\zp��,�-B��`h7�+��hn��'k'Y�,L�9��udH�t�9�r^ȼrJ�}d�o����N�+��w\D�j賅Mn�ڂ� ����t]D���S�U*xS�7t'`�P�4إ	�cOD��nrY�/LBy$�����Nz�������X�%p��=s#��z��qc��ƩF_^	~���wÊ򩂕�$�s�0���`�чL�u���N���<e	Ur�ﻹ��P�,�FM��W2ۚ�< ��)X3FvfO�\���F��6��N��)r��2y䍨�C��À5��~njtП{�y�
�@�4�]��0�7G�YU�Lo)0�w�Px�;�X�']E����h'L�j�k�tE���T������d��]�<�7m^Z�!������"�7W!X�셮It�S���^�F%IdƷ\�Gt�"{s׺�vp+�`�0���m����*ōq����#�N~|o��֎W2nۛ,\��a;�z��h��EwB��X򷭫Z��N�+!/�'�:�1!�-`��R��1֔I�g`q�.�jpZ����w�g#8gv��Jx
��:�ۛ��S%��L��ٓ7W=5nm	Ftksj^��1��3f��.�{8�k'`t�5ᑅ#���'%V*��Wj+x���!�6ȷ��e�0�9�oz����f�uq�m�U��i@���x���Jnx�:�n�xnВ���U6�L���wǎӦ6=Dp�
���u��9 ѳ��=�O�^�%�>=���.	�R9��.�+��#��ԝ�O���8!2�*�m�Ժ0�c��X��B��<k���c:Ie��A�P��1�v�U��s���{�j�"��A�fx�>�&�0�(Wd_O��.��@��[��q3�C��U�����iu�#0E�Oʉ*	�&L zM�ۮ{M	9X�Θ�:�m�����;�2�����~k���ѱ �rv �A)P$���Pk�=ϤwE�/��V��E������e�"�3�����/n�
pT�D����LYɭu1������s��ȁ��&�=�T�#������;�||_�a�O��(��T ��IoVMv�>~��XfY��4|��\9�1c(��9�p.��y���jQ5x�!��K�7&t[���1ecs�cyyqVLFB��Jl99a|~������q��,Ϻgd���D;F����١��U���aS��a�FΧ�%;a���s��VT�~�N�gWLwa��n��Y<�-̆F�
m��Ҷ�**�OE������-��Xh��]Ef���%wQg8�I�$��`���[��H�}uͽ��aA��(�kȾ���|�Z=��|�Ѿ���AM����U��ݱ\	P81-p'�&�f���`<�jʇ���-�����O������*����Mg1���9NVJ�ҹ�CT�
��i�X��Ct,�ǉ�B�{XWe��|*R��\��{݉+��]��q�DʺGK󪡦��C�9��E�|󎑹�&�H'$���@B#nP�_J����y-�Ր�F8�C!�}/����p�gع7�F������u��CNd�*8B��`��w�tq�Qu��qP��UB��@����\K�Ҟ�F�5��3=��fsq;Mck'i�������àKE4k�~��,�GiR���v��k�tf�"�'{�Z�ǐS��;�y˴��i�2�������^�_�7�~Ol�8l]����f�Дb��Տ������X��y[��$e�W��ȏ�B�o=}��:{ZͪQfP������6L�'$�+n��v���K��Νd]}P�WC�r�ۣ�q���i�d��uv��jP�ь��5�u��+*F�ϑM*�H��NDt]q�H_� wI���Q?o�>6�!2S����[5�|�\oF	s�V�B�M�E�P�����z$p�
��<K��~�<���b�ue;�J�R����59Ӽ1ݳ&�#�N}(8 �!�L`O#7zg��c��� �1n�X�rv�`�9��x��y;w���gfX�J!r�<���=퇓��S�I	���D���X*WF߶I���|�9��r�!狡�;�'T��ԫ�T�_S���U���
��`�* �zD)�0�0�ܕ�`o>ۨ����n�iƯû��{t�ga�@��Pˎ�M5X\���C4�2&d��Kȱ�(�.��)�l�o��RG�u+�6ϔ�y9`���M+��t��1Wd
�}�7j��4k��Ӛ�V����͎/�#�P�p͍�w�<��"i�yM�h4�r�`�q�ݷѽ��fی��׭��
r�!\FW��q[�A�D��|����I��-�/Z�e|�?vv���zKu(��F�;	�z��u`W�&���׏#HΉW��D�^���]B��=���Wq��,�; ����m��伧�k��y; ]M�Ѡj.ﮒP7�rXڶ;fa)�j��y��8-���ܢ2|d�:F\�6ar�Y�꼇r�#D܍50�GX� b������(���~;��d�,.d���Sٜ8{qf%SM�e�mx\	`�My��N@}P8 ��w�L@y�����S<ۼO_Nd",���:�M�F��^��\6N�k�`�=)��>@V��}��n:�BT��r�Cg��w�'\�!š��7��"9�m�"_�2zC�B93=�xu̗�Q`�I[��ל��X�u$O��N}x����Q!5H�
iGH�8���$h-�&��UJ�S��P�x9�Hf�gO,VA�,�����/����'C}v�k�	<&���rwg��^���(�T�q~��0Ж�TrV8�)���9�D��t����`�d�E�&v��m��M�J��js�.I]�x���(�rn����jW�OW��2ޮ��!z���=m���6UZ����P��J��|`�*l4����ƃ߇�{��iDFrÃ "8�C�q~N�_��� ����L�J��3��2h�$�^��k�W{�#Kω{�Ҧ��jV������v���6K��^Q��+<�*fr�>�[Y�s��KgX<��D��譼A�V=IB���9��i#'
 kMf�^�٩��I�wS�;�ǀ.�Er'3�7��w�LZ��;��A�O(kjK����q�)��l�s���hrT� Hk��ߛ���Z�s\P�tC�H�.�^9����֑�e�c���;(g[!���B,��i�%�}�ק,��3�sR�N\�4�g���r[����T��p��9�b����ȣur��vB�$�r$񖚲y9"�(Ք�����Bk&�z��X/�b�5�yL�
�da���3+h.��>�y9���g�*��Gg��Iɝ5p�r�GJ�U�h
���tj���Z<NJͪ��B�G�y[��BB�)��ڻ��3Ӫ�#��V8�v�Q�^9!�]E�/�
��ni.�Z�%d�g>��D�]�DR��r0*�mΙQg�|�[��x��f���ueLP߃�����˩�k7R�7DB�q?eQU��.	�R9��r˷J�������}r{.A"&�>��tΣq�-x�q0�N�wQ;�%���@vVo:Ie��A�
��yOe�,��js��\GK���B�Q3�p%P\*��\�ew���7U
�Ÿ�K����Q�����<�����f��ٷn�ĳ��Y�D��\�p�Φ��9�n��;$ǵ�|��a�΂�V8^].�ǸU�x�-ڣr����ڍ6�]���t����ulm�ڠ��rI�t�j�mN�*��g���vH��4jۑ��C��2.\�x��e��ו�y��Cd�j����&�3d�;�U����D���W��00�6�ᵦ�Ln���7ǊT]�צ��#ȋ��(!:��zly�y����,�1�x��o�nd�b�,�Sa���.�MJ���S(�t�}���n!�QcK��r��4a�(��t���7%NM�j�]kF��!i�{Oa������H�Z.��Z���|TT73%�+��+Dñc#�B�(�]�iշ�F0n�'���C���Z�U �{��u�}&�1��oa��[e�l�Y@ܥ��^	r�A�� �;U�ˮ�&b+Z���}�M̮����oT�Sx��'�w�u�s�b���*J�Μk1�L˗]Qm`iS�`�w��!����R�����*K�pR�O]n�mn��E,�Iql,�e���M^e)�J��{A�S���s"Gw�K
��G��`\vԙ�|�WxI2��;���ko�dF[���x�n7��n�(��md���/�7�9�����<���q��:�0Zur��-��ʶ�d���$\&f�׼ݾ�g�ps����B�)h�e�AI)�Z��v.�f�GW�N��z��d=o�=x���94�QW�-�XT�O�M���-�gʈ�Q�xJ�''�έb�te<#�ϰHW*2��
��aa��$�4l�nh�㾥���)e�(�n�	'r����C���2��s��>|��T,�(gP�N���F�inGm���;z��Y�r~D��o�'�eyޑ�9ڈ����r������,��7�e��"

�׿v$�.�;�e��F��p��j���^K�"�Yu�I{�5m�q��Wqt/��E�֖��0��:!SDJ-�cAVT�`كb���]c]�'͋M��yb��ʻ��J��Zܦ��ۼ1�6$��&n�� �vsbw�倦�hun[O���n�KEk��X3N��S�*��q�*�NM(7*]m��V��yWkf�$J2����{�]J�������߀9&n�
F��ٺ���8[�J@./�Ɩ[��%j]e�vk
�̦_P�wdݓzw3�ɢ��i㝮����zN�٫(\�u����Q���ܤ�T�uLU�iTan��ib�f���L+�#ro;�uoP,��j�W���FeZ��ںTr�,VirՋd�E�.�c]�\�'n=��a�x�_.��+DW�sZ j���U�_I�RG����d���
K���Q؍t�
���3��p�����+MH\�#]q����p�D��R�B�]Ĝ�6 ��9�1;{z����
~j�����Ql
Զ����Z�`���p�V
d*�B�sr]J fR��
6��+Yt�1X���[3�al�P��Z��*�[suH慶TYX�"��R
.eJ�����E(*��Q�QFD�[C kAkZ�K%�j,Pme-�Ub*��E"�a\�l��AJ�E�V�,��Df�m�PF�TsF�R�B�Q+-b5s+:т�aP��e̓�u�6ҫ*-�݌:�Z9�mbۭȂ�$�� ��Ҭ֦�Pm��ԬiV���XV�mVe�Q��ڢa�@��VT���)��뵶�0�:�mZ�EZ�V՚�EE2Q�\!�ء�X#�ئa�vK\&�D�f���UV�f}��U���9$��֢���L77"BdᎮR��v��<@��FF�pr��7���WK+k&΃v,w��1�j�8�'s��Y�W@��u����W�x�$4�UL�s���c3�;4��B��o0q��AJ���$�\�N�۵ܝ�"�b	H�;`�Phǹ��"Tj�NeK�<�r{Uز�bw��pD^�;�N���,��/n��*,( �	:8����y-���nck��js�E,@�*j�n�C�ˠ��>�snT%�o�LBSZg|�d��;ʢk����`�S�6��u��V#�	��L�s���}�9[a��(U�l�U�Y�.������^ׁϚ�wp�y����3��!�yx┥��=�թ���w��GR������|�w�y���4%�i��d3`nH�Yӄ+���r޸��f#U�s�����̓u()*&�uN@���l�x�ypT[��n��6.WQ�Y�gY!�3����[��S6�iE\>�e�aE�8���-��Qo�6�//>}�6�vwVk��PYj���UP���/bJYՆ��{�'-H'@F;�Q����uoMF��9�GMʹ�wNV�"(#�0�so�����=:��Ѻ��<o#��t�*Q����YB+�Ttӵp�Q���"�[�ۑYA���7�uˤ�@�44>�3�т�W7�ɵX�SG.�`�FE��U���ɚaXL� �۝�m�ԑ�H詞�GlA���8t�N��&���緥�L���fv�$��{x�!�"%��4"8�x��0�{yC���8�>�u��EF�#$�D6�K�6��c��K"/�I>[���弖��(L�@������d������u\2	xu��|��h����0m^�y�]n�1 ��\�SG!�*��͑賈~���˽����X�wQP��y��&H�Bԛ����w�L�}��J-ܛGI�2���wjI���$ߦ�e��7y�Ӭk��qǈ��Pd^1���uxD��n�V<^��V����!N������� �]~�Ƨ#:ڶdؘڄl'>��J�7kkZؕ\�q��� �H�T�HH[C:�U�NҌ�9΄sŜ8k�۱�s�r��66aj�w=����I����A;>.t��l=��!���r��{���m�i�a�8���s;u�t;a��uLۍ�8\�'�i���-e\[�>��4)+�������S����I%�_(ǆ�&�(s8�=P��[y�5�IAO��+��K�mR_�n[�P,�1�����Fd��Tch�zK��X���J��.aJ�����)g7�i��:6�Tr��qsH�}}��1���Ȭ�iN��ݩ䒈�Z$��n ߓ�6��,�j�����MzanO�T���X~w�1'��/9.)���Ԝ�(�{>S��i�@�]s�� ��vB�2�|�P6�@jj�Sw��R���P�4�f�$U�����\�+�+�h&�^ieɛ�q
1���Ư��c
^�ӥʴ:�Lq���ˎ�J҇�/���]M<����z��[����9�؀��i�y`���������G�_X]1!
$��37(���������5�ʲ��̙:0�A�eΞ�h�5U�.��7�	gk��s�8����v�%�S��ښ!�y���n�A䬅f�q�Z#ah��B�kg,�r�=ι[x�w|�cl��y�3a:n-ӤE�G�7,�51�'d-�fM;'�;�[�o�0��{W�g�~���+jH����F!)�d2�jQ}�
���b�V�ǉ$��<u���Ozfv�V�3(;���"���/U2�8/$[�y����_Fo����ӳ""�y�EnLX�#'����(���f7)�3k'%k9W�����/�7���u�"Bb��!y���\�F9�����IL�yK!�ySy �ěb��1�N��P.���e ���cPQ�n����
��U��U\�2W<rQ�4��v�M�d�Q���U�T��2�B��n�T���n3v�ʋ3H1��s��q�� �n+c�dC�9$�� �)P4c\l�=��9�~��()I�PgA����-$;�~�-'8<+Eo�B�\
)A)W�� �{"��:��F�"�w5L�g&/���[w،�6�Y�\�!���'R/|��8*"
[㵋%����w�<�3��L��*�R�=^��&���C���Z�v�����,B�*�N!���=+�s	F�b{�ĥ�d<��d#~IU�"���MP��zn�\���9B3�3�<���f��f�@��(/�q̋�D:�
�tԅ���]��yo�y&C�ź:�z��m���iW��:6�?�o?���
�����f]b>��`9�b�[�>���חٸÙ3ƺ4��ق�l�$�{���q&��Um\��#�nz�6��㳧F1�5�X.\�Nh�c�Fd{|��*�xV��s�Q'�X�	,�Y�[{V��xt`�&W�׷q��m�u�1�V=���g�ⷘ/t�c��
��,��nv�籜�Ւ�R�3
��,t*��&l�A����_��h\�
]k3çxứ7��Uu�γ�⇳��M}�ܵ���u��R�q�H�1J(�#��3��u=��F*�j3Ũ��wǎy�鍋"���0m��5p���籝NL��d���PRu��#���ܲ�:�ؿ<6�{�cm���N��/tv���� ���*&FИ��b��^ɒ���Vt��NCh9W�bn�&]�<wl�B����;-^�t�C���x�>������wM��=�#Ʀ���=�։�Y��teP9fs���p�H��N��T*<L���CJD�s��XK�	�Ow4֫Y����u�Pg�3��#���S{v���SJU6A��׎|����4q;}�z6��Qߕ�����t�$ӄs��4�dD=�#<*+��r"<�QO��z��o��q� -���J_Gy��ˤ�x}��TzS �i�|�yW��Y3�mɈT�2	�:��C�2u}{0��d&�0�&�gk#2���2%{%��dꂼmO%+JK8�kq�!���A��.w]�X(�9()��)�
�(���q<�=Q��[M�ʽ۸�B݇*V��,�A&�ֹ��me3�^U�8��Rw���ç{_@)��r*ժ8�^��s��dɹl\N����fvk����h�2X�<�gv�5�_
��ىE���f0�vA����Ww�}�\��=������1@�+�	���|^����]�u ����-o|���݁��.�2�TK�3�cd-�_Y��6-�㈾<5�}�W�~�av\�wUd1�C��L�{4��} �"�(������.�&[��:�J�M��iM��!�ɳyC��qG������S��=W��fNXR	��is5��;���}��V�p�
�V�n��N���Ⱦ��:�:���M瑿>{z*(
�a>�ypRK�����E��Y:�F�f���:�30�{~�ěι�R�kz\��{imgM��N���Ϲ�z޺ٍ�\��":QW�3�T�}3q.7H6��r/�h���j��$�Uϰ�1�a���|����jĔB0bA�E�1qɀґ�-��&e���W�Jw{|sT��G���V�V'�ßi�H `�MzɋU_v�nC�_iK���P�w�������	��q�r\/\q�)��ȱ�eA���ܳ��y���A���p�]����U�cx<�:���T*��c��nñ�2���/@+�K��W�]K���Aq׾-�s�'o�3Qq
q8�ٮ[ŝ8<��Υ�9`�u	G��F`ON�zx:�<c2!@,�Q�#��eYI�g�S4��#�J���W��̈r�.�#5��!Z�\<���m�^j8�	����.03~���u���QD��"auE��PG'iFs��8b&�nq��skku�}6���x� �?�|;�$�
S[��d���_lPV9Pg��A�HR���S��|�o2�#���U@�M�c��8\�'��h�:⮧Ns�(�Jg�=}��iN2�n��+�m̷̞��ډ\@�_M�0�2tџL-����}��3��^����'h���u'xeg�b��4���� ��vBӰ�	������O��|"���Yoc�P�p3[�=�ΉO+�SV	֖\�Ǘ3*�&f���\J��خ`ݚ~��D]��+ۗC��I{�R�<���[T�����N�\�ٮEs��K�-�ٌ�&���\i�G8��y��,��ӨX(u*�N�'ۮ�K6�%����a;��Ý�hW�[U.��T��+!����Wz�,[�\p��.`�j���]i7���v��=�|�"���/a</:P��!\�@'U<9ً�]�l���MX��xѦv������r"9ɕ�)ŵ6��jZ��b���U{dK��b&��4Ȓ�"�EzTs_7$mA}�(�w��1T��Q�_�w�y+"r0�����U�̿{���qV9*BS*P�$c>���Vz8�ͧM×(��9�~�"LtDH;!j���W�GSf�e�4���X������Ձ�$M���׈Jq�2�jQ|*Ҏ{`ac�rQc��*�.�\tUK�m�q��dBt:�Q!2�<��z�S,��%�yw՞x	.j��$+���u�E�	؇c���č�E�tX�����X�j������܍=��k���"�^-7�����a�VsȾ�����{v!�rI!L�)�k��ROlg9�-�^a;�_q���Ғ���R�=�"ӷba�QY&R�R�$�s�U�-{O�߫(Aϟ4�[az�U�۳��l��q���t2�sX�`���
f
W�!<�z��΋�u����Xd��W6B<���&�@�y)q�	k���sZA����m��r�S���ԅL�/�2�T�TG8�D+��d"������N�-H��rD&U�}Vt��8r���E��ѸQ�"���e�:����ܧ�-;kS�'�8�7��U;�6��wx��4#PƩ7d�`��8%R*��5�[�������$�8ϋ�I�7w�P�����G_lǅ�z�s�R�f�����1�+��p��{z�^,+��d�B�b�� �8ja�ȿT"xd�q@����yݑk]�"��#��ˬ��i>�=��-�4�%O�>]mXk|�1b����eHQCWb낪���V�cM\_�9�����j�5a�-͘*��q�@Dn�;�؇k�f)�� �N��>$����u�G�
s��戠*�<k0�����axV�7�݈�dcv��3�-��W��;e�8�q=�/��UT����M�9�Ӧ6,�#�&(�n�n��;�]:�w1�2Y��.d�PKې�΢���)܌�w,�*��}]�a��a1^�Ȼ�N.�"۞�m]��]�Α^�>ghV�Hx=��N�˰��{f����3=������}k�4X�d�����Z*����L�q�.$���h�0t�DAױ����yYVr���.�<*�/�1��P��AEx���3�%��<�oj��2�׵]*h�[s��tk�D��	��Q��؂(1�Q#dJ��fB��C��=#s�݉3qt8��f��]����[|0!���s�'�|�PΡ*q����:ޓ��yy��u��5dn+�}m3J���c6��{�(����,$���P^��,����Z��էEd���t�&JFѷ��a� qzlBT�8"-�;���Bܲ"���"��Qj!PNA����-l�֤���&@'@[��SP�q��A;�}bہ.�uږ�v��,tq1�Ƕ8��(�!=�f�]��n����>���o���s��'ԧ)(�̍ �z���t�8�kq�9�U�n���λ1.;ɹ��P ������^�,8Hy�Ě�5(8����ux�ٍ�7�<᝸^�a�F�C�]˲�W�޻6�X*��(!5D��Ȱ|ƅGvJ�_^�a�l�����ׂ���cV�O'�ܪ�3��@���e�J��C��aF�ȟ>
]�lsj��㳁�O��ɞ��s�Cf��*�9n���
���P�O��z���$-���❱R��{�e }CUXt)��j�"�CQ���@�t�N0:����o<�x��ª�"s9�n_o�E�l!b�|x ��΢����Ww������?�?�?�����O�ҵUWA� ��YC��UE��Z9"
�'���"��^�Pز���7/�������˪��k""! *��:B��'������N!�Y/�?���*��ZQ$�1��m�Y[]�z}��
㞠�R��kt\J�P�tj�|���}�b/�9/�\d�,�l��PUE��W���N>���xET_0�������@�%�����zS����^թ�����p�NE��a֡C�r ����
|��@3���P��V�Z�6j�1_������)�[��w��w�!0�]ʡ`��"��QUE��2�v5������,���J���"d�H�W�
��Ja�k�qe�P7����.��|���.�q����Z�v�H�5t�525�w+��[�9}�P��禳�-:B4Qz��Bf�^����~O0�B�i��v�qZ@�_�}gPpzS�	���^{t^e��^���rDQv'L`L}\F@�z���B��I��ް�DU�:C� ����>B�|��9@��dx����K%u�Ŀ]QT[�͵�B3PjH|�G\�UUE�[Ql`@�CxX�22XZԔ�wK�2��U����bR��qk��|��eAUQP���ݨ�8"
��}�Z��ͯ=�p��?��v�{̍��kM�Qν�wQ�=�k��C�~��s�<=Fԯ�~�)���
��e�6(��#��N�AU��\�	�S��_����hb:.�X5�;0[\���S�B�0�Q��N�p�:�a���(����#
��KiwHYUE�n*��6�ܒ�S��"cx4���h�n�5R�mMۋ�ZX$��"�/Ղ���
��P���a��X����w�#��x]��Ǎ�xQq �
���H/jC�(��2�^�w$S�	�F�