BZh91AY&SY��� _�`qc���fߠ����b+_                   �                           UT�  
J
 � ��_\�u��f�5݊�m0�Ϡ  � @  � � P � @ �  �	�EP$


��P �  
 6�P*� R�Q
���*�D ���@(RT(J �J �PVO����  мPـIR�(+`�$Wwt�\�O�w���z 1������ܞ�^�=�y���;� y���׽�y�Q���   ��E  �T}�tP}�{ۨ{�ء^tl����(��k�R��h�ϳ�R�<s��x>������Ԩ�4<���S�;�٠k� �|�U�s�R ���EQT�u�(W��Q�W�� �������ܚ��;;�{��W�ϯ�G�(��_[�h)�y��}����T�����
��@Ya����gEp  ��<�R@pv����w��@s\�箩> :n�>g��0I��릏�����w�<����t�n�����}�<����/�����  ( ����R�="�QIaD�ɅU� n��dW{��`y����g���>h+�����`<�v��>���{� �><w�P���}��  *�}JR `>� ^�&�;��o S�;���g!��{��S͞ �K�J� ;��{ z]O�� � �@  0�}%% 9�@J���(*�X�_���������^`���� ����'�-�"��`����<s ;�JG�y d  ��G�։H ��� S��d�xٌ���y�� w`�x��
�lz��s�;���= < �4y�I% �=*�*�JRN�*��'�C;z�=zn� py��fh����C�O&{�iW�$y �0   ^|�����X���4>� � ���!���y�N ��x��{�9 =2 }�D� P�P  ��� 
�djR��SC� `	�M S�"RUS h      ��U*�SҞ�M4��&�  �Od��IJ�FF�M4���I��T�L �` �M0�  ޥ��J��z&�	���M�hz�=F����_�����'��I:�=�-�|�Y�V��g��$��"}��?{�$�D��"	��I��H� �?���K?�����������d����9m����DI�Y>�D�e�������������T�$�u1d��LSI�9$ŒuLY&,b��1cŒb��LT��)�b��LY&,b��S1c�b��LY&,b�1cŒb�,����8��$�1bb�,b�ŝS8�)�$Œb�,�1c1UcŒb�,�1LT�1LTŌX�1�1N�b���$�I�1d��b��)�����,b���b�����ŌS�1LT�8��*ucŌXŌTŉ��dY&*b�)��������*b�՘�ŌTŌXŌTŌX�1S���1c�$�1d��,�Ŏ+Œuc1LS1d����Y*�)�b�)�����,b��*qLTŌY&*b�1c��TŌTŌX�1c�LUY�������,b�,b�,b�eXŌXŌXŌX�LS1S1qb�b�*b�,b�,b�,b�,b�,bՓ1S1S�LT�LT�1LTū�,�ŌS1S1c1LSU�b�)�b�)�b�*��1LXŌT�1c1cI�Y�$��1Rb�Œb��LT��XŒuLX�1cI�rI�$�:�LY&*LX���d��)�b��,�:�IŒb�,�ŌT���b��I�1bb�ŉ�$�J�1LSI��LY�LS꘦,�&,b�1d�LY'TŌY&,�Ȧ,�1Rb��I��LY1R�b�Œb��,�1d�c�N)�$�1c&)��W8�,�1Rb�1S&)�����$ŌY&,b�1d��LTŒb�*b�,ud��LS1d����LS�☱�$꘱�b��,�1d��LX�1z��S�1LS1LY&)���,�b�SI��LSI��1dŒ�b�,�ŌY&*b���V1LX�1c1LX�b��,b�,b�,b�)����LXŎ�b�*b�)���c�ŌS1d��b�1S:�8����b���b�.,U�XŌS1LX�1X��LX�1d��1Rb��N�,qc1LT�LXŒbɋ$ŕX�LX�1c1c1c��)�XŌS1LX�8�,�:����*b����uf)�1c�1LT��b�,b�,�\X�N��b�*LY&)�b�cI�1LSŌY&,����8�,�b�VI���1L^���1LT�1LT�1cȲLTŒb�,��1d��*���)��,b��1c��b�1d��)�b�1c��I�b��LSŒb���LS�1Rb�1cI��J�,b�1LT��1bbά�8�*b��*b�1\V)�S�1c�1cudŎ,b��*b�1cŒb�,�&)�b�����b�,b�*uf,qc1c1c1c��ŌT�1dŌXŌYU�bՓŌY&,b��1c1LY1L\Y*�)����*LT�Ŋ��b�)�b�)�'Vb�1cI�&,b�����,�qc1LTŌT�1dŌT��*qc1LX�LXŌY:�T☲LS�1LSucI�&)���b�Y�b�)���,b��LY*☦,b���b�)�UŌS1LXŒb�,�J�WŌT�LS1LXȦ,�������,b���'�N�b�)������9��LS�LX�LSuX��LX�LX�LXŌX�Œ��&,b�,b�,b�,b�,�Y���V1LY&*LX�U�1c1LY1LS1j�)�b�)���b�,b��b�,uLY1LTŌTŒbάb�S&,LSŒ�b�)�$ŌS1c1j��)�$Œb�,�'X�N,b��)�$Œb��XŒud���Ŏ,�I��f,LX��1Rb�8�1db��LSI�b��J�SŒb�,�&,b�qd��)�$�1d��1cŒq��:�1d��LT��,U�1d��)�$Œb��,�c�1d��,�I�$�I����)�I���,�I�'b�ŒucI�b��1bb�1�#:�T���1LT��)��LXŒc�I1N)�$�1Rb�)��N�I�LY&,b��LSI�$�Œ��&,b�1d����I�b�Y�$�I�b�Œb���LT�T��,b��1LX��T��:�)�$ŌY&,����1LY&,b�Œb��qS&,��LY&)1S�b���1d��1LT��V*LRqf*LY'Tŉ�9Q�$��8�I'LPbȒbȒb��*I&,�!�	:��⤒b�1Hb�1I$ŒI1P��LR1BU�$�!�Hń����Ł�"1b$�Db�#!�T%Q�X�LT�LT��$1R�b�*b���1c�&,b�,b�)�������œ1S�b�,b�*b�*b�,b�,c�&,qdŌX�LT�LT�1LXŌY:�b�XŌXŌY1LY1LTŊ�T�1LY&*b�*b������f,�LS1c1d��LY&*qX�LX��)�b�����b��U�1cŌY&)��LS8�S꘲LS�1d��N1�꘦,�I�LT��*b�ŉ�I��Tb�:�☩1cI�b��,�*��1cI�$�1d��LT�J�b�ŌSI��1d��LSI�:���?KZ�fX� )ɨ_�Nx��۵U2Le�čm��5!�f�k;�V��P��2�D�bÐ�B^$hS'-|�#IL�����	�z%���A2����PASJ��eZ��%Ǫ�-�* sol�w���5����I�n�l׮,?t�w�.\$�+m���/m�s͵s���Xs�\�Q�8S՜�h��I�0���Co{~�ІT;v-�4t�ȹ�Qa�q�,�eD������˧�0�S�ޯ;w�n�fi��n��Ď�-2\!�q-�&���ὖh6�W��b��抉�5��V��G��W�%όS8��%�&���Tܯv����i�p�vqc[Ol:������ʔD��+���G]]4�;�<%��:�#u��q������:"�ov�L�ʨ�ew/}�p��oYS7DG��9�nw'���6FU�%<�W8���tx4f5�-ެ�D�{e�W�C;8�%U��ը%7uN�j�1:��лN��WN�e8;�{���[�7K�C}ҥ���J{���!�cj��2��p�nh��%P�Y-��ppf�Ν�kN�4Z���p�H��Uۑ�S�w�=�5���e��4�w.��k��ӏ_u�+�&wL���1�I��t��lug-�uI�'�'�rܡ��v]]3L{�zD�gɘ{�,^h�"�;4�9��a51@�:[F�נ9U_��^���&`�-�x^��;�v�6�"i��q1���.�c!���(�7vm���e�aq�8��@X2L���ʫ�_���0���Z"��#�0>�s��#}�,�Z���r���Szݗ�^�}�������osg�C1��Z���.Z���Pl9%CRsb,<f�\2�3���1��9�ӽ��{:�����)���ܻ��;ϑ(�%��S�b�ێ��u�5��.��f�5ְ�1j#	Z��0�2;ov���4���O+z@��,{P�V��n�;V�m��μ3�%M�N�7r�.�jva�D���S��U ��%��;���Fi+C��� ���/�E�\��wN�S�s������$�ږhT��4Uz,�yS_l�0�j������*5F�A��;�\ޔ\�w�������vۼL�V��5��_o�]�T��U[��X�~颳h.�:;kx�{8:i����C9w[y���.�JEݑ���pU�7yw���Y�8�)e�_gNe9�.�<l#��٩ ����i�=ʱ��\���'q/� ʓ���sw�bkثp�y��g-˶�r�ϳmB�>�74`Fl�*!]��kKt�=K�72=j,$��p��3��9�vB"�@���kt4M(ڧ!p���� ���
 �dZjv<2om#��Kr�Ā0%OB'��b`|���ӇWV�$�͖L�۸���#1�XTü�xShZ �G[�T��b�T�q[�>�2|����-�z=��]e3oΔ�qFTV�V>�m�؞<�q,;��ڋX.�U�P`�9�(��^]:8��Gj1��7"���t��z-r��cZ�a��
G�ly���(),?;6S�ū�o&�wu�ZԂ�n������6��'fvT(>Ѫ��>
���F`lݠ�Z���r�eֆ�1�}�޻�4�3L���%��5�wC�\Hf�)!�������,N3FnË��/��݊�gD3S�,�
H���40�I�8�t�ԝ��%�[�c���ZvQ�G�c՚%��8���)E�\�r��	�n���ey.��*�>=W
�C!gE�C�D�/.�7 �q��v�/ָ���%�Y`y�.mRoJ`�χ1��ݪ`�vn��� ����Nߓ��In�m������^��x�w	f�O{5����"s.-]�/�HBI_��)��N�{%�#��lAk\���h����Yӓ�׏l��5c�jZ�1(��/A��X͇�ߐz�ͻ���Z4�ᨃ��Z2Ğ��]�"�,�<$[j�b�V��u�.8��v��� .f��Ǜ�[%+�����J�
򨙊�罊*Rza��OW���5�����Q�f�V�Dׂ���.��5��ޢ��ɲr!�I���[ǹJv�c�����n����u�B�7	�Ã�n��՚��
ُ;�JW����<�n]�sVʺr��Qx��<"��c�s%�-k�d}F�����ND���т�n�x˛Ѽ*jn��2�i���o}�>G��6�JB+Qd���)p>�7�;T�֝�XgS]d
]��obV�K&Ց����76>90]l��� mp��˰�,t<9��Q�tV�|�7�ՓG�t�^%��f�L+�c�.E!�&h@kT��;_27��P֓�ݎ��^�c]zj��q���e��fv��2}>�K�x�v�>�t��i�ͮׄ���T��۽�`�:&otШ[��/l�&tS���b۔p�o�=@�Ď]��/�8܊�&Y���q�
��,��Si>C�A]��V��r�i�3�|Y�J��o����;����w^V�=�R��p�Y�1�t��Z@�#t� �%�ߘ��ev�ޭ%�ssV^�vI���:]�v�$K��H��F%�m-�q@�ᱍji��@��N�|lw�قw�ˡhCL����UT�7��>{7Gn�3:��C޺���k��,9�X�Eٝ�tpo`Yf��'.�9�����MTm8t��qnvFλȳ�2GgDV��cY�m�����,��7Wls���a��}������f��!���L�덋��EH�y��/zݠ��6�����7y�]O*գ��oN���]�u��*z��W�{p�m��5�x�������(���S�O>l�P-{bn��n�;�c�3b��oJ!�yٿ ���zP�9��%����ø�b���f�2lz���;]
.x[�lZ�!��v��D�
�: m�����GK�.}ؖ	���Y�N�m/�;�3 ����r�ɐд�5�ht���UOWF/[�7f߸���f�4�7�[�O�3#r�n6\���3z�onw�+~E����ib��է,-Kػ:�6n�`L���Mݢ!��ƹ�1b8:�=�	���bS!��Bv�8t=����h.��%��3C�"���%[�hns� =M��o��2��dp��8�g +K5o^P٠ry�,*�B^:Va��������k�5��w>Z���E
�[�]����5$�Z�`̮�w�3trN��Y�uS 穑�q֤�M#�x�J47��N�u�ܵ�/[�H&Zu>�`����,X��w:�-�`�	�s������ w2 �>���O��eʹqzEH�Dش���N� �N��sͬb�}t�@^��!z�Q/F�L@
�)NAHirn4�T-W�w"1TV��I�݇����C�ͭ��Ð��̔c0哔-��e����r�j�ۛ�┞SCȻk1���� ս��MT��v�p>�m��vG3��e��Z�Dd`�^F
�@�u�]�tB;��s;�MUw#m�Ĝ�87�S�Q���"�<y�CVi�&42W�wJV�����&�Xڻ�JbȚ�\�a�r-}�l�r#Q�=t�۶�Mi���d$���t��bU�&ί�q�؎p#sU �=���|�>|��q���|�_!��F߻r�U�xT�w�i��UJݐ|-{�`�Q��4�k�OI��:$.�b��y	&��߻y�
�{�u��>Y�(�0���<����Y�}ݖ��`[�k��Ir�d,`��$\���/`=n��o��o'�@9`/g��_Ht��+�״�G`(!Ӿ�{�d��SB]�����A�u�=zBUN�J\,g��LҬ<*�t�&U2�w���W/h�I4wڽ�:h��,8��0�;b�8��'5 �y:�t�h˹�m�\����MC��j��k(�\7f+D[�K���;#p�sם����������[�괕�A*{@�h��湚��t}�r�eXú�ㇰ5A�{YɀtT��ij�24n� �.�=��%1h*p�����h-�Op3�M�Õ�����s"ͳp�z��g��S��-Ouk�6ٝ�	%�ڄ�wT8H�j�sn�2,�lɗf���-!gV8懭f��J����)�c�q-ɻ��h���|u�鴈c|8f����5�v��VoLh��v�Rj[t��Nٺ!Ű�wOx`Q�d�����ږ��I20�˼VCܫxs �Cኑ;����N�w}�76���xf(�ܖŷBX��'��qLZ���zD!��n�ȠŽ�1�hA�ۇ��F?�v1�2,��Ƅ�hkAڑV���Z�έ��ZcYz������x�Y��Oz2.׫Gђ�`��ԛ�T\U�
�'9۷nu�w�&śR�t��N[f��(/k�=��'Ӝy�X��٭n9��՜�on�J:1��cSo!'���=���lWt�.]r|�waY���N����{\�[qܵ�%�&t�����D ?���}5gs�r>9ں؂x�($�EhT�KomO_�4��wQz�ُ��ИNu�9�h�����vJ���Z�����Hq�ה�.�N١1��BѷK`�@�p�1�@�
��
�Q�+;���56�ӓ��=��q�q��:H�߁F�vt&��N
r��nA��c�� h�b�Q<��e��Ob�*mtƕ���H��	��V�v�v�운RTp@���]�1S�N�7���{���[�
˼S��N��	 �R�}�&n���D��.;d撗n��{�q+S�Ń5�tM�,�V똖�cn�t<Hn!�#�O_*��æSeӶҶn>�/�ov��?��N����H��ݞ|%�)n����2�o`�6m��ϙʀ1G"Kdm�~�q������q�k�YĽ�7k��&l�:�!���^~�x�>�vBo��2�jNݤ=wo귢D�̉��-Ե��<�{��ۇWq�ƞ4���C��L@��O��Jn],f >�n��r]��H�8�)h_N�i=�=�����8dY�[y��z��Z���5e<ӱ����=���U�)������p��z�OL���{���>;��ɻ�S��콻�Kb<�J5�w��k���P!�� �½KgV��dQ�7Y'Z!L=��t�����wG8ςW0�`�c��Q����?A�B���3!����Y�)&V��>7�1SS.*��T����yZ6��s/�NrK��9��;U!�.��#�N�<��Ǧ��_!u��ыT�|��R����+��
��D�p�?���f0!C&$�6��]��Ệ���w:o��)䯶#Gb�9#�ƹ{��eS+��'��yF<���S��0��܆��}�&J*����*s���6"�������/>t���ݤu>�ݯԾ��������V905�� ���7�u"
�K|��Ƀ8{�;W�o����Xp�ዷ]���V��Y�x���d/7&�踨��PXFڐ��r,��*������ٺ!�M���iS}=�R�)���+�7��کJ���t�5�l��ꚼ�����?�]���<�{��|{�����������wϽj����{zP;Q_ӷ��Yϕ����~J8���=����y�	�`�X&@�J»�����0����^f!E�5��L�-�!<��o��Dj�X�5y�{��Ź���#9M0q#C$<���_�V��O�N��'�W�2rkě7�ыӄCqJ nOR���6��~m����7�r��/iv���͖���"\\�3)�;,u��Q��f�1*�A�x~v�g��6�淞��;��"�H&C8�'�R�����I�B\��}�z�ъ�u^��26�Wp���e)qN���.W㨳�_F!S��*ʸ�2��d�G��	��'�XP�~I%IWX�o�:��R���+�1mw��J/�a�q!Z���`r͖6�8����o�3��8�[��a��1����k�����=^a~�ݎ�b��+��#W��T�gxh�45��p���;Q�����#��Q��A�q2��&o���T��N�t���qO�[��cf��_����ԑ�����"�)sw�Hk<��Il��Dߖ�R¯;��ô$|�E�Wj�ո�v#s|[�[��Խ�&�j3��K�a�g���盘�iU_'�`��9���~5�ɐH�Dz�+�Um�UI!4V�U�.:L�!#0���Xl��i�=�����gYĤ��>��ßd lm���Y̓Woil�d�X4�$��C��Fob��=0TWo,��s�d��]�ȋ�Ӿ�|��F��TP#E�X����'���:q��a�	�Y?���%n(�s��fzi�˚��σl)���.��n���!`�"H^�-�n��p2=-C�}�=��*�t���Ս�8���!�sQ����<���๼��a�Oky�J��/gv�6�|���M��B�k���w-�d��r#ĪnZ��]��0�<� `�����R��[,VI��xy��]m2ߗ��U�K�Qi�s��Q��!�N]���ZŊ�Q��L{#g���9W��,����<wӒU�O埅�<t��Y������.�]�0g�w�b`̚���r����6L'wpB�ᝓP�x�7]0Uò��)���gW�H��e?G��j��JR��ow-�R �6y�ܫu��i��q��}�y`�t�ѥ=z���y|d���6z~�㹷 Y�����Ej�b-�,Č-TY@�6Na
�=�S��x&k�Q������_��>�?��=��vn��	'�dE�-I"�Il�B�!lA%�Z��$KR!jD�%�D�D�ȑ-�D[[Z�[$��Ԅ��Z����Ii$�����$��-�"Z�Z	$��jH�Kd��ih�%�-�Z����-	l�����KD[%� KR-���- ��Z��D�[$����h���I[$%��Z�-B%��B%���-DI-BKa$�$Ij$��	i�-�!l�H�hIi�?I뙗��;?O^�����n�����y神�����k���÷J�,�׻�A�Vo���V�щqǔ<~���6�|�fb������v9�����K(Y15�8R�k��]��䷅�/aFٝnX�fV<<�r������@�5n g��UQ��.�g|5�9KK��OT�q"�@��re�����np�*��qǃ��Lr��;m:U�o$�� �ah�龃���fB"�N��� �f5-���}�|��Pe�����,@�A8C	���t����h�7[���𝓣�� ���sr�hSk)�C�|�͇��l�]hca7$q �X�
���yc�k%��f1)��;ݭ�k��K{���gq�F�'߆������m�^ۛzBi�����I�X�/"�r&[H�p��Pn����s���v�=t,S)X�zb�}���i7	"�[����wkQ��X<l��Q��kt�GZA�&�$�ab y�˃��x�0>�%��>'� �M6�͠��g T�K��|��8��@t�M!fLk/�0�̷[& P\'G�?{~<���+��q���!	�ZҖ=����s��lЬ]M��47kyC�
�h0��mgio`oCF/��?k�vϰ�s�\c�ކ�BIq����NT�%�!�zGټ-��Xۭ�D0��\\T���`� �Y�
=��7(�s �P�<%��HM�aċ%��cX���1 �H�|Qj�>b���?���i㱏	���j�jX����n5��B����mi��9�|ᮏ�Q���3u���,&�\��M,׶��Q��D"1��^�L������a���8߮�Ξ��!�/n��y��Ǒ�t<��F��D�!��`�#��||����j��j�|���d�c쭚��'�G�ۨn�	�����9�
K�c��z�Ϊޤ�s'���`0&�L�|�����4,@=�`��A�u=%�u��ͺ�����vw-l�
������*V6\b�Z��M�gz)��m�<��<�3Ლ��F�RxQ��MS�@S�63VL	�P2��@��L�s~��Q�a�0`Ή���1��A4�-a���=CY-se61Ĳ�!���v��݌kB:W��6�'�B�Y{���D�		�~s�߷D!?=�e��?��'����蟀�"'������3������?��}v����v�bz�s�ڠƵn��tj�����vC�a��=��b��_v���ix�+"�oP�ۘ��ݍ�-Z	<Er�-�k��#��H��7�eT0|�J��3}�]�W�vy��"qh�ʹTm��3+�4y{K�Bq�/f����zy���#O5�.���sC.B��M]SG���y�u�X`~�a��0?�9��Kk�a�qS<�S�p�����;���;E_+�!��^0]�ɇW�������Y:�{�����7%���� ��v.����f>Jpյ�#�^����S>�w�G���':Qa�!���̬��_�,g��]�Lx|1��k�VqZ�R�<��jos޻���[��3`�[��e�=�!2W�眂�V|V4�t���W���]ݹgq��ӫ8�K��~)�@��XQ�|3�Lb�/al��!��w���E�؝ G�@��#iȯ�k!l؄K����uҳ����tn�+}g]b�5FP6.�	�����-�d��3���M���
�>���Ig��O'�T��"n�����;���>5������kcZֵ�kZ֫Zֵ�k�Z�kZֵ���kZֵ�kZ�ֵ�k�Z�ֵ�k�cZֵ�{kZ�Zֵֺ�k�Zֵ�kZצ��u�kZ׶��5�kZ�ƵZֵ�k_[ֵֺ�k�cZֵ�{kZ�Zֵ�MkZƵ�kֵ�MkZ�Zֵ�mj��kZ־�5�kZֵ��ֵ�k^�ֵֺ���kZ��ֵ�kZ�֫Z�5�k_^��Zֵ�MkZƵ�5�c���j��kZ־��k�kZֽ��kXֵ�zkU�kZֵ�����l�m���t���O���s���;���2��(��rj,tO/����8p����N瞷�os��99�J��/dͺ�,��C�0{��W�G͊������*v��;:r7�{��_U��6k��`�,if���X�o�m#���^[ק�_\�~��̾�в�i� �xn��Y�)e9���Eo���\V^R*{6�%�>P��5&db��Oٙ��Q� -82�ia��e�>�Tj�[{��Oz��.�3�类�bX�O�L��}�_b�"n焷1�3��yҫ3�{��ϯ����m����Z0j�;.�}�/#F�_��||�N��t�FS[����7�M"��cڼ������s��M�Q��������ޝwʿ+b�ۛ{�~��9�gw��9�HӨ�{�F�x'�ta��`�P�/[z�P����.�N6w_8��&C��!��V8��`ᆤ��];뀬��M�/�$��s�N�T[�.�v�3vk��>*"/�&��GL��� ]�����;���m�ĸʳW�˳��a���F��cW���x��+32-8�tj���y�jջ���W�����=%��j��϶Н>��ΊFDH�ٚ�z��v1��9	��Cc;z|}}k^�ֵָ�k_ֵֵ�k^�ֵֵ�k^�ֵֵ�k^�ֵ�zkZ�5�kXֵ�zkU�kZֵ�V��k^�ֵ�kZֵ��k�kZֵ�k�kZ�5�k^�ֵֵ�k^�ֵָ�k_�kZֵ�kU�kZֵ�q�zkZ�=��u�kZצ��cZֵֺ�k�Z�kZֵ���kZֵ�}j��kZ�ֵ�kZ�Zֵ�|lkZֵ�k[ֵ�k_�ֽ��zzc�{kZֱ�kZ�ֵ�k^�ֵֺ�k^�ֵֺ���kZ������/;���w��q$�N0�̯�g{e���J�Ϫ�kHCK�b׳����ޏr������I����C#F�E9P��V��ꚯ�tϳ3��9�ۻ)�\1w��E~>���F*֎���43�y�� �mg��bYfwUp�;K��o��~ϸfeC��k�쮃5x�ϝ�u`X��~�V����}�Í����a���|�znN�	�e}��i��}:EF/T�S�\�
Z����ކP0W���� ���4�%�
��v��<����s}���2�����}�;���;�,ۍGm
tB�O3H�l�G��s����2͞q)Ҽ��?b�'{8�����z�9^����c]���|�[a=QI��E�z3}�]�x�zg��������ۦ��Go	�k~��eJ,�#�{��39�_}�|���rk/v�����}=-F������k� �{a��C�S����y��:�û�����߾�y��C�muɪ\�f��%sM�}��nyɤv��x�Mu����@).ki���hG=\�]�������,b �h����K��S���<�����>�����>��cZֵ�{kZ�Zֵ�MkZƵ�k^�ֵ�kZֽ5�kֵ�kZ��kZֵ�mk]kZ�Zֵ�|lkZֵ�k�U�kZֵ�lkZֵ�k�U�kZֽ��u�kZצ��cZֵ�kZצ��u�kZ׶Ƶ�kZֵ��kZֵ��V��kZ�ƵƵ�lk�Zֱ�k]kZֵ�k�kZֵ�kZֽ��u�kZƵ�k�Z�ֵ�k�Z�ֵ�k�cZֵ�c���]kZֵ�|k\kZֵ�k[ֵ�kZ��kZֵ�mk�3������-�ǪG�zVz7�`��M�l�{ȭȺ�U�tp(ܡ��<}�a���Ӓ'��X3�b�{�^�]L."�M����;�P*��[x��y����oOnͳ�G>��RY��hK�Y���ʂ,�ؽ�<��cJ�}ph�l�`�{��4Ny'����v�\L��'<��_�}�/�
`�f�7��h���=���3e�N.e߾ϴ�$����)^�^�Oq��M:v�e+VÛ�9�{��֩�9�2Y�ãƾF=����²��V}�k�=��u�)��N|�=C�ܼ��}K������3NHN{�v{|qy��y{��3U�s����v���<��-+ʗ����5G&���mF�Q�.n��r��]�\���F�ެ���]��1���g��ȍ�|�.y�䲮B�i·�8$>� ܰ���o����"��+6U��@(���2U�a�Y3&F��D�0I��~μw�{��||1M����C��$ӷ��V��T�����A����J�*�8 9���rXW~������ֵ��ֵ�kZ�֫Zֵ�k_Z�kZֵ�}j��kZֵ��ֵ�kZֶ5�kZ־5�5�kXֵ�zkU�kZֵ��V��kZ�ֵZֵ�k_[ֵ�kZ�Ƶ�kZ־�Zֵ�k�Z�Zֵ�kZֽ5�q�kZ־5�q�kZ־5�ֵ�kZ��ֵ�k^�ֵֺ�k�Zֱ�kZƵ�k�Z�kXֵ�zj��kZ׶����kZ�ֵ�kZ�Zֵ�{lkZֱ�cZ�kZֵ�kcZֵ�kZ֫Zֵ�k�cZֵ�k_\��=�ɟ>�����8��������{�D�1��S��s�v���'vo��rļC:�z_F�|��O\�)�s�x�cSM���&��[�F�s�_.�6	�16>c��[�pNW��L�>�(=�sS�z��b�^���H'<�ت��-�Ĺ�l�ֈ	��?qUW��Sݥf�x�ܻ�k"�l�0��g{� }�Ux���~9�	b9�����'�虲����4|H�
p�3i�=�wY+5�8pw[�I>����X�;���,Ӟ�|N�K�Ƀ�;thWVM�&�f�s�,>����iŖ�ێ��'����]��گ�>�Ґ������,eg����s�� �Ўk��	�3K2jYAS��Vx������V��}���S�ជ4.���u�;׳b����A}M�1���2
�����F�6�]8���K�m��͘��Y����y>I�q�v�#ճ��$�Lޒ!�����,Ͻ�{�{h�	���tnv��U~I��t��&�>�LFG�3&����=��u���P�m������O�Ǉ8���+�=��QN��f���]���}$ <��h��=]$�fn}�������@�uZ׃��.�ۑe;���DY͈Q����K>j�@`����f�~?2��F��|�*颎����K�Y��"1���V ��Ӻ�=33=OI��9�Ν��8�ʗ�����_\��]�d���;�31�X��?{�e�k��ଖ���mVc����}�! c��3���E���DE�����|�w���[�BN�q3(8u(�y0E�)��%�30��iP6��H�n �̱�X�,�C�P����Q� 1����@�S�O�6���N���Y��G��ýVfafHzc�P��r�.VF{^%�{��raXO�IZF�C%$�E��J��%����7V�N{Ď���S�ƐE�����RV�፝�	6�L� j�3�]��9�e2?�>�~-�&s��E�*�W����[{r��<�|�E�B�xu�-��H.��I<��z�g����u`	��ώ�@��ص�ј���1BJK���(u���g�1˂�⯦@^o�&-ħa섎���$@[15L$��-Ij4��9�v�8W�n�+my7����0P!L �;32w;��}yFU95�.=s��!�y/��q��^���}�4���<<ޝJ��*��ˊ�`����f��Ǚ�϶ǚ����-�)e+���cs��m�}�E�:��f8Ģ��c�K�M���z�evv�zI������Q�"�^�@���qn�BRREV�]n���@F�[���5��"6lK�s��@G�X�dy��~�����������7�M	��������zT0t�s>�Nq�1����j3<8ѯ۞Rn>}5뽾���}�[��#���_-���Z:�3{�����E�=��ˍP\1nnf}�)�zoٙF��\�[��wgD�[��)��;�0��;$�M�Vk��ϝ�0İ��}������<�-y�T*`I|���ѡ��D��áL臁8�h۹7/�+/lu"����^���O��>�QC��yzo0��x;����C���(o�sxޞ��sC4�bnh\<��ݥ�ÈCf,s�@j�lU���Ͼ�2�gQRG���~�Pg�(mMa�g�4h.�f1���S_��QbA�%�{)^/��4��3{�y7��˝_gٽ�s�_o{W�>�o��*�W�I�X|MiN�ϰ���N"���V�
}�8q �ISXL�VHqN��7��{F��6s�x>�So���� Qݪ�����G#tDM`�- ����8G�.k��𼵞�7�:>�?f\�8-Ը(�f�}��{���yhL������/f&��-��V��ncg�ŋ�,J����ri��ssyD���k~��Ǣ�Hϳ/�PyQ�B�{�b��М�g,�ƖvS��c�X�&f>��l=y���������ƑD�7�x���\�۳3&���眎܋�A�a��F!}��G��7���}�C'Ц{��fO��~�+�&w��
�x�bev��jyh��>�����
 ��ӾVӫ0#�*�WǷKs>�-=h���jw5Hz���=�ԃ��f���G��;3wY�1Q��u��\�(�bI�u98�G���#ݴU ��3���&}�N��/?�)8����vj[�v�7Cї�����$���ۍi^̗�a�����,��-z0����`p��ň���%���t��r�_R�����O��n.ط�?I�v���c����a
\��s��]�5���{\}�w�
ש�b)��ݖb?|c�+�z�O����Z�wz��΂����q�Tg�2���-�n+��S��z`�/�v� ��ʧ;'M˙��{s��V�ct$�{L~^vdn+�c0�|��G����'�O�^~���v��H�y �Ώ�Nn?����������|�j>�.��骭Fy�G����?�;t|�'ӏ�!ŗv��x�z7�uﾙn�cx��������V���J>�����]�#]}�|.LG&D����~�=�j��۾�{���g��*����/ڎgk�"���9���w×�/�yl�qPh���]�rxc'�W�<e 2z������9����fk����G^Pɚ�Z�*�ly{�vγ-��������	��7s_�p�4�v8;�5���x��4���VZ�X���%ޗ����c>g�o��Q=�t�ϼ����:�7��╩8�&7`��Nnɉ��ݍ��ac����9�p;��9��u2z�b��VE�pS��qݫ��>�^��3��F��Wm�Wo��;A�^��;<!��fd��}�H1��DOػPX�_n���a��N���vy��fCO����)�ݽ���ڛّ��/�s�ák�7퇚ӝt�6Soomˢ{������w�X�����]4b�����zU��P1��{9ӝ<�ݚyyo��Q�=�x�{��b��ud�ұ�^�z�r�������������t�Mή��݃=|������@�.xH엳s_ox,�~������^5�[��F)v2���[� �n�SC���,�r������4��;7`�
n�`��Xڻ�O�;�s;ݻ�P��I�*�r�w���]�{����8�w�M�b[驞o�+k���tz���wa0νsGN�����t^�B�dxT���L�  � ԃХ��(��	�.Q/7�lJ��ROPx��I<�ߥ�M���W��v���g�RGx����<�X��r�9��q��ˏ��^����W��<��G�{}�.5}�k�����74.�)���;'�Օ�s�ƿ�:F�y.���ܖ�<���f�� �G���!ԟ;TO�1ӽ�3>��0�R����x���"��JL���?wvJ{&���3s�~�"�ĀG����nk�AAi��籫���}�;�
��rp؋~�{�@`^�IY-ɉ%n�b��>��������W���$��['����������� o���?W�w�U������!uT�	�@�HT�h�+N6q�,� W�F�!��ڬ�<��Xvy����<ۖ�`����2\�#��6ɩ  O�c
 X��ĖyZ	��f (9e�׈�}>���xY@0BX���E���6�-�t�iK\�܋�Ym��5j���n��L[��U!C���;C��/�ݱ׸��Pf�q8�v:^��'�ԏ^��On�qٷ.��^XB�EX�`�m���d;W��9�ު�́�ɕ��e#tQ�/+���m,x���9�.��9�8�˷l؀�{���T�،V���Dl][3�񷓳p�İ�c�i�2#�Muf7�-��3C�y�Q�c��t�*�d��m]/�lG�-�-!.R�����P���p���.�d�j:�.��-�&���&�X�;X�-��&t޸�:�W�W]b�p���Βc��C�n��<�M�{K]��4GN�y�X8�B�2��7;ú�%���k��w';M�'��n�k����ݘ���3���qp[���w�����:���:�F�����E�*qϰR��ץ�{]vkvU5��$��LC7%B�K���ո�F��Ƚ�L�5n{n:����>�㧴Bs=y����4p��;\� <wk"�5�v��D;lO�-�	Щ�.�e1�f��lø�
�,��x׈=Pv�	����<[�Ɵ3t}�^��"�`��Ek�G.�d�=���s�� 6�^oe5�؎q��W�Bc�-��G��u��5ۘ��6t��X�]�7?=���h�v���t�k�q��W�x�]� o4%	4�����T�ƣ6�ٶ8K����kv܏R��]��+�pv�1��1NlK{y뵹:��Omt������5��jc�F+&�e'�pr�97��-'7�w����b-K�8Y��Qn�;6]�Z"�LD�P��ت�����e�5�zۢ����Eۮ��k�4�k���mČ<�f�y�M��x&3�.�lZճv�z�u�mhڅ�%��1ͱ�6�.6�N`�r�d��5�ڂݧ6����@��$ԕՉ�m;x#{pv�C�^[�!ۚ��=q�m�1K��ǰ�%�������n@����ޜrK8�p�.K6�N[,h3���D���,���H�B+A��)a��2B	[)-2�eB�嘣1ʌ�L^^Bn�^F�Ҝ���n����1M[xC@�v"�mq�&	-c��.=]k��`���d^�
<h'u{]w��.�f�m��D��f�$%���&��X���1�dwd���=k�&p���֫��p�GMHֶ	ICi@	Lkn��prS��u�.Ϯ�bM�e�e�w�30֑���1�ŭ��lM�&��M.��+&K.��<��X:�L�e��_��y����L�S�{.�7]F�N������nN�<;(\xu�a,:�����tBnqr��koE�	�lq��^��4*�9��5��z�'��+�8�獨�<jP�����㮱u�� j6%jʭЪ�.��..՝b�wZ3�a�ps�ި۱�m7�60�	��4,�!q�҃�X�B�f�A;�uYku�����rzC.��@eٮх�c�5:��!�b�3p�tq�ݍƎ�(չ�&���QϷ;�}'5��`u� ���w����Gi��i���+ۯKs��c�x���U&���c[mS���8�q�I�c���r
u�k��(�u�H�.ڎ��d��k����k�s
�Te�JL�&�cM�n)cKx�RjQ�+GW����ZV�c��@�]��[�qX������p�s�ыk��f���ͤ{מ+����66�8N޷$��NK;�-��\ḳ����6(6�w=uY��r@\��:�=��UkL�+��Wr9x$�O ��T�˸��k����9������W+0mkFvɼ�!<��q=�Ős	��(b�@�H�������`�W0���L�ƀ<ыWMSe�`ˤQ��ic���q�bN�5��n��=������$�ڳ�-���#�s۟cc�X��B�Gg;��ul�n+.k�RGo34rƸ�<b��f��!)� Л�[K5�Pen�v�1�f
����e�v&�b�Z`a+���^@3�7�|eT���Vjb\��ƌZ)��\r�%�SY�Ty�U̇0��UͷiN1��KA�K]<��b�ܛZ�
y��W,�V�-�n-�YH�1�0׍�t�ڡ�+Cmf��0�8@\	w+G[i�M^wZ�՜]<�gS��b�q=��JbJts��\�p�Ҋ[�,��n��oZ�t�G7��ۭ�j퍹⛅��F�����;�0N��N�6�n�\͸n��._[���=�zwe�Iء�8�j�X�mէ�A���*e2^r���@���<��{n9��>���|l����i�:p��kA�Ll�]��q4����4U�ƫ����Fb1�Ҷ��\�[Br���<<��N3(�B�[c�5,���{�9�ɻ�l��ѹY�8�ۦ�"͡ck�0тG8�c���s�=�;�2<]�I�8wY(1���e!](836���eA�ŌJR���դ&3dor[��vq��g5 ݣ4 �WFl�����݁N4tv쏣��<�u`A��*A:�u.3雯8�qh����<�A�:Yq�N�7n�S-S�I�z������["��fhVR� \�0�[4�Lvv�N��l���x��7�:3�\��v�e��H��v\@���R;��6^ǂ�q�+=�y�|)۰qvA�MV�4��H����L]���L�K6��G�^g�@�qsz�܉ѱ��\n�X0��
2e��Zi��-�P��M4!JD�4	�L�Me�l�s0<38KHh��;[LB=�RYvn;XnV�����N9.�.�v�,���9��8�HV����eĆy��tpm��.�{)�X��q��8�s3in �4��C�7.c6#ۻ�
'r�J��
	�B���X��^��p�G:g���ĭwB��m����gRQ�4�/�: �&�G\h���n�rl!�{"�.T�*Q�/v�ۡ�l^g�<"p��.0�8��B�ڳc�u���fN���ݤ�E�M	���p����7�Γ�3��<֍�n.#�JDB�	,BЕ�@�t6w1�rqyVMg�%��uY6x.�vÎj�FA��4�C�-�]�b�`L@���T�r�<s�F�[=��FБ�=�r��q�;X�&�M�z'ڞ�zÂ����q�=��(�W����v�W��t��^��n�=	�gj��l]�����2;���dyu��P|mˏ[�.m�۬u'h� &�r�BS�+���_g��i�c��tve��.�.mIE=lv{�7Na̛�un[�z���yl+�kFhQ������ �f��A��I{fln�e�aivK�ּ���[�pv1y�m��0�0�q[r���K��,aBA�j'mIϋ��K> �Yӣ�V�S��Ϙ�vqv."�spl.^�;gX:`��@cs�����sp�3���	E��x�ѹ���uʶ���z;U��31�]�:���ֻnz�[��魚������j�����������ꪪ��j����������������#O�c����n����U�N�+P2��+B�F�2�a��1�����:_k���eG��fe�g$�Q,G�\�X���#�*G��#�dC�pfՆ��1ti	��u�_��]w�OZ�t���6%μͺ�����M�c2^�uf�;�{�ѻ����;�$�"�*��ta�:wk��@p��n��;�Vqx�ׄC�&r�ע�h�dh"B���8�#;��`O瀬k_���E��"��/fԺ�ͅX��]��^�l�>y�
n��n]m7�n�Tc�ܪ��X��)�j����Qe�mYZ!l��D�B���nY�f�����ƵZֵ�k_[ֵ�������5)�6���)hV	ƫ�)�%7s*��h��Y9\�'-��1��}k�Z�kZֵ���kZ�1�c�����iEU�FcOU�#_r�n�J�Պ�iS�F���뎸Ƶ���|kU�kZֵ���kZ�1�{z��e�Ys��\����̠�R���D�G�;��9,坩��<|q�1�}k��ƵZֵ�k_[ֵ�c����&�b��e�ut�I[����=	.jɬC%�`�\��(XbS�	���-�.�q)�eL{��R�e�!�����HTGH����`,��Y�����3BHc-TBE�Z�G-c[�2�@���,$R�X`�K
VZ�־!%ıTY��	-h�I&�SPP%�[d����Ҁ�ZT�DP%L|ˤP�j�BM2H�ƒ�	�f0q�2�BŐ�Y�����V��aD���ᘦB
�JHe�ɀ���id/�f�,��D�Q���)q��Mf)#P�+q�Zf�12���WN,
�p���������-����a0Z,ljbd�"X�H��̙>�q�8p� B��&(��%�L�%�ɄJb-x�e�}s%
4DiJo��]�z���#-�����Qd;�e\��,�m��8��T����-� �54ft#�!�M��H���y��++�=�^t�`��m��/��{e)�^8���������\������[4\P.���׽�1b�ݳ�#�x'���:;6�3z0n�2@=�y��z��ҁ�sn�pX�0������y�t��X�un��zF�ӎ
�MUp��)�3VT���CW6�ٗiM(�ؖlۭ�6� �^V5��÷�p��Lv�����Omqͧ��Wq��<Bv#�	y�9�]zu�M���L����8�]b�7[w�zVA8��4�z�����W��Y1nW����O^�m���F5d	��}r\;�g�m�;���Zʯy9S��F�iˠi�Fn\Ҕ���K�a]!HjS���,��*�ȜBu�E�d�ǟn���=��sh2@bݺ�ѕ�D��%��h�-�vݫ��rUv޶]��B�;M���aiD��2FK���stX��*��-��iaݹ�K�[O��:Bu���!eq���)��L�1�@��v���GZ�ܥ��7b����r	>zp70���noɳf̧gƑ��Ə�w��b�`��Xc���yW#xэ�����.��>��.����}��s��t��˽�Ј��0+..�Y�*�@n����G�9��1�tN��c�&׮w83�y��3��j�-,B��0�����7����ԕ��J�UUUU+T쵶�s�Mrq7�e������К�����n�q]\�:����w�&�`�1 (@�a�g1k�֢Ȱ����k �Ԁ0���
#j4/ala),!�����Z,ya//(�J �����,b�A����ڵ���а[�H��T9Ym� ��l)b�(XѲ��(��H�@h�j���˭Fj�@=w���-��gq�n۵������Ԣ�X�D�>c��|���8��u�^�}�+-�O��Nl�,���CԷ�|ʚ�5�-�y���b�[jdk�^>g��OZ��y��ߨ��s��ս�Q��E�̏���~��W���Tm;����{����ųm^�#j�( ��!Xj�l��a�xf��ML�ʮY�k*�b�ջ��r�O�Ǥ��y��[�cNM��������eF�ٻF�r��M[��z_.��z|\|�A-�M�1j^�rEQ�o!�a��kMm6�߿��Z5����:7n�"Sר2�pa��(�&��=0��Ui�ߜ݃�����N{�/@Jmk��U��w@X�|6��x�=>���i�H�Tx�Z�!kt~��4��W�^���s߿]ɋ6��xԉ$�d+�� �m���1b�1b�V?�ʟz��'6�ooKc���Bfa�=z��1�)��i����v�d.Ϫ'Ϟk�~�z{}ٯ>y�v���MC>5۷��Oy^����H ˰� � 1�#wZ=�v�,�|;8ʊ5w(���MH+�vH�d�����[U��ϐ��^h��̻�A�m�k�G�v1hP֯��[�Yk�_aGK�s��
�ե$4���L�ұ�ь����2��_�7,��ę�3�|�L��y�iV������l>�� z� �
W�q�(��������dۭ����UZ�)�_��4�$�l,���2i���|>�D̍���)�����7�a�/wW����c�'dSyi^��M1�3<Г�+����{9����7���}����r�U$�USd�r�f�k ���n?��c��@TϜu�õ,9>y��\AMʀ3)�o23�5��{��i����駬�6g[e�����p(������}s��t8v�r�2��,�|!���P�`	&W�L-"����Ȼ�̴j3]�����>���.��hI�HZ1�hUDs�6�E���䷞�}�y���9�%�}5~��5���I>F�X�9-��-�d�.��I�i������U����N�$��Y�s����z3+�X�kY�,�b7ow���$�!�a�Igg��Іت����UPo.��z��RR�-2�5�j.�H��'ؓ�MRhH��W�>�����&/x�~�:l\)y���v�m�_��^�Y�^��+�0���]ުi�Rq�<���ŌS{�����]���xt�\�w|�lV��BF!�3���Ԟ�b*�y��<��M_8&Zz��ߤ��ߟu����e��������F�Ah;��E��|N9u�j���"��gF�i�*gu٢ ��C�����X]o�׀�5�]�KB��y�Aͺ�9�v�
j��цkv]�KS6���>�A�*�y��T�g�X�3�
l�̼�����nj�4����fQ�}%Yڵ't�lI �h��-Jd�_3��4�f}5�3�9��^� �a��&m��[P�q>{9mE�����4�E�ۭ�����DB� f��@�	@@�*��S���!)���ߥ�=�[��[�Z]�f\S�UC�5�g�r�-<�Z2I�yՂd+"�����tE���ޢ�4��6����<l��'�Uk�p�S(/�ic��J��1剻�$�L��s�xM7�G��l
M�Qlm�U���hx�m�h���<f����7I��1 ě���Ꚗ9�z�>���5۱n��ű�����q�K�3&Ć�Q۶�k��b�^�V#<#�]��;��ڹ;����`&�48��GH]��w��qg��ݶ�6m�k�8���kI���HiX䨋L+ͦYa)��+6�ٰ�E]ƀ���f��٦7:��ƻt4�5�>��ݾ�sS]�H��j��4(���v��6��mb�7|������-N1���VW�g.sљ^d�bpc�9��Ґ*�	k�2�m���ݙv�I�o��`箫z���U �N�W�h+�8��$���Yd|��N��ʍ�!��U���enj�iD����j�O� @b"8���}�w�505W�&�'6fr/=����;z�z��<�c�<�ŋ�E UT�����-J��b^�������Zg�oy�dF��g�Z�3S�5�v��؅��3t��{|X�"���m�����ٞ-�B唙���m��Iz��)�n9�Us�4IS��y�'� -w]��f����3�kgD߽�`ݙ(	L�f8����A^�ěZ@�o��ڈ9�|E�����g�s���9k��o�s���y��$���f�W�]�|w��P�8/s�צZ��� bcs�Ծ��qw_zI���~�����EI�f�`'����L��2�p�%	�Ƿ����:���3�U����E�Ii���@&�P�UV�?���BƦ�b+2��e�.�����Ɍ=˲^�t6g�\�ܳ�RM+df�
�3kveN�y�17��$���2��;�#���w�E�@qQ<O@���cz���~�h�5�.fJC��gucvY0vsʓ�hӞhj%��eD�O�[�=sZ3�א�%�t�,`m ��3�T����oQI��G��#؂ktQYV�D߫ٺ�l��|����w�q&��($�!�T8�!&�L�/Tf:!�Qu�/+�b���j�8G2��|ɠ~�����~�S]�ݙ�����L{����
ϖ�{Â��i�#iik�����"yJ�gw�fk�c X�,@,C^+���S����I+)�	��
]���������Y;:��<�;�Uj���El����t��2�ږUӸ�
o5ݦ�Pr2��$b����n0@�{g�����o���{yiA�K~̭�R�y� �y�) qo��'ɐ��]k.1F�,��ʷ44e�]�˟<�J_$���8�;�3!�B���I���>�����Z�'�$��L\3�i$��6�q�YrІe3�X����;g=�m��� ���C�#�����9R#[t{qcC;���Ҽ��0-[��� �LS��T�+X�;�ּ]ݻ��z�(�������L���kNP&D3�Q�{�)���@S��ѭ,�����n�x��>��bR�҉xVs�vf]mљS�u�l�l�籎�a n{g_j^��y�hZ�1���/a���_*�+��C�����A�bC%�}��q�m��ro�L2�{56�l�*���9x��@�V���3�	j�Bb��޴�K�NAp�pW��Z�)�Ko��CL1!h#�RƜ��΀n�b�#)��r#%���i?���fU����;=kĽ�V�g;h	�9`�ܲ�kdn�0n̬!���&:��&}��/y�۟	cDk�Ůҟ	�00)E��@�Lc)XA(�UM����o�wDm�^-��kKE�����	�j�Ԅp���v�l����d�D{ok�fUm{7_Ϩ5�>+��5d�c�ݷň#Ͱ2�Ls2��}ݷ���^�L=m�};�/y�۟Qh�&T�cww��5k*���/�ǅ�G&�^`&`��A��Dg���mz/f\=�R����!���^�$z3U�e���5Yq>�2� z����O��CC�Q�dg���q�9UH���qǾX�v�sp�
�<o�B������1��	h[�ȃ�F!#����nr٪T�)�����́�Ҷ�(���V�=�ہ�uP-��t��ዷ7��k�D[Z흸�6}�kq��G�#�f��@v�	跥^]�\n�B_!
�z���!v�&�j��UY�Ŭu�l����8�t^ݳ�:��f��h��8��+��:��¤ٞ�2�C/�e�����0ֶ6
�mtI���Y�5����y�'�����(&3(yzj�G�v�{`��Q�ʸ@Ц9N�H?�&�t�o������
��gk0�7^[2�}��>��%�L�{N��i�.�֌�ă�ji^A�4�b*���s4RO9^�2��s��M2�����Z��]�WO$��%�@�v�������?{��}�g�#�/���Fi�3��\�L�ؕS��[���j7���9�M_:oy������ªVvl�϶1j�t�����(��F��6kr�X��M�<�߳��o<��-v�n=��/����>jϵi�%Vi����i�E5�sMQQ������&j��on������G��K�y��zO'���|�����ю�r�����Y���}��*
/ш1�A����=j ���F�V�/lCz�5B���K���GiW��[	���U��z��ފ�l���lʩ�f��?�fQb�2�T�H�W��{ߋ[4�+ |�����>g�vݜR�����ng�l	�dы�*P�B��')$��[U�qUJ�ʒ����b���s��b���;�SGX�G���__�5՛&Ia˙�߫���9oi��M��Ϸ<c*�0Rh@���]zָ�6n�*���yI���i1�T�S�VJ�I��{7_��j� bjl0�H(JP�I"��R�^��o�N����������~��������؃P�*�ׯj��V!8�:i�*�&���3 |��T�:L�ݫ�j�������U0?9���d��z'Yb�����1)g��%����t{�"w�Q��>�Z �'����'{�����}�2$��3��=�E�˾po�F�Η���->Y0v_<��D>���}@���u^}E"�+��D���h�}�˕~aR�L�����_��I^�����髽���t�tޫx���	���xlɋ��"^��ց޹�]�׹��Y�i��W�c=�O,'ؼT�3��S1��nF�i~f��O�=t �N�����N�z5�����	j�Oz'�J��:&Y��xq�י��M{'���;6L��K��˓�����`��%�~��qr��=����=ヵn���f������,�vL��;
C�\�������'`����92#DcF���{��nН��p����p�zG�Iޓ�w~��������H�����p�x5�3ot/Gz�E�|��o#"����. �Ş��r{7��o����~��z��i�oP�f��<�V���j��z���%��C���g�I�b�/�:����!�ѹ�w{��w�٦��17}�[���#�8]I��������\g=�î�O@F�;q|��	 9�[f��y�+���y*<rng����]�ǔ��W8�r0^#�XcSP���)Q&���0��}��̫��V9S�L]���ٽ���4�1 �I����Neb��*��D5�kM�2�)}���X�������Go'\u��<kZ��k�<x��Ǐ�#Ƶ��뭏sݑyg-��vq:��~�˷����,*n��Q�*ؙlQ�m�����m���u�׏�<x�ֵƵ�<x���x���]uּ�>K>s����~�٤���9j��i�ݶ)�����%�UMr�C��|��u�׏^<x�ֵƵ�k^<}y<x��]u�Ԟ�g,�S��"���\�߰��gĆTSe�5>�t�PH�B��b8�3V���NM�2jd�r}<�O�ֵָ�k_�^<x��]u���b�"�U#^0Z���`�֣�m*�	��nX�eUY�B��UUkP�|�QDQ\��4m�ҳWm��%cp����3j6Ղ��n�4�)���
(��q�VڬU�bcj��\M��m���Ԫ�!���UTX��j)W3&T�4Aq�ʎ2�ZR�eT�Z���ӡX�R���ծ�b��n��c�
��<�9[l-I@EUos"�%J���\��,�b�"�AQ1��Eb��j�X�Q-��bɬ�*
-��T,��~Q�9qR9��W8�w~g��'ko��o�;�A�b���h�a��v= ��C�Oz�si�T�$��a�q����w��k�＿��/]پ� �c��b�uw��ֳϹg� ����9�Й��/�u�/;ut�E��ˇ���3*�w�O������QLAj���DL��S���Q3��+D�*��9�Oc������[�l�;���jq�Av�@��b**���/W1��ӷ�������Ē�yo����ڵ��'�����4�6H�hd�3���B��cop���E�!��j�b�rC"�d#5��U`oZ��T�-�����R������z�m���"�b���]��],��}ݶ�/�g�pD|�3�K{�ǀB�R��]�=���>�{5�#ٜ��ME�J,PT�ZaN�5��ȁv��l�L*�&b��䁌@�0��5K�燞g�k����-�ǐs�pu>�j#�d$�Ay�[�����b���g_��K�{��O��}�����]�����Gۯ�P>������icH���2��-���o܇��̶q-���i	�`$�oy����&"�3��J�/[ٍ�,�S��#�����y��4����#h[��O_~�W��)�ց�fCE������giw��g��L=����ǀ�ud���S^���G����1��Zzc�gxz?0�G�������&�2�O7\��V����k lQ�M,K��8.�ھ�-L[���8�A�~ld�����C<z,C���u$g`�Y� �*cd���0��,����x�f��t��e뽛�އ��c�L�I�*��T�ao�q� ,-g���}�0�Q�Ȋd�3��jk{|����}�����>�1��`�zЦvL=�2;���y0�D]v��r�����l �4�#����g�}� �;>�V��Yf,�UC	^մl�-�9�«��j�Y ��-^ʸ���S�0a���D�g���/��w��������?_�
`p|iX�()�E��D��`�8rxN���Ow�#]��f�Ԛ4�{�Om�,��g��73	s-1ֵ��~��X�2Ƒ�2I��a��ص�q,͘4B��,[l�2v������ҩ�C���uc���%m�*��vj�����'8��,\z��Ա�,�U�k�14u�p��یv����ὧ7[lpu]��;=��kS��nJ������JF�5k�f٧�:�]U���Ϝ�8���[Z]4`M�̓)n�]v�<��1��9�"�#B��a��*�b�C�K+�U�.�*+�7��)c�K�%=d���3�M���0^r����D{�'��+��� �N���41q^zcL�������}�Nv�!�8Bcl@���n�r���kk�^�	%�|��!n���5�6�5Jڏ�y��H֓� z*���]�� I�-A��V=� �jzNe��W����Զ�7�%z�}���<�W<�h��X:�5	��&涸��r��?	x�{7=�\��M\h�{F�0E�� &S�A�/z6�0��90�yL5��A�g�����S�c� �$�341�Ȅ��	ӵ��/���h��CY	��L�RΘ�ԃdON��wͥ@/ ٸ9(m>Ld�3U��( �[R�C�qq2�R��'>�ދ�= ��'��4�������Ǫ�o	<z,�E{�v�@`��|k.��v��;��UÂK�u���w�=�V�_Z�](���Q짛�\ӕ�(Tf�<w��p��5{#�ݞ<7�|F}FX�����!F`�3lpxb(�xʺ��&b��{Ѐ,S;.�d�R�5Z����ɪ��HxIG��8|1xMC�z�u�94Xy�1�(�;�=��>�ܹ~u�CN�|�U{�7n_���|�:�[(�13���y���)� ��Mw(l�X^��߾����ܥ�Ñû��]�ȣ���-����U�6<a6���D������U��x�%3��2d��<E��`�����D"�A�� �X�,�v�CU=>w�:0 <Ń��ܜ]��V�o�Sc�Y{L�i��&m�
��֣w$tAz"��)��0b��>~���g1�S\h��%\aH�̬Ȼ[�bTJn�o�_���'b0"����1qv�&����yڬ��4h�*�FZ�0DcAK�pD�"�i7i��v!d���_�B�0j!����	y<Ǯ��tǪ�o	<Xk�X��8�XPG}��S>��y����Ya�u0[;L%�4i��y6!�ZZF{�w��A.��(�ʸo.y��v��I�$��nj�P?��JL��(J�|�WA���*n�*����X�/�nd���K,����Ǯ2�x��f�и��^h!��NQ�e<�y)�t�T��OuM�!�b,�0AN�����������h��l�3��)���b�F㳵�ľ�"�`x]�䷽�0MS��{�r�ڽ���������)�]���'Ļ���#ϩ��빐�x��(����\���� k���;;����	uX c���5Ҫ��۲� ���~��xv�W�O��"�<�aDsZ����]��Wvozm��=��Z ��#ɱ��RЃ�Wi�ВI@��|�P���<�����>U�\�����2�Y	V��\����g՜���x>1Fxೡ��w�7o�:I���kΪ��]�����ƠŎb�ϟu ��_`�^���1�k�� ���I�n,�,��x*�$��#������x�.XK!9���X�56CKH9u\���Ovo�],�;I��5��f���9x��Ѣ�k�4&�,葅L������`a�<�{�/_]�+�^����c�6�'#H�),��e�!���%g��*�k����{l��9�:l��Aزb[��
��ט��(`۟f{��}Yϼ�F��͗b�R�q4��8��W�|8|<��U����Z_Rr����6X7"i��e�k���]c^;%�\e���h ��H�L�cF��Mf�S@��No3�����b�K�0Oj�UM�c|���񓽧'ފ���0���S����0i� a�.Ʌ���n�w������.�@�N]�jL�I������2��^����c���4Y��p����y��Nv���Ug�},~�>���lx��N��̇����PdZ�"�+˪f&U0h��&	&v>�|��\�~����k�� �ıX��䧷��-�d���<J6>O����E�0�Z��c`N۽{�3Y�|�/e]�&j;�{и��*C !�R�YG'��&<N]���*ȵ�l�6œ}�����2n��0OM��l�����.��T�{b�18��:�,9w�c�b����'���{7b�m�M2XU�F�Lk�|��<��9�<�/F��t��bA5�mه,���>��K2RYf̎,`,�L���Zhs�ۭ:�鹋���:G���[��i8����h�A�Q�k�ꁛ5�Wm���]���V���s��8��x����,�QP4H��m��3�@�"���^�؜ccC��v�&Ӧ�]ڵ���݁�ힹ�'k�ػD��͢R��k���'>?���9�L&�Й�
�1HM�˛n� g��R�}�ܳO�����Z.��`@�zc/=����UgF�3��V�+ǈ��U�	`�X���.;�������u
c&�.A��z�����Eb����*+n�o�A��0{d�e��"�FvǕ�g������'�j���S�}��կ������9T/v�γگ�MV�f�Й�E �Ʃy&fӌ�Iq���bs�	������[�:X ]��v=�o\Ǫ��zX��8d��E�*'�݁5���'�;/{t0��<��{�X��R�rv�,�@@� {�%� \�ў�⢶�v��d��A؀�s-����An�z��ڶ��;�R)ӹHZ�wߔ_�fhѡ��j�kO=Tn�=�ݪ���:�u]s�a�>��D6�#3��ac�p��5;L�^Ww�����z72a�宜��Mebp��Ʌ��N���)��X� �=\���UHj��]���iqy'��G�hU&���¯_-ܯ��QQ}��8Q�P��x�Sc9~����#�Zy����!M W�a�kkg��Iخ�r�8��뮜�l�%, �jH5��/�*����mN}�Ѫ��E���0��g	��J������f����d���G�,C��� "�ޣ 6t�e���]��0܆2�}���#�0���"s�"o��:����n��\�P'a6��ϳ�=����e�Ge���}q}��z1j�go"�l"�#�w�0_7{�<I���a��������;:�7��zy�"�	h����K��:7�5c8� ���RA���v ,Mo��O����!�⤨0�տd����_����B�Z�Kh�hL�4!SCY�H:�4	o6>.b18#er�v���h;�s�T׮��ۓg\��şM��L�~߰�}C9��Ĭ���x�K�����7ٜo7@oJv y���gbQd��O��z��7��&@TÐA�Y�
�7;Gzv�����&��v���!��pA���-���\�>x[���1�z�?�����_�iK��I�^k{c�����K&���3�6�<�18�C�p���770
�p�ɁRI���䳮+��
-%���� � 7D��mK�Nto�F���U;4ԻA���M�ˋ�vC�/c���i��<�G؜ݨ����S[WϾa572���Z����(CG��%,�Y���!�i�
��p��U�{�ױ������PH)�}��'îo�x��U$��ڠXIo5��TCg�_k��e=������)��cX��$���>S�oɇf4��4J��JjC!�fUͮR�7g��H����.��@h;S�v��/���h�ý}0�(��Ao[�r=KH��n;+I�]�b����W������:�,l� #{՛�Mm_>�A�	�*f`a���F�k�[�ԑ� ��'IM�Y~KnG��s\��s	���;�;,h���Q��7پ!�EJ����f5���{۳��-������"�:��0eX�L��>,����վn�ez��7�7��Ł8Bb=��z���7��в�^N�<��U�W�n��l>�;��'�ٽ�<|fm<i��r~]��H�:����\W]��U�a�U�H��$�%�ؑ��ч��"Y{���B/8��Y�nԵO#}=S9����{����*cn����oB�0FR�,$�c"�����6��>�%-��>	��}��%ɔ�5���v�kz����Q��2��A<:)�R6CSZ���L�HC���Q����3�>\E�}��'��y	~��x�Qӓ��Q��0�ޭZ �G1�,:�=^?��K(��{� �uS�����M�o4o�fB�ÑU�'e,u��)��N�Q.��"��g��T��1�e���1
��w︩�]��� ��)oS�@�p�kA��چ>b3���l���0j W! �1 9����T�W�G�.o�x��!���Tؘw�������.gdZ��n�U-��N̳��:�/W����|���21�Ƒ���&��{ޙO�}�?:�Snsx}G}�5f�	�B ⛺����n��"�b7�U"f�L���W�̆�;FP�t^����ߗ������'5�v̗^n���D��@��XO�M3��a�gt�T���w/Qٕ��}� {7ٳ=xzE�J��>�W����&M��}���w8���^�ux�|�m��i9ئ4��>���N�}�؂��1�������[�={��g�f����.��ǟ�%~x^���aZ~�^���w��ܢ_������y�̓(��Nz��/{}��w��;�c���6�;\͎`��G����a���Wa���7��*m�P^O��=fh��|S��g�www>���w�����=��{�)��ú&U���3�	7�b"3�ٻ�[��GUGJ{.4v�;�������|�M����������4F��K�;;��NM.7��=���S{ؽ�-��4�W��	�/�k�i�wz�gnv�#{A�x�b�ۓ|N/n�s;G����FOU��
���1�f�s��@#p��E���:˨%����}�'aꤙ�v�a��=o�V���a�WY�>�����F����� �E���ۄb�� ��\,�E\l���p��w�7����y�Ϝ		D�
��.����4&���9mݻE�k�V�xAݹ	�o{�`v���|�t-�4[6��fM��/Å� )$� h��4�t�1���֣*�A�J��r,�j��i��q��0%0L8BY�ð�x�}I��7��śp%���1@�Dς���sNI�x�z�ś��9}����ca-˶���b�kLc/U"-��)-��:_��*�ln�Ƭ1/k��,�����,H`q��%+L$��L�$o_,KkH�cB)��N��b�}��D{.2	��X� 4b�[qg{�<�w0	{�CK�����6���2���-�>=�;[�ҼF3�aR� �³~^�Y�q��XF[��V�0ez���3qr�s:�4v�,�~k���?`���A�q���h8�}S3-3W=�?{�֦�**�m��"�~�PQ���b(�~��rr,��y'/,׎:Ƕ<}x׏Mk\kZֵ��j��ǏLu׏�=ڨ�3fpj
GMR��YZ1ijT+Y(�֨����˝�~>��>�����Ǧ��u�kZ׶�Zּzc���Y}��Ϡ	��Ds1�T(�,UQ~��TUAI�E�~��ק�}x��Ǧ��u�kZ׶�Zּzc��|��;�W��KVYl[j�V�Tc�Y����[l����,��8�����Z׌kZ�Zֵ�{kU�kǦ1�'����aZ��A�E(�1�u�U-B�.���[V���������#$c�"�����ģ�JI�*��#�Q8��
��QA-���X��U��(������.�X��m�^^�[i����wk%TE�QQQ���Ǽ���ùTT���DRڬb(��X�V(�e��ENR�R�b(�X�Q��\r���
'.�mDDb��q"���t�h�U-l
�hΰ����UG	a�*��EmC�fO���n��QWy������ܺ.��ۚ�W2c��������?=����,�\�.�H'�ݖ�kћ�K�NP�f)t�L���8dŎz���ծn6LX�V3�g�z�a��1y�������j�BQ�,�=�-���#��`C���7/K��ݩ�g87b�L�ܩ�Pح��63M��-^�u��c]X���9�We;c�E�ח���F�n{8u�3�ˀ�H] �3
h�5n9d�Uؗ�[��6x�=�jq�Z8�q�p�%���Ps���C7���� ��^=k��/i�����{U�9ݜ�uγ��7V�v�q�����v��8���囖u�M�^�xr�A����V	m�5���X䮮�!�/'>�Wm���JYd�z⓫u;B��֬����1\6ܼ�Cv�� FY�d�5\��p��烊�Er/v|��n�=8��ᠣ�B\�B��Q����g��*��c��:�9d��v�8M����1��S!\�����v�x��R^M473%���ݪP7UeJiڞ��6�I�X�]�^�q �ѳ%r�%������7.}Irm��hc�N�C,��@܏���8���r��Mvv��6�gksRq��[��̜����q�;Z��ۃnh<��]�lx�pg��i���v'��r4�`ǯ�kqM(fXԲ�e��BfkM4[��/��,�$�]c)�ɹ����]S�/e�5����UUUUUUS�u�=s��v~����׌�g�سy���;6�	��$;�n�woU\�]��ä4��	�,g� ��$��#�K]q]vI�I�3&CE $&�����ºݳ۲qu����k�8�4.���Q%f@�+*p�Hh[�ΓN�myg���q���WPh��u��F��A��%�e*�0�h&�h�E� ����<8
�������ʂ[==u���g���ی:Y�R�	ӵ`�s֔ݦMZٍP&��ļ�l���Ԝ��~�}	,6.����C���UlQ��74gc'��`�� �lV�&��8��ݡ�`�g ]�}�1��}�c��n������Rfy�x�XT������!���ٮ�}��?&�02韘�%�2}u��.n�yys1Y]  ��U�F� �.�?\�(��|�d����V&����g{�ǉA�=���#�������̨ٿ>��y�ĝ!؀�ݫclBH5H4_�I'�1Y�+#��q����A�k 7�X�19�[�*co����Ѓ��Ͳ�T��	�Xu�)i}���59�\7u��ť�R��E�`��偀��=��gW/���^\XK��Z  U'#Y+��M����7d�T
�gI�8���;���Ć4�.B��9�auص�8�4�L���l��_!�����!T�"a$��é���L���>�F�x�8��.��H� ��a٢B�w�i,�4ԭkUu�c���8,��N�WEeS��Z���q�
k�8+�b;����^���w�}5�sv֧�wR�{ӽz�����8A�`�*�xc^p����~�Fr`,�]v$������D���-$%�$쌯Ŀ}󲥻��߾�ߊ�߳|�,u�� �z@6C����'z�'�np�}���ɶr�=�ghU)ld,�v��2-���b�sw���"�w5,)�?N�]ݢ�{yt�7g�{�������V�7��s�����#)ê���Q�}�L8�	������h���A��Q��U=Ai5�@�Ja��`���Q�u��{ً|��>��-����NX�	�}W��dp�0{%@B� ()Z�ߤ�}��d��>��k�Q�3&��t�秥�В�-oʁ��LA�vj�v"��.&zk��p����/? A��=wy�!�x�4��؀��4��L���!M��Zf�M�o��c�"����Vfo�Tzo�y�y��(g@v��|)�WWצ����ަ�ė�x�d��ř�{�I�YP
N\��1�o����VG��F�*�a���C�5�Q�;��|��jd��&)X�s(B|j�$? eD�����q�uԑ�Yq]vI$��!'l	;#�}����^c�1o�9���,�;QX]�s��3y�k^f�5��M&#|�j!�V�� ѵ5]�xdUvr��-R��Ć�ϼ/����'��<~�`�ܹ<1X.
0�����8�TG��7a���g� [�n��T�s�y�@B؀H�S�V����l�7r��Y����xt�c-�ܜ�Ͽ��җ��WR4�5��4�+4L��&�6be��\�]f�=�<��'~���d\��cR��5����;ً|�b?}�Ϸ=�����'�j9��şg������~ٖ}��'r9>|��W,|^�l�}H���Xm&{L��j�x�Ȫ�����\r�i`bu����]>�2S�� i�E����{ �?S#ؽ�ǎGs��:�g1���1�E�<t�Ns�&B3������S<�{���j0�n�>f�}��M�|��P�-��lh*��ڋ̮���f-�sņ zP6}�6J�#�$_���/�a5'w̌맊��}���=[U6㝏�^�<��y����nN�h�� ��8����\��S�0o����jI%�N���"'W]"N:��	�KK`O��l��st;�<JD����ߕp�t�|a�3����q�>�&��*��	l`ňB�+��[�Gx�ɻ����)�1��-3 ��uN�wR3@TX�D����/�9|������0M��3l6������CK�a���l�����9�{>0���1����Q�����	\��ռ6cl����}���ra��2}�W?7�⧹|��nϿ>�ϸ�#��y܇��5h����y��ü���FS")�=O/7��F;gC2�}H�![e�Abؙ둵�qX�o�x�ʻ���Zey�0 Jv!��N,��Q���$�-Õz�5x���PpX�v��(��ks���Nto�A�ڇ1��#DQ���АEqd���F��)z����ݢ��{7�&@=+����g�3Q�N�]��ry���C�/ڰ�9>�1ЇS"a����l�Ovƙ��K�z�M����qgɛ�9��3y�����9<g�}??~����2]��iY����Zq:LK��YW`�ݭ��H�|�q�/:Vj�&�sR3����m KW�����θ�i�c���Ya6ǋ]i׵�w�3;�����U�Qu]vHv���:��;R�Il�-�$���^��y�[V���QT��Fܽl&Wq\�q֙A�&�r��qcm�-qP�i�xzNuH��(6Sn���n����I��@��+ۥ��j��3;Fq�z�/�:�#����1�Ύ ���Yḁ�c-�-f��n9{�i�����������<�NY���ߜ�x���`��� 1�Z��]�K�Uj��=N{����2��|'7.�ׁ�aR��&��J}q�<2��yy
rAW��ج���Z�ɱ�u �!L}�� HIڙT�Ӡ1���{@g����L�}h��}��^S���K3�	�!UF�/�HK�`c���u��d���G�kx�9a�7��~���b6�x���玛�;��Ѓ�����t�#�g#�d�2�0���;�=0l"��`��p/	Zޫ�}��+/��/.,�T�2Lz<\���5���%�Q|����!^���ۣ��d��v�����͑C$��r�2d��22.���^S��Θ���;4.�;v��e�����f˼�v����۶w���'>�����5uqe����b)�fN�f�%�i�:n�&�;�O�~����1��;M*��[YǞ:s�7�#v��.�`ӂ}�'���i��g:���,i����O[O[�-4�Ӓ���;�e���4*�c�c�AM��&l}��M�t;x[�A�m=$��O��oF�������h)��n�������I?+��;�W]�ڄ�밎�Z�q]v;Q-BE�) S@s��}i�X�L�MW�=�#u���/.-R��"�igT� ⬏O��f�ɩ�qF�ܦI`���+��YR�޽pe+��gk���F��s��D \!-"�waU&�7*؎�9��+` )vpX�y24 �p ���յy����7���=9a*�ݴ2��n�&TX;j	[���RJT! �+؇�Q��A�_�������BX�(�d���4����g��!����%���-
���[5���a�"�'7�=����4�fP����qb��\��^W\���ݟ9�xn�T�)�t�@ Y1�B�*���':7�Fs�[,����0n �X���"�wDsk�A� 3k�r�*wC6 �[�al`r��noں#��f�b)���Гk ��,#��l'c�������2���<�~J?B��pE۳�6���:�'��n'b{���A[o�p~��uy�._�O�=�ŝ��0�g�yw�"�wW�F�9yg=�����⾺I'W]	8�서u]u;$��R	虿G�]e�����昀h�q�XӎNbqO��TxdM�I�ǝ��s��L��gLt�,\S�1��{��|2�w�9�� #M��X�e�X��In�mYĐ�.-���F�ōڙڿ��fj�F]no�"��n�G��b� �^4�$���z�z孾�v~� �l)
��N/ߗ�'����v�#�s���U�&'��b�U�����N��ԯge���j��������=u����g�X!&�ojO���adŠ�V��g�-"^�I(e�1@ܦ��{���2,���)�S�3β�et�Np�G��H�,�b��#��ӗJV��a������;5mr;QҚ�41a'�G�@!ϱ8�ha�l��-&�8�.=�|�;�6�vvtD_���� �/JaM(<��*�Xb�����rbn��Y��ƭ6����o���z�+���1&�I'�nS�9��B�h�T�EK��YF�z���1I�+�5Wi��g(k���g��*/+���ͧ�Xu"��/v]k�S��4�2(��|�4��K#��ԓ�"���du]vBq�u�E�#�2�~-����#�G�y;��Ⴠlb�X��n,/�^D՟{�'y�CS*�2���/FWN�K� Ɖ'��0��0�L��h�>f�P�8�m8����[��I����~O�f�5��܅]�Kv��a�M	��k���FF5ޠ���*�b�ݮ̜�r����& ���N{��C�Ab�TF �	̻��3}�	e�సL�����c��ez%�Ԁ�LmL�v���<�.�a����q�N�J��K��+(Q�lͰ���B��_��c���a�0�M<� ��yc�C��� ��>勯�O�|s�OR��!��&�d�rhb�G3�$HZ�b�+ƅ����u�Z`�&L�>&k�ʇ]��r�����!��C#9|=o>�	�Ӽ�a{.��y�F.��e��b&���'��[]� s��z*��٫�򫷗��;a3U,"Hj_;��%%0�rUĻ����9�0��w�CR�_4���w{dj����E��������'gLA������8dnkYiD1ct�p�k_�}%��yܷ� �k�>�.�����G,��q�Ő��2̼������?J�;�u]t�8�순u]u=����/y��P[�n^ba�a���t���m���d�J��e�v�7j�<tI�y�_M��L�S9��ָ≴^7pe���cj�`�#,��o
��kN�8��+��J�o6�a������E�	��
���3e�q�s\J�j�Gk��m�{�;�|�����#���l;P�̺⛙�[��b�0��D��ݞn_��2R���?F����u<���^��V����ӜU:.@��H-R���5��e�7j�0�����z��k�a�@9��Ws~�*�����G�vS �i$�����@������[��ˉ\\u�!�Zɤ�`��N�ðv(&�h�Q�Hʘ�)�+ʧ#�V�˯o/.d��I����A�N:$HC2G�ٮy!�����[���v�Q$�!5�^իo�'�y�80g`@:B)���t�F���g���O ��R%>�c�l��!�42�F\�z��e� CHK��fw*���Ry�d�/��0t�伎fc��g����<�Zt�J�J�����-��nf�@7n2�t���W�2�f�\��~���g�q'��q@��h!Uw����yu��ˌ���cg���̥����)@-T��������y�c��{*�L��Et����7+uɨ�܀|M"t�K�>��.��N�%_��8X�T�m�<!�}�"�g3i<놬��&��'�������D�$��N����d���I��HH����g���/;9����}�\��=;�9�A���j[B�p�is�k�,5�s������L@v�Oi62l�V��e2�n�)��w���l��x��IJP���md0�]�o�X���\:�}���"a�'�P�����B!�rt�b���:���E�W�]���	�NXE�_�!�1��}�{��Rc���;K^��v���T��]�0|p���ūo�g�x5`��T�o�'Y��5l����c?	}��~"~C̺f4��L4��G4}{����������4���a�Q�.�r]����X5ɸ�;U?��c6�{������u���*,�͊mv��q�⎉�q<��7�U(}�����av5wvJ���%�0�L��L�t^��yu��/.4�Ʌ�XY�Z�]��4o
�AR�I QO&�u���+�~ہ��g�� $! ׹��{:<��:6�fYG ���;O���\�B��{|������ܸ�O�ݦ�I�;`��`�)�t�4��f�T*rW�<������s��ҥ.�[�_so�3�@�I��Yç5��Ӿ�OU�:���k�jђ<��Z��W�G�e4��
�����Oj΄�D��n��
�uq��)�����^�C��Ç��  ��́���s�[�b����.�]�0Gz��/����k�����޴����fz���=ǽ�/&�оqGO;|+���h���wЭ�r�>�=����3�O���4:Ǩ<�{�{�[��x��)}��7\�^��4HS�I]�������A��n9���5[/?�V_w�<��uҍ���Můw^�ڪo����\�{���O4=���%�]x�sA�sf,M�K�'f�v�1���z�W�xby�{�m�[J�Wyg*��0y,�����绔� My�X����;�\>������޾/6,N�:���= w��������݃�[��n��-�#����j\�d�{׾^���9�8r���XqT ��	Ŧ�Y����d`��X����l���� �#3"�)Ev��a�ڧ=��z͸�G)���<LM��6�X`���S�Ҳ��Y�K�i�.�k��6�-��]�:�i̾�I��S&�@�v�����0E��CN�AS�-Ķ����d�Ƨ�T5۾]���S�ǃny�Y9˷L4��ڛ�MPӎڒ��#����C��-?h���7�Z_��s�:q��ٻ������ZAb0�6���"�k�ȁ�e��Rߗ�,�[g�8��=5��ֵ���kZ�֫Z�<c����(zʨ,����E�ւ�lA� Qm��U����k�r�d���X�����^1�k]kZֵ�k�k=1�>Ye��}���ej���UT_I�P�J�t�1�#���R{;,���O��1�kZƵ�k�Z��j}755>������*�U`:ʪT�ŊV�x�H�=�$��m�Y�u��oO��ֵ�kZֽ5�q�c1�$�b��b�Ed�K1T��X,�@�(���%Ryk�.��ob"
i*��Q���ƥ�2ʢ��(�ea4�F��oZ]ڪ�*f���
��Z"&���T�IiEF"�u��93r� ����"��XVE�**�TQ���#=OwM�T�8∊�ؚ��mh��F�UyheNV���b� P߷H��b`���
n� XY��ʢ�(I?>+�Ď:�����q�\t���KD�T$������|�����jϜ6�,�;!QT���1��L�
�C��!�@H#�& z�A5H��y�k���C����f���#/Ϸ���D�I�\��6����̱Q�`
�qR��N5
L����ǔ�Wn� �q�(�',�La���k����5��܊����;�'٫.5�j����*~�.q�p7���.�Gh:������:�����N{L>�!�%&����'i��;�/�g�xc\1��yhs���n�ñ�Yԝ��L�/Q)��Y�SϾf�7�%w�R/�^����;�b�q�T����r��I$�@�m�"6��d��&���9Oq�Gz���e+�n\��a�����T�Æ�[�v"��)̮�^^nR�1�A��1Š�bAP,Le�[�$ō��(cb�\�M�}�[Z��=;�V�tEmC����'�yz:�b���v.����b���ǵ@Wj/�D����[� ͫz���QM��)cr|��E��8��Y�� ��SR�+���"���$��\v$�>w�9�;��"S!�"P�+b'H��[�����Y>tv���=}'s�[::f�@��A]�	�?[�?�,����S��6�M�Z-��=�����*��湩�f��ڠ��ge[��sn�&1��>p����匱h,)ݟ��Z�!U�q}�Js+���1a/��<4u�c�m��c��sTG|��%�g/\�/�矯g��L@�B"�8��_��N�U��Y�SK g���t���d��pzm���`q,��wo�;���W~�u� B�^Y�������--��ݘ���̃�p���)7�X-Z�ً�m��U��<ǋ���L��gk���)̮�/ 1�+b�Zr$W�i!��4��BX�f��v�M�i7h5����USN�j��v���zw�W���4�-E0�DֻE���u��yO�[���k��v^?�����%��6y~�^ݳ�\�bZ��`����&��=��Db�Os��,4�2ҫ�1L�5� ��p8�,c�7�-�f�;�B�[JA��Rگ��'{1y5��̘H#�,ʫ���g;���̞��?��:�+���$���Q�q�	9��~w�����.-�O#��H��%Y�WU�[=�<٩K0�]ض��)cj�tiLbhѬҷYF�s�t�e�	k�պ�ci�:GLKP�2��Kq�ˣ�M)j�y��u;׎���2�u D�M
�q��F�s��x�5n�ؽ��d���U7���g�~~�g��.���ܐ^^f����W�I]K�^z)����jp+T��$��9��u\� *���5���;��4�T	jl�Gr���I��{0�o2v.ۮ��$Ā�^�`���t{��!��,��4����دw�������nd�qv���s�
�F��m	�%���	�7��>2� ��!hd��������_U�a�����[t�X]��	.�s*㘰�����^$���ۼ��q�~Rŝ���K�@�.y�{MO�<�s�	��-��vdf׳��Vy��� �X���3�s���6d�>��p�.�UY>�oy��vɯTV�������3��t��K&�-P�b�'��8�_���e�s5ԉ��=߿�Rm���uY��:��N�7��4X�L�+��[?C��?v��Rq'��Ym��%Y�kv���zw����v/�<=9�m�KqT	2����ّ7�J%Աal�Ui�1�A���u���!ۣ�N�<�n��Q�Q���^�ʸ�!����z8�>���?gs!��'��P
����V C����1&2�DCL����$����~On��$���W]qЮ�㰉;b,TO_m�磾������z��ڟ��9��DtÃ�
�ÃE��ѯ{�ka��	�Aq��-(;b�T�E;;M��T=��eg#9���������g�0��%�f' ��б8�23! �מ�'k��O���3 ���EOui�E�Q�1��h��G��m� ��T�U�)*2�W���K@%�f���%��XAZ!*�Ҋ*X�(�H�R�
�6e
,�+��4"�+��e>�	=x�>�-����[0H�*�y4����݄�G��y�G�<����zb�ĉ�t�P�,O�noF���CrgFI�� �Bs����Z��kc�C��X^1��N���3ݜ�o�#��d%�\Iav��E�U8=S�VT˿qJ�n"c�9q��߄lF����� ������j��wOT7� �,P�v�P�E �����܌�Wo/."$U��z ����'�8Fh}��Sިf��in�t\�i��d=@Q���f��[X�hb��H��W����xK�:X"��Â!����L�������dݛ�;�w�,^b-�:v,0�T���j�^��t`,��y�e?�d����٥60�9�ϹU�<� D�Էۉ��h�սLm��mƣfv�C�i������y�e��~Mc��W]qԒ��ɝ���ɜ9 io{�}S��u��Vd{�'4�c�<w`�2��y�\e�Qgc�S��h2���w#7�����Z�n 8;�8�ڞ�6�5���K'��fy�{�w��}M��Y.���NM�D`���[�Me�I�}jm�a�9�;���2:�9����ime�v�b�g��F���A0JD�B%�H��r�Ȟ�U��5��Ǫ���t��Q� ���{�}��__G�����PXT��_z6_���o�#�Sd{:[�)l�!,�=1�p�$�`@��!��.��1}�a�������G�-���X�L�j�/����v��2r� ���M� n�ٺU�lG~��i���_|���j\��X�L���/U##{��dz�9��=�ll�؁F:l-��<I>�Xsw��\�k�|2��0I1s���j���^�l�wk��<�2o7���쮷׻^�����;'�dw���{��&u����{�f� �[a�w��eT�o�h,����º���\vI+�����	��?��X����G]@�!� @�vDOl��i��`fF&Br��{�#7��� <��W��q@� *���|V�tx��\���e)�����*},ڛJ�.3��ɵɲ�C.�X�iӹs���^��ߧ�w�����+��Y�`]���������U�p�����s����cfCb3�[�$;DB) ]�.�y=�wMS��O9̵x,yc =��̯lzO������˱a���\�R�I$��7W�ag�:�v[j]��+��ST�)n�mvֽyLD{�R�����
�clz� @�NA�[ab&h�p���>��b�5nk/m�Iz,3cu�/7ױ�59�v���.BdR�gd�0r/�Ꮠdj�5RM,��X�F�G���B��}�.
Ӈ���������ɋ���5�g��Ա�{O��FW�+}�nz����Ѧ��:k�_ݾ�Y�T�Ͽ~�=|�bM!�vvY�:9����n!� �/I��p���O��9wUk3�H���=�����Ҧ6���5�V1�.|�t��S�yXs(_#1L&��#j��ͯ���$�1�qԊ�;$W]q�+�%�B�Hv���(裘�j�4�Q�, r愬���.,���������ݻ>��:v�!i�t���5�t���6���գRuӖW�YB�f��s���ź+��i\
��wH�J��6[g&�z��y<֫[w����nzmi����Kq�ض�.[	VnZ8�چ+U6ߧ~����~��C���l@)�P��"���݊Lc��R����g5f]��ȪB��'�ˋ�rUy]������g���eH"	0��T���4��H�"L�� ��`������,U��`�o�}����曂���(���B��L��m;O]���ؕm-��P,�ZA2�&�MRg5H��W��^:��g����˷!�u����M&���;�d��+�d9X�{|�]�@����{e��=J�!1���F{y*������Ce ��W�k��DGkA������B��x�E�wN��ZK�D3�8v�TF3�Li���w&8ŭ!{�����;U9��U˽�H�l�Lq�o�a��wm5���t_�6ʬU����'���!��b6��xΏ�"3�Rў�3�Gs�k��z7�2�/��6K�W9pAu4�E�4{����`狱�÷�=}����>yߋ�휩~|����f������؁�����u)��)�dX��K�Q��]���q��:g]������^܇���qE{\���d�ɝ�Bn:�%u��+���I$�w�{��ł@&Br����%W���ˋnS� #-ؠA�V�<�'y��{V�∦,�:�5 ��N#�?����s��B&�כ;u9����HPɅRDP5Ձ$�$������O�VI�Jy�T��pY����I�)hO�Ǐwk��[%�7��!þuz��iZ���q��̅�k,��ÑT��s���|aDγ�d'��}�� ��f�\C� �h
���@U�P{,�o�}�i�%!L0��}O�����4�z3,�1��.�:�&�t]i���1�[��Oǯ�u�1�H Q�*�E`����r�<k����5NX�1X� �-7�8��*�=剓�pG��b ����8䂁��������`�aM̽)��1s�hWY�{�fJl���!V�h-,i!U �ԛ�v�x+��8$��̳y�]�mк�Ȼ́Y�����H)�����l+&���_�+'Q�W�}k�w�Nre�K]��;m�~��Eu�"�뎤W]q�D�~���[��� �����N�Ml��;[ x�S9|N#�Ɛ������վ��a2N8r��È�=^�_�g*s�cT��1Hsi�se,ɋ�4��,z
9��ٜ|���*)���,��O�:�c��>c���U��G�����0!��L��E�
�P��aT����i�q�F����x�<>ݭH{cm���2Z�nʻK�5k��g����仇�2����O<9�Br�]�)���,b0{���lξ0m���&C�Ϋ5ڝrI-�Pj;�k9�p������cXX��y�W������YQ~j�g�S��A
�r�ݦ^�|^��#�2�@_�h;��^X��,(�T)������ه�}Gd��r�a�����e�h@,�p���-��J����;�"���X����\b֥�8$����}�Jo:�.>b�Z,X~����4��
��ř_lJ��Ӿ)����X�0``s�c������yɜ���54����f�Q����(Ÿ{�P�ZK3(CH � �ͬ��]u�Eu��]u�c�"O}͔�޵,E�@ݠ�Â1��-��=1���g���0F�5�<A�v���Ct?��	�$��WчPX��P������nb�mW9�,�S���\�c����e��V�"�&�R���5���N1T������[ݶ� �Ք�W�ǭ�/6�؇�R�`�����4��	c�,��K�f��)'��^�X��Zg�R��{����4��C\� �L�Jfoƺv����[rw�x$8��A�1C1�Yk�g�=�hK���B�dt�����me��5W�)��k�!��vp�Rd�ʒrºL^h�i׫^Ӧ�p����
���c ����j������3�Ɔv�֚q��f:~|n����lVۇXS��CIGQ�����9�y���0b7LJ���F/����<�� e	bw	�뵛�<ݰ$! s����i�w�!���<��7��������h����x��t�7˷���>�z�N�]��kЏ���78g����qa�u]�Ho�m��=w��g�q�>�䈏���7u��<I[����v�iƎ=J�#7n�v����rv��
�)�t���V�r�ٻc9�۬�u�Wޘ�:C��vJ��j����e��l�R�ߖ��q�sW�N�_j��/Q�(m� w�q��0����mv�yB���U#C�pR�\}ټC�,�ṱ����:4�����C��Ȯ)��g�� of�s�I����J���>�;������7�t�hpntĚ-�P)^	ޔg����x�e0��{Hʳ��/cDd�)|&o�ȴμ��U��N������|g�F��O��3՞/e��*��N�Z���xg<���G���l��-��S�g�P})���ѰF�����gm��ټ�<k��f
���ۑ-����}����=�u�a�mB����\ݍ�z�S��C\'���+��C���w�K=������B�P�U{=<��7�6���[b��*�'�n�+;O��}�}�Y�L5��K�æ�9����������p(���mZ�K�;�rg5��,Y��9���x��G� ʤJ��b��3�p���C	g��3�mopV�y5T�0�'S|h���q��U4W�,�*�������.�[#��f'���A�&JB�%`cn�� ,G��RdÂ���Y� ��VX^n��]Z��r��
]b�E�w˻�t��7���)�*dD�f�9V�=������_#�j�x��k��d�B�0F#������{����-��6�^��k�2h�7=�4�<i���Y}�r�"�6y-m��ЮVW0su�̄�Bm��,K4izik3/m���?�Ţ0,,��2cl�qm��ǥg�٦�s32�Ye��Xq6Ԗː�W{;c��m@pb��uC=�]̑��g{��y���曘a�P^JUQg�we������c�f�r�TF�,�kƸ������^<cZֵ�kZצ��5�c�1��ϗ�y��;.�pE&%"ˊ�5GP�䷑��1����mx�ֵ�kֵ�Mk\kXǌc�ϖ|���-Q�g�5�y��1gʓHc�Ԛ��X����x�Zֵ�kZצ��u�cǦ<||�l���qj���U*[5j������S�����^<u�kZצ��cZֺ�MMO��Ӽ�DPU-JB�|��Q�鰬-l�*Q�#9X�����<J�|�Y�'�m�dQ=K��@�Q�+'��l�'2��O
VE�6["�j0X"�PTH�!
��1��Fҏ��V0�wj�=�ҳ�J3ƌ��"�X����������T4��*V1�((�X��[���ܘ�rN���S+��a��+�̣�]���.H,�Q5��hG4�C$t�6,��*��XE��Ւ缝+�F�<t��Y�UܺS7!Lk(�0LP�晥�K^V�\h[�`Y�M�4o9Y1����q����]�����f�({.8�>z����v1���s�iӠVm��/4�m�jLK�4C�<nd�bAi��v`^���͵.��	�R�B4]3�ڊJcC��U�IH;�t6R6�x���IC�ձ��k�7f���uw
�R⇉�.�a�q���q:{0Թ��4��lh�/d�i䋗��Nȓex�k�k%�vc�ݠۓ�Ѻ"�N�v�����[���@�Gp�-��ͳ;0��<���-b>�:bT���.�H�m��XWk�af��B)�v��]���X�Q2 ��P��j�eCe�Pr���{M6mg�x�9ǉ��1�8��;=�x�^���;uOl]�BY�p���E1�8�[M+��Т�Vh�%&�V�J�s���^^�V|&ś/cI���7�Ink7kR'��x���\eĘ����L�K;]c�ڳI�!��3&���2��6���t����T�S�7kFx�Y�88�sn�.g���S��Y�.�{Cq����ѻg%��K��S��84�	mܡl:[�ļ�K �K��e��C96��ֵ��!�K>�����K���H9v�\
ltnl@�ݍG-n��jj������t�D���hӵ���˝���ic�3�=���i_^�kl�T�Y��g^��K˹�)��cyp����7,�d�fH̙,��ɒ����<ZU�W�;�je4,Y�fni1��Ь9h�!s�4��7�h@�t���ۉݵ�$t�9���k�y�y��cq�b���e���!\W;Y^{ss��y�8K�Ń�yBp�r�T�"��c	`��Ռi1���*[�Ƨvp]��u��6���J�cK�����ϼ��F�v�x��]�{H��Ӻ�ݹ!D�e�8�9�����݈�\9���!Ak�`*�ݾ���ǻ���^���(iÑx�;ԃ$ʩA��њ�3ҽ�K�,&[�����wm�g�b�XjA��]9b�h��R/�x����K�ې��`n�
�i#�}�����پF/�y�������lD$�T��dR������a�m�;Y���a��������������ǻ��I��!�X�y�NP��u4!T����!���y �2���vA4��K���~�;u�w��w���m�g0�œ,H1c�N�D X�qsw>O���*˔�A�ؒ�d�H!�~z�[�d]���M��;$mX�p�35���M]_��� �%D�܆*����Tk�}����Ct�qs�_o��z.��x����@9k���h$�Ȼ�1�,�ZDŞ��;�0���Cn�k���:z(	�w����R�0�>�ݷ�g�n��o2�Nؖi(����F�Ï�;�뎢�뎒��&p���p�Yx�ξpIO��oE�}�gm���Usւ
v iƘ�ۇ,"��B���Ǔ @�L�t����; \ �٫@Z�]E/@#�^w=���� �O�.O��Ќ�!ĭ��i�ys ��߷<sg4¢s!��f��^�������d�9	�3^�f�v���@��5\��ɂ�p��ίc���y��,\N�v���������a<L�G��]�Ù�~��-<�o�ۇ���R7��i�r��"���c�n(�HkGAY�xDڶ5T�	����=��d�O�[�l ��R�>��R����C�v��p�\XHT�y���{l���oK�����ai�0vvT�Ե4d���1٬|Zg��^L�����#չ���f�\�)5��@{TnZ��
��pXU&h���Fc����M�c���%�d��kVC�����<�ݎ,�!��ڈ�tZIۃ"��&�2��Y��-��4�qS��\��_����fB3'\v+���]u�Q&��7��7���o������Ń�1搆C�a�p���u��t���<zݙ�:r,�b���Rp�~�[��O� �����n���vy�1�,����ΒQ	u5�B2�c�"�������<)��gp�*l���xE�ntyqZ@9Z��e��ѷ�W����4��]BT�&�H�gg����]\�롳�6�\f�	n5����g
���s��������{��<K�g)0y�����{�j��a�c��H���mܦL�[�փ(ng�T�P U��F\l7y[h _��O�;��p�F�:�3�9��Key��K����qyjWTT*х���1����i,�T�Xf;�b�&Kf�,���5W�=��8�n7)�d �h�A��N�Li���fHxc}��"�;�;�'�.���+�s}���2�Ts�p�gd�k4��Ɲ�gR3Y>O e$z����-ͼ����~��LcMm��[�f�[{cciD���|X0��Ο����zk��]u�U�\vW]q������,Կ$�?"&nw���w���鑨_sƟ���q�X;�������Χ���;c�3E.ief�	��F���}o�R�G�2:�a��ϟ��ƣ�WD	m!B�q3M����0��
��A���럧�r�'v2��{�ALn���;bM���_�A���G�7*b���j�cf�b�ַ�JX�21�u��d7(��xzO����![��D߅罽��2�|�I?1��#�q����n�j�&5���m����'"��
�O#�k�̳ Y7�����;&=ٵ| ��e0�L�f�
��$�)�a�Xnӄ�N	�΢7�|���q݋u\��9�����:<���RhLݨ˭�-����q,��,�~����i���NJ�uq�{��u�{{;NV_����c�*d;���1���@�v���wM?���j������<�S��<wi���.O���z����������:h��z��SDVj)%�NDZx��v�F��i��ՙm��b�ـ�a�ø,� [P���Tmշf����5�M�%��3&K2ɒ̃2d� ��U.wWWE����8�W�9"'����ܾ�A�v��۷>���S�4@k�(�gٺ��K�Sy#��Ol��觋�=�{d�e}S�[vj�k�����v���(\:���&]����wc;x�cƩU8�1�|���������l$�vuB���!)Y���'�<33���Ym�� Lз'=���C(�Q |e~ A3���R�X
��}����x�Ss!��1{�=|z���p{\9����c������*�����Oj;�C���!�_.��`�A��Ώ ���AZe
i=D^���h���YƆTƙ©A�Y�źl��[8�L-��|V=k��o:�\�s/ A� ���TK��y�ɒH��.כ7��[9靼Z�bL�&�Q�+�g�3�Ign=y>�,��;І�����+cg��rˣ��s&K!c����;�>��_<�	�M��_�������ŮS�AM��'��^"��� �t���I	^���	m�<����Q�M��i��]R؄�6�fZ�ɢ�+��]��C�����`���,F�kA ���ӊ�w����r���豸�z������$=h�j!�P�	�I���ND�]�z�������F=߫�_��5��kW��~ʗ�O]���H��2��=z2Sݝt�r���,��W]qԮ�㲺뎑3�,�K�9�(�YW��Wٓ��xI�-�-�D[�4FSｏ]����)�쇆( �
�Ñw�-3�(8���<c�%r���oks���&�M��n�F21�I$�̱1sl�����e� o���!m5�6{���ne�C��	����1]�g5�����ޙ��"���$1��(��L�n�	��5>���㞓�ϓ�d�-��8 ��ǩ���=>Nr��K�+�Q�LB�d����ϒ��M�Z�&�hM�qu��Z�fغ�Lc�;��c�XDb��VC@��"����S�2�3��V�l�1w�a�!p �,D�V�y��
�&"̂3h8#.D�1�.���/T�^���[&�oogA������e�;1h9oO�++'��g��!��I��Ik�m�vtX�'.��R]4�:$$��ku>�I��*^M���b״�7�|k��/ޒ���i��$j�yQ��a;�*�͙��c�`Q+m��c���Z~#�u�8��\u+���W]qش3G�k�I��;"{�fY����!L�Y�q�S���y��2*�G�;�6�l\aJ��[n�L���؍�v4e;J��{����?�q�R�[vܹ����o1�Z��Ac�;Q�
�$h�kg�lb1N,�*���y��v�{��af��;��0E��p�M&v��#�m�!�B�Ht�%�;�B����{�c]X�69�3�`��b�&�&��+�s���=�-����!Rv�MTU��}'�9��F[�v~9�7�Ժ�����jg�,H�"�;�3d���l�9�!lS���Kad'�W�Gt���?ʰW��!�I���"n�[s!�#�p�"B �K�!�W��&��`�%� \�@�&ݨ�01UN*26�fW_[���텛����	�%�n�ȪwE��J��G#x��{T_s{֨�"�fn� �i�Uw�}'�9��E���#��A^HB�m]\y���9m��`�����q~=�2�t�2���{��WN�_T4e����8�b�ɝ]u�d����:Mό��/�r��p�2�7R�*�X����o�}�ola��{�����9����G%9`m	7���0 ��X��y���Yet;�5�OS�������Mr�qv%nd��B��!�÷k���"�h�Hp����#9�GX���	�5{{Ͻ�����X�sz�U
�T�L(.�_ۘ΅�CÄ��*�ciڐ��$��VAL��1j�3v2)��@X-���{�}'ޜ��G�b��N $����hl�O�!`�>��|��R��|B�X�̱���;�+��W�w�O�漡�ho���w�9ܞd��;�c��p�Z:��.�;���7L�_S�Y`zU1�m��0@B��m�}��}��;�pO6�$��NF`���P"�ݎ�O�%J���w���=��ߕp��yfrk�YT;:^�Wlޢ�Lv��R��;�vO�9��֩������hN�@!T��i���|��P9�<�ܩ��o+'%-�ͫxBN~_��d����:~���տg�쳤S���{$��<s���s�k��0@Ծ��
Vʆ\ ��.�M�/FQ���� ��w�	+�kE��:�ֽ��B:k���Ջ+����od�#2d��%�!ө�va�cN��O��ܼ<N���Q*P����u;�{�S�ܳ���]u��ݔ����X��o��H ��5Ů����VP��d���u�WB�!@�����0�\ɤ9�6����1�\�onMtb<�6	v�eƣRP`�C8�[����d�����{�'�E6qb�JKB�lڥ��6�1L�5aU��>y=~~� �σ��2�r*�:jp���������y�����&8 �dbpA�M�
@{B��m�)��3�����<B ��G�q��}���^�S�pA�H�p�EQSA%�[R�8��ύ6�"���y2�s̆r���WR%�k5�"nON-�Ί�%�p[hb�2����D��Aṟ��S�|��A�mB��U.��}xg��z�ׯ�z-On�>\�JgGo�d�{|�y�V�Fww:~ثQ���ϧר�}X�_�weD>�Na�ѱ/M��_{��8�����\!n�70؅i�g����^�U�&��F�~~=��;-�52��$ t:��0��jCn&��Ͻ�����^p���v��N'�����~�x O�����CH=��X��Rǚ�x�(����gm"�o2���Z��к���j{x��5�z1S�'���y�j��u�����[{қ�U��^���?'^9'U�\u]u�a]u�cw'��|�������-On��䒸:Ȁ��6��O3E�8��xcI�|QD$�#��9�8�d9	��S26��A�ɋ�l�>�y���6BT��"����e�Wj�x�Uk�;@�#�0��j�a$����n=ϕ���'��X�c ��Q�u����c�HD�ru�QH��,h�1��}�c��ۛa�!BdכK��_�g�y���Jg��P�C$/���&��~�v��S�iE��[�Ͼ��`�p�;J�1��iw�qnK�ۭ���4]b�������M�k��s�jԛ�U�y̼��{�q�k�߃�G<0�@R!؈��Ce&�-L�bR�ER���F������mL��2@ֺ��a��쬞�	,�-Ϯ��I�O�Q��{������'��(�A���$ÈD��vv4�����R�|j�
z�˘�o�g���[������A}�čKs���x��+�V:��콰?^�?=�V���{��M}B��s��p���̳9�����|Amć�M~�)�}��ޤRR�a�ːqa�ۋ|c��duN`A��yg!��-���+ǽ�⽻uK�z�>�
Ǭi�;޷�f�Ŀ=�rD9���1;�n��ɽ4�Z#����l9����ݥ��<S��W��k��v���͝����|=�6� s��.�ڳ�v�+�}���VE���s�e�߭!u�V<g���ux���>R�$t����U��h�_�{�L9��sj
��Ѓ�h*YV[��_5p�N^�����6�篕|o��j�ݞ]�"��y@1�1�'�swW��J�v�z�4��i���NŬ�毹o���,>��tX��5��|��p�J��ݫ/R�a��ϝ�
�r��!��ݹ�{���t�a�ys�[;���p��C�qf�0Eݢ^�V�H�̵,��(��	�T��a�kx��%za��G嬛/I7={8�l�y�&4l��u4l�I���hT�N��Q�$g�!a�h(�uc��yខ�(A��yUڧ�Ӈ�Z��QaDĶ;|j8�7$����0?O#������:|��h�f�<t�A7>xX�4�x�;��3���I	���<�����6��aFG

�l��QVEF��d����r}=x�Zֵ�MkZƵ�u�c2};�u�;w��C�d%�\���l���$��_Xǧ���:ֵ�k�Zֱ�k]kǌx��oKU��#O^��W8�󓝳�9�>>�u�o���׎��kZ�ֵ�kZ�Z�1���e)'�R{!���"�������c�Z��Ƽq�kZֽ��u�kZ�1�x��l��Or˺\i�Q!Z��*x�I��1:���+�TdTUj�)X{�EEA���D�*
�K�V$��9��fQb�R� ,ic��e!�1Ʊg�5_2�����"�S�*`��4�T-b����p5b�uf�,��EU�i���E��\�Mʕ��i�f��pCt���>əV��?�d�Ie��X�؝{����۽悾���zN0����E��oA���&�Cny;�� ���
cT������v�ݮgt[̸K, :�A����Z`��h4be���g���%27kw2S��-���oxlb�VOO��n��{\A�wvH�b��'�0���I���}I�	��^�}��5M5�.&k)s���\��X�S�u]��B�5�B�p	q�Y;c����wb-2UKo�j8On����k���t��W^˖ykdt��@�R|�IqDA&�<�s�6Z	����6Q$}p�]~����V�p�1��D �l AZ�t
eTj_-�4���AD���k��2�L��$�3)��鋘ƧWr:-{+'���D.�9�����!UL��So��޾���r���AUK��j8On���E�2�S�k�r��x���T��@���jz�i�7�)o���[v)�~���{���|X�.�;5
�3���*��b������ ��;����2d�K,�d�fM�`�?��k5˟ު.,���������'I������^���;�sBb��$�A2��Jk�������F[a�
TJT(,������bi�7^3DnW��Y���f&��+�s�>s��z�E�b�v��JNwoãWed������y-9�؋"�*�R7S��S�t~p�0GiA�:����h���lxg �c�L�5F�8פ�n�r�t��ԓ�k8Ty�Q
�Xw-���y��fJrٴ�7���*o����U��G-��}��w�d"(�t.ݜi2�N֛���y;������ ��ʙ  �&�ܳ����j쬞�x�d�m��^��Q�	\��lr��S�.C�p��u'$U_���#55�;���^�=���L�jNvӖYd	�;�}b󹎞�-CA�zL�.j\�W=�C�p��^��
|�V4�`���}�߯���tѐ�f����/*E5��QS(T�TL.�<�;u�k�M)��w��gF� ��,V1f�����xX�G7i�yU��\�V;K�]���<��p�RYe�3&K0��M%��u�t��zn3u룊yg�9��n/F�:�ayV����\룎zB�$���aT��A�f���·�9h�fЗhrf��&2���t{jKW��>�ۭ
��v��&Msؤ����s��_vŴ�����c��&�{5�1�Τƙ�旘�����S��hU�GWntɵ;�X���9�[��ᚵ��<�G��>���b3�sd/2�/h%�}���ݸ��<��+�ś.�W+�����Q���p�i2leE�ER�tg�o=��K:���2���Oed�𓅨�`�,p>+#�tUK�!�I'H�Lt�F ��v|b��q�;��z��I�n��b;lc>� �,�s��Aܻ��fذp���/؋c�8F���ȑ7Uo�}ݏ��̡K$C�ܚ��ׅ�x�~���;�D��v��h��yǼ��:����W>��{+'��'�QD�h�}T@qHOn�z��<`��������.��U��~���~�H�X��68Ɣ:����Ƶ�K��9.�Cä��6���F����E�+��hsVޫ�5�3۾-���VB'$y�^]"���O|Q�X�����ض��	��0� {{���~BD�պ�W,��8��힣;>!��} �]Gj�x]����6�M������Q�5aE!��%���k��쮺��;"}ξX�L���꽏��|͞n�L��3Yp�]�u�A��!�j��:F1�uӄ�[G7��&K]�xuo�{�}(��^����c�,d�! A�w$�ZA�d����A����_̈́�b$����0����Ղ�.e�R�nh ��4����$bmʯ=n����x�7"�0屐Uwq��j4(�d�y��"�P,��5H#�*�Ú"_��y̃���lp��|͞g��H@�(&"eñ�Bͧ�Uz6G�Ԡ��9V0J���_}�쿾d����zf-`㶠E��ׅ�"0��C��'�X�*�v�&@�@����Wn�=n��^����pAFS{͹�֌("}�1��dGt�}��ԭl�{M�G�S�3�Ђ�%5�޶d�Zgz���xϨ�n��b� g$� �%H5>l��� �;��$����n�,e�bl�"��eU��b�I�xߥJ�uS����'��eǽwsv��٩���"=�]��.B�@�����,�}� k���3n.���5<�V2�1�2R&L��1U[������>g�>2C��J΅H�H�/M�Z�e����-T�yz8d�VOOp��!lIF���:�^	�j ~���,��>
T%�R2uI�s肠>G���z��>�=���x[	b��R΅2	:<:��a�h6|��0�^W�^�Ľ�ղ���?|���]��kF����T��,���)���X��j����?�Σ��/�f$�JAt�����vFn�Q�,s��+��|�iAY;*/Q%�W�Z�����t^=����sm���-��i9^�����I,h��@#uiD(��i��D�gE�\���@�A!,P���X�
L�g�q��vX�=Yz�c'(�����<vS�dH;mQ��U�4.��y���'={9]�$�}�f �lb�Q�y��;�3vxrd���E��%Kqz}wԮ�<q���~͸2m��nŵ	�NW_cczc"rz��Z�:A���������3&JK,���0�O���1�����$3��7q�T4�����Vb�lz�t�WL�5v��ˇ4}1����J_G�Kx��N�YZK)|���/靠��涆M+�s�٢3Ff�u��t&��~��M�*�h�z&��G���n塚�}����2�M��i9��I��jy�����)��Z}ٷѣ�2�g���*I�5��K[��C�Ϟˇk��Z�Y̡$���73��.��nR鼮���-h]s]��6>��݁�O�A��k�c&T�ע�Gu����r���K_&�b�^�$�,]���-v�]X���=���W����[��]��	L�L��i�w�O�.���V�j���;�fm�+gdw�wp�P�-�c�O�:�5eE����uf�>�v�KL}te�Vv����ٶ�o&3ˣ������T�C�'=����B��պ�\���b�RLM��^�ճ�Ը��R.~��RYe%�RYe����f�n��<�k�]n�]��gfjR?՝�N�GWLR���b�^��ҥ�N��[mc-N:��v�:9��Yx��k�)�a�o,H�e���af�*���n����k+�;�ആ���'8&+��ǀ2��fЕ�%V*:F]�4U�6�=l=@q���U�>�C�K�f��o3���[)T�Re"83�E�Ԧ�P��S$X�����I?�fݯE�t�p��Ќ�DB� {�CD`$B(�1�v�Z�^�����Ш�p1���}��J��M��lXM^����d�GϬ��t<��$�5���y���4b'�:�o��g��Z2�U���^��Y0��?�0v���=zo�ע�g��S&�.��|���TD
�m�x�b��'#)�5��IH�v-��"���3�{Y�=�+�w��,Z�4�㭕6Im;s�']kF7��P]j�5�h<�����}�����Ζ�uZ�uͳk�<
iR������ӿxO>�����4����+}u�<�6u���BQ�׶)�\
��D��	�{C��OKٿ��^��m��~��{qy5�!��j��P�6+f2�e���\>GÁ�&'Xsƅ��v}),���,�,������16�^8{s-}��߯���2��i��F�{�TZd�\3��I"��� �q�I(��Uq4{��{���v�{6�w��.3��UI���|+�oq̏���F�y�k!�37��o]n�;<�C@n)�A���s�N��^G�;?�t�3�y��M:�������!�R�WC�뵱yQ��C��4E*ʗ}>���E��^e����{O��@�3�����5��z,�/Z��C���<:O#�j]7
b+�gk��Wq|��R�6|����&�a�g�ŭWJesZ;(�?�}>-�ol��G�g]��)�0���e0����B^���$��l(k\������O�p��v�uL�ڷ8����s�J�x�t��{V/ǅ��q"������P�����m�
i]�A8���#x�R((�xu��T�}��l�����}7,�2d�X�L�3�:/+�}�Z輨����v��@K�Hƻ�Ī�}�>���`5�&������;�+�w�y�N���0y�Ej~����}��9�K�m�쳽쭓w��Nz���@��VoL�>�����4�U��V��-,�K�UG�̲�?eĨ���� �R�V��!wϐ��Ќ�6Vhm��k�%ے4;��[�t��!�H���)bC%��g��\�GKy5s����X�C�@I�&��*��5W��{¹9v�eh61�^E�u��������������b،�U�URn�;��R*[:���q�Wk�M��{�7��{�+��ݞU�6	"^��%Ūjh�.��I!6H��W���/1ۚ��y�Nf容ʎM�@�� j�T䔞R�=�"�A���l���C�=�������+gl���<'�M��!�\�͉�f��O�NJ���A�&L坝�dɓ8M��薖)��	�m���66e��p�̃,������|��u����&�7��U{�j�"Ď,�N��l훠������Sef�b�~���ѥ��f3�%�4\���w3I�Y�T4��;7���yG[̴� z+��𽮭��{B��ֺO�;�W����X�,��0)2R�"��/�]��y���-��Ng�׮r����ݖBgD�Y���4�.
I�R5��$��ihXOH�rI��y��^�]{�v-�I���4�	P��EQ��"��f�S�;L<ԅ��f���n�*�M�
��RvF�ӷ�-��"��2�@=�iAC���Ě�e������8e�Ī�l���5�2�we�n��W�kft9��qM�T��;4���9��\���4D��Jl�.v�c=U�������i�+ g׻5�cX�of�wc`��Juu��;�W<�{D��Y�$[�G�	��i�ьyoT"�����־��ej��+{��m�o3`DW94V����z<��8*�8����V�P�Ǟ�y�7�Y���pi{f�9�M�f���/����W�=x��O;<���2��Z��&�{�W��hŶZ{��	���bm�����U���"��=�|J\A<�rv�g�0s�4��yvn�_gnN����Ƃ�����"y���2�����&Q�Q
\=t_v#2�`zP~O���t� ����9t�^�d{�篱n��ۼ���{݌����Xx����/ÐG(�B��{���&�v)Y�o��jWH����hrvwN��{'7���hvU��A8��=��$N�_{Q�Ixw��l^ҽ��{���Յ���g��s�ǣ�瘏��|Vi6���4���{;��v�gg�s�l�Cܼ�Y˂ё��M��y����1
0$>t��da���-ix���/
�08`�}�H�^U����Wh��\�?N�Q���Q2f���9j`�z�ݱ�9�e���皣�J��0<s�!��(y"XH�T�6�֑@���e Xpc��r���(w��Ҝ3ݭ�� @W?H���4L�%n$�׍a��@|�V�|ö}1`k6}��!�)gދ�q\�T`//b�Hh㲧.V�=b[o{z��@�� �rZf:�١t+Ⱦ�e�����VR^f�y�m۵v�н�K��;V��U��i�|
��T��X���X0=t�����r7[�!L�6[����Ķ��a-�cƳ������m�]��b�Β�ֵ�AՍ:���Ƕyݛ�b�率����ю�/SM����S�V��P���[fW��k���o���s�y���(�h�f;�{�i���
Ԋm&8���1g�]��"�s�٩���Ǐ��x�Zֵ�{kZ�Zֵ�SSSS�ÌTE"È^�@1�e4�S��b0Y������ֶ̧����������kZֵ�mk]kZֱ�c3�ܲr�.�K��EX,ձA`��g�b['%[l�����=�x�����ֵ�k�Z�Zֵ�cǏ^��>��E3�a�P�¾�B,U�Z��Z�W���{9579>}x��׊ֵ�k^�ֵֺ�d�����p8�Y�0���Ɖ|��X(K�~����VUM��"NBj�mAA�b��Q1�aY�6��-���d5��1a���XV����Ũ���Z
��Ot���g��WVT�<h����ɑU�Q&�!��m���n�QV(1lX�������g-��U��3k�E�
ȶ�2�k�5�n�c`fQm���rfkeҗ-����	���=�x�
C�邍e�,w�$&�{k2������W.�Y��uѶ���5�i,r��&r���UY�V������]��)]2����%n�S����-�i��ڼ\fЦM�+GucN�Wb6|Ol��J��8Į�[p�����I��\���]�f"�TL��0��j]�����s8n��ݛ{#�'LL-�YНu�mɥ"U�Ӟ<�ʪy2�p-�@`K�Y����l�R�0R��\u����dw;ưu1ۢ �X�J;�36a����=��xa�cl^�F{ɰg+i�Z2�������.���df�5��(-<��n����}�rwcMåg8%�)��z�=U��<�`�ã*:0��cP�t���L��P�E��n������X�[���dՄ>7v�z)\�t� ,͈1u��[\���n��N�r����cd��.�ǲ�+�F���H�)6�����6��¦΅-�v���GA�[�<��OZ�#�%��q��ÖK�GF �4��-��0��.�pc^[����g�1h�A�|]V3R���Vj���-Ic��SS��=:��Y[����g��u�r�:M�C�l��j�쵓\�.�^�${��e��	�)�
���a�s�"aW�Ѵ��wk%��5����c
��I������B�YYKN[Y�n���δ�R��$J���'2�IL�c�3��]sp�=g�u��UUUUUUU���\�ma���b˴���ąŶi�5�}t���.�㓚��^��Gs�e�+֝kMq�7���vK1�2RYe�̏<�;=��=hX�m�3h:�E̬����(Ĝ� ��y�y���!�˵�m��g�h�DD^y�㇑7R0A����fKF9���$2 ;;3��u��6˱Q� ��Y�R�=e8���gQ�{8ő�]�,��;�
8�q�q���Mv�5jm�}na�u�����}����d�.2s̥�d���ە��䊷C�q	���&���6J2��Y
TݾVǗ\����k�S7۲}33.�œa�Ԉ�A�j���dx]���&��x2���z�g�u[/6[��e�x�HƐ5/5���Yy�v�N<��YP)�z=��(��;���^S׋?K]|.m�M�d���Z�	�FHm���ʯj��������b�3�s�j�oksKpz�cf;&���,��
�ڑr
�h������}Y����2�K"��煕n���������*�K�J���c-}�������s^ix.�/�r�Z����+VWR���=�皓�$�K��>A��[������]�Ͻ���ڦz��U��]V��+p�dG}��kZ3KY�|S՗v��59zz]�X'�`��C�=��ˊ�)�lm>c���|��!}}Fqtf�v�c�E����Ɍ�M��+�b��Գ��2RYe�̙(
�%_�����o��/�W^�n7�y��RsF<A$���0�keIU!@]��d��e���^��l��pv���.˕�S�K�HEB���16���V�ŃmV/A�z�����e���-��}�;�M�-�ۮ*%�'X�4�a���U��Ae��L5ڿS�du�������E�'��u[q�k<9�a8Ss��7 y>��O�[�x93lc�.ӤRi�]�su����g�I'�]��h�=�����k{8Tl�lr�����V�y��{�T;8�Kż\\�l �ܽG��疓 ��|��g����z��5�f@Bf�F�jq�] <� �{�O&���	���$�ס�U9J3O7���Jmǖ.�?�݂G���Z���{�Ϭ]�Vu�گ^2�-=C�*��O���fL�c2d��%&\�^��=]G�V�|5�z�[o!�����3�$�r��Is�3�)�{6:��ikgS5�~�"�9҉��c_��4`3Ӗ"�LxO�_�u�Pv ���;yt�yO^p;���X���U *-���X�͇2�@,�1Ě�3N:�C�^~��ܴ�!\���%��	���+q��iB���g �o�{��χ<�9��]�����>�Q��op��T��<x�k�����=��g���I8��(�����_Y��Y}�͎,�"E�5�k:W�y�,�EW�������d! �I��y&Juϥ�x�5=�}���?u� �H<��z��%[���S��wͼ��>>�y�`v�t�ɩ&��o~�������ꤹ2?�r����a۹�Ӑ��5��G�8s+��/m�tN�{7���=ṽ)���u�u�LL_ӳ�Ie��Yg�1��9ִZ>|�[�ynŰ���w�����<�5����_'ױʸQ�L)��!vƒ������v�	�<�$g��_����LL�Y��4L���f��@�vŭ��l2���>�F1�5���e���I��q�yO<��l�����I&�u�c�K�-R��[<�����[M[L�1�ރ��z�xy�� ع��v�;��*�9n�]")2d��x��3�p*�סc� :�mVu�ٮ��]�L���^K�l�-l�&�#Ӎ>Ե��뉔�Vv�?�q磺C�����*�5T5Rfy��5W����&�m�?������={M-�X�S�;�����9'���>NR���S�����=�w=ћ��vV����.�K��d������X"kWdv���@@�-�p�H<Ւ ��)՜�o*��N�����WG7u�w"O^ݰ���s88�i?N�,�fL�K,���1mg1%Q,u�j٦�Ri[��hN�N�6H��������"��;]j	wW!�u���;��ϛX�sJl���Ѳ h0�WlU�F��gqպ�l����b��OM7\<�m����l�l;7@bZ���۩���N�VϬM�-Fi����������G����0�p�KBn aQ��CKL��\��^g��Wp������U����"�4 �6���I9r*�$�WAad(ǉ^�W��s�=m=|��2�c$�'�@�5mf�eU�X��T�>z�{�����^�o-��;� �:5Q�*��e�Pf�	,*����ۮ��z�&�6��/x�{Ulŵ��H�"����g`i
�4���:]��l����lfE���;�ئ�5�n�C^Z��C�5��ͥl���?{�%ņ�dB��N g�<�]�6�q��Ax!?>6�6�D�M2����S��W��7p�{�,�w�f�&�mv� ӹ���G��h�	�q�q���71���ǂ�����F����޹Ĺ^�����Mɇ��t�p�f3a�$Qj���Iht����2dɿ;; ɓ&pA{���������}���.`$��B�@����>�O�?������C���#"�~׼�.�����;K]�ob���7]�ק�כ�F� g����VF�)�Y��d�EI�-�S[�o&ȹ���CQ�M,k��}��}m�X�on����G[�>�l����bm
lm�v�٢D������}y��A"�Y�eޛ5\ӭaϓ��f5��k6�u����]J��dH���7g���Ó��s�K[8�ȕ>>���|�zy�$�W��iB���Ļ*j�aR��:H�����A��!;�.}���Y���BY.�x�Ӟ��IT�Qd�K(�)��كz�v�&�Zr�J���{�
����E��v�����O9ċ�����!/��6��=�+޻�ݷ�W4������2dɜ���Ŷ��g�e��]���	����ZTD6K����!w��f��8�̿=,���d�N�w@ �`�z^1�!�˲��鉤�1DϽ��ւ��O������=���gkgp"fg�o����?'������<n�lI�{�~|l͗pu�G]�3M6�ͦ4e��8���G(�g�Ȍ�S{�/{u����w���C�h�S)�I&Y��2-�7��J��X���4��Qq+wc;&_%��t�3�����|�Ke[m���כ�߮��SV߱��kf`R�]��^{���^����d��f�v�k:�������=��`8�7�p��\tv "�G�-��rv��������gm��K�����i��ƶ�� L�h�����i���XN��+�F����x���v�9�UCUؗ7���:o�wɎ����V@���s����̡����e�.3����{#��\[oN����~����w���Nk�+��D]I����j��"�Vk)K̅�|q�����\�mҝ�s�<�܀��� P���J�,�b�iR,Y`�I6��c$	�(c�X*�"��<B�dP�m�1�7�����ܳ�%�̙,�Yf#C��o���CUO5<ۂծ3�p3�����3r��}��1�!��MT��=������1|*���K�2��޴jێ�<����!I���tm�oLGX�hX�6ҍ�nek3�{<�������L�&.�;�GY��=U�j=�3:��j��p�LΐKK
-���9�7ύ��/"n�|^��9_�Z�zJf
��&*�2�U�i��v�$PX�iMT}��c��S��f�<���r�y��MU���#]y�H����m�Qy��=��X��ŋs{���cki����p�p"�nd�Rlj�D�*�r�ö`�@���/{U�W��4��Bg(���f��{�.��4!Q3G."K��Ӻ?��<����z9<�yƽdf����	e��u��6��e0���X�'m�;|c;��e��[-�2�99������d������]�� �Lӹm����|���&JK,��%��ǝ��F�7�M�s�D��\�h�sV|]�zQܧguև"c���s���M4\�[�K�42�����j�ug���a�<7
��k�6�f�|�u��T�U\k�r�MAe��2��6j7N��v�ݞ�a�=jx9�Wk��W6lh�GiS5�#5\�����?VbW\�b��-))��f�:���b��7	�ɤ�I�<9�g!6����<��F�S�O?p�S�DM�.���!j�@ɯ2� �N�6b���}t����λ��OY��7�����3�[K����7h�@�qoKf]�55��q��������r9X���(���L.�.� �lK�;�uH~E���ɉi��z{cٔ��|6�b�w,�лi��@Q�v7.:9�[D���Nwfө��>�v�����l��H�/HzU� �Daf��"�;���$i�e@Í^U�Ɩ��Heb��R�C8�>��?~�Iz'{'3�Wj���/j�c����C���^��l���-�����a�E<�i+��$��?l^���o�,>�O�ڡ����{���{�ʘ�e�bۼ�c��@�O�X�7L��As5���2o�;; ɓ&H���l������y����A$�m���`#�]u��
�4#�	 sx���8�{2������u>�۶��,s�� R��D$�uKZ|�o֧�X�R@$�L<�476E��o(����+�n�k�@,Z�R��-�RzV��ȻB����U�������ۧ��~� T�:j��WP/�����8/	�z��Z�wl�K�h�X�5����L�m���ј>O>���d�K�nb���]FϬ��qئf)��x��F6��i؜ ��C<��e�9Uakʘ��q�Tڪ��wj�����}p�4�j�|�=�}�@H ��e�3UX�*���*w<��Z�)��z�n-��/���wr�'�r�L�7е˟{.q�N��6s�Ù^j�\��W�y̾˻�fB��~�
�~z�{�o�彜7:q�z��:s�vG����7����;S�ݞ���ۻ�ۓ�	�C�����u�n��`�˓c�d��^�<k����(��j�c׬=<6���N��'�G�ۆ���ξɾV�x��o��7��.yٴr�zwf���x�-0w�^���=sҩ��w}���]�oМM�$w���H]��׶�rM�%K=�n�k��<sH>�ԺPy_��=�g��>CS^Oo�
��4�r+�+�3ʷ�0�YË��Q�o�)Ύ�l����sV��M�_�;��M���T0��\,�9vO9D[Ð��u��麺�x7{t�y����C}wC��zj�{���wꤍM���{:�s����#ݦ�&?����0/_��<'�7c�W��l���&�����J�|4w����
�sr��ψZ�x\�MB�>���I�\����g��1��ǉgZ��]��'����s�Lm���6�.���`~7�t�خ];��`����j�'������ydFCI�<HzɃ�혭IX�0��S�E'ʒ�x�:��i��)�&1v����ηv�w˽CLSićXvmT̲z������@�ֶr�ѹ_�),&����n[��n���=�
���q����v���I|eͪ���쨑v�ܘ��X�'=׺�����LnX�ݷ*(�j�ڵ)�fx�L��%�Wu�{����iweAު�[�8�o[���䷹�����}x��Zֵ�k_�ֵ�cǭ�ڒߖ�;���R�4E[h���2��X�S_ N�L�l�+_T��l�������!R+�2յiig��ɩ���}<��+Zֵ�k�Z�Zֵ�c���+�ByJ	�_,�¨�[�\����Ŏ�kKk�r�U���LqE�CYUE�fD��y�33��9�r��u�M}}}x��Zֵ�k_�ֵ�c�z���N���{tn����մ��S����8��O���zu����x�ֵ�kZ�ֵָ�c�={���YlET���L������Lʳ�f��15n�n���\`��<�b��4.��\���(u�Vy.01YXZs$�3z�Z��UG(Vf�E=sS��\�2ǣ�1P�5aP�ƶcKet��1
��2��YR�SK(#�
�/u`g��L� �i��˓X��F�
y e(��ȳ�2�֭�m%�e��ܸ��j.ڮ%���w)�]�W鹩Ie��d�@��g,f��c�r��߂X�e[XH2mY8p����Iy��ʍ{mdM56L��u�˨�����綋�[o[���<��4K&�L@4�N��u�^Z2|췴�V��+k<������9�Q�����Y��3�%��B|xW�;�Ya3-�>_��W]G�kq(;q,�1�U�aX;a�D��jSw�}w�}޺����eR�uO���y���7�c=d-MM`����&�6f;^���t=J%�y	�̾�Q��=��c-�zfH�[>��Ma��K�� v3/0=���5�oǶV^_9�4���Nzn�"�Y��p��\
�v��ږ.�N��
0�{f�k�^E5oCv/K�ޞ�S9;m���mt�����m�շX�#H�h~����p��>�]1���J��T e�:@Y�H&�w����@������(K,��%��5��|��@��ƨ����~(&�g�Q��}��������
����%$�@�����w�Wp���f��-ܹ�H�&�W�Fc�ϟ|�M�Ă���P��G�_����"+k<���$�۬K�x_�h|��d"���Ա��<�f)�t� �T�q�>�Q9<�m��`�]�-sY�v���ls�� w[co5����r�������Gu�����hUdC�J�n�|y���Tv@r��Xѧ�ם��[Y��|2"�f7�R-'^�!Я+jL�J*��IF��N���"#ٽQ��o'����k�gv�r��^�Cg"�RzQ}�>�tw2Պ~�
r�/�M q��������(��Tz�..��A���E��}�ԭ>e�W�}IÕ" ��E���B� ��!1�S�e�<���1+c��:���h`���kg/T�4Gv�<J�t�@.W��?�����u�#�8�u����ϟ/W�v�m�لӃe鎷5R�]Pֱ���ė��P���6�	6�����e��ڭ���S/j�z�[1u@�����^қ���\$*hLb]jMR�\5\m��8��وAya�	n7.)��ms���B��\a��gڤ���Tq����Y�{�ɇ{�|�� �3gG�/	���f���:-%̭D<:w�6���=�A��<������۶���$���KL� �wL,�1$����F�Ͻ9r
	����C�mg�����e �sT���(=�2hcq�*��􄖙Y��yvo�꺍ӗy=�d
��T�u������5���9�����yӴ��v]캈�ۥ����rb�Mk��l,2��R�]�-73ɳ~�<�'gET���ⶳ��u�)���$���娾�?,�^��&#�g-���A�n�Y�vܤ�[@(�ciV�	��v���	�#�����6%"�WH"�����G˼�����V&��t�LG�'<��M�}PќĂn ���֦�Lk�J��oJ�AJ�H�w�X�>��^��{��E��K|,�t疳�c���}#~�z���=�b�Eb�4Ո��I�����d��?��%%�Y�����g��T�q����u�����Θ;y�����ߣ��pA�"�b"Ah��2�d)�i��9��k�jH{�c���Vs�����ɪ��MJ�����h�ɯ�Q��.q�m�Kv�nm� l��S9��%������eF�˼��憴�둛V=3���W�;��e�T�2f�@=���zDw��;�A��ڋS����>u���{��>K�(�WMS����=}�o>��5% ��̶b]�-A�%̹X�r��P�;<���ղ�IEb{L�j{����[]����wd�~ͦ���X��(Ļc�۵��_���W��!�ѳ]�7.�:;�b��m��Mfm^��e�1k� ���l�E���bD:'��c�*�(D�Ӧ���ˣ�9�.L��[���"�eS��}�>�/��ʔ'N�����|Y��L�3�vvL�&Z=>���Q�}���3�ih�d�I�p%���V{Yǒ�S<5&�n[�<bkk��g�ɖ�筜��b� ^JԅS��U��Tv��9�A�*�*4n]�p��2�Y���G��w��3�f\}����L1��K��z�\BN c]��n�BO�PB~z�1h<�j��S�՛	D{���Ƣ���k�w�����Y�5���g%^g"i���z���15���L���� ��ʳ�_�_�M������1���.�]������,��z��G��#���b)L��$�U-ٺ�Z)[㮃��OUWY9�J#�ۼ���zT�����c�?~���Fj��� ���j��Θd�1n/d����n�/�������Z�v$�������XN{�Ea)z�F�%ȗ�h�HC�4f�3/N�L�Sk&����g,��&L�� D����]�Z�S.��~T���-R��<����D�׵�gC����2�w�;^��A]�BCI"�MMi��g���Y��ҏ�w��:��n]�q�\���B�)��AP��wpTTMY)�|!sv�
�&e�"�z����GGm�à�����55�!^�A��K&݁��͕ծi����}ۜ�����,|鷭��)���GB�I2�hl��Veܧ��sV���;*�ׂӒ}�Q�"�'u�g�R8YE���[���ɮn7˼3���gd/�g	h�2"������GsI�%����څ�7�t5�{�����	�܉�6�8�=�uyLD�h�\o�'�p����m�5��f���T����:7n�v�rMv�g�t/=s���Fm{6{vKn
�_3��g�8z8��$P �A##/s�p�|�;;���Y�qFc�ԤRk����r�hs]�hB�����u&yF9���K?��%%�Y�ɒ��Î���hA��OX]�Ph1�5͌Z��c�p�mʡ�$v�n�v"��^����v�,`]��]�4+���N�؍
�<�;R:�h����:�u���1g�N㗲	m��۶��V�c�cc�ոӍ�l�C��v��nٝ3GY�NN��cAK�~����Y��:��Ir��]�Z;%��Ⲹ�6�=Q6|!��Y�1�(]�ƌoWo�E�n�c�q쩁���/��1Je�)��g4�qY-�m�_����~�yzI5�ؼZ���;<{鶦��M�-�4Y�m��+����#�֮�v��gE�v��ޗ�޷�OI ]�!J�c}Zd�,�!���� j:wwԞ��8�Λ�k�n��9Y�Л�W'�I�yi������|�3�:��2�|Z;8 �t��L�EA��qޝ��^�K;�n,v�?|���i����r@�wn�x���0g���Q��D6�_��p�b�S��T�y$�\/�y��'y>��s����I�o!w�r���Dg�J��w+Y�M�e�d4���|χ����޹��DF=��ʚ�;�ȭ5y#^�Ѓ�� L�Ie�b2RYe��k_No���~���N����r���Q�CV?z;�����m�O#m-\Y8œD�$�g�k=s
=1�eM?f,��Gv���kc�2E5ہ��AW}�8��M4��f^$�o��w�ɓ��Yَ��CM�kMv��|au�ט�^�7+���N�}W����H(
�g�*�UWX����\�1[x��|�Ͽ������k���1���M[i��3kp9�Bu*�E5p��I$����اޝf,��Q��|z�'nΠ�]�Y$��U��ј�T����,[7��ٚ������H��⼮���*Oՙl��4��,
ə��Et�>���F��!�=�����:	�މ��w��Tmسf��.�wY=� �7��d�ݛUwM?��
{3��`�~�1�awa�/��~��C�왓&A�&@9d߳=�J��{��L �4�FP%��o@X2��*k)�*�N�?�y�1e��w�uw�b�Շ�mh����6t�R@�����^��Wc�z��ik�W�*��.��}��v��z#�ހ�~ʊ痻wA��v��A��A�mN_>~�o>�&bZ�e��)���C�93ۤ�q�ڨ��:��-=S?�)���Q�꽞����1���u�@�q>4�CM�CqL�雦���;�t��zn+'��ŗ���1�3�6��;�<fM�K�%���QF�H�@t2v�6eϮ�z�;�^��Y^Þ�L��8�dԄ�etEk=�:�r��U���|���Q��׷������~a1���=²�:�P���	�\��UB��!���b�x@�o_�E!�#_	[�s~��EO@��to�=~wSq�>�F��#d�����|?��g�2d�,���,�X��Y;�x{�I�k���f �/;��qz�ӯ������Ų���gvS�^;�H'���N�	ۈ��˘�b�v����@tӇ�\�`���E]�@�ÖPB�=5suk8���Wp;"��%��9ۍ�4�������c��?-o[UȆ���-@�wN�6�k"*�����g�ݢ9�1h�&�\�w���TW���2REd��mIl.ä��� 󹞞}�F^O�� ��"�T	-2�U>Ϧ��^�8������7����t�1v�΃�a!F���-�H���CZ���]��eo����,Sם��;^����	�!T�UH`Pk۫ё:�y7rC�9f������n�9��{#]؎� �>�<5�
�I׏��ۯ�b�h�v�>>����Ua{����]��c�Ky;��|>�n�Xw��<����6���$�d^��=�!8�q|wĺ�G�(��OFwq���������4%�ri=���&w-�r�/3�G���P�S�0���f�J��m����Z� {�䱽��-�S��L��<�{?O?.���+*���oo��#+w<��;Y������k7�G=Kd{�� ���I�ã���Os����z�ױ���ճ�L�.���9Q��L�Ӻ��$�
x� w�N[�Y������J�xw���*y����bG�%3��w����P�hD;|>�g�����}�4�F���3"=<��������]��;���e����x�������p����7[8��݃QM��\��._| {w� 嵿-<v=P}��������*�0��F�o")��Z���j�*�]�*W6����`�S�;}��v�(�7��p{s�m��wRc9�����ˉ��pX�
p[���Sw�O���v��Z�m!؟��;��<�u��l%�d�~��Gɬ�����6`���`�D��c&��F��Wg$��F7�w��=A9�[���(���J>X%�jv�BX�%4aoF�G� Eۑ�T� �\(cőm���H𓠱�q`?�4&����j�� z)]ì�b�� ��������7�~W#a�"�������p ���Ia*1?\�ĳOm�=�^�E��f�F��0$חI�EF�Ӂ�V�"�L]Ucxpaj���qc��FŘ����1�!��y�N�U��u�wL����6G��������Z�xp����=�>���R6��S\��l���&�зq,��a4�C�7~y����<ib�L�:5���� s������%d-��ޢr�ic6��^�b�������H�vz%�Ѹ�
g����@o\�$�:����B����:���ٙh�kK\5rS�s��
z���c��R�����LJ͡QDa�9�\���9>�8�������x�ֵ�kZ�ֵָ�c�=OVw�0�\�V�F7`^$��F�
�
M^�A�p	f"#�t�v��>�;�5�u�<|}x�׍�kZֵ�}j��kX�1�~���sݜ�ZT�DCWV�)�%���b��d�+OsO2���n^=<��ǧ����ֵ�kZ��kZֱ�c����e�Ԝ���-�-��Ԭr��U���E�[h�c>&�MNOgg��Ǎ�kZֵ�}j��kX�2jnq�K�^P�c�2,��7a�Xc4�ޝ�
q��3�i����2��R�
Q��题�DE��\�!j�Tyv�$Y��պ��b�lX(�-�Zd�k:���i��H�T9��Rxɷ���hiS�\-J��р�VX*T�J�,�$-ZEm�ѭDeZR��ֵ�hT۴7�m��
�ƴ*�b%}h���TU�Gv��ц1��#��͞`�VdlJA(�I�a�磲iV6�nk�u͇�Ĝ����Gvˍlm�o\:��������T�Y�����dN5���]^�v�Z�㛭��*��:}�6�m�!�Js��Ξ�vu8ٮ1(�,ư�X�"��ɹv 9�}T"r5�g�*�����\j��mtKR�%�`��WP(���c�W��фN<\n���En�b��1X������T�@�6���vw8�b��5/���{Tn��u ��*�\ц��ЍP�l����*��]e�7\�-�"
�:K�f�ma�1,M���Y�B�K]�5��Y��	�e.�����R��skkR*�m7,���I��C�����Ntg/=w^��`ƫ��g�Gq�Q9��������8��p݈;=q'>�q��n���ڲl��63�����=vKY��׊�y}����wj^�{WgQ�v�$P�Ѝ4�ΖP�d�0��]7sQ�]�:�WtVy����ѰX11�t�b�!���������X��E5�?pd��N{on�7Zj�NR�ɺnNv;p��mT0]�W�;LEறf�r{=���(ʭRNޅKw^i�u[j��0uS��j���(�h&�sG�B˪�$�e�8f����j#e�����Q����ϲ Sb-˞ۊ�al��)M��Q˩�@��� r-Ķ��Z�3*�&ٳ�Irj���Z���Me��k����fqA�����y]�l^'��u(������yg��y^�����;�p��3&JB�(b��o�E�S[tf/.���'�mխ�����6�.�(\ci�,M ��2<���[�N���aE�	y�q�ԍ-���.��N�:�mWn7=ckg��6�2쥨#�j�h����<<�msO>�=u��ٖ#"������yd7+h��Uu��Ȣ���,r�[a�����UѢ�.&�ܺpH ��,t�T�&1V�R���[�%���%�]�sc[�b�*f��}�Y>���{����E�P�S2�*ZB�|��{��Z ���X�f������1v��V�k3��NNS���12��^�lcqU�H4϶}\P�r��ksu���u���t�-/|�ZH>m���4�m�؞��+�Ze�ڍ�v�egTw6�(-ф?BDzm��������m��LYL�*޾Μ5	k����5���b��
jd6Vs��6;'�W�=~���
i9	�A���տ>K;]�+Jjۋk�j�1��D��"��M̂-|��ϻ�9�"��y_l�{�j�=wC<�7t�! -��)BY.��P���'�fa~S���H�_Sķ���Z��X׿V=�~��j�ߙwj
7T�P�X io�.X��&-�@LC,�̋q�,�K��\�?Gm�U�Q��CT������G�ޖ�e�����w�"<�x]��UŽz��u��땓����oB{��U-k���c+�ͭBq�lz�3�=��s�lW^�+�J��%�*^;<��r����W���׬��ʿTs�aj�*�Bk}\My�-�Ju2!Ġ�����r��(9e���T�!6�،ѱ*3A�-�H�-^��d߃�~�dy�,��2���f.��z��oy5�l�3��qlp>��C�h����ga�,�9�ٮ��W�a	-�Eyw�E0�lmj�AȺ\�ʪ��h�Ů6����(\�����&\����G0��B��|e��o�ѹ1���آ�ѨA��5�e�=��[��y�:���# Čee�V��}��z�*���EO�cD�۰s�I%��\n�/��� �&cn.���f.��LF'g<^�6��`ƨ{�ăm�,m!3QX��4�w.�1�#&��y��Z���
h�,�f�W<T}0�E���li(��Mw>v��o��故�.�]B;����au��\�G8"a7���/�����<�����ǚhN[�\�.��� �Ɣ�����tC�� ZWX$�fH�BZ���X/E�h�g��.��uf?n�&���f ��e<�=[��:���x�hPr��J	��,�^Ɔ!���^c�ڻ�5���]�um�پ��WM¤�����̖��F�^�1�\Ňw��Y��o������1�$C{3b'����}�s@�9�pa�E�Ow�=���_bڻ�{�7�'J�q;���:�[�6��$ ��� [Į�#�Bđ�*����_`hT*��I���V����d�/Deg9�:��gp�Ly��&�&w��'Т$Wߣ^�0|�#"��Zc8@d"gXO^�}�>�66^]�XkW`��	��vx�2\m% ��6 F�h ��4��BW��[��7ճ��Q��O��_�=黙��.�6���0"�]�lk��ou��̺����*�����~���2gj0˫m��]��ͽ�ζ'g=�v=W���,L3���[�$Psស/�C&��=Odn���7ճ��t�a�s��X��-�oR5���Ҷ�qY�Q郗w\��;�����N{2��u�����&pi8�s�9�q����;�|?G�fd���r`d���!�^�:��/�v��ʧ��⟗� �	9�����0�2�)3�3� �D�m��� |��w��e�]�$��w��5�"?I$�FF�$Dr6���G;�mw�8v�]�Z����Čg�BČed�9yl���n�sxiq5%]d�fU,�a,���	��� �66%�����e�fx:{q�ӳt �j����Y�uk���Αf�8�]�M�!�Bh��g'`M���x��%���֢�4srMy��X�t&.���dm�У�`�nخ�Z1707��T5�}��?_=v{C�:Úxy�+���Y���o����쟱'��9ޮ�]^9��^?n�y���q$�-pK#�p+���3,��}7[�z�1��!����R��?fp��}[<��L��L���&��z�+MO�'�,�QG��~y�G�eļ*���˛ۮ�o-zA,e�Ї��U���I,�s�j�r�q�����Cz33\�u^?k���l���ʪs���\G77d�&�ݦ��v:C��2x�`��پ��V����Q��,�j��Q�\�Z��|Y��f�: c|������+�.����L���K�����qF�P��[|�z��4�d�.�pz��}�7�~�glÛ��}��c&]2��z}������O����3��h���¾}u���V��ZlIU��z����#r"�^1�E̹�Mx�1��-�Y1�d�&H���Ik�#=w��:���c���d+\���[M�=x���K[ �V�fYݔJ�󚠢��<.���V�k�T��H(KQL*�M5�{�p��j�m  ��3x=o�}�7�}�M�ۧ}`ћ3 ��^|�y)$QM�-<�n��L����	����Q��vgً�}�s��c�C���O�ֽߒ&��,,�o�������*W*�
\<�H�����1��-p�ף��W5��*/���ɿ^ϕ��b���)�@��0�[z]�Ϛ��|O�=R�*#/T����.�ǭ�/r���8[b�=߲�j��g��QJz�L�4	!�廊W`lg;�]��C�.ڧ��D>�v�1���M�G�}�r��1�"rŪ�ʁᯱ
��'��@��'�%���K�(�Rg�՛��M��wt����G5SM&������n@��?��L��Fp|�����M�x[�<��zps[x�%%&�{��\pzv�o�4?�+����o&�zݮ�5�CFS����ɦ�Rq���	"`��5���}:�`+�imY���^㪸�����`�wd\�0z/��rIy��z�^WU�{w�e-��ˬL4�`��I�*�RUϭ���������}[=oňy��5�
�r�4���Uպ�.�Ѻ�JJrY���_ԓ/>�77.d���i"��Q�#l�O�4�AǬ��������];=Rs�R�ݮ��즖�0��S9�=�x��k�{w��X�0h^K�~��W��Py!M��U�]��w(�x�CI��;=��0�tݛw�|�KI�T$O� ��ɐ`��	I�K(�Y*@a���xgl�A�M�-�n���tg��ݥ�����l߯g���yBb����>����>���Y-�K<�DP�[�{�=��R���k�[�9�UFh�j�Z˩��eϞ[߼����K�2�q��^M��cv�
y)-�Z��p$��ж�ܘ��"�6Z������n�5:�Nz=�X�"��'�wҧq�p�e��X�8��i���|*��<|'f��y^��n��-�Os��X�2O�k�����g�Tkռox*뮼����d0�tw�y�ױΑ0Y�� �Ҭ��������������K�杸���s}���
wn�MB�[��J������U��͜�2��ǌ���,�+Y��Ҡe^���9^������3F~~{D�h|vL!�J��BK���oL�y�����z3N�������z9�V������ثhv��r��Xƨ��4kaN:�;n���H�F21!:k[qL r����`A;9������M`FΓ���m����W6���@㭭��M����:b֖�qj��I<����K����c��rF�\m^	�kxΰ����Y�˹����BJ��`���-��������r<��r2��l85��>�?�����d���=���E��A6��Ta��(f�~{��y���p���45T��!Ufގ�u�<���ס�#<��S��	4�t�ty�]�|��T�%^��ɯX��"�CI��=9g�I!PN�&S	�l���i{W�X�������k�a�N�f�bI��5S}2�ы*{eMRC-��k��xhlq[7٣���v�+�B�A��Mjo+����m"j��!�uP�U)�'�Iǃ�װ��ڏfV�Uz�:�N���+u�Yx���}�c�9�q�K��a��J���z��U�(���eea
��rS�d���D�^v�޶�5�*���X�m��3=�mY�#%%���i� �U!���Qy@����z�G(̈T��>gW�ǨNy�՗ۮ���Z���x{5N�߽��p:?ۅ-���R�Sbř��  J��3�y~�Su�\���<�UL�
�ܻ�peMr�~gR�^�A��%繫�v�36�n�^]m�sY�M2��$	�U�nP��5r.T��^m��3:6��f��^Z�Ks�yU�Mܴ��-�T�=���� �E�(o/Vo{Ʃ���c�pLD<��2���3N���^���4���5@x%7�>_�����Z�^6R9��(<7i�RgDm5
���|����+Y��Z�⽫�篳�ٕ3�z׼���<�w!�C0�A"�d���-�=2_�3����mٮ}Q������~T�����I�z���TE�cx��v�����;; �����������֮��\t*q w�y_{���$;.{�;Y�d��m���N�>�3��OI�L�+� �]��y�7��q�щ<��D�<��c���F�=����sZ_�k�%�>�#2g��vz�ԧ�7&p&�˓��H� N���?c˥���I��N���>�z��@�3x	��/����ݧ���+m�,QQ���x��n�/�1e���1�Zͧ��!��{i���܈:�y�q�f���{'-V�{��w�iR�����/-����dx�>;}R
�{���h�any��zp^�����b}��c�8���˷��{��6f��%�P�U���06�ٽ|�{9Vy���j�O��{{ݕ`�M��6l��5&`���~��{���el�y�E��s���Sh�d�n͞���^������9r��uws.��`xS�yy� ������1�ɯkA�v;���#o�p�7�P3�o��c�4��m�X��[Ҷ/-F'�l�,���pC�C-�$�Y=�4��P2�����3�k���:j����٬��sq�1������&X;��(�x�5�}3w^��={4X(|H+���O����Ł��[� F�^��1泌�H��9�]��ql�M�8{ϟ�j�<bi>���{[1$�3�څ9pf��&�������^\߳��Qkxyt���P�>8�QM8�`��ܢɉ���=�����F��kZ־�Zֵ�cǹ�}�y�#�['}�14�1&ZX�B�bT�aY4��鈋�)S�LIg�Q�59>�O�ּyֵ�kZ�Ƶ�k�57��J�~sS�w�&b
��F�/)�ҰӦq�E��%���:��=<x���Ǒ�kZֵ�lkZֱ�c���rT��\�r�Υd̥m�g�f"�R���+�7�16�\��X̚���g��Ǐ#Zֵ�kZ�ֵ�cƦ�'���}CN��[W�SǮ�f�6�U!�F,Db#R���$U�U|e�-�
����4EXW��TE:��
�+�ʩ^���W7Aed���L�Z�*��9�Qm���b:J��U4«2ؚ�J�҉�f!Y�Q�M6�(�B�i���T�S<��"k��[m��,m���PKj���kTf�&"AEbڴZ���eFnԈ���ԨZ�Ux�K��-E�(��+6��U�������u!h�d@b�X�,Y��ꩌ�͙��m���Z�5ۈ��A�a��LFd�4C�zQ|�fU{.z�9�؇ޢ%{ֱ�޻�>E J9��9�׆qT�z"=�"i�dTd^�zٙѶ�T��)-3Z]ThGȓ�?S�y�X�i��R^{��|����GN3g=��Nk��F�͜R3eZ��~��v���\9U"����u��b⳯�;��{�dW���=��y��U �	,X��ni�!�l���`6�k5aQ���wU�d��c;u�lafd���nǪ�L��3�EJ�U`�g��3��VC�flm�
��B�Yt�= ��̖ѱ�~�s�6��s�4��A�ٛ�y1qY������>���!˗�+�MZN��[=��Ϣ\�����01�����M����.��#��fM��KFn�!U�9���ŪU��G�=w�}Iɿ^>䯿k~��o?�*0��W���V+����]�
-,�C�)������꡸XIF2�E���������+;��ݶ�6��1��P�aa�����<����1^ڌ̭�����똔/!Vu���jhkQ@y�Z�D^�F�8~��ً�ξ���vi�x�p�ߨ�����2z��G�A%_�p?ߵ�켙鷧#�_�ֵ�E�3�[��
whcO6����[@cm�b*����ס���~T�л���ܶb�j�GY$��cJ��_���;f.+:�#�Ml�v�z50�,X�Q~V�x�\��:�w5كenա�N��E�^3D���Z&��|+ȉ¬��HL|�Rō�I��MLD��/��/N�������9}s�_=:��`�,�D�6`M�K%�������sg��]ʴ�;�`�q�n��1�BA���i96E��2�f����F��%����]n�Fm5Ux�5�4�&Z]IlT�Y����M�7�$�,�zv�d諍��ɂ3�5Y�`��{R��כ�<.�=+�qgu�a��j��p�F��EV��v4�ί�_]��GT�W�b�:$�d
&��~�bD�!�X�g�\ʊ��6��%��4˞�'�y�O�bPy��}��ӑ�}~�:��OO�X�$���U�^��;�</�U���l?�3�lπ�Lo��G7���A>��;y�H���gd�z��O�ׅUe�͈����n��%ݦ\>I�Gp~/��62��v�9^������=�<;=Q��Z�Ǿ��I������=rN>��IT���sP����z#יѷ�J���5�<%�Dp24n���D���TV=��7JE-���L�Y�x�CeA���]睰��?}�L��[�ۯ�ꮼ�=��}��۲-��n�� �̧W1���Zۺ���r�EeV��H��w�/s�{��y��ty�-��Q����ҽ���(��e+
=U���(��3�` �}�o��A�bIu=|��f�y�{'+�#������swhn�nM�p�/m�}!{�ȉR���]�~�us������ɉ���ŞKKr��l˶v�O�x���>�fhߘ{���LS&3cj7-��(RcE�p��^�sVom\��ܙi$�&t[*泏�.j{o�ݺ���k�<�+	5X,w!$�34�*����>7�t�I�m�윭��]����^Z��1A �5��W�L�ޝ~�8�Y�))�/z�ޛ�a���~Q>�l�t.���U�L���Gr]�Q���q�U���g��a��wbjY�L���^=Y�^vO0h�7��55w��7i��W�����QD����\{j���.j{o����ke;Zkk7s����۷��"v7Eb	��L�Qb"|������k2��5?t���8`^؜kS����E���e�T��9A�J��_%�G�.{�h�<g�_]o���#��bI5��~��c=8�e��*k<I3wL��%"�<v�*��s�w�j�q3���m�V�O�9W�t'uN,�-�$Q	+�Ğ"�
�ݞU��m�j�U�ȹ���c�"��V ��7j�z{�%݂��.Q;��\���/.�Y���l2԰+�]4���fq�SR��-�g���qeV�R��?d�t���9��I�[!xD
e4̍j����|�9�<���tEf���}��u���Z����HԠw8��[H�@�e5kS'J�5�����Yy홫㾋��m�?c��d.Ъ[���^=��ڭ�������}':�������,�k�`��`�<�쌵/~�&��=�N����Y��'����qMQ�����)%�a�)�聓/VH�� bI�_�Z�����Ѻp���d�bj��k�S!��ϐ��Mm|�Ѿ�W<Ofs�cy���7� �h��X�����%�-��'n� �ة�lWy����R���]n�XP����	��ƛj�l��\ ���~������v[vÑ�~����um�il�l>�g;o�ii�d&�R�Tݝ\n������^6.oӏ���DEL�8�L5�!��]�mc�_5ܵ�_}��̄��Տ��{�e>��w-�T��W���R'I�ݠ�����W�ɟ�lV�>�ݱq][}M�-�N!}Q�#Ɗɇt�ӭ
q���c�ӇO��Ӊۙm�����p��O8,z.og����$��:HO��#SIꘪ��NU�P��p�]+��zg����;U�R��E�G�t��h GҮ���Z�� _q��HǧnZ/�C�y��i܅1��Kp��]:T(�(	1ׇfA�<���2�0�nbk;��U맀ͬRN��gtr�;n����ţ�֔�n���H���I���㡕-�u�f���4#�����fh�@1b��*a�:4�E�x}IfK���lZ :�U,�(�q�y�2�xY��z��[��1A��`={��ٕɇɶ�\�n+�]���X�<WgT���zy�{�9t�>;=���4�Č!��p���Cj��������Ϗ�D��l��$�[Zj�.w.�KK�vգ�s|������W���y�z���#D?S�~bS;Y-�w�JD�zjj^�V)�A?)�},��V��ظ�����[�����_٤��P�o@o�I(oz�z��=�xH��ܜ}��i�5l�v��>�c��YT�#��(����f��rA'��7Բ�39�]��c��llku��
���Z�W���3#"O_˄cѬsr�-v�=׶�9��E�CE=;�j�����$"ȷj񰧿_g��$����F�Fk1n2��qq��'hl�Xy��w�)+j��E����u�7�ƶ�v|�=j�6�d41���}�R�x�<\�p�u�g��0y۰��ٴ���=�.����_�d"��������a�5�֏����o���b,p	�d��T϶���g=HeI��)��f{/��E$�0���yB���w��xyl>�����+v�)�4���L��sRq���ީ���g�A�.����OzOd�t�E�vsY�z���hg�����)�2��3���jH����3	��v���^s��oI���ZZ:c����<���|w�N��i���mt��z���l�Yk33�r[�\��C����X��� �9�T�%�wec�>��m�dt��K�HsEJg��0���RM�a�|.���5�z��w��ݜ��}\	(�d�Yj��*�o�'ёl,����YX)O z�sR������A<�g�� &:����^���~׊+E�Ks�b|VZuv^�G���24TFh܁s�p��L
g�{���D祹����!�ϫ/6�\��=OH�MP�U;P>j.��<���J��[���V>���n�#���y�e����v�ґK"[�4MXԅ�Ѯ�o��;`�D��t]�e�W滖ວ^���;����g��|�'�ܸD�h�Ԗ�b�١ͦ��f+�^�Jw�&���sN��4��w���=y�R�c�0�{/���,X�� �5U@�Ʃ2ܖ�O�kc&�J��w/���������������oB�Y �F����h��k�͠��õ���ץ�����k�wA�ťݦP,��ŧN���;3iX�ض�csm\0�v��̓޹��z��ճ�޹ٜɷ�Fj�T]ӗ�e�Zj��5n3'd{�v� ڲ������W9[v�E�˜v�Ѥ�R�w�/��������1#Đ��[��"h��t���uds^'k���os5�f}{���w����i&�2�a���q���}�e(ʡX�/��y����Mq�H�6e�-aA��]�VlT�r��*
**����
�$s�ӹ�/^���݂����޷���G4�H�;V���O��CxܡV�eV[���Dul��i����#�+��)1�ƓS;{�4��DT5�ԵM�4Dz&7�I�w�7��[�{}��m��1�dو��2g�1$���o��+G��������W����{�-�5!^������0Lzi�:Z,��K=UPjM2큽q�$c����D����[2�g��I�0��������&��I��!!!?����'��BBB_��t0��BA�g.�H�F$R;��  �c�`A"H�R%YU"��$�V�YUB���*Ē��VBUH�b�*�X�D�jȕj�K$["�Q%Z�R*�	,@�#	"$#�B1H��� 1��#D�F#0��-Q%�$�eIBX�,�Z��$�,D�*K�� b�b@  �%UYIdYYH�E�%X�)$�)Ȳ$�$��ȩ$�)$�)$�,�K"�K"��Ȥ�Ȥ�Ȥ�Ȓ��"@� ŀ��#$# F��I"K"K"�K"�,�I,�K"ȒȰ�Ȥ�ȢK"�K"JI,�I,�$�Ȱ�ȩ$�(�ȱ$�,�K"�K"�dIRIdXIdP�,�K"ȒȲI,��I%�BȲ$B !� �"ȲI,�I,�I,��K"��߿q��%�d�YYI%�`�)$�(YI%�D�E�IdIRIdRIdP�,�,��" ! �I�,�K"JI,�I,��K"��ȱ$�)$�,�K"�K"���d	 B DYD�E$�E�%�D�E$�� MZ�"bHP�I,�	,�I,�I,�"K"Ȓȱ$�)$�$��Ȥ�ȰYY$�E$�E�%�I%�dIdRIdIbIdT�Y�Y�YIdY$�E�IdRIdXIdY$�D�IdT�Y,�I,�I,�$�ȢK"�K"��a%�%I%Y$$�E�DL�H�BY"�	d�"BY"�"Y"�BY"�	d��%�*H�d�I"Y"�H��d��$K$RDK$R$K$P$�lIRN*Ae"9$T�Y"�$XAd�$ĖD�G,�bAd�,�a�, �E�H�"��Y"ȒȶE��H����;"K$TId�D�E�%�l�$K$TIbؒ�K[X�R%�(��"rX��ȤB A"$ $R#!,�d�d��,�dTIb�,["�,�E���b'd�R%�bJ�,T�%"YX�Kd["�"�ȡ,�bة"Ȱ�E�Yűd��b�$D��	I��B$�VU��I*ՁVŪ"Ŗ(,Z�UD�H�VUYb�DU�b�IV�Ő�����O_,�����)$�Ii"�!�f	 ��8�7�:�����?$~�������u������ C����Ə�(�`��O���ӟ~��٘ 3�'����������D��d���I�����K"��G�'�S�i�S�?D��$�����~����ԝJ�������O�?�'�D��ORN��?�O�'�y-���DH�I,I,�J�,�,I*I,I(RII%���Q%�IRIRIP���$�$�Y$�I%I%"�J�RID�I)bID�$�I%�JIRId���%�IIa%JI(�I)*I*IR$��IbXI*�)d�[J��ԒX��؉j$��H��ZH��$�Z�%��[ꔐrȂ�$��Al�-�XH�ؒZI-B,����@� D 1� %�%JI,��J�$�I%)$�,�J��K"�$��KT�RX�QI%I%I%�IQ,�,�d�XJBY$�B�dId�Y"T�X�RI`�$�� � �I @�I%�%�IH��ٝ��K/#��߿�?�!!!-	"%�H�Kd�$��DK���9����g�%�o������l��O���H� rO��������	�S�g��?��Y�d��zY���?G�H� }������|�1����D�?`�$�I�����$HI!��O�;�J�Iܒ�8��֜����D����������`@BI�ğ�����$����[$��=����������~�=o�~��I��S���O��q"$���������rDI�$��䟯ԙ%���N�Ꟊ��=O�Iy'����}����g�'�O�n�S���>I$i�d����	ē�d�'����?����&�~�$���1d䟏X�C��?���O����I������
�2�Ϋ�z(������9�>���`@                @                  hR�P� ��R��()B� 
$��(UUP�%@ QI
R�PH%UEU*AA@ �ޅJ$(�JA!"*$UQER�"T���
�D�RH ��IT�(
��U((R��EP >    ��*�$RJRT �}R>�˪:9�
e�fZx�]�fW<���^��W�{��v*���X=���{��+��"�^�P����Z���/��@>   ��%�  ^`9:

 R���^z
����w:m*�޸\�Wi�������y�"���o=Σ٫]��"U��u�Z�c�ΩW�@ �P>  τ�E�!J� JI��}[k��6�����;۽�)6���S��3�QR9����v`�k�T-����«��Z�ڋ�����f���٭�{���(n�  c�o0�T� ��@�9�R)�� 2��	�QK��Τ@�hR���$  )AA�  u<P(��AB��TU���;���d2���ͨ��� U������Ewn���d�J��M۠��$ ���@:w������w	(��Nm$JfhE]��T2 �pD $9 >�q� �@P� |y��*�**
H���I@D�� �z ]�@7`�� 5q�	p }��T �`q��n� ,H�!� �
 ��|   =�<G  79*�\ P�}���X�9� 9w �0:�@�;� � 8)T�E)�   >�TT�(�JJ�
 �� ��� h7` r�H$�#� ��D@n���` ��ǥ� ��P ��:�  R�  ����Cw� <nRT���q \��� � 8� a����� ���hJR� 4 E?!�)U=C ��UJ1� 4 4�*@�� �a ~�%STچ�b10MB�D�&�~��?�����w�$��$0�������I��+����8��ݯ䄄!$�G��R��	  C����$��BB������ I������/��+����)�ܠ.`���,f����䫹��Ac�YI�ٸˆ۩���q��L`��k"��]qʽx4�1�ܓE��ֶ��������e��p�(d�[����:�	�F��� ����2�۫/`fҡ� IՌQZ��U\���,��[�MLa+".])�_]����3v�.Ƽo��g[��f���ݗV��W+����T����-n�$M	*j�*n�_ݭ�Spv9�2����Ba�R�퐢��t(���US9�Hh�����T&��ʕEV@�v�I��72�W��r��p�!2f��x��7HwǸ̼�+q��).�{N���J�׺��aX����Y��b��^}��]*&m�h�Cvk���L�7b��� ���c^J"��1-83*[��Z�aݼ��d�vcvw+*�McR�oRآ-&'�8lH�д,�Z�e�F���ܰ�6�m'A�P4+-[z�'��s(.Mb
��h�1�f˭2�m�k9m��� �Г���
JK��o�*��i������יD�v��8��Se�GiĎV%�IjYP�wv��I���f�k�F���d�I�s~Ͱ����ڀTݹ	��gwn�,G r�3e
L̖ڔ��igr�8أ6��k6�������f�G��wt��V4T;k(3t��J1�!{�4����q%�����me��di�B���#��ݼ�C(�"�;�1�0��ܶ���hkF/�$  I���� /N�slfh[�%��������%)\ːZ�DPx-�-L7�h���ѽF�����r�IZf��X�FV�w��Q�Ň7+˚0�OC{t�d�N��;�i	�Lq]jZ�g�ZP���6�֊��4����5�j� �,X����3�8�<�3f=��;��@;o0�L͔r�+�O/FVJ���'" �ܺ�̰�d��Z�٭�4-SY��Jv�(��.d�˧�q`C��,�!i�w��Q���˗[%���)��n�����a�s0E��HB�2�e�j$��(�J"ʕ���ٷ4r*9Y%'x�;�If �F%V ȝ�Om�;�é��4N<,Fnn�-e��ˣ,P��u�&Ú�݁M�;��Kڏ6�GV��f�1�5��(l�Z��5c��)����Y��V�,K��U�2ؼ8�2�+c�C����Y(�s%�z�!�{j�n���Ժ�v�5nA�wB�(8�ܷ/Dʙ1c��rwe�j�0^��e�wS���Xm��w�����6��i*��SK����mՁ�-,؜K�1�V
7Z�l�Yb�i ��ɦ8B`S��&n)�����51��u�*1��둃�X�9tU��U�����]�K>�����X+&�0���[f�;[P���[J�Z�nlU$�Fк���c �B6���# ��Z1Jʳ�p���aZ�p0p5�&$c�6�`��^�
��ө[ddZ1��ud1Ӻͻ���	�p��.h����qm=�b�lȒh"5X��۬/`��&+�ڦ���.z��ee��Y�.�����,?�uL6t�oS��K�ih�y���ֽ�`7��DU��ܼ�rM!`צn�kH���bKmZHN�;��zCl6��wr⠫m5���ߍ움��j�	9�K1��N���T��M���a�ݣ4�MiblI�vh��r�2i���`�
�ܺ��^�)X�F�;��۔�2�K���
e�]�p�RI��l�;�[A��Ǜ5��d[�^l.<�^c�E�/-Z��R�e����6'�օ�j�[��ժQ�t����˲\�{�ּ�J;E�ͼ�r��V����9dc;��ǁ�����2�0���O�V�֜5���4��'R�F���s�d��Kh0��̽�Y�VQں���UfbY���*���,*��gAk4��Y�7��װ���-�%�ke,U�,VI�pʕ���k^����c�-�p,0�~֎���-`��񱦯*kUf�Q�v�)xh�/2�����P�zlM�U2ٟ^�[XPHˢ�Օ0d���J[hE&L�	��b�ASq�3�e^	�mmhwz�f3B!��O3��ݺʃv�t�e#��:ro���V��CUF�����Lm�m�����m��4w�b��P�tܼ���ڀh�����zj�n\5z��$T��Ղ Ŷ�{`�f�(n�ȡw&��CN�����W��-Z6��4&Ա���5��Rӓ�Wp�]5\Ӊn̩�(h:v>����\���W+~:�XXݡu{Ya����-��T�o/(�ۛM&���Rͽ�d��e,V��YZ��f�X@e�n�f֒r���XN��9��6
[W/U��׷�ԯ-�ŭ�u�Hf�)ly�XM�f�K��/l:�(���U�4�;��T����̏e�V�!D�fJ�lJ�e�&���;T//Z��V�\ge+���6�Q9��`�w>z�n0a��h��X������z^�f�K(M�ب�'Z�Z���e����`vV�Y�nXP�{��[�K���`�Oe�Yd�*\�ɥ��a�,��*�X� ��T�e"��d��l�W���I�9��C/2����wvVʱ���ŰXh����cX��v��q^��|fc���/%Ӻ)��s�X�����C�h��r��ׇ(̹���$�+1���M9P�����Z�"���٠�fK����Z��iލҨ��.`ȅf`)Q�i��msu[�7F	k��E�q�f9ib�yPK���@�-S��+[�$����W�5�{7307��D	F�V�-�[�Ͳ��w�f��{��B�r��M�v��Uʽ�/lay�+(�bl>�f��8ؔث�w2j"���R�nTX�-%���T)�/"9��NU������,��,]�=���4$C�#+!�\z��$�v6!�F����� Iy`Z�a{H��dl�Y�c��o�w�n]F%mY%����E�n�6+U�C�'�t��w�z�`�I���h�6���*�Uz��vk-&�,u�Gs]�W�C,���DV�A�V�b�kf�XEQ(��7�&kč�ؙ�X��d����fC��WSK���$�nV�ہV�E�nj�"�4F����-�N�fii�)/T�LYtw4�i��������٬~�˔�ݴ�P�mkS���~7�E w���Kq�ՀVcw�uU
���D�j�V��7�q#��$ז�&d-B`�/2ɩWd��+Rn�܂�Ÿ�b�T�ͼ���G��&X��ڴܫf�nX�%ym��*��I�%�=O+Sۓa���m�j�M��(ЋB�C�7f��[��jiB��G+M�!��W.! �L��[�o)�l0�3��;Btd��R��VJkjTN̤D	J�"�b��n�Ff��EV��++��|����캔�^�)h7(��;���[��(T2�%�^ň��R;y�N��b��0��n�L
�S%�hK����������X��,!uto0���Cv!;��u<�fV^"r�tӮ��.�'t�:J$�Ҷ]�ͦ�6cj�Ze�f,�^Iu�.@����̬e��Z�i����Ol�����:ܹP^�e<"�,�v�D��:�ָ<�n� o8	xEѹݸBn����$@9f��u5V��60�*����0#�S�73*���ZQ:8�Ty��BX�r�މX�3�QU���0o�CA��kic4��kM�@�Qsl"������Q�;'�{�p��c�1�	r�`���ͼ2�;Y��V�Z��E���WM��F"q�;z(2&*V�i�#����B�8�F^fڭug[�i�SNY�0jt�Y�2j�Y�RS�im�@��ٵ-}{6K�{bn�b6A-�B�w�,�-��dĉ��1�RK��d�w{�������F;[Y̻Y��g1��cu���ȦVm,�r�3J�͠�̻cK�p�̸�nbG,X*ܥ8�K��x�͡�Y�n^`
#7� �����:�fk�hIƾ9A��pl͚����YY�G�J1�{RI��	5�c\j��5cF;v��u �P�4�Xx���(6U�9�7�F"�pf;���P�w�M���m���̱5����]��VYJ����e�aL��k�����%7� h���d�2�sd�2ӗ�(pիA�ɻ��[����-���l�A�{/�+�g/b�e��o4���I�fx�'7F�D ���T@�#3�s/��M��8M�n�M޺�7,��F���Yd��S�B�ଋ(Q�WdG�)��<�2��:�Wn�*���kFe����Y{ol�4.�h͑�ki�j���P��@�ɮ�+vY��SF%>�LK�Y5�!.mkH�݄Bp��h�>�ѥd�a��6Tb���Y4h(+���P䘒3$����Yg@��Z�q�5.�@!Q�y/^T܏0މ��3V݁���L%��ۡ����4mՙ�e�2��ᚳM�I��A���j��?L���Q8�e�4 X`V��w+qQ�N�РM�2qd�ڳx�*�ѦܢR֘�Mi�mJ�@au�y�h�8��V��5��sa{X�%��,��
n��F�tf�d���[�F�fT˶]n�l1[�q�D�f�Zײ���Fݹ�Zǖ	G1Ye�M
�yYj����fd��%y���aB�@��j���܀�k�+>guk�W���up=1��D],46�Z{��j�2��M�w�un� U��4�޷�@e��dZK�B�����g7��A�'j2�q�VheLu��ɔ3$ِ��p7����(�fQX*ktQ7;�r��P6�X���kn�1�sF|�VP�Iޙ�݅�=/�`��[T.i�c6�*Ȕ6�Dp=6V4c(:D
*�����vK����)]֋�-�woJmZ75ɑ��vo
�U��Z�ݢ�t���82�34��\�׀�B�fc�I�7�x���F�ْ����t�v��j�E˨�U���謐1�nBB0ͧZ�M�Ly�����~چ�s6�(;��o6��hٙ{���5�R�-���0��ԥ267p�w��q���L��e��^U�U����@~���2�L�����Z�̈d�ufk7%L1�-c"hR��Hm���q�sQq�R��W��ie]-x�[5�1{����d��Ȉ�ѕ�B��	�{���/,���R�6Y Yo�Nʋ���i��%�nŗ2�VJ�],��������I��.��Z �
�W���2��x,�iRi*폛�m��MŮ�-�]�T�VYW�of�����TUvA��z��SEO�&����*�8�m^��-�{F��.!n��*�R"�Ra��{��B����w3n��Ts%5h8�3C�3iS�蠝Ca�Z��h��u������&�����H�i���!iڸ)h�ͭ�p�X�+u[�(RԨn���y{Iî&�)TR�R�����X�&��ܔ^�d2YE��S3B�ڙJ�Ů�R�iJ��n�1FS��-̷��Aiu&��ɶ�n-�Sc.b�+`���[x��O�\�u�[N���p6�2���˘�� =��əX�,sfʅX(��heCf���������GA����-�w�ۉ����L��4�diQIm̷��dt��/q=�{�pc�!֣e�M��%m���2��^d̆�ҽ�����8�ݣ��(L��	��re���c&KY�ø-*)f��i`!�]5�2�ݽ;{0:*�o�g~xm�����7iitnB`��Ұ��jf �ϥ�GvQ����z��(��h,���ڨ�Vi5N����YfI�7U�,����T>WuMAuz"�gd�x�rF[z�A����o&i�̱��Y���YX��`͖h��2��̭ ����@r� ����j�k1�N�հ��Oб�y��ܫ�}�n�$7�jA��J�f�{{)k�"�/ݛ �M�rR�2l��嚼Ѷ�)���Ao2��e�΁��t�Yi�Z�ej���4�bV�YF�l��7��N��f�n<��l���w����GGE�,���1:�hD�����toTB����g��ӬTn̊� c��Z�y����c.��j�� .�@ŗ6h*�)H�hI�S9�͢Q�`Б�3b�'�`���T� T�űD���`'C&چ��j��6��ܭ����\`2�î2Xj��b�Ǚz�̏[ݰZ�@e�rR�����;2^���gD)z�H�B�q`Nj�����NP��cnG*P63Fh��wp�6��*Pux3l�&b���`BQ�m̨�,m�'�0sVXu���Z��)�D5jũ�h����%�/�+-룒VGN:��C2�j�����v�Jڼ��T&] 4��H�K�qt4Z�Z�ĆZ�I=E��eB��vα�@ov�T�̠V��&<|uE�32K��|�wL�6>�֮E�)��
n	hJv�j4��"$`�tL��j�l�1+th����l!D���YKq���)]ed�W��Jy�@z+Yh&�s��u�7�rS��VS	�;sC��Z۵� le�9Joj^�M	��JO�8�`�I�C�-S(��wR����氵ehz��n���80�N�h �e:��~�9!>�{��ͼ� [�o%mG�B���u�w^�ɛ��Ӎ����iJ��ӕ�wj'���d���teϲ&s1��a*�á�u�KUԊ;b��4B��Z����]�Vm$RT��ۡ�>_m�Ld���F
Ӡ�V`�B�n�m�6R�[� &����i��F-)RV����ˋs*=x�Xmh�ᩙ{&��6�7/3h����h]�wR�f���vY!X͕c.�77Y�0��)�������F2����n���o.b�7�+O�	�   � R@P��$��$R�$�`XB� �����d$  ��
���	BY B�I	)
�E� ,�($��"��
HR@P$	RY"�"� (��$X��AHH� ($ XH
 )���H �BH,���$� � E�AH	$Y(E�" H���H��E� B(H$ )!BE	��P��P� P Y$�Ha ��BE�!d�,!$P B �H,�I	�E��H���d�����E�H��,�,��a�$�!	�`� 	!�H��I 	~�����N~6�Z݀q��q4�E]���iӟ��v�E^КCD�YS��%�P�"m)x��d7W�z�Ma�,�tng�*�-GC��H2{���嵔�NM��̈��2�
��7N���ZV�����ˤ]H�X��P�H�[�E����^R(�сgn駷��a�ޛ]��Q����u7�Uk��6�O�/fEW�ҙ�&e�<2M��^�ہB�,��ӝ��u��$T��Ż��e��;�����̦�Ht #tZ��L(	]��y�e�:�g�*�LKd6�c��\+Y;;��;����Y�g��h65�<)bI��l(4�5��Y1x�v6�ѐ�����Wf�%�t���{�}��3GL6�f��Ĝ ��-*T��]���Gv����$C"�t&ŭ�
�-���'��	A#1E}[w*�e�M����,dBōxe.��&���|nL��ڄv��h���N��u&<d��T�T�"؛��'�9)��`��J�O{�����y����b�W���O`�����}$���u�Ŕ���k5����t���%Z,:r*uL��7w��S�n4兆���s�˽�7��|�gum�xhj_
l�4u���@���Y��n��e���.id23��sܰa3"���F��Q���I��7f�	��%qW��>j�7~+;]Ğv����xb��<�W%�q4:,��*BlI-r��}i�l��,rC�rU)7yPI��Mg̗�^�gmee�Z��Ss.������a�Ж�dfZۢ1�'�/U.=3Vl�1�e��:}al3r�f�In$�7�@�pټpN�h����=R�2�P
�[r��˨�wXj�Z�� ��Y[�Zep;װ����0��;�Y��.����{�@������L����S���<C:iX�l<�-���OK��P��l[+P2.5� � V�omJ6�^�W��c�� �:���oc83t��
�u�်�H�%���tD|·:�@���WHF���}Xi�T���i�`;$�j3}vՑ20\���ʉBk	qB�1C.�(e�@�.���3��U˗�R����N��ѧw,1�q4��j]%��`&em����7����cps�w�-MEwu��&�����
��º�f�%b�։�g�Ґ䃓mmW�![���bu�J�y.cmdi5�XkU���!��z�:4�x&�`^[]7� ����ȝ{��*���U���EdPZ"U:����hv&���P�0�<�Ekw��l80�:���LḺ�P9�1��&��Ѵ�c��-�h��Dkݣ�^���/�zEہ��g8�,,���b�n��a@h:j�N����.BZ��\�hʺ����g����gN��fL��3P]yYk_[X�5�M�b�f�̻	.��
%�G%���n�.����(���<�X1^�x��]�ʶE�Is��2�n�Nh mf���w��Z%����J>�|qs��)�qIM��7A��rj����_TiS�hU������T�Z��'8��C���{�
�P�ub"��D	�q�+���[�e��ʠ����.Q��2�"����^J�>:��[����m`��X�;u��9L)���uj��2U�&�*̻|D��i��.�u�i�|���zJ$�9Դ�u����,>Y�-��/fNCev��묣y�p���^C��r��l��A�;wX����T!�*F�2�ZB��Y��nfL��xF
�omM/�7~���H9xwww��f�U�X:y��n�K	�"i	7v��	V�*om�u�*��3��5�������DNA�0�7J]_�Z�z��lޜ��zq�/��.�QŷFh;���AQ�-�UM0�D37��W �����|�氥���Q^�a��&����R��[�n�ތ��q�9g��:�PҌu��ZBF����8�(��Qb��畛�J������x�-�9"*d�F���[��6�0�_m��u���ZkH��*W��뾡U=Y|��qr��`��/���x̱�a�-��U��^��1MI�UܶB51�Ҩ�L�R���;np�:���1u2��b�uٝ��"e�w���	Ս�����L�����o��U��"��4�+W���>�Br[��@JJlw	�t,��T���,S��Ҁ]ҿ�����71)�J�ugv����E�HV�h��}�o):�7ED(�;��V�ꂵ�A5���St��gC�	
�B3Kv��0¸ʘS58bu��q%ٻ�T7���0����c�&uȍ���o$JY��ݪ�T*��]����HA�e���(%ܼ��g���)ofżxV�����4+�MI;�s��N`�.(L�i:T2��% -洘��f͸~ۡ1�j��)��_Y�hd�7;����'��gjrn� m�O�N�����&5��!��aѨ��T��s�z��2���)S��X�wqd�lg*,�z{&�6�{��+��b� ��9f�K��wR��b�F��b����7�E.Fz�΃K�k]޶��P�:Ly��7��֝ mj�Nvɉ��}���F��M��#wG���ڹX�<�	W	[�ԏ:�V��qf��Wwy�
]�͵t�ѹÒpVb��R-�-U�-����lO�Z3&�]�wR��<�8��d�^��[;ww[Z.��5;��ݾx������Ӕ�����뜣`&��:����C��i��v_nCLV�rU��ɘf��q<
��-8v=�V�oj�r�q�PA�u;wt�v�<:q)H�VR�+��!��+��[�$!=�\�ʦW:�DVMl�I�k�÷Y���Sp]��m�q��n(o.�a� �	[6j��w��S4u��ɹ;c�w�6o�5i鹍tR�MY3q��qع�7 1;ZbD�$ʆ����4�F���D���p�p���"�I�d��w]h���۠�t�4�#gm���mğorhF�X`�����A�s��X�`�t�5\ ���oh�):YQ��MB��h���6ŝ�F�qV�ו�:p�P���E����K��5oj91��u��t�V5�Wrb0�$53K�+�x0�W�0���V���#�MS5��w�Z�P���3x�/&P�y���6�c����+I�݋��ZZVa���5�7\{�Df�8��U�ۢ�;��ƌ&�BN��S(+cOr��Fi�
��}&��u�DeҸ�م�W���;�ܫ�oGG������0��b��oVb�pe�nF�������e�I��+��:ȣ���Umc[mTY��J�i:��ٹ]Vh�m����+T�Z��X�ljF������9�	���mP��jPW��b�:�Ҋ�clS�L.�] ���&*6-)Ѭ�of��d���+J-�wne�L9B[�Ν�Nc�/[�F�|wwk]tp
zS�.�9SuD��R����U)d��U��E�ݹZ�]��;��w��͘� �Z.������`���+Wҋ�NΓ�B%�]Yw�&�#Z�Η9d�g`�-d��h��O&�h����w2ƎcZ�r�F�q`����U�e����0v��)Ժm�ZH���5�+�f�B�+/Eb���b���7q��N�d}�{�ͳdX�ݱԀ��B�W�E�68$��f�ݬz���rs��s�<�6�bW��km��_<� ��D5��ὶeڨNe}�n��Up9n�|P��l�ԏf����!�e�)ۍ��F9��:*��!�����ʰ����b[F�hGb��/c)�ڈZ5i�J�v�V��������qe\6�^����u3HxG�v.�;Kv�l"��J�5��3/~Ћm^Z�ϱ�1�Z�i<���k!��v\W�3hF�wQ�6�6��2�2��I2�W�N�
���@թ�Qrnò����I-�u�;�y�Sj�e�a�-����3�K��u�m^�Y�^�ݱ���ed|�����]Y��!����E��r5χQZ)5vxg2f�&�7�r��\�L�e_7��΍����[z�����V��nn�륫����<��d��(X��xL��*4�G,+�Z�\ �1.�=r�՟;�-Դu�؏�����Z�*��H��\�Φ���w�]MTG��H�f6��/XӉK2جu��bn���F�s��Ȫ��Ƒ�������7{/��|�Y(ܖ0!݂h�-퍠󲞷�1��0�3Iv���Ҿ��7�m9ˬ��X�*� �X�/'=daԶVV"94~�s�̫��ӯ��&r6�)�zk4���0�+��4�=@D�dF��8��������r��s����<I���[�{�r�6����rwO�欖>��*�P�P���E�[�*�	�+�K5�I�
p�m������V;���V��瓞ZC��826�T�I�/Y��w[u����jЬ�N�2V��F�nS�zu��s�N;��k�s0��}���0� ��t/�i�yetݽ�G��ʸ��]�Ā�ׁ	�S���m�*h��LtI �	N�|�qh�A�f�U�%��uWN�j�**ҸӖ�+o�sڗg,mwG;�Vmh��
��L��ӛ�Q���}�[�L�r�+��T�p�V�kS���M �����[q5�3~�p��S��n�Yӫ�v̽���SԷ�ƨ�����A,�b��om��3@������u��\)q=�%卽���P�1X�͵UyJ�TSb�aQ�z���moQW�<$C`ѳ��3g�#��;| �ܓ�6C�v9��b}1�6*�x��y���$͸B��6�L�S�`�'ȧ[�ffq�Ы����Q�L5���S��4�Hڎ���ǳO_LܫM�;��#4��MC�89b�0���%�إ#G{g1r,�e��j�A���Z�+��u�@1�k\�a�n�6E]iQB��K)`�@r�NBO2\�2��*�X *��,^�q���Y�]Ι��f�z��u�� ��R�����U�[W��SO/n���b���Nu�,�M����V�,Շ;37��,�x��Pfrt���03�Ѧ�c�
JL�k$�Mܤ ��3z@ї��hI�:�h���-���x���u=�qgf�n,�JhV�ga�G�7��-�7d��ӓq��Ҷ7�L�̄�J3.���]fmNϤ,f��������N*�*&���qQ��B�<�;�a-+�\�}[ٺ��ղ��[[X2%��tai2�`��qWd7�(�\f=���*�&��Nh���#v�f�[6ƣt
Lܘ�kYv��[os�gj�w�{�o�!f��F1��yՇFgt:s�etU�]�P��D�]��3FV�Y�k9�"Xwv��s;��t��4X.=�� n��g-�K��1S)U<�-������k	�C����8���M�Z
V��L�Q�#�Up�W&]u2Mu���4�=aI�8�),fS]��x��ү_*�%�~д����s�z���cUeӜZ��J�nu��^�G�Ѻ�Z�//5R ����vZ��4�˻ڼmRQN�	��4,1YH��E�T��DRH!m<�{6a��Pє%P�4A��v�@S�l��r�W`�+��w7�-MƂNK�X)�6؆���ٛ1�S���x-_�D����WG��]�{\��h���B�:M=n��9U-��;Ys4�ܫ��Gv������=��)\�.���DŊ�ب�D��
�I��,@׻�Ct�7ܪ��-q�H�)�,`�wL ��L���5w�x$�G�Zt:�&���r����grd��S���
��QS�")�?%Sf4Px�i�L�rGE�������P�Q&̺�^Bb�ښ�)9
��9�ܙ���/�Y����앭�VH�9[w;��FZ�񭰂�z"Z���f�
�x�Xkw�]NP�V����m^�=��9󂑼��9o�)�ڹQ�B�'Sud̡-������U-C�\�GYS���}:�g,�ø��a�v�6����*`m3yN1I��ZSUF�fZi]3j�ĺ���X��h���A���Fވ��;�}�`��H�J�*q�k��p�9��͈s��nr��
�{@hC`5¸L�w�e$m�*+k!�c]0�G�6���ovޕ��I%I]�J��ԁ��6�7&�㼒�ؓz�)�䆢!^�,����
�<M+}Q2g1ܳ�[��h	B�w����F�����Y�ܫ�����g_]p:2�^X��R`Y|��nKA��#����>j��*�ዑ����6:�S����T��"tը�Q7Q��F��uיx\��e,��w��oe����(��N����H�9�����(��cM+�f��卽��Ó���V�<��B$p���3O���F��۲�f*��C�/s�ul��_�w%��M#�*�m�XjTCB�ӿ�gC�;�
���]7Y��]Ba,�-e�� N����[@���e%+���7z�:�PX.�պ�az��ӓ�;{n���h⬾v�7{d.����j�X��N\{u��,f�U�|~����+ҶfuwMQ�fF��V�{0�����Ͱ�,�S�/k��{k��`��x���D���i`�mw.�;�c����PsX}���������u��h3]j�Oj�N�w-�n훦w���b>�5Ѽ;3�d:��|l�ZيL�m�u�UVĉt�$��Vƙ�T����q�����j���s01���i������KOBŮ��wP;�n���R�6�Y�Ȩ�-Z�N�nh��Xv��f�`J�����ofe1�*��7�8�fIa7�y͠װ5q��un&�K��lK+���2�X���7��7uJǳF��-.��K��×j�5Vƛ��|���j+%֤�0;�Q?�\�n^e�SS[��06����4��Z��m��V��V��C��..�5�7�HҮ�P,���7ZMi��»�A�r�s�ޛ��9�<���t�?؄�!$� 篚RfWL�eI�l��@��0�N�nuuÎ7E��vP13]�p\�Cl���]���f���d���F���t�d��/#Q�������3M��j�EEf͆�p]Ό���ni��*	m��۩mH�C���,⎭n��	F1)fN�uc:u�n��U��]u�#�B��l���$r�ͳff} �ø��r=�:4[�l��8�^��Bvbݞ;��r�-8��z�ɨ]v�pKBӬ�n���r͖h	����.��v��]Z]��"=�3v�VͨΠ��6;A�h�.�pr�Ody�N���.��um�=bܜi�:|>�<����V׮n�X76��SŎ���2m*�Xv�WWZn �SÍAF��|3�O|���9]�����i����K@�M�/Y`n�$u7u��a-��\�s�1�#Εn��^�n8n"$�]�\�i����m�r�Y�%ˤ�x0:h"3�k���[�yл�㗭�N3�qc�&�����IC���[����X)5ڴt�34����1B��� ���g˭��WXC
�t�:�n���m��m�h��ZP�J6�bXRE�b6hiIKc� �0����vk��G��[f���O�a�]��z�d�݀�j�]��K��^�ڌiM�ǋ\�.:�[`��^�0m����7n��D�g��_��l��X���b�	Xa�H�x13�h;f�Jͫ��@�8�	�q�[��híɎ5/D�̛Hq��`��]��΃ȖM�3���qZrӆ�mD��9�:۬�D�q+�f�`FxyK��XK-r
:J�%�h�b@j�0!d`.֧�{�7Z�s�N��-�u���ܜu����:���uiۗgPn�]=Ѵ�ͤ�����alV���C+��uD��J&�֐�@8q)]D�ݠ��ѯ16D^y�Z̺8�9�A%��\���Ipi�u&�r.ͧ$� 2�Su�F5x)��9����yz�s.�7۳�u��A�q9�7&{��ֱ0=��]���L���%
�@]�Y�5bM�LK�ɛKn�a��$�p�j�א��Gh��mǱk��$�n�]h����;P��7��c�r�n�̏k<
v2:҅6:v����vrk��z�0��9h�9��E��^ b
�l���������Wk��)�J��g�w!�Q���ͷ�݄�F@���cU�����@N��uv�#/p/6�vIN�atz�ְu��(ْ��u���lK��ID��p�f��(at]�,:�v��g!A��q�e���&�0���u�<ջ,.q�vj�8b�\0Rۣ�:��4��QdN�"L:]4׭��Jk�5�σ�.N�����+ejMI��&�Q�y-��9��ƹ;�f�nT�9(��y�Y��+��:��cs�x����
���i�CY��$kl,�L�s��>�Ձ�[׍jWk(��Y��z���yj���̀� ��PtvY4'���^Y�ѹ�R�Jtg��ܝJۦ� �f��9�C`�Z=�5΍�Ӄ��ݖ;G<��ni�q�Ýv�1���y�'�H�Z�ή ��cK�����l�V��q��]d6�"�z��f��_<���h�3&@	��h�a�le����cj��OMu��A����7.9�ٽ��ٍ�����/���i�m ��<ݼ�ɻv���[s�۶"md�+GiKR��T�c�]��m��;9�3�����c��6�KnpKI1��DfX�b��Tԗ&�&%U��JM� z�nѝhwHq5�gk!Fcd��ֺ����vݬh7�k�yË\q����6�1�B�r������7PХ	v��	�e�֏
��ܠ�g6��ܻ�υ�b����MX$���b�+���G�l�0sً�&���JZ���2^A��kom�v��f	��)+5m��hS�C��	v��t�gH���X9{��|=>����ոᖭ�ҁ���k0��#����z���.�kuM
駹����j.�8�|4��nD�pV�S�}8ٞ#<��]Дl1MT����o�V1f��k��p�(2�3�p���7f޸���qn�-e6�ɃS�5��[��p�&g��Q���\s�<�tv}��F�@�ն\A��]������h�%���mB�Pf�ɉk)eѸ�9�t�:f�;e���x�&涍������>��Wn:�q`wl���gn6cT��y2`��è1����4�n74nX�8��B�@�,+�<�k��|�u�j���s��e��I�]Uf���.da�	�u巍��pd8��\�n���KjF`n��$Q�v5�[��/��h�t�y��I�-�ɘ���� Jk�f��k!l�'�%�� �n�S':]m�"k-��5����5�7Bb��뫨�o!��d1��nAܜ�[�Aj�:$��뉡��ZЙ�Ŗ�F��u��.+oW����M���h+�MY�K/mI|���0�Q�0�-�9���v6�7#r��c��"u7N4�M�.�u^uК;l�.���i`Itd´uV�s�[Z�	�ŵ���4�y�nو�9��7��;-�x-3�nڙ�s͎H��Q��յ�bmu��CQn^v�φ���5��q>t�.�s�P��PSjC��0�y���'6����N���c�c��nF�ڲ��8��w[����Q[��;�o1�nL�9�5���:�� 	z��.�m���i۱ϫ`mۋe�T�e�
P��\O� �:}'�s�[qMC���aHF�k�z�lf�@�X�_<'��f#IG0�v��nư�C�Y�vF�%6(q"������m���Α��H��mn��t�x4ښ�$b�[�)J$[݅ݢK�]���,6r���Y �,�7�P8���٧8�n9��l�^c����n��6CMk]��ݜ[Ps��;��)�z6=n��Ŏ���;�GJ(�v:���y]����󙸸w���{z%y1	8�+����BX]��۷m��,-q�MJ�X�᫷ 9�Ok�,*�p�6�h`��q��K�)��ڑ����f��u�����{g�q��݀�z�m���N8[6�	�X��R��kI]K154ͦ!�f�f��v�G���v�=ve��-��p���I\F�w������i��:D�ܦ��.�:�T�{�*�m%�@���v�#1�@�Yn����GX�v!6�ԛ��5�h�W���JUhY��Ncۛr��y�P��j�{\j���zD�l����R(�])��&p�jƺ���t"���F6f��&�Pޠ�չ����$�z$a(ǫ��YH�+pP����7lvN���fQ�NvG�1�AƥhB61�m��f��)���2�G`�3�*:r�#v����ݸ�ƫ��Cv�C�<ݵ�H��S������]�9��ˬЁkA�0���ݥ�ԴJ�	 ���q2^Ԛ�ru��s#���T�,��݀v��k���nnv�[�����$�5:�;8dSVZ��.v�棰nT��t#m�C>��9� 2\F����-�T���ҁe���Yq�'sg�d�r���W���v�����J<�:i(�B1+��3]���˭���E/+
',A�V+�'<꺗�f����u��i��@m����N1s���uM�ks��b^�	v���[��f>nk��=��U	r]�����Z�'���ڠ�u�Y�qt\�-p�h���6a��k��{���g�#Tٶ�ilte@��g f;�b�N��V�i`v��y71ѺCt�v�s�sc���=]LZ�&&y���1�箞㺝�cj2�)p��Jv��g�f�1f�!lٸ�����mU��
��On�!�1h��L%����kO�Is�8&�권�\>��ةW�Q6w[T;]KpX@t���":2mh��Tiez�Gc.�x��vk\m���`@�,��Y�Ĥ�s�W��\r�<�Sl�{�'��+4�ظ�sv�����Хq.���F���X���S.j��ݧ>��A�[HN�8��Ͷ�<��3���ѱp�\q�V{�6��-�<m�ca��]m��knuG8�{63��P��.2���,cڭ�8ꀆ�9��p��=��cj�F��Ȇ��v��k��n���y!�Kێ�^&�f-�8�lk�[�0�mn�(th�y��j8)ɬY�#v"��V����u�WW*���e�gO��Zx�ZF�f�9	��e"8���4��D��u���ku�u�[[mu�A4�?|>|�m�;X�벪9j�!��R��]x��R�^�5�B�X�N��L�z�3W�j\�q����q�-�[�qn:��r�a{U�9��U<+��潎��m�[n���݈�u�	�q�0)�ηB�a�ti��V��6M��ص����fx���r�ӭ�pc��b�c��h���ԙ�D\q�);�H�J7�9'�g�'Ip�����ɑX�'F7�OS�v7�n#��W�vݛt��m@�W��4���#���hy�w%���H����h��2�0B+���.�<�r�v:Ka4Z�u�F�.خ���ɍX:�l1u7cP�;q�	�pJ����r�0�DD�LZ@K&+�����eqpF�z�6�1��u���J�Ɏ�8�G=kjB��A�Jn^���6�u[���Emɬ-��`���9�F�qX`�6�/>̑��2�b[SJK���e3R	b܎
s�c�,i��<�I��Q�����]y56��[dn,>r��DS�;eMj�v]�s��E.�Z$1����OW�ǟ�`~qi���Ak��Ԭ�	���uѶ4X*'�zj��\���u�.l�3z�\����y�1�]�1�Zn��6٘�]k��?+q�8)���i�ٱqQ�6ׯU�h�N���q�s�.̛�Z���34:����[ڮ��u[��f����c��qU�9��춻�����t��mf���&K71��61&�q��{X��4l�5�I��fs�{�Ͱ5i7T��WujL�i8�U�Y��H�gV��^��0��-fW=n��N$��^8��Tsj�T�q��+��9]����,�]y�3Iv�L;5G&�d&�K380�S2��L�ՙ���33ZuVuN��6�L1JK�o{�8+Z�c�{��7�ժ�m6��ƭ�PF5kk��`���&�*b�um(�[Y�T�h��R�[�,�J���3��X����^�0�ד��hT�Y�7�o[Y���6��Ì�7<��v���iZv$����%�ZL�{�87��^k�3��1�.'V�1ж�s��0I�qcWL�{׮�kZ�clө�z��-�%c��u���1��F:�e�N͇5kz���謦i��4U�!0�;0��o�����a59h�ź��y��n�B�0�ϒ�z���`xi�Z@�u��v��Qe1����윇������T�[#�!4լ`@���KI���:��l[�� a�ָ�K,���0&�3P�K#0�cit�!l�f��rr��pWe:s���8m�:5puɣv�ݭ�J�f��׬�����dnp��e@�6i86��8xF�.��;��1\MN�#��M��oF{(�si�����Z�m���h�]�d��Ƴy�&3�Fv6�v����/l��Kv��g�l�v�:�9v�=����c��t��]��p�����l�v.�u��G8�e���b��	��\�1\�b�tu%G�%�0{.ћ,o(�����ڑ=�0螱B���+�Nzњ�C@v8��D��Sib3CT�;:�u�����]������cA�5�mL�%˱rj��2%�YB[pL9�,)Rm6��G���&�����m� ܖu��l;>J�<۪�Ztb�1݇l)����jz��bJʜ�46m�l���$٬8�=�Z�v��@�{Q���nh6�`�<V`剥�W�#eKm�S8��ظ>?���=ɣ�q��T�TK�Cm�m���dc��N�ՠƩ��\��F�4q��GZc�c�F3�s�3�uW,b^�ێ�Aͬ�[�	lk����f԰.���[�[��J�vד7�tu�]K]V���nn[z8ѳrYN���㭗X�<�#�t�o=���	�oXl�#�Z75�Á8�dm��r�% $K�-zո(�iX̉u�e�l�*PU��w��wV�<�q������0F��y:M3R�b��nyP@%�6�79��G^�8:䲦h�n���-���\)���q�i6x4ه�v5���m׭�����f�<��n6P)��w1���2��͆K���������$��k�vu�$�n%�!���eiIV�֋6�2�*E��VVV4�)���:�m�	KX���z��	KN��e,�k��0+J���V��j0H��(��hT#^B�TYl%QXuJ ��l�2��Hq֋Fp�l��mX��ZZ�P�iBUIjJ׭�-���2�����}`	�Kmv�16W;�H�&�!/cc!:|�Ʒ�!У���K-���4����t(6򳨩םK�ۙDwLz0ud*��-��unD�4���P�_� �B��cuӇiw5����졤\բ���R縶^*H&��A��Ƅ�נ�)K�Ґ��{+@E�^
L���esD������[��D��ѥ��p �}�$���:D��!_D��CM��B� ����R#wdO�"�����;-t��U/�ŝ���w�?>��4�wy����g�f�ȟ�	��0 Y���ok�����3�~w���ق!�J����n�cEN�f�nV�gf )"�����3��&��s�j��^�Z�9�-jg��s����x�cRA�3�H#L����Ӯ�9鬸� �r����a��PW�P�X$֤��n�����J��讋����v�_�ʖ�L��7Ve�;E�I�ۼ��9�k\o�+��$HJ��̹�F�U�}�7,3��B��{�}?^t����9\1�n�<A���ٽ� �L��|��~�S��~���z����$��	�<}yHwt�e�ה�<Z�*O�؄�z>�wuI���4� ꦳F��"��_P��$� F�Ȝ�:�s����ۥ�KR�� `/MY�/[�c?M����Q�RK��$�ʡPUI.�ۈ���T�̬����z�p��J�x�z�H �9`�wvGn�f7�SU&y^J`�Q�$�����n��Ŭb3M!r�e�x�\�Sy�X3ӕ�ϨP�Q��+��P���ztw��-O��M'��R�UӨQ���^��P�%�A�>�_�̯�����WH�,��P��W]�j�[�-Z�N��'wU��W5X6@r�O�Z@�wUwvF�
�e�U��6�Yvj��1n]�o�s�����rp�����W`@��wz�uLo�\-���a�'&�<�킘ܻ�\�}zm1�M+t����R�3F�?��'㻪H{{�B$I9�?_5��� \բ�뼥��5<R>5؄�F�S��W�Wg�u)�H#L	ݗ�(}$ʨ9��c~��������+[����تY}�Z4�. �F� �}�$��#H�.w;Z4{$� ��P&:�8g�r��Ӻ�.�*��;�l�ۑ�ُ�æ5'�S� ��BA� ���wvD��^���fOS�k����8����^�(|��#;ED�9��r�"�i+����GU�L��RA���sV�k�s����z�hp5؄�O���N���6���\Ȑ~g�z���H?l��싽ZF<�N��fů���] �n��H��Q~�y�^!Ɠ��a�Wj���;s��`����}[�"~���s;�3��u�#�� ��3�3�[�ƪVs
�4]ݶ�ʃs{F���p4���h�B:t�=�c]�1"f���5�\�iՋ�����B^%�#VB�͚��ϙG��<�.bq�Ns�c�r�WP9���lV-�<W"����^l=R>�Mv '��A�� ��C4����>��������\7��)�K1�M�n�.�<.�%������4�J<#.Bk��h���^�|�����χ�|d�Mt�K_�3C] �n��#]��T��v�f$3_Cܑ �j�@�����]O�oVv��X6u�
N!!��o���%[��@ �R�vdg9��};�/���3��;�o���ee	%�

�PE�)f+�"�~׺����m��P󜼉�ř�ov��]��<��Dy��ʕ9�Y���iO��m��|*�?
�y�ۼ�~}�&���I�s&y�Y�����D�*�]�$P�|�QW;���:�p�OU)"�'��vF)�IJ�GU��t�	�ɢ��Z��6�ʣB.r�Y_]��(�y�ٺ�^���QdvuBEs(�
�\Fp^蕕c��x;wR�Ov��:���Y��B�s6���0����Ύz�l�R#ڝ�T�V8�ZFy�ݸ4��kg�Tj��z��5���k�q���C�6�mB9�ZK�������5�EMɡ�ԋ-U�FR��m�3�+�,e`�Q�L�i�l�tSm��w.��lU�Wv�sZ����mu���F׮=B���դ�L1t1W-"�R;��G7X���ϛ�����\�ٔ�"6
��$��q0�p���,]��fW2���8�o�S֢<߰ǜ�����j�ӧ,w�9����ʕ��û��ٱ�%�}x�9�0g*P��/>Q����u��q?	�)�ɧ�Ɂ��Z4�/�_rwu@4��4<7�(�<�&��̑�S�U�����m�hE�]5]IǪ�Z��O����~��q=�ِf���-���6��s�;�kY���A�#��F5h���9�1:�}t(g+�B���C�4�Z��}V	���f�Cڴwwf��Y��zO�4����Oד�H:�[��"�h��e���A5癹��'�����=�-}MX��\���h�R93K��v�c5Tn5�8�2ͬ�� 9����~����YXw�2>C�̑#�=os�/:Lc��G՝����y��D���3Y[�X����L1�f��p'5 ��{*'!'D��ty��^vX�����r�;��,��ʤ���G��uy|�@����;le:ՑӦ.���d9��3�5|俽�
�j������lpǆ��w�.А̈9���L9��7���ڑ��H�~d@-¡C��V���Z�_��<L���ᓯ��j��X�KFV%�?_@���~!Zv号���n��5R�yW fd�;�������Ɍu�� �z�V� �,|9.���;��w@G3�H� ���9��y�%K�0028��ϑ{�R��{�m�@�� �Yd"fH�<'c�bX�F�}2!Fg��8�8�iM7dyíQ'�튩i�=i�8ڮz����g뤽���>-�]/'��;�\��Z2�/��el���<<�G����0�}��H"�-�����-����!1��j�X�^t��_.�����������B��i���]]~��P��3  s1H aW�)�ۜ�-���`s'G�e�w7 0CWAu9��������v,%y��d�ِ�X��iVT-U�Ƞʩ�k2B^�v�i���܋lH+� �_E���I� �>JQ��,KEС]VU�?�+q�.����(��p4�".��^��}���>o/8�nܱwv�E�n��W*`��Jx2�\�}���VRǂ��:�tz�y�H?d}��I�����^�=�lt��!F�՗)�[oY��e��\��fԆ6���8��
�=�~K,��:�p��b�	v��G<�Ѽ��Ă�!.E�>*v�oE! AdG��B �d�?ad}�5�W>ꅢA�b>=�.��ܾ��d�v��/��  �|���3�9��4q~퐾��$ّ��o(�U�+O�i^��WnJN����Ey�ʱ��fԨ��,wv�'��3�}^]����da`�&�@�b�~#.�{���{�m�p;hIӷ�.l����4�Z�ou5�S�%�5b�pd��:���U<"�+�pS������+�x
���u�R��Xz҂�7@|�ቭ";�b3wp����e�ޞZ?���z�.�tl�νeD�K� �A�_fb�AUY?:/k��.�R�mv^��<�x�-�$��v���;8�5�#J3X���u��f?y�b���"<�Qݫ�d�weYK7E�c�舋����9ʱ�{�	��`���F:�s*�^b�Xώ�R�D1wx�ܦ7��6ؐT���C���@���6�1g|��eGv���mTM�:T��դ��˾N6Mg^��V%�4�� s1H �F� uS�_K�����w�����H ���$p�}ݵe'�-gj�< z��=x�]k����>쀁���`��3v�#����~��g՟)�H�>կr�����bA\�vП��(�6(So('�9��2�D>��:1�U���׹z���mY�K;���5�or��jn�7`lf'���6���@��2��Ľ����!2�Rٌi4pŵ��� \�.m\�I��b٭¬uA�/#o;�9lP*����6�b�t`Ő��З�˜#-�%���cK�@�bkuW$Ɋ8&��H�,HXm��&T�- l���⭥�춮��0�jEe�\XL�
�	d02���5X�i��N��F�OFt�{e(�S��:��a�c˛���ߟ���x��x���5�v�F�|�d�#] 2��a[F�F9�]V>f}_���a��nч7ݭ˶�Eg^�1�p#[���Û��k��潈�r�~��!�&�.�ف��E�˜�;0�"�dHb3��j�OtZ���|H�\"�H��؆HRxf���C�,����Mi�e��x#�o4�o�6�w�1�GR��|-�lH+�&vГ�?fD�Ff!'�!�׎�s���Aul�?tG�f!ՙ;v�rZ+�Q�H�@�lv��!_��
|�n��ݳ`�P����U��}���}�*���ɲ��X�¯�} ����BA�">#1}� �z�	�"�b��lR��!tqdE]v8���vC�[I�q��2����o������ݼMk���7�Le�-�@�m��$EqSh`��P;ʱwp��T.�C�S�}��h��������\�b�%�Ct�h*�v��X��N�wMhӁ��ͨנm���CMԖ�q�s�S��2���u!���������Iuu]����c����ъ�K���s1T������k=���R��W���0.��'�B��k�i=�K;*���O\"���e}�9��yOlTV�oIH��6��F�ux��Su��lP+��BAc���� ���5�X>dРٺۺ��v,����+9���f9h��m�ĸAc�.��v��S1�D��*4*?Yu�9���\/�չ�M\9	a(�1�ɒۤ3�,]�uW���б{�l��n�������i=�K;*�����폲��;�Dݲ�wo��y��e=�ī��˽_48M�G=�c.�1m�p;hO�ȃ�{Nq�&����]����mTݠ��3v�faX>��G=����"�SM�E�ve�#v�;�Qw���R���!fT��	�h����G3�c�k�nG��a�d���w�^���Q��޸��V!Z��HN��Xz*�,L69�>Z4��zl�m�Y�!�s��7��1�Vx��4�Qv]���$�+Ha�����ƶܶ�����'�T�w�~�IE:,m����4擡�����\�v��"�l=�C�\��qV��OJ��gw����8�o�^�$����u�\m���Fn �k%�+(n����8����k٫Y��*�wVr���M�qL�\W)�*+Iy�j�X���^�Pw�nh����0��u��+�c�*��A�3��V�_A��A�!.��i���������	'�P�Ks�F.�N"�U8}9ǟm�ǺvĬ
��YA\�۵���=�ٓ��tK��v�Ni�k���8�Z�Y������ѣ���$�d�W��3JXh'\Wu��@�9��>�Z�[B�)�E��"򄼼�R[�<+�ZV͢E��W*�r�x�P�2�g-�Ii�鮒���R95�՘��HPs����y���վ:�k�f�59y���عm��oV�'\�F��#7\DنX� �}�TМGm��8�Gg`���5�zݘ�;�Թ+��u���йo�4��ss�'�ԽK"���3Pj���V_�K�����Y�7/2��!eU�b�H`�-VHӠ�ړ�)T��=�*�α=1�����+���ѩͳ�ދU���A�ک9��3!���)SL�5�:f8�Uծa�ٕ��tُWfsZ��'Y:4骹���;սhf���4��%�cia�WU��6fW(�d�;Y��&���q��rӉ��N��n6��g盽����v�ŵ��s�n8�Z�V��cet$�*�&lc��Ev�d�����ʻ:�籇���Z�gK:���ei�Xrh;�7�6ad�e�u�*	Y�X��`n�k���k:t�L��g1��)q�J��`���Z�fc2�͝S��yg�a�41��fVH��f��&Yls:\�a�``��V��aµ��Nr�Α�ie�֔�1�a׭�q��{+\ls+�����8�3�ަq���c8�V����0�i��&6�,5�`d���:�f)F��T�hR�M�����s3c0�զ���H��T��PV�����Z����}���z�|�1? RAe2R��R$���~�ZAa�� s��x!I �* X��Xs�8�Rw�����_���y�����}��Z��$��s�f%$)s�x�X�~��E��E,�ew���b �?D�S�P�Le$�y�w3���������<H,�
��]� Ԩo�H.0)�嘞�YQ�������
�.�X`~@�������x��Q��,��?}?����� C���޹�s�[c���XVP~H)�혐|��Z��$�@��Bٌ��P�7u
#�O�%G��/����.$�L@�D�3�s��9mv^��U�uhyF�iE�r5�)���̼����W�0���X}ʅ�c) �Psa�A`yH+ʁr肐Xs�H.~�y�w��k�����{m����,��) ���o{�������{����T
C�$���;P���P?olĚ�$����bRAa�Pdq �s�bAH)�����gs�;կo�
H)���[=) �PC���:_�����{w�8y~o?���х�����- ����� �<�$�@����{�����ܿ�)ʅ�C��H�l��@���d��@�,II�9P�����r�I��R
�Rw^o�w=+���}Ϗs��O{���AaYA�H)
��혐|��Z��$�
a�T-��I
�9g���
H+�ai%��;�7~x|f_��k\���ZAH(oۇ���IyP.�#�b>��>˼ۜ~���fy�E{����b~@��ʌ����R~|>��`�K�,ɨ��*|!r�U�Cgi�����7�ŘU�����mWv�����\�<�l�,�ᝇ.�e^��w3{���)�Ǟ}H,?)��f$����C)��H��Xs�H)
��嘐|(�$�
H)�9P�$%s�o�����s���ЇD����w���.��Vn�? ,	����	`��~�C&�(Ba�@�s7�g��3�/4f��˘l�+���ӎ�A�2�v]����`�9�%�u�Ke~�x�����I�)���$����bAa�� s��x��$|	��@	����s���ǅ����AHVs���^w��혐v�RAk�i-�}څ���!�r�#
H/��RTB�s�d���P9�ݽ����|z�X��^�,.�)��|$��2:�n}�Iyh����Y -�b~@���d��
BĔ�XQ�\1 ����r�IU�W^]{�H,��}`R�I�v�Ă����,Ă�R�*���s�fFJH(�,Ă���oߜ����z�7Oodd�{[Z��%�0���X~�B�2���^��<H,H/�Rr�i�`R9�1 �{���|�;gd��
H)�7�H,20���1'�RAd�S� Y�_yÿy��~;�ޟ�R
�i!��;�bA�Q
H/���?}�y�����H)�0�ꅳ �I
�~�Ă���.0���Xs�d�RA@��9����I������x|	��[	#�L�o\�z��������Y���(d��
BĔ�XQ�\1 �s�bM������?�����1ފ�42Z{^�.f�K�)h�ܭH��e<r���`n�jc�+!�4*�z���s��j���?!\r��@�5|�e��e.���\�\wqOu��S;<����=]�	���#�a⋂=tEv�Yz4��M���1x���k�e��c'�H����l;,����B[�OKq��j���Ry<���۫˥\;�\P��yt��u���
sL�"�4�%�l�n�]Gc4Tet*�� 95c�x1c�1�"`n��;$�f��ɞy�8�/8�7`�i�,�￧����U�bd��� �����u�3b��۝F�3Y�͂&u6���Ζ����.��HUP����R
A|�ہI,@��B�
AC"�,� ���~󑔯�*�o�}�>� x�D�~��y\�C~څ�te$
;��Ă��H+ځe� �C��bAH(�,���)�������������:y\����x�Xz0��lĞD) �P�^W�A !�q��x_W����a~P�
B��<�ى�!I���QB ?��#��]����(���Ԃ���l� ��0����
H)��T-���H(�s
AH+ʁ�� ��*�_?jg��E��s5��įhY���@%	'��*2R��RRAaS~�bAa�9�Y�<B�
A^T
@�) ��(0q �*�w��ݷW/n�g,ă��Z+�I,@��Bّ��
9�1 �� ��~󡔯�+oo�}�>����B�~څ�c) �g��ߞV���r�U��ߟ$�I}�]R��bAr
@�9f$��J^T
B�RAaD�.�X`9�Y�;��n��$MK�|]������y��g�����?G
B���f$(�$���RAK@��Bّ��
s�����E�\OJ�x�!*H�J�!<G��R�p��.��)˴�c���B^�5�SO�- ��ZAIB�ߪɌ���_�w�����.�)�#�	#�L�������9�m���Y��@��˯��x���r�%��HtII�}��
A@���l���@�^T
@���Xs��AHUP�,Ă�R~���i��j����k�q�Fڮ!ylX&��״U��I��x�{�2=����C�gn؝��Aꤠ�Tok�GS��{>��yg���W��S�0��Bك��G���BH���;Ͻ��������=�^	�B �y��:���[�W��O<��8�;�\wv�"&��56�jo��ѾU�����f���e!��ݬwl�k<�����#���2�l@:�X��]�g9�EdZ\A��0����9�q۵$F�#1 ~9������>�Փ'=��h�`7��^�R�\F�Gݧ�
�yX>f�͚�&�D�
{��3��1�;f�f��)e�Ŵ�r{&�Ĺ�-�Ϩ,�͌ ݅�a&�g��T ���3���-`֫E�o�f��	�Ț�f�$C1M!���3$I� �Bg>���v݅/y?3�}��J3;%ۦy�rc"-qL|6�_�O�r���t����$|���s!s2A��B�Oo�n��5��'�In���
F7*.������(s�Z�ӵ��ja\��mƃBiF}���N��ª��bQ��TV���}pi��S�_lVf�DW�G�w�+�~_��/�1YV0��rx����5|���:��:�1n��Ƴ`� L֡$2�a��S���Va���L��|ɠ?[o+�n�i�}F_o��R�7}���`�U��
�u�9��~#1�����Kn�C* (��6�Vz���p��*�7&��ezy�\m��X���6VS�y+�5睳A�(wj���3�ӽێ�t:���,�Qm�b;�p��EDݹ��� ��"_{ｽs5���qW��P���={ԟ/Y�f��@�;hH ��ّU�&�Pu=a]���;��D�܆�Twno�\�pӪ���p�t�1�i}��0?[A�RA#ْ�e��_>q���b?D
��Pm�g�w��]�<Y߬W��*bk�{�1��̠�nn�e#�b��ڑ��x�ʞ�^4-5{��	/qc���<��ж���6��m_�I%����{U;�-���5��.;����b(0=��'yS����6w���BAD|s!|Ff w�Ȧ�R������2��L�*be@Q0P�$����j�I��=������c��g]��l����6_o$H?a�b��W^��F2"�.`I��w��Aϔ�H� �ā9���7�OU�����@�� �Y�'`�s�U�^8��=f�] �p�5�"O�"_X[+�H����9ؤ�� f ���$»�0i��u���r�	��2pT4רf���V�͊��2j��L��'!��Q��}��5��`��+z�F2"��+c�1��g��9�|9����ݻ��f"�|.��5>�*8��
wzn���jA���B�ڱϷ�6�Mڟy�y��F��ʗ��\e���eFn���l��;�]���v�z�/����ɇx��'��T|pg.+�Ǜ}�[<r�0	��)�⊸`�I�������uȨ̖��'3m�t6p�/f�&C����;�NѦ����`�:ĉ�wm��H㴩s�fG;�v�V���������X��Z9�NPl1n.�:k,5�XCB�
,2�Z�t����3"���[(9h�n:�ݽu�j���F�ݢ��k�=�.ћZ�u��q-�6�Ȯ�k1W)�E�[2\1�L��+X�4-��%���_:���[��v�[*���0Bi��&f��X���,R�N�qvuD�2�{��~���~cf) �0��x��/���l���ɳt�G6j��%��"H��$fԡ��O��9��~ݽo����Q���
�ҷ��DZ�$i�-�G3Q��!G���0Ch/��A8D�B�o*ߕ�xf���߀/R��k���俊�ڱϷf�Fn����/kή��N�'�_b�A#	ܼGy1w����6r�j��b�FM�,yV�s��#5�����c7�T��d��S��:�B�����h�%_� �4� �A|s1} �<�Q���%Κ_�}n�}kQ��N8���'E�@�z�2]e��6�nG�Y��f��6���=�Y|�����A�t)�u�};ݸZƳ:T���<k�Q&���^�(Ur�YC�O͟�v��� ��j�. �	 ���I�lS1�*L��vh�Yy��'{��Og�A��Qf9IU"'b)�of�+�Q%N�N(&���z�e��E�U�k,Ǉ�  ����/��bo� x��gY�j��r��n����r��h��a�6�F3b�o+1T٦vEws��"o�Q��\��d����(|�u���d
�p���dd���5@����ӽ7X�d�V�P�C�D�	��u&\X����3o".���n��oy�}���q+���nn/)�	�h��kP��2=���_��2�?y��#����^v��q�l�k��:yv�x�f2# ����Lb���e���?���S|���4���Usճ�d��o[�MTl� ����A��e��P�ۡ!)楻��8n�$��ӽ7X�d�V���P�<��tԞ鑻�y.���r�O��9���p��0���G^�������b��&���!`wK6�u��6�9�������f���P�eMz���{�C_=JN�ٴ�>e\d-�K1bx�a�dl�����̃��⼮�N(����q��l�
m�`�>��GR��`��Ȑ�f!���<�l-b�����J��+�����>�����Bn�cݰ�ڔ�����%������Ss�3�6�'� ��U���|�O{0']a-�<+��=�e�l\$�6�t�=pc�m�ą@�c]q(;il\�Ұ˺3�}}}B�����Du=��ȍgZs�޵C}WV(�{����w���ϪS�գ��dMe�X��4���#���c�f�n!���x!vb:�k�w�ADP~��v/_���!g�)�)d�BH9ĀA fd���E<��o��g�����ՙ%Cյ��P����~�ց��e�����}���3߯Z�B��]PR^|()g�"5����%`� �������F�ucy6�q���T6�(��{�N�j��־�j$h+��`|q�#n�4����l�]��HV��W�w�5�ڴ��e�xp:jo'&�:�#wh�و�
�NF$����9���������ڳZ%�ڊCB�"�̉S2k��㠚F#h8�nU�B�eѤrb��?z��ﾐ���d A��A��ڦ2�e�;�"d[��,���W8�D{ a�c�-�����y�϶����9���x��[���S��qj���dG�(whϼ�o���v��Z�������㘁��dӫ�ꪛ�B5���O1�Z��ľ�Ag/�1XF:�����|z����=�ͩN����'�ٯ�Le�+���xN� Oh�r���y����|�g6�����R���ݹ�a~�~{thAG���+93����\�����3#��B>mET)�j懵zw4{�º2K�*W9q�d�Y3I�R������ E�*iD�ɮ��G\뼎^̋���,�n�\��Vy2�n��s)on�yև�3Q�m�'�<�fޞ6����ץU���@��fό��l>=b�V�C��wd�ז�V�`�*1�[�Ng[�T�7;_Q.�p��'b�^>��d��bg
}��w.����u�9�G�h�Nƨz�UqG8�u�1h�������w0���9bb��yXد�ݫ� &�������a�V�9����(f�&�׷�I��gg�n��E�#�����3s�\��&�V��)R�ͣ�ٝ��4�è��l�:UI{F��(ܤv��)$Oe���c�ܭ���=��D����z"d�g9T�_�$(u�E��Q�4 �ڏ�N��E����+0�B��*�fO�Swe����HIg%6Q�U��L0��O\}�>�܏�W��,�M�Z��:O(K%��dn7xlX��YPs6*]��q�X���ec�`⼤�(^��~��W.p�1dɶ�Fj�X�ˬٌ�|���&w���R��Q���9��b鸰[Z4ˌ��ّ�x�8d���Eb��]�تvJ�l���9�۴�㸞:;mrv��gp�	!}�YWd�=�<y��ECn��_i�P���f^�^����4|pFey��� �ݵ:P���]�a�oVd:��r������!=Y}R�
r""@��^G�J���BCZ�*��c�4
�nn%�{:��1Uc�$DMM26N("'4��K6�N;Da#~n��leu.-��FtTgXiR�f��ý@��γc��fo{���e'O{y�Ns�V���޷��f�M;i�\q���g����n�1Z�i�nU�w�����M5�Ί��4a�nf�fN5�{���Z�8j�E�i�ݍ���貊�3�m;9���l`�6���ey�<;գ�m<��^���c��.�slz��ۛ;�n���ak�qZd\J�M��O{��^����{j��m���Ϊ/{{<ڮ����ΒI6���[U��+ֱ��f�&�a�����3�9뽏Y�3���z�ݴ�c���0۱�ZN�b3�n4'���Uݍ�4��Nm{�w�7%��ɪ�Z����R���~s�J�tיf���(n�U�t$?�<�x�`��ۙz�x2�h��F�	[!��b.A%˒Nƍ���0v�e��d\ѹ[��9�W	UCF�rvֻs����2]A͍� Lk��@�vX5�TZfB�u��c���z0t�v�c�BN� F'S�f0)pDR�CAv8�$uu\r�X��c�����J��U-��j��d�3@�2�#q�����/\����n:���� J�'\1<���s%�q0�d��K��6��ָxfdח@�4!����vd�^��`X��)O%�UV�QM�m�0�K�r��a(J��M�.q۶�������fA�9Kr����m�֎�u��1a���2�IC�	�Z<<�7:�h��ذ�8L-Ü����Bg]�,��F�Zi������k��%��+�>Vͭ�*�g�<�Ka�0R�7]9Nn^�&��m׳h!؛�A	��t@�����W�Ķ8e��0]�����2X�,Iq�f�`�M�:H.ۣtq�d)�+����sd28^N�u�`Flm'='gŝ��W��.����v79�A�qg+£�=V�$�6��lnn�6j�X3WK��P�)�qf��2�2r��40@�����rT%��;��gW;��æ.M�u����'A��%�/4���qj]ez\m�uj:�� �]n�NI�Yf�5%��Жۛ�H^d�b�q�t:9Ni��'J�qrv�\���$v�kv.�ݔք�/3!e0�ʑe.n�n�i���@ ͪ�kJ#�2T+�][��s+�хĹH0y�4!`��yۍ�h���^��M�\8Uz�3�]u�f���1FĒg��z�;��'G%*m�Ʋ�Q-^Ii��[��K#�m��%�.Ι��껭�n�*�ra�s]�vn�v�6�=�UvǓ,m��/Mp֞p.�˺+z��Ѷ�.'g��u�u������L�GJ�U��]�vm��>.kpu��HZՋ��e{-͝��u��p��W����ȴV�����w�����H�`�Xld��m�I�]�ì�[�$��N�[���\�b��[]�Q��m�1��0fj���h���ܚ���"���f:�JT��g���pg�}��f8�r`�z��>�h��"^����ޮ�_"kI���<;Gj���j��(L�����5 �����`,�i-H�f4�reW���X�).ؠ9�-~K?��r܊�N"-��]�En9Ʈ`ە	��s��U�ffz[� �j�}�&�?��J�]x��d�b\F8�3ݫ��=G�Yo�ۘ�TM۱wl�;�'�t}5W���[#�dN��o�.2��ѱ�Ğ �v� A} a�y�y������~��� �TMڛ�~��*!/�-��oW���b�ëӊ�ʞo�}>�ݬ��2&���V����RS+(W���W��Z}ҏ�H;µ���q���ڃ҉��1�Rn�b�혉���s���I%��>WN�F{�
-=�\��D�_#�a��n�Ɗ��ё9�M'�ڃyz��{㮱�,ĮwZ�dn�n^۲�3%0�N�y�_�C�T�Y�m��A�5j&D��ëӊ������p�z�ណ޻����=�Z;��D�S�V�ev���w�n%�[��+bsF#�1wh���3�7~�׻��qۑfzY��Jɣj. ����4����݉1���٤G�ϧ���@!}�8�j1��Ya�����¿e��Z�ȴ�~:@�����+�����8���	Ͳ�{�,�fԧv�E��=����t���Ji����J��F=�����`��1ݲ㻷�����T��A�#}�H �
�����6+;\Z�k����jv��`�؋��~�#ϷZDwj^��5�������Ǯ� _{�z�J3�N�w��"> ���� ���\;=Y�\�7�?;��kQ�
���A:,��K��3��lh�8ˎ{e��eu�U���t�7�bq�;��Sn�*}��Ji���%z��K%����jĨD� � ?����@?Q6� ut��a��RA�������lVg3j���'�3!ƪQ����Ô�|C0Ar3wp5�ݳ�iW���w־���y�~�B ���W��|N߭���q�Ll�yP�7P�tfOVTKu��.��=X�LT�e�Dc����/�Of!  �Ү��y^�����K���#9s1O��"�_/�n����<�Q܆�E�]
m�eB��~%czmr�J��z}��R��V�k� # �wF� �l����8�u=`�Ģ <o`��5ٱ����\�BH#�ȟ�9�#��9��ަ�X�`�)(	E(S*Q�s��q���Q�C�֜d&-Ƭ�h�ݬ���o�A7Ј}�H#�bmxޏ+�{�N�w�]�^�N#-TVi�I/�Zv�wl�f{��+���=��̤F�!=�{:��2��gG
�8@ �����df�}��iZ�;䳼�Ǽ�Ȋa�3G3�Agd���y'D���7�E��O��k�wX(|<(��С�o+>2i䦐VN�.����D��#㘃���r���/Y9��"�y��t\s�{^���6��s0�/�1	�]��E���u�M�B��*f�DX+/F�X3����#]
Kno�+���%fJ��gv��;9��|> s{���u��dwv��n׭��>W3���ز��\���Jƶ�R�[���� ���2��� (���ZW���1I#[)�9�<t��ݳm��-��J���&ƤɋkB��2��3�6��zЉݹ��=��Z�d\�o8[~�s(o���bJ��e_v���pw�b&���(Gv�;y���lfF��!����W���W��|{ή���"&����ݾ;��g�M��tN4���y�`��P;�/w$2��a+�N�������b��>yV����3h*;�\wv�Ok��{���c�W�}ׂ����L��i���������*r�L���Q=�Z'�sjP�����0f׽���L���������GL�-/Y9����g �f/���V:�.֕Xaq���!�H��Y��9IbEN�b�����ڽ��pӝ{3��̇Yy���zv��I���a��pk�7Ó8���wt�O�}��i�A�Hra�푆槴�h�H�p���6����}�m�.���2ݴj�:Q$��9�6��vOd������A 6vY�G]3��t�kۋ�ng�K��8���6��u��Td)��uV�]�` �L�-�䁲܉�"���Cj������fB5��M��%�{�RT��[��nذ�7 �Tƫeځ�~����E�Π.NE�Tb[/j���v竞�*��6o�u���>@��В,���B �d�7�/���]%�/C�w�9�.�jO\a]d�2����-�ۘ&��G,�s������yp��Fɹ28�o��lwX(6h%��+�j���Q�����2~�:2�����ꙍܯR��^�ϓZ~�����Dքݻ,�YN{��w}A�����p�7��3$x'3�z5�r��տ}G���}�ט�V�ͪ�ʛ�~�SZ�;�X����z�����=B�`+��ߦC��=������Y�2>�̟�-��
;����
���wE�R*�q�z�;j����#nb�e����/҄~ږo�������F󞎙�Z8^�r-/����*�u�G�e�{˘&�w%�;�a~n�T��9׽U����%g�7pǍ,�t�t��Ԥ�[ک��2�$��PU��y'�����g�
��FM�W
���St��M-�� >��x�@@��/6{�F�e�c/G
���Α'�m\7u'sW� �.�H �0��w�LiU�{�eڦ�/����}������b�ͳ#:�;�h�fH�~��wZ�.i⃛����|�F�A��~p#�bX�烦s�/Y9�0�����*:f��w) q�3�bA��s#�eCf�ʭ�dOF���FҬN^��t]BΑ ����m�þ�n��'xW�N^Rڷ�t�!��-����X����<n\�j�]���_����i��㻷���_��Z�s9]���Ġk�=w�ilUM*�Ζ���c�Q�զ��7��ڴ�+��Y�V����R���ν����S�e]�������#���y�z��{̱���6~ϩ���_�#:�E���T+�
�g�Tu��T�Ƞ�6c��A���a�ݚU��7�\.���mf�o�*R.�V)�D�������<�-���q��z����ݦ�~���'���۴>#�Zu8,�錡B����Կ�S��ːzB�/pۡ��c��{��W�2�}0�
�ϩ���b�o>��F����̧�xR�zPCc��:g-h���]�n�ɭ;��ݼ��k�7��{����d�8��hec2��u��bͮpm]�P˴����h\U�fItfԵ#�����^���_�m���ʁ9��]�R�p1?G@�\=k>��s[n$~��'��D|s@�b�H��S�nk���a|1�υ^Ҍ� �<^�C}��|�ٌ�7h�x��پ��t�s�C�U���c6�3v��/9Y�+e���~�N�m{ç���m�Ȧ�~�㻷2#��4�Nh�b�-[5��_ �C��
6�[�ވ���0I�>>��i����y���j!�����% +b��Z�h5�ne��e%үB:!��ز�h��σ[�,�����u*ot[Z�)R2��h�,j����<���G�k_6�|(P�>l�|wVY���s;3��fs�&�݋ɾf�5����h���(6�ߗ��f���!���"�#��vr���� �?ޯ0��;�e�{a����NSS���U�~��23YF���{�?f2�˻����G��t���=yr��~̟�'3�91TŘT��o�lP��++Ź��<�؄���������Α ���1Z�G]�ܠY��ob|�&�ݼ���_k�}�2/�-h6�3�v�굖٤��sl�=Jڱ���{��_�{x]
����?�wWXy3�<7S�H��b\$a��!ȸd��s��C|߯�&�Mݳ؈�Twj������r��V}^3������BA<d��S�*��~�mFn���~�n�oI�U��=����?2�:b�ڗ�Rͥ>0��׌��]`�¬�X�*Q��	�7ev����������i�y��H@��}��5WM]V9�w؛���j-Ͷ�Ihir-��kǭY뛺C�'��a&R��֝�/��x1��F䖻��7n��Ư�����N����E˷#X!{���mw6h:�=c�����ҽ�Lj�l��+�\�ɋ�Y�-Dq�zf�7c1�v���v6�N�;�������vv�r4�L��T*u�w1�2;��[�#kB[���;��Z��\\�?������!�u��v�[�ێu�zv��5GN���D�򩮴S�&h��

@��ͻ�P�Z^`̹8������-j��q�HP�p���6)�u�>b�lأI�3dg}�wk�|z]^&{���*x	8�]�ޡL)���n���vR؇�JZNmػ��GR�v�Fn�7�l��cz-��^��UZ7Np��uBVr�a��b�3�路��J ƤAa]�1��{TnMg3R������ǻxNHX�N�>3F����ϩ��G��+��<k���t��eO'i�ۿ�15��Yq���5h����o���߿^�뼊�����5I��m��G9�z� <
\p9�A��UC�������<q���z�̈9��9�"A�����Uh�9�~\
�9�ﻎA0�Y����76�P�B�4>���)N�u��}�����A@$�v����ɚ3n���$�X}t�
��K�D���a�C]��q��,��qv�K������|��ǊA�
��cen��ܪ�3T��v�|~g�e{(�j������wL���@>7��������^�r��e��-��T��;N����Mi��wv�	�&�!MÌ6��ő ۄFf! �n�V��r��h��?O�f�q�"u��n[�Rg��Vw�B���M�ͻ{���aޡ�i��=��c�fv��U������0F�ڱ��}^�ư����Go���p�u845���T����V��t�m]u�s�֢2�kS1�������,��|�_���wX9?_?�T�$�w~�Z�Ԫus
�eX���6�0��f$m�`�߮+y��G���
�3�9=�q�Yy��G՟g��7���3�1;ƻ�;�X���C���n��#^p���:�U�
��Vm��sP���lup�=;Y��p��;�.GMV�<��}�eru�ҭ�Ii{H�"Mՠ4k���ë�^5���A��LҴ�b�Egg��*K�DT��c��+�>��)���	Ч�7/N�h�4khz�R;B�gR��|�6�H;�iJ��3�[���m�su���64�W�{ռd�[��T�M����lvbY�]�1�j�߳�]۸)���̭PG`G�]mw5u�^t��C���Zr��a�2��Q�r���ձ�����BuH`��X��$������k;!�w�Yð���|�bb\�[� �<i0\�9����qc��:���ݧY|��.��W\���l�ɣ�5;���3��.hZ�j��v'e�uܷ�,�v�AO���2qG0v�Oj�����3X�aK��ʴ�f���ؾ��i�bG��\�R4ѱ7f�n[V��[���E��AMl;;���	x��˾i���}���<���k�����q������:��q�QԺpfCKmv�2���ܫ	[.0�%�Ud�l���[W���!t�?+��9ӎ���Oşjõ/3�ݚ߆�3����:�}#������[f����I�u���f��|�\P2�w��v�B�@�SL��E��w7p��v����U@�ϓ4[�V���\�ˏ�][)���������Ǘ�:�`-AJs�u��o] ��y/h]��dc�.�qi�YM�A�֔��,ZfX:�j,�����1j�J1R"Z�e`�B(m9[Y�w�y�s|�iU�L�TE@F�-)/:ޖ�%��Q���F�[L�5�b��5\3�G3`���9�O;NՕ���޵���s��-&�:������8�34�*8�S�t6�]X�fʱ���6sg��fq��Wg�;zѰ3;�㢜f�9�Mvs68�f�39'a�� `�YQ��֭pS]vl3��c78Ø���3i�V��.`sj�a���w3K1:��θ�n����30��ُX��b�`l���kU�9���VU�޵�ه9����+P�s3c3��0+M��gc�CVф"]R,�)a�O=��e���o�}�מ~,A�v��n�"n�3h*r��ſN�Z��O|��9AQ7P��9<�u�z��pr1. ���V��7�~������&�؎�ق#�N��M�pFĭ�)�`�'��αY͐�'�� z�EoO�*>#1�u�{���z�_m��dt��v���8��:��6�]�2�%Qr�f��f��9w����@h	ƛv��J0f[���=��~����������uU��*�w�g��<ι�ý�k�ύF~��}}<��������������Й��GT�����32 ]k���)�M��s�7X���B?U窽�=�٪l�۷�xQ�Ql�Tݥ���T��=�$.������wqƦ\�R'n�nj��nC��qʳ&�.M�J�f��Ňf@7X$���ڬ�z1X*=VT#�M�:XšY>�  ���{Z���6~m��#�W�S�c�}~��~~Y�������Tۺl���饗����vծ���]i�4�nڻb����(Om���N�*����^��V.��7�6�nw�LcÛ%	�^z��jm%�Ë�����l�6��l���8�9��H���_N5iF�s�\Ǟ�r��X�Ӆ�cf�]\[�g��M�l�w��-{��)K�k1�T�@G�Q���M���6k��N�z��={���nڎt�6-�͒��=�{Ma2�r�p����n�?Sm��.s�'$�9�\Ǿ|r���5S��?6Ҿ���hf�����:�`���ǥx��}&����^ďO�+~�"JS5[�-ٓf)Ð�'�*��*�~�����<����OZ8}������s	�m΃m��������h��: X3��{v�puǮzk���/H6:�	-��x�n9:1��u#���[�{��Y�k����k�۴�6�4q���0��k��38���%۞q���3���O�{E���e��g����s����sk��p6x�I�W؎�:��n,���s�hx�vYM�C{c� ��v稗��ڡ�}��3�h9��=�K�s�n�|��p�Q�V<��BQ��1&n����z�w��~�~ϯ�zo�J~�8���<��m[���[C2>́�f ʫ�5u042�oo6ż9�T>���~���//%h���u����e�Sx�x�vW��{�YG9�K����Ս[��5M�n��_Rd�K�Ծ�d)�퇴z�tg��w�:��_=Hs�L�����g�ݶi�S��J��r�o����+&Un��������Y�b��X�s��a|zD�$�',�ձt�۫�&���%�2zmΎ��P�=��[���~y�2ۺlե�8�������\0U�U�|ۑ����24r���T���k�n���u�t��nT����}��6=�w|]ʥ&���\�+orh�N�0��;�mn�G�bŕ��!�aO�N�ե1�� >Uw��7o���N�����݀3�2�_l���Mi�4����m���M4t��b����/d�}�}�5Z�m��l�n�Uw"�t�|у)��lդ���ͼ�̄�����TL�D�����_fG͚��m�{o��h���/'��,g�J�qUH~~4ۿ���x���Kxv�ྡM4��It�k��C��3�$��3�ׅ7e�^�Za0�H�31�;q}��d��f/�;7���X�Vi;�T���V��3��H[����3pN�=to��[6��xը�0��Cs=�ʿ}�_�7�}�y���;(PŽ����6�ڦ��~ݹV�lh� g�����O:��8�"c5����Ҧ��c:V���6�-Cӏp-�O�.
������t��\!*!1v_������7gp�����"�?��5O�n�o<|��u��i�Oƽ�M��\s������'�����^�2_��_ש�� y=�S��o[4�Ru��r�K�̟���_��G��[��۞�v�6�z�E����{kj�R�T����T���͎�]J�ځ�����W�����?fk�t9��4y���O�]������?l������r���l�з��W�_V��_���F�)�'���{M5���B�NY]Y�6S��{s��6[w�c}��c���'�F�ܿE�2�����ʦݶ|R��v�b��?}z����f��t9��4����O��?m�5\��.J����[u����͹N4RfX���,�!�sN�L![;G�Z6eA�C'�QUb�1DÝ�N�jf\˙���Q�GV�������b�3#ᙈf@���]:��>YK�<���Jxu�'���W��Ms{M�Ꮪ�^�F�OhŲ���tyBlۨ��c<V��WM��(�0��*BFT��P�"R�L����̯� +�dÞ���.��}U���:�fN?(~m�Sg�n�R���iu�����?f���w/�i�q�}!����~�<�c�5�V3K���g�����⺮)�9�~}��\y��}�4�[f�-���Х�&�>�}���=�٫^L�s����{R#�U��7:�Q�7�r>��2>��8���d��1�M�lT����8O��4��ۺn���� m�y�7�f�k����S�/Y�z?D���>/�=7r�:��=���:��{jv���)�ϭ�BS�{o}��f_��;������Ŭ+�u�͗���N8�L���u���:^�9��m��p��0ּ���ΧMhÎ+5�.�{�j�ݨ-�=��w���麎t!��v�7\�L:�'<�L��x+�Кۮ���f�M�f�a,��eʲ�FQ�usyd�)��Tu�j����z,�#l9$���Ş۪�ݞ�Q��ʎ5�(��]r�G��ɡY11������ߑ����Z�*�
��O�Z�v뙬�n �J�a6�в����?��=�>|9��n��������U窹tE~�U����e�uM�YJPB�,���M��?�ɓj��ݓ�YG�ҿ�q�c���Te����\���{Tسp�e����M]��7/\��2p�}����6[;�Sڻq�!��-5�j�hS���ǰg&+4��
x�����I=*���2��l�6[e�_ަ)��l�y>,��)�}�9Ŕ}�]|�y�6�J莬�T]R�G"$D�%"dIRfa9]U����X�5q���멬ah�]+��u�?�I��?�K��Sy�t�7/_�c' ��p��e<�'��w]6[?6�A���>��Y���+��t��
0�Wg)�˫�b�bn[U�B�}���v��@ڽzb�������[H˨-�U�}�ﲽ� 7�
�����������W���m]�yZ��	?_+��l����^��щ4��;0Ľ�}�9Ŕ}��8�6��m�b���=[�Uv+���ėG�Yz���2pIW޵t�~`���۪��j�w�e���J��Ĥ����R��U��־��5M�=�����ƶ���u�n���QZ�t\�\s��6�<���]mph]�V`�"��5^f�w_6~^i�����ݓ�YEtq�s{/:�^-�}��Fj�wM��?9:�vvx����/Z�G�������>�C�>?6�5�"F�x��j���uM��;5�'��W��i
�=�N���jNYc+�w:�b/�ıH�x�l]ң#��2Tq�G"�Kq/�s��``�}y
�
�Q1!Z���}m����| �mm7���e#���9��#Z����-��g��[����Sf�J"�%;�Nqe}U�e�����h�}�?Uw��g��Sn��&�
>m��꧍8��^���8���soi�31�甂�"��ݍ.�V�'�Z��톞:����5�zx���GںY���{�S��\�|ۺ��s�\:SۅJܜ"{#�NT�qC�}n�d�̯�v���T�]z��=�vI�"�>�����4ڭ��}x˚�g�����m���7�vȯ^�1��O-̗�p�T��ͽ��͔p^k�N�YS�����u��Kb�T�<\�k�*X˓n�x��n�(�mn1�47aQwC���&��F�b��M,]]��5v͹��i���#0�����_�$��]g����Ĺ����������-V�鯖�H`��|9�"T}U�_��l����NՅ:sH6I"7J�P��%12�l�-C��hJ�n�Ck���ae�֦c��}~��gO~�[f�4�W��<��3��,z��/}w]s��@ffO�3�bX�ki�̳J�� ��+�5���el�h��<\
ƾ��{�o�[2�#^���5M���6*�<�:gү��Y��ǝΑ*>�J��ϛv�.Q����O~Y��j�+5z>����{� g�8j�{2� }�q[��٘��̉��w-���V���7�+f+EV���:��Ƴ#3���k�Q�9����2���j+H�x3kG�?�:ѕ�� ��̖^�Q'�������&5]d���[,�����h]�[	�5�����Wi��*�QN}�5
M�;�X��;|{QH.�c�lڙ��U����'y�1�|9�!��Ot{�=��k�����t^����J+��W�R僶N�V2�n��M�T����e�1sB5��),�N���3*m��]���儫/������'3V���q7R>�;+k{o�8;k<U~x�1�JWlU�+����T��x��\w�u�}�{2d�I�j*K
�.��[�^e�E����fone�le]��S��%��5�Y�jre��'32�Jl�T��[R��#j�I oFcp�W'l�m�d�9�9�nj�kX5���
����R�t
㷃�e n֣����n���,��������
*Z���ڤkY��+z��2vb�?�=���ڎ�Pb�+���Hd�t�i��P	�T��}���ˮ�$N^�7��ֻNU�s�v�[��e=u5�)nF��ܣ�h�Z���$��!�5;�|Oe<�7-��@v��	����x�ã{�8�ne�ÆC+k2��6.|��}g�*΅�:��joL�/.���(�^�u3(�qV#�iqQ�GZ��|��Y�Z���9�0�"�b̧{i��웕9����4�i}�3�$_�W�_alf��kPaG32�v�ά!R�NT� ��Ǝ�
b�r|��wt0�Qڭ��s�^|���LP����V2\,2(�t(�N��+c:#�K�{/3~ӹ�����\¯ŧz�Z��3vvm�ڸ�6�f=FV�����ٜ�g1��k��{׸͛07��_:3�Y��ٞ��ꦛcqŚ1��u�&�pg:t�N���l�[����`s�Fc�����z�IX�=Y��6�\����a����0�Y�	t�g6��k5U��YV;�y���1��6�� �,cj�������n�����z���c��羮����=L�=�ɞhٰ�Ů��WU�nu\3��6������Y_zo,�m,�ٰW���4��L�cf�d�z��1�W|�g��ZL��ׯme�%�[�X�2Y��z^�]`S���,;{�l��3z�����:�N-,%��m`�J�In�$.�>���`�hmt��t�j�$3]ŭ��S�M�g�(wF�,�$g��'��ݏ.�=�c�����kO�'�k��.��������fۮ�րy�Z�A�k<��q�l��	'�Vޓi3m����(�<ݮEٳ�zSv���hpν���Uj`��5��v��M�au8Ce�R��nkTJ��+ٻY�������al��PwZ��ƠFisdT��)usu�bۨf��M����ln玶��/o������D�6�A��XXwI
|'6plm���y�뷱jC����X����5���9Y-�wkB�s�X�A����z	խ�s���]%zr�%ս��@�n���1v20v�hq�5
*�ƙ-qr	Oi�;[�j��[v�i\]��n:	��2�����	X�z�Jn�-�j����C��Hz�������=���*�K���L�s�%����m�a(��y�+��wM-�w��u��gehM���h�$ݺxW]=��s���n��j�4jm����T铫���m����y̙�'��p���C��ͱsН�<�R���f����Z�v8���ص�ͼ2�7l�,1\+J����.�K4W��0�k����W<ITfa�1j�4%L�]q3e
�tne�<u�x�gr�ԅ�]e{Ml�E���nêB�[m�B�7CB�аcM#2A�;��`xr�F���Kf��5���>>2���r�܌Ȇ�{]����'m��R.��̻5\ <Q�K���Ӡ��ң�;��t�p�V 8�+�i��EK�b�)K�k�9(�%*�!+��6�6�ceyt;s��Eh��5�W��hζMع�h�!t���]�͚6:�Ee�M5FbQ�Q�Ў����mv�,��-W5cK�A�i���k)�ҔFv���{4R@��M>���ol���)l\���#�,��k'9&u2���Н��1ۍF��:]���N�T�A�sb�i��;m�j�q�D����λm���$��0P�c=��'����Ԋ���݉��$���ˡ��޷G���؞(��M=xxsW	�i�Ř�뭎��9����e��;� 2d��NN���.��������m��'=�H�5��nz<���E���|sɸ����UU51)��j8t#
2��l�c���ܑ=�WNZ]�v���R;b�����mlE��v����	|�����~�6T�+�S��]MSWS\�ڗj��Z:��t*����EJR�1����l|5�f,ʱ�����ft�Q������rJ�q�Rn�?Sx��{��qKͪ���+5H�O-ߌ��8 ϩ��M�?s�gQ�}�Fi����|�LyT�U2y�f׆��S�J*Ȇl��W��q���6�p^]�]�\�|��ISf�R��)Y�ft�Q�jW��	̮~���V�4��ߛ4ۺn1��_���N?R�w�=a� 3�ϋn�Be�}������:�K)���&c �M�7Wl�4e�$�PQ�,�U�Z�K��i�T�����I)5Y͝W��s��u:v4�����ų�f/�d�O�UƠ�P�]�1��4Q����4��q�� ��"nV�w]p��#��k'xw��
��Tk��u�͊��慟�}����Mb�Vj��Dމ~�ov�Gwk�p3*)]B��ݧ���n�-�En'�zɽk�����zÜ e?S�M���M�ћ^�}���O7{�n�ɍ;l*�ꀵ�Hez{u���5O�6���6��1�~��vi�Wx╝�{�J�����M���N5CO����F��a�yuv�5U�l�F�����{�Mpab�%�(��lf�k�n�D�(j��t�����\�R�w��Xs���\q�!k���5���6[?6���n�7�I׉͎N��Z��YU����l;Ӵ�^?~��_��-���������_Tm'�0�b%�R�z�>����ɦ7N�24�taP�f�E�~(q��rܗ���4��TJ$�KK܈�bn��ͤ�2ґ�m7����5�5�އ]�^m�^�e�f@��k���\��u��٫Z�ϊ�w�=a� 3�p�����!w��+��m����|����v�vwu�݋��ѳ�®�{Oի����Jyh�߷v]X'�ˬ̠b	5���t5u�s�@�<Wn�:{V�u۬n��8E��?s?6���j�'R�|�D�=Ws��Zյ�陏����{�e�.��Or��w�j��x��S� g�N��n� �ͷ�0�0�wT�y�nx{��G�zM���rּ�5�y�i�W7�6[w��Cݳ�����+޺�Ρ���š�c�{v'�v'$_]��X��P�kD�p�^=έ�5�Y%�2�y_{�b]�܎3jv�ޞ���p-"����+c(�n��}��c�ý��a�l�6��c��_鎪3S�n?x��S� g�N��n�<����=�����p���qUWl�|WZ�#��GO ��nml�!J�?L��v�љ��vn�]���s1�Va�u�i�$��M���Q�sy���W����VkFo)��ۉV{��>-�c��� ڿ+�>f�v٪n��6ָ�+}#+1߈�Np ?|��|[wM��e�y*f3^�Q�Sf��1
y��춦�ob�8J���)uƍ�����|k�m�Sg�l���L�C3u��9-���;��y꿟l���Pj�����Yyd�t����y�oK�l�(�0Wt�3k��S8��I1i�8Ă�&N`X��-��-Cs%�n���А�����۴h�̺K�4�Xۨ��1� �e{r�N��xl�#�� ˅��n4�ջ��ݝ��%��훒�  Q�5�^)�%�2Y���Z�TRf��`%�ݽ���fx�xn��n���6�[���v��ʷH�{gt�n��]ڒ���cXEm�z�F�ɹ��N�TF5�N�evz��l\�'��#L�O1�7a�~�g}�~?��N��W2��9��ت�5��G-��VK:�Q��0Y��4�o[5kWy���~"z��>���eN=��xk}-��wf�W��a.�5�^�I�HN�N!7�o�����of]Mp����T�٦��}To�E�\�%W{w=RGnE��ҿ�-���m�T��R4윮��ߝ�5�ِ��cV�߈��8 ϾP���^��]��򿧈̀31��n�K��b��f��tu�n!3_�s��:����g�>�,��ؙs�Ym�I����nmbf�z�م2�`9w��ߖ��Ƨ�wM�Ze9�u���ηT'��J���fxvkϤ��g��S+��{��=�'�J�N��U�˪���[˞b��:���l���-�>�˙��W�v�$�L�rb�j���F�����w�oE�^��W��Q��8 ϩ3Oͻ ����ŇVN4�_͟�5M��~bN�W�}tKyY�v��T�8�hf@�31	��;�؁t9���ր̫��5����n�O�_g���=��s_fG�2>�Řf��;�۹x*3����yۜ�N.��C>���~?Sn���Y�{ٝ�h�n��4�1Kv��]���Fc�K�j���/!��n((���U���؝��?6�\���	�\�7W�s�S�
Ԧ�|�>�9���l�n�J���(��P֨���WE铻v��TJ��o>��.B}�*�ZF��m��تsP�m���v�o���.ŉ٤�PYl��Ae�M憲���n���w�磮�t�+
�z�]d�NͅK�s�>��]��4Îx������I�W��G�s� g����?�wM��15!��s��s=ͻ�_I�-s�+f��,���4�sE�'�t5U̶�ڦ�nʜ������۔���y}���	�TJ���|ۧ�]ճ�x=�R�aó��;M�7���[�L�Γ��nv��˱����`l�A<�w�F����;������p9�-�z���Y5Գ����C0��odl�O�����5[;\����\�wWVg�����˔�Ϻ�n]�S���}�3#3�<�rmS��۹a幓�v���>-��w�g�A˺��i�k�����?^>~�q߈�s�'ղ�FV-U�x�SPtVȳ<(�ˈ6�r08��9�i�El�mҩ�wj�E�_^�hgf��mj<��v��o׉��Qu����T�2*����}��5|=����d�����ܫ������&K՗�ƒ��~w���'�_Uo����>��5���6��CWf�@q�V��c�j�e�	��p��;<��e�t��i�NKes�;��{�o��xb�F�<��{33(f@E)S��4���y�f�qt5��+s�fc���Mʡ�nU,���T�l���odY�*�ֶ-:5&�K�/�^���Kl�6j�v�X|t��~=Ϋp�z�5��y<����2w%Y�د�O�*l��ו��8�\��٪l��nF�y��l������ӎ�G���>�~�C�6���̜��q�ćq��YJ�w�[0֭�$=l]6�4���"�Ό�%Ԕp�%�ܣq*�&�v��+(8��X�������M_�W�d�l��4��v�Vz��.:�gd�0��]��7`�q[k�(wnz:���B[�m�q�������m����_�0�����h�k{k���� g�],$��\��KL����G�hM[�CY����c�	�Â�f�Kw6��g0nr�i�`�: ]u�,JQS�2D�h�lD���{����[�2ܢ.R]���wYf�K�#�<�g��l۝gs����~������~������yh�<ܚm�V_�C�}׀u�R�3�V��� ́��ν�\n��j���	WlO2r[)w��ܖlW���7�s7��P˨�([v٦���0;·���K�0�R��2}�d?W�oi�M�����%o�����m�c�w��3�7j�	\ �i��KVbY��=���6i�T�����<p0�٥��f{��K�$��{��ϊg�m�#�j������Ë}�4úڲŘ�&F욁ؚ��ֵN}���9f�#0����U�z��6j����^.�kh�v��oY'#��܉{2b'�[@6~l�ۿ��o�}�:�Cv�x�x�fN�S�O��FZ�&�ES@��xx��0J��s�l�z�{C/p$��Ig]�D�s�W_��}��^5_�j^��,�\nA�Q�w�Tn����i��k⦟���Wq��ͻ���?R�Y�b��}y�K�zI��V��%t4����m�d��3E�2����&�scjtLg�oY'#'Z�Z�nLZ�%��~l���t��:O�$�b��ޞ��`3��m��;��Z��6~��M��ɘ��Z"��\i@0�k����c\ݽ3but]���jQ�T�2�"R���� fb2�\<�K�_zI��V��閨4���8���ͻ��Sg^���ck���@.�\�Ϗً�u�w��N 3ꩥx��˞�p��"6�Q3���3 fg�
u�X��(b�D��j�ft����+c4��7���\��̧j����Xi"ޝ���pE��L"0_V7vjf������]i�oM�';����t�;V6�ls%��68���xi,{Xc�Vxȩqz������<����:X�Ǫ�rfu���|i��׿i�����xoo87K-[.�t7�fs�s�:V01Ӆַiѓ;,}�$:��}z��t/��(�+�Y����zI®�DO�o�А*eD�� %Q�����ʍs7M��vN̻q�v�ze
[0�x�r=���gG\��G��.�La��}��J��e�S�l"�7(f�K�c+����j웝�����,ѽc�3#/e�ñ��Cʕ�Ee¦dU�&��,��\3�@}ʯ��ٕt�4����g�q]ͨ.#�l�$`����R�؉̾�h�7]̚�tٵ!$�Ղ��v+tsY�A�ґ�1m�	[{�#�?6P�n�vk������X�PZ�:r��t�&��xA�ңH�&"����k�;��S3)�Ds:^
�ZZ�u�
�X-G��M��E^ʼ,ή�����#y�eu)r젛�1�بc����X�*������iJiDxoH�T7*�eS�a��ȡ$U�kT�i֋"6K��o�[�(]�rB��i�������G��zM>�[�+(b������c�V�ķw��#[��S4V���]�Tsj�V���3��o6���>͛32���&&�ȏ���b�P���dk�C~+;�;cW{{i�9�s�i���2z�o��-z���f�V�L�{\�c3��xvzם�k׈��X�A/�%��am����	,���z�'ޠ։d/B�@��RY\����͝喴7��}OT�x���[z�eB4���Ṽ�;�]|�=�'���א6q�X:��z��Zί=d���ǫ�֌3��zm��7��Y��޻+=���ٌ�6g_{o}Lc��,b�������{1��35�{/��'}�x�u�q��Ι��Yެ�m5�g���N����e\�o�fm���G3y���,�z��c*Ӣr�� U�Z�:3�[�ѷ����3{�b��G��}���z5�sr����V�t٦�ͻ\f�����)�����/']�X�we��\ݡRހf[�����ݷ���8ӳ�XD�2}份y*���Y��^{��M�l�|\��>��g�]-�.t�XP݅Imq��Y葷���j�d(x
�v�?�yW�o��K|[?|۽JN����	S����cЦ��k����UT�����x�mK��5��'�����}�&w%��Q+��r������<&fw�u��%Ԓ��U������oU�����N 3�W�d�_G.������u�;�u�r��j���5��Y��p���w=_w8�S�ae�պ�A�|�j��gÈr��i��F�G�`�YZ�;��63*��AI���gC.�7�;:��ɖ8W>��{���2�n�Ӕ{�}\{�ܝ׼jII.CRA5��[�A?���7����}�&w%[�_��M��z�'R{J�ٶx�^�/b])e�DZ������/����u�z��K�[�MQ��P�f��v��[�3����Q~5���>����Ñ�ԣ����~�%ԇ��@I�j*���u��u�}��D��ؕ��n羮✺�y�5�r�Z�Y�߮������H}(��$7�c��k�$��}Q+��r��]I��f&�U4i�}M��Pݙ���	_SF�q�}6]Z{F�f�&�Wu��R� 7wvss59#�_u>�Ԅ�9�4Vts��~N\�ꤌP7Oei����x��n�z�3BoK��b�ц���ư'Nh���y��jF7-��:�{K����ک�h��{{�Y�������O'���Ӏ^Ê��K��Q���^�md��^zʌ��5n�n��7o-dc÷�cCb�ax�ʽy��εo I�`s)�i���� �;�����-�zh�B�%�a^a\��I��kdj�]r��K��.4�`:{k�S�:u8�Y;4u�:Mv�q����V��օW[��y�^S�Lt<F��]r�'na�;*�ֶ4������>���i����IQ��(i��X<�]26�@�!��&�hfݱ��������6��]y�f{�J��q�rU����}�J�5?
�C� ��7uط`�[��r��|�[�ӗ�(��z�}�}Se����%�}7�ת�8��"�C�I:跕	��<��)�Y�ct�o�+s��qN_�K��/���,�I}�H��_�K��C3�JV��;����/ol��!<�ۮf�Iu$��}$����͈���c����L��NtB��X�rr#��Z����wDo79k�Y���ZJ���υ68*k]�d��Ig�R8�t�s��L0����[��]7�􆤗����˯oct�8Vd��_^!=�W.���=@n����<�ٌ��K��4�u�n����{�q��Kh�n��B�c���3&�� U\�M^6�ol�M;��{���0/Y���nè���}�����;>�5ޑ�r��}���O�L���?��b�T��Iu!��v�<�ԏ=v����[�����E/�~2K��\�������jQ9PF�H�hpx��9�f�=�3����:N{Cb�6���%�I$�:��}[]�;�����_S�;/��e���n�W
v��/�cỼ�:�ʋ��>" ��t��������u�U����ؗE.�	�s6�Y�+7=%~�>O�S�IuR�"r����,�vO���-T�xy����RK��RK���n�}J����uCr���k*��9�f��k3�w7$�t续e\��Z��)���%ԐK#��t�Z�k���Ϡݗڌ�=�ԃk^*a�B�*R�� z���us2K|-��%��m�;_��*�]�2-�����R�}�/ݷ��ȯv������75 �Gt�� ��c��6�aN^jOAW/�5.I���O�E����ז�5u�ܹ}$��Iu&6��Ü`�!]�������5Z���}$U&�{�T=��v٣v�(�҅5"��[M	���5M�s��m�KX�XcSm/��o��<jIT���3�\�]�w,���>�{��}�[�e׼j��$����)�<�$n��S����U��K�r;�u 1���b�����whf@��n�*��e	�b��|��̱9�q�S�k�Ɔ`n��Z��5��/�������pL��0��,��u���S���۳��n����w�����ZA��.�dd6N=��T�݉!����y�z�̼X����x�|�����������ʒ�sp��
��d}�����@��|AmȒ�_��po�W�|� kcw�����~�j\���Ŷ������Ԃm�<���]��g�ED�$�`J��ZD�;s^.BѰ\:Jn���k[�9�����@�Y��~�����܉�/7���U߅f��^ʥ�=���<�:�H �9�_�|A�@ۙ�[hI��{^�}�Yb�׊Ao��z�~��9۞���x��b�Fo���]���#wû�3�EP�$?]I2����!��ܧ��/&�.�W����q�r|#W��@H�A�_KnD�Ck�!.�n8xr>��3�Ϲ�� �t�����6�H����7w�^l�d������}�p#1�hg�<$�jH'��s �m	 ��@��fI>�r��؆�˼^�/��޾Ý��n���/�1}�h`!��-���+���Zw������Q7&�d�k��RJb���ʽ��NFy��hPrw�9PR�ʇ!�p^q��Q�����u4�v����}2T�RPH@�c�)R�c*V�L�cn��#���nv{Mv�h��Ԉg���VtL:�N����L����s�����D�X�S0:��ö��^5�r=���k��UI���=�S�ʖ��ؚvT&�j@	�sjd�a3��봬��V�,(.U�uIT
�
�
&�M�t-u��8�]�As�#��Y��Kg��U�{u�ޮ���|�@_Ͽ��n�z� q����G��Ϝ�(��<\2srE�u���uɘ�RJ�J���|��?ڐA �M^�̛Sߧ�'�1xH�Ud�xz柝ǐ�#��$܀݄	m�""����D�f���r'�ޏywFfX�6mϲixA}��BKmD�[�_�&A�B@ ��m�܈�r��OQ�6��m��[��׾��RFy�$6�ŷ"@-� ��ol{_�~^�Y���,��[���q>�mK��N�8F/	�BA@�:�N��4�Z�G7"~!��ԐCnD�'&�g����\������fe�����T�?о ��-�$�{Y͎=���4�H+DJ�$$c$��đ�)�$�Ol>��=�t�Q�]]L�� �w9	��8�ԂnD�[a>�fE�ߕ�t�y�{��Q��%�6ǧ�5P �F� �m� �ԀA��������[�`�r#�4j �^��N���6k�)��]f��#*P��;��ǚ�G���W2l�+�������C�57Od]\\M[����[(/�=��x���O~�&�5���W����xF/H%���~� �m�a�`�v�ы��5���ԀA6��/�hW��"��?R�u����yty�j}s+�|_B#7���m���p�m�5���ZS��7h/�o)��ۑ#��O�ّ}��z�/P<�_o5�V����H�[k��@��[knϡ��z(��m�+x�N79+�1{����/��R-����+�&�;*A
%�`���Ք*kX�<t�fK()����p�s�Q&.l�����{ھ��D���|@mȟ��O���>mڟ\��p2��g��C��*�~�ya����bA��В�������k�{�=m���2-��n�^��s�@oMվ�Rg}�k�؀Ώ�um} ኝ�E��qd9��br��
�${"��:W�|0�ݳ��������*8&R�ote����u���2����:�7gPw[�� W���9��%p�^�Am� �������n@n����GV���j��� �h/�hN^i�z;�/2��U�^�>UF�=#���P��q�� �Ё�$���͵M���'�u"@�����fE�ߕ�t�x ~/1O��r$��_6�8l<ցg��K5�0F@K�L���6&�դė�6Ӗ��u:ْά�ڵ���Fgݖ�@>p�{�Im��*��eo�����s��#��S5�]6Y"]_Y،��,w�����bw�Xǽ��G�73�T�Qq�0'������'�������6�W�J�_B �3z~m�K��=�o�~���$mm}-���������>ڐ��#u���;�/[��k� N�)ޑ?��|[r'��RF���,���F���-����nff�������s��#W��� ��y�N'����Y�)xH$�Fd�By�Q!�~�L���n��D�8�﫛�vC�3,+N�d����5��	3���+�nM��vq ��=���(��W�?zD�Ch Am�rwu��|���ؿg���'��q�r�̯C�j�jW����8�D��R%���ɟS3�A"'�B�5���v���ݺ�ʽb�b��B��EW(�(
fLJ�����!$����Ԑ�C�Z����R���r����B��7�s�����$�/�hH-�$�"5�N�HR>�.�9O�[\?8C/3Y[��W�q�ɟ���	�F�m�^~��i\��zr@ۿ� �)܉!��!�#}{龞��{{v�'<^�U�R�?�D}"Km} ��B����fD��J�T���G;��nD��q��1Oi��r�yw1I��]Gb�/E*���t���n>�r$�ׯw��
 �}���o���+��&|#W����A�S�܌r�n�Ld�d`�79t�N�e�"��+vpf����OiR��ͩ	�w!��+9��ܲz宛֘y�:ؼ�7�����&���N��yB���i���C��
���GJ��G6�C�s�[nr�e���@omf㵖�<W�( Q��$��U����	q�N�^.f�췴3�,���8�=�w��:-Ԥi)uV4;P�4���8�s��\j�G��e�_��Y�v48vk�c�r�RH=K��}��<b��-�2��y�M6n]L"�:Wm1�Acݨ9���y!��vX����X
��H$WKwu&��>��y�Α�Ġ/0�]�^<��ܫ�����}����P���$ ;�����q4�]�x��Z)&Ç�!\�f��.���vx:Gc�y�di��X[�YܜF=իb����+�L�`M���[rh�ݲk��@۾�n��u!�@L��v$�pa���i�J\\J�bc>d:�F?�A:ؖ�ups��6��Ŕ��6�,�[y��^��e�\�/6��v8)yvlJF7�ZU��P"p��b����jYZ/��Ȳ���}��^�۬r�iD�')�o�o*ήy$5�nʛ�i;��o�F�䳨�ç�݉X�2;D����{6��vNs��e�m>U-����W3�a�'%nBmL�a#�7��9��w�s5�
5(SfM�E_U���5��.��Ֆ�h�>�D��8�a[�Y����32�8x�X"�@Z�kR��V�x3/omoD�"=�gR�و`pf�^��f׬��Uͽ�}��u_)�v��!�d�{���/{���*Wޜ�B�z�l�h^�tׅyx�Hpz�,��܍.�� /"0�}y���̓'u��z�i�V�V�����_}s��jit�S�5����Z)e��g��;��ƙ��������z��:h9�Dwmm��q�m��e�{گ���s�uֺ�O��eՏ]�e�����e�v��j�����+C��x��3�騇�ͬ`v���U�kڟ{�jX�{{�����ƾ���Z�{���`fc9��W��|�s����>����Z���Vu�䵾���9:g���I���m{���췗o
����KN����ɇ�����)kUuY.b�m{�{M:�\[z��R���;{�Uں�œkNZ�%kz�>�F6!j�7�K�P��	�%����7n�8���8~tөNx�0!�g���Cn78�۝��b�@#���4Ў�;s�'E7hyٞz)�Fbb7G@�aab�h�, �kc����M�[���p��B���j�Lݴݹ�n�&Ŝ�԰�X�,��k���Ŋ$%����d�su��v��K����)�9EM�cERcOf�=9�"��b6S8��'�sc�vwZ�L��!��|ѽ.��0��gb�M�+9�>:1�S���\�i4=Vڵ�d:�;VȜ�S���n�{���7F.Є7o�;��lh�v�6�-�U94���$m���Z�N��j��MɌ�&.���f����9��#����h��F��
ą���Ѣ��Gc[];��Z�ŻI��J�=:���]p/�Mk��],� зn�.�j���ϏH(��~�GX6�d��	���ED���еKZ�!^	{B�t�K4�̡��2ݳ��D�Ul
YJ��	FiJ�s�&Xi��ᗏ/j���2�ՙ���a��u�5�s�0iy�q�Ę�ٌ�	��aJF�lv�9��(����gYQ(�N
^�/�� ���cc���S�X�#4f���,f�Å���ؓ[ �\�-�ͥM1�S94F�u���&0W�2rm�;'to��������x�%�n��6�ؔ�]I�[����6�!���W���pq[tI�#���fH�����kF8�،4v"-Y�c6ft�V�I.9n:�c�\X��mN�p�bBV.�ۣR�s�"�/^b�ҒX�n8�Bmc4Z�-�u��(�Yq�M�"�ʛ��89w
Q��e��ƈb���(��Ύ���\����K�$ҕ����e�s�It�n0>��)�ɜ�b�b�J����n5�qX��s�,��Ș0l]5��6�DQ7:�$&7�Gjih���pOc�2<��Y�p�m���d
�����I���lL���� ��F��V�MF85#c���g���A=F*������\��+׏< (����-�D>�C�:�\<Wv�<��ފ�i����f�]��Z�vB7Bf�vx�J[�����fz����[�n=�b혫�]�`m`O,g��8�튽\M�t�[�7�(����v����F�l79�� ��<�H��m��[ے�{zǝ�p;�5�ӈY��:'1��W���a[+�!Mv��$��>�;�X���c���^ɛ&�����8t��vе�ؘ�R::�O޿̽|����t��}m�w��w���'<^�U�R���ם���/���k$Oǟ��A���BKm�z�zpw��Ԑ@��D״�}�Y�{O�[��5���) ����G��ɗ��P���?A�B ��Im� �⺱����ڲ�cw��O]t^7Y3��?n�$��[jA6�O�7 ��q�Va��k|���$�y��/sW�{���g�7q^�+����;{���en>�}�����!�"A��А-��-��Ѥ�WR&�K��u�3�}��ρ� N�/�Z��?6�q�]�\��9ނ�B��Q(�e
RDƍc6�yc�w�Lb:k����Fb����w�?�ۄAߜ��_an^n�[�7��7Ng�5x	����E�qq���퀁��A�"A�� ���C|�?U�{n�P�*V���bde����� լ�Y;u&�K����蝘�%]1�bU�v�G��M1��"�y��$�oM' ���#|�_�}"�5p�;ux��7q]jW� �B��������]��nh�sc�[r<�~m|�V!�#�����H�ۮ�[��3��u���'s�A�r$A|�B@-�?�����"ET�Ɉ���s�I��/�^n���(��F6���5xH'u� �DϢ��1�|k�I�ȐCimHۑ?��z��䢷��Bþ���uu^��Cw�R��~�A��$���A����,�i���f��蓗�2�p���;/A�[f*�vL���].ؿg���	�j#����nD�����2g�ѭ��0:8_Ρl�fdon/����͵�ma�ۛ��<���~ ��?A}/7\l����F6����N�BH!��m�Sb.}���tȒ/��y|�Cn>m�3�4NuJ1<͉����La�sx�/&�5{�Im5�{�J�"��v�q>��6�Z�P��D�z����V��Y�WY�jq��.X���'s+j�c�n�JW��>CH��RA���bE}���������x���H-��\>��,��5�s�ς��)!z�C^�&�_��bAԾ#��'��S�� ۑ%��=���>kRLp3�]��ѳܥ_�1뻟k�	�hH ��m��܏U���ίM�Ah��)h`e�2�6��b3#u

A�gF�8�����IDD��M�A�5����Ci|[r/<˞�w���Eu)_w��x�!��o�$����?�R��!�"~m�$)�pzbz)�A���ޑ#�a��ub��8׮��� N�) ��ȟ���P�O�܉7澟��B�r$ڒ	����q���M��}2��{��#���u�ܾm���rv���n^Or���w%�����Yۅ���_x������=ތMU���usJ�0Lu�j�nWE.SPB�p@f�	O��J޳�*���CEÈ�[��H��;�w����w�E�����6��$��_���O��8D6�A����@ڟT���P��1���{�Oyƽw>
<㹊~#B~!�����c�;�}���}cqߥ~<Dq��x�CՔ���(y��<s M�)���f
`��+�����%����n2�u�Ϝʱ绮��G/}"s���}��e�R��A sܤ~mȒA�m���|0�5��Er�}�Б[���t�do�u�^�z ���H-��=㧅���.���܄�͠�-� �ېVUh'�2�I�S�ڵ���^����)�~��O�6������_{3�!!�ڣ7f$���O�ܰ��!�����s���No�9xH ��̃�秇�2s>�^���;ޑ ���Ԑ[r$���ú�w��{{C���R'��Ͻ�Ց��-�W�ex������ޑ%����/�Wo�
��\Ȣ�oGZ��+ӑHg��$ei�%cj��d�.f��"J�����ck�/
J5�f�P5���o��M`L�/�1>_s��
�Ѯꐱi��q4�[�mhB]  �Z��N�W�B�ˬ�rj[�;�MpL�1�Z�H��nzێ�@��[�����#;��ݺ�R���t!(Kw[6F�MwcBg�c+Mj�ѭϟGLj�<���y|\k��u(N���e�&��r�:,�N��� �|�^�.��s\pg]�s�oKU�C�8̚N��}pf5��Fً�ʰ�`�����+A��P�{0�t��hM6�g���x�sZ��b�M���&%G�u��ߚ!��m�!���i���,�������P�q�u�Qt���ٹ"H�K�ۑ%���-�#����w� �ە�0ep����d���s�s���No�%� �u��? �m�q��H�3�@��	�� �ۑ?5�ŷ"�Fٴ��i�{��#]�n��S+�����^���XA-�ʹ+nФ��!�׈_�U�@ܾ�ۑ=�9>�]�����s���)U���2����:������k%�D6В�J}U���
��nW���?����?u+��n�s~���x��G��m����nDU��{�~eW~{��kPq�V��\��d͎:��P��Ֆ�.�PΆ�F���}����}t�ϯ�$��|�BGc������^��+�2�Gw������ ��ȓ�j~?76����@R��z���2�T���5b�� j�mwl�1<�y�����g(�i��M�1�4�*�
�A���uM��}�W�9���~9��aM�+�$�^9澐3���i���/y���������s��6X�{�-���;{��\��׵H �[��'��R��D�&njT�ry	���W;����rHx�����-�$܉!���\�M(�?xk��/��C~#z>@6�H��o�ޞ����n��S+��z#�ͼ	-���+�_5�w�r'��!�-���w59�S�}�*�s�y���gu�s�Ǘט���9n>A�"�_���Pz-���s���d4�5�䭻Djm�ҍ�>u�}���n��Lܬ�pYM�ɒ�����,���3���5�ڐA�YON��֮v?njs~��9�+-����$��� ��k���_kjH�WL�'ɎB�p�)�����u�/r���^��+�2��"��D�[iVJ��U��9L��K�@>�B~!���_O͹>���Ī�'=���2wt���O*�l��Rw,��O:�r����Aۚ��(��s�4sw���g^(,�V_h��=���ݫ�-�����f/�� ����ۑ �ԀF��N'}����Tix���� ��,�ӭou���njs~�x��z7���S�i�� ��zD�_ ~-� �ۑ$6�6'��o�z/�\vH�ލ�O�t�z���W�exOzc�mI�r��+%�P��3%�׭a5u;S�u�l��gm�@�1iru���n�S&Dʃ�R�H?g���͵`�ۑ#���{��ާ��\߫��k!%��C~!��ۑ �Ԑ@-���>�&���DK��A��9�t��������;���?w�@��n��t�+�Rg�x{6D�ڐ ��$�r$���ۑ;��%Dj���Cb/2o��s��-*�L�G����ڐA-�!�"C��Q��r#Ҏ���� ��yH ��O�����>�8�o���b�GVFd��A���7��W9%vvG4�6܉�[��oXf��ذ�쳃{Ee1�8�#L�wcx����*\�jν�;��`�qz�
�m��|<Gt|���-�q[r$�u}�txN�;q�����٬�����q�A~A����5�r ������Aу�BAN���KfEY�c�$P[��ae�f&�����`̰����A�r'���nD�=��>��s����z�W��Q�fn�l�|��?>����݉����*o"׼�+���x�7�#<��g��f��<
�@�s-H �� ��nrx�W}���z��-� ��H-� �[��=�Ǧ:��*��(���vk*+�a��^�A���$���-� CnD��@�nws�i�~��־-�9�>��.����iW�ex�z>v����1`��}m�%���k�گL���>��ں���R5��=���Q{����x�Z�=�g�7&܍ޞ�V#�S�Dl�фNF��U�=�\Bi��J��r��V�ȼ��N+��.�Ɯ��S5Os�:�MVD��0n6�z��DNQ"`�24�e�(f��h��SE;S���py��q{�V��9y�T�l���&���pmź6��:�`l.������B�J�΁��x�x	hP�j�xNEn]��Ks�X�\�ns�q������k���F��OŹ��ݮ5�ɴ��%��-��8���7;=x#���t�W@��i�U��C`~���hO���F����،t-˙��B��5ɺ�Wg��DD�d����_� ����$ڒ	n6�5��+*��a��<� �ʨhK��HW�/� {�I�'�AmO�w�{��"��K�_/��nG���4��Sl4��ex�Ј#���̬�^j�����l}yw �^�'���-� ������\���g��>b^��u�g��k��z@n�ʹ$|[jH�|�^�)kϯ����'�w�I��Cv�uǺ�^�/nŹ�=(x��H#n����={�8K{��Gs�?�@��RAmȒڔ����e�q��-Ȑ�#���]'�M�ҿT���ބ c�-� �[�Iߛq��o�.R�
 �� �\K��n�J��ۨu���X�'Kl!�i��ɚ�J�e�o�	 ���-�$ۑ9��OvxN��^|�8Z7���>��kԚ�A����h/�mȐ[k�-�׊vH~>�]d\{-��j�N:ȉF��{��-�;������V�fbYa�yݛݽ����3�� �֍�n��*���6n�* J�h�T�-LQ^��ɟ�Ѻouǩ�{R�������7��/�mLv��.�ETȐE����jA6�I���
f���/��j^�&���Å}S+�|{ЁgzD��RA-�6��W@�i~γH�j޸H� ���-��o�x{���ou�:�3��2�г�	�S^"Ǭ)�=��|��OŶ��[���܉ �׳���
��0�º=�㫸^ԯnŹ�=>��q	?G͵d܏7~���F��&|�<u�gz���;.`�� e4�A�t��o<Y�n��Д	
N�V������!�6�_6О{�}ˤ�w[��W�BH���h�sQ���BN���Kp�m���BH�2v�ڽ�(�������'<�L��a����<u�k���~ ���H!��W�X�q>,b��>�'<ԟ����"~-� A|M-1�z�����vh�e�F�TH�{�S͡:���i\��[����Ź���.�*+�x����W,�U�������P!�vk)bu�^*�MB��o���}d��1,]e�G�p#w�/3��×����7P8	z��q��l;\�#3.։�H�20+�����2*�YJ*UN����7���n �z�w-��x8�o`�|���̌`�	L��[�p�f@�4���b��廾Ӛ�T��g=r5���4�e>Vss��ИVź�6��VT��^�9|;�{�@�'[~��lʼ�Y��A)=�����Ħ���c�iv�q R�'q�}WX�<ʣ��ڮE�Y����*{zbћ����v��^�+S��YYaC�2�*��t����ec� �� �n<�WJ������6��r�[ޛ�t`K��Z�XL��]��9ڰ�:�b����މ��*�-9�ˍ�aUgڛ�+V�\!��B7�D�]�tA���w�������i�!��"���D|tE8�.AU?Y�B���7K0k�û�kF�K���,�'��Ӳ�s�%.�j�՜ë��R�;Ekq��&�O��¬���p���ٝ8�]V�p"jwp7tsA���4hfّit2�[�$y�˼�RSۺSo�;�Ֆ��tET����Y��5'/tT	B&9�VZ��k���;Ey��z���z1��K�d�Zn�4:iH����>�SUfHt����W�,�e@4��ͼ�Y��No�ۛQ�M���N=�>��A$Ԍ�y����Fl$Mb[�q�R�Z���V������䵝:�d�Le�%u�G+�U3j��['��Zج���udy�ͼ�릳�K��Ln��U��J�fXl��7i�Zʛ2�{��v���oX��]��Z�Ѥ�:�f��.��^gz�5N��Þ����I3��kaT�ZE�@Դ�מzo^ٽE��9ѫ��J�Z�s]a)�:�ӣ*rk�r���y��5�1Mi��K6L�fR���N9ŀ�Z/.f�׽�kgD[��]6���Ӛޡ��Mk%Mu�Du��p��v��V�he�GZ�M(��.���N�cZ��z��E�y�t��ĕ*вX�R�,�ƪ�,�nUU*4Ϊ�ڴV,�ͧ5Ռ��vms��h�1�2�uk={<�5Z���M�e��N-%��mba�q�k;8z��\��of�Rթ�6���bH�3��Æ�N�mk2�&�%�yޮ�~�{Z��K��mx�9���C�����BA�P7��[��쎞���6D� �?6�O��t����m���̯|A�>U��c�>�cM>RA �B6������[A���3��GF�+�"@���χ��&�q�^��H?g�"Hm�m��a�m�����S��K��W*_�����f�+��핱Q��T�6n��߯���Y}}e��zD�ڟ�?�n��q��/jNm�^{�H�����2|� ���>�)ې�ڐ�1��m^v�Dm��=�F�K�jb{+[f*�fP����"Az���\��^b~*�/���܄���m�܅&�ʞ�K������M���^��̵$��Ci|�BKmI.m��Mz�{�\�p"�� �����q�3u�Svv�՚���}u�x>��KyB��e��l2��$�.^n�LR�����vļ��i��ʷ�>�C6� '������ҹz'�
�psLp�?W��s��ȟ���-� ��n|~�]���u�oG�ޮ\���b�ҥx�_���[j~ ��w�;clH�ޱ�
,i�N��-��.��@����f�`npX�fdDL�b}Hx�jG��RCm�ޞ����&�q���H�:9��^� w_��r$���[�G�3\����]mDT���� ��7Fn��w^¯Q�Ƽ
�} �w�����ͭj��G�*D�3`#��~ ��H7/�r5���=�:'�YK��\��ي�J����|��?6��p��:��9������ {Z�nD��{��|���ow�����!o�ƌ�Gɉ"�>@v�mH �[� 6�H-�Wd�֍�&��S���5����xH&�Py�-�$܈[#|���{rC&6��� �w"�*!�0�ƛfÐȇn0Y�}�U�݁�+�旊*[�����u�o2X͙�	Z�i�-N�q�ߴ~O>M3�<�$6��Q1K(�]L:G�4��0�)��r�Ԝ��-[=�΁�4�V�uslv�#��m�aR�I�%�h^Ҋ؈�l8�p��՗M{��,J�h��l/e�Vy�A�۷/��en%jh�2�,�uԅ1��E�&��H�������&%6!�B-�gKK�k�(Bi:gp�ms��܂ � �[�3+��Zl�(��m���sk��e�J3�f�K1���U���Qr���J�LA����34[u,��L֤���$����܏i����aWm��]��^#�����HƕA�r$�@7m��~m� �^�WǞc>9�R#|�Hݽ=G}��	��ok£� ~9x���H��l<�z���w|��"@>�) ���$ڒ-���׽��Ș�t���:9Zׁ�C��P���@_�RAm��Ŗ�[��TA�J&W^��_O>�$o �!�"{Nww�.^׍���̯|A���.�lyLtS��s1I��6����@Kh [i�D���z b�͹�9��w7[����_fb�;�`!�>_r'�����w���W+g$vx��C��/,���;k۠���N�V�2L��Z�~�B ���-�$�f���:�z�V���zB�b���qS���֤Cn@n������z~�Y.���t�(a�����9A:;�NY��=~<7;��΂�Ρ5�]�iv<J�/qɝ���B�_�Um+>�V�K�
�"�{܅�i����k��f��3+���,�Oʹ��W�9/I��'�y���6���@�Ԃ͹�a@���}�鲺�d�܇�ww[��J��� Fw��/�hOŶ���w��huH&�8�d���%���p�i������^���x�H&�P�=���>�oپL��v�m�!����fC��#~uL�xq�󮘊�xٺ�L���B�H��mI��2,t<A��9x5�գv%���jCvl)r��m��;�sȍ�I	T��R�GW/�9ܾm���"s�zxV�#���6[��|����D�ɿ�*�#�Ȑ}6в�RA�_
�Xw$t�x�T��
��������YZׁ�_UZ#��Q;Q><ԡ�>߰�'ܩ���D�{�	�Ծ������(~h��WW-~C�ni��yqϠQ��kb��9�xp?�B�R��������V����jfmGkX*R�ɵ��l�9��Lx����ͽ�N�sl�_�e{����?H�mI��_��:n1�%�-�yh#��-�>}<'}��۷�[��/�b�EZ�1�����xY�/���m����'��[�n�D-�GW}��=���8Ǭ�V���{���{�"�RAm�w"oײ}�?��������Kb���]�,и(8U�t.��D�j����Ά�[4u����[�����Ci|�B~�9���鈯7����̯*o�����Y7��k_`-�ͻ�Am� ��gF��bo�,P4�I�H����9�9����/| �� ��! �N�)s]���]��L���K�@�r'��@7�y�kv���k#G��^��z� ��B~#ހ�mI�"A����V��C�gʈ!�Ȓ<�_ۑ�;��t�"��l�_L�� �{Ё�t�����c0�ں�fCr�ˇsr�>�(��a���{YEz�+E��7�s�c*Tc��tv�w�kw7,�љt_������"hIm�$�ʹ�z#�'�W�g�Ǩ;ozxN�#��o'[�
^�|��w���mȞ����������Y�ĸ�<nRSv���m�|,��t��&��+Kt�d��Fo��=���6Y��9[k���t�h}]Y�~�Yzׁ�𐯲����rz�ހ�{�A�"A�E����}���B�:�/���D�i��~��m���)����_6�vpޑ8�B"��A=܄�h mI܎{Yz��Q��lO<�7�y:�xR�@���3����_�s�m`#�h�̭����=�"A���Kp����������e��W��A��$����1����X����r$����RA�6�H!��[�=�Y+���ٲ%�G��݂b�O[�7�2�~��o�OŶ��	n%{���
ڂ*��}s��2�&M8�c��]��B��	��ڸ7Ճo-l�ځCDwB�qtt�s�,ٗ��w:�S35�q��L�����3����l�66p�T5�a���4���S]ۗ!�.���[����b�6�lpA-���(�������(np��p=�u����W8�wnŪ뱗�+WR�m�<g]��%v7m�]u&n�[DB\�	h�m�v�+rh��*X\���\�v�i�"q1r8(ݺ����ں��[x�]���d �d���9��Q��h������������x��	���	�mM�,[�K[��IM�l�ZڙRg�����P��<�@�Ԑ�Bs}�<'}��sהۿ
P.���f=+�;��G��H#܂�����_H-���wyx���&43���|�������O��<k����^ $w�@��	�J���4{�_��RA��"A����"�H�ym{���-��������Jo�ex�ބA������A�D6�Fxn8�=���w�h ��{Z�hH��t��Gi�^Sn�)y�_@ۯ���ʎ,"㇈v��|�H-�$� A�6����a�ߢǺ�k��t,�e�U_Q�Ǎx�	���y[jH#�܃��4+eBI�e)���MGmDir�
4΂˒��[����X�ű٥��@���ӻ����?6�H�����&+��v���W�#آ�d�ݏC ��H�{��~-�ͻ�A-�$à_�+�vn�0�4�bU�G7�7�c��W#mrR���T��͈� Ev)oŜ�;Fø�����l_]�-#F�w��V�uQ7PD��r�F?!#7�����;r'�M����=��������3~���,��p}��!F��q`�ۑ?ڒ	n&����M���5����m8�.|�Y�Hy�-���ۑ ��B��#�n#Nw۫>ݑ?���܉�k���LW�u���)���zw^ɏy��/�ODxI�� �_�۟��BH!��mh�Q��N��t?o�N[�z�����e6��+���R gz@n���܋����_��{�O'�>X�|��sH&�"��$�zxYkV������.��v��5����~����g�=�}"~-� ��nf����c<V���#�<o ,nⓀ�$$�� �In�#Oۺ��{w�[�"1������:�����1]Y��+�R� ����$��U�jħ�����}�ېO��O��@�ԀAm��;�>�Qv/8I�Ge>�+i�ٽI�ܰ���&p��gPb���38�9��Y}j�[���si���v	��}2<�u�����}F�?�RAޑ ��������FNߑ\!�{ݓA�"A��'��}y��_59�|//]ǁ��������sՉ�@�ڤ|�D�H�Rm� ��4t���
/�M!�Vn�{_�J�Tf�b��W��s�D�[jA�	?z3������O����6+V�KM&�Ӗ�K���,��C�v� 髆�Wm�����Ͻ�����4 ��E���A�1�>����z�=�\�+��T�̷���ϼ�ܗ�6�H-�?~-�"�����5;� �I�\^f���&��7��ぇ�$^�$��A|[k=���z*�:1����D��G��+��ۑ ����ۑ�znrt�x��wۂUuF��xA�B�r'��R%���H��.�d�ۼ� �A�RA����Lm�+�g��ς�/��H#ʱ��ř�z�^�E)�ct�]��1V7[�'g`�e�'m=m�f�v�zr�S"U`�L����:B��R��Xϫ�X:�tҍ�d+�Օ��v%��"Km}?�[s�m{��,�Ju��_�Mp�7������M{�� �-�?~��#�O�Ӊ�>|��2���2jT�f��F�kAnRs��ŝt�q[��@���2X�@z���t����_6���]پ�+��n�����ZQ��zE�Bw?6�Ÿ@���ʹ$���X~�'�P)�]�I}�9���S�o�z�z޹�Y��^)�H��+c{�q���܉ ��R ���nD���An<,>�}U��ɚ�\^^����{�G���hH!��<7�aoe6ǥx�\F�! �K�ۑ�ܻ�}�Wm�a_+���z�Cb��3�Lq�yH ��6������h"�]�����g�D����U���g��><'���o�I�ʹ0|>�Ff{��KZ�7�kw
]j��ԦH^���w|q5M���Y��A��O��GN�`[÷�^Vse�crͼ ��
%��ON��Ro��7cb�Ӫ�ݤ�m��[I�|B��Wo��J���թ�"�V��Z�ܻB&�2^%�D��_W1��/E��(�k�1����n���'�g�ڼ<X�f�����9[6�[:R�86bF!�Z�v�t���#�t����'w>Uw�n*q��(7��$��$>T).���/w/j�=>2�.\C���J�k�|�i�7��M�+
��QBI�w$3,���q���9�Un3uUP�s;,��$���lQ۸�PLF��~����k���Yc,���#�]2���0�qr���3��`�]}��$*e���ne���x	���c=�����=�����l]ɼ�c]:ˡb�hP���O0uq(7�Pc뤦�f�m�6�k{��ܽ��~(�=z�m"/�C{-�M���u;�*}�oS ����YWs�Z�wU�R���AN�i:$�+T���/�r��tC�'5��T����Ͷ��ok��-��iޠE�Zѽؗs��Y�6�Xu��F�{�Y��p>ΣK�흶boQ�k|P �t=9��j�)O
���U�����c��6b^Z6"i�����]�=�׸.��70,�+Z	fMg9�!��N���P��p߻G7��n� m��6�)��b7rj�cT1E*Ź�.iT����kwk*�,ưC�a���tFԇ�,Ň�%�Woi X�F�m ���U�\���O{�i��#�M+�Uڭ4��V��œ-��&���շ,S9��i�4�i��u�WCOzޑ62�ޯV�Ċ3:��޺w����p�W%k���)srk4�ZceN'�y��y�o5-5&��6trjՔќή�ue6�9��e�K)γ2o[��լ3S{�{3�m*��ֱ�i:�3��k9��,�Gyq��m5jɩU��i�Ir���,�Z�k���a��k64�4��4��A��z��k����*�Fd��-2i�O{^j䲡i�lev7Xr�%�j��g�lw��ֵ�k����O&m���y�R�
��f3��Ǫ�-t�9�j�7�{I3%EW������O=�{1SWL�{{{v;M��؛���U��n4�15�i��d���F*´64�g�=��,�{�Y��m)��ٮl�N��櫂N3uXl�0�ٞ���f�]�{�3����ꖫ�4�[�{]���,aJ�����3�<���0;R�2�)ڔ"Tl�R����f�V,U���ԇi��=��l�����d�k�%3��l0k���}�`K�b5����3��sy�,HF�@�m*�yj.�	���n�q� �I^Z���7Ip���h6�v��N��>f�]����U/0�s��BjE ��4Y�=r�)���]�{wk���b�6f�ٵ��S]��Z� k,��b<����N㋷.r�xP՚uNH����ѡ�Ymp��[$n�7gsm I*�\l�//>2K�ܬ�@��C���v��d3ْq���u����	|�?��=�35Z����{�6 p�GK�5�)�=Sv:��P�ݭ�v��$cm��:c��qyB�1�m��p1R�"Jl��lt\�\tV�st���s���`'���VM��9���y�ʱ�-�j�%+�Τ�#F�X��\ʎ�k�()m���Y� i������j�B��6^l+jV�f�#7Q	�m#��1x�ً�u��K�m�+�l��Q��y{x�=\�Kf8����-mp�(<&8t�4��l�k��.��5!@���R�;.�.qe2e��eɝ�b��[*]H�h�oFI}�%��X鰼�.U�\���0%�p�Θ`+cn�zI�ݫqV�ۺp��<O=,^"�IiS����[i]W[\;q7
>�<"��1`��x&ݬ�Bq��:��l�	tqo<�]VNp�>���(��Lx����]��t���=�*cLl)M��˯.Fk
gl�PFK�-Wmqf��s�^Eث!��pځ��H�0��c35hŖ7gluh.ֈ;
�żOkvS�r$���3���&�]$Bkl!���d�Me�c5���wSf9��L����)w.���j���'��M� F(��,�5�U+c�D�<n�\ˮ{nt��Ju��^��nG�Onɫ�`��[
R�CZ�����s��P����89�Ap��<��\�<�]��L��tڪ�Bؼ�/�1��=�vڂ�,��Ƀ��&Η\��ں��me*d�mt����1�8�$�GCι9�kGD�et�]Yy�Mtkh��9_sujܷNz�K����w�]�U�"u+��bnM�H�W��.U���F�� �s^%.���e�F�mC�� �c�%�t�mq�:�w7rK<e�w7H�!�ٺ��2`�Zq&�n���YW]�������;N���n����w�"���y�Y[�)r���Z�\
�������@�;O͵���!y�7_9������q�a�F�e��١�܃4=�R-��Ŷ�����щP��4����D��.�~�+�+7XW咾��!�r$��M�f�,>�2"��~�y	 �����B[՘��}�w��n���V��mς��կ��o�O�6�_�r$�ԑk��1L���J7���"NsR~n����p�5�������	�b���9'ՃNw)ޑ$6� �Ԑ[r$��c�ߘŒ=�˽�~2�En�|�W�?�"yȐ[jH?�y�����s�f�P�y;�/=s		����J:�{j7�x���+3i9��d*L��A��'���ڰA��"F{�uUm�-��mς�*��v�D���J�/�	o/�͵�m �}����n�O.�>SFa�3',o^����O�o�������C%�Vc��vN�f�9)0e♨�hf����zD+��7��R���/ؤ�{��1����3�z�<?	�^�$��mE����Օ�k���椂ۑ$6�_6Ј��*����Ef��+W���)��`ߖJ�� A7��mg��[��h-���[�ö�:�'�	�u�$܉����~[���>
�x�b�8AZz.7"t�{�A|F����ρ��"hIm�Ʀѡ �Z���rs|<�]��-zA5�BApŶ�CnFa��� �Y�T��DPB"���T�'�n�٣k\��^6`޸ݱX�\ [vk�ߗ� ��Ԑ@��k_/�nD����u�+�+3X7咼���=��Ϊ�2x�X ��ȟ��r��?�s ��BH��/"'V�_W�����S��r$k���~[k��>0=��� �3}"Hn��<f�[�5R$��'���BKmH ��D�m/W{WG���ɺ�W�%�+q.ޝ�s����6���@(*��J����՝`	�F�S륻S��sEjr�=I+ɳKmΫa��m��Z��^�$�/�k��u���eɛu���;=׈!ۑ${����H����׌�h��`ߒ��AބG\΋�#=	I���A�j@ �о!��В͠�-�S��q��v`��~�{�ު����X��s�����?Fo�I�ʹ3gu�O>z��=�,��>��1�`@�l�41�fSi���K]R:::9�\�m�j�����e�~�~~r$�Ԃ-��u?t�v3�m��0����&��B�����ې�͵$\���S���U�`����r$ws��u������^ �{Ё�_6���:�}֑���j�	�{�_6��Cm�Ld�w��(�~��ݹ���۞>يH9��$6�ŷ"@-�����uTި=�"z���r�A�W������3�m��-xO��BA���4�0��O����vS��z�2��/%���^���}GQ�Հ<j�Zj+
��3V�7Dl�I���Ov!�:�em�؋�v��
=���H��m|�-� �ۑ ���6c�b���U���������5��咽���o�Im� ��@�W�A�&�\\OB�%����P�&�ȷl��z��8�=�7�2 ̩�3'���$zА}�_HmȞ��魷�[>���\�l�?e�� �J�7�D�G�|�!�"~-�'���y���Ž�#��w�� �B���K��|�.۳�a�A5�@N�m���(��3�s/�����}�Rm�$6���r2gX���U,��K}5�Nbw�^k��W����r$�RA���r/J����3}��Y���?CnG���k/}sKg��<.|'���{�cG
��+|f/��H�[jH%�Dۑ%��U�B�*�a�0�_d/t��C�vݟ�A��Io�E����nD����mw�J����g�����ؾ� �ĳڷ����J�~}�g?b��ӾY�-t&�q����zJ�r�&����]K�dК�ʉD!f`Z�$��V���!�WY�V�7�\Sc�"����zY�-�M�AkZQ�L:�1��&飠g�/`�`��h`&�K	���9W:,�٢�܈��)ӛ;h5�j;�b��x:���0�Lv��9��ܢm���:MH�K�����G���^y����{�E칓mX`:����
��E�,l��M(�4314q�����ϦP8��{NB��e<솪�rm9���w�wnj J�_L�������R!�H�_6БϟO7^�����`ߖJ�ʻ��Z�{{�p� ��"O?)[�m� ��ﳢP'}"sF����~���m>��u��������z�I7�$��c����~�l��缤�wЈ 6�OŶ��[������-J��Gao"��<?	׵	o�/�mH ��H!��u�����x�v�m�<��y�T�����d�G�#�(�Sᬉ�W�xg��;Ё��Km	!��[j���'t_�9"m���[n�U�n�.�޼RA�� ���ۑ�nd�C2� �~˅�tL�tn�q��W���-�p�+E�n댗J80���I@����oЁv���k�\!������Ȭnρ�� ߹m0��A� ����BHm KmI�g��ߤEQu3oVT�ܕ��lӌ䀷�r�~�P��#���ѹ��=��5j:u͢\�8�Qu��^Ǫ�(�r�d��Y��G���7�s�sپ�3�r�X7�%x��@��$څ���E��9���Bmzd�� ���_6Ќ��3�bfĶ����z�7�����@�}�����Ck�!�"@-�$B>���;��+v3��H�s��A �nf�~���|�+��Z�M{P��60��ӻ�~:�O����	m��r$�<����9�N��{*D���^��Rw��ɿ+����s}"Am� ���뗶���Wz��^AB+�n`����Rl�0�*���Ɛ�\�m��	'����̐A�H ��AڐAmȑ�z�Um���U�u�7�"�\b1�=z� �d�>��hYm� ��"1���76�lOd~^���P�C�o蜳ߢ��>y���-/��<�"�N߰���՞���H����� ��O�܉�������M����p�R��T�
��X�k�IT�H%@���:���X��w��^�Z��Y6�!T
f��'F��J�@16e�f�nt݋!�i�~�(q�3|�m�� Cm
�S�⁯gk��(�/���A�"G��|���x^��[�	� �>�R�3+���ܔ`�k&���3�|Gk�%���n>A�"~-���U�jȥQ�@;л�Q~���w�k1�Z��	�jA���m���#��s^��кw�AЇ���&` T�%�k��8��U�sƮq�Vͪqma�����9�澐7zD��|�mȟ�q�~�����My\��}��<�z�<1Y/U��q{�9�) �� mȐKm	��h�p�?o������zD��7ڮ�O�������يA7�H7=�{F_���!gs�H%��ۑ �ԐAn#�O?��}[�l���������W�^�$G�������"Hm!�#��8й�-��H���_�mȑ����t��_�f�k��}��A|{�y��]I13g�q�iu��h�}8O2�q9Aޮ���h��-��c�R�G�`��ߥF�]�WK�y����� w�!��AZBK?W� ��s?6АCp-�B}��*�x,�"}�wݪ���^��[�� O��ٽ"Hm����v���z���|��g�Q�bb��jm5�v�ͨ͜s a�3�:���5��5����O���}>��D�[jH%�[{�?>����k1�uzG5y
�K�'�u��{P_>_Hmȟ�m Am��:�rk(_�'�9�����9���7�J�ߕ�k��x�_���[i���}�}/i���|�A<��[k�m��S��3��������/]n7^~@�f)��3zD���|[r$�Ԑ|�d}��ӽ���{yI��[{�7݋���c����H&��I\r��5ӯ��\A����m���ۑ$7ۓq�Z��s�̏P�\��k�>��7�y���^ ��"?H�[jH%������y����?2-��G��<�+9$��·{UJ�gbl;�g8s`�hDQ�D���=
L���k;f����ʺķu	Y7��R�R���������e���°ť��Ve�յ��D]4¼�I6z����]�oj�k�RqjIv��;mf�6�D�L�3���h�"�/[���m�F͝�]�Sj��sYE�lX\�K���g]{8���a�Zb�R��Ļ\m�DKY���7!ܷ]v�9�c��ۋ]]S=q���FX���s�ݺ{Fr���\��\Z�11A�������v,{6`�� V��6&��Lۦ�͹&��iX��CiRdЪT�S'�:��hI��[j~܉�k�S�{��n�.�7F��t-��t�/�ڀ}{�܉��@-�)N��GnϷY�^� ����M�b�9�9o�:�$^�'�A� �mFɚz�r����m��"~!�;�O�܉6���܎����o�zfb����6��^W(����?6�	n!���=�[0r���/�Z����Amȟ�ޮ�s�{��n�.�?f)`հw��'�d;K���� �ԂŸD���IiǱ�8�B������9�9o�:�'��! ��A�Rm�GN,�ý�?�~�����$��Ѕ�)-JRU�֐��,��mT*��m��g����>{�����Nr�$�iwIZ�]i��:~��2>�o���DE�w"Oo��p�m̂m���|}}sP��&eNM����V7�ks�v0�g�s�7�v������I�K�.1\4S�=ut�$��HCJ�q蛚�$�`�y_�����D���OmU�����������$��'�UY[V��@U�$�H�"mȒ�R�*�:�}��RA]k�{���c�k�H&��H ������|Ch!����)�EE�e{'ɐs6D���������>��=��C�r�%� ���0W�vT�`�<����Cnd�m	����bEg{.�����o��dH����jm��dzs����ׁf�݀�m�ٛ��E�>�����%f	QW�7Z����hN�8qѦ�=��Z�,am��`�T������_^�G~k��� ��е�d��~Ö�ׄ�d_7�v�HP � ��jA�܉6�@��R�Q�������{5|s}#sw��ح�֯t�|�W��"�������!�����Gޭ����CpŶ��ۑ_}}Wц��g?�N�vf�&_j7x: |UvZ9���g+I�,h�����Yb�ft��Onh���j�͖�|y�
�n�V�C�����Յi׆5NN�ĩԴif��mT�S�,�i-�Y��p�א��N�dͭ	"�ެ�&�fMu:��h�5XkJ��R�3�ϱ]�&���Q�9���ȗn��J���y�iڻ��J�%@t뽜�x���9�?��Uz����췕���b�5Y��͈VX�>����Y��uo#�u*�F҇e�;^G{29����h���<%�6��1��w]��I:�N�.�|�Uv�f�����0��̗�2�
v�2�c=��0ɕח��	�b����+� ܻG(��`��*W:ݨ�w�a^�D+����f�9֫�#
+��F�VXv�B�l���*nV'�d��u/�O]t�ңpP����voϳp�f툪m;��vf�J���5u��Z���؎�c�`�[v0�ú��N}6f�6����2n�p�r�i�n��ݙÎb�������ӄk'5[�tS�9��S�ݞ�2֜++ ���f�X�wgf�}�\��>	�>�b����/t�B�f�m$�0b�¤eP�a�MÉV!Q-�b�uҗ]yq��N�Ȇ5Y��a��a�3��]��7�ify��5�(�9��V����ΐ�R%�I��w{����)�F[&�f��2���˙�nNL�,�0%uDR�Q���N�m+�ӯ�M��ͨ�a0-��r��x^Q���T�$�N�� 7�����4�Z�X�U5fZ2��ҷ\9����c�ڳNiԊ���;�̳�^{����T��f^y�ԁKx��o�X�ƍ_g�Vћz����j���+���<�{��;ks8�U�-Z�XmVt�hf�y��=y����6�eGU���un�	��SV�T�l�^�ל�6s��Z8`X��j��
�Wd�1,c���`pj��5��јt:�h��mc�3fgz�͝4ꕪ��c�[X�odq�s�;M�F6�Y�sM���s�hXl�1�,��<����a�Ms�׽�+�ֵ�QV
�T��YuF3*��8����ǖcT
�&���޵mV:��/]<�jta�:������ٜ��Gf�mZ�33g�kVN�f�`Ζeq��:�͙�޵�]�9f#8�f�c�vl�$`$��u[3x�w!������}����oH�m|�!�"KmO�[Ε�`�ْ$�r�A-�ot-~�����xǁk�O��BH+���zLh�n�����"Hm KmH �ۑ?��`�����P��"@�z���z<��K咼���Im���[���
����H(_�h��+�2�K�).f�$�pvpX��&���\AKW��egϸ`���Xa�l��{x!m���}Y3z�ۑ�1��w���o�T����^���Ȓ<�_�s�ma�{7��¨s�;X��_I}�е�d�g�#-�>�	ױ	 �E��'�����x]y	��� 缾m�k��Ϣ�>��}8��s�z=7{����^ �� �1�D�ڒ-�6�A�j��R<�E�/��#����MmO�#�cu��� A��$<w�;�~>�9�S݆�Mۺ��lݰ�VB�F,%hWq��F�Gv� �T��$\ϝ�T���](ۭ�q0�#w�K����-� An�#��K�}b��4Ds�S�ak�d�g�1[z|5����?? �mI6�t{���FK��������0�.�ʹu�-�4�41�,�ֶ�N{.#�Z�4GRo���z����Yg��!��?6�ny����z:��K��{�#xJ�r�^�IJb��W�^4$��O��|�B�m	#�<#}�Uy������) ��#�Ϻ�M:�nG�cu�w�����$��*Ʃ����p��$����}~mȐ[k�-åQ�L��T>9⳯1f�Fb���~�A�bC�[jHm� ���vt;��Av�w{�A�H�%�mȝ�o�6�^����y\���}�ع�¢�b���$�RA=��m-�'�mm{:s�������G������r�n�]� O^)#7��ʹ*{JB�Ͳ����;F�+�R[�N�Xe�؃��M�f�m���b�%�_!��1b|����X&���6�˝E�K�����ލ����c S6]b���f�b�a3qc��6����Tu�<%u��췮gXB�C��R�j� �ЦY��몆'Vu�:+f��2�6��n �Q��6f[�5���#��Tq5.�fm4�p���h�����Fǥ݋B�UN`�:�[���m��h��&���e�wS<���;>�8�y�,GOb�
�`oϞ��}�3�J�HE��ݚf;P=n�'L,������q�2f�sm51W��ޟ�/_�G��� ڐ �y����|������vzQ�~��IM-�3��}��?6�I����Ԑ���=Q�ԇ����%�>Cs�����к�t�\�W� �о ��ޑ%��t�Nn��ǂ>�@����w�	 ��@�ԂnC�5�ž��OH��t�k*{rN7^~׊H9�"Hm �!�"Am�:�;9��U��G���$|s�}%���P�<Ow�1[zx~�M{�GxW�5^�����!�H�Cpm� �ې�NF���o�5"E���M��z�F�^����/� A�=�m} ��%ZS��R}>�~����W��Map� �vu�G����c�$4���:��I(ʉT���O����BH~��m� �܉��ճ4�z�=��
�6m���hN�4��Um�#Z_6П�mO��"'��9I��Ӳ23�ZSB��91;���a���&�n�[�aT�1lH9^�^eL9��Uǵ/~';�u��˝+�&y.��Z�L�������}����,�����w�x��>���؀����گ{ϊ�����>��d܉!���܎�꙽ký���<���:��znW��� A�zD�ڒ-�!�2)��%��WJ��o��ۑ����Uj�^�b��_���H#v��φ[u�4�|$����/�k%�_[r$��r<Q�33bAW:q���:w}7����a�H?�! ��_6��ۑ9���<���@f���H���0�g2��m�`�L���F�6(�f-1dD�k������	ﯟ>) ��"~7&܉�s����нW�X�M��;Ӧ7�v}�G�$�H[��w�[hI�n��#{��q�#{�H��}[*��^Ǳcu�WuZ� �ސ��I�"!Vg���$�jH �?6����A ����I�BNv�5����Z-mX�C5��8�l�IK���d۱wV��Q�]לI�'n��߂�1^��2�2`����f1Wr�T��\�w76szo����C��!$�A|[jA�"Hm|�Z&�x����y` �f���|[r&����O�h^�ѬW��x���v�>�wf�dN����Јm���BA�m�{���*�|}3%�5#w}��Z�ױڱ��W�	��oH�K���n���8��|��V͂��k��m������8*�|�ӟ7h;S0�D	(⼿~6��;H�[j~?7e�o�:s]b�y�8_g��C�U�o�k������nD�A[k�7� �R���a���������ҽW�X�M�� ��#=�'��Wsy#Ngr��y=�LW��y2�u�$7ڟ�m�9Up�{{~��ܚR���j�߅_���jH��$A|�BAm�#<(:t4i�K��=n$�5�D���$�p�3R��ە���Z�<?	�!$6<48��51�^��ڹ���n�x=`�V3A�y��z�E���i��ZyU�B��l�J80TL�1C��@�hB�J�2P�}u��;zD���mI܉!����QHk�^����ț�Ͻ.�N���F�^�����������pf�;�5��@�~h���"B%@�����{;n�m+v6B�9��Ԃ�g�f�Mt��ߦ��� ��jy��-�$܏wj��Jc}{�)�~��n>������ˈ?vz@��|~mȟ�mO��"M��hDCw�]4� �35-��ܽ�^�k��0� �^�$�=�-���jsK4DbC��8ڐA�m �?6�Phy���E��N��[ӱ>�ѬW��x�_B �"@-�?Kp�!� Hk��邎b�F�|���ۑ#�ѽ�J�{O��=���Z����;��}�[{¾#ޏ��!ڟ���ɷ"Am�G}���X���n�ja	�ļ��r��{�#���M{�/�j�-��g�ٍc���ac�l��:�>�u�b �vpӺ̽n�B	��.���XsJ&���[J]Y0	ʋ�ʋ�!���R?T �|���=Q(no2q���n���q�<��vB��m�춺�<���*Z��ݶ�1l��1��H�l!,��"8�%���4)�؍���koh�k��nV��3Ʊ�t��C���莫���N8�hb��h��	ku��Y䭮x�I�;&w=n֡Fㅀ��.
�&�j�p��z��S�&WnSa�ƞ�m��= ݇���}w�����Qpd�;�j�I�r�Yͪ�������.�bm˖J3?���^�O���w���܉�^�_z]����^�b�7+���٦}�j�z2��Q?��H�皐A��݉��BHp���{aҭbO���ۑ=�ݴ�˯i�ԫ~~}�jH��~�\��E�1��Mȓ~�${�[s�m` ��f�72D��M��M����=ȭy?H ױ>�-�$ۑ �v�q�M���A�;�O���-�{���ﴝ���'��xA���y[�W��m����j�	ޅ��	m� ��"�Z����ğ9���,;"@�tw���˯i�ԫ~~_uڒ��Cq��պV-�� ��b �x�� ��\0�CdCl�3(暁�u���m���������8��"�mH �[�33uO���l�r+^G�������n�1/��A� sy}-��@��S�"ß����剃�-	1�#�'�.��D�������\SYȉu����+�Y�;���`Gt?8F��r.:�vw?�I��.�<E����$nv����'f}{���_x�B ���OŶ���F�-���:>ז$y�[A�R!�"�,���>��Fr���*��/��}9� 7a|�BAm��=�w0�t��L A��ȓ�jH �33WWwl�Ϸ"u�x~�ױ	#V���̜��ߵH �D��|�W�6�Ԫk��0W����7="Gf7�K�i;3�ѬO��x�Bo�H-�$[�S[�O{6�M�-��asz:�'��0搋�.tX�hv�8��nq���gT"d�O4=��$@� �����ovJ�;^��R�����7U"{%7�{�;u	#���ۑ?ڒ	n�gzNf�t�G�xq��������]]ܷ6}��#��xH ױ	 ��m��ޝn_�zk��{�
e�Ƿ��[r$�|�r��=�I���5�Uy�oq�������<�� {r�))��J�]����omk�f�C�&rt���3J�j�����DF��br�\��T�ѬO��x�}{��m}��r$O�j�����!`� �y�ۑ<ov�.���R��]y}v�RkWGs�j�-�#�/���"~-� �n�ۑ%��i�O�A���8~�6��}��#���	�bA�[jH-����'����6O1Ӛ6���)�^�.�%4�ͪ�1iYk�u4�4�7��_�:��{�H!�ŷ"F�k�M��uO�t�>W+���j���\�͹���}�yxŸD6�A��АGnh��ޡK�$�O�~�9�ݽ�H\���mJ��u��>�S� ��!�q,r5W��d�HodOǭ� �w�m�͵���n,/^>
�2���c���{���p1ސ~5�B@ ���-��m���Aʒ��w+ ��$w%����k��y����t�|�/|A/�|G�ݞ��Y�Z�+��o5Ʃk=Պ���+7Vr�q������h���ɽ<�o>���#w��akC~k	�2���*k���+�f|<}~@o���	m�$�E�����t�dg��MJ�~�m!n}��Q:�.|��jA��n>�܏W���W~��B	R)a(�T��
���������:���zܾnX�����xA�B�o�OŶ��[�U�[��YknF���c���m����[������=�RCm	6��Ԃ0{��:��@���o�n{_*��vo�KG���A=Ё=�[k�=��U��#۳���rAmmH �ۑ^����{��-�W�s�;-~
�'�jAn������r$ڒN{ީO�j�L2�� �?�*�>�yK�ql�\w��{�D��9ٿ_�p 眉!����R-��{-�G�'���n�}�rk���R�A=Ё���9˞�9_�	BI����� HBO����$�BB��������$��!!I?���HBF�!$��	BI��$!	'�!!I>!!I(��!$�@��$����!$�D$!	'�!!I?�	BI��HBO��!$�����(+$�k%�0��;k0
 ��d��B��        �                          @ �  -� � (�    P ��@ P        ��� T	(   �� �A%$ITU*��)AP�	H�!P��"� �DR�IE�B%P	J�@P��J���P���   	�HR�R�%UR�P �D�6�
-� e���\�F�=�VuP�����&�F��R.�P�I2eA@( >   !��t(9 �$��@���` =;� =���cԔ�  a�
n��=�D�  � ��  }��Q%R�J��T�IIJ� xn������K��{�]
êA�������O`�R�vr����IY�=��mP  *�� n�}�=�GJw���{��u�#��z{ z�F�Gw�T���h��2 į;@�J�@  w�*!%*RJ��ETU�/ ��P-�r c��o@qJ����獀;��"vJ��@�{�$��lu����  �@;�*�I�U�.�AC�H��w :N{t����UUI��J�t��)S6�"���
������{5 
�C�  �ҁU%IJ�JR*�(��������*�2B���\�C�=z����� ���w��)<��.�w7DI,��@ P/�   X���^Z�}���(�t(ww)��X�"U��!BfԨR��E�P;�D�Uɒ�*�T���g��( TS�  �D��E
E)RU#�J�\�H��)�p���z
����։@���)R�=� �:�@����
��E��HQ@�>   �-IT��J�C�%��R��R�',��U���BfҊ��Q�@��(P9 h9� tn�H��T�2�ҥT�@h2d0�?i)J��  �Ѫ�)$ ��4�*@�� �	Oԥ*zOU10 `�L�=MT��5 )?����������BIq$Q�|p���߹�ǿ��� �$�����%`! ����I_�	!K�$ I1@>�}���]�����ݺ�Un�������d
Xչ�Pn�Z��-��M�n��t�KTc"���X`��IFV7���pem��nS-G���&������ʫ���:��������&^"s�X�Tݏ�Z���]��9(%/L��R�^����ۅ�<�n�GbEi]�����/��(�Sfb��35T�VX�ʣN^P��xd�Y�ub��g%1�l�2"+FDMF�^S��\���ɷ����J���u�Om[ۢN֦V�ysE�M^�6�،�p���檳�_#YZ+!
��/*Q��m�kj�kmj��P�J�(���8����+ܦ��#���cdKU�����I��h�[�:f���R0��f�ܻN#N�WJ�Nn�!3Aʫ�]������*�-�1����͙V2��/�F:=��ݙ�F��y�VNT�T���%h"����^AnE@�LKz,�����uV*,����Z�{�;ֻu����3��a��^�kG2D+$ߥ�y��X�Uu�S�E��j��i;am�bQX�i�&UТ���%������Q�$�nBj�5�eY�S��b¸�+t�4���J&�"Z��Vٷ�Lv4��bL�Ib�oQڰw�;+.�Y�|��ݽH��S����4��m+�	�����cHG���R
�An�)����1��X��q16m�-Vmӌ4k1����:S;t��w�֝WY�A�ŷw����)UV�L��1Z6���C�֡Wz�m�!.�8�f�iA�9�A�e/+ۍ�U�Q�齙�U���;��*�j�f���b�HG2+V�)9t6,����E�`7o2f^ҳi�ߌ�t�Qsiؼʺִ���Ђ���D���3*�ء�Z;�reT��#ǴB�m���'hH�5p��if�B�G?�e��F,j�`ֶ�pk�s-UCy��k�ʤ�U��Ym�;������]jo^��ݴ���z��F�'����MZq�A����n� ʰ��nXy��Gq��UX�{�m+�p4FVJX�X'E����-%VLße;��Umi4�tm�F�]����L�x�'e����ʀ���+�M;�QT�4sl���)�q	�ǁnY�B�ѡy{���h�('��`D�b3��	FG�Ў���/azl�T�T���n0n`uj�Vݶ�bR�IS7YN�ӷ�B�wD�ޙ�6)OoX�Νd�r�3#�2K��r� �X���Xګ/�V�
z%Tn�L��Co�!�d�A��;M�[r��ͯ�V��'*�eU�I6p7��`�
<w�h��:���*����Ϩهj�;�0M`���Vʴ��5���l�W�F���<�+%^�ϭb��H��$nnҼY�`��U�U$�uk
�$���j����&ʔ�=u*ۙYt�n6��:��j�#lVk5Z�wo-,ʛ��!�DŹ�1���kU��u��;ua"�w�[q�[��*�N�c��͢�ܲ�F�������ѭn��#u�0�U����
�*��)��-�SMK��؆}7'� ���"$[C#���]�	H��6�ǵ�����Ygtm�om��ܗ��f{�Zjc�����	^l*�\IiJ[J<��C��ʤ��K�!v^:�J�nU�H�M�ȵ]r�A+ʗ{y�E�ye#��mHiU�uVZh^V�B�+n���-Z�.��Z��'K���4��e�(�-�享��+�:�j�lH�yjK�9n����Y��=�x�l��&VX��;F;ٌU^n1���ғ	G�Y�6��[y�F���/����`�܌5�a�x3(�+32,�L�4��{J�T75ϐ���9G5i�f�S��7��p�ɗ�x�܁:����j��WY5�m�e�-��Hb���p�2��׍�aR���=2����.��-�h��1����L�p[�0CZ%]ic8ʾꋉJ댋,��V̻)��]��m:TJ�V�M�ؽMɹaY5[�-`֦��N��^n,W(k�r�YLtŋ�VY�7�7X����Ӓ�䅆��6�e�w�6�3�90V�T��ܼq�Q]�ڽ�7���yz�X�[b�7\����G���CYnmՂ���P-���K�Ue,���%���#e8UU�f�=cr�!���5*��Xi�G�UJ�bQ5�v#�;�·kt�HZ^��{yA^ї�c�Ӗ�����̢)�U�v�7w����TYz��Z�泛���=��ʩ7 *�wG5�x��z��I�M挼���l�,��#`��/Z���\jہnI���̘�!+h�h+U0]jT���meU��`�w&�VP�����xF�sk,�6��j�گ�	L��t\^�=x��r��]�kn4�j�s.���&��C7�%d�Skj�Ci�c�ņ��zث�Z3jj��O2"�a�k%�\�0=7�N��7�-�H�75��)��F^*�9�Z�wvj)76�b�D�(i�,e���nA��KwY�Y�hu6�Ju�B�mT��^��Ť�%�Kqc��)�*�����*�*M��)�f��gԖ�\�	��T��N�tU5w�ҫ��U��Y���5�ۼ�	J�'5�j;��r�K4��J��Õ�q�Z�ڭ42��a녒֗�Y7����3��kEmhh��o#[g^�efC�n<x�@�L�x$V���)1�˭�bSr�I�K��˻ܽ��(����i�w���gGx��4R����݆�{������Gr��yR�{���u2,9�F�pefL��L���h«V�Z�1M
Re�)�t�J+3&=�<����H*[
�u�-e�E;ۙOl��u���p�+qޫh�E[x�)"���Z��f���
Y3m���6^���ǹ#�I"J�T�'ɭX�],(E�T���6tA��o34L[LkȪ7�Iy[�kŗ!{�����@�e�+rݛ��YlаA�H�x��e\�lطgq�-���VMiv�����.�kdB�mVZ�'M'f:�[y�f�c�A\wr�����ֹ��3-S,�F޲���m�yu�A�۷z�
�ܠq�x�ʶw2��vn�f�7�mG	IP�����k�F�O������f���bk7��֊�s%)+Hi���͠ꈢ�?k���4%���MZ��w��Et�c��"�U�ٹ,<�oLnM��[Wy�۬a<��K`Ss�f
v��	;�T�C�٢@�G�֠t܎Ԃ���E��z�f�%^�Ұ�N�{`��un�]o�Kt��^�F��X������Kv%;ZU����S���'�miH��7��H�V��Јm(/CV�G+3�k]��f�h����.�v�n���;���Ta�{Ur�3rM!�-���x�~b��x�	��W�k35��
*M��{!7pU�����B��E�H�w�Įik��&���n�آ�ʓU�al�w��bI����A��IyuiL{���������8���t*��'
L�K7rJL���rZ��W&����5F��[r������ض�8�,Suӭ���q,jDn9U�H�N�����e[��RU�ɴ6f]�$��z֚׭'�y��P�����V]�:of�_,�;2<�m���+nvT;��l�EW�]XüY�*j�%��=8f��	C�2������ҹOi���͗.�1�[������$(�U���
��Yʰ��)��Ř��SB1a��s2��/-�*�ݪ�0Z�D��
��qbq���B�=�4���Z�Y�9�{��L���lGj�\1fm÷.�^
�^;������J�̬���^m
eTI�k���F�l�:拳%�/+w���i,�R��TMҋ��b�U�;z�y�[{{���4Z�MʪՋ�x)�[n�&Y���u��*�x�j�{��xq�ܲ���{�*�Ҫ�t%��kH7��1,q��7��H-��6�fY;U�5�{��%O!��,�,]��kI ��M�gMVJj�b������Т���U\V)�c1Z�?SjQ9l:$3�A�Ú�!{a���:7�F�ٵ����6���4VPaّ9OM%w��^����<sN�TX�*��m&V�!^VX��|���5��ʙ���z�ꖖ!{xΡ���4�Q����I`�vl��y�����5�3v�ˈ*�ח�k�����h,�׶ӄF.+8���;��en�7�
�11e���ѹ3i[��v+�$�h�x�B��V��H���6eͲ�e蔵K�j��*,Qjh�ڦC�bON�B�[�e�]�nW�Va ��̔T�l�"�姍+��m�x����٧vU1K.�L�l�Н�+'F{f�YXp�v�c(%����U��X{Y��EkU����I�9�͸Pt�[T��Z�}U{*�%�S7f=N��yk6<����޶ˠp�T�GI4�X�d�UUUn��_I��ԛ�C�v$�*,�l\s.�x�a4�PC"�Ӭe]GqV5z
ͦ0f���v��h�qM�M���uu�P9����[����	��7�ơ6�w���S-��V��U�RQnU�7iJ˨wq�2�6��t<��H�����p"h�4�e������zCY�B�F�-��nU�1Ej`�N�nګk>�Յ\�`ӧ$�L[�s�K[�v�Тܫl�Di�2��ȍ�t�J�bOn��!+ĕV����E1��W.��j���$�[40�J}��V-fԟ[�R�P`8oj��Ѹ��^�۱ol�m�tj֬�o^�nf����ݥ�a�]	�(���cTx̫Kٶ�V�W�h��gjaɚ���3
��k	h��{�/�osY����.�U5zb̔���̱SA�L�xhZ�,TGF�SJ�u5�2�ZtJ\b��օ��wW�+,φVd�fi�>�N�U�V���f�-���<�K4��Sv���?�Y��j���V
�Όț���w���t7n�2m뽢J��B�:�l��M�)�Q���z��A��6ЮJ��Z˻��mb����1X��Q����5r��ߛ�?P׹�׋iI�f���"i�Uh�]�m���z��Ź�Osj�;�]Q���UkU�i�"�#+we�n��%�9e�o(�7T����t+D��e�ʟe�T���&ɒ7�mJu755�
اq8ռ��%֧y���7�����ĝ^��k*��2lXp��f�XV�Ukš�n�J�jk�v��]h{h#��Z;2�W{11RVPڻ�wF�j�""��=h֕U-�`�n�,��Ǩf���҂��%�u+7sqQ��e��fm�z^�	��؎��(\���Vt0��'�[fܧ`�^��uq,6��^T`��,������U��/�p"l��J��j��7w2�ڵ�Kڭ#~nL�Ɯܪa��ˬ�C
.�2���m�U9V=�ފ��t.��W�0��J�v�Լ9�1 �1�Ma�Z�&��auJ]�T�0ZX��k^�.�ǰ�/+w3nd��bm�[���Ad��*eSY-��f
Q�gXt[B�n��C$�,���U�����XB]ǆ��ޢY������F��U��U����3"²��b3C��Ȫ#�d�uF%	���0Y���V�6�1��-a�֕V$J�s����4[�����]m��*����i�jd:�u-�E$���.���ˣx�:�R̓2e���۬����J!�ЈkRx5y%�t-���Z�`�t$m�ه*&!��zӴ���M�~tq��vB��p�ʴ�+������YzJ��ݣ�(Rʻ��ͫ�Vvo%��Cz�(+��4me��A�Ayb��Y���r�(]� V�fq�	�)ٕ� ��p�LmH�w���\�!A��m�V�HSu�Ajͭ9U/q۫g-�j���S���R������'-	����H#YX��Y���H~��V��⽳-=כ�BU`6iſ*ʪ�w�x�=����8����z{,j�vԣ�u�6�L���!0��D����N��
���ӵ �5��q��T��n����u5fL��*P�ܳ�b:�VU�eޔCuX3����'FD����|N	voj)v�!*��x�7a����aa�(�1V���U�TnP�F�Ղ7��D���x���K���m/�⺃s\V-*��rR��S��J�An�ʪtd��28�F"3qc� ���{��k3X ��3O^�Q���ӹ�XS�$ޠ��Ս$T#X�:kX���B�@3ʧf픨X�^c	U�;*�ue�4m/��W0mxf@�uVB�F�x��.JZR�(\��i���م�l5�)�C�Yj��&�^�TnY�^aJ�:��rVE�ne�v�*��>V�\:�lڷ�\����e���a51��ֻUK$�N�꘯��8�k2GN�m�3!rRˢD�dD�KU���f��Uw0�6�֖��l3.��4�F�R �IzUMȒ��ӹ���u�jh�����ݻ�Е�j��Zȯ�9c*����ۺ�-n��G5Mr�*c3-\W�^Q�[�S[����]����iVQ���hӦ�Wv�jw0�,��%��'/r���K+i���x�]�df��U�b��K�X��6^���:��i�]Tj��KA�Эͅ��h�<�j[�Vy�S�uF���ꪫ!X�R�N���Wyn�z͑���ŵ�Ff��4Ea��Kj���ͧ�e�R[ �dbL@rn��7I�ѷ{�-�3t����4��0suR̼(�61����^*��Q.��!�F֋n�*��Z���GcV���u!l�jRPZ��T	�r�wJX0=����V����[Z/\�4WW2��ڙz��5��W��$��(U�Ǯ�ِU2A�����%���^h5Vڂ�BfB���˭��̂�*w��i�Xo1��f?��������a�[y�yf�UV˽�W{��w/+!U�0�1��W3saT����Ú3o2�@y�M�@�!&�H@�HB:.긻��;��껸�.�������ꋺ��㻺:룺���;�������:룺讪�����;�������.��.�����;���������躺�껣�㻸�;����*�:��.��;������:���.�.�亻��ꃻ�����븺����.��;�����븺�.���;���:��:�����:����������;�*�::����������:������������ꋫ����@6���BG���%��?s���+�XhE�t�~cI��W�1r���nٹ���oʄ�)6�,��m,���e�VL�i�@�۴���Z���n��s��_-�!��]������|ʗ�/K��WrV�PyV�X}e2e"�����f�5۝v<�y�Z�ъp귲�C��M�W{��m���F_<.�􉝎�f������y�T���2�7[��k%mq����vq�9F�W�*���]U���U�<�����#ʏ�v�Y+~�Wf�l���nN۾���T�l�Ϭ����nw.��@�"oru�{�VoL	�yҮ6;�vv�FL�j��+)�T��h�b^3-� g7K�+2�����y�&�]�yۼ�RԐ��gr��-t/fT쉭R!<%"�XY��n�$6����2��ؼ����w�&�V6aS�gʰېG�EG��߰����ѧl�[���{rY��r�}T�1'nɒ�
.���ֈ�|+zL��]a��X/c�ÉiVh�a��5����{�wf�FP[)$��k�v�/v�@�vbU�f�r���(>W��J���HS-uv��L�U镃��(tǉ>�:�۰sc��J�n}��nq[}J쌇Y���[����X��TF�T@�w��L�eA�d�ܒΣ�*�C�f���*�(�qU�-Ѹ�齄qZ�Z���TK*���L�	�J��^ ��OBۗk�>�����5�r�\bL`�7�̳nC�L^�i�s`Q�LhK�պ���	o(te�W��J��:���Zʮ��y�j���=CR�Y�n�>�{Ъq�3,�𕷵]��BS���hҽx$�Ӥ�l������d�^۩�M.��+:�ޓ�OrN�2���� ˻���B{Oi��FD0��53j�^(xX�TǪcUP���^�<O�ӌdU1���٣4��)��!�;zcoV]k�ĸIGk�;����Щ:+V��[ۻo*����n^u>&N�xpխN=��C�,�R�W��6M�v�
n�,#��v͚ގ�=��:�����k$_sELbY���q�7G/(�bmYѺ���T7�TN�W5X��ݽ%�D�c�y��`���8G�����c'7.�cԅ�|x��U�^d;��,p)ֆZ�]�Ay�����Ⱦ4+ui90CO�TYt.Uݷ6�fu��ko_-�ՙoC���J�f��j��� �]�Wj�����1�.��{��]r��mv�d�e��v�3���53��)���`��N�q��^M$����˽ѳ3h���o]���+v�ߎ�b��:�KTԦWR|�VK�j���iZ�86�[x��w;����GU�w�,V�Cɍg�j,��;CWuV��ӥ��.^��W�}k�Z��V�]����Ɔ����v�wׄY�K�&������t�:b�|v�X��FX/�}�խy�Y$YX�nV��>=wk2��S�E�-�X��PX�a9EU�L껫CX��%�"�f_^堻���L7j���MW^�n�U�p+hq�b`�1���t��Af��ʕ���2���*��J��m��4D�ݩvs�i�ce$���={{��.����Äe�Ɲ v�yn9z�Y�+s�^�+���X�/�=�sS�����t�fb�ud�B5gw��N�v��0�g������@�TY�.⼩�{W�)۸���Z7��:}ms��B��)�I�H���w��]/��e	�6G�jzU����,g��%!UX̼�©�/D��:��y�_*�[Z�Kq��{w�W0V�+;�A�ڪ`�aPuX3�s,����ױ�{�e֍5�9�L��Ct�33�/Y[Bw,����]}[[{�1�Qyz����[>Ǫ�*����.���6�5�ԭ��ųۑ�WP�;oN1i���BlQ���U�ꮛX�w$�Xm݊�x9��eRbtY���*���|�{���x�C0��TA�����T��ۛ0��S*��2|��B�p�+�=�EVV��ή�T�x��1B�щ��e_PY�Qc�϶�r��9}�>;�6�r©��g�
9�trf�(j�c-���֦��XM_#֮64Nr�;���6W^�չ���fZ�7��f�9�Jb�e�������ɚk�[�Z+<9�d��L"��Y�8�ܼ�#��HöYB�l#<�pI�I�^�+��ը�������*lڍ��+Kw��2�M7c�]�U�ݽ̻cf;FP����}��s����� u�K++/+a���Y� ���<ni����T�����Վ��ѝz��o]�b��l��<$��I��������u�mPt]��Z��TEʝf��twhmD�o�%��qѬ�^X�x����^��}T��� �|��MG�;@�9�y�"����GR{/.ڗGe�"f;�­i���<=Hhfﮏ���o0��&��^�:��nK�Ļ�j���ԥ����ݫ���#����ԫxӚ�u��i�ڪ�V[ϡ��D�X�</:�*�L�b$�(���U_Y+4���[�<�a6z��cV)G^�k�)��]ZUr-˨w�U�����{J��Y����k{jL��U�{��`���o)�U�]Y!y[B����5�Veǂ[	�cX�y��>α3/��5�Ӎ�i�Q,˥�Qڋ)����k8k�j�7�B����%hv��b�#���Cw���KbUfy^�S��w+����f��t�7�M�6�7��U��+]�}4l73^J�t�.�8˸�!0[,�Uk�s�^���p(-�kRդ��M��m�"��F�j��������mwl�t�+jn�BE}�o:d��P6�*R�f���V��ZJξ����p�i�ڦ���*n�d�-��w�9��r���n�Z���ޡ�Ref���w�j&��^�����.�m�/��g۱�;���O�BV�Q�ݬ��n,&ژ�V���������Uuܭ��Q�f��uӖ7L���ʇ5%)�_-#;s+7�M��2�$��֧]Kb��/������f-r����3��<KF����Mf'&{�V��Z+�30ͷx��}HnUǏ��ic�WI�	9Z��v
zS=ne�]�Y�[r�n��v>���"B��H�r����v7�CU3�Z��'rm�۽/�i�od�Z��t��Rf�v,Xf�)�0�Z�+�[���T.ճ�O���v�Ӭ2�8*���Z���o��VVqA;��fsO%��ԻZx�N�d�p�ga6Gb��@���к��}5ͱ�8G�=9��a�l���]P(G�m؛{�z6ͻS�匣ARJ��7�4�e�Ƶ���sQ��z�(���wk7��h1�S�N3�1��U���}gU��{��Ӂ��AfJ��ky���ivV¡��b�a������:��ݍ.�]�Ïm%�}43]KaK걛�Su�ײ��]3�#�S�Қ�wZX_�xE��ڴ�S�s.�J�:���˼��3;:�r�f�Ї]|�M�����].�ND'A�K9r�TR �c����Ų���t���7"Y�~R��R[p�Rŧm#g��9(:��d36�z�ne��8��q��J�5Do-V��I*�&Yf��j��-�7�ώu��0�_^��ffެ5W@�VW����wY���Hutw��v�7/85��NR��(�e%n�X���U M�����2�)�O.��ȱһ����PK���)���tC�o�[]V�f���!]OQ0�,ں�X��Wd�)��jf��o3L����F�{�i��{N��A��JC�fU�Q�-��VE/a�Bg%�𞾋XD݊��8ZE�Y���圯�惄*r5�3�w�aj�f��%R���V�⺼�%Ty;�ܢta��R���p����-��Fzce�0�A������fI/l*�мK*ԵF��b�lߛ�)���T��sn����d��K��+lU�s��=��S�(=*I�.��&a�T��ڗ�b.U�&�U�`�U��b�9�N7�F�hՉn�Һ��s�n�L�h��1w����|�nӀ�s�S%�%Uծ��Kٶ��n��]ͫ�x�!�S!�͋l��,�j9I̎%��lԬ7CL��Ǖ&n�u�v�κ��(�Qh7����W�-V������h�d�aׇ+�>��f�=�Cxv9���i�CvJ����Τǝ��e��r��P��/��|-+�1`��V�1��qq�Ă�K�5ڲ�o�|na��3]�0lʾ�fZ�<.��QF]�Y�n�[�f�����{��
-y���R�3!Eu�k՝X����N����p6��%��]�/�y�Um=�NrW��dd�s�����%�Sn롶w)`ˇ0].�i�Ƿ�c�4�B��Y����}Ѭi\67���#��V�Ԋ�5d�wu�:g4d�\��ӵ�7U��f��W`w4��V�i��4�RN���x����5��8vG�n�ʑ�-�pY���"���n�ɘ��-h�3�)�uYo���X�厽̹yRѱ��B^,�5
�ھj덚��2ԧ}���[��&����ѷ�.��U��a��R�`�Vlu��6(�d�ջ)�|,��wD�)��m)�e��Ը*�u:-W,�wT;�L�S�q�������܋!(�K�1�;����׭�����QwJ�����(c0kڪ��H��e,�u6���󷱊]P0ͽ%k����9�3o�c�y��*��6�ɢ�QuC�p���ْ�]�ǒ�]v6�;�Npc6��o��)���@�W�}����ڱQE�$�(X��f�6���VR�
-�wM�w��>�rw۸��d6�+�l����/e]�&��%|�V��ഏ��������0��x�vH�r9MS(ڬ��.b��&�����VB�k��j�E*�i8��B�vn-�F��u���Э��09���![�^�v	gU̻��ƛ�E�<�[W�b5~��p5L[0�k�+q啎�F�ܝ��Փ"r�3cnC.x����{Dۖ&QC��}y5h+z&�rV�x��Y����R�����鄖-��F�άB���m�W�WG,at���ȡ&�\����{��q�wr�z��ØC���){w�Ƴ��i����똄�f!�G�e�z^f5��5wj��3��ʭ:*�U(�b/k8k�����K�k��q�	.8����ؓ�P���.:��5*���!g���G�XY���zfvLU(����{T�T"wQ���T:��N�|�Q��������V�r˭�K�^�'LF��\z�uCy�p�n�@�4*j�C��ʖ2oup�#�ƻV	g)���v�Xj��i_t�|&s��f�ɺ�5�{���'�TJ�oF+��`�T6H�Uq�d��y4��Ν{!���ܡ2�㕑k���W�6��~�=�.��mX��Ɍ���m+�{__Y�%*64���K�˻\U��W��^~)�^̼	�rJ{j��*-��UoS"�(��z��3vn5���Ą�ǑRz�*���{�.�����2�hUyzּA��nMO7xc���-�j��]U*��~�﨑Mk�A���'{[Fd��b��b,G�
T��|{j<�+1�ݹ0Az��2�B�v�]��዆���:�cVJ�;��l�ɖ����ݹ��ɕ�f:����'iU���M�i��]��Gm"N�-+{A�iVgb����GdͶ�d�N�)e�]Z-�ج_^����M��*��uF�Ċ��sS!�-6�s{���c�>��
�z#uR�ۃ*fn�qʃ6faB�,�Ɛ�y������������M^IU��Ѹ����4����O^�j���L��2 ��\V�h�\�uO�����{��4�}�V`!eb�v�$������"���Z�i9B�%|x�Բ����ה��i�gn�_
P�u{��uh��#��.ڬ���ۛY����ި��HNP�k�\�T�Q6�՝c��AC)-�Zʙ��<����S�Ug�z��ӬMۿKAɳ�8am\RUfP���M��ݧk�i�4)�:�����+�U�^�be�-8TC"�k&����*�u!]�^�-�K23�+,(� R���pK�e�rwz[�i�Zr�v�[{4�4����]堹��7u�ꎘ�e�д:�ȃ�6�'ִj>9�16�]�S(��c����%���=M��;�Nv*�m�㩄̼ʄ�f��[����y�-��MȞn]K^��6Ce_���͌�/6LeYdd�J�)����I�u#��s�ݨ��i�E���}Y���s-�w��x�X�J�J����s��^U)7Kw7Z*aL<VE��ml[P���'j��+&>�����7�ۗV���M�V�J��.��ʺ�ٵsT�Knuvj+���S+HoR��Q��Q�¹,��ygA��E"��&1S8f]YyPVr�|+���+�{r�7�wn�o2UfS�AW.�����F���(���|M[�|����ц�����ے���-���w������B�.�/sw6��?'�i�/3qN�3J]UM���ś�r��s�9��u�n䩸�	P,�oJ�J��V�뛒�^�������W��}1�ҥ�)Ѯ�c}A��F�����_!��N;L8S�N����o.��fU5b�i����[��@�C�W.�5xv�x��е���v�>N���].�8r�v�h�q�eg�Yl�Rd_^��Q�]`Yr�(��U�/3��p��a��[�rQ�J�f^��f��]C�2UV���s.1w�[�`m]
�z���]�L���&YC%f�����ڲ�c2��q���]]�'Ћ�4���Z�7}�QD��W�lx�j�'\媙�<H�6�8�[n�T�@񪤭�T�I�w>P<��)gTX;�|C9����h��hvf��W��&*��7o=�&[3^:S�=��fZQ-�����m�r
5]�,b>6���5djV���6�$rT�-]�I����r��d�b���v���^/�TR��r�ߡɲLW������(>豷��5��}���IQ 7�m��;*�:2�;�����0���ٮ�Ym*9���(�5�K��2�`̭tق�v�[����\��MfeG3#�n��J�q���n�4��L:� ��c��k�MpX��u-]�͜��¤-�ݒkvSuɱ�)E�i�Tƫk���X�����ض&)�5is��pF�4�,p���WsY���PINR����	k�<��EsD��&���c��w%6�+�[��c& ��-��60ʱpB�\E��۹4Ѐ��e�Q6�p`��+pi�T�tq�cD�-qe���r���huQ��j�sE[m��4hڕ#.ڃ	��+ih�,�R��j�G�o!�<�De�-Ia6t�cz���{�_��$n֕/X��.�+�#0�!-���M�V��[Jn
�Q�ΰ�g
ʹ�K���*��H\���hPU��&�3��Ū��Rʴ5��jjv����e����+f,N#��`����J�Z[�J���شH%m��ci�`���2k���]kM �tF�\��mXXqB:;#�A@�]�.�VYc�Y�(` ��bm�-˺� �@a��"M����]�%���m�l�K�j�Wq%(����%�:�f�u�m�-݀�pV;i�&Z�kt5f��o�ėk�m���l΀�ζ���b�J�V��p�c��%C9֖���mvz�J�`�kչ[��P���X۴33b��Ʊ&롣؃��خZj�KD��	c�Y�36�E��2����� B�֩�c;v�0H-��KQ�ȱ���L��զvMX�Y�����u�kK�+�M��:]B%5(Z�f��e�J�!76la�����ڹk+n���Ke�l�^�ٙYXq7����5�l*�S�˚+�[[`ff)+)��0�+�RhGIm��_�/��L�v	W��,�=5�%M�3�n�+���z���6�v��]�V��sr���֖��W���6�S�3*�vf���.��`ID�XG:��XFQ�.̯eS[�1)���%n4 ��1@��fTr݆���Ze�bU���MԱۭa6�*jK5"6.�mH6���7��<g;�p-�9�V��[	��z��U��6��U���f�GD�iv^X�1v��6kY��f�4i��t�Q�b�Pt�ZH��K1[���k��"�5! �H��1�#څF)svͬ�V��b�f$3��Y�Р���V,%I��-iˮ�.n�laֺ0��&�)ia��s���T��H��,��0v���F�[,��#�XЛD��V�.Ԗٸ��K]�ae��X�`XE���������ؙ]�a.J�,��8X�(B�K�*�Mqy�j����a�fkyn�ι6*l�.�Hi`)f��X!0�-h��"ˣ]�Jd!�K��ar���])0s5�Kڑ�X�a-�a�h�P�) �iH�.�f�e�.�[��Ы�]��s
Zcmb��k	t4I�a��U�#�9��h��$+�vf���H*Mq,�i��M�l�#�va�-+l�f-gp��jE�1�l6�+��n�˒VT�
��@qrC���6�lTp�m�G(��9��ֵ��;C���j6n�a����jF,+q�k�qc��pY1�m`^��"���Z]vH�)Ncp�,�q��<�gWV]KMk���� �tqx9v�M;l��� Xiu�q��XP֌��(:����i-w��2+���۸�`x���>h�>6놘�:��(�7d7l$l�K�Ѻ`]&�72�oeB��H�F��iK�����ٙXF+f�)���`WK4�m6�JcFlu^
�V4�;j�b�JT�����uX�b�,�:��Gi�@�1n%��1N�a����HV�NQ����Kl��_�\��4U�5�Ύ4��`PL� �eʮ�Fp�X�1KI����&��D �.�L湋�mi���e���nfbg\�Մ#A����\cp7[2���>�F�I.��^�n�D�v�:�idj�S�%�k���̳`��v�D��nk���"A���K�� #uq�(�	����&��WQ�p��m4SL������fntrfS&%�����T�f&�`�-��T�k�n4�r�p]WD������
ʶ�*\��0�v��[��ґ6a2m���t!B�V�U�qL�ґIh�vs��I�\mpX<�A����M��4{)+�Y�"؍m�$C(��1+��h�Y�CZ�[d4X����9�aj*�mɝ���i�`�|���P��cl�WI�e��.X4J�غ��m����K�{첤�%5��g�h3s�+.�[4���$��\"�i�����T2�H�LJ�*�4T!OG-��O��[.9�Y��
!�_&�4���m�,��XT.����
h�n��ea%�X��1�۶��1��2ό�G
f�G$�G&T��L�"�3t�he��jfP�Ib(U��-my9����a�أ�f�p`�U�a���u!J��,��X(�n�BiEٰB���3ڌh��1L�m��c����Aىh6�c\�ү3G>y����V7�h�)��b�
W�.��ɶ�!s5Q�g	�.�iA�i-�P;X.Ĵ�D4!vq�5���K�:�쪙��ʲ�e�*@,h��A��R7F/k���`*�YEBk%K�Kn�M�7j��[Jɮ*��M`d����W��)E�r�1H`�i�w�k7xSP�Cm
]�6�㲆� �chڵ���M��9bЂ�<�X���(6hM���ָVj���sa��lHɵ����v���Ռ�i�A�D����`���X�AZh1)��Z�]f�)�������h�4]e�l,mà�L�(�t(����팤ͪ�h�*�#��lxZ3SE4#��u#D�Y��UGS/b�v�ֺ��e��J�2�����l�`�ƭ#H�a�srr�U��#ځ�h!.p]�֖�M�m�MR��aV�73U�L^��9@L�E�"8���F#�cؚ���S=�H����2Jb��h�!M��q�m�5-�E5I���f ���n�1�4Gm�������I4c6P�U�T�it�\B�J�p2]�Wei�#[���,ҹ,bA�^؉Z\:�9� ��G	j�B]�KA�3@5�V��ʶ�E�m�]-t�R�K�؍e�3E4��Z���bܑrk@��M��Ƌ7B���:G6�����[(�ly�V1�la���f�dF��d%;7B\MRn".0Y�p˕���p�ޭ(9�)R����)��h�Ɨ�-e���Lf��4t���n6�a�0��\Ri�B�M��h0���1y`�m#�v՛�=M�G��J��me��I�Y�Iu�k�y�KQ�H�˯h� L�(�� 	��5�R�X������ՌGM�Y���R��/$�4��$&�:��u�a�Ah�Y�қ�p��@�CDHX�HCGL�i�.Y�D6	Pv��=u��
���2�i�MZqce�6��<m�qL�B�ԉ�٢GWE�8��X�v�(Le�����7Z�M�l�[���IX"h�6kj�f��l�.�aٚ 9f�7V�l޺iveG� GE���͎�*lXv���ՁB��Ŕ��;�d�i��ѩ`�R����/&Kf���[c��R�i�ĵ��]��Ƙ����@ڑ��f�j��+����f\Mb�C+\$T����n7jױ%�f'm�cQ�89��)z�T
�
J��j��`�:��cJDv!+�!a���B����W�����	�1Y�I��)ij䮽nm�����kyH���Kb��pm�B�٭�`v�X�Rʹ�TSR�56������ҦA��$��#��bRl�����k�Z�R�҂EF�cHF��e�;[�K�V���,&5X���fkZ��;�v�)(�\ư�@3jҶ�CB�0�*𽁙%�8ըln�,���WY�50/륊2��e�F��k`�[@R�VӉl��tõ91�!+s��LP���@����f6��֤�%���K��4�҅�ԣp-�W��`t
a�-��AF�P��)�n�a��\t1f�FKn�3XRX*�سM\"WmM��CZ�"X��L��G hh�I�5�-��7L��\�V�šf#Xʲ�W1BR�V��]��\��K�`M���r̶&��#nlX%ˬ��m���hE��P�5CYfMj���un�]��Pm5r�	�tX.0��(X�mK31m�UΉe8��q�9�k1@�U"��f�ƣpT���a�&��k[M�6v4��aK�n4cb#��Cjي�lղ�"k�Bd#i&m�mj�.06�4� gR�c��6�U��l�Mq��ˬ]VW�֙�k[LH`J*�I|_<)�4���)�q@t��y��]4�5nM���*n!9���vt6��2�64�).�h՗ZTMZ�JnЂ�fJ�M	KJ!L�Z��X�6�.HP�2ƈ��j8Yn�d��jW1\�;u7��R�O<ecs�Ԗ�.��̌׭�n��Ěn�0[qf��!�Un�Y�����ܮY���Na�t�icS6�k��i��pkTp���i��ݛ��Si]�
����X�\[J8�LV!.Aqj��m���bh��ݵ[*c	�3.��l-�z�6�.�ˋc��@6�r�ƪ�YJ�X;�]�:���d�+�r�mn�N�0�����j8���I�&.�q�pJY�j@t3�e� 3p�7m�&�G;k�mb�Q\��.mt�&�Z�j[�����í� �.�r��k0��L��E��vc
٤͛��Pj��D&�1�kcI�E�fm��6n��
ѷD&�ĶVcJDɫ�6B�U��T`����Xcv�8m�^x�`lÛ);��`B⻳���.�1\���F8S.��j�2�bƵ���l&�b�A�c4e�smk�mA[0֌�Uh�2�?��$;�@�.���)�C����%�&X;����2mw�Yiٔ\ ۷;�����mF��Gf%E�PGB9C5"�rq՗�z!^ۺ.rn/-"R�;�+,��A"$#��^nmgN̉�Ye�Rq���@H%�r�\�e"T��I8�kqmȨ�*s���g)ͻ�;��m�ⴸ�/<�(���1$�"�(����ّGtV֫"������6�l����NBE��4�̢ۜg���'��[h���v�8����'ye/M'{X�L��@�)8�)�
.�$&�9�C���,�Dt��9�դQ9Ns��"�'Nr�:KƭZR$��-ӓ�!q���H88J;���:I.�׶�q"E͋Jw"�����[�C3mN�;(��ea.N��'�bTp���;����%��8����U��-�^��Ocv�(,��K.�ju�s̎�Ʋ�9��hHX������)vJ��(\���$t�*͢���hie�@�G�头�[�W�������ppݱ�Ev�����h��:�ks.�7e��K����p �W[)q
]�8c�Z�2�VT�!/0�����u��+X�[JՖXQX�k�!Ա�3Bٚ-�"⒖�u�Ϋ57L'3^è��4�{h��$��3��6�1�s�7b�k�A�{WXXGX��m��ka���l�ЕD�h-k��*X���*U�ź�xv�S[7#�񕸺)��H�3�	�ٵ�����t·i�]t��*B$���\��-�ͫ���Yuqol�[�ׂ��i3�X�"C�͛K������[N֩��bm����u�auR���9�(Q�ֶ�3l���;XgFԢ��-sZg�.�h������h����RTPl����Q���<&�m�˩IZ���$\��#W0�l��MJ$if�-���e
%*c���U��cu&v���Z-՘��T2		M+B���/��#.��	j�-\f�#M�%�ɴ�X! �E�f8�D^).a�VV�tDjِ�
�c�"�t��
���B�2٧[��¦`#�Ͱ��8���@4uf4����i�B1 �D�X56+��@��h�\�k��A-�wjSK2K5�t� 1]�,�H��4J��f�E�@�ֵ�cA���	r۹%��c,���Z�ؠ��9�Hŗj]�	�ي�)-N����ц���Z�pdM�
:�k�V���Ԛ��ame��]�� �1�b��!�Va�k�U�s,ˋ�ؘb͎�mo#�M�Q*W�^��]mip�v5�z��	Z�.�֨�ر� ɵ�\�h�ښV�J�	�s1v��s�����"�+��F�I�����V+�k�F�mP�.��:�Y��i�l��I$cq,+�
6� ��+-:Zڨ�mE���0�z޲�1/ EV�-T8�%�m)!`�VED�U�j�
ז��2�
Yob1!Rez�X�A�V�cF@ J�T
%i�������5�A �,cYh��#Q��-�Pd���[J�U�A`ʒX���ʶ�|���?�&���+�F+��ë�Ҝ�m�H�+I��W;T-H�j�t�|����	��{������*ẫ�s6�f�]�����o]y_�K�,�qf0�3���	�G�L�o �;��V7���P��;k��]y_p.R#�A�ڽ<;�ev4��z�}� �$t�/�^R\��x��[Y�d�Qu���&����E��%
2&ME���+��\���a����J���x��]�·7tS�0A�Atg*U���Tp� n��y$`�#��"F�I�zor��%% � ����:k��7}��.R���ݠ7h��[����UU+�_O�K�i2%�`�E��ձ#+��Kr��4����5�P ޠ�=fH�D�=�d�K�8noej���C*Aګ�7R���~�A'�$�FD�&D�#���R���粷K�kk��(�C��AN�\���r�i�����A�Ǫ�PԜ��)h��{��Yg;V4Zɨ��6;��:�@ͫ6/��3�wo:��_����by����gԕC���o����>��� $��d�,y����O��2��+�.���/�k�����E���0D��<����䆐~�a�zs�AF�׻ƣ��{*)��'� � �36��p���o�����dLd�(�Z��u�hX3�~˥=��[�;�Vǎ�~�a�$u�!��x�Nh�B�N�KU%A2�I�%�h�\kl,MH*JDX���J$f����/�����0���h�0�3e
պ�}��gI|o��#ԣ�Z�ܚ�_y�>���O�$�@��l �y��4��ߣ��a�zI��Y��Eϭ	<?�P��:��w�;���� �{� �����l�:�޴���y�w7�AKJ�;��w�:g��N^���o`u�27a��:�t[���Ik�����Y�MCS"hy6�l�̭�;�W�(w�y�d�����3�v�:�C��sv�y���2'0�"IB���Ƨ{���_���r`�6��QA���<��YJ	�20��>X���W�?aa����ϻ����{�QOP��	���y�%���P���AV����h�L,�1
�%����%�%!�8��,�Y���q�6��D��p �ڟ�$��X Ȟ+}�u:���C���1c`s�yп��h���Ǝ��g{T4>��i�tv�Y�=֫�������/�ta��x�Ol龖f��+��)Gta��YU����xTY�#�K�F��������������Km;��p�;�.������C�� A��dH�%
2&������ǻ�uW�"�D�J���g��w~y��n������N�/N��:n��G��� ��~�U���ݯOY�R��=�1��Hk�-U�0n�[�;�kl�8/B��O9`��w�za�r�';�� ߕ�����a�D���: �#�7���E�����olŽ�s}���y�\� �\���3�HAݧkwJ�l������e�ٚu�i��Ы���Y�b�k�L�4���A��O؇%=��: ����O:�J�<g>�2y���w�{sҶ��9E3ުO���Ki"��]��aX����j`��a���]�̺�v��~�y"y���~��[1�P���#�N��2$A|wu��$�yb��ni�gL��%�qx~5ɐ}�FD�?��%

�Tw��_��w.U��!��7`䎁 ��6	��ٕ�*��?�9�Y���!����#c�D�B���A2&2J��s,�4�9��`�b��f횞��{�ղ��	؀by�d�� ���7e�%�R��,�#~���Թ��edɢ�f��	tӽ;\ι^��/����Jb�_V���+Y��k�W��/�Y|�>B��L��-Lf]\:������M����r���(	�����0�6���p�c\�fninc�7<8s3tƘ�aQ���X�%�ح��^�2�	HЮ���j��E�Z@��]]ٴ��"ktWF�l��9�k�X6���cE�B��kI�rLT32ܨa�$�vfa-ׂ��6h:��Z�\�]W1�n0������߿������@%����J	-���:���ua�6�+�/{l�q��y�;��4��$�7�k ���uv��ƹx�j�ܽ�r�����0~�2$��}"3x������n>3"�Ȃ�wN���l��N���ל��=�2$�1�y׾�r�D:�[��v/����$7Z���%�f���{�ղ�;�� ���&H�IBfY��}[�-w&?l��NA|~�0���4v�u�f�=�w��H��˩O���*�C7ܟ�d�D��~H� �$_IuV�qzWl�w\{��}��s�4�W}��=훚E�>���0ȑ �"HǺ�ֺ��m�W��2��)|��T�,FkQ�BS�F�F&�<�^5�nf�Շ�1���~�>�ݝ��"�A2RX2�<g���혳t�u���o/��v�="`�$�0D� L�?����w��i"����m��kƆ���2�Ԫ[��7]Ԉ�#-R=F����=s��z`�{,7TP0nELt2�ɹ/}��w��^�ݑ�SG���oF��u�;o=�噾�B�~�_!���wtT��O1����� $�I��qf�G�>�ߡ����3ޛ��t�������,I�e%r�z=�Ovo�,��Z:�v��r��7Υ�^��y_���sD�đ�>�{��<9�{�W�����Y���q����bH��o���X�kv�tm�f��Y���ƨº�4�&1f�e0��15э.�,>m�G/Eo0:!$rG��m��Y��jΩ�%���'zN+.���������L6��Z�g
^O���\�>Ρs{	~�N{�l
��n?�A��{^xU�u��9�[����&d��1:(T����S�\���t6{^�~:on)�����و.��`��T�L>#�k�㆜��]_k��T�IY��rê��LY�%���.Uv:^{c�&��|�{�����$`ʥ�h��%��N_l�I��;�g�p�9N�3</#3A^��Kվ@f�I�	�9'.n��i��P6���V�~�NOq�����ވ	#IZ���Z��T�	I���"�n�HvD��-�8و��&�M�u�H�50Ҿ��~~����$_I��Y�>��z��K��S��޻9�w[����$BH��<X��>�}L:���E�3�&����\���w�}�ޝ{�<Vh���EG=��w�w>��$�>�Ds��y~�U\^��p9��=��wט���_�F$C�ݞ�X|m�}��r���E�1�Z�|}u��oq���+�u��7���&��>9�y�d����G	��捘JY��4ŷ��gx�b�g^����I�K���a�3{�ײ�F�Ε-*U]�UJ��n<�~��I�M�J�����C�^�޳�{4糔�y��}��$uo�X�YK̖*����Z�Kp7;8-R����l!s�h
@3.Ͷ�M�"��9#L�{X+�v�Oq���T��ߗ��ށ�����I�m����+8Խ�:/�a��{���V�Ey}r�(�n��}Y/�����j��k��r/���'P���ٷ�q�C�5_g)�6��^G���	���i������L����h���]�.{��g����;�W[�����K�IG��-�FX��yW!�w˲d����+�CwP�]�<��{���Nxj������Qt%O\�8z��Ol���{\B�/m�Y�*{hf�!5۳�W[�;gu��Σ�ߩ�_�-�қzT����ڃw*�)�JRab�����JUSZ�no!�n�1H�^̡*F$��Sv���4u�*SJ����aL��&nh0��4��(V���H;�G�c�g�fh�%�r�il��e�-ve�kaR�F.l�^�ZJmSe��4��.��hn� X��B�14!0�R�-
Zkj��(ĵ�a6ɷ[��pFi�{>|6��Jl�V�Y��%���m��u -H����T@�[M&M6��Nm��PG����v�o�j�g+�y�+7�h�g�BWm�:�u�[��������������h���]��{��o�q��53]���q����9�I:y]�K��-]N�����&�����P�z!��)#�/g޳�j�뻻�#{�x��ߵ]��Λy�c��Ǚ׭���g�P�	#�D$�I��&�s����|�Z*z�mg�H��M���IN87����c+O�UMA �ESL$)�]@	jV�:��F�,2�Bm0��AP��P,+��o�%��o����=�U���[��˽���HĊH��1]��
���/��!gp��lT�cE��Z7s3����k�y=���Π����ee�z�ض��X�Ž'����Z����(��^z�h�vU�����_}y���`ʪU�����;��	�$�H��#��V�`���f��W
�eͬ��5�q��_I�?�B�fM�����oO�n����������~��w�Q6�+o$�6�܎�/-�Wۺ���O/}�]U=�ާ�H�g^t���e��6��f����XC��yh8��
h�m�%2���)��)�X���<�E�R�\���J�WǭpTC'0$�D3={�Z+��7/ä/}v����[�I��O0$�X�wP�tq������2e��
�w������MV�=��(t�n���]��.^�e��`H���$�&�9W�~�E�s2�o�yzK�ge�"<��˹�>�̜.���%p�7�.��_a�G�n�;t�ytn�JN��hR7�K($�_�����#>���w�i ���u�׵8뫬���L@�6�{,ࣧ�>O�[)5�+ܡ��<�]J�9(1$̳�AͿP�-��B{<��d���hJ}|�v��*��G	�Rȸ(l�����������x�*X�O����ZT�(�W��uR�or�
����^���Wٛ-f
�Y�t���n�n�ud������`��Q7W���é���j�W��#63{3�&�s�u��������]U�buu�m��ALE��^�ޠ�Z��G�4��[o�U,X�U�Yrn E���w~���j���uSj����v�RY�!�u);�uF�f�(��B�UO#�i�9����7�-��ﳯsz�p�i8�M-�N�Z:�9l�k�bv���I�ѧ{:��:n�\ιұ�5�:�p�	\��ҭ�:��]�n��y��W&���.l�7��~ٲ�*e{�R�SH�J�9WB_�c�G���Z��ԸF:�?hy�d��1C�܎����/ͫn�_|�q��� ���޷0��}�(#.�S�2�V��=pd��M�ݽ���X������[�[�ࠟ�IR�Ί�,pm��͙��Z��̢o
7���9.����{*�}fF�u�J7�y�\��r�[5:���\��V�U[��ڭ��8��ˣ�aČ[N廲ʭ�U%n��*��J�^�Hn�{���ff�6l�ɠ�/Մ�n������*\UU�4ot��>H�?|`R)D8�����rE�htE)�������@(�#���9�	��۝�k]9�@��ȇ�� � 8���99H�@��8��mv��N��Z�����t������$��R)�K.ɝ��q�� �!�3�s�H���9"�. ��(�9�:J8��3	���(�C�	J:��/:��m�H�;:� %3��A%����Ns��(�������E��P\q��Np�$�NN ��$�N'C���6�8�B���:H�('P�&�rp%M����;�"9"S��8�)�r���(���.�H��m �	�$�'�����\�*p��o=��`{�%�#�1]�$��!���dg��Y�۴�W{.n_�H^�	1��izmx�+'�ޑ�"�I�1'���1d�Yx}��/��|*Oo=�޾w�5[����r���[�����Q_;�ZTB�%P8ac�;e��K�b)ۚZ�qh���ƷEj�{��I�H�f߶^��[S��M���W�a�Rk�f���I�	�9C��d�v>���v�1��~��Y������$��{�L��K������$r!$>�6�ZWy��߯:�wG�}r�r�s�H��}$G�϶��ƨ}�]�����m�e�G�</�m�ۑ�2S��ws��HӻĽO�ZwN�F�t��b͋k`N��Z�ѩ�SS��D*$kv��/VV�#���V^c/:]��'�!���}��$`H��9'��;�/��^z�gR��u{\&�w�|��I$�p��wV4f����iؤ�Pd�2f�RѣT������v�Mˣ)�iS���0��$@I]/6�߳=y'��}}b��UAu�Ʒ������	��$Eѧ^���>͍�m�TۯG�<.t�����9%��̑����uq�G$���R����퓧����侾R���$bH��}��m-��.^��>�I�$at��>~��f�E����\�mL�{���u���@IF$RIU�\������y�~�u��O�6��nF=�r/��������a���!�c{,��a�2̪���Yb.�dV$n��+P9`�uv2�e�d��u�p��e��^��\���--6�u�E�l��3A�"f���6#J���i��"[�i���8����:2�6 Ɣ�Պ���f!jitYj��iV�2�J�2��4�k�g,-,���+H���H��狩5�6�iDt�P��&�q�S���)�F�jb��U3��6i���M`O�y	�0�0�v@�FԻC�.�*337 ���j<��f���gϵ[���a
Rli�Z�MqW:�7UC���[�	ua[L��cT��O���I�}"���mu߯%��HVx<tA�N��{0
�����I/�$a�뾭�hUI�ڛ�2�C��3Ǘ]��7��\��9@t�w{��%�+:���	#�I�����o���������xfɗ�����!$�`�L�Uʪ�ou���s�	eg�m�w��~�R%��y���wx�r��	�H��9������k��ܥ[ڐ�>̯nΊ�u��
��9#)���7٘|(򿏠o��M774Y���ܐ�˦z�t�@�Z���k�ٶ
�L�Sq�����H�F�6�������]�/��)�O��7��$bHĊ;�{�S�i�ڈ�^ZJ+�3	�Xdc�L�.
۾�7vVAtΩClPׇ:ÏK�_C�9��eR�B�=0�UG`o����j5?�������K&�[�o�U߾Ϸ}��]��V�1�)9@��w)�
IH9Wߵ޻�߳��� ƀ��H`ze!ZhCRKXФ���IHj�M���{��\y3��W������}[��߷A�B_M��g��hRJ�Ba&��$�4#|��~�}���D�R �n��`���0Ch�P�{�;ϯ%�Z���;߱�h1����B���{_T�}^uy�cB�4&�6��;(8І��@���Zm
I@{���cϫ6ο8�i�+H
]����U��ۼ�u��V�0�	�@�hC&RL��[4�$��מ~�O�����?̀h����c @)�u��-�Hn�1/W �&�E��a����$�קK({� ,�z�4)4`�IH��ο��{����uu����4#|���y�^�U �h��=�ZcB����I�IAlII(�߫;���m�nP��J ���9�J�9��}Ǿw�y�h1����B����X4)4 �/��>!0�;H�̔І��i T�ЋhRJƁI�p�v�깛�W8��dW_����{�g��[8��I�ߨeD��C�9�"��neI�����h���<�&t�W)�on��}����M����~�[�p�t�ĔܠVІL�"�$��!�D��,M珜��^�z�7^=�39HV����4)4�$��˾���w�s�<��ޤM�hF���u&���W<�[B�2����sH
LIBvP.d��S$��}ن�c��V��~� 0�~���/���*�����A�B���hhC3�`����1�������T|q��=�tU��k��Nͻc�i�l)i�`�]�T1���ˤ�����6�� �HF�����I�r���n��}�n�9�� 5��1�|���}��A���B��"�
wԂ�!��% Zh	4l	%
ϯ��_��R�^������)4�R�/��������s������1l��RhF{Ԅ[B�P���xKy_|sDB �}���-�h=��ZhCRRL����I(�Zf�ߞ�}>׎��}߾�ze�W9;� 7� X��
Ƅ<�Z �@m4!�$�����PZhG>�;Z}�{w���ei x���й2��І�M 5�s�Wu^����6��� k�PcB�I�cB9�oZ�P7U{�ݚT�v�Y������<8�K0u��{�Q�}��S]]�o�.�>�K�ʸ���wu��[)|���k�7+[�ލ�P����@%�~!���H-�4f~R �H�JB�hC�X"��e~c���Yoy�~B:=�R����>�������uu����`І��h4!�{� $�&�\���{�Y�ۭj�;v�Wc4i�tn�e�2Ŵ�`l[f�u �&�eJ:�el]O�I��I}ܠVІ�)�`�� $�W�������L�n��߼��44#���t��^o�I� ,�v��}�(hCa$����Ƅ0`I�TЉW�VvW+�Y�!з�PІ�&��{��}�{w�o��7���� X�	9@���HE��>oZ�'�Ǫ�"����ɠ��6L�+hC$���I�(hCa$�����j/%��W��f\͝��� 3���h�z����iI�I(,hF�����d�}���R ��!`��H-0CMJ ����޻~�gJ�o\�{� 7�4!��ԅ`Џ���W]��Z��x����rJJ4!�$�*hC$��[B�P�_oϟ��P������%M\����m�����H��V4"f��)% ��h�P�������<bg�݃�h~�4?�e~]72p��ԫ�]o%@��nN����7����v�_V�e��{�n{x�7O�s?��I�~���o��m�����.��C6���	���i�([n�9��S
�4.k�l����(���6d��ڬ+	���(�C.oT�WZK��0�R���`kŸ���%Ƌ���Ue����a�,)v�S0qpY��@(��Ա���i[5Ѯ�N�B�R�:YW�BR�f��f��ف[�FS[�͑�z�u��C7X8`�*�t6��p���c?|�����\�B��fhk�R2�f]X�JUF<k�{d(��:H~$�%�`ne!XІ{��E�)4�������p�����w;��s������P�3+,�����/4!�e�Ф��$�c �P[BA$�V�;Z��W:��D#�`�ߩ�Ch�e ]�Ϲo��L�Y���~����З{�B��g����[�y߽���Da���=�&��i Q$�$�84!�	4��a�:^�;��Ͻ^��ܫ��߹��7����4!���VЇ2��Ld��!�I(��$�RhEJ�~߾�~�f� �7H]�5���4,����0�R���:}���}��k�������@�4#��J��_P������g����$�І4JcB%!0]��w��ڞ�$t>ܠW=�[�>��<�����b|�cB]�ffX"����	% 9;�O}4�=�<t�~���ز���͕R��&��r�k0�X�tWm,	s5l���u��:I}�|�N�&�SB3Ґ�M
I@[B	4����z�ڿ��}�g�{��������Y쿦�������<�!�L���1�IHMƄ4��R���۝�~B����P��&�[����o����V��Yb�ԯ�K�53���%�ʮ��ٖL����L���Z�ޟV���ӭ_j_�f�U=߫�$�����#�O�Mi�粐�߸t��9�����[�@o�H0>�@���Ф��}��ﺄm�=�&��hC	=@�����`���ƁI( b�߸��+T)?g��%�P~�RI� �44%��B���HM������Jz9��V�g ��M��Ph�@Uo�\�o�}��3�o��}�����9���|k���\���`���(ƀ�H	%!X4"IHM�39"���~
O?������n���t��� 7��Ƅ1���*�{քXФ��c	4��}�W9�����k�����.U�8�j2Qs)�]0鞵�(Q�Ñ�5�@�]�UWN��S��D�g%�Љ�!0RJA`�)% ]�ͺ��}3]ǽ��{� 7�4!��5�z�[��!m�o(cB�@SB�IHM$���0`I�T4#���NWy�y�4.�(Mi������er��{����9�� 5�(1�h&���e!��z��$�0�y�9) M�64!�32��4!�,i�I�$�|N����έ������n�o^�s'z�pX��n�qh�8*�<n�Xt����ZlV��ᆫ�v��g)�ܧӾ�Ad��v�@�2�U43u�ۇ�������u;	꛵������� o�A�І0>�I�=�B-�I(�iH`J@���}������Ǎ�_(�Ї;HE�� �mJ ��ouþ�=�{�N�b|�`І0;�HVЋ�\�ަ��>�[B�h
hCa��@Zh	%�cM�Ї$�"�������˟B��Vvbz@Uw�r���g����9�� 5�(0�	�H�R �R�Ch�Po;������k�>׳�"ݎ�҆�ck�\ (miVY	�͸[3�����.����*��א���w�B��>�,bhRi	P�IH
�}η���K��m]��~����6v�h�C�΁phC3%�г=@X�)4���$�І�I) x���}����<�9ߩ	y�3(��|�5�Y��=�wϱ�h1����B��3,cB�@{7���f�s�j!&̡�� \��RhD�������1��� ���9\��5W��)�K�w����p_n���P+ɔ�P�I)��P�&�-B�|����'��x	��,��=���a$��>�u���=��'~��bz��1���*hEOnq��}�_2�w/��!gN�n�g0�Ů���k��yzu�볕�*�R���Z�*V�������U��ӓ,j������Een*����%�A˼B?�-4!����$�����P+M�HIH$�}_�?˪�A�|� Z�=�ҽ~~�7S��؀�4�9�Ѐ�3,m
MI�0�Rͺ}�xd������S$�!"�td)�A�p�%�-�
����SZ�T;��4�uz��x��AƄ6�@�4!��hE�)%m�H
+|g/W�}�}���p_n��f�6L���پ}�5�P.�}�B(`����!��% [@I�
�JB��j�^2_fw6��`з�Ml2z�|�|~�k7�w{�߫{���ޠƄ1��� �=�JZ��w��F�s�@S �ܠ��6�I@��JB)��Rh��;������������ݼ~�sz��~�����`w���hC��[B�@PІ�IHh	%���=����t�w=hE�,����I�V���/W�}�}���p_n�,�P+Mz�<���_"C|� �cG�� I��І��R�!�,m
M�Ϸ�7����FR��=�׬�'9��������!�M���zЋhRJ�B�M =���ΙM�u���.�-�)�~�Y4O;w�$t`�`>~�7̙%Q�#߼��hûJ�'6ᬭ8)M����|{�M�!9�gׂ�-彵d䵮�h�5M��N�3]�tc��'��ӟ�����5�u�Q4��m�"ȷ�b�_w�+��5yd��K ��;+���f_T�*������V��/\�aPZ�]��n�in`z����c��
̽��kr,��7\����⫪��`����G��\Գ�i�{�%�ղ�+�𥕉�"6�zkn�J�xJ���̑����U��i���x�v��8^�I��V�՛{xX4��̴-fS��Iv�ʣ�:�ꖪ,v[��)]����^�c����ٛ\�Q�5�{hs����]I��z9�+������mf\~�g]��uǖ`QH��d����-t�E챹e�B�o^��A�2�귻�'��9.'���^��̲�X�������z�Չ7/-q�K��I�H���ܳ�.C����œ�8�/����*��Y�:mB;EC��U�Q�{ٶ��f��]n�����K���*�y�Ք�X���+2�?Z�v�˭RK��nc�����V'&�̽8JB�@��|-
bnm�XFo6�.Z�>�I�y��r���M�N��yyX�$֥l�{~�`t��x���ʬg$X��]�D���v�:��1vY�p��w�J�;��w/S�{z�}3��E��Uq$�3m^\�Xjk��ws(��E�n��X��Y	���*���ￛ���''K�Y�2Aӈ��Q�nR9Ͻc���8�S��8�� �$Bs��G$re�E�Yۉ:t�N;-Ӣ�8�.	�6�B)8mgBrIG%�I�j��;��;�˞֜�ts��	�'^ۏj��)��;��(N��NBH�Hp�;m98-�.#�"R�w.tP8�D:�I�
 �s�#��NAoz�r�)�.^v�:A8��	)%������:t���H��H8��6Q�NJ9^h"��R�$��M�{]�������v��������qPB�f�9�FZ�� ��) �z�R�vŴ�V�Y��Ә�1�N2�aΆ�[nfl]bm�]��J�l�$K]�jƗj�k)	�W,�ʸ�(˦��Ɔ�"ql33��1e�
���Յx:�^٬�Y���uy4Vh�fis���4tR쒅�P4�mn��Di�kڸ��-���$�#F���1C ����t�F��n��TF"*� �t�5l��%�,�0�d&�*h����v��i��.ڦ�c(+N��[z�ԃ����)
�tڲ�y[���%a-�qi�W:[hP��ia��t�e����\�[J�f76iI�u%+b;\hL0�d�n̹�-Gm�]\�P�#]���nQ3��`�JƊ�`3\9���g54X1f�2�0���(mճp�,-���a��1e��G,��mi����Z�֩t�bbn&�IZ��@-��՘����_��M`��1,���U�%s��	�Kʲ��K��oA�+�1�,��\�,�
up0��7:�M��e�4����چj���g�B_'�d&�ج�K��&\��͠j�1��b���o*u��d�<-�Fh]��X��� K���+R�%^R\�c\)���^��j���e�R��YY\�Ɍ8RK���0�Q����ZY�&��l�m��%DM�.˩M*=��������!�\]v�Ό�+]`E���C�,4�S!2KU�1�"8�H�0Tۂ)��HR�k���U�A��r�* )+��k��5�[lЉ���K���a��Յ	y��҅C9fٙ�q����[k��k��!e1�W��Fܛ%�NZ�tV�Il3�2k,��cc�L�Qp��;KRtj�c�[v�^�Gו��S�щ��wF�Ync{u�F@�9hZJ	��[�L[�PXĶ�#n����i&��r����M!�V l4Y@������b�l	ps�&�9�:�P6VX��	tv����9�ح��:�5��]��J$���glV��1��WwN�Ӥ���<!c���[�EHj�B]�ͦ��ٺ�i�a��R��ִ�,�`�E�!5Ijul�cu7;0m���|��3"�]MK5.�:#�1ŗe�c@�J�u�;5̻!�"��o�@ie�	+�hg9�A�Wf�$�U])\���l1�Xe��e�Ԏ.e0(���u��
\�˱��,�A��6�m0 ���f͌f:X�>O���X��KZHl!ƴD#��\+�`�ķ*�l!��(��oW_����hCh>�H�JB)0RJAl�D��.�>o��^?^>ks���|�>�Ne���]>�B�f���3�B[a$������M �ڛ�}�m��!h^��-������o�z��>�a7��_n�,Mw�cB�B(`���;����>�A4eJ ��9�
hK�)
��I`�CB�@P�)% 7r��M�}3T�v��9�s~�������@����*hF{Ԅ[B�P4!�iC �PXЏ��w����y��(�[9��CV���ĿY&J������<��ru.�[�7��9#E���|�,/}���bJ��_���;$5~��'��9'y��-�z����QM�%Q6#C@�Z�6�gY�+��,t%mز�͘��T�M�=5&��n�Wv.s�_K��m]�9�϶��2��{_��}$�����\����zU��5�� ���N7��n1��H���*��(m�]<��v�����P��l{,��gEx���t�g>>��V���xa	 Vw7II*����_�P���r���������t�?����$rG𐚽<s۸��y�v:^ۿ^v�_��o���XG��{"�����zZ�J�wj��_3wۙ�-���>��o��{�cr�fF�I�F>�I'�\��Al�ء���U��r��}�����$jz���_�2��,6�pei�6&�Rg�4*SL��+vQa/.���	i�M�M�D;��0$7N�:}2�~�]r�	]��)�̪Y��,���G"�1��=�]S�g5���W�]���n�ft�n�y� ��ݓ�J��d��J}�^�`w�K�9$
{�s�{���o��<7t�v�y�$t��n�Bt��2�5WU(=l�Cc%x+ݙ:���D]����x�>]��z�+ �g/��ڳ<��.���r0=�9Hđ���N�����WI;�+��MWL�g�\���o��5n^{j����3c $�H�q�#�gǹ ��q�w2gM��s�{�(t���Cw�s}۴�=�x��!ڹ����^��v���F1�mjPڛ�]�-\�k}�{#�Hđ����{��K��=~������ۡ���_I$���XT,�8dk��sWU�ӭ��o�W\���m�_I�-������m{]�����!��I�	"3�f���Vp˛��Uy�S�W!��$`H��1<��[��W��:��G�3w}O�=�ͩre�܏T&�������]V�X�;/<GA���˶�[OCxwl���o9����;�%Xw��:�j�N�B���tt}��.�D�V��R*�K���|N����g�)#�I���Dև�/kS��e��"��{�O)#�P�Y�i���~���}Y��V(CM�+��ב�F����C	��f#XN��ڢ�b���X�zI$}xuo}��{[���I޾�����Y�	<��	#�H�E�՞��=w���zs`���~��VmK�/=���Ċ�{��Į'��vn}����#ne�Ap��/{��e�M�3�a��}=$�I�|��D�>����oWۺ�z�Vp��/���_eO}�w^����᝕^��_��$���$�&�Mc}�o��<=&���{כU$��}���$@I�u/:i�����
i�RXݷe�%P9|����_7w����Y׽��{(^с综6V�Ps���8/%�e����ߏ=ʗH��|>�I�y��`�P�&uttpj�F
̤�]R��]lC*ҋQ��[�k1���q�(��@u�m0,7l����[�c�[nu�(d�p��,��iW��j@��H�.�U��S��&����Ɋ�-zҒ��خ��@Ͳ�U1#���幌CL�G3ge?�e�ω�31��iM��H��ktiu �y�
DAXM�{D�ˀëw7K�a�������S�6�b2�һ��G)��B����jWQi�h�n���
T�<o�^Y<��7�;��z_gY������S��WlL�^��0$�E$b.N��V�}{������m�K��n�[��9@t���ޥF�;~ą�����I�9\�W
��m7��*P�fmT�/<d`{�bD$�I�Fo�n����f��zK
�3����ۭ��>��D���d������G�}$I�EoO]:�kn����xz�m���=���{�����u��jߎ����O~�#�q4���$T�	-�n4�C �^Ѫ�b%t"j�SUO�=��tBHđ���:]�{�~�������f�����$�=/=)��7������Z�2�,��������]��
�)���&��7�3�(����Q���n������]>��#��գ�>��7���o�X�=��ޘ�^�y�byI(��uܨߟ��1�������v����K�J	�7�z�<�ʞW/tbH��I=u�=�]�]7��f��wh;��y���U6��dnﮏ����`���%���$�"�1$Y�<�c��J��_�������װ�{�`O!$I;0������)erf��l2��ٳ��:3���[3+(���2	�I��X����KH�{��������[� �C��6�fc��}$IV}Yo/v��]G��b�f�{��w�ܽ��׸�������3l�:�ѫ�}����$bM�Q������j�o��sn�z$��{~W�]�[2L=��\�k�#�ݩ��hZ��^�A�n����z��Ӝ5���G�2���W���$��f�
ۿ_{"�{�s����?��E���)~ϯ}�7�$u]�G�r����-�vT�ȟVlɻ���u�ُ�t���0$RHyg��Sݽ�?��6�]W�i��y�s��/����]{H$�i%i=7 ��c�.���n�Hl��k�	EƻX�H��%��&�ò-�_}�U�~��_{jK�r�WA���$�]�wox�[�7u	~���S��x]y�u�ӹ�1�ӗ��\W��s�W =�䜵��g���wy����7��$�ĐY˼�/�ݺ�����;5�M����7www|��Y�_�>�����.̷�j_z�qwn����/�S�1<�殏�b��{Ib𻺃f���(l+��Y�G��l��5*��Z;�ge!]e[V�o)]��xX�U���e��y��n�Z~5��>��������ĈI�9/����fvO�2㕓�f�����Eu��<+��ӟ�G����
���WG���s�a0�U ��u�#�U,.����H�b	VѢ���LRZ;Z8�ʻ7����G��^#�׾�+ݚ�K�0qH��3^�
�:Zث�������nߩ�A�z3���	Ro_/��U.����No�ə+/��!�������be��п!����$�>�k�,,�J�*�{r�b�ɹި���羮@zs�I%�'�i�=s�Qx�v��$W�g�o��n���y�cR�|�=��;T�đ�$BI$�����ո,�_���yס������$�	"<%V�K�N����eQ���>m�鵕K"�u]kq�:��WYv�[r�em����g�&��{G>ߖ�=\Ug8>]sWr2]���		7��Q,�?d2Űq.��S8�7F��K+��a�t\ChԬ:�Q�9%�fպ4j��i<M���5�:�� �[ к��fb�`fq��΋ԫ�Di.#6�`����Q	� �4��[."J�v��0t�+(k����V\Cf��b���[�-�W�^oX�(]AKZ��ZDf��H��[i�jڍ�e��H���#>|�?~1-���c[3����t��[ĺ�i��-�D�kg ,ت	Pr�n?��IIWn�ּ���z���˞��ug��L[`oy��	$���zx�����OV�}3R����O�������m�7m��������:���U^��z)$��)W�m�!kٗ6�<w����f����/��BH��G"��8��[c��}ݾ�n�nfw���.s֝�{�ʲ�J��I�x=�9�����BI�x�.�V�7�
l��"���N���=�;������ё]�����T��pD�Gq��v��Ƅr�2�%�|l߾���bH���^V'�ν�ز�R42�P>�T�����;�n�ݯ��ﱷo7�US����~S���5�ըrO(���,.����%���R����cZ���X6�F\�*���^��=V$ ��f��z����[��߹���:�ʞ���H.{0�nz�G��[B��۾	����}��ؽz���^�3l��x곥�1��s�D��#`��� y.��[�!��2�k��󄹱e�J�^��y����	��_I��3�=��c7�F�.t���;o�R�geO}\��9#G/�ښ�)+NN�yὨ4�l*4�,�E7L H���hU����j�2۬�0�H�T�%E����/���%z�\�{�OR�so�{T2��fn)�Os�|�G$r /�7sA���5N?w���+�����jy�\ز����.�7G�����{��1"I4��c��v�Mp���ձw����v�um��U^k�%d��t��.��������]+k�ܳ/��ޢ�RoS;���e������8{3*�m���zί�vXQΗ����'vط�>]�.�
{��Ț����љ{7u*��g�ufM�Yn�D��u36������ͭ�<v^��2�Lsrں�o���0�*�mq��i��f�f��j�T6�*eU������Ul^���VQ�T�ߩt�*qX����7gjH����wu�3ft��K�mn�grMܜ������T6��˼�۴&]���"�MY�/��Q̤vP����u�ޒ���Θ�R��r��칽f5�-Zk�^����c��#Z�Ŋtj�r������޻�78νbw�R�ƞwKTB��xE>Dk��.5�@���}.�<�`��4�����5����n�K�ڶÂ�Pe��������]�C��N��/h���8J+#�/b�~���C&ط^ۛ=
z!.U;W!ݺw�ao6��̏u&�EV��]�r�o	)��%W�Fǒ�KƍfM���gWFc��ji�<UL�v�#WA����Ѷ�dx�ǅv�⼄�&P�rh����aT�A���J����[��Hܳ�p�ܾA�9�1_,�
�=[I&��QX�	��v�6�d��ג��_; ��j}�����>�YJfл6w��r�E�:,��Ev��Jq�l ��nDr���ե��U-\��b]�Q�°$3F���X�+���5�y��n������ϯ����j�Q������H\H��r)��miD�9Bw'��"�%J@S�AĄva�P�I{g9)�*Iâ��� :�r(�\�8	@�	�s��D%�g%)���"E^��'9ܓ�w|Փ+#l��B]�g�$IGC���V����ZqYo�	y�NT�qs���p�=��9'|��6Љ+�;��rQ$��a�ۭ�o���$"s�+�9����b�W��/o�Ҍej�ݝ�'u�kI�$"k���ֻ�ۜ�޾��sw��9#I%���O�����e�t�U����OR�so��۞�5Fb��(�I0H��1$8Mw)��߈@��oZ�����vos���?��������A�O��?oϲ�0�sR;WU�4n�����k����I*h�.�2���3{��@a�0̕�H���6��.�Ӟ�y<.��c;tɝu�(� ��a����A�D��	�/���h�c/ݜ=��!9|�c;�Y�&z��>V�o��'ש�A����WN�����|�;SwF?�� �"J�x:6�������v�u<�/$���&�&A�"$�?��������=S��W�W�H��3��=���l�jf{v��)�����@�|�eC�Ʈh����xZ9p۬s�%�T��cx��7S33ʵ.���e������xJLeH`~���x�ս\�6ϫ_>�;�&$���;+5=A$��2D� �DI7۟���t
��}��k,WwM� �������^�A��2W���4��ꇌ�)"OHjL�\�;9RU��e1l,����2���ڨ��%��%A�?��0D����iﷵ<�/$�����
eqɲ���{Dd��$_I_Y� 4����TMmg��`�&?�t.��.��n�^��x_�҂���$H�����KC�@w�� 䉂��/���)�v��-���Rt�t9�ו�/2�>�L{����2DȒ68vM�����Kn�P@�lA��Uי�=������({��0~7q?��?^���e����݌3%"	��奈0d�^J[��K���1��1;��o���fzu�O'��y��A��0d���Z��yub�خ��x��^�.��/^RufZJ�4�rS�S�!���v��r˫Ăch��W�a��}Nr�g�}�MS6}Ì�>d��@$���i�9K�8�C�fH��u`�,+�!�9�-�e��s��i]uhc)�.�2�Z2XZ��2۱����cS&�P�W�"m��Ҧ֥ki��4*�lؓk[f���\��X��ȨX�X�F��ڪX����^�Е���Jfa�S%�Q�hق���p��i�"�t�I���TH.���Y����w6�v�!��IP���z�i�~?���ɴ՘b�ԚKUth��u�f�UGA��%��RtRi}W����S�F�Dy�n�d��~kr��n��߄�"=N�?����D�F("=�a�w����x�L��^e���ڞ>$��b�7q?�;�	$����2^�}y���Y�D� ��U�~�)�/=�۶�׾򗗙�/Zw</���A��0d��D�/��cJ?�|��%��e$��2F୽�������m�W|A>�L�PEo˒��]�)A��L%�H�2E*��{.������Θ��ojk:���0~7q0;�/��7�F7:�;8�_rC�"�H���R�fҨc�*L�,/]s�fnSK�#i��˴]�VoS��{q2�IV~�'���,��g���Y�2��n`�9쮴�e
d_IB�"��%]9��=gI��<��쉇 �Z�;P�]"��glx���o�K-���Ňٗ�c��n/RE���Ӓ
ڈ�����z��'����=2�W��;��_����3o2���&A��J��WŌ�0O���ޙ���ޠ�� �2DȒ��N#�5��ӣZ�kj��Cs�w��&A�A$����H�2W��ٗ^�0�U3w[�&/���A�;�ꪏ3�v奷��&��	f���V�S�ُ��A$?���dA$�z��X�ڼ��
�a��1d���Uյs6�+� �L{��d�$�q���\��L�8��06��li�J� �*qb�!����Kup�\Wa�i���`{("ݼ�H�r {3S��:{�9	���ҵmm�^O�0��7��H�J_A�&G�[��8G��n�?gD�~|޼��=:�-�Aޡ�҂ ��a�"Ļ�-�d���?W���'�&P_$o�$ct��{�$H����M�[C?]Q;G{�o��Z��[�c�F�L��K<?(�9D��o��Tj�E��0HjQ+�{yW��s����c�9J��a�d�AH�I�{+P���m� �o�"�� �^c��ojkw�l����0A���?[��Ƈ��k'A&0���a�)2D�D2Ui^ᾯ;���#Z�;��=���ܡ~�`�J���,]{��ʿ��Y�Y�)fC:h�BW�r35"�L�e��,FSG5�$�T�j��>�� �A D�|đ���޽^�W����_^�=vo��\A��?��G�"`$A�( CBs�]���1}%9fc��驽�����n�`�7�DI=��=Y6�z{�Z��_��`����d��"X��W��[ڱE�����R۔/��0@>�#� �2D�DD(�h�1u�}��ڂt����n=��]��f���'3!w��ZezjN�8;+���ݛ��}J#t��,�������݃���DͬO:��;���G�s��J�V�t�RM�W��t�?�Iw���j��걒K,c�E2H��̋[3�����z��k��tn��͔3}���&#y�7�Ȅ^�����ג�����5��36Ms�^�X�ŲhdKr���c<�ј>������>�� �HA�/_����b�f�:[r��y���;��;L����_d��H�I���0Ccg��5K����lX#�(
����B�Dڞ�,x/�6V����O�������	�ޠ�穂;5}�B�"H�2D��.��{9H�Gׅ��vkO3��#����L���"H��IfJ�<�&����w9��G�"z�y��W읎�ܡ~�8�P@�uU��mD�����r��"�#��d��$���{͓�uW�"
�e���f�/5�W|A3�a�%"ǻ�����P���^�Zbԕ!�v��M�J�f���=�viT��}��=��t[{!ڬYԷ+n�����~�y���o�A���kZ��TkT��cZ��;��q�
��s+�V6��K+���)i6�
�h���`�Hj��L�C�tkE��t�%��6cf�g+1�%�SK(�[ �fsUr+ڱ�1v��Ƹѩ�j�jVXk��6!�Ĩ��9���[pͩж�2����q0�V���,j�Xk1��T�L9Ѡ-��K-�щ�(3:W0�#�;�7O]������⁢��撍�QVRiae�rJ�d43��(M��n�U��J�fH� Ȃ��^�}�y�7!��
C��n=�?j�{�W�t7�:s�D��d��2D���]�QE�� ����z��;�ue�6���(_�����a�$V='�Z��y�z����D��#
k�a���Aw[�RǑ�z�c�^ ����Gw0�2W��"Hر�[�#��B���9����捺���u��r�y�n�`�<7�.xQ�T4�����fJC���?� I�Q�9A׮�R��ؐ���rc}̭��Y�d�em����J��A�"`D�Z������'���F}���k�$���Vͻ���'QBت.���@�a�M��z��������L	#�$�0��s}ַë�j;�Y��W�a�v�?)���ޫ �"$a�d��ؽ>���PE��]����+�r��e6�bn�.��S��=u@b�;0�Ӡ_�\��m�U�������{�j��ʱ�  +�َs��e�o�����]?_�F=��7q2�yK溄�-B��͆�@oEd�3%"	�.Sۭ.vV�V`ڻ�V_zV{�.2��������a�$_IB�D*�%^Iy��WoP����?��n��9c�Ѯ���W� ��tFd5@���s/X�oi��2$���I�DuV�Ch�`�h]I__�o�޾��{��w��7� D���2G����W}���	0b��Uf�fvR��YJ���nP�tu�k�����i0�?�w��;z���a�%"	�'~�Wf���_2�%�BS����u2�^P�������DI�$L����y�
��6��{�&��6 ����Z��j���y\A3�IX=V�Y�@�~L��A�% ��0��&��Y�~"�u;��iE������1>C�T�6޾ݸ�W�V��GW҅�h#T�̞���n֒�/h5n�Q�;���ef��$M��}��}(�~����ʙ׿�&���I��$a�%"17���'ի�X�?��&/����������~�� �PDl�YHIW@�'�X7�y�����X`�"`�"$�`��U��]��݌7�L�����mTw��+� �L{��%Y$E�*�Ug�CSl*H�E6�.��\�J�0�*�2�
��\d��vR1��OW�h �PD3c� Ȃ��m��>��S!��U�>=a���v�?	�/����D2R �d��FUmm�ܳޒ�L������vk��{=9�۔/Ӿ`�J�;�d���B�%�`�$LdA$��$�q�[�Mq�v������
;�W��|s1?�=�����d��$��e���j�唍�����"�^��w޾�ݾ�2�}@��_����Ք������9�68�UNu��ҫ	�]n�p��v��Ŭ��z�N�fN4i�ݭ�Uo^��8���֝7bϰ:[K<�گ��x`#;�$���"D��d�ۖ�k��U�h��:�i���ڽ��3���8Jws"`~!��;�Wk��L����{fwm4u(�b���[�Z<C8��0v�+��]�{|�с��ل?}�I-�d�,������qpQl�y_bᏆuH;dMa����"H�J��w�������<�o��}��2�y��&3�G�f�g�=f��A�?����9���}���e��յ{s�C3��A�{���0A �F�\�3�w��-�L�o�P���XIg��5�v�\\*��w�������{����=����=� �gr�I�%H���lo\�������PY���T��_o�L�k�`��_>�E��H��0���C7�@���[��wz�}S+$BYm6W�Y�>����Q��_ct�����^=��ɴ���:�;��xc�uw[���2>d���hcm��cѸ04[�v.����;��Ys*�V���uf=�ǲ�蝃��r�,�vk]�Y���j����{5�]T�����Vɛ��s>ٻ�j�^y��	��cx��W^���dy�d�z�0B�7�������j���؊V���))����I*���Pd����\�ň�#�쾴gh�8��MܡS�:��n���sP���)%���U�%;kX䪬�B�=�5Y���eS�-Ȟ�[���r�و�	�ܢ���\b��,5x�&����/���&��{1����e��	�$��:��[O�����!���T�V�lH*{Tr��ۦuV���#:t�h��1=�r����N�����n�n�M�����wvŎ<��7][�HQѸn�o@�a����;�4^ރ�뽛���l�x�f��֎Tr�^��t���d�U��__ڡ��+�$V��o3����P�ε2Z��"��cemE2!U�G	��fU�g���,"��h67��n�n�T��.�Ы_`��v�77z�F^U�N�e���ʾ�g��s,%��hw�Ѽ�W���8E�˘F�:��ʔ���Z7y��JeȇN"��'VwS�c�yW|��<6���'s��5�V��	i��
�L=���dܧ�)�`��WN���D����X�g)��R����a�-��t��=�V��1F}����L�^v�$�Ǌ$�$���쾷d����=6Nq��I)3$[]��C��f�HKktw�����mY9{yz"p�e�rK�U�NI%�nt9ŶB�L���׹+-#��<켭����W�nӱC�+^��ol����m՞מG��qY`%Y�<����r����3�qM��{Ifh�yG=��M�G8��8#�����^Qy��Vp�z�8gkmK۬��m�Y�
;�gy��OmC-�qi,춍�Ok����e�x��;f�@]��=}���rH�]�c�����rږ�m2�9c��!�iIr �K���!�e2%��ك�Aڪ�5��tWT5��.5�5Q%�T�u�ѥ��0��hE�xsb���4�K4���Y��4 �Xqn��jDM��&Ѵ%*W*K�0%˅])X�b��6���#&��iuIa���MvM,��y&p2�gыQ�*@�(j�aZ��n��JQxtt"M!e�J�MD�����nж���3fs�W]it���9�hrM6�a��ՎIH�8����l°҈)�n5+�RB��8�0�)3*��a]�4��L96��\4���зb�:��8�WPP��ѫ�]q���m����#�Å�X)�r��)tМB�]!��A������[���Z�ԁv�.sj�ґ��30mh��F�0�5&��kf�Z���9v��f�h�\%�G�TbECXF-���X�B�l�MH9z���0ڲ�!��TR7&P���.�F���UY�,s�Ɋ���-��1tmL�*���6�w�S&.Rf�l�7V8m�	]v����j,)�ٛ�KE�L�FE��Ա��9ڲ�Q���Fnip����a����hi�j�cE��q�"���$��K��1�J���pٳS�)B:"]WА�BS7Yx�JS[��V6I�lY��iT��	#�fKT]�)v�0�bQ�Ԅ�\!E�Kf��GY��uҚj�ŵ!���mpE�1#h�)���E�).�Wl�۝eo�`$.XLtڮ���d/a�Y�[�j$t�֥�U�(QtG2ꮘ�R0 HaM��7Yt#�]X�ҍ/[������Qvh5�e�v��ےī7e43��u�r[�i]����f��[6�&T[c�Gkm�\�v	��i�jM(�b���jK���[1ŕ�(q��6��
ij�d,�EI{(�lWd��	aZ�0`7[qrG�z��k"��gEh�]fm\2���lS8�Fj�3el.R�emW/�ӻ�&��y�t.��pa��fL�6�ѕ�ݰ�26�-u̶�J$�xX�v���	H�W��bW;jjG4I����4n�R�l	�fi	�A/=f�������p4����z_�yBk���R 7F��f�R�b�$Lڴ3R���69��h�&��].�lD��� ��K(��F8ku�JB���S[��2�+�����Ŵb��v���������id��nAu]Տkr�G�5ɮ��40,�c	�Y�}��=~�����2Rd��]����c�{��۔.��=�-��c�>��e����D�2DȔ1�5y57�x����;��u+Fz���56o�+�٘�#��fJ�p+��7�]�0}��؃3�"���/��!��^>���UY���y�̄k�`�n�0Gu$��H�2R �mԠ�t�"��
�S��oU�A�/_���|��{�u�(]�����p2���VW�� �A$a��0A�D"I�ҽ��~:��9�}<��|wL���MM�����3wr�HA�'�ܟ)L/RY�oGX��f�F��3Yi�-�1ln6� �d�6n�H��f����;("�3$L�"u��jg��]�v�%o�}H�UGtWJ�G�*�d�A6?��D�H�$L����=ar-���+k����6`ћ���,�;�1r���D�a����$�,�#�N�Σ�=�H�b��4LoHM�}d�ןχ�K������`]�v���n���긅ޡ�҂ ���3$O��O
Pؕ�B=�r3���d�@I/���H���
��-3�ڳ�X�f����w1|�w0̔�&H�"H�c�Q��R�<�X ����w,IC�ߖ"��OOy\�#}�?�LO���JY�=�/�j�K��H�bH�J���`���?X�{y;�]�S���w��{��J��H�P�Û�ǽ���2J��ham�]0�.ŋjm��(�UqN�ve���st\6�~`����F�$_9#���쾫;�9��/�aZo��X�i��}��< �c�eX �d��$a�d���]��&�5��_?�A˻YE����F�9�n�2���f�]���	���w��})~992�0̔� ����.��B������MƬV�K)|��b�8�v�1+��Grňqg��*gv�B���m��͇u��C�SY���fZ9^&}�K�t����_k�v�����W����AGw0�2E�D�͵�n����uEf�����	#��4_�����[7ە����E��7��ە]M�6����I�Ad�0d�SR��uÞ�m��.l���f���w��@�A$_9#x���Ӧ{�h���&ht�%P�4���es
m�еƴ��n��ak5�J�b(m�������ޯ�rd�$�Ǭ[���<��q\B�P��{=�
���2���a�� Ȃ�$A�"�GxQC8��|Fw/���x��o�:�؋f�r�N�/�����N��=�b��O�=|�w�����&"D$�/ޣ���U�`~����f���8�L|Gu$��0����;D�܍�o���20�;)A�'��[��z���W��e�@���9�G9�����|q�谌ܸn�'.��fi"��r���ky�N�$�����<�DV�:lb�\zY�F����U��{���{�`�%ڒR�%�$���ڒ3Y�q�ޡ���]��}U���q�s ��a�%"2D�>߭�����w����,�]�X���J@c�,%]]�t��p3]V��w��i���G���!"~؂컴tU�w���v�6�����j۠A�r�3y����#�J�	�&Df��u�)|~�vs���[y��<�1w�������"�A�l�`xw�@��A��L�$A$o�$���s�:��払ꕳ}{\?�O�w0�JG�"�I��-���W@h5��LD�.˻���zt^��q�����"�+S��W�!�?������ �$_1$a�%x�Ֆ��%~z㽳�Qo�.�;\�Ρ�=@�� �ޠ�2D� H���X�f��|k|2ݝ�|��Ξ��ظ�ٔ�^@�M͵Y��;&Y���l�^q���k�T�ϳ�k��=PVX��{vT��ص���>yߨK���*u�&����\����#�t�WHL�˚G@���R���U�e�3+M��CWe4Zv�٠�kŎ�ZVaڸb�Wb� �T6��6#2�Y�+4wk�b�Zb�d�鲓G�I�]�l�;/0[b�ΰ���őڲ�l5�(LPu���Mŀ0l���)X�m�J�j��K�Pغ�����	��TAf��F��QK#(ƚ!f���~���n�c5K4���,�n�jX+��R L�-J1�tl�������������~�����1�qm�㇙�+f������ߺ۬�ZS�&rί��H��``�%~����9��٫�#bv]�O�Ӣ��ۏhg�?��2�J�tOY��9{���=�� �ؾrF2R�W�B��ތy�!9�]���X�1w�����$x"F6:C�W2b�ĴG���H�=��*���|��Kȼ~�_��꼨f�������zP5O��?��J	#�,ά��^��$�w���;�y��q��C��&D�$?���A�#����'���Е�QaS\g<h�Ͷ�ż6;�"G-Tݱ۳We�}��i�v��Ie�MP��߬<}�e��j���.���E�4t]A|F_/���J�#$L��x��_"�f��U���=����m�fXW�Ub���YR_T�,���o�;��:�ޏUo'��>��.C{Zb��������Ij�g���Oe��w�Z�o5��eH��������;�����\�!�]w��1@�`�x�'��$a�"`��b�O��B�e�).S����{�����n�2�"H���`)�ѳ����xZZ?^�����$N�a�ޞ���5o�q����Ҁ^�c���_VMO�6PDI`�"`�( D���G��m���a����{�Xy��Ro�k��bdwr�_ �?SϞ��=y���z���O�m8{B�Q�Z"Z�8&0.6%��Wَ�5�2Q�/��~����`���(!}wxO��wG�]��C.���hb�<Ok*����0�#�$a�%|�2E����U��p7)NtL��Ϥ�+s�ֿ\b�y��A|A��0d�_�v��{�F� �w���D"H�rFNu�B.̶:���,�gA����I޽{T�w'>͛zC�~�pו��o��pz��Wx�J��r���t��_d��L��޿~�}�~�����OQ��>��~��fG@�{�P2R��d���0����\⪨w[Ή�dA�{�K��t�n�2������w�j��N�߇������2R �$_1$a�%E�V��'Ѧ=��I�V�M��s�׽�J�NID�N�\ڔ���l�s-�t%�ѺK
�0���ۛ���)
b���XJ�f��ո�s���S ����/��O�fjK}������{\EؠJ������n{n�+����3�HL�2$��(
�U�׎�A��^Z�A�A ������w�̽���� >�_>���&��Y�6�/�ys�|~~�0������c�U��޹/^Wwr�y�/#7�2��?��&2 ��6/=�½JNۧ�  �j���#�2�-��g���>�qxA܎��<���Uv*�K����jﱬr���Oe�HxY0At3q�B��ڳ��&�QW�o*�;RtK{Q6vi��˚(��W[���yªW~���"��\�jg��I.Ԛ	%.Ȇ����\�u����9w�ק_t�wy�������ȝ@I,?��.�[�A{ߟ_[ܬ:���L�Z���hŲ[xE]�`d��L�b�H4�b��;����|��IW�������[�c��.���2�<B]@_�`���Ȁ�[�$O�.�����cw���ta���k��g�}Q)��\A9��c���W��s���-��G|ry0D�A��A$A��?�2 Jx��b�Ǿ؜�U���U���
y�@��_19$��Ⱦ��ΆN�=SO�������?�JDd�߬t�d�V��X��{�0A����V��oY��i�������#��#`�"dIA$�˽g���[�����/��u�D��mp ��O�;����\hi�Y�}�2w V]ױ8�/u�E�r��7�˹�����Y�����nf-�.Z���z+��F�)�j��|�t?�ӡ��>�-.dt˪&&��q��q��bQm[��52դ1�]Qke���.sJcL�Ėh�-�14�T�m�ٮV���A�dfg5lq��Ɔ��Xb].HX�(,�lB�GG:k��e�-��ce��mK	�2� ���`��U&j�1ɦ�F���z�t�b�Z�u%X��զP�j�f��u�˄���[i3@���{!^яh�S����MX�\唄��4��E8��dk"�PYl��0��ग़ݱ՞�?������0��/��&�ٔkӯ����]���������dy�SL�/�@�"��#�% AH�l��9�N��aͤ?"b�c��LT��E����?�("ta�$GW^�<��U�ʱ�� F�0�2E� ��7�1�S�4��x-轗��Ms���������\ ����3%"2D�I�}�C���hi�o&A��^#^�}�7w�����z�}n�$,��UB;m������ �"d#+�,�+ܞz	�b�}�,~�ǯP�e��dL$��m���Ͻ��E7��(��Lm��L3!��#�����LJ3J��hY�������{� D������7���:��R,��=tH�5�dwj�PEdI�J�F��n���LKq�O^��򜺸��vcCF�(��v��Ʌ押`�A0EU�Ԩo)eex��O��=ڱ��*��+_Ooݺ��|��_|�������#��Yd�)h�B}'F��H	�ɀAF2R �d�8՟k�J���qҽ�V?\b�y�.����fH�D"H�è؇+���Y�o����#'/��g�/+#yؽc��%"˯�����{mm�������&o&�/��d���"��O��և�^«�_kJ]�A������?��F�2F6�F��j��(C͊�K�9p�U���qCGB�ћg6��s�qjj-�������U�~2D���2�j��m�\b�y���\���B� ��a�؟�DI"`�֜y���03�����0�YyY��vz�$�Y��A91?�"w0̔=�2X�Tg��275��� A�H�2E��s�����f!oֆ-�l��f;xWweܻl^��N!�d2�-��r��c^>WZ�=;(�u�;��t'5�UmwS�R��]f�/30�]YVR/k��{Tb��}�qP�;_n�ӻC��o^�()��6�n-̾6�"�g�2�����#Ww���)���N�zՌ��D˛x���1xd|�O�8tN�����^<ϞA�i�9�ɣlj˻g�{{6���deK�n�˄Yِ�6�
�+�X�v���C+�V!|����!p��d�w�V�0��s��6�١J�N�ܿ����/bι�Fg��ehr�h�x��Z:�G�w*�GnӛU)��앦��x�Էf�ԙ*�nnwUN#6I��ml=Kr�vM�C����h8�ਔ�w�Rw}�V)�/{g$\��%>�ŜܤVsrcY����������S��"\"����]s:T�|ΪpzI(��ɵSX/ZY*����.�"b��mJ��f;kL9�f�i,]Uѻ�31}ge�Z����N�Um��/�)W�Y�.��S�������N\��k|5K��NSnU�L^��W�c]va�x�c<%w��5�}�|�{8޳o*��k�C��J^�j�d�=���8U��h7l�R�Kؤ7�`F�W7�+�U`GĮ�k0�%�n�}V�m����+a�Xa�b��:���"_l��Πs���U sC�Ue]�c���ڶ��=Ǧ�6��A���xgi�]���!�3qۃ�1����o��Ro3�:�����V�Ќ,~��|��M�O��)a@��	 pޚ���2R y�f�'nm�2��v��^��m���y��mv�<����j��ݰ֜2m�1��[�l�4�[8m,���vl����7v7kmdl1յ�^��^�,���2�Չ^��/B�F��ӫ�z��8�@��X�K,�8,o����ؤ�ZaЭe���-,��Y�qW��lѥ����A��#B�ea �ZQ��BT�`DXy��a3ngyeydmklv�6��2�Qͷ�)<�m�V�f��{km�㌶��m���ob��Y!I�f�S�v���$!e����-��t�~��h���t���g� ��2�� D���"H��VEfｘ�|�������H�$L_�w�˃���m�\b�P��{����Y����H��"H��$L�$A|D�Υ<�j�FC��e�S2�7sY�%"y@^���a�d�A ��J���������X�Ir�hk\XgQ��S%%.]��ٚI�5t�ٵL���s��a�vD� Ȃ���}�����A�����8P{����A�0ȑ���P�����LAL��V��ǉ}.��vW��].�Z��[�y�/'����=`����x��Ҁ�"���瀃##%��`vi�6�kyز�܊���r���Q�?�&D�J��Q�� >�~� ������X����K�W���/]�M{W}W~��
��v�ʴmC[s�kȄ��Sn�t� ��*�Ͷ�_*eDf�19��{3ޝ�k���9�G;:໙u*�.a�捡��v�9f&Niw��c�uLo���{E��Xa6U��7Wٔ7�k����1��)�Y�/#7�2ތ0d�ꑍ�(��7�>�׫�,��1��#4�B�*5�1��X��e�`m���LS*�*���5I����ׯ�����wXW~�i�c�=r�)+�\����O��5ٔ+㼟�"`�%}@�d\��o�2:���߽�:ץ�{h=��߱2'P��uNj����ޯ�:���� ���P�dL�dCծ��b�y�h��w��p���q�f�`�|�F�H��"D3ޝ�]ҳ}�;Ѽ#�G���$b�fg�-�mn�o�'ܯW�q2Kgw�WU�u�( ;��	ؾ�?�BD�0���V��A���F���؞���~�W��	�bd9�K��*VR�FY�4��N�ڱ�r���7VRV��e2]-�eu%�*��jl��ѫ�C��UD��=O�/%��e\�=�G�~l�D�D&J��A�Rn���C8��֗A�ˢulYt ̐ڥ�����@���l��ʤ��Pb՗*����j�(�,T/h`Υf �[��n�*%ql����i-!�L���p0�$����K4�c��j�In��7�J�J����t`�.�+n-A���[�Z�f��&!��4�f��l0f�9Æ<�1���FVa�nf�>}?m?�8E�Ga���t]�[z��XԦ�,�+Ll1E�t�������}&A�P�dO�	�;���� ���-�P��f!�ng��~2b~����ψ�� ��:#��tGjU�`����bû��Y�ǘ{:�)+�_p.����1FE�]b�#��kD�#/���A��?��� ����-1^�r�j�����dW��	ˎ�w�$o�$�(Ⱦ�RU��fu�w�j�A����ȝ��s� ����g1{<+����8�-���r��~2G@��	*ǡ�3N��g1�y���ٵ�{:�-�쯸�D�Fݯ�ݮ�߷ɭ��~��`ek�F�Z����@��t�L&�@+�Mf�t�ZJ ��OWϑ�<�f!���H�"��h�~���u슢<ǽM�+�;��> �k�����2&?V+�d�f�5�R��w�[0(^�S>��M�(�ڕ!�0M������k���M�⣧�u�3\�˲w�d�0��sS������Gx?|f���y[�\�d�{���9���@�|� �0�2F��T3��Y���Nu�F"F��$���jG���ў�.Nr�_x�&>�FE�DȒ1�{;��] ��G;�#v�s�0{���o�D*y�r��"Z4h��!�����B����L~�W�!�[��՛�Hw���sp��uq^���� �j㻩�A�A��d��^t�W�����n�BlR�sSC�(�CT�i&�4�G6�f���kW��Х��Zg���t�]�l7w(��g�{��R�^��7i.+���]�� �ShP; �"�I�	�Γ�>x��A�L��7���w�ꗴ�����/�P��ݛ����z�e/��t(�'���%
D� ȧ�t�]�xs.�b�M�,v�b	Z��w��D����6�T�J���I��*����@�����md�6���e��F��垾��{���T9[ݧ\�:V,�/'�}|��B��: ��H�ɶ=�}��S�7�v������"IA����`}r�-�w\?�_l=�,y�Wf���ގ��&A>��J	� �a�#���`lm衼�k�&
�y�-vEQ
���{�a�#�D��=�B\~��}��=S�œp���զ�v��֤��X:���Q�-��Mk��7޿x�������'ϕ�A�ȘWQW�կ��Ҏg!y<(��}Ŕ�� ǵ�����2$a��: �S��sZ�2��XdLa�FoP�U��;��>��Ke]�N]"�`�ӛ���'�边�@�� ��2F���,��f��xN3�������r����=�0�2J��]\=SP��*���d�� �ڮ�V�o�J9���cǱ��~���)�o^1힤5w2�CT�gQb�����V����v�X=W1-�w�>Yz����q��ycݹl�C�̗-�̪&����>����"F��:��$`I�1A��.�I��B�u�{�}x�W����w]������ A���IG.��0W:}�/�c�L�S-���Wj%�.�,�����4pn�)a	��%�&r����' �y�$xAF���:=~�;,�"��jsG��@�뺖gy�"�%��J�0AD�#�8,������`ܤ~���}�����Z.�^��z0�2G�;�/M��H"=��	��D� �?�ۻAg��u�䝃��z���Vʻ� ��Dt�?��#��D��
��7�q�fhg���=�|������r�����y�븙��}�:�;�峟۵AݤAJdW}^Oe�I5����7i�����ʵ}��r���2�";h#�|��yH-ʽ>��E�p���|v_���F��k����S7p�G���T��\�f���UP�ܡ@��\k&MwW��y�����86R�N�d""&�����E���\[����te.
�%�4)Pn�1�#C�K %�a-̶]JA�қC�\	p�m5\ ��0#��l��F��ѨB�:��:�QGl72�gh\�¸෶�a�ȉk�N���[�[0�b	e
������/)mm+�Ƕ����X��lġ:ĩK��0g7K�F.�[�Ŧ\Q�+�C6�篗�غX�w#7��"�m��;Ii
l�lԌi+FfgVC�|����@�#���$�A������^�#嘼�������r`�<�|g& ȟ�I(W� �����Md'��ɼ<�Ls��O	��r��͎ȭ��tG�����q�i���8��?%
D�ȯ��Vh�G��Nwa�{�/҃�����:0�2G_~��D���z��4�t+]�a����P�W�9�Ţ��F9�w_w��@��0vM�箻��� �L$�ȃ ��0d�P�w@���qi�8NU�.�7�!�|���#�F�_n�u�+ |�Kj�xA��UX8m�1�5Z���Im�2��jJ��X�%hm[���������{�(ș�D�X�u�^����A�su�y�<ǅ����}���A��"�2G_�sxb����ŉ7V_����#z����ٙ�*"s�y*�{��ǯ�/wΰ�C�N�R��̢5#E��xssU��W�m�{v�����{_.��	��������Wu�M�":E��`���H� )�Я�A�A�G���!�{ڶR��`��%��9�����:#�A�#�#d_FS����R�k���(���ȫ��}zc�C���2�/��{3g��Ab��9D����� �����mWzȍ/������|;ְ>���r�^��{���a�"Gn�,"�L0ߓ�7Ł
-�S�A�$��L�,ue�e�2�f.qS2���^
$4�|�#>��@A�G�H�[��G����a͗dV���׸o�]�{�g0���IB���N�"��R��;4��~c�R씃����Z/�r����.� �ڂ ��y�?e�}�__޶�������_da�#�#�l(g���y�����:.r�-i]��(�^X~�k�g@G{ٺ�7�B�[����j�\��𺩈U�nQ=�'t�k�	k2��/����9f/Nb`����	�$�n�2���S�+k.ZGk�|��� ;��0����f��<���z�X�c�YgG�? �#whT��I����sa|m����;��3�ೌ�B��(�b����!���N��a�n���Pt誢�H����"h0�L�d�,���k�l�S�
�����>��~a�$`?��PN����x�W���r�^",��;����B��'�Ⱦ�1�`���>�^{��:�c���=^a�{�9�>���"L�9������w(P2&Aܘ �(P2'�e�պ~̓�+�n��x,�/����P'��ц��FR3��M,��/���ءw ��H�W����Ǹ}�Q9��x~;��2�ts2M���O(���r�W,ǽ�Uk�����X{d�H�B������Wj�r�_Kcs�l���5�����b�Up��Jd�t^?o�"IT2 �	fH����T�����d1_���8nԴ�7���`Io�$�3ݯ�6�ו.��	��H!���A�|���E�Z�c��ME�za�����iTYco�'���~��dL~2'wq]����|e�q�J��@����k�w�|A0ȑ�H�Y�SB�l.M�����os�s�S����+il�ep ��H���c~вƽM{�#ohW�`�#�"3{��Ƃ=�qE{���-��0M�?�w�[��%
 ȾU�S��6������u��_O��0*�;��r����P~�8�P@�U���Xg���J[�sK��D�w�P���U�n�ߴ���P�S}9J���-��W����`����"��<*ז��:8*wk*�{������ޞא�˻��2\颪�^V[|Fޞ�0^�����݉R��%�[���47Z�ц�߅)�Zj�eژ홓�b��j���,]negARa����׵deX����P��W�h�����Ś2c�.��a͵
�	���G���*����
ݨ��r+���	4�٬�8�D+��7���:VU�f�qs��s5KB�����Ցʪ��X�X�2��EQ	�F�&�U��X�+�혣8�v���Rr�:�v�D��%x�j�n��[Ek��9�b�v�Co�O����2Z�+�ĳ�.hN�.P���ʪJ�em�B�쵲�֨7�lH��<�ܿY󫡕3�mGewvO���"�^>,ef�3i��&ak�U���ܴҖ�+�Cb3w��ג�$���^v��j�;s��G�ju1����ё��Uy[ݖ�eiສe6��t���{�VX�9J��*I��1��5�y�y��n2�K��[�j8�K�n�^b��k�uW=�p�H}x&�VI�s�V��A\�<h�tn��huU��i�W���*��L:�3�v�x豃���2ٶꕒ�^U���ym��l�*-V�����݈!������6�fV;�l�-U���u��U��Q=�r~���o�U��6:t� �e�T86��ڨ�cv�'��9E�0ר;�'C�І�s�tW��� �oR�^���7
��{���^�58ó|,�3���Tz��w;<����O��>f+v�V-����fr�,�#�,�{����e{h�m�m��k��i�ܻ;q�ڷ��ی�i��r���-ȝ;�{Y��֐)����xs-mnK�����qk�ݝ��b�m���i���[���ɶ�9.#8�%�K[�u�1�`s�i�I�mke�M��Mmi���e�=�^m�mӶf����њf�f�����N��G:ii�w��'I��m�N�KlͶ6�.ܵ�ݣ;HN�;Rg����E)6i���!��i���k5�ֱlccv��'{V��m,̲�l�^���M�ܴ�ݲ�M���Y��	m�im����u�@�m���f�E��d������l9�f��m�ٲFY�ݹ�f��n�Sb�cd���ܶ�j͛���2(��sV��z��җ����Z�[M3F3v�iR1h]0ʕ*f��0��],"��l���[T�]J��p��i�`M��:��ki5��� Mr$�ѡ��H�M,�bS5-]-ƥz�+�#�\gJ�b�]Q(m.�#	�6�ʸN�4�T�ٮ:)�Pu
�J�l�����H7����lL�4�t�#�l� ��e��a�&�ږ5VY�u�!��M�v摽���l�f��ۦ����e��K21	��%�@,tyi�#jXaܩ Z�\/!CM��"GKN��4ccw\��.���2�\�&��1HLh���.0�h�]�G����0� cR�l),Y��(1�s����Hk�\)��e��SK��Y�]D%�0A\A�]u/h�7�����u�a�&�bˢ�z5�*lC�P��0�ͥ˝�+�l��j����
�ym���Q�����]��rŋ1sc�\\��4�*%��1�K�ґh-�yJgGŵ��BV�+�%�Ck�	Wk6n��G0y��M4(<����Z����gh�ԋ+��a�L2�cv�l4��&a�T�k	�le`u�ZB�;4������6Q�/R�JUN,�u��$	e���/=�M(��a�\���E��8�4�+H��ٗ:\�Z�Z�c@h�Y��a�.&^���.�f��T*gd�M�vG5��K\�D��T�%�%�m�x�ݣ4��m�]Ll*4N f�E�cP����XČ6s3��&o)�l���\"�e��_)��i���\�x��%�H����Tԋ�M�l\���G.ШM�L��!�ds��s�l�Ylc��Q���K7SgSB��K:Q!`�lƸM�I�S]�l���թ{ѻ7mv	v��mqEt!�6m��SG;b4ci�pVi�#����+�č�[V�l��q��iI8��hh8��ve�ΥFX�Z˦���N�5C<�GQ�t���Q�KR45s� ���lS@�36`�I�*�"�6T�9,����f��v���\����r4c����.f`�6�v��p�f��H�T)Cۺ��	v�®�q�#��Z��¶]����˒NI�^am�e̬4�j 6P*kR�5 ���R��s�ͩfĭ��D��e��� ��.&Κ�)o�#���-ې�1�fn��i�@����9�M�Z�.�M�p�,���)����`�9�M�� .iK�������ߡ>���]�YD]s+A�]c�E#��E�"��]BښZ]��T�,��k�~�
^���{V����=����z��G:��{�8!+��u^�ci��ɀFj����JdL~2'��*vz�{._J��ΤA9���Z^����|����A��a�#�Iz�8ꗫr��0A�da�$o������]�fl�1�_����R�^���.� ��@Ș"dI*���Ӿ�7�׌3=ξ �����j�|=7���Ag|�������5z����w�w�|E�N��Y��D������{��������׸��ێ�ؕ��U�}@�|���D�:$cU,醼,�K������X4��"���i0٘(p�d��Pb�	��v������O�/��z��H�:��7��n���S��W�>7��O�S��a�e��ɂ2/�����w��*�o� �n��8���.���o5�Hs�򕬜�9z[�\�eo�֝�I�h"�b7ج��5���˷B�𙲗�f�+^OY���2�|�~��������s�ܴ�0M�:w�]X�h��IB�����0A�P�dO�2*U�S�o*�;uU���+�/����P&��FH��#�$l^�w d����: ����$�_:�����n��]��x��_fu��9N_3�9Ծ �zWۻl"da�����4�^��a�����{�ܸ3��8 O�&3��$�%����ܣ�F��,Qn�U��m0�L-pL�*,Yk���6��@a1�1����.�O�0F���"`�dO깊���+��+�/����{U�UW��X��A�0�&A�u��	������L��ޯ��#'��o���������@��1_��T;���,��=��L�P	�@9�G��J��W^z�����wVVp;u�_�-Z�&�^�Ԯhq�3�Tqz���$�%
�Y��-Ҏa�5}�wh��r�7ݷ�clw�bN�+Y.�����Z�0Kۃ=�Ag/��|��0� I(P2/���ܹ�U���`��_�P3� �s�Ϳ*��+�/����A�A��
�վU�߱� �<�"G���0�W�I����ۓ�x��w%E7ֳ���'"��N] A���(Ș �mSnP�0"��4�h�L��K^Y��(e�62��61t�&�VQ�X�p
�c�D�1׾��k�x{��c۠��yXĪ�QV˯G?z0���+�2&�f�Q�u�{���� ��N�c������J���*��A�A��$x+^���Ud3Iۃ>���?�|����?�����J���T��lٞъf�=�v��]����'���+�"`��0D����-�pOr�;��F�{y���Ǉ��=�8 O�/��KI���W]՞�����i�s"����
}}�����O*:QU���A�Hr���]����ShꩻOD�m����ܛ`��zP�dL��0AJ�E.�C�������jS��������P_~�a�#����Q��5�Yy�Z���@%u�L��d���R6�t��/Q��nˢ�G�Wp	��@�=dH��H�
���^,��o�{k����}dT�W�f* ���Q�_3"dI(W� ��D����[�kxx�|A�s����w��}}�jb|�79������2:�cڌ���B��0A ��F0Ș �"����k�x�-w�ݍܽnv|e�s� ǣ���D����%{N;��xA�`{���1UW�T�[�Lu���E�A��'�����x�s���7�k�����#d@9`����g�jMg�:������C�Ϥ8��,�	���}�a�#����)��..��fNՠ�n��U�K�̉�챷VP���®A�f�͘��̌c�)��W�m�4v�.�]�(���T�%�S�p'�Xx߬n�v��s��,Q�u��޻�\��eZ���3ʈn]v����C���"3[ii��E��	���P�M��Bn6�1�=���X5�VF�P�Է�vR9I�Z�IYt��K��+-�6D��nE���A�%e&�*Gau��ɪ��m�X�B�5[{&� .�
�uQ�Ų��4t�+���b�p�de.���	�pF3��|���B]��ݶ��Y�#i�x+4Ga�cF\-�8���,m�q�˺��|b�0~�?��뱛������/����>��>�����U���"�o��{E&w��}�j�Z�/J�&�w*����>u|uE鵽�[��{�A �H~ޏ���Ƚ��� {�|�F(}� �2G�X�}�"�&y�[�Vװ��$8��,��n/��r���$���z�<�\�b/�^ �����ȭ޺��}^�B�xP&��T�|��cOt_l���쎀"D_e�{s>�U=��+�+�^��]6��$�7�� 6׾ �=��"���;���&RT٣T�����4X��[v�)6��Uk6�W���a(�XjE�;����r~��`�D�1���^�~<=��m�YCf(w����j���A|F��H�"`�L��hnz��ݩ��g�]�7��s�?Ȯ]�馑�X��J��d���n&��f�^���h*iL��w���y�e�r2nǲ���⼊n}v���'��뱛yϫ�]��U�}@�|� ���2Fd��#����F�Nt20$���I(G�r��Ó9s㸫�=7������f&�s��dL����){4;[�` ��=9�#ח�}J�|._�똃� �g:!V�΄��^W�x�[���dL~2'��%}"�9^���@����y���.���.�0@>� ����A�u�H�wue{�|�h@��)j�aan3[,��h��E�ɛ�V#�J��B���e�|��,����>0��1N��F��2{N�[��/|FH�ߪ^�ɐ{v��L�dL�1@ȃ����r��(����,#%	�ǳ�^������8lL��#u��+8���t(��#��&"IB�2&A���<e�PZ��hm^ou�\�6��p��kK�6��v�ۙ���UWJ,{gHOM.�߷5�<2ȷ�M���p�o6u�����#��n���U�P � ���$y��`�c����"|���F#|��I(UU�����Oi�+{�"��'�N����̽wc�lC�L��L�%
ȃ��`�E�o9���Pb�T�^��ߺ<[tp��&A��n��wXɖs�;�����^�}Xj��A(3M�m4�$Jay\���v�K�L��,�y�XLd�e{|����8���C���(�ȝթc6�W��E/���'��]����V�/�P ��0wy�"D6�H�`����#M�!�K���é�-Ώ{�%�]�ؘ&��̤z,6��-e|�iq�	� ��2GD#�t�u���ӫ�_r1�e8��;k\��0M�:�a��|��P���	���'��֪4�쯻�ȟ�V����}^�u�B�?�!A�����΍����=.��K.�f�7��+�հ�!���{Ժ��8D�M��=E�4&�)R$��Զh�d��b�[&Bdצ�WG3��K~ �F?� �|D�2$�f���ܯ��c'$�[�ofQ[�z���A�P�dL�"]���B�o�Q@�t�4�l��RMjXو�\�Ε�R��61�hGM���,[�	�A���H�daŞ���]\6���۠��/z�k��4}�n��zQC'iR�{E���&��P�-M�t�������^{�G�U��J���}(/�=� wuG�%Y�������Nu�	dH���$������I}�53��z��ܒ�W�����(ș�F)U90$���%���ݠ�y�9���7��ŷAg N\L��ݥ�Œ��g ���ta��K��D�I_H��e��>�j�17��c�����9\��s����D2G��,q��p���C�ڵ~�i��z�	�W(�������-�}�u��ޫ�w���%��n�6L�-��(��H�AZf�����o��A�9�#�{y�l:�R{}xi,�������M��tt�PfvSW��MP�nԠ�T�+bؒ� ���1\��b:��̪�Ŋ�	��皞Y�;]��V�r�ح�V�e8�S�)j��ʶ�5��U�D�4ܐZ�՛XG��ĺ@,�-���ke���BҒ6 ���l����nkV���h�R8�PHRmA�tWV̐�5���6����M48��GiB����&˒Y����~���4-ځ,#65��i�h�58%�]���2C]��>�?�}��Q�2$o�#�r*碒��T���_rY�)���a�_1�l?��/�'v�"I_P&Dg=bc��k1���,�{�U�{o\��0N�?��g�IpFn�}�*�(��AD�2J�E�"��L����� �\;��]\1�\���~7���#��0ȑX��ݘU�1C��q��0�2J*��
��5�aOrO\���.��8��K����� ���$�Q�?	$oW�Uy���<����^[�=7r��[��u���"F��1���
��w�<�D['܄%].�`���%�a)�kQ�l�Z͠���3R��/�C�ۡ>1��3���Xݿm>�Ŝers�P��hY}EY#U���tL�7P@������zc׾)8mW+�&t�X<jY!��NӮc;a$Q��]S�E`����T������qI�nT�vn̸���g/�g0���_A�{
{�z�w��u�۵��&Fe6Mە^��ξ��?( A�u�: �#���bQ��z�����pOLݩhV��΁�"�H�|dH��oƩw��e A��0�J�|wj��2����v�k�=��ޔ+k��]�����sF�: �9�D�0L��H�"F�N�y�\����nq�Y���R�l��\ u�ч�ݤ'v�o�������)��gQN�u�U�ٰ��2Ф�B�[���T��)(%͸ �;���}��r�=��:"Dyz�,���g�n�����*�ժ����:P@���ݔ+�"`�"��{ڥ(�r��+��x�/�3�w{l��m.��|�rs�	�A�{P_�U�U̹�|�� �"� NdTA�F/��PϽ�߶�,/ұbgfm�t��j�KF�jǓW!���{�t+��)���_vVǜ��Y�w��,�������w�TVrKz�W=���>�8�mGk��˃�$�����S"��Y�cY�����z�C��;�[��.m�,���ka
��w��mf���`J_r�{vV��."���\�S�ۼ4�P�qm�2���e�uոt��������OK:C��ɒ�W�"�$���F�|�,O#���V�[�t�;����r�{�ڕBE��9������w��>��+�q���/k���b��!�����H͍�3��A{5M�/��ɤۉ�0.����Ve�V!S�ŵ��oP���G5V+��j�Op����m�Ui㴻�2�e�YK�V�����y�]ƛ򯅕Q��t�1��6f� M�8�:����`%�):�U������۵��U3�1P<��Up�T{ K鎘멚9Wd̓UUW)����v�1��h�tH��v�af�J�%�[��#���׽�tj�q�k��@�ޚ/FT;8*׽��mZu7���w�z�>�9��w/y\T�C�5K,R׵T����W�oZc)m����^U�tT��;ڶ��U�͋p��Z�S�Y�U�g�o	]k��M�����*�ѹ�{oEl�
s����Y1�(�Y�m�Yu����:���Y�y]d����W����)ԕ���x\�^�L�Ǚ�r�����+M]p�,�]f�w�rP:�����rACJ�p��Ƃ�o1+�zt� ���0�0Ԁ�[�Y~���]P��A���QE��f�n�f���Y���*ۙ�:pvkF�lM�Dmmf��R�c�+rH�@[Ggg5�-�DmD֋-�$2mkv2�C6�G(�n_�{m��y��9�ԎK1C�k,�丐����V�Lf�kfuh�]��3!8�2�[m���;6،�;Vnٽ��^n9�$��������f���e���:�n�2�cV6�k�Ăaڶ��!�e�s[�Dڛ:�f�5�m�h����co7�hI"������Dml��t��5�f�t�f�����Qpg;m9j�K4cdN�[Q����q���-k--mX�d��t�׶����R�a32n�X�Ӳ��kY����ִ۠��vջ[D�ե��+f����I3m���h�,K4���� N6i��o0�@�rFݒf3��:Z��z�<�m6m����M������� ��)�O\� �t�"����wi�$�K�:�@`�a���#�����nz��^�KB��0A���x�����3�{�P2/��0A�IB����+\���]�:={x^𻎵��!��PDv�_�L����}G2�Q]����df�0���\b��Z�҇5m�9���5�+Ð]Qi������H�$�)Ռ��o޳�d�J��<Z���|�Uӛc����(�d"`$�����kӻV����z0Ƕ�}U��J{�6�н����:��;�?�;w��{������g&�1FE�2,�]��{c�r^�.㥰�{;���?z0̑�H�H�����ݑ܃w0�"IB�uc<���z�n�d���� D^��]/�ng�ƹ��У�X47��P�9*��W\� ����@��^����rc��tu��[d*K]�xF�T��w� �<�J��2 � ��9��؈Nc��}9��e\��vv:ޙx�{8	�D� �A7[��$�o=Y�*�K��Ӹ%��-A+A�`���u�;Mt"��d1-�ʸ�
�#��̥ �&#{�+�"`�dLU]mU���8]�Ka�pX�3�v
רP �`�s�A0ȑ�A�?�������V!�_����O��9�ڗRd����?Z`~�u
Ew������E(�L��@������ AF9Q�Z�!�[�ڬ�i�ݙ�օ�0~7��]�"E���DȻ�mm���VA�(P>��􊝹o�h��z��E������?D�]���h���lk���;���Ռg{E&w�W=���|��-w�W3jm���\~�R�������追�F^״puf�����!�)�P�U٘���)j��2�^�K�[�w���3��z�y�b�<�u{� ���U��QX�f�+�#.e���.���3pV�[L��Р�lI]4eơ-!�afa���̲\١�6GSaF6�3YYk�����z�LJ�C�"ŘЗ�i��1�fe�WY�gQ�-���J�NJ��X�6R:㙜�i@�{��6��37��Gbf���9,Ga����Ύq0kB�F�$F��m*iYP+��Tіh�_g��í	�P�K�� `����a���ܫ(ƈPFѵ).J����o�2��"v�猪�{b�vf�Z�%[
�_g��x��Ț�#c�$�FD�>{�����x�H~9ԛ^�Ǿ����Ɣ�]A� � ��fH�Me�-����^�h�|���"F��F�Ax�2��7��NM���>�'d����������A�Ⱦ�1��~o��8����� ���;�)�ܵ��m{�/h^��	����oE����Y�dv0��y�"�	�?� l�(ȯT�o�%,X7��U$ٗ�}~[9S�!�����}�3$tD�4�U�����)�I��9��Ű�r dt�f�f����p��L�]�
pZ�������#u/���~����m��;'/���iߥ������
�L���D��"���U�x{��"�X�t�/�5@k<V˫����E�D�
�=7���^��>Yk����;Gr��msv=92��+���|o�n��=������{~�0�e��������9��E�O��bIB��0A�ȶ�m��h�C.�n{o��jB�`� ����F6.�.�o���w0��_1$�N�{N����m��;'/�k�p�M{]��^ޢc=���Ս��(c?��V	HB�Vh=�W��{���������r?���"F�"IB�>��������j6ơ�Q��b g:�rY�RåM�6�UI��ýt����ߌ�Ș"��l�Ѿ�l��]�:�:>�S�\/�h�0�o��#�#�&�h���4&��=�B�X�9Y����{�䯻�ޯ�H����Pm�<��~�/Sl�(��`�ۨ:ޡ9uq��������}��K�|�P,���:�Kt��u@��s�ǽ�ϲ;ےj�꧴s%NF�9e!�>���ܹ�V�i���]N��������B���oc��� �/��W�,����ņ��d�A����?n�-�o�=�;ݣ\q��|� �� C^+����q��h��g�g���DF�H�&H� ���n��/�c_x>�v2��=F���;:/O�2=���`?H���y���t�>��N4��9�9���J�P���\,\h�B3�S�LB��#���߾��/���$A��[-g����׷ԅ�d
]�W����#q��?��P��� Ș")Ԗ����\A2$~��쳝��q��|��P�܂;���jF.��bh ��@��H�"G���%�2N�1�Bi���z���vt^ �Z��(�Ș"IT)�J7� ��;�dc�{s{ۋ�������`�{3C���[K1Y� ��g+^�F)F�נ�4�l�r����Rh]��Of��a�h�2�F�cE�ۛ������ʛnYnj�*n�.R]��lb�2&&D�2JdK�M�Uo�A֘9S�rn���q�J�0O��܂;�����U}
8�_�o����$U2Z�L��%��!jGΤR`.��{M�kK�ΰxrQځf����k�6 �7�J�ӱ�O3V���sk�#�gp��Ufꀉ-�D"dI(P?da�u�{<��}����+S�=��vZ���z:��W���"7]���f��nq���l0v�|~�_1$�@ȾfE;BpDN�EWyYrn�gbq�J�}��wS#uD�1�m;���(�y������UX�29��5��I��x~>���ҽ�i��޳��x毙��I+�Ȁ� ��g':�[�Gx�b���m�λ\�e�:��׫�����IC�^�c��q�]T6�e����M�Snx��p���n�1��s�V��/�n:�3v��a{{E��ߩ�l�(��ǊS)��o���0JR�#lI�D�-��6��)��7U���BU�h���Y��)^�Z��%�L0�b�id�ٓX���iSfÁ"�t�5vU���V�h�2s���:��g)j[�G�7i�0����vXJ[ipj�ga�4A�����<fnaюiU�4&q�!F���u�af@54�hC��fg�ڨ��E���u% ���F|������kkeHe������R��C]e��a)-4iFT-�PU��K�b`��1FD� �"`����Z��v/G=(7���ګi4�]A��}��#K`�#�;�����y6$��(UU��1�o��}sv\��	�R��;��v��s���G,���T���d{҅� ��G�D�TY�I��㕌�����۸�n]�B�`�y��y�D�?��W�,"���gR�(#fР}�� șus]ﲽ.��^sZǾ7�%I#��ŋ��G�la�D�0L��F"Id��x���P��6��־�������Z�G�> �m�k�����"C(��u�Cp���!�K�+�\��\�h�-�X"�6R]]?o>J�|�`o��G��#,׽/{{j�g�:���w2�Րn�DH�_n��?� Ș!�[�;�����Ӿ�;n�Y�fq����U[�s������j�#`��f�{�*��gOhz����w��=J^���^�J�=����9��ݫ�����}���I6��4l0Er��_$@Ia}��>V}��]���,f�L�^)����� ��O��P�dL��0D��X�>E�r��C�$O����N�jvǛ�����>�L�s��VQ^��`z������A�?�2J�E=���x�=�_C3������V�\��w���}��:"D&k��Kvr��(�G[1c^^yp����at���INRZ57l!����*�F��~�A�a�D��#Uc:�Ζ����E�|y��KͶ�7�}��eX ����l�@q*����yׄ����j
��wj�8oc����M�yy��_��N.�J�P���r����a�"
;�������T��:C2fW��L'~�YJ{*��CB��W���ؔ�}�ܶR(��I�2߲����	��u|�Ρ�E��j��-yyWY�-�Knϧf�t��-��a�?���y�d�� � �l��NX=\����#����𹦳�;ʲ��l���=�G�Rvϑ���!�LA�&D��"da�$h�6.��%o+�w��o7�����t w�[��%9z>�r���/� \�5���̚1�R�3��2�6mU±s IU�-P�r`�6J�|��?�c/%��}[�b�	ͮ;�Tk��  �{�� ��H� #�2߸��Ϣ���ݯ�o0�𹦷�w���6vH� Z`�=Ҿ�3)/q��϶��r`��@�"D��#�F�C�݈V��y_�mO.�%��wP񼎁��E����2�6��kE�����P�90ADˡ3�%g�o��'k
���@r��FPB����]�M�J��)\^p�^�5Z�5_I�0���Y�z&n�����_{2�x'�.�����ӭ��i���^0:�+_��a�#��d��Fr&�ޕ��*����rޙ�+2���x��?�#�P�"`�d^�\A���g��>Y���ސ"9�ȥ��/X�mk�kM5����C#
��hQ�w���ϲ��F���H�a�_5�o�=�7�Τ&�1g��.D����=�Ma�G���(X�{�C�uMjQ��ծ/{\c~��:���%g�o����Xǎy>��$w�]D��K)���oG_@���}rJ�s.�;��W{��/5vl뚼 �d�B��0A2&�P��^~W��@�y ��9<��#�ߚ�=|5u�D�{C���`���z�h��#��(Ⱦ`Ș �(P2*�����g�9�5�X�ޛY���Z�ڂ���	� y�d��?�5�c�E�Qy��ouWb�m��.��aP�P�S{��6�E�s����'N^Ԫ|���t��a�*���k!¢݆IpEi����q�(,�(��"�w�>���d�6�,���]����yL���PםI�)ܮ� ���[�*�,c�|���+2����og�ۖ/;��G�+Jq��j���,报�)Բ�vA�Hͬy���᳸��ӡ�dɤ��͆�R��w�蹺�b�j6����ws�e5����x�ؤ
+��ѶL�����T۷]�͕k��L|��ZNe�R��^�$k�j�f����)s-��p��sVob�<�ן�U������={��-LmS���g=�|꺷�j���;���,�[�D�ۢ�����Yuj�7�p8y��Ҵb�r���:�g:�a�]Ek�/�ԯh1��W7�(�����U�r�h��M�7����j��4�$�(*���P�%��6�\�yWݨH��oQN^��8ڷ�y^��e�s\��X��|���r=ك[����j�L����us(VY��g��7��V\灤lTJ�Ngf��x�E(���}�b�*������qa�q�M��+���MQ3�$�^�H���{z��]ꔽ�B"�������#�������x�p��2���J��zxVh��J^�ޥzj㮎�(m�;4�ʖ�p����ڛQ>W�D̷a�ދ���'8�f��9��W,n.�r��Eb�z�l��Ak�e$T�7��߳%�,I-����Q���h���6[Ƣ��|0d�-h�mJ�͍A�$.�>�tm�m����fBY�Kl��s��R@j��fB��H��c7;}��ۊ��"r'���$C��M�f� 9:5��Xٖ'H���'K7If�f���GGD&�{v�q/kr����nёi���s�(��@��8��;���S6۔H���9'8̉!(��� �39.^zs��Om�Rqӑȉ+n��f� �9I9�N�PB�t��������Й�;5�����vW�i8���6�'������K� $dR6�t .֜�gn#��B'�)C�E�mBC4N@��t ػ9�A�G'��rB;�)ā�����
(�����u�3՟�4B]�J�b)s2��_������h����U(j���Yn(-FmS$#]�m	Fn9�Cjj�ЪV�u3a��L[a2�L�X4e��#�a�!%йP��40�.N%GVѷ)�<���ҙCV�cI���-e��`F��V4a6�;�WQ���+[-
vm�`���ut����B��i.���Jm��X�H6m4����hiVɒ�E�u��Ż��c�0��h�W��m�®��b��t�]SGWb�J%����BĮ���ڲ��%2Vı���*RƷ^س;�N��
R.XJB�f҅GAp�hˁ�b��Ac:�tպhfcD�����6u\˵�Ђ���Y��M�fYD������7�a��eD�E�E�5�tȌW1ɴ6-n�.�@���Yt���T#�tM�C�v��+cC62�l�\*]p�{W�a-o�:��i����l	�bkM:�c�+�����ͪ�i�̚��aد.�ܒ4�j:��Vm��@����G*P��3á-�-�f�k�`�L1B]s� ���u&�M/7�"�3P�0����]m�l�E4�s�,	u ����m�EY]E6)e�:ΰ\]M�$�է$ņFV�U�:��q��̂^4�P�����3�Չ�#-�v{=pB�X�\�bL�I�%�Hjh�i��]�� Z�
	1+��˥���n@��Kc�cP�4v�8Msڥ���U���p@0ݫV��И���i�mP�:l���vh�-��I��c`��M3[F�h��"<D�4]2���[��뵩*�n�dX��.�ض��Pڨ�v�ն����i�D�K�u��]`n���V��7L��˴a
E[0e���RU�<g�y4aNr��Saʉ����mjlܕ�3�Bi�6jCF�M��n42��b�p�9����9\ ���6Օ�i�]\�ff�e��!s���c;lKM�u�{�ե� ٠�
C8��`��t����1���]���횮c����R��R�h��\�hXG�n.c@tɮ�	D!YQM3kؖm]�wZ`�2��������4e�4n�6f�B�կYt+�,fM�m��nVi�Kqv�����f����c<h�JjU�B��61�uYHV��i��M��B7D.�)��Q�g��o�~�%(Fa���њ�:�E�%� %�� ������u@URI"*~�0A��7�	-�d�(UX��]&w���{��WV%_��m�XA��{��A�2$�@��;ٷ-��|=���`��D��-.�^෯2'�}z�NA|F��w�}�yd��V�_e]
��A � �%
�ș�E�ú�M�գ�^c̗���ٔ)��y�$xA�F�H����d�A�	-�d�(UX΅{�}x�m^�yu��z��{��ꪢ�x?���㼘I(W� �2?���
����{�%ݷ\�/p]/r/ECw�@�����#�$�;�!zV�(U���U0��[]4,É�]�ʍ�Ћ]�@(�q��vS3_=�_q�'��b�2'�UvMy�y��̡K��3'��Ԯ]Gy}�t20���?#�4�c��<j%��K��ڏ�*�(fҼ�w�wM⨣���7.#��u��n�Ƹ��%-��T��bʽ��c2�`���⍱)v�v�������Pop��m{O\�'=��5����vic��f:�#�P�� �"D�: ���`����ʏ���7#�T3y���A�����%
2&Er���hR
�IݒOW���A��F����<��u=Ƿ(���r��u)OJ�zh@�tA0ȑ��H�~����8�^�	���P��=Ӷ���ⓞ����y?�=҅"d"7�"�=͏�B�1h�@�;[il3D��R-&q5خ��qD�t	
�PLGs���A0̑� �#e{<v粼����66y��u�2�1��xg�����IB��Ⱦ`Ș!XgG�5&��!�Ek��_0v&c��&�{o|�mL��W��2y�d����d���w�<�$a�F��"IC���ז����/��K���D��初�}�)
�u���ު��4�m�]_����g:����+�Oi�pm�C0N�B-鵜:�9��k��(P2& Ș"I_PV�X��u:�*�f��7�|�P_[���r��$7x A���_j��*���#61_�Ș �(W�E�;ϥ�Z����o��r�3����ܠ����Gu}������<b�}EU��UD�4�"��X�*�^��.��`���-�0`��G:�]�
����_u�dڀ������0�������2s�_F�7y�mZ����(��șJ��@�y�m��h�;���#߽�K�~���lI��7��#���>�ohU7�W˺��_`2/��a���ӿp��*`�&����m��Ak�X���C������3��I���^�W�V��Ә`���P�V3��Wj����׾ ��Lw[�:�W-��L��|�T�������ӕ[���:������:E��~�U��:�j�K)�^��ؕ�jdJ�4�ZGMf�yj�.����?����%
��$wS0{�q���ߝ��wsG������x��tA�0ȑ�����g*�'�I|l���BM��
�Q�M):a!y�:Qx�u2�lG�A0�}=�z���vJ�	��3=&��o}NeL��
�GU�N�}�x�NtA0�0�2G@�:�:��:�ӓ�A|GJ�z!'�yä�pS�wb�W���L���,���A|������A���d��H��l^#�7s�'���W=:>�bO|��:��?����"IB�2&�sεd;��"`���V3=&U�o}N�L�>`����������������;#���	=�X��z�j�SOO�6%W�IpS�wb�W�Ԉ;5�ݤA Ȏ!�}����=핯S۽k��-8�v�u�k ٹ���	�Y�X�E�x�3 �v{���v��D�հ��Y��*�`���{�ϫWQ�"���t��ƣ���۩��Y�t	P��uf��]��Q�+�s�isDݦ&�����òC]��.LF�î�R`n4�u�"��v!m���6����q6�e�b��f��b�r�+��h�4���[�n����)��e�s���E؎r5��M�cq�41�˦f�m�,lh���a��f	.�8؅�.��Ǭg����_�!U�v��P����3�����[���Zh���������|'�#�wu|��	vv�|����E�Ll��Q�f�+���QC;()>����m1��T����<sR���y2�rb+�&?f���ʝ�hq�AD��C9[eg{�:l23���xD�0D��D��ʻ�Wǵ9␗��7�����mx�}i�A�_H���2$��K�Y���sv��� f���F�	K�ӯ�u��-��C��&A��_�y
���}���dL�d_9%
E�<b�z�š`㜝�w�f����}�7Lx� �0�2G_dc$K�e���Z�i���s0�s4�#G	3+Me�to5��Y���u��a�Z$V��[���c��H� ���Ow=7�����m}Z층�m��~�}}B��3��D��2 �^T<*av� ��xq�̭ŀ���#`3ݗ[�~�����r��v�T����5�ڣ{`�����?Z�*ݬ�^6�Y�y��]q]��(%3�N�E�n��Զ�o ~7q0A�����jߛ��ք2�A�L�#�0?���1�Uq��6Xu�ؽ�{��K�a:�Nr�#���D�+l�U����ۚ�#b��(UV��w-7�p��v�A5�����8��<�*��r`�DȒU}"���>�K�2�y��� ���:������m��n�d�"F�I(?!��_h�e;�|�up:�B�lS8�ȑ���Y��m6u)l5LY�f���k�޵> �n&A�W�,"q^�1{v��u%���0B
�{M��{�Bc�tD�2$l$X��EWu�D���5���f��ލ\��^�}���D�}�^��U����h�zRz��'y� ̑�H�L�^���מʡW"���:O8�n���9Ŏ�F_R�UR�Y��\�4o���x�s�F��N�11c_h���j�]�#(��1�w�������/����d�(ȟ�d���[����;�o���}�X ȟ�^�a����K�a:�rPD[;Nc��a].�`��|���la��:��$a�'{_�ˋ�}��P��:1w�W2�W�\%�}$B�� &E�V٪#���]���� �E����]X[SZ�c�����-&�5Ǝ��3����&�Tn��X����Ld�>��c;�(���u�.�w�&�Lf�C_���y)> ��r�Ē� ���C��mU����i煃|�frxzl���گT������@�?���X��L��������da�#$�=��ː1^W)���xI����NWk��k���+�dL���D��
4�`C���:>B��?��:���0���_��,�;]	<�3���Q�9���R��To���YQE��aN���1^�,�j��嵪���}
Y>��-UW�)����7/1��Fb���dL~D�I_H�L�ڥ/���=4�٧ۻ���>�	ׅ� ��a�$T�/��_<}���~��vbC�.%�9%A��n3Ɣ�v�a6S�Z�K��ua�W���My��A�PDn��#wX7�T�2�];�[*�\�u��J��=V/y�� A��#�Dkps{ڗz]�7] A�%�c;_�u^-�6bcs���D�a�$���W�n� �ߨP9��AJ���Eu��הS�=3Gff'�5Lb�C��A|Aۺ�@��D��/u�OH]p�ǿF����n����T�R����Y�� ���F�GBl���,�;���x�%W� � �$I����꫈6�W�7�^Ư�g�΄��g:��;�	�����>��e����ǡ,UWk<�=�+�����?n"�v�{�޷s��G!.�e�R�iG�s%�l���x���+l��h&�HmUJ`��YZ��
G86��Yy�a*\®��+�n��lF;]m��@M+�2�u�픅@�3�֫1�� �Tuuc��J[�����508#��cZ����[�hj��>$�;Mm`�
�Vin	hmuĳb���7�cF�� nհaKr�n�M[2�w`k��r�;�[���̙�Z*�6�ֺ���=P���(�������4Pd&�L�;bfճgH�`Z�Ma�ˢ`)�I{����i��	��뙣�7U{j>�ר__�	�j�*��d{Pfz: �[�$L���pZ�b%�ۜ���;�cΩW~�ͫ���z�]#�v��bk»I{�|o�#&РA����_Hù��o���yu^�8t��M��s��#������6J��E�Ue�v����E@����?7z{&A웪��m����L�����z��?�с"���\�Ҩo���}�+��gQ�~�ͬ��{���C���E_����y��щI��!�B������RҢ�Ѥ���Tz���>���[�@�bFP�[~#�R�A���܁�7'>���yi� D�|d�+�"ddL�F�����7Y��w�'J�b�4��Ϊ�:j���=;$����Q}4P����Vz�k$�m^aׂEJ�t��'�V	6��<�+K*���(��n�Aؘ7p�L��3U{n>�	ר9�B�2G�^v�f�����"���o:#���$�$J��j�.v�cݼ����-�.�����H�; �dL�%}B�wf{�!?_0�t_=�9]���~�x��&����}q}W������ۊ���#7�P2&&E�%}"4�d���f0�7ɞ�;� �L�^ۏ��u��A��0�2G�H�e_���AS9����k�C�4���WS��l����0�moSDr��
��5�n�>��ߞ{t�0D�?��Pw��vo�<����u��<�X�f,l�.���K�2&D����A�1���-8�뜠7�B<�7�[�x��3cbo���`�' ����aܢy�� 7���X'�2�W�, �}�� �%��^�g9�WMՖ�b���0%�TG���o�V��%�Y��\u{Xt2�6�c2�R���k�R�uo���4� ���
fH�	:0&�X��v��Yʣ:���7.�%�wU�f��"���S u�m�E����^ԫݔ�Kᕙ0��ıԩ��.�p�O�b�p�A����Vk�,V1�5q�;�T��eh��w��&��dy�t�q�ݜ��x��9�����Cx���.��$]�ϫ�ψ[�-�oLJ�Iѫv��v�5��u�i<�ڤD��IK����F�Y9�y�T���n��}}b�oH������g(�LWrj��9���m;�I���C���܀��߯��u\z��|�ʃ���ڽΟ>ڻB0��o��Jiur��;P���W���̓rGr�fLܯA(z͌�D]=���T�O(7f-RX��X�7~��*����+S��(̼��<6�V�,]�#ת��+�|5�wW27Ij�����tE�*�}�2���G��1!0M�u����T��՗��ٵt&kvi�c�����n^'1FS����d���2�J�%V$]!w�:\Ô##�^�X�r�=�Y��|���O6^�wO9��p�>i:��f��آ�7+k��eHl��Q��f��7e�N�U��ہ�C��5;N�9��<ej�����>[{��ݾ�݊�h5|�t��e��nQU��ڹJ��\;Z5l���Hn�]�h�G/�zZ��t_fd%V�oI��Kýf�N>���L䥎g]V�V�0h;�Tm?� ۷H脎!q�s�ݹ9��D�܎]'$I$uC�A�Nt���%�@�*8�8�'%���H$A�η;�[a"$��0D�����).$.+�/k@HDF�p'$������8�l��:#�Vb]9�Gs���yv��qC��C�8���gn����Нyd.A���۲9pGI	QBqI"���AH���8rw���:9(���m'r�t�����ݬ�GS��a9��8''+78��8q	H�#۲8Nqy�%"!ȑΈBqG@�"JN�����NH�8�$^���/-��r�s�Y��e�$$twG8���YYrQYh8����	�l�s��N/j��� <��mVOn�,��������Bt�u�8�P �$�������wd��5Wm��a:�@3�`�=�3$T�0D������>M����G��d�*�ٮz�f�sɹ�C.��=H�]��*��{������'��D �fH���\��Ǝh,{�7�+�{[��;��׫�9"��������1��h%MS�M6��F(ȫ�m#m�]4M-\uu�aR)a�go=�~�ؾ{�P����dB�N��=�5W����Жh�]���X<���?K_\���#|D��d������7\���W���a�Ků�^p�7/5C.��\�n�*˾��&��u�6<_R#���{�#�H��#�	=Ҹymؼ�ّ�;�wU�0M�tA�/��P�6�#6ǐ����+$�x�Ka��@�dB�{�f�l���Jv�U^�r �euA�^��0��B������*�dm���E4�A]�1��z.�m�[+2�R{�7h?K�	^n�nb�����Z۪��T�PL�g�qp: $���� ������T`���N�;��ۛ�������z����;��L���W�~ś�챈�5�%��DT���j��4t6��%5�kZ�̐�B�m4oj�1�o��=��#����WI�O_-��d���bi�д\oo��"�}rJdL�dL��8i��q��,�r�n��nA�{Mwm�u��D;���d�K���x&�_6=�?�H�"F�2Jd�WeF�����Od<��Pͮ=HGla���L��D���]c��ê?R���xA�F����:��9�guP�_U���S�g���z�zt���a�~�J��2'�IB�2+iu���ۼQ�x��ET2v׺�w�2�arg�y��A���d����a�{��a�;�j�6�s�v�](�3s���b��j�>F�>W~��w4J�{ܰ�]nS;�K��=O�
������`I��z�I�eL��g֦�K�V�j�&e,�f�l�MY�Q�k�Fa�phZ(�4�ЃT�hk7,r���)��w$�cJ��)Z��3KfF�
2��ڰ9��3vum;&)T6�cm/\Z�A�Ҥ�MT���t�a��L2���:e��u���n�0��-�<\Tx+�,�(h�飗Z�.��:��o��c�3")�Ḷ��b]e&�����ܤ)&�����P�&+���pAL��CCk.��h���@��"�ƴ<o��D0�2J���]a���j�mq����l�b�׬a�� �"�I�P&D#�ey�^�`�b`�܇)������vF��@���� ��"7p�ڝ�yf)�Nϟ��
9��Ord%
2/�2'���1]��LM��y{���w�2�arg�y��hp �s�H�"#?u��r��uAO�{��#9/�u��]�:>�&m����x�e�����C���ÞO������D���?���ߏ�W'f�6o�@z�5��;#bg|�ש�@�a�#������{3�q��<�%��K���#����B.�KB)a�ٹ�`�6�Q-֒I�/	Ș �+�@2!y��������<+Ͼc.p����B��iv0��GD`#0L���r=asG.�wޥ���pS�=>�ÿrWRܚfg��m�v�j���ܘ�jc75������'-���6�;�oY�lo�k�jo�r�W�5yv{Nt}�L��K��}�z�zs��噛y¯���}��@��?�#�$P1JG9�����1��}�����'uP����G��H���%
D�"������\6����W��O�2&�����3U{Ogm�vǾ3��4��K܆���	�d��H�I�qbW�p��Z����s��2g�3}�mw��c����c��ӊ �ٮ�����fi����!���V.cXD�ݝ)��jFR6�?�	�|�'�NA���A0�T�����롑.{̠�V>n�#1Gs$�FD� v�w�}�G������% }}x%����^���a]���2�#�*��7d!���ц	ݏ�0�"F�2J���X��i�U����4w\��������p���T���y%ڙ�)�����2��Z�lu�F۹QL:0d�T]�=¢w�+"ǥ��p��S=���d^ �\���(ș"H�n�ӻ�i甅~�N瀉~�$���U{�$�����0G�V��K�Z�q��G{�(ȟ���	%
2%��w�W�K�`E�@�z;=x�a���@�9D���1^g��۝�HC��XI&��Sa2�M�Ao�b����,��U��ld��m�2���Ϟ{�'��`D��d�֎�w޽��rl�2/ ٞ��nQ}倍�b��2�DȒW�;�">/=����ƃw��dA}���W3�Vt9'����ש�r�7N��{M����?����ܟ�%
D��v��U��n��3��^'|$��W~������fH��$!��S�v?	@����a,��s;��/۹��v���":Z�Ǽ��uOQ�}M�k��ɕ��Vu��7��¶���`"o�=5���س8Jsk8ԉ�_t޲��\��w�Y�L@2'�F("�����n{�S��z�c�N�)\��Y��b��_z�?��A7R�wPk�˖�M��*�PT�����Fd{JM)�+��K�i\�����F]s�����q|���(Ș?H�_^���ͪ�	3<���y�pf���/��3+��VAF"F��:z���[�4����0�#=(UT��$��s�6_�����wj!�>�>���XN�vr��bF2GD#���D<����bN��5=�{��D=���"F�F(Ș#*^�炳� �e
=ɂ	ݤܼ�/���I�a{�'es9/'o�a펁�2$l��� �@�ٽy��1��~��%63'=�ߤ�|v/A�L���P���	�0���5!u6������0;��z�^rIFE���m�ː>YX��o^^�C.1gm�����a|��-n�}�|%�Ƒ�Ƹ�+5-64�)�uX�B�j�t"3B�SJ�vq�(�v�Da�c��D�õ!�RY�8`�q.h��*��K��F�\֮�\P�kT��jM�Da��l�m��-�pgWsۘK(؋�Gg�k��u��,�MxM�#�c�kjCLT�p�II��p�)�]����i�vT�]���[�&���@�Q�����翿>���"]�J��J�h �m��1��X�pݝ��4V:��A��?v����g��H��0�&�&�7Ҕ���2!��nI�=�L�|V�3��w�0���IB���2&]�@�wޙ�yE+���O�?�nh��������7��}9 �`�h�����}L1���a�����F"F�I@�/4��8zN�7ss\9��\��0wi�L$�C�FpzLG�A��̞tF��<���JS�d����0A�������;�*�������AE�JdM��U����T���+|oٻ�~�hw~�L�y�d��F��i��gd��}F�S ��n�AR���jD0��⍌%�[�h%J�b�k�u��[�o���� ߼����H�rJ�V���\�uss\7��MTЅ��Es�\�>���2$�("���m	=f��w��Kk&�!�H�U��[�bC�tNnSiz��]��5w^z>�s��o`���]fF�v醯.��5w+���Yg����v� ���y77})N�mu��0A����a�$¶P�>U!?[ݡG�0~�L�$�(�"D���2���uz^f{�I��{�'eA�0d��20ȑ+>%�k��o> ��a�����$�U��!��}9�t�|r/A�L+�o��>~�g�؟����"I@P&D ̑����qs�X�+�	������}��T�	��6x0~;q����0�2J�e<�KHwSI!Ȥ�\�0m�YezƐqPB[�#Ϊę�u�/)5�[�JH��` ��� ���+�st�w��ۿ�4]_������:WR9؀�g�����H�H��H�qoK<�����}��M��!�޹9�t�|r/|~�O��u
D	�Ns|�q�߶� ������2��#���X2����Ɋ��9B��Ǔ���U��j�D+�CYyi�-����R^֚�}�.�;����'T��:`��W)����Wwe�)s6���͡�=����"$_I�/�l��Ij��3(P2&A�Ȱ��rە��ݿ�4][r��OĚ�S6Ŝ�P������#M�>�����}7X�ʡ��v����w���x��_?�:�|dLA�{�׾���zF1}�mWl����8��a���3*���V�6��S2����ƙ��7�����>��I�!:�H|�g�ʽ�6���:���_%&��a�Gy��JdLA�}At��A�B����bc�h���ͼ���&�w��A���3$y��e��غ�#q�L�P���"F��()y�s��^��F����[�6_�����G�1@Ⱦ`ȟ�I*��{��s�e�{�}�����A0ǥ����L��Cu�l����Έ_}s���y�6�R���N�V�0��kj���Pl�K��"�,G�V��D��{ML�ۥ�NC*�$%��{�خ�MYBZRI+��/8VJ5�È}_!۬0v'� �$�_C��hX~��X7��:�U`�f�m�t���g ��3�: ��C�B�uN�� ���� ��"�[h�fR�;(Ia]����^[��u�;���}� �2 ��K����>��&��Gy&K㜼~�Ћ���+�u
 �LA�0D��}"��K�Q	���|rj`���޼�ԧ�n�]9C3�@��� �܂#t�;�,���+��d�'��I(W�D��(޿L��w�1��L�;$�����@9���� ��H��ێe��e^������|F�sDŽ$���]�����.'����L���J�L�$a�$g靖~oʘ_-{c؅����83��YOhfP�� A�Fb_�� �$����%�(B�`$�	/�$ Ih��%� I_�	!K��I_���%��$�	/�H@���B��H@��	!KHB��	!K�$ I@$�	/���%���$��B��$ IqH@����e5�w]��G�Ř ?�s2}p!���           @             P          � �UP	*T�  �@
(��I@TD�H	���%R(��)E�А!
����UB�"��*E	R�AE)JJ��H���J�UH�B�T 
RE$%)*��  }�%
%EH���H@��l���J������*��sz�;���CN��W����:�ޠ����罀�"P��� �� k�˺V�W�)^�U)�ǐc -�=Q�y�WOz�J�t3T��w"@Y��Ei� <E@�|  =ꢪ(�%B�U")UH�ϧ�PQɡ���
<�O=��Oa����PR��*�΀J��A@	,� � )����X@


Gy�TNS�w����{���1�
��   `��`�.�tzi/z�g����a@��u@S���ۍ�*��:w{ט4�������t�x�t4��T���W�  �H�P�DUJ�UA���ҁ�� ����޷Jٽ�t.9R�Сޱ�S�ް��S�P
�y�үx$t){�9
gN��U |   ��/I3����9�@s�� rT{
���r ��� /{���u �N�z��B�PQJ�   >��$����*��UI���{��@�� :;� uwH�9���{ N�0 �w� �&�JFz wwW�B۽`t���  ��0�����窪K�=�����u@wg�=4�� �y�\ -c��u� ��� �*�EH�   ���J�T)U(���' 2<�n����kP]�Tl  d�� �:����� ;�:E"
�  @9 4�EK O���2@=��8�E�u����A� � x����I�� )�L��(h#@��T�)P  "{R�Jj���J��(�a�j"m�" ��������_�c�s3�������Ǽ4f��Dܳc׈�T���>�B�ӗ����$�		�H@��B���	D� ����[������(w?�V��p�K�Z(�G��yI*t�Yy�j�+��p�T�9���.<�PTz-E�>��P�t�U��e��]C�k�E��V�O�a�{F�Im���>(v��aM%uM� �f��S5�%.>�gg=��[?g[�rft�U��,����9o#�l8s�v�d[�VL@ݫf!�RV|����Ӹ���Y޹N��"ֻO�aӷ����iT�W]X��I�	�Ұ�И�4m;&�6�#�c�fl��n�9wv�>Qئ@v���շ�O�LW��M���^������OVK,�?�yj9�1�{�kWwE؃	t0sއ��s����b�L�{�n���w��t�;�ǡ86��͜t�ql6���ӳ�$��ԠѶ�2��KU�u�u��{y��|ur���R�����^�|m]gG���K������gi��V�Z�C׻�u(�����M��i��cyD$d׋���V����4<І��-��;����7s�w���W�y?����Z{J�E��z��,gIa�����F!*}��Գ��8Y/��y�m���bQ�1�8�x���6nTA+�@�m1��>�|(�5�e�\��qq��a�!��[{&��Z�v�����a���2���=3X{�'1�]E�B���C�5,�=����$�oX,[0�ss���wh�w�4݇p<դ�B��Z*��'8_�{�x�Ǹ�Z+Sh���Y�9r4AE	vgt��'ml���T)l.Y���i����-;z䗃c�͔s����2��n����"a+�q1w��j��A�@xp��s\dc�,k�s�`*W(֣�ot{qS�wf��{�s�^Ԡ|�ym���{�=K�6t|n����\��ԢY;�8�z\��$oKpV�[�8U���*��c�����u{dY���@�	*�Z�����=�D�.�xj��uoa1�tI���v㔷uŸ�h����/BП"��f|�.�Gˮ�,Lr5�7rz-
yF:8�V��{v� ����\��9�ܖ�H���z�خ��~����b֟�8����k�wx�nvܹ��t��F����
.����}��a㽻�l/�\;w����j��;ۼ����b�R�0��:c"ݣ��؞@����`���l�,��Lm�U �
���/�3�	��h�Pz�sJݱ�s��#�!n��E�Kۛ{YK-�@���w�qԆ�f�s8��n��@B���KC�����׃�T���T�����Kr�L6J�*�{�)��8;���t�y1Q�ҵ���Vճp��b��ٍ�j�:�j�Є��vC���L�ǌdGo�P/��9�#���N���C}�r��n�z�W\�{����Qc�� ��3{.m��uu�a���TQwi���A��wD��{�m=]������[���:�0�[OKƎ�E���u2{,g�-\����<^>��z�&�z$tcނ�]�h��d�Sۋ^"{y\���w���\c�N����;1�-��ىj.�t!���t8ñ�y'P�q�`�Y��:��[��j���� ѷ"y}O-<d���e��-f�F�7]<�yoJ!r�	��awj{�Rp����v��v�!A�to'�p0����/<����"��x,��3��*..��s^N��p-U$6��X��([Mhn(fX��:3�_wj���S��S��=�T�(g0�9!�hYҰ8�[�q�)����cgw�ۻ�'aT@ߪ�����Ӥ�P�TO5L!ˁm�X��wY��94ٶIq�u���fN�ٰͩ�\����݇Z��7��5vu�M�v����&i��L����ʧI�BN:��q����:��aQn����v��������sNZAZĻy����uޱ�;��ݼ��fª�.��ը&��t���xi�xl�}!�1S�9�p�ڥ�9N�渀���rp�X0��t�H�mo:Gt�k3Fq��!?��%xӼ��郏uR|(���[=hJov:&riqd<ZP}��{U��{`�����3�ɉ�P�j[������ �V��hI��L\�gr�{��bir���ajU;�j���d+A�r]�`��64���ͼ���p�䮻�=ǳ��{7�3f2��)�ʧUQპN�e\��cx���x�$oKy$�DG�9�G�.�d��!��%=
��>ۺ�7E�hF�{ʠ�!U������N��k��9�b�����-iZ�.A2k'o,�@z���H��A�|��&欼��1Q������7m�ndf����;�t��ܡ���f�&F��F@�/C6)�	�U�(�����PP��<��� n���Ŷ{,��G]��:;�b)]���Y5��ǆ���Nv虤��4���.U���M���_��pv!�^:ݏ��{��4DŨ�B��AɽH���&���wh�7�9⩹��q�%�RZNv	zᣪo7M�t/���nݺN�4p2����G)�y˹��l7:+;aÇ���OMzy��҉���6BJ�E^���_rp�	I�.H0E���h�FxO��6���B������Ghԓ+�P�%���N��:i�؇j���j�°sC�u�L10^��� ��d�m{,�ږ��� �M�ۃP���0�h�Y����sz�hFZH]�d�L!B�R�z�ʃ��n�9oC�X�����4���I0���ڎu�
)��4bG�M��������gqFx���/n�0�ڲ:x@�8������ v@-�̝p#����C}���P�d�@ڸ��q�;v|Kvs;�y� �g(���DX� ���%���^���w��Á��Ѩ���{B����)�݈��F-pw�:�#L�)�������i���Ӎ[�� z��L��
rF�3��2N��7�N�UN��"!7�Vk�8,Y;�yn���I����[�)Qԫț��x�x=չ��+�eC��6��'c�6~L�0�z���)<���.�곈���+��?֐-�<]�����`hE��(۸�{�����zy��z�ᗶ$q�ܛ���j�]z5Q�7E}pt���a��H�Tl�=\߇�ymݐ��"jÓX�7�r��0mh�`��K�G�Q��O��ή���olv���[��.��{z2��پ	z��wm�}ܲ�a����9��X�l�1q���es���t�Mw6���qjx�*֋�c=p�w�n܉�4wm�"Ea'���_���:��`���1���B�K��r볅�RO�;m�CsO�Z��q����(�
�G�b�7�!7�^=&��	X�E1��&q'�[��ݿ�:Br�6�(�9��KT�#-Y��K�q�unQ�~]3�J�N��rѲ���f�����ɝ'I	IK�\ A��Q���@�k���a@�ۋD��lW�Y1MSI��>K�w$#ׇ ��`�`���N�.�$@V�kK�9�c�wv��N�&��q�O�M�Ky�»MW��`�V����哏$�ׁT_�=�NW������+�,���;�0�t+��Y1�2w5��JB��ɬ*kt�r�x�C���s��=+�<�Wb\"���0�ޣ|ln��W��μ1`���m�)/!�w.��A�ȯY�x�t�L�3��U��(RC�%�E���Y���K�>E�Εz'�Ncs{,tnc����խH[���$��);x�u���YC^������|	��W��p)�X��ݜ&v�'J�x1��k;8���qW�N��5�Y�7�,YxƇ��ͧ�M���own�<��wJ���q�G��A��X4���E�v�
�0F sA]��z�0�J��r��$�xև��"��A������Aaï[إ�8��dM4-Y\��;�� ����w�u��9q���ðmIvl���j��
�^Q��,{S��n�Z�N�X9�NF����w^���$f^��=�U��5=���r$�mZ�s��H�iu��>���9�*�R�6�� ����o�@��7��sxe��s�� <]�+L��
nT�ľ%�{���;D��-���̮�m;1gs[��;��R�R9����8��E?NG����R�P���Zn��j��Y���v!0�=��$3�h�mǠS�f�CѼ��S��(��OvqZ��c�h���4e��4�����9�07Ce�"�3t��!�H,�:���F���@��#�����4j=Sr�neˉ�݋V)���3��@����-]����'f��P�	�4�+�\�J� �ö+�ʵ1��CXC��E4෴�u%K����a�t��8!����@���]���������4N՛�!dOQ�zߚ����扣�vg${�\�����`Ԩ�y��Fىq8��_;�:u�W���0��9k���A�ѻ����.ލVi�>wKގ�ׂ���l\�����#�9���Ö��'������/� %��:����r�8:bb�Ւ����HEIJ���w��S{�2h�Ǯ�8j�vr�@��)�.��� GWfζI���3����֠;�C�^���0�2M�")j}Ӏ9�b�7{��i��y�g��|s��3D�tt�S
���4S�H�yizhɴ��.�Nb�˒�����V=e��4�%V/�z�<`d�Yu�Φ\��Mۦ$U��Т�H�V�"F�F4'k�A,Uu��t|ws�	+�Y���>���V�p�of�б�ۇ["�r�u��;���]���rn���{�=��u.1��)&*�w-u���'�i쫷����1 ��D�5a��$�l����Hv׽�)I��{6�ύ����կ��[s�$�[݅J�lagIyF�8У%Ȫ�,�l�h�tn�Ä�U�sh�9']'��i����I�6НÍ��[�
J7 �ʣkZ���Aϗr��	i�;u�0�\����up������Ǘ��Bcܺ��s��NvŅ��X{�=$.jl>)���&^�G�,a�4E�$[3U˷�%Ɯ�p�w1oL`kN�A�ɝ�K��SDd��A���h���z��-,ٔR�aR>ގ�4ɑ��rHv�#���x� >,k]���Oiou<�1ŉv�H/�a��7@�o��HtQ���{������u:s���V�!�K�Kc��O�m#���侲���j��4��wn⁪�{-�uRun��6� ,E��L|D�L�|��
�s����׻pD*�Cz�	+��n\�i�ƝQ�zn�A��-���5�����-��3^V�v����ǥb8�j[� m{��8����{�OR7�qg7�������j��u ���I:����˸d=�]���.�@�YFN�dxY�
x �����ܔ����B�"�ǫ�^/��3��=�zc>����^�,}�I���=�X�/<�bXB����5n����ycȱ�;`Ff���,�P�w-tn�*-��iY#j\�u�w��'c�IMju{���; �4D��ݗB��
��L�.�㗫JV��cc����>h���A:�OS�wPb���ރ7b��r��B�n���B9�nj�0�7j�@W�J��8YҰ�>zp7gM�|V'��qU��������-��3V4q
�2nǣ�٧\����־Yz柏u��V��[���;;S�pu}{�}�M�苐��M8�3z%0'X�mʻ�<-ŽԄHa�wwm!"�����=��.�۔ �E7w:� �;��Whck��W� ���¦]O=���<@��C��rJ����gl=��Op�q����|��9:S�Ǯ�ԄH����u@ ����:A'�A��p�+���<X�5���nȲ�{e��7���i�+��D�lD�C4��R>ɣd��`�P�k(��������ށ5'�tc��q���'�uuf��!� �N�3U�:f��5��sd5K���4�Z�۶Y�*1 ֎���.�n�A2�r�W(p!�����\�2��"�����&����_r��r�{��^%_[);�������ӗ7�9!`[� �V�֦<hN2�-.�ԁ��K[{���^���ʵ�x_�7q;��L��Y�4�x���p��U橔��u�
�u�͌-�3F�ܰu�M�"\ȳk	�R^w�DC��4��jխ��}1�&S��He��r!��:�k��0`�{����y��r&.qa���s��T�.N����{�_����Bݝ���8nvlƴ �,�zӒ�}[�ѷS�P6U��O?p��Ѽ��P�+q^Ͷm�������i�N�[Y�":��aq嗜�i��w���M	��M2S�e�Z��;��킍f��V
���3�8��q?�v-é���j2�:zfwQ���n���{[Ȃ��y #�v�F��¦���p�^��tyڣ46�#� P�������7�.��	����IVmR��fM\���5�1��#ri ���b��8�U.�Tn׻r�x1��t��e��D̮#��{�]���Y4�������QS;{W0Z�D��nAw��w�q(+걣��H99`�*�u�9WFYn�{��ۀw�/���$H)	@I H((@P�E� 
@�(
BXHB,�IAH���	 ��HP	@�I ���$�B
H@P��$�@�R�HE�AH�A@XH" �����
 � E	d��� ,��!�Y���뮢���AI$�������I((@�)	 X�,�H)$ �Bd���Ad�Ad	$ �H��,$X
@� ,����,��(@�$�  ) ��HE� d��A@�) �$���X
 H��d"�B(�	"����EI��� ���I	{����~�2w��̉�A�͸�([R33��z�W�d�*7{�3��� $�e�O��W�^Վ{܎�V�=|{��WX.��-�FYwImd�ɢu�Z�__Bx����87���i,��B����ٳ;�(#tٸ��tbIe�L��.��{k{��̪��U��!C���A�+rUP�N�5-Qlr��)ڽs�[�b���8�\���=��{�}L��'e&��<}˗�(��~=�|�s���o��V�'<}t}޺�3�{7?,�������߮lz����c=�:��wo���c�mŏ6�yv.dQ�	^
��O>4��6�7����x��b�X`Ǻ)2���g�=�~>�*����6�ᘆ36<^,;q�e,���vԼ�-��� ����b��R�WIF����ʞ��_-�8'f���[t�4t�no�=����3�)9�vz�Ϲx*�.��ķ����P�Fg�&y���U��Q>����[���F.�y	�/Q�H@��N�F)��JQIa
�;&EKq^�� �cX�b����������I&ϮJ�J �Z�EI;�V�6viP�R���o6I�L�7�� �T����r�L1?�-<�Þ���s���r�}6����KE#��i��e�N���N�O	��0�x���,������?nQ'Noj����I5e�.�7vp��|z���<[��g��plȫ$���O~�؄S]E�ʻ;gc(n;����K<�~݇�^L����/b��ww�߇�[�A. c{|���4�N�|�'/��nt��y���b��� �o��|���Wea�-:������i�y|kys���㥠�(yx/��l�l�Čv���g,��Xݫq�H��q�e��Ykx��0g�s��t�!���B����H��<\N����1�
��
Cr�,`ݤ�Bbڄ�=7w�����AUn"i��c8�rr�<�n�r� :�+�I��e�<������X���W�i���V?e>�^�w �����M4I��_.2ӡ
a
?ty.^�w�_u��ύ�u߶�[�f5���;��O�|w�rx0�W4V�=+��Ͳ���24�sp�=m��:�>�ڷ�rΏ&�Ž��a�|�%�r�Wp�׳I�o��`��P�eo($�qP����Ӵ�[)>a���[�l={8��±vw�c^]��Q��w`��w^#���4�C5��7��1����O��{n�`�YM�v���m�0����nR�n��4,PUb/���υ���kU]�QX���;+�nC���ͪ�S�{v�>nߎ1��m��)�#/tF͗qF�/��=�<po %��Z ���7�@+=փ��Ğأq�o���+u�ɷ޾%f�u�1�M꼞�Z��w|ߺ�b�-nt/���gs�˞��?j�m��ޭ�8��9�&��{�,�e�y�yg�mq+����K�+�k��v������j�ЯyWOT��T �F�Z6���Z�	��B\影u&��;;��fN/���{4�4�� 	:�����%LzsV�}�J���g�i��;�g��v��v���+lm8����EŇn��r��pb��=�:F�y�ũ�|��f-Oy�҈�{x�wm���}�]�h��o�|k�1�ӌg����CՎMT���#`�<��׹q�=~�ժQm���ͺ���f!��f�tKMF R������/E�+}�͘�Hq����kcT<�FM*w�Jr�gu����0��0�5�� �_?����dc�8,��	�ё�ͅgLc�W@D,�
�d�k���7������{7����M���&V��, ou;��uoH�=O���=��3�@v�����\��+�tw��c�:qp�jA�4�S[�~|�	�s����=��~��p���p��I��u+�[{{[=�����\�/a^�>��ky^s�q���;�Ty0�r2܁єr�Vu���KB�
�t�7�Sm���-�ͭ���Z�j���WY�3��(�H���	��F�fE��X�$�nY��w,\�kO�z�$mwL"ӞL3��7���c���sm�E�*@,�;wq��b�\�  �L~��:�v�8(x����n�x^�"�3쇽�*ε�#��mk��/R��ב����eKQ�Cx�#@��m�ۇp�i,�f�mΒ�0��P��2���ʼg���g��f?����?�ɒ6l˼G���C���Lta�]%���=��e��[A(���ʚ�7�r��Ҕ�r��[�M�w�~�_<�,���v��;���ֳĐ�ާ9?od;9�~�>g6�=���q���+|�{ɺ4����T�N�V�Kn�M]+S�B-٩(����7V����$��N�Օ�Ԯ���;{z��V���`3z�FM>�x���Q
}-�s��}��=���m�����o1�� ��6H�@��U���d��O%��l|�������'�y����E��:wc�b��s�_�������Xso��S����f�I�&ˤ�
4v��a��U�=�nG��;����vj��%z3}�.�וx;F��JC�p�D���=t=�m�[�-unn�x�,�Oeŕv�eP3L��t�ɫ�v�sN��\�T&�#g/$:ARY��:�[�ѻ�=�G�G�ၾ`��/)/j���h81���rwG<�!̄x�1W�/s��2�}~���"�(��("X3Ϻf>�e4���D�a�W_t[��^p@tz"<��r�s�\5�H�K}%^Y����Iݫ&| �$�p7��'b��ׂ�{��/��5u�q3���C���t����A��uS��כ�&mrA
��������|ea0e�8���@�ۓYqB�nXg}(Z�� '��1�t�V
��Eމ�&2!����㺞�}����ϓ���7<KR�s�u��h_I�w7�(����E�0ۉ򉽁4����݈�u�u�}�cX�J��� ����#r��w<�͍��=�'L�	�8 O���]���,u�q!���)
n��U�z�7=A]�S��6�3"j�������]����o��7������Hm��Y�V;�s��ý�a�a`�g�K��ۧt��[�$7D�B�ޭ�gU�K6���c5dL/5x��(���G��\�Ob��/IZ���b*T��Su7n-�2�f��:����xy�颴�p嗶�N�)�P�
ASjf��[�ea۩��ѝ�ޤ��U��o14�{ڭ��ާu����r��y����LX��.*��L
`��Ơ��ld�(c�+�f�3ޮ��M�w6LE{��oi�d{ٸ��Xx��=�n��z�{ ʆS,A�3�yT|</|M���OS�|-�M��.\��K�˻��M`�_N��=�=X��nkĔ�GTU��|V�L���h}���f �W8����w�+Ė��Z�J���[7�U	����r�S����N��7����ک������p���K�ۗ6BQ-[�T �T#o.�M�,9�:66*�\�5�j�:76��J�K�hi�	�{+����j/���E*q�j5���°{��m�v��N�i��A�#ż��Fz�nYv��	���&�0U���N�R����}.0���9��+�<�彋ֲ��q��g4`�@Ň�������ַ0^4���/6FB��D;�x�g�=��0ޯ���ǝ�� ��!�d�,�U�	y#7�-	�gM���b�kq;���ݺY�%y|bC\���㳱n�rݣwG�6s^I��y��C��%�O��!�ç:��w-�OIs�g�<5��<�ޮy&hK|�jc�[��T�k������M�jkdo�c�����&��]cя&��IV^>�Z�袵��3;ػy�J�R�NU�jKܹj%F����$S-G�T����,�gc�A����:@��+k�G�48��>�=s�c<p���ѯ��ʹט~����[1��ύ���T<�yxq˰f�ө�v��}�Ӆ5q���mM{���gS�����*�?o����eZ�	��9���>����Z��թ�p�nǺAFe oΙ%ʸ�(�[Xz_�D��D6�ڷ����6����='�K�ބ{4�xOy�9v�Am�
>�س�����;�En`�WE�j-xѵښp���AӖ�YO����{P��ja:���{4l(!/g�I��x��ׯ'g�}p�y1�,*_^����c�LGq��)M���%<�G�i�K2	�$sw�U�|�tN2��+�	ޚ]�����1%p�=��0���X��kϏmE��+`�1��҄ʊk.�j�[85���PF�*�jh�ZW"�S���b�^�{s�;|1.���CP�K�+�l���z����v�Q�z�8�������#h��2\ҽ�F���u�c�z�w�v��vM���.ԧ�t�Bl�cNx�RW�/�1f��5Íl�pI�d8p)D�nieצ�]�F9Ew�sw�>p'��Բ\�F�р������'�,�����Q�:���f�X�BL������+��쇳�9�r��{�~&W�y�j�zzv���v�Vxg�����>:��9�j2��"[�ldy��ɛ�J��	�ͺ����-���p��W3{� Fh�	��(�y5�r?@q�]+�;n���7$i���uiQ}����D�YK!9��u4^3��\�Ç/Q�h�=����+�Ő���W1���y@�ZH���d��[�.�����$�G�un���S����o��-�Ta�|�ڶC'Q�݄{e�
FN��B�wt��v�����"����z7F�1�\���LPW_���y-篩~/�dK���-y�W�٩��Wr�a^RF�\���Nl�sY3��"#8J=-�	A.�/nT}�kw]>�:�<O�(G�tnF=����s��'�7$͎�^��u{��ޖ���Xt��V#�yd���庡y��i�I�eX�J���dF^躕���T&pl��e:ɡ"�P��Sc�\���şX���M��Č�{Q{a�w��x����{��;�Щ}�JPtL͎i�vv�׽�{�����Od�Hl�=��f�g{�%��gM^�H�@�`�à/�g=/��Yǹ�=�yO���<סg<�Rl��x�ǂmd����R�p)t9{�4�ӌl)�ye�/[�}8]�w�*N�k;V�עBLR�WPr�����A�����v�y�ގhҽ,:��9�����K0���z�綰�̼����4f��-]�|���k�z��-�����*6b��Tq��=|�ag:�`x6�>P��y{��]�rL}���Q�;N�Y�6>( z�������;9�/
<�2-�՝���:�&BA���/rs�:����I������i4�Z���K���k�cǦ/{��t��Z�`�(]����x�i�)ƘW���=}���z�z����&w&�Jg�^s�^By��c����sh#ob��t�~RC	Qy�=����B�āX�OU>�;0"�s�ǳ�IdZ؋k�w.D�#��.��ˇt�}��-��)0�c���y߶
�4�L:��k�^1�����#��'�9!-�bc�?i��D�^�r�'������&"��}���9n����1��e�aEL���f�7�q�U���w譄ͭ���͖MVԛx����x�^ki	Z{:|n��ަ��x�uBZn����Cr�#���;��#vy3�zm�{�^��C�-V(��X�X�t�1I��L	�"v-�-N2,�ж%�Q��߁KǼy�f0��������%����u�w�vwl���=�X�s�/�M81M�(}�����U�v�^�U2l�p�rn�ݿ]�$��r��{��d27��}�(��
�\<����g��D栢�G�7�6=��ɞ�i��=�oR�㾑Mӧ9E�l������ye��>LO	��,N݇�I�ߺ���1�a�ۛԏ{���B����ǹ�`��o�*⻏}|�ԉtE�������C\�U�QcN�Y�3�"����7���g��Zc�Z�ؗS{V������φ>�{d�v͡r0Ř��w�.��O�,[�WJf��ilbݢ/5N�ljܛ,�gG1
�>�1=�9㯅��{��i΀��k&���C3�����[8�[��Š:f�����D��b�=5�2F�i��LMwR���Z��/xn�^��.�f��=	K�6�lR�E�K���<6`=gr�/�?o�x�#��o��,�(�I�E�Ë�-#@�3��������o�&�ݹ�bl���ŏ{ό	)|�� 哷�X���f(����zB�
g���P��À�Zyh� #��/ѿh�����/8O�r8��(��i�>��ys��hwT��Ƃf��Ȼ��^]��:���Q�kB�h(C�C;�E��T�|ǫxƳyL�F-ߝ��> c��i㬧�X�KUb
m��n�e�',�A�hj���A��"��5�����1��=�:f^dML�PB`˳��=s؞C�E����zGB>'Gw�"��%�Ht3 ��<#�z�.�m+�ĳa�����~���NQ��U����}�[��
�2.�"��R�YƼ��47���ڃL�x���/X���{c��=�[������00���%�mU��!.���Ed�F�q��6��ُ}������Z����_��5j��{ͻ��au[�ƧNC@nR��N��	l�5�^��qG5�@�3�[�(|v�hٹ�O`��"�ۉ�/�輺I(�����ϧ67Y=�ḁx-~}���.�n�麴�dj>�`�:�)K���Z��`���{��wv�����y���F.R��Þn���.�FY�N��R��q���d�ě�����R*&Є�d�n�Mn��Y����fX�P������1f�׳��V1e��`f-�f�6�bgkj��Z���[H�;vh�ƺ��;��F�g.ў��;]���.%#qL�QldfmZ�F�l���5k�<�$�+�rLK��U�:V� n*�fP��F�rK�k2@)Z�0%��)�T	�kub�6����:���3\a]j��d��->��b��=���^g/A�u��X6N7m�nd�ݻQ���]���ez}/f��:�pm���\�SjK��
e`���6����pg���t���([.l���.H��۱�nPB�\Wj��ۮ���u����u�P:��l�� so��IL�k�jl�,6j[@Ŗ�[ŘR�5ꮵ��L3ml�GK%S.d�G#	y�+��w]�,n�Z���X�J�ֲ*!�m�R<LL�v��t����rW(�[�n�t��Y�����ֽD����@�<��=����{m�8�V9���cc��%�\�Ǘ�{u�e��t\�v���(�h�KsF�^qk��J�����)�i+��1�˓X���n�dQ�D�ڷM+e�B�\���쵲�����eٵ	��[C2��vv�h�� W�m�&��H`ػQM_	Q��dh�X���lm�;�\�mϋ���Ow!f����%H��k��U�5�M��Z��K̐γSDQD�Z�-�04�捣�\����Z���l��e��&OQ�@q����k�n�v���۔�-�
 ���5(�m�[e	�J+[-�,�p��sŀ`�b�RR�:e��G\G��]if��3p�0�c'c�t��xݰWS-� !�G(M��l �<O�u@�r�O'fwu��t]-��<�йZ��bK��[[Lv��[YJ�����m�>��lvv$���aTΎ�nUv�0�:	a;I��K���b{lI�L�4#� !M�sk��r�"b�;���Ϯ���T�$�^�ܥԥRb(�m�ny8�p��M�7n��c��z��l�Aq�^����oV�\��t��� sF�S�Hz�majCk)01� �&��2�tY�c8�-2�v}�$�W��.�r�ݞ�Iõu�
:b��Gfk���$lKh.4�����hD,���rD%�n��\��Te�&���|c����S�cX8�w!��m��3�����!r���c�����l&) `moKH-i�ٔQp�V�j7'h:m*�tHB��֊��+��a��0:�vĜQI��ѣv�iK-˂�J��*�&.ڄi(�e�z����] ��oO)���9�`�r�5�rb�*�f�4���o!�Q����m��e�k�A�����nR{]�4�X�T]��em��}&��\:��9�v�Z��g��<qv�i��n�+�ͥ�͌����P�N��mT�bW�pvG��P�.+H\�eL��:�XDn��f]ÃKG�2ۮ�͡�Z��a��nٶ�瀹��[r	�����V�@͖]��+6S6�Ices� `QR���=���H9���Ʋl;؃=���E���\\���i6Z�K.LԠ�0���q3tR��1Q�ˮM��5	Y�Ϣ�+��d���oB�҄�a��K�Yt����0��(B[
׳vنwm��\��JЊ��qL�4.�ۘD����Mqix�)��N����Gdn���9�������:��q�<�k֨0ƺ�U��KkK����JٰU�!��]�1��4c�C�ĳ������-�ܝ�� X�ǣ�i�2�mԤ,Iq6�1��d�֎6��ez�T��mc�fɵ��J<q�Y10(ҡ��۸�W<�$�=q����F��q�*����̣8Ze�m���]i���c:_`�Ȝ&ۣ�l�g�q���n �V��0lΙ)DSQ2�Ƌ<��p�6Un�o4�M%�M�6�!�1e�c�k����#����[�x�RԝV�I��>[��&.h4F��+���3�w�E���:/>�7]rs��<Oc.����ϦRy�l���ٚ��&�%�
�X��	�-0�b�Y�l#�V���ȗA��	[�&^	�[T��c.`0un�2�L\lm���P��5�Lao�K���V�C���n�}n�9p��^��z�e2[����^Q1��#Ö�m�)�K��f����u	�+j۰*��L٫L�e��e�v��7��y�IP(�v��+�s�n�k��.":㝂�Y�ż6�
�-��"3e��P�16�4�ƭ�M��yng�2U���-�����{L���<�vf�8ڛf���:�d��(JLt������fʨ�\�n!J���l���Ur��ME�2;�ld��y�a�:��e�ÚY,%:��|C����9�v�g%�Z�5fJMh�(�-z��u���b��L(�u�����t�6���L[6�=��jy'�B�e5�/6�(#3�m4͔�vMO��y�z[g�ɾ=S�-J92lh��E�gE8�&�Ù���Ƶ�I���/�(���,E{]�qp;A��OhrN;Zwn���1���GMl�Q�!��TA7n�ݵ��6���������"�%�����+*�Q�Kr�M�G�%�"�c
�Ћ�3AҦJ�ы�Y��i����,D5l#V�-X4L[���fm(0X��D�i`F�5�����c���;Vf���q<�:z��;v�<���ۣ6�3wgG��W��-�oR�Ъl�,,���ĔJ�j�\.����:��
�m��bͮa�x����x��r"��D=@�#eBfQ �M��3�R����J��nwg�h�y"�m{)smN�KW)D�9�v�=%g\l5���w�t�nN����+���]��#���Q�+��\��].�A���YP1�i�ٽ��m�"v��霜0nm�x�XR=���
5l�c�Y������@]Vb;�u��c��&pRiW���C�+�u��sU��s��?�u��(v��qKsn�n;.9�IHK43-i���lY�5VZsM�lc��p��z��'�b�)��oY�.�3`��7m�.�4�t�!�Mq``���su���WF���v�a�!.
�q'�Aۧ�Ϩ�mn0]`lu��[14��v0�,��F�i��2i��ٌ��cu��
;E�62Ƙ����$�c�XC��q#[�!�1K�s�ۂw��'Ymb%�!���5z�&�a�$w{J
��OPs�[V��Z�]S#STm�rĳ/0�kF�3.�s4���+���u�m�(#c�NK�p� Eq-k�c\Yf�c1I,*��m�R���g�ڑ��(�6�i!��^�m��>L��py$qs8�ooVL�<��@s�@0�݋f���bd�A,��(:h��N!�i�)�#AN�9Ǟx��
7E7lu����������8�l�*�M����
�rnۗj�[p�D��Z6���n�46��x�%O;2�<F�Y�s3��CiZ\��fI���7)ex\fꉮ�����C�^۞�������Z����#���Ŭ!/S�[i1lX,�,��c�ԥ��a�J�K-��Mn�v&�Ғ��#썠nP�����us�c�	�E֧(GC�w�]+[�o<��,�
*��,�h7n�"�Zx�/�d݋A�f�t�\3 ���M���-�ĸ��svA燙�w6i�s��z��Q͞׋��L��x�q�k��Y���p���X�e��;�12�0�c4��^Z0�l���p�n5�#�-4�]b37�r���BX1�\;h8�bd��ű��ݓM�7"stGk�f+2km�]l\��l ������uОn6q ��7A�ka4֥��oS8��v��H��
��,�e��a7\��w>8�t;2l��J֔���CL�
�R d�P3V֚9+]�w7`k&�`�;���.��
)X�v�.�vFK+<����l����2�]s�N8e�9��듷mX[���ͩ}���ٓ�&�vU�rx7Ip�`m��%�vz]��I����8�n��Ms<���y��V��-p�P�A��X�1��vxw<��5��x ��e l��뵕�sl��M6��U&�M�iKac��V̰n-��[�Uc��Ac6tn�c:l�%o`�\�^�/�o���y���ݩ,Ԗ�35�Ī�h͙�H��J�R][4���-�Bծ�Iq�v'���2n�R�4I�uhp�j*R܁@ZJ���R)KOG��n��+;2O]�WV���c�om+!n�ҥ�:�Vg6�[k.$u�k��q�Z��Jެ������D�/5)D�����ܮ�%z{n���٧-�!q$�[NBi���IY<|e�b�\Gf�i��f�j�(n�Cl���T�8{@�V�0�6-��8��t�G1��9�.P�&���&�1��PD����f������ؕn��R����ѥ-���8�s�րz��3�'m͝g۬�p]�݋����p��T��\\e�@m�U+��$ڥ4��|�ͦ{h`Ld�D6۱���E��[G;�[�r��	�۵�s��.�6�f�|�m�fdr̘C�X8�g��,��\���0W2�140��ɜf�l�"!Z���CZ����F�inN�;��{�#��Wиږ�3�	Œ䔮��ꋦ� ܒ����$�;��[8����i7.9�b����X�XM-f�m+,��� ��� %�	��t�2�=���{�v��I5�} �)jw�	ك�Ke3h�d[�F
��ƳL��c>}�r�QΞЦu�A�#�paA,l�V��5Īبy���x�Q�L��M5Ynj�X��j�J	��.�r��ƺ�f�������I��2��fr5er5e��ݯ^��C�@�q%(,�+8ӻү ����)*Q(P�mu�e��ހL��<ӒN��	��$���=�Q��=���tG�$NJ�YK;�#Ͷ��c޽��Dq�M�C�r�t99ŝ�Е�g�;��G�'�<����)�r"^^'�ܤp�/F�.tr�q���krJ��y����޷�a�m�c��%L� ��'-��9����xZrͶ���I�np����mۜ �c�<����3�"��<�Om9N��ؽ�y���ݵ�圍�����X�� �.��^�I�Eb��0#��$�e����҄��Ć݁$����a�ʚk)f���V[e��Q9�����-�ck�[�%�E�m�v݆q]��GV�n��v�VR��(��q�4�\2�������ppgv�{[�
c�5 �f�خTj�ڛ`u�h���c�B�[�mD�B�]�Z�6֔�V܄�p�i�[�X�a��&moe�s����XW�:��\��<U:��	��	n�J`��'�`�+	�&�΁cl� ��\�v�[���p�rg[�tݞ��l�%�9|㘬�٫�݁�σ@t�ȍv�Jk@��,5-�ĥy��D�=�����j�n2V[��DY�:"0�,c�&��\�X1)aaڌ΅)�ՅqaU�nl�U7���`2gǶ{r{�����l7l�ůj�XĆR��F���YcB[�p���֜d��W�y���8�����J%qv�����Z�0n:���Ur	��m�Ч�����@�69������X.4�V��C)���ʈm�4�$@u�j�Y�0ܗk�0�NP�gz�[�1���{
��H�������y�8�tc.���0V��1��h�Y���1jbb�#�l���o*nR.��wBu���Q���kp�]��[V�!0ݵEуD̲��tҦ�-�4�H��l�]f�9:kIy�������'�� F�ٛ�6m��R)5 MiZS5Rc�u�6-�[�v��U�- ��� �hAU���N;��gxy!��<=�N�$UȉM�C[��=�[��������.���׃]1Hh ��3ePt�1�٫m��ˠ8,�n�J�n��/^9��R8���V�	����oQ!]��W)Gj�U��mC�4r�K^&�I]�	Ys%pM����<������L8��X۵���� �R�@rl�5��cb:]#[�H�f����kr�	�͝��B�39͠��5C@,f���7XЕΝ��i���=���)�	��q�v����=��x9\C	� =����s�ϑ<�]�&0q���W�����N{���`vO���wcȽ�������yWp��s��=�a}���콑���9��Ns�=�'�&����=�q���w�!��<��Ev�{g���__��]���s�&���h�:	M��nJ�9,u�/Ju�+�d�H4 Ho�}f����N}nȈT��b���*�u����E��0��1��Ƿwv��xxÍ�s��]�ۜ���6�i�-s�<7L>�!M���nۏn���u𷱙z�����V�'T��c��ݱ��Q��)x�Jї� n���FxW.�3�[�����ޟ�@y����2SmV��N[(2��o^��z)���{Z��71i�}���[_s|=h��{�)�?b�,2<KoF���"�������2j2�{B�VQ5���Q�_=ˏOv���%�xK��q5Ni�O)�=���^9��/�6���&��N��O>� �r�������O6id��G=�ɔY�Ɉ�#r���K|�L�zj:�Wv&"ic˚�Z/-�6TƚI�	�f�^]��"���ڔ��p��|������<1l���ݨ{���Z�j}�v ����i�ͅ��V�eZ�^�8�nb�\�n��#vΒ�.��c�K���Iu���t�Oi�5�O�j�� }y`őbqw��-��M��}׍����u~2V9���������㙓��N[����Y��<qҙ��K.�կ4cA����D��9�lq��7msT�u\ �ݑ�:��������cxO�;�-��ͯn������dD13�B��۸�\K��z���q=�4�xc����O�-�� �t[�>����wF":깦;�M�:X�/SJ�2V1��6�^�B�Fyon/^���{2��<K��{\�r:I�]i}�ŗ���N�g׏׭��v7vFVD�ڪ�����#v=���;yk��'s�k�,�����-P��n���j����2�߯[�=̷��;�rg�t�OU�5������K�*�����m����a�g���I�>N���*�m�uE�P5lJ`�D�����o�O�?e�OCs�*���s[;����WݑM@��w#:=��#v63a��$t��;�:�����\�1;���\������[{]D�c�5}��݁��Q�އ��uU�T��X��'����[�����7V�L��7B<z��;��{wJ��p�����mn��+��J�v���B�صŘ��xU��X�z(��oi};.�gr�#�ǵa͡Q|�����͎��Gj	���I�ڽ�̗ t�E�q|cB��ݐ7`n���@�y�r��!�����l�+'���_)��Db鸱0���{��y�kk�ZMe�ms��^�,����9=$�[&q� "0,^37�g�+N}i�?�w�����4�i�|{2nz����n����761��[�Q�ӟ���SP��1[[��=�dn���Q���G����ݍQ����Ͻ��X��k��{ˆ����'s���>��7vF���j�;7 �r�{v �T���s�Tҙ��޷*�Up� V���7cۻ>݁��n댚��<�T��b)t)aM����mn��V��{ww0nZDU�wt���:O��o�Y۾����\G�:
�n�y-�ӯ-���{�~��T��7��z�3O"H}�8��X�%�2"7�vNS�m��6m�n�5��!�ɚ�&n���U���[�^��/e#v��D����8��fI�6�Xzû-�B�P�B�
��]�4���3�l�u�xls��z�إD�L��R�mX�9���a�k���8��VDvv�8�F�N�箝���{۞t�;,b;�u�p�|�fK�M�\�����u����~��`��`�vK�����X�'gh-�y �(��Փ&B߀���>݁k����s7�N�=<&&�Rm�' n��v=��s�9�s�d��t9�E�RL�y�mS���>��u6����:}��5��VZ~����
03[����յ�~b�����.�e���n�ݻi�.��o}�OO+c��O�}��ͽ3��O-s�g1v�U����ݠ7vw`������K�q捶w��Y��S�3Ox[��7vF�j�|�8����ˡ�0�È�	��a)�mfvt5����K�ke��rB9J�C���s�z�5��ݓ�>��ܝ\"��D�Dq�0볪�7`n��۱��D�j��{{a.i��q�a���2�`�̺{�#�s�h�wv�n�wywU��=c�Q7�ֲjMn�"&k�ʁBW{�GMw�s�'s� ��}�x��'�^�����^��Qo�B!�sF��U�6 ��i�ɪK++osOWEc�j���S�}���T��9�D�.q4'�~���e�U���ϬoH��wvj'��\��+�kn��	����&D��4�s�����G=V"r�D�9f������>���Y�{3��"}7X�\�1p�bw1#�%k� �>:Dn얱�Ԃ�uz�g����3�bT]*&�v^%�!y�\��9�۴�	o(�Aݼ��~:����c!��� �z�m��qY��S�3�{"���B�9�u��"n���sQ�,��P�nϵԇ]�����@"]5����y*Wx�ݍސAG�#VРwb���L��z&=V�xP ��ݺ�f������-}�����Ɓ<�[w�&��Kv�3T�ХK2K�W8�L�v14Yf�F��o��QI�']���O�AUD�u5�C�+M�rqՆ��sX��C����qȟ"�wf�F��j��������E�Ǡ\.oO[�Φ��[��qǟ!zk}��{�5�ˏ�G������Hb��Ş�wT��c����5�cv}�k۱����=Uɜ� [yf1�wF�3�C$[��cۮ�O<qu)��\��	l��V��%Y�����}\O�R{��牻"}-�p�{��cFw1 u���eNou���'����^s���.�<en*�L@3IV��J$4�-�7�泩�ǲ���}j8�z�њ�M�=/����x�"�����\�hF<�/�w�v�8Y�W�|����C��L[v7xH>:~����J���~#-���J�;�*�f}��n��x���_q�Ӝl��!�q�h\��g��EY��]e��ݬ�+3A�'iC�3eV �zxw7����?9��ὴ�y��_bLa�dȄ$<f Ogla��E��#��}4F�� ���Рwc�����N�>�%)=P�k:ڜ{*}og֣�AG���j�ӈ������H�P���k1���j���p���u�ƭ���R=q�O����ݽϽs���s���׼=�����ݍ��d�Ɲ(��(Q�A��7v���5�Y89����W^>}"e<�Þ�N1�;����Z�#\��:A�]j�9ų��4����wv�x�Ǵ��S�z�qB���vo%ӳX��Ǵ����{IG��ϯv}�
��N5޹�t�:D�ݘ�|�l�$VݍސA�����;ɹx��Ǿ8�F[[�҆��-�ۖ[�7�+�n�L���:���2��8O_'�_,B�80j#xj�����۷�r������ũ��Y�OeY݄`hn,ty7���]|��d�������"�`�ܢ�qTQWՋ���s��ߞ��4;��F)���'.СfY��M�+��F�Z�j�r*.��m�I�w%����K�GCA���n&�c�K���n˛��k5t����b�)�4�N��4k�-��u�Y[����!
s���X�ltЎ�ZA��zL�����!�L�:�.$v�k��&t0Fn�!l�^�ms'Q�s���]�muƫ�h�r(8��=��>���xs��Q�f�.�F���X]��.7m�vb�YE�PԚ���~�z:�~��ؒ��������v8X�����o�i��;�?d�k�ӈQ�E�1��!Ƀ���(� �y�М��|=�U�Em�݁����[B��s��C��6�~�6̂_w�?r�T9�nj'9g/�6ϺЫ7�d^,�׽��6e,C�>���`�X�F�����~o�������q���<��ښ��+1ӏ[ޯc�mJ��gfm����wvh�$����%����1s��Bݥ�'n��	��@ ��^<�2���'�ږo��M��ō�M��燵�<��g[��.!��Ma�����O�f���w������B�wdL����^�o%3G
�Rx�]3`��[�s���|X�Bb����׹�������*J8��n�qu�+uHs����0pX�hછ����w�N&�m���w�&��m��^�v�����k��{�0��[���ښ��+1ӏ[ޠN8�Q�#ws_Q�{�}J @=�4A���H�}���s����P�م�|�����>��[^݌��#wk�*����K
b#O���B�F�m�p���d�i!�p ���#��,\=A���s@���t�<A�B��8���\0pdX��f�r��ֲZ�v�����$�xn��ݟ�6���q��� ���IM0�p|tn)�t�U�L��qQ���Њ�q��K6�I>�}y����E;�4')0_3v���;t7x,�r����:����E+�;�)������{���CZ�WW�Ջ�����ֹb�b�Q���P�"N�ۻ9Wު�Br'��wk۱� �z�,^F���9[��Wqr5U	.]�qts��4��c ��0.�؎�1���a��gW��ǲ6��g0N��:�WQr�*���d���#{J��k	�����g��\<ǔ�6	]�'`��G;I%�ǐ�e��;g��>ݗ|��<#�KO���)�K�\��8�p��	x)}����<]�E�ׅy;�P���B4q����1���g���Y�hn����7(�������\R�ӕt�(l{B�cR��b��FX���L���4hR��K/�:W}����j�UΪ�rg�<��Q�n�P��~{�qD7�ku�{�&��|����^ݾ�k��=��g8}����m����-¿{۫Ǒv���^�C�78���:u��⠟j�������%�����Y<�/�,>"�{<�8�=:�^���S}z���=��JF�a��]'ή�wG�T{�xzl���8*-V�5 ы�����v��wL����=���A���@�����𾺽86�E�m�&�:��p��Q��;.�
 Nuv3|xq�ꐝ����n���\�[�4�w-R��L��{ۅ���sv�8J�İ�!{lLۥZ��e,�Q����*����8}�A��ç�������۫�������F�H �@G�ា{-�ƞ��-�s�en��p�x������p;���E~Y��1��DwZ�����t<�;�y�QKgۀ��|����!٤�yxMӃVs�����w�5��ﺽ:Ý��
����E�K�9Ē����N��)8�lt��r ���^qݗ�ZK�/m�۱�YGgi@�:Eiq'@����y�\��N;��y���8��浩�tI9�aDve�W�GqeiٝDm�ģ+��G��Zu��n��\��A��[�^ն�2ӤK-9:m�tQf�&�EÔgY�E����:8�Ύ�m�Y�a�ٷZt�ܬ,���/#��gMlmݶ�E�������;5�w��lGv[�Y7��,�y�V�и�B�J2���٘Ts�<��&?�{��n��+�d���ǭ�ޯc�#�m��N/�~�Ûx=���Ɍ��E;�59I���y��\	ܡ��:}-2��k^�,q$3Ỷ{v$�6= ���N@�n��X�"g;^��Mob�b֣�)9�:��E;�p��/Ď�"��7 d-<8[���ϡ�M,�mӨ(4n�Y��3�r[v���g���;<t�ou{v0�6=��]��fK[m�z����ȅ���zGG��5�^;�$"���!�͍b�ʧ�4\6D��1��K��o���Cw����5m{v"��.f�Ƈ�@"���#O��ݪ����mù��j�[|֭x��Ũ���S���r'�H�Awf�ݑ#&�uTo�c�P ��E�Ic��[[�k�䵶�G��
ۉ"�"�N�Mا�qP��CE㳥Q&����+�w�^P�<����q��܊����Rvwbr�v`��㤗���(�$'�k.{;s��G����<M���w��d���',�V,;������H~���)�C�����ٿ�x�>? F��.��z:n�ٖ�\\��TN�Ga�J@`��{X��L�v<Ь8�~������=?�Ž�����e�1��UR�ݝ��~��[�@��s�,^2�}]m����`�D���M��k�䵶�G��
���
�A��\�5W�T��%�̽�[ĠDy�_m��w2&�/-�㰴���ѝ��ސNAK�����~82��?�'~x8�k<E�}~ݑ3����{�S�KQ�ầ�C�munɌب���Vm� �� �ِN�����)u��v�?\{����yVKT����������F�x��q{۞X�I�x���l���N�=�!�ڈ��.m������\����7�s7qu~7�f�[�t�[��WZ���>d��4�j�l�3~ý~����Lћ41��K��� �w���%��ҋ���ݻg��� �����Wt"ha�S.lۮ,�Ǔex�l�um^�͉�QN�9�Q8�{����>w\;�ziݓ���� �i�`��j�RMF32�`��0B։�P�U!��mv ��6����MkU��ͣR�2��<���Ʊ��7��setE˶�4)��A�z��߯=�������z|V�*���-y]���VX&y3.�MJ��Y����/B?z�H�9��')�Þ-.sgv��z}w�7���ͳ�D3��̯�9R���#�U�\��d]���i�x��%"6���kxbs	j8GAI�ND��x:ԓ�1�o������M���(9�h��T���b��r�|Ohs���=��%�M�M��y�j�{P�9��y�,x�1�Ϲ3]}��|�t�<@�ݚ��{.x\���ѝ��>��!��q%���zFg�Ǟ����'9�M�U��*T��q�R�;��z&D5��'JRG�A)9��>:D	�٪������Ϸ��~���pZV�=���s)AG^{M��Ћ�T�QٳZ��4�7��Y��u�}|{��@��_u=|1�)�r�y��7��&1W[|��mЯ��G��vk�c'����43{\e��CNn�b� ��4#��(��>���<��t$l��m誮�ɝ��� ��u�����5=Q��X���r!�^�����"'>SBs�\���nf�����>�F��Gv*��+����H���W��D�F�A�>݀C���b�弬�qv0�:�I#��s@��I�#���ϷpH���\TBG�=J��;�/�������M<�S�mĂ*\��ټ����y�:�B�#�jx0Z��୤��I��}3s�f��.��u4fז�X0Q�����-?,�~>��t_>����O����K����L]Xh9ƕ�u�m ;iq�RZW0�	��c0����������^ nȍ��8Nr�
�����8��F��W���ֳ�l{$Ig�wf�݁'O����Z�y0�i��p�8��/_aS�ra��O��
q$�F����c3|�$H,�� ��gۧ&
0���W�.�)�~囝�NjEų���;������7��I�)���aн�w�ק?ޫ���%�B��Z�WT"��Sw�7��M���xtf�i�Z���3�Cw�$��Aմ(�Đv=n�P��ƺ+4_tQ����n����&���I��H�A'5�]�� -��=dMM7fA:}�n�
v�F��)1�]Y��a�i���y�	�!ǆ�دՕz�;��	���)a%�q ���# �т�&�&������zn^-��F��~�.h��S�"�������k�V�r�n�݀�D�%Wg	��(�$6=#wdP;� �K��o������5ȝ�L�]�T뭝j0���Nh�{O��L�|f�{f����'{v1�
s�4<�K��V֭��
�v|�L�ӹ�<���/�)9�kQ���B}������^��� � � �����l�
�\�Шݑ��A���q�:el���`��*�G`:JTf�"!Y�[��[�:3��'���?:ʹ�'���:TPp�.�暵�%��_x�{W�G�
<7v����n��5�e�;�dO���F��u�εG)9��HH�n��3մ�\쳱��$WU�MaVjf)\ʕqv�kk�Q�D�B�D!,Ͷ�������:8�D�{S���ʕ��_'�e�2�N���C*����
v/���u�"N�wvh5>�b�YZ�F�">/6kӝ��G
��ˡQ�#v t�:��x���e�p5*�����Qn$��ỷ^݀�=��>��KNg]ъu�εGx��Rs@�܉:DN�ϷrFi�c����B�v�Ǡ_ub}�_(�-��O;�	�E �]_7�����}�Q̲�%Dc�r�#�>���"g����3�hJY��8Uw1���s�s�=2�Ng4j<�\D�D��*pJ���0��M̽Ǻ�H��p=U3س���Յ�H���e�~��� zV�PS4W�§[pᝧ.��UU�k/&�3yr�)�{���"*�� �M�Oe˺�`v�̻��ktkA�ɪ�,��f����nA丶�D:5���y�m�hd�6멶��3��Զ��j�����iz�][C+v�V�Ip�F���61���B�D6��׮�Y0.͆�݈N^Uۮ-��[/T�X�����.�r�e��.����i�nǎ�}����ʝ�k'��6.��\1��陱����Ƴ�Iɭ��m=���Ѳl��5/Ku����T�d�
s�{�'���F�Яn��Y��]�]��Q�W#�mՌw��7flF�YA;�4F��'O���h��0��s9{>�Aq���;�/�i�ڧ~��8���wU��S�6ԿlG� �y<���B�?ڈD����<�nAV����WseШݑ���AV׷c<F�A�^���<�V(O����29���5�Gr6�F)�{:�aA'4F\XȞ�V���k�۹�>�Рwb��CVau��>��w;b_li�ڧ~��^�8�x�ݪ����x�'��9�'	M�I ��^�*�k��:闝��E�h&y35�B\a��|�y��x��"|t� ����|��.�7�F�ޑ;7�j���s�T|��P�yD�FǠ��b҆1����L	����Ĉ.����r�\�=݋FΓ�vF�ۃ�E�v�R��0�BL����Z2fX���ڼ�z�&0��� �|E^Ux�~� o�s�E=�ݝw�֜#�%'>��I�)�\U�z���]�z���,�F�Я���J�A��]y��	OcL��;�<��O�g��B�@ݑq�Tcվ;��w����x��9ɩ�yϮb�8�j7dn����UK��p���ؒ�����ؒǠ�ݗ��Dg�8��2$>��������ӄp>Iϩ9t���we�쩫t����aI�H8SL����b!p�"�kQ�Ite��(*0�KnqXb��������ؤP;�$��=��	}��Sj���Yv�������O<�ba���mLc�W:w&L��p�>��S��}7\�˨�ݑ��A:} �["�wa�D!L% �x[��|S� ��G��گ��մr�r�@�*���v�oX�wY5�ʭg�`���xs@��'-���WWt��8��3c'wX�ڻ|j�x�J�;��yI��8ł�ڊ�� �5����s�cq�cxp��A)9��>:Dx�wf�ݟH��U�.jĭ}@���G�$���ݻT�K�e5)ߩ��w��u�����@��U�D��@wvh�7dO����c��*���MzZ��鸺�]D�����["�҆
s:�k�}���aQ׿������x�n�F0b��zF��n��A�v�@�+���o|�L�/d3�D���n���ݑ?#y���u�m�2G�W�b�-De��K>� ��	����	>
�E'Ұm^``���Ǡ_[�O���FSR���H��$C�G���7�A;�1�܌��Yn��wנD�,��Hǜ����ҩF��W=٪�H�uS;�7zA���/W���0e?�՗��ٝ�8#'B �����U�"CF󳛌�;�.�xd���9�1Y< ��Դ5�BC�2��T�� {6�Ukg��.´o�����76�w�]s�v�������1��a��&����"�n�F�����������'9E�e"�4i�+���V��,�G��|�����aL&�;�<�@��$\xn���� ��{$d��U���c�iLdҦ.2U#��2��n��c����ݕ��yx�<r������|m�����Awf�9O�����+�T�l��&K�tj�u�ʮ��&�� ^Đv<7v�@�wbHq�T���Q�} �����[�j����m�8�^9�N}�@{��uL�XgWM7�A<} �7v�x�ĀF�\G9�
�"�5Z���S	�N�/:�:����wg�7dHH�A�C�N	����_T� ��x�����N+}�f����3�#7� �} �	�s5�B��MtO�.<7v���ǣ�n��B��l�fN����w|�����i�0Gx�� �"|t� ���x]�!��z�3�W@�����2����Nu��iȤ�Ξ\��e�[D����H��=��ü���<�{�Liu\���=�)x|�Y�mt{�w�v�Z�{�{[ü�d$V�G���m/�ǯ�נ�ٓe�ܹqe�s[���:�_R�ٻf��u�;�d���m:j��S`a���fĂb/ۺ7�g9��}A��ԙE�7V�{F���|����T1�~��hݼ���Êy���:w��Rp�1.�r���n�C*qӚ�E�j�B�7�풌=� �	��)�6"ڹ�;��c�����*�כ"7i�T�On�{�j����Sِ3�1���*]0��BbЉǑ-�d��K6�ٌ�FB�o�^���F���۝���A�.���h�fq��^O��^q�⸩�x瞌~_$Sz�>��ѣ{n���i��5-Z��{�_Q�g�:�q�E(g�H{���7'sKx4(��{8NA3�=�N^��ɮ�˴u�3୴���ـ��z=��RCZg�����w�D����#�w�˾'�%�N^.�>��>�j�"4ɕ�!7�ͧw~gwwAcz��.$\	"���Ў���LèO%��z{&���xIW��Q���系<�[�*�oRP}��OK�xFK���8}F�_zc�q`��{t�=3c��و79���O{p�J�D-�'m斳�6]�wwuҼ|��v�4b���B佪�G״S+�nhx�]s���Nb@;8b\�D��1ӍE���So�n<��x�p����"�1��k��F-{�^f���,��9��^^pSL�l.;[I� �8��cHF�Śfr[o7�Z\ݲ[vm�:̱+mt�Q�۲׶��ѵ��а�m��t�9:�0�f�лN���gn�&ќY��.�lq�i���L��g7c�ܶ�#+m[n,�;�18�ֶ��$��β�vѶ�첓��8��ee'i�8�:̚�D\�kn�30kwv�
m��Ȭ���6Ze&��Vm����6�m�760觶w^tY�[��j��U��Vi6���YwgGu���e����_�Zy-��	7$�b	��:Lr�=me��	r���or��Z�[[aj46 �]o)�h���]	#�+-��)���aè��f�s��1���'���Q�D
��i8�xX?��`�|�=�=�"s�n��y�S��!�]����T�eQn�]l��c�AId�B�v*���\���͠�[U,LK
����0���rr��	8���gV�=X]t��^��&�[	����j����� �6sf�筨�J�҂�v6#W�uʯ3�7-�e�G)-�BZ[fl]%-�[5�V��F��9H��dn�!�sl�1��\���2�#��es��7%nȲ�Zp����]f��9��m�t`�l�&�.	w;v�܂��t�Y9��]�4�"��8�2��������rwP{r��6�k@Z;;��ڷ�q�
�R��l�i3=�s���5tL:��7�����Us0�d0�ۚ�0�/<��X��,uˈ��n�R��B��[����=��V�F!�v]�<x {�ܤ������a:�>|'|���n��3����n��o%�$��&E˙r7
dp��㮰D;b��og����,F�l^�� ���Y�b�g�x���:�)Ű��:S��.Fz9��i�n�ڑ��ns����J��%ƃ�Q���Qf�XF���C6�&�z�.�l�hE��Pi��ٽm=�n9�����ү(��2]��ɦ����-�{��w.F��瓦��Sm�b�cl؁�&F�j�ͬ��!F�.�G�o�!�r�H�{�b̼�k��s��o	�W���x�����T�2�֡H���
D!z�f��WC�pPG[�Yb�;jV�a�
�I\ѣ�8��e���o!���Ǎ�w)p��P�k��[U� �,ˌ�ٴ�05F
gv�f���H��/7Q��C/Pm�7R5Y���c�i5fѰ]�8\O	3��k�[���;5.a��vQ�Ypc��T��-�|��w{��{�;�{��'-�ն:N�ck�x3X��g��cr���p�5�v	���j��b5.�T�F',����ip�)�l]j��m4^Ք�k���6MŸ��:��x�=��F.]-Z�#5jh�L��^�\�IE.��j�s����a���A��՛��/*���n�	�t�n9����waE؎��{V��5�A�k3��c����?�r�bm�Z�b��m"��\�ݗUɛօh�%�KDl��j}��$}}^݌i��t��U�*aCIߥ�
�.*d1��a7��	ڕ���9eǉC9�^��g���,��njw�wK���G����� �}�hQ̓�{}�Т=c��'���)�����aJ���e�7��+��u<7/�n���4-ȟ����r��}�����Wv��|����k�h�ld��B��JG� @�L<	�n?���ߥD(m=���S^���Ad�2�g�����X�t�g/Y���AH)9��>�R��i4 S*�[%$���`i����2�i&��U,�o�W���ϼw���A@��"sdG�X���wM^���U�f�DxXfP~I!ET�)��I3�`i �c%0̨ZII
�2�H,5�s��k~���������Dsn��*[6�Rl��z��m��m���GI[]�zH)�{�4�R�T-�RA`T�ڐX4�S3,��#�� %G�"�{��3��6�~��R
AC�������{��ٿ�N'{���II�N��I&����KI�Rfe��ƒ�GI �2�H-�) �-a9�����}J�PB\*�ϓu���/x^��7�y+s"�dU�GVejx��d]�Veڽ
��r\k�ą��־�IH]��?�%0�j����Xʥ ���~���~絮~ӕ���w�
AM{�I���a��ZAH,�Ԃ�R
fe���U̮?~����؇�����)�꥖�I
II�e��6��ʅ��B�T�X�H)32�(�ͷ��記���y�gj�}�U����}��H,3(?�
B��j����
T3��6�Y�Ja�P�4$���A�])���S3,6m �p�ƻ�|������?vq�ڨZbRA`n�H) ��~�4�<	�J<$�BLV��螯��Y���`]R�ђ�
AOs��
Aa��9��9�ې����*�K����S��L��XfPi�AH,�Rq�I+34�62Sʅ�^�s_��s=�䂇��<	�|�������M�_x<	���'��=P�%$z�H) �fX�
Aiʆ��$JO�|h�;s��18�&��!u���W꺥s�b�1e�'���\�kn9����K<��P�%&�v��AH,6s�$��S*�Ke$�$$�G�]k�}�7��?Rs~�<	�J �#�����/ng_UtC��1�� ��
H)G���Af�Ja��-	) �C�R�) �fXm�Je0̨Z������`󯞩���AM}�f肐ZC�P�AMwO9������[w���0.�gᒒ
$��=`i�) ����Ri
`eR��bY.4ȼ�ԟ��@D���H,=�:H)
*�eR�[`RAL̰4�Y��L3*����P��])�}���v˫/���+�<�eQڻ��fnէ{��g��~�g629�6�C5� CW��z�F���=n�uNj�R�5H�6�s�;�{�����gsU;���N�x<	� ~6�R�B�
A`y�����AL̰77D���$�@�4�d���u�W9��~�m~�<���I ��~�i ��B��d���P))32������~��>��|�-���Aa�A��
B��i ���!����j�޷�ހ�@�F@*0s�i��Ka!
Ns��{��g��o�XAH/"\xQ����}�O}g2��]� ��-���P�����HlII�{�$��ƒ
AH)���O�7�����W����A��\�����`�ԦZ�����%��yU�D6�-�����ݷ��$�T4�[�R����ld��CPII
a�<	�����?�F�eD&ӯ�	��> Y��r>����>�����xI �%$�H,i �s��肐Z̨i ��)��2�%$(II����JH,5�~����]�����Y�q �؅06�%��
@H�} 
>�Z�}������)9�Q�e��AHT��֒c�
Q����͌��2�hf����5�e����$0a����S����H,��a��@�%$4�X�AL̰4�R�3*OEM���g��Ut���D�g2�r���?��R
{��4��RAaG�p�AI�)��2X�H(���`i��4�XfPht�R9��?i����i �`RAJ���H,�d�ꅡ���
0��|'���_|�7�*����H�$Wd��Ci��S�B�5��=�~�����M�fk���W�#VX�3<g�<��sٕ+4�Ʊ6bwv?%+y0۝����������9&���9U���Y�^꿒B=��Xƒ
{�4�R�v����@�U,�JH(RJL̰4�ReB�
A`eR�[s������yO��$��#�� Q�>���NN}�>9����H,9��$�P;T���R��h���2�hr$���2�H,(�u�~�{��w���^!y��ⴥ�p�u�Yn�r�!m���M��F��Sm�H)_�a�H,��a��@�RA`~�Rƒ
fe��� ��eCI5+?q�߽W��y��ϲ��05T���I�~��,��0�O׫HlII�O�\4�Ri
`eR�c) ���L��XfPh$�P2�H-�$�v�m���{}���L=څ��%$)�])��������Y\�}�_{���������Ad���ݨZ���]��m$�����k���=�t��]!�T4�S@�LU) �q%'��Hm%$�H)��K&�I�A	) Q��/���A��rq�?as�����AH,�)�$�������Ja�P���P��R�
H)���m �k��_t~�������{ꅠxJH,
2�H,i �?v��肐Z	G��H+��|y��vr�d� 8��R
AC�������Xs��������bAI�
`}T�X�H(��~�4���Aa�P����U*����
Vfh�m��fT-��9�Ώ������
�L<	𑶟j��w�)m�����H׾��m ��B�5���Ԃ���AL̰77D�Ѐ�xQ��_��F_ٱ�2��F_�W4��<��9=;U���8�}7������\����ڽZ���+���+U�*���t2���˞t���������#�[��"6��~&��Y�R��8p�SqE��� ㍎�������۷b���9��l�ИL�z�pD�x���s���ۖ2��Դ�����n�9� ��ǔ�7]86����#YG`tpX�ų"��anՋo���]f!�"^a ]���"�wa�ظ�%T��
�u ���]�f�ƎSR��A�f3\Qu`Ͽ����Yh�f�Z�j���+�`;:�{j9�� O/L�SG<r�����܆��=��w�`����>�4�R�B�
NS*���P,JL̰4�ٞ�����y_b��!;�I�j�>4G�#�㯺o��R�$����6�Rv�hr	) �L2�H,.0����a���%FSʅ�i) �>�Ϸ�?��������R�I5��7D���T- ����~������^���Z��U) ��y`i�) ����I&�)��K'���Ng~Z�8�P>�����AH,>�A�I �;T���
Vfh�m��fT- �	��S�|V�ˈ�_F���ߧX��/;�����߬?m ��B�4��X� �-����`nn�)�ʆ�
A`eRͲRAB�߹_�Z��ַޒ�_�XC�%$?e�I&�)��K%���BJ@|��|��O�c�!;�$xXfP~$�P;T���$}Z�D���D�W:�p�O���|{�B�В�
��ҐXX
fe��6�Y)��2�i �)L�<	�BJ@�߾��n�2��)�C��$}�?��{���^�����<���gᒒ
����Hm%$�B�
A`eRɶRA@����L
�?�������ճ����l.t"̹�jh(���c&Zm��rJF�Z�	b�Z��K��XwuH)*�~�R
AH)y��i�d��CI) �2�H,=���r�~���a���w�)5�XH,����N��{��a�*��JH,
9v���S�큤��]�fT4�R*�ld���$���I �{�o�G�|6+"��G�wqd`��w��y��uUϺx�K�X�R����L����,e`[�����[I�Z���eI���_�W���� f��Ă�X�Y?���� ��H��ޯ�������;!	����Β
B��eR�[��
Q���Af�)�eB�}�߾5_���:JH(l]ҐXX
}������L��P�%$eڐX4�S3,��
Ah@�xQ��b���F���>s�6ks>�~���~d���$�����AH,6{.H)4�02�H)Ĥ��L�$�H)|���r�z�~���JA}�R��4�62S~�ZII
a�JAas���ٗ��?~3��{��R
k~�4�Rv�i �>ݜ�8��7���u��yH) ��偤��^{�$�02�e�%$���`i����2�i �A>�ֻ��h���?m���G� "�� Q�*A�y-��Rwz��'�T�:H)
���JAm�I+9���͌��2�i ���])�:�~cTu��� �Q5f�DL�mi�c0�iuF�1�/&�V3\fv��������t	���bH)��T-II�GnԂ�R
fe���RHs*#��B]"�~Z�M| ��2 �|d���������{��k��4�Ĕ�XW�i �U,�I����L��XfPj:H)��JAH)5߾�e����@�Ag̔Ü�ZAH(i�������?g9�_�c��f7��~� ����m �P�a��-BRA`Q� ����`x�~ϯ�w}��_D?j�����0>�R
AB�R}����II��$��U,��H(���`i���y���kR���>��TJ��ߧ�)nG^�呕cs��;�^�XR��F�/�� �o���W���}�Ì��!��7�|{�Ȍ�����xxx<�9����
N��#��fP$�U@ʥ �0) �L�t�62Sʅ����*���R
fe����%_=מ����7�k�l;u@�JH,�JA`[I9̰7� ���$s��~̯W���2�׀�꥟�) �I)=�XH)���gm���~����6���u �*���R
}��4��I�e�$�U@ʥ �������i�)�eB����_w���V��AB�v�H,3��y������i��G�"���@�<��ݨZ���v���S3,$��!�P�AJ�������M>�]KT4fV�Ś�LطS&�*�hŹt�DkZ�g�u��g~�I�Нtv$��}`i����p�AI�)��K%�RA@����L�w���M���~�Rw~�<	�J<$�G��>�\3�V���d����R
k�٠6�R�B����*���R
fe��H,��a�P���X����v�����I5���ReB�
j���_����_s2���<���gᒒ
AOw���JH,+��i ���ʥ��{?o��H(D���`i���Aa�Pj:H)�ڥ ������`i �c%0̨ZII
a�JA>?e��輵w��k�:�Zo>�R
k~��!���@�a��-II�^�Rƒ
fe����]��$��ʥ�) ���w�q�����~&�����?$���9P���B��R�R
�I�� ��,/��U���o�Pw>�<	�J��AHQU*����
~�~˼r)�ذ�Niͯ�c��!j���p�����?NknI�_\��X����q�7�kxu��B�X<�֕�������]C�֧X��2"2f̅R~������Ja��CBJH(S�JAH)32��Ad���2�hJH,
˵ �,H)����>���F��?w^ ���CI5+���?����ٙ_o�`}T��%$)%'��HlII�s�$�B�T�X�H(�3,0>������?����նldBĦ�y�s���Q�75G@]��ˌ���Y������������ݤ������R�R
AOw,$��2�i ���])���<__�#_i�.�y��#��Y��#������W������Z�RA`eR�X�AO����� �̨i ��02�e�RAB�Rfe��6���~�k�o��$�B��R
A@����X`l�w߫;�_}Ͽ|��e<����ä��XT���R���H)�eB�p���yۻ��ߏ��ׯ��A`~�R
AH)�}a��Je0������ʥ ����`|n�)0	G��H}�F掊x5���z5V��̯���U,�2RAB�R{��4�Ĕ�XQ�\4�RhB�T�\e$���`i�����2�N�
C�sV���Ͽg`UR�R
AL>��������~ʅ��%$��L<	�}<�}_|�g�\�m������?m �P�a��-II�_�Y��[�m�ީ ��ް>7D���CI5)��K-��
AL̰4�Ĕ�XfT- �U,��+_�Z����׾zu H�EvH���֚��y�����H,3(?:H)
���JAH),�w@mc�W�}��ާo�o:ibp����y��h"f�����k�ɭ�*�.0�4r��>���or�T�������{wcwu^��ռ�;�% h�[��}�f}���y���d�ݚ,s�%MŨi�k�(�͂D�!ƚ㉑���6:�i�R{��:�St��M���(`8�t<�]����x��fS�=.-�-N�wT�[[jԌ/Z\�����e�z���u�ں�eb� �\s<�^�H`Cjl�uW1���q����L΋��C���ڎ���7&W���k�T�o<�]�����p\��ƥ��B��Y���:�)#
�T�YrkI�±h��j�������q� �ݯW�ݑ>/������Ԭ�dp#*��mM�{,���DA�٠F�� ��:��OF]��row���|�-�F����M碟^�A�?e����ٲ�-˿]�����S>�"|t� ����[�I��>�4��5��^�e���,Yi��
>#���J��lz�ڡ�����	/�0A= ��>��"|y�����-m�W���-�Д�ʽ��z�d|��}��	�QoAwhPv;��OH�'c�22�Z��o"�]7��r8��q�#wj��j���~�ʀ�~���YxK�� �esaC4�8m(#�H�^86]&������F��ߕ�@�7��E|�κ��ު���E�:,����4�ސv��X���2��`�kx0Z~2���^3n~/o�M���'d��2��Sur%�щv>љES�r�[Aۗ/T�q�6;^�T�eV�S���`�r�d`}��o��/k����� ���x��7�+�T��Y?�Y��^; p-���9��WV�ń��VL_x|p`��JGȅW뎭}�����U����Zq:��S�,� ����j'9e�CY\߹���k�w�F�,Yݚ��R��YR8 �F�O�����Y8��u���(�Ϡ�ݑ^;�$i�7w8�yB�����n���AY�)^�#� �sDr'�Hwvi�|'�G�c��OY�:-b��c2�C�me�8��y&�[��(��,R�Q��ߟ�}:����#c��R}|�'�Z�E>����oo٤�KN�0g��{�_;V'�P�	�yv֥�hӉB1�2�y]��j���Y#s��i�մ(��d尧*��6= �ܟoG�lz�����+FVT�9zi]N����̦�C)�X&�d;�ڶ\�S.&�H�WVa)qR�(,��R�u.]�QcC!�0���B�b6���3x��s7��R����g���3F�_bҮNد���O������Q*�k���G�{�Ǒ''\��P���xg�.�������*�')⬐iӑ�ҧL�=J�|�oB� ��fNe`�9�Bm³6d]��M��NB֨�.S�2Vד`�غ�{*�t6�d�Ľ��q��b�V�w�˦����m���:;w�oyZK��oʘE�=G��D�ӻ��5W�����f���o��j4fm7����r�wQ!�	�1�T�1{82"����ڭnM��1����bQf��]�ؽ�\�n�>��q��*��E:�<o	�7�u�K���nz�=�y+z^9��:�:v�}��ƳWn�d�8D�x�_�͘{��+���4�ة����c^�l�l�����S�o��8[읾���w&]C��]��f�� x�sۗ�&�3)��Qg��O@��/�����Z��83L{B��E�SU�5�C|�L
���B��7�i�繶+�W>۔�V�Q�w{�Ç
.&�:.�:�Wý̔�*eG�+��|v.�Ш��ٜ����ta�
�=�|���k�Y�U�6��Y	��F`���aR��7E���#_OVt:3%�с�F� �sq�Iأ7J�������*E����7֢^�g��1�{w���ڂ:ؤ����h*�Я������;9�Y[n����2ٌ�&ݶk[i��rm�*�K�9��Cj�ͳ��nɳ�gdȱ�2ՙ�j�ٽ�ymjV�����7q��Z`ein�2��M���v�n��imjkGrY���s�9�E�K���lX��e"h���ՇBP��[n7�i�ڛۢΊmF�;+jv�e�k-���MͶ-�r0�j�	٧cY��4X�i[j�M�"�)�۳���=�N^g#�"x��ۚ��$�9K[p���f
fY���5�2�M1�l�:
fI���"�;�n�Y�kY�b-�m���i�Nm3eq\U��n%j͓H��#�=��#Kem�M��&�Zf��ׯ{���!�:�oi��#�A.����D���wf�F�p�h4��h8>���۱�������Nrq���S�P ��^-���#7j�VȐt� ��׈>ݑ'H�oi��n(>�"����u��yη�e��g�s�K�*"s�ѡ�*�lz^&����B�A�:`b*f�ƀKh�3��f̓5�u.x��E�G]��Oqq_��mD��z�گ�"|
犸&OZ��ŘGx��%Ȍ#�u�x��C���@|wvh�"A:|;�b��:ӆ�@�G���\�}|��v����|(^���z�b�>ٔ�*�';��3�"�橢ݟiAwg�rQK�ͭ���0�H܏a���۱��=��n�P��r��H��vuW��+�*�\��׋0� ���Ϡ��O&��� ��=3�yM�x<�$=QL�t&�ު�*�*qz�Uc�V�̗���d�ge�0�Uo��6�������w�t|  x]稁�{�@�ِA�� �ݡ^;���W�K>T;���9_6�NҖ��O��=������xfZ���	�|�5$Y���$4��t�h&6���r9��C7��D,����\c���A�sD=�i��٭���Nn���<Y#s�����)ZP��h�t(�|0}O�[_�����	����%���x��b�%s�\�DpŭμY�-�� � �(�CV�!���Dk���n�;��ދѐ&�cO���ONҗ����S��C*P��559ʜMD������e�$I� A�ٯm7�����G�$np�N��Șvg.������춯�7
~�l�V=;4�$��[�c����^,�;���)��ݞeI"oP"��b+v��rb�p��K6HQZ��{��l�#�LSՀ\���-��w����q�J�ee@f%�',����?{��	��D�j0)��4��U�� �mW��*��dE�
[L�)+5������j�0t��d�ֶU'�4s��gH�jg�烜!�"�M�.���*�0���vA;b��.w��-.���F
�j�b��B��]����H�݌np��e�Ϸ-�,�
���n�q���ք{�9��l9L)3�8��]j�Bi���Vn����O�]��p��#c���r��9��9ѭ�,�v��(5�=[�����7�n����ؒ�=��������eK[�ޠ���ִo(آ�z "�׫�nȐ�(s��4��ev�q�R.w/[M��qu������$t�G�
v7+��~�0�9�����A�>�n�LOC�q6v��bze�[�μY�q�w4#�:D�ݚ��$\3U�m�>�BW>݌�GG7���nFʗ��#�{����Ɯ︌ίW����^>�����
�AM�<).��mN�K���Q�����w���֘0S�c�-�����-<R	��biK�P��YEm�0���s���~o���b��!@���:=n��v ~��y���ӝZ��D���}Evc��΂���9˜�,G��4��Y�����h�_�T=�/<���kަ��9y�rRA��Jzn�Lj�V*{��bB��f�ˊ9��< ����>�=.=���_���ل�}��� Txn웹V7�C�lL�� @/\����0j�!�[Y����^�ӷߥF�*a������@#qH��#c��7v�C}�Wp�e���i���m���/V�G%�Ūsw,� �h�5z����L>�2�� �{\�����@n�;�x�䇡�G�)8�pw]�iT�}�������^݁�R����]Y����g�oM<K&ZW)�A�pR����ˑ��LX���<�/�w���VO�zD���wf��i�ӑ�Ą�1�#n�j�Ö���'#c����0cb���Èp�������)r�f9��i�In��}X�O�Ӄ��p.��C����Ω`�G�mY�v$���"��v&�P��s���"i5���^�כ�ܸq�h�'����R�IC��y���d�i�]�;'�x#�����^6��x�K��S���H!G����"N�)R{}F�	N�N���"��^�[�+����ّ��:|*6ŇŨ֡)���L�C(�-�� ���)���nvj����{*�V��3��V4�-[�q�hqO��GweE���<R;X�glk����V�1�l��ņ�ˌͅ�0hX���k\Y]��١ǳ�=���ǿwBc�K����.�T��E9	�R33�=]+z�|#�(O��5�Y`�)���>ŗg�������W)��kE_���ӗg7�����,��U}ָ<e��g±�`��Ǡ�ݟn��&Y�!H�]k7��j��+R�#�%��P�"|� ����#�Vp˼.��'�E�$��'guR�oT�{��}_{�����x*;пߙo��
��Nu�����Ң�� P+*�ov�-�f��t���?OڋŃ��34h�kjʕxq�{~�}�git�ѯ�y�H���39�����<J�9�\��,��9���5�}A����7�����v1�6dnw�G��,���Pv��:d3=�=�k�PPŤ� g8Z�qL��7L�R����kA�v�ĕ�e_'��aǟ.�'�׉�߷��!L-���2��NV%�GTVK�i=�Y���F���P��	�\���}r��炔U��CA�Ǡ(l����ީR�}�P>-D�Q�n�r�[W�}Ả,�6��#v}�P �wvK����7�tn��ccfF�H'O��B��{O���)�E�}y��!�AQ�w:��aogwD�w�9X��A-����O��A��7W��;���e�������/�z抎��
)��Q���k�/w�NG�AG��Ϸ`,��یl�fr��z�v8t>�<�p�^�>p�����,����[�uzi�����D=� -7���C���;JDj
Qi�9�<?���O���q*��vui���J��pz6��6ݹ�8U�Cz�t��Ϛ�[a�����<d��+���qT"�vi�YY��]�Ρ(��Xv���2���}$/]��e�nx�K��[�j�3s�p��^xcD���ls��P�1�c;g��	\UИ
m�7hE��v��A��g���8�J9��Ӆ6jH[f���������g�9�3��[p�����!�eGdr���V�g �lG���	�B���{"N� ������G3���g6dnt��'�U^}"�w�H;���^݉#c*��Mj�s����[���e;Ɯ�%�@�[ɠ�|t�[Ww3�������~����`��bR�Q�p�f����:�\v���V�N�H�r8�IG��ݟn�ä	tz���P�!��J#2<��;�5������b�1�"��'�}s��f�L�X��q>!A��i_O�e��W���&��w��9��n��e;���%�G A-��:���bڠ�?�����%��M5��9�+o�ep�n��'��b�1q(�K��"R�h˅����ǫ���T�sS���NT���o����[��4��N�ͬȈ� �2�J�Ϲ�j3��ǉPE�9z��՟���.��ɀ�U�E5��͝:n4DFMx�*n��os>�&���P~<��b:n�0��t�֠hVl�o/R�#!7*�P��{����{ǈ�A?j��߸���b���"�x��7��݇��J�=�w ���	�b�tzFǠ���ݑĭ���98�����n�:�����/s����ǈP�D�&BݞvTݟ/|��wG�l{�:�>-sqN�{"i�
q�tޥ5+1GJܗ�v泖\x���r��r�ޤ�S;�l#ݳY{�s�;�N�s'fE�ؾ��0Y������Y�����G��OQ��&�F-�Ne�ZlC4�K�%�����q�妲9�37��!����$�����ޚeO�0�ެ�oV��5(�{<cB�s���3�:��s���r�q�35�-��V.��[� �}�u����Ne�{bi�[���=n�g��׏��s�~>U�b�Q����~���� �ѩ�?RH���� �^�ם�|��:��B2��;;����\���h�=:���RZ�hJ�)w�<Hٸ׎��?���3{�ݕ8䝌�N̍���<eDN}���|#ʔ'9˚��z}�q��G��
��
{q>��ڋoVQ �h�$j��ԫ�("�y��F�� >������"��2��q�鬸棗"���lM>	N$@Q�[u�i��������ܿ�4�&�ac���+�����4�X�f�E.68�vh(�ю��</�|ܲ�'H�A��ٯV4�:s�0v3�;2/xH/6w��dj�2)l��`G�[^?�(f�-\#s���~/�x��ҩ���W/�#��sD�D�t��sW�7�A���v	�O��n�
;�$��㽻�'9l%�L6�퉧)Đ���ݪ��'�H� Wj��fK��pkr}�$IDA�wfq&9+�ڃ����"���O����ckxR�Slb��u*�_X�-˸XA��ls��3W�}0*�M� p댜˜��Vl�]J
8R�7��������v����_~����Bs�քyʒ6=n�t��F=���z�w���w��m��G|]��=�>:@���6.���z�|/�s�4�u���X䵗jጦ���6�;Z�K�Qa`��lնgu��hq��C�ϯ{�}�ڧ��wK\1T���lM��Unf�;�*����3)������V,a�`;�5�/���3��|q���Akf�g&9��ڍ��d�H͏a�}��Pv2��zzϥT���օ��9R���Dݑ`��
�t���o6[��sm��8;sD�D�"  ���@��sk�a箔�N�P;�$�GK��-pͩ���؛s�Q�a;�1��W�C�O�<�
0�>���0Z���f���7`�ܦ{�qJ붶c!�v�f�t�#qW�c���4���%���q���g�s�hts�_����e"���ڧ7�{�4�b�T��
nM����Ɍ��z�?bi3�4�+�z��gZY�t��ٱ#L��5}^p�V�>�/Q������FJW,�koc]Xɖ[y�؛�9eUу�i�PŮ��	 �OH�e^9�����ͻ��}g=�%�Em �g���C)����G��pUjS��i��=��ӧw��W���å��Mؽc2��3�g!ku�<91V�Q0MR)R�nˊ�����z�<E��}�9h�r"����n-��Uy��r!Û��$�g�J<��f��Z��ې�; ���ԁ��~�˷��;+ؓ��ی"�6&�i������&Z�8�%l�3|�����[���:4L�	��x3o]Ş9.�����a���2�Ƿ�x������I��G&�y'�*�N���5����)�mmeϕؼ�������;���C��<f�a;R����&	�2��X�A�V��ɲ.P�g��FWl�k���o�}�z&���9/�������5w�۽�0�;BI-��/Rx5&ܧ^�O��9�^Zr����liǓ��L,��e��Il�³{:4��5z�k���G*<����P�2��yW/�5�2s��&��M�N�>���=��c]�G�ד�^�G_W3z���=�%5��_��G����n�}��m��)�q����Y�����������]�9�|��z�Ӹ�Xdu��H�剱�uM�A]����MwL�1 $�ml�'���&��q���[n�P#�E�gJ�$�ݖSZ�r:&�9O���m�t�݅c4��%#���ܜ!���Z��J[;6��2��֚ݣ��v3���3���ݳ;N:2�f�IͰ�mͬ%�m�����Z��P���e�u�X����[kZ��i�KfЧ6�7n�6�)i��m��kKlm��$٬��Z8J �gg9�[am�!�9���te�AFu�H�֛����36cd�$�Ŷ�c-e�S4ss��彌��l�,۶Ւ;mֳ��#�mee�ܥ��H�$�;ktٚ	m���kv�;;$jM��3ޭz�dDز��mh2���Ӻl�ٍ��m��8�Fl�vI�E��,��u�MkjKl[)C��I�������֦^�<u�P^6��,yݎ�]�v�.C;h�9'�7�٩�M�f��-^J�D�bT#M�K���kV�g�g`E�W-A�	�h�甐�c�f�G�1�ˁ[K��N����p��b㓫�n[bSiR�nm�a�5i5�c CL�K�<.niXt�yՆk�b��h71�;%4���&����8�6�g�x�kiA�j�b�n���,�� ��6:����8j��>�x�7���2rv,�Ѝ6��i�g��"��� `�F9�-�j�Q뵱�,2b���xmy����!u֡���nX��n��E�h��y�q5�`8燯2�e�PO2��뭸�:��;Y�����06����7[e�N��2(Pm�8��M{d�.����J���ƃ��_NVaG�����X�3�DĆ2�wT3lK,�2i��
m����i��f"]h7����K��`�e��ˆ�sύ�+�'v�k�����-�p��p==�w^-˚8�����)�+!��2؂Fc�����c�����h|�]R�F;�c��;��JB�й���\/cnɷ.;mR�r�ܯPM��m,J� .��$�5��ʌ1��һ�#/l[��y�%�=�kT�]��α���	��W6ϳ�qy���lY�ۓ:�G�T!m���<�u��T�c2�"�c6�7p��ۑ���lڞ����y"9��P�p����+˞��R���x݆u�pg	��td���}��y1D;u�(����\9n���e��Ai	voh�	��j���fŔ(���\b�e��<�w�u1��1���0��V��dΞ� a���l�͵ۮ�-�L��ɺ�ۣ[pv����-��-ڜ�JL�[���,t{-��j,�[ی7�nP�R�.f�*�r��S1�3�Й��aakfAR5�3����]eY�.a�̹tˊd&���h�m�l���Z�qh���"3�n���_�{��=/�=�;v�'\�l=l=3�s̳e�c�2�6Ɣ�rZ\�iB�kV
��`\ղĕ�����/SZ�X�SFkZ���@s�)K\�i˃B3R�L\E֣^Z�j9�ې�9:�C��㓓��\m������g�Rq�nc�s���\�^8�݆�Ы1b�2�1�ivsy�{U�Ay_.��Qfk�¶ک��������� �5 �� \��n�tG:��Z1#� �]���4B`���׃��~\~?�����VH
Uc��,����W$�7�9PRD�ֵ��'>������9˱#�QXg��U|,���/�AǠt�[���ژz�튷�	N'����څE�;�N�����%�r�#9�-��vi��퓙�x���n���ls'jFlO���P;�$i���9k��@���8�x�Ϊ�ݑ.UcI�YE�Ҋm\����y̪�������|Ӛ�#vD�O�}��(��T�:��'�Ǻ*M��U0�9�o��Ă
�@�kVW[��I���i0� �\:���K������Ŋ1��]���)�BẌ́֗�'�0}IMx�� A�ٜk�T����l6J��$>,6��[r�Ο	�t(� �>�7v�@��Ve7y�ћ�iBB� �����/��X6|Z��M�-���00�Ut��RTd\�uӗ\�ة��]!�=��yr>����FwO���*���e{J)5pG|U��^Ȑt�B6�ЁW�@����>���; )��Ooa��\��R^';b�ϵGx���wo�����{�*35�tgV��}�|Ȣ	�ٜ��T����k�T��A����"��=��OZ�}#8z9ʸ"z��sf��*��)9�|ov$mW��dK�X�|Qw��W�iO^Ȑt� �������V��E���6���fk�]��E}�����6�ۮ�,<��&SI������3��^g{��3�<Nv�[�^�����ײ�<�=f�����(ݚ*�9�E��r*���	��R�����ͨޟ�d��`|F��֗�O/>��ٟT/�١~�Z'*P��.js�&�/#���O����[_m�ɶ�k&�;`/�|1l�����YĜ}����1LMf�ҰR�	r��E6�F�\e��V���a��Km%x
�|���]�8����nh��t� ����ܐ�'P�ɍ��13gȄ�|�g�#cЦX�=ϙɄk��V��	N$'��-*�K(�3~�7��x���H��ݚ�t���l��a�F�͵o���ݨ�.
��q��n)wc��_h<��S�o���ȸ�h���`TC�E0D��Ju���Bn��`9���{����;�w�n������>�X־(��qI��8���jVs�w/>KF�ba���m_[�|FNlS{haj'����Gww8��k��V�p)Ǥ(�7w8ml�8)�"}�~X��t��0Z�
0�j��v�r!�-��5ٻ���U#����B�wc�6=n�
�s]�ݻsq�*<7:�^;�:!=Z�+��i�6�H�	V�i�R�(Ѐk�)�ͦ�M�����D��!�tӔ��A8���v���n��K--f��jT'�V����<��!���q)�r���ؼe�ݯn�}���{fQ��H��D�7[�0��s�*�
��AQ�n�
�V���z�݃��e��a`lKX�ܵ�γYutj]�Fg hc� jxy�L�%�MF���D��-u�F��vc\�*�-�����>�͡@�A���e��<Ҿ��F��n{�����)�O��.��Sj���x��D�#2;G]e��F��	ȐA��wk۱� ��F�p9�i�P�/j*a��lU��Q��F���7dO��M����M7�^ �"K"���y�x���[����m�[���A��
���ң�����Ilz<F��]jt�*�D����>
�Ūp�;�����?��g�R���4v�oME�v�b��C��Y������oE�R��ú������/�����8�q6��=���Ul��y?{�K�.<Bi�����Q�z`l�����-�jfVݮY�1K	i���d�ۍM����at<��^yM�z�D�����|�ݴ��o2Q(��ڷ/K�����e4�`K�.�Q��=͌`�����շdDV��tsk��Gm�j0��jAS\F��2B�M��M�}�R���nըR۔�JW�Ϥ.��]�'�nNݕ�ۦrR}����O�in!�z��j��r�f�l�e�S82&�lYl�sl+f��j���X�2�9�Y��*��G+�^���1P��s�*�z����uj=�q��q��f��֜X(Ã�jx3Ɠ�,�cF�"<A%49�|�nmd>�p��>��^;�il4�H��G��ʠA���ݱ^;�0{��&._�;�I1�J2R�[vC��A�O� �d+�,Y����)Y�-}pf���'��莖�}���Bg5�X����q'��WYrf��Q��/6�x�r$" >�٠A��:FP��<�����5���S�{�q�ڀ�H>:| j��I��`y����|-��7�K4x&lt��Y��֞؞h뫷R��k�,H�n}�n�|�B>�F�ϫ۲$*����Z�����Wdw�=�N;wr�͐CR$@�wvh�A��ou]�h<{��Rz*H&0ъy���5Ajw+�6��<z���N�ͫ�0�s��ř������(\ճZjq�����H|^Ǥtz=y���b�3��,S��Q��z<F��R9�Nz��p0"��ݑ'H����]�fn8v)U�7Ykp�tbt�w��a��<��?�[^<K�E-d�L��S�Q�nl��dt�����X򶓜J�� �nhF��lF�qe�k+X���Q��ށ9�,xʈ�ѧ������b}���t�%�>F)K��Yb��q$�F�Ϩ�)�?��ﯡ������;�9됇R�+E&�����i���\<]+מ�u�ѭ��������ߧ�"���x;v�q��[�����	@���wo�AqT}�_9
Q�>���|wbA
DFH�OMk>���@ND��[͞�)9Ī���v��Hє��]�������o�,G���sB�݉��>�*vWN�f�k�}R�鍻ҍ�c%M�_r�l��r�qn��B��_WDΞ��֠lx	�f5ê
3Kv�ʹs�3�\���)�9���[�%��#wk����t���hc�9v�g2"��@�p$"�vivZ}���M�5���:|.�hۥ%Lq��;��ą`����<Ұ`��2� �lj��j�z�ut�y�U�')<����K�4A�9��@�wvz�v�w
��Yϐ\Xݸ4a�N�m��谎�A��=���e�'i���)���纼bҾ,x�;;�xE7G��V����
�ɭ����|0g�[�ᖬB���j�Ӗ$�W�S#A���<��A�q��V�j��;��x��!��>�\b3B��c�A͉ �c�wg�����N�ۅ(��MF;��y)U����C�t� ���@�ّ�f�u>ǁS'��{�`#O���.{���n�%yb��
q$].�9z_Vȋ]�c-U��Pi)�T�r8����N%��!��;��[�s�nD�T]O[}�YF3!<%�ZZ'(㌑�n �2VM�hM_9<%��MFs.q<�/H���&d�;�d w�kZ��=��n9����}��xŧ�>� �W���i0��v;%�Yl&��-"-�v�!?�<��O,��MkEQz5��c��pG�JNs�5r�?{M[M�w3z�R� gDs����Z����% ���v���pC7�kV>�A䠼uD��=ݢ��>F)�8�劷)Ă�xn��Iӫ�7~��>�(�m��dI� n��y�NiG;��o7u����*���@ ��zv<7vA�s�T���#H*=n*���T^�o�k����J�� ��h��Ti� 9�4ݟO����mxŧd3���Ä�s���'��<��^X�r8�G�F�Яn��FQ�y�sY�e��⛹͈sm6�,�d1�V���c���&C�Xxtz�air�♜Q�lc�95�`f/Jt�,�V͹�v��7���Ph4�,$C��7�뱅��7gq:�E��iY�G��iI��^sKeC �4�9�l�2�5B�A�h�m�/"ɮ%��3R�hU��;A*�:�K6��vv�X��Q�$���q���X�I<�y̢��3�x�q�+>�n��(����h)6�*	0V�%�4�K��1���!�i���K�"��u�U"��۪��k��8����}љ��I�B�Θtm�3�]�bU�G�a��-P�k��K���� md��H��@ �ݞ�k;�w�6�*���;�[]����A��^/��}^"ڱ�J��Z]��{����y��ޑ/�7��1����VGAv��:B�5'{�4`5�4��>�;�B�݉ � ���17VjÆ�2��Y�k,U��AN$�z�>���G;�/Oy�:�^�����c ���c\�G^�ێUe} �p�r��/ެЏtIG���+�v$���#mz����b���췽��ږ�s���{�ބ{�,x���9˪��;]��������|e�q+�B�tE�ê�R��G6��bȖ�4dxu��z���}:_?1����|Whqo��N���Yb��}��u˛�ݛ�i�4�mϷc�F�N�ϑ|�z�*�b1C�\�,s�#������&�xW�*7�uo�-��g�7�����-�V�{yr����R�����NӇUc)D���A��sK�_.ի6�YC_	����Pv4�4-���y�z #�@��O�;�u��uXN�(��V����2sw%*�8�U��8�aφ��?�Zq��m��}�}D��7lx��ž�:�+me��#��*�UՈS��G+�+��'�H�;�5��dI�'1�VإP�s^䷻��X���U�5�@8}�X��0S�oPb���ߏD�$O�Y"Łc�X��a�0آ�%Е�-cYX\�x��]��u�����=�$#�n�W��c�]ݕ�9���Y�v���k3tZ�T�o�:�����Nr�`�w��b�ˬW�`:�H.=�C�}�
u�V��n}�<����0��
�'�$>���B�9�j�� M���9_��s���Ĉ����!��TR'5��T���H�{4��h�����#�p��n/u��{�qx�z���f�@�Giy|�׷v�Ӈ9K�[pP�/n�ۋx⶯z����G��wj��mE�X{8���^�����l�����)�]6�贘=��C�t�ܳ��yO/it/L��^D�IO����T�3|?w�K7|g�����ܻ�.p�� �eE�����	�M�q*��wp`V�7&սƸ]�d�0!�;�������^�q:\;h}��.��,���'z`ฅ~:ww^���U��$�3݆l�N`���:xy��g�]��)��Ɍ8��=�Y�)O��J�{&^��GY_��_k����^�3��ʋų,�
���z�v[2W�U��ңN!��E�ܙkw�Ly�y����k�:Mᾑ�K:��8�r�sJ��)��S;:ě�O�A���ҥ=�����x��N��l�{
ȡ,Y�1U��FB,Zļ�.-eb��m�#aʱ��F��ZC�2��L�x��i�g��4wPW/u�1n>;Ӣ��z0���{V�7�ڷ�I��<�G�]����dM%֫���{��z������#�L��A6�.��M�k��S�oRW������I��{�C�rmȀ�ܸ��"h�V{����V��o����3w
�&ӏ}T-{ǀ^�b�������2���1ա㛤deu������2���%�i�2m^e���E���Q�,[���}��*��=�����%T�&Z�ٻ[��&i��8���{���m�����:���m���8h������eZp�6���ն�����A6ʹ\r[V��٣�S��͉��y`%�m��m،Ӗ�i��)
hڰ�&i[�첁 m�k�ZktYΔ��Π��dr	��̡��ŻjK&n.m��{���f�b֭�$ێ�W�/I�-�볯,�L��۠��;ZԶ��iіF�3D�&ۤ��;�HM���"Nf��׽��Gy��,�mi�����6��9�d��M��@�Hm�S�"m�w���[�`�Β�[s`���$�q[d�f��P�k��/[,��e�2w!��!�ۉ�d��fw�����g6av�vp�NpPFڳ�e�,��gb8�m��":'m��T�����.�fڙ���������I�7�9,Ue|�����P;�> ��@#wj�#*L��+wb�A�� F�B�F��w�wvVl\��JUdqnh×U^&�X,��׈ݑ ���;�B��u�9ֆU%��Oh�����YEmڱv�p+�|Aq�#v�V,���Ɩ~�j�D<�% ��ݹK����Ój�R룄ڳ60sD�ODM�qȓ�Aݚ���^,]�Ue}"��y����`��(��B>	+�Jh�Sy}�A���o��>���W��o�s6nsw%*���!��8��KWkZ���\�e�e#33F�3/Q�>�5v��;����`�yEmڱv�P%>�� ��A	swr�8f6'�eyN����~�4�IP�D%47s�z�.�,Ue���O�:��)ŚY��v����Y�E���?j��8;/i��ƅ�<�{��Ӭe�{�wG�'|azS��Ħ�
$��@���Nn-)����E%4A
=$�l��#�dzkv�v&���f�7rR�#��>��
�C�;����e��u_�2q���0��WXF�f����X�¦&ҭfքh[f�J��I��1�v{�8} ��W�S�|�����p*��ݫV.�z�Hŵ���úv��"n�'s�534hJ\̹{�k�!���5^d2�.������^,]�X���G��AIТ��ᘤkV�GH�u(N{�h}�ޑ�Q32���|պ]��w0f>թ���Nn�V|)�R(@���$�PUD�.z>�AmР_t��zWh-��S�;�j���^O��
��q[�T���7]W��",�RS^�
(������&�hF���&����>��k��Yak�P ��|��E%4!G�êظ�N��0r�7�A�T�����^�~��n�\�Xk7�EV��s
9uڊ-�>v��=��~J5��o\����i��g�^����w�'sn}��KW[le�%[�S�ݰ�U�*��E��0�%u�[�-���"ŚZ#(p驭����þ/ga{n,8,���V�,7m��V6��	��pBL걥�Rv�ol�۝CI�$*��v�gq�s�-a]3�]��q����$5cU�J³6���4���I���b�ǩrT2�6��.4v:`u�u������6z�EU:�ػ�I�V��]D{mр,��׎�y����*h�	�X��n9�A���!%>���L^�}ϻ1m���JUdq�w��tE=�D�=�O��#����e�f��׷��N^P�]��x�9�
�zK}��a;��X�]����tx$�"��d��R�|ލG�H�s����48�s�RfUΔ�A�^sloV��e�������A	�RS^ �	+�	���Oj�c���,FG���W�IP�+w>�ŗS��)]�����dH�ڝ��g:ߴ����IUQ�IP���8n����u\�@�VKIw	SN#v�ط�@��h��BJ|���@F��<��>��}���1�Z�cvj��ݪ[�D���ER\s���1ɧO<r�F��ۻ}>7�>�t(@���	�wq}[��i�*��'�6�&�8}8�Aoc���6���H*=$��)�E�����+��R��PũǦ�n]�mUPŬ���w�ܜ"x'��Ё"�~�dA��m���	�a����y�ξ�S���]��|۠����n��fnJWdq��^kS�D��j7'8U3{P=�4G5T	��!%"�))�A
=>=����qm`���bTӈ[X�[��Nxz=$����E!�4��:�6i����^DX��	���{����*��7#��� �r��蒏N�r�@B�A	*�jS�|P�w�+]^.���fР,J�M�mڳY����A�k'ٮF�D))�墻�A�9q�0P4:���"�*�ؑ�upM�e	]��f,��9��� ,`�A�{��(Ϡuu
))���DV�ny>�����]�yޡ/s5���)s38A�G����x��
(���׈��ē"n�����kܵ>�=ks*X��_P'O�Bn� RS�����C�Θ� ��"��@����!G�J��$���o��Բ�º��]����1{�]�W�V�i����v���q~��;6��`�W6n��.����O���S�ԋ� �m!�K7��R��{6#B�Zz�r՚�ܔ����Y4A�t(� ��!%^��e߶�k>@��"��s^!@�Ԝ�O�����b�u���@�i=Jq�ٛ����u��	�
"��%B�DT�bC/)�E�M-m�:봫�R�N�z�W��7^IN�
�=�(N�ͽ�q ��
�є�tԆ�V2�Qkh:�X�T2�q���m���Uz��_a��פfT�33SQ�T+�'s_>��vk3rR�#�C�E';�31���3��x� �⒚!%U�|&�\�����ka��6�}AG�jO�e�
T�z�[�	���tz	(��6g�7L����m��^�&fh��9�t1�y�ۉ*Wi;p�������@ ��W�RS^ �G���B'�ܣo*Ng3�;�����F��IP�cs_>�vk36R�#�A��_�f�V^��=�J� �1g�a���e#%�-��_��f���i��j��'�츘�	�cGM����;4H�W��m۹�аY�IM���@�|S���/t���q�R�9җ\)�n��n���wMz=$���J�lွ��g.T���\�a�tstN�[����)��m3�-��3F�$�T:G|i9�sT+����M�>�����S���ʎ��x�/:E˦�!@!%"�IM-]wF4n��0x^5^��^�&���J� ��O�\��DzUx��Ws`x�Q �@��wv}@v`�4��a�y����K-�=T-�
�t�#����_>�x�p�	N�Xr '�:U�" -R�7�S�Z���;a����_(p��B��M��%t))�yG���,����:"2���wB�p��.���/�il�%ښ�f�
 AIL�;3w���=0S�sJ�]�ȚՒʧ*�+��cr�ɝ�o��Y~�V�A#��hk�����^�G���>���b�^�=�B@�$�&�V���ll�m��[t#$�+����w\�U8�� ��b���#����h��.GA;m�+���W�!�6m+��[2���!`����m�5�4��)�J١�ԫ�����L6�\D�;<0J����xå����b��*kI��a�����֭5�Y�%׍����ttU� ��&�X�5q\˜჆�G�Ŭf�����f-4�F���5J���Ū2�+@M֥�n�f�����w�z��{O��j��� �G�T�O�K�,�P�P�r!��tt���˚ �#�IW��$�W�"< �����ʫ6��9�GXgH�K]4;|���o��3���� �t(����ד�th����^��>Q�$�
�	*�L�Μ��Ϲᦎ^��ٲx�S^ �5РQA%>Ih�=a*��^���B�k�!EJI�u�e�bީ�@���DIӦPQ}~�D�O��@� |RS@�U�C��UQ�hɝ>s�v��zP��_
��St(���q�W|}����{/I��gJ`�-�L1�`�0)B�����@��ŕ�����n1Q��� ��B�/���%b�RT+������h���-� 0��T��E�l�϶�G�@���33����e�{��u����b$딶$D�k+����6z��@b�o���YB��3u?y��������9�r�fͱ�tX��{���x��O����]�]WY�nM��k�	��A�O]�(���Pr3vO�f�
�A��BJ�@����p�������}v��h�3���>�A	�RS�Q�$�VtC���r= �ު��J�b�u��2����[8Gx�ZɠF�	�mp���ې�"'��U@�}$�P))��wF��TG��ֶ]WY�hE��k��jx}��!$��偡��h�/�e�S�Y(��l���2���]�\$m[-^W�w<��nJ���8�~����?~��u�E�@))�<m�w�kx4�*��qyy���]��'��GȂ)]
�� �	+�JJh�TeN����/��T+�ͪ���ow��e^���8�ܚ �Q	m*{�X�ogϔ�<}�y%>��n�mZ��8O(��W/"6���D�D�Z����y(�o��f��Zl�4�ݸqG�S.��O�*8V��!�P����j�w�6��"�R5�@��9�z= ��xW�J�DJVVlm^�� �t(� �RSA�o���[���V��:} ���Nv;&5�p�ovh�<��BJ�RSD(�QAŖ�s�f%�U�*+C���<ʵK'�A/rk�f�Q|��q��V/����r��c`��C���C��zy.�m��cfa��7D�P�Ѐ����uW�NU�Б�)������Q�V��î܊�b�R��Lշ���n�#ʔ	��P�L�ѧ�#���bU"v���D%�"��{|����ka�a�����n���9�xz�5=������A
= ��
�	*l�CQڳWm�Z�<ʴ�'�A�Ϩf�QIM����{��#�>�}�(����G�ծ�)�u�b��
����x���T`I��6�����b�q#:�ҵO+d(����{�MY.�9��!(c��닇�wӍ��9]�	��S�~�:�z���"������prlsڠyk�V\jk����uԷ��4D�_P'O����$�HG��y7O\�=-CӶb����FLԣ[6�,�F[5��ˣ��9upn��Ȏ�$H���9�
�A	*�T+�\+7_p�b�U��8@�U.�b�8NV�}y=�tiĤG3/Bff�#�rs7Dd7�ncK�>���ϴƻ��Z�S�!S��9�G�J�?1��#+ff��W���@�A;�k�$�ȁe%6ݍ�!➚��-�תh�v��>��$�H#�= ��h�ɮ�ݙ�]�>���#uϩ%B����}��n�V\a�٢*�"�2�#Ԥ^s��33F�q����f_��H�5�,(A�����.�8^���T����A���W�R�e�T�	��S^�z�����wMN(%��9�ZlU�7',ǝ�
�`f��{j�B��eb��M�M-�û��_�q����+M�ğpwX�����R�b��{6c�ܞ�]�n��|<�FGS1�]& �6���|d"˳G�z���6h|�ܠ1�˚�L�ԭ�7�����rЙj��f	��A5
W:�Y�wA�!�r)�b������/�osXNZ�p��{��t>�N�[m{s^�d'F������5������;���'�m�ve�y������ߗ?q���tNX�Ê���2d�0ei;Vw+u�����g�r�(Y�����o�11���BgY��gC涥 ��#/�=e������K_}�|�.�
>�����ɹ4N���x2��%�yI�f(#�U
b����i�î]R��ܧe�nog�%�U�bY����>�|4�"*��^�j�D�x�M��
� �H��4q9����>]��$yF_��L�_d����_���w��C�W��n-�t��O�_!X�.�+s�<j���a�6���o>��ؔ������t�^蟳[F�N�.o��Ѧe��KBXn��&s�.���b�*B>�#���5Y����4�;�x/��R9|����Ӑ�����U��w���yi���#3}������14\�����r��jR!��V!I��Znŉ\o���3Co�p�Έ�w����~+�g����Q���OmHo�\��PnS4ˡ����Zj�ߎ�O�ٻԾX 3p��@ r'Ƴ���(�: ������k$���;k6�v�۷[v�mٵ�
ڴ�f��lr�Ir�L�7Rf�2ݶ�D�L�,'JYa5�98���d�9o{/L�nY�e�fI��e��Ͷ-���fݶ�v\�]��ݗa[la��9�l�,�9[b���)(��u㎦Z�-�f�It��"���"��lÌ��m���&v���F�q)�d�����L�%#�I�3Y���[4:�tq�k-�R	γmb���lչs�9��p�H�ևN��-�v֬͵��m	�7Jki#�km����s+q����LKC7'hrB@�ͤ�YӒ[V'6� ��JP�m��	p��YYqe��slr*��նv�"�.@�-�Y�[b�l�vu���t��PS�HK
S�@���V��-� ]v��ŧg
@�����v�tu�SM�V�l�c�*�L�oa�{)��J�<�Xs��wY���rl�-�/��b�B�ƫ$Ыڈ��P�S6�2�B�e��磩���b8�8��)���ٮʷ/>�8,�V9��g	���n[�V�L"�5.t�ַp�X �L���^b��D�onA���%���r�h����8G$a��"\e���Ԏ�u�Ei���fݺū��P�PVCGk[�6,��W��������7l�{h��vݹ��n۪{*�pp�.p�F`�2r�q�ݍ��v-�����f��+L�`�K]E�bs��7Z�Y����:jlm������Rv�
uf�d��@Kq�Q�C� �pP&i��5a����`,Ԯ�����c��U
�e���13sEYz�`�[H/0,�����z�?4�;�T%��><���=�vx�^�!��R�c�WV1�RZM(�����Y��an$���\�6vMib�&��`��XK����Ps6�h�$�pgv:��N��}�������6�ѣ���.Yϣ��ݻ$]t��7�'+�����7Qs��0�B���2�hZ3ghhQ2V�)�����a�Bn4t�c�ЊMHܣ�,�Zh��as`�niu��%�֖��	)�T�çn���k�P9��\j&�ls����1����Ԏ���ɗ����dڭ��rMMtux�� 7���q�{�컮;9wM���{rݸ�����w^m���ej:S�U�K���GJ�R}��:�'����Q��ˁ^��썫qq��v9�g�uOh �yT{�:G��b@)�`벪ru��+z���jQ �_#]-��v���h;*���L�)Mց[�X�а�
�)��V��ɹ���.�{$E�Iúr3ʞ�۫c!'m�����ѸܬX��.v@�r�%����i�R������FZe�YU�T,s۴�uϣ+�
�+�n�nJ��3�J�n[u�VX�И0R�=��+�,�lv�۝�*\!e�9m ۭ۩S0z�d�e�e��tj�Z<iN�u�v��pjo���
0��)1 L2�V�r�.�F`ą��1�ņX���xJ�s64s�c�s���� V�&t�u�7�t�Km�q�\��*�α���Ɨf�GJlB[�KZ�S(�0�-�c�������o⣣������$���88�-��J�E��S;We�hїJ��8��k����sF�J���z�ݷ����rNgdӰ����q�e%(SO,�g;�@�s@���T(RS�ʱ��Aʅx��Ш�+3_p6�[�՗G�4A��FF����ln��#׳�ޟq� ��y%:AG�.h�{%�v��yf���T������$��RT(�V�ls�6�̰A��B�d@>IMy��K�k��4�=}@��������W��2ft#��D�A	)�Jt�z	+�.�[zN��Ӑ�;�x��E��������f�A�k�E�*nX}�����2�d`@�D?�Y�ݛ\ccƙ���9�P�.���j�M����O�O��U��Tz=����]�vFi됩�LDm׺zs�N��= ��PIP�D|RSD*�ea��Ή��Ys5�0��"����ӗ3g����v�2!��nX��PS��ˀ�Z��N;�������<��>��5��[�[#�" 9��t<�]�]Lh�a��}!'"�RR+r6�t���."�G�fX�O7>�(�Tx���������g.Le��yq�p ��45РQ ���	*�i�ۇ{
L�a�>��AG�m=|�;9�5��B�ޠOs� �--�ƜǄ���cT(D	IO�%^D�+��%��r�o��R�Z�Ίv��Y� AIגS�}b*�Ղ�̒yS�	�d@����h��-�Qɖ:cM��-��W��;;[#�����P>/���BJ�x�%B��O˸M���q�����Qg�'�\vt�[��"��Jh��
�A�N8�[NO��� �G����»�Ґ�z�*}@�����@!%��z�^9�B�� ���@��@� RS�obg8���&=OE�������;P�>�P�A��f���m�L8�Ĥ;�s7����E�a�N��^ۉQt��HZڬ��fme��i�*ORtgC�_
�>�|�РRSD�T(G;{|4�O��Aʫ�%B��y=τ���\a��4D�Z��6D�'4BJ���|��E%=9�ghb#�[٩��8$�[�C)��{�׈=���+�$ϣ��<���7���n\��,q^�֓iٻ�ؑ�����<��%�3He��˥�m�RO�~}M��E ��oo�t�J�Iѝ�=}C�;��y<|4oe
=�5�
��� ����F���q{�Tz�ByU��N��'��H�Ƿ@�^��5��Q��������i���iP�AG�A	*RS@��u�����-W$aU��HU�t'P �h�=��!%U⒯",�F�^�����:>[�(D@))���wNt�ĥ�������|��"f*�]��2#*��1h��yGNU�(��k4���q ���%:�d.(�Eށ���y������2`|w����x�9�|���S��(�I1�蝳�ohP1�y��
���=��8�^��ٮ�@�RREm��6D��cm��n�Of�n9'd�0r�;	ء0��`,@��r����=�,���c�>d�|�xm���!���HV=T2�
��6���P�S����U��IP���))�*e��əC"  �^���nwtgu<t���=}@�} @Z��)�u@��wp�dx5��(|��IUx��F�v.F��"dV$���Ka^�ۍ p/vh���P(����$��w[1L�՟Qr��s��G��k;�wq��
Ǫ���P%� �h�b��=�C�ܦ+��@���$�iD8�謮�'V�gK�����շI�AՆ�P �� �-t(�SD(�z��GD�}��*����M[�n�s$4G$���"Z&p!�T����a,U`ػ����B$��>�`��ƿ~�4gg"F9z5�k��n��B9�YatV��l�3]��q�i�2��'uº��1�n;;��H]n3nہNz�.M�b�!��d��q/;1��ڧ]z5!��e�+�jYNuy�k��-�[��V��H��dr�4�����oYP��i�<sM��� N/=s�A�㰃�f��@�R���jN"�-����3*(]l{��-�t���۟Cq��l�*c�c%�i�Mm΋�8����*�Q]@��Mx���IO�%B�����|+�7��#H�:.�wT�yvh��3/Bff�0q�ױϫ��h9˨qy�^�F��˃�����c�AS�^�sD��!%7u	x�y��^(�w9���P(� ������V�v8J^�%9���bXua5ޠAg�A]
%>�(�UA�s�_M��&���o:��
1v�z_Ԓ�׻��q�f�g[���F�
3H3�@�h��} ���^))�n
��ry1�����y�����+}��sD��!%>IH�"ì6�#;�Y�\�[���r֮.���SI�i�|N�N�,]���(GF�&���=�ѧfe���{��+�CL�f�6���󮋫��l���F�{/B9R���hG3.s�I�⮐)�?y�KV^h�!���j�jV+�Ѕ���7m���Y\��&.Wuǚ:���)J2�*u�rE��"5�Q��M�W���+�.�oK�z�)�{�:GA{�@��"�DsΜ�	�c�hodP<}$�QIM AQ�'�I9����n�!�
�z��|����S��J�xDx��/�F�t���̋����ywNO+����Xmw�}R��7��y�Ox���%`P ���z !${i�t���W��K:KR�kskH�/vh�H��RRd텲�p3E��URA뫴�Y6R[�{u�^&���O]�ɻ+�lk��r�hX)*>�S��Tz�{ںN^��R^[����	2�5Q9�3�grwfȳ����Fff�%D\̽&�Ɯ婋"�[��`�74!����s��٫_P>(�>�t(��4U�C��J���B?w.k*��D33E��_��~���^��������Y�{㻞��ZEʛ�v�gv�w��7���N��v,�>mC�bN�fb�,*��ǎv�%/r� ��f��E��$�z�`������>�A�u�Jw�����.�����۰��Z��f��}��۟bj�@�RSD$�ȋ�Vd<MI����.Z6��6k��	G�;���� �G�]S����&��R5ҭ�#��0�fk4�ػ��5�y�Z�pK �٘���0���3��O�>/%B�n��8u��Kܼ�#��
���K*vnM��("  ���!%B�
 w'#�Ky�.X��{O�u��rk1���=@�S�!�A�Ghd�]BnύeУ�@ ����T(DJJo������[O�\4m�LV�G|7\��IM AQ�!%#���41QK&�.<V+�%B�������������'��U��\�t�@E�5_��n���ў[�w�wv�G�q���son�l�;�xΛSN�3�Ʌ���r��^uvT�,=O3Ǟ�D^goDL̳@�
33F�3.�DvT�ұ`��:�<�P���wj��>Z�A����W�IPuJ�5	����>V�2���6��1���V*P�^�qn:�̐«,�m��!���C�t(Dx$��:y����p�������Bҽ�4� AO�Q�s�
=$�P))�B�n�.�y�=�����+��>:��R�/+�%��F%B�QJ-�i���"۪} ���$�@ �7\�5�����{G���xc��T>�K]4A����W�U�E���]/�bt��� �u
<D|RRz]�q�mzԺ5�k�@���{OA�=��=�h��BJ����μ�r�v13���+1S�;�{?oKx���� ]�׈#�@����W�{?6��\|�j;�u)��r�O��y�f����P��"�*��� zof�P���*��fRV�9.ũ]]�����\�2J:A�&�`LE
�:��M,��#q3�1�W&��sx������MC�����`��Lr������q� h:�nw%Zh��[tN�u�ks�ɤ[ZuLL��-�55���z޼���c�3��t�\=xL��ztF2�M���\6l�ҝP�-��K1�n6c��;���\aA�L���W�3j��1�at�q���J[t�M�IWr�WA�3�-k���R;&�.��Fbl����0�} ���P))�Tz2�vu�q����ڰ�����w�%xO\�}��ߵ��48�s�z��z�I���Y�n�:D���o�G
���tk�ޠA�� ���P))�{�}�@�͏AYB� �t�G��$�¼RT/sC�0-*e��	kwT<���8A{�D�P���A))�BJ�D�4c�5R��A���Nt��G��vOQ�q���a�ž�D�큶�n=���~�+�4�W�"���)*DA��q;�_a��� ˚�m^>���޵.�`�r;�O�����)�AQ�d:��M�u�L�w�xg�>�poBQ�[\�ծ1WUM�6��[������Mk�V�C{�52���5%B���o�	�Y�����8�=Ѷ�ϵ���"o��Cԡ���fe�e$�j�8�����:�I��PV�Y��r�(:=���8��0�56��OQ31	�"��4]-'jv��B�	��
�+�bu�[�^ ��m[xz��;���mXx�W��8�	,�܍�雏.͏�3/B!����D̻�qz�u�k5��m�R����	������PQ�!%@P�l�#��d��x�����RT(�����/��.� ���g�mY4U���H���x��ٗ���hGH�f�f$��W�e�I����}}?W����|5Xx�P%��P�� BJ�^!%^u���||��~���qX�4��i�\�.^���-sf��'2�7�0]A��O��߳!;]y,����[k��8�)tk��B�)G:'�DH��)u
9�>��R(���1p蠺Aۗ}^^!S�^#9ײ)[�&���8���#���٢%^D��E�C��A[SD,u@�>��⒚�(� ��.cT���yW�4����Tx�f?w�C�zu���Vq�z�����؍���C�!���ъ��U.}�j�3�2(�ZSa�T�d7|����Zh���+=uU��,�fҼLCk6��7�f��kr̞�w��SM����K��c63��d��7��ٵ�^�7ڷ���V���{61��T�ښŢ�������@z
E�����'2w��d7�*��AN�ڗ�}�^�u��t��w���ӷ�W�E�AY�=�&�{��߉���>�=kpe%	�:�l�<}�{ؓ�ڲd�*�Űp���`?g_n�/�M�z�WR�Z�w�EN}�M��Ë�
wZ�:Ħ�r��&Λ����J��.��3�9��NҐ43ݍz�3�s����#��z�N���{��aZk���X�a��w�=�Nئ�r_XJ�{�'F����7b�r���i�g�E�����o�)����5�vUV�h? ��A۽�$��z%�3�{�w��oOjd�ֻ��o���$���a�샢�=7��ϼmM��Sܶ�����l�ﱽ�헧�z����7ӗ;�C"��5�^���>u��e���b�5o�����}_ft���?e<��/�Խ٘�+*m1�6V��P	2��D���z��o+Ɨ��v��_�-ó������7�X�y��kT�x��p��1���>�亓�gc�'4�+���=v!���:�b�'���{d�si�A�qc����8p�
'�7�4�)�W����is<Uǫ�_6ث �G��S��E�A�s��_s_s{�ٷ*�Q#U)R��X�Z��Jtr ���6Ć5��$�w$�m��vP��m�r�'q'E�j�9:93��fq[�`��'N���;m�u���6$��'.�
R�
f⎭�-����
J%�5i���$�9�서�Y���VDp啐��9%�˶��NqI%�6�:�Ҏ&u�8�9���*̉S;2���M�8Y�*2�8��ƴ�r"(��9'3�f���9aۇ[X8mAG��[n̑�3m�I��fRr!B�q��[4)9Gpt\qY���p	$��n�l�iܴ�R���E"J�wrp\�Q-A���f�H�㒲�lq�gg'�rYMhαН(KK
���mդ�s�E�ڲN�ܣ�>e�ک�H���3j��#�}5�����PIP�@�"�4�goL˚�'�(� ))������q�R���#�:|'U�
�bib�f9��W�=$�����BK,i\e�^��YB�;����o;S��W�p ����;�<>��Gis�����&6�v!c[��k\�ʁ1b�V[�`�/0�K���#ㄓi�j%�>��>mP�RS�
=���b{�ޫrͫP��@ƾ٢�<9���RT(DJJk�-�s}-�\p���ڛ+�>g��z��5�5u{O�n�RR�M�k�����ZS�Q���^)*i�x�
Xm���r*��qUJ���f�#�U
�(�))�JED����;�{�ϸ��]B�wMTz'q�ꘞ��nY�a��P>)��#0l�k�����Q��8�g�8ʙ{���B��ٌ
̸��'W+-��:;B��,�l�]��=�^X�ilxE�c�b�Ӓ�-"=�!wP�o*�"� ���$�ȅ�z��H�옜����vq�R����	��R�@���A
=�#��.��Dt����0�̖LZ۫�]x1�73���y�#�)��s4����������C�tzIP�J��_oqʛ��檕��.��Y�:A�
 � AIMT(���2\���Wu!��^#��q���2�-�,ڰ��[�A�BKk{Х]��Q{��Q�<�h���",-S�ѯe������#L;:�)tk���O�@�T(���>Q�!%T!EM[aP�&W�G�BJ�^!%B�U��슛��檝�s�\u��6n������A��z%"�>�
J���3Oj�
0�
I�蘞��nY�a���}4A��I]x�����/��,=x�eF�@����K�`7�@h��-�-��<��?Gz҉t�n.]G��_���ë�����3�9�x�bR�,��L�bfo�7��ac/l�a�nV��t9C��9�^���@C�1����v��&���㗧�V���d}�1����J�5��.nP-��p
��Wu��\h9U��8��h���31�1�51���Q �XNOJ	�;��e�� c&��(g���']�$���c#��rr�N��۳�\�L]F��fWT.�{����VV�ıKbԃ56f���sYJ�W��1n�����69_�w�y�O����DAII�w�]pvu�R������
��e�\�G�A�VЯ�>G�$�
Jh^캵��󯏸��@W�r(�O_a����54��A�Y�D�P��QP�#]Vt���|4���7tW��R(���G��d���J�Ḑ�]c�uXx�P>-�׈>��IO�$�QDA����W�J�A��(�#��⒚�V�w|8^��\�Ѻ����=g(��ѿ:�s��T��U@���(����0�M��vc3���t(�v�OU�o9��x@�f� �U�@���!b1}Ј�z�r�X �B#��̩o�@]��f�15E�\��F	,5]f�%d.��U^ٜ�>�u:
Jh
�ms�虗�v^�+W���a��k�Щ�_g�TOs5532�&�32�����h*�C"�%��I�;9��Q�4��/0[�N�'3<��宼�N���9�����Gӽ	���d�ت�G6��;��	K��#m�q�Å��K�Z7W{�O�����)��[��/�쮺����,�SDQBJ�^)*���U
a��qʫ��sSJ�w�͚� �T(�`�
J|��P�J���@��mm
�榁�"�w�fe���n���<[�F�).��eW�j�F�A�IO�R7�#Nj�M��E�75}��|8Zk��Ѻ�
�">�T(����f�ߗ��k̢I
c�gtu	���+�3�c��A�+x�̴4������~��_�K��BJ��$��m.�5y��j)X��"X��3�6�V�R�!�H�8� ����	*�D@"�=�*���^��/^)�}�m7[�f_ar�[��<}�^��^>�#�$�ǥm�����M�	I�RT+�# �
J\V��+�J܁��9��'s�b���A�=�����:��s�(m�o�z�GC+��[�"�N�s���ZƯ�g,M9>ô��Mbu1Z7T�#H��U��D��Aa��GL�Қ��d�oHB �n�x��xͤ�FM^f���V0�>Y�@��7�`�u�0F  ��4BJ�B")*�Jzr(jō����������oD���+�P }5�G����%"fL�Bz��w�
�
@�)��\�f��:�nNBXx�*�)�f�+W\fnn���c�0|m����"�A%5}����Ӵ�TV����\��x�Q�����D2�&fkC̽#�����\"�P攊1V��uy)t�K�#��>�J���q��M���_����!@�τ$�W�Jk� M���<v�.ݧ�&%��VRp��o�@�}4A�U��JE�T�"Ӭ���S+�Α�H�8����v��'���i:����@��@>R��T�L7�&������Tl��`~O߿l4߱�Ǫ��vM���G�J`][���"�����I�re]T*%5r1ȵ��^B~������١�f^�#�32������΋~�K�P1]��s�%.��v0� ��4F%"�� ))�
�J~m�i����np.�Wv��Yr5kR�]Č�.�i�m!wzU�{Κ%������ 5o�	���J�N��𡑖�
�I�%��r�'��F��W�3F�c@�s2�3Eu+�O[�؝hnj6��OW��uSZ3W
�AuP�RS0��!����W]P ��	DA	*��N/+/�ڷ���ٞ��K��]�<�͟V%@#dRS^!%T!��oF��>KhQƧ�Q���1�}����U�k�@�}4E�_��V⽛� ���W��B�F���!%B�B4��ܼ�'ǫ��e�o8��	�f�F�#uH�
Jk�C�_�{�O��ͭ��Ar�e����Y���Ǫ!�dFiE��8��Tꇅ��te3��u�Ua��D��uxx�a�5�jm<ń6�)	5N{W�m<�ܜc���7,��c�llr
�{��npQ�5���T�!����c�9(B���Zͅņ��k�q��͖X�GQ�+a�v7� #�&���i|�����k��ѐ�@�g��p�۔,�5�����Y��;ܸ���h_6J��1�5�d�G,����hdp�k�im�0KF��)�����"vvn.������p�z�#�+G�`�u��s�9�שqW��y�y�1��:٘���(�٠}�G�IW��%B�������d�fU�<G�Eb���f�׻B�C0A))��U@���>�f�莍����Q�#���&�p���j��p�|y��>� ��u��c�><��,� ��4AIP�B1�|���η�C6�^�L'�ۺ�њ����B�Jh
�A	*���F�ֈ�sD�׊J�x�,������
�� �{4�le�
 @-��Kh} ���@��n�Jܖa���z��&��18�aڑ���8�	*�U7Ͼ���|��rV�c"�X�����]�^�|���qɂ�D%X�,�'�w��Hkt(��%5w���W��wSZ3W
@��w�V}���@湠*= ��P �����4GF:y}�fQ�_k�z���Ԋ��	����%o}�
�t�s�p�������ظp%F�c�_�=R�����qD�6�xkhH����J�x�,����d��
� �{4AĨQDfLP��*W��DnmP ���
 ����T���q�	��LB�N5Xv�
Ϧ�=����JE Q�DTw��U����Gs�E� �
Jj'o[�\5���'E����G���W'�؅��BǱMGG�J�����إco�r���:��ĸܻ̔WdB�#����#X�8>���p�an0�X?~� )�T2JݠuQV����r�Tے���X,��U5�O��оe�{�4�e�ʔ{��1I�˃���1Xv��6�Rg;_[��Le'ݲ��sF��B1�*�U��@�������@� �y)�3[�����cq��u�G�f�RS[��(�jg.�1^���(P'w��(�T+�$�`�(۠�_f�ٓr�*�{e=J�:���H�W>����4�6�#r���\���8���$��+�j�S6
���cUvj�a\�ː�ȅZ�F9�^�?fh��TDs2�35�a/�����)�� ���QK��G��Ϸ��\��q�õ�	��DT�!x�O bW)��{������|��RJ�A�a���<�Mzf�����,��ތ���>�A�k�$�A�J��0��b�>���uS�P�&"A���k3s��p�@�&��Ш1���Xhc�K�|���0=|��Q����IP���u˼�	vD*�8�S�q�]��u>`n�y`�RS^!%T	G��#�n����TƂ�C>��ۊyҾ^��õ��>��A	)�)ȧo��1��
(��k�$�P(� �����#��,�ۙ��cRY-����@�>�k�$���{�$�
�M#e�%,|���}^IP���u˼�	vD*x�
��!��}�iX�����1�$E��޷ba�N�2qq�V��Q踔�.J#`�>���ǏI����4 ��98�n��X����w��% " ���@��Y�n1�[L:���#ms�N����^�x�:]@�}4'��BJ�x�����_%!H��I@�Q0��Qh��s�χ�\��Sek,2�6�[c4���O��,�k�^!G�Jh	��]��v��KfwFj�C�T�':��#={B�s���T(RSDez�cc7�S�� ��
��k�B"�>r�.t�ȅcO*�h%B��\���K���]
ȂIW�S���{Q��5}��<�a����t���Mx�$��%��n�C)^N�t�M�M�G�Jb'uw�8$�[3����=�^������y٣y%~�J|��շru�Iu��u˼���"�{>Ĥ�˻�}�oj��bGò���)�`]5~�@���o�h�$���r�|�t[����V�{ķC�/1��D���U-�z�Ň�ի��^��J,�*�ֈ�biZW�>#҃��W4��-��v���z���C����^���f�j�����\��_]�V�z
g �k���,�`o��f��]�|�7��I�E9ճ��n�][̸�f��-����Gz^c%�ܹN�3����e�2�ۑ�3;v��ӚT�ۮĵ`�[�uζ�H���ml;�}�mw8=�3�������"�;�^Y<����}�-�v����� QK͹-�t3^��7J��*���[;�{�4���`���b]�����ׂ��r�@�#5�P!�UAI:6���L�{Eُ�r�������wh�{<�!�s�\0�_z�)ǫz�\9n�����2�s��U��}Ǽ�z[=u�I<�=���v����F�p�'���}��wiȖ����Ϗz�U����]��	U��E=6��n]��jڡufYJ.l��z�P�2�a=�}����5���m�U��i� q
�=4^�'Ʊ��~𳣊�� s�!�v	�j��2E��]�P�����بkB-� �in�H��pm��L�褽�U����c;��Y�C;
z���`�ˡ�Z����{��a�t��͊�oX��F@�B1i�$�S~�o)�jgӉ��i{�J�����}���p9�����q�2���BT��� nocv�1�"e��r�����ש�[}H��7�U���Kb�H�ʬW�U��01H��t��&�b=�GtWR�k9tqȎ9GC��]�%��R�9�d�Kb��J-�M�,ӎ8�)([aD�v�DppgL�t�:I;j�u�T\��۠�FZ��j��f�NEn�
N@�3'.
;��38� �Q8 ��H�.����-��m�r��̉;��������9�Y�I	q��NpNk�� ��;:�ڵА�w�Gs��$\q�efu�'$�%Ju[j�m�IIM�m��V)v`I�w9�ɖ����D��]�we-j�ó���8kp��[�&e)E�"�*r��H�&��s�Qӓ��X6�m�4RY�pmi"B��"�9)ēmٕ��8���4���O�[��/e:�)�fg6\1mrۄݮ
��7o��o��v���睵FSź�m�kq�]��^{*���W�3t3e6neha� 2�hjhҲ�\Ųiv����l�54��h�����V��`;�m��1�a��{]���Cpt7J�� �_4b �eq*B�kݛ�^��h���u�zt=�M�<8ܵ��b��*f��y�g��ہ�K����nO7��i�娛h��q�l�鞱��Mn�c&�m4-	ur4݇�04t]c�胥�ن�Y��Q�6 �s�`�X0��\8����LX�u����EK\%�M�ւk��N�]��s�r=�;��+�X�S'm:_]nͅ����.���@
%F�0b;n�sūc����^��3k�ҽT�m���"�x�����KZ��t0#Ֆ�˜R�+�n����}��;&#0X�0h�8���u��j��]��t҄�K{��H�QWRaz�p���\�\u��*nHJet��9��&�#5�B˖��k���̕r�ĝ�E���F�8�Wnq֨�v�����c�����N�(��Q,)� n^��7$��X��A���ܤ��K�ǜpz�e��\<��:î)��(��m�0��٣J۞��u���e.0�]A���ZKU�Z�B*FӵL�*,3�s�8��IZ��]��8-y�lf�6�m���ח��t(E�go
`Jw�۷��WD>�k,��������XU�,�Z���&.$ݸt�M\j±'���\8v�e��b\\eKI�����o\$�ƯZp��WX�Si2Ģgl�`ga��㌃M��{w���sF��+��=�9��^ŷ�:h2�s]aF�@m:S��-��{�1ȼ��x�Wlh$ܻ�.���ݶl"�h^5��n�޸n4�1t-�N#k��hM�f�F<��4t ����%�&`�+u� eЈ�Q�E�JMrv8M�y�r�ԃvv����.y�V�x��3�$Ë�>��\�;��r�Xݛ-����L�ТC.86�HF��V0n�	��cf��vP��N5�D�o�<��n���]�6w]J,�q���].�pm�1�B;0íg��7$�8�d�g�W�H��M�6��<@���^���b�Ӕ�bT8\����C�/���\�����wa�fP1����1ηT�ػAJ������.Y���9��=O;���:R�����<'P����W���>�׿~���Ͽ�������7��-��eㆻ�1��Y�P�̯gF�$�(% �x��u]N<J���ٮ@��I�=9�%�ٝ�]�p됒T����[���T��jRQ����x� �Ю]����8+�Z�(IO�R/yj )u9�ù�b��H]���>}{����X��nW{�ܫ%��U�J]q��ېI_�RITߩ�\c-Yx7����i�}\��̬���xf��JBF#	q�mk����1pl\D�4��jtխ��;]1���@�H52hP�H���2��}󄔄��cWܣ����xan��*���B;a4���I$��z�]������=cgWO��ȿ/MCgI�U�����&=�x_:_�,웷�V�xB�vlK�ˆH�Ѣ��;;�����y����[�/�e�r�ot��������*;�v�3T�$��$�s�]���Y��nk5�n�$�Z2� �<3\�%>	BK��3&�I�M�����$�I��w��9ᅛ�W�����WVN�PӐ����IHIl��!�� ���ۻ��m �9]��;�%!%V�gƃN*!%��o������ô�qsM"]��!��^)��W�H��5 �59,:�����)
���$�^�y���#m�3a;Z��(IHIO�V�yNћ&����H�]��;�����^���"��v�9#���ss�n}��S���I�K:Q�	��}臿l-�x�z�Y��/���������I���ԵW�%�k(�zu�VIR���B���zo�]��\���̓�i��=z�5�ƶPv���w_�RRV�1it����� ���I>��$�^�y����f�\��צ6w�j{��%>�J@JJ�2Ec������3�9��W�١饻�W��HJ ��^�1u�������y,c�!�of+E��Z�Kv�e������5X��������J|�>��M�oƶPv��
pTnڊ��8Ww�8�S����%!W�p��:/a+�q���%JO�!����/1s��R]�(�Ѹq�i�	@	)	)9�ۚQj��k`[�7��C�Kw���{�%IHIr�6�{=��=�)G���&�7�ƲPv���.�*#� <s���:�&�����4~:�8tuo;��(��nb/
��#*YUrPU[|�G�*�$���i�5>	9(�J@IHJ�j"g'E�۟e܈��}�2�J����]籚�%>Km���iC=�~�0p�Éad��P"T�؛\&�UZ�x��v��M��&�q�1����
m��_wu���+��;3{l�4�xl��{kn�7�ŗ�;�}����"�ҜG��;b���&�7�ƲPv����<�K�;n+��J��9HIO��y$2��K���TF�󩞦W/f��kI`	G�T�O��{�݀f@��<�%wt-��������^��WH��sP3�����$���19��+�o3yj5����!�y%>	(�4���k5���h?
��o^��K=M.����)j��XEc'V9Ή�U��KQww6�k�����5?{������ǂ�(�;�Wac���I��Nŗx!RDzhp��ν��>n���[��(����!uu�fT�b��c�&v��Ti^���������h�b7]E�lPƴ�q��V8�S�m˵ȯ<JM����5��,#�.�!�L3�t=b�98�6��I�f�0�\��LV�	��9����ஔ��nuRˡ��0�bkmA��F��/���jM��|�������a!0 �`�f|��~�b�`��!+�]��3<��M�%���fk���(�d��B�<hM�޴�nR�$�Dm.��	,����!۪kngh�Wt�(	)�IO�5D�Qk*�7F�N�t-;]��E�Ioy^�T��K��m�T�̝PJBJR�W�=��댫Z�7���Pk����	)Ij��2�DFC�Mr�s����j���	,����c.)���Bo �r5BJG�S�%$j7u���wu;""�V�����KWx+��� %$� ��ᒞ@g�k�f�j�@��hd��F�j��״"n���}�M�#�^�L����mH	)J;������m���/�g�/ve=��P��Հ���x$�
�KT�-OY�ٰ�F��B������ǖ8u%9t�7GmF�,9=0'���jf�^wF�{J���b����Y��T��YJ(fs�ȷ���iLF���5�%����}�7\��uC������୐+z@O�%	$�v���E���Y�w/(p��\<�V�(%))�x�a��0f�:�������yvg%�jc��]��#�C��*yS�Kwܔ�(�J|R����p����[�}���-X�K�������I`H��&����c�K��f0�r�wVP�Gj�f�нFXV��� ��P�QB�ȀH�bc����В�S菗v�7���p�oWz��F�yM˯s���$� �Ҝ�{U'1��PO=��ڔ�q�k��t�В�Њ�\=@��x$��G�J@�[n���汿Z-��N$/k��P����+˙~�k�I����t�Ҟ1ӂv�������Z�xK�����B�h��j]^>�n��y$���;5�Y!V`
�+ILG>�Wq���q���[#wi�Lճ�e�[��|���R��u�"�o�����obX�ٶ�XO>�@������5���B����4N�n���6P\s-c�g4�Z���m�l�BZ�" �\�O���P����wDt��Վ�:�|"w�[����=�|�J�R"컛�G�X���3y+��K�՗x�iw����%�y���EʝY 7	)�JBU�}m.e�W�x�4�m�����������%�q��j*���o'�J�.���Q��ux�q{��F
F����ee�5��ݥ&�Tf�"Ui��w=��'r�/Vm�%����G���h��4����e��ũ����y�2�-n˱��$,���� rIX	)(%f�67cP777wR'��oVEnw"�c-��U��%a$X��sw,�7�"�QL��%�(@�˥4����둘�ڑhJg$0@֬��os��OzRS����]��N5�x��ӊ���̝K�ۂ�5�IJPJob`B}�ɜ��\��p51�K��:z�5c�n�p�>Id�f��@dj���¶��7 %IJH�ନSݷ/�iۚ]��\���b�
�}�$��ܴ�Y��q̇t�Fs����ƻ�Z�j5��C�} J����B�m������%>�I.s�SJ/��^7�"�oT9��Ձ�sx���\�$�'�R�
k�p,��r�7ۧ�W���v�B����P�p؄!m���UPg���V��ho��|zm���I����u!;��y���i@㕵̨˺�����Jh�GWgF�ZʗBl$f�Bbm��i�a�b̰p�{�䧮sʥ���=�bd ��]��\1��BV�E�M�t�#��q�\j
�P�S���Cv�ְ��ZHУF�n�)v��	�KKt����af�m�ѭ��g��$.,7��<���tf���(^f�^2\���w�뾻���Yd�8mґ[P�k3uaW5 �s�ۮ�D���5�{�#��g��#\ ��$�C��ʲ%��\lV5��	u�vx��<��$�ģ�h�}�b�O(�}�<��׉�BJ���5��.��䑨.�L��ې��%	)��*h&�m5>�����j��9�}��-r���R9_��ڗ>���Rt�>IH���ʲ&��\lU��U�Sz��+9g���J|������&��y�㹕>����%��E��>wO�BJᙝ�����6e�f����������6S"�r<c��9��elj�˰��Ee`k9d�2����+*�t���n�*���1P�;j�Gv��Ҕ��$��h�{zv��\5Wө�,��瘞S"K��z��Y�J��=���5�k��3�o��������f�
���~��S_�Ĝg?ٞ���_g*țk�q�V�yV�Z�"2�Q�Ck*id�j�����%�}4a7����M���5�<P�˺B��%!(���[�)�o��8����HD�O��OnF�����' �</4go+͑�%!%#�BK^=~����e�z�"m�E���\l�I+I[��.�FA3���4<n�`��\Rxu�T��V[��7%�E���ociBL��jRS䣺��_[���(}F0Ik�T��C�7�|��% $�ނ!m)���K�G�R"v��=�ې��z���N���Iz+��co�\=�Ԅ�$����n`��V�,RFu�O4�v��M�s��C6�.�rh6��ZZUAH�����żk�ڋa��[6�h�0���o4�qsJa'�mh�<m����s��pot[�=tk�G���i��)è�x��>��[��8ּ_���t��ȡv���/+.З5N�)ۋ(�omS7+Ɏc*�n��g��n
4.��ξ��O�鸂����Jͣ�0g��7�f�rZzb!sD�H�{�W�@��z��sxu�)����r���խV����7X��d��/x���ۧ���F�@wp��ό�ﳦ���.!��3�΋Fq�-95�)�F��($m%Ma0�F	05�n�SEM��݅���Aw�Ϣ�dHٽ����"&��V���3YE;VhnܸR���Җ��
&�-q[k0��2ȗQT��/s�L�Q���� �rLy#9N��H5��,=�޽�{�����W�ש�ȟz}�=:5�{�^����M��{D������ D�F��u��Ɣg��B��,.���z����ʥX�2�{�E�U�K�2!�zُUM{R�f�B���0�m��U��X��Ua�^ݘ�
uڶ�s6`���V��M�7�\�c����k�Ʊg1�����Ƶ�Eŷ���r�=����{�٩̖���ַz�-��~4,�ۇ����Ӷ�t�^`�zn |�f�#8�C�/�mHh��=�D&u�Xg\)ׂ)� �2�٭�yD��=�=��U~z>��NB�����||�)��N"��$�nHD�8�r�ps�$�Ý��@�䬻8Kf���Pt�&��*N-��\p�8R�F�8�'(�����:$��H�̒wH�E��G6��#k\�'I"L�I$����q%�\P\ ''s��GB$vwYngGDs��r��rH\��ͻ.��� Vi;p��NqAH����X�j�%��8�kwfNdKj�:;���eYI�%�rEf�Ç�NY�Y��pG	�')�mƈK7;2�N;#�ݖۑD�)ȸ�K:.-�vhn�G:�kD�`���Ŋr&�4\m͵���I+IJJ}�n�q1��N�K�g��e�9�<P��O�6��\F��Ԓ�䔀���r�_Hڗ�S�L�^&z9�JZ1���N z�X��)�q�Q���f��ڼJ��(͠�����ඌ,����+)�:�Q��(����ry�J@IH���9N�־E����\zz����fd�G�S䔄�Ď���t�l����k���G1��xs��NRHΛYC u��y'>IJPRs��bw��m�A)�^���.��я^>N<��IH	BJ@4cd���u<��ς��Ғ��=ٽ;7Z�sovs�.���{�ә����礉������s-�)pv�?d�nsܲ���>�u�/J�w��&A��u�əˣ"v��xsboU�˾�8ԥ% %IHI>�q�]�f5�*�ޣ�������$�%�e��r��A�r��ݘ�ZLC,zͪ�h1�2�%e%u�;Y��mS�k'�t�IO�����t��kF=q���wB���D�/z�H�Ҕy%!%"���r��w���R:g�7�f�_"�nm�yV�J|���D!�0�]j��������)�v:�OrvWn�wr�+1ޣ��ҟ t�����$�dvu�U���gH�% B�O��K���c���p&sF�Jf��ג�y%>�JG���U��'���UN_nt���"�n�oxR���)J 	!^��"�o{W,2��w���Y,Cs���ޭdg���pn�@�q��Tm��.�L��Q"%waǱ�0�n��ӳA
�[w������}��>�>}����۱��,�!��e�ZfP�J�E��ɸ��k���F�q��X��pg��BO^M�-�m�N���|��Q�Ĝ�<۝0�������qn�)��ȶ���y���s�nk��\sq�r�˶�㧬�]��ơ$��nJ�=���Π.��u֐ɘ����s"T��ۖZ����n�`�&�nnt�Rˈ��ÃB&Q끓������~��n	6O]�N��(���h���Fťՙ|��O�^������y��ƻ�f;hk�����Mr�z�%^��IO���Hh���Dg +�-靥��_K̶�c�����%��B��$�r@|��BJ@I2VF3"va+�]k2�j�\m�-�{>Ԥ%	)	)���Fp��6ǲ�^�	@u����Z�N�/T>��2T��wL�zqσnR����!�Q����/ڙ��5���-�q����=r���;ǹt�����	�|�I��5]��(��­k�s-�`�[.�R�5��K�M_�7����̹��O_^��;ܡ����U7O�ü�fcw�������qDDθE�X�L͵�*��f��\���1�F��t'M(o��[��PN����hK8jq{�>��+4%��w��\,�j�Yb�\�=��D����ʛK4�P�a���8	+L���n�6:����BJR���/�dNZ����g3W��[Z���	Ǽ����$��U��eHط�� =rI�Ou莣��+�[��f�&L��˩�[�dcS䔀�J�H�(ͩ�m��9[י������v^�>k�pr�������t��ߢ6�i"�-�8Y]2�����3:�\K��`�d�J��1�������G�R'k�w�{������h�7�ͮx ���%	)%8on.�q��3&<�Ϸ\���;�G{�8Wu����R��u��t��O-����%�G�8[.�3r�{TT��9��9Q;��"B��.Qj����d������:�D��7S�7Q�E��;�78�\]�ۏ59m�H��{��}#���IXq�
�WdVUz�'��$�Kw�zn[V����٧""��W=�{ҺJ|�J�K�v���r�*AB2��YIՑܡ�ˬ[Y�$��!�5E�����<����K,-A&�e
�(�MXYqy�H��KPdѪ (I�+C��$�%����Ҥ�ڇ�x��ݽYSU� v���)��IHxf�d�S!��n��M�qjz��']f>�p�>IgGKܸ^�W�������� %	)�J��%�z�nD)���H��eeR�W�I+�JRS錪 ��ޘΘ]r�O�Q��ƺ9��"�a���}=R��".� ٸ��㷒�N�M�����9�n'�E��lb��J� �3x�ӿ�c��p�H4�����V㎞u��f��ت'�W�;�W�I)�蚋�h>�Sr��8.U<��p����	�\���\Oť�c���ɝ��Zx�N������&��h;k�x�,+��*5��(2^�c��%)/�'���<��o����.��0������J|S�=:�f�u6�n�P:k��撤�N�݇����Xpvn5��܆(����I+�HhU�L�Ӆ�m�]Jt�8I���'�֒����^
���w�,T=�F�y%>s5����#���l�6@U1|�h��4�S��J����32��V>�"�fc]�R���{���t�.���$�vq6\E��ۚc2������ù�󞛜��x��5ַ@�|)!�7��03˃y.W��ಌҒ�AO@�n8��퇦K���4m�z�y���ű �1�%���Ef�g���<�:z���G6{S�ĭ����vKk!b�n�+� �])ب��ˋˁ�\j��U2��2�bF^B�P˵���2.u��AZ��I�S���Q�7vZdl����A�;:݁�^�s��tI:.�%km�RԼ��mH�6p�R��d��\�@Z;;_S�ߔ��fAR�@�&n�Ie&v�Q/i�T�r{�{ܜ.�4(&�/��$ot�%#�վލuP���S���Ѵ�usW����Z����$�y%"���P;���O��zf��A���r9+x,���)QV����[���JRRZsa��F�W�G4�R����}�@]	)�	)	@]�I�z(gt��	)��o�F��K�q������v�A�[�.�۴ھ��ֿ�?�pο��=�jO���,����-��݋���\��·���� �h:�^
��p�J�vE�1�Kk����P 1Bj���ہ�{�`n�r���ڡ'�[Kv<�щQ�y]��7vF� 7`p���t��*p���By"��E�3Q�ޓ�	~5�^���|N��V`�ǽѓ�t��p����'DfT����S��{_v�wF�WB��=��ڼ��os�8�_>�s�+�pӫo�w㖜��2-	���2��>�m[a]Rʄ;3Ug[g�)������-��۱���$�Gqη���v��;�j�ޚ�[��-sDs3��׻�7cwdٛY}�.
�'[�6;o�CnS�o�5����uv�����Ã�}�k�A	[�%��pY`�j����\S�&�n:X��.����̑S�</�@΁��!���q5���+���n����F�@Ώn������Z7L�R�i�}>J<����9ޚ�Zw������i;���~m+^9mV�����{�6���]���i{�q��ӭL�9m�{�v���2���(U�d�ͧ�5�f�6�,�D~=9���t|�nM^�a��^D�J��x�Z^�t[r�[|���n쁻���!A��R�c�P7v|�]��k��%pW+x-�!S�sm��lk��vǷ`{v�6��]�i	�K4&��M���������݉��j
��y�q�;0u�B����y��6n�Q`0�1p�֭�\$��4 �dNFz�<R7whCJ��客�T���}Z�	��"j'�j�>�ݡ���#�D{I��;7���Q¹̫�����-�n�h�B��n@���>�6���\�؍����95,lm���7\��=�ۻ#v<zt���͓[��Bq��Zc8<Y�Sj��\=�;Å�����E[����}dT���S��ěw���o����� ~���~=��Ű��H��W�R��?'}�L��+
���M���k̶�̴�j��8���*�jg&���)�y�s��l}:��ډ�޽��,ߡ�qI�����&�Jㅵ�`䲍t4l1z�-B��l�Q�.C|��L����ݟn�>�|;��5,lm�ز��F�S�;�=� ��ݏn�i�(J)ĻKz�iS�k��۱��tc�u��LoEt܁�݀7v�,��;��e&*�D�U��-�b�v ݍݐ#�b}p2c�^ɃJ�s���]V�wm�j^��[��-r��ӳ%vY��v6&/����7wuxr�=(��b"g�,藽��UI01�݀7v|��z$����$��HH@��B���HH@�y!!I����	'��$ I?����$�����$��$�	'�I	O���$���$�!!I�$$ I?�B���$ I?�B��I	O���$�	!!I�!!I���e5�	�'pN]� ?�s2}p!���                                    3�P� ��P   B� � �*� QA@�D�� PAE�Q@�)@@   o}
B$�"��**J�A@P��BJ�A!*�J*�$�
� RIIUU	T�*�A@�R�$T�  ے�H��%IR����� X 7X�n� ��E*�z��� {��x�s 42 s�)W ��z�
R�U  ����́AÞE���Ӡ;�@A�u�� t�TS�;��z����� �c� pP .�  x��
�)EPUDH�R�$��{u����
lr /)T���C�<���A�� '�� U�AAAAF�tD������ � �
P��  �� ��h���PPPRz�<���((( .����h.X()y�4+�\��s��&��/0�`����� R����  �T����EU$� �*}�6>�C{�(S��� ����� � ���tT��
��9������J��  ��|����� z�����Gv=P��� m��G 1ĥ\��A� � �
�AT{�  |�JH H U����wpPw`�t	�*)p��A�]��݀�	� �Ê ()R��   `�{����&�;�22�4@2 cȜ ˥ �5Af�� �(�P�  �*A UE�
(P��=L� �{��@zw��Pz�� ;�h�`����<l�X w"{�s��z�)  ��   w�;�Hw�� {�R�]�B������XP7{� ��Ω)W ����`9�����* 5="��   �~L$�*��?L�R@�i� #Ll� JR�  S�*�z��@1�&�)�*P�G���zj{������s��W�I?�Hp���������m۶�??А��$�Q��	K 		�HH@�bBB����!!IA!!�>w�����?�5�oO��,���^���Oz(5��NT�'g8���(&�WE���������o#V�]2��f���c;A���l6pnr��f�=� ���*k�=���|�0���|c�Qo$���.�Q�A���׎�@|4�_��ti�p�Of�.'�}�e�B��J`h�Ls3����	
v�f��ශ�;XY����YY�V.�=v�]]�n{��jԴ˻��o  P����EZ4��r��RFj6s=p�{x�H3�M5h �=��nl��Y7g%�2c��j	!K#;�;�<rU�G�u�7=��'�0]s���n\:���l��^A��,��ob�*��ݝ�1�t=��ѵ㵞���dL��e�1�p:���{p���0�&����7L�_Q�.!��|05J;�۪�9�J�l��ʻ�m;�����芘0bܧv����]����6��t6���u����-J���R�;��ww^GA�3.b���<��,�ݫsW�AiY���H-�6�t�y·]�G�=K�nm�즞�Q�2��!C�"�����d��R���=�c�k��3j�ѻHǊ)��}lr����a]��፥q�o�u�v[��6�G���,�z3MC!»qM|��˧��h�ϑ�Wdk,��3R,eK�Ux�\�����e��wN����r�ܱ,yy$wA�� [������ zv��^չ���vL)�LE�y�L��nBeӷQ����캲���ŋB�Hf��f���ʐ
�걾�f��{�������c�lռ(�	ɫ[-Jiܙ��6��bқ|��8mV`�Wz\)�2\��9�w�J�0�)*��	З.�r�i����v�����Wgb�8�v�^����Ž�+w���)ۂ9�E�sz�bGE3I{Lݐ��']64D���-� �#$.q�R�o*���x�;NR��N�����H`ۨ��u��! ���e�*�Νܷ:���F'�O	��b�K\.N��vu�mo�.��N]�ĳH���bz�J�Κ5��u^86�Sf��t{�a�� ҖZ�w�,J}ܳ��F���]�����Rf�^�I��^��e=�&��ò4�������5Ƽ�ܢҶH��L��7/`٥w���jr�.Or�%m�ZB=GU;��5�͝��`�,jǗ(���x�wWEʝˮN��:_;ĵǾ'y���6fǋ��[K��paGk�8�j�Hk�y�vw���]	V[�A��=�5�{��:d�S����#������5��s���r��z^�Gb9�j �y>�Ž���\�/m�Քwsg9���
E���|F^]�(q��@Àvn]��5�Wf����W��K�$�e���kB����{�̉R,�Sœ:�Xg>�l�NjX��@r1�Q��P(�Ї*H��7st��l�kB�oe����y�^��w��F*��2��+�e]������7LÌʷsP�,k\\ҍ5��v�q�Rr��)܍��l�^1��������(�K���e�15i��":dcĚ|�56W:��8��v��w��<ن;�\!t�L&�^SnF�t�!�>�*s)����"فU%V�E��v��5	^j{���w��2��E�=��Vr�1Oq�jq�P��O�}ػI8qL:��H�����Uv��E���hC���d��p�'��R�NmI�����'�
y����,\0�}�r�������磋|	��v��Vu�k�zX�0�Gn��{\�^o>�Ln��({Mf�t����Ն�Q	�δ�θ���,�M	{8�Z�%�}��������=�,��կ^s(����h�m{�����	)"Y�L���Z*�r��� �7U ��Y;���ۻ�vEN-x�>��e�!��b���_e����Ƶ�������l[[�r�S�`�/C$�����JҔ�z�����ۼUʈ׺�,%����;���h	��KN5Y7��n�ls�t�O�՜��I7j�:��zXc�!�wC��q&V-�%�L�:�&/U k'lH�.�;_9:]ت�¥�%��6��P"6:z�]9'���!�����e7��"��{��&��n����Ug��f>�m���t�e�m[��F�UpZH# ǧf�٤�쳃n3@��w	�z�lb�yna�'h
�њ�K�����1l�݁�É�Ñuݯ2�<��x���;;y��p>L��9n���[��ԫ�v P-�t��unҦ@��mn��SE爲[�5p���/QC����!��,�Oo���J��e���C(/,\p�Glˉ���s���$�k����n�x�l�7x�1��J�`M�@�G��s<z�<{y�!Xѯ^�{A۸���e� es9�b�ۚ�R>{sa��5�hUC^���j�+/8f���{��y�q$�\�����ߎ��Z#����Ce�b���!�zq$3�6��eK��p ���F,����$X,8�-�3ۊ{-ׄ��)]�Ԛ3��0Տb]<ƣ���8� �ٕ��A�vjGa$�{�47�t�3�ȵjf$�{��ե����*��{q�r��BӢ��k�R;9�:Ś͖18��`�~j%>��n\��ltjD;x�K���q�'T�Zx�P�a�j�e#��<�ec����X�[�s���E���'�f���<�>c�ίh"��_<���q�=����/
���S��򮛼dKL-�Smi֥|��Z��9}�6`�ֿhR2�Y�q��ޮ���$a�Yм޽�f�R-7�v���]���'=t�p��n�G^�A&�!f�d��0k�ի6��4��
qŸ	�;2
 �c [0.�Y21^3��Y�-ܜu��K/�#\ڹź�ph�K\* vͺ��<�����05w<{3�՝����-('�89�n��NL��ܽs�� ���\�򉍙p�5@�ä���4�Y��[z��u�<�<�Uuu���z�D�hܯ;,�(�<oY7bKTd��f���1�M}�Ʌ�;f+�7;�����.|֬@m0���&�����E���Q;��)�(Fu�	�/��{���BI���� �)K�E�I�	$�XV��+@�n��BcZ�8Lɺ�frܰ>2>�cF��B������.�An>�f�ܤp�����!&�n^GL�5������9$��:W9�p��v�9������x��e���p����ZsWs�^�V4J�gl�i��F߅���-��� ��g.]�$phW��<�=�����;z�4Z��ta˓����|�c�[J��&^�%�S.4fѹ9wsy*+�]G���;�NK��#V�0k��4��Ig��j��ޡЇ�{�m������9k�L�Q8������ʦ�l���������qܘy\���nw���4[�
=ɴ���:��/�NWED��c|q��.Ѣ�����h�姭��n��x�-Û�r}���\Qh;�^�Gii���]�I��8q<Ѳ��''׷���ic��K����҉.��k:�E����n�	Ļ+�7��H;Ȑ��� ��{{�h\�dk<,9gk�GG�P�q�Q�ĕ���ܼc|���I�fD�}�ݿKwl�CejY�f�M��m��3�<{W�GQ����oK�3���1�Wgq4T�Ը�m]�.�i���[�Vi�n�*@��k�C����xa��^��-��G�X��ۤ@�ݣ��ǧ�O5�i��i&Le�k`v��� t�.�m�7��TwJ<�<a�#'J���>2RtG���`��Z29��wL<�e�ۖ��S�km�02_B�����%(��]Q��0�����>��uc�;V��Ʒx��X��c�4'_��Y�K�U�׆��6i̳��':��, c�ziz�cF.��{���c�""��V���b,u����:ң�S�E�v,}2��$���<y0k�X�ӧ��h8gwv��n��S�p���Ɂ�aKh��{�@V�pFq�7I�b�ǰ`�(q���u��@�f$ ���밇��t�L�g������:��(&��xj��o���H<wGK�n��B���}ؕD{V�5�F�X�X�{'�⪝��Þ��K�)��3��#{ ��DB�wS��ܶ(�C���wȡ��{�ށ���/q�������χ���\3X�g?�
�����h[�3oa�ü%ʖ��G�X��u���3�G�Q��s�ka�Ҵ<���S]��Ou܍]����/@F$����b�sF���!�&��]�^����lŋ]���C3����'f�H�H������C���r�ޢ\��싲lWy�N�� 6�ovf�ø{��P˃s[y�Ma��[&�����Z����ڙ!1]�5���k��NOk��ĦT�:[�œ�;��װI>����lO׶ޫ�f���_+�S�'~��P�"�σ괾��^��8�qi�Q����9�[K4i�"TpO$����s�f��_4��Y��C��%�qVN�pg
ɺ�|9���}�}}�v����cxF��OH����X�L��-�4�nӫ%[�����C6p�(%��(5��oJ]'��^���,�|�s�;:��1�_o4JwN\c5���;�KL�#+��n�=��fZf5�ƯXy�8�Vn������l���]�v��Ѵ��H�>�G]S��t���\Q��E�Y�Z/3��ڎ����� {�iҹRs����yGu��.�k����@�dO8��m�Ǥ��2����J\�U��f��EZ:�[깋@���(����)�V�X��ref�����[0>d��I��m�)�d��jƏe6�@�ok�N/Q��5��� A��^�I��r��I��;�L�|�&��;3a�pB�ΝځZpc�m�Kܼ"nI����4l�릻Z��`��O+KC�w&�Y:����.;�.=>\p�F
>�>Bc�u�ha���Άc��1n��YL�Y\��sJ�L��e�D��c�p��������u��7u�{����o��������=���8��q����xy�Ӈ�ick��3k\q=mYܦ�9B͉(��V��w��Z����>�[=���J�z~�,hս�fq!����:d.x�d�6Y���:�w6b�H�/�Yp��,�\<C��ե��cR�����M�_%���O��4��5��c�t�������vn�k�o>�׀���U�,�+���^5��Ͳn��AIǧ��GL{�]늝��U�~U�vH#��!Z�ic	_%�òk>Ws���]���b�h`[w;	�BZy�U�q�����S���Q��n긡8'}hsK�z#[/4�[����b88��{lW{5�����r�Z3T�:b{y¸��nΚ��7��m�t#�I%F����$aA�;�5�lm�;�N�7'&�K�V@�9��g�K�r�:c�}uƾ�����aE�y�7�;�$��"����6��)8c��d�1�ĵ&N
l�
x�����W.�����.�Q��� kk��H8gM�wӕvЬ�ّ�;)7�'�����U�Mї��w�L�e\ܖ�A�'r B T!$.8�I��c�����Ww�=�F��7 �h@-l]}�3\����#���/u�U�j���I�B�k|�N�w%�`ʪk�h�޼��Ğ�<�2Ǔ��fGsG`lf�y�&r�p��P���
���YМB�s�Y����7p4z�$��9�wk:`j)�v�H�H-ŀW��$ʲ����ζz� mwf��3Q�R������U&��!�r$<��������E�Q��B��Ԕ�$K$��O�s��t�d�lY�Y����e�	�xY��	��������V�T�Rx93��ws��#J������$gK����.K6�mZ8��"�/�2u6�[�d�gNO�3��.�I�!�R�ݪ`�i����Y�:ǭ-�#Ƒ��zm�m�*�����v��0�*����-j:˨�#�BO�-�D�w+�����}�H�`:����}̝ӗ�B��V�Aq�G�T\C�F�yuq�R7$�0d͛-g�'������w&���g}�[A�h�н�+��O�*V8Ti��sVkW�c��K�ww�iͺq^&ZV&n�{�1�������u���6��6j�����aoq�oI��-&U�9K�8��������{I�tp�͘�9��`I��Y���&���u�$���{��3��C{���g�N<L��r��p�z�^f�0b��-�`z���Kz,V ��������;w�;��!��	��Z-d�lA�v3YCh�%�oh�Y�un���M���T�5vN��N���	�lT�����Rh�'�(Qi[ۭ�V�>=:�]�GM���Ç6Y�Z�V���ѶZ�!8H��-�'m0�ɭLpz�+�Ϗ���t���]:�4
f�z�F���DF���1	��\���RT�����q0xNtȈ�w�Ͽπ�I@�I	`�HIRI ,�,��B)$�������닸�R@RHE� 
B)(]GU�E]t]WQWtRB �$�P���		"���"� � ���@�������$�Y  �$�a�E�AeT]U���]wE]�	 , ��X�Qd *�*�ꊎ���I ���EXH@RI"���I(B,$�� �d"�H@P�� 
I$)$P!�)I"�I�E@��H�� (I$�@X (, �$�@R E��E��BC�$$ I5-���̬��g����n��su{��{���-A=-	�����贈��f"�Zl�Hn�`e	�x�����W&3�p�Y.�=���ynB����)�_��.����KN��q �W�*ɕɤf�yo{��Y�lԇ�7������wFL���������vf݋Y��;���f\�*��y(.磆Oh�1�Ї���g�������u��c���5�s�cG�h�x�n��
�t��&!���<��ީ��kj��`�SiR�o ������S����:P��$}�6��:|�������|�����zɩGzy׍�G�"gۼ�Zث~"��6s�k���f�v�m��\��P����ֆ�
�{��x��
oK�.�D��3��v��l�FE@���ʶ���\�o�&���ձO�$�~>�zL����P7"�K���\�;!���&
����qd����7V�p�y�����i�홼�`�{���26N;�������|�S�W�g��=L}N��L5�9F,'�M˓�4��fp8t�;u���;+d�ѫ�7I�����1N�g���$�~���q��{��,]��>��V���`�3�׾�˦Q���e��������~�Bx�<��jK�ءޏ��L=�7����1u��A/6I-���g�"���j�96O2�LReO�q�X�i=�i�;�4�P�F}�}�k˕��l;׷]#b�	�.�7#��!�oR�:��f�#�����;T���s�|�`����&B��Q��u ���T�+]H��׾yV�x?7�WG<��*B�Z��vxw9����9���R�C�v��-�Lل�W�.q�T�׾L8��� =����g'(jކl#�$9n��P����_���͊��79�*6Ԟ��g?yم{s�u�T�������Ӹ�ɳ�3�｝�sb�܏<��;���:E�G�x�k7sG�d��޴s����B�Q�7�{Q�X�}�I�._1N̳Q���>|.�L�qdW�!�����̊gf���g�[Π������:�v(!�B��A�#l�#��sAkã�he�+���$�j}�on]�A]�ty�͖ג��mk�
j�y�}�2�rQ�#DD�\[���J�"����L0�ǳ�j�=2h�D�m�GU�LbLs^�z!-Я���>�*���`^٧�|X}ő���=����*Gj�2_/,~7B�vQ��z�8Q�Rӆ���j��F*��9��kKИp��;�v줿v���Ρ�x�>�?����E�!���S��TVv���ΔNt��h�$�"�*2�/.���%<ж�ֺ�^�nm�w�&�YG;����,{�R"[�b�_��GN�?� �"�w �h߮m���=ث�uΘ��w�����{��WM�l���-�L�F��b����e��K���;R1�׮2���8_���!~�g�|q�[��!jv�*�y�(�sX�P��3 ��^�]��&}�G;N�D�UQ�I-���-�4�m<���p�>K�x�M�,Ӿqr�[���{�ΧJ����Y܃��ܩeB=J������ޞm%�~=�0�\�8�SJ=�P8z�^"t+�g���ІO�l2���B"���r���6x��ؖ����Te�M�莮��|���Vm�:���p��`9�k������j�l�拞v厲�����@��h�$��>��������k������<iEn�aۛ"���ZulL�b��@]�'w����=�k���ȥ�kg��k��W��o��<�qk�* G���\.��LH<L>.r����SaH��w��������(]��w��j�����J��ݢ���fy��~v�(��o;����\!�Yy��:��z�˞;��o�N���8���6ӳ�h�dFk��<G�v.��ǳع%�vNмl�	�����]w��w��D�J3�G�����5�@��������&�K����Cp�0zo�܄�>N����w[��{1ڏ��4x�Pݍ��+9z}OҾ6���x�ޑnz����ފ���⩋��a����n���N<����h�����kܸ���`bYOxYc&���Y��mx�{��:�BE{��zm�[��z�s��wd9�����c�@��t"}}�=5g��垃<��7iʡf��vr�1[�Y��l�L�xg2�pYa��9oy��w������uC���^���g ���/�7���ג�/OGa2f{ܔ��b�6�������ݢ���5���U���ڹ���^Թ��n�ۆ��V�.)�uXА���3p��(������א�;K��3^O<C�=��7.<d%	J]��s}��uO]jU�\���#�-���D;v�q<��qi_�T�9bܽ���VCr�Y�Jp�/$�Eg�װo�7O��;�5��*����)AE�fպ{Z[����w�5�+���1F��/,��Γ�و_g�=Ǿ@E���^���L��P�n�b*{��W釭Փ�Pk�xL.���tW�ķ;#�;�|���uMXy�,c:�LS�QB旇�9$C{ܳ���n4^,b�wF�b7��{��Ў�P�2{�S�@�}x����F1��-���ww��j7���>o:���>�o|��̈́ �n���)�t������Z@x��m�r�pd�P��۹�u�-�n�q^�O'�=���������v\[�ଋ�8�#�Z�Hw�2��F�3��??3�o{��6��pw������O���E{s`��V�ҌD5�*m� �����Csp�ZG�����L���x�w4��x^Udn��L'/!Ν�6J����� K$������>�:v2�{en����	Q���)�и�p4V٭D&��װw4��|��>{��o0N��]w;HIrY�f�}��xt5�^y抌���wW��}�ܛs���5���B���>=�F���7`.u�۴{س�R�&O�Շ=��w���͉:��Ψ��t�I"�E�R�/���4>��"z�w��:� E��0`~�K�J6�w�."]x�W��׿(p��4c��w�{d>R�9O�h�쏷#M��sQ�t�{<1�S�g=��l�Dâb�At}�aJ� ���p�����v��S�oN�H�3v(�;2�l1������u�����W:�:x�~G�n��8�Y��r��<u�6S��ӽ�do^�*�� �FS;�BU������|c��!O{V��y�Sӣ����{9gw.L�i��V{&6�ۺr7���.H��2��T����j{H@���{�3��i%�v��e�����k��X��SO��*X&ܳ6���R�1/o�P��f�v���U��ӎ/Y��Mdd�ʂ�Жag�LT�o��k�Y���|�({_�@e^�ܘ��	
�ě��܆ق��[�V2�D���]�1���(�)>����Nn�I�E��M0�i����AO̬���/G�\�ٺ$!����#I�p0�u߽�6?ey���#ϩ:xnnW��g������������k��j	;�Þ8;e���=�����n�V;�K���:����w���"���7.?{c3At��h>~�յ��^PF)�OYr��|5��&�����J�&���[$�y+}��m��c�o�Y�JͶ��e�(�_!�nC���x���N����؞� ��æ��:`��hP�'��q�o��]���g���YK��o��E���S�Y �����1��&��%U-iLz���2�[i�'�9��Ụ�jh��k�#Uw�]��APU�����~�s_��f����[�}�>{��l��We+u�ˇ��55��%��|%�h����^���๡�x��� �3w���G7�w��A�0b]�c�LG��9��=��S;Fނ)�QS&�'2��{�]�t��7��c��k���� �(f��ӱ��	)ئ�!]N�{��ԂG:�������u��(@/M���]��Y��\쾾^я�[Q��x�r��W/bC|�����p�1ǣ<k9��B�	X�Kz�Ι7�4R�	����r�������{8:ķ��0v˞\ǽ�OZ��{�^��f�(<�q/4���4)W����Æ�j�g$hKۻ�_{SΤs>�>Ʋ\�t3+��K�A��� \����y�>]�����\;7��k�am��|�{��^��\���jMx+{ņ��t�s��V�b'kn��Ѻ�;P!DUjp�A�3x��{v���=���>lh����E周�5G�z��#�7ħ��2ͅ�����\�s��b��ݳK{rPo�\�� ��ŉ(|OuD<J[Ȕo���ǎ!����E��l��12�e��gsM����%Vh���N��W���[����+�f駱��1�q<z^�������/��;J�@ ��������ֶ_^�Rc'klET,6��#�֔�p�`:���o���\>�{o���מ����r&���sZ�j	�/H�?>���;������u��h��vH�m¬oN��;�L��0n�]*��7��s���$��
���9�M�q�>��Ί���7<%\��#���/w,���d�Ut�X�}�-+���)���qѝ�q�����,�%�!=��zx�]{lR��ݠ���r �8�k7�+���;}�]^�n�=G �� Į�G�k�lj㚏��Y �m��wAb'�}���	@b��.C��݉	U\�@�L>:��6M]5{t@H�6���kW|���F�3��f�+���L&�Y�6�j���L�[���@�6P���*�e��Y5x	�ځ���q6�,��'��|��a����_R
�2#���*Q���u�|�s"��Ț��hK�ֆB��ڽ�{ޭ2��h�Q�K�x�x1����p�Baԅs=}���zjS����ɯ�r�[�
���3�ϔJJt5���~T�+a�غ�ޤ��UE�Mi<S�=��[��K��]|!8JH����x�M�`�'`�{Zw�-���K�G0����8�t�ސ�_�C�]<����x���A
�y��uM�9�=����~�X=}wH͎�=��z9x��p͜��GB&W���'Պ�*-���:��J�_{��Bz����	��l��n���c&�I��{�Wm��� ��iP�:�ae�����ċ��KPV.�|C�dz�K̻����� �s��v#��.g�s`]����I��:��v\9ʜ&BP�F������q~H:�CjdLɴ^��R�:�+F�.��se.���VF�΋��ٗy��;bJ��0�TW��_g���;P���2�%�G���f^:>�_#6�}4{�%�H�V�����,x�V�/C�\y���)cݙ�{�[!�������#ղ��k���3����t2v�5m�"�p�wy��"
xE``,��Ag6sTvq�����F�e�#r����)�	�j�����j���5����C&l�������<y^�^��/�}g�ב��^~Lk=������.=���<�F�;�nL� �w��c��O*Q��c6	��zGB�P^V�sCkz7��i]��!Zf5�z�[��D8�<S��
XQ�JmG=w��|P7�n�N���m�p��"�w!HX\�0�~5�q\@gެ����fޞ�ke����.�{$��j��������z��w��X���֟����Q�i�3��\�#�ú�yz��,����W&��؎Z���y3��ɶ�L�=��j���Zƻ0��Z��������8tѐ4�|k CJ�c�E��]���Ox��KwΟza�;�]������m��/�'_>�zm�R>���$��G���{�cqy�<��� ]&��mP���7M��������L%f�/'�0�3�7�Ԗǒ70��"C"ftVoca��0�JI���ծhM���jf�V��o5��y1�O�4�����3|�t�;�Ix���!�gޯ����9�ex���:��ϸ�:����c%I�Ҷ=lg�0�Ml�gt�8$��,�w/���f�A���p2���>ĭ�<aG9���&̶$�\G�+!�{rr�z���kԝ)�D� �CO���ά���[��pW��W���ny{<���D�ӏ�'jW�����cG8z/Y��JG
���e��=e���+y�T�ED�>�9��[�y��|�����?g��9�u�'\{��j����΀�������~�o���[G)��k�����!c9�-�I��ţC�÷r��
��<��p���
2r؏�m�`:���+:�f��rn{��{�=̯���;�˦�K�v\��~S")<G]���08���e[0h�V`ۮ��������M�K��xԉA��=<�SD�R����;ϊ��z���Px���E�y��c��)Ýy�j��:|��#�^�.ʻ��=�9|~>�چ�h6��gz�Y���s��i���~�$���F�{#0�/{r�W�Lcs���}O�p���"���x�k�[�p�:.VG3PK�P��~}�}�΁�����-�|�eGsg��.��w������7����Ѽ��h�/z��>�Pac�.? u]M�oOiu/w�>����h�!j��
�t�4B�����>�s��wul�o>���<T�;���h:��˦1��'�������~�A����L�E��w��ĞŹ�j�I$��l����7r0p�\k���8���+J���!J&{r���&I=�E���V�O�x!�K�/�E\z�yv���zC��(��;������v��U��!!I� ����N�X�����Y�Ct+��^r���inlԄn�%5qk\^������Ş`q���c֚=S�I�27N\s]��F�nD�1��/*us�'���k&��]�j�(b�Fn��;��{�ngi�Yi�q�;�Cv�Hvv[�n���yؚ˫��`�ځ��v:��b��-� :y�3�P��-`:�8�����A�c
kE��xՙ.w,�Kگ��Y<N��c����N{Z���.���Ć#4�ȬƼ�B��=���h��3�Ƶ�
lbE8�SV�Yy���6]�q֨�<Ju�^�:
ĲL"�oe;O-Sڜ����cm67�
�u�Ħ]4�sb*0+�˱JЖ6��ң�c:�GM��]�Xu<ŭ> �[u����m�T��=���"]����\��k+����x��ޙ��7
WX�L�kڸ��h��
-�Fq��0�ٖͤ���473GL/ >�K���n-��=�����F�C��wl��g�uEko.�YD���q���ƷJ�f��^����&�/���j�h9z۷	��ٿ�y奤<�n@����NŨ64֚S@n��.����`�s�Z�,�.Rk�]�zW�>��b��=�R��� [�])�4t���g�1H��IV]æ��m�Yi�h[,6z�ֲa��pF�m%�3==nw=nӸ�iŞ:z:���;^�����-�xŢy�^<g]�AeM�e��������g$K3��r��g��ֻ��[��-���;���y�Y	�.��P�fL�	�����$�"��W{yxb̵�b���j3�d���\�l�v�h�f�7F�-�aB=`�s�yI=���-06�F�
#)4*M3{K3��i��B:;Y�T)D�1U�t�Ɣ�Jꆠ�ILJ���R�9�����[���w:`u��vK�)!���4WZ�on _���š��"�y�gt����Qq,)T�S�m��"�p�IL�7YY]XFC�3Х�.�py[�[3E��׎�m�vZd�	Q,5e��v���66љT����/IK��[�ג
���I�v�\�Vх��rR�i7m��3Th+�Pұ ��`Y�@uڎ�!vu�&+��f9�R ����!uf� �v��2a+C�S=�G�әf
�t��7Mq��6m���a��&�ݸ�.�c �S����bۧ����x1����ٺU��n
�"�j:�1�1\=b:�0���٦�"Ʒ�������A�m�7 npt�V�xn�����v��\/=>��q�8mQ�z��	��[Q.�-�'�ԺD��>���}�=@}��ն7�����Em�h�����E�ǜk����.�'Vاe��,�nie�X���q�lƥ�m�'�)�ܖ���eZ���^�N�(�+�u>�v\���dR筡�N���s�wh�Q��e�@%���9ٱJ�<[�N�cڭHn[$�uMA#,,��z��$}s��k�Gs�v��^p*9	kp�[5�M/�<�4�x�|�~���4v}jp�ݣ���筦77����zŹ�ґ�M5��t)� �v{X��RB=��Q}���M�[j��&1�l[�%&��ƠP�8�����X�]@�ͬ�pd��6��2�q#���84-�4)e��m%��+�V�tn�v�cm#*���Sk,���{<�=���F+YW6�[��� 2�ىa���a#��9e�Ͷ2vX�C���RS�m8�i���m%�vz}�٠�t[�Ԓr�{�����:�VNz�כ����n����l�8��z�������^=�YNĜ�==��k�88���uoNQ�k�Ykn��@�wPD��#�Twg{nm�nd(�k�{M'�Bpf�I�D��X&]fB�Դ�#����2#�.���斛f�b�kal�����Fa1	v�y!�[\:�j%H�AM����*��#
����c��ӡd�֒��r��&̫�Sm�s�Vh��1^h���J�v	�ۆk�K�j�������]�3�V.��E�4Ж���mWK1س*$�e��뎬u���>NwSk]���s���������`��,�ydd�ka��L��(�]�ں��ͻga4��V�	�)AO5�0�&ٺrvKk۬^���ƙu�+Ÿ1^��p�j.�.��8�k�w�Ǵ��\���Ϸ^.{u� в� ֳ�5ф�x�fۜ��lh�3�:�qg��i}�g��{p�[�9�H:��k��f%G[���g`�8���rc��\������v^�g\�V�j��r	q�S��ơ����)�vy�bbՖQ�3]Vc:�Ae�����Օ�H��*E�nJ����0�S�ƎΈ݃�R�[cQ[�T	r�2+m��,έ���z����\�R�Ѯ��{F�v-�ϓa�8#��|&�R]�e㧳43^5vW�RX���^'�+ډ5;�V�t�v�8�YKb���n|6��F��xôc.�v_Q�Iѧ�Ln(���鳵Ȧ::4lM�i_�v�b��c�]mEW����x���S�:u��t.�h�Z�3=�.&[[A.���ҔXg�ãy��P��Z�Y�,���63�79���s�Bq�n��mtvKv)5e��E̔�4��\�Ġs������ҥրEn6)ncԪ�Ι��Xm�n�)� ���dN�+j�%g[v67<]���-ۭ9��hɺq5�=�r��F!��<s�ØvMR+�k���m�+�wY�K�4b����Yn��(��t�A���#�]�b�F��s��ۤ��(G-4���e����w#(��g.s��;a�����1�R$��[fR:�p7
�Ŷ0���a��� ]S�z��8ڙn�n�m�Hv,,�rKqXҺ��p���tl�<n�p�:ݺ^��+ɓ�s�^u� �[��b�z�f.���s�-�qE�b����g4�M,�V�:�[dA�kR�Lpmuc�E�Z��f�`94���l�
::fB��<p�V��$
�u�Ԧ�7;�q�z:�n������`��b�A��� �����B�M5*�H���4�د���xJ��GCέ�TY��܃�-�爒�Cб`��R;4�kUs����ė��GM��Q���ֲ����u��b��8m�z���Y�:^�D�j8�H3+f]-e�	��:;�7�ޞ'h�f� ���-��z�rb^#�D��`M�6�1W�^3�)m�34M�B5�K����Z�ܽs&fqɑ����l
����Z�^6&�wZ����ὒC%.��q(K���F�˩�g�{�xN8:�3�v����:fs�S��W7Q��t��d�\m����;Wn��۷M7gAʍ��=���p'�&�⹕��5l�`�s���"V��LR���x��cGm�8d�㝋{b�X6�a�[���R�Kx���$�<')��(�$���.�́u��h'[���S�H�X�	��MH��t3`{k��;M��IdU���&䇎����^!�v�y�X3	n�p�pr5�^�p�vy�V��I��J�'��Ngη*X�zz�N�
�&�lcu+�'\)�]����U�!}����v�+���5�n������\)͐Q� �(��`�k��6_X�/vy�g�1cV�e���lƚ��V�A�]����ã74��P�� \K�5�����)a�E��2B7g!�;Ys��j�n� #C:����k�� �2�SB���[k7Fۓ�4c�Kv�ږ��}�;E�I�b�ʹd��7��J-�ns/h'w�=V�@<�֋8��
d%T�ۣ��5B,K��Jl\��=��d�T��L9��,�h�;Z�"�6��c���e�ô�����"�Js���@��f���S[�;��{cve ��F)����۴��Vh�0����vy�`��ڨ�q�l2a�l=sҼ�%�N�I�҅�;�Su5u8�����n�3q۾~��4�%{l�u1X�JC=f��٪�]4i���p�"6'����f�LE�4�dW���(0e-w3�-�Uά��܎u���Oy�n_,:�]��P����a�Vxl�%Y��l�:����\���;��:Ռݣv��8��gsZ�z�m�#��\^;���Ҟ�r2�82lp�Ø=��Okv�0Q��q�)&NfX0���F�`���*XۧW bx��sE�-��C��^��R��^8h���RSxR=u�v,�)Q�Ӻ�t����Š���W;}�}��p�g�㓳�����CiB�ݐ�� ���^:ն��R�M[����jS�e��tm�n�7P"[�dܝpcY�ܜ�&Yݫ�ζy)��3���i�sY�.5\�%؇*n�{J����u<�p�r�ƺ8qc+rn˨�����}�S�8�:�F9]�Y�	m�kE�'������\k�{d��qÝ`�a���M�SRɳF�]7T��[q��`�;-\6�����U]ή�"n=<��$�ɜ���VU�A^@�j%�&�1P�Ĵε�h;��+����4��)�o1���7x��6ܣ^A��iю�6������t�ZP�Q#�C(^��d)����f6��*m�&��%�9:n�3sQ����拡H��'��q��X�h��I6�t1�i�[i�vn��z���R���/'u�
���$9��Ml���P�������mڜ�Oj�$��lk�N���+�Q��-�;��6��\�sU�l���g\�Q\8
1�l-�͑s	�5VPi��n�˅���b~&�vݱ�HY�cp�6��x���i�ˍ����nƓXꞼ��q��h�fI���=y�����C�9::�"NxZ�`��Q8J��8����Mkr[u�!D�����C�r
'	@�9�:�N����E�a���j��ENJij@BINff���$tBP�8��G)�f��q"�$����L�Yn�9!K�l�:p�sm.'#�������	�tu"Y��8�irSk��#�4	Ӝ��!�\R���m���F`I �țZ:qID�8�#� D�fVgȂ��q�1�$H!�D��IJID$�)�`D�-�����I�9�ĹHp[b��tN��s�ȁTR",��EQ�� Zd�arv9��k����78�n�NM�e�1�܄�نŬ�l*`�J��vG[�59�DK!�s����ꂎ	�gUKh��C��{Z21�u��T�� �-fvJ⚖�36�pp�!1�`��Cr�����p.]�n������s䇬H�F�	4v��q�^���%�a���x�(ݙŵFP�z4_���>��zWm<�V��y�"����r�8��Xi/`��l��:8}F3e'����=s)�T��ی�ƫ.���V,�m��c3+)\as)Q""��%�2	!M�4����cD,h4pئ�%�u�o��h{g����i+�FS�v�#��8�������6�=���/>:�u�'�r u��wg�Q�Ǚ�{rZ%�����GkP��t�:����s�99�q�T1]-�v8ܔ�{t�s�p��K��Y]Lm��/5!� e�9�b�"������ܬ��a�e*�[�v�N�^�,p2հ�5�MGiJ�oUù/E����.�n8��h�J��k���JД"=��P%]s��[Hn4ư��FmLM)h�t���e5$v4E�b�{{k�q<8�%��e�GfᴃHҽM����5��ꎬ��ݭu���P^���6��[F�<�Ѫ��bese
�t[a�$e�ɫu3-���)!f�k�]0�-�7g�=���Qk���Ѯ���[�"vmD��v��A�ƹn� 7n�/$ŉ5��hTlH��i�kW��\��v�K���)-�nNg36ݳe!�̯:�ۜf�C�a���جݢ)1K^��g\o#�c<1uЀ�v�Q��j+�X��*���
�M3�#��&�Vj� �͡bj.�P�1���4�JX���B�`Ϯ�U��	;�v�NN�<p:Tɒ1�F�0�n��
��M����rq��=�t�c=��U�ѹƮ�KOki�nL<����ct����x=��Z�K/]�Y�I��Y�.��wwwlݱ���A�Jy�e�ԖD�Xڠr%�)B�X���i)���$���4m��=m��[͋�qe%���p�xDvM�{�6@\�� h��KA��T�m��4X�B��F���lZ� �z�c)YV"�Q/6��zb�kE�%*�[I��|�#�A��<��2���	�˸e9�p�
�pӽ'n:m�X�Y��ctn����D���&��Ⱦ9ɜ�6�M�x�b�A�i��Gz�u�4A6}���|ۚ>pnE8�N%N���ϭ9<���Q���Fs�#��������ݸ���VY�sS~>���e�4��حW\���{y:��v�������"��"��6�܃�y�p�LT4#S�D7�!k�,N���Ƨ� ]�� 쬣�sV�t��w��9�k����"�MȢ���'qF�BghSÛ՛�*�:�h�J{#�}��(��W�,��l?LtF���#�B�A5i)��J�ֻQ�L^�k0�,6&i�[�-Й���'�W9�i[s�-����o2yY�v����t�����r,���l�܊�����Ȏɚ�׆/�Lgu���6���!i5�R��G@�{�I��ű�ʖn��͍�`���Ou9�wVafr�٨���ίW�dB�59��=��L\� �Κ ��͹��*�t��� �nE[t6A�@��yWF���*�s7K�R6^�)�
�3gm �^�Dۚ!^��WDi*'\�O�f���滻Viݼ�Vr��ў��M�H�6M�;'���7n�o�F[�^!�"�fmȠCo�Q����1��]Wc�c5�E�{<AH�۟P�9|�>��|�z�M����4˱siuD�Ԗc�tkZ��Շ��ccf�5�Rl�o}��y�2|����f6�Sg�挩�΁��1Nde\N7g]D����B��T"nk�[s^m���N2(��O�[=�{z\��Trm�ў��|
�^ ��B�f#����F޺�|�РGb�@��!�B���x�F^��*�<�����.�/�q�b�X<&�JG�E�#`_e����py㞹s����k���㎵�!j#P�1�"\�tw.�N7�m]�͌ב=���M:Dۚ�׏�;#m��5�(F�@�0AmЯ6q�nn���B�@G���n󫗆��n�Fk��<D۟Qm�K"m�����r,�R�_^�.3���x�g��+�@���l�܎��{��~=��|z�F!�uڍ�)z�mQs���
������\��P΍f��}��izY�� �:�tx�D%�PC�.��ٱ�p�ϙ(n�썬� ��AKf�%�4�܊NDI݋��1u,20ǁ�Ey����u���ahB���f>��m˹h�n��jb״�g6h�� �ϛs`��۝Ov�,���opy�NM�z3�G��Q>�C0A�@6�:���g@��'���
#�P�Y����<]Wc��-�S>���`�=-��,�k��A��-}Hk�{G���1GP�~��q�]���K��v6�z��ϑ�gv�*+<z{�����%�w��g�{���˲8�s���x8�[r(ۑ@�Zx&Ef��
��(oO�h������+�C>��mϨ�|%�6L��z<�hG�0)�]���Y�M�Tn{we3���6y�f:���.�݌z~�o���{��>6A-������6����B���!G�P�+0����A�����t(۪�`��zh_��B��!s�mm]�z�L��3����6� ��	mȢn�x�c�6�9ܓ1�w�l�gn!w]g��PW< �FvРCn�^%�6���Gb�s�}SS�as�����}��7����B���9�"�����tF_@�Ţ�`���+�6�Qǈ!�@6н�[N�Ϥ���A����a�[�&xA���"m�x�mʕ��3�b�.:5L���f���q����[w�DC�qUYklI���Ԥ��j�Ti��k�Ω{��Mۉr�W��?`�#h�'b��;�NE.�s�v�۫[�aM����3�1��yJMV��&͌6�Ś@��,�2w[��=e@÷n�����v�O\c�uc8�F��oq�n�c�����v2T�
��\�W6�X�$�*k�L��ܙާVvs�5q�.�q����^@�n���N�X��4�BWE���T.��:��!����ռ�f �!�ݒ]�����������Cl��Qp��n<������Y�B��ὦ%��k2��*���������0�8�<�(P	�۫6�V���u�Pj#:�w{��`�s�`��"<J��r�"��
�(u���`<�}@�9�7��66N�!uv�t�O�d�]�B�fp�9b�ڈohP!�Р�A���Ĳv���7R/CmuM��z�L�w�� ��͹�|ۚ>q �;��;���!y�G ��Re����5�p������`rv�k.�U�� +���Am�x��ۚ�� ��;e�۪�R(�ɭ�כ'{��y�W��㝒ޠ�Am�Ǫ=d%tD�������t=������<iz���&IG6B:#l4�#3BL�L���0F>�D6��"�j���=��z�L��LA� ��_�� ��׏�sG̈�-�C]`��o3^?���:5giI{tk|��{<Φߞ=���]�b��<��{�.䏴�p�=�C�b�z�[�r�z�P����	���L1N��U]@����Cn��cEmS�d@5{4A��٠A�6�� ���t�"��mY��\սN��{/�
��C0-�Cn�ezЂ�����г�j����x���cX�6��V�ոfg�A��S@�_N�M�(�(�t���8�6�Qͺ��`�"�:���L�N���S\(�A��x�s&��z�X�Uq�u��M�PӳաK�:��Kp�Z�۶�^ú�bh��kuК>����A<���t��>�ۚ���xu��&jާ��Ӛ��Fb�@�>�ۡD6�!� ���=G_n#�,����n�b���×z���>�S@@:|۔v�H�'���o��Q���AK�܄C>mȝZ�Q��99��6uW�<��j��zxYe�+�MqԶ��ޞ�+����1"�&ܞ��i�wٷ����� +�"A��
f_�ˢ����!WP �`q�
!�>�ϛs`�Y�(��͗��>�l�9�>�ۚ]�f�=X�Mnf�^��A��j��B��OBN���mP��B�m��,�[ٴ��:�j:���+U��33� ��4 �[sD۞�V����A��Wf��;��Y�":���'O ѫ4W�m���۫�;mk���������O~�;q��r+�}@3~6�$۸�vFpzS�AVxv9�4�%�(�ު��4|ۚm��8�D���D]4:��f���Um�^�	����f:f7�GT��VUϤ/�Л�D6�AdCƎ�U����9Y�r"g� �)�:D�׈>-���DI[m�����7�23���x�`n�H���L�d>ga1
�p! �y�P�%mT���#���)[��W:�\S�mb'��jWO��|sx��@�soO`:1k��Zк�Oq	w��3U!�׫�Ǐ�sd[s� ��ܦڗn�b��ښY�gv�V����t�gۗ#� ��^!�!�"���b��j�A34jA��wI�E��%�l1�u�k��۵8�n�s6�Z�����~�0�n�M�x�ȇ����o�*Õ��"&x�lD�Lf.��A(�k�X-��|Ȃې&�.XcfD�C0A��^i8ܸ��b,��cS\(���j��2���`�eϨ�4A�-��8�z�w]��Xi�(�N�k����(}��(�x�n�ۡC:M���0Y@�fЯ���k7g�]�+#/܈��	�SD+3�P�yIR�>ǲ� �ۑ@[t(͑0ټ���M
�����r��`[|65# �5m
!�>�ȑg����m�G1�9��(d�U�ٵHϟte�E�f_P�{����"�S��"����s=�։����/X�Jo�N�>�s�Jw:Ӿ�������z�7jktfb�Lѥ�e�V��YsAa,M��Eu�5ɚL�V���э����i12Ƿmdu�@v�eK��F�K���	��-�%Wc{c	�����Ok6���͐ƜqG>wEtv��ĽE�ۣ��D����qp�"Pq��q����3A�]�����u�c�E�F�v����Lua��F��X��m]C�276�O��B~+?�� .�	��eҵ�v3�E��[s��g(�����v1����|���l<[s@�[s��Z7���N�k��"���)8r�`#��W�� ��
!�T	�!�Vn�JuFn�x�D��z��ݲ�e�=Ff{��4A:Dx��9aߥ1b�wt u��(8�@���
!�!� ��N�ؘު�����{q����Mp�A�n���,��5�:����m���(O6��A)�����w��c�o5���{;$Q
bu�F��ۚ�8�A}�(��
�-�� �9���կ�g�l���[�{�8s/1�33� ��5�:Dx��A-��G�d���/���Dɑ4dT����v�8]ureB=f���=���L��W��-��"�>Z�W�f  ��RM�e�'����l&2k�ͱُmj9#K �;hQ��x�Yn}@��E�l������s$_;�Rp�U�������e��;��.�3���ʩ8.��u5}�r��af�t�T���-�k*�#��"R�j4�d�ʞ ���]{ۇ�yF0jvֺ^��NvH��+�3՛��kZ��c^����
y���9�۪���c��{{ ����V���9�����|�"�nk�͹��3�����n�F��B�� �ۡM�w,�g`ŧ�c4d�P�"nm�$���$
��^'H�۟Qm�AdG�nU���4k���`F�&�_.ý���3;k]/_@';$Q�"���C��f9���Y��Oo�˳���774q�[�.��1+�������5�C���^�}�Y}|��Bt(De��+����y�Y�� ���jn��q���p�{f��nh�Ǆ�[r(���B�{�lQ`^��z��"�E��ahɮ�HF9�B�m�[4���X�7 A���9� ���� ���@6t�p�d33�4n��a�ѣ��f�:s*�8i�0����V([�y����dW{i��d�z��5o��W��nl����ʤ d/�M��}~���v�m�ѕ7�q��I����hd`v�k�����X8���3����ׇ�?Y�!r��y�J`�����6Ұce����7t�5S��ֻ��&�x�Iļ�Sp��O/�LS�&"���g7�y���>"|�vT�y�)�+��g��?M��Nw����/��%ы���R�rbSޤ�lf��#hjUj�����ѝ�͗#�d��{ý�j����]�+�R�����w����;l�(`>w_��Â�=Vze$���"Wr��=7�uV(��s]�X�m�J`d�LKئ�����(�R�9m���i��3�ȍ�x{��sf��(���8�>6�GL�u1xN��>Yox���i�=�2�����>�~������w���_v˾�ni��.ʳŵe"Oe3�绰�C��>�s�i����9�'�B�P$F�o����r�/G�8�<��r�'�����^�V����A��<ϗ���]��k�"T��"�m�/��lS�����r��x ԣo/ay{W�ٞ�����N) ]�,��B�Ľ���5���L)��n77j���p[��K{5B��	)�y��^�SS�%�E�̅u�,�+�9i��\��<���p@ s��^��}V���P绹��3T��lY~�t��[�-��2���s�Dx��¶u����sγ�6ݝd�6쎤��e��fS�� vQ�I#7N QN�p3'vڎf�8@���"t�-�.R\I':���2Ї(s�
�s�����s+e���г����䋎r�� 脜��s�%ed�ȅ���E��N�I$�$� �Ƞ�(!�s�$��Pm�.��r⸎��m�GT$A�Vk-;l��(�%6�ͱ;���6�q�sn�!ˎ99:;�+(�,�]ecm39�!q�tڬ�㤖݇QE[nJ�h�Fڌó�)��݉$q[`���J٫..B�.#�b	b��j��{����~�xL���K��9�"�#��P!� �ۡ@۪�Ϋ�G&=X �J��P�2��Vz�{`fe�=ff}��M<�͝��$p7]4A-l����܄gl!#����\��k�e�.4���lf���(B>�{B�!�U�Y�rWS��XP��TT�&$G:�M\u�Hj�M����u��{L첗]	�3���}�����Knh{�{Fwnt<&f�[�,��X$�Vk���wm
:DCn�m�@�DoZ�-�����:=�o�Y�}�FV^c�fg�&�O�tzm�F�v����w4B>��D�
�dG�>��H��uc]�.i���5#�QAǴ+�6���znhD���
a�Ԣ���4 ����������n�(Y�	��G ��(CBF���cd�S����6q���L^z������˲�h�i�!=;9W51i��Jl`����R;�p�9�Y�Ĥg9�0Ns� ��*�kf�`tz��+�O����M���Ȓ4�
J}@�t�K"Ln�
������>� �L�=���fU����\&�ɴ���=,��Ƌ�˫O?�A�r���`� �n��ӖU8	�ح5!�f˸ۤH=ڨ怯3��m�|[s@�[ب��я���Ϩ��C���s͌�fku�B�x�o�Ex���+ő���&��Q���mТu��=�F��ܫ�ڼ�ٸ}��\��}�w~"1׷x��Js���9˜g���ܣ�3�` �*�`�t)���N��|6+B��@���+z��s�j���+�}�4A-���nl9�h�N�rnk�;�盓�&ku�B�7}"���B�Yt3z6�M���������z/x�"���
�feAuh�m�/�a�/�Mv���j��[�Ƕ^�׻<s��+ �8��	'��n�ೡ��;q$@_0,(�X�Ź��yFǁ�ٸ����[���q�q�u��3[nu �ډ(i�0WZ
G���d�'gYk.�8,�Nae��N��p+�xp�W6e�n��Lv��>\>V��6ݷZL�V�Ю��n0ۢ�X�=e�����D5l�����aW�9��6h�n�<j�	=6��;�z���h���=��e�����֗WJ�����سg�k1i��"�1T�ΰ+l+ m,S:%��,�ki�Ϟ��[��Yg��(��
�>��v�җ��Z��z�L�����)ɚ��׵]<>��x��� [sD3�-�F	6ۂŵ�PUpg���Si�����lV�5#�DR'���87T<��f̩Q�j��s���4>-��F�{j;��pn�^nodwnnK3[�����W�(���(�n�x��
lm�e�O#���B�z�W�,�	��UM��J�1�13����"S٬�����>���x��y�"��@3Cg*��}k�^�����t6��1Z�z�#f�
6����!팼�7�a��0.�J�±�P�D&��lH��"�-ˀ*E�da�1U�,��f����m�-�����/e�����zȬ�8.%��'{�#H=��x�}�B��C>��j*�u+mn6nݕuA���qHZ����F�@��5w�!㌸W������Z��5=�z�=��������-�#g�j��-P��}>�x�����j�O�
mc�bdܞ �"nE+��������1��^�/��0D�9�D�B-�:	ݎ��ӎ�m��N��؊Ц��# �� �^�Y[s@����!����o�����nkoU��ngK3[�ez�@>7}"�#\˪<9>
��Ƒf>�t(ۡ@3�mТor(� W���//mWFLr6�ꈙ�A��SG�D۟P-�M�V���<����K�jE�vĺ5�e�h�X�ܪ�;�Ө�3҅��6�C����[�|d�~|�x�`�t)��6�]ح��v"�)������b�5��,�-��-��D5
2	i��A���UwOS͆*f�V���j�E}��(ɱyc�\v�+�
jڠA`@mТr_�<���{xǁ�&~��H�F�Ws�.��!�;N�s��;�.�O^�͙b���֜��L�`*,[8n�Ik�W��Z�`�Uq7�1J~��gd��[����6��12�O����[s^ �ۚ>q�_��4@�Y�:@Z�
i�n�&�㫗v+h�݊�
/�F�1J��R��{B�����ۚȀnH'��v��{SJҾ���c&kul�_z��>����6�D87����at�iɍ�"�~e�{�wn�r2�9=�Zѧ\���=q\n..y��VdG}#�>0F}�(��W�d@��cZy.�2b�ZǨ��/�&��R�(3csqj� ��s�hAm�8�܁t�������y��F�CݑA6��ʹ��\\�q}@��sv�|���Զ�����v��۹��r�E�P�[s]W��.*��>��a�3[�ez�=W�(���Am��
{\��רp�M�ȣ��u��|�dBݍi��ɋ�+�<Ar��Z���]�J��ÔQ޻�˟�l��8��PK���s�he8������`h�Z�sh�ޛQr\m+�N���	�>~�nd~�r�Zr(��� �F}�3T|r�>�A��ZQ�0^�K�ѱ]�� �}B�!�U�dOd,�����e��Ԋ$H�g�l��5�4͹�p��J5r���Z㳮�v���/��4'H�[s��4^�=�۝���ݗ���t�{M\�`rT(�<Am���=F�u_v��ڠ8���֞L�91}ec�bg��MO-���|z�}CA�ɡ�� ��9A�n�g�ۡ�y>����Hmv;��F�{�F�p�|C>��^!�^�"<[s�g^T�Q�|�2 ��@KNg�Bގ���fkq�YgH�G_M���&����3�q����t(�6�Q���]ӎ��{�a����2������Q���:}G��nh�[s�ܘ�ܗ���Z�:fp�o��������/3�yVl���B+M��Z�Tjgt�3{{�`��7H(��[X�0I-�]���F*�g��y����'I$W��Eئm�/g�aQ��4g�/�[D
gg$S�9u�]\��p���t����lM�#�J��`������]ە�<[��ύ�B�
�Y�F�$燂W��&vۄ��U��ԇ�\m��f���Y�ӗ�� �Fc�Y�J U%����T����Wkhg��Ge(rn3���ls�!gow6�Ǘ��@	{�>ͳ���WfN	xu�j������av��C&�d2cv�kX�b�&��i��pdݟGH3�%P��[�uȯ��P�� ��B��z��җS�u:6*E�M�nzWzf�5���;"�!=�^#S��,�� 6�Z1@AdI�s^ ���
��[�۝��n=��� �ΑDwt���f��P,KT(�K�Q�s��s2/�Gh��~,�q�����;�l����Q��>\��A<Dx��%�4|�C3��X��r0^�F�� ��&�_)�2���i��ة�_M����!f�E��換s@2 ��z�Uwh&^M
���{�tk35��_��Y�(�wP� ��N��0�:��dUUDF��])3v�9���]�6�l�=�t�����;%
�a�A��ۯW�,���j�Iܙ��i�1S홑��a<٩�A��s�}^-�؀KnE DY���C�f��%T������Y�{���j=G���t!���-n�S§��=nR<G~c��薝^��{�b{F�7��O^4�&"R����wC��
�I�y��:WΖөѱ\(�A;�Q����5��z��3��Jsׂ#����*<�P-�����mӳ�Sv{Z��fks}�|���`�����Ns�b6�P�LgVY��B�"�ʲ�x�[>���kn��ܙ��i�1S��Mx)Y7�67�Jk��vh�`�m���0�}���F֌b}�f�����/#�-�S�b�W���B�Cn����O��ߩ��{��MXA5�1X�'j�`e�9�s�;�؝.�P���2��	��_�e���h����mϨ��4�V�|�u���[,Y�B��{uP-go(ʐ�;�B�� [t(۪� ��sl�弰��f�V ��+�8����˓�3u��ꈩ�r�q�*������`Q�S@�0|�dW�>mי-��݅d��&���{W���^�י���4�NM	[�oLmXb35��G7
��R7Z�3����)�y�suF8�X�ϼ������s&+�t��S�b���"�mЯ8�۟b�h���Yҧ��.�r������ծbkql�g�>��ob��{�+/�d��P6�P%�6�Q�Q��lc�S���v^=q.Od��[�"��^t� ��@-��A�0�s����P�&A�f���6�cbh����C��R�c3����pݓk'Dײ(�B�"mȡ�мw�S[9Ҷ]N���E���;��"�>�t(����܀ۖB�]��10U��>�f�h��Ӛ�����V���ŲŞ�x�t�[�B�!���YS5�_)�����@�@��
6����9'Ғ��ww�[*�8ژ왛�ku���5�G����A-���b0�\�hΧ�3L��t��ۡ��w��N�9l:���(�@"�b����#�%D�nmTL�GT<jc�2��R�������"{A��͟m`����t��t%��w�`@���lp<���a��s��u|�BHI�������<�q� A-���[sk��P��x�A���k��]z�&��x�r�Ewz�xD A��#��8���\O�H����M�y��he���Whgn�踮ݺ��y�ՔF����"�(��z�Ϡ6^|�:�ܙ��ku��*��}sgz"�,תx��Ao��%�>f�A�m�
��շ^�T��<D{z�{�����m�r�u:O
� �9u
6�	������yd+'�q���s��"�$6�`AΛ]	��s3[�e�>��(���̋6�W�mР�����j���r�D>�����nLnLM��T��%�M�z�P�Q����!� �[r(�u�C��ެ�}��f:�Fv;��������C�����G�u
6�\y�]i�w�+�3�
��)����
fx�dur�Q5����p{ް3F;糯uӺ���t�]�O�'к�;�AR��' ��]5�~:w�!��ܻ�`�!����iǀ���.����\8"5�{  /U�zg�x�<oo�S��� ����x%wX��=���O�z6��ΧC�A��#�̓=��2{̏l��/�+Jզ���݆
���%��=ˏ�
�{�;�0�n��	�Th�q-�j�jb.�]`��s���>y��&{�WJ�K<T&)�a�\���FP���f�cU�k���	���r�w;�� Fȏ��n�hS�|M�i9�c��xk�X�g���jvn�4G=��K�A��)�y�K��|<�n�gy��y�h�f�9:vR��R]�?M�z+8�g����e��Z��s�7�m�w�u綾{ o���<�N���˼;��F6�h
�e�9ʣWn��O2d�ɡO+���b�D�ok����k���^�r<��E�1�=�Cu�s�xz�/m3��3#Nh�o#�D^,�A�%b����)�Q�?rI��{�cv��v���)��%5��Bj��O	��S��r?f��$ Ƚ��JgE}vR��g���.��w��6G:`K#NW��|��V|~�}3^}٢��=��6�'][����Y¿vr]���yG��>&j������caFy��f(njw_g�g��$n�}R�4;���U	"ނxz�Tkع����[:7u�oE��� �]�VhNo�u��Jr���nq�TRI�A%tT�qE�q@�%�Ӈ9�DTBI�	��w�TI�G@�tHtwEpE��U�%E�E%qwQGGwNwTu$�QD�w!�w(q�t�uArtG�qu\tp'A�t�w'�q�GI%Dw)�"wGqI�u��E�q��Ew$�R\t�twT\E�DQ�EE�!�U"�t�Qqtu�Q�%E�=^U�<m����ǋэ�.z�"�rݖcpnm�5��=uk��/qx|��e��ēj=�gA����L`a�����0��Śx��i֔���m� ��(��$�du�T%Ѕ��S�:�����UW&<p����x�z�X!��m��*]
��n"L�`�M�wbRM�1�0'cۮ����N�М�ư���*�v�ǡ�$���,�90���(� ���mƜ�[̹�Ķdu��3fZK'S�q�����{%�����Զ�c
X�;cYi(������f��y�h"�`%�m�ub�%�ّH�]s�b��b-��紌����y��$�ׇ5�5�9������v�M�ОR҄\����D�,���x%j��[׋v{OB��L��u���)����}��8�ѩ!M[��vM]��ø��S��~'����Ԭd�Q�o	mA۶�6x*Y�x-�.<�^z7k�q�m3��\��)�kت<L�mq������&��v�X�mlP�V�"͙�^G N7��g1����&ѫZ9]��$}q;�\<;n�m+��SH۠Թ�-�:9�#]�:��Ÿ\M��z��nN� �&&��^v�[�d:і�*H�-��2M� ��}�K���:06&�f���n�Bj��xx���sSgE:���!�L^��`�S���0�n��g^5�.�m]0�UH���v!-,�ޖ���04s>��/;�T	�b�sx��ln��"������� �����6f��YS�%4n%�2�`��,��#��&��hL�5�k�a��v8�Ve�PgOn��Jbڼd�O`�W��<nKte�7@��hR��[�!���}d�v8�v꓎rmv�
s6�V2m�o���6�SD��'QXw��ݴ�����Gmdm�ml�9K����vl��F�DgX¥Zmț�`���oG ��淎�=Pcmq����������'I;�WO<B�Ӎf�n�]��;6�z��il�pe�O�Z�sI�:�уuЮ�:��,14-C;R;Z�IWa��Դ�M�)��C������XS+]wFRh���h�s>��K;b���K�6NBObKY���#��m�PuB[��f��6���#9j=��,�99��u�E�D��(���7d��6����l�9Lى����y�y �k�ҍ��\�Ԫ/�V�r�]���;���0&\�~nk��Am�6恮�M�vu뙚�Q�Y�Dm���o�q<}��� rT("  ��Q��D:r*Q��U�+,�W��O9�u1�bo���r��:=�<nT�����x��o�˚!�@/�@m�E�ۡ�@��h@�tt=�ɪ畓�u�hu3�#�<��t+�Ǡ��#�V��SݸR�} ���ۚ5�)��νs5[�5�>���@�	�z���Oe �ϨQ��D��^!�U�2���a��Ĝ:5�"o���s��:hz m͟6�Wz{�?l�]:^���səS��Hlux֬�eZ6�}���]�Y�'���̈�}�<J��1ȵ-��˚ᮣC��(c�{��n}�`a��0�5�{��2nlKnk�Q{�-�q��d'Z���&W���٫�U.W�.:�U�ܷ�{/�Խ6!̕����\�t�_zd����R	�x�C�7ނ�u٧C���� v��k� ���F�ei�{:u�Un(�� g:E^�
��3��y
��t(3@��nE�u^.=W���;4Lytn�bX�&��{�<As��G��揚s�l�*yG_Dc�7KƩ���G��CnEx'"԰��e�WuT�H����Abb�(p#�����[sD[s��sl�3�3M0TTH`�٠k���_gN�����<}9�(|��P��
HU�g���^l�33*���SU*�kޭ&܌m-�ܐjkfJm+-��+�hs���f�=��~!�>�I�n8�+As}%n�E�D��3�8A����^>mϙ�|ۑD`��'���Oe��x� ���V9����&j�k���xP �A�B�Cn3��l}�C���"=��yA�r��vϹ�iDa�^=�&�#w�){yA�:3�1:1{Q���}������}`�+��B{�O��i���z�=��?x�*���N�
�1AY��>�xxxu�Y���5;x�XG�	��A{�(@��
!�B�(�e����{<��A��Cݡ^>q�M�'�h97�S܈���3�&�b����^�=A��B0A)@�R(�%���9;xq���H�,D�}S�]ƇS#�x��ޠj�|���*K�Jg���3�~5�v�լl3ƍ�	Gj��QK)
M�w�f�ݕ�����w����*9�ȋ�rk£uN��d>f�o���H�UDLft�#s�Q�6���K"�w's�Um#���ǡ6�8tkAɾ��p��N� �>�ې�������k�m"���"!�s��9�d��w�X��S�2�C���48��#ٽ@6�y�@-���*��a��M�S�������A�5Q���_d>u��:�>�9�+����N��o��@cc�]�->���`�fr�{spo��o�c:��^��<P���7vw�-\��w��o� o7���J>��u�ő |۠s4���`��u�wgB�����J{�.{��}]�[s@��ۛ�p�Ӹ�@��1ޡ0`̮��\$������ Yu\�1�q@5��t%�TO ml�#��@� �t('"Ӣ��]�wW^����9�嘸�(�3���k����[s^>m�^�D��W����A/vhTn�������֠ϸΐt���bI�^7B�!�W�>mТt+��7m�,ʊ�]**�]5�M��\��>/���=-��%�4C0�3��(B[^�,�ۡA9�T�nnxk��⺁��B}�J�y�z��܊���{O���A-���zm�p^d\��f�F���>Nz\m^m4� �t�!�O��r.����^nK��-��f�M�ٷz�i�s�o�!d��J�'n=���ې=��)Q��	���B��}��ې�)bz��Ws��I\�5:�{�ީnP�13BQ�HV��vq���6��zF��]=�9J�<�X�^�W�&Gg�AAt��=�q�h�;[�$�b*��f�5C$a��g�E�1�q���s�qwgp��M�]�����̛7w%u�:HJǨt��ncuhY�ە���n>���h瀹���볺���!e��Fbh��Y���gY�I���b��n5Ό۲Ctt���PƧ�������Ƈ��c�+��mwcv�*b �����h�vyAmn��	~
��@ ��B���8�6�|�rn4*���ዞ��B{�u:��]8A���Ϩ���� �ۑDa��K�C*�a�;��"�N�E+�諞h�q\(x� �u
!�N��¢/z�9h>ۏ@;�>�yl� �Ǡ��>m��5�{m�u*����ͦ�<}9�(_u
,� ��
6��&������jܐ5�Я��W�=����&�B����"2x>S@���c�z}eu�-l����W�!�B�!Dn����(V���CyvtU�['C��(�G�>�(۪�>�������;��~7�lWUօA6+�v�6�m���y^(�Z�)�i���~���l�ￎ�/�F�� ���C�=y��^����ϲ�3�M徐���q�B�!�B�,�#�4�����m"Tҽ�mX��}�kN���'���7��:R�Pߙ�C������A7�Q��ogT�x-�D�����=�t/���:�>�BmG�Óq�W�q=Ȍ�>|����[s3��4��戳�;�ECn�Dr��3|2x�Q�Z��h�жN�Y�|�����'9˘r�9ˏ���j��pݎ�U3��:= �t�ۚT�-�,p{W�O<A���G+ִ:2�<�f�ȀA�����Ȁ-���$��W�6�*w�����qi9���+���"2xA|��=�[s^ �ܱ�/d��Wf�&U&hCn��9��^�É"R��6��C�+<h���� ��r(���́~mР��i<��q|����r�ȼ�+}!" ���P#y׫�8�x��ŷ4�N��=��y��d׈ �٪��yN��8=�ͧ��p9]"�/�� Y4�o/�O�K�@��^	�n@m��=%��S�gv?���\}���A����Kx��˵��S!�z�ַK;���O(�OMv���9�?b�pd���s�| ��������ɕ��{� -�����-��۟3�3x�c���#k�"  ��
N[0�<����gd�q}@�"
D��y��\�x�ޟS�s`��4C>�ەbY�{k�[�]:W(����y��3� �9�(���́a�B�����Ҥ�U�)��3"j�Ȣ����II�Mm���sq��u��kq�D�G��u � �����>a������\'�b�#n0n�!�Ω���x��@��ۚ!�ɹ�u���"�I���QG'"����y{�+������<DZ��Kr�l��}�:�_�(��}G� �} ��ŷ.5u �؉rSP�s�f���	���EȀ-��=��8�>��F�^���4y☋���Or#'� �)�E�3���@����S2�I��3�����.�7�+�F󽸟�9�f�]d�ʖw8�ާ/��
/#be8B�m�'�=�l{��'�ޚ!�[r(�t(�(cv�7g��@��+ݳ�.��ܸ�\6���<@��P�ۡ^gװ������ݵ�����k:�ܕvC�x/6�5��4YYA.Ρ�6�ɗv^-^e�˾"���*<�/@[sT�J����36�x���nOM�T�R�N�Dn�ۡ^d@"ov�zE�;F:�q��:�&oD��q=ȋ� �w���=-����R%��4vO��'Ȣn�Dx�۠��/O�����n�v���E��t8���t��u�} ��	F�J�N+�������M�Am̸һ#as�f���x�WHqN7�.��F��>k�W�i�YmȢw�\t�+c��=ã��E�M�߇����j��{�בz���� w��4���L��{`b~漵G�WH�����ŕ`�n��&�ɦ2�}��{{6��z�ѫ&��!مz�"�R~�jS���.{���h���{�wC�߾�I�r,0��Y�[���#��E.l�r�a�p�hF.��3]Msqfc�]݋�;Z�h\s�/��Eכ�v����iz7n�OG��	˫ˍ�W/�	G�-���90ca�'���p�޸Ѓ�N�U�oU��]��|%��7c�礎�q�la�y�[��뇛v�n����.]l�e&�G&�P������K�@q7�>�'���E�hA��b��V�w[�n�4�Q��b��I�J̆����oD$�IK:T�U��f$Q�I>�lH)�
aڨ,���
�{�4�X_���ܿ��rW�h���x7*@��dAd��e�_��}U�����[��4�Xi ���Z�
Ai�AH)�혟�$P�I����4$�����}������M��׾��R`� g=f2he$Je'9��Q X��/펅������|6#�H)��޾��$ﾰ1 ���v�>���ݻ�Y�nJH(q��4�Xi�$�ܰ�CI��S���[) �Q��$��S�큉 ��v�
AM����yM�j�v�c�	��R�q=� �o���$P�I�`bII��PR
K���bAH,�I����	I�j�����{O~��p�}f$�������$�0��,d���!���$���ꗹ}u��G�#�����$���,�2�
s����g<k�����z��䂐R
{۰;5D���)-�;�ى��I��I���Ă�Xk�pR
KB�;�ٌ���+�{�w�������R'�F���U�y�B������G�aڠ������7��Ă�`RAJ;���
h)�j�����w��I����M�Օ�.���QT��-�P����P�DeM���&d�3=����<��YF5�bAK����i �ʨ,��H(s�bA`i����lj�)�!ۨ).s��;å��f�O~ 2 ��G�#��^#J�+�vt�i>�X��RAa_]�H)�����2�%��{`b���AH)*��{f$L
H$T}3.�c�W����3q+�U����yVpX�]�{gL��Y
pDZ�Ģ�⍙^���X�B�d�Y���q��<�}��~��X��դx�~	!![��$� S�Ae�RA@���bA`�;���_�q���m�8�Fʐ> ZAd����,��H(;�a�����AN����y�.��� ���
AH(׬��@���S����4��
;w ���c'�e$JRw��1����˙g��"�*�>��k;������O���
B�����H.�$�߾�4�R�Ag��I�혐R
AN���i �:޻�o��/s�0��ٌ;U��) �Q��$�I;����
Aj!ۨ)D��k&�U/���� 	��D|@) ��)=�,H)�t���s6R淫����)|�f2i��Y(e'��4��Xv�
AH(�lĂ�R
~��p$�@���͛�z���W��O$1k�i<	�)����_M�b����È�$l��4�Y)���,�2�
w��I���
w��4j�)�;u��8΁+D�bL�s�f"&�;R�I�k�f���F���An��ũ���3Y���I ��큉 ��z�
AIb����H)��}n�(�/׿X89�1�:��H,;U �3����������fY������}�`H)�
a�T[%$(C��H,5RAN���i �P�`��L��H(�f}�g�i�[��y��H,F�
o��4j�)�
�B�
_{�W=åk�f��� U���@��ʌ����!���XQ_\) ��
@�{f2^����m���o�����R}�� i) �yAci �o�Y��`RAJ;��H)��L�) �,C��H,����p��q9�Ϩ���-u���5�U۽�&s��ޅG�eվ)�|�?P"ln�+��(����h�8|0ٛ���ψֽ�����"���o!���n�{��}M�q���b�\�<�-���be�oE����K��3zs�+��Uϲ��6y�y�{t  b|� z���ws;~��;�Ȯ,]��'yy,��w_@���gsg!�
�Ws�pZRB{�;�s��܄[�	��$�{�-���z�E������{V^��R٭nA��lꨙ3��4�4��ê>i�Qԛᩊ�|mޙ�7p��K4�.�`5�t�'m�զD)ۨ�:�^�s����^֫��"��\�Ӳ���X�1��hi����U�w�;���n�:h�<^Mr�Z[t�̀͵��Gn�y����(�ջ��,��ͻ��dA/_;�Z��!�},{�_����ق����<{;L�����H��jW�7���/��a�R��c
d[3�5ÞE^?XXo���Id�v��M��tf�\K_��~��}����s!XNI�Rz)��Gv��1�@�Ωn�w�<��;x5��2]k\l����=�{t���>����i38��9�H�7rf}b&a[�jm�@[��'-�	:o�_�޺�B��Og�#��k[�w�>�v�[�f�|4�7���Q���/ܩ�ۇ'�]}����i
�[}ط��������DH9�#�9nx�Ć���p0�.�*X��l;;���(�肭_l]{J\�����;��;_���^�2��/w_��AVA@DP]�pQ�q�G�PEp�uIQ�ԝ��qt'P�ˊ�[k��;#8�N(�*K����8�:r�γ��2)*N ��컵���TTqED�q��	�tq�GGt\\ugZqqA�\]�'eeGQ�QG�.#���#�8�$+��;���).S�����*8�-,��$˻$��[SZv��pq�QG;k��E��X�6�ʪ��0��%!�^�]�2������q�H)�݇�$Je0~�S%�������H,F�
w��5� ��+�
H)b w��
Af�s��~�e�$�k^�1$����B�
K�R��1�L���F������>���V�O�#�`����
B��3��bAt0) ���~�\�쯻�_��AM S�2�) �Hs�Y���R
w���CI��L�)��) �W{�4�R
AN��_w���Z�=����RhW*�R������t�x������
��b|�I��I�}`b��X?T) ��
@�{f2i���A��� � _|>����g��w�f���7m+�D�L�\�����;jn����7BawycX�a�) �yA��
B�P��1 �`RAJ9�$���B����
�{f���/���o_���ANo,>�Ad���}ϯ�z~�V�p����R
�?{$��
}��Q �{P���P;�ى��)���큈hII�f�~.������o�\סI �f�Y� �q��}�4k�k�ݷ��p��w�o9�Ă��B�
C�3��bAu�S���Ă�@�j����3}��������P/;f$�) ���
A`��L��RA@�{f$��
w��5� ��
�B�
}�]v�\:e����`�C�U̔�� d�(�G�ϙ)=ϬCI) ��_\) ��)��ɡ��Y*��{`b���6�R>�k��S�����Ă��I(��`H)�
`��L���
�{f�����r�g����t�H)���H,�L��l�������חZ��?}��^�K2�?��uR$8�[��*��Zf��z�����G�j4{����e���o_�gS]/��\{�͝�@	'�>:�R
AN���TAH-D+�P��� R{�14�I��I���Ă�X=�RAI�
@�{f2s�~-N�ܲ��x�Q�U� � ������w�����|q �{P���P/^��`RAJ9�$ЁL�)��I
�{f���~�y�z���USC̱-�m$[�dld��>x���'[r�^D����3�� �s���AH,T)��RA@���H,$�{`jj�)��AH)z�8�4Ga����߀�"rE�	�����g��ޯI�ֽ`b���XT��
AI`� }Ϭ�M���C);������õAcI!P��혐]0) ���{�W+��������>H)�����JH(T@l�#�����F�f,�m���<	�X}�AH,>���R
��I���
w��0��o9���)ȇ�PR
\@�}�14 RAH)Ͼ�1$��»w ��)��ɨ�H,�I����u����u��^�F7F�O�#����I!AT�}f$Q�I(��4�R�Agᒒ
{�1 ��aI;��hCI�]tw��~7_�ru�꠲xI��{$�I;߬H)�����oS���3�a��  L�#��I�2R}ϬCQ%$��s���~������R���ɦRAd�Rsݰ1 ���$�P�lĂ�0) �w��4�SHõPY����;�~�vJH(�Y�x�j+��WVb_
���#����� ��TO�I���i �44�S�큭Q ��T���}����������xvg	�RƝ����^�V�(�Uk�U�T^un�@�EaJ�/�fK:�W=b��o�v�ۇM�A5sg/%`�v�c"V��ͽ;�	 B��|Qy�X].��r6��$���X�ud�z5Ƙ9��ܯ��t�qc���p�2e����-���.�8ێ%�)-m�F�b)���(6j�Nظ��.rn&�0��cAu����u���gՠ5[��H��pk�и��Dk,n��r�H���jd"F�x,�+J�Aoa5�\�li�Y�X���٬�d��Ba��n��u�����ؕb �G;qG%�֜��j�R���!GE�U#��O�B�7��� RAe2Ro��1	) ���
AIhR{�1�Q���G���ݐoS?9����j�H,;U �;��5ϱ����H) ����H)��3��I
�{f�) �;�&�S�
d��H(���~�>>��:�X�I>���Q L#���<	ձ�h�9��0�߀@��f'��(d���X����XT���RX� w��;�����v�>Ϗ�$M�R}���Rt������9�Y� ��{`bAH,�)����P��{�G�>���5q��h���W������t�H)��a�CI��S�2X�H(;�a���R
w��9� ����) ��
@�{f$��=���������vM'�`bRAaU�
KB�9�Y����<	�ݐ�������Ծ��s����H)���
AH)��z��ۆ:�5�x�
m�?T)��I�혐R
AN���Ad��`��L��H(�lĂ�R
w��/Z�����[׷G�U��)�
�B�
\3���}þn�޵|9�w�8�w��O�
H,�JM����j$��«�$�!H�lĂ�Y42��큈{�����~�v�
6;9��Jh��
gZItBT��i�f�VeR�p˾�H,�RAHz�}���]0) ����
h@�j�d���D;�٤��F��{�~�׿k���C�;���CI����W�������>�`��S'FRA@�wxi �4F�
s��
A`��I-�;�ى��I�);����JH,��{�+^�~_Գ:���޼��9!�.H\��{�n=`{��Y%�{�g�=�F���;���+��;����|����Y���;���K�$���v�d�>�<	�� 
 �<�7��R�nk�s��P�6�RT�}f$L
H)S�� �AH,:���s\�
9�bAa�aI>��!���L�aL�RA@���H) �{���
Aju�����ɇ�J����w�v7�3;*��k���]���
H,����}`b�) ���B�
K���bAH,�I����%$B��
A�=�q�{�{���f�\&�u��!���B�s��������j��߼g@9���@��C�������j�k�ygsw]?$�H)�v�֨��Z�H)`�H�l��@���S�큈hII�XRAH(�l�Mku�{\*�g��$OFR%r � ����u��ֻNkV�2<	��
H)�P��1 ��R��� �AMì)�2RAB��vE��O�)�w�f.�>�������I���%#�]������`�33A͎�H&��iJ�5����$�ܰ�CI��L>aL��H(�{$�H)�����RQ�����w|���ٛ�k�7���*�Y���I����ϵ����O�݁�~II��ZAH(�lĂ�R
w��1�RAa�,m ���bAt����������5�o7{�����AM S��\>��H��(�|-=	�ꋛ�K�:}�����4�Y)����l���G;�4�X�$�{`;���s5| �aI �_�ى �����lCI) ���- ��)��ɨ�H,�Rw��1 |Ϳ��ۓ���.؅T^����K���۔��=�3���ߔ�Ȱ!� �ɾ��U�_��2Q�Й��7qVQ����d�Հ�?�����A��������y�\��A`��I!�*���Y��������$�0{P���P���i ��
w��1 �~���﵇�{T)�I��f$�I>���D�� FǄ�H�z�;����U�=��.�Y� �ᒓ}`bAH,=���_s7�u�RAIb��}f$��S}`b"RA`����
A@�{f$Q�I;���R�
g��s�7Z�s��$��P3[�Dx�.l��w}�}gG��G,��!���Q����L�2�
��A`hi �y�STAH- FǄ�H�|�s�j|�?�_�c�Ep�v���Y��[�z�7���aB�O3�qR��7�1=) ��JO���II�W��RX!H�l�M2�%FRw��1Z���}�g�}����?kH,�|�AHk3o>6�W3z���;{��$���$�0~�S-��
!���$RAN��CI��L�)��) �}a�����W�^kg��AOs��Q ��v�I/��㻻��i�i��@9"���e����!���XQ_\) ��)���f�s\���)��I�n��	I����i!U@{����I*w��4�SH��B�c%$)��i ��w���넳�ȫ��m�xa�U 
#�����) �w��
AH)���樂�Z+�
H)h����M RAf{��Oړ�k��!�%$_\) ��)��f$�$x7v@@��|�gyv�ז�4���B�
A@�z�H) ��\
w���q=$��x�������q���O�?�ػ7%y�d4�/���E��V���[�	�>ݦ֡بo����$�0�
H)����I��RAN���Ad�S�
d�RA@�w�i �4#���� n~���ve���H�&� G��x$}Ϝww��sOO~ �_�1>@��ʌ����!���XU}p���P;�ٌ��I��}n�(�.�.�5b�$�����F2Y��v3\Nu�q�f���s�Om�X�a[8]���5�g�H,�:�AHQT���H.��R����
i�=�RAH(�lĂ��wo}�g�����}�����S���H,�����\��^��s����ʅ$����a�����AOs�$��
�B�
X�H�l�ЁI�2Rs��1$����s��ڣU����) �� k�Y���) ��ש}�4}�g뿾]�5���3} k��DsƬ��R���̷B�]@��[t(t+Ĳ1��9 ��uyy�ݺ��c{�>�szh<D۟QM�2&fImQ��u"�A���r+�ok�9yz��`�ܞ��7DVf�1���CN�^%�&��%�4 �#ž�k/*���]����kz�l�~Q/r�9�-/>�L�H���+�3�m׷_�����Dݍ@��|��o�s���]�oU����*N+a8�Z�T�kvõ���hfB[lBb�^�.�8������Wٙ�WŨ"V�!���7n��}=����0q�<��ɛ�'�q��e*hQ2��Q`J�-���79���AHM%�z��D��E�SF����il*k�G)a��54���#������=�n9�h��7f�N�E��z�l�&5g�-��n}�5�q�gQn�r��_#��q�m�B�K�s�;pf��&ݺ�Z��ܱ������+v�ѫ����k)n��c�]-G�֩^,�@wT&5�q�U�@�B>�5�mP��m��q2���i���Cw���ڈ��3:";Jo��1�9x3�O9�1=�x�,�"N]�F��&�d�=�h��c���C6dqc��Тc�fmA��iD@9�4'{f��m�Knf2m���ֳ�N:ɥ�t漴�Ϣ�G5�3��Cn�M�FTof�ٷ3�$��eͪ�,��m���*���x�d�� ���:++Ɂ��д2}O'�v�8	mȢn�������+b�B�s�Q��ͺ�&�l�H���u�^>,���n��`7(D���k���&NxC�::͔�E�r��nӹ�^�`MS&T�>���[s^ �ۚ�����]�q��F��V"�~�����9�a�s��N4��5��@7wNk��$;#�ˡ����$�
�lRf�L�j�?s�_�&Ϟ~��C��q=`�A�vmd��]�����G����>!�iG|��T�;{�2}�7���[s��`"gg0a�٣��r(�۠�m�b'�jv���dfR	�����u�M����m�x�ȏ��!�nUt���,K".�Qm�>U'�eήz7�^| f�@的֘qs F��5�(۪ϣ�mТu=��5��t�V����m�S������@����jwn�Ӑ�^v���@��w�t��(DjD,[2@�㫴�,23�\k^�e^��{"�#5���B���gafe��i43f}�w%�|��>n���x�Ȃ۟P-���i�j:����r���/�s���#�3}"�7�=�v���f�Ɇ0]B�Ĩ
�ͺ��x��Q�UgV��̎�^'��0��;v^���Y;7�{��X���}x�PYj�!d:N�+1w<�]m�l�V{"f�N]��:"�!3���?x ^sQ���t�:{�2~ ���� �"m�x��4�8�6�ڈ��)E�B�#O�ͺ'�3�V^^�v�C6dp#�&�"�X:�c�X#��+ǣ�nh6�!Ǡ��w����Ж$�dש����φ��H3��5�(|�W�!���Og���_����k�Җ��c�qwhuUt��U���!Z�h;$h��ߺ[��O_v�s�<�4㹍"�t�d� ���j�+z��X#���}^�4���P*��ɜ;O�r� ��^��gt�����&����#� A	�
6�U'���UO�",� ���@�"n@m��mGd�����K�tj˾��F��%�}�8S�f-�CnA�5b��ۉ#�xs2�o��Ĳ#ΒLwh�ʺc=�>��MZ��V�!]��L fwʐ��H)Z��;�=���O��l�����I�GP
�T�j=4���*v�1��2���z���ʔ#�r�'9�2�/��É���y�:o,��w��O���xP �0AOhP!�^�Y%�<��7���li�R+6��+G���%,p��ԼY��VS�]��^.QW�f�����H�۟P�3�U���F�Ǟ�+v���R���� >�� ��
!�T	�3w�ë^iv�<�1��4����v�,��1��1�����O����ۖn)J�hX*jh�#�	mȢr(�c�6�2�nfM�<Q�T+͹|S#�}>�D6�K"nk��Ʊ�Yzb�l�+vh�[s@WhV9�Z��7o3{x@ �t�#(�Jj�n���w��΅x��P �|ۑ`���F�TQ������h����=�ĸr�㗸c'���@��4>-������+?�U-~��ً�^v�ҿ]~"�ܭ{y��d�jRQJ���I��Y��]
�=G��d���(�{ވa�ɓ�ͩ�/���O��.��	uI(*��f�8���HO٧[0%�	�V����V�{1#2$KݻU�6+�wxѓo�kPd��	��h����%^��=Ν����yb�t{`�(�)\��Xadj�	}{�o��c֍yw�Ka/�}���կ��^�˓H�-J�s�����ط��~��Je�&wmk�c��l�\�^f�2Nl�>���Hj4�u��a�i�b�Eŏ�h��r��0;�������Y�����ԍi@�fY�ݼILS7�u��t�j��S� �����e��	��&�ղ��\�V�ܻ�w;�^=����x�1����V���~��I�D[���Y$��ξ#��7=�s��<�A�n��LT\���0�*f��s�&��џ7^X���q�[�����i-p������'���4��$U�|���e*#|�'{�ڡ���7;�廆ߴd�4)[j�y���=5f��ٹ��\�j�L���и���и����Or��ve嚈�ݗ|�G�}��0�o���&�dI�&��u~�{����kPYӾ���z��?HOI�p���!����e��;'ta�(nE��C/�Ϧb�k�yOk��ۣuNO����ɪ{����Ռ����������w%`���0��|f� R��0:��{W��YfDޠ�*tv(��ʣM/w���}���^�:9!����%,�WN�-�Ve�0�G�#�I'Ы28��p�䌪m��۶�G6�ȶ�gq�I݄QftQ͸�㲳;kR]�qu����E�gvYV��#��Ί΋���-;m�]6�]bqq��YgGBad���FwgevVqvu�e��YZq�s��ŖvwBI���6����q͸:��!2��K,Ӓ����Yre���٥�k�7kE�;2"��v[����GIBHt�ͬ��qm���D�[[�\V\RiSjp�(���vu6:��Z��v��(��m��9�v[j-�wm�::̊�a�dI�h�;߯�qߟ����`����q�,w�P��)�b6� 4�v�c`��=�f����,j�	��X���7�͔�8pj�7�4��6�k��N��رn����=�a�
d�� ٩h���W����IvK��x���qa�m��z[���=7��Z���	u�$�"�֍��
�z.)�}��(Vp��a�]�8]r[����n6<��L6u%x��L�lͣ���V�ŭ�#�%��D" 2pg=[<oYb�<R.a[b���h��ˎ�i�;��we2U;��qp���;u���BP�����Y��XY��>;����Q֧����V�;`G����i�D3���)����6�Y�r�}�T
��W���<Ņ��+*P�c���B7*ж!.Ix��i�h4�nK����Q��9&���v�5v�V���5�V�lK��X`��v���DK˟E��q�x��u��'��!�}�VJޜt��]���Ǹ�c��g;͢����[������+CE�;v�(���6�Pn#�����k�n�S�����԰0����*e�+0�N��N�ϨٴZB�W��1��SS�f�����>&n�����E���vwW�B�[��m�JZ�ƸeN,BM1-�P��˵
MZ$DAƦ��r�����Tq̮�\=�7w8]uj�cpv�S�j���F�����`�J;H�t����[`I����l!t�Fq����j�stX�=m�,�؂�w5c�tnNݱAqٹ玞ֈ;z�E;&�H+�]fى�fËq�J�>�qi�+4�q8�c���WΫ�k�=�����X#R;����&z[:α��N��7�p���<�YcI�.��c��y��u�� �ug�Z�i��^�w)t]�e�6v!��pm�yF�����s��8�r��sv%ƱГJk<�@k�������C���-8��L�!�vՂ�LÍN�f�nf㚞�q7j�6���ޟ�|4�(��ܔ�R2���1a97��;E���N�G�k����v�c��;�$O9�����'c%����Wn6�	��Po<M��]�����Ua'f��K��-����h�+j����ϥ.�ΰݜ G���4�e�GV^]!.�34ҀVQ]�bf�J�X1�%%��=����`xn^.yݨ�����9��$V���3߿[�����clZ��p7g���׮ՙ�W�W�yŻV��յ�c7��s��M��`�i7BzQ�d��%���z�a�lA�WH@��� ��>-��*��V>�S`6�]�X�]j��ݼ�y�#��H��C7��Y
�s��Yν@q�[t(��
�{h��޵
VU-����\,8����}����-�� 2ɅgK��ϛr!��l�md:�3g�G"UǕ����N� �p�t�-���܀ȿܬ���-X4�)��hr����wR�y�>��C} 3��m׈���>��<�ݦ����댱�e��A���9�\g��9Lx�p���2�1�+�{՜M�#9�a��s%x��ux���d�����᜞]*0��"u)�%)t׈%�4�G�r(�5Y�㜵g6U�_ �=����xn� u������sv:��&�Ff��v5օ3���t,���W;�
jff��yxG�{������8��t��x]|"�l�G�P�n����Ne 	q)�A}��,��m�|[raA�͑\a�(X�N�W�=�pk�W�-�
 �`�ۡ@��
!�m���F#��Q	�
���ϔh6�'��9=�	��D+��+&�^3�4 �߄[r([t*�5�N����B���\-�r��u�(f�P$q��mרE�ԕo��f�����޾Gh
�J�,�t�*hK�IX�5@�c�4���:���^���x�n}@��;���]�iݵi緄�r]Wg;��ݑ~ �9РC0!�B�m��	��8�Ox���ˑ��v*�Y��۝�ɶ�p�ON>� � ���o)��={4� �ȠmȢ�nF��2��n�m[��"jUs��s_u���`�K�}F^rտk�y��;Ÿ�G�A��"8��.�w_Kp�CQyndk��^<.�E��
�
}B�m���mϊ���*�$婠&Ȃ��6思�H��k��j������u؋�.��#�{]
!�^!�@mТt��hB�I� <գ�s�� <�����A)��͹g͹淮'�z�>���K�_p�/�b��ZF)�v���,���P3\�����&�e�/�{%������B�C0AmС)8��9xӎ�43fE�A��j�e�&H#+(W�յ^ � �� �我w1Ɍ�d�7N@ǲ���Qݶy��ڝKs�ޏW@��B�EWN`�U�DX[ $�P �0A�R'�$�W�DM�H��L��T3�{$<���NGAO���R����G/=�ݘwT#sdW�ǈJ�b��^���8�3C6z��#��q�B�+w��t��Ow ��b����ܠM������n�n���@'��f4�mv�^��n�U�tcL���X.^ �mx��R�RS@�
"<R���>��N�:=���=��in{z �@3z�x�`��ZƼ��e�d��FZ9��R�f�&�m1m��Q��u���q6a�qI��������j��=�摞�&��21DC�h����:�o+Ud{3�}w2�|�p��ݏH))���	>6��yIˑZ�LQ�_@���ܔ��Ɯhɡ�2� �􀒬��ѯ;�ԫ���*�E��x"�)��� �{���u��#��U�{^�Լ[����]H#7�Q�($�D����kj����"ԉ����D�av��byZ�#� ��@�̞����᜶MG[�f������w�-o{�ms�gV)	Ԉ��{%h7�ӎ43fG8�ϤH!%>���
6N8��[fkw<�^��OȌ~�ߏb֯���^Q����#��۾�w'�Ջ�v���zR�B�	�n#WfV����t*ņ�r|���j�E��ц-�]x!Fï����0jY���-]�x]�o�q��W^�w����:�؝ѵ�SWj{N�	87m<�N��8Mh�n�FՋ�opv�	ԓ͜Q�ba���w���+��N���R�ن�8�T�ŷe8ك�Hl�:�H�6�>.n0Dt��l�%�3#	��4�j��Њ��R�e��\�$�% ��ф�~��i_���H,�ɶZ.=b��b�l�{gh��t�z�wJ�J8vm?0N������-S@O:*;�����KŹ�����ʈ�A}�(�>J@IeB `�xS��O��!ձ��#�5��j��p)��ǈ��9���v�̽�8�h�l	bR(�x��g��܉r�v8��7�+DU�P��4�0A["A�'��s#ع��FIۜ��}��b� ��9*;��u��KŹ�� ��@�e�Ϝ)�B�B>NU@�� A	H���ŨbWY1��soO.f�nq<������h��x�)D�A�))��]�K��=ۥٱ#H��i�e���s���b6扖�җhh�Y���i�y�����Т�BP#1F�*�x��94/g�Dl�ȇ3Ӣ��t�-Ȓ;�W�(�AIM�X��\E`�����|�wP���{;-,�2V�Ѹ�o��b y��{�I��ۚ�|0�N��Fo�J������$p-D�A)���EGuw׳�/緄t	ޡ@�v��|��~ީ�����JD�BJ�x�D�XmN�C��
c[��^�\p ������ �A))�(�up3� ����S�4�%D�(�R��i�����P>#���vC��z}.B ��U�Q�zAIM" �MN̵}���%MzwE3�]õ��KŹ�� ��9�@#`��Yso���}>���ݿO3F붶�iV*�o\�80��:q�c.'�HLT��8s,]~G矴�{� �rJ@D!�{�=�0��4�檸�M�]un>���ܵ<A�� � �����"J�Q}O*F��0A�"r�N���ً���#��쀒˴����yÄA��ovh�%|����RП�?̗]�b���t���2D|���i�����=��&�a�6�Ï�i��,��_h��ð�W8��{��ͺz7\n�4�=� o�	��B0J���P;���1�H���$�[ "-���L�i;�Uq� ��k��:!>Q+%�2$�w\׏�@%(AIP�[����D��Қ����ً������dI	*�Q5�f�u�����A��*dD�٤ɰ\zXW&���2;�jv���Ɏm��#��٢O��W�Jj[�wҷM4�=�gPכ���4�����E��	!%"�!gN�;�]p!P��ȏ:�зv&��'u�W|�M�(��sn婪3���4i�z�gj�v�7��6�;ݝ}��m�U���;]�n[J���={3�B�{�	`����W�(�)G���Ccr�q�S��ȃ� ��K���F��X�߷�s`H>���l��+�p"��U$Fo�^{��p���u�cnu����ٵ�C.*2�u�twU�ҧh�~�>�`ۡ�aV`���H!% #d%"A	)3+^�s�}�v��X���[�q��
ޚ>�#�(�����������ܡ�2 �L
3��z��oR��p�����pc��.���2�ǲPk�In*B>��HU���:�s��c*hnOPQ�Lᬵ�Y~ �UH�F�R����3�f2���~�'ّ�>z悽�����i�m��i����D]z�5��Y"Hŕ@��
RK+���*��^r�z���u��IW%N�f��㯦�}��G��%4�@f�\t�5F���$Ŵ���J�]Z�֋�M�e���P �>�ݕ�(-U���U�B�����AJ$JJh�QJ3�z�f�\��.�hy�v���.�[>�+`H5�(�R�wv�Ń6��5R���e�ޯ���ܐ���C�c ��O�'�Ǘ���DQ'ڼ���=|�Ljzi��Rd��p�r��B�ho�zoq�-��Ќf���х��z	'q�ڇ9G�2$��FИ�&(k�mAD��K��n�+�`���R$tk����rD%BLv�5P;q���٦:p�=#��D��,tŖW�E3We�]у��QGa]��=�-��!Q�G��iEђEv�f�20m,�C6�\��s6���,�B`���	�VZ7	5ƌ)�u�ғ|�/�߶t�n��T�x]���x��j�	�X���
�*�p����m�+����u���	$��DC�o�{�01*����qE׌r[�s~ ��#�\zJJh�)@�A�CN.��� �"|���(u�g�{*����F� ��Y����Ǻ�������x";J�{ݘ��u�m��z/l�kc��/`�F��%"@!%^�|(Ż�܉<u��M�=ܘ�rT�vn8��ϧʒ3<�d�2D�Q �c�>P No�[V,FJU0yMÓw7$�W���ɽ�sCrz�i�>{"HIP��ݞ�����_}M���A3� $�vlBڞ74.z��zy��[(�L(,kvO���ud�� � ������;��I��o@�%SF��A�<�@�0AJD�T(B0��m��7X ��q�%�\t��,�{DNL�c81=EB�5��I���<��g���{���Z��fn9r��)]�DR�8��6��j�^>:Dy�oa��_%N�f�><�k��� ��ӶR��\oR�s���U�X����	����ۈ���w.C���MSɗ��F���F�=� ��P�)D����;:��Fv�D"�tH ���W�b�cx�Z)5�����	"'j�Up�#�g;�@�0Bp$��P$# ����	&�e+�W�őOR��WT�$���x�y���� �>))��R�.�s�w��z��߲�"KQ�h�ܮ��xLޗ�����`�@�3PKt�5�V|��$g��hQ� ��JŏSB�GZgud�ܞ���å��q�WH��j�@(�)D�|RS^f�5���,��H �[�{�+�7��u�S[ހA{H��(�K#p��a1 dȟ.�@g��$$�����%J����N�q����^���M��N�'�������{M��m���ٺMf�NF����G�V�:����u곉8xWѱ��򴜞���y�z� �ϴ^>�7���<�|w�/,��Y�h'BG܏��zw��a��>!��1��L~��iq�7E�:q;�2�&^J�9�7�M�ĺB^)梨��F��t�����;�(��/Y[�:��Q	��E%y�{Ig� mý���x[����yK2���6�{���9�zzn�{����}�%m���=r�;���;�{NiV��F�aLh�jFj)`Y��mj���.Q���j�79��$c{��=�l�v�s��Oi~W_ ���[�^�j19b3H���=՛�6!�j���N��ٞ���t�5b�k��E�3�H�Ԝ��Oz.�����\��-6�Bd�^��h�9��:����������;^3b����x�
z���Z{�h�;���&i�{64iŞ�S���|��׊�� �{(��KZ����vN�5T��K��<�fN�w����6�+Ya7�w2���,���/hCP87��H�|;D�s��{�ݡ3���y��{�A�S����{7=�z�;0�]P�u������lΘ&�6�Rdvn�
Gk����}�=A{q#�I���Z�g
�n�-�u�ᱵ;cyj9��N����������/OP��]-�o����o�}�|�:n��һ��.��O���  �l:�MY��e���dY�m�sj�EYm�\BG�A'!����L��l��N����2�3,�;�
:�[jʶ�ag;5eaնwFY�Ee�F֔��E�5�m���:�����ifvwgE��nnj�F�6����b�����[]��DvvQșm�J³m�Q�n�嶝:u�)�nQ�k36�6��ٔ�Xpu�lͳ�m��6�hӫ-�QD%��md��qs�C�$0��+;9(��f��`)�@5�b*�r�ӊq,�f��Ⳮ;�k

i6��e�*�SM,EX�

^V�p޿\,ԝV���O=�Q�䢈 ���|�>.�Rof� �5B�fJ��;9�S��3��dnO
L���"\uѺ�����D%;�X��{�v��u���]�O���i�{-u������)��o��uu
#���pi�b�_��剂f���y�ާqn�.���+��&dsw����w�]����eo�Zo{�!�8[�d��I�k��a�e�<��QъY�H��H>IM(�JP'�1!N\�]��`@jD��RZ�Ǝ���ɑ�=@i�>{"A	!�BtJ�(	6DN$K�4A(�(�	IK4���i��emTN��Ƿ�w�Ij��%"HIUy�e���%�9��\�f<A["|C�U��i�Y�«2��uZ��>+�h������>Z�י�s}�>T|�z� ��X��,�����yi=A�o�d=�zΘ��mp�����@m:�;
�{�G���7R��踎��16۞���y�Cw�'ݙ���I�Ց"�dq`C�BJ}Eu�Ȭ���� �Ż/6�&�cv.:K\Z�,,���1�� vz�a��uE�]�]���E���"=f�X3iM'{c�n�]U�5��#��3�B����*�
3�Q	*�HF���*�/�[t(D�ķt*�9����W>+�hq�P����٣�D�$RT(�`���r4�ne��ڷ���oVD����0#�dI	*�Q
Q$\��n�
e�{���}`�(�))[SǬkⶪ'Bkc��;�$�˝�f�΁g�!%"�ǈ!)	-�����5�^�Z� �pk0�\�rn�U�p ��4A����
Jbؗs����Fљt��C�N00w���2����8=��=� ���JJI���l���e˹����/�������GA�w�Հԉ��(����-�A�]�g�Gn4�\����<�3���-�olL��7A�� �u�� ��>`�lhS�.�Ŭ�^�lvK=�:[k�L�ʻB��Hp�� ݴnKpv�����Y�T��)2$��.Ԯ��hkvy�M�q�%�p�N��9��sG����^����JGd�}��}�򕍝�u����!��������<�u���0K,&�u�Y��5�%��v ���K�.%��}�gp'�[T(�`�ŷ��^��E<�4+g�U�D]���yHG�H��5��(w��G{��ٕNUW\Dծ�R�`���ŵ)�������5����FoP�Ѿ�/��P��$vu
�<A�R$��
����V�coC�օ#&�9��Wq��V�׈ �R�H))��B�2��F�l>�@���^#�����q-B�ObP�pح��I֑)��sZ�y��7�fF=J��V�
Jh�Q�P��:��ˍ�m��Գ���	��it	 ��
�� ��[wӹoTտ(�L\T��b���G�L}�#���8a�ڷOK&�+��0�X1��4a�֌��Gx�0�D���W����8f�9��Wq�i���x.ؿSp�l�H�q$�׼|���O���u�����\��������|L�g�5�����U����/��
ٚ1膰\fL�L�<r��nx�+8^;tC�����o�5xaޣ8�0{sŭ�=�C��b�xP � !�	!$ѐΕ+���dG��I�5ϫ�%��Å�qͼ�0��"����aGA��l{x@'z�FwP�Fy)%��5�w����;YK�$n�� ��L%�t)�7���껎 ��f�E�Jo��`���s�,u��7E��b;���&�kg.b��y��/h�b���l����&���v���׹_��zn��S9���4(n-ѭdG]�l�<One���붶����_g������Yo�	}��	IM�Cz���+���l{z���̔�DT�^��C�^!�%A	*�A�+s��537���[^�Q90�=Ч�g7s��8A]�G�D��rz�s�,� e�>8�		*��JA�z�3�0J3	g�t�d�n��(U�V��ݪ��2�׬k�>۞4US��8:��숁ՏK=�e�2�U���)��Pf6�h^���N�
���0A��$���
"<R�D�Oj����R�j�O@,�:(AIM.������VǷ��}�i�{))[r4ϡl� ��
�(II�9�,ۨ�����8k3�w[U��s�(�J�t�$s�����i7��
n�d��Y�q4�:nK���,6��{8� �5�����Pfh�Q�u@�BIP�N�u�W�	�蝎�_o7u�w���%	)�9ʨI�]uHb/�º;�v{�==q:έ������	k=Vnf�҅HД ���[������tv���99u�<3����Vz6��Ko1��/��%7�[VIW��m�b��މq�`!ϰ�V�H���k��G�/f(���cZ��� ���3�{p���B�1���보uGf���2g^�"��ʳ\/:qBQ����%1�׼{'aWFL�䅭�N�9�aƭ���;�% %V2�R'�FX��s:�vcE��m;<nT5�����!�p�����ݚ"j"�U&EFV�8�J@J=Ʌ���p��'.����찌�c�����f�~	)�Q�0w0r���ڽ���{1V�l����S��.;�`�	&m맑�{B�ϒ��y$GP��o�7Bۼ'��C�[�z ��J<�y%!�[�u35�*={u�	F� �Q�w���ڞ9��3��r'���JP�JB]|��������ٺ�noE8�=�7`���� �T�޳tw�2��1�4ڜ�YY�V	��now�Eb��� N�;�~x�o�j8)?�ד����<�"Ue�P��P�V.;s�8h�z��A�����M�<V�mÀk�ə�q`]�ɗ��`�T���mVb�	z]�1s�2n�u�IC�&�'���cJR�z�I��$f4�af۬gT\��ABgQ��}��W$�Bv̕�mb�f�6FR�4&e���
\{<���� �5z�����S�f7��煃vv�Ԧ]���CZGk����Ϥ�	��[r4X�:y�t ��<&��lW��)��ܤvY��{�gٰ�$�bg����&���V��%�u�U�PI_��P���7w�@��s������5|��[Sz�{z�yu����2I�'��9���S�'�pt�W�;�u��m�����S��nǒR�x%��LS]�1���rJ��K�7��<���z7�2���]�Ԓ�%	G�BY�SYT�j��7͌x7��5|�s[U�;g���$�OT־>�z�����������k6��\�+���ۢ�0�dM�,2�a�޴3u�%���ݾ�|��ߝ��]���5<�V�q���=�iY��y�@�r<�� ��Q�RaN�i9�,�Ccn3Dn�%��j�&��۽��9Ä�h�a���d��j �/w�$/P����5��̣���.�7o/�o�49ձ���!'�eR���\)��ݏ%	)�J���q�+,;���0��M�mU��o@JRP��i}2�c����[#� �fJxwP�3��ѧ�uf[=�0MV�N���JJG����/��H�.r�'/B�V�oxxCձ��7�grV<�Ն�/��i矼}��K�s���,�Gh$�v�����Ә�����7kd4a�֞ϟ{��O�I=�#�Cl����Qؓs{T`��+6w���x$���*H����K���G��fO<���d�rq������	#�s�������Ҕ ����s0�����ud-�5^�v�D�,�8y'���|}��;����B _I�&���=6{�鞖��nb�s�=���K�xa�7�D<�;�o@��	G�PR-a-m���T{�	kf���c+�$���w�zw�����<����(�PR�E6����05�[��ۂ"�=�U�����JBW�es�1�O��	����]T���̕������h{`��\g�ײ���ld����%%�>˾3�M��7N�Ȁ�$=8�-�]zZ�=��%)D=�bwMtM��N�ٱ��4_\����\oH�e<��ӈa��kڷ.�簒J�	n��F:*����0k�\�ɪ��ǆ�y%)%^�z��ا����tJq�Y�;��������of�84�W=�Rv�u��qk/oj�d%���v�}�[�	KUuPI1tȷT�t��ݳẠ���B��	��d��b[�js ���k�����%��͚&6 ��zw�4g\�M�ڮ�#��[]k_�s��ԗ�D� �
�z6^��2l�����X��f�vM��hyR�\��~�Tv���G�%����b"���S�܀�I��"�W@�rP� ��]��7:}��4�W^!��:'x����;�ތސ�:��*8��䁛��	BJ|�+��U�f��RM�ڮ�oN�%I%bZ��ˢ����r�-��#]��ݱ=��70�7��QL�X��v����$Gt�chu\���X�w���{�{��<�%a-I�0/��Ȋ�܆�P�1�,������l;�ޡYMT���fkKRLrr����I�~��o{s���	�䚩{u��ș��Ѣ/g]E�e��Ӈ]�t=�Z�%n�]I2z��{�Ml�P ���yW�k�N$x/Fb�Y��ڽ��`�g;�c�\<���7�I.4���Ħ���a`ɯ~�\�i���z
]��>��x�k�}�-M-'���	��'����)h�KofIQ��s^Z�	4D;W�_��Dg�o�a�s�B��C�vdG��Q�.uC���P$B�*ᗃ3#l_{�+��ۉ+q&���ַ�D{���&=d�ͽ�ߌ��O?p/G�[o1�<��X�YpG{ve�J���n�W{�;�$��fE�}}^x�Z�h�C��ۜ�sw�#0�����q	�]�I{o�.�n����j^�g�u7u�'��=�匍�ON~Z�7�Ƀ�����fY������8�ѝ��q7s����nϽM^�5�\y(����*wD��4t����DcwQ
Z��o]�:�q��;�V�[N�<X{�i.��;��Nl��T�[�$L:�V�`ԍu�y�v�I��%/G:�.��zV�b>�9�m����JP���{'X!nQKѳyIOWr��aK�T�w��y���H�8o'��ȕ"�e-��Z�[��w�b%��*�_��������޹wG�|c�=�+���5;(A�զ�Z�2
�cu�D/s�^ɖ�=��j�����P>�Iw�۳>���)���4	[5��Ƿ`/�YJ{�)��Ozw,}����:�j�z�Z�3w��*E
x�؆q�rrIA�;mNF�gqA��l���fqE��A�K8��̉I١�Cj1,���t�K!�%�"t�β�"�;���3H�̩�3�ݙ�R$Q8�$�m�̄�v�w֛m�2��:%"�j[Z��H�8�$㤙�$f-�t�d	�tq@BEe��E��%$���+m��L�rBv���9ܴ�.˲��,Ӥ@��BBt��:9:Ve9(��r��m;l�"̶�\��$���3�� ��88����Hδ�(
���&�ZE��j��$��m�f�쳛wn2njٹ�Yh߮�9���2�j�if���K���g��d��V���9s���c����n��ָfW�G�̤!��kIa��[���9��u��lrA�"���A���ӷÀ�����G:R�b�e�K�aK��a��cX4��Df�F�ˡ�ej&��0d����z�i�����:�x����([	La�M�Q�yH�[�n69v{��sV�+�e�l��`hf�D���iHb�,�&��IG]R,���M	2YNІ����q�؊��^*G��痋�n۶��3�e��3Yu%T �h�ե�>����=�K%�c��>�.ݎ#�{7C�&��= {s�ݗ+���+\�]�kE�V�st���؋���2t�'7^���p�z{gn\A��r�/<�j�p�b�s�-͚��Z�9�J��x���CgVi@R&1x,2ˋ"Պ�̵�RҤP�v��u�@�fa��8����Rj���<�r=��q�B�͕��q�x��p펗��f�
��{��V�8��&�nNx�i\T�׶`{Q�G]�j3�tj7lF��ޫ��;I��p�\M�&lɄ>�i��1���B{���;���NR�9 �����ͭ�^�Ĺ��ܑ=�z�� uW��m��t��y�q�Y�%��l�J8��dn�&̼cn2��-��.�ej�����tgJGT�A�M�q̹��ɱcjz�1H�pۏjU�l���i:Q:�s�=����Wsn-��J}ٞ[�g���i�.�bvrk���۟`����z�Լ'"�\68��ۍny��\�(�Ff��p��m88-�`��=�y�n<F��C`�q�MA��ɵ�)�lJ i�n�e�j
c��d��h�M��.e�:٩bI�a.9�N�'������ΰ4�h�m#�T��wB9�:��l�O��3c��4�F�Ew+�kg7Dָ]�P�u�|�b������8�W�������.5s"����{����c��`[��6^�}n��wXk�xsj�>�Z�z�$�̍���8<��Q���ikv9���vˠO#���n����ֱ�=���^<ɫc��ѣs]v�q	ueKz�n��m��#����ml�յɬ� 4�����ݶMp��n�j�꒷K�i���ب�%�#�Z�%�'m3ЮH���Xu),r5��]6�����Ҹ��r��a��v�j9+��uFr��@���e�Q�%
�K����O���$���Z��1ٓ�6�j��#GO�-
���x�m?Zu9�Oh�g������#�n؊��ٛ�iw��	,#7�75�OT�=۲��%4v{��t���"�w�e�=���w��>��$��F��y`�C�ۻiG��|��h��ěu�]���,���\�p9(	@	)Jk�H�;@��.�^w9�u���ݩ���{v<����rT��C1J�V>7�$�ٮ������<�
�,!����&Cf`DM2EULML�0�O�(J IHHv�Ι�=�{��25FJ�׀k�VPS��x����Hop���[�4-�5�'U��W�ȏ?n�w�9S�b�P����f���*�;i��ϏE`ʖ]𪌫�&����pp$s�W�
����	ǵ�Z���̔�u�]�ӽ	=U��T>�>�	G�JR��+��ҲD\h��"�����WV�������IJPP��BN�CY#.1@IH	i��;�`�'7wc�b��̎�X]k9G��JR���%x��L��Y��:¦�U�W)6�j�7���Q��Ud.�3,�����)k,�p�m�ɝ�3�%�r�ۏ:v���Ԥ` ��	GE�=�Zm.o�~ٝ�=��U����4�����	@J IHMF旗Ilxb�K��.1�{9��8>�%��*-u�g�(��������%>	]�}R�u�*҇+$x��a���P��cgXɶ��-1S���y�=�l�=������$;��.#5�/f׮v����s��W�\�ۭ�����	@IO�� ��c��=��d�[�wG�Qy-�N�.{ov�&x'�6�#u�8TJ�7����(IHJS�/�qR�ջ��c1�w59���'�_��t}�k<�-GVFU��ؙ,zu�U���f�讃X�B
�	�0h�2a)��=ڒ��.W�k�B˔�u�]�sciܞ�Fm�t{x$�((L�ʍ�˝V��O:�=�s�{;Y�8�I>�8�ڽ;�1��)	@J�K^j3ѓ%*�1�y jswv8q���J����jgLi��s�m��it��_"��6�m�{;�6T���l�:�Qq71-,�HYyIF�/
�����|}Ӈ���Sq��2�MJ���i���2�CH^��66W	��[����$��6����X�ܬ�F;ogiD>�q��	)�uO��۳7<W�i��{b�f� �b�ݞ ��y����g����S&d�UD<�.�@NPRf���=����ݎ�/�,m"�f7�d����%�vun��mZ�P.�=��VT�ӭ��3�@ބ�s���:�����?��l`���zҥ7���{�|��R<�T듇���'F�B3�w턒Cg�8�q�T�����<߭��6���VPP�/����z�����o���,�O���gv���$vgA��)���J������a�A�=B4�-�[��97��҈��w���'�l��)��{�yyرl��J?Be�ݾ�>ke���B{�	��=��<+������?�q�Qhݸ�Z���� �)��%`�ச�K4�	��r�dŒ�e竜اO'a���9�#���'k]��!���԰���ix���`�-��eh6�lp�K��^q��j�Q�bz��&�D��P�e�͋� [.�h��,�)Tz��XXb�h�Ά��j̑�j��*�4l��,�Gj���Hd���b�m�%��l4�2��}?���P���k�Yt^f��+]��cO�����7O�"`MUTje���sJ����T�Ȯ��6r!���p���{�w�W��%!�M˽��Ǟl�����ǰ1�wc�'�QW]'�uY�F�nX� %	)��{kMGq��M����P��<N��wH�$�MGoQq��}w gG��y��uK�ңsc" �:�i9�Ȩ����,���% $��%J���M�v�e��K�w�LV=ӽ�{!(I����|V����Q"���#Xra�B�W��燙h<][�V�v�d2�r���<�I$�����e*��i����ib��F�o@�	)�PYg�U��4V@�3�����E�E�V(Zڮ*:L��{�n��D�V��K���Td�>�g�w7NF&����z&�X�a�Y�8k��/9�O){"��nldC��݀G�J��P�5>J<�x$���t4^ʭ=�H�z���<��P�J�ʋ٨\������%sY���ҩ��N�����9!��[
��T��y(%>	C�ڒ(e�5���������+V�D> f@�IXJ)�;�ըQw�1�h��GhZV�3�
��Jf�@���;%�	@ukfي�����}��JJR=S�q�<��u���Q}�{/e��(�����%	)�Q��){�"�{.�O�@C����2�Eeju�|wOt%���2j�K��Q䔥K��ʜ�ޙ頲"��Q�`Lݳw��8���5��L C��Ųxv��Q���ӵ�|H��(<33QR�X���z��r��:g�*r]˝N܌�5��r!�#���) % % ^���sb�����]�I��{��oV9��띩�2#���n���BP\��٬�u�.�5��c�\����j�;��P��9߹{�n���Lֳp��H��~Ҥ-�8�;ruv�v���7�sr`��iM-�
a�z���=|R�%��7<��Yt��!�CXb�w�i'cr�bJ���n��
�����������.a�Z�xn�I�Y<���YkeUP\�\ �y%>J���i�;c���eju�}����	G�S�%Jj�����r}{��(���V�o)�۵�����+�".zQ��8����l��U�j�h˧q9���l�OrK�\[C63�kȬU��#�Y����� ��p\hP�37�Ƚ��{i�܋Q/�e�jU䔄�)�qMv�:ue{�G����;���w�#��r�%�(Z��4�0�:@�"D�"}˻�|Ic�LNu���Ζj\��M�"h_������%~Jmo˴v+�YZ�m_z���	�=}�C�)J�qe��Ξ�Y���湾��7��۵����t��Wwrn{7ϢT.��P�$�kW���V�t�E����Y�����P=ܤ%(%>�!��ɚ
�i?M�͟$�k�>�2o+[���ގ�1'z*�\���V�y$���o����5{����}7����;v��!��@�$��˭�tT�ӰD9���u���Y�?f���͝�
���1��֪��[fA_����]��Ơc��u��YX&ݒ����=|�5�μ�Z�a<�@�N��u�sE��X���:���6��\\=����M\�fF���]�@��l�vN{f-�l\���a�kOh�^^�S��l������\urtr��v�����t���4a-R�n�te
/gs4���vX9��n�ύٞ15��5cֻA�nlK�Z#����%���Y��wLO��}o�u�u��W<�մؘ��P������h� �mQ^�R"ETA����BPKc��:6V���u�������B��v�I%a(�M�SS *��p�ky�݊���nv��}�7��Z���m.��vv��6@<�����L�����]z�gT)۵�������J@J���3��8����q䔁�3GWttt����j�����>�n��n�%���I_��%	-2����^�m�{���΢n��;W޾�z J I,2d%���}vt�a\m���SbgiG�F���^�X�& :U	�3Pj*LΞ�T{�HJ�������
]������t��Q˧% $�k�l���$�Θ�x���ҜF\\�$��t�j�8nE�N�%h؜����2~�*����-����Z�\��ͽy�JP[P9wGGN�Z��o{ܠw9	F.�78�M��<��y(	)!*������$��Ý�Q3x����_t���)Jkj�uEi����#���szڽ�Q	���ľ��gz���pq1��|�U��%(��]�FۍR��'��ӰַU���敥�c��Y�;�&��W�j��32�n��kpY��'nCg�im��Ү��͸�c���_�%~Jӏy�םD��n6s�¹���Ѧf�ݰ�R�y(�Ν~�a���Kc�c׮����ۉ|���IB#fg\�e\͝�����$�+U�ߜGߣt�¸7�oRr�AcFK��ۧ�jC��� ѤC���:0xvqz'A
����q��t�٥�t�2�]��.���3�a�(��<��zw�<d����{_r;���h#����)w�����ȇ&�i\��y�3����&=���6Q�PpS�<F�nG��9-�]S��"r{�,]�xyu��ۃ��v>E���vus��q��z"a�@�Կ�M�]�6gl�E�޳��Bo8l������vzge�^��á{��<�O��7#���>�2�L�+\�5/?[yrYb�y�����)����u��(�i�s��w=�r3���M�ٺۛ���,fn�l9SXq �͑/x���7^9��¾�K�¯P�r�ŪL'}/�_z�u��,�t�ԟ����	�dnu��`�^����[r;4{����wqU���R�r���]��w��2g��/;� �224Ȱ)o&���9
���F�w�V�u��oe��ӹ�/z���_����ח���6{`��Ǔ<�k}g���ugq�H�n'#�:M�M�r�����P�tC�h�@O�t�%�}�c�ݽ�'�Ԗ�*hKC� [�d���hmh�G6u�%��NR�7�Fv�4����	lipY�c".Vڟ9�Ę����6�ߥ)׸ÇQɉN3L�������=�񼢇
����ry�)�fu=`�d�����rc�{����Z���ފq%�f�����ź���͓��(K'��矷f��ۄfI 8D�9f�q���J��qrF�nQ����s�n�rA��nu�N�Fi�6�Ѷ�#km�Es����!'G�՝�I9[g#26�A.N�L܉N9"Q��R�EmXi��`�	m6�;l�F�8$(�dC�NpY���s��E9��;�r%m�%-��씜N)·s�����H��ku�BYk-8�:#n7I�ִ�ӷL��s�[�؉
t[ZI��e�&ܜQu��� �f�jl�p��eȄqH�\��r�����	@�@"�)ĉ�n:\�[IBR9��3���H�tN�r:6�h��$t�#8ݵ��N! q$�q2Ҁ[m�Pvݶk�g@B9�Yړ�Q��"vnڲ��[`�#���P5%��mT�w�#���	)���}{K`%t^t�%
�s�����l���Mi2��j��Wl{��%(�JBU�%TC�R%G��'15w��1���ľ𵮒R]���^��-����٤6�k�P�gnW���/����ު+�8I�4j8�Z��~��s�S���ۿ`S�9wGGI���N�윷t����y(IHJ:a�M\�N�Kג�y[����|.Ncl����p���ݚ����$���f�����Xp��9ǚ���Ịݸ�޵\��(	@X��NO]nuǱG�Jp)�ωޘ���N�سz��U}�6�6���#�J�a�w���rü«�E �Cj�i��\/yl��7�vv��m�tE�=�<��`�(O2�V����IH�P�$��\��0P��U�>\����I���_t����̕���xg�F��<vqɫ�3$���NPݼ�֎�ӈ�`����D��Vǯ�J/[��j�.]8�ڊ}�T�3&���&�=s�%%':��]��F���{��8���c�wu5S���;���2����� ��n�[8���#v�]E��+�����֩���}��*�JR�it26�y1�=fG���Vۛ�J�.][���j�}���s7��t%%!(I5�UNu�.r�J��h���MT�p�f�<���uut۴��d���P�s��e����V���ԥٰ�L!��f����x5E�EA���V\��O�VO\������؆����n�(���Z��C9�#+�f����pius�]m��l@�p�����ڷ����A�r[�����.��ݡH�z�8y(��F��3v���gZ9��Ϯ���;<��z�]<�Kc3S)��5A�����Ue��4ebjd�nJ�++�#b�J�>ɟ<%Gt��;4
B;�9)��toi,�V���S��}+�*��V��y|���8����ΰv�1M�!�a�ص�sCC�}{�����%`%
�?��u��KTۍ��f���Ǵ����۶��������6����p�z�u����%ѭ�1O�Y�	+C�Y'S�p)G�9�P���w˓�Ę��3��OF��j�7���s��%"nf����nI��<۟%-����T��m�����ܡ�9s�ۛ % % $�(�`�¹������������3O���pS�M��f�����}����m��\��b��\���LdL����rTW.�&EU�T��뮐��$�b�j}=O[U�#%!��.�N\wV�9Д��(	��~�L�R�ה~n]�N`��g.���4n��%����sF�ך����B)���ݵ���	3N*�ꀔѮQ73+��{-����s������;��;GmF�P�����=�<R�]��� e[��
{o��S<���3O�G�pR J<�qɭ�K,��a�J�!�#7zvOm=o*3x�ra�eY��� 7	)	G����GEm��+#�j3sOk�2��':�}Ӻ��V�U95�rM�����5�v;{H��M��=�j�:vçs��n��h1"$&@��	CM�r�uTOi;{�i�t�˃�P��!n�IRJEV��Jƾ��L����d[�Es�t����󐕷��Q�����)d��$���/:�jb�B�v͚K��^D���d�k��S3���5 �x�n�crZ�zi�Ӳ�m#+��h��c!ĭ=�u�S�oR}�)nƽªq�s�p����J�JR����Q�Ri`�PP{��U�Q=�b�MS��j���2#f�<�.�}�(�J@J<��є"`�ټF�f�N�\�];9�d��$�)�����:cFv�ɣ3Қ�jܙ��ٍP-�5����Z�:��;�I5 ̊�)怚J��}�����J��)Υ��/����]�f@�%)@	X&���Mm�;���M�WUD��d�Y 7	,sp\@u�$��%4��!�9D��&�6By��{�����>s�(Il��Xث�}#Ր�g�B�����*����Z�/�b����V:���0��bm���^�R�6�ؚZ���oZ��E͸�U��{������'���-���#�:�T���
�:�+,�.s�%%>	\m���*�P	r%�(�c[{uR�r'tܻ��$����M�풌�"CGҘ�c;m�W[N�Oi���LK꺠�v����i1Q=ݒ3�(�JR�wl�%ېݜ޾̈o�X8���f)��,RP^l�{U�y�W%��[�����+�ۄ�Z�/zG�R��ȞN)mI�!8���IH	G�;)aȎ��b'R�7�7/�"wM�� p����H�r���X1Ǟ�IH	l\���j}��9��9C5��M;�.�BJ@J JI����7��5�w3�q��+٫)޵޽���P��=%�ˁ1�U���Tq��YU�W���?(�--+E�w=W�g�xt� B������w����p�s�zFݘL��\ANҳ�|p���5�Nـ����,󻜼0��j������5�@6�3�V��\��λ5.��;�&1�ݶU58zn���&�0��Y�˘c��k�9�{nx@���%ۚ`��f�n�=h�O2��K�z)��BE�I��q�bjj�*�c���@%�����
�����s��a�I�c���G$�a��-�k��Len�]:6��ݐt���_>_ߩq�k���v���u��K���[H��8&��̈́�dɏP�L�M���_)J J����]�>܉�6��T�]���a�o�z���y(%#c�o!�[��q�[R]s!�회o�ã��v@|ҫ��l�Ħ��=�s�	@IO���YZ�0
C�5y}�ɮ�9VSZ�z���v����A=��o�{��� �|�5Gm+��ױ;��w�dyB�utw���wO��PIZ]]�NOt�<aH�Td�}�P��p����#��J��v�����ed@��&
m]�>�w�v8���Žr�f���ڭ��[�^q���*q�����I$���1�݅ue5����R�~K��S�m��֜�����U��ە\{
6�n�%���k�@�Q�Y��kYk����F]�,`��l�B��o��ţ��ou!���d�s{������#K*�n5��}���i\[��;��vd{\$�4F�\�3�&6d�Q��V�y$糮�L���5��i�{����=iZPS��j��&o����d%[}��;˶��5����H��./�V�d��O �!($��$�qX������>��P�:����ӊ��̏{�$����a+*�s�DDlUTW�#�f:�)��M�rf˭�x������k�n��z�p� ���--�m�(voF���3C`ː���$�E9&�"Lb��b������[�
�q�O���v���*dlһv<�J��x�c_�fҦ�	�w{x����֏/;���JZ9����zo�&7o"��LZm��`�'`E���ߐ���,~��������(�'H��.�7D�[y�&uE�z6�T�2<9��(	@bl�#c�(N�հBJ|��'�v�b�b��܃�Db[���������(I3|��89>�W��2��lB��ǩ����r�����sR���V���N��r��hh��t\m"Cd-�ƺX��\[�K�>���@J=�oo7�D�ܼ|6�T�	܉쾊8�)v�a$��)9�qv�FpC5j z�.td�����QL^���R�*���}v�I�T��	@IH.�pN�rT�����9�q�vϷR�R�z�:�*�v@�	@�{y�2'+e��r�;�zyC�ϘaQ����o����s2qi������˄-mN��7C4�7������#�`�|�y���!�A�O���WP�?a�_8S�n��n�]���%IJQ�\��:��w
Yެk�6�m;��S���\�~�����|'�ǵf��ڵ-�Fܔ��al�����<��wZ��E�Z�'�^��~�I$��[��������{�M⪻�}���xS����J@J<���;9�ɟ]n��X�]�t��5��&��8e�Ԕ���}R�*a�j����$�$�iR]���u،��;�o�E1{޽��	@��������Q�!،[q����Og�J'��w�y[���˼����@���R"r�U��_��N�x��@F  ��
!)�ʞ"��∋����f�x�I�W*x�VD��Y<RS�)E����)���J������;$\J��VαP�yTٓe�laМ��{��4��h����R�S�f��P06Nup�����f�w'N����k
��g=��s�8��>�i����5WL������t���;��ؘ�/ �����4���0
���P�Ig�7�n��o]N�έ:��H��j�Ϟ��c�~\�s��lWۺ��%,s~~���?v(\vz�ٸ҆������sX��t�W��u��6,������ݧKy��	L�[���� ��~����M�c
P���A;�r����!QG�:�_m鐜y���%�Yo��^s�y�&�k�}a�]>@�����e��e��n���7���g���3ܑj���#�HS
SwVgY{p�ɩ���,D��]��q��t�;�7a跗tڏE7�ǧ<���7G��k[�t����2}��0$]'����Ӟ<������z�G���"���F�Ⱦ�I����p	��S�]m�����)t�(�?�S����3w�~�z&Lѻ[�8ҶԲVZ�/D�ѩ��Ճ��^�q��t����2��9�_�J=����z�<2�^����ӷ5Q�ӓF�r{
}��˗�0d��L�Śǹ�S9��7Y��C݊�\D�<iă����2�}��!���'�C���Xa��G<D���E��g�:�F�db��G{���ߧ+��n���P�����7���R���#<�?R��sz��k'�}=�zP��·<�n��z��m�����߻w]H�r��IPX��[j�n:7TJRq;n�E:[h�Z8:
"�3$p���mݹ�r����NDee6� �Β��0���H��(�;��e�9:qf�\���H�8mۄ�	�!$�㥵�p@��	
M�L����Y)�3�p�r@���8�)E,qfCM��Xs7Ya�����r��㐢�#�G
� �'rJ'� NQm�P��tp�\۰8R:I6���QN�㔬��9�ɵi�C�GաY�2�Y6C���mi��E8��9�����.#�� � ���!�r�"#����NBu�N��t�Fۑ)"Ȓ��	oK������s`�XT-a���j3q�flH�����]��D3U�=X���q�S/��D,+	yJ\�i`2�*��k9-í��M�1�)��)�������rB��<��lC�C �X���^������n����H�F7M�ۀ�<���31e$ۡx��������{�8]�Z��EI\-;q�<��k9˫%hڎ�r*���	j��m�b��\9RXv�cE�͂���E�aK����K�v�
f��l�#�����^���vb���ѣН`x�jɓ�u��tZ�nc�l[kOg����6�x�+�;�x��xK&�� xx�a�	���y��|���0�����`z�1���'lk�F��`����6��alk-s�i؅Vn{[�.��<�H(b�s�+��$ާH�u-N��u�	n�S�Z-F�iy���M��ܤrJM��Ϋ`��
�y�i� TŮ!��4Ķm���M�Ӻ�P����NT-����y{t��Vc�В���=j����VN��5���i�Z���4�*z�:ݐ�ʜqcr���v�Q�����q�|bQ�l.�;J=�ta�����)��e����d8��R�Snڒ�Pa�bY.��v��q��\i.ݍ�sE�a %J�:6���h�1 �6���6ܤ=�KT�k`��,�Y�.&$��V7@Z��ͪ5���]9�}�Z։�e�\ݎ)6<���R6�'����ݸ�.�ןmɎ�\#�ѽ�
�'8�j��j%y�[��뵍��[�#e��U��h�DvuKҩ�k:��\���]8�e�ۍ�tq��c<���W �,�T7��c�M)�LM06��K��k'VP�;�t�y��"�/k���ۧI�]E��=�g�p�]c��%˞vRB��NW����\�\����c\;1fJ�B5���ݭ7��h�:�v8�V�d��ۊ���Viyk\�1N�ƍ=p���l�<�Z6���E�T�cJ��S�P��IZ��]����gt[�m�n�kͺ��)�ə켗\��uZ�T�X�i�/M��A�6�TU���k�lxsF�Í�k3�ԏFK(Uݞ�E���͐�u�ч������&�i�����N��u�o9Ϻ#�=rg6��I�,��y�<hD,�m�>uJD��V�������3l�M2�������5]��Me�V�n:Tb�d�ߞ��^����$�`RT(s`ڜ��.��U,!�ޑq[]��mZ��(�C/����l��Jw��#�3���f%�����4�5�	΁z��1��y��Ϡ�@}�"HFpz��x��!':�΀@���@��||Qi9<����uD���MZ�S��
ȟ2 �׈>)D�(����6�'E[� ;�����*�lS����|���3zA"���������ڳ�k�\_%����ub.ң���U�ڈ�v'�f$���V�6r�7Vy���l��<B0AIP�5��gk+��_{F}�b�۵u�����s%�8ݖe�G���]�u���02`X^9BR'�� b��ޚ��u���\��D���=uz4M-�A(���AIH�C�����N�ll�Y��5�qo!�L��fv��[2�$LT/��ɜ�rH2u]\TF�3��7&а`��FU��;�X�,�j�6ɵ��]'�rXC6f�r(��.'vaq�p� ����v$J>IM�|R�wu�þ�|����K�6r�5��� ]�+��B0AIP�BS"UR�.�/�����ΐv��7��#۾꩚]�8U��>��<o�	"���r�>P �� �"A�
k�tܠB{B�6�9�ˤ�Kf�H����,�����w�g<I!f�H:I�>�7��o���sqo[��B*�5t�-�\�B���j�������K����H��� �R�=�ܔ7��ʼֳτ{N�D�Y4�R�r �>#�RT(�$�BB�ɣ|�t�J��~#6g�DOs�UT�:�3­\��x�D��Y�Jbcc��<�3����@'yH��	!@IW��J��s0��c w����Vf�uOa��3ݻE�B��8��U���tG7�,�m��]#4b�3[�mJ�!��7[WM�Y,!�ސH� ��ݡ^!)�Q�Jl5<�	��F��Z� ����� ��I��ʽ�7��Uy�g���0����3q`@�>�^m �!��D$���ۖ�DF�vb���[��Z�S��2$�Y
Jh|R�����?o�����������G-��f:ť�$؉�aۈ��y֕u�q��u]�[�������2�G8FIH��a�|��C�Cf�����}e�f��1�����S�(�24�L�>���橢:�^��^�7��uy�g����n���'�1v�Q	O�C>�$�Q��Q9�ob���R����U��<A7���$��A)D�|��PY�b����AȐC>��
���]49d0���@"�p����Yrg��A�)�ض-j�� ��T��r��e�7�瞢��[��%�ũN��v	�U��M̨��ݔ%MM������M����7�ބ`�uh�iN��yݻ�'8\x�w�Y�Xզ�ky��	���ȐB0AIP�;��H�̵�n[��wZV���x2SJ�.܍���v�t���#�%X�˼(o�r�,SM"�����X�3]or���<��;V�T�NŞ���Z��X<}y�~ ��H�=IH����Z*غq@i���\��.֪Z�CT�`���(��y6{�~��Tu�^����)��x��׵Zl��m�y.�T�4���[�/P�{�dFs�Zm�{�	�ܳ��w��r�hG�2���@�Q1���1UBy��v�L)�|o"|�{%M[�ZH�o�� ���
��)���!�l.9�!�U
hpG5n�S��8��$��"�	L��Q�ew@��g�x2���h�n�n`,�<V<Q*���j�"N��6�������f���}��s�z��Ǉ�Wb�E�[����X�۳���&�z��7���|���r+�\z螌-������TSl�7�t0K<rku�����s=18�t8N�ѯ\�����rE�aa2hXR��f�h ��ZW6��n.�}n-�[�1��[t��ܠc`� :�;b8�kN�F��=����[����S�i�M�n���6����;�3�~����l�H��54j]�gDj:간����ݍ�B]��ݡ��#5EB�}��I��Jl	J'��gkP��û�k<�@y�\��η;B#^H7dhRT(��#E�����ڇnD��D{��R']�'n�q̉ �D��3��ؐ}� �nER�$#�������%���w5S��8��$0�ٻB�!)���S`���M'�vDb�A� ��%(�Ν�Ztv�/5���5� _�T;�}�x{6���$�P!.{���9n���"=ٷ��梌���ژS���A,�%7�*����`��o�_~�dY�|
C7B���&w6������,��m�Ύ�#(h�<��m�z2<�H�A�$�}	*�l�sWkU8�#�!�ޑ�],l��Q�c���A��РBs>%))���˓L����D ��
᱆�y��m���W�2)��#���;#�]�8�8����[�E(ъ�"ћ�3>�ڈ�Dq��'\Hq�:���-�fkK����^!�	"L֥�����DnЯ�@�H�䔋 ��||Q�SF����5�!�@��k�۷0��#�dzAg�)����|��s��gZ�J5H`����A�J�l�s�kU8�#�!��	`��3k.��D�``���∀RS��J DP%-�P5S%k"GE�S�Ǝ��e洽dp5� S��U��>�K�@��q2�f�fśi] �t���z��U��������t��C����g�Y|��
%"|AD@��J�:�p;v��"j�Q��3sjd@/6hJQ (�J� ,��"{�G�9�B�2Q\�Z���V0��� F=�@�����zr�"A�S@�Z�IG�)����5�?��`��q;��+\��^���	*��}�Esu��Nh��w���]�|~[�D�f���d~^f	�����oW��Kj�{<��ۗ=:����1z̼֗�� �}"�#vD��A	*Jdo(�VJ�����
#�}> �"��l(訉�k�۵*g� ډ!!�B,e##HE���q �D
JE� �WR[���P��JP�n:T�N&��A!�'�+�-��
3H�+�ya�.I����9��w�w�<�6�{@�Wnj�$G6%t4�3hM�ųN�t�q'�D�� ��\}����E�n��Z^�ꍾ�u�[��8�Ȣ��B0BJE� ��
���/&�nEQ�������:D[��W��v��R�}�ډ� �D�ʘ��Ɏ�P�l��U�v�������B!��Eb�̊\{�j��7��S�8�CWH$# ����$D��"܌�J�؄'H�iO�����{�E�t�浞���R���Q�!,ɽ�V���d�����jS\O���]t���?/^z���+��z��*Z�7}�����b͑�{�N��x]&���{J?\՞M"Oox`��؉�����ˬf2�r���"��%q���k�ۥ*g� ڏH,�))��.vhx�|�g����p��&+��:ѹ�ɤ�9�f{lk2��`vԗg{ߢY/��5���2�`���2Vl��t���Z��Gr�ÈTwV�͐kr�1ǧ�$��%(�6�C� ����"<'4}��;Xb�Kj�^g��k�� �vD���كT�¸ܮ��B�̂B0A�J��� �!VW7�!�lnc��t:1]Mh;t����I����J$�;o�i�[cD)R+�!8F��%B�L��S�uX�-j��4\�#��ۗ��1+�a���t�%5��A�>IJ<4GB�0h/�6��ŋ�+��_@&���"A�%B=��IH���������s�l��c��xj��Zt,K���=bk:�:�Vm���(�}C�����q���d�A�Kw���a��p]���4a����w~���;��fP��^5�3[WbK LG�Eҵn*�0��\dPRԩ�f��3��鳅��$�v't�݌Kj w�:�jh�k4�Ò����l��;�4x�l�mj���ꭷ��Z⸒Ć��BX;��i�P�M.3	A�ci�<h)6�G���m��t	0Û�֬�ұ������ul��$�Z�I��4��VZ���b��|���������n�X������ț�����BxEug/TB�"��R��x�%y����s:}E(�(�JEn��Sr�`�`^:92WBN��[�)hCW	�h�T��w V��H|�Nx������� �(���y�7̸�ó�V<�u���W9;�$�`��^!)D���n�Q���z�Q�)��{=∁��4R�+�8K�S
{�آH3K����ݑZVT�E�*ٺ(G{ݘ�vX�t��چ�!nЯb�+a'|�q)hCWH!6�&��0M�ˋ��!�o�9��G���,ea �)j�x��Ѣ����B'1�)�{�mĂ	DG�dI�ds�U�7:'1f7Y��ph��A@�sNg���`�T+���A!�6��m���U(��͘,V���٬zU����F���2�2��326�X�(���������c�$�j[����sؼC�G_�	��x�S�>>���i	���Qۥ0��J$�Y⒚s�Aӎ,�F�$�`@ �� ��I� ��J"�y���
���9w�JZ���vE BQ�(�%4E�x����kc"�S@��v��s�nO
��5���=\�Q�jV��#9���Y�Т�H$#�%B�	^�xӴ畔ug�"kJ!	���Qۥ0���zAdG�Jk��A;n����Y<��Bh*"z�We��6�6�V�cq��-����[���TE�:<��QT�# BJ����M�9y�JZ��C��12p�� �R�DnǤD���J$�w��vi������^ ���9���ܾ��N��G]"�:�H!��!1�1�˹��tX�i���&�e�v�;^���X�ȼ���Z�h+ʊC�n)�������Pz=���Ѱ�������:�UFӗ�iˇ�N�BJ�ѯi��ŲOyϑ�q��h����nخ�'S9h�D�ZZ�㼡�B� �3aq��[���=��I�*����ʇ*'�wu�5 i�Fl�9hx�L�]��^��6Gw��q�e;x=�N���SrBU~�����������7V�f�X�� �;5�7"�6�d�N8:7~�AQI��h�{�C=�MɈo�k�\5A%��2����s�nL��5�	��%���,�7��/{�<<B^o�P��=�ہ��&L)�(7Og��w��r��7�_/m��"�������M���A;+��կ�P���P;ӷOz'S��^�x��;�s��c���Ǽ�\g�gE��S��7��7� �3�ќ��g2a����}��d�I�]<�'w����vI�D���WM`�#��������}�j�-޲�A�É������t���x}�ӠC�Q#��nS�w��Ѥ�"��.����sG�?UB�6�٢-��[�����D����>V���C}�ȶ�٧��]LD�|=�������E�b�)�W*�C�aNs.Us��R��;F�=�#`K�C��h�7E޼qO	��?$r���}�Z�3��>�%^�F>�q�u�266����{�%�.�ݷ�_e6;ȍ�cé=��t���%���ŏ˥�M=��~N�5�`��<7�. �ܒ4���Ʈn�X*��/V��� ��Μ���Ӝ��+k��:��8m�)�G�	$�vvw �Y��qpD��[jA!"8̳9$�%8#�m`����K���gN:Y�)���8	8�[����!$�m��%��mi$Yb"Y�Q*H䕵�prNt$C2NNӔ)kh��$Fݢmh�:"$AÎ�w���αP�����ؔ�9� ��-��D�Km.Nf����H	��	��A�9aDe�e�#�D(��*C�Չ��m�.˱�#��p9$�����P�H��V֜�u�,Y�3���G99u�[rH�M�qY��BE� D��6�(�� H�$����B8IkY9H��QX���XR�9���}*�w]��m(S<A(�2 ������.]nڼ�p̩:�H!��%B��X[	��o3�KC�H$3 �/�����h�F�$��A �A(�))ꐎ'Vr�;!�eď>�;����
Jާ9�>����D���R-k]y�������l��a��l�1ݢ����pݸ�h��t�ٷ=�il�a�1�C��Yg�u�Ͼ��BR'�D_7�B�g+�b�i���ul�Q�x���P)@
�
J@oc�^G��0mN̉#�/vFic:1R��g��5���
{B�K9�߷G���A~�z���V#7R��w����Dӎ�}��
����V����g�&�H�uȒ�y%@%�M��]�#���]ϟ��
n����|!r��+j���2�GW^��a�y jL�Mf��h��!I�������]5���#�j~�Ŏ����p.I+�7��
��[�oG1hQn�J�w��c��y(���s@�V��))�R5���4o�t+�AMK�5��
�k� ��{ $�Ģ6��N&[��/��k*�� ��y�������3uvJ�|��9�k4^8�����~�z���V�Ԩ�)�|�K�Fn'Q[|),�N3���z�W2�́ �`���@��h��۬��sD��|vO���O�$Aɭ�7�Nrg� ��> �ȀRS�S˚�T.��^̀G��E��!%AV��x'%W�̤j�z��@f��
!)" ))�7�Ftm�]���"��(��Fn'U;|%-Z�g��it�>3*h��Ի������>�͡^!)�HF$�W�HŎK'k	�w����5�p9��ri��ڥ93�JȒ	d@))���75�B��S�h�Vn_d*����t�P��۹\;{U�w�,:2"g�qri7���ݭ��F��)*
��՝�W�J�D��i��R���@(hF2-!)lo�yob���thc�k���ӌLJ�t����qܔ�Ou�dR����<Ը�s��;c]�e��� n�t��;�8���8�3� z9=���&a	ef�b��0�t����Vr�]rk���ێ).�
u�t�s&�[]5�=�Ɯ4�䋹h�AՍ�md1�])v����7ܮ{5-�~��N��-�Wha016�{g��y�&�A�5˞����͖��Bl�o{��Y|��7�)ȟ��$�P��t�-��v�C;�B��_���f`��׈�y�0Oz���*;���Լ(��W�e��_ys�{;�f�sS��Rש�z��K�p]j����~u�Y�0\���m�|���>>(��2��<%�sO��j���A�� ��#�%4A)D��vl��"��A�R$�x�����t�T���A�����C0"aT�����抿a��j\x�;��dw��Dv�
Jk��U"",'ײI�W_E%�[��p�R�B�W�J���'uG��~Z����6�U��(�"s���ׄ�66m�Nj��
l��=�cL������v�in�H�篫cnT����f�i�x&�H � �S@�
P�IH�&���l�^�1��N��'�B&�FwpV��SẺ�h\�O7v�m��f��	�?b���*��=�	XNcM#�%ő�;���O*�]�ԚZ[�	� ��hQ	���n�`#�@;�4A/�O�RS�"�(vR�f���gx~'"������z�g��z�H�["A� ��Q	L�����:'N��#����B���> �-.�0p7=�[;r�&x��I9<Ho-<� ڹ�x��x@%% RR7�JS�
������<jZ��ܵQ����	�{B�J=%�<����=��}tx�ڦc,w6�ӓ�.j�\���9c���f"��Bj��ߗԲ������G�IM	J'۲3q9��镭�g=\ VI��9S�"�>$>��
!)�G܌�[�Fpq]CA������n{��v�NL���H �D���O��T��y�#��"�>J@F�!%CTUYC'�vd�
�75�۹Eœ��a��R�n��nm��F��c��/nЧ��,[;e�˅j��m�BV+)�ξ:�4�����I������������f��Ϡc�(�D��]��-X3��#��"o��R��3oU����ֳ��5�"���o�V�M�#19J@�A�J����$�k,BZ�D �]�{
2d
��%�%4��E��v�x~>hn.ms�nٍ�^�����앺�z7�%��=����&V�jR~�b!��f��T�w($��|����o ���ȵִ#d����(��IM)D�_E[=B����'�Fn'�u}p�Ǭ秄��+d]���ț�P!�� �RT(��|AD
��*�{���LEf֭�s&�kr�oaFL� ����D��R� �TU�1RؘЕU��AnD��1�IP��<�<c^>�!hc6 G�D���;ծ�������N�l�Z���t �f≹��Bɖkv�2$fC�@���#@�ܙ4�6W�6��7XCԭ���sm�#�}>'H�RS@�
Q�(�))�0w5��ߧ!>�=�z+/�m�9�� �Y��'�# ���Uz��M�o�<�[.4*#-�c��7:�=�݂����+�^��l�a�ST����ϗ�>��{���
"���8�t��N���/����UF:Dݚ>J T ��@�'9oyV9��}�?�<�
V�uP�Ƽ}X!hc7��Ǵ(��4)G����x�Z��J|�J6�&�z0��le�YM5�礎5}"�+dH! ��Q	O�����B(�N�W�JgĢ-����Ȏ���њ�T���{j�F��q9y$@7�}@����Q	@�B8d0E��5����VP�����B��l!�c�BS> �23s_�k� ?]U��7b��Ti?�Dy��ل�
��3 �'�����b���/�b�"��4��x^���w�O�_���ߵ�<�7��6�h,	to%5�6�B�0{l�e��`v����|��ےU���d�e(��(�]4t�����mҧU$�v�ȉv&�J�
qց�7ҜZ�ĳ�b�Z�J��&�]�rs ��]���g -�� l�3ׂ��g�;���V1��X;��m=R�ۚ�	Ǻ��>���t�0&�y�K�]�;hƶ�kI�{�����iv�0J@��<}���Y�=��[yY�qgT#6+uź>��_��%��������+;,�m�9�� �=ק.�ꑀ��"A� �%B�!( �w���7�j;��3$O��#��|
�#��3k6Td�x��y��Jr�󰋸�@%� RR$���g9.����F��svoj�cm���1��0A��K����RS@�96�k��f�Ȃ�MJQ=��q�՝�V6�����M_H�&��#e�<rqpt���(��z�f<AmЯ۞9����\�{��k4ȍ�ͼ�Q� U���'H��� �ܳV$+��W4ƌ��ÝI��2���v��,�S\j��w9f�Q^2bVVљyUl��u�Y�w��"q�x�
�Ϊ�m��B^�3g��/h����� .hP��5�	mϮGU�6�;a:��\���ޛ��MX�ɂu�ņ��f���Ъ��5��)�A{��}�NW�V�h�e����S�@eM��N���C����+z�zH�W�(���Q�3�6���b��H�u@�8�t(��
�,����4��j��ppr�3�kU�93�o:hA�����nh�Ǆ����ƹ[�K�Gz�l�܊����ص�hK��l�A�e9�����=��K��|YnhAm�|Y[s4���`9sc
ڜ�#�\���*�z�zz5} Sޠ�Amз��T��{�>�����mYn�cLGQ�d4�;�j'�$��,mM�;6T3�Y�侼��[=^;翴(��
�,�ץ��<oZ�v�&x0A�f�bu����l�-�� �ۚ ��6�n���+.��F�Kv�@e�[AӍ��Z����%�b����c�Cmf�SW����<D�4 �5�,��m�	m�m��]⛣�0MOM�Q5;���v�3[���կ]���8e��ߡ���|/K�ȏc���G�4wQ����)��/�p%���z��oVf�[��w,�m�9�� �j�Ex��P!�6�Q�,Z�إ��	�AݺO��|Y��A��<oZ�v�2}�ΟQjr�����䔱�:�h�Ǡn@�ۡ@�a1��!.R��Ho�u
�q�.��E��B^�-̎!�gl�!�^�����T'��%z��Ý1e���������v����RSQ4�V�E��j��s++����s%9��F<nky��;��ESoY�OUĝ{�:0.�>��� �tm
�3!�L�y��R��U!��g�"<��Ay�/�Z�k&2x@7�>��Am����;"��rF�w4�k�D� ͐ۑ�':��V����)ص�pK�Ź�(C1�vРCn�x�DۚL-k�6�m�Y����"<
}5��nh�\V�nOeM��=$q��E�%w�84�C��䢱N@�ŃS/�&��������������	�;{*r_V���k�t^]d9�YmA�6��"��D-
���$q`�1�
!� 3d�
���h�Q��M9��K��KK�u]�������A��}�@-��|ە���������Ј�c�uo)k��,�nK/X�3��tvH��̺�k������Y�Ƣ3�t(;q�;�Fͮ�0�!jz������2ȓ���D.��D���nk�^&�8�-�{T����\V�nOeM5�=\#�� W��
!�9<&M�i#bv��H�C>�� �B�K!�ʇ�ni��k��E̪gBs]m��Z�L\�Du�בz��Dy�^8˶��C�y5�!�B�f���V��y�6�)OP ���+�g!ם:��dx�󜼈��r�"<Js�c�l�k��8�b�0�hkU�[�ܣ�7�����uf��p� ���>$$ I?ܐ��$��$$ I?�HH@�T���$�2BB��d��	'��	O�$$ I?�$$ I?�HH@��HH@��!!I�BB����	'�HH@��BB���$�����$��!!I�I	O�$$ I7$$ I?�b��L��n�z
i�� � ���fO� �)�                                     |  �                                     ��U$RD�*("""@�U�U(QJ��T��(R��
 �)QU"����$T��T�E*(|  �R�%H*����Q +��}���U��ꂪ��T �Cz�hp<����w�� n��{  �tuJEV^��G{t    �  h�c��ɠ�x�En��k�9(떀 ͊ 25�hn�*�8zw{�`7�w^�ػ�=z�;��� 
  �  |��*�(�UT� Q*x��ay�ފ,����{�y==��m�y��x-����k��:h�`���(gTT�:v@�    � �`� Ϣ���R0� -���� a@�(*�  �a�= r q 7�  �  `   � �W�����
(T�UT�����q \�@��O��*�,��� m�����*�n�e�Ч;    �   �� >G�uP&F��Oz΀-��!�w�9*�s�]ЯmW�PT+;�BUy��F��ꔪ�   7�(  /$��A@U�Q(D���.cR��/�W��B��	�J.�R������]�tEC��f����OZUC�
)�
znmBR�{��   �>� ���^ڈ���Jt�K�P��b)FZT ����H&���*;��S�zЯ{u	@�nDT.��Rs�\�P   �  �� �$T�IB(R� KީJ��E(�
�-
���t;j��J7n�z4s�v�k^Z����J���UQwJ�^������   �  -�;:������;�"����z��w�=�-����6��:=�TK���2����y؝�9�����M��R� &LS���)J�  ��R��$���M0�d�%I  ��IQ2��  D!�R� 4cS������I����A�!$���}�F���y����������	,)��HH@�� @$$~�!!K�I	_�HH@�i �HH��?O��k�r�����0?�ץ]�}Ru��w�ϳ�Y{��i�"�/&Z
�'wT�cnލ��Kچf��{v��5�7����Kn����_*6P˧YE�!E��ED�`;�LfW)�ҷz�^˒�y�U���U�Jͷ����ٔ0�0	l\�B�n�`�S=w�+E�4�T�-\�)'��3��e�����Ool�Ec�w��]�[����xq��H�W���h��d�c�
n�9�%^f*p���:���UaO,V�/%�Y_a�����VJ[R
ڸ�Y�0��=ղ]���n����t�e��f�ҷ���/]�R���W��7�"�5�^�f��U�І����^�H�:6�;EBf�*��*]�[Gd�ѫ7[L�
h�Ҙ�[D����+��	H��wFd:�b�qT�[�6E�T.d�UE��NMZ��'M�P �/l�IH�f^b�U�F��:�V+wU`�@�%cV��V֍�fʬ�܅��j�!@�X3(Ì'��mKL��34�W�]Ɩ�n�Ub�E�{eZ�5S-EF�ͧ�*Vpdw��CN�1ŪU����x�;M�%k4!v�Q��$����d�6vp��������6&[���Ib�����"un�[,�{yv謼���V�+ۡ�-U�k3N���V����	J��s�`�*�̥V�7V�۔�o6�򫺎2^����A8R�6�^�Y%��Z2�"���4�n�[����j����@��#8�b�n���(���k��}-c�ss�mV(�fn#�2�osH�]ۥ��2sV�j��m�FT�բ��f�l�7.ͯ���BGA�&�˕S R�BU�N�G���U�����Y��h��hH�LP�[�V�eZ|
ӹ��J�BF7�Z�J���Ⱥ�3f�n������-k5k3n�[���-�ef����uZu�����U��ac�Z!�i�Ԫ�L���k�w�:6�l4���U�!���E=�Xt�����a�T��L�[������;	8c�gvU���mP;W�Ew2���\�N�뙅Y,�R<�㻊�]�z�L��뺛��2�VEX�p"Ipn�F�nV[��̻'��I�]�����KTܠ7�;�Ja�����i=8v�=�U��Е65uLR[��%ڒ��,+ǒ�2�KV���h.��n�U8�b�%����DM�w31���{�5�̀��d4ol�B��B(*�LD�x�f�JH��L�Պf�޹f��z�Kv9f\F�j��3p�Lw�ؽ��ۏFS��v�׉�Yj����dۼ�,]]B]���D�UyE=�h��h�U�"��1�q�LV-�Ef'[Z��AS�n�ƠW����ja�����mk{)�Ԩ�&�YZ���&���ֈ�&�C�X��դ�۩y@Օ�S���Y:�ӏv��֌�:*�h�
Vq�ch:Mh��n[*Beg�tY�������;�n��bJ����)b�r�aJ�R�$�fBH���6�Ð��F��Z�%�f3�M��'r�M��.��v"sa?L8rZ�U_X��V�/�������e+�Ы0��w$I�2լJ�m[�����&3r�j�o2�AQ���F��(�4��l�C�ɔ�I�X�5�n��-t�*ZN�A��6iZ�hʊ�����\�JT��޹�Q�hùK,�S(dPK����Li��U�&��f���D���͑G�[��Z�bn̡mA1��**�U&`�/lfc�hh�W�Q�ޓ�S
R�iY���b"��Ȫ�s�5jG,����j�Dpн��a3EPܺ����`���e�YTc#CՕcEhƩҽ"LJA(�f��4���N���X�7f���3e^�TU�m��Ea��[���E��sd��+6�d�_!�-ӻ��]J�W�%<���eh�`&ap�P�n%F�P$LfV�;x4R�kF�K��.dQ�V�UƖJ�Yv�'j����*B��KM;�G5�R-uj㊎��T�e⛕+DjbNҚ��E����M��Mb��f�Y�z�u�,F�Q��wn�6�#���ʼܚV�c9�E��G�Y���&V^`SD��v@����z��x⽢�1|\��nnZ�8��;��6�3�e�W�
'.<Y�ټ�q���ܚ��*݄Nf�
�0�1^--�]�]�nk4sB�ث�TΫeRz���bU�v��ŕA���~�4a�o
���J��Ҩ�2��ݹ���j��N�9�"�b����*�뻗�U�t4U�eZ��yL��n��J�Cr����6��R���i�.�t�+XD�lb�7��)`�f�ˠ�u�o��*��ۃ�ysU�y��.�1�j�ڧ3SZ�)���&����i ��g)]�Α������w��X��˼�Ř�kEV��n=�����d(�m��n�ڸ��6Lj�eV��sf��m7�W&��9Fӭ�1&U�U�%2�%��:�z���n��/�ఖ��e����%���%��EU�����z�4�0O�dܙ����5�N�Z6�(�D��E��5P2ݑ���U�:	�V�OY�X�.�5n]U���sK�wc!��o4���WV+j��J�H����&b�W7x����2����f��ًf2�J�&81�(V��*��ݲ�^nZ��Y�F-K��6�f��x-�;/m=XMj;��5�+mQ�p$�U���У[�(�Ae3�����[{�FT��e���yp�'ql7wu�Wb��L�F�n��S���V��-٤S��e�V�C`x�Xݭ#nkT�P�u�VF�7SnfQ�;�V�Sm�~��(9n̵N�NƳHrS�٬��6�V���Ubf�]���Լ�Xc����.���T�4�?��?Za���Y�ooX�ĸB&���7[�0�[	8���D�m^�ܲbbc�&�^��7y�m�$c�Z]RܓY�nг���u�MR�Wy��V���å72\V�"��1a� 9/(ݝs
�[���3`R����V	Q!MKf5s\�eQ��ص�H��b�9��<˸�i�"����.�ⱴ˦���x�r]�F̳ ��������30�d���k���e�P�6]ˊ�-�m�%'3qf�vi�x�E0i�v�J�9vK��y[B��De�PT�U�آe����ZufET ��ʷ�ʷC�6�n��N��,��������Tl;W���f�*��}x-��t/���tZ]�Э�4�%Q�r|oi�q��9�ܬ��!�Cp�e�TC7��#���6M��;�(e��F�Q0ػ�4/A�vLᏝd�S���,M�0���v��Zś�ћJ�T�2��u�_b��Kܸ�~�x仡N�H+c���/��D��2��V�h�Q:�V��X6j��QT���SZ�]Mw�F�����w2֛"���kf�Q��_�Rb�Y׸�n���m�D�7�fY`Ԓ汸V
0��]e��b�+��I��ʻ�,�UB�^����߮���������Uj��wSu-��a�ҋ+]e[���+i;h��#,ܫ����2Lz-M�b\wf��3i�,T��T,��6)�����sj�U�;2ݢf^e�TN��Bؙ{ʑ����1��%؆�9�|ԛBH7H��+DX��QXi^ǲ�g�v��
��*��;��k�ŘmVk��;P�ӹ/7�X�����
���XnLl�?^n�¬V$�[M)T�l�lҮO�*Wt����kP�+G^=�Kjʭ;-Yq���oN���"g1���R�v�[�&�&)[T�r��w#"���'�R��2fù
�Q�ŘkV!1Ϣ0�cMe'���-+�M1ɑ��YNj�u�J͆���x���6�+�R�r�f��sF�OY�Y�1��I�5��v�YR�j�V~����+2��ćP�)��wJ��c�*�J����G��%�!]!�)^j��X�a�V�v��.���U{���K*Ƭ�e�Kv��m�ǎX��Y��~%=Jg�x3j�ͻx�̴FZ�~4n��YB��.n�Z�q`)��2��Jϛ�7�'�I�̙[�k	�z�p��Ij�5��r�0�Cs(�&\Vd�x6�c�t,��*�Q]��%QÕ�r`��X���UV�פ�p��n�-�� V�W�VU�v�f����D�\e��[�7!l�C��1�R{w���ͭY��hPCN�+Y7�y%�b���m)��{�$Z�PwSl֜�V�0�o볹YU�-b��}Ϊ�oV2�/��.�̴j��o6��B������VJGf=:pkX�X()�[Ö��u�Ggl����
-5-�v�۫�蕴%�W�e�::T��"�SD,��P{�H��7iE����&�w-��^-aKV��Wyu�V�CH��G2�YtĻ��K�Gf�j�T�&�ݪԐ�`MR�z�d�+b�P���w�7�k(����n陳v�Z4S��e��{�����M�� 4�/57��Tƙ��6��i�s7iZ���˵q]����P�oy�%���BX���̈́l�іj|Q�k6����3��5�]6��R��哒Yu.^a�;lV��4�'Ą&�;[��̧�b���,�ˡY)
�*@I��^=�٢�ˁ]f���B�a[���:t��{���d���FɊ�aC*�v�M�,�֊F�j*^�P`7�7�jʭ��h[uw��4V
��Vf��V�1�����Y%���Х�ڗ�TvPx.i�@��-:����8lSFOv��#�Y�ZÔ��M��c�:d���fPe
r�Fr���r��O^M�4-�S`7u�7o$��r��e�f}*�a�\5�q1�&�٣��T�U�;�������1�cw#���b��<Vffݪ�H���In���{U[p`���)�Tњ����LkbV��3E�w%�A�N��nëʼh��s4@Y�5�6�Fe��&[W4P��îi͒��5�3Y���ZV���z��]��[�p�i7T�׫6"����6�O�:g1��r�6�S �R�4��7]�W�)!x�H�z�r�۶�a���uV	n�/��*���T�M��"YU��i2��[�E�3�i[�*��c��[Sd���E&v;�ݔՖqT�#hh$Kb��w�U�j+�Ӣ�fY�?c[.Дc�qaQ��m�l�M��%Jo#wt���W��m�j�̘��:�1mK�nn�X��@��R��L�˛m-љ�z��A�b�n��u�j�,�!B!���Rn$r�jP4��!��]�EK3��a�	]R��r�eJ̹�Z�;���V��ۢ{�)��gF5��af���h=a��*�a��[Jn7�u�U5f�UDRA�B2��+�O4��5�ӭ���(fCdԄ�����؎[@��䪐�Wґ���U��QB��əe͘͜�J�;�g�M�$�#35�p^}"4�-��(��L��쇗A�0ae4�rfi���*�8.�,��X)IU���VMlS0�l�N��������κ�2f��̲��0�mb��VM�7�1y���+*�N�[H�/,�V���m4����4.�)C��]�ǃ+U�Ϭ!�m�i�&mAR�Y�5�ӭXtQ�n�p�i�.����
Y,MT�+����
T�U�Jt�]شs3Z8��l�ZS����ب�ܩ�1/��w�ڼ���PX�/M��Cn)��S/��z��m�]S̵���t�EN�^�[)��fK����/m�Z�푿b�;��j+��]��f˪�Nd�c�̕�k�r��Ei�bk�/n:���њr-����Jl)��F��mͱR�ѻ˵��)V�*��m]+aҢz����q�d���b��-]U;��b� ���x]��*�6Lm�Ө����ª[o3(Y�Wyu�]K�Cr�wB��!���1��%Hi�dm���
f��#go�/`�
��+3.nľhW�i]lX�9zm��B�`{Vj�C�L�P�*�fZl��f�֭%S��V�J̻g�P8�:Hjܯ���1���������3>���S�_��x+?K��U���o.�m@��w�s^=ȍ	[*X2+��T�B�%l��I�����AFk���lU���h9S��$���5��+�U	ef���ej�ݖ���T�Va�Be����wF���N�31UM��sU���ע�ϕ�j[K�i*Yg%B���r��]��ikT*;�O�RZ��k�&�T
Չ�U4vЕ�o7)�uO2�S�F�<�nLI˃h藍���Y�.��V�5TBy	`�N�͕UQ�yA�ef^Y4![��ۻ��"o�)M���5C4��+�3)�&[��>�Ri��F�Nb���1e�{u����h��v�Ԉ�d�wdiCP{���a(��ח���
Y��'^�3��K��o��R=a@��.Z�e���fni:�
G֫DhF���oMb¨�Z�`��Sl�URL�&�����Ct��y\�)�*\]�7AZ�Z��*�N�32�l�˳u(�Q��ܣ��y�!U;7U�d6�3T��m^h�yx�Gn��̻��m��R����v�%]d^oكc	�S4��Ӭ[e7i�݇���9�Yل���՚����ߠ��j����x��j^;{%Q�+.�غR��^���WW1�y"�yi-F�+�������m���o��cNV�n'sf��$@ٺFD�m6��ͭ�[���XViV]�]� �u+N�f��yj9gb��-�o4��躵�(cE�UJ����͙�GX4)�+*�b�f��Y���/D��J9Z�t�O]���-���������edhԽ������qc��71b�t�H��t�ö�/���t�{���t&�RxPTr����jiv���[�,�X%�'srP�/e+��j-P���O+%j���r�\u�U�ڗY����hY��^��[n��clm���U0�UN[�#U��2�D%b57�/��vn�0s�H֐��� l�����*닺������.늪;��������:�뻻��:����먻�+����;���;�����뢻����;��⻮���:����:�;���.���뎸��;�:�.����뮎����������:�:�������.;���+������뢮���;��.������������������;���.�����ꋪ���:�;����:����+��+��뻺.㺺�����㫻������:룪�����@� 6 o�� ���$$ I^խ#����~s�A>�<v�%�=|�ݫ�>�T�=�l1���r�i���]@�Tp^J�ۆ��>�NnV��p�וw�&^�m�3J����t����#=՗���9���vQ:����W.�A��j�J���W�"Άe79��ʮ�&�Vl���}��a!���,�k��f���	�j���n�����=�mJ��l��1u�n�/�9*���co��[?wK�t[��<�%Y�2����n��X2�3;�5��X�6�:s]H�v_�7r�~����do}���'��3��>�9Qk2�T_t�N�7�.�עԗ�D�����2ɤ_]�&Q�j���1gQOw�=�z;�;��ɰv��U��e˺w7�-����tMT�WU�iLg3
���W��������5�t�6��a�����n+c�-VEk����v�^*��M��+ӥY4
��A�"k���v����8�`v���f�(U&���s희nQx2P[C�ְ��2��<�+�w�i֚���]Sk�8j}�of����̰q2��O�QR+ދug�j��q��X�J_`�ׯ6]o�2ɸj���w��s3ήRU��l��
�1�-�*m���8w.�2��Sunqd�7F�|S�l`�.��}�Vd��黽̺Y��n�-���_�r�v:L��~���x��5^�zA��S�hr���-��`�-�������a�p*�쭇w-,��x]��U�ÃS���3F_T��Lt˻hi.r��7$���˩V^s�\f�+��si�GY{w���z�����j���FSuJ�Z�Ӝŕ2��9q��pv��マ�3�2�C�aq��=���d쭺i�����(6KD�L��՛"��Y�ׁЗŴ`�(�Ҽ7�9�Շ4k��u{�6�n+(�<�2��k��|�oj�KoL���:j�gv�:�pb�l"�DdKs,nbK2��6�+\���Ǖ3�m�<͊�Zй���KU�N"{f8�VK�V(fƁ�����E���'�����2��ݗ/�$;W��vT�/&�)��n����T�vB͗�hu�����U�ʗch�3��Ne����	�هz���{l8��i�2[�Y��nhT�6��Cf���Vn�NY�ΧuQ�.�̾��)(�V΋�������>�\�l�RS�8�4L�5�m�z����ݫ��.���aL.:�����F�ը�ʘ��l��(a�����+e$�!�d���^4���z����c�wCxs�_Ugs�q�v���P4��]�W�*��)fҠ�������m�Bg�]Mkj��`�l�Pv�WI=�ɾ�b�$3 ����؅���pv��1��u�����Ca���[6���n�9��Ƿ3\���f�3jZ}�W[f�*�b�R˾�N�&wT[UM1��h ��Pg>��]�f��]av=p՗]��k�-	4�l)q�*�*ܻ���w96y�a��F�Kxj��oj��q��M�),5}���po����iO�Wu1t#}UH_Y嘆�[�J���0�f��|U!8��n�ӻgsm�8We+��Gr#*��U�2ﳸn��k+ �'3���r��S�_R"�sZ{�/s�o��6�j��V�����F[��n�s��,�t�J�vI��dIm�p�Tj��z�[�Ӵ�"�'�$'�����.�-:8&���
�Ń��f���Ś{��S��w���4d��ޗGj�V�ו+k��75>�%ҏ�t�u�7�l�ҫw5�.oز�}��2�s[�6�<����%�SO�D&
���������YJ�����䬋jŖp��yw�~��6Z.�����A#��Vr��f��գ���qw���\�6�#��6�n�k�\���vkԬk��t4:?<��-T��h�]�8�X%�# ��.�K�V�b|\�d!��H$Z9�VMP2�&���С#9>&��n�������( o:G\]l�co��lņ�'YZ���8�ȴێ����/�;�x.��Տ8��\3���펡m��㘳���Ӗ���^`��͛zu�[m����w�m.)��:	��Y;�FK�T��*حr1�Z}y�.�wK��u�ڙ�`��1:?R��K@���g;���ם�O}���;m����j�/M�onZ̛C�o]�NMZ�&����x��u��������`�wy"4'j]�2���#_װ�v�k���:��%�ۻX9�r7q9F��kEbʺ�GN���8Zݴ��G1�GN�-e���-ں�K��n��*���hp{�2wZ��F����V�-X룳�h�wu�6n��v��vr��}�ur8F�f��i5bgVl���=�yԦ�>J����3��sC.��,�V�v���V�|jl�і�;[�S�Z2p;{��B��曻���e�*<nK��8��ͣ'M"F��I͜4uWi(Z�:st�*�qq���&]>�z���G��%��"�̣�Ǫ�U����qZ|gZ�yN�n�P�̷��
}\lvC����"��ێ�f>;t��H��,7t���|o�j+�Ƥ�L�2�Ck]me"�2�A�n�-�t�ߍvL}�D�++���fM�l�&�*N�9�9ʔ�:���~�X �9�Uu]M]{w�q�u�U�Ṣ̌wJ�	�&+�՝ٗ6�5׊��m�g/]n���y�Z���$ۜ�U��SG7���R�{1��R�����Y�Y�̜��A��h�s��7�77�U�[�0��_wv�>�cbǺ��#t{�z��m=z4��z\���������(K#�*��3�!���ci-5�4����]\齂k���,�䧽B�ԳO�2c�L�)s��ne��zj����V
��*e��yJ�к��*姮�WV��׹r�m�uE�G%�Ý�L��{r45���5N����Զ�ه�e̹}fՐ�tWEL��s�]�ÑI�u�t�&���G��{�٪[;[��R]���Z{����Ɏ�1wM�ӽ�]��� G]9On�%�:9ww��NX�e�����_\�6�M��C9�ʬPP�ݺ{�AW�fqb��b�9��]�b�h'�ւu��,��K9�`�޼99L-��]������\r^LѬW^��Cd[CVl�|7�,I�[��up�2��U{9-���Kw�I^���]I��K{_h����Ѡ�CNE˧:���-h�v磏k��))Pv�x_JX�Te���i��7Az�^�H&�r�ÜrD6nҽA�"2�P�5�8�[&��1U����:�>HR϶-m}���<�n�)s��a��娰K����wE�}b%��X�ڼ���Fs�TX鹐>�;��S�rf�P�ڝ�G:�N��X��=�} =���'|�n��☫��*? ��:�-抳 ���Z��1���h �&s�mA��ct]A6��͗;��Pg�8�LN����evA���veҥv�V��K��nK&V�ի
�ǖ{����Y�4U���ǅ�<�g�O{��+jJ�mW
�d�u���0\�3-���UV,����}G;1r����Jg׮�v�3��}T�d����ܡѾ�����ػ�eV%���e�p��4�yݗ���[[�*뙼Mj�]U���G�ۻf�ʱ�e�]�j�|����F�:a�{F�:N�;b�.Ϊ�ǵ+�x�pX}�Ӫ��:ᕹ����eݝ��Vu����Uke�A��N�ܽ;7\����
p���F�K�[�2M{�u�GA�ݎ��Ieت���T�Ѫ�ݫ-�N�mY���p������A�ȑf�U��U�*�+Z�r�&�=� Y�����QnM]d_;��O�m�TTפ,y�m���^\ߪ�۸���Nm���݅J�m^nJ���]�"�.c)�-�
J�lMb�O<hu�ѕ�Jh����^f��eǽ��)�-=Wv�K����H]���׵�9Kme\��eWb�@V[5R��:�.�ZO���d�R�7p2ef	cuj�Ty�1��yb�❷���
re^Wfe32����k�U������p���s��u���T�sZ\j$�H#Ջ��̪�WW�pZ��^rঝ���}vOuf�ʵ������u�������ڮUßcȷ4�F�6.��=�	}nW
&]��7���S.��
�Y�^�e����2����u\J{�֝m��Sn�3*���ʬ��+v_f�of����R�8�T���j�{v�
��uV[�e�6����x�mڲ2CPN��̐+�ӘQϨob3:�2��u�a�E�E����U69��t	J�K�=��I-6����u��.H��o���;V<�ka�UR�uןQ���;X�ݧ-���^'�+�o.����B�-������rͽ�g�ne�۔�������Ct��{Ќ�+2��J@��"�=.dY.�ޖ���tS�{��c*�l�B�B����NS��Z��}���ߣ��udZ�0,�C��X귴��;�93N��m�7�]Q�m��s]i�ofV�u�����r=޳�����ĩ��Ih�%�46�:�Ɇﳳ�f�U�%[Wz�w)�q�988����,-}��Ǯ�;c�;��qbs�Ģ��F���=+Qyi�7��,F1�P��U�:W���뾹yXIf�}��X9��"7��L���F.1�Z�����3f�z�f�u�},��7�j����T���[�������Bε�M���a�/8d�]��,T�d�D�(���u�O.��b�%S-�[غg0����w�wU
�=YK�ݮ[xgN[��ݺ
b���n]_:]QU#�
�=��J;ᘕm���PH7��Cy򸹻��'U(O<�)�	�юim�R�3]W+H�y��]\�N�;h�n��2�fLy)�j̇%Qnt����1h��z͓�6b�.�i��懯uބVA�8�Y��|�fö��,Q;˲�{�����4��)��}���o����U\���ݫ����FQ�D�Iz�бy�T~�[�&Y�l�«-<�.UCr�j��G�ݛ3���Y��Ϯ�ˆTr��d�g���+%1��[U��%ܙ�.�b�T܏������$n�&��](�Z:k�"�s��V��nҮ��дѽ��/�]���J`(�H��kCY;��vC{G#�pP=n��ܔ�]�N�ew0-����"��(����p�$�9v������Zٙ�rmp��������°�8&E���3v_Y
ΔSfڴ7M�믗#���T�uE����[珫NR0�dX�7WUǒ�V��)qBM������F�[�)��p�1�A�b˺���|e�{*���U}��>��Җ��K��lD�4#������W�mgS�L���%,�*��(M��V�x3�L���Q�s��8�c��p��k��mάX�)�/�5Zq�Vc���SK�Б;���q^��᷺"��ܣؗr{�A-g���N�}�MT�-XŻu����{[�p�c>\�n
�����m-�e�Ԝ�g=�M�iE����X2K�X�E��ݣ���yeһ�,�{h�ϴ!l�!'.T���J�s2W�	�9��i���-7ʛ4w_gU
�;�^̣Rb�{sZ�]��B^�����������uC�p����[��2S���p�w�6���]U.��R��}M�x�T��E�,ޜW��]��YF�|Q]\K̆ء�����Ui��e��r�5�h�r]�p[X�¡x���T�S3��1Uā�����3r�`q	���30�/C.Y�����vٻRڲg]e�@��Tk4#yO��v���2J6eZ�;����v��@嬷�qޣ�w[�i����ڽ����ͪ��q�u*�*���g���i�2N[V^伨�S��s��+gGN�^q����)J�:m�v�V�#&�h��������T�Ub�[���P������*�:$^��Ws,-��κ+'V�����ol}�e��h,[�b�Ո���n񤨒��6��u��XgV���
����p��d�����bTz�h���mR�r�D�tp.Y�[�%�\�\m̲�v�^1|󯻥�WR�r'I�N�l�)m�����Q�q�Y���_,[��ޙ��Ӷ�������g:�Q�����WwL��*�u�0�d�"��u�n:���;�o����6��]�\�<P]�Ў�Z)�6��!2�P� Vp��Uga�)Z��jzt��Y��e�Fmf�4�p�X���F%��H���F>�s(�<Hy���f�۰���Ӥ
���7o�ѕ�7����⹷�3��gQ��`�g;��8#2�\$�(T���f�;���y�B�v4��!f��*�E�kI��3,�wn�T�WJ]�̭�!T4��v�H�T��y����Ɇ��21d�����ש\����k;���7�\�¨e����c��d'f޶�Mvnv����,f�>9�_�i4XO�CrG�!�yP��Β��k�s������j��k�P�S����U��OS��&���oW��5Ϩ�rȕ�(Ժ&�esFV�V(^Y�UZj[N���1�����]#��w%^8ޓ�ݖ3*g;�k)٢��-3ve]sҺmZ���(�}ǎꢷn��o�f�ŧ��Ě6��V*[Y�}�K�3���BQf�m�ɛ]|�p�A.�I���e�
`a1�����;����F$pԛ�u���x����v�˾+%3t�M�̩�Mu=+CWeSʪ�O�[�[�3��(�˽]�[*���Ÿd��v�f���`c����P�P�s������켬�V�];�V��Ԇ�n�}�ՙ2��q��L��@o���9F��H�hT�V����tFNS2�Ul}�������v��4�lܻ��;u�uan!s^[��g����:�Y�Z�c1����ugh��K3�u��w97��!��Gl��^K�i��-f�6T����m]].�N�ʻp������@=Ys��.K
녋6�S�Ezn�U��8vT��cQ_c�i�<
�ʳw��d��^�p ����
Y������u�i�ރ����2��$��	- �����ɂ"$�.���o_z����aн^�ƺ�ˊD0m�avl�{9Yl�6\%ݳB�(7�JQ�����ؚ:��� di�8���:5k��b�0fHCFWJ�M��s1�XD�6��XFSX�U����CZ[�c
*Y����1��hb�%��b��"�\S�&�p;S(�r�e�CR��3����k)`�R��5�R�\V-�Y��RZm�F\��6kjFejj�CLj�h�WA�i�Mǵ�0�����#�	W�H�eRR
p�t��هEcYcNe�i��t4tnV9c�H5΀�gR�.V]�s�D,XaZ%д�[,��WP;[Y\ڪn�T�c-�l����\4�c��͈��W�m�`Za6����Jli��n���*,X�Xd�Y���*ba4a����Ћ8N�p3MfV^�GC������Ji�,h�������`]��ަ��	L��B�.��-�ͮ��дf���u�n+���i*eaH��h�L፸�5ڵ&G����348A�בv�2���R�cv��u���Š�U�g��8�tq+��仍&ua�A�!*Fi���ڵֹ�*�(:�lB�49��im�Ss+m���-�GGC$�˳��Ե�b��5�YZP�\�]�tjdB	n�칭f���v��[��,R���і$�����X�6;�%bj�],�tF�ıG�CL���l�kl(#-n&d-���1�]�ό��Y�ј�
2�U,����
�	R�j䮻�j k-�e��)q��S�0#���a�SL�v�,���Ќ,�ڔ�6�-M��)7m�0\�[`�0�q�Xk�36�V���� ��a��t�)�.�d�+A54ٶ��M����P[Ia�h%%&����AW[u�]	��f��`�s#�R��T�UrؗJ�Վ+���%�ʹ��5H\X�fhG!�a�3��J^/W�.j���g	ve��K)CVj�5܅�����]H���3s�er@��{�{�baD@���܌`&Z��K*IL@�0l�+��b��b�,i�"��cB�mn�a�r]*f�ćd	GЬ
�]H�n��h
�+]%R&��0�0	�͈��k6�1�me��B��*�Ѣ[�a5�%�К4ߞg�.�e�Mu�iz�J	�K��E��$ιb�n$6�떜nf͍I[`�ՆՃ�7h��Ɖ�w^ѱ�+Ջ�����,�z�+\�IM�V�9�c���rj�M���R9�F"�끶�!H�#2V��C(��f�5":-&���K,Rq ���Y�l�CX27j�l닌�PT��Bc��uVnLF9HS*غ݋���+m�`��U��,kcԐ���+ �c�mX��ل�R�Ytˬ�L��7Y��R9DT҂m7������<� m���)X�&����C��nJKL%���E�\�4��'9FWmݩ�)!4�k��F�)�,X�X����b4Fi��3F�,6��m��mܶ�6ZD�E�˒4�灙X[\��Z$��W��XKa�j��9��q�����*�R2�yҎp��KLً��]!��]UR�kԹ��bⰕ���bŘq*�W(�5�ٸ�(D��ٵ�F���s�l�5�.�3���6�3.��T�Z@WChT�`�Hac��Dr�uu�f��a2lWZ��T�`JR3\*m�Sl���bk1�2��W�a�&p�lDY�@�m���,e�9�6�(�B�V[�W v��[�0]T�����P8���:lA6�����l�l�ư���Q�%./�
5��6�*n��bh������%�S6�h�i���bX�+v���]�:��a1Z(ea�ܺR������cU�
�"���{%W3T��W]�M����&Ք�@ɴE.f:�
�ZI�6f*�\��J�u������%�1���6$A%沪�"%,n�Y���lL����A!dH�9������X��i��霄-Gn����l�)XSf��D����i�a5�R�P�ld5��`���L�2:�uI)-�`cmc�Ǝ��)��A�*�t�1�#Vi�"]\�i���cI�E�m�$����u�70TNB�d�Hcd1��)k2W[�-�7
�Rc+	��c�)�eb�M��*Y�������k��U��HW2(��`��R�l�Y[l�4q��rKMs5�Ű�5-M6�����i����b��SB�!ɉl��ѵCK�����s(͑Ue$0P̴��!kn���X�ے���t��TW�C�hՃ	�����W7k(g-`������e"�H�2j�^���e��l�B�����:5�@Np[�cT-ͪ��OK�)2cA�ٖT+�9���"4q���p��`���aqhn�!3�0��5�Mt�[���P�1��ǵe��	c)�����X��v-Ŭh��W�uB�.����$ÚocI�Ҧ-�Ζ��a������XL3j,Ҭ�
��5�Z�:&��؎���d*�⚬�q�Q0�tַh��R�.���J��2��j�E�\�֔525�@9
�Q��v��b��[,��5�T�Xl�������jfg!��Y�qlmF�l�7:[�1t�҂{o���t	YCYt�C[L��f�5:�ձP�m�,fqͥ��̳%k6!�M׶��JVõ�,��Ve�����kq'�3=<\p������%�2�n��J 5���%��,�E��ژ�f�sH�J�CI����.����v�ŭl���-����:�����U��R�mF��n-W mա`#�V���ʹ�����֡��c�u��JR]��"!+S0��k�쫗g����R�.��juҲ��n��Vd�M��3W%�֚�	����&�+�Z!�I�ۋ�!��6���J����M �H �R;�iP��3i��r�+�����9�)f%����D����fmZ15q-
�Hڱ���&��&�t��iSa.Y��8%,����G���Vԙ����e��[,������.V�Á��Mm�tT.�6��Mn�5W."�����8̃��r�g�K'�e[�v��h[[����1-�ЍPk���Y��6}tZivS�+�х���q\�e
P.&$�YM.sۨ�[��f"BY��&���5"V�7M	 �m�4GF��RnEX��E�h�:+���D��B�k�l�з`��h���-�iؙ���6�T9�Η�	+i�[+���R��EZX��a��pZ&fY�Fˎֶ�&J!��X@.�p�Y16�e�W��)�fS]s��K�c�3��n��S4e�*1#-�ᎃa��ѹ4��Ʉ�%����)2]f1i�D�9�j�b���q0�[�ɣc6��m��6��i����!�XD	8�E��u���-�%)v͖��s� �WY��lNl�����@�mjL�CD�����҄ґ��Ylֱ��:օ,��bBX��QХ���]��nȦ������u�Bf�!.�����Z��W�vr�́)�è�F�6�͕P�Ԕ�Zɒ�+��cSm,͚l�*ʅ���i�ĕ"k�\DV]�K���/f���"R���Q�;�;3H�ٮ�]�-fָ����0h�6��9-m��d�̶Ü��jc0�6�\J=\І�0��%��ı{f�j�\Q�`&#2�����rQT��Yy����0�+3��&�E����%-SR3>|���M\��5`���*h!��� ��+�u��hJ�R����\�iҒ�1�$�� �4���f�˓R�l9Ki������f�a̼��\`����bc���E0�粛[�u4ٖ�044+p*H�k�B�ļ�$�A��@+k˭�܌E�Z���`/6���P�I��.���`�aM70p��o#c�c�*�ٸ%j����[P.���nڦ��6�P6� ��R �+�0�J�!� ��cl�B;
!aVl�B��:�k�IDXP�Q6�%˯j�ؚ��-6�-��-Qa��Z=M�+J�0�i��P!L��P� ��,`0����J�!,iZ��+@��ţuu@6���Jpv],��f/d�n
7����؉j��{-�D�۩����P�!)n��Ri�e�qB<V�ogK������uYhv�ilLR�b�DU�tu+Yi��uE��6s�c.�SSJ�U��l����i�œq�
�+GX���+��Zh�m�mq,̩���2
����ńҴР��²�Z�����U5��=�.P�9��鹚:n�²풶� �e]HmfP�f���P�����1�0&�a���՚]{\X�T�j���mh�9Ü�Ǜ���,1 v0��n�Kn �ƃI�7Bc^V�.koZ�kXԲ���[#��6fX\1�l��K�ר�D31�M]�[�He�[I���i���0�8J�c6�Z8m˥�[.� �5�;F�H���˂Զ
E�[�؁4G�[I�L(a�Zm�����c=T�m�2���,��F\f��3fք�Jh��AL���-�Gaو�uD�������+�(emH���b��f� )n�"/Ь[�+-v���;\q���ٗ:)ú�.-��3�nIm�Z͢F��2�-�.&�6���a�hf�4�M�"�[1�38�%t;]�o���L񥉊8�YQ�X���ϫ��/:&U�-v�3��Z���L9 ʛQ�m�r�p��r#Q��i�+���z�ք��Z)�W]-�J�*h�0Ա��V],-4	�ńH�s=c��e�����bě4�ca��8.61��źT1�p-,X��s��x�Եtq��f`�[�.k��6c4v4P�af&�	�qp�b\�JYe�h�GT�;k�2WSjlhE2��j�c-c��*.ʻYvb�X%�n�1�=<��W+\��c3���V��c�3� �IH �N�8�e܁e���BȊãkN���YVwN����� �pJN�wge�.&���䢁D�6�RPSm.H��&��g(p\wg`�Y�';X�Ίl�KlwdY�����f�:��{oq�ge�D G%�t,ܶ�9#�Gd��j��e6̵
ڲ���<��:ɵ�sh��*D��Y�oY��tte���qYf��	N�Bҷ28;:O;!;�B��{Y�����m�qprnNt�m�rwc�Β�D�K����ťb\%�v�qbr��8s�Ryd�y�qD�Â��#�C�;�ku���ݤ��rI$ޤ��I�l@�L�q�\Ut��ZI�IMa�i&��[� T�f�kh�����������gr�@e[��Ȁ�4P�-U���m5Hl��MP��jv��B��B͡MH3#�Iad�λYe4�"	�\�Ѱ��@�skFYvl��ˡ�7z�mv�:�\,��f,2J0�p3i�����M&�a������/���fnKU��օ��Ycq2eRb��T�Tq-�b�i�u�@�[�R�Gb�+�ЕQQ̪��]e�l4ƱCF\�(m���f6�X�[�M61n�9�;��PK.�9�eJp�dk���c\�YA��Ylau1J�i��h�u�m�v�)52��*�M��+�$͌�9f�&]fqv��8�!J�J�5�$o.��23](��XRh�m�" %�Y�͡���\X�݀��D(�������3KFBSJ�݅�2�S
s+�i�+Eٳi�a�i�4�)�Cie�0�Q�-��X*@��Q�=h=x�,��j���[�C�F4�����p��,�A�"e��|_x�zb�M�Z���-�ճ\���2�T���8I5���aSu�v6�"�7�f���5�J �	�g.#�Ut�ə�������0h��6�@�M	�%`n�.��Q����Im��1�oT�&Y-Z���%��6�g$�h����i%�g�1����3�&N�Ĕ�.B̶jl�m�̳'1k�.�$�6���Eюн�K:�;��K�F��M�Q�ƍhi��Uct� ��g*:���%��XKU��l�T[5�.�`�Z��1 �ѡB11�R���G]���].L���cC$V2��th�SX��8(+�ia��B:�j��[���2�.��$X2���1�#��n�2�4\M�n��f,��cq����˓`�1�J��l��t�nr�X$̮-�	[�k*���[���f�B�X�.�*�d�H��Z��Ũ����RQ:�[Kh�P
<P��-8j6R�$��@���Rb�A��6e��*�R�h5�R,#^��P#bA�cxl�F��
�`c��=yb�Il��5�ie(�0����`���4�U�qj����UDh�RZ%xH���y�_� ��c," YP��Ku�0���iJ�u�hZ	�d�)q\.슧���39 �/���-��T���o���k��0�*0#�%Wꀂ&��~_"��d�A�-������cᝆ`���}�5�)��O2!d����=CN����.��.R �,X"E����$a���˒Ծ���<6N����?����$_Y����(\��e�}�J���� ���_I���Z�aO��O#��͉q�ާ�lz+�h�7d��d�;�V�R"J�$Y=+]-��yx/��6N��71��ܺ�u�!d� d�A�XYb�ܮa��)Evi_�va�Jh�-�tH��ef��
�X.%q��Q���Ң����w���ՙ5��N,Ȣ�	
�d�����ru���2(�k�ر��-ݞ�J_%�{�:�u����)A�
�|μ5_U�3�����(��,d����_�{�m_h6��¯; �\wQ[ԲJ<7)z�F������ډ4�iJ�`��[�﬽]�W���v4̅\��u}����ERi��H%}$[�+��7��"Z�k�����34$o.�̸Wq����)2�I3{��K�����ݒ��
�+�֚̕�ԕ�I�71x���H�B���磑�޲S�٠c�+�Hӻ�)��D��9�� �>������	W�s����۠�f�'Ǿ�M4J�̜�y�{�m���#9��k�BD���օ$�!��$���.�G2�lA�KL��F���M�H�|���!�|A�#$VAJC��Z����{�!H7�?�z�&t���ʸ�+"�� A�Ib�"J�%"���7��2%ǙX!R�@�U���{�Nk�v&���2E�����Vt��Z(T�$:�A�d���í���w�/��Z\*�T�D�n��+y�OP��BU�*Q�B�Ա]�51
��<�";i\{t
f_B.�6����{��jZ7i���߯,]�Vo"i��ȽƲ%��2Ed&s�i{3�L}����y���7r�=_]�*��ȟyq���׾�6w�{Ԉ?k�,"���Yy5�Wg}ۖ���lQg������+�3���� ����H��%&�LR������*ѻ��J�+����8c,�X˝!as-���3\\�As�b���_c)��,D2W��%�r�U|ʕ��g}Ak��z��r����2�ƞ��\#ܗ�H� ��L��f�[�y��};��a9I;��f!]P���R3P?�;�@(b�hg}u���ő9 OJ@d�,"_#Dg{��ݥח�����:n�/A�Hz ��+ �)$�73�mZ�%�ϐG�}$Cg.�W�T8��V�s�<}�������*�b9�#�0����U�v\�&�E�n�,-Y{{WUM5:������U�P�gw�_��Ǌ�u�X˫��y�]Xj��|�#܂�����2R �$A"��̋3:,��8��ѬWU�{��U�R3TM��Wh"��A�X���9�p�^ɪ�U`�8P�v�fkA6��]�&��
�Z@��C-��5��mE�A��@������dH��Ȅ~�ח�"K��75x:<��?�m�u�}x�}����H�@�"B���޻��g�8xt� ����9t������O'������w����0$[����m�J;$�n�c܉c��GwsLn�_'n�	���岯	�y�©fj���X �ܾ����$�)�������L�'Xھ����K�.[�7��n��S�D�v�s���A��̚Lo.%2D "2 �����ᬼ;��s.��s���S���>=�gh̡dH��ȃ�"�Z^W�K�<1*��	�Ս�ٿC'Q��/�*��m�2��a���]ЈHI��&�j�m!���w�`��&;)YI��6�i��R,�M�QU�J�R�V4���A$Z9�5m�նh;K,-���0@cҩ�c��E�1t(,#i/%���1%]2,%����5�B��Ժ�Z)1� FfS9J����[�`�p$I�\2�b6��r���9e@���\kb��"��ZX��[`���b�f�e� ��;�`KCj�D$�qf5ȥ�9V1�����L�A������A���ٲ�[c��e���*�v0���htͅ@�RIY�h�y���H�""��&J^p�j�r���3:Г�^+sV��q�/܂� D�H��RW9�|j�^l:� �@_��uZ��]K��7u{���":P_"��b��S�Č�̌{�!wS��wrY��h*�畾l=�uW�T8���{�ί�+��KD�|dA"�B��e	�9���ߓ_S��S�gb[x�r�'��ݷ�E��4�ȔO>)1���lC���gXo��) A�X�D��'��_{h_���^�}؊��:M�_x��tA|d����G<Y�{5M�f�UFŤ��B���M1:�&�q��"6ie����!�.Q{_��Ϻ �����J�	%�r�U|�C��8��x��M�2��dxc�{E32�0"��?)Aq�i�F���K�P_�DG��˪ɠ�T�ּ�V�^0^l&�Q�ڷ��0t���;77Ρt8n��(Vl������V.�Z훧�ǁ��`��3�y����ո߼�u�'� ��,�;�@*v<+N�]�|�J��X#����I,Y%��E���w4s3eg�j����"�_�I�����H@�2Ed%}%�ڳv�9��D0����W�D'W:����s����/�'�_N:|*ݗ n�br�$V~��D�.�12
���[HN�a��ո�<�v!%|{b#�}%aD��~�.���J��WD]�UB�Q�5Uy3�X3\7�Y��J;.�WAc\%��cO=|{���},	5|D�/�����vY����fvtc����A�ú��{
�S�l�cwp��7wrS7L�VD�묅&{(��3�*�Ϻf��<��D��v4��Tԙ��5�<���nEg�ԁH�H��%W�<Vo�YH�Yy�B���ڌ`n���������/M��%{~���Ӆl˫=*lٕ�Fq���V�6����W��D����0��y�[nNg���#O;rP��K��cWwAw�Yɝ
gG�����{������D���k��캭���f�����#�d8�5�[����Ou"$A� Ȃ2UγWƾ�xpM����Uu�w�O
�� ��@�m"9b�W�H����
]�{�P���[,u�Mc�i�+
�5�W�-[Sf�wS8a6An�R�D\m�s�����_�% 9����ն�<�v!'�B�Y+Ƴ>�}�o���"I`I����ڲ^�^�����d��~Al����v^��äɫ�A�H~辒-��Z4�,�B)��!`dA%|���u���2���恵�/NS{���m"��&���}$_jO��^�4�������X?I\��y:�ߧ3݈ICǣ@l�G2w�X�J)#QZެx�WVZ��]�W)��R�h��^+W���
q�54���tS�]��g�x�vݫ��>љ�T9m�}C�3)[����� �,X"@se�2ꅇ��!�r+�Ǔ��-~&M^�����}$_i����/�?��Wv����[�2�]�-��SU�ت�c����A]�Z�4'�_d��}f�/|����2K:.3����O
�� 졛9o{�Y���c|�(w$�w$���	���{X��u�}�Tҹ��6���~��v!%� �A|d�D�zo$���B^�=(h/Ԉ2K��R i*�Zr��^'�����~&�^��c���"�2R"Jr���7�A�Ԉ�!�\g+-=�x*�������T&{���!YUO:Zgve3rU��Z��˹Ww:�es#w�_nW��7�����by�п�?NA d��D($���z��(zZbP�=sE�V�k6ݯ:���2J������߷s����J�x<��V�*�<�4����ޫ��(���^���3b�Z|'��׍v�QB�,brbS@Ь�����1����T!�T�@�Գi�����v�)HۃZҼm�-H�L�͈�
:�jK.���\Z]��M.�L�b3:<�h�������K�\
8�q4�2H��ncL�K�gFZvíe�r	#���-��ۜ�KSKZ ��X\�4NE���aW;1���ep�Tj�X:����~+���l8��(gKv�P�2�]X:WJ��a��j	]��H��cv��~�A�`I���-~�]��';կ<:M�}�<�W��A^R� ��+ �%"$_�� �x���]����R��/�q���{�<M�g�'�H��X�$����X����vi���%������\�H������Fm��k������z4� ����%�"J����f*E��{u#ޯ��}�]���;��xt�Z�n%��9���ڬ�n��P�"S.���YD2Rh"���t�/+���;��\칾��Y���K�]�w*U������w��dl*VAHU�B����˹�BAƱsZ�͔\�KW5`YS,�\ʿ��<���������<��V�O2Ey�}F�	�J�|��Ȏ4��Q��d�,$�������6�Wmy�e��3��4~+2��懨fwC���u�Ȣ�V�e�`���:��^��dfYT%�x;�̆m���Ң�U�_]��o���Ak����syަ�údk�|vR���D2E���6z�,��D8�'�@I_IS��Q1d�zn���^�oI�sy벳T�=�K��(w
K�%��=��h�T� ��="�A��Q-�b���'�s|��7�>3.$O7�ܺ�]T^��� ��M@�d��I,Y8_Z��[���h+�{���syަ�údk�|vR#�}$Z&J�L��&>��,݈�"�SM`Q�3�Bf�u��b00Lhu����]ݫ��p�>@�g4� ���|��Uá�3>�c�^b�b����庻9u+����� ��+��%">�Za{�l�sڬ�g�y����97��=؆�	���4*��/R�k0hͻGr@���2K��BD3��hx3YX��V���g۵Q��u#��ڪx٭�^����]���zeT6�7��K�YT/z�d�Q��Ejս��u��Jl�ա�lv�C��mO��P* �'gdOm����&*A�75�Jk�s�㕊��3UV0�����/#���I���u���@e�*����r��x�{�,��6�g&M_l����N���0�ӥ�3jR���H�H�U��jsvĥ�S̪�j���p�lč�7�-�Hji����]+R�wݺ�v�u�ژr�]�-�k��!�tR'(�Nf+�KF�:��x�s�+��ܬ]��+vUկ��պ}׵Zk�\����7J�}E�Sp��+�{�^i�S�"r�D�z^b�[Э=����uU�(2�^�;+��#]\���g�'b(f��c�A�E�7���������v����,�݋��v�{����
�9����W7��:U�5n��\�W]'��|i�]�K���hw6U^H�K�$̧�^>��:jV�nuy\���:Z��3�b��%��������B�>>Z���8���������wr�T�ì�r�QcP����r�oj��<S]t5��5�J.܈�	��?3n���EbKVv�|�}�Tk�8���жOij��8����At��Y��OA\�t�k��ʛ�:��-tY������e��Yq(�^�m�-]�]V0���V�{�T[dt�[ΗfwL��ز��.̴�)qS�bJCp�}{tt����ͤ�����e�M�> ��1��7u�N��ʩ�]�-�۰��I�;-*n�����㜯�v�b�N�A������8�f�s�9�Y�s���[4�D�v�D��p�;��8۲Yg]�m��v�t��t�ˁ I�e�h^ۉ�8RR��Y��NM��C�m�̰"՗-7�֎=�^��
H��j�r�&V�f@��η���$� �Oz��})�Ҳm`=��/7n�t�_.��}�{׉�{n�%�D�Nq��8�d���N&�9�Z��(t!^�yw�۴A$���%!"QpfJD�>�`!��t� �y��[v�q8�[���)�w(6�Qŵ�8�(W۲y���Nr�pバ������kc��H�!Ӝ�q.t)yn������������7�;�F���A�H�����P>s͍��&uy��5�� �%��3�7{"�U9�/��>t�#[�{L�����=������ȧfJMd�A��^y_��+F��i|3�e6�G�~��݈l�@�z4u��_)%�yN�}~R>�vj���ٿ�Ȫ�Wt#cv�F�e��m�c55ʅʻi��0 �ޣ�e A��bȑ|�����yfk��Sy��25�2ڻ7�ɍU��A�A��P_"�4(}>��!ܤD�*GC�
��|gvN���F����i��X�D�vק��~�y�����	}H�"��d�3ʩ�푎ʯVb�<���C轚�|f\T�|	����fEMf@��c�Ya���L̕*�	.��^9�׭<��"� ������|�y�+�+��"l��R���j+����Oi�/��wS��%Hgf�f�ڜ�v�˶�S̫M����2^+��`�Oo�����?���~��@����2/���쿯FXe����B�X�C��q�EL�'P?�D�]��W��޻���z�|��>X����M{V�^F�"�S�Zl��f�W6�J6$١B�Vm�{�k�����+?IK��8��λ���W���$��ܒ^d)��)�r�i�Č�ƫ�3�����(}cH����/���]x��^��úd���� ��}$L��UOC#u�_9C���ADJDI]�X�	Yә~�>�۵�$]eL�����>�D�,	7��D�*MQ/L�\�6w�ӽ�'���y���t��8��}]؆���4,Mv�3��'��V�c�� A�g�Y �2R%���>ǽ�׋�Ǻg�1����^9�ۍ[��w"����_I�����{��ֿ_me*�����Q�W�^�N���׮c0�Z�޿h�,n�7kK�sمio��.ܡu(fU�q�=�m������u˱��lHGi��Z�l%u�v�RR!�b$�0�F�sb�b�X�ۘ�7�5ff� �������չ)(���Lk�k.�f8K�hV�i�f[*M`�Z.�m���)P�rkt�f��w�z�����81(.�:�Jb.�s���W��d�Ly��6���7X�	z������	B��O�L[��K��r(:1�T���?k��jQ��t�X�� �Ƥ�Cj*���k��]QT�ͪ���j�e����辒��$�T���UL>3��gŊ��3D�3Vծ�[�� ��G�|�_I�A��#g�L�|�_۳4h:�Y�:�����^op���^�Q>0����3���3ʨ�d�n�n�V�Je��]��w'�R,�~[�<=]W�iq�����ƭ��;�xK��=�E�%"$Hi��.� �k�+D,z�����Ҽ+fs�}����i��z�z�v\�dv��#܂H�L��2 �2Eh�?=U�����g��n�����x�轛Ț}�c��� �%�/���y#���s��a�W�2(��B��h�*f:d� ZnL���
ͪUt\�Gz!dH��JOq��׹���<�E-�����\���W�% D�� 	~~�E���[3��{��=3(��O�j�nv*�8��Yշ(>y�ƺѷ�3T��	�m$�uXqcdd���h��м��EQ��q� @V��%��V�<�����\|Go��+ �=�H�_��L���M���;���AجO�H�"�H����/�̺��myMwΝw�yN�74���ICfJ��j��]ʓ/�xMC���;�ő"_�A}$�<���Ɠ�w"���D��C�`G����}&|�2D/�����K*mkZ���/w���PW�l}�|`��D��}CH�� f�:�f�F�+ u-�b�q j��ɵ�b�k[a]�f�V�P,�!�J�]��A�@�E��i)}�zKɅ�٧����b���ߌ}[z|.�=�dA=H�"� �2R#}-�zw��orǻ�������N��1�\��~���^����]FH�G�:r�kԈ��_o���"�J�2K�5���<<q�c�k�,����x��o���X��!i�q�N,#�۹/P�����'��0�|h��se��;�ѵ5���8-&>缒���� ����z󧑉�Nߐ?m"r�����Yl���*�VAz�-�`�������i��Ϧs�����в=�R����v}�i{_ �X�D���KK�]�fvJ���\A9=ǖ=�\��sÝȼA/�z ��Y(׷2�jf[	�@�TM����PH��,���]�nf���n)�N%eeMM.c���y���ND�𸩧{O3�4��̥H�d;S�󧔤��Y�x�G;�v-���,�r_FH��%"4;ۭ�����4,��cZA�������~�s��xؚ���T�Eg{��̹F-���ߖ4�����2KM�$C|)���묮���K�qn�Ǯ�����Ԉ=FH��d�D�
�o�����!d� �3ԁIc�t\�Iy'��yӄ� ���<Oi�j�=H������j��\/ա��˒owr��ʽ�˻�҉]|��qc�V��{�Pɫ�T'��m��V{1l58��7-����>�����|{� d��?)��"fT���Ì i�?W-���Iݯ�zP}����/���Ic:���T�V7�Z�>a��yHZƔ���:0�47;-b�.���1j�Y��e
6��{�e"r�����D�wu'�n6m�w�||"��	ߺ'�_wb�ފ��H�����w��^�}�E����d;P+�=��8N��H���X�D��X-����Y��^��i�Čj�U��XܕYj����x^V���]'�>������4,�A+�"D�!,�Lw�����W�@Nо2 ����a��͹���//��^{.i���m�7�@�cV�R"D�D,��N<Φek��Mb[*�+��C��3q�yӄ�|�=���!`����v�L�_z�`#N��S��f���+Υ�7r�Ӯ�;6���5J���.��Ӕw�)��}�}mގ5�#|���<�䄁?n��StTLӁ1l�,UM��3..h���l�m��Z����5bB]r�
����	���m�l �G!@���e,o&�95�kc���3�����u�dk��	]�Y��,���Z����B�ƥ�^H��1f��d`6�(֓]Ybl���̥P�/�U�R�L���k,ՎJ��X���CM�ʩp�ٗF�8����~�� 6�NLZ�b�.�6�ev�e-��;R�Y��Dt��c�B�����A:� ���2D��gW'��I^ާ�A��*���M﹠�r��%�"D )������`V���m��K�=�/����=�u�f�5FMi�;;MI�d��]fo����_<�	��/��d����G\��T��Աz�t��ҭ<��w� �� �,XI_ $A"��\��^���W�� ���<��%!��\�zW��\�w�z-M����_oVq׻j�ő"@�%/�Ib�"Jk]�؈7�
�͞�Ku���S�/�� ���tA"�� �[��3��.j{'����-!���te3JZ�s��-����jm�l��j���P��F>��Rc2�]�]�U�,�j|m���,5E���S>���[yU��,��|�A$V~��!���N�e��ɝR�d]�$|{�҈��nih�r����ްb����h�I����W^z����)w5�7'��[+�w]��I	sz|�~�Lc͉^��K�ɏoi���ƨ�{�&��2W�c��;w�7b�#5|��/�� $�����0]կ��t�ke9��}+��x"���J@"Ae��So*f�A���@�"��˪�u�y�[Yӄ�	��T�?͞[)p�=�|~qd����_!"��A�f�UԷҌs�>pOv5܆����)y�K��Le��u�=��9N�s7��_Nv4v��e�`k-Z�%A���,\jCq��A�4�fOS��̽~x6}��7Y�A|dA}'������NxN����*���S��ئ5�$�m�1����	�!`�A�^C�]�p�w[���q4ׯ)W7��v��v�|`���i� $���Z��]� =V> �\���/��}`*�F�/�ת�b��s���J��N�F�����9WSrQ����j�5:�*d��2��7y&�uU�W��h��|�����{oi�@���Nn\T�h"�y��<̥C.�I��a铱Q�Vd���S.䐹����o6jO	ˢ� �ԁi8�[��sPV�"d�YH�2U���^��X��NUu�y�}V�t��T�yؖ3=tP2�BS.��>r�|������u�VP՛FѽSWCi��;*a�,��-��g#P-
mu���ޞ�~|9�1��<l�d�9�<琞pOgj�����^7ATG��QX�r ��/�?	%�"J�ƯfV��
��"Ԛ�� E37����Z�r�x��}Hz ��$'y��t��Gʉf�T��rJ5w"2R �$��������6�����罧k����&���4^EI�Ȕ�̜�ŧ�͕H�T�N����@{��2W1��E{x������TM'�q/�A��]���凯՟��^�k2���9��7��%.�꾝�KV���z��Y�/�eّrp�ݸ����>%��2'v�]�8�p��>>}���)�i���!`%���,��E}$������Z�9H�A/���d��2V�s��5��,��*UWF���k
d�x*��B�dl,�y������u��gr����M�qSN�(�;O��J�C	d>>�ŝ8N�^9W�h}[�E�B�� �2/��A�_Y`͞��z��T8�j�4��/I��-!u����sr�4�A+�_��/o�1���~���$�$��!k�j;�k��][�{{m�=�rqxA}HD�H��%}&3sj �;�n����I#ۉ��܆:�|}����Q4�w��5�<G�p���2EL��2 �� X'+3���s��x�罸:r�s�l����B�?����!@eR����JK��?7�\�D�70>�P�b�.��)\0Z�xbO��,�W4�C�����U8.W�V�k7j�h?`��)l����A֞APf7zqv�N9�ƙ+�:��wmj��n�F5�B���5��/9�wU��м��F.�e֍�}y+5��5o��sW^M�B���5�	�6�Ec�1���MA�y��dG���W�쬡��2ㆥ���3�Ic%�5*n؆XT{D�\�:�g�J�O2�^�oO�o1�wY��]�$$���k���.�v��iS��n�.���r䯢�aE�.�����d�&��L�v���oOy��Pݲ��N�ݙ�����!v�V�X��[�F��ǚ�[ų-[�w�a�9Ա��[�i�*U[9oW��|���F���b���ý��+w�O\Cj
�Ytct�R�;+V�ݫ�6�k�ޖoY�N<��=�sCv��;��J�r�.��X�=��SgL�M5o�V�l&f�Kܵ4/��}|H�j���b�OO��+)b�ۖ�R��s^L�8pʡ�!�
�����J:wp�������U��ݘ0b���z4E��<�9���n���W+eZŉ�|�!�Ц�q�������yXx�s%��D�΢oU��.�n��9d�qu�)+:���=���3���wwz�����<����^n����я�/��c��κ�ݴI&���x����2>I��y��k�p��S^u�A�:�fQǕ]vj��Gl�ź�U�Y7��{ȼ)�\}��z����i�lm8p�8�9'JK�G�c�8rp�$��j���mےs��ԗ$<�7-�S�JBq9I8H'r ��t�+���)3u�m`!N�N �9$␝y��\�p���������9�k"q��v ����pBYY�;�E8�l��ܝ{YI���[Y�"��;��Nھy ��9 �����@q6���D��{{؅
H� ��砄�;�h�����y� ��kI ^�qNvVN8��HEչ�[o���>v3�PfS0�K�%.>`���:*��� ���9��H!y������w���z��{ʻ���ث-����kT���m�f�Sg(�쮋9��-3��C�n%��T5����F��.-�' ��i�5[��e@�k��v,f�s0��L�?��x��,5��v�[ER�0KHCn+��M`Z�.���n���j��B��w6�Kt�)q)]S!3����ܚ��f-�V�uZ�Y��#]�3� �\-��eJ�Y�.%�lb��4v!
��m��e%��ɬea�gE+��X�D��m��䔕�ve��񠦐ѽ�z�B4�.S3n͗J�i���#�T01j�Auʨ�\�C#ô\�c��nIcFRX4ĥйf����Vmp���,i�s��h�6�M](޽�`��Mff��f�����v���]m�R!Qؚ��K2V�e��͸�\�s\�keR&r(�[�Y`�X!H�QMc�����'�DVX6�1�7@��nm5��"���EZ�n)f�v�N�2����k``�\J�Q���0)ZB�ؔ��XYBR�їd�g�����GZb\ۢc3�t�ٶ[��aaP�$z�& ���VPH�^�����6�5Ԍ����Wf�$S3[a0ы:W����]���"��x��ݳ�n���P����)�Gq.Me�b�����&��Y�n"f�ʔ#���-#�7�L�3���LMO�����XBX��`�kC)N�i�Ca���7&��:��I�v:Za�qHD���ĩUGr�(��:�ce�1v��麋����4�<���kjb8���MH���al���fmIy�vitPn�1P�VZ=�xꁬ��;k30����Џ�ҵ�dn1ka�6�k�{XYo���F╪#,���6���(彛kL�p�kVf�R�J��KGV0ɋml+5� 1iK�m�WE�b楌��R3Q����+c��/�lK��:�n�	�.6�Fm����H��Vҡ���;@�0� e�lP������n,2]�:�h�V\
٥��"�G.�w����wI;�.���P�h������e���m*�����P�M��.t���{[���U�
��N[
-y���)l���W�b�v�����haXYu�i
3��se`��64&�f\�k�^65�
��r���&5n��n-�]K6�2�A��ibM�f��8�1
uX�H;f�w:R)vZL����=d�t,�%դ��kb �2�)�4�<�����V/)*�m؛6�XBf��+0��]�H��ԅ�P�h�n����@�߬X"J�J'N�ON������*���Z�ʰA�# $���@�"9=z�=s���}�����O/iRa�非�x��	���@�9�D�I��@�#$���T<�R��]ܮ��	��,����_�F-!u��٪'ǹqSO�JD$�dH��K��_\;_9�`�y/��)=;�=;3��S�g'+�{~Y�Ō��_R��(#$@\� d����z����ر�{܂�]�h��FQ6{��^RY��y�K��g������_Wd)��^�a-	[�� ָٚԔ�h%H�Z��i�Q�JG�������\B�(����y��,l�7�#������!����o-x����օ���>� AJ)�r�]Ħs{�#;S���U����6{�\/|�2�^5�����3�E�乥���T9�s�RSj�T�p�΄q�]8��Gۙ/;�T7�K|��Cn���L��y� AQ�|3ޒU�^d��דm�?q��^����tA$N0ru.k;,a�H���B� �")D��B�z�sXײ �W���7����F<�)��C.��ܒ��ha���(��3���ӽ���y��ll����Ǥ���{5D����������8���g��L��#N�%��街q��W�;��]"���l���z�Vh𗓚�����2E~2W�&���;��ѲZ¼h�s1I4+�K6�](�\5�â�۱f�F�Һ�0��ˑ�����ܒ��)��)i"�����т�TG~{�O��GJ.�������/�)s}�w��~j���A'�:X��>ߕ�	e_`��'��Y����6�f;�B��3vdc͉5wt}�˹:��ܙy�V�9�s7�ӣ�K�8�2Τ5q疘�CM�Ϳwa#GՊ�]��Y�Ӎ������f\����(��[�j%�Q���oc����\Ɲ�o{�om�O����|�/��~ �)|D�����5���!�@Ƃ=) A�X�w\�
�'Ƣ{�`��D�=�ג���a����4��|D�-�ȷHCh"�%���w��c���Wx`�����Ut�}�g�orJfd+��1�wI��o}O���UT�;C+�e�"��J`�\ܳ$ՄЦ��WU��mZ�~@�)��	+��D#��U�u���/���C�Q�P���%\A�[A�VAJ@�(#$@Nj�<5��|};(^I�}�>z�U�°ꪲO�]<��a�6{�&��K3���V}���@�j�/��� d��2V�^N��zs���nL�T�����@�o /�d���X��P�#=+�qT ��)W̊q�E^�%�{]����d�A���G��!���uݧfV����P��ѷ�YCI�v�ȵ�̾
�f_n:�X�s�$���^�F#��h&��%��.�۾��כ�{��u��X�}������>wf��!]�U��Qw*�>��6q���ag�b�;��v�,�Q�7ӄ��H��X�$K�(xըwn�i����
� k�K��l.ъ��mvf��Y�֍UH��Сe�E"��1h �:D�}$ZA��K�p�=����O�h����w\�:]�oݱ���nI)�ăwtpu�¯e	��O�5�y7"�/@�׼�o��'S���Ԉ?tA$Awqi1��zk�,݂^^HUܫ��Ʈ��G'S������I3�g�,:�=�cL̥Mfw��FH��h��깾��� �����s;�y�o���>_f�������V��=��V/�:!`��%}$@Iv����?z}�y��ܓ�ڛ9�2u8����"�2Eg�(�bOY��H��|��g��^��Ɩ�<�p����R��'{�(�b��G��cĺ%�pd�v�ꥣ�T�/�4rX#�(��=\��gj��62��	!$mˉ$�r4�3T�aك�*�jc$Ή�Ҋ�Lm,3��Q[�k��S\)m��mZ�2�cj5�՘�e��J�0Z�aJVe�]���e��3m�l�d���hih,vH蕅�+4ٻh����l-Ж�V��˵��khZjJ�:�B�i�f�Ό�j�m��l"��ke���/i�4�+��n�٦����*�ڨ��4�M7ϟK��)�����ź�Eh�Uf9f�*)���W6Cm��	h˪��T�O
����rJc=�H��A��VUFHyj-т�T_Q��;[��S�ɶn��u1�����$�����r��;��z���X����M3;��{7=���\���@���A���)��1l���a�~�kx�.]�#�@�)|AK��_H�N��:�pݓS=�N���K������~2R"D��yY���*���=�r�$�\0�:��O���F��v$��Ȣ1�g6��e�/ЧvIww4���L�A"T�n�ڡ��/p�o�/���a�{8U���vJ2�IN�$�rX���{A�X�,�wv-|��B��6*A��λ�X�Ս���t��ڴU��R�pAg����v4ՙJ��d�k2)�%�x=-_�9:� #t7{ݳ_�]R���}�#$V �_I��� �+2���e�lZE�H��yv��:$Qow2������z�:��)񷷵�Z�a[��L���;qPq�j�#�:���훮���>H@%[�瞉����� �˙�?��F���������̟z��F�̋H �Ԉ2 ��X �*�ؼ^�3����m����.y}�@N��J@�$�$�lUg����v�J�A��������Ȧ^�%�x;�W��0��~;��T��a����j��)>i�Ƴ$B�E��(&��I����>�)w�[�U]��7��/4���ă��`"_>�)p�[������Y�Yh�
��8`��o2�S�<k
-L��Ԏ�YAXUj�ט z��?P@��2R�9�e�S����������	����yA�ZԈ?	%�&�~2R���wm�y��C������
0	-}���j3���o�bhΩǙϴ��:��������K�1��3�B�H���H$�y�`��ݤkj�`*�WhO<u
�o.������{LVu�U�ɐ���0��V�����.΂Nq9�s5w��vuv�c`�V�s�S}���$��g����y����^�H��i="�%���+#޽7Kצh���Sy�ޜ����1Ü�U���Ua��^����MT��yݥI�cO�5"�}%|���cYh�C2��P��Dl�KFl�Xy��uo/@;���H��	����-N���^�ӥZ,We-5(l�����ev��Wd�8���v�5�Dp>�T;4 N�@X�2R"H���՗].�{���'x �9�iv�GՍւ�nő"_""�~��?>���ܻ3�� nE`�񒗘�<��ߋ����-��=�B� ��#%s��>���"z���j+�"H�"D��nѝ��{3f���l���xt�O�� �Wˢ�H��d��$-�n�w��{�� ���=�ƚ��T�(;>&J���t`����@f�W���7�ț��{�U�{����Ҵo�T�o�ݦ6��붋���h�����r#G�]�,g��Y�r�_��}U��zτ$�\���2��)�� d�	+H����$^���?�}��:�i���-�{ׇ��/bl��M>ay��Y�Hn_{��|.�ޭ��UG@f`����%����;,l\�ū���ڒ��0l3U�u�@������"D���{�����sä�|�F���nw�N�y.�����w+ �%"$_ ~2D,����;�:_Z��w8��\�(;>&J���O��M��ȩ5��xokWd���
��و/��+ �JD�A$V&J�k�\q���h�3 kv�/Q�ɢߗݾB� ���+2KMN�oW��ٴ�w�1�d�ذC�|dB9��h�qf�>'S��;)���E��m���r������nee3F}����^�C'�d�/�����}�W�H�er{�;ج��+1m�V�cnj�;�7+gU�!��S^�Ͼ��,�T'X8rV�sŤ�I�˶)ڻ�^�wv�L�n�W~   W���������ցDX�[���"�B:;mc�Q��Y��6H�cQ�ڜ�`�(�@�\JQ����R��z�f������HL����Mei�Ȑ��36)DvK���6нn9�b�bSB֢e�:W��Z2��it��`H���F1��4%0V�!5[a��̻h*84�h5��bYZV:���(��K�C[M�.�B`�fQØ�|�����GK*�y��t���jĄڎ	b�n���s�\�u%���b��=?�Yo���|��Y"�AJ\��
�i~�#ݓC�3��8{_��n�A���_)%���)��5��;�i����wrLf�Y�=G��|�A ����H�{Yʭ6�L�Mq�v5���f�I��O%|����V:}��vyd��Fwq5ӄ� Nz��"J�J�|����w����+�<��d��ub��n���=�4<�@�{|��y�e��o7Ŭѿ�|��ző"�d�� �,X"On<ts��{��1ܝ�1�9n����r�� A�FH�@2T���ʮ֯������e�%3�*�Ch�eW9�X��;i���-F�U�������A�#%#$����q^��q5�O��,|�܉���m���	�,�|�ޭG�s��ٯ���e���q����85<���c�V�h���n�}*��kL�87��}r��!/sw�Jߠ�����c���e�r����$l8N+Ǎ��k�tm�o�͐N��Lڣ��D��^�Σ�=���_6���n�V�晚
�&��Sm|�z���Ù��k�~����c�xm��қk���7^���v��viu)�x��ǲL���_	(7A�[�yns�g�=�n��ݣ�+�֚k5�f0�#\TmF]�U�]�F�m? �}�����8�aػW�љ<����������鶅�W�ݵoe#O����љ��&�7�������^L�����_o7a��o��{����n���F�xY��Q.�WNJ[%�WE^�:ݮˮ�Z^^Dw.�u�_T�*�卼ń�z�\[�7(�9O#��h���afxj����>AY��ƫ�*�s:��Qv6a\�n�bҫ/Mf}f��]��kov�9sF5�ǐ毶ԕ�ɠ��O�$�g�����§_1#ΫWO{&f�ι�otm�ꗺ��Πk���;�,���˵uُ�o*f����h���5�q�.�iS�4L����h��j,:�۬#�=����۞���S�ztfg�R�A�ʡv���6�!+4XD�J�r4/&���U�Ե��'1m�"��-�ٙ��=�3����9}�9v�vWGKoc��Y�tx�����,��GF�{��UEQ�]�N!j����l��ʨ�;q_|��;L�^D��7�.���ή*�5����N�Ry��>����ڪR1�����ᦇi��0�JGwL�w����AnV��V��XE"3n��鶁p�0n��tZ��ca#�h��V�)0���9h���\vtN���GVky	���R��a�ޮ�ş��n�ۭ�&bu�9t$���Jμ
��8�X��T+��R�%ul�N������T�wh̠���ޭ���nf3Pg��Y�I�����	YC3�fe҈�m�2�c�Gb�=Xܵ��������jO:�X�ȼ��n�CK��Qsm�[��v3�f���ڪG��cɕ���ݛ�#v,��#t������ڐd�{��B�t��dա�Uڷ�^�P�_�4��=�r�66&��-EU����}�u���9�tNDr������b��L�d◵��s-G3qJ)9�ċ��ݎ��d(��Z��ǝ����$�E���S��9 ٬VhN.����׵�R�K�H�u����1e�����=�mƢ��{�n�8	ٳm؎D��O�;�¥��"��1�����"�=�N�6ܹ��-�����sM������9��0��}-�b7��}�{�h�o���{��XjB��B�J��Y`����{V�;gd�[���{���O��Y����͒�,i����{�E����k	�<�˲w�����k^��8�Xm��[l���}��y��"���)�[,��J@��[��S-�����瑜p@
R[	Z��'��'N��<�g�!o���3���RSu�m��^ro���3;&����8��Ƴ��
�O�z�=�5�%c7P�n��ۏ˫V]�]�܇6�v_gh���]��ko~��XG]z�ҥ�D�V~WB�Aq��l\�*�a
jt�CC@lu��:�������W�y��7B7���x��^��.i��W���7�~�W�Sm7_6=��Cݭ���Cr6�kK�Ʋ_���L�� �A�35e���ou3�2]�����@6��Kι�iŴ#|�`ח�ۇ3�ƫ�~��lM�m���9�n7V������$���|��ww3ý���FR��A�y�<w������t����{�aD�sQ��,vd�/&���.�a����Hg
�
2�Z�"�K�}��ο_Pq7A���M�g��d�g��U����.�T��Q��}�@oSm ��z��9K^VYҴRFʱa+DRM
�k�nX�4S)�-�\�WB���p�M��w������a��p��1����5]�����]��7`�����o>�5G۽+tzr�7ks����G^_�v��te�����3�l�R�t�2g=(l��A�������t��b[���g9G;i���oP����e{I��^ok���<'eg����L�jTN����]� awk���6��nު�ht�
���������{�K���~A���m�Og޻��<�Ҭ�W���W����g���t#e�c�[J�v�[��}�݉魵W��3^�H��j=�n�>��}�A+W����+����$���S������T��k���aλ3&�F-5�b�`J��G�b(h�c�&��A�s�Gi��Jsn�9�4)�G'"���R�cB:ST)��j+JK��Z�u�"f�̣�e��3U(���m��bM���X1`B�X m�+�.�`�X�cXcF\LS,�f��Թ�î��e��ܶ�Z�EeL`Ѕ[B]5��fk��3��~������8�0��,�c�[��2�	W;h˛.5��Yf+��[���|�����t���CV�<���X�ۘ9ǳ��' �|� �R��D�m,a�|�O	�}��/;�j�=��;b�X�uλ̯��+��6��o˽�+P��^��k�Cg��_9M�m��Y*{�����n�n8������gmt�{_mI8e{xnm��}�A����t�M:�u�/r�~ٜ���vggh���]1��(֛n�w��78���t�W+��a�)d\,��렔�M�f���,X2�CUWdU���Y�h�6�����ðM����C�������]F<� � �M���������y~��<s�>Ҳ�k��+E}�oc�Y�r��\���W}C�O����p����Ë��n�'>b�r={*M����|  �?����"W�����p,� c�m���/j���|�H���������J�gq:s�o�����\�q+�o�ݔ;Zn�n�}�i^t�/f�c=݀7Z�0K���3O'};W�ƯUl7���{{�NA���=m�C�����T�'%~���p+���c���m�s���"<lжM��	�0�����khX�D+Z%\.X�E�����3p�m{+x	��6�msú�hW��t͗�fp{%O���鶛��*���o��oވ{�7�Q�2z�[�����x}%7�Q����w���;���|�o>l*��Cw�w��R\T]B�L3+NF�gP��>�&��7�1��
a��o~c3��2��wN¬a��;]۾���a�7�Tsi�~���	z���5�Y{�YU̗߾�C�ot��|��N��m�h}�:�`W��t��ݔ+��9�=�L���:��6�����测�4��������s�S}��C�)�6�%CY|�o�����Y�t�Dآ�:�u5[tCp��,Ըb ��jV�J����J��|��4��=~�+��,�u��{��f��UU຦��u�tk�a��{=�}�5����˅vl��/ãn�L� �ֽt������C�鶛���U���d��^@�z�c�~�5�x=��%�6��A8�vM�M����\�+��}=�Y��}���ۜ�P��O =R��l��=~R{���nT����쮽�Lu]̻������w5��gt��st�g_����_���݆�x��R/���:>�{���y��.̓ݕ3|:��M�����׏;	󡶍Q5f�vjZR�4�5��l�ƓJu�4�i�J�Cf3Ay��_P����od��e�6���i�s�`O������|�A���/Ij��W���w�/����F� H_��Ȫ>�;s�N�� 9�!�4!��n�wr���C��#�݀�B���T4!��p���\���o?fi\=�u;ȯ�~̓�*~ ��І�m�)hC�e!��%�4]�����
hEsnlO���9���"F�}(J�p���^?��q����o�c� / >hK3$�{ݧ���o}�E4*�F�40�ܠ)�]����\hC��"�+�A�}݇]�ʯ`!��� I��בTn�����u�����І0/��)�nAЮ�@��]������LMmq����7�U���ܮ�2@�������aק��֯)��$����ϫ:�et��9/}�g��Nֱo� >����虍�G`X!� Vj���8X�A�e�0уv&]n�f$؆a�`iP��ͣl�e�@K�I�ą������B�!662⅖�)�m��%�E[+4���bmWYa����1S�M�D3�R�LLk6&��0�CA�&�F��P�hXgF3$�j+%dF,툳CXb�茩��l%bf�@�e/k�Ԇ`f��X̺�9�/��??��v��ft˘���h ��c4юR5猣K�̯[��7M�D�q����~4%�l���3�(D�
���w(
����l���,��ؿ�=���wh��>گO{h*`�>�i�vH�!��� ��.�B��0`]��B69̩����iq]�����B��@��6� $=��bcc�_����g� /!�`fd����P�hWpp�IꚎۏ!g=(
`��H�z� ]ܡ`���CMp�}��g�	{$�O9�=�n�箝s>@srC�І0/��-g�A�����1�� %4���F����BrDdƄ1����n��5�5�=�z/�v�0h=�����G��?�ըG��n��̀4��SB����HЮ�@���z���}x�LB��"*s���w��������
���B$hWp��`�/����1[��<�ض��Մn��_Vp���5�%��V�Ʀ3S[��#ѕ�ąqLj��{��ƃ�@)��"�
�H�h��	�n^MQ��z��3�7$>hD������'0��4#�6����������0.D�~9�Be���Ӯh��Xܗ��kwuu��	������7K��Ÿ�X�Fg��	��9E��*b�]q�U*�2�y�97C�o�>| ���|?�h\��% ��͔��̍�6kvk�{�=���hC�@��B)����U�I�u�CM� K@{=!HhCL�]�"Z��4
�8�����a+{�4ݩ!�ν���>��E��B���CB��"Z�)���� ��1�Tr:s���W8���^hC>�RC�	KE� M�켚��go�r��3�7$>hJ�RЍ�ҫ2�^� 	ܐ5�W����pІ��T�˹B%�]��	�.r��y��F�5�5�.��=����(hC7�H�uƋ� ��.�2��ݿ����GF��ank3P�"\���UGD�r#�hCq*�
�5O�+$0�v�hC2�-
��
hCaw	>�ͩ��q���o��<�y�hC���g�liX��Mf�P�hW�-l.�P�.�%�h.� g9K�r�"u��$`��=�(�f^MQ��o�v��3�7$>CB�R��� ]܁5<�4�Ȏ����i�v��	�� �hCWr�J�)�awr����٘�U�b
{���g �;��ǂY�����syb�ۨkc��]l�+��]ǞG��-���Ѻ��Ǘig�G{}�� �*�y͚ܚ�������1%�w�HE0Wp�Fmp-wrЊ�>���y���h�!X4!��@ߤ��1�� '뼟�cxr��{~��W��@��(4=�}�y蝍��#�6 �4!�/�(��hCh.��wwHE0Wp��}��s+�`��	+��d��w���b�� 9�!�І\!KBːD�B����p��[���=1��=c��<�_�{�g,-v�c�X-,F0i3m���\unf��(J�AhhWI��$�~��K@�􂦄3�J-
� ��]ܠ(��r7�٬�����q W�>��>sɬ�Ӵvy��)�
���]��wrЕ�d��s9��Ǽq�#�B����@w뼝���g>��gy_ / >���AP4!��B$hWp�������#�������h6��Bwt�.�S1�� 9�k~�f=y��ۓTn9��_�+�����|09p�#BːD��wrl.�-w#B������o�}rɡ}(D��	�w(
��r7�٬پ�/츿�+�1%� �hD{�Z��;����묛g)X��8ON�5��Yt.@�Gs�k�rsrV��Yj�5 ��tX�&rU�Sz��ZЗ�}���
��B����Bhl Jh����1�wR��܂$hWw F��θdr�b;�ơa3	����f7�u�����|�����/$ˁw q4!���@gw�O܌�US����s��#-m��r]i*�t��c��r�i\���d7u��hC� �hG���0Wp�X!�p~�̚�q�}��=\�@srC�G>~���{�r{`r`@b�d->������l��TЈ����/K���[�ph\�)�a~�@U�_Ӽ��fϻ~���� ��|1%� ��o���`����v�p�����F�g��`{a
F�;�JhWw RhCL.��3���,����ɘ�r�9߯L�W����/$B˔"Z�!)]ܠ)�]�KB;����m�|�'y��P�nB	`�p7��ɪ3M���G��������B��G�/�?V��o祥���/� y�Wp���.�$hC`]ܠ
.���]��s��}e�²�G>��w�٬�Wo��\_��p�>[�"�+�A#6�� �#O#~��B�}��}2�.\�sv��e�2��tR��w]]%����WU�n��s*��p�\UO�7TK2�M�A]�"��7w9�0v36�����*��Wѻ9{�Le�_5���Y�o+��N1���z����+evڙ�Z�b\,Jɫ*��]͘�:�9���B���͹j��wU�o8�c*�Q[���3�Wn�5k8&Գ����Lq�&2n�)�,��̦k
Y36�ݫ�����USw0��׻�p���W��ˎ�MR9U���V�5v�3�����ߘ�8���P��3`��9��tx>�M�=�V[��괤n���e��w!�U�*V'5�w���:�d�ٴVg��r�b���d��,LHu3�n�7y��'r\Y�Ȋ�����;2l���p�Y�s K3��!���^]ԫ{�j0f�=�Xf9k�+;�0�Us�%H{T\t^���O+]���v:�iՈ�e��u��w��Ob�̾�A�]�}yMwbB��k����i�	^sGn��a	���|�^\�݆mɁ,��f> ��.ʝ����h��K��t�s-4�Y�"�8;�弪����k�/�<�v�[S��{X�\� �Y��c6fQ����S嗻�n�h�h̡�n�+{��á]�Ӳ��8�h>l�̣����V�v���P��_�;z�u
��x�,4��q�x��.�F
���n*�/��#����7���W���oQ=G{u���[�vN�ٷS_.5�̩x���L4,�u���簼�2�Q9;��<��c��X:-�,x^�z3�}��_ƕh]�.=��&H������Ge�Dr\[f�߇m��n��8\m�Z{^��o��<��5��v�m� ��[k26��}�^�͵��������ݳcSn�2�-�f|�Mm�vj ���f�[v����-�0V�������$SG���6�;+;56�;n�̯��%������%����Э�'�<�$ͤٝ�i�Y#��[������o1�2��X��؏}ﾾVq^Q�6��`O-N��h��;0!kY�Pga�׭��ٳr����Y���
����Ҷ�Z�XW�w Rà�Vu�FB��v���{d�+,l��i�E�n̰S���e�g��ۇ��e��ٙ��Y�m�D��ݚP�m/���M�m�Z�q�ns��k�ױ��ץ�`�9,�.��`�=Y@�8�d�KDmen���kS37}��4	��c66���[i�%u��J���X�Ût�;Z���SY�[c[)���Į9�ֹ��[k\�s�H�Jie�tl�#��lL���v��\�/�nn�P(��Lp=�٦��S,[u��X�h��Ǝm+����4�i�-�&͗�5n�Vқ]��Z.,�h�?���OX']�ٰ�i����;dlBmV;qln�UQJ)e�6,5iW�n�d�W�X��8�a���"�.�v��x���ʺ�5]nؘ�r�{Jf�5Cm�D�3f�F(�GA�������af��,ƶ.kU��h¥TL�����3T4
���k�[uنKj[�$:���9��C����L#��� ��L�[b<�:�����j�F�[B���LF�Enł*4�7E��N
&���ْ�.v(�&���ixcpd1`WZ�Z��`92l-�[���"��Ͷ� ��MH�P�1��a���ٳZ�V�Cjƻ$�P��5�ؖ^���%-�6����lx�[HSR�ת�M��3��i�1r����LTT�IT��,YR�&�Q��ʬ�q68��[mz��KfH*H�M���KkM���X�X@���-�.K{F�]���l��a�b��U��L���Z\�نs��oR�ڰ��Y�x�؄��	��Z<E���������[���˗GL��3�X]Kj��Mw]VgA��m�,0��2�]�kl�-���l�[�`�;-vIU�V�aL�=��-a��IE�-�Q���B]7\ V;6�u���Dm�#I�"����ױ�.ՐMqNf#fA�^-���nVS��4n��n�IB�6���&a	��b��-`ܵњiͥ"�k-SVh�aF
�-\ٍ�/S���	+�r��P��k1-[�A٘v�Z���S*��6�V<��Ǭ�>srU�X+�m��-�4�"�vԎ��{)]G��tG�h���r�W��qfCA��2�.��gh9��X��n��7��;ń�l���[
�2%��0룭6pT�A��M�e��<���Y,�F�눌v���AM��^�2��f.���UJ�ԛk�tp���ꙴ*&@�A"�ví����fSl�xXm���h$��N���ɠȨAr�.Xl�J3
B�wn�*K�\P@��n��S6��5A���Xa�c��b7V�2����,��������������5�.f]�2�a����Ќ��`+�C`��]Г�����І09��-��"SB����p��˼��cyʌ�~ߌ�W���[=��I��ș�ot
���ۄ"F�� KBawr���.�%����R4"�܉��9���L�LrK6�d M�32j��k�����>@srP\!|������z#29��b�P�����H4%�r
��]�-
� �І��� G�5*�Wէ�Vv���gE< ���}��Sw%�E� K@]܅4"��a;�|*�hC�-
�% ]�s��L�s����d��y�4!�2�APЈ�f�����������\�"F�~�%�a�d����h.����@p���}Q:Wr�+� 绾ٚ~�+s�G���7$>hK�R4!����:4!�.���|s��;��G����43��6�FܣkCE5�^xs+-2���),��U�q��@cB��@�"� �І���E�n��{5�uw��n��v.�\_���|��;��P�^�	w��:Е�!KB7OG���}�������wb�6�fyy���כ��u���u�vUb�N�ms��*o&���������oh���ꮩU���>���^~?wd
hCa�Ѐ�r�ꉝ�9��o�Ok���B`m䂡���"F�w o��٧�I�=�Gs�(
`�Z�����h��B)����!�]�+����������+/����/s�| �r�B�RІ��Ю�@�І���p�d=68�{���������г�Z����n��{5yuw�gn�@;��Y�
PЇ�ؾ���mӟj������ ��.�B��6�!HІr�.�@�;���>���B-�n{���g�s����|�{_ / >Mco$4!��-
� ��a$_ ��i9z��>m]ݫ�
��/�Mf4���Kv�EJi���	v�V��a��!̈́
��ˀRІn�!0Wp�S1�� &���3N�6��\?w����4"����y~����]�5�H"F��P�&p��4�����ASB.�,�G���`��a {6P_ٻ;���{j���]_���ml��=�RL� ���f�z6�Ah�F��d�4!��!HЇw �hWw SBaw
�;q��,�=e]Γ���P�H��1��7hduU��eo��r�L5z8�G;�v&�����{��r(oU��ۻc�ɶ�:m��>�Jڤ�fV=�x��� / ?��Mwr .�	q������#���FS#���A�`�!��H��`�4]�߾�ɚw������>@wrC�62��|dW�t�ȏ���D��d�M�a-w#B�� ]�ѡ]��uwTg'�߷���������ս�V{yw�g�����bK6KB�)�
�K1�� '��k����4���{�o����tS���fڋ"\��+�X����:`Ťa�]�n�30م?Β{ߺO�@�}�!H4!�d#B����]�K��f"w��W����U|����hD.������9��y���/���P��#B���I�]�HІ4p
F�o{w9W}o�B-� �hh̀	/ۙ�4��k��Gy� ;�!�І07�(T��d)�fd�]�}����7P�9������%4!��$4#3%�hY��c����t�)�W��ouc{2N�s�
�d>bK6HЇ���S����� ��fTlz�M��W7f��{9��N���2���ò��s�G���������ӽ�ÙӖ^+5����/���;�{�Y�XNh�-�}����n�]�u:��R�\�������X�iR�"�⳷��%�7:JE�R������·�~_	"J�I$�eV�@�}�.�?����nu�����$�I4'�}��F�=�5kHs2��`�9����@��lX� km�nm�-�U`]m����!%}$A�wWv�z��t�3�u9��ב~�Bw��P�!$�ʇjb�����76,3{��~���Y�}��l@I$�y�;l��Hn��T�IWO	O���j�c���(�u���N�`�!%��_��]'��H�ԛ���=�Ӳ,���e�U��ص�<�E��$C�"���t~̮h՚�d��k�Ε�+ن�9��v[��v�$RT��l�Ö<6�-��8u�[�`S5+�lX�|����X�ň���v}�_`�H��(\}l�#�[�#�!�[�+�o0�Λ�Kz}��݃G�o�������N{ߓ��5�����(�mZ�⋴��`�.rPv�r�M��7j��G	�$�ih��Ƹ��%�3���J��k1�	k�H. .nY��Q3arIq5�����Q��w8&���z�kLB��Vf�r�\s,�u4�
/��0��v�G�k6.L[ f$Ҋ�,� ��FКͬ��Ye(ٹ��Ō0�S*25�t�U���Ľ��6qb���O�Z��kƬaW6�L�ƃ
KYY���f�D�k]h�f�܂�%�{���}�I�	2I&+��nt%�_D+�0YY��j�n���z!$�>H�>�5��;w���x���/�f���>�C��$�n*.�}��������}T���y�OL�5�X`�]�n7�e�|ք�%I�D{���Ư:���=1�BJ�$��N�~��]g_O}���g�];3����d_I_I�E%��z���Sk���o�Wv�zg��vE��:��ɢL�~�>t���*�F�A!e`�e���;F�i��c������kC$�4�WDt$�<���'�D$����/f]9�{m��;up׳��� ��3�"�/����0j�C��|��gn�ڕ���w��k�R|����5Kv�՝~�޾��I�Sb��I�y��O�S��:.��/�.ʳn���)��]��?u[�LX?wU���]g_O\k���ӈ�̭�Lnߦ��H�����׻)}T��鸼��wwNɗ��uϔ�	(I�>ٔ��g��,����E���>ٗS��a�=�К3����~}4vW��9�J�) �K6e��T��̳��~��ξ�Lk��$�$��܁���&�p��ȋ5VUY5L��6,�jZ��]���n^s��Ճ�a),���LV�}����RT�|�ݸ�ޙ�fxq�oR~�vǷ���%	"M�b��[��{�_?O
����w=�a�=�ք�!p�M�Q���<I'z��I�tk�W^mm�2�ʻ^j�_`�oi	MB��B�g'g�������¹�Sxl61�Ga�J;V!�R�Ђ�8�B���a�u���|���f���{�`ξ����uI�D$����-̽=�*�[����ޠ$�wJ鸵����س�����U�a�/��/��/��$�u����^���^��}�{�{m�MrM�J�I��9i�k%ժ�
ɥb�S6�jPզ5�S�1Lh-)�^� �!b���93��ߟk�=耒!��ܓ0g�����r��O�S��{�5�^W��C�"���8,�#����V���}=�3| {'�o0�|��ǻ�{��0�G��� ���$[<�]*���/tU��]/7���s�MhI�P�/��yd��p뼡����_IC�f��Kۜ �]=�Ǜ^�M^M�����ԟ3v�՗öIx�~�Y>�u�}Z^�n���U�G�7���4x`���ٻ�y���z$�[o��� �����l��]ܫ����y߯���5z��̜[��}=�4�y3<'P��I4H����{�"�tj�F�г�j�i1���a��Җ��,4�G]�C3�l���h�LH�����2�w=�����d=:}�gd�}$R#���[���*��/��1�&`�wR^�����&4u$�S�����)�D��\�$_I@I4޳l��ʏ��?n-{��;��[��u}ϗ�E��$E!J���ovwוBH�O/b�K��_�m��5�]ƃ��mX��s�$_IBH��Th��۴r�}�e�R�C�o�*!�����:���%��sK&���+-W��u͝�n�V�tޗ�K��-.]�[8��4�3�w�$�oEpgk+`��c��K(��r�����Ų�j���W��g�y[�y�G"��e��״�̹�e[k������0���m�chs�[j��ҡ�"lй�51�M?���2�lj̷��^ݚm���dy�ʛ:�R��9�����YXX31c�\X�ړK�,��%�p�m�L�a4pV ��Oai[�ut��r�ڢ1�	���l�՘�6��4"�uf�v�ZXJ+��C:9K��HE5�e֓o�/���ݫ�`b��t�R�Mr4�r��r@�F�#k����(!VU�t�����@��D��a麟ƞ������Xk�����ɂH��!M�i���t�a9��C�~�^ŗ.���{m�	��Py�*���.�}@ID$6��zOm�[ޙr��N�.y����G���/��b�zЛ}���t�$Cd�{����gN�.��N��ˢW?hA�tC��&IW�F�M+9�
��\��x��,����g����Z�)(I-�i邵hUFq`-��s26U��ZCh˛�ͫ,���V�B�sJ�Ҫ*����e|�!$RP�;��7=�!�����W���3���fE�ܑw~J��iŻq.{I��7��������^��
�5�ZP���|���T�z��us�#&{g�OVw_d�K8�y�u��}������v�F����y}�����wI���u��B��������S���ܾ�w��I0I6�xō�ݣ�>]�/U�پ�'��#�JI�I�g�W��Q��[�d��ņ{���p�rr�_�=��ܮ��k��Koe]»�A$BON�|/{�D��͝���پ�t}Ϧ^����$_I]�����b�*�����0��+��0�0���&��K��[ˑ�*� 6c�7�����Ӗw����Vh��g����{Q�s�q�^c~�\��+W�������	$�i߈k��z��;���f��,u�����5˧��Wú�����f:�8Gz=��I&|$����a�<�Ή�s�jyUY���%�۽���B��|��lTSlmc�۬�r��2̽AQ�W��AY]�*�L��˃�>i	o���̆�}��k0ӳC� t�;�Է}u����`��X�}cu�����N�6��Zr��{3w�_u��lgV	�ܬo�^d��y=��k.��6O��Ө�Om}����۪�dU9Qv�K�33�^��7��ծ�ee�Ya���n[�w:����7�]�Z�uϻ�dH�.nI��1L�������������I[���×��5+<�+1Jq*�h�#�5=��+7;j�V7���vmd�g�����g���<���;شG]ǱYǸj�抾9��(f�M͋��s,>��j�e־�f:�(���Ü���X�nR�-�1e�wsH��T��[׌f巪uӜ6gmw]�V�{��/l�r#r�l7�m��̱�i��l.wk8��9�5A�P�eD����=9oM�/�:|�8Jo�۴Sv�W;V��uYF�tų94u�Y�{NO=��3�STX�uj�2�Yf���^3_�-�8��K�6�bN��3>��a?G0����V���D��]�YvH�i��ƶ���o�S���&��͓Uef^k��1o�����<3z��6�ΡQ1^�A�k]�\%P�W�K8����/��UBؽ3�Y�mW^J̫}�Ae�)���n���$3/�1axc�r�k�ښ!y�,���y`�X������К�����UY*�2��Oo%��}�F�K�,ju�f���ξ��]��m��4����ֹ�]��=�Ȗ�R��Ƙ�j#c�{[�e�3���q����މ��{^�SZcvs��;ݷ7n��[C&��M�M�h������m���w��d���(۲�0keo�i�{|����6�ktM7q��v%�Z���N2��mN��{4�wm�#��^��=gd�Ɩ�׵��/2����vZٵ����p��m����ٳ΀��-�L�DG}�^:�Iȳ3�w޽Ƞ�n�!y�NG�w6ŷ��n�̶���:;ν�n49��q�g�����ͱm7K[�^�YfY�gKk[v�������'8�ntu�V36Ҷ֓{�y5-mf�m��q�fc5���٭�����y��h��l�ѱv�_k�k��l7ZY�t�&�l�^�{�72�޽�6IE��ךr�N�ͻ�i��^��-m[5`�g-kI���6��A�h�t]�{��b6β�浶�l�l4�H�)e��vv�2lM�" �c��J9�ˌ��w=����L����9�&�*H�(�K%:}Q��_s�}$A������fG��{m�5�^u�gܼ�o.���)"���/����OW���7T�۸��qW��O}7P�"J'���-�Պ��]l��%������J��Gt��6`�6��\d6&Yz�W`��B5��m|#�%}$['N��{�~��;�m������nkQ���oD>���}$C�i�hh�cӮ�}=���}�>~9ג߼���k@G�X��f9WY�Ƅ���I�}&[��[�'�����p+��J����7W��$�	"�J �wS��rZ�Cg����өv��{ٜ�t���w!1w[�����`$X[���啚��ydमz���;zN~7cپ�s����a�⛐�<�}�+M#��R���,-�W����{�}��I�}$���Z�W"��%��0]�μ���]��k�l�����2�v��i�����e����6dv#z�K�32l=JUU���}vA�j��ᮇ��I�IC6D\�s�S�t����եm�_(����y��RE��E%$_g�
�g�����=�;W����x�^�R/'31�w��=������I�I)ߴgt��d7��l]��^z�y��s���8��I�H��:b;S�k�o���?h��l�97'��~}F��{纆ח|�Nw]���ֹ&��I���B��2IԻo}ޗ��wt����8���&^Ր*B�^]��tx_��u��UBW{��T������ֻ�F��qq�}6����3��gh�pvQ<xn,UW��O��]���ͯ�|��'�*^hM�&��7K��I����r�K�d�r.Y��q4�f�\b�fYk�.�1SsrCL�襡� 1,%�),�"���Ķ	,�\�.��e��s\�:�irh��`hGX[q*�qRV6.r:\f�ԻC4��4uq�/fR�����1*!f��lh72���#L�t��2�6(	&�P�µ5�Mt��ni���L������!�p�b�mBݖkr1��ћB��)FU]s,X&�
�6��~o�d�$~��엎߹Ŷ糩��G��s�JE$RW�4ur�xث���ެ�rnN
�y���麀�$��|6߰{ֲW��RD$�$�����^���'�C��ov�|^ e{xE���řՙ�jZ�y�����R��0�fd�G��o�}�{�������un���e��T�M��I��D$���-.��T<߂�7'O=:�ut��C��$�	 򾗏~��|qe0����Rk��+�����%��P�]���UV��ڃ�RPM���ȷҺgI���r��*��/s��%	"HDj�Jx���`������*�J��%��ɇm[A"�ʬ��Z�n_
��]��WΜ,�:-vi�j�WW�q��<|��.���e}�>߱�To2�u��Z�sÛC�䐛��`�d�3���>�_I$�Q��^z�Ϛ���AT������n��$_I$��S;q�}�s���Y��f�'���s�0�½���\[	�b��٫���H�� $�"�����wC��v)��;e��ͯ���*H;�q������o� {���Y�M.M5�\�cA�m.�su+,e�
jgE��t37h�Iw�޾O���)"��͐'%��T���������=Y�3~��ו����%���M�~��nZG��'=�c'���k�/
�V��}$/R5Z��z�v(�	(I��k�#�!����6����[��ڝú�8���j��Z�ٖ�lq�\������1_r�VuNju���i%�}!��dn��� 8O���z���{�~�@G�>�!$G��6��{^�����6@�w�ªM����u.�[Fm���6rP�u�;��WU�F��Z���{ޱb7;Գעw�s���^!��c@EI�9L:�1���{����R��S������+Mt��ltn��R�{#�mML��Òm��E&D�QT6�g|R��J;�$�`RǨ�U��}u����Ξ���G���{f$��ݺT�I�'���C���z��lj[��8�?{կg�W{���dPȵ'�qSXuF�1�����ԕߢl�p��X;�I~�w2�e�������u��^��y�9\a�������J��q|�_zs7g=�)VwQ���P�(����'x A����Y�)��v����Cn
�"3��U�ۄ��e.x�W�:�rú��B��/hv�h�λ,5�K�G�D���j6��PeG�莮�\�����w>���h�y�4c̉cY�E��CMt��"ASaט�o)tew��W{����3i7�qWxN<�c��l�C���`�[�]a]VM��6���k(W+Y�#q+\j:����D�#O'�^_�9HͥM���r��r���g�yҾ�<{���S7�i��sM���h
�&����꘻z}u}��!ݒ�MRǨտ|������xXlO�s%&��J��{�+qu���^{���V���'�"���\��Uٛ��ֆ�b{��<*���
�3ì�OX?�M<' �i�)W�ck=�3ݷ��i�e*Ma'�s2�r�Vᵟfd���'җ�{}��������_���I��4*�SMQ0'��X�V��1÷,x��=�.�I��׻�w�I�2WЊ�	8���Z�R�Ѥys"��#Y0U��u��|�w���ݪ��spKת�S�tu��Sk+z���?��C�q��t�����ӿ a�GG������3���R��-1j6������)�F]20���32��L��gV�Q�K���]kHP�`����ܝcԲ�e��&^WT�GM�"��gG3��-�cD&U�۪�3H\�6��04�Y���)R��Y�����@�,�2�n�HSKmZvX�EsX�W5�{b&��w!6�C[��{��U�L�n�K�mjQ�t]�o�����	�����U�:P�ī�ٽ�YaX�l�	�q���܅�!�sr���|~���Y�*`J|�������Rg�Y�.��^�fg�N�GM�/b�͔�Rh"���������u�����M{{ɡJ�n�_:�6��,���Mi��ؓO�R�>���ܿ�r}{��vq�2�>0ة�D��;��^
}�.�^8=xr������;�>=2W|Ф�ܜ|�0%q���gy�N����{�(�Mby�=��R�ox�I�r��{�B�"��Kpu�yR~	�X���4���h
T��ZIM����)&j!=�;�^��s�,ˇ���os���&��L;}Y'k�'�ܫ3{�r���٥ajX� �P�R9�pi�J2�F[�����ff��<���W4ȕsH�`JMs6gw]|����z�xN�����ߢ`���V�q�
T����^k��?]7VSv=<������yc̧]�s���}�{�蓑b��c)R4������,��i�Z�G
XCW�-��t�4��?�|zǜV �Ծ�8)S���o�d�:�chX �<�3�ov���&Emx����ZM���Q{^z��wD~w���O]�Ϥ]��Aҗkp�I�)4�v4�����}�WwbZ��D�6r��K6�u�����{�ü���4_:��v������R�0%&�Ě`W �&�}�>�ϫ��a����R�{�TS���B�{�M��T�K6(���}J��ro��#���ם.�3V�e�MtAf{V�m�B!1jW�"e�CUV�+w�@�]���2���.wOx��~��q���n/ C���x^^��jT�Mx�T��M6�T�Rk�#=nO/�,��Y�*�u����}�a���%.4��R��������j�	�*O�"A�4�p�vyP�ZFz�Hxd�=u�Sw"#i�oc�:�������m�q�[I���ZVV]Ugp���(/Ot�Q_W{!̢~^3o�]�Te���R�l�-Ne�(WO��T�|͊q�)4����gq�u����`��biٔ��;�"�n�J}�^N|���|})|C:<�����X�<��I��4r�`EM4�(�����d�Z�̑��{���=u��_���{���%4��R��qN4���۳���~~��?|*�Y�v���n�҆K��9hf],&Ø��A��#�A�����q����y���+���ò�s��-��K-��6�����^觳�ص����'�L
T������ݎ��廂��[�N0)R7\�O�&�}���_�SM'���[�*`Gf�z�iغ�Ͼ�Ri<͊�A���H
L����q�_ڳ�Y�G7�Nx��C�tVA�ӬX���' �L	\ja������O5���`��b��+{��ƥ<����>e��w�I@�ܸ�v��������E!-`[-�XU�EǢ�vq¶Q]C[iݏs����3��:��O��{}�����n�ڔ-\�w�⚽) �9L	M3
T�L��Wt*��,yaﻼV��u����<@s���Y�����P������P��!U�1b˝��Gh�#-��1�\��%t��SIb�X:Wj�n���W/�Uƚ�(��h
U��r���
�{���	�-���e��;ߢ�'���⦂N4*L	\i��=�g�욻�	��'UJy�?_oZe��f�3�&�ꉁ;�w�:�e�>������y(�a)4�����*�qV��y	��N�`Y�=�����[^4�;|[�p	�a�ƀ�R����뛽���ZxE����KHmM������s����@�3$�~���,ܜ�b�0%&���Sw���r��7���w�����hWOX&l��Lآ`NR���y}�}��6�<U]��z,v��n^�\B��
��`2˷�<�`�$n���9N��ﲃ���n��E���w�����nrp�ukh�,��׮�rK��{rS�W]��+��r���R�9t�����e�Eu�
��6�g�ϯ�n	Ɵ��ݹ�Ø�מh6��|򘠕>���ƽ��8kُ{Y�gl��s�Ao�t��3��f���:V*�VEvT[�:�)kW�(�k��Kl�V_0E���n:<�����&ժ��|B�J	�˹��y�Ԧ�;���n%��C,�n٤>"ů�T��3��M]�-���y��,���.�:��i��3�,�S:G��ڹu^dHӓa��	ȁV#�߫��'�r��`�g+�4h��]Y����u��s���u�f��r���9�]����c�w6�f��:l����I�M�����v�#����^*�Eh7�=B��i�,�Ss2�aG����2�9|{/u��;�v��7�II��5�ﺌ�o{�D.f�)*�z/-�g��҅9���L�g���x�Q�� ��j"w1N6k�w�L��:
挏�]�˥bl�gj�IR�h�4j��[F�/x�]�6R�}�1�(���޻�on�[#�[#�
j�0V�wX�"�M���z�{{h��Ru��*����t���]Rl��ibX_^u�0��6�̽�o���Ykf�ͽ�yyN9�s[ê��*����j#�����:�ݪ\��y�w.����{�Or�{:�7��-ԥ��8]gKw���f��%�b� �/�������͵��j)Yu%Q�o^e�ȇQ.�y���N�Z�G>��&l�>w���ћG`6m�m�lŦ־���ڙYgm�{{�[6��e^jRR�m*�^�@�Y2_}�l۫����3m,�bVKn�[���vѾ_{�}h��h3������l��gjp�}���囋}�G��ov�2�y�[A�nv���-�^y��k:��on��M��kXC��μ콛��cve�fa��;D���C�ۛYmڶ�`���Xܦ��ěv��-cN�9�"�E����.y��֖dIl�l¼������gZg��h�l�lq������gd�3��Cfsk5�knN��3Zm�����q���C�m)�Z͚-�6h��4�ۢ�ܳ�,1��fO�W��[��������kk����u�toj{tX�~hv�דF���g1�A�\F�������vZ4�q[l�Jܙ��������3ME��Ķ�,��0��CZ�fy�؆��{V���l".�;R0U6TM-\�u&[k���V����F`�픍�u:��V�ia	G�F���m���B��Ś�X�1j��
�Ф-F6^7,���̈́��3�ZKibf�1�ht�ҋ�����b��U�q����h�̲۱
���ˍA�ԅbҨ��78!Y��.��̙MM,s��t�mlfi@���ƕ�V
���A�p��kf����`�1��CP�3��-ݝ�t*٩[+��Re�(�f6���݅ЎҖ�@��*��h,��3v㋢�v �����m�Eq&��� �i�����疓m.���lF��Kk)Ha � 15���k-�n̵�����ct%��5"1�v)ui�D�Yx��u�B&��ŮG"�©��{$`V6l�\�5�F�%�L�Tm��ǹ��{&+z�
M��@!n�T+�a/iR,yı����%\��u�	�hil�U�f��nfSd��;2��3K��28�QM�.tZ��k�s�s��Ae	k��+�l6�
�xM�ж�hX�a�qR�T�͙��m6�.mX��	�P+l
��Y�f6��\س,n�Tu�34��ka�%�nR�6+ �U��б
�CQe.3+���m�E�)�Y��#X�v�iJPT��ݜY{i��х����!K6m�2ڼJ��5ky�l	�,Ҕ�aT0�bv԰-L ��[]i�[�f얓*��*]����B%Ԕ7i��8	X�h0��ej5�Q��Rl�vmU�i��[M0 ���-�.�ZM��S$�ԥuPٙ���8�M5�8�VڶU)���ٙs�nv�W�]2��ke�-םnu$#
���P�P���� :�����ћ7J��R8{XZal�5��k� N�A��f33Zlkb��ۉ��U�A!�{V�W9��XFb�G#j�*��.#m�h��v.+Ya-��5Ҳ��\��J��3f��b`���[�\������[m���ZX����]��hhY�Ph���a���Ŋ�X��	sm
莫fP�F˖�:�v�X*�rKF����
�XX�J�Xֶ�dFk)v+��hL��!D�ؙ�R�1��5�8&)�c.��2�Բ�Ԏ���%M6��B�j�2A�*�����F:�i�\�Y�K��@�M��E �*-���@�8�
md�>O~�������_�m*I��q�
T����|���ݯ���\���OC�x�w��-f�ñ�)W ����Z��ש}�_'�d���\�Sj�Ti����^,:�铔�)Q�fJ�G��{5/���`��X ��=�b��������M�����Ϊ�߽����υq36�O=�#z����`R��EȺC�}����P���d�4����5��*3suϔ�{���|z�W/��/zYMw>���f�i�=�����EI�� �O�=]�*J�x�\ۗ�&�ʍ7���ņ����\i�R�����o�qvm1.�Q��Wv.����;��۵wI)P�F��P2�#&��l�նX������4��W ������xW�}�|+������/m���DCMi9{��&��0%q�KG(Uk��}NR=v��fU�Y���0�ub��B[T��qY�����hḲ�%��ֿ�u��Gje��&���(,-���:�2���rʪu���=���"�77\�?��l�Pz�Nx�R��NB�=ܯO��ҵyL���W��/q<͊�|����߉��i���Z�����9�w�����*h"�*`Ji��:����w���ە�ݜ�����xW�~�>���R ��/�"HC]U�_Ty�hCo�� �6�&�(��O�R��W����\闶/�/}>�[��\�?���/�=tW��nv4�
T���QuD0*�%xZ����6f��s,MBa�Fb��h�3b�Al���:c[���J율����Ri�Ri��SL
T��ڛ_#ۻ��.��]�ʺ��w�[.}Ư�5���@R�0%q���<��VWU}������w+�����;g�^���\Lͤ�w�*�L��%_|�u��k7w��U*�ZH�0��B����c�+���#�B�AP�wBVk��~6��JZO�5���W�=��/)XW��[�����a�y.G���i�Gʄ�y��nf6�i>(-�e`�;�%�����Mi��ؚ{�*L	�fB�Δ^o9���Ȩ�{u��)���f�P�Ho{�W���໼Vo昬�s\̎^^O�5��3�����i�bi�\�S�����w��'����&?l˳yd��X ��,{�F�4����J��:��7�]�v�j�LZ�3Z�!�ҩ9u����֤1
�)�Y���u�J�T�)4�iJ�A�@R�77\�O���m�=�k���fow��+��}��=�SM�bM\����ț^�hR�,�%�B�Ed����n�J�������gV�铕�I[.O���>����܊��Ĥ�y��i�
T��|a��U���mv��׉�_�a_xϯ���I��&��D���MI��W��Ri����5�'�#77\��H��۰��W��4��/���O����yf�V;f����濶��F�몈�m��i�dWX0��j�c��U��̣n�B��,���j��9��r����QRf�mw`�5m���f���-~���O7�ԟRM4N3�n�L�~��^�A���QW��������f����M4�)SA�@R'{�߱?>��~�K�ai��2�X�1FYp�M�����n��i�U"M�Wd$hD�y�m"$���O�;�0�7�e���v��z#ۛ묪����zr�M4*h"�W�{�3�ܿd�bk�'��T���W���j���W�����M;ҕ0'�Vt���.�_v&�ԩ6J�E8���<��3�{wfw����n��w�ƨ����Ф��S�
T���噷\�-�V{+/}>�`�����<N��fk�ӡ���{�Y��@~����씚|��U��EL	I�*Ms3.��f����6�+=�������aw�^��os���JT��i�m?a�|+����f��(�3m#[����"���;����'ɝyE����K+/��{-V�WC3i���"޳��f��*�A�L%�.�Fq*u����15���\JMM.e	�a,ń ��fg;5t�[�J�*Z\$ڪH둎��f���Te-�F����MDu]�Y`��6�tn��H�aA�������4�*[��F��BP9F�j����0Z��QR-FSuىH���c.z�̹[(5e���K���4��0�&��1K4�,z�4*ZB��ia����Pf�c�����cV0jh�qU
L�/9,�#GD.�W@�6l��m�RMΫ�����Y�^`J�MKY��W���N���_ygӏ�ߵ�/ S�m*\kvrp��+�6���ީ>��{_X3�{Z�'���Ǜ��&`[ݣ���v������f�Uٴ�&�'�E�5��D�vp��y ���JC+k��_s�~9yh�z���7�{5��;i攩�9L;�,ǾR�zٔ'[�ƞ\QᲓL
T���f_W������z���W����=�]]��}��׿/&����\Zi��i�
U�a'6�]^ܞ�7���vf�S����]�/���;.*M�r��k ��|�Ok�	Q�uWf�*�3&�/YX\��UˈD�ȓ`v�����!������Y.�Whҕ4N0)Pnn������swۋ����d37�ʼmV�A���s	\i��U�"�5U������{:<i {��������Țs/w����m�zA����8�sz{G��}�=^���{wՋ|���
Y9��했����"_���ohݥKza�w�`]��Pi����QC3"5���c��Õ�)�|�i��NJ����}�g�fI+w�U|��/�K�4v���vdT�6(��ƚ�4/^���}}��G��!��W�J�F��
T������z���7}���Ҿ�<��_�	nK�N,~۔�og�&�*�|{|��i�����Q�+���#�s�>���_ț����)Rh'���Z�2y�����MQJ�]��TB��ȫTH�z����.İ��T��G�B��X��� ~}��ϛ�N_vr���ow���4v�c��{=U=����X�͊$�'+�RA�����S�!��7��>��/������W�}���oos�4�JT��!�<��� ���������W/s����rl��'}�k�O�,V8.ϙz��]�o�0b&gW�m�n*���0��X�磗ůb�Y5yvew&<=�g٧&�^;y�����[���7q|j���MnRh"�iJ�R|��~�y��=�%Ղ�X�畂	���:�{���Ϯ��ۋ]�4d��ǞNh������Ҧ�rp	I�"������Q���W�}��� 7�Wԡ��{Vu�����Ɵ3JT��M�o*������ŷ����̎ ���.-�bؓQ�����.�����i�[�p�����ɻϾ2o�X��������mY�=�__{��}�}���W|˺U��D��0&�7��K"�}1�W+4u:;f�3�� Τ��ԓOs��{�M�'cB����+�i�ޘ=]׍�f�ł<��NW �\h;Ȁ�.��0��y���߫�Sם����g�7����;O��*`HfGP�̥J#n�%I���T�c쨝��M4sL6?�{o�,3=�_��Ed.<�e��zƚ[���p8���7�9gǜ݌Z�}���,��3�yr���p�F�
f,��
f��sɑV��b�2���}X�/�������L;O�
U�������C��f�{��v�}u�~h��'��"��F�)�d�Y�Gw#����tG�TR�t�(�cTjd�vy�d���:܍ݲCF���*M�[���|"oK��Mf��zp����{�}J�������+��n�<��Z�D������i�x�6K.�ԇy3m��_�Rw�����*OM6}(�o��hf{�_���f�IL��{�]<�N�ۢ����M��4���	O�޽��w�)gv��g�V�9��q�GS�~;� �b�	M4*�A^�����]�'45�y �\�{�O�7}=�9�����})��˃�U���|���� �&���L"�0"�|�^�����t5yز�X��}����7���䤚in�4q�
[�mL~�����*ˬ4G�����^Y�)�E�l�8��6�{�?TǝEm�?a���R�aއ���03�N^�����U��rS���<k:{�#*�÷�77AX"���M��M��7vu��Z��T�J���hm��I�e�+��Պ�օ�+jsS6������)��B1��i��p&�ʱ^�&�u����IF��u\鴦��^2���ٙ��׳[�fmβ:�F��I��\��]��0	�b�k�H��kmlgD�sMJ�h��o�v����7/���6����+r�CM���I��.p!6�����{;
��mF8�sf[DU�j��.����������3g �O�;�;�^헎���S@���vd�F����hx����ݞM&�%8��v����;.����jMnw�sM�I������j��Y�D�"�&��G}�u���'��7��{���y�.�[Y��4�{m��o7��{�G�g{���EM>n�zq�J����J�{�k{�M5�R����L;��L�zYK����꡾�IC+����ͮ����U�E0"�Wk�R��W]<���r���[������Y�O/��}9��v4�
T�r�	������ױ��$�<�#v����L��䲘)��5)�{e#��XMr���7GkJ�&�U��w�*M<آ`J�L
V��{*�7��}�#�3���/���Yu	�T�i�̥\k	8���I�+�6�!��
��^����Y=��&�4M��wj/6�Fii՛�y��Ad����2B�-����f�Ӣ���n�4�sG�w+�ԇqW��\��_�jO�4ѳ�K���|W���E*UwJ�E�D�II���dw%�w X��P_��ٵ��Ņ9��6�g���os���R�H;�&��[^&{�oV�=���pݞi�J���{*�7��g�Glgx L~V~�o3|.V�٫�5�'iJ�`J\i�c@EI�/��'jMX��og2�d�
�p���������4͊0%4��wHz���r9���y}a*6n��,U���[m�41�
��m�ۦLa���w;)�C�����Yw�4�MR��qN0)W�7�}>s7������料{��~����i��R��II�;8��M0"��~��ћ[u9칉�{��=5���o���uk�T�{9Kp�I��2��J�����\=s��w�E�����u򬽯u�T��Z'�ϪhmV����b��]A���*��-tiW)[W�n^��hWt�����0#J^SGv}�{Vf�!\�WK2����{�x��v���몖�^٦~�˯�\n�Ό���R�ɰ��T39僆�5@�����aj�ǖ�e��Y�u:q����,�q�n��ڪ�e)��kf�w�w�\v�������t��ec=w�O���)���KTe�_[�a�������V�fi�3�]걫TWۛ8�qՋ+�;�R�u�]r��]�� �"�͖�]R��]ҍ�=�Yǘ�d��OU�*��	���G�G_��ps㢦�M�y��ମ�SsAݾ�+2Cs7w9��D�ز�z�;͵8f�o�}�-,��8e�h�#X9�mt��sy�v&�B�U��앇]��¦�7����˫���w��T�I���U�0�^Y��,c�"ݽ�"ɹ����l9JZ{{���ַ��Ęn�5G�6ku��/��A�eS��6�	A��]�퓭���v�^B����ղţ�W�n�z�7z��m��Z�_evo}��+X9�O&5�`�{��U�
Ha���q��½�Gk�:_3����k+z��Vkl݊"�ڽ�c�8��������5�sz��s�Q>�*?B&�^����8���/s[�)�t{�p-�+t�ȧR��܏.2��_S]u�pˇ�u	n�Z]�MV�ެ�l!47�N�b%7��30S�Y�̵�)寧����w�Ë��X!׶�����q\"m�2��[g*ed�r�+;����0���g!�#�!��M�P�!�sͷj͵f�h9XE�?Y���%4��{f�9ͦ�&ӌ�mYN�����ltY��i漻瓞�l�0-mm�,���qIx	5��nK&8� uY7[�p ��mmnQ�m��,JN�/;9�ݞl�p�G6����ebS���il��Z�ݖvu�̳[BmZA-Ĝqy�X�Kku�m[j�(��4�.�KnɶY��m՜3p�t���k1�Iq�֝8I��9ȉ"��YE�dei�؋Ψ������qYX��tt�bQ�w6�kYȇp�n�Duyhym�ȗ�t�G�p�GGI[j�N��&���2�������َ�C,���mN�*�^b�;���m׶��:�;˽I;�":ˬ#��w";x{2�ޮߖ_4)r�JC�`JM>I��=�߻wy��NU�`N����X�{ެ�1Oe{���ܚ�w��k|J��|��{9�����h
��*�L"�0"��h+�r}6-�ԩq�o(T}��yz^]Z=�'�^��kp��ӍI�������fHo�+�P���ژn���s{F&e�p��V��UH�8�UWj>��M��&�e�q�aJ�����wT�]8?zu�w���<,M���3���4�أ0����(�Rd�7��~�L����)��E���(b��/oW=Y1}�/Ԉ2u������ɭ����Ƭ�*���\M>Q0'3�V0��7��sUA��}�y$��h�uk/g)n���`R����wd�����_.����}��3	M4ñ�@w�����_����ȩ5���q�^�e]��w�a����Ϲ�;�p���l�A���Cۂ;7Ϯ�!��s4j��W��Ų�0��z���)�K�Z���5f�I�ꉁ9I�P��&f��sNǽ���m��o9镻7�Ozg���|w��>f��)4~=�;}��n���PD��@�Z�l��l�p\Y[fX���V]���F�	��2ܨ��_��R|zdJ�lQ�8�:�YE���9ǚ;|ӊL�џ��� #'�Y�S�\Zi�ñ5�*۞���F�\VAuwut�R�M���z�Ro�"�4�b�	���S����Z7ꤋ�"o4��J����@R��T����yz�y�1u��z�uM��~~�k0�[O�;h
T��}�/��t"�4_T����@R���Q[^372��靃G��W��Dpd̖3v�����L;�*�`Ofg}�g���zw}�w7d�z.����_�EI��g Z���*ޯO,b�<�2�רv�F��ɧ���#v�?9�Ρ��Wj�E�_���gl�Vk�՟}{��M��fŮ\�H�"�$p�-MV(�FD҃vR�6l!r.�K�͗f+��[m��nW��!n��������K�����4�s..�iM��Zce3T4e��Ga]ՠ�+.چ�M�2ؖ��)4���ej��R��a]��QТ�(�k@�%j�r�i0���Ț�d�Ai�(��c2�$�&�T
(����7�����|ĭyѵ[#F5�0�LU�uL�]-�\��`�L���R3y4������e�y�J�A�D*7M[��_L�f���L�驯i�[���ؚy�R��vRi�� �A��/�*z��*^��}��NdW���J����E}����／j�������,���e��B�f^��͡�+����+�Ki��Z��Z����_�rV�f�����|=��7��Win�8��+h:���V\�W��5�4N4*�j߾��e4��zg�M�M;��D�Cٯs#�z���}Y��毸�Ԉ��U�"��E�㹽�&��E�����>�Q�zgޯ,���͔�kp�\h$���Ѕ�/��s�^�ejꊫ�$��;B7Fcj�.A�np�^p�7��EM��l~����S�{O��*L	M6 �vf=����|=�mLX/d�Zi��Q<	M> )SA�<�'�~��E�̝�?��T������y�X2�����ZU���M�`�T�ZF߳o��jg�M=�ќh��O�����}0r����W.����r��V��WУv��ޙ��Zn���>`R����kz=>T�}ؚ�eW76*M4F��@R��S���=7��^�{l���C����� �N�MS�
T���:��|��n�m&�>
T�%&�a،�a��z.�����'!����<y��?�N�/���)RMQ6����������,��W�4���U��>�Ͼ�x�5`W ��a�O����z>�2�'}ֻR�s��XZ���q�d5���a�bU��B1��Le�f,�Σ}��N�E\Mi�=ƚ���S�u=Sd���=��{*��VA�t��a'��)4�Ě+�E���M�'�Ji�;�e��^k�/�|2�����{���Y���d�)���SMJ�	8�-�~��{����X������ۤ����=dw��6]j�Y�$�e,=5�fʪ�#N�j7��ܴa|��J����Q]���7/��y�f���A/Ծ;�Y��I��v&���.����^�̋�5�Q�l�4�����ڮ��ٞ�>��uk�%&��ۯ�����G�<��M�ExR��ƛ�����6���gp�2����ó��{�*�����g�e�&rrǼ�=ܬ;���ۼ��D���������nfz�4m�W6�t�6��16f�"UL�n�7^���7(�fL���;����Be�����U�^#��5�gμ�/��rsBol;8��p�58g(���yFW�����nI��vvv�/`�g����l��Ji���Me?�[���U9�W�R�=	I��oy8*�R ��^��o��W�����sٿt~�&�x�����Q�+�>J�AU��6z�W�}of�s��R���)�"�O{�1������W1xK� DּPc��wy]v1{�᫥Ou���1��6*�Ͳ5%���_e2WQ��e^�x[����[�4�;�&�2n�uw���qL7�U�.{}~�N( �&�y��MT�`EM0�&�W����-���)W�6m9�=y��.���$`�nU/nQHfd�VfI{�]�����޾����ɝ��a�.&{A&-LH�a���g����o��kW!��O���!?��c�l;,�
T#��5����2�ܪ�os#��/%r�=� }ܯ�wX�@E`J�i�*������|b^���==��;.g{y�f���~~����b���Z]_���f�-N}ؓ[�T�w�Uƚ�SMK��n���g�a'��䖩emzk����C� ~>�W�+ҒN&�����T~/��w�4���Uǆ�|�f�1�n`�_��{�M<�5�>���
���W���+��iRh"�Ri�)Rh�����m���}�_����X�e�����j�k�7{ؓM`R���ue���߾�������k����iP���w��?TC���,lmu�ں�or�f>�Nm݊=��ӏ�C�7q&6h�����Zx_������'��ip����
 h��̰�gR�9��i��c&��T�$�� n�3��nR��]��Ć�I�,��T�����Ҙ3���u��S)K.��XD&�%5���-ˬ݆�e�316�*-��=L:����X1�30T�,�뵱���m3Sb�ԷQ�,�\n��9�N ��U2��M.�cAnh��]Xv%`���L�����ߴ#4M�B�b4��zɪ��\F�@����m��J%��Jj.S=��o^io�|f��?1���@R�=ݝ6���̛���q�Y1\;�v�����%���$�VA=ԁ��kw�q�޵����`Aӳ�Y�S�{��ᗴ�x��L7d��2y|N��g��9V�Pw:H���X�yN>Ksח>���.d��Ȯ���	�������2ׁ�@��T��ƛ�4R��_���}���^M="�i�J��Ίj����o|]y]jQ4�rW̢���V���*h����J����0)W�U߳�OtC�Hdo����ys�Ϻ?}`�����݊&�����߯	��u?f*�V61ׅ،m�5��R���Z��6��H���6]��i�|��\M�\��Y�J�	8������������S-x�����Ͻ~=�7��Ϸ)S��M4ñ4T��/�'���|������l�{��e�w���8��Zip���Ǌ����ݛғ�/���0n�Ya=�g,��-�o�(q��f�T��׼���X��l#�������^W]Z��Ji�p�\h=M����Z�~�\e즚f�q4�,�__Ǻ���AC��.���r�h~������^EI4oT�SL
T�������t�ş3��72�q�$��x��R�Y��oǾ��ϪkM��4��z�2fͬ^y�)������N0%Z��w�0'�r�D&m͏k�3}y��/�+�Q>2�RM>n�����T�o����X�9�M�XC]]B7Gk c6eeGl���#[�f{2ntƬA-����:�/��e�iJ���v,0¨��+�[
+���]�X˖������~�X+�"����o[Ƞn��Gy/��7�7T�W����{�=����ӽ�i�0�L	r}�w�]���RNﳍ�I�H� �0%&� ��ޓ>S�.t+\�}���{.��į.�ޚ/����`�<�Jʨ�.�_�^Vͽ:S%�d���tHr�,3)��|����De�:�^�3�+����SOp�M�`R�����b��Y�0{�ݬ�}��,�VC�ŀaP��+����=�ټ����*�i��/}����E׭N'��^�[A��`R�4>�oE[�Y/���Wf��Խ~���z�w*���{ɘW ��'����C\X�d�V�v�Q��^V8i�l֪�L�L\WU�%��ˢ�jO޿y2n��RM5�Q�)4��̏]m��t���+hy�OC�x.��g;�h$��&�0�)�����g�=ۜ��{0*;�w��_Ǹ{6��aq��b�0!�y�����"��ʒ�z���&�i9@R��)ƀ�wp_{����u���Yc�ٞyٯ�K���~�A��_�	I�ñ�
�)I������X�[�D��M4*OwJ�׿eo�Jy����������=��Iw��/.���Ѯn�VtOG��n�B�޶�]�"j�#]Sta����'-�u�t!u˻��\�gP�lUbT�,Jf%�ok@�'�[�*`JM6�0)Se'��L�;�u݀zS���k�V���.��GG�}�T���Q0%&��>�4�=��}����˭E�0��#J[��Ti<�q[�����y��"*���	qÛ�4:�Mkw(�fL�*/p�>���z��UMM|��k��}J��|�4�
T��+��ؚ�I���Rg+�y5|�B�.w�i�e���:�~ɾ�)�g���pܔ��"��
�ugY�1�v��|}yb����=��}���w&~�[*�Mﺭf4�==��z�U�;,���.-��ȩ4��Q�9@R�GuL��YgR�=LG��{W�E\/p�>���]�2�kM;����r<���K�=ݕ���ƀ�Ri� A�A�QV���y�wtyy}~��>��0�����Lܔ���I� ����r�y�x՝V�Uf���� �q��;����R�J!KWJGpk��K*����M-MŶ76�B�!g�/�9T�
'n�.��+Ӱ��vg`]"�s�|s�'weT_^v�]|u	e���x�r���ZO�|�H��M�}rC[��X���p[�sVX�^M�n�ѹ;]jFì��¬f�x��N�tk)�v��Kʧק��O
�B��ٹ�Ʋ��v;qm�+�ͻMP��ۧ�t�,���𤫴�ѻ�cQ�K�c��v�Y��)���X�V�nN����oo�{��#���Oh�f,o�_1V�-�ӿS��ɨ���ų���sY��u�9�Y���OAU]$�*��̅���^�Gl�Y�Mo�ClB�+��l���ղ��v�f���S�)ݜt�8�!�P�c�W`z��Th��-Wj��������=U�6�n&QD�w�ٛ�є؝��ÔUF��j'�rl�\�Ǘ�x�
�f�j��m��fݱ7 ��H�ŷ�.*���Q�$���K�;Y¬�}�8�E�Z8�%mХ+wk\�:�D���}����t��1�<y���FL۽m�]8ާY�3����k�/	�unʺ� \6:ڎsu���7i���,j5��N��eiM�b7�a8+Ŕ��C�S7L�ܝ��h��r����v�9�4��z9��lVH��'{/�F�z��V�*�j�Oj�o�Q�He����B�����%�Hmb�J���m�ќ�E��'�خS,�䷩������N����z���������g�ds�^Yܝn�ft�����ڈ��mXH&d9���ۛ�;�"�09�Ҳ;��&n�8���o^�㳰�,��#��8����s�;3�N:���ӣ�{onú͍�Y�ܻ2l�`tf��{gGNu��-��G��'�Y���s�����p^��I�4sn+,.���h'^��*L�:�Z�;���K	����Ө�[�$�lg�mlՙZqGt���vqm��q퇭۩9(rH��B�ʓ�V�ٽ��.�Yf�u�vѥ�ZW��u�w�[7[j�"s��ݥ�e�F�VqNIE����$yaXu�i�qXm��΋���N9��vY�a�'�yv���-�(��3�}�_��+l�"������Z1M��Cl��c�1�&v��l�(Y��s̢�v�M`a	mJ�帎JLe����.,�Ae��4(� 0B�tЦ1"A��
iK��8��Pl6R�0�Ys�0̣a�JY[�������n,h8��^6��u3`C���F�u�JL�� l�L���Ml1bdf�̹uRk�ָ1��������!npZ3X;3[0ˆ0�;1��+�Bc��L\SSe�]l0�����m�Θ�t��P@j�(Ě�G���n�6͗p.-;E�J����K �k��P[�:�!Bcl:Q�clA&d̶]��,P��2ݫ�D�d8\i�"��-�:�c���j&]T��iF��W[� L�kj봴�\$�"�15���M���֥�]�+5��k���)t�Ś� :�JQM7ԥ��T 	cB�Ⱥ��u��mu�2K�ӉvҌ�^��x���\\Ё�g2��R���W��[�-�c�.����y���QKF��LLl�v�5��r�!�y����b�#e�� 2��q��tL9�b\��X3[�cؖ`׌H:[l��JT��E�յ�4�G��Wb�QeK�T��,��[r�L��L���usu���F2�0���MP(Y�i+mM��\�5���Pi�,��УֻE����w$���]�R]2�FgѥH�.r�JJ��D����	���witM��D	���Zf	A�ƺ���e��20�R"K]`9BKu���LY�#�A�I�1����t�`�[��tk�-��ie�f&��Y�Y]��֛gĲ���GPEGb�r]��Zec�m�st��ĵ��vқ���P�Ir����AX��auh�b��.�rXE��#��b^Rk.?��G�{RP)j��Ri�j1�@T�v{&�jA�m9Ε-�$BUu�F[\��l՛:�V�+5��Ғ�T������1eH�#����YX����(i��U�U&r�`є���2��u�	��!N��%��َ�c9!��j�D�RZaųT,��m�-Z����g%���#,&�!,$,��ܶ�u#�]�Q�ˠPwmY������֜��j;2�CZ�,VX b�$�ZmDQV�G5��j���X��[BӐS85ݫ���9�Ti��ZM�fŖ��[��N6n��l4N\�k��:*J����Ľ�.̦Ø��}�>��J���b���%t��FT*�Yh��H�����UM�d����i攩&�q�e���5��J�α#����i�.mh�!I4��Q�JM0)SA' ��^�cYʏV�`�D�|C��X������g��]�2�oM����OQ�ޢW��1bw;T]*M0"���`Jh	ˠ��'�lS׾�C:���d��߂��+p�I��p��8�j�sm��]�;�4��R��6Ri��倂�z;��%�:ď�	��1e��y�����h!�6�(�SL
T�����n{۸p�l���N�����ݮ�����}����\`JI�ý�x������k����[4%����H,SS
@��L���6[V�X�Ir>Ҫ���_e�M�SO6(���`Wҫ���x��+�Qv��vō��>i��Ҥ��y�%��;�y�~�8<W���f��Z��GD"�������v��1�I�^��(9M�]!v�m�gz�Zu�gX9��Y�(<K��wV�{�k=���aج��w�޹���f^���SOv(��ݧ)���_����*M{b���J�@EI����W%��k���=O���9�w|�E.׾?o��)R`JM6��"��l���m�M<����i�
T�ҫ����������{�Um@��T^9`^��:u�`JM>0�M0)Sw�����|�gs���g��h�=Xyf^���"�5���i�K�`}�����/bq���cf��fj�٭ܯ/U%VƼ�dY�4^�ZW.w����S�\���)W��ni��g{���>�]��k��|�AካZ�R{����y&T�7�b��wc�,���
T��Q�W���#3=�u�4��M4�
T�y��߉�/�r�Kȼ�^�Rzw�
T���|a�O�o��j�7�k��]|\�f�9�#캪@�ϑ�ḶF�����u/Z���=�����Gܫ-�;���&�E��/G���gvu}Z1�������̽T�x��[�Q�8V�A�=u����Vr�W/T�{U����oy�R���5Wm��ݫ�e�2�s_����E��~�)y;2Ri����I�"T�(�X���SFu�_b���'���:��|nfg���&��I��*MS�
E�~Σ��{��w9Q5]t�,�XÉu�ሢ��s�T����L�`��~��&��5�EI�+�4ó XW�{g�[s�M�_Ț�Um�g}���}qN<6Ri�) �"i�JMg�}������֕���R�ni�����r��&UMM4����&�VYB��O��ƽ~�R|xRh:�SMK�h��-z�Lȼ����N��n���=�)���J�A�@R��׽���B���lY���{��p���ql��[;D���Y��r���W�gq�{2�^e_^R.��ڠnVs�fЮ��:�ߡx��������V��6j8wݻ"�/3�Sߖ�u<��E����H�`J�MJ��b�3�ڷ�7����(��3J���nצ��˛��C�w��*I�+�6�}�V�J}��<�"ٖl�T�T��+nU�l�[�
�ʺY�m���Rv%�:�}��w�*M0�&�J����ӽGۇYe�\�G.��J\�`f�9�]Ҧ��' �M0�k=�/ڎ6���=Wk)>|�A�Jwp��Vmv������}�*M5�Q�&Ww�߹߶,kv(����4q�Kwgw��~��S>�WG�6�Q�dʩ�O��C
T�SM0�h	����M9QG����:��H;ݚL��)���TY~����C^@�~VExC*��8bÿ,M}�8�v���bi�J��VP�v�{e��HOH"�7����d�f�O�SO�E��`R��]�X��V�cY2sg�l��;�U�ʲ�Ϧyy5�{�=�V�S'���Yft��X�K_>�b^��m�	��k��7cA~��~���'�M������X�����G83u4�o]�-�$ (�t44�ڰrCr1�ZK�J��DΆ�Yl�	a��# -3pk��T֖��9`��n��A�p�#v@.���i)+	�єM���$5����T���DKV�I��kDM�9�c���͗�j���lc\�,�r�RV)4�z�]+�#�TG�K��wik ]5c��>}�feu�wXC]J@��532�۝Ρ���7et�I\�������zhA���'߿4D��EH��i�ߏYߌ�&UN[��u�����:�7=���[O�;�<��EI�Z���/����s+e���T����ӽ��fy\ؚf䦞�J�h�o�o�ʕ��ܖ�ON�\Zi�0�m�M�n�V��:Њp����Y;D�����&��D���@RA���γ6=�&�͊�k	8�*74�}�_��t}�_x�6��laΌpÏ��o�g)�bh&������N�]A圪�*{�U����K3�樛/e&�7
T�I�r�F['�=���|p�T��,��&��"��L����6���v���]��r�T�:���[M2�ȳ
T����S��]Q�j���I͡Q�������4��S�se4��I��&��Ϲa��;�����Ta�cYt�kz�9��E�su9sD�(�}]�Js�)_e;FN�S��6;}j�"�x���k���v�]J��&�E%�7�N<ݥ\74�}�_���2˙U9��{33(������w�Lc���ޔ�6J�L"�`Ji�K;O���^b�}^��������լܜ��RA�ƀ�-5�ݒ���'�]Ě�⧡)>lQ�ez����I�f��X����n�֟7v�q4D�������]|^���.�RW��O���/W�Ys*��{{i�J��O�:���ܱ�>~��l�I�/31a(ESlƅ�r�k,��a�R�8��4U*�⹻K2�*�I�ɤ�h
T��T�z?�G�y\���w�w��>�#��wn�w�S̥�����yR8�����l��f��]�/���G��'`�!��Y܂=ܽ�~ܞ��,�v�{(��o&���P32IO��,��]�N�絔�5	ٕ}��z�ui���Z����5�O(6������}��y*�Jpe꫄]RK۪��]hN������gG�K��;�@�;��&�4�a��N�񣿩w���<��݊�h��4��MK^�B�{�����}.t���١�l���*7�)&nʜ|�iSRi��i�\L�nwI^��}2�o
��S�<����؅4�0%&���O��L�'�~Y��W��M!�+kqa�<�������6��K*�N���_}�O<Ji�0�I���
V;���4��9�gG�K��%����Ⱦ[]���)S�%q�ó��)Ri���B�:���B�U�Ɨ����c���T����@u��Y6'��l�n��yy�z8u��r�Gn�s�>��K���0%4�v��}_;��~�ǳon�hյ�����|��U&���4�0'+��,;�Q0筴|�%�Ś���ԩ��8�*F�O���E���.eT�	�R"���}8^eﲰX�:ڂg�䅼�^��0s�9�!V���5sQ����V������]<�{������g����]ů�e&�{��8J�(�/�	������,(�J��ɵ/{�=���3<�ujg�Ri��{��ϛ��{�����-�ߜ�A�R���3t�cb���)�0X������v�[�Ȑ�{����e��l�y��L	\i����b�/�u�>Yy����^f�m]sr���Zw �w��AH
UƂD�������y����^Mo��ksiQ���ۘ��^�Ye�UMwԁ�X��w*ڣ�]�b��Y(���M}d�[O�' �i�)w�{�:g��*ݽ۵k��N�D^@��/���$S�¸�חb������!�f�|a�x	�Ŕ^=�����36��;rP¶��{�n��MO6������������,�2�o�&�n�_��fR�n�n�F���]eT�4߷���*`J|�9�n�=;jR�>�K=�g>���Cu�U���&��Q&��]k�J}��ҌU�D�ub�� ���9*P���A���W;u�N�s/�o��� OYo�l�-d�f#��)޲��M	+Ժ.���7iQ���k	�`c`���k)��2Xd�ι�P���l�nf�(�kf-�0s�\M�أ�a���aÅ���clu5��ڎ�f%� �Բ�L�6,*U�YU�-t��cn�İL���6��r����]�Մn��]q�14îX��i4,h�3/�����n�.2�[�tuk���6S&(�n�oM�E�F���8F(�W��;�q�D���)R��λ��ם�'G�/��@�{~�;yJ�͜�`R���ƚa�|m���Im�3������i���t�c���][��H��lB��PG����59��Ů��*Mg�M;�r�)Rh;Ȁ�7暾�3�3=6�T�bt:�j�������@W ��i�bMT����~)m�ٿg���Ϣ֟>Ȣw�)�*���wOկ=�'G�/�y��j���g�wJr���R|�,ȣ�����y�P`ͥ��1]��'��s�7�?礠c6���X˻���C���3��=��U"�al�@b	D�b1���m��U�cK཈��Dr���h/��l�'3�MT�#���d׻�w�̝H�H��A��H"@�"FsS;�X�˫�Vn�13����4��]Q�go���TU�Bd|rê�x��d�T��Y�fJ/ֶ��{��GoU��}}��m8����\�ŏWt]gҵ��d��E���oD,$�g�=�vk��VO��sv�/{y�D�2SM<��hZ+��Z邦�W�'V��7�	�hXD��H~�X�D��5��˞��\-u|���D�/��>}�u�01=���n�9���C�-���徹�0y���� ��2 ���:^=�7d�hფ�c��ˬ�jy��;��'�H����$��D3��f�TUA�����h�7&�d���VڡB�!�5Dƚ��]�"�|��[��D�+ �%/��
��bx���������37*ЄzP@���%�"D� �K�7=9y���h���@/��O>�ۘ��Nw.׈?� ���!3t1���]ڱc��|�F?fICw*�8�wrpX}4m{L�<���=wN�e���F��=�QM�i��͝�M\�8*�nSԉ�G�X��2���M��Ki��]�e�i:R�.���iLª����uΧ̊'I�t��f,��V�q��=A>¯�VUі)�f�jp�p)�������hge�VN��q����aw/������\�S�cDڸj�G����u`��ƃ3\Q��K"��er�Fw=.�nK�� �R���+wG"�k�R�!۷�:�I�����6�2�k��G��Ҹ�{��������uF���/]c ��V�͡��q���:iL;���&[���絛���nn�z���`�f��Q���9+3�;^�ܮ.f�����y���z�PC�q0�R�T2��nt;��ژ�zʩ��s&�b�b�A�)me��H�:;��T(�̬��:�'�KO(�t�Â1w�1E�����P�{�3-�S��E\�ʀߦ�+��q�m�aߡ��P�������Wʝ���p�4�J�NɅ]�E-tl60,�f�}�%�y��l���jS��:Δ
��'J���n��<#�\���˺�ִ^���6%�x��f��R�o3��5ko�J,�%��˾dco��1\Zڪ��M�������k�D��-9��b��u�v���_b�;����{�o<�Z�f�s;p��y�щm��V]��ʏv7G�â������l[7���8*Q*�O��r<�.܀��]�ym�K~&�'KGB5)�����
W���"o��6�I�m��Ycn���-K���dE�ì�α��t%�'!��+o���wf"q�i{v8����r�8��жΑG(��%�췽��	��e�Lˊڷ,�t,�^��"�Q��8C����d�@�kn�%I����HrE��۰�ٲ[fv�����q��Fi�fGq܎t���ptBql����Y�h2�p�k��ӣ�8H� �8��N6�yyל�]9	�m�,�q�彛m�p��k���v�z{bt���^g�
<�����e�l��e�Çeas��[u�yvC�u���mvYDQvI�E��Mn�4��BF�wS7)P�TU
(�HE%y�}�|&>�N�[ؖ<��C.�Jeܒ��ʾ�͹�O3����]�4��ge��feB�k�h;~��B���5��vϝ�:ŀD� A��Ibȓz�u��fw}@{�Bo�z��`c�&7��e�	�W�D�+��%}n�d��V\�$錒.ź���JL�(D#2Р0MQ��Э% �ph@��*�CÞ��}!G�Iw˻��Fd�O���c�x"��J��n�TX�^�����B��@�� �H�p��m�ӱm#���M7gf�"�;����w`o� A�п�=FJ�7��lҭ�N�����7�7�
B��]ʔ˹̔�νU�7o�뭙��xMo���^ �wԈ"DH��	��%�N	��nH�ա`�t�2K{�Z���s��}�^���W��u��ܻZ�T�{�R�:�/��D���IbP�w[Ϻq�^�UZ��#�{X�����U���x:�ǧ�S�2��y(U�o�pA����[�N��P���$VAJ�H�H�h�x�+lp7�Rw�L�/1<s���7�3bA辒��$�3b�oy��{em������6A30Bj�^&��QST��v�H-�5��("v4��܈��=�w$��$��fT{9��i5��s-x�
>��u�ц� �j�����)$Hd�Y��pM�0��Î�i�m!�����a���M���g����[�\�s�*�}$��ɡ�{)%�+%�p��z���{�~bx�����|f�,��E���I�$Az^Q��!�dH���_N�+�}�j�]��}SRi�og/P�F�������K�$Ad�YP_+{&t�^�T�v/��>���w�en>�^}������2!�6��y�)�/\�=s{���W�}Zp����3��~��t��Ǵ�=�4\7�w���ܮ3Y�3��/'(ꬅƪ����g^��|wߞ�'��%�-��6�3M-qDb�,\��[�*�vR�+�ٌ�e/3+)�CnYjW�-C[un��A8,Fmb�� 4�3iV%L�����{B۳&�v��Ĥ�Ȑ�\^�]��s�6�
�P���Q("!p�9s��5wii��m�ࡡ�]E��#���L6\�ËM��h��{�thY��Fhf]a��Ȅ�I���.�|�������+55-/'k��q%�1�]�uRPZ"�2�UBs,�U߽:�����$���i�<Θ��u��\%���y;�-��9Պ�n�5�g� A�X�$H%}�&�u�����5|~q<����`c�&79��^���H���=-Ua�p�3������@�腀A�� �,{��8�Ov1�wS��ݕ�g;hJ�Čk=�}	L��]��ׇ{�u�d/�o��Ưz�O4�ƛ���d�g��+��`o�/���;1��w�>�|���/�$Ad�A�X�$���U�0���^|��A���wŎ���s1xN�� Ȃ2Edd�����}~��D��2ꃚ1ΎюfJM]��P��ƈ1�) P�֦�Qebd�*�П=}�Y}���A���X�=]�u�?S�{+^�v"�@���Lca�r� �=�`��J�H��%"�~qx�n�ݮ��7�s�5�uu��
�f
�o�vw;����޲k���j�E�W��i��q���}�3�W���ww,g�q�ض���Շ�;���|I�ϲ�����{"�4Ǣ�X32�欬����,�� ~/���H��D,���ۃ,�����B����s1�_GC�"�A2RH�w{psjK�hi�ǥ/�"Ib�]�u�3�~�{9؋�}�J�w�U�n��"D�+?IH�� d��=��:��7�7�Ce�s���d]�{�#��͸Wq��wtm�]��]�ϟ=9�h����L&�[R(h	�f�1H�@mZ�6���<��|�Y~~e����	5}%'�r�v���з9��^^{Z��il�%\A� [�AJ_"@�"˚��2<,R�%qN��L���{u����K&���v&��J�w��ٻ}!B�%n��1���z�]Ťd��,m�΢���گُ�������Ȉ�����R����u�U��;�Jž�O}0-��>������oKcI�-��ǹ���d]���f�)1�nU�pc.�e�tfNKn&"�G�����2)�,!۩��/U�S1x�wԾ#
�;�{�W�B�Š�;謂u/�� L� �@�@��x�w����F'��o��]c���^@��"9����D*���G�'W�o��]3(ʖ,��1FԘ��RZ�gB��i����׫��)�M�g�c{��z�wsL`d���q}��:~싺ĞB��"�iܹ=aL@\����X����2R#8�o��{��7�/������V�eԧ���o1x����~A$FK8���;�&OMu�,��^�d����S��wru��+����}�A�߽u�{��~_g��ϬYW�	�E�盔e��u���A����;4�����Z}�)foL͈X"�RU�
uxm�*��h*Z�)�N�Y�*c7Rr몹V��;�貫�g�E��e�fpE��&0�����s\����Ne�v���AYu��z����˹R7w�]��v�.�gI��-�ˊV�M���Ǫ�W�髍>�|��A d���R���:�W�dÒ����e�0Zu6��m%ư���ii+3Jf�V.��<3y�4���2R �,Y��;.��z��;�9*Q#�{k��@wr�J$VAJ@�el�^-O>�v,~ݔ�3;9������>���f��/��)�c�{�{<�rX�gR%�"D�2!bߵ^���9~��3n�r�N����A}H���]ʠwq)�s%�]k��qf���|��T�X}]W��>�������'���>�7�&z�Iw*��c%|�A$X�g����,�R��n_67�������FJ@�$����8�9�Y�WҾ<p}��g������C}Դj���k�0��e�ys�Yu[��Sw/H��Uvn��~�[�N?7�{�_z��~�-�Y��#+J	Gi��;[�s�1�De�ʅɛ�b�ՆĤ�y�h�͇CL��f�iet-6m�+�辡=e)��2�	��  ,��� e�)Y�h(8��#���m�W�<��[(�K+hf��c�ٗUH��7��޲��p:]&ִ���C�[��4PJ��i��ErK�����)�򄴹5�CvE4��iR���H������Ϧ�f9��b�!+H������ˆe�]b�f�M���D{z�O�|�2��,%}%�r<��tN����7��v87��� �})"@�"�'b�٨�Vu�8�R �"w	�t���Oy��3���� �>�dI�G�u٤EV+�_L���A��iE��i�Y�my��=z�b=[��<�Oa��>��ր�辒��.�]�'������ۨ��wh�e�)�Ȧ�
����b�y�����ƛ��q���ަG?�q23�$���FJ���M7D��,_�x{��=��-o>�&P�>�@�<�ł$K�"
��/z�v�5�f��"� ��h?"�:�lH]TetU�7h2�E9zƐb$6%#����}���p� d��&JC�����<�Oa��>�w{���R� 7��A�Ib� �2R ���a=�Ch���[Ph��.�X0"eꐭ���m�;�ñ=�v,V��6q��xA�藎9]��� ���ٹ��g���_|rq�E�a�b�y����֟�ƌ�y�+�P��� �JDf��;܀�"�J��X���K���3Ѝ�6���bg�@�m"���/�� ��/�fn��L��ſA�������Y�'���'W�5��T�8w��ލ��T�a��(w!#w�wrReۮ�+ynP��Ϗ�h^��m)FA�v��/|A��R �_I�AJ�����O_?_�q���a3]�bm136����!u�r�mpF�U��W��M6�#B{���e���7XD� d�AK=]�WY>�iooF&y
�^�.����� �2/��A+�7�����m�,���zWI�iL}y�_T�� ͈�d�j�bM�W��ݶ,�� L�� �,X"J�	��^U�w���T'��F+=B��+����U���������P(��u���՝YPjnĬEUŏ7�Y��H��\۸/ɥ��8l�������HGD�/�%"$Hn}պ�9��,�r�c���+#0��g�����-g�D����6���gJ�����G:�H�2E`��""ݗ��
���@<��j�={��_T����͈X#Ҿ���%��Դh�{=�ȶ�L:�hj�fpJ��r����Z��S]����:�����.�+�I���)��$��p�M.'���;oo�-U��w�#�7j�A���_Y����H����<z_���2u�]�WY��g�\��	�h��,y좆]�#��?lǋ{;˚1�D�2�U��X�w��w��&�6J�+���K≧�ȕO3��X�$@!�K�Ú�[�C~BȜ��D=Ϻ�-��xl������_�����g����w�c��@�A��u�L��]���,�g;9^�ȱ�^u��ܱ!Y݄g��M�CH�ML�Um��8�V'�H$���h"J�Z7��lz�i3�������2WL�qǱ��'�K�>�`���"ܡ�.�y�%�6��D�Vh]�j�Քm��"K���m�´��58Ůp�ȿ��B��Ў���}��K��Z�:�7������?l5Kb��U�9�"�Xh%"�>;�^���#u��/wwZ�v���d��^?l�#��H�����w�:Dw%�����}%`%��#_]`n�on}g]I��8�0�}:�A���D���0����gs(�BّGa9I�v#0n�^��oB���;���Ψ�w�{��)ض0��(eܒ��YwrS.�/N7�w�I	�Mn�/[�c�7]��u���_X-�䐐�%��!!K��BB��$��	($��!!K��	_�$$ I"BB��$����!!K��	_�$$ I|�$�HH@��$$ IpHH@��RBB��I	_�HH@��D��	/�HH@�𐐁%��(+$�k,��B ,[+�B ��������>�PH�P P
����IUP)J$ ��QP"T�TT_c"	��x}%֣$��u�����פbb��X�Z�R���j
���Sm�w��n��Jx,�_9�o�{;뼻�vH���2�����nW}>!N��vUqA�  l`�6�%)�s�E.IN3*���7Q�
�AR-���n��j���u��mAA��y�$�lw9]V�,XD��b1���6-���P    Sɠ)II4 h2@FFЊ~F"T�4���0��d �5O̪���10L���!�0l�P��i��1�F i���%=�L����C@ ��� ) �&M6��=SOESd ��mI�zzy��=��� �b��(��M�"(�� (� �b���Co�Ȳ4�����f���F�C���]���`�&��@E0���q@�&�@�!
 �DQG�O?����k�Y����/���"�Ob=y4Z�4�A��}�w�>�t�z}�||�L��1\џ��ߢS~���o߾��ީ��k�eC��~��@[�5�
�6��U�e�f|\�]�{��K�Al:E^�l�������XQ�,뻛Y��E�[�q�(h�r�-J�@q7R��Rɗ�جT�;�N��y+F�Gp҄S�Y�*Ƌ��M[�����u�6��. ���Z
*��#Y�M�&�l+�����[��x�:4��qyB��U�UaU����@n����]��ЫUm�̫�c����Yk/*�d�@i,i��N%��Vd�I�����Sb�n�#\�qʲ��g���ɍE�h���D�����֬м�����O%X�xB������ڏ/Ff<�9�c1n�ق�B�1�6Un�J��TI�Yin�)��.H�Y;�N`�9r1�x�pC�p'.Bk"ȚX&]	�Y��ܔ7L`�4�Ĭ@�j���X/)kUz3��� q\0���Y*��P9�7d�w��Kn׭�,ѧ/i�m%��َ9��Y����@��mo�&�,��f�l2��senS��l���L����D=g.kOrV<�\������D���YȆ��hd��V�T�����m�Zn�K6Щ�&�X�P�{0;�Q�#Dn��O�����& ؖ.0X�b�挱��vp�H)Ok]�r�`�`�lf$���ۤ��Yz.�b�3LwVs6�
�F�� /!������km��ͣS���@���M���d�����nnX��^�ӳ7S)�omۻj��<F�����ԩ�=�&�4PV��2
{gv�c�$�aVy�̋E�^hb1�Ң8�b���v��+ǂ�ӭ�ȉq�����I�I�/$Զ��	�.a� `�6�r鵭@7�`)�{oA��Le�y��n" d�e1�uDF
ܡJ��YݹP9�q���E���ړ5��31J$ȭ�9�wr嗇]�.�[Á�`$ ��u��a��Ki��C6]	m,�4�0�DQ�J���-;EGCdຸ�i7���y�ӌ�12�(���Nj�p�Y*'���u2F8�5�j�١^�cnCXd��0�����6��rHQ�f�B�ܵ@c�3Wmm���עh��h\�t�\]��gJ(*�(���S/�D�Z�7�LC�6.޵9�``a��I�v���O�LۻڗK�t���."��l�۽iڶ�v��zQ��R6�����2lY�*���Y[��aރ�6���%e�i��=	:�or̛FZ@��mM <�IGѹ�����8n�ѪGs	�J!����-�+4b����p����LYW��c���X
��R�ʧ�4fj�n)*4M+� <��!���Bb`LR���1�Fg�B	�.����d�B����=���A�M
�m��Jۘ��p�b�rkԴ^	�Z����8��z>T"Ь��YS�X�#t����Yq�Ĩ�V��D֤Ի@-ue�X>��7�F˭����,ͳ/v��V�蛪�=��Z�c*�4iV��Ҩ�4���c�&�4\�Z���|;�pq���6�~���g�>6O�F�^�q��!�>�<�N��~�C�'���:zzu;�N�*{!i
P�V���
QB�T�)@Z@F��
)(D��F�@�hP�Z)T�S����|;z�g���N<��_��"�wH�����<uҠ�Hw��VO�M�DQ�q=O��{��9��s�m*ܸm�,���#|����:�V��kN�"�L�OR�k*�S�ZA�����+20��ˣ����<A��w���T23Tlm����]գrΫ �����5!��
�0��$H�#p�v3"�2����̭�:��H�i��3��T��,'�9����;Xz	�����'iEC9w�~4���u���.�ٳ;^�ǖe�d��a۠��.��%�IzG�d����
m���Gi��pV�)b\/xbIP�l��b5H���"�쭔�=��	b��.�J��:P]���k�3�b���A�Qz�̌)	�Ғ���7���-��U��0)ǮS�m>��>�E�Q��X�L��K�GC���D�U�j����n�.�;�,���PM�~�,��<� x��x�3g*h��������,�<J��eh�SL>�;d�q��X��J؁�S�T�hh׽N!ѱ��ۭ�X�+�L�B�ee,��د(�ѐ���5;�W'��n���X���l��`�6��pM5ʘ�k"簎���Ju��\�LE�U��*��㈈GS��)y�@c6�����Z��b���pi��;6�%/��qwt"}��C�GkO$F+&i��f�V
W�-���X��S�U��3�h��Z\c�MN�6,�U�Yf�K�}�rL�~����l綝�Ȼm��݇�$<8h%u"X�P�`6/^y ;����^���RzFy@fi��H��U�.�7K��|��'�0뒵RRN%��P(k7���X�ҥn����^�F(ԭ,9�-*��)7-m%�{k7eoC�\��o+2V@M��ח�[0������]�9�Z0���ԩ��v�tw�e�6��|(Ÿ"�N5tj����D!K��.�'��B�$,���f���L o�K�3J����Q���Qt�Q��p���r�H��"�JPoGPM�GB��\w;-n8�*${�I�YP&c3{�*+��`e�iɇ�1T[���n#%R��yN.t������u.䩥fZ��:0�ŋn,w׼��n�:����̍�:c=��X�@q�k4����^�ܽ���H�ܴ�A��)7��җk��tU�(i�o���Vp���潽�\O$,=��۬-DK���Z�u�V@�5��b�ب@��o�t�_�:��:~r�5��4��n&�N@&.6�V��6ӆP+`�u�^�P��;
�Wz��p�w�>�6|�ٹ��b������n��v�ĝW  K�rJ�)��P Y��z�@w��2�����)O�����)�-�<t�7xX3squ�f�$����v(�E��/�ݴf�O�"�{�s�04$OVm�]ul^=;V�]v��u��{{Y}�e��e}������)�c�l��6bي���5fgH�)Jx�r����jq�\�����$�;h��ɂ�%oD�/k�
Η6�0��B����P�3Gw���vSA��ݕ�i�m�M	 ����U���Z���Yܕ��[�nH\�Dy�ݕsH�e^�bh���ZS,�ͺ5ڹ��� <=��P5���!Ҷ��K.��C��Ľ̰�>�/l޹��Er����`�� -�W[5ԍX`6�l�e�]-KXPћLke�mr��`5���w[��6fb�å�qL�#s�Nsq����Ņ�h(�WKP����H҄�C-Seڢ3I�Ѝ�m4̵+[L�S�#leT�s�teZZ�ˉmHu��dD&m��9A��r�\�s�-IXm�UM]�S�M�p�ض�h�1R�1n�S�7���Ci\b�-�� ���$W*]�w\gv��M��`�e�+��)s�����]���it�u�(S��#�	V:u��U�X����9��ݣ5k�2Qm�-ƭ�f��8å���E�@��E(�4f�aCk).dl3b��ZTb����9���t����P��v��P��!l"�H��Z���YT�C�f�ʰ�;0j X�.�it�f��fVŻG����n�<�A])5�)�`:jU�2����V+��Z�g���)�v���;6\�뒡k��\J#pf��s�1�WL1�F��K����fb!qLLf����7b�����Jʶ��663c)4�%�ˮ� �0�a�[sbWLd�1MM�a�F#]����]fjKf�iG6gWMnl�e��ph�`�@1]��pM��&u��]\UL�g%{�Ƣ�S���q0�.����gr��]����֒��1�35�Lљ)2@]��5J5K-YL�M&�kMM[a�^y�����5+�r �0��к�Z�ʦ�m���H�s1�!.&2�!6r���76�]R��k��suA6AZ�� v�8���q��[m��iN�HpL�Zޙ�d��[�.��H�ff�؅v���¼\��C(��Y����4�+�Z�nh��"��34t�Sf��%Pv:��EH�h��lݒ7k[��+����4�R������5̈́]�B�i�(T�eX�4�+��[�D��l��	ˢYuat&xX��M����55�;Dq�e�-#�qE��@m��:W�]u��v1����[i)N��N^m��TxԶd,�m��)0��5��K��e5%����k�8ڑ�.*5V�kMA�L��1%)v���Iv(c����S����f�"�j)n&�":�bU�A��f1�YP�#rEQ�US
��z�/���u�n�EȳkJ�E	jފB�4"K ް	mQ�$ E"�l-�Ky�֒��K��*q4
�x�-�m�D�"[�5����ɔ%bBʵE� �
�%#m�cBK�e����5��bJ �+@o���?^v�K˲��ݲ�&��j�n�csXjMCh��Zm�]KjR��ňF���K�R9��!Ɖd�fnj-]m�ۄ��Jf炬�X�DH�3Nci�3Rm�c�qmQsU�;M.��6�PЖ�[۵��P�&���#m��#۬�ZRkf2�4dtά�h�u�:6iF�Y�:V�kJ2�4�u�`;bؚ�c��g:��%"�M��U���u�n����\�0E�vj͓�I�a�c�aR-AYE"J�C��+m
��F"э�P���>���3�Y�Zo����x�ʮՇ�4�fVM�Y�6R�����Ey

L�wT�#G�0\���E`����-�؇&�i�q5h����Rϙ	!�?��)�١�5��]���4���y�V����PD"�:��w�Q]h&�S.Y3e�I!q&�^�X������(��Pӈi;�O
��5���
$��f
N��XW�(���x/=gɋ�\��|��d�}H�%�*�͍�u-�4���u�'�y0ְ�i��:���ξ��%�d��x%��QD*��YI-�9W���?E��mY~�.��w�C�`1eɭɢd�6Z���p�(N������t�kZb}"�����~���MjEhQw�ŝ�xA'G\�|����&�)(���w�������?,
�O�u�>�/<�mu�R�IX�˚�S�6t]ò��P�n�pƪ��J.���mYϞy���5�rWпY���=�_7��"('~��d�(�+���oE�S�7~�m�l�KΘ%q��PZl�!j��Tڒr;�ы�h��v�@ﭹ��O��+���}�8}�̖�i]����E}v����RU	k�l��S�É�(�����_�W�K�1;��E�W�Tv�"�n��W/9�Q>��,��/+����II��v]$�c7Q��l���y��O\բRIsp	#eģp�2�>(�7u6�8auC����tܦz��Q�'^B�S�`�9c��i�=F�xNs���w��C,��pɄ�稦zk�늂�·���SV��)����I&]��뻣����4�������so��t(�;Q�+�A��X7t�WlZ3R:��kvx\�i�`��A�-]"d�0�6���g������-Bx��E\���I�����Ś���������Ix"	'�.�LIEQc{��R/GU�L�le�8-C���v��WmR�K6$s�ޅY��X�=�=����4#�k��#�p�6N�f�.�sV"�jJp�Pa?5��
K���E\e$�� ���Uߒ��#��(�߾|���/������f���Jj����Ǌ_��i�Gz�0	E��v R�ܚH�]��e�I㗉���[F�v���[�(�QU��g=�T�:͝�z޼�κ�z�ݼ{��k:�����i�^],��݇�f9�Y�Hf2B���<�s���<�*�,�S�{\��v�K�۫�*���'
����{-��{�	%��%��b5%BH*$����s�� ����-���b 2E��b�E+JXA�Z!X=KX����E,#�0E��#H5~̲؅����k[�XK׫Im�!���B��`�� h�]���!O�}՗c�Je��I����^M�����X��R��W����,��H%�_^}wH^��qv}E�o=$Rh⸊%^�Yٳ,��`�;o��&D�*���}iy���o�,R)�R��4�a �)�����5�\ݛ �-E��b�Dn�U�i��2Hȷw�b�)^��� �k1�ia%��v����7�I�$=��>@�Ě�B�WPu�"эSX�J���4�-��#�-�s�	��V�S0�y��L5���.�;��(�1��+�DіNG��o��_>={p�c��zw�^�Ԋgg*��*\s;hʇ�.	p�Q0B0��	D$�.QSs�F�iО�ё��;>�W�eآ���U��sp�Q����Y��|Ny՗�E�*�A����XPӂ�5CN��o"[���=3�1�W��ex2{b�ۣgc�!�I��d|?C"����))�j��7�9�q�$�E�*���w���r�@�5����}�W*��Lw���T��X��Q; b��g��w��X�w�D�ͺ�nn�G��<�h"��7�~�� �9�D6�a�7��x��X,Z��l���H�$*<�	 ��B��.t�W6�j%�㑊%���bempG�3�\X~߻�'���q��c���F�k�+���u��-L�nk����[\nk`�d���bP�-��{����a �)������j�&���y�
�{6�٣tL��}ޚ�ر"Z^�S��w7C���o=�e�a��8ɳ��k	tJ������[��N�J�T,?������Q�߿*�(�IC�ߪ���bQd]����C��!vh�r�[ά��oN,ӊCl�%�e(s����v�N%� �JގS)��t�hc9��v�e�Q�����/������_�٤�t�0��J�b�:�q ��������ji�7j�&�(R�NYS�3(���&����"��bSo�=�W��9�C1,�z���$�
���{����Z�矎ZJ8�}�e8`�pCPZl�q��ʺy�9�>�*_���eI�"d����tA�o
�j"
[*�zn�W�h��ܨ��5�[;��j�0�r�hn��l�o<��V�e���o\�]����p��b*��hzEw>ة��T; ��㾘"����+ұ_��;�vn>���Z1������ظ� o���Օ&�p�Яqj�wz3~7E
�Y��r�O�W�Y���y-�e���0��ǹ�
����_9��y��;���=iA�(ѯ$aV�[�P-��[�(��*K-��� JJX�D��(�IKbJ�F[ccXXJ��-lK�*�L���6�ڢЈ�E�qoKz�Z�n.V���=��FK�f��U�(�R��-�q�;���H��3rB�-���e�1i����nc��6u�[�C.�+�`B:U�1�i�N��\�,Yv����X6��pi��V](Q@�Af��rL��jf�0��������wWk�d��f��\D��+Bj�L.ߧ+��@�uM-��f����K�쌡U�&+jm�����b���`l�[t�s*���إ�V�uvc\l+�)�I���Y���m2S$�kV%�')��mY���,�e[��v��d�:\��ζ%��}�O��~��X��
'?^���s|��7l�[��Z��R��� EO���&� ���"#:`�I�h�WC���}W&����nH6�i8�xʝ��-D$�d���l��d����_~�=�*H�>�yXC���&���<�0I�e�;#�d$����9i%g5�d6!&���S&ϛ�=�o¬��p��-��dMk�"���j�E�s;�={�~h��Ó�W�1��I0����}�Vp��5E�]GSs��|�ٵ�)~���mbK1\�bW��2߲@nf��k5���]����v�I���}�՚���|�Ѭ˒�|0���4w P���ɚ���(�6��<���Y�D4�����Y�I��sq!8S�w��[8z�[��DWsP<������������1�.��Uv%�]vavɇX⤷�h��L(`˳�|��FP�X�o?�~�������mM�:nҗ2򎊄��A�Q��u]"R�n���l$�n�Vʆ�l7��R���KW��fC!%��˫%I�O7�J5M����oز��
z��A_e?��E�6S��/�*T���ه3V(�������e �)��:g'f��V �AFP�j'閉I';�V&��26M�\��{�U�\�k{�$ݛ-/~'
&�Jjܹ��YEp=�dC��*�s^v���d�ܘ�}���"�'�Pc�i���o]�qQR����]�,�MV�&�C������w�H9�ro/���m���^��0��
�v|v��jUՏ�5Yܒ�{�l���$�|A�W�s�u���͙nm ��
��</��(��,߽� �|��7�L��J̥��F;�)4J\E6�Kf
k���p�SJ«����g�	h��ӂ�?�!���|�1-/z[WN-N���6�hD�9ޫˈ�u��G�~�9�j?{�w#(A,q\�d�����Q�A�>G�"Um챈(����bn�����A>�;��h�A_S@�H�!�ٽ��:�n#��I�1pZ��>y�I��b<G��x��I����m�x����cP�-��)�Ըr=G����C���S�19�^<������ρ��G�=��)xAK�~�ӯ�}�J�t��H�����]�l�Բ�K���<�ʾ��&��[�\��2�:�m૳�رb.�]�Ց�X�y�.��wҶ�e!+��\��������[Cu:;*��|�Qe!�^ҽ2v��Ǡu��۶vL�ҽ������kl��u�ˇq�\��������>��>$F�B��@r�%V`�I
1VYm����YE��i�x*-k%:��RA����"�+XJ�b�cKJ-�P�e�l�E����	�[ZԕYy��V�,x��ZJ�n�kUZ� T��{���VI��o�)�����}.�nkRQ��0��}�1@�.�wX��Y ���T�o=m$e4��cH'ă+�NMl��� �sϝ��@:H����9�<�$��������������D�yr4,�U~_8h��ؽ���+kb!��U����=~��Dx#�|$pΎ�^�9��Ė���y���Ǔ�lꌸ�3��B"���#\�>�'��L�#�����Naˣ�:7��$��-Y�׶�H̉��a\:��<� v�H ��t*���OO�׼O�(�^%����̩�QT\��jA���u��� F���#X]��n�����X�S���Yt�)�v�b@�j�i�%�����k���~Ñu���M�̯�8��k׻N��L��FFI�c��:��^y�N��5&A���s�]v��)Bu�t�Ҕr�[p9幂��甩�\�������g���ڸ��8���񰗽�ٳ�#w�#�}�O��ɸ�E�D⭺�(;s��v&�� "Ad&��y(���w���y������l�;��3�<l���^�7lߞ�x
�.(���׏˝&��i�.�;9��zS�@�5&�,^�G�v�'�b"��<G�,I��d�׬� Q��>D �e,���(vˮwTsz�F(���6Ͻ��	�� |��$�u�9�t�p������bw`
TQqH�9n�{��v *(��9ʽP�-��)��.�Y��F����zG��d���c~��>��9�o=�g�:ȜAqFB"��u9Ϝ��;L�AL�jr'O�m���o��#����Xid���t{����$y"**����>DS���m$e4��Bρ"O�Bs�����O�gȅ��I�¹S��v�N�|���}a�v�#�zn�����8�2&wג��̃h"	eU���|HQ;v�
>�@�)�y�G�ǀĂ>��e\R���
��>׵q���������pL��,@��\;b3�ؤE��m�U7K��aH����p�W�>���9�#.2��)�����o��NIN@���ld��<��v��dn�73�^����=�p:s$���{�Ө��ν�؈�\����!�\��v�O��p#��>>'�K���9E�/3��;�X�fq���-}�B>�S=(�}Ý'/pVCu?/q��+k��>|�M��\#�Þ��Y���28G
�/N&D������z6��p#$����_W�����'� ���1C�m�&���0;p>o<��q;c�"��9��bo!\\v}�ngH�<�p�$�Ȁ� n�wX�S�FbU��;�:mT�D�=G�� ���u���h�	�d�d�^����,t����.s�����v�N	 D\���oe8`�2\&��݄}�M��e�Y9%9)q���;s�w�LJ(2θa\������[�t��H�
{��p����ҾC�{�o��}I������߮�5��UH��$�7$�ӿ~���<|(�T��T6�a�
o�\9���9���6���p���$���wC��;�����x�\9��Mp9�������2f��R�}�"Wϭ��;��3
Jk-��x�~�����Œ��'ﾩ��:]��\iS9Z��=)ގ⬎�>�]�:�#�����v"J��[�ӳ��9)�ٛ�m`4nb�B�V�c�˽�.�^�r�os��	�OY�"�vu]f��B�����y�J�Xkg��؆�{�����K��dSf<�����Ee� �U�+5�b�/7WgP�^�)Kw�ۋ{d��y���nV�S-A�#m�_P��H#��T*���KY)Yd���
!(��^�Bƫl�"JJ�U�F�r�*�	K #��GlX���9���6���Zix	`�l�6ԣm��c�٥���3�D��Q��Q�"��Z��]�X�Z�Uʺ�bJ�+�\�(�db�Kt7�0������4�z닦%c����u7l\D�e�֑R
Fl��,,u���"Ɨ$�IA[�n��A$�6�qI����M-�%+��:��1i.�c�̬R�0�rk��,f2�IL-�m��iX�)l�.F�m��v0Y�nb�l3���Ӭ<1᫭����n�]*ؕ�U�ˆ�d�&*R��g5���I�":�����6�-��IÐ?����7�r,������ǻ(
W�ۀ�H�����{�������9C󛆸w�tq����1�{��e����X[.��D&�Sn�Wt�q��D����aҹ��d>	��ۯ����a�6�H���� ��}9۲.�'�H�W�S���i��m���)K�7۝�w��M�n��='۝�����)x;�}Bυ��x�=N�|��-
��^���[��2�ݡz'~̩Ӂ9��ùמ�I�O��A�AK�L��oSv)&��]3������������w&@5ȝ=u�:qNu�tq����Gݕ^�� |�ڈ����M���>8q�������y0�W����3�"�K�)N��>�!��O�(�S��v�ӑ�R��(J{s�m�z��(JL�P�%	C�2��B�Ν;�׃�JN�t�	BP�$x<	��쑻��'�*�'3�7��q�
���L��(J���!*��(r�Rd%	BP�%	T�L�(JMI������(J��B��)9�&�)5&BP�%	UĖ�9����:�2�6E�s�8��m&BP�%	BP�HP�%&I��%	BRs�����s	T��J��o��d�$�J��(J�
���2�!��%	BU!BP��ͳ9��K[�BP�%	BP�HPx��������%	BP�%	T�	F@d��'��	BP�%	T�	BRjL�i�J��(J�(J�Rd%s�<��<��%	BS�\�
��ԙ	I�2��(J�(#!)5&BP�=M��J��J�(J2$ԙ	BPj���n����s	T$�J��2��7۝��ۃ�JC,��B��)7�!(J�	NK�!BP���!(J��C�����B��t߾���ɐ�%	BP�%t3�(��Rd�!(J�D��ׯ0���웚����M8�*� `�<���х��I�8(&�E]���@�f���r��1sQ���j׿���+V���]�xJO	2���L��(J��(J���2��]��6��(Jv��;.�BRq&BP�%��J��(JMA�P�&f	BP�%s߿x�
��ԙ	BPsBRs�{u�9��(J�d�ɐ�%	BP�%	��kBP��I����BQ�	N�%	BRjL��(J��(JD�u9:w�ߢY����ps�v�q&K��%	BP�"�)��.�&{���a�<u*
)$�\����u���}���J�_}��&�E�SI8v0�I�@�ʹa	��>��Q��2�euO�1s�7�xh����O����G��5�q�w�߁�S�0�4NF��u�tv�ؒ��Q������O��=.<$<����K�(dBnNc2�4 �M���� �DE]h(���@r͐|��nͺ8[z�����^Q�{��onc��)������u���	��n��؞���-���m$�Ť˘n�$���ao�Beغ/H�{��M)m��3�!M�ZQ�׷�'k�׳>��Ȅ���T�(8�h�C�bI��0�έ�Ih��~R"˼䰙w�Zi!n6OV��6c�w{�ˤN�*K�qH�����elL,j���N]�ߣ3퐽/��+ҍt��bVPh\���[Br��++mC#��E3v�UL[^?��?�#(3 ��ߟ��{����ʗ7�I�����!�o��j'��K���j�wR�$�{�К��r��a��Cn;��FS�2�%C:���9Ց�
�#�o燀�㗽S�CTBD#"����E�IȔ�7�]/*HJ�[q�/j���W��˳�A�r�u�t��D�`B_y*��`�U~@����3'�+��j�iS2i?�,���Z?#[1�en �r������:Z�r;���P�}
�]M�@T����N�[�A_��L�fveF���\ɯl�(�0����#.1��1�c{��,�R��4C$��'wQw f��M�Y�W�Vf�Vi!���D�"����(�\����6�%�F9�%EWeE����@\S�����b���¤@�b놡�W�t��1̎�u���#�M�]CM��ՆO���}K��?k{�c#M]�-��n�B�����ZAJW�aC"8��0�t(�D*��wpA�/wZp��k��'x,�w��s���oGo���9Ww��X� {����G�Y��s����S�	�[Am��sv�Uջ!%�~�i�풙�MQ[~JB	�݉�A���2��	"�����BO{s �A
}r��J���=�	nC� ���	�T�jF�kT���v�ʭ��]B����9.�QpmY�{>�e�v\�ÿ^7���)P�AFD�߹,V�f H�\-�ش�K�I9I����|;ŋ<�:b�dY�����i�Vp�uщ��J(�����nQ6OF���Ǡ��p������Re� ��,(��>�a�&f)Wt�"���M��a��Co���M$��4�Wc���a~?ơ�H��Gj���V��62�2νD^�{�YuW�H.Q��Y�j�I��FNuآ�Z\F�Nh��)��:�$�7=sx�Eu3.'���DBKۥ��}�B&�`�#�e�;�*U�3o��a]������_$�2(�r����C!�j
p�P\ؤ�U��p4nL��`��/��!�9�E^�����I]�
�uΊe�A�h
K=�%E�r�9���W�+�6�#�[� y̜Y�2�X1)T��DlZ��p��*�H�he:�qL��GR�F�P.���=��u��Ϛ-U�u�^I
w������Е|��I��Νx�"L�Գ$��*9�\�i�95B`�e&ӂ�;}�sr�7�$if����3���Wn�����~���M���ծ�|c\0O�_�ws��(�������� ��1	��C�~ŕ�L˅'Э�HW�w`���N����׵).�����}o�(��V���A,���7�A.*'�̲o2�F�p����0��L�/�⏉8�2���I[9�3���2TwL��oaHp�1��VT O�����/W�roV`������O��?�m�j��"�A��z4>d����{䪀�I wݾ���ӗ���Yqg�t�V�6�h���j�*a�o���H����.����.�ec˹��:D�T�V%��x�F�;<��;L���f��u��]����Ϭo5ئo@G
���g�q�sGa�D^h��SF���%7Gw�B��ݕ�����]�$�����I]D����5'Uׅ��K��j,\� ��`Ls51r F."�\$�*�Q��]E2H��8�H��E��d�x�Il��d�����&ʛ�������M���Kuu�M-�0�Ĭ)p6ڐ;V�-MOG��_�U�4\[F�k�d7&����s`.,�`�<bՖ�1�*n�&�\�L�厔��K�b´6���ڥ؎e�����n�0Ŕ1�h퀵)3V��[�$F)�T��0�!�D�c5huZ��vŔq�s
03��M-�����,���,s�a��i-��%�+v.)s�BƦ&���-�a�a�2�4�Z���L��R"�eh`h:��q�!n�46�გ��+�L̎w�f�sKf�@Q�nH�q6xvT���uҎ�+�����*:kXe0b3�=���l��%���7:�ƺ��&���eeJ��{�@$}����?B���׃�u^�pɆZ�Დk1�s+�`�s;��e�����+�7s���{֣��}���:��	�S�b�ȰBQ��rA3`�aQ��-C��;.���A���v��Cd�SP0a��!0d��$�B��[� I37z��b�W{�AZ!+va�!��6�.�)S:��w�>��}�$�DRAgs�B�3a���~��>ږnJM�ڨ���>?�����c����bb!���݂s'�d��ω�=UM:� �pE�ݝ�	��	��qY ���'h9�Nv]{�Dh������(ki5�mM��v��\���:�7)�3n�(�AL,��l3�|�ق���SI�>���m�K%�rO�/t�Wu�X(���w�L%�U�"S�*p�,�%݂���nF O�p��,���$�C$wv^��-a�e�$`���{%�����ۖ�ZޘpɆZ�Დu� �ݱG�@!.:Y��_Pez�!J=���a^�"�~���{�F��m�ϡ"".-��L3��ʈ`�e8e�j�"�ge�WQ���D��Y�lם=������Zɾ���O2������iϬζ�±x"kg<���AԢ�ճ�����J&�����% �ј�;�}��6)=�y��͸FĹ�9�����ed�'��έ�$��m �.
a4Z���?��p�pŊ͒����G55� j�Hmn`�y�%�׻�B���m��N��(X(�bX/�L|�>w�v���B@�'y,۫�^E�-y�5�ރ�AK��v�����ﾾзߧ��X����NT�Ͼ�/Ѥ��ŝ��d��s@���U�]5�����rP�i��h�.�7N�+�%���~ߦq����Ŷ�0ǤS$�1�K�7�F��A�;JV^e0�3�)�ó�&����v�J�9<{�QXǍt7�&��Ҡf�L8ñI�N��te�޷�����|d�q��4)�J,̼�ݖ�0�ݝ�M��kò\��^�Oh�KY-�C���y�E�<���͒.��������0�5��N>84�'sik�(@�M�f�Q��ޫ*^r���.cdq�il��6۩m��u�ĥ����$׭���J�^z���L�ey� Z�VҖ�|�0T(�|JS�ݒ[h2q_�ט��*]����j��M�ߦd�@u;�n�l�#T�C�|��O��}�g�����tE��0"t]E"F��b��dOM��P�p�Ajռ��KȐD���^5u��9/�"�Cb��:�Y��6��vKB�Ĭ��b�����e9��X<�fb�]sƮsU�5Z�ˌ4Al&Է&m�C��i��� ��33}�~��.��o�<�:lJ�j*'�����S1�B��x�>~Y{���c�W�3^��)��B��n?N�;����E������_�9�v*޼���۸vt�W2"1s�J&��oU�Λh�U\�01ӄ�'�K ���i��fN!���՗t��s���n@'�t��)Ծ[-z�=�mc�㩿`��RyM�����F��ޙ����2�����*� ��=j|�#c���>${�[ׄ��Afd�7����C�ʃ�
�S������S��ݹd���5�E6��Z�Დjɋ�$�D^�!����9�&Cw��<OE��'�5�2��j���3ǇS�(MSv2���Y���6���u�3���.��m�sU(A*�ц+s6ڦ+���k�0��\H�e�Sw�TCCI�q����vU�D�
mK�f�<y:s=	�%/���]�v[����7�:{��;�F�v���ӨW����X}2�|B8�=�=3��X'c�m�]� �|b��L�s	7�E-��*�`	J$�zJ�k�,]�wwy��(n#�}��`H14v}&WΥ�� c7C��󪊈�!z�vDV�v�M*�>7}.uq�H;*X��蓄�XP!�M�i8�0]=���f	7كb:��t��-"}v`V��8�F.�r����Z�m����ffi�BAzj��`��f��Sp��%Asd��/f�-�[�� �V9*�X��(��d
Z�^��pI۾[7w|K|V�n��	ŵ%
Qt^����F���8Ƌz3�k�nJ=�OJ���AwZ�jP����ʰ�����ϊ�ɪ�\�d�X�N�ٹ��CA�a��wzq���r�x���
<0�:���5�jQ�k�-i��{��Wݯ@[�Ҭ��k��h���'aO�����X�����Z�-��޵uG�O�6�o�Il�S��*�[�H#�B
2�l�����2�N�Z6^崐A:�VԦA�)�6�e\��aF2Ѱ�K-,�V�B �,K�e��XDQ,�(��JA�я�W�B��V��j�s#��e�Dk%��Qs0��`�%�Qg׽||��㵌V�mf%t���E ��y�9ܹ#.��j�d�4\e��+t[v	��mXǝ�8D�ˑ�K�S;V��X���f�n��p�Ma��V3%�9�*�71l��,P��hJ����3�(���j3H����o��!M�\�ZT�p:�.��#,u5]��,�Ra�JWQ�JKV�*�R��E���/��\��͚��Û.6V`4#SRb��(l�3�Ȕ�ii��E̥��e*�@�����f��溂��JbٝC)�|��~�Pa���l���Lg["�ߐ=��vw�%Hy=uJ����0��$I�0%�L����MC*!����8��sV�=�,�g(]0�}]��r�����)d�X��5wB�Rmw^� U,�zI[��x���l�ߗ�|26��T������کΛ�3���0:ץ,eWGWڬ��m�y|Iq�Wt���1��n���q*"!�Sf"Q�3�2~y5 ��f#b��ɐ	.H�T���Q�����riͶm3��6c!�Ndc��|b)����(ٽ���i��fIÍt���j����:.h�Ւ���M�鎞��W	���U��&A��zI�B_��䨤�8p��6eM��VⲸ݈���Vʷ+�4ٮ��R\Y��־wߞ�7(�5m�o�)WJ�@�����P����$ڄZ����7q�w����4M,�\l�r�C��y���gVqlzrp�`�1��S[ �g����1W�z"U�Íy�=޿�M��\~���'�d칭},��
��A����[�ܻF�++}��Y��J���:�	�Xcrz����"����>���s��c�Ao&���0�������#h�@UG��Ւ��P&6t�{sՀ�p�`݉��̱�+ç�o��W��WA�y���WNߎ�s�q��l�و���^M��_���#c.��,s�$(��/�էr�i���(�]���{�
���k8�x�M��[U=GpFI;�Yߝo5R��eKP�ۉR�Ɖ����l6.�G�s����J&��Tu���}�b.`��2���!��˿��{TI_VL����@GF�C�� ��������֭!1�9*�.�;;X7fś�WX����M)}��	�����U�/��GqaS���G�v(^��%@A���S5D��	5��t̤���Ge�{g&�����a��&�i��H��ڷ�Ȋ\�HB���(��_�������J=�/��k�u�$��iu���:�W"YyݨU� �q���g.K1*Q���U�C�+3�G8����l��Ɛ��� ˦���v7:�zwJټ�VN�$;�i�(��H:;`"q�׽\ ��I<X�!v46�tϚ:��rV
���A�;[��p��A]<� $o[e����jB�H��JD�o"W�Q;[r�(�$��)cF+%�ETTdF+R �,�`�X��QG�D�F�d�fF�dbZ�b.Ta��`�jB[��q$d�,�HARȹ����?Pa$޺��D$G*��B�;{�,��
��A��7ib�쾪0q��ɲ^c>h��9d$vs���<���0��]��ʀ����f�d������[�w�u���?{�Q�!U뻬������>!�N?7��}#�`<�|�GȢ����*�ˌ%T"X�Τ���I~0^G�#F�ËeP�,ݮ�k3��۵��[�5�,Hpu�p�Ym" �YCGj��M��
E�[A��B�����@�و��~��eg3뫾�ř&�N�1V���d��zb{{$���%UY�w��I.�n��$�l���4�&Rp�%s��[6M�{��˵|�xS�I��.��ّ�!>}��	��\s	�E��:a
�W9���aQ�RH��ls�Ǘ� .�pۊ���cu�|�(����ʛL[mT����峔�ٷwnǳ�4�CA�����J4�W����6��Q�!C`�-9�0�KP[�Pn��TA�c>ܱ�egQ#}˟�{�2<=dI�ݫL �f�Ѓ��̎E�;nZJWE-�)�Ai��M����˺��Yr{�O�ͅR|M���xO���12��S��V�'V_g/9(���J���spXjy�(��bӋ��;��	�1c�a�
E�e-I�7bb�@�T-0�ʑ�0�ʎB���~zej�!�Q�V�vU�
$����E�:��$����&��k�ӌT�R�QF�u6�ve%7R�z�(��P�p�?���}uW��ML��Ub33�n^J�ރ��Z6YՔ�')���j��	/4�U���l�n_������������I�r�8s��X�wHDܼr>RF�o4��M�9j;�c�����ר�~$q�>6p��D�!D��2y�$��������ٮ��7�ly�ܻ�R�"�ҁ�7��f<����p��R��!���J�r�@��<���t�Q�$���/����B�������0��Y&�f�Abh���Ј�K�Y�H�)�b��"��YT�i�j��K�PEI�x�k���G��������H�a�TUP��,PGV��@E��C���=ݱ?FH��a�i�i˗��7a�'�����θo�z'� ���	����b� a�d���na3��@����r��p������P��?qx����N����{��p=����;?��F���۱�h�]&|7�����@�r��|�C9�}.r��h�w웇;���TG���������s�@ayW�"��yPQG����Rb������oQ<h����?4?M�?�������G������Q��~
(������Y$D=�SA�~D&�Mσ���?���7B��njD���`����Y���z���&^s���i�8c�"���c�幏fM��4o��"4u��
(�"�m�:�8���<9�4�OӃBz��q���s�PG�xS�*�a�|�������#�?5�5o���y�A�|D߸��+�A����������=\��뇇�gQ��Y�h@�Jx�?�'�䇗����a�ǐq醇��<�}>�=}�#�w��5�z.�~��|���k�_W��>���<�g�@E!������}C�@�Oӡ���"?ho�{�!��	���*3~���j�us��|�+����p<6�ю��'���A8<t ���z�) ����y�#���� *8��`�<�"{hp���N��vX8�Y�����CJ�Ï�u&`�^@�sc����������=���=������=�(��> �FE���y�2~�������'��{����!���b�`��������[��O�?$}�������o�����=_M��K�T���~_w��_j��8����ź:?�?E� ���?7���Hx>�:<D����C� �O*Β?]�A�5|0>G��௯�����N����������M'#����?�ux������m��>�jZ�lp���G�u|}�>�<��0���{:����n���r��?�/����H��G��<ޞ���"��}�֞i'�x�����p���ۤ=u���Jb	C��"|��=�_���"�(H5 