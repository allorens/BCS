BZh91AY&SY�H�cݕ߀`q���"� ����b+_                                           ` <d      � 
 B(  �D   �  �        ( ��@@3��R��T� ��)J`� �IIBDT�P �"�J%U@�@   � �� � : �(� �0� ��c� ���{�x�@[�$0K!��݀:�Hp��+v8��( $(<t�l����ϥ�^�t%T�0�H��ܼz[ȩ֒�u�O,�D���m+�h��g z  f�*��k@v�� :@ `P  
w��  ��@R�
R�P��� mc� n�q� 8�  5�x p ma���;h<�r=� ��‮ �x���p   	�Ҁ(	�}� �y� ם�U�!�� w�/ w� �y�����G��(��zu��` q���<c�� PA���h�� (�QB�UAG�� ��` 蹀� r�{� �������ϠC>`����� ��y =�O �W� p  @��� |�=���w� ��R�����9t ��z�׽�$. =��O@;�=�ްW�� pP P {�H �@�RT$ (��}� X|�������  �� $u{ ��=�� �f >7�� lÐ ` @o  �p;`���t��`#�u���� 8�W��v<�9 2 �d�   [�   ,T45T
����lx�b@��2 c�=i��q�������u�[� ���r��E  �x   09 q � �pk �@������@� M�@� n�� |      5<��R4�F  C&!��IIUd �  D�2�T�id4� d��F�� �����T��� ��4���S�I)J�A�#L��  �)���)�dM��D�i�hf�&'��}�^}�h���\����m݄�����o��"+���T](*�)� ""�y+�ڠ���b��g���?I���?�x!����������3� T��������r
��"��(	�I!�CD(&�M"�$tH��� )�GD�B��D ���� 4H�h��!�D
h� �P  P4@(h�P�
��D�D.�]pJh��D.�]:$t@�4H���WD'!p��(h�4@ ��]�]�.�D�@�(h��h�� h�4H!8$�a+� � h�4J���D�h��.�$tB�H���D.�CD	� �+�@��C�D����(h�4B M�D	��4J�%��CD!��h�4H!�x%4C8@� M��]�!tJ��#�WDpB��D��D���%t@�$1%t@ �D!��h�4H81CD�� h�4@�%tB M��P�*a h�4B%t@$M��8 �B��+�WD.�D���.� �� h�4B!tJ�D�B���WD�� �(h�4H ���� � h�4H$M&�D��$D	� h�4J&�	B%T8%8 4B�h�� !�PD(��:!	tB
h�D���
��@GD��SD�B�$4J�h��)�@SD��� ](� 4Jh���WD���� 4@���"	�Q1?�x��C������ܽ�q����&-��'E��G5pb�6#g�{���(ƮLf��3��B|�7zowi�rt&�k�4�:pT5յ.\t�ƀ�q���A�4�\����e����~ft�d�lU�����d��	k�QS��gQ�����sV�W:�Ik��H�gHfLB�w7D���t��� ����-�s�,�CRk��lǯ��I�.��@��כJܔ��؊��n�?N�bB�- �{�#F-��;���rr�P4-��ʨ �Y�ۛ�@ܨ2�y^�J�A7��AVY&rz$4�E��Gv�ru�-ĭ�Di;��o&ìQVh(#��Gps�vQ��n�vǇ'Wp+��7��w;DzYKu��({͆F����|��CXX����	��NXX�cҮ�m���i5L�{r��G��gA��M��;Ƨ����'
�`��F��}"�3F��z�;�q,F:wd߹ͤ��b�mխ�p.���n����;����_M�	utg���Z.γ"��t�n�T�Xܙ�X�쑛9�AiU_gJ���9���V��#7-Ƶ
x9vױՖ��N$�μ�ga/���L�L������@P�����F�=�[E�PL�C@�è�&\3�%�Nv��4#�;���5ƍ�F�幃x�kN58��������d�/ۗ�9`�̽��Ή�;u����� r��6�k�����h��4qU-a�������h<�L�������_C~��=�;�$���
˥U���8��-��N5ǣ�4@�V(X���̗�5�n��b�1;Ca"b/+YX0U���vB7sMÛ�rʘ��9ҙ<�`�pp����]�x�_l�&�N��f�!�+@�B�w�.<]Z���:�2jvnn���ڋ3_`��C��M|�1$h���mN���{X���<4mQ���jԳ�8Vwo<<�P\���$G�v����Wq��gv�8u�u5�.�קZ~pͽ�7p�� X���gR�o}���.���{�:;^��7�G��	��V�y^�3��G�6��V�О�@�e�x<��9��r��	�;����I�9��D)�Iv�^�������˱e��v�5B�����t�����R8{A�̂�(*�v��;��5�u�p��9d�m2�#����6j-�]��'	�-��lx��^��vr\���}�S$@LdFs�F8w qA�c$Ȫ�S(�9L}������q�u#X���> ���ѡ�Wc�mPО9�L5�qmmJ�ŋd ��6�0���)�F�'l��1�M�ENửJ�W�)�3�r�ɠE��˰*.�3��W�Lɭn�i�UE3��ັQ��hPs�x�w��3�Zf^3�8�t�ۗp���ܶ�s��F���mB�:ۂ5�:�Q*9�Z.��:�6�PFkl�axi�%�4�[f���k�t�<�!��Z�s�9@ם~{�⺸�ɄG�2W6]��Sy4��K������tݦN]��r�i������ߙփ�G�֠��E�'��u��,����.�P�G����#�o]��2��w�=��+�!��oˍ�CMÚ�M�F�cN�#$�����9'i7R�hݽ�j@�o��3���T���v����s�|_����d&�x�M�	�v�	4w.vӍ�Ls�5K%i��u�~t�q�:a����o7�L�$
�,�suA�˥�\]׸��^u����q�\�:�t]�XǼ�G9��80�sp�F�#�u�Uط�*���av:2ub��Dz�E2�T[�`�����k��ø!�s��m�-Y:�nXW2q)�,�Oal�7@���ێ�������e�u��P�2�'t�8N��Ը�ǐǛʩ��fA�*p6'��fX��"L74�>[�r55���v���O�Ѱ�㱗�I7G]\ti�;�3��w�yj�>?O�΋52�n��lu�u�P��F\��%#���R,銉a�:-�u�3/�T=A�X@͛���Q]�72��ҎG#���s2`����c gg5��n��l����C�,^Nr��h���`'ĩ�����sy5v��C���\&׉�C���6|�<��L	XZg<0`snP�t�8^��4v���!AӀ��9Y�d���9gu14�^���V�LJ�(�jg�˒��7f�v����[W>G^�:�7���8c*aX������b ��Ã驍�9���&����JR�Q:��6X"�ܫ����gRx���-wq��Ǭv��X������7jƲN=u�����4csE�P��R��eO7r3�f���H�6-NQJ��Y�sy����1�廨��Q�km�es�8XUqy:�j��Zӑ�庁��'���Vi]�\1s����P�H��h����e͝>G~��B�on'&��y)��Aր.]�Ɇa*�f�a�&��6C��K����S�K�R9[�P�'
*?MkɈ��y��_gN��|�ѻ��gh�r��aql��p�vt�#T�ܤ�^���8��.���dP�קe�wN�qQ��*]^��e�wi��D����� ����נ��$�Y�p�E��-����Z�f�HQ*�Jtѫ{{� )�;r��S���s��XvӦ�M�i��֞��,����`�Pw�����[�.�u\���` ]��R����DlN��حڇD�B���Ӊrn��9�����7��y�Pk��ģ�i2�v��;6$�B�e�.���8R�sre��4�kZ�>�r6�<��;����/:Zo#�I��EBU�c�Vr��&�|k;����9��.���s�ˢt�W��R N�ئ�׺����yV ��[�ڐcfi��_��M�7�S�f�d�u`�;���E�Z�%M�n���j�U�s�(DȎi�u\��F��nk��G��Gu#ɓ�ғ������C�t��n�:.���w�=���DK�,��2�X�y��kŽٮp�t��y�[�.͇gn�s�Ig)�1�۳�| ��E�+;&��<'~���"��k�Mrd]"�8�Zn�	 ��VUH��n�w�xΘ�˸�+�$^�g�ܛ�Y�Ǭ�к��Ö��ƙ;��]�DMp}�N��ho�����\�Uc�u��}�;�$�d�5��d3��3qk+q��gw�we�۫9��O���� nnmYD�뛎�W&��`ہ�a��k4i�΄��*e�����5����	��qK��(�SGs�dgk�lƐ�a-ͯ[b'�7xUa+e�ذ"��<;���b��X{p�-�9�j{��aKL�w'�i����v❻��E�3���h�n^���Ge����").%c���$Ws�~QT��s�YK�}�ީ�Fw�OY�ʷ��	ٗg'��q��&ժ�M�ΫD,������\2���C����ߥ�wGۺ�T�{9L�\]mR�ڴ�ܵ��#�Z5		�F�R�;�lY�;���la�S���s�p<e/��n@��I$�k��N��"�L}IA��M-�Z�"���k�1��� �;7��)b�%��B�nL�vbK{!{�$p/x�˚ׄ%�\�s�AHtsr�� �E�)غKhh;X3j�p���9�J�w�#.�X%��A�۱/��^lU�m5��jow���+r �^���	ܚ5��'��$c����:��6�]��u`�!ǿ��{��-�k��J`�W9�x!z���z[/i�!N���]�r�Q�r5�ݯ[9��g����2m�7���&���Q-[���][q�;�.8�����<��P3]sP���6�p��/:̖a�&�㹫F�-�ɰ'UY9�dzn�G+�NJ���8�X{�J/u��7L8]g��]Ҧ�Lŷ��r#^�ܺM��4�H����P'O˝�m���v���WL���WwM|�Ϡ��Ͱ�+�Y�Lr��x�@Dö���z�5t5���Y2�۷vw�\xq�볦KS>;7�%����C�F��)Y�ѪQ5�z�T��u�9p�oD7���Uv,�ل����Z�F�'��c����(�%�U9 <zߍHZC,��QѴ��k;���5������NoG�N���VIp�:`�DB�]��h�<�:��
-5cck۽K��z��8�rws0ܦ�ۅ��>V[��Ri�Wiic�Px�ц��V�o�A��킦B!o,�o;Ͱ����͘�B �Zu񳃗F�D��qf�Y�����Aw^�^q�Y�u�v�J(���G�(;p����)4�wik85h�W��;9��]��=0����S�,�����2�)���!�ň3ȗ�q6N�`'�YwGf���A�;��6���ӧ =��j:2����|��^+8��[��OӧAʜEO���Q#��L=�v<1m��ӎҞ�U�RǛ�'. ���bΤ���A��G���Y6#���ӷ.�3p��S,0�/�]w��Χv7�q�ᵓ�������[���vH��: L�o���j�
�c5�	�$4H�W	�Wy� ���y�5�4�}GVlZ�y�*�F�>�T�arj�,lds"�Gf� ��f��p�H�]V6\ -����U��� �#t�i�޸m�gH�6K�)C�1���-˖E�#F$&O�|3�:8�]���x|����;�C�fC�N/Y1���w�c[��NE�:dt�3�q-�9$�f���o��a*u��xr�41,�,�'v�����r�\93x�T���͋ecqӣ���v�y��BO�8�A�ȷ��먒%�̣yb�����9��T[�a \Qi����xa�boR�Vʛes�kq:Mk����Wڣ<1R��G_A�N#�\��7E�A\�SJ>�wbYX,�հV[y��שq�e�3j�i�2v�����Y�P1[�K�]q�H-�a��-�Ԭ=�
}&�C�!u�D����6��oŎY�!{3�S�����d�-\�:��z�y�Xlc�5S�4͏u���M|�7rG*m��i�<aڎ4���x��ga��.�{S`��vڎ��🠯*�sk��2�^8c������Ø^{����r����uޫ6sO#��ac6�7��p�>:��݆��>e2�܇�'Y�mJ��\�� ���(tm����.A�C�uW�؊��(i�pd��5�u.���'���� �=�o(y�l��g��ۛCu��b�����8�@����ќu����u���v�ڞq�ײxYo�"��vJ�\E�4�M�ޣN����̸�<ڴnj��)�cᜓ�z�~�w��j��=tp���1�bΧ��nCR7�Zg��]�2����PZ0�Q8�� ���s�1�VE瀅�^����[M�	��R�&�[yXA��w�weV�����u�� �ɠ <:$M���(�5P���������M��X0�5���sk]뛠����:�`壊�T�n]�7Mp<��T���Z�y��u.K��:n�Ƚ��=�1�{I�T��'��׫Aނ�H���$��@��w�L�Xۘ�s�Km�j`��9��m�n���E#��^Ѱn�z�*&���tH{"�wBh���o+���ގ���f�\�q�m�á�th���4�����=;�D��J��1S�ӶsX�r�.Q�kk���ü8e$�F7x���qטq��ͤa��x���5�#z-��JAsSx�ǖ��;&ӝsZ��aZF!p�Q(A0G`��)1B�L}׼�C@��bg�Y�AOγ�7̺;u�����ۮ�۳�'K�9c+�aYC3R�VO%��z�۲�;9(s���;7'n��&8��d�Ѵg-3�7<6�.�3���}Ŏ� �����r~w[Ů�OPK]�3Y1�<I�g:�lf���v�h����i�`�m�v�e�~��/�f<���B��g5�v��@Q<�h�-Ǥ��Ӌ��(yMH���*�n�x�3g�Q��7Wq|
zSO�U�����KG]ִ^����ߗq"��jº�����*�ܜ��bf�:�P����ws�7���a�'�i�¿]ID�ӳ��S�A��G	��
��r\�R���t��I��]���h���Zr��bN����R(�3rj�gDGM�i��o�:�����Q��X7�H��9ė4�Id��g(we�|f���87�坃Z��2������owor��vt}���Ł��j�����嚙j6�u���j����D9�82M�k��ɥ`] /�ĖJM��]3�>W��R�r!�\�����I���mK��Ԛv��{�Xt��� �g�Ӆnf��7���9\Z�a CN�
D�l�l]8���	��R�
�+���kmP�7M���tM�����ݽ��M�2!��J����D<^�8�.�u<�"0��X����܇c�69�I94b!�Hc�&�-��d,�]�<�CY,�1Q�pͅ5�v3�Bp�N��!ߗǲd��5kշUf}��l�w�@���
�?��'�j��=VpSy�����h9�Nп��?<��D~z�v?� ���	x�#�� ���(P P��T�@P�))�C U� �@��A�D�A�DhJDJr ��
U � F��TrP�E� iU�h 
EJ@($�F�ZW T�T�J )(i@Z@�T�E()JU(�Eh�DJ(
W$� � 2Q�U�D�JhV�ZQrUL��TrP%(�JTiP(C!Q
D�2E\�D�@�S @�U!�L�Qh�@J�F����()C$�����D�D2 ��V�O���O��8�k��Y�q��sS��݅��/�7��U�c�Q:^��,la�RO�AGv#����u��y��Ju�՚�X�,�7Xmf��;^fukx�ZYz�:e�����n:���4���L�5z��u.�����yX���% �]��Aj:li�������ӫ|z�	�W�ݢ��f�O30d��+�qI��;��f�Ͽt�r�x���#�7�Ӕ��Ņ�7�l�U�U?���|���ǿY�o҈(�Q��o ��������; Q-��������������k_g!L�W��^B'1[�`Ď���^Fx��(���5�n{ϻ��wv�k�T�_i���u{hI�<�z��W�����n,��w�l��m�+���ה�p�)���b~���}���y2�e+F�ݦ[��-��M�׏�&7�O�~S%߽<���xx
�|:����br�헵?x&���N�ՌӅ���v�hq����w�-�A>���I���c��4w�����+)Hx���}W�8�'��G��AL��D��j�ˉ���ݽ�#}o�T�
��Og��;�r����A��AXX{p{�l�FYO �o��ǻu�V�f�i�2]�7}0z+�S��O���z��x�xf��n����ׇܵ���GN&s�3�M�e��;������Y�0b��0_���K�����x�+@� �g�w��۝�z�x�ۢL�w����aa��_|�c7��[O�L� �@!y���x��Ɓ������^%��F�;��/OpL��ƨ ��%w��s#��w�yյ��g����o�wg�����q-G�4�a���ui::zq�q)����3s�#�ہlT�Oy5�������=3�s~;fG��yo�?`�g]�5�wd]�|�ܾ�|��|�x��-�$�x`@�*�!��0Ľ���Dp��R����N��]�t�qlsB�zG��f�Hqa�
0!�0`��0`��	0@��0`�`��0`����0`�y xAx�%�*�_CW�G}�=s�27̥�.�������,�`�s�̺�w�&��w,z��祯��&_tW��Q��0��pO=�=h�RP�g���=�q�N'T����i��W�
q�ԃ� Ս����;�;�=�"񉃦�_�^�;��Y>�!ü�ł�ǆ��7�6r�Hu��[�����\C�:���چx���b�`Q�)�w �/�����{��5�uN�'ۼU�oq���8�\�z~�i���+��;g/u8[��᧴;�@�Gk���*�㗵>�X'�u�5���4>ö�$���Z��X�Iw9��T�&O<�L~]l뙳s��u���=%ܽ�7�N0bF��|p�<��,����������7�`�uQKK}8f�Z��{�P;-��g]tl�	N�N��>�11�N�Lr[ Y����+�O9b�ǻz��;ۅ����i���{��y��Ǽ;�پ��x��=�]���I��X7��s�s)!��{G{��J�������}�P}���_n�%��7�Yy�4���௞�D���k{ۇ�=����^k�^u�.Afͣ9{ݾ��dQ{7�v�9RE��yL��.�M��s��*���(�eI����/��{X�.�3V�l���@ٺ{���z{�/�$h9'I��_[�o�|r{��?z�I���������;��ox�7<�O����� \g�N2���
P��0`���0`��F`��0P��0`��08��8p�3�4\V��d�ز��_��Q%�w}�^~��.���o�'N4��	F'��(��gy���n�S�h"��&��d\v��aY�!�5�7���蟕c����Y!!�L;�jE{���������� D�I��`�8N�>��X��ZD\R���u�\� ���=snD��Ԗ60�"Rm����9O��x�u����^���&{�|`ո�r�<�O����y��O��� 	W�ʯn{������M{���Ɇdc�U�F�.��՚�;�.�������Q8FA�	�R�ty�|~]���b�v�
��gЭ]���kמP7r�H5���C�N�y����8u�j��p�H}u�}�������C�d��w^�xI2�����]�[�����v�f�X����Ļm�k�vgf��~]�9l�ya��R�"�	k���J|�m�.aLE�h|\������o�U�����~�}��F���Vf�DU��!�E�h��;s�!ɤ4�
��F��n"~[�S^���~95vl�g��w�$|��u7��sg/l�Cq6=f�q���,�%��j���]��}������ꭽs�_�Q*�0�}���<������t��m�8��{X»TB,�NIPp��wއ���U��[��ڳn���Pҋ~��s����B�{d��A�˂�,@��0`����0`�� ��0`�� ��0`��0`�������ʅ5Oe�̃\�L�"!RE�nH�d�ދ�̫�O�mԷKC��5�������<g&��{�|�c���rf�ָhg!��%�!�X&���c�d;�V�-��̨d��sQ|��{7=��xbѕDG���S�=�8vS5�="�D�uM#�C;N<��/���;.I�×�*�d��.m��q�O�c�v�F`!���}�z�q�9����^�W���~�Ŏ�ܽ��w�O��O.��Ϳ.ڒ�7��yQ���^����s��/����K)���眹�}4š,�<;}�<����ݷ����9:���=��ٮz�h��vN8v��h�B�m=�o'�{l�x��a�4�GaX<������x��+��1��j�X����i��������1�F������{���k^�O�9��;��T �XtOx󧳍V���@{=%�Ŝ����ſn�z�
��{ǳ�w�×��ɦ�~#D����G�"����g���F�){ٳuxk�oi�cV��{�_,�}V������5}5��'�>;��%�<�:װtey��"��@��ki�c"0�����.%��x\��jn)���w�\n>��w��	�Py រ����:w���I��]���{걩��y����p���e�v;��n��X�|���8�I{GK���ݸ��o{u�l���Mʑ��E����N47��i��4�����0X�(`��0`�0`��0`��0`��
0�0`�c ��0�0`��uoV?xu�&o�{qm�n������U6Q��S�d4z5����0�.��^��%� �Bx���ԣ��W��s��y`�3��>�㻟Ω�/$�o3��{ܚ�}�ئD>�ۚ�ɗdْ�!nw7�3����k���?׷��O�(�<�~���±���5<`��x�Gww���[ůY�G����~���{�}s��0N�W�{֗��S�,�g��
d�I�f���az,x��FL��ׅǽ��{qu�7ؼ�w����r$����/�\`�K�	��k�Gx{ݽo��d�5�S��p'�[����H�v=�>x2�Y����cDn�����휘��F{��tDW�Hܺ�ǽ7�tw�e<d��)< �Ȏv}��{�v��U�);��}=�6��������o��-���Ç��� y�\�{$��S��/�kO����vu]�����[���B��
"�7��=�xˇ�C���ȵݗ�}Lge����^*�l�<uwfH.	��t>ow��K�@�Ҝ�j���K95=꯽���9���ĵ����\u�ۃF�p�'����xx�kb�׹/�{��{~�<>�ۛ�p��K[�w޹�ס���[���k����9p�a�2������:]��/%�^,�9�h� X�c^��g9 ���J=�FE:*q�ܞ^�Wx׍�����:V� ��	�=�>;�	�K�`�0*��(����̱���Έf|iYv}���ȃ=�r��m	E�k��CO�{}�[���h�V�1�J�=���K����:��k�'s�Ӽ�n/b�9b,�����'�jì��՞�n�O���ja	w�>���Ю]Oݾ�ڽ(碓=�\2������{_����nj��B�6es׷��&���/�L� �z�;�u��l~:toS���c����:����}�w�щ?w�����ظ�o��|B��=��A#9gX��?��OnEt.��ѐv����|2l�Q��ǀd�'�OF��{:���sy^����G,(<�.kXod)���h��)�>��C�X��D�4g,CH�绞6�@?�n��Iu��a~J�9 ���n�E��j��[���z�ڷ<;��(�u����Cr�����P����Ѹ=h�9�P�s�Up��K�$y��Bd��?G�yx�߼������v�}D������z(yq�{�X%�Bܻ�'y�g�3�ҚΆ�k3˾3�l/�x����yX�fS���NX�����,h�����<�|�y���<7㞽�࢖g�����6	ü���u�Fl����rx< ɜ]}q\� 1wG=��Mݲd �����qN�n<�}��W�?b6�ڒþ �Nb�2�'�I%�� ���[s��L�~5
�uW�yr�w>��u���s��#��"Of���2�vS���7�ɶAww��j��[g���7���ܷ�q�o}A�)"=�C�]:7���4B;���n#���5�DQj��U�x#`�Hu�������2�;ys���'�-�CN��ī�I�NS�����A��Q���b�!?/\�?-�}�d��N'�]d��ós}���6����f��;ک�o��ޚ&�'�`��Q����3W�0A���1�=4�jv^���gN,�Xc�1�۵��P&K�$��%��%���^��K^�j�u��<�q��}��8�9=�����ݛ�����	~>z�Q�Ô'��lf�\�����nt��4���v�W�q�ĘI�Ɇ�G�6H�n�WU���M�9&����ݝoX�$>�_F*-��ŰZ��J7�c�B�l�{�N-l�b���fn��)�D�:����wg��p`Z�n
�D�=
`��w|۶��2��t�]y}3HCY��h��i��<�o`�S��>�����=�LEX�U�lQh�]�8�峼 �i�'�nk�B���_�˓������}=�q �������*4龝���'G���g��0M�Iy�$GF�)��nm$��M�/(�2��f���/�v�F����upB����w���G^|�������o<�8�ێ���M̀{�A��8.,M�k��;1׋�;�Y#D��S��g���m�k�^��{�-����7Ej��{:�+'�x^��HNI��A��1r�x�i^��Sw�L����.xl���;F,co\g����]�|e�.>#����-���v�Fj���ŧCZ��,E��{�g]^��r��:l���MW�ݪ��i�߀�=�t'}�c�<ǌ�
󌅏w�y|��}Ʋ�[�8�l����o���7�?TWD:�>+�ny��]~�鏮B���{��E�\���wM���y�7۹w�n����]�g�t�Z$+�n=w�=ڢ�;�\�v��q���M��C��:��;e����<�gW��}���vһ&�͍bמ�X���3�޿8�>~�����/�g{T7�o��{}}��"�v���ۉ�W�
�HK�4��=/���ro�nҼ:6<� ��Ӗ��79J��ߛ~�/p�g}���<�	<�sR�0�A�M�fN��>�4�H��FB<����=7�z�>=�J��dO&mvM�3wt��d�)�Wf7�ͽ(;oz�5�ѝZ�V���o,�SHN���;�����gi�+�[�v/x��(�/���k^~;3w��E������ƌs��{A����OM@��o.����[�^�񫻅��9�^ȴc<���[����+p�۫x���E�ܞ�����{ڬK+�Y����p�~�G����g=�j8����78��=���`=���.��J��S���k<	��Vq{Q�7�2��2U@^k���I�"oe�;�z5�{����T(����z��6� '�����@ݦ+���`�VO�\䁍���o�咳�g�KS���	=z��Z��������˳w;c?r�^�{{p������J
E��eU�b����L�*�/�R����7X�<�O�����Z1f�����_v�/'�G���;��  �)��x�,\}N��qNݸ����(��^�<���V����pk����{/%��#;�f�}���H�Ϡ�����\�0a靾L�kv,r��|w���ĉ�Q�=��}˳�E*��gv�=��F�Q�( {Ε�/���=Ő4n��p6��x�i���ͭ��X�3�A��Ǟ}��i����Zg�DF���}�b͢�}L����M��AV��_�❒_D��?Gn%!��v��>�M�rx�z���s����>�7�n�Kuo�Nb���:T�N��U���㛫//�
3s¬�\��B�T9��q8%��#��@�~�!y�@<����o��70���b��BNB�L��Le�6^�?+3��XJ������ųy
������\zV>k1m9l�,:��7|��V��{�/��٫wig���e�I���8����0���°���H�|��K���D7^q�x	�Uڷ�lN���/x�s�e�g�l��뱌�o�P[����x��I�{���^���UC���'�uQ/F7\69�ܲm��Y��ar���)�})�eb������V����ׁ�J�r-�b�"����O 5�we�f���`�Cx��^|)7��s��Ӂ38x�V�f��0"�.��J�P��%�ůq�yBγ�����7�����	�4�{�ڄ�.�#�ݻ��=�ך�	�o���ū��W�f���W�����.^��v�	�{��&Wn�<�VXϭw%�5��˾�!����
�|W��gy.zA�w׵�<ʈd���]�{��}�{��^��V�Ƥ��W�<�ű{��;�"�������F�8�<�����k)�`W�\`X����w�LCB���V_u�G�����V�g�Y\���{�����g̫E�X�dİ��9��dm�8�H���n˚�}�c�R��f��YZ��{N_rg�0R������0��j^z#^��}���s����ܛ���9���[��L��$d�%l��_��̧y#���死�Y����cl�\x#ǧj���g�]�� wb3��Ww�[�����xd�8fw�z�=�:Lbb�v��s\s��c׿][��E����� ""��?g��G_���j}W����샀�ھ�?Afh�Ʋ�7/k�d���h�i��f��:���Ʒ>m˫n����Y��x�.
����xqβ����mŰ��n�����Tj��CS�����^���-`t�,g����x+�܆���Ju4�j=rv�熻��I�ٽ��M��"�� ��u`�'<��I��ny��7��p�[��7 p�8��ʢ�x�r�G�k1�Lm����.v�n#6-��\��l)�E��E]��H�kR]��R�sIV]����4kY��9���l;��7l�ͺ��k�Q1��M�:��]s�PL�J���"��q�����7I�U�Ģ��'��lx���=������qӛՙ�Fj&Џ4�M�/i<�)ݝ�et�v��n�Q�ۖuO/Gl���v����=t��_F��Oe��1A�6�K`V�f�c�%��>��u��%"�q�X���B��Xˌ��Ұ7G�/cxjks���-�c�Ҹ�ާ����y6{GvL�z^عϑyq�v�U�:���Q�=�7M�jю�<���cl�3�t;-rZ���><d�x��9wC�� ��G2B��b����Wj�֊T˛����8zi.݋�f��<��Yq�5k +��b��s@��j֌��3.{U�M�Ó	ښ�`L3R�#���tX
¸��P�sU����#�S�!\�؎�eaQ����^t�F6θ����uՒ5#c��͐�ѧ��!��Ǎ��u�͞Ez�瘶{r��@z�&���\Y�4NyV�V��{v��F����k��R[W��8�kvչyœ��f�S<�1�9�*��N���N^E�8V#f덏<8���e��(6�M�]�52��m�����,���M�H�q��Zn���<ü-����we�dG����z�r�zJ�6 }��N7�j���3ەd�M�$�����F�Pt�l	j햶2��V�=��^%�ݞ3��}�:WQY¹�H�w#���v����|>7"�j3�f�v�8n��Ņ�k�a����^���hm!�n)+���h!����5�at��<Xd#dٛ.�1��n޺�7fns��tg+��n5\�t�v���`j$Ŏ��N��:��k\\u��4�ׂ9w����j3�^����6�L�U��iJbU�Qm���Üm����3�=��B赹Đ�䕶kJM)
�x٨��-�d.�ͬ]�R�zd��&0kk�H�Ý\�vt���=S՚;;�sC\��umG#�=���s$a���\,�\��s�h+��bX���"W���,Rh��Bʸc\�j`7-b�7.5y�.5^�toWI��)��u�Wl��m��&��2f:�c�pQ��&�8�s���v㱊t񅛨�v�c���0��]#����hz����@om�r%�H��\�9�8��y��n5'4����͸z�vzi�/�W1]&mC�ݴ0D�u6�++����k,(�tmڶ��a��'�7��km�-��Eod��-���a��xX�y�a�G7j�H�cZ�2E�6k�1��Jl���j:f,[#E��^U� H<�Sf�gsѻ�x���M��/��� �e[p������ùY�/��;œ<F�;��r�w�	�9�%C�nn:�3�<hn:�v;e�<ݷٔ��fe&YM-�6�:dN:�p!�AyD�<���WZ���GT[gJ嗗�8�����ظ���%��[[�S\ekDk[<M�nδfᑡ�gT�M,���C:<#�b�ᱮ�WCL��f��Z�n���'cm ��׭�ts'f�Bs�%	��Sh2�r�`qX`�m�pwCY0Flt<����8���s��b��|��ƻnl�A�\A���jXc(B[��a����.�ԅur�62�Eu��hyƍ�ͣlp����J˖.�Q�R+-�4	����MZA�k�U�M��mXe�Yccb���m&Rn��w3��f���;������ �yq���=��c�n7��KN5�31�IV�Ø␛q�aeu%t-	ts���CL¬�ɡ�ݰ�r�"ʪ;��k����/;7ty{Nn�l���7f�rӸ�wA�����2`��˶ᣣ���FӐ'���Oqg�����	M[�rff���l�6��&�ɲ��s��+����Pa�x��`*sV7�i!�mڜ(�v��o3�7���C��z�gEѯg��l���AO-�ر���ר:C��+����g�q�Y���]avX���KF	�&�[�v yHwcm/C�Ͳ�)�̣tn�tEղ�&͈�����u���<�˽;2Ē�������3���me���=�n4�D)]\yM�.�&��[�A�2�s�73۬CB]�X&�,ek���X�����q�n���C��Q�{�r`Q��8MGI�[�ͷ=�NX���U8�Ꝯ�'!L�v�ڱv�XLi���P6�ǂ�ٮ.X��N���x익�4ss5�,*�Cc�0G7vK;pjI@�:��L�=�*q�5c3t��8g����M��^�v-�(}w��L�[r�+Sоn��.1� V�@��=L�[PMU�Q�;45׹y�݇��D����t!��Ir\��Ҏ����q$�7A��7vx�[��-p�ֹ���ݫ��np�RZY�WcI��M#^�

��y^2U�Nq���s�cb�Y������nx�c�@[4]4Ô%*;�h�h�h����[M(�hp��N��&�OgGiZc#��؜�^��bF5��g��<�'Gq=��Y�:���Fg]����v�!\�qvjϮ���/uC�0���+y:	mtpH�Ώ
m���I���ܖ\�\��v�>ܜl��[�wC��.�y�X��%[��3���%��:O'�L�e�u�)�,=>|����cun�qHn����b�V����r�n]�ֲݎ��M��y��=�WY{���=`E;mE��n��ۍ�75ڪ���AoV�����7/Nl��G%u��%�hKT��T�3&��CC:7G<��X����n:�*�mHfy�)�V^�\J�6��crܼ,íӒɹ۳!���Գv헒�n�kvi�#�a�B��pp��6�p���x��g��n��u�6���ζ��}l�i}�0u�Q�6w�i�Z{�X=��2=�uj;�;+��3�=/�K�E����D��8�6 �j�l]�j�����7��V�ݔpブ=s/y�\a���k���R�#&b�RX�*]c�CK6#��j'�6�.�ws�i�F�{9x��M��K�Q��9����&6�u��Ў3�f�"�W%�	P�HrQ�ҶS�k���+ysXS��z��}�+mn�6�^jjA���i���Q��k=Y����u19�۫Lb���,�
;Bj+��H����ۭ�^`�\�#T9��4%�Z���%H�+�����lW]Mazw!�����D�8z^8�Y����Q̸�sf{�6I�����<�e�8��o<SuBk�$nl��iJ��;7K�n�X&룙wi.x�8�;g�K�P�q��uԊ�u��K�Y[=s!1��Rr�Y���磳80�	�rYw6mj��pV���9̭eq�Gmy�M�k������hNT�[V:WDe-�%����ɇ�;��u����d��L�ݩ��<㶅���ɹV�ۥ:��v��X�ۭi�a��y�K�|R!o�6�m�w=,Z�ooj��]y�v�̚ݬ��g�7J��y{PuF-峋�a��XO��:�1tn��b�q������Vš}�BvS�Q��[�}Dt��3ݻ�B]�;��t��Vϔ��OW,<��Mj��Rs���8,�+\�6�upٞC�㓴�4�3ˮ�I�%�Ǳ�\�N��Y�X�٘�J;'F�O��n�;�p�ѝ��70�qx�X�ˢ�<6;/��ث8�q�n5��=Y�����h��ᱸ��z\�;���A��T�Lq�u��.t���OrTV�Y�Z<�u�^�:R�ާ5����:q����lK��-�|ٽ��Íb�V�s�=�t�n��:�<v5��bXy��rSp�	ö�ʛ��=
��a���i��D-\�N��d�����&�[n@��]R�����]e�Ƀ�����5s��嵋�yi�
'G	j�G�ո�]�P댑gn�h�\S�w��Fn���5ɇd\kTSL厨.Bi��si�3�a���/[GL��j�4[V����$q�N�r/m;�h�z�ٍ��j;M�%q�Ǳf�3r%܂���3]]��;XB&^gA���rhy۫���8�u��������v��s�t�<=v�mqS�Y��� ��9��nɸ���#�x��Fuu�n��(�:�m9�Ĳ������4a��P�m�-qC��G�]�u�L�]V{C�v�n2�a��7(�.��9�&�v�%u��V�n¹��{e[m��N\���]'Fz���t���ݴ��l��nc�Z��!nk��:\�]z����4t�	t;��� C<���Ҍګ˩
�d�BhN��n����Z�K"��v��s�C�z�\�,ܰ�h�l�X��n@�b�l6�ЊͮqG9�	����fpM���z��>�Ք�[&ckh�f��Z"{X��v1@8�Vmd�t�ۡn����!g[χ����QY1���d�gW�=������]WBWZ�m���RI���r��:�հ<�u;��$[�g'U�{v�gS��Zt����{.�m��Nճ�$�ڠ;f四��j�W�,����֗�a-���'�b%���ulӦ�:4,��]���GgAI�PxI3�2<��*��$����g�����S=�2]#ʈ�**���3�"1����?t�/r-�4�s��B�"�lI,m&K�Te.DDT^W��R�a����ǾQ��W��>��\�/#�<�B$�����jSK:غ�E����dUDr�	�x�~=�+�Ԋ\�p�R����*$����7*�r_l��\��V�Uk��R���	����q�"�%_[�0���4�Lӛ�x����񑂏)�P�8��������Qg�E9?1�竦`d��}f�h��ai��If癚Ʌ�½Ȋ��"%��#ҡ/<�L�")ل̈%���*=�2A(�J��R#����2S("PZ	w]Ќ��4D����P��3�,�<H���='WC�R/*z�yE��ʂ��*�<�( ��*Ȫ��'���B�e��^AAШ��Od�S�@���(�0�*b��u�!&�٩s)��%+�H�I�c��vKv�m��^��c/���Y��N��l3�{*&�ƍ�p�NOF�U"`;��F5t�k����[�G'!��{�r�s���GL��[�mF۝��j۪rm��q�`�(O���;�8���^��N�=���a�"k�SRR],�,R��yW������ڞu��s�W'.v&m[A�p�.]�nf��V����M�������[Z�J>ɮ��ې!em�Ga�=v�}�	7n�˵ۚ���1�y��s��=n�Uc-�ɭ!l6���tt���;DQ��pg���qɭ6�K&��ͪ�$�/9g�i�8�.@����!X�t�%�K<S�� Oo/�Zɣ��K�v]�f���Ʀ���d��0����[��}�n���Txܡ6^c<�wu��f9�q��ҽ����K���ly�v#��Z|������a�Z�y]��uq�y6�1b�p=��KθIzvٮ���:��}�R�㠰��y�c�z����[k��Yx�[jx��xۙ���6;dx�8"�6x��U��p�A��1���מy��S��4c=�6:G��R�@��պ'��o	�\�odP�5�:�Y6c��\��*uc!��	���9��rd�GW��<�p�U��LT����*��d}4u$(	k�6�ݔ�;m��*��8�n��1H�U�v��sb�=v�B��T����[�N��d8qmmMV�I���:ՠ�V7WD��q�q=����V���VCs��H��T��o$G�l�ث�k��[݈=��u"�\J١��]R#�/Y��D��$�����4]b��z:�0�'<��QNN�p�4�;�N3b����[��zgo<,7l��'�0���X�k�ᠻ8,X�ێn7nq�H��16݄)�(�^I⋑*mO��ުFۭs���Vٸ�d�����9�{G������{��<8h��6N6f���i�g8�kD�im�c+��6���l��t���%)6����f��Z�g+C���,���[fȣ��enՍ��b����Y�pec9��]l��I��Z!��ۤ�Y؛�e�֮�f��6d��ź,����6g˷S	mY�n�i1�l�T�p�v�a�m6��YU��y��?�Y��Y�'󗿾}H��Ɯ�$�|������Q��&̶���ہ�g'c�`�ֈ,���N�hJ�[S�7eNE���	�=G�
�� �HT٪	>�W���EHܨb��1��N`�����$��!�$���+q�U~�O���G���PHv��18�&L�k����c������T䃬�	
U�IS�.�嶌�Sާ�D6�z���w.�:�[T�x6z~XŐλw��~J7� ����N�� �3HB5T���x	]�\�;�V.G����v^D�3-aq)6�f��M��Ņ�v��:3�IgK���c�'�R̀��H�ځ���r"$B�Pq^%����E&"Y�����=�G���P<)Y{����?3�)���Y��՗Ɇ�ǁ�L�r
h����a�Q��Χ~���!G����ׂ�Y�ഝ.*1p�|Fٷ�_�3����	��M�����3�6L5"	fg,���Y0��-̇|�ZT9��jӵXH+Ub�2��Ap�^C$C`d��;8�u�br�L2m���AЖ2���#o.	9�re��CÜ� �^�e@%�X�ې�3���Z]�x�I��� &�nG�j�1��X3����G��-��JI�Zp�o4ƻT͌j%�K�58� ��75L<�2!t,CmϾ�����2�����1�̧�H%�Hn��i2�F���:خ I��q �ׅN��H��w�񝍈 �̻v��{ʅ�a��Y�<O�6v Ej����,,B3�z����LD�!w(�|��@4�< �"���vd=m3�j/A\3"�ρ�O4��v1�p����܄{,{;P������yٱ>�p��\���\�+bS�x�h�TJ��ւ�{Y"@$;;�@!u)���fr�;��jV���5�5mR.��C�����$^VD�V�T[!�w��e�WC��q$X��b��8A���Ъ6� V��hQ�`�N���"�{��Q!��T:�//��/���i��b"}ڟ5��]c��f�m=I�6ZK�����C�#[���e����Y8�!Sn�`��P(�>��	�s�	ͬK]˻�΂�LA�1ڡr���S5k[�>'�Sq �X5>��wX��5#KmX�Nɕ���D��w��b	%Z�A�ȩǍ[��uF�	�>$�ȀJ����L�LD�:b�(w�<bحxɢ\���	�%�/%�Mv�I*vfKbp�9�Gj}�*�ؠ�o�W��=�)fO�\:�")�R�鯆������y`�5zx��+s��_KAS�{�Mk�C4��"FY�fXL����Q�W0��-��3:&�z�8��m��HГ3m�^U� �֖�m(ݭ���D�_���4f�H� ��[5��-&��@�Лm�ي۴a矼�/�h��38�|��,W�$����c�^b�Le����
$6c��I�ŝ��<E������V>$ُfڝq'��p��Qz+a�T^d�c,�.���gPd��$W:�$�/;���M�CKm�$6���|N������R�g$��.�&we�;�-6��H2� �7:�A��y��Qx��g���`@�dRc��]��0P����ba�5�pXpn��A �y;<I�P#0�	
L�Ϭ��鎊k��1wys����D��揆�8��ݞ�{�H���9Ž��%�S_����$deL�e����A��o"�����0H7hI��؍��#<62:�f�{vNSY�|��zN93�)��2;�lv��љ���0G3ݪ�6��n��P�f�u�-�.7ضQ����{�a�v��e��M�������! �D��Gl�L��Y�\g�5IsWa@���1��S��3!u���UP�Qj��9�ׇu�}W��T:�Sn�qYW��v����
`�R���ьv��d q��3�ܶ�r�}`3b���6��2�
d��WC.�'ĂN���	$�S&I��O��;� �o���p�g[c":�R1L����]ˈv�z �I9Sp �n� ��س[	�������ˋ�	�D���0wI�L�w�'oj ��b�!�7�~�ʼ8�,�H'*n=$��lnt�i$G5,~�9�n���L�����A7{Q �O��`b�f#��� �c��͟,�	`|�0~��� ��ɊM��j^��ߧ��� �X�H[�#��f�v��Q��I;m��Cl�hq�Z�v�z]���ʑ�Vy��>�l����Lp�K;��ݸ@���ۀ �	[q��WWh;n�X���A$�Uu A#l�1�>I��:�Q���|
�u���'4&�x�!�>S�UF¸�g��l���:K�<��;���K#=�{�jo�ߞ^������m�K�f�������'r_n�v�_�	$nu@�	��HWU��-m*��ŰW���p�gp`�9-�� �A�&��Π��F�`�5YQ �ջ A�r��l:fr嘴k4�{ѵ*���m�`7�K�=�F��-	���SC(��N��A�N�A�Aܳ��6Km�E�ۈh�¢����7 �-���8~^K�x ź1�ny��c�.�NY@�^b�S�.�G�p�ŊGg7BY�'�*=^��kw>w���,. �%�7^6�$��`���6CP;�� 8I���F3	,���;�� A��n��3M�Tm$6��N����"gEUV<E���3p9	2r�gR*5����N8�@$�gh'��`��
�P��JIg��zۖ�Un�<ξ{� 	��p�2{�n�&¯�����$,m����D�����gZɝ ���ǉ;S� ��61E� �����5;��$����6�	 �wv��&lf��g�9��0#@��~Ż�vL��X��;{Q��z`�B�l�m&<A���$[���f`�8������5*;	�ٌ��+�4��E'��zn�:�W���#�����R��gZl��D�\��I�ڈ6�;��E]���H'�S�0>$X���p�$��,�.v27`�BV7����	$w;��"�T�ѯF�c%�\k���%Z�����pe��<�<��DA�f�"^�׬�ƶ� �[��H9�QbsK�b�Σ�oj�.�x�I]��D���6mS����Ā[/\c�<�sA�Y�;���o�������ݖ�b4�L����K`��eXB�ud��Q1X�M,~�����9b�jJ���U����בVf��&ƴ$�%^MlQgD�vp���X'��V��H9Zr��50���@�F���Lx�3�"����+��r{V��k[E!�Ғ(hb�MM�#�)4f��F�gϝ�~&m�Ym��4� �
�!��Lu�	�5�ffK���>5qq�,&4��"�;�Π�cl#�xm�y.����I-��`�;4�qi�OY1$J�ф�<k8p���y{�>$��d&��5nK�g���*�� ��i�vCn�b'�;�k����#Q�X��\`w�x�`oU�����)X݉�ϟ`�ۈ9F�6 ᘹA3���l����<X�!��g����Ǖ�a�IS� ӓ�%8?=�FOn��<��Q�I�j(�v���o�L*� :y"7,m� ڇ��o����ww�=�n>��#�:Q��������&��K.GSxG���[�={\v�i{lf���Èn�X�I6�ͧj�^.��3��cv�S�v��-ӳ��F8����=O���ݖ�j���f�\�)����lz��k#�O1s+�	�Z��s��t��Y�9��ŏ\un�wkÍ��J�-n�vƕyr�G�<��i���+���s��� �v��gscCT�*�`��ڎ˃^�
�mk�PŘ&�8չ���cb!f���K4�	R�j�d�n9�M�a�\V�R�a�s>}��D��.aft�	�s[��{���z��Ru�Ώytܰ�э}�@%��L6�h������`�؋� �J��c|�2�����jvH�8owvb!�����C��~��Ԏj/0o��� �?,x I:���+w�zw���6��D��N�a�m��p�'��z�ݝ{ȭ���Aa
m���$n�C��Bכ���L2G%& ���x6^�˓0����<�u/��J� �7g A>#7j0ȣ�I�s3]��_�6u�uH^:^D�R�J,	ں%;>eG��8�\w����N�l�`�ΨP�����'ڐ:�N5�ܽfl�ܛm"�7Sp�:lEtN,x��zp;wŅ���g�:�|r�{�{'��d����!j���s޽�����7�y���y��N+��h��p{�7n<k06f!E�Y	����N��z�g+�]�
4��Gt��n�����ݨ�H"S���Ÿ�5'Z�ǉ�>ʛ��N��aq����w,�:��m���#U�v�\f.\@���� ��}7�"�f��^���;9. ���wtR ���� �K^�B�
��ߩ�1W� �|v�'�X�z4�[Ͼy7e���~M��Ynp^Y�����c��]d�*��%3l�SR�me��~�y��X����:� A �̧	j��;��A�|]��|f����b�`)v� ��Tyv�����fS�O��gn�$$	v�� �]�c�Y[3n$JV�c�tO�gʂH-v�H#�#���m��7����n��s��g�ǽ�ͧ�����{�}{vք�k�y`>�=î���T��_-��^��ԓ�{�N�L豂�5
�ڄ�e�at�yB_s����2�}�HXz\���N!��<�5-��AOt�c���#��{�n�'>�vr�I��׵�tp�<=E�B�Vy�zR�پ�e6���3�E�܁,�r�Z�D׮��w1�ɽ���R:9��:���|K �i��{j���y���4��N�^+<P	��ǳ�=oU��:f���O�ok�;܉�Q�Ks��G�q��pE�"3�$h�O<����^n]Y΃7}�׏������+z{�@�zܰ���0=ޚ�Շ�g�D�������}p�Q(�`mڄ	�%�I��A�����Z��M#4��c����Yw��. �
m�sݔ��� 1��L�V�R�?''%~�+ɅT�߼����}=D}�׌��֧�=��w����x����)��q�ײ��e�?��0c]����vɶ�ZZ��2x?n{�t���\z�]�=��;�vO>�t�o_��(<��ފ��y� � ��^��}�$L��,HyN]�xsNf��\s	�����9�>�;���ݞY|�m8�|;/@�������{/+��	�vwg�|�6)]=|b/��lZ=g* ��������������<g�����Rx�����܈h���tѪf�ql��C�&���d� O��Ͱ�[��z=2�|$=�nІ��{'��=����uEΊ��r��0oy���D�*z�Dy��I4B��ԫ�Y��+sȫ��n`��C��؂��"]Y<��N���}�i�Rc���VXw�;�G�������W<�������E0j����{Qr�]����a.�Ҳ�S�k:u1���3O����	.������	1�$�Ʉ�17݅��v�t�C��q���o���Eu���y�$#՗�
Yaϱ�ө���_t��D��*�e�o�N���c���W��k���/g8]/���w?{t���W�ؗ��t�l�:v*F�G�Lx�����_��ӑ��W�l� ����[o�qK�s�����2z�{���Rfz�XQL�Y��v�I�i״���[�}��0����'�@�t{\&9���Y�b�L�P�c�w��n�k�o!�C�����f��D��nK����UP��J���/f7x{v����Qy��ud����C��az��n�{{m){aPn~L(����%��<!�Qc@��s#�TT]�DTU�~�yʙ�yW=p���9螌^ֶOD,��"�&���Ә�"�Y�K9t<Q�Y��+����:�msȔ,|�~�"90�D�$ �O��،*W���)�1�D
���n�._�k!�-(���/q��S�Faj^�TDW��� ����J�<����AR�j#ϜSGf��{�r'���d&ˇ�=��ބ�R��e�k�����!��7��^���2wdY�xY��`�NE-`k�<�\��N� �\�Z�杄��	rL�$��޻�rR���O�y�����e�gk�Ls � ��|!9��O��NG�{�߄KI�ve�)'>pNM��x$����q���F���:؞�	�y���&�)��k�5��6ːa.A�u�[�p��E�W^��A$ǁ4�y�;��v�emh]�b5>:M���3h��f�%8Xa֎^�}�����ӆ��5��	2:�ZM�n\�%��^��|�'�JC�L|�ΦI��>�@�wS,�N���|��y��+pk�|��r6�z82�yqf�,��cl���N�� 2�;k�Gg���\���=K�0�.8a�9'�{�~lrɐ�d�2�v�A>�>�1�=|�L��!���D��]������L���ܥ'{׮yN�%)L��}��5�<Dx#�A 3����%@���w!�������|�)A�\���\A>�>	N.d��r�:y)Gs�I�V���^��n_D.']��yv�Ja!����u�Л
#�zSx0�7�xG�����RO=13�8���Q;�c0=��햤=��6g�����{���^�ٸ�Xx�h�eY=�ƞ��L��\y�39��+�:�>��Ҕo�w��G�Y��\qq�����������8K��^zӹw��y��lD��u�䔘|���0��}�@s�~�s��? ��c]�r�Z�[`�	tWS�b(3hm��RL�Bh��1Sm�~�ߤ��3vn��JN=o�<������9�uﾵͲ,!20����=hNcr=�����o߇�8��\��F�R�� �<��nM���{�k��q28�#�}2}O�'�O�	����a�I�	𝎎]�����B`u׾��&�Ey
C��Ǆ�^�%<��5���^��lހ� #&���Ŝ���<�\�dNJQ���i�.��F/qI{�-{��5��޺�ֻ�2�%��ߝkr4�x;��$If)� �9L��IQ𹮈��7F�ދ��j�}��$88�9׮�ͷ�<$5j#$20��u��I��a!��NG:���4�?�V�3�L/A�=��Ȁ������q9�纴�D�͙�'s�9o��܇2��2M{�yvNHf{�����w�{:���Bo�}k�M�JR��w�|z����$ׯ<瑣a!��J�+e�x�ˮ5T#^�<M��aw�}_�`��ٺ���珽�~'\�Q�~�jq�������F������;�4bM˄��mx^��'��!n�˴œ�B�:5�k��`ł�[׮�z:����e��&vPkYȄ��n�	6`T����k�n4H@���m��p�Ɂ�9��rj}��:7f�tm��n�csD��c��֚�Z���E�`�����g������C��9��͟��#Î��Hr;!m�qm�^n������Q�wm:�U�jv(b�7��x�����^{q���ņ[S8��M`�b���Ki�U���b��}m����ggf,�<(����}� |��r;�=F��.JRc�]�����{ݾ���s�:����4��2���1��}��@� VN��1r霹g�#>]qQ���3{ c�U��
xX<-�b	�G�(��}�H�梇2��;c^��|���r\��F�D����\�A>�<���-�쓱h��[P�<��:�5�rnRe��$׿~s˲rC2C�O]��\s�����	a$�'"'9�����'�╌&XA�^y�F���Fz�e�Ɋa>� ~ݘ'�0ڨ)-��;��g�e�9�d���u���K�aI��y�{NK!ܙI�h���2��y��4���S�' �|��	�%{Ĉ#�z�[,AfY��7��d�oל�4���:��|�[�f�޻�}!�F#A��唼F���#^���F�a.A�:.�=�Y0O���|6����H\�*ǈVV�c���`�A.-�]v��_i��{v�u]JmLVݿ{������η�����"N�~w�s.�2R�]��<�)Hm��$xO�#���]��푒}��ܐ�R�	�A���|�$209���,hdΝ�i`|@�+��	����G� ��nܠ��H�0�ŷK\řm#V
���gr��������ϯ��N�3�r�p�U��F�j�
e�؉��^�wI�RcbF� H�U�!�2�I����hw&JR�=������A�NHq��^���Y���ux��I	���1f.]0wL��P(�?m�xIG�	 ��d<;+b	�<@�B���9G�MM��b�R��z��4e�2\��Ȃ|$�|���:.�3���#�}�H�](ۼw��;���o��x�d'�ߜ��ǉ����ֻ��Л,��%1����7�q���Y�x�g[��J�, �~u�F��vA�p`̂Q�L|�Y�a^�ݎ�'�@� D�X�մ��I�5	]]�}wǵԞ�r^��|�4;�!�2\g���|�� 0�� 8c�����>�$���j�3w4�`Դ�<��1������ݮz�2��n{Y�2�d�T�`���N�,If]0u�G�|#+c��d�f)�`�z�y��d�)F��^|>֋��
�q�>�+=u�F�r�8�'���i6Òg�m��r�.u�g��=�_Y;9>� #�sl�Q�xy����//1� ����d��8���{�	�!2�Ls��^b[��#�m�IS�q@v��1�D(:�����ӹb�C�ȿ=k��vI�<O&A������Ͻ'��"<��n���)r��s�Q2�[��H��޾,;w��	��L��Xx�X�}�k�]������^�L_A�5��Yꮽ%̉����3�g�3>��6:��d�>�|����5���FGϙ��Na6h�^�x��֮k�S�x��q�5_=<3XjG���{��y��&X�dd�F{�����d��c��~r<A�.tg9���s�wϵ���'�|�I��:���L���/3����ֶ���8A��A�{�~s���������޽ts!쌁�<��ݒ������s	�d�l�޵ߜ���3����߷�/�����RY��u6��P�KMe�/)a���f:G�u)5��#nUWo~����Lf���Ǆ|����dN@d.G����Rd9&'�9�͎�܈�N���+�a�VxQ��4�L�O���#��*e!�b�`rK0r郪����䦝dt;��"���]\	�I$;_�I2�r{�Dי$��,�uy=0'Ӂ�Ƶf^�;�Rw-*BO�6��I8`�5���N�U�ZmngN���ȓ� �oL!/D��%�Ν�l���Fd�?��[sǙ��	lSԩA$���`�I-���[L��2 &,������K��ޕ�{ڃ;�q�3`�9f��f��3�b�Q�g[aNQGZ�ccgY���N�v�,�w+ͯy+�.{�%{�&e'�9�%��`����>���3V�� �F����:P��>^^@V\I�Ix$23"%$���D�C�clm�-� ��
>wc�.�dC�%����KfL���j�\�m�IMÃb�ڳE��{���P]�v	y�K�^��Pȑ��4�^]}2$�:g��K�I�`Ȗ��a�$�`��]3$ ��D�H$��������lw�R�I!q}) ��]]�&Q�'D)!�	Gs�.���7�U�)�$�yݑu3HE�̉I"z�`L�Ipo8�{����`ȱ���&RAuvH�JP�\�{<�)ì���ՇU���A�i�I$��Q"I�Wl���Ix-�5O#�#Q�/+�Ia
���$m��p�ӹb�@U�s ���(%��2��A�U�J$]�������İH���D�E �{�L��������6q�-v�X�����5an����۫��h󞟛^=t�L��UtWL���N.0p��g�=�W�:�xg�vg�K:��m�έfaA:���\�Q�(��Aڽ�OEGGk�:�<�ۖI����v8�A�+^�������UA��&��fB�Ñ6xv��:�J�W4�G�q��;=d]��s�:�I�(GKv��ٜ�2��2�F�v���5�溹ᳬŒ�fѣ!�]hʝ�\�͹�v;5��fv ��U϶ɪ��mNֵu�&v���6�Į3�4��.I	�+�2�H����m4�
�H;q]nZ_g�~�х.싺g]�aėI@f��`L�N�<���=:�5�[n��bx$�Vt���(>�6`]��y��+�����_N���+��z�b��@$��dI2�-�4�M���	�rt�4h���kIr�T0X�L�0��h��% �	gcɉ	/%Y�g�DI˾����@���dH�W�K�������Y��Ⱥ����t���mXZ�w�ql�	{:��I.�?tY��#>�n�n��Yy1��C�ΐ�ǩ�P 8h�y�{|�)êj�O��!JI%��b][9J�omcm��FߙdG@�	 �
�b�p
�!���Ғ��?c��;��Z[�f�l5�3]�x��p�n�S�N1����\�[\ѻ}�ԝ��GgM�}��M�r$JA$����T�$�#!���%;i��nvn��M$��D��%�`dvE�3��-�ע�>ګcT�j����ޭ�̯H�~܈�7D��2�,��yb�:�׺z�����Ӟ\�n�HZGP����nk�X{�R6�a3C3�n���(C���)��K{�L�I ����Ԩ$��E�X����	��ʖ������3̑EV���J���'�C$��N 6�!�x9���ߒAvlI��Mf���R\����&�q�"�=�����&�y���%�:�(�H�v@�5�y����$wE��u��<���vE�ݨ�n�e$��l	�7=9�W�\�A;�bԆo2^���D�}��%C��.�؞�4C�]�rd�e��8m����]�>[�I��V�]���	�]���w�Ӷ��.�Nsr[��|Ғ�,�m�d��3x0K�]�"HV���o2��t(��z}>�(����eHI<�6A���ˇt�B�˞�D�@%w�Y�P/=C�<�I!Q�Ҥ%A���糪	D�l�iz1�jS�Q�HX��ÁE1wd��:���Q��	 ��l	R��IEgX8����Z%���	{53��� ���%̈́#�~��K���g��>�K9���׎�WWK��%k^>��qP�4�-�8%�r1����ū�
�����%��`W���z���^s���O.�:�$�^�G�̉A%u�"e"W��D�M�۰wce�5/$�9�T���i*Y�c;3$¢�_t��"I�י�S�.n*��T��ݴ��ǩRI ���@�
($���$̫���k{�$'c��.��MH:�JK�'Y+Yz�;�м�N�k{m��h�[in����y�y�L�������K_6�)$�K{�L��;�a��0*m�����ҥ%���	����oLF��˳'U�UE\ɕ�7�>�N�̘��GRI!u�"d�I����X�O����v#��^��#V���tq��g.�5
�=̉�JJ��$�(%�F�LoGtt��tF|�X�� H*E��T��pӣAI2wd���L��k�n���l4�3g$K��	��A*��L��{މ)�A�m�TV��K�^�8��O�k^iV�!�L��坳0����{��Si-�����IX����}ⵣ�{�,�\�-�u������E������x��6;��� �f�L�OuM�9.��g���%ׯr9���Gt���OO��Aۓ���8�Kn�D�K�$��D�&RO}�&BN3�B��@�('<坙ӂ�ӊ���Q<���ٷ]!n,�mQ���9��+ʲ|��L�����͑>��H%��3�)$^}�>2��=��W=8�g]V���©�$X;d4I�K6���0,�wgdj�\W<�I%��)�3l�n�<��H�Hn�I�H���g� �v��^��B�wj���R�;&#B!���Դ��Or��D>��K�bY*QZ�t�����AwdQ�%�|�2����d��wN�(�z�L���>7c�8��W��T�J&d)A$H=nD�"R�����(k������AU��Iľ���ݓ�u>�'η��H���΁}v���I.w�^�H��bL�4�/N�H�)�`=�褤]#R}�b`�=���K�K�K���!����,���νg��檔�^��{��*���7�}�7r$5����Z�G�Т���	��;���m{K|2������+ˎMﭚg��'{=e��y��A�aՉSRz�Ḗx���b����7����(g��zeY�����C�e��Y&ɉX�pSc�ޣ����<��W��+�t��o�����`�u�|{\�t��P��y��Vf��y\��^�������{���`bx��(���Y�\�}pz����sq"+ݑ���-�}Go�v=�_}ێ�@|�3;t����I��{&�:{��R�7y���|���������R"\�mjz\��q��ǻٿ�>G ��\�ɾ���|ԹT����
o�������}�)�Yj^�L��q)/��ޡg,d7�kx\���iط]�ZO��^�q���;���N���Ydw4����A�bQ���I^�<���`�����}����I;�=ٽ���,��}��/i7�x�g��_��U'�wd��Y�^L�*q�G�Ѧˁ���w}���|���vY;zk�f禠=4v,y��gyU�E����{���!��,@q�q8{��Oz��T�}F��;~zcHm�G��c��{���n�7�zt���x�������\rTt&�w"y==����B�W}�;}��^���;����}�����}8���l�{��nt����R��b*�6���iٲ����q��a�Ǜ���(�đZ�~[�(���P�zZ��c�^��wӁ��l��N $!@�m��1Z�!�L���EKl'���	��|���<��x�R��H�����yG��:��E�5~K�U����ޜ��zL��J�����)���~s�V���9tsq����x��n L�o,>��d��6�in�'��#Yơ<��yJ�D*�2���JW3/<���ϲ�4�}�������S�Z?����W)���{+��$��4/y�dh��E��u"��Ǐ�ᷣ��a�Vd��za�QW����Nd�D�
��������z�O�E�{H����&Q�fyC9%��i�hWPI�:����q�O��޲�B��&�QzM��dVeS�(me]Hќ�����G���XDG��!��\/�������Wj��W�xTw�2g��TTE�H�w8*Iz#&̢"�HIy�Ҩ��Zϵ��.�g�Pf^<ʞ���Wױrk��m"��򁪧�u
����EPDO5]䓅��QsqY�MK�4	��;}�*�R�η���;C�ĉ-7I F�`F�i���Q�e��3X��g���-��	�rJ ��x�gn^�vx֡�q�K�����kk��5���v���,����j#��tNY�1���bڡp]%����dp�g�ͅR�n+���7S�.]�Y�ŢK�˞��pJR���Gt���y�/6+�д�\�ьn��:�ucp�7��U�rq����x2�{
�8x�|�����Cܻ�;��.����3vϵ���!�k��pT�����Ѽ����.�`�yͧuθ��ܽ{o�.6��N�l��y�dvn�^�l�!��hq��]��'o��,SGc,��3)�#ͮ�12�2Gr��oY�GMI:18�<�k���B��;w6�ٶ�\��3�����Z12N��&<Jg����c�I�ĕ���*����{��Ӻ79`�9׎�1�a��.5�l�^;w���l�=*�vI�Y Y.��]�-� Kն��7c��A�(M�L�@���i��@ a�
�x�88:xx�f�j%���V�h�7�R4�b�Vj���r���m�e�lەY����q�TY���|qНv��,أp�MV��	U�`��(�r]�nxK�{=�:+l�Ç��N�Xԗ����D�D����p/[�*;]���H@��g������1(طK�r�����"��ҹΞ�ݸ9���������E}ܦ�^���n��5�c�5�-q>���p�[h.�d�:�\i�� �c�]�;ceiիMWr��F�mEm��,�'�����op�cf�3qڋ����uլ�Ac)��k���utOb��n�%�K���	���af'������X͋e��M(�lx�ۛ�z�����p�����S--ѻ5���T����y��#�J�*v���g��[E�]�i�`���[@��Pl�۞ͅ�R
]�`Z�CI�~|�#m
�J��|��`~�8�Ys���z�ၨ�u[�,�u��n�e�a��A�q�v�;����Zj�6s�6Pd�C��Í�RoQ����������T-,ô���q�xd]pr��@�GG��S&���u����i۸��79���5�s�&^m5�d�6�:m�$AeЈ��.���B�'��qg��vm#h�I��Φ%u�k���\�]f	�6����;)��4�k��׎�-��.��\�hҚ�������I���g��+�ڐ�JI�5�}L̒%���>J�͚���*���~��BI�r$�	!�R�b���̙��L՝"e ���m�j�fi�$4��`�;^I$�@�_H�E ��Z�Gqˀ���⃣n��"`�ܚ�FM3̤�D�n��I"^�`wv3�]�k�Mz3zfę�D���%)Xg2LF"�	3�jI��zoF�j1�"s&^$%�A$#�dI$ϖ��&�U��f�6��Q&B)�����;�jI�.D�)��n��n�̌M����6쀕Dc���AGfșE$����O�s��Τy�Vm2��`A�7L��k�l���eZu���j�j��.<��F�U6��|��=�m��w��ǯ]�<�I�R���H�V��)ĭ�K&��N�q�6r$�I"B@(��)?T�8�]�y�y����SuHiA.�ۼ�d��k�;�x_�ˢ����f�����]��m��Wq
:�?hkuΛ�����/m)����}�wk�{c	�U��ڝ��{�%䗤NvP�I���J	�S��of�N��]��&��`jY�CLɜҥu�"D�'9����J�kfx��Үb�fl99�A$n��O��Hw��@��e�f!�݉��q<�4�*c#�ޫ��	�#���DSi!��jN��{������,-?�Jz2D�A�0�d���b�$Ω�$��rPI�{^$$��sB�ڒ���"R�	 ��iH��(��	'z�Ӣ[uU�^��Yف+-�����4*㎘sA�k�w�۔e�c1�7�C��4,�N��˂�˅pM�r'җ�A-���ҀR��H>oD�JՋ~Z�RedjjΑ2�	%�1�e K��C33��;�KoSŋ�d�����Lc����Iv��I�;����k|��if���O�L��:,�0o3�Іn�ؠd��e�Ĥ�D׀�&Gf���&�+S=�۹f����N��z��C�clͼq�򞹢�K(�r��W<��j���������ϸa�s�Y�3=�z:JD�w9"D��M��&BH0\MK"�|��33�T�t��//�����W�ڒ�I�j$���$��L��I(���3������@��]-Q)�����+�j��$IFc����Y�'n&��u��!�"I��A��%�$����"W��x�Z\ŋ��/ B;�cF��7[^��[]$E��<��1㹱���+n�|���0C<��)�srO{Q>2�H$ڳb^�3$��c�D��^kS���l���%	0~l�i	.�xa䝋�r��,U�@�J@$��p�%�4n�DE!x�c���&T��Q$�'G]�a��ŉI�?$33;���N�B%��fRH����H$|w���\j7�R��v�32E�6b|�I}"}){t�,gb��`�g��B3ӑz��]m���r�I$�D��S�fHFwHq(�IoWL�Z���r&����E�1�U�.��`g�2�g�е�������-��h�RX��:����Rg��y�B���8����vXMQI�����$��L��3!q5L���Y��PU]�|Iϧb|dA�U�w��阔�7��0jk�%W�ޜ�"WF�3�w0���ZB2nu��@z��9�{b l7F
����<�c;�����m�;��;1,�˳�5��{ڙ�I)��%�CzzD�H����03\�ى$Azw�D�B�b�!�b�$��)��t���A-k��Z��=E��I����3�AwOJ�%�<��Ebf�VѐL��г�ٓ9gI�*�n�B~��2�I���D�$���g=�D {bv$$B%5�"e�t�	���S�	b̝���'TG<�FJ��a�.A*����3 �^T�!$���[PX�y�7���u:Gg��) �ȭwd���y��������C��L���.����HN�H�JI$d�$��`��[:�36��&۝3��u���5nӻUV�Gˡ�h�vZJ���=9�_~�Iv�kj�M����ވ"�6T��r��n
D��3?���x� ���>~�o����l�m�R�Bˉ�֋��k1�ng:�K�N@ͻl��7��ڴ���Ϩw�lPi��OXz�q��u�(��� �B]j��u���{�-���hNg���ܤ˷���l+��.u�������w,E�m��K���k�š1�^��ׇCa��&�����ύvΖ9���{I­4�V6gb��Wx;G=��E�X�>^���rz֮������Ⱥ�L��쮒@�d�0;�`�r>)�3���Wd�6D�و�IB�3�K�Ib�Ku��M2&Q%yWOH�Kv�5�f%��vwF���Ꙅ�om�*I��:N΋����HvOH�X��?t���3�{�nT(���hB�S3�]$��X�옳)Xo#��@��	F���цE�I$�"QA,/�L��N9fgN�;�Ri�W!�$���`�	TOD�!��$��gKJI$���)�9;�=���H�^@�J@@q1��̘����\�.��,I���t��&H�]��i'^�hN�%Pݒ��Fk��ԓ5�߮{�u>���#]e�-�a�/; �#���z�(ڈ݉wM�����{��{E�\�e��ς]S� �q�l1'���@�	L��m��l`�L��RK�%�%cX�	���2v�maf�H�H%Y� ��!��TY�k3N]f��`�_<MkjD�V�ߑ����o��sf���k8�Lf���l�0�����x���廷>�}XjϠ�
F b@�� ����Q^I%n���JI$���%.4���s4t���K��5�f%���vF����bNy)��)�K3֣��WC,�d�I{��e�$J
k�D�|�t3��$3�K���X��˂�����3���ڪ�{1T�$�dI3�fo.��U�Zb�Q�$Cv�JH0y80��Y;��΍��ӷ"})/$U��&Dv��c�Z���j�be$���H�N���dA���>vi�
�Ƀ�,��;3B���,�i�!k��k��st6�Ԥ]�W[��������1wgb�9�c�D��3`L���HoWH�	e�])�j�h�|�!$Jw2D���;�wp�y����T�O��y'e��&[���ڢ�/�^���3�ŒI���5j��D���.)�W$�c2���!�'jT��dL���I-yؓ+� �t�u�*^^O?<☩����z���s+;��񃽇�t� :D��{��8^]�fu��/��kO�{<�X��΋m����߷ǏG[���
D	�ʂD�ב�+���^Jo:D�$����#һp[XwѧwPդIJ����w���ߧĜ'�`O�/$�]s����͓�Н��pf���]#�2K�vD�P�Zd̆y�tS;J%�&=`�Iy-~m�euuf�n���lI(�� S3y$��H�PI~~�>K"`ކ���bԃ32���ȗ�ѝ�i��S�r�ۊ(�;(<��8�4��f�/���`4;wt���e\��`f�I�vHI�>�J��ki�u��m�S�r'Ҋ�IgNșPN�$�A�ӱt��$6:�'� �dd�'�z�^��D���!$(3H��$�I��$�K5�~�ѢR �U�G˻�p�Ϟ�vc����K5�@K�`�M���K�� ���Fג^Iyv�H�aW�/d�D�^I�(3Iy8Iڕy]gHlQ�;'|�I�:$�>I$�FdI���IN�H�ӊ���kʲ7���1��r�C��a��C�����]]�ww۷�`�v�	h����&�զW��;X�e�����]���]f�F�����A>(D D"Ċ���|<Ï���&ݤ$g�1�;�$ɜ��7v���>_`�%�|�%i�:Z��`�i!y�&I�$��̉2��D#=}"eL���1���6�|���}fs6�4����04�n�Xݗ�kڅ�3K9���`��r�]���涳��dn��q�84�Ἐ�}׉�H$Jv�D�IiYj�x~{*�aH�Z�y��=�&@IY̑<wt��ػM�r$J%�*��ׅ0�f6�E��RU�RI%=}"D��L�����r���8�hY��wN��s2G[̄�&o:��%)A��F�Gc��,��K4$N�c����H)��%;�c����8^g�>=-���9̬��� ��S�2�A%;�"g� �]�<���^ҩ1���U=q&@I8��eb9	;R�u�"})$�Y�;-*�l�[��>��AHdI�݁>�a3(yߔ�S���ٜ�Y�F��l��g���R�^m�F�����f[�|5`=�Jο2�t�p���Q*
d����)�$��UC�,4���܅7o��T�ކ���NR+fbD�H@�|=�J�@�D�)����㵭��XR�n�a�$ι ��M�����jF�CD�W8�;�V뭷JQvU�f�W85n����gj]b�8��-�ź2����k��,a���*���Spe�����Iٸ�����l�ew�t� g���']Zu��n"z����N��G��n.N*����u�$#��s�y`wk��ٸ8쥗�:u��ډ�Wx67R�J;��ƦĘ���֚n�n.9A����`��f��3�wF��ə3�vF���8�)$���l	��%w<��P�y����*#)L�D�I��t	���a��1c�0tS;R�����ZR��G�� ����w�x��(���$�	%���ex���N���i�41���H����394*�n��"Q)*析҂H��r�7����H�RH��@�E$��y�"Rh:0�r�9t��c3�������e��)��D�% I*�RL����M�i'L�I'��'�D]�c�����^g�>1����d��kĥ�W�n%
�0�d��dI$�Y�<�O�K����^Q�(x��#��%�Y��m�A�X���y7<��Ԛmv3�ջ<�K����m��'�s]%����'u�e���o3�D�J���.�[>D�
UW H(���x�spb��̙�9wdj�_K��D;�3lr<NQd�#����mh����}�ۭ���8� x�=.��F���.헂�x_b�=1���Ș�LY娛.|<�"Dbbb������^��|7�������	����ϒ&+�w�
H�`�������:E3��.��PD��K_9�BI"e�z-h�r�A$=m��Tɟ���@IUX!��wt������f�?��u6j�I?a>����0=�%憾�2�&d�zdL&��W$�]/r�JA��ᄵ˧�����]/$L�l	��閦6���sDw��J��ϒI -۲ZBI$��>��z����b�]S�.X%2.�>G�\�qs��װn��x-��[�i��5��r�����Yû�����%6ӫ�>N�d-�c!$��=�"d.Hhv�:�i�� ���H�PH�v솟$���RC0�\�E;J�u�"})$�����Sl��0=K�햔�K�z�`H�����Y�"`��C�ܨ3���vff,�ݑ�U���C�A)��)���y���MͩH��u��J����	^l��
d�L�'}�!��ג��������2?�}��;s�ZW}�|�ud�~��/z� �c�;�R��y)�-�?Jg?	����Z�e���y��n���a�j�	�ݹ2LgD������`���j�����æ��|�ܗ�{�Ȅ$-��wc>�ss�Ypx�禾�̝Wǉ�˻e췑��N9���C�Qݱ\y��i��A�P�*��m�מ��D����;<=��{�{�
$�}�4oy����V�h��G�`P�� �3�LF@�̫7�~bPzg�Ac�����'���ؕ��w�F��v\'777.�q� ;����������{9#���dP}�h!�C��w��}��Liqh��n+�,M<��Xq�w7R/���/���!��h̀}�H@�ƈ}��l�^^>�������uczy�/�LI��
=��w�'�'���vo���ӻz#���>������I)����f�L���K~���g�:s��ek�f鎋���������ע] Sa���U��9Gv���Όl���[.?5��#�����a~8�;�Պ ���wBj��pȱj�`��W^����U���sf|>
��%_��=������x����X�J�{� ^��{��3bo7��wS�ǎ^�}�92EAw�=��=�ٽӹ��w��A���?E?nk�6U��uy����o���{Q~��^����3z�ݝ��؟@�0�z��lq�Rp��#�CĄ�"̟9DJ�
��>������߿���_��S��(����((1J�'?�2dU��.� rOg��4�}�E�AT�B^9�a��"����(g�@�J�*�NT��lه�M�j��*��gB�"!��EL��B���Q�'�E�oc<�DO��hѣg��1$I���.j���j��dEx��y�J$��DI�>��=~#�>>?y<Q�F)�D�/(���ĕ��ǵ�$���y�Ԣ�Bw�vʧ���_Rd$EAyAE�~{3�6	yx��a�%ȯ�\�*/*�Bj!]*�\���1�/��-���I<N�P�QD44U<M�U�qT��څ�|��ǝ��}t�zʓfh�^��]�QO'�#�h�]E���I�����O�\^eS��d��?$���r'5�<���ly�]�(��}�hʊm
OF�Vg�'m�&}O��x"�,uq�S�@�D(!@*���翆f�u�KO�!���$H���I�����
B]-6�^yO�3!�u�$��Z܉r�H%���T�$K��W����̞H"�`$���ۦ���Y`�E�ӳ94*�uT�2���%��R�='���-�^�y�iff	 ���L��Ao?J�O,e�˴o	�%�@��.���6t��{;���<n�Nd�Dvvc�M�qA��UM��;>�B�q�2�Ӽ��׳/�T��@$�I��~�3�0�g���΅�:�R�A%�5�"��cl����^g�����CI��ʦy��1$�]�$�	(�R�`�w]�Er�1r׌MbɎ"�)�D�yz�:D�A"w�`A2���vͮ���3��l	 ���ϒK��@�Kٸ-5�r���POk�n��F�^���K{��I'�+�$I2C���޷%#|�G��6��b8W�p<z�y=���:��	��z��Ϸr��๟xG�Y� ���Re�S:fq�&e����Ă�
@��P"R%"H�J�^�><\��Nn�LX�E��Vy(쨐���K]g��c_p0���ز�I�[="d$�Iu�H�B���zZ|�sE]i~��%?-��o�x�� �.%@����+uد=�F^��=�M�\T�u�l�Y����o�~șH$O\tH|�H$�ۺX���;z'+�\��$ϕ�t�2���*3�N&5KaWL�Ѡ���]ef��u;ۑ��X���	��+]�'�!*2��9�d�֧����^:�1�p���3�����[�>�H%�y.��c6�H�|N��;2d�I����.�7���BI������Px���	c�Ād�H67t�JA$wd�l��y-�'h/��_�$ủ��vv�&LY˻#wk"[&C$I(��)���V�<��h�Y��T]H�@��MW�&|�	/(��vc��n☈Hd�u���h�Ƿ��Ǎ�+^��K�V�{����=��og�<�;�dg�4jFe�S���ECS�`�ٚe�Y��'�Z5�3��| A��$D���V���(��>5���l[��Y����ο1Z�y*�<3��]�vI�*#=�`��'��{]�(}�Gݽ`��֧ >J5�Oj8�ܦR3s�L��qu\/����;���mc�xZm���hֻt�皌�ң�h��H]Y�b�`j|�Jɽ�m�F�����3
�H#Ի+�ea%��!Ǒ�vvU�rk6w69بN���I;1j�k2i[���pS���8�\�+�Z��}����cc�]�é�۷����i/�%�5�����ο�Q6L���od�'��v���a4k��ͼ�>�RM��RB���Cp���p�Uy?UH�)�HsN���m��($�M��B\3 ��$O�PLʶ��D,�1����ɤ���仇d�HQ�o2I�<g�$��㕏����˺��!$��e"R��"R�8N��;�R]S�v(n;%�P�31$�f�Ĥ�I/(��)$�[�����%e�d�\�e-�0'S�f!$�
|���A&BWѱ �*[�E��J��tO���J;�D�+�%�"D�OiGT��ZM;��̨8(�b����x�@x��u]�/���#�����\��쮻jշ*�Y�6�ɓr���rȝy��I(��O�3�2��Lw2��lI$�
3�D�pp��6 ��wv��%��$������{�����/1/3�9Vj�W�wT_&$�*v=۾~����'�xm�X|W�l\�<����z���Bs俬���M�c��b�@9����-��dcy��aKc{���m~�78��� $@�D�%(@�@@!HY�}o\�3R^I{�{�$�E���(���o=Ftt�<
k�:B����K���P��3�)$�羁�X�:H��D㻽�"R��>��$�L������j4INK�vLf�~�y�zss{L�uB%���Af[�H�t���u�%�L���$�Gך�C<��9{����	�<V��N�3����TN��h2�I&�׉!�o4��u���u܉&|��轑>�P	 ٽex,�u��X()0wZч����c��3���� �us-2@�q��׷@ȣ���N�Y;R;5p;җ�I\nę%fg~�|nT���͉����e�6rD�C;,���30w��\6��e$����{��~�u���/$��U��&C@wA�2���I&R�%u�[�3�$L�Cnv`d�FXC`:wRҔnTO��䵃1��I$h�-�P#�*�oυc�M
���T��oy'�	{tk=���[{�w����/�^�D}NG.�H���~T�F٢�.#Y�/9�7캖��G������U"@H�@J�bAB�bV�zߞ��bA#y;G�M��I������.�Y��E�&+�w5=j��Gǯn$A$��ȓ)/%AO7@g,4�g�	�.N��ޑ>��H�0IN�r�|��̤�I��Ao]���De�%�j^	yy��$�K� �o�H�;�������]��}�~鉍�]���Ç��;vP{7�>Tu����h&7Mʃ�U�����=���L���^w�F�-^	/$ٚ�L�$���&R�poh1���="`K[��v$�IpN��ҙ�8b���J�ޑ"Q6�b�<��X2�A&��>H��D��Y���,�-������}�S`L����#Tm㞄� d�H%=C	�7�H���t(�v��2�p��I�2$���H�"@��4�:v�vN�ZR췩n�[<�9BW�$�X�!%�	Gf@�	 Attq�ȗ�S��m�z�E��O�Wy�{��Z<7�|b��8|�8��hQm�&7U��k��Ў�	<cV�@fp�O��$��|�z/�{�?}�|��h �"D
�P�E&TH�L��g�]��-[N�TY9.�ɒ�U��5"��U?HR���2n}k�%U[��$���vȂd$��:8ϥl�4՜6*"�|$���n�l[f���b��G%��]�v-E&dLj�Ʒ-/>|�S����Ư�]���ϑX�J/6�I%�����%(�*�y�OF�һ��L�����3�yӎ�çwpw䭤�����H�qŶ�Ok^��t�JIz;�D�IzC&]<�fl2`�:��Pg^%1�~{�<Vs٫����]���A>7[�$J^I%я��)$�m���l����0�)}$�K�;2D�T��e�OG%����f���-�Q6�<��XMq��9{�$�(�]�`��f|�-�k�M�M3�+�G{q#�yӘ����3b족-�z0L��>�D�K�z��[e%鍹)���x� J)%��d$�Om���Jgm��])	_&��
ޙ%X	��$@��j���˷/���)l@��^�w�G�z�{���4y�r�MY*>��v�F<pgp\q���D�ФJ� D �(�B	�NHB@�I.�}_�kcL�]Xڷe˄�]����0k��ny���Ps�uuCu��Z�ئf�1��0��-ى��ĺcR�WF�v�)�vAS��\�j�����=�(�0�:�h�GXˌ�N��X�K�u�y��v��.ۗ	�{,Đ�k�N�2�ѻ*�"���=v�s�Q��,��£2�nwUy���c��K�ء����1�Lt�k����t�k�E	���mkk�m�,g(�^9�v��_�O`��t�pϼ�&�H��ITc�@$��lމ2�Í��zn_1����>�|�5�dJw��仇,�%P�슠^K��QzVi�w��ۘ�)$�B��L�H$�;�I2��yU�̜/WBB^7?�$���]xe�����C�׼�L���I��|��C��ВIyt_H�(��gtI����A��;����s�m<l�u#nvh$�y�&O��&�ǃ)hI���8��0=u�$JY��6ff`�:\.��� $�(��f��*ޣ5����x��Ct�ݨ�I$�m܉3�AGgH��bY�������_{аg�5�.�̘��[5��Ҩ��Gs����n�df��&k]�����c����������H2���M��%����t"|
�>�dM�=<�A-�׃!$3� �H�wN��
�'٩(�U�Z��ݡ5������#UEղ�8�\�������!�xUe����1W�7��Ov�A�����i>z�95�q��>$��	J4!�+2�� ��Ĩ(R�H-(�7w�|�mᙙ���^���S�}"}(����O9���H;�Z��Jr]���$�y؂m$��t	�JJ32�y��^��fd�;�	3�SY��!x]˂�݃7��U�1��\�3\68�.���C���	 /cdL��H*������l��,�극S༬B
Q�N�;���)W[�$JI8`�ϛeL�'��'NCv��2W
�R^	��$�	H[=� �95�M����m��V�ATżpLP���cXp��nh��H�ha�Ź��筿�m�k3�������h%]})$J��&|�\�n���;��zZBP�=�"D���ZA��f��CHK��$�K3i�顔�aRI$'�dL��@.��(��;��U���^�͢��"��:fR'B��ԉQ)*��%%����Hۋw�l�B�Y�͞���>ZFM!�OT�g��=\����Yk�������>;����.�͏5�&�7�ùK�=�z��V����>��������(A��A�@�F�I!�Z@�
���i@�f��|I �7dH�R^At}�$JA�j��S�O�L�+au�O<���;p�	t��`O��%dfș��^KwCs������ܑ2��U�r��wA1�.ɘ~�RI,u�V�1͋�}��p���
��e܉:y���ݑQ	-v���5hM�?KEs���s�f�6���p)��5�JFZ�f[;�toq�v�������b�k%���w!���%��"})$��͉2|PKwCHI��X2��"q��M�ȑ)�E���ssc�L���:t��=���RRi��(2��=�srb`L� ^�f;�&|��!��-) ���W �S�t��6s֓8b�����%�ue$����>��U�9M�F�zn�q�%*��I8˺<��Ҥt��;�Lʘ�tT�On"#H���H��ED�+�fKá�e�$�F{:����Ug��)�2���pn8�c"*nMk��޹������VJ|��r3^���]��٢!�w�����?�~\k<y�o�6�X{���'��e�Z�U�dZ ��h"@
U�JH$ �8�q�3�L	��q��0Iv�Ι�VB����I)���Y��ܯ't��8.sdL����>�O�P�΁D7_^;�P��z�M�h6\�جW�.*Ke�0�mkF�TyMp�v�,]j�����.4�M�|�)>u��a�d%��b] �	/	��)�yN�v�7��hɑ>�I�]��#�7��[3��CnԲ�dG��f5��ޠ�n۱{Sd����e�)��Α"W�g?�Ȝ	A��MS��^�69I��;N�Qk֖�t|W��́RC�5�lDC'�bl����D�*{:X��C�"�gY��vTԗm�:�H�����+�i�B!$��d��(-���$64��x��/�a&��� JĊ;��ZWMH�I%�;�A��ic�u�	�$$��ʐ�)F�H�J)$�$J�X{3��y�j�e��,���Z3K�����ٴ݌(�u-�����e��������C���W���Hb�g5z��)�~m��݊�}z�Òߴ�� �x�}�j��f���vT��s�V�'{7�7 �����#��zB�K�/v�U��kI�{<���~׉??S_�z�8�:rg����k���:g����I�[�Pi,;x�SHǚ�м��g9Q3�9}��P��m�yL�Ӭ����0���R��Br��l�Ow�輳���R9��;�i��K�c]U�7��naʹ��Idd�;��s���7�^��[�*E�߽�^��� �{�=C}��|<�Lgx���*x�w\[��9{��x�s{����r��c.�DJa��̃�V��&�q�HK�C4#%��$�xv�1�g��S��^�M-k|f�?ڼ~�A�&�v�!��e��v��-}��nb�-��{i�K��Gh�=�����B��Bpv�Lv��y"9
�wG��;ǋ����Ak�{��l���}�yY��޻2��R����΄���NG��=tP_��;������X�ɿ �ՃU{�n(s���!�����I����@��O��bz��Bx��v.�-��w��:��Sq�Ĵa� �X,���a�ޔ�5�ޛ�n�l]��0c��^�b%�����m҆��/[*�+��7�8����'{4��y�7��/$<;��ּ�w�]�͘�3���u�p6zpү_8{�	�h���#��*�x���I�δ�b��/M"����!TD^TV��Pqe�N�,Ƃ�5�q�I	�ƪ忑����N��O��:�N��p歇*���>3��P���OfQ	��Rv����Ǐ�ž��%�S�E^Eyza�2/�98�{��d�r�AE߿`�%$	�1�������2�L�<�µf����������q�� ���0�h�z>>N�
/2?���a��i�˲a��("�	��{j�vTM/\�+�?�Oj/7Yc��U.A�SDɬǑ�aM.L����$�>N�Y������#�*!���Tf��*�'���+��������̑J
�)�$iFn�Na*EI'%U��͊h&^W���TDTPY�Y.zd�O�'�j:��`�\*z�C�L*#�>�*�KK�W�CV׏l	
G�J���_��m)(\G�;uXJ���6 מZ��R �F��H�z6�^y�]1�9t$v�mՎn���6���&�mw�����.�v��C;.-�ٞw+���J��#�Ŷ�5t��8o�/P3=�E�=��׳�9���y�㣣�;n׮�P�m���EA�"<�3���0i�e��u�:�����+wlkg��u�G\i��&ȃ��\h���kWcLH;4��7����upӷ7��٫(J6u��:�Q��e�[q����&v��*@rB�ێ��q�k���nc�ja�Xng0���d�[c��KtqBjFXV���A�������O1������nĚ�睇�	9���3����y�]����<ڰlGk]���峬�C)<sG�W>�1s�6��4��Zx;����r��G1<�ԥ�E�8�PŚ�i4��К���]C��{f�ts��vc���g:�mn�Y�a����]C�ZC�n�f�"�q�MF��*��"�B�I�û�-o=q<y0O�I��@��W����U������mNt=�`ȩ+��]�u��
I��15v]1����I����9+��ve���7�y3�&��Mu&��0X��Q]tF?/::.Mi�0:�: PԽA�������.y�	��\[ǎ���ղ�F�\^�m�9�ۧ�=[/�"L@#�4t�f�Rj˸FN9q��F�����L��mԓ �f4n��m�!
ZKJ>��5{�Z��8{U�n��;le�+6R�p�{@�Y� �]�jѮ[j�Z�M�t�0�������6�X�jz{Xы9��sZF���J��*i:<��7S祻n����@�wi���[R�;,�cW���e�s�Dl:�u�+�i�q���c%�vݗ��)�r[R�n{&�WeX��%5��7:7k7��`|��ٻX����� �u۵��2��;�pܷl�G��]q�=V�K�֍gf��ָ���"D�ČH�	Q D
DL#JB��ЫH�G:y���\ktU�+�6{�m�:�,릌��h��ɋ�/=y�	��E0\
�[��h6`j�͛A�I�6nv����s\;�!b6�f a`Gv����7ZM��<E�㸸��Egr���{�⸆_M�ɻZu�)a��c���\ëu�4Ź�kS�)��U��ۑ���:n}��[0n'��%�cn�K�ء�������n�l&��\ԽJ( "n{G84��k��ݺ�9L6{G�����>��_��`�����O��2$�Q{�&RI$�:;�L���R�*	P�s��Gv�� �,��
/zD�K��V�ӂY����RS=� �!�:�[�i����� I(��!%�$v;�L���i��g���������9L�1v�MK.:D�H$�]�&RI&����'�����E(��%���s�,��]���vt��A\sT�\�[�-Yz^J�.�^	�/$L�f%�[�襝���7wAmmȟJW��fg���KJ[�Q&I�-���Sj�.xH���I��!$�[�H�+� 5�T�!��j��C<d�Y�!��0!��G������Zz�Hr���!e����ʮ�i�����?~�JNӳ1�<�ԉ�H�Q��$����*R#/+�$D�[N/��'BHQ�"���p�RIv�9Ma���m�WL�C[O6�A�B"��3l��oh��eL�־�Y�A�&�M)�ShҿgQ�t��^��q�>�.ïj��':���O\�[��O���D�Б(R��B 
"P�@�@�J%$J�ͨ	I"P�;dM
f%Fs�*|�"�>[��ٌ�œÄ���N��)�����*g�DJH$�ͱ-!��%�F+S�i\�)`f��ޑ�Iy��%H	.�ޡnᜧr�J�u�"��J�w1,[ua.ꘑiQ�I$B���R�	�����3^̍F���k��"U�%���3�.Δ�ydsTϙ �J;6ӷHoF����J�2D�H$�;"L��0fAOgH�Pr��;�^�b(�.��@A�`dHlGlBme��2�58�Ț$^X��m�Ͼw�N��ܻ-bk"���$���k�>��J7:DϒY�/���0h.�ų��+� ��e%��#IIúvf4*����"@��c��<_tt��̩�2�A$�b`)�d�K�ozD����d�aW��?�����̄�L^�H��U'�י�I$�nt	R�D�Z��(n�WƮF5�'��r����j`���2�0@��b��&/M�d�T4�����A�ڧ��{2|o�����O��(�)��C��5 �RR�(W�3z`w��$�l�bI?a6�i���I�jӲpK��t�.�*��1(`~�vX�]��I(flx��K�$�Qג&G�I%�;���Ɖ4H��[�����ɣ@$�d���wD�w!˵#�W%��;��[�]�;Zx����H����M$���$A2����B}-9h��,��t)�z�j&���P��.�r\���0ƛc�]9t3=V%�]��2t��,ܶz�d*��3��&Q)%�i�i���n(K�ƆD�i}�2�,�[="D�;� ���)ùvT��srPK8km�]�7�YO���A)��)$��];o4�(���X֧�.���g]/���f�F�úvL(Qgف`J% ��ސ"RD��m$�V�ݗ�t��N�	/$����	$�w�e;���A.�wp�z$'��]f����$��5sd	RIy$�{d�A�$ٍ�j�-�V�:g�Q9f��h�j{<k�	v�N�޸M�w��u���Pt��LU`�бd�FMɷ\e�����Lũ��|��x,@�#4�@�-(4-P��e׾�rvz�ƺ���p�7��:i�JT��D������:�22)�N+I!{�"e"M��h&R|�x3��5X��N]2�	`�*E�v%��"TstP�׷g��s�u�!I��)6f<q]w���\�]܇,йw\a�K� �;��J�I�z$�I�(��	i���Q�bAD�����J��lc�wfN���5G�du<�H$t�9y�&f�4�e�c1���/$�V�|�I3���)Jv�;5(E��>q�JBD�Y�X���ܻ+k	jɶ�2	X�\�!$�K$���Ⱦ9� ��Zӝ.}(����O��$�F� D�$��t�0�4y裢�r[����$.�I�V�(�4u�џ$�AG\q���s�p잂�$eNcO�;��2+ՇK�W��'ğ�9����J��n�%з��4�4�D��<P�̀Q�fT��Z�Jh�=/=�%L]��{��2��^v6��78�s��#�r���{p��~�U���nh���3��³M�"T�Gz�	խ�����:π|�""���F��@;���-ߚ��Mc���oy/6+4�\��;Ff���c��ݮ�"��r�cY��.�[{�����{9s�}c�nb��M%��{�qnz_Lq�g�+��k/g�5x���\��9�� 4ob��E�X�"��b �us^�á͵-�T������i�E�k��z 8�<�\R�1�]c�7u�с��r��3��ˎ�kj���+)6IBˌS8�1�8� �۶R����O:x���@wW0R�g������汝7�L(��A�I&�׉\���8̤[r�z��ω;GcO���dI���A A7a�����%<���֣��3�(�Iy��$�)/(܎3�(��,�X�o%�<�t�J^q���3N��v��,�����+&S��`�Ix%#7�õ��C&�RI&�x$�I,��� �ع)ùvRҖ������S�Oͱ��r�(��&+_�HI$�7O5����$��*�L��q"�ZÇLP�E�^M�K�$�wT��V*�Lm�`Aߪ$�)%�"e����y;��_G��ι��*yg{XK��3a��XKy�X�k*J�"q��r.u3���0�ܴ�����+<�s�g	�u�	�g�H��e�	��H$�7u4���r��cMe<	 �
3:D�L�V���:o;t�T��r��V2�۴���]nk&DU5)P�L���Xo��:]ܐ�%Z-����.l<�uOOh��,|�����]JL��ļ�ǿZ�z��,��>B@�D�$J4��BR
)�uf��$F3�L���+����QA!=�O��-���g�2@T0Z��pK�'!��
�zD	�6��y$�:�kz{c��}4<���G����M"R��Ή�];:E������tպGI�� �U\�e$�j�؂Dyչ�[Kv��4q��C��zd�7!�ع)Çvi�㦣!�%�3�A�����p�gp9�&g��F+�h�>-�}u����w�)=f��^�s`ݤe6	�\ݳa���
�v�݂@# �&�q5in�O{I���ó8qk�؟�!��Vu��:�0�c8x����FoT�	�i���k}l9gwL�e���A �ы�ξ�z�7dI ���4Kf�L�p6r����P�[��U,�X��عo;t�>����۱ ��r'��n:GM4�[��i�]�3�N�A�NcAI��4ݹ���4pY�.�a�wW� f.����u[��\0pG��� A �|D�DI@(P�T)^BMUz~���M�ϯ��VS:	wd���Ω���.�M5�H.n堒[z�d�c���7X_�$B��|t@�b]��,����TwT��v�L���sQ��Q�}K"Z>$5�tωF�T�a��k܄-��L��ŋ�LI�ƭ5Ü�ڰb���u��lm�j2��5����#4���û6�2�Ál�؟A��2{wRI��U�M2�I-ٻ2xM� i%�8N��t�Ϥ�ëLǰ��y���w���*��O���8���cF0!n�����K�+��t坝3�y�ڝ���@��I,'�|/a������h$���$�I���}���:.[���5Q���vA���z�燾�G��@�Hw�2'��3[ڋwR�(v�ۜ���L^^�n������J�k�}����;��ܔ�<y��yq�T��Ä�"��%�l���Ï��@ ��#�$@
PPP���vD��x+m��$r�2n~�>$���½��N��IV�w��1 ,V���O-�h'��3� S�C��HC��u�q�E��8�v�Xk��n}s9���Hx�j�rҝ$�Ea��]�gt�����2	$���	 ��g�P�[l��UXΌ��I�ܩ���(�g�N;�DW��N��/,���͝q���4�A����A�� �z��5]u�ZC���&��P��YÄ��%�f�H'Ǝ�@�w캸9�onj�u�H>�����G.�h'���l�vr�Ιü�����޳�{t�
^o�	$�K�O46�@4`�fwrn�!�{b}��/�:.[���5W�Ꞇ$څ��4�����-fFH's.�|H�9�<��K�_H��p1�!1t�(˶0��vQk2��#eچ���u7T9�d:�z9�����fx�w4g��.�wFK�o2�3�����7'q��>��t��zm��r!$8s��+2�@@��H�}e��gs�G盠���+��i�����i�s���cn{&[���$�b�\eq�v7=��>5����sE�)%� B&���XG��P��ݺn��6a�6 9�3�*�W��栲
&^��zz�[4�c�G��4�@$�V
�����.��)7D�6F�v�M	��n+�f��;�����eu��v��j���㍷�:^0�Y��a�ܹuHF����ʹ�!.Tx�ع�[n�吝�S�Aw.B[��ͩ�>;�uG��>m�ύ�n�,�P;�����(�Z����衉�g.�3���F�����Wn�EQ�]�"H'ǹO( �+�7�f|F~�O���+�苓ٰ���%�g%ݚG2�B�_s:�K�p<qn��z�(��:��O�:�d$h�
V�K;������i�>�&��-� �ܻ  �}�� �I�Π�v9����d�?b�:��w��;Ćʞ� �L^uO�NN��Y�-�-z"�re� ��ntϬU�b�}x���i�(#�("�@��f�f7nSB�{iz�3��!��n��u�^4x�fI���r΋��wM���^�ē�-�S ��p�c]4b�|co:$�k�����x��!(�%]g]	����L3���_��<D�9:b��fJ{9B`���ә1ց���y��K��rc��j,����޽��z�ц�=��'���B!�("D���JU#����5B���!L��\�|� o=:4�N��2v�	�r����A �n�H$�`Ӭ��KW'Ҕ5�L�H1���݄m��.�.��'��\Uλ��1T�\H�> �oT��ݲ�r��
��٫��&��fI�	���,�JN	�%�f��|I�S���{�s�5�6u��Q>$�^�H�|{T��ns�4�)��(�ؙw(�])�r��Yݱ{Y�vi���e�[�宱N��c�3�gwL�߸6T�'�/6�H$��g�	�q8S]�=�O��$������~�w,�o;t�>"6z�:���&#�t�d��|Ln�L��O���\�h�ms�5�������V�ΛΝ9	U�ډ$�}؂d ���:�:1����G�E��ر��g���������@�E�@=����A��~\�p�8z����oHѧ�����F^㰃!�W{=ut�O�����/jX~��i��mΜLkՋ�=����'7kV�w�^�}<��h@���A:-���ˇgEI/_����1xww�����~�u����s�f��={�]�lcTj�@x{��}���{Q\w���w���ʭ>>՞�W�. �ٗ֙9�&�i�����x����yO<�N(	�7�Z��=dM�[�p���������y=e��<�����5��hQ���kܑ���=�"��=`*#sQD+���N�;|�ޗR��ޤ3���;�\�{�X�Ԗ�E�6y��<��5�ީ\��	=��A�����������Ϝ�BĀ�w�L�2�^c�eO�˾�6z��rr���,��MfDDݣ�,�<<]l���&�O&�|�>��<c��G`��ii���yo�����W��Y�n	�o�{�ჽ۴>��8`�w+sY���\�^�D��ً��}7=�o�uA�5��f"*�3wGt���=��B��;�A�b$`H�p���'���3��� �!�P�xox���oDbg��f0̹���xRX�Lf:!�P+���8<��������"��'	�{sR��T�˄;�{�'q�4��V��_.��k�G�̝�g�^�fI���x�w.�����,�P�~��B�h�2bt��1��uJ���'�
!�f>)���5���Ć���^c�4[ظ��/o��~[O4���wS����)m��
BS���0���d�WǛ�AW!+�Q,���t�CY؈�x������Xi	��'�M���}��$�O{�υ&Ԫ'����8�����������z�G�W��m*nBzBj&x�^^��$~?����N	i2��7.���eǂ�L2y5v���}O�fɒv�g�U'�Dv1�����򟣽F/Ū� �oY���_3ϪO�R����(7��(�p���D^��s��uB����I%��`��kEk`�B&<�6����J���i{�{��;�"d\��4g.ü��3&乓��z<��$����YqL�4m��RVŢ�F�fBR4a���2d�"��=��'dD��2���-�4)��
j\=��Ģ���0���M�(���d�a�FBfa\��4$B��H� �)��׽������ y�����������ſ>��z�t��3U��D̀ۘ�*ك�����U��A�1x�sSs&��+wtK�g��d]|X ��lH��߹��N�MVU�$��<x�O�{�gū���؆���p���ę.�+�%�f�:Yk�	3����<6�u(1��Жq}��Ե�,�Jv$��D_zO����ׂ;�$�s�����l�r	 ��x�j6Y��fp��CmuL����c��T9e�\�/�������Y��g1����xI߮��r\���:i�h��Il�ȒI���k�ύT�®^�A8/9�Ēk�D�Юܖt�t��KEQ�~���fޝ�]$�۳I�i�蓡!-�/Ht�H��n��ׁrr�,b��;���GD�T�kl�!�Ht�rl쇻��٢�C�`Է��5��)�w�q>M���F��f{=�WB�盼w� >�KEB4���p\�ɇ���i�w��0x���0L}�1/���w6�s:(��8�h=^�ω%��s����	�NI$�ཌྷtg�g1v�s=���S�A(CK(��ՙ�vs��w	�vp�컈ۋ�$��݁>����ǻ�8TK�Ѹ����O�=�"|:N�KXN�ӳ"Kt�Ȑ�m$�6@xA��M���ד>$�!N�T
���"�qR♰.S;���8g���	E�L� �N�8�*�[w[� �^lO� �oL�]���'%�y�3��!�{�#����5p��=li �DV�ȐC��nUn,b�C(JA���G�U
��gf�;y�ύ�uL�H~݈���	��1����u�D4�l���b�fD��K��h3}<v> ��2�ۢ�l����U�v|'EV�/�7�3�̝C�7or}{sN�1w�m�gѺ�m��$\M�J��5D)/U.�����������!P�(D"��fg=q��ˁ�;�ųz����淝����r�WC	�V�9��t*qq��zdٸ�]���͆U�ە�q���,�d�{��vkr	˫p�n�s*�kfɶк�#4Y�e�gdϭ�Z���d����:3U���H^�ֶ7�V2�C����s=�gN�n2�YQ���]=E8�)���Ν�w&�Q���*լ֮��]�f��p�j�B�Biy�.������u���n��q������?���p������+c$�،!��4u�n�N������3�A��3}��ZY���.`����D��a�T]��6D�Lh$�c7�d!���A��[L���tf��M�Z��'vI��n���^�yA''V�����{r��VtȐIͼ���ah������<�m멆��u6�h$���$�V�L�|ޙ�z��U�u�6d�~�wI�t�NX�L���( �E�lѺm�`�=r��968`z�ٟ8H5�H'�9�d*z��G�����N�;��32�z��| �v.,klv�	]�椅��W_�y��Z�y��y�q��	}��G��Y�i���y�� �>��K�=����ŧ�;�d��D�GL��]W�Y�!��J�!Y�����<{J�v�.��n{�����z7=<�1ާ�:��$�eQ�<Y�Q�[a�^w�?=�� x��H	z����h׿�yr�|HQ�L�B�oO����ym�&�p�]3�we2�5� �[�>'�NL�Tl��כ�	_-���AY�l�����gI���=���7fB�����3�����0&&����|z�1[����~�*���.�+RgE3�ល�v0�A��r�&�8"���������	���E�cm��`���U�*�9���K��`|v����9���&���˶.f'^=����2G����o;��`��.�|5Lc<y�;�0���F����e��;�$@��V�fs���̪�gK��i�/!�\���'�����$���i�2��$�h�6	�<.�p]�gL�g�6d�y�n��&۩���&N��3i��C�
S����{�8��0���R񌥝�ρ;���UV��G�9����6�.�iq#-9��˳`"�&�!�)H�޼���{�r>�� EnB,��ӄ�ݔI솶���֭��"�y+�n8	"�r �я�*��kr�ʼ�%uwL�\�A\�&t�ΓA蝏A�1���p�Ul�U-�����	��܈�����4u>G3��{�a��}�r�q����.��<i3e�*��.��Vb͡��Ηm�0��i~��>OE���<�71��s{"	�`�~�ƍ0�5��}2H'�wr< �}�wI�.��L]�@0���H�s�X��%^�!(m�@��}��I V�~0�n�;խPL�19�}��\.��/39�wu�P(Gd��9��3�ۡ�^4@x-��2���A�̀ 	P�`��v��Ι�>m]�4.ξ��T��=��N�6$�;���ga�'����\��5�y���W>��Ч:;�O%��X�8G�hɵ�CQ����u=�N��-���L��z|�v�� <s:�Z5�/z-z99�h��%�X�����A7�E��ӄ�Yݔώ��� ��_D�V:)��͚�W��DDA��Bwk�Ak/e�hh쫭���Y��\�n���6b[��`6tG@4�e�i�b��88��u�Z[���?R�4����3� ��ClyA3�}(HX��J�Q���J���}w�<O�K�]�E�$��z���s �[o�-u�ͅo^�+���� �B�_�@#�dA�
���C�r\�y�w)�.��L]�M�6�D���� �I�\��Ftu�'����|0$���2z�r�Cw^u�cugR�#��)T�\�I97�"A ��Y���bS0��η� ��hؖÑ̍�ٙ$�{7�T�{�8�5gn���$*wvdOv�z6id���?��5Bz���Z�lؙ}���$JcQo��h�u�徯=.�Bn�5$�6l��D[�҄�2�hS��,Sm3�ŉ���@D1
w�ə��kNpp����ti����S��UVK��v�0- UJ�s`a�>��7<�j9�]Q.:�̜�s�&�V��!�ݺ�qj�F�b�6�S�m�v����tP�+���P���nx���J�B���V\��n���Y����T�U�n�]�q���I�u�p��:#&k�_/l�M�k�2.ڊ%�Z����HgEY��ױ�wL,\��Yu�c�T]9MT��m�T�Lָ���[��p��;��n��V)]���z�"�����}���Ú_I���6�L��Y������@Ae;���qFٵ� ����$�ہ �Sy��[<�㢌�q�H�x�w)��`�3��[3�A�p�"%�m��M-��Y�t�;s�I'�nz�S�;Y�:�U0���΅�`�O�� � �n<@&z��i�؅ϔ��I�f�̓�9�'N����:� �t�����Pɉ��}]I�l�	ޛ� �w��AΆ�e��A��'~�ɀw-E �# ��t��{[#f����vζHf�`��l�ge�O��{?CB�K'fA����̒I�ۀ ��O�a���c�� ������d����]��kr��;��${k���d������lԧ��y%���TF1m�sGY��I,5l�J��~���`4^k��"Գ�X��1�^!`��i�>��$"�[����>4S�~u�%!#�� k�t=�4r�qr�6|O���3�1t�9L���=3�L�6�@��*p�la���٠�I����7a��$=�[�EæN{^h���|MU���]m�	|����ܿ�^��^0Dk�Üc}�e�`Agܷr���N���3���|_3�$��5{k�1Z�"��� ��'X����E��b�ْ�B��l���^�+��ǐ�v�X^^Vg�;|Qwf,]�+x��D3b�	;�2U��0q����h�	"����p�7��p\3�zͫ���?nmG:��5��e���	N��H'�9�2I��9�P�֎�-�!� !7��hr��8d��D�{��%볢|AċM�*�(��������M�M��%�6����}��ຮ���0�/C�׹j)*#�$}�O;o��}������s^�|��$@D1 ����?=�F u�\@'�__�!�A���3Aܳ��׺#.�/+k��E�S�%�� H��m��p������'��	yr�qIæNYy��=2>��m��j2�\{�<Aם2O��ڈ5I���R&X���O�l����e�WT�S7�a0c��Ax�����6�0B����þ��;�XWY�}'͌|>6�{	�ڈ�0�5�ڑ�ۿ8�^k:d�=eN����r�A�ځ �xs8̡=�PA ��lH ���k����2�Ş�p$	�V(%�"�23u�2��ǵ��j��n	�·������Y�� �mG�J�ؐ�Xgd��L�k��V�޳I���$j� �H'�* F�s�1�ޅ�Y\�M�"�+�L�U�w�e�|��͋��_قm��r-�P}(nXSV���,�O�u����k=��w��r���?i����_�KD1"���ﭛ>n�8&b�;�p����D�'c�*��6��Z�7�z|��A9{Q �7c� &|>/��<�x}����"��Q����Ѩ���e�蚺�n�,%L˶��q��|��<�Y��N��^�L�|��ǉ#�9�."00�i�GF`�2H���A3�[�O�v%��uTD�s��,�q�狉�֮��O�#7f 4�	����8D*��wY�Q.�.3t�5�NSgAʙ �mG��r2<䌹�+p�FK=�8�^'ă��<uls@'��
�pȧL�̋�Ι�ڠ����A�ۈ$����}����3Id�u�/a�*�"�� �\��vI8d��d㫸b��ؒ����fu��H�N�Ȉ���##o�A�'�=u	��/8j|J/`��W�q����}�Øg�^��!��X}�f�Z�@������:��������痨�W��g��Z��I����K�=k����-Kw{��9�o����)> n�I�w]�����u�d2���&؆��uTp(U�=�-���/n������Ý幻��{Fm~<�9w=�﯉R��4�����s�=�B��~���<|�+l(M�0yh<i����}3��#g�N��E�W����q/$Č�%��Pܾ{��m��m�!xl��za]۰=���^sA.#է؜�/p��M�_�7�u\[]��z���wX���QP�}븪'�$�ö������oohM\�\@%���4����үjX������aO]�R�w]Zi,'���v0G�;��l��a8��N�������/L���3�&��;2�A����#2�>E=�Ӥ�P1�V1��ʲ�,�|sf��;�rK��m���g����ݺqޑ��X]��5?����':c�{�)�S}MKÖٹ�5j���O���Ν�xMԝ����WnVo�:#�g�t��o�{���᫗���`�'{��飼v�~﷽�?%s}=��b�@ʃ8�D(�Rv���=���/zyE�RhgV 4.S��gC�qrҳ{Ƈ�g��ξ�Ỿ���zGާ7���{�8���x�.��y��U!麌�N�����g6��t��)y�zf�훟�X�ܛ!W gZ<���]��|(� ��f�͙��d9x�Y�y3 ���d�Br��H�7OX�(��7�g���𵱗��'��*&|���"cOgS���	��l(|i!c�!�k̭jci@�d����.R$:*}r��&O y��<&1���||�~N�h&y��i�uR��W�T6��Ž� |�&�P�%|$c����V�2/7�v�{%����%���'��]q	��!�����||~7�}@�,���Rö�~|��^^�3�w��z��6�E��؞��M{4K��"�0�B,'�rUHު�E9K��\����Wn[�`ӳ{nA4'��*䘌�׉��P�]v2)*tǓk�I��=����I&ys��PU���"���A�e*G�0�y��5��)	�-�_nΘeFQ�#�9� a��$Þ��m*�z��Q����Y�m��=l���U2���>�{����煷�^��=re��68��c;ۖ�v�Qo%���a
ǫ(�pm���WV^]�n�VU���ɧ`]�7QK7hf,r���wB3�˲jˠ��E�Z:�[s�qfR���NbcÛ�궳��ϝ�*��Ģ��7�Ն��\�4,\���6����	SBH��t�#C̢U���*\�y�l(Ҷ�t!V���Gs��lю�vY^�2�q�	���d�On�pm�ںݮ�u٧ӹ��b�|���iywb8�sV-�b�4�p�
����R��& ��p�Muz#���Fwi�g�X��%�b�\�B�j*���3�-��aՎ9�	��ƈ�;*��x-!���8s�ȫ]���΂[a���1��U��!�qp�e�G���F� 1]��6� �Fh�i��M/�c�%��ǸtY^ֆ�w�!�p�&�AnN�+�n�/S0�N78�F�A�X�m;6�6�8ԫ��/	!�U��WK�p�ۛ9\�rL�a	�s^:8u��f�W[��a(����l�Y�s>�Y	�이'Q���l�u��Fے�ugrv�!�;����2��Ggm�퓞��GZ���C\��:h�Yyc�Î��w=�>x��$����Վ�ȗVݞ�i����Aٳ�|�֨o.�z����%�o!�b���:"����$Gl���s��������&����y�X��v��@A�{9c84�Y x�u�W
٠bSv�Ӻp��Z�i���!N�v�5��0J�N�ru�8�N��H��+�!-�lZ!5ёHԳa4���u%��SY�Bu9rʉ�s
:m-��!L�.ai8�`L��
튬blZ����������`�\��mɉ�u^�"Z�.��\�$���8	yJa^kr�6P#nKy�b���`�<�u��M؍v�ǲ�E���j�q�N�����|����k\�e��r�;`[�Y��}y�խّ������_G�bX�%z����P�v�+#ZK���<؏l�wn6�b�\��`3۶]3�'`^�81f���;=���u�n�]Eq��b]�¶����	��{/#��Yai]\��Wm�'V�B��瘎�}���u$�=���xۗ�tJQ���/.�wθ��\Ptt`���v.KN<22��E�y{���Wjӎ�ʷ3cP�n�w}�X	��0������qr�����x��������.̓����S�A�݉d~����h�:�f6�dNZ|��T�#���c3A3��ĻXU�L�K3�I�d.驐H2��nY�L��,ٰ}!"ᵛ�aF�uI>9��'-��S{+�|�=_8t�gbX�T#�1�#���I��o�����c�ƍPH�o�A`�\t�0vt��c��v�6tG�R�����/w�!��v�6�V�,��]�9xWJ].�E�vL���_c	$�m@�x��ڠ�C��H�j� ���Ι$7�}�u�{�>���#=��!2C&��RY�[�0��kn�,�2І�Q�ѭ�y����GU'���n��1����O��>�mD�˜��M3+"���I >fd�'gJN�3���>=3���P�7"J`�(�f���W��R�djq�
��(����QԁI2��|;B^�kM�س=��gTigdV1����g�s3� ���n����U�<���SXK��e�l>9�8�F5-�G6x��dΒvx��="@$�mG���c��b����u�΁�ݵ���û�Őv�L�`�����aى��|�Q0���$vvDx�}��i"-�:�U�]"\<�:L.TɌ�|�!��P�N����LE��$��m?�S����ܗ�E'`4��X�p�ny�s�o]+nlN�%���-�/T�U��__m��\�,��f��ɑ w6�C5?(2!�7Y��s��8f�і��k2)�&w1�-��PKm�ZJa
߮�7@�O�� ��#9��^�<��ѓE��o����y�p�����5�u��Dڎ��$����sk=���Ԫ�	Ͳ����?/��6=��U�^���F��SO�Ꮗ#�Go�́�����e9�j��]���G������%�b�x��^�|)���:@��<H��-�)�2gI;<�h��{:�T]�x�4DA�$�C�LuwC�Z��჆�$m؆|����3�b��.�c����5
+�T�S��EC� ��� �}�:&�r^�:�7�w�g��h�kW]��:�b��^u�4�ڶL����M��f<q]~�y��frٓz�ڏA"� "x ��z$Sn�M����݈�gC�Nܭ�	�vL��n��D�I����ښ�Z�Ot��H�j��d6z�:�Ȇz*�pmܸ��A�]�-nJdS�L�fKu��$�Ή�3�E:ڈ��$��n0O��eoL��C�k2p�3�2(�Âj=Ա��Ƶ���wd�"O��;�I����Ѐmt���&'(�[�f�"핬t�.�B�hdN�Qɝ��y��[dkʓg�B����)��C�� �A� ��> ��O�I2�Ao�S8fw	;?©�*dI �jdn��0u=lx��OF	1��A�O�{������l�UiB|'[��\�7c��E9e ˣ	�4T`7b���t�$�cB��>�����7����7P�� $��ؐ	�'�i��u��w%��jzY�\�I�":�&|Hq1Zĺ.�:,C���Xf�����)x�xc��-�H&+w�h�|y��=�t�k��4�u���&�U�;Ļ&`�7��3�=�p �o�ڪ�C��l��ۀ �}�N����;�
q�_��)ȼ�ȟ|k��6�Yg�w�H٧}�jzf$���39A#>茱 ��ť�YԂ���B�<N\�&��� �6���/��Jܙ8J5<�ZISo@�C�ZS���9*1������1�ޕf�;v�l�{?j�������yjsMSt�Ȭ��c`��/%�>H{�7��P�q�� L�F����j�ߧ����PI���8��g��Z乓r��{�k�=d�v��Y㤍z��=iѮvL��sqD�g[��=k���w]�ج�[��u�GCڴtԁ �N��qGLv�H<B��d9�."ܴ��p���a��f=x�i6�2�����P�m8�K���Z켝�g��PU3ۊ�L��U����G�qk��:7qy-�	�77tc��ը��z�vh����?y&p���?߉�rd	7�q�>$������u{�"��3�dD��>�4<v6�v`�y�:� �C\y`@(Qum�۟�8�H�ڈ`�H�9ߌiH��1+��(�g9�p��p�S ݘ��}��A��oQ�r.���t�nT��Fܭ�HNK������N����ă�	 ���8$H�������F'6	��|ko"��&��L�8d��gź�� O�]�D���˳t�x	� �*��� �FWt�3�|¢�{�ݣ���������r6}�ͣ���'�!�b��%��x��/6��_�e�М;����v ��1ս2	��Pc,4M����{z_Lj�9��;�.��)ߺd�����j�&��%^����o�r��ᱨ�Y�`<3�]vk/�2�ʪ.1�TI�ǌϹ�M	kg��pl~ ��{biu�\��C� �����S�|s�sc��A&�V�ʹ`�ՙ��!?ks;3�7���@������I'.s���k�;f��	����ކ�ª��p\���U@�G+�'^N�ܩg�� �'����Sflp4B�ܚl~ٺv��"�o4 H��\։E��b�.��rfD��$elR&�{D��#E�ǀ	���L��0���%p����5� �Lr�V��v��Kت�=�P*��.k]�罇�#SR�c�a/��	w�	��oN�x��vT���K�����Ι&`�:�;t]��Q�g�n �� Z־z(`溘$EWt� �v�@>)A�N5]�i�S��&���&p���<�|��'ă}�� ��4�t�L9��aGU�=�ʵ|����k�F�=�q�@M~Ѻ�׺H�WԅB^9�&��Yg�I���:��\�F �" /|w޾'����� �H�b �������8M�`�d�ϭ��T����E�Tē�@'��1����jgI��Y�s��D�qSz��.Y�L�����H���["Ti�ƚ6�I �sg�=^Q|� ���#��8l�SYwr��);b ��B!i��ٞ�H��]�<R^��mJ�j^&�[X�K���L_��:f�{6�A�N�s�������՗�q���^TC��-�ȸfd�f�Cv\ �]�3A�3�ص�}H$_<Ǡ�>��:����	�w[��'1�N\'$:2$�����9�x�[�k։q�u�	8�ڈ�Q �o �i�;��᝜:fy��#�8˺�l��͞]��@>$}�H1�}qUЅ;�l�D8.�{����<6�UEӹ���*LE��U�x6'ڐݘcr��"n���}�N�V6RQ�&T��b�haP�|wF�qyA�	%�\;�C�&�;8���x��B�9$4�!���u�.���u�:7�̧�/���I��6$̸f�x�gXd��^nڈ �W�H1�}�}1�|�b3�������c;��2e�|mlR�jMʹ��6������ᱶ�ޝ�憆.�k��N���]!��l�$�n�L�f#44��v��������Qm'�i��D��;$��n�fd�
k)�B�Mυ�	$�趏	����j�&�xn�n�C�N>z������2.�;��V �y�$f0�-�Y����	���B	͎� ��V����L袕
]8e��.����<�r	'�9�2O��fm�7��\��*,���3�vp��|�#fI�]�O�Ir�@��*�$�������:$K�ev�gu��$�SL���%GN�EW�,�Zߩ�Y����n�S6{������wۋ7��Y�h�U��o��ή���1����p�?�{ H�����+Rx��u�6;p��ӊ�醕���7==�۞g��Z�-j�M�#��/fhݑ:�d�U�=��y�.w]��Q�8Φ^W[��<>N�,�*��
۱�99���붼
z'�^#FmX�6f]ıs��c���.�13��lm�gǦ�g�mʤ��4t�
b˞$ �V�%��,�]�T��]3;0Q.��a�N�5g�ՌQ�lWg�
xx6�kg�>k�φ��5+�?o����R��ϧ������&/wbA$�ݲ�#N+�u,$7GU�R{��A"/of|e�W8.rK2v���b	�}��,�p�S�H ��]^�I{���()����{lE�]�"�0rɋ�
ofgĂA�فWfAҹ/o��H$E�t��C{a�7���d�.�;��S�b�_3@��|�	���Ȓ@$���	��.�h��<�:Hj�6r3&I�&q���r��Iڜ� �5y.50���^p�����I �mG���"0�CA��	��'�u+V��v3b��O=���Gf���)�=��d8X��{���>���h�æg�X�s>'��ͨ�I���Ǌ��F;.�cjr+ĀO��ʁ�)�ݙ��M�`�d鮘��'���FK.����}��U�0xT��U�N�T3�3/vt�n6����"zk;)Bh�}���w���݃Z��w�",R�^�Y��cC��x��'������� �-<�/����U	�p�:�d��DV��$�옃� �D�Ζ�[��A ��8�G�wK���b���_��b�9��7}��b#'�,�g#1�I6��
����D	����U�$��=ފ���b\32w1`�귂@7;� ��bZw��$d�D I&�%�L�wL����mY2]�T���+	��H7�A$�Q�CCgqx��[	v���K��LcZ�N����
�ðtBZ8��#k� �&s��#]>�\¶�8�8G�9�.ɱ�w.��S'",3tt��l-����µ�wl�Ѐ|I��x'��'��A&C��3�>P��Ӎ����o;U힌��݉0
/��ټ��]p� U$�&�ˤrj����\D6Q|u����<�F������=�m�-}�W~�σ��{�ͨa^C}�{�wT2w*q@xd��jU�&Q�S��K�8wxM�]���������mn�{}{{D�����g=�.r1��+��2��s���h�_H�e3|���1�ӗx�o�����
0q�l�������+�6^��Cz!�����K�~����q]�ZXߒK�x��,믆���M��֢�4s��[9ñC�s��zr�(�ڥ?��?�F/�47w�)[�ys�(;l��'^K�����0����Z����x�F���6�b�dyڂ���	��O�c�"Pv���Q���q��o�g{T�*��w����pe^6�2�����tI�=C��-iW�^�N�s�!R����xF �}ݼ�)��/^;3�*�г������[�oi帱��5����~�99+�Ne�J��Z{f����'��!2Ӎ��?iA57P�盲]u�ZbĲg_3f�};���tp��v�V2����4N�<����g�V�
w���}�K�����,�w<�}䞮�E!Vе�\���4�ճ��pR)�s�Y"�ر�d�:F�7�^uw���o7��%�_�3m;��+s��1�T1o_Ky��N�=�/���ߚ�ې~^9����3�mh������.6��9t�6�����O�o��>G=>xNư��OI�;���8��}�s����D��kJ�Ĵx�h��q+V@/-�1�J>�^�=x���a�>G��#����7��BC�?	Ė�awsX2B<��H�wi���Y���"j�g
������<v{�}�-��8}�ʨ��d��_E�E޽�}�ʇ��b1����?<#?.��g�D�=��[��ڒ�!�'�/�Rh��Ƈ�]��߈������E�H� �O�:Ð�����)z�DԢK,�d^|P���'#Ȫ#���F<|~=�̟"��a̯<���vp�9���<öv(�1Y��U	�i�|�-�a�E�m�Ŷ��[$�-�YW�0K����nT�"��n6F��irH����0rv2�/v�Xۃ�Sۢ��Ǯ�P�t�	K������+]�z�j_���S���f��ELِV�h�����WK�>eh�N���e��g�A3�D���'�\��Ǽ�ˈ�D<���1(�>��7`(0�����ѯ&e�W�3W�D���&'��}$M����/>��H$D�}3エOk��w �gi�����=��H(��8$����ݖ�n^f�5s'9�S���̛N��ŝUf�T�E��2�ONʜ+�n{�H%�F4L_^̒�ˈx����SC-^A�v�=]vyj6���ͺ�c�s\M���I����B�F���}�&%�&L�B5��L^���;�q����87_]�VfD��B�3'��BOT�@`�Q��h5�n���b��gƂQތ� �K#���(���n���"�M.hhE�˻3���Sll�>��	/���Z�#4�~|"��[A$�/3fA��;�q�)�ݙ��3 �:�MGek��M5�&��.��^'ƻ-��;٦�`j�����
σ�x���{��G�.������+�
���f��=���{Ӳ���0�`�p�f�~����ϱ����~ ����������L�U����H(���xXP9h-�yl>�޻��E�I�9�jS7���� ��|nlk���	�,�m�f9x�]*5�	�h�-�j�m����ΪP��>���S H;�P!�'ض9���N����s�g˗$����#fH����3��rʆ%���KL�
v��t��ܨ�A�Q�Дd�s� ��mf��B�ɓ�p�ASAj:<č��Wm�Y��8P�A��q��Q�M�(����p�<2��:z{�������w�]ߠ�A#u�=}��X$������vfr̙A��;J:�|zsv$��o4�+���+�MSO���@$t���1�NNꞓ���!'���X"�8�b��Q�;�w��J�۳�����7o�wt�>ʷ.��b�
����]~�t�)�L�b�X���!�>��� JE���h�<���,��:��N�+JE+5�Lf-`Flh�AE����E-������gV�G;��j�΋hi�S��3�ݳC�,�h��6���V��(sYv������V����Z�ڄ�;-o)r�vߠ��e-��&G��^1nJ�K�u˳\��
�,H�1�T�魷+��s��:�얉�ĕ��D���9�v��q8-��v���,[���$�G���vtҜ,��u���{��;bC��;G���A>>7��Gē���%�S1<�)�h� ��MCُ^ɤ�JN.ŝL�V��	���N�-�+`��}��'���l$W��B�xT���d��3���g��d��H~��D�J���I�7�������އ�
	����$4��%�fd�\;U��꜡�pz�O\�L�dZ� D�H�{c&I ���,&��'�P�c��E�Qwwgd�2y�sDt�$@H�mD`�7s��A�~�$�mz0H$L��ω�헱u�N�����sѣt"�l!���:��ұ^^T\a!`P�Щ��[�,��ޥ%������nwfg,��;X>P�~$��tI`P'{b ��.��f'!��nwy"<O^D�a�N�tȹ,]&w��e®#g.oG��p���F��N\k��sێ�SZ���5n31���4��OkI������z������;
Gh�ˆʍ�s�.2\���l5���#���I �fL�6��۲��>�W�M����S��1��,%㭳�G'W+��uҮH�"���A �헏H���3�fqTz����<�7��	<���l	燏0H���jر�&ٟ��g��5ゲ�ɝ�p��Nf���7#�*�uMx%Gq�K0��S ��&	 ��<qME��^~:��a<�|�B��͖�a�H!ֆ��8��m����Bi�̶��Fi�����~m�];/�)�2g�kvcр�H:y���Mi��a���B$�����:L���:�mGDoh����@�I�1��s��z�)�O,�[^��Ê�.�pY:L�!����[�DL���s��^�S����
u����W	�������tpk#b�9�]�w�N4�F*�bb��ՏM^�S[۳��8�x;<_�xI�zb O��|��H��&��'�;e2"��p[����=�I]� G���x �@��鞃j�1���� ���!��0/�L�O��n=�y�Μ�|�ۭtY�m���ȏK���vP�$�4O8�7�[�\��^ڗ��c��8�,�K�(&�x
�g���3;���Fs�g,�3���<�I�� �rz�d�Q�$���+[�G �ӈ�~��TI�)9wwN���Z#�I�����*-�|e�$��~���'�2_��gV�f�Ag�kgd�S31v�A�� �.{v$ ��h��s��c��m��"�u����&�당,N�;Ԁ_�wc�/�%��H4l�L�gH�GwL��Z������dTaABlM�K]ǘ���c���iڪ��j��l-z���x�X�f����nKE$gq��z� ׮q��{Ob�����;����y���&ݙ'	�v.ʫї�2	���\6a���E�"����]���F�L27�Bo�冝d2cGJ� ��J�^�;��Y9�`ܧ@� �-1Pn�u�w߾�{-ų$�t��Nm@�d�lH$�	�����*���@$T��ω%�����'��B��x�Ǉ��l���7�����ɟ'��= �6�����G�Q��$��;�wdelGL�H�]�$#-�꥜�	�*�fA$���@<v�3�p�3�� U����)�]�
:bI ��ă$��O<kR��5BQB�`��v�L��k��,䔝&w�/[1�E�c�Շ��ۀu�v$�N�L��[�p�'M^u[[�5T���@���S˅5C�d�V���7��vh��)�>����b!a�}1-�^�vw���=,vסe�o��{#�����lSv>�S����N+�#1usI��3�x����x�/f+���v<��c�W=��f���6u&��Q��(s�n�gT�V�F|�u7]��x�=��q`�#�P�뉬J�l-䠲�.�1W@l26�Ɲ���� oj�p��pDsbh�[�,nׁ��.�=aq�=�Ⱦ��s�D{��W{t�������Yۉ�u�q�kL��P�Ⱝs����#�rzz1�9�O\3��b+[�^�Nœ$�f�X�p�'b컀����O��و>��㝆'n��J�4���2I'�fF�	�39H2d�I�q'fS�<�gU�_�'��/� �A͎x4[�X�97]��M�t�8g��B�ً�A$���H�e����wj����H#�%�pHh�O�4�����;N��yEGN��S�2}7�#s6=��t���Ηz�*�zXL�g1\[dAfʈ,����:d�郴ρ�r�g�H��ؐy�;��j�fnN�>����$����c��$���{ه3b;�k�Q���^M�8�����e)7U'����x��Q�cm�y����j"��}����t|��ʁ990� }��>;�z���>�'�= ��U���L�&	ػ,�OQ��
|&w�u=�HtfHh*�3�NxO{_k�9����
7ݾ������������y�^6&�������V�) ���7�I�8��`(WV�rwzdz���h�i����En)	�39H2d�dv�`�E+�Ί$�Ď|\(m�5�=�Oo�i�H����I��r�	T(��6����Y�_ �ޡd$}L��$퓥J���U�]�4I%�-�m�6�3�t�>
�K������c9�Y���`	79� �2j�d�|{�^w���b�g��S�������*�T��bl�Xx۟8��$����\�5�L��ΐ[����b�郷z�����݉�Ov�3�X����g��O4�H'�w� ��Y�1b�)�-ǡ�>5��r�mt��Ot �|H���A=�0 y�a��꛶�q�[L�3����m̓^$m�i�]�e�/ߕK�#�^�kf�n�0��my�ٛ�y`��ј"��W��fV'5���ˈݩ$EPT�a�P�x��d��ψ>;�0 ���4:gp�d��P"z�Դ.n
.�����1 �A;�1$�s�[��cp#K,W��MĂG{':L8vpKP����Hˎ��4�b�!!��1}�8)B�	 ��<nŦ�����U,@��2����v^%��g��7�:�l�/��vt<Ԯ�홰���k���غt�C\l�$�͘�}�_��u\�c̱��e���$M^�;�:N�Ӈy�F�^Aj�U[@_k�D�A,�Ę����H��<��m��ξ&�gNŊA�;F�_�` �G�!ρm�v�C?<b���v�`@ �[�H�
�gt���gLg�v�gUs�Uc�b$�j�<H''������dE��<�[I=-;�,�k�����[u/�v
�>ۇ.��Ӌ�6/��G�<�lC�`�_mUX��P$�C��8�0=��l؃y)&vgp�,�(�N9$���H=<Έ��
� �/jɶ�p!���1&�t;����MU5!$�qb�;&9&���v���ֻ%4	�ܛ/T��:�箈�k���5�`�ó�[��ȃ�	��c�A>$t���6&q-��z�$.�ـaI�����Ėn���G�?�3�_˯�*5@U��7Ă@��� �;W�4P�B�G���u`��K5�����8w�<j9� {+v$��Y�Vuޑ#��}�c8!���H�*��L�؆D:gk�
:�5���󥝦㶼D��9'ǲ�"I �혲��2�@��8��|%N3�L'gLbzsngƃ�ǳb �*��nP&UD�x��܉�㽳�Ma`��m2%ky�����Ӣ����|��y�����^�"ְ�M�n�vLS�LB������C�}�{���i2�щ�6�S�	� �څ[�>�,e� ��v.��C���<D���Յ�Z�y*������zh�.�m��ܼ0x����\�ў~�4N�{��;T��]�8V�����3����,�T�׮��ݻ�_bM�.zq��� �n����ǔ���nm}�=�f�Y^W����0�y����!��ݿ�/��޾sWwh�T6cO��c����N�����0�x�Nv��ܶ�N{x�|<������
�1M�����\��<��$�hg��h9�{۹�
�m%�ɞ�u��,,�pn�H�;���Q�f�e�����~����N��WdG�hʖT;�ܓa_	:������@#{��t�f�#�>�ck_���+6��p��e��_5v���Lti%=�BS�<Q�rL;�v�����ޒ��3Ͻ��7;��=6��M3v&8����]����U~�:)��Ney�Z��c�y��[8M��z}��3;A� d糽�1w�cl-�R���nY[�"M��D�M�B5�(���-z�: ��eu{�I���|���<�Տaj�+|���vz��?�{��k¾K4������(���-��H~��I��o�������.����x)��&v��d�;ݶ���O0z�xxLk��3�w�mݘ��ht�5t�k%�Y�\���q���kG��k($���`�����A`d��������r���}��>���	?iW�%��b�p�-vX��^�OG1n��Ý;�ӄ�vKb��۴-�0�sj�$	��^=t�m�{�S$<Z���#>?�o���=��:$Sm��V��*^U�uvIUUU3����F<~?��|��̊�5�(�jْy���(^2N��//ma����D�'�w~1�����W��z�>m��#W*�\��bg=-N�S&t�*���x^O�F<~?#�R�I��!	4�/*#��ܵ�]��T@��%��K�p���40���8�UQ��SR$y��.�*�:!^F�ٲeR�����I���r�]#�0��=�V��U�FR����^'��U+�Vf��eY賕m��(J"#fˣbUf�eE�)T]0��E�tWH�(�����!'AleR�VX�&��j��\���S�����f���q�m����2*(��24�̢�ę�S�ԷC��<���WA R� ���Y���>q��4В�\v�zǋ́Wb�2�rm����e"ੱ������wbC���m�oj�Z:��0��^�qNE�GF2[���n��Y���tMn8�,[9��#���vn���MH.sm�����A�6����ZI���[sn�+�Oxa��v���cX��v�j7vA�d:������u�0�$���m��`^�n��ɷ0���Lli��q���3+h�vf���51`5��}�<������6�qz-�vEu�m�ws�h=8y�����S�oc�Ҷ�4�r=F�"��-�q�g��qN��8b^wG2Nv�l2u攓qzݞN<�	�}c5���-���.�r8�,#�0�,4��t���xǷc����	k^�Za�s���xb��G�muC/���٭�˹:��n���p��ݏ=4���<p��9ޮ{*Ϟ�8���%9�\�έ�Hm�ͫ�0�'�Mި�o��1�{�����ˎ�q�km��Qсnq���֭�����Y7���K�P�t�̱�p\X�V���h�n�D5��V��ѣ���"Ck�Xl���]v�7Q�9�%3�1,Π�,UF��Ff�ڂg��n7Pq�6�>Ԍ�*Bɒ�\�turV�ǫ"g���y5БbM���V�͇z��s��%�2h.�Y9�:p*�ܼ���=����%���n�Ky4vYt/������L�Y�uX�V��
��v���֙�qˮrێ8��@�ny�w^d'Hv�,��͟k��l�N�+�6��v�y��ӷs�����Z��㨳Ys�Ɲ�W��&��N�r]�����f���v{@���e��2�0�v)-�AP��`�X��V�v����u�1�ceי����Rf̭Ќ�6˒i�ʰ��9�E��@N3pJ�n���[7�cT�f���'��1-��7�#�MM����s�u�q��ؖ]ֱ\\�dڭ����o��L=�97uo0��:�0P�=q���;n�;����p�3"�J�n�˖!k�5�����n��k��S�,�ۮ���z�6m��[��u���9:���71Z�&%�1��xL-m9"�]��+Fl��3�6�j�9��8�s��q=D�{;�Ým/-��.Pҭb/?��=uE�[u��q��u&.ؗF.�'���ۍ�]�n��4����v2�ǫF�a;;2�V2���j5�n��y�[�(���{0�v�6$�I#{f?Y���|�歘[��	��"PHh���7"�Ä�j�l�LD��NZث������P$혀Oo�b��ۦ�y4�B���C��gb��y�g�I�e��X�u�J9�4�x�ž`�$VU�ρ �vLB���:N�˻��G)GfۣMqbؓ�S�%�@�m<	�h�%���j�M,�|�{&I�6�:pő��!������
bM#۠�#З�\�ω'��l��Ir�`��U�z!�[no>��~���R��v����\<e�[���3[�g��q�ݵe��;��|�-�u�=�Gw\�ݗHۗ�=P���cNI�kͦʩ�	� ����f�JN���3��{-� D��j�1	��i����޵��
~X��х��=�@9��������Ōpi���ۉx!=��͈��c�Wi�`�qm7��w�϶� �@�و���~0	.�ף7����-F�nE��	� �$����A����9��5�3:��*k��	�f l6r���Wk���8t�<Цy�ar��|A-1�sA>�&.P$�F3��zޚ���zD�;���N��r��<��gCz�;bM-#2�S�eݸO��"	%��{�w�\q��w���G�Y�#c��4.����h2���l.]�d�at���Jr�.+��<���T�ҕ0��<cr`A$;y�#�7�A}�%�I�qt$.l�����kA=�
����'gLfc3�d$#]Kn	�Ϯc^3� �ukA �mGt�'�3���k~�&�)�'�*wD����A�8�4Gna��=A���/:d'E���ºZ�b��o�{�� ����v5������rG�g>��@�^�dAb�*"-��;�'̫q��'�g�|K�}8�j,8L]��=3�ye��ՀIc���^OH�	 �uԹn�l8&��4��wk���8t�=Sl�̟WvD)����0��x���$OfWL��wdDtt��3Dȩ�S͑�O����(=��|��Syݤ��ja�����1~y�x✋�[�Iݝ;�`���4�Ǡ�����$�{�n\�x�mA��aY^;�� �or~���?5�4�7R���D�k�Yiwy#���z ����$ȟ.��xƚR݋���k�6�+hI�ِd��1�~ڌ� �{7"	 �j�KbڝVu������́7�Qt�� ��D�G�\K����F�$�>LI$�v��vs'��F{))P�	t��1�`u,#2��FVK��u��%�����=������Jzt�2snv������|B���_���F���1��8���Ɏ�Ä9i�;��cY����0l`��[C��!;�S$�A��@ �2���D?S���;������p�nXx@,� ���0�zz�tY���^u8!�â٢��.��:t��c&G�$�vǠ�)�a�%n��5XW�;�D�}�C>��.�'vvt��QsO���bC^��1k*vr4'�q�Ė;|�H6��E`!3�<�F�V�C;�R.ɝ�A���� ��ƀd$x����n�&���$w�A>e���ݠU&e�C$���Μ��n�mTGI�y�$�e�Ie�� �D�OKll���1�5Ol�zĥ;bQt��&%�L�X1n�8 ���H��im(�����Ɉ���~h�'zzdy�Xy6s�h4i�So��O��t���T������bK;�8ovN�<��M�����鸺�GGe�DI�����-f,���s
�\�ID���YGq�ݸ��[<�,� �)��n��^x � ��t�ŉ�-����m��YL�F�U�5�X���b�����Yc�")6�^��pa{g`��h{dX���Mb�f���h�h��djk�D�Pc�m�\A�H���G�S��M���`�I�ϭ��O��t)Ȉ{��u�紁�9�v��V����q4��]��2[�D@kv5-��܊M�9@��-ͺ)�8x��+��&lL���ӌË"�����q(���`9�D��L��.�y�?6Ԍ��n�@��r�	L1e���I�w!�@i��N�c9+D8�����!!
�	�ޝ�$��Z�V�<,��pt̝��ك<�c��ft�O�&��Ի�4}�S�C��@$�l�IB�+�!��)d��(Ot�<]jC��_z�g���u��$�wdM��`�1��!�'hI�c�;�c:��	( f�By��%��˪�p� ]�t��;��>~7�W��'H�Q�p������zv�=����VSJ܌	�y�GlWR�{�������L8�8v��I��؟A��\A�1MI�CU`%�m��u�̂D��4�\8A���>=�PX-�c͸ò�+��x����5�i���?^�G�׻��� ��e��{P���	�&~*\�7C��;xj�˖�$��i���EnOH�	 �uǄwm?R�	>�<�oU�i)���Y8)9.�<�Ǩ��|k��� �dn����`��5k2zD�G��=��+Z�&t�ك=P,f�nSwb���\>�$4�T��f�F��$2��L���o;P$?>t�&�'
!��)靦A��x��.z��ul��C1`r�n�:d�I��,����C�`9�σ��V��̶��	���"Z���Bn,��^I����[��s��Z�Y��}Z��Wl������2I �m��!��Q��1�)�MM�ܨ�H����A��J.��ܖ`Y��5ɢ؃hvF��;��d�hn�D�ZZ�@$��g�/�R��	�O�-:R. ��P�j#b�gCFt��(�6��CHn�=���nm�W#46����O��2��{�{��6������L.�.���J�$�m0ϸ���5MX�^�S�Ă;6��s_($&��wbRr]�y��畑OZI���PH�'��OV�NT?^�Lpou��A�����2	��v`�ZV�E�NĀk6e��=)�C{ā[t'����_Hq~�v~���y�.hZ�)f�e!l#��`�V�j3Yp�fp1�@U]LZ6�����[��u��Ɉ �[dy�	jw�Av����l0x�nЏln��|	�����RE�Œgr�e�:�I9UW��==�o�#�}|� �.'m���G@���I�@��s]e�PI,Y��VI������ ��tI%j�l��ڎ�o�Al�����R�A"������N�v<��@��{�PAE4gL�|A>{�h��A�߰nįZ�ӯ?���^o��AHY*f���9��o-��vΠoׅ����1��4+��yu����}��@�T��]�^H��`��V�.肝��T���>$�]�,6��ǊB�gx0'2;bG��wdxGQ�;����{�(S���-�+�n������v{
vx/pn��F��[0�rݵ�qz���}�4�����ŧ[s#v$	'�� ��]����C��j�<`	�{2	\Q�Q('fv���򭐇�|�xl8AΌِO�=ݑ��;��r�ٸ��Q{fIF킭��3�sU��$���@��y����C���a��Č�����cr݁�;�Br��;�&A���<cֶ=\��2�uM���݌�Azv�9��/������B�W�$\8A��� �F�Ij��v�n3��3@'���2	�]ώ ݏ�W�M�O6 �7(z�A��\��<�K*��C?޿W�k�v�^���|����'�c���iK��ق'T3c��k���﹯ާ�>ޑ�����<��@^�m���i��r�N�ӌ���tNsǎSH�y9x�u3u�Z����ˑ����&�R����[�۬�|����run�\v�D�1��Y덎h�D���8ׅ��=���x����gAs�^u�Y���5ł�vR%;m�.um�#�<����kv�v�<���=���^;����;�x^prݹ�δ<N؋�����k�x�ۜ���۵�JͶ0=<�1Ʊ�˥�H�KT��T[
�j����go��Έ)ػ��|�fB@�Y�	 �7c�|fGQ��1=2	$�vDy�U,)"�ܻ0g�-:��ڣ}�fO4��8�r�q ��<|	m����r�����E�y���SzQ	��J��h��Hn��BX���s�Qr�T}�����`HK��V�l�I�ܹ����d�J�M��9����dA>��隈���v��,=-� :����IbŸ5e��a�M�gD�7��N�=��c�vDI��c�~�;�)�^���S�t��7FO��mXCM-�M�Зj2�v�k�avw�t�:�L�ƴw>���e��}�w��#3��D�}/{�%ፒz�2v��{����%0�C9D�b���]2O%^�>lG#8SS���jkf)���Ny���U�g��W��w��<���[ڸ
X^�vG�z��f��G5qI�}iЧ�}ڽ��@�k~"	��oL�|�ȋ�Ƿ�ǀ�yr�,]˳y�9��I9��aL��F���I����\I��	���,� Pr��Gl��2�^ƨ��AT�� �I���zD�]�<*�p����$ا�x��R	��&N���}]q���{6�E��hN�VH3y���ޙ�Ov���K� ?����t2��M�x3A�͉1tZB��J��[���v��g� )�2ffw���;�`�8��!��"	�A�O'&�ղ^�<fw�	 ����$KiKЋ�0r��w��f�;��[������}� �Q�ڈŔ��z
�/��P1X��Q)ٓ��}���&��o �f�v�e�3��0?��Zs%����px^5��}���K�;n������<~N|�����q=O�����NS�E8ùH�@��� ��W6!�]GNɃ�W�W�.�JZW^y�Ñ�&3����n���Xk���On�=��i��ȆXݲ.��p�늘�-��2b�Z�ު/^������t�k�(�]�}���ڇF���d�����&�R��z��;�l;V�9�!����[�U�;M�!����Y�-)h61M�ca�g��A����~���`��/�ƭ[���c�̗��/:=<tp��#.T&�3���I��@����_3����wfI\;鏺H��M�h��)��2��:�w�q\Q-�#�nB���m�"���=�
}R*�vҳ����s7ڻ6��{����bϡW����|���2U��2z"Y��u�Cҽ>3�h�;ڛ���z[���Uo���$C��'��ʼ�W���
�o��d�����2_�r]���޳��5^�{uy^H��K��|�[��|�Zz��ެ�O!;�ǽ�v��,s�s���Xg���,��7rw�V���w�&W�aͽ����/�e���ίy���980�Z8�i�,o3/#1ꕬP��#!��b�cT�?̿j�}ꔞ>�7�d��K�ܱ���K��N�Y�_���+�s���7n$���37+���?wY����6�b���/OBJ����2�z�x��D+�5
m��
�M(8��&,@�|�{բ^p�����=�f�Rv�̯&)YE�.LD<(�e���@�I5Ћ�8T{#��<~?�o�����byG�aȱ���7L�\�$+Vl�\�<��w=3��E_�G�����r���[��^W�$�܂U<�B��7L5/
�w�#?�|��u'}�˛n0���94"J������*B��L�)vo�F<~?���W��s+2�1R%E�ɍC��4O"
�4��+\�A��v�z��*H�HAE���!�Ri�Z���`���!搭�Ur\T̫0�����g8^Q�F�na!��w�xt�*����h��b��V��$T�UDf�y�Q�\ɖ-d�R�$�0����=<�ƺTD��Ģ�)$�-J)[/Id9Uqt"���q��t_�y�_Lr�2$�S,�'$܈�w�%"�#˓&]K1�s:�E��^k�T���E��琴�:/0`C�Gҥ�Dq�W�3�L��H{j ���AЈgwN�;	�tS�v��Y���1� �O���ǉ$��E�u[LU�>���x\�ab�'H�j�5�	 �����Y�0��#=Q�3�|H=�. �{��{=�8^E$�ߪgCu�傶�p�ظ���j��,�ڞ�d������3394
�`	��;xF�d�$��I���7�&u��˼BߣfIWl����I�2g,�g+��8 �e=p��G;�Y$���|A.�|���H��vo]�L�:�X�R�8"�����-�|ێ���!�hbdwY�~�j'/" 3c�!F�C�D��_�WTt��.�3��;�H9�� Dw_Keԧ؈��r;k��r"�*E��R�xh��Zq^�k�a�N�[� �G����uHIpNs=�>׵ie�ؤ�M�Y����VL<8<,��wt��:�b.���؟���4u���j9��	�w_L���w�[�ڛ��(@b�W��`EM�(�WnK������W%ϝ��\'����?�ߕ�d� ��i�f�^ ��ȂA�}3������x�ĸ�HAOF<���J	�fr�����H��%�V���!��qă{���ު�$���u6�U����A���fvg.8�2v� rO�]�D��K�տs<�횎�'ċW��3�р���RC�X8A���G�31�I�� UT�62�>.9d�[}� �Ow]W5��L`$򩦏�4qX88t�N���@&���A��"!ĴRn�tN�W(�#��D�Ow[�#9h*~FTvAЮ��9~k�Hc\� ؕ���/r'��i�^i�{��,ݵQ;�/+�{�4�w�s�O/�)���un��:�Q:3�,k26��qf.����'=]��z�c>Ex��� �3���91m\˹�cM��f��k Xֆ�MƓ�y9�k��Z��k�2;���/I�͇��xt�֑��dy�Wb�Gu���t��{�ۮb�\B����9�=&y�Z�\�\;03rEb��sq��\9���^7��f�\����=h�j���-�s�5�iw=�\�,�l&�a�R�]��j��@멋:�u�����{ms��N|�Ę�݉ �I=�qT>�]l��1*�g��Р��D��B��k� �;K	��q��],g6�4�\��0>��̙ �w��������+��儌�
�`��;
��̙ٷI����N��ޔ,v�D�w��A���N�&gL��3����6�J�ݯ�H-37�׶����Ȱ���<a/s^
ỻ�$�jI<`�1!�X=���}�C�A����6�ЍT�̝7{#��j�PL�y�;+c��ߩ�}�YD���3eG�ժ!-r�u>hu�s�ų$�lZˊ�睯s٦X97/pM;��� ��<[��4���e��A>$�m��N�&�!��:	�-S��;��S�?n�ǅW���Q�t�b��
h �_u@ٰ�=��w��S���0F�k�
�!:v-oR6�v��1M�	9b�ө)Y�X�>$�u�� Alm��Y�&c�ٱq�׽�XTU�0.�S�P3�>�A$�.� �n��v뒳���9}g��q �Hln��F킩�3�N«/�'?6(N��E����31,�������I~Y��b�&g�~��'d�~$=� \�搂L��&q���.��$�܉EB���j�$]��|H-v����oL�W�R�:��� #�p�k9ckpSs�8�DMj��-yva1TP!���nbI���A8`�0%�Gx؂O�b�P	�u�ɶ,�W��V#����׊	�*��@�E��.�u�L��{��=���۹1 ��!��	�u������qGLFd�t�`���x"�Ӡ���]���������5�6��SnI����#�����!��<x[�sZ��=��^H{�ۃ�}��}�i�mX����~Y_�=��$e���]��Ckw!�o�A"�dpd�t����|g�Y�Oj�\)�u G\��$��9� �	�;�)��N��ga�/� �WP(�M�3;���T=����f3��;���"b���$��7�${�_0n��77��j]�����~0^'�C�+�eڀ��=��tksF���\��-\���m�Y���;;�L���L ��6$	�;�1$T�M;�2.Z�	���G
~D.\`�2%څx���>�/�n�~�@�s'vd�G{� jK�fNs	����mKP(�4HO2I6�Z�p��r�i}��h�	�y<("	+�`A�T�<0�G����O�Z������uNY]5�
̗�A-\�v�)�oy��ӓ��d��o'v.���b�tn���R��Í�^���u?b�e���g�=�q�B��<k�/�Ů��!�j�r�`5��q�x.�ə$SX� ��@�	ڨ�\�0H*��Zn�/�92�~��v� �A�ُG�j�� �;�7g6�%a�V��]-Ef�fi�+1na���9�v*���:�dY2N�6
8q�y��a�ۓ 'sj ��CV� ù��[�k��L��ȟb�o#���]�2w-2�Y0	bn:���k�",I"�*��Ph ��{Q�f�76��,��L��X'�v�'�2@-��	ݪ������0"��$�̨�|	M��BP���p9@����=Q=�0�m����HA�]��Md@'��<���ޛ�KUd.�вy;�w!<���l�o��A����|5�"z�b=��u�� ��t�1Ί"�9=D��*B���9?��۶~4���k)�x���{��c�����bj/c����ḫ�i������5��v���J;��
��<������M�5�e�K�ys���[��'���Ak��Z�	�Wn��2mr�T9�q���+\�{<��ٹk���P�m�J\�a�Fܣk*��iSq������aŷ�N����&yy��G����7��{E��Ae;����-�]bٰ ���uv,�k��X G;dwnF1�Q�N׷�מ��;��FnWT�z�]7mƯc�w6�v��b�e�"�#�]���9v��y��«�e������E�LC�\���Lz$�ca�	�;�]"5�_Z}�Z�(.���!	z|0O�ΠQ�\�ggb¨0~�ʯ_9���O�vA>��H��>���m+~�E�[����gB�IN��Jw5@����O�^W@�I��d�k�f�&7�z��$%�jb01`�2%�D��ɕT��9��$����A �޶f=u:�S`pHV�`�~I`;�A"��ޜi~��$�
��DV�!�MߪA>O������D�]������Ƿ����>m,.�sh��u�6�fc��c����f�u�%�I�+mϮ?���3�!?p-z���y��>>��x7�f�2��n�� �7�rgČ5\���	ڨ���[Y}ʡ�ЧW�T��?<%���?�*���ɭ�xlа�[$�u��2l\-�\���d�!�/���jv"v_Z���������Cʘ�][����6�Ă�y{���	�q�7lS!�4�}�<	��Q,��d��۹q�${v��١6ׯ=�p�ҧĂEWOL�I���A&�,D2��Y�̃N���m�0uzH*��9��lˈ�C.�n���ǔ��q#�F�U@��i��őp�K��<��Ƿ ?VX�qRk�A>�����̷%}����������l=�Ɩ77-u�S��I�����;v�[9%�D�{88����Jf���$�$:H�����2A7�qĉI��4��wُ뛾������ ��u�x3���Јg.�<�,{n rU].��i�`e�:vb�> �y��"C��a �<%��p�ꭢ}�3a���%�.�#�/�I,j��M��������h��@�`/�^Zt�困��s�OOkɯr��.��J��h=����-�o����~���x��
B�WJk��
�h>}3v��&��y�_4�@�BY��d��*�k�KM,�`��З�ah�A<�D|He7�$�ul��؜��ç�`�d��aA���3��/=�$̞�*����*`��ѡ/lwD,���	2�����e�ދ^�×r,.\p�t��@�H�]{[�����5-��79.0��=���N�v��;�D"N�T��'+��Lt�F�kޣ�ǯ1�YVcG�#C��6�������&H���xwU���6;DO�eٍ�Z���&�2�U�~�wz�B��pY�Q���g��{��p%�1� �Vd��u���4�C*�a ��;� E؄��.�&{�T_3���$��M �پ�$wu��Λ�H3��+ʋ^6au:��݅L�5�_��~�ie��]�<`�v΋�L�O�����Q�+U�9o	uT��g�i�#n��BS!�;�&_3�d�;v�����9�p��`r{ƀH$_N��'Ğ����u�����{�.�lD#��<�X<��\��m�H�@�m��<�w�[k�,�w�4f.��9�$ $7� PM��\Z����H���H�u��c)8`��D��A��%sC�x�8 ���$��댑�}Ia{�v�F~	`n%�)�����A$�θA>4�s����O�����A�)�6}'{�=pxV��,���g���,nW�q� $�]L	��. Y^�6���,� ��ɹ��H�zX�C9ܢ]�U�[��K���vf۬޵7h�0$)��a��׾NX��4~��~������}��}���~�T��?a��*��߯���y��H� D D���� ��((��@@�$�  �kc�蘂"(	@	@ �� �� �Ph� ��@�0��xd2 �PH�@@�E�PQ(�PHDA1!D�QD !θ�"""! �H� �&C	p(��L�����V(��bb��b�E`�$�\("%��X� �
Qa��TX	`-@��@+
,��� 
,(�"�J�",����J
,����(�
��4Ư�DU�H"�"
�3���G�~o����i��}?���q�O�νn��������OF�?׎�3��?�_?��O�� ""���~���C�?�� DE{�Q��? ~�y>�������������~������8	����?�������]��@
,@���%
�R�H�H(	�*�H�D�2���K(
�2 0�� �
H J� ������"����,$(����H�,���",�"Т̠��-�}�""�?;������@QhJ R��i�'c�}>4���n�������?W�����8���}98�xi����m���G��@DE�������ٯ�=��������?a�\�������=���C?g��Ɠ��}c?����4x�2{t�: ""���Z����@DEt�Q�;�����>}����{~�������a�����~�DW��/�?��>���O�����5�}�O_�_M�""���)��BG�x���{y>��{�~�DW�<���w�"+��������{����d�Me��7-f�A@��̟\���0   @   P                  P �      (� Ґ� C!@*��4�@h�C@2��R��UQ@)T��ւ�
 PKMJ ��i* �;�    �                              !@R�    �  
	p �� 2 Q� �  = uɡ �hDd b� ��� aօQ 
 � (;�� �d*�� "�2'�U+�U����yx bUQE���(��R���UR�T���媔%J��EPQSX8�UDP        4)UJ��vd��8�T�H�,���f�JR��� ��"�3a��R�s4�s4(��j�TJ��p 9��,�"*�����%JH�)���P p1: 1  C;W@�*��� �p 8 �� d �h�(J�           � $E ����x  $9�\�Wf�s��ԥrԪS� z=+�s�+m��:��@���   ��j�ye�UJ�W ���˫eVۛ*��e�UQ3n��p .UJ���6�j���mScs5JD�m��@�   �        z�Om��Z����M���n��T�iT� r��nvp���wR͵Nl�u��%]l� �)��eZ��PJ
Ex  �/7��VYͥJ�� �޲�^N�kl.m�1��6�՜N�Pc��:�׼�<,֜]�5�N'R����:U&)@ �o  A        :�ʥ��6��m��;X��u����q� ݩT���5Isnڬ�,R�r8t� �Unn�ekK���� D �@w��זVշ;�S��� �
��I9B�j�my�@@� 4Z�  H4Hd ����� � �)��R��   �LM0�b`&���U��~�  ��S4*� i ��IBd`#e>��/������s�� ��/?�����G�Y���IO�'u��$ I6 �	!I� $�	'�$��	" ��_������y������a��9b)�,:�?]qӪ8~��mӸ�䌄�!��R3����9%b��^&؂�iM��2�`��L���F�$��������K�$�Ǫ���dhn��aQtVM�V��N�W_<��\�1�͙�e��P������h�!�m�N8,����k�gE�X.{Q��+����u�)��YK���U�Ǆ'�����Or{�9���#j�nm�Nk�R�s�	-�޽m���i�1V;��S�{8BԫF��݃e���FsTn&�(�u��jcbIY�I��E�=��"0y&R@ݙj�	��a��Q�Ѽ0]⽖s`�pU7V>�:y]9���$wj�ҀQ�Ǵ� 
�$�ԡ��_7(:�����'S]��g�z���b��0�`�e�j���Uș4�h��� ڷ�G���oB���=�-� X�˪�= ۀ����Q旷c�xc��i���届�&�Q��(GfPQ���@\�V��ym\��.�J�l�Y@��{M�]��w�/~׳�wZJ�v[v��%˲9�	�Bm��ѝt5���8d�g�oi�Q��6��v���Y8e\�q��{3^�w�@��8��E�r�5�}nhBnw<�B�\��%�
��PԨ<���/E�橝wF�Ȗ!Gw5[��av�m��sN�(y	�I7,�-N����^�T\����;֮ĕTf�i��F�.vYݶ7�����F��ws@���"��Tq>6ں0d<��"ɻB#"��	@` �Q���;N�3�S�;��D�i�\Ȝ4��M�ĵ��V�d��J�k��r�5v��e��d�	N��;CRО�Vs��ʁ[��
(l��j�G�pW2��ى�ݔ�$��[�p����E,�[��'N�n��.��f��d��r �3Mn���<�� v��]��)��׻� �{��u���y�d���K��]M�C�x��S��΢�YXD;��b�3{6 Z����t[��BNΤm���,����$�0�5�s�<��F�1�d�,�8N�����:���=tv��9��7&��[�ާG<mKw�,\���N,�7���b^��z��.������&��3��Ж���T'K�ˁ�L�����J���j#s�G#S9���"募q�hW+� K+7�;ҝ�ƴօbՅJsg,}8��0kf�ӕA�ͽ�M�uѷNX/uT�3R��ٹ1D�aFpǇss��C���C���@{pFPs^E��h�n�ã]�N1�OrIF�����7�m�[�ZkT�9���ov�� �����v��̼�ۆ3�n^ٖqI��B���n,�zOm 2Iu�m�$=K��dC8v=�5���Y�i	�D�Y����F�4�6sS�� �gl |z��5�\��eܴjs��t���7{*8p�3b� H]��U!i��b���-�m�i�1�lye�	e8|�?Lv�3y��4k�f��i,h�x5w�m�q���p��;ӟ.�#�۸�Z�ލ��sI[n�8�T#�ޅ.���d�{��Pc�	��J=�uJ������y�6ױƻޫ��&������Ӗd�A �3��������W/.�E��o*��s�ǫ���{�lٝ;���nPur'�u��&��oi�m��o�%+��7 �ʬJ���7�����-@�w�˙�(x��ts��yh�K��0	ח8b�"]�u��D/�a.uK���z����-}��Xt��·�;�7P����{�k�Pc����(�}4�(l�y%��5܂����I��_&P�z��˻��7)�851w�*�Q-�#�Oi�LE��A���,}&8�㑩h�]���R�-[I������"G����]��whRܺM9�c�8{sCOm�*5\�l�sl�03 �+`�b�e:�y��÷������P]{�VcN���֖�Zy�E]�ע�B�\J��^�GVӐ��Ժ��ꠗXl����"1��s�$9�tG$-�m�-�B�n\�)�n�[k�ٛ�����a���Z���!��ٝ4����w,��e�4W��yr#�g��w{NMH���]ۃwb��Э㎮�8�jh����/;{U�.ӂ�R�l�:vv)q�Ŭ1{�\k썓�oD��a�
��Ӵ,�fvʷ;�%@��\罹%Vę����.�e�r����T���ۓu�3F��h�Ory�Ջ:l�`��WoY�ON��xR��o�|�\JM�x}���sn����Ql+7o\�b�u-�ŧ͋��&�9����hw gT��Ɔ����"��K�Y���v��yn<���MR��u��{��v��w�Ϊ��3o-�W���#��5TR�7��ַa���یb�Yش�뚗p���G5.gŕhӤ�5��:��h�`��ۅj�W�hA%��ɼ��uUnM:�%��kD��]m�N�����E��M,�����ZF�)c���{y�
2�5e��n�u�w6���s���(uo(Fpr�誁� Bʶ��F��8��O�����=���l
�Q���F4�E7y��v,	�1���	bv��z���<����f�D������-�Y4�T�_n�/j���?y����s[�}�2�J��y/60Ճ��9�������e�cf��H�rr� 
��t};j0�Ã9�Z9(���>ӱ�ªm�F��x���ڝ�q���Ѷe��3�V30���s��k�u����,��{.t��P�U�v�۬�oW���	�"�ǫ]�jM׍^D��$\�Q]�sxm��fLd��Ve�6-��\ �j})��v�s{%�E��={$��&�4l������"�օ�(r$,��sd�@�`�Q��1��=��r���8��
4���Թ�jr�SÐ��I8�СG�=��A�T��$$�]�I| ���N\ga�i���x>E�費:��|�9d������HcN�u���Zj������YvH�:x^ ��m]J���qa:�\��`�ɶ/8�;�#��t7h��Ęc��V�mz2T�M��׌��ۃ�ۣ�m���[0t@f���p����p�9�s\쏁}��v�E��ٽ���p��g�:���ql�rk{�>\]�l�1��Qa�$�A�Su�|k��_���@�	��r���wB�ܮ���ӛ|��e$v�I��Ø΁��zX�f��Lvf�(3n�W� q{{�/����v�U�j��B��>�6�� cM���|�FQQ�%۬b���.mR�%��#k`��og
/R��npŽ���u[å��9J=�wJ����4`�a�z0&���#2I��PO��x&�0^�Q̷��v{i��OCb��]���*q,�(`ǧ#�Va���+���:I�3��+q��'����M��48'S����uj!��ܻ5�$��1���w�>�{r��3�e�gl�;r�>op^���5��9�z�k+,���wt����c�j�vjxk�� �m/V�x�3�+x���B���I3�mt:YX�D�+��E�9ـn�]���1���Û�ۢ�4�Ei�0��0ݍ�3s��û4�ĩ4-`Q�yű�;ڡE��{�kC�!��Fc�L�F��am�s��|C/MG�86(���݁t}[A݂��u�\�i��Oǟ*0io&u�s8��5_����wn�OT��}���@�SV�'k(׹
QgL�̛0la����k"cv2��&�S4o۝9��}���7Y��]�F�F<�c$%I�	]-��9˦�䜒���ր��f�뛐���[W(�;�-C�˗�ok���lRw$s���������J�  8̠��x�6u0G�b�U���^�٠6B<�]�f�͹1�^G�}���:����ݨ�ѝ63z��:9��tG���t�]��}���F|2u�͹h��I���أc�ٚF��l5���>�ʷ��omS~+1�KX��˴>����Qԓ�^#v^/����$3�Rњ�'#�LD
3��X8�˹f"��|{q��b���R/tAb��Y�鮽�d@��U�ܩ�J�4��{س7�[a�9H�M�wP��̾)U��D����.��Ѽ�a�����G.�S^闶�l�rnt�� ?���튷3M�E���3�ND�"�U�	�T���*6�񲞴��0�+h.h����#:t,^h�U�Q]u�\y�l��Yͨ��Ś;�-/���c(�9�m]�n�]fb�'	^]٥�oD�)��ZrM/�s:�xF�t��X3W
�e�4ٛ 7_=<�s��G���]c��� ���WV�.�!��a��ۇ��ѡ���l�h7����W(¯�t_P���Vv{[���V��&a`X�X0�����h���˹��J�J��ItN�gY2��s��}��4d�x�\��0�o)�ʰ"l����̑u�N�T���6>�{4���#� ^Ǆ�#ޟ��rO�V�7B���SM�v�o����2���D5P�N�9:�w4�]jꡌF�Cs{g�sC��������\o&�o-_VӅ��}�����w���]�AUoD��L���^C�=���,}�9sb\��y' ��Ҝ��]xݔ��]���G7�a��#*q�ܴ*V3Gm0�ٶ������㛌+��`�.�+S{�G݅�=��}E��{��I�Q<��y ��H��`�m����ܽ������os�6���L�D����ְS����y{�����W�G�J\=�f�.A�z%��Y�aM�&=�?��1XS�T��4	��vn#����	��ذv���h�n�k�unN靤��x蝇���A!��jޒ��8�)�"�� (x�1	��ݴ^�k�NAN]
�(�]��CxLygc[���� ��cr�#� ���h�����C�m�Ǆ���-t�u���'!�Y�5d[˾�~�}2��C���V�[5�6���_ԭ Pj]�����H!�!{�gWy�J$����`�^����ޝӎ��Uǜ�Շ��C:{$>��;��ыwն�1��w]c����3)�=X8�58#�RC�xu�DJ��2&!���j9��`�+�Kí:w9��}��}Ո���xe�=��ФǼ��~{2��E�����M�(�/�'+����0:��4e��h���!*�����J�0���{qt��qYڰ2����q���	K�9�s�>Vs��6�1��.��yz]Ӛ�=X��5���ck���f�"56r�k����ح�\ý7��!p㡄���dF�����of,��=|͔�7X[v�'�3S���;QRo�;�vˀ�<`3\�Ws�%����k7����4���N
�y�nv�:�e�f(�\Y�q��@mKZ&n��o��lރ����̸A���9���t`�Ջ8޺oV6f�vkN����#Ze��S�5U��u7��T���fؠ��E�/�`��{hC$5����N� �oI�M��j׳G:nwewhD<���Q���N :�Z�x9�[�pJ^PHV�q�0��M[hpbe�l���jy%'�.�����T��������X��Y��=�'*��>9U�7;/GvYf��;w���=��^p����L*w��,�a��u|z�eӑ^�v�t�;�w�Z�����5ݢoE��:z΀�H+��SV���sK�㍈�x��ç���G�j�v��\㥮��;�^j'v��4G���A���Z��!�%Y�E͓�h:qt�׾��]�9^��5���wdӝPtݲյ�6D�f�=�L�f��b����l2�Z�z�0���ы&9̉����+""�TY��&PT݆�<�_r��p`Z���P�s�8�yY�`��u�Kq���c]��J�Y���?ax*�^�i\���uG^6[@���j��5�q��gl7$�;U���9�t����e�v��^0�7q]
2\Y����n�5�����@�����Zq6��%wFM���"o��Jn�8v��eߖ�_,�^n�T� 0�A�Z�͇�5�Vq�eI�3`��5�Z�cr|�q�N��.�́��V�lusՑ�󙌤��c݌aF<m�z͓̲��a�å���7E�Z!S)L�epk�Í�4=�=� �=�.�dQ��'3�빋ow@���V�;��rw�DK..����w[�q�bJ
��y%�t��|8���SൻoB]I�����h�uM���("��;Fո Q��W50.����h�X^H0>�21ܷ�p��(��n�n��9�4�U��:sp�������>�f������	�<7J�V�'%��S�����)��p�A�6*\�L	rV-ʚ��eS��4e��9��C���bg6�K
����O�P�qf����fw$��9b{,�Ys46�7�ɹ�		�_;�c�� 3�v>ʻS�:s\�Q& 0isg��8�^��<����Ck���y7�����vt�7e*'7�1��W�˛���T&���;4<�_>Ҥ���.�����U�&r���7�� �����@+!$RH)AIT!
�!$"�!�Id� � +$����X
BE���@��d�"�T�$�P @P$�J��I		R*H
�,�H���$��!
��� �� �VIT$�VI$�@�a,�"���@� !	��+$�E$�R��HT!$YE!@�HE�d ���@�XB(@��%`P��X	V@!X�H,� P)!"�$R  �d��! Y!�T@�Y H� ,��IP��!$��%HA@!R H(R"� !m���A@?��BC�H@�s�����s{���������T7�l���-{Hм�F�ᵩ9Ze�	m���Y���BI��v����ٌ��N#���߸�ʷ�{�5=e�]M��V	���{��!:�XK���b�7&Ԙ�Ѷ��c���l
{)F_��p��3�<��`��#����95�J�@�w��7_���Z�,۳���IQ
Cٝ>3*4���d�ִ0^�PM��-�lK�U�`{����狯O|���FuȲ�s�'���g;�h��8�/6󉧏����{�j	|�(���������u�λY�	�i�.3�P�;���˭b�c�bC�{*�y�#��zp.�<��4�xP7�;��4'��Ik����[�`^�H����Պ�Ң�7�ĝ.��x]��=��3��2,G��=.9��LjCI\s�a���|��ۜ�oqO��7τ��f�un��+��������q����ڻ�3}�pY���k�CՕ��;��K�9u~�÷�+��X�{*�}|�����o��^��br��x��e=�K�1��F���vt�����j��݌}rk��xݐ�Y��qzp�O
�������qq��0�d����0��H6�Q3�>ɋ��S�����4UںS �.�١��#�Z����>�[G�!Ga��Dx�f�p֌���sg��T�0�v�a�$�=pS���^��dӚϙ��c^=Dm9�n__W������x�N����R�s�2����c���s��Q�V��kc[��I"֤\L�O/y��=��Ҥܥyn�.�方v71{*1o-��}z�����W���R�'$!m͋:�SNlFBI;�1�!���1���tM2�z��97����)��s�;G��Z�����8�-g��`qa��ڭ�K��Oz��M��(����/S���_v,�B��<���ޝ0듰�▊�Y�M൤�R��T�]��4LRk��W�ga�T�W���o`�M����as}��^i����t+�z�7����W{��==� ����~Ђ�kΞ��w�{�J	K������ ��'C«���H{�S~��{����ӣ�E��Y��ݏ��x��*Z��W���5��y�[��OpR��b8901޹6sէ64S�؇4t̐���i��)���^�߻����/��V�v��3��+ć�d��zj����z��T�k5v@�}���F .{��H�wRd�����
}I9��1��+��/�n���kL���?{�4lw`�֎�~�.�3�����$@{ݷ�^»�>�O{Tپ{)�U�;��9�v���Ѿ�{ع/6 �����6v'����|D���s�b˰�q�עH/�q�M成�d%�M�Qٹhj��g��w	[��ռF^�}��7GQ�;��쭾B0'�K�d��Z�,��{��Α�N�L���h-m����l3�Q|�eP<�����ܵe�h��B��w���n��FF�&��(���6N�.�nkj�S<��;�O%ٮ�c�o�Ƿ�0���������������4���+�I��k�#�O#�sKzv���<���a���+��ֽS~d�}�:t]�Wځ��:N���C7E[�Fի�zq�2���,'in��G�E�_c�l+;�t�©Vz�����zyw��vp78
��kdr\xoUͯT�ۙTSV�H^M�����=��vÝ��6m�И�����M�{�N��GjЍ�]2q-+2����k[� �ۉ3Y-�8h[�R��X�3ccS�J�ht�ǯ��.��-y��F��Ƿ~�HA���n�����WW�_���=�R�
M^�}.lE?��!�Wq��6*�4�ohH{�`�W�O\W�Ҽ��e��t���{z�r���:�;�5��@����R���M�q�f23�=��Ep�9��^9�w\݋k��Ei�0��A�-�-,�!>#�r���������V�bC�̖V*��
P��F�9����� Yj3$h�)�����G;�-���>�>$Z-��es7�1��␾]]������Jp<|N��S�����mk��{Ц�A|�.N�m2����g�.�V�q�]m1le/&u��(�L�Fl�`��׳��7�4��ޒ*�@�(XvR~��:����L<7D�gfڄ<��!:z���I3�C/q�����)�Zm�58��g�����z��fzw 5��ˊ�x/
���z �A�����`�q���^�pXy��Рm��$�ۢ�tm0`�H��Ƃ�Y���}�ӷ�skZka�w�:����V��6��w�wё9�;]�-���fOG�ܒw}0/U^:VAq{'������ͳ���p*lyӰ2�X�ש�_t;�P�ޗ|<��ﶗq�Zt�m�p�N��4n�7o�(��ȉ�F�ܗCz��l��ע�Č�m�ĄЬ"�٪6��q��u��?��ݩջ��(�@ �
i6�fޝ��%�2�+śgт�_C��T�X�/a�������y���U��Ox�M
��v�!/z���1�{�����E��·��dzw�:�2A�R8f��
fl�d��^��ߥg�&��n����7e�6���U�np}9��=�$��}��K7�^�ֶ��7u���nخ,\ҝ� �,���	r�u��t�U�~��ⷝ����=2z�>퓸������ ��u��|�F��d�]����z�y�!�x��p~HN�Պ���׉xtO�gg��\��%ឯK���H��"	�S2G�",�S��gxÔE�Uթ�+TN���3��R��
����Tn�l��j�ʋVM@���λ��W[Ƌ�D�վ���aI#�ݕt�'W�b��:޲j�9�o`:Qe�h�9i�s`~��e�C��ǗO6I��S2����5Ut�zzD���5gr�����7;<�Pỵ��Z���a��X_�ژ���iY���<8w�n{U�}�<"VUE8��O�n�]Z�;�(I�m$t�Ǐ����F�������sW���{��5�K�h�n�W���1�o�E�q�*��0�\�_�N�~\a3ܻު��=�Q�h��3�J,}L
k�*x%]X{5��9����,���C����|��{����:�Q�nEz�%�n˺���&7XlG�g�z1�%u�x��f���n�N�{'���vD�w{r�ƌ��ݐ��b"��h�[%�kgCH58�Ղb���Y<Wv�n��	K�x%ׅ��Jf�8��FP��<o�v&z;����]�n���n�%R~��n)�=���R/r��Iu�=th�=�ay�Ľ�|w::k��ĺ�y��(K;�ཁ��qjE�{��76w��!��]�}�.����;����;<x9�԰������P�W�}����Vг�ۓ�����<�����<�no,L������Gi�[�Hɼ5zL��e� F�'yO 9{��7��zp�=��74�9{S��<��"}������.�� �P�0Z�Ldl�<ft˪y����[��x�{���m�Y!��&���b�����Ǯq�B�x�a5�M��������"����ofٵ�i���83Rb��Ĵg|�Rt�EC̬�e�w������7�Dē=��w��)W�Ż�6ݧ�MiL4D���|t?]dt��v�F	
��ս�L0`F�<v4��bkr�=��v��#s�b[���x���ۀ�b��������X�Z���le��1�����kS�O��"���GQ�]�y�H�6&73���n^��ئ�P�v��H����n�N�K�n�N�N�m��^�,�ng�H��9���{�74{|�j���.v��c�'{�`4e�>��΋���nڨ�&3�Fn�>��v﷏�(���y^�eɣ�b�����I�7�(����A�Z�3��g���v�\S�K͞]<��������j��b��(�l�]�7UF=���"GYъ*�'V�-H\�u�3�L[x/b���~>��}8�w_h���ka�/$L�	糪�*����eFSS�nٛRy��s���"5_a}Vv�ۯ��7]C.2g(ޱ��������A����^J@�SE��7��W�6�� ��S���ޫӱ�u���0��|kHe��D�N�k�#�����p��{��@��hq��os�/�2$�F�����ݾ�bzc�jձ4�������l���9�q�]��UR������7v��~�=���U�
p�;jo_n��+bn{��w�)|jʀ�g(у@�r�t�H��IN�e]��V��p����
�Q��}�ܡ��w/+�$��v�؟>�ЍEz�8;��i����ǩ�Sމ.�]9���(��!�t���f,�د�݆[����H�%��q3�Q�P�������2��j�:D�4Q(T<JpNM��'�S�n�&�U��]�z�w�@`�~�Y�tܣ7�A���BI������^�Z�$}�]�;Z�D�tk�����UE���oi�Ѻ&�C����8Ŷ��}n��b楤{��%���GQ񧠏d��:�f��j=u/7�-�Oo��R}��.ؽǕu3�Ԍ��q�m���=����FԘF�'�_��=��z��p{��Ps�SP�o���v�&/���;s����>�.�������u힣�_)4eǽ٫�s��>�{�Aջ�M;��>�c��z�0�G�j/>��3�+��ya;�F΃MP73[���h%��r�7k`�s�&R�X���~�7�V�%&>��+#^�$f��Q�;wK�++E��Xsqs\�8=��9�P�;�Al������S	w9��v�o|���:���ɴ����ir�r��n?ik��c�Cb�+:s�w5�}���R��2�7ڏn�P=�-Y��^o&܄Q��_1�>;�Xw=�y�u�ݜz���j��ž�re�I��S�$7�w�x7nu
g�a�w��T;�"d�V��j�{}X��{i��3���cWfɌU����m"��K��Nܝj�/սs�rf����3F̝S��C�{!�B�� ���a`S�����%б�p<�(��3�G�ދ��Ӵ���@��7�{(�B�z�o@���i��Jug�?$�'�7��x,�s�Gڦv�9��`��p�v\3}��ԩ�]S-���;���#Ȏ���e_C�L��� ޗ���~=�-y��V�L��}_���\�h?=/*C7(�Z޶��\��Q=N�{��w{C������h�R�F4�ůK�=��՚3Z�o�Ӿ5�q�}o�ay9���^�@�9g��t�y��Z���������3W����wq��E`J6��U��mN:��ѱ*�Ul�r���#j胳s��
C��v��\Q�T��Z��4�����w���!%Fs[�~���,��0z�딝:�����*\�����P�-{p�[��4�ɸ��̧���E�wm�9{U'y�r� ~�^��sg��������/5��@Z�1�V�	�X�n�·���o3sl�V�o5��=�l�U\�*�)�O1�sی������zewt!��{������<�����v���@�T{�.�x>��Q@�Q��0j	7.����v��D+0e�p'|�l�r��K�(ArY��+S"ړO��ݜ*$=�4ة؍�EY��7�{�����c0�xs�s}�T	3�}�j&#Țk/u�+4����&�:nf�-�:8]�zO!����З�9-�=���qs��(�;�Ay�]o��mYm]i�#F��C2aCח)9���Q��=ܼ3�WA���N烒5-|���V��K����l0���Oo�*��(l�(�^��=����Yqf��3c6�T`��cr���7��>��
�dg���I����cט*^�Z1�{E���A�s�
[L+�z��]�<������qC<�Ʒ$/L+p���c�%:��^���wW��nv����n(D�ᩃ%PVe������{J>��a�z�����{���C�L7��#�M`��������V�M<k?391���'����ۗ\l7_��yu�vB1�v��_��ޛ�^�1y�2L�a�_N��n�~�F1|��%)��9gO{V@`�.{��ٝ�$Ux�۰��M�x�n��Y��7�=���/��jl�_�&��ӓ�%^���ɓʗ�-N�)cv0���	�=[@�dܬ5F�;�b�P��.������m�K��T�ڰ��\�wV(���;�#o$������{��&v�˶�nD�o�w��[�X�F9e�̫ڄecx �^x�h���u.Õ�/��{�7�Z١7^�*����j�[$��C|m3|}X���y.���Iy���	ӡ���᫝Ȋ��*X�l�i^x޻�l�;;+���Yk׆?5[�*Q�0��&��q�o\�s%�^�;�v��vp�R�w@�DV�u2�̕�L��eN����ѻ:$^����'2�-����Յa�ۉ)�{|��w�5�v��jΪ�+h�d�X�3vq�^�{o{��%=�|̴	������ۭ!�>G��#�w�;7}�}�N�z�@����_t�%����ע�:���y�R��۞��s���M�{��
�'h�1/ U�(\Dn��U���aJ<�J;��M�����v� �;�9���wI�\����ٴ#rK�-�w��+��§��qIb���w�YfY�����w�����&S�3RN�Z��x���ʱ�G�lV���Ӧ]4})���7lٞ�=�c�(sA��ɐp'_9lT�.N�6)��[�ss�MȀV׫RN�ڻE��,��q��z����t;�-�n	�M��C ���;��w��Ӟ��3~��{����@�$�BI=�}���6�FB��î`�^rs`Ds���n�y_k�k�6�Ÿ,�<l�\U"򻘷(�=:�Yv���@cv�v,��h�2t�����]����CU�Ok�\�h�2���7MO6�)-^\�h;s[x �"�:�O+���Z���m�j6N��r�v�;��λu�K��n���>����$i�}��<��p�<v�ћ)7�c���qT��k���La랣M��;z���sk�˻k�<�&�6�h�7[X��l;"��nC��{���r�x��݂+f����N݃e�C�ŀ��3ӎ�p�u
q �X�`�|!̸e�!��5�櫆�%�"�y{;ҙݒ�V�/�������}5ږ�甹��=���b��R6ڷ<qF����ok1���x�)�0��:G
1ū�YNWrcv4�Ga�qr�ZÞ��u���O��t�w^mi�Aa.'p`퍨�'=���Ɏna�od���Wm��f^ٻm=y��<O'��;�A�[$�c�丄�ݎ�R�q�p�#�l�ās�]����k��ۣnn�yw�#k3xٻu�s�յ�50��ݸ�vGo^�`�x��Ƴ]�n��<��ު�P��m8��r'�WA1�-�r��rvS�v�0�pN;2��a8b�ݞލ��=���6��n;5�J�!3��p�֕#]r���n@�#�'�7JM�8�:}��`�]Qpʷ
f���t��G�<n۴�5�vwns�;�h:M���b�&M���h��X���ںk����E���Yzq�n=�Tuv��v9n��ۅ�n��&������9I55h��z�T��;�����b�2��o!\���Ej���b �zNT��&�f,�;[����[�:�k�	�Gm�_tE��A�S@�Uv7x���r[6��:�5��m�z۴Nx�NV&��]������q��[st�۶]\s���ˋ<zħ=��pxz^om��9��^�z���+ǎ(�z}iywm��ƳĜe���7n�$����$��[ ��F9:ۘxG/d��n�]֧�u�E�1��jScZ6z��9�����⦊����.7\����.v6u�iܸ;V��H;]���Y�6��q;/Ogw/hSpp�Ir�{���`�O]��j;<�W[V{Zd�3�����:��s݊�^3�!ڷc:�ݷ�4��{Xq\�Ӻ�on�-qڳ���֪t�vY�34q��n���.��Nx�ź�ݛ��V�u�ݫ��^�۵��y�<��\3�O�8�ۈj�t׶���t�q!ƻ9����wW�[���[Wc�.z���װ㞞oB=��������Q�5����jK��,��i;d�[�ݹk�d;&�xq��.��\N�b4򀮴��K�e��A9��sj�l�v(�<�l�0���.�qcg��v�q6c�l��g��z�����ƶw�7N����Ҝ��+�`�'��^ۓ�͜��&wg��6�G���Y,���]���ε�(� �x�j]��xϬ�y�;'<���q=���)���۶��t<ri�rv��㣶�zk�'�5�Y{�fl�t��<�:�]{�����A������c0�y{Y�Z�#���z����n��G�x��m8�[�&��O��$�Z:Ku�&X8�J]=�v��&��zz�޸�{q�p��:��b�u��v�+����.�^�:`oT�}u��f��ۺ��ۮ��N��7�c�ք��n��7=n2�y�Y��g��9�՞
���q��Kno'���\��|) ��GJ��0�<���=�ɲ�h��vnt��1n+��\�vʾi6{;tn,Fn^{rh�C^��i�v�ή۷,m<u�,��u��m�8���/B��y^x�i��ܻ�u��h��1�k�pۡ��� c�����ͨ{U���+�9��s'+쎦����/[���\���n�W`2��ݱpLa�|
�����m��C�7���@-�{>뭂���-�]���x;Aچ�cuL��Y�\js�og7d޼�aی^�dz�^Ik�an��2s���Q"z�.;B外�^��z/Y�O�%v����z�F�c�2&Ѯ-�:vy�nb��6�dr�n�n|�;v�{6%$x��]��*���bZ%Ǟ.,�S���׬�{$��۹۴�\�e3�zĶ�x��ԣkm��]����m۵����m=իO&���I���v�t['k�{Gn<s�M���j�v�mv]�vp\g�x4��=��z{�u�m��s���mЃm�k�P�9ָ�rmu�JHW/3����t�۴x���Sh��О�JN2+�:����m;��n�m�e�wn��ɬ�]�v���=v��@ݓz��r��m���M���4���/���=���s�^K-��sw&r����Z�y�`�{9��7���3�n�6[/-t����|���A�<sk��U�d����ZV���7R7`�x2��c����\[�^M�e;��y]�n�m�f�A\�M�ޥ��G:�	]rv��˸i��qh���5z�v��![��Dq�a�:9�Ýv{�&t	�]�!6�웮�ݓ�V�Ӱ����fN�8S��Y���kIpe\�Z�U4<�룳��`)��a{�{nڣ\s]�s��;K����n|r�!]b�e���_N���!,k�[��8|��s��v���1p\��q۲�w�y5��՛�v�rv�=ha� eu�s�=k�ϴ=�ku��]9�eK:�ݺL�l�3�@��.�'Ը&8��p���au��<�[�;��8��v(�c�:�i�irӶ<�v��W���S�������`�����8j��ek��v��t�h��;Ύ/]�1H,m�V$��n1LS���8��=��`�!�� �v�t�m�ˮܒ5��A�S��u9v�tvC�1ϋ��0�m���z"�^�_��j���t��̩Lz�W��[3����m�^�,Ml��FL�lPF:���͛GF�L���e�gXb��Nm�l7>x�����HqǱ%���$�Ӫ#�vr׋W���c���n��� {MBL�V,��u��v�uÓ
z���m��.�Y�z���$�z�9Fm�i����vCgS�cg\CO�����B�nKͮv�t-@�e^pb��4��q��]ڎ�43��)�
C�+r�`c��Jg�\K�v7�2��r�a�8��������{����yW��V��m����i\f�G��6D�ce燥zg����ӷ˚�u�+�A6�Vn�j瀺LQ��K�P���x����� �x���;k;ձ'F�8=��c���׷+�0s��[��[����a��r{ny���X�s��e��z5���|SA����lV$�Ǯ��L���vƸX1���^O��V��+�\�v��P�s�]��5�%��qn�P����e680�,�G]��>�.�v��v�n.ζ4n�uì!���R�y���g�+���wb$�N�����j�Nc�u�b�m!�����n�9���e{Y��l^9�+���6�GS6:�ײ�t���ꡋHn3l�R�F�DU�=�j��Vz�#۞��1[i㸑�n{��N���.)9qc��^�keCs��W]/,t��uO]�jm������v��&��Sc�q��:�v�ە%|�nn�� 2ms\&��f�$y��l�`�6�mn���kl0�ٔcN�{����:�c��	�'k[��6���̮��^���n�����)����8�[�ݖd�gpv뮸���ϭ��]]}{-�v:�6=��#�q��:vn#��HXG��U�C�:�n��z�X|s.Kq��-�#ywf:⽈�	�;%v�=u�T���q�f�⛌������u�a
�����>�`�9��[�^��\�hz���q=9ź�퓤���oO:�Oc�K���� �h��,��+�s$�$������r�ۄ���[�lW��M�E;&��q��q�L��۸Z ��[�uᑙ�6^�͎�s��4���Ú�`�%q:㕂6�O[U�=s�nT�P���p�,��4�ل����C0v�ۄ������b��Ǵ��9]����쐽l�غ��mCu-�li��&�g�y�>/l�³����sٞ��ƶ���\��EǍn�lh����׃��n�9���aW���l�n�/l��g�8��bc<�[9�(3�")��͓Zk��Ϯr��5tnw��:��;EC�#ˬ4��٦J2s��s��ӹ�����3��wd��Q�l�lm�q+�f���aN�s��0X�'W3ւ{���=�hq��˵^y�n�>�>wt�v��;�
c���]Zf��>����u7����<G�n���ogh'p�t=a ��3���prg���dw��5vhos��F��N�ݦ܃�\n������\�Y�8SjQ�pj�s��ڋXؽ����(�آqsk�7�l`���z�C����!0-�8Ź�DM	ϒ|�h4��˒��z�[q�Mڥ��f;Mv6ktΎ���@w�q����)�;��"n��2�{Y��P��v�)f��#��6[v-\j��ӻ[b�p�� �h�[�g�V흷;5nh�x��U�j%��Cτ�s]�ێ&E���zvh.�q���i����J�۝-۔��G���d�>w��������D���2���J�x���Z|�ţV�q�x{cOn+�9��kcK�գVe��&Q��ۣ<u���)�t Ej�;�����Sn�I���T� :���wu�Ɨ��ʕ#�n99��\�p�����I<\����6+��#\�hg��ݹܓ�����t�\Ї^�%̴U��h�5�qT�^-��B��>�e����{o(�+|As*c�DE��q���Z"�.	�V��a��4j��\�2�R�  ���Rңir�Ah�*�[jːp�G��w���cll�J6��J԰U2�Q�DTFܶc��A*U�2��[lTqYKB�aLs
ZT�iY\,�%�e[\jָ\�����\ˍƈ*9�#U�-��c��)h%��m̕UVf��qneq3+�N;�ݎ�&G�S�ݑA��Gc����������ܥl��4K�R�&��q��9ɷ q����ݳ��e��e�2Z�V��D�G,�e+�+�L�+s0DTƵ*"��\���������UU[jU������h��b��ѴlQ+UU��5�*YLa�A0�q�V�-�°J�r��,PbV��9\�Un8cE���q�5���[kYQL��eR�Ls	q[AL����n5s2�cLLr)�1UR-J�e�Tq����bTD�V��-2�L[DE+U�������n�z��V�M[���n���v�Q��..x�;N��S۷�L�$(1���@�y{v�?___KVs�zj����".�W1l�u��g���ؗb���cN75��5���8v3��z$�ۥ��=z�v8���	#�s�z듭����|�����;�^���z�j���n��m�:nxst��m���P2��l�����B�n�����r�z-G�9��힐���	b��v����N�Go&�:�zz��K����ɻ[��X�a���v�����I��3�RfWF��.S�88�b�>��WH��X���ڹo\Q�u�؎8�3'l��ruxꖗ�lm�:�}6���ݭ!�u`T�&Hwmmm�tGm�>������8�m/i��|�8�lq�=��)��u�����p�]Fs�
X#�˱�x��EWZ���1�ޮ�� �m�����I�k���`7n�c�'�݁P�!(k��pYA!�,�=�55�xʇ-mɮ�Ļ����m���J{c�ۍ/E�qv�v�	qpt������k�ّ������6=fwU�Do+�H� ��Ab3��K�:���v�:Q(U���>^gC��:ݹ����:���9��:���d뭬�� Z9�k�fзm�k�=�r��+���-�i;Y�t$W#���ki���mმ����@$�[�N�Y���#�7ٹ���pt�lv�ں���61���Y��ǵn�v�ez5����6��qĝ�u�^��v��pr����w��u�=���/�q��]<t77\n۵�3Y{.�Ļ]2������:�[c�ͳ�\;C��k�[��s��9̰v�u�^�~�u�>��H;&�h��{@��C����X춫�=.�<ݼt�lnP��rX�Ah�<҆9x3��I��u�8�:����n���ܷ3�c���$l�m�X�^ݼ�j��H�un�ծ|ώ���y�]Yd�k����{ӹ�:�W��s�y;{l��۟eC�*nw=�{d=��(��s+e1U�̃2����8�2��'ev}����'m�''rg��۷�;v���ܠ��vvy�=���x���ʛd�)�������q�v/g�x;�xy�l��U\U�8a��S���)�\�Z�1�r�q-�4q;	����L�d�2��n����?��
	�� �j����͚��۸�os#3,���qS7��Gx�^n�
����P�����Ol�gŎ݄j�����wEt�$����@�A��p'Ǖ����|��;[���J��҆Bb8����I �ʸ�A.$Vk����n�F��Ux�|x�\�j	�I��=���R"�8[�'ź�D�E���>'�]}]�%����C}39U^7V�h��&b׎�ː�9W};�6V�؁�����y�@��*�	����cb$wLN��x��Q!�^p��i�b�8�f����v�E͓��\X-�!0�]��l��n �%ޛ�ʯE����>$_]�W�wv����N�A$����F�9dB�a��5@�eu
&�N�lV�yB9�Cu���طw$kֈ���xns]�{�����T�T�F�<y�"Vo ���j���22d����x��]}��XȝowgI$�[W�^��Q�M�]>��&���@�J.!DI�Ӳ�>z�*��0v�ӌp��	��p$����"jU�6�8q\뮆-s����o��"A�Wr�$�뾡@��ު�d�5D�Ƿe��V��i$6L��ۚ$�ޚ%�"{*I�� I ]uuW� �nf�Q�࣯����`̈́�"'��<�v�c�ٳۧ��ET��y�Y�i�oU�QN���a��M�S��۹��u�� �}ٛ�F뢜��Q�ݴY�6��3n����l�YL��0��wo�� �'w�{i����	��eW��ު��<X�e�D�9!��r�0��0�9;�=��5�|O��Z��dU���NaR��G�'d�V�����nɝy1�⹥���s�l��gF}�ދ|�G���#`F-��ݓ��qs>5�]4s7������a��(�����8M#�N��*�Vg$z/z���GvwP�|���(ee^O0�-��`&�^U HR�a��b!������$���sŜq�3yJ�<M��UH���I���"/�Q�J��q���D����B|�#���[٧UU�8Ks!�k�k0�z�Լ��}|����&E a�FMmuN�oMxH<^�Sd&�*r�����Pر{��	0���x�܀Ɍ̓�v�� ���׉�/n=��k_7�/�M�-��..	f�t�$Y{r��&"]jt��3�� ��t� ���Ď�v�-��l� *�g.�H2Ӂ��b'�_MI#�ۉ#+��¥�\j�ር���E�Yő�w��|��c/4����Ŗ{�g�si �����	��ݻ�E8�=�ږKo�$5���XC:X6!ln3~���ֶ4	��QDCE�f;,2�����a�{P��$9���A���NWWUxӉ���Wr���� �;a&�DP���9��v��P�n�60\���l�v�>?�"m8�o2�����`�FT�U�[��{W���*����g�_[��-�R&|v����������O.$��=�D�[�g	�j���lc�����X`�b�<r�@d�r��h�1¹lwC��'ě/.C2����\��bfJNm�R��r%�W�-=���A�S�TA{�F6�FR�dY$1{>g����q�l� *�97��$���t���1�ni�u� ��9�@�.�z��Un��wl�x��v��3T���ٽ���P��2�5���\豾{�|�eG�hl]����S���>C˂�Q�������ϓ����ﾶXJ�s�����/A�<�n��#�<�[gv��g��"޽�����t�Ӹ��RO1�n��,cڎ�ѹOBqk��/'�:(�x�OS��ۦv��3��>�y%��x��yz|Y<�5[<����Cl�dB�t�{Drv:�Gl�6&�9��8�mj��<xѨ:Vڈ
�v�����m��3t��K�Nm�wV	������\�;u�P��$�T���֞(����q��]�.�ڶ�|ߟ�4/ڱ�2^\�A��H�����������5U!�HS�T	�T��a�4L�8���u@�Qª=G%�	�Eh��.�:��.�z�x��N�u�,a&k�2�Ɯy6�(��2�ͺ�<O��oH�HS�ˬ*�C��F�z��h	﷪�NE�Ћ�lB� �˼��Tsb��KzVa>��hQ�z�	�쑶��"hE̓P(���P��Kd�~!��n�t�>6_d�5�X�Å��jh���I{�TA���%�3P;L�M�n�&"��ƼMٷP�=��d0��<n\p�z��68�;���~��m���#x�M�/{��$���D��u���WuP$ם�D�oh�)��L��,��%�}c9��o�m�4��\_Z�p��b�L��ݴ	�"�cY�ۜ�܌���؅��լ�n��x��A�F0l��z�V7v�^��ʪ$����@�|t��츭[c,����b�gC	Â`7	�P��uD�O��ω#ф�Bک�rҗZ#�;��$�=9,��zh�Kl�r��wgh�$�W\���D�|	ɮ��*2���F���������[���Yr$���xS����oFu
~8;���`�� ^~��Q�����P�K���B!	�%y	�$o�]��;L�'=3���/ܻx������m���.���ʯ�,�ȐI#&��Q��9���13g��gU�:�|϶ޫM&ߛ��X��v���+�N�~?������$r�$�ޯ�љ`�D������@anI�
0)��|d��F�vUfk"���eh���m��z �=��RV��t_[̒��O��XQꝎ�1S3W�x6������]������o�"1�C([�yN� `�5���	5�U�J�I��8����g�f�%���$�ޚ �n����hF�ȸ�Q��S�ȅ=�z4J%�L��{uD����@�������ҹ��I�ڢA7}�T�ى�kg�����j����5��9�G#k�x���Iv�ku��� �0�1��K�,@,@lB�����$���$]����} ���}^s��@�����!&kv��	$��F�0Q=l�A=7yB����6 >�\Q���u���y&���x��EQ�Y�^$��t�$9V�b����-��F�_U	���Ha^Q�JP-�l3�N��N�w_N]���MM�wMN�`��5�&:������k�������P3�#O��#%I{|��v@�S��Z߶��z�P����y�ꈟ]��E�ga�{?뉞�&j��0�bÈ��}�T	$�y�q�2���h\�C�گV�oUO��,(̬��W�%��L��}�����p�Z�ۜ��]h��F{��A���kn}��W����\ϡ�`�[d��̺�'o7��$�q=�;WY3{�38I9y�B�SI_X�X��B�<r�Y.#���m��'&�$2�z�N�!���l�3�N$c��x7�"�C���5#�憎�/rY ����W-FX�j��M�oU	���%���7 �m��5S�"bl]��{z�$����x�Or$�@�꽪����#�v�:L(��m��}� �M�Up�;����}}�u^$x��Od�U&n
�!_r{_�D��K��->�X������y�^���Oq�$�!�4;�.�b��N�P�}���lo6��'V��z��E�"!Ya"�0�����1�mӻ%���]��u����lk"ip�u�c�ڇ�{I�Z�Ev�z��+�g�u��cg����0��{.�O�����:KdR�c����2y.sB�$wn��*t��H��l)�44��m�q-m���\�h5À����nF1�%��YF��M�v۳-B��S��&��ny/l�3ha�@k�
l�f��Ȭf�C�'7JK���scl�ڪ�}r�#������X+�9�q���˪'����Kɾ��YL�Ge��$�e�O�fq���D�h��ܺNt�U\�P�U�=�ď��� ~�?v1&�^�a�g<˖��Ǡ1��Tx���3�I����H5#3�/�zwĂ|l��	���P�ڡ��H�I������sI����"�Y������^��k/
#]K$�&����Pp��(�Be��	:���lI�̌����sO�\�H�O��z����b뚞�0�N�e5�e�"�kq�׳�j��9��%�N�=��1[,�/2O��
�2[E���$0N��P�A���o�ErhL�t�t	��o�W��^�Rl@A��Uy���|����k�ˌ)^�P�������)�v�Ѽ�xz.��Phf��6�@�O��J�<:��nn�{����J*��R�k(�g3��}TI"�7��$�A���� \
0��`��]Q$�f�� ������y��|��Mx�}��@KE_c���B���b�h��wO�v��	��U�A'ܺ޵s����	�]TDFb�a2�(`�;[}B�&�ܖ�&��ɽ��!EV�UI���H$�{�����/Lo#��m�B�Nܾ����pgJ�s�B��X㣳��'q�l[_����2T��[��y�3S{U����I��zcGd��'}���@�2���¼�
�2[M9Lnϙ<y�ճ��2﫨�H'o���H$/r�ac{I�U��7IT�)C0�i�U�S��|x����he��
�����=)�W<��Д�M�U�hI�֗�[�sǢ������l<3��]+��}�d�E;���j1\���D�=����r����Ր�8f��:O��9v�]uZh�Ŏ�,��[����L�͊�h�ҹ�8�;�r9Y����_��xi�Y.z亸��niڧ�Dlbt��s9S<�J���mo�o`���;!^���=��#xÅt$i�m���>��
^��4`�1~R��0xO=#R����ܯ9�̾�b凣����f�1��\^�LY/^Hf�:�Zݰ�=�Ɵ{-u���:g\�=D��̕�Y:5�!��b��E=�eY�&Eԃ�la����<��;���\��ۢ�0�t3��`�Wj�V/������C7k8�������+2)�Y`����lg��ܦ��0�@��\֢ M�
�gf������Bʛ�D�(A�ە_{��I��.�y�u��nn#2���� ���ov
f��!�}�;���|��J5���y�OLd�u��uQ��A�sN�=Ğ�s��A��=��|-��m�w��?7Ol�n%��$YZ���� $�3�{��3S�1���iG������Gi�P��=)j[�	W�3}3T�\��\�,�Pm:/n=w��ύ{˧Q������ͽ�W
wr�����&�Vɚ3T��s���y/8:��l�<8�|E<Ӥo��|��t��4���rS�W�	gL����y�Ea�+�jΚ�D������ߦ���$|S�9���\n�J�j��[��9L3)��&-�bX�(յ(�F�kUK��`ᖹb����+,��aRZթS0���TZ���ELJɍB�R���i���4�jX�WTQ338Ь�\s������3.6��T������Ō@��̮.2�eJ��/�6��<��r�.��x+e��aB�ѥDs,ĩT��⣖��[El3,Q���+f\�T��[�J��ʋ��
��ZQUs1,�����[�!`��ѱ)m�-��-�J�h�9V�Ɩ�X��j���k���s.	�e�(��
`���2�kD*��
��KS)*�����rZ)KDlm�.[��k-+F�������
���F����Q
�kFڋAĶеƘ%��8�pcv�'��7�J%Q��`�%E�U-q���2��*�4Km�R�ũrՆ,Y[n\T�U�.�kJPl�R�*+U����TV��e�ť�(�#JX�ۅ �HEfw+��#/7�����O�g�GكP�
wG~���ʏ��fπ�����"H>͛��
��ĵXn��H��ڠNSE^�c���B�N]�������� ���[���A 
7�����O͎Q6�7�gn�QH�d�:�2��l[��Whr�]/e�'c'!u�sɀ��nv�a�*�]{w�@���%�A#:o�����c����+뼪�^d��:!6؀�p`�4f�:���w�\/�ٸKy�D�H:^�Iٳ}U�M����ɮU\�s
�(�Ɇ�92cv'ă�7�(��p֫į*��s�<I�� I9�}TL�+��PɀKm*����ꭥ�!�X����2H&�o��$��u �}��A��.�����Py��Z���	���^zC��/<W/�^8��c�$��O�&��2Vm��9J��'qX��;Ƌ���B�e�!�d�$m���C���(�I�N��$�v��Q ��ِON7���.&x��7 ��	���nݭp�����qq[��pC��6�mG��~�Ǡ1��<��I9s}T|A��wU�dnᭋjk�}7�^$�n�i�q!�����
0B}�v5��z���@H���O�y�T�P�(I@��ݦGc���`&�%�x�NuD����A2�J��t7r�4m@���%���,�"VVh	�3��!Q�F׎-d��5"�'�}�T��a��af�( �>�캠fi{�A+@X5i��Ө �+��N�vL�;�b�J�|!��W�'�y�B�'����y �{z����3�H��:o��B��,�h��fex�*w�z������=�>c������}"|6M�N�v���c�.��]Ŋh܊�$��=hv�zY5��Ss��)����z�ҥ�,�^^��;\��L�9���pki�n�8��5�3��wg
��뛆�m(]v�[-&zv�̓*n�&�!�c:��7N�ɶ��ۓ�����銴vc.�jy����\Z�\`��۱�ɮ �X��՟9�vz��.V��Y���h��{uN���i��;�_G��QI�{uƻtYnHE�]vZ��u�Z�n5�6{\X����P�a��Z> �Y1g��uGĝ�ޚ>#�D�˜����!�Ux��n����"���D 8�ې�]���N�Wi�w9�|H���A �����p�sв���i��m���!�ݻ�O��Ւ�&n���'i�}�O�_wMN��z�h��jn" Te�q��{�p��=�	5}"�>�Ց��N�T��t�]�ܒfUQ"��@I@d�N�<�Y#g�*�kC6=��M[��D�9Y>`�����"��y�t���}�������x�WX�Dv�<�v��P��ޫ��/L�V%۶����6��7����0xW{4f�^�����_K��{bad���TH$;Y,�p���;��^�aek����*I��![���̞P{	
����#.'�/�Z���ؕ��^+F뤶�3����8:��{�u�z�r]�oy���~$r�ȒNO_O���gv0�.�����f	��B��v�̑�w�D	�z-t��1V(�;y,NO_W��m����a�k��Wm��A��H<u�ӷ�(������}j�&���O�m@M�D�8���NnwM�<1wV��o	�D�|MN^�I��BC���Q��`B",d SM��m¥�s�Yz�ug$�ݥ�c�v�ݻ�]�Yݨ�/xAPP0[�św!��o(
��7��9p��H��[�$�l�ܰ@'g/��i_C)C�)�j���Gw�SKT=yXr� �{W�(�/3z��g��AWta�^t��R� �C�P�3 �n]Q�'�w7��O��.�)ݗ�A����G�s�n�y��|-��7h�f�t�n�>|��{;LI^7�P�d��oD�/����������m^��o3嬨=-|����T��5="E�x�HekݯP>$n��P$�����ehLW[Pb2VϢ��t�Q����N	�!����`6v�@pˁa�Zp���FM�7��E F����F�,y�(�7� �x���V�ϑz�9漴�;e�-��n������@���	���D@/C��ޣ�FvwMx�I�-���Y�is.1M�?��
!����Τўw��n]-�xI�Ϥ�H���}�1K�u��}���q��*�y��}���ְ+_o�=��H]��}�U'<<���"�U��bEf��:����vq ���|�?2m G� G��S_�8��}����7����%O����:�Y:ʏuvl��� A�%��-��8�A�O�}ْ�"�%�A���A ߟ������l`W���wI���O�#z����#���Һ
�qr��l{��Ԝ�o�Y��^�߼a����taS�6�݃'_=u�%/�1$T\Eu�C���^�4�x��~J�C�����Ԃç�r���8��0�y��0�׿��$��ID+�y�|(��[�Ge��Ͼ���}3߸u�T��_��=�Ct�B���>��|(������v�[�u,J��v�4=�%���xͱ�\7��nY�=%�^�n�!]�J%1ٿC��11�|G������YFJ�_/�{���B��T������!�aXkǻ��vI�����:�Y:2�Q���结��@�y��6�"�D@.���O�:ߤ���Qy��8��ӫ�Z�]'��B���������H,�<��}�,�ϼ���D���n�$mh�oH�	+�<�..8huu��6Ã
����Ib ��ϼ�gc:�YP(%@�w��|��<�������V�_���p4�yH[a�>��ïX��o��u��Ʒ4����}�6u?z���+��̷��d��%~���gM�A%B�+�?y����*@H�#>��E���٧�O�_1� O����c+��;�8�@�y~<4����]l���߽�a���HR�?{���8�{�Ǔ��w߇�q�_/;��i8 T���{�ۇђ���
!�߿}"�G��y�{ƻr�ʌ*c2��ӗ����W�<��������ޯ����{zOd�����޺�~���_�<�i�{�.��5����Y,_�Jc�x7�A�\;$�������v�7\�n��ݸ��u�#Pc��\1�!ن;�7p�����A�x5����[CtZ���:��n)�ZO6]�읶M⣨6�&n3����n�l˳�v�0.ۅ�x{z�]�.��ȅļvlWGoh�2Wn��nً��1�M��]�[�g�m=Q����Hɞ�^nr�A�>����l���7 =F��ѵ��ո^����Fz�[m��v�f��7VCv��������5���C�?��{��6�RT+y�nd�*�P,<���u�+ �٭�!}�oa�Q�Y��
���R	�u���f����	�1
"1�D{���E�#��*�^���3~�]_��g�hT�
$�(}�|�����%Ͽ~�gRu
�YY=���K��W�6���z�@׳�`&ۄ�Y���H,9�~��q��jB�@���hx"<	ڽ���]��|�WW�4��
�YD�}���td��� ���E�O��������i��	>Ww���no���zo��m'�*J!Xk��~�ѝd��J�}��p�R���~绁�3�ׯ�����R����g�#4o5�Pɟ��z���:�++%ed���=���hk�����7�*IXS��܇XtaXQ�@���}��:�d�+%e|_^Ͻ@� 
r����ݰ섈�	���a���14����;�u�p���\]���F�ۜ���L��_@��>͐:��Z�����߾�����k�#���� �����w�S�
>�W��ԂβT*���l�IX_��o�����8frH/����z�i*�oqϫj�k�\�v
�[�;	�؀tc>Q��:�]� g�&؎�nh��1�Ɯk���h�w�G���po��(P���pj`�GJ�0Te������~��3���Ĩ{����@� ���}�M�
A��o̾~�̵3����#���C͆a�pT(0�>@��O�y��:�@����2W��}��M�A%B�+���~�?qﺿp��}�ߟC�=aXV%�>��Τ��Gȏq}{>�x� �{!�p�q��@蕇y߿l>>�Û���w���������9Ґ��+Fo��}�'*P@�=��{�q�޵�c�9�$�,d�T<׿}��tIX]�L����ֳ��
����0�A#����dY��{>���7>1����S_���:��*A`V���������������p����s���O~�鿏���3<r��Ǵ�f�'����w�\���-v��u��H�&�����ñu� 2���M��|���e+(�_מ����B�*IXX{��{�u�A�>=�cdO}������=���ϤY�����Ͻ� j��>�u��pԂ@B>�f���H�z0n���� &�����E �.�����Y�=��{�u�d���>��o*��;n���x���h�|���i�3���
����Ì6�Ry�l�gY(ʁD�wϲ�3������r�Z?0��
�"}��wV"���sv��Gy�Wy{Ѝ���G����m�(�rL}	Ԫ����;jS���FDR��j!��-۷p���3R� x{�=�����
5�F�����7H4�-����nz
٬�߳N]C�!8.� 꿤Q�.�O�@>��YA���s�6��*IXS�����~>�@��H�=��Pz3�Ad���A����w'"m�������E���] !�ޟ
>�HP�|���8�q�߸_ww�������{�9IȁR*}�<�p�Ae�y fo�H�<	𿦢���o�?jd��
]l����gd����s���̃�,�k�^�����z�|���\������Ww���I�
��V�����:�FT��d��}èJ�ߟ>���Ώƕo���F]_$�����;织^�l���[�F��旐:�I�~�͝H,��Y�k��y�^c���m�ַ��&Щ*%ad����!�V�@��}��;�������U㾱|[j;�e}]>��$ �\4M:��k5x)��{�͇�X����!��C�|+;�g���
�;ן�i<@��'���gY+(�P�<��u��3ޏ��:F�с>|,~W� -�5�G�G�
�Xk��y��:�P(���>��H,��F����p<��|�<��~�+C�k';q���>����;	��/{��?uJ�b���)��\G�1�5�p��y�M�{s]{M{�κ73EU�2�fn?{� 
�<�!���g��=�
�濿�K�.9�X�*q'߻��ΧD
�YFJ�~�96��e�}�����O�V�Ͼ�8ì+
0�('�{��:�����Q��~ﻒ�@��S��1W�z�'~dd �F�E���;r��Y΢2��l�S�n�86�k�����i����n" ��� ����f�:��Z�P=���ăФ+F+����� E}���D� Y��W���td��%@�Ͼ�g蒰�_���!BO�7�υe}= P>D�'{�?~���>����5�Ϸ2|2�T������P;�,k��~����SA^l7!8/s�'��|8�`V�~��ѣF[sK�N�7��y��؁YFJ��_���g6�T,IXo�z�k���n���<a�°�0�*y���l�N�+%ed������8"H�k PmD&��(��o۲T��w����|���$�ot��B�HV�
߳�}�'
���_g��g���\��c�F{�|ϼ�C�����V���>��ѣ4ᙸq�XW���l8�i%B���y�΃�>�
��쳢�+}$��@��oP��`Q��~ﻁ���=���|(��� 3�w|>7�]�T�guMX���`� `Y%�ns2Ź�ơ����>�^P?Y�O��ݕ���M��.�m(f�AS7����we������N/�����4��>h�S�S!�=����V&�J)��Lz�ݲ��{m@�>M%��z&�����,C�Qk��e�7�vgv���g�<�$���)��n�ʑ�� :B�{�1���of1�aӻٓG4V�����5@��-��3J��][��y��6_���c*�����{�:���ݵ�����B1zM��g>���� ֑��`\���M���O�v�����8�Kݞݽ����|d��{
M�흦�B[7sw��gftnk���q_M?n+y���ɪ��>�6d�4b���vr�������yw%�9Mp��;=p��½��:^���&Hp����.�B�=��]U�)��;��ݰ�-����0=<��tÓܖ�4H0�ux��ދp�ç�2$u�=������u�@�=���Q�}���X����R��x�8y�y���:�o�ݏ�,~]����G���0/s���6[6Ƀ6ۑP�����*����SU,���/��N��x+;�v^�H��۸�u�f�m�DӴ�(r1�.h<�*$��1�AS�N�H�H�L��WP���ꫪ�sj/(�'GW�u����b<f�eI"�蠢7,B�<�B�/x�����qZfب�uŔ ��C�E���<=�`fp�=ڷ�^������W8�Q�;��u�ZR�v�pԹ]�|����'���iw�!�}z�y��p�}��m%���=NQ��mmKV�e-�kGܳ+iVU)i�qD���r��m�*��H��ir�2�������;�aW��˹|���1�kX6�j-Km�)�KQ�eE-���KL�����Vڃ�-��m�&5�V����G�a����e��EJ1�E�s,-�S3�����
�������es�0j*5���f[lP^l����(�{c��\�rsݐ�ˎy<���v�oe�W&2s��ȋ���ێ6Ç�DW2�R��D����Z��fc\�bؙmr�F�
K�)h�(�գh����ť�Z��'m��&��x��`^���m�ڎ&\r�QiFZ�T�Ɔ+kR��W���KmKTT�QkD̘2�ʴ�DV�.e�Z�R��h�5l˙1.6�d�R�cR�Z+��ܦm�1\L�h�ƮfL�c\�L*R�����ib�)m�h�֫��DknaS"�*�$J��G,�-�8�FZUs���8b�7As��i�[���GF�U9Nˎ;1ڶ�/�ۊ{n^���N��u�����u@� TA����k��l����uv�}��)���읷W��yd��B��ږ�nbx��9�[�X�-��� nD�W����b��s��;>�5�5�
��b�
n��6F��q��]Ghc��ŷ-�tu�Sc �8y�f�	��^7g����xc���3ӌ���[�M�`�|���ڮ����#x8ב�;n��<��\�y��+j��ͣ��u��N5&@<�k{�����ۗ.^�[�:֞;k��[̗�y��V^��vγɤۍ���2.l(�s���k�9y��쎌 6��u��ˮ��l��`啬�0��J����k�;�NB-�e�)#�:�x��6�c-�cz�����kceו���u������46��P��� [�ổ6Ϫ�98�	��-i���nݹ��6p�l��$����y���{dn��$M�z����$�yܽ���ͽ�܆�Н� ]m5Ɛ7��5�w.ŧvY۶�bH"wY�f}���6Ҏ<D�ۉ����]]�I1��sm��,H�Q[����r��۶�[uǢ�`%xP��0� npa��F�v�Pd���n�6��`3��ɥ��s:��A�ݻD�D��[k��c5��G��p����s�����-.lPt�m�9<e�7n���-��oW%r��08����t
���;�^�ݑ��3\��a����g��s����c]i�ݞ��v#rg��,S�l%�ݞn�k������K����=�8ŵ�i9��}
ѐ�v㤥�gckv��$�w(�ۇ��m�>���.�a�WnSmyd��� �-Ůθ��r��ܗn�1��wV���f��ͽkku�6z�s�&�zr�c�[��;�l���Rj7Oef�\�������t���q�x!V��s�n�.�t.CC/��:�O&ma���R�bݣ5uҁ0����I.H2ZJm��G'IN.۶Y�>L;d��2�N�@nl][�#vD�ȹ�sx��Ƶf�6��;g��Kc׀�q��;��s�8(�ݮEh^��y��u���[Ǭ!ț��DhK��C�u<��v�8�e��li����ۇ��\��E�q�<Bh�˺�F{R��qn: ^����ͫv��۞Oj�z�nW��?��K���g�]�a���Zͳ&.(��K&�{��Ѕ��[.���]u�[r���?���C�.9�X���S�y��{���
�J�����8ɴ(���}���dx�>s0���?)i_��"{����
�YR���wH>��p�֝[�Y�5è�;���ïX�����6{������g�HV�
��?w�@�AH,=���p�=*A@�}տ]����@���F/�y�5�te\1�M]k9$W�~�x0�J�H,?s�=��u �T�׏;���s��>�3��� ����@u}{�� �H[a�?y��׬
~V�0�$��>��=/��F���W�Xp�Ԃ�+���g6�IR���W��>�@���(�E���z�>���H,�W��|ܜ��
k:����kWW��X{��<�z=`Q�	 ;;��V����˔mX�$x��� i �q=�{�u�+(�P37�Q��>�����WB�(����ۮɃvwGgm=/&�v��4��{]3=��ij	Q�5GȰKC�b>����G�}�Ì6��*K�=�{���d�*J�g�{��:��+Z��z�G�4�|� �y������!m����w���E��0ఙ,�'׀DW��vg�u: VVJΟe����߾t��k��?�hƌ��/�c�ݟ���F�}��q��(Cjf��D�0C���H�!�:C����ى��$���ca�n�z����<|�����M�RT�����{�u�c
��%O<���ΤN�{��������ߗ�GTuϽ�"H��06ZM8���dd#�w}��� �,�|��q ����{dP��蘛������2<	����χY�J��P�y���l�V�p׶� A�曊�g�2�t�vJ�����|��s�T�D*J�a����Ì�����~��@�J��R����}"n��B	 �*o2|,�>�Tw4��a���Mx"������@��� ����gM�����{���IXg�w��u�aF%O|���:������e|�����mϻ���~��}w��l��!M˜���FX�sv�5m�]E��`�ŉ��w3e^'f���?��v9�9�]_�V���v�+R�?y��s�!iHV�
����yI��"4wuEN1� ��p��|(�@2T��C�=��Τ����[�u��es9�����z0�J�Iu��2�v�w�w������Ȁ�H�?}��u+�`V�]��p9�x<I��Ø�G?(��ɋ��g�"��Â�e��^u��(� +(�YY+���vr2m�
����V}�/�.�}�e����(Kq�/#=��R�� ��ݷ6;s\գ1}�[��$�[��s\7qU>;���۲�|�=��o�����BG�߿�� ��aRX�����I�
�Y(2�o����� _<�((l��p����O�M}�Nܽ-D�q��>
#��M��" ����m �
�����ì`מ~�#O�C# ���}���A?l��JW&f]��Mg��62
A|�̐=��֟NF.�_L�vn*��@�^yϼ��Ĭ
`X����P$�G���O�l�Y��!������oﯦ'�t�OOdN��
:�s��G�,b�7N�Ƚ+A0�74��?g�d��P��YD��~��������d�����B�*%a|���:ì+�7���_}x~��T����:��VJ2�VW����N Y�}��f�:֝^
�?{���;����߫�:k��^��l�!RF}���ӂJ VPO7���gA��8s]����e����#�ɑd#��(��l3ŲV����Xta_��惌8��Rw����:�A��P7���������7�s5���� �(����s��iAxd��>l�W��Æ�e�5^ �Dz{��E}۷�D� 4��#�+���G#'���RVo�}�8��|�G�۽�#�����_$f/ߟ}
����ɧf+�.W��iupU�B��;�����o_+n����xwp�Ÿ��lQp[��$v]	�;Wd����w\�����=��3�~>G�@�U{>�$ �����a�a&�H,9�~�z=`Q�
���߾��x/��иu�����&O�ETO]xG*Q��~����u����
����E�,�#�;k�5۪�c �ѷ6.�-�4��[sp��K<ǎ�ٽ�8׬��]�����>p�.������0����a���T*J!X}����q��*�Y�w��dd#�>�5��f�j~��|�k������K7��w����q)�p�I@b��`�}S�H�/� �����;�/�D���3���<�쑧�i
�����＇R��IS>��E�� #� |��������몧u�����r|&�.�����5qִ��P9��߼�a׬
H[@�￾���x%�<�n|V�!58��di " �����w�v2T(�����Ρԕ�~���Ӭ4�cu���8ñ�_|�3.>�d�J�wÈ�^ #����Ì�P(���}���u+��c_.��p5������N�wH[a�ٽ�6�F��4�M0���	?s��l�u��VVJ�w��82m��weHꉼ��|&��
>|�A�ID�����ԝB�Q�����~���6��IG����֮�OB���<[����ޡsMO\&��8��p�#@������Ʊ4�u8�'�B���F�G�ruN3�x� ׵�[���k���7���K��9]����OTnם��n�8Z�Fv��H�WU��d�H[6"�i�M\�Ը}y7:Y��5F������k�d�1��q�9����h7<��Q���+��g�V���D�^�⑺�t��K��s�l�uO�m��a�n�3�w
��/N2z��q����vn�Uo"��k��u���D.^7Aj�K�E�L�շc<\�q%�ˎk��Q�j��,����#	�JM��È�ü�l:��cR
�����!m!J>��k�2(#v���s�L��<���R
A@��>�g�IX,���B��ه^�Rt�G�������\��G��ɩ��>�>DJ�~���p�D� �]���p��Hx(��\��퉕�|n��i�|*j�t���D+�Y�=?O�"ȂβT����ݜd�$�Q%a级�9������a�
�RX��{��:�Y:2�˿�ܜh�=��!�.j� 
#���l����ǵM����:��R
�y߶s�!m!Z�EdOmxE#��/���>}������9�옐P�s~~��;V>����Xi���+��u �_{���OD*J�a����Ì�׻�3���y6���~�~w�P;�+X�뿽�M�)K7��w�`W��g?~�5m�����B`7d��v����$Ӎ!�T�]Y��p]<�-v�	@���Xp�Na���>#�W��ΧP++%ed��{���B��T�����w0�
�z������
��}�Ă��+%_��ܜM�S����f:�K��S8u�Xw�����F���*�c�}ظ³uSp��&`ͥ�Ζ$�Oa��֊�wۗ[K��i���E�� ��pDm�� ��+G9����~��JB�B��[�o�yI8�YS�����Ԃ΃%@�sO\���śu� �3�i��>}�_��i�sSZu�CL8¹w����AH,?k�|�8��ʐP;�5�s���w~��������7H6��������^�+f����n�4e�\�G u���C�}[�~�9Y8t ϴ��� }��|�͜��B��Q%a��~�p���+
�������ԝ�}�yނɌ��2��o�����<��f�:�i�����w͇��jB��?~�g:��������!���Ͽr��J�Ybw~����td��%B�矿}���>�]d�T���h�] �CJ�\���ʮ��]��D�:����N�Jcr\h��_٥2�2����<	��r��RPB��Ͻ�8��T
%@�����d`�|o�������I������K���{˯ߴk4�Y�i�kWp�O߻��:�Y�JřJ7-�B>��Q���U�#A����D,IXY�����Xu�aXT�<���u �v2�a������~�~u{�����;fq�8A�D`���gHz��H[@�Ͼ�g;HT��]}� �v>U��7b�/D��$�ń�!�o^)�����jp�/2֜�qu��8�M�ߧ����U������oi��� H���@�D
�@�>߿{�q�d�
!�߿�u�+
y�_�����?C׃>�0��B����_���<I�
��V�{���u��T
��翾���X��w�π�쟺O�e����<��ﻲ|,�>Z��I�b��dXy����@����d���=��ɴ<9���sy�8$�)��߹��*J����u'b���VW��=ܜM�k7�,F��뻉!f0
)���@&.�Mx�(�u]�ݻqi1kn21����Z���>��s����J����͇^�+R�����9Ф-)
������}�'#��{s�1S��pa9�O��Y��+%B����gR�k���f�Y��+��u ��?wp4��B��|��y�g���9���gY�KP(��<��u �Z�~ﻁ��)
c�Fz_ٞs��:|*"~�2�Ca�ֵy@����g؁YY++%}�wݜ��B��T��}�y��n��~��Ԃ��%O߽��Τ�d���#�����+��)8�
 �P� ���:@ȯ���mug �<	 o�s��v�����{缁���_P�_}��g�	���	�*�IV�G�`��N��53s�ߚ��o��B�s^E^�T���7�=����\Z��1q���n���L�_u�k׺{����Lg�%@��;��!ؒ���g��i�sS4k\��r0�_��a�IP�*��y��>��e9�ad���� " Q}P����R��绁�t�aH[a�>�g�̓���oʏʉ+�B"�P�}���=X�6n��]��*
�{l�^J��zGY5���[����'
g��cˑD|@�J��_��=��M�����:��llv!p�s�H���y�#�	 �Q���绁�]}屳Z�3Z/�X~��y�q��jC��{��w��ծ| ���"�!��C�|+c���8�R�VX����:βT�����zF�`%�d� p#��!��J��2�˫\�C�;W����pa��
�X{Ͻ�gY�JʁD���k1�5�5�<=@�+��
�����t�A��6~�g�̓�Q���(l2�j�"����E���d�^�+��8����~�gM�D�
$��;�^G�>� ���G�g2�/�v?�B�ded�+۾wrr&�({��}r��35�S8u ����퇯X��A ���<��*����]��Ă�s�I? Vߟ��8�Y��P�}��u ��k��������� Ӿ�-�~W�<��{����̗߯��s�N���@ϖ���GDjzj��w�S\��=z�}�[�B�/4�m�-�<<=�U#���C-�����\�Y໫��_������������]�vtӇSZ��å�˜\�����	s�[r����'E�5�s�f�PY��Ѥ�k=)�lt������X�qĚ8��r#2�B���펷]���7��=�(ɨ|�v�R����s�q�k�7�Q����;�r�z�^-�<\	�	��@oh�6��=�ˎ-�V�+��ل���en���k�G�1��f��6;������6�W53F��CI��9��IP�*�����Ì���	P)�������|��4��il!�oI�����7H4�-�ߟ��:�0+w��}��8���E�<�~�E�2�Vk���<�３�.������
�����}�:ñ�H(���q'D+%����k��o���']������p���D�Mff�g ��������Ƥ(Z�}���$���]w�|2�{�~��y��@�x�R�
�'�����Yђ���
!���Τ�k��n]a��Bi���`yU�6E�4�-��I�B������vu�d��*?~��u�R��������Mş�UN�F��C�%�}��fπF��-�SlBPڟ H�G���$Y@�2T��|�ݜM��s~����}&!�����Ͼ�:ã

����~�gRv!Y(��FW����ND��_&�d���Y�B$l$&YE �N���s�fAv��=���l��.Z� ݎػ_�?w��N�Ɏ��/Ǩ%a�w�v�+R-߽���v���+X�������@����ڙ��!�>�y���g���d����q�+
h׮W���5�CL8¹}������e�-�UO�/bv�]�,N���Nl�ܙ$�w>��(�9LN�Z�";�PH��F\ƩX���Kݛ��$�����}��3����@�{���u+��Z�|����A���ϋ��u߿S�}�s�����ux#�0�^ȰG�鿤Y���� �������hX$�X���؟�N[M��~���'�A�Dݿ}��;��� �_>�p4��p��A<�!�	 P!ϯ$��_�RϞV��P9矾�ă�B���}� i8 T�e����ì��Ϻj������?I��%B�3���Ρ�%`��שp(FF"�,�Y_��$y�O'��➝Pr
����$q�����hou��΁FZ�)�I2L'�6�@�G4�ֳ��uڜOgTl�;6׳�^޻�����-�SlP�
u9<I>8orC$�O�(Qni�EG������$3�5�- �B\��y�v2z�rwĐE�܉�>&��Ux���w�:��`Z0J0�7
9�,�>̚�'��b��NL�*Ly�[��v��<��Wv�_q2�v�={8{j��~ղ9Q�M��OS�~+��}۩��v����I���wb�^�S����)�"�*\ǧ�х^������n�E��6�`�\df��E!��..�P�I��$9��ፓ;'a�ws��Sz#g>�d{7��q���{��;��@ �h����f���-�����C���c������5Kȫ�"N�8�p�HDU�,q�N�Hx!X2�;�,�/mēSWY���E��^A�O�W���E�Mj�cZh3/�6���BU���غb[�8>s�ߺ�,��p�o��}�~�����]�ҹ�J�i�%{6CעTfע j�	d�D��/n�(�k�U����j~�l����Lź��j�.@^n�<X7>��[�a�5!)��deY�q.�1֙��)����1�ʽ;x�כ)M�l'�&L��҇������we~���>{�$\s�{l��C�O�[�aN�oMy�+�H�-j��t3C�d��XD����:��JZ��$'����<�h^��y��\�N\wځ6�ޘ/�wv���/M����M ��(=�8̓~�6'V�kh�����'w���G{k�*斊T��ZD)��5�ril|&1r����G�\<�؍jݠ�ЯOx-�?�]�����cs�ڙ�.���{w��0-P[j�k"p�����t5T���C����?h���^Cg5�n�;!���=z莴/�*��a��f�Ǿo���ǍD[m�)a���iJ���Z��R��m������q��ڴR��)��0��Z��m����he.4C�Ve̸���jRTQ�9{��s�s����;��������U�m�p���=�Ǖ|)�Lv��n��g�*�`;v<n7 �;�c)�r��1L+�fW)�S0b�Z*.Z�ҥ��,m0r%��V���l�˕0�2�R�Z�m̭b�.ckD�������\s�˶��)���lpvm�)R���2�\h�#1.���p�o6��7#��̢R��n	�\�0nQ��ʵ�h�B��ܥ��q2\��Kq��me���8�)ceZ,TkE��j�JZ��asr�ƮU��.9h̴�Y�-JUF�+�q\�Rҵ��L��c�h%�UQVՖ�+*ڣ[KA�j)F�Z�Z4��ժ[n\�Ye�ւV�kJ��֥����Z��b�E�[D�Y�R��*�F��֭L�pZR*��4��e�����c\�?����� �I��\�	4��$9��a�aCQ�U�ݕC�.⓴�H(�̲"�vUI�v�V^\�
�3���ɼp<O��]2(�i8�l1 ��]Q����Gs������@��� �@���v�MFM�O&�r��-;q�|0��+v��;s��OC�6V�u�-Y1�֊�k'R�n8_��?���9~�澿xI9s�T|H'�۽Bz��(>���Jڟ?��T	
#q�l2�6 �O�{ߛ���:�MM\�}�)�� �r�	�n�UI���!�^m2:x�@��d �L���ݽ4H$��ڡ8��p���I�������*�F��?C������V*�8]���|�͚$3wz��f�jy֍����(�N�0;h�jofp���{��^��v/�n�VMiL�1�ڹz#Q1�q'R��)������ݯ��<=��}�U�P�f�GA���ڄuK���$��$9�;�\XZ{��I"�fУ�������p���uWƦrN�O��m۟��ip�Y�<6���4X�C�w<�����י���|�����������UУ�A���I&��ĂC�������	���O���!CA�8QGL���g��إLkyT�w��{�z��7[,[�)t�%�vP'�"��L4�6 �t=��A8n�Y$y��v����g��ww��"���=6g�Z6��P��j�����ݙ~$۽r(���b@ �>�5�[�Ff$��7��Tg�@�lAHC�0�H(��H���*�Ξ�0-84VumW�a��`��>ɯ93{��D�.�wUx�UF,cE�n��U�C�٘vS��6+�g�@* ӂ,�ê�h�zm�\T�yλiU�"�*.Tr��{��ݾ�U�]��q��j�0���3�<��Y�r/g�ǆ�0��D]6�h^�45���\X+v=�z��:���1�y��N�':������x^��;��ֽ�n����t{��;��3�j2k��'�97#��R�ǩk{=��]��d�'�u�+�S�ss�{r��%ښCq�Q�;��;0���[�����#������h��368��l�&���nGK���]mϛ��n�]k�o�߿��:�3)�_��9TI>:f�C$�E����nb-��A/"c�3]TO���7�%�\.�CjO��VP�X��=�"d�$�qM�I_>ʢLl%�9ڛ��g+lW�´�H��QK��vh�o��c ��/z	���o��y� *�~_�P|�;\4f!�8BF�ީ���
�$a��w�d� �n�;�rdO[���'^�"���R-MF�ƪ�k �v��=��&%���q ��{^�P�{��@��7�b�n��9X7P�.���Ƨ�@6��7K��ޯ۬�F�A�.t�D�?C����I=�2��I���U5gJ��u׋9� 0A#q�U H���[Pч�.�ʢ3�S��/q�nͼ����7�1a{=\gJ�6|n�^Y}�5��7�9׎�v������Gn��s[�ا+���B_9�|(��k���W�{�����f���X���V.�Cj��7�A'ww��H�n\�',�.��x���(P&�w��#c����P�8Q@�ʺ��م��w�@H$��mP$0A��_cEJ]���~�>`|��Hn��Cb
p��ޜ$��ob`=�Q�M��_7�`o���0�<���b]w�#;"z�D�S"S.!՞]���c6A㥶�\s��F!� �Hb�vp%�����j���DA���H$ٛ؟�t�<�s���l�F��Ux���@6!$!���IE�� �X턻aZ>Jo���w�W�����Q�ySs�����-�hÃ�T>ʠH#K��H�K��Э�D�`���'ck�c��T��5v�O��'�u�݋��C�LΦ�*�d�K�z^�U�b��T�i�5�z���d�ם��;=��uA��8�(��< 9δY#:��A6]�K´[
A�l1 �eaN����o�d>��ɻ��I<��H$���W�hB���c [m����ВI-$�ǅs�px�+Գѩ���(g<��e�K����Z�H���<���WjI"p`Ҙٝ���A����۪S�I�s�5���.?~~���Cb
p�s��O�}I>�}�^=�r��37B�突�w���\��A�!���x��\�J'�++�Ed��N�A>$bw� 	���^;���:ﲸb�(�͆�|Qy��$�<�|I��荼���|	8]���H�}�^'�7f6j0��a�(��=5ՏI��AFj���G[���'ċ�ޮ��З����B��y���l�`?C����x��K�s�!��rߔ�G�i��E���N�s�>���o%�v�F¼1Ǒ]�\N̈��������t����_��Q
m6�{�̯Q#kw���.b��:.�W��۽���ު�m������Q2�=���qs�ۊ�8g�=vM>�E��;0=]m��s��&Q.3���M�b!D@h��=w!�	7���	�7]�THt-���Ai�9>2���$W�G ��ЇA�Hܚ�Q�`�Y��th��d�|H��.�z��v�4�܌�������A�!��0*����M�wM�:9w��鼚� �gu
��j
H��a�����}JN�����
$�ު����76�6�71ϗ�s�����n!�LBL:�.}�+Ă:�$I�i�wjzhsozE����[o���p ��}?@S�a�Hs].�E�=L�B[��k�F{�vX����S��m"Y��ٚ�V��n{�fQ��y�W=�f�����3]���O����3�}Xq��n9�]�.���Clv�C��e��cUq��klu�&�2�!��yv�ݓ:�c��į��{86+3˃�:RP��l(q��r��ڊ�4fy�sӇ�<�mڻ7+��H�.�v�����ntu������<�rv��b����5�<�h�-=q�ns��ֹW���um�l�Ar\�����B>ێ��.=u�Xn,��sۤ �.w��v�r^K�n����ƫ"<u��	�D(/s�����P�4�?x�fexW�/zh���rpn���R��l�}�D�oQL�B1uDvչ�_WN�3p�t��x��uP$�FV��'�Q����qU�3IQ���A��0�	���I$enHA ��!Ft�3�I;��B�$���=�|�pe�L
�59�L�oa}fA;!�>*r�kĂA'�1�}�7Ս�6*�'bPY�v�uP1�`@�	$a�XmψOvD��o(
�7��P6Z�k�jh�<E�d���}T	�,����돭�/��W����:��v�\���]���'6C����M~������d����3&�O��Y�$�N��U r糪��i��+��\�OA$ufL�rB�,��-;�7����B�?6,��c��t������GKfu��:Ω\��k����o�u��3��L���{L�M۴��}4C�s��f];��xxxNÜ��$���$����4H0���Σs9��p�e�Ci9��w>�	�w��������]��$�2�_��n���9���m���'f{k$�+���q ��H�	�>���	��ڞ���Ng&������.w���I�A�͟Wv�ͻrmA�n7�"��U O���v��c��U�i���玍�����h����ip�^kci�{j:�n��R�Ah��Y�5BIa�~6�� ���I��T
�#x�Nx���$z�*���q�Ä�&P]]UD���{5sB���$seW�$f�mQOO�8^u��"�4H�X`�(Bm$�e�D��� �ؐ�!����v�-TKP�tFr���=��v+粴��s��W���k$V��Bj ���7�en[�+�\��T-�u+����������7��$���mQ/xN'�T#��{g*��R���x�gez� ����^$�E�ꑮ��Ϻ��&.�ꉈ�Aci�ᖔ8BF���$�F\���[7�
6�f���ɢA"��j�$�E���M�s٣���A�������D��m��'�m�{y�q]������m�Ꝼ����?~x�2C0�009w|(�A��٢I]ι �TRy
6��n�Fx�^�mP&l�)BIa�rY;2Op�sy�n�:�Q$�۽�@	 ����c�p�6\�_Mk���/EE�$�Ra�)��6�$I ��Y�Gة�I��T	�w;>���C!B�h?v�]Mv�v���-�Ϩ`5�"�� ��9 ���^Ľ'��} ���i7��t����w�&�U�F���M-N9��#�֣]��S��v'g@4,e�qt/j%gp�+��������E����|2�&X)�m����-��e
��Ru��#A]4�]YTO�]�1 6�eP�f8\�hΘ�BĲ`��,��0��ұ�y�sE��ܓ���2�=6}V���w������-�eC�8]�uQ �2�\���e��q����u���$�G]l�%��� ��I�T��ר�Mq�6&jS���|}�\�	�}�^$��*���5��`��h�E�b(I#2�n|B��I=�2h�zŵz"��d�L� ��@�Io��Ƨ�3$�Ra�)���w��S����Β� |_o��࿽zfu[�y�a�I�Ee�������B�h1>;�y@Q� �ntћ���̩�Gv�	����M��U��|���+��5��'��B���k:<E��JG�s��xV����g^�cv֕X�ݏ���WG(�G�c(I��f7���p%���/-��b�>�K^���C� ��/��+	+�V�4������3�f�<%/���uI�(J��}`,禌�5��Ӹ*	����{��s|6>ה�#�C��������"�)�x<Q	�T�PG��˯�)�e��������#|�!�͆��uó�F���v3��j����оW��m���'��9�^ge�Y��v�����l,�eRɇ��1�~λ�̝nڋOx���Q)��5������o7=��-�?�������qf<C��j��>ZO��7{H�*�air��ysޤo�칇K�/_q�`g8�Z�OOn����x�]9��nz�V���`lD-��bb�I����z�Úӓ^ǜ���$��\dUcb-um^��T�t���!,0��ys�����Vf�����9v��g��W��`�K;K�M	�wB�E�OwsbCҭ�'��ƾ�d�{ܐ\W�n�,����t�Ku��ucL�/:��[�����U�}�e�A�/e�UsH�u�%��4�*����kk�g}�,[{��`�yxri쓰_�@w<��B�j��o�eB�SP�~�z����&2S�@U��>Rѝ�6��� f��Đ��F#a����Qi������N������fK��MY�f{*�>�y�et�W:eL:�y��$�|��Vp��{�ػ���\j�{���ØN��m�JV�DFҫmTE+U[*���Tj4�l�ciERձj�j�Ҷ��TKE��1QЭ[-��ҬV�b�m�����*-|L�lmaJ�Z�T�[I*�m��ZEP�Q-�+(�[eaܳ31D�TI�R���QA)Kh�iE�-�b�Q0b�j[K(�Q��B�em+Q�m*��jZZZh�+n�V�ƕ�l�emEFڥ���V\aQJ�գ)YU�����J�("�l��ڱJ�,ąk
���T��ʭ�[ZQhҶ���Yjc1HڵjUW���4�[V�EZ[l��ЭEees2+���U�2��b�X�TU���ZRբ#kBҫJ-�fU(�m�6أJTmR��Q
�+ZV2�F���j)e�-�*Z�d`��V�ƭU��ҴJ�+h�EF��m�֕P��b%��Z66���Z�[K[YieŴ�)�ST��-�B�#jW`���w��7���:�l���6o5Խs��U������gu�n6%M����f�V�۠Nt����`�f���q��{]��=�4�[S�+�i�g�㨫u����3�]�۱��c=nwי�g�]�m�>�-��\��y�s��z��uT�z9��d2]��Ѹ;;q��=X�@���W�F�;��\Y�Zf0����G�tl�uY�\ʱ�N��i떿�^�ܟ]���v�Up�7+���2"�˴���7$�qB�tk�u�T]�����\�\��8�on�1Zڹ���S6}lmOY����mi��<l�A��3��v�����$]<sF}�<,p<!;���&"x5HL�0<���x�m/��v�=��q�:ð�A���컮��\��q�x$�;�S���j~�u�8�e���徯��H������]Bl�wK��H{v��0���M��ݺ���q�TΞb�$�u�ز��� �Y���h�:1�)gX��X;h�p���L�=>��n�ٳ�v�`��s;8�\g84|�ۧ��k�kNN.]��)��ޓ�{i��YW-�"n}��y��L=Z�\9y�x��;<8����	�n�9L��=��V6�)^��N-�(�2;���k�g���[��-��jM��g�y���V�s�p���b��O���y.�X�-۴�Cc��遲��v�X԰=8,�[Mmv���V떄�w`�w)�Ҕ�7�s�H�^����u�#c�]k��O\uq���Au��,�q�Y�¼�rl�J޻��3���5�Hm�z]��;y��O�O-�G�sW.9�MA��n��c���#k��<mf�+�95¡���{u��8y��r��J�d���;q]���7C�7�s*�J���O��}��Ц7`z�N�[hM��u�a�بur���v�>��h^v5�5����;	�9�����E���ѻsu���]>�yd*���y{룱;s����;m̶y�9��i�=���HYY�nv��i��^�ےHBr�3-wY�C�3W��L/m��nx�a��|t��ıKnp���\�{N����ee�<�^]�.ֺ�1��.kv̇:�up�p��z5�^ym���8�zH;�v�]��a����d_8:�E�Mn�%I)뙊Ňt��\麼�k�����ce0����z�i���s�aٍ���*��n�α���ku��6�r	���D�[�v���t9.^��sul��E��1�����?�;��%���p�9�컑$oe
 �O�w:��7���+%���/>��g��k`$�H�f
6T8B}�[u^"�C�}[��WtؒI9ϲ�x��Π"��7�$�A˻��I�����a�`Ux�OmQ��nt�$W=��k.���|�ēz�*� �Κ �9,�����a�>!<�U
V��]��=r��	��U�I"��Ԩ�=Xw=�;�B�N��f)6IJ���F@#j�g��ʻ}�۪�"⮪�$^�uP�]^���dV����������CeV�g0\�hݛ�a�]j�9݁�g�Zך�W�ٿ?>|�λ��9�sj��{{=�"���<q8���p�n�(Q;��Tc��L�Ba��9��n�"�T�>z�T���1V�TMt�EE�f;�O3��N3ݍ�ѹ���jûŇ��"�9��6����'E�<��]41e�^1߼ ��3���A��kďl���Oh˶��\�r�O�#1��A�҇H�κ�	^� 㣷.��q�l�{/��	6j�C0/�`���I�A����N�ٍ�|]��׉�5U�O�$n�ʑo^9õSx@'ު�ʠ	�1TBH�d0ېQy��$�<ɉ���:u�j���T�Q$a��9ϲ���f��u�ەb��SR���|����[wGld�ةۆw\��mj�Ph#��f��)6IJ�V�*�Ǎ^D�Nk�5�;��a;;TO��W�E�\0�Dy���^P�G��*:�ime���3<	$�ʯ"A ���T	�'zC{���=�$Ff+i6�	��uG��O�� �OeQ�8�\i��B���g������<�{��}�;�;]���.#Z���2��9�Q�u�� ���Q(��4]�hvN�%^�L��1�TfϜ����O�;�H$5�O�$�g��P��:��� �-ChN��Ԫ�/�	v�|x�\����s*��[��_7��˒0��=��	@�a�`U�ݡ@��ޚ3���/GEͼ�F+ށ ]9�D��ޚ��G��W��P] �P9�
	�R �G��K��k�p)Ʋ���q:;!���8ٻ_߻��?�P0�a�⋻��l�PH���k7#�/``<g2X>$VN�Q36cI��d��:�����񛈝9���A"�o��7��4H9t��%��ݫg��0a������ʯngt� C�������b����wW�^"�7��>�k��� �Æ�:�3�Wk'�2o��ΆH6�*Ex�ݛ�(�;y��RZ���'n�h�8tJ���s��4橐I�c����o+\-���	�4N��¡w����C������ {�x�q�:�,f��xx`��y[U�C�W2�!���'�;��xH8v�|��8^�T(l�om]Q$��uQ$��o%�'pUt�MW������м/;S��4N�&x煺�ضG�j��<u�s�kˣH�SG�{�F�N=����$��ޚ��H���qf��cJ�36H'ݹ�TV��l(��P��n@0vvC>&H��Gl�MW��E�wM�N���t�e�~<nDU�f.�F8M��J���=^��/%�J��RZ/�m���I>���O�<v�|�KC�oŴ���v�#l�>�I�q ���� <l�;�2�O�s��N.H�.} �gl�#���b!�uG��Hd����U�z�3�8FI��р���� �ǯ I��飢w���؉Y<�j��l��q��*5�E)W(���]�֭D��*��7
����qyz������}5z c8�g��?@��)��a����ۢ�ִNx�nO;8v�n^1�\�nM�nkU^�s����[sF4��K�,-ػ&2��k��89ݬu���-9�7k��Vm�����V�=�m��>S�q�l�u8g�r{9l������S�=¬�x9Yv�0���ɤm��ٵ�;q������8�89��������Bɸ�_t6�W=rq����\4.M�k'c���g���բO[z�;�u��#V��t�`�\��o��[�sDD��2�F���쮾�53DѠ�{�� ���d\�d��
�Yu��'5��at��$���ȒA���Ik�=aq�Ӣ'�^|��I%�(r`��N�^UI�����8�NWh�I�9p$u��@�cc&�D8 �il��C���'0Lg�(��	�릉$^n�f6z)5�q��g��V0�/��z�(Q��v���A�"�rx�"��@�}�u�D��y��F�u���-&��
��$p�C�G������t��!jB;us�9S��{<���%l�ێnݶo��]��8&C0�㧫"A �]u
#Ă}y��G2rW4��r����7�,H��ⵐ��m8�BF��$��辘9wn�E���]�����NХYj��+�v茅n���4{/��}�^��޲>#�R����Թ׾��U9��zԪ
{�� k8���$����|H������Y�x����p6u�Q�K00(L�d�+s:}@�W�~�����#L�[W �>��� ��xÌE���d0��0_l�oU��q��l�o{9�!�d>ʍ�Mֵ׸d�J�.f�BwD�8MP���
OS$�K�fK��'p�,�e�hI.����q���D ��F/XM麲�#�`0RHD8EA��f�c���N�U��g,����iI�������u٪���U���m0��ͦ� 2eK��ږ�]�� dvkPo����ȇ8e1U��e
����S��Ůʭ`��!����� /�{�*�P��5�uNkBI�z.m�*�/[������iЀ��鳸�y�L�~�s��Aѻ/��pi.M��w����ͦ�2�jb�Ԉ�I����䋬��.¦��]en�����2��  6;���� ������˫& B,�d��J�:�:Ks�'��u��J�r� }���~�Wx�qw��;�PV�O��� L^t�
��: 7�i���E�����`x��,�FF<o� ���so�E��7\.�� �@�!��1	�([��x��Ō��� +�n�ɮ����������$��,��w~�I$�W[� ?O_̀�~>�hФ�a��q G�[�',]#���i��p�P[ٕ^��BE�Ɉ٣0��P �s�,"���")����ȱ�R�s�ȡ��Z�f��LN!t��͟Ffu?� ��MVT���?m]S��>B�x�d}�T�I���\�.8�@-.v�='������4=o��76�!�\v��=�1�e�S͑=6�B&�n���5kL�1t��#S�X���Wq���qt�PiA����r}���r=;y[-��b�]�g�����}]4$X��0��K00)W�VuI�$����f�Ets�o7k�N�
=]n�	}��C���Et�U]t@]��wC�+`�
�"�xu�{6N{v:�cp�8�Ƴ��	m:�9�1���H�E'�l��B�n��A!v�T4�3����Ǯ���3t�	^n̒�C�E�`Cd�����m� �P�2��uVҞ��h��v�� H���������q���J���I{"��N��*���*�/$ ���t r����ލ��3���<���D�H��٩Z�tP�pfL�T���:�%E��ב����{�M0�"���1+��_��
,���J0Q�����4!���YpCl�P�.��n� Yw�X'���Ct� |tf�QWw��_�^���q�r��8��`�鱕�����D�諸��������o�H=���{�Ql�Wo��x��f1sɞ����{��徾Ƿ���:r���[��N{^8�'g�v�Ӕ'��9���:�s���N6�t 2l��t:�x�)��v�7e��n���`��gk�:w�z��!����-gn�k�Q�����v�Xy��l���'KT]q�Q[7B�����Wj�˶���c)mc��ԷOk��^�i���uu�k���[��S
7I����ϵ���O��9X��t��O01�۔7I�s�gpGm�{��&h���1�������=����7���>@ ���t"��S�*"���s�U�l�F��򠛌�XAA3!��x���އ������ ok�� 
����/&�2f�*;�y$3-J�Xb6A������� ��M�F��gu,�M?n�w�$dokQ��lE�:-��?'U-��7b�P�Dt]eL0 ���L�k{7�Y`Zj��mo4���bZ�f�D�y6�m�؀A��O�,�d�Oz<�;��LCö��.��i� ��a�YN����]B-��@�ᢡ��԰g:u��V�w�gR�jrku��Ǖ6�;������)�����G"���.��$ ݭ�
���w{�}�8u�D0��a��O�^�$�1���m0v�nܯ|.��hK
�{YN�m�oz�y{w��.�6n�u��z��}yh��E�͚�U�^[֯w��Z��5� ��j{���uܶ��$�]��$�Y�mTC�K����Z`�rA{cg�G�L�D�:ix�� >�ڨ �=�y���;"'ս�An����D��B�M�@js�F����5�z��}���s��i ��[h"#t��Ǟ��W8<����m��P<��\6\?'U.�ʡI�K�f�������7�n�T�WA���l"t�~ߛ�u�Q��s�u�Wڷ[ۗ��N'S��3N�exh�����,�-�����?���۬�t�ʢ���� ���w���"M��s�^�vυs͵� �����:�.l7�Q��mU4���w�v�j߻�Mn6A���m�Dlnu5D.��]��^.�m�LR��>�{艟��cCy���E��S�H�5�%eGJ�a��p%�Nn�;��BcIHǰ�t3U�,K�Zl�����淪2��]S����ֹ�=��|x�R�UZ�ɳ!c1{zFFSBҷ{�
%��=�{�R��'��%�-y2���N����k�Tr�=�Ǆ�oĥ@�֬��秄����8��=������|����?�+7��i��_Iq��5�jE�ՙ����M���cF���2)e���j��t��)�����S����������}�C ��M��t2�8��#66�em˨�-PT����;�$ZA+P��n?����?�k�?� �Lc�ʸ�E�N�L�U6oN�m���-��Q���-Vwjݝ���B���/s�v��>G{����c�g۶�'Us����������{�]���<�g���A�<�#�4* 竢�:؏�[I�=�ݞ������~�ޯ8�/vzA�i�	f�	���F�jа�U���Qv׽[��l�LŇ���̈́+~�g�.�R�dy��%��rܙ��e�byr���=��DZ#dMI�okH�,f�{���yA]l3+\R�wcD�h�F�b��Ac�cF��':�X�q��s��y���i�8����(7Jj蓨�v&�.���Nz!����ualL��n����lTl�7'%ku��-i�Q��Ϊ;��o�J���;/`2y����XXhİ�^P�V�
�NT	�Z^��",�;���7}<*&u�g��y�=��5�a��ŧwx^J=x�(룓qyKU.�\��B�mm�j�(i(�)Z��F�J�ZV����m+Kim���*Q)h[+JJ���R���
(�����[h)Fҫ-��-*T�pmDJ6�Z�lU��Z���kh�b"����UhR����)YZ�
�ؕ�B�#�*�j�ũm-cL�pR����[k*VF8�PV��Q�A���%���FZ�6���R�[iA�EF�E�-ҕ��V�Q�t�YGM��D�G��2�Qq��el�cmV(�[J��*�Z2���+��*�2�lDj�e�S��0D��8��J[K+h��TX���ZR��V��j���TQ�f5DUĹV�F
�f2\��iH�R�QWX\TQKF�V5�Z�[m5l�Qm(�eDJ�`Ԣ���҅AkbQ�h�ֶ��b���W�.2�m*%�X��ũU�KjV������EP��KE)e`�u��IR�KKm��J[j���h���us,-�m�D��b��I�uuj��L0��ZYg�$��^e~���������FO�!	6ZLEM$*s����VglmV� <ͦ�F�fԴ��TN۬��Ey$�UW�Cc����� 5Tz6��"�s�m�꽪������_�+���� \gkt@��Sg[�Sno����ͻ�T#Z���<�;,���ܧ�k��R�q���;7������v*�tD�U����l�c7ja�@(���"��L(/���٫���������]"n
jW���*��A��MN����u� q��bX�*��PKz�v8j�3�M�:q�[A�/L��g��5����>���| A��6w\��n�>�s�� ���I������i�鑍,�,T��c��T  �c�gg7+vS�3M�h+��JWyK�5�ܳjrB���5���|�K�l9��7����<��S_��{$��UDS^��"����'��H�߾���yŤQ�	��L��ؐ�ͦ�5���n���Ex��- ��SL���UA,5b:�wu�r*7������7:������Z�mh|F6�S��:���������8���@������W�$�Y�*�H79�M�Q1�V���!���2��Wj�RlC�K�*���*I++�"�ѳU��� �}��3���T�b枻씇E����F�T��X�g��uT0�y.P3�>^�{�q}̜H��ɠ)C7:��8�M�pD6�&���R���'�G\AO|
��M� nko�>���~��ǜʙ��I�)�UR^0hL!>�
|���o� ���Q��wuwE{n����t�A��T����Y��u�d6�2Π�nS�\�d�{��y�>����vl��W�'Y�O'"*�U+~SVV����[�	\�g��%��4{�	�n��:�4�����߿Y���s��V�1C�H�*t��yr�l�OW\F��aܜRj��r��3ێ��źi�\(7^����<�#����+�E�J*p�H�m�C�q���r:=�*fe����a�,����6�:vm�vrf�N�p�%��=�c�K���σx6n58�[q��\�]��:�δ�1ۮ �ΉZ�r�����=`4/X��Wg���z�u�˫�
<R^v4@Ztc�ݺW.2�g��aN�7k�����e�"bQ��u��vm?� �ﳟ���/nb}e߅��m� �Ϊd�v!uj-�p%�[¼{�y���Nݣj�W���Ā�73���|^���d��z=�V�}���L�rL�Z�!>�>�
})�wf6� �pͦ�A"f��rǤ��<����M���TI&�_L�,Cp� �UI�˓y�{���D�
�t�dD@�=���H+}� ���4�(�`]m�/@qڛ�����M��ڪ �X�nW���Cp����@zsa#8�nH>
�ci���z�#""�>��D��TY�^��N�-�[g��ͮ�G�O'�m�L2$�&��"��p�3[=@��:�[�t�w��2z��x����2�� $v�ͩ\d���J,��I�ْvm�c�2��Yto;XA�3{�O����� �-����,�w8/D�p��[�jLAؼ��D��b�ؚ��$Ih?k�ۧp������w��~�"������o�6�P	N�l�7��W�������@�U(�=PI$l���IA1c{�w�8�y��#Pi�ڒ >��QƵ4�0�1&7��՜��]�p�,$NP�[�u�7���׷^oFf�$�r��itZ�f���%�����������BUz�{ݓ�BE]���k�u���븎�μO���%�d�`��!B>,�@��	����m��Ք��qA���s�����ͮ�ع���>�nZH��Do��� �!c�7 ����`�X.!L�]"i%�6�*M��p�dѥ�}�v�I�Z��S�X� ׹T� ��븋A��w`Wx��EN��<��I@J�jI�ؐ���Ղez�*���3�N2����ոUa^���[�m�,��/nx�r��O"S�Ҷ����5��ܼ8(3`X�s�WN�\��$ƅ�3��~@ ����� >������7n�alA�m \��虬Iӎ&���Ј^���� ����"���{��3�C��gIں�z�&�p��	�f]�@$�[�(��8o��Ւ��]W:`�n�]�fw�j>��β��S��"�y�A�Lwn�k���q-����jx(�t==gI:�q�]�������nG�$��~Ho^UR	 ���U� �gN��)ų�b��0U������7���H@q|��a�pKqD�q�F|�W���� n�uݠ��dCA���,鋬V���������fh�3��Tt$�Y}4!b�e���r��nwuݠ�2���Д���JPd�SI
}��\_K���&���ݙn�> ��m�H\�Q�ɭ�<�ǂ����ljP"��t��N��^>W[#���cwj��ف&Y��v�cz�tʘ�B�G	��&��9��ΟI���΍���=�	*��ۻ�[\��؃�@�M{�7�m�k1�Ov�}UT�Rz������"�]v6Ȓ�� �u��A���߉��a����6��N�n���Ltc�M׎�� Ip��գ�I�\2K�$�ۺ�����k�@}WΘDu�-e>��/�70�I6~^o>C� ��K�P�|����gf�7��6#e�:8�+�|���^B����`yQw*{��N��$��r����4��DRA���� N�w������� �]}����7�&�-��,0��[}ֲ�U+}��I�o�MD�� /�~����E�q`�H���怫�g�� ��?�<�����wdGM�:Q���I�2�� ����@�w]��ϔL/z�Nw��/{�C9�2*Wh���7�v�1�X�,�ծ~L3��ۃg{��8.��ه���&	�d
u�qF��<��|>Ͳx����ÉȊ���7��[#�iz6��q�W>���u�fN�[��l��p��B�4b3�n�$�++�A�ɇ/]v�:�rTOkj�����'W�&{���7y]�7�g��.�^;WS�5k�ջVՅj�h�W;�,�4<F�W Y[q�8v����[�]���N��1�盄�8
C����si�on�ږ=Fv�mv^�ϐ:�N�\݇$�|��y�����񳹈�^G�h��vC%�PC�^g|��1Ci�5_���.!� -��Q���]�C���Us���&�封 .���,kT��\2K�(���K�d{\�ܔ�Ӭy�M �-�ڦAy��� ����L۬�v�@lZ�j�1�ȅ��]�y�g� �����Dvv$vD�qT�^i$�C]�W�U��]�I@q\�2�0�&���u��i�U�f 3M����wh ���\頻�ᛈ��Cjn���� u���Bω���xJ����w�RE=�L۝�w 6󥰃�Ҙ��E������DDx��6SF��K<�*N�v��):lq���WOmtD�nz1������H#���3���N{j�gw;�@ �u8a�wqde���)��� fouU����[�Ci�5Ek�8B
�`g���+cx�?>�q�|_�y�')g��y�V]�yR.���;�!��^Ͳ���R	���s��F����{�� �������>#o:[Oe{W�}�zdb�{O�Yk)��4LCAl�eѿ$O^k��I(�-C�طk�+B���6�� W��wbA#��漒صc�8pc��&U���8������R��뭸����B�쪋�}ꈈԀ�]�vR<<LJ#��J��hݷ-� �{��O�k�7�n�}�@|��������m � +��ٽQ�<�n�TldO&ߖ���h�� ����F�Y�g��9�L����KX�(&<�;��"0�E���V��ѿ���� \�: ��Ϳq��=]�rHI$~����T�,I����s�T�ӽދ����X �[���	
��C}���EMn��M�m��ֶb
���jJ��$��N{m6 �6�P�w�}?&�Ɣo�=۳���bq���Κg�����EА�����&�x�T�N��E�{E��eAܔ���F�,�{���"?|��~��@�W?����/b&`���U�ٗB���Cp�=Ť �ni���"�1�H�3��&峍M�5IX�6���sIb�b:pc���)�]��&�������o۽��_�@�L�S��
�q�� Y��w~I���*�H��n�A=��@%�{U�WS\;��Ջi��[�éy8է��]���\�u�]��8�1(��J���_g�~ d�4؀��n!eU��P<=Y�o�|��MR��4H�Cd���J�{nŤ�j.�f'�ݿug�� Qs�����$.�{����z�C��ˑ$D0L	�D��
�W����iy$�@��!w��f >]9�Q���v��N�2�����P�:�\��V9�T�7s�� fg��r4]u��n:�h�,�r5�	�3�͚�2���b���s��4��6��{޹�׉z�0/C�s���hR�T��#�	���`e���A���6m;� s=�׏b���#���u���΢�}}��v��uT.�����["�%��@�>1�[>dWu��M.������*<��n�PtG7B��|�?y��}�JzG�e�n ��v�> �g?4	Q��iWd�W�UUh;�����1\�6�D�4JTN깜�I��]�z׈�Y��V���n� %���	�%�-\=�3�&��=Ix�=��B�D�J ��>�۵`��:���4���W]�� ���A�uP/<��E�"
��	�SI
}�U�<��ԡ:@$��v�>�sٯ�| ��gDg�=���Uw]��-��̡L��#�y��c��s8�����Pf��v Fa�^��`��Rg�3��nX�\"�,%�U�!��j�ٝ[���w�����rh����0��C!�ѹU�.`F6��SE�>s�4Q�Рѩv��5&%�Tl�q�'eh�i����L�JDշE��N�ө!f签�pK��}�w�v��yz�z:x�8{�����anso6h��F�/U-�NF��ٵ��Ѷ�3�LS	һ����8!#�"7t��o���pC'[�i�`���]�`�V��x]���'|�g{������=�=�o/2oNo���͉�GQ��;�4�$�\#")虪���g3'�PJ����S�V#�X��xv��~8�zI�'���h�I�͊:��i
ɗz�3B��n�.&�Al�=n��3�{��=�l�� ��S�����O�?V����:��,��2䞅�ۋ*Ku��ay�3Wn2�y͝����%^6ef�2Jv�X,�u�S0�^����췈�e{S���ށ�{�䣭<�m��zuJ�nOv����%��oZ0A*��f�5)�](���(�y~8�r��oD�SN�ªCj�N�uElmnd���D��;Θ��k��ɋ��)���Mo9J��V?n��<t�箋6�T�:l�ᢏ]ܒ��O!}���o�����$�_9�}G���I�#�|�y�;�3�)]"v�� ������g�p�T,�Ff#��}�|zg��o4ǩ �K�-�����7U�Yڲ�8d�dO%5;�s�wa�ۣE��i��UJ�eEfV�`���V%�^4�ILD�E0E�������LS��VԨ�U�[mJ"���LsKt�b�[AKkl�V�"�V�up1DE�+m��*�kQ4YEr�iT��-*-j�ikqDĴlTK[kj[M4�FTkr�LK4�D\��J�[*�A�Q���F �M�cF�[A�����E��JQjTR�F"ZW�*�Jղ�,Z�(�QJ�չ�ke+*4eb�h�K��W��j6�[q�1q��V٬�EM-����+Z�����ӊ�+m�"�+ueq*�u�9ceJԨ���5�"�m�R�h���*��Ne-��[��j""�(�-����R҅`�F ђ�"A�#F�墎VR��eA��Tb��Q�mZ�QD[V��Z��)��u�5L`��al���V�ҵiV���ԬX,�ږajƋ
�l�m���J��2�QF�Z*���U�1G�+R��L�f2��+*Rڋic�`⨃A#�v����瞷2��G�FN`�6��Ka:+E��=q�A��r����+��7a��׎Ny����G����ڶ�֗qO�C���X��N@�m�%/C�R�mlOe�5��Y4H�l����c�����n r^��5�;�lb_v*�z��n�<���q�گnS)�gp��m�RRVz�h�3�����\,������U��@>��l����0�m�n�x��c�?L�G�ne3�ݖ��y�mۺAݛ��f�rZ�1�1���N�GHaɘn2�s�n��=u۝����8 ӱkrޣ!)g�ŧ�{�Jm�Fx6�6�QW*���l���uiGt� �`�:磧nKV������ñ�-��̧@r�q+�S�8�]��:Fs������ۊyͻF8$;z4����m�1��)��������Yקt�\��	����.+b��`�2d��,��N;\�1�v���ó�$�g��Fe֞K�@Q���MB����������U틶��79=�]Z�bۓێ�T���ۦ��pI4r9w�y��6�k���E�<��s<W������ls�W���r�q�%�1�u�ηF�0Bv��V�}}_V\cpg���Խ�y!�	c�Y	�.��A�Z�=�`㱝�7����[e��X�N�s�v7g� �����d���l)��gr��uv�`����wq6�.:6-�@O���܂�A�n�[B]�v�M�"�G�V�s�Ž:ۜ��ʽMCc��cm�;���L�Z������[=k�l��n�Y���bҥ�n�a��pq��������Q�I䱹��x����$�Wmz^z�N����A�y��^4]c�;%/�n�e��4on��ݮ��]���_U��[���ǝ��cmc9g�H�t��1�=����ʳȹ�a݄)�k���S'��sМ�Sv�q�`v��l�uq�����q��.�ɸlvsS��/"��0{=�`i��h����!�m���ԗQ�kF����n�x���G;n�D/��#��*���x�p��f�ˆ}�Unq`��z��"1�e�:�7a5���u����v{.6XK+y��͍;��';\��˭�q+��n�j���/���Ł�i��m���qt�lۨ)K��tE7C.��]��7E8�f�Ӕ��a�]�b����f����k[;c��k��h�m�9�i5�S����y���6f��y:�)�dz�ԝ���x��`eخ�ٮ��9/��wĲᄡ4�1_���]I�W���.{4��sz�'�0�����H�,٦��-X��� ��mU �ܼ7�UB֟��O�m� �#6���(!o���\p��	Ȩ�26����I��&!�R�wU��IOcM�%���f�;��g^��سj��A"-�MR@gv�h��N�����ٝM��4�]z9���,�����<����;�����KF$
Kp�����y�6��;��W�V��ѻ�����=�H���7��+��� fosq�#1���8�������^�^3�����m�16��s��l�����GZ8�>|>We��z���f6��t�6�ٝ�w���5nj�F���$ |,���e�DÆ��D14��$��ݎ�&b��s���������n�p�4\�,��%J���DU�\��s�7'�u�!����@ܑs6G�����Y9�O��fou�� z��o9� �6��)?�ԁ�7n�l��f4؀A{����� ��}p�V�t}$<����B�̦�>��n ^�t{�E�CD�+���VR��VhIĐHc��` �����>#3=�%]�d�UfBe�d�Uz�,��-��$C"��=V�3=�ׅywH�����]��3[�� ����#2�ͯ!��:���`*Ɂm�!il������o���t\3�q�<�'.Vԭ�XS���������!{���<���ƛݽ��� �s̈ݮ��"
m�rd�����[��[3�A�J�UB^
^i�z{t�)\����n ��I�\_��@	��__��Ԡgo߾`�e�D��PG�<Jm#z���Dk�m?�]�Ն�UC0�Λ��Ur�ی�B�7۲
}q�!#={�Q7�x.}s^�
���oq�:��єxbOo<�k;���$�W������MA�ov�� c�sk��Ѥ!�ŤZ��rz_�]�T5���� ������1ߺ��@/����t���v ��G��s	Y������ޒ"
G<�d0{;o\����{%K�- �q�������W�A�ʡJɦ�8b4�=j#�!4I��t�V��az�-�/e*b
��N�7c��ۭ�ı[غ$�h�H�4���Z^I%�~�k��=}��^��q>}�c#����E�{�9:�Ƒ��X�Y���������ۯ�^���w;Ve��""�����d�n9�ϳ��ڥ��14@q4=���(���i�"6��ml�,���� �w�ɠH[�4���,�a `4Xm�wq潝��h�"*7.�� t�:�`-��od�Ӂz.g�.�m�YH�_]Ew&3�����56x�����v��Onֱ�T���dՉɔnxxf��ު���dV�����q?E"G�j�qi�l�����p37�݇�\^�n�A�� ���1!\�SL�����@���=X��q����<�G!�On%�s��M���;fz]�;Z8�
z��&��LF��Ҡ�h��%J��Sj� .���ݛ�wiyC������kg��IA��F^�h�-��S[�tIk�=u�b��3=,�ˬ� ���{��㶖x�m��o%#Յ
d�
 C���$2�i����X ��9Zz*��}�$�D���H��7������U�B�Z 8�Pvz�#Bo)h�{����C���� ��w`|��#��~�Er�S� ]�����"d��yI��ޫ���C����G��:�˴���n��+����ן�xv��/y���9��u��O�D����IV�ɢv��l�
Q������ί�L��gc ?V����Gk|!�{����︌�~ ΄Q�=�GX��Z��=N;coQ��۵Sٵ2���	�<a�G�u�8%���FmʖI����4;R���ܬgnk�Z�vu�����O3sZ�Rìs�x�ި'@>�����4��>s�ѝザe�b|l�t��M�`���=p����=z��;ՠ4��u�V���Sr�/k1W'Q㝷H�Q�{t�:x������M���n�u�����.]�i�tVu\���:����ri�0���a�D���"8C�Q���O��ƛ> ���v  |�nU�6~�Rms2 �����0�i0)H���*��ʪQ.uaj�nB��@�[��w|ڢ"�ݼ���#��I�/:4a4�d�b�)���E�ST �Y��v\[�uM��u��$<{2k�R�$-�(��Dy:y]3��"2t}����{�� ����, ��W[��i�_$�����������P�A�JO7�@?����\uqc��b_}��d`|dm�j���m��q�s�F���X���=�P�^����]g��2�F�\�`LY��], ��
'ĵ��YĶ�4J�Xbc=m�� A�����(��tû��t�7��0��Ϯ���o�ڛ�bՁ��cd秫���L_u^��_B}ڲ�_�^�=ڼG �o��q����X�3��t��Bf\�g�]�����վ��tJڳ����4�U�'B����c�` u㖀�]�6��ug�^�n�za�q0)DG�@��tV[�`|.�� ���0����r��e�Nv� G^7�]�i����G��D�����������ӿ�\e�4��n���kۛ�w����@J��$���کC���B��҈�yZ� A���������v�ޞ��8=�KH w~m�I?���HO=�9����� .݌��pA���.%��[�^��-;Oew0C��=v�Aq�]ftt2�*h8��6�Y�m�4؀����v��Sq�W��\o8����^l�!~N�����R�GO;���K�W7wwN�  �~|�8I�}��0�vD���>I���׉�'lE\Z�EiD-X����ln�;� 	����s�y�=N"��]ٻ���K�;Q{�t�Op�0�W[��gq�H�������!�l뗽���s�K���[���k���e�6���w &\�<)�%J��9u�-d��\�oD����+�޻�>㣯d_��x�]9��te"%�MRFvz
h�e&AE����޻�����E��S�O^nx���t���n��#��)�>���7���|��Gv�[D�e�]�.�NI�l���]O"�"p�	az��$p~`���'խ� ���j� ��ʗ�oD��a�t{}�^��� ^��ݠ�g���B�Z!��L��T��z��[�b�ͪ�� ��m�25�5D#��y�T�Yk0�PU(����oi� >�"_��LR6on�� �o]�{N�joǹz}�dH-X���s�];�m�V�/ā�z��� }��r�">��q��t�W��ٜqw5�U'����巫(D�GzWk�蚾�ۓC<��Pe��/���	��s}\�ݳ[����ݤ������Q>�(��� X�})��̷��b1M�븋@zڢ �x�L���N�e��~������p;g�qqI��"�Gj�ύr����O�_oAML�(�g���6��)-={,�I$�u�I/[�s{;r��@$�\v��J@�H"���!� ��@�V��+jf��o�'��g<�v"�޹`$Bμm�|����L�:���}�Nxe�*l�B�Z!��L��P�I#��H����Q8����H����  Y׍�Hvm�a�a� ��PQ�Wf�Dc�#�ri��  ��*��w����no���ߑ'�(V��olE~Ũ"tn�g��.���� ���wc����<�Ԗ���IGu�ФIW۽vK�1�B��u~8���{�<.����b��+�:P��<���A�V@$��.�Ȉq��Fv��m�(��CHoj�?c.��}�� �w'RCq��;p�u��EԲԮ���2�p�Vb���XV\�"�,�H47�Yt��ѕ����f�v�xc�G�nI��=�c�h�ڭ�Yvl�N]㊻b4��=mu�g���՛k����Xü�c:�ɲ،�֋x�a��Х����n8."���p}q�t붡��\H��������\Z�l�E[�h�+n*J�E�P��,D�v-�sC�Y{n�N᣶n�n�q�w�p�&	.(_+3�L�I�ʪ^@��]��c���ۍ���[� <���I�cv�&�&J!�X�Am^�݇��nc��}n�� Fu� +�޻���&���Z��Y��)�HV��^=�O��:}Z�> 3{yݑ�:g"�̝S�o��4��,�ʡH��y��v�׆�)�����fz:z����!�r���k�m����whFF�ʿv';��D��B�T%�\��0�Xb�(ޫ�6 A�����1P��j�m����+:��3w�� ��o�'oٰ���p���ۜ�j}���{\uLѣI��"�S�1��:�/����?��B̄���.y�6 ���ȁ��h!���y͑>��H���� �������ZxD���Q��lV[P|����3v�;H�Bt�`�����
h���P�u�;�m�t��;�f�B�v
�c���MFIuۊ[jFL�W �H3�;+�����~r��5޺D
�w���F�7D;GRdTοz.�PG�n
d��(�S]�v��	i��t ��徊��V��Dnwsq�0��W� ]�B�dQ�ji*=:�[���Z<P /w�� &�K�� Cד1��X�6y$*���ǒ��R�L��)��=L�9�!�����|�5Ѿq�i%Z@\���@ ��� �0~��+�~���:[� ����t�b����S�xl���e��'%vW��}}���Kp�a@,1\�&���Iy-�{0i ��*_�����S��wa|v���i�����PCQKH՜����	*�|�s���Ȁ����q׍�g�:D�R}®�蝀�P�
p���=mI��t$ Z�u�v��3Mb��db��c~I�L�E�\�p�l8Ǹ��շ�]D5ɘW�f}���/�}���\��Ʀ�����A�=��z]�����3@������"x��y�d��#�	"�e͢��S$=4-G��|�;1����j��6��c�=�$x'��|p�-޾�+�H8�<�����SqE3׵�|�o�zd>޾�z�1��c��1��<Q�5`��u��&��ݽ�:G�רK;:����A��jBo��������䧫p�nz��t������U}����p�W?=�h���x󦼾��:5��c�}�m<��	 ��.B�S��Yy����X����G<��x��}�oH�O8������`�yǻ��o\�(9ɼ��yw��r7MM2Ŷb��yzb�p��n�@Ƨ�(���v(צ��i[�!֤i#�� ��|��`蘥�IN�����zA0J��n�����@�]�g\�t�KǦh���6(/�Ǹ='-�9Ӧ/sxM{�����j؏�]��k9ﭛ� g���x*�;���I�����V�\p�aM����d�G�`0����<��iW��zϡ�\�޻�ɡ�SܩUFΗ>z��]��p|��wlJU�6g����e>{�.����S��ķ}<��K�f��z�dI1[L��Hj���+��|����;Ϲ����#b�/n.g`ܻs�56,�VQ6�V�w��r�A�?,"w��+n���\{�nWb�e$�R7r���۳tX$� B@�ҕ8���Om�F��`��6Ī�F�-��,m���q�X�X���JԔQ*V�T������Q�h��ӂ�h�X�մm)j����IPDVXe*��V��JZ6�Z؊���KlU����(�[j,�h�Fڨ�DX���Z�TQB�%�
�+m����m*Z�TZ[Tˤ�ԌKJ���V��l�Q�̌(��[k�X�V��Qb.�QQP����\�j�mbԱTm�Z#r�ma�����fV�UkQ)]!F9j%�f86�Z�Bی��X*e����.��uk�R��32)�-.fecF������Pkm�mƸԭER�J�--�q��Y��V�kZ4���,�ER�l\��X��,
2.Z��L����0��V6�Ъ��.JZTEE1�e��&:L��U)Su��j��Dm2�ܘ�kS2����|�?�%�Y�MR�]�^���ʂ�0���{}�yۼ�4�>��LeDo����� X�� W��w|����	*�"[�A��H\�
"�
��T^���@���++��8�q쯽*�=h����� #!�9�`}y��v��f�nm�q*�<t(�! ��F<؄b+/n:�fN��Ha�wh.`,[�A����ύf�6�O�W�$M��R �y��Q�+�~�$�F��~�,��A¿���$d>����B&|J�yD�N7���	�}G�XjTȩ�Ӊ$K�^�& ����iw�޸���9x���p���p(�;W�T�$����j� ��ݷ�g�߳��[S` >:ct@�
�{�� ����x��	=*	�t�ٽ�3���(�A.35^�_ ��븋@|dvk��ک����w�SEnj���k��J��낝��F,���/_#^�L�=ۭ���~qvJ�η=璘A��/c�\"Ş|?B��uR�/v�&IE�� �D�Wuo� �f�T5��:����9`|]��wh�ٴ�T(����ښ�ߵ��:�ѱ>�Wpv��8�.���n�B�*�C%��$���!'��s��� ���v	 ��께���`9p��eT�J���IջPنB�ZT=�T%��2����ݚ�I� }���v����mQ K[s�}=�Me�Kʶ��[��
a�=�Ϭ �:76�� a�K��S�/Ϟ�����n�@��ٛ�{�+И*)�����{1��o"zh�\�	��w���,;5�@|..���1��1������ ��3p�Է.��=�(�����b}���)'2��H$����@�O�F�֌����5
Rr��9s�գ΃7\��Y�j�;�6 (��ظ�77*J�V���;'��"��4zKB1Fv�XW����$j j:@	b
���K��u��u�Qr�$�u�;a1�\�9�id�S��m��Z�ta��t��#����R�X�m�:Ɵ]y�_ ���2�l��;n����i5:��q�_d���a�C�;uܾ�a2�]�S'7�rE�����#���q�<ջ,/g�/-���Ѷ�.�ʹ��ͽug���%�"�����V�.l�>��P�Atѝ�����6bC���\<<�����ҳipf&��kt���4o�}�˥k�ɀX�f���Z%%��e�	$����E��p��A�I��������4ʁ�o��ubO���ݬ�.s��Fn�wU�c�dA�q��XD|ߥf2]>�w���:��^];��P�e��U'���)�KM^K&��sȜ�k_��$FF涕 f����eƢӈa� ������q�����Q;�� ��s���v�%t^�m,��Iqy��[vb0&"'��A)���ƝD{��ҳ���FvV��#�v�:ۖ��}��� �w]�To1�Gm�d�ۈ��)��<[������:�6��V��]��&z�O4v���~�q�0�p��d���U�R�I��d��I+��f;5���f/%�M������t��h4��_�B ��d�s�P�n�W]�q����^�GQ�������il=�\zn�b����I�P��{\�)x1�����(����X��>�7�� 徐�=�n%���%3�!Y/�a�
&h��n����n- 0⵸�V�����0�	����A$�}�@%�u[�t��[l*�'���6""�)�I%Q��t| >��@ ��}���]c�� z�_���{ҽ��P�'���X �co)�FoMo��ԛ���n_� ��޻���2;2�1Y̘��s�`��[_D%L�D!��dFde�ލo�u�}Ct���~e����A*�$yR� �7��$�N��㧦�/9c�����d�Y}�L�f����Z��|�|I#Y�����ʉ�� ��� ��۔ɠWD긡�wW�!r�L�т�A�F��g]	/%��%�h%9c�k�� ��~}�Ω�����p���7N��dn�O藐\��&ﳄ>�t�%)�O�|���ڷ���)�̽ٶV#����emd� ,�޻�>X{v�JA��~p��QS^J��gT�ޫ�C���A�y�����` ���Sj�"j�Y��.���wa-�y��0�naM*=�T% ��]1�Y�7w�ע��[]�wi ѻ������̈�UX�0Ј ���ͽ`�w�@��Ϛ��:��}q�w��gq�3���Q�O ��.�~KN��T �>�/����݃=i�=��Ia��f��و���b�1Tx�t$�Stn]f\��� �v떐 ��D �3Ax'�l��ߒBC��*%P� h�Zj�� A��� ���u��3�>�Ȍ ����l>�0׎Ʀ|��I#^�9��sWKېנּ�c]Ӣ �2�K@ >���.:��etU�o5�I�\�/N{wW<�T�������7���V�W��ƚ^lL�O<*�vt�A"G!��(��~$�=6�	H=��l��	��$��ܪ%%����e��ir�.;�(��nb@�ci� 33z��%�k�h��NT���Ӷ�oq�aܑ���kv<���nwO�t�
s;[k�܏iyӵ�����:q��K��T\�uט�`�o7h3�̨ڞ�#��2�&3j��^c0���-��k��#��ޭ�U��w��쮠 �4���A=���3)��m�3�[��1�"�E�$v��RH��ޫ�J�C)1����>��d� HZ����f�]�I��0b%m��h��U�޵:�e����,t���o]� ��Q�9�P�|e������������ϔ�z|(c6�z�_��n��I����LV ���1���� ��n�y�ұ{}�o�.<�p�MN�Íx��x� ���d��D��q<f�{�G,�[�<���G�/�v�ȼ���~ɞ��
����6�C�א �E`I-tǖ��5�v���Fkv��,!��Rv�u�'gm��r��m�{����z�ݫ�k� m��(��ny�Y��m>�q�T�=N�hl�!�La�aѸG�Ɩ��wC�A[�����\y2=�7=����ۋ��q��\""���$h�e��מ�Y�t��:M�(Q/�ti�q�bv]� S�+��s[��r[ӄ���*��.�<ݩ]�.���qө�.��r��3�k:^���o�����O��S�#�\���7G� ���j� ÷\�z��ջ�۬�w)��|d7u^�RK�ݽwa,�Վ���MAS�X�;��֖I�qw�:> ���v����tDD�v����{�g[��!�n �'s[½��2 ���j� �VÍ��g=t�n��Ԅ�;z�I��*�/kvb8&"�Kq��:6���;��C�7;" ���j�� �w���!�=��Ӿ~n��I�ܭ��$���P�2T6�,*,�נ�4?վ,�[��-���V��GN�K$���]�BS׏�3eg�{�~<�م뢗1���]f	b��vՄ��\uE���'��u������Sm�d5���s��q lv�5@�,c���ì��	@�9���]�I �Zwr�Jv�A�X�@13IQ}��-�%l����E�7�:?(����f��+I"��-�����=�@ox����Q�L˵�X�o�&D}�]�O��1�[#��� ���ׄ�$Ⴛ*���]y�WǱ>�"36��|�Ğ���$��w[tD6c��@�i*~�1wgo`�N�����O8��^ACqQ��_�YG{�-��Fî��D=�1f�u޻�*�8������f#Bq	��l�A���:�n�s����Nx��i�kr�H��������썙���������ؕ1Q#g�aKn�a�Gnͷ6
��U��k�ٻ������5Z犎6-�t C�:> ��������a�� q��ѿ���Ė Q$�M���D��3�M�J�|k:hJ^D@�w�b"3���@ .�]0+���
������6K`�*i*/:�RJK;������Of����L�3r��F��,D�ƻ�ђ�(Z�w��mV��t,��û����?��΁yo>�T��n�mY��/i�����'R�� l;�� ��������G�&`��U�Gz�N��#7N��x�^KK�n��@}y��v����}�Fu�%m����$��R9�4�J#s\��J� tf�:>�jb�g[c�C�r�@-�63��/�Z����� t<s���#���g�1kZ֪v�GO<5���oa;HtA�v�߿�2��R��ݥ}�tfct ��wa��u԰y7��D]�lK��|ٻ�w`/t^Jh�(e��OY8=)y*(b=;^쫌oS��ٻ�w` :3��Ey/��zn��[�0b^X�%ަ�%$!�E�*�޼�h�t�\ץ$���i�vFMV��b"v�|�@#�:�R��`�%��T�h���� �����h=�����6ܿ� E��SĜ���L�D�~"�»"f	[����l4�������罒��J{�m6b�1l�g.����]7���l�{m-�'p����;$$瞏M;�a�I�lq��� 6-�N�h�o�ۼ@.�˻� ��ζ�|.-�R��D����$�VX" 6ʆ�oS�=�Fڹ��t��$��R�u��+��?�u�	Dnk��9�$'	��s�$�-�3�h{�]=1��ݠ :3m�������x�Jl6/2���[}g�]e��wa�FnT��@l�tДIɒ�:�+��o�F���&�^����E��k(�w�- ��\f�H�][�@|���mQA��S/q6�$�M�h�U彙�9Z���3:�=yN��þs���뾭���6RԐ\g��R��ɀ!�Py@�q9�Ѐ��n<�]��F){y��p�\�?�;�Q�v�]ߒ��4D���7���89����'M���*;E���t�u�FcN�����%gt`c���{<hR�ޛ1Z��<�'�%�,���Uȼ�WU��vm{�nN����so{�a�c�z(��r�d�3X���6,X�+)��}�e�}����1%��������c[��T�4�rg=��|yw�*�܋Nܠn(F�eQ��k��{�r(��#�fj黝�����y}�����cs��7"˨��/�u����g�L�K�E����=��x�@G5����]X��>���u��=�<��!��}��[�ېk,��l���|#~��ld�;�|��@}�DS�U�Tǻn���776����#�޾C����Nu��Ѭ]ʷo5Gpj�[�݇[���;T�׬]��p*"���vD<L��T�X� d��j}����v/.ڵ����>�
�Ƌ�@�YnYsFn�x�*{ɱ�l���óc�?w����x�o>L���ͻ���Ks�]�8�[;ytf�"`e+�]���(�[��f�	��G�z{ޔ�b֌#���隧��t�X��gnyN�(��'R��hS����.�d�MY8���Ѻ$���P���M^䆗����_|��_.ξ����)I����Avqu�7��{�L^Tn��*j���	0����<��n��U˔?lzi�<���Ǟ#���)�d�@����yy�3��;i�n��u9���6"��F��t���	ӫ鼵[����N�f,:�fMq{����B�b!7^4�|B��>!$�c�Um�1J���U�����4��lS.fQ)�������b�,�ո�iLʢ��Y��Z�H�c��WYm���PWT��"�՘�5�Q�E31L[h�V�
�"��b[(5�L����2�"+��������,Zآ�Z"�n��IKK4�U]4cZ�J�S2��K-�RٙE2������Yl���Qq��YKb� �[Q[V��5�1jX��Ŋ��օ���#K*:-Z�5[r�ն¢8�J�KEE�DQJ�e�T[s[r��1�(�b��X)���h+�5L�Ԣ���)KU�[u��(j�Uf6TV�EU2�S��DHcV"ƶbvp'X�� `��vݷ�J�\J,-(题���5m�F��+�j�h�W31��̩r�c�W3
�bTY�L��YEfZ9j�-m��ն�[-�ܦ-���k&&�GV�+����N���g�v�������1��[����qs�NSq�x:��d�Y��I�f�>.ۊ���8Ѳ�g Ě�I/mŞy]r������Z��Ҵr���3��dqh؞z� �y����<�.y۶��n��mNM��aI���v��j���a����e��5�Ű����흫[f��5�iw5�p�ݭ�V�Ϯ����u��3�ō��3s�x�˷C̺���7�T�tX�l���eY1a����m���SYM�z�Y��Z�O=pY�9�`�=�ǎ<��Y�D�ʝ��͍�luQ����k��xΞ��6w6�q��t��=sa/j�m�ϩ�۶����m`P����\y�ݕ;GV��h��ycu��ۓ��t\�vsk=E�g����Uw�q�� ���.����.qG 3�՝��*��ӓ�z��:5�bzvs^�����u�m;��렟qO6L�h��x͙^�`��T�)j�[0sF�e�]4�s�:rQw�;�;ǚ�Ύ}�G'�c��n��u�s��#��J�'3۬��oll<�5��;s����]�A9maS�Q�M�v��]�<�*vW���۷Et�qd�[[��K�ɻ.��vD61+nĳуK� �q�H����]��l��q�7rrk���s�xMk۱��g����{�m7A�qsV؃{<v:x�q��c�-�tk̡nb����[�!͎�t�|Q��ۮ
Tæ��}Q��5�n���t�s�͛��:�pv�����t�b�g��՜����[��3bl>8Ju�8���s��7e&�ׇ���/�j��v{0�G���ܧgt��X�z�[�Um3cGX�t�n���%�*@����s���3���A��%m���%z�.����g���'U�ZF��i�{e�6�d;�^J���@����'g�n�ɮ��kL�އ�۶m��S�x��=�c����8.�ɹ�AМt9hg�]��nk��tu�����c�M�g�9k�p�r���1zm�+�u���]m���>�X'�e5��7;��7!�sv�+��^��\�`Phv�UUyG������"���zͼ��:�K]��]��E����읹Q�x݋Tc�/`Tڞ<�z�����6:�s��Ob�@\\޺��#t��V�{tV]�SY���\����ą���m�zp�up���h8^������øt�v�%<��`�v�Y5΄4v�
"��{IG�%J�=�C��ڠ�Z�b ���v��*~.���OT��$E���%1X�[0���꼣n��X ��󊖦�Q��F�V* 
<���2N[�~�~&�r*}�UԘ�3ђ�cvb4&�1Bh�T��̪� ���Ղ ;k���zkx�Vd�� >;��@,�޻�t<��J'ȸp E\n����цhu@�]+�I$��l �sz�"��n�(ۇ׻wmܙH����I�z�l�TCp�*�6�����ݦ�}�ض����6(@}�]0��޻���c�[R����SV"�j�PCa� �a$#���֝j�N�j�H�I|���ssA�>{b���ߟ�9�oJ�z ��NoZl@ ���v ��{��O�d�U(Yg{6�Ö�π�o]�@-�;�<�|J�(��68�m��'���<";n�(�Y{�j�)F���ӗ&uK�j�b�V����$Gy����ܔd��8u2nw��R��a&�Z�{����w`i�٩Ey$:.h밝u]%銴x2�x���-��W�vDF����tWeE~��}��o��_7�	 ᧷j�%!mو����!b����k�Q��x���Y�j�"=]�����Ӥ��HmvT�������$�I�������8���n�x��Ny��x�����!8G�e��U��`@>:;u�DCB���L����m�׽�}d]r�O3f�&4&T��Ӹ��Mv�y�8;b��h`���&�$�n$�8#/�n��۴�  �_c��}��VD{s�yV㻻���ݦ�x� Ⴀ�3^HS�*�J$�Eپ��U�]ϟX Zn�� ��� A��O{���^��@%��}���^����GuVP �s�i��������DL3���Na&l ���G������A؈�blD2
l:��\�}�C��$t&L^���K}�$�N�Hq�������Dw��n�Dk�m�<8��(�����=�}g��^1�Ӑ*&���y�����r�fg�8�ĉ:m��/kvb8z}��)�[����������p�Z�����69���.{���>fwU_�sً����[��F5���9��y|�ͤ�����n-��[X�E\G6�E���Xm�x.7]T%$�]�6 �����^�!��ka��y�R�	 ���T�/q6����Jb���ݫ ڼ���+.�P �0{�Z �� ����ۿtz�qQ<��+^JgҠ�AT�8�֝	 ���X  ��O��cce��2t ����6�ߤ����U,Ha�7	I8~�T��W��Gm�B �����������uD�'�SqDJ3�qN!��2+�-�6��<�q�yw��m��ۊv�ۨ�[�VS�w��-Қ'r]���#5�$.7��
�I=$�{�*\/�Y|�N��m���P�4������ ngsv��,�	�������	��`A�r�����ܬskN;m��l!���Md������#�j�!1?���
�H%���b�$�]�L����#�3��E��J$��S�+��A��A1F�ۭm�]��q�����Q\��ݧ@�3z�� ���M�����{�L�:WQD���)zf�l?��iTR��۱h�F��ɤ�k6*�i[ϝ$�
�;�� �;u�{�BjR�����3�%E�����Ʒ�&;���h�����Qa�8�ʪ�v��b+�$�F�d@�!8,%
�
_ 1��y]���"w�ݰ{y�v ��[L�����L;��^�6�.���o{��\(K�� �"x���QmT�z�=Bu�8y�B��A�C��C�#pOO���5���j�*�0`@E�M� '��>ٌ����]�L�of���UڣL�obN�5��^۝�R5�g�����z�m��)q��\h�%��s��ѧcD�;bq�W���mq�F㵮�>��Kw��K!>�4m�8�[�s�v���+�>�Vv�ǘ��{�q�۲�]�3�٥���ω���E�u��]���l��h1\<��Ż"�j3�]��t�I��[@d�F�Y����aR����3��cv�3��~�6ʂ��_�ǯ[��[���`��堛�Gᐥޙ��d��������<��QP਀�&*�㷒���a<�m�_�������須�����b�1ۼ+EFVn���uu�I�&ڄ�JT���pж�:�A�ו/�d`��x���e����j Y��� �����1}�~*Ce�QJv�����ڽ�D�몈����s÷w��I�{���u�	}y5�O��ĥ3�Pz �`�k_Ώ�oo;���<P���րJ&n�4� ���1���v�/�dUG�}V
�D��@�{Tɝ����v�9�5$����[[u�xյܰ���A>�A�x|��cm����ƝDn�7`��W]���������(.=yT%5X�'��J!&��7Y��/bg^����b�^�f�?��V�Z�ۭ3�)��`L	�\�R9��ȗ�Ő��{��o|��y�և��LY��Z:'in�UG >���h v�]�D(�=���T���ۨ���XMC0��bI�9r�Է7z��� ����nqM��oݕ�񑷕R�I_n��1�;jE8�T��Ko-�^[����@�n��" ��w�� �z�I��q�8��yq{�CҐ���n����*����Qԉ׳%wL�tV(��;�S5L�	nn�v Y���I^�F�j���V�w�y�:ک�0�]E�p����͛kq[���i'5�8�������`�%l�J��P��A�����@|ћz�����Ȱď��A��o��HIt~=Q@ �!DB�B�z��.{`P��$����^��Ѐ�w��",Y��� 3 `��Wp�]�[�N�O���I�4o<��@�w)����{�L�C��c����)g�Y�~HZ��k�pF���~�#;�!��g�s�F=�W�1J5{:[0�����HT��H6n~<���p��ڛ�� �o]��wL�l�)& 80�M1$�R��8�q���� :��`����q�C@$du㽄a�؛����}���e��J��@�O�ވ*�޶� dvcN��B7���I�W_m݄@,����L��9r8��ە���Z t2P�G��;wl����q����k/hF��]R/9��x�v|�ngCp""!6�W�ۻH$�۴� ������EӿnF�{��Ā Yۭ���/E�JI��43�KA���C]�V���m_[ϬAG{v��I ��}�ɠ��м�^�3$9x��+����Dz �>�ǆ���i�	E�4� �����fO�ՓؒH��ɪD���eW��"�)�%��$�k���۴�Y�����x��]7��|�#��*Z 3���ꛍ�:˜,�*���w�xtَ�L�
n�r����~آ�E�Ż�d�rl�`����˙����&�����vy5��iA�'M�����^�s��u����N 5�1$��)$���U�hč���6��H�����(����b7LbQ�����E�lĽ[�+��@�ۧ���؟M�p����\\n�߿����E�aÈ%I8jvxJA$�w�*W�^	.��� �ɱ�q��gi�I�U��K��m�����E[��~�af���nc�������j����� v�sq����QQ�~��JOJDM��iЀ��w�� ��c����*q  2-�* A����$����$#��j$[���ѡ�{�3�|�org@H6'y�Q {{���H辶����R��|����"޶�����[0�ê��}�~��^GE��T8��z+q8��wS �]��wh"t_[j�IO;G�S�x��^{N�7�N�@��j>�S�����]��wp���<B��d3�,g_ ����I�ׄ��{�w�d�]�x�K��B.�Ճ��I��;�]p�..܄�Pn7i�ˠ������ܛ��]�\�l�
�ضMp���nú��g���h۞wN	���C������F�f���g>Q���rk�cGj�uG��5ۇ/nq�m�yn�v��u���:�N���ۊT���'e��[\� �q��8�n]�Q���j�b�[m�4�8���8;��z�έ����t�7:Y7R���NֶM�n�,R	����oo5F��e�"e�'M]��p^�� q|ܿ�nvp�yU~��wͪ H�޻��+]�J��A*�yq�ʠ%�r�iu�X���'@Dgf�݀:/����}�X*y�;w5)K��m��B��h*���۴�> 2/�: ������O�-��I�޻�$I�}S^��X�E�^��Θ8��{Ue�x[�
xu Ufk�d@���` ��|�7��::/�_3חv���Ƽ�^��l��Ѿ$�O�o��	���|/����˻@$�z�bE�o�%%4w'���	r�&
��A@�֤!�"�����ÜO>)�f/7Wey��������Dyz�sYwXFE��$@�V=�P<��(6�;w����H$e����m���L��Bl�T�̯
���&�Wq�q��=�u�_"�g��Im\��)6N��;e��Oe�|��FDN��\�9�Ύ�sB��AЏK�cwb2ډ��=�u[��j� 
6��D0�|��q����533�X��Kj�a2\8�T�9�L�I�S��$�Ui�)�VV�� ����" �ȷ�a֯�-�E"պ���������H$�Q��W0@ż�av��߽�����%��C��TC	
d�6�]���ʅy�������@c�Ԑ�o7 #�8�q9���2Z�KI�����9��y�Z���uy�o��t�t��ݷ�o�9˻>��\8̶�m�r ���AX�3.o��W\���T@.�ͩN�f��E��"�sAs�˱i�Mvx����^�8ǵ�}��� >��7���/$����W�(�;�����#�0�MG�e����eSI!�sz��	���[�."�̩���KE���|�>����:0�uC�u�����W�g�u��,�����n������U������rE������N���|�.�~���{Q�����5�m�F��������|�ǎ�o'R�������<kT^�<{;'�f��w�wIv���+�?7>���j���lG���eInjg�+�g�	�oω}�;���m6�t������|�n-C^����3��|&�m�o�ؼ�|����g���C�a]�r��?;����I/@��|�-op���0�iT]:�:��;u�e�σTFn��H.a�䈷�M��݂��3�gr؛/r���eD��CI)z:$��,6y�Y�d�=wG=�3��1���~�7we���^D�,g��Nb��q��;�{�ϻw�o����-��ݣgD}�8'��}7��}ES=��C����{�x�F#�����P�M�1���7=�;�|)�oU�|���y�(�{ڛ�� <m3Fv|ທ;�l>����Y\W�:��Y���'f�\F��$���{yN;)NI���Cf2���/*D]n��7�i;-NЭ(�2�-=A��̛��Y�wZ�N�2�fnBݦ�+�ƹ����hS����ofp��Џ1c��U5��͋��j���j�.��ܞ��/���R�\��m'@R����Y��vs����K�H��N<8���s~ؔ<���]���j'�'n�=�	-0�������8��{w�S��4��������gwc^[�[�R�R���D��E
��pJ�[�2�1J�+r�P�hUmV�5��&)r�L�SX�ۍʆ[1�c�e���s,�q���Z�R�U�722
ٙTTal�
���V����J�%*T[1s0���*���Z2��E���ۂ��m�6�!�N�nۃǌ)�3)2�əJ""����GeG�r���[V֕�qȈ9J��9���0����Qn5PA-*����iX�7.
�V�\���0R�LAE�F0P����((�T2��h�q����iQƫr��K�k�U�iq����\r�"�W��������d۲;�Oc��0;���v��9Î����9q�-U`�q�%qm-
屈�"�es�1�6ѕ��6��ɍikKYR�mU�\Jb\Jb"�2��W��n%k�±�b��r�"2,�r希��C-��W�-K���Eֵ�s_�i-��U�A�J���I!�Xa2\5 ��/*U)���v�L�`|��s|��� ���m:��2>�/.0K�-gU4���m��*�;�ժȀ2/���5WGY��] �}����7�� �辶���ү�9�?�߿��S�m��׌�wt��X���79{Ht1����0DyS%�X�-̨a ���%VV������X$ _[������5�mvUy������	X�.��������=�7��O����
��*\�3	$����$�@��9� N�����4����h�R�S��무��N� �g�mH_d�d���Dg�}ٝ�v���l����1�d�x�1D�,���_�_��]L�e�L��� �����ִ���$��7����揄?ۓ�r,o�CŹ�L�b�9��g�wJ��Ot�j�U����;�'��*9o���:?a'/wz��@�y�L0Ul�Ues��9���2���nS}wh ��� �,=��i�K:~�����Q	.��j�˝�P4&\Rx��$�6·nǋ��F!���m��'�[_f��_�,��� ��s�ٍ�cwW�.g�w�v �o�(�Y���0zP)C���{��r�Uv�Ug^k�M���w���Θ	�W6���հ��G V�ĕ�4`��M ��؞�m�YX�r 'y��p��"R��T�(���Lf�ٕ�A�	R��w׵Ӎϵ<�) 	��i� ~�~`����dF���^�{p�~���'2(Ҹ�պR!�*��̡RJ	^�uQ�P3'm�7Q��FK�Q���mQ�����MŜ�1/�(Km����l��]�;�����z�gη��/��TCV��_=��]�1;w����7���>�UK�_U
�٭�u��@��-�C��Av|�I8䞴�:챛�K[��ZH���ͻ�tX������l=�Î���g�͕�q����W=]k�ۤ�&�b�+���\<�^ţ��z#����r��-���0Z��<`:{Z��h�qI���'؆�c�[�<���������̱e��L����ۡ뱩sͽ���,c=�p�6�/;�X���v{6��R[��������=��h-��5�D���` �-Z���r�9�t�l��p�I��ܪ��Ia������n"<�O5�2����aI ���P�����I�pE =�ۿ��v�u��/v:ߙ 8��,"�s��� 0�k}���F�c�fJ42���v��" ��#Lؾ���S@ t]cj���vM���Q�,B���+k����[�eJ��R�D�7��� ]uUm��s����$�-�ؔ��/�a��&R�w�D�GS��I�<�� I�`%C�s���7��/��\�L�4D�����s�Ǡ���E���E�����jk��n��m�4�F������s��j����}�RI7��V- �I`�;����[5�>(�z,,7^�Mvf�݄����0[%0\4�TH�9I$�Y�!I�(v�a�����*�z�:|�ʻoI�#NO:����O#v������ͯ��sg8�E��_%䝧����˃[���%}��V��H���Ey)�r����җ���Ce��A>����m��  Y|����?z=[���6�@_n��� ���
H��V>L4C
��������W{% �-���e�t�@"��9��+�;����ۻ@+Yʜx=�+ǽ�
��g�6-��з6��P��'3�=4��� �����`"��UJ���\�� Q
�P�`3B��r�n���C^��1ny��p���|���߅uz&"}%ME���V [z�H >��9h6#�Ӹ�9�뽻���u�uI-�Q�8m@��A-7�.�Jm�^�8j�t�<�|�4 ��S&�EZ�x�u��Om��$��`�`�'�Ҡpж�C 2-�N���G\�N)�~��S��V�>XAڈ�x�cO��D�Z�d@Ɂ�`�I��_n������Q]��������U/6�9-�uQ��|�R�!��"p�QJ���UgIu� -�ڨ` ط�1 ;{��uǽ��֮��=u�]��`�\gũ���$)C�2��!����v/d�\9�GQ&?��*��`|qo*b�.�o�����4�Q��-mU3-�\3�R�l�-��9H��ڌ���۞e�������?��������;�u ���4�A%���v�t�{/#bF*�=�	�u�F*�jl�%�	����'�X��O����舅}o�w��j+s�xoj/����(��8m@��u�P�H7��4 �����*�-�'ח]T�����h��	���U�yy5���f6��@�}��@�H��Cu����ѷ�)�Bnj`�X�ћ[3�^Cs��ɝ[;���M�l̹��.��^�B��9�@*aW�LPSZ���f�S՚�fj�5��۹�D��̈l�I�\8����uW� E���EZ�gJ�Xf�X�uٕD;���	umȝ�ܣ��/1Tl�p"#В,�� ��0`6��M� lf�WLvˎ2Q�F��v�ߟ����έ��������N�wH�x�H�m��Z#:����i�O*��/;���mB� ��Q�7�>=w3Y~=�UM���$FwwP�@#�m�5��.�켃����*E�l��&��P�꺯|H#�.d��N+7��g,Q{��ۻ�^$�:��H9�Y�f��{,C{n6�';���A��� �.���,��f�T�L[��'�V�,0�q*��s ��Aʺ��T"��.���$wm�Q �GV[H����ү$h<�É5���������z;�d��j���|�_94�oh�vye� ��0x��yW4yW_���Im�:묉"P���x#�WS��lK��I�����7B,cY�mO����v^�Kh=q�6�v�P8����z�+;l���qѬb6ޞ�泸��u6��d�Wc�oBt1�6Ͷ0[��:��;��g��/F�ё=v۳k�6R��º�E���x{#��=���㛃8�ӡ��Ƅl�o��o�.�]�۷��t�la��]�͞��Зdy�9M��ѻ�I{m�V�k�ɸ��BVׯ�.
�M�_������D�È	}=Y�(�u�2I ������
��z�tl�xH"�nd���z��0�,*�9s�D� WV8&��k�1�5�H$��� �E��Uxm=@ɧyXW�O�a�>�QH`;�q$���Ω��N�VP�	����s�%D^fܬ޿o�������r3b-�	8��tu�n�q�����	wT�$�յ@��ۻԮ`���ȝ �Fm��H��ކ�bbN�fP�M��H�]o��"�v�H�f���I������Ox�c��d9㜔e%�m�p�6�{]���i��hغ0ku\%�.SuӍٻ��������8`��F�s�Iʺ��|{wzDO%KA~;F-o��o��� ��R�@E8M@Jgkz��ýX�b��zD�^�ʧ,z3}/5������'s�C@�.�鏧��s�q�c��
�q��x����e����I/xr������}�w����T	�EE{�Y��[�~����0�L?&P3�;TI=��4I&d�!a�[wv�N��I]{B��n�U�-B�!&���'v����smN@=�@Q� ��ު ��vԹ�b���ֆ�2��"���m&Ä�C�U��uD�w>�Z�J�Ӑ�$��}U�A#7��W�<v�|�gI������� �AOy쭣n#�J6�"��$�T�S֜I��؋��������<�r�Zۀ=]�TI7��4	 �[wEX�0Ђ.*�WUI��CT	�Ⴄq��q��7�/^���9TA$�v�
�x��{Bpg�$l�d�"Tw&�h�I�5)���A&��� Tj��\�X1Z�*�3V�B#2�c��޷�n���A&���*Y���2�pS��%��/������UOw.Z�^d�նN��7m�s;z��O��z��
	�����	���Ooh��ʚ�$�ˮ�I��ޣ�'��6#���ME��@��DB��'���v���z𧰽U�wU�|H6z�����5�&'�tꋓ��!4ಁ��=P�1bQ����8E9u�a��:��+���0f�i6E�1�[ۺ��9w,�I��ꢞ��7]=fof1��u�TH'��]ϙ�Ȣ����!�2v���X�LN�ѣ�}����I��$7U�U�A[u]���mz#�V��b�CE�!�ոg��o�V��`�e��F��gh�O����0@7U�4	��Gbm��a���ާyby�k�%���U�4H$gn�_���w�:2��0sl�Si����8����{��N��dR�;xI`��`*�`o��z�z��b��n��w���G},��<,a�0j�㽡@��ޟmvzj�^��8��$�H���Nn�UX���{0���u2₠�х�@�p�l͗���Y�`n�զ�9����Om��|��G�1	p2o&Y$�V�� ��ުjtq���l��$����U2s����Xpي�$��}צ��|�2O�U�T$��ޯ9ۺL�o��n�g�`U�ABnB!�d՝�D�{��@�	:^� �u=ز��:�	��U�r��a�p�0U39mw9�:&�A��������A��g�\j���<2��X�X�`�٪�BTv��d�ja��N��W��g���>�Q:�y3�߻�����=�ȱ���ٯ��$��H@��I	O��$ I(B����$��$$ I?���$�p$�	'�$��	'��IO��	O�H@�~H@�P$�	'$���$�`$�	'��$ I?�	!I��BB��rBB��$ I:��$���d�Mf[ `�m~�Ad����vB�����\|� �  �                  �           ��  ��  ��
 H�(�R@)@�� P (�U(AA ��$
�P�Ͼ���%$
R�D$�@HP�TUP"E�TJP�
�UR�B���IBQUUUT�U)T�R��P
*� kZ���
*�J�*PH��n���w (w`�s`(�D�t݀�����RIwp:w%QN�݀ �@  z	��(�4)�y��BA͔���� w1�Ehf�)Gv� ����`�<�QAr�R��q��E@��Sz��@hEQ		H
)*U�)!��n`�@�aЗ��`={�P�J)�׶�i]h=�:)鸌W}��>�F��b�q���Z6Ϻ � � ��iQ��ʯ{w��F�����"�hP���TL|�[kB���^�v(uZ7�{ǣm�X5����=V��续���4{��|���{ճZ���i;�q���׾�z�lj�n���e�[l|P �� (��T�EUPHUTED��Q+W��U��y|G�NG��]�GGl�}�z�շ��W�ܯ>��y�z������9]���:G�|��w�/��3���w)	P��| �S�y_}wIG���:#�|>����FX����wUOcW��*Oc�@���/��.F>̎�q(��*�}�}P   ޠ  �H��PUDH��
�D<�����;�R]�p�b�R=��I�!'&*(w`r#�J���%	[�*��T���݇P�(QA+�E >���R�m�1T��$s��	��U�
E�TwRp2��� n�(!���HH�HP(w�@��¡ ����)JTA�@�1�ݹ W����&���z��ݹ����iDF��*Ku%)�(9� 5J)@ x   Ʈm;�Ҭ�à[��Pr�r���
wI��de@=�pJ7w
� |>�       ��h4��R1410@��0&i����%%U       OF�Q��       l�$ĩS�` �L    �	OD��R���     "	��b1 M4hI�l��A�}?����~��W�5�d��WS���\����5xIɓ5�}���..�?�P~�T���U0"��'�*���PV�)�����P��EP\
�W������O������3�#��q�=}����H�Ң*���R���{�UT� ���"�H(���?���y�`��/�~�(#�o�����1𻻻�Z���UU����UV*��5UUj����UUb���ʪ��U��wk�"��� ���(b*��� b !���"(�(b	�
�"���b(�� D� ��� ����b(!���"����b-�A1A��"(��b
� ���b()�\Uj�" � b�� "��(b"�� �(H(� (�  ���b*!���" � b8�	 *� �
���b*	�*� ���(b"!���""�7WA�b !��� ����b ��*ECK��b����;����N�����E�Uj��UUTj�����\�?{t'�~��[�ۧ�(��A�ȓ�Co�G����j��v_?|ͳ)aEY?7���Ly��?n��{�|��
�5U���S�5L��P�[�Zcu�[�y��0DY�?ʖ0e��q���!{���;X�[Ÿ�م��*�h�mn��?j�ȨUZ�i���cN����
f����N٨�L<���fVͬ��j8/2���7m3Zٛ��Շ)�w��/)��d��d$�n�įF���	�j=����'^]^�$��HX�`<Q��(��ck��ә��C[L���'18n�2��GLGUVh�f�Sۆ*�2ƻ[,����H�tR�Ks3�hV!W��� ��U֜%�)U��:n�!O��"��6ڧ��"�آ'\T�&ɹۺ9[ܣ��X)�z%����q�Pò��Clql��+[fcF�m�%�w���J��o[��jF�/*"M�ii� 9��^dyi���){.���WPlIj�љ�f���ewf�^�wh��ø��kE�bӹ��5���ǆ'n�]CX2 iQ+̓-���+.kcQuq�i+r��S3H������)��'�0�����n�]�)�m�,�6�Mm3�2�+X�tTF��o�hש�18crJ̸�d
��n�]ۇ
r|5Ltd�+��_#���;BJ�r�s�(�b�p��������6���i�l�CU�}qˮ�H�N٤L ��c��<���"�f=��3[Pj$L.��<t7ov-p��y���QV�.�z�����wE��Nb�)�����^v��E���l�8���ձY7,,(a*m��>��j��jU��o���I�+m�ERl�� ��J������r8��-5u�eޫ5&��v���f]���` ���E�&�4UY14��-!�֒�t���st@F��rn�' X8ݙ�f����iLf֣���(volۧ�]KFT�uȡ��Ii���ٽ��n,J=�VT�Rd*���m��<���[��`I���SAV�cu��anŧ�
lL��DRk�u�n��6f�k/76�����M��t�w6�
p'L޲��um�L�(d���c>F��)ۙ{`a�6R2�\ج��;�7~�8i�T��+�
-���t��nX͙	��$��ڼ���M�]���3����#����ʼ��'\�����0��Z[�v���2�ٻʙ2�5�X34 �QJ�V8����,�Q^*tP6�m���ڑ5���	��G1\yP+T�wZ�J�j^|�M��e^=9�0�h��$\�vE�˴��װ�Lt�R;I��Rj�v^��J!d$��E���ŗ2����W{r)�/a�T�����s2���3.�4kc6KZ���2���Ҭ�[2|j�Pд���d;H,!L�k\�����2��P�i�mXv��.��+*QKVh	�R�7@ʉfR�!�ܶ*�xB7�A�1k�[�Uk���-�4΄vd���û�LWO&U����w��m f����Qt��6i0�R� q��t�s��#���z&l�]l�2�t�$��	P��y@���x�wYz�ʄ�W�X�e2ł�ŵ�U)�N����P�m4�^hjdYn�E�J��mͼ�R�/Em��g�˼:�����4q��tذ2��1Ӽ%=�h �z���6�e�U�D����Kw�-�	�o�7k�6�R�זU�q��pܔt�u*}�{��I�j�u2��y�q&w.�j�/@JB���חy�J�R�n�o̊�
9V�cz7�*ؖ��-��3v�KQ�i˽
���웢�yq
��(�����o�"!:�l-���&�@���c����-�h�����h��@�����(VK˛����@z�x1��2	Xo�y,����l�I�C�q�;sN<�2��c�)Y�qY��=Osr��5��; ����X#�jj�WJ��Yb7��By&��en�l�(�%��ZqӴ�<!Y���ww:��j�M0�+Kyn�Xa���������cŬ���,ޅRҘ�EX��Y���ܲl�y�v�m �����R�t.��wW���r�*9����kFޚ��!��ڳ�,)�sY����k+IX4��eJIQ9�V(���-P�X~����Ӊ��&��d�c�u�р�;X�e�#�T���e3�)bŋE�Z�<˕�*�y�F��h�cj���;��j�5��-���gE3��߃��VBEL7v驼ފ	�Wu�F3��'e41Q��R���{K��%��Z�-�][���p��
X�ek�MwG0��3cc�ɶ4-�{�]��ed�� ���O�*�D�����I|ΠZ�� <��fCoᕂ�@v���ma��3F�Q5���?7.�ɑU��F��t�<N-M���[�#vëݨ�������a���m�U����ӱq�0v�nY�Lި(��uͬ$</EU����FbZ�'Z5��b�Ah,t&Pek��Pf�������w-4��84��fm�+U)�L�P1/V:&�)����;z\T��7��T�L�0b-刁w�f��u^B�j����t^B`������1�
n�ͶPڦm����'h���֝y�me[�S(�7w�4,�e�����F�r��B9�iu��f'��;WsL�4�ۺX�e]ZÙj�;N�R3^�ذLToԘ!�&Y�;�VǓw`�g]�`u ��"�l�H��ˇpY�"���Ce �w)�r����`�a'QWW������v�E1�w�GM-:$�,N���b8MoI�yP8��mq��n͉%/.;��ƫ�JS5�&ou��՚g�;�Xw�{��"�6�o����۶��@m;4�e:��� b���N��Qtlm��X 7%[I;�Q��1n˼�#y��Z��6���V�V�oMC�z��XG`�wS˽�w\�>�M��Nmar0N��-��߅M�whL��b�ɖ"cn�2(��1��Y,���i���H^<o_�Td;{�x�K��[��ӥ�U�*ֳ6TX+c��e�%t\��l�r;��y�X�2�8Q1P2���S`ҳ1���֧��K0f�(�9�|�[ M)m�,����JR׷{�������ѥ����"Hhq���"�oً����z���N)Z�7-���+�L��K^F&�	B���ܕe+�)��+7Vշ��f��1���Ǌ����ݬ��� +D���^ʒ�V껇é�튡K)�T�im@���]n��,TB� ֘���y2,ZsZ�a�1�dfZ���)�C3UCR��Iܻ�D�8�B�;�*��L]�T�2�ه+U
��LR�y�5q��Z�Jm�{�%�L���y���j-ܼ!b:L���yHVH����Sv�6�5Trj9{�ݧ2�B�m�x���a��vA���T�V�6U��șI]Y�FDU�a��Zߐ���fi�B�0]=�r�c���P��XLxJ7u�ݕh�I@��������AQa�ʺD\�H�Z�A��y�^�2F�À�
��w�����%U�183]u��U��I�Q%۪��ED��ĀW�$ލ$�T���X0����@JYH,���d�!��M�sM��3Mk +&圄]�k#���2S��+>U����F�]k�C@�ڬ�2Hn�yPٛ��͡�n��󪱁�����(�^H�X�����6F��J���ͰFC��ܣ�n�r���Զe�H���NnEn�����N��ceֹ�J`��i��a=ܢa����v���8�i�ͫ2�RP�0e�MU�ę/#N �)����^iCQ�K�.�0��oR�.�G3���uh��F�[Ke;��ɗ"
�X�(3Vk�.��c�w�p��+�b��VYm�qaA���aZ3h:7��zس&n��ՔQ��3�;�mk�gE�c7���;WyR�Ai��!Y����"��7�.H1}��`u��Ӄ��cOyY5�Z������ea��y�[��nެ�L�	vu� ̶j7���M�G/����Uhֵq��̻7q���h�۽�W3hfh��-�Xp���r�9�&ἳ�"!J)�$�J[p�	�n� �%��t�E!��f-����X��ه]�c��h�r���(�n��ѷXbF��5�;���<Iٙ0V�36��]���DG)�X��HZ��d{�Ԣ��W����˖d���LӺe�ɺַ�����F��,�L�����q�򔩠rf)2����V�b�����5l��,^�gY����:�^?��ot���K�V[B�#cCD���5u�w��PG��`�����]=�g�Z��5��L�[ -���-��P�2������`b�|�"�U{�b{x����Ż�F�{z�Ɨ0eZ�[Rպ�v5�Ѭ����EP�mk�j�*�
�Ǣ���,(�kE	��b�ͽ�+
O)b���!���fб���lm���*�CQ2Kɚ�ٓ�1�q��8坌�%�0���;�ۂ�i��.�V17zK
�����M�+q
C헦m���!DӒVs0nX�4��)����@�n�[�f\��U����Ԓ���A��
�{J�w��Ù������^4�-�.�G�Ҩ�-�9s�3vc���u-a���]<�W[|�\���۫sA�:����돭�ŧ/vh8�)c#C��el�N����-+ڰL�"�o��u��R���#��R���jƇN�zpH� �5��-�7.au2����BTF�."���.�\)�R���휟g[�U����P�w����搨��jj�y���L�
s"�
i�(d;�j��1�y�%���-����C�-�0���L��uơ7w(�u�j2�F��|n�6vᥢ��V䛺&�h�fS6�e��5C"�V"(i�l*�z t����N�g�y@9@�9u�5�Չ�X��G	�rlwx�9j��b0�*k��KX�3�n�3g�ЭYA����D���P2�Y3K�@����O��Gf����Pˍ<DɘۣX��gQ�JnRLibU�l؅��X�U`�6=#��oJ�~U�)�5��u�xNM���T�Vi<����wH�(�<��������5=��X�^�tg����1�l�1���sn�]-�o7��TSJ��h6/t���,�x��gh:8�b��R��NO͕w���vV^���1����&m��k͓E�+L���5��Rd	�����ҽO��R-�e�Qn��L�㸅���b�fJ�k+��X� ���[��iOmHR;�H��"I'���D�kkZ%͕b]������x�Ve\�v�W0�B1���ӛ�b�#m��eV�H�&�6�t$��������@���gV
_2�pSP�x@�D�0�԰�a�u)i8*�p�ԻF>���x��&^��@���OPɥ`���c�U�T&�;�
��mٙq��@{(ٵ4��Xw��f�70k^���TrL��8��-TwG�u�b�t�B�P{O�ޓMҰ�^�Mo�wf�Q��w�ד�j�4�Ol�gI��1JkwPұ��5	nA�.]9v+H�%�%fi.l�5�y,���\h*��y��'4�nf���(D,P��N�%T,�+���r�!�@Y�4�]��;�V���[��^�0[ɸ	j��Sg�m�m�,<B���Wc7J���R�v/+[�*V6�I���V�7��ܶ�˙����uk8^���%2� @��%�����Ku��F�mmcۂea5w��k���hm�Zw)�7Q�Jѻ[��`��+1�ӵ�<8���L������X�D�^#�v��@ʗ{FҠ�:(ǲ^�ʼ ���U�M�R����jS{�����7�Ke�A�l��#�7Kl#c�c�B,A.EwnX�gCb`W4������x�1���.��;��v�4G��ŲM��B�n��ٱMװ�[R�c4�(υʛV~��D��^拔]�6}(���AO ˻ת]j���f�N�d�QKZ`wR�]�Y�`�zv��+���ٳ�ER��Z����s%$h,���^�j��JȐ[�6�~�JՒ���:����ܭZ�K�v�_;�*vq�~��hM��J�%*:1K��f��CBQIQ�R5�����SFc���lO6���d��b�-��sel9���i%Q��	��(B���w-^�E�)
���u=z �V[�z���;��[�7*Z#So[Zcr(P�V����Co.�	 i���J]��R-���1Z��L�w �z��n�LfGkj2�VpU��R��6ؒeO��a��nӐ��U1E$g$��iw�l�0�����Ǐ2䥭��+\�2�t�,����h3;Kw��R�-�@���{�V�n�m�F4��eEB���-��cYB�b�t0'��*�4����;�������a(\ݿ���'m�=+91��&�����F��}B��
�	1ݕa�e�镐��N*�����	ղ]s"DW���<�^g-�q������7N�~�玧T��Ͼd�]��˰wn����z���}�xy�.trWxO3�����1?MP}��F;?	S���}�Qā������࿮g*F����;�}��v���b�,�D_��"�H�?�YD
��$���*2 � +" �EB�� 2 	 2 D���*���*!PEZ��D��H����"�"��(� �5 ����"	  �� ��"�"�QB@Q��DD�*�2�T" TD�"�H (H$�	 ��" � ��
Ȩ��!"��!"
�   $�� � ���"�EJ�!Q�
�" %E��"�P��!"�Ȫ$��+"�Ȋ2 �#"(�"�I
�QD�H # �� �"�?(���dPBU
�������_C�>W��o�k���&�PA@Z>$�J޿s���oÆ���>T�U�2(
��S�?���?6�~��1��tHį̫x�?���!�u
&Sd�Z׶����̚Y68Ymէ�5�y[���r�iQ^ǋ[��Z�m��\��*;�����T�ׯ�^�}ǵB�G��*�G����Q���jp�Òp�S��;ի3��>:�f��,����)N0�Xs6&�_�W���Җ�����-�n��A�uh�!l�{�^]ft����z��Z��\���z^�gfSEj�/F�q�gZX�m�E�U5�*�ni�f.]�X��҇V�9^��R1����|��V�w��6/��vF}u��u�|��%ϸ+̂��g3/C��a�܆.�ό��(��n}ٙ��UN���#4Z�L�F�p��k$���[B�nѺi�m����Fbr�z�!�e����̚7�v��k:�S$u�YoN���$�Վ��ɻ�_e��q��]Xr�;ݻ�V�VY���(M1����Y-N�WHm��d�w�H�7wN6���!��ɸn�9���G�Э�(c�3�ٷ�;"�
ϯv�M�+/o�#aI[-f�[���d�f�
Ct������)ڮ��N����:[U���tU�����Q��R[����n���B�*� r��u�ذ��#]BY�`�"B7c�؂�^t����e}����J�*'8Ӷ3A���̛�����ۖ�nۦ�:m�m�m�m�s0�p�]ؽ˷��գH���.�D	:�r*(�+ �[7Vr����m����u�2���v�w:�
���.�7,�fK0�iE�_[aLWy����.���XK: �u^?���w͝��%�TF�꺂E���1���A�W�M��\˘p�x���V��٫��k�fi��̱p$���Tt�wu���`��ٸ�]Ԣ�gMm�ݻ�QZ����+�u��uN����Mv�n�rf	-�V0ź�t�r��4��/�<����:��tU�s@Xg6�t]d7��!z�B���E�sMf�2��[I��6�r�ּ�{�aN+nTܑ�]M�^�O_H]��yp��RS�4���#�I�R,�����׋t�E\�hb������GA5��:q��r�afe����w�yn��k�8��]�P7h���!�oT=v���V��2�m�(Iܰ�FM�'F�n���"�e�zSs#�V����@i�;$��Kq6L�/�ӛ!�T/T��Gmq�	_&�������{����x�������k����Xnf�Q��V\�K%oM#�`u$��p]�-K��+��Vrv��>̬���[���T5��B�@G���� �p\�����}t��P�4�̧(v��sMc�+DڽNAx�S ����t)��r��:�E�m�X,��Zw�[m�m��m�n[m��m���m��M����WQn��[.�o�K|�YH�$�v�3��Q�x.G4�{+�K��l(+��㽑�mf�s�fw,BY���������NIĀl�%v�_s=3���#��=�]�S�{��d�m��4�� ��ו��ٙ���veA'zʜo.�x�̸ѻoC���9�LP���Lˌj��
�wl��}[��Z����fn��-��L�x��)ś5]L�r�i�ʽ�LZjֳ�K΅�^VS�7�a!x\�ۦ�gY���\��ӗ`+0�nA�����}QQ}�8�S����䬗�wW���L&y4=����U�#�@`g9p�w̅��SVb��D�<ބ�u�q.M�T���%Щ6�.�Y����Myٗ3��|h���;,����Z�5��˭�d/��Orr�I9�H�K!���O$_n@. $��\������뱳��ru��G�}��O7"��Yw �&u���,SMm�c�v�-Wj��y���6mȓaS
��
��7��:v�s%j�V���b�ڲ�ue�d����ӻn�ܒ�$�����M�/rꖞ�\ջ��Frl���J�e;p�rWn�~�R�vŅb�Y, �jٜ��0�����a��R�h�h���sn���ܽ�WsgvMwy(e�Rn2�L�)V8��m�e��m�m��a��o�ۙ��m�7SpТ_p�*f+�� t:�օ���
� ��͵L���"���Ω���K5K���-�ne�U�0���ܥ%ŜD��Z���4->(;�+c �+d�c
7b��l�7���-g
����b�t��v�w�"�Ŗl�˵��?���CM�Ei]���s�չ&tV���ڹYt�&C�g%<�T7�����ɍBK#\=�Z�.�T��p�D���Ƽ&e֌��[��]���W*n�-,O�#�x�k�yoZ7rŜ+�*���m���jн	�sSt�]ų�۝�4ԃ%NQS����/����j�"j�n�[�V�3kk56���fei�:Y�T�F�ݽv^<��I�w�e��bĨX/�Ո]��P���V�˗9���}�6�B�P&��մ�D�)��5�n�����<���9wU���\��:�a�'*du��Шnn.���au��\�-���'I�&Z2� ��9��!Ѐs����y��(������:����,���N�׳+&E��e�Y���;��ۭXGl�ɥYܠ�5S;vU�yx�r�:�a�&J7Mop���[��h�7�l�"s�0s��2�=����*����"�CPQ��v���F)=�f0���m��m��p�m�l��m��32�m��I���Uq�UG�Mܼ��a�yzx�m0gcOz�qb��+�wm�R
4əl���p��pa�վقa�W�N���T�{Trd�OU�=��{t��o�&Q�O[��i*ܨN�(J8Ra��hL���@�Um�M\�p��{O�40�+GRs4+���tv���q�c=:�J�b������Ȕ�C*M�9E���wiY�`�]������`e�V�;i����5��l=[,�Z����5�1)��+W�enGO<��e`���׺[E)�T�Blŷ;��5��f*�h{�^|�k�����$=}Ou�v�0ۗ�4�cW`�U�*6Ӿq�w�*��W&�UV�%���}A�m���Ғ�kUs�t�w�����m�6�_I��.ޘ��+v����'zBR��ӌe��I�WٱC����+;N�8{mX,X��o� V�K�.�nFҗJb�W��J��z�����ElU��WG�i��sg`�Dʓk�}w��^+9i���΂V�;�If2��λo�����n;�ݫɑT��R����i�Re�1@�+�Ó��la㕹qS�]WH��0�-��MFi�s�g��.V_Y[���s/
l����g���{hٮ�O;�[��́J�Fʺ��'\���O(���gk(	+�L�2�3!�ΙB}w���������/�;��˾E�D^�0M��ˇ(���ӸĻ��sh�:Fe�<`�_gfU��r�Ƚ�E���7���KM	�
�A;7��|�7�{{o;����u)�͎=w<wJf(MIU�l�#.����N����I��JWX/Jw��J@cΣx��A�kCEM�U�oj��PIZ�_st����
�G�b�*�.��/�±�Z�f��n�kaV��{*9*��&,��˚���a3W�D[{7xve�C)��p����8�n[����KOq���j��x]ۄ���®d�m�8&��r��Z�5tI�˙�nA�8L�B�hR[����!�J�b̩gF�	��Ț�7[��A"d�V,�+��g>��Y77c#6]h��^��s�;U�5�h��4i�oD��nӸ�!pإb�­Z�V�ԥ��TD���Wsi�^Ip2���<�
l�p%�f^�f��~��\�ְ�yٛ� WAԮE��x�ܺZ�鬌˝Eb�h;uy3t�-��J1��tp>l�X���,��'%*�#�I��)�y5[q*�bus貥�S��9O-�t>!ږ��3�Av�^��mY�N�d1��g-�%a�G��y��E�n���ͫs.��2�-�?��j��/uVs�v�}�U���Ԃ��W^��D�S������32M��˴q�X޹\�(�d��y0n.���zRi�v��3�4ܙ�R��n�[���[�N��o-Q�b���Q�a�A9/���D��:�t�µKcr
��.��'�{z��m��v�x�0m�S�����Ƴ�h��[X-�)K�Xz���S�R��o(^ހlڷ{������̮#)Y��3gV�j�Hŭ�j܌uI�Z�7g#$��an�iuj��I���P�����o�kkO4�J|�Y��>a�7;5���uˤ�w�h�\oV�1L�S'Ë⫶�K���h�RFp��ͨȫ���,5�w`;3+{q��=�5r�Li���R'���/�SJ������;8o��]��F5�zzXܑ��ya2d��하a��Wi�]�Uc]K�y\�.pW++	���!|���z�0B�fԋ�z7���Z56�5t�R�&��N��c�r�rś]��ƜVN��j0�0ė3�cj��r���a�yYZs[5���ֽx���,9;*��Z��	�!��l+:m)}&[߮^�}	�kFTY���3{��U��ɻ��Xwc.��Y]��Ķ�"���7v&�K��TW�ov�a����w�����X��
���(�d���\��3^�}r�b����m_7ҟ��j��Y�t4�S1��Y�N�l�V�=��L���X3��v�K�ۭ�!�Ȱ��{Y���Z�m�\@��9��X@��P��v �;�j5՛���9ݎЅj��]ڢ�`��6֒�1ttۂLS"w5�Й#&�����#���.���,��כӕ�yool�.�}%�ٗ��3�K�/y�JΣ��
K��л#��񶞇)*�
8ǈ����H )��@��J��+`�m��=��P٪B�'�75��yu+k9���k�Xy��1�6��:jv�j��@��'�R�b&݇JA�230Ҽ�@��^�10��6�lC��C��	�ږ���O+Z��P(#��q�S�xA��a���+.��X��-)n�����,�AGd̶�;ު�F�,	y��P��і{9R�3%�L�n+��D�Ѳ�c��Vu��o��B���c�����Ҙ�S!d��6��c*�;�u��S�k�:l���i5��e:�9V89��'o(��n�(����E�ڗ�%un͠ɛbU�ԢHzm6�;.'�Z���)ſe�]k\��>�j�������5hG�pn �a�d�w�p���HiA�h��d������k"�:�!S0�1����x��ؘw=���Qj[&�OD��0[|!W��y+0@UcS2��FU�ړR6�Λ��)ԭ�_d��u���;�и��M.�v�(���kr͜��kD13��'.��8�1�y"�	��a��K�6T��礇��+���)W[^^�ݮ3��uv9e&N���(_XYy�e��4M��u|+7)�WX�w�n��W>��vuv1��{v:A��h�/�ѭ�/��)��̸�=D��^I|�A��7�̉��8�IX3HW|�O����<�9
���3w%�oNjr���{zf�d*�����I[[N��˛��U�i��3���0v�[�{$;�a_-)倗Vq�		�F��yV��-gh:�,��:����T�Ծ�.m`;[ws��t3�|�ʱ\��h�C�^�#�;��:J��G�z��Z��pf	�MX)�5s�^�;��L��߇c����$3+�f�����n��A���zS�ұk���݊Q� �:s�j-��}���S]�}ײ�N^3��I9Ȏ���7�������ͻ jP�pյt�r)Ղ5�q��V�K���������2��W�Zo�>����y��:�<���Q*�I4���{8�r�nB����ޜ�m�p\��{]	��fүE�4QW��j'Kx���u�M��+�Gٝ�h(1�Io�����L��4E��ol��^h<lV�'�,<o,ӳ��UF3�R�<�0B-^����@�o[�9=U�&��,�Օ�'&gsn�=���\������&��=��dz0�!X���ˬ�[YhT�� z�IR\V�b�E*ގ�S�(�f�s�Wc
>��e�6T���&�k	��,D:V'+�jc��
�ȷ0�"����kq��^���jF�{{��\+D���=VM5OkFS�hi(�|�f�(���8�+b�h�A�]G��ٮ������_q�!��΍۽����3u{@V�Cp�K�+�7��gEN���W%�k�&��(�6�LnAԵ<��[d��U������&v9P�f��9l�H��Q��h��r�j8�=��o]b�fY�g��=�/�����y�Kx!���O��r�ޢf��]�{3'X*�9 ��C��(����)���Pd����Xrq9¶p��ɟb�X냡Ɠ���mN����`7xj.%�IӷPtͺւ�}/m� ;�d",3�wu���j�.�۩O�).����B�L�s&���*����.ݙ�2�.B�N��&U��j�-�a��e�;ZA`�0�9[��c��X7{Ʈ���~�DT,a $�j<Pr`I�$�*�A��|�ߵ�6<;t�laJ���x)i�i�;�3�N�9zI�۱����Tu���ѣ7;b�U��h7�����x����:����f[y��a���J��cla�q%̲�b�6n��A�31��+w1Ղ\l�5�����/ql�ʫD����!��a��h�l��f 04��v�卻�;4a��۩���Э��#��j�)i9���aG
µ.�cj�k+cI�y��`D���M�-�ћp�/neP��٭q���H�u�e���c�cm)U̡�pR $nlIL�S$�]�a���av�sR����ؔG:��L�f��\
�̸��k�+j\t�����Z�m�R�*�U��`�c�,��/LL[�y[\%��	-��"�ME Z�/:੫�q�#��r�1[5
l�ɷ6�V�b[G	����e��	6K�Ɩ�����b-h#�pTqMFh.��pk6�p�h�H��Y����"'Y�Y��``�8�����ذhn0D��ۛT��=����˅ђ�R)i4�6���kx�q��6�M���A0\E�ly\�������WX`��b:RX�#-Z
�����x���a���-��k �Rݦ$N�ڽMIb���8QH�)qnv�.`�J�Nvk�ga�(il� �jcpj2�q�M{&�l[	b�Uk�"[]�.c(XJ8����ƺ����5������p���105WI��f�-�%���kh�X�9+B�����ԪJm)H�J��0���aaq��L�v),�]�)F�1��-i,�K���ܖ&��Y���.�Xf6�6�jk5�[�I��m�x����õ�.ɵcsR���R�Mvc3�$+�\��f���kkr�J�(�9*K��1!K��ؗ�[tIu� �\��]a�t3q.n�
��\�q��BU�nn�f�^���-�[0U���8�-���,ZLJ�Q�rY��E�3����vWL�l�16qNƊE&&�3B����5Ɔmu�E�j��6;�(	�x�5.��
2�Q)�%1L��7F6�����a �<�d)(.�2�j�.&��,e\6�`�m˔��.]��v�(:�b��n5�(٫{h�@�@������]b��[�0��X�E�l��,1�!b����XWW�n�C��z�dH��˦RSF����r����ch8�duh���+�^K�\Pnν��8�k���rT������Z��
�f��kH�.[K
k3fQ�5�h׈�f�Q�����5QȸS�m�a�ˍӛj�����cB[�nP�;$�Re�0K�ak��^��-M���.4u��&�0��hM*�WU�Y��������bUq�c+�Q��ٴɴȗ)L�4�CM�i���%���	��.��c�c���cw�2�78f��Li�8���D��h06�*��g��)A�鉠.��x��Z��rI�3���ktV��2�3@%1c��R�4�
#�F�$s.�Vmr��4�VMm����y���I�,R�Y���Wcsu��*��Wg �c�XX���KR�B��%����vԹ��-�Mז�s�[^��\�a�v��V�4��\ˡJ��	a�+��ZTiayy��Kp�R�fT������nI�n��\걺3K���إ]���<he���P�F � �-�6$.��e�5�9�X�l0%���!k&p� �)�Q�*���6K2��:4��1�n�K&��[l���F�#LG�Y���&��(J�sf�ܔ�s����\u4b:�	(�7 ᅌ�Z	f)	q5 	M&�5�3Z"�e,5�nŤ`6Inh�,͡f�u�gV����d�yjZ��\��2���=�%v�j�5���� V�e�^]��fZR�f��4m%�,�2��e��2�vư�n���c.B:iGKfM1XP#t�i��k��6m�� n�B6�-am�r��طXF��Ω5�B�E���k$fjg�M�9,��&e�t��`Ұ���,�M(��jKl�F˶���4a�I�/\Ɋ&�Utx5�x�60,���ِ2,ЉI��ir�����cLD���RV3u�l�X�LT��[��9:�%@ ��`.�,�Wk�/JTK+M��s��4�R�P��^��m��XgK��W-����t�ӝ��:�P�s�e�	n4���G:63<j��M2�b����#V��	��B��eea���b��M-��P���(��bj:��[-�\V:�`ku�+�1�����heu�%1Jca�͔ݹ�ୂǯPMq��e�kb�)����%y�!rjT�۩v1���Y�W&S��ܶ&jZGfJęWhem,��j2�B�11
�͋)��8�l�JKU�[� �4^v3F�	K��)�R�͘Cu��M�e錛U+�����6M4�I�v��V�\m���J�š	���B&�H��n�J�f����у3FĹ6'$P��@f�"��8���-���&�gYy1,���bYi�,hɍV+[6���[tBSlT�ێ��1�9#�h��r�- ��B8Qmm9*��c�j1�P��B+����X�\8�ځ�XXt&�5uшc1l+���K3E�,�ץ�i��/ki�;�n+�LT�#��Ѳ�&m��W�Y�bL���].+�D�t�H�t�F�Mh0Lds]�����`k�Q�Mv#uAؕ�%.��9νT���m��%��.��vE[��-va���hܲ�6WF"��%5��у6мSW1m9�tc�]�q�a+JD����LHb�<�E%���t�JL�!t�Z��b�3P�4#��m������\��bj����5�\���E�L�Ԗ�Z]nc��[�CS�`���]vF�p�kdh�-Զ�$%��Ka��]�J�*�-�l@!p�/%���6�X)��1�JIX��i4ahM*X���+�l��\-\7E�3Ff��`�Hm���KJ�EƪW.c�f��ꍴb:���Z�n��v��H���ƅ���f�I.�U�4ɣ���Z4�]�94E,siz�*݆.&HJ���R:P�[í�L�-�c,:���#��͘\+)\òٴ��ȗnĦ��Ni6 ���!nM`�iۣ��c�֑X�(��2�j2�ek�̴e�ؚo\�qiQ���¶3=�+r(b�)(�Sv"U�a�vv�)5�iX��*�3P�^K[�v���*-��irs��
�3�[-]�6�\��r�Nv�wj�-ԙC�Ib�.�l{Jc���h:�k�,Ң%n-IX"�׍YjA��Z��v4��Vk�Y�nÓ ه�kqYe�"鮘m�L����7B�Y[{X��^��]�e-�iP��`%e.�@��L�m��v�k��f1�*i����a�H�Θ2:��a�)v�HS����h]��6��i ZGK��9l�:�g$���z�U&)���+(�SR�[��c0���1�ɫ$�n�a�Ps,�H�1�����\��]]��u�3q��V���0B�%����-���.����׬\
l[W#VXk2b[.t[5�%��6%���#-��KHKu�f�:��ˌ��NpZҎI�Tɬ�u&�� �ڬ&9����H�V՗e��ˬiuM���H]�08Cg1[-]36�Rǐ,���E��ȭ�欸�bb�-�e�:���6�tWh���T�lu�mlM�95,�s(��-;%����d��kkT8+eZji������f[U�Q�[1�n�L�C�nD@u��0X�N^��v�]R4�c�mEe���e���:�j�t
��\bb)-��MM���0K]��\�h��u]�I�ꉯmaEcia��51�\M4˧8�VS[
D�ST\B�4�{E�m�t�Z�] ��s��� ��\�k��b��9ZЭ��t�nLM�١��p4e��╬f���%�Q�ʪ�h�kM��GD�֖딷9��d]s �]�fh�9ai�&s)��V���C�t%�j)JZ��.j��n�M-ι�6�s���Du�-us�Ѽ�Mm�t#6U�Kh��V(9ئ�Ixʹ�i2���b��f�EE����L@�i4�.���nt͙�Tf���b����!�˂�3K1�̵5ƺ*GA�2�6(Aa�m!�-�L%�a�X�6,Ќ	������cm���K.i�c�\�geݖ�S�ڒ�ț[��F���g�*����mz��ll9�����ȬZ]
�a�2ka��w+lK�Y�kR�Lec3A��
�f�쐊i�r�	p�s�v�7Y��Յ+�69�����ja�45�J�a:�L��.�n��i7ʸ��B�)���	eA5a3kAhf�mLb�y�f��6�of�r;$mҺ�0�-QUU�1��ek�[�vV�UUU��k.Y��ѫ��Tn��
��,%�e�ȇ[�tp�a��� )i���p֘T�ғXXk�,P�Rc$`�%�uEgH�6�����Xvq�����e�T6��glLb�9j�ub8��:���,n�r�]P3�ʹ��Y*WZJd�ײU"��� �˴��
��\�2�[_�}I߿d�$1����j�T��FC+�Q��ȑ��c��1 D".8��˼�{��&(��*B�A\G
���$X�E��G�1V0�,�\H�e�;��=�AE�!�)�(�EN�V$DT�O&F�qȕ���|���E22HH�5.ؑ
	,,���jDH$U"�%�DpM��;s��$S�qrHB"�;-Z�d��6�f��W#	Eb�d�B1�I�*�"癈���g��y
��eJ�*�K[0^�cI�a�[Rmywa(�]0an�(U$*[E�+��l�RpqmF9����t�����6.Q�c!ȭYJ�%��rŲ�&��<��F������/�),� UZ[,]����Є3-�km�K��!C�j��B@Y6Y4��"XAl"�H�:�Y8�"���W&HA�8�,j�es
�� �O�xs�?����5*�@v���V���w����M2"M��R��1�G\P�:�t�^�2��%)f�Hd�3p�V]W�3�6�E���0n��Tt��鮘�æ����var�d�"*兽��иH��[H��20D,�e6c[v�lc.��f������uƘ��!fiT�."0�ebGLfc f ��#��$+eԗqo-%el�٬�V�D&e�%�3h���o�*�V��l�34�F֎���ҥ��ms�e&�4��n�[���1�BU�36�j�gq���R��S�y���`��;i`M�]�j���Cyu+�c�J�շ��:mj�*��3)���J6Z�"��n�|<<�.z�I����g
���aֺ���a��&��6��m��1��A��í��J��Ҁd洤�K�Ś�>3�.��5�)��AK�Mj�QIr��^�m�n��WV�b[��3�Kly�oa䅳mF���Bh2��ƴ�l\q�m�jQĨ)��K�P�0T`�ZRln�R$�&�DV��#W]�A���Ů�������r��j)�g6�0�!p��-�M{%5�6mz�[�`m����4b)D�����rn��j�/4���-����୮[�G�6m�&1i�� K\֙!��$����j�W��9�̌�g�f��c�ɖ;� l�a,�m�ꅉb�]v4�f(iVݘ@%.�n�V����۩L��8��+�t�R\ ��`[��n����������[IW%�:�[X\�40�J�Wa�غ����*n\�5�ʱ���f0�JbW�j�ʤ.�	E:�̚��۝M�apřæ�R�]�ss[i���Ur�*�����k�*Yk��2�cRcLe��f� ]Zֶ�s��I&4�����)�,�YK[z�P�:�h�̣a�C�^��Q�-����cFV	P(V5�+X�Q�Т��-�lB֑m�T�
F Ť+b'B����D�^��,J�dƖ��ՄA��D��icP�*�HJ2�k��XAc�V�`�b�YK$h�(��^^
��P��U
������Ͽ�4?�����)���]�ΐ�۰�:��$�Cت�;�~~ڶ�a3���I��m�[pS�ՔB��5�Λ'�}b�F-Y���T"���[~�� =��:$�we@{v��ٽ���O��f��Z���
�D�~�J h�&k�L�$���Oym�=���I>�v܄$�'��tI���Y@�p��G����{�;|I�%� �$M�I�>�Ia��;*Og��e!��.Bh>�YDZ-R���,t� �>��!�[Ow��U��뒉?hOk��$�&��{$�+���6{w���>\�I�e�!4F�m�f�[a��p
���5	��"�V�V��{�_=�56�a�6re�!5�ʛ ����	O���-n�x�OL�RŒh{9�d�4A9)�J(󻭸������;�Of\���u��֌3u�@F�Z�����M�2;�B�`ͨ��Y�%�s]q찱-�y`�KW��p�j�5Cs�&H�y9U4O�0�Z��iʄ�z$YAQ�(IF�<���4M3�؟h���p��$=��?�4I����P���4=�RV�V�
�OK�zK��v.�G�k��:d�I5��I4w���0��!5����I��t�&���HQ"�8nwF �N����}yӣ{���"���30!��w �D����	�=��n��Zݚ�-(��5e6��r�R�..�h^�P�M�6i����2��#�(���]{(#B �{�~� �W{���N���c��t-�I�;���R}���*�T�C	��������'��W���2L��&��d��I��u�A$w,��1��-�Gݹw:��(�'-*��i\�{ْ}��[�I'��'X�5v���U��*���|���5ܔ?u�?+�����n���<�|p������bu��s��^�4� |nU�3A��;�Zq���@���$�����.?�Z�`���(Hkg��D�N��e෼dϦ���""A����%j��Y~��v)�Z{%Bk��{���"�
����=��$���Hz�ב����uD�I�O��/㗯��$A��H���U��^�F�,=x;f63Y�[�E�2�a�Ю%����`�J�R�6�`��$&�/5�˺$=�)@ #3Γ�gl�7�M��=�H@���T$/
޲��*�RF)F���d�5+l��{��1��	�$�kם됓D�����	˻;�nk��p籱>2}�h!tE��RffvEĒksʛ$��U�Ϭ �⽘��ğ�^o�UBFg�'D��F	:�Q7����G��8�W"�10jѹ>�Mg��+�A����`��z{)�h�k:L�U�X43L��;Y��sU�#��:\}��g�U�{Vu��ub�x&��n4��~��ǃIE�f��D3�MQ�Wsb�<�`gEL"�$A�:��x2h���w��C]W}��o�q$�Zܹ	4#3]&h�O�;�$>�JC�1߬�6���]�*v�43U�J�:84�Ե�,3���B3$H��JWY#F�A$�)D�"6/�P�I��T� <�l��z����&|ֺ�3�9s%�fY��T�Q&��� A6P1ʣ~ΌBp�������(�>P�$����$�9��!���ry#8Y�6��6��	�:��e(�ڤ�R�_c�ɪ$�Og�ʄMf��n�z0}.�Mvj��D��k��y>k�!tE��
��1ٖ�+ih�}���@W�W�$�sݭω4H����&W��ҽ}](��	5�U'N�כN+TM�e%rQ��IU	$��}�E@�����'� �k�?N߽�!Û-�ת���7W�4�ȧn 1eF�J.�h�\z�q��G&�eD��PfnS4]�HM���}��ܖ*��K2�_S���FR��^�%��Afع,Yl�rG`�S��6�D�A�[KM4�G�PVbǶ4�]bKWE	��i�(U�R�c�^1IV�P�lf����1�5�,�Zܚ!4��q�kE�洦�:�թvr���XU��7WY�+�2��5��	s�X]LS[��6uq���K��h�p֙��j2���c�K��S\8&�v��%��i�QE(kj���l,�\�ѹ��̚�]�:������L�_�P��Q�D�g�[� ���u�N��&5��eݒN�쐖��]Z�I(R�"�D8��W�X��d�k�f�[N߽�>����l۷è��
 4�R@�Q@�>7��*D�t�(�xb�~�V�/s)a$��풪I'o��Ġ��O��(�ڤ��>5}��\��'��$�zؔH���rfyR��fs���?T&?�z�EY
�(@%t�Q'�&�<��X�~�o�Ĝ��BI=�Ɂ	#3Γ&{�+b;�B����H��0�	b�3Π�D������H����r���ψ_��7�����l�Rzȿ���N@#3Γ'١+�.��Y���%B	&���R�?d�ϲ������G�Hi;�~'E���C��[�-�=�PW�����O,���h�8Y�Ӣ� �p^^ʙ�Y&U��;�f-��"r�^x��^��l��w��HI$��Γ$�)}k�4��K�qj�4H#)B� �$�[ud�+sU:d�]�Vg�ʮ����/<����I$��ڤ �Fg�Z!�p��v��(�c�/l�5gޕ�`{�C]%8~$�Gf�N�$�>�l�B��髁�I���ү>*�Wi=^�O�OĚ&v�C��x�«l�I��R��Gkt� ����>��X�V\�Lx}�D6�^�7 ���eH鳈���X�.f�<�ku�8̅) ���f�( �8D�˫��+�ʛ'�@=��%Q+��vU�|��A�wt'k��|�#��D����yǰ��r�{��w�Ǵ�@4'k��$��nP P�,Kڗ�����O�]����k�᧾t�D�3�� 'q����<w[&�y�V<�o��2a<�SMWx���0ak���J�t>z��h�uwOF�gs��,���S��;�:�10p��kI�/5I%�]o�d�P%�-yJQ1$d��j�jL����Ě&��S��� �d��$�'{ڙ�sjF�a�C7Γ��A��ڱD����ђD�Fo�|�l���;�ͽ�[<�2MN{vHl�Y?��S�F��|w�{�=>�&�]q�+����a6�F��V����2��(�UՋ�~�wχ�Y�l�}�5y��&�$�n�%h�G��Rٜ%�㧓�:�:h-�s{n3أs|낁0D�A���˫%n[��gVz�ʐ�@?f��>$�>�j��J����*;�@�]�p\$�B��Js#:d���$�{�p�$���͇��:�Y��	����~�$�C��{�>��L/)��p��A�u�G:��$c3f�!$����RI#ێ��܍5dz`�/{JO5V0��vg;�����r���S����ޕ9�M"�>]Zk��`�����4jn��hTO �ۻ�2	��
��)�4=��N$�Mf��~B�#���'r�ڢO˽�'ĀI��R~�3�ATF�h��q:7��ȉPP�@���|O+5�3��F��Zd��Nfy��6f�_�^�8���`�W�1g���&���L %n:L���=�v�=<1��9i��wGB̫'�}�j�	��q*���H!5�2I�����G�·Q��ꄒh����T�H{q�tH[�}�{�Ћ�ޟBiϱu#B��*P�$5�>pD�x�z�@�$F-��ق�z�:�DDA=��!�&���:$��GCBT�_Y��J>��l�l���þ$������ �5G��<�ٺ�X/#  �ܘ���J��Y��O���6M�k��Kin,�	�����$gk��$��r(z��ayA(���-�X�zߏ�b�E�j�y��:��o	3x�1�{/Z�8[ˡ��vU�r̬�l��P�VT�o&`�����2�"s�p`k��%4/�$4�J���vΖ�:���L4����gQ�Wb�V�6RXd6 [v����.����"Z0��l�湲����T�t9�-��V�R^���B1��W)�^����\D[�3��e�֗-�.�:��G-������9�fP%fK�7L�G]�,֑1T�nS�ٗ5e�����J�[rf+K���q�����	�b;MA�CE���V�@�v@\��L�޾K���v�݊��ӽ�8�kwU �$�g�@մ8
����%=�*~$���HXV 4��Հ
A߼��D�Ԯ��ϣ���uf�ܩ:$�O�vHA����i����Bh/��Ī�B� �S�W9���	>������ه���k��#w] $��������W Ϧ
+�J��B
B��4w�A�k}:�M~$����>�OĚ�}�ԯOe��B�a��׌/�4�� �WGCA�����{�#��G��Υ�{ʮ5���$���d�h���@��jc�����*�M�A]�t\�3�d���#�1rD�U�:��d.�������=�W��m|;�k}��̀I���ЀI4{}�B`�O��\����HI;��T%.:7ƕ�WdP�	��NQ&� ���=5�*un�{�}W�7�t��U��76b�����8m񫬳 =�z�o��ro�.|C�hz^[��m�+U�{���h���$��D�s��>����'fq�2�&I�p��V ( b�b4I$n�g� h�������l�|qK�ZI$љ�	�$���1W�z��WH]�k���u���)� �x�.ݔI>�E%�fyҠ����n|H���	�}�i�*�T�C	���	 V�!�����w�Iܛ$�Oğ����4I�fy�d�qү��z�ޏ+�Y�2.f&ˑu������B �����!R	Z!"���@��D/��#l��Q'�G��$�$�3<� ib�u������$�>��>��d�r�+�H6�+��u2I�^{ˇ�9,�!4I$���!4h�3<�:$�M��al���BR�!Ѿ4��X?
���Ύ I��T�^�J��C��'s�O�*_+=�t֋�f��o��9�牀"�-<N�=:��/�W���S������W/Q->��Ц�յ�R�ڷDe��w,��N�.�{t4�C�`"�s&�bS}F:c6�)��ͭ��t���.c��#@�Y���I�Y��� j=� r�P�;�:��M��ɽlѲ������,wk]J�ޖyu⡒�#;�M�Ja�כLPV����r�3�Fm74Y�/���=pPo5��z�k:��v�D��9�V-��4Gr�xq�P=�����s�v`�0���7'R��'L���я"[Rճ0ԍ��]�"�Ep�iJ�Zim�.]�E��uK5�tDLUۛ���=��˚�㪳Ы&�'.�R�f��%N��+y]�������U���QCn�F��x�
Un�-���{Mtɫ4!:�y�ɷ���F彻Z0�X&�蜝�|pQ�n
�x:X+��vg uu��,���K��1.T��/�Pդ���7���o����� � �����e>����k�݃�fܬ��%0^<��bj#^�7��S��B[s���k,�*b�d�v(J�L#\s�!SHN#^	u���� ���:���ٶv��gL����=�]u�v�u�![��uh�󗝪�n��f9*q�@�T8������p�w�P��m�N�S���U��n��P�Jw&��Q������ �_�m��ve�ME����Ў$�6b�k"!�25�Y�Ē��kb��6Ns�^v9\����d��l������C:b@�7�X4�c�\s$���J�5+����y�89��ʂI�+I	k�Tc�"�5�lb�)Ȉ�ͤ�Î��$�l�y��S��|J�%r�� ql���v�;�xР�J��qqF��f�8�q�J�Jsh��s<s^ζ[ ��X�p���*�´r�L��i%b��rW�P���9�$.�'y�""f��L@�!��#1�q�&(��1���viDָ-ci*�G)�rsvrLq�jD�Ҙ)�6R���(B�Y!e�M��#��.�#2I			����((D֣���&Y\�YX�T#��XD��jj,��La0l1`S�u:�6�U,�]a�6�9�)!*6a��R�TRB��G����V])\���T���+�)�d�j)���[q��Jc�RLL�a��&r�d��d�"�H׉P��*q�\��k�U��TGf�Y(v���š��p���$��L���V�����*�D��w��$�E�jy׸k��}�I3�r�K�APs$�}�;�e|lFGѤ�r��=��^��HFe"�]d��A��$�?���C�'������N�&�o�HI$��� �{veaF��W�/�C�l�|�5�蔺l�l�(U��K3�SW0�L-E�[�ʥϯ�z��51k������$�NT�$�k��$�ѷ{���}������vn���<�2n�\�A�����#cIv��W)��&۸3=A\G�3�����&�7�^g?�p�Y��nU��D�k�Tk��A��k�	��_�S��_X�x�dY�4I����$�I=��*Ip!ѱ�]Z�~ ����e �j����]Փ�'��wqOwڰ�ßC����bN��Q��p��&!���
 �*a�a��_q���]a�W��nΐ�WN�.`�c+��m��/��$bg��M�Γ$�� ޠ
�-S��J��O��o~��T�++p�$��U�Oď٩� �I'w�HW��(C�}�e��00�P��CD�m�v+�Q�rS)��M��\S.��*����e%��{(UDG�"a��ʄ�H���RQ'77E8��Lln��$�I��n�	�j�F��
�P����p")GY}<��_2$Ҟ�v못5����I$��~���J똿.���R���ۦ�)B��������}	�$�#��l��F�'Yh~��}�7N���)mI'��I���'�}�ܧ����/� ��8k��S��q.��&r�ͯ��r�$�_����I��Ε�՝�Ij�Wf�ٱ���C�c�]Z�~!?���p�+f�t��m�tO���$�D9׳`_�7>A�o}����&����q��?a��*=�.��gw��v���ssh7�0-S5U-�U[m�R����]����gV3[�o2+���O�9���f��`D����.��0�R���ƭ��wYc�5�AZC`Ԁmh�F��4��� �jB�s�vŚ#��2�ZmUنA� �fDa�E�1+ջKVݢ朷Y�h�8k��4if����:�"�v�WK�y�l�R�]��� s��M�e���Pt+倦��v�)�Pfj,�ڢ�t��2�:X͚�J�[Vl�a���sA��Q����W�]��iM�Uб���$6t�1�ϯ����$�(Ư�-k�����׷�f�?FO:L�k׹������oa �>ٻ�2�i{�A(��#H�v�I?���U���
��Bk�wD����r?:O�'���c�#��
�r*Z���aj�0�W�'n��\���h��{��W,�qN���d�$��O�0�D���I�M�~�A�������&C9d?��g��	O& ��_ɒ��=��VڱF�|���?ڥT&���R�M���k��T�$�3��1�۾5 e/b���5R�>�%�����%C^g~�=������g�Q���y�Ȁ�j����������3$ar�����ߒ�ml�/
�3s��H�����w�vHH���"c9�uʄ j��L�AJ'��Ub�@����$&]�璽nF}����M%$��c�D���t��"br�[��Eීs���8�ܖ4�c���W�`�i-��}=�w�R��$��t�$�����0!'�7� �q�\�x��%2�T�IB7�t��B���L}�j���e[�Sg2,��ӫfw�q wj��$�O��tc*T����h�j� ���}R��gx��z7ʝS$��&n��$��uw�d�d,�J ��AW�g%b�0���Ḥ�ْB~$�����ڞF����Wo��tw��N�$���ݲBƉ9~����y�＝�}J�P|Ec�Fl��h0��]1+ap�[�x�%⼹��>�w��yH�m|'�v�H ə��&�4bOv����*��50�2���Јr&I����J����ȣV��M'�~�򄒠��ٝ����9V�h�D����e����r~%������j���{XH�UX����/l��_뺳���|��M��ά��5b��1.̣r���jGm�"�Sk�Gb[�f�`\�{*�3�¥��w��NeV���IL�(�߹��3sK˷�_Ǉ���7���A��*������o��T^���j�A$��������?k���I&�O6'�h��^�ܔI'��_��U�,�>�!cn�&���MJ���WvP&�W�;�\z"G�(�c�k3�Ӛ�<�I�o��d$�#����T4|I��ݡ$�tf[]����*%"����Bh���S�+�k�K��v���feu#2�;g����~e+�6��6G�I'�|w�쿬�M~=�I/�φo�v��u݋���}�`\@J�2*�"I���Ú�D�H�A��-��ߦ�:������?W���x{�v����l�n��WZ�5j��S�O����� �:;�4I$��r,�������N_�ە5D���un�뻖��G�*�ZF�YF/ޚ�H�6�b��IG�e�d�G�&�DD�����֏�2ԗ����S5eM���@i��5��T���.�|���oq��ʬ�3D��[�'mT��sn�� �����?F��`\A���j�A$�J0.t�4h�'�n9�B�=B��_ku��Z��r|I$�;�����?da�)Tcq�`�PV
T��*�h��M�a]�����&�c���Z\��g��}��Q��(j��grE�ug�ܩ��,�2du}�v"(wW�O���^͋��g!�	&�4*��2�O�%(ϴ	��r� Z�|�Z9��BI$��V��dc�ʫ5��~j�]�b��B~J�yB�$��I��::h�I����&���]�g���-~S�Y=ʮh�G�~�*B7C�|F�X?
�D��jn���v1��$�O�;JD�D�O߽�|I�I����PyZ[��$��ղH��<�a$(�ǔq��rX��?�"��nd� �q�+�Ò�d�?���ےh�v��nT!t�Sޏ9_z���#B�D�X��s4����
��q/s������gi�]L��"�܆�H5�F�ً��������Ϳ�QI��ԋ�Ѷ�o<GY�B���y�Xime"��q1�`̻��Z.���Wp8�+����s)P�FU\5���bh�f���*�譼G0k��aE15��X؂��Gk.�J�Fẘ��9��l�Xe̸U�
�sw
M+�� ͪ�5V˶rP��k�X�F�te��T���ɫ��A�n�[0e��٭����є:�`2�	���$�@l�q���@�in]��g��~O�8V�/�:D�D�����U��~��!"��u���]��/[�$�3���Vw���1���@�Q��%&ţ��~Ua�I��;r@%N_{n}?7�k=�$��w�v"
GNġ�J,��$�<v�P���I�W��u]ʻ�]����@���܄�_.�Q�I6�ã��)�z,fƳzM�L�I&�����D�_���oU�K�n���srIP����?��A�`�+p���tPN�N�`���7��Zp��.ɭY$�I�����mϧ�ʵVO��ճ8����{�~��S�[,�ie����\S��^%u6�GlС���l������������K�����O�����P�I��}ҭ�;�(�Mg~};K������ە,��V�6�w�R�$���?��{��ۛ��A�'�b��p�\y=�����xx�1v%_E�$��Zf�Y��Z��0M�ׇ8�F��)c#��ϴ���9��MQ&�5���rQ$��{�\$�1��V_*�."lYu:"L̡(FG�2��J�wVj��?n�4��q��A0!�����D�3�]%"dFO	@���G���n�:'�=�{��w����BI�O�t@Q&�g��Ӄ���h��u��7L�r�D�k��Ū�Y?h���ϡv���5��ے���'}z�Oğ�_��ِ����j�ۖ����	�,�1����5�S B��̠b��LW�L%XѢ~(��Ǡoz!��v�������N��&�j���!ۭ�`9�Ybٗ�{�� �'���΋$��~|����
�sch��ŕ�-!�~U��v�4I�޺,���?�����I"��+��s��Eqd�D�I%'��CD�|I����*G�ݞ���ju�z���Uب=<��.Q+��;>dާ���x��-�^y�� �v�5�]%�0���k3��a�mْ��������̉����t@��g���c�	�Pb�Q�wj��F���^)�4E}y��$�3�JVh���ID�$��~��`[��|��3�LW������A���B���9�����h���o�>݃GgE�'�_:.�5��`�I������swB�ﾾY'�}zJ��4�p�VSs5����[���ش*�"\\[��R�w2"48��D��a�'�"�'7<ؔI�N_�m��2�7ʵKa�un�?~9��į&��I
�V}'����G�ѺϜ�Ť9DDDD>͒I{�l	���~��گ���yD֭���A/��Z��BI$��m�� I�7Äv+BC��D�u��8A���rAp�<j�]��J5s�dz����/�M�w\����m��&�#}����ȍ
;�F\_=�D�q3%!B�:n{ɿV��Y6��3G�R���{��w�j��pZ�1T�5`��}b�Z�
I��y!����$	 ���"/uܨM}r�]~�uv�&�8M��"��M���u4<&Q%�Ή>RI�$�����	#~�Dr
pE}��J���d��y�tή�A�R�
@�%֨���b��7lﾡ�_�Qwi�w�# J'�ݱBI$�3���Y���=o���m�g�#����ֽ�ħj�=���	6�Q��t�	2#�mw$�P��k�.#�g����I����d�sp���(�B'����.��!"%	�@��GGc�dǢ>-���$�K}��	��ws����M_v�hg��d��8��A/� ����ՙ3�?�oĒ�Eh�;��N�$��?l��\As���]��&���'�xxxՔ�I$'�j�m2h�O�v���wMo�K�y�y-��2��M��lʈC'�ݘ�x�=�@��,�!��C����8{�g3X�nK����LffY���knlw�,��v�n{3*+F�tf�uU�4s:%܆$���z볱�J�놯V�ۇ�{�>����{1i�þǲ��V�ǒ�Da<��&:�Ҳ^�ǂ�1��LL��,A���3",K�+��{*޷��4g�ŕ#pɥ�^DA�7��S��#e&�xnksu�����[�J�7)*͜pܕz�D�r�|%:U���l�����1���;�LLY�Y�U���*�i��IPh5ك.���ѴF��a�2������k\��#U$�,�cLܡ�W�7DH&a���T*�wJw�6�mv����^i�ܲ�_f�8�v�b+>̍P���%��;�X�퇸)�΃�E�z�`=X�-�dҭ�s�˖�J')���t�f�vwL�nE�����R��9`������B�9���پ.�횵k���kr[*�*sJohэH��]�M�"$�D�uy3�l���Fjj��Kg��ts�u�;�YJ�v�y�l�p�]_�	�y�:�5�#�<��\GvA��	u7nZ��{C�h&�ac�N;��/���)�64�q+������)��x�&ޞ�y\������m=G71��D\���[�>�݄�wu�R.�`LV	#,��
2���/��@fMf\��$"����C��L:J�"��!I-�`[@kN�nб�,b_�kz�l����t��7hi��f�V��L��h�{�|���W��q��5�28_��}�gw��y���}�e�r�����K��j!6�,��HA�^� ��-�PzP�k�J)3]�VHC5�T�.Vo�xq�,EW�W�j8��қ)\�AX�R�H��1�
�%�ԍu*��[l�Ud4C(�*�T�$���7X�H!�ȱ�HԶ
�D�XL�`�8V ��,=�l�����2���#�u�&y��]*D�+������a��#�X��l��n7e���@R��&,r�������2C<픎�� �L Imm�h�pw'P-�u��e�a�,�ݚNZB6QqAqE���\��4p+a6%dʕ�PPQQ@�fA�AE�Q���� ��" �b�Kٔ��Z#��*d��͐Dl	�Y��DD]ClvaE�!fBL���TW
Ƹ#u�W""�"�H�Kf5��F �0�.k��\�rɒ�Z��R���R#�5�Wl\�$-�7\Y+Ps�-I��L	dB���X'R6��������n������CH{X�U�f�k,�3���L�D�@�`���!��L@S��Q���A78���5�t�,FZBYMnCJ7ZJ��]kAu�֐�H��4�A�e�@X��n��� X�LE��`�3V�J��K�ZX[e-��`2�̀�[4i�s�e-��h⑂scYv-���M��a3������t"��]uH����MveX����ы��hXa�X)+Ʌ�ڰs�&��-��ԕ4sa��nΩ�c�X$ɍ�����#��4��=V��=Ko0l�6��.�tm�x�kak+3&n΅����V�*��U�fMe�e�Ah�V��hcj�R��Y��.$J6�����(��F�݆���k�h��A����m����J��ݓ8XE�B�����՘��,J�ʢ�AJ	��ƍ����\� �����8fV��嶂�U�2�P�]��*Jj�-�eZ��s\���9ԅ+��u�6�j��#4�F�Z�r������Au(�V*l���V�6�"��LXI��b֜M��\vW�uL��ܶ�����ʵfj:Q8آ3mM���3�N�(�D��Ĵئ%(v��U�ѽb�h���QYcũM63�u �x���e]-�P@���-tѺ4U�t��f�Pa�땩rB��cĩװ�ͅ�,e����ԅ�CWl5m��sM��X ���-����t@�4��+��6j��2\�YaV��hR6	[3��z�@n
s{8�m���MG�Pv�-΂�uut��ȷ <j�&�!��U�Kp�֩���[@#�L�9&.��N�s+K���톥��R#���\R*�V!v�t���+:���R�m�l�0�`Gk�V�+��Ff��3ř�J��6i�7[5��+VmH�����Ð��A�Vͣ�ls���ʹu\���.�R�����E��0Ԭ����Պ�I���y��N�'��!���[G�n ٝl	� �([lHE���ƍ8vpk���D��-u������L6��#qsa��p���z�tpP�![1�]�a��;�YJ[��Vݗn�q� K����u-�e���[q��Ź`�VX�R-�CK\�]��.3�b����&��J��	�2��f��4r�%��&�B3#��+c��ː�����J �Tmڎ��c���Rj��v�G!0�.k����￿���]�]/�i�^>=B�G�����wv">鱣���=��G�2��o�${�:L�T�[w�)X"��3�Od��U`�v��u������p��f$��
���������L¸���̟��9(�3HT�R�8xx�N�4HۮBI���^�����|_:
�DD@�ݷb��_DK!"%	�@��)���fp��v m��uv~$���Q&��G�/�ku���~���?P��@1�~QAK�U��T&�뺳��U��{�޺L�I;�vHA�I��a�׼I��Õ�BRVm~���ª!��2�VKf�%�%͂Z3�l-��Be	
e�:z�AL��?e}�>��$�Oݿ��I ���	�����|��lZ�I��'�뺾����L��������BKW�K����s���P�3�P��E�c�.�>�i���l�c�ugs
@=�|d��7X�P8�9����[��}8f��]W�C��H���@�`�ڂ?DD@��쪸��t��k�����N_z�+AG��ԽD�tm�QJ�v���G�B��z�%�H���I�xz�k71u =D�3�%O�@�>��L�ԴI��
��J_	~�
'v�\Qۺ���*	'u{�F��n*��o�����ч1�|^��T%6�7�I
HY���7�LD3q
��y���&Z�X��O���tw��2��d���\Ȭ٬{�o����.��գ�; �l꫐��)��uwhj02�4�h� 9cEَ6|�����5�{z~W���N��O��*�+��������Ǯ?y�8�}��d'�z���$�I�;�Y'���m�exOڱ��4H5v	$���HM��whkط�o�f��ܮ�F�$ݪ�U���D�k��(TDD��칏�JPd�.T��-�mQ��})�{ݢ˹���+��	nVy�}b�n�j�O.���EnOkd�~��>�#ĀO�}_�l�Q&���_�/�d �F�k��5m�r��E+$]�G0����F��v�<$����i���V$���v����n�~��������)�iX��t����z=��"h�3؛=W�q��}���{�r~'���J�I$�߻c4*�s����?v}x��e���Bܚ�iZ�c2\��ˁ�mKh`��9
�*��=���d�׬��%8w=4I�'Fꦥݓ��w���z�0���.r��]�!�����I'�|B(�_[P�>�D����yL�O�Wd�^?�տ�4I��ݲB ���\[��;}�~��W\I�()R�6�heR'�M��rD�?�vm�xR����c��x�ul�I>���FO �ՒU��6_�ʱ�@���?I�����Y#�~�OI?O_�e��J=����Df�I�w�3W��Q�1�V�N�qi���jTzlZ��vl�Yگ���!�J��8T�YЅ#��t9vp��	�d[�|��|��c5T-�o��"��.Q���H]]�'���)EޠwHV+�J�\I�r:�H�.����	}��2^�r��Я: ����p\9��2��ˍ
ԅЙP1�m��Jۊ��V�l�Mq�A*�R�?Ƴ���2I$�\�I'�N_�e�K�x}��W،n��&�?�7�2[~�/��!g�X?�[�q잗Ba��V/�E�&��t���߲��Y`�.�g���m�Y7j�I4�{@�x�Q���Y�?E%BI$��e�� y]�9�u7ҭ�O�'{��}�.}	�Y�`J
T��#�	};4O���#�� �v�Y��t��WC�c�O���;$��s�MJ#?mF�$ݪ�J�o	4O��T�>�+�pn�5=���,��'������F��I�y���_*c��Owz���̳��g=�6l�F=�L]8��'�c]�6-�;F.[|_B!�%u�~^�����J��M�]c@�K�ƴ\�1�����QF@Y$DC�[=|� ٪�7]&[2��D0hWM�iR��e���M4i�3��cA-
�X"�]��)��ⱶ(7���  ���6Yu��D3Ֆ�%q/i]v\�1�/1��wP-z��rA��;H�;=s��+�f\hG0,���m��5٣�,s"�����T#�Zff]�s5n�ʊ��Yq��Z�!����X�X�EacU+���0.�]]�1F,Ji�r�jf�ar�߿�����P��|�;2HE���s�h�룿�Ru�>߳8���a��f�P��ݷ>�O��&�%�L�^6F� ��Du�Yu;�>�������?����Mo�T�$���&��;���"����?Z~4��>η^�"V�B���xcl�>5W�興����r�h��j��$�<�� ��Q��������fW;]�&���e)�*H�j�~�I�$�G��e=�Ŏ��~�4H�]��q
+�`J
T��,ۡ^d�h�{u���^�x���z�\�rQ��$n��$���d�sU*b�*X���;M��M�X�&&]��G@�4�cA�X�[t��v�Tޢ���*�}�6rI�O�j��]���������~�����B Ѻ���m�7G�	v����ّ�TO�;�Z����+5��h�q]C��K��b�¤Xt'����N�o��l����i{ih�y�b���`��=��]W��M_	���H�H"� ޺q�d��!��9\�DG���w`Y�ug�����˲#_��&��M	zػ)|$>XuD�3��	��N�S��+3yfN�\�I'����h����?]�����hY�Ԅ��ޟ��)zm�$�>�M@�{7d 	G/���FԐ i�:�D�u��;I#I}x�����Q<{��_�Vp��m�(�-��I$�g~�>�ha���,��{�{���]r��s)�J�j��ZMl���{���ʆ r���k{4�7dZ�j�B C���?��]߽�Ͼ�D����n�K�{�9%��n�D���$2���(�H��PfQ6}$_������f�A{�=U� >��K
fDDFOv⳱����ѽ=��d�.U���փt8"�"��3>��̒���g�N�@ZE�b�|�+c�Z�Ur�gl� �-k���K�F��Η�K��Y���7ܵ�9X�.i,�-�t�솷�c~O��� !"�"y{ޫ��Mw�������nUB�$йeL��KƮ4��Ѵ��5#p��2v������{�Bj����a���k��Fb��܊� d��	�Z#�m|օ��HO�����$�ʝ"��7��,��$���J$Go��� �j��][�fﺺF�.��ʺ�pAY"� Q.�~��m|8�M�vuP�2%�pd�sn6���؝O�d�s�����~�D�>$�t��V�&�����ǰ�TI;{�"/<x�eR*�CQ��zTDTϺZ�����$�'�vۄ�7����|Hf�p��,����[�\7%)DB�},zaGّBI�j��4O��]/��^P��$�$����C���>�V���ROu���$]�G�H��āg�t��$�$��v��Q����;�w$a��\��oY�=���S��91C�t�ջ�ȡ����8�m\����-���'���yX��>�ȊH �H!�?|I�^)�^BݲM?uwwhP���_�E��{ӦUC��e������~�@" Dq�BI���O���=�^ҝ.�>=�߷�/y����T,13�DQf��Jf̦��m2@Sæi��~����)���{����}d�[B�DD|���8|e͎u�"35�����P��5 w�\&<c���Kӈ��U".���Hȉ7��vhd��ǵպ$��n�� �5���k���2�^6�<�	|�6U"�$"�Κ$�?g�ʄ�ݒ)~��%x�jf(�~Ӻ��ĒI��d���;�R�H��P��#�v"`�ZJ��w��MQ<�uH�����ܢ@�ئ��96g��D�R/έ�&����a���n�#�G��$ Fw�S��I��g�Ǩ��B� ��ӟY.�����K����ɝݳ�
������94F��[+�4N2�.���#|)�LyMA.�:tj�*f����!ͧ8 D�GSto<��3���֌U�O��Q�0��0�W���2�ɑ�܋�ZZ��8��փ���K��*�Y�`���Cl+K�ɍ%����2�sA��`�T��݈���p�V����Tѷ�b[�f7Z��ƃ�5�<h񇆔Dǉn�WR���![yf �Zɫ�W2��WaGaƺ���K��ar6�ƣ��m[\L�2�[����e�Ճ��j�e*K�˜iF��[c�b��V�4
:�n�rY�*[3��s���l/��]�h�����t���^{�eBI$����Mp�|�����~t]I'w�@.#ʕ�r�0$�'�3�&��ʸs���7�y�;KT��$�I���$���I=��>���`�ۼnN��$��wauY�~��������{$&�$�wd��V�yn�˱�Y�G� C��d�M���T$O�x�ٲ��B8b<�wn[��6I%f�_���$�w�ITI?8�"�襕��"<}��n�x����*�eU���%9���Q>G;%(���[�g��O�BMI���f�]��UR���=�K���^BŠ0u�3�ѮƁ]]���I�T`e��4nq��w�������7v��|vvI	$�=���I�T_ĵ��^X���0���5�~�� >�����g����j�_W����%u�׃�?lm�o`;��^b���NW&�B�q�Q�p%n��r�U��媔�B�o/w����4��x�.Ʒ��/�"�
��)"<< ���~�&6fa��U؈����W�D�v����6V��i�HPT�V>4��=ҩ��Wd��ʈtI�KU�W�������{ГTI'�ؘx��/���V��K���K�h��V}��6���;+O�l�H�$��ğk�.���~������c�$��~���x�ٹ�ɷvw��<��
w9��fer����=�56A�nt�f�k�Vð�C.7K�<�I����Q��/��I@��Ũ��þw��M�~^oO�����3'�5b� �2�%�WЍ������,6�`ty��k�R�y?=��Č��6��>9S?r�ߞy�<z�e��q�n'+�g$�Nb�j-F��=�şz��'ÈD^u�Bu2{�'�aߴ��Z�o^�)��t��A��׼�IC�ʗ�����4�2ۻ�+�9�?}�x�x@�n6���٭�u�/�q�+��Y7�w b7�l.7�߾�D� ��d��[�7�y�qvn��W^��I۵"�l�E��mxQ�FzH����3��VVݧ���=Ƹ{?y�
u����t���cQu� �n�p�	b�9�N����k9����h��8��W9ñn��/���r ����]�v�l�bqL��F@��E�vG#���VE҈�mY�j-ыU���������޷W�lp�N��������Crf	B[<	5�ab��yB�]��%�C96<������S�D��R��͗��@^޻����gZ�'%w1� ��	��l�uX	^�Ug��]���m�s�f��%�ZY]|5��i�o{8H�"-�-&QQnu9���iYwYo6���a�#�˻�=}��uD,gpe��5�T�e��6�^u4$ ����pj�^Uy�x��NVQ�~�|���=��Y���o%h\��y��W�>��ûjm���x�_}4\/L;����έ4�7$�.�u���=#}w�ۅ�0#.�oS�S��6وu��|��6wa�E�������y�T�/7,8���@T�=��yw�����Ḗ�g"�W�$;*�`L�5�W�5�[�x�wsLR��0�Ԫ�4r��	8/����`��g�}��^Rn�,�p��d�|������jΕ��r����C�`�f6S'M
��q.�ʓ�k-�2���t�.�V���7�����ͩ[9X�{f��`Ӻ8%n��87,��f�`�/_jc��d��uc�u/�A���;X���:�y����D9Mgu�'^]7��:�)���1�D9�so��*�Ӕ��qU��)2���j��9��d��{��vk�����6�("���\�
�&AU+62@�A�A#�����H��`FU�W	e�^~������mʨ�"���ڸ�F,v�L։\���05ȋ�*�/�w�75�B=r����A���lCd�&.f���\��qr"�\�;+��[���ͻI$�0qW�FaZ��AQZ�jO�ZqdE�d_.��7��+q�H�%�ոM����B(V1�D5�M���V$K�U�$P�[!�-�ʜ�J���[ԭ�,�J"�*�T��4����� ��Լ�F��m��b���)�Da׭�+dZUBH���!H��J�d�@��-�#[*��[@TNRK�ӊ�N􍷋�B7���0��F@\���F���JԂ�K[cA��V�1%�0���ȑ��T�QEQE*Tl�Ȑ\Y!��TnF����R�U�q`䐤��*QXE�$�	"�"��<�C1�>.7���K��9$qDn7 ��#p�y��]F�l�2v��`��*O��>��A�uI�����<�㘵���q1Y�9$q��\[�E�%��wq�����l�/�����u�~�}��=�+Fu竈���i��/|��Op�T��祊|�Ի�;��q<*w����臮k�"U���s��M����o���yF�J�L������t�L�r���9�y���鸵e7吸_��2��\ȓ����}9������6��X�ݑ�\��UͷrZ�.�+Ų�pŅ �\S���|���F�f�&����g\���pS��2�l��m��9�s��;��`�nD����
>�0	>��[�|Ҡr�o��$��g$�b�j-F�{�<�1��bx�p���>|���m���3ƹ$B�2�(��=1�>��쏺 �覆k�ؓz�9'�:�r�qnXB��<�9�E�j-F��j��)���[�K� #�tu89+,����#<|$�H����	
A��J�ҏ��zH�ma�0��d���7�y��)���q����q3�S���|;{�`�K���q��]������7���ܶ���3���R��Y<>�n���yˉ9��$�3�k\��u.��Qjֹ�M�w����,�&#�a�w��3�dK�Ũ�m�s��I��������6��On���cq�Pn_:8�op'@��d�ڲ$�罹kM�$G��u�,>��UwP�}wsz�������{��|Q�A�$IAH�!�|� b���|�7p�my����묷'�穞�ʓ��ù�Gqn鸶]7s��I�u���ug�<ǝλ���_g���}�����j-Ca.-���}�)��<<��jYO�ψ~�O�|$�Hi�
ܠ���J��M��l��V��i�Qm3�)l:�M[]s0,h�1�__�&�=����󧳼����]F���ln7
����u<�q����LWy��8�Q�4^}��J�g�G�l�;湍�ٺ�V�q��J��Ͼ�>'�eM����-��6I���9�OZ�Ͻ�^9�˖�k��y�3�rfx�����]F��j-C���1�|�f;�Q��q��Wy�� h���b8� k]�=��m����"�1��������4��M�>��dr$��ܦc����qj5����#��4���2D�zH��@Ӑ(ꏗK�4�q|�m��wE����u�Spn7,�������
�N�~Z��6����.:��\;�|��<��޻�|#�����j�w�M��w��n%��q/��5�G2�pn\n-�G{�cq{���b^�6�
��7尸coܦ�2��{Ցg��!m�<�g���k��ILŸ���l�[���cSd�������3}���=�\]�#P�w��ͦ#�<�q��������#�#q����7{�cqu���{������E�];�P6L`��R��q������G:������i0���壙7�B���Ө�4�"tIy8�_�DdPADC&q�[^@�&Ѥ��&T�p�a��+��܌c������W(]��録�B�h&�αi4ҦL�[A����j�\��fw9���y	�<y�͓R-�hmX���tk����G�C��KB7���H3M2�4f&ɐ�����E*��%NڷV2���fm`�&�]�4t��Ʀ`���isYF����k�!��!��NF��W���7V�Q��]jeti�I�5��9
�
��?_���0(۷o���K����;��L�qj5��3�h�1n\.-�!qnw��w���Z��<�։��c��3z�2�����#q2�Z����x.jtp�T���K�]�����x8T�������$�H�����]�z��7�C�����n%���K9~�Z$q�P��Gl�1�s���NB��nw=�G�u�	"7�ׂ>�>>F�ߍ����4�v�|s:�5�g�{�s\��r�ˍ�Kp���j56A��-�q�w��=v%t��v�;�� �|}�>�� Ln7_9��8�Q����Y��w�㇉���W߿�wY6���ʙ�.7_w�����M��n��9��/n��wM��k��#��5�r�\�|�y���7.-��qn6�c��S��bo����q�d�e��d��Z�C9Ƿs��і��a\���<޹������Z�C��y��uޚѫ��ۨ�-F�zv��H�Q��������7n鸵aMŸ�<���LM��[���/;�[�?{��t]+m��R��2�v�ne�봫c0��{ns����_m~��J��j.��q<�oY$53�wKq����1���r��nĸ�,��4�}�ރ�>v��e;!��X#��tH�-F�i���\ns���l��s�w��%>�w]�ܾ��z5ʟo����3Ż����%��{�k~�S[�ɜv���K����a�MmEH�˺ڱtJ�iU���e`3fol�J��;>�����6�1��}�Y�O5�D��9�?�����# + �i�&�~�$�S��\[�E�_>|�wp�.-��Ÿ���Ϝ�n;7Kq�pn7%���.O�%��P'ȋ>}$NMp�0��\1�3I��"\5�}���5�Qj5w�0zGq�`\n-F�sZ�[/��w^�8��\n��qn���s��e7����jw�a57ŸY����얶i���|���{�\6y�x(��J����NU	�u�fi"S>~����Ȟ_�����ri�j-GWA��ַ���Cq��/Bq̐��f�pi����2}$/�0����.��e�q=�y��"��n��h�%s7����5��g~�qw���,��e��{�q�Z�M�n7(�����\�29�I�Ov�����2J�fZ�P�ѷr4Ub�Z����6��b��3�ʪݎ��� �̥�}�ނ2�+>�27�P.7�y�0n;��\n7�Q-���h��]K���&;�q�C0�F��F���qw�n-[MŹi�������Oʗ�ެ���FKn��s=OIp�}�޲H�-GE��{��������y�{�NA�n[�p������Q�1�wKq��W|�I@����2}$���۰C���8�YK���#����ti���b۝5�<k�?y���㸷t�[.��9��(J�IDj���ÿ�T���f]���ǵ+FX�u;j��_@njdVtL�%��@���w�b+ޗ��x���D:%=Ɖ7�i�� �AD�U>w܁�>@*	"{\���#�-@�5�o�9��	"w8��x�b�̦�r%C=ϸ��5����kS��; T�Q5Y߹LE�j	"H�|���"	Q���4 P�sf�O�fr.����aBTK��ܦ&���{ګ�W��7n�'q2���x)�&��w�y�D@�w���^��\�dOH��ߜޓ4Ĩ4@��=�3�E�j-F�����0:#��U{����u,����Ł��f�pX�+�Mt5e\V�v�����[�;/�����������'�����L!!�� ��ߜ��!PI
=�9�5@*�d�����
����Z�b:�-��5 ߝ�rH��&�ߖ��6����
������0t@���xje�MW;̜#��F������"��T����0I��.�Z�|�z���\ϹLA$;�D���32����__n_�
�j	!�y�D�A��D�����]kՕ��>�~�G�@>G��z��k$���MB��ZcP���P�?^>Xl�Vܼ�p�;���̗J���M��� Xꁿ@�PI)�T+���P���&���-!�� MI���?�Gu��Q�?��U�y�s#�u��u��1�rv+Fk���G}H��r�f(����yȕy����v*����� �n�5���� �Q(���]H|/^��MĨg���������������yѩ��V� ���Z։�J�H�G{�`j��Е$����^�D^n��5�w��F��vCM[����+)ڀM�K�es���7f8w}����+e�웷�	���
`�	!����u�5��JM߽޼��{���{�|�n}�G��2�H$��m�Ŧ5{�0`<��6�K7uxu��1���y����f
�{[�A�>�ʠ~��x �";���5
�y@\n_{��"{��.1����NΦO�t	�����7��aMі���\�O���P��Qj5��u��]F�B���ۓϊ���w|0|#���9 t�Ԏ`�o��sz�D��8�y�2���R � ���"��=��Vcz���${��9�505��&��w��M*�.��;�d�|9}��o>ֽ�pIi�{�`�4s�ч��hۗ��tc����8D��)�_g���7BT����qM]���L�
����A$4@*<�C��k)q��T�D��IQ*'�׆������s��Ǧd_�圑���cqS5V�9�J��a��j7ܧ'g�7UU�FΫ���Is7k4����̏��1���_��YED�As<��9;��X�+Zn�[�l�Z�m
*�@m�3MU���a�"��.�f�U��92��ܥ�(ײ4m*��unc��{D�4e鈪.i�D-�u��2�mu�����J`b�,[ir*Z� �:dq\��1�6J0pA���U��dÈ0k4Y��K��a+��t�!�3t�vTJ��沬��X�[,�\�u��cJ��M��T���\u�b;\�v�n���ֺ�gW�ϟ��~��r	!�|��PjA$Nv������H�y�	"�|ߒc�U��dxl@�M .�x �0@�_w�W��N~}���u��z<�;�Hp�TRF����w���Lqd<�^`�@�D��Q)��{�%��������IQ��Ƣ�櫼��d_��zȲ �c��b�(L$���C�Q/���7�P�U���5BD�c������~��s{�~�:@*5��)q�Z�L�P;����w���v��m��*`�ʹ �me��$���� ����,�y�Dq�5�T���"%D�%A,�;�� ^}�$����V7��	�~����W����V~��t����;��$��H���\2�hD��c����v%�q�g��N��i.&���Ta��Y$]F���z�����d�%�r�YZ#p���@lt���.�0��2�Rj�.��%�(��K�鵛���?56٣._.f��)pN�JUP��g$4P��E'����;��IW�����������Iq�-@�@�s��IQ*%��F��wv��<p��'}����=  �պ�Y��V:*�C��u�D(�2L�99q�kf�_}������T���f}�n�ff�71d����O.q�q\��̟֯ �E��A�R7��{��E�5 � ��9�!�Q
���s h�̆e�~��}|��;�+�����셭��ˮ�N����{�N�D��-C������Q�Vs^�j�}�R�'��H�$y� �@os�.�Qi�A$;���P�B�l�9~��&P�I�O���~�� ��ˌ�50�I �Ϟs�І��#�w�P���5��R�7�wy���(���โ����mѶݼ¸z��;�C�L�G
�9��95E�;�+Y� �O{�kD�jTA*��]�f	5BT<����\��Qm���QP$~H�nȤR�vH�mL�a�\�����3 ˲��e����s��_~��~0�t��0ta�=�@*	#��7�`�@�D����ֆ�h�Pf�����{��s���כֲH��D�`�O���L�u~��g֦�4j�� �'3}�R��	���`��c�{����#0p"O{����D��C~��\@��Js�W}Ϸ��w�\#�?s�����%Ǹypj��`4@��Qj5��k&��}�>�<	 -?o�;�[u򸝹�n����vl"�X�m�(p�x6㼬j�m�Lz�b�Y������5q՘&�����ס�(����%����w۝���dddP��$C䨅��k���&�R�o���0�����'�Xݮ��@�_�y�B��o}�3��1j4Ũg\� f��JbTJ7�;�%������=�y��/}߹q�W|u�Qi�C�tΧP'�~�j�n�n��z�z���yLA(�@;�s9$K���g%��:�/OxI�g��� .��Ȳ=�*P@�D����
�\Ȅ">;�O���"O��k���R1"k�% �ۛ�y���JFP�����̪%2�j78��w�O�/ɴ��m�~�S<�{���L TZ#Q;����c���Q
�S��v	�`�
K�em}o�9Ǡ���;�3 �+T%J`w����׹̓�tn�]�t�'���w��T�s�d�3�˕.��s�{�3�j%D�����\A�
�w��rH��E�5Ut7���GΚ Q w���(���z.X�����GS	!�$�s9&�J�
�D*�^�ל�w[�����';|�R�-@�@���IA�o�Ւ�rLcU�)��"��@m;�w9^}�x��<	��j7}�MGIĲ �9��H>��ƀ�u�����Ԛg���������ǻ\�
f��{+(�Dni��������|�^>����V.f!�K�1���9�� {� 2
2 ��.G�P=�7��^��ߩ��7K�n��5:��{�H$��-A$>y�ph�����ҹ��w����*%oxߚK����A��;�k$���9�p�Kcpwϐ��-�\�3<��"�,N�Uѣv��)�&BiK�����[��,��2#e�5E������e	��?>�`�N�e�(��	EP���I���Q
��*�ẃ�$���7�hD��w����P(�P��g$��%A���n�e��ݽ¸x����\:��\��ݕ�S{�w�߼��A$�P��g"��0�H}��{ �����^��QT��o��?mxI�|TLn��]���<Oϟ��x)����Ũo��u�)�Q5�1���p�/��}K�ؕ�}��3Q�$�
}���C��H���7�>��mћ��>�����U����~z}�HN���X3�LB�D*�<���B�}��)q�fkZ��{�׫�2!���\;��{ϝZ'���U�C���P׹�P5��Q��#�|��^��} � ��h�юba	�~{�t�0d0�bo���4D*���Wy��j���s�|ũ"!��8Q2��^��:{�w%C�-��N�Oa)����[#Uy���
�m逫N���,H��&Ϥ�u	-�S;�P���sܷ���̢_d�1�˵Qu�Y9 �� 99\�r�L�X:��0�"]K�/�Y���Օ-�{"���Re��'A�f멇a`<�`7�)��AxQ̊��b�U�kiM��ŕ�aζ�`3�4��z��n��(��,�H���m>Qu����z�9���b�N��mM|�$��Y�fD���@@����j�_ٙdc���z�>��Yf�&{n�7JC��_#ՠ�֮Aұ`�궓W��i�LLK�ر��%`v�.M�ns2�㽵�v�����p�9�6#z թn���˲�px�F�/��a��C��-�vBU;=�1g���f��t��^A6�7N�w����"@���ג�y��CJ��:�eBnNb&�"Kn9��髰�iɻmL�IZ�'dg��8�ӽ]�6mwJ���}q7�1eMQn����7�t��K�ǅ&��c�ʕ��+6���A�/k9u�isol�a������x�g�b��M��¬Q��6.0T}���f� fN���t�NM��J�!a�"�����|�R+�.�(ei�.���[N�7�B(r�5T��53.��1��n1���3:��u�6�wk�XC.�/:�nt���k�`��v��{6��%t�l$��;qXR`D�f&!HK�w�M�h���m�._��O�r������[{�� 'B��),��6d�v��X�${w��AS��#\�\ ����qH"�#ZB6H�c"��A����<�\8rT�Aq�I�ʨG	c(�\��j�HI$eH�������#�%ɍ�r��c�`D\(��a$*���B��%qow��uF���!�$a,��d�F��pZ�aD�d��`�S#��$$cc ���V1-��h"U�-e�F����D#�3��!b��#	�%���G+�
[,/@���ap4�jX�(�D�l*�6��11�#��V�W"c%��)R�R��V$B�%�Ycz��% BuH�R5�����L�S��Aa,�H*�Da�p�WF�#�ZH����)jI�� L|��Oq���eK�f�R#j+(�\XJia��
R��T�0D��:��llWi��]�͠Jؚ�i1�YY��]�bu���	��t̹.L�.��(�T��K���UKn���a�����#)�SfF0cb�b�X�6�U�9�YcCք,J�Y��%ł���r[	�W^`Dh�R8 �h�$��Urk���,�@u�lR�Xm6���hVʲԬ#�ü�\��<��I�֑��D�Z��Yvv�3B4�µ�A�A�%�S1SAKvH��"ʵ�κ�Ճ6ژ;l�3Hf�ŢG[CiRR�1t����W�%�0�{:.0���[D�
r�-�
[J6��S�����N��l�5Q͝r��MM�iK2B	�I�[U�ۆX��w8�P�i��н��)ڈĻ�+��w](��)���Yn^93)�56W�C��T��m�8� ��cIL!L��McEԱ����qqmu�F��`�fjGj���چ��U�u�K����L��ny���f�F]��V�F��b��%R4	����c�(��.��L��F#���L�,�e�������k�6��^���뺘�R+X�BkSD��@�)N�
T�ɪ���k2G���#HX^o:�����Pd
YCY���Qof�D��%-�k��h��UL[��\۠5���r�����v	��Te�u��集5�WX��A�t��P�1F�l�oX])2�2&�K�]�i˭���a��Y�L��0Fd&\�:���Z���ئ��!��ڭ��k�!Um���b��%��[6XG�B	m��7��B�@�o=P��0��rY�\h�5��v���.`;Bcl���RW5n`Z)ɦ��iq-�Z�5��p9lW0��՚mn�4��"��Ԧ�i�h^Ȉ鳪`��.�Ur����Af���L&R+��ݦ�f�L�(�&m�jBUv��T<�����$��9ɧ�Ut�ZMtk%ٸ���&L4ڦF�ڗf s���Z�p�XT��t�4�n�)@��6�U$����5fJMlY-н�3t���cb�.�ي��fl���␖�j�4��8�MkfGCd�Y���%�d,it֚]U�sm��#Y��e7;l�&�*�`�c4���.��Q����iX��i�%��*��Vٙt�j�)��#��lMr�,��̤�S.���.Hҵ�3E����?d�驙�d$�7�pf	#�E��Z�<�04��$�I�q��.&�T����ɹ���;�B�j7�TZ�;�<��w�=��ûf�����0\'���=u��/��[���sށ�cx3�DB�p"y����"r	����0�h"�
�P+Fus��}�0{�j%|3+fa�ABbeFxI���u� /��P*-1�������"�F�B����.BU��UW�ϽG�G�#�b��`�$J y�wyK�"�2t�
&�3(׀�0��#{����{^� �zŨ�Z�3�`�A�D�%D���Iq;��A��y�Q|;�o��|��������5��9�w�N�L��������p:����d4�A*�ȅ��c���P�1����9�L<}�$����N� �=��yK�E���@��D��΍�;쥑��r��RR�J��l5�v)5�
�� U�b.ڥv��l�j��}~|��8�l�r'H�y�p j
�H������"��H��`�CR��~�Y�o��a�L����L�C�����^�Ɏ�;�>R��weٽ
�}��raq����
��{���6��'�R�zZL�(Z�z�^� ���5�XL7���+{�u[�+x�+�� �1v&#�;�<������FAY 	 ��w���A$D����b'6R\ T���b�5�q��}߼�^��:�3|� �������������0�����*�J���0gE-FE$��C�3�֫�W|��:�Xϝ���\D���b	 i�P(����5�4��+�=�D� �ʋ��`�Agb��bH��Q5Z�2��H�Q��0f!�TB�A*���� zQ�V:s�����e����0����^�Oy��}�Kuwe��:���;��rc������ ��	7�F2:����_w�&"j%A� �����"H�F�����jgwU�f�>V9��L(���q�⡋+)��nً3շh�p��Z�`�2RJ�0̕32����H�'�ⷫ��*���7������T��B��� �<	5s��}.�� ������I��P;����&�φ�!�1�QV�&�n%C]�0�P*-f�8k���㸞V��Oc���PB�w��&��jTA)�;�y�5���%���t����Q���Q�v����I|������]�vo@������N�D
�1j5��;�A�
 �J�Q/�_�˝E�N{G�v���f��h�7*��%o*Oj�[�/��u�Zn�o��(��Bۺ,�����W�g���=�Q�yZ�|���$����>g�%��D��L=��5�7�<#��F�3� �\ާ'/�c�����h0|'�̠)?�Hq��^b��M�BUP�����")�T(���5�� ����yK�y�sg;����P{��5q*%��g.v���n�0�8D�ϾhtC����}����,���Tv>2�@f/&����Q�7�7�����y�Z�%	R��{��	�!P�{���u�ZM�H�i�SwK��M����f��aK]{D]Kȑ���g8mWϯa��͐[��I�t���CA�\n-F��<����Q��%_�ޓ5���{��앺��,�f�k�w��E�4�(�O~}��w�w�Y���n�^���E�G�����q�헼���o�߀v��N~<���Fc������
 ���o)�$��5�w��I��w���%D������vǸx��N������H�Ƣr����s�
�@1z���c�v|�Z�������`��<" k�p�P�	%@����bj!P�k��ɔ%(�
���z�܅���8��`쾁��DH�{�:�"a"n��򘉦%A$�|�0j-�W���_��>8E9u�l�).��?��͠���u&$v���&`�� �T���ḱ'�a���gV�0fz	�W8n���D$� �EH�_�j-F������Cp
�{=����.�M�m������A5T=�0q0^k�l��O0+�'��?hLi�Th�o��)��-A$
��`�f�8~�?^��a�ǯ��]�Q���%�usVZ�qu,76ܸ�t34�+�>~_�����n��WÄO<���u2!��Ok�u�Ds�
�@+�;̚�jTC}s�{g��{\�Oj�w=��MP������y��p"}���M-��n��l`��o��F��w��%������Y�Jx���@$���4A��گA�.��,�s���"J��D��Ś���+;U0�+��^f��Pw��Ē;;k��_^�d�P��_b�&܋�?Ghӆ[�15�� ����:,F������ѡUصR�J�5SΨ	=�(P�LS����R�i7�EݻTDۋ=�0P���� �ܼ{u@'�����Ʃ.����W{���7�B[��mS�5w4�:�D�Y$q����x������� ����f�9�ݍ��V�vFJ�-�f�U���ح!i�^M/��/��ͺ�ڼ��#�434�lT���!+K�6�t��k��W��m+B��1���j㎶�X��]�6�ZiU����!u�����%��� ����\Mjfƙ6���m�m���h!���i]u�3�v���G(8;E�-���0*��F\1\��k����XSL;4IJ²�^���
�R���4��M��ѓ�,	�E2�������e$lu_��N�ꮈ$��5BkS�.fj3�kĂC��V��_�@%D]�'(ztt���q4��쾦�$�׵@��r�s�7�\�@�~��j� ��:�R���v�3y���H>�n��3�]:����L�QEr��F�$	��.�(��D�O�L�%/@����J��\����S@U{y�� T=�y������J�����3�u`J�g���Z�t�]y<!Q�S��Fr	9��(@�}sFK��Y�]�w~}}��Ϥ�4�����Y.�.�Y��YQ�Q��
��u���7f8Wׯ��X͌�vk�z�~�t
��n������~������nW��R8rX2��&T�w���YP�٦M��4d��(k��5vxl����dZ��C����Zx�i�5�w��켌;1;��W7C2Ԝ����ȉ "�=�	w�7��H�~�s@��C5d���U	�<R&�"��.�m�I G�4 q�{��v��X��� ��s�����PA8�(�T��:�|:.]u�9R.r�ŐI.7.MD�������< �u��fUJ��Fax�������@�z�����sǐHWO.����$<����tE�� 1ԙ(��:��2�ߛ|-˪f��)m4�˞+�6p5~}�>L���Ok�Y�w.Ex�OgmP9�a�Sg���H�ܹ�H�]��2��2�MT�"j���K.��|I�r(��T	"�i���VMuS�GOO*J�ZPvOGH =۪�P�\�ܵ�=W�Fƺ�IeJ��˻��d��GX�ll�뎇��i�tqg.AƬV�]����p�*t�bK���0��D�>�Ed�Q}�k>>N�w������N�X��v�c�:C��d�4H<k�kĒ�v� H=������"���/f�9A3�	HRR.���|E�{b��u	�s��*+jkē��ڢI��߮]�JZ#��DI�f�Hf��5�[�^n�V٭��9��\6#].ˢ�޽{�/˛-�,�O���������9�/o=����&F�犺76hK���P�K
%H+��ƟS�,�g^֛��\k�#9���H���I����d�ǾdNe��[#�8D�RT)R��W�� �{7��`������� =�j����ݐ*����eID̩G)��f\>��~�'�k�$=����>��ʿw�Xn��&�n&�: "�6���F��ğ[40���v�}��]�&�F$p[h�oh0�ꚦ�7�s|ϞLi��g�|� dQ�R@< �'o>�BhL|?BD�0feD��U� h��ҷ&�C�ٴy�:,��}%J VIn�{�f�ߕ����6h��*��5GC]ͨJ�9�qk��)�i��lՍʯϩ�|�؉�HI$�m.�$�o�_��	�빣IY��މ^��t>���ʅ�����H)^>�����D������w:����'Č���G�[}������BI,(� ��i�;��Yۺ��3�l᷹aᠧ� ��^T�8y\�7:"T�����rt擻��h��u^��K��'��� 3���c�_��Av�	��B��ژ�3.>x���d�_ā�sc��Q���ܭ�"F��}huE�r�!fe�3��y.FyI��$JA\�c��s���l7�!}����td�Cn� �}�Wȡ"��� fᩝ\�c��e:��<��Lgj0�b���AR�2�:�H70��6T�[��
 ˍ]sqڠa�X�d3[,]c�(��V�a[3
˖kr��96'i�zU&��ʔ�+1@8-̪n$ۦ�",qk-X�v(h��`g1��WT��L�j�k)��mW�	e[��dliΘ첫.u�p�+�f�3f�cJg2�J�sٚ2�.�m��2��^u`�P��9[������~����L��� �yt�$���GT����̪�j =�n� N�ܑ�A3��$���u�^2vF떺��'�U 4nKa�+���
�
���k��˪�	��	/G�^ב$�v�'�it�V���{]f�	�n\�!�j�	<�W�J�W�Y���n�g*��5]�Α^'�v�@o�`t����.�m�P��6-]�JۿstC۽��1?Nsuq��<�j�B������ɿo���g�1���Sif��(ZkZJ�[t����+���`e���R��G����`��O������u
 GK{w�w|�Nt��;Ā�v��* ��bfE�J���=�ǝ ���Nf�r֌��z�kE�{S�P��w��a/VVFT�=;&�#R��xGb�]��&�_�u��p^�{�d箞d�<���C�$T�FDU�s���B|�|�fw�9�M���z� t��]xV�Tv�*)I$���wTI���Js��9n�'y:I�z��H/����U(ץ$�L����V݌�����x�z-v��$A v�m�#�F�ْ��׌�gەD��^�y��^7f�S����חh��&v���8�.UP�A���H�빢�(�G��}{��FhuGmQ�sn�b�٦���+a�	a�敬��.~}}�=��΍Ew�.y� ���� �����N,��_���'{{n�;�L TJQ�MmH��C�);�mQČ��~�du��k�,������z���}ZU*���Q2�H�%@H:z�>^��ELY���q)�Q$o�d�q;�8Z�u�8�ɂ�ᇩq�P����ɚ.�o]�()���t�aQ��DoF��Dcuu��E����N�q�F��ה�cڠ%Q����x��0"4�H�W��76�sm%�^j�6��N�t��,<Q��2a:��m�y��.�&��L|��)^�/���;#�fG��L���y�v�!<.o4�]V{K���l���f*&���`thcj4��'T�.	��[̨�]By��+(9gVQ!�9٫V+����
`]��*�
y���w����b�+N�l�L!P�Ī���P�j�2L1��0���{��b޻2f�P�Sz�[#"�m[��t^��B�c��͘4oOd�wSv�����va�v�Y�ŗ�i_gc��(VkTv��hwa"J-�����k�$��n9��篠@=�w�zMtħq���J[�TO�X�"$�<�_���c�>�U�ӭM�U6�9n��%�*f����l�/�ojjR���y�,S����n�41e� V��u��$Lt7(���ђi����#n�c��鹐��' Xg�ʙ��ɵQ����s���9S�4蹳�6{�;�=�}�Q)�	�}��V����s1˾=WW��۸����9Yts1����a��J��U��vÎ[۩˂=��= �B�G�Y������O(���Ѷ�a�Ji�����h)�A��@��cY�1:��	�Gv��2/���Q��T>ڭ�D��!	*�!X��a��Eݥ!�aU����".FE��;��D5ζHq$fEV"�HFL,�V)*Z9a"�2�e�p��Egw��N��yj�$qI���"2pV�X�r9H�0��wyޜ�"ҤƢFAm��(��ZQ`��FŊ�Pdɉ$��4�
�{��zɄ�E�kZ�;+`E��2�*Ed� ّT�b�� ��$�G"�Ąc�	Q�#%�LErB�+"�4Q���.9A��T�2[
1)$ƌ�q!e�%�r1�ȋָ�T�������*B�<H�m��D�c"��E"���(�"I!X�l��*�L�"+�$�ɑ�P�Y"A�-���K W*JE���TH���t�R��
@d�b�8A%�DX�I�9QaZ�I���H�V�]�	*QP���Ȭ��	 ����g�}���`������>t�y�RI)=�;�������q�-�d�{=���9۵��>�t�� ^L�șD@�״��W���/�.Wn�c��^�`P����<��'�l�S7��6��7\��T��hطA#��8Su6�m]��/߯s�h|J�������,���Ԋ=��D�"�p���<j�݊����D���I[w�t����zlC��Y��t_d�$���6�fL/�(ך��0���8w��@�0���e�ܟ!@f�P������μ�y4xzCR���{[����J��l�vlʻf�a+�0GdVW�	�ݡЁ��v����&����=d/����l8��Ǜ�M��c{t��ŕj�����X�y�@��Ҏ.HeL�w엒�hz�(|�Ȳ! �w���޼��0*W�T�
I%%~�#`��Β�L�ld��'j{b�%��U�
��N���d?�)����cn�L����(Q0`��#M��	��3�%��Z�rAQr�����L�f�p7Q�R|H7�U=ݎ���r2b�r�b(j핱@w^��X+��0��n���v��w��sۍ�$v=�����b�,]V��4C;�6��`%�oB1�!%*XA=��łxW��]Q[	'sv�	��߬ܝ>�b�D�HJd�^Hy��=�~$I���H'�S�"�xvK-L�:�U	�!>Q1
 mJy`��U%�B\�v*uuT>!��B�"�ߙ`�oWֺ��ӯQ������Z�uvg�fRv�;�y��Փ��Dw�\�f�.vlx�E�ve�י��jg=�p�7��'���$�z�9��b��YRZO���FV��_!��n�XP�	�FUP�F��aWhA��%�Y�V�A���u��r�S]R�K�b��uKV5qьnq�h7�/�Jݺ-]����+Q9%�Z�#LK��A0�Zk��j-�0^�1�6H�e�3��	�9�r0�7͐l�L�>m��s�Ƣ ��3n͆�^vCAh�͝Jˬ�C3f�a�R;%S;��k��Q�Lv�Į�I��>�s�~��y�$RJ���u@�O���vAQ�jzD��_���[o�(3w�@�T �U٫�A�v��rz���oi�H?q���Iʞ��I��o�W.s=`
��ɫ�> �������A��v(
���+���h$����,}�=P*Ⳡ�33�!%%sC�b`af��
y�w���EA����;:�����UA���f�D�H>�t����lpq�o+��*�UI�$&��F��T�{[�v8�w�~��O�CE_��$Z*���F�H�����J.���M5���cnR�1���?'�X�X�l�O��� �s<����n���e��unX�@$�w	�AY1&Y�D$��k���F�8�]DT!����u.�D�ElX:�J�%�'1�a���Z�r���^D�լw����S
aB�.�q٬?�{��$�u湯~:}�|�&�|��cUw��Yov�r� *�I24�2�"�T=� ����M�9�2�B�^Q�y��`'��Х9�F��%E|�u�׸i�]7`���D��P�H=���2�\#3c�Q�ؤ����M'Ƿ[�eVg�\��;�@�On�Q>!�n���uy�1ȃƠ� ��`�4ܙ	���֪�t��a6C=��Imab�v�W��ѶxڡtM������v(Y��=��"A�:���O�G)q��.�n'�|A��k����<UB��Q0z�IP =m	�Q5�"b�(�3�j�>$|���8{stK�n�uؙ�b��,��I)+�����|݋ ���/���.����0�T�tgJ�g�i�zＴ����8��B馺����ݫCwC�8s|��Z����g�@$R@:�v?x�O߾�	���nŕR�"F�S0&QW��v�^lJ�o�ʶ ��+7y݂A>˞��ۘZ�.�Gvz��yDE�"�Y�%E|$��~�@�c��nL���B����IϾn�2��=Y�p�盽� T-$�4��a����L��YZ&k,!�Qv�q�G\������lVē\&�j��$�|�ω'*z�A�n�����N�s�f��.&DD���Nc�p:~��z{� �7�@ �~��0��:\Eç ^x���̥�J«�l�L�d�
�s=��<����"�w�߈>$�m߬r��(�7D�g��IhݿH˭SB�ל�{o�5R�H59�`Y'��O\z���'����xQ��he(w7�"gha�FE�N�� �S�W�V4s��/J�ImL��c]�uk���hK��Xj�+;��o�_1���W�K�� �H����B�?��*�D�3eEx���hO�3�[�}sz�P'���w�Ir�)D_gPQҧr�����M) �A)�p_ۼe���uLշ��74^3�6p.}����f�������[�,�Akf�H�ίe3Z�.���J��`S.{E���E���AT{�!l��m�G�#i+"��dgUx�#|��y�˄���F��^�ЂO�y���|;5˱mЕ{L� AZ�(~����Bs��%LB�;T�H�s;�7ނIy���|y�H�q�9�8� O�%Ɖ���,�A$���7B��g���-�N�o�w{�S����M	�B�>/;��+v�!gP4ZC[�e�%��~N��4��p���eAy��ښL����jt+:����Ա�qF��db��Zk@�Lg[�z���M�ܯ�"Ȅ� �ۘ�܊���l]��i���er�V:�U4�ZX�K4Wb(�YF����Z*KMsYC:�
B	�̰�5��KAa`�qQ��z�Uv)**Mkf�8l͹ ��VE��,%I��L�2V6����RX.�z�r��F:�����2���4����պc��i�v�u���+.u��p�\J� .#&WJ����[c�����ݢ 5�R�Mt��d��؍t�.�����,g�2��A�-��'gyQ>$yݴ�ݺj�)���Y٭���M�����{���@Zo8�N݈�ܮ���F�:�I��b�Sl�eI����.|fI2$��SU:�$�z��ǈ�
���f/�9���Iyݶ,��gL�H��4�ܿdO8�D�ԺŴ���*�on�>'k��s2�ڎ�eP��u@Ruy��aR��K��"�z���o���h�7�|�|^���W,4��j�{�w��t	Ή�6.;"�b�RGv�q�P�:��KD�U���;����J�̓&�$"�I�u�Q$�o���|N_,4���j�]P�H=��W�P���	�A�ӵ�谮���ݒ�t�LO���S�0�d�O���W_!�����Q��9�9�dd-����{P��m�]�,��U�,�Hȯ<���$��{�3z�{�BL]hQ�}p�.�0 L80��p,����M���L����-詪 ���.�FO, ��M�V�VRX�^�H�Y�s9�oeL��5`t �k8��U+�ؓݟ�	K�X���9��"dDJH�.��	=�G�..6��N��ݒ	��@!�mQK���Y��N��0�憦���X���X$.�Atm�*��3"��9[���.y%
FG��v,���9B	 v� _Y�����K�`_��y``~��"���!i%�U�#��M1߱𠉬�L0 ����7�j�����{R�ѡ`(�WhP�W�F��ڨc>���ň�gn,�onyn]��s��n��bnFu�q��ಅ*X]�W�]k�.��a�����W��Y*���N����� �|���z>ϖ��o?m#B�0"Ll�I^9�4�q�sy��>�Ӵ#�s��A罥��`�{yy2FE�.4H+w��&D�*a%5R�P$����mop�'�k��O��ݡD��{k'�r�s��cpG�޽�M�9�"����G`Y��l�A��E�Zڲ��]>�_"�
����a�k�uP$�[���V�iۜ��Ҡ�j���j��KFD��H^fb�
����j/�;��G��j	<�:�`�7G�7�F��G�VH�ߐ�����#`Q˿�yg�U *�Tao�c��<kK ��D�@<�:�U � �b� �;Q�3��aR^�Ƹ�O��λ'�!�<e������u����ӫ�;]ި`�uR��z�٬o�q��7S��Ak �H�����{�^�dԿw���{�{����Ȥ�#�k���dD��`L��J������� �����*k3*"�Φ���:S�$�oc��;~�Sgi��>�>��ݪ�-���j��ۙ���.��`�q]ع4]��{�������T�𩾪�$���b� ���7"�"^��n=Ҷ�ĂD�{��ȕ~�i�B"RGqw���Ձ�D�R\I$���
 xᾡ4�\:f�Ѽ]�bz��-R��(�:��(
'�� T��]*���������7�4H����!����V��z��2�R���$�_d��9>3=9H���'�6�]�4�b"h�	�A�ƻh/^g*"a�ȼ�r	���Mu΂A/3���-�i�]fn���w�tL�c%��7��B��>���˵���i&�	�O��9R�5)�ky��'��1�흜1�}BE	�,���e�S!@�f%fAJ��xy�^��H0X�jkl�ֽٸ�¡O0�{�e+��v�r��h���nf�Õ�`6:���8>]fv�Wt�AwZ�f���Ւoۈ;$�W�r�j�c1Rt�is:Eb�Bh�&���ou�wO�SnY�}0j�Y��&���b���h���^�*���G{tVG[׀Ž��q�k���4oq����&��D�{���#���>���9׷{iN㤎m^�j��㛵`(�b˻z��M��|���(��t8�b��~���Z�1P�dQgG�4v� //�<���V�R�;������|2;�	lR�ʺ,���o!gjli�ٗ��6f3��Ϻ�fح�Q��s�!՘N���q@Y��鸘۽�W���1g��v�����1�v)�`ǵ7k���f��zNv�ul��9a��%�u��0�>�����˸�b]�P�{��%ٓ�^�:�ry]|1r��oxD����4l�̀u�a���ch!]!�cMQ�i��B��黝�"MlI�������V�	��
�5*��k��.z����:�VAx�ͫ��S��WY�E��[�z�tU 	n�O�O��۫+j����&�˭ [Ye�8@H�<��鼷J��> ؒ`������Db�E�e����j"
���k��p�R�*�BY�"8���H����B��e6K��{�I:�[�c�.*��	��r-H�������W
Y![r�sl�r]�wy�c1TH3��c`�@d���Ar�`�*vM�wy�.����V[q�dLT�"�j�[RفQp� EE�Z�@��\��V5�r��,Ȩ��#dRXVI��ʘ���`��0Qk��$[1r�H�C\��!���$$c!�j̒	a&G"�L��l�f
I ���APP����ƈ�f2a#��ɕR�6`Ql%��B㈈�0���E\[$FLQE���1Bd�"@�.2fUɋVAE�FLl\lk#K(��d_����{Q�v�&�\l�ni1�]�{O�V�JGQvp��5��3x�� wJ*m[WRE�hbJ�[b��kÔ�MI�	��Զ�A5-�cM�!�KZq�pDGV2��i���ư^D�2���XWl�Mb4�e��bsDD4vpH@PaL]#	[(���5�1f�=.1���mpi����B-nY�� ����0F�M��B�m��Yl�-m.]���Ci,c\��J�Q �@(&R�4E�4�\U4�]\v�mIZ�B%���ՂЉ���H�Ĥ���FҀDM���e��*��m������KB�K4u��n��R�ݦGD�H���X�p���epU�D��eh����+7��JO&��4"]m��WB%�V�ٵ�	uF=��t�f�و����ٖ5R���j1�B�[��D����#�=K��`Z]2ʎL�[�u�`�B$1�Ł7���n�]X4�W�7��ȢœeKj ZFV:!n�+rSj�k���\�+Rn{-��zk4{[BgF:�) �)]�L�cv6Ym�D�F[ X\���.1�S�s���G9bV�C�H�L���G\�Ƭ�XX&乺�3	�e[���k@���n�X+�"�V1�!l@�\n5"ݮ�v�1l���s+���,itV5�`.��v���YZ֐|Y����8��٫X�-]&M4]L\8BW��mSCK���e�[It{"�k��nT�M�уZ۝Um�p�˅������MhB㱨��5�T"@�+r�b��W��I�s�pFn�,.X� ��KtѮ)�J�\#1՚R!.��Q �	�T�ꢓP�3K�ٍL�ݡ�U#Y���f�FmV�u�b)���f��c�U�nd�iPl�J,����*;V�,.�٣��%�P�:��ʌs��*�UWe[n�m�abʎt�y�Z ��(�ju����n*������}c}]�(� V�!]@�hF��e9�2H�lR�X��k#)Ƶ��f�bR4���mu���3-6�I������ˣ�.���U��i�ee��F�����*J�W�����g���M���F��N����%�]0�� �%����2�cl��u�]Wp�c���5I3[[Ε�Դ�;l��q*�5֦�馦��TJ��
��:e�D����XG.����m��l������e���L���Hy����,��!�{^Dnj�e�tD���b�C�ܚ�%v�	�(2���<O�۔���fwwS��[�����S�����~�]�|��;R����|�H�"%$o 0^e@'Ǟj��|o<���]�X��EnMOfuQT�%��@�!DQ��H��^$񕔈'ā�:��{�����v۫ٲ����<�ם&�)+����Ă@6����|!����^�D�Nd�@]��` =��oޒy��>�{����V�Z��+l��0V��hf3v�����
�**�{������[6HG5�>̶��=�Vj�O6-���
��l���Vh�iU������Y��(��nج��n.��}|�>wZ�R��]�q����Wu��噵���ݩw*�#�W2�������� 	p������@�?9��X ��&�DѮnlM�$��
�IMz+]P��{[v,�b��ʚ��8A�j�����
���)�I	@t��>�[$J O>L$��� 7�2眕��^h�k��ݍP ?D.�t
�T,m�I��8OcS��X7ݪ�>;��ł��8�8>�Xz�����b���u������`eX�A�L\JX��d��ۚ�Rg8mϟ~�u�h{�6W����k�@U	��J��Ɔ��lB&����}:���6[t,�����L��8���i���g���߯Ut�n���}�@��crv�ƾ��142����!+����~�%�ܤA>�U�D]�qī�~����\s�Ex6�ի;�3��_9z����#�ʹ%)7���^;��C�ݔ��%,�q0����y���C����|~���ɀt��@�ӢA���+�����؇������A@|8OK ���3m�����U�>���=�J@�bRF�/2}��o����<�X�)��{�d��vg&+�;*��jo��
I+ V��VBX�f�if^�6xv��ԉ�&����ъ�]���ײ�z5�EPD�9�}�v4���N�����[���+���wC���$��u���^ �3�')�>� �3�t����m�Y<�<��e�\�v��FұWh�+Ś����+Ĝ��%[n�n_M�o�ӹ~'ļΪ��c�L�
R�s<i���g�����޴+Ɗگ |��� ���jQ9;��t`����Ld��֟C�l�q����μ���^�:����b���*6vߦ�z���N�͕51���tR���e�O�~'���>��'xJ�vU�%q��lP����'���7�|H��$���^�y�m�وׯ��~G�m�1��p
�X����F${G0]��xI\�z�������5}z��_�2.T�̤A%�j�I �7��en[�jg[*����=��W�@�]"��UM��wf�`�f�}��������{hY���vIo�ggT٥�蘙�
}2��}YT	"��ز	�;���B-d���{3������yҬ�3�fQ�U�GL�Z��`�@$�UA�}�}B�Oe�զmk���O��/ѷ@|fÁ0"R���vr�~�	,����q:7L�j�ז�8�<	./rj����+^z�������2�pt=Z����No[��I$�܈�,�bx���=�p@vB��R�R��nu��S$</���e5�lbEwi����m��j��B�&�̎��Kd���z� �:�a�"�k	����C]#]���^� c��S���L�ZʶX�%ht�a.o:Ue+����n�������7��޸�cv��4�RTCB��q��͗AL�c�%�%WR�l�k�tLݲ.j�f�:(cͦ�f�K��î2��U#b��˨B,2���@i�#a6r�[�H��V�X���F`t�}������RJR��k�$�wu� �6/�����.m̩g�$�x�
P��l�5+�X��M�s�֚+��b
��(�n�q[-Y> �5�݁1�����%>�g.�"y!
PP�Qvo���3}t ��Lq{w7���߬Hؾ��i:��K�*}���+�05��دJ`	kޟ@	��^{��w�4��^y�� W���#n�Y&���2�"�f�kȂNfr�5bU�݊��#z�]�����6�g:��NO�Mr�hf���J�e����$�SCy���N�]74^3�L�%)Y�L����FW���[��/�Oy@"	$g��P�MO�]���Z)}�J ��)Ѵ�]ڰ���/|�P-f{E/:���H�6�`�km�i�h�i��;Z6o�l����a�=���f�DK���繷xX���͌(��6l�ʻ�M]rŷ��#��������?A����	Z�A7�~���1أz�����(����(Q� ٪�>'��وV�Eo*t,\؟§��:#;'�Ue*V�"`��K1)F�Q�fA�M�Q��m;�O�rn��e�w[D`$��B�ezf'��>�IX�=��ȁo����疮��PD��^6N�!@�[��]�{{�wE+%Ɉ=�r�"�2�ͥnĳD��pX��B���\�LD���&��3(�-�8�cTO�#�7c�C|�m�����TD�:�j%X#��ʉ^5��S��u��&I�p[����6�H<��9Q
�b�S��X(��RL�Jf���v�udw��w24�ۘ����/f䴪%���W�A�]"���@!�/U�p+h�Chv~�$��g,`>���kv�U�<�w��5~�4�VO�}��	#�����M�<Ԕ�^1*U�]�_��(��>U�A ��[�d�_\�1ȭs�]M���v��ԕYJ����랎�	���U�;w�3֠����}�@@�9���6���G�˿Z5e}aj�"Ư0��0DGf�
d���E�q�e&�c�M0�;߯ϼ��>�I>��Ĝ��Y!�ۚ�@��#�_T��9��&�w�}v�ث"��FeE�k�y	�>�\wZ�\A;Ο��	q���Mi��򾏾7��'�W@�%hڠ�}�� ��l�(�Q���2v�<	":y��7�"��ӡwj��i]�/|�t*��vVM�>g�T�W��P��%ˍɥ�hzj���Ɋ��5�&MK��F
�ݝ�4+��]"u2�c���LR���T�'̆�5=4�bQj�����������PH$D�����TP���IID@��*��L=؅ '�ja�1��5��y�<�C�3��<m�*+W]\`���Р̩�D�0����)�1���S[6�i��2cj����r�>z�}�ABAJDp7;�vA%t<T��$�Ϊ񳒣(�g�c�y7�[���X$�ne��?���/�i)7��S�W��͵xtf����O�.���&,��p�����8k++�J�dA�J3(�,=n�'�3�I�{�!v�goF<�c|Y��BA��t�(W�z�H��d��"�����(�v��gU	{��ڴŦ���f��}�FM�Ё��$J��k�+]z��mشvb�Է�XNh����z ���7z�-ܧ�"��e�m� ��� ܎|GR�pѱ��ύ=���!���+ar�s�F��e��
{��6�v.t����܊��]b���H�X�f�˲(O��� >���� �������Ա��Մ��i�+�v�[7/*�9�Ź������PW�5�M n^X�B�֘m�.�U���5q]�5�݆�/�MWYM4R� �b.�TdZ�s�8��X(B�f�-pl��.i�l�6�-apB�p�%��-.��qjb�̯:mh�YF6g+�7Xa֙����V��4.�ME�X�Z���j`/��a�f�&��j��ih;e>�Og��¶�ns�ϯ�� t=��@�H'�w��ܑQ�����؞�OfmP$uZ��(��
P* t;�Ɏ2���/jt���V|��v'bcn.��f��RM�]�*���i,���o���Y'������L<�	��x0G�}c��.��F*ݡB�xd۱׻):�$"H��@�I#��n�Hp�f��=�\���+n����`舎��_��O���o�6R����N8[�TH���߮
3�ժ�u�{����z-׷���Z�Rͨ6�`E�Y�#4&�)�RX⻱rh�3g|�����Utc�������Iw�аF���:Ŋ�V)N�P�{��*
R�o��j�$ڵ �'7[\�},X@W_�s2Y��H��jIPUi2%S��`��j挠R[�rj��Mؔ��,����ŷ���$����� ��������x�|�L���y˻ vdÕ(��
P*"��˻$�^W�P5�%P�����$�o_m�$�w�.Չ2ZQ�e%|խ='C�g{���8H9kv�A�Tv ��z���HfB��nő350d��TL��z(��y��2n�%b�л)�����Q ����%��}MFڢ��*-�u �!,j�6�t�5+#���4֎CWqU��&%;b 3������7v@$��I>�Ϊ%�%0F:{*�ݼTM���12�	R��T�Ut@3�1�WtI�ލ��g���[�^���(���T��v
�y���+H�IJ�`".�{]��TA��V�W���X2��ڎ�(PU�ʲ���Ɉ��N��v�]�b�ND�qe�	�,���8�Z�k���3�p�CGa9���Oh���9a��9�_:�v"��ӥy��2ْ��f�,8�����O��6)�L-���xVEr�XÔ,:�,r��Zw���z��&����!�Aq�����\w�45-��uڎh��7�}y7T����"�M�A���}��#!��V�Cڥ�Ē�����;җg`���J�z73v�^ñ*۹;�{:_fl@����1���9��eU��ֶ�^mo��r�6fYFY�Q��P��+�$���e�6���n��O+*'Ã��W=�Σ�7_p?����V��Vݔ�6b�/���Z
�ӽ�	gΈ�q�B�YC)��)��e8�/.��լ7���0�xk��/n�t[��S�r�x����,(��T�c���H��������*�e.� ��┠��Wp��;��QǺ�؇�OX�;����Rn*���hu�%�'�;�K^���*y�i��Ču^>"U��r��{R�췰q���a]���V1m�ͭ�Ơ�2��v ݡ�����`�҂��5���n�g-S,���wX~�!�NYq�$UnV�"�h0"�s$f7�ȭpr����t��f�m��-n;���3���W6_۩��m]�`�3g������n>&�D3ۑ��$�\\sQQ�ж �I�*1m�JH�7B�m�;Ü^4������ݑ.6Y)Q��f���P)�qL��A�jDinW�.�8�q�,����d��9l�k�8�R*���Hɶ�"�	R���W���_@�����
@����H19�EE6bI20�*Yk��&G�w���	EfF*L�*�Vq�Ra�1"���"2Ҕ�$H���"�bȤsY#�&d�b"� �2dUX�E#2���*Y\ȗ�	�$�� ��2LH��2$L�0��
�""(*�*����`� �"�q##¥j���E�(ɒ1H".
E`ĵQl%)x�����K
��KP��.Y*A�FHH�&F"� �+��b2d&AR8FC\����Xd�bE�6Ė�E��1$j�*?BBE�@9�o��I!>w[�H(����
���mZZ�j�&P��!(�x!�$����H=���$��on�<�
��M�O-+>�h_�N��'�� R��=����2w��i٬9g��ͪ ���I �omDd�D
�zR_f�#K���D%͵�h�Z���GC��u��PI�[���=D� �X切�����o�R=Y�<����Kx��g*5-pB��^7f��~�O���ރ���O���a5�^�>ùf����+_�*��Q��]ۧ{́@���łp���֦da�J��ƨ�=�l�>��iI)Z�Q��:٩Y�x���e�$�sT �׵`��bw��않��C~ɽrC���a��t��˲�r��u6^޹ ��snm�f�U����[iE}�x~#�� h��:�*�=W��ʄeJ�(g���W��{�X(<�br�eLܽ�ݮ�߉������;szy]ާ(7ޠ��U٫$��,cC7ubWT[��4K��K3m.j�m�J)4J�_>C��d� IW{ez��󻈂	���N��$؊�[��<�T+���>RFKVZ�l�Q:'Ͻ�� ��ԋ4��
[)Q$���V	$و3�Y�Z0UfSLDx�h�������v�{�@Q����Ś�z��@�a�۰A>/��>�b����)�m�3�2Ȯ�aЗ1�{��f� w���JV�m]�6T
}��E"�$�jAFv6(�k{PK]LDR�H��H$� 9�6%��10�3�n��V����7�4䩙�L��y�P�hg�*�5�Y��y���,g����E�mm���j�MY�\Ε�;�gw�����F��]Rh�y�!�tBhҠ�d���DZ95�W�F᭡�A�����)���#�t�JܡRj�Wf�e��Y�7mEr��ŷ2�c��:(�at[5V�Q��o,
�l��l����J��.�Xs����g5�2�B�11,p[1F�j������a�ck@��؊0�j�ɝ����7�e�F�v%Tm36�څX����*9K���:�Xc�.MJKIc�s������߿��v\�:\���]��� ݻB�$�Vw�@�d}���#�f1~>:�j�+��H@2����n�2��׸�w�� ����'�Y[�Oew�-�.�.�ѻ�n�P!��A؍�����x�U�;׏A$��¨}w�U�}4� ǣ��S+�wƚ�S��@�� ��CK*�G���Я��nxn31�s\�AW���P&T��r�Aǵ�w�w����B#z��	z� ���h�k�qt��tL�Lz�TL!$%cy��t��h�%̶�؎��-E3�j�>�߯��Z[W?\DveP ���&� -�]_��4���ׯ:F��I$m�U)7R%Lʕ*P(����I+ty�w;�$�hא!A�.�-T�3Q����TN�Q����)��P���U����*�@��gj%��ܢ��3��Y4ԉ�{�o�A �2��D�����X'�K;*������u� ��&���q;{�I�91�8]��^��o�{��>���.���F�
M{Y��T�c�~$��*�xn�\� O�wԁ�xF��'ҫ�W%N;�%%2�t.��dC���M��Y����A��B�IwօoHRr��}��m�Bx�̺�5�T�1Q�+`�6ZZ�`��Q`4�V�PS0�[g��"L�Fz�
#w[�yب�|�-�K�ʠc�Im�����DR����N��?��@����Ϧo+��@����=���ɤc��}���ݫIZ�H��y�� ����@$N'XQ�1�/0G>���"wgg�jv�{3���$�+�r5-�OsL7�֌��dYta�[��cFV�ML�dU�@)+77�ff��O��m��}�Z1�|]���>�uKRa! �JN^ǘ��l��]1O�P�dpP=������w;���_���S"fK
&QQOj�/93LsQ٣G�����wt,��B��P�c��>�^AW�1)x���u����GC�:l�4e.��/̙���+���#��BR��|kv���H5�c���������kn0��<�����w֨OLo��2�Gk�a��?EН����(P== 	=�LH-�y�n{3\�wʊ	 IJ��t������|�Yev����A�N��N�:�RwK�Wv�%j�!�[�֌�X�d*�2��M�m
����H��R��y!n���7krСB�b�FҼH ��Ru���U����WUGd�T)
�մ�Qo�(��p��x���&F�0��e%}���p����+��b����8�|H}��@-�v,Ln{ս��h�$�ɱV����кEZպ$�Y^��0���i�̒��0�[6t0;������\AE�ڢ	3���؅JF��:����ʼI�ƨ�W�d�J��o<i�;A��ҳE��A��n�>��B� ��lX&�]��6��_́X�?)eJ0�?��?n�ݒ}��=���%ˉ��W����l`�*6 ���(Q��ؾ��|I�A�i'Ďm���_Z�|b�l�N-��uR�[�<��U�V���	o��>w�B��wpԉ��27�������63N!z��R���`@���NF�h�g:���1��P���������aџz�)ju��(��(��1+�NϬ{K�1}+��"�<�G�4��5�Zę�؉q�qK�k�(���[ڢ���a�h����B���l֭8��4�� m�]�5��Z��T��ѻ.,؈����2����0nֱ�V"º���MV��b2�Yf�b�4KZVAd�Q�,-��B�"�]i����b��ە�ջU��,Q�;�6Vj���X*�C<��Y�M���DY��fI���g�RmV3T�˽���Y�H�2�w��@$�{W�o�P*�6�̫��Nn��������e@k�yD����`��دĒO�}�/ĝ��^;3f��@���B�pψr�)�A���wd�onh��ѻK�M#]��O���n��8œ^%�o~0R ʄaX/*/��Y��C#y�r�ݶ��buVz5>	�d�V��a 	)Zu��e�ٚ�~��"ѽ�od�P�3r� }ٞl[F߳�u����Z�F͢B�6T.�c�G[b;Y�l@̹&�z�V��nˑ��z�����\�D���G+	᝭D|L�7C[�lr�
K�gP�O��ܚ$Z���`�F��v+Z
4 ܞ�'�Z���YXJ���4�����6�I��s�`j�W���=:۾'�F��%,��PG-�p��Iep.0���'ż�(`�,�rӃ�n���Bb.d�L� �\W������>��ʸO��d*� �p��o�j�ăp:'�#QJej�4�8��h!7��uB����T �[��K��Eۈ�e��f'@Q�{��@��E��}�������+E�ݶ��N�mQ��������,���H)I)H̸�klаe37t#��5�
S�Kt*�b럞����."!)W�wk�%��^$�K{ڮ�Xo;T)��eڢAwҀ$-�3bffb	@�ۻ|n�Ɋ
yآI7��(�[�۰|^��.��܍�~'�J2�Ք���RV�����ʔ>0��'�B�.�Y��;����8���>0F�ڜ3�gQ�vٻ{ ���|��#��Z�x4�U�hdɫ�~�O!�Á��\	 ��U�I-�m�$����eE�v���&M�o�7mX ��ŏ��r�r.�U�;2A�ȩ�D�\���;ܪ�M��Wd����|s�m��N�b����*����u�ۍ�3J6t�0*k�1�)���"ۭm��݀���Ut�����h���h�W�߱���g�}��B����'" �m�y�D�-�m�"���&BD�BR�v��z�c�|�'��Մ�B��n�_�}��>�����
?��q��*��ƭX*�JTh�w~�O�w�B��;\�x�b�c�7ݎ�I��T	J	r&0
I]�Օ'�m1љY��%ev]�����ǜ�YC!�s؍�q3h���b���]&a�h��dbO�Y��]�uE�)z�ᨳ�b�w왶��aY�Nx���crxU�{���@� ��
���k ��b���<O�K��v�Q$l�'A�"���p�)���Q�&��hWVى�Ԛ��#y�8�Tї:ر1�[j���zyĉCFfew�b�`Y�;�^�������ZvhЏu����qP�;l�$$(Z(��6)tM*�	�/zx
 nv��[3͏k���9X,�XӼ�L�v�(
 ����&0�`�9*�;��Hؽɯt@����fd��V��
� g�גo*\���͹��v���U�ǽ9��wF	�⣺[GM^�YH	%6ߖ�6�|s]ul��m��1]>�m�x���c���G��ß�;�ֺqUa8N��u�<#��KG �&���m��aG��YZ������R�O2Q����6���Wy�Ö����;�R�N����] �w��n�Ż`l�J���c���a��be�h�MK��˱"\DşJ����u)۶hn6P3��0���2�j����*�У�CdM��3!�Y�e��Ֆ��]�Z�e�;�p�T7Ѹ蠳n�����8�6p����ScD݌#.�1�e�A�.��!�o�#n6rN�v�e�3WƁpLG�v^9��A�{O���Q��>�au�oM�^�M�����6����F��o%m�(��7}�Q �<��7wr<X\%�
��*�^y$��N18�ѵ>�2=6�B6�(u��đڳ3$����Dхf=���z������}ٗG6VuK	��\j7��(�juf��u�wZ'+�q��Mroҡ���6�w.�v�ݧ+��6��[2�ת�4�ÍX&(�z2`�j��v���72�d��w(��sz��eռ|;8�	|���}�������}�-����v�i�i��|%m�6{��B�b�K�����[���b8��c� l
��s�ԭi]�1��zt⤄�茣C��N����Y�}/�s�zH�0-����?��s;�,�n�[btս2�ک��*0NL�N�I���-�
�F�-�ʳ6a��D��Oѩ����BVx������ӯ��XҦ�ͱI�ǹRKݨ˾:�HX4�fM[���q�;�
(orp2����,��i��xy`V2�|���'o�EUR,_Y��c��W �-�A� ��Im��df#�%�~��H(NLach�AB`�e�*�H�DU��-"�!�]�n��̃��$��H1W"@Qy"��,���HT�X[h����H�u�y�o$H2,���H��4�c2
� ���<J
9Ta�!#"��fA;e�w�H�$����X�NKX� W6�M��2.*k��
6E+�,d\c�6�H���{<�)z��^��u��m�@$KC�z���e��b*"$�$�$bLQb�alT#	&IHH+��Ql����A�9(96�"�Y#1QJ�Kh��H0��.�1lc1F(�rH�rHI`�ȣ2d��DW#��1�H�$��L�H�⨱Qb�"%H�!3a"8Bd�����\ �����EB*A�W?�}����t�xf݆6ZF�r��X�q*i�HU����0�Qф�m�4�\����	�(��Dь�#�2ò�`�Ҥ�^j��
�,(����u�RQJ����l3p[HX9J�R(mV�-q�6�Qz�	*�u�*kF'm�qe��4bHR��'.е�=�v���b���FM*�MR�J(��WG`3�Lf��"Dѭf
A�L.��ԗ�Ɠ$u��kZׄ��.k7;mah0���R.Q@t�X�ISR]�E5�eR=�����l6.�a,8!n�9n�-�c]�e2L烔&��e�A�E�V�vJhf�3&]aY���d�*W+��W2̻j0Sb�����
^.v���2��H�[�G[a-LF7;���5p[�%mJL�-ȭ͆��534h&م������DmsaU�Mqθn-�Sf�%�4�M�2�L�q���3sK1��Y�d9څ��U���J�S�L۞%��V͚R��CYdRf����"�uJڳ9�L1K[�,aZ��P�f���u�m���n˦-�j��1�4k+j�$#+-qͲ̥&�gu�R���R�c��G5٥ց,I�B3Vk��-Xd,�(#SM4��!�rm.��YTُQ`�s,�Yi4Xa�����ם��e�Sv�v!�=��Y[
iS
Y�V��0���]�⫪�c[]�cH\�B-�֦�i�R�0�1�@f��h��a���;W+���qf���0���a�3�	n��8�F�
h;5�5q2cT�]��Z$ųJb����<AK6t[�!)1��Xs�Ét�n�
lr*,& �+yks�;.�� ����Z��`�L���8�B�Xu6�lvV�h@ݓBX�R]m1��QӳD�f����eŌsW	MHM�)�8�0�$rv��;gg9����X:�uc52+��0�jۨś1�n�m�WG`iWvvJ4���һLE�n�V�Ύ�F.-&��:0�j�� c�]-̼92�mv�\��B�aH-��Ս�]%եh�H�-�L4H�y˭���q+`^CR���|����Y��5a
۶�����]cHڣR�m1[]ͺ�j����EX�r�l�2筦4Gdd�+�R�Ŗ4��!]eTmn�ֱ�˃ ص�j���/VRXW6�FfcWB�ܑlu֎!Q�s�߲_�a�S2�#�[�e�B� �=�i�X(��by^����&�����7D�h�̢�5=�����Z�KK��M�u�T O�grI��v,7��7s]ڥȰVs��R ʄalu�>��ݒ/�:MvA�P V��؁]���H=�:��X���S1��`��z������(�;;������vd�č~����sV��%h ��*'��vR��v�gUA'�c���e��i������;�L���782��.�X���	PM��m3h\��ۇZ)4J�΂��R�I*�Ǖ@�o;:�g���8�ɯ���=+#h>�>\ܻbd���`j33(��Wn�_��U���f];S4c�^��{*��`���t�����Nf��2�n��ƨ�,P1ӎ�%Z|b7�;�C���p�DZ{�Gq�>$ns۰A/�h�fvT҈Q	�b�J$��ffQ����Y$�{��R#�Z�S��U�^�>$�7��Y����1 �A��B[6����C�A�T˒1e�� ���'�ם[$�I��(ܾ�ʡ����D%*��y��ު7��$"	!:�$���4�f�W����'���*[i33*n�2j�IueƊS5�!�iQ��5嶭2�]����ܦ��T%�/k,X%�yAH%��cl�N?#��Kfb���P�����[D�
*�4JJ����?����R��7ٻ��I �n*'���U�yĝ)ԙ��<^f;��H��&#���� ��_m
>$��ʉ���0��[]��ʝ����ɫ�����el,�Ml<-ʝJ�-������Π�LjWY�[����֐�t��u"6��ݔw�NJ�7J���A��B��Ϊ�Tѱ�"L�Ffe^�]���Yp(v	S'�S� �r�����e�����/���B�˞>"�
��I���� 3��>��+\-{ �/�P$��u@�O��컮v����՗��v>7Kr�����ڳl9.!`��k�@&NF�-��:aDc�����{��Zkjʯv����@�A׽�f��'�8U�D��������6빡h�hY�@�s��>2�r̉�Q�z�ע�go���Bi��gL^X�Rh�7Eh�	%6�-��(Wf�%T S�8��o^ȥ M� ���.ȩv7�d�"�}{. �+(�S��Đm��(`47ݨ���G�a��v6�����D@Ci��3-`8�5�%�ۡ�r|����(!����w�#Zr+eȩ�/�I��TI��z$I�,L̢_���ŐIw*����EW=]ܪ`[�(��y^��������2* �Q0���si,X+`;/[�IPI�&�ҍb[X�h�1����=����&JQ���6 }�v|	$��T������a��¹��TI'�ג �پ@�D��8 �ƅP�4%�p��=b^�d�@$/���=rhL˻��|Ϲr�bE(�*LʂK0�e��������@j�'��^P���
 g���� >���`Sh�]�M��˱���wI�G��E�%J÷.���/c� �r�� |��T�J�S$Ĵ&� ��q���OS�sp��s���>����	>q��D�z��PSj)R���<�Xt{/��f����eme��7�#���y�4��b�6��u^[6�CzK��Ã��*�F��g��|�O������l�X;��Ͳ�	��Y�-�M�9+.��r8�6�tF��5f�kt�(�nb���sXm���{el%r[���3]�а"���FWiV٦sbd��a�ۙ��`&,f�3��덁�Z�M�MX#6\F��f��U2���r�,veb!miv�ݡJ�]��ť*�j������,�m�Q��J��cl���sj�,Kl� 7�)���+�ǌ<Wb���)t��.f�C9���VdI�<&fQT��Y$��R �OVuW��r,'�B3���'�nH�g2����X��>g�[��q"���=�ɱ�|z��x��^'
y����Osr��{�QH�IJԟ/�����N������e
{p_μ�̀����7J�X��7a'S? 8L�  �}�N����dR�Y� �ՃD�t�h�^�EZ&�I9Z�� ���l��ڻ��S �`���-�H�M�t(|7�� '�n������[c�5]�1a���e0�f��M
飬�GX�d)+TQ6���݂n�P����ԀV5@�s���B�yeGfM�{T	�C2$Ȗ&fQ�k��92*arN���y�'2���\�I� �fY�m۸gj�A��1����]T�)(�+"�t���ڴ�[�.�@���ͺvk�o��$��P$����~>�������Ӝ$�u�`� ��g,'�g7��I��"3z
޼�����+�����,��ټ��"a(T����Vt�ߪ0(]���|�{d�C�;.� 5JX� ����v�R�
TRI�՗d�x�g���nԹٽ�H�YB��o~���OE��4�95������ͱ�t��JժWD4�
g�Aaث5�1y��X)���˳��ݶ|�J� ��<�k� ��ذ�Fvȉ�7~�w��d/����
���l�(ݚ.�&\(3�+�q��G�^������Y������Hz��`'Ĝ��Q�;�M��7z	)�D��fesr�bω ���(����G
�Ss7X^��ꃓjQ��6�ޡGiM��N^F�T�
qV�{m�md���"L��2����Z%XU������}��=O
Ã��W���B�X���8���p���� >� 
�fᆄIW�/^˺�H�3�/�}W�|T�@�P����x�u����lk�Q�YH�/���ĳC��?�
�����LtƳ\�ˬ7V�B艮��ųj�µh��e�tiv��k��#���)-���S�!I'��U�d�k��$�����b���v����9�*&�����^)%|ա�7�Ӑh�y��`��;�U^gP�uo�h��<|�4U�M��,�B�
��S �y����&��������W>�2��<Ϊ&&��&$蘙D
1�xg���Dv�-�XDy����ﵝ�ۛ|�v��M�WS�(K�.f�Ç�J����m����&��e՚!��#��e�{t7����~gW��μTHoL��������ͽ�[���R��O����/3����߅�]�I��*]�N��HL����T�������E��ŉ����Moi�m�M���N;Ҡ�)	B�"32�H-�@	�mߏ-<yڍ�Pn�B�I�f:�|�NiJ�PV c��$�3��45���K=DN<�	 ��{n�)q�}O��e+�`�WQ;��Ax��`Օ@ >��hJ����I��wn��R�;9��a>��9Tn�d�~(�(P�+��M@gtʢ�M�Y�N��b�$�������b��$�k� o�h׬�:&&Q��\�Y$�r�	sƪ�@�n�Q؎��B�;}����th�K��c�v'-��;a��\7a�Y�wz�������w{xOm����~�����lufX�"	�<���MN#'H�� �"�j���W6�ڳ5˓mB	��V������CWd&!�2�2�M��ҸJ�����3;l.�,(pk��H�Z5K�C��-$s4�0З�f^K�x1f�1(K�r���Y��$ٶ�[,�j\�)�C�kv�¨fYU��Z��H96��ؔ���2;�f�d�	b���X6�b���UE��؆1�ۘ�n�4�)�m#���%�tp��,YqX٣����&P���a��d0R�_
�ʰꀡ��P�Cg�:׳v[�?K�7�6� �����W�}%	E T��Ȏ�U�Tz7�6p���鼥��I��dw;N�!In��&���`!(@�P����b�']�/~�>8�Us{b����B��@l�����meJRx�!*��yyb�'��v!^%�u1S�(e<yd�U2LA����A�v�F���S�[����}uv,��q
�Ρ�άDׂ2��e�2�SD�E��� �Kmu� ���V��[�v�B��J��;�DQ&��	{�����X�
�́��鶱��[���y�w��	9���B�r!�("`��
��mv�MD�taD>�B�O!�
�
�gG�9��Ƭ^����61�ƦtF�o���ν�8�;*2��8�L�Jf�ܗ}eD7:��OfuP"���7nzzز�a�%	E �QWdC��
$���Vl�XoL���1cu^vn*�Ay��u*$�BQ0�5��:ۇ���D�#�ZwB�'۹�D�u�nD����cz��$]Q�H�Ax�J���
� �o�W�4b#� ��4׾�}��t	!������j1�9nc���%w,��CC0�%�6��5,fqڸ��6�V����b��U�&	��	�AE��@��5@�I��vem�E�]��ur�I:�i��C�]����(I���7��1�l���tI'�:��>:����{����w澽��� BD�w������3��M�ϸ�xz�`�7|c�%/o% �U�׏<�){`V=˔�1ݛ��u:\�m���nļj˵,��L.��oQ1F��`���F݉�G*�v��N�bif5y}kn�w�-t��=�)�`j���[�F<ٿHЦE�غd�R�r�N�L��������bwf�w�eBY������5��]�.��Gox����s+�t;�����@����a��0p�����:�Ge�T��6�]�p�7Q�l�R=B6/HC)�}��6�Ӗf�|1i<vհ�4��f^�Z��F{$Gq^V�B� �Q�9}v��mLC��XS3`��=)�@�6�ȑӲ�:��|�4���[.�VW\�oq�\c�;���I��k>���,l�h패���г'�P��zP���d��lŏݷ��(��ٕ�������I�^���֤�kyy�LL��ޔ�Dv	�U�*+�����٫�fj�V�f�������x��sC>��v�!
0����t�L��ClNt�7��^�ύT�˟m<n{Q��z�i��TlLVmEp�Х�/z"�6�PS'A^:���eC�M6�촲��˯�����2=�ef������bo���n��{�X�A�9�p��ʏM�[��6��3%�q�m����{G���׸싼[l\"�M���<��ݜ@�`�8*ً`<YaU�nP70e`(�(��d�읍^W#l��|�9�V9�*��YBB#"��F�[!^�j2K(XH��&(�q%��;�8�ّ; ���2=s%�P�YPZ�T�H9[j�!$d�(8�)�Ǎ���q���vd��8�:�2H�W�Z:��c28��-��bF%�pBRR�v[���q�A��$�.@Q�&-e�QZ��\b�H�\a$cٕKY1���Dr�U����w�����l��r@\��3$#�D-�T�F0�Y�d�bXEbɈ��H�Huȵb�2	&.#IC��G"D�E�E,�b�Xń��FH�Ud� �$U0qm�`�!$qd�(�
�#
�QR�H�N8QT�((��AP���T�A����ȤV2DW1!D5������@d ��$�TPg.Z�k��G��rI��Ld��D\�$�1`�D�cq�0��,r(�K+�Eqr$�,���[�2�.,c"$�B1'�����H$���W�c��(J)����;ξ���R�W#i�	 s}�~'���v)q�5�H����r�LB��WH�DP|�@ ��c�1�<T�VŹ�0CY�@	^��� n{,��
4�{%�bf�1b���`bf��q�Ǭen�)a��ͬ	R�b.h���� >2e�2�_z6����ڲ(V�:�NĎ�Lפ�t ���Y$Q�0L��D;��%/;�s����!Ğ��D|^���I�%���B5{�e�1g���m��{��oߝê�|������߆"L�߽�H��IC���Ta>"�
(����jcfi�H������P f{���*��Z�/��$�h*�~�Sh
�zދ�������^L&�D������s=+6�L����G�,�!��:yU$U	ڮ�%mV]�T��%	JS(��"�U�y�>��yahZY>\������D���TX�16�#Nt�#���1ku�.e&T!��U��qW9���Ƽ�զ]�v}}�q�Q!	%$�����ov�^/;h*�5%�Χ�O���	"#�H�F 70%�2��ZI���ss�V\�9*���Y'����T>��ns�V��3'�Vp���&	��	�AGu���M�j�H'Ĩב�i�S��>$��@<�[�i+&"#��&&es<���c�C�C9U��'�ޡ^#1����El���ڝtW��t�HP(�T��y�I��l]��9�/�=kI$syU�I �>ۿ�*�);���bU���]P��k���{,b�d����os�1T@0��J�M�0�*P�oZc��:���Z�k����5�uD�v^�鉮��M�6������.���.���4n@�Z+{ Z�U+�
K���g;%�`�0�D�v`��!�Kd	TŬ�H�v+r.&!�0�ǯZ7�	n�Eq�j�+��AҒ��K���\4���Y�Mԕ�h��3^6����؄ɜ�&�-�$M���h��&��4mFl�)�R�2�ݶ.��7�-�6n����lkl�J��b[Řt�f�PID�2���P��#2���:o*�'{qW�$���n�lʍ�����fr�:�*�!Pފ��D�!$Q���N�`5hO\�H�;�b���6��|F�{d����{�Y}6���l�뺴��Y|�i ���vI0L���K]4�>$w[�$�u�m�ԣ&,L%�"X!>�׷�zAo9�X$�v�H's�lX$��,Njs��)\�0fX��`��vLL� ��ԹزH"��Nb�l,H�z������;�A ��T7��[�c�}�t6�Welإ�ER��F�!��t�#1X���"�ef˦Q�}|��>�ma���R���H9��X$�b��۝Biѓ�[W�@�Fk{v���%	J%	�f��P�o����(�{�qi��m^J���]�C��m�{�gM���ٱK�z�`]d���mCá��Q�a�����q=���A9�_�^�/�*fX��;*�PQP��l}x.�>��B�&qj��"0����\���	��(
��T�6�C.dJ�e,���Q�d��Uo��SN�3;�=��Pa0�|_:���&,L'B�͂"�Uy���nK䝼b*"�� ��b�O���w�G�}���갢~��PeG��P&���֘%c�V��̻�����B1x\Ͳ�s���K/�yLD̢|v���d���
 ����';koF7b6��F�b�f�r:HH
Q������3�:6�-\�2 Ok�@�ۛB�q�]Sevu�j �w��)D�2�׋�X皅@�p>�s-���ǹ���K#y�N+j�o�M%-���Rfژܥ���PYn�o�Ǚ���o8O�gb�Gfy�N�s"HJ�X��p鰄����Qg#�I�j�Q/3�P$���_V�ۇ�UZ�M$n$�HH����B��$^om��=�u����T�㝚��F��ػ��eP��<�	��`H���[��˄�a6�E�v� �Ŧc�`3&�vΆ��G�0H�D"�.�U^c^�}����n�o����^���3s�T'ɰA#�yY7v�
�����p��#��UڼtqX�$�&���%h�Go�ې�D��\��W��e_|I�>���EZ9F-�!5D�9{~[nh�C�'����wU�� ў�N�gĚ=~{rG��}ް�%v�Z#�VA���^�2��TO�G;.�$���=�(��&��_�z����}4:�c�y��z�ݦ����2g��ѤM>y2�*N�E��Ճ���w3�A�yq!5���E]�]�]0
�ײ}	��X= T�"�R�d|�|�4	�k�ʛ0�o��<�jfd��$����ܨ@��RtN{ȣ�.��lF�+_#j좉F��M֛�0�UĘ�0�M�ř�����?~�{�|+<l��ώl�Ģ@��lP� �t�7b���i1�[�k=$ �I=~�P��R��CE�Ap�
"
��i� �ɯ�?��{n	��*N�ۻC~E�u٨����5j��I�d��)�x�t�@	5٪�tI����=�&f�7ϸ�TI>����~$��:N]�h��� �V���ӽ�Dr���֪�����"��+s�&I$�g��Y�lt�BM~}lA���*�#j�c���Ӫd�I�}ۮC�M|���,�M��rQ$�C�Γ���$�=�Cb��3F��_<pY���N�)�pv�M�X�/9wZ�Y0Y�����sso��ݵ����)�}:����?<��{���hy�/��;����֑HB2��-v�Px��`)��l��s,it�m�Q!L�u�H�+��gf]b�hf���3cV����v�� �k4��R���b]V�.ep:��iac�b1[&����%M�9�T�$��R�f�֦Mn�r�
K�/x.*�-B۲.)���f�%ha�E2����i��*�j�|Ŭ�j�W�.J!�;b��U�Z�`��Fa���6�Fc&v��������&� �>yj��G��W���$���$�F�I���:�lOUg:@Z^d_��i��ْBh�_fG���c� ~$�g�+uvI4{=�T ����������/��H�*�+_*Ch��3=�T$�D����}�!�}���~�]�� �4f{cv`�LFʙ��DZ"O9�戛$\����*��:d�h����	 ��^�7Ǧ��I������J�Z�1s�6" ;�����'a��$�;��I4w=�T �N߽�!��~�Q�ߝ�m�±��2%̷R9`ʄ�5���"�X��hӨ����I]��o�*�"�ݢq�2*��$�=���'ĝ��\�Oue�x�C�n���I���'В����"�ҥI�"c�,+�DV{f^NcAgfQ��P�"�\�D!f��ż���tL��fv��okKw�����9���x��i���T�%�{R�4���:�9���[��$�����B�B���Զ�kʍ�Z�B�]�X�ѱ�Hw�nh�VW�t�犐�}��B	$���s�M%�vIF��hP��l�5Oz*�|O{9ʄ u���$�I�t�&_��5E75�KT�9c��WwhP�(��J I��Tٻ�[��uD��ܒh����e�A$��:@g�����>iy߹8ѫ7We*Ll���v�����b�m ��#�h�͙���נ>�P,�/�>Q��$ t�e�TI$��:L��u&v�X	�>���G/}�*C���*ū���c���ӦI8�}-[Y�~��К$�߽�'��uVM��?�$���C�޷ҡ4�����ҥJM�L�	?[�T�d�I�t��'�*��F�wo��7@_��j�WfS�h��u��Ҹ2L��b�1�fs���O,��]q!����[��i�|"#���of�P���>�����R!|.�9�s�"΂��/Wo o����R��I&�f�O�"#��Ō�\ȧ��l�� ȍ�}r���@4�B��k�� �?3��P����s���;�l	D���:$�D����ϰ��]���;���x[1�cH-8�F%l&ae���2��1�ݠ`&ݐ]�8PRbPz2"6K�I)�D�茊nʹ�~��M�I�$׳�$'z�H���Dn��`O�43<�2M=��
��V 5v�״b�IP�g=����b�.;yD�$�����M~=��>��f��M)�]���绦�Q2����{tɢv��[� $el�������"� �&�<컸�*��D�0DHA�B�'��$�}:d ݾ� �h������w{�|1֏C{Y��y�:j;�P<�".J3c��޶c=`�8v�Y|�X�j%W^��Bu���q�uF�t�Q'䣱}v��i(��$��I'��b��07�Y��Rd�Fo��%4���B=w����~j����X�dA+��i�q�sX�&q5-Ω)��qc.��Ϟ���b�
��!�4�Λ&�3��@2�������x�t0-���I� 	��*�Hz��V�ݡB�'����|�䂷�V�I ��I!&�}�P�D�4���u|w��@h�x�+Y@��_�� i�ء$�S��c�mC�T��O�W��� ��e�&�����Wh�V8�tJ��P�o;�UI^�9 �{�rh�;6�Y����&W�fDr�6T��{^��7J�/u�ģ7g�I5��M��t�I��(S�Ĕ��B@7-��$���5U���?q���������*�J��I Ȗ�(�Q���*��W���U��/��a�8
l�E����0�U���p��].ts`})�(?�`�B�&d L@�B�BH2@��?��{ɢq�� @$��&b	�  � ����E  D �@  A � PA@  A �H**�J(� �"� @p���sA@PPPPp�]��Ƌ�@?���C?� �u��4I_J>Ҵ:JZ�(�_���� �*
� �Bn=+�?7��g�c}K�`4'������:����\����~ph+-�~������6��*�}6I�%I�q'ܔ0�Xt�2���ǞB��EA��q�_@�����v��
ҼP��@_��~x������BE	�l`���c���?8}A���>�g��~a?����?�~/���@�~!��� ���*"��ڿ����O�����Č`CG��z���A������i��O�T�"�'��ރ���U��"�2aj�ٴ�O���~p�Mϩ��u���CM$�����R��a���s�e�Ƨ�1���	���� �&lET�TU�UBA yB��Ddb%hh,��|i�)Va��?��H�O�����ܟC�UD��H� )D*�R�RF~����������ho�����p�u���S�4?pi�}T�D�T��e_��ꖿ���)���P�����?�X��7��C��QP\��i�>�����A��?���?��
?�Q����Nږˀ?�~�������~��BN�~���H�����i�?�}�g؁��g���'��q��"��n���gO��?����!�� q�d<#��@}??�I�4�FO͘*�����ਊ���?`�x�N28��
d�>���p�_���y��N��4������PC�>��$dH1z�aG�J��q�|a�� -�K��^�؏�}���/��@���!UK�J�<@1��7������(_]��h�'�L�@(�,
)���~M��?k��}∨-dg����  w�������h����?0�x~c����'��+���)���G�8 A��_����a��ϼ��(�}��O��!�C슸?jZ8?�����P=L�?��DT�?��d��}��a~�e4~���`�H��DT�������C�@�@8h���C��W@��?j��Q?{�7�;4��b-!�Y�!Z�O���F�� �?���~�����6>?�Nq�a��}�k��i�w�G�o�>�I��~A��
�.��?���$>�g�}��F��S���C�ݰ��}����G��H??E�-���4Q��2&>Y��Q&�g�zT�b1P��1�����`��@�!�o��}刺P�?j�(�/�?@~�>䋰2P�~_��9f��?���5��E���M���F�AJ��@��G���������]��BA��\