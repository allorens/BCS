BZh91AY&SY��/ ��ߔryc����߰����  `_�>�^� ]�0&����{qGҀhJ�2S޼�٧y��(H�����}��x��8����r��ڊ�� ����Q(�${aI-v���������������='1��e^`5^��������u�:{`�T;`� ���r}���� v�����'�      @     
������р��M0 &&�0����#B��=@        jy��J�#&�     i�j��L�0	� �   ���@"��D�45d�)�i��h�#O(ؠH�)Q2=@ � 4�<�O`{$��ks��(��X�\(��PP�?�En���(���o����J��.���|��Rױ������������|,(�}#G���h	�lnD�(
K�1�RIAU���
 /CrD��J���   UK���E
�V T^A:�~>���c���G������W�_xs�ο�/��R}�w�Wi�;��֞�󲬕�O\錑D�0�k�L��D���#"%A��ICscq���̝��"gIl�e�:�A�K��Q�dG�D=��_e"�:a�aݲ���DZ��nldӦ�%;����#QD�:U��+�8,�����(J�<����ĿO>�Þ���<Ζ�,�2��QHf�:��.	y0nX���tw��#�'��2�3\fK�/T�j�&S+cE�0�8l��\3&/[��lh�:t㬾N��2D��65$Ӥ�JM���nRm䤩<�wB�t�r䷎W�1�Y��U�-�Wio��i/[{��&�W�oj�gY�f5Zጢ��[����tG�b�[�Og^�Gs�]�=s�7*U8Wa}
�=�a=]Ca�,�K�'�m�ա����p��źfk{��wz;�0�hi`�4ǭ��}�s�M�W�'}:�g��O3���'L����`��H�6��Fԝ2�A1;����t�Q<�� �N�!����D�q ��M�Jh�iMzMd����4�J�6G�rlK�6r�Y�K���jz��z�z�`�CCCAj�է�������MO���WT��X�Y�=�Y�7���7�2�K�Q�Ô.�A���:ꒄ�x��V�N���%�2�g}6������KU�t�[+��0��ù�9��2M�Dj&ڔ�y)3�؛�L��i=�:n�Vo�:���dji�#${4�NdG�:�t�>���WNc+�*�u1��Iǔ�E�p�80ı��K�%k���kV������/�/�ᵖ:��i�M2���Γ��l�Y��7I������o�߻m�l�V/@gV�oe���#z#�o�:�B,"�%���t:FD�ʡ,r:�ȓ[��"Z96'���rV�#�y�Q�"F�L�q�e�u�L9�0�v���lu�]g��r��1-�M/L�f���{L��w�����k|چa�n����q�\��9��W��j�O�_v?�,���}������8��=y���uHY��B� ��]����P�v�|�K-�d,���)���-%pT𖦺(�Y/���]��qZ��7h�n/�q[��M�V5d��e�^��ۺoz�|�d��n�i�Y�9E�,��Oz��D�Ζk7MJyY�9�ܙ���Y�Yxo��j���T�l�Te쳺s�_<ݾh.��T��~+�ja%F�c��9��y7�+[5�%s�6Q��6�l��G�^�E���ի(����G�����o-�e:�F��U�!�W;��08��ᷛ�c�� ���׉��a��:9#|�Bxొ��ySF,i�zvU�_��a�UK
�W	˘Q���=��4N�xЋ���嫷n��n�6eG�tv���$z.t�)���W�桁
{�7VZ�Ѳ�=�텫�6w���O�{6�Y�rCwL�+�b�1$a���e��xa�yꊭ��3�����-i���t�)��d>�gn�믎��_$/ZAҳHAiwL����E���_��χ(�"	��R�

�pE
�%�{c�i÷R��ݭ�aY$�x�V�Y�Ԇx�-Ì���ym����t%m[��ԷE�o�=�𣱼�(�dE�����!���y�o+��d������__,0`1��r�.���.X��8���>�@0`C�m<�ªr�뛔�6�}V�D�M��NJ�3�}yg���*O9;  �0��	e��[˄6qg�����ˇ��9Wt~���'3�r�$�1�	�`>�o ���]�`ݍs{�Y�5W(ʲ%CzhAl+�|�"�gV��=��:����q�&[M�z��cn�ی��P�ΰ���>�I���P��ͽ�H�UC*e���z����9
�a���f��VEV_ɕD�tl��E���3D8�Y(����Q���N̚6�B������	g o1
'�ƣ�O�-c\ɂ����k�-p�4���Xabf�!!ӔO3����T���uB�i�㫍U�p�>ݪ�1������2��3��l3OvfT�W^^�Zp�y���-+�ړ�������m�r��tb��FМ��d������᯲��#�dw�;��fȟ�^�#@G���6��~�/YKӣD�����6�t_o�h��$�C�6_�A�E^�a�b(����VW���,�W���G�o{ܩ	��#�G��m�QT+�K/��UM���)k��E���Wu��Q9��T�*Fm�'ty6(<����fK[��-Nu�U2k4�C�-pM��+k�J��ے�^�yq8��ecӑXY�K��b���A�����"��-6�����]:��Yn�2�p��4ç�E��"/\C�,��x�&�j�mסZ�n�X͕tM:�i�n�Ȗ��w��:AtE�}TTڡ^cA��)b��Sԍt�[b���`&���)Gr�+)X�GeΟU-�G���B��ޚ@	@.��K�Z��й�8�)���Ě��d���HnIcB��~@Jn��(�K�4w����(��d	�g�}���L��"�x۝�&|-��;�w��RTOԏ��}����'�����:<�eI�(�(����n�w���UWȭU*Ҫ�V�Tz�*�սI.�&��BUHV��Z���yy��Uz�wT��UqWj���U\x��B ���*�$(ҦPUphѢ@ѐ�jBZ֧(�U��گ�Ү+N�J�گ^*����~`� $$�d!�Ed�֑V�Q�- �dD$lG��9���U�j�y�mU\Wj��UW�|�h�IU�� �IP�M*3Q^f{�*���W{y�UU�Ҫ�V�U_1�\�Ԝ9Z�ѩ5�]Ph*h�*�3�U�v����UU|�UW�UUToZ4��!"��8"�	 9�_1QUU�w��UUUUUU,� kW5���d9r�����UUw��b���*��b����UPUV��((!4�y��}� (FB�_��}���}���;=<����(��'���\᳅�A,�$6Y�8lD��(K6Y�%�b`� ��<"'�OabB�ؔ%	BQHA>k�j'_,~��^���C��M�EDE$���;ރ���,dm�X�E;��,VFN^V833yݒ55�,>�u��+�Ɠ�L���-L�)H@�G9������Z-�2���dɂʝ
�f.��}^!�c���O%I[�TX��>��fnft���u����a���U ��vg/a�Ee����*�Q�q�M�Np��E,prǖ�o�,�q#&����f
Z��VQ���ݵ�%�K��-��:�9�@���"�r��X��X��Cgo3��n	�M��-%L���V9�Btk�y"T�Ica*-1[�2�a���N;Wu���9���DsiA8������Pܚj���(Î�f��+&@�
�t�S�1Ʋ.CZ�#i?����'\кֵ�kB�kZֵ� 	�kZִ�ֵ�kJ�kZִ����kZҋ�kZִ$p(�h�����=Ē5S�z�e�V��������)]�9�a���<f/Dl��m�ڱ�.��td����J�
���^$�b"�5:��鏉�����.ݢ����S��M�$`8���^���rU�����Թ�B#h�CG���A�Q�w�%�2�V$!���`�D2[�l�h�Z7&�JR�l�B�
9����6h�X��{6�3F��Y*Hڜmof�̷�ͽ��o,(��7udf7G$md��e�#c;A�qmѳn@�����<��od�����v����9���Õ�q��Y�Ӌ���!�ݹ7��&id�f�d���ݙX;DPE��[\�w[\�X2���#Z���a�I*֖m���b��R.�$�a�=�����v��Z�%t��*4Z8(�]�S��&���PE#%M��]�]'I������0�5g
,,���Q1b,Ä-�*`�gK]\"@m��$#�*vA�^�#�͍�\k��w���n�ӄ�s�Eޯ�J��4s�T����@��m���pA����m�+F��H(��B��:��T�<�e$�
;#i�TҢ�錬Zm�Z%�D�t�A*L�A�I�zx������Ѵ8D�����HK��tn��$��
 Q9�u�b���G$( �4�RAK�hcE04���mm�Se���ِ�X�BE��M�2���8���jSV��t��҂����xa(�<G��'��E�&� x�	�a��h�
0�F�`�xQ�h�=��Dlz<A�dy���GI��a��0�6F�#C�
%x�: �$y�#�$@�6x�3��}��=��^*���'���U}��y�
��*e�]�}����:�	�.��A|g�}�A#�u�#QM�|�5�ֵ�k*���s�$RI^)$���W��I+�H�!�$��Y$-���p
�4��X�b�`�D��>dT4����Hr� �m:E!���lf�(��	LD��iu�������1;�E�n�8X�B�J�Z^�B�a�H��Ɗ`�By���2Uk��L�Om�ab'}2��)�$�Bzh��\ńZ9!
5 �$`:�d����Jॉ$^�!� �a�HM����8�hV��K���TR &��G�GVV���&�����2IFB�z��S��"������E���â�]�Y���$"�h"�R^"i��܇pD�d!��"\���ĉD�Pl�d�� l�0ZN��H���b��t�)b%�wGM�BZl�LM�z�9��m�5U��赮w�L\0�y8�6]�rY;�X�H�䤃 �%�,$��%�2�D�Z��O��i�D���!�Y,/D�/e㦅�� HH�2II�M%G,C{��ۻ�LT��;��������j�ˈk	��`��4�m��`����B�5-t	0��/Ls�P��r!.���'�7��t�ud�2����$�a�����a)�f���#s6�S�^io��X�KhY׮�Gah+e�41H�jo0�H0M��%��ʆ8��t��쵴X����Z��a!ϝP�#)��a�+pHRh�isH��s�Ç�w���	����ג��wM��gH4l%i��y��έ�B]&z��YAP�!�Hv�⠣2!�C��mh��4�\��Ft����,:l'U��� �#[h7ӷ.�N�C��݃$�wC�*���ܓ��+)D�ה���iZ��F�J�ժ�>!��-&4�(�v`���d�wgma��@�gi�Bm��B5��!ձ�8m�q㐸G��i:��Ln�p'I���A�T�� !A�HnϤ��[ dxfΑҌ������ÄQ�����:L�6M�AFC�(�0v<C�Dhz�#��x��z3��x�L ��d`�cфX�l���0������l���A��.����7�!���a�ʣ�V���S.Iy��}Jr �ܒ�1�n�7��ΕX���ճ��D��kR�����^f!Kl����&15��$i�l���!������|�)����@ɯB���]^���v�싢�S���e�9
�������CPq�*Y�ь�&���n"b���7�v�F�k�$�(�{_w�=$rF��G$c�G$bH�	$����A�������,�mK�͑=ř0O2��Hնc��ex�Ք5���o45�m��#�w1߹�,p��x�t�W�)pV�o�ʃP��EL_�#��r�Ъ�N_�i�M��(:ur��@�HƛY��p��X�l0�����V��$�\<�A��m�p��ToA��E����e�2�(4�3@�
�ٗ�˥�S������H�Y+�\3�9�J�L�UQ�sf�N��89x�Cma*g	$eXXeE�)�h���xj�~�ί@1���B�h%Q����6zN�A��˪[t����H���(.�gTqJ ��A%��L�m��&S�K�֞wt5yi$��KB3&���V��T&5k��k�Aj%@J	$�����٢�"pg�x��n��wɭ8"亁���r/s+[�d1�J�V�9�Q�92Uݜ2�,�,S�.���oW8����ޓ;e�4F����<Z�ֈ$a�`�B���!����3E ���� ��RD��n�!�(/Iʐ�Ig���-)�whT�`�މn/7�Wyw�f;laܺVL�n�V�kr�e4I%�� �-���ל�#�Q}E��9l-*
4hr^0/Ԅ��l�&̴�*.��A��+�Ɂ��Wnv���@Β��$������ɒw��z[\iA��T�-[M��鸛*|H=���B�e �N�қMo�l�Px׋e�!w����
����	:��u}? �x�'e�
�+�i�U;Ĵ$��
IJ����qqk�0*ík�'D�AB�)�,,K6�z��)�I&�D��#b6 w|șʡ��w��
)F�8ID�X���=��mb%(Ki�%�8���)m&J���N����$��%K�	vs���|�yp���&n�%+�����!Q5�� i�Æ�J	��-4A����	���`F�C0�ǈ��x�VA$�?E#ñ�kŔL��4;4F�$��Ğ0���=����G��6a�%`�0�yH�H��6ag�!��左�|��r���7v�0�kv�U�b͚2:UB�QUD�ڠ�X�t��G�>���O]���^w%w)$��T��IR!$�"IRI$�I$�Xa� a��|�$|����*e:�[�1�Dy�V��\[x����CFH��k!��$��ݢQ��B������� myҍ+AE���bw��l��J0�D�l-]��ڤ��c3KmXBҒ�
�tV�	�F�N�	�X�B)baC6�6��kѰ���6�ѣ$�Af����%w%�)�Z��)dRETT���D�!n��b燍�omZ!�n�Hm�IU�L��;4��,1iq9�T���-n��v�m��p�D�ͽ�f�%��������m1Ю�i�D����R:�h�[�xH�(�$+�#��͒�B��6��ZE�ٍЉ4B	Z�B�
E"�.\��;��2)��PT�n�&�������P��E�I��2���a�2g�h�Xѝ��p�i���f6i,��s��l7ڈg�I&�7��E�-�ғ �����v3��(6aI8�a��
в��@�2��o�nN�䌙0��2�4X&u$��ƩV�ԃ��Ŷh�\J�١�*�)5F���G��d�M�m�(��<t�C0,u�L��
���j�)By(�AJ�tnƆ�'%�8��RLD1�%�1uh�B�R3��I��8�N�6��ՌTl��JKF�8�g�U^MX���!���$��Y���b0h��h��W�Ğ���+ѤѮnL׶���f�*��)�M��K,ޭr���ӂW�`�X�U�Ν;�D�I��X�Њ�6:�9��*g%�(��F�瑱w�h���L�d������lh����R+�¬�d��	^$�9��ݔ�F��IA����=0�:h�-j�Qob-3̚m�SN�6<4?(X2	�	EͰ醱Iې;ld���v��--�*O�4��ܝ'ő��p}<t��Q�7��0�"IFQaa:��(���6;6F���x��Hä`���xx�O��6?A�a��&/!�R��L��pp����F��q�}$U��X�sh^/2�X(�H.]�����u..�#��72ؚfI���@Kv^-s�ds�2�Q�o��|�k�U^&��0C��J�v��GPBS|��E�SUWA$�>�E�K��f����,�gP�˺Ѯ�*�gŒ����c\\�u�U�ψ,�D���Iɘ�J��*�菑Q��O3,Ȥ��M^��D ґ443hTJ �J�WXRKlZ�L���.I$��$�d�\�I!�IrI%�$���X ��� �}\U�	�ʵ�q�a�&1y奕o���#�缃��.���;V!�!l��c��@-8'̻:<%46�@��.�����Y�x�T�j
5$J�'���fv��ٳ
��r��qhF��"ͫ�:��r#��53%�Ӑ��d(Ѷ�?C�MR)h�$�$�����v#n�8]�2�v�pX��)�K68�a*�=�<��Ak�#y��-)N�K6p,,������(���՚](DU�V�Ŋ�y9�6�Jք�j�kZR�-� �X-%)O�	�>zǲͦ�:IAakp7��l}Y�uh�`�0q��1�G;�i����o�lg���5�.�يU�vi�:8�Q�D&)+g��6h�`�,�d���m�Ŧ��@K9�p�C)�#73k!��f[����&K�3��Tȱ51�ȨE:.��@�3��1A����F���Ȥi�I���<����`[�nV�.q|�j�+�+��_:���I6%�r!�bܝ�T��^D���5D�U���~<��%����amZ4yF!�K�����-�2ʵ($�XY�}q����8�)d��7�u���Ƚ69C\ ٱ�����f\��3��Ƌ��v�H��
=�-��h4O�>2�(�(�m�0�m�*[��ݮb�2�6b%Q�Ť�o%�!g���؜M���d���n�cGl)��M�nL�6���,��M�ߕPФ�ǍV`�+���Q�qi[��2�_$܄���6��3#ڥ(8� &\DqiB��`�45k�Q�z�n\6ۇ�4�0R=���ś$�XY5m䖔�&�$14�,�t�[���QxA(��t1mT��#�j�;eʂ���
�<�B�<)R�T��h���=�Q>�'����4a����!Ʉфv:"�#C��9���썏F���z�x�<���#��I��?G��EE.��H������p3�y�r+/Oor�%�L��O�ӅV.�Q��k��ȅ��>������ft�I �I$�I$�I$�I$�C$��1�c3�2�IT��ș���2���)�x�!Ĺ��,�c����$�ύ���J�-�8A&��h��2�ED*ᣤ�Ph,�L���YM��6܎M�GI��p�0ƻ[�EpꡃXuAf��w��*�X��ˆэ�4��t�����ż#��i���<&�����v�!���vIVBQ*�"m���l���&!Z����fѬPI�T2R�ɓE3���,kz�Hh����b��ڃ��̿u��c8����<I��Y�ޑ�҃JH�,�+Q��	$��!k�.�(0{F/'Cm�!Z�i�1�&3��d���X���N9""�]6��r\�71��ӓݦ�&nHܪ:C����$KM��#j6Z����=9H�������%5�0d챀�]��:�B%iy���qc3��Z�;�jOEd��(D���۫�����*��K� ���p�ߘ�G�m�ږ�	%;��
����6h6z�+�S���j�~W.��ǳ�p#C"��
)���ѝh�典��X�P��^�J(���H����� �FZV0X��1�ܱ��n�2�(�Oh��ZZ6AҎ�y�TU�{�MC���6����괜H�Y,�h��-*&`q���YDAKݧ�&T��ֻ̣��Z<IdXx)V�hC�"8�A'�����<��J��4O\N��6�F��f�M�Ԕ�l��h�J/Z$w�&]�w��<s�L�;��%΍��V�驣댌PH�
8	�$���A�(L��;x��7�w�\ˈp�U3$��bjB[�,:�6��k�G.�8{H�S�5�S%�� 8W�F���tA�v>�#��K��H:a:����a�Q�Q�+a2aD��x3#Ѹz#���l����Ğ:G������������{#c�D$�����(�rEQ0<V<5���������E������K�8.���D������u!�C/jzJ��Ś[5�&0�ݧh+�V�?u�+�%�Kţ\�]�w;JRN�˖�B((�]��V�c��i�ዌ�tO�S_1���f �+Ȏ݊z�e���#jR�R��e�|��.*��A��.-���9�RD�W����$�	$�I$�"�I$�I$�I$�" �ɐ�:��>\��xT(!��)��%�BC.ꁰ�L6�I�[Ui^��2����xy�\U#�\̎�����#�
�DA�~v�K�"p�q�o��[:6A���M����{=1����c�"�GiZ4���8
6���`b��lm�n%�OSGL\��o�5�z�H��/�\Q�>�����F��y0����è�ar�S�3g�����5��!��\�&��󊟩�i�����5���6XXQ�ql�k8��$��r��_F؛���׉[N=\�YI]�f\NǑx��̆��������۞���ǽ�ټ��ٱbUW�ۓ�'+Er5Ta��~��c���{�ͱR�� t���6ݶ�"�Z����ջ����j.�R�iZ�A��K��玘�!x�7|��w�n�{��4�q3I��g���4L��:ON+GV�Z򒑵p��f�1�qB�/�"G=�Z�M�fe�����l#k˒yH��tth<f��u.n��&vL��H��,�v���pCP@1�Kj�Md��v��o6�a����BY���'�M,��IW�,q1`1m�'�6����UKt�A�..Q�%X����Иq�<6�	6�)�vԝӇO}�ҋ��T7��,�,�]u��Ls�(�mĬ��M��Jn`�}������)1U�pc�~�����\غ�i��~Ӳv�V���2�h�u��͛00$���h`�4�
�'@y1P�q��h�Y�L�h�9G�JWWW9�?D�YD��A-I/b�K�	چ=�ȱ�G��a���xa&�&`��0�0�(�(�n�Q�aa:�dP�l��c��p�����>o��x<������p�#c�D$��$x92�&G�&Klx��%oȃ�J�/i��D��,��_gsƖ7��ޝەH]�ZK��&M���V���}]�$�I$���I$�I$�I#G$�A`XjJ�m}���Հ�S��4��v�<	�<vs�I#i�G���K��ͣ�yUR�|6If��I����TJ�#)ak��U���ٌiƬn��9�q���#���c�FѤb�0��q>��;ޮ(W7��)RF��,�����8o�̎ �-iȝ�a�um��9�c�� ��Ch��F�\��|[]��ϵ�I��]]�a�:7���n[�#��ί,����t�f�4WL�.��.j�Y��J6���ť�i:��A�i��b5Μ�j��9�eus�\�1�v�Յp��I#(qm�46�d&��������;�뙂_&!�'dL8�m'�,%f�WT�ҕ�;ռ:��*0�`I�<pѵ����j���[cq�5�ŪX�<����8��i�1��t7{��x��_���O..�Ԣ�~:-k�0�� 6)#�M;5dS �������LS1VG�y�#�ڙca�H��3�D�^ͦm����ӧ�fS3*���13|qF�����x������Q.X-�e�y$8Н5�m7��!�),��*�Q�:��pL��b<���[m�ٳH�Gml�e�h<M|8榕s��&��=ȇh�I�B�R.��P��Akt��F��K��0�'�m�e�-��[�J?W��;�e�kCsI�N9��� �L���n%���69I<=�xل�xfd�2�������VDDX��0v6aA���=#C�<x�#����~��`�x3����=��[�$$����&C� x`�jb�L�}__�ȶX1۟��}����r�����&��V���(�B�ˤ���_#�Y���Y����K9u/ b�Z��m*&��׻���-2n8��,8�t���e��JB�ǗY^�rY��n�k&�sh�0��7�E�汩*
P��\� m:�kB��`���[�����\U{/��g}I$�I$�I$�I$�I$�I$�O@���wŴ����PK��v��R?%d�b(�����$�#*����r�ojf^�H�F*�j�'����E�1�r̓pX�6�R]�[��rV�[K(�ɯg�鶏as�Rԗ:���
N.Qzm��A �J�|6�F�6d6;���l`����$py�o�����*S��o�6�ǎ,\Z%:t��۸��F����[Om��bHI�8h,$���L8�s������I�mNZ�꓎����[g��J���k}G4l�l$�;Ѳ8��\P*2$+'-L�v��|=�B��;4��d�s~Z<�#��mu4Qg�EY���QK�B��7֞l�0;1dE�}W�ڻۖhN'4�VW �.��� x��\��v`s+����ҽN������ť�D��nΞn<�yJ/��S
�#�H/��y���J8 6�:Q��Zc[�-��u���&��B��d�!F֚8vtJ�e+��̼��i;���=�Gf�����*E��SjN_�ҵ�HTo��@b�Jѵ�e���f���A�<``l�}4Ce��wU��*�P��q�x�oG+�;�ޞ4^��͓��{fѹ�ot3����Ւ���p��$x�P7��d$�eb�2Rb����H�R�PX��\�4��SB���
�h�iѴ�`�i鍘b��=�F4 e����9D���E�c��&a��5��bs�׈э�յ�u�勑�;l�2�;h۽&䪕�l�������|'��A�0؜6"pHlK(���%�4a��0�L0çN�4a�F0�0�0��tc:h��s����y���j��]+zn�z"T�GfgBE]��ٯ�^��ݫ*�"�E�����wl�|��o�K��*��3#�v��ewk���8]���D[2.��]�4w@�x's��r*�wuk���ӄ��G�.ʴ�ӎ���|1v��;��|x5���n��+X����(I�7+o�I$�I$�I$�I$�I$�I$�P"|�)��j���:L���ǉcsU!
d$'{4�Z�h�xڒt�q=B�K�HY;�NrΖ�;pi�N��l�X�������rީ��<yA��r��B5K#��y�`��"��R"!Ee��]��"4�EVUd�R9"j�b���Jׂ�����C�#�m4���ݰ=i�[�{^'f����ᢈfvJ*hӆ<6�vd�&�5�n�VT�L�'�d!��p|��6�Z�F@�:��uSZ��3J`�f�l^�x.�Wn&PDF���D&�{���xѻ�&��N6(��b�+o;T���(j���X��Q[\�v��m�'m�<�:0ӂ��rBM�X�	mDם�&�9u%�nJ��16�1D�4�@F�J�cl���6��	�6n�m�Q�J���&ݸ���C9/&K�;�Y޲�2��H�=d�p��3R�Lj�8�B6�B0��FC1R�,F�J�:{K+��R���Yh�{<I��^����d����I&#�r������P�m�oNۦ�y�̦�X[\$�!�J�N.���S~U�)*�1�āD� �H B�d/�4��y�G�b�%Yib=�>���������hd{*�2TI	$�A�  �bQ�~��>���%����dtx~�,^�
(��-�T$@�1.3� 蹫��8�f[T�V@IA�$I���6P��h"�"� ��0 ���� AHR� `@� `AH�XT� AHB� E T� DXU� D`A`E� � Q�XP� A��P�
���"� 0 ��d���PHH ��ĀQ )��@i�B`H�B�	��L���ŭcE�A�2� �H2��1�D� $ F H��k� FH F�@H H�%Ah�D�`� H�D�����	d���Ah F D��PZb��AhH`�ĀE�I	7EK�� �@b@"@bD�)L,@"@h���@F`BH�� 4�!�IA`$HHH�F`�`�`B�H1 �a Ă! ă�J��.H%0c0c	�0cA��d	"A�c #0#0�B0B0bA� ��#0� �� ��#0#0X@����$� �#0"A� �	0bA��0c���B0B0c#B0XB$B$!0��a��"@�#@��#@�B0�"@B0�!���$ �0���b���b0�E�&i$B@���� A���6F� EHB��  F�Z�ZBBFE��K�m>��.�I�4�^���@uk�?3�%�(
$H� �F��|)*Ǆ+��5��k�9�>���g�y~���a-�r�{L��z�<'A�~���H���ٰ�Ô}�C=F�p���x��������諸�%1�)}ޒ}$*>�F�������|����%�Ӭ����(� AC�D��� �E����9!��[��}�
/�� �EB?�! ��$"� P��/�/�=���~�Le������=�D�O���=?���9����Gg�|�z}�?��@tz��C�"|6~H�(@������T�H��9�t�q�q�R��l�z��bd����?B[�6'��%%%��x�PcF���F6�5����=��:�/ׂ˄�0�F���'�l�����)0���U,b�}�ȆB((��tB�D��#` `@qv1,R�R���*T@�f��a����(�R��.���86���s�<F���0 � Q��(H�� B ,�"�PEA�F 2Ǭ��A�>��=��`�	�zi�o�/��"d.�X���1?d|Q �] ��Qa�D,�<O�B'��YE�2ߑ;���  �d����,�����?A��&��=���Cײ��;=Bh����v�G�-� }�)A���h|��	�`���A���~g�C؟"?hy�[�O���}3�8}�=�򢀡�:<��bY�oW��X�ȯ���vvh���@>/�BQQHC��,�"���(
���D�����'��=�k)�,���=C�y�!G�p�$,dC�ƄT\� H�$"�6$�ط�B�C ��R�P�H�}ߖ��= �D��a�c��
T����R/��� ��N��NP�h��r���)b	�p&b�	�P�K	Cװ�����.|O|� �{�@P���?�`v�����<�XCݗ�PO����������x���g�?x\l%�OOX{S�^�|��HD�=c���������"s�������v?�>�1|��?(���qmOH�%HA�0�0W����Ԋ� |���NX� ��� 8�~�<��=A���z��'�G�A��O-�m#T�!�>>�|���`CF��,!C=�c��
=d��	�}"��I$�t\?��~�Ƀ�8�6&�2&ȟ�>>��6����A��-Q�-�by�����j�E/��2@����G���4���! �6I~�׷� �R��$� |��bQ�/���'���Qn�kw��|�p��'�'���;N��t ����=���p��d=��\�F�4P�灮D>9���g�	jPP�̈�_�����/�.�p�!qz$^