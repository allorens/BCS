BZh91AY&SYn֏���_�py����߰����a	��    :   l=d   t�� �B�          P.�4�   � 1����c0�   c��v�/wyz�F;�������g���N���������;�jlk���/n�����������}�z����{�{����s8뮐t�'�����5�����m�5�=��� � 6{����Ng�<yz���6e����=W��mv6ܫ����ss��:�c���-zש��g����x��r7.wv]ˎk�ޯZ�w]���9]��7t�����[��a�Ɵ@ ( G�/��[K�=�x��ݛ�]���]�����\װ���wV�v�#�F����=Xp�mݝ.�.m�q�`6��ܽٱ;�{����G�  "�+�����s��wNv�R��&u��tƮt3R]��x ����{�^�{��}�]���^w�8�A�y���|��{Ou��˼ �=  A����okM�����m�׻�9����]�=��w;wwY�8T3�{{�� =�ݾ�>�����s�Wp���d��W�                 @�z�   �         @ J��7�R�D� �  	���S		%)D4� ����44d���B4��3I�`S   0T�""��Uh444   M D��hS�i=S�i=���I�~��� U5�J�!�2@d`&��4�����A��)�ڛݻa���� ϧ��Ϲ%����ͱ���l���o�����~"�7�����v�Z����������l�G�c!)���o{f�3�>����s�\���1�h���>�$P��Z�E����W�a�?7����[��_4J�<7����^�-r�8[�&a�H�yߊ���B	6���D����}�'Ӊ7��I�؎���	���h�C�Pērd;A���jM��:���c�8gy$���͑�4�F�H'~rNw�d�	�d��NaxɈ���,�7>�����ɣF�'��2h�5d։��h�	������И�evY6MHm!�KV��	�Rm5�4a���$G�	0LHgɉg��KM�ͲP���GY"g�"aNH����D�La3���a:w�bl���
Æh�w�D��I�4�:= ���,�hӲU%Ĉ������H�1�>�͒��$D�"u�(����n	�H�,�ɄĘp�d���5�"Z"u0I:H�CZH�H��e��舊p���Z"bYC�DI�;'ɒȚ�&�"^$Å0�!8�����DI�6k�	ׄ�f;'��%�+I+�)I�E}�D�"j(~���$N�xJ��X�����J8�&D�h�7	�"X�0� �`�&��%�'d9��'ւuN�p�&��"u0��G����Bh�&��"`��8F�f�M�Ƥ���M��|w�6���D��O$N�0�D��a{�~0�,�#Ȏv�s"pD���N����'hG�99S���7����K)��!���*'GS�ocS����Å��%:�G~�ϬF�8H��t~�Z�ϑ�BsD�,���~��bfN>�kj�ƾ>z5r�M���ӿ�\G�h���q�Vt~�dџQҤDyuΕ�#�I:'	�YZ;A5���tjtΜ*���T�L��n��<u�N���R�%�f�p��'bv��$��*Ěv�<jt��h�!�.]��*�ZsBw�,uڈ�f�|�5���bU�g��#�Q8m��ʈ�:Y�}�"#�����hJ���:���.�#"p�����uQ8oq�TD�':�P#���"p�AU�&֥	���S�E�F]JL �TN�Ƨ��L,vH��I0��j�"��a��Bs�NQ�C����˨��*"oMJ ��&�3u*Q�2�'6Բ'Ȍ��_H7ʉc�TD�ʖCZ�"<�DE�D�kR���A��pӪ�#.�#��T"kmJ ��#�TD^ԡ�9���y>G��4M�e��Ds�0V�w�8kiIӝjp���?�>���7(�{>G���
g�;��d�J9Bs�#&�З�;D9�,������9SGuҸpy¨G�N�j#�Ʀ�NmM�"ϧQD%CT;��� �|�L�l�w�$��8O�y>A��϶ϧؒ\ѫ�D{6=����.L;'�Q��R�t��wmN���Ĥ�%'r������+��G�������"�8��˄��oe�����y��8���1b9�l�6�KZ6!�gֵ�r���|}�k�>�\�ktJԝ��Q��<�G���*=ʉ���&t��F�u�� �u]G����{�[ڔ�̩VI�$y3�����{��9�;MO�MNT���j.�,�����kRUԨ������0��Le��t�����|ӅI�b�'O���T�����2�K�$}��w掮��d�mD��'z��=�*F�s%�I�M}&����9چ	��N��j]K�M����'�Iک6k�T����F�Q��<�9R�gmf٩�i���7��I=�W�IŎ��3��6H�r�Q���G���wMNT��jq�/��Ծ'|����:$��#�jsR���ƾ���k�y}��y��ȚU$5�W�9�>�$|�9&��:�(~FDý6u,�D�Ҟ�fȖ�\jP��B:������/�(�D�ڮ�/�â�+"Q�`�D��_""r��c����A)�NԱ�&�W���*U�DN2DG$� �"<���8h~�8:ԯ�Ȕi�&	H�����Ɇ�R������:hJw)��".�p�[���K�+���+Q�J��YDϢ&�JD{��O��"iܤD숋�XX뒾Mh{6"k��bm�k)8oL���r�4�R'1��F?L,u�_?,�4i�"[�H��V}2�"iܤN?DEԬ,u�_?=�B&��[o%"me'��|�R&��D�2�h�ۘ�(����ȝ�V��>�%�&��܉-ʮ	�eP��ԥ�Y���'Y�U:rM;ܪ5�<��U'���|ep�/R�sf�F��v&d��ȝ�V��C���r�T����Z���5_W��F����H��ep��#�+Ȳ٭'(� �#ɾ#�/�t�56%��V���`�j�C����)�9$�l��d�rʑ�9"9&�ʮ5Tt� �%���U&��ja�A�;�$9�9 ���SY���oSV��e0�K�</�r	�&A��T�ʕ�R�))�[�mJ�r�䥜-������UܪnU7*�yU���%m�Y�i%�YR���\ԪnV�J{��Y[��2�$ܛ��\���9��ʓrjKjS��%,�}esq:kr�!Ϸ����I�U\ɔu�V2����檪L+�����˕�󒒴���l��O��"��>�����Q9�;���mU�q:���I߳��E��;�8LG�'K,��"wghN��z:q9��LY�,�;El*�N��\���w�8x8^�a+���G�p�����F�����Z����������H��U1�y����W�܅���z_�ӈ���{��槥򫫛Rs�:�b|]7���t�m]����O��o�O��OJuW��~�_t��<����+�ߗ2���%P���e��y���K����>�o}�I�:�{��g�����"�����=����Dn���Ĭ�߯Ӝ}��T���i���}�t��ɍ.km(���^��|5M�)ȭߗ��>�!�Ũ�q���\Z�G��{9���9f)[���^N����_ON�v��w�3�Ԓ�:s�L����Ny�7`/����8��l}��}�}�8��ݝ���\����{{���澙(������.�������L�k�c���9�s��o������껾Ԑ��>�g�����s����1��'�aΤ���w���5ut~���Ko5n�^H�s�ËWx��E�dG���Py�>�i%⧮�~Ϫv�k��jNm�1�����������v�T��?-�e}��./{s���o�\�'׼޻��o5����FG�|���&�.��_zz�W�!��W��3�/\��b�������J���5��8��[9�8��~�sˢR�]Xĭ���[��S���y{�.w���8ԕ�Xߵ�/Nռ�`�8��M��_���E侱o7��r>�}e��������ґ�*�����}��jxs{=yw����{��:�>�}��zC��^�8?��N�Ƽ���T|o�ݥ�\��w��������#��s�z�;9��w���ȯ�"��_�+Hu/\���8��[��!,b��Ȣ���$�%|�&��8��;yf��~�W5EϩW�RRG�M�ߟ4�nsi�h��li�.#��|��h��p⭢�z��.��j����_���V+�w\��7��=��K��[ē��.k�y��{����Vj��⯗���s��GK�˭F��[6�����!�x�EǩK�q��qT�e�H�5��M4�l*h��m�}��mYh��[�؟�H�����隐��#���sT��p_x�b�/t}d����%�!oP���1%-e\�Ww�Z%���+����J��OŻ�U�2-�����w�s����s��^5lͯ~E���ʒ��:LqWR����r����Ko���<o��9I�볔j#�r��>H|�~e',t_i;��95oQj�Y���gz�^!vg��~>�*�V��USD{�~[�}/e�%+l_GX��hω;�y�j7�X�$�E�K����񬦛�'��DRI��Ew�ayN~�������Q����V�R9^�s7K���Ǧ��l{�>Q��}F��9��5�R���?sfÊ�<��4��"��M~E��ڒdKa9��1��hך��U�?�N�u�b��(��6)�NU�����ҝ��ے<��i��7�|֫Dlic�����\e�ko$d_�2v���/��������[��П3��۟�#�V��J�~c���w�:��6�}���F��>ޯ�r������������;z!{�]�O�����5�Y�!Ϻ?��Tn�c ��\�:��7���5�e>����g�ޡ��}�� w��w�3�G>Yɍ8��>p�3�Ws|�+�g)j9�9�2=7Yx��ś��lG>d �J�Jkӱ�'�;��7�w�=�h�G�?3�*�5p�g>�����7{��>GWG�*��=�:�6��S��Њ-c����4W��
�SZ,c��J�l�n|Ơ�9�����s�nc��Qu��]y(��8� �g`��������9�������[����I�b���#����h˝�66G��2
ieܴSF�[*�-�P�8I	nJ/��s.^��s���L\�������{���Q��>>Y䅨jY?"��W�X���UNL���!`���ҝ��)|��r�m���~o�y��$��^���x�i���>�!���d��>
��q��)�א;Nw�Y�};��y����O��p&~g%;P���e������	��p��I�����Z��/�v��M�l��RU�ɣHuC��AFV��CvM��=��F�b���s�2�!ӈ�E�5�k>���9r����Ջ����N� A|��<'���h1^��N&s�z�9�o9�n�J�m��E�/t�m����=�w�{�v�<_n>����x�ԯ��M��Lޖ��s��qwo'�'���gw>����t:+�F��LeDk;��r��K�p|�X�{s���	w>�bB��,�߇`����"rg��H$�s�>�iϠ��}���Gx��WMM)(�!{�=�ut���t����j'xo����xj�N�}J�j7�,5��>ᵜ�������Opr��r�pܺmrY�oaϼr���6��������nm�����4%��-x���4�3�A3�~EIB���Q�IQ��!���hË/xG�;�~����|LӰd�Ũ\g>�oIۯ!�RhI������%qK�o�/ݚ�?�O1܆����m+Һn��i��g�3����0Q���𾧯��na��j�R���j�	Օgt�p6ߴ�g����A>�9�{ӽc,��*#Ӊ���ߴ~��:��"����$�eﳺj��ӊ����i�C�9�T6��9�����W��GFNS|�S�����G^�=�,l�Y��Z���7h���)��-��5s��잜��:/>N?oK�_-ޡ�Ts�Ž�~��~�����*�'�-�����9}�_���}]�Y���9�������9�Ͽ��D�����6���$&}�>?�N)���>��>�����?��7�N?���e�Nɺ��&������5$���I�������yf������>�e>�^�w��d��޾���rg[���}/��ٕ}�G�,�M?�/;ӟuz��#^^\�G��W'7}M�S��$W�"IF�Y�5n��8�\��T��_v>oy�������Q�W�`�Mb�4w� A�K���Y�*�_j���띹��n�y�����ǐ泳�Ր�Ş�9��Ի��no��ξϻ���XĻ��V.Y����iĸܓf����c����g^�ݨ���{j��<�t�ą�1.���.�&�Gk/Z�y�po�G���J�{ɑw�bBK�y$�:�����篖�7�כ�i�t�\^��K�iY�s��[�!CO}���zo�^{�54�Đ�F�_9�y��\��1�;I߽*�uʷ�7���4ܿ-{���0i�>��Ic�A���w��M=?�_����	H��XX���el�D�ܛ;�\I���5����YSdr$�Y*b�(�S�jֳ["h�+#���-�Fڍ��Ֆ�$!�nV\yIr�V���lZm��hMʲ���ȩb�T,DIF	2e�u�ŉ��<����']%bU�+�X�5��m�dKrH��˖W	�	B�J�䊌���Q⨭��(���D��jԅ۶�jR��/�9�czKe��T.�E�n�$E����T��Q��EQ��۫JK�VT�X������Er~e�vJA�(� �vI&�"�����*P"��b�i"�ls��Q�C[)HݬVX[B5��-v�m�#��׭���������e���X���[�%G�吪�9�M�*V�*vIPLvj��Zբ��;S��M�Q��kձ����&+���dI�\�5��)
��8��&�.ѿ�(�c؋`�U%��,V�LJYJY"M%��5���T�k�;�k����j�ULh�IUJ(��i�+"M{e5Ě��h�R&�%Uֈ"����݌���U�UT���uKv1�
%���F'`����C;�8�4�8A�p���&(�B�I+�6�/ҡ쭥XБ(��o��Uǣ�s�����Sֈ�B"�'��(�:��_&�IwFN8��QER���N�w��&���'.��-��A��^�K�[�&0��L�B��2����ԇs3$-"�{3Ď]���)�d�Gk�b�V��*���:X��C�ǆ��v1�욊턔�-�;��)2WU`�""�V�Ԣ��n���
�߷x�9KkeQ����nH�q(���D�i�&�P����d#T|�u1D�T�Uʫq�R[cv���A�9<����%�l�=#z=P��(2ʢ+��d���wI���V���b�Ĕ-��ŏ�Q-C�l�J�ĳ�Z��Z��ƂG"U���
�R��%q��j�
Mym:\���9��:�q��8�Qnˍ]P���k�Z;G��RQ4���jV4�c�y�����Ƶ�h�y�_� �O�O���Y��� |=���=�>;A��?<TB�G��0��W��?������G�O�dR@~ح@*�*|��?��?��QUUQUU�*��iUmWjҪ�UҊ�UҪ�ZUW��U^+J��b���U�]��Ux�UWZUW��UU�*��<WJ�*��*��*���vT)$ڌ�����ugI��m�����9e�X9�V6�jQ���5�UŊ���UWUUQU^+�Wj�����UmWj�j��Ҷ��U�]��Ux���ZUv�ڮ�W��U8�UUEUUV�U괪�V*���ZUŝUU��}�����}>�a-�$�$
fڰV|I�I����|�v��*�U�]*��Uz�UUb��V�Uz����Uz����U�V�Ү�*��UW��UګjӭR����J��Uګj��[UҪ�WJ��]*��#ʠ$��RE	�FC�J�<@����{��Ux��V�v��U���^/*��*��*��*��*��*��*��t��U��UEb��V�u�iUt��U[Uڪ�WJ��ZUU�Ҫ�V�U�)����+7�7-��͹3u`g,��VlQF��V(��ۖ�)�Z�6+7�R�")"�%�~?3����TU�A�`_�����w�j���
a�C�}��a�FΟ�t�#b`��&	�`�""aӂYD�b"tDM ��B&	L8Ȗ&�؛4!�"A�DL�"%�b"`�&�4lKblM�BQ��$�6$ �5""l�,N	���Pt�DD����� ��"%��0D�:X�l(AA ��4hDؚ��|n���@��{���2�)���Iw2Jr����ڰ��_�ÅPPlb#ܣV��B��)GF�"Q+�Yd��	��(�b$6��J��5�FGD��@�U%NRR֧��jX�D��M�	���*��V�$J�ے<jy�!ݮ
�ѐh��A�4GjJ�s�TRXZif��dN1Z(5%Q�<���#�j��u!��\X����Lm�D".�De��A�)�Ҏ4V\A$1ڛ%�i4Ib+Ѕ�vw����`�)M��xƭ�l*���Q���d
�7�1��TŔ�(İ���-�B
�&!4i)YD7+T :�tq-�*��U���x̆#���cN;[����R9�����(�Lq9E�mvI���b����)RI� �T�SMX�����vT��H��LQ2�:"�U%r�F�#��E��&ڬv;D��D�qWjm(��A�GS)b�Dz�ɤE 2$�6�T�U���^2�*��u6�'�-��R�yJ�A�X�Օ��(D'��ʄ*2I}�h��R�s����U[�������������{�*�����������{����V���}����{����(��wwk������i��q��Z��μ�Νum����G��<��I$�Oӈ��;Wl���Gx�D�V�����H�|p9ȋ���3+l�dO�-ȓU��mb$�"�ii�:��C��}q�Q�U��I%:w������������O�l1�P��3���S�������0�F�ǌ���3٦1�yKY�w8^5!���^UQ8p���FFUT[�;��4��-�B3���%ܓ��r��H�/�(�s+��BH�Q��R�e�����K����II&�(١�N92A��<~��Ν�p�0L�`a�:p�͚Nz7������D�K��S�~+���T<>+8��HA�C~h�a��C�,HbT�牳Mx<������B4�\�#����}R�x����Ņ=�#��A���)�cPBF��"Bp�9�Z�Ν8`5�[�`�H�U��u*�&�Uz׌�:Wպڸ��EH�G�8���&	�00�8h���WZ]&*H�&�d�ϴ��I$�$$�.�IE��5�Y�Ԓ�L@�Λ�٧�4�w$��I5%h�:ˈ�c�^��	9��I�%��*Wp�����D9L+c^�1e���	ےH�b�G2��d������I�HD��J�ET��Ә.�p��gڑ�$��4�Jx�x���:&C��[�l�$�7�/�I$��I�gVw�R¤~�̚�!7ƙ�~��1E�r�&�� eyk�⎻P���UD-3L�!q�{nHrJ�0�luS��zn�۸8`�d��8�0b-�HL��(xdz������(���D�D�dtaf�4z�+�+<�'�	���a�4�LԲ]#�4U6Ҕ�I�����l7���pm�n�2�W��"[�e����k��e�DZt��R�X�Q��71���Ra�W_+���-�r�X�$r�Q"�Բ��EE���"���V7Z�����H��'yĕ[�紣��ΕN:�IH�L�^�i�CFp���p3DBC�!CӃf:v�ܓ5[��yY�i��l0����u��e�;/�p�s~�"D�+T�2T�aQ����{��2��z"����6D��E6ֈ(�[),J�!9��$2��e]���)�II%*����[i��O&	�00�8hǡU(%d$�*����U[�����j�oYx�8�ZWoRI�GU���xk�����3$s2�J��W�|�����9\�I��P!u�J툇y�B��&B�b���m&\����l��GQ[p]o�q���W��+4�r�N�$HJVs*��0�o�ޭ�y�\0�0L�`a�:p�5�jNkD�z-��j)j���I%��C)�i�̚lh�ե��x��X㻎N�:�h�`Qa
}�)Mz�D�+��M,�dP�6DFT�f~?���h��[Q#*�;�2��8qݵچ�br!*�Sι�rtll�s�XvNJ��1+��N	��^xzl���&	�tL0�N&˓$<�F��r�$�-�T��I#
�"�tX�r�δ��*)+�1�`�E)*ē�KH�����;�gs���bI9�T�D�'X(گpf�q�c3|e�/�H¹[mXeY"�vȈ��|ҵ�kb�CC�bJ�F�{ĚK��{!Ǚim���[�:�:u�q�Y�+�<�1I�J�(�ʚU=���ٌ�c**BP��(JH1��DA1�e��BI�CQ&�2���B[v��Z�[R+���"V'bQ&WZ�"(�nI���Id�j�Ԣ&�#����J����,4�e3��9�sv�rZ�����ZIC�1�H���ҴU����+X}Xf������}[U�]���f�~�!�S�
J���)��,F~Ő����s2?8�u��xk%BD���1�s�M�6lɳ�:�8�]Ge���)*��JFU2�K�\�Ih�h����Ӡ{8�[HAE,�/�&p������̨�F�;��xɦi�,:>T̈́�3����6��Ɣ���#�i�v��ς嬕��(�UbŒA7STr'��*�HX��_��}V6VC+��S����]�pt^��$�VW{��E[�����IU�w52?	��;bS�d�!�IN��|ͱh�,��L?-��~O%����i尴���u8���ZZ[,Z�:lzN���=:0��+�=!gG��ZZ.M�ii����ZqlR�rtp���L%��0��:N�ۑ����8'I�t�zlRt'IӣgG��:N�g��vu��H��4N�d�ș:��#rtK'KdI�'K�sK�W�%�$�I�q�Oj�ah��F�iV�C�4���0�&I�^3��c�t�'d���N�ӣ�����N�����d�='I��:xɳ��V�\�u�v�S�^���)<'�^V��|!'H||:!�>�'�0�Oj�su>�J��qu�י����5�e��w_Z��|�޳=�BxfX�m�<����N�y�o�kt�ۻ=�7Z�%G��ȉ�9U�7��fsy���k�s*�nm�������t����Ӭu�����f����(<�G�������@Y�����QU���_���|����g����{��ޟ|�W��{��xUw��j���z{޿{������{����|YӇN�:p���	�tO"CF6o�Y'5*��Q	[*%RT����"�*U%@���+q��m��:���+%`�j-9'�`�2:�\x��d0C�7a!	ALL]s%� �"��b��A�Gj")�:����~��2�[ji@�S`��ۑ�&�dȷ�6	C�%*B+a�ѐ�ʅz�4�Fg�P�d�B�J��J�=��j��'�#hx��)��B���Љ�[�ύ�;(@�TiPDa^TiP�����GQ�����X���5�*�U�a�2�ZB�_S���m���~q�mՖ���.>]N7HY�K/zUUQ(�R�(��>dēW�Jb"TrT9�G%U9T�b��A�>��Ĭ%�L���Y.AU�Y
L����
���P�yZm�����?G1�#����xa�#BHI*a�c*)�>�^�T�jS?��b�ԧa� ,`�Q%ܴ���
���G銪��2��T¢ҕX%<B��J��.N0J�i;��7�q>��4e3D���F3��b� e�h���lb��n����H����m��'<`�'D���4t�P��������E��H��I(�,WYwf��f�DrJ��n,��su�"r��N��4Z\eǉ�\�9���sF^ԟs�Ώ�z�z��$p�Ʈ&��beB�ͩ��hqJKD4Mav��^y�UU�$��p@�
A��Hdv��jTL�s̩�:D�!��<�v1NG�1�Cȟ>�M�VP�uH�i���)��Ն+��q
D~�bh"��ܔ�A�]��zi���7c��:�l��VB��;b`�ՙ��Ÿ@<��
�!�H�V���C��;U*�n�1���=n��!�H�v�SN-1H<T��Tq�P����t�!�C�>�
�*�0S��V�[��~8xO�	�tL<%h�W	z��,�EUUD
�*|�q��ẅ4��H���j��%?uYUb���ی!YQ��+�e��`���C�l�"��3R��U"�5)�0�u+�@���x�Y��w�UQa��Y	*�:a�RT�AԧC !CD
�@����I�˻�샌��Cq�;�e�9��/C�n횩MF[e�V�Ԫ�B �hYp@JA��n6�����润􏰛<��5�>T+U�p��%A5�}�32�+��9|�|ڸ>aU�*��y�'��"'D���Q���3�ʄ���t�ʕ.��7��UUJ�h���v`���44%���r��1��Z���3�a��!\������G-�;�sox�U�������//��Q�-J�³�&*�;�*��	U�b���7���uu����ƈJf��N,Fn#�n3���#����AI�С�0�9*Q��'��a�R*J�*�w=�9��$���J�����0z��6Z`l�K.Pl!^"�תc.���*�֦�oI�˕+*�f>%+��8Jn>�ȧ��,%:��~i����6�����<������g����6M�u�Z��'vN<UUQh� �%��JT-���'$�t���K�h#��.0�IY(}2@�{X)$����~��-#[�B-��)��жW�Se��faq�32H���<��Qu�U�ъ���b�ba�9�j��Tk�I���*����q]%9P��S	U]FZ��$�AQ>+�¥a�D��R*>V!��J{Ҥ`5Y
<�p���#ౖ�F�?*U��.SJ���U�v�£(#LD1`��=�&���!8mV�*ەj�]��R�TU3�1�0�b����������Ϗ��?�Ҕ����M�V«n2�F��V�Ɲ�M��P��k=rFi���<C�P���ѼᤤdB�����;�]�H�ʙTl��5j�[,c��G)ȅ�wfY�b��4���9�S�w�u��]ePF��ћ�V���R���r���3�F �<���л��-j��d��-�aL! ��ZH�@K�!���h2���(�2��ekL!&�̘�!KTp�Ua���S(��6�Z��%5Q�'w>5�Պz����dz<�Z�UҠ�6î0�f�j�L׳&Ta\���1�u�?��X��1E�}��f?�¡��CM�Ѻs��bu�Zn'�:f�ǌM	�|��#�y��������E|�[lS�Y�|B�S�ӌ��Vk������?"'D��a�f�|�p*O2�u�N*���^2�*���C�F=;�������h��łD*/B8�V�;(�gRM���t��c[������*�X���~�V¶p��EP�Lc���=}�4���L`�EF�/�Q)"Y,j-c�ǋw��2w��Ӛ�����aɀǡA�4�aZ!�q0�0��8��
��4J��|��ūJ�T��U����!�����!�G�F6W��U��Xy�[u�����מyǝ������q����P�W�2cU�1�%)�CV���F�8���~Tb�`H5K�A��G Qs�F��_�� ���E8�XC���c��J�Ui:�hiA L?��ϙn8��奡�_^�Ӵ8�Ɗj[ ws�e�n�	�����b �04ѲQ�\�� mˍ�F�}7�N�q'y��H��*�^�B�;�%aʃ�"��}h�Ө��֞�ծ�odEa~mk~q���מyǝ:��g���d>>�&̊1����k�����m��c�FS)��0<��,��W �[��t 1��F���՚F�]TUl�o�~�8�EH$���e����UX|CD'7I\Jb0���9T2���_�I1��OTy��J}T�0J��*�QO��U?#�Ee�!�eX���U�Q�j��I=��b������YW�4��%a+�t��U������ǭ�ƣ/�����(�qd�d��=iK�(
4���kF��Ё}�	E�h��é�J�m?�0��-�4�<�G���2�Z~K~c�[������D���Vͥ�Ţ����n#--0�FVť�bb�ҭ�-�X��gD��~!��ؚ'��0����0���Vͥ��ǖ��m���ZZZelZ[lZش�-.N���6ta�鱬:&���ܝ'Kd��4�J|"C��tHL$%uI�ʞ׋����{O��M��q�+Kb#I�ZWɇ�+�u2�:=:ΏOG��N���I�I�W�lZmlZ[ؒ�䴷�[�6��i�t�)xO5^j����<'�^)=��8�[��x����7Hh�!�G��\���]���\ݒG��i%Q{D����9��*u��3���~&�|w���G_n����ĉ�*�zׇ�&��M(�t�ݖڤUn���c"����.���_;�]lk�"G�+�������{�\����ǆkM���UUCV��b	I&I֬�:��x���2I�
Xe ˏ��6J�%oy"�!X�
4YyG�kI��8@����L����d��t���R�`�<�M�!�\�3����~�N��<f2�Ty�:w�!�{�J"i\2�$�y��z�dؐ�$a�����$4��!�U	�r|��ÄD(�<���j\�kFAf���r�D�����rV�"Bʭ)Rq����g���F�G��o��zh��AQɤ�7�ɖ�:L�.8qf����d6��O��:�:�[1�^�<�SY<�-~N�睾���]��D�c���;s��v����c3<^�YF��\�ʤ��q�ڵ1_*�����!�EZ��(B$Ӫl�R�,�9��(�F� �YY��ѮmdC��vW��vj���D�+��Ol�V�i�آv�\�!&:�E�J��Sjڄ�b][u7��ۼ[�J�N��H�$y�����N�bm�E��&�\�mSqIZ��[�jX�iF�Hbb��U�y��/sb+눛2E� ���0�v��T�^M�����w�{������W��������{=��{׽�~���Uz��{������~��^���{���w{���}d:�n8�Z�y�yӮ��q���}�ҪKs�թu�Kr����шBD�7
R�Ɗ�q��n�o�p�Z%.AA��\�h�2�vdc4�t����H���I�iR͎m��T�� ��e��f5��d/Z!�*��{�n6�yZ�D(�f�
����P��.�
U��C�ã&\���h�׵HUZ�lw���	S8aM/�F[��x`�Q�X��U:�r7�:oY��#|���0�A��e$mrNLV���d�+(�+��>�T�@�E����H�%&/`���`1h<B���2RN\l62�B������W��K�T� ��!��ei6�d��B��,� �J0��Č��5QV����~EyPe��RNU|����������"tL0�O6feT�̪�UR
<*P��`|RPN�T�F�Cf�D(�Me׾���w¦[`i�LJ �H6H�O^���(4�	g��	�K��c���.]��X�b�iL�`�Y���(C��t�D
h���+1QcC�ڑSJ=�o��Ϲ�l�ä�͇���ֱ����ZCWkK��ʳ5����� ���!UAu/���!!+��
�>�P��O��[�-��V�����8t�IUCr�BY	�S[�UU J�[+E%} �D*�/��5���"o�[�M��Uy�v��>���/�ҧ�+E�����648 ���fFQ�զ��/k�� ��f�К4]O*%ݰX����Wao���ȮRS�N`y{ʣp�a���
�F�<h��l08pX�/���|HIƇCq��r7!p�$.Fx�����(��e2�g�Ѐ���3"��� )rp�z��qOL��N��i�`�O8y�ߜ[��y�t���|���d�D�-XsF��UUR�J
m���>t4��A��B_�.{.U�UY���HՋKIdl�&n��+�X��-#>��i�R��.��\�6)�$`A�<쵌��_ui=OW˫d�T���E1ZV�)�r��\h$.c�)�3�IAp�a��z0�#�:��C��۷C֜�L�v塄
���K��ӑ�H�Yйp�������LV�+���o<�?����00�<tٳ'�IP��U-E�5ȷMek��nV���kx�,�WY���2���!.K1�+���H��R���Ɯ��6""��9|W.�Ɏ8�Q���*�jUⲪ�XH����g��UT���\�1J�R�*i9���B�Ԝ�(|x�)��q�чvD�]H�	$l٥�X�	TQ�&_`�Xv�dr:�=������!	`��g�G�!��<X���m��z�C�(j���N �HS5�$b1����jD0��b�%i���pP�е��BU.>0�i�|\���K�qq�mi�4��܉(!��Ǌ\
����e�B絕b�v���"�CJ¢�*2j��YΫQ���䦊$�R�I6�C��l2�ߖ�����y�t���;ܞH@���䕎Y�UT�gAS}�&�7f�i�Ɉ;,�����j���]�0=d.;�sNI!a�x4�5q����%���J6|�+�Wۯ���2sQB�J$$��
�B���_K!Ļ2&<t��,.6��A���>y%�9�C���&4BT�,�E����
�!1��(g�۳hӐ�0l���n�+p�g��,˓O�	G��Y����kd�\iH��h�PiٲMʘ�z�Y����m��֚[�<�疷��������+�Q���vrNX�J��*�{+*�UYIWG�r���D`����L�W���Ć�7Ĵ��g3�:K>���d3s)�q����Τ!����"L|j�U����c
�Õ)]6�q&��Ǣ���^W6�g�Ϊ��<80��kGH]p8�2cM�kN����ޯM�1��XI�'T�0���¹�h����4p��N�8zx�Ν4J��l�,Rk�*lދ�����5��d����YҴq�i]�H�4�����5(�2	�d� ���i�Ɯƞh(�o��x��F#@�Ѹ}��*�!4�!��@�3�ԩg��.S
�^�Lbߕ�r�8Ȍո�����m��������B5	 �L4�����~ϴ��9s:u�^����0�N�Q*�M��\7Z�~un-ǟ��ַ��Q���>F؎FI�*Y*>�YSJ7���!F�1����I<nf�7HK��n q"lw ϙ7Q�"BB��������,�)ɺ��f�jM&K���Q��E�$�ll[-�0`��⪪����W�����p���qN�/.���s�����tYP$~3��4Jѳ~��y_f�@���ڬ�J��4�|�Ɂ�\ә��ۊ�-_+׫��+2����H�a�m�.�{_I%G"G\�)��U�q���:�+KWk�!�2���a㗹I
��#h�Z��c��kfǇ�8t��B��n86ڰun<�����ߞZ���:�8C��u>E��J����iI�-ڪ��>��{������#t�b1�Sh�a�\}/%c�M����HU0�e]V�+��v�Sf�M*՝�#���19�4?~J�;H��u�aF K:~?���f�1g3JWgS�]���!iSm�<v�y�ƛ�`B���7TT�bB��G��0�G��;�0�-J��OQ�+�Hx��O�'��x�[��8�%�KK[[����'I�t��*��,X��O�Z-�-$����kb�7%�V���4N��$��=:8h�}'IԷ�f��m1�YlZZelZ[k_I�zN��tO'Ge�::'M�T��t��'Id�c���)!���}8�JO�-����������-8�BӉi\u���4�N��2z0�|'KgN����<���:h��I�N�Η�t�:='OY�O%���|L6�6��)u%�H�/*��'�˛���I�v�Ht�C�a�:J�:C:F}���g�a~�5��qU�����S�5��z����:$�{'I��yY�F�O?vB���.<���wu��:of�����\]S|��^OM?i�n�c%KWW�*g3��j�<ն��B>�k��ɓ;���5׵̫�᩼�]����eV��y����fOCm�5�o���������{��U�˻�{�{����{�⴯�˻���.�W�ҷ�]߽�{ΕW�ҷ�kZ���q��q�Z��ַ��Hp�d|��k���@�t��24?��z��ҭU�Gc��j����P�$��<�V82�P��C�2�t.y�7 �߽�������� 5#c��%��D���D�g�gs̚��pA����xF)�F3�D�� j��e�dh���6prVIL%H�S��L�
ᩓ�)��W�ȑN2F�n���O��2�ο6��ykYç���,Y�I�c&HZX�e����*�螐�T�HCE|p7��)��Y�b�Xq.i��aO��D�K	��5�+#�#<��!	ʻl������+��t��>
Nס�����%p!��>\8"�U����V�#�DnyZ�;���1���z��'"0�կy"&&G%s���U�e�v�d�l��zUS�!�Dpl]$��=�4d��'_�qן�Z���:�8�-�w�ʓ�	!��j�˪�x��Q-�s.�ik.@P�W�#�*(D!����M��:�N�����aM�]��N��!Dҟ�.INےVHE[���DMG-pP��9R����h�T&4ZTB2�˶���UT���M�{�\˲ZZ׹x^��<dn:�g�d<~���[d����#�=�q*~�%��ސ���|s�ě�ceː'�hrQ�'�l��&�m��V�Yl`#�;�.`1��z����q{��\�̙@���H�#�Ɖ%���KD�E�ʐ�V֭�Q�<i\V�<7��ժ��}�T��ڞa�ַ�~Z�Zֳç���,��c!wF�⪪�.����e3�6 ]�'�FJ�0:aI��pll��$�C���(�c.�q�Kѱ���481qa�tϋ�v��ǕS*(gy��������VT��*X������zn�>�OjW�grg���>ϳ��f�4�2�珛"2��*GϪՊ�o���θ��x���D�4{�W~�jW{\��ܭ��Ē�#\AԿUUT����`���c���x����=vW+�¥u�CX���öD;��q}Ӊ�%r;1r�s�B�h�`�8tB�L�AS �#�h�A�^npz4d4��:.Xpm�Ü�T�l���+��C�OMf�V��O�d�y!�[r��qF_x�	��j��y���I;_�iP�y��TH�q����y�V��ֵ���<��Y��J,�Ze7�r^dy�UV�b{�@����,�A��έ�JnX��Xr��`;�+�X����ǉ��1VZWR�Y"2�����H�T�3_3�e���Ek�499\ؖ<��\B�˖4���9T`��$�|b��e�oң�e\m\�?t t�tm���C pG��8h?)),����u��>DG�2��zz�`�k5���Xy�_���~ukt�������0G�i����nr���7"��`�.ݼw��AL4�D���&��D"�ℎLx�D�3H�D+�	-wSKR�J-�9b�%#�n�؋��
�,���&Q*[K�b��"^~m��@Ě"���ܲ%�%��,�.�Xź���U���}�Q��3��0;4ظC=Ԟ��Wd8<n`3>�*�u���{.:�-�)O}�7Vt�%�0F�z���CP���۹��F���e\��!!��I�>V�фz�)��֑�����#�Hwۺ=%	��ax�F��"5Ug���G8>�@���!
4`�����F�?8��Z�ZַV���8C~�����uo>��O��oE�5����UU���U��+Gƍ��Ie;��v����[6nil���[��,��Rt�E�Mt�]u��V�$��֪���?Vw�N7l8آ���b�!�ĝ���HQu�ہ�?a��˅!�znp�4�pX��6(��v�������Ӈ��4l��<x�!��ګ����$�e���UU��U���ᕮw��9y�小���TT$�:��W�V�����;Y��W��"+��{��R��< ��T����<+m'T��8(ي��u�"!�oM�T�UD�>V�DB"Q�r$�Qz{���#5�a��%a�qV�Qſ�?-o�����Z��]Genr�eR�^�^V���ع7�j$k�U�..�����nO �^�ᆫ<|�#�&�2��-�f�a1\K�9��d-)+�a
:)S�ʲ�܍�s�8g�M4��A�F�Q"2�#�Ef�T����7�&&���D.��>�a��� Wk��I-�^���2�>p!��b�!
�}k�EK]W�.�T*�PH%z��4�_�USh�-4�[�X0��$?	G��C�W����$<A<P�,ׄ�	I0�'�a�6���ش��h�m�-���4Ţ�iih���Z<�F�5�nN��D��D�t���'D�}!�G��<:t�L��tЧG������~>�#�>�����G��[�����h�:):lL'I��,�,i�ysO��_c��sK�'�O"�J����%��V���p�N���e�&ϙ�!��C����_I�t�zt|&N��v�D��:�ܝ'�D��N�	�H������^�x[�S�'��|���Bt���'d�;&���N��:J����:�{��ꐒ
�ng2)�����[�=B!u�[�7�H�"�uT���5��/5o8p�EK��7�u��x�Jpf��]����"�����_�޵��s��G�������99O-�70�'%�e�\tsto�}�:�<qN_?z��WU_/u��o�������r7��>l�\����8Cr�8�p\��6h��A9[D���4J'Gğ���l'#�l� ��?}���j�Q��$5HR����}�9��e���tG�t��]�p���:B&2芕T���V���n���^4q�3������f�Dbmee�&�g���Uo�>��Y=}P�r�'���&i�dCU�d�f��]�h����`�z^M�ɚ<��=�VL�X�F��{��dcz|�È�C����AG
�(�9����^��E@�qTn�G���/$%5�st����ԍ�jӬs�K`^�����A��zR^��\yo�����7��Tj��jѮ���l!~�����wyo�[�%�z|׵������{W�~�|Ve��}ި�vJ����t~�z�ZGD�}'!d���!d�tS�%i����lNږ1�I�Z��-h�G�T�J���L�����`����P�F�A7�׉�Z��^n�ejh�UI;b�D�%vESr�H($$+b�ք�,�U�g]H���!,J��>�Y~\Ubؘ�z�erʞF۸��̚�B�!7!eH��*F&Kd��lQ�PڸɽT�ԣ��5z���z��{���V��ܻ�{���*��oܻ�{���j��J�����{��V�t�~�߽�YӇ�q������]:�8�-}�oҌ���f�-$�j���2�iM���#�%���CЈ&:�s�'!4e��Aqzm&���$,Zꄑ;mR5\H'7ePojr�.u��8CD�%�VC����o��z��s&J%!YaS�&J�mQ���5��q�R|�>���k6-^�
�+�#�`�
<%�a�~BI���6�H����;]u�%��+���<\�X!��՗���U2�7��T]c5�\I%$P�Px�F�C��#����B�م�(�Fh�"���"C�w)�s�R��*l�W��E�τ1������!��9�ȯTE�ӯ:��-張���Q�E����UUZHzT)+��!�ۯ�W�-�N��ū~|���{���m��ժӵ�n$��H��a�ᶬ��D��H����# �pL-������0t���c����8]�"D��%�%��-	T����b�88�rM3�H�I8�R`��Z��Z���7G�[DE{M�����Z��u�k:x�xO�a�k��͕-R䉨*d��UUi!W�]YKJ#R��C�����K�÷2B�u��X�|l��nh���QgYba��pB����-��/*4E*B���3<t�̹ғ�`B�Y���m�I>u-8#tBL�f�W?�f���9�|��Y���E��ǉ8��0�ć�-��ո����[�uӮ��2���a�cׄ-�\b ���6�m�b��Y&XUr˰��Ǻ\Hd���IQ�~�������]o��w���8J⥘�#+�:�-ee�%\�r+�W���B�W�Ҵ:9����DGMZ$ڧ�=�e�v��z�*RTH�W�eHm�}�0���!�7���~3�t:Q0��������$ C�R�C�Q>w$%˜446s���i����V��y張��]:�8�
%�b���Z�bM���k��~��]�7&,�V�H�iq��F�a(Ɔk�Z��B���2�rd2-��gTB���!�2:�1�1��V'mRљ*�$��9r-�^z���C7�ƨ��[�k��&Y�:	8<e�'��:�Q�^�d,clB�9H�����R�6VSڪ�#����|���W��q�6�m���7>^��<!ط����uYTYH��٢�|v������KQ	���L�4E���y�m���*li2����)�B<g�?@B%k�xoԚ��¼:l��m�8������t��L���N�M�wE��zW<�m�������(7�"GӘy�/L�#�a�g�R�f"~F4m�v��h�h�<zX�\�B�7CT\,:|CDD����	�D4���ڷ1f!�X�L�A�'ǽ���6�*�E�u\��E~x���X���z�Xe�Շ��Ҿ0��>�I�_�V�v�N����?8���Z������:p��ĳ�����z��M��ˌ4yꪫI*�l�$���xz鹒��$��QM���<�K!���a_����RY^���¦e��Zd����$���%�*Q�H@d2�֕�WEH���4�W�!H��g�g��z�J!��%��c�8x�pw{�J�rp���yʎ+�Q�gU�I�㌣u�YF�?����g�u�f�ڲ��D��s1�4��R�����-弳�������,�IZ�UV�jO�,�U�^�+��a�~��#�j��i󇑻�V��{��O������EFE������R<�x���|0��f:�*i�ȑ*DiٜBr,"�v
[�l��,�i���rx��d4C-�7KѶ���� ~ϳE��;RĎ�?�p�Pn�FII�m��6.l�g�6'���0�!ӆ��S9]ߥ}u��8���6V���n��8�օl��h��lf��i�U�Cu��g�Q���=�jO�J*�eye��QȤm'D$���m$0�ul4�UU��d6��,Iq�%��şr�xU�&xՠ���k��tI&1�m�&��Q�%��#�>~�*F>w\b�"�(��yˇ��\xa0Cw�w���.Me|l.B�q�d��Z̡� ���_s��!��T8:" jdN���) ����Ѝ�&4��h��D#8���o>�t��ݮÇ���������Z�Z�u�]GXq�Zfe��K�e���1��UV���Ҷ�~�v�[k.��禘a��SqD.r2K1������y�--j��h��IRk=��n��Df��b��l��XVB�����j��������"Q��qĥ���{�.�.�lc�f��l����|��'[��h�I�d<�3@�_Y4B�z2�!u�_}+�},؝0O��0L�0L0�ç6!B"hDN$D�H"hK�DÂ,�X��4&�١4A���	�B�DM����8�blM�ͤٱ6%	D��x�ȇ�yku��[�-Ŷ��GϞel<uխ��kq�4 �D؈�(D�8X�l�A�Q�2&�Л?���&g{%���+���y{�8}�-�S^;*uv�η�u}�u;z��[��䬷sU���q�쒷Z�ݎ�D������8�������j���.��^q�������U�Fm��Է��V5�o޿��7��ퟝ��?sg�ƻ�]�ֵ�͘Wܖq����IK��}�g�Z���ܻ���{��[U��߮��{����ڮ���w�{���ڮ�t�w�{קm�mŭo-o8뮣�8����a%H�UU��j�*JJ�#��|�9�Oʎ�7]��a����ZLQ���1��+���G���h��F3;�ӂ>;���װF�22e�Ր�[�7���b4�U�nT��[�^j��y���on�xazK�#���@��{�4l���u�yj����iVW�[����O�x�0�aGN3�$�Ѣ�r�1ޓz��UU���5�|c�ɠ��N`�ilܒ���՜(���h���W�:V�cR�b���1�ge2�#�M��n����U������A�¼t�,ɒV���D�*Vnܙ(o��.B|��G�ʌ�X�rv�'!�*�����������|�W쥗�0ش0BS�0��y�����N<x��e�<��ۮ����l�%c��[��k�4�ɖ[�2JHJ�@�<`�������5QU��(��,�"T����حaf����L�Z�vd���*�KSF3ŸƢB3&)��*� ږNz���CT椲&��-�S%�q�f2�$U��*j�6{�Z�M��_��ߑ�A�D�W�@�0�C�c��X��<Ԭ�3�N��p�U���$��{w�2�kW M����L�g93/�FM�01�bc�8��0�%ܐ���|n�i�E!f����u�D�0f�ڤ�-��$�X�`}ݍ<Ć�%N��m)8�͂0�LXi����uk~yky�]ua��9O��\��I2,!y<��UV�2x���.��Rs���!	8QQ�wcА���m��.C��\��?}}d��J)#�I6�!nf�l�X��d�^s$��� ��b�<%��[������HC��'�U4O:��qە(�>J��!#�����D}\���T�%F���GH��p�brXj�������0�&�|�����~yky�]ua�e���dI�.�0�%�[⪫I+F�T7��C�6i�Q�+U��l�ꆡ��$?Lu��U����hS<g��������H#u.��G���d&B2Ll���n+p.zs������B��ު"����h����>�ʍ���Q�m�!!D.��$$4`b��9��_+�"鈕��<~e��i��[�yky�]ua��[rC��ɑ��z���@.��}�J�		��Ǎ6��́�GD~��'$����"��ő5QHbc4ϙ���2h�i�	���,�?f�j^�~2�?��.�0�oC�Y�Q���'մw5�,#�����ڱ��I�TZ�a�Y�V0�~=8�%F�ex���	{�!!� ��T�ҴV�Vi�u����qտ<��Ӯ���ӄ0Y�4��k;��u��6d��\�u&B=(�H�2)���-�J�sy7�����R]��z�H�!�&&Q�b���{Ϋ��}:W�A"�m�#��R���	�\U��c��2҈Yq��5y��m��x��)��JJ�$F��!\"�n�R�F�K��g��i�	46(�����!�����(�I^6=�D!�K�X�0C���M9t�����Ś^�:r�b�3N����!E�G�=R�\�,@�f��D$�.#Ɗ�UuX���K|n�G��X-��WR�����*ʘ�v�hK��$v�ӂ�Q�nܒn�;L+����z�T�+J�yY|�kx�p��<&0�Qӆ�g ׵��Y�nW�������@ke^�4`لtcrD#��W�1�W����àz\���S�;��1��%�`x>�BBS�����c��I�rH�˄iW+��M��QБ�<M:Pi������	Hp2��W��O>+)�p�^��3_#�czb����u�e�T�}_W�F���?4��ͺ��疷�4��ӄ8��:�!\�ow���i!�]d5��PV��]��+�{���x	$��BX<O��a%�T+`�:a���A�c?1��؛���	A�c��91�]�Ơ�#QE*Y�
0��d���)��r.�{�x���,���[W�#��""1Jڴ�>>�iW���0��ݮ�1�NW�F���k�Ȏ☫�8ێ>yoͭ���<xL,�aGN5֥rUOJ�zc(.- �%F&as�UV���<�4x�Udt�E�\h�w��sDpK��DB�����{u8��l��A��F������nB�8����8$$�)C,c�G�n�
9�r��.B�r�<	Z+N�!a¡P�+�Zk{F�ñ��tl|X.h�gm��'��%���ێ���Zq��8����`�&	�`�&�Dât��H"&��'M"AB&�L
6&�؛4&� ����'MlD�"l��&��,KblM�6%�&��rO�B����M��-m���>[(���^Ǐ�x<x��M���4&��w��,�B � �"Q@�&�؛I�����o��nlϤ%s�Wb��8\����ǧ�s�E�|��98/{���✤|���h���$&�v]�\:ɞC�/.ꤺ�����G7�Ӟ����$�8Z�9��c���!�?W��:��Vے�_7�x��̶rڞ�=��|$��ECMD?Sbh�6�D#��Y��O>���ѷ�|���؏ۼksc�BR�I.\ۿ��4活9��dɖ��X�}K�\�|5����e6��q��|���1��BƗD�Mp�5h��8�bĴޓ������sM.i�td�cz:Hj�}�8� ����b.��Gv����街j%���4�rhq1�f��o��	��Vl�Ո����>y���~�>Drx��-��#q��м�����p�!x�)d�L������f��H�����	s,��[�.��ͷ�/���y��m;.����2��fk��;���=�M�7������4���BY2},VJ�TW*��^ET�AF1�YT����2�n6��b�F���
���=z��6��u�(�%N'���?n��ks�H�i����<��m:�&�tD�'k��]V�'j��R�������tl����gV�e��E�NJ��t�kB��:��+$I�2քrMX����|��Sۖh����g��"I��(�rEc��sSYy}qګ���r��{���Uګ�����{����Uګ�����{����Uګ�����{vt�ÇN�<x��<x���Μ&~�6���x�Z��\F$��G�H�EeF]UBK��TlEP�R��ˉG����.+�iQZ�E�-(�D9�M�7Bnj���J�m�'+jA��#J(��6FTĪ!(�IK���k9⪫CXn�\k%�;�ġ���i�#3�gƚ�1O�\G$�2��V+&[�s���Ɋ�^Y��gW�$TVH���Ej�<+�%��/��Z���J�Y#�BJ�2�$qg�����6uAa#To.:�������,s�?)ϿNgC331ʕU�0���V�$������N�#�:p�*B?l�~�W�Au��kCF���VaR�=̦P�%����ÆUr�Uܫa&2ڑu��p��j�a��f�m]Ta����2�<u|�M���A^w��DE�bq��cQfE �&A7�0�3��U��t�㿪tm\r�E~R�Ɇj�����*LՈ�Ų��mkqםZ��ua��vݓ�V� Z��<��UV�J��e`nH����N�0m!�����p0(��x[��*�#L�C�h4
,`���ƛ��0�G����++CHX�'}+A����;D�h��ca�!Eܔ]x�G�kEm�D��|:gL�i�t�Ys�u�0�.]8�έn��έg��<xG�t��ID��`�n��d���R;UUhL9�HBLJ�*Z���Q�X�����q�E�}ݯ�$2�%�vJ����q���VW%l8n�����۔�%IRn��~V�3j˹eV�`�#��2����$�iP��k ���ҁ�����S����(B��K%�VJ�&̭���zo*�Q�~J��Ti�y��~u��t����N�S'�֛mTD��\���ˬҌd��l2a�ZA��+*��CC�&��٬��B,�Չl��
"�7,1�RM��v����da�m�V[er�.U)-���
���m��x1���e�%B�(�0�s��d�"z&��a�{�KSo*�e�Q�NE��H���j��x��i\Vh���^�ëV�k�ē�>y{�[�̑��Ϡ융U��[,l������T����[U�o��؟!�.��I�q*&0�*"i�n���q�yky�]ua��e���@�zUUhO�5�nh�(�V���	W[;~�N��sE$\����V�hh�_rN�x���$h"3�Ʀ̗&B�=�ci�B��-ʙ\i.c�69�~�����i�th(�!8%Xl�]XB�'�Q>U���RJ}�\e��:��μ���e�P�N=�Nȫ��	d��=UUhe�g(i�Eqe˙�|$�Of͂�L�$;����a23(1���="��ɍ����85+ �x�G�@O�J�IR[f��j�y]��Ѳ?��~�a�jQ�֓i���[��9Ta��b�1,�]"ބA8��v��8��^m���-o8ˮ��8�s��K2��o�UV������< ܃r�t�ƃ��Rt氚��bJ��q,m21f90��� �)�I�:e�]�B�_b�Q�$�%a��|Tkg�Ia���Z>'�`��JQ��7�ʪ�EKcrH�o�%����i������u��2��#jI�,z~�x?)��77Z2�ϟ�[�?<��[�2��Μ�0���(��em�q7u��Uy�q1k)������A9����򆚢�D��A�cA��.��"�8��$\"�﹪����6�M����B��HV���nVHe��Rfe�U����Й*�9$Pxș8�n�8L�Q ��Q�x��s>5�t)�ĭ|c�Wj�i=u2�ʐwF��"$e�$&)]��J���`�U��{�E�x}���q����X{^s�ߕ��fYu�yYV�k�W��$��	��l�	�֐���akknˑ-�+t�w��.��V��O���\��&%"�~mźӏθ��?-�u�u�o�Fq�0���.F�M늪�	�@��>�Ɂ�g��Ltw��&��W�?vc$L`��n�uĮ�������9����<�d,���I��8�^+���ծ�!�0��J��j���|,���A�'p˾ܪ����L���x9! esg��C���!{Ҽ���*�xÆ��L??&��`�&	�"&:'N"C�&�DN��!�D�4"X����8&�؛:lК �D؈��҄ �,Љ��N	blM�d�JGDᲇ���p�	�"%	���tM�<p�e�xa���DD�:P��!�Ǎ�<x���	�0�e�f�AA�L�e�b#�SwT��p���{�K�V��<U�n��=Ûx��g(߽mm�w�f�sECP������q޲c\Ԭ.���l��&����>���O��4�l���;�=ɮ}���V�,�;;��Z���;y�=�{�,�_>w�8}�-v��ۼW�����iU�ww����{���t��ww~���{�����V�������{��եU������pçN�a㧄�<xN�<<!��1Ҫ�F�ee]N��+e�u��;�����h������Gɓ���d�s���9a�#�,k�E���!	Ƃ9�LM1�G$Ș��`⒊��vZ��h͎��h:7��ͩ��<9,h=�q�_V�2{u$Gw�!���G:�����1���b�����W�v��ԕo:l���O�`��	�FC
�8rx�"�Ė�۞��۞o�UV�M\�XT0=)+��o��6s����B��pZ%'B��K���p(�RF1#7�IWC�u��i?T�!�H�w ;�\r8�sc���2`����+�t�+�I����҈HI	ik��e��Ǟv������|iOw��n�m��Z�xN���?��0��p��N��f!�(�?�![I�jPmTǈ�����Sy
E�)X��8-V��D�J&;u�r搤���i&�b�*�>��[�KQR���dJ�<]Z��)�$��8h���+x�f��x\ÏUUZ3sp���G��r���c�DTƃ���ߪ�ӻSJ��ſ�1QY��1��4r8tT-A!6q���������pr�.�f
�W
v�.4�����٠lr���Th�HH�!��ﾮ�.s9J��uWZ��.���a�]WT�u^?"a+RC/����]qo:����:�g<!�{�����[�j�r	a�:��Ѳ��W�= ����+��z]$�~~l��WW^��h�_��U��[�#��&���dHpo���!�S�Y�AM���GIcU��yJ�j��y"�����p�KL�86��SUQ29b]����=�V���9�I+�:���\'DL��:h�a]'
�}����ܒ���ef��UV�:J��������P�!�L!s�t%ۖ�����D�s*n�Q/�tM�V.r���G��$���~�E.��]��2��,�2@�M�n�WXu����+7̦Yffc8�V����Z�U�^3�Ն����Rw����]=k_jI#��>:p�a��`�<'Ma+���U�냉��ߊ���.�,��zgH�UFC#�
�g�!�K���fʠ)��UIG�����~I��x;�g�M��(x>h/��<�v��Fy]>�qX����\>�
���I���u����"LF&0�6�:j��L��}Ky����?<��[�2x���������Y��|�1	���X�`���-����k,�����-uW		(�a ^R(S���8%6m�C��g	���!(��q���]����N���(���!(��Z�6l57�m����C� �c��5,��U%�(q�l�x��t�{��d¾��X�ݞ3��]7ӳ����LV���>�~W�"}EH|z��5��s�.�|�#�iu����`k0:w��V�"��d��,h��d��[R$�$$�����=%t�TѪ��KT���5ZW�:xi�4p�p���0D�'J0�WI�{'���&c~*��s�+����N�F�Q[�7{aՃ�},;��+{4�8�>D���$��}��x�2�է8���hclN,=�C,�I��h�C{߲�a�@a��k��5rF�^mÎǲ���;$۷Y6;�orf��o��X����:"`�����a]'�+�ujݼP�N:��j%K����m��r�%�c�ɍ/�*<�p�g�x��Q�8Wk*�v�W>����Ο��*\q�VۭZR,�%�<3u�p6͇���Weevt�;IHO���r����[�{.�ѹ"5�D���Ք:�5&��;�!�Џ,1��9�c%J�<�q��<��u�~quc���q?�8>"D�Cu̒9��L2�����jC�k�mՋq�Eh h���!%�:IyA!q�wHFJ�h�t=���K�K���>��^\���Z���V4��KI�taƂ��Ҫŗ�I���L�q�VA�=�mkf�8��kDlo?T��J��O�X���G�u+Dj��I�W?+U���_�'O�O�	�"`�&	�`���D�e(�b"""t�(�$4"%�'DDN��6&%�6h�H"&�DD�:P�$b$�&	�p��؛4"l�4%�i��>A5��Bp؉�GO6x��x�""`�(A��<x��x��ǎ�(�Ś(AADJF�M�f��z�*��w��Ȏm,��9�^�v��%|�G�j��9j*�T��L5���<�PR1[�ӕ�v!*�ݧ.�5"2۰�!������ӽ��!����g�u��w��7���]ۣ����Z9�g�ӨzpKU�vF!$&�wl=mZ�$��XG^	��p����օS�2D�ń"h�V�T��%��e�{z���Ka�E	)1n�>E�A}�:i��Qy�!vm(���8�k4�L�c����ۗ	��� �e�4�\6}�"B��tAs�����H*[�^XB.M�<ÂZsZ��8�¢�9sd7B��x��k���ǧ���?oP�t��A�֭ݻ9f4�+�\P5I�Z~�f�a�]{㆚Kk�ji��J\n6!T�_�f��y���v^�.�������	y��o�ۋ~⾣�N?s��7�����Sn��S湯J�&V�h�!"�Yj�j6�UWD��D�T�,Dd�S�88�k5������]_75<�Z]�N�T�%e[Q�&�l�&���A��1*�-��&����"X�����i&8�`����:���ZpD�;���s^�c��
�AB���;G�۴�{��m�IdHUM�� ��g��ߩUn����{����=ZU[�������{��V�V������{����V������:t�O<&�~:#Ǆx�����I������ёrj(T�#b��2�:$*'2���!�6ܴ�����n92��7Vm�t��+U��ˑWb�18�M�V���1Z��9vsx*�7=�UUh�j���ڲ]B!�B��n�B���]�C�%��d��Ӧ�6����*�Y�ׁ�W������M�>a^/g�˕�&�[�aZ6�NE�\,��8��s�J��Ẅ�,�j�e=�g����sf8ڶBX$��'��Yx�W�����OJ��^/�=${�ɺ�����&4'�<'O<��:��:�:�-��ꧡ��w5�g�E�y��#��b��n�7�m�"GOx��e����{2L0хr���Z>�@���%"*Z�0w�<�ll5a�v��%�/EE�&R�`V���e�!;!U�4�́�� �ͅ���t�̹�4�Ӱ��ϘK�𿝴����~y��yמun#���=�����$��C��DD�����������¥k�&$��l�l.I{���Q���ӱ�Ҏ>%F1��$&��U!�2����v6��;t<Ԓ9��B0<��"�ˁ��7�Ι���QU�F��C.K�j@�v`z0p�<��a��a��j)���d�\����	�L<t�C�8j�kQ܍�zd��ԒH��B��nȹ���l4]nH�SD|��b{K�1S?j-F˟��/^4�
%����葱TV%��9>��"xH5o�$���o:���0���c�QX�`ė���b
e��'������n>�As�#!���װ-'��0�W��n:�ߜ[�<��:��<xG������F�'�Q��*�m%�v(���%3�F�2[HE"2N;1�1��4"3d,
<Y�-�D;�xģ���X-�a�4�(�>
�j����A��*[�'��
X:;M[Bܶ�'�I,#"4P����I�sh$<���EE��ꎴ6�}2��<0ؾ3�9�ذHI����06
ل��4�L8'�t㵢�]Wa�%h���w&���IT�U�h�D�ȸ x���C��}r�=%��e6��R����uUnD�Æ1�9��Y�-~q�kuż��:��Q�p��Ӳ`�C�RI,��@5�!�E΅:,��.z$���h��U�E�a��;��J<9a����q���FFU�Z���s&�h���+�z:r���բ�W%[���2��������¡�[�h�0?�6+v�%ۋ�C�nt�=�f�&T�3�?F�
wP��gp5�J�:'O	�&:C!�M?F�H~��6��)
��I,8����.O�R3l��I{WO�i��]�NoQ�1�A�o��,z�6Y�IХ0tJ����x�g�m.���I2X!�2<l}��๰��'�d�t��I�q)��+d*��9ʩ��+5���:��^uż��:��Q�m�911+&;�vI$�T;fvF�^��l\`�����)��F��+A�;RO�$$!	�a!��$0�~)�����	���jՒ=�C��	G��~�*-k°x�<�%n��Xh����x6�߮s����C��x�Wp=3�pv��燡ʪ�)20�@�Y�Ǆ艂&:C!�8}�f���P��J��#S8�V�#j*\Y�#c�e�5SK�M�U$(Q.dB�8pB�wh��4Q�Ӭa���gZؤ�b�NǖSV�i�D������Il�u)���$�Xr���v�~�R�U�sy��l/N�a�ҷ\*�8}��p��p'�����W+���Ҽ�g��������)����s���RN8a�_,��5�!��P.�!3K>ԏ,�AƎ����XzgA�x%S�šq\��$#n!�et<��:g�D�ʬI�T\4��ki�ƕh��-����^y��y�V�:�:�-�^��O]ʲ�Il�$�m"��K4�H�ݤ2>Ctcq�.̌2�ۙ}�GXAaɚʿ_���"�þx�cu���"1 ��l!ī+�M�����T�$Heh���!Lc��2n���q��9&[O��!�j�^t�م`xW�(�����I\W=&Պ��+�U�n���2�4f<�O"�[�?D�0L�����b""`� �$�؈�8"`���؛,�F� �DK0N �Ԉ�Ȉ�&	�p�blM�I(M	D�T���'�lAIcr%�4x�0�<x��B�B"X���V�V�6��ae�Y�Ǐ�F�bh�8eT7|�r�Us����E�ϪBd�.�w������q�oU���k+h��=�T޻W���9Z�y�N:�\5׎r�PYÕǖ\&U�����[����������'Y�^_����_{z=�#jK����׹���=mH��wu펞K^�k�{��w��|�����">��T��D��޼�Y���-�ݞ~^o�ɚ�_^o�5o9��b���[ԓMˤ��;��Ϻ���﹛���g��gE�*ec���(���F��}5���<ds�w�w�f�YW;u�0�_��n�=�b���ݾ���{���b���ݯ��{����b���ݯ��{����V���}�Μ8p����u�mg]G\e�ڒI)�f��BMV��C��W�|˯W��;+���;�Tl�}=�<��ZCL��!�.�ЈN!��`�;�
J(��ǍX�k���:gC���
�s����xϼO���8l2��Gj�htdzq��[l0��b�����<��4#�r�R���-c��:"`��C�8>�Б��_=�I(ᇦV�����ګ�+��U�eWq~ۉ_{y'���db�$�.2�R�!H��-��f���DTH�6Jk⮃��gj(�֒Aó?tgC���g�����$��c���gh&~��H��YqF�a��Oq��RZ�e�dA�>Yá�4�~�_�醍�Ç���"a���æ�?W��'�{k��K��x�S�Z�l[UH���t⤮�
�R��a-�I,c�һ����=$����u�NAG3���d����-l��o#�rrn�k��X���X�Gv��KҢ�B�Wb�6��s�$���b��<Dp�R��%�KTiF�(�$�i�|�"��0���:��%=�$��)��f�P1/�CK�F�*�a�v��4tt6>Sۛrj�j�_v����Q$�p�[��*i�Ц4!-m1����#��pU�\��B��҄ģYU�knD��#C[d��!�o�s'�M�����X���8~�&�p�a�<t��b� _u6;G���,yUY�noI�㖯��z;w�*�2bC�̏M�\�lz�f͹Ĉ����'~n�y_4��k��@�g�~�m�êy]���"O4bߘ��H��Ȗ˗v)`�'W�쐄a���M�<r�;W4�34�$���$j_U�n�]G�:���[���0�4s�s�UUk@��K��p�I%v���+힬`�2��(�/ts�@�hB�L��g/O<�O����I��q���M�ĉ��A�eU��1
�2�#��Ɣ�f���|��w&NBM-�M�%����%��j�r������3���(��5�Ƕ	�����LDu�J�l+�mki��,â&�p�a�0飃�zW>�UpW&��L%r@�I%���}�Zg0����Y�m�|��I�/�9/ZI�0�L�0I_S���I�������0����w�4���=�Z��ل4Hɦ�BX,6��\��6�TYu�6h7AҬ�[������ysK���:h�Ǝ�8lN���:'����G8�%k�j�<�D�ǩ���9�B�L�)e�F���j4���[�66r�����VC9��2e���f�h��-��nm�5�VM��X�Tr�FDQ1bSaMF�
��7!��I$�������86�Bf�իP-�Z�ktJax��<]dt�l.C�4UU2=2<(q�d�bH��Q%�����OO4ec��S�7|d�5��(���v�|d'u[�9���V�4}s����N���s"g�����K��`zv���������X�o??��<��u���6C��B�Ģ|�m�i$y%٢]I$�̻?C�V늶�I$���\
n󃃫��O\K�Ūz�^�k��u_��j�z��2�u��W]|�p����q�C���;.Il��p�(2ѓ*�]V�+ĝBj,hm~:l�),�'�D�I�!'vCs7,!�p1��~��$���IQ:j�����ߝq����yǞ�!�%��u�rS"T�e��$�:w�\2@01}E���L�6x���x.�7�Uhxl��n�aT�P�9~�^S�2bor9M&���)7\5�'KlQ*Ć�	���>)sK��4�$�@SwI"����g�}a��&k���xvu�$*Q�u�N�9Xt�}��x�ˍ-m����<��<�����R��I��|�!y�����$�w�_���>2�<p��Ȕm��$hr$仌Ycl�ܴI25��UA�C�0l��&����<Xv]���5��h��D���3sC�K����0Y°N{��+����7��xkJ�H��i���]a�~�_������	�}RJ*���6�q?M�������[b�~���������4ѪTUQ������������6�!�1[����M����I-F�ZZM��ZIm$�-�h�-E��&�D�id��4�I&�F�-,�E�i��KD�4h�MDI2i��h�$�dD�I�#ZM"H�h�$�4h��%�h�����I-,�4�D���4�&�d�Z|��KKDI�ZZDIiiI�H��MK$Ѥ���H�K%����tI--"Iih��Z-"$D�h�ZY&��e��id�Y&���4��"h�mh��MZe�K$�h���dɥ�idM$����s��D�I-�I�I	$$�M"M%�A�$�ii$�H�4�d�I��K$�4�4�HI!$�Ȗ�,H�I,�Y2HK$��Y$�I��-$��i4�ВBI4�4�4�d�H�H�I!!!2I&�&�I	$�$��KE��I�sI-H��I��Z-"Y$�I�KD�$��I�L�ВM"M$�dI&�MZIL�h�i%�KL�đ4��E�I4Ii��D��i"�,�$��h��Gn�8�X�I���F�$�I��I)�I���I-,��4��i%��5��I-I��-ZIi"$�i"i%��$��4���DI-$ɤ�E�$�I�I��$��i#��4�"Ii$�KL�D��I����d$��D��$L��KI&�&�d�I�""&�-""ZD�"h��4IH���KKL��I	$�I�D�L��#���B�h[m,d#hY�6ІB�����d-�B�B�B6B�ж�	�B6І��n1��hC!c!��B�hY�ms�n�n,�ij�:��L8!��B6B��!a���F�؅�!f!Bbh[hM�&�@�F�?'6nhXж��24!�fGQ��	�d-�M����-�d&#��2�l��Bl�ozg�B̅�h���[4-�d#!m	�[:�k96�B�pq��BhHZ8��&����BB�K&�"h�4H�H�5�25B��Ëm�Z5�!-""�dHЉ���E�"�Ȳ$B$Z-�h�di���"ȑ�DD�h��"&�4DZ"&��D�#M��D�F���$B$B$H�D�D�D��"#���G�8""D"E�"hЈD�DD"D"�Љ���������&�"""h�i���"h��"&�m�������6���F��M-&�DѭD�dM-&�շ#MB���Ј�&��DE���"h����$Z--��H֋Bh�h�&��D�"h�&��4k"h�h�&��"h��"h�h�-	�	�"�"ݭ�D�D�G:��k!h�h�&�"h�4�dM"h�&��h�D$Z-Ah�D$Z��#Mh�-DE�M&��h�DDi�DD���#Z��	�Z2�E��2Ѩֳrn|��h�F�FM	�M	�&��"h�FM	�DдMѦ�hM4Z&�4&�hZ&�E�К2hDMBh&�4&�і�Ѧ�Dдw�]�74-д�hքAE�h֌�&�hMF�&��b5�H�kBК$i�D&B!#M�ЈZ&�"��D&�D�"hM&�Y��ƉM �&�FMB�4-�&��DѭF��M��M4�h�-L�I��i4Z5��h�kH�4�E�i%��E�i%���V�������<��sa0�iL�)�Ӿվ���U���A1��_�|�������Ͽ�?R{����Si�?�~�A��>��ߟ������"/�4B��pp?�������NH��gP����/�2|�_Qbxq]�(�E�O�������5��X>ϯ�y�PQ�QU�j|��<O�������4�"'�H�G��coÜ�$�p��w7�7�]���϶��?���?�H����.����?�p|߇�~/�����Ň�Q>�⨪������`�Ȑ��DE�����E>�~%#pg����B!��9�?��D�������4�}���!�P�T��	���}v	x�0! �ٟ���܏�����RR�U�fd��QP�D��)Aj�f��w`��i��2�����άl��v��h�����D_�G 5p����~�����f�m��?m�m���c��L���a���3m��ۑ�8lm�������>��A���"/���&���k ����������~���??��2p`|�O�<��|�DY�����۟�`�PO�h��}�/�2k�jm�
����D���!�?�l�?�� �����& ������Ը�� ��H}�� ��7��	�����**�����1��_r�����~ߴ��<��n��~C��
� �2�����R+���O��?4�R���Xr�����p����a{�M�X�tܯРDA2��$}��%߯���g�� 1,��`� �"Xc�kE�RP���R?x}z��T^��7v��6��\���#��r��9�
�ǈ��4�A�M������~�� O���r���y�+`~�����O�S{ }����?������~ߘ��������jR� �i��������	���������"-~D�~b�P��~��=����?#�t>*'���w��o���e2�
�YL�B�Z�Y[V+j��e
+P��YYYZ��������eee5eeejՕ���+VR�e
յe�[VQYEe�jիjյj��ee�����5ejڵmZ��B�mYEjڲ��+(�E
Օ��ՊԬ���QZ��jՊյj��X�V+��b�X�B�X���m�j�)�+1X�X�V+�j��b�X��V+��3Vj�X�ej�
�j�b�Y[Vڶ��jZ��b��F���X���(ՔVV+++��P��5l�YB�ղ�����+e
��B��P��L�PVյmEjիSV��EQMEe�(�V�SV�E�Z�P�J)��V++R�j(ղ��e�������jj
�MYEjjj55
el�X�Sj�l�������b�AE
�b�X�PV+�(V+��b���b�X���V+��b�X�V+P�V+��b�V�j(յ
j��j��jյjSP�Jj�թ�V���[V���MZ���ڵ5jj��)�SP�����V�5b�jSP�E5jj�թ������E
(QZ���Z��V��5
)��P��R��(VVVVVVVVՕ�b�Օ�mYYB��������QYYZ�eeeee
�����VV��ee
�j�ը�����5(��Sjؠ��(P������B�jڅ
+e+++(VP�B�b�
յ
�)�+S++++j�YYYYM�SթE
�Q���ڵ�����eY�+mAYE����V�5mYAX�V����)�1[V+�
�l�[V+�
�b�VՊ�SV+��b�X�V+��b�X�V+��j�b�X�V+ej�R�(յ(���YB��)YJe+QYEe��)B��jS(����mYEe�S(�QL���j��+(�����)��J�J�EeemJ�VՕ�+P�
P�em�Օ�����++++j���څee
��VVVVR������(�����V�Y��
V�ح�(�eeej�Ԭ���b����+V�VV����[VQYL�ըV�(�)YJ��ի(S(P����y���_����Qq��A�C)��m��ԧA-���UB�}0���c��B}��?x��!xK�^��,0����(��~�.��~n���䞂@�t�<����	�	q��n��~�¢�G��E~J�����p���?!��Ken|�?h���}a�x�>����#G�ތ	YQ�=����"�����?Y � ��#��?��
l��Y��S�b �|��%փ�p����/��4�}��@0���!�~˿�$a���p0��>B��]��BA�Z?�