BZh91AY&SY��`�)_�@q����� ?���bM��    �=ET�ƀʹI6[[f�2(I ���`�E$�*���URU%T��l�I
�T�Uh�e"�p�8�3f́L��eZ6eR�,��KE�5Y�f�YmUU�6)��Tf��3f�Q�1i�5l+T��dR�m��M���� y�u�mcM���R�UZ�J��ժ�Z�X�Ӭ��lfƊ�ʁQ-����X��SL��)2�����CJR��*m���e��,Y���WJ�L�i��w�
� ޭ�U�R�+B�u�]t�d]Yَ(�ښ�j���v�@��:W]�a�qR����9 ��k�l�v�dܫ�&f��LRf�V؍��_>��EU	 ]���ղ�a��D�q�� �N���{�=hPm�{ǯl�ݭ{�=R�#���Wl�K˛�JQ@^��xzJ������OB�Zv�OL*I"љ�-P�DQ�   z���j��^��xztTiz��ZP	�������4/+���*	���= O'��U(Pw�k�=
W���� � ���Ҩ+���f��ћAZ�Qjl�R�  >��\��}5b�v�R�<w�o` �^p�h�o.���M/.��v��L���B�{�< zR�'��l4���=�Ɗ�5��R���6k[&��d�Z«|�   y�|}�5����)T��Wn�Ef�o���
��<=*�9��hYg����)�Ҽ�=�( 
{ݏy��AB��{�OCJ{�����v1��[	)�M��   �4�@Uٝv�ý�l�:��*P��wU( -�%�rԅ���h$�Ζ�{���[{Wr��iT�n榆�ι� wj7�ma�Z�e�5����|>�P S�w�� *�x{����z��
z�gq�@QS���AB�4�]8t�6�8�T�Fnۭ�ݴ:��Ptwm�thP\S�����5��lJ�R�[�  q�-���q�;  � �Πt��m�WCEݛq�
1�q@��[�F��Crv*Yh5�P3c-�6����� P���
���ҁ�⻀�iծ
�؝�p �iΎ�uwA�Ѩ�T(��(u���GZ�ih��*Ph���   �@=�P  .�� (��Ae��@��@ ��� �-�ӁT�XP��      5OlU)U� 	��& �����*T��h� d0?%IQ�     ���J��h�     ��RJ��M4�d`�i��i�`�Ԙ����F�)�mC��F)���J5�o�UK���o�u�;���4����^��o�|k��'|]�9�ڪ�+��QYAO�PTW�}���+���{?�>g����v�D?���+��O��Ѐ*+��,����D�
�����O��?q�G�$$p���0��G\$p�0��@�S	�\$$ !$$L$�	�.�  $p���W6Ha��@�G	!p�0�0�� �p�0�0��a h�0�0�@J�0�0�p�0�����@�W	C	"C	C	\!p�0�0�0��a a l�0�0�0�0�\$p��G\$p��G	L%"�@�			\%p�0��p�0�0��T����������l�	A0��@�CT$Q0�P�EQL$�&��!@0��PP$p�D��"���!0��EC	$0�@�	A%0�� L!0�D�	�0�D�P	$0�P�T 0��DS	�
.":!Dp�Q�W	A$0��WUp�	E$ 0��C	A%E�E\ 4H+���B�l�P�	AL!U�Q\$E� 	DvB�%@0��Ep� �p��G	!p�D��B�0�� � �	\%p�d&�$!p�� �G		  0�!p��W	!p�0��	\!tF� !p��G	$p��S	$p��8H�� p��	\$_����ײַ�����>;�����ں�M#1-��56P�ca[���7&��oX�hyK��a>m�Vj��«8�����<��i��R!$�5�<&&�1-�^�o�����e��)��	��<7�U
3Fl� ��M=p��+#K�iٶ�S(��0I2����m�$�j{0��m�M�F�_��C4k�P�=[s��;u��b�Տ��$y5�4�̠�X�����wȣ�Mj�g��<%�1�	(�"�obʳ���ɶ2(U���0��:�^'|Ǯ�d���/�0�
��Gni�"�f�F�#J�������&�1�h�cƄݸ~S�}U�Z2������}��36�RO&(���}��2���Wc��K�%���
j��<�SPGltm�0_m#�ksM9�]&n�j���e�n	3qݯ<�w1|ߔ�q��;�h>:�����3&Ob��.k{g�k~A�;��Vz�3I�,�hmia��kXB��j��P�-�kr�#���$���d+T��ۨiCpWl�<��.˞�ٺ��X��H�H�|6�U�ؠ�����U3�eV��Ù�%����C�E��Lo��4ٯjg���//  ļ�P�?7�ŒD ����ԋwYtQ"����o��f�7qM��F]��HMt���/^`KEp)w*����Wo�z���建}�����
��C	Q��1�=�+��^n�"G��x�vǡ+Ёr��Sؕ�f�b��ش+�<x��z��r�[E�ã=4��
�ǣ�s�sA��Q\��P���`��[��O�F�pGH92�Zt��;�o�0Ͳ�v�[âb�Y�dxVn�3X��Zܛ��y�(�fH��
�R�Ғ���F��q�w_.&��i�o�u���o�T�=N�U�Ͱ�0/2��P��nE������Z��R�#��p).�}H����i�ɹ�r��}-Uxi5�u�눡���|���lҳnk3N����Ɠ-`Z�{�c3ۃفW�d���(�6�o���{B���K��@jP��[��+����'�LJ���lDS��#s�Jj�j�!a�2��ѧ"�EVjX��ԖU�;B̨��.<зnF��=`�@g`�m�0Qy�5m�)<��f���S(�Q�k	���V!{���-�L���-ѹ�|���f9<�^�Җ�C�ؾ�^j���4��X�ee���,�),3/q=�-`��z���$�T��+%F𫵍�փLј�����Ϫ�WA�P}�x>N�|�"����^x�wZ���X}
�,�En��=���dS=}<��M���~,�v�ޭ�TY���ZO5������qO ?�V�%	F��͑�U�Z��.�o�p���j�tTa��{�ێے�x"�0�h��K�LJ���wt�Ч�bz»�ۇ��r�}�a�b73�>̤Z#�]z�zՕ�U#��+);FU�I�T1��%��f��X9�T�NEDQCDpK�ˢh��k{��~�a����ް��G��/sn�Д��3�'j�^-���*#�S������E�n���ȖU(� ����f����V�&[�B
��bE�m/*/o����3d^����P�&�2/k;p���Ő�-w��w�<"s.�C�P�;��Sک����#�G����S^F6�������=!�w>aM������j�p�S�.�vb��)~�Gi�(F�Pn��Ӆ�d4V��	��*1a�Pl��Y>�3=11�~�$���ߌ���~���p�i��?J��2)͌[<�����9EH*�Óh�h��)�d�lZV�o��Ӛ}7u=!��`J�w���[J��<u��FAs9�H��#�8��©���F��ā�B}�ݥ|�c�-�Ibf�<)>(�2��t�"������L��+=����ic��L�ly8P2\�NѾ��g�:�+�md@r�ॵ��[H��Y�i����<�s'�7�廩�s��hN�yH^�-T��3*��#�~���ߦe�}0Z�J0f~�-Qv��Bh*����aG	�q�)����7���,쭹W��z�v\l���,��6�����ٓ3o�Hךf��u�n93d�����"�w�#��� ��+����(g�*vX�j��)P{���7d�Vպ��ZH�1,%��su���m�~���_-վUU�L�h.ƔY^
�<)����<s3��S^��!�6
��+xNỒ����D���FP��xn�S�5�j0"�6�Ҵ]��&��HFM��v�n��Y�7D�ܵz�
��6��9%de�<6�(S��M����K]��J:��L��Q]�!�i�^��Y�&�� �.�v�n�툮*X�v���l*��)eˁ�Aϱ<�"36X{�qAH�Z��b�b[�A�����$�[O��
�'�۱4��$K�d T�Ӻ�6r˙�ݚ�Q�s��b%�*�N3^��n�Q۳
[�/��@j�KK��@9�g��qp�W|��Uk]�J�Ǝ�±;m�Q������h�
�뽬�� �sm��/��K��E�"�d%���C���O�vy�t�vH��@��}u�7�ꩼY����}[�r+�1��֎�V]��AF'��Ϟ}yr��X),�2(�!�>�I`��&�ʐ����.T9�(B�b�[�b'=��Ix`f��=���:�Ѩ�&�}���_ii�na>�s~���=��ö�����oQ�[��\JUPj����0�n���jH�b��M+��\�>Z����Y��Fm�˂ 2�|r{`���1`�_H~٦���L��1���{�嶨�9���a�ꍒ���i��zF��r�&��}� ���lờJ�r<h�b��S��������yJ�h{����eEh��(�s%�>����� v(U���f�à���i%�Ǣ�:k	r�7,XzΊ��A	l�5D����1�s 3dN�ō���/�8h�5p�4�c%�**î6�����3}��T��.�f�7Mr<���P�ᤊ�M�Ҷ7lz{&z%�P�q~�7^��s�-ũ'���dCA�E+�b�8�I&�WB��{6���[���yk�c9�Y��Z��t�������2W��++͘vt�r(���J�f&f���e�Ӏ���z3q��:n�2-�l�j�4k3�P��L���tAg��N��/�:3nXR�^M��rb��X�3���k[�N�ns�O��$hh7OF��-�Wl	�F���Sa�^�<5�5��˙������>>�8�yws�T��v�4��sʔ�������,wtx�����n���o<���)��Z�DE��n�����p�|}��M����$d�$�6�
��K�烘��l^�Z~�5���su��f�p��W��r�ܠd�p��zg��չ�
�+��4�zi̤�'2�"�!k�g��q�z-��������Z�0l��wvm���ڲM���p��6m^�ƾ~L����O Gw�B@H34��L
z׺J.�Ur{���g�b��F>5ϗ��[�	�v��XH����R�}Fn���_��d>�	6P_�f��kg<��}�6	e"�ȓ��.l�0�l��g���ðV��;r��l�3=���e��*8�׿�E����:8�E�4�����LB����{�$��9盂,�V9W����7@(X��{sv�$�ei����J��H�5}�I�g��WS�zISsA�}�ᅓ6ƽ�}f�nw3��1b���^�{m��N׾����r˻�M3ƨ�~Гwt��s7`��mm���-�C�Ɨ%^ Ӭt��s��C��ծ��$��Q]Jf�ǻ}�m1�ݵ��%ji�(7�z��bHP�ؼW�_Z��M�n2�yg����E��&�h���
��xn�Y�iv����ffI��w�`~[��/���&��^���3R4^9�W�A�{��d�̆J��8)�uQھmj�oks�Z�y`d�{cy�J/M��C�C+5_sD�w�!;����G.77�-ىF�X�^�o_�xl���`�<�S�`Ŧm�n�%�j&n�Ị̆.��A�5���׍�[���H4�ˋ+��8�gi��e�F�N�~� Z����ܸ�L��7�l�/;d��(`�2730dA3.YN�Tuz ~���os�1 T*n����6�)��`���A��#��	�B�;���z�bX����J�rzzV?V�W����d�'�n�m��f�`���Of����e��l��vA�z[/��Ǵ�\�W�D��p��'�O+%�L���^�W4Q���ڱ=��^:�Qxj�O�4\r�+ϊ׍'�;�s-1�t��z����ѱVТj�a@��%K�\7��4exl��҂��dz��IE��.���b�
�&L�wml�uÀ]�]��d�f]I=9$x2�Cy&��t��m��B�:�Z,8��r��Tt�jf�Jӻ�ud��&��������+^�9�k��0SX�����fU�=1g�������7�L�M^乳u���Ƀ
Ww=	/g�TH��<n��s�M�f�A��Uċ,ɘ�X�o�
m�G0��9�iL�SX��֢'�^�|��^!S�Й��,�33��
m�7؇��2b�+zXc7/u),�UG6�����(e"�I\��hܞy�5�sO��d���Af*6�vz�T�1"C�f�$jN��w2��)�ն|�nǻu�BJ����N��׉�	wU�� [��`��n?[��5�F��'2ֈu���/*��(3L]��:&a��A�W�J2iKF�eKw6Ǹ${��ѷrI�|�׳#���R�f$MS�aY���djg�V��n���Vw)�y�ùg�/Z)�'Q�(�1J��!mê�����jY��3�4�pd���ԡY%�z�� �(�+�]Şd�v%�1��_�պv��ƀ�b�b>�]Jʽ��<sAo�S�p��[��&�y�8�����Ce�_҇�gs���ckFd�ӵ�Y�:-�u4p���Cs}2
�Sի�
�&k��S� ��O�]���~lї�$�M�7�(T��oE��f�sL�BgrZlf��y�A�uV�Z����=�k�$�����)7Vv�#��[M�,Ͱcû6X0ٴ�����(�C���^sd�4e��6Cۦ5u
���_q�I�ܛJ�}��,�k��sn��qc�/=�A�kl�7����Y{��;�l���(֌DfJd�u�;c+�Bl��?��R��*�a�^i#r�h�h7/n��kI�c^���HY�j����F�o�Z���~����]�Č6C}�OXBu0�e0��9���c�J%J�ϔ Z�O����@�-���K\���[Z�߲m�Z�G�f�N%� ���F&�w��)�R*f��t���Ug���;4��^k�/�Y[4n�1��2`i��^P��|Ջd,`��f�X��ǰ�PZ�Z��OlS\[}�ِm`I�г����1��e�ƶ���h۾����l�N�ƻ甤�fx�t�~ib��ߦx��0�C��Y�DAZ��R>��븴�^�����V������f?%�$�_3�&�7 g�[�b�R�,Î�'r�w]ܤH���!�mA$��T���s&Q���Tas0��
��Of{|��o2� `ͳ��	]<�F��DB"(�ui��]z�fR�*���S�
]����&�	
ld��}�wv���컇ͦ=��Xsf����+�*s.=����ӷ����� wq�%g�"n�����<���^x%"��J���
��NR#�ݤ%��p�T�/��X�֐�sg��g�i��Ǵ��M��/ek0d,� ���siCP4ߞۭ���^�$�Y.�H}!ly���mQ+����W�����H��W����k��^!��h���4V��n�<M�9�
��V�9[�e��'K���ͭ�I��3q����56�.��yb���u��e�ѳ\Eeaˤ73}6���HO��8}��Rܶy��?B~�(���1�\�w�H�`/Pp
$h6��d.��Ȥ3l�n��M�+�7t�6��'u,�5j%��NLhEA�
�[)Ւދ�y��l���:��="���p��i�Fjk�� ��>�'�\G|vBǍѴ��F����������*�Y}�M^~"�I<���˶�zA���2�߳\Ȑ�^A�j�!�L�����&e>��\����iT�*�Ӊ�l+�4^�#F9z^�*e��3E�D.���3|5�Z��H[�B�Ʃ�$�ghm��d����h�q�BX�[1ʞ/c8��7ےcwTa�S���Dka{��e�s�ePj�;�'�ۯ�Ufؼ����;�X�pv�[�̊y�V۴���*�JD/`Քʟ���T���p��Z��@d~�6�_FWQ��3"�i~��w)��N��~X)Wۀy�Ւ���%}��_����hX�u4Wh����5M�0��c�.��H�^�ѝ�H���*[�7���h�hj��st��]��eF��g�靹��4���J�F�LqOn{�\��2�	p�&hv!6-���īf����j��/{���]I� �l�-�cj s(�+��'U̚6���?2��"[�jX��dUGn�:k\!ڽ�{��=7CC��餩:ٻ�h�k�E��-�z�oe�6h��<Ȋ�q�<u>y�]M���}�?Y�_h1�e��\�����)�dx,,m9k0�h�)l�ջ��9m���[Цn;�=u���aϯ�@�������"3��>������xbE�y\cG��Sr�-7�w�[���f��)@�=N���#q�y������yT���W<�~h��J�ᾏ�2��j����k����z.����55���i��3���-(�����rW!X�pݙ���$�-a���K�JHs��}�f&v�wf��7��L���Wge�-�ۯ;|��h�����X�g5m�����s�3a��G�磯6M��h�1�.o�yI|�[G&M�\��\��.Wf����K�\L�Vt��N���0ͳ��Y���A�:�1N&��܂l��,.iYKf̚��凍��N��М�T�s��R�w:!�KEG|��:��d��|tNRwu����Hgq���ǔ�r-�d��±Hq�S�6���s�E����6��
�,І�*٭k�^.٬�.�B�[1�QH���[� �{\�oA��W�x-퇕���pL��c��1�w��^�K�(L�YRS�O;s2�����B�ݸ(J�Z��w0������Vr�&H���lX�4ye���f��g������h����-i�D���w�r5Ba��˼�����y�02���D��+����Sw�k�J]-���]������u�O���m�I\P�+1���ܧ�*��B�����e�ξ�J��{q�I�[U��r�������H�]=�A�G��*3�Ǟ�q��~�Vf�n�,7<�(EI�zW�dއ<s$��;�S���;�9���һ�o�j�C��v�Φ�-������Ӥ�n����vG��Uw�k�YD�Ó�WЌė�^�x�w��<瞶\������_^�x��=n��l-�mYi�k(���E�
۲�SոfVY,�E�#+6��5lj{Ə�`���N�^����d˸2���[�j��Rn�n6��#���Q���ʶ�6�ܴq��������?X?J=�;	��Ʀ��O���sb�{fsS��ʮ��~Vgz����3u@���)EN��)ν�;uRz��ն�1�]*�����Zx�cfTF1�d�۰[��1A� ͣ��<�W����N6O*)Gn }Z,�f�#j֌��MU8{�����UE�pб[�������}�t��34�� �����>pO;�����~��#S��v{�D��Gn�ƳMA0�k��M�s0�/l�U<v��\��w{�1B�)��ˆܖww�#�H� �Y����Q�u�������	��c��^t;|���=8��L���7�\�uk������aY7ݬ��/�֔W�{/o^^�v+�0���7{q�>��KG�˜K�9P�߼��YfRڡ����}��ӏ���T���䓷}0����yCd̻ϳ�%��
�#�|�{�ś3/UM��9T�w{�yCp�A�c)��9ϒ�uFL�	[�?u��D��%[X�Ž�Lӗ���L�1U��J��V�T@��p���v���r�/31��VE�(e��X������m�?_7�_����v���'�*�v�)���V�4v��[��C��9K�=�Z����o��0�.�/�H/yU��:��OU�i�[S�f���W54�nv�h����ؤ���z٪\�!ڤ�7.�����H�G��vm��r�NG;�6%��.�<��y]��i��G�g��] e~��{.�SJ[9�Y��}�%pwۉ��WΩ��XRS����Y��ɣ&��]V���s5Tצ��i��3��J�D�)���&�Y��&�;[�u+ۇxf**��r��bI]wصGY�1�V�1��Pߔ�{ǘk��ZGyw�"X�n�2��EVS9@�� ���7�һ5��^	�����ѣjLEJ�6�� �`���wv��>o9>�04����}r`rG`�bQ��7Z�܍C�6s!Sn�>ȥ�<�:�~���sp:@쥹�3t�خ��=��.���jC���C6��s2u�;���/.�����W�7��U�q�9��+��xȸ�z�V�f�B^���/QC��M'"x*�4���U4�a.��ȯ�mJ��EGr�2��.���qoq��W�1�5��9�p�2����<���������Ӷ�W��.������R.�{u��9#d[�(*���p��9��`�b�}&zV[��d��TA��5�X�R�Z���H�R&�r������P�![ʈ�rUg*�����<e����c�M���ڑpkS�8ȝ��d��e�鸼���`�W*�c�קi`�,,�'dy�܃�gwb^�n)w2e��Ҏq�Tr��+��'5�����N�Eڂz�W-�gE�
�f��u���:�������Q��kw�Wu���|#Gz���C�LG��Ѿo��Ω���a���$O1BkŔ��x��e����Ђ�˶���^If!�ᕌ���/�ҘBj��w�gk��n������������+�f�=��J�׾�u��v<�� �'n1�R&��2��:�VV�{�؝x�(RO�UQ{�+з��*�I�ih�LTF�0�&V�\[�1;(f����sT��X��Cyo&�a�5�U��ط"��8^g뒵r�Ą9Pk�+��ɻ�+s~t��¶*�HӕdZ�c�h��*�^6/�v|��GOt�*�w�9s�x�kZ�v�v>9׭��ڱ
��0o<�aî�or�m�<K�yO�滽�:jݽ夻u$�&Η�vLS;��t�=;#`�Y	9�nn3�>���eKuY4�׺hv��7ܳo�t��趖� щw�o�C=SϬٌ]�f��Q�<I��a��G����hi����
�a�o跱���RN>́�-��
��GV��u�ú�Z�w�oH&Y�ѽ�N���z��`�8����֮Qб�N�u/s���4�)W�EXS�.�X�y�z�q��'0m�؍���yg�..�R�U������n*�}���ӏT=(�챴Gz�ؓ�����$%v���Xvěsn���h��P.�G�;�\���ǜ��`�skJe��!I8Y:��XJ�/-C�؎���y�yf� z�d�{1�yu;��/�vj��-�DH;��1gpb㇉#$�jfw	��x��z�'��g�b4n�ވn7��k�a��a��k���������{b4
_���4��$
#���E���	��T3n��bV){nvry�j��Os/�	|�n%5���|�a+m`�I3Vf
�sj��O�>mW����`�i�2�X����gfIP�d�=���P�$�+oo�ξ}���|�/L���T�nE�J���cu��f��i��@���k{1�Q����Y�p�vZ#�N��t��R�&��9b2��}����)��o ��:=����<FG{z�;��jO�W,|]od�Vþ'#/�䡩g{h��OY�U��[�v�ts����=}6f�=U��B���U���v�z�L4�f��M�6�!m�s�y�YR�]/��0"k:��Vo7�6��5���n\��WS
]��K�*F[�xc���w_�����;�c�,��Ӎ��]4����M�V���.;���2p=tA��Tv����=�[��������O�#���$�w��xM��UaojA�D�ơ2�f�nvl�=���C#�����[߇���p��*c��=�U�w�h7����N��.��:�m���L��R��?����V�k�[JW,������64�@Z�V1EDV`���#]�å=��y�L�MK�u��\�Qft�?6����bF���٘���ٚ��������
�� �R�Zql�p^�K�W�=�ǭ������V�a�n�VOL���ܬX��.$��2�� ,<?b���|����SX�G��x�9�#3ЏYUc&1���1n�.C�-w<Ri<V3��;��b�.��n����E�C��G���p}Ⱥ}Ni})�9�n�6��d�I���w4iR�=�'e�����پ���Z�&����zl,�=�s�+�M7�En���H����8v�M^g+�D:�֋L*�͈u��#�:ʔ���|^s���3�Iv� �V�gC���al�+N��9XȲ�z	h��x�[��>qۺ��-_j��i�q��d3vlMih��57����s��Cq<�g�h��q��ɡrt�q�>~G��w�x����#�Ja�/N� ���U�<g���D'b5�kĭ�Y�Üh\�:��;�B��PcfƠ�2�T%5e��ؗ;iK���v������w������z����ޕ%.��^��O�1
�엤�8�)�i`g�t�	5����9�M`�t�N3)�;�;Q�1�(z:���eC��-;�x��3c5W��Q{X1�bomfy�b�K��	{k��;�,�gZS3([�,�Ł���)4�m�V�cGjs���ퟥ�Y�c!x;3^�]��QЙ�}�K.��bg��7H��99Z����x�F�q������e1뜴��C���6�����C���;��-����f4�{[� �����/+遱���-�c�Dk�'��!��9r��!Rm��l���Z�׏����{���>�,˹����W���q6"�Ő�g0��cNe$E������$B�nf��)]�7��$��⺷6Y<>�3�\2�"Wj�{���=�5p>�$�ež��\�h�{*�1`��H�h��zS�n�Ɔ~���L6��//��xw�|&<I^	Z��{:���sb�S�u�����PO\�04B���p���ƍ��u� ���'�x�σ����FnW2T�l8*Si<��Zx�rV����f���!f$�n^�/Y�0棆�D���l�X:<����׶d�y��P*z�v�
ZOWV��f����L>g8�B5V��1jE���Ru�u�t�i��\�Õθ?�(5��������mjz�`�(���^#:�7D���v��w���!��aZׂ�{��Z#��ǈ�B�Á��j�	�bΥ���Ud���!��fC*��}�a( VX�OH��.�q]dl�;r#ub+���U8e>��X�9:�&Y�9��/-���K���ۗD�Nv�NE�Σ�p����H�p����`ܱ����4�+�9�؂���K��s��3����s�*�:O7-з���؛	Ji��
���%pٹ�+�E])���ސ���krm��Jrҷ^#\���Ov[��Mx�������t�)��U�X�KJ���OG8����&B;uw%h��	~�	�6G�n�ݿwS�U���rN<^Vi�B;�x�sz���35i��F��oI}����� ��EntA=�υ%�W��#N���d[|���`V�a���
����]����L��ْҽHauI�D�dUs���]�*��I��/^=�\�g��,B�r���4��5��='Ip�Qq�L�^ś�^�̇�.Ǉ�{����X�4+pv����H<��seJ����O����c妽��(�-(���>�Q/<ѕ��"���"�tz�Ͼ�̆��8e�jL���gJ���ipWg��E��%�2�f�J)�Hl4��r�ѹN���Usp.@7�J"٩n{��?=CgX�z����m-リ��p��,�9������5�d����ِ��_J���C����ֺ}�)�3��o�ޅ��k�+�G�_L.�z�79)=��Vy�$�3ں��)�SWwf���9AnVv�X�.�#�c2N��VC�&����P��78Peojl�5��Ӵ���,˃s(�>#���%^7���]
6��hZ%Hko�.
�f�:�y��-�������,;
c����y���z49�3�{צ�f��+;��l\+�ojVHZA9�`�0�.ܷ�Q���Ys�UR=��x�8����M�Ǽ�����Lv�w�~^j���Lk!N)�����mu}�{Y���s�ѻԜan�������E^�lJ&�5U�Z6h�Ż�A�HZ�u������XU{�z����Lv�=���c��Kq�ѳ��p��G��
���E��Џ�̓���NA3b�zb۪���j�4�9�q[b�}ى<�nI��2�������ۜ֏=�\\�9�S��i������]=2����]�5|�ms�^�[b��r�Q^3u<�o�y���;$7#�6C/Ȯ�=�u�y��%��n��XԠ8s��rs��ѐ��I�XU�,�S l�;3�+Fr�Uf��:Rݹ/��:�.�Q&ƶt�Z��+�p��ey�$|7�[��}vm�i6*C%u�YmgH����Ya�D':oNwRoFB�e��E:y��Y�F۱g�!�Vo��O,�d��k {�OO;
��V^���YEN�]�CB}'KL�U��K��;�\3+�`~_�C��`Jn�:��"���J�Z�j=Mbr�Ru�i�O�ZG�<A�]�u���h;�Cj7��Ek\�^�\��t}v'+�50��o4�yz��y�v\�	֞U�&ZW��P<n��Ӳ)Zq��cx��]�J:�1��MpM4����*^�N��Je��i���걵�E3;3fEM�Qɕ)#�X�&�$�2l�U=�0-nL������6�=��+��X�@j5{z�J�Rbvƪ�j�=sY��k��:�Z�i<���sk�R��&�γk�qr@�@�o��LL���-��s��~���'e0�u~1�q���E �泽U��~�"�<b�zݣ������n�u�r_Oh�{n,�nB4�(����Nڳ4��%�I
M$�qƁ1���T	ʉm�)���A��� $��j!�*���j�-�rO�ec���8i����Aj��h�財o�� J�RB���(V���Ht)�)nl�5T�./��	1@�&�*$��\�Q �f�iY�%гdn�̨�x�4LwҿP�m��Q�Y�T!C�$��%��#�J9lCr�,F�O��\��$Q����n���A��T�"5N�(�!�hs[�h
����V��z�����<����������߯��}g�}=��u�ru�?��Q�{F�k���]��FV������fRբ��Fߞ��B�@.u�)3��+��v:@t�[*�3��P�FŚ��@�\�#V8��:{4R��+pV�.�z�@�r�����q;�e��.������$i]l�?q�]�gLy�+�����yW1[�䑧Q��ۻ��-�i��t�<��LG��'!�3��5��!��O�]r�δfGU�7:�� G�v�z��}Z���M�݊���k�/ac��iW�N�L�ʀC��۹)�ۦ�feD�γl�l*��� ��~w����@�!1����^h�*�n7ԧW��p"�������ꗦ����uU���u���3B�H����vgge�8���;CҙR:�y;��'�U����̫�G/B���X�^��.欄���<Q/���g�#��뉍�\�V]c�sL�z�����܇��7E���v�;֏��(ᙼ�Z�/����Ί�ꦷ��;y���L��r��r�P��x���{��XIzV�O_e�"d�#nry��;Q]�wj�6j��FE��I.�J�)2���臂�Y��Q��5Gh���y���>����u�ـ��]Bn���(i7�R��gz)"w�j�t�n�E��`�uo���U���{w��i���A3�R���+ke#�{�J�K;v.썍��8 �P� BA �" �� � �AA@ � �(`S��˃���I��!?z;^����.2f]_b��m�'O[�6ѹaa��C�cL���Us�7�_c�[��a�[\��|�q�7���yF��C%{�zSbN{,^`���ѰÎ����5	�5ې��ު�=�Hk诜'p`��euN�U�t6�q���͕YP=�ɘ�:��/J�P��M{97�u������~���O9s!�:�ά������C��v--�c��û�E��[�1����p������0��[~���Ȥt�8� X���^H�U�����2^`�o�C��w_\t\��U��ͮ���P��G��_"���ҏESU�j8��=��&6������v�r���y�]Lfj�B�n�[z�X�bv̽�D��O����ve�z7����v^�6����&�.����O�>��;Ww���0�W`�xxm(Nֆ!���@Nk��=����]\;��k���_��嘎����Aw�+���&la��-]���W������Y}�xңۛ�G޳.?N^l�۝������;�d)�:��4n��M�}���wY���۫�h�'ű]7h���/�\綿{G/'7h;�H�Y��A�0�9s���\�K�b�/nLh�b/�:��oO>_z�3kR�מ��w5���5�ĽO>�ݑm�n2�y1M�Ο�=�Έ9�S�7!{�R'�=*릻�,4,X���A� �AAAB �ŋ � �A� �� � � �� � �yH��d>�?t��Z����-N3���๟M}ۍ���O'�=)#'��vC�f,��\�_�Q\�Ɏ�i��=�T��v���}�q�=_}e`=��`�#.L��]��0g^��A��MQ�2�m������]�Y�V)B�a�k�� WV�6ܨ�U�t�'��q-s��P,ac[R瀝�f��{���p:��eWdc�*.�Nt��"��@�q1�U6���㽝Ƭ�u9�m/�<��r�靘�L>��/��S!;J�͙�ye��4J��[?C�7ًŭ��x������
6��]��c�b��gMM���@�4n��@�CCLu����ai�L��x�)�p��6��uȎ�4�޳Y'VT������/c4j�>	S��Sힿ|��pw�ج��RK�\���-.�./�v��i�6��˭g���Ҟ�U��Tr�۱jh��SϬ�^��WsY|9z󴼞L��/�l;o)�ѻs��(>�6��j��gh�
��׊�"M�1���g*/��B5j鋱˒�ˍ�n���{��l�
��Ӱ�6А.+���E�Ҩ���=5G|��v�4SE�j#Y���f���2�:���څ �pgh�"��F"~ݾK=���*�k�'�ud�/9��4�?�B��PG��"j1� �ل��}���q��EK�Ą����ӥ-�Y�,hB0AA� " � BD AA �A��"�Ah��q]���B�����Rs���h�s���U��RC��=է��ǙZ�YX�*�l��9;z���<�n���Ѫ���G'^TX
J�	�X��P��PK�+�f�SP�������Pq�}���t�>�mk#��>�Yϣ˜w�"xڰ��}�}z5���3���X�LZ&�\�O;�ԅ���ռ;���V�:� j߹q��{+ڕ\뙪�A�`�K�^u����.}/ʫ�V7G0�N��]��#w#��u��rF�#!�֔����)C:gu�́P�)�cog�hO1���AK��_���zb�x�;�m o#wzf݄�4+��=�}���c�0L�]j]���i�0�E�ÚsZvee�δv�T��eǡ�����*����_a�PN#]��p�t�Rٛ��&@;�4�og�w"������:a��7È'���Iʱ"�-���j��SP<�UߖB�t�D;�ug!v��zܺ,,�\v�&y`5�O#5�۬��;<oi�/_a���g�n��y�l�������=�����܃�y7'��S��wh���}�~�,g���}|@�Lf�T�5�����7�j�x�wP���
�z?'�"�f�Ǜ�9��L��4��F{�sK�5a՚����o��5��0On����­̕U�$ivf�6�t��V��BE�co�ro�+���Q�U\O��AA�4Ap�,AA� �AX�D � � " � � " � ��ɕn������]���E�=�i������ܛDL��P�\/u���:�&����6�x{1s�X�T���,�q��]�6��z�_a�?K�;�ƚ��p4,�f�豗v[�������������?I��'�s1D��h���q>�\*��4��5[Y�����b]MV�:5N�n>�M/l�mWh&���7վ>����T�Zr�S����(5�����qxB�����o^��r�����&����S�yn_j׼��z�Vx�S}oaYw>�ye�d?Z���tS���G��nR׵.]�) ͊�KZt��"{}ɾ�wo��K��)��"j�c���4�b��z��Q����0��@���Z`�*����(����ߍL�Pxk.�[hnMC-�d_>G�.�X�j.r�;��O��;�IX�4�Ĉt�7�sF�XON�����VdOY���{-;WpO�1�I�@�ˍp?
�v�m�iԶK� �_�b���Ŵ*��O��v�wN+�4t8M�d]�Ԟ������;���Ҍ4Q�0L�G�=~g;>=3���[/��ޝ�7	�&{�篺��]�$�|i-e��ug�)�|Ļ�Zu�팑	�p_	+~��C�B�Ob��*���s�!5a��eöhnک:���?�u�M�N��u�z��Yv����#|-�zJ�2�E�(qIF:[�#z�S=����H=��-���6���gp܁�ޫ u}b t�"��;���
�������~A��6��y9��z�҉��A`��%�sn=��jL�Mpw�ri�9G4쵖*c#gO3Y���z�x(��$�\~կ`u%�őHuWi7�iw��mio�f �g�ʼ��R��/<�<�o�a�e掌D���~w��yD�a�z�u���o�#��]��L���X[�+�nm���6��u6�սD��<H�B;��B�gz�/q3�͋�I�ƹ�=����=�ve8�k;4{'�7h�0��.e��&m��W��a�x�l�ٰ)-����B���徱��&�ke��ɪ�����`�*����y��;3:��;��1l*l�3�J���ŗ��!!���gL[-����(έu4���vш�Gb�`�c����Y/�koI��^xv{�^m�1o2����MoH����jN��b�&�`�ғ$�z�����d�]�A.��bu���.������	r���q����IQѝM�`=k����>5��B��J�4m�<��0�S�6s�e}����ԤcZ�rޝ��Դ��Ppc����=�4�<��!6�rH;�^ȍ�U�n�㛾��d�L����\����+�ۅ^���o��a1XƘ7��.�r�O��o7>����?-���}<zxkþ��px��_��T7o��L�n��cgS;�v���Sc�}�Vnjt/���h���e�j�ٷs�3/@b����9{�ݏwW�����ˇ�x���rm�l�;���վ8���B1Դ�-����l�s;n���bO2��� �J��̚�'=q��P�6n���W��.�ipL��x]	nu7���Ws���$;�E3��-��K8����v������"s�ƖuE:���r��G��ϸq�+f@�؎��֎]�\⻫fk)0�y�CN͝�xlho�BUZ��1CvG�I�{���ovD��?�Ts%3��ޓ�d�n�q"�4��;��t�>�VQ"*H�t�xN�⺻ԹnB�� ��M�w<	�|���m��L�m��&o��^W֢{�:#��1(����79r�P���3�·�U2ʊ�t�^�|�����|D���r��Qxz	p�1}A2�.ƞ�/o:㙪�V�1Q�	���ź���kIb�c+y��]X���A�Z9���Wv�r	��	��Q���s����T��E�ꠝG�o��U ��2Ptظ|���v����U�p�e�sm��{*�92��;�k�=S����|�fޫ�~Y���|���T�럮���ncs�,��nG�����7���2�j��o@��1�(��q���*[|�݌s�|2Hv@`��C��{��u�C�E�f�8.b�V~�bں1GmM6	�a��9۽�˱(<&9�:R<�QO{,�[s�ș����֖��zG���l����n�Mm���eU�6x7N~�Q5t�
����m���wL��:��l�v�;��yDY~2n�1�U��q=w�Ɏ�z7��oy]�78^���JV-�{IW'?ja���W�~ܼ9t��aM=���ǜ�^���g�}��'���Wc�7q�`չG7�����76,��Q��{��ƣJ�1�ba�r響k�#�MW�[$�nۮ������ٗ��ߍ�6r�n�PS�+Վ֪���K��!GPZz=�2Ș��ú���~�'���8'�`��/�{��0]�ҖYs<3S癯�S��^��R[Y���5ϔ����5,x�y�����=�xN�p�t��1r�q��A�(���a&��m�΅7��{��'=��ʗ�͉�^�������3�����ϖ_rۗ9�OX��ӈ�{:N�.�	�fze&}��w��:y��oi����Q|���c�ـĪ
7�����z��Y*�
����7��Qw|`�b���C��rt�=����iG��a��A�M���ozj4l�6cR�z�(r[u�і��k�x�K3���[�����|�0�s,��xy}�0����7�OH�Bxp��a>�>�S�7}��┚ۼ%��O�p����=�|:�:�V�<��v��T��Q+<�1�jT�pz�4�=�iC<���ލ�/�A��jv�]ͳ�e�{pU���j#`A��e>_w4}O,�uU���	��7o��LtF����Tt=΃A�6Pa� n�u�����O&�\m���䬡lG6��ݶkK�W�gH�����@p�w��S�<�V\�t�嶎,�U��uw�]������TYMi���$�m�{��<���$��a[Sx/�i��o\���[�㌩�����3N�I���ޢ��V
��z�|U�q裏C�ه�g��YX�N_�W�Q}�⺼����K{�����ݻ�Sy�"t��IX|��3���{3I�3+���$/~x�-�q�g��c�;���	<nV�׸�F�7�b(�*�5����XUT���2���Yz(��ֱ�S�3����W���<���J���Z��e��x\��9Y�pb��":��^j��݌�R�ݑd��畈۹��t�	�j��@�;�X�ӻ':i���|=�;��{���p�	��q/w�	�l�X�qvH��P�Pn����K�u����E��/E�!�#<�~�w�t�ݏ�՞^�w/A��㬍*�(���dx��hV車7��m;�T�)�P���ä'	ۊ�`U�>�V����ө��A��� ���"˾�˚�P=۰2)���iX(��H�c�$j�-�q�[�	jʹ�O�UM�弼���mW��'(���� t�A�_	�a�Od2g��Yox9mm?AFY�#�Y��^^ϰ��2�=М-]�b�H�����I�sw��O\b�S�m�_(V����̭R:u�Xj�fB��x*$\zi��3(�s��R$5�K��]�:��{/a��`��NK�UG��]�r'u(�s�������dmD�7=Qۙ�5.}��۹�����q�og�Oc�%.|<���^φm�_��C����w���]+:��Y�C�΁�� y�#��V��}��77�u��t�q���mPY��/��]()��OE��7(q8.�Uv��¶h� ���:�V�e�]nU�@����r����
!����h|
`��QA������>�.7}��k3���ys�
qvA|�ΟNcC�_ۜAgX�|�1#>oW__�ݮ���&�=-<��"Y�*Zv�wwqL��3¡����+�d�dˣ:�������@�bFe��ܭ����<\�Ր���;�v'X2�E�%[�^u�ͺ�?=�y�����_^=��?vz��n�U������4�؞���B��������UE�������/����~���|������?��A�4���S�����}��&�6x6�g����.̚���T��9��eI��ӊ�WU62W�����
sԁ��Q��.���INK	��J�gcL���[+���oD�$"�SF�fv�q#��Zq���*�u?��"��%�UH����PSor�K��&��J������
�����kW��0���&��ҧ��n�����;%J;Ӎ�#N	�7�nY�5�i�z���z`��s������2��^n�p���]+q��ʅcճ���d���S�W-�bz�iﳁ���c�VqrP՚Y�A��_�"�H0C�ps��r�S�f��=���h}�e7=�%?Ir��+3ۢu�����ֻ��.�5�--��|ҳ-��������S�1�2Z�
uN�#�n��C7��.��,�䆲@e�'���3kFZAtj�y��5��^���iǙ��p���Ժ�uc���������I��
j�\���&&�U֬r�<�P��$yR�ҩ�'/+�>�#��N�!Ӿ�Tou��y���Dr������z��*V�j��w�hf��2�pE��K0]��F��i��<�n Gjͫ�4�8��� ��ne��X���Uvh�UdS8	��g�[��6�=6:	��7�aO>�*�z���<��At��LRA�����$�wof�yIv��f�ս٣*,�Zw�#
�fq��5OϟC|Wo�x�����n���E�����6�L)���j�zYs2{B��g�iI�IE'm�o?����#�"�M%D��ߜ�c%J��ۅ�����6W+,��\�3Wc����������rB�(33C�+?�e)e�l��B5(��[b�zZ<~?����l\ ��lnq�I��f�m��tUZֵkZi��loF�-/+��3-J�n0�
{��x88<��q��N�N�U�SE\��CP�7�=H�>����Q�Ea)hQ��fa��;K4i�7�7�Y�U���L�������ʳ{-�C�ff�	O;O+'BU��t)�;���xFX^QG���n���>vF����<��*&щ���YazAE|Þ���TUp��)�(�d�&x��������^�MUW)��DO1��E.rh��D�{-Z�<nEVa�ԚQ�hf�)����_� ��3d�)F/*��U^d�"��4p^�L�fq���ݚ�*���糬��tge��dK�wjY�U��y6m��$�B%��b36n�Rl/'�����M�wV�{pwٱD�b����'�x����#X1���ϟ���x)�{���6����y:r�H��U/{iۯ~a��
���`>���]('`颰���Eb��+ ���x׆��ip���W��p{��Kn�Zf�Q�0���tp�������Բ�<wL���`���Gj���h/`�M��yT�R�۞U7=�7ްvzM����!���]c�B���2�J�篪�����̒xt�=�w�<�
&��0�~���%�XiLof�N����z�(��=.~�7���~�k��5A��e��p���)#��4�1v��*�<�AD�e��rǾ����qo�=�~�}<'�/�sC<³�[}�_������{&�N���R/j�gc��2k81�����[��:��:���vT�Z�.'�85q���p]c9��.��\��C�CG[��k���M
�w^���j�����[�.��W0u�:�\�=r��R���/��h��e��u��Z\�*宕�[�f:�t�38��z��B�DoAK6�hX<��}��/Vե��t^�_z+G�W�.��dx*w�t|!C��~٫9{¢5�U�����P��m��a~�ᜑ��{�'���!�B6����|�A��+*�53+Ue_w�����÷��^V�@s\y������{�;�j�e-�d�\~W�Yܲ(iC�u|'v�}wJ��.$=��[��>��}��,�}H�����)�f2�����`���j�X�!{���w,�
�,�B���&�ܽ߼_����?\~�J{��_��I
���\��Avg[YF��W�||%ũg������m�{t��{^��G���냳�_����|�P��7�給�k���]J:�ݦi,�YEdu��rU��$A���Q~�ٜ3ϲxYXo��;�^�:9i�u$P3h���a{�����ٛ�_���a4�����ͦ9��\�2�3؁�A٬+�Z\ɜ����\�q����x��	V�iQ�a�ݩ-��Y�.a-���X��q����ŴTԝU�y%qWMz0��O^�_�|�j�� F��\�?L.���I�0}HM���~��6/�� 勖�%t�]�.��Ǿ�WIW*ʾ����[�z���~��0�1�����b����|p	�ɻMJ��-��l{�v{��?�����0f��݈v�7���t�n��D�Ox%����\ǭ	�Z�o�����m�`a��9d/LY���M~�[����tt�*v�E�([��)���ǿ�[��b��� �����]Oʧ��ye}���R��.;X3�r�����&�|T.�U�׾H���ŵ=�'�z�jQ���g���b���qt)I�1ʗ$7������`�ZsB�5������<�{"T��w�hC�:L.�~ɉ^Sp�3���z~�P�����%��"?O�}{�f}$/�()����R����RFR������~�5�`�w���_~��6��_߷���6�Z�����#w.���{���J���bށʷ�E]r�ֵE��X}[[.�&�Na*���I�Y�M��n^t�K�zU�AF�n#����+U��`^{x�]�C�If�����	7ѴU��lK��r�Y*���ɈT�q��J�֗)Շ������ǩǦc��'��~�"uE��4��^����N�v������Ü��ڞBz��$/a6�/X����y*�͉�}&��/w�Bû��]��.kBc�v����4�F��~��[ߟi�k]y��Q�o�~��m��.2��
�pW�v�3�֒$����mDn��謫GQ&��A�8nB�� ��+:���>㈫�~�u7��;�mZ$��w���x�~�N�"+07��{D�5d����\���\ϵ�tq��w�˵z�zL���!�lx���o-{���?��ѷރ+qw����f|R7�.�T�n�7�_�@��	�J>{����\�'S�Iy{�F�!�����ĥow�yvNe%3�@sN~�Eb���K��M,_� ���*�My�^����9G����{6P��6&�A�F�>t{(ЇηY��,�ƭ��s��0���_�Q`i`�h��(�61X��3�6�l�tC}w/���P�9&��^�p&��[�Bʹ����X]NR�ێ�+�ݯx�#�e]�j	�FTv`��Y�h�F�M���M�U͙����W1[f������`����U��2K�?H�wG�_�3�w^�\��'�὞ږ���������N�7�O��*f�K}�~�kB��C��:1XY&� h5A5;�ߤ�c�+�_����jN~���������eb�3m_VJ���F�?`Jc;�G~���ڧ�e��4�_�V��;�힥kr�$z,{�8U�ߺ���f�z=�K-W��v���_X'�>q�V�
p{���6����7W�'�"J�І�G�k�є/"xvQ�6�`KDgQu�!���zz׍K���G�����k�����ݿ��M���:���D+�GoX�~����1�K�FG.�ݥ��R�]��J��)���rvǽ"�BR�����*�X���k�e�}����q�y�G�&%�g���{ɖ�ɂ��?�a���gG��Ca~-�:�1������4�C�(M)��w��X��B;����ѳ�S��M�Y�`���tU37||�W�^j2��cn���rE��k{�n�N�ƈoo4Ҍ�.�\�r��ϲڞ����:ӯV��or]�wF��Ǡ����>?l/4��t��]ޓ5,[js7��w�<؞�<�~46*V(?g�,�*�	|�,Q)�#w�	3ٓ�&t�"�d��7���=��\����cS�.{��G��^�����,~��5�Y��ɾ������=&���:'n�E�E+��Wv}��N
���+���t`r�!y�W�=�>��/yL���Ξ,�D$��"{���~�G���RP�%pCҊ�ߖ<H ����Z?^#�}����xq���,r�D2c�Q�����DW������T��M��������nr
���l�B�*���j~>C�k`�x5�"�gY�ś���'m�{��es�����4�����o��4���Mt��ـ��xeZ�6 ���=�P�����ݽ�$!�nȀv��3�=�g�:�wc32�.�9U��z��7ۚ{��aǇ����_���jۂw��:��05�̌t�xe+��^)���L���N
7�F��s,���k��5���:�̗뙙���<�o�wYU�"��Yx�ze>���J��ċ�]�p�|<�rU�/aT��۫��}�k�T6`��5�9�
ݍ�.��$&\�c8%Vۨ:J��Cֵu����60 ���t���|���:�2���`rɝ��7�αޝ����{zx,��G�Qc�e�O���BH���{bs�t�u�(A�����.�+�ۿ�օ->����V{���{��y���U�jdr�|uM��P�<<��'L���ro�{X�Ko_��Ø�D�E{�)��~Y�ϳ�"�;���}�+�d�8^4��z.��!���XQ�:���t#��+�7a
�o��=��j���'�5�Ud��0~˝ַzQ��\u���g��5�7Zޛ&��O�?K��x/�������)m�<ԛw�&X�������9Azpxٗ�b���WUK�� Y׽��/�¼��.[��跂������ѹ��Q�&Cz|�{3�}�;���>H��(�]`�6�W�P(j;Ư.yA��*6����C{sY[�B��+�I�[oleԫ:��t����g��v���T�۹6�л��f9�l[�._Uw=g�;�*�e�����3{�K-/�����JNF}ɝ����j��mMZs�<���azf�@����yp�/;�*R>s���6���&������L��rCb!��ix��X�+�sW�y����a��P��s�ެ�6Gv�p7 �{|'m���Sy�c,_{ZY��jG�,�
l!��f#��/�ޭ��!8mi1��:C�5)��7�v�9:��϶��V�١*wm`�Գ�,_�����J�ם�5sgo|=��(%����Fslm����������Y��X}�O�e��s��i��w�v��K�Ez��^���oTV�����X��<�����=���k`������ihn,����>�v�G���� ⶟Z�{!�<���<:H^��{L�RK�2�τu��f� ��z�r3f�Jz�����0Wi��@I�u�o��GT�RW�VLu�vIX�v���5�7u*�����/c��n��'��K��yG���ұ�Z/�����������vxG!�3��e?'�6�n��ohk7��ҭP�k�����)������N=Cx��X$Bi>��@�IT�׫����̼��ìpٱ���Hm� �gq��v�7g����}�e��eL��ٕՄ5�hs�U�y�:ՒD���z��RÈ�D����T
�������Ҹ��pU(9�R���9yi7y�e]�U잛��pg���k���B5���xQi�k�������9�{"�����^�yvNJG��g�95Dym{w�g	���;�!CO�Q��{��z�ƣ�ޓ��ŮU�(�׍��{���}�Rַ �3|7E+�,z�4V�����þ�$0&���zAz�m/:�.zu�!�ᎪZ��D(t_�����`6#���M����2�r�����!i ��:1_VI�ϴ�0�;>g0�e�<�c{��"�)��,���;EY	I3m_VJ��^�#]����g�RN��]Gj�nm����ޞ�����1�=�s�#q�7��w��J^�:���A�BՂ|,t�x��:A��-V�k�e���S���'�ߠ^�7SA�z�&:mQ���<�!{��8=�[V���x7L�$�[:�\���w�m/3�m���{�XÆ�3���wr�N��DMKs�j��5v�w�o{=�����w1aҤ�zz&��Qb�I�i��ΕR������]BD��1���T�"܎/	EO��������o����>�~<Ƌ&�ؾ����`��=�xwZK#�_�� X�g���c��;��4���^����c]�5�lu����*ǽ?P#hJ]}pDH�*'�����~r�]j�FnvOk�"���V���M����Ab#�(�V�%vޏe�x�W |������1\�p���v�V�8�Y��{Ȏ��C]�P�c�3�S�O;���`��-Σsڂ��*;|=g�3M��X��q��{6d��}=��D����tm�n2w5Wfe�z�w����+k!W}p�8Б�Bv=���Y�Y�+Qn>5Oc}��U�s߹��=n<M,@īzX6�j����~�ݛ7<��P���45�{�����q�>z�Q({����(�Ǖ�U��/����=��>�p�3�B��3�O��n�E�ߜ�ʿQ���<�
�_Z��{�-���|��8Hx��wSL]�Q�����w Ou�>�k3�Pd |q:4\) �ʹ���7i��i49�-���^vV8e�j��wɨ�.�˂�D{j�0W1L�7W�PT�S'/���2�.Czs����>�}��Xmzv�3\��2��V!%�W4÷	��ͧB.L�
ޛU�N��Gڨw3�N��G�;:�#���uZ�e���"s�8�y����\�kۼ��u���gͬ:�{r@>��{8G�|wʂvg7Tb��yLM�)��Q��zS���Ãp��S��R�W����97B2 ��W=���HW�u+/�'����y'P\��J�Q����8X{ٽ���h2���'��Ce�<��qN��CHڮ����I��:h�NY�jswJ� j����D^S�`�����@���qչV�e�W�����F�G�l��^�-+m�����A��[4��}t����oK�AR����7*����:� �+�@�~86�&�^�!e'���ܖ�@^�l�2�|Y�W�G/�r�#v�ܼ�Sl�pp�欋��C�s��SS"���avSYP�tl3���:�#�{+>�ft���^~.h�F�;����<s9P}ۖ���{�4A��==���H"��}�	�����D�������"M���9�*Wxo���\={��r�ǖH�<�>M������p?��W9'�"�s?�G��hn��h	�������WOU7AU���|�q
�����aRAb7[�8̴����A��)�9u��&2E>9������m3�6%���$���7��@�~Δ\ou�:.��_ma�R���:�L�:��%�ǻ��K
&�J·T���]�.4�-)��l�)��bs�O�&}؊��zr�|�q�/xZB��4&�<��{���`8���}��5MX�Y�9�Y��!tЊe��c���
�ؘYW�Sǲ�������eGz�q�۬P�mm3y���	k��<�b����ǿ�<�^����%{X��fG�_�9�gU�:���Ǥ��=ۢ�����nTz�I-��ŝ�Cݮ*�<�.��ַ�JĖ�1������=W�����^�noc�+���ۚQ���'�ϡ7wnewJ�r�,2&X�&ULnθ!���Y�;i�k�֍o[D�H��ug�]��{�-�2�1D=�;ud�g����\��m�bF���k۠[۬�0sF��v;f�םn��k7h��ƭ����f�9�֌�r�N�	��T��d�0o;ᖸ�U|���<V�X�q�p�ZMAx8�\vDutGi��#'	��x���z�=�����3>��whf����:!��m��u}G�]j��n��Qg',�͘�LNA���cr)��y���Y9��֮L�k~���:u6�[޷Q7��f����&��6f�\pf9/%���޼a����E������(xP�c�b�v�B��J8C���)W��>���G
����\\n�A-�ӑ��u��`�Uj��^|��q{ĦM�h0z�*�{����1�����*�{�;G߮��*�`6�{lj/r��{֔�S[u�媣8�鶶��M��-q�����������A�0ه�����>�N�\EG���PHZy썦�	w�<�r�O�
��e��.x��j�7Rs[-Yj3{���#y���n>>??�C�d��Oٷ�aQެ֭Σ5i���2Ƞ��h�3,C��_�u���Qm�o�f�����"Ә冇F��i�=:�=�?z���\�%�*|�>�iӨ}������o��?{x����=m��ݩ�s�s��hG�G��m���rL�df�0�����j�ٛ��	��(і�9�m��#z�kOlヷZ
�>k��f��y���a'����@�y=��IUI*����y6Z�}��:�m���hhd�Ջ�L��F�G�{÷�<ȁ��a��y��uDh$�ѧ�w��m�x��څ�v���gϖ�)�������|m�����2L��_7da�>�o��6��֢��4옵�Z޴j��խvs��3<���n�R��	��f�ki؊�LF����kj���Y�kȋzs��w|/_J��]�<��6�RF�պu���}�T�9���ӽ�V��L�UΡ�?Ǖ7"#>	�,4���#g���nV�j�d(Y�^��~��~+������C���.U��s�����j�������>��Am�=d���e��d�϶�����ԡX�,����<�몟�*뽆[���@�!�V{�
.mP�\z�y-�/s���I�}W�Z���77����B�}�R�����)ߠ6o�>��B�zb�/�oⳁ�4�>�oM�tUWW�+��s+�c��
�x��Z~Uk��!�]��M���!)�46E�.w��;5���#�bUp��	��!����ņ��VW�R��c>O��ad�����^��ϕ���rL�:]Xc�q�&��r�i��ld<	�q��Q�1��,���Lo*k�GUK�k4���H��D騍a�\�v�n�X�� ��Ф��V3��J��������Uy��ن�W����^�H_P�B���dA=[��;���N>78Uk����l%>�/�f�k(��Y~�Q�R�=w�):}������@Ⱦ��ft� �<���T����Jv���I�fTlz�S���c�:��f�æ��!��x.�<�Z���jE�K�!�duhK�󨶁k�߯�U�'����$��ʐKΣb��	L�ݽӥq�0-������9�a��n�N�[יDq��I�s ��=��L0�1��?�>����ϦASS1�𾊁l@�f�aɀ��2�,����1�_���b-��z{j��/�W1�97�b��B�'#,?�/����G������̛�S8�ڋ�P�6y�x���8���\�F���7Ђ��~��
�`٨?p��{)=�މ���]��yuXlt�UOA3��B������\��S�b�3�'X��a�:&G�&+���7z�D��59􆢝��b�R�WvX�l�$�|��%V� 3	R��y�W���'3j2�".B-|-KO�a�`p@3���������v׳_��%���a�9�"|��
g%�o�ȿ��?n}���7ʹKO��`��yF'�(N��S�3o�;�Y��}�\�W��rΉ�U�`om�MW�����T~8��x�ߐ��&�9C�x{�:�N����$��ۤ;�͌j�s��,9�?P�x�Ή�Ggр{+jVȈ�á�'�ZS�S�Hأݛ�ǽaa�l����΃�ͷ:%ׄJS��i���^c���r4[R�V,h��9��5��ϗ��Yh3/�
$�ζ����O{A�[VH����|�o�-߻�� hݏ�{�2�~C�7�7G���vg.��GFd���+��k�G�y�UZ�tXp^��st�L���ʰl�Q�����b��=�;0 EE0���M�}�L������MЏ�Fȏ;'����˼�r�V5o���=��7���1sP���rd��u�Eף�X"�+'" uJ�/\�����Y8���S@8Oxz��9������H��=���xҿ)ɟl��40�z.�'�, �P�x���,��t����4�7��H�f3C���Ar�!�@ŀ�͎�o�&�|$N�|ć�0�>9_c�q{���~�{h��۲�O��?S3p~ն�����Mu�3�Gl��!���	p�����}�+��~�$G��{{����B�z�<���V�@�'��F�y�'�+����h'�P����U��E�R�ZO���1�v��d�Övx5�} �l΄�)ا-H!��ce{��x/�uq�v^yF�U�0N� ?��1"<�x�}��(3��H&��j���ϼR��_���O#�+�0Q<ǡ��C�s�Ӣ%�
���
���d�v�߇������7��V$!�kM��yP�(����R�혀�ި�Ӆ]�A�����Y^Pj�1���O���<�U���{��z�vr�ϰw3�mt���+>@�������z�x�W�i%(}�|��,�d�@S"���I�1�u�n�X1ƳuJg2�[�Ѷ3�o�
ΥV�5��X�5m�چ豋��� ��7��ګ���z�\u���/ٝ�ߎ���G�d�)�� `�K���@���{�oB6��>��CşXT{I��i���J�0y��ߐ77�!�����nn}�g�u)�Ր�Q���M���TÜ�=��4�豵쟜a�ږf�Nnw�`����Ɵ�jot��=����>+\�}"���rF(���g~�!����ݮ�>�������<��͝���}���^8o���4#~w�n��>1�P�Е��s��)�lS;�5Y�33?ms�;�O��j4���T!��"П��A�}!>vc>�ŸIZ�_�B��p^�7���[��g����Pg���7Ez��Ξ�Ӝ�g�6 ?NԶ'��] 8�蠂�O��-�W�s1���R��.&f������?O���r�� �� `�Xdd��9�蠦#f\�<��=��в�VC7ZpV}�wJa��c�,/��<���j_��C���8�~��/W�R �h*:��r�Y�P�bx�cJ�^'d[��W
T'��#��_ΤY^xnsUk�	ʄ�ک1�EȘ~��]N,�^���ǫXl@��E���D��/�u�p\��I������۰L��zQ�ʬ���u}6$�b�՜��,f�N��C��ڭL��=�U{ՑMs�����r�u]�-�[S�Kf�G��p�p���|��̣F����i���1����W��駾���Qd�NR�ϡ����~]��4U�}B�h7y��)�Gۼq����}��9��>�H��B$�wc}��1,-�6vD��	I��@40EЗ�``ܬ�zb�����:|��gv���2�Κ��{�1�gn_ُO\��T���@AC�0��{� �Q��>���Ӏ���3�W�#.<�ћ���ֽ
�~��:��	�����,�k���>��`��������@��M^S;s��#�e�w��;���㵎6S�b#�zғB��В�B�Y��c%F��S
��s3A�0�;�j&3��K����!�Hb�ߔ�ݕ�ұ	wg�:�J��H5�?zf�yF��}���y�|E��W�LE�iŊ������\;�\Ev�P7�j�H�1.j���ڈ;���2Z���of��se1a�~���X�/H��-�;����'ty[�c�P"�r
)����5Q,���/����P����X�y�Y����[_Yo$zC{��gû�S�PLռ��Q�����0kW�w������9b��ze�#O�\���{�p�r��N7�8���q59R����R�����nw�<�͇Z�����3�;�#�J��F}S���,Ѕ��M� ��L*��AwŲ�7(���9�ĵM�0�;���f���'�	��z���_1���\�6SDĚC�oH��D�����i�:%D궡=���r;����4�ڰw$Z�g���k*���j�e1��<u������x�]o�:�^�=��B�
Ĉ'>H�ҟu���_��@���,�F`�9n~S4�6ld<	�q��v�g��ږ����Χj�8x�_1��b�o臀vh�$K�n`;�[�m�r~
��D>� ��v�7������*2fr��L)�Sl
�
���N;>� �=~�S���>��pnpZ��'�b�Uv|:���b%����|��}W��=߿��B>|`k��"lp���VJ=c��g��*Nl���]>'=�s��L���W��r��$;�4�xQ��X�D�7S�9+�e��b�d�m�fp�{;������^��eZr�|���oF;��R���'f�
����#Y>�	9�k`g�ٝ���QCh����<�ni�D����� j�:���3M}��A�ͱ��v�x���_��Qb�G��ݕ
{�I]m�Iʼ�ӊ�u�>Ϝ���Σ^��'z&��w����j&�
q0��*E������6 �w�
J�O��s
YX��vr��S�[٬r��E�9�nof�>�*gP������b��{���v�&�>��'����9��l;V#�+��R�T4���f�F����'<��[���EG�9Rj��^VR�A�8��5o:�_7�S�C��S ��1Ծ��t[o�NU˔�1CU4�J��NA��e���рP�j���c%ï��U�(�/��h˰����i�v_0.��m��~��R X� ���ϯ9�]���ko�1���6�)]E���s�opU���l]�8	�����?yX����O�zǇ�}�T����0��� `�LC�Om�^��J��g�τ[S�$�y�����)�E��V���_m+K{��N��ۏ����i�=��0��p�5�^|��c)�^���'o�޵�����f��v�'���G�5�ƞ?��b�)�->X=�8m�#מ��(WV��ɻ���G�xSc�c�T�#�u�s;�0E�[�e�rUU�zX�ʙ�ʟ`�zl�����R��];� �9�l�WE��ċ�8}sA�\x�6���ySRa��.��]��1W�lf8��
+ߩ^�ɡ^ٸPa��L 䟎XAN.�p���T�6���mw5<V��[��u1�/�sJ�����T[�6;��j"bL�H��b��R�>�w׷���|=W�XsD������:���l�Ƭ���w������|�D���b�,:�]�g��_�3�����5���>�X�����~Uk�n�!�(k�l���_�w�g+A}�֞�9^*�x�_\�'7qbs�I�ͩ����A�3���3��(cr�����o�Y^g9=�T�L���jf8E5��C"�xQ�����?��F�� ��v�0��cKFWW)��1(N�٫5a��q�ڪQm���o*Ԉ��]7�Q�}π}�x���u�C� D��H s���z�-�1?bL+'�E�4��9��c�+�uo��)6��y61��=yMH��^	��s�βDd����3�Q(_�+�`ҏ���Jϯ�a�|{��C�y�C�1��2�Z�ib1�Za�CƇ�����W��D�0�O��B��v���G��@q���O�2	�n�;ܫ����0�w�J���\+aa�e��Q'�� ɡ�/�]_ſ�!n=Y�U_���ն79�"��@��ky�6��b,��Z𭇆�f��6	C��-x���O������N�y��ͳ:3+oձ�/���ؚ�ԅ�3��W�d�˂n���������/wo����K���E�����)��(`]�+�<�Vgo쪆�+����_��yb��t��H���������k��e�T�dI���S�;�Fc߼.!���\�%q��%a��nR�7>�B�u��C�R��M��;`�ߺs�9�Qc'bc�AVŀ�Z���6/����|�����G0	�;2p�w�#S����/Bt-@q����ջ?{�=�86|��b�}�X#�߾-�۹D��Qʃ���m˘+��"b��}a�ꓕ�r����age��}��A�:�";yF��%��q�����@ĭ�E����u���4���/8�'�b�C��֟�/g�s=e����=�R]Y�=��7{�Q�]����N�W�8�뎳��>}�@�*Ĩ?}=�>���up�0�}m]�/�M\7/�5��V�5�F	ݺs�=,*���j#�G.�ʽ�7���O���R_E
\���ϫ��5,t�%��Y*7�"�_z���ῳ2��5�DyWߐWPb��)CÖ,]��v:������Z����(Xͪ�3��V���O�ͤW*�c�Mt�N|���!]>�r�e���u�5'j��v=�Z�^-E�U`���Y|��Q�oC��ʇ��p���h��z~#���WPڔw�1F�ߝ���ꫯOT����}�EK�)۝�F-n\Ga��&�6 D��x>�_�����&{��V����F�R����C�9=�%_N|Uلi���Q���	\<�z�P^y��ڥқ�c���j>=�zW���Rs��GX�ԝM}hN���V}k�d(â��W2�YTy1�� !��F����}�*�����җ������J���WQ�<6~�})}}����>�opk��|-z�`��5g��x�xq��c��"+4ڀxo��C#ؒ�|��N���סP:6�=���g��� ��KJ��)M��J�ow���뒛Lx����(�ɜ;Uv��k*8�ؙ՚��b˾�Cd�;6b�v�&��U��k�(P�uUN�;�Fa[;���Ļ�b~ݹ�E�_u�����9����"A� � ��K��Bb1�H��c����������Qqx ���t]Wd�Fe�f{�Y���#�������j�����.�F+�;����{�AVl��I�����,����Yu_Y-�6�*m�X�s+<��M�\f�U���!f;S�!��x�~x���s�Ve'埭b_��	���4`�{"ͩ�����/���_���^8c>�L9U\7:W��[X�f{gc�v%�<I����}���5�u��ub��^x�<�EҀ�xN0֔��V�9��U[����x�����������b���Ǵ��J`�b(_�;��υ/\AÖD<�`5�u#Î<n|VX���L���_Dɭϵoqk:�/�Ӳ>�_����X�-�����/�ddh[���)u���N�w�n����\Z�(�����Ǜ;���Br�M��H_#�M�!��|��ׇ!�ܬud��h^��+bR���k�Z�g5��q���ǡT��!��D��z�Q��eT4��9+Ygw$a������fln_m��ձ�Omи�v�ѺM�*4y�[7n��˸�g[�W]j.&��O����������$���qYj�;�ޚ�0i��.��lf�̫��l�p[����f+�����(��WG�C�f-����h�f*��
N��9��K+o����&>����u	I����{�wh����k��q�M~�B�����]O}ve5ov��7>YZ�9�7�ϼ{���	T��*��b�r��� !6��Ȫb,�@��i�>��&�k��i��n��!{�*��_#d)�A�q�+���j��ih�v5F���;*������S�\�%*"�oR&�@F��B�Dj�����ϷO�ʣ��$y:��5r�>a	�w9^YW�M{>ͽ�͆t�'��^*��Z��j�v�. �d��e�5����*�Е2���|��{3�ϭ4�������w�1���vWp��@;qXk�D.���pV�m⾮�˅�qk5(o��$����S��SL�Gj��#�z�]{����w\�%�z����U8�~a�^�qw���<���kWp\��iSF�V��ZKpf�]F��Yv�6���`cN��gɓ��mM�{Jg�G|�7�^�+���rtM�o�y����s�������Ӿ��L���Y���P���yg9�.�y�^�rfNA.ce����DQ��LW�Q����v]6��k.h<'j�/�"�`�&:��+�A��Hvރ��`��Ժ�{6ʭe��#a\V��S�S[����-�(-r�3�Q�}k��;�0utj�!�g��h��!�˒��Q�༶{3QG��R�Tćc�	7UM���~�O�R���祻��:z�'Ep��9�r`�9�/8<���q��.�۶0�N�l�7�QԳF�k�
�v`Ӊ8��y6-�ܯ�i�.g��3:�]ʩ��2fglBE�Ys$X�=҅�<��.��Em�cy����C)�b��q��鋇v7�
ÝΪ!|ay����b�E���&�xrՊ뤠�����[0�]Qcς�J��L�Su�u>A{�N��f�[��Q�I��IVf�{=h�8��D`���;ZlP���}L�p�z�V2�ٔ�f�w�ᶙ=�y�Czs��1S�D�"_M;�M5/m�ݟG;��	.�v-�{`�&Q�d�ܻY�J���5����O����s��;b���TL7~��d^�E5���|�wT����t�)$�Z	x+�������G���h���Mj������r�Ld�3w��N�pZ�fJ5'ZC3��2J�r*%�M�C�ڂ�>r_U�jEl�,��2�u�:佢a{�@�f��:o_%Wp<�%o��r��Yϋg���u����k<��_��2���t�\;֭aJ;Z_5U�܎gYgq��(�Y�k{��6�5�Wn��Hr#���-؅�)��t��86�G�n�X�sI�0�3P�2���|٪ؾM_��:4)4�W�\�ڧ�v�}Y�q���lK�����.n���1jp�#��7%���a����ݿ�����S���9ȩ�C�(ʡi�V�1��&D�}�z��م4�K��$XV���U���Qx1-�C3ҧ+�E$�������&�!�k�(�6O�ؚK�)��QБgr<�Σ<��d���n��0��5�??���w[-E~r">q��,)������}튻��ey��@�ױҺEo�:�A`X�����~�? O|�L�RL��TQJ�$WS4H��ȥSEЊd��l���05�����~�W�
��D�2��ȿ�dY���DEE�a��H�4�*�$��K
�3܏7@���e�	�I�D��YCb�K=�쪨���=ICR�
�����BʏDK�J�4�#r�!CB0�։b�]s+/��^��~�;��L���{3P�� ������H܍J�WW��	5״�������S��{4�47���.jUY$����U�i�DVk6�u��֝��Z4kM"dE̅P�ɝ��>_G=1A��CDʉ'̎��������QVBI$���l����yJ.��I�&^^�sBET��4,�Z�V�)��.c�����\}���4�t(�0�ǟK����sk2��0<���;��r�[tJ*�g�����ָ��o[�=�H@1��ڶ|��wt!�O�:R�s
{�Vz[�p)��ӭ�ڬ1�):$xA�3��Ex?l0��W�f8��>��+�%F���0�����cr��y�qa�:�ں(w��/*�i��b1����	�ɔƇ�E����M}�ٵ�zN3aw���LLU��u>���s<y�a���C"}��ʹKO��`�?��QC�щ�n_�_��Q5�����5��_�ԫ�b�\E04�9����b04�0Z�*���O�6
I�<ă�����Sӻ�V�;Ez��jk��/���Y���I���pB{|�	�188����@C�������a�=�L/54�����]K3������՛	��o�0������
�ϣ=��+�:}7}fަ�z=4s���Sxu`xU�G���ŎW��^�g$��:�r���=y�Dأ��X��{z�EB4%�v��� |>~��G���ȏ	�>�$ӆ�~UV�������Y���T���ô�n����Ȥkc� ��!Cc�?W�dGA��g��Y�lNo����1ɛ���������vӳM�u[�z��'ims6-�r��@�l��P��3��q���ܪa��(�$ସ��v���.ݎ�[� پ�r-1�������.�<x��LmQh�abqɻ]W݆.��\�u�'w{9�����@1*E� @������$�M�Q��t{�G�-��e`Z+�8&}�P/����߅JN���y%t��sa{��7�oKU7LzG*,/e�9�{K
A��@{�r'��e��!��O�C�,vG>��=�gmxA�`nV):��1j�p3����5m�7�ڄ�]@�53_T�{B�G�~�ڳ�d�^����]�^��ٔ�,bJ�t�Г�>���{�<��	�S�ٚ������F�_�K�$M1*2��*	��^,'��eվ�T}%:V�c/9�m���(�Le���ͺ��WC�Ή�*'�+�u��	���� �\�Cq�b}����vF�?n3kp]s*~`#S�0� �|�S�Έ�j����*C�����쌟�|��a�a��O�}=�fzo�y��8�y���S��.�*�hv}_��_�j�?�1'�9�V�����wW�k_k^�����r P��X��M���t�i]E�
�y��f�`�Z؅M�SڽӞ��^��� +�4\d`�O��|�W�����Q�U0�>Ol1�4���ײ\p�r�K�N�F�kD9W��z�g��;�m�kr_+%VM�E�7O9�e:Iз���T�ِ8x�R��}��/��{��F=����l��]���\��a��6�j�gB�<n���m�͓�,�W[1/+�p���[\�p���λ�x�<[狭�����)��@�>���y)&�g5�&���JP�8�����L�r멉��=
R�5�pci�3�)��Û�)Z��VK~A|/�K������|�7EOh<���~���.g�P��ẇ��~��!_�Sߖw�+|���sb��,q�5xr&( kb#$O�]]��"i(�=+��خwI�$�̕��pe4�wX��̴oz.�P�/���|'l#�Z�c�ȓ�#�������'-D�5(t�&��$�Ƕ���=��������8�u^��9��"|�,[��u6}X����ڗ� �C��*|�d�΁Y}q�Tl���}�E��H��uDz,W
0p�{-]��b�s�q�C	҅b��b����^/L�
=ϟʫ/{���k�Ј'���C�P%GE��E���,��~��r��Iٹ±����ܛWټ���;o=�9��-NH����A��C��켎{v�!�w��b�GvM,��I��5��&u:K�۝�F�Dw���&͈ �A?���h����Y�x�~W��^=����Dd���W�o^���v�{�UV��u��ۋ�-Dr�FzD����Ipq�d먫Nh��bi����ݽ�B[�n��i�Ȍ����$�i�W75ٙ��݋��G�Nw�su�:�4q�s���u��)�X������ |�5H�������|����ㅮh��%�a��f(b5qJ��AG����.v��tϘ�x�Ͼ��p-�u6���I��b#��ڒ�~�$��}���\+!F��ٟi���rȉN��3�52�	� �*�ꞹޖ�X!X��	���*(!i,������t/o^K��N�}�7(��<}�{j�p�'�ƌ�ߌ+_|��w�����쪷�=BP]Y����:���{��������ʿR�:YT,>0�|�*���S��CrK7�ϸL<z�=���֛����dC���
4&�	ϣ�t�Xe'�����/�����w�M�gӯ�3�������U ��_V}a�-Ǵ%lC�~W�t<W�0#[�φ�V��牛�!W�}����'i���
��Y���<�O꠼&���0
��d�`9U\7:>M^C�k^�����ȗ?~�3[3h���A2Xdj6�W|+(�g�A>�g��-ς��/~f�C���}��~0�˝��os�Dd�p��Ԝ��@�F��wGgݖD5�0�u!�7>
��D��SN���qd�OLt;�	%=��v��HƯ]b��hd8U
81��oF�7�wr#�h8�q�W�-�3eJ�/i�s���UO��N��y���[�8�,���������od�h}�7K�^G����cMS*��aN��L`����n�qz<s�}w�w��ﾋř�޳���$R R B$@O<���;�����=	���pg�ה������"��a����)��ˤ$�ǯюW:������V6�uW�=�&2َ�c�[�߃�	@���7����^�'��D]R��t�35�.�i��>�ʃ��%G��P������7�v:N���� ګ��5��P7�	&vrm�%����9�h�8�<��Rt<���+Y����nTy�Y6��/~���O�R@רx6��/��N�fVQk�t�u��o�2L�9Pg�]�d:� �����7�Z�1�Nh���ԆUN��F�=ϼ�ps�A�l!JX����sǕ�$.��-r� w����DA7�kq��z�O#K�p}���XH0<�O��_�<�`q���;,t7��f�]傶��\V�_,�}��m�"?;��=�ߕR��l'�*(F.����/��+��&2n{7���P���=�숤����!m+�����8f�igXɟ"��@[�5T�ь��ɇ��l]�x�����^f��=�>��g�6$j�!��=�#j�'��|=CJ�NT����OW�-�>2�����9�ʧ%��>�w�:oF�v�MɆ��������n�MU}�+vϥ����#�)3bN�+�������'&�q/�w��;�ڗ��:M�n�od��:�p1��9�+ž>k=�;Ծ��h&��f�=4��}/���{���� $�F$ �U��~�y�{�B�|�Ꟛ�TE	.��uf�Rz4ySq�����tNGg�h]슚�J�z���}�骓�"AP��E[�캡f�;�q��jrM1Ҕ��Zo�SVE8�H����Ιo"��C���*VN�Зs�q�M�X�\����I���Aڪ���گ���k>�g�{o��]~�V�3^��!;Rؑc�����옱ٕ�J�����L-+J��:����9�4&s��,�k��T�L�;�5��<	[��H�p��d�1å����ϟ�T_��m�YKb��6;�/��a�J�^Ʈ��F�C1V7�����3e����w6er�`ū������f����;P��ʀ�fb%Dd�L�e���1��d�ժn`A��I��T&�̾Y��T]#Rv�c��6�ǝ�����1ޝ�=�Dk�'��vD�"�OA��b�*p��c���#���} �
M�-817=QM\��<�W�	��;��t��ta�O�ʿ��(!_DHC(�П9Y���>�ؠ�S1ӣK�c��b�^�mH�+�<IgX���6���ٕ�ux�O����5�Tf<�*��U�<�h�(Źh���"����.��q�fo��U��m��6���᪭͐SL�c�t}{�����A�Ȱ۲�a�Iq�)�~���B  T����<�y͹��[�ޞ��Jf+�V\�X�/{=I�ao�������-����/�wH���q����\�~Y�Ά����S�W���U�E����c�*p��c�/b=��˥#vf�~KǏo�왊�0��AD�@>�jD�HKr�Һ�^���MB��~����uV�z3��i�hR�V���+N�lwN�z�Q�M �{a�igё��ڊ\	�<�U_h�¾�V~�q�Y^tV`f�NxF��T�ٕѝ�{2�c���HT�=y��/3����
��v��PT�� �鯫]�|���h>������u��+�v��t�fo+�Q����0��s���Ѝ���6j,d�LS
�,9���6#J^j��N�z��Q��a�q�R�(�r�v�2���R�v����|�(!��I�c���[�$�R�	��]:s����X&�~
j�~�Y5n�D^�'޺r��rg��{׳t�8���4l�c��
�;hB��-�^�S`��ˀ]�R��o��R�"=Bi2,j������6�2κ���Tp�:�Dr�N�7}��
-�S�h��T���*w[A3++����9DH�A��[7��u���/���h���x̊���ox9�y������y=�qܰI�	�h�UM­��^��w�|o����QbPbbQ }���������D3�H��uDz/��E�;�a��{-�.�R3��s�qɃCe��ٹU~}�8�7�.�>��5��~���?��_0>OP�C6e�������6�K�������~��zDO���g�)W��/�r��4�	��~������W�(f�S1s皊�wǯ��aFٝN����tb]Bv�����c����ٛj��f���?/c������T�U�p�4r{BW���Tc�ۈX�DL+T"$��5K�31�Y�9�)�c¼��!Y3�;�eB���0L���QQ?RW���V1�9���-��S����ϸ���5�\�}�\
	�4�T�vW�[J�%ݞ���>'�'E������4��;�},V{7�.���X����K�U�c���>��TX~�UӼW�ޡ��1LE[��	^^��+��<���&�@��,xo>h*�^_�u��
c�~�s���,������!����Z�R��_l0;�	؎�LC`���Mv	��s�7�4��|�2}�y��q�3j�ON����&���ޞ������|n�e�v��:)�k���y��y�xX����A�?M�m=��J�.��xz�J\�owL�9k7x���`iʆh���w��}ڥ��m���tg����ޝM܂�C8aɨcp��Z�e<l��z�Zտb!�X�!V�����~g���������V}X��;�[��s�⾁���sg6iNǦO��X�fFS�c��q^>��?
��p�]A����I��U�s���{���6g�v;�#`�����;�ij$��ٛG�U���]8�K���ќjܷ>UV��62�#�
���2N;�۳�Q>�pa�{j#�Vܮ�k頪#b黈��!����/[�m�s�0I=6n'2���E^,���rpm�{L���'������_Є�9�<:}��O�߿����Fe���U3�C�_��tZ�5�S`�f���	?N�Z]R�����MK����=5c+�<��cso#�>8cWSShk���S�d�>�ML��P2iʟ���lT���^�q�v]Lt��0b�����g�t�nTo���{�����#�:�f#��ƻq�B����M�r�8�D��Sb��&��}�kߝ[�s�5C���m��U�<�z����׸�Ƀ^;��c�'�3Lzè<%���D�G�����'B>�%u�!85p8I��3j�����j��k�Ƴ���ל\6�L���d+|��Q���׉.�4�P���:Keś�Tǭ��D����:vV��ޠ�Vum���z�2t
v��r��G����'�3A�^d�ز*��G2�čB��sf�G2"3mRy��k�u���}��Z�~���H�>� > D}�����a8��-�g˅��� �2�.(�������rĎ��|N�c��yL42�ύfqFz���zo�u0���R,.�LVM,I�������}�R$��č�Uv��F9O>W��]�W�&Ҙn�ar��2��W)i��m����&wַ���$dHw������>�sC��u��w3o�z;�=ੱ#5S�<�!3^�_{�a�ޡ�.b��e���Cz�KHz�L���I3�zr]턷��f�s��h��H�}�k:'�	�1v�?��X�V�.�����t�	�b���eM����Y��M1ӡ*�/+��+���/Mm�um|���uU�����6������[ ^?�^d�_|�ȏ���+���:0���O;<�S�ǲX5_Y��5�^�������0,V�< ߣ갅z.��"��!��	i�*���93�����S��Gዮ�N7�<?Kq!F7�9��X��=�϶j�ޡI��V�߳��sf�-�=����X@�>���ϗ�TY�[s�VC_Kb������3bL��p| �WNeB�3��a�g^&�)�:��m�r�ki_p�)��Y��eM3�����D�2����=����"�;K��^�V�v��@%��8�V��>&P�l���[���#m�X�jՕ��K��R���]Ώt���;}v�7}�))����O�(��v?�����n7�\0�!d��z�:��ܙ��;%[��
ӕK��{j�ǈ����vq���]�r��qɉ%�̐v�I��O���x�
���%��@O����tv��"^�ktMe����H��ۊ܆�h�9���^��|L�v�x�0!�M����
�I�WKYĲ2�8��U�b�sw5���&[�����ͽ�7��q���g\L=�{q�1�w�sf&��V��e����U1fX��.<���ݳW����u4��,9���.�n�jj��{�I���ɬ�+�ι	i�@�n��7��2;BI��l��N�:��gH�B��EFBV������FN"���fR9U��!��.�Lb��v'&^��xM��]�3����n��c
��׳Ÿ�\�ƛٙ I�~qKABS�uIh�MX[��t��5$�{�/��)A��1�S޾=��)�����C�`�|�d`��W}��})͗:�Y��9TÁǙ����/����5Ɗw'�7������4⢹s�~��h�i�}^��Cii�9�e,`�ާ���t;X�V�l�7̥�����rs��bFp�D�V"�ո,��A���I��>��8�����������xg�9.d���t[�{#sw���:v0��6T�R��l�L�\�{k�.��Δ���?aU�:ǝ��LFg��'�M��]�l�m��4vi󎃬�0<�=��C�����.;l�2ϗ]D�x��r�1�to�![��٣Vpc�洣�#�F��}=Q2�l[�B��;���4�3l�R�*e�C�edr��+#�`hN"��n�I�vU�P�o�t}ZB��|��|�4u�%�h�ԋM��Eۘ7�\dO]�#>ՕB��*��;)�M���oS��5Ga�Sw�4,��.\3�w0y	�r���7_��)�z�Z��"kw����:�M��5��11��L��3A�ʩ����~�|�RŲt^��^r9��܌C��u#w���xE�����R��]�=�P�2��i.w�����}Aa���k�u�>{2Z��-�ġe�2:�� �P˺�͸��UNF�ٛ���w�:]/��&���߶I��aB�Rz3i��<҃�^�h���b��Uu�#�����Hiv��Y� ��!�3��ջ������?L�����O���bG�6���T��>������vݓ&��S�:��!�o������K�w��b�:��sq��E7���0��+�����}�Φ��#�ݱy�	�h/\gH�p��Ŏ��Ra�/��UQR>>><~?������59����E���x׻�[t���H*�^G���f�ix{�~����l$���W�>��R||||~?vu�GlY�]�e�߽���f-�Eޮ�>"�`�m)����������e�Q?VUO�w�}C��w$�K�|��|�cv��ޅ�]�U��MBQ>I�	���>>><~?�RɰG�w�<k�
��T^�^D�h�8����H/���zn��£R��{�*����i���R��/z�)ޅ}�}�{���:On}���s�跓^pW�1%�v��B�"��,��z�=��]v�l#2��̧ͮ�]{��DD�8a3r��OS��vQ_;k�=Ny��Qc�T>�W{B;X�1 ��'_A(��sf���f�kZ�a�f�I��[��}���R/L���cơ����UՇ��G�|�ٛӼ����fi�5���ѕ���E=�H�(kɶ��r�������{�J��#	L"Oz����L���X�0���.��5�sF#�_z+�7�q���S5�x����i���|�t���ш���L���d���=� D�� �"������o>y�Ǟ�y�գ�7�ɣ����D'8H�R�X����l��j�noBv�c]�F�z<�����%����Q���;5.o����bJ�k��g�iSK�3�I⁀k6a�2��"g�=��b)dJ�&09�C�@�`��8 OA�\?�c�;˫} �NlᄽY3�'Y�����R�k���_OB���Ƃ]�s.�)�+DW���Yѕ�!	�D�ĵ��Fx
���:�/���t�U1}��1�>S�%XV.f�T&�
p=�4&H����o��Ǵ�)��D�ɸ�.�(	M)�J�N|U�.���[�Sc�VT�t�	�R��8]�
axO�/�Sj}:��qvq	����Kr��T �l=O�����M���R�x����ZER��A}�
W��������z���RBj3�4��ol1٥z'��]-O�gE{3�$FK��y>���mI�tS�b��� �W�����P�#��fV�g�6�]M-����=��^�oL"~��j�_��p���ȸi}j��u���2����C�mec�|z�9]�70RU6�J����Өe�K�����Z����v2d�i�E�O,*�s��A�|o�*M�\���5p��<���Y��˽�Tś��忤����f�9:���4dMªg9�ֺ�:�k/�,�x��¨{%�X�%�&��Q}uתK�i�M5����Xp�����enǺf��V�� �?,9��'�dҌr��y>�{�]��G�� �Ɯ�����ʱn������@q-;;[�����͏���g�2�mEgth9������%
�A�}�|��&�~SW���xX�`�Xd5K��}�fr�8cd���`�R��PDz�g�B.��/��˫���ڗ����N4Z��f��Σ����ԽH����T_��8g���z�����.�K�ԋZ�{/SJr�Vnc�л-�DA�ga��0-L�Ϝ��40��s�B�韟��mJ��Ǫa/�F�*��l�W�?Vqc�u����&]�ǀ���-NH�����W@7�B��H��3��x����W�M�i:M���~�Q�];�H�3��SCbtc�ܸ��vt�$8s��=�#���N]������-�c��eE�u0}=�Y��ㅡ��ԯ��*��v�*���u�Q=�*x�r�b!��	��r�6g�tvT)8;�Du�[Rw�5��9�QAv�>L;�h.��Rt����p�fzlyW�����Wy����ߌ6p�T���ԭ�KUo�:�s��Sh#�!���3�����x߳�޳?kR]����ڹ���K5C�w�|��d]P����r̅�;��m�f.E�GU;�B�"�C��]&�^E �$4���/�@H�Ba� �Pb��I�[5؊bje�c��T����k�%���O���ީ��^�o�%��ݞ�1d�Bm���Y��z<�2eLT1c�\~�~:)~�n��L��~0φ?՟�:&�#�A��Zڿ��+WRŗ}|��Ev��zo�<orᆩT��V9�7�Qc��tI��aӋ�^�F#z��_c����^�[��7��0�Dv��>b��
ɾ��+�Z�~���3B�| d7d�z:A�v�c[/�|Wn��X�__��zz/�>�K���!�|���U��o�>�͚S��fM�+�}%v���S��X8^@�����b"�0�}&�r1*�nu5y~���߳&���U�yl�c)0�����N��2<f��o]8Ϣ���22�ۖ�ʪܲ4����m؄܋��zLT����x�cE�>��Fp@�aTG��7q>9dC�����n�^�|d�fD�;{����7G:��j��~n�>� �%^S��� V����!.;~� ��.�t�C쨊w�x�ݵ	K��?IVK?_�K�l%8ʛ��*�V���}�ϯ\�"G��s'��y�`��ΰ����[qC�z`3�J��:V#ғw��p�UXlf;]�H4��R����^�tW�񣢰n���Vy�~:$VΟp6y�}�s=���u�e�x!Zϖ�w�
��UCmrTU]�ʝm)ټx����s���Z�}�>�Y��H�!bA(Aiy�ή���L�#��up���=yO<1�[Sx5��u8�g s�l*���^��i����K�ݳ�%�"X���:��Lt��0a��,d,V�o��&ۗ�@ػu��Yw��gw��'F�(�����阌���%@B��T�KS��3�*�2[�p)�}��4��|����ʁ���{�{KQ}g�Z���~������,��>��54�G����-�0�ʏu��T�0��A�'Xc��������OC�>~1��/XڃO�e����D^鎛���qshGK��=ߢ�u�lw�>0{��=�ߕ�Z~��$�*+�чENz1n��C�uy����_���l��_m���M����a�ϚWQ��~+��8ߴ<��)=�TF�
��'����	�E'k`�+�w��ω����M����8��lFj�'=װ�oM
�嚲�ɳ��){����e���<	>0YH��3;�h��_���~J�r�"����^�-��v�v�q;IB����aȩ����%b�����9�C��S�k$��c:sjk�V1w���r�W�]Ć���-ZV�29�Ϊ={�vfv�4�����~R���SW�t�{�
,��)ɫH0.����R�D���?;�Jw@��9d9̠[��e��ĉ���J�.e�4�Тf�J�M�V����Kb�D[�:)�{�=�>��P"Tb~�3��[}�v}�6�d���8���5�u;k��������7R	���Ԙ"p��9w�����I/x�ئb�ɣeLӖSX5��19�
���b� o��|,!^��Ď�s��/����Y9��sn`������ǎ��ߠ��8�X��<&}�P,w�`���Ymn���3|N���t�p3�����TY�[s�U�5_�P1`�S�h�xgMέ�*-DϺ�ڋ�|�Mˑ>�"A麒 �Õ�R��k�c�������m�����B���f��y��>����;��2>��%��5� ��!q���(*M͙��m�Ԧ��g$�@�7MI��[�W�}U����%n��l2 D�=�	�1!N �P9`�V1�Iޯ���ݕ{��y��!?����NR����>�Кx�K��!p�C�_�ϗ��
M���d9����g�nc��i�� Ʋ��85~�T�����21O|��`�&��v�-����Wd[���]x�9�����Rɨ��w�@JiLw�\B��U�18ȯC��lK��	�z�`�a�}�����Ʈ�k�Oy�}����#?yN݈�)�C�>�IeSS\}7��*���=�J�Gs��Y�{{U�ḏze�к�A�I9ΖWG�rMO� �M�寓�����t2��v'KNB::fV��d���/=[����5�4��;.x�|���(��(�)B�Q �(�(%
'��r�|��8���`���3��4u���'"{ըO�M���1WQ}��T��¤(��[�~'H���u��_0J<ğ��+�̯�YT�U��xg��$&���
u���wF��{�MD�߂f}_��R�C���\见��a}��<,��xk�Fh���s�>�#�n]�W^|��_�TD<׸1�x�B��0�q�^�tW�|p���!r>�o��A���q����n6�A���(bR�ڕ�5��^/`�F�Ӏzsf��v&)�[+3/�o�����;�/�lf��t��`�Y��ŸZչiҀ�}M<�W�ޜ��M93�<Z��Y��iNE��/�Oߠ#j�2��}qQ`>Y��vܿ)����A����8	���'�u�ޫ;�����C�^������mR�̛�!p]-��{p�ӎ\�-�y�g��ޅ���t5�|FD��k�*|�d�ϦA��9���!F��b�`#T���f�޶:Nʿc�/�/��c�[��S�	�U8�"PF���_u��]��KNΘu?Oշ���{�k%�����om�JZ4��Ar�Woe��֒�͊T�_gOv㱊W��R�u�I���1?1儇ݥ�j�&>�v�v��8�qNN%��y)�빴�c�W�I�x�E�^��I��Y�'"���$��oV���x�g|w�w��2�W�@�J�� �"�	(TB�D �� | �)�����O�g%f���w��x	��9NH��$Pb�� �ʅ�f���w=O7f<�K���y���hK׏:J�I�:Jv�~�>0z������� ����~9��&�m?��~���P��֬�GC_gWާnsG'��T_IUF4v�䞹��~ድ�+��څ�1�(D<�N))��lϔ�eC���`��S%D�HO��]�
�1�S7Q[P��OB��!�&�a��T°p^T�
�R/�yO��񖒱	wg�L^8�gd�;���o�U>�/�)]B���uVT���e?��~�c�Y��]N�_��p��ȱn�˓��b�0���Y��p|��c>j�H��}z��٨�:n&��1p×KT�决ӂ���;
���2��K�VFro"9�[�?^�q���9����zsS��t�U��u��F\E���g�F���M�[__
W�	W��$�n=�+bc�s����N	��u�q����n�ї�Ϧh �{F}�y�!�;�}`���6n�r�����g���R&p'��|�'ڶ�,p�нT
}ä��V((N�[���=Tu&�[�r=�����(�,A��M�n�j�
�;�J���ҥ�@O[7���h�ww|����V��J��I����r��t�R=)�ڪ*�D�[��,�\�K����4b�L������?�_��� �4!@1 �M
�2����׭�w�^=z����3�OҶv?;���ٚ9�1B}��谅�Z3i�s\�E����>�[�wou�^�};�B����_������~��#b黈��vY�.���<�\�995fA���=f�ž����|���~lb��	N��'���Ӱ1��/��8���b�t?%�[|f�~%x�G=7��:�u����*��~���>eI!��Ȟ"+`%��}n����먶�O��{
�
E��������x��=ﳭ���c���tL��9��?X
�d�Sۛ�XfQ�3ٿk�J"C�.Ԍ/���^��2+Y���r��Rɵ���f�����@�t3��>�޴R6P%eO�L��"z~��P��� ��T���W0g�����p	S]�&��B�;��˻w�>_bw��������+B��������ߺ��u�G���}�|B �P^���NB�zi��p�E`���U�����Dȯ��M}LW���]?JCv:�+��'�ܷq���<pA��χ-�o�s
-*U"��Z��d��X��H�|}��tX����_X}W�(vqS�I_P\�z'&��݆���o��e.N���n���B��t�q�Wvz�g����6���f����(:�Ǝ9kwj�~�����k�^s��6r�;��WӉ�=J�0�X�H��w·�n
A�U��7���ky�h�q�:��Z>_d	B��1* "ҢRO�}��(��W3�y�b������;e_{VDVm)����+���c�7�J�ǣݕ��۸#&3�œ�LL��Lp��@N���Ϳ��ug� �Č�LG�}����4�����M��R]_h��7�,�Sʒv9������b�0h���_Vl`.�s��,9�ᔹN[ҁc�W�.�>�U�5��:>��V���}B�%|>a��B9���Ot��q*�퇴龓~�&ѩ�D{�L݃I��=1����~�9[R�o�Dt��9u�.��-��B�"პ����')���C��J�ʙ�,��kט���ׁ�P�v��&*�x<-W�+/�T����u<����~��$FWQd���h8O~�c�e`[J�N	�l�+z�Wlb�wY=��9�Įc��v&��������u���*���*���p�cS`�>�ȩu�G��|��߻K3/�\ɉsbD�RM�*P�gV9J�Ů�v8��-�ȵ��܎s��{{��X+o�g>�W�����ȟ&�/��Q��*���V{��`ՠ*��4Z�2�wsw&"�?��ײCuuϓ{���$��X�핹J�.�K��d9;�:M��_� ��������]�xlA����(����f��;V���<ׄ� ������rM!�q��N=���촬�di�%K������(D44�� D
D% DRJ0�
z�q,g��2���xݙy����	��b��?j�p��.<P���6��z?�U�p���3���m�s�^6G�R�IN����F���`3�d�4 H"��C�����n��u�����=3�^����T����97C:����²�ǹ
���V
��*���&���+�_�kW�)�c½��j���e�(��%w�@��Z����.�4)��\'!mmD�]v��m�${܆0b},d��pt.�(��a`���?{7��B�߂u��Bq�D0ǵH�I�o<�"2UC�vr�r�?V�J���$�;�1��U�:7_�31��3�|~����k��Sz���&��;�a� �����T������� X_|�wr������ܣ�m�+���T��Q����g�X��,Zm�������T�YLS���t�U~EJ����y����w��_kϩ�ǹ �N7�Cɩ�r�m���t�YUi�J�>Ӱl�����ͭ�ϴ���`W	U#�@g��g]��%�p��5n^����SO�z��`�>�7�_J�c��?Y��y�/��C�WԸ�z5�:/:���j{��#�'K_7�s�`Z�Uz�ds�f�;{	O��L�Ⱦϵt&�X�d���c|A�[�Vؖ�����iTK\��I�P,(6��]�,�S3V�+Ef��ӧ��l��a�j+�Ս�r���n,Lٵ�B�W���q�b����ٸ{<�Z8ηV�
'��^SQ��IӼ��؎Λu"��9�t������η=|���2�i��u�,�2V�vi�s�	`Tb.���{ݣP�݃��|��$�b�YTP��iQ���R��܋r�;(4xJ�n�F<ܔ9V��g�3�ˑ��]��*V��Ol�H3�>���IȻl*�M�j_e7�]ޕY�����M�ɥ�t{ǰ��D� ��Zr�w�>
�ݬ�y���*��u��2���R��Tͫ��]I2��tCUs�`[x��w�ݘo7ͫZ�̴�G2^l�q1w�����������t��Gd�����{��˱�1:�+x��S��2ys���I���۹��9��=_�6��Ɯ(�He�Vz�n!�Q�-�\u��;�;���c4�:P�;�v�s�e����3��|*�ù�͋�;.��NA��/�_]��HEEz�UK!ո�]5s;1[�ɦ
p��ToS�{�0V��mʷ[��Vj��+�pְp�h��$�c���p�k�Y�}2,�oxo'l-v�V�A=ƶ*UhJ:�do-7`�*Nf�����]0�͂i�v���K���y8��&�����^r��)�ܧ���A�����x�x��;*�9��i�]�-��U����y�%'�]w������;�l�(6���*�;jYv6���$S���y�/�4�}׏���q�����;D/6c�J���/�!�}��{�eΏ^�g;a�Q�VC(np͡��^�'=�b�8������b}��<t���{q���.��w��od���W=�_��4H�� �j�7�a�c�f�W�������/�M:R��(*Ɂu,f̥�S�����Ɋ���%�9JAK���N	�֘���;�J�d�K��o��1;���R�k�m�f�Z���x��3�zt���V-yH��d��E�P<��=[ڷ�U�/EM�rl�e�ٛ�5����ekL�M8hξ\�]70���i6��I�e*�#�Vc
해{���om��B��3E��I��'�G_Rj��}����G�S���м�9u!܋�xk�q=��"*�����/Ъ�D��3o���r��Zm�8�]����nӻ������0)�ϒH���'l���+�4�����w |�zI�j� X� �X�1��oj3y�~�uhy;����t�#���2;knvIz���ɚ��r�����=��9"���M.,��NX�mu�j��<�M�G�^7!��p��~l9#����B-M����k;k�m庌0�%q�G�$NJ!�6�u�FaVE��ٻ����b)[��'�r��\ⷼ��-�0�(�����a�g�E���O�ɨ&M�>%�5P�F0z�>�ţw�ۥ���-���6ۑ�N���<|~=~|Es�z]^Y�4si��~��Ｚ�Q{�3��W������)��ڦoF<�4MD|||x��?�Ğ�t#Fض�£#M(���=�=���(��-ӶG�7������9�~>#�������/��"B�QQ�]�j�]���֍��c
�&����*K�����"�ǭ�O90�����'��T(=W�`��M�!Z޼ak��Ũh�9v��{��$P5�<��{�2y��4�>��ԋ�͵�P�z�aN�˭o���Rp�^���h��l��#עϕ���(l���S�5yô�gR��7��s�g���y;ۗ�lڔ=<��=t1vfE=}��3g��3u�9;����F#���y���{�U>6�@m]�l��7&��[7�x�g	��n���!g�Z�����״��G��v|�*�8oH�%]FM�j�t�+z�������]������vJ"���;����K�l�O���i�Š�hټ��JBB2ġB�HD$��D}���+��i��JmO�fh@��9lO��9ρ�PB�>Y�5M�Q5Jpk4K���;2n���3Q=N�?���]�ʀ��Ks' o�}ʺ�!�=�b�/c��}X���܄��C,!�P�&��Qs��gX�Y�*Uʎ":hH���O�G�E88rÅ�{�L���21+���>x����竰���&5:P�3j��9"h.�=`��ten��E�������Yǵ���R����{/�c��7BO�k�eތx	��8��T���A��=#�_*�C�.��v���P����^A[��Q��;�H�2��9snz�n\H��[I�Kz�}��wƐ��S�g�
�`v�[��5��Cpnx򽇡��~sG'�%_IU\s-;�{ ��g~�m�׻�iw��*������
�(�ŞW��ߗV�����jN�5��2���%<q/���6�Qk���_:��<s��rs9��W	�un�N���K~JpJQ�|uR��}���.�����f��y�j$!�%�
8d��U�'>�،ؼb�.-��`j��&���~�`=^�t.���R��3t���"�d�>��"�z?Ea�}�h�f�Y����ܶo��T�~�k��꽭S�w#�:NR=��A��V�ӝ��w�v�.N�L��4�rl�qV�.4�e�ژ����u�!�{w[w���/nrËP�ZY�o����b(�$%a�"Qh
V%ZT<�λ���>=k��]��=�`��,���M� op1��T�����T9KL�P�,>0���gB��%E���3�-�t����_��U��97��y[߫ 8�]�s�z�=9�N�Ԕ�1��,����z�_|^ڣ�3ᖳ�߅�g��%q�	[��x�C�~��w������s>���h�E�v��'��d��8`7@F>�S~�<)��0�`J���|$�)yPC��sৰމ���7ذו��tm(��թ��K��}������5:&ȕ��+�u����5Ve�62~�<�\���m}@s�Ǒ6k���N��"��k�Qӄ̝�O*�n`<�ԋG7>
���7C��A��S�,��VE����������[�bsN��w��ބc�tDs�ъt��/��pnp��%��x0%;�a`�@�hI�$��n���,�O��^K�C�p=F.��"����z�	�}W[Sx5��u8�8�� �	Dz���_U׸w���<�1�`L�����?PC3�0�v�b�~yc!�w��yNTo�j�͖u�\Fu�2��q������T��4+��tmLwd8#�~=�oމC��+^��\t�z�;�
3YyG�ʦA��ea�A�z`E�on��mk�{��F
�3��ٳm�ӗ8��*E�ʻU�XqeH�rV��f����uYs�]�ݮ�׎��H�(
D$2�*�-* �@'�z��u�|��k=>���Gl�C��$1&T詎��ʃ=��-~u{ ���v���.���^=ۍ��0T����u�0):'� ��`�P��
���T���7�yqP�JJ�f�_A���Wv/�T���x���S��p��^V��
�X��Fޓ[c�Bp��Jmi������aAzN3~^X/W�c *�ZT�xFAk��zm/�:����;���_�=��N5}�`�"�蚟f�c�(�M�C�ՑM%0�d!4���>�s'�wH7*��bv�f��x���-њ�li,2.� z�������;�w��}|�T�ps�?^��mԫ��[�sD&H����4��Ύ�1�+��$ŏ02�k1Q��������|�����#\�I��ߣ�_ ���_O{�*>/OA�Vԭ��0�m�R=SFcy�C��珲���x��Zp�O��%\ў9��>|�cט�H��}}�������Mb�}N��m���t�h~ۈN�{����1~�������N�UV��M`��ӑ\�dA�쿫��CN���l�����ӆ��n���������fh��l�Wx]��Ha/���1���g�b��ٮ���K��C��G���z��?gj�犄Z�J��ٛ�/UQ�=��lW��f�֤ҕk�{|.�-�v:�����ALK�]���{���}�#	$I �����Pn�/)�A8�S�H�tD,>��"ϳ��Q�n��	��+�W�a��$2 ����[q�>Ɣ���Ca
迪p98XAN.�p�y�E�e�9�^�R�
��mFOX<}������y:��L���L��0#cMԡɹ�+�{ ſ��f �l�П,��5�n%�Dg����2���=j����%�Ʊp��!|z~l|{ʀ�xe��`ճC}��gѲ��k�GՌ�Ǚ��f�?��(��c$Ot��t��ǅN��>W9Ivq���'�]���4�\��~Rm�ߓ��c~����Mr��rp_�b��.ǩ8�����ǝ���V1�:ƅ��.�q@1�.o2�7�:UL_aYpc���*0D��0�������0dv8�=�exx:��&L���e�7/A7mw�}>^s����B}���3�U�^��mbͨ��?'$5��ę�����]��P5>XF�x~�~�C�����+�v�ӹ�1vo��1HX�����;?���ϰk��|1� �'�+N�Y����}۪����f�.AW0��{� �y�.�7�ޜ�Y"�C��¥1ֺ��t�l4'q�7�ܸ׬�w^��&�(qZTje���f�7��wr5����a���0�x�6����}�K���:�p3-��"`��u�M;%uK4\{�Y�r�l��p,@#���BR�@%(ǟ7��^n�x�&Y��TC�Ol1�4�豵��ڗ��٫X��Kr/�ݼS^c�Ny�YY��^N��T}�q���a��$y[�5�{�x�D��~��7z�&�㢴+f�Α^7C���o.��1R+����}���%�q�+�bܐ�-��:�����d���k�uڍL�.��(0)	������>B/��f0Ib�-
jܽN�)��X�g{.,f��R�|~}ڨ��|)ZL�+Wx+�n�
pl�+���;�f%**��_G��
�+~�D��k�<p0I�2#r�,���N%�rؼv�s�I���V���7��^>@��zg 2r�-�:�{6����KĐuXAW��$N|Ǻ0��ozd�/ވu������	i�R-j��z�\�NT%�6�E߃��&��������:hid+
��M�����u����ܼS�����\���\��V��&_�@3�)��&���^�P=�=���]2@� m}=��;/#��q����@��ad���S�;�:1kp��<���O&�j'#4b3���Tq���ʸ�vV�x3X��q��:'E0��o#8�ֻ4+�w�V�S�4jҡ���=��D	mꈞ��N��Ꞹ_]�����Ʃ,%�ۏDoK檭��_���_��"3��۬��������]�|o�y=�z%�(� �* ZJFIJT��o�z�}8���2�aH�%)�Lt����1ޜ��o퇪�8Z�O%_W����t�ǳ�v�x������N��X����0J���2�흅��ۯ���U<�=�'�����쫘���9�L���K�E��U�Z�Y
	�FP����XBK�b�^�ߎW�K6US��pf�J��b9��΁1a*hN��ʋ�O��������^,�~%>j�.����_ݯ 俷+L������<��m@M��_H���s����X鸓Q!��I��&�wwy4�C ы�W�]�}N}޻�Ϲ���V�<װbk�Nu�K#tz�c�.�w��4_�d�!#cDs�����3���7ϭ$-��BV�=�Ҳ5ҝ����S^Sb����9M@c]o�Z�OUX�!���\v �����῭}��h2�x�r`��K=�:�+�����<k���e|�+J!�>s�ǰ]8ϸN2���l����f�ɫ3�}�/~f�C��8��;f2}[S�/��1�M��̝�� �W"��i�Q��M�#�ɥ�| Ws�afu�����=����΁�,n�j�7-������*�מ��zhV>�}K|����Į�3r�N�Ɗ��{T�/]�λ9i�Nt<���x �F�C�{��Y���Y�3B�kӍ������!"F b	�$�}���.I���G~�M��J�{�<n|��)��61pߙۀcU�9���ϭl
�1.�a�C盾'H�a|��[�o��A���b�\�z\����%�A)_qv ��w��t�éQ���|_e�������~k�!�%rέ�@�xcWSSk]��wT�fz��Y]c��ѕi.�U׽��B��/���!�@�����2�,���Z�F���r���z]��^�^�~�6��Ɓ;}�lU�t��T��~��N��d�x�
�.c��Õ=����C�3ö^fc���`�ٯGt�k��-V��蟍�jp�aa�(���5)|S���H<�Ψ�>�;X�g���L���[��h7�8��a�5R��S�dP3Q5�
11w���^�����א���):��E�?��yX�+�0�QS
8%J�O���ʇ)i��oP�Mf͙�$)�K$TR�X��R���d�	��{ڲ"��Jc��#WP��&~�Q�Qӕ�}�W�����i�}$�1 �xA�p��fm��{�=<�#T�.hy�QV_���zfw�������Uogj���2k�x ��3�99��a=1�Я���C0O,͝�u���[j�E�Mˢ
�]�0;a��D0%&$���+c�}2쇣z��o��ceާD���(͇j�	��'�{Q��m�w��޻���AA(����>i��'��=�}��{=CbT���V҃�١��G1Cd�p{�����j�^��>���1dzz�D9��5~����0{+jVȈߘt6�U�ϭ�F���Z�����g�f�����H�0J�!�u*�-�m��ߣ�ڗ�^���R��Wt����.�|{�x�-�����`Z�&�7*f��͌M�'#tW^����b����pꂜ|{��S����[��DC�똯�'��,�x��M	�B�@M<�d�;��dt���]�����X�{5�c`���u,�8r�B
s��.|���>�ns~*��yjU���ޞ��M�����Be��3�o-ޙ�3�6$N�|��>��HA�Õ�R��k�v8fy#����}�ݼ�sv�oq��d������m:P�k��XsS1}S�"}�83!�R~+��[��0�o���?1���Y���P3�هz1�΁�)����6��3�i��OP�����W����,{����#�@Ǜ�[���A!I�g~N��������a�&�4 { �?������ћb�S|߆��Ê�s������Fn�5g79%,���:�ҜO�O��|KWR�Y�����y���Ke��)9�oA��Y�W��S����7��aڧ-��7Ai3N�s�\X_G}��狮\��و"�-+k��9��Q�5�տo���$�h�" � h�>���L��F���I2������0��'&�gV�UL_aYu+},w��ZG������=324�hp�"'��S�ȝB��;+�Q��d�{r�G�����=�T�1i��u��#%�01��� �lJ������|'�f)��Nz��Y({լMl}���Txx�v����c�K��A������g��-3��	��~B �'�-̭����_��׵�b����?��q���4����ˏ��fn'|���E���y��P>��!��Y��SY/2�go�.7D�t�;��z�ž���o�/n��t�M��nT�8Ŝ�	��>���#�<F釽bmCĔ)��V=jŹvv�����!_0�h��y�s�x�ၳ蘤lXr-��]����x;0��c2��-:0d���9N+l�usOwܦ(��"�ޜkq?*�l<j@��<��,�YCÇyg�M�r����DWm���{���]U��zƿ��C��8&���ݺs���-1�V@fp�!b�oc;S����&��ڿ�<��T�V�\
�6G��IV:��dH�U�wS���$��h�O�bX��O��*Մ��8�L��ˉ���g�*su�oW��I+��L	�ŝ_:绡[;Fd��7P��	�N_\wy�ֺ����X�-��L�N�Ɲi�z�׎������"a(d��]k�u�֗O"ߪb���	]5-���**�/��:�
������>�1j]�"Z���gqD�1���b�z�H��������c��N�)Z�R�H�Au	�_�n�B���w��$-��\)BwV����	r��<W9��&]۰L���Qr&��E���Ο�T���OV�!�|g�$��켎z�Q��;���KN������F/��S�{OJ"6J�߅�!o�k�0���$N���h�-�yS����ۓ�S�}�;�{r��8�Y���3��V��W� �Bhp��ղ�^���U$&�g��4�]�m�h��\Fc>����؜	��Ug�
�Q���X��h1.�s��n�建ޕ��c~������3Z~~��}+�}�+��@�RL�'�Q@��$��YDL��j��n���T�1X����ioa�y����K �AW�k�:�����,���j���c�R'}X�W�3�5�v�&�}~�C���پ��E}a߂�Cl�0VWd�̿�N}޲3ѿ�";@�!�V@q�5�&~��N�o+o Ok�[�b6J݁�tgw�x�k����"�@��bZ�,��[�f,�6V����q�c��USW,�o9����}!���j�X6^��lnLn؍�d�[��um#\/�^"�P�\fZ��*�IN�u����IcY0e��Mtf�;m��H��Is(&���)��9��K�&��k���ICn�:�������|R��MGt�c�ΧF�B��Tc�s��wm�]X�rAr���;�S���$�I���藆T:��iw�o�0��M{Y�h����Iz�r@DW�H�7���k/�m�\�Z
�=����e����pf��P�ALD!\)ա�c����lv<G��Č(BpdK�8=����M�2L���3���5�^C��/�*|=M������a��H����<2��s픎wC"	�y�f���>��/�엙Q�3�V��`�u�pn�yޘl��H��HiS���w��I2JG{3{�z/ ����n苅�Q[��u��EwbV�:�F"H�X38�6o/���Z�����W��#=���ݩ���.'�O_t�D�؜2]+��!q��_qe�&���V�Mu���;R�����UY������ӭ%�K���̅u�d8|�x���7dWM;�a_E�N�;��<������t�`D�z�b�q��`��ҽ�؃��A��\���f���3J�;��5IV���n1�?'P��uS5t$P$#'M���Vee\"��JX�"�Rq҄cS<��9�Ь�����ݾ�eLY��R�i�|���� ��幛e*;2�1�v��]����Ga��/t�������T�dڮ��w�?���s����u(XLKWJK�[�0i���%�E�k�ԍ�E�����L�.��5�_+�A�ښ6���q���qq�+�N1��m���qK�,鶁�Y�֗E*n�i�ꓭ4^N�7�wtq	�0P8e'�QO�m.!�4�_9ޛU�gNh�HE�s&O+����}t�O{�V곻w�i��^�TG��9ZTNh�t��*�ɔ&V��6�mǩRRAHNT=,��W���,���>)�5}hMo�'�LWǈ�D�k{�~�s��r��H���ђ�=F��dQ�{��Q'������s�� ���<b�(�w�#�1�F��J��ߐ�Uy-��P�� �'����[;4��PT)���;�EV�-��jPhr�"t��]��E>��;{Trits]M�2�̂����,�(=j���TUk�Uq(z���̦+.�wBq˔�<��-��|ڨ�.=�1VisUU��^��wG4v)��	e:��*eh�NZ��x�k6��z�t�A�K�ݕ~AZXnt�/�=�u^��[7Iv2���xx,���Ã+'`Nk������ܭ��g�4L�w]|qE��"��gP��i���v����z���R+�9���UG��7i�&(0��{���{���ҙ��F�u2�U�1UUoM�zњ4�ekM�����~?����Nh�gZ���ɔ�ϽQ���zP�T��G�{
Y��MfEA�Jz,��E������|~>?	��*'��dh�%�3*d˞h��}�h�C���9E�^5j
��+Z�"�dB�4�9'2�{yD���������x�>U~o�5d�WS��(ȥ�3�h�[�	��C�G����疵���G0��������G�iҌ���)��tTP���2"Ts�T�5���7j��l�K��Q=�A��4�|�s�4C��9+&jS��:(Ra'3�E;�?D"���ē�=��;k�ie�Wh���t��[�n�Z.�zE7jj�g�ɹ�̳PM��(�Rm���%�s�P�H�uĨ=��#ˢ��l�'��
��ģ����y�x{g�d�f$��F����'��В(��",�Hg��v�lc�t79�����9	��GZ��8RQT��)ʢ����gm��g&D�IVGF�4�hùoA�T�Nn��R	����$��"VٴioM�=rfY�.������x�G�י�T��&� �9TH���ji%w{}%�Ԩ=R�fᬦı&l�o�~�(~�> } G�{�˙�7	����9�^��d�xHح�ح�������t�ġN4�B{bҘڔ��� �*�Æ�k)��g�����+�S)_�z�%{������N�PHM�}a�<1�����!�79���jq���W�\��W��q�Uw�~����i8<�A�D�G�1��|~�R}����}�Z�pxo�Rܩ�r����xX�ch��g��ڗ��E2l��o&Z����ɗ����|N�u<	}Sp^�R,qǍϕV9O��Y��06�_���EM��������.~��/!���O
P��B�F9���7��.J��%�C��*��M�#2�������:m�ܪ._@c�����W��JE��W�^�o^D���7Q���}��C�ƱɱۆM�m�2P�y���k���/�C��:rD����fZ,d,
�z77ʃ����v����ܼw9�)�|��ꐜ��]�N�d<�~x�L��0�.�N�����wI��DU���=�7�ޫ�	D�?O|�������3A��M��8Qq����Gty��=�
�d?��v
�/c����WF���V�3���XY�\+������]��3�5?(;y��1}	hv��/��{Ϛ�����N	V���)�,G{���z���4��R4���:&糕�B��q{�S=P�S��Z�~� ��R�Her�g���=���r��`|�I��$�^@ρQ@�|Ua�RFʌ
tL���D�lGC�|�km-J�A�L?W�jO����BZN3~^X/W�cW0��T�E�������Е��^._4�o���,-# �-����� �����^��?1�Ց��Jc��#���skǻ�~���i��8=~��q����s^%��W�P�����3o�:ug��[���'ϯl��m]q��<n�b��.|��Ҩ�g��1�*�r��y�
nlT�Ӑ0]턇�2E��~��ϼ4�URo�I��/��ޢ<(��L9A���6��s�Ggў���+~�á�4U�<���Eg�{���j��:��c:�	�ϯ�L�b�CU�[�b��|E�����xR.�ȿ��^y�?���]q	�1`������1�I�ʙ�,��z����u�	�#A��|3��+�����}B��R��c�šA˘B,+��q���p�4-ϳ�`U{�4��{��OU X�/ʒ�L�����x|��uA�<�{�\5�u�[s��s檪	�qa!��2N��;��+�ݙ	�Q��{�c���o�b�=K�)�DO}M��Vbڒ�'�&Z������7�f*G�7?=Z��s7/�zV�5aOf�vw�\��w���\ł[C��wC����VSwd.�y���jIi՚B������oߦ��$�}qw��<�=c�W�|���#��ͅ�zf�U+�]�E$>��B	�+�${$њ��r��3��{��3��W�n3V�s{�w���m2'�H���"��/�@�������}8�0�vq�7so�s׫_��e��V�F��@Z͘w��Z��:hr��,j��9oS3��k�o��P[�J<����y`סվ�uI�gBt��h����/��)�3�ݵ�8e}3�����O�xc�-2s��\z�sx�7�:UL_aYpb�7'K��7UuP�b\Dd��_�:"yЩ�!К)��b��$��\Crɨ�W{���l��Q��Ƚ�<aMK������d���g�B����TI����hy��,"�\�����Q�3��<��%����������>�OM�b[��pi[3���s��E��`�~�;���=��S�������۵��};it�>��=�,MF�@��04����ˏ|n���5�5��(�.;y�^��<ٻ:}�懆C�o:tfW��2�c ��3;�LC�5�{�x�D��۬��p���Ǆ�i�g��ZO�yҴ���	��	22�y@n�Z0��\�
��Y��|���8X!6{.�����S}����l����"���?dEC:b�d�Y���Q\U(�St��kQq��6V�C�)��]�f�`�ex�����"" ��2�M�Χ
���#��fza���6��K�#�%A�-ס`�:�{�v�t��ş
���{�_{�ێ�3_���0s�!hO�]şg�E��f2L�n��/���rȪ���Gy�w!ץ�W�ޜ��V�&?@�6~?|Q�x|�
^Y�[�5J�d��؏__���ն�O���._��xk�Ma���t磣�Dz�g>9HB��橛�
pF�콉�^o�T]106ǟ����:\�/�k!��>T�TD��rs��!�9�H�%���7^��]���y��
>�[��u#3���5V�1�҅��U&1ȹK����"�78gݦk}��˦C���cp����+~Y�=F�Q��9<W9���z1�&p?P1�W�����^�y���k�vhH�)�v :���}';/#���lF����@ϒ6����S�7;���3L��'�b���חZ���Wa?��a�H���;�����U��}�W�FZ���%����tɔǍ�}8�ٌ��,U�&�B �"o�57S}>S��Os�*{|cc�֒�}�z*΅�ea9�~�x��U3�C�nn�th��]��2�,���n�.<Kk�fl.3����d��4�8�Y�%�1�w]Z
��U�֎5m�U�z�l�XPRq��O2`ʱ����p�h���u�{�{�{�{������O�"=�����M}hIQ!{{ο{B��:�GӜI��hY���5gb'"�z������:ץ�+�K�K+��@��i!%D�9%��?_UeL�yEP���ë������ͯ�`�׫��Klª|w�|�4$���y쪶:b������T����s�f{���^0"�ne��{�>|���)�������\^љY�뽌�Ȏ߼��x�{��;F�(���Fz]��[���b=��W��7��?����!e�^���§Մ�����n=X|�z|xlZӏ�OA�Dz<������v/&��g�-u��®�Cbx���G]L�ȭ���w9/؊3�*��G��HeU�s�5y~�}_XF�7���++�FҸ<�|��84}j����jvr�V�2�:�<�����8$չnT�9k�ld<mc������zr����<�k9��X�q~��<n�"L?��qσ�".���z�H�8���)�B���3��g-&u����o��O��#�gߎ�����С`�~���_���u��s�S�0��H���p�����|OVOjg�k���ǯ-qdVf��;��e�.��$�+�=�9fޟ�ɕ�*v �{��p�/.�uy_ �oRq92��w`���<)���w��l���w�mڣ��Y��<�����`7t�ݜʭ�W�o�Ma��H�~ D� {���,�7Q�R�~]�N���[؀��J=2a�7�p{��1.����O�ީ��Y����T���9q�T���5� c�$���%�fZ,d*ؼ��:o½9��{ʟ�
�J;ʸɇ�l�����R���'`�A^��y@����봈�Ҫ�����^<���g�Ұi�V�Y���C�ԏ���Z�1�):'�L58A��#z�%�;����T�8�Ogǖ	8�7!hU�E�M��$l���D	������N6��r��믁��_�~3�u��4�u��o�;��e�Dx�\G���!3v����rCY/�٣�)�$T}�d�ԧ/��=�����=�YD�S	yk9�׾���5�l�W���_e��⫡�]+����%{��y`�5Q���m�>�L����>�66��&��t�gY�B��!�U�c{lF ���Ͻװ��6%̓9)�� ����F��wڣ>�꓇�T���o���`뾬�Ʃ=<����<MgD�ʎϣ �VԬ�á���r��VbBdXn��U��U��J�wnx��æ���%����2�~Q�V7T�}>�;��e��n����"�����V����۠Q��pɋo{\\WH`�+<7�R���X�g>�|k��}�d:��NgNV�U�S}j�\sw]뷭oY����I�(�����]�}�E���L[83��Գ<$��:�c���n���~�� �mKU���HVr&xj�q{���bX"�}�j#t]s����}Jp�N��U[��5�^������r���i�ٮ��2Q��:أ��ޏ���LH�!��±���c�D�	�L�c�;c�tg&&X����=�y�Gl�P�W��Prp��� C���1QEK^�]}�I3��	�����͎ϑ�3�L��7"v+�$>���&p�c��<Ί��+o�v:!׽όe�a'��X�f�fn3V�siօ)߮�?���A��<AT��~���V�̥]�|k�N�����b���jSK�3�O�Y��tS�'�쉯�D�,����g���O�^�R3_�01��WT���^�V�A�Tq�)NDS���`��Q�>f�Y謿y�}8��3�e��$��ϨO9x,��q�]���\�85~�*�8d��dj���c�=�ź��?���_+d�$�����	5��ˈnY5H]�P6r_�I�8k�2U7�(����.�q��_�g-����[#�r���i�9h�SF%���~T<>�7sqȰ�gָ"T�n�6��w%��!�IV�mXM��r�� ���hQ�f3�#�qňewt|3����.�bX�+O���}��^t�LT�ُ�޸��UUG�g��������|<�г��,(]�?{4\ƫH�䠲����~1?��ؚa	nCѪ��+a�$^zn�hU0ȼ�_x�P/%}.�*߯�O�Cӈ���;s��{�X���M g�g��~0[�_��5�s����fzХ�|��o�mX�P���}ٰ���p[�]Y�Xf|��h{������@�\]JyQ��Km��7hԗ��2)Q��*E��CZ/���	([�jV<Z��\��Sb[���?j*&r�����81U�h�FǇ���	಄c�����:1�p~���'ux�Cwݞ��ռ#�ߧ��ـ� ��������4�}3P!g���`hx|��I4O|�JJѾռ��W���t�5pܿ5��5� ��!J�\*���Ȝ���Gܚ��F���W{&cVM1�<I�p�Ί���U'�n\/-�~�A���>9PqR�Q�'��5�w���;���KsO���6p����|��1j�u#0/<785V�1�:P�mT�p*D���d����?o�¬�͔�nT�C�Kd���Uj�ƭ�A��(ǩ��xŕ(��U��M�_�׸����g�_�낉n��� yS�꽎�?���-��f�ԑ+�	!���p�r�w��D(�!�)һ��c�^_W�����yT&��}��� @�{Ѝ*��}Z���WƠOG��p���v^9z_�(ϗ.��;W+�tL��x	��ap�<R��p��X��Ll=��5����] �g�%t������(�z��6��Y�6�I��4ֳ�������?j�X'nVGd.��8s	�>�4`��#Mft����c�l/�Jχ�#�Y�����Y�t��]�� Gn!b�0�P%�<�z�H�Y�Y�Q�9~�qk���ַ��me�:EC�l/YRuM}hN TSΧY��Ed8Ţ����bT	�^�_�_���ɷ�>ZA�����ҟ�K+��=bɤ��X&��K*-I?X�{r��5=u��@����ŵ�V��\xT�'8V�ux�����"��6�,����5j�Jq��=�QL��w���־�-3>P���V8z�Xh����Y��]�g6���ʾb6��M[�����7��WWo�*�fC��`Tl�U��?����A��/���n �w�צ�������36�4��DN���lB���^9׊�#[�ؼ�R��o���b�("G�r�n���=�~��Vڸ*�����ݭ���4d��g�o
觤v���}��?ni��YxGS{���9��0����1E7_�z_��;�/���q頹8B��-�ʬK4S2,��m����Ն�����1��.�����̩}�t�;�B��z���������]�ս��S�,=�Q�U �`J��M^C�og�]��a��s��;aP�=>��U�g��7�滭��E����,}H�I�r��*�r�3c!�mc��}f2}[R�����缟�����9��bǪ#bx�C7HCAu��N�{�q�s�U�S���l�@1[�)�e��E����y�\�r��_K��V��a+��P��B|{�tk�]T-��s�V�-�8^��C.X�|7�,^K�9�"1��ȓ�V�W�E�R��`u��3�����LC�P6���F����{~��������\�G�&8�c�Cc��F�˽�	���M�Z�v�I���;m����g*L??OZ������Br��H��Yx.!��cc��^5U$mGno?b����*�>x5�έ�8��N�����م�~'L0#s�`�뉸<�1��ZYRĿ�+Т�TyNʅ=�!��'q�\��D��*��|����b�L�S�w~k�܆2&C5_p�)q5/e@���'�/,��^)��s
�������W�]�J{��}�g�pP�v=#$��[={�u'T�a��X"�u3#Ix�R��D�F�a:gB���b�����~�/�/zk
Q���L���<3>�m�ܽ�*�G���y���}[�弩��}�q̶=�g�	5��c��0��3�sy}y�z�IE���������n���Ckwi<�83����LU�X���g:WK���\r���W�&z�'��Ro݃g��Xz�Y���͝�i�u�<@����Vh�-��}0b���%���8� M�d���U�:a�Lh}A��Aųg��r<�Y<�S���OKR��x(�z��z���!P{����eC�Qd��S�g�$���%�[˦�|+<���r�CaY�t\��S[�髪�Fc�E��%�yn�S{��z/�/������
���{���f�v�KjnΤ�j i�]Y�v���R�y�z��Tã�s�7�뤑�w�굘������5N�H��D�/'�u��>�Ţ��Ȁ��� �X/fX�5�Y�x��c���/��f��G��6�:|R�k�Z���N$2[���D箅�3�=�`+&ɜ���c5+���	������.{�s�ٺ�쫰]�>���_iu?�\~�O��Xk�(겵\̺�#��e�Ձ���?�7m�5�1)�I���n�=�H@̩�彠����)֋���A�xU�y���1�%Xr4�����[ޤM�D�WjQ���:#����N���a��;�)�Fm̏���=ya�+휾Gn{�Ű?7b��M��8�W����P�շ���:V���3;8���	�bxPc^*L"
J���Q���M��:_�z�Z̏��jn'/�u��j�4	e�GB���;�e��B.ǳS���[�Iհd5<檙���:�e�Ѫ��{��U��T�j\9��̋!͏gb|v�:�эx󸒓��.MHW���(^���P����s9���w�jn�^7!���d����"a7. �������X�P'���y�J�g���Z=^ITϚ��|x����s<g
��fb��#s�37<�iYg4�/�,�2�w�u#��#r��Gc#�qj������f:�����<��O�'3���*c_��t�:���]96�A�D�C��f-76�U�ͧ(lȵ&-�Z���䴻޹�j��J&qvTމ�vpeQ{�ⶥ�y"8ƊpnۇS�ul>�ԖIL���;��wZ+x�Zq��; �s l31����W���ОZ��-��쏫���^�;سt�����%��M�2�4��r4�Nk}��ܘ�T�kr=˥�V*[�<�ߛ�S�ba{���zxt�{�	�I���׸7�%��z!{�zo����� �nw<��Y9�5�p3;2X����ƥ���G�yӲM���{�^N�[����¿4��	�d��L�E�и��,�r;��O��~���}��C���>����>Wd����)����^�#F\�ی�sM#�<-����9}���a��{P;�OZГ���{6�M�5�Z���;n�+iJ�����}�)��, ��ڽ�ox�]G�������
/�2m'�O27�ƭtd�4�ҳҭB:%{�y0"��i6ɑ��%Fs��܉2�������~�QG�ݵ�/J��
��KB<2ʄT�Tݞ�V��TF�x�fl�3y:�I�������~ꊇ�Y�*e�W<NO��!摐�W����9TI��QQ�� �F5]"��=-2H��4����2�HRj"HW=�D'��7rT(��"��l��t�Ѓ�Y��H�rP�?&{"��� �h��J��mO��dAW�Yo��D!���rɴ�Z:^RXIeQG��K���fF���e�*��%�N��y��g�[���֛V�kӺh�M�jrm6�D��TA���=���͠�H"�R(	��H��
D�h_�ˠ���Vu���"�[�,�-��;�^X-��>qv'M�r��$�DǦ��l��[����-��<w�����E�f��=AD㻖6����G�c���9��XX��Bf*8l�Ϫ�zr�������"+/�20qP��*���x��m���V�����Y�Z~���c�����[���Ff��k5zz�{͘�+P�i!9�@�LC���`M_D���dK�93CB�����=mLG�*�1w����7*����h�Vl`�L9�߼��8�\<	��''c��[R�DCѪv�sY�Y1[��}-
c�_�<���b�_B��S3BM1'�U�=�n�c���kљ�EC�b���Wܮ����עhX�Wʕ�n]71}�"ϭ�"w�p�ꪑn�j�?O����=�kR3�w �N��V�,	gG�0P�~�-��HC^��#���	�n���~س��;*�Z=x��`�8�4
+�W�rg�5��Pa��mJN����*Ǉz������`C��^�ʿ��wD�L���ǝ��,�3�
�����T[�6;7�p��S�
�>ԏ��9�a[傫�4�^$�Ž<ǳ�0��P3>^�f�5m�7�;P��*����>��܉�vt�)��lYa�?��.լ�����>aF������=����Gݨ�������f)r�j�$t���K�^N��,xU;V�vn�{�T�s�\�&*yO�b��6+˫��ݬ��⦮o�Qt�k�WM|��4p�[m��n�=�ޭk^�x�{���!�"A��^n�c^\����	N<�R����~Uk�n��@��ه{�<���=2D����iKNY�v��.>����TY ��X5�uo��I���N����X�Qx��ҷ׳R�]����C��3�� ��"�C�Ĉ��}s�Z�a{���ro:d���;<�.=�y}���s��GC���*±s4B�5
j�d��!�h��'^�p�V��|qI�8O�y�s���AWu��1eyOڢ_ �hy�S冏G��w_��^��{���v��.����&�a!8�!�U¶�����DO��k20�ub��R�w���wO����>� �_��n�#����~����lB�Pc�ig�,m{%�u�/5�71g��?�n�[��1�ʠ���`[�+�9H�,��FG}��L�1>׸1���3�Z�����F�]̜އ�{������"k�)Ǣǅ�_�f7�_C;��\�([�o�Xp���{}�0r�ފ��^SǶ_c����M���nN��|�����x]����{��f�}���\����c橬�U�t+����y%@����b=3��{-����s/��%n|_��{;D�hY�-��<�����"��.ϸ{�6[6u�,�5[cf���������\�l��Z/�V�o_�_�&6�R�ḝ0D7b'D����2��J���<��W=�[9���~;��>b�%��^3S��Mt���Q(�����e�Q7������+G�p|0��E�s8�K���"���޿�j�9~SW�nf����C�N�Ӟ��XU��B#���8UE��i��K`w��Rq�_ĺ�JٿK���j_��C���AR�}LE2�R��|i��O��\tG�p��Q���.�Z�H��y��8��N�,ک1���l�Mˉ������3h��+�@�~_��0��v^9z_�(\�c9'��>�v�auf��\Э���I��3%�T,�;"Nȑ�
��_P�/����>��(�z���<y�C�ו���}�ܽ�eK_��+��=u?����:
9�ǅ3��Nϐ��ү�o��A���e����<���8v�O�+��py,ˌGn!)�ʄD�B�<%�������B�M����kҽ/�P�������'~S_Z�E�,�߰.��;EL+5s7�YX?<$�����߯��}����ѭ3�+�)y,���&=�4���B��.q�����yC�!>�U��yy#:�B�}�ƎJ;�õ�v��cʛöx�RIU�aG$s}�[q4�#��e*�*�i<���`C��D��J����0ev�2�M�57�E��;��N�[d�bWj�����)��ǝ�no��a��[pK�ʹ���
�il���"��@ﻚڶח���j}�W\+���"=J&6���o�W���c��"+�P�yY�G��g�r�ЌuR%���W����)�~0�������/X̿��޻����{ݥ�.b�����rق*�Y���
Mv	�V9�Nl�4.g|$l}@h��v~�4[�B���}t�I�y����g���LC���/���P�x�Z�O��%���08E�� �3���Wt�Z�w	c9�"|l�	4Ñ�U�s�&�!�7EWz}2%ϲvgx��U��ÜO���ј��}�>�g>�V��-���8ؓ�c�S�af=w��PSN0��Z�]?HS��'q�vY�T�|�n�X'7>UX�?A�1�:��Q�k��'VVS���g_�
C���Ԩ,��C�)+�	B�}u�:��c�\�ש����MxG���ߠ�_���c���s�2��8��Гp+`/��mJGT��.���73�3;�1�����zv<戒�;No}V#�ܐ�x�|�� �Ui�0&D�@B�P4~]�gԂ/u���|U�-���@�g�pP���Z��o�~�g����d���2]Ʋ���&B�lk��K�7^ܨ�.�$�Os��W�Y��ll�Qn�����E��s�խ�'o��9̉��v☢9[sv�,vy��Ԓ"�v*��͂������a�Z�z�^8�����1}� ⅶ�%��}���Ǻs�e�����F���r�~�V�n�}�幑��$��.І��D�}b� ��bz/�k�r�rX��:R�yP��+�Ӂ�Mt>�	��U�0):'�8*`����騐�$|�<9��$�8B6%�]
,T���
{><�I�,nB�*� TP<Tَ����|&�q��U�O4�#;Xx}a���
.����q����~{�'����+�0=��]�WfB_W�0f)�\3��E�Ǣs�7�K>�0&��q\6�MKr����v��7�'����5u|:g�D�0�+��So��7{���5���?{`��1'���g�>�.��	���{"���4}>��^��Y0��1#>��q�?c�=����G�+	�z�����>�
��qtS��T�9.��=�͌�L9��<�����\3�oN*[>�{+j^k���JO���U��O߰kA��C*9�0o�C��S3�i�K��J���,�p.#|�_WAwՌ��7�0�If�l��Յ`����̛���0nDxv?�.:������'��Z�6f3|���f4r�_����H�@�c�"�oD��
��Y�g�<�M#��<"+s$�����Og�{��?mA[w<���ǌjqbWf��~�}�'[�>ܜ�筴^J��N���>J�l+w����eZ�GW��x�8x~ ~��#� @x����K΢�������]~�`V�, ߠh�MD�bGu����B,�uqV���ڱJ}9v�#�7�ϣ���c�L�E+�9�϶`T��1>�(9&� ���<�1�^����ک�c����B��s�
�����͎�o��4a�][�#�g}���Q��'{�O���(���%�ص˱�����gڶۛߓS���m6��%�ƭw��,��~�Of��w���1�v��F|��+G- �r�ޑ��O�lý�t{D�Fh\b�0�3s��&�@�!Ap%G�.���;><�k���H;�l΄�)����RS��e�L;�(��Z��H�L�<h����"�?��:L`�>r�_\��֠+����҅UKt������9�EK=S��A���{=I���-�+�omu�B~�|4��c��>7�:csq��qc<��g�yy��w�g����
�奥A�B�^S/���d�w��=�7��Wk^������7��X��l$'��4���¶W�P�������3�t�=l����vA�k��9�w}=�T~�hg!����ct�{ϲ�%����1�Z<�#,H}�0���ު�z���������$�ZN>�{�nO�iU���A�:��Ij]x{ϛc�r�8����{|��t�Ut�y����"�yG4����(��Ys`fV�v=ӱ��$&����A���|ׂߣ��\l�����r=Y��}�VT�=�����|{�����?���H�����3;�LCז-�{�ljT�nq�����w
_? ��� ���
������|�|���6��]��9�t�f(mtu��{茈C#X��Z�˦j�Ui�)YE��yك�'�W���	�_!	�FRCշ��p��c���ں����biJa;Pe4�nׯޜ��M9��υ��'�z�%9�\�9gz���I�C�NtH���ω�nY
j�p ��)�����5�#>�ۧ&:#���W���K�ϡ�s��#�P�>vE`�Sc�Ԩ�,�ezd,�X��J^ݧ
�_����K�"�
�����#�`W
0p�˽����F`^xnsUk��t�Ob�tv��w+6��1�F��hD���/ޢ����z{c���/�b����^+�q�T_�"&L��f�C�gn��R�GC
rD��"��� ��$K�=uqρ�Q��j�k���Q�<'���֬p���&��</|�vv�euC���:u��P>ꮣV���mJwvl��"�J�y�N�{7ݰx붌��.��]ŭ�G�c������-q��[t[�UM�έ.�7+̞�'�l�~�kZ`��[�S;��H������T�w�@������S�6��-�N�g@+�0���Xt":�>}�~�NW���	wm6��^��3���uO�ۄ����	_�Ӏ����B��DL+�P��	��Q �����j����>���g^T#��c�����
��U�j��!}�qcr�[��"ywO��V5�КZ��|ށD�c٪l���L������L*ª=^�<�rAl���0�U��	Z���bЏ�{�D���&O޾��/��F��s���^���_�����|~��������O���q]b�����ema����W`����oZsg�.R�l*ǭ������6/��~����dz���Շ��۞��_�����a���V|�#����Vl0�g&�u�G���o��s��.]��[��"��|9��|���5o)������S��"b��%W5ɑպAg�����E^"��N��h��$��l���m�;�l���z~�ʚ���e0�Y�sͽ�������w��(����9��5���Ov�U�|�z�+s��.\w)��>�=-��C����1R�~sǱ���2<�-0��$�8w�IM���a�n�t��������K����a�߫�pޱs���(g��~���K����;^s_m�ʅ\I���6 ^�^��$L�^�[y_��O_��a��fP$ߧ����{r�Z"t�����O97=���z�{9���XRZ��`�T >�8��q��fk�"���r�(i=��BW���NI�Ϥ��T��|��M�u	m�����$��c;ӕڂ������g�r�ӯ�X���l�~��|Ǽ�^��{I9.(� ���$���O �3�)�ؑ8v���o��P�F����<z3��}qA�N�z��>>Qݩ��M�*B���^���Q�����2qC=a`bb�5_�	T�՟z�7���U�mFL+F,�$� f{��XM%=�#:���~��P�%�k6�t���
�E��]@�59ډ��u��Z-��������]q#B�jS�"�~+�*z��}^�:dp��:yT��}U�I��p���{�9%�@�����hØ;�J����]_��&�HU�Roj��Z��&��p�F�i�Tἒ,�������w9��Ǥ;;.鋎A�y�{-���*7g�^�۠�ǌ]���;m��y�Ӽ�aja���Ƿ�Cϼ�z�>7��H�^uݍ�|�=�{*�<;�v}��<Q����������近����+�����A8�Az�g{���_�=l�@]�@s�g�ﾂ��%�иڀ��~�(ؒtN�οj&bv�b�n�Vlh��Hm�lWl���ɷ��yUyb���-_5ǵ{|����һ���^��!�ln�����Bdo�E��TƮ�.���*����~��� ۴�8$�r��,1�}(3�_?gN]�J	<k�k��L������|��;m�+e(,�p���>���o|>�w�'��ފN!濧���������3W��ɐ�e���Y��
�x��]N�q�ؤ P;��~�ݗ��G�K-��Y������{g�7
p{0�dF�w �rP�Tk�yc�?݁J�w@�7هL����j�M�Z�dc�W~�*��Jt{_���'\Mg��|�w�m�=-%?vf�7\������/�=�g\ݐ+W�<�5ʂ�V��ϡ7���^B�7)m5�n���t3��D�[\@B�oٛ��J�_?^֘�`��Lߥ���V�wP7C�H�紐{�g�����MQ�R�
��^�e��Z���c����=��W������i��\�-��.�W��8XwCz��)�=��+�:�v2��#Wig��9H8s�(Ե�a�uN���Z���5-6��Mv�j�=�{4�Da+z����#J���ZȺ�6��Ps���������&�ps��/j-���^���$��$xY"OCl��7�U�y���վ������E'N8�<��|:�K�u����/�"wk���f�X��@֑c2ESk��-�y��`�i6w9���r%�ˈ�8���v�r[�b]�Oq)<�}��X�8ܨ�ù�پa��x�ޏY0R�)a,�g\}j�Z5��Ԅ4Aʇj�ɾig�u)��s��D�nz[�"كw����=�!F�W�/��o�Ɍ���˜�Y��������1�3��Հ���_����A��{rG�e�v/2<�3��ܥi���
M�S��eZ�Hތ��l*����P�ɹ�f�É����{�hCK[��t���0q��`ŕy�e�m��;B�k���ǵ[Î#t89`��ܬѹ��M�|ڒ�����sr�p�Q���b����n}�uW��F�D��G��
wnO�sA.����u��ja�>�ǒ�l��Y�ʊpQ�?w�Q㸙Y��u���EI�.�6��2^kŲ�s����KΪW,e��+����1=���Mgj��lnK��1�3{g�."�h����c ��6�fWf;�o�A������}$^<�k�T�m7yC��ޘ�'Y���@m���9�t�Ȋ��;tquu�tz�Y�h�lJ�sU�e�]�Z�&��ٌ|nf��h���_���s���3)�ax�f��ڲW��;�4L=���a��V�y�nF�}�t��%b]ٙ<}��s�����]�'�ꎺ�T��8)M�N�K��0�^�n�j�͏ly�wVf;J�f�����=	߄I�{&婑����.��g^�ϓ�_]�ΡL�b�^nb��)����V;Wt����I������[R^�7*�2s	KWl�閅���Wv�sO��짯������)6y��Ń^T��CoEkHMY3���N��o���0K��Jnʻ�ًse�d7%��Z�v��u��x�/	�mD��UT�K�ݝ��1��լ�Ea��@�PS�9P�z�و��Ϊ}\Ь�Ƽ��5�́=q��Uŝ��9j#5��qH�ܣ��@y'�</Y��=v�3w}��Dd]7j]`y[�hm���
Nb�uޫvvE4,M�Z]�d�^y6���a����vj\�s��<8K�ĂHi!�]J�)��n�Q��UTahYEG���P��ݏl��l�����xV�h��zQEI��=�h,�l\ߵ�]��A���*I���F>?����IFLBL���m9a�H���������v�J�n�è�C�������Ea%i��J.nbU�.5
����K�,7J�%+�~�2K8���|~?J��~�*�����IOb���z��!Y"���G]	��	��Õ��Psr��E�fJ��UyzzW�a ����_F�]t",���b^�˺h�Q�JRDj$�YXy$�0�llЈ��N�T�������*'�.��̏�
)4�B&A(^��
`v�9ܨ�4vҊ

"(��6��jRe�bT�.U4d��J+E�=;�eq��TPyZ�J!{-Ъ�,��ETR)EDi �jQY:U�ɞʈ�D/�L�	X���@�@_�?��H��k�ۤn^��\}�NH&�2��6ٜsA�CS�W.���/Q9�1�
�&,�8���o�����N\�9i��})�b�����b�����pA��p0�������G!0L�1�"�ޛ��7>������3�<�b�
���Q#����$K*���|k��^��v�aռ:�>��+Bʅ�O�\1X/g�����^�~5�Q)� ���O��S� �]�X	H6Xh�����ѷ�}g������(�5��>? Ļ	�=ޚ37p��w��ЛP���B�D����xs��:}��FQ˛�A\H�Ά�	��ְ]����n�Ǜl��v�dt�4����r��;���^\
}�4��L�������xo�_s��䫖�&i/L�����4��kV�;[�������y�0������
��Q��O<li�+Ы��T�2y��U����yM<ɡ����e��4,�=�t����o	��{��P���A������M<{h��p؍�p�1&�`�������*=��v5�����o:�v��w,9�Ƞ�}�������K��.�VE�v��X��|�����L�&\Op���|Y�����pb��|g9����.��H�7��.=9��84\�J�^\!'C�����J�q����cDdU�p��5���d߆�2���~�џ~>i�8�����k��e�M�6�����{ζ�-{N�5y��Dd�_C�BI=�HG��x��ל���Xqs��\gYk�'�^w�H���-���A���di��Io�L�%�����V�z{��^�ו�Hor��u�f���>�,q� q�$>=U�Gz�r�}��5
os�����-�y��q4���Q���&��H1? V|���׹�#*6�+��3��v�� T��=~ωw�U�
�X �*\uj�ɋ��3���̡B!h�t�����8��I�0�]Ep��y�Y�Rkf��~����D1��u��Ճ�|ނA��O�% T/��'K��=<*�B2e|-v�%���u_1������#����&*�%纽��
�\�w�����k)�}���VJ����V/��u>��f���ŷr0c|��uö�z~�4[���,�i5HV��k�^�K1��O
X5h*�y������ĬU�m��|udO*�f���f�O�WNbT�0d�J��S�i3wu�����n�l������H��_���%�J,U�}:��&DLTNUQ�<f�
�����4��n7����cڹ{�\N��ap�ӯGMz|�Tt��׷�����������d0�<��z��:����j�^Djq�p������^�(
n{�/|?	���iSg�չj��e����wz0z�_r���͉��P�e4��G�>f��m`3IbO͕��\j�'2u����G�����w$��mKb�D}�Y�|M���Oa�rc��yw��̻_G�_��)j�ޚ�1������ �>��o�Z}q��2:'����:��v�ҫ�e���h�!�?t��[���P6C�JVgw����lՏ/2Mf{�oXï��Y��t�$3頦(GlkÏ!,�Η�����<��"�&�YXm��T�-��ܪ�����
q��:�������R|�Wʇ:T�����mI�
y�D٤���y�[���耠*�ʺ˅s�4�����3�*�����t��Xg!�����-s~ܲ�j��|J=�޸ �f���}'t�Uv;��Z�z}�4�Q�6F'&�H���V���q6�͸����Rcu�~f�g��7}ن}=9��Dd���j������|��>�|�Ʀ�|��������ΑUa���FE����F�=��<����m���#&�v<�W�mvq�=5��Τ�|
S@.��*�C
lz�i���?Ez�;�������6����7����m)�����e�"<s*�DW��
���wE�,�υ�n`����&�������L���˅�ٝQq^?���h�h�������̧�zN}^��M���~ӿDu�"&�}z3�2��2KW9`���-��S��(kֲ�͈(=Ě�R��ɞ#�yzc��������}f�o#F���C�=�E��vgf�}�易��_�,&�Y�81E�i����ｲ�z�?T�6��w�Q �d�TK7���)Tp��g����%��ew���n�%��y����$d�THL���4+�N�t�L����sE�:�������߃�zl�S]T��^��*�G�jGk�V�x��2s:���{1+�;���h��M�:��9n�d�/8(۽]��Ob
��V�p�Ѓ���l+�Lge*z
��;R�![vٷ���<�7^���:����|��<��LX[�A���ClUVh�U��W�����G�6Յ�7�����	�`.2�C���v:��G��E�t/����k���]��^��x�	e��U|+�_9�d���)DU��,6���;�Ϩ�'�7/a�a���ܾ��^ρ�9����������<����xT�<7���
�W��P�*�,�WO���=C���^*{��j���U�B�w^7n_X�so�x��:��={��ڋ���T-��Q��z��'+���p	�>|��+��n��=�׾GI�����HX�S�@�>�y|l�8?\�V$����xo�XwbT�v:�p��=���D������	�:g�Ͳ�ib�և��?W����N�����;������ͦ�#辞��B��ޑ�=�Z®���Q����e~q9��./6|�W.!R������=W����>�=���6ŕ��"S:ٳ :������w�=�wc���C���}˕XS����~��a`���e���V���^�����UB-��Ӌ�SZ}%^��~ժ�'b��kڹZ:�C2��I�,~o��o�צ����NM{�ۃ��ޏ5o���|�����͆�S�BF��O�"��ϝ��\��ى��a-�$�O+kJ-ঞ`�n��W��S�ٖ�<�{�Ǣ�����RV�b�iV	�ހ����ՔS�'�yϹ`mX�>�1?>��: �6���=���(<�xe_�֓.�l6�w=sy�Ҷf�&=�w2�ɾ�_
 �����������{ֱy�|���3ۙig�:�gp��"��eIj�|�:�5�I���Iq�b+ʯ:�2K���b�g 5q�0k�7�d�z���}�k�����LJ6{��}//~�ş��w�Kgd(�ϭ�7Cl{����%�`�T�[��n�\�����җ�g�؋�¨�c@6#�vjn�K|���񼥮����Uᨮ+Y���*�Q��Y?uʺ�E�x6|��N��.����J�ӂ�.ޘݩ�C����s<]����H�5j�����~!�˷p��qB~�(:��ѝ����AH�H�F�������R�ďL�\���e�G���2�jy����D�F(]$�Ѕ�#>G<@�~��h1,/P�^Y�X}(��Rmg�B�Q\��E�t�1S��8�!9#��A�_x'^P�z��s�����'�6��}�+c�4���W"����c�+��]1��x%�a�{�[��9�R�e9b���۽�LWh�3��|���Ҝ�d�K�\O� ��j�V��[��fr�����m���,++��E��ǷG\N��L������t䨪����]��|2)���|K~��v�V
>x��ٳhG����ȝ�|����E?]y������'�[i�d;V�`E�z�~ޟ���]ІI�y>c6&��e�i��� ����(}��7�^��h����9���Ożτ���*�)��_Kb���`��rl�!�3���$�kG�oo��0h��A�7ȥ�n�}�g��A���L|e�}�zyVb�\�@�aaaC�*F���wXX=�,p��Æ�N�[���zx�C��=\se�k��5�e�뙓�K�cs}�2��L��
o�T�\]�<&�|�oE��g�uBR'��Ts��*�enٺ	�S���ɳ5��Ә�sb~�͉�{�T����[�d���6Xx9F���J����}%F�|f�ώ�]�����d�
���_U���X%�\��G��G�f�{��S9/|�=Ce���x�����~T��n�>�X-:,y�
���	��b���s�_B���N����U&s�<�>H���anT�Wu{��\���C���B �J�,��_�ˬjhǻx-�H�K�)b�jŵ=��}3����VpB�Q=�P�bn�m��/�Fѓ�s�Qv*�O :�=� �)M��Z=Q,*����ڳ�f���s��#���E�i��n!^��
DP&$�Ń�d��{k76%�x��x�Yt<P��7K���y������XL����z��EJ��Zz�����o~ɪْ�L����әg�z�^��m�>҂���vҏ?@���n)�����fWq�O[o��0�+���+��WO�8�ݦ� {5#}'t47��ސ&��o��z��DY6h^�����*%���nN��Ħ��r�d~~�=��v��5�\�ȱ���|�'�J=��S3o�*�Sf,p��Sw�{Uw�x+\gB<)E����C�䈡�Z��`��i�7�/�'G�����Fz�{z�|m����o&���#A�tخ������]�Ӳ��0�+�}g���x���x��grJޡa������8y������ٵ�Tǽȓc7¯�����).2�z �L�����2T����&h�}���3�߻�D[��X
�GΚ�(��r�V�݇�tvs=�V�݊�$�hI蹮�[佂������$�^�d��+��+o�%/i��-W��=���T�r��ݟ������ @>�<��]���Z��ˏoy˚�&s�qp&#=�m�3�l-γ�'�P�P;��Y燖4 ����:kM�2W������0�u��X� ����_���k��x/������*��93��K ro��*��5�Ǘ�`�� ���;9�㺚��|2�5P��DT}i�#��]���O��]P>���w�#�=����Yr^�Iޕ7��.�ex	�ï#��eI�FGfPY�ets�$���1Zz
�d{
z5��ۄ��i&��WJ��x�(�U��凜z�u3I��\�����:RD�Z;���ǫ���#��W�Wn�V�����U1k�+��Ni�����\ǹ�(�xC�`�SG{�g�V���ID �a�$\誩u�oX�S���\fs�D�dܛ\H!U ���n�^n�z����xq�s%HS���*��7lVN������X�`|>�ݿ\��c�C�]���_ku�_=�ȇc�m���{W+�\�����j���g�����<�⊬�%��n{½U�D��	m�o���7/%X�,-Q��2'i׷}�i�w8����b��#��lAa򖸢�
i�{3Gd<U[�5�oV!��&&�1Aj���aHUϰN�}=���ީ��R�q��9��XٵW�Q�'<�FI�'�H����;v���,_�q���Nʾ��w�3���ŞF�:lq� d�������8{ְ/9����o;s.ETa�H�J��G�����:�R?8;�]�y/a��Vw����d���l�e>��|􋗂mkgҎ����z�d}���,ر1C`�aorZ��׼��q��Y����[�V�� ,�=1�:��~������r���/Yyv�V��E{�O{�fv1뾣��o��笵Cjx7qz~�c�Ңm�~#_r�7�3Gjнp�[m�%rj��Oy�hn�a�r�s�H]�gqY���i<��i������R�%\�r�Ɇ.Fst�/F�>��1��Kɸ�B.iu1����;UƝz��g����g��vȉ{�EH��;L�뽻��w	J<Rʩ-*G(T[gt�Y�Z�c:+)p�*�R`����d5��͂#V�u�{7/4����ebp�A��j�d�/\=Xmw��u�}�Fp9���o}���,x�w��ЛGS8�]:�$kt+�;2�u�s2z�ۯ�l�|n=�A���f?n�8Jx����O,��}sӶ`�0�wB�/3xya���ȣ�.����C�t O���= ���������w�v�e�,IB��]���,0F��rm\�F�f��q�|�h�:Vhe*���:�YM<,3I�W/���x���"9UO�������}��<�HW�w6��"��?l��1�Q��7������rI��-�]�le�k��'sF}(>�;��l�8�3�r�xb/|������PQٳ�%�`��N���������S��~�lxw�/ ��������7]ѽ�J'ge��&�˃�^vf�{���μ�j��Z�*��xΡa�0�âO7����w.�e�r�A0�m�wWU�ת�ݧ�_r]v G���٬K����	޼st�zEy��i|�����;�cYgzi�<�����G�K�5�˶���h�uLg�
������=����ye|�Q��{ݫ�Mw7->ZLCT�ݑV\u�\���R��\]�z�vn��[��>Ξ�W��0�v���iG�&��F+Ŋ�r�ܝ/v�9���6T�q�H�2�;���;����z���)J��_a��f�LhSN�9�q��Λ�JT�ڵ�L=����� r���/��{|���~�es�c�����e =Ѯ��5�Vk�Ίm�T3t�4���jQYU�-t�|�j
6[�Ҕ�.v�8!^۾m�*�`�T;3B�����ʽ4���*�R�*{�1\�C�7�z����1�%e�<���K!Դ�l�"���!�g'pj�gQ�@iˑ�|wk8���L�r���Cm�<U��d�޹5kl��{�:-�
�ҧ�ݧ�'�p��c�[O$F<�g\�+F�9:�I������g�Z���nA�5癒�K]p��Ӛs�#���x��';������T׵�C������R�ۘT;7[��ݜ�[l��Ou�r�ڻ�+�l�e8\eIm7���N'��~�h�פ���o�����%Zi�%���I����&�y�b��g����)�ܖ��j
�֊u�ջzmkf����!TԑCD�ҋ���V�QM�,�Q<�,�j�E6<~?�����T�ƵDQiզ���Υ�d�&r*�B�$�S�Ӭ�hy����~?��U�^D*&�b���뇔��l ��H#H�+�_���x�����]D�H�NEx�TE�fZ�ĆJQ����Xgls�T���W�Y&�9�H#�FuŮ�Z<�=t��=5\��`����U�ICQW5U1(�L��u�\�T����J���Բ�+#��ڼ���R�A9�Q�\e~�"N��Z��7ozx�EE�U;#VN�|�0��W#��
�	+D�C�E2�ŭ�W���:dK���n^���$m�����J=�G�~����%�惐jw�7��u����6���~/D\}3ŗ��"��)�-��t����i ��<�%K#��E�ue�o1�n:(P�]���5k����Vʒ�L.�}��~�#��I�!U�7�E�z!{�QQ��wz�M��c�(�:���l���}?0U@+g�z	l��َ��;�;��>��̓G^����ϭ����s�;���El?m��6�;��L�����S";�
�w�y��O�ϗ�"�E]^�Ve�P3"<��1ww��j�O�8A,��c���;��9��T"�Gd;�Q�Q�ۯ�Ld�1��DtAw���G�����uj��>�df<���Y����Z<W���C~���!�k&413ᆀ���{�B���Ǫ��GMO���\Ҭ�`�k�/����}Y*Ǯ$h5L0��ת��q3������xzp�S�?�շ�&���k��oې�����z��E�����+�_��n׶ϊ�^�%��좻Z��!>�蛤~�������o����y�&�q�=�'ݢ��(�~W�_N̺����f'V�"��V+T煂�3[r��'^mk�]���C�r�eE�Xċ���q�2���9ˡD�T�p�N���}�`��iD`�\r��}D�\"��
9}�/��>Sez}(��U���y�:��On�ϙ^f�g�[i�q}<��ڍ�������m��{*Čء|!���M>���l}�����ZR;�uu��=U�������̞�;��r���+�C��u��V�½��w���V#j����W$^{��I;G�����騪3*7fe����7�Y���4;[vU��>��}�d��K��qz�j�<ԭ弓����B}�fOKۓ�����ۤ�,�k�T" s����ŦI�9��q���W_<�رR�R��ܫ�)3r:_��d�s��~B6H�ِ$/�x{�|G�Bj���}�ڱ�W2�����[>����&��^	�<u�������0�I�X+���-!�xm����UK|����K׿��q�O%�F��W��
����X3��D�5]��n*��}��Վ���NJ�18p��8��k���j�ߖ�2؇��,��Q��6RX^��b,�!��d\p�,|�!�:2��Sa�\:��m��T���#F�r�.Z�����9;c���+֘c�e8�۾��}��]k�?:��{r\�������{xs^�d�1ȥ>�+9
��'�:>�JN�c*�_���ӥq;ᶄ֛
�x�s���P��-�)%��5�����{m�۹b,uGh��z,,U��S��F��=���}~M����w�OL�?�&5��Jg�HDe|q{>�q h3�8̣�z�}묿���4������ur�9��e����.}W���g�N�_L�A����)T�����UFI����́u6}����夥��+/0.���ȟ�F��6�Cc7FF�1b=
�c<�r�+�+ZiD�SN��;���,��,9����ݏ3��|+���+��C`e���$�H��M-2�m�O�*�u�����s�}�ȏT�޿a�'�F��>+��u�:僶����[���*ד�7T��Fzo�QQ>�}t8>��ٶ�/m�>nO�g�'?O��|�o�[H'����_2慠�2c7�����V��\��-g���u�=���Fo����I�J<AKn���0��N�z�pz|< ��A�ޒ!��ץ�ފ�i�����S���o���ֽ=���µz�������ި��5g���$��{0q�ge���I�W����!~�8���0_�hy��{;��ԧ
�򦬥��}�]���%�o����z����O�7�K\%�U����X�����Z$�����]^��yvN=��n}�G8�tz8X�	�ߒ^^��Ĵ���X�߳�ʽ�»���g�HW�x+�2���w?�]W�K�4��~�$��X4{�����!��^����#w���ۆg��O2/F�3�{�D �������4~�A��O��l cbDEy��v�k�C���V�R��z�Hw��V}�7�rj���:A��>��ܶ�>gw���6��5�S��9o��6�_�w?���������(o�g6��c3wG��2wɇc;��Nw���}�1��ҽ����v]������C�|g�Gǘ{���kV����r�V��7峹��+[�]�CwnL=��x�\ҍ�^>�)�Rx6L�y�ɫ+�vKM�������	��.}�{��)���o�L�9	�V�.--�r�vN�w�\-{7b���#^y�\hb����ȱ@��̡�f�ï���E�Ŭ]�h�<���
�Ws(/
~��.��}�>�[2.u�'I�C����þT� Qd=����>݀j̊�܈[�3�]d�1�nD�A�H{�EPo��@��o~�����۞0o�'z���Sj���O�����+�5} ���p�!�C��5r5�񛲺:���օ�^f/��P��	�pjKL���{�޴�d�ڣoN��;�8v��}g}\ms)�ʒ�JD7�B�H��W�&߯f�D��{+0�v�I�X��}�`Al1Č��{����fG�=sq�}�r�9<K��f���-I�����C����]�]p�0V[��_*G�H��u�������/b.�TZ#(d���G��Q��Ԉ�(��X�Rq$`r�Z$�����G�RmW���_(W��I��&"�d��c�pGDP`��j��z�����{��}K5�;龨Q��ӛ��zEP]=*�����&e���NFe/+Nk�D97q(�k����T�7���~
�O
�eo���(�s�ü=��m�F��[͉�i�F5R���gF�jD��s�TU�M;���.=Γ��{�8]���6/��Wș>�o�X'�'�%�X'�����Ż~��g����Q����&�qk�-������]/A���'�;X2#p���̜�k�^^˷o�9�ɱc
���M�8��P�)�O����#��0��A��z�/6Ez��A�L7��Q��O�|ޓ�_�=�{Zf~�{=�~�O}XE|�N����O>Jۻ�
�����z*��!���ͣH/f�粯6$PR��)�}�"�>g۰�{��2/�6���^��bt��y������4�lgޢ��K����ۙ���*����V�0�Q֭.g K��ޚ6Xcfcg3WV��|N�.��ڲ���o�hv��>+z!��O���vL4d(^͟b��x����C���H�G�������2Hg�:�҉wT ��S�b�H�Iݞ�:S�{��,�����ͨ@g��g���}��m��WwR��Ko��]���k%]d�Ľ\�/"�pt&��W���R1����v��vm'�X&���~,nt�����&@ڡ2�	Fd�k;����G�Fl�����Բ�W_<6�`T���~��?~�������R?xF=�|�LSv�y}�=��jCj͟_ü���>���!�q���M��r�]w�^KG�8:�4UX?G|�6$���|h�/��������-q$d�j��J:�|T����VpB��D��ǃ�oَ'	g�]<��|s{�y���>S����d�q�VR�\1����He��M�w��Y���^���7՚��-��^% ��5�/�� �r�&��s2gm{���T��#����;�e�o������l,��Nئ7sor"+*tU��Dd����y'��@Ч���Y�.�����}���.�Krs;������t�)t#{�!yUc��a�^$P�����Նnwq��&��Ѽ=�8�ai����پ��M^D��:C|�Fk��F�dߵ��G���߇��P��#�h/���vS�%����$��G���V!ݢþ�u�a7�'{�E�<��|����~[Uy�\��Fs��ک�/��L�b'w0ȳ�+�Ŵ�q�7Ml	��7�Hajc��j�"Y3��5kӍؚ�������=���-�*i�	����v�g�*�<6���7�I�Om��4-x�۲��`���im�݄ʱ}NQ��=�P3�(�� �l�`�P����l�^��.sC6����C���"�J�T���O37����{��1�'���3�i{+��h/3UC£��s��9G�}5|*�������tR���E�j��嚄�g�5{��M�|_�SN�qlO��>�ϛ�v�h�	q��g�;q���D�Q^���]v�����~��>Ǡ[+�v�rT"A
:����˵�r�Uc-H񯄨���|���97�S��]g�V����|��6�>�>�tz�Q�}`��^���R����֚T�Pu���y׵+�6�;܄�kɷQ@�V�=Y��_{ڦ�HW�1���~C}>�^�f��H�_�YN�o�S�9)��]QM��:UX�%������K�YOU�"�ui�a�h3�R'��}*|���`At���N�5����"��m)��9wT�̬�_�z����o�fK<uPN�	!Ԍ�2�dh'����<��`>�;��!��W�%Li�
ז:�p��y��~J���L��''N|>�M��I�g�[�8z�^Е���v�=oՓ��f2�پKgo�me��l��L;�r3q��/A���
��,��H�{'�/3}�B�K�eNz|�{���J����P�@�Չ������ut?�q�v��X��B��7���#>*���/ ��{��>y!��~�qO]o
]�������%�v��M����xz��F��}��"�sp�����t!�-?�;k���̤Q�lQ
�l�I\�Y~��s/�݂t���X��'M�
:��_0Ĉ!����O�z�����m�uO��\|vk㧪��s�
&�\d��\������w�O��;YgoG!uG�^��~�Y�����Z�|@>���e�p��qd�eд�t�?���B�7ud�y�Q���iǡd��e�j�׼s=���1F3��>�pOwh�Hp	��<~�>�Y���+�{��ۿG�d淊%o�xDε�v�mQ{^��O�����3yc�����|��c�mqs��#$���������`�w�z&�����˱b�T{�jH��RY�(���3�)�	j����x��O�ϰ/oȻ8��,�N�.�g�1��y(��ŋ�9��30��{�����|c�4b$dfYc���z�������}�}eQ\-p�$1!��pn�����ώ���S*A��S�Qsc���9��BG��|1X��6=Q!���q�8�eu�VU�x�:��zqh}#w���Қ��ud���i�+O{��TP^�U]{�Mô
ds��̠$��oEm�lX�¿���5����	��5:l���Mk��~̢��{��>џ&��Q���	0���WF#�97��T�x�'7y!3�[�׷��0A��{(������'�O�P�~"`���z3ݚ���+Wkٷ�e�͉�(e�������z>�ׯ��]�ɋ���z�I&B���h�T�&�lt�4C�c���zY4Te�IOj}�y�'�n��5������)����D6�Z�_�ر����Kej��0�p���Z�>�*Ś���ĕ�t�%���L�����^�.T����v킺��건NJ<+�op��D�.ya�G��Z9��k�=�a߅��v}�OW�5:v:Ȝ���b5lŝ{�uW�v�R���{|wj��c]h�z� �ᙙR�o��^H_vn�ƪ
8�6��+�Jִ�O��Gr#A�
`�W���0^���`�Ц>q`��އ�x�Y.Aqm�C�ˈ'���|n�w`ܭ���rK��b��k�1�)��&$]*F�����n����}:���t��y)���`�F~pT�p�
H^�P�.�<�{N��(��'o��:���[�Ezn��4���x�+"��AP����P��s�_//b
�r��:�������"�Lt�.�=�c�u5\A�8Z���pFtd�N�F�E���Q�t氮�fR���	��W��m�{|�^]C:�ˬ�,����]8)���G5��w��/O/K�C����>t�o����'G��嶡+���cv����7+]j}�B�7|�;Q0��KCՕ�pǲ�)+0wL�:�v;Y�x��d�s�ә��r����2]7�U,���u%5F�����ҏov��[�����%]S7��s�nV:sV�*3�s�%9���$�}R�es[����و.<S-�
A�Ꝺ��g�P����L�[��<���G��ś��NR���Sm��wm��-["�p4�W6�Gl�}}�Ï���s�ۇ{�-�@��-{�q{�ՃJ�^>'��;fś���O:4kyzv�l;�����O�����u{p=�$�I�T�<���F����/c��c�v~��(�̪5s�W�$�7�`�M�E�1]^���س�=�vwI���gew�)��9x�{3�R�m�ˎ����}��n����/'��ɫ���v�)(s���&����;#���U�&d����jLe�t�妑���e�	�r+�>�����ΗN��b�a�FG��+�Iw��v�.�tW��x��|�>[�]���|��z�����W��M[�X���츟)��\�b����(f��K*��{B��kU�X�a2o8�Ʉ�,�z�Q�u�o��[ �j-�mt�f:n���;!P�*�kC�s9@pw��6N�sz�/��I&�q�6�ƻ%�wD����[�*pO����(��z��>kkm&��y��������Ϲ���Ҧ+�c
���rUz���ń�ݏ��%�G3:K��vP��zV7�g��/����{pE�]׷��2�N�:���/t�8�0����goP"]T�b=�m�zN38>ڭ):H��ӯ�ZDF��u�멝;�;f_l�KQ�Dgl.Kr�]d����Zc�K��$�DQU��kr��JS�䞧͉���)E%��e�U&*b��x������"�E�DF�TR[!+�dP���P�����Ǐ��������5*!������yB�\��u�d���Ǳ��^�\�]U������R�~�6�%ū=CQS(�q��Oa����꭯W����/��U|x�~?�~"g�{L�r߱�sW�����EG����{�l8i��r�9غ.����X�_m�� �I�1;ѲozS
5�&|���C��%�U�	�S�D���J����^Ǔ�{�:BI�U.)*��F	"��Fw]y��Ԣg�����>����F5�a3�V6x�,#Ҋ�
U9ّ5.e��l,5R�<4�
==sz�>H�\���4�W�Y�R�4Ʊ�V�bh�T��QV��5̾���c��Jj�[����o�������6��j�����=ϒ��NO�[ĉ�~��TV���dڸ��Q��Gq�_ͪ��L��~��b��=�6�Zi鷴v�u~��q�K�_��m<��w%�)���1�����TA�̜�/����h�m�eh��is8�#ޚ5�D&��њsw����[n�>������V2��}_?t��[�Q������f6�*0�{6)<;�<9�R>���v��[t�4��꫎�*R��ҔG�G>O�T{ꀍJ*믙���
��>E��;����Q� \��LIU�v��;뛁<��~�?!N?¿Bs�Z���)Ou_�G-�>G1z��:��vd����<�&+��}?�>h�m���T���q���?�r��$uI��8]eփ��_�*5��ѩ�9�P�_
+�w��t�+i=�����
#��+���W��P�>"��,�"<���+a��p�, \I]7�5�w*�B�Y)m
���[Bz,�
�7�U؉��Ůf�������}-�{���|�m���Õ�&SŐ�x��u\����n�q	�yQӟ��Dr��K��z���ooƫY�(�{4��lPt�K�b����⛏Y/xn���p��:5��LT�6f7��{�HN�~��3�1�wU�������L0Ec�k|c֫~f}t^�=�oc����DhX��C�3=����*}V�'�3���W�_g��
Z���5Ѝ�ʹW�tJ�&H;�L�����j6����q&��ir��(wܯf����(ݸGm�p@�������Zυ��z�kT�xN��V`��c���Zs1�EnGb�a��gou��������!����{��H�m��ʜ��hƝ��㢍Y�b.Mr����z��o�|��r�;m�ܭ��gܶ~�#v&�����a$L�y�)�>��A=�!�j׶�����+���;M���s���ewV��@�mq�l��U��"�}<��Rv�jh]��/sQQ�g�w{3�y��T��-ΰrz����w���;I�Y�(~��S���+un��t�0�����HpQ��
$���p��7�6f	77 �V�/�g��M
��
u�dVZ�&]8����vyzS1#��Z���{Z��q�"����	���Efz�´r�i��)�5��պ�"�b [R�������-���4=�ZE�d�V�]�,�s��i�.9��O�ِ��j��S�vǵ���Y���9W��u����&av��Z�þ}�_�}�H.����Po��=@v��+@�Zj"|*_S���l�e紎"2h���K��J
~᪦�,׾�׾H*�ޝ���V�j&hGtT���wԗ���=��)MJ�Ί��I���j�P#\�^n�%��Y��W��8����)�l/b�q{�z0{=1���7C��IB��˱�g��gb���̿Xݬ��߼�w��v/}���Jꅱ2��q�]�퉾�ylH����K�^����Q��%��kV���]�^�jwVoTl]g�Ё�Vx�D\�oᾉ �/xb�د���z�SE��:�3ٕ[��2��ĭ��d��s����'�]������X��@��Tp�G�(}H���mZ�ٱQ(�FMT�Swd�����:'撂ȶ"��6w_6���s7�K��M�-ny���}�F�XQ6�:�R��d#4�?�?g��z����T�K�CqmuS��U�3q�05b\�ڡ�qi�p�Uu�7������m�Y�Ƥ��t���8��>߇<�DQ�}KU��K�bC_J_>����u�O
����˱=3Q�id_��7�=Kz �~��	�v����&~�Z"V2�o�:�kF/"M��z}g��}^㋚k���6�QO��Luk�g�;���'$f9�5��z�|y�$���M��;���(�짏ʞ��}�D�Ǵ�հ��5�	�Us�vh��	l�	���ݎ�хR�����s�ެ�$F�Y�K��e�G>��;׼q�}Я,�t���=�����$�:�����_�c�����_ް��Q���G�얯<x�]u�.�p��Q���?t���j'�#%[箩~���^~�ù���|	HX*"d�Z�Ւ}1�%�������ѷ����]��ش����R-�S_f㾤6��:��o�1�����-m���$dC��!���o]�':�[�p��O3t:���7���-��r�Ф�d �(�9�=�o.�� r�2���(�h3#&A|N+��)fj�Mp9�ۄ�p�a̕��zm��h����m����iΊ��r����g�>��g>�V�&���Mtjos"m�y��(޹�¡�r�1��Ogv�[�x+��g�P~��$dOq�ȸ#�w�1���C�^x�X��v0C+�v�"(s�`N���D{��sr�&�8�ǝ�����ڻټ�_��?}A8C0}M:�������16\x_�\qK�E;d6�g��@�K�ߕ�W�c��(e��j���W�������I4�fYYi.d�y{)#vP2
�][ߖ��#�[��àC�'�	�8�^�8��o�xV4�C&P�z�1��}n����.����__���8�]�� ol�:�u�X�ۨ���&,de�^�{�"n�ƥ���#�� #BYV(���.�����yW��Ι��������Ql�=�=�`�P��Y��}s�q�$]�on4��:%u��7�+Pv�nɖ����S����,�:�2Ϗ��' b�gNt�Y�oz�#��eW�뼒u�C�b�9��B�rUZ᥸�:Z�P���o�&�¸���Vx�_���v���J�~�t�0�F�Q'Ns�P72g��V{'<���3�H��u��'����j��ö��B]t�S4��,������w�~]z�8����<T��b����X��Do���G�Z��������Ĝ86�+A ֭V�,G,�7��o��q��g؜L�fF�N��u<W�j�4���ַ�P�j`����W噐Ǖh�S��3�$FL�Y�rS�S�	�k�ng��~m��IsP������D������#6���vƅx��;�ޣ���2;��_�����:��݃J
��o]�9�R��(��{Z)��/7�wZ�|������� ��&PM�V^`�����У�ވήN.(ZB��"|�(S~��6"��,w���Z�i�~�VF�C-��J��ub��ȓ��7��2w�[}h;>���/�ވ6�����؇�̾.2Ͱ��*�.}6�9R+�5�$;Ah��_^��d:��.�Q�9���2(�>'/H���I%j�8p�$]e�aZ�͡d��;{=���gK����^J.;\U�[����/�!��W�P�V�������7��Y�E6Pe1Ġ�)�Q
4�͖����F��~�n3%��#�)��@�*k\�SX#}sQ���ε��1s���9�\g�#f�L?|�>�3�g�d/�:�>�UE(���~���W�X�&M��˰����@��By�t�λ$U��@�^��5��-���a(�}ʘ��-�7��<��t�f�(���:o�ˎPϷ�+e`<���}�N=�lZ�g ���T(�cс��G�3�aġ�_H�;}�����ɿ`�^���G=K��iW�[���מ�b�4!��j�׽����P�e%K�e��+m�U��1qEv�7�e_ƢXS�U4�`�׾kIA�<�ݛ7���g�]����lsJh/��rtư���}8�U��8>���x�^bKT���aw��y16�ZD�����ƶxX�č0�5Q_}Y���۽��V�)�n��5ں[F�Mv�4�k�����d�����pe�����uU����\�.�;�d�o��
��B	!\���(�v����ya�tή+K��u(��<~mb��껴c�=j���}��]nvq��H�حQy���m97�?��W_��ig�&�&��gc��w��Kޝ�v^J񍵥�����kg� �b;.]1�̑^��<�-�j���Wk�}�3��ϳ�a��e����m�^�ǎ�>f���5W�'�t�v,o������y:��>ݿ� м�q�<%�z����/:�݃�[�Ou��{<�5�Z�QO>���w��2��ϳ��{�<v��K�V^��3yy�*�����������:lB��G���S�O��-�n���p��Pk�m����b󕯫Î.i���6�k��޷f�kkw�&��3����MO@z���'�h]��M�w��]��c�ʱ�۱w����n�b�%�X��}!���|�v̜^�q4��B3���n��#3�1׫�&�o�c���4 aC�Ӟ�����q�Ǥz����l"�{
����c_�f�/��
�S̼`��3F3�rr�ވq����Y�DGfW��[$f^��˵�R�m�E�C�鷕E�����̚z�,igh��-��w���\��j�$zE�<�YS�4eb鮯���,b�FLdW�uwI;[��۞����\�M&
v�%��^���1RD�;�dT��3����3�c���N,�T.*O�ˆ+ ��$�Ĝ�h��=d��f���v�:��<��q���9��i3_WՒlz��X��uX6r�|������5�����Bo���7�[Jsm�z�1g���Vz���g?7�í�=�~����h/F�U\�����_�����4W�9٪�3��ϐ�V�_o��m;yZ>�t���~o>�W��v��ٸ�ӊ�]��%}���G}{y+ ��w~�G>o��{��yӳ��\�&��xk`�o>M[��}w�/o�s�w�(u������;3:f�o�uuX7�'�������͞�%�<��'���@�e���Iڅ(��^�9}ǌ���'�p7��`)�M��Q�V�Z�y��?�"�N���4_ۈb�,g~�-W��W��+P��QD�Qs3f�3K��V��P��@ﰌ��BN�ӳ�c��>��@��_h���z&�Z�-4Aw
��퍑�&��*�:0�<D���	�/FN�w����/���J�H23��v/�=�M3Z�g���A�`�w�A��+:�[w�����yW�*+�{n���G��uT��6�B�ê��s�{g󳯫��E�gn�_e�Ģ	ɉ�����l3�0;cX�|��eOS�L���l�.��"Z���߯\^�ˍ���VZtX����������BBjlA:�ˊ�ښ��Ǐ����s��I��Wu�I��#����ٓOh�����ܪ�Z����.�|�ך*:��WaT�{�Y��G`>ίU��5�-�Ί������M��Z�XS»��X
R�dzU�e����ۨ�y��'$��%Q<xl��i���k{�o�w�
U{>��	�a���ˑlm�A?i3��9��sC��k>�������)��G��h�I-��_2���_}я/Z�p���[*�X�l`J����������S�y��քЪ�+��
������=������f���4J�J$JH+
�@J�*�"�@J�
�AbG@B ��o����V  ��
��$ @
UX V�@  �:�t D� � D Q( ED�D�A�f��Ċ1 �AD��EQ �D�" �D� ��Q kHj � � � �P(�$ `�@UV&@P ��  ,� 30h��H  �  @J��@ @J$t�� i! @BT�W�1��� T�E"Af/�?�����?#�z���?��[����g��G���=���>O�x?@kO���0�<���UE��?9�?����*���<*�" �������A��������}?�UE�g'�o�G������:~�o����������������+(
�@ 2��P���� J��"�����   I*�	
�#  @H��� �   @�����,���` @BVR  ��U��U��U�� !�U�@ �Ud� (@� )UL��Š�?o���
��� �#y�����w������8�#��>����
��N�5������?������g��ETQ_�����p|zw�� TW�QE����A�����M�����a� TW��O�������޶��:�|�D���ppUE�G��/���B�(�Iɽ�>O��g����F޻{x�`����QE}��~�UW�~�m�'�>�����~���GϢz�l}^TQ^����0J����������=�~G�QE~�����Ǉ�z�UE���_���zt>���(+$�k+�a ~�0
 ��d��H�>v�!$�� {�(�(�()I"KY*ѩ%*Z�i�P�*m�@�AR�"���"Im�P�(�U+S�ʜf�U�[U�5�l��KJ5���Y���mi����m�͚ʫ`[UKm��Ȗ�f�E5U�j�u�ʂ�ƴd-2�URHwr��km�ؖ����(�V٪Vʛ66��m�5��5��ck)�эBQCL�-e�f�h�-f�1�Ulԍ�ѣl͑f�LX���kA�������ۓ��U���  �t�ye��]�Og�Y�[�n�w5;��lk�M�����v�W�.�nܸݦ�uQ�maUWT�V��m�f��Ҫv��ތ��\˚�8�km�C���y�e�Y���[Uj1���  ��(|�mH����}�w�c##lH��[�/C��N���waB���}���P�Zi�M����z=uBك.�����N�vV�ݳ[L��z{Ƕ]��Z�l��v��Ω��M�;���w��khT�V���*���ڭo�  ��:#mֶ:�S�i��Z��>�{�wvm�����:��j]�Zڻ�ڪ��Fj�Jl��UM
Gnݮ-�ۮ�b�h��Uv��f�Z����^P������-����  ����[av�Jm��R�Z�V�u���՚Y��+L�O����,��6�ڋ�[k���ZE.�j�����{�<��,68�I�{Oy�v�ݶ����ha�d��V�����  W��f��:�iƵt�������Uۓ��$ٶ��v�u���Y�ڮn����n���j�v�����w�/S�[�t�X���du�uI=�%��l4���Rkg�  ���\Z�wu+skk�v����u�mϱ�5��u�����k��d��f�um�%.��gr-NWru��qǭ���:;[�f�N��ŭ�����Um �  w_Um���]����E�E֝�-�ҭUekoX�z�:��\+4�^�{�;��i�\w� :N  ���Pt���I%i�ef��i��%i�  ��M��Cl 5�� ��  y��  'v��C�L����Og+� ��S� ŀ@6�J�T����6+&���  g�h�n�� �L�@-���� ��8 n��( 
�v��(5��m� `�
�{��P
���՚���6��J�U���  �� 3 � ��  �`  .F  d����  T� �@(.J�  ��)��*U#@24Ѧ�S�0��� ��~J��i�R0 �E?5)*�� hh��&eR�� � �)P�U)� �~���#���ܿ?������ߛ��>���؍C�ő�1}*�Yϴ��� ���}��=�����06����1��6?��1��p`�����6���{?~�����b��im�V���/s�Yh	U�ok���q�A��)�;i�r��Mx@�|�ø U+Xʶf k.6���j�5�(�;@ly��'z�KEiiQ7%Մ$Nk����q�C,+HHX�����\�5�Ÿ�U�3��5���B�v����D\t'�<���=+�#�,Y��n%�L����M�+k�{e(����r���9�(�������KAZ��sX$�M���:�B�!a8'�h���K;���`9�q�A��	�f�dI.�O��󧛝����,�kz喣�֩�l�0�F�>�ǃ�v-Va3oNJ*�PUٖQ�@[!iۨr�4�59sE� ����U��aN�IK�uɽOb����;�v���Pȳ�R%p����wY��@�-qP��ud��d[�SCc�6���qX#X��`޶C�@K����{W��\�P�?��in��ڠn�c�)�b��Ws(���)��9�ic��,�ج̬r����I^+�q�7F����|��;�-i���̡W�$&���Xe3wr��-�0	xRW��9�� ��<��W����.Xx1�V��)�6�)h�r����X�iF�5���,ˎ����Tr�1Q�A9���3�v�QB�ɂ�Ʒps�8eK�������ئE�SIYBX8��՗7F�^��XU�pP�QR@����vͻ7+Q�o�i�).�w'�9N�$D7r%F��;=�U�-V��P�Oodwj�;r��oፇ����QL�0����
���4��*�6�G륊��,n�-��6*{��9R��Mp�1)�k��d�", ��+j]��\ϧ��ņӚ�^��B�,�9Aj(�C����%d��Xw�P݊�Y����v�_A�v��?��L�f�a3&g��,<�.U�.]�Ҷc�ڡ�chL,����Ӳ��%]�3N�Dr��ڗ���Y��hu�����2�ߖSē:#xP�YfLl����j�HrwD�[&�����rSG63��OWq��t,s�'QY:M�<	��7ao,R��CME�J�Ese7g2��n��J˄��'��+Z��b����!��n��p�%jŒ�EK��2n���0A5,xvP�q�wj�M/��N�&�-٢E�>�9���^uM�.O�u�m��7&�E���\�n�In�������9V$0ꚱ���j�U��/3㛖%G��7-�OMkM���^Ř���ֹ��T����E݅G	ˣ�ST	9q$��U�b��{�6ģ�����r�1�i�\%l7vѼ�kɧ\_X�q�O~b[N\,�Z�$k=�v̈́bz���t.���trպ����Z��B�����F�4#�9����a����|�^\�T���F1�e�`Y6lq-�B�V�w��%giT��Y�m�CvY�uL	EV,fِ�ci�we5�2Ze܂��x����BX�OkL�"zA�/]�!K�km��D�����#�dTM+���薂z�,������Q��边Z��1%�t0	�R+˧��� ӭ��o:��.�,9D���ek�d^�E�A�o6��$�D�h�s�ˌ]�t��;�e��ޭ�-U#��k�>���@��x�G^�pS�Q<�vP�"� a��W�2�Yi�ժ����A%�[d�@
pt�m'Ha��z�qL��4�8�r
ۼ-���/cVt�h��^n!��6\�n��9t�&���z�*8DV^��)�&i��ʟ��D(�7�-K�mTX6�Ӻ��e����Y���c���t�q!�����li��cӮ��L
���.�B�۩���4Y��r�eJݸ�CMF��I��I���N^�ɹ0��e*��Niำ3����S�^����Y)��"r�F���+����l8�H��s~n�T�͔D�0�˩m��us�F,A�Q����Ն��rD^12��JiO5�{QoxKa�̎��&FQ��zASq������!̩�F�HUY:�nӬ���!,5��Y���O)79�e4ٽr8D�*�Fcc�dL�C�nr',r�:ŰS��V-u�흹�밺�.�f�IC0��YRf����;�=r�I$��7f]�t�ջg-
���/9��5���\ƚc�lYX��*+luZ$s��ї��S�ʧ#�e�ժ
�)�j@y�@�OV���`LW��+Y[pٹ2����*�3kY��S��f�dz�N$�}�Md��۫)�p,Ϊ�!l��
Pq���L=�}�^n���31�@}u7v�r��W#�O��)��	Xa����H�����B�AX֗T�t̳9��둒qAE��cCJ�p����ЩJM�{[4�jJ���(1N����Y��=�����su���d
T*va,6�3��2��-y5>��4�ü�]��º��`�S�g��̫3T'Npo��1X[$H�G����\�V$[4a@��,��6ڽ9l���f���g쫜��ܗ�Y�QT���l�K�D�`e���"�@���vV��N�i\P�;�ӣeģ�n�(b�ے��!�C'F2s0��TZ�GV�'8���.9�lE��.6%6��}�jV��J�0��B������O�4B���QHw��[�ǐ�e\-Vn�e%݅�4�K]�s��eأ�W&��C�D2:����>��̩�;waF�\۹y�EC�X�fȣ�=��z2�mǰ��W��h˳X)�/�FiWxQ��Q�ԋ86r��Z4.���8K҆r��m�� ���$�K�+/�OW�lK�kѲ��VnY�
,1ڡ�f�YZ%�9P����qL����Hݗ���V���a0(׏�_Y��Pf�2�@Z�8���T[H\�H��%�]�9VK�k7�oB�r ��Љݲ]v�S/1�s@Ϳ��̡FE&l�����k�ie�s]���kVL��ݦ2����ֺ��]��AV�d�K�_:{�՞�ĝwp/qWqA�i��p���O3v8��p�P���G7q���D��ҁ�j6,@����=a1s%7cC�c/z
lrV�P�Anө�0��l��S�ԳEcA��U��XU�Ŵ�B�V����b]�@�X �o7Nc-,3r���/2���Ƙ7���|-uX�\�a��e���2�k��eǳ0l.��4BދwPIfKa�-��'(�<��gp��B�|Yk�a������0XJ��L�F ��x�]d�ѵ�lV���X��d،���S�99;�Sjq�$8ҽ�S�{1��s���*e�Md���_�H�̤��z��*ϟ��C�U��w �ʽVպ��EL�U{�;;,�AsS@�e��	���u[ѵt�n��⛀R�&̀�Y�>���XoY؆��!y1A��WRՒYY������H9�����&tz���a��a�aQf���+a��Z��ܸ3Sx�I��ӳ(�m!�,�����c�퉹/�	j�\�B����~m�˱��ˊ�t�9�c"VrM�A��F�=�ʆK-ճ������*m�ܣ#�6���:��kwL��xf�e쳊��2Tr���7+<����qۓm�͏���SG{7.���kQ�[�1�Wo�/vL�3q��է5�2�x4����%&��e+IϜ=����mݷ	�)������g:1��,��8[n��i^bhr�Z����=������x�Ń�nM4A�i/-��B'��h��Q�5��!�M:g2�^����z�Q/]f���g.�A'P:���o��xKn�^�����YYw黏�O*L��0d���JM|�vl�6�+c��!<�N؃�oJT5 �5��f	37AȆ��6"�yL�X�ȱGk2�̽'(M�m���*�ٰ]��r��Rbkj bu������6s	Ҁ�q��LT�9F�/od��"Y���n5�0��X\��C:�nљV�*M�밑�X��s�����ꗖ�e2]{~�XZH�1������j�ˀ�:���-"�C� �)�3�6�TU
L�o=2��H������^Ganr�%.��6{y�c&eUNP��&Ë�Ŭ��Ch<��%N�'���+� �v����CQ^��Y�'�MۓZ�ɻ���,��t��3�f��9�s�͵t�ܦH@�QV��G`i��`�,,&�Xpl�QA�Ҡm�p� �U2�K�#��K
@���2B�[�-��b`z����m�=��#���sq�3FHFk.�s]�ƙ ��б�����yf�1����Vk>��#͊�P�-d�DE� �1�:;B�-��%M�HH7��,�����4�t���뒙ƒ��Ű�ib�HY���}��L·k�D��YL^E3\�d+�����A�N��is���DB^�i�79�S�
ٛY��.*�{DYǺbV�I�z0�3J;��Jn�\pV��on����Y�f��6�ݣ��Vx54d��]�+:@W����c�9O#$��t�Nf6EY���6�bU��{�s�m����)q�b����3&�˴��LX6��d̼�(�F
�h-�r��u������c�����9;��<�8�֡;f�\���6o/4�.K[��NJ�����N��&6�z�.I1�E��]��Ncqc��wH����HE������M)88��5�AI�z��If�m�KT�,�;3�/F���YK4G\WGzъnm�v�5[�
J�!3�nXNi����/A��H�ɚ�)�<�-�UZu�e�h�j���շg8�gI�(��44��OJғnF�+!�R����0𽨜{
�R��F��1�[8�kS����Y���ÃV֩)�VCI�	���,g�ڒ�,Lɏo8v����ά�DI�Ks�T˸[�n�Ђ�n�I�,�����5ֻܔ�M
;�{m$�m��KT
^��co�ck�m��1�{7��n��kY5|KW!�wz�T)��q3�-P��e	%�bS@��������7y���h�ߜB2M��ͽ-�N�0�Jg��d���S�svYy��*�\�teeGP�kC̆�h�Wl��c�0ۢ���CQx�`�;Х��{o=͸[�cԋ0��ϥ
���L.��Ż��U{�h:��x�̇�Pd���� N�����B3id^C���_b�.�l$��!�we�v�x��?=,�R��ͺ�CL"���r�'sy�:��Uɕ&`�چЄZ�c�B�&F�[���.鵦�Mu��v0���]�3M]�1��[w@�rf`�ۼ���F��Qf*G�ї4��x�ǂ�6�F�H0�%,��-��\9?�Ŕf$M�����h����g6̻q֛�`�B��gi��4C;nۺ���^��P���]�%��32�)B�� ���Xsؙ��9#7,��>�"�-�R`�ƽZ"����Y��a����iܞ��۱�Sܸ/%d�ǫ����v����1��g`2�
��n�)��v�;�r��4��Q+�!����<��֑c�ݤ.;z��"j��ۄ�M��\��`�WR��e�5�5q�fb��NS9dh&�ǘx��	��Ţ5Nj
Ή�]/A=�d�اW�i�{ Ա�xʒ='���������a��wXPH�(�c�	���Vn n�Х�:�q�ڗs�`��6��B�*�)��Av�z���ޭF3iհ@��V�㫈�ђ��\t�4�Bs�,��ͽ��	gD�Xz�YZD�<ګ�
\��I�{x� {�XښK�Hi���ռX��Gimb"PfdqB��V4<Ii���Ֆ��� �)��\R�E�3A�j:w�J<I�b�T����6�ҙE�@�ȵ`�g L*j�/JKD����-���`��r#�Ȳg*;�n+a��ef�ء&椔{d{_��ռ+�X#\��K���j9׫�t=6-rl��5�"9��;����L�x��]x�We�T:{s�a�=zo&H����#я3�e%�&��zB(�Ƴ3[˺������@�+�l�%_����	��c{x�jũMѮ�>�7.2���2��F�
�˼6 ���k��VǙ�%Jv�͛B�0v@��n�+�]�D��OL�gŮ�ݓ8 ���j�o5{0j�3�(Zѓrʆ5�k��@L���������s+vnP�v�L"��a.�\f���+%�һzU���opڂ�$&d0n�RH#�2�ɹ�v��o`���p|�-�x{6��-tP/�yu����pZh13�C�5��dZ�ؗ�Z��XZ�^QFQn1lÁ\�t�1�Z`,7X�;8Ő��PF��k+����҆�	�	���˧\��lTn��:�m��0�},��x6���Y����5�;r�4Y��Lq��[;[�*���3r��n8�b�Z��ղD��T������/���)è�C�Yٝ0�P���,��ez�T�#aa�,���H�Q�)|1w5�P]���lX���!�Сf���ݧ�m��Xo.���N�:Ġ!KVʶ���e�6��l�u+�5z��z��up^|�y�"�V]�gp�t��|e����kSƸ�ܻ�R�6`��3�h[ي��a����'b�(��-���zkd��8�ԶA�l�-͡�P�j�J{dC��p��&�YyqU�[����G
֢M;q9*�2��\����ARfo�u���E�\�HGuB�\���M���g`i|M`��7eKW��]�$ټ��<	��4�ʙ]��.wٴb�s��{	�j�HGB���~��ʋQ�)+GI�kG7�8
V���|�coO��_�܈�Y��U�)���e�Յ�.���}�u�E�s,��N�����_E6��RΏ�ݶr9Y[�Vul��\Ucѯ:sǙ@�w{� �ˤ�\�:�5^��O*wYJp�Yh��l�/�Pj�08�η��3bzFݴ����)ty%͇tҽu��2CbrJk��X%�r�x]Ĩ^Z����W�,mk���ݜ�w-$��}F��
w�o���Z��/S�c�1.�KG����f�Dͼ�V�����0�m�b�eѭ؛|w}|��û�zR�V[ע|w�%�\O�ԑuY��뭐��z:w�0p(��XtK�W^��QZ͛�59k�a�P�S��3�7����=YMB�,��=�[/ǋ��}��c�lQ��������gJ�(
�7���˭�%%t��~�wȼ�O󺢻����Ưᚂy���՜�Bk1�G.�A-��g^�6��yY�I���˭�?���{�(=K���m*9�k~{w�����b�Oy;�����
e���=�<!{$����olsv������]���Lv���47D�c�K��|m��-rs��S��tx��MX�GA�ZM&�Zޮ����U�5m���:�Sy\(�ټݳ�l��X��yO^c}H��x����q�.L�{j�}��YZ�/?u�D�U�b�qK�zxb��2M���y�s+��QUw|twZG�<�|q`��ߜ'}8+JU���Y:��R�Y��0]�-����q|:ݩ��̞�,l{b�7m����j8w��9ݦ'8��5SHp��c��Ԛn��	Μ��|�g=k{�h��-4wi9e�Ve#1���4hE1cF��E���BBwV�S�Vݜ�d=�:���\�'۷0Eq=Y�MP�>��@�gR�Xo�+����˨d%]��ۅ&8+���{=>�A촯�SFu���v��ݗ�|1������-~��7��]�i�X�Un�pݽ�wc�nu�sRn��O\�5p��Ɠ͑����Lbv�	��R����nE�D�f*�|N��ٲU�ra ֥��(�7xm�9@pn�[��	���1ۦJ�Tj�|�\��GY����^ც����SqH2J�p^��T+oA�m4_\�_r��=R�z�.{���A�:li;GlJ!������M<-�l\�1\���m�X��2(�Hv���8�\]�,�B�4L�K�o�^̈f2�T��X�Ԫ��&�^�1�+�B&����17�����D���C�ef�%M�+���*y�pp=y{9'h���׺�]�7�[&�bN��ɸveťc��!rwd�Y���ӶAq�Z���-��	!���0%�3���@3��E+�:�G�k����7�"{+:F.!wxAQ�w蛢�|�hÎ�,X%:f�.�y�Q��	����2�/�8\5d�|�hX\��J�P��F�t:)��&��ϻ�T��b��ߗ:F;�n�選|u��N�l/�|��,J�q/�t�}���wL`��t�{��o������[�5��ѝ
�zK����z�>j����svu9;�%�Q��9A�N������z�bw���NB�y+�mݷr���B�X�5�8T�o�E7���Dd�����,�����h�Wfw٫/kM�J�E��Bh4��A��B��E��%�S۔F�(��/r]�1hҕq�[#�[��f�$���9��^�:/j#8��&��M��Fn�x�Ϛ��y�g@%�k��2Q�3��L{�e�#!�g,��6����;�����g�O]�[���F�1�r��f1����<s6'�<�9e)���Љ�X��8���TLe��ŉ��(����S{���iw5��{8�M��{�g�8��G��rSL����.���au�:qͻp�2��޷|"��޽�e�A�(<hG���2u�2�C�	[f�J�N��^�h{�9{��T,z&e;�s��鹌&�����3yGu~�>����o�f�in�/S2��Y�����栓=��3���c�	�hJf/W��PQ��Gi\�p����l�ґ�I��y	�[0Q�#�1�Ԅ����%�[Mp�����H0�g\ީ�O��P�s"X�bq�%W�e�91��r�μdE�����x�Ϡ6�H������4ӝ�o1�Ԍ��ۮ�"�Щ�_��3v�WM�U���y.�Sj���[|1��+�m\�̵4�:c����E)?�d>�5,'�'Y��;�����.O>�E��5�t�2�V���G��<B��N�����Bu<����"����q�'4��J�;���k��� ��_!
���h�%��ֆq�&��o^�,�u��h�#M���e�^����@̼��D*b{5o����f��7��,
g��AJ���"���S��89��{]�(�F�>�Z�p���l��A<�xg_n���$7��XKv�:EN̠�Ħnc]2lW���nh'}��a��1�����o�Z�[#���B��b&��u]7�Y�e-N��b�;���/$�mջ��Xʽo(�r��,��̷[��"X�Sv�j�S%ZT�<�N����/������0�]����ae>�nw*W��ʗ�<׹���'�q���	�l36�sa�j;�y�����T�0j9�C٢Q���	�n���}+�G�ON��OX\+��f�0��e��&�u�g�lfdy����s��s�}�mV�����v|͚�ѕ��HR%�n�yѡ'-Zֽ�o��"կ�R=�����z��J�֘��⠑��[������)��R8�����R���s�Ў��9�9�m��b#^���~��W��d�Z���ny�H�|����tȨZ�Fm�s
~�3�5�F{�M|��4h���j�����[����)�&uw��F>�r�Ӯ��=pp�Q*3m�sJYM\��*��Ѩ�4���J�4�1CQ�9�]\�2��v�N�щ䧼vC����ї3B�I�*�GQ[��A��v�q<<�ќG�/ϴ^�|�`1'�a��lcf*�o��F���[��ծ��0�y����K�Vg�pQ�Lk��fv,�C5L+��,�f����l%5��G����w��sfA>�g��W��5��xyZ3�\��Ok��7��}+4O,ѽ���l�кyle>�/w[��
��5���L�tW9�Ʈ�J�֐���FZ���-9Vt�--���p�)�d�zq���=��p6d�ѽ9'�t�;��G{K�
����9ٹ�XԎ�A�[��r_:����F���%�O���sĂ٧2N]��F���ݣư8���~�S�l{�ݤ��u���a)�nizEкĉ�s1��n�-rz)����pc�i��uʁG�e�M�f�cmU�� 7mzI��3���-F^�����>�ز�5�$+1ŭf���@(��F�-��lI77e�3�o�s��0;��S�A�r�\~ks:�917�ތ�y�tN^6L����Q<%� {��e:���{�l���=��+z:5Iױ�`��08�}�+���b�̽6a�˨. 3{S�,M�V\�\&��8��U/���ʷBZ�|��%��R4�4�_;�1�7�+'u�8�����oBxI9Z!������xh�:�4sm���]K���2`����A��κ؈<��|�"�����+	��q,�|	��s���xW���6dv�����tj�������n<�/��c��Q����^Y��Id��(֨8��5��C[��Ϋ���]ӣ/���`~%���Z�{{Jpi�P�E���$}y�W��{x1m�d.a�1+�����QL,t�t��Gh��D뒁�v!ϲ�zϻ��<�66�6�����9�LB�m�Y�Y�O���Y͜niF�6�x����z)+Cx�w_|��S)��+��"�3㽊�Z ž�姙-��t��۸k�E��<�~K��`s�ݞ�9:�+�٥� �X�%Z(n?�\�{�z��&����j�[-���u{*�hY�*�x�?5���»��Vz���J@�ݺ=�1K��_Ķ��#��� �9և�%_Ma�/��n�Ր��5��ڃ���G��X[������'$V�jz����+/[;��Wv��63�E��e�[��O��F���u��e��F�U�E�����M�!��m\�������Y��$�n*1�2�Tzl��R�P�^Es9�k�{Le��7����Lz������-�s�N��RGMdx�H�wU�Ι�uټ:d(:UifK��TtX!X}����{8�Wd�!�����GT�Pϧ<_�nڝ.�\���Qs�5�پX͸�罙oSeD�ZD��\��[B�gd�w:���u�����JXA�V��K�r��̊�H��[��g��=Y�Gf$h�2m�`k�r�}�'&*��1
V�%_�74������ջ���/mvk��ZE$�^$�n���L�/7u\�-M-q�/��7
�M��9�HWa�+_E���/��r�Hm�ETر0X�Kf�=W3].��T��h<u"���HE1�70F�Q�5�ɗ��a��]*�/ ~��aJ=)�p����MѺv<�4�6�J1rcb���r��eӴ��������u��	��
G^��i��Q�|(mK�ѹלD����=$�b��PlL��,-����?^������}���R;.H�Q㳺�;m�'�k*<lvu��E\�>Ӛ,s�1��XoTC1x7��94����v-`G�37bt0��u�;6�^��j�Q�%�e
7��FnW����0��i�j�A�龳�:��i�	.�x+�5��, �O_/vt�x�9L1]^��vjTh�"3�t�{SD}�3 �;��g���ƣ�!�	{ci֋�l3�_m�(�|Pi�vl�z�R����]�A&aB5vy��"e\��!u��q�R��=�kl���i���aW�k���F��9al��(Up;�EF�c�;��j�ݑ�ܼ�v��n�m�M�ov�Ϛ�-!n�R+���w��s[?	�G6�q�;_nL@@ 1⅋�z/�#��9�ݞ���4#���r�1��IWA'�!P�uu�Ѯç]�����z��>5xF�ٹ���\�I�f��%A��Y��=����u��Ժp�a�!R�5�-F�$�k;.��l�v.
{��_]F׻g1u��ýi�����*�.I���f`s*�}s�m���;5������i�L+�7�5�<����+-f�2��e�R���Yy�8Q�l�mZ�sY��n�f�)R����I��Y;�T���Pz�����s�z�N�(�Z���:��w�-|�╵�z��.�N�k]��ܮ��d�{����Vl6fkйCSF踝+���L�u�֫���!��s̍��\��-z�uEA��I�S+طo�ً���C�����X*)r��z�.O�D��,�^Kh���.Z.����q�I���^���L��9I��ݫ�m�&aʹ.��|�4�]EY� �)�T�c�`��{0Ꚕ��z2y޴2�o��!��{��ӓ���H��v�W��##}o�u�f+������.�9�Bèix��ޯa�z4C��I�s
/���4bqq�)^����m��]}�-;bX8�6�vχ|��!I����EN�աЭ��V-�P㺰��kR��$�+j��/;N��:G&,�Z��X�D��ؐ%.p��Γ�R�ns>x�>���m�U���DO ɴ���|2�b.���Qj��yeP˚�Fv����h	�;n=��lx5��&j��b�4D�ڂ�!�`�ܻ;�C��w�蟐[O�ʫ�]���O�� ��<�f�v�v��Cp`�v�ERnk�d�!>��kb9u�X �<b�0-�y�n���S����n�lɖ�k������b����t�@�ژ�J�i6*���]5Oc�)B�u��Wlw*��n�w�9G��*"�w.U�;6��ގ�����u��]�'X����`g>2��M;�}4oqC9;1�GE?���}�0L�le0|�n�X�fou+�:����a�ZΡE��%���6�
��j�o4�#jnb<��Y�ʰ�̊ ��v�^��݇�o4��0C��.�U3s)��z�����[���N�G$�6hX5�=����w�'h=��O�^��^���R��ј�U���B�Y��
T�z���5Rv
%Œ�bۦ��:�a���Ak��搝@�ԣ?>vo��5��o ��ұ��V	����CC��φJ(!�rþ��0>c��-�w2��q��C���Y�2��];u@��|	�bn��ӧ�������Ţ{Om%O;�sc�M t�ՙ����i�޽�0���j�9�,0����o\W{/8��6GŚ�qZ�8r�x+'Jͽ*3�=���^�+6�:�z�=����c}L�˔5����r��/���{����a��v���R�֮/��W�Į�>X�y��I_u�`J"�1�/+:���bouͬ��J��1�ׁҔ���M\I��������3�����j��P��N�'Z��Y��p��o���me֊1X��Ӧ�k!�d�SU�Z0�K��e���,@�m�]�4�d�lss��d��Bx@����˕v�WN���h�x2��Se59������K���:��v
�܊�*����+�F*H�a�y�!�,����S3�|��Rj���s�Ҟ�γ}�:�7��<�q�<��u�=�R��&���J�y��V)�)ݴ�Z�`��z��ϯ����cm���l�z������?s�F�0W`騌���W���v�!���k�����6�0
|�ל�� ̷ȱG]NU7�u��V�Љ��f�٩c�V�P�a�-�WgXJ7`�J+Feep��)ݯ��]�`���t�(J�`^��Т�y�(�R"8��#@8e���7�P�޲7�㨱�ZX�������Sm輊�^�+�T��4��]�^��dQ��ܜ�A�����61�����ø=ۆ4�pZ��G�6KԖ�š�W����������(V�V��o���u�zF��P�c8�=jn��ݒ�������<�[��*TP{�ʹ83��ͣ�	�Zԭ����<mIY���Iv��k<\�έ��7Ox���ٳG���e+�UẔ͗�Fu�jN�2�w����������1�pr	�g�=�{���E�R�ج��;.�M3VHQvY��QO�mdQ�y����TԖk�]%��Xvr��r�3��n�L�{��5���{U����s�L��P8��Ѵ�dٝ����X�"�d�<�hG&X��Ǳ��&wu��/���on3}���j+yv�]p�n�vR�[��i>,�)[�a��j��^��6�9:�o�-Dz���:nqT��Xڴ�b/s*/�(c�r�U���/6C7�Z�p��h��5J}NOz����2����OC���qix�ǳ��W!|fe�[`����8,W���|�
��y}R�U��_fxI�r�^�#5�E��G�p�]ᄄ���hE4`�Ì����Z�ӭs�Ә@�J-^n!9�r��,��F7�:Z�Uq�ε�m��|�2�_V;�Q�4|����\R��Θ�xd���V�4�K��&��J���C�w�L��ҞmB4����;���U�h��Ei3_'E��թ< �]N�
�6���Q�9s����g[��z�RPK~[ut^29=$t�B�̱jc���ۢ՞����˵���y�w=��u�[|r�u�6m_�� ��U��e�u�q��q�a�f35ɍ�ط��ee���}�_�)�w�.��/��+W�?h�}��Fo8�j�-!m[�ӽ�ٮ�G+c3����C`���(*f0��dR}F�-<��qt�#ն�>���A����K�E���K������XF�e0b�B6vi3zZ�h��u?<^�{m}�E��vvp�}�|\��ZP!�����:�����c@آ��������6�s:�.�Ȫ�f��L�(b�U40ki�x�������=��nɹ�a�b�����1c�}٢���q�yTu�J��p1�N�0�^���9��0�ZZ�+F�aZ�=β�lY��f�f��٧,
���e�\pI��\��o�e���1�Q������_)c�%J��$���V�+�l�Z�L{�����P	;�Om^���/K�M�Ƥ�g˴�<�t3�SF��K�nd��oM=�H%C��
�Yۃ�@�^%e��Ͳ��mF�h^���!�^zs��ŕJ�Z�y�)�])�kJ`��!&��*[��u������[O���EI<�8yӸW6��K��O6��@���B��N�|'�Д��(`9�7'A��`��:����W1�-C��I��٪>׳Z5��u7���%5��$�%B�\ѣ��c�7�V^�0���f+o4D����ۻ�U�ʅ��A����vW5���yY�Ӱq;���ܞ�[%����S�[E��,4���i��r�WF�cn�A6�]�.Z̋�]�h�^��o�S��C��&�e�4���C)`J.|����@;Nڡۺ.L��gc�4��{91��TF�ǒcFHWunY�����n���)M���7���/
��y��o��Wwi��..�{p��}\�gO�Sqh�ٝP;
Vd5v�t��JE�67[tL��RVw<��ʅ�^ �=oN*ݢk: �QU�b՘Sd�~�&P�1�Yw5��PF4:�f�O��0�Y��`�T��"ffpu��J���\b���9)i�Z�{�W�t��9t�d:Ő!b�YǴ;���2n��{��,��ڟ��q���L��?��Bw�ۧ�+��
Νy`��k������z�oa����j�[&Tﶀ�z�`{����Z�������"~��Ե�)���:s�µ����.��f�n�9��&i�rf�\ۢ&r��Z�6�p�1����ΰuy�����������<�=��s- ް�l��E_J�\�}rQ�LQ%]E���KN�z6���N���Js�*�λ��[�X������ 5���hD�֍j�+���ZS�x"P'�C��-Ň_BΕYH|�r�b���Zk���S�]A6jMݨ���Ԙ��(��۔�Y7��ZC�:Kk������9<X�}�o�cō$l�M'r��])���MVX�Y�b*�,�`u�9�)ٝyx9��QS�����vM<%��U�%{J�4�
�5uqe�5GL��cN�쎙%]�f�9��M�'�Gr{ڨ� ��G�.k�;�l����Ƭ��3c�O�W[���vK�k�ʦ�do ��WmY��t�>�f���*,}k��k���Q-��3����J^�ǃ�z�J��'d���`[��X�6�2��}�N��,�"������jwll�f�ճ8�B�,�@���喡9p����m�kXT3�����"piďS��8����YB�����A��K傾��K��b����H���S��-ȣӳI�mfA��ډs�\E'��6mk,��'����K��Y��Q���ͻ�;m����P��Kѧw0<+�I$�\�ɨN�?۱����=��!��ʴ���x?X���8令���,�r*e���t��ϱ����զ� tù�n���K* �n��:{z�Y�E@\�<�qkGszv}���E+ǲH�
y�3��3��*�LE솺��ąi<f���R*�Է��pz��̔Ҁ>Vd��NJ�Gu�J�������s1����03`��իV������u�wЀ�Q
<��v�N3Y�*um�}��\�ؼ2��B*�`f��M���l�=E�ޛټ{CfN�2$���k�+��:�m�N��g�Z2��r��"R�}�kA�G��z5�kwXZ�\��*:�������O��8kd���*���}�*�����J�TW�˻�5��7^�5N9�Q�ј7ծ�B9O݇s�}��Iɐ���R�z�Jy����v��V�xY��I�璭7���A��Y:��+�8+������]�sos�\���u�����Z��/-�52���˕�Cϫ��/�a���즿_h���{9y�aX���-��:��+0J=�@�}�d�Bx8>�m�0�Iβ�txn�5JXzi1���ab��FC�v�Y���St�dp���v������CYŻ\D�����`�;Ϸ.K�y�M�n�k��T�M�� `��ћj�ʮ7����+eY�l9N�N����,�{�.h�ah�3�J�%�ܘ�B7i��c��\^�y[ݖ�(Y�:㺻��S�V�.�N��zdl��mvT��-�r]�y)�����\�r�؃�s٪Ѻ��;I���_G��_��5;���hW�`��X��n�-�=EE��$5�X�s���Ⴒ')�!���!Ը��Ҙ�q�^�Z���n�tI%u����q���WB�Z��\���0����_S���C6���=�������m��cO�(Y�E�ɯDV����.lh��Kn�
��n��.�F�q��W\�t��U&�����y�s�Db^��G�|)�5��m<��*�v�nP읊��ʧ���g+����#���$CH��{�z�n���Rv]*F��5�he;���5�M�|�G�e�E�u�G���yt摚�������}x۾���}�+�u3�p��[
�`a�ʯ�Nb����,��i��'}�6�VSV��.�D�����}����27_`�Ӄ�'�.j�}���y�)�a�`>㦺�ʖ�	�MeXC�t�(}w]ggN圃:f�t-����Qvӣ�W ���3������9������g3��-��ۆ �z=r�r�
-����f����[ڂ����iHH��짶]��\0 ����{�i�k���0f����KP䯞{����4���'m��ͣ]�7�5�\o6�͡�Q-ʋ�.������3�����D�v�r"��
��7����}G[��N�0r�}.]Ż�3|�\���{��]���n=}�_�6ىR)i��[�ob�/wk�0ny�]��S��Wn5�4ͥ�+��������x��':asF_-�h�����U�h�凡|�vܭfl���0��>��]@�WSRW��u�#:q�������wL��ZBi�ص7q���K�gu���S9:�.�6�u �gCsk[�kI��8�Ϗg�b��RKA9���Qf�up���Ý[l�&���bǙ$�۳� ��i	tJ�2�����G,¶p�[;��ÙP�����H��.��u�\{N^B~�Y�H��Oh�>W�4Mk����݁����O��GNQ��p�+~��&��=�s���w8�\1�1�>�<f�����.��x���rL�H걎���m�����.]��8�Z:�0��E��+��������CA��t��(�I��;�cLޫ�ܭf��H�P�qӕ�ia9�״CR��Eݏ//�/�
������Y	[�N*�Wh��%̍wf$y��z�`��wm;�y�N�L#&#����6��n������6Fi�Ia5������.l��	���6eA�y�{�+-��ylu��;���!���>T/[-�����9�u�:�=Ժ�Y9V>�;ao�e��$%��]vz����A*�%bOL�'�.?6�ͤ���LR86���V^˛V"��\B[1׋{Ex���;�c�4<Q��H�:
	Z�n4��)q���z>��]���-����㴍��L
u8V'�Mp� ��e�v��Xjq�|#����>��q�P]�y_4�1����Gˣk�4T�f�o����oDwκ.�v��fN��QE��O�Ah^㽙�:���[2�&��h[�o�b��\0�m��1H:� p6��lّ��kw�ș�1\8;�n�o#*uEh�g���&�J�g��)�2fz���ٝ��C��_G��n�X4�J3-�`W���82k��Y��0{EZ�$�Rf��V+/���Ў=��R%�gs{�|���JM�lE�o^�Wı�����0Bk��.sJWc��5�����p�\��=���q�N�̓7��1����ıyK���\�9S`T;����Wr���:��֞ɧ-�%�e�f<GE��RU���叓����[�N���� �J�k4V�@�g�.�;q�/7�(��J8呢a��{d��\]�\��քn3�72Z�m�$��VL�O�3�<�!q�f��з�@Ke�ڸ`$!{�y}w4fQr�F�trSe-����ӢM1���SYQ3�m�sz�!�f�XD��XNB+0��nz,�QR;��ۏ"��d���-l-��v����f�+[0R]�­%��2�I7��d���-��S���h�L��n��JG�Wn�qy����{��0T[U-h��y��ͷ��������Fm�ׄc�)��u�D��3��Ę����i +�U�o;�B�
�fy+K�]BoE\B��5�{�_t|�z��v$�u	�����[�;a�#�S`���H~����C�	�o��X���d�,��{`Τ)�7ҼD��ge \~H���M˚�19rxu�����kh�F<	I*R�7�pj0���<k2޾�}����N�P����4�9��Go�c�t"��U��R<�ŕ�;�n��s�����[]�&�u�^�"�l|�=AΥ�s�xt]g	���n�\8��9:C����oqp�l����j��D�x�|�B��o?��0�2������oɸ��ۘ��V1u��f�q�kr��ɋ�59���#/eq�F�w.]�B-M���N�h�]�ri�-3#��[��r�w>�+������ձ�[�0t����I�[y�]7��3�2��
lg����,Sn���qv<v�z���o���E�MwPaun���Ȫ ������<*"��
L��Sw��o|�Ϯ����.R�ǻ@@�K�XݛH٨v[��6>��Iǘ��ŕՙ�yG�r�O{�����ܺ�yQ�؆��_����������\f&�n	RE��2��MŽ���}N�{�hU����oL�Àu�P�#b*�"+��x�3hRo\u�62��6f�z�������|��� 0�������$P�����A']�L����ڒY �m��h��b�c��a����(���_۝Z%�T���)������CI�[2�Q��+�r��W��΅B3��u��J)^�Lwt�N����i�s:P�����^y�MI3�]dux��5
J���r/oz���o�tA�������a�#C:�,i�=n��K���m��c��F{���Ŭ�O޳�)��_@�0�t7�s�m�k�$����/��7���kv�g��Z�թ�v���ό8���R���������d�Z�ކq����@�㊷��֭#�B��qSxC��̾t��o���l��7��Ȝ��y�wL��1C'�'���ل�ښJ���\�N�c�+��V�]�%Ι�k���BꡛF��h`~ہ�'�>��sh�z/km�"�}��a�Ɵ�*t�F5�+9��-r����lPSY7g��Y{��_�}�<�����.�z�8'� ���}�����.���	�)^������3]�.֩���z����u<L1�y[1܃*�X��ؽ��"�]p*2�����}Wx��j�K5��՗,��$ˇl�:�mZ0�	�8���{������_|��]��x��%M����m!+DC8k�n��Kv��5{��J���"����_SM�16}/u��V�����j�m�gag4�o^��b@erYz��m�|�53���=wǑG~�BP,Y]�^q]�*.�tv�>�ڝ�&�d�1T��N��z�F�k�H�;:��io^�Rf��ϸ�/���s�%��7C�+V�D��
�S�����dΑ��]ѓ��h�_L��=�����ot�o�u��t��}�{6L���z�kp�Z�٘QQl�����}U�q���X�wn>�ќ�It����Ze٫,LK��,J�d�c�u�:�h��Ƞ2��Z���Zt0�ޡ��$ܙ���4��
+t{��Juj�v�j�Ce\sG����۴c�fgkUyM���4O<CA�4P�zV�?l����ق�V�����T�6��;�r�Sc��L�+x����r�F����u�V�H*}\��b�ne����Ai����;t  vSr��Y��07�Aso{6e]�}����xf<��ca.�X^��s����������O\��ٛ��+��s�W'����|�)�;Ɠs�[��/��|��%[M_�Y���DD]M%KN�z(YEA'���V)�r8U�d���tHI-$*
n����Q"��$0��R��9b�;�Q@Y���ah\�3�� �TcU��V�y���GD�5
�0�e$��+6G.7S�*�J�	�ȯK�zY���&�Y�Dt��"g��r�9�Ҽ��9d]:pT��:	c���be�A�3gK�ujHI�(�"�G8Qr*4% Β(-��I�Z�iUa��dQ��QU ��eӖae�L�BQ"P۸�$$D*'R¹SN��#���J�ws+j')"�B��Ȑ�D&t��c���F�g+P�"��6QZz�����!2�Z�:�9Y�TH��EJF�udF�
:d���34�R�1	P�d�ՆQt��jA&h��
v$�Y4�3dJ%t:B�\�I21)33���;y����޼�=�2'��A��Ky7�g��Nh*��[q�-����n����9:yv;p�k�����[���H��j����/��
���D�U&
>��}�*ȇ�+�\+w�]_Nd;0��x�����X�ݫy�1��F��3����]����z��B�ۓ}���:p|)^#���#)���֓�^\fתq�f}��/,GϼwmA嘈�]K�:᪵�p9�*��+�޽��w�3��������;حΞ5��a�`����)lA��
������.i�*�OѪ���8Y9�t��Y.��_:�gS���j�����uvI�Q�5bs�ǧ��U�
~0:v�/���vK�2����]y���-��n������>9{9w$u{Ǌ�=��g���״?���P	g�]���7$R���}��b/!a[A��3��t����o�]���a'N�=�����j;::�;��w��go�oo�s�0�"�d��	n�쪵����4��0u� _s�>n��<���锇���ݻ�����B���r���S����d��M=a\�u< C�x��9k>n�Y�tY�M�S�);���Y���ӏs�J%/����=�O�0M�o��<��Dc��%u�]I[v���0k�)�����6��D%���s�!�AαJC��ʝ����Q�Zxq�G���n��ǝ|�/s$;�'&45�I�[�{ʫ4���}4��KJ�#�^KeC���]WQ�9��VYx���ONy�3�T�����o,��E:���FW�y�E�P��I�j�Q}�ɢV׆�lN)�'��]}���P�K��7��3|���8w���}*[H`0��t�	`lwg�`�r3��v߮$@�w�_~h�G=�k�6�<�}�f���x�P�ť}|�͋��9����� 8W�*7\a?e'�����5�S��?I�Tγ��F���u���I���Jq*Y����=�s�C\�XqA���?]��J�ھ��cXd�V?��cf{�Ü�hl_D��=x�x�A�1�w2��t��Hž$A�[��X�b
�-��$7T0��{��K<��-�Y��w��<���{˓s��=W�V�'��P9��Lo�`7��@
�:�. )s��w�xW�e���t��+�����h]��wl��FG�V�IO�@�ۉ<���$Ң8h�Z��4ǕFe��-��'��m5�	v�l]k�8{-���/�5L�0S��M5ܽ׻m�FQk�7v��c>^beghШ���v���mγZ�IRm�W������ؔ	��5���(��k��tFq�n)\�h���=sFզ�����qry8�_J����Î�-��!�j�x���c֞�w,R�<����Ju���Ӗ��<ϡx�#w%�5�YK��I%���}{w*���;�םy�)t���.�!$����]²P1O,�q?	�>�B�P墏N"�*R`�ʓَܻ߯ԪЌ]+�9�̩F�\�	Z鏶�H�ҁ�l8�N�U�}f��\��|�����R�-����f@x��+ @���gf7������B�K-�SF3Ώ�x�UZ)خ/6�M���>��À�(��<Ku�x�D����6�v�.`�T��p�nTy'͚{.wDAC	��P��7��H��T<~@&�J�)�)�V����;�D���8�����o��e�� 
�{����ɚN+T�I��t�ϒ���.��-;x�[ׂA��vu���3]_Ab��@f�6�}���q��z%<]��TI(aҕw��<����w�˩�f��~p�	�4d^3P��SV>��3�R��I����jb���ɥ޽����m%��t7����hݫ���@Q�Ț��`���<׫��gJ/+�nx��pRU��R�zs���Z`��!m^d|�]Ĝ��;�r��vܼ�2\�b6T��Z��S�g4e�N�M��B��J��pи�u�y|��ºvK�{�l�&��-��.����,��7�4c��N�D&F̴�&��{�3�P�3��m�̳�c���Y^����v$lκ�T����4Xje�bt�u^�$e���دztDV��*a�]�)����׵Ƶo���WJ�y�3���&���ھ"ǎ\�u�4p��Te��ϣ�K.�e�uߕn�x4Ǭ��`�����L��~FO�6�=���{��� �����Zi@l�[�ǟv}՚�1]�p��Pc�%��
K��n��x[���\�Ҽ�%����E
c���/�n�G�i�����A^��>���*��32����ǌO�`�e�����;/�e�M�p��X�|g*�a����CA���������)�ZP��^UG�⨮p[��y`�?H����4�(C��ɚ��a��ы�L{u<�>M`�dÕ�c+�#܃����ق��nm}��)4�׊o^[����@!F�ba��9���:
����:��L�Єg�Ki��;�+`J�Ss��ͣ�mۓv���h.�Cn{,X�n����o׳s^"�Nu�T�J=��3S�Z-�%��S�aY:m� *rV�5���"�)6�jG �CeR競�:r��<=9���] #���kQ���e]v�5��Z�u�+uܗϜj��L9��J�;N}<��Z9�U�M"�χyu���
n�*�[�97�ě�֞����6��`���gG�S��`9�h�1�*u-�2�$ȴ���o��q��q�ܵ���)H�K���n�;��r�lG�1N���:��R��$�e<1��ft��;�$��U%��Dh�qڜi�s�����gh�I*d��偯ߜ��+�Yq[y�Ġ�`8[PD`d�>B�����s窼5�f�AN�{/�*z;E��4�������틸�ĢO���3ׇ 3ƇTK����^�=����5��?=���k^�zV?kHȞ��ϼ� ��z���O.��y3��':���}ۇ}i$s�ǠM�g+�x|�{����K�S�=���И���^��2k!������p�W_��!E��v�J�3��p����Z>ڼ� ���{�5��D�wF:�gS�����b�1�O�]�s���/om���Ή[����N����pi�X�����22)'�7<{%��O0w/<�`����`H���mTȡ�ĵoh*^�ɇ�k��ܩ�O+�X�^�_2��H����/����F6�<��Cn�Qaf�Y"3t�;yے0t�g���r�jT��t�k�����d[����O0��]�Ǧ�Ы�"��K@�/����A:��ú��*�t}���[��wZ��%�;[ұ���>=3���l��+��8qŗ���K/��Eϝވ7>V�]��˵�N�;�>*?�-U�^��j�^`d$f��
'׷����o���&�q���=��!Ŕ���ߌ���B��Ʃ�4��ȯf����;�g	z���RYzpj�������+���k�';�`�̮U�{�bi�E��P��~�uX˧?NÖ4`k-+�r<U��TyT�;k��_�"ק���ܢ��F��֊!���ۯ0]i�_>�}j��V�X݅�r�ef�
r������� b�D�f�!B��Z�/�q��]�<ׁ��	R�A��ּ�G�z��4O��נ_�]'D(�Y_6�崊{R׀���g�y�6�m����_p8��)����O����T�'O�AݺUu4�%ŀ._*3^mWx� ^��w���Yw��ҬW��	;s��F��N%K�OA2���J��CɜPS"��]��//XR�d�JX(_�78�r1V�>YY:�
5η4uMF1;DV+�N{���FB�yh���5vwAz��(}��8L��	~���'d�g%H;^Ø��]�=;9.�Y�<ѵj�)��8;��ps��fe�t�O(^ܼo���q�!�+fӈ�����yGD��_�?s����J���kp9����X��4;��d�Ŷ=3�.s/��Ɣ��W����KԆn�3�񅺛��},��c��ʔ�߰s��n�g�{���<�c�g�J��r���Vg�{;q�o�,B��W9}N�;Jwg����9^��7���y?[i���T�ϣ��U��<OhU ��=�W{-R�\7��b،���JzO����䏅_Z���X�6a>iL.�{P�l�8C�^�+S�Vڽ��~<��$��8<M':��<��L��:���h࿮"M"xy��7��o+�[��Jc�'��Ѥ ���e¢)��r�O�dϷ�T9i�ۤVج^�P��W��wo���<
��{k�F�T�j�(M-v��C�->�M\=��"�Zc9��3V�[��x�8=�x��X�����@��uם�S��g/�x`���j}[�0�e�z��E���ȱ�>(�P�cp��|��΄��Y�C�~�w�����K�8����M�]�^
&�㞳G����턄l`�*�Bs�1���*�+�C{7[�9���:ϳ��	i�O�ǜ{��|u�-�]�W"(؛�1�I�m6$���0"!N�(���u�����VelRP�5�#�5y�G��c/u��';�o��Pn���%�9�]�VRuĒ��0��n�x�/��d���.�^�{�Ӥ��-�I��zUi#=XV���'>�����3��Z��@]	��N�ŜF�_^:1�w���ȪE��6�}��	(q��%8~%�uTYȤ:��9������r����R�P ��=�guMX�Z3�����nb��J}����L�l읩wg����͢Ip���]�_��c�z\՞��y�1�͡�x���^p�#�m��=��s�-C��>�	�CN��O���n�g]z*���CH���=tV�5�.���d�Z��KV�����ve�<a8���7GuԿ�?CtҬ��O�rl7s��oe,��X �^̿���6��Nuׇ�z`����٘=8�Ux~|-	p����$=BeW�v�N�&��mz|�ϻ>��VD�<lt���ֱl��S\q(}��`n	~��nJ��d�;bm�E
�n'ௐ�u��p�8x��� /�V�OE�6m`�]��B�N�/*ܷ���:E8��W�w��	;��a�7e�h�9�}�Ö�7pɓn�z��a��i�o��-�u`*t��S�;����;��p��`�v��6{[��R\�w"�yפ+̎t���%]{t��tA�̡�,L�����~q��+5�!��LD<��*LE�)�u:��1��1����X}��4 }t�@����|������W��_7N�:K�q���azx�����4G�'��(m��UlϞ�KOh��.W�$�_3�u��|:Y�j��>wG��=�0]g��c��p.Ͼ�5���ߵ�7����@rh���!�x�WًBDmw�d*t�K�2���'{�.Qw,�B���:�I��>����QDP��.ḱs"h�P����}0¢�z�9�:>b���֍�T�zZ8\�M��fB$�;u��ck[��Nص�R��r���>곗��;��)��[2�\�P��77(��<g3��rl�V�����5A�5�A2�����^�ffǔaϢ�_X��K�dfC�.�*{�ѶM诬��u�G��(M#֫�q�w�u9���GX��k[��-���HFKGD A!�a��Lv,z��}������G�^[�^�������ҳש;���s{��]]We<����6���/{�Ф�t!��#4��^.ٽˮ����v��.[[��
�Z�6�0l�o�+G����]D-���Ο��Y]O�i���V��	���+��m���Y)ֿ���U��:^�2�\LI���fg��L`i͈VӻӞN�r� z��N��ؖY�
ઍ�:�����]0�r�A�1�B�;����-��j����*w�xN�q5��c��Ɖ�(Q�n�-��_��ڳ�ڊ�O�e�X��%N\o�__��c%Ҹb2N3����U5A����uuy�~�=�Q��x��x���Ъ�w�<!D��� ���ž����g��b}�˞΁Y���+룴ttg����Z�?X�|*3�-�`�]���� ��j�����vҙ]�T���W��R��7��r�V�U�mft��0��:k�暀�/�Vn���z_�A,ꞡ�sMh���C�p��e��m!��IjL���u
���ٷ��Ty��i�����"��X��r�t�����v���π�lmT�w��x���9�i��oMf�k4�����7�9_z��V%C��>�f6��u<�~���o�=
�?Q~yIFb^ʽ6_���� ��#�-���K�!�><%ǟd^��y�>��Y
����Ծavt�70 �(s�WG�t�����A���J�1�7�3��v����Eu�o��c�".�v����"v!�u�{��R+��u/W�A'8L�G�i�`ܱ/�T�5��N!���]1�ⰲ�:d���Ⱥ�qH��f�:�;�:���@�9��9�����.U������V�aF,Z��7��z�j��� U�Y}!�y��!ȥ=��2��J>*��]���ݗ����ӭ��޲��ԗ|ͦtW.�#.2v��6쥀�A:��ܑ�-�%�P���O%���Yx1e��%�J�a^�����h�F1=�(f;.eZ�z+ZxX���FYޝ��a�;�,{Rvoq��k���IpgJ�Ɏvp�� 6uS,7�/����<�;|^ɚ5����"��M�ۭL>��H}���k������o(7>L1���^�!׮�ϰ:��ث�tF��\P����\q�k�2�����7���^�hB�=n�җJ���k����F_y���ڒ�$٧��u��6�V��p�u�r��#��D�0!HQ8�Q�Q}����ӂ��x��)[i�&���>A���\�Ƀ�mq��v5�k��zpV>׏jH�8��%k�[z��؊����c=�z�=iJ��giKif�y74�q\��X���G}g*r�k�
�V����.���ɍ���*;\b����Μm�0ܷ���s��Â�㝷��l�Ě�ODNh��*j�Ѵ���J�V��V��]���`�N8X��B!!�j��*]SzMC��m�F�
�*���:g,�H��YR�ˎj�k�5wT�y���݂V.͇�j�n�u!\��E&Ya��q�6��LM�h�r�M��ВU�T|1���l{{h�:���*Vۤ��-bIŻs[� �D����S���-xg!�Yڝ�[�z�W+���yX#�OSkv�##*����{��}���n�8z��Xq�׈݉j	(b���:��t�I5M�9�����'�0�Y��ݞ�B�im(w�ި���g�0�%\�i���旼==��Ni���d�u���w�Q7�=+h=��a��O��C�-�Q��� ����.��X�Cs}-���1\ɬ囉=<�g��Ǔv^�|{ĥ�ٞ���ɪPn�iYyI�6�	��|=���E��������4p��<qnO��Sp=�]v�,���*�[ӈ��X��Fe��@��IZ�r��},�b����!_�t�U�Z[P�[�u��V�*���=��N�X���$��tn�긖��#�;d�׺ekE����v�V��G3.c��l�]�v>�B��ޤ��o�)۠��0�D��ٹx�������� #4aZn��s�s��(��\�ßv�V]iJ�=�f�]��86��ρ��.��b�u�*�b���J�!30�#C|�9	e�Ք�*X�fuYH�SH�"���M�]%e��a\��+�!sRQ8r�Mbʮr�J��jX���,��p���3�T�%�*E&dhu�e�a�U9V(h�#9V��@R��%G$'2��ir(���^i(��YUE'�m!P��\P�u�$�R�B�e���΀���J[U-j�R��S��D�MC$	J��7P�gQ�*����NU���Ea˩���̕+5=��l��*t��U�Q �Ê�p̺vS*���\�s<�J�J+�r䦰�:l��1"�U
���JF*�h�E�&�JB�#J����EkI�Q�w�.ŨY���(�
�Մ�Nj�J&����"�P9rJJ�Q��ei���VZ7S�EW�Za-"�1>�T�";���2n�oo�&~o�ڥ�����#�`�L��Yֿ>-�'��SY��(7,Iu�n�w9�-^��<�{��ݞ[�^�#����@�(��
��=��P�����:�N��C�G�۷'&ǈ������P�=~q�*|v�F������뷯}x]�� i�����>?C�ȁ�{��c��O~������v��M��v�!?�;���xw�[�ߠ��OI���u��~y˾8�G+�M���:=�x�����=��yNM�����&��(npG� p����M�̹{VOE������[[J�T��DE���@�nv���~O.��u�&��w�ߐ�;_)�}�$ސ�w��_?cxC��?-���8\>��&��������¸7_S�yC�5������N���Nd�mwB� ��E��D`��;�����P��w��x����Uǣ���nBpy=}�c~C���������\N$�������M�	���n_Vܜ��5d|T~��dg��� � ~��ޓ��5g^�]�H�1�h��#�g��o��p>O����I�!z��{�}O���`���H�~��~����
#�ǿ�<l����9߿���bw��=￨?}�(�����_}V��@�-�����̧�w��8轼� 8�����90��N?j<+��������󿝤��\P��v��C���c�o�O�o]�σ���;_~����zL.�����ؐ��?�?h��$�#��?T�@*��M�?�.�{��!��(������<�����z����r{Cߣ�<&w�5s���L?c��/����4S���u�!�=�����k�z��ϗ��z������o�s��������&�뮾�E�_�@Y�����xv�'�w�}����ǫ~OI�	�Q� ���s�h{�������t~w�<�w��zC�o�$�|x���7�99���@������~çD#�-�m��P~���|�H~�q�/�o�ɹ��S���x��~�y@��������ݧw��?��;��Ϙ��]�&���z<X<;�o��ý��������ӏO�9��wʞh��1d���_�B�q} ����ｃ���ﯫ��4�v��o!��o��ۿF�����aT��}�_�p|BL>�۽����;z}�'�o;����������9Rv�|B]P���a�=�~q�?>�n��d{yt�I�'tcB+h5�ʹ�dl�ÄQ7[�49�^���r�K��IsG�j��B��mJ� �%aWs98�8�ٳ���iGȱ��;��ך�MQ(T��<ûS�s�^m�I��6�j�ǧhu�?�_|�);)�[w]�Xc�#�E3G#���돮�h�r��v�
o���~v���?x��~q��7�s����xw�����q�I�n����Ǵ9�Xj� ���!�������M���.�����z��7�����u���Mվ� ��g��C���z���,��<����E���Ѐ��DB>d}���C�H���nPgﾄ#B�?j�ʢ��?��}���;��QC�ohH~?�w�܇'?��u� }I��ƻ���ߟ	�!'��p��S�z��{�S_��o޿x?���@��{�ߝ;��vs��D_�c��W#
6�x���<tJS�Z�c�/�Y#��#�#�~���?Q����<��yL.����Î~�ɼ�
��㧓�ĞN��Sy}�rr��˾~�ﱿ���o)����=돐��@��tNy��~�Fg�mJ�5�_}� >c��:#�~����H�ۏ���o�O�nN�~�c�i	�O'�S������u�?S�ĝ;To�9T��&>�}��{v�7�{�,�g�D~#�/��j�1��M��o6nk��.�">��x�(��~�`"�$'�߼����9��[���/����{��=��;]_����Bt��<z�I�<c�xv����>�<�x@��y�>�>�>#��ztu�ώ���VpoE~�??~���#�G�(��|�}���~w!����raw�<���������8?~�7�$ߐ��w���o�rs��< zIĞ���y~���O����C�E��(�^�����:����3?E�� x�����H����D��,v�����c��o�s��>v�}w��}����F'~M~���ü'&�����?'��C���q� (��?>�_a�������ڪ���ޛ�%rw����MχnNO��;�[w�k�	����V!ɇ����㷕w��^?�S�~v��'��㰦���v���<G��� #��}�=h|��)������(E�t_�Kaf������j�tD���F��~ǿ�����a|����]���<�q�;�s�O�<��xL.��z׎=��L)��~M��q��8�y����	2�O�?��������|v���}� ������{=���3�6�#8�>QN�v'o�ǧ?�m���V%�ܥ����ҏ^n $C+��5y�:��B�n���h�ڝZ2NP����
��Q1�-�}饛o�g,���D�d��+��gh�?3�J�����+p=�N=���W�x{��%z�|�
o�����'o�x��?��<.�� s�����.��!�<����É\z���}NNC�ǜWz�N���rI�i�0���ޝ�ߝ�v���o
�� ��� �����՘/�f/R[��#zC����׏�ސ>�����<bO��oτ��}�ǔ¿���z����!�0����q�<���M��~O�:w�C�xM������&��O!��?��G�~��R����r�w)���D�?n����y�������C������(x�����I����������7?��;�<bw����>���S
���,x�����<�r������~O���}���9[ߓy׷����ﾂ�`'��xO
�Szw������;�1>����b_}��,���>��?|�Bz��w�iP=���|�;���~��yw���뿎���raw���]�=!�O�^��߳�*�u�W�.���`����`���ճ�	2�'��u�Rw�
]onܛ�������]�{���!���j���~�:�ׇ�O���|��~O.?8�޾��xM�?��ٹ�����s<F����A!������>'&�����ÿ!�=z���BM���S�ߐ�Ǉ㷔�;ן|yq�>>~|8|�P�¿m���ǔ�P���/��m�=;۴�8�imeD��yl<�]w��F�ﾺw�~��<���[{O_�w�p)�;�ϣŏ(x����X��q�������\rs�~��ׄ®�)�������_?C��?}�?X�~�?}&�*�V���85�]wKSF(�}�#�aT�~���o>�!ɿ~��?;r������y@�O���}߸���7!>���Sʸ�|�|�rw����N�m����'}v�=j>���W��YuŎ�,ڕ൏Ew�G޳������ϯ&'{O�9?��_��zL.����9>!�@����ɧ��;�>��c��~'�߻o(��;��<y��nM�<����u8�|���?|���@'=�>@���e��nt�1��;I�x���˅��7�}�	�����'T�#�!�D�s��4>��3�����(���j������F���xW�N<�w�<������x��!ULQ�����f��6�Cֽ�CD�����GC��͎ʕ���.VƤ�������Vwmd�gr�a7���`�����|������P'��zu}�&���7.��k���Gr�iR�q!x��7�d@�ZW��gf+��\��I�ۋ��x�@�+��u�����\m�vy�K����,��o�����	�~X���r ]�_�?|ȳ��F���E��ߏ�����xM��������p)����<zM��bO���~M����9�X]�����Hc7���Y��r�3��0���`���G��	������O�o��n}��V��~��#!Ʌ�x�=�_�xC��շ}��ܮ��gϜP>�����}����ߐ�_�獼�+�B��v�p3�*U�i}�U�B��#��ۓ�[~/ݼ;�[|?מS�;Tx�`��r�v�,ro�;�kw�����Q�7��]�c�	�������c»�i���z��Ǥ��	��ƚɓBM���T�EOF����߿}�V��ɽw�:v�R����o�I;{{����c�.��!������ɿ''8���\�7����wG�o��'��~w�=��}���gcޑ���̫���uv�H����;������
����ݽ!�0-�'�`x�~��z~�������~|/�P�¿��p'�ސ�z>A߯�o	��ɥ@�����{:���G�Db'�zf�r�X�o�*��>j�Syx�O�ߐ���޼��|y�;�r{�����s���=x���®޺]�@�F�(���|0���Q�p�+��=&x�o[��{C�<��T��q��DH�c��O�I�5GA����G;r��������+>��'�>�4<>���ǉ���0*"��#�D�WF:�gq:��j_�rn45�7E��e`}#��w�� ���X�֨C@�q��O�CWd��AI���ԛǃw��K������_f}-hu��i��	��,���E��g�<M��f��0��]޳N{;�^�#��tʄs�|a�u��n]g�M%����_ʝ�u�"R��<<p�����	��QYܱ+
^�O�vת�DRm+z|�%��[�(iw�.� ��ح�V(�}Ӻ��*���o9X\&��{��SfF1t����lO$^����L��W)�њ�v�Z�	+X���Z.�����R�-8���r����#���{^�r�ŕK����;����	�C�p��e����
��t�i��.����8�1[ە�=�e˶�2�QpCf���'(Ҋj�W�����J�xV���v
=Ӈ��<�#�hq���1��b��]9�Z�N�mh(�x����fE���Tƞ��;��!��Qh$����RR'WG^��H����Tw��/j��m�]�O�f�~�&9���`zz`4���@�\�n�5�Һׅ�3}���ltE�t�D-+`J�ߣ������$0���%�92`�(�Y_HF�-M~f�)]�dߩ�n_��+W�y���؉X�_=�	<C6O�wn�_SK���Y������(ߟ	�7f���[kuNM�_�u#>�N%K�����a��!�*A�����Np��Vj]�G.��}0|��ja���g�U|���t�n�K���Y��~雉B��؞7t6�1;`ލ,���)V��@�����!<�o��z���L�:���++g��P.����y�Q[�>���Ym�D�K˝�(VZ	فVGW��ǝk�gT�#D��+i�Z�y�`�_�}�	�گ��up�ƶ�M�ޫ��X����W����G��y�l�[ޣ|�oc���Y*H�^	�d�S��t�wk�&r����W�WՋ&q�{�	�_��ì�k���_I��
�a�����@�:��fb|�<9��U�z֬|��"�vVŰ׾�Ln����~���(N�S>��J�Y��nt��G����$qt"�m�����Q��%��ɵ�������kԅ�a>iL/���9AE{��gox߁{ԧ�e�`[L�*���tS�_�������6���}��C�><���Zw~��ͼ�{^�<���%W�\aa쿞 v\+>�S���ɟn!zQ��r�ty�k��^�g+1+� ��*�
����C6m�T]�T�<�f�K��z!��ϥ����R�>�l^n�k��|�"�9�$�¦M|Wt�8UwK�����}��Vdy=[��mM����@75��0�у��㎥дa`�'Wʃ%�Խ�C�~�w�K�5�vߟKj��:���=S�&�ʀ���N$b|@���A�y�a��E��q��˳���i�E}_$�#�J�"E�ߊ���'%a
�uI>X��I�͏1��U����DA^�Y:��I͔Ӫ�Im�%@F�+�K�ϴ����1P�����:�;O3I�v�hÄq�(�q�#�t�ݦנ�k��{6u��\��]�먻�cS9���Z7բ�<=uŻ}h6��[Mkq�RJk6$r�Exu󓤎���}��_S��<��y�S�9k��uܴ��ʤY��Hm�c�m�h`3l��`��̌�\��A�M�+����С�U%�#�֪��j��s�h�
r�B�m�T�IB���xv=;*���P�>��"]i�<����2�ʬ��oA���|�s2��F�pu.�o�4n�qk��c�H�TV�J���~�6e�Z�]�et?^6>��$��D���� ��:��l�u��
�Y�U�A�,�O�Xµ_�ʘ}vЧXa9B�x��S�?C<�a�
&��3���F���|$L�������y��o�Kt���U�TE�P4�d	��z5��'�{'fu��ߌ�;��,��I�����tQ(��qǟv��`1��5�����\��c�L�,�	��T�Z\���1�Xu@^|v�"�u�B��n'�|�꯮N�Y�޿,vw�A�;�]� k
��!���*`�0]2��:��e�0o��9��¶ih4]���{�֥̏wQ�A2����eSVA>ߗ�*�*�g/m���v~���بG�l�f�r��'�8f��3nA���*쳓+{�^��y�ϱ�^�FSBڄb�)��fd{0a�����)m�7c����j�e����E��O'H�\��|Q�����6�}��T��@!�#32�2�l|ޛt�um��{�>���iƾ�I<h������孴��4
��ɉ�2�7��Ղ��� r�+��N�U�Fr��m󡾩R�vc��1X������R痾��CpzY3Vzu�����P,�u\��рq���z,A<˩�z�ʩ�hs*$C�Ǒیuc�r�qeEܸJ�j�r��Z95L:���8��n��y��Ȣ֯R3�n�5��B2��{kF�m��s�������K����l��q?[�jHe��_tiy�Y���؇|�f|�/�����-Yg|1ʉ�����'�3M�wD.K���(Jv*��[T:`5�A2�����^|;���lyF��nt~K2rὢ�G�j�/ 9`kϠW��tE/��'X(M6}����J�^�ee\Mc��θ�d��ub��|=^���a`,/~*��v~��'h����c�d����՝�hw�[6�VT:�r�s����,v|�����&T�����=iX�
��\|�~�)��)w��]���#��ò���Ngx)��_
�������q5��L9{����dЍ������}9�r�y+aYh�֨�sF�$�8�s"�^i~j�\�fe�92����׬�fitˮ��?IށJ�tl̫�=7��tޔ�f���ƻ4w����4�Nv(�����m�jn?Gg��/3]b���m�˜�gu���������úbX瘤0���Z"�����f���7����ƽ}��5����o��M>4����Z�^�z�b��b�T��0e�>�2���(��т ��_x�gݺ�;��S��x����=U�ʗ�6�q�g1�G�43�xW[��	�d� �cnz����'m�F���|f�!��]�.گc�~o������hc0��@�+
������;��v7PhLZS�+U�&����=.j�:D3�l8���ެ�=��HP��KGJ��:�LF/{{ws���d�s�7>�wg�<���5�<��(�-?C��'`g���
���H�����6@ p�x�=)�1Uc8���QXс�t��r<yn׳�6ҧ(>�j����	���3�S~_�D�F2������E�"�No�^~��JY�j��r{:ת���9}�zKˁ����k�-�������\=����e+`�r�o���\��Z�I���T���a�Xr^��d�N��Hp�!)���@k�L��j�g�wM�Z~#�������Y��lA=�&\�o}焌
U�D.IZ��l�=3�ܟ`�9��e\Ғ����"�#,d��]c�ˡ�v�r�+�S�n����4sƁRg*�|��xv�Y���Vq�h�]L��k�uidl�tc��| �˿m�K^�^��g���lnv"V$��O.x�g	�ۥV:�_QE��=}A�Ϯǌ��i�p?<91�ߠ^�f��>[k;�r�����q�7��J�|�z{�g�r���ھ�]��\�ٓ�Ѡ;=�X���Y���V/<����yc��3�'�kkrxm���"X��W��U֨~U圁<���aV�{]q�5{�]g��<�,��>�^N��W6�'W]�G/�ޫ4zeV-���+�b��\WaG�wl�c<���{�η�(�������U��g�՝�ᾯ��tsSKw T������ӾRT�3����wc�d��� O�y#)L6M��ޮ�Z+Y���4�'��IL.�mU����g�����d�?x�Wp!篪�bZ�tS�����W�(q�+��X�2��3%�t�f�w*Q�� z��Vj��mWU��!oe���V}(���)�����f�.h��{��O�c��ճ��x��"�*B
�־��{�Mc�j�}2�q�ϧ�F�6���m��x��D��Z�e�y�ڇ%4�%vd�}V}��L�〕�҅}��Q�!�va���b��h�U�VӚj!��Om�{�b6�����]�yg;P=�u���Mm%/�>&Uc"~�)�r����*�f!���.;v�5V�s+P"�44}k�`ky�x(�Y�!z6�Y�c�c3�e`� S��,��g))�D�����m�~d�rYu�[�'}3F9����a]����R�%w-��x�Lw��Ů�:y�tI���# �_nų�7J�����KU��#��:_q�i�za��Ĩ�� ��b�e�� ��1De[�Q8vKq
n�w�ZnT�hB�h��r]����[�ln�ع��+��p��$ͺ���#�/�^<q>��suk�jރ|��� ��N���v#��W���Fs�Ioӎ��hRe�]
�w/N���7��^.������z���bi��&W�j�vN����*���ݕ�z��c�/@�Y�È0�+�Z�3l�YI5��C&��=G���k�΁��lF����N�����5�h]�5�1��l���}j�kV���4-��w��Np�����D(�vt;]��K�9�L��p���}�w����":�4�i;�5ْ�&�x���ufb靶���w���Z�������e�X�,��FrGc�H��f)ۓ2��j�XN�ha�"�q[���T�8܎_f�$��(��`fS}��H���r��6���M9�{k��#[�W.��u 4$��Cr�l~��ǐ��s�st��ܩvV�r�X
m��(꥜6KLa����L S����;"�Mg�H>�i�UmkU�5�;������F�%.��׷��r���ب��޶x
3y�y�(����ŭ�7��`��a틟ʬV��F��}(��=��fg�$Kr��e�9�f]4�a�2w[G�IM!ni��P��C��xH������م	��f�֎�˳m��|ul��d�'\v���/��Ŝ{�R��T��3�.�B���`|�t�Su��JĲ�^B�]:n����UA�i�uM��7��_��H�2��"�k��[�p�u�֍E���*qp��bD��f`���lґ�L�UM��<�c|bzcWVl;=�_=�X�H^OO�J�c��#i�t�N���X�_i�ْu+|�!u��12z�WS�Մc�S�,���twA�(;�#�F���3`gDC�=p{�M��V����y�������A���#��-�����)J�u�md��}��k]�U���r��oT\.�];�${�e:Ȃ�W�7�ۑ�{vي�19%GwL�a[�L���z�8upl7F�eu��j�c!�nF�7mۂi��y)�m�{���+i̽���8�)��)X�[�y=Z�br�eȍ�Xub�:�|0�@�>R�Y�(���N-օ$fuH8�դ��Y�KV�V����EB��Unn�r�Ή��!4�u��!P�V,�b*HX��XdQQ�(�U#�f��j�D�i$��������UEr��R�%$�hU$G"�N�*)\Į�I�;�-%�*���eQQ$j�)�U�Ќ��Y�j�����ցt:U�dH�ՕGT�u$��D¡K����縐F����m���*�Ƞ�
�,�9B�V�Qf���%4���ru$%K:˜I5e*�9B�j�HjT�S=NT�VU��ډT�B�������V����BT]2N�������&dI�-@���R�	��5�e:aM1a)�uT�����/�!$A?�@ow__]^V���Ļ`����j�jV����71�	��JS�;�:~�7o{��XyV<�������������]yjn��n�����܃6��(F���<ʀ {��jCq�>�޿g)�F�O����P�1Hk!w�|8+�;v���~�A�MޤH�s��q��L��g]����Jh_�N�t�����vyp�fyP����D�O�� �����;��~��l�.��&.����CO��etOw�D{���7-��*�����X��'�!4�|��l].	��b���U5 H�=ˈ\�/��Lߎ�ki���4C�2^XR�ž�.`���3Յ���B
�Cv|z�l
t!�bg�KG��3?���`����\�	�C$펨�+G�\��T��u�}_m�T�-Nu��G�7�����	��d;��nq�,Ə�(όhʫ��4�:������JB�;�����uן�[C�����vCD	��F�*�y�3ά/��L>�hS�0��c�t����t΄��-�ꦕxV��9�T�<s7	��j�'?]xz7��\��������j��u�z��0q��J*��%O80GY�η��&:�e��S!9(���n������n;u���D��t{/�����-fH$��d���_.rn̅|^���Ot	���Γ9j	�jJ7{���� �d�w�$5���N�s��N��������_n��9����џ�7�!0� ;�	��E�n �ϻVj�Ƙ@��z�����{��I�	1A���.�ᎂ_y��g��!�%P�^��LL�A.�oI���_��Ps*�������
���V�.�CµD!�7����n���I�ֹ�sZvq��� .�C�T�;�;�A�1�R�՚������o[��M�����/�������q��+��	��q�Ϧ���<-.^��N�T>��0�ټ�:�Քk���<��Wz��]w��~��Jw<�#����f��ӭu_=*��w~�����2�+{�s���̨E����;ü��bڨ��J�j�mE�dc2����%��*O}X�7٪��'��
�F����`�8������l��|}�����~o�8�x�����VJ;�|P|��~���B�y�НSf������5�c@="��/�H�! �Q5�O����(���'_�*�X]�����/�jq�w8=�}^��_�b��J�{:A[I2�Q�$�d�L��]���������Eά�Y������}oz�ڬ�-���U�i�Oxc�9�9���X���8H��$�W�b�C9�<�=뜱c�I8x�gk���?��+�h�Y�WzO��X��>�}� �{�\�r͚�8Y�?~��L���^|+�a:�#B'� �4�Q�:t�<S��X)7j,�xļ40��02'L�x8�)`�m�`x�*Ňgᥓ���~�F�M	k�o|{J�+Y�_V�YM����0�Z��b�Ό�ʠ�غ6��V%�o�o^r9]����i��AZ���n��;������;ؼ'W���⎍  p�_��_{�̫:)�ϴ�5�ׄ_X%�X�΅r�{;m�c6?}R�E���r��쫙�.�=�ҁ0Oi��T����(��+�`VV����꽱�����}Q��7��F�g�U8��;�`��z��`����f�w]�A�ny�����'e��ߪ>4B���%v>����u��C�bê�ǍO��m��BN�;Ǻ�z(�~��w2��ϧ�(4��cZ���J�L�C=�i�������a�p�`�\���̾^������l<��N8��!9���H�.�QC��N^ҋN}��>��pq�'Z�L��Z*{6u�X��=��|�3Mޱ�,��K�T�}s5���gZ�O<���`0�<Qö�+�n�hun�e<�e�EK79�D�خ��ݸ�g�4�vZ犂�
����Ӫ����sޜ�]X���aJs(��vOu_T���������$�tＺџ�`ô �L]⮇�#���]9�u�0[^v��3��+���_@�&y\�����B��t������!|�M$3���E9�|4^$���.�-l�:�ҭsZE����2Ǳ:�K ������Z�[��jB�����۝S�>�r���m�7@�Z��m�񒥴�|bNJ�;�ɂ���s�~������Nzel�r �p����K����y�3����b%bI|T�����,Q��u���;��_c�τzE�x����#���ćY��9css���a�N%K>rY==��#�qe\�u��z�~��[Dｔ��8�)�#��ΖM�ʣ�i{/.�On�K����x��;/N�XK����A?w�l�3
�uƀ�B�N�
�2'���R7i��mx�����O�ծ��!�Ww!������X�0뼷4� ����B�y��������Z��['ap&*��x����5u��9������'vʩ���k@���ϝ�����V�ܶ|�"���"m'��gU�-�58������h��y�+�DV�� �EՇ�o�[�N�?Jg��(VĜ�k�n�&#hq���;T����egp��1���ӗn%EtR�0��FǵW^�Ս_&�J�݆&M�ߪ����Z���_�ЇD����� N�O$`�BD�J�&�}���vV�ͯR����S�{h;�p�#����幜<3�H�ve,�hꀾ*�k����ϡy��t߲��8-�_z�9s��|�*q�+vI4���K��~J����_t��l`2��r�[#��P&,ز�A[�2�~4�:(���A�`�>�k�^9]��1�Agӽ~v�^7�}Sh��Mee��� '��ϛU�m���Dq��D��ϊ�G��yaBg�9OOn_3�[���w�T��ǫ�h�'�4�Gˌ<V-݇��&���IT�$ZJ	s�G�-�W�M�X�OP��76vτ���J��[��g��@��L�Q# 5��Vm���Qem̷Փ3��u���|��G�_�x���r�Yg�8_�M� �,¤�+Vq��|�:��4{Ƨ�鵟$	�#u>Zw�qx�C���%,P�!�+�)�n���7~��۽�>����:���z��AU	0���h�g��j~]��pP�������a�;0���ڏ���ۣ+TA�7QΕ�j�nf4%�� _Fn�gp��r V]�����g6�a����y��{��e����j1����!\��뮦���`��+�As���aN=��4o��޽������ޕ:"�ڵK�r�نX�cjb���M.���o�*js��?i�5W��ʉgD�;���ysƍo�g�ve2"�9P�Q�?eo��^�Ն�o�n��/,��WV���W[�����,���LgNy^(r;�FN�2��X>5��
�n�D`D�|�e�\F]�^�dё�]_�?x��*�/}-��Z� ngS��6��N\~�𯷦��?S�n�<G�_3�
0�q�����4���(�U��u�Q>��>1������w}��q94�N�FW��p���^=��f�����e�?mD�Q�)ѝ\��/>;ba��T��}y=w�\�C{\~bu�ߨ�5�q�a�p�{���+LL��N�\b�|����p����Ǿ��z����c����9N.���8��5����	��*U������y�$)I��<ۋ=��O��%�0�9��Pg'ޖL�/��®��UgPp�}Yc�!ω��Xw��l�X�[ǥ�J�_:��s����z���۪��("{�@��ǯ.'V�����4	�6&]s��͆�6zp�o��j�A���]t���e?jn��PF�,̾��+mWq/��mM䙞��%G�[���Vܜ��̇�{A2WW$/n˓c��q�z��ZK��b���l���M��6/��諭�����~�fxX�~�|"�)�u���>#�xEܢB��(��2LG�:�O2yo̜gsF��b+�^HKh�>1jG�S�
�qu7�ʏ��ρ�^�0���3��On�f����AW
��ۮ�_��Q#"�-}�B��&k�}�5P�S�ڍ��{2�V��V����r����x�c��*W�Dv�Uް�4tyfq�MP�z�"�6_��c�9>���0�/��q("��f��k�,"+�KlE��=b텝�M�{	Yշ�Gviz��K�!������e����7X�����ಬXv~�Oݹ��'X|<s'��^�|ߜ�8z��l���k��9�N��7P�����'@9s��~�Byv7=��lؒ4�N�?UW@���qq�絗����
���4�����(��k���0<}3kד���w�;c(�_V5!�Yz|M`�=�C	t�3����� �����[P��9]�%�}^�d��^�g�{ɍޮyƳ֖����tU@�{��xl����j	��˥��,�{Sx�1K��n���ƴu)�|o��h�<ݹg�G(���J�Vw�q��
K�p�5��k=�o�W��g��Μ:�6`�쬰��c��p�QV�x �o62�)\�{���=�k�wu�L�*�6� Tǘ]J��q�͠.;S�]��}i�ŏl�$�������-���\w���8�3�����hg����n�M�Ӟ���C���m��H��7$,:��<�!\:�{&���]H˫P��j�G��W��%�zL��&�p�����!�i
i��0?�5x"��5�~�����w5>ߋYw**>�M��.���a�`��e�!�B���F���P٫�s��4������s ��*�b��e�}��w�.��/Ǭ.�Id�=]`;M��;�E�2_վ�\�rZx�:��������z����r����~��A���t����
Z4�M$3����-�4�x�o����e<W��T�Nh�q�_�_���u�M��0-Y񨾯���-٭HUt���{ؐk���܂c�WBθ��`�:�xϾ�-�0|bV���&
�1����IO>��W���nR"
�\�Q6�87�Cbs67>�b%rK�}^^ h��q�Y�=��{������.���Z���ЏU�~�z$����:��N%K����H��^T!�6nT��6-��ӹ���2�Q�u����#E疜U�Z�SQ��kl���w��O�.c��ku@�AX�_;��b�7����Y�
r��GT�z�'�^������Kb�,�e��ҁR�M�h�3g_t��N�/G������9�u�d?_(3���$�Ǆ�z����G�3�+���|Q�_s�����'C�0n�/k3�u�Lq+�J+A��n,�<�� OP(>7����^A\��?�ο��&;�t*�u��Ȃ���r��5�:�?�_˦ٽ�\����#>�XHW��K����g%�[���^Ë
�:glf�_�/,�S�|j}��9���_��w���q�V{'���4N1q����*_���.2Oc�g��H�J�&�GZGq�{E��R��4)3��u�V��Lߔ��{佅�r��;U֪����Pį�뢝�Ogм����t�Z��g��;�Pf�����I O��//n�Pϻ�B��<;.�P1O+�g[�r�
�W�ܸ֕݃�����+��<[� �0 k_Z�봡�j�Sެ�Z�$�^T�=睮(`1��}�&-���;�VE��#��y�P@�y!uG�Hc*�K���I�(���.:�x�/o�=f�{���-�|���b���xRj��uA����Ӽ���hV՞�<1:�����]�te��E�v����MYE.�.c��j��u������ʖ� |��Wlٌ���yε[]7�t��u,��NOD
��gM �n��h�"7*q�\����ѹ7-=��_WqzK�:�� �ջ���\Rn�${���e�����/����z�-���^yP��p'U1N�
m^����m��A ׆������>�DVqM��i:H����|_����w��f��q�9�,��'�vb�I'�+���(ȸ������W$6�씤C��5�����M�+�z�'&���	�Մ�W*�����ʨt���b�h���T���t���7�VJ�W��}��ZWHA��T�Jf�`�-R^�����V<Eo��iY���&o3G�̉�϶{�`A�f|�}̣��]U�*J�kη��/W���S���??�#²�{�z�6h{^S��}��gN+���<嘩�	c
�`9B͎̺"��I��S&_�ٹW�7L�|���o���ø��H��3#�3q��lg���f�N�h�WQ9���=��Ȝ�cz.M�y�X�aQf�N�g�]<oM���4u���O
u}HQȶ���)@��a;���	����Y��l�|��_s���.1�Xu@%�5ׅ*����KW~�w�h{E���X���Gr���5wK�b���V�S�V��D1LT�y��1�pvVgI�T�28�v�_t�!�J�,dʱJ	|7��#����:ZpaU#�0p��my(�5e�#S>X�K&���t���\=��7�ЛX�����0��[]w�5��sL�
 ��@T������*�m� ��f㬳���rZ�h�S71t�7���Yz�膜�.M�u{��C]hEl*Jw{�s)�;��s}�Z �{>�a.��tK�ݶzS�z�au�Ob@��%�tF|$���x^�\7s3O&ؓ��n�M��.u�N
U����n�\F_� �o��}��Va��.∶��.��p؎�6��wNR�{����=_�r����Pb�*j�sq�t�����gIX嶽�}�}z���Y�����hYG��Xcr�:u*gxe��CQ*�=�� ƒ6Ҥfc[OH[�zyǱ��G��޺�����Ryn4��I�g��U�D�l�r>�9�/����2GD�wF����뻭���n��N4�]Y�y�[I�CS�jX3��q�Qf��9���K��m�Xպ��n�M�����!&��%�ez#�]�J5zA��ou�gWEpW���?�KǠ=mYF{�f�0�y[_��rg�B��x8���Y͔:�C�f��#��]�E_���gX��1/ht�Y��]Q�� �/DV�7�����#�Y!��J�wK�p���{U���s�\V�u�xwv��]��z�J�e�]���AD���cr����+�j�2����v�j��|*�|;H�m��������aN��`�^�B ��B���M��	���H[5@�DU��ɴo�q��=�-�YO����eV�Je&7l�Ӣw5�|z�3\R�B�0����B�-�պ�5��o�U:%�l�F��<�q�#��-.�P�� ��e�R�I��z,��W;���o�+�h�]�P3�^A����(I���c���ej����[W�.'��b��5��I܋µ���=�t���>o/�L�����k���Iϋ�Nw�4p�`_g1�>�|�\FM�nf@��& ��خ�˭]��2��Lk�}fWr��]7��ف7�mv2 5"��Ӎ���6Oj�ӡ�Tz1��g.+"�G�WEO7�N�D]�x��H���������{g��h�{i'L�A���T���r�N���p]���t�Y|e�/��1^z)�=ܙ��6��'���8�lv��K>���w��S�YsίƑ��L��Yw��,%vi���<��gi+Ph�yv�8��ހ��r2 E1ϴM�Cp�guc�%7Hu�q�{';N����\�O�N��"�k8�m�����0eȇ���f�fy�D5ng�o����7�ͩ�ΐdwnS��f��<ɪ�Qtx;�H q�Xf���V`�kw�x�G�2�r�e�M�@97���<����݂���x�w�4�K�U���2�d����h��fEUr��H��Y��Q
�9��4YU$��H�"i��ʍD꘩�4���8Qt�1fCT�#���Eˑ9�˺�j\�3�J�$�lDupK�g(�U�B䒠��9QȈ�s�\9UZ�gK�k�y�(��
���Ü=F�DE:�3�������҈�K<�V"IU�.D����ʂ�UQ�4(��9Uf�Y��G9(Y,�\�VeX�����G*�eR��ʥhN��E9.�Z(�aN�T�XUkwe{�S�N�!��
9*E�̊ԣ��J.U DD�Wwq�WVS�8\V��W)Vy�UQETT&\�G$#w��N���N'TMG<�D�9DDAW"�@R?&��d\�P�����S�v��L�k{��\���㧊���;�Kn� snw5�L<y�dW-���X4]o���� �������N�t量�_݊���p�{��:`�P�Qc+ަ���}<�:��� ��*j�	b(*C��kD�oP�>��Y� H��]l����6��4��Or�O�b�lKy�?�4��a�� <����q5>��B$�Y�!H�>�eosޯ��Ys�r&��ͯ�S���#����f���Gp;��/*輖v�mf>�ݓЀ3��!�!���y����^��x/���J�h_w����Y۪�쐢�
�K�.��rp�H"���ܣ!)´�+�3�Oz��|�d�?7S�5Tv�%l�ʁ��]�(x�Ia{%�To�T��
��5#��uY�|�C�j���C-�B��)��wVi}��78��%G�"FD�?�E'�Dv�	Wz�Y�GG�ԗ6��-Nz�KQ*�͘��t��5rce}��q("��f��i��--�*�՞!]0�+N*�����V5�­yR�W��b)k�c!5W&� 0�`az^b���B��	/6������:�.O<{�bĴ,�E�8����$ݙf��L|ڸܺ�����\ �֥iZ�ޠe�A��W�F;�G�ظ���,�/�@d��	eY�b\W�^D�00Ly�f��+yPt�i�ۊv�HhT��W�v�t���}�U|�i�a�α��j��|vk`��A���N�}XGcs3���&T�}��_i��]ͼa���^��%"�p�J�k�pTmxua�ma�Z5P�@ pw�{7���6p
p��)=�/g{�uX�`^�Y�St�gD&�T�1`��3����� ���U�'w9M�c��5l�g��*�:7K�!�E�U����B���֬��O�AuB���<,�8��Xɕ�;����,�Ѡ,U���I���RgUOه~��f�ZX����W�0����n�K��=yX�J�
��p�h� k�ܑ�,�nuܱ�V�=�u���FRc]vx�~�2�_d�8}_#4�+��KP䴈
kCט�=.j��!��a��p�M(7����~�X��w�xHO�qIjL����_]�!��((�衲���Oz#��7�|3���5��Z�Á�Ʀ���|����r�I��&M|yw���?]do<r�~.2��%�B�!���Ҵ������R��\�y,}�ʠ��4a}D�|�_#SIOz,@�%aܞ�F��j}�Ui�{��{�á�߷6me��F�&��d��aG�;=W�Q+�ުߗL;������b�nfs��k5rer��:=۶��띷�R�%�����C��7i�S�9�c�;��
u|��K�����|*⨊��E���=�UUU��-9����\��׫G�C���g<X�Bu�M�zLV���D�ԅ@}]�w����ntC��)m�S�ܪ�IΉíǌ��R�C��%a�zNL�*���Q^�z}3�J�l�pϳ���y�_Z�/�5��ϡ��o;+�_<c��@������/Z�p�=�	�̶�^��~U@�qg��ڰ<���:��r������㰍���J���9�!j!l��4#�eغ�VI�P��8����]��_���4���S5{ݒ�R�/��7e�ws�+��T��D��:���UY��o)_m
�
��G�zn�9���aI���C��>��T�{n
����&יVl�[�8�Ͻ�XHW$�w�=b�2��>Bs��yB��|�8��bԬ���h{�D������������(7ػ��0T�Ƽ����>߷�9J�3=�EW��4y��>�H�J�&�}���vV��c�/G=��}ǉ�^�h�D4c�2��R�;(�-��kbz��c����5����B��[w
l�Zì
�n���RS�)���y��$�]W'J6��Y�I�K�^�Y�t�R�MA��B5��s`M��ݍa�ò�n�9 ن���w����҆�����}�/;;ғ�#�{���=��O]w���~��fsb��}�|>Lv�1�ئF��8�me/�I!IqwA-޷䫜A���Vy@r�ۧ�����U5:�C�����Wx�] _�P:Z�׎}ٍC���-�c�����#X�6�}~�-�yBb�q���d_X��_r�.�* ���@}���P8��9aӞ����'[��.g-b?�9Ưb]4/�:��Cꚸg�����hS�~�}����0b~�o����x������^.`�W�r��g��J���l�ۙ#�&���}��f׾� CK���(�J�)�H�M�_�r�Q/��|<�X^�a��Vy]�Em�V_���0ua
��%ܰu��	C��\�/iN(5rCn>�HU=����\��W�q�s�! �B�o	��y��'A�44��w����E^:i��SH�Pnօ;gu��ժt�P��E��jP��s)�]��1|�]���v`���������S���U���m>�3>g���������BiX��~��tU���_���=��5@���I3$��2v6S�%
'���]�ag�No��oz��%�\��!^ա�-h�n�z7��{�1sŬ�9]��qN����E��>������%v��m�Që	 w��x�oU����']�et��ǃ�\��������ַ`�z�,�2�2ʇ���7�>5j�;�F9f*r���O*c�HT
�����z�m=W��(;l{���ս����ҽ��RfZ�_��o���k���e�}H�*�0�:C�/�x9z`����z�As�\EeW���J:}1���(β��b���U�gI�����B���?C0��z�`}�p�0^�旙�uE�=�>:�Kl.�7*x���o��)�����X.�3�|c1B�����B��T�i�<*u;�#��i���x���N���υpՇ�ξ�L���]�2���Y�X}릳�@���qQ<7޵��V��g]���9��D�5T�ݭ�#arf�	Ƅ>�K&n3� ��=��ʞh��0�zk�Kv�,A��5�.�W����[i��`������.ϡ�,ǯ �q쑙��t��v�AO3òhZ�y3��,�z�F ��"���y�xw��y�Qw,�B�{ �t�fZX��^TOއ�`���'�*⦑Dp'�w�-�|p�8� ��7��rel=l/e(�n�� T�{8�����p�)�2l[^>�sqvSخ�C�W�vT֑�PoR�N�]_���Y�wkd�_<�s�B��ٱ�����v��e�E-���RuNz���*oZ�97&1!�35^=���x�n>��������������#�r���0EBn��fG�L�jOɍD${ܘ��׆�a�~zkڠ��.z��bݜ�j�o�d,�Tx��Hz$�y�J����*#�A*�X]���^�<�y��+=�z
%ӝf*�m0��"��}a�q)�*���	��E}ɓ�e�~~�	h�=�W!L\>9�����{A�����.q�R�(I����]��|��H�\�h^��4g;'�$}~�ao�>��Xo�ok`ּ�#Z9��c}XG7.�v�d�W�!���ߠ�N?/��40��m��=�e�j
�@�\6��ڬ;�F�
���S{~S�|Ͻ���.����5�+�=+_	��-��L�f�L&�Ѩ<�b�-����A�Ϸ���r��ܞ�QL^�5`8o�!�]+�#N3��X�ٽ1�Y�kL�QU�0P�)�>��^mm'����}�Y��N��cw�22�����;�Kn��kC�ƴ�	�A��\��ƒ�
[�Ž'��}�w�[��5��J�S��s�l�?
����ḭ�y	[h��^�J���#���ȧ��+����݄��׫&P��cˮ݂�ц�J�@{cSx5��|.��MU�Y�����.Ӥ|1SZ����o)W�>�NMme�����fe���v��R�hbZ�.��R'�pk��և������ҧKo'�[BٲO��/���U�_�jP1_�^`~�������`���.]铧`��z���g����ɯW	:S'�>��hC�PQ_�Cf�s������EE����������4s��[�c�	[O
¹_L$�o�z�*�v�?dJ�U{o���\�����g�^�����1���O����w�ԁ���������e�Yy��u<]=�~�;rTn��v����QSE���j4�m`��4��{1�Y2(�^�Rs�|_��9����&C���	q_0~!}|�K�����h��)�gk��}����>��E$��l�Tu�\S�=Ն��bzګ�����f��y��ϧ����7�{+t,��r�X�z���0T6Z49����f;��ޱ^��5I�OܘKM�_�=�%?B<|�]z�{[x�2���ByU�f���/l@�UKًb�G2�÷���DRru=egN��vd�A�C1��}�|l��ụB�`��Q�i��_ޣE���}�k����<o#s��wŘ��]�m�*���5��}�=����n��ڐ��y�F�oI��6`Ep+X3k�����j�כ;� `9�s���_p=���Um�~����|SY��^�#�c6����N<�C�;P��P���؆eb��,w��a��x6��}}����m`���P�G3��z/9��w��sk&,J�Oݡ���՛G�r4�q{+�;�k3î�J]�G�A��'t�+��)���XG��==G��cY�l����y@������;���,I�o_ۿ8��/{��v_��{���P����\'hҁZ�6�N��y��BM��	�fw[w�����sX���ۋ�['i?�<��R��ԥɼ�(��v�e�dȮ��7�z����=�9��`����	�bS�SX�YV�};�w{�[��}��2Ĺ����}��y8��t��l�}�=U�l3��M�t�>������Q�"H+d��'��Ϋ�vE����i��p�x/bou{�����)�FV���,����_Ox5����lE�3���ILPX#�z��`�-��)��'�X�g��R$3\��-G3���0_	r��;z���Li2I���Nt�����K&�C�0l!�Jo�Ѿ{�+�M.�j��7M������Cw���r��a+mP��Vf�Fr�:`�����ŏ�| kyΫ��:�����r�P��)�L�'K�n�q�y�:.�=��Z�἟��N�T�'��}
u���V�P������%ۉo-K1������0+��]�֬6�V�l��G���q홝T����y���J3�k�N�=~�>�����ǜ��N@��G��Dy����JLJ�f<�k�۪u��ݨ��Q:��=����y��2���w>�nJV�S�ޓ��,���dZ]�X}6������^OA��f�.�C��yZ�y�.7|�"̿�_L}���5�������nr�N��
=�<1��}��J�u���b4q��t�w����dÕ�eDs���%C�V��cVy�n�Y� �&xW��b��z�sz��S3`O(����7(�N[V���gz����뷀�B�dΑ�ϥ��
���g��g����Ӳ�}��j|�����öƁ8�3~���up�NՔ�k�;_�!��q�~��N2ΧxN�p.:����#׉oS*}/�%K�goe̎�8��hU�K�pl}��oORv�*$�E���A�a�oz�n��Nq������}UU_|�r��w�ߪTΕ>5ꢫ��	��~�A6În{���"�yF��ft�=&��a��m6��Թsj�9�ǫ��V�/�u� ,)�1�s��Qɶl���I�[�ζ��;����~*��U���.�+j��Ҽ�8ͨ��T9FQ
w���AK�Y�f��/t,RO=j��LT�#��/����62��*�W)��H-�8�
�z➻�˫W�"nǧ-����a�=�F���u�r��
� ��F�l^ە�{]gv�}�$�g9֭�N/9D=���~�~�+��Ƭ�~���ܝ�a��3�Ե�MI�N�MǞc+g�Gp��Ng���)-��B�9P��h��$?4�u5����P�ȍ���۹�¶^˄�.���UDyٺ��9����9�ovz}�JF�������.[OV��B�{��S��m\���x�`�:iޓ�k/��q���W���m��=$U�N��~ɓI��a e��j���7V�r\^�V�Ey�����0��A,�O-�7'�f+V�>��M����B�{��.�.p�j���5 �jfs�;.���%{��x����TY}"I��#����:��:M�U*&�a騪����Qp��+x]d��,h��ԛJ�0���e<NՅSf�ti��Zp$�Z�(N�&%I��4o�#�>`V.�WX�L�reoX�g	��IrG(g|����2��n鹾�@�/1�Aޡ"5v�4}�o=�<�ܝ��k��:�;���v�����]Vp��k3:��q�NG��\]�}�W��(eH�'[}�g�a��[��QWO��T����I�����tL7�#X���:�o3�D�Ya��Ԇ+Ŏ�����B��:F,���x�Z��{�.�&#��L
��$�I� �y�e�QX\�q,��,����դ*�u�5��5��:m ���I�/k�B��y�#�Pӳ��WI僑ۣ��<�q�S/�j���bV�_'�n,\�RtqpKU�|�-�e�\e�%�2����H?�J���ׂ�uu�<�DP4m��:`}g�W��a3/1i�����i�K��x��U�S��.h���Hżf�慓������	��̺6����4���X��񙏩�{�@���/��s�B$���v�»����βi7�gB	��\��%)wO�)n��e�9�S�Q���-�yvq�;2(1���LˌTo�sd����[�bD���aWK�n���F?%�y��OZ}F',���c}�i\��cZ�d�v��vQQE�*[�k���b���2�Ѧfo�/3Ϗ�ٚ�î ˻��Dbf��I�V�z/9-�/��K�����j��:_o��5 �v�,Yݶ���I\�[3ܶq���T�zN�	 Μ�n�]_�s��3X[.V��e.��Z��n�Y�7;z��vWJ+5T4Ge�V��У��o]��y���K�� �zrS)�$�Gsv��ux�p�c-%RƸ���V�݉��.��3����\��}���a2�闟��3e��:��뒩��$�un�*\T{<�v�/22�]\��k\Pv�>]�̻�A�6������CLc���ԑ�kYz%�r^W�\�5�t���d���'.^!���g�Q���KV�W9�������5�W;��]HvM�����j�A0(�#�I��2�;�Z�<Iu��m88f�j�i�뗀U�8�d��|E� �G�V��o��fЎ��քS���v���s;h��-����C�FQ����^ҙ��8����M�����u�Vk5�R9�up<ϛߒ��yu.�Xޮ�m��0�6���L3S�S������)�tk;N��:&�\K�ʃ�(�)*�O	9"ww#�r���PJ���E�Y��IN�g8�!�*�"�U�9�&��+������+�'
d�&)s��U�$=v�eHr2S�&�r;(T�s<�XN�g��T�<�Z���9PEV��.\�ADQ��\(���:EK��I�8WXTETK����X'I+�W�:9���H�Ә���ݔ.�tۊZ��*#�!	���OB�rS���G
L�I;�W!R祚��grr����Zt�u��GU@r��K�%s��Yt�*9Q�#�L՘l* �R�U��G�̓�<�=kQtNQ�Tw4�0�ȯ"�r���U���j.B\����j�Zʊ�4��ᑷu�8�mY�C��aqK�+��i]#���պ/��X��J��qݙ9���Cm��ś2�LHۍ-�#|��������������E�z���e�5�.�9����(y�%NL{Q��n�30���
��u�K^��I�/(���S�-��������6�K��/3�y{9?V��R�՟T]<Oz��oz������J�w��J��]��%K "g���Ky���RX�΅�o����K鳜=����oxc��8���;As���Q{m�޺|vD|��]>�����:Wff;����':�9���Q{�1˼����-j��-�?o�:���]�x����X|ʅ͇ì��p����ld縭��wӽ�a����"�z[<��2�r�wL羫C��R���N��>���2C�آ���HQB�0����9��(S��J��չ���B��[���	�[c)�2��Pm�����Aj��g�.���j��0��̀�T/hʄ�W��<a7q�_>���
�����ϯ�n�l�ۍ����V_�\*�؟� ���
��ቇp��m��s���4&J@�Yf�'6dȟ<J˖`���{l�=x�+o�{<�jI�R�y<����x[��ũ��[&��3������ot�6��화�����gJ	�϶�w99�o��+�q�z�Z|��
�oc�,W��prigC�S�k�7��.ْ�{<��u;��Mt��h����V�l�]l�y��q��"[X��c1��)�n{�,������,��Ǒ��8"O@�����1e�6\ʳ�~��jl�f{=�8�[�9��?J𾎭c��k��g\%/׉ǚ�{Gj��8�v�ZV���NWt�x�G�g=�����+G����{�Gg��yzzb^��f�M�D�O֬��YMX����_A���u6��3ïᒕ}� ��sp�sp�~�s@ׁ�8oB'j������A�2�;�ys�+��o�1����^��M�u�Y-6�%����G�_n�ά�^�d����m���9Ʒ6�e�������U��7<d�|㝂[��^�n.�d�2�P�AV�g�����0���f�^f�����g��w��3����ջ���n.Z���U8����T����ɑ�竪�1���!�ЇA�=��Jb8�6eؽ$��I�����x�b�S����2kx�g�j��f�K�����!:2�������>��^�v�瘶廫�����~��&ێn+��c�Wx���Oy+� �����v���b�!����%ͫ��G���uŽ�Qb�k5�no�q�IeX���;�zF�x�/��uwҧt9;��i�9/�{�nϫ;1l�\t��C��4V���Nr�w��(���=��CO=��Qd�v�7��.*h�	��S�Mt���٫�WP��?Ki�o�^��$�0�f��3��+���I����Xn���k��Vj��lN�[�j�nI����ѡ��|q�L�������.)F#Ý��ؤzi>{O����x�jÐ-��w��G��If�Z>��h��١�]n��[+j��Y<�oM��ɂ:��y�ɸ�^���f��`jJ(��q�?n�f#o`��G�/'����D�tUm�q����W ���k
�;���Nܺ�.��q�e��;2M6h�j�gZ�6�������p�-����r�J�����VԾ�Vu�wJqm��֡%��y��,�gM��Q�żǼ˃;�'%|X�����ڑ�S�cw3�sK������5��*��T
��}�'y��_|]��l�@���{&��3�v�R�%zR�L
�e�ld:Ƕ�ݸ��۳��3w���^X�{&�:u���:��!~��v|��C�[���wu�^�A�U�`J���x�+�Wn\��a(�;�kyp�{:׶k���ά�N/Q�X����1�Y?�O�Mz�u�����{&�=��M�㛛����`��䀱�����]��������+��!��Ӕ��ת�`��W�@����!v�l�q��*�7~z �l��<���΂5�;��p�s��kn��s�&�8=�2C�����}�a��zlq�����ʸ��se�C)nn?�����Y�|�_9fa�9HƉ��b��Mv���GZ�r'�N�={��ǧ-����a�=�+�L�0�}�])�5B>��}5��u^F{bu��r U���=R�_];�5ۦ��b��~�����󛸔��D�I^��dЎ>�����C�W���|'ES��=��׮H9��D�p�ɐ����(�m"�F�Z��<��d�S,�3�uvz-��I\�᯻?������NP�{�)�9����VN�ϻ��9��R�ۆa�l��)t��$(�{��U͞�F}0�6�e)��W�m�������8�X�Y�.R�Fi�F���tX��˾�F8���Fny-�?E��͝}�(�BWn%��N?�O�a���r�VUG��lW;>������4k��r�O3|�@ �woB;��WMjU8��.�o��]+���[*�O/dsj9z=����g��H|%�v/w���BڝiS��������ӑo|�,=�>ʛ����=��'�Ŭܭl[��N�z![o=l*!�ݭ���#��x�햻i<��ضR�a�;\1��w����>�n.�M࡝~�ԓ׼O����Y ���@�t�x��(�U"����X�vs`���'��vY�t�5��C�r�����N��漛�<�>&��\Y��3Y廏�Ϊ�pm2͛��2�K}t f�˸�㒎��ͫcUp���9�BR�g�e�R�R�z�K4T{p>0P}i��>���O��W�;̔�����j ՃyS�J���[Y�\R�c�.T�uʹ̸��x�8cםȒ&��j�.��ܹ�����.��yIV��W����N1�A6���M7�����P�rxoF�<�w�c
@j������U���뗹my���ڶ�X�آ���v=6V���7=m�q�ՙf���\9i1~x��8��T9f��k"��0so�[+�^p�pO�Qe&�5>Z��*�{FRM+�^��e�2y{k����{<Ve{���ǝ�V�3|�.���y���];�>�'�����E��; 3F�����gE���|�*���I�nw���?g��^��E��{J�9�.�l�k�ڳ����D��_/:gz���%(z�b�˒v��ǃ���8"���[a�]��ucdZ�s[m��M���n���J���;ᙍ��c�����N<�=����˳lk>�y���<����=Gu��v�ԧ����(_���u=���;��ԜZ�t�QjI�Yk%x�����/�A�v'W�N����N{Z�^��4?,��^6��o�{9�z��*���2�#ԓ/7&t���wuF���^�:�oX#+{(���]<���l7{Ua���հ٣��Og\��q�u/���������˕���TD,�����V��<:�JU� ����~���/��@��OIB����h�7��u���xv�oNs�c^f{2m9^0*C��~�i�;��{~��HI� �?��X����E����	un���o�nx��9Ҝ�+����-�� ���Ә��E��x��������n��I�'��'�8��
�g����k��x�S�5(:��������jn��������5���fս8*'�%�ǲ�{N�wJ��6f���'�zF�x�)��3k��x/G�0�s��`�z��D�	���r���S����	K yk̪�9juN93��Y���{Z�;r��m��M�9g>D-��|<�jNݼ�tto^hJ��}y�M?{ڶ����'��`vg�����gr���Zmv���+W*噴�$A/Z�`,����Ft<jpˑ��y2��:��0>�7(�Z�d��lp��K�+�Eӵx̫*�Kӗt�{���2�N��g=�Vp�ؕH�kF�$2���]ßG�rc��㋗(���2g,�р߾���5��z��НW�S�o;�����i�
賈]�q?y����̬�w�μ.�aұ6��QT�y�����yU����p������>��(os��7Tn��˒��|ե�Y�md���/7Ϋݞew�ä�����Q�_�vC<�n�$\1P��fF���)�;g�^���V/G{�'Yo}T�uA��ײo���cZ7Z�er;���	��r�߆�D,�W�7/^�&���=�X������ߧ��j��-��*É_h�՞�����9�Y���Pl�����Hr[�����gŐ�z�$��n<&�ءoI��Ӏ�ɭ^|#)���ɜ$s�ts�9.����t}�#5i^G�iS�bud��
�V�+۵��__`2OM1���v�߱�^�ǬQ�pk=_

y���s�+i�疥�sj'2>�r��R��l�u'	���d�[r�;e���+�G����^֓���5�ʴ/�����m�ߛ���v�sf�՛�W< ò��N��hnm�J��;9*>V���V�6���Gip�#}:»��z)X�ͮV�3�A����_�GwֿG�Z���V�� �P�����H�1����%1'�$��8n����������*���9�+g�>N3j�QQ��
w��,��c2VPN]�N��`z.�=��m�����6�>���U�dT���K�[��k�&yA���l�JZ���X���֭����(uQCmu�z��M��Y�}�{L��)��k���z;����:�n�2�Yw��;ޤ���x gua�}]4^R���f��摬S�S�:yx�{�f�㋘�6���0q(r��0�cf#��U�7<�����nI��~0��y��0�x���Kޯ�-jr�|A}r����p�^K�/z������ߔ�'lk��U�����K�n1�{G�Y���אKhw�A�O�\n�.�x�<;��a�m^Ih�}Y���vOz����~�kf�x|Nx����n�ӎ!�D{��,9o;�t��6�<���Cf2���H�d߮��=�d7��Y��2��1˰Z��E�a�Ok��I�9�yns���G��X�s�R��l�D���.-�����j�5mh����cщ.}S�i�:�:/��}��mq
ŶHK����Ϧ� �{�'qk7+[9-�����k������/n0x>��{��t��̵TƷ̽r��=�B��d�33V�������q��d|���^���8�~U��Z�uJ3~� �dފ��b̶�ˍ��&5c�~P��]�����#��=޹��C����c�9����eTs�8��������[b�g���	�[���r�ۥ9a��$�j��,��=[x�ç�P��5�y}����2�r�HY�]o�ii��@���g��#[xkgn}*7l�;M������Ke��:�s��Fw��)s�Z�x<�����o>�K����x�}&6���w�~���Q�[-�E���7)=�u϶��Ng|Ѝ��H���{'�f�%����_�a�q��x+�M.gApm�{꼾�Py�%���Ԣ���sa���9vQ͛
�br�c(��ov�lE Y�*������;}��>�ܐ�5����k����Dcm�N���P^��[�U��{K�R\�C�L�L�vh��-hluy�y'e�r��<���~g�e��%�{Ӌw1H��}��(�a��n���Ǖn��륓h��}n�;v����V��ٯt�5S[Ǖ#z�Y�Z��L.}�w:n�b��k�X��v��L=�#�b����ږ5�0�s��c~нY��\���m	-�I�ڷ�rjvr[;�.���3�odRsfmj�/V:F7b͹0�W\����{��<����jd�}�c�[ԥ5{5i������͔��w��3-)6�u�f5pDE����6Q�E�-���B�r��Bx\����ec9ےT�u�"���]x
����4\�� �3���6
4�,����f}�^W��Z3��3�ȝ��Y�#Q��^�5v�U#C�x�$A�i�B��m���F�.n��Pzٸ�|�v�;�T�7
�� A�a�vb=1@39u����8��NP�eX��7D�*�<��Rg�a"�i٫V�;�M��1�{�<J�^U��зs'dt~��a�������@qj� ��)<���:�lȪ�ْ9�6	{}���sT����8!R�ģ�`�,Α�K��L=����[��]˼��ّ�=W�o��[��G{�b] ��̓�eN���n�i��v��.mKu�о�˜��H�J��)
����٭ul:]���J-n� �}�R)1	}�^�y��1=F���d����@U�!��ނK�~���u�ə��u=�3r������A�9��hl3u���h-��/��Zk��%g�FҾ���,�e�?no�C�y��3�pfH_q[�)`SI�"��0�j�۴>���J�ۺw�V���a�A3nT�2���gb���з��[r>�нw�+6Exm��X�W*F���~��ˡՊ���/n7�J��ۥ��(Q��۷A+��8���ֳ��8jg^YT$͗'m�չų�&nu$ �w��6��ݨ��Y��u�#z��J[��|��q�)�	����]��c|8l�T���R��!�\�[�����Z�w-�*�ԅ�IS�q�Floԏ#^#ގ�(ȕ˞�EW�r�@g���;�>�M^����;BI<d����ܙ�\��z�˚\�=x�}7}4tz���AC�Q�sT�9�7+ 1c�5��r�.��{^�<@������>�
]yS:�n�����Y0��f��#w�ࢢ��1��cJ7gJ<�Qm�g론*�^�Wn�� ��9��:��bP@f�+���cP<�F�ˮթ�H�F
����n�͖8p�Y'T��X�I�8�DY����u��nU�h���j�k/������3��F�Y�P�A�S���n�h�(�ޜ� �VEG"��/��;�����VZ"i��H#T�'P(s�Nw]�P�R㻅8t�*����P$�99,�;H��G��H�ݪ�T�Q�H�(�w9HwQ%�B.�.�z9G��L<��t�+��Y�S*8A�r��K�簈���xQNgV!�L"�F�D�yd���!�L'%M*�QR�$8G�PU˳E��G�r�\��u���T/2�݅TEE���S"9\�a�u�r5M=ZI�*��s�!y:���Q
,�]�/*B��ȉ�RwS����e$Y[UG�(���稫I�Y,�6�Ŭ��'E�h��Y	z����L��f�T�p�+"춥TwP�D;��N�mK�2��­g].r�x��NDY�8��l��+��Z �痬��9dvTV뗄br�9E�D�.^z`EIQu0��YE�><?>=?=�gl��F95��P���|�=L��3G���
G��:o�����s`�0[© $�J� �Ǻ�%s͜g��W�sٹ/�A��?���<�ڰ1�U� م���s;G;l���<���I{��S%�5�k ���}�{����/������ʯ;7�5���q�˷��nA�s�h��ٝZ߫9-�'��T�{K����<��S�*��6�֌�|7J�1�s+��b�[�>VO��iv�=��Ѩ��W�Ɗ���������;T'����ƿ4�|��m�A��2�tj�:�g�X�J��a�d��δ{��>]� �G����M���W�q�=��@�:^\����sF1��$=���mh�f<+���d;O��7팲u�Bz���O�O���ݱ�[�R��Ƥd��p|��o�͊xG�އ��w�}w��=���^v"F��'�o����Ԣ���f8�Nw���~�A6�sq\~�4�Z�zN��24��f]j��eAD��ݿ�U��}^��5�~蟩IZ��N���k�Zu�f��"�z�42n/+�x����Mh	�k�B�ݸ��k�V�䜺'u�+��l*�`�Z��=Yɲ)�m�\�s�)[����ٛӵ��AC�ӡ�[s����țtN6v�5҈/ Ze�&�C�`o2�u�d�qv�5��%x�>%���q�Ew����G����oHޏ~�{:�T�l�W��y+t�c����d�=��Ӓ��'�w�W��F����/��s;��k�E�9Y��jrb���~�����Bo"��3�"s
GT4	�KU�����/A��g�}��o��+�I�g�z�௃�'�C�5݌(�<�����[�+�SS���m��Xu��T�zqx+e�����˔C���l���z�{WȊ�^��I���x���=�����r��*��uvM��씖�2=�r�\����K�o�9�*s�~/O�W�<އ�-J�<5-h�v\ i�Tq��Q�f��C&�ɪ��)�;g�Ϧ��	�wd-��yD���Ȭ�.�����d��֖��˗�qQ��Žo쳭N̓;�����7�Z(O>��!���;}�{r�w�c2�n ���6u��6o3�������o�o�Ᏼ���u���wBd��痫tC�C�*l�?a�	=Z�;|v���+�w�u�};���ݜ+h؍�35�XZ���Z��Nn9Q�ۼ\����]>}z��3�l�K�)�4��1 [��%g'�Ý�H~��)w�����oz�cf���.R� ��؛�s�����D����:Z���\�,yұ���X�m=s��g��`7ʫ���N=��_��<��W�ݮ�:��I3��'�ucC۽2O\�ϣy��pCjl縯xQ�	�	��V�&T�}��Q罣v��r"���.sx�&���7=��'[��g����$�$�1�}�T�Ư/_�k�.F��K�/u�{��'�m��(�ЈS��C�D-Ҟ�{�Ѭ�{3��~};՞�%-+g<�|�Wɱ�Y@)����/ ����Rb�	�U�N��n���Z�e�w�
ø��6�ʭ�#�rU����\��g?f�a���7S��:���$�y���)�����r��U�����lpWu�_t;E=�0��3�e'�k���{@�y�O���W,��+(7�uB��FiA�ǲ7I��)f>��-�Yڳ�T[?`o�z�{<���kp)��}���8�w$Y����,�U��Qj��̒q����WՇ�J}���ӻ����]�	��{�4�N��)�\][�i>�v�v�m�ݷ�����5�������"� ٟ�cf#���8��>αS�^{5�V�!��zZK+��&�uj�i��bp�<����<��G�ص�3d�S���a8�����>�?:�^�������x�T��n<��9u~tiy͝V}��c!���^�ݶ����ҵ��)_l����;'�k�j�=�m��ݸhk\dے �g���W��oMU�ۇ�^uzR�s�J�Ô���w�/F����1�n/]�:�O+��ղՍ�ώ�H)�q��;��ݹ�q�� {�j����ݶq�N���t�����Fu�J��͚ۯk�BD�&��v�1����7>W�f�P�N��0��U�Inu��*�7|��tS�p<��%˫����c��nN~4��=C��M��.;�
Z��"g�+g=��YLm_zq�v���c/o�ך���3m�~r��[�x�:r�x���|����.�����!\�޿b�]&���.��c��I�,&�_S�RY���cwe	o��'f�t���>�)�s����=���{#�nR��8�HH���TL�I��{"���_����d���k��Z���}V��ʛ%${�����,�W=�����y��ۂTo�{f���U�
�hx�@��A��{��S3���>�`Ojkg{r�����RzE:�<����Gy�Kw���4So"�31��
U���N�N��<�Ӻ�cKkss�֤�.�O����f��x:iW3�S�{+�����[�Ⓒu����o�'OLqڱ�¯� ـ���Z49���������W$�q���1{�<�sJ|���?N����W�ח�=�-��.�塽��ȗ=;0z���tO�uiMȐ��:O�����g��R�������� ���OxҊ:�ٺ�xfWŹ���m���{��cL"���Q玺Sr��Mp7�:^��ܵ{a�fst�c���c%@�3<��~����-�o�
I	x�����f���3��)��SW��~c���y�mJ��Q k/�!���0C�$
	�%aa�Y}�c8��H�ᏴMw�"nn�bp�6�Jx>i곖��GXA���ˎ1Ѷ��C6wR�̔>���=�H���n����v�S\�Kb�gB��)��\O���U�e���I�u�=����7�B���8o��M���/�pL�7�d�|�_��-�}z2\���Ք�/]һ(�n�
^r�
�V�4�oy��*2'�Θ糝N�W��1��!5Q>�.�nʨT�ik~����bk�z�x�@�Θ2�=/ڣF�wk����L {�wvt�,K�W)�s�N���Y��G��׆D���%
U ɧ�)�E����L"ޛz?x�7܍T��<����o#�5އ$ܩ��A�踪�w]P���ot�Hr����v��0_�}��$o>{d�3|w�t̢�K>�= n*�<~r���M���F��=9m��+N0;a�q0�CȊ�j���%��x��Wr���=ܟ��k��w������7
�N�6���^�[���}�o>��p���#X��J|���?N���ꆮ�=���Ɛ�x��w��>�MC=�{J�`ht⾑f2��v;�M���fo9#�{s�_ur��5��r
�O?��e�y^,-�g%X�M�Ԥ�c��uGK��u]#{�l���b;�� e�n��<�X���g.k-m�q�����ë����U{��m�@��sdhJ+�ս��Y
�Ð�����/f5��/��ߋ���cQv�yVn�^�Wp����W5�Cڮ�ݨH:��U���+�0����XbK/��=�A.E4iVjŶ��W^kF�X̢�`v%S���M���Ռ�z5�u˽x�~4�����*Sc!�=���׽n�V��7Ɯ�/uGeH�zb���}�ɋj�J���(�����t��*�z�^�^4�g�}7t3=n�e�7jͺъ������P�@�c�7��zf5���Kp��<۬�H��m�O���R��v�r��`V�-�{+�>�{שy�u�q4���R��9ҙ&�A�M��pW�`=\��	�g5�I����hC�~�	����W�f�ڂW��$1�A6�N>�M���P���\T��8�U�nyY��oBLz++[U���뗻p�=�Bq�Qm�e��tＮ��cB9i`_��S�t͝P�$'L��<F%��Z�N�׀S���P^����}�ξ�_�b��@�'I/�il�ʮT}��u�O����q�Wv�pY&�=�O�U�S]f�u�3sY)��c�6u^����R�d{�������ly,gMPx���	j��,څ��Z�����BleC�H�t*�#Bn��^�$w�a��s�Q:���=>�����^�a�
��s���amTN�a��MÍ�3Y�@-���WV>�����g:�L���aU����Qd��C4l�f
rѡ���A�^�Ȝ���/\,����6ЧI��s�ܒu��E�9�/.�b=x�t�j{{&X����]���1)��~���I�o�z�_��q�tǱ��*8+���k2����ў{��J�����-��^��g���S�z`S�VOD�Ȱ�\�_��ew^�3��w�t�XqP��\o�V=a4����%cx�W��������H�q{��imP�����2�`��1]��e>��k����1}W�:�K/�n��w����-����k|ΩRu|5u��~՘�RF�����dzl7տ]��ؘ�[�7p��2.�׃PFL�L_sٸ0�l�X�H�Cu�ݣ��w��v9F�1nM�
�]\�f��*!�},�	�V0GF�js���x�luwǻ�۸i��f�c���Y|7G�C%7z��09�Lq供���n/]�v�Js�[Qw���5|�*O�i��]�RM�5��&�=�z9�%���z�6{�;�TK���&v�,Y�u�p�f9s�dC�.��.�Nss��=�A6���q[b����n�%uc�%��OP_Op5o��RU��=�^ߚ�[�����^��s^l�Ř�g�Փ��pfP߶P@���kY�f�=���J��?z�n�7~Ĳ]߻�!`���}����3�������du7�_�����L'���8�q�'�g����qW����n�ғ~��'G���Vzm��̭����V�UϜӶ>���q��6a��gh��͜.�Һ�;��~�=	�I~�X;��}=1�j�7
��^�h��tv�گML�u��g=�V��rAG�+�U5V�S�������O*�j��5s�7;�ow#x�tE�Y[��֫�~���b�W�u��l���ѓ�YQ�1�$'��~�:�^���ޫU���5G���W9n����X���GXJ��[� }���w2t��U������X���Q2���9�.�M�b.�h��UY��K۞Kk';f��nm��M��Ƿ�q��:K�Z.7�!�gZ�˾~��T3#W�h�u�)|��w���ig�nT��\��x�͏'ke����u��8ק*Ëpw�,�KqK�1nM,^�նA�q���j�x��T/(�u��s�{�
�/����k�M�Y�������Ϥ-��~=�?{c~��!n��{�L@��a�̯V^��L��V�k�V�6*�����)��s9q:��<��efj�eM����A[\��N÷uo�ܜc�z	��%=��^;A�=O=����΃2�����>���k�!}��t9]��E�q��n�d�=�u����oj�}�{�F�I���L�3����!����r�л�k=���@�i�D��4]w͈l&����5��V��e&�ev��5�q��UUlCP��8�n�{�Ƒ��z-:����}�6C�q�oQ���G��M��7�T�egtl��b�2��ћ�v�N�f��Ñ:r�ڽ1$�:�ͣ!j�b�й��P��5��ךn����V�X��olk)(� �#tE,�5���Jd���)wo�V�{��ˏۅ��QC��R�g���S��\;��+�Vj��Y�K��E�!�2�)�s ��/ެ�y�{s .e�O5c��A\�˦'��
e�{��Ӎk1>�����(�F�>�ӘT��+���TsU�^�Em��x[��ˮ��KpV�l�Y�S�%�"�w]w�����0�=�~�U�r�R=lu$�ѧ�����E���]x/w��4p�GX���o�%�W��G=��ez��9���j��I����]��MS��b�E��]Rc���7�ڬA}T�TO-K�''�'Wtcu��k$TE�Hf����;��o\Z��R>U�f�W;�痈(} z�A8�phE�k�.���໦�*�;댤�9�Ɛ7�fL&�$���)mj'EY�q#�E���Q��>�ۤ��x�7/���tj)���l��r#��e���õ��c�����'4��zp��	���/M�)�,12)��j�4� ��{�����ՑzK�u|�|��V:��k�������6��ܞ�!ݗ��7_��>}��[E�B*��\�1�̣��o0�ʂ�%��-}e�Wm���eʂ��_{��������%/���j��V��ǫ=7]QN�gc ��Q��j���o���5�\y]f�yA�/2��>�F	Ocz����d���w�j�-�~�"�|�s�4cE�^�`�}�W����ٙZ��DH�O�q�̥s�.ˏj��]�� ����.�l���X|꾡���D`� ���ޮ裭�B���rI����ٹ��]ƭ^'{�+8��PL-X�e���d����r�� �s�m��8�k��Н����.�ʃ`���'��p��`�Iz��.�H�)R)C*�,t�9R�Z�`� {�{e����L�c�]V�k5^�=��glP��HY���WM6AEg^6't}�Z�Wb�{N��յ4᭼��B��5u$��6֌�&%�p��!�̳�s9��E�5�3���4��&��e���BK�M��� ����U�+;}g���1u�a�V9���>8�Qh�d��<=S�9Z;�d�A�e�;�Dw�-.{�Vp6�7Wfu�kQ�κ�3r�r�j�{��^��E�Z����j�ag<�K{T��N��o�Y�wC(�M���y��r>�ȼ��Q�/z�Z��i��|w6�Y��(T��k�3��|W%	�b�*U�����'"1*��[/6�F����µ�M��XfZ�Y�e���A���Q�
���=��H���)"*w�S�$�ប���NH��G'	ԏ8YU\�O0�L5Q�,��n댫�r�2�wJ9���ks��&)%z�V�@s�G/tI��p��[R����e��N�#f���^��y�PzʠU��DJ�qQ
̈́N��NE]"+��M�I�P��Ԝ�.�E�'a�aQ�U�K�!]CI6���P#Rs�xd���z��k���J�4B�M��H�EJ�H�TN�;��(�Rj�1FU�ݧ�I�bRCr��xm�:��Ap�%P6�,H�K$R�ԳTR�X��J/6�M��PYj,��jdn�;:��%�{r��֞B��W�(��C�$ӕI9Q�z���^��*�Y�y�eY��"���^��^Nyi�����d�gH�,�^x�;�/wj��D
p㈹&Iy�ib�q��h�l�$s
tDwn�2ˑt�VHu	t2�$��L��!2��)��8[����YAٙ�f��+�ֻs���%R���͗;i2Q+j����w�Ke��gD�b���i��5��w*t;M��/Vxg�W�����y�PpJD@<�Y�=W=�a�Y�|��ۼ=�~8��k�އ�p�4�L�'�6���l�Sc�;�z�*1�˫�~�}�:�����$�-��*�}8m���tK�x��������y�_��D��c�͛�9�ȝ[ڠ��u�<�;!�/%S�4-��{-�x�����b��b�?G<�����$л�MvWC���}F7���ϩ<�۳u�L�C1���46�u�U�x���R���ꞝ��Ƈg��˧L�⧸j����x���Q5��ة���(���9�����>N���K��q�`�ܖ�Yf��,wqV��V��=� ��k��|����#��5��ܹvz����C��12��T�O}6ϟ�	Ό��Ke��(J<�h��B��@�̠%�J����&�����M�Qksh��np7�r7��f�A���ı���֗Yh����Zl�}�/l��ެ#��M|Ni��t���wW-�(���Ol�M��LR(�y���}bD'_N�4S9����yގj��n��3���ū;7���q?}�{���Tg���kW��uϟi�(��l����:�g�������m�7�_��W2z�a9ح���'��/�X���2���A�O�Y�r�[A�c���-)Q�9W}���1�x��L��3q��2�B���f�ʞ�|���8��	�mD[c)�3�!{'2۵�Z�1�4��C��|����Y��������9��
���U�-��>�jf���uv\|�zR��٨�Z��7Q�NW�kV���].Zy���}Um�wEq������-���gr��W�c��\�`���YW$}��z5�m�����0�6a�>�o,s�i�?b�{:ǭ/�3R��w����m��0+�&���p���=;���Z>�z�Ƕ}�7�Zv�:���Fs45�
�o?=��cr��������> ����>�Ɩ��;պ�:�N*5�Y�@���e���OF����ŷ��sz�T`<��@h�7��]ыF�Bwj��Y�� ����P���:woD�]����E����v£�j����H��n���c&�sz1wf�e���+�|gC:V���_wf<ұ�9�z��n����-�������5=�~�������u���ᦵ�T��FQ�W�f3�#1�M�T	�2��(�z��[��f���Ow�%���!����?����8�uy�]YO
�=zO�tY�Sc���G����>ݺ����8=��.�˥�e�%tV�v�yݽ�_E��;!��s��	�<��p+����N�˥X�f��Q��L�*G����gR��ˌi��N{E��h�ܕfnkͽ��Ƕ�=�N�7t��U ����c�L��'=����S�(�:�i�lf^۫��-F�y%q��ۧ�P��?{��'�Q�o��k�����)�q�Ϡ�f�﻽��#z<`�u���%F��poP�}UY�s�S����;M���Ĩ�/;�ƛ�.�V+_M� Uz��n�o���鮃$��E���
���(<+���Mx?W�'�1�m�ݮ��l��v��3j�����6�2"����Ⳮu�31q�n�Z"�ec�e.�.��q�wve��4��k*h�$69rG�^�sx�v�]J}�m���gC��ʻu&Ov�����zE8�3й0h���)������e^Y~u��kKJ�	]�4��=�go�Ϣ�$�`�zqx(:iW3��)�+����K��9������#٧z<������7
� ٟU��W�ue��j�>��y:��Y/n܉��+�|�O��Wz�<�AWy�^ۣf��������F}N\ʽ�iM��%���>��^��g�u���S�4$���������˳o�ü��uJ�����q�20�x��$(l�d\;����[�1e���z����A]`x	B��̜m���4��rϠ=§�����7������U=\�Ӱ�������VSZ;�����6�0Ks������� �tGx�Λ{(eK�*`롻mr����� }!�����s�LT�exp�^z�#ي�ٶ~_X�X^�qw\�stȻ�`�9��5�]Q�]��btx)�o��}3�:�
�ؠ4kb���2ᔓ���z=��Fs��C��NA���Hᛥvi�Ű����B��.t�����Jf�J)9�\�+L쒱���)I*�t��ޮdv��;I�_; V�)�vbv�ݾ����'�x��%����c�Tٯp+�4v�]��M
H~������dL����]�I��2n� 㛃�N��|�b�������k^.�������m��U�"��&�E;�/N�3xd����4]��2�M�"{��e�Y�T�ۂ��7�P�J�g<�|�T&��2�[�ŏ`s�V�
�9�*N p���V�{�Nzr���ē��=�]n�)�Z�ْ�{�L?%��V$ګG?f��[��>�Xs�X�v�0,Z�{o�{�߂�sc�,Vø(wZ5����=���w��Vn,�\�cji��в�A=�#G֧�\�m�#��h����J?=�ꌛ�ڵǐRsB�^���OSیNW�}Q	�l��C����2DB�W�g�4Nx���ܩ���1���yn߈}��*�)^��3PC���\wپ�+�Ax!��e���/]�x���չ����ee� F�*�_N�9p��>�3x��K.*���.[�:���&�땴�*X��{�]��xV��NŒRRwJ�8g&n��"uq� ΛP��`˛#��޳�����8�ɍh�}�ww�����{f�V*^�Si��ʈ���������Sa:Ƿ��_k�1�2(�{S
�]2�z�.h�ö]:��bv�+�ΰ�	np�������]w���#�Ť���__�e��6�]�������x��z����嵐?t��@�G��v+����L��y�^/X�N���6d�w����4j��/{���'��I�sp+޿�������~��r���R��x���<��R��������<��^�p�V�+�IW��U�{�X�6����=����\��!?m��;�Of���k�!8ͫlc+d���j�ǛMF'��b���?��P=�M��?F{=�|�y����g�y9�{D�⃜5�aU1s'�-��7��Kmx�-m��x�]�x�`P��)ړ�in$:]�̗s\�pVr�݀�0/p:"�x�!i�uȚ�~ð �L��h��b��A��l���"���-�����*`;���t�� �ɘ�]!-ȵd}B�'�wn9F�yK�0���o4>J�}/LW7R1q���r�6��\��E�u� ������L5\�������U�>�����?���W����1˗B*C��ƒL;���K��@���:��Fn]��y����wL=���e�#�׎����9�/.�b5�P7ޗ�����Ϭ�Q�/_=�a�X����m.�;�����'U�*4G��S<�c�Q^�l��w�s:�wz�oN���m������?��Z���UYې��4����v�Ǽ3D3s]��)��A�WZ���k0o�c؇u���1��~q��]�=hM�c�Fk�_Pi�n\z�t�\�h�R������۸�sm{�[2�*��q8�>XTΜ�>�	�ca븳K|$_P��}�&�z_�g��c�n��n&�K�tyfU����8.Q�^���t������i���?Y�N���N�r��I�-FvV����{qI���P����~O��;��g�u�fo�u,�#�m4_E�]��ƅ7��f�a�2����QH�*v�STѪ��vzY���-VE�����F����[��q��8TvE�ܛ2pi���)rW��8��3�|ԩ������:{��6c�J��Z߮����ͼS7'[.L� kV�Ng��e ���a��yܱ*m_Ҝ�G��zz���g��߳�W�>2_�����b�ZDUg��7ZHҸ�A�y��:o���E{�'�mj��.[�}�>�4��3�`�2T֐S_�&WV���h��t{u� g�`s1�Wz�f�����=�EG��������ޮ�}��8��'E������41���ז��ͅމ]B�γ��Oq��*6���7�<��zxo`u�T9�3"�vrU!�u�uj��f/w��A��fzQ�QZhtF[���*zm���|������2o���7��Y�{�Փ8}B�ނoV�2O}���a��D	X`�M���T��}�7]U�5>��}!̃�p�=R*�WaZ�ʤsk�x(n����Ī�s^��\~���?V�;������J[���2�V^]�u�:"����^vՉ�>�X�y�#.=,�W���_Ąs��e}���cY����L�� [��_$`v©GW�'�굯��ϺRP�;EN�������H1��L�Q����boRm]B4�ggJ�%�ym~��ìd�&y F�B 	������ �����n�A��Pޗ:��rfhNuc��A�lԩ��Г�W�=�m^�V��X�h����jz#��z��^�9'-K��/�d��'���)w���v�$���DK�P����*u�K�l�Sw	b��Xl��O��c䇶�E�I���?��x�����������F*=J�),���6�.<3�_���wb1J5S{[}"�g7K2��}8hk�������I�۠��ޫ��p�:�{!�>+�~v��{���^��w�k�+��T�vY'A�)b}2���ʉn�Џ5�~��3j���]eu�N�@�s\���w[�х�'Mid�<��Ej븞#'�*F�/��u�;�S}�]^����gr=�#qʈ�êa�d��@�_I@HJ�v��bC��]4ViJ������uF�y\U�WZG��+�>�gu���f��,�B����٘;�^�{�]��qjtZ,{�ϑ�z�6ᾶ�qͮe���p��=q�|d^D��[�T��e����S��Eq�=񩆮"�Zd\V��w��q�W#o��}ܬ�s�q��&g��M���ϳI;b��qo�z��|�K�<~�p�¥���l�#����3(�WG7�õՄ%���k �b�jI���c�G=�ėw��]��sP#��;�O����OU���>]��8v��HnWu:�8�ނ[y)��:�����us��b�ZN��*�ݯi��#�3�}�*%�u����A�k���T���]�	x-#��n��!�y���:� ��]�5
Y;��1�{^�Z�S��ۢx~���
���{x�!�ܪ��wPn!��o�yV/{*AG�^�p}0�"z�����tr�#�:'��a�)����ˋk�������GnTN�C�e��&��KMA�C�?s6j����ίp\��VW
��^'�i�7�ڎ�5�0��u=������y����M�4��:��"�x2��T���r����\M�)`R�,�.�g��qY^��%��̝�8?��&�c�O����+�˲���<O�fb��^�."�Mx�T��S�y�/���s���E��x�g�]J��<پ�wZ7N|�bo�S���'���,4gj+�ut�� 6��؇��mgz.�u�T�x��i�3�&unPk����&+|'ZC>gĝ$O�U9���j�W^��� ��sը+�pd�w���s�Tv����u�i��:ᦧB߁�U)`��'�w�[���nz�0�QѺ:lwͦ�v�D�j��:˧}׶�A�<a跉S&:�ܕ5->�$Ê�mS�2�X]�@�$wMa�}����N'"4�v�g����e����!;�(Wg����A�*^a��=H���F��7"�/��ʌ��ll���n�� ���n�7�� Lɩ��9r�͵W�z�COp~��]'���M2�M�}�Љ!Fng�w�n[S(�`:2A�L:�������{oy�x{����wc�H�A]�xk]�/����ZsV��d�g����.7��e���.�/hɈ�.�PZC�]�*)*|9^k,:�<�5��V���ҾL+!n�@�\���:�i����Z�f��u��̐a�ΤN��mpCOj=$p�]@b�H@ֱS����e1n��v�m�$ƷKet���\�����}a�L׳����p�1�)ZZ�=�̮����5�ukK���6�	� +۹�z��@��(�oNyf-�H.س���PY�5cj�8%եuݬQ�yV��G�N���G�H�;���\j�]��[��g=-�t
�����=���N����x{	.\���������_G��v�)�pM�JGS��vŽo��	�2�"�z��Z��<)�2�;räSSr'�0���
2��?d~�=o��č���P�zF�;�T���;ti�O�|��*B�A]�CwW�
D ��B�e��
�8 VXò��ք��v;9�I�)�
AV3C)�rF���z0�v�f���2��Ҩ�޲�a���x#�o6��jHc�s�i�c�U���Sf<o�n�I�f�� �����R{h��^�5�kc/�ێ��v���Ŧ4Jm�:����J�A��<&��qօ�SW����o3��cYe�KsW�8-�5)�>�Ɨ�ҭ�;���H�i�[���x��MCf��[��D����;���l+y�7�(�9�%�g~�&\(���D�����Y?�^�LMG�m�UK~�Ǹ��j��Ͱ�ut�T��s6TPv�s"�Q�?qXs� �(t"$5��Lir�rwv����5�:�K���{�-��5Ե���Y��L�n�a"��1����3�ʼ�Q��5'cU�;Qon���=;��$
�us�J=�w4��Ah�#-�y�{/-/j���lO�:Y�hj�&c<���"4q�Z)��큨wf�N��rȨ��;�\`ɑ�V��Vn�#8��)�q��]��x�앣�%��9�dg��ɜH�逭��;��ִ���K��O.G1����,����Q7��D�m�W'�a��@�e�A��o=��8򸠺��n�K�[K����Bn�+s8,�jN0q�0�H�f�ư�e�#4�S����[#�85�Z�n$6�fgզ����w\�f�1�$~:O�н���\�O{3#�}*�f�-=2̥C�_(���y4��0��_m��E��)�G�_j�����������-ɡX�sC���9�u/uuiY�]B�p�IDYjqEwp�9�T�bD���s�F{��j�%�2�ꑄa$f���D��D�.�R�$;�p�a����8�J%Գ�x9tq�u59*I��(�Q+V�{�QQʭBfEU���QHYX�n�TC��̹W�,rH!�s.�s*(��[13�*/S����$�0�(��ji�f{�W��8�͐�Fa�LV�L���kB�H�Lͮ��QL�'-,��̂�DeU��y9�9\�BU�T�;�I�����B���/!�J"�"Ȱ��I�W*���- �H���2�6r�5�X�4T�ݹn�W'pwEI� ����m�pHΜ��T��,�*Ԣ�s�벩u�<Τ����H$h�O5��v����Jr��B���f���)�"�>텗��G�VeY}1��}�s�h����N9QI�y��ob��*9�տ���NX�Ge�����밴K+ǽ�8��+�\9�]�6
"�^=�č̛����,�#�K�3�'�P=)<�q���������Ϥx������{���J˪7�<ouS�1�rx�l7��&K{$_�g��
pm�޴4g�띱�����vr�O���vjɪ[�S#��{���
ةE`4$�\����g������:Ƿ#�ˍ��П���5��٤�]s���:|8�}8C�q5�iu'�yR>�������D-�	u�}����)�Lw=��q��z:x�A� �H7��'���6&R�]!�ǝ^�أ�u��\}g!���k�qϝT�g��Ϻ�����\i�(�ӝ��]T������]�h��ٖ�{�8=u/���+�o���+���d7�h�G�F��<���Q�H~�e�����J��or�$Ζ0�t@ɍ�8�T�>�֓��Lu�m�p�n������	s��	�սW�v�/rv	��X"|���ǋKw>T��n��~տ+w��}p��<�[�p#|�-�Xr�g[�R��B�)뇠Ez�も�0Z/���LȮ�rfTВr��D��6:9�:*�u�j�sY�j�=��d���w��,gQ+�����]G3VX���i��;���8�Z��s��Q�RsɲR��獩�)S�}2��#+�s��wU��ظ:���u���d~�R<oM�9��f{s�֍�{���bǶA� ww�d���Wt����7�V�ȇ���3g$��'��%٨3�~o�X���W�;5��+��랁�p�¡�L�������k��x�?~;/zb���� "&�u�������?f�_�k�ǿPJ�ҍ�U��^[]Xx7������9��|VG[���3zkz��+�Wdוv����{�H=Pg���E���|1]Բ��
�]|4drL_zOf�z�����6��ӎ/��W�o�+�rx�/`@K�F�����.��/���j���>��e[�{�J�gy�y�C�P�\�j4����9��F����<��[��R���m���W�ߩ������m�����;�RNwI�UaL�5@	H�E��Њ�{�<��T��F�s5�e>�j<��څF�7���tw{���Ϻ���d���F�<n�����V�2����:r銸�I	Oq���
�����7�<�㇧��|`i�ȵ�#�T�"������Ԇ�R�O�;��T8���'�>�r���cW�zmupNI��8TP��B�I�{5~�M8��D��˹\��ם�k�$*$�e]��G�����QY�+_92����cx��o&��I~�Oq���N�|1V��W�š��u�l����#����~��GB+�j�X�����ϒ��ᮨ�|��Ŷ�̗Ǡ{���e�����댫~#6ڃ��C*��Xx�Pɇ�%a��63��]���Lm���|�]�0'���[~[P)�9{.4�L�C��'y�
�ʑZx�B����-��x�R����U��9�c%�CIs*�����J�0g�a9����3)��O�C�U�w2/=,�T@8����++���l��W��f��:�zKf�m��U����.9�D����Q�9'.6X>>��^�xe=۷��9��W0�"�����(�K��Σ�D��d�C��;���Y�4���J1_�&����b����,���P&P۩T|,�P�8},p<n�>��c�q���
.n�xH�ytn�t�t=ʞ7Y-\c(����I�F۠ˍ��:x�?��\!�Vgf�̯ø)"��<�3��C_z��ĝ�0�����ڥ=9�*%�;yb����*ǲs���ZWXLG:=�m��;ND��V.J4�$��0�I�P���l��j��$>���t*����)��}���b����*ޫ*���ӺVm�Q9�ܤ��Ƴ7���f��o,�[��.�/Rf�\lw���\
Y�0O=֭�7�d{�u���f���;���\�=�����T��X�6����eޮ0`_D��uǵ�U�ܼ��T�=�����d�?u�o��Dz��0��UB�)��,���3%j��0�WP=�Y^顈��.�OGL�����:������3P�Ag�4F���Fe�t��;zs�މ� �,��̱�"��Agκ�1��O���A��p���7Ƿ�l��Mͽ�<��̎��<��50ݍ�&"Jjh_ԝ.;�fxu����毃<��{+ɝ|�R�u�3Z��H�d���d
�uJx����.��;�*%�u���o�;��8N?G��j�o�{�}q�Ty��;[�'���_q�>��r�v�M�ʂ�}���\v�/#d{Q޽��֬qpz/>�[ήM�>����4�@yV/{*A�<J������W��ՙW�b�:j�$sQ��]8{��\Z>�/M�.7�h�y���;r�u�]B=�9l�(��c�E��2z�֮z��|2Xs��z�i:s�/��ڸ�5�0�O����'n?Vx�>�B��{�ٸ3�ɜ��^,����n���5h��#�h���Z��W�Y�������gxx���v����<3�)S[�5sq�l�O_T�I���.Z�\��r0w�a�K�	�r9E ��#R����4s��.v,���:Ď�9.D������BoP�f�-!��7;1��v�󔧳��3����]�@���;�^��{��턵����f+���Y>�0�>ȱq�^2\��G��_/;|d�Jt'�{f{+���U�C��+��N�ۙ��Yd�0���v���T�F۠ڿY��B>�u���H��p��Gw�wN����u�D�h���H�ܲN�����UC���j}{������z%u���	���Ǻ{v����u��9�[��D�hV��K��(��h��Οv{޼��M��@�TmӪ�,z]O����x�r�����H��r�{�m�^��oX9(Q����f����W`(� fq��)��-�<�s���B�:�����m�0�{�g�vs��^�>�^����tl�1�.K5
	QtDĖ�H����Ͻς���hh���lUVzR3,��1�;�.Ҳ�s�js�'�;�����P̖j��:LLJ��7����u~!��������z��4'�`��V��O1����>�������Hȗ��VK�`K�ʵ=�*�M������LTm�j�M�wR������2��B�N��2��[���S�d����Y6���!��+[���6�N���v6l���kx��� aS[}�n9��<�h�F=��TQ���V \.���y%�);��񈕽/�-w@^�+;�\�!����e�6�'y�شM�7RM��ܻ<'c�t�zF�X�:��L=��_�Ʒק�[�%�����]����M�9|L��}���b�Od�C��eef�9���l���t�NXs��T�	�mp�������'�h�y�WI��O	�(g�jaۍ�ңe����2���(�C&�����T����u����3n�87=닙��;�O����Z�u<-N'4'���
]�8�TKw�-�&����+��k넚�0L���r�FU_{'j�
�`�U��C��/>�V7N��}s"��Y>�0�SNb����#���m�߯�����@| ?7�"Y]�_]Fv�B�H,YZ+6rO����2���[�f8{���37���3=yX�J����]ɾ�P9g����o��q��ݗ�εq��vZ���37����;�������'%ᮂ�
ⶩL��ۡ.^��hoW}�<{�!��+>�w��ʊ�W��=� lyj�l��2�E� �`H-.���Y�,�sB����܇Sl��ۦ�,W��o����mF��ן��ͳ��F�$�2��R�pv[s��u���E	�(x��6�/�>c~ ��\�a�(���c[������k��îߣo��.zYՓ)<�z1�SZD�ō�ņ�F��f�)o������y�l�u�dV�ˢNutK&��s� �c�|�u�؀��1������Y��&f(9�̊�����g�O2�+q�������gb1�ʭ��'�l�oP�Wԁ�r����A���BI|� ���6�H�]Gn�w��^��QR:2�s�q]<�>�G|���n3����SQd��� 74zH��)eO�.�,�5���@����5F��m��s�}����ׁ��~��3Nd��`�+�A4DL)�`9�y�{�zY�D�T�]*�to�����B�y��+�y�q�'��� �|_��w�`��,ߵ@�~y�S2���f�62\���i�J���H��]ɋm��&W(��¯������*��
ހ�1�'*Ψb�u��?��ޅ�_��jc��wx��o~���);,=[!�2�G{������'o�y�cz�A���=�	��)��E���}{��~��yl�� �29�v��Ϩq���^@j���\����:�}�ZY^x��ډ��U���'ۇ{Н3�3�'�!�n3m��{:e�ǚ��wQ>�e�TF��� ��䠦z�=�#a1?���,��td��%"t�*/s���,��s�w!�Kf��#|缞X�I��FD�)����,����S�k��no���k'�I���gw.������}��*�Fk�x �kp��t��t�2��*9 ƙ�JB��m�nˊ�gl�X�]�
��B�����D�Ѻyp�#��ևh=�'ff_K�ZV?}�#�m(1��~��΀��)�>���|�K��t���^zM]�;,����m�mb1Y�S�YD�2�T:X����7�۠���a��W+��&�\Q�)ףszތ�N���Hv��oLW�r���k�0���U1V�)�ϖeD�ݜ�����WE���nө13��=W��q�������M`\�Pd��Á'�C�����:��&Ǣ��V���=��qW��s��s��;M�r�=q���X��i���@WEΘ5>����+{��ܝ��E�X�9�Q�=I�>���q��G�:i�>�_�`��^�ެ�x��#NԪ"g�h66_=�f|���H,u�َ9�̸=:��P�96�����Fx]b�_�9�\�$x�)W�Z��G�Pk�k9�Ԍ�J�b�2�w^2���IV����㧠��I�Q�)Ө�R�ځ3�N኉{]Fp�齄���eUؓ�UBW�:����dX��}θ����og��`��A�,��d=#�c#=5��w����N��A����'1s����܅ҥAMe*p�"uF觻Y��Z�v�d��|]r9l*��jY�:u�@�����۴i���>G��({�~j�t�|��x��M��JS;R;�X1��rY�K��i��qcV�tc�X!�]Wi�j��Ǣ7���:�8�@r�}|���\oeH4��P0=7\cA�TjTԤ-�_N �E�Ք�g�iZTF�zsj���zsϨ�9ە���.��1�:n���Q^��{Ag�΍����S��z!]='NG�_��WY���V�~�w��5D�cҮ;�zY�_�W��g��E[iΆ�G�_�䭏�;��+��t�8]��j��9l����!l�o^m��j���î�l��*�zެ�T��S$
���O��M,���>�ՙ����T;�7K��~�ʟ�[�xj�C��7��'u|�#oU��紤9\\��v݈y���"ߥwN�����Hp���h��R=qr�:k�+��F�}8��vbYW~�U,�Ί�&���bY����x7��s�O�G����u�r"n�+�^�gjj&-�����a�f!�}�>b�u�M�u3ǫ��w'}��<_��t�;y���V�n�j+a.��.� ��e�0�3p6[,g�׸�t�J:�����m݌������Ә����=��>~[C�`�أa�����}�L�=���ɚJ�Dw6��		�p�YX��#��fu�8�0�f0�F�U���hPᡐc�(H��/�S�_k��"��j����$��{f�c��^]���t��Ȇ���X�Ps�:��;�rY����D�%��. �s�>
����O{���!Oz���NkH��9Ϻ�o��-';������d�P��	�beum���lܛ#�����P��wv���lgOR'�t�q7��q��P�ze@!�4��|�ϠJ�̋����Az
uFY�}|��q��ǵ5}&���=�������ΩɚR�ѕt����½�Y�6�m��g��௥�𫈬���ĥ鶻���IQ��2m�P��yv9�f�j˚��L[���r��fL���4����p�_b�����~���No�?Ok��۰W?~���9H�l����~ipCdmT�bk�߬��͟}��U2a����wS�>�֓���_ٷ~��s�eIL̏r�snQP�U�К��_�U���Ղ�.ʜ>��at��ev�.|5��5Kif�on^ :;�ֆ}=]~�>}[������ʑ��s=�xh�{��r�OU@���Vqo|������{ z��^��#"���=Sޝ�spL��:�X�ݯ�k��<{�^�c�x��.f���q:i�;)��;��q`���B�7��Ꮞ|SMԣ�f�2�҅��gޫ��r�F�y�V?b���_iӻ�k��/k�8!$�EB~w��i(�;��r���E�G�k�/��5�%���͹{�6�}����e��g����e��������[��롆G�m���e�a��"�&����q�Xǎ䀫��g�����zU�ɹ};��vJK5�k�;K��j5���mpR���58^�7���2_XgX�d�,�A��v>��
�:����s��������Nz�f�"L!�<�:��lF��(eI���T/�yXn��4)�{XwO�I���Ck.qH���p�7U�����{{!���)>�F��u�8��g�.4�����ֈ7vz5���Qc�mM��Ww�==�Ц2�߬!t�v*w6��d"��5���;�j�)���r�r��XXy���Iܕm���[�ϑ�K'E���5r�*��wmMŐ�s�3�o:� U�c��ǝc1�h3�v
EU�d9�)/y�@���e��[��m'JdWJwv�h5]k��4	�o8{\4��=ķ���.m�p�l_S&n^%�w%�T<�q� }dR��i���j]� �r�����Y��t�;�<I��͎9�T��U*Σг���*��3x�ʟd#���s��tj�۵�Z�	�VV},��{���A Y�Hv����ӏ�r����ۙp=V~]+��{6��mv�z�K�Y��ysn�}ش�j�V�+�@8랫���%޳���v|>Cm��q�؈ԮXB��b�OV���R�YG_K�9]d�rv*ZK�W��֘[x�
�ҵ(V����8�#w1�%N���#�=/�m�a�J�{sq�i�ec���r�/��x�-Jf*q�z'OtZ��֮E�f�����T��E^5�Ϋ�V�[���K�m�"�n\f�%��Qud�O���:�,��u\h#*ҙ��*���d�!�T[�d�m=�)еc�8"�3n{� �����S��͓0���9��K�xu���p�%��=�5
6��>�ס�G9"� p۫�m�u�;��ͬ��D�{\nt��=Yx�$�}t�ʽ���l3L6�#K�)�7MnJ�	����{�6�q���c2e=�9(���m��V�g9��R�w¬�Y{��r�`��ٻO��2��k.T����iZ�*l��d���f�K�z����ھ"���I9Q:\��bh3����|YP�Ȅ*���fI[eX���f@�U�-��-�������|1S2��zP�qZ�]�I�C��(K��y��f��s*Ʊ9i6�T魣.,�]��/Um�&ғ.�V>p�3:X̾�K�.�Q����ҋ_/��2m���r���?!�3��q���>�1.�6T�,{�b��㙕*� ��7�`�6H���.Qh"�S'�U��0�05BY����H�9�U���n��%�r��B��a�tLΖX�ФRd�F����K-����r�W'�$BB�TJ2�wr�3H���{��3�I�QB��Q-D-\���:A�*�!�2�"�]:⸎JdU!�G$�I��0�T�̃+��4�ˡQĪ,.S�^j���%	�2RC�¼Iԍ3	E�w'g���T�UZ`,/v��*�'S��;DLʳg0S�U����Y��j�VZ�e$�$2)=�s��%^��c�zI���sUH�k���ye��Fb��H5��T)ea����P���ul�TsnG��bHQF��S�{�JK5@� �h��UOv��24R2���tS$C-�&A5N�QB����[$E�)�wP�ey��RR�~?�����{�H�fr�>ɝ�&d���x��hb����<vE��i�j*7bE���@[�ݢ�BN��'q��F�}�q1K^��Y_���g�2��n�N�P9�g��t�;����ˇ��Z����C����w�]~�̻�v�$���$���	�vg�c�n��{�A�������/�gbq�	�5Ri���[�(�]�X{N�nܐv�2��y.���w2λub���9��T�N'����� ��Ώ��w�f�Ê%8��`8.����j�ཀ:uȍ���~�"j��
���O3�z����@��s`\�i��&u��>ڣT��������?QO�:�#q����X�GO���>�4��;��_U15d�@ ܕ�^��u;9�.�b�+�;S��+JΈf����*5��ˎ�����=��o�}��/��ϧ��.fǼ��}�Z��ɶz Դl�"b%�B�)SGF�|n;P��毤�t�'��OI�=�ǹ`����i���;枤��?�'�J�~����b�/�qrK�Qu��ܘ�b���������Z�@l�'�N��ϠuFTF�Y�iN�{��ĵ��Ȋ��y�c}@�p�$���Pn�`;=E�M斡�o�nh<�� t�4
�/Z~�\mm��^Qp�{
�[6Ƿh���+Z��[w�L���=���B�
��:�Ʃ +�F�q����":�7�g=:&K7zl�9�%�n4����IFz�ڭM�Oh���Hﳺ����O;q�<,_��RDl�*�0��O�k�o�l*;�S�a+M���N/՞#����u���6��ds��9�y�2��N�}�k2�e�Y>��q3P �~�z�?���	t_VWq��^'��qͧ\���L��F����O��e�o�oT����,��F�-��/�g�h��m�Ux���l����].<Nu�q�Σw��鞬˽���#oq��=�G�2�d��L��N��EOQ�N�),���7�t��%���&9��������<پ���n�F3ng��Y<��,e:X���;NC*=�AA���P|Ӝ�;{�ߔ�Z`WP!1��s�|VG]!ۅ_�iC�gĞtU{�eG�(�-4���W�}6�;z�W�]��}~�'��=�m��c��M΅b�P�$��3�5t8�*j����V��Yђ�Q]v���ۊ�u�w��s����g*#���`�*���V���g���Vx
�nb Jz"O����l�^G�X�9�Wq�֑�s��P�G����#Ր.����?]<ʷ��e��:��g�E/v/�(�(��ƀ�˧
�_^!sj�T�a.�U�HR)%��k\_�>ҩO��&�ř�m����A��˔��<��4c�ǔ��
k���7��D=�sA�]|E�C��P
�C�XD��\�J殕rp���$�j��3�:d; i�}艖�A����ǽϑz�P뭳��fL����X�z�.;���!�	�S���������I��d���M�N��3ïܮF�fJ�&���Óه�4Ԍv��"O���:� 9s����&au��0^�Q�Ւ���]F)X tȰ���'v�\����C���w"�\Od�zE��}w �)d����P�\�-wD��_H^��z%ua��\v����v�}���i�
y��{ <��� �)�S��&����'�v��4)�986�׼n+Ҵ�>�/M�m���o����}@t��յ���F�~Qq�EK��K�~��Y�;���9(+���w���
��:s�/��ڸ�s]�	�����������Y��^h}]���/�6�����3��|=>�*r���?��yS���#��b�u��ꜜ�S��z|��guX����1�s>>E����,N��T����u�����k�mz���_##>�]|G]>+��N��ʟ���fa�;P��r�~M�bT�~�eL������^�"���*d����,#���c6�)[ۯ�!��sCٵk`��;p��&���Gy�٨��
,�ע��Y�仩�BJ����� ��I5�S��9с��,��eV���ûӜ]fnO|]g%f'�oK��a.���{;$f����߯���T!�wQһ�}��1�#����V���[g< ���=� /������^V�����Ϫ6��ɸ��BY��뻇�7��{I�ٝP��u��u�Ug�>�}t���ע�/z�	]Ӏ��3�G)��[T����.�����b�:���z}�q�\w�	{2D���ܜ�s��=�xa��7�l�( r�2��
W�-�2<��":�����0W�ti3e�]}Yz� =<���*����Y��)D�%�_����H���n�+J:�-�� wV;T�T�O!��Z�����|7����q������j�� 7I���մCZ'���S��GV������y_��</����ԉ�ド}Ӏ:u�s;���A��u%�G<���Fu�\GD�ӣqNR;y	\w�91Q����wu {W 7��� s.L՛�0G�z��^ս��N{��~�$��fq��}+k®++�픋�Mw�9󪒣�&M��7��s��w��#�iA��s'�َ*h��ہӁ�^8'���m=7�������1;}>?8��鎁0c��P+M7��	�&���̝I&x:�K��uՀ�:g���,�S:J��~Z�U�0�B����>��C���爆����;����|\���|KFTEf�z#������¡5��]d3/��U�[�t�λ���^�P���uy�qNj��g֏�Vʍ �))�	�s�Y����q��U&��z�����n��Ϸi�]]U�CY�����������+��V'oՂ�.ʜ>��A�]P'�0H�gp�,�R��u���~jr.�\����5|2%�_�ϡ�o�����:5~[��vx��!�H��O����gp����Ε�ՕL�T�D�� ���$e9]�z�/�;� �΍�6rO�zVʛ��
�����7�%��=��2�6�Uܛ۞������{��l�=���εq��{z�����]#�zQ��<�|�rO���Β�΂\<�/�V����u���<��\zO�fo@W��,o/V��F�h�D+WrޚGp�7�Aڃ,	�E���s�!fT���
�Ď�5�7^[]H�+�X�\=��x�w�f�ÿ��F��x���&K�@�ۛݫRl]�.�^��c�#z�_�E�������F�q�Ht�Q,�" r�0í�B�uw���Q�����zN��1��{��#��!����w�>�4���=q�LMC�.o��o�_m��8�;���ח�d7nb����l�¢H�OZ�~<mc8���wr���K��G*�\R���-�˹G��-}����;����90L�q�w�,d��HU�&�E�F"y�{Е6���)�ݭ��s��ُ�^�җb .F;�j�7g��y��#qP����/�}�����^���~�3�p�ђ��yw�en��W�FY$�"JG���P��M��P��毤���Ȟ!x�@[�\��H�d��k�TO� ��y2�O��^]����x֥OM�]Dw�R=BV>��ݢ��Ly'FOwO@���3OQ�rd�D�{b{TK^����i�J��L��S�n(�=#;��x��R-�2�`O��y�b�7����U@ɇ�}���q�LX�ua�̸:�����p�������cE�m���NG�P�/��O����b�fT��d�>22�5ٷ4�/ٝt���z:�qYI'�N-���m��u]�����y�Ds�����1�^��]yxk)+���:X>>���PT�u�Ux���E�D/s���].<Nu�q޺P����Ц/{4���"}�w�X�Fɟ�]'��,e	�
���>i��#ŀ���b�]�*̧Yٳ+h�����u�g�u��ygZZX�?�U����:�;NC.���{�MĐ=�_t�<�
��`2`S�h���+�ū�I��>�ut���P����n���䮷�b5Fz����E{�i�kK�O�q/mQUo���ǜ��:�/��q���Y�C��m��Ih���
΄�7Xk�dٗ+V��MR�K��~���_ߴup��|w�t?t�1Kr���$��Ơʦ*�����OW�v*��^�Hz%u˞��Q;qo,Cς���=������[�&�B���EI]tх��F_�ǽM�޼��Ny1�\��{w�㯶�:���s��w� w���Dz�S��]lFNqVy7��+���� �I����e��άyw��:��98����[kF�{�Y���Z�C���������WXTTVE��#�%�X��Ǽ�z�s�َ���x�Z��T�O)Z��B��<zw��uA��2)̖��50ݍ�&J�4.���X<;�Q�~�J+�E�)�ꦄ�oա�Z�����\�VD�$�؉{]G��g�R��w�3nϒ����M�u08>URSĸe���q�S�N������eJ2j�{:-e�^���O�"+ґ���w��޾�\��}@9��_����\F�T�B�Z�^�xC�����ݖ?Px�Ʒ��W���>�/M�m���o���P.r>���u��_�gX���?��k��3����݇�\�Y����^�dt��`�n��[$@Þ^;��he��g�iE�E�����̿u�n���S2[$��VLܐ]��!F1�;�%B�j̏qg��ʝt�v�-����h������)Z����j<��C^����ԔQ���e��^����X��;���t��9�|n#6��g��y�{��ڽ/�����E@��s�]���?36}�?���K��Z=t�3�ˏ�����._���[C�s��	f籴���g��OWvp>����c걻�Y�+;*|mO�fa�E�VMx�TP[����0x-O�j���pt���o������s�|R��x�s������!��(9%�%W-Yו�d��ޮ۹7֨��؇�=�d_�һ�}��<�8,��ndz�WI
1sJ�赈4I���k�=P�+f����Y~uP�|7��r#�O�mC�n�*�(��w��E��U{ z<�������@���45P�f[�	��񾾫rw�s�Rx�>\\M�ģYosxݽ��t{����]�6
4����R�����w^��ԅq����/;u�ׯ�I�h�,'�OO�vۨ9�T�;%��A*=DLIod�;+�����1LG��-t�U���}�=�4t�t�o���-&���>7]Q5�2Y�����Gј�@��
(��!����ݾG�Me�[<
�{�G��t���S��;"���m��7f�t���� `�C��Gwv��ڐ��r�f�<�ܸ@�
%��R�:�{�����%���5
�%��긝�sF�P����Wy�W�����jsm8�%uQ�];�l9�j<�H����OR'�t�q/�p�뉨s=2�����i^��w�]
g�I)R�(���T>+���D&���wu { up{�6ϻ���>�/lUX���K�/�L�N�Fg��Ȟ���\v�BR��]��j����ɬ�׳;�u%���W��{;jF���as%gdYc�N%x��y����OM뼸w5�U�
�:F�#��wf;yEt���𝿟_���{��ĩV���޻���;��@��be�vr���Ir3���4g��#>{�7��9U��M��*pߋ����'<a��ߘo)�Ǉ��u3ƽ\�� TE���K��q�Gϫx�sC�;�:3�dZ,���>��fWm﫳K�g��Tzⲫ��g�+>� ���$g�NWt����N�t�W2�_V�]l��~�fr;�C?,�.�����hK�y��nS�v�ĳ�3�wP�U|�z.̶�m�\pa�5��%tnv�Q�9'��-�'j&Pt&t;�ڮ����B\��z�<�����ɝ�C���j��I�+�;8���9RF�.�5�����cz��Yf�ٴ5Jq�GS%��t��wY~����0g'���{%is��`���[T�1�,�| �n�$�x�ŻK�p��U�/���dS-�]�]��Vmz���^Ej9��X� 8��=�r���Q�Pf����F��$�`�,\Vҹ��Y����7X�g����hĞ�{hhϹ�=��G��>w��{�(�<IU���L��n�U����+�G�X�_zԵSz:�4P���_�}�k�^ޡ�:�>6��;�\�j9H�F���Z���sEos����9o hzy�Q�n򸮞V���r;�Ԇ�y�Dz��$�z��oVO�ϳ���^�a��� jh�"~�u���h���5F��Q��6x��l�A����y\3!TWes�3�
��9��r��5�$�D�����K�B�"�4tj�q�Tm��_I����.j�O���׵֩���O��ȁՀTC�s2gd�U���?��#��5}ݾ��F�����Ӯ�,����s�2n;��od@uK~���~��%!^�?S=̻���CFf�s&�:�X��o���ۈ޻��'�r/Ps7������xX������U@ɇ�R�����e-�v-lb�c�1sr��Et�-{U��q�y|3�Wi���e�Չ�ߟz�Z̩�:�g��w��9��lY�������5s���.� 䁭����:���,Cd	4�����v�>Z��~;��c�C�:����wDp��%a��V�il֮Hܬ��9���})'�ff�P��+��KL��n� �3Zj_lc%����v�)wl�b�-\`�\���}i�l�{N��Y���ؓ�B�`c6R�ݕ�%@G}7����3�i*��1K��y��6�5XÁ�'��bm)9�[9��u��ǀ�6� .m�S�WN<���2�5�<1=��V�v��� � T��lv8m������m�W¬Y�R"V�m��QW�K�ݗ�)�c���nds]�5Yv'T���,X��X�z��#�T�S��o5�ō�7h	%&ZV\��]�.,kˉ�i�fa�k��/e:M���>�ۅ�z�q�}w\#��bƺx�i�&Ő�GE�=A���y�4c�V����0����9V��O=l�%�N}=UJ(}K��AL1�O�)>պL~�ZO��r(pYװ�ÅER�S�+2��;�ДW�ӝy�U�,̌�m���o�p���?�5��wJ;��8�q��\�i[��=b��+m�u�ũ����%�H/y�6}_�[�6z�t&n;�e;�Ct�|*AMJ	C����n��ZN��V4���`�v��{�yP����W�<�e�:K��7�4��|j�2_T
J=��^ǎ��i��dB>n�wq:�o���u�SNޖ�@����(�K�j�&��%w �'��˭��B��RnnB����4�T��T�1��~b�Ep��I�gP����MG,V���֥����(o�k{MB�^�ᖘb�ޚN�<���j��V�u��3��qk��+C]���Aܧo��C��yy�����)	�w!T�pX��,v�^�Ӗ\��Ko���:�
!f�Q���t�֫	(c�M�(��U��&����qʷ����"0��)��l4�#��۬��"/��B�.ٝ���9������J���B�9�,��r̹�-'{p�$�lZ�儊A̡����%]���	[؅�����ѓ���i����Zz��n�^��Uk�0�e�\���eqK8��:�������cz�@-�勖� R���6�c� h�=�sм�f{�&4J����ҷ=�ԥ�n���94	���:�W� Af:���$��]��9m,4�]��HW#B��̗DP�wL��f�'�y��4�MW6�k|x�͍V��Hk(*Vl�����b�M*�֞�%���}Pd3�܍&H����cO�Én�i�ww�a��q�[`�bb&Ugj����畽�yj��Fxh�=B� =}�5����g�ǫ�W=��+�8x#��ɏ:��DQ��{A�jd�鵋+AΎ]�	���0-Y�Iv�3Oa*�6wm�ʋ����-�������4 �@Q�K��D�DE�=;#c�T�I](tO)����S�tM"�3n�'2�(S���*�H�ĲS�d��V��H�,TQ����S���T�=S��r5�G*��D�R��T����w#�,����-qD���i�Z纹9(�Y^�z�Y!��A{VG��#	,NsK(��'aFeDb�w�R䎆*�R�/"�%4���1CD(���'�����w
�Rԍ(K[*U�n!D�V�T&�:�jE"���$se��YJm,:t�'B8���)45���]=���k��p�e�]Ot(˩!S����$�ݹ��-�nG��d(�'��BQ�B�f̥49TU��N��yfaEF�JmB3+���0�E=[�b����g2��\�\҂R�Ȗ���H�,p�@� ��?|E
[Z���ۢ9&�fM�Ѯ�ͩ�+�Z��5yFd��4��E���A�Z�չ>Z�i�.8g�M�U�\ʾ��];�9z���U�ro+���s<�at�~C���g�{�3���r9�D��@9^���MH�[�����ҁÞ=�3��"��L���Fs�Gt�\x�����7�t��H[�7�j7voǰ�L�\.���c*΅T�4�r���X	nS�sD 6�L�L�W�uW�:�}\��/�����܇X�VnT�ݖO+�,e|�bvg��9f5!{,_���%qr��ڰ��p"߇Wc�|VG]!�i�}r�,x��U{�?��䴩
�b^����B��WU9S��Q.�v��<�.����=������}Lw���Т�G�/[��R��6�D���@���q[M����'����qW��r9��;�{��q���U[��O�>�9tW!^��k�>�U sQ%�!��cKe����qW]i�qZw����{�h���Ϫ��V�*7ѽ�G�:k��Ag!A���s�ƗŌ�sK�z��tz=� ����^�r�洋�f9O����N���Psz����2Z����wh��+�и�N�U���W16��H��R�PJ���~̃����kе���a9����*�%��d���Gش���+>�_vڲ�0;��o2E��u0Nz��>��I���(�@-����|�ԫ��G�M}4;+>ⵎ���bԚ��䖖��+��{/m�}�:���~�|��c>��g��q/ uF@�t�&��v��.�;�<��M�yu��H���WU��Wl�CUï��r8_ϕ܋m�����σ��+��r)d��ߐd�̜��{ox��g�9�-׼r�-����p��k�_�ήN>����i�*Ǯ;c��߷ձ������H=8O��pv�����ϰ��/O#���m��o��W���K��z��R磧}	D�nYئ�#C?R{2��֕���ag���G�珇��t��9��_͵qӍlL�9�����W���"/��tF�e���N����38n������P=>NI��_���}��B��2�u{/^�'���ݐ�DOS��z�8�}V7voLnvT��,�z����O"Ɨ��(��z{|�d.L�ƺ����`T/u�22)���_P��9'EFnT��d��d���;����j�^����tS=z�.)��7��x7��<���WJw]��g�u�{�����t��2��}#:�	,Ԕ�Ut�I��rĲ��C_����<{��p�H�u�냹(��v����3�h��R�C8�v�U�l�W#R~}&����hGLjeO	�f &�T/��
\,	�7�oj9��	�l�)7ںMUiC ���PEi��ͤ:Pݮ�fi�LNYgvoGt:��l|Ihr��wmM��=��.�Ib��ju,�?�_D�xm���K�%�p9T;��nxz]O����x�n�Ϯ������P�f���H��C��Ͳ��Q��9���q����c<��n���j��L�;��)�LT����������#��>����w�,�( %G������Gr&OCe\��t-��]�R�9�W�ֆ��:������-&����uuD�K( ߃����^�3+U�2�ћ�[&:Uң,�_�uw����;c�J'��&�ux��/r��.n�6=W[=��U�:�e�2!�
�tU)h��W��&*6�W�{�P<�W 7�l_aq��G�Q/ S9&p�|8̦l��R��*����l�_������I�^~��w����${C��%?H}��_�{&J0ʑe�l@�������y�x���'�����"�ѝ�]�����M�zxN�ϯ�tu������Ɇ��������*�Q3\��qB��xJ�t��ۿ�uۑ�z���G*�;~�\͜�œ�����f�樰�Ѷ⛕ҹ]K�u���r�����i��ٳ�FV�����I8,�ݰ��8�A����M׭׎m��T6����~X"}�u�O�&��=tj�L}M��'�nv7��/T����V�[Q���L�@%1�fS|N��&�����߼ux�א��_Eew�4���m0��+���e���s��#rtVvT�y��$6\d���DvH����a��*�d�Ĩ�`��Hϩ�u�+���N=]��1��зΧ�9l�E�����v�]o]��.2��c�\Keq�%6�r\u�,3��[}Al�����n7]��9'�邏�(u@���+j�f6��s�z�>��h�q)~�){oޭ�:��_�|�_�G[���7��Gp�7nH;FX93��W<n(i��=�s�Y~�X��u͞��X�����c��v����v���%�x���Y�+����{sٓUKQ��� 3�g��]A����B��_�s��W��x��@��t���,����r	&j��g��R�g�3[�M��l�z��6���\GW,C#�������W��Dz�Ld��<^W�w�񵪯�Ot�� ���&%��ll�{ކj<���*5����-�wQ����x�&�w�T��=v��t�3Nd����͝�&_Rt���P/���
��F<���?\����a�Jfle���v��OݒA�yw	�.P��t��)���٢Of{�w��M���R9"BI���1��|���R�MjoU�]WՆt0��=���w���s2�*d�]+�U���xK�q<yѻ싫����8�=>W~��j|�<�%#:����'�A������s2gg��]p`�s�h^[�����j�5�5�}[֢����}�C��Wrb�m��7��7��_�z̓P�'c=�	�1�j=��fnF��H]���=��+�v��m1����}w#Hs)����<,^�T�Q�Ħ�#L�D`&��=[������@�Fӯx�R����_�y|3��U�|�GO��N��ޫBve�騯w��k.K��Ӥ�����z��er2K�8}e��w�"]W{�}�7��{�1ip�}'��9�4����y|+\䜽�����z|�Ui��\J9��/s��Ώg�\=OT���P���<�s���7T*�5��g��]'��2�P�Ю���Y�C��q�7<����5�d���7�K��/��v�7q�#�3�A�� ��4�R~�1�f��nj��Wl������k�=���ë��������C� �酷2���$�r3����Ԗ��yZ�]�A�V��U��]�Kt�'w_�Gh����P����h������\3���b����'Ӂ�˺�F�{��\Gٵs.���>W��;�����������{�G�����ܕ
�3ҥ�o]�c���|6��_u�tٳX%k�Ur�w��Xd8H��|qҥKcձ�٢U����7��75�$ʾ��e�Ԗ����C��٘䢑�O���߂ M��꼡�����e�۸�=]����9<�r=�if��U�n<���he�Ǩa�/��\6���R �5%�1��o��y�V<�C�W}]i�culR5ƺ�k-;��/O>����=q�L�D9�YP+��D�u���ŏ{��ȫ����q�������Z��Ɋ<���m3>��}�|M����2+�2Z��S��\������7�y뮝Y뾉�
h���
���m��_8�Ş�q/Td��J������q�]/�b͋�s��:'�N��K�z�p��w#��U!�<K�<�q�>��g�.7��H��n�v�UiJ�Ip�����m{�+��v��p������>|����ʇ��i��]DǠL)xn+��t׹D�h��Q&����x/�����/�o:��j���]��¯���c�[��� x7<�*'n9�,!�3~�g�DaaFk+��]='NG�_����;�2�,�t��w��3�c�uo��w���ƙ���x�|O��u9G��ȋ�ƆJ}4+�Fa�/��&*�U��z���-{�ʡo��l��}��t����������Ώw���k+L]�iGK�lc� zO��6���;f1��M�0ǆ���%_2�gܤW"��l���XEB��a��x֥�کŋ�M�_a/����dpϥ���}�u׸���cw>��1_geO���a�ƞ���1����^��gc�~::+&���m �|=L�K��Mu�=R��wHn�����r���A��ݺEb��B�؇I/�f2�6�]ɽ�@7�B�{�ȷ�]ӵ��'�hpG����9��_�����3�/\�}(����U�k��%��z���ޮ��'�cN<[�2�2o3=�wsѺGCW=
�0�&�B���U)�Iڙ`H�P�>��nx;��*:��Wox��g��-*��ҶP�g���{NG�G��p� Ͳ��Q�P@�Pe�!J�66[,n����w��_{:���o{Du�!W]hxg=�h���+;�o�T�;%���I�;�jdN�z�B�����H���g�=�CF}���Οm��|���y�p|o��&��,�?p��J���'lng|'	��Z�F�y�|G������:a�OR'�t�q6���!�y�1�Lz�en���\�ODt�L�	�&%�u�R��ϒ�|n91Q�	��7�H�uG���*�s�ox��6o�~��eA�(����;�X���}���*��!0}q��d�.�׻�mf����-#���+nӔ�V��-�;T��S�h,���C����h�r�a�{0��qT{9;�2ڭ`���	�D�G.����ʏ�,�70�v�͑���ժ��rf��:*��pT�/g½YK��ĥ�k����`0�̸���J���#:���ɒې<����^�ɒ�2��%���Ӂ�EJ�����qC-�N���8^%b��,��X�������s�c>�讓}��;o��tu���<J��\W��~��{������Pu#���'�J'��۴��ۿ�uۑ�=��������P]s6r<Y>�OמRz�3>Y��yz�OF>h¸���piׁ�|���ʸ/��_�ϟV�yάn�����2��h�v֟<5������������*���*�n"�_���`���K;�O}�Q������p#$P�\���8�5��ޱ�)
�6rO��xg�e�;P�+z�M�ܸ�A���{���˸8�D�MK��e�R��wz\./>�W���f�I�I;�C��%�����%W����4��������bD��p�:w��������Q�Pf���e[��`LȰt>�`�Gگt>�U��<ʝ=NhS]\<;�C��gm:��w��0�G>G�*w���(|v��S���G[���\|�o�L�6�g�l������̆,,��h�����6{T�
���/r��e����c���n��C�N�L�z��=�{Mu5ws��lo�tAEMoR�N�l�5�|%��0�S�}[ �t������*s��b}͕��}��ّ<�����}�(t���k�[���K{��M�I���z�I�i�h�q=�0��:NA�\_�G��{��yZ�W#�}Hi9Q.p�^��������}�׸�wʩ���.j s�=$L�Zih�11�W�Ly�7����f,�-C���ي}�m�@u�H��wu����5d����͝�&%�!W�*h���#c�Q3��#:em���U:��EP���[%���zO��σ��sNfEB,���]aV�����	��u��*������twS�ˤ�O�ܘm�+�z�9��l��&�N��&��!�]���A����x{�Wﱯx�9���cn5��a>���Ps7����y�b����nB۲ _e߳=�"�[����Rg���q���p���8��f�(���:�ӑ��8����u���P�v��5%Z
�d_l�>�q���P�'�ڙ~'�i|_ٶ�s=�2o��j��m�T���Z���Q>�ׇ�zrNi�p�/�z|�eV�%q(�|}.�#�~�ks��`ܟ��y��yb
ˊ;�R~��Gc[��쨙|�
�[�)�ڽ5f� hP3OK�M��������T%�[�qb��r��ʽ7w������í��{^<K�U�A�2^�b�8��+�d�K;���ےP"��� x��s9A���mco��EJ"�L
ދ.XL�6Ϻ!�K!Vi��3ผ8K�΅u=G�הʩ����yuŞ��
1S��\x��|R�5"�j�Z��`��?q���򮜵�_�����m�cy<���2��Z�ˍ���W-�up�C�|VG]!ېf��-ʔ{��m��TK�����4�3�"O���Qz���j����2�]÷�!�]��v��>�u�o��ӆ`ם�<�ٷU��`8���Q(�(��f: �0�"��W��x�u��U�;��'���Oμ*�v�V�l�z3������6J�� RC�<[)�Տ#��\VQ~�j�19�^����*���t�q�>}#�^wY�,Ϣ�,�zHؖ�A�/�蕵�}8�����I���ak҇��dt�o������o��\dT9��٩��d�z����+}�����t��\���q�W#y�������8z}ļ�uF@��:�E���U~���or��0���O�]�.�������/c�0�h�ͻ�A'x;O� ` ?���1����6�� �6��l�@m�o�l��`��� m�o�l���cm��6������6��l�}l�@m�o@`����m�o���m���1��@6������6���1��l���d�Md��!H+Q~�Ad����vB�����o��:D�d�4160�k*V���"(T�j�$J�P���J���������QZSm�+[[Rd�6�A��ɶ[V KLլ�6�}��UM��Eh� ��Fm����m��m��[)�aX�����&j�+4k4,���hPb�m6�Y6��;��/�k� ��=�	��Q���wps��Ӊ����Э�	�p:X1@���U�"ma|  �� �P �`���   �p   7��   ـ  ���6j��=�[hV��b�>  ��F[����j�w�{�h�w ����և�� �{;�ޞ�@�������GD͵[e$d� ��4;�oy�:�� ;�z�=�{ހ���C��k�����zw�ں��{`���;<��6�U��1��ӭ� ���*�ϩW�S�q���=t����E5���Itz�w{i�uή���4*�o=��t:h��z��=�]����V�4�  '�}S��݋��� �������{�������7���kڛ�g�
�ږ����q�w��-�{`�*�\u��K�-Z�� �a^��wiN�,m�ֲ�7v���k�u�W+U���]1�m���{a��:�r�j-��:�.�6��$جU��� ���u�Kf��֍4:[vڝ����յev�뙅U�lmn�5��v��vq�Vܺ����9[Zښ�-c@x x�.� ;tpEU:�d�1��Ahj�sMf�8#e�Jt�j�lك� ��{�͊�E��
�ݧ�9��H���]�� ga���9�_        )�aJU*0       E=��*)(F�a� &�"������<�h0 � #& T� JJ��0	�@ ��  J���J	B`i�  	� �&"�@&M4ei5<��f��&�z���*���/�w�����8-��|��d�,��R������a(?`*"��� 4
\PQ~j*��/����D> T0�/�~ϟ�����t~7������G���y�q?�'� �$�� >pP��.@:���.���z"'�D$d@�@PACqO��������c�G�����?����7?���l6�n��m���cmgk;m��8u9��T/ �PB�K�/�B��Ao�PB�@K�E/ �[�P/P�T� 
�^ �x������
^ )x����  �+x���x����x�7��x�7�"���^*x��"�(^�x
�
� �x"����^(#x����� �
�x(%�D/ D�EP�@o�~�m�����cm��m��k;m���m����Y�m����m����lm��l�m��l�m�۷?/�t�Q�~w˥����`\�	���Y���5�xX*�b�M�T�9z��Z��#��O(�9���On�+)2�S"5�--l�ˤ�%�V��Bon+%��e�n85Cxm\z�FK�3�Fn�GRk��oD%��f�bh��vY��v=�D�f�Ջz�X��70��ɩi�1�����T��&�ve�ST�\��.��@�^e�E-6حqL[����n nhɋ"ջ��v���\"��nF^U��K%�{y�T� �Lj݈W٫YZ��zҼ�{���df�Z3���茷5�#�NUąѕGE���yGQw�N`s1Z-�jU�.�]�Cst��%m-ڳ@�W.h@A�`�Fne5�3m7J��o.�Q�7���7V;�I��u[tHBU�CEзz�b�ht#�E�v��e]�C�1�dV!Y�2�1�K�1;���R��`��^�pQ[� ��+�����-,��N���-�ʽL:uz�:�j)�����0pU���Au����1�৆�M��	�elo��/f9voieLM��0�e����;��ckP!R`a,��!6�[�Y �Z���)�D!���F��Wc$��R�R������t�ih�y �[(N�y��e��mm@�kj���n��M�v�ުj�fA�)��b8�Pt����� �v��ĵ������/7��n�&�:�Ӗ0�3oeGtXqn�f��]F)Ï1n��2m�+6�ǣn�a�����T��p�+���ލ�D@j�Q����fT��i-Z�գb֥eɊ;FAE��n�����5�1�wT��&[��S�]�3\���:��g�,��4�Ii�14���n��UlÙn�����9m��li��հ��e3X�Lw����m2��qW[��M�:�n�����AF�����V�V�̫����\�>d��ٻ���<y����)�jwB^��2��,S�f�Z�+��3U�HA7lDv��L��a�{u�wx�ᚷ5�Q[����ѷ��1p�CT��j��43t
<b�t��v�m�D$�w�VB��%��r!E�S���b�R�r�����&`�䭂fQ+d�1�0�(mY+3��lX�.L��H����H]��Q��@-�M�D�>�y���9K$�� �cv��e�I�'v��V:�a`C\�  ��cH�׉�*n�d�ʸ��q�{JV�X��ѷiJ�M9i�q=�{3P�b[�2]��ҧ[��U��A��4�|��/!�zn�aTF���1eB�����Q�|��[y��Wki�m��x����l�?�yJfWme�$�.f��a^���It�졲!1�N�opT�57�U���aQ��G�"F�Lf�Wx�����5�;�[�ۚ�-N�����ۻ�s���Q%,�#i �ٳd�?nLgZ�ŋû�Zt<y$ׯi[�EiN��斨+�7��[u�@ܧ"M�ܨU�f�NEx�<ݣ�dicn1&���TҡWt�Ըs~�"�a�b�U�Y��W��5�M��)�ٙ�a����c%�DJ!@���&`�Ų��� `�ݦ�)p:��;}M�;���3.���u$��d�n���zi,f�y�m�꼔k18q^�k-1V&��T�d���n��J��u�,��H������^�9f��g)L
l�:���X��n����ք�nK��}��4�ѫ(My֦�U
f�շٌ�y/4]kCwhƃ�K3U�1�u�mU��[��u�v�ɴ�E�˵�R�x
����F��.
z��=�K/F��k#�ݍRbT�(�xn�m���b�Lʏ:���Q��iQ�;��N�6�F=K��E�Y/[y[d��nO�������FN,:C��:��T.���T��R�w�(���(#b��Y�%mk�K�"�:��v�-�T����U|���܏�Ci���#���D�eR�=�m���jT��9��f27F����Ȇ�6�U�_�&�Ln��F�̪YH#4k�t3(D��꣏]�r�/�eU��l˛HM�ɧ��kB0�;�[�"-'��'x��s�x�;3LT��W�RЂ�M�n�4j�q����9mҖ��7)轑д�
�X-IdK�Hn�J].����vʌ�&޴�M�uc�N�Lܦc˷�TW�N�%�s^i���Ǩ!"p�,��8/D��b�bparג>x��y@� ���V��6��j�������p�F<�#`�R��'T�L��Ҭ�r���鍳
����)��H���n\T�J�H��16�P�L\����Fm�÷1m��ԋT��Ԭ����@ɰ��Ʋ�<�̴wKO�*mH�l��Z.�hKǊ�.�d���̓j��r-*�*�Yۺ�Q�wj��&8iU�AȠiJ�P�L��r����x�Qܬ���a��В%(�K�ïo*K���Ȭ�P)�D��f��ֈ���ꆠ�Q乙�75(������p<ي�k�mb��捪�XqPu{���9��ZG��ݠS1�5n�x �5��mh����׎��c5�ebh�h^&0諫8�ؐu��m2颰%�!Nh��Hܛ�൚ΧQ�����32J�bT�T�Sz�6l�4��s�t!9*so*�T(��$ꄳf!�Q��]����kڊ�un��a\o2�p�\��74aĢ�n�ee䍤����ٽCq)R�Hd0�/z��N�5H�[��&

\W�$%Fr����B-uc�;,2�Ӻb�C~��իV&�+izԷO!�MCF�8��$�vٱE�R��1�ȷ��ٺ
"ԧ��tep2�{B�Y�4�
I�SX17Sd�͙�6��~v&,?d��qY�&���FB� @��NSdf��z�^n[��rG�j�Å&e��OE驃lkhɘ킮�l�ٰ�mл�N���H��̋Q����*��vJ7Y� Ř��-��{p˘�6 C7s۱{K#k*:A,\NS�H\�KJ�������XE�M�u���uW�Fږ�,�����uS-�%�2��L�E}Z�:�[���j-�V�XՁ�]Yuӥ�L�n�,��OTAi�(1k�E�.TN�X�`P=�0�|�wn�+]'l��lJ<�P`���Zh����-��%E��t.�,<f7LI �7%h`eH�I.�b��O,�FPh�+�ve�r�=?&�2����-��x����ր�n�J�me�ehx)��ĥ����4f�����l%\Wz/��"�wv�ऺI��ѱfު�ʹJ2>�o�U��O�%d��(�f��\�����E�DS�܇V�4���}�ONn�������U��-Pt��$�	f�eڽ��\�{����o�I��jê�;{���0����Lr�"��95��W���-�k$W��v����J(#YY�ƈ��1J[��H�i�o%=E�畵�r��KHëD*d�M��əV��11t�V
��#��#��i�ڂZ�����b�W6���᫡��1�j�O�kr���k݁V�VݹYOULk��9�F��+�UfY�^��Y+7i;Q�Uf*9[�+y*Z�v�@9t��h�y2�Ɍ�N��Xx�rT��Tw��K�[�Hi*1^9��(j����1�ɭiP�Ǩ��:�3"M9�oc6�U��w�nܩ�em�$���X�Y�l��%��������׺�䊑tne	�J�) ��#���g,�.���^;�$fܻu��jK:���J�)�˔��鵷q�=h������ZZ�#xN��-�W�7U�q����eCld[b��$	ő16��2�Qm�h3ut�pe%y�aB�(.�7%�`�t��u�H��aMaF �Al%H�X	�y{��R���$�z�R��`��0�ݡo�#W��(���"�h7s�7NH�õ��I�Za7�.���k��f�lA��S�$��B�ˍ��d�Dqf�i*�^ |1��vST_jd��kv�nw IX�7PKdD
82��YRLz�{{��d�6=�:[���-V�d��6fݛ��m+qu�N�j�Ϩ��ԇ�ԦK;�/p���GI�61�̥OH:��c����e`n��5Vk��mV2�m�k��d�E8Y�[u��ϋn�4��ZFS*�jrm=O$?]�: ۗ�kD�FFbxn�����<�e4l<�u�A�EZAL�@�{A�*�M�
��Rq�62�G�m��ϤԬc��sX�{q��%�����5f�/뗚��42���$Rvq��4	�
-��ZDKQ�-�%|@�)f]�%2��Ђ�whޱf"A1�ݍ�ߗ{�c���Q)���=�0YD'F#*8�,��;�[��6-d��S$�z�CZ�]F��#���ڵ_~��x��y�M��~����y�����|�����(�@���~���r��Mԅ�F�i>N��x|~_-<(�h�Ѭڴ��tlj����wU���;c���I�m��u��%�%!ǚ��ó^�[��EZ
s.����c�w2&�x�^�� �ֳGb��d�u�����-7���&4YOs��+�,^��w,8��Wl\�[�o������}�2�g� M��,BY�����Vԇ������SCFWVW�:��Y���ڙF�w��mu�-�n������*��;*�Ǯ�����-�`����;,oX��y�*s�r�#P� C����X�N���9��I�fm����1�y����k�qI����6�����4Ŝݓ���}7��U�IZ��sm��j���י��Vɀ�����4Ū�9E���inr�=�	�nuM,���U�����N&���m:���nsW�̵܆us��rq'm���C�U<ɝ��W`�5��}U���H^���/z�9D�C���5	��>����n2�4�9k
�H�{�)�'oD[�T
������7���|t���[Bj�#��S��6ir����а\B����l�J�Z��9���;���|� �p�gn<��9�fP�zM�{{+�lD7{��Ѐ	ϊ�,�Bt4��<�퓎�\Y�F
�M�]9��`�֫O>�j���dte�\�fvYP�3H8���)��݈&����]��*@X��a��ܥ��ծ	UHھ�b�7��r��ck*�"������[�֊���iڽ/#oo��UԞ�+�iC.�#�����1XT]�����;^�m���;��~�s�+C�&���jz������1i����Q�r}�}W&40�&(��m�v�1WWu�yR�Cϸ��4��.j��Jv���35�T�gk��3����\��kݱ�����q���wҪdمbr]K{n��{ɉ�8^��z���(4��u(C�Gyp�zc���E�x�����zF��P�S�о���1l�@��YO
�ve��y���v\=Y�hu�����J�J�^�g(˘�>}�c��f6��#ث���=�������4�,�h�V��Ê���Fe��![��ھ�y���k-����� �%a�Y��hͨ���W��'���2�O#���<�V*A��wWZË&��X���͇pkv��醖�+T9���WN���9n��
���}�:�ɤ�;+�If�`�+h�3<k:�G�;4��R�Q��ہLT�F�-}v��W���������a��+�ˋ������b��+s��75��"0������q��d���֢����4�
P��WBC����}�+��s1PŢh�5շ6b�N��f���$1i��2,̬�c�����[CuJXu��\*JƠ�e�̼�N��OS�х7�eu�!N�a���x���{�ؔ4R�t9�
����9�)Ew`���)f�-y���T,N��ѕ�V��a"䋉�r�n�Lf�$���N��u2d��T���Sw.�܇��Lg��N�$��:����Ȓ�:C�5��:��#[��W��kh�*n��Ӳ�|�#40S/׸1U�y�l�'ѻ
��ie`֪ɇc�!�o����3z-r�R#�с�ݾY4�	*�l����5�U�)�^�EhY4.F���t��e�P����+�ۧ�%��,�"p5��[\�p�.�ӭ�[�fA/eAbD뉤�|o6��X��K��f��):i&d̦ki����{� Vĳu�ʾ[aT釠��)�U��M�>��` �*T����*��YGCGx]-��1���r�i7�-�@���b���WqQ���b=��wd��laC�a���lG�16%���zn������m.��9]m�p�kq5��±޵}��b�T\\Q��쌠�mk�Pd�na4R�)�§{�.��C�M�P�s��/Q��K畵���]����[B���V�u�AC�wv�٢C�2� ti�@�j2��1^��4W5k�ڢr9Knė�Fh����L�jڹ�GL5��}���ٜo�D9�L�UV�jyA��=Sv0�x[��S(f�,��&#�+��yN����R���2����z8�m�D��6zm��R�;,'�L���7R���rYR�@�u�s{/2����0C��p����v��<�-G{@�,Ζ�X�'4(�q[Z��W{ƴ�/x�ի�D�kQ�Ρ�P#3]M4;j�إwY�AVqN�e
�y�:�sN���*[�{�mA4+wq��J�c�]�Q����-	W����LG%\o�����wۘ6���ͽ��#�I��Q�ûZ�j��p�+)��R�A9ڏiub�u���*ܫ#@�}��.�0$M|6�wd�3�f��&ܭ�/�<�t��$k�Ak������qT�kD:�ւ9nٽ[j��Um�(�����f����>�S�B�I�l60�����:�sy��J�Υv� �3���Ǜմ�1n�;Ա��8 �S/����v�"��#͜�S�8���N�j����Dv-bMˌeX��t�7��J����-7S�[��d���*��(���&T�t��7j�f�tG�+�:�R��+�5�P�p����p]��mC3�v�;�v���y��UHȁ,U[R�}H�������m=����e
��X����*��ܽ	-}Ӗ���M�Wf��V�Bo
斡���*畣o���NF�i[!����uh��w-KOw(,�%Fz�Ei���e���Փo
�^��3�:+wu<�yH+�bʀ�҂�<=t���t�ś`�LnĊ55+�01YUgw��m��Q%Ht��.,,�Z��8EՀQq̧�g]�F���H�K����*jN�7m��d;#�,�mS\����ټ��ƀ���c�C�WBw�ٷ�1��t��d.�^by��Ue���="����h+��<��n315��A�n:#��T�ّ���f��Ѽ�I���RE�"�XЮ��ɂJ�e��Y*�<�Q��a��J���;6�H$��IJ�]V��
������\OM��r�l�f�ɽK�5ݕ8�ew>f���j E� �B�R��ܫ�-v�!�mi9�o	���U�U�)e'X9%(b,�.O���kR};u�Gj���/xd�H|+�q�[��6Ɋ�1]5f��k���^��M3hP�c�����]�X����lK)CO���6����>t�eˢf8ƻ;D#xJ�������2�)��Φ���7%�uռ�MF��9ż�o+e&�������U�BUw6=�u�w	�W:@V��w��JM1m��n�]b��]n<�J�;z�iLf\\�hpl4�9�]��ʻ��JIWG�����d6r�6vQ��ס�dJ�K�(Jj0ħ"�eG��b'�ۜ��,dz�����9\�IoP0�z�p9����ɽ�=��`��n�Ce+�sl�WY+v�������N��z�B{u�N#�%J[�;؆megW���8�â���uIg�+;�%}��C�������H�Ȅ��\�.�IU65Ŧ�lN�=o�JfU�|���+`�s��	.��j�W�R����$G��K#��"�N������<�9��Ҩm�9��`�|�5¤ow ��g+]���֘1�f�	ہlHm�gfq�]�f>�_z�w�Ί����{��@Z�F��rٵ�r �Q��ۛ'W\W��뇉�m+��ȧd�B?�`�6�A�w'A��Mo��-�{_)q*�:��Ov��U���<�hټm�h���[�PȌө}�rȩ��e��ó2�h��^��̽�ч0����*�S�u��	�d�v[�qZp��Q����$+/se�s͙wj�0�)/F� @6��Ás�NJ+Z�q|�@�ٵ%lB��\ͭKK��8"8v�
Mظ2�lۍ��(�?v65Ͱ���Ez�mt�0q���̕�c�L\S�o�H�S:��DS�\���S/��%����Y���)F�.s�i˰[�yIȆ+X��8.�ښ�n�Yy�q�-wq+Xp��axj�	�n���ڥr��MsR7�d�̍��xC�״F�z]�F��s�ym��F��'2WY�M;O�����sFh�ꁪ��=���A�o�H�{(P=v:dV���ܖ7J���ɐ&�� NI�_L����������������E."�N��r��rv�N��]�m��[���S�	��5%�擕z����I$�I$�I��އe乹�c2��zjs9E���#X�������X��dP*�h�t:[f	1�v��k.�i��5v9�#�~�~�s���/�z1��i����(\���+9��* ������ W�C��QQ���UP=���O�G��A�}�L'��{{�%M/E�S��R���VFt��<;.���\�[���yb��m�^Q��	
��Y��e���33��%l���a�ŗ'Bj�c��G�]uK�������0��G5#�yY�s��"��"�}/V������kp�7�Ϛ(��y�A�	�+��Э}�֐���.���INjSE֎���6)-�.�������Jdͬq=r�30�٦�*b���X��Yr��vΰ�^B�����q	�6�ڕz����W��0e���!R�}�Έ��������f���,��uH�0������6�AlJ��ikvpu�D,�^Zd>��Fr}:�2n�
8Z��\�S��PEq�Iӽ�����FѤ�gS���=�)���˒
����+�iJ���u5h�m�QCȘ�q�8��D��[\���|#� ou� �P[5���.�-�r�N�M� $�I$�J�I$�T�I%����t��a\��XM�EL��9�n����0�{�䊴vl���,�V��+ԲӇhثR������ڑ�tF�V͛����/*Ʀp�$��:��!g{�Z�s�P����&P�/0dxNWZe���2�����;m{�D]+*q��l02�9�٫"{��)w��Q`�5y�M��P��L�B 깚{8�wGeG�n�Ѷ/*=d����=w�Ȣ��3�Q��O#�>E�b�^�6,?��)ٟm�j�	Le�:��2� �[��_ZF|Ԗ�^��k�F�4؛A��M�EΫL�p�9F�k��,�[r�qv�̨D�Zʦ�;�D�e��ɤt��>Z�2��<�Y(r%e����pX��:��X�Ǵ�:�ݝ5���H<h3lb��*t酼-�xQ��+B/:��M�w�W1�QѹbW,�WFB�CZ�xSw�t)����!F�T�I$r�32I&�$� �I"�	$�Sǜk��7�K
��Ӹ�]�%:C��I$�'��J�IԨ�Z�h�vE��s�
��m��$�@����{ՙ�q^@��	q�u��N^�J��u
�;�Ds"\5b7���E�H}��c0�}ᕼ��뾖�r�FT�&.���(�H�xiǷQ�Е����wV����A"{�B��33&A[cL��e �<���ޗ�������s9Y�eDV�ڻ��n���/4[䲲uݗZ��4C�n+K)��v�NX��yʋ���9��m��nu�W���s
�fjd���
����K�D� l۴��wd���ݳ�8�
T2X��v��qR�c��o:k&�[)@Ś�
Q�HH��)iR��v�v�.��tB;-Y�l�Z3v�ҭ���xι��*��]�CHY/I������B�el/*̓��I'I�I� .I$�I�I'I&�$�'�����q=v�畕����ɤr��!�fj�r��5�ԩŁ��:�Ff˝��6�Q�c7dT���Wt��b�X���c��QD��EkF),���gc��^����ڈKɭ��Qǵ �5\�F�1[����v�X�:�4���R�ni+u���P%R+��b;+��ݎ	9X�:�#��B��O-�*�a�C*��(68s�.�n���*f�тI8���fﳒ�6���ma�vH��Gǅfn��cF吟P��K}+����z�����'J1��!9�JN�+!�e�n���8+y3��*kOx��"�<�P�:;�j��XNCt�\�N1T��w�ܜ��IH^��,Q��i��J�Z�Mej��H���J	����iF%��䴮���	�F�l:J��dj�"`�>\��D�p�!�d�M�I�A3�$�E �I$R	$�A���h�I8��|�8+&�)��U��%�)W�:��.��p*"t�
ˡB�cf�o�K�HG��A��ȭ�ur�q�H�}�TB�1���X�����z1�b�[���ɛ�q�#�[��,h��^U!�s�w�۽���$\y�㳢�3�/zt���Z��%m1k*�'υ݌-:��Ҷ��m1%�J���c�s67p�pA�N��f�l`�7�����j�jۢŬ��Z�e,˲ky����̉�ڊ��w��aGuh�x�ym9��N�@��GZ�}z6���Pv	�r�WuI�zc��m+������2QɇmM��w�Q��a��1l��9��[dGY�d�����,�`�H�%,+���9�4AzB\[M�wn�$���u���2n8w���N��PhV�WMu��YE'�й�۔��҅�D蓻0j#��Q�/�հ��DP�U��r�ۥ\�r���e�[h'�-��2�,�W�݃ܲ��g�;-��@�yE����27��l�2�-1c����nX�1�q-�A��앖G?�����n�ֳ��켄M�X�:�U���7��;�֡�d�^o�ō��+f���be*���E˩ټa]��V����eR�aGu�96���`���sY(6.)�K�L�y��������w_0oN�u�=�T]/Ds��v�W
��jF7�C���-���Z�joE*җ�k�UҶ����{�Q�]�uJ-�'�U��K�zb�8[����6�J�!e�&p�i��ٔ���W��B�*�N��Y�*�S��n��]m]��R�[�LMvA|Ѩ��爼����Q[;�w�L[	�ʬ0.�D�\�܈�"DhQ���>qJ�0���!���;�^ +�5,�[9�~����
�IY�	b��.�7����#��XQ-�C憭�h�gr_=R�!�S>�vڗ��w�`�f0�jNI*]�h�@��[�ۙ�t`�y�lE�y���uC��5#5fo"���pQ��t��:|
0��9�v������ܥ�+#s{��i�����!�=	����6	�}�$.V�.�$0Se`c/�;A��<�T]�{�Szڬ�t�mՉzΧ�������c�./�.�V�ϠS��,8��c����(�J
�{�G�]%��S��i���=�K��m��5|��e�c�t	wn�7!�������v��JYA7�¡0�XE)�Xͩ��)�Ċ�� �kSu��&���d�ɳ��";v���͒hv�ƕ�R]���lv+Ⴄ��ĭ�x"�q�v��veu=	��vBx�ze)�p�ri���eΖ)�_
Y2���DC��PC�y(a�}>@�R�ǃ2�k�l���%��h��s�{e��;�H�-���
K3�SE>��y.;���X� �wv�x�X)�rZ��ݓE����c��Y1��VvA�s��]���KJ2#h�]כ�G-=�O�G�T۫��hQ-�9J��}܅s��,&� �2��=-�E���ۖJ]�x ꒀ�k>ҳ7r�ʹ@�y{�V����}�����Z�Y��e�fv��g!�{�k�jx̝��um�gtk{J�nD��z�Z�7G*���n���ҭ���h+mm�iGd��E�3 �(b\��d�ŋ9�A�%̏6J/u]��5�>��{�Whӆ��8��Bmf���:��̣qm����qf�xݫ��d�A/'1\N���4��k�&Ec���ɻIԼ{��d��Q�m0"Ŋ>�9{��'4���y=ݮH��|Pt��Ψ�y�YR����Z�k�Ӷ^���<���SV;��>��r��Ȍ�e�Ԍv�Z�[zI��ѕ�i�I���+L{X�W�e1�a���G�U����|�҇s�˲4�Z��Z�
rnSR=��%���yrI+Z��:'t6�}&��B�Bɯ^�ѫ�];`V�i���镇�Գr��`���ž�5�J�eX5�D�.�(�"�:W]o���ݻ��n�;�Ӈ�|��=R���>˘���؄ϴf_ (�㹸j^ŷ��=����*���oZ&+$Gǭ�����\\mv��כ��\��I��Π�ҭv�'���ϬrJ���}gpWQ�x��v2ov�c8��I�3�i,��*��a=z��@�7%��&��Ճ{�>�}�19�R��L͡l����]��'&KE�
����ĄZi^�y�Ҿ�AiaS8
�cQ�pK��U���vS��)L����̣/�!���z2��r�,�ᙪ��SZ�*f�5�M��δ�=���B��ʏ�wi\�n�DJiT��t�V���q��r�';���}�؈�:A�ް9V^涉h=νa�y؂�g�.{s��+�DV�+;l�۲9с�V�z�Ń/��,�ZM^B��Bf��ay�׌a�s����R:&�{3v��$��Z�n�v�|�A@F���^�Z�2�0�l�rs�c�:�w��{Ck����$qϹ^D�2;��Enᖴ ��A�4څ�A-���&m-%ʛ}�a��ܬ�zH)3rw D)M2`z��%�E��W�5�q{1B|����|p$�n�C���v�J�j�E��bc���a��U|~����*c���N~s�8��}����K�jߞў�&��p��zI���rs�tߧ��?Qߡ��f��x�z���l�3r�����Zc���Q���ȋ}k��٥�����!�kAL��o.�I�n`�`s�nK�X���v���z��|��Wa��b�����2�q�oAëp;j<�laJ�ܻ�%A�X��"�5M"��sz<��J�����=�=N9Vy#�5����-�va�z��3���h�%K��&xpU�����R�]ܖ���W����6k@�o*nu��`��8I�cz��+�YOP&Q�)Yo �p�ƹ������F�33"�l	��XV�ʸ�Xyۛ&N�g��2�b�1�_�*ř��.�j��9�h#�X�L�yk���t*L\-��y���˸��v��m�J��ޚR�R��B	 $�,�yxjȼ�͉3�+9��B�m��wqt8WW��ӷ��$G��=�D���% �<xD�Duq�35QZD�#$M�r�1Y��?;ﾃƳ���Z�md�䄦L���K�b��W{����²���"ĈU�yJ*�Z�����U�7�����啤�, �dbXI�)�3�
��F�����L��4S�)���B�Q�͈�͞gf6�)(n~:�Yv3��B�5̖�Ɍ��<J���9��6w�;���"أg+mm��-k��k>�;ۏ�ŕ�S�Ս38m��*�J�ۄ/(vUԍq�M��$��#X�H���m!&QjK�\%�����̢=��@����*I*�y���p��P���u���@���������ڻ�l+��s^A�,&�q��n8�r]}[\.7:q_ߪ��}�gvU�	|bz�!s�t�.�����йC��a{es�A�Q$H�Mҽ��N(ҋ�Z�ũh���@�&{6ca�ii)�̱7��]�vBu���&v؇]�0�*��������B�7��~� ���p8�+#x7Y��T���(�:��x�Xz�V��\5JٜSt������i��]��\\pdޅ$�@�ݑiű7�� �3�o\��Z9U�B�oF+�X��ǙQ�㓸�f+Q�b�}���z��Z�B�利��Jy�H�%�dX�Ӱ)�Nَ�Zɝ�!]���ՙ�l]SV�>�}��\U���gg}�,�e�֦�9��Pq����.I��@JUG�9��l�ky���=i��(;����;w<R�Z:Djo�����z,��F�蝌�`q1}aζj���3}��&�u?�7��A����ȐvBtc�ܣ��k�;��զ���3>�V��n�w�>��9<�����ݷ�3)E�L�vaAe�7�v/F�݋&t�9�<u�.茜qƅ�-��r��bD�Sz��]�~{��4�m.���&f�4O\����X��)�G�4k4<lZ�8թ��~�wt;xi�y���;�uN3fh�s,A9� �3s��7],���]]���vL�Y��lg�����<|9}2h���d��I 9�F���r���ɟ>Dtݑ3\���4os�.嵽\"\ \-a)H�yڸ�x�e�>s�k�����͙\ګw�w6��
�;~�)�B����Ky��S��E��Or^q�=��cx�U,K4ӫ��"�8�-.s5�L4��ȑ��Pg��y�-�ո ��
�ŝ�.�J9o�
�������9'�����rJ���H�q��a�'���ʄA�,������(/]��V����R� 4�i�F��qak�1�}Km�Ӏ�K��ь]�OvS��է"�;�r�Ć��S�q�YP���y�@t&S���m/}�:/ �V�v��-�R�;�����7�'���*�Z�2�q��GnB�\QU��q-"h���+:����^��w�fSq��޾�3��Ѥ��"���E���_8�H��o�s�δ�Z�ToOAT�̀�5�*���h�ۍ�Q؝��QB��-ɵ�W��I�Oz�&���xX�u�㭙J�׀�Gܣ��+���^�8�lsW?18,«��v���L�� ��k����Gְ$�f]��j�]�re:�po��,8 ��/FE�B���VsP�M���Y�����ۈ$�Ĺ�]�|�����e��E�k ��cլg��&��0�,Fs����yy�����	CO�[Y�\��2�̘����)�x������o"�Pb��o�j��R�zfp�l�7@2)S�u���B:auۭ��q�����erE7�jIYs�*
'��E������s�+��,!�)9��;�<�S�:y��z�@ڜ�Ci�ZN��m���q:�p�T՚ ��}�<�k���t�}�jwP�9�cp�W��^9�zL�;e�B���Ԥa���䝾�X=u�Z�N�]�*w�=��O�/J��M�L>SP�4\�c�H{���K�kc���z������ �s�Or�:ʼW"��b�-�3����;��u�VTG��ل��mL26�A�[/,p��^�c�+>�9d���Vn4Mhw}��X��+!��P��Ցݫ-BVJ!n5�g+�����ۧ<5G![w�c�;�w� ���
�Q�,�L�����S��Q��drkxx��}]�.�K�|��W���7kQ�)�Do]�����y�IH���7d�W�Y����as.-Ĭ}�Aj�W+�A��e]�걋�Q�	qy���k3���
2c�SG32���?z�OV�S�죧�VA�aJ����~����^�\��{=�gh��v���2���eL]��Zٺ�1<SZR݊���~�[v�7&ۊװ��1Z8�����V�/^p�:gw������+ ��HOm-�V��Ȅiv�^�������iۣ��Ŧ�|a��l
1� �����$U���L�{uL�:�1���ə��vv8V��kVTq`5��,�3v�"iZ�ӫK�L�n�m�sBd�-Ɉn���og�|U���[X�O-��'u�����]*׹ሕY=q ��̠!�2�c%��3b��;q0�⃰r�q:ujj�|l����/�k��pds��6�F�@�m��[�	,��}�U{��.�0ڭ��#��I����v�+Ρv6�CI�v3;� ���Z�+��G�Ϋ�r��XJ]�Q���iVh���<�4��7~�A�$���q�Zz�@��^R��!��lG|s���댬�u!�"gR ���,�"krxͱw<��9VR��Ml�U-ߧ�r(@���$j'���x�� X�>�d鼼��P�Vu�z���5ҰYë����.,ʀk�4�%�9MƌR=qrĞˠe�����h���`�7"��L�Ԝ��=p[��l�]�4]�60Z ��lOl�ь]ķ�%�n�3�zξNS;v�f�K��9�V;��"fxĭ�z��>�E�)�dQX��b5V[�RUVY��k��ϡ̠�RhQV��,�A�v37�+�ޚl
[m�a�B��x�XQ����:�\9���1�e�b&��qyvcR�	.3�n_�yl[t�@�3Q�x��E ����ӓ��)�?V�d&�FȠ��g���ɥ��V^a��,��s���-���܇u;�j�9�c&a�"D��t�{���-G3"��{˙vd�Y�=g�nC4�|&l#ju���B�v����u�������{a�w�"(f+��eR�|i��Ȯ7�M�Rvp���-R\Û��oo0��3p�{�cH��oem�ʍ��.�����9�&�{��@H���Z��CQ�N۪��mU���5szp7��S��s5m9���p�S�:m��h��E��fw����γ��J��t\7w�-e�vI�j����La":d��]��"�����v����J:a��4�˕0�G�'z�@��L�gFl�2�}��N#r�ѫN�>C�ڝ��;,�8WSy�zR�c�l�g�������'\ܙV�(v���lE�k[x�3��w�o�5�q�Z^H�h��n%�Gԍ��/U<�#(.k�i�n����XZN�QP�f����|��o��E�����k��7[�
J�;86H�{�®۷�T���9�)0ו\e�T�dXF�y��ֹ������n������T�[å����#Cd��{Y��3�
D���EӀ"����ɽNq��.Fz9U�B�i�ڥ�v*Ʈe���Ĉ�3Z�1����L�ש����(H3[����N�k>��&1M�ń�X�9���������39��c��T ����~
C�\W�_����p+v�)�me.�fu�n��ضS��;j�˦�Js������f]���l�G.l	`�}r�Ͳ�����g+�窡����Vk��=����Sc�C4dO���CN�"�N�`��¯�� �53{�LF����K�Ɍ�j���w�r��n��$��ɷ��uE4ܡ���<a7to�"w>�Iw�gϫ��y���j*j>���G�v=��+n��f>��v�b���&B�,h&�WEܔ��FNYq�d)m���Kf�ށ�;/A�J9�� n^pyE�d+��b}7����vP��{D�ak��7}A#Ů�խ��܈�R�9s��ji����4q�)f�|`Y��Ё�j`��R��9�L�l��<q���T���-�馮�/oKD���hM���S��t�R�i�at�60���YX��������̜�mݗ���d�R����J�m�ۺ<m����h�$��E��x�ڰ�6�%w-�]9j�����h���.I�����׸��W�wJ�g��o��
Lŵ���K�����ǃm9"�^��JLdRjuO��;�j�͡"� ��j�Pɜ?�qc�jFR*0�nK�bUe<��_T���mM"����6DG���]Z�4�D�Kr��},Ûw��I��-9� y�zІ���-VX\�}�]��5%m8]���K%1�z�w" spd]jecֻ4�!�x�3�,�8<u��c�Õպ��!+U�է���4�u)�앴鞒��*b�U<y�l1u�!�>o0ӑU;��Q�V�ڠm0��K��Jںp X�#���$t���
��\�|p��]�)�ªƜ�L:yc14�]����W�%5���P3��Y.������K��]H���wG/kyEl̸�V݂ʕ��[N	�̡g11u{Y��|?�U�!u �$$��ix�T/&��/��1q)x�]=�߿}�lo�hWm�pF��� ��Ԍ�v'\2sR�}�0���<������$�:��V]����l�p�2�8�<�	�� �Ëi���������hT�)6��5ĵ�$ܞ&�!K2
}�]Ht��P�%���F��3L�)M��Ñ�̨�6�q�9L�]�'+�uRIIrQ�A+[)"�QT*�E��5�	�'�PRx�]a�"��MgCƁD�{�����sFs��q�[�6�#Lĥg�8���4��E ��+��nlH���z��v�25����<�$So�~,��-�æ~�ګ�r�z|�����a�G�n_L*�R�Tn�frIt��R;�\|��]��.���7dQ'��~��*z��x{$id9v��>^ݷ���sg���j������,����T�'�ǽ�s��Oaxk�ƚ[M�����q��OǢ�T_�Vo����Ԯ��}�TB$yN묤���3��f����z�;�ܻ���c���Ž{����S�x��+חx�i?z�����x&�+#�����ۗ�Cï.�,5|7������dŰV\����v�bo���-$Rqn&��x#�ۿ���^�n��z��=�����m899o5���)��[�~��`P��>�x�R�G}�f��S�*x)W-���D�繇'�S�㻡�M��ǣ{��ÞQc�5�v52#l2�r�73o��B�یA+�;�RRq7;�nVｽϻ�P�*�}¥�{Z�9��x.>�*4T�#$�b�}#%�ըP Ud��(��v�K�y���o������۸���gTt�sW����9�q��Z�bs��E����~#�E�;^��>-^���!oB���4n��͡K�Ⱥ���:o�-yg����_��ڀ�T�c�����^��u5zA��h���_/1vz�j����X�ue`�s�m*��]�Uf�ʂ*/-ʨ	\��sQA����U<����I�`���)�~O@i9�8)�i�=�������~���K�w��5ٺ�L��vƲAki>`Ǜuw��q�$|,��Dr�����ILi���b1��ἅ5*^e�ۜ=�KQ�����,���0�/\(ڈ�5�4 �уXg����:A�l��u�Y���g׍\n�nܓr�����
���˸y=}.���߳��q�g���� �.�{�2&���_\�GF�H�{kX����L�^�|�j1[+b0����MF�ϫon��p�q\���7[�Ȃ��g+�&��iuN&	���q����*�F�/v��>��O_��{ Wϓ��pq���gy��kݝ���r{I���=�Q��VԽ5Q>ϭEXc_��
+`�y)Ph���>I�g�'#��{La��k��Q�Mԧ����ܦS�� �e��2����˃��k݊
�ّ��ǌk���_c���@~����z�aBP�r�f��6A�֭���5��J�\s2e(S���Ĥ�%`�y>��������С1 ���J�A��Cٻ`o�Mg�5h��W�Y�{���/>(��;��;����β���u�� �{ۻ�ׁ�>qcܥbU��G�+��ǅ�N�2�*v&�q^��W�Qf��̥O0�j��ϢFLeہ;�Fs��9��[>W2 t��"�s����a�3�#Y@%����]�i{|���4kZ��,���/�u�z��[���O5W�λ帆��S1B@�D����v!�&�������)�RԴWY�{�Rny�{��1�ֱ��pSȖ���;�y�zb��`\�/ba؉�� �5P�i�v�pA����a�]�{��Q��	ڤ�W1�hM�oF�CN�76yB�p;/Ѩ��@n��^E�B�u�3Y��^;'���5�^U~\� �Hܤ�{Y��9V0��Ks/�`*n<���C��x+Q\<�Ú��n_z컹Wr8�a���x�P�&8��;V	��}3DE-����l�y=j�R�;��P��Z�C�v7�	�`y�M@1�\������Ӹ^+x���,�T�3��۫_��8j."�T�����!sT;�D|���d*��	�Kb��M���q	>R9�ș�o�w���g;���D�5S�=��Q�/b�]�y1k�Rإ�D�S�Z!�RH r����A�!�c���s�����Ѩ6���;��K���pu��^O"�."��;�uA�� �)D,U���_ݭ�{<����3�WE9:��^¢��/ d��]��935�b#�5dŹm�թ�0U,�j&���<�{���xu��!Ҩ�1���/�xZ�qu�(7���KC]E�s�;�sE��I9}y�ܒj�w�ռ���fz���E9�B�!j(\A�;PC��^�"�I�/`_'"63\���-Hr�E�{s5�o�3��.a�^��3�oe*l��Oh��G����RvTq���`8� nf[R���1W3�[�|���">@3q�F���"���yaL�Pj/aQjȺ�Dw�Nʈ�)'�Kc�3���u��0zj�7iF�<�_������Jn"��*Pj�Z�Aq5��!��5q{z<��S�y����
ׯX�n�?�X:{t�t~�M���8!E)y���wsY�t�d7��C��܈����b"ǏZ��фp���i9�Q=dL7ֺo[���xT����}�`H!"-c9��7�N)I5��!��5KȮ#QQ$�7�7ڦ�]A���� �(d_R�\ԙ�q~ߘ�.`��P9�^6�E
��Z!�+�Z�D�D���pL�/�C�[�$����;{k��9�Z�y�w���M�y;�G@�����<�X�":�؅�h���!ȖsC�P�(��D�^B�n�&��Mk�_|�w�Iv�u���x�b7�D;T���R�Z�!�.���R�M\����/�T�9�U�����g��1�g���]<��TSp/1q/ �^��.)|R�.�c��gb��;��F�j_��@�S~LbKb��w<�w~�fuIh-�\�������vy�<�y ה<� /�CʧP�T/�T�y��ߕ��|����@��J�b)�|�sp3F�Ch�^�D|;Z�b'b�S�x�y����6��o�/�s�[�X���jpq����P50yC����Tq;��WQ1E��#�R�L���]DU������͛Ǚ��x޺t/
��=�h���]��m<mC���D9Q;q<�n/`st�4	��b��+��5�k8��ƻΝD�f�"�,�1Bf&�*�Ej�{���{Rv.b��)Ƚ�@��)���.�����u���^7���֚�QX�P��2}�Xd�$p`���l�\�v|V�k�?>��>񽋓O3�,Z�]cKz�q���7$'x���YK��}�Q�����uw��)��ַ��tLA}�r��s��+�jԩ|S�pd�H�	"��:�Pj7�"�^	 r؛���nڱ������MNL�w���{/�G1�[�3T�@l��:�P�D�/a�)�Z���+��\�oi��W��/~���]����y�B�;jC�[�Pۥ�;���h�3A�.�j���Y��������g��Zc7�3ٱmp�LU(s�SL�ȯ'`TT��w�iDs��ê�j�BDu[ݹ�xǕmc��nE�!ڤ{н�D-�&ཁ�������v��W*"j$��&�R��g��ֻ<�<�X�;͝@�چ�P^E�|��v�<�n=��PZy�E;ϕ�-F�X7O�C�M�3W㊚�|���Đ<��)"^/^���%��e��o��d^�D<-@����Jn)k�vv!hr�ȁ g�o����c����ռV��Ѩ�n���TK��$NŶ�`E���ה�#�G1R^+y�y�T�Q�v�7�������/9��\�+��)x-�y��w -�u�K��yq|"��^n�Ew�R�.�Ȏ�""v������l��y��pJ�������@b`��&(C�-�P�q��j����ɘ-���x;��;��̱��ձZ�B�PZ#����]��LV���e�|��]v�qޭ5������.*�=йDn4��/d��[�1S��}Q��W�������-�Q�d	kk��:u�$�w�"���3�[ߖ9��#���}Q�^\�<���B��P�NE���R�;̒�f��w����z���CQd �nYO!�$�b�;Hf+k��ȡ)ME�*Ds�3�7 7P�^�H�'��o��n�s{����t���\�����@}@���j�3�;��7�D�^E��D�w�2g��|�;��ɨ��w���6<��{3�ҥ���D�<�	��^�p��<�
jZ�����C������{[��n����j9�nhj"w4&":���.wC ���^ʖ��j�j�+����Ǜֹ;���w8��j�ȼ�_�E�]�@Ú�<���.yd9��Ñn�D
ͬ�@l����n�e�V/[��/��;��.�DWQ3�A��yq{�) ��3�!�&#v�����s@w���(j�z���O<���l��]RȄ����/a�P'#k�rTWp�ئ1�<��j&P�9��@/�\��_7��w�;�s{����E��T�����\Z������w��b���y�:��%�@r�|����{�s��1E<�u����)�-��j~�00b��l���j�U3�W��;&�Jn�B����k��@7���u:���9�%����qY�w�Jyjm"1�;O��L\���r��6��sWƷ��{��Y $EP毐K��;� g�.:6M���Y�U�Oi�6E~:�][tiS�����'=U���	�Ҿ�#;/-j5ʡ�3�p�ٽ�lU�e5�jr��Q{z�Fb�~��ϝ:���Eq|}K�{�E=�Z*G=Z9U����፴�5�F�`9��1�j8�>ە�nʒ'��I`��G1A]]lr���h�I�ɹW�&U K�Iq����kc'	��)J�pNi*NÛ(����Y޼*�;_����p��F/z�@6r)��oNQ���FH�k�G���n�(n]r��0u���e�L0�m9���$�4�z,�Pe��;�j,���r ����
Wm,J�S��E`nu��֔�D��Ó��������긌�+�_��޸�����C���qk�^x�5r����)�즍@���eA������v�,��sk0�~��*U��[Ţ��]�����S���sg9D��q��l����������}vr-˛�(�/x۩Ʉ�������zp���2��/.7�frN~T �X+A0�ݺ�$���76[5l��]��7k�]*�Xa+vg-2r��nm��#1;�݇{@�I�#��r��ZuT��T���y�Hf�������q�_��̟�+���'���航�4���l��0��4)�ʈ�8!����ʛ]as��l|u��i�]'���L6�-�fal�b��A�p$b���	���મ����7z�m�u�ٺ���߬��A�u�,[�C���=�Pln��@�Ct�?Z�c<�ٹ��S^�n��䱞AB��S��.]*�����Q�B�4���%L�@���'��;#;k��o�Y՚�z��R��vB�ZT�F.�aG{(mn��q۶H�ݼ����%�ĴX��"���>��̥V8^��42Aʏ1#���k�^��!�@��͍�Y;{�զ$�ܕ(=Ρ�'1t�+);�	'N�Z�m���Y!̣�J��P�S��uS\ڤN�̰���]�b*a[�TG*��<(vڎZur��������ڭ�b�Nw2��8
�*��q�(i���ۃ�e�uk$�X��NhW�3aTA����6c4���XS5�-���m���6���pX��F�d:�9��w��EC�=�ʤ��E��.�A������|&?�E��N���^��o�LL�tB�2�=T��Nd&�dѐ�WR١üV,+b;8Zf=�"��f2t����N��'WAq��L�����;*�ʐ�^��B�7� .,���rBڽͳ��'Z��.�iN�eeJ���H��^�,�y��/�v�繓�S�F�Nz���Y���7`�@����ϋ���m9�*^߬@b��2wE`��C�6]
��=�;KNP�+��	�c:��O`LV�y���4��u�՜��WE�ՙ�n�}���!:���+p7ǎwu�®VH�*�m���Z�F'U��x�u�@D�"��a.܁�؟D�r�^r��Q{5�ʛ]%�w��2\a�@��)S�ɛ����])����gU��+��q��q�l3{�-"�Y���Ѹ���Ue�u���� ¹�9��i'����~�n��p �+:��g��.&KUma�dEj2M�����ɓ9pK�t,R9ۍQ3k�CS0�r�X���(�������&�_S��&������qAx�+0�!k��]߾����EB�/��n���)#05�Ғ��7�}��2�~�Z�j҃���*9��:阴�,٥M�k��m��f�M\�f3�R�D�#�ʶ��Dwl����i���t�rUH��l��!T�p�tm
Z�˰"5�H�9�Z	�S	�⦹i��hʪ�$���g��l����j���E݄������rp�b䨶�ޓ��S,���nd�Fl�ƈ�0��%\tk������N�����CGz'��vN�<�*��P�u��qgV����������纯`�����"�1��\�5og��9߷��w���A�9��|lU����<��>N7�7�����s]2x�� Y�y�������?�Cn��:]��c�fg:CjJ��ҙ�>Ǧ'��;U��|�din��s�B3q���s���F/��"JgK��{�lJ�x�OOq��1k�f�,f<g>}P�5���B�\[~���}C���� ���^�M[�M_f��p(�1N��a"��U��=]��q=�KE(9�.�:�5��ma�M@������UY-��l<�hu{�z����o@����Nϯ�TQ�����pp���;��A�<i��f��'�r|cjqz+�h�;��]ڭ]�[Zh�]�I߁�m��b,ym��mLc;7�|�5����A�FEBEP9o3���y�{l�\�m�L�`��"�-��T;}��؇�`�Bj�;$��Nl Q����:�΋c!v ���1�PE*^�z�������Nc�x��O�T�z��!�.�=�$�m��*2i�{;yVFA�{�*��X/)*y�+b���DT#Q|���V�FTk�5Ou��7=���{�=1��f*�P�}�9<��G0��(�V��ʷ0�Z=�λ(���Y~)w@ќ�.�J��zw{ŭe%�[�i���Ύ(��-��_jNɫ�V_f�����;E_CC�ͷ�P����S�\�^�`{�^��5�}�j�������7�U�Bf`�2G{��3e�R�[���̳�Þ9,����;	IdQw�5��*z�<�Cw'���W'u�T�MْxU�n����[q��r���Ěrm���@���-��7[�� 88ٻPucf|+q~���\n�=�<�G����Jw�&�o����w�:�r6�f��pY�g�����f�@��&�9���['�BNB��g��)U�yL&E�}��P�Xr[�{�k��e�F���[˝��Tn[10���Cgob�5�N�)�]�Q��s�����D��r2��o�����*r�D�+_t@�pT�׎�W���j���V�D��7X�I1�0�ӶL�XwtnR��k�ٺ�f=�f��Ȗ�]@Rc���[�f������qMz#�jPǽ� =DYd�D^j��u����Y��a�+ؼ<h�����T<��Rc��wm��R2�X�9��<bׄTMu���9x�)��|7�Qp��v�f��o`'��-�Ӏ�p���V2�Ҟ���x�#���~��uZ�܏��֞d�F�P����;L�	�k�H��*z�2*E�7���9f�Dm���kS��σ[Y�\�ra4��h���Q�1��>Ր��'pDL�h����9�q�m��<�!�%[U��l�B����M�.:ΰj�C�3ш������}�WN���)8 �K�i�.ܟUҝ�%��pQ��L�QU�.�-������퍢����>�
p+&�
?GFv�jJ��ܵ�+:�1�V��>�QEd� N<�Z��L�[w'}ʦ��`C˸�U�PTL68���u��$s׸2s~y����3�BŒQ��ؚ�|�V�pЛ8�b�ӻk�{��%g[��8{�?�^���=s�������I���ҳ��K=��[��ח���)��\�˯��;��dhx�gp�d��2�����f`P6()�Y��|/;Q%�^��Ѕ�.��T|��{,����J���M��l�hXf3>��"`^]J�ٌr+c��t/#=����j���&�
����ū�qU�����Ov�=������I҆�5�d�`�m*�s9��
���:�y�!J���;���N$`��rE��N��̕�o���E�	dD$UG��}%�`���!�7�25.G���i��o��߆��xֻ���b�C���4�\�:�T/�mŵqO��[�9�ٍ�Mn�d&!�U�B����}��@���yAX�s�W��-�8��ql��u)\���$�Y5�[�m˺�/؃>ռ�y��,W1Q��uq����?F��5��	�m�v�߸E;G�a� ��3��\vE�}_^]�C>׮���Km�#�Ӣ�-��H<�^���L\C�m�
� 2���<�������LV��3���c�5˝�*��]�mEZ�^%�(u�S���+y��ٜ6�֬��YT�7Sܶ��гt�H1���e���k��q(�hu�L�~kx�g^lַ�H�� ȢHȫ�|�o�zp��N�� �\n�Z���	ti��[y�<��k�U5��`p}��� и��e�{G�24p�פ�Wj[t���76�]t�n����qmGlv%] =�����44؊�Ö�i���2_=��Ock�f�j�!����oi�����[nM��{��g������U��+��:�|$L�TN1�>��|I:%<4��a�rq���b��l^��w'f��$q� ��L"4v+GI܇��b#��B��3n��i<�E�^0 �|%�VQ׹&�g�Ÿ��M�t��������y���1�tʱ�`ެ���#N��k��PR�jt��{�*�����l�y��ٓ�oJy��BaǛD��E&$�������U�DU7���k���Ʊ�uo[���˼�1�!�3qK�m5H&�Z�V�D8=��3{[(�V��7qg���hh����Q�wd7�y=Xu�TGf���co ��bM^;�M�R�罡�M�Q�O���A\U��,��KF�2�'-f;�|�1�|c�[p8�_]3n.T�,��S�e�XSp��x>1�`"�w���=���\K�鍎9"����qܞ���a%Q�{���ֻ�`��W}'�@Rvd�M�����Y�{��}P?n�� �W��ץߕ]�m�ߤ���$�%�q��q=�W;Kv�:U	�=EK���6�sV��3>{�C|0�6��谫���ܾ�2I�װ��Y����W��"�* �*�s9�}�������S�
�5����b�IvBa��0f����N�� ��s��b&Cα+=7*�f�-��q<��腐������E�(�����uJ`���N�������E��i-��b�_\��q��!��Y���c�"G|Ynn[&���8�7�6�5���;c{���	�n^��f���n6���<������Mv'����\�������(ֹO����N)��o�I�|��~���#�^v��>�B2��8f��I�M��e�
�t�)��s��mOWl�F����5�b�6�j���/�5g����\���Ť��C4<Au䍧��"��/9E+�嗙[�&)5��=ARD@FAw�1����݅�i�ݲo*�$YAM������^�k~���H��X���T#3���w�tE���,>I�μ5R�;�Cc�f�u��=�>�N<��uh�&�\`d���k���8Ӿ�X�`�uF/����n�J\�;�Lq�b��C�n��^V��THڽ�'�� ��X��q�q-Ug�n&�����\�������_��|z*�c]�h�޽���'��P*c���S͊b����{b�s���uС�M\�v���}���U-��P��B]ꙍ���}Uw|`�hs�5�������P,��nkT���齦�>xzBCxoo��R�M��E��L6�n����j�yB��`v���ה:�F��H;����"|[q���R�o�QK]K���1�*�։�\���H,\�/�!�=v����P�w���kW�k�[6�L�u*����l;�^摁���A��4���иlv�h�#����U.-���.{5��o�eo�CXv���l�'|8�i�s;ݵ����zz��];���0���Rk�؜�9U�]��{� S8h��$=jj�Y�vˌ➳�wT�t�ێ��]��Ua�!}��n��jM`Ҕ�a˵�o2EY�*�w�O�q��Y]-й�c�f;����:�Ҫ憖AY�r=�he�=�|�t490(F�d/o(u�ui�::�rN=c-47�%}�����R�ᕢ�w:��|��D�4�,$��2g��L~{�;U�v��̳�T'���Qv���n�2�A�jML���`�֍`�qN��nе��;�s{vS]�`^Ԡ���ص��#��|��r���;�4����IX����%.�����o�9�|��ڍ9[��7��z��+:B�cUɵ�k��j8��&�����Ƶ���K��v�^���A�κ˽��m5xg�D�����9-n�R�̜h'Q՛�1�Le��ϙ�ٓ�퇨m��C��<�Qv̡�@�j�g%W3���VS�`��b����Fb\c����v�|�r��6�]�4�D�]u&��>P��fp��®�]���}���V%��w#7�z�NVN7s�W�6oD��*ѽy3+zo%�@J]��#�c��'<6�q��k��W��[e+�=uy	�!.�"�X��gN:c!��(�-�M,���߿��ъ�I!RI0Lh�9���ci�ksmj���}�}+�D|Q����x����x�W#rX���ގ۷LZ+=��}G���­Y�f-�y:�m�ڹLsq�Uk��ҿJ}�ᘥ�,�d*���G#'�:��V(���}q��~��jj�Qa8M��꽘�fZM(��q�R�˓	%P��l���I��#�E����ʋAa"n���3JL��A@y�iE$k.d�zƙ�vm�B����ĵ�mK�TY�:-d�:�am�T����lv�ӭ��t�"�ÜOw{KB$�Ivظ�3����L�^봱Q	�$AD$�'�'�����\p�V�����5�6��q��J2��ʖ5�n�����m�ַ��y����Y	fc��>����~���6kH�WI-?Z+p�y �Rl�g�k��P���}cWC��&�%��'�q�)��;����Q�Θ�m��S7��� &�U��v5�ڵ��qsuZ�ڣ���<�W?�Mz��0}�f^�r:j��ԯn�Q�*a����¹�3ђS���G3C{��2kL�x���[ lƊ��"�m��O�N[�n��/����1hjcu@�;�����̶&���w���'s`�*e?߽�����ڭ�+��܋o����b�9�ñ�&ɘ,�O�AeYI��4�8�屧�o;�O�D�k+]����s������8r���^o
o��5屣�S�\=����������kߘַ�J��"�$}��G�OK'��6�W�.�|$O�[��Y�.��yfߺ���қ���G�j�����CY*��槶�>�=�_i�c]Y���aP5 ��%cgD�·�/���^����N$�80�F�բ�\�N5¹����^d:c;.���&�dl����NV�����?>�/a����2�LvQĝI�M7������Og�ތ��&ET�^��7�}��C>�΍ALm���w�D=Hˌ����E�>_,u)T�V�/��O7�Y��'#]C|C�Z:��f�:����)��G��&��*����>��R�('H�9�s���V;����+3"����&Ѕ�W�<�ŷ�+�,R�r6��ğ���_�_W�v�ȂH(.�3��{�vc&&��9�ܶ*,9���a�޼���՜���m�5��!\���KS����ʮ�<;YNr��<��t��i�B���������N�wqG�lQF�`�r�"�ӥeD��ȹ3����:��'8�y%ˮ�"k�:փ1�{�ʸ��o��k��g`1�Rt�r.6e��q��]������z����B�oq'ͪ��\<��Y�Umљ0"m���A��B�y�P�;��&���F_���Z�wݒ�s,{+p6�6x6L}�S����4.�9>�ӢṴ�WN�.�F\ط *��B�"���Y�LE�x8�b�4��.�j7Ц2���R��)º�n�2t�@��8�~��ۥ	II �g��7�Ʊ�5��^j/Ǔ��u(sOf��ݧ��Á�h�B�(_硷=�U{��Q����ߕ�柎��Ve!����c��&!�����qw�5z]C�9�5���<��ܞs�o�@r���m2�o'\ .!uE��
��Fg���3�sx0�+|f���xX��FW^�6��{�w��}�rT�f�=�=9�+��Z[���3Pn½�q_g�
��徛��>�3�t/ƶ��ۋ�o�5����^a��Ĥd��S]��L�<º�]��<�B��]�A
[U�����j���VVݠ�\����N��w��Q��Zq��4l�l�0��q�u��tNe�z*޷�@�#" ,��V��}�e�G;��\P�%�٬d���쪺��)��X	��,�D��e�"��h<��.p��ɗ��f� �\��b*�D��}F�Җ{���u���% �s|���Sv$`�ʋ��Y�����y��=H���*�gU�c����A�6h�����I�r3{NG�.s6���d��䝚Bޫ��[��=�l�s��A[�r4��P#��[�y�V4Z.��#糞|����gu���Tz�#���bz����C�+�
�b�vnzw��'��eyur�?��=����6��(z�[�9�p���v�D�+���rB7γ�N��҅��wu�p%z���b¥�4m�XC�E3:����*��2 �+ (<�����܅����ߚ{���c�gz���n�/��r��/�����Cy⎬ѱg1�w��ļ⸥���9�S�ø�
��r����.^Q�]ٳ| �=��Ytf���}\�o}F�nlq���t��syI���W����?n"���u!�y���NN7���<e̡|��{�28F��]c�
�[$�?+��<�UF}6��>���N`5�]�n��M�"�{g�xC.�M�w7�P���T�}�w�rC�ѵc[.��o�r�-#!�87���v|E�x��[�Ԕr�����U�c��t�_ϊ��X󘻪`3��o�oq!2֦�Y�-�m�6����w+U)r�R^��o����$E�VEAs����^��/�BnT2ۍ��'�"�t����Y��F�a�y�s'�[�u���V��3����-ԭ>�:�aF+ߟ;��"�Q+bk���s���˕4���~��V�X>���<l�������n~��o�ǋ	D���|���2QUS����Q�ϋ�3�۩|�o4��u��MѰ� @�ɩ��:����&����ތ{U�3ݰB/ɍD�o������Em}�u׻g͞�t	o��㞺Qe��B��� Ězh�U�vwO
U�`5�.�V�N��pS�÷�������W�xo-K��G�ޖ.#J�68!l��⏬k�k޵ɳ	2�~�3-�u͝8$���ކ�#Z�Օ�^��bBf��ʯm�<]�99�V�ni��{W(�%w]X��-�������5�oZ�7榷�B�� � ,�� ���w�߅�I%�=m�T�����5�!d�W���a��E�!os���a"Z�k�cM�4E�斡���H�jE!t��A�	OD�6g�	S2���υ5Hn�%���Hi ���&���^?^�(��9�������h�2�:T�!X����k�TWi��-��,|����lh��%;�T��f=���4IK�F��ʈ�La~lH,b��U#]Z���鵕<�]��!�O�9��3Z�/���Û��+��Y�}^��̱�Y&w�qj���)���p�)�6�4�uF:�91��i\��cufS�+�%/����Ac����yاf�4�KgYr̳�9-쬫#��c�U�f�4�G#><F����5�N���Ś��!|�\���5M�nb8�A<�.�7�
��{&znk���U��ɥld���ZU!�KQ�)i5wb3M��&�')�P��2*H� ([9�u����V������o�~\p�׹r&�4,^�t7^`�i���?T���{���N@4<p����z�� �V�2�����pȍď9��0���B5氻�.�g�{���4��uI���R�B����od���ۤ�����X+�[?1�H�!Y!����q�*��X��2�b��a��N�O�i��.>�Ʊ�i�����,j�z���2%��n�=?8�u3W�ϫ�Rd�� (�LQS��l�p�BlZ�����xZ�/��9O Oo�N���]���!g�e:^	:���
"����3ʇ ����"��X�M)�N�,Q��t�{���z}�O5�Ra!�S�)3^Vx��A�����%�&���h�R�̮m|U3m��+�r��rг�	�:!��؏)/���a2WegQ���ۃ���:�Vcse`��cz�f��5�z޽"z�2�) ���3���U��z5�g_U�[���y��3n���^:`�o�?z+�-Li�O0Hd�N:�1hY}_|; ɉ�����ZB�^v���o�������ӧ�|�j�!��ݹ>b챜� h 49�&�e}�2�P��6�b�.F��/V�F�H��WL�������~�����Ƭ.��D7���-�-��눭���v{�h^��&��ě;�� ��������upn�?ρۻ/s�OphW�Kd�����S�e���|�G#�X��1j����������y�z�e��+`�@���z���z��|6� O��?�ٿ��������:8xB�:{F�!��׉aT�gB�|c��v��R�Ґ1��. [yq膞�4��ѰP������	{��M�\˩0v���6;�rr���/Y�7
fʏ��k�:#(�>���uolZ�f "Η\�/+AF�]��*Ȭv�(�u΃�̈����m�0]�sfE��\r`���T�#v��h+�M�b�nE���ޅ:Jp�yO 7�ӥ����9zp�M��%����f=-t�nJN�*��L8;���@|.�E��<�H�� �]��tgۛ��L���W�ʴ��m���s�j[Ӏ��p_V�-�,�)M��ƕ5G�w33�Ih|�ݻ����W+�;cL����]�B��ee�IOy�tv�/o8�d���޷;Rn��g`�.k\z ��{'%�oo}մSם*
�ݭ��Lp���`��_m#.�o8]M�Pt��K��)�m�./��m�T��;Y"�K\�6ꞣ��t�Pt�^7���z���:�D�v'j�[�B�r��H�Tl�dKr������i��_.F������`���ˤ�$�VfP�K%�ׯ�8�ߘ����u���l���Os�jöѨ-�dH;--ͭhG�fsV1
]��Zדmv�O9���>�{Ʈ�%�����t�@oVXV�D�x7��5M4����ZDMF7\b�o-YY �])%�������*�7@<���{[��z��1Z�_�7��<�30�AY�I��0R٪�ZUgl4�eYد���w�5�r1EBվu��l�㫠cQ�"�ŊX��5n3d�I��H����/��oI��i��we�I�٪`q49�(��s����+icR�0�5"��#�b�g+vQq�4�sR�<�^+2-S΄,��h�u�\Y�t��gEQ�U�yN �,<rQ�2��h�XXҳ9Çwq0��Z�R���`�Vpݔ��$[�h�(N7��Ǻ�����#rG-o,\�P��XΌJ��\̝r={�o��ˣ�B |>#�F�%�v��1lI���$�ʖ߯��ϧ��&��=��K��<iF�m����w���Y�i�E�ŵ['W"�= ̅�w�_}���^g�-���z7x���v�����W����fN��w��C�:�[�fv���N�ۨ����v(DQ�>L�����l����yw��E�b�+�)�l�ݝ��Qֻ�ש멡^�u���z̺���D����w��u������k���u�OL�T�&nl{Ǽx�[��!�fwgJ����ױ���N�s�ۓ+)r�-�ޢ��`E�"��QyֺTdH�[���Y�G����������0
����ߩN�kk%���Ҩ���Ƨ-�.Q��d9)��Wx��_X�o~�=����*	�cY���~��?��덑B:�|�� |��-)j��>��c�s����rNJ��~�p�$3@�O�'� ��~B��N�`�4�=w_�[[m{w�BO�^�����x�A��|p�LХGQ^XpV���^wqPٲ<:<⇍�냨��~R�E+����ۨ�ȝ���u�.��>�9�E��D`�8�8�ͺ�]�0����3�Æ�]��Rjc*����ه��uГ[���eB�SP��<��o4�����#�;c	�|N�yf�B��J���faɀ��$��8M��1S;n�����>./�N��`����㞜�c�A��M��f�ÿ����B�1!>������E�H�#Nŧ}���r������3 �C���B�ɛ$����7���~_���鯵("�5~Y����Яiy,G���XK�%�����ka��%����B0in�<JWc�'\�)Yݢ6�y�0��v��e�MD�o���J�ߪ�������	dk��:�{寏!�Z�i��ƹcH�OQ(c0t�-,/��7_z�~�����"���^"��x�+.�d� �O��qxjN{~ �HuVp�Տ��g��F�i�4���,~�m�9�t�<O������9��@2���xӮ<<��x��%�ģs��4Կ ��I�4t�-!����G^��)��������;|VW�H���q��eDC��(�:k�┄#ǵO0��*�!.aTѨ�ܙR��L�*�ȔCp/B~zF����=��E-�.��>�a�{�_?���=b̥��g�7<0��m���k<j��_�xl(p�P�d�z����@(����~Pb����b���e㥍^>�����_��{����i���2�YNL��|k���!��~	�-�K����{%�\ާ6����b�f�'YY��Dh|���MA�C�'L��V��B����(�";�1�����4�#��
����0�=�5���L��޽��K�v�3�S��8\R"F��T�����-�j��(����ޤ���9]!�;�>�׊��X)<ϰ�[M�S^�C 0+\%�+��+,L{ʵ	�j�����J��G}����hiI���->�|F	��j�.#�9�E����W����ޙ]{�	#`��(x��B��ԫ������{t𒵂���w�W����$*g�x����q�=�!)@֗|ú��k�����(YDn���O%��R���(4!`��*xnx�����Ѿ�$F�"�X�!���Ĵ�N4|x�]{<�yy��o--xRE�����k�4�%������a����#m�c!�%�b���X�J������ʕm�qGa�K�q�����rǄϱ��7a��<�:
�)	KM\GQ]3m�Z�7��[�� H! ����1���~+蛇O��	fu Ο��Yx�ӥ-2RQ��u^��Q��Ex�z���@��si��Ƿ/9�`��{3������!@�~^!W1���^~�����c}��mFm��sjB�dQ�j'�_e"G�<2�5�g��gL�1��{Q��W�<��Ne:T���:E&*x�r[02���{��|)x�y��i����&[tmN#MX�{S{�*
�>A�g� ��;�!��xzHg�챞�hws����#����	1��lx�z��_j�P���u�,I6�)GP�B�\�3.�����`?p�Gt�zS5�����9?{�`h#9���"2�����{�$0��?S�� d�G�S�~yA�fq�;ZѼ<a'�^�t8e��3��S�nisd�sL��q'�Q�+9����ï*�ZD�9���<C�Ve�<��o��5��Ҟ�	"2�<��������?�xC�~PhA}���jA�:�\Y��e�1��쭗�_���A��Tf*?��_+�q�d@I��z��y��y���w���O������kv_��(��Ǥ0Y
��F�����׻�(��n��.#Jr��."�lx��CO1�i��h^�W���F�����F��R��;\h���jn��7?~o����T�hz�;���|~���'��yW������?W��|���XI�yg�φF���<Z���#�}t�6�~K�}����W*@���LZ�.�\֮�3[q��(�����S���W��j�x6�xvb����8�n�7f�����#���{��H���!���+M�5-�aAc�н��I�ý���"7S�g��v\�ºLcϸ/1<Ǡ����eح��^�2^�TN��?�y1_�<qt�w��u�8Ҽ%�ޮ �ދ+�v�δ>q5ì��r�:�EE����Ȅ��(���u����F+|S�I|��4�-$��V3Xc<�J�c�l�g�n�2=��pzE&�{�}�� 1�w\0xXb0y�f����{ޣ�}Y�{��>�%�d!����j�-��q��3��4�϶|�f���Q~��T��Y/�E7F�HY3H8�΍�Z��ɜ�m?o�X=M���0C����ƢB���I��v.���K��wJ�Ŧ�Xz	��=t�r���_cu�MX9�U�'o����=CO�:
��b��(Z_�E�5�\ʲ��y���y�é�=�jP7�F��\om�VDu	R�<![���L�};�x߀~�5hu�y���R8N�!�ls�v�)�	�u5�[�r4|5���X���63#DP���=c_�=��u�g�x�m��(zk�O�������4-埑�%���o��uys�C�L��-��Pj47��,rӅ�p�����n�D�-��;���O߫��H���7~�:�{EOM��J��O+�O�j'�ސdJ!��g����^p�8�u7��9t�qXj��m�ײʪ�i�Rrr�.iG�sf�ЃQ�K�-9<�u���8v��+��V��q�P��pve�{�R�^���d��CHX�Dl��䃋�� f�)�^���a�P�>..	1��:*z��rD;�;"]
�Гښ.r����
��� C[S��b�_��Ʀ�?k��~vX�&���=Tr�SyO�8r�A�p�M��	B�&]M��|���jO��`I1�"_��2��^�0���

YOv�EF����z�!��×1�ww,gK�/b��JL������4�Y����{3���M@P��BΜHO(UND�}{�e|A��9��b���� ��D*��Q�q'I�KP��	vF;޻{�ް�����Q_�n3��퓶�6�H�ќ46Pw��e	�:���f�v2��0&LRܞ��BE�	M�c;�{W1�z7Er֠����^��4>:k�'��X�p�t�`m79P�!Jnjv�yr̺�4�R��S����G���-��w����Ѩw�6F�?P�<����xI���b��?xzvw�@�cȈP��5�Y����6��4����/R��V���_p��R���<k�_O ������K���|aZ�Zr�<��{H�~����V�.s�9P�l���~��4�-���ъ�z{ǀc��>�!H\4���\E��C["D�2��2�����{�p��B�
��
�Hg荓^�O��Vx��7����ޏ��� �~�A*�7�b�%�}��:E'Y;���ݮ-�
rXv�:���.D�#ֳ��D_e��hA����g�-%���#�b��jؒV��^�g^Ӭr[6��{��I�X(ͬ��*=ͮn�ПAY"7	}�@��ur�k%`�X �'0���*�\Ӝ��!=M���<߲�@$INb��u��X��=����ܱ?�{�vg��2'}P-Y�Wu���Ի 韶z�u�.a�V�� 6�"�jx�cם2����g�"�=۾�>���>^h��O�<���=¸�/+$�:�,9[*���	��V��+�.�dI�+Ol��ߒC���ɼv�a�������������B�,ZԃZ}z})��3�;�֝d����XD$�k���_7~�ZD�l���gчН荬��+|�����L+^<a��8v��Ⱦ�A}ݛ�}��ey�pH;�a�iM_qSs�'.�]P%gt��.q��m�RF��:!1z�� y{�U��"���y�����_�k_�������H�	-�I� ��V�i�\��K��HS��a�BT�������}3(Rۊ�v��k���Ѧ>p�Fu:��73g.��!�����b��<���\�&9��ϛ������$D|�m�����?��X��d����<�E�1�,.bU�K�a����<����ܷ����������*�^+�ǯn")J�骽~>�zL�n��|E��ǱZ�kQ{��g�DI�>H�w�S�ʾ�����$:���zaɊB2E�[pg��R"��w$SS���f�n�U��Iy�3�-%���w�]S��S8�lJ��~�j��SיL��FV}>�����T|jh`w��Ǔ�|1�����k��H2Q4�������b=�GY;(l�]�䅟Z��tTѧf�%��M��B  �WL�Pw�r�<����x���+�� ��MQ�/zE�z�ā,#J8��}�ϯݾ
 ��ߧ���#hz��=���]��A�1��5�>�m��
>�_>�v�x�-��Gu�P�66�v�.&ûJ��:Lc��u��a��w�u�B�މ��t���r�n����tD2f��랝��\[�i˴���[���ų-�0�����,vN��W���>[]���
;�@8Qr��.�9���d
��}#�bzP��W�cX�He)0L��	9}���Y[{6:\�XYkz��B�񤥬���1��W�r�!Ζ鞙OCզ����Q��U4�(Vu�>6�8��Q�3{Jq&��~*��]�[h��ќ�Hѭ 6�7O�^ �wO
	�A4�5�%���`e8Z.'X���2�e[������\u�k�����Ms�DT
.{C`��z�ʹ�eL������+�X��2�N���d?C�f|ki1���9kjo@�ƥYf����$�i5�ΦC�����Ei�����T_c�ϫ����R���R�W
ҳA, ��-S
�tY�eJ�y p:�ɡ��M����?21Nl�|�1v���7��J�Aę��o�Y��&���y5洢Ǜ�{��3`��:Eҧa���	J�V���v�ڧ4v�O+gw��j����Y#3@��RQ��{�P.Lb���j��c9�-6�,KQ�x��^�ܵVor^p�-Ѥ҈fL�ttE�@ʶӸ�/����ܫ�#\�N_pE^MAFe�vԻv��O�h�0�+�>s3���.v 3�	��&���yNU c�one��N�ru���"�0�J�8F�L�} �}�B�n�]�!��3����1{6jX��#�����e-��[|P��囵��D�%��VnP4ġy���i9Y4Ky:��t�)G���bءMűr�	 %�Qj	
�s�H]J��<�FW�J����b�3�p�(f��q��ؐ���Z�b�V��1h����;�ǽ��v�]��诽c�;s�K#ٗl����M�����}ը�fԒ/D��ǵζ�گS���ӯ\��s�|ǐ��~�ʂg���P�<��:�L0��s������~���'����޹Jy����U{�OolvY|��;F�H��u;������U�v$]q���n-�'�J2Aۻ��M���
��[��ެ�s�ʣ�1]�N���'����!�_u�;2C"vˇ�S��Q:[]��{�d����rG��u��y�XU���ww��w���9(�^�z�Gu��z��p�ݲ�!���ܜ󩓎nk�{CkqU=�ǔB��O2�S��i^��ƶ�緻�(�v��Ǟ[#�G~�����~u��ՙft��5
b,;Z�5 !��QFm�������(�w'���n��@�Qٍc:�;�;��j�u3�(��}�6���3������͆|�~��߻����D=�גK�?i���Di]#
u��,=�.zI�RA�:�yq�5�'W�6�#��K_r��7��D01� W�âQE�az%�{W�mG��������/R*cS�r㤞�L`L*Cp#�4�iz�|�R��������ޔX��'��J�8Ejv����u��A���^(���Z�hPޑ��{�PL�����}_v���P�eI�{S%�(��S�����;#�?��~}��MQ/Ӽp!�04R?p��lW�����%�
�Ȱ�qz����e�|=WY��ڜ~i�#yi��{-6��z���}R:f���{nB�F��\�P�ʍ�f�lw��9{�f�'͕qS:e�MK	٬�1y;K��Tyf�����6y/�f��y��[פ��F>���%��<&8�5_�����=E��U��ե������V{z�3���$��qT=��笜ŧrޟO1da��o-�1��i��~üU��?{��d0h�-�E�voW���qy񚽊r�(M������Y�۾J>����r�,j2�X>>E��(h��D�{�jX�����*."����G���\_'�lB�N$%+AO^��ﺭ�n>�_?>�(��tP<�W���7�ԁ!f�u��w����]�B!߇�!�ZC�a�d�/�Z=��u��4�Wo��Ԭ���B�C���t�!��ica/���L컫���x��,K�����bk	?@8�$�{i�c��o�0�$���9N��<��!C�z����a_��k���O':s�L��mc�s�`�M�qd`Z��N@ R�.�[�`������N��ˠe�8�Ϧآƞ�2���a��fmCs{	q����WD�ZD�-��U_�� H(�X�sk�}�cy=jė�9�nC��B�����w�6ƶC�������h2Qns#��_ưR��5��8}D׭\���&�	�Z�������[�(M���5X�a�T�����)���*1�w��5c���V�u�{�[�+F��Ԏ��Zq�{�]#K�_�C�b�i1Y�c�N���z��	_nT���操�qΪv*���:IM_,�8�����1�k��r�ZJ=���?r����<8xm/1��c"�*�}J�����^��z��~��7O�f��A�H7�a�����ʯ��G��.�3E�8�܇�l���M,mkRyih,=��#H�{����o��bB�zF��_1� e�H���Cd�e���ď�'���q(�k�E��]K��(�ĭ�����ZY��^h3l�������V̵��g/8�땨�eL�6�c����o߲���E�1�������Y�q�/>5�:�0����YDPk�zE���O.R�3���K�����=�/�b#I�?."�l1�Ǘ��
�7����3P�̤@��o���T���~/�@�~���d�f�S��G�5�3)��"$�'A9W��i��Q�wߺ�|j&���4�f�*�B�5�ǋO�UO�;��X>�&�׽�L��Ex16<+�}�����uڬ��8��\��۠oެ:>D�z+�}1E�ވ��qe�c6��8�{�+7}���$+���@��yl'm�ek���(6K�K�����7Fab򴴓ŗk��~\K��9�sO�rg3�u�{�����y�#��;D�I���Ł�8wJZݦ/��ޟ^��U���#��y�Oݚ�����/x�4բK��ä�&�k�H�������"%`)H��ܼ�4M4�k��汐^*��ѓiD�NR��#�	"2���k����1F�ss��%�dPHQ&$4��aیd�t3��ͥ7�}�=Au��N�PRf�%��4�  M+��&.�ë��8�\}��EU��Tp�ނ/��J���N�]m{��|^, ��L!�kk~�p���}qR䯕��5��Je{����Ѣ��%��cK�,mcr"~�j`L)˨�(�v��IMnӺX�|v!C5�%��4�'�#I�	R���<v��@O^˚���:X����2�8`Z��|����3s|��!4����4�4�Ә�ɕ���X�u�>��v�]nf�F�b��"��EL`�O�9q�Oo&0�������w�=�I	�zB��H��:���%�����u�{|��~[k>'pɽ�f�F�1�k�u��Th	�Cv%�D�즹�d<�veȵ	��"�WJ�:���t����f�xMg8��Y������^�dBE$���_f���Uv�K�,>����ӄn�,
�-%�n�õ���"�~ R���F�P��u��Fl�&k�=��� �>�h�8p��^�C�xQÒ݊����غ{�PgԼro83��`#�%����0�jA�1�fj���~w�3�@��|�A�/n�P�5?.ٱ=!��������'7�L�ze,=�
�F�j�)xn�� �u��UT����p+�'����[�2~|`��V���A�%����\��(xgh,h5�ԉ�^:!��;�'���y��vߴ}2�QѨQ Y��Z`�&�Q��Q��yc8�!�l�o�
����+Vyq��y�tj��P��||�<�`�#,��c�u���r�u�n��63�ۺ����u���bT��P䫼�E���%����)�j�qY�	�����k���r;آo����/P����q��W���vȲ*�-�k��;4I��fY!ɍUC���E(tT�R��Y���l����0�����48���C���!��i��e,���
'���P5���[&������i�#㥍���_�$�g���^
F�2񚦈t�V�<_�^��甬�v.�㒼)�j���~\lD6E��`�������w�O"������6�eM�3�0��,ഁ��&�j�!���)��|_p�ؼx�[�}o���^���=��Iq�_X��RZ�3&`�싑&vY��s���z���"˃Iܩ�*���J7��=��TL�U�p6��S�Y�8U��}�R5���\�iD��w���7ԉ#�s%��o�]�ŏz���}MU���1-��	bߞ���E���'̛b��
v]ޑ��q��sg%��X�إZ�Y�x�C-h�\���]%*8�5���~��U��U��}}OG�zog�7+��݉�۩�tg�.c���
q>��`�"���kݬxի���)��d�8t�PL��`X���y9�w�U��%r;c�)���^�����1�A�q�����W�W����B�iQ�ZD>	
q�`�/�w�m�%�Hi��>�Q�>����N�G�8�/Kŋ���aZ��,�A�:'#Vz_�|6��^��������'����a!L:�����n�H/|k��֍�Ht>`�쵈!A|�pR���AW,W�Y��*�������iȑ��DC��^�5!�~��`�|w|<Ku'�q�S>u��x�x�����k?��."���w��$�ݺ~�{��F_��^��P񜮺+"�0�~,�D�&e�9�ȗ��(��e'[ү8e��}��#��<�=�f#=M��S7VE�`��-�̊�rq�wڻ/��Nn)��N���n�G�歭�;�5�k{�'��$� 3�|���_���D��Q�JFm�w ��¸Q��^7'��K�`�ӣĊ���D����iek���,���v�^��&!S�~W�45o� ?TU��)rg���������5f� Ӝ��״�vA����0����1+=���^7�f�sם����m�|h����	!e��H;ZZǇ}��#�e�ݞ^ÜH�x֌5�ET����t��͗'M�G-/����.���z��s�h[Tp�ނ/��B�9�0�o�bO��'ޡ��,�,�\N��1��T����9�d8�_��E��^C���{�a�H�D�,�O�q�(m�Yu�A�,�"z*�.�NU׳�hC�1tH�7��L<ּ����ŗ�x�	�y�p{Ӫ�l��p��LWTB��<�������meka�M��ӗFi	��y��o']v�����$��;�Q����.�r��M�ێ�C���Wu|�����O�P`ҝUr��'X�+�w2��G_�NP�n�󼆗�gb������Io����Q���zy�z�d��vѶ6��E)S��-8pyqcP'��Ϸ՛k=�����Ib�ğ��x�Gߔ���qؾ���pB���y2ˍ�?���T=f��1Z\vs�ן���)������pl^~��he���H�<_M?4Y4�P�����[{ϫ��M}���e���T/��.J�ׅ�hs�S����/Fy�@���pA��j��^0���Y�=�Y�V�h]���"
�ٿ�٘�]R�H��c�>�c�Ś����^D������\꟦]u�[�X��j9�Z-K�\t�'�c�Wz��utiݠQ<�UݨE�,��Otвvkv���r�`���};!z8
�;���/,�˖�,�ؽޢR��ٌ�:[�r�ȶV)���:*��.�pm�-���v�f�y�,r��r�ܥ�xQ�c�7>G!�k�f������$ wt��؎/*U��'>���p5��^�]�vb��8�+.����ն��q෪@F� l[I��Z��7G�,g�Q��u�飳n�u��{�� ��M���v_;�Q����[�p`:����Da��2��ycH�jd���X�+j_��n���4[nJ�]҉�#�kiFt�Gsl0]:�n����9Zfqug�.�&�o[Ĵ�G�S���o�][Z�k7lan�~�<E����xL7�]��#��J٤捖if]�k�S(c�}�H1v�Q�:ͭ�tgf.	ư���=��b����F�s��;��n
�J��ȫL#D���g7���0]�4�T~m��9>p��/�7/&�#u��fll�z�;0W.l���C͹�E�f��ѐΩ��%.�J����y��E��\۝Z��g7����W�wn�-��utg����GA�!� ���.��Nz>�ķp�k��'��O�����mt������}���$�����:����.At��a�t�X�!dmv��Ũ&�<�Ү[rY4��m87�C'0&���<����8:t��A���Ĕ�Y��RG�x��4���ɦ���n����6W6r��N����1@{���K��ݵe��缜����]��p(����9�l,�-�ĬvGY��=��4��z��VnC�Af�C	цs�C-�ݼ��2=f�k����27��$T��FN�+T�9k�1%���z�.F��"[�R5�0'rM��u9}��'J�v�򕶟)��(R�ק�v"�?^����>��rA�4*L��@��"|����ǔ{�?����"/Ϝu���ΰ�뛏Yz��sΝ�Z�G�u��_w���{����ˉB<�Cԑ�<�\�1�r^dbG�J���������=x��*D�c�����s��7;]H��6��/�������D>B}Z<���.Ҏ��v�R]����(���U�
v�\:��pG�QPE�^M����[����.���\�K�z���1ԗ�>�n��ɗ�"���ظ���.�V���v�Ԟyz�޺�v�ͷ�	��5{׻��О�s�N�	�c�G�z�+�W}c���Hbx�,{���jQ^��}���n^у�wb�u�Ɨ\�
<��{��|:�
����)�.o7��N;�n��Rp�!�%>�pFW,�(�a�o����I�	�~Y��?z6+�|3!���r�<F����,�.>�|F}<�����F�+����]k܅��MhK掂8gM�1s�*	n/�)�n����e��\�u�~[/�����QЮ��X/!В�~�P[�r���W�[.��\�^�5���a��.59�v�3$�W��p13�T����q(�S�!��y#�Q��?�\C���#F��3������K���q�0���F��q�L�FO|.ɍl6����s5�v�J��I�;��5����<Y�����]k�I�
�6Q!W��n�VEZ\p��/�y]R��:J�^��)�{���d��-6a�@�3�;�g]��u��u��R�<�׌���B���Y�@>x@�3�N���H�U�=�e�w�T��;rn	�7�R6LAQ����.��YB�$#I��`	��խ�+�l�hE4�>p�rەp�ޫ�9!Y59���ۺ���ǋ��p��="N�~u��.��a��:�%Ċ�c$έ��#Vp��8}v��kϷ�3�r�w�z���_�vw~�}�R�^`�4��������>�b�/Q���.����{���~�_�G'�e����Ha��I��T6�J�Z�v�%�JJs�ɑ/�w6��C��m#^\t��z�8�
�
��$��~��(Y@�c�t�w�6*��T�@Ţq��I6v�s�~� T1��=ٽ�S>	!��6ݚ!R���m:��p^R
��cE���
����/	"\z_�]��y�:�d>U��)eͿw�G�"P��^Hu��!��u�L�p�Ŏ˓m�ܜ��v����d+ְ�|y܃qA~a�iM_uxK�1�>Y��������C��j�2��h�[a�X����b�����o���Ʋ/B�����w9=c��nB�\z�� #-M"h�sd΀t<L��1�7��M��_�����s7߿*ц�!���4�������A|�tf]�N�W�{�0mxf0��:O-#�%�r��=Z��~���u����ݼf�uB���(h�>WZ8hBLR�02+�G�ݎ��q�qN�W?g�Zp�L�*==/����W\)���R�~�F�qN^^Q��Hnӑ�{+�͂��B�7���x�Ip^��U�����ɥ����t}�Z5T��JY\/C)2�el�Bc}07������W�D��� �vƗ=�q!���eHq�x���|:�7՝�B��٘uw G�� 1�����qz��~���0y���g�s5�nx1V�P���ѓ.�s����\C��*����LigN��e	�h9�L�d�C���9^ƙ8m�ȥMR��S��C��ym�J�E��QU�Y���[�t8�{�/f�u�0^E+npdI.#��e��iqfY��w��M9?n��g�Y�|��3����L�R$Z�8����;(@�����C����������}�p�-!���d���^��\ǭx���@]Rb��#��\��5�j��9u �sC���C�?ǱՇ�w)t�I���ꌏj_�D��קb�rI}r~�3׎r�wk	�S�7Y"P�ur_�L��w�y��y�'��y��!�]U��[>"c�����a!�����o,�\�5p������ޒ�/=,E)q����z���N��>��/}~	di�痙��ĄC���ӏЍ5��� �Ҍ�W0s)g�ף왾���T��2B�1�ʇY�0�V�z����?�[Q��н
��X�7Ml {���c��Bd��%�jx�.\�zrW��.�	��MTv��1Qh>�������w��(~)�y����������_]<u��;*�&1%�e��8�;��H�(�A�jE/~����(ṫY��z����ƶ$N$�x��E<a乫��3s���G�9�+�Z�Mi��	�}j��^���|p��-�'jwN�rS<=�9W�엨;�A�
�|���i�ÜL�%Ǫ��h���x�H���rW2f������<t��z/M:�on�1Ť_7�+,?.# \G���ىx��e�?�q��.sn\
�X]�u3�n�Du+"iKa�Z�k�)2�v]Wz���+���9y,�_kڂ�V6�bF�����
-y�+A{�u���m8���О�Q���׃)z���� �V�2�'���v��7�`�	�<v�hPUк�~�1�UǴ���<5p~q�3��%�T�O)x��mX�c�x]�	s���5�'��+=���#5Q�]\�3,hsVT\��\���/3��+�`l�)��6j�#������ɺ���Wt��J��|
��%/��~��f&b>�����zs���=	a�YIb�U��Q����;S���Gl�Z��*��f(J��.jt�$n�gʌhJPZ���Wg���Ts}�y@{���揸 pzxp�X7*];F#¬2��r��k���T�m�BR�y�/Y<_-Hq�Lq�N��}���ǌS��*�+ь�a=H��q����N�V�:j��d����D��C�����9��:z�/K�1�I툲�;1��Z���w(MC�
�h#\*߯�g@F�Dù��o|����!�Bҳ�r|��c<��F;��� ,8a<Քr��~K�}����wO���k��E٢�����z�yƹ�d^���
������4�)��n���V,}a�9�^�zJ�ah���LˀmmL$.���c,oh�;0��v���j�-��Ϋ*(/'ݚ�4�H�,ʀr�Y٠gRRJ#�K�~���&~���#��@o�g��=@64������Q�Ky=���a��^������<�*���F��x�x������(����S�P�_0�������BV�*�,�8�L�3�1U����<#��k�<6	.ƙk"�ge�ӝt�ȉɊ�n��EґwpEk���;W�� �=^�V��$o�N~�<Q�}�Ɩ6�:FӞ��F��FM2�T�������Kñ�-���{���W�"=����H�qk��g�sz\�2��)�\I,V
�D &D7.��"g���[ړ�z��x�Դ0�Xx̧}x��1����5P_<�s�V�W�H�>^���lL�Z�5�T��	��^Vg�s������u��]���|����D��<��=�J���q�M��'$⋷Y��/�� ��:���e�C�A�te��$�+|qsَ�J��n��9xV�-���lP5+S�S��r�'�[ߥ=A$	�ǘλ��ZnoU����UD!���\Xs���Iqħߗ�=aM�f�������Y��m�k7���O$��F���p����o7|wG�[p�Y�����*P���ٺ���S�ڐb���[n3%�;R7.[��1�R��}�Z1�*�0�!�d��9W��g	$��]����8c��T=��]|a��:ؠ橈�������܉��>g��i-+<�yz-S+�s��(�'��[��ݿh7 W��ō���t�8�(nVOb�z��I^���/�ɉ^N��!��l]B8a���L1�ג��#O�s��%�3�;���N�������Tи|���g�c�>�0�FK�h�y*����h��>oK"��B�'�.7cI#N8�)
G)�����B��Oq��s�<�:�h�M�J:j����Q���*���m�76�.�p9��82�[;;���l�����!yqݦ�!���虉����"W�?�i!��xǠ����ƈ�PkO����q�����kbcަ�����!��GRlyH��41�D�)/t�u�ܸ�U����k���Z'L������Ƶ3�S�m�����Wi�b��`.��h���CF2�\g>���r��Ho���f���>�p
qiĞ.=jG�R�^�lY�������Q2V���J_;�:��*�0;][0>���֧0��q��z	w^_�:����m��U�!��:}��lx�S "΃9�f�I�ڻ��:��MEz໷1j�G�-���2��*p�|��c;|Un�8x���VX��+��qm��/���{*1=�۷��YU0���r�ϻ���6u����q�#ZցU���r�nj��^�b��j���-��Bv�4�D���ك)�������ͮ�6��Y��%����t���g�m���˒�m���$����Rk28�*��S�	����:���_n�mP����@/����O�[�zk��̀��>ۇ�T#��Q�Y��6��%�JeG�/y����\�`��0zR����xs'�6=u韢�@����n�,�ٹ���{���C��Ĝh����W1�<n�\��rHeS%��b܇P��L� r*����BO�u4ח�Ma//T�y����<Q�����5��3#_��S�`��m]f{)�����ol��נ��%��¾~?q85��5q��"��=asKw�:���~*�4P�x�{`]x�% �k���d{z~
��F����7�N(�k�7�s����l��6ť5	�ڌ4�OY�G�Z�ܸb�Q�� ���A���w��6of�º���8��T��zc;!�ϡ�ݎ&�׭d�M|`n/��6U
���/_hZ�ꊪ��ك$�bB����B=�!�M�+4��tz=�l�[��S�m�ڮ�E.K�ٷζ�������B�˱wC��24pG��k7&ҕifn�%ElR�۴!�[@�+IK3FXNm�����!�un�J���V�Tz(�7P�eakX�ִ���`�M�n�v�n���J���Ȧ�·t�IGkvn�Q������@,�[�i�ʞ�N�u��Ɯ�X���M=�MG��7i��=��ھ�/ms�3��
[#�S���c��qUPC�*��l��1����]R�}Z��{��ܨVu&��G7��7��q�p�Af�2��;;�E��j,�i�2�2��f����@[��}ґ�Ϊ���^�w{CkV��$�v�\�;�8���VS�|��^Zv�8_D6�.�F[����oWV�=)�!U�ˍ�^'6N�6=�ְ�gWƥ�V
���w��>ۧ)J�Q��4�N��w<��oj}bV�Au��&�j�F�֤HV��4xC),��*)���[.^���*0e���eC���e�k2i�8��	�4�]6ᨯ��r�X�F��)[�+Cnl���/������e2�<;��X�vV����$�c�;��5Vtb=��v�l��,���I���w&Y��2M�QW�T�3V���n�֭��:�$tH;�AcY+��:����M�\<�^����ن۵b���c٦�ԡ�T�A�)v.�t^v�U�N�ܩu�2���&�sť��{z���-�zjuy�+j��j�ܐ�A�R��F"���)���,�m��8ŚHܐ.W}���ӑ�������J��9��@�I�`�|M�B˓M3���\���OQ��K!����7�S�߯��O�O�����nu�f��{l�v������nfg���}���|�\�nK^Ҋ��Qy��:�����Dx�������5�;���U�@�ۅks��Z;ӻl�� �hM\{������:�m	;
g,�ԧb�b<�x������Ƿ����.P��nOٰ�y��lfR�
S�Im�JB_y�z/�S<��㦚YY&e��gq�8�bfQ�����;�IOi:�4�u�n�Ї;�m����la޶�d9��ZY��^u^d������6�z�ws/;;�y��	��u�1<;����Ӧ7v��;��M�wm�v�ݻP����S���v"D��pe졻ή���1u�n�ߧ��F�z7�J��smL�\m�6�)B֎J8�7q�%tGr
J_�����q�c��1��x��(��G�q��Epw^��.��w�/���k4�c<��ݖ2s��C}��$�m���f7�Y.�]
p2�$1I�"5\1�,3WpH��R�$��K�<%{�ׂ��iAKuJ�Oƹf��&�Y�$N�����N���e��Xn{�H;���}F�����k
�+�v��Ŏ̞<�=�-j��bXZ��z����;���s�����yxZ��O�A�vR���"�%�^,��#�\`�2-��7�0�=�
i�����CÅ����?ș�iH����Y~,B.�T٤$s�����b����(��=�a߫r��Eh�X�˘i ����U8�/3\\k��Y��߮:�Ĺ�SUZ�F��Ld�u�a�U�X�8-cV�������<�*�}ePe̩AӼ<���ז�[S�^#&�d��c'��n[E-�V�q���B���1��N�[�T����g�s��}7��ʵ	\�OP4���I61Y���������
k��ay�Tǹ8�xͧ��k������
xYN2����4u���ЃUZ�y�Ǘ�-5i�����L[�jt�׏���D{��0k�_A��c'��D����W�y��Nݞ�6�(�w98Չ�F���l�e�5�g�̞6����������ߙ��$�X���ֽ�y,#ɿD�TY7����ݝ�����,N|h��+E����Ϳ3>��8 ��4�e
�����||6�1c�慵�H﹎2��dR���r�]e�𰼙�`$MoU�jH��{���\Y��}[��r�̾Y����k�)�~ +��Z+B'F
Ԧ,p{C�2��IQ�<d@�����]��>�z�_HE齺4X�y�g���ʱ^�������x���e�\ޜ9JU��9]�lgF���t���J�I6�m(����$���KzS#�}��E��y�kX��y�ûqbac[�����u���8����1��ym.�gyi؆ֿO
�Q`;���(��W�"���ϟ<���;˼��d��ڙ�e����5"ɥ�?|ޟ����H:G�Ǎ���$ix����/4ۧ�����TI�.Cٯ�.���>h�5����2b�Պ���S�&g��@ʬ�x�"���1�(Ԋ���z���㰣��<�y+d��8�1�2��Bu�ϯ���S�K� �]sϮ7��T�����9QC��46F�!���_�����E�c��de!���iğ�K�m�.Z�	\5��$^NR�����[�7� �맯�B��2�e:���5S��|s>�'�mO8,n�r�X�e��tgI��7r�z��x�v��kŉ��軞�*�+���L��v	��w(U��C'3�K�����9�%-��I\]�[b��W�c��U���eUo�fbڸB�ۂF�Od�����d^�z9>e��KX�P����lR�c�ʘ���@�� I������-#3dM�(yq�i�.�LH�����5�7G6�jx1�c9�O����d~d�c�������a���f��q�@��y/j�XB�����-�����w�~�hf�C]}��6f$律�C=L��PkK�^�泗�3��.w�����ď��I>Ň��x��&4!v��(r^yr���~�k=���R��C����J5��IŵGǍG*��z����go�tÃ'�j��t%�"����o�����R�*��u���W�/�C(�x�D��,��H�GѢTl�uC��t�P�8�T�Ia�S�sl7��Z�ۙ��V�+�1�u��dr�Bڲ].&$t�d@	��tE�F�B�/R���<�DӖo�f��6J԰�!R8뻡j��G5k��a;��q:��k��!FyK�U/a�W�,B(V����[\��;�b����-Hq�M�S�/^��sf�`|���י��� � ����X����w3o^�?)�l��>T8R7��0���:�-�t7�㱕 ������u��z߬R��|��8��ӏ��|N�P�EZ�{�އ�^��T?~b���do��O��c/�<�h
WY&W&�s��{6� Ww�#Z�\_��8֯�=���M��#����#�`#�3T�]Bya�dL);Y���YI���sʬ�C�Y����S��~*ό�/o6y!�ms�[��J�lh�*��-�\�/%uȷ�ÃwSc����Xvy��^"�VS���|��z�d��b��ޕ��Ev;歱J�e��t�[�K��Cr��,�(����ǧ<�6$Z{"/E]�l�|h�|�{��,����\c��}G>ԧw��ʳ���t�<0�Cb�'�ˮ���w�{}ˬ{�f�3��>�ǎ�丫k�[c�Wℚ(X��� �Z�^o[���ϖp��rg���5�/ah�t�--9��y���J��b���D*������|�ʼ8�	�^�V!w~��z�
��
W��Px�*�����hY�I8N��JT
R-�R{Ա��8v�����h1ş5�႕�����}ے���5��ã`�0��U�k�ߏ_�������m˖��I@c���K���j?���;]s�,l���$/���8�{�Ӽ�����C��c�a���l��,�K���S�Ȟ8���}�#������H��8Ϲa'��y �.���ǣzG�rx�'k��"��ua��qMޥ�Z�.a�=N���SUڋ̚bA��56VB{4_�Sދ������Yg���e�՘�$2pػp��Lm��y}��Ȧd�6��G+z��KNA���2������C`͞ņ� �_��4W��S}�u����B�P�c�|��s�Ǡ�eEZ�����:��pgtNO]���)صz˛�*�T��#�V%�s���c�wF�_���φ�@H�W��y'��XKM�QQ�>X2�U<�T`����ԛe:���;!���}��q������F؃}US�>y�[�t辻������,�5�"ڌ2�^����5/%��#�J;Y�Y��"7W�Ӳ���RӜ�4A/�/�T�pVj��d�<�v�#����~?Q�� �^=�48��>�q�/n4��v욨>{�U"�%�=���)q�<g$V�}�a���,_��v�0�����O���	��!Ձ��BT�8�"}�" )轼�p�<��:�8�JU5��b���b�Ѷ��l!���o�;�7k�S�]z�v�ڲv����"1�)��hj����S
P��yT��vӏS�9�.9�����<�{��AwF��p�Aeg̦@�<��p����y߷��������i��Fm��xk��:�\g�~�62Ƨ��w��}L�r��VG�1��bE�x���E2��#����G���Q�4��pu��}jN��:��5q|��{N�ۆ���_o{��Ig��e5"��P�^#k,���0>j�E�������om�R����ɿ���a�{~�8�9��ǲr3:t�"V2[wyW:��K��Л�}���1��i����ŶŠ.xw�.~���RL��������X�̛:И��
�֨���v���P��H�e�@�|��F��ۦ��B���9���V0�Sj(T�5�LV�E���=��8���Z]��Ŕtbr�H::�^/�[bU}Rx_zn�%J����Vv�N&BA�Tʊ�s��i�o��Rf�w��{ٯ�9���W�e6&��f�P���'�&��nE��Y���~Qj�$�k�u�3Ԙ'�G���6���vu����C�x��B��$f��[\9'K��#j��_�c4q ���"jaD�VL����,h;5ضT�(�i�;��&9���_xU0��g�|t$�,阉��4C�hR=r�����$�Ӧ<9V)^`�7�'~�0�%k'�jl�!ڶ�j��7����x�2׈�y�]� �D>��d��Z���jS�/|��o��M��D�_e&��Z]&lZ��jݞ��-)��]Յ����p�DO
��O��U°��`"������qY�ր��䦮�I�����w⥆"�(��G>w��3��|����y�n������&p���* ����� s��HaN�Mb{�j�J+�5]�]ǃ�Q�k�౸��U��{�p��Y:b�X��D_p�2��$v��;���XU!C�jf�5�N҃xMRDdq��\���ۻ�.Y�iΪ��P�,��T��h�^L��-#��v�c�v���شR�SX�3���fP���#���y�Rc+�D����+==�$4��}O��Y��S�	$J���p���wS�N��qa�����S�E����m]��I���ޫ��-��h
n���V�s��z�(:!�R�ݼ���72,�b����|"��%B�aqI��x��}q4T�jg�ȇ%�[�Ek8�Q�n�m�!�Ѵn%eT)�3��4 �����h;��Z�xfhzu-�(W�6��״/7Q�[����
���E�f.2��NOL�z�`OY�뒅+�=�Ć�f��p-5��������])d�\b3�t4�$5�Q*���oX�l��_���7�_%��kz�P�U5騜ܜ��%�eCI°\Z�Y���6�s:2,B�mJ�n��]�b��[�un8/{Su)q�
�4�j��6�Wf	k:�W��:gr�T��\vR�`����ˉ;������xc�"��ʃ��ҭ�3WΝm�[x�"�E�h�Ȓu�1�5�m��Ō���RI��2njړ��P�n����f�������6�Zwf���K�&:�[]*�zsy�`D�j��V�L��h��X�M��FEҗdn�Հz�w�׮;|�-�FYm�;�ڧ�VgL�¥���������Z�c�;�N���ÕQ��op�����n�PI��
m�[b�	��������	+8η�Xw%���!��W߇hT��ɼ�"Ge��9��ZE�-�? �4Ea����L'�2��㷷3o��ci�շ�v\йν���]˫�C�[��&ܧ��MY�wk�����.�R���[�	�q��EF]�0�U�s���I�s��|�G�y�e�O�Jh�9#�v��I����3�f��R3*�&�v�f�{&�Cٝ��p��1VoR<�ŰS���^t�Jmg]p�RG��=�����=Y�ۚn�g�&�oj�X*�9�˳A��㊓���6��#�������wѾ��<��Dm��a��*w`�����uA��VT:,�[f��ُ9�mY�!mNpF��#=q>=L�󻟶��
��Al�o��]V:���eaϛ*�B�R��uaP�M�m�_oM���-��%wk���kI���*��&���Ibr�:�0���;������SzЭ���cL��٦���b{�#����'c�ݑ�$���}ss��<�ά���7t�ι��z�g�q��2��d}���}�)2(�L�Vn<z�z�ot�S��i�2n����ﯶ��2?%��kn	��J.D�퓧RQ�p��r�U��}ﾋ��'�⼾��w1qy2&�xC#2�)Gg����}��K̹cMry �G�V�-�;t�ux���3�����y0�k�FfC�ll�U �ԉםp�vX̃C�TQ�%J���.���٫�᧗�Ѹ�%E���Pw��D�U:�uW�m�fn��������L�A��ӵ�������d�F�v�W�{Y�5�Jj$d����/۟���{����F�Z��d��Σ|v�:��� �]
�^�Q[z�Bq�p�8�U���g�}���:�vKkb��GPxK
��<�v�9M	�:�F��͙��@�{g�n��^k&Έ�'w#2X�m����k24�m1НӔ4�+y-�a�ukWkP&^$�����l+�&48�_n�](��g&��i��_�^�Y����}V5׏�jW�ۭD��ͳ��R�L����!��q"���Z�����&:�	v򭊺�l\�؎\W&�^9޿���M-�D�^�MԎ�<p��{�V�{:<���C��i^�?Y{\S�UPã:�^�g��w�۔�i�iIږ@�)�u
-v��h���/����q�#��I)bR�\��!�l�	�Q-6�)����D����Da������hǩ��g{�X(�s)ŸW�{r�v-�]pZȒK؞g�?�3=��Q3��A��ËئTLp�q� d��أ_�@7�6:���Z�-�U���MQ��N��eNU��no�6F8}[,Նo9����6a�mað@Q�,v�o����e�W�oY��z�9-�����#��,�W������p��qEW3����H�ۑ��bE���f��^pS�"�dh�VV����5�J����nT�^�:����I���i�bw���Ƴ��b�iZ�+��3&i����ɸ;Y*u=b���=����Ƚ���n���]��MK��2<��7[
���`˝��5
���q�5(c�����,�C5��E,Y}b9� �����xjk�'�b�@�d�Y*�m�'DJ8Mĵ�eGk�����
}â�NE�g��M
r&���(�Ll��C�*�8��{qGJ�D�����Ұ�EV8���{����*���_L�����m���R��Z��? �ͻ���9�*)�$�é��Sl]᣹A��ܥ~V��{�x�,m;����u>�p#�}1����jt滳p0�b�gd�J��3gW�++!���^r��2����0m喴�v���P��
�a�9��g����W��RTgڒE�f��켷4�@F�����l[u���#&�}���20�]�tfu��L�����$��sQ.N��=P�W��^pԺ,�^�s!�Xv�+-��=��͜Q&�W�^�f�,�Ә����drh^�$m�~��j���Ɋ~x�]F�^�a�}ro�"���a=��XYW�<��ġ.Fx�I��X��'���3U������[�6zVY������&wI�ovB�Z��O�b��LmOѰ���u�:�FI���F�����-����*D�+`�'�+�--���o�t\���Cd���-�G먑B�9Tk�F��WZ�����ཱtVR����P�Y#����'���I�e���)q�F�9sI\KǱ2STF>O70�Kd�h�l��v�br'�+z�oEw-q�($4��J�p��ڊ�cr#���lI���2�g���9��!I�72�F��G	֚Pf�V۹�Ő>U�C�J�I�&w�ο�Kn/��=*�ݫ3=0��ig�����81����yԫ̄��uv����[e9=��|��#'7��w^�o��x�*�\nu�h>���v7V�;��OL��05>3�6Ů�[9�����j��;��M�Z�q�e��(��q��,��)AT"�'ɹ]=N�4WT>b�L�ήg�/n��r��v�ۄ�kc$w�%5�_���}.��V����ayF�Tu:5 �-hLWXb�[cFѹ�+�\���u�M����6��GR$M�u�`�KY3h.�-˼����*��Ӡ�Q;Y��)��i�]Pl\�Jp�g��k�r���xy��^�a�/���N�,.�[���y0	���佛�WC9��CY�&Ywx��3�^���q�s�y�G��[b�;��L�6�vʗ��{3Q{�<��r�g!<g^qeWj�P�ȸ���Ӱck��ξ�3w[��n/A�g&j:I`��/�)�cg�wXWL�;�k;'}f����䳼��]۫�|�V+*L,(����7#�����y�3�V��)�َ۠b�����jٜ|����}�|G	}w�r����&k����-hK��R�-�Ûe6j�,����&lpvM����]���������8vN���ٲ'�jh�y$L�bE���I������QC;&���l>7!,=���TӬ֋��/g�9;7ZƾW��7z�8��I�Ju���z���Cz�>j��y����nN���$^d������h�vȵPBص\�ٲz/W'{��.a�d�p�,#
/��]q��Pع׬8�e���<�h�!}����J*yλ�nɻ�C2$�������-Fn�1��_8U,NrO"��°<齺:WE�ٔ���R�۩$��PG����'y�y������U����QzOc�E�4.8H�p�|���qwi���Op�+5f��NLr�{��5��&������w}w6Ɣ��p io�t��I9���X�k[2�Ĭ�7�
�F���19�k!��#�mC��({�G>�պ�9v.���Gٚ��ͷ��%��j��2��0��4tl�2��3ڇp-!]=C	`3U�2Ӵd�P74�2&���i��qc��������c���۫�C|˕�9k��ؔ�����u���W]��')�"n{cA��)���z+렆�}ǛTmƱq	��G�=��2�/qW��'�fQ��bSxNZ�>R�c���/I�n�u/]�Yk�j7I�n�_�]q��o�f#
�ʝ`d���fa���MCA̗�~8��{�sQ��p�_v�Mz�+r�Y���dH�I�e7��U����E]t����Wu�������G<�q�i,����|�R�HW3"Z�qt��b]܂�����В������W��N��y���(�4�Ǆ�%=�Y�H�
��&�(DqG�'�����9�~�ۇ�t[���Ae��I
cf�m[���ԙ����/�W4�m�˿��ǫ8��z��R�b��a�I����SJfb`��a�j6g�S����^������R���s�G�U�U����׫6���4��3Rz����ʬ�B�`wq�89����J�؃����Ԭˍ=��b��}IX�hEz�O%�����aG�����~��`�)����X���l��_�3����O]�\�7C�KQDz���N*���1��
2<U��7�+�M]�� �ҙ.��1��P�����q5(i���7��j43�� �.i�3NIMƌR=9���TV[�\���/:~FN��g|�ef�V4&�d�NΙ��q(�;��<ˬ#f
�'Zu{n^]΅��}q�)�u��wB̍ەv�Nsq��6kD�"I}aβ�N�n_fF!��u��F��J���V�Q����b��Y�N��/�9L�\����[�0u/�q�k���~5]��C�I�Yh�ܳ�yx��vw�T��k�E e��C�dXE.qۓ�ޫ{~��7I��3����G��.�h�_#��s����٨�#��yk4�={
"<f�����o�!� 2�wp�p:�_ :f���z�/�U<��f����M�}�Km�Y��.��Ypn>��c]���k��k���1��+��ʫ��[\��`n�T�e��,��W}��w5.o�J�!R�-<��8B�p�7�ܽ�q�AY�a�,���Sb[C*�wuλUl�Q��n��
����;]bI"�Ĳ�S�q�v���)�{&���=����r=�j �v;T�n��R �_T�z^\F��{sɜ �ͭ�R�QP�#vl�u�.�Z�:%w>���3.G�����jP�WK��Zc�ͬ,�XQ��O�9�q�:�BX�"�:�7ݎ8���2�VyH�C�0�qB�C5���t���<�<AΆ��
1�/_շA�V�ӻa�bo{��1��̭כ��
�X�CɛzVٝ��
����SHn��*�[��T�\�Z]���S���i�ΕsY�ټY�ا y�[h��m��U�1��X�y�����ծ�t���
[�wt,NV˾���w���`i����/��+��6��gd��d��N_w:�WDdR��Ri:Ww0�ol�ãG6���|��a�R`j�fZ��"*+o�'k�{�*���obv���z��HS{������ѝ��_a�q�nZ�3���Vmqw�%1�\����]�(��N�:���v����볩i�J{SM]ӫy&]�:�n[9+��KhlB��q�^)���-���R�C�2�%TtuN�B
N7���-v�R��c�O]τ�)�t��� �o�Nʋ�k~�)˵j���yw��2k
Xd̦9H�#�t=fAKΊ�󩹖�Q�7�jXv�_G5���^#�錙̫�RޥqԖZ�u3YcټY{
u�2��T�`��4�g.qq�#��ΐ�Q�m�>���\��������h�ֈQ⓻�}�|}Zk�� $^#;Fdx��)q6�񪸲l������U�~j/��y/�2�h���w����
�x�_�RreI(��l�s�Z��o�����5*�\���<��9-̆37S�3�j�E��b&*g���"v#˒��#Ju�n��TW+O��ד�UB��e�9TKʧ���Zx�'u������W$V�Y��J�!��.�zH�e�l�j��U*U�hk��̤�b�UG��Y�C;Z#�]
[��"����RH�+�In�v�����W}CBF^�ᘨq�mRܢ�s@z��"Y-D�(\�ܔ��H���`W��|��m-��z5��I�l�-0>���W���^�Z��4{����=,':�*�����P��Po�;NT<(�rp�.�;�Ӂ&��';!ք$ݲ�1�m�o�5�R��%&�w-�(nλ�Q{v��/M�3*���2vo�q*s7�-;�+�������*Iۼ�l9x-On^�dJ�0^�%6`��v��%!y��o�,g?S��^^�ᝇ} ��G�`8en��rH���������)ͤ�]�����b��ڛ�f�'ݔΐ��&m�.ň�B3vI��os�իs�������*�(�v�v]r�cut��z�^�����/0�)�N��b q�P��Nu��qUZ@x�C�qJ�g���q!X��x^�ݎ��d��IRz[*�0�MF�|}P]�WnM읉㤋�7d��{�)��{��<���}�Vh}���]&�i:��J�]w�m���� t�[ݦ�3\~�v����&P
�&���u�ٱu��x�TuQr����L��F�á*;{|���l��sW�ݛX��Q@�jV�\���t�����B�M~�f]�r�3�o/��ᢒ���!���;���1�����B'N�ݕbU��Zm�"�Bn[c`ݒ�,��S=;Gc�����r����6����J�ub�F%&r���f8	k��z��X&�|d�C۸i�R��{c�|u<��i��������D�K�h��ځ]����5�����^/ٷڌ5x���"_x��q�̘���ZaEV��&�+������PzAqr�p�B�_8����ܡ8{�u^��[�%�;�5��+��dN�Ǹ���b�-o3�+\%��Ew�d:��1�"���4��+�fᎳ*}�WI�/�[޲�54�Y����͟3��E
Yg���Fj��� sF���[�_sW�1H�d����X|�O����2���[���]sE�^��9��8W2�]t����}��^�\QP��r^��h�U(!~?I.����ue��e�Y�\������c��S���B�sY\GV��tQu�ğ-���Z`\{�F�Z��Q_C���lvWF�[G���]�ܤ�[�<<#�׹F���I�g�{���y��O& ����x�vN�U&�.�kFf��IѼ�_H΅Z{pl�ٸ�ga������.���pRm#����ɞ�Ә��|���8ع9Z�¯P�-�1k�2{CJ4�./;�E{��C�b<�8�w�I%�*�ݕ������<��������W���J���z�w8��N�^�Y�D��9z�k%]'"qzA`�.�
K����P�G��Dȭ��曊�m��+��������^
�´7q�8�@��ͣf�^�������B<�34u��A<1��ꌒ{��[�N(:�#;��lX�X��`��P�yW�2����Lȣ̈́�%o���)�V��X��'�^�qh��)7z��!�-�s��M��%�]Y[���<�y�T�r��sQq�C���Mn��>)��]p���G%�ȋU�l����pmUp�-���j�&��.g6]	��fd,S�@��Q��J25�P�h��F�4㈘N���é�|�����]FxOk��P}�)g;�gl���'���c�oaMj8"��&�4��6�<�q����O:!��xU���Q���J6�I��m�͗v�G+Rv�/�:����Ѕ
I��ezkL8���F��dub�F��՜7[��=,�g�13S{H8�̳��wVh���i�B"$9[���4L�ӔӜ�u;t�� :�)e��nF�1V�B=!:��ޚ����|��M���VVT6$���������wy#�ʷ#^5�'���p�|��f�y��/ԌϬ�}���[�=�o�	U��gY��֓ͥ���c�}:-+�7{��Y�ӏo�q���l{����j:f�M0�"�,�=�����si����H/i�.�y\3�w�\V������XxJ��ag��HGPM��w�	�&<ռiy3ݥ7Ä����t�D4�VI�����{�lfF�%�Q�.��j�!��z/�nL%�k��۴ *��ثb��0vJV�x ����>|&���t#޻:���Sv�5w��N�Q�VU���`Hz1޽	wI4�Y��.���,X��\��v�p[���g;r2����+w�e[��Y\.���b�La#j7o�r-�C�1��Du;pjԾ]�y�ɷ"]6���)Nw3|��ӂ&eė3Q{u�t��Wu��*�^�\�K]`̑���U�����7ۭ9���o\k�W��-熰�}�f���Tnz'b�o�c9�J���B�r�<%F�P���3J��N���8���쇘Va��)�m�K0��l���=��Jr ޴���Ȑ��"����1c{I�ކ&��rvy�qfO�(����x�+�ܟ+W����E��6Ϯ���5"���v��5X�S���r�q.�iB܎���B�E���nA�NRNR8�7�-��f����_�Ҙ��{���V��,^kPܭE
�5��f�ˇw�ŗ��2��SW�<�E�������6|Ү�����M�]����
���n�fu���_�dF�;<����}��U�(�U͉�/?a�5ꌨ��;/J�ӛ�y����b$}��̭@��A1��z�����A_'�hz�u^���*m�^ry��^t��ֶ4�և���-[-���'5�#�ͬc4S��:Y<�[���_#�%m�Ĳ������m�@K�x��b���� �D�f�[b��F@&����jׯ���no�������aN����O�t�"%���J#,�^�Nev��7T�yj��5p�j�*8��愔��<A�}�$�#|���ov'�$�� (rN+� T��Wiw.�f�iI���:,2s[/��?Y]�� X��Er���[�{�����\W+����&2��Hujɲ{�QS�%���&�;2���F�6z�b���4!��©�by'�P����7�4�b@͞�jwm�$�e}�梂V9�����N�^^�z�\:����'bS����#��u��j��m.؛��$ c���{��Kϊ:�n�=�3X�U�j�1����&Uj�J����F;T��飺�]�:�]��˦�N�2��|�R
�}����y]�q�N;�StS�5� ��K�ju�̨��ȡ�C��=��~��1
/j��K*Q�ʐCZYq��d��w~��_8]����Qa�>�%f����\��+z%C�e��ytO�k�U���GI��ՙ7	�I�ܤ%�ܸ΋�#mQ��Zwq������|���853?`��#}���0zs���os����#vyU��g�Jr�8.�ۋ��8�|�F��zX�|m��ps�m{����q�w���ߍ>Wz��D�ᙡ�3f���Q��НCy�돛���gu�'�B¹�t�w����Y6������a����(G�}��ʄ>���B@�$�K!
DT-
?���
��B��*���щ�?�h�X)�c��h�\
K���ܻo�j0yz9w,X)B�)�)T�
E��TTX)DT
��@����
��Z�@���������
�� B��$�H� B B�d���� B� H���� B`B  B`B��<�`0�MA�� Z�J���W���F`�W��)%-ZJO�?D~�@@T$aR�Cؙ�N��W�x�ų��o�!AP>!p��
���B�/������ߘ0-�A��h>��4�Ӑ�oh���$��!Y3|R�I��1�����C��~ο]Ϭ� �O��t��
�"�Q�DQB��
F���?�/��>a�P���x�O_��.?��?�>���f?����XVQ��ECA�_�S��'��X}�HF���H%�o�L������`h�F��T���X��P�?�TZ���<<.�X,e�o���P~!��s��<�~Ha���O���x)@P�φ
z��,yOо\( 
����Ĉ���D���
� V��
��b���Q��X*�����^��{tԹ��P=��(�0@R�
T*� ��>'�!�!�����'��_�?�C�>�]�+���?��C���,~�����d�?� ���~Uj��?:=h��DEC��Z;,��k�G�������~�=�����G��㟅�z��ψ����~?��C/��c'p?!����>'����t��������5��}���[C��S�� ˞��Ϩ`@����G�l�x���@{~����O��QP�܀�������B'`����
d�>E��p�P�{��{�+)K �Q��`PAC�>�D��Y�
�L& U
��/�����>g������=!%�!UC�z�hV�=�2D.����E�%�(yr�`I��%�فEB;�>���~Ӡ?$q� DT+������E��w�<D�����x}g�����>#���>G��O���>�}������."}G�}K�^���jX�y�;���؜>ȟ��{�[��,���`������P"����xc�|��4F��i �?O���q#� "*��2~������a�������B��Ǹ�����3�52!$������.-���G�p�� �����vьS#��S{|,����&?w�>���v68_��=�p{�P��C�G��zK/��F��=��!���Q	�>��=)�z$_M�)5��(�<��G���L�O��=��� ������X�@���hw���q�_��>������� ���#���A��ᔷ��Xp�0�m��5o��~e��>	#���>��?�"���{���\��rE8P���52