BZh91AY&SY�m��;$ߔpy����������  `�~[� �UU�U@��ڀ���TUJ��UIQRH�@H��)T Q�d�R�I#8P  ��U ��/��s���ҧp��v�ծ�Ǫ�픯*}���=}�V���ޫ�{�l=n���zӸ{��u^G�{U�e@;�  >��_GF���P���h�*/j6���c�yM�i!_u���G|9އ�r����M�{�z�ٜ�[р:�} �)��|kU/���,z�����l�ގ��l���窣��ݝ��7��vv�ڛ�N=z:���=rt�8�(+�����5}eM{����ī���׫�8��0=���;�y�*Kצ��pz5�rk�p �A���o��I��Ï{�R������|C�^2��8�����5���������8    
�  �
� 5 @ ��T��)�I�h ���2  ��DJ*�`	� `0 i�R�J��4  CF��)� ����`� bi�  "*�50FS	�7���TڛS�i�i��Rzb@��R�HѿU0&�A�0�i�0 ����:��QRB�F����� ��6�EL��" )����UTO��P������˅�'�ḁ!"���B*��nB���%�%�� $v�m,��d�[m��D�@U@7���~�~����������(J �茟�?hm�,@�`���d��E��f��GYn�v��3�a� �D�a�s����Y&�S�i�vND��J�w&��"���2��,��^��N��[�$��pA4N�I�XM�d��#Xd8fp��Tfj��P�MQtw��/�I8�Ĕ@OA8Δ��6��+͕�uZS�)�Lњ.΅A�Jl����M'�sm �n�F�\��%�`�,�i:�V�[;$�t��,0��F]���q�L��'IcQz��]��I���ȦE2��A�'h�Eٱ�@�uQJN�)Ij
Vg����f&c2)��g#9dfu���U��M2i���ueM�P��E�I�̄ɣK����L�d��l�`�~^.��.
g\��u�g1��q�F�ݝvS��
�K%�O�'JXR�����٘���溲ط��z)�!�M��U�;�2�I�*��YO�31z���qt�/��u�uTsKM&!�����gY�e
��(�|��M�u\�y�&i\g1����Y���bV�,z��(`d�-J[��%�q�p�a�;��&V;�S�,�H��x^����e�I��h�E��'ZIM������M%��i CpV�^n��Ɗru�L8,d���Tf�"�IV�%�J�a��h���)8'`^��LS�q�XN��30!2n�1X%�u��Xp�����Y&Eڐ�U���^nb�0�}�&^7ϣdܛ�Tfj��pS�|�ﵐ_�q� ��0���h�i���l�êґ�)�Lњ.��I�w%S&�M�&�Is�*��JJ���-QKL<i;�V6vId�JXFj52R�O
�8�N�K'I�/e'(�E�Fp�eh2)�eMQ�3D�)їe6l&N�VV#XTN���F���e�F�/RPgX��)�x]d�d�J��I9��ˋ(Qb�l�K01�T��ILBV�'%�[)�h�&�	`���̊f��e��Q�6�g^D�K ���XPT]�G%�[)���5H�J�C��يҭ��Va7e]��l�<γ1z���/WnqԶs����6N�K	����JR^����U3����`��M�b����f;�3���I9���6�,z���6XVvCz�%���.�l�S�L�pSA#l��D�Uaz[:�g\��$g�\�Ѷ��l4]v��I��\	&�M���X�X�NN�J �I<���d��3d���N���.��M$ta�IeN.H�&�E�a��3'
ܘ
��vS�+zS�IV"�:��{f���	�F���+�b0���0�B�&���SG��<K�Aͤ�A�%����r��m(&đ ) �H ��xX�Ҝe`�if2��~S��b8b�Σ�W�o�a��N��I�E�_��d�*J����E1.Ҡ�ㄤ�~b�%mƻJO[s��菴
�m�ǋ���:�{��|eeF�>W��a���I��!LX�+ō��4S�&�m'd0�a����k[15X�NHLd#��<,KiN��f4�T6H �uX�Al����&�e��AΤ�+�3��w�)
��U	i)��)��p�
��5h��)Z�4X�MV��*CZ�L�0�~g@�>�4va�J��Np��+FQ�o
bޥa�ōE`�Xu):��5I5Ey��01O��=[�5���7x�o��cK)�E�����N(�\��>lɌ�V:1,&7�[ղζgK�)��fB�FXvXzw/��t���ņ�]b6o-~�\ݮ��13a�Qf�8�qz������:]p֨�V�`��r��0p�Ɍ�X�d��IѾ�e��r��X��2b�(�O��8wX�|=`؜�^I8 ?`xAb�8��
x��pQm'XT��&�^a�2Ia���H\�A:J�]�A�c��b����/4�,j4-�'tT�7&M�����F����3��R��LOŋi,h�5�I�*nja���fO�Ɍ�V:1.�IW��Av�:)�m*�V�Ɩf��'-�Xg�����S	�r���#�mk���Z��gw���f�z6�q��݌�냄8��zY��a��ְr��`����k&6�bwI�`����A�e��-o,k�LU������C'i�A��AC������<7�0�a)0>pa�0شPb�����8�`1%�����ƂEn�0��a��ؑP����,�2�ka����A2���1��×��Yšva	$D׈�x-y�`-��"��I�l+�(F���-ӭ�佔�N�ҪMI�yI2]x�2�f��lݲ����)$�)'�ޥ��Ru�X݁�.Y9B铘�8� 籒q��d��ɹ)��/)D�{Fh����]^(�'å�C�g�H���I������t�:|�|Y�W�����q��e�7��8ͭh>>3�m��}�jc��a�x��69�y�=�aݱ>wO��6�: ��7��=�����S,���F�wI��qVe�?b�0b����֤������6��RAD��9U��Mږ�R�\mQ�5���j�o,�k��p�v��]���3y �n����gV�Gz�w�ُuٻV�w!$�9��r�kT#�"ԷEF�n%jz�{.����i��K��dS�2ِ9K[�.�}&Y��d؂�wU우j����(��wN�����{��rv�齛�rr�7�d�ˍ&�N��=�n��e<���?JS'u��}Cr��.�(�1u�]
u{S�O/��Ok^xL������Z��f�X£�7�1g)Қ�1P�U�U(XaH�1(�&-���ت��30_J{3S�f���8>�.�;ɭ}�cε����{�{��,�ρ�:��΂tY�6.�ŕf�L�$����Q��>��0x[�W�1[~&���w1�o3T��f�Fՙ��Ңo�@��9+	��}1
.�nLA97j��Z�1�ǦUS�S���R�r@�{���A��������a}+�O:)]:N�xw�?0�Ϸ3l,^ے�a�<�ҫ{"llk��<��˄�s��MP�^8�gU�R��0�rkN��Ibf��]U�
�}��ea���!zN�0.e����c.�3��$R�l�r�]p�����;��g�wج[l�Q�Ys��a�}�6Ͼ�0���wҬ�4z������\fg<�ݾ��wK؅HMe0b66�zfa�GEVc��c�蟼�ӏF��x�ܒ.�)���N�:�,�0)ɺ���N��V�f�i�ςw�6N��i܇ٱn��e��^n�����f�b���1Jil�"��ls���tڵ5qQ7Ʈmn
w�ziT1��2orx·F�ˮ]N�=+�zz����~f�na;���{ �w�ڴ7��~:}�?3��ېj�˟����M�(��{�c}͜��5d�J��`�ɃWu� �9�RQ�F�ŤA�dm�T�D+Ȍ������>�d�Hy�TW��f�����{>���N����d�s�`̽-Y�`INj���Q�[�h�L���ȅN3
�9t}8kUd����`�5�b&꡼�I�����QS.y�Is����n=�痘�Lֵ�����$�[0�o5�Ө��Ͱ��ɞ����j���ɷ��P��l�)�6I]��f]$Q��Y�D��;.Eu�9���{B����/����2aUՄɢhU(	#\�=��wo}z����t��߈����իT�キ���j�n��۪SZc"��,��Uue���P��z�r�c9�5�'�B�u���ۋ�׷�l�.�Y�a�3{�๔m8����s;,���{���V�fL{7�j;�ä�}�v��l�&5��c�2v�<}N�MY�E��݊9��2'}�ò{g{�����w�6\�Ǣ����Z�sl;f]ɝ狥y�֙���uoK�Qx�͸Q�v6�T�{~�HW2�p���&�O,8I�ӕ�P�ɘ�≺�K��g�z���gOf�w� ���;���W�<�;�^��H{d���OUމ�� n�e�O�t��N���qB@DH�r%![C�d�qY�l�3v���@�S*gM%1P1d��$��u��Q���y�aҢ�^;��k��>��{���O����������Sy�:�{�)�ȷ)�٘mNT'5�?�������+�&���P�#�w&`��waHB��A:�#���S��C/D��0A���W��7oHع79a��d�(�;�R��!4�M��Ñ�I�i��inj��p�������x߯sf��M��e���D��S��;��N�$��{���2m�}���������U�-�$�WSFw9���rk:r_�V�}��¸�����b�O���?����i����ꃄq��i�3�,4I�Ɋ�NaD� �F�I"�������Y�Y'`d(�z�مquB���,����)F�ETmE#��9p�Vs#sm�Ht�9�jR?����o>�g.^lFdNa��i1g���v'1I�̈e�jHԜN���DB���ZdZU�����w���GB�dD(0MՑ����m?/ruvc�����v�K-�RetTtFݝ�}uF�bb.�Ý5�B����m�;>G٢���eޏ74r=�,�, ��{V{{)ե4��vl�&]�,���Κ�biڳ��ѽ���M�V[�v�m��:�ȟ]������C]�l}��4)x�v�����2+;�܈ܓ��ӭn���;�=l�=[a����|�*�y���&nu���{/.om/q�a�w[��a�{3_h�ഢqIz<)���b$2t<j���w�7v�"Q3F�B�������F�������Wh�\�����o{$a*T(��m\I���̡�oZ�7��9\�<i����K���Cl��U�"��N����7��o3vP�Wfv�G����GF�_�@���KC�6G�s����܇�H3hߗߏ��C��Lҟ�n�~��_�	��!�R�ig��O�����<ycr]fK��K�_}�
��Z������-_�z��mD4�Yc��[sl��9Fcx��Vy��e���	k[K1�@;\�_���+��s4eWD�n~\�SwWK�Z��.H̸�f"0m�cΗ{,�٦��Km����B��ӟ[3�n�
֨�ZH��H�[̓�����SΙ��b�>��V��d���U���S�#}Fq>Z�U2N&�v`�F=	�Z�Y���
@��j��ؾ}��F���N:�,�Tw���)U���	$e�n�H���d>ӹ����E��6E*u���"��-��5�?�����rҒ���e]�;ˋ�Ԋ�ҫ7Z��,XǳI]hݥ%���b���6B�e��ܯ�D�rmx,�7�ц
���MKU�o��3��O��32�nY�7�[�^�+�(]ő3q���8[9(X��U�k�ۢA������O|Kh���ꈕMK�[1Y\�ͣ��͍٨�_[=�>b"�;^#�on=���b�.�t�H�w�����k����@Fbm��N*U�:<@���eqWH�k�#Ī�*�3��?��|�y�볕I�2����uM��@Ԕ8ե���a.14�'��.�[�b3hH7Hq�4佾���z�mc���ו��!�Kv'h�✬��3�����6J�uJୟ#1>Y�a3\y ZK��ĳuHɉ��9$���k(���d���uAD`0�+ZCY�7fV�ţ�����жCBϬ��x� ��vD������R@-����g+��V�� hH`:A���j�����4�!>g�Ƴ1�� ��������@EAs���O��� �?�2�?�L��~'��~���?HEQ����L����}�m�m��m����m��cm��a��"oM�۶�6�t�r�n[m�m�m�l6�m�d6�n�70�n�n[n{�����m��o��Lc�{����{�iPQU4DjO�� m��6ܶۖ�t�p�m�m�m�m��m��6�DCm�e��oM�۶�6�n�p�m�m�m6�o�m�޲�m�m�i�M�N��ζ�6�6�v�T�m���������� �����<�� mĶ�Zm�ݶ�ۦۖ�r�n�nm�m��&e�ް�m����oYm����m����ݿ6�m��m��6�m�{�wwu�a�m�m�NffCm���fŐA�xA��ޮ��}���m�i��vۆ�m�nm�m�m��P�m�e��oXm��m��m��m����m�m�L2�m����m�a��{�www[��m��D��m��m�����,�t�oXm��z�m���[m���m�m�m�D9m�M��ݶ�m���m�:�n�m�-�۶�0ۆ�n�i��x�m��tn�����m�����m6�o+��	ʹ�o-�ۗ�7M��a��m�m�޲�q�m�m�m�M��ݶ�6�v�M���m��6��ۦۖۆ�n�i�������ް�m��32�n[m�"�"������UD�!���/��_�����O�����v,��ҿ��6ۦ6۶�v�o�z��͛;l�j���������n���ƛ=m�ͽv�Jٳfͱ�6�M��m�����|�;x��m�����|���6���v۶����f͛Wn�|�];m�M���f͛m[m��m���J���_�%��j�Ȓ�V�͍�̹/��qQ����v�uE�!<��5xђ�',N����QU8��� �"�v���ڲ�m��n��:F7 ���L��Q�,j�DH�)�L�@��JBU����ϗ{q�]�5�*(�V\�=��Cs��p��12�������G��0���jO�m���u�M�`m:�Fr���3&c*�K\�8��?5r��볶�2�R��G��eu�T��q�t��hH�厊� �9c���C�Z�Tu�2��	{P�s&r'��fTR����k�~�>�Si��G��bh�&"h��@!8��R44�%�X�3r�k�#l��0�B��2�:�2��vՏs�[�M��iT&����+31�����~�s�l�ޒ�����U3�{�C��x ;�����xoq(w��;�����xs�P�xx�������fE_{޿{9�1��w�+
�#A��<"'�儋�6��Ut��X��]4�hѰ��J5�.�{7m����(�6�6�s��W�R�^YKx*V��V>���+���Y���I�����R[)P�7$��I��Z�^�
i��u� �i1���!,p�,Ĩ[Í&�O�ܨdR��wԅ&��,4�b�A#9�F��eQ�ݕ*�Qֱ��0���I!�&��-�o-���:0�1�U|ϗ��]/��7Q:��TB.3�BLp�Rq�	���Z���{2�\�6�-=		0��oH��i�~)k9$m�U>����h�%�%|qR��VQ�tk��؎�����dЈ�6YB���h@�Q�ޤiAM�.��TV\*�IFW[��M�1�$�āG]_]4��j5*g��3 8-�5 �� m9(��P����l$�mƍQ�����k��F3�I��MI�	��M��!5`��U	`_����R��+��CD舛:YC��;����k9�eg&�:���oZi"y#s��UJ7�k5QE�� �Ie��\x��{��N�N:�M%�\9M�n���<M��F'Ƃ�0��~G������Ǎ1�f��）����mWm+$�%���ěo�le�@�x�)���dej���DE7��}�X��r�k	�#�I��h��X!Z>�Y��1��Y%�P�H�-��䅅��Y�����:��A�80��q���/Sm=L��	��!����v��1L�8�J=��+����Do��#�U�ڵZD�isNR=M4'�n���d�!�%���֌˺.��<�2��F)���@GnS��9Zq�\��Za8}��L�5]�%�Tr�.��H�Ձ@�#��UzY�s�I��rP�h�a�A�� �<#��Py��öc�Ut��1�ZXu��;t�>ό*,�n�d�Zm3��݁0�c(}��pJ���"��A�)���z��މ�)�M%�^)�Z���`d �4��Ų�*��Xvm��,��,���,�#	uD�\N�vn�;WGp�n�Y �wwv[r��Nu�`it�N&�`ܐ�k-��*�e0�M!�M8Mg+n3�<�L��jd�R���f䔖��ԑ���Q$��~V�!������_(��)�Ïߖ��Lf�KE1�X�i�ȫJЈ��U#�����F��p����q��D��[1dmZӛin����lP�z�����ư����YJJԪNYH����S�N#WOk���Քc]!�iS���� �Ŝ����������@4?8}����$0�:M��qx�m3]��KQ}��h����H��Ѫ��}?!���`���j����F�za���s �6���D�e,-�`J�`�,��,�Ǐm���V�V�C�����j%D��ʙ^�t��x9s��l���Z�dæ�ϼd�n�{U}5F�&���D���7KE�uY^�V��Et2zI!�E���؜������0RV�Zx4���6N#���c�~_�3K���{_�������X�W�����ұx阼+�	��x`������������8���{^6�3K8~�C���N��D �S�?`�~	��,Oõ�N~�O�	�xp\���I`���W��}�����`��{�$��pO&�Ɖc�D��|(���gptp����8>8M��x�A�^-W��x���{q�^+����D�Tp�@~��S�������g�Wi��T޹�����w�=g��UI�ۺ������JH��Jd]��J��z+��Co��`�;ݔ�"��P,��P�b��Wy7	*z��F��}����>.�J�&��1�A.�ǀ>]�uUR�s���}����USßt(�GwwOUUO|�A$���������ܒ�Gr���������QW�����'�Ye�l������(��YMQ�&���JRdJF�u#Kͥ��9.+`���:�G�իZ�R�w����q�	�V�>HX�����]��$�o�;4�����l7R����X��kR�[�H��/��p��L\=UUD/4Aݶ���V��	U� W�kO�A�u(k�G	��[��Ċx����)@���mF5�U%�T��
>�74��馊ѧ�v|Ye�Y�͵ɍ�`\��m�.�����H�H:|$�ۦJ�1�����QB䉈��	��D�,���.��w4W�7�ZK���!���%��4�)��E3$O1�����XH���!i�� U���N�I
T��-�B$bD}�
v��J|�*� �4J�Ha�ئLBL)`h
)�&��6�`��&R8�
�|(��,[Ylf�'���gU����V�Å�Ye�����,D?	�D�s!��i�7D��$H��/$+g��η��؍���s1������U�)P�)�ݹB��3���bk	�}�q&�eu�,V*H\1��U�2���1)��#�SDR�+�����$��D�2�x�>��B�i�(a��v��)6�"D����H���;�i��iHm#��̜��HlqI����15=�P:b�'w>�'0LS��]�%��ʖh��Tj(��?fb�\�5,d�c	D$�c���Qm����	�#dL�:�/��M��׳Ƚ�.b�����M4�`�4�R�(��EJ7WGV�$�Mk�%Vp��!�Ĥs���%�p�=g��0�"}L��X`g"cԀ{"�"�Г�%J!UTG	�!����	�t�~|��)?X��g(�jQ��0<4��P��p�b`��ދ$F}F����w$H]Q���kF��1Zcf;q��i�q�ߪQx�(��A��W��o��������	!�v�a�'���HU���wUQU��m5���	xO%��c�~"��������le-=�ID�m��N]}$�v�6�"���怭��mC됙z��8��l�xLո�U(����0��f���=6�Xi����i��D�A�P����\ER����tB�a&Z���� �9��F�T��[b��U\����,��_'���l�g��<sJ��|�y9~߫�v���u��Z�ڒ
����͖�3�9%�g�Ip3�؛�`D����U<��~0�;u5u=���ڰ��1��(��mx��6��~[rC��q���F7l+�Q��������2G��%��^���1��d�CP�'q����k���R�>���&"G�V�"�+�e����z��a@��qi~�`�<|�ˀ=�0��9ET�M���D�9��y�&[Op	��p��I�`�Q���W�37<{j�q��}<h��Ŀ^?c��x7�I�������Ce��m�IrOe�i�5�?٘B�a�䞟vP��q6:B�d�|�|Ye�Y��֑�$�jj�5J!��~�O��}�5 �f�W*U˖Y�/R��'BL:vh�G m#���VL�6�TQTI(w�RHC���ȯm��t'�'�७)/Z1�4P:|w�Ѡ/���ƀ�n�?f�J��!!�c���y���
���^y;ug��;L:|�<b�ǆ>q�cNÇ�uQ���|Ǳ��a!�BI��4�N����o�ϓDO&a#-�x#�<Z|�v���5ݚ�v��U\"�n�}Vq�T�g	n��g_BQDq�y����T�4��@�O���|���M%��L"=ʹD��s�6�6R�{)۵a�V8i��ctd���4�)KQ�j���SF]~�]CüN�5�E;RIK�l���X0iV�I]r�,�Jp�|�HƓ	��JnG	\�T�:�0�������FA�}G�{�X�}�����[�1�c��d��f4�k)�z��a7�l�`_(o��K�R����<�D�D����><J�Bl�B$��{^+�Y�q�'�+k��]�2b�j��-^*��V?�xQ�UGL%a	�~4I�/k�q��b�������~_W��d�>|	�G�!���l�{�I��>�3��a����~0�>��d���<v>'ǉ�0|8x�O&����8>��C��x�C�6BxQ�'��Ό���=����p}���Œ�Ɖ��Q�>|>!��|>!��|�>9G���C}��״|o�o75�\5��X����H�k�Ʋ;�Ύ)9����sVࡸ6�m�+�T��KM$�O��nl�*�X�w&�r-�l�X��/.ލM毯{ݡˮ�ʽ�Y���dNǢ���썝��{[(`�6 N����6��脢��w �^WY1���w�gV�W�����R�3ӫnw�Lc���×n�2�l���j���vN�׳\�������m��F� ݃�Xo�����YZ�z��C����}}���ù߄n>�v��_{:L�ڢY��r&��m[˳}���l]�d#�t�2�[sT��FMۢ�,�K5ǚQ33	��
\$���{:�٫SL��N"�;�1路3"�m���V�o{c�ۍ0���2������$�c�ݯ ��;�kɖ�|��_W����N���n<ۻ���ٝN�V���˴��y3�3bz受ن���;����7�pn�Ј5i����7�w(��Td��e�1e�\	�5�
���n[h���e��J!m������^2�m�+ilBۗ�
u2g1��FdCle�LYv����Mؽ����X��52�m#a�-e�GBL�BY�z����6�6�=�ؐ�������\H���뻻�ܒ����Yww|;�$����wwwû�L�wwV]���I3���Yww|;�"χ@K,�<x�B���z2�QDY�F�5n�ĲۊLl~�<9���ԉ�r�+T�[�t٤�j���]�dKv��̺���:߉:?���7��K�jbًQď�}(�<����~���;Gi}���	¿Hɷ/���H��>L�����Jq���Hv������m����M��v�9��� �]$:���;Ge0��/4�5���"}��)�i�[��d�ɀ1��F�8��vڰ��c4�ctg9o�=!q�@�r\�8v�/R�L�����7�$�M����<��P���^@�8l��q7�G4h{h.��4��F�GYM;�4�����.�Զ��髠�&��Io��̣���{3+�*�<.��?h��M�d�����8L�t0!�aZi�vi�lcttyKgub��5�&�㍀<>�3�S���~t�~0e�a������H��O.t��C�NB�f�\������1�h�S�b,Iunp\���p�L��IЪ�t���z�E�z�}M���w)�d�6�Kߎ� �u/)!��Rg����N��fEi$6�XWm1��8��cN��}�Ӫ�Q���qd��'��˺]0K��y1����ci��i ��G�VV.U�.D�M�Uj	u� �+OC�0\�%�X'�suGػ��16��0S`l�I�,4b
O��0�n��H`���Rݦ
���F���[��S�� d�}���0����Fd�3#�cr�??+
�!��!Y��K�������ɹ."�KT��9>�W��9�{��̰ȫl�w, �븝�>q_�45\%��Z��#�6�𣶻T��֫�HL�M5C��HHF/'��4ߒtz��j[�R���m��'�I��]
�4[�!!^v��#��{��N����DJ�y�P�+wvΦ��<lh�l�ܭ�ʕu�Ӯ>�Jl��ơ���0� ��M�u���2����4��P�06ٺ9h�}�Չ,^�<D������JĪ��KK�yvU����[�L��2c�
�N�ad!�����f�f{/_7 �
<4뛣�<� ��TX|j�E��~�QGl���=9�d���ǌ}r|�k���\���}�j"r������O�`F����ҋ���ec]b�V�we�Un�ߡ~�I��x��I!fS�Ą$� ��dC�ӗ���]��n��K�*Q+�<$
�1���m:<au���G������!���C�܁�A6��a㑃���gQ�i�w��X�︟<U�p���K��%�d��%D�8z�����0��nHg�p�/��U%��' �����I�I��"���jV�@�5���7G�V���4>Y�{��nId��x��K<"af�V<ƃ��4��#����J��m�lr����LI!��I�3��tN�H��帉�C������B(�-��@
��D�>Jk��&܋�&�����d$p���0V�<��RV �()6��ױ��;ڪۨ�������z>��h���XV+N�Z|�򊥚��/V6�7b���S�����yY)j��u��g ������·���[��jPV���eYo Q�k���k4��I�(�
X�U��%��B$�"*�]��U�?Q�g*��M8}D��9K�a��&9J�x���j��F�Cn�����f��*�������0�q���1"`�9�W.B��r���z� R`�����$�9X�V�sL��X�d���*��֪��{����+R[Ê���R��aX��*��U�Lu�{�G%BL��ག[�i�.���t��d$i4�)2� �i��FG	�XN�$h�2rI&2��aM&v�Ҕ�t��3�����N���(��!>�[��)�2+�Km3�& �i��&& ᩊ�HU�+�n�A��T�6}����F�(�zC�&&��������W3����cV׋�=����Q��JG��Q<*��&a+L��+���W����lq[^/���:q��-^�����WOG���^�'���#�x�xp|a�Ǒ�8>:OG������>?���x��'�8:<M	��d����<'�<=,�'OG���^�gJ��\չ�L�xW��xa�<>����0|">���P>@��v��Vf�)q����ٚ��ʫ���d|�Rʙ�Z�֭�i�VV���5���iʘi��� �!�k��

ADؐ�ɡ������wwχ�,�wwV]���ȳ���U�w|;�#�����.��wGOwwuV]���<�����o}�9�����Ǆ��K<"Y�Ś�1��v�R��S�ژi:�A��#���*T��m�h���}��j��}��T�J�x� ��ł�R� $�QV�tp�G@>5G(���P���%�6�K"G[�%I��6��ߟ�����ȩ��a��a4|"Y�����s��ml(��h�!:<��:j��N�!�)�O�_͒4�4�R�47GY����K$��B�R�p�ӳ���{_C<{O����y�o>�UIQ4��r0�_u�ND2�� q:��tx��R2d�)�x�XV+M���/�U/�<�H��IV�(�;�M5�:�d��3*R	�G38��=ȳ��7�c-Bq�#�2W$�0���(��s3��L :�I�k+.�v��dm�pA�e�������!O6�=�Z��BF����O�\�J٩!I�¹#)��iEJP��1!��2��!TS*��(���2l�2q�SAKԆ ���J,H�-��rP�,B&��0��Ľ\��ٛ�L��N!UMl��9̄��q<�����r.֭���+
�z�%�"tѠ�2voۭ��_9�e�
/�ĳe�1����#i��-4�/��?S��G����6��e<�3=�y����I>}��E�HŖ�1��m�ĕ�i
��B�7o�3'ϓ�����e�O,�t�p�~����s��u3
�XV+�D� �,>9����ͅ�%|x�X�R��j�BM'��8�]-�"
,j�L�B�9�DI�1�����}��e��g��a���F[4g.4��˒���I�l$�Qo��*HH:GoD�@7�HA<tK!�	��|�W{��n�c52l&)��ˮ�"q6��P����D�����T\%�l�Km��"�����WEJ���(�(�:p�m�v��Kb,)�[��0�G��$6�{���˻�t�<�$w���p��aX���H~ ���=6�}�;��^�������}ڻ�͌��ԙ2
�mz�M8���X�^(�c�վ�{�H��[Uˋ�X7�5��l�FT�7$��,q�� �\K3sS��1շƳI�������)nҒ8Ӵ�t�N}�X�T����Uԭ8H���Hå���e����g0�8�i�d$2�2oԪ�}F��p�<� Ȭ"�tJad�����v�XV+oU�m1�K�Z�n�JR�IQ#R�@�b"e�P���QTQ/F_q>�Lz������prFI���f�^� @��ʽ�S���BKY/+W0L��8BBhw6�7��׉�>����:���>̝ژ�&r2F����ch�׼��G�y:����в�W����Q۵���ZO�|F*�K��������ѱ����R\��w�[.K�Eh�ɧy6Ӄ _�<,����G��-8�t��UUi<��G�HN후�h�-�!��9E^�OE�#o�N�>V��|��1��?w���LP�h\��r���;<ucI�h�'�˔�S�ƪ|T�.H,��4��ce�kO���)C�B<�v@8��� }�\r����o�*�T�@%%�:Y>�M)Ȧ�	q=��5�a��{K��Sd��k�xU�*?����S�	�6:�Ѹ���G�<'��x��t�]�=
'�_O
>�F�S�
���&E0�e���c�Oõ�C�c�<'����pN�����֨�D~�v(�Q������x�}���<|M����yr?���|N�����<a<����:z5���gK�iy�s�������_Ϙ�f��x|O����N����lOZ�x�����q���W��~YW���0Q��8n�y���I]ە����Vث�I�Q&�h��kv���;,��aDKvA��Sb�r5�$���4��i �݊��eC�����݄����{�v�L+�X��{v<ggke������F��1�����k��\�fL�V
��y����7=%����*�X;,��y��scod�k���/��Ф�d�q���x�Ǜr�4k�m���M�4���p�b�j��I2͊=�ۚ4b�tosqd�0����c�2�V��!f`گJL�&�^
��f(ZD����UuX�����,�;��Y�ş6F骩,t�y�J=���
kY1�{�6m���bƠf�l���z���ߓ%~�������[�J�F�J@vl�����&q���]���bT˂�rF�Ke�B�#��g&b�`<�U+�"c�T3��ϵ5LjE#S(�e;g[˹� B3)!B"ҡ�G(E���w�L)�A�]
�6��䙖9,)�:�MLh�V�*����U�g2��V������U���l�{������q<4�wwUe���xi=���Uwwø�{����.�q<0�wwUV]��xa����O4xHCņ��Fr�"˓,ֆ�aH�k�Ф�B�FGktmob\��+�6����
�U�Z�F�#z�\P��=e�S�t�����9�ZB2I�5_���9_�~��$'�ǿ;|�i��&�V����ɴ�ei�Y0dk4Ԫ��y�$#��Q�|���cUԒ�r\��.�!�N�%oLH~�O���mR/ß]]˪*�=
:B�M4`BXw��9��hb��+@��`�>|}��7	)���4��>�y���8�j4ku$$�B�O��i0��2�:N|��2W�J/��f��ld���-�Jն�d�-K��cA��Vx����^y����ʝK�>�Ȓ��j�����1]�����;{��aΓ�`aM��.ݥ��9��[���Ώ�!Ҟ�v��s�]s�����ݕ1�b׮��<�L��$NM�al��-
K�쌗n~��e-;y�rBG���͆NQm�Ǌ^y���#�:���;��Ҙ�yy�Ug����*cL�˜�<�ܳf��b����7YA@���V3���.�E�9��䠾$(;1�	�3mD�j�{��A��&S9f,=�H���u4��z���M� B	a!pC���S�5#A��������Q9XF�B%L|i�X�ڤ��l�7S
5vc�1`�\ɌOj�t��Z���~3g���ڛf�n�ű��$�sy,��B��9ms�"��Lb+
�	i�ru]� �+��}��)�n���X�!����q wJ�u�z�I��h�(�d�8�cf���9�u��{
z~�a�o�9t*��X��X����G3��"����V�OS���8�Q!�����~!�C�e^��Ӊv&@<t���:HBSvZav�(�ۄ�WG!ڪ%CO�wa�Y�4��-��O����C�9>%U�U�-�Z��R���A�w��'�6�Q1�=N1E	]��e2���2QvWL1����j퍱.��~�Hٝi���̭��I�����X.]����m:Hi󤷅[f�hZN����Q�7F�Z�K�k �!U�	T�BYԸ�V \��ag;$�MioE��A�vs�Nc8����b�N!��':O%'��������~��G��=8�1V"C��	SK�w˭q��k���:�ٴ��V�.�B����\Ok�����i}�K�A`���&Ғ��d;I�;�a�S�c�BBy��uy�<4f9>�з?%���NI%��~2�����L1��U�]����l}��X�ʘ�6ݙ��u�fG��S[n�Z��&�S.^kLu�W��"Ź!�]l�X>PM"R7�U�Jj̹9'e]I,��(���Z�*���½���ߝ�}�ȞNXp#�suEV�i4�zI!�˧��!4׋M�$	>�!&���M�}x
�I-1��XK&�0)��O�k���>(��ʻ��]B��*BU��p�&1:J8}��I��� �!����[��֥��U!�TĲm%��џ�zm0�$)n�:��	i���	T�"C�m9`��0Tm1��ש}�8��M:�"}2�*d�r�:e�^�Mof�[U� ��3ϣMIF�O�)8O`2���a6�2s�
q�a��(�
5���G�	�k�	�6:���W���Ç�C	]����
'�
=<@�Q>OÂ����|Bh�C���6?���������5Ӥ��a訞<H'|(�C�xl�<n>'G	��}�ã#���r='��<t�>���	���0�0|?OG���Z��h|6>��<D|���d��:L>=oI��tx�����W�����qq�q�⸼S�"8"|JGD�Q09�~�>l�* �֧�ڌ��Z|�TV'"T��N�l��F�C��r�b�5�H�H7�^���F�5�����{ݙ�E�T�t�p�}Fa�^�[����"(걀�����Fo��a�<��݇�(qJ�&���DM�3	{	�[E�f��t{7L^�Oi�W�>umTϘ��n����>'����˻��O$wwwUU���xa��˾������UU�|;�����UYwø����WX⫏��r���4�O?�6��a*���
��	�	�j�%����^qjϺ�&�,U�+x�+������i�7�� �ȓ����`�0�3��bt�J>9d��������?XeQGxuQ��L�4�1[Uc���\��|gxCƨ�R̀l�de�����L�FN�2l��Hu:���lɠ�ɮ�ae����+	����ܫ��Ɛ����z�l�m�����$�!��v�F�N��vQ��'���y�1���`Mmɣ�'JL{��?d���l1�ҫ*���[�c����E����w���cs)�U�y3
�ֈԓ�(�ds�\1�V���Z Y/s3�����*)dD������3��i�S�fQ��Kp�(UQ���nH�D4��%9y�P>�+�?8JH5�m9��P9��)�D>��$��$�#�+x�?@Q�s�_2��R��1��R�\e|U�YI,p��]��]I���V�˯����Cd�x�Ǌ��L��WA�=����[�0�(��)�4K�ӹwTUSaN�i��c�����h>/�*F~G]ZFf�%�י��#�t���A�`�"�S��G�{���4�����+�$6"~8�B3���6�Wn��@�kWwZ.���I��	e�i��I(��>��·��.�P�R��K&[l�#o�X����Q��(���������%�M�ŧ�g�)����!i�����������b�&��:�Y����+�|��j�<i���Qj_nK�e4r��'+@�k(P����d�G9�Ꚍ�*2�挥�{QGUZ0�w�J�𨨋��j�4�I��A�iI˚�,r��i���HmLM%n��G��b?u0�,y���aڕ�]��ڪ��>�sr�r�Ͳ�l���,�l��nwx�2�#핼Yە��'��c��]MZ�s��9����KN�@�R��g
�&��84גJ���"���V�Gd�Iw5��M��ҽ	LOe9`}����SH����y7�HY��ONB����Ԑ��}�`!�i΁��A����Ĺkue�ѣoԑ�Py(�䓾�m/p��@��+�v��ʯ�y7+�j�Z
�ᇮs$�ܦS @�	���nHh�x��w��b�PD�h8��ñݏd�!���i�>�ؗxí*(���V�FUI�	�����,�A|}���!f��TІ�x�ݷ^V�����B	�4"C���/X�]��6mDD��H\Ui%��v�ﲢ�����j�є09+�	SU����)�X�[�U���~@8�)ә�u0ģM&5C���%$�6���2�y�i0�i�~�324��}^WQ�F)[WJ�?�e�@P�%I*�Sq�!�2H�� %�����5T�%��($5��$ 4����h�����g(�!bp���"�2� [�C8��܏�y�H�a4�~-8ϳTԪ���Ҋy�ו�L5�*ą~�&��?�	�|*�%a	�?���,t_��]�1�^�1�qzmƛWJ��A����G�G¯���||*�&
�A��?e�����'���Wn1�z�/kE��>ZQ��W��6x�6OE<t���0�]�d��x�/������0�&�����9<M��Œ ����x<,�!���<r0�<K��$<A�G��xg�x|h�~pD�*84��Dj��D�xY?
X>�8ՐX�/��N�ރz�뢶Lv��#�K�K���1hTB)�g�U~�7�o�Ǚۄ�o(F� �R� b�Q��:aA��(R2���9��TZ���]�[��������ԏ�M��֩�v�S�ִ�pFTྟ����-Y2�bZC7yBY��\�0�����2�H@��pR�نL1��:��Q7�5�b�7���E����m��m�]Y!4������汢<�(&�fXe��L�u��x�˾���X�ڏeyy]N�*�to��������n5S��WB�u�f^�0�+	{��P��$i���Ǎ�E��f!nm����������ժ�h�ڃ��MU8�:�uc��� ��-u#2d�[kZ� ����{f\�m�H��jg��Rc)�T�'Z���2z��1�u)��k"�%�%m֜�P9�Ø�S��� f>`�>������ꚩ�*���Kj-d��$$�"c�˾ڪ��a�5û����.�w\;������q5���陛���Mu���33�ø�����33}ø��	�<"C�'�ݓr�#SU�%���:��Y����3՚�B��US��e�<j�HUE��GYz�k��7Ԓ��C�6/��qH�è`q��!i��°�8��䅔�yD�J1�C���Xq����F�u�� i8���QEP}�6���9?�B�hiѦ�֮�B�����Y-`��8�<�x�ϖ.+?>���Q�*�ab`��L4v��ބ�#B��ƆCv#�bX�0����)bxل>v�9GO���*�>2�~Q9\�!��u�H0:���H��`H~X�����F���O#q���m�m#���4�L�b�!�!��G��)FH-t��i��I	 ���M4�x#Q����zpy���L05�7����Z�ܱZ������]q?mU!�����O��F�ģ|6����S���Q�3N6���ӎL0�� JM	����*��z�X�U��w^�U*Y�
�Qp2���bi4��O��׿�a�̭�XC2�ѴkF����(�=U�f"��|��mt?{5�}	)!����a��4D��Bi,<1��ٿBB;x�&َ�*�À�>l�ZԐ���k���$ޒ��Jڟ��Ǔ��]y��[l�71<��1c�91#8���x�t�ja�E���j������,��ۍf�|2�/��M+m��t�ԕ�eƷ��s,q��a�;�%���r�ˮwp��)�m�"O�}�QEJ'�&����$)8���L17E2�H��r�3����PK�Cu��z�	����t��g̳��#v[p�ݲI'�o�]�(/ʰ�x����8\>w!S��m����S�o��q���:`�BR[MJ���'!%��8M�,��E*����Գ�i7�e��'�9�Qvr=��
�];M!��G�󛦄�:a$[(���E�d�T�WL+jz��1�>��3O�K⫕��樼l�f�G�S	X$���o�Oh�W�s;%V�9�/�s�������`�)8�UW�d�>m4s@u0G�K2���
<���>:F1��1�`��M�lO�c
ҟ1���UU��Wwf��$��Q ���N6fҢσ���������ۣv�4&Ѻ=t�4RCc�)>N���I���(־�E�'N�������2�2ťؒ>�I����!i�%�DD�,Cx�!�vz|L��q���Uّ���X�o���c{��ప�D����N�+��1ǵU����e����M�U����8���dn�eh�m�Ĳ�~N�j~�&�1�ۚmįbBG)f;Ʌ�YQ��i��I�	���d)�e���u"w�Ws��U�p����9��Ri0u���%�K'HI>���5[mjb	h�Rť���wOt~����I�/Oc�*��Slx�1��s*�Q�qB����2�amHx�.��.K%�Val~)>6�4i��u�RoO}��ە�Fd�h��mYbM,� �r��u�'S"b�&P���}��-
[3��H�)��QJ�����W��m�M��k��o��j�Ep�Ç�zzzzz�|�8ӏ\v�{]��k��Vϛ)�ٶ�cm�m�m�m�lm�lx�M����|��6��;m��ݶ��cm+f͛6Wn�v�Ǐ����mX�͛6l�fa���h� 5�dF�Fj�c�"Vh���T�U䣵���B�sc����}���SV#����R~͋d�r�93X�ˡ��-յB'J�ٍ�*cgd@�P+(-�IL7�vB��w`��]�$e�bw4��W�ER��B�ڛ��Ż@�f�0{�
*�En�a^��>�:�;������i3V���{|vq<�hQ)���Bl��8��s�e$'�&�ff^�|L���陙���L���陙���L���陙���L��ꙙ���L��ꙙ���L�p �a�)�8�1Ǆ��d{��n=�J�^ݚ'Tɧ9$;T*O�m2��m5?&��(�lî��ݜ�z��ي����V^Mӫ|zC���dӔ�Z}��)礓�`�^�#�a5�G��cB[�y�D� C����C�gkzݑ�D;����o=�$��
��p�YƖ�N�p*�2��rJyfP�7:3��ͅ�a�gLq-����&ϰ�4�3�?%�ɴ��a�r�>=�$��N%�=�$�4�,��)�ɗyL�	:���l����#�W�*�d<B���;U�ۑܟ�m� ����k���v�!�X*���8L���UK�AlN�H\�/J̺J:6nil�m��(j��pJ�I�=��%�,A�%�*�������:Q����d+��ֱù �����]Qf�T��G�+�NQ����Ѣ�SB�N$�]�������G�S��擩���h���d6B��x�#c.4i
6�'�Ӈ$�&���n$���xnI!�����3���q1F����y�5;G�X�Ѻ��Q��[A�D�ђ��ou�4���),�t�z�q�]1f0d��CAՆ8����Ǭus,��S���[O9�|Ru6�+�L�s~Z�q���1ˎ(A�-qA��5�$�Ϭ�y!���8M�5l�HJ�ʔK:�)r���t��V,0���;UWl|�1��~�2a�$h�=p��7�BJwc����n�?o��FYK���fhԘp^11U!0�	Dq�d�f���^$�L'S.��h��!8�}#&�n�d���M'�L&Ĥ��	izL<'�v�1ꪽc�1�8��X�eT�@���+>�C��W�6C]�UL�X\UDV�9�/^�$�k�T�0!�̢"
�U�����b�@�����	��2�2`�����|T�5M�7�!�*��F�G��tc�	{Nw�8�>s�$�6u�߳�JMi;٪)�8~8���$�wR�n1�]˘��a��BL�M&��S���4�9FoLߦ���p���pDO�Et��2)���j$�0�A�]�(K0�0�N�I��E8N�_-{&�'�tT��0nHq��u�x�}�\���/��n��Y��[���!i��S�2�%��,�������G��>b��ʿN����0���:B�>�5����]��M���|P��$~�Ve�� -���qk����<�(�3�����,XK�;��6���#����%�_�q=dd�2����f� 5��tψ���|s+���>�u�ȼյ��dS�a�UU�1�x����h:���P��R.�:����i��e\��^�3�z}N��$a>@ۄ��,���O#�4�L�JO�#�˗��}U����n:�<1�����+��nݺm�޶�m�vm�V͛6q��������Ϙ�8�q^��m�v�Jٳi�j�m��t۶�x���|鶞<i�m�����|��6��;x��n�m�ح�6lٵx�m�x��n�m�ح�t��76�x�m�۷�O��i��	�J�NQJ�ͩ�^V��Va`\�+�̑���еM���û+�N��?�;�d�lƪȳ���٧U�&�pY�s�A�;�7S�a���[���l�s����Ϋ�LlW-�SV�ݝ�w'�m{5�f/��L1 J��U����%���\��=��\��c^w&!�W]S�mǹk�n�T�'͹b�ݷ5���+n9d�*�,R�G�;��.���_�kI�7�XfWؠ5-w�˒�>=�6J
�=��hm�b�b�M-�"��;B�����&�e�,>����5�֎W#d}�8a�����h%x�<�F�R��'��޻i���\�\ܤ��Ox����%<1aɮ�\^��.��8��=�ay�}U�\N���T���ƋDIb�K�#
��YN{1�ū���o�<PU�U%�U��;J�ZCY�	5�L鱷����lOR���,P�W1A͘$ݝ���״��0�����	���fIw��fg�p���=��33�ø��=��33�ø��=��33�ø��=��33�ø�����S3�ø���8 p!�<B���l�����nEI�X��'6��t�.�ˮqWn�ih{mR��a�!j��dn^t-�G[*�bfxI|[�]6݂�X���䝓�AQ*�D��G��#�O�:��Y�I	�����~�=w.�U�שlN�mٰ�zHZc�'Ѵ�G��F�D�_�S�=U�Q̺2~��?qa*�J����?ձB���Q�ɤ�i����I�C�c���1�|�QՎY��Y���o�0Ӥ�|�r��Y���������9!�|�_g2�_���z}M����P�n�R����ZD��MW�ta�wR�1:��OQ�s��qZeez�g4l9Hl6@���:B���>�*$J�� �C��x�>��	���8�:���Rۗr]�Q�=S�YD�����~{_�-O�U����˒�L��KN���BꨅHe0�J_;đ�JL����Q��UUy��)��1�c��My8�%�j\�qoÃ�$H5��㓊����w�q5�5��Y��G���2��(巍 �/s����&�`��ip�N���+&>M'\���� I��O��e0�Mc�=L&�>->�M��\�e)�c�Um���|�s1x���'mR��X�ş�ռ��xN�"�I�f�օ1��w�t��Z�mp[n����x�y�є�4F^���, z��3����w���S�Yy���[�+HC��t�@u&f'v�Cɳ�FIiFICi��6�x�1�䭁��H�i�����$#f���?L��I�9e�ݍ����O��U�mյ�Qҟ0�*��=b�6y��\n*��E�K���0o��e4xS���L��G������$ND�4��z=Oy��}B@��aNS��{�����[��L^UwQ���<�!Iig��Z	�S9��%M˅]�1�����<�v�l����vx�x��!����u�$&��ݎ��SD�4t�L��2�d�!$>�l7$~xz��Q������[�H��!Edb
$$<Ԯ��D�F�(�4`1�AQ�e>{�?R|�S�4y�y�d?v�Qt¬8@���8B�_~�Q	%�	[-črI$';��	Vp�r�'��[���.��Z���p�5�4�@�C_L>LQ��-��FR����,�u���2���BB&#�O�OZ�F4��h�cJ�ឌc>g�y����^�e.u�֨7w����[^.SM)�����Q�����0æ�v�����f�hWn������K]GJ�y�lѲ��5��G�.:N���n�3 V 
�cS���ބ��S䴲�(��3;O���HϬ����"d�q�a����Vi=f/��)�^8V.J��1�U�R$�,%�kv��H*=?_��ojY���&��UW�;cl�=ڗE1����:�|����u"e��<rRG=#�/�h����b���(�Ug}E�Ԙ��z�mZm��2w�UIU5�@�Ti�Ӈ�坭[�,l�ƕ���J���[]�m�޶���;6Ҷl�fͶ���||||z�\q�/�x��>m��V͛M�mX�n�m�n�m�筶��m<x��m�����|���6����Wm�i��b�lٳj���Oz��ݴ�M�[6l��m�m4�m�����h������X�t�f������fy�6 L��dK�Ţ���q�}�(VE��\3u�L`�x�u�d_c'��<����ھ�-f^�2"����/����=z-U�ϲ�/'!���ꛋ��;ݾs�&�[���"r�(a�X���/��CԽ4z�G���qж4���Jz��e��ç��wUL�v�ç��wUL�q�ã��wUL�q�ã��wUL�q�ã��;��g������q�⪸��8���&�ZzI8�vѴ�m��{�Q�S���o!sU�e����m%x�:a�q6��yRU*�&⧡���$�k��G�ݼ�G}����;1��T�!�C�r�-�rVr���d���j��}{=ʑ��1F��vFۥFZ����7u �T}���:8i�����KM$a�:l��q4��1�I�@x��d�Y�^�Wt���0Q8 @�D�SM5�|_�����c�.���pf'��8�Mɦ"i.��-��A�S;r$}��̉�|]�择�x�	C3^������ً9[����YJ8�0��ଶ�9l��D�͆j�撔�z�ev���s��+-#<Gf�?_7~�ﹿ�<Z}I����O���iz�Դ����̄�So�bp�k&�#�%��M�O���v܄.YKb��y?cǗY2?F�����6i�舟�C���E��R�~Ҏ�uI�@��A��r�|�:�)Ӥ���<t���rzʬbK+��֬�q�f
�=��w�Kߚ L�}�'�����n��t��IG�5����=�_F��*��;B3ѷ�a�S6>+U��yr[i*���f!��x�Đ��)�ø��l�UA8c���A#7Ow����0��X��6�s��{���
p۠Đd�q<�>��6PPC�"|C�!�Z��6ҔGB*+�T/�],8*ԭ�=�����ݹ�C���Xz�m**Eo�4�0nۻ����ҏ�ن�$����LD���� e/f��0�2�i0�����e]���ah*��c��H CB"~!����Gv�U>��"�p�����^� ��S�ܸA)J((&��}��|n�Q�y���K-(�#c�v���,�iwi�'om��kxW'�Zr���- ���.�N ������h��5�B&N�N�Jۄ�q:�]���&��r�������߼Mf���cB�%�ٖ[SF*�ߓ�u�<�^�{�*��l0�"&�p�!�� �9(1-���֗�)l�{�����z�&���Re�ܧ\Pw�0�����2�̐�&\��	���9!�UQ����v�op�n�̢痨�o��1nfy4t���1�4C�!��]@��k^lwW,&!�i�N� �:��t�o<f�/pKE���l���E����yx�dJ�]�He�c���1����]�F�bn�y}E��}uaв^B�5������ərH��4���u&�]$v���|��%-0�HD����Dߨ����򩫣�n$�����Į��wH�EI%�v|9�%HBx�Hl�6�k:�B���4�! C'0�m:~_���O�$HD���$�I$"��QG��������?�O�>���t���4+DH29���ZSl��#B*��{�@�H�'VI�RE"�)AH�
E�R,
E�%�RLDT�%Id%�%��%DQBQIX���jITEBQbE$QBQd�E�%$XeH�EBQIRJ*E�*�fYFd`���F��Qb�E�-(��Ya�#"��X��b�E�-(��R0Qh�E��Qb�E�-�`��,��,��b�E�,��(��YE�,���T��(����`�E�X��,Qh��E���.U�T�YE�YE�,��QQI,��-(�E�(��,Qe$�E���(��(��QI,Qe(��YE�,��(��(��,�b�(�E�QE���(��,Qe(��(����,��(��X�Ȣ�RKYE�Y��,��,Qb�)%X��,��,QE(�E�IeQb�(�E�X��,Qe��FJ,QR�QE�YE�,��$���X��,QJ,��(��!R�(�E�TQe(����Qe(��YE�YI,��,��(��b���$��(�Qb�"���,T��X�eH��A�$�c$����(��YEE(��)%�(���u��X��J,��(�(�E�(�eQe��ʂ�,QQE�,��(�E�B�QR�X��Qb���*%�,J�c�0dc0cR��R�dQ-*R�X�����ZYKX������K)b�KK�X��Q,R�K�R�,��J�X���T�K�R�,���JX���b�JX���)E))d��Y(�Xk�E,R�K%,R�Y)b�JX�Y(��R�J�X��Y)b�d��Y)b�)QKE���b�)d���,R�K�%�Y)b�JT���)d��Y(�)d��Y)QK%,R�,��Q,R�K�K%*R�K�R��K�R�,�Y)QK%,Q,��K�R�,��K%*R�D�J�X���K�KKK�EJX����U,R�%�Y)b�)d��Y)b�JQD�R�,��K%X�%X�%Q"�$"�����+BE��U��U��U��U����!!!!Ud�*�V*�UV*�UZ��X�Ub��*���b��X�b��b�U���U��b�U��H�`$`$E $`$U`$T`�U`���APd$�TIH���bIH���d�H���P��Y�X�4��4�0�$)H�B�DR*
E�R,�R,�H�#��r���9�����愡4R��4���b ���I�����g�?_�/÷�Cs����劉������~R�W�������� ?�������p2��Hb���	'�������C��O���������Y��?�����)��
/Ӹ�<~*������������h?���

��@��&���������O��1���`���C�����)�	�������t������?�C� Ç���O�O��e��$���-��(~���p���lOܚ���II���b(�@��k[�p?A?bo�5�?��)�fY	 ������(ފU"��YHD�A�F	"e$�2���"��a������»�����ӃaY���w���N��IePIh��U$I*�2bHI%��*	 � �/��������hN?�k��P?����rA��@����|1���Z����sO���QUD��������k�:��;�s���~�d�g�3��a�=����c�����������!�x����!����~u�?���<��g���EU��  3��_�d?�⿷���M�?��_�8 �)�~�����~��E����s�����f�?��k�������|�F;�����*(\�~da��d���	o��F%4���i�;I�Į��ID?�JhO�@���z������ߵ�\�x'�!�  �+�{��!?���#?g�\��*����L��R�?S��~7B�?������y��O��C`����]O�?П�)?P�����3����?������#���?!<�EUD��G����X���W�W�UQ6��~��l������`�����������t?���H0Ȥ ,���� CF0Yb���7_���w���� �_0��܉g��k�\7�p7�~��TM'���C��HS
���O������
 ��~V?�x�����O��)�p$+z0�s�C���ԜD������PP
b��?P쀟�?��'��pPP�?4�Ta��K��oSe'�~�}�S�?�W�!�IT�i�����/���H�
�]@