BZh91AY&SY\W\ݎ߀`q����� ����bC/�           ȑ*D)P�/c@U ��IR	%�D����RH�*UP��%Q)&ڪT	W�I"��]�UEt�APBU
�IQD���U ��D�DDB�"H)�T�*���UR
�R*$���T��� t޵R�� 0��EX ̂*�� ��H�()QDT��$��!T��H��@E)JQ�D�	RT�I*s��RQ*X  �Ҥ =�1�4i��j,U-j��1;�;`�����ՃZ6Ն�[
Y_g \Ұ��ܕE ��v�Q���) YwϪR�5y��{���R�;�]�*��W��*U(�/{Դ�T����J���z9���5J��<�t�*�R����_>�ҕ�'���(I%S��T�UH��"�$)}���;|)B�R���J��+�{6{�D����{��r�AV��;��)Qy��<�R����ǕIU*�Q�z@�ҥW�^g��[�y�D����"E(P*�QO�J����Ҕ���{z=PQ��xz��)�W�zP�����P�)]�{ޯl�����T*T����Ԡ
ޞ���J�U���%R�v��J���f�H �B��) ��}N����S�>���H�Mʂ�]2�N:�J���n:UA�7T�JR��Nt*�%6�[�P)�R�҅+����Z��*�$
�meD�J��|�&��;�ǩ(T.���<)U$Oz����*���J��-��U��U]��T���*q�w
�
�c���U{���l�cA"����@V�U)B�A}� �=����Qw�wG� N�� Ηh:Pp{� �{���p��ڻ� \��� �J�*!"��IT�
���J  �x����V���z�ю��ܮ  [�� ·5J s���8��AC�0�(�TR���RJ�A=��P /<�| �� ��r ��t S�z� y[Ը� 0@ ����;�=p=h�G p��Bƈ��|�����
�}��(x�T� hw/w�����Sp���p g����1� h1�  T�AT)@  �������ɡ�0�4����C���0 �0 �'�
JUC 0��hj��!���i�#C&�F�1��D�U@ �h    D�d�RJ&�5����i�F���S���O��?��g��~��옯�fv��{�FF�gy���<���nUy�}�@Y��( *�(����@@U�N��b�@_�v	�?�����������S����RI$��<U ����EO�D_p�_�������`���`��6���6�-�[�l[`��[�6Ŷ-�m�l[`�2�6�-�l[b�ؑ��m�lضŶ-�m�l؅�m�lŶ�b[؅�m�m4���-�m�lK`���m�L-�LR��b� �1�lKb�!lض�-�[ �%�# �l��m�[�1��-�[ �l��m�[�li�lR�%�`��-�[�[�-�b�-�[�[�lBضŶlZe�
b� �-�m�[�6Č`��-�`��!l��i�[�� ��`�`�-�l`����`� �-�-�[�6ŶĶ%1m�l`��6Ķe�-�l`���m�0-�LKb[�6Ŷ�m�l`[Ŷ�m�l`�ض��Ō`�ؖ�-�lb�clZb[�6��%�m�l�Il`��6���-�l#ضĶ-�m�l[e1-�LKc�ضĶ�-�l�6Ŷ1��`Ŷ-�m�lbS-�L`��6��lK`������-�lb�ض���1-�l`��6��%�m�l`�����%�m�lb[ضĶ�)�Ŧ%�m�l[b[ض��Sش���m�l[b�bF-�m�[ �-�`[## �%�m�lK`��6��-��b[ �%�m�[�6Ƙ���Ŷ-�m�lb�2�6Ŷlض��-�m�l#ض�-�l`�-�F%�b�b��[ ���m�[�lm���`Ŷl[bŌ-�[ض�-�[�#lB��Ŷ�)�[�	l�S �LR�%�[b��1m�l[`��6Ķ-�m�Čb�J`�L`�[؊�J`�� �U� ��V� ��
���Am�-�-�!lKb [ [b+lm�-��Fب�؂��� ؊�ؠ���
�P�"�E�
����`�lV1E�"��V� �@� ��
6�F��cb#lDm����
6�V؂� [b�lm����"F �-�-�U���Vب�[`�lU�
���Fآ�[`�lQm�lAm���� �6��"�[b�lUm����(��V�*�[clc`�lb+lm��lAc��A� ��@��� �(6�V�"�[`�6�V؂�ت�blAm�-�E� ���[b�lb�lEKb�[[`)LV؂�[b+lPblm��P-��� -�6��؂�[b"[[`��-�m�lŶ%�m�l`�ضĶ%�1-�l`�ضĶ�m��#�6���m�lb[ض��-�`�)�lb���b�ضĶ4Ķ1m�l[b����1�l��m�lb[1�%�m�l`�ؖ�-�l#�6Ŷ-�`��Ŷ6�0m�l[`�ض��-�-�c�6Ķ�-�lK`��6�1��m�lKb��6��%��m�lb[�6��%�m�l�Klb[ؖ��%�m�lcLm�L[b[�6Ŷ%�m�`[�6Ŷ-�b����ؔŶ%�m�l[b��6Ƙ6��4�����������|۹vd���v�����E��L{(�Z�`�[�T�3��sX���V�m�m�9j��P��7�ɻ��$�	��QuN�*������Ϊǒ�`�"Xd\�a[w(XKU:�+0��.\yvq�t
��R�n6nfQ:�'Z��ۡ`#H`�l�[yxĨ�tģ�]�D
Ƶ�te�T� [�L�Z��32���L�q��oih1U�hmj�m�Mh��9��D<9n�a۲c�1��m��
�T$[��kئib:��+����/!2�B������u�ٓT��d���B��"�nmbt�i�����$p��.��L)��.��Xo����!B���*^�1س��[�h����6�(̷M[���0kL7[� Q*�`ڕ]ǫqf�]o�/Q�-�����+��n)��&�׌Zp���D�ɿ*�7b[D�ef멗�c\&����i�G�μsUڠ_Qs4,.�լ!="�K�*3%�&4�f�͔E]v,GYS�x�L׮�[��]Zb�)�nQ��l�f]�B�]d9[JzЖc�{CjQ�y�U���ג�(��u��um:I�Q0�r0�%y���V�ð�*�S�h|剪mm����M���P�f�m��L�lѢ�e�5�2��¢@*�=���4/-'�ʨ�5 J��dzɆ�1ep���rcY{zʩoF����Oa�[��iJC�e�e�W�����ڦ���Ջ����,i�Y2���ʐ�acj�n��X��v@�ЊQРm�
`�ҳ`ӵR\,�s.�
��S��8m7q�ݠVm����&���/ژ�6*����4ʗPM�ڏV8�:�7b�HY�I	Lm[;��n��q^��b^ l�K-�o\2����kap0To ��sA�
���f�,����,\�.�[��y�Z�X*��C�ܘAE�xNاB��C!�[�f�4��	Y��=�l�����Po���˴a��`��ְ��k,ݪ0�l�J�T]rl��# ʺ�]�C^,"�X ��B��)[�Ř��r��1j�F̐\��4c)kx�b*�6]u�r�E*ɻA�=ܤ��ò�1��f�K[�E�	�MX���.n�
y[j��ݡI���k���apR�z�fnËY�X�@��[���"��U]	��:"�fPEVم]a�x.=R�OJ��ZYe�ӄMZ�HkʦVU���k�*�U��A���)�^.�V`\��R�I��S�\�F޲e���hܙ	Wo�ZAN=�f,Ra�W���i1eZ�fZU��8��0��|[
WW��iohZ't*ú�ZE����{X�ѥ���J���˗�mE�,�U�n�H�wMdt�Rw�GS0�u^���82�[��:�9*�nЬV���6��́��$��$R5a��X�V=Cb,n;����ڭ4t��[/�!b����E5��$���wl"F������[z%ݸhA�m9�`#�5MKY�{u2��k�Z�Vk�kHV!���3180���U
�$�T!�7-�НG� b��=��,YZ��0�%!(��s�J�,��,V�ڨ�Րc���nS�����f�0��1�����nYU5<n�b92%v�6�k�a��N��e�8�,�7Bj�X2�:�J�������Um+�4^Ԫ�oE�H]4F䢱�۞�q����JO7Z���v��N�[
c��[H���G�&FMm8f�M,f�C"���[KF�a�fM�g�[R��ڢr�m:�hǶ4��P�����0@;%đ�Iң�`5�#��1^�3Jt�h��TY�-������P�R˧eɫT8���CyCC��^&d�(��.�4}h<� ���CZ�6�y)�A5f��ْ� ��Y[��R��ԛ�H�W0ݩ3B��Iǭa�Utݡ��ڎ���7Y���Wp1O�۩�&ef��,Y�7yRC ��lF��MŸ�R�Y+-��6���	�L���E]kԳ�r���Z/kBܐV�0�pE�7G�55Z��vҕ�fn^³�=���6
ź�3�ݷ6�ZP`eݡIK*+�Ve]#�@��0<��ʎ��ng$jcK�Z���L�E1�R�&�Kr���nl�tu�櫻���/DД��E,�V�3ɪ"񵦀xX0�v�(&�����$*WV6�csQ~I����A�okm3P\�h\�G/k%��e��JɆ�,,�sP��OP٠��Ij�� 7.��ҧ�E3!RlX��ۚ`ڵ	�Қ$�G�3.�E�X8l�gř+0�x.�^6&�d�
��H���,���R�\��է3w|��Rcv�a yr����LZ��{�<��iD޼QX$KVc�/^J�4e��i�Y���(�p�"��x-��%.
slYz��K��|MZ
�a	V���G9��Z6��? 4��5����ݥ�[�P������#�����ݛoF'I�rhɈ^�kX�l�M^�ߴ7{*zE5�aҠ�Ps�L�������F�4�,���;HHR�p�P��4i��<53e����˂Dŋu���p9����[g!sb�Ql�v5km�`����`3d�v�׸�X�#Oj�	���+tql��Q@1&Գ0�)]�ڽ�(,��8"��Ay�J�K@�7,'t:��&=7,��nd�O6 BS��䱇L��q=���X�(�9r����[���]Kf�M���Ʈn��-�
�їLFi���5uo֢�˒�کY�YDаq��n�,^�5H�D�S.�x�(����Ve�q��)��3T�1���F@Ţ*�yw���(�!S{D�M�"J�f���izi���%;/�������ͭN�D���$�؏�`:^����f+���e=J)�$��5�e��������*�u��ea�M:i<
�t-^�R�V�(�$֘Ԇ]iEL�0��f&���ȳ�c�U�e+vP ��E���+^��y5^��0�Ť!O�mG�t��APJ�^�,At�\�WXX�K̫۬�m\��
�6��D+���v��t�u%-��n6n�U�%�ͼG2�B�L�b�<�\b�Nֳ�;�ZnMӨ��$�f,��[�Y�.d-�fy�c"������B��/�TRK�a�j�	�|%˕�^Ռ�QN�kj5$�qMg�9/h��8or�'�%A��L1��\i:SDs�zˤkf��ua'Y�!�^Qm�nƂ����-ie�p��{v��[Fx&��y1���I{��%koI[ChB-��90�aV�d�45R���*&�`��A��{��2��R�40�kl�`�S�^2%i�D��Cwiڷ���tM��Vˇjí��gv������t1�� �������,�"�XtT�c�cp=���j������2&՞�����B�n����v̒ݜ������]�qe�2l�{VL
��*���SM4�㘩�i&٥���وe-`��QV��L�Uq���:�������Y+ x�&� �2�%ZSӒ8�]քu�ݹW����m$5֗��LR�֪Z6$�=����c�2=�퍑�q)�8��DB�-L��z4;�a+eӖ�`1�b���r�,G�q*�${�@���Kj���$�J�G8�F�����ɝ�T.P�1�Z��+ZM����[+p՝WN��
�.܌����]���ݸ���hӶ�%J��M�W�t�LF�۴�S��2߶�D��6Jz��fl7+�U��we��`�X���4)70]޼o�l�+p*�s�p����a�R�pـH�nɦ�C׊�͊�6�M�n��(eL;��we�Z@#K[���ɔ��)He���q�,�ݤoG��M���eZx�
��6l[��,vn1H�X�*�X2�=��F����E�[z^)���`��Q�����w�6�Xm����w4��%	A��j
y�ަ�lԥ�p�HA3�R��Y۲��+n�rY�d��
�wtjm����Fj
� [���۳I��~S+Gk���dkm���f�e�R�w��ܫ�'j�+��6�7z��n�b�Y5�
y�U��ʱ��6�Ēn�q�6�Qu�)�Jט��`���a9�te��b9Ocr�͙�䢮��Y�G,"#���#m�a����[e~p�U�u,0X��.�¨�D�7�5ڨ�en;�pP�T&V��̼��tŁ�P�ظ%&�%a+5�a%M���Q�ǆL;P2��h��e곧&�u
��
)�kjQ�5��h]�ܛJ��B�+���&`f	������m�fȩ�O,�J�*�v�赴f[�!d���`�c�AȈ���Gt�Дu�Z�j\�A�-�cuQ#�B��Çie����M0й4@�l��<�uu�6LJ� �["&���fc6���I����&7YG�Ⳅ��ں�nnY	5'F呷2���Q�D��I�Ce�N�zˡ�ŢK0S�]�R�@��m�v�k.%v��:s�,��a�I �#I�Q �=؛W@�FֻYxkc �@�MSM���̩I� ^,۠���B���N�:\u��Ф�X�f�x�$b9Q�"]n�5*������R
��y�][4�Ws�&,���܂\U@3���W���j�57���gu0��ͻ�Ok.R���.�RsI�p��HVĊ9u�c���Ի	<�n𩌛Q��o(nҚ)�a�TB����e]À*5fA��5R)b`�z�5nXZ�.�j�k̫w��YE���R��7j�LWR�W��*�YX�CJMI���ɢ$op(j��:T5��E��ң��E]LVZ������R�F��KT\��b�xQ�l��Rz�VhZ��43]jԕh�*m⤈7�=W�X����mjݙ�A��M�Z&^6;�w&8��ʙ�qJ.�<U=˙.��w��GF��7Ȣ��V5&jJ[h��(�	v�Ryt�l5�,�Nݕ'^��ݲnnưР�ڷ��Jk�t��y��MMu.�r�kRզ�ًڱS�VުD5�ȫeS�Y��i��X�T�ӌR0��]"��s/pH�5�hSy�%12+Xݷw��GY[2("�ۣ!R�mj����B�U�D�ѭ:77"��f�}�{�D9q����S[�m;����nͅ��hG�u��bŕx��֬"�0���wV n�DU�R���]-yJ�d��)�d��$A|�0�
K�E��1�1z���.Z;B�E�r�e�ŉH5�S��t�[K3|b��ɶ`E0t�'� 	-�+mɕ�FZdM�ʧ���!g�ee��ڬfY���ˑ��@��:K��ZU����I����Sw�@�� i�֒T���T��ۊ�c� �ڔC��`�5onS��u7`�EJQ܉I�7@ZgP�I`�)][�XѺ�Ww1�Zr ��s5iL	��H%���Fx�Bլ�iJ�n[�xh��ݰ��� Iw���R�or�Gi�ٹ2XɵXO&�#�0!�+�y��)@"l���S�bN�%��[X�!*W�bA�Z*%����ť	�q�ąe���l
RlX5���-���u�����ɐ�ec����H�A4kq�����m=n���;�C؛`�3nf�G��Ä0(�q���˘�t���DRY��b��F=�ּU��c[2�:�޲1�^�1��ad��1LX�,x+*VʺD3p�+7E��gw���6�]'j�g+����ø#KI�p�g�:
-z�Ūd����q=p�y�"-1�+J�	���a�Ԗ��ÂEZ-m̺��X1���y+!�(;��T�B�哄���.�Z%i|���füU��qǞ3�����h#<��L=����+���S�u�YZwA��ä�E���DWm���U�A«a��(d6KǕ���힠8�d��K/~���X��}��'p�f�a�v_�2p��]gH����Gt�=�Y��m���A#�=�.�oM����&�ݫK��(�d���_�ދr$B���hr�=�{fae�(-.�a��!�Y(�EC8�]�P�	�f哆q$ޞ%qnʲQ�o���.��ٶ]��qZr���N��d�p�����1��:d%����x�di�8L�	,�;@i�u	�I6m��"�!�k_hޓ�YP�!���r��+�C���8�1N�41�OBy�x�Q(�WN�t.�]ѱ�Z�#yY���l�Y-жʡ�*ΓP�2�$"a�{3�:i@	��Ų!�.�Ys"Ӥ�{��P���&"�l�v�$��l�l��"Y6E���˹����3m�w�3�n��e
Rdi4�t.˲S{��W����e�!��gE�xOȲ��F췃/]�\Ƹ�%g�Μ3oMG��7���	�,�&��se7dЈ�Q.���jק�F�g����8���McTk�K4\DA�]���M��yBY�.����oIga0�,���-�@q$�I'�B��-��������9Ǩu�L�V���n��g�w�iU�	D�,�:IG8�{���:U�f34�9��P����V�^o�v�&�<a;�(<�y%�f2I8D+��ώ�l�O3	���'I0�f��e���.�����s�͗���d��0����&u�l��)pLE�ah�:�U��p�&�F�¬�oJ�\}51�j&�h�΢ZR+	�0�r	'�i)��ׇ	�h�{���c��*f7t8d=f�{��(�n�;&�;��y���xp�k��9	���0��ɶl��a��o6Y-�K-�f����3�qe��b(���2�'�P�m�G�����1��_�� �3��D��,��Re�_3_f��gQ���h�+G����9�ޕL"IM��������g�E$��=��������+�0���&���7�7t�wv�Y�؜�-�ݘ���P�w9a����X�כ24�,�2��<��܋��EWf���;�J�v�V��_/%�$�Jb��t�\�oVm���������"0+Rvk]Z�[T�`�Z���=,�B��z]�74
�%LlˆgeOw\k�3��8����td�����ٽ6 �v�i�dؖ�Wo���Cm:Wo7]-9��W�}�a_4$y���ɀ���O��ǝ	[Q2�R��o:���G�e�]B��t\Jw\�\Թξjf>~�$�4����]LS�s�e���Πt�F*��#%e3:p��] ���V0v&�31�6II1�@L�p�W�mw'��1�U�}D�f/,�|����g���l�ml���@
ܜ(��Ȇt��3�fwp�nئa5kw5�c2���p�vȢ��h�D"FY/��Ӻ�gu+�n�Mp�h�8�iZ
��)�)|M��g`	g��kYW;i�#���=�g5N���������K��t�v�x��~�F"s���n�k+rQ0��(�"zBQq����+pI��{{{���\�0p�3&��5SSW��M��d=a�ל�l]��r��������Df�t�b�r�K|�p�&��Tx%(W\J��!"����>�A���V�h�4ڙӷ9a��u�G�"���'V� ����Ɣ���:��̔���ީ��a�%��}�[����f�d�6���te��m�N���R)�S�汀V䷋�1ڵ��ZԴv^s�Ƿ��[��.���7���V��S|!p���V�5[E���eof�W(n�b��:>m2������4	H��;�ω��Cw��o��]��
�ǝ��뻝%:Q���oPN��%ْ���d^r�C,��1��q0f���D�>��
��#gV�;��R����]F�s����;B������f�*"��vG��w%ʸwb�E(#WJWS�;U����ʹe�}m�M�L�|�!ՙ�_Yו:^T�Nf�@�q�Y��5m��V�n:��aU�� �V�Η�q_\p�4���ބU��(�fYۮ����+�
v�^9.W�i��fd1��	�e]j���>&s"
6׎��%i��u��_d����Sr��̔��l��6&>�m�OWi�����f��3
��]�w�m���+���J�iܒ��w8h��M����r��ۮU��y����;P�N�
�.�Ij҇�E�ܵ+F�UA@�w����e3յu���4u;������vw#D3�Q������)B�)M�j��d�o5c�'d���q,�fpe�OaNBf����Ů�X5�s�]�ȡ� �vf`�ׂ��M"x����n�g+�t��յ�-�S9�d��KM"�fhY�t�ve1洐�K�֨t��w��l�ɓ��9�����Lr�:�YWPi�<R�M�%��#3(�s
��B1�/L׭�.r\�ʹ��h@fs�&M��r�M��3p���{`R̞�	��ҟw#1#Wk�<���[��C��G�2���cd�����t��f�қ��ǹ�ڥWݔfT9!*#W��g���w�ԗC:���%_5ًv��-�c2�U�6��F.���m��H��6*<����l��;�I[�፭�߯c7�H�;w�����n����1#��)�L�\nqg0����b:I5v�Z�.N1t��;x:��+��n(�O�)�E&B�����i�x�mi���!I7����&@^7]i���p��	��]`*�)��--�{l��Ս&ާ�$g�XT"�f5o�g\�Y�]fә])��wnT�<`�i�����!�R���mc����Q�0�	\��sE�bZ��ΰ��7�J�g[�8#�Zs^<�c)\��HDjp����,����I���/����f��8��zr�7Wx��Y4��s�X��ҹ�њ���K�O���g��f�F�3Y���d��5t��3[L*���:��ˮ�n�(��j*�5l�+2Ն:�v�yR�qcsg],d��;�+`�x�T�Y�9��u���̆�<�Bn�!7��n�wY��O$�\Gq����U^\���NC姹�p��
;�Eַ�{�e,f�7����m��Q��P#���ү�ز���<6�>Bw`uZ�{3괰<-��8�2�v�n	���N,�J)����=A���^F�V8�L�lNe^j�d�Î�!�B �}R�:��2&�Xӕs!�0 �d!u�i��F�Ń;^*���^�jj���S��7�W51F�O9���5D�t�o����V)(�j{.�G��l{��x�0!�ՠ����;Y���w����8�ts�;H�B�W�Y�G��K��8����`�xV���5PŀuNꑒ�as�U�C��ٲl�1%q�^�ߦ�_ye}�﯋�����.��!�o�6�;ֹ^��:H��4�j�bO�@ȥ�m�`L�Vm�̡�ύ(7�թW��F��ʯ+���L��+��,�T�k�:���k�LQ3��=)���m:�vv=��r�5L��ٮ�&*Q�z�^j����ѓ0�J��u��H��iCh7�[}�=(�Z���q�Q��ttj����2҇��}yF�qu� buŚR�a�.ޖ�ض��gmk[Ǥ5�ŭi���͹�#�\�"ٗ�0ZF�.���%Dg@-�D/�mhᷚ����>N��gJ����X�NK�R���BǕ�_Mmt���-#I�^���c�e��G(Si,�[�骠��Tκ�i���W g'|�����C�7��yW�݂^ɉIy������ԍ�k��(Ѯ�W��;�vT�N�7��-In���۫�OU�F�>c��l��6�u��.	�"���/aȎ�و8�G�V�;��	i³V�dv���g=��[����SY�E՛���r���,QN-��.�sX�:�[�h�?���ȏ�@Fm���S�Dg3:�&;v�hT�m�������x�V�U��n��l�2�:���f
 7$��.N��V��Iof �{c�]k�7��6�TVK�H�\k;��G���8���X���z�mu���#(F44/4�󻻋j�y̝H_4���;��u4|4�[��-����Y�ʕ�AKd:��sU{ �G+������;�
̧ի��7xt�k�]+��V��=�.������`XV�W�F�{��i���&��A�k�b�m�G��.�͖�����AB����I�,�t�0�$ޓ�u�� ߹���8W�Ck9�R:Ϣ��wZu[w��8Jȋ}�Q�X;�C�YR��ζCJ�ӑ����5t�L�t���K�Z�r�t�Wi��^AN3!�3t.��Ly̸78:6S��;r��"E\E��M��{�MB;�2*��TZ���5�L�� vK��]uI��V�-�H!G}���(B�J�f���:���j�I�����&=�@�*�?bgYY<+�!�=7�{y&�e���t��w������tK���1�s��w]Z�r�v�M��8�ڄ�6�����V�:���wB了ش�h4RM��}]\9#0�\{jas�:�r̰�>��:�q�:Dƻ�f�D����Ņ��t�(�`G�ua�.�Eܝ�a�A��uK[fS�h�㽣ԆB�o[׽f��%W���Fk�<$�g)N�A�88@��v^�B��K��Lbpe^b�ϰp����v�ȲGG���.ۊ!��8���w�s�i�LvVf���i:��OIW�Gn�+��`:�b[D�:}�cG���\�"���ۼ�ۣ-t`rN��W)��Ô��4K�ɵ�v%�ؐ�{�U6�]��rfXXRg�d�]��e"�n۠�)�G��9t.#X���3�Ytz뵝��\:�nS�R��'��0ĭ
��a�zd����]]=�iGr�us���)i4�RND�7���m����Р���v���>8Nd-�N��7���T��c3m�k���!�\��"�ܵȕ�£�z\�l	���o"w{&�E�S��!��6�۫�\��>i�7�.��U��ժ��냚t�"�l��8���b��[J���0�F�[a3Y-ҳ����S�k�p=;'R ��ѧTy�u��O7�:4�A�Ɇ]u���̏k6>4@�rTp�fˡӲ�I��`5]��J't�^S2�R��w]oL;׊=�Q�d���vG��ĩ�ϰ�:mb�Pɺ���v��Qn�}�f��#-���аc�:��S<&����Y���[��Q�ʁ'���YW�-[�^�)�#���;*'��vA�n�kT!'%-w��q�*[������3��^
���GE�i��[�l���pB�Pi�csg��#�%Y{F����(�lڶ��r��ՠ*oe�ն�|^ �"��;�yp=�Gq5s�/���Os9�#��5�ܹ����M��0�����M������p`��mJ��]'�`�W��:�ةM�b��$;]�c��9쒝���v����WZ�6�D��镠�y��Fp��\c$e�/<7a�.�.����2����u����y�.�b�ƀ���:ãx�v�@�F�s�(���*
�յ;M^��x hgg���d�����u�\�I]}E $�]��C�Ė��#���m�y��;U�i2�I��]��I\��iåu�� �0��'r��%5�}���u;ޱc��0��1:��AK��YB�r��&��Q�	Ɵ;t�v�:(��uwږ��
�G��&�}~����:Z���֢�㜶�:���r�f��ᗵk��i�v@q���#����P[��kS׾g�����:Ý}Ό��x)e�%�ẖ�W�s��������[,�0��k�,t2�wp�G��AMiZ̷ �Y���x_�P�y�^m��9�]���'>�7�p��.��wf���1/�8��L��g��_r[�����-���<ò5$�ֺ��/}{������m�̳�W�]��X�4�6�n����͎�,zyj�l�@5�ݤ�.�ꜙdznX��׷��]d�Ar|�뤻+c�֎�\�����f�3P�R�WWW���;�pV�7���wir���1�`ru��/�
��.�!��9��ܱ�eH���Ӽ�wL��*�ԔT�ͫ|�Z��kZe<�ټ�r/+wJ�T�Q٢�g��f���	�&�;I]�ᯢ<��8�p�4�!��v��x/��p��iu�}�8G��cL6��5���';� �Yok*�7��n`��:&Pv�wǅ�ӢSG�nҜ��i�̲Qz��"��k�η]F/�N,[IX`Q�)���m�*�����.��Z�/jAe�)u�D\7b=�z�in�J�ǅ�:�m��w%�Gf�
��Tb�Q"�vۙt�t�J�P��`�-5�����O��E�1a��s.�v��Fw�Y���N�mY�u�Z)��p�9E�������n��4s�_Y���\�D��o�aŃ2�C�Ө�(&��^��;Z/�3OT���G��UD%|{�{Rw��,���J0fu�}ճ{��o_$2�o�5̘����aˣ�%*9Q)!|�s��"��i�Y�o9QYw�c��!�㗃�:c�r>�]��S��qw6	�����v�\���E�C��!�Ѯ��Һ�/��e6Q�eu�T� �ge*T%�*ʧ�e<{׳[�y�V97�o��q�u�}I[�=�F4���E���;}�����g��Wùv�c�ډd�S�8���h��㔱釶��B=�1�@�u�V�n�N�s�WR��a��y���,�CΊ��b�d���l�.�&��kI$�����L��I$��3&^���Ԝ��ij��}��
^�3��TFX��:�h��ѯ]g)�WJ���f6y�s��BZ}�X��*���-WU^�7�{.L����`=���P���nv �eUQ<&o�A7tv
ԯh� \�kܯf���(� \�o{�
k��5�]��pCSsQ==޴j�����P>Mr��jr,�YC�&��A�&����ީ�N]	�)/�Ƣj�����g�<������E�P�בG�y7�y�"��V�)W��|���U�(M5�����y�O����U@M'·Y�++­Mr��P%�v'5wQnq{Jd���"�����K�j9n�ȷ����N��5*j	�]�`���Ը�{Z��T�*o̽@���?���DPT>���ϭ���?p�(
?�����>�����g������Eo�0�f����rb�H)���ck�ܹ�H.�<���	���٭D�b�j���oFg<�ꉪ>r*)v�B�"��d����_Τv��"f>�7Y�X9��;H4F�v����[a����
�����t�.�.��53h��vTW��;���"�/2�C�2]���|\գ�l�*���W&s��ּ9X��!]��*�s�����'S�ݔ4�<�zX�t�'�En�^a��Q��j�y�Pr�����Ej�OWC��.m�5����J:Vib�Y-������K���!�A봵42�k3+9E`{KR�
��ab�2�wza�Y�ە�A�r�dv�2�%�Mb�MX�k%�r�nѱ0�S� �hA�vY��hB;k�ot*@��~V+��7<�[u�p��y2j���Im>1�elU*�eJ��׽�O8�^s`�o�f��硝wg��J��:�Q�Z��U�u:
�{R�mb����P��[��
Z�-����0��|��U7M�%O�+F��M�;��)齒���]G9nwf�R���!�=��_vb(��ĹV7
���Z"��ty��D0O+��{=��8㏎8�:q�q�qƜ}pq�}q�\q�q��q�qۃ�8�8�c�8�8��4�8�;q�q�q��q�N8�8��q��iӎ8��>��q�qǎ8ӎ8㏎8�:ppq�c�8�8��q�q�pq�q�q�:t�ӧq�q�q���8�8��i�q�}pq�q�q�q�q�8�q�q�Ʒ�!%��a��s;�P�T�W[���ł�J���7Y�S5}�㺀�<i��mQ�YP�t��K��R�A-�:�˳���ҏ��6����!I���o\�T�{ht�囻��B�B%��!��4�����a��X���v��x7��Īt������X!��ay�
�Ig���mgwk2�]1n�����y��Ά�0*pj�&�7��e	�m7��ҍܩ:��ݣ�ݡ���XʼUz���˾�(:M��BKI�u}��<s
K�l������0iUy4ܳ�9W*�I������-�^�-O3�e����
����G�%be^L�8t�ļ�,E�N*�[[�3K�n=�2�=ʔ���賷8��Ł\�.��Q�R���5/r���D�r��u s8�|)f����G1mtӸ�M=&g#D�<��ရb´Ѯ�t��=����;n�b�J�K�vR����*����.�D�;MS�+0fG'
]�k�6�@�ҧQq�ʓ����w�j�ҏ��'�b��0w-n��H3�j?
�vC�x�Xh9�UC�_=��j��&��с��u���+���m3�8 ��;|�V�Xlu�Z��|�-�9��vtͭt��I�Jk�zz���������㍸�8�q��q�q�q���q�v�|q�N6�8��q�8�8�q�q�q��q�q��q�q�q�q�q��㍸�6�8��q�qێ8ێ1�8�8��8㎜q�q�q�n8㍸�8����:i�q�8�>8�8��8�q�q�t�4�8�>��8�8㏮8�q�j�3�'���nry��!�dy� CGuᏄ8�^a��e�4�l����t���W4:����0�u�J;���#X�P+p���շ�{��˻�"�B�qon��'.���R�:�L�U�^ҍ]�V�7�y[}BGIƶ�;�)��������N��lփ�W�W��oO0$�{@S�*�'2L��.���R`�a܇b`��T;}vj���A*<̫������5؎�ѽs k�U������0��XqJ\�G�V��}�o]��zꯂ��1ݘN�y�e�ST񝾎1s�SgT�x�[]���w�M�A|f��Nv݈���+�ݩ�'2���ɏ]�٩4����*�]�+���=x��7;-�{��[�,�ƢW��O����롹;r��c/qD�3g8V�)Zv3�)�C����e��6�T0���o�\E�,�yl�-b��&X�M�c����8�qڒٙ��Yh�\WA� У�p7gOn��2�g3r^������Mc�2&��!�����cP=:����d�A�1.Q�$+U�Z-��9{g�
wV֘��}�l��z�H�T�6)u����-����u,�.�+,�6��̣�lqC*�<�������I���3�Vѱ`'���Fkw����V$������㷏q�88�8�>��N8�8��q���8�8�q�q��㍸�8��8�q��q�q��c�8�8��q�q�q���q�qǎ1�q�v�6�4�8�xӎ1�c�8�8��4�8�;q�q�q��㍾>>>>88�8�8��8�8�8ノ8�8��4�8�;q�q�q�N8㏎8㍸�7Z�z_�߹|c��
y���Tɶ�,in4���9�L�̦-�=9!j�Gb,cn����$���U�x%A�4K�ڻ����T�����F�BJ�}9)-�y�`b��u
���ǃf2�����.�F�v�mS�,�t�_m�'�V���n�����}+E��W޺9��t�lu���u¯�NK�Vi�w��[puއrG��=waR5����nI������)�N���6ңn���� 9�Ix�f�Π �0
�����vD�̃���	�r.���KL��y��T�KdtS�S6�ѩ;Iot�Y�8��ܡB�X��YW2�.E�v��`-kF_Y�*1-������AƲ�]**������ed�EB
�5�#�h�w׼�e�u��e��i�?UU!^ƠR����R�1���7�W{n�M�J&�\����j�9D�MZ��6ޒ�<��Yb�7aq��Z�%⎥�t�U�=蚔l\�|�L������6��:f�m2�;�W����u��"�V��7���ac�Hj^���X4�����Q?B�A[�y��.�y2)}/�n��.�yqS"�6��u���^3�^�:|+6M6Y�ƨ3.��*Ѻ~���͊X�ػ"q�[b�$���C��T����eJ��ژ�a�eڻ���+(�÷���uîv��v�uy���,�hc��T��ʺ�!E�-��� �zڮam�t�h9�*�5R�V�{��$�%i;�'Z��uڔ[T�0^=�v�KZ�;+;}�UvD�]-�f���M	���V��/��Wet̺
��;�n^�V}�;�j�ˤۈ�Rjl��9�n��x�z[����#̎<��|��vwV�5`�܁\�����%M�j�Z����cx���ٽ������2�u��RA�)i�6��u��Z/�sԃ
��"���Un�1J�����{m�|�5�79Z��9N�1��!Yk/w��r���T�Gfr�Q驘��z>:�E�;�(��xUM�6��f^l=1�*�]��z�"zvX�󚧤0ǵ�bz'xֹ]�3,��h�⵩��|��u�k�V���G��H㬻h�୴��$$4�U�.%jɓ�Z] ����q�{k*�LI}J�^����T��T��9��}�{v��.Ըu֝�W���9͋h�Σ����vJK�)��~�W�xҗ!R%�F�b���U�o+Rc뽎��n��v��-0Ҳfm�54@MmF�A:6�u���㢭�$�mI��A�*�'jW��N�Z١{i��>�zp��w>�X��E�
����j��,
�z0:�N�z���y����Btᖕi��gv�W�*ǡ�M�hJ.�5Ӏ1ʪ�=[ژ����Ȳ:��]M��k<idT�oI7�4��&]̚��e	���&���{ީ'�i)W��I��L�շz�;f#G����8�W�Z-���]����l\��(J��V��q��ݯ{�+)�<�<���u��bj�CN��ޖ]j#�,�D�� �5��/ZcL/2��{t��;���^�1�ҙ�E� "w�]Dz!����J�CY��'c��q�21]�|�ۜ��U�-�um� z��W^�;��̨��{O*�g��le@���H�ӗ�pq���V�R:���$V	J�U�D�/)��Ҡ���᳔"��=ZQ�G����|�.��;*�����s9"�m��]�Z��*cG��h����A
;δf�cRZ���@jl^��K/��B�]뙙48&е����m+�_;N�J[Ru�w��Wk���36��.�{�Wr��P�xp�"�^���uϥo�T��R"��$G��^;�S���M2��ѱ{ާ���`�qu�=W��9�)}��f�g*�Kj���,�&��\�/��]���V�ؒ7j������v,T��%�ĢӢ��W,�6oT|Л�l*�-�n�Gq���3��^XW��T�z�kP��l���i���F3��{K��@���Jh�1f�s�1%4��0j�z�m>��!��Y`Γ)h��WƏY�]�k�S�Q1>4ٚ[�f��G�4�Tt��.a+��a�sE�����ȺM��W>�I�ؔ|��ê��<�0*xz(o1�9*Lj��;�{�QF�C9��d��%��-V'*�%b�e��c�I��
�<��L��*�#��Y�hY������#�we��U�; ��:�P�*˼Ѱ&�w�04S>��x<�1�U��>~��*�����ʯr�y�0�G�2�I����+ʐ�f�5=�N<���qgnux�E��]���Ku�{V*V�e�`P�9��^*��HM��f<�t��
U��.�m�s�ʦ�^[�.��UW���cF�V�|��F�,3�վ��#{,X�R�ʱ�+J-��n%����u�Y*�b�RڙX�82X���%P��:%�G��=$�'�KYU����2H�v��n$�ת��:���3��Z�r5r��3�T/U+�U��x��[ddO'dY���'Xp�{2�f��(�&��	:)���Se�#m��<���5Rc��v��*LW�m꼣�U,����S��F3�N����1H���X���������(#A���ht.*�y^=֫x�[7���'u�=�����|3�:��ٝW��%5B��|���Ң�mn��W�8���>�d�r��Om`P�q�]n-���a-�Gq�܉��{��b�Ԏ�7��di�;��{#L����쭪���Z����2JY�x��k�ە;5Z�Y��27Uu�&�Rջ]YqF3� �8�4�׍Q��v��)�	Q����7k���ѭ����s���UeI4"�9.6&�ʊ�^�ܒ����Df7�:u�ޚ���f��fTlс��"�
6Qw�&��n��#�*�����;��D��t֕!W��P$��٦��J)_u�<�s�垣D�$:~甭Bn}M��z�Nԑ��=aK@�lڋ�\�R*Uγ W�ʚ���t� MnJ�p���qn�Qz���b�E(�³%�cg�M���0,u����cs�Ǽ�����F��M]P��z:�[������%vM�,h�[5�I��c�ö�l��S �N���z���k�Ԯӯ�9ێ��Hʡ����GW�^��h��,��AyP:�ý���D���!C�y�3���YjP<�oGR-����ĥ�$��v�s)�4/[�0�!`�x1��j��89��Wlə�[F٫Ι�aD�!&�o����nU�7A���2���e9m�.|cԠ�;d[-S��f��n��!=�Á&"�5���߰{kO
����/^�C;|���>\zRV�oJ���j����
�A����u�R�6+kEv06���;E=��o��]wt�X�Q+���ʏY�7�˯���`X�f�B���P�Z���HQ��5��lTP�����C�=׻���ۯ�և��Qf�+�-̤���uH�SǼU��2����U��n����Hd�絷����v�%�P�����gՇ����yv�gY������u���Q�-ɗG�̭�DT]����(ьN�1'kշ��k��*TN���jtI�W��Ŵ��`���muqc�^Y�V�Nf�����ggN<Q���	�}0.\ѳ�	�ѓ)G���W��mqY�����ޠ�L1_�KJ���a�鼩����X�jK��� &��˳2��ɉ��|U��9�!�J�|�y�	� z�C�+5���$��gt�/���`��4cƃ1�t9�u��j��+��Uk���ď7-�ݝ4�qԮ���ff)t�l�I��-ԮYj�3�y2�iҡ�V#WX���F����y:�f��m�cZ;pU��j��^�2�aױVm�hVv�k�R>�5�$j0r��v�m������V2S]*�y�X��,x�չI��n;�b��CY���8��;��:��`w��I��&�6��">�4Z��Eq�"���8�Cv��N�qaak;��J�A_���wz>�[��T�*�(:��6�,X���R���G:���/;z��WD5 B��'2f����zP�)��������p�P��٩�ca^��k5�a�*h�Qs��:���۠4�/Y�<������{��]Mέ�O�ǽ�(d[��uH���!�^�P�kX/���m�6u�����۹6x�X�3�&ug,]�N��������f�;-q7���wh��*[�־y��n7AV�}K�g�RH�X��7���먻��]d!t<�u^�K{B���a��ؿ)}{��K�<_S����s; �F��T�J/GF������w���&āR���W%0��p�er��)�P݅[óA�����vM&��2�žx��X�1�E�Վ�+Y���v*��}�jaR��/Ae���gMή��7-	�n��M���\�;�-�a. j��a�R�������Zߍ,�G�.��hծ��.j�Ӗ̶2�g���	]�]�uUCڮa=�a�Q{���[�=����E 	�?�������������!�$�(�yZ�Kj���SM�!fH�l1�O�))X�y*Qq8�Ѕ�d$�LQf\&�ͤ�J$����0��QS�"h�$D�A.D�ˉ�?��hJ.H�����6���>�j��j�#%�Ӑ�э��i	��_@d�6Ѐ�j �1�#/��D��#�7�10ci?�R(�h(̒���6����E�!��1��\���鄣H�1��&4�q"�.�Q$�r#���PP�p�%�B_)#����W�4�0K�%�z��H��	��b4�Lv�����x'��_dr������("GmU��݃�<Z&��E7�`�bZ�:��5�Iv��.�Ӿ�ZugM�]�V���׸���+�绊��r��en̢,ӗ���1��l}kx�c�9�%�k;������s�wT��g:5�TX��Bfb]:I������ݩ�(ī�X0ԖR��|e��ۺCo'6��\]^��Tv�������;^���
��%�{�MǋU�cE���κ��F�������6*��c��ڲf��Z�0��Hx�oR�{Ӗ=��Ӈ>(��\P�W�@��	�9*&og��ŌL������{GS��qw+��
�d�b�S��ֺ��g�]_D��4��/nL�:3�{M!��e��]фfm5���[.���X��:���}����o �Kz.�b�Bm��m�*�noC���rŇ�uwj����mi������XT����8n��.Q����ى�E��B�n�.��I,��Mٕ�M�����u.�U�J��5�ut�4q�|S}�2�q����^�bw8�d+T�ֺ
R�n-!p�9�n��]4��ǩ�d㳇K�;�D1@ќc%�p0Y$�Q��P��f�I����a��!��n3)�LM��L���G�M|�dH#H��(��0�m@�E�|�)�5��
aȒA@�H��p��R`F$�MPr1H�H$�	�ԙ�D&A���dO���2�D��Q�I��$�8#��
&�i�g�"�$�DE�C Ě�[�$�1"3��
dT��Q
���R���&c.$�"���d��B1/�(��*H�a�(��>p��!"CiSi�T�&
p'p��r2�D��Q�[�B���E�!2�-��%Ab"`_DHN0h&�	9�!&bM���j�Ñ$�
%>���'$@A>)�X B~��$�ZI�SC
C���(�M �3)�L)�#LE	H]1"�II-g�}	����	4"�BM0�	��HFYf|aN2�E$�6�(�I��d$Y�5���(G�4�b!� ��A|�l�*8���"�,4�¸hB
��I�	�A����w��b���ͱ���Z�[r׫�4��1�ć\x����q�x����:�o����hҟ�hT[E���m����w��N���8�8����:mӧ�	��|bܶ,o3V��j$�	"H$ �8��\q�q�<x��M�t�uq��I�
����u�$���x��z���3.l]"�[���HY�gwK�&���MI�Uɻ�Ԑ��������U�ӻwp&��˲wmW0��mD����)<p�uݶ���p�_���\� �����X��^U�o{����ɪ;���5gwe�b��iwnc*�<o$�VX��j��t�d;λ�&��.MD��ζ�x����7��)wv��q�es���ݹu���w]��v��byO�&Qq��ML
�c�y���g"���N]�wn��*�2殳iM���ݹ�o���Ϯ�+�r���޷������#K�޷'�p+��r��Q�u`}�J�ꅔb&�Q��HrC���B"�P
$*6H00R	��(s���U�W�����$�ٹ���̮�<��]�7��I��'�ު]z�+ !��,�u�w��DH6�e��1��FB��Bb2~@��A�[4�f"S���J|��NG".$��j!H�BO�m&���HJ6� t�
�"�w�������U^��gׅC��,�z��z*P��[�L�
�L�W�UְI�*��N<ֺ�=�<����i�6{i�S�Ӿ#J�ц�:4�s�$^b
haJU�eP�� ���3O�b�Z���ոr��d #t��s�6u�A"�Ί��4�hŌ՘ڬ����	�x�M��V�F�3!z�U9���/c���O��2rnU��K��:sT�q@V�x���0�Q7��*ڱ5Ml�$/i�a�/�|���O�3z��m
�a���:���䙘�aN����±��0����#M-�$L���=�� c���a8���Bd�]�2VX��P�b���J1>����S{&���Sκ�gP_)��uϊ�@7�x+�����~�9�t�+vaJpf.a˪{�E�����y�k��38��	�3��[��T��~�!U껲��Ѱbf%��_l��w�fc�t�[����撝-�cx+{����n�%H{��{�9P���wH�����[��e�Gc�_U��,_pW�hn��7�oVk�v����s��-r~ʧ������{9v�	z�n�,�_��{s.���3��r�0h�m�QK2/cN<�%��n�������auF��#Ml��$�y&�""C�Q��E#���m�7���n�+j��l^2�k](����8������t�w���T*���[z�W��5�Hn�G]��0�Ī�����*
��Zf�TT�iZ�vv�f/>z�i#o�F���A�u��49�CχV;��]*,�U���sL��bE��>�,�Y`6m'���O"r�>����g ^)I�
|im�6�D�<��:�	���4/��c�Q���5�f;�ϥ%(��C�m���p*%�}�;��j��@�vJ@[�*ļ���زY�>��q��Z.�;Kq9}�g,'����Ï�F�m6��E�+l�E|���\�)N�p'sU\5����+z��8�b�,�ڸ�W��!t����x���{��13 j��s��H�O!��V��!����w�_��
����\��V�H���������W����UﶪK�0��l��|;�I���W������`I���D��ݯU�bh��&J�۸�+E�t��ȴ�2�g��Z	�"�R�ܘ�����I�2R�d:H�:�)[/u��/�4a��*��g����`�{ݬ�ͭN�I͎��B1�q$_�$Ey��hT֊����V�e�x'j
�
��Z[cH������]��@�f�pߛK�k��m���7�=�rU
ݰ)N�X�$C�Bk��tIW�A>A��|j�}]E��W!�#�Kq��/MnߩA$pr�M`v�*�r͆gw|�Y�PaaD(U#b*"fQ6+4Ȋ�.�r��6ln��e ��*�3��٬}�oL��e��+M�g5df�u��Q.Y<�'�^�'U�3�s�r��z��k��SL��1v�J>�<p+0ʕ19m��B�N�|�>�E4=�x���[;���ێ��w��K���j|�Y�a�C��=u3U��d�I4�J[m'nD�u�>���
}T��ܥg��\��mn,Ȕpm:T�6�I"�84�B*��ٖݕN���.���ql���"K�|�s�Q��u��)9>U�+������12�f}�v�gnJ����'4G�ِ��Җ�,H��6"D3�ʩSy���	��ǲ�q�KdA��G�ݖ�O�v}�}/�{0H�r㥲�Z�N��a�c�?� O�hB�k�zm��+�M��L7o�����q�f}6���H�>(��K����,�Y�" �^L�Ywr�0�K\��Ui�#B�**w}�o`ש�}�3Ѻ���&�5X��[����+��,��d
Ru����&�Boi���m�KM���6��'Ө���� 8U)]b[@���{�:p�	�����{~��2h\�w�W�M�|n�}�2bso�j���Q㴣Ad���W{\�j�=�n���0*[�]c4·�yOd���
���]�Pf;0m�k,[�6��8'<�q#|�����u���_�z����"}Xߺ��<<*��W4w�q�a9t��b��R.�ћ]ɽ{y���7�{�|�:��\��F��w)�lh��ty^���ۄ��8�J[�� k�X�ʦ��O�R�#�����Y�b���S��0��ƫ*����������6�O�Eʓ�s�B�"ϧM��@$��4<�̈́�w� G�*��OKb,��X���<��瓸�Hj"nV�lS��g5�_X���K�}21*����{F��f_�g�L���ӟwXw��&y��Y�r��')�*��j�"l��A������2�B�n߬�/. +ƥ�;�yIT�Y�AkhU@�C��V[S��J�ES�l茶�W����'+ �7z�N��?�S����%^�"�nBGKTDڭ/.�s�4�F+u���L�"����R��������l(EF:f��*�"I��Ze*FQV5�Jòٟ0���U��NIҡ�;�CD��A�Q!xAus�/�W5�t3P-�UNL]�o�]�J�FkT	�l�F$;my
`����R��1�l�n�����Ű�@�K�ت��ղWG,eP��5v��h��U����G��$|�<<*���=�ް��_����;���^�%f� ���ƻ���U�5)9��=�����+>�r�M,�*@�V�d*c���\tP����*��i�
w趞z���%AP|͑��W�oS^�#o-��Cn['y����nj�
���b4�4b�S�q��W���7�o����A��y*6Clx>5��m���=B��hLJ����?[���ފ>����5��5���|�󯫊��E���$�WV������x-��g���i�Aܨts=���[�;)�#�k����[¾.	�t���b���J���L&�?�Fb�gl��;�p�c�cz����M'�я@��T>����U�-*���ߝj���e͖�A-��V@ʬ�lY,�?��!Q7��B��:h�j��(�n�4d�to��w�+���
��E�;{��۷c4�Z���Φj+EnT�]��!l�<8�m\�$��r���GAf`T(�Ww/���ᔌ�E����epY���`2��H*��I���#rE�V��y�t=�/jVN�<�����P��F�f�cC�0&]��(K$wQ.oվg+��N�{m@���4�!m���V �Ù�3�Q�Is� N�/��a�-@�7�s'ƛ'}o~�S*�g��󧋛%��s
7�%�ډ�x+}iT�VC6���T5��c+��W��c�ԩVI�A�16�l��c8��o"��а%�5�|Ŋ�~�����߳�u��/�R4%P�E>ǥle�M-V�=�k��U9��#M�55n��̩!5��F^h@��|^��흫�2mlM\�ˢ�Yo�Q��ʕ��>�=��P��E}�J�i,Ts6sFt�j#�����Na
35�1R���/%���c����k�8�!b��5�읽�$����������R_P�fA������`�7�k�X���?�����|����'���{;hG� ��'�-_"�klYƬ��e��+-�p7X����������*I���K���ٻʵ�o%I*��~nJ�E�%K�N�Z:�|�!ۛ�u�'x����܈�����r��f�b���vƧjP}e,&�ȯ��^�P������������(������S\�I��s��{�GX�O�#������R����H���'ꭏ<�nM`����%$2"W������J���ʠ����긹�1:U�^ϩw�E'���'�}F>���۸�y���-X$-� VR��:0�+h$U_��Yܣ*a���DY*��ܪշCsA�J��c�b�\�?����5ZBYp�j1C�d�r
"I�UnׁUz��E}�_w�E�n�¼�*9�-����p���mB1���m�[X5�*	y�M~���ȍ�-�{Ϙ�_3Y,gxB�1)�e�~t.'���1���ҕkʥ�Y�/SU�g^�G.�6�
��]נr��4_��MHfm�3��n���[ع�®|�m8m!nO�>�U��g}���)hYp�(ƶ�rku�6���#�x�nn����:�♋�e=+}�=i6�#}��4��z,��ZG��eMۊ��X<�� +�O�����d��Q6K�'Zt����К���m�C��ԁ�mj��p܋f��׸���{D��B�1�bVS6�$h�לW'�t�;^j6�.��f�*^e�@�ַXVT���V(iޝ��%��Z�ħg��e��-e�*�̡-3-@락�/p�}(V%TLy[�����`-P���L},�-n�_�"r�Ru�� ��j�������O$��T����6��%tp���*��GM��HF pKڡ���oK�LV�I+6�ec�Q���d5+� ��{��@*(S�,�(.%h���C�1WA�j'a�����V2��|a�SE#B��3�P�bR4�*��9@����G�6-��A<`��e[�hg�g���[)󶠩��2��~$�����U�b�2����V��x��z�& ���P�0#FF;Z.,��Y�ȣFA&�Wz7�x���$�'���-[�\��vt��R�a�cʒ�Ǧfm
���FUR�l���s} v���=�]t{�o�a,�4_���+CWMuݞxiM����}�eoT/ 7��9,B�Ø��PKf�ak��;�|Pℳ�9�޼�;�itҗ[�
��������AX#�is9˕�f="���6��c������^��f���`�s��N�eVV����(�!���dl��	)��/0�.������A��FS��@���%ZD��c��W��u�� �h�3a�����I�6֊�V1�ၨ�Ǖ�|�Z֌����r6�׵��)#d���J��+ZV�n샶e�	��$��@l|�S���M{��R*�m��y�ѦU�t%>_�}����RC_;���"�5�p<��;��nV$ה{Y[� �&|�+%���vu[�����ϊ��V��-���g���H}�N��Q5
w%�Б�����R�;QK*�g�'�ί��[�d���n���~���k%[#
�"�!j2|4�|���C`�n�$�q��8�%�Mջ���%-����\;{+�Z2Ke�����Bݜgqa H����H���sΫ��1`�Y*r�]ΐ7�gW	4���r�gi���b��i�O.���� ��^s!%/�R�gWa��G�d�S�E�i����7��a��re)n�Ňq�n�n�>��Ǆո������Y1�;xja�Z��:�g$)�\�L�Iܦi�Za�E��7D����YoEEWs�����(9/��n�;��R]��fZ�d�%��8@��ި_"f�Ki2��7��iɚXR	��MJ(r�^{��ky���W��Ӳ6>F�����d� ��3udu���;��l"��&�ѫ��C��A�L1HpΡ|sg+�+)s����[��M���m�5\P|�E��;p8�̩�|ĺ:NA׉���O�WɆ>wY"�/�ĵ�/�.rr&����.�c��I�]���Q���3S�z,�l��k_�YT�k�<f��*�n�<�i�T���ٺ�j�7�M�U7��9no\�x��o/������gg�1�S73�U�r�Ȏ���],]������^5Aj�G(�IO��om�5s�9&Y�����g>�K�Tx�o>�Y�(*�x�h�fSe���2��+�Ş�������n��Mn��	������,�3@�V>S�*�vz�!��Bx�yoJ��Fy��'�%Mf��U�p�]�ޘ��[-�x�ݼu�L0���2P�QH�F��#@¾��K����[C���u<���|_!�!��f?ޡ㚄v�n���[�qR[��a���	xcwZY.��htm�j��*�+��a��Mt*�j��M�K��Y1����8�X9e�9��V�_�;&�;K$t:�Q���N��}hѮ�w�&��*'ܤ)�ݗy�Հ�����i����ׅ�x��#����!У�r"L�Oں��-Q����N�:\�hɓ.�^ЕI�v���3�Nھ���\��2�/2ldb�C�k��.,�Q���'+{��GroL��������ڔ�v(��d�CTu�vnC������ ���+��l��m��u
����󭰸�Om��^�K���u�j���vt�z�0��-�����vb/���p�;U���X�կWC&����eU��S�9]3��e�M����Xc3.�OA����k�f䊖������5��uݱ%���䩐��k^�Yy�y9v�b��ű��X���r��e��+;�Ns�&�ł�
����7%Uc�*C,L�z��ci�ξ�ʐ��6��ބ�//��ȎY�݇3�](L]Ո��`� �f�ᡬIك�v�>�3�ϩ�7��:.��Rce*��.;������ W�"�
�=@x�(����ݱns�_�1�8����z��__^�z�}o7��ݾ|cE*)2k�\Ţ5��6�}./��]z����o�z��ׯ^<}}q��nݾ;oA���r!
�[�yG��l����1����d	$$BD�z���n�i�^�z��_^=z�۷�n�@$$Gp�#!�>�2e���_[jp�Q�F�񹱶4F�5%�n��R������Ư[��or���vE%3�\�cW�r�cQ�������cPl�`+��眅��\ɾ���μjᤣ\���>��D21��"��!Q���M�W�xT�r<��X�%e#_*�
���;C��bTm��ۭ5���:s�E��=�u��~h�=�]Ot�i���hi6�߾s�C���z������i�6��ݨ�^�3���Y!�U�v�~N�NB�J���>����lEC��@�}ϓ�G-mν=M�t����`kH�B*�]�_�������L'�z���X�%�f��5%Ko< �qfս�\�߀=��w�jz�--�8����es����3���ˠܺ)�b#���A���r��� �ܟ��|�冊�v
I�a|,��J��U�-�O�o!��lݘ��X�;pͺ�Mk��5k�M�ln��7	(��ѩ�1�ޭߕ@�/��������7���O�r�0f�o3330`�N����^���]�a�7�Ys߻��sz;�N�}ņ�U�~�>
�v��0����(^��c^���g�����x����P����	�|��E'��
cK�s[_���Iȸ~/뼮��EJ��8�<��p������o7�a���]ρ��35&v�y�;i0-A��Ve0��$�n��U�����J�UN��+r��-�B9��`�t��[w |�Oa
��=�n��N�}�7C*�1vt,c��x��4+~��"s�l��	B4j����p۵�	1-�/z�*�qx }�sU�N�l{{�Ox��s*�]x��]#[$�W}�b�����Ui99+=�.�L�6k9�z�uy/mP����D�����{�iϲ�U-��z���xy������*.&�_*[�S��W9��qo@�k�J}��zݮ2���x���0T�9�Vy���:.l(�ˮ���_5bA�4�������1�B���p��$N�C�Ch �͇�ך�%�M6� {�z��=Ə�/h�.T��tn��yA�(-l ��p$C�x�jv͊�d��D�����}`�ǁ�K�v(�`S>�J��%�g�����@��,P>�h%�}t<WwV�Ω^�!�cp����7�t�Dٓ���=��ǓS
��v��&=qͼ��p����Vc�U�ǀ��Q�~�XQ��~7��o�w�,��܀���� S��[���d�O��`e��;�[��1[;�;T4 -^Z-Yz}�"O�@�-t��?j�j���ҧ��� 	?fYP���0X��9�{�����07�� ��|U�-=�O�(`�hv~=ŷ'�D��5f�d��m�3x{ԟK��]0��R�>"�i���X��N�JǗ���Z�ڢ92�Y��ub�3<��Ɯäl.��~���>ѻ�«ϸ�5��qs�Ѭb'�m�μ���6w���� �)�8C�w�{b���`|���0�ʀ�>V/�U�`x�.�y�MV��)���`�vطv�n�exx\�<�(�s�-�+��Pe}Gr���E��{�b�i]G��5�'��{!� ��=L㒗K���e^�u�^�̸����o���1+����&I����=�̺���u�]k����T�0`A��0;�O�/>����q�%P�������L�f�����'>���H��B�Ô��pD
�9���:�t���Uxu�\���f����N8^K�î�/�xE|`(���@gƢx-��@྿�n�W2�n�V��/\���M�A8�p������$�!��\���	�^4 |kEO����cè	` ��]��c���ζ������/��7'������u�H<V�4/��5t7�~�9�̽t"��n�b{� on�M������"�rw���p�cv��>�����B@D����E�ð�LRu(����y�Hkk��yN�G��8�zK
[ k�+�XO��w���w�0`���}i��x��n���VW���>ko:q�i@��2S�#<^�BOms�a!mN�e�C��:�Y���b@s~��ς}ϒz)����+h��*Ki���1��}H����#�FS��{�h���ܢʑ�b7��
=0��	C�_�>�m��d�T�H�{^!�o�Y��ݼ����ţ�Z��C�ע��!h�eF����-�h��}A�V��dS�� �m^{��/D�G_n>���V�_��J��W�sj��1�q��q��bv�U���`�ut� u������oL�`��.��˧�Ɏnd
�	�,�ו�z���0#�<��tR����Jm^�!��e�g�OkBz�|B1��a�!$���Ҕ��w��f_Bg^�4=r����}@Dg�;<* � N|4y�$�������|���F��=k��s�W�퀋��xj��Ǧ��g�o��T�@[�q״��K}}��G~���J/�m�Bl#2����������� �V�Bԥ_�FŰٮ`��RZyX�s7���ڭ�E?���&��y�q�O=�r=�DsP�D2��^�����Q��
����;�|��z��)YE�yك�B�����>�5_k�-�{����{&��T�{�n>'���4��6$�B��ܮqX�`aMQ��Hqls�p2����v��z���z����d�8K�;8
�6����g�Ih޺;�>��uu���R��P���F;�xkd���v=���nWQOx�Ζ@=��ߛ��b���uIO�^)�}c��B��f�`;�O���t�Q��7|<4S�s�X���X��Տ��ڍ������I��*����bі-}Qb�X���p�z�7��&�F���p:�i��B�%ԥ��}�)u�_/�n�{Ӗ�",��-VJ��a�͍����JL,�z*��Ws�Ԁ��.�u�+�u�Ǵ��G&w�-�5	"l7��S�T,�����/��o[{Q��z��ME�������%)�_r
��7��}ٺ�3c���@?�^�q�(T	�c@��4�� �=�ݸ��}�(cp���{N�?Ԑ%�A�Zg7�@;>|�x��T�q�2qt1�-�m�~�������u*y������� �GX~�!��G�Lh�2Ԯ�9��g7����S��w�k��	���O�G����Ԡ����)�N�Y%a�*υ��vZ1W�]}7[o�i�o�w9v�综^w�>]�`&+/Թ���>jc�o4<t<��.��>�\�Ȃ��������p�x��i��q�@?!�z_�xt�o`6�̫`�/��@I�g�` �K�J5�۹���Мɛ;�f~ѡX��ӆ ׈���U�ʮ�BW9	�*��{T�]�ЦY��[\�v�9��U�E�d,�4X|0���4�W�ف>i/�gwP8��?7��)\׼zݩp\q���'���K(=f������R*|,/�/Ćꧏ�~����и>�6�7�Tڽ�;�~�ߓ �����A�W��Z7��U�>�V���lh��{� j�t���é��Y�*�q��3w��pS��}oA��%�{]�7XʅWm�f��֖�J��)Y�c�75��<�=�Zu���AM�A��Z�GW&̫��}�o��!��>��l�6����>92�nb��x&U���m�j�ej �+�⨌�Is���3sL�9h�v��N	�׍�M�nh�W�����sw���\�~�~�cJ���ЉcAQID$A��9���B;��+��Ͻ00�pE�Pq�d��>��Y���t�[u�\�� �s�q�0�:�^�U��fA�K�[x�qL�G�C��j5��
|.	q$�W'd�s.֏	H)-᭝�Ka���Gt�k�1W�]���HW�yK@^,@Y�_�/��(FCl��O\��-��PE�mצˀ�dg�m����/��^|:�M0E��]�����k��4y��gE�Ll�ޡ~�N��sd������6���%��׸%@�����O��%��B�@:���{�r����A8���5]#bw
i�]�e�z��ƫ�s{�^m��K�|��H2�㴃����<� �%�!s
��x�K�ͯ��.��閮�bK���[���)�lF�;>yh}\߰F{\d2��C�63�Uw����;�tx;6g�Y�T":�E��d����@9��i�ydy���җH9=w�n]X�x�Z�($6&S��;��/����w� 8�}��
�ޯM')݀Mӭ.ެ鞳�og�՞��ʑ>�z�����<<��DG��q�)�7�׎� �v| �K�o~�+M~��ۛ��oZ`GD4�Y��#z�nr�� �jL�]�!����N�����Lp�
� 5��>�Wy��F^Йؤ�(n^��/��Bty�X��4�ޛ�pΩ��V��i_rۼ��<�7'У��UcLhT#Lh*
@*	"�Ǟ�y�w�{�hP�?X��r�Z�53^�u�����$}���e9�{��b��4� v�'ƾs�yo[J�d3>�<�l��6N7s�kzk$ιS�D���7|��3���Y�K���5��r�ױ-����/N����aa���=�m��2�� �'���E�&�=n�^9>�	�J�	eA#X�J 8�nb��lx�9̀�}�y�"��3�g~�A�7IR��^�]Aop2{Su���{�	��T+�z�
j�|d�r��n�!�7�2��oٌ�?s�x��P�ފ��u�`n���C��|���U��5n�� �)��0�ݵ�r�t�=�+_"��,��`Y��??�@Yz�P�&�7H��!�Y����M�RĦq��YGm��{���=�"���צ�lw�L�c�=w�&t�w��tqi�ŝ����F��G�uWx�����sνKO�`�>�&3G��5ն��M���9��1ÞZ:�e弮� li���SF����Nw'��0п\�@^�&qS9�"`א�c���V]�87�U-�9^�|Ú�����������ٝO�v�RaW�,��aϨy�邕$c2�����ٛ�'3�B���J�=r�ZÂ��	M	�Ҭ�<C��3b��Q�n~Jz�6W��څf���k�1uk#^T�Lh8�l����sWWr�[�qJC�I�O��6�$��E��ur�Vt������8m8�0����D�i�($i��i� �QI$=�>_���߀��С��V�Gu\_>�R+��?����r|ꄞ��,��u˧Q��S��{�g}��t����q��|J���@�hv��<g1������Wճ�����ʉ��I^�z���$��|=�����������X%}��H���]�#$j����v)����u���3��Ǡ	�I�\�m[��)�z�\[:y��EE�+�Ǆ�ݣ�`�M�{��������w�9äav��C2BN'o2WZ+�|��@��cG��{[okn%�����˞���y`;���W��Y����o�񁧻�Ϲ����{n��ŷ���2f��h]v�|�v�xg�����x�
��X&|��.,s�<-�װ�+U"R[���v��n�ξ�x��T�7���Y�g� _�����\8���lvG�t���T�n)(�2;&p_m2^J���	\��v��ަ�������P�2�ߎ�HX�����z���T�K�n㞮St���]�)h�������P��^�]B�F�c�Z���5�<h	�0�[��O�7�Rږo���v⛛�<�����Y�����7<z��oJ�N�����p[�	����D��Q�E�n�h��J���y
�#�����jj,ܱ�z�7=����;�6��(m^���`�ې���NB�Ob��N+}ݘ��W������/7k[�kѴ]�7kW5*SLi*
�
� �'� 8�Υ�<�w�(3�����u��Y7����ܫ�P`.)��9�O��$(k[�{�M=�NSl]vt{�+��x�~�c�=�rs�Ȥ���w��t�Y����09�L|���75�n���Q��Z�{�[ ��>�:5ׄ��ٳ>�r�I�&^�P����tP��GY��^���b��0��t���
��Tz@䠕�s��Iɮ���3�k�W���	>�������߀j�d�X���K>�����L�B�Q�4?A���S�J���O_
5��D��2�1�S�:˼����wEyt����W03<b��$�����;6�5óe�
]j�ӌj�8�j6��p5��Ƨ�*G�^�O�܉ ����5{A��D��%>��Ѽ+"��5��w~Ǉ8�#�����b��`�zZt��%zǥɫ�� ��D�����Տ�������&�Ç|Ay�PNr���>��b�gŨ;�����Jh�S⥚�[W���KsF]�b2Pü��s��٦x"< ��u�U�}~�A��
�τ�9)��7�����V�uS�V����]�p��=�:0�O���o{|7co��i$1FS6��+n�v/�c�
|V�k}�[a� �y�]5���]�yR{�� ������w��Y�ق����ul��������f��@5#�4QE$V44 �=n����6��j�mmk�����L�߀�\HN*��g�,�P�xH�h�о������~Uϻ�}�"�n��]�|�[�d/��6r�鯽������@V++`��y����ܟ=�G�y�cu�ES�xOEھ���;�)���g�a�����&�x��7_�8E{�1U�?Y~\�H4k~�aj$��vW�mK�&���l�cG�#C{�V�I�r�n�<���}_c�Z����[�K`�k��������X��
'_��ư�V@![������IX�������G�զ;��hE�Օ��﹑e�ow�8�jn��}$r|0�0,C��7MFלu^��PJ���Ϟu~�e�<�>�{��C��mK*s1T!���Os�	�q��3�üǝT?���cF�����+�p\��O1t���(��`��mHFq�ZԎ���s!G�{_��fO@�)���γ��!���[G�SL���+�4v�*��|�۔gB��p1��iO�cS���������i1�e�ӏ��[���k���Lsf[�4���݆�]�5�:�-�#&�a7���2S͵t�UL��UF�j�W!�� �6gg��Iϯ���Y�"��rcs�t Y�<������J�"'�f��9ٽ���� �޽K�w�rko�����4�-��l�k���-�:hqk�Nn��E�e>�/�*>���q9��K]/�;5�w���{����b$����֜V��l�m;�wWfv7N���f��h�1�������r�fF��b��]c�>�K]�����YPZ7�軯�X��;`Ý�1�e��`zk�t���ҥ�\do2fu�!Q�}O�(T�Ⱥ�F,�3���|��6ݍ���6+�1�����Oc��1�݀2�PL�C��Ժ�����(m̭�:oZU��<L�V�*��cd˛gK��]YI;#,��{Um:�jQ#�Nm_>؝��sC���kkh��7�X1��U�{Z���}�+TzH�j��|8���<`ժ�
�'�u�9^��up�� ���rqKڼ��-��D�F��30x���ڊt-���k@m����9(�"޽u�ɡ�A�ܗ0ͱ���N���O)�UlC�p��,ow�v<Y5�n����2�� �D\��S˕����#M�Ni��rVBc��/Z�[tGU�B�Q���9y�j�[�Z��ar�t���۩kM4o�C,Ý:��[|�oV޸�#d*G�b��U�i�p�%Z��hޚG��f�K˰7sj�Ջ�H��#��B� `�( ��3q��`�gU����DX$�Y�L\6��5j����"AR�������'P^�B��pj�I�t�2o+P,�7�����U�ڛ�ٹ�Wa>#���n�ޓ��J�2hĨ��J���-��aCט4��t�S���';jg%�	��P7�e�řB�u5Q`�֪��b�Tv�s�I�E��[�\C�/��q��[�K��f�/l��m8r���J��Y:	����E�^8�~v�쫻�%#ء���H�]3JI@�7&W��GjW|�va�m̀�w~-���.�	G�{;�Q�F��{XFL����E��|��3DG��}�:e:y��.��+�z�A���S#x�;��#�{�KȏPX���Į�2��\P�}v��2۶�����Ե�v�o7,�,��vH��.�8����V+aU*�|t.�P=�2��
���Q�w,s�M�b5���Q�����XH�ĸ���E�x�X�h���f֗ʦ��Z��r���Z돛@(m*r�R_6I����U���p��;vv��2��ts�Z�b>��0%#۲��!GL��A�޾�ʒ�u���]b�j��뛝�IƔ�u��4pU��﫚u��7-f�JwK��2��Em.��^�w9����u���z��usҳ��#.�V,ɋ����D�z�E�_5��f�h]ݼ�9�j4�s��V
�=�=���湧�[�ϭ/Ί�_�?a(]ŏ��v��q�ׯ\q��ׯ]�v��ֈ!## H�-F�BE$ID��F��^�x���N8�8��<|z�۷n�:G��-�X�VH#F�+����n�;q��q�z�<|z�۷n�:MD$�F�Q$$��j��������E��^5�uʾ*�l2��v"�m�V->��Z(�I�=�|�^/�9�sk�!�p�߫Ǌ��*��}��M$s֯&ƣRDO��*7�sE����x�*6"�M%�k�J(���Rj"�(��?^/�<���i�{�NA�|����*[O�R8Q&m �AFۄ�P6D|Io�g�))$���%2:��t���K���ut���p������L��8�U������m��o&%��v���o��`2[	#��\a n	ys��y8��o}:����u.�"Sb In�-�A_� SlH�-�����#m� F�M�`h��`�~F6� ���#$�UI��E��n�I<�<%~��(G�Р�ТT@cCH�Tb�T�d��|����z5��3�ǿ���Z�c�X�xdV@��up�a����4�l̴'�� y��b�Z_}%�2���
2=J#[|����5SmWM��8�1�7ងsvL�d��Ԍ�ٯw@9�� S
)���oX��L�O*��]�)����J�A�&SJ,`� `&�k��c��C$3{Z�^&%?o8��n썽z���0�� �ݵ��C0��(��3��\�������a���pc�.�'�^b�o��Q�R{�5���`�xeyD�p�A��yK�����{N���0t	A�-�-�8pb+;C�[�v�<�� ����)�^i|����A�P]sA�o���������yR@X�6�U�vsU��bهG������-�"@�t���['�`� �� u8�L�
5��zK{Yy�j�9/t�� ��^V��6���o�B	ލ@,9�#O�}�l5�3c�eOz�+�ʼ+�OQaL�j�{�=wYm���-��P����֜�~???O���X-�OHg���_�D��;&�.���UB;_$�.�Txj��q\!��l({r1�W�����г纅5�v}O���`�4pk�^�<���:�"O�G4�&�x��$of�(<�Np�=�����R�(���0��7rIR�3s��EXQ�W�PW�:�W��>KA�Y��q̻��k&��Ů�J�x�*����N:������ro�{��Noܐ׆yy^Oj��Q)�Qhh*F��*H������"H�\;���4�
p��h���z���PJ�2 �a���1�<��Gx�E=>`�f�1������x�����K�:�)�p%���1���^�3E��<M (�"�{z	�:b�3w�����2e���'�I���ze����P�qS4uz&n;��U�R��3�;�h� �<��wʀ�jjl�v_g|��]I�z��e/�������Q|GsԿz�X��g8��+bL�O���+|���n�j|+����;��35|�}���B����+/X��}�Oż˳���Ϻ��s�������h�\�'H���xf��r��z��3��fΌp3��"���-�l˼�ܜ3�/|:!���9��d��
����}r�oT�X��ciM��5���vE��ZY_�gO���~����7�I� <*'�^	7���������={2|p)(1J�ł-��^߲<'���W�ph#�c�w���5  v�ʢ�ThZ��o�P���@!j5�q�����ڸ�gkk���q^��[+�..���u�!\s�����y�µ�y�%�O?q�����|�{w�v��޽��T"HH�<�d"�  Ǎ _�X�O^h��R>)�M�]�K��U��:#M��bWʺ�{I�\T�3=���k�Q8� 44	QQ#C@��AdIV�>o�w5���5������4/yv�E_���s�F6c�ɼm\��ѩ�#h�����bE�a�k�8�<�c����;;��O�3�i�{ZO���+2�߇No���e��*(����vKk�D~Q�`��I܊�W��:�Yд>�9�0$
�����?+}�W&b����PR��Yz����ջ��[���F�>��'jI$��N���V@�L����&Yv�Dָ�v��Ucr��`��`Y���S���9�%��Nw��h�TEwD�0����w�:O�����⛫ݪ��5�yYT*r�e)�ڽ����k�wL`��9�a�m�;nz/�L�O\�t&O}q�}�}>dv���gp� ����!y�0�?�̛=F���J~�0X�<h]���N��.�o@�ou�"X����r"]-񕷴7�����6�/��|#���AohGm	>�-����54�K����Y{�Ït����{����df�0�_0�~a��(<Zm�������ڷ �ׂ�%oO�)��2v:���]��ac7z� �.�	�X����%
D�F'b�������]c1���M�8elT݉%�C ��m�s�n�t��+z��-q�^tD} ����"SCB�M�'s�(x]��%��M�
F�|��
�W���Bn5�z�dlg�`?H�}���ۗQ�w`��>���/?'�v��k<�W���+�:�
��r���VF?����`_%���=3����B�$Q9����௿!|�l�&p�2Cd�l&��	=�P̧I��xY*:�\�8ӕ|4���uDT:��,��e�[��wUEV���O�]v��9��&D]���X�Ȟ8 'q>�w���t��P����V�W���}J�=1�E��ч*�fw�i��������Cw�Ag���b����-�a��V�vZ�x�������w�m��ǻ
������sﻔ�
F3����3p�uV[��-��oa�#�����.m������\7�a�nOar�n��B�ͽ����y�Χ9i�7*������.�}��Z�#�'.���v
 m{g��1���S��_lneN���d������fi�
4�Gt��I%�Ϗ���G���[���kV~�� �g��ᠺpě�۷3��^��A-�'WV������V�����'R�h������uj�
D�澔���޵@�Y�Q]-������hQ\rNux����o_����[F�F�:X����q�n���xx��
hiP)��R��"��)  �(��֧�K�k���ܮ�^�m��j��w�
�XI�9�١6a�1f `�Q����<�#@h�~�t������t{Ӭ2C��B9����.+�)�_AcdD)��K��Y�
���2��ȴ��X��^F� K&��¸>4{��Y۵��^�:�c!u�Ұej��e��G!�jG2���K��ăM.[�1ώ�rA]�9�V��5w��Iŭ� ���Dn�k%�Ͼe���Y]ޯO]H�P����8Z�M�<9'nfm�ǅ��7��N�΋���ɵ"��Y�Nǥx)�3(~ �q���,޽��.q������[���
d�}��Mc$�%۟$_{|lm�c�6��M ��A�K�R��	��{B��O|X<;���k>5J�$��a7v�&�#$6<�@ޖ�Q�2ܲ�a��Nr���ɣ��f�_���|gG�H�1Ѓ/�ߌ���U�ToW�r�����IKJE�f�́����+x�	�X�b;������R��rP��_��8C�u��Kܕ���{7���[?%:.��P��cƷnh5���ø:ŕ�KӾr�,��i11o{�Cf�F���)N�`�Y�h}ss�����1ԣ�f��N�_^N޲'_c@�f?U�|�GwJ9�V�ք��W6Ԕ�g=S�u"�K��L(�yjf�ɸ�8�l��f0Yg|�7�u�~� Cx �(��УM
-AU� �.x�.��x}�������\�@ބ��7!��C"�f�҃�7O
|&6�)�]Dmө��[�I���t�%ó��s�s[c'�!����|�WO)��v���]ї��#�ub�����!ѝ�鯻N�R��C������ا�XGDZm��9�r�92�ץ7�k��e�'Ҍ���څ��'��e�|;0���YcV�	�n��b�k9����X��U8�õORm��n�/>�^�J�k�|w���2`G���xáړѲ����88OÜC)�:���T����ۓ�.w�K��vWU$�**a�5���e_3�˪�vgB�/a�=�,�.D�+�U�^Z�\�=�Be�L7��xw	ʹF�#���w��4ft�V���$-�$=;@6Rz���^�-�2,�O�l��q^�2YM����g�S��w:����ō���b����p�!t��}^=�c��B�|��Kc�ܲ�A�Ya�"�u��M�Ѭ�k�/ld��h���P9�Gn���<pt�Q����S��`;kD��H��r�ٶ�T�O��U����.��6��n�#�F���)Ų�e��.���; >��N���}�����%�3f�� ��ʱk�aLT"��$z��키�m���si�}a�sz��fo��x} ��G�hT���hiZB ��{��ﵿ��ꤜ��'���#4��1jF4��ԕ��D�x��#-�
��h�&�|�,�V�4����і��W���T;-z#�'�k�Q��ϟuD��`��xhI;�3��{	�Z�R�)ӳ��v�d_BPb���/N�Ɵ�xd�՝u�W;�HZ	ѣ�H(=� v�U	z���[��Uz)�F�i�*��F�-��td���w;���+��y�P�a���_ܯ+�b�"�}x�C,���sU΅���V�28g�c��e{k�
�����xB�X���}���d��=mq�9�W��Q�M���)8���uЮ{�(PF0cս[�>�e���P���I�K����{�O5}��I^!��1�>�;��f'���|~V�`�ɘ����+I������]a����{��l���F��ƚ�^��3<�`/˞��7W`��3�ė����j��ܺ{��k~�<)�K�x؇A���p��1I������⛻T�V�o�b!B�k�_�{�vN����|����6�З~���ݘH���,]��׶qI�=���(��
�.p|���fX����x8�T�D��f�nɎ=�.�u�zZEv֗�q���j�nw�m����{����҉M#CB5I���o1m���6�BH6��Ə0�,>�fn�n`R��)U���H8|�R�[�]>Ck�f�G�3Em�wUm���ִ��������ӆ�}������4������[�؞�2��8�7t^%�Ϗ>?
��Q@�^� M.�@x��CY�y���<5q����Of��r/sy��<5��õt����{���
�X�+�l7\0kB�!nS��6��ܕE�7�&��vf8����*��}��O��_|�}�U���T {߇�H=����.��Z:ZGNudGVK`�b�Rp4�����@�� tE2O�Hlƕ)�=�l�wx�g����D� �v&��XCB�>w�mg�EûG 9+*�;N�$�S@]el�j��놩�zV�=�Y������Q��s�'<e�-�v�wF
����Uё-��J8����c�X��Z��ra�5#$�
�lg:gI��
v�=������G���5����[t�}���{q�S\��!�C���i��eYɚ��[�v
J�hX[��B�:�N��2sZ� b2FV6��t�tYR�3zvl�u�|ye��ϵ���26�	�u�vX�h���������8�[ 

�Vƶ�emu$G�����T.X�ei���_�春+x�5�
�:���� +��v�s��A����y�}
~��
hhP���D�!"X�Þ׻����</{�d�����?$�J��m;VS��1���3XYV�Ӱ�N�F���g��\>�r<��O �a�pnl�r;T�
F7v��%陫$Z�3�ա��)�U��[X~�"X2�@�׫ )�Ƈ� ��=�}Vu���V[�A9�������%&��m��*�Y�����"B�YӋ�0a��>����L��0މ�(��Lu<�+\�in_t�߻2������Q�<{�[LwP�!׃U>����]]��v���zWv5�5[�LOyh-���b��-ת}��!�4'}(3ۇץk7,�R�{V�R5y��p*9�^�E��� �ix��0=���4Vxz\T��@���l�����v�{i��&��x^*C�Qy��C�.�^�>9�)�T=����lP������^o9]��KAXwhH'��'�r��Z��es���lWO�*���طp�@��eJ�e.}��m��g��=0�ܞ�;')ᵲ�	�bK�^6����\��L�T�dq��T�-���K'���T7;��A���ف�;���j�L����Br�V�:��s�bfz5��b�7	���4�
�~���è�N�u�XN=˦�^�+0U�������{ ����>�B�E���j6��i����l�;i����p�(�܂�:�p˭�g��}�U��}j@����3�V�f��y�k7��+���4@#CJ��Т~o
��ϟ3�>&{��ٓ�L	�)`}(����ɽ�lF<uW�Cc��O�ϕvef�M;�pމN����"G���UqY]���#ZF�[�ߨJ�I*��������b3w� ���W����M�'���7\��5;��hyY�T�m�����:7�J��,�5\���#��K�-~���U�5'�q��d����L��X��E^��*{������JӁ^��A� h~�v�yaqp	�sm����nB	�8�Z5��÷�}���=x������1	��x�}S�C�5Maac�>�y����U��TC�N����+b���[
d@���;N�;8VP~??��kugևC���7�ӘӥTfjtt��E�tD�+�����𥎈�`v^�ݘ~p+,-!�A��ϝ��%� 5�^g�[N��7�q�
K��M�Z��rT)�,�5��� 
1�p�W�I�*㚈gH���D�<�E7^T�90��4����y�1�exs]�ʁ	��PT�~�K���߲S��Kb|��=Zh��x�ɛ�Rǹ<s����=�#o3���~G��\�-�u�3��v����U���}Wy*P�&�SA��aQ "�,�+�8}��6�Uz��Ά�\�gג0�	۩R���C�aP���R�gcnŌ� �E�9Jn��Y�/�;+�NƵ�%��=�mZ��7�%mg5�s0�Ftڏ����{oj��t92v�j}��H�8�ؕ^_�^�E���=L�ٻ�դ���1b�՛;��%;(��k��`g�rR�,�<�:J��ac����Hzv*�]q��a���Iɹ��͒�[풒c��u�걗�1ڮ�<+����W�0�s������z���e7i��Zͻ�7
P�|k���]�씨fd�Q�p.�W|�=�w�S����9X�Ҵ2��;���o�k/�;��1����rNU}���<��Ί9���HazGm�_L��T�i5�&�Ǹ���Rb�po.*�*h�uX�b�#��0Z#`���,��M�+*���^����(�`8&�
+��9��pS�w�5�5"��J�O*G^A�y�)�.�[q�Vpw�o�d�2��!�u�4a����4Ġђ���>o,��G�t�S5r�K�r�m*Xf����[m�F�-��R�ۢR��e�R2�쭠pc�;�E��GS$�-9� 1��R�d|��=b$�Q:5\4y
������I���K��}�K;jT��tﾶ�����ώ�� #k��/h饌�:A<�ѭ��)��mz록2r�B���@� �f���Mm����j%�N���~�QV�6�GV�x�z�Ŷ�j�׭�n\�x�a��H��w�u�LЩ�!�X�*��|�x����e�Z.TVE���T"����w|2��{��{{x��v��y�nn�q­�xɩ�Z����p�y4��ݯ�kv���LQ()�+@�2�ci���	V�h����Uݮ����İl庚5,��,��N�*�#����]�z��u}�u�N7�����	4����9�"�+U��;���|eӒ�r�fY�fU��S޲g]熮SyK�Up���J޼��wB�:Z�Q5x/�}�~��f�|�0gͤ���:v����Q�P�P��ap�B�yXT�nv>�L�E	�b6/:�̳1���xGu�o�W\ֵ��O
�	K}7�o���b�]�{^���r�5������=j�3+
�җp��r�f ��
�	���7��wsC�]�O+�l+ι1�.ת��^y-�>�U^$5��)�m �ӳ�\���������仕=���w;2��$�$���J�ЃlQW�wU����o�����!P
��Ǯݻq�n8�<z�z�۷n�:r!��A�#}+�{\�`$YO]�z���델�8��<m��nݻoĐ��D$	@�$�,h���`��uݹ������O��v��q�=q�z�۷n�5zJJ6���К���Q`��s@���ō�Q�m��������u\��&��sd�cr�G�r�o4���_ԓE�������%��}}y�r#�����Q~5�8���Z;�u�W#&�]7!w;�~v�^1s]w�\M��r�b"��5r�-�tn�Ѥs�O;\�p	���J���(�Tx�"��q�6��s��nj��Fs'�x�=�w�D�3������Z
EI�����{]-\��u�^�90�Z����4M(SCB 
�G:y4v�ߜcG��n��8-H�G+�¨���-\�=�Be�L0b�^{��S����ػ�轤�յ�)�E�bk/B^y���}fJqv�RaW��Q��	�������޽��)*v�Sk6tqRXA���hk���;>�"���,q�L�����)�F�')�OW����m�5��A��z<���1��Y�dd�\�F��/��h#;����*����z��z����	�x�~.f���	�*�e�bz�L�m	�Έ��GvS�+r����n�}�fZ�wj�I���vc�J��|�8�y}����ǯRݧ�D�y�ҩ�_�y��{�Sる2�{�Xs�*n:�zF%)vX�e<i�C"I�n���6���笆ޏ1'��3P����*������E�^�i�R��4y���������Ӻ ��;f
�F%�L�HcB�B|��y2D!�@���o��ݑP�:*�n�I5<g8��]t��YɄ[S~?G�:�a�.ƿb����|n�.���C4��&�9��\m�8�dr̋+,r����][Y[���R���i��V�.��F�+�����J&���~"Ω��NZۼD�ռ���:�6m�t��ʲ�׋��H?�Yl�#�VÊ��%��~x ��h���A��y��+γ���^.����<�x�PE��-����=�8�sϙ��u�Sd-����qb��yO�jO��Ds1<�|�B�iﶅ�ϓ1PⲵAJ����(ы7;_c���}��7�~���f��H���;�=�؞%�?��ܫ�1z/�f�Z;KErʌ#N3���q�w����B2:E��䢥��'��\^)�m�y nTD�U�Wc֎23�S퀰�"a�:�ߗC��1����\��A�&]�,Gf([3��ZFv_N�;�z}_m����/C<�\�W�-8b�N������a~ǚ��nH�ӜE�4A}x��s�*�R�/�[�t�\��i�zw��������Á�^��ϳt���yCA9ɩtȖ���
�*{^��{��]ޑ=u#K�\0m�`T��a{]g�=���H��hh��D��R����H��y��S�נ���"K�gc�Z涺rZ��_n�Ld>��!��^��8fV
���xbG��Qh��k�c�t��墶;s�z%���Q�ף��K���ż��Q���%�ua4� �]qk����J�z.]�Ұ�4��ݻݻ��/fݹO.�Me��Lф���'��%.5w�l�	ݹ�":'r..��n���&����4�M+M*�9�����7\�im�T�c�@P���;z�����!��}&�*�M��ֹ����]�(�]M���>���кC������@q�*�Fs��W�=�c�B��	��oq���������5����a��HȌk�uP��W�������_L�H�u6���f��X>�����ʠ�zu!��Lu�QY���>���_:Ƒ&� ���ݘ�:�K���^�P�f87.�a͠w,����'9���v
I�a:!���;��v��ֺ�I=�-t���;#ݡ ]}��zj����B�~��}��0�����j̤���&_���<�r��w���9�ÄZC�W����\au�wN��өJD��F�38e�n�{�OmML��On�����D�b�!��g��� ���y~>�wPI갻W��tu�k�7<�w�˜!��-mb+ŤIȸuF<�i�wH�Ct��Xt��\UF�[/��+ù�/h�e��՜K��z9��@��ou��,������0)�M<���=uk��y�"''����J�Ky7{�I�L��z�<�����6�Fi�.�0����.�u��8+����Q�-�̨m�Zz����e"��1G4�mC�B�-��8�!3mμ��.6v,�_9�0]9%���TA��:	�]Xn1F���滽�&4+� �7���(V%p���n�q�;CLf��ط/.�w%�>���4�M-AcCB�E7�:�i���-�އ�K��TK+�"t��y�Z�̡��t�����9��bM�.���I�9K�p`�����ݳ"K�	�,f	6���M�|d����W�]H�C��`U��=|�[�ԁH$���D�����E��ߟ��\�Ⱦ�
5�bK�^5�^�3���q�λ�+)�wK�����Z_���b �:OJ!c�&��"�ג��e[,�-���:cN_&���~����ɧ�=q�� ��G�<?[�8M��o5���R`��^�L���r8i�碡�ϩ�)�`���+�9I�A��s=����ݪ���{d�V�������B�����I����R�)�:,��£!���~u=A���ge�X�/��aqly�/�f����P�>��[�4�������7��/�tL�<r�z�C9~	��4,:/ Fz3�_� #qMg��ڷ!�j��es;)��MfX�Gn�7�߮3�k)�U_q�P��a? ���5Y�-c@����%a�'&�]k�dȮ�gX �&Z�~횐�۽[�N4�']gۗ�:�3�f�Z�n�m���a��hU%�,Ӯ1�dκ}D�.Y�����-����"�k[�{����˘-b���79�Z⤿�y���󆄦��C}ֳ������]���������6i�m�����F�VVO	���b�W���[�.�ܺ�\��yԖ�)7ɬ�:�d��Q��O�֨u�\���Y��I�,�V�����:�PX�4R%�y�\����5��wH�>"�*��g	�}��):Gdp�e�>�3H�q�<�(��v��3���w/o�4i,f!�~�ђӹRy쨦����`sOiy^Fh�Y�E��[g-m5��x���!���hp����%�ԉ5��*�9(������r��`�8�A՛��>a��^�6�H<ֱ@�l!��6iz���(}��p�N-.�����XltjHn���xWW0����Ӽ}�+�a�$���օ�|6���0l��08Lٞ�m4yal�Y�\q�/`wB>Q�<����=�.W��1Z8�c5w}<Cؼ�6���R$��Z��Ûq��|
m��@��U�\&���:0�'����n��ȉ:���a�57��|�O��8�okH�޹�S�,}J �E2.)�9��~���3�Y�q���ǰ��
%�2��	�<�Ĺ8ʗ�Z�4p>�z��`�2R��F��ph�͛�jS��jԝ[YA�f��o����̠���ܬ��Ͽ�_E�>��g�H�{�8t�25�i��V�Υ�wv�7J�P�iJ�I/��~�@SCAM ��[���W���E��x�j���߮a~�H˷E#2A/@r��IJ]�(g3q��U�۔6�0��� N�u��U��}2Ц�3��/v���{hp��^�iܥ��:Ý��+�p���qB(��i��
YK�}� ��>���
��,�A�R)����)u���P��v���+(���Bk֮�J�}͜a"�o�ת��O�4Ae�Zl4���k��h�y�k"y�[9�>%5��}C��%����voyC�@]���3�VQz<���wh�4��aWRb��
�x;[�y��� �_Y�x��\�϶�P�"Ϟ�л�f*�qYZ���>%��o���s�,�u5�ѯ��]G�Acآ99�xb��ѽ`Y���i�k�7z�����o��>���uǘ���P�M���r���#�a|�y?,q*fSLqdp��o(l��C�B�M^1��[`��0Ä�70)��Ys��VI�vތv�5�Р�~�NZ�Be@q�ކ-]P)��`<��x~������U���ZTfc{�~#�(��0�\S�v��|3 �D�]w�j�����H��TU�"�3R4�����|����}��{�����ڼ8&�ap�s��ט嚎�]�p�� ��b����A�N��V_w<�>��C-44���9�̳�_`�x�aq=��u1t��ZXylVWJ�d��H,�¹��@�m�g�ݡ|��G�|cH�~~��'�x <^��P`�͒�p<ҤD�qں�x�����b@n���
d��`��Y� ��Oޮ�M�ʁ�b�d��`ٍʲ_��N���2�^z�h�5I�á�rԧ���ɴ7��O&�l����T�y��s���SL��{��]�D	ތa1���5ÞU���%���|����S�Ζ9���H�Ѐ�׼�\��)�jBSߴJ}߭����s����`�S�'��3m�_�:���ٙO��!I�F�Al!���b��޲w�}o���Ms*�0���點�/V��E��2�0�7u�촥�=݈К�%�)����pE�Zr�I�,���a��\���B�7��[ͷ�m-��#I�V�����zhF���l�h^�#Mn�(*�L�X�����u��^�Im{��Y�h$J!߼�`v������?�!<֌pnj��ܧPF3;чvb��_-B�<�_x�����t_?��P���u@=�l?��P� �K,d�K�Q֩����ʉ�{Ɠ��g4�\�7n<�	�ݏ���\�m�?ď��<�i4�֩��?6BJ���j�mۚGEG�:KҺhw�7�њ�璹B�y��6�VZY�J�s;��ޝRg�s�]���g��>�O���CCM����k�5�Y����-��V@Z�+I� �4�<�5�N!�ڿ�:����}��z����ڷ���ˤSʹ��ȓ�p�_��c݂5�vS�Y^���V92��Ή=B�q�eJO�s˯��WWtz��硓����ڇ�xtz��sYN�w��;�{fws`>Ѭ?*��|�q���EE����v����a$�r��\M�<�E*���z�ccP.:���ۗ�C3v�f������%���wz�p2�l�[��a�����:��pځs��������`Kk�x�k���/��Jz��򙓼ĭz�dc�å�FM�4�}���w	�4�� Afa��0w���}��m�jEqx,4��,y��g'���&�����t��æ@Ɠ�������d��]}���ŐZ����EDL�̶��Y�"��p��4�&vc���<�hOa�F�3��	��E{�K�M��@��O���-!��,q@f�nܯ_X�LO:�vR�4%,��)����+�r���!�dz��p���Gc����G���7�s;���`��R5��9��Z8��;�t3d�=�[u���� �hP�4>`z�ӱ�8 �^��A�ݬ���T*���w09�ϯ�����Fv�H�b�x���}��L�䭇�q���J�jӜ��w������zk!Gk�Fee\��*�b}�P��#��)i���{�:WbPZ��pv��ϯ����d��|�+��B��������)�WQ�^��w�ȗ�ƫpon_Sm�ز��b[��}�ڻTEl{�r�6z9��ې�{��½���es8k�6�A3GLѻ��W�q	q�^�0N�B��yB��M�9k
�����>�P�U߹3:��f�/��+t�6p�T+�OQaF���b�� ��8�ڼ�؏un�q�2�Q����7��Ѻ�ዌ�u'�˛�B�WU.q�/mc
;�ԧ�$+;f���7���w�1|v�A��	���_ �=�7u��\�;����_Wi�`��p�n�V�W[�����]d���ݴd��T�{�QM�,=����sPÏ#K*cc������}�m��`I�]-HM*/B_ݿ���U�7�>�d�4r��W�J/-^�`Os���ǘ7��5�Z���<�
�1�D�P!&������^S�(=fJqq��9�տ��d��q�d�~���r�XhK(2X�L�*�q�P��o��F:���w���i*鶺�P�h����Uk|2�^��zF��l%�t����`Z� �9�>l��I��9�]O���*��W���cQ��O�w�;�ǟ�fS�sYﹹ�8����i���k��������� ��{]!�<���c�-���"��=w��Q����8�x�x���zh����W��j����k��S�j_��zM[��i���"�!٬�cl���s5�`��U�\&���a�UH'װ=���w��\���n��h��E����{k�;�>�M���x�;�|�E;��%�Z"�Q�V*��y���D������[�(����j�MVB���FK0{��y��bO��D%�}J{Q��ř�v���<���W��Я�c������V_­��{��7�܎hn�Yi�������C%P(p$ך��pv:j(S��C��n�>u��^L���xQ�����$�m�B�S^��,�����=�,�2����q�OC��|�[Yq�7����3�w����lVG�_�75-M��|�O9�YS�#�ͅy�͌ҁ��P}�/�6I�*:΍B���A���b��,�5θ����L9�w*b6s�8Rg5��`[(�;ج��M�ζv�d�}"t��i���\��dl���p.U�J��N+��6�]2�;9=-#�
��]V�wB�uMn���]F ��ϳ�����J;-1�d�뻮rv�H��cM�)�8#�As��mB�E멃��p
C�M���H��5c���%�wc|�����^�z8�_=d�����u �^�+��I���sR=���v�\���K������:�ouoN��F�<���ə�X�ҳ���#�hMՍF���o�
�����y���s)؄�EmI.��b¬��دwG0��R��ur�,MA���[�X�/{��2�w*u0Z3�PΧ���H��zpU{W��q�hf�u�R1a�6�y��rɜ)���[�)ub�/�u�uL�x���U`hX�D��C���_e�(�b�@n<F�鍤�-�U�elN�"�q�=X�$�<H�K�~�]Iq��l�>D���q�}�u�R.�Nm�ȭo4]�|�+p�n��;]����p�|�;�\������e�Uݗ��@@�Q��
,�K\��KX��c/N`�jT�8%��v��(<$N�61.��x���E�j�*R��#�(å��;c33u*BX�!Ok�C�7�z]D.��g����Q��\��5&T,D�i�Kb��K�э(�Ј���K��	  4Sg��@٥îT.�V%x�3;���`�|�I�z;B��{��#gQ�!�y�J�q���t]�v�ï��p�I9��c׼-�W{�]�,����]&�Y����P!;���:�C��R��=JM=ԹU��1�\Vqݳ2���2��4&��G����s]Z6B�tw�&SU*ƭ��#S���l��{�j�}/OZ����`Ng�e� {����j;9�vT%�_e�H,G�:���TI��R�sj7ĢED�b�]w�:�WI�5�է�_K��榅--�ٗ����]w�4K��^evL�Nױ�U��s��I�m#.�=��3�;�G^�'FWކq-暆���c�U��s�aA�m�{(;�F�멘1e�t�h�t��L��g[R�U��]<ڊL�$t�7+��B�mC5ak{W�ҝ��(�5��8a[5�6A�WϸȲ��j��PX�㻐�C��&g74e����g�6A��,����U��I�X�5�5�7���WSC0%y3e=h'��a�I�Х�����ެ*tk6�H�]g4�]6�5�;`N��kP[�ٝX��t(L�M�8��U�Ϸ\Ы�Re�-��8 ��Kc�s8r��wK޺���Wvp��X�i�aA,x�_W���%N�Dms\����C%U-F��Ovۧo8��8���6��nݾh�A5&��eF��HI��y�o'"�͍y�HF �/Zz��n�����8�Ǐ\q��]�v�ւGR�HB�V�~|��{��t���7BFUQ$��O|v�N�x㎜qǏ��O\v�۷�r��P7�W;�˻���7���E˻�^ ��Mv\ع���׊���Qr�s��2.n��x�^˖}S�n�wb#��[��������R���4V���r�wn���nl�t��W'�\����S��n�;���N��o.ur%�q��J1yu�>�A�����^S�ۻ���.��/^�}��7�ќ�susx���
��~�����u�Q�  ��<@4|Q#\��h��%�
J&8�m4�LG"O�"BIp��n�$��$���IDY$�LP�ARM��d����e�pV3��J���sͥ���N���(a�M�o@�^Χ};a�핛���'VU��1�FRB�~lE�&Dp��,�A��m��NBm�I�	�_�Cj�����>p��Ɖ��D���Cf�N&�()�xBjP�* �(H� �A@L6#�%�Ƞi���G�|����8��Ĩ��8gk����Ʌ�x�"��aQ��]�N	:�ŔUa�(��k�.�!Ŵ'��^�	�հ�3��zF��'XĲ�1M�]�Ў�x|=��m���w��/�~���<)YW���£L>\`v��I�O�"��-1ގ:ٲKY��O$����@҃����k�SO�1ͷ09�E��bm��;q�r(����R�/��_9kѾN�S��k�h�#!�o�y�ck=��y��y9����V����D4�t��J��_��{�Z]*]_F����; �*�3�I��X�ֆ�����Խn�J�}��~�Ozi�QBdKt�ݢ==�k�3^i�u�?T�(_�\#���y;��Mb����x w�wU�|���9j
�T6z��x�}�T�u�r�i���ƿ�ڧu���S�~������	���Z�g�p�K��N�&�=���?���F��x�O}����3pn�l��"8[N~�߶�=������[%�ӂ�K��9Ѐ�!�/UŇv����78�.kz�R�Ń�oBOI4 �f��)���\�1��/�}g���-������g/H7�~-����e��J�m��"EV�kib=zof�2����#Ԛ01�F��{'l�iYp+\����qӟ3�垐�w��nC�eio�7R�a%�Ve�p�0��仜YQ��T�mΠ е
s�\9��{-^h�:��˭y�s5u/�}u�i���C����k��o���7�O���������=>HK�z��Zfg~t^8��{'7�Wi��Uw|�k���,�����q3g�hU�A��M���(=�7�C��Y3��wg3M<X���/���oA�5��^}�{`�G�y	�c�sW<'�ܧ�?Y�����̼ה�߭��5�[�]b��Gz����k�|-q�y
�X���Η;�{e��/�O==��j���Vk�+T>v�!z�����4K�-����笼�+e���~)��]"��r�c�|7 ��._�Ty�p��0�摴6�
���}C�Cp�^n�����-��{��B{k�ﴬ�뮟oH���I�d�Ӂ�|�<l[:=���n�j2p�`h�pu���b'�]�M@�&�z*/������A��r%c<���t�j�P���p���:�D<2ס1�.�Cת�Q���V�s(uμ�sc�����ޙuͷ�����I�(���~P!oR?������.��)�ct
-v	��*��O/,������8�����Y+9�Ƕʭ5�>]FҺ�o~�ĥ��E���2,,Z��t���?{�Mc�tWAy����^c�5D�.>��83G7`$,l��w5!���T����DX��`
G�&��[�t�h͛��F�ƃ��Ǜ�|��]�����VB'>ߍ�/�u�A��A^�1��GV�P��3��XnV��eܝ�����.q���������믽'OR��(4y�A�
�zzScr|�ϛ�����u�|^��O�8�	��
)��v����u>~m�ø���EzD&v��XBz��=����m��15���� T;&��3�侵3�"]�6K���#�!�8wDѺ�@��K�\{��To�ל�|�̾��M(��4�O醐��ۭln�U�W�����ͪO�.yd��(hxC�y\��U�3�׾B�����ݹ��мe��.�];�9�W��:+%Pb��T��X�u,�f*#1�ۣc���n�<�谒ܰ�i����1�q���׃��B������G�9C�BW���_	���ɟ`����d��7�V�o�y����x�_
׳�gԼ���v�t�ԥe1�����1{���i�7� �Fp��zS��.Z۟ � ^Ø�~��C�7�������ɖ�Q���V���x.���nrs:k;c%e�w��Y�_p=x�0[\�:r������n,]�X���Z�@3��>��*"�ήQz��:!GW��(;v�-Ƀ�1DP캝�jd���P�w3%�;�qƦ�#��G�-�T^k�֘"|��8�y��Ggt����f����9��`l��33)	��e�/7u���W?pHoز�Iy�s��=�_kI���?�k���C���n�fKH̩<�T_��?hk^���$�&=ܽ�\��9� E��s��=M*/B���w����g����?
�dިY�n
[&-�E5oRC\v�ዧ�x��#��A��C��_����L�-��o���'���5w�u���W7���ʲ��{ml	��X0i��e��F��8Q�]6^F�J������C��,W��K����\�=�K�'��rûju�Sᆑf����5��t�ɒ���k8lOއk�s��O9��)�f���lɗ�<B�3R�z�ٓ�>�z-�XzCM��Z�=��D�}I�bS���R��s�"����ɴ�-���Sgz�[9y���>t	�ܽTB����!!]ϥg�,c�T9�/�樒_zv�	ő�w�+�B0Fc�N�;�	�bM�D'����*�F��4 G�}�>�B;���?g��sӟ-��T������Xb�n����y�9-����GK�j�-��N����+�O�t�<9<��9s.�J�1�K���3:P�7�����'*���e Uˋ��cqu]_VF3��V)�8n����?!����½7�p��mm��3��>s��\�nZ=�v�d��#���;M�u�56�K�&��`;�a
�k�"�і�����,�����]�'"h ���f�Y�[�3�W�Ot�h�R-��87P�tP����l7#��p��� d�3�]V�ڻ؇ӣy7zBy��r=��8��b2��B����c1�XV�^~�=�<��vr�3��[gN�k���l{�l���׆>!%�LO?wBa̽���J��oOV�^���P��ցJ�.*HE8�{�	�������E��,�����wN^���u[��#z[9E�<E��r�,�����Y�/����4��躑�p�̴YiS�/(��׮Xr�n�xe�Xhu(8��6�zh:=Ȁ9��09�;zr�%���n���n�"�l���*/���BeC��r������>=����g���ƛxfmnw�O(�9ۄ<'T&�z�������P�A.{ M.��!����D�ecy�o�[�����=�@x�4Ķ��`����1��$�/u� *��L�a
�޼~v�(m��V��.2�/o5.���+{�[M�K=�4j/���<��6}<vtg����Y���T0��O��_-�p�p�*�'�o�8���g�y���������UĬ�<�N���������?�y���8��~쾖 �`�Bݍ�O���A�y�W���O���y���c���K�)��]/����@�\g# w��~���/5Þz�ϓp�d��w��P�5u��v��#V3N8�/&���FW�k�b��E�����]ߐ�p'��~X"ûu��v1��[���mԳj`���Ԧ�4����>�/�/�7W�|��4���PZ�:�:���t!#^�ׯ�^���{]u	����y*��R]ċȴ�o�I3(T��b,_���V[��s�lo���@Ү�l?)J�n�}~}����X����;y�n����{Za��v�,���J_i2o�$��_,X[��'��vF��ϐ��Wե_�������_>wc����9Q��6���Ζ0��xk��<��a�.�c�T7����uB�3�y�N���9�9�7�y��E�O[u[,�T*�>5�[Bz��LA��z��������A��"��ʅ*ҷos(�IӼ'�;�Su��|�s���@;���/�<Ř�`��s�ݩ>(�ٔ���s���5����a�^��q�sj�#*=��w!QEX�-�3\/�9�e(A�C�汫53G�������]�rcҟ]C�aa����y)8��K@y��s�<[wÈ�f᳗����=}�!+�}��<+��׍S3׮P�İ�?��Oà�ɸEĂiWs��]e�����>��6����<�b�]J<�ۣS}N�v�����@�������[m�t���}\��ޑ��g�Ewh�J����p%U���O��[��c���Z�$Ķ��7��-H�s�{]]�g�i�^'��G�XTZ��t�;ǅ�(����B�Tx���	����}N��ݢ�~&{���6b+{�=�1m���+��*����H2���b �ƃ�����z5��H��6�Y�|����W��]��̵�LzJ������8����֐K�� '������f�Z�,z�ɇ��.�{=�.{ݒ:�8$'3L
�<�U�>NY4��� xg�`��պq@ތ�e)������9�sv�2Cc�9j���vM�J�E�qY]~l���c�/�&u�h��c�8SK���7����3++~2�ٺ�f���yK�_;������/z��9*ڵ颓��J:��P���VDT��+�Ē.�Un˭~�|}Ǔ����VT���C.��8o+WJ^�W]��]2UV�9B���V�}��i���V
��IP���u8\b�NƵڽ��;�`C���w�k:�s��-*I�(��Ӛ�6����
uw)R;f�'c�N0��S2r�z5�g���X����(��>�W��p�q��ܭ��W��I���e[+�W�򤝎�O�X[�5v��h{���>�cuQ�Y}��1�J֞t���C-�k
�>�Y���3���XɁ�!���gtӐn�ך�v�I��l[�ύ� ��qx��W��
�E�5#��Ǡf.|)�8Bop=��̄��R5c���L_�E����M-o��2� �^sVn�����+uϟ&2���tN�<�+V��[���ቃF��k�q>���j5�k./ė�u�rg��\����:�P}��Zh�t�6��3cq�Y���%�L��'�5эi���(5z��nT��5�����Qh�u4��cz`���C-x�Uiك�zn-�k��^�ҁ��a5C0��Rjk8�ehP{K�%Pu�W8�e�L0�wq��nC�oo��k����З��#Ok�!C�foa�U������s��z�
�K)����<0�� A^!�OW:s��K'��f-g�+v�p��7�)c�S�%�{��I�Иv�o�:keAEAƶ�B�d���KU5J
����^U�Z�ˢr7����SM�-A�2�Z��E�f�RV�Uh�<l�����{�
�!Z+��λ��HH�������T�U�c�o!�����T�4^K������õ��)�����c��v{���{��y�K>����g�G_l�+S���@Մ�͙���Q�*��ȷC2s�u�T$D����[�\�ͷ5%�i����k^�*����6ز��9m!,��MM���nU�a=���Z ���?|D���N��P��p�Qn{�����wh�X�W�����8�Z	.���Y$�����}�$!�VB�Ͻ�2ۦ~%A=�5m�بb��x,t�`c޴t{�>�t�� M���Zy|���GD���oDF3��r~t�����~/������ꐅ{Q�4���La�Ƽ)��0<>�aT�mrܿ-�D],�"9=z�. �H���"گa�C��PT���h�����1L�ʉ�O���yͳCB;��xcA�A��v����|dO5ީ�^�T+����1���zTg1��77�������M���t[&{�	i޿@k����%5i���Ҙs(��Q��v��ߨcyٙ���S���Z���!!�0j�.0�b��Ǣ��>��3��A�-=��u�m��,��Y�`2��)�.o*��绘�k�Š�D֑��
蟁 �|׾�p�&bp�u�dAΙ#�OL�%0�q=�E����
Iob�N��V�4���ٵ	��z��/\�Y%d������8v��[��aZ�J�㝏'mt�%�[<��уt��y
��*]p/�EB�V���K��灕�?~�Ƽ<��ܽҢyU��������9?p/�[�P�y����a*/��.���1��~���m;��Ywt����cAQ|�wBe��yP�ß<��f�z|^�*�U`�B��7 饏����(G4��uBa0֑{ʅ�]J^���P%�}�'�y܎5y��e����i�tE�-�����ڎO���m&�T�������n���u����̞�rW��k�e����)�t�d"Ys������V�:������c=H{Ť�r��m��'���}�	]{�h-?x��p�'V`�	����-}�[�q\A���qx��,�o5��ϸ%��A#x�OB��!�~T�2�e��F�_q��.s���ܫ`��{��ŏA�B_V
_Ln�|c�G�z���__3<�m���2�Hŭޅ���*����w�A��}��n�<;��Ilhx��v�g�����K���ټy������Ȱj+w�Z�u`���b�f�7.�a̸܇p87��4�r���7Uoۑ��2�V#��A�|�S$�ֺ[��YM�Pyuڗ!��ui�����el|�����B�B5ܭ�鎷��K��f4��ˣ�Q�5ñ��kV͔^O��慽��1�ǧ�d9P����դ��6.�vswR����܃�`�ՠ��b��C�7�c�h�R�}-��/�9Q�Vc�Ţ�6�ջj�1)r�=�yx�[��BU�\!Bv������2np�(VG`yp�1�.I��Zs/�^N��+{�8�NW6ыbyKe���������O+���(ő��;y6�H%t��u� }�m;��Of��<��Kw)r�3����w��u v/yƉ]]���YD��m����8Lͽ��5~·n��c&cݨ��S���6�ڙ�&S,�h({v��+�����kܸX����N����^e����.�[���	��ۮ-qG��Rmtw�~��u���r�3rFf��2��J�1J��)c�}�N�s@�㜗wnpC����7n�7��-��%�/�����fs�3��C�Eu�+U6���Q-6�Jxv��6u�S'.��m�ū��65��m��+8�����p�[��8�a���VL�Zj]��rT­Uö��YQ��,0��=~�Y�aWMʿ]z���vu]��z�W�w�w1��������l��r��C�x�Z�u�t2~5��B6���r�i����g��j�u���j�(:K(�?1�Etcs��p��O�"�6�Ф8���z�m0������;D�b�-VѾ>A�@�&�.�.0�\�Y�m�̋ڻu�k9U]�s9�F�ǲm�����U�Ö9"�2�������W��7�-���2^��aU�9�KH���L�Ld��v�+�v��S�P� ���umG����NvG�^�2\O]�@t`�n����}ٸ5M�c��8r���8T�ڡ,�TT�w��u\��'}J�[)�;n�U��y�Q��k���u�i�M�8�p��t��X�)3<֬:���}����ژ����WK�n�-��1c�wf\O]i���䨽{�8��[��8�^��Qԕ��'^NZx��2�J���)�`�ك��f�U�$�l]�e+U�ն���VWlk��]����u��Y��U5�
�4� ���դJٴ+�8�<��p�TF����u�&i]%6��ή�`�ݼF�\�x�Mh��O3��3:�]�Z��yO�ࡧ~��r+�ĸN]wI���Fo,ݻ͜�
���Sq��R�P�p�!콖��'ٽ�"�le9�>2NΝ"���<�Ѯhv�<ya[����ÓѼq#��ӻ���#������2�m.1M<Ld��\�k}�n�66���ۀ`����+����:j|�;�v���U�I��*e2s}��%0�D>�^y��wt���WwoV6�I"�I#㍾�ӧׯ\qӎ8���i�ݻv֍B2I5(�$	8w�E��0wq|��
����'��!�n��iӷ�8�q�Ǐ\c��v���	$�$*� $��y��}�����ĒI$�y%')��k�];xӧ��qӎ8��Ǯ1�ݻv�P���T�8gp�}�ӻ�t�n���{����Ly�^���췀�i�B$�m�:g��ö�(�t��n�>>y����s������wx�Ν�;�w'�/^�MyŤ<j!!��h$���m�8Bi��W�$�e?�)$�	��e"��HB>ex��S&T �R_�h�e��$�ʹ�@�BD&��=��A�����$�_"!����a�x���P_�D� �F� ~��	|�\w^�]�����uq@��뱢���;�D���	�tE��H�Dg���Ѝ�ߜ�D�a�<M p�4,��}�9�X�Gx���ټ�uUC34VҠ�꾭�ʓ*f-�(����������A�z侨�!�����<�a����9�ûo_X��Ͽ�E7��0������]�+�^��
��1���6�bQՁѺ�1�㮒�a��ޜⱊ�9��5�X�a�-!��q���w�m�n��p�#"����G�p�ۮ��=��u��uYZ�+I��!�~B�G�rK��T����3�7����z�+�����ϖ;�E7B�\���;�y���6��8��[Q��uCP|�z��:}��S%s4#�>mf��Muw>:�e�^EOwR`Z�@�P��z���ѷ���i ����<�~���nsȮ��>r�9O\�{��An��5ε�s��&:�_i�fWS�\G��S .ƅ��xu�;����s/�B�G�ja����_E��F�t]<�Z-H�b߼���I ~��=�W	{��w�H'�*-���[~�4���D�B{��{��_$�uy}7�Mz6/+�RH<p���u��-�_�sY���z�W|�[�xj�by��^5���_�����H�:��Y���}�hu<s�Z�� ��Um�E�͉쭩ڜ�H�л�I2'U��$yހ]�5wF9�����#n�Il9�����u��>)���� 6�#wazv"�3E+L�M�a�ڳ*ގܩ�bJ�`r:w��:q�z)p�(�ב���}.�������\���y=�|<���'��0fl��es�|�i��x���b֝�OA�F<3��V�Y��FoqMZ'�e��
[k,F4���@qw/�f���+U�kGL�d���:��1�����{Q<H��d����ߢ{�_5F�z�����A��h ��35�;�¹j�Q�]Bő���NZ��O6�kf�Qc�&��0���+�[�AN����|�}'�/�˵��� ������]�����"@v~�۬���R��`�Ň��7j��8&1;�`{�����Y5}ܭ=��n��۝�#�e@�KݖW<��K��^��Ѭ^���B}���lƅ�8�rè�s��ֿ>A�=�-�v*��XK,����뜗�p1�,�q�����w��k?n���3�\�?\,x/���_s��P/9kow�6��;���FͰ�8ڸ鸇Y�S�'0n���ށ!�\��t��%C�g� �t�Z^9����\��b���q%���]���j]�D�a��������S��E��_j����̩�T�u���R�+t�����o�>.@���mJ�S悢�X�����2^�k��v8����N+�L��`n��˕�6��N`]�
��Q;��S��� [V��;G��5�� �4Ey��Cd��eM�v��c�;���m��X�����^�c�f�?�𝂿lJ�\<ciۼ��c:q8z[\o�A�`$pJ Q�i�RUǛ���9f��[)�W�N��e��n����^�4pp}�#W��*a�A;Fa��t8��|)MGz,���a<z{�Z����t&T8��0TH1��G���-<����Wo���/b����6L�.����:���^�s����
��U�=��W�%=���ӟD��}k�7��j�5fsv��v���㛪`��W1��jF{^��{k�G�+��@��� ��^��������=���G���J�H��:G��r�S�r�F"�X�\�h�t�%���k�{R�p��|��#~��Zh��%9�v��1ٲ<o���LJu�K�����]���21�f����6�@ZYy���|�]1��|�q����t��%�����GHzT�7i�z�|P	~�z��Dg�;3���3��%h�}�-8���z/�x�Tؾ}��6�a��y��i$�[��v+,U�3���f��!CQ�4���O�b.}�,��b��:S�ܡ�v�}$-O�b��ܩv�q��[^�����%+*>l�	��k���`�3e1�r�W]�x��J��<fvW*݋n��eqxm稦s����>���3��৻K��>*�">�+�B��}�Gg�[�r3,��iY�V�$��wbl	fE�3d�md�l��;}+,�tP�l��N��=��y��8���ǳ�ݾu,�8��X�t�� �OF7v@��-��@���&��#��U�|�<��U���m���4�{|���ƅ��̥m3��,�!�����>�hэ!�	-Zby�������:�yՃo����>���L���:��B�<������6���E�o�TcK����tAF|�W*�w��h=�(ք�v�)�'\�2}�wմ�꾡AZ�5O��š�.8���-���N5��2�����:;�AQ\���*���Y��UAA�L�^ý4�F��;�/s�#i�N�=J�Ú1����<fS&����An�L��eC��8���z�M��U�n]�u��$	�����A遧���q������R�/�YE.�K��c�� =�M��2ǯq��VĶS
׈�����k�>�m}"0���(w�&��~��s��� Gl�k<���	��6-��\9N����!ٲ=�p�S*��P�\��9�a�7�Э<�i{��>�z*Hno�@��G��48:�x=�G�'�yH���ǽ����y'�lao��e�p]�Z�EC�(u�/i�ǫ!�i]���A{w ��Ѭn2��0�X���߂����9��,�(�n�3�l-�me���b;�f�Ѩ���Q`+V�Y�H�:��]�S\{á�$���^���|�ŋ��;��Z!����o���zZt������m#�g���FB�^� ���P�'̍۾%���I��n��oV�	~bec���X�7O��|�\r�����D��ř:@�cZV�m�a�ۈl��֐7U��m�1}>b�v���%��P�\皐&i�W�"��Rkyc���O�ՐL.zf��;J��ӂ3<�V���|�����+���츆�n"��~��`�������`��_��oO�N�?o�$����a{�Z��=�}s�o��O�H��&����muN���9�67.�׿�{ޮ�+�FRk�>D��Aa�+멘d_��8�G�4�W����3k��o:��]�Ͻ�(����َ�VV�F2h(�a� {�^k�7��f[��:F��7��������&����<�}�"��r�kk�s^c�p��1���|��^ yy���*���Q�G��d���H�%�2��ϝ@ˬ��WX����O}d�&.K_WU(�U�yӖ���B�>�A�2s�:l�=�w����C`d�8Һ^~{l�>�!ԟ��쮹 �T��X�"Ej�PV]\2����]�
�"ɣ�u�[�f�Z��h��j+ay�fwqN��TG�U>�1�a�+���5�$���1�)�㙘���Wr��Sv�mi�T��;B�L����I�2���&�t��xy���=��z�$b�v�[��0���{=�ޅ�ƭ�W:���`��M?t�ٯj�o��OӜF-�` ,<��~�ꡪ}����|XQgqB�#5w�U0�Z�s[n�Ĉ���k��U�E�qͅ��u/�}{��)b�}�o�g��A� ���\!��H|�>[��J}ݽ�e�xӝ��;$WP�Sxl�n�Ҕ����^Їm�a.��3f9��1�9^d�5��cw�����vO�,�����87�'3L(��wrF����v���e�=��|
UK������;�G�e���0R�\c�AlJ��J5���GQ?��~u} �Z�ʝ�[\� A&�|�c��������Pe�`q�j������>��WlK��%�S��I
�c�p�p��WyT5}��5x�O�9EbO�;!����+}g�)ъt�Ӣ���j�̱��ӫ���GMC����HkȺg�0-��|U%c�W��[��|6�#���J˞W�w8
�k�-M�r84�0*H�?���|f��T:���;@��3�TZG(;p���L$P��Ӝԝ��ᵲ�w;�E�`�øx�՜���f��M�NFV��V���ثiT��ZW��m.L��5\��ʼ��r��	��9�^�[�)�}���X����\���a0 }�{��>5�GƼh�!�������'�������C�L!{�"�e��$S*ڶ�鹇l�����U�e�/�A����}بWGIa��ە�f�!��S�S�ɥ�s�R��g�ޏ\t�xa�z\	�����7�~�����B���)����w�f����u0^��hT��M�=�3������}<_Xc��Z|~���n�r�*�R�x�'7#6���3F:Gdp\wv���
Y��cXm�<���-`��(�g�5���9ޝF�����k�Єi~���~�}ng�iyJ��e؃��fhC��� w��*�^���|+Z曚kr�|q�J�U�(�"��Z��{�t&\T��w�aĝ��l3l��O�ȗՋ�̕�5����:�*D&�%8�.�¯�����	����}`O��y�R�.�s7�����xV���ts��sBT�5���U���Ƹ�z�~��)�=ʜ7�R���m��o:�;:��M�W��T(�)R�!{+�k!�8�aٺ�Ä۝�'3Z�8���%<����R�j��t��:`]t
��#�pk�i�o��q��PZ���9�^"-{3��-L�):��tXyccVq�:�K���U�ŋ�AZ�$��Ͼ��g-�{u�>�o+�`��Rbȑ�;��9{�MJ�H<�d�ͱ�hvL>36lJu���.��ǍW�z'{M]0+/;��Nw���H+a)��%g�eN�*�~`�/��zｼ��ǜ�/�b;����q�-L����֨��G�|<�SU�_:vwϔyG�W>,<��O:H�w�7=Bg����(�   ��4��k$4z���q\Ӹ6�m;cѷ���D���l�����yC��������HlgL�쎾�[�O9�85l�i`���͑���p�q�/�*��(�=�#2k^:�R)���E�޹�Z�	(V��6q�ov>rʃK�q^=�:�z��EO�;���a�LK�L U?67u�,��~���#���P�|̖��s+u�WR#nRܼ�x�>��&gְ�Ǉ�9��ʆ��=��tcH|BKF����5������v5���4֪�ós'���&6&��v&b�++UR��Yz��*sI^l��8����X�U�ѓg��!�x�\��+�k��
y�kָ>z���U��/.�%W+UU��߷��jQ7ntB;�wl�"ϥj��~ac���s��n�;U�ۭp;�ׇzn�ܑf�����Wx%w��Bk�01���\����/@�Z���0��g8�yI߷%��Z�`Ø�Sm;�7�� {o����a9�e��"��χn���SN�#;���ǺL6��*�]m���N�s:�5���qg:3ܖ���Ʊ.Qf+�<իt�� 0�w_Wwu�{+omc�N�H O�>?����.�_<9�v��$�I�B?4z����!֟C�~���Z���Ժ���溙���������Y���;.P7@]xa��kWߺ���v�p�В%��d��z{]�v��d6{C�ql:ܵz-�|g\�(q��a�.�@ȇ�� 4w��?p�ep�֕����m����P=����"K�gc#`3h.P��
+��<N�c�iؼ\�:�.�u���%s�x�z2�7(G�9MG��a���`x.��˵���̶���:�"v{���c.��Hm�ʶ�v�~O����,��_?��P��RZ&�m�L9f5�(��gA÷���� =[Ұ2|�thMn�k�r�o���8�v���~|oF��f��.��8��P�>��a���FL��^P��.ov��wC[���ט���w���o;?�\u0���H�}��/��Τȧx���,?)��\zy��.|��z�+���i��&�]<5�D��r�aA�z��Oʻ���h�2Xp��*1<���T�>�+q~*V�9i쩇�i����J��:�LC�m�y��ŕ�u�nio*���:w�l���J��ѻ/�� 
�@�uk��S3d�wOP����ݤK��_J��e�U��n0T�	r��kB�s�UK��oQ����h�7�y���t��+"Wl�?t[C�\V�I�(��<�Ut|j �����}3b�m�[�r��m����zc�V��(�\�k��x�˪��� \�s=m���m�qb�L7��³�U�S
��B�t@�j�Y03���X�I9����O�ehW�y%�a��*9��u����[p;`AL�{h�CJ�_��낥�٪a�.�/���,�ؑ�.��o�c`!��������}\�F�"�o��'�e掵� �̈́�b��L��L�s����{�qY=�ޑ[o�Afݵ7e�U���]�v�s������5�x�Py��vVɦ}���ᙳ����G?'���g�Ӄ2P��S�F���u��AFB�ix���᾽}���L^%x���`�Oݥ�fU{�h����U���&���6k���\�z�x9כ�	leV����Q�[�`l��<���K�%�����~�M��^�p��Oi��fs�eq�Nz-���h="<ײ��}U�����E,�r���N�[���ݼ�E����%D���ǣB��i�yp�VvVQ��;S`�1=ys8cͧ�7L��c	Nk����efX.�'�X��,M�s3��{BkQv뮠`�IE�����V�8��,uqx���f��]�n,��کH�� ��)'J����]tO
�+Z�.� )����D�~��W��]��7'ؾb����wK'J0�ޭ9��[��M�6��L��{�@���&%�R8�j�4��<z�<߆s1yZ���Wײ�L��Q�Qn�wH��}�����㮺��?:�	;�7Xᯓ�[����b#��$�q�"���Wt"���ƌ'%s̑m����;q63rk����Gt7�LH=O_3���UΑ�6���]e�2�v���>����+qi�u��:F���q
����ˎR"&fW�)xi۾�s
�B�6N9��f�l�k���#��a�a�|ณ2��ԫ��� �<�@�T }R��9æ�_�%�|��j�O
��^���Vot�n[`Gԭ'�q�c�����<i�oz�ҕI���cE�]_
e�Wo���[�6��Q�ݫ�M�5�"�!^���k������[��5�&��(S�ݕ`x][t�fj��b7���K��h�St
>#Ԁ��:E�i��˭ű�p�ȳlP�f��39��s<3��9A�C.��:IK$��X��gr]XۣJ�j�!1�Km��y2퓉}N�2�7A��ƕ�Eщ��z�ۡ�²��'�'!�*�b��Ĵt�N�ts�OO!�÷<^��|`�}�|-�	r���e�s�;r�\tq���sQ���p��ϴ�zS��Xu�``E&��!�cK�Ͷ��x��]ӎ^O;״YF������չW�����V�:��.��P�v��#���;�ۜ$��ΙM��y�6W�<�q+�L�M��C\����m�������N�x��g:elY��V�F�R���V#��1��p����ǲ6VK�`i�ʈ;/*��k8oprN�Ʈ�Z��qh�+gq����:Z��Ҥu��F;�U���{�Vh��<����p�۩MV����#�Wa���̒[s0;z�\b8w������{�����ɥ;���ej�ۨ�ٛLc�˅
��'P�ܱ���5ge_>�lIWq������"��r\x;/�6���n԰�'�5�=�u�N���Y�j!kq��`���Bb@ݞW+w}5��-Q]ͷ}Pt�zĸ�s�������Bv����W�V`�G�
�*��BR�{�A-Le.���I	=t��t���8��<x�_]:t��h�h��(�I4�4�##!'7D��T�B=�,%�z����\x�;qǏ=��t���y��k�HIA5M���ĝ�B��A�p�����kx��o8��q�ǏG���:z�j5�Q_:�'Oϝ_��&|k�ۯ���׭^1��w��H��f7w��{�ہ��M�&0D �۟�ݩ$� Dā����]�H4����d�7e$�whْa�\�p�(�a(�Ċ$���wh�"��ґE�VCA_]rb�L�bP#
���k�� ��B����R���шW"4Pn\�oU�����R^*�L�Ů����DF'u�`��D,Ȑ�dBf~���F�A4�	4�����D$xP1�Δ"%�I�1�>I�����|	! �I��"8�eHR)��Hd��0B.S�i�;p��tպ(!��4�˛,ﹺOwy�q��z��iH�Z�9t��L�p��{�ٲS��9�0���,�Sm�a����e@~i���(2I��qy*�d�L6�R��$���\*	@�b(���GA�D���h8�L�JrH!��|�Iʦ	��%4A��|~? ~#����9��9�2��,.vQ�����X��	u�M\��ܢq���|%�e�H�W?A�8��|?�}i�b���g�sUu5�z�����Ѕ��h%�	�~�� ź�aO�{�Us����6��e����#��B wV���{|�?-�_^�6����".�M�wJ�ɮ>�����Q՗������ϲ}r��<t�Ug�p�W�뙼�+%�ٞ*��4S1���z����GU���v)��v����K��6M�:���4Um:Z��`�|��DwG�hO\5�$�>�\i��hji���5Y�U�3�C3k:s] ��+۴2�_g���8"�c�8Z�Fk���&Q�n����J^L�����\�Z=�M�]���=�^qTi��LN���m��w�̼fR�vQW�~���l����!%�l�c�V�iӏ�(#mt�X�R�������W0�'�G�[�k`2������8���Y�_�ZK�F�L�"���h0�;�4>:8�7��O��oV%,s	v��5LR캞[ {J(X[�8�P|�4��=���sǜj���I����.\i����������޳i�o��>>a��{�����]�z�م�u���`�������4�Om{ic�x�NN�|���F�A:�y�h��ã��I�E��S��d#��Q5��� �ln  ��rvw�n�1��8I,��叀����@p�3��1Hp�uD�Ӹx�s9Ѯ3%�g�>��!�Ijf��E�gu+��#��q�@1f�.�"��N���U�ƌң�^�Rh���Ns���V��+��lMZ��9���LJ9w��Ѷ��=�ff}�V�@��
�o�ھ��θ)���s7qE���BI0�NjO5wud��� �8�^\W�3n�S6�:;8�4^[<��u�]�D9�2��ʽw��Ҡ�m�&�.&�]��?�hqYS�ީ�dl�"�}���}���&�
�vP!�#5��:�!���i:�+��r*i�j��+�Ot0Ϭү�`�V���v�����fQ��j뚏o�g)K<�T�l\�UӇC`|�V�[-���f��ںW� K��>O�{WL��Q�:v��o����w˵�+��l����.�~Rx�*\������,{
�%��,�6^N�/Fyy_V����B{�w=��<�|�G�����?uG.��xnd�u�� �Y�����X������X�0]:g���P�)��~���E��]��5������%�&<xn����Oa�۽�ɭ��H4gTn�vIx4���hJDwlَ��mlf����Jx����az0�gdK��:�͐7Oz�Vǘ(�H�6��;���<ԗ(5�\-�5x;Q�����͠m��)�i��q�]�#��|��4�Y�P�Q�����36PH��Vf.}��#|�@���!��L��Y�-��u{����l��ׯazzv��[5�>����ԇ+�J\��h�w|Űυ�U!m�d����3�ឿW����F�����W��T��Ɓ\�ow�h��)@}�� ,FZ��t^w]')�{Pm�MZE��x��c�1	�[�$�n�J!M��z�S��n�r�Q.X&M�q��͑}2�M"���٢�m�>�����+)�)�\���g���8���6T����N�X<��өK;�H=��XV�>��8Cú��Lg�ɯ����+�¼<�߁��p���w��Pρ�)G�;�hE\���3�9R��wyɵ)œx��v����D䵆�_��p��� Uf�+�f'#�(�L�&���Z�u��h%|�"��6�����h
Y�c��X�h��JsDL��3"�6�xxd����o�Q�l��t)	�5#�7���B-�?�uߥ�+�_�{}θw�	�<P���V���ׁua>����z���׻}�~�a̴D�wI��[^���,%c�t_6}C3oP�Bq�1�k^ǒ��r�i<��ꑭ�sK��&�w� ����z��u<�M� ��������BzѦ�c��H�6o^�'2���ش�n��!\C�FK)�z{`e���)y��m.�E5����֮�7S-�-/��g$�r,���p)�6�7f1����[��d������^	D��r��H�^&}��G�s�7�m�Y\�x����*ub5����ӻ���(V�ʮk�o;�v��z��'j��Hkge��H�&\�k�Q�����+���K��՞������k����zEn�AHeY	Q��\�j�<�e�Z��z�ǯ�$?~��xxW��Q�VC�!��>�^mC[�>>�;-X�f�/L��T��S��7m�:F�@���k?��܇��%uv鎞�
�$m3�<�i����2�s�Sy+v��c'�'��̩������+@4O��^���Lq:Y6�q���[�ߖ������h&��Y�)�;R���|Ыs%�J��\�9\��v��g���o�hf}���<+U;�87H�z��{��ؗ��cQ%���>Ty`�����P�=3���?j�9[� g\t9�ǜ]�M_f*s&��IHK��O&�y}F-ʯ�h��p�������Qx�i�Ԧ��y(��S��ݽAwW	����zߔ5XE&mwΆ�ʗ*&�f�0��w���� ���� �\$��#qQ.��%7���;�+��5q1.�HU����G��eЦ��8�(��v�T�t)�����&���%�Yh9�"���=�HW�.Y�c��vpf��<�B��\#N�c��wd �Vt�F�@�Z�UƆ��tE�,�Ms��ظv�Y%��au��Zt�j��t��;���p�]'#�ֈ;���	V�=]k{i�@P1�;����������/��7����r�wZsT`b�]���~��hh)��@(������+���w�U���r�����]�0�G�x�k+�nv+:�kJGe`�n���u���⥻�f���s}��od��r3��=��ћ��FYP3a��w�ޮM�
�o��\��v���/���a����D{���督dD�8/޵�"q�i���Ҩa�����]]��L�i~��ϸ�4�3�u;U���kݽ�0�
*ۻ��fR��uUx�_�;wB��[���9�6�X�[�*����aw���D-����R��QD�[���5��M��[�r���C0׊YJ=�a���-�+�uT��۝Ź�b�)�}�(�e����������9�B�Pu ���f@���,���Em Ͳ;o'6s1UF���ͅ�)�JGzU��^���Bȵy�Ŗ�4�"DV��O�3��k8t�3 ��I	�y�6�Izu������a�'�~�kQ��o1�
�����T�u4��$$�k+*�%���؂��_��.�m��7C�iȴ�^V����]��ia��re��;Y;���+Uoz����r�Ǘ�)��ܤM�f����Q�rm��h�����©���w�.�q7Nw����U�@�M�v���:���H����Jn(GfC䧷���,WXʧ�}��){�U�s1}ʫHR�����M��kW$��{q�׹ssNge��ؔ�:��۷b:^eNS=�m��Z��e�oB6���4�j��+�vM˥ք[������Ż�@1B�� ���.��s��/�z�o�-�<���	�R�q�vj�0i�[x"w�:W+/�v�*@H���̵��`�[l0~��g���q��}�����_�����~�M�nkܲ�ޠ������fH�S�
a|{;��(�~�*<mlH�]�ܕ�֔����_����Vf�Y�j^:��-�W�g�^���{�ply�t�;7����n�H�
�˩�Bݬ�I#>W�U4���\vߌ�:ހÍϛ́��Z�Ź�����7���'ł�k>��nT$`���o*�z��V�ٌ�M��碑9�)��{�>ϥ�Dq�/��\=Z*�DQ`���]H"u��Žl�@��b���L��}ط7<���P�tz��K�k�����DH?�A�^jn[\[y�׾�y��`)f�#l�e��XR�owew%QS�\�6��|��C�S��{\����=	`�A\�od���+�zv�+f��>26�jꐥ޻�a�� �p�q��8��k��ff�\��m���&����BJif,�~.����c��/�k:�z#���o s�k�-�P�-�)�jf�$��TJ���hO?�%��t7�Y��ձW*�����"��F-���e�D��qr%��P�x��侯Ƒ���T�s����+�;OQ�f}�/2�����U�K�������g��,rk��Xng�5Z�g{guja�F�
���В5�{�̸�X(0�Ԫ,����l����o/G�`�������'�����em��?,<Ѫ�觺Z��+�e�?��H��Y��Xe��:���\��ZS��EZ��ܠd���\�eٚ�h�
�3X�+���$�@�5�W��kw�!��(u�eK��Z}m� �M�F����^��9<���5��Aڡ-�/ut	\3-^�<�;'92W"�i�]��2u@�]F?�����¼��H(o�@����3�1���$�6ƥ�N]f��֨́�e�q�<k�
�y}��[u��5�oM���Mw]�<Qˬj9:���ޣu�����{A#�AQ�|�����u�`�6�<kt�F��ɇ=��{H(=��<;�m��\"�3l��0_�>@����-�|�*�����uL�od315uW��=� N:f�����a�i�s���uFo5��)m�c2L���'�R#���'��]�b)���-��������ߤ{��{q�ݬ�]Ϝq�9����ե�f����G�W�A��4��\�(Nrv՗�<��d���~��FGlz����/���;�v��ߵ�[U��M7���!��`Y���Y���`�7K}�o����e�I8�2"�|w�	���L�1���z(c��f�
ʧ���3��ӽ�޾E����@�Ze�{��cs�c�����7�5ŭUbrs�6X"��m��0�P�v�|�4���zZV3M��o3�{�*���oV0��Mkvm�r���l_WU�8��b�cò�`b�n�s{�a;ع�\r�gb!��������D�,b �&��U{����Ƕ��(p\DU�W��;�5�����:i�B��y���� U>�w�*n�GQ�f�M����u�LNS���zh�ϱ4�1ubpW,�1�4*���	Wa��*#,i���袆\��79���@����}��y݂��t|P�b䚐��-.�� �/�պ������*���rߧ�2E���t:�O��2����y2l��6_�u����h����p�s�d9��Z"��e|ڈk�j��%Z!ۮ!���@�=
j�r{TqK�������-�,4Nf��vfP۽Q�����H��
Q�=�ʨ@A��]�;�������ڢ+��wN�5m�%2�k��(~Z�!vz��/]����ĨB{v#�x�Tq�ʝ��u|�=�C��"+�:�O2G<��:��<��#>���n��Pąb� p=y�#�BqP���Zo�5¯��+z=I�N�|��f�S�#}�c%*;�T|�cѽ�ƙ#~����1ii��p�~�}V9J���`��&9Q�9t�';�h  �K�#-tc �X��F���=Z$U6s���uN�/��ӷt����p� ���G�\!퓩�������i,�l�ީ���f��t-R,>���yȣo�Պ�yc�(T�B]�����ĺ=Σ�M��A]��nu�^�ѕ9�\v�e&.=��t�A����q5�-�������!s:8ި.��&�����T�eY�r[C���\!�u:Aǚ��ҭZ/x�)�p.��ۃ+/BfU���5�|�6����1
l$X��֙�j]w*Ջ�3
ͦ�7�Em`9�O=}P�ie˲3i�'�����줙��wp�5WSEw,�9���ήsZzs�m�\Q��&��~�ՉK����k/�֫��u�����$O-j]��ft�z*_d'���u�w/K�z�=��Aa��s,٬vo�ۺ��G�-W٦��qF��iV6��S�Jt��K9M]�=
���^'�Aa>��g*���w�uܗv8!�.H֝/'tӣo�Hn.E�5�{c�e��de�.:6��'A���O����a3]h�i�sL�d,%h��*�V��'k*2�*wD3V+�]>���Ѵ(Bɔi��{7�]f�I�����0�����}�z>gJ�� ���EP(��}c���sZ��N��B �2�=l�Wvx۝I]��r�`�HZV]:S�R�#�v��u�+��I޷�3�!�f���Y��I}�����ޔ)����ݳ�su�����Χ�4���f�wCw\��Li�'���7&�n'�c)Ѝ�;�]X)����Orӵ0a���	ͺa�kSà霺��+N �Wj1�p��:�#a(�^[�-r�	vp5h��˸73U1>l����=Z�t�ɅC�6�9�ܫ�TW<���c�ᠨtNY�if=O8X,N� �y/m؃)uh:��{KB�RG[!�l��յv��M�Nk��vko=<�I<��nfYN���_�p̾��]I�����wdS�4b;�2\����ru᳏��YT
��a��wԆ�0���am y�JG���紭�/;����}o�<d�u�V�I����>�WڏS�S�*���N�]W�q�X�f֮�.e*���ݫqWRA'Y�� -=B��]�宥���udd����ˊ���j��Q�W�� ��ᙋ���(h����[x�צ���q���v396zG����w)S�]ӖU�±�����H��ͷ�������=B� M!x�_}�;�0cIܠ�H��wwǑ����ӷ���x������|���O���c�)��
��wrS)ݾ7�bd�(�z���;v��8��<x�z��ӧ���eI���HFHH�۹:�r�6$E2��&�oV��r�nr�������;}q�q�Ǐ=�t�����H1���F�"2D`ĥ�������V�\��t��m�u��^/D�p���]@��"��sDb��:�~+��z��wv��n�\�	1BPǽ{��Z<r�wD/��M��q_^y�("�L��
�
�\7(5�C��ZJ*IK\�ؤ[�)a�(�Q��we$��b1DQ����x�!��úq�&r�P$��Ń��&J�ܹ�Ż�� ��sκ�a2/[� ���q)7�׿}���߿w�}|�{�c#�H�z$[��m�Q�r�S�I_R����kGk�4�[��q���m3��5������«�T���'�d�Ļ=S0i¡o��2lj�qp��=@�y�t8�%m���O�́�5ҽ\��^�c�'ӵNr�B|�@��>����Ŕ�©f����g�;��/Rq��х�L�L�s~�F�[��C�{�C�ٔ�n�*9��Fܻ���^.��	��y!@����^\����
ּ�{����ʢ�)-���lp_ j�dF����dU�� �$a��yj+6xU8ʪ�4�ʎ������B��Fe*���./�]�Σ����$�є3�x��I��s��4� �SǸG�,wC�J��^xlm��@�׻�/1���9�^K�U�
z}S�%]܊�o:��cϦB�Sr�(G�����1�����p�k@�b;�=�����@�n�4�8�o-.	��P��n��]�?!3���c=9+�u�n�V����ZO]�۱�"*�+m��;1��E1xѷ�Ʊ����T!B�zg.N
c.�#�d�d=�Yx� ��V3Ho
`�%�1O���9XS�%,wV����[�n.�V\	[��B�w@�bh��T{�mN�<��̾�� ��������TKw}
!U��܅�zc<�\�G
��@��@��r�]�����u�Ḥ�b"��[�m�����|v^���;p�;�]er�kcE����#�S�\�m�Z�bZ�Lm���a�t>z7��|����Տ��Ft�)�ˣ��2s�$u�$|M��u3���x�_�a�)Di�ɍO*�N �{e��pp�Ժ����)8nJb�񗼞��^>@��u!�32�������88;�������ZT�$am>�x���y��S���o��쇅�|�Fz��d@�-q�Ķ�s24��9; �2�i��P�X�'[A���;=�0��y��=wp�{t^��+���d�kFԢ�E���d!i���'�����wQ��uE\�^ʺQэU1�'C{�m�B������l�����s9,�lòxj7[����Ix40�I��j�t����1��vm�R�Ǽ�z.5S1QT�,(m:�$��f��|�6O�{z#�:9'"�u�it�Lt(O�E��.�W�N�L/EvVl4&&�]W���w S�n���vڥ�� ��9��I���r���g�Ok���1�|y���
ϴޘLȵ|lr��y��q�խբ9v㋜��m9�Cw�oyby��;�����]ԹkNmt�?W�5���c��Mܴ\rg����87#��ïM^�K�F}è_AM䫷�d��M�[����gK�U�k��ıM[Yk�e*s���d�v�Й���p�5u�Q�i�z������|�U0�f���������5��2�>�����+�t�f&`(����]������n�ѳ+yſ��g��$���ﳓ�pKZ�;���$~<m-���t8u��>#v�t�!FL��'��3y)�z���v�f�I��x7�]��ӹ9�/V=.��U���Y�!V��mlQ�P@�&[�S36��s���z'vNir��ms1b�Mlu�C���^ruP��>�N�}�@P=ݕ��]Oo����ؔ�M��w�>�!�:*ه&M��R�WP�մ_{h�j�=�KP���ת�!Ȭ�Uj*!��i6�
�[�BKw�I;.�wa�D�k����jV�^�V��2�n7_;�>�b���]�X���O���f�7X�by�&f�.h�r��\�f��g��QsFL�xv�Sb�ݢ�Β_n1��FCw�����y���׻;I��j{�� `�+f˜��_�v������_eW,w9%pv;[x�6�+;��)T��lt��������v�����d}^j�nuܣ4�(�w}��Qr	m�H?�����z�4u��#	^�!~�V�+4<� ���滒��Ԥw!�@=���kӂǓ)�=�M�\�r5�tQ�3x=�W+�ɟUU�mi	wW
��,�U�ּ��ӹoŝ��B��n��5o9�h��>��`�P{��Z.���Z���{�Ȃ�i��*����r�s�Ӕ�ʪ	�xH1Ͻ�� �:6ذ��]{[������0	an�M���z�U1 ӝP�U���1OM���c�]x�s�������1���q8�1(=��t#Ar�t�P������#2$[�u��	�78�,�U~i�~C��锫A�u��y��HW!�^�f?��f\O��5LSW涒˛{,ΰi�f���7m���
�C�O�k�C��k=���m��5����t�V!X!� �!f��k1?L���]O�����+�V�n����T�z5»����-�0�ޏ7��<�m��ZC9G7�=
E#rz�<U�{�uq��W�L6�w�L���QhY�^C�,���~���ʀ>[F&�wP�&B���$:��ύmm�9�j[NT7������+K�q�#uU�}�Ĩږ�_"A�D�yQ��n�[C6<aܝm�h��&����ky�UE�7�|Ǹ!�<�t�[:d߷���1��:u@�nA��k,�Y�������mgx��[��J��46��8�J�xV����d3��^||^��B�Ni�a�my#�j�Z�b&��)�(u�_=�"��R"��|"U�EbU����6b8HH)4�=O���\�ݷ-�^���oK�m<�41�m+�K�y�8.�¬�H�Q�H��7w����YU�7
�R��]��8��{�N��\�W��;�א%��N���,�f�j�_m=�	Օ7B���NT8\�����1@˫��C���f �a��v��,E0����$-�(�:��^���?ʶ�A��}���;!��m��k���B�5%�/�c�uIO��ɕ�������y�w�E�P�����ϔ�p����/�U�	6�y}>��S��aSA�_�;��J�gi�{��w��s;�l��z�CӨmf�J�Og�x�5S��l��\�N[��7�sZ�r�r��]B)oz_H�/ݩ�]M�V m7M[@jL��ִ�Ӧ��Z�;|���`��:`gO%`�.�V����i��4�vjj/��3��xs�r�dƎ��E)�G��=)wx��̖�̆z��<9����j��lcT�=�9���k[��o��[0xȵ5�JVV�T@����&�j^�����7�ggJ)̎@Lm����m�#�#� �-�����6�f�&W�%K�Y�i
��j��a��Ӳd����cZ$򬢡�N9���%�r\�|�*�J�B�������7t�u�g`=N���BݘZ7Q����+���|��[�K��߶/W:�f����h��v6�m�{���U�P�M��##w >�nx4�b�:_��=ƚ�9��W�&]nQ h�+��`�Q�0A �~'B	:n�G9G����̥�2�ul���m�t�ǜ7R��W8lؗ���Enh��;��c2�6rʹ�I!d����T<<<+�N_n��_�*.�M�{��b/,j����p�K�8.ċo3�(�M�6ya�E���[\z��׋��-�$�9d,�Q-\��IU4%��.�\E��	���w��C�F�	���9���r�ݳ!�����9�;:[��B@xWZ�i��U�m���[w<b\��M�݅�t�U>B���yJLS�,�@C���st�V�̒F{3��S���S,��w@�C���zw�jU�C����]�M�hsܠ���l���vD9:.��I�a'��퀺���<:k�O�7�̯U��&a7����!�v�a���fСsc�{�,6 Ub��j]>U�f���M3�:�z
����}���HN�����l�׃��d�h7�d�%�������3��,���#�"7�<�u~%�Y3S�22�p����[�J��>��x�qKf<��:�:�J���lkEml��̋6�,j�7�~9ډf��NbEmξZ9��|��&���O�[Fr�ﾚ����ሟp�E{���yN�>�'!�W�񽫮�i�������f��E¥��8
����r���]5T���t�,�;���y��`�g4��J��F �䦂��b�|���ǜ�_NVNkS�cW?+DLﲼ'�D#��ރ�{=Pq�TϷ�{�P�JB8�&f�[W_f�L�{&g�c�gww�A��y�2F��m�$�J���\�2|��L������l:9P�#�*����>�rا@��ZGx�:�؁Zk��3�DS�)�i�j;��v�F�d9�U�+�[ݳ�o�0�� �i��I�w�0�A��=���`5��`�шpk���ݣr$� <7�s4����)���>�cҕ�33�B���GGWpX����NɒV���ųlIs&������H�C�O�Npo�'2W1��բ(�©������L=�4"�j@�\�н!W�\�\E6Gn��e���\�yu�C�Y��`=T��t]ot� d������^�c����M�[�����v�9�Z��Q�h����uΝf`�;�܁f�Q�*p[r�vj��;;����צ�R�>ݮT� v^�,��89t�{1�m��L�7��.�s,I2j�[���S�Jj�f��e0?zxz���������,[l%�te[⹚P��W�2��WczT�Ǡ������v����|&�Y�3�w�|�2A�x��?c�\��2���ך�<�R��71�ǹhN��7��aժ��}#r�ώdu0l~���fl�*�T����{`x���%����Z}=ݥ�"����n�Ӗ �+&�r�Ƥm8{�1��1�tu��nQ⣏-~��0e6c=���j"�v�F�&/����D?��R���ʖ#��w�>�T�L�*���Wyo�*�2}���h��|Zj!s�wu?�0��˴gZ��������7d�'�f�w- s�G�p��{{A��x�ψ�,�Ii��u���Ӎǆ���t��$Mtq���w����<4�q��O5y���Xa�Nԅ�n.)�-{Td��Ĕ�W���Bie�ۥ�i�ʦ'u�p�9}l"@�T}y�V�d������6��8�9&�{�t��e�b[�AͭDê�'/�E���ܒ��*m�*��y\>�ؿ�H];����;O+��Eu������g8ฎ�r����2q*k������zxxxxx{�oʬ����j��(*s��*|SJ�	25[���&6.`SGMgFu'Y��@xU�!�V�໺j�a29(Ay�tۼY��heRB�) U�h�w��ŋ�]��F��E�N[�9W�v�e��V��N�B*����а,P2^�O4��RS��j��绕BǦf&��T���j��Sd�N�6L���6] 2�O�Y��S�o0nS�P���-�[q5�Q=�wPL/s��^����q��V*R��8 = ���Ż��jX�Y�/�4i�s��}���1�A>�����O.��~���|OW���sJ�����(Jz�"p��9-�t�Wl��}W.γ��;1�ᩎeN�Y��u���=���v�Wݎ���F�6�|q�p��{@%>*�9��M̡��p��Col0��Bx�F�����V�]۰R!��)�ji+z�i��Fc��-�}gt�Eer����sWK�zeA���&y�W����v�ڴ��L��ˮ�;u��\朧Zr��R���gͷ�ʔ+*ջ}Y�{C�}MN�3�b����	c�ծ�D�ɅZ�!�n߁�.�w.�s����
�E[K+���Ms{N�S��o3��-˶�D��n[[]��V� BJ=&�+��a	�L�t;�ϐ��0m����h'+��u�W}��VB��ڀ��YrT�f-D>@#�'0虻m�B	f� ��gf-�S��)������أ|)���� ��iT��-D��^��C��gOsi��\0)���x'U��[ڟ^������)��4R�:��%�ou������S�d.�3���-5V��Y���gR�) 7��%j�����{)�/I�Ѕ��o'om��:����6^��]����WL�v����w.c|+Ax_dt��Zs��P�P���Tw3l��o��u�3�hc{G+j������8V�g�:���oi�{�t�C�U�g.\*^���s9@��S�rWvRyw6���gVgwF�up���S7L��ӻ��;�%1v�ۍ��X�d��w)_va�u��1���2����RU�v��&=��(�*7�ʣg*wWP��G��\'H�����lP�t`���l���
�*��LG �[6ϮJ;�݈x�Ƿ\\{�i�2��f� }nRm�B�a� �1�±W�YD�"B�J��{��c��S�h��+��'�\��u��X�WvSK&.��דqA�E�������q�1+ ܢ�+�M��Ꜹ_m�G��*:�e:Z ����k2��]#�r����
	�W%�/�[�z��IҞ��Y�ye�
8���5uwK�+k�����\ж��]�k�:g^��e#�OE�q�%r���ݹ��T.�2�)&������NmoI��c�8c��CxS���2��(B�F���I]W���׻;�58-1���j?�v�0�qnRtt�K}���	��֢wڊ[WcSa�����MuXO�]��|�7ݻ�q��	u/i'q<R�˺"��Yc��A� �Ɇہg���Wn	�S�+_M�`�@걕��t�%��&��n�+P����O�$�W��
�"qn_R+v���']ͫJ��)WH)v�೵@whZ���	렖Gv�n��T���ވU0l˕�nI؍�c�%�el%��0�{��v�7�9W)�F	��F���Y�����'�+Y���]��Ae��ʯ���3x�n�JV6�jG�2�(Nǅ�Y=��Uܫ�G��V��F�$��K�C�Y5-�{q.���tap7�ɩ�#�ݲ�Ʒ��{�wk�<ַ�~���!H
$`�' ��؍�����dH]�萑<}t�:v��8��<~�X�ӧO]�H���Ik�r�O������W9��,`�r0b��h�w^WKV�xKz����ێ8�>���ǯX�ӧO]�j�XU%B���	"�@��m)bŃ�턷8U�s!mˆ������ӷq�}q�Ǐ^�ۧN����|\�]������t����������11�M�Q��0,o������wu�ʋE�����5A^7/���� т��j�7�f�Ħ5(�Ů�@�nENr��6,L��ݴ��ط�љm�ݒ6*����65FŋA�LD�W�W��DV�k�_�űjLO���Ko�rxۖ���nkr�*r�2f�m ��
�"��ʛ*�5���YZ��^��QT?�p��2H-��hдҐ���(B� BBNDHt|�& �7��ǧ�W(.�َ�k&�j����NmsP
�]t�)ês�.��M�m� ��fq5�ݒxÒO����J6Ke%- �e1m8�AϘ_2
D��"R��Ñ��3_%TD���qdD��hBl2�!�� �J�Q�,D�	� �B�mDQ����ꛂ� ��^���g���sw���',_N���/Z���h�԰�]����z�/�Ĩ�Z䧊�A�:������w\v���D)�5�2J���ꢹD�ay+t	
��
��7i�^w�;S�=W��$�̞�;1���>�ux���TT�0;٫�$�a1ٷ�\穪r+N���@����@ˏR����`���8��L#j#��b��f�ʫ���%~�a!�O3��~	6ڸp) ����.f}��0ʄ.T�+ǒ.��{�����``I��\_u��n)Em�c �݉wʡ�
�N^I�4�l_��"�g�メ@z+��^J���w�3[�-:s�݈Ɠ�+��(�
�Z�F�i�cǴ(�9D������yg�)��Md;�;ѽ^�Bz�Tg�e����\�����K-��ͧ����¥k��m�pD�����5n	���A"�1#O�ЎS�������3RS���_>WJS�tfH�wk�X��snR��h6�NE"e�]��n0]I��;�=���D���]�Ta���1�J��M,�<ʙ���ڊ�.����݁�����b=Ru��춆7s%iX�Y��^o7�����F�͢�^�`�Q`FTz�u���n�F��) �G=0rG*�W��`��nV�۹޷���@U��B>��#E,�7r<i���ym�����YMn��
�5���c6n����õIp�z5󻮰����gy䚽�G���KF��X�PIq⽍���kD��:�҆���WR�r���UF���x����,s�p���ӵ������ә��F�B���O����t�=�#�W(�;�㏉�}4I���T����xYM0�wW���h����=\�j@�%�T��+u��k�zW5�K��C���M�luȦ��U3���CM�.S�+'�c׋�m�2<�}5���m�c˄t�'ە[!���7�Gs�@��V�1���q]w��gol����c��Z��z� �����(㼵'�k���J}�V�Y9nڢ�}��ӣX8�isM�|�>�|���k�}W��l�g�ҫv�[��h�h�X�b��d�s�n蹙d��a�QF�����Q���T@�A>]*j���������ُ���T�<<<<=TZ��w��f`������n��[L�דjA�x�@�m1�2���e,T�}o	Qi$�2�H�g���~���s�'{��|�I��{@ź�"�ϳt�a�h�DlE������ ͑�5in^��.�_:B�]�tƙ妠{l��\�W[���fq hX;O�E�'Ķ�yM����{�ˊ�x_��垻1�( i����C|i��8��_h�����l^`վ���M�|W=ig��I�	j8��Val-꠷0ļKP���r#�IR���;Ŷf�k4��ǜ/%##܉����̴�|���o�s$^��C<�]v=��:���B�k
O��Y.��c=<8�m�.�SY΂�+oe��o>�*ss]��|P�5����&6��j�*�����S�Q�׻븮{�bo*a�4ǐ�(+ G��m��ʨF&�w`�h ���7�~u��`ي&m�
�3��L�����k"�q���tȾ[.j����_|�`�ٝ�.��_S�l�Kኩ#U�$b��4E�_r/;z��R���u�9�3٧^ڭDl����\�4	:�{n����q���ﳌ�:�\棬5F�Ėn�y�o7���Jh67����-~���+ϖ��0[��w�����.�$l�i�ˋ������7�ww(�=�!^����Yxg>��!����gE�&l��vR�)�`'a(����������>b%��i��jw��6����g�+FbprR�6��A9���2I�RXѻ�̊N�8��n�'_�D�D�y���"^-,�k�>E1�J=`�ֳe��#J}�|�T3�3�_@u����X2�Z�$�W9>����6���X������>�gR�8���k��ܛY�����Lc��7}�9�{e����؟n�w��nT������ǐ�k�V!ˉ��0&���:��]w��a% �Ƒyw씽��CQ"�W����Y�[���|��3�'�[x��77�uޛ�|��8ܭ����B���E&N:�8�p^>��G����*�����4W��=��g2�7�r47\��_�v��3�!����}pR!)��k��2�m�	���*p��9+�����B<�5�6I����p%�{m�}^�1��&�L�2w��B_��M{V�wr�c��OxR��$Yٛ/�S�&`[�k���/��z ��l@ϰ�rG�������\,����]R��iAxp5,�N{H�5:G%e�wl$��si��+/[	��+tg+�=�l��G��c�\x��%#vOvu[��sk�Vw��8�akY�mu�p��>~|�����t;f(߶��� p'���ت�;�n��C;��U��Gz���s����Gݔ��Y�^Άx�˺��T����U�O�Ev _J�W�U��I��ӂf�?Q��V�1R��nq}�"O���'2�v�U1�����;M�n�u�d�k-�D8��@�rc�c�F�vV�;I���࡞UT*�G��O�T�$����~%h�^�/�1��x���P��_@�����Jy�U�i>�m�WB�H�}A�]��GsO��w���=ⅰ��,���p�)K�>O���V�w��Eچt�޷�{���qR���|+(-t�y�7>�]���Z�Jwx-T�*ǫ�O�+��J��V$9z%I�&�J=�C_I׳���(��O�=�7m>;�YLΧS�,��j�������P���|���Ԩ�~�JRe�|��*g"�qڽ�Т+��\*i��Ţg�K��Z6�z�5
��T��,z���S�%��;i
����P�L���"?}�8��hV�=�GF�׆r��;@j*��wcH�����[u���z��R�X�O->Z:0w_��z�m[�y��t��R��LZh���<2�e�*�cMLKڬ�h7W��~U����m��R���jõM��-�46���I,�OyJ�p&ߤ
�x	��U1ʳE�Y>#)�fs�_U�!FHY�^���
�F�mr��C������
�=��9��ɞh�o�Ko-�I�_'��T�.�>���˨��q��A�xoï��[l�cӛ����&���AS*�{/���Uǭ�{5�هk��&߭��F;3s�Ζ��EN���s���+Tɹ�lв�Er&x��x�};U�v�1368t��W��:�G�jU�"���Ҭebz߉�ZzҌ��-k}�k,*wV*��R��A�.��6�	��ۮ��_a�6�$��#\�7NnK���Ի;j-�[���nw�m��~��o7���qH�%.2e���5Gޯ�����#:D)��j����m��b\��8�?q��}o F�`�i@�k��n��= (+\���&�ҖU�q�K��e9����`���.��>o4�0�9?y�tsm`�E�&�=�X���؋���g�j�d2����:����G�~Za�	�.�Y��^!��+�wh34�2�H����#W�ֻC�5dI�Zk�:ym������P�Y����;�����w��� j-��-m��y�&��|r��f_��m�8E�ݥ>�/sSU�mz�|B���B�m�-sx��ee�a�d܃��|������qH���T���{�"n��b��#Yn4f����X���«�P�?�\ؓסuξu�8�ޝf6���Ź�
�6������!Z��z������-�XOI�Et)*
5<J�ں	L�%�u>�D-����E�����&���������� 9��<��İ!�Ĥޜ��);]���N�����j�g8V��b�R�j�Z�Lch�X�pW_fI5�s dՆ.�[ۛ�k�d>�*���c���N�}�=|��	��|����C�t�*��/�rߤǌ+���΍���Z�;�)OР
�(�:�:�w[����ml�"����KЎP�&b�\?����Wwuz<GCv�z���)(7+�ȁ<U�_��kbضv�}7��Gne����� �_�NDs�d��.}͔`��:#�
�w��]l�)�.3t�9���ϸ�m~p����vz�򞑽����}J�T�3c�J��%CGn�Y�����4�~���À�=칙y�����-���������w��D�X����K��J����%�3d�n�mIѹ�Ŧo1��Z7;�c QgKx��J|�2	�ܥ���ǵ;��0w�p�|�yW� ���NrD�RS��v�����m<���154&��W�����G�"z�}u�orz�6�V?����@���O�wJ�H;���fRh�s|�;��+r�u�����E��l����v�^���嬜	�+���C+36JU¨��(x�/Q z��"��DؙG�K���j���_����-��RJG�us���&�-�՜�PN�쩪��,[ы{F������V]��Wǌc�p�'u�/�����w8�p���h��b�5�J��|8��Q��Y,�(�p���~�&�лm�O�x*��'֭l�j>��Z�d�;͢�Ԙ��hw�Lx!��p����<�����廤D��p��ԧ<�%�#5�{7TΧ�L�p��]�*�g�}:4�?B�vq��:I]�)T!�۱Q/�[�s�h.%�%g/�؜���2�.xoMϟT�bۍ�>�#�_PˠG��C喈�_���63�k �}C�ZO��ӤG����آz��2gM v�^�:��30�3��h�k�M� -��r�#8��
�=�Ґo<;�����'��Gv�.�^�]>�v�>�xm��ֽ<3YQ����"�󛵒[CM��hܼ{�lt�&6����I�L�/^4�E���ap]eŻy�e'�zu�ye�A�+|�J��x�A<bE,�V�^�Q_w7��(]��u��̵�7k��?e�F�啺�):��Eu)D�Tw	��r
���d-'{�福�̳6�΢��N(x�K-���WdY��g&Wa����Z����eH���C��λ��tSy�����7�u��p��y��`<�*Q+'�x���b1H�-�Nݫ��� ^-�h�Fnh�[�֨}9q��������6��e�0��م�J���'e@�/��od[�ތ��ʶ��i����S�=I� ��y�7�NkՓZ�VNr��9$ϴ�d63p[c�{�z�Fw&i�M�&��َ�֪�G�is�=��P5�������!Fz8�>��F����U�ӷ`�F@�HN��WK^n��X��Գ�K�i�����1EM0�S?uN�7y�~Y"����"��UwR�#6���/�ͯ�q��]׷ZXK6l2��am��zeZU���]\;��a�LZ{�5ݫ�:��/���}unhPN�M50�vuG��YQ�x�X�n�MS�6�M6�9��%��fbޝ���q�uS�VW��5�[U�yc��>U�ަ;�7Jγ��n�ͮ�ȻK��4�b>���a���pi�Y��f�vv*�{����9Z	��x��e�ߛ��ň"��|D��+����.�Z<*�.n��K�QV"�2�
sr�Ӈ=V���;�\���u��c�%�Ԕh� U�^�.��&�۬l�9�6̻�f���%����r����LoM�ݷZ���m��:�O����I
�͎�,NV��^�;Y����ݚ����`6'a�ުQ����T����;Y\��$��,@�s���u�� �X���lgN��]�Ye4���:�-J�o���[3��Ջ��-1�a�Wf�@em0z�s'��:��x)���PX��SU�C��8@�#`Yv�O��/�Hw"�=}F�pR{c������Q��z�*^uc[ojn���Z�x�|.�{��X9m{[\��u �}��u.!L�C2åEC�h#�۽*�n<:3
���������������uu*�)hH�Z�p���ރ�W>9a#HP�	�o�:���]���Ir;g9
�5�2N
X��.ܥIm��k(��.�u^�H(\�C�ze��S�-4���t��[�˷sT��4�!��e:U�Y�a�j4�K|7i���s�(�v�^hrCSz�2�W���3
W�C�'D2��7t:MO��n8�Mf(6�+6XOC���M��$�	�)�Q����>@�PCO,��I���.����;���_ǪhDI�_?Xl]�f>��`��\]&J�����jUu��.��役'�Z:�T1�E-�V��aS��+9v���ͅH5H�dzT����l�_l����R��jҬ����mh"{�j=I��4�,+�U�u�%J��n;�5t}v�!�Ea7�E�/�=����Ԃ%67��ʚ*#�|&���oTvm�i�T����{�eb�=�7%%B���:�L�������t��|o�f+hl���v�
�@�-��й�m1iM5f�u3˵<Wt�7/:��b�ɐ��c��3��ֻia��5��mt��a����:�u)qGjv�i����X��!{N�!6[Zϰީ\�������V�eg�T7��#D�� >�\�_CaK�9�4��]�6zx��Iwr�r���D�cmݪA^�'��������
���.=Tr7;E����[U��ٜmY���T�G��Z�y��r��E�rjY,��sV)O��H�+ֶL��d!>�T+��J���sG���N71�]ƍo(7Ub�YL�/��*�ܾoٖ��h�-�.���b��:Y��W|�m�,]e`���:�$��L�d��v[+z�2þ{����*^vk���8���}ܶu�ӖJ]�ן=��-�ߝ�$�E��U��m�^�F�Qb�U��~��:v��8�<x�z�N�=w�B[��#⹱��F����� �#"Ȱ�z���t���q�<x���M:t�뭡"H�I���*�6�75%B!"���H�u�ׯ��n8�8�Ǐ=z�N�=vn$���HoϮ�ǕKw��d�!�.T[r�Z���y`���4oV�Tksr�%F�QsWF�.j�b��&(���U�M&�T�W5�Qb�Ŏj�1��KA^�j����_��bf׭w�m�yۛo�wTj�I\���r�5����c`�k��i�W�k�X;�?4�4��W1����\���L���E#E$�o9U���.��9̨-��Ɇ�/�����-<�w�Wcu�2�;]�?6p��&O�[�Z	s=��9-�c�o7��� M���P�U�7�f$�x'�]]@.o.��=�[o'6��eˏ9|�f�M�B	�yg�I�ݬx���R���)lǁ������O��v�0�j
�F��&;��%�����Xn^=��lgK�=��������5��/��7���[ў��+���9�:���9��=wgR'}�[+���{ɽɹs�a�g����oUV�'��23Jm�/�2�pNH�g�#����yrs�*緢��+Z�2�D��l�{�����D�B������� ��E�r%�I��F߮r�����8#M+8yqLW��*X�a�<d2��p�ӻ"�I�i�����s������9k*9.�0c��zA�ZZ<RA�rF����Lg%"���U��{���tkv7?5ʅ��/���wp<�s]u<k�j��tq7ۯ*BU�x��ʈ1Y"�=���6�d���!�5��Pĵ�ڶ�^ä�
� �3�ׯo�w�-��u��lN���i�FU�ɻ�N�B34;BS�JݲZ�w��&��x{��N{��1���Y�w�t�}�=��zs���b���<�L�r[B�=�|�i��͑ǜ���7��$@�g�kӰ�cʆ�US����S��&BE����0�E�n��+AO�vSy#m�� ��7w��;C�Cz�qq3����'"Rq���0�U�.�aoJ���{�ktm��nSV����W�-��38�1�ܸ�*�9���?}�Y+��Feq��ؓR���p�m��1(�q�t���s	�qU0.N7����%������c��%�����4v�ʾ�^�E�z�oO)�U��yP%�!��2�P�;+���g�M/�q��F��Hp��*c���7��s5�ih.3e���L�.{�a8���(0�b��v�w3Pr�`�MȌ�w���L5��p�Ҵ���·�W~��4�m!���U:P{u��_SC0��%@XK��Ȳ�w�KԱ�{�L3`����w`3O���vs�5;[J�9�6�Қ*�j3�+A��U�4}�� {0�duЕ�I�Gx�7����/$|�j
�{�՜�ʐ���R��b�O�<ܸՆ���U���e~��=���fU�c+>��nq��\y�,I{!g6�I]<�s2m�I����m�A��Q5ו�ƙ7��j�QQ ��-VE�W���UC��q�=����->�|�N��n�Ш7wj�6)0[:�>Y�@�:�P��h1������8�؜7DV���|����o k�������gnXw��|�y��mp/r��IQZ/��SZ�����9�-��ɖ	>///�	h��ݷ*u�9x�Y9Y.���o ��I�d%(N�鼾��6=`�!�]9�:7����v1�ɬP�1�Nf!eJč���Wޭ���Tcʮ�F��sI�������:�H��uQ��W������]��p�+b\�%�j��v#b"C�����Ck�7l��}]������Gq�{��t�w�ꪾ��6�nNF�v�D�8�f��tg����%�ץNZE^l�����5�y�SC$k>��f@Vu���;S�E���b����Q�����.<����nf�t���Ы��Cv/> ��&���(9�iq%!��%�cy���� �S\�_T/s�PμD���J��\ԗ���0��o0��s��.�|S�+�9�����p�[��uK�\x�ݦ�S[�%���i.��WQy��; 푞N�|8�ThCS�V���t��Z�m:c3;�wi2���4�gp�1���(�{u��e��wKsD�<�����F�r�{w7�E�b�)q}7���m�-��|�W��X�2�M@W�/�M��Dt>�GW�\�<�I���F��i������z�����~�����R`��Q��V�fk�de�V��C��QqYS�UT���]N=̓��Y����'wJ�Q7�#z6��[{e~��-�N��2h3��C�� O�pn�X�5_כ�?ǌm��.���� �I
�ؕ�Հk��h��/��]O��aM��:�X�3~ޗ�@uz�MOFg�j,nU�S��V-k���-pB�n�T��ͥ��_���L��#��s1�&K_�tĬHJ:�s��G��&�0wcx�����s��>ϙ���._@2�|F�RuoYO9w#V�6��I;1[��+����ʲ�'�����sw���1��/��>��v�C�aQJ�(����c[�V���eŮR+G����w/�SF�1���r��S�����u��MꝴdV8���Û���S�Dȩұ�S(���	,�ӑQ.�CP(A��_M(W{����X+-v�L h�=��er���v��[��n
y�Lr�����
{�owt�r�BJ�5��k�T�����.�u��@���s6]�r�ʮ�!#��x��_v;���U�yR-'�4Y�5۽�~P�o�g>��J��`��^���d�<zۯ���|}7����mZ��+2�����O�넂������靹�lв��3UΫ{f����PƾD���KDnYo�p�[������Z�'$�!�Q&.w�'��t�)]
�6Y�|���g���>���tX�,^����j��2��U��E��hL����/�Սs<���u��R5��͹A��K��e��+/���}t��q=�.���n��(J��Xg d�}Z풤6哌�QY��鲯����qg֘�N�o��]5ݍ�9_�g����x��f�Ue{W�:�ڵmMW�i��M�7��#�G�h��R�Υ��Ons����Z�����Gd$�r�<���`�jJ�w7�|9�
d�p��S�z���/����0��X�'8$�e�!��R�`��ja�f����J|�\�ώe���29N�ت�����8�͕���{nK��s�
M�j�"&�j�W#�v¦w2�˧��tvb̝�=`}1�&����r�"���2�0�Rj*��H^V��6|b1��ՙ���{�\�U~|
.*%Ԍ1��P9iu	���d��3��	��J=[���?�4uV�o���͞���jӔ{�*��B%���X׌�;�>�B��Y�Lwp��i��^T�Sc�-�+����N;I���`���{���g3u�G���|���|lk��P�:�.�d�n�|��}���&�ݢ�M�wX&(V�y��RNt!(;��"�Kp�6��PR�o[0��V�|��m	����b����]��I�j��Wl�uu�@�o����q�`�����T��P��}��,�{��Қg!��������{���c��]���e�U��˖�&9�L�k���j�}u�N��qU���bU9��s2�a��R:�CT��<:�^�=�O�zw�&H�����4��u�U��I�����['�P������>�0)GR��m����7j-*������Wv��K��>�d ��\���L���Xs<����O��} �Yv�,�Iv�	N�v���w�j��.5�\4�o�j	|�י��x��D��L.�\�d��Q5�<�#'k]ᙻ��v�SZ��/ef��Z9�r��pj������5@$蓦��5�-5�wEʩ�Wp��xi�ӗ���kd%h
�D�~�1c��Lc��X�����c�J���vy��#�����)�o�Y��Wk�Ϯ�jo�)�Nn���d�yk�B�
��/ϻX�дWN�YuUy��Fw�/��Mnč��zHën=���-�a��(vx�f��q�&&rz�_.���vw����|(n��, ����,��鑟�vM}t>�k�0F���������t �nƃL'*����yq�{�/��=�W%1$���/�����<��W]�(-��\������xy�o7��ଝ�UQ��Պ�#���+�h���X�i���.�.�'�d�Y�t��"�%������Ο�gWu�����dY�)�2Ͳ5[��p��-
�~�^uG\�#��]�ϼQ��Y��56hS
�g����d�̠m�i���W�ez9�l@�iN�
 0��w(��F�Ps{����it�⸹���*�?(���ݱ��&�+"���x�PnR��˨'��g�r�|C�p��8r��6�����Qa�5GvͿD�O��\p�O�iy�gu������u�Ű�_!Y��:@�.N�YT	�W���U���	}|t����p���ek<z���b3���0�'��K�QO,D����Ym�L�U�iT�/(Y��:x�Xx��%�+</��^��9=YQ��W��s)O���B��ӿhզɶһIν|ڬ뻱��p�wOzB��8!0�����0]�����P�KA�E��� ���w�rW���"�&ً;b��HN�-G��&�:Θ���ѳs7�F��k�(սTSv����{3�@>�>C®�]����9D��ʁ�#5��q��R u�n\�)����8��ݟwb��x��X��A���"��;p&�|��y��]����[cӊ_�n�50ۮ�n���!^��e6�C:v���qTӶw�6����?wK�%W5&+1�j-�֣k=]�$�;ֽֽ�O,�i���������N_�w�!��t��wuK�;C����ܞڼ�rvX��8��i��֌�������O�`�rMF,�/L�}8����
�u#o�î��p�J��M@�ET#;_Z�c���b�PN0��P]k�a$��ۖ��>�.�篿9WH�4Z�u��HUT�/\F`�cXOq�����n�z9�%�>\��l7�ۧ� nm[���Vs�e��:N��ݦpkӓ�U�ar�/kʔ�J�=��}um��\XHj�z��;������*�]��(@D�t$��]A�c���\W��{ ��� ���Â-'��Ui�,[�a]ktt��N+�]l6k9��Yv]Ot�(l}}3or��F������s��y��/|�����c��׽�h%l�������\�m�����'����8;u�cM���qU�VF��j1H-�\Ldv���Dq��O���/t�elD�eBx��lQd�$1	.��2��Ḯ���������a�:f;���Z�d>�"���R9�U��Jԑ�J�7�*�nx<�w�p��}ٱ�3=Fi����x周+���s�M:�''i�7�䖪�}�D�ҽ�Rtm�?o8Y*���k��UvJ0�@-��������J�}��R$��4�+�3�/�YI��H�f��$��S�x�U=�*�6�����!/��<�<�*����'j�Ix�hQ�CwE��X�U��O���Dp�>�O7��G-O;�ZDXn�:��s�H�6����4�R۴�ӽ�Zל�>��~���uR?r� �V��������T��ae�A��tn�
A��h[5+l������X�m�2�,em�L�i�f֚��mf����,f����L�j��-i�����2�2ڦK5���V��[R�j�Sj��m��jjmic6����Z��[Rɚ��U,fښ����L�-��m���ԵM��MKjjZ���1f�5*�R�55��֦�ڛY�MMZjkSSZ����֦�5k�5���MJ���jjm���MJ�ԭMJ�j[SSZ��jj[Sk5i�Z���ԭ���56��֦��5+i��M��MMZjU��Zj[SSZ�����MKjjV��kSRښ�i��MMjjV��ښ�b!�P7�����B
Ě��ڦ��5-SR�4AB!�P"�U�D�"P������-EZ�KSkU-M��jU� �E �P��$ժ��ڪZ��RԫU-MmT�*�KR��Z� B �]�!b�B �-KZ�jkj��[U-MZ�jkj��mU-MZ�jj�]�W-M��V,�UKR�T�5�RԶ���mT�+j������Z�E ���� 2T�֖��-KZZ��Ԕ"P�D!
�Z"Vjj�SkK3-���LY���Zd������Z�jj�R����b�VX�m1f���ZjV�R��"T�J��Z�*� �d͵,�Ͷ�3mf�Vb�j�3mLY�����}}�����D	H�I!����������ڏ�!�c�V��G�?��+?h|����Q���~iT�_��>��ϓ�*�
�����?����"���ADW���?�| 1G�O�������(x� ���C��N�H��=�I�~����"s�+�����I�G��V���V�Ԧ�*�jZ�T��5��6��5*�֖Զ���mM���iV���M��M��k-���-i��*�ZZ�6��֢�6�mL�KKT�TԶ��I��V�ej��dEFAIDd@dU?$���Q@d �-Tm�Qj�Q����T�ֵ)����U�֤�h֣Z��ԥ�R�5-��iKT�jf�%�)����Y[K5�i�J�ZZkSR��kSJ��*�Y�J��Z[S*�٭M�V���-��fڕ�Z $5g�J����Ͻ?�U�QQ$�R@@I����������@������=��_Ђ������=���?��3�	��H~ ��h�\M�� p>�?j~_p���>P� �@_����=?�3�N(�"���7ъ� �����O��<�((?�
�i<>��Q���x* *ϱ���>�?���� ����=��������O�<����D�_���*�
��f����T U� ka��z��D�W��ZY�(8�ʃ����8��'��B���rF1���R�?�x����z�~&u~Ȉ�/�Z٠DQ���g֟��AH~	���
�2��?���$&������9�>���=�*D�%F�mU�"@QH-����UJ66�j�Uk*TJ�U��Jm���i�UJT*��
DT����5����f6�[4M5�e�ChQ��fQ���ܭL�VZkm&��6�c-�Z֤mR��5VJ�)m�[M���kTͦm�����j-�mRY6�-2��e\�wT�ر$ٴC1��K4�f��ځ�Zl�,̡�J
-�)bĥf�+Y��Y��hU�JC&��%�PZY��j�,�1aZ[0ͪ��ukk&�  r�z��Ԫۺ5ur�w<��lm�a�m��s�9gw���WhW\�u6�m���Wkm�ե�)Z��\�ѷu�]�ug��f�n[�u4V��u��5�[�l���Sk,mU�@��|  �*���klP֔7>����t>��֔�CJ�|���*�ZQ!��#�z�W�[׽�+�0ʶ��h�:wF�uJ�f���`��W��m[�ۻeSMի1ӚVYu�Us�[T�i�-�F�fڰ�m�  t<�Cj��vBܮ�ڛ\���mvڶ��wNچ��ۧ[mv����:�s�]�G�*w[A��]nuu)Ҷ�hm֫W;�J)�aЪ�k��͵�LT��,�QQ�  ��ʨv��4u�gs\�C;�u[@���kB���Fͧ]m��C��M�`hЩ�knˣ�(�s�ݍm�DmAY�j����ɰV�  ��G�f��[��::�:��)��'}u�	I�m��V4V�[��í�ѪQܻ\6�h֦���Gn�uj�S�]����Kj�ikdm����l�   Z��֨���랽\*��m�rt����̵E-`*j�Et7kn�Fh\�P��;�+�Tm��yf�gJ��*ɵB��l���  �� �{Ԫ{jHn�N=E.������

��vM��$��{sG�^�+�㼐(��w��R)E	ܧt�Q5��zZ�ٛ6cV��ٴjX��X|   ��Uv��v����(Sz�y�
E=��(�׽�J�7^���������T�*)���Uj;�0IH��l��I�J�l�kc[Z͐bZ��Ko�  }�jHR�����U
��wy���!Wq���US����v�W�<�� U�N�]�U ]�m���z(9�PN��n{O]B4=��k,ś3lU�mb�,٧�  }� }d�Ǉ*����)J+�zp<�A����*{޶q�J(����<tT�.�x*T�Z{�g�I�����zRT)��S�h2��F�di�M���%P�C#M E=�)J�  ��%*S&@ ��	�R��@h�0Iꔈ�*�4  f���?����?����.����s����o*G%��aب*g*ً��@IǅR�_U}�}_W�}������z�����֪�m۫kZ�ݫkZ��Vֵ�mj��������+��VҼ�o%���$����X��p
o.f(!97M�i[Orf�$Ee��bI8��r�f	�G�����7M����j��Q͡�1�W%uns,�YWN$���2�,-ǔqȎD0����Qɖ)Ӆ�&�m�j����lQu�cP&v�tn�`g(��/즨����[�����.i3���@|5�`���*X�u�L�����y��q(*&�i%�6��J�mZ`�ʕF�M��"]�
D�+�(�jhܹmɴ#�a�����������)��pf�\���e�mnAEZ˔�86�V �:��(}$Z�����U��^;@��W®�������6��YR�M� ���
�ǆ�:F�/@�8�Fn�m��&�q��"b�8�%�v�fmf�tB�.	
&�j��q�kE�ɹ�̺��t���t�i�ʘ�+U��!�5伥Kr��O&!��)�φ��2�c���:�щ�����n䵎[�8�7lr+��ä�A���*�Yъ\���C/fڨ�D��m��w�f�����*2v�vZ��	�YOq��w���t���R�H�k7l�9R�I��@�،B���@
a�Z%/u�m�؟�ƩnԬ��/^�Ƞ�a#z�KZ48��Neb�P7%eCm�ӷ�En�!%`J����i:(�1X �r<.D��5��eb�pB�	4�d&���e�Y���u%�ڷB5zB����.�K�n֝�'�c�5d���i�2�;���P��2����D6E�i�.�J�`�,�W.^:±����G�~C5#+Y���(K��
��2nde(�Ɋ��4���m�d�X]�[y�jP[<q-j�"N 둥i�vF�a�H:ۮ�}�z���ڵb
Q��셟(��4�BA���庒nT����KƖ��+hE�ۣ�I�R����U^�1�/@@��yu.%�;JХ��@�vYK���l6�®B��#-[)�b�D��j���$k3c_L4(nE���rД��M�����}�f��e�6�[���v*��)�;���y�o�Arʃtt튻�Y�4���/lX��ju���lf�J�Vŕ�,۴1���EX�r�[J���f����Y�Ill���n��E왖C���XyLn�X��l(�S.�F%E��kƑZ���D���˫��a�j�f�j�6�GLZ���Tv��U����5*8�n1n�Uʌ�k3"�xs5�0��h���*���F��6�w�5��m�� +�R���2�ZU��gZ����Y��沚�5m�72DI��q��I���ͫp��eY�V�E7I�eZ�B�4��@�+�MG�YL��Q����69T��/-��&���k%@1Y&���%���llr�,tɶ�F��Mn�Q�h{i,��iF�-�7�em���n�[`mZv\mj}���^�oM;ӊ�O`@�{c=Ǐ�1��*Z�vQ%#����0����-�Jy��b,�@S�`�f;������u�4,d�]c?[�z�hјZ2V�ŵ��o�c6���ǶB�v Q�j�w��w�P���1��W��
��b-7���jQ'f�Wu�d���&��lV�((�Tu��T�e���+jl����Q[m-��Gy�^���Uը�)���ۛ�d1 jl��f��e�Kq$9.����J�,(f*̨^3#f:)<&����2�5c~ݔ���]Q��Z�N�A���n��tMH�^^��R�0;Z��^����HT��{��E�t�fh(Rhٵ�nTf[��d��wL�g�`iyQ�N�KP�͏2
[�u���![��e<9v7 �r �;p,�A}p�+6)S�ٮ��hP�L�5���P��BC�C���N+�����PVn��;w�љf�A�e���̙�d��1�u�X�G� O���՜�X*DEhY9�A�P��E�W�K�
�G:�`c`d�h�w�60��pc26�kL�]�w7N0&c��A��b,l��,�%͡�v.Ԓ�آq��c�g0'!�jP�Cf6uT�DU�U+�s�$<����{�2�E)
i�̩"kR6�љJf��WWyUgR���D�H�2\Ѫ�H���z�:5�I��ځ-������L��JT�ր�H�^"a�Yu����gpܼ�0-]Ɋƨ�u���oj����� �鸯���� X3�����#�051���&�viT�¹�<��n���ѧ8_j�Kw�h6$Ɔ�S$rP��Ѧ�/T&�8��z�MI�U��A�h6�
�C���ʽf��2��8��Q.���q�G_;�Y�`�����NUԖ���jUzɬ^��W�,ĩ ���6��Z`�1^�d�8V�j\�(���WGm��ݔ��%�t �� �Də{��u536r��#ә�hȬ��Ѡ��EI]�Y��-��v-AZ��.�l��>s[�s[Z]۱oh��x�je�cS!G�ѓZx�i3[@5775���&��e
��t&Ne2!\����X�V&���n��@Jp&�����^ժާ��0H�1�P�y�TN�ګ����*ù����R�kV*���|�q��j�M�kn����dVf,����u�M�r[zN����ƨ^ASAc%��`!v�<�+M:�����o����c?!v���i˷��XMa{R h���#�kr!6)����X�E]�
��i#�Z�E[�Ζ�5��T�˰Q���Z*z*Oh˗�^d��1��C.�oeēcH���E+oҢ�j�6��p�G%=����8-ѹ���
1�-cz�hw�2̰�"Z�+.�640] ��mnK�e�z��QKP��!&G�jW��i��E!W�`���Z��k����X������6�onK�BT����u(@:f��r�����s"4���阎� -VP�����4�;�K�L�^Y�mH�ȉ:1m���v&�h�KqeU# ڕw���8*HbT�6�ۣt�Y�pۭ����6ТF�1w�!���QׯoF���VI�}��VfL����������'6�l�A�[�*l!3LT�����j4 ��ۄ��&�h��Tv�Q�2����n��R�䖰��F���T%�Xd-�J�f�_��Y-���!����7l��.	�^̑l��0��2\j��/q���[('c0!b(�V6]����p+�xf:���(X��J
5�dZ�
��0�	�p��3T�E�wu
ͬ_1�t�P����r��a��f��I�v�q ����-��jR�52�L��t9��f���SA�Aj�sY�غv x���u(팊tdA���>D��NTn�Ƅh,���+�S[��a��So�%��(3G7%{�
[�fȪh6��kV��m=y�f;p�M�g�� l��+EM�W%[D%t�)�����ۦ1�X頳h� �"j��)��fIW��fk\n�#�8�C%b���jy��l�K�ѬEVQ��4h�H�Vh���b��w��%4�si�F���6o� ��XSq�)!.�4�7k
���M�Z� 5����3W�i`�$��Y��/�Y��O
����*X��yDp���q�e����(����F�:p��I�P^��j�X��q5eJQ��r�جA�Ua����W��Ej��Z��-m��«q'�e��iٰ���V�w�LCKB�'pb(�{�F#1�Z�с�ʽ��H���Z�Q�5j���z1��oY�JI���-a�����l
%ޕOYr��\�=`SYX�㰣��H����}\6��`Z�V����Kq)M�U
љe��)L��kq�#�v-S�b�%,K9�mT۬��p�`���ZM*ݱ�M�Ʋ"�!�%��X��)�r�{�#%��M��[�֟�Iy`�Z��Wh
*�Òͱ�[Z�I�����0&�WQ|����\c�CBn��f�
[�,�"fڛ2l�.ė�Ĭ��L"$�d��vM�H��ʻL�{��m�k5�^��.�=Ŋ7WRҊ�Vt��dzѽ{J|�ɂV��ʹz���/�!w��E�3�{iLX�`֧`��0�4f�VN#N���M�W�G�SG.�H�㥦�Yf6ыtZz����,�:�Yt�$�Iݔt3L�cq���@l'q�60D-����<1�jk�"i\�J����D�wt/�Y6΍ۼ�X�HQ����Z-ÿ32����fM���4�t>Ci.{e�p<�W%�q�cn�N��4�4�d�|�vd	ԫ!�w�����y���`�0h�<�I�E�)�Q�V:�R����Kn�i!�� y[tr�`�Q�dTf)w�t��
VT��/p<�X��D@E�j�ґV��~�)�j���O�4��6h���f7X�ҹX*=�e��/,����8������Ff���qGPԙSn��[�X�ȍ��5� "ʕ�Msw3U-�QnQ���XeB��<�a`���"r�=W03 �Q���K`�dn���lK;5̤��"�X�����%�ז��тӬ�EL�43�q�HaWp�� �t��}�9K��%k�b������Ejڴ.l��Qɭ��A��B6l��h0ǔ��B�co [V�]�>
�b?�=��0&��&����:vи�nMn�`E�oM6�2^L�M1)-rfK����3Nܣ�LRId��k5uj`w�,3h�2fT[y�f0�k��&�r�V�AX3�y�+p�4�:�T�%���2�l;��ck)�.��r�I��ee�Rh6��'n��UGqD5�(��vT bt��jG��/[-����6!ef&&YǲE6��,|��b +-�[hƍ��wN��n��X�t�:0-j�KSlѣfF��+���\�`�[��d��L�1��[�Tǒ�;8�ߓFf�CI�I��քU�p��%��L�-ѷ����j]к��h�f��KR+^�N!�Ӆ���ʹ4��Ӓ,���n�����̂�'^���4k�� �͑C�Am�r`�X]С���4Z�v�����>Ϝv����֩$un�B�[B���P6�'�Ԉ�Z٫(� ܤFZ�yP����dF�ۅ��P.L&$,c4��)SX�%]� �d8j��ܽ��3h����[�"���v�$�ZZ�*�V�J��Z԰�ʰfnPA��Q�WA�zYAa[
�$<����vS/*[�v�6:�k?S˖�w�u��c%/������
1��r��gc�Z~�
�wx]ر*liVؤ�1C%g	j�9[�LV����{Vh��H25��B3XX�f�����їpkXs(��3�*!z5�V�����5��ԓ�I̘t,"}Z������:�񔌫�e�{(��LmG��'¬&�hie�Q��Q�w6�~����ӗ��4�ުfLu75��a��1iRh�B�	����*MT�t(U̫f�9��YOJ��+��(	lf�o*����Mf����h������\Շu�e�v��DŪan�!PXM�kl�5P�T�5͠�X!�.7Mf�x!xe��E6�ц���"�^h�t�n�c7�X�E�f�p�61sM`3oS4ڛcPD�*V���3�p�7��J�j)X�#"т��d�[� �x�4^d��Z���wq�$��t�_ &D6�Љ�DAJ��+�u��J�u�"ƬA�KV�d)B�S�T�ޒ�EC*f��t6�֭�`nh���T�t��}J�P9�Pl�F��Wg2�zUa3L�X�SMc:���{��8-��U�Vf���a�oqV�[pAy)��ªTs!fS���$���ubzU�*�0Ѱ��p���$��mca�_]���&�a�(�.�;�^���"+��Ԯ��4h����%F��4���r`R_�Em�^^�TM5S�����dj��#t0�9��f�c�7�/[���mPG��Gi0��6��4�����z����ol0wO�줒��{Yɶ�))E$�4mֽTl3]h��:`ˬ����ي���H,�*"%-ٍD�I¦�;p��F9ai�4�nXB	�›��4�öҽ���f{ P�+6l���i')�Ռ EE�هN��'D���PeM��-1�L�Y�GW�*�i:C�t�j��ڋ
�!�;P��KUu+4�[����t�Tݫ��B�K�hѥwX���pnC�j����v�I3�[lm���\oQ�隡)d�j��R��كp�'�����'M��m�t6	�H��G&�KۛcB�S�]�Pe��ck��x��伢��<R���L!�4�3p�#.ث�[�.֣{2<LK�e)����#񐣅��Q��~�P���>cE�Ɔ���T���nQ,D�:řlZ���SQ��ymXn(*Ӂ`Q�omh(d�{��]"pU����T�j�hf6�&}��#hhZ��fʔH�5Ѕ��Xh뼍�x	�+py�q>�ߘt���i03P�Qޜ�9$�&�\�a��:͌9	wSF���f옄�\?K-� ��J�闻t��9��	m��bd��[l�( 7�(�Eڥ[Lݨ���[p:+#{�E�
Ɏ��"�K���eCt��@��nc�#G�"e;N^����ҨԨ����u�!Aۀۥ�lK�[|���Y�W4)�*��)��9��U����ڠ ]�R�*8��0[��$�.���,�i:Ҧ	Y��pIj<ɳ
M<�y4=����f�2�r�P��;�e$���ӥRH�8Յq��M���!��B釕�$v�%�������@���z�9'N�n��[9�㝳�G��=q�7x���ow�\�gun�����w)|M������Å��bOS��Bc�����QZ($�ce��Y�roY��|���lz�1Q���s ��i��xV���a4J���u%��Ծ�q �*!��ЬZe���ouΊ���/�E+�o��H�]�G�nWe�ԕ���-żx�33x���r�4��;�ȕ�@�������9@$1N�[0Y4
[ZHe���ٺ7�֚.Y�#]�N-�����m;|��M�h���7R V����:�NE9�[ܯ���#!��[��{��{��hL�;��"�y׍\�]�k�B�ڹ����o�KϢÈ���նPl�;�K�a�Hw����wl�����DK��h��mm� w�s6h�v$�Ņ�o��<�ajH�Cr�tN�L��u�w���`�5��2���Hv>�99VpRfֳ����f�t%�nt��h)�6�ya��G(�,�u��?��u�C:��0z9YY��g+�{�F�revϔ8�[�<F�g#Rb�s�Y����>iQ��R
DR��Y"g	Ֆ6W��S(��5���f�7�!�:�|��D���L�Q�nj��u��AY6}��o�n:�Ma�/������|�NlS��X��sT�td�S^M�f�bt6H+��^
>�q�{��ޮ*�e��ܱ��6��(�.��{�������P��y\�I�x��KM��̭�-�����:bޠ�
�����Pv��SD�ij�6lUoHA٧o�c�SnW6�c����ɭ�7�a�+�����rL��rI�]N	/k����V��錁e n���F'5|3ll6,�C���B#������z˵����y��[+�vq�K\A���vt�Ym�V�S]���I\��.6t���*��qv�qQ�qߕy{@6N5�Qz7.K�[��� �f��u	d�pk8P��t�C.�M�E蠬�<�{�X尜kRm3č;�p�rt/�3;�4�Pd?$`��\yK��jh��䡜��-AtS��۔8�E�|��o��H��i50Ic4wh��j^�T��n]fV^վ.p�G�]F�Y��[�e!�m?��GO|�AO��tUmQ�=KZV�^��(��1*kWN��f�&�"��b��;Z�q�4<�!��;8�n-�[N�T�k�3�q��¡���d�3�]xxQ=9���Os4�ۖ`l�q�:���Ǒ��;}��tM!9d:��j_u��maR�S�a��ڻvq�%3�+'w/�����~Ɣyw\qRoH)`;�D�̩�b��Q����>���j���7�_(�".�)�{O��ppͶ��ckv��i'vrCl�Zc�E�J������h�ŖU�ѕ��MW��E_><t?�k9�+�M��:c�dS�Iv��%�ݾ�L�HvgE�^�6�VH�[(�[M)�R"��0:q��
Lb������b�5s�C:]Z�fL���x���k�^Qw�n�Invsʜ�b%�����lK��TyX��!�2{t]�y��UV:�g����F�Q���F��<W�b�թ�bG�W]e�ǔ�k
�9b���X���ZhwH^C�&��N�2޸�Q���]lg��D�0L�������؝���1$�ū������2���;A"�삱�n�bw��qe�� �uQ�*�ݤo,�0��&��.����Zܸƶ��4i���R��#WʜX�#jo(����g ��n:QK	G������]/��0��˥�S�k41�ta�3��$�z���kxd�{)��Z�e��T�w��}��;^��z��E Ť���Üq�7&<'$���).6r��v��J6��,4'Y��;�Ug�*���]��L�n1֨�s�Je<�}8;��uOua>T�]K*��Pm��h)U��2J�Rɜ�ſ�S�X���q��.�<�Ѣ�v�l����:�I�+1�LX��J�;�pn�N��#�6�-�%m���e5[R^�]�K��]uYm��7%�J%ɷ�ՅW�8��A��/� ǷN��F���@�����T��]��#a��^e�Å��Tn���:�jDY��Q4Nז�k��h=Si7v5��+�a.��l^F�����+
�W"��K�T�o&�ۺ;m\+�K(�q;�Ԙ{x���I��n����=�%�R�^�����k:�Cj+�qvgV���em���f$��+�@b+k�'L�-ŻC��n������ �+��kz	-?�-k�_b� UJ�;F��ee"�	�&�u���kl����n��O$���ϜK��ӊ3s�t�q�O1�$L��w�>��k3�A��Z��;�#r�+��h`��a�y��=2ma��PB���(ٱ�������(3|@�pW@�<76�>��K���Fq7)�:b`�KF��hPϚ�R3Gp
+�6��2A�JRmĲEp+�Ga-nX�����u��y�|�[M��)V^�b�w��YCh�j�Z�Z�a^O�Q����Ih�hF�7wۙ�u$>U^{U��-�����	�����#�K�mR�N�]Y�j��_�4d���d+]�mu}��]X�T���\�5s3�*�ùтC�*Mg���y�t���V޽�N�[����RR��[}u��6�6��7o�g&���|��t�f�D9i�R�5�%��W����[EGP��*vQ�z�{K���'��e�o!�+_��,9�����c?vsWGwgLy��0�F.�6ҳ��<����(��s{E�|n�Z��:��32-��`�8xa20�OJv���i� G��
�N^^H�%<���@�C,�)�]Gn�^=p��;Gd���,���fVX�
�W��2��]}abӎt�R���@=�1�3�uÂc�ݴ7�O	f��kh�q7�#�RR�Y[9�wN�f=�²�]�k�EA��*[����/pJܭ������(��WODB��EY�y`��w{�B����J��|���s�7�h����r^>���;�PU�I]��O��:u'�X�a��)�M�ٷ-�R�4T��N�FU�cj]������a��|�s\�b�nm�h��Xסu��)��� �`��Sb�zRC%�[��	�p��ӭ��'���[��y��Oo��qN �ǚ�:o��9����a�Nm��y&����v77��8�e?��71f�]1:R��ju�Wn"t]X����d$#�̬��1�t��`,�����P�0r-�!��3/d��x+�7�Vx��,�Ԣ��GU��cVB͠t�"^J�I)K9����[��a�[p�T��m㻔N��2����-�3E!�(�x�V�t��0MeT���+yt��u�U��)��3�MB���gG4LI ���1���
��9@�Wl9�/�<����yu.�Y�HoQ�� N����&�u|V6^���ѭ6���+���o�(�oV�ֻm(��Eh��㪯zd�t�h�d7IQ[�so �E\Ϝ|�$V�\	����A��ͷ�+,�i���FdU���
a��(�٤����zũ��"�m?!��YqJv��K�Kk����;�"���a��k�b���fc�^5&W�K.!A���9Qh�8Z���ٗ&|/^mj�)�F���M)��^�M�b���=�1w'�A��8�̛WYaV5�窹�+�Y]��C ��(��UYI�f��S�G��硕���]��*��$r	��Z�}����]�G� ������8'��ͭƣ�ov=���._!���~���$�ձEx�D6��f۔g%����ާN��:1�и�c5z��S{v%a�n�I5�ơ�Ve��Vk���vӮ*�X�è��r]vU�앨��T�]3{K�AC[tҷf��/���jFZ��Q��ѵfewW,����a�	��$AF���iu����P���MV�7���ԁ���Z齁[�I�i=G	$]_hF��g�f���F�9��09Z�]Z��1���N�в5�}��S-K/A�a�P�#��3��ԭ��%f=!օ#��df�����^d]4�Φ����1J��$WX_ŲěG%��hc��0ށ� ѓ�qS�{�;ݔ˟��t%Jm�D(�N#���׹y[d�NY�_8��dzu�r��00�᫞�ǲ����Vq��tz;��9�_c��!����ΒUܛ�M���KX�V��NI_U��=v5�&k$Vs�A@��ۊ:�ٜ��+���:��gbikg���۩�q�ս�Ka<kH�n��w�Rrn�{w��ރ�i�䁮k�wg�rK4�BCˢ��M^��s��A�5z�(fJ#�(�E�B��SQ@R"|���8��7�����d(s�Ѿ�m�9��z�蝀�E1���"���71�e�r�G�c�D��$h9��:�(0�����>[k���9��L<i���Z��)�N��D��wlƉ�\�f���q�Y�����kQ�i��{v��Ԅ?�QpF�>Xց�<�mM(����%Vb�f�3��\Ȼ.d�dH@ۘ���w�j�p�}��&�f2V�����Dj�-���W@����F.�Td�!Q\�x]����R�R{f�U�9Y��q��:9j�ѭy*�6����,�\<�]>S�쏒�]Y�Sɦ� �}�(�f�'U��z���u�7x����Ja���f��$w�gE;P�u����K�\�(��@���Y��ӫ,��,�R� �h<Je-��嵽:�|K�T��]ҡS2�Y5�����آ�#���y���l���!lr)Hݼ��ޱ���KyM �u:���Y:S�NC�oeH�r�\�nљ.���{��/�Sѽv�l��r�Q'�l-�ujv]g3mX���1��)��7��[���)w�!Ͳ�K2���)]�v15KISQ�	Z�{]�^�C�v���,��#�}.;�M]���d|��<�b���;��%k���˜Շ���i!���m8BWt怹��/��U�w�.�=�������dv�V{*ڬ�>m�v,m��|� �!�*,8�)n�tFW<��\8�CD���̫��/;���P�����X� tװ_o�p,��S�g�;��s���b�=���S��zbv����=�6��7��M��T߆Ħ]/��Ô�o�,ʜ��<�яu*}9;v�)f9}KkF�%�\8�%ĪV'���m����1��¨��e�Ѻ��z�sJ(�X̔w|�'HGw��ۜ�;�ۖ6�q+-e;E
\,Bm=��Ii��C��i�8�wD��ռ�<��i�0.�n�N�(͗�u�K�5��S��㲂v#SJ���䖗Gֶmeol� }���ʐ�*C)���й�%ՎRp]|-�5;�Vm�ԑ���!����.��;��ǖ�cL�*qc)�ʽ��Y��҄J:��9�8Q�t��	uc�V�<�T9��U�i^Y�ܨ��I/�p�+s�$��!u:�R���	���<,E����]i��Lt�ӧ�gu:�w7�^��5�0Re���+qVNS��(�r��ȥ]JX�i����cB�I9!t�q��0�v�rB��>�\�j�c���ϬT��:~ğ�j� w�³�A��c�Y���g�In��r^0�-�{9[ذm�IvR�x:�\�(��JD��o����.��ok�jb��a^��1s���t\�-��'bo畗�MG5Yrq�s����֨fҢ:iN�9Z�3�-VR�w|j[�򜜩�jp��S/M�8 �B�[r��{xb�&,��β����6�����.�8�AfԊ��R�+�$�*��ɚo*�s��F�M������ۊ���(V?�-�H�:�Ɩ�؝�r�9��F���E��!g��0��R����>n6"ȵ��[n�y[*X���o5!&+���'Z�۸�Nѓ@\�Q�G}ԟ3��);��$��Um�.�L�У]$�Ki���j��7�ur��ĭK&B%�}Xݭ�a=j[�u��1VT7;��r����=�C��D��J�1.����&>v��c�º�E�Z�a7v����k;��
��p��w-�
3�C���Z������v�[[۫�+�j�7Y+#t�s��.�6���Śe�4�|�I����ܬ�W��m�R:�7X�!�+�&���E�͊���4/�W�s����u�)M�9&խ��d4U��7� \v.��BR폯������5*:�2����ZYNwM��{��Ʋ.���򡘇j}�%Xv�tn.m��\[4ب�s�)����^�=�wmN�r���i'5k�6,k���xBQw�Gnb�QAA��`��k���]up���w�j��P���(R�U�]R�(@]S��)�eN�B�����KX�[�WM���Ȋ��G2�p�b�`���]����q5��/n+�9��N+"�iRs[w;Eb���2��K�R�۷G3j�%.L0�!������|�9��xo\�pt��1;�:j6+] �F�cSZVQ�ݛ[|.�Bl���ٗ2�ZA�Ao[��d��bЩ�x]!N,�Ӓ��!�¶e��Y�xU��C�Zx%@��n�H'�:}���/:�"�-{֮�n���Q[�bvZ�bR�u\4����Cv�oL�2޲h��܊fL�sq���[�3p	����)SZz��`�w_iu��N�w��Q��u���]���qP&>���tcTs�6�u�(��L;6�TOf��B@z_q�;n���Å�lNx)�9bL��+�}��aR�##��Q,T����6e��}���9���y�n%�pm>W)7D�+�Z�T�3��25f�t��a˒�L�����������Jڪ���;[Z��������ҥ��z/״�x��}�o:|uK�9>
��/�}Ҝ�i����fgGI�h�l`;��uAQ�zr&��t%L�4�Q�W}�5ƠN�X&J4ʘ��ݢn��N��YS.�X�r|/{"���E�ti�x����'�oy;Uń.\����b"
j�/l��S3���F�c� A]ε��C*i���wA�2��w��j�o7"R#H.%|rq���-i�&
�\6$��V�̢��]X0Ӓm��wD�3+��}�r� �ٶ{C��n�c{J�uݴX���1�����e�t�=m����u ìB�t��,��=�ؽ���8C�x���+�WZ-MSၞ#�T�	*��7%���,ED�N��s����"䵩���FwZ�+�������K�*YS��J��2���
L�(��T��|FV�	e�{����$-��y�9�9�6��6�&q�kVs4���}Iǲ�x��Q��Gn`��=�bt�k�����'r�"	�ltι������`Z|)Ժ�9�{�.�Y%մ۳��t��qj+)Ն5QU�|9������*��+ji�,}��[��\y6ļ})�mu�X����p�q��>�PU^҇��W�u��v��Yx�[�4H�Wy�Vdv(m*}3z�(�ն�h��L�^��:���������i\}�5�Mp�y�O�	Q�|6�_��^�:��M�p��»+��e���Q;���F^�톏fb96i娎[�N�<�s�֑]"��U�4�Gd*:s9n�Xq;6���ܰq��2�`��'(o*x��ʖ��E�(���m;3�ػMfռ�f�%W�Jx��J�h���a�S0o�F� ��0�����K���$�&� 0��Vw��*vm�a�[n�=� �Z�$�=C[��(�Y�y�;@2w
���!	��ƥA���R<9�e�Y�<#p�$G
���Y��O�������aMr��n�
`��i.喣�Ne�r���ce)�]/{(l��p
�����zƪ_rC�l���Yz�v�`����)��fl�H_�7�٣|�[�>ε��!\^�1�b�7�3�Tsx�!��S)����Yz!k��ƺ�XQ��l�H^��m�8�k��@L79@��*���t2���7[�uf�	O�=�Q��m�H]N��/�n"��$#S4^�#�$8Y�ղ=�8Wb�E��o!�n`m�ھ�k����9��۶i����B�Xͫ�fN�&�Y�Eܩ����IXPѱnV;Pof\�YX\C�JNU�b���5a���}�{38�{{c�i�ӵ7}]�ޱB�eR�b��[K[�\pii)dY+*��
�ʴ���M����)����95�Ǧ�.��A��� %�*ZW%\�X��H�vD�Q��w�F�..�JCu��V�8�i�	YXm���]WN����+�,���C���.���N6��MjN�|�m��@h\:���/N�x�A�_D�*�cb�g�k�ԛ��m|���s*� o�v���~6�n ��4E����[J��(̹u.�:Y	��ڠR%`�e�lg
͖�R;�	N��s! C@Ft�H�D�4Z����yc���3���r�[���t���^,Gtw��  -j�ZY�xܼ�[$�Z�}��V��2��d��/֋�+ t'o��Xiȴ�C� �&�.r������z��H�s��׵�O���9.Ŗ	ئ0q���Ҽ[�M2	��]��S/+�����5������0+�$�Y�^҃kWB���\�-�]��6+	�/��8�O�qb��Q*�����
�-�^%�ΐ��%�U���E��k:����:�82�2)�Fl.�U��s� �������f�bv/�t��n�J�+:W	��܏7K���Á�tz�jl9̗3� +�rkZ�6 ]n�q�a:�.u�ʟH�����ҕ\���v���
���X[�lL���yĎ����\��rWl�P��ث���Dz=�b���z�	ZxwoYe��7�FQ8��u��Uru8�0ϛ�;��;�e+�c���oTy�7��s	��W2]
�Lf�T���6��Jg`Մ��	3V��֔���XӰ%E�PI�oa$�r�Z���=�}O�Q��KN2�Z��D�5�:�k)D�sޮ�UK�k�]�����n\ �-& ��B�t�Qm�c��$�P�KB����b��ʹ�{;��R��i�B��iU�;8y႒�P��������B�d�]���6m.��y�y���
�k�����H�;�ܢ��1v�YoI��A�ҢF,+J�������8CƵ�S$@�:�G��+ �1c;*e$7�ۧ{HǦ��"�xz`�{����V��_[��a]�ֶ�I
�L�PX�������:�9`�.˹�Ra����RCv�uE�d
��[��L◆�r#[9(j��4:�[�hpĬ�\AÀV��q%B���Qw��� ���N^K*WN���N�9ԧ7,����J�+���R�d���R��N�*�M	�k	�8C�����,
�r1mݻ���}��n�I�]Np�j���B�UٸK��e�.�%�K#�W��k0����e�M��HI1r���>r,��FU�nD
���7�q#�*w�,�s����x��^&�G���/8.Gp��W2���.�o���}�N(�s�Q\���6dv �v�2��n�� Oh�1�6�&_�##n4&��F�έ�f�cy/6�UԾ�N_9�D�[�l�ꜥ9�.GvZ�C�˩�x�8���n3�]���*�Xr��mj��l�V���m�N�̈́LW�V��%iǛ��p���k��^���F�r�9�h��1	@56�t���+j�d7����Hk�fI�l[�"%�j��.f8.J���O�[m�Am3H��t�f�sS��%��3�)b���m�x kz���ixfNnK����W�+r�v��u�*��)pq�=(�����Wa+�7vT;I��.#܁�]�Ì[m�H�\������=w�:���:łi�綧N�Ɉ�@�k�����mK)̇�/�Q���Q�g�2Cϻ5S՘�L�U�j�,&�(5:�H��>��̋!=�@�[��7^f��5��!��S�qn�A6�un��ӕ�slr�չ�8�{�^�Nr��{�N���V	wu��Q�ncr^BY�'���'����D��X:E+� ��j=JoTԢ��ZF��
Vƫ�}a	�r�h�Yۊ��w)�94JV��0��z�]Jԃ��m��b:I�2e�t�P88�S�@��|��qP�����5�&	א�{B!��1"�� B�m\jg9�n,��YwQ�65S��%�˱�4t��چ�Ȩ�L*C,R��NY�ި6�U�r��)j,���;���j],����5OF'��J&?�<.�m�|B�Y��Bqt⎱�8a`⊳iVc��Aѓ�֕�{i��s��������{/뱬��4����[�082�R�	�޶i�,�W���P4��͐*QU�;���m�Z�8��:���pη5��f)��ެճ�r�ik�@��x�6,[v�盦=�}���4�+���Iw{m�HGK��o��ᙋ�&��Ɩӂ��&�z5�t�e�����:�C������k&��N�f��sla�K!Ԗ�{-+-�3�U)]M�i&��q�d:�xW;��V	C�CSU��z↯/`6�*Ƙ�/���9�V�2gc�T[{�CE�D�v>�&���c
�s�lw+�w���}�KHej�b*�"q7j�_T��P6
����5����R(��v�6�i�9'�r��uڛ��˛��#W�VŅh%��Y�j�΁E4�q�̫�7Y��r�n��T�!6��{���v0c�sx`w��w|��C��r�h�*Y�\X�w]�RӒX��E�q:���`$�hw̅v����kh:�te�2�`�`uF(<}�E{r��46�AG%�p
��VQYݵwL�Sr幋c��ɐ��ɩ����wn�**�X��7�@S��]��-W]�#�>��,ƕ+�"|M��{v\�jJ,��u��"�*>gsj�k���O}������B����5T�D��eL���\�,�;���),":��^�J��]$6���Ő�!Z�\�<��u0':��:��I�DN�5��n�6��U^�V5ut)�5R4����X«�T�5�Xj��%�M���Ӽ6[ˬ�P�r��a��'FS[/�-��<Bτ�#8f�Lj!�����B�f�nkh�ٌR4UCp���@�.��b��9�Ֆ�=�U��Ф�Th��oX���_J�nȚS% �B>���*F�n��g5ѣIfbg`C�`�P̀����Y���:��ѩ����e��2;,)�B�D������"�*%���3����н�9��&����ÚG�� U,ރ%���Ӕ�^S���A���pM��,��E=u	�װ�����-�5`L�c���e���)T��ESOΥHH9b��90W��Gf��j�m_���SIQ��jѝ�!&E�09��ҀI7��X�s�.��WM�F4���z�Xo"bAٺ`��l��	-��;�Ӵ��%\��Z��}6���gIZ0Z����NX���Cʳ*e8Z�J�뭀q�@t��[.p�����r�u��H^V�[���VR\�UZ��X4(�V�л��^��z|%�n�q�ʲm�u��ښ��b����=B����ji���-�����[��R�+��ǜu�Y�V����b��y�@�P��81z���\��E �.q��Ms������k{���^����F>:Mb\�Č�-V�{�g �KoK=��Q�Jfk��}��6�a|�훸0�=Cn�޻S�ov/�Kk%��
�]�c_S&r�����Ȟhb �_^2���Z]9��KC�2�<7�RZ�Ug��PRr?	7�oh���#Y%�EM��7��K3v�i�n�i��p5�ɰm䢐qi�s3w�X�s�F���dK�m�X7I�вvVD!�ԥ��uګ�(��Y�H7�Q]؞�.I�b��ҁ�v������55�U��U��[�i��AQ j�y���a14��i<���zŚ�N�C��P��P�gX����';vv��5�a*:aWV
H;�u��ҙ����]��t��&�ׂe�ʭF�����>� ��F�|�*X{bT�(�kn$"g`!_u�B�a_9#�U6�uwQ+��Qg�h���$���Њ������b� ��e&y;��e���g]G�c�4�]��5���C�X^�[�Lͩ���g�YH�[������Tuh��ڀ%f� �3%j����ϩ���d�n�! �9x82����R锪gaV��� 5��OQ��d&$!.f�h�*�>=��X�ghJ�ڜ֫��Z��S:�@��v\5��I�Ⱥ�Ȳ�ku�!ݹ��-2E-��VB"6y�w��)�\{/k08�Ȳf3�s�(뗍l�:�q���"�Fj�8���YLw^;
�g9�b���yi.�s\�A�R"Ŏn�=�ru@�`��ښ|&̍�{�(o%�}�j��L�L��	�D=�λ�:^���\�wE��'�VPi���w�ev����Z��9�np\{"�5��bQ�BY�m]�s y�V�z��"�P��Te4���M*� [����"}�롻ۡ�X?kC_;'A,e��:�yݼ�Ghu�On3��.�ۃ	N�H���U��]t�����1���'O[t�,5oC̣���Z�]�Ý�E$��M�I�ǹ���-��[X���r�ߠ������j���V��h�����n޲�3OD�೤R��c}ݝ�<8>.
s��}!G�`�j���pڂ��wV�9���V+�hX�},:O_���@Ȅ���K�8�s͜pf2����p�)��yH�����\�R��'N. w_;N|Tz���=.�C�u����M���T�Ɔ�]O���}���CgU���Npm>�Ʈ��ˮ�im��]�eԃX�Ч�3>���ME���ov�1ί�e��m1!�,�Uj���
���,��	U�K�)dޡ��""W|��H�:���C�J\���*�����:-&:<T ,�������AX`-��-���u��:hc2�U���N�Q+/:�>�.p@i�A]���e�^t��νWE�.�&��
}V��Emu�wf�
wI�68L�&���ٻ�,k��}Ŭ9�j,U�N����2��h����Ug	�(����Bs37i� �:K�ݸ�^�⇭��6�u��/2�ָ�)��K!bsd�W��m�ެ��1gw��U�" n(]d��֮��i]�.�պ��B�}܆�"j�5k�D�Օ�Ν�V&����E5J{j�7�p�9�1�����;w|C��k��V�O�jh�o��Wc'lx���O.c�HRđ��O����L�{��Ҕ�y�bƠu�SWg;1�JXN 2Dpoy*`s1�m�����{
ʊ��%��m�v��$��=��b�_Q]�t�YM�=T��L�Ƹ�&m��۬k]'Tv���N�q;˺�!S�y�]��76|YoZ�ڡE��͵���.��q�Tkx��T9�ݑ����g��\po��Pm,���ّ��$-�I�̻�ݘ�G�r�����MjJFR����ޡz���%�ۊ�_@�Ky���ݪ ���Kc%�\�)�\wx���e7ھ+��Y���ݎ�t�#���t�h����:��9<N#�5meXf#�W�[Yr���˱��e�.�un���>yHr	ra��k�6Ow�K��*G�����������}�*�Gپ��y�Zr:(ǍW�
}�.*�	��*���d�eC��@���I��67g�v�+WY�N���t
��z1�]2jKkQLӬ�k�k/vA�h�C��	��j'h���owd�Џv}[Ӎ���E�A[l�S�.9�V����%d���\�;ByH�x]A]W �6];��OyDmLt�8�I����8Xl�wn�]���G2 ��r���ͩd��&>z]4pBJ8�^A��
<�[�.߅sΩ�fP����UG��;�E{��_gX�C�H{�E�zhmu\��g��m�-Ƒ���i �(B�T�1�}VP̺��](q T�9rjrc���ī,X�1i��ȅD�np�%�;�V��Ե��F�k��ub��[�)\�-ʾ�W��Ѩ�3r�H3�kRY\��mob´B%-Y{��2V&�-�ˠ/7�T`P��޵��u��;��m�Ec
����w7����4�ح��w�M�)�*=���n�d���X�z�n8Z����Yc���]���h�7�ڦ�Yk٘��qf^dF��}�e�R;��9n����X��r������s�m��I'{�ĝ��z�GWH^k�7;w%�������w�0�y�NdS���ʮ���ؕ��L*�.��o��� +�˥��\�s����fsO:�\k��o�j�;2�L�q����P�q��ޢ�I0�b�)ͅ4�F�*����R\�&"e�pL��$���Ӻ�c	A0F�BBFJ�B�wuI"I!1 ��`��
�c2L3wq��A�#�#��D�wv$�d�sB9����))D�� �� $�Y��p�h�"1!a��Ш60%wn�&H�M��Fܹ��VY�%$��QeݷJ0L�1�BBH	ؐ�FEAj,�Y	1h
#Q&�i,�Q����3�!��I!��F��4f��
z��6�VU���OFj	|��GjӹR�f'�l�:�N�M1�U�Gx���Ev�媥<��4������~�ऑ��w����^�a�4r��Ϩt,�Eu�4�m�9�R�Ӗ~�l���T(nv:|�S�4k��/Ц4J�Cܫ���B�:�z�{���f���+��P{���n�:G}�`�<��32��S3�Bd�_Ѭ�U]��1Ҩ��.�/����b=��J��1����Ԃzo��l��#�C�18=7�sKU��Uaq�DI�f�"�wZ�uҦ��70��$��d
���^y.��Nqv~���25�c��.#E����S^��5��RnL��{oh�G��iῩ��C�>Uθ������B��ϛ;O��r]�1�p�X�ܙ���z}g	ݲ����\��� =5x[Xx �s��{�~��:�ELg�s��߳5�;�(�{l��Y��Q��F��WP�U�𗧘L{�Kb��J	V|�OOmHk~�L�]Qc�>F���5-�v4���n�n^�3V�f�������v+�+�u,=}{�*}F_x���p��� n�t4��~�)<�^��QW1�ྂ*[�x�Ğ�ħNv��K����9�R��C�_gh�&�#� ��p¸�kB7�,ڵ)��dW��nLG�xM���f�a����G��bSBJg�;D�t�k\��)VPe��O��ff�J��z{���N�Q�Q��]�^˺~6��U��epQΧG\et����9��h1��,�e���OHF���̼�Z ���G"B����٩��.��%[���l�o}t���/�p�x])e�����}�Cu�@hTg����
�r:#�y5jr��F18�)�]T��N�{<��p{ˠZ��TdHУL ��$i_��3�������]u9ב��Xh�P���=�l_o��9��6�);�"��U&6����6i��/B�!�h�*ե�9���*kd��ي�A0�M��y�fLu}s5�ܳ���
����o�Ǥ����x魐�sù���H�p���.BN숷���������� `b�uƢ��z�u�ExwOz�r�����p�5�Gó�}ji��v���쮱yQ�o�E�VV�z�C��w��$��/XlW���e�HÅK��aM�6E��|뙱E=���ވd�V��L�{�{ۃ�<d�M*�Y��\:���/j� \����x=�\�t>k�N�6s�>Z�ʐ�6���3��q�ԣi\~j<�B^�_bx�-탠y�V�ﮧTT��=�������b���7�#�j��/qK�iV�9)�֋PX��O �ɝ@]^.�n^Xr;R����K�7NC�����"k�+�7��쵞�t;t�z���"��@%�IfuT����5^���ay��l-S�/��>�Ό�2�����~S��p��Y�x���0�'������������M�,��?]���S5���r�E��6Aj�ۀ�8�L.P��S��:�K�l�m�;]	\nLd��=6M$��S�2��pʜ��P�ч��>�ѓ
ysE�X�y'�kI;ꢰ@�>Ү�POf��X0�hT�W�k�D<��L4Ԭ���Y��$r�����{;C�r�ҡq#2C�����LV�qWI\t�4�c�����	d�}��`�Ͼ�P��x\����Ѐ>@ѓ(R3��uϱw_�v��[�Y�ާ\/��7��T��j��{ք�LRʮT���G��@���[f#��+j�C���m��>E����!�������:a��� �zy_����Dt���Ǳ^���m��bNr���3R�%N������}
�M?rN��1���)��2c�@.m�t��wF���l�@��wNj��u28�����[3�v�P��5�e��Hّ{�'��{7ˬ���Q�t^�<�UB[Tļ��-�y�u}-4���d�=[��Ї%pd�@EW������X�J�㣅���f���M��o�;o��k�D��)��w��5���HaX3
n����I]��ʪ-ә�hW�3�Q�6sncv�g&��F����M�Xj:=��W/��a�����Pܵ��g�����1���V�{)�M픺� 0jk�ܘ�]�m
~��cС!�_}];�n���=p.9G}��}���yp$��ff�sY��f
�v�E���H�c֭,5�'[�p�*�谩�T������4y	���Pn��X7�6o���LvJA���j��k}6��ӝ|���9R��B���z~=L�*�ls5s����S��4/�����;=��|���9�yͰF������5�/�Lz^���1���1����g��@��({��9*]a�֥`�d�b&aP��G��iz|��u�%�u�ޣ^՞._f*�Θ�\�ǐ��/�f
d�������0�,����y����.�=����⎸7�Ŭ�H��u�u^S�ƻ�`��@�ط�hW�f� 9d04>����0�3Ɓ���O�S��0��n7�)�Q�n^Wf=���;"�u��Y
�<Y����b)}^7�S� ״�Cy���F��fZi��>�7@�Вe�])���K���GԤf�5ӵ�^�vE�IN�T@㖉�Gt��υ�V&l�Wv0��][o��H`�Nr���A쌮QN���p�C��>�S1�-��Y��r&7�x#�T��	2�Jp���'�;���P��^����Z��d�����3v^��j)4��s�z���ɝ`����������9���M>9"m a�C�9�=�n,v�0��m�>6�s���"=.�����3�ia���;��MĮu�M��g�C3^���{��+��F <������3u
'����G��w�k��\)Vo��wrl�jB��_t����uh�Bg���67�"k�0Oφ�ڹuո4����5�^+�ݍ�&�I����L�}��`y����
��y��[�1+�*�z{"r�A�M��8k�:@���5��g��z�p�N+XZ�sK>�)�3P���k��^K�pr���i�C����s��gy���J,'/ ���������g���E�[�ֈ��x+�MKZ�*ߦ��)�h�QU��d0:wG�U9p)��zD�G�D�C&5���ۣ�ܛ�9�h���$ɤu�u�2�wXh��
�[Y�hCK&����<��ub��z���FzW^^�_s�̺s��T2�0]@ٙ��������u��xԫ�7a�7��W�+�@�ou:��m¡�v��qDv�K�p\�jJ�*�\��:�a��$��X�{4��*'EF|+�j�xW� N[��,��Ô��]�[��Z�."�S����эm�싮 B����hס��N6O��֮zƧkbu��k䲻�ٗ��:�0؅M�����f��J��9t��鏨.�����%5�X�}C��G��9԰�dh�N��ÙB�}��l�;��A  /��=��5���҈P���T$.
G�BA�M��i�u:;O׿6a�;�C5�D�oN�ke��s|;��P	=�X�Q���¯���B������M����H���d���J^�9���A�]�6��dT|_ЊQ�ɀe\=(�K��e9�`xy�(�̺�Hਬ��Y�����y+�<�՛TlX��2�����{��/�h�K�n���s'{��F��'��x��r&�ɚN�ȵ�<�X"�u|��k�wMzg�˶j�m+n9�������I��&=� 7� �_X
���8����1�W�f��<�,$v���
4�G,8U�pbvp�I'�ަX棍,Q���5�p��=p�U�ge64�yO�Ǳ0	8�P{�\��N��Ar�n�6�_4�Cp�[��a����Q�X�JRK�/_wQN\�f+O���Iʏ�]�Q�Ԕe����֖pͮ��'yp�'vD_�k�@��8���No3:&O�pr�u#^p_��d��LۮTk�x�Á�,���&,p���+:y�������MUcʌ0����Z�D�4���ȓ���C0�mSU�X�㯱�ዷ*�n�����W/`���ֶU89S�0q�O��,�d|��$����Gu��V��ͥ\ ���ۄ��\��U˚z��mB�p��u?��v�|�o_��R��K���֣�`DU{F�<C)w:�v��ū��,�(OQ> _��p���}�<k��l)8��:M��&T������͕����I9�jK�K,V��a�'��z�¦���Npl)��h68_Tk�[pVk�d���"�6@u��Mw:�Tf˧?tc�T�@s(i�W�:�֚�/��:��D����!�x��(zM*��IA<���/U=K�)?e�݈���U짫��Q�DE��b>�"2&R���t��U�I���b��U����Z����
(���V�[Q��,V�=t��8��~�B׷B�:,���Eu`Ù�]e���(6�CM��i���n?k�KW�d�ڝ��J@���<�X,�;+:�a�n���O��דE�w9����H�sV_\
�(n��.5Y�Sq�|eEd�F��"w�㨙�t�|�4�� ,|��&P�g��.�<O�3Ӻ�X}}}�T^�����6[�L$3�X���hK���W*D�F�Ed�DO�l+�9���͞��[z�s���H2�H�F����σ��6� ���&8���d�� J�;�U������寽O�V�A�4�����F�_ܤ�c�v�uQ��\d&gȪv����ODZ� <�p$�t���"i錛�O�
s9����+�7�eU6| �$�a/x�[�����}��r�В�Fh�]/����n��^ۥ�p���:��h���d �E*n�jߴ4VA�E���[=VЧ^���ܾ�P��z,�Ɍ��b���&V��`�6�o8�۝+���E�͙�s__%�rὼ�D�}$1���77|��`<ϭQ-�7ww��e�@1��g��o<��E:�u_f�����F��zF�ʧ9u�|����x��Rn|����ߐ�]i�
��8�������N��k5�Rwot�@�V"��X��(�Кy��������I�6���S�4_.��JV\�2��u2"@W{������.8/ĵ�SO�vVkن�K2I��M:�6�Mo�7��>r:��%��t)�D�+�:������Bl�]�>dW-R���\[tEd��h�@�:�|G�br��+����s�lvz_ou��(э��6e�F`����t�������EG��旡��
�U�%�a�^�ޥ^�C����c�7��>v�XR��Q����L�bu�ßB�/(��hy����7�K�q�(}�5�=0y�D2w���9�Z|��iw�	�ܭ�=�~��{fl��Ch>�-����.����I�-���s���p>:�ׄg�:��1m؜��6��b�D�	�U��6s1[�젶�
|`�P���|��Ȧ���h�n�f<f+nݰf�i�[<�-�+3��W^m&�[�g������b�*���O�;ϧ��mXc"$M�g�.� �QI���؛p�U �AqJ�����ML���ˠ`��(����7���g�vV��Qn�Z�vPגox�E��"�#s��U�E�
��`�K��r�a�*�{�%xX���k�{78���D�����x��0D�F
�|��m\�<wE��2$!gqc�I��	�=S�]�)�=i��B��a�'N:�c��B[���{��E8��@֭]�m����W+���c���9_!V�㕉qx�:���#Ԕ���ˏ�����1�+i����tsw��ę�ru��)�XI��+]+�I�qp���d�KhJ�璘Ev��ۇ��g�x[�H^V��J��*�_����o���Gs�N���J��ޣO@Ѳ��ܼ��z���N+XQ��4�] �����u�5����a�w����f�5s�1�)V�Nf�-�D��|����W���)�b4��£v6�w�d���M"���ʀݺ*�T+!�u�಩ȓ�L��7ŧ�9�&5J�QnԂ�i;�x�_i�n�MƵ����x��� S�E�<�g�|`��	����3f(�_Т�mRJ��o¥�80o�_ҳݶ��P�G����Y�3���}·V/{��:�4��êA2�0��O�)���6"�.w!���H��:@j�f�_C0�����oN\w5���eL:<����c������q����V0�'kf�H	P�۸3*;��S�k@�\g*���S��~A�M�s�ibpj�+��1�f�mE�#zݜK�N�]�<,dL�o��� GT�O�J�y�B�wK��M������U|&P�hڲ6�����|��*G\F��@p&�E��) �?\bӧW<�/��>泻ѣg]���M8��[��% ����ˤ���Z=n@P�F*�k5�S�1��|9`\��[�H�8����!��ԨUa��#Ip�˒�.���uu06�ѥ�Juî��|079������Y�y�P�(6Z2�>و�:^JS���S�G����������v�Wτ� S;���J�I�����(�4l墻�ֱ���k��ee��3���z�_qFE6���A������
��C;2��&qG��j�d59ӿ���+��Z+Y먞�J��#��d�Ha��[X��2=	N���|"��N��PLJ$���'hv��Y��(����&GwR����-�K��G	�.@N���L�_�e�u[��,�R��.e�ĉ)�N���Ɏ�m�.�gs�s+��#v��Z�{��SpM	w��ͅ$��Ey���Q�����=j�Aheff-�%j;���(h@P͊�h����'vs��b���e�����K�Vr���[Y6P�:헊ȑ��3-��z�`�y@��U�JqQ^��LA]6������s1����5�3�r*��+T�q�������[�+
�x�R�S敭�# �(�ק.�V�u��͐�n0�s���@�|���v찳ft;z�O��VoR��dϚ��
̻F˙�n�ִ�� _1� ���LZgؒ͏d{[wj�qW��5e�"l�Ṷ�#��n�.�"�&/]_�q�)��Nq�m�pԷ2�W ����S��r�2
*J
�ViUi�6�q.�/���8@1�����+�(
��W�;_mbeP�1^�G[@ŭ~�Y��Ɂ���9�nf���\�&l�tt 8f���ad�`�bP<��Մ�d�����&���I�7A��`��t��5'=����pfu��2V�o`�\���;-�q�H��Nwe*�A��u�=d8�_3��Ȧe*"�Izs����C/��7�X���*��1!{��I9c��Y���0��b)Y����D�]�$��kE�N��e�ݴZe�Q�,^�n�,W6W*!@f#v�J�p�X+4ɕk��*tx�&�4YUHR����s#+����B�����
sq���ge��*9���J�y�*Y\1RX�T�D��n���1�f�\>+%>�n)ϵSx�w}�T�J�p�sr��WZ<��2_w!IQrS\�Z�n� �&���-��@�L�d��:-v8�i�|9>	c�nVt�#�;��t�mt9���RyHgUϻ.�_�X�����K�̨	syY8��]�b�;��y��Ȧ^���[��W`V��\G����Ay,��r?fVM�ɮ"��Źx2Tkw�}�+y��:4DQ_�ᕥ�w��d,�U��7k+������/i`���PQ�PJ�[��9З*��p��{��_��߷���^ș(�X��H�RiL�b1fF �2c���H�s\*(���"$��͒R&�ف �PDˌ��(��%H,�)�+2d�P�&���,f B�F�&a�6 Ć �H4��IeBY4�r�i�1�]���$C
�-��`QI��L�@����SwqI�,1���H�;��CI�(R�G7D\�"�i#Db�˙MÈc@)�)-)u۱�"A�k�ăh�\�0b���Ć�F(�� �&��O��_�����������[k��6���d���b5�.']sv�wYR�-���}��KJc7N�k�.�
�h�4I3��[\B݌=tg������zk���������_����^�^/��owί;�77��{��Ү\������m�W.W��[�~��o������_������F�*��|�?}�>���Ϭ�o�Lnn����<�^/��o��[��<ſU���/?�}�k�~�����W���Z7���^k�v���W��s�����ߝ���_��Ϟ_Z�����[����|_�x����w�} ��O�p'��ֺש�J���H������������鷍������w����}��j�W7���s�|�ʋ~��7��|���޵������[�������n|�����k�������}[��B�#je�ݖN?A�у�>�B��~�����{����Z�{Z{��!G��\c�"$D�}"��?o��\�/���������\���^a�ڹnoW��=��n���/K��x������6qM̽�fӹ������8���6��=/=�ߍ����yo���o�Q��#��>𯘱�o�v|�p���>�^��W�_��x�~_޽lE|^��}��K?|�}#o��X��G�h��?}3`L(�1<կU�pܰ_�%��D@\ۿ:����-?:�k��7�nU���u�����m�߾�������Qi�$G�"����A�Ap��{꯾o���o����������{���z|	���g=ǫ�E�P�ٳJ���>�������#�"##�1�H����w_���o���?Z�W�O�~W��,}_ͼW��_7�n��[ү���n�����Qo����<��p��G�#n�4%˽�b�ߵ��_Ѕ�����W��痦�ۆ�u�����_潍F����~��{[�z߻��+�+��_�������o��o�����߷���o�r��uy������C��	��AyVk�糙������W����������j����}[�{�}��_h���\y�ѣ�x}�F3�����x6��׋~���W~��^7�ߏ�zo���o�����������	V�ŢbHs[^z�`v �� 
�����j��lno��[�\���������*�;��_w�]��Z~u��k��+�o������ϋ��m��6���ʿW�������m�����>��\QVh�&��]��K4�N3h�.�޿����9�;�Jx|�φFe��jJ��1Z�j��s��[�clvȾ�fv�j����+N���8��ǅA��,��"���#T�nn�د6�0��oB.5;@��҈�p�Y�iB�
�����T��)�p-���Ѿ�����>�>��:0����} !}m�v��\����x���{��ӻW����^7��^/�{^?>}�W�������}�������?�+Ư�;��"�
���(}U�{�d��yY��w-�����y���~�͹�˛_�{[�v�U�\����k~^�y�����ߞ����m�������>y����ߍ���h��ߪ�z���©�J����s�hoĿ ��M�Ţ�����[�^�o?��+��깼U�\�5��y}6�W����ץ�>5s^�]�^���w�߿�>z�[�ەz]���o���ۛ����&��9��>茉���[�fQ�=���Ž���?��7�~<}��<�������������|^,QQ��7�����v��������\�^����7ϝ���+�z^���۽޿�}���1S=ǆ@�M�Z5}w��RЯ����ۚ�����^������ϽzU���o���[����Ͼk���Z����߾W�}���үϝx�ۻ����Wv�W���y�ϝ^֝������/�x��}���詭���z���:p2�����zk�����/Ţ���-���ϥ��A�#��NCJ"0E�}���m�����_}��{�\����u�zm�ϝk���^�z^-����ۛ�p��YϽ�kЬ^?+�"r�v��|���5�j�z��_�⾭߽�wj���W��?ޫ��Ѿ+�����}k������� ����"ژ�Vc�"G�~y�j�˚��|����_[x����_}W�_XC�>��W�j��R5�+������^������~�m�ەy�דo���?{������o޿{o��^-����z�ֹ�-�_=z潷�����}^�����ޕ_���_<�{_@���G��+6 t�J�Z���%)�|^��W._w��5������������o�{�����Z{�}��{��5�?GB��>�'�"8A>�g��Z-�\��|��o���s|�m��|zHG����7E�7�Ž���	ؗ#��wm����瞖�_�{���OޯkN��������x�5��h��Z7�����y��^-���ս?Z�W�~W�ן:�c��5�^�|\ߍ��O�~��oJ�G�����S�ko=���i@7=�kFeE+��ŷQ��[v�+�S&f8a&�S��wR\�:6�i��hM�N��)�ә�}�o��z��FK�t5�K����:��I�t�Uot�F�Aס���堾HA��s�%-���U��}[:,������H��
��mDP�>��ш��s}C����5zom�o{�����^��w��+��/��k�w��k�꿛��y��_��h���~�����x��{����G�"kh�t��vP�9R��G�Z}L}B"D8�k��X��Gх%�H�>�U~k�Ͼ�j��ڻ����J��z������/��m�{�}��^�ޛ���Ͽ<���w���x{��W�}o����?z����,��g�hR�������=��E��j��o���x����*�FE�(�b>���yL���#�DG;�7��m������׵���������}W��z�}~6�o�n�o�}U�^׍�j~�mz��W��$+4���I��d�G�����u��E�7���/?z�2(Ǉ�"~���!q�>��|I��K�
�U����^�����Ӻ������񾯭x�7�;{\�o���}��~��^-�ȕ/�j������䌧��#���W�l�����}��zU�s~4]�o�o}\������}�F�+�;<��~+��ۗտ���絣sntg%��f$}}�;����b$Dx}~n8
�Ih��^w���.�<c�#�#��ׅ~��x�^��|W���_�ƿu���k��=o;�:������ү����צ�/���5�����+���m���KzW+�n����>����o���,N?�a&���d�g��)P��>���~}����m��o|��}o������~���Z����<���/{����k��^7�޼�KA��u�+ŧ�׿}xޛ���*�����o��������E�ٹ�z$9U���}*v��DX���Ϟm��[�[����������!A��HxcG�!F�����_�Qo����z~6���ڿ+�znm��>/K�\�ͻ��;����Ak����(�N��ά�y��h">�1#�u)}�G�!��Dg��Q���@!�/�����D����(c�o�rb�n���͠���0T	൮�Q,�{�K��fv:�%�"91sE}|��Ȋn���Z1���񘭿�ݰf4̾R�P�\�dD�F2�9��
��p������lؾ.���H����MW��;,5��Y��;�!����U	1x{4����<α
9��S�ʥ-�S��aC�q����[�֚�Lس{0
�I���̘s�����t���jD}E�l���B쓵cѰ&cn�]������h��� �ڰ�H�@T�a�F;e�f\�t�L�t������렀��Ⱥg��uX�{$hp�:y|<ׅ��D~�Oϯ}^��Ǆ�@��E`��>|���� ����h����^������>"Z�l��G.f�����z{�ٺ�:s:�S{�q�&��q#���6�z����pvn�}N���M��LX���0�#�]���̲/��ҙ3��������ӟs8����W�*���}�e�s`(;�ƚ�UM���O�G|5�9�Qb�S���=�M�;w��b]�Sn�5�5�b��r������Yo�����a&y�b�޺�O��=n\˦1�q�Q����x+�TL��U�P����i῟/VUθ��q0�E9��|���}��������9�6v�X����=��&-�7��*������ U���S��[��m����g�]E�.c�)���ƺ�?c[f{"�PH��B�.��E����,�L��%�d
pN�o[��������$�����^�)��n�{�X��+�%���3
 ���)V����-�z���Y������'.��5��r��e�rk�s�y{�Ԁ�X�c��r��B�*+r;�t�$t�菣�x��i�_�OP�sס�V��b/�h�܄v�u*��t�^]�Y���N�A/W�̭쮲B�t�!HB�������:~m\9�/�}�PV��[F�Ҙ@��緭�m���6�,w*D���}����97�=v���S��8}oeUM-Pȴ�׫˺�ث�Cl�ܢ�* �� #�z'��s�BK�_�C��*��ߵ��\������AJP�VIt��ܿ�z���"��X��={�9�	SC�F�T���P;6Fnt��+¬Y;_{�z�粝���� i��g����7�6�4d��A�x��p�ro��0�3�M����J����rU��q"ap#j!�:�[�o���b��Sk�z���q_R~9��(�I�E�l���`�Ɏ��f���g��U�cd��r���5 �ΘsssQJ��Urw)h;ח!'vD=*�1�;#zxZ��>��9�5M���m<�Gxe�[B�8���4�����O<��?`�ߵ���<όT��NȜ�ɫ�Frj_%�ش7g[����V[��74��W|�j�]�VK��gjg.�����rS�:�Ҳ��bjj�T�e�;���*�w�!($jY�0��8�m�b;��0:�ѣ�dI�7��{��:��_�ﾪ��W����89S���+���-�81� i����]mW�t8`9���[U���U�owU��>�rM�����YΌ��x��S��8�h�*	ݯ�9C��	�9����t�l8��̮Zz\B$ڗ^
;���1[O���b�Z�P]v�#!�/�ȝ߱{�7|By1��t&-?c�s<+��i�[=���G�ȼ���Z�5�!D�fK�׾m�ꠔ�^�����#�΀��64~Έ
s��m:R����Cs_�w��[j�>x�<����:�w�i�Tf�e���8eN`s(iQ��f&���y��'`��q�_է�y��P�<1�\|��y�^MOR�9?H��T5�f����K��t����k��a�G�囥@I`i��w.� З*T��k�޵��ӥE�FWlS�����|7a�'xc3{���Cd�WL̩���d|1&^[���6�F�#,wf.&�0cu�a2��.a ����5;�����Q@)F�D��ʷᣞ(}���%b����OU�!�����d'F�%�mm��}��	�4d��q���T�&�<�eg�rs�i	�{��_
r�Ӄ͆g*��-���x����l���"�h�v�S:-/�W4"�M`��q��s���Sl�p����DG��r�n��Lǥ`ك���C�~��B<���t��uV�Y�ٓ	�`�D�d������E4O@�}Z��C]�Kʸ �	���{���U�hA䝆1�Dc�OL��,���J�;(tci׾������H����h�R�7��6!Ng3󝄕ٕzj���{6u'6���
��S����ۡ�[�Uk+�}y��{�:��T=y+�v�$��!v����a�7Y.9�s��`�reVէF`��,��� ��$\�t¿���is����Ӣzf*j_�1��{}9T��&fa��%�vC��1	ኜ�����L�7�=���c�evoPRZ��`TF��U
�}vG<��E:��K��g�_���F�"��j�y��dVt]�|�
4A06Ư�6�~C�_�x����^sƆs��Ƕ������'�D��ˁmJ�S��W����X�\-�+O����\�/��7H͠2�[�𣹪p�Y�5ˌ���������vD
���5â������\@��HA�^���OY#�����x�U�.��ǯ��wV
ymP�#;�ڴ)�) �.�ɻΔ뵶x�Mu	�Pw��)������_B����L$ܘ[��]LeJ�:�/GpxMݪ"A�Z�*�z�
�7�_=�{�b�xC�7Y�Z� 7�F)��a{�D.����ꪭ������r�|�}�B��e������UuҺE�@� �+��B0E$���{����SX9#Ct.���K�8�x25Ա�`N/���ط�R9f)`/,�>�RaM
�n�4�Ү7'�����im�\U)��9ZѮ�cm�&�6��:����ʯ����,K"u$'r�c�T�ԴbO�!!��u��E! �F7Q���V���|F�LQ�@�Oy�r�e�cѶ�n���gjaq�_ϋG�{`�{��}�e:��=OgN; O�d���W�k��7Q";��N�"��4���䖇�#v�\�����^�by\�������s:�f.g.~@�#>�@>��0iq�.�9Q��m���2g����j0l�������$l����Ja��jEM���4�׉��B���s�*�lR�T��\<�
[��qx}H����M���\��"�0)��?Bd�^�9UlD�A�w;�����Y���|������j<��4�<�Y��h��-py��d������W�1S)�d�����C�{�W4��{S��}��:rh�u�/p�T}H_���4r�6][綇W�� )�Y�fj�/L�q�Cx�n3�w��w�j�;�Z���|�fe�/n��š,�	\�]����7nY+�њe�W0�塨��+�5�n@������������w4�T���w�&�T,t�x���X^R�����
r'g�k�v�;ƨ�!׏�_Φ�d�ӬW��a�yP�TUx*��n��t�x�	�G�L<����FkWv4��8��pɍ���g��mi�kl��c [p+�㪣��(W=���k}~}����E�Ffa��f������:������:�v�>�	0�{�1UfM��+�[K�.��I�(}q:��ʥ=q����L)ui�6"��q���H��:@P7�ncT>��"�7ę.�V�kU�كC����4�Nތ��R�њ>S��p��
������c�sr���}b���MD��+�`�r�iT�s��!��O��!O�o�������پ����Y��04a� ��*B��[��`�~�,+��W��\�/:���}��ʊ�"�'7�t]�p� ����=(���0.�^к�n*�Y�$޲���E錨R�n��xy��+����.���N�puк�F�{�3���U�池^V!���u�.�ܕ��kT�L�9Bd�w�Kʒ��,"�M�0�#K�5W�=,V��)!�]m<ֲ�ɭX*v�\�)\��⓬J&�Bs��8ʼ��v���a����e�+��Mp}JP��I�k�+Dw��y���� ?}_}�}�B}ܜ6��&��^���E���t&�Hx��r&Ќ��N�ȿ���U"apY�
sk
�^��T쇺��@���La+}����Ƥ��"�m��y�=_\λ܁X��u`�>eIQyd;�U\�yY��>U���y������'vD_�k�@�N$i�
�ܬ��3rr����t�L����D<uк�3�^����_#eu���'�}\5�1��U[i۹$Vl�Op���%F�d�� �[ϴՆ�r����݆i��Z.w� !kء��S����|�1����:3����N���4x좫�_�u�լ9� �<o�-Ǫ{6@���36�:�0�nC�]M�K��C����R��K�����qPU�����SR-(���pDGp8O��u�HT���Fm�p��G�b����
Jm�:�:@�8p� lـ��[JEK�,W��<�38�3}��4~�,:�Y�1���ogL�h̞�((�P�f�\#
�Ҏ��)|�¸�˟�2�G�0��u2�a-�e�1�)�x�����C���h��;"��c}}{���8��Q:s�I� �j�.قqu�d(���f�VձS���N.4�}��"��mE�oY��PT�rb�^]I�{��5�m!�PP��;餝ċ��ju��a��<��|�R7�Qs}��tF�(e��$��o0+w���VVndcb�.o��A�Jť�L��W���ϵK�}fh��n+�R;�;>�Qt��lV�k�e�����3���
V<�m�4�9˼F:Z�����F�K��Gl\�yW�5��r,�ַ8ab�V&4������bЖ�9�IC}��#��m^1�]y�@�j�.�EQ��Ǜ��۵�����N�uܫ���8'HrqG�.�G(��.K������:=u�wo��C�ZRl�A��*�]C׼����ա'��u���*���oE�|�h�H.���5rJ�U���N�)w.Rk�KeşDЖ�\���3oL	Eu��4b6e�9JS��Mi�y�@�p��<��� ��ba�[i��c�;��D;��=�M�i�@TGP�r�j �K�*�N}�f�
jǻ!lh{������մ�sH�ܭV�tmb�ZP�Ŕ�M�5h��:��8�v�#����iT�g;fUވ$�宷�;D�s�S�)3)�{�#S(�yr�AOBS���<[8x�4���Q��ɡ��k�$�xkSՉ��H��|l�����@�V\�a8��F/�Y�����o;��]��|�{K��R;��tK�{+V�u5^JE�.C��.��
0؆��z��;s^f��E=�]V�3��t�(Ү�Z8jx���Xn�1�|�s8%��U�$��4f��2�,M����l.�ӕl��t���MJ�2т�o��em�f�X6J۶j��=G�R�GxɕҜ��v	S�ñ�ߋ��d�^����]_ks;c�Z�4ؕ���r�D�U�(�<$[�{�Q[��is��FU��_�P���/C�0���Y(,^K���}�i6~�ת�_���6!���q��ؕ�_w:�,Ptݭ�M�=)HUI���t��4z�<ˋ��0��&�S��T��1˓k��{� ��pg�l�F_>���c���V^Jwr������^�ӝXeO���GV8�x��";�Q�z�q������K�ָ�z�͌ 3)�"T�sb��n��r��V5̧���x0+�&�n�V�m�ȋ3TQeu�,ڌ5�έ)���m;j�:>���ҙ���1XGT����/vT�����@��Ci���;��h�1��U��ƧH2�|�Л�8�P�v��JL��D�mf�����yO0)@ ���7�ƕ<��/q>k�@sMl��B�o~d���.�;c�oҬ����]�m��[,⑥L����2���k^��.�r�i�ɵ�I�@��n좒�<z�s����B����t�U�fu=���B���4��4�F`!BJL�b����PlE$j�HƢ�1�(тM�BXK&*c1b
�(�lFCQcb(�Jf ��I���$	��F&��@�I��-�QD����fQ���l(F�P"�3&i�J33J�#@ʈ(L��%\�3#a,3bS��b`H҄!�M�wLL�Q$4D���Dh���t��Der铗$�D��A�'uɘ�ە��DD�� !�3\�(�l��'u�"3!-�A4<u(P8��(�j�������t�N�w�+�Dj��[V.|�Ѣ��>`N�ŝfm���r�
'�ⷎ9��
��������թ[��m7�K�i��3?j<*&*6��|�YwPeݰ��'!`��X��Tk �[����Rog%�hE�c�CnGH��fp���~�R#bO�#2`:HE�tp�y=�{�=8(�Cb��>�]#9����q�;����AM&����SQ��L ���ܘ���E�Ά���i�ɨ\1w�:���H1ur6wS���QU�����C�)�櫚��YL	��9��9�!�84F#�[C :��r�(�0vgE6Cz��v�b�����N#���(��vC{�Y��ׂ8L4����$hu�S�����Nm{���^�$u������o'�y��H���u�t�]`<}e���~��'�MuC�#�щL��'�^ {����V:{,�.���t���N�J�y�����YݮVf��s�'gT�r��M��71p��`�reV��'LS���hS��c�lz;��N۪�=�8 �R��d���Qc����s�"^��30��.k�{o%��*m��x��+а��Uh|�Q��^;~Ƣ��J�U+����7�.({�Χn���h�̻��8�8�����P��{�N9)fI�ļ���}�9D�����h&r�dv��7��o�(U��}W�B͹|���
�1:
M^ˊ;��<i����S��������=�������~E�_�$C�}s�G���ul�1٬��Mc���+��}Γ͔�F�{��t�RPc���mO��WU��_g8>qy�U����k���X��$���ID�Lako|j�y`P�¬T���o�i�?&)�b�׃�i�0�Op�C�Kw^:�m�q�%$�!p�����8Amm�r�P}���G��^�������-��U���oS�-L��Nn�u@�6��/�>.�z]t��@� �+��B;�]嗚���5�cƫ%x�7>��k�b6��feh��T�3�󸁪��� ���)�S}q������m���렃�+�<rNʲ`Zg�]x.��cO�݉���h,�c&zuwJ�ͯo���v�`��Qu�@j�w�
<d��-�켦�z��d�B&�}��N(����z��7�_�.�Kk��* @�@�jb�*������)�ln���8H��mybh�����z�N���w��E���(z�a����U��+�Uo$�`��(�M l������0i4z#Ao^���u��k5�zy�z��]�n��̬�ɡ��M�x�k;a�5���=�<���}\dӷ�wt�|O�Y��.X-�0��KQZ�k���L����VDVz���ru�3�v�Ԩ��菾��V�{��F.��'��ۯ�u�4�9�yLd�Be���V|��C*��N�F�Ǜ�ܺ�V��!�QBU��{)��o��f�g��� ��g,8�Pц�>#�2^.����h�dC7��C�j�7�3ZO:�HhB���ؿ����X�6Vr�b��Q�����9s�n���M]ҿ�ګy����Ts��cM|��{E.�S�;��cum0eԕ��A~�9�f�b$�?�xE�Ń����� luܦ����q&]P��[��z���ޑF�z�6��c��q��d�u3.��+!�ݧ�q�"��o���W'eu��s66ʑ.8��'1�vC�|�گE�j�[���&-�h
{G�BbL��{�㛣˞�`,� ���M}��7D�sl�ㆺ�8�ٞˮ 2D���<
��u�u�ҥL�g}���10�R�ʧ=��gp)�.��lE��g�꘵��K�5�˲g'��}�缴�΂L�V�νt�S�|'�U�^�:�2o�t�K��/p8p��v�����:�JiI��7V.M��+����'ۭ��>��V�$�Um�ɴĥPZ2���X}i4dO)���y�z�7)p&�li�����`�p�j�o\�MZhqD�;�*M�W<����,=�-�ĳw)�@Ɯ�c�GW�޹�\t.k�U\~�>�>��gE�%2�� �N�<-�爐�P�~�}%��j�������s�|��C����7+�Up�+�Fx�(�H}�0��G�z�� U@� ���<)\�B�{*j���-�q.s�n1����[���p��W ��N�0a	�j���d�4���+���:����r��(S���?rj��xy��#' -��7��2$J��+���6A��pΰN��/�ʦar���Ț����W�àa6zCsW.D�!3_'v�V꣔2�����/��q-�JϨ��M\|i��/BѼ�}���<�0�m��y^/ �o�o-V2f�w[i���T�[3Y�G떯>�f����vS΂iF��$�ȋ��|�A���&��� ,8�X��%�~�
K@c���~
�s�^Á��5uZxc�8E�4�ڵ���� ���|\�ܸIT�K��WX��ʌ}",:�`Sk�خ�^ѱ*rFC=�W1wT��7���;&\'f��R"�H�u�Ό��+��,�uzc%��u�8Rϣˠd^Gx}�����e:I��U�����f�Fn ��9Sݭ&�6�����n��V�����r�O��,����ShcC�,�8�m���kn�V���n{D����s�;pG]vԡ6K"q.q��l�:�.o:[��>���ﾪ����=M�v��'�Px������&.�w���+i�c��Xk~r�(,�^kMu}��q~$�A�r:LD.�� !3[���H��=��qWyW^��V2��y��Ӹ�´���^#��Q>�%��>�����kÌFbOÐ2-:l(�����K0�3[�f������q�G�|� �W�`�\Q�t���Ɋ�^o�ս^�e:���W��erB=罹ן����P@�1@X>f���	,?	����M��m��TdeoMK��9ɸn)��:�5��5�w>�!r��L�ϽP�K��J�p&��]�^X�\U�%q�q�V_�l����g�
h��!ա32���zba��[���7�W3G�Y�1;M�rj���N�
 :Ʉ�:Òf�yٹ�κ�6�l[��璵o2��`�f��3y��?PZ�K�у@�ˋA@u0�Q1����8�lc��d��{^r8J�ʉ�uC]��W��p�kx�VH���F��w����F*��8�rT�*��/ ~tg�ᙘ�[SmJbC]��97����=׶�F��٬A�#2�U8�^�4a�K̀:�"�+�T� ˌ��7W%�e� �>Uv˚`���8&:�5K�w;�C�8�$䁚�Ԣ�G��舏�E����ʚ�#G�TF+�38&Ls�ȿ�"*P�j�v��x���\3<�{i�ʂmgq}$���%�7vf�s*��NfZ��S��Y�5�5U�����c�Y�lx��e�#<�4��	zB����r�l�᳓*�|ǋrŽ��9궅zK��Ȑ�b;E��bkr�?Q�ڞ�x���\+�	⫻V���#�'�
��\���os�.���$M�Q��������`�N	!�����p�&��e酼h�"\��d��9�4��C/���D�8m�������×�1�CW�M��>|����_-O��4��w4Շ')�Z�}UV+5p��cv�^�W[�C�&�W`�<.���re���C�������s7��%�R���Γ
c>wM��]/dE����f��>�o��m/Cv<'����{���j���٘����^�'5EC��N^�?,=*d����0+��	P�ʶGG#�1�S�f��C"�J�8�l9�
����@�4����E��K�Y*�v�Uǅϵw;$w)���ᨚ�����G�k���"���0���-��+�Vݲu!uhc�(��+��)��*I�>ӹ�κ�^�.��nnT�#�dKXv��C�l��o^M����gd9�����U5���}Ƨ�}UU���O��i����#�P�����/�T=�}�t�*���P�p�&c:۱9��"�bڂĬ�o�a���VXΑr&t	��UL�JF$Ȏc�!hؾge�Sv،�-5w�� �bJ���*z�t�LV�u|�|X�smq� T�@�jb��ʼ2�����=�+��W��xOw-���f�K��2D� �6��?:�pB�p t�D��/�{M(x��7C��d)]�{������rwR���&� �s:��ɚ�L������ >��S6�nm����b1�VC����ʇ1�����H�9�ȓ	ә�Ԋ��0D�F
���Az{�ڥO��[ءt�o����m|t���/��oA��[�KGs��C��f4��3�nī�T���I%m8]�T@��k�X���/<5�D�|i��ܯh����k�`Z1�[�i�ڜޚ��1S�#5b�� #Ƽ"�u��??�,'.�p~�\j�@��Z\�ɭkUQ�7�??�g��t|\T��ڤw���z�������n�*��\�bm�&�i�Ր:r�Tfp�9{Wb�]��^��VR�*R^@a��N��ru|Y�(n���|�w��(��!f���ƽq��^ˮ�j�-�7t��9j�ԝ�R��B�˕�D��z�\��8��]��wBm�/�(ͰF�FzSS��BW�_}_C�|y4IS�g�;R&��D�2cP}^�|��E�j�[��i�b�7���P�[��}I[��L6����B��X����F35��tv�sqL���}ϯ�e��K;����K�b��ORi<^�̾,V��P���tO!�9��䩅.�0��M:�N�Ԫ��*{����of+n�ѯS8	<�-P�u�M!:A�!D��(�v�g:�����x�Z���Gj���h�2�mc"'kf��J�!|N��PT��"jx����>4��;{@��Z��[rØ%S��3���{+½���� qѶ�P �꞉���/���(�Jj��~���Qyq�}5/���q.�t�Cg��z�+����BbZ�3�p34Ӷ����:�)��yd�z�����n�$�θ�EJ����18m��un����:�g��B��yj�烈�H��5��a_#����9.D���ϓ�r(M�_T��(�z6�@�7}UD��~_PzT���������*y�#�fg�c)[=�����xH^Ko~���ˡ7{d`l�[��
%�w�!�Y�^�g�1�/.$Z;W���� �~ٍ��\������v�6�YY�oI���,�X���q��r�N���L�����g,��|$��C�C2/(��opub:cvv�r\V����悔�%61��Z��_n���k����a��w�Y_<���s��DU���F}�ݗ�z�Egڏ���v�[s�i�6(���t�N�P�0���~����>�K";Z�'�7}��7�g�������s35&�B��	��v�j�>�����;�wQ|b$g���O����}���U�P�����T�b�7�=?��,�d4x�s	K&�M1kv:���.���Z�FE��p���~�6�����@K�Qk�g*M��p٢'1��n���p�v�Ϝt��y�.�+Bf�8��8���j	�i��~��ؙ��}�ʏ>���2��p7FoL�s��m��3&��o���-��g��N�;�S�eRXˆ;\�k�'��F�T����-0�{��0"*��Vd���D�	/(cQ�����n����a�y���i��0�[�2�ܪ lY��&q��.G-�DU�MQZ&u1rX�'o�-Qº��J;s!w��VQ�n��Q�w��G+H*h�c�w:R����7b��70���ǯ���M%Y�v��JD�N�zݵ���c�w�I\4��ϴ�Nnq�qﾏ����d>�q;��	K=�	K��%[���4�[s���KP�ˋ��P�Py�	)~�@�%w;�Y�}��&��K�K"̒���$����̍��$������;�C�F)k�|{���%��sy�sf�a�k��'��q�#x�����W�Ak�K��؞w�JM^�{S�P���i8�Fm4�ʸa�;�2��;t~�/��_�.���@u\`�O'�bV�7O�O6�4V8TSq��B�ƸȨj�y�ȫ�LV�aV�R���ﯺ+�VTe�[η��tm�6�:���0�C�1K�£��������~�^�ʵ��3�e�W��IƼa��{sD/Mڞ��P"��*֚F�����a��S��U��8q@���\uW(�����])YQ��pe^�}��#�t^��i�x��A-��n�8t�W�+�:Q�q��Т��׊ݕ2�W��eQ=�D%����%[1V�c��x�&�Q�˕�I��'�w����<4��@d�a�|9a��)'�r��ȦYS��j>�s�p�F�ʝ�s�nƢ�֚Qf.�7��R�"m�p�I����"�-�{O��x���e�X���B��[��o���3���NM��TƝ�4N�c)�WƲ\�m�mLt�D24.�gc�Z���*r�w֍��E��܏��%9��7����;[�I��@����U�������SN�K�u⬊�ؗ�m<e�Ye��:uf���P�2�V3�̪�Fn�oB���a���9C]}Ы�86��5��8n�;R��߶�8f���Y�.�a����JrR�.�a�Ǝ&��.�LҾ��s"���c�"qV�Z�h�o.�fV�N��po)\�*��]#<rk�)9�N��{�N*�W��KY���Ssq��M�X�:�F`�p�2#xí�n$�Ø�EBۮ��nI�k��͜�WYF�n)[�Xk'*��f͆��w��v�����Φ\+�^�h�g ��H���@�tw�X�ze�M����ڦs�%"��uA��&]n���ڡ���]vǥ�P�R�����t��<1&�"�5F��\܈,Ř�ք܌��*��"�*�/�^�����$g1Sc���yel��6������I��|��9"eC>�0��4-� 4L�g{pF�,NO0��t�Gvĳw8�IApZ�$�5P�e`1�ќ�9@gƧfW8h�t�_KfZ֤W��c��@��R3;�cz��,jm:-��ծ�VB�Sk6u@�{����9��uf1a�������V:w3l�C�������4���r�u�z��,wӶ�[mb��n��fwqy��Q�}��������h�'V`Ŋ�5t��6r� �����1ڊvqt�)}�WwH	B��l�)r��������s�V�*<Rܾ��q������U*���%��N�A1N�6�-࡝�r\�]�M��:�׎���e���ԱR�5��
B>�c��6�p�
R�O�j��΁�6�l��Ycq��:�����x���<V>*��v�q�)�kE�3֭[����ж����y�Eu:�"�2IF
��D����xL��a9���\����yݐA�a��ai�b�y�˭X!�2��ỽ�9s4�3���w�*7	��Í�u��m��+�*�'9�^Q�f�*�dp��o�A����駥�f�̤v�X��|��5�E����X��XꆝG��Z;�<�ՙj��s�c&ܴt0�)����������*���%��F_-Zc"��%r��9e��b��}Z�;N�b�ۗ8�'�tM�腢K(^䦀5E���5P��+aR�_e� L���	I�e�S���ɘf'�9
Ӯ��6Mti�h�C����߾�=�w�������$i�II!�f��	΄�0RFJ1��� ��`1hҙ3(����H%4X�1��H�<딲l	�u
%�fg"wq4�湘��7#%�F����uD �Rnw:���n�%�t�����&9�e%!�wv��wu�ǝ�1;9��&#+�s�)������ˠr�c�\��2Jw"��.�F (M�ww)"�"D]�d�d� a,�y�<�K��˱��v����]�)�șۃ����/7�ҢL\.���&1d������%'��^9@�U@|M> @��[8�j*��%�q�
�v���R�x��$%���2l�q���+%c��v�iViy�s���vU�&Xuڭ�O�к������׏��>u9�u(�
�]��u��kk��v�q:��pP��5��1�nY{�ܑjEs�U�����O���gmh��vc��9yq����������Yk ���に��Byx��i�¬�z.y�(�5�1��k�M�<���~�H�4;��I�Dk��,眶�cq��x�q\o��̲�K�wEQ�y��IsʲN"G����|�\��r������:3���'d������/�h��Wҟ���+�~^�>��9�j��ɝ�t[v�2��y�9n��ca�誠�G|�ФC򼸽����k�������m�ь�M���K}-�S�����
�?p��m�+]U��{=���C9��j��u�\�5������˔����J��E��t���i��7�~��b��k~I+9�MƻB�\\k��opΆ�,r�@c��$a�e��CˢX�t	ǵ/��:������i�#l�wdN�
B_sꏩ����f��Kv��!�ZU �Q�7��6jÆ5�O�BK�[˪*Ұ�&1��8�٬c���;��յ��S�	�g��;��ěb�VISz�G���}�Df��6P�D����gm�ϩc����6�;��Z���ډ�Q��Lr����^��T�L}���&����s͟�9�{��\�n{pۼ��G)U::�Y`�Y�*Ḇjw�w�s%�Nb5oM,�1��D� ��e�Q��:R@,���F�{����f���ݖk\^�Y�q�»V��&v 0w���t���8��OWcy��w}�eu��[p.ěɫ��v��6aj�T�T�k�S��1�V������ٷ�=G��]u{��f��}�ϊo@�����4dk��K�
*"�Jt�z�����fn{�s`y�N�W�^?S��mc�DG2��p��R17���s�ӽ�{cw�M8W��Л�0�����!�a�~��쥃m���ALP��L��k�%:zM�j�ۊ/C�[-�Ѣ埗܆ӡ�J��E�*��O���9l�xk}��!{�uxa')�83f��E��}4+�3�r�ʶum�o!ʺ�c�;'�^�$�+=���|V*jŧR�[�>a�ד��E�b\<���p��ì�T������Uw][Z�}sOpb7t/B���I)�������?y��'����|��q*�n7�%�~�P)�e|�}1�j�Wu�n'�B19o�U�ڋ��&�3������.��UAB���uNۦԌ"kŏ�{][�r�E��ys���w[�p�CH��/�݇�yM$d��aƉ�?N��]�Y�5��q��rNk�7��v��Qv�P��Q����IN�z���~�m��2�]�G�YY�����3�����\�B�;��q�[q;�^���dj���b/>��d�;�6�aԬN�n�����f� ��Z����Cn�?s̫��9Q6���$3i���5^�ھ�p�g���r�3ʷ3��O����F=�e���Q�5���yv���]�&�����z�w�ϝ��p�ŭ���9�Hx��M���<���(�U��wn�}#Q�U�C�Q�*o>qt{�����0c��z��E�ay��F���z\X�<H�iR�;�0�["6� �}���564(Z�O$hpu�uI�-��
ƙB���WF��s���+%l��l�n�
��t����WZi�ɛ����\x͜�%1;���N�U}��US/}/{R�d^o|��w��Fm��UY�˕u��HtKv�����v�ț�}֡��=��k��o�L��N>x�c�As*�yUw�5t{!�XWc�[��7v��mB�x�ki�9��>�	tU�|3Q7��e�.{����Fk��5S��*���^�)�E�+�O�}�"�3�Lv��K��D�������h%����.�E�t79�-������.��d�*l��$x]�2\gٴ#G�)���B���B}�*�,�3&$�FcR���w�������������´О��.�e�EW��\ё+pȊ��Y���.Bř������р���p��t���R�N��6	ͥճ:t�f�[4b�cM�1�9vÌv�E|�\T5l�K�:k�3z�M�s�O/F��UU?�e}�wb�I?,p���]�!Xc\dT5`q�+j��S��3�}(<C�zc��h��4)I�s�&�m�7�g��W��XϯFZկI%���^�u^�wU�Dnk�Ą�}Εw8w��fTngOJ�-�q�{�R�&��9E��ZN��Pf���9/����!R>������:�5�;sv���Y5̯着��&�6�jq\̿E<��{�m\o3��-p��(m�Zc�X1����
�ۭ,I��8�3�_a�y9��2Ϋꧩ8�l!�^�#��΄�[�[J�'}�Mw�T����p��ϺQ��)�<�
f)�Ȝ����(�i��v�F��f�[��A�D�#u��P��أw������_ZK��cmN����e;�o;�ݪ];3֨��/)�^������Wun��u�f�c�\c��\�dC�����L��N.�	ь���S]ׇz�|��*oqо?R���;����	��6�駶�9\h�U �wxs�3I�F�u��ٞ���N�4�iT��I�놶���9h#;��9ntˇ�$��z�ʧ��Th6/��3�.{rN"G����3����<�ciҎ6*}�8k�VŏO�F��%XO��,~�L���FC�&Ҕm�O��x�M�M�ŖAO���La�.V��y�>��,jG`�����k�ќg����Bu�"�=�Y��dk�zk2qnV>F\�Jp��#�/�n�v�J��K;>i�=���!]�2��r`�w���a�vJS+��#7�䔢h~��>���Zx���s{������쟞1���|��1�.�LO=��Rי���b�6K���e��ِ�&&��[�wZ��FëtB�:ew��n��o$ļ�K^]1<�_d����{�&Ìw�E|��?*�Q�N5����0���� ���fWeg��Qř����4Vs�)�֤�箁����+&�e{驈���j��Y���~����J��-���'�"8S��W�X��^�X����^�E𾎆g:��ƻ:��UYn�^!���U���[��;�����O����/m�f����X�s� ǂ�b�U\:tp�\�QSP�7��Rٴ�;�O{#_a��e���쳓�������֮��&#sOm�ޫ����3�p����sYݍeu��[8e�]kzf&�E:<�����E�J��������ޯ��m�=B��-^�E�%�䥏[!�N�٤�̷�n�H^��S��j�)QO"h��j9�n���X'��u^G/X~]�r���q�;���b�,��R��a�Мp�z����@DGS�v�z��ɭ�9S��w3zTz.f�P���Úr3����#^==��;"��g��ʗ�#Q���(�~����S�M��q��n��V�fa^m��f��[�A�ǧ4{�S�pU cy�H\�,���eo_C��1��'�4��,n�w+�T��i���*p/�`Y7oj'v�<z�I쌮6��o�qy�8al�z.Y_o`�>�����[߆��*OW�7�q)�-���U�܈ovL<cM2���5�[3W���W5��^���hƸ�qQ:ګ��m_h\�J]�yfI����3M�Z�̧���m���H.2���DƉO���˔�/�#���}.�c����iN�ӡ���b�VÔ��]��Q�Y��Kj�1׵�����Q9���r�+vi���!q�s.��ُ��m��/��]�p� �޼�L��>l��
���N��u��q�_k�d�19��S��&&��*S����m�<}��^�˞lO�)c2	IJw����
I�fQ#��ŢŻ������s6��Z%�Zګ�6��%��Q�sH�a1����e�ڽ��VSW1-�OU�v�m��klj���`Z��̭�zD��Ve��ћ��B��n8��5AN�W�_}�^�����0�v�FY����\�â�4�Ls̫}3p^��}�`\����y@�N�t�vN�<�սT�n|��6�Z��+2I��:�Hqy���Iy(���5u���8�D_>v����������G�É��S�C7�N>2q�^S�[;��$o���W����}J��}Oӭ����|P���.�WU�m�S��KQƲ���q
�F�A�P�����U2�,��(�⣦���y�)����r��!6��=���nq��>v�e�o"\����;dqr����H7�wxᬸ�Oͧ�g+�(��S�p�΅[���QC8�cs�Z[,����mㅦ!�?6[��r��0�����}��4�i��O�{�~�]I�e�o�D�A7�w�;M�9R8܇սt���J&��<�~�H�$�
y�Њ��4�I�j��ߜ�2�7�Khy�:�r�=�a�}�����	�艜�;���Z�1�D�p�h�;�C��&;�ڨ��hZ��G���*)4B�0;���՛OV����ŬL�W:�I��<ŔOj���ƹEהE��� �q���"���]\�{�����������I+�N쓣�Hu��]C�C��'�Q�������C��\�4��;i�[@��ta�Ǫ�{}yF_�S":W�/Y�o[����t�NѶ���B��&4��F#�r�q��ȨN.*�����vc��ūq��	�X~5��N����oRF��
�n5�B�\dW;��-/hN+����}�n��va���oVVY�q��-p�E������Q�:#q�5����{������Oݦ�}���;f��)�9ng���V��Ba�9��҃�;��Y~���\y����F���w�ؠ}eꛮm�$2�uoSI%ʨ�Joy��z5�����z\�ye��ίl��f����x��*���r}'�r��M�ȧ{������3ݰ�Hձc5��3a*gn[n�mi@���WvK��\�c���=�|�`ՠm�����MF���=I$&���^�T�^%i}��n�R8�;�	˚�\�ʆV[K�8r���fO,�0$��g^V��ux���n%��[7�)�F�<�s�:!.��zF ��*��VmohG�nK)�Q]̵���M9��Pva���&ؗ�u#��N���O���Ͻ^i���3�!i���]��Y}��~՞�Nz��j)��v9<�w��Xr�ܙS�>[A#�ʐCq'�ᬷ�H�Z �Á���k7��}X��O�E���|��9tUغ��2�˞�4�#�)u�JEm*B���Ĝ�31��f��9�L�1r�|��B6�;Ϫ�/���͵j�S��2���mܻչ�Ɉy㮼ߓ��<��
�'���XԀ�\��}}�ed�y�<�=�M+�[�nJ�m�V�L�`���9w��W��,�6�A�n�s�8�w�	s�������=q�]��D
��/|�9�R)��2�$��'tΚr�'����׊�F�B�sG��k=3�o�	��n��X'a�FU������ؒ�4����K��\�f�߱�$Y�I��r�$���	����(k������ ���3��z�p�~�|E�*����ȁ�7�0j���"��`���u8�/���h-$_�Ӓ��S��@3�nvx�f��`{w��U�X�}-��5����x"�v;^l���̱�|x��I�w!�9%|s��ۻW\$�l����G�h�E
�fj�3��Q e��^��k#�F�J<e��u|��M�@�B�����{u��m����֧v���&�F����'
{s8\��s��V�M��̫b@�k6�H�&�]�H�ֶ��AI}oh�N����Ӌ��Tq�Z��+p��x:4�o�Q!Q��ROYC*�X�ӹ�sN�[��W+�1f���|~��yp'Jo�"f�X&����@��1W:��m���]���70�r0T,Y�9eI�Z��{W]>۫,V�]�3J�m\��u\+��;�9f�����L�{�bKYW+���Jٕ�Jhcy���-czf���J�m;7��$gu�jo\*lҲ��MQqu%�ʜ�~UB�# 5�*�ۮ -���9��O�o=����ImiT�/��ʈ�r_<�5r�X�vS-�6;�uՖ%9�y(�z���2�1��ڼ�ۡkR�U�v-�*��#�2c��33���兝��]0X�.�.�!-RI��3/w��g-�2�ĮU��ϲSR�e��29]ƛEA���sy��!s�������U�J@����TC)"��X:łA���(�ҺJ̳Ғ��''�X��;�N�~ __^P�c]mZmbZ�OT9��N-g[=%����[��B_n�:�H��2���9gL��H*�=i�Rl�"*��]�i<�]H:��99����=֖j��wj��v�ht�--*�a-���:�цV�֭M�CF�]-�*��&��^��L�8��\l�B;�Z���J.�]yܖ�T]:�BM���i8"31;�ӝ]��kel�� 4�ֆsI�@m1���FNtn�p�J�΋��귅u�i	5��F�.9ʨd���
7)��'U����qp!{H��,;ŗM7iV^�Ѫ�0r��o�̞.�l�����i��76���)��1�d������"��S9z"fʓ�� �\�z^v!P+�n� g[�w��%O�`��p> ��%�x[+]��B��[GU��$4:�Z�QP�R��Rpf��i�n�r�YvTQ4UcVGYK��y{��MeN��X{��Jq��	V;���3f����:���
� �� ��F�]��p,RO��LQ��&�R@V���hމ5ީ�Q���}ѧ&@p�G��A+�V��*�g"W]<5R�r&���wZ��
`����!+�d�DEm�
�
]˶�c۵���ٕc�
5�64e,-��t"Onoem�e7�ouR�fK�b���.���(D�E*QZ*�Xv5�.c���'��4�KZ��L=�H樜E���)b����]R��I��w,Im�KN�N�R? a2K��qtWd�$;��FH2n���8lQ�֒4t��'t�t���;��ww.$D.��%��wG#��Ne��ݛ���w�nx�s�t��r��<o	vac�K�u��죗;��9���#��N���1���Qcp�u����;�y�+ˇn�uݓrӺ��s�����q���Q�w�y��f\��r�fw]G.gu���M˗	:b�G(.sE8��.w9��,\�wiwN���s�ip�Q�î��Mw]�n�WCw�nn����]!u�!9N�]�p�w]�]�Wdn�\�v.�3Cf����T�4��S6�>��ݜ@�9.����F�h���}�lEPr�Gx
kf^Fg���Z���9f��4?}�|Wj��q��t�~����-q���q���w�o�n����1������MM D���ހ����^�q'�����7��yYm���8��P5�F��}*�@�/����{q���t�|�=]�7����Ʋ�.��'��0�����C3�F��הk���*�ճ��RDg���Zip�	�0\�V�ץf<�=X�vc�B<̧4y{���pO^d�w� ����Ak'C:���^��#�釮�*;F��:FGIzu���gk@����sRj�5E_cJ��LCi텍��atʨ{��ZV뷗��������ն�Q��?o�Q�3K�a��Ƌ���a���r6R�y�L=�bw��VTL��u�*�n|�쟞1�)�'A��lF�c������5"�՟S�[�Z�em}}��ҿ�޷�fI��ƚ�������� V���Is:�7�n������9b�;I.b���(�w�u�a�=��u�p �*��訤bs�q;�f��n�wO,���!vE��ۙ�K�[2j�Ͳ^˦��+\�Y׹WP�η;������£JN��NM���_}M`�I�uʤ�F�~��m�-�[�Ju}�\��\U�Q�6��S���'��%�3�� �Z���צ,�ϳXO�L��m]����ͧ	�M�>�.+\\Ts�G�����ٗI����w�x��0��eS�����4~X�Sn'69�q�Q��q���b��Vf��r��Jt۬ŷ�.�Ϸ���p�Ų��3y�U�Ϧr�}��a��햊[�!���9�o��ќ����k�����c���6N���t�>D�j��{;��3"���=�2/�;�U�-S�P�'���MJ�����$n��د)o� �̠����\�>��C{k�wp�7���of�(a6�3y�'��5�Ձ�1�
�g�*�F����Dߧ��N�R)?�q__9N�o��=B�[X��t|��
3�k/�4z������Z�cS�f�nS͌H�N=a0bO��z��XyWHd��\�����7hP\�aꢾ��oD����M�w2,j�5�U�V]�:���n�w"y+b��(
7�e��m�
���7{�P=�ʑ�H]3�$F$2g�F�i���֕荒�pK�7wᬿ������Y��d��Uc�W��6'��\S�d���P�~���sC���n8Y�<�-�X��=r�Ʃ�+:�[=��ia7=>{�	B���4��-���%�D�}��澨Sq?^:��T�ut�b�C=W��O���IV��EkJm�,Q��}{N>���+�a�ln�|�ʿg��N�؏(RϨ�ח������������]#E8m�q-��bԫ�2+��Ԡ�L�����]��T���2���qY5UN����\h�N[���2*���=L�<�*y���o=���V�8(8�o2�<��4�W}*-��hV��Ae|�8cn��4�
$��S?[Zs͟�����o�oOW��P�k�cW:��Y!�9Pz�(�LoL�Z��}>��~�v��cFr�s=11h�3����s����4Q��B��H+��^x;�+N���nޓF��l�J4�[�,���Yj��f�I����G\qR��!�Iƻs0��f��F��bt�����9�U�FaސL���m��n������2`G��N�m�5Y�J�u��wO�ӷ�]��EߔMM��b�а�Vynm�]��v⶜n�Δ�ʩ8���n���{Y�LOy�w�Jw}�↍.�a�01�K�:�8�M�ȧ{����EosCxf���a-~���W֭��2�d�ϯ�7X����W����`�:uVM��y���=8\��P�1N9�&/���ުi�N�^�
��z�H���P��z��9�dʳ�7%Ý'�W��.e��a��Т~�sA�~�#P���'�"����=&U�=�d�LkW��r��K���3�9�����M��R�b�_r����������u]��1٧��iH�ِ�|�iC:��He{�V{3ו.�F�.h�Z��P�u�bp?�k���'����]�����1��
���L���V'p��
I�[��b
i�n�"C&��Ox��+,	<U�����yeߺ���`Q��O!�5��j��(�6������	AB,:�0��b�5y8��wL�:��"�|�]�¤)Cr����J�r,�g
|�\n�h���˜��z�b��
�A�Y��1:��	.u�	���ž����)����N湆�iv�ZGJ�=���{M�^�I2�����!ৌ���Jz(qw�:+�g��Ȩe�r_F��ه襎�b��6�4�h�<;�� W'v�ɸUmD�b�k�%��TN�3��S�&���X+q>X�^ø��^Puo�nC���χ��!�5��8%��Zl�o\.ކ+gkS�Û,�wT�y=x��k��n���R���/5��-t�X����WXi)��/�Nu>qp������ʵB�]r�����G{�"j��?W��PJ�r��ӝ^�T�[�ueN\��$�R7��7-�<v^_}�+ٍo�%2�N���wF;L�>y��s(y�i�2ar�8���J����OH����j_<���`5E}�m}w�u�b����˰|)����х��R�Q�@V󩶜�8��q�kC	VV!��耔��.��.�	��zf�����@X�.��O9r	(\*'�\0e<�㼒����r2��!QֺM#i�������ݾF\��d�'��Z�r�K#.�M��Z��[^�7��q��4 Ջ�.��ꜧp������~��ˎx�f��y��-�F��Wܪ�m�}&���ܽt�;�0�w�?OelJ]�����=�9��^h4��}h~X&���	A��Lh��'V����}��M+�]��Ux������$_͋��|g�Łe~�x�jF?���ފ�v�]򹧝8�~[#Z;]��:sFؾ���:��2.r�p��t���S죋#b\��ި!��t��1v3��|��0۩�N�z�f�{�i��v��pudՙ<���UT��f�W�r4ac�M�����=N�yX�Vzo�\�-�	�VF��}�5�e�W��>��[�3b��wD��.u�TH�RI,I��8��cݱO'1=����:�l����Lq1T�{��3�wbX�V��b&c؂�ۜ�\�γFL3G7q�s]���b«i�x|@����������%�ۀMR����L;���I�p���}��J��{j5բ����J�k�����l����U:�)�Й\�����kN��mo_-B�8��3���xMΫ���䧨<o�`�j#��]�]�ty������q���ԍ�N��(}�:;^^�,P�-g7��>�Ό�F��_���)�jx���ѝ���X�~��/r����Oۻ�*4������/��I��)�ۅY��X�����5�̣o�a莉<�[p᫋�E��RJʤ�[6�������{p'9����k�{}�-�K�ś�@/Q���PH�P�vU���5��8Za�ו_���/6J����:S��*J_4�(r����~	w\J���>�p�7b�F�*�v�����[�fܪ�#��<�|"�iJ7k����b�zo�o.�}'7��|��3$�li�X*�#�+�Lh���~�Z��'�=�}���xÇӓu܂B|�ķ�ܕ+�ȨN����::f&PY�H�}{��y�m��S�W̆�Cf�N�@c�ϸec�aܨbS�h��&kij,�4;q,h�I� x�#rf;~�3�}�=kU�Q!��Wh�+��fے_n��A�^<�8��j�nqN�GH�o�4��vq��N��v\�L��HZs�����.�1��3�3	q��$��1��Nt5lv�\�9y}YK;���MOc��+���?F,��x�F��
�n5�!X�Z:*�݉|=ɽԒVM�!�=)���~��6���d���aEGE&v�<��:�W�9����+Ng�����o�/1�ӧ�k'Y7J�c�Wn��k<��oq�n9co�W�R�y��#����7��z�s#�FO�ofא�|��U�/���n��F����m���[���8S�]�yhArby�=��?����]<�J�}��v��1�mu���"b��;J��&�2H�5���1и�>8T_.n�oCՌ,��B4S�d��S�;�$��������vE(�pw�Ɉ��n���!��ur�f�:>r���732�ԯ��tL�eQ���44*A�I�+��n*�� 	a �R�B[��!��v�2V_ؼ������Tb��{z�����Ǻܦ�S�ٱu�ߦc�%m.��[X��{��mE6���S_V���z�Z�xU,�0�'���ZJ�ܬ�Iǅ���CkD�![��.�֝ڑ]^R�֧j��N�6���հ��z*�?y\A�*�l�{���~�ɛCjq��m=����)+m�]�k��m��R���f!}ʄh�J2i����n����.�=�u�_-w�m+�z����i�K�
�#���K��wx��"M�gU0c\D��r���B?ri\����-I���ҧ�:*9�j42NoR(Y�Ph��cG�/U[�c��.tS}.����3�h�q/��8;y'j�p����וs�yӹ{b�e�>=z��Z�.������٧�cR�s�q�M[
�����5ه襎�Z��&2VF�Ε�9ڎ�9w�9��\:/�q��a�pɯm��\�?[|k<ڭ�,�S'#��<	ٚ�q����}�O���x鍼u�;ʻ�}3�~�cm8��:�{ul#����p�^���[7�'���O�"5�?�׋>�\�^?$���LBU�-��a�S�d�̐�3^�~�=�m@��6�u.�%ǃh0�V
[F*�;,^�j(+j�%���3���n�^��dO��Hd�LM���!��h����-*�s`�G;/FA�%�.\Gp	�=�]��]�k7�ȼ�Q��#V����:ΣW:}=S���|�����bʠV�R�A8wmw��v���v:^Q���Vz��=J�b�2�B����n]l�����X]5�j)��������`��g�*�9����Գ������>m�P.o)}W�m��^[/�Ut|f��G��2���iuI0�,��v����
��bo.#\5��8ZbOe[}��atʝ��ǌX�i,J�s
9�nK�u�Ҹ)`0y|����8^��n�\��'��������VR}+���u��+��Z@�+*�K��U��ovLC�5����4�N\RQ$����LD�:���ھЏ&�3����̃_o%����6�����3)؏(R5By�}qwm���
�:(��x�j�sv�ݧ	�1n]��Mۓ�%q��+]�O��ԶQh��W��GF��Q��t(��^<�o��Pv��kz���N�e&� ���u.�G��$\D0,{U�#��b<��f9����T�x ����b@Ax,iD��mk�Ӕ��S;W��Gc0F�9��p��I|0G�㋃�-�����A����qՋ灩����z��(�<ݱ�/i�����l��@-NkN�82+)��Y� ����	��C/��跹;85m&�kwS��������0 r��'(JTW7��tC[C2�	��K������Ф��'B��J�8���ƶ�^�n��|����!J��՝2�H�]r0�b��6�2匏���T��ڏ�n+�JI]Ӧ+R��\U�8�.��*'�f�a�β�z�2>̫&����R�ݦ�A�Gf�_ r�A� �t.��Y� ��� c����<A�.�X)?�vQj���m����o�G��w�7B�=F�H�7]�.#���q�Q�c�}V֬��&X]m���p�$�V�ʥ�YϦ���4�)�˄����g�b�ƒ[�m+�g�LB�gr$�IL��Vk�o�odZژ�<ʶj.��Lmj޺勸pp�0�ޢ�JZ��p����4P�
�D�.���6�����1k�1,��+�����eU�[KB�w1�v,(���=��K�ۑ�1w#��]\-��o�쐬�2���I����{1&��[h���ј7���9XN���+�Eg�	�dy}"���C��}(����(��|��h�집��8,��[:ѵ���h)����J[�M
-�xWGiks�����í5]oY��^*�����V`5� ����H��˓/_Q���jqެu��<arʮB��6g��/�u��0Q㨘�é�3ٱ)eM�f�'+�9
E���5��(�:�M},!Hb��J�+�lЊ���W�k�QfQNTr��XfV0)�d��2�4��0� v�@.\��bO0
݁"H�5XZ3V-���=se�u�¶(����K�c�..��]ٹoYZє�l�eT�Q��-�aB�Ս��X�휲�p����l� \�2JE&��ʾ���Q#��R���e���%�+rt�en��8�ô%ԙ����@�������������@�B2e�u4���7�N�TlQ</5]���!+'p���T��Z!ך��LJ��6�%sU�p8�C��N���L�Ү�s0JéV��X�����nJ�9�րc-*!�5���͗u�F࡙���V�,�	�]�$�ݖs�NXBO�G�vo=��WefQUrIK�/V���Cor�X�����@��� ��j����Wx+�4�� Z�/D��M�Ԧ������Qݵ솝�����i�nZ�&;S\�;b�w4��_sM�*��)(�x��ܘgw�������T�u�d9�ܝ4�s:�.�����9r]��n�r9wn�r���N뻇]�\�r9;��rs������u��w]��wdS��t��.�9��:��s�]��(wN��]��G&BA��˸܍�u�ra]۔�����N]�G;�\�E�̤0W;�\�"4Hܺ��Bfs;�ܮ��n�3��渊fK��pܮ�t�9I�:wnS���9p��������ݻ���.nf.q��&��	����]�nhw]�r�:L�r�]ە�qΙ!�w5� �뻺3p5�bK��d�u'we$�;��4��f��I��f]ws��a��uӹ��"뻝s�uN��t��v��ۺ�)]˷sr������ߞ~��\�q�St9C���Qi�c��p�5Q��$��h�0Z^N�g���ɖmi��#��D��Bd�⎅��t�91����|ۍw\Tk����n��v�X�)K�ٺ��jw��Zc��f]8�Y_Fq�w3F!c�E�Uþ�g��T�ILk)�����)%n�x���!��[9��9O�+��sګ���m�6�:�Q��n�A[��I+m4�z��b�\��g�ڥ�1���_e�W�Kf�I��j�V��Ǽ�R��sAz׫�<k�.K�v�X���S�[�u�_fEFGm�!���=j��JOz��N*�<i�<���Ⱦ��UX�s��u>��Rk0@��&(Z���A�o.Qpo����z�F5����?q:�O<[T�"�v;D�֔������W��[�����o�Yͫ���J��	��UȒ1�Zb��]ΐK�47x�X�i����,��=��F�>{�WF�r�vs��F�s����������Cz�v���yfLQEV0�R�k|w��-ң�9ŵ�S�ř*��K$��֙.��wy�}�VWR��TJ�&t��"��B5�ie�����]l�m��bɛ(㥭Knq��x��t�[�e�ǆB��vIc��j=Z���{�y�ͮ�Hq��ksE*t"����F�/�����对l�/�Byb��9񑰪�s���w��tgrI��}fc�S�i��2�b^��T��JQS��_ҷ�=��U���n/j2���w.�,c2L6ƖK��*��uJ��ƈ�}C�p�Mn-�oTsqx`�O��Q}����\K}-�R��2*�D*c�W3R�����g���j��[7�9�Z}��K��'.���bqpݘ��6z�Γb�4��<2g1�N�s/�O(��+��%U�*-��J����G���2��FEoX�"'-�������6��j�Q�i�����ӹ����<5!��,�g�&��F*��y��`i&{j�-ҵ��۝)7T��i�<a�����C�.�ت�MM�ϧd�k�^nC'fnmƨ{z㪹ħ���^�ǥ	>��Ⱦ[V������壓�aS�su����e�4����ee&i��-Y�"���v0�}3gZVM��4Rg��L�zc[�o.+�q��V�>�}J�
` �H���Z�R��O3��w%IJ}���Ɯ5z0���Ϝˇ�JtlV*F���,�mɕ)r�ej��GRR/��n�wp/�I���m�w�7�c�Ⲙ��+��5HD�8��Q#t�S�1�q����
*�su�;o�)���@7r�<v2��'�W����t�>fS�|}����<,��v���5Xm�}'�F�qMv�K�6��2�0�Dy�$�Ϝ�a�P)h�F�&�{[mJ���r���%�{�[��{h-3*|��Tj�b�zK=Lu]�����r~������9��}�3L[s��JዖWܦ6dƦxtRDkݭ���NÜZ��^�=r�s�z�!��0�?2]UA\_���8�9O����?V9�>���bw+��B1ɥq-��bԖ���PoI�q�3��IC<�AW�.��"���ח^t��fd���i�`��=37�53w�z+�nu�*���/�镹Y�Q�f�SK�5A��L�kw�j�L%m�Z�\ g5�ʀ�WӶ�ۨ.� �P�0����m���ʛg~��^����xy9���(�7�n�F0�b��1����j��."'�h�V��P���B�5:q�WkKl��>��> ]�fۼ����8�«E2��ʲ2�I����3�����kRk���bK���Wf�����[��7z�W�Ã[*�&o/��z�k�Fډ��u�\a0�g�'W�ZL�r�B��w��t�M�����輍�}k\s���x�Jw�o�n��#i�K���N�����b�9�uT�Aj��[7���O�5�vŅ�B����kw�9��Kg`��k�Ε�k�#�:��:�������x�=G�v��U+��i�.�����y+d�����\b�>1�:��щ;��&z���S7��B[]��[T��zm�X�wF:
mY|b�r���#hB��U�ŭI�Rp���r�\&��tB�㋰+=3�6�E�(�@2��|	���YZkJuY��� q7�ᬸ�p��������T�jeU����\�;$���;�)`���<k�5�iy�͖�yA��[}�����o�3EsM�\�H�V��w2� ,�{'X7�P��>-u��7!�Q�&�
�Hx�)殰�ڴV��c�I&9�es�bܥO�[��V8Îf]i1v�9Zs?�l@�f��o�˔�y�|ۼq��q���-8==�ȋ̓�m��Mgv�~����2�T�0bVlhK���o���� D�x��"|
߸=��#���[&*_5��Q�:���+j/�#ɥ�|���̈�^���f��43$�{[�
�#R��h����R�˔�ܻb�蛪�[������r��X/�ۣ	��l[���>nܘ��+�*V:�yL\F|�k̻5{�p2UU7�Y�]U���m�>F�o��}=~Qzz���]�6){�u87�RyGgQY���c�E���a�q�Yx�*Ο���nТI�nM��?S�1Kެ��j�z�-p�[(hs/���m��l\��{���{��c|뻥b���m��4g*�Ζ���:V�O{}'1��vh��3�O�K��]��a�s�(56�/7\Uy\�km^�����I����z�7�����V�r�ݸ	e�������~�F�ś��'��a)J�C�����_��=l�}��]�O��&����e]\a�[��>���޺��s��B��!��4[�����Z�'�s.�h�w*���9���:�gc�A9y��$Wd�W��sRb��9:8�1bGw��`QQ���6�>�y����WY�����S�,x�}ƭ�n���l9�B��8\c)������I���ƫ9�a���f��R�3xc�v�N�Q93��Ďf�p��I_��pլp��i��S�jZ���u)�8M����;%�?PH��pU�@�n��me�mR������iִ��lT�ԆH�h�>rʢ$��*ˋk���\���^��0�}�O}|�c�L�Zd�r��O����XN;��#^��$n�-�S�fCI밚PΤ�̓�li�K���?uJ�1�����/��a�btӮח���з�5K}-�R��L��
���l�	�!I5��@a��q4>��TivV'���K�䜻�������خ������(�b�t�z%q��A�e��V+��x�䑣+��`S3�-�\AD���N�eN4k�
`tP���Y���Ɛ�r�7�'M���^�27���p�;����S�Jam����GsZj
����P8�p}�&W�5ۮ�oz�A����`f�Y�&)B��;�ZU�ٮ`�ޛH���7m�9�������N��uu�)JS�nJ�U�c���kَ��~�sϚ+�l�+�=ﻝ���ƛ�V���Ls���o�6��9�ռ1K'#�OL����q����'�i�e$Ĝjx����N��s�T�%F����[}[�P�s�Z6������+]�Ur�	�n��k�0��m�7��fXelNg��"�����B�����=F�@���So�)���{�4B�n*�(lֻirD�����;����N��(]��ʎ�\�c��]�3\��/v5�f
e��fG;��p��@�h�:]S�v���XvbZ��|�Zq;�cq8MF}=��q*0���ڳ&}g�V�zЍ�2�7�|��{#.�M���mㅥ�-�u��Ӷ�ܨo����n<f �q��p�忨bw�쿹c]��4ŷ8i�������^a��6q���2���C(v���H:���S���oL� :�-��`Y�#oC���Z��������=P"�Pu���c#�bF��;rcy�L�Q��nH�cǁ�W���Q��8�)�Z�Y�'�&�V�Y�+ ��w̶�M|�J��������}uҜrۙyK�	���M��z�6�˽[��ɈxƘd�W��6#cܭ֙B��>��PX�����i\K}.ص7Km�Z��e)zi�(�X�L�C>�G�������]�G����%κ�L�N�����a�����ֆ�%7	ۓ
���/�N���(�I��e8�<��J'9�R} ����4Vs�1	��p�Y�q�_5l+�K���"�2�gÓ���۶��Z"�]Uv_�4ھ�yk�E�N?��:�	}3���N�1�N�>uqʽ�WiZ7����Y�O��9�e��;ʸ!�.�".�F��Kfo�9�_n�<�8�DYz�����r|�]>�g-u��T�;ޥ*xs=�Kś0fo�z��':V�����s����$��j>��y:v��X�cԽR'�]���o���Oj�o*�y��T�r�Lb'ye7�]6�	��O��	y)�X2T��?{����Om�B)��*bZ�"չWV��\C�����p��u0�����w5�_�O vk�ۇr�.��5 Pˌ��л�gIF���TVO^���=Ԫ�Ƙa\Fq�v0�W9[R������y٫�M�E�?����Kn�͸���@!�TϪϜ����~�g^�ɷ��:�V�
/��\�}SOn!Vv.��0�Uz����h�ѿ*�^�Z��b��RJ�CwѮˌp���������t��o-nm���6:�;3��p'zjZF(w;)`!'��<k���C���Z�14�4�n�ɔ����O���:���#n�M�Q�{G�ҽJ�H�OCQY`.3�h�C���lƈ�'�/Z��F+˺���5ܳ�5�����ОΑ��]�YfKo!��D*�1؏�y�\]ڇ��g][�5�|���ɺ�A8O��K�bܻC"��&����S�w�o�g��!3�;��W�F#f������n1�0����p�g��M���c�m9iH';\���W[�bʌ�j���h���{ޡ��Ϫn@ǒ�!{�����k5)ak�33Cě�8%i��:�}'����:>PRHP�z_|f>�[.ya���a���<�3Q%V�0�Ts�da�tY���+y��R
�VAԻ�97��b[ʣ؝"�V��[k�˕ۏ������jG$���5��j�C�[|j������ꛞ����O8�ͣ=���Vo�pr�8�˚��$��A��A�Q��+OƑ�'g~���rv[z���b���v>�rM��<���֓�yV9��7�>Z���vT��g	�pB�5JϤ����_���^`wv���9J�.y���L^loV�Q�o追ڎ�&�_�gG���d�2K���tj��8+��k����|י��:l�!;�ݾu�b�1�R�B����<�NI�`;���j�$�kt訅2���>����T ����
�9�ϯ�׃�3~1|�w���r�m;�<�M%I�8 ^@�
E� �؂kҞD[�,u�[��%��ƀ���L&������RԪn�c<O�eK��Z!À���FHli�R�2�#�
�g�h�.��^��/GE\&3'r�{=2/[�a�F��{��;t	���l\A���32=��Ys�^�枠��"�\K��eͳ�9�ö�"���q�m Y�Ƕ&@����L3��J?��t���A[�IS$z����i�n�iA�Z���8�ĵ(>]jS��K��2�0���.ջ]�#��+a�V��{F[>1�L0/V�#
��O=)���ˆ��Vm���:ŵ��]�Xս:xDI���JLa�&���#��(x�z�iԬ�ݭ�����|w]�yd�\n�ae��@�ف�S,���Ĉrު}�t6;����I)�P,���W�4���~�At�d�Ћx��S��Ǹ㩏bD���	k�5K������pd���;��0rwR�U�n<
t9�wI�c}L�ns�+Tv�G\�w�V���e.a�9�_7ϻ�Sc��l�� :�Z����5b�~�o����8�#Q�'Tf�˸{	�/yV��Nt̲f���E*����T��U�Û�J�̉Ge���A�tGM��X�Rv�OI�f��/�f3B�K�Hi�hl����vy���K����Q��%wd]�)�u�T�f�I#�������8V���(��6*����荀i�K#W*����a��f5�m����h-��x�Edʁ�;�&�$�Gv��З}��TQ�)�9.�r蟱��ӰN�Vr5m(�Ӯ�+_.dT鶠T�^�p�y�͵����BB)kܜ44>+;���k�@2�_],�0LY
b���̠��`PWw�6�����^kxt��6���0��V刑1N�ˁ�-!:q٣�q����n�W��}[څ�n�b�� �S����La#���S�4NM/��9]��O�����X�_���������:e��MN�fg%/AZ�c�v �剎����ۗp=�{e?��
�Z�P-��dyA�ZL�1����w������8+t��f����c�Ǜ����u��S��E^�d�s� !me$�>�nS %J�ۓM���'���ƨ�:M�(���Ga�g��ܕ0�A�W�r�+��=�{6��ɠ�:J8���q�f�������`����m=LGx��.�s�9ʯh�3�vʬY՝|X4 A�R�]�l�$�(���<����\��]���μ\�JHq��Ї!u��\�J�lU�.	:f�<��<9��쥙-�x�5�RE��]�U���u
�3JΒ:f��}�w����J�v���6��N�F��a����;�9��z� 	�}oDkZb6s�i��tv�kl���ٸ%�AYg]����`gvyjUa����l����c+��i�yX�R� �H�ccNXX/*'\Y��k��"��,��l@��N��4w�4�f[����{G�"��̦V#�kp+-��;Aq�wt���b�;�gQݾ��:��:���DK��v��c&Va�"�$۽Mc��(g7�gt����V9�f�V���YnwJnN�e�9r+��Q�>U�V�c��Ԏ*#:�P����r�1��b8rM�������^=��ܥ��/6������!�^u �q"� OĚ4I��]�n��B�c��#Lf���ss����Nq�Jv���+��ww;���rwk�ܹaCH����N�Q1w\�렻����nWJn�tu�6WwK����I����4S���,�λ��쐨���a�n]�.��]���;s��˳BQݺF4�w�]������9]��N.���]�\�sX��H����ۥ�:���3�I
R
 �bC�;�4��29���ˈw]
r�Ld��uɍ�&F���r�`̘%˥�),l��s�Iq�J.�:�nFnQtɒ��f.�F]�&.�e78]��v�e&Nm���Ϋ��+�!(��wv�ȹ� B)G;2Az�?=y���y~枅e2���v����>�(�����x�dT�R���V9.�0�[��\&���܊6K;K�}6[��U'&�.S�s�fVI�!x\z}�O�،���lg�g0�m�NӪ�P��%<j<���ݕ�^^�Z�s��`k��e	e�X��T��w���Qf����L\��n�m�e�/)B9'��r�)?I�H[歷�w��*Z�8�jWR�I��O�%�X�99�N{xWg�ڃ��غ��n��'�j҅=�0�B<�*��Dg�Sܩ��7�������[��3lN=��4��B�\e@P�\��� ����a��^�Oa��4�>
��˧��������o��5n�	�jFo�h\�?I�M���������dO�f��M^�)he��t�F�����8^f����~�	��e3��nl��c?_��C�*q]�5O��\x*NI���'+'�����/�%�����[�Z"�ٷ\6;��RP���y���)�7��0�|'<|+�r��' ?V.~�ux_y?;�rM��&�n�nVnO���s��S�>��b]g�,`	_¡�"�ïU!�]L��S�]����&W�F�*e*U������@�\fm�{��J���=]wK+YɗE92����r��$���E��Ѯj�`��{�՘��V����4��ʛy�։r��ehm�ΌSU�A�Q[F�6m:Z��vNZ\��ǂ�&����]Z�q�)W+�����5Wrn;;��x-�b��O���R�� @KC R0��.%1ѵJV��@G����j��V{�vo�3�q���L��3��+î4͒�!Ґ5]3S�a٪n��辽�����vw|�g��])���O�k��i��#����C�����bx� =�t8Ejrn�6�y
X�Ү7�#�9���2�M�w,{���u��/\�;_[un�؇��xoor�4,{�q��iJ��Sx�����xj��\K}\.���6�I�x�'N(��X뵊�Y}�~���S�Q���Es���)�M���5ػ*\�B~v��PP2����Lz��D��x�ݜf����d���B�hX��.|4�i���=⣽D`�y�/I�:�[�>��Qq�0]��`wV ����+jb�P��g>��d٧�e����.��^(�86^������"���\{���ȼֆ�+znK�6;ѭǼ`Om+}]�y�ӡ�!f.
�{
�U�uǼ�b��hչ�i�C+Zh?O���ۨ�saSPG�p
Λ���w��y�,V��E ���8���h�Y�ى ����|�f�F��;1fo5�R�h��z�R1�;Tu
} �Uo�qֻ2� Y���m�1�UЛ�Nv��X<wc��p�s�nh�.)�g��7�ӷƢZ��)��7�)��,a�V\E�Dݟ�˪������㵡�7�S3���i�b4�d��ǞF
��9�~�JT�^/�rĮ3����=4�p��E׺��Љw�2>^���ɫ2�*z��_D���s�ٰ�)�mi;���fuT=8N�!�is3X��+)>
��.oq$Fl��b}�'��V��T���Sq�gHY��*����(T��x���]F�]�wV�	5��|Z|�1H����q��������
J �T���qt>���twcsޥZO��E`��xg���-@Q~�<Z7�[>��ꇷ�a�T�t��v*ȪU�c��Q��gZI��tR�Z*�y��J5���q�ᗍ;_C}P����a���j�٠��*M���d׫��h�t�}#�	!�b��)^Ϣ�͚������B��0�����hPsz��D��9�FRR�M�Q�*O�"�|f6����/
��A���*�X�z���K_c��<��p��8�ܴi5�cR6Z\'9�.j8�HH�g��@��9������~q*=��I^���u/�TCҺ�� αY��)ɥN��24x�1q}�{1��p�r�n���M;�s�I�}b���ٜ]�]�q�Bd��G��틯{�}�;}WP�ͼm���:��Pc��&���+��X��y�p�Ay�ɉZ�����w.�๽-�s���h+eTrJC��h5V�TD�%B�N(�8��{*�VƷY>�_�w��\y4|B~� Y��Ͳ]��/�V�=IɯL�޿���I�uY�y8�����P�^Y=�FkR;��#��E��p5��hYa@� ��ǽ��I%܋�jcv��_K�V]/
��xb��U���ꐯ����`�@a�P�̊fv���typ�z1Ƙ���bn���5�c���a�G�����Z��}2���t���*^A�Y�mz�Fm�)�*���6��-~�M��􋹎�P�a8k2*��#��+1g���(b���I�/��g�֓돱���k�|��h��u�Z��F>�V���rZ�Ɖӣ��z���R���o��Fm���.��߽ڎ���l^Mp��p��ė����O�8S���{�Q��凪�:�0:Zl�'u��:�1X�)x�{�P��C`np�r��6�O�^��3���3���q�G�(?TF�}��W�g�	���X��F%����R��!&��s}@4J��o�.���]f�`Q�c�\�D�w�ט�xlߖ�#�x�V�]9^]6z����	�y��TJz��Q`Ɋڝ;�m�d�o�BCN�FO;T���C��Vm�,8�<���O�3�J��A��{FX��xIY�a��Eߏi�ECBB�9j�ץ<�f\��xط����A��|�M+(�{r_X[���>���\2��/#���� Ȩ蚀�����$�y����b�dH�{���Op��N?��;M|��FSuL;��6OTt�=Ң$���P��q�8�$��k��V�X�[��U�v����i�nN��茗+��6�,�A<�d�q�>]��1��=����9���U�V���u�b˽��g0�������3p�4�sB�%����櫻�>���Y�.A�r�D.�g.c���Ԏ�y1Ë~��Ù�'�Q�1[�7Bi �_㟦��.��S�T�=F�BR�S��EK����ƥu.n!�vf�g�yguB�o��s������n�KS%t�ɟ%q&��E�@yf>;���a�0�j�H2a���Gm��k$*���S�L.��Q�2�>���g��Q&�T&�#�^�f�g��1}7������u&�|������G'v�Gk@4k�t�N�:Ck����h�,��c��{����I�T�	�T���>�0K�	a_,�f'�z���X���ƻ"��}}Q���b!���Em�l�ap�VGF���%���;ngGEb]�9��\��咟5R]�^�̓Y��Q��T �h���6�����3%��r\��e��IN9BZ���Y=��=�.���yJzb���7�&%d~�y'ߪ��~����߯��V�z�⼶��x�t5��&���]>'0�){n�D��9O��g�G×x�éw��;����c9�7�D�z�&4�ci�'<xR�Xg�ۋ���W�����M�����F�p1��/2����vǵq��zJ
� ���x@�0���,��j�I�J�u3����䗸��m����t^��ҟ���N�۞����R�@:�@��a��/�!Ħ�=$t�3S�����x�6Z�_E�G�;�u�m>Lm�,��3d�t�|N�A�GgU��ڱ,֭�������bM�c��,U����ީ�|27�,uǵ\>�r��p6lO���l��F�Z��I=��@;{��Wr�5�^.=��s\�;Qm����g�����n�sy��V��I�.2���2 ���[_E�ֆ.%��]�p܆��(u���y�����CMuYP�)q�"��t*=���i�젫��vT����������<==s��*�L��(A��?ku*#w��>^��6�^�h�ү&վ�`�{�rTƒD��2�TI.�v�����X�������y�H��(ʫ;ט;�vxT���/�P�jK�m���"��'P�T�&;Վ���*���b`�o	��64��sZ5n�Wܒj|	=�4��h�=�b�f��0�Bp6V{���ʊ��stѮmxq� �q�`�0s���*=2_���=��N�8VuC���v���zȤ[>³mGW��j=�̔jhwRZ��ϕ�=7��M��+�E����u�jz���pٳ�*M�=U��ϒ��}�F�������@����O��5�~�o�e$�&������^	��>-*3|��;\�s�c���׋�p�~uq=��q�/:򕛈�I'2����c�Zzk�]8Wы�t��_�w��7A?8��H$S���'wk�;��ѵ^�@$�^B	��L�=zr�̿TmkdG1����s66���l��c;g������k±��}�6Oߦn�3�=P�^)؍��x�3uX��g�Z<��t33���u	�������AI� �T�Q���2/�W"��wG�7�;�U���%:��C18�Z>�-�\'�o��<k:}�x�c23��I�����Tȭ��f�-���<)u�xL���L�L�b����
�Meu�w�
 �!�"l�9i�.՘hv��2�c�n������ޥQ�����^�
g!:�}�"����y�m�R%v��r�y�u��I*�D ��"G1�4���t�2:o�1a��ᗍ;P�T=U]���T����7�|R1N�- ft�}! $��6.R��o6jn)�^�/i�	��15޳55@���{��5Q,qO���p�wS�w��E��"�A��{�O���v"����}5�őJ�;��E-
��2�?�80�nH�	�p�s2�~� }+�F���(
�ij�[����Yj���z=��%�s*G��]�˛����`4۬�i[+�����U�3�go;�"s}���*��oXMOx����~�1��M�_�e�L����#"z���kf�+���H5;ב��ҖB�-PS��(K>��2{��w��"�~�C��N�0cc'˶���LR̠�}��RR�Do�b5�P��巳�]{A��7�Wy.r�ٛ��2�k���Y�;0�=�Fkj|�)�\,5���-wFO��S�sv�k0�Џa{z�`Yuu�pwc:L���|���v�I����)�T:vn9�^{�g3Ȁ4�#'�X�0�!d=@K���UN��ڽ���T`��CI�`�N��J��Z]�,F� n�KxcY�
U���w��� �*L��P��ђk�\14�x"�4w=Q[z9>$�P!'>\�R�s0��ݸ��ѬTw'M_+kͪ��W,���2�q�cv*} ���Bb��dQqκ�_$�I���f�ZLO�1���kˇ�Aӷ.ʃ������ͧ��n+=��	>dV�����G�Mb�T>�>dD�[�۵��W��N��q;aN�:��h�$���5].�"6n
�j�}2�4;�<�k�'��}�'u��q�H������?c�y)�r�F����t�S/ơt�>�!�~�� (�pt¾i��զ%�,����H�)7�Tu�M�ׁ� R#�
��$���=�ԇ�ڠS[�ꢋ�ў�{���y
a������ϥ��1l 0*:&�yw�سT�25��p@�C�:j��~�{=�+n/\-�񿛐�v�;M<��S�͓� t��P�P)�\��|�S�����g}�<Eh~i��\Sv��/�i�7'�[tFK��r!��g����N��zGf߶}��06=S���piQ~գ�'�w�ws9��n�v�U2�ӈP*Fx�"���Ʃ$��&W\��TH^Tfˮ���G�]u.�W�s>�#��Z0 c�o)�f	��n�r�Xx���G������[5���Ն���V�r��
�u<��/jy�f������/�L�RF��t��G�^>�w,9����YκT�V�SmbI�5�j����`�ju;��=��-���63��[H�S�հ}�8PըNvWI�$?l	B7�ZC[GC�tjWR��Wfm�"}r���9߳Ѯ�H�xN��΁�q��9�(�tѨ�_�A�P��f�gF(�9�Wv�s�ƣ�g2�h����7D�� y?��K��(^������������5�}�x{'#ՅU�����ǡ�b7/.rwh>�L���.k�!�C|�\�� >�rǔ�O�{eSד�y@�l�zv�4�/�,��)OL_����Ɠ����/��S5�߻�~���Y��&��,b�d��Sh��,����'맷/�%����د�5O[��]��w���Y�ע;ox~N��끈9Q(迋��+�K���퀉���.�_~�ǁ �ė�������g'�g��Sq��P�V*:ʃ:��KƗH�H1�ܽY�/%��^�>��՞����>��X{-hដ{jn=��R�.�#�y�JTp�B�7���U|a�O�sވ�ʅ}~����o�i�cn9exv�D��.�i@:�GMp����?�©����T��{��ur@uΝ�w5^g3���˺cM�n�: �4�_rȩa��xd�ch}�]͍��t�s�0j?J㏜݋I���kk�������Jt�JoX�c	o.��i� M�lU�r�vc����
�4#�'yP
d͘��%���¦ܒp�t�m�����1%6�qB�ϑ�̝���ɼU��%.��olv)�&*�q�EYt�WY�X�%���֥�(k	�7.[]�:���͘��ΕKp����v�q��*��wwV���#�1��w�{��l{��HudFC2y'1�殮R�\nH+_4f��*�%���y~ǧ�=Z�=��di��J"�cЪ�y٨�3�)�쩲��l7B>ko�kn���J�1�yf��U�j]�|�fV�f��u�\k��%��=�6��K�ƨ� �\�7������W$��֋V�	P����|*S61�:Œ����)h���&�Y�����ޑT6yPt�ճVBN���՝��"�<7�QKe�QJU�P�ΠeB����^^˳���[|E�v1(K�[��A4uto2,u�>{N���ܧ
�׏��ʘ
`,�Ԭw;��zcA��ҕۉ^�/���,�N��t�Bۼ�dGJ	K5[N�B�ϳO���m��Y�nr)�ݽѾۛ)�S0��t,ї�(��R��n��|�XkH��Ǌ�`ͥV�K�aV�����{�z��w8~�@sU%�e�c��i�O�k�I��w�ʚb65Fݍ�H'��D�PP8ﻐݺЩf�)z�z�s���5y�G��B"ev�@=].�܈ʺS���pk��5�r)rjJ���Aԓ���(�S'l�!�K�����%��X�waيu޸P4�=A��&�WXW��j.(�����`u��-�o�YJ�'k{y�ƫ$.ec®�w�vF��Ǳ���[*�:��)`��[�C*Ju�>����J�t9ܞ�ػeZ벋�Q�G-��u0nCt���:�F-���"uu�V��t+�d{�m��[�w>��N����a�*�#us���&۬��CY��V��� ۚ��J�^m�]�`$vQ�J�X��[��g�" ���!8�ˬ��X-��\����v����ҹϟk���Ǩ;�y�-�����]�P�4��뙤��7.�J��H�f5D�Mw}�����QG.�R����K�fT.!#�.��g�t7��j}�g,dM�ܤi������MC�!<p�S&1�Ղk�����WJ�ԣ�0p�wB��eKX�.��8�0��\z;���q綫H౽1:�}��^���e�CNG����n����u�f 5��<3唞*�s�J%����^�Fy�6L�
*�	��5�y5��y����]ȱ�[�.es���P*���L[Y�fdd
����J�z�Yl��k�Ӂ��-P֣�ٺ��b�)������))+�����^ur���v�p
�v'!dfy���w��'8���b`�12$�wk�`���wX��b!'u�cD�23d�wv�u�6���wk��]33���IL�����t���ҹ��I���;�;�r��J�sns�7JP0Ȥ79&�ѢIb�$&4�t�3�3%�q):v�BY�Rwu;�LF�
Lgu�L�2*%Nv�K���wwb��2e�л�q�S#t逄Y�Wr�a�1�]	.�I\���d���w7@�a(\�κH�I�)n\niۂ�JQJwW'.0'u�*BwN�(�f;�wt�s���h���fI(��&!���p1d�����vE�n��wR�9����F��)��L���Q���ʒJ(6�r��K]� T����L��i&r�0;� �('w���̼�rn��\z�/n�kAL��]-,�8�6z�� gh�H����:c��'�W[�&�a���8���`�T̥;ij	B�F3?F�5^��׋c-�b�;���!�ӌ�8�T{:�e��f��z�?e���uO>���07_�l	��"'��i�OՖ�٫���;9�{�hlk��jۨ8����b���1��ׯ67�yb3�!�xZ�2�EL�HlL��R�pW�Z����Yw��Mk��`M�V9�f=Ok}X���N�Y�W%�Qt*�ߐ���ML��^5&(=yP��#�*F�/����=��Q|�K���O6f�P�Z5n�TrI���{Ɖg�ښ4�iŊ%��ɞFq�dl{��Eǹ����h�sk��e0;��;�L�S��4vhe>�Q}��ױ�|�u�N!M��kÚ�C��H�βQ��9�HekC�tϰ���̿O���S����T)��x�U=�Fz���斘�k�Ѩ�s��7Jv=q��.ɫ�y4�Y�惟B� ��~��b���/	��d�5uV8^�?\c�^���������{SNT�P�����m��@ہQ�f�D;���8�����Fz�ؓ;���/��o&�����KB�i�����}���2q�9�Z*�;n�$A��rYut��̚�Ќ�����v���DU�'--p顯&� ܙEV�،ʰs��e͑gr�L�t��B҄�GWi�z0��f�;�&��_����w}~�*¬xm?t�k��9��}��ˆ֓�fa�Ps�:�ZXds'�o��Њ�ןi��� �|�DTyrLNC'��V���+!{�M���!cà9슬�bq�x�����3B�7Y[�c��>�q�D���d�ɕ�Y�lu?�^�R���
J ��vw��=�ԗV�e���I��gF�/f1zG�p}����ţ̶w�ꇷ��&���/L�s��og�i'tgK�� �3�L�xT)��/�;](t�s�0k�</�v^v���o�Q�ʏgWX�$�*gV18iP𮙩	3��ߍR��ׂEDOs���Ә������ܼݯW�a��a���xNn�C�RY�3�Q�2GR�F��LIV���fּ�=����q.%�lR�sͭME��ڄ�MsJ\��@�A#L�{�=^�k��Oc}��wf�eE�J��k�����l����[j�s4��d�n��J�X7�Fkᙛ[����
��j_q �7�3��SF����Ù�K�+ ni��p���v���e�Z�N�uqQ��c�J�C+Ղ�c��U�]¤��8�(�hȺ��g#Me{��y�:�!�:�x��"�겕��x5�=�)�4�qe�9�殛L#4mʓ^���;Ȱ㹚������2b��]�l���>Y7v����ڑ@�'ʇ������#Ø3^���zoxԶ�$Bk��q;ֽ�83NuЧ�#6j:�,��;��.�5q5� �[{9״�s�U�K��I�ؗД{�L��"z�8Ԯ�M_R����u��Z�t��d
��9�:�5�j�/n5p��zi ��=���V׽轴-Wx?���n;Z��j�N��9C|��
~�M��l?�b��V��I���n3wsB/7�i�����uxzf^�K��I�����_s�����h:v�]�y��y�n�Ӯ<93e���/���βD���mڌ�ޭf��)Џx����.�����>2�p��fŨ:6��-�r����F�י���gy;�ݛ�"iG��5��j���%�E�+�Nr$p�)��_.���(?W�z���T3юb��{V1{ir��Mh�t�����=��Ȱ����"���$.	�Jy�˗�i; *�_���{��(���m�@v��<>�X�:��6� �TtM@�0�lUd��Y/�Y��#x!X��7/hEY�8�Sw;F�\޹���yXX/��*�>�l�&cӸA�CC/d�M#aSkf�[W }�:�/N:�k�wwwHj@N���Ӭ�a������#�&�W3W"�����S&f��G4���\����`\�н��=o��^��ƀ�5<�e7Tø�3d�t�=Ҿ�:K�퇕=E�V�>�ꁝ,��e����<�������L����j-�#+��q�m Yu��1�]R�]��x�Q�N��f᪉���)*C�qq�a��"}zR-���Q9��1>�'�3����=�iA�JY�)#�P$���zP�:��,y_��uG����ߨ���q;>��e��� �����������Q=)ɯ�2Gz��(D�jh��\���g�R8SOGp�i
^b�}�w�cA��S'��`c��Q�s�P<�4}�$��;J�ڳ�#��]�Z���
�����Y���G��h���ʑ��ƀ�\遥��e�q�>W3>�hv���c���=�*�y����c�OɌ��A��z�1�斞�րh�S�q�#5ȹ�����W����0��{ht���:6����M���V]mG_���/���7�sK?~���ާ$<�͊�ﲷ4�>$�䜜���򁓁ɹ81zY9Q<_�u��O]ߞ�v�
�"�z��`�,����U��r\�kd��L%�6���6����NZ�N�<fh���j�p
�bzy�wYX�r؛h1��R%�I�u�T��:�&������^*��Y���ޝ n��.MS�L�e���c�N��ͨ�!{i�:��$�]<�E����'kD>�5ãޮ�Dz�kPsg(�.�|�4���Nԉ�Ø�ۋ�뇛V4a����f�Խ��U���������|��l�T<Wv|J��\7R8E��ї;�W}� �x9y�h�O��u<;\'^m�=����}u+"� 4R0�k�[�o���$���ZN����+���ʽ6*�#Ż�Pߦ_K�Y^qf���� ,�h���S[���g���}�>��S<���<gs���!��c��i�;m��^k����b���:��i&��}gQ�]3
EĆ�E��O՟E�vj�S��ﭡ�ީ��Eb�p.�b�f)�\^���+�f:��x� =�@ـ{����V�5��D�����j��bv.3V�ƇD�#O8�-�k��Q:i�:�\�O��|ԅ���&��0��Q����p-�r��^�t�368�m��:���&���I��=��f�f��R���q�詰�N�eg�T:��SF��^�C)�1��V ��0k���<I~���F�7�_�|;:�J�D5���X*2*�����cx}n�n4��%�ƻ��]��� ;[C��B�fq�6@�}̬�\m�Y����1i\bt��Guʊ�-��z3$�%#������%
���`��̽]ɱNC���1��-J��O��ɠ�0���/�^Tww$�Y�J/��_	�z�Y�@�<f��5-�P$�r�ע�O\�d�4�l�Az}&�i�1����^�B3��h�����v_�>�T#2��8~S�9�ft\�* #=P�ml���L`���.�����5U=�l��i\vz��k�$f�[>�3�#:�i��w�����R�7_�|-#^��̿�ցZ���yԯ`Tz����cW�'Zǚ~sk��9�k��Q���mi;�â/��V���]�D�T�ݾ%�����.kV&�exK����Q�iR������!g���*��@��/�¼��8Bנ���薅ƏD�����LͮQ�v�:�ۏ=���#ᛆ���#���XF:^��z|RX�>'�3���i*�.�:��3q;x����������j�R� �<�p�;�x��O���HG�]3Rl�*n	�'Y�[�=5���k��cF7&��
��������Jz���pyc0�N#Ǉ�=�t	�}�B.{�|�|<�+��H2�?�$y���P�ҐO���F��7ߌ�zFi�z���ي�0�58�z�.�1]yuf�F�#��Һ�Iu�5��Ѣ4��	v�J�C��A�m���h��)b�]LJʊᓻ��[7w�Dbr�_�u�}�e �n�=�u��"��#����ʹ2h=i��g���s��A�� ��>>ϵ��k��p�����h�\Dr�1�$� �30�ۖ�ԪȲ��S]]>�C��\U�&�L��!��x��6ܑ��W	�3.w� Ҿ$i�����G�����Nz'���x���֊���]�˛���/P۬�VʮII��Xe�WuJ�d�ܗ�h��Y \���h>9�.�j�E��^@xx
d�}�`�o�jWo}��y�I}K$�${ђ�Ĺ�P���UDd��Ԏ���R1Q��E�H���O+�XZC���FB�������0��{����c�}��Lj��s{ʽ�!يp�ֲB�;��n��{�z�2:�{ ���k�d�Lv��1ښ�4�azJ�G�w�;��v[�>~��9�d�2;Z���t��9C|��
~�M�Ǝb����f���Ӄa��&��x�Lo�]��K�9��#�
�v��󭑣U��������Zs�;P����56:�V��{���p+�T>�:�����pݨͽ��T|��f�L,����A�q�e��c#6���<�^�\���K�T���h�d�:��;ӧ�n��flP�����{O;߰��إ:��%�
���
3a����*j�����՟3�pK��{��A����nF�O{s��5�Z��L�O-\�:�;���'6S��X?}��f�RX1����^gE�!����O�������i������I��L�"��d��L�z;�B=��C"� ��s�����j���R½�>W��6�xP�a�w��qx�����	��+<a��^�
eH�!!S���$. ���o�q2N����s|�
�9�-Ջ�q/�g�e��޷>��R�8a_� "��k�/�;�����o8��/Ƕ\)�f�֠����~rN�4i�y�#)��O�8V ��̧N�:�w#n�Y�I��v�!��5�3Ǵ�S{��4��lm�9��lS���;[�vF�Uu�{�MT�@Ѹ�1�@@�9�P;N��V����w�ws8G�E<&O���o���B����i�uU���(���P3���7C�*���N���U�sً��w�|4�ۻ]�,Y���E���=|Td�;u
�zS�^�#�QT�Ds��*Z�8��*�i9��}�k1b�����`�rH?w&K�fX�(�3�]@_G��F�d��GiB��Y�*�Xu�գ$��ޕ@�X1r���Z��l�!���2��ʾʻ�6p�ɨP���Ð\�-$���OH��_�U�7����iNtː�r�]jf�$��;D���ʺ��F�����*Ú͊ĩ���!�hB"��J�9��41����sT�=RB$�P|�N�a�z��JG��s��q�P��P>W3>��iWH��t��e�w7��3�\�p�n�^i���+.���|�o��5�p��n���C&j+(�X�#�F_�:�_z̩Le��2�NP�xd��ٱ�}�[Q�R������bv�>ܶ=�:3\f�{�>��~��?�ՠP���������XF��_���s5�e���%<�N7�S�TF�j��=��H�U��{Ί��v�E��jt�s��٘v��
W+.��x��9����v���������p-�ߩi����ҕ��Pȱ�%
������AmoD8��_xz��k���N��	��V@/�ܼܬv�~���4<*z=��R�"� 1A��b��Ӻ��.�ױ}���q����. �ؽ���aj����1�7鿓���ܲ�:�͓ΪD��k����M^�NK�|�&h	���t�)k�n�W���xn5��|3}R�{Q���j��F=B���.Q>��Y4��)��5*��<�E��O�[����N�'�����}������Ջ�V��yg�
�E9����w�e�_��wT�2щ�����C�/-W����I�NX���P,�O��{!c2�w0ÌÂM8Wf��C���[���]uE��}��b��EW`�s�W�o^��Φ\�h���MQ�ε�F
5w�ԣ���`�%p6�>�7%����|d��� >~�����Zǐ��4X/v���Я�.�xn6�Ix�NuN�WܥO�����`��
$��jN92��ݺ��Ӄ���w!������ľflq5��T5n�\C$���B�	�Y^�r跾劼����H��a�v��tj@�m��ׁlK [��(�t��䭩�mdV��|����$5ල*��4vM�|q��s]���$�vO�(�m��C3��C-�B%ͅ����%)�C�yX�Ղ�ʿ��%٥�f���7��j6a�^�B2!����G��Lf��y.�SYR�$s�;i�s~T G螨j�N˸R��ӄ���Uc��
���mm����&�,�pᶇ�o�r����P��;�Vn���Pf���V���t�8��u�2��;�^EO�̦��UH�T����9��F;�C-���٘vQ�(�ONDι����ұ��q�/�^�T��bj��#�'!���}�*VB�Z��|���@s�>�O��Y3*#-�׃J�DA6�5X��� ����2��f���ӜΚ��R��up��_"���1�b���B�K���Q�pb����	u���/-B�]���������ݳ[�}�i5/oaO4x,H��8���
Ά�o��0�ˊĮ�#qJ�67��n#�PE,��60檂���7t�` 3�9��p,u�����s�e��/������c����7V��-�9�4"����>�ueQ�A� #V�k!>Vd�2��ᕼ�-ؽNa̩�6��nC�ji]ݗ��c��ī],�h]��,R՗�xȉ9�^L�l�t>�:��S��Q�+z\ O'Y��{v���9>f[`I����V1�����= ��OP�'#����:���<!7ь��cP��SV'�#�[|���g��n�����c,sI��H�3)M��v�$�6t��gmH3"���1�J�4S�8��x@�%�٧�B"f�Z\���d9b�h�@����E�h;�4�C(u�F��N���y 4���Q�n]GP���b:���X��1��m�ָ2��e�fC��8N"�l�ӆ���q7[�ܳ�K�({�0Ri��rٜ�n��JN�:
�Ҋf��z�0>v\�N���(v-�I�K%�Q���u��޹w�J��U�l�T�8ӈ�QQ�k��f��$�dNrY�y|`����J���4��<�b��4_CIj�:��̘OT���'�e��+E�"��:���S)Kۭ�p��Ⱥ����Iv�t����v��"�E]Y��#(e�:�}R�3o9k]�]���� �9*��w�[��@e�������b�tw,8����r�ȿ��K�F��y7]�Cي��8�s����fo.�U���9�����^�:�'b��g����F��a}N:ز�@%,]�1bq�;;0����=}�(t�3��WZڕ�ɵd4��Z3V�K�3��27�M��Rs��[�mּ�Y��8S.���;�\�
4�4Ep�'N�l��/�$�$	WKQ[5��@>��m���\h[ͣ�E$eFU�qY�ȓ�Qs{\��}��,wP���	B���uc'B�>�a]!�R-�f��O;3Ú<�ף�:�؂��w�����(���U�-CӾ.����Z��D��=ͦ�Eӝ1$�F���Y��s����5�� ����������D����\z�h;I��;I˼�8D��x�Mw]�8멮�
��0>�kD�C���C��;�j�r )�+l��v�`<�yU)sF����ޙd�R:���kp+`��<��RQTP����ڇ]�ʝm�-j���H:\��`Rf�-�y))�wV>�f�z�3*1���]��U��R����v���!VLpϞ�kK�@���Ԭ�KU��Л����Do<��m�ڼ��G�>X�sWr��а	�����jP�ĒˋVv��sf̆���������~z��9�1w]�HCB1t���J����)!+��.;��w]&LhDZd.�bćw,��J ܹ��5��0�1�)@"���;�#�ú�7A �2��]H2s�bIHRI��.E�)lwk�.RN��6,\.L@�\��ܹ���]�ܸqI3� B�倧u�.�rwi#sv�:����%�FX��d���3wrI%�'\��F�w\.\̀&Y���d;�]�r�I�35���wwv#�,II�C
9ę��2 �RX\�9ғ	�f�s��F:n;�w]Be50�r�0 4�wWv�]�u��;��I�fI(�Pwp�� H�wn��I�d��+���wl]�b4��9�q݌!�t�*��
|(
(���rw<e�[;���`��R�l���� �WYQ\��і��S��R!�ҹ!< �7�ռm��a�R�n[�:fg�c�@�0�x_�(����J:�1ɕ�6�Gq���c�o��z��
Qu��ț�����w�Ώ�z�>t���%�>UԧW+�l�����1�1����8��j��S���՘)�}�8��U.ᖨHFt�D� ��"�ɯ'Yn���tŃJ���<"�ݏ+���[���u4a�;�ϸi\0�GLĤ�=ƾS>|vE�t4�o�}!m��xH=ܬ8o��r,���5�:���xs��Q�438�ץ|�Mq���B�3�tW�C�7��U�k˺���x��j�Dm'U�k�R�����5�EwQ�Vy{Z�Ɩz�e����iW�*:�λ��7�����k��`+ez�J�T�	�7n�Vf�x�K�M�.���ȗ�٧�gr$?�v��̿�9�d����/�d���*��s�=�r*j�v�I�L��CUӬ�p}KA�����5-�I��'�n���x�ߣ�b�N[(�� g�qQ��E<�BWQ�s]�5���^�oi��k�g3��*� %��6����0���yZ�W����f�g/=H��U-6g�V�3<�Ho�%ؼc�4>5b
�3t1uo�����_W*���iW
��wn���;2]�Ԗ��$qcR�T�S��
���#���W��ѵSy��f�J��M��\�����r9Kg�8���a�q��td��n�������A׏��ԍ-Ȫyh�����}3�}��eT[T:vo���wt�c�$�ǥ^�ճ����oA�q���j��3�e���$�I��Ly��i1>�{x+��GdT�K�%ת�j}��>�7�^�F��V���Qz���y�.%���a��qY�Xv�rފ��\g׆�թ���j:v�f��:=jZ8*H~��2�C���k�%ڊZ�E�9�p¦s���cK���|2����w�F��(+W��\٪�԰�hϑ��\��PX�{���II�P/�3��='��6}p��{qҳ�)�ʖn��>Fa��������a�MX]Sw��*��a~�ԹHa����Ջ����c@v�7\gJ��=���a 9�P��yT�	P>�5�G3����j�-�������G��ӷ�4i��R2�n��q�a>Y�cj�;�]����O��/�d�D�bL�����k�qW�7i	b��D7'����ّ<���w�@�t�����Fi5WNW^��w��+��w<��j�w�P��˰Of�*���h�ʕxg5�j<��M���s;�wj!R��!yë+g!۔�Ō>��P���$"�d���z��WeN�dgX�k)��`�����&����NӼ۩*�������m@�<b*�z��ds�)9��KȊ~��dg[c��G2�Q�nJ��wz��=\�+��Ww�f�&�T��|�(W˧Y�{b/�R:g�C��3��*�ە��'wǣ����Mq=�Td�;u
�'�95�;�%��M
�������`q9�~�WO_[�p�v]���#��z�wK%�2��|j0�s��t�92K�;J��<=�6�g9�w<�S�0��1��^���萡�@r�_�8�Q�2�(|�f}1�S������/��v=��;��͌��i��=�F]]G_��U�q���K��?Y�W�zu=�v�=KiU�>��~�3!2��Ѳ�N�z�м7j�{D%�b���y����N�	��Յ�4�f�9''+��чd)�pT/O�s�On8<[�z]����Q{]�͙��[��Y��r��k[f<��Kg	�ߌø9��!\�3���	9ez���IR�Ϣ��h��'>����ao'Gc��tl�z��u�vc�<T����1�^������V��Δ��{��j.�QiK;չ� ��{�n�&� �J���=U�W���eC��|���fh���^T�;�nm�8�ǋ���n>H�"��n�:��>�}j&fA�2���78-�[��%팉�v�\.3�lRl.L�S����W =ɑ���@/�ܼܬv�~�����Y^�eH��S�O�\���S@p�j�6�ug$��|g�l���>��j2g����W��-�:��6�&6�9ex3�;������Z�ʺ> w��� 0:E@~Q�Ot�|��q\g��rv\k��i��T��s��^T-������F��ߺ���6lK= v��`z|
�_t�D)�?VE�vj�S�[���.�%�c��lp����F��PrZ\c��Y��%3*g�$6&H�^Tb\���wӜ���O6=j._��˃��k��9��!㨝5��*�*x׈��P$��R&f��Vÿ�{�6Q�11�~ڐǹ�x2��-�C��m��:��G$���'�Z���s��E�c����v���c�/�pG��za�ԁ�pڶ�G6���S c���}��w�g\L����)����2�4}j�=�C����A}/VJy�F�a�v��;�����%m�5�8��eUG����8N�!�#���(����|�Áw��9Z��ƫˆ�������b ը5�u�§t��1#�FRͫ��ʰ�ls��1�lm	��F�v���P�]eLtJ�V�Yt�n�/�(a�\����V ؚ���ʸ���}�MN��U�T�]�����pL��K�D�ٔ"�}J\B�s���Ҭ��&��7QwO��u!��0���$�D�팜�^-�̟Ҍ����9?g���{�Zv<sO��C=�q����-5�<�Vm�I8����	�1�r�����k؊IUu �fk=~�g� v��O�[��q�h7���Y����z�s�H[s���E]; �C�,�}���p�N%f��N��"��QQ�k̋�����������Q�$��1#��m�i����|R��81���f6\�ȉ.�Q���̞^+�)�6;���m���'ݫFj����A>S��t�NE�AKÝ���K�*^#�p��^t�:�-���ت&8�_����v'���j7����Le��Q�>A�EMP�u�n��I����fzﻒ��QV���یhq�o��|y`��6��x�'���d��:F��`�J��o���:�m��x$TO7X/�9|v�Ƈ�x�'i�x*H� f��@�Q։Z��-c�B�w����|,�z���]6�N���|ڌ�m��'U�j9�.}5N|X�<7BN���n�J	�l�}����h)�L�{�t�����}I#K�e۰CZ�>�f�$�A��k�����p4-É�ڕ7j��*ƕk;���R������W���U��g*7�t�d��&.\�.�N�/{��j��Z}/$���jj|Sr���~ #����ϞP���95��\a���p=Y����vE�޸ܛ�*-(��'N�n�
�T�_�RRX��ސ ́ӢTB�ac,e_�v��M��^@x(>�sR}콎�ܒ`%d9�>~+ [�l�D��צH�T@�@��P�v���9�Ԏ�
��P �%u][��}A_j0��)�p1�qQ���d�i�Q��Nуۊ�.��Ud5��F��	�Sy^c�(�q/����$�����`m}u�����td��Lv���)�P�1��P�΁��Ϋ-��q���WQQ����h2�ڡӳ����T��>��{���Im�ڵT��x<IؿoTl��d��l�Y�*2�k���zo�,y�Ɠ��c��[�kv㮧�NO���6�"I5�B���'F��ӓ�Ҵ���̑C�-~Q�&w���[�Z���p����j�K�f�FF�����j�ތ�1*�Ct��t_�����b��v����E�sW����X�������;�ݾu�-��ӱF�ݨ3�h���<G"��ǐGK�����i�]vj,ۨ��m�+�K�z�5���UpPt7B�U���o ���(wiԺ��Wa� fDr	����7�	0�i�_�y�b�|��'�`%Ɍ�ICJD�� ��8G��A��&��bUᠫ]�u%�t��.S�����G�>|��BZ��JT�^B����E��17�6}.|q���5>�� t�|2qS�My����wc|���2,o?�ԇ���X����F�����ϸ:�R�Oa�.@)���$:�B��ؼ����I��f�����q�3���t������C��r���Q��S�V��tX��Ư1��jSD덐'U�3&]$/�+���^ۊ�n��'Y�l{�4s�y�G��Nv�[}d,�)µL���<z �툙fr�X魐�gz�Z����m�Q����N*1۶�}#�h#O�ݒ��:�֒e�M1!2�	���Fn��ܑ���F�9��oku�5�.B6���E��3|MCj2�n�2��H�T	��jh����Q�U�1�}��7��6%)ÝF{�"{�ԅG��%�X�j0�/;��x�/ū�h>��R ��w굅=s���È����f�E��9����T�DvK��04��2��P9�������+syxʕ�M��VYɱ��a�{����]Go�Z}���ܹ�)�q��ˮ��r}#}kf�4T{���E)�'5yiÔ���� ԗi3�j��)xzPڹ�(1jI�(��R���`J��t�i���]�댦��a�t�(�|��Y�֬���<��m,�$Ew�f��yp�Bg����{kȓ�^4	�s�܌\9V��&GBP)�U7T$fBeGF��|}1Q�@ Pw�cF�����ECH(�z�n���7�,U���*������~��|?0_��+C*���Cr_�)�P�\��M�Ff`��CI�
�η��ܦw���a�Z����:��|&��7_���د{�o&��b�i�d�w���mX�6ޯ
���K�
'� �Y_�H	ە�"��*L��uq��O��7ơ9�_b�<� o�y�Y���u�^y^�eH�e���P�=�n�o/I�'��'l�aԙ�5�=|k&X�}Z��-������c/)�*���\�=���-O�u`�Ґ?Ut�5P�%�x�3�}�t����3�sK������HV{�	�Ɣ�{�=�yc.4ؖ��b�f��JA���,�/)������ze4��9����E�
����:�dY�[P-Cu\c��,�t=��l�=�v|�*�M�;ջa<������dK��^P}ޯ�����a.ډ���(������ w�� h���= v�ώ®,�m��.��%:Չ��#7�_m����b��7^Ξu�o��wd����J`��m>�ًz��|؝���9�Z߸H�h�ˡɉs��`�Zv�m��G�v�*���o2�=��N̖����2���WJ� g6q�g�kAD�.(\+];�Q9�?|��P��~ۑ½ϫ��:�`��vk@�j���I�a���**���ǣ�������P�5�ÿ�W�.!��ba�~�Un!�|��\�ؿ^{��a��˞jUD�/㩆�k��^��/C�c{���X����:�bCs0P�
7��}	a�Z�Q�=�,��5�RǪ͂6�^i�_d�꺇�^��쎼ܯ�H�^y!\��Lz���s��7HekC(~�O��&;hb���#l�g��u��nZ���e,�{��ᾟmC�փ5�q��p�J�|�$b��j�s����&磳6���m���m1q亴�r~sq�Pzo�Ǫ�:���CkIݰ�;�\DuĔ�w4�:�ⴸ71�i+4�x���������E�Lozr!�^����}�#^�פ8{�+���ꪯ -*��ƕ�TuW7͇H�g�n�϶y��b�hGb�}S\pc��H�qطmO�[:B��(#NQ���f�ʢ�.�����]t����۫㼟쭦�	D/�K%�-�w��wo0��F`��f���8Y�.�w3մ)��a=�c;ej�U���R���r2�T��`$�ұ�|�Ve5�8�̺A7`�R��z�uN�l��L��Cxj�a)s%��S6�WF�+l�d�x!�~�~�0��Ƕ���ȵBB"��$y4)؂k�ֈG���W{ބk��žn��x��G�}P�b�G�õP�L�l�4X��9潲DZ�\n�GYp�py���sV6<���r8�x�'Ct��B�"���'`����9I�?T�=h�.�"=�>����=ޯ��wQ�j�Dm��ۚ����
�^��.�eշ��I�Լ 3�#���>�נLv��P��l1������3�{}����7Ë��3���}��|I��P�L��xl�4�zw$?���p��L��*;��u1S�ou�b�׷@CΫ8�gc��l�A�NMzd��T��(T#�fϙ�������]mm����TU9���b����.>�Q�v�5��)f����}v�:�*�E��E����p�.b�j����
�Ƈ)�nXQ�P��F��G�ѓ�F;i��.猛�̃��{Ds��[f�x}���.���5��q�U}mP�پr��Ґ�".��P^yb���7����X�KG�iU�:t��QeVR�J걮��.��<ƾ|s�j\�l��H��CTԈ�6��[�QU�����R[�]b�5]J���ԩ:��貯�yM�d�ub�p(5�+����F��͉[�v�t�<��3�x0�����rX�Av���hf,�P��ѝZz�K���I�t�j�̾�b����y8
�7�Ic]�X7AU�S���/��.oV�Y���m-uy/)E��ArSH�V�mT��4U��k�
�C~���PSg�;�_;�)c�dԆ5\���MHpB�@�ڛYՉ��J���m�z����E<�s������W+{�`�F=f���OM<s�dR�I�P$.��v�:�c�ǁ1j�m��n�q�9�C�էb��jk�,�t��ߖ]�ܴ����D�B4�T]l��N1��r��1Bv�����y������w��hJ�H���ǵ��o&�W2���)��
v�|:�E�p�a�\Ɨ�NtJ�h��^�
���S7��ǻy���1�����x5�M���[�\���%����޷9�'�/(Ov�,�*Am	c�	ʍ��3���{e�wYڜ��А�j��>Ժ�F�0֬ʱ:qh�d�lգqV��(�y��]Yʶ���#V�7�Um�#��&%��h��Ek�v�c��a�P��(ӱ\��׳�����J+s��4��"��R�d�]ZF�y�n;ޕ%�����ÍTI�uҥ�ܝO:5����Ǩc����n��3]mrƋō�9^��0�'�c��o�k/%�1=z��y���O��*�*��b��g+c\�.20l����'��k�ԓ��Y6�otR���E�[oi)@ʼ����K��/�Q���Rw��	������9R~�`���o��0#*�Fb���T�_�����u%Ka����i���:���u�)Х�mYx���}�5��mA�Y�û�{r�sf��pOLo�.��7�G֍v~��I���o4:-�hL���g��}I���܌��$wJ�<u'_H��ԗXNZ`��]�V������u'���T�a�����؊�7�͇�9�!/Gٱ���]��F�35msZ��,;5�-�Nc�ܛ� D�Ǳ������c]W��-���}g�LFjp���,��p�+�ltEE��`V����: �1�آ�Ќ�$���]�ifV���L�]�[er�C�+#ܔl5Ҵ����7�5�h-c^��,j+F-Et�ԙ��A��{;�s�`����oQL8,-=�1b]�]jk`�Om��U��9�����k��ꕒ|1]�<����WW"hX�Kv�Εj�9���˾ݫ��I-=�;U��E,����[W�#���W�
+���2�T��[`U��U_L��O�앉�N��{�aI �4`�#��."b����-�wn��L�`��J(�d�\h����$� Ƌb�G8�Bf�LX�IK����#fb4����1�*f�wt	�,b�ɑ�u&wtыW.b��e��L�١E,��5�b�32��D�1n�v"��k��d�h9� &��g8j%�)4H�jBF�ͨ���s\�&�)#Q�6�-"���]�QbҖ`�WE�( ���1
"�);�e�t̃HlE$b�J��]ݤ�����JS Ԙ��I�W$�n��w�˚3;�ц`�Ƀ.딌4�!�wp�':�!%$T�`a��$n�\e2u�Ww2�5��@��4*�� ̸@U��}�����L����nr�N��J$]K����+;��!���[�9�.R�wM��"Bv��88��-R�]��]�N7���7�Ys�Z�!�4n,���[^���1��1�9���f��;<J5oTWG)�g��}9�D{Ʈ���&K��Ј^L`q5�뇐������b�'�%h�y{�<S*gao�3k:��F9�S��IÛ3tzԴpWˤ?Ma�2)z`��~̬uw�~�����;���m:l�>N�7o�h���]-7F�ݣ>��0�%�񧾟ul emW?-�{ou�ʄĜq�A���@
/���-��׃��Y����#��_��Y�@����^�Î�Ec�$֗�<;�1H��a}V3��7��v�7\��ïᶧ����ʌ�˚�$�7�I�@Ӡ�;~�Wq�ixs7]0/�M��9�q���<�3��b�C�k۳=�Iw7�B�*����隉US�H_�W�Z��U�v�Ӭ�Zz�X��f:4��-�����@��n�"�eqq͂�GA<HQ�@@�:&���:;t��Mi��ūn���r�+{��u�79��6�'i�S(W$��x��P$�|�P��N��Or\��ې�Џq~k�q<E���eŵ�+���@�S��,�yyYv[
�+Ks~�(Sc��2k��y��7�^z�s�%ֿ��n��K�r���S.^	Y���L*6�V�X�!o�<�����re��V��k�P2:�L���h���%�s���: ��,�C��&��}��B����צH�P��ݙ���@��LH���m�\ϔn�E��{%TFK�yH��=�t�}���w���?eįY���q�tn߫�줤���f4vo��0�C���.[l���c�}Θ_"�~j~�?z���f��V�E�Bx\�(��v������߼�o��h��B��}ʣ]���y	��+ڤ[������A�Pnxz�N����S�N�>eF]]G�e����ag�=�{I�����s,N��ߩ�M2��ě�ٟ��d��S���ӄ�2�<Lp�����^}ޙ+��o�:g���5�_��3�ֶ�z�TΊ�'v��;Qsǁi{�5��q�ԍN]�p��c.�բ���Ҧk�Nԉ����D�2}ΖǼvR��N��((��-P��p�Q����).8�.+���W��Q<.
�;��� ������֝xh�o���:�5n1&�����oZ�I���]h�C���^B�q)����� d_�x�qΡ�L���Iy>��#�Z����_�³�6�}�]�v����>��.�_��>{^e�Z�ma$�KV�|���R��tAΧ��O�kw`Gw2v�6�qѾ"�J�p��E*Sű죚]L�4�Ӵ��7��[N�&ŏ�k��e�]eD�rR��w4R�B.�7[ğ���1m��eB��隈�#��%QU�Lt[���s������\�Ƕ�Ǣ�9��9;\����yc.�l��5� �:&�R�~���. �%��s/��f[�o8��\�	q-�.�]㑮F��ꃔ�S0�M��@ݦt�:?����ۆ�-�:�r��C�bg����V��k�=��&�:��Q��G9R�qMs[�U�v	�'k��J�48=h >�1��m��^���˵���gۜ�:�����r���H���/IuMO�xP~(���3bj�.�5M�mxpʰ�n���U״�f���8�v��+n���}3$�H�%��F����P�j�Q7�v(ϭc�Pi׷#}`���J/�P��`�օ���Xk�pjX�@ٰ���a�<�$�xO�Ff�?<�ym+Q�g.�o��t�Tv8\�7.�5"�5���I�1�P1`�/ r�7/���_��Z<�q�ы.�ǅ�o�z��jz-�1]��px_�۶pg� 4�9Q�(l\dYq���B1�Nt��= Tum!S��Bp�b�L:�Hl�)���s+�M��C�ƕ�
�D��i��P��=8&��e���&�v��������n"��.|��Bٽl����R&j��w��S��:;Hj�P��-Ž��"�>�I����9G�#^�U�;Y/ʌ\Yu����V�qܟ��k��o����v�ݒ�\��Q/^�̤��xu��Q���<��F. M����Iy�|�ޜ��x{C0k��>҂.�w�q>��j	�w�X���-'F��7d�����z�=��<�[�ȼNNo6s0�oo>�WU�z/�;����a
T^PA\U9���U�u-UFϡ�뚃��l��y������8܏E�9l�_�<�Y�M�i�n+�d"+Ҍ�A���T�Z΢�gX��99�/j���y��(�~�u҃����8i��o����;�v}�BDp��a 3�swO��o'���p8S/M|�X��"���X.<�_�hq�x�'7N��i�x����lp*�Z���R��������@(��ҙ��Q[���{�~z���m�j�DbЎ�����v�/E%~��}���_�L��f$����ȉ�|.뇑O�؟�ث���:�Mi��_�BPn���jwЬ߁��&��F�U3�+�I�4����__���J�:=�u�V{�%�/�h���LKD����ܕ{���H�%���j�aeP�Һ[�{�X>7�V=�"��u\�n�E��k��W"G�y	w:�&������;2�!����49��2h��
]��Z�3���z�����\ �[�l���p{�8�����=l�DsV���NMG�H�F����(W˧�S�odK�0��^C�`���L�~�U#�h�����@Q�i�^���;FF�[�����T��Nox��x��*�2X��X���+���k�偮�Bî.`g�ѓ�~4�F���o��O�8���c)yf̞.�.�j�o��ʨ��t��9Cn��pmL5�R޿%dс��� �#%!ctó��.z�>eDe���<�z}�@�r��xJ�n�edm�C�B��&��V=�F��AÕ��''R���>d���2��GJp;�*�Ӿ����X>�����6�f�,g���N���GN��E���m�b|�����߬,ܷz�
���B��@�]�"]x�ß��q��u�,'���%p)��W;���^�F{�+Ӻ�)��\\+���d��Tau +�y�	Կp|T��B.#�{t�E� O��<��2�j֒�,�-
e��Σ�V�b�:'��Ƙ~����r���w�&�L������J�$
�-��X��t�L1��?X���1�2R"ȴV���xej�\�W��j_=[p�'�]Hm�u|�y�jf�
cC��3�ᕝ�vr�r�0q4s^���
e�n%��sW5-�|���*u3Q��+�<��́��z����R�K�8I�f6�~Q�qϔ��q�AW�Sf��};�@�5]MDꮝ��:;�Y�o��v�.yJhS��c�%�ŢG�3_JF�SbȤ�[{qA��O%�zc��s�>=��\VA�h�N���h�؄�q����Y���� lwLM�H��Rr$>yW<��Ӷ�/E�E��-�f,���-��|��NӪ�P�IO�A���|�P�f�mC�u��5�ڋ��B����.��\B~�.r~�͹��i�Q��P�zS�^�#�C!�nym���NO�9T�/�|�UFO�ީ+�ΐ��ľfX��5��=�-[F��]�����
��(I�#A'0�;J�X��f��u��k�wr�k�ɂ��3½.�n��+1�Ѱ���u�j��3��A��4|�����;C�~�yp��v����Nl�
�(��.���;:�Eg����{�{�߫Z3Uȃ��W��.p^)�'G�|ɬ!f*��-�8��1S�?��~1��u�s<'\~�H/��S7�I���&!�����Շ\{�jJ��Q"Ok�KŽw�32�
z�톺���Q�+;�MN�V�ՁmB�ܡm�'�,�(q�"�S��~增���E�"���	齪ՋOց����u����t��qjZ� �*'��C�wm&��Z�-�RBh��م��7+n�M�#�nj��9�Ȩ�����_kw���u�o\�w���cZVs��Iݸ3���7U�����!l�5e������������I�O�#�;)��*n7Ϭ�W]xR�7캌��9�I9'1��� ���ɥ�_.��X�y �}����i����F��9��-�ՔK���q�C��A?�ڐ�.�A�#�A�.q)�Ҳ]L֑���1f-�2���f3��e��r��̩����7����H�隟#�RU^��[��V4�mz�3w���矇�=O�\wHg��9u�P�ǖ2�Z�����r�]��UF�ߋ��r������	9�]�ˊ�MO:c���q�g+�A���8�h�� �lA��s3��5C���S���(gH���\ƫ�*'���g�׆�kt��玢t�:��U�s�,�q�֤���o��Ӿ�4����$
{P�a�;v��#�{�W��k-�b��m�2��\ז�(wyj�\�A��Ě�)���E��n�MC�1���i���x��85sY%��+3*�
Y��__�y�D���T�S��}l�q��AA�w��񷷮��1>=^T.��aY�$�������l��G=�R��Yp����K+J[Q>�#+R��!+̜e�Ç��׋@͊V�u��/�p��Ǜ��9�i��moΝQ�JfΉ�J���)e�E�3����T���AOjaT)~8����ʎ�/�6�l�]�}W�<'��E�d�\�_	�25�d/5a�M��=_�
z}���">�E�>9�!��y�^�}8"���eﺩ����n\�jE�0���3��'N�~���>p#]B�|����{F��d�����3|��/���\g�خ�~�</�^ݳ�>��Sթ�v<Q\���7��艬�gB˭���.e�\6<�V�w'�7��AϧNK�m���ޯw�"I5^3�����!XsU���G̟V. M����䗙�ޙ�ū۾%��w;���,ע�B}���t�ϓ<OdUf	P��'EK��v0�(����:MS�5���׼ȫ���<��vy����±��|���1�����r���=�~������u�~���x9G��+�ţ|����\{��Ρ{��W�Z�!��FE �dl��:�,䇯ћ���|%9�7^�;�K�,^8k�_����T=7�C����0hRG�ʷ�L�خ)'z؃*r\X�W(�p�<ұ�Q�]�%�Gr��g1m	lm�#�L�Ÿ��}`�3���Z=~�Q�&<B/��wl�pTM�x4�4
��
[FoDOP��ZtYy& ��e���E��b����6%�ԙ��1��wE�\��}�>�lt٪LPW�>��fEOs�p_�#�<^���P��.s���s�b�)�L���'Ç����0*6�y�s�iL�a���Q5=޿�=i��6��/��#�.�X�8>�Y�S��ۚ�H�ulL�tb��ى3����}����S��63�_����P��ޡ�h'6s��N,��:���2��RxzI�N� l��^
���2��:0��ɹ�m_o��*-�m�|l�~%�s7��`dsV���NO�#��U���(N�>sT�}YU|6_Dؖ�N#�YQ�����b�=��C�p1�Ϲ�fd����)~Q�]3�f|�ԇcRU�ބ�&��`��Kª2X��X����
�Ƈ)l�1��B�Q�1@�6�5���}�p/<��hQ$�P�"/=[�=P��5�����W\/|�x�kA�߯�Y�(�y�����ޠe8%g���u"�|�>�a���1GM˳������V]mp��I�yY���NL\	Qn�?]Fm�����'o;oG;X�[�AÕ�~#�ii��M��=b"�)��A��˪��%�^��@�4�!�m�r���U�
�5d��5gxed��s۰��%WN�4��F�D���5�ܣ���@����iXk3O_E8���Z��\�㸳h"���nofx���k
lG�
��Y�7�b'(�Y���j��[?W�W���𿧚�7���Z�3V�F�7��ۙb�@���7'�;�U��dWV�W���X)��G�7�����`{��ϥҌ�������(e�+�;ݎ/r���u������ex������A��T ���l,��l��^n ��o�O����ܟ3ԯKl�}�����LR���' {�1H��ʆ�tO3��0�i����in�����:7�}79uH{�H����FHr��
��}��k�ou�G�!��R��gʉ�5ܼ6�e0�MI�� {�D�Q)}M��)�[{qK&��F�������n�)j��>�|wK��N�n�ʄ�q���t�ā��00�|�3Ʃ4��1��I�:p3%�5��k��u��[s�M<u��P陞9�-���6���X�d�MZ1���i��ʔ��9q�<<��mH�s\8qo�Y�s7��6�6D5n�TOJbb"{G^�E{��ݵ ��~� (�s_3l���UyFw]J�I���<�b���#3�菾��m�����m���mk[o�umk[n֭Z��kj�_�kZ��Vֵ����ֵ���[Z����[Z����[Z���m[Z���������[Z�۵mk[o�Vֵ�����km������5mk[o���ֶ��kZ��Vֵ��յ�m��1AY&SY*�O� �PY�`P��3'� bA����R���Q@TD�%�)���*�"���B"��(T�JB��Q �I�%QUH�%R� @�P�B
 �U UD@�UP� ���JT�*�-�	J�
H�z5%"��*��v:�U@�(B�QR*!���" �ER*�*��BT�QR�!T�")
*�J*UU(
�BOZ��$D��5%R"�AU({
U(��  /D�����C�ltu]�;uFڲf�Z���+`�B���b�C��Z�Z�Ԙul�+uWnm�4�ڒ�)EP���H�� ��:�ڨmt���[���A�(�Ը� ��(��wOoQEQEq��P���(���PP �wE�Q (���8�(��( �ˀ��(�tvT�*U@TR�*!I� ��V�ۨM:Qn�겂n��jmJ���t)�V�L uT�+��u�m��7 uvmvS��.�ۄu7[j[9Ն�AE"T�( ��w���M�v�Wv�Y�U��[[����SZ�f�\�1��n��\3]���n��Jܕr�ln��T�ۺ�Ӯ.�wf�N�V�.Q�T�eln�Ѷܵ�5��jH�J���*)4�� ���hó����:�v[ln]U�U�I�V�r��ۻ��f�v��ۻ�m��k�ju�[N�6��u���(��]�ַg4���N�,����v�U���:�*UT���D�J^  w[ݪ���;�n�6�5m���v7N���W:N]m�Neݸ�K����v�ή-u���]u�ݧJ�v��حԖ�ְ�s��5���*���n�\�R��$����(�^   ��s�u���+:���Z�ְ�;��۵����hf��]���9�;m�W[n�[mMihk��v��mw.�&��[����ݫn��FS��M�6�s�v�%���(ֶ˶H%u��  w�[=�ۗvwSe�5V��5n�nӲ�q�n�Um�k���]��f��Lf��ݭ�Ӷ��]uݎ������]ksuw	�*���\�u����e��]�""�H�*\���D��  ���N��uN�Y�r���̇p����9�s�-n��˥�mە��ێgR��t��]5ջJ�wB���tݲ�]�wv��5r�f����mJk�;b!T���P�O  n�Z�][p��w]ۢ��vt��;��mv+�n큭T�U�Su�U�QS����v��s�wv���K�p�+�u�]�U��w	���Q��OCC*RP Oh�JTPѠ 2bi��4�E?�)�  T�����M4  RD�U$��2hl�������_�?DF~����O��ټA��6���^���~��ík߼���AQw�� ���QS� ��������+�@* � (�����_�?��ٞw�`C�Vq�n�3	DI�BY���z�H��.�K���kY{!��N���4�:ւ�+Q�Ď�]���)4�x%"u+!�?�kK�M�{XB�GT͢6鵩��Nօf��� ���h��f\���V�R�h+�֤�W��{����&���8@:�)�ػ۷���A`����I�oeA�ƖM(鶮�GIڬ��˥��틣���Ԭ��:4X����6հ�����MX'�1����qҟK��`��2_���=�E
*IrɀՄ��e]f��"�n��D�c��A��̽6��o%n����h��M��Y�	���"+R5�.��
��u#��fe�O�n[y��X�Գ���u�NI����u)Q��ni.�&,�*�c9OiK�c�UӬ�r���ckf8�TOn�]��w*[ּ���-C��n�ܩAYkn���-B5�E*.O�
�<u�1�h[�/�qE�RL��n��S��PD�
ʱ���Խ��Dl��s�O [�Y{qi�ޗ{�`�X)X�T���Vܵ����J��Į�=��X6�џR�! �JJ�7p����]�*�q��DN[�`�b��PQ#��1��yY/.B����3-hV��ڬ��y���j;ba��V�z.�C��7K7j[/
ԫ�a:�Cԧ�R�S�8�P���ǬL�#�Q���+
m�$�f�sM�u�5�*�jt�jұl�X�*��2De=-+��6>�R�]���z��Gf�J��v�(�4�O�4no1)� �@~�ҎΚIk�Hlt�% ������t���鍤ZbL�X&G��+b�PI�ktmހ��V֌۔���1��P��;���Y��ikT-IEeln	��E&�W�;�yZ��*5x��$�z݊	E��՚o�`�C�f��jeI�-�˷���_d��ܭ���q?�99;K�+ �BR���F]]�pM�NB�[_n�Y��-�3�NyE��6 2ص��<�dMtl����`��Wr�t�6�T��".��D
-F\3�B�ؒf��VF�]P���"7��wB�]bb��0�q���p'w��i�^
J��4������ڽU�+k��2���IX�V&ܴ��ݤ�yU�M&1Q��\ʸ�bR^���k_M\.,#���YW����#X�wͨlU��Q6�KN�͢����r_=w�hM�n-1�����Vj� ť��f�Bv]
��wkZ�n�����C%�^�NK:�Na43�30���llŬ$۩u�KB��lFM��#,� ޥPb@e�+s���=вZ�I��jY�����H{u�F������E$����9)TET��"�%���򴺟IN�υ'u5TS�(ш�����U���ڢ��ըn�ۭ�3X��â�:�+A%]��՚#�ŀ:i�Um�j�%��EI[bQ`�ً#��&J����Qi"��Kn˧rn�,�U$.�r�ʷ�[瓟�
�(�����y���-E�����[Ms^GV�Dڒ�sKv݋hr�!��S����R�p�zud�5���]��zޙG6�eӠ����i� W���V6��g"x�5���&O����{��n`�ƥ�̠�˙��4,��4P�B���U�l1��� �w��͟Z��R=Dr!�i�FQ�h��fX��`�әuw�2� �C;���	Z������m�m��ܭ��y̛����S	nMW2�VJ�at�Ÿ��m�S�)��'�	��k�v�!CG.Ҳ7��o�5��ֺ5���[h�,c���@n����5��D�RQ�vF
���aSZ�Fh]H�͍��G���Y���2/`J�r�M�r��	nL�WC["U��n�hđYXK��v�f��ت��rT(n`�H/$�B�b��5��i�;/@H8�1<��e�x�chG�5��|��Y�n��q깩��gVlDַ���V`p)��Y2;[���"��T��&�H�������趥;"��4k�%n�椵�b�Kq��pbV�p,B�ytRZ��v�c(}r�e�:��oGt��5-l-D����w1]U�0V�aJ?]^V4L����Ѻ�� 
?�:�e[j�H1m-;�,��2��(+`ܦ�%�;���c/k&�Y�t�
�V݈Pυŀ%{NP� P����+�T//�mJҢ��=���Kk�IT����;���T#�&V���(�(=VD���,�QT��בܕ���`'f�8\"�+�D�m�W��{I��	J�C��x������(��J���F�+D�f�*��lJ�n�j�#6-�*�C��=�MimT�X�B���ml�h�C<���K�J�2��n�Kiá&bI����uMxi4�A��Fo-UJ �ec͘�@cW7,T�F�Cm�E����)��z;�-a��]eX�ZD�l��5MWx�:��^@�۳n��d�%�e���^���?�n�.ٵyٗ�)Vݥ�p �"j��3C(ѵea��a蒸�:��EZ��[x���"�(FX�B�-!Y��c(�7b�L�MS����V0�v'�^�z���Yyc	��)Z)��J�ڽ�tF	f��m�kN�r٭�2"��̠��Ю�KFS��U�nXMg�+e]����,Pl�$��ny%�3�u�7(���^C.ٚ@^X�mn5v�mGX�(���A�a��f�	v��òDВ5�����aLYu�bă���`wR�v�m0�[g.65��S4\8���АӶ���K^.�7Ebm�V]⥚�0@v��Y�m�aV嬐�X�/`XpR���ݸi V�qH��!�[��r�-X���T�����P�Ød��Cj �
ac[J��efԚ�#$wn4�	�o,�6VȵD�����C%��B���㙺d����b�7F`[{p�J��6��{S��L�)�Q�N��r�����Mvh�4���ܽɆ�Tר���D�Ub\;�*	cv�����9���wL�д�寂zٸ��-������-cOTV��D�D���߲,�eTȒ3iZ��vv�[�����4�ڱYUw0��ĺ�n�V��'�4p@�-��d+�V]w�͝&[�Ͷf��l67�
%�nŃ��X�b2��mL�V*F�^�v�z�Ej�b5$��OFϵ�J�Lͬ��*N��r�T��H���x�%��r�HŚ�&8&)��N����(�r��:�!t@b��Yi�9p�[x��EdF2��[�#^�Q�)��ɣ��{.֡iP± ���
��e;�%r��ǆTP�X�I��l�V�LH�W`4thǙJ�K�n�;eR��XCI �
�j÷���f9�J"�����GJ�`��$���T��L�V�i�qA�E[��"K�]��Ld�K�WQb:�K7 ���I0ؼ�Zt�\W6�
��$LJ�&�ͼ�b���-K���mZ��Y���,���&��*V譈S��yz&��ѐ7�mZ�JXjXϭjPn�rd[vQ+@42��q<�L��.Kw����]��R)�b,v"���yX�eӱ�Kq&��ܬHY���J"��˥�!`e"T�6j҂����P�ͺ�X�R���!򁭑kcI��旮�i�5�.櫒����Ě��J�v�ֻ��ٌ���F����+o�P�F��9�A�!)Ca�%�͘XL�I�h��E�[�)�7,���hb�d�0�m�tVSk��x����T���Ȱ�{[�V�9���+Fd����J5W�����.��3-f=o-:"�5.��OD����Y.�;�VƀYYX����7-c�Ks�E�mnS�Q�U��X��q%��uʁ_؍�+n�E�(��h;e���I�0�:��[�U�# �mXi<0H�`5+/i0q`�r�3%#v�ДW��n��T�i6������b��I�]M	��M��t66�/�#�kn1@غ�*e #��N�Z��B����T>8.I�f@�`�r����pZ2ځ_-��f��,6�G,�X�Z��驆,Ҿ��ں 9���Cf�Js�V�bP����%��y�2f͢�KT4�TݘlM�Z��O���&nMg���R5tIo,34l��(�*���K	бwNm^pe:7*��&���=�5�2���R���*5r�[Aj,�"E�,\G�ɫ5���-e�`5>+PX�(	%n8I`��iF ��#N��.�A�Ćc0\��Xmn��Q�E���M�7�㖪���=f���m^��B�=�،eǛ�1�T���LP[��Z:�Aj��#+p`P��Jx
Ů��!%=�w�)J�Hh�v ��Kk2�[NQ�9��F5i���NSs%�A9�wFCϢ��ˣ��m!N9�X��]a-��A��l-VpSE'��ܭyBɡ�M��kk�m���w��(�v�Xq�MMڤ�7w���9P\�
kv����2l)��� �ޣB�=�7!��Bp��k5=�훁-yf<�I�p^mxeT�Z��7GiM�Ɇ�J���r&����<���\Or++Idؔ.�)ch����M;yB�IFH(0�MH�H�7�[9Bɭ��dn9��Q�1:4U�-���h`c2��h��JZ�7�.Q14D�2�:�/VL��#N��2�7˘���3)l�)�]Z���V5ͅ'f哛�E*N��P�p2�J��jU-��jd8�2�++E�(�G�*��0b��7�cٳ	ݡ��k\+d�E=��c�E�� m*�i�h�����Kp���M-`$�4=5�P�G;��;�oq�x���5V�1�MD��V:w��Ĭ���з�B�q���%�[�9a�`l�m2c���6m�)G-V+oZx>Ԧ��5�\q��3�B�l{@nfJ�7�����x��5sUm(@���Bc*`vv'Y{l��2'y!Z%mcxk"�ɚ�d�Y���%��m�	��̍V�$f�\��`W7j�r���%C��]˘
�%Vf}�w)-�9��F���#Xyy�$���+�[�bP���a-806�]f�wh�i-$�܆Bq�VeA2����7F�9���� 2��ʼWC�Mn�X�U޸�c���S[Ԛ�[��n���Yu�j�L���F,��+2u� P�k�&�
�IFk1�Z�4��m�%��-9>�p%�+����uj�=e��Y��*6��l`�h'�W�[��oC���V�j[��]ec���u�%NE3#������\��B)��k�N��\�cj�`��a���3
9�$���l��˧v�:^36j�VV�f=�ddomֆD��j˫��)]V�P/pBH�8iE��	�FH���+-��r�����˳t���I)r���r�aQ8Y��6�<�n�M��!M{cȓ��ԓ`WZl�u��@��e��v���򍴁Ͳc�R�ȱÆRC,ᰋ�@-��0�nR̒��(J��)���e�v�چ�`�bPutc߭�ۛk5�
U	T�܃v�tQ�a�K-U�b_�2S� ��(�WYMI�N�a3��4���S%]�=u��F�mُS�H��ϛ-�)LT.)�Ǖ��6��ڻ����0[sYıCh�`�(�"u:�*����VLV=&��ֈ�Y@�ITI��kPL���n��QP��[�0 ��q4�^&�l��S�i�j�ј�-#kU+�	�Um�]�R�Oi�wF�5$n����x�6&p�/j`2$�d��q�1�+譿��1��4j�ӬpK0�Ӡ���d�;��Zc�(�
pݽ�Q�WJ�m��"���-��37-�O�ٗeU�L4&��f��b����͠4��T˖�[��{����ѵ�L�"��ؼ&�,��M�V0�Q�����Z1��noN�[��Q� ��[6�;M� �¡VV�Z�عb��G�����]+���\�qV�m@�<&��;Ux�-l��qFՍ�Z%m%1�+6��+u;���j1��Z[����yFؕ��#SD�z&��0�nhJ]��J���FJ
I��Ҏ�O�y[�L	9�,L�7�	qh�Xq̗�,%cŃ^5�����h�3n�`��-�Z�į�u�w�mpй{���u��_�SWN�d���Jq&Z&٪�WZ��IMH�7L�A�f��"Jbkf��2%q��j�x�h)�	N���Ǆ=7�:���ۊ�i��Ҍ�6ڹ�����z�O\�l��C�
�6M+�s౥Fka��v^���֛����e��Y��\!�|6�_K�kb��H)Q�Y���WPpA��jS�~˳J�)b��m����y*l�a�(�9,�W���F�k��i,vd�[x.�&���o�P=�������x�+L�
ƼF��aT>�&V�Ӹ�����E1��(m�~����-Y�R���f��bb"�Xp������赚�jz���[w��J�7�U��*��>�&��Ȭ���yz�e2�(aux�Q�09[>��8��f�Y7q���MM!B�k��.�U� �a'
7.�ڔ��ޢ2,l\+54��Hi��%����JwV��ne����,qC�	vٖ���C��	ѡ���[�����Ջuj��"�@�2*f���7*�b*5�daZ�W��ci��-e�ib���4�$��S(�-�2�,ù�9��4e�[(2q� �T�KJ��Q�>;�V�JA�	���au>�$��u�1e�B���[˩�)<���-9������u�5�awX��vh������2��kI�fإ#��r�U�]��OY��A����s�����P���I`]Y�y�(*�z�kUs-�.6��z�h�2󦭵>�u�4�����Tr���A���mܔ8}9�-���!��l�Bz���`��#;m	���wJ�ŏh�k��7{J.˫��ZtN�׽{Y!*�J\�g}���IL�[E4u[�]K��t����n!@'K��z���@!EW$�	E������*�����d�Q<A�д]��4x�f�f"�4��i^u�E�Wy	ot\}W�qv�4�Wok2�롽��"�g-��.��>ټ��;ҋ�6��{Js�8n�v�� kRm"0
��������Ž-�|h|�OZ�h1S�O(nYY��+�D�gv5]{�U0�L��XK����V�<��V�CO-#�c&��w�GYK�TT�[�nI�&�f��ղѓu���Om.����9�[n��)7N��#�'2#BVj��r���aM��fV��V�N��k2h:�9N�a)hj�]s�3��Y�� GV�6,��]�7M�HL�����������Vi�քu��r
�����w���K�ơ�MI&�]5PY��O(z�
o[LR�]�a	�B��0�u�n��5Ƶ�b��"�@�:�ݘh=�fM(�������Y",���X��!+Ec�P�܇S�-�om�wK��.�<H��yr�#>�/\���0��`!��}B�Q���F��gd�'
P��`�Z��x��]O�J?1���W5]J�N�oE��	ږV���g��f�GN�]r�B�;����Q�yz�s.�"�I��X��iڵ@�X�4�F�}Yvd��j���V�������Gq*�$w��� ��t�\�:yͩG��ڭ���ut]-:���Ӗ�KH4k��V]	G�]]ܲ^VhVsTŃV���eF+�+h���b��t�z��6<�W�IV��쉲3
�����!V�Ӂ�QuY�c^[��>}Ԗ;#\lN�m��M5u��T�TW��f�Ċ�R�V:�6�长^Ҿё�)Xw+
 m���	Q�|aV1��D�m��9��(P�/μF��5��rm6i�*����]9�� ���U�}�ҋ7��c `\��S���|V�L`�����xѧ1�;�aR���8�������.�U�Q�:p��B-S`��Tn�GWC�l{�:��]h��1i�"�"#1Rp�Ww(�Ɇ�D��-muD���V�oU�9�ސ��»-�̮���"2M�f]��������ͩK��ҺN.E�x�
��\aV� ��ߴë��I�2��=/�wq�}�N�sI�7"�v�r)���u����l��x\�A�>��,��.{:�s���M�+���8u��x��p��ݲ�ii	A�J5�-)\��: ��+@�{ՕHu�}x�p1�4C�_]$�%��Е�R�/�q��(�v%�{���#s[�6#QT��oW3*��2}��7������z�iR���%{z۬b�Rn%C,���2��՞H�~��ڗ��h�'B�W�KWZ�ՠ�;�B���}-�i�v�no�
�{օo.�`�ˈz��� kpt��:�,�]���$\c�T�+�{r��PJ�S���*����.H6א(���4{GE��eee:P�﮶:	�C�2�{4�t�]�@��3�U���&�[t�����Y�&7n�kխ�M.��yyv�ץ� ���t]#F+33�t�+�GyKκ��v��a�V|���E���� /-���8�KH]���l`��0~�8p{
.:�:�8��v�kޑ���D�+�y�r�]p�AEs����Ju=������X���;E6�y9�6�=L�z�ɮ��Wlw�,��wit�f���k���4siT���Ov���M`�8����>����&:�O���ݤ�ET'1�l��5�X���
��#a��qnu���R��5ӈ���u��j���wBPӈ�A� ӎ+�);秚���Z�4Xg�9�B�r{ >�G�ǘe�خ��q��!�v�K&Y���޲�/IW��l�v�}���Uq��Ͱ�%�Ƨ�4�fUq�\�"������/�
�!�/�ږApӜ%���k�j�h+ªY���p�<�4\3n�)�c7��Z���э��r�s���g(�KU��Qw�BU��˨��C|h��"{*v}4�҇�2���R��*��V���h�6�Q��h�U����|�K���`��|��'#T��Ɋ�9eL�0h�ZHe�WRZsb�1;p��mX��؏*";���ǻ�D=�N��u�����j'�n�E���Ȼ�%o �j���O8�β�m.�p���}uز�}�wGP�w�}�m�h�0Jاؓ�����1W��R�Ӫ�N|y�?</Ef֚ν�p�+pc�(�m�^]M\*f®��oR�X955橘veO����dZ�"�]c�u��
�n���e�1i��_Z��f�52���4.���[j�3	�lm��tq�I�T�һ4�u����t�=v��T���Q�у@iIn�kl���j�t6��Pl��r���K$�\p�hw3�mAol���ƅ�}�̥;P��w!S�����a��#�X-���iU��h��*Ɯ/F��@NR�����/F��I��C��Y	#�gt�o&���>ﯞ��ĸn�I�Bc�.�H!W`͉\��%'6��ݫ�ڝ�Q�;EŬ�gh^n�C�L���7���C�ɓa<]7U��R�pηTU�S���u�@�#���KY�\��D�vo��7-��%O9ʶ~�)��r�.�8!���vٹ6��U�2�u�զ��2��uM��n"�����e���C8�RAH�;<�VC�W;�IV��}Ǯ�}�F:�07(�һ��Ɋ��=@��[+jE����-\1v0�vΥ�2hiި�2���vU�dro��.Q��sV�#z�\��x>5b�L�\f�ʺ��]{r���F�����)�b:�`�����`�5���ʾ�O
}-ܫJ�ӯ�\�O��l��-��=�y]ې6���^� ]b�]81vr��4qJ�2��H�w����֫F�K=h<'C=c+S�R���Kz��ҳ}S)�i�����.F�ڴ7@�jP��Ս��W�=N՛�4S�FR:�D��k����w;z�+\�-�ku��t����Lo(oc�|�&�:ħv=��RAV�iz�Y^1���ҏ;M1E�]�j���*�/b�n �0(^]>�cG�>�ӎ��r�Z�h�|M�ݗ�y5r�-�W�eJ�x����Dv��w/ZWu��vs9��̖N����`0u�g��}N0��67��tkw2�ǽYWQ�ڔD��%�k�������g��z3�*��rt(+b��n@��5��, +�}ս�n���wzby�}��J�p��l䭂'���V{�>'a��V�����nK�N��&/u��9|:V�����C7����gN�1su@���������d�2�i���3rz��,K��� �t7���+�3���	�v�E&�F����}3>f���]g4o�<���,�:-�+�i��`��코xT=�98����7��klP�����M�� �vVs�E�>�Ԧw,]y
��5���('N_j7��]Y�I�}(1Aug���|N�o�x+Nn��f%Pq��B�C�~���r�|��21`��³�#n��9Am���w���j�\���[���e'W2�'Fjې��/s��JK���͔�]b���א�Z�D)f5��[;4�q
)���gh1�˼,��Q�71)\����G(���}�={mRӔeK���*�gO�]�#�KL��bKp��M����J�"|2��ȭf����/��6ه)�NUܹ�Ɛ�'�:V����+��s��bN�V2p��3%%s��BLwvn�<��'�5�w;Pi��ay��'j��O�-�[�RU6���a��z��We�o�c�v��.�:$]���w9���/qh7�\G�JάVon!���j��:P�"�j�.'U����_9�.�������� 0��5m!��t�j�v�YM����6����F��r���*��oj�V�Қ]7��5C���@C��(�Ÿ$4�a����<6�Lbd!��؏|r�v�X�Amg$�U���:a��FF\�����DZWy�e���Q���ɣ�[g6��%ወ�j�(��<j't�kxn4M���K܄r�.&�HdU�'d�qXfvP<�E.����'Et5R�5V*�5θnTYO����qg�.�����e]��h�vS��Y�V3���������Eo8�)�lif��-�A�Z��p
�Eԫ�
���d���B� pܧ��Q��L�/gpI�[/�����Y]�аU��ǘk(�d�G�u	6Vn�c�ܧ�8����u$��ڔ�Bud977����݊�)Y�z*�Z4T��QۇM;��poיI�
�7�<�����Lr}�m:e�Ӕ�����N��]�^Q7d�!;�	�s7�?)x!O'hͭ2�G�L�
f�H�D�]�,k��Q"���۽�m̸����CƗ{-tg�X��c� �K���YF�n�9K�MT܊���w)��R�L#[�V��N���k��:�v��/�  ��;T���`j�m�]�Y�x^�����Z���pO��ö���C���PIo�u���L�6S�l�x�s�U�W]w����G�I���lBT����^N�t��+F%8i�:�iɫ{hF��dYm=ur�L���x�2�<}g�h�v�Xh%r�o��n��\=�����pS�0�����4Qp>|hLQ_�8�k�Z���q��_k=[1^��$��}t�VY�y���{�q.U��1:�� �cr���r�f����=���3J�e��L,��[/.vhV<ɔ�*��2��u�ݘĻ#c�S�_GťD�������Xxg7��N���F�ZT���f+�+K���P��D���Q���^2.�+�~N�fºbh�;;8�����4���::�Ůf\��8=Bv�X��{�I���s����	�\ū���mBηح!Bd�ֺ��n+��jpH4���K��{2wW�Y���qY�VXK��j���-��,ݮG�T���2�w�N���{3FQ�]XJ�]���CsXY�U�l;�y�%)�R&�@\^W<�+���z��RV��7��#6x���p�ޠ�C�}��+u-6��:���3u"��UwԨ��r��E�r�o�6^ !�X2�A񽮮r�/m��9+�"���<���p��u���}��gl�]}D��A	u�X�nP�Iֹ�*�5QE�nO����i� :�"��+��4m�>[-��p��0�>}K�e�Ø����s���;�rT����s;�N�d�T��ּ���dGaH]��[f��;WV���<+��Ur�G���8/N�:�7��
=��-�\�U�0.��q}�8��� *��GC���O�p�^�Tk�4*��ۡ�΋~�$����9OI�%�v��]:��utwhE�W�(���WS��_ܱ"l���KCǠHr�w#}�xZn�t�k��u��7ib���]Yx-mr�\�}�����z�Wu]A�����F#{O:Mb��|��Qct�l�z��|��h��1)�k�Z�3�T|�
��淩CZ3�Hօgf�+�<Jf�F�9]7�(5u2d�:��O0�����r�\yכ�EQŊ���BR}�lY��� ����7h`�ވ}�qtj�;s��s���[�Fwf�R�GZD�r�:���V*o��u5�Yy&�l�u| �L>n��}[�$���s����g�yr�GN9@�m%�����O��,�x�v��w�.�S��R�Šۢ^r����ݥ;�oJ'��V�
��U��H�:�J���+��zs罣��9ĕ=�M�h�K�&"��w{��f�T�&�}iL��N�VN�`o�������|n�������K?���he���C�n����&c����8w"��Yq�ykq��,�NE�^��^��6�F��z[t���i|��*�x�b�����R敭o���nX�5i���]�t��'}7�������k��՚T�@����3�eo\�F�tЙ��+H��L-]��`V@���M":�RV��M���@�X�R� ^S���n�9Y-
d��b��[ʛ+��P�#�˧ǟ1ۘ��wI�ӷ�T�� �f��A`�#*2� �����]��N����>%�ܲ�9dVm��6�Q��F�	Q��tj���Z��R�{����;|b�)��sD����.��^.+mF�:��ڙ��q�2d0�X�Q��-i��φ��(���A*N�@0�E�)V�Jմ��͡}l�{eX���n��ꘪޙPV���
�Ns&�W��1���r!%��d����ۻ��;���$R�	8򰳧V��a����Y؜�&u��f�aa�q��;���r�Vu���������sE�s�ъ���}�얲{��ʹ��mp<A@�5-����f�{��@��v���p� p��ɲr�v��*�.��I�c��.q��mY�p��[��{�����`�S�	�u��׷�9�f���/sl<o�)��%�|N�ː���)X���XV�>��q-�:B�Dw_i��6�σ���84E��_L,��`�ܤ)9%�Yod:� kM�}�X�QśCJZ&�*��Z��ԧe$�#<����߳�~��>�����
)� �����)3B��	ee���o�=G�5:�om�DK��@���B������#'��]��C�:{���2k9[�Tn��`�nF*x�+)�����ŷ����Y��k��u��Xӧ|��VR�r0�=�W2����I%�÷���:��ģ˵���U�N6Y5�@��d���a�S�n�p�ֻo�R��#P�}�yn�M2�p-�:�T���2�(i�
�l��h�ZP*0��ew-ŝ���U��q� ���P��E�e��*R۹a���]�«p7�ݝC���(+W7h�Q�T��pˠź޻KP���*�-����]����+s�F�E�{��Y�ً6�fC���YMF7��ɘ��D6��y�s[	���PA������j��+R��r��F����w�7��cyT�͠�	�r�r�3B@�J�]�{���B@�D�H��D���6@���0<�n.��S��u���� E9j��`�΢�hq�v�Y�8��Z�:�?g3"b�e۽vͭ�w|M�N�7L��;u	��R��]�B���@W�`!	��U�*$�k��� �y�̹(�SN5
z
��+���*n�U��U|��mX��,,�3�wjb�5�꼇b�%䡱)K����֟���0�G��F��m8^u��􄘅�K8t��&�6���Z�(Dew[� 9�5�Ν��:]К�Š����,�M�Y*Ue��3N�ш���F��/+"��K���%6�sQ�Ղ�Mn�x���=U�V^d$$ȹsC[z%=š���{Aџ\��ʅ���ի����O[��m�#f�K��J����\<��=�6f0�w}�G`e�|7��3��A��,��3�I�Z4)�L�uAZ�6�l9�	;t�b�������1oJ,��G�-�P.�"ق��L�%Zq݀�V��,wZ(K�㵒�9u�B��2_*T�f 9W3�geЫ�'&i�V񹖉��#�]�U�fh�(%��1������Yt9T7}��Y m�P�JӺQ]Z�J_+}5��+���ݫz�r��������[��X��k-���}���;H%�s�.�����=�ܻڼoo(wf�7Juww#w�R�����&�Q-�X%I�wZ(+ZY����ˣR�
�6������S�������)��&^P&�)bT(㚒�%�OZ��DE����ད�2��Y��e'z\6��]�eu-����=;F'bˏN]<�4���/�d;G�_/��Vګ�$���І�d�^�����:�GxQ{XM�QT�CN
@j: dv���v�ut�*r��x��� �	16��wV �����;����YN���j��M���-����h�MU�FydЩ���^S�Ec���4�yF��<'�@�vn���u�����aȲۣ�L\V.��ft��vR���h������/]�SIqֶ0t-��+����1�DdW���S
�vT�>��%KH�� Z�
4�8�sO9ġ[����s�X�e�5���v}4b��P��͹��Ǝ��oI'sԅ�6���qؤ�H���4��᷽S�G�����C���4]f�f<&6oF�%��x�k�m Ɨΐ+�Rꓧ�u��\��p�X�>T`�-�w.uԂ$ۣzo��p��IN6Du&�I�ԅ[)J�A��3*�J+�p�ϫ��N���T�3��cQ��Z�)B���]�`�Ŧ�'ۂ������Q;��J9M��o����d��´%yq0���oǷ4�q�.�(_7�*�oWժ���v���%�n�9v��C�����2�6ʭ{W� x�w����d�ɱR��݂R`><�Jq�S��j��Z$�.�F8��D�I��S.�@d:�&�p�Ѫ���`Գ���W]\�)>����� .�8�
�:<�nj���B�����I�ܮ	K���6]��x�J��"�����
�˩;�Mk��1��;Ț�p���W�E��Jm�/3NSh"�P0Դ��hͱ�K2N�&���Q�&_vP �G�N��n[A�>�gy�q�'���xڭ��oS]�A�����HvV#��nu�p)�X2<ڀS�V%X���W��ٻ�o��0)A�R�R��,�b�����3C��;�M�G�ec|���lx�DX�8������M
Ö�ӑK��`���p����"F/*kOe���50�폯�T�Z�������c�&��"��-�Ҏ
���ST�5m
_n�scJ�O:q4�εP�]��3�J�<���j,w&�YIf�D�}:��Z��XMi�z�%�J��/�;\#ד� #�h�	ʰ� ���bW��1cK���n�J	��ȳ�fQNb^"�q׷c S������i���'����P���s9FMܠ����n��W�5u��"�����\y4V������Aύ�0K�f*�Rf��������R}ڠ�j�-9��!�F%��]x����JX���U����u#)&Nr}��l獥h]'ur���yN�X��v�7���P�+u�����T�"��`$W����<غ�V�]2%av9�������ū�����̠*�`�$�T�� 3v`��]]��:*��s7���i�ŐnR���3%2s����ԥ�g���y]F��%�T/�$��i*�F)���gd�U�c�b�,�Q��ZU`�������p��+)>�3��Yre2Nr�c�-��x5��`x���P�=u�d���D���k#�k�V���� bp�zp��քLl�Ԍ`I��̔aIt�5���8RY*��$qh5�C�Q �1���&�n�P�X.r��':�H٨v�p����y�tC���$B���"���Y%��:�;s_Qڌln�鋂l�VJE�j:(M�a����qZ[�Z��\e=Ĉk����0-RΞ���Mm]�}�p�LIh���K�o�h{�E�����6�bѬ��lJs�v{��!�"���Ɋ�UM�+�+K��>�/'*=)m�]��1���8g�`�k�����U���&�)&:���#��uث�`��q�9֌2-�q]�� �p���*aEU�b	�&Jnd�t�W[�3Z�PU�]tj�$޻�X�jH����[y���� �)�IR��ud}�5e�cr� ��2[wu�M=nq��#BS�w��(i����=�]I�f9CNM���u�y2���͌ Yj��(�c��h�MKcn�y9��V�R�.`��Pӫd߻@�������8Jre�u�r�f�_�`��r�D���l��q���V;���;0�vvا�8%��,,6�6�8�f��ث��k+J�
;�^�P��{#]��I��pO��������4��z.�閥��f��ak�7ar|kk��Ne\|�I�}��@ڵ;��m�˵#��v�|��g�=:���QW���/�H5�ivi�ݷxˣ�3���\�t���z~ͳ��k�
a�쵟;�3471R�Xeª�YNr�2���}�P��3�^#"�D$�O�,�;�����\��=Ф����d��M�g���m�̭.kj���ՇO��	qR��aNp�"D>ь\v�ٍ9m�b�V����7 $H����\x��Y��P tÄ�� ���>,��4a|�ܹ�ܦ��km�ἸFD�5}J���wj�-�6���S*���Dg��we���X�s��*���8� 㔲�����8fa_��xt�˙�E��Wlt�����ˮ�D{�T/Z̎���Q��Z�<��qV�N��ۤ�5��iY(�GF�H/2༲'rbm&�HEr�V;X!���}�����A�*9e�]�X%���U}�4����Q�mj������բ��΢]o��m��w�+k3����0�h&ap�"�b�ܶ�Vs#C�/�z_P6`������qʲwh����R*v�g�u��x��t����u�U��m��{�F�u�k]��u4Ln��*�	�Rj��Z�:��Dw��wR7z��p82�&S剂0�k�vM��[痹k���M��L�0E��
��6�P쩎�����U5�=������5v �W!��ÉVu�e&6tZݫ��7	�p
�\��]r��d��\����)�+9W-�n���2�3�N�XN�7���Æ�5ڌ���v�C9C��.���U��H\+o%�>�[�Y�2VQ�uj(�I���3�{�0hsJ�E�wyj����Ƿ�v`�[ET����UwF*'�D�`��U�& �[�^�j�S��<g�,ӬIB^�h�X��aY�L)�(�/���S뺇�#7�'�Hv�N;�K�4CΫ� �=��K�Le��������Ք+,%�k��]u��9(j�b�u�5�.���*�j�χ
�3�Y�A��-��r����¶^
� ��CK��r�p���׮����D���f��f�u3w\i���ъ��	N��`=FN�Bv*�]��s�sc�� 
d�a9)�/4mp�����Uө_s��&�Y�' �j��KN�"�#��Ƴ��9�W�e��n��@]%�-F���]�Y�mp79]�)X���^�U��{��w$Z�U�cH�%r���d+H�ǅlK\R���V���#����eլ�48`\]d��g��.�u�U)���l:�i�pFi���b���@]L�����ݸ䮖o)��(Fmb}}���V�a�F�1԰�y����P�l�z�o�)d���\���p���T$/i�t+1�Rﺻ���oq�ȉ�}L��#nW�P>������V���~Uۣ�[� ��Lw�����v�qB��-.��[Y���,Q��0��N�YË�i��t38���:�,v
2����r�+�`�����X�vL&�
�M
��N�`�v�"E�O/���$ɽ��v���eq6��X��;uA��l�<��bm���ժ�4�Ӿ��m�C�{�4��c��\{Q���u������u���&K!w8�|n�%�v����ږ��#�[@h(��S�0'^U핵!�+8G�r�c�z���;J��#Z9(�..�Bj�i�;��Vj=�+��WG�2�{�<�a'^	cy��q ��0�}Z�]A���[.�cUp�,���u����LUҩ�k��|Ҏm<C(FY���n�
�_]�*�po���:x%G(�z�Sx4۾F̎�,�{x�'�t�'�j���0�BkV/i�sg*4.�>yrh��^<�\�$�S=��X\���e_ןkS3!�Q��L� � �}WZD�zJ�����֥*v!u��]bX�95}ujr-�,R�Σ1�ߓ|��c���vF�ή[��<۲۠�gVռH
���:��e�����*���;���5�Pi�����E�r����.K�.�A��4�Z�u�{tm���Ρ���G�VK�'8�l<�r�e��ݦ,EӉkr���уv���lLl.��]�MF+hTvZW�Vi��;^V���ϱ�����a�x��	\�me��RX��b�U��5��f�ó�lR�i����8��wl��uL7�r��rAF�1R�j1]�CZ�g2V<*�r��춏�N��͂*X�㖸�Z��l0�u���<J� &}E˅�z���Ԛ�E���Z�@M��f78R�x��yѮ���:���H�W|jp�3��Z],ljr���K
+�cѮe�E��ӏ:�8�n��P��NgG.�oZz[�à���c�4>�J��Iq�m]�EV]���2�5d]����8�%UΘ����&��6��\�=\�z1�u	L�Xj�T{l[�޸w�[Fo������PL�%M7n,ڻ��&��p�<E�߭�t�]gS�I\]K+�����É�zv��Cߘс[��R}J����&)�VR�	��/�؋\^0�׆֙yyj��JQ��h	PC+1�e
;�z����u"L�1ڜ+e������5*�v7NH!ߘ��o�L3�&��SF]�`��yr���x�aT��ݬ�G�p\"ͺָ�b�wi豈���_|���ƶ;&���+�@���Ed����w�J�aN�g8�2��zȴ)C�]m26�`�-��L�����Uh6��t�;0���	ɒ>ش.�oA�Yu���הq$1�A�:̬4�<�Y��$߲�Q���c+r��,*k	4,�إ�}vUlU��Qd�B9�W�5����r����u�|�_!.�@y�wu�Powe��k���+/�~kz�����M��?���\����ԫ�],��b:_u(2��'�>����N�2�=�yDLgN0J1bt��A�죡�΀��$n��__� �jCe�j�y1Ky�ia*�>��FV*A��!n�լP��f����1��-cv��K�����K4]���:&�4F�h�o4ѣAV�j���6�vnI�,j�6�,n�@XZż]Gj� �6�J��B^�"��b���f$/��Uj�z��9��M��[�:�o.����ü�t��z��H<����cJ��Q=
,}�V��թ=��̦�:h��,�R;Ż�m�v'f�ޖ�X��CF�]a�9Hs�N!6�`<#�{
C�vsSobͮ�\�����uhY�_�73um2������ �OC��]�.P���^m�����X�
̡,���q����v�n���J�/w�H"b�u��v��Gz����+呍GO����ס��;�m�Z>�Y@V7c@�S0���)�6���7�|D����%*:�4�25��w�EPJ�gx�E=;{@꧴v2iex�a	[�!i�Cb�֫wV=?�꯾�z#���Vl��麢36��;Շ�����jH -
�Xw(n+�窊4��֚�Ғ�F��o�q[ Xߚ�����#K5��L���)�ig��������h��xWigO�ޤA��ش�9O�t3�\��T#����f9�w��9��|D.���Z�=;W%b� �p�*�3]�b��Q��mi}��ʃ�l��ͬe>5�[�ow���cq.q�����i�:ˢ���j�`Z�Z���.;������m��Κ�b��!�<��[�u��o��;�r o\/@1�򎕁l,4�XVQ��΄����{g$I���N��:ut�\`���k8?��7K�uD�pَ��V�a��:�t��V,�wOf�܈)���$��r�b�3�m=��$�܆8kh�P寑��K�����V(�{�C#N���������k0�՜8GRU���.���q�˺�l
�:�V��'�(�I�1C9���Z"��B��:���W���t)�#&n��ĉ� �,��m�������Ñ�z�ՂR���Ư�+�J5�j��w;�3xކ���ʷ�Z�;�[���er�2�ͳV�_Jәw&fCr��_>y����,�S�l�&��Kz�]�6�j�\C��pWr�b���<��+��	ԙ�F��k�����.{B��Ѿ8�n�ɣ�A�s�x�v4����4���j��ZH��ih
!�����J
�(Z���&�R�"�iH��B�i
��rȤ"
��B����JJJT�����JJ��(hi(h!J���
Z�B�$�h�R���h�JR��h� ��)�����,��(
Zh
 �b@�hhh
�h���������h� �����\��(h

i
Z(i�(r!��%*��Z@��i�3(JC#%JR��R���Ɛ���%J�R �$�bZ���|����~+�}�s(gW`�ܓ��Ί��3n��{,P}L]�Þ�f���s�ak�O�S�	t��״���h��:�y���rQ6��Zx�9��٧�ݮ5�Ȋ��Q3�
�"~#ƦV^��fy?r���.�(g9��<�j_�G|<�2��d�:s�7s�E��\�}#�<�e:t�A���C3\�V���I�lZomѶ���d��nw�)ӌ�Rz�3q+z��A�G�8�o7Zݨ��lq�]��S�|^�_��Oja�~� �T�C����xQ̧~�r*3�
��&����8{&C��������<��N6���瓌�J/*�s�{:�e"�϶E鯶G�n;6x����Z9����q�r�:Bב��x��2V����]���q��;�Mv�vmB�۬�W=qY&�VC5���"��R�8�\e���q�G;*{3^d[U��F	Tu���1��L*��di�]��
��{�7�0�=��&�����������A�t���V6D�F3�V)�z_n�� 	�/A�Ja1��QZv�쉗u����6��ru0@R3:T��1CW��bWW-G6��7�@�9(����1ʮ.x�]�B뭳��9A�ʺ�Jf�@��hF�I��,���ms�����K���p�UbK�ƪ;@~ڪQ5��<���|�GH�����;��"���{�g6��:���F��]+���qN��W
<�6yĨ;���ڔr7��e���'Î�잴�]�:+õ��;��Ô��S�۔sv_e@^o����z�;���q����6Я�3Z͵h�/3s:rw�P���޾�s�߇5��+��UqM�E��F�ܘ4����{��7)��=��׊'�������253�
��!K�<��]��e��j�S5{=�r�sY|6fb4$<i=꿩�Y�3V��Z0�QκFxD�G�\�r��C�{r�4*A�4����W��Acn��iL(��2K�hV,�hۈ٥�vŶ2�6�)2�:8���zn��=�7���==�5j[�-�ϩt�Ã���(I�1d��'���r�s� �q���w�eҲr�Op�����w�w�B�h��gv�q��M�lA���
� ��(Z�jd�+5��ԅC�v��vn�w�;�9u��|�$�77hbY
���W��s�e���L��1�8��6��y�Ipk7Bj��iqǰ�->/ ��t���y�E�8>	���8�zv�9d�r�f.�#I
�Tr�'�ٺj��VZ��yMfҌ�x���&��V��b�A8-M�{�'Ջ�z�O3}.�ҰU�^��q���C��M�/rgY�^o����㈥��6�:�����}Eg��K��[ޓS��T;51]�Z+zo�XSMnz-�ү2�!Yri�K�jjcX�7eD�IN:δl8:�7Ϡ&���Y�!7�}K%X��k��[*��鹗f��1�gA��n"�I��	��p�<��'��ܻ�â���o)���m��'�1O��m+����(\��*{ܘ]oL��L��]�&(�zoSpW��V\shT�lθ���9.̅��r��͚�{9��q�|�n�������EeO\��s�S��T^���gb��"&m3p�6�<�ӆP�$ͼĐ����L�9ЎR��7�e{P�Y���!^����vDopּ�����8y'�����Ⱥ[u|�����is�ׯ�1�Ybj#c�Qwd�u�H���E����n�ޔl-�yz��-n�u��jW.vbPt��r�v�n�eQ���}G̻sp������X����t��'����R�z��׼�Z��t�\����0��d�Β�VS�u�*O]��y4���v�6�)w�E�SJ-8�M�wM��#���ʱO-z��c�Q̪�L�u��⑾�n��	����)�oe�h�4��3��[��|��>��7R�ʖ3f����p�<��X��\k�_3E�����id�0��@|s­�ו�e1y�/��4D��%��g?(Vt��~�/A�y����mU�t���r�Vui^c6bqw?p�Si�'�����ky?x�ߔ���ߢVn��gf6w$���e��k:f�qo��q<�
��4���U�*�^ϖTa�p������}F�ASX�=ћ���@�����r
x��9�^�t�%f���q��vJ�#:1[�l�YC�hl{)�u�Y� j�Ӽ'?b�ѻ���mj�8�Ҭ[�ݣ�<r���8
�n�:��{�%}/����xN>*��*��Oac��0�����꼡u"�*��)	���r3
O����?�w�Vz�V��><���$��{���F��ӷ\S�wۜ���[��YӢ�3e����+�ㇽ��.��u����u�z=�˴��aݓ|��;=`��v�C�_WZ�����a;�*i�s���8�>���w��&�w��Hp�xP/x���۾Ӹ���e՝y6Rx���Tïʱߛ坐˾����*���Y������N#Kl���*����NE�z:��e{7��G��<�h�s-O9�ZaZ�NS�R�=�{��D�yɭ�U,j��j�����8��ެu���.��(��O����.�u�'$T68ܭu+��+��ݜR+y��7j2a�2�n�)CT���W̂���ez6�)2Y��5����
1�N�\�Sq����V���^�ځ��ɕ��8׷T}�'�;�2�c�"�Ut0;�ٷ�J�]1��$��ym�S�ƅb�c0T��Q!�Z�"�rT�_\s^��[���:����]5u��|9��}�U����듺�pT�E�g�c��dV*�⺅������mt�8:L�{q*Q�.�t�%k�����uA����Znu[�ޗ�w�;5<����r6�QYW�ٹ���������Ū�9��e[����hYe��[��v�םT�8n��Fe�<�3M�b�\D�*������7���y^��{�\�޻K�K�lJ�{�l	��1X���.r��[�֣�y1~ĝħl���Z����;��ӝ����,6{_��l�s˅�I�q:�)D��0y!�C�Ź�J�ei�`�q}[T�+�R~����zI"����N��T���V����ő�sq[��������i�/�gxN���!���y�R�Z��s���v��2�������vw�k�EeN�M'c;��s�r;������"x!���u���7���K��)%Լ��J���M�Doow�s���B��>Sz�0��Y{�~���g_����j��'��`��>u��ϭ�u������h�X��d"7����)���4�y�;��Le�(�`��V�}Y�u;�fq��T]!��E;�%&&gư�[�&���ES�Z���ֱw�'��ٶ�]�=B���z�5rᆯ��!�DF��_u!:�ɽ�O$��O���+o$r2%oU���aT_�պ���0��^7��&��٪{��n��H��Y�~Sr+P�~�Z��K��+,m�f�p�v�.�/$̛o�Ѭ�6W�p��l�0��}ae��6��1�L�N���ZJ����'.�9���I�N�^l�\s��}Ѧ��t�U�J�COL����Jb�m��w�E�8S�p�Z9�kӵa����)���Y�B�d��.�2zi�^SF3iE�p���&��V�'O�7?8K&�S�{R��\�gV#�[.�^
��%FAƢ��;hOj���`ͺAw�SR���Sӛ~��F�ɳ�7���m�G+�ެ~�UG
�p�[�9��t�����rv���&�ܶ�O��_�!Y~�N��P�
=Bθ��3�hN�/3C���O�&�y�Y�ɽ��Y*�p�OR�� bd0[���t�u�u����N�t����Pײ���p�c7�3!�-�V�٢��^��]]nL��v�"�Ɣչ�.ǋ�����ٷ�r�)ɞ��R�ա��؍�X�F����_36��e1��A�8�)˙�[�c
̣���L1=Y����gog��떌�#T�7�9�&��;˹�QV�U��M	y�;�*���֗u�R��9��1���긅ox�auT��[Q���h�W�t���ja�����c�E�+��9.+q���g��Z��a�Z'm��'�Xm
�x�	�Z/��{2�G��.�#S܆z({Nɾ�ܦ{��W���x;����'�WOk�B�#�6ﴱv�>sVN�w�w��(�b��۾��sl)�,d�:p'����#\�:�I�M�[z���g�(�_!*��汅=s�yj����1�����Ǩ'z�>�7��vqH�n���Q��� ,��IMi�����㾤0ת��p�R5�Q̧��lo(>���ڋ� !��g,�B�e.�}�t�qcg��T���UyMa��gc�62帽�C�ivt��\�� �L��k R�#/�P�}]��xa�C�.�BL.JV<����<k��̨�_
`a��lu�M��kRb�l���&���ba���f�,
*�V���&�Q��K25ȋ�1R<�*��ɻ�`��ۦ�Np�ؓyq�
^�u��ǝ����z)�K��ߥ�_/k��:���V�̑�ڹ���Y�pl��;Ӊ�q�ۖ�o��i�y�Gz�%` Mf6g����t�ޭw��s�茾W<�.kN4��ڨ��{7�9����Һ�[Yn{=�b���@V�/�ټnXNt�q��Y���]9��kvn�Ffƫ�vK<fXY[�X�:�7͗��O;��ѩz��[��-)���O��ը��ǝ���՞��~�]r�QMa�P��<��P�s�œ����ԩ�.e�\���;=`�l��:����2[iI��*�/m%��;���U��*�C���g�;�;���g� ^��:E0��j}я9�s�'o2�7�r���Y��]��g���C�=Ɋ�c�"bl�*������1���*��Ә3d���u���j�9[���A����FY���{�{:v�@w 7"OT�UTB�<g%sw��.��n�Vκ�DC����b%��9�*��u�Џ���{kw�\�\yZo7�/��9�_j�nsn�"��7Dޥ)cГ�]�1�L���oDPU�c/�{7GE�V��wD;���cu��h�b��b����������>��r?w�JY�'���ι|6�Q�|�$V��r����X� �vqH����`̘��]��x�nQ�bf��%�Ϛ���;��g���4�xпz�-V����k�cZ/է Tsj.+A�QM�3%��\pҺ
��#�b��޷�K̮��x�g��z_{y[��O}�\�ͩEt �;y���.�?Ks��+;�V�9��V�;�MY{�o_����	��}����u*��O �����Qpq���9QI5�kc�(�|�-�2f��w�����ޫÉ�k�a}[\L\F$�t�F������gy�t���q��Ֆ�l�W	��J�g]҉����$�=�Gu�J�����	�>zq�m�4��ș�t럼!C�S�l7��QӞ��$��:#*�	ϲ�T�;���X+��3ST��#t����#L�S��w�L��k8ASt���\���gl��F��a�:Na�}�A9��13J�F�Bc�o3��6	o%A�N@�G�R������Aun��!�B����|����wZ�H��mі�-JD3h����{�#�e-������1�2��*�AƭH�k�"����}K3i��[{&,�����ڀ8�=+L��?ej_Ҡ�.Dev�M��@d��[*ƄJ����h�z�����:��8�fp���G����im����V�VS���<L�v<}���J�<���P�ל��/�f�ͥ9��ܩz�K5�{ǲb�bsk�үhm�r��6�8�8�J�	EG6Ie�ʥk��1���Leq�"VtV�uu�n�$43ԦÛynf�ފ����A�(t�<r��x���.�&�a*}mw�\���I�{�R��.��ӫ&���U�ڙ�n���X�J�:Q��C�9#ukB��7\qRy�.�e\����_b���R��+�Un�C�{Bu��9܆�q�-��L>U�p]�g}�q\&��~Ⱥj�=�VL΁�M�� �����k��Di�+p��Y�`X��qcj+Ȫ	�]kC<�!x��$_eN�zk���)刕֦��q�;#+j�S��a�wt-}E���eB��rB���ͫ�����Ӫ�x��|&��XE��:�uն �phK������]�3)J�D������J6���Z�c��_f0.���/��V�N�N:�nvp[�v��
e�N���	JE��Nv)�m鳫:`|Wm�x���u�R9�N4jp�25Ƹ+CY�5Nq��"�+P[����Ꜯ�"]�tgw�{}�k��#�WS^w;y�F��*�V��42������n�&��g���������z�=��;�D,��� �IM�l������;Ye�:�Gw7�-��;��,�l��MC9�e9�DZw�hX}��ږ
��}>�M�����u��7q�����Sy()V�ZZK�۽&�C�q�q��o��o�`�] ���Hٚ(m�ĸ�
Q�*Ǘ��e�S�V5[ �#�$���\}�_g5�nhmج�C�)�˒�NhO�q��2��ufN���4!��o�$�8�����S���*����%z�;rT�F4ӿ�6���$1�y�w�����M����s���c�b��;5k��i��>�3G.��Z��*0��-M�����@�'t�2�9�顜O',0������G7�-����e�\�Z&쪈C�X�M� �)|B#r��k;�f�[|�rV��^�v�� 5ʋ5�sٟIz�̴��5��w0
\טa�y�$
����fY�c] ��9Z�7�=sz�����={�▚ZZ�
�JJ���!�h)Z����{�
b�Ī�J��j�����"��((���bZU����(

��2B���������2�("h��20"Z(
bP�hZ���ZR��C)�JH�����i��)����JR�$�*
H���i*�rL*j�!��bZ��(�H��P�(+$�J
*�*�����ihJ
��+$Ȣi*��"���*B��Ț��a�")"���12�&�h����*J	���"����h�l���
b���((��))2L"&�����0�0rL�?G��	���������lW���xP�չ�D���髡���U�'o#`�WR��|����,�I	��\��t���������q�;�~֚4�:E�_�|�C��ό�'rᎌ���W(��	;�Л�V:U�;��>d�*�w�ս�)�O�y�Lw��˄���9�.�.�W��!�_�e�<�v:�p�*�m�,��뚍���Y}V�/Q=83)��+=�/9���[/����yEUا_����ek��,��bN�3����K��F�y"���[�t����/�b|ߏ^F�)h�Os�o������pV�rm�<%�h�;x�WO�z���,��'C���B���g6F�k��bÃ�X�'�x5�e��PO}�+�\sBV��l㋾w��R+����龃+�=u}1d�nץ��b1��:�n��|Y�s���e;�z/y�)��L��h���w����z�V��fNU�9^�j�E�4c6�^Yw��6�Cb \�'���fg�ۑԼ���Ϭn��5e^���1k�F6��X��棽�٢���IBӽoZ�X��\��ڻ+�|�nR��
_�abyScC�W�r6���K�B�}O�f�s�i����8�1�mJk����.��8���Y�&�I^Q�z�_w x���w@�\�#�IgV3�[,,�E�(�8�\e��{���׊ɱꎰM�����I[Ӓ{|J����J�^l�}�s�]�3
���x޽�Fs����JV��>��kr-�ү2���^D� �F�q:�n�oƣ�í�Rb�Rw�O��Ma�=97�ԲTp��X&��s�nΩ�1:��|0�XqB�^�O�zq��=ˢ�zZ�7�]M�gA��n��邁��s�S���½s��#�J�l�u�'V�[A���G�ٶ�M���ʜxP=��C��fu�Ǜ���6��w��T�ŕݵT��Fϙ�H��nb���I���u{2;�_�af^�W7�-{׷鵙c�L꒶�z\VI�P��=#��{I�$ۼ�.�����D��sK6���ۉf�`Tj-O-��/.�ޓ~��WI�7Xa��*�M�ج-V���4YOh�ᓃ�N�Dca��<�9r:����󽜾�Θ�㼜�k���z����bw`�D����f+�X��� �t&$����k)��م�ܜrk۷j*t;�����M�"�O����gx�v6�9z��)�	�l_�{q,�<MIWd�ً������5H�a��*[�7��+=�풮Kb�MNjVtB��<���!Υ���j;x|eC��G8�{yRY���Ϋ��ܧg��G�P����/A�q����<�j/v��j�V{�]���+3ϝ�1�B�Ti�9���~,�	����x�j�/2<;��s7&{R]D�7\��C�2�a��/,�γq4/ŧۖ�[=��:���^	������އ#�z�j�88�5�oQ�}�kr��*���롱������
��Xqt��d�l���s�@Ma{�V�6�;��{wGR�Ɨ{��پ�o_����%}���X�����M�����˸����J]���G�{�F��~�~�����ë����]������>�Y�|���ϴ����οt�'!;�Oc%�
N��ù�%}�q�X���~�u��~�����=Ə)���q���9�o-r!��9�Xv���ac�m�|��ٌ`V-~{͙�r��*�5�	�0�QL�"�kE��}z�p]�&f��d��r������飻�b��6�|�t�]�6�U��OJA�Ζ��Z���	s�8�����)�y:�Ws���W�O+O���{�~����P�����/dz������nG�ϵ�;�����u�����'Ҟ�a�2_���0O��^Gn�_!�c�b����{��7�B=���w��|���7/��y����r�y��r=K���{���'��|�;���y��Gpvs��]A@���%�
N� �>��y�����gƬ���s�w�:6���y��J�:�=�~b���p����}i$9o9��p��?iy�����~�?Op�o�t� ����
��=�yε������{��;��C��r�~�q����=x�W��x�×��{��9��|�zC��7�y/r~���sK�#�B d3Q�Dh�TH��>_t��Ֆ�\j�)��D�{�Fa�z�H�y�#���xk��/�W}b;��:�Y#��=�r����t�GQ�;}ޏ�=��yuQc�cѢ"%?��6+�s',������޿wĠ�.য়��;��{7�}��O�ם.�!z=�Ò���w/�����rG�:��ܝ���{�";6���B$z>��q^/U�|u��^����7��?p��=G���_��9�i(7/�S�0J���~��W�~w��.�Ҽ�}����!��_���<:�wz#��1h�`�1�����d��⵶��θ��������WS�u��9+��oz9.�;w��w��~>愡�^{ގ�z������?ih���L���#�4{��I�8�8o>ϻ���ߺ��Ǟ�MJp��r�'��q#�yy��A�h��G���~���|��������<���>�m����:���4z=bd\�M����Ϸ�k��š�ԅ'R>���;������^I����Ի��;п�������W���oG%�dg�i�%��o�_eθu��w��9,�P]~T=����#VR�{u����ol�F���"���p� 
�K�QG���fׯ��Hˆ�qx `��W!�\��뵥1O��]Ъǡl��,��WK�e�I��x٤_���������ح��؋x[׭L�)~G���:�<�A.+�G��G��t?]H���h_K�d�W���C��Ի����/�r^A]�ށ��ٯ��;��ގK��=k������$@��f���D�#���<��ߺC�}����=�_d;=�C�{����|���d�W����J�{�仂���?C�y9�o@�=��\��t�S'��v��Ws�G��=�K��G���r�m��1y�>_o΅�Cp}9.��5�~���vkJ�#���J�����d���i�D�狶�f�b=�<G�G��Ҕ������м����wy#�綐�>_K����G�޹�K�y	ۘ�K�AޱAԻ��a�_`�jN���g�VL�r*�Q�(��ЄP��Gΰ<�����;�r��7�R�O��G/dz�����~�#��֐�/��ϼ�5+�o�iu!=sA��=��Y�7>5���t���3�D1C�B8��R?C��Oc�]ݦ�9/��N��ܿK���ޔ�ܛ���B�.�Ð�{�[w���^���&�~�6���?��"�W�F��|����� D<�`�y'N`��~�!~����'�Ԏ�`{//җ��p������<���}n�~�O%�1cy���+ݛ}z^�nWѷ�{�#�����:
Wpvs�:A@�<�%�2\��>C��h�w/#��>�sܞ���S��F�9��oX'������eS���=�S7Ks��`�p����=����_��@����_�
Wpvo�t����9&K�d��7����X���:���$wA�'�����{�}s�O�S��;̵֛��X�F��=DW�?I�^~9�:�p����Pu/�S�b���s��)C�뾗Q��>���}�@w�]���ìGr�>y�%wջ��kϺ�3?;�6Z�H��OAw���I%�����2[��zm@/�hȉ&�ftᵽJ��\�|�֨�C�3S68�6��9��:-��8:��Q1�t�\\���쫗��h�:�2����r�(�n
}�kT��Y�f����c���ż�^���{ފ��O*��O�о�ܟC���'���%u'G�h䜕�,u�=w�%��=�9�2!��?t��o_�]FI�S�CD{�:������3k� ����>[�@���x�y�?Hw<��<?y�J�2N�>Ѹ)\�7�<�pP��撃r�'sBP���e��G�{�qV ��g�eMq�q������y��.�п�������������`;���G%�����z��v}�H�I���9+���z9/ђ��rn_#$��~��7������UU�8�f��z �p������zǼ[���Q�ش?�$:sr��r5'RnG���:�����/�u.���$�h���k�3g�uuk�y�����w2�P����}������{�sH{/�����j�/�����������=�f�ܯ����'$܏Gxy=C�(��%���>�����4fV=߾��Y��z=�<DGՕ<D{�"1}���2S��4n^K��>w�!����y�|������y�<�e�=�;��2:;��/��;ٜכ�����ߞ����k������ػ��~��:�~��z��F���>��~����kp�w��w�/$>�����_$;�n2^��{�)�z���G:5�=��Zs���А
��p�z�D�}b
��{.�$<?`�'%�d�~ށ�<�7�>�y'ٽ�w�?��7���w�/$=���[�ԛ���Y�_
�۪o>]ݛ����!��P�!=R�22p}>`r
G��7/ђ�~�����oJR��Ǟ⼓�ގC��^{b���>��}�<�d�7\v���(��;}��y�4߽A9)٘NC���}��22G�wu����bn_�$:���~���~<ޔ�ܝ��o�z��G�B�-����Q��ꪡX��F��5B��Zc�]٨�{6�C�䙵�cA�
o8��3^��ez�+����M��֦�s�;������K�)��x��<�nU�\�\�f	(�h�4c{y�]A���g1�Rr�.++*�kH�Q2���:j�J�+��/�{��z=�>���_w��:���_<�g�w�zMJ�ѿ{�u�����(z�C�=��ۣ��p}:������~���QDC�4DJ�|H'���i�{o;����:�h}!���r��y�/#��w�?ig�w��L������PP=�����zu�nOe�0���>�3�y�_ݪ���돷n��8WN���w��|���c�!�{7֐�C�;����|������_a�����;���~�(]���y��_g!��B${�ꘈc���B�O��]��O��޻�^{�?Y����qüOs�z;�����<�O����<��~������Ի���懓�?AO�w�y��k��
G���C��;׾�}]�l᾿s����{�ζw�j�Q��?��_��R>��p����/�w����G�4nGS�;=ޟ�rW��j]�B{�i(�p���Q�Dp���BX��>��~������k��~���އS�>�斗��Z����u�b�Hr:?`wy�?Hw��<����:������z�}�ŏy��#���}֫3#4�����9�y��%�w=�JRy.�ގ�y������W�����_�:5����y��M�~����K�M��<�<�����#�^oό���u�w�Y��ל���q�.G=���w	۾i���2O�sBR{/^s�^��^��y���W��x4?�d:3�C��?u��;���#�y&��~Qy�w�������{�y�!��pW?{�|��;�����|�<�s���i���2O��h%�^}�_J�/�o·ۨ^���ג��'���~�g�{�s͚_i��ޝ�Q���ǣ����"ǽ�
^���} ��;п�䝻�G#�_g����w9)���7/%����~��Nsξ��C�~��j��<��R͛�����P�D��*e�p*o�p�܆���^�	[�v3�P��L6� ����Y*�ݕ��BS�6��s�\�B(�����;+y��KEA�f٥��ⶣ�T�c��2��Σ�ǂ,>N�օ��{�u�c����\ �5�g��Q�{��M�|��L��?F��?�X���t���H��������<�r�2;<�H�&����7��?���K�qǜѹy.�D{O��|=�{���/�%�������|k��Gr=�C�{��2S�ԾϮ��G�2:��P�:�A�y�O�ܻ����~��p��r�W�dK��{�g�����1�V��:~����z������w/��{/󿴼��m?hu�)>���?A�S���z�J�#��7#���&����>�c�b$Gc�z ���lQ�eqK�>5�[ϻ��xjܮ��y���rG��u����<�K��iοt�'!;�Oc%�
N��9��{u����gX��ǽ�O�����ȧ����;F�VwgZ���8{�=��ګހ"!�7�Gײ=Kٽ��?[��ϵ�;����u���Z\��O�Ðd�AI��	����ъ�&��~?���f�ֹ���{������{��sX���اn{��]���<=��C�v��[��^�ޏa��_$�o�Gqܼ���R;��u����2_`���=����y��9Y�Q3��s�]�`��D`�P�����{G��Pyd�����y�)ٟh7.���M��!�>9�[��~��x����N��~�?Op��t� �뿯����J�ʾ��77���D���H�}9@ne�0�ܾO��r�]�]�{^Ju�w�}���}i$~�y���'�����w/�Sז������P������������G�D!�5%~�{�K��^}��!�r^�`�_e���Gp��<�G�<;��9y)��w#�����/�;�,��^f�λ���k_y��Kܞ�q��%R�=�9�y��λ��W�~޼�u��n��؇z�ܾ�˫���}�;��ܝ����/p_{�nߝk�������O�S߬�nRŻYďή�4��I�d���� S�������^�x��*�ݬXƃ/�"�O���XKeYf����]`<�e�]]J��� ��}AL_����U�\�{T��;آ�u$"u"p�������]U5˻��G�#���Ǜ�zWg�{�"G��cyC�F���w!�o�J���}�	C�s��;�䟍��K���?�Z_�b�ܿC��5�Gܵ���6����0�˛�G~���y��ѳ荎���{�J�r��G �r7�9.�=�4��>�A�0J%���G�~��t����ش=��s�}��׉�*�eTZW��ܛ/ЄDP�pc�Eϓr�z���^��?��#�yw���9i��9+�����F@��C�}�����K콼�ξ�����������]}B�~�P�����6V���
NH�O�u ~�'�y'!�y��K�+���/�7f����W��oG%�d�c�<��0rܑܻ<'-uY��{jRo�{�{�f���>�~�~t?]H��š�}/q٬y+�d��!�w�j]�K��_ 伂���;�>�qԯ��ߞw�Ȏ?|�7�Q���E�x��}�P��Ǽ�þi%�o����}����>ڇ�|���|���v���9��)_�^�9.�����NG���yΎ�hD�[�<��Z��q�#��VTp�=A?�������|��a�4���o�[�|��xNKԟ��OѩwkJ�#Pn
W�{�6���D}�H�\�g��#�DdǸG�C��v~ޔ������f���H�N{i�����sK�Gf��K�y	�f���'�d� Ի�ѯs�-�������y�}p�^��5'ѩ_.��_�$:���<�~`~<ޔ�ܝo��^��|ޞC���ϭ!�>_K���t���;7��]C�M���}��3��~��M��}߾�}�5�?A��
Nf!��q٬5#�?GgX�GR�]���~��ܿK��=<ޔ�ܛ���B�.�Ð�{�_s�:����?yg���\��':�p/����2���*��KO��:`���0ص+?~l#e"�:ۍz�&B�G��z2V^ŵ�[�g4_f�}+��Y+r<�KὊ�M��P�g	g��S��|��5*�r@q���{��-��g�u���<���jW��y�}��z�;�%�
N��7��{т�����Gs٬e��R�r���|o�	�$��5��^��:�>Ն}پ��n�s�u�~pu?��N�>�пGr��t� ����
���/ђ��7��8H�^GR}d.�<�����D�C��G�!�药�ݹ��e,��u��}{�>���e��9�'�~�����w/aοt���?iu#�rL���~��}���Gw��0z>=b"�T]͌}�w;�%�<�/%8��H{��f��NJ�|�K�|���i(:��)�1NA侚��=�]�����=�ɒ�~�T��{�=�`�̎�VL��w��5��_g���pp���9{rv��[��d�>��rrW�f���'n����_`���Й��s��{���c��z�H�{��uLƟ1�U[ϩe��pir�%�/��}�������pv��?O%���k�����ϴn
W-�C�(M���|��q�@��Q��~�*�w���@���H�/<���/��b��~���'$>���~z�w)���9/p�O�؇�Լ��>�$}�$�������>�&pc?,��U]�V��q�9�nF8�Gf��'*��x"Y�Z�^SF!<�է�s�{C<Dn��yq�
^�)׾,�܄��ΫǛU}.�V
��"�S�gz����j��f��1ǧ�ᄚ���ȵ�����zsn�V�bsHa�L>����Yf7`��X���W�["C���UǴ
D-#�޽�;39(��P�:캙gR�t+]na��CH)[pM�q�3]��>#q�[��@�N�=���{u�r����̆��$���}��G(��J�IWC�����RAR��'���km�w.S��m����k���K�4�eWu����1$U.DϲY�qD�Jl�*�v6w\�%�`�X�2n�(!��.�+:vͲ�ŝOD1G�b7W8����oGQU�0����j��^1MM�_jL���T�'9Q�L:k+�6�,M��f�p���+lnT#�v���jn��\��&�xm_]f�|u`��M�Њ�.�|��f��1�^֫��ך���SE[��!yw7��_q��;���u�+5g`;��R�.��#ܞ�9��dp��[�z���)(��ya���U��v��i�)�,Y�	Ce�+wZ�u���g&��2�8y��,��co�]]�#��1>ܷ�6�~�=i��/9�j	9�Zb�0C���
���%f��c2�$�J�Õz����I=�]�*ە;�a��2���o�&�R
j>)���g8�q�R��t��Y;3�W��e&p�[�h�.7���r��Tʹ��6���u�ʾi�=���yιǗ�ni;k9�븭�Z�g��;|�X�w�P-t���Ԋ�`[�Tl�����]�'%cqr��d\ֲQ����@����|�tM�͵3&&�d�>��9'u��먣EV�x�ٕ�b��P�X|�M�6�Z�g}k%Y�>"u�s�� ��yZ���,�3��^���O�2]ry����������xn�ͽ�wۑ��]4*	)��;X(ꕭ쇩�Y�$�L�al���M�I��
5���V�c�F8���4NT�ɵ���.����RU���� n�8��7] 5��y��2�4'9$��� �It��]B�_f��G����3f��pWZN��,U�2KS0���2�������^T��|7:��E�c�N��f�泡P7�
��r񍮦����8S�@�wq^d�ZCO����U|0�UvUEu����)�l�5�%�����坦�|��i�n�GٔC\r&��b6Xz�rgPt�kk��`5�G�3BYE�\3�y�^�����:�ԥ�y�މK�\���tpŸn�����IB��^lZ�%���̽$af�-��k���2-�|hv[�0�L��5��0OM��(���@�s�=I��:(�-I�wƟ:t��k���N�=
��B\���.�農kc,m�������*9����u��u=h��x�.���N���CP.B	A�U����Ԯ/E�f�]���
�}���M� b�Y��5������U��f�66:���0i�[�Ң�$�OWy��;a��S���?yV���o+v�@�@$�P�HdD�Yd4�SIIK��%HPST�P� Q��KEAFaFUCT�2MSD�AIE!AME$KQQfDM@SHU-RD4%QJPUHD�QIC�STE�QMA4��%RL14�MPEAPIU0R�T3IJT�44�d4%CQU%%R�AT�D�R��L}���;����{�\�&m��7�8����ڹvV��;��0$�Yӊ���Dr�A���mvT�u��f5��UU������?!Y�/���le�����>]���W�p��O�[5]4�턳S6�9�:�𨽉������Iߥ>fk�w�{��ɲ��fX�W[�ת4��˞�\��\+ǚ��R/\'�+w�b�\�Ů��c�;��}��JSO{]��E��CϦcבͦP)���ǋ;�����0�]oL���C�ᇶ_�s�}LμA�f�ξ�[��qowۜ�r��m�,�CyS�K��h��)�����$������TН���vD*�K����}E�w�&Ȍ�1�^sV����Q�g�y3�U�ʌ���%��Xa�}��f��]Ҟ���X�yk.�� m:[F���ƥ��әLhТ��%I��U{�\�z!����T�r����'� �+�]��"�[�Z��NB�(ţՁ��U�ǛN�v��[�S+�.r�-��9�L܎�]�p�na�Q:�b�&Ft�}V}���|�-��)F�(<Zm�y{�s;96����E�-��R_�x�V.�]����lWc�lH�Q�m�mv���n��y�Ҋ����{ވ�N�xS&Vd�~Fd-�ey�l%��5+�J���ea�vg��j�ƪP)�nk�Z���Ϗ�*�2��X��3%�(;�3�i�w��N�2���ܥ��2�.#;�q���]�:ͱ;:�y�\/��ɕNc��We�J4��&oj"�/�����s�1��e�۞�Y��h��Y���Q˪�N5�tv�L�v�ɗ����p�sй�\֘ƚ�ih�WpՋ����4��Ud�~��r�Z�Z�\H^$�%>vᘺ��}b�i���;Gn�Ցrv�S��=�S��X�:��^��9�d�r�-�y&�/;A���|\��gxNn�x�N�5��kQt�,���z�z,�ЩW]�y��1�A���79�q}bo��;<!�%KN0�˛�pk�B�?Z���1�3�׭�*�w��rwbv'M�'��:˔(�U�)-�T�UD&������h�uzth;)4�2��_.U9�
)u���&m;���]:� z0�,f�C[�|�>�a�Y��qqN������i�vwU�Q���^�ԓ�=o*�'eΏ�&&�h�oc�BC����ޏG�=\K֝m;�&>���LwTE�w��䳱V;o�v2��R��u+�b`v#��U'Er���q��P�������]���3}�Vo^���a��������oC�c�w;G���ͬ�s6�*��>oꞛ�vsW�3}^���y�Z,I6*���GY�^�Y������o�$��ON�Ө��n��%h�ؿ����d�S^^���!u��44���Hm�uu(͜qw�p���#9@I�(L��k۪<�rn_Q�W.�l����W-�X�+-ʕ�O��:Z��E>�Zs͜�zqH�j�R��+)��NUÃ��m����m(��*�;��
sf:�R��ύ�C��E�v���Gj�w+zھ���_+�ـ���1�VR-��6c�{�=���7lm���*XOa
��S.yq���a�3�_�U&�'�YT�6��g���]puv����$�l���;�:�J�O��Ge�{��v�j�S�W�e>;;3A9��%-�ۓ��r$�t���啊 ���_.ﺟc�u5Th���ϕ�J0��s��}����Dtu�$��9֍�����ϰ�i��[}�Գ-p�q&��%n>�Į4��j;�?Wf)1pT:��8Mzq�m�R��������6w�32N��/-��dZ���ی:�j�ޜk���	���Û�_���f�s���޿��v)�������oݾq"���F�c�^�GZ��[�� �����+>�~���gm�S�΅X�����ff��]�UO�Z4�k}��&�9�4{�9�_{��j�*�FI��uͬ�]׶rJਿsW�QwJ�v�k��^�`����B�;��mF�{u��%���7�1?G
~�h��ۉf����K^���X�ec��S��9����v�{47�p����j�ޏ��J�ao`�;�uK�!�+r�����.����P)&�8XW�㺼����
���x�i���M�׼����i&�\�b�\n�f������R>���<w�qD���e�hZݠSWv��V/�"�@<zkr������$�:+Z�p�e�����]���l�X�.�#� ��ܹ�t�D�S9������#6���F{�m��Mյ���i�\p�)�c�{)�g=������rIg<L�q�^��N6����r�ʸ�9A�U���4}�J.�59q!qӯ#^Z��ͽ9�.+w�h�h3j�˰���T|o���Gw���s�ûދ��s��в��ȵ���n��9�L���jf⯟>�Ñ�|C���|��c��_����a�i�ȶ�UP�Ff�\�%a"�bW�N&�NϖS��@\����p�Ӿ.<�Q�/PS�];�O\u<i�̗c�e�R���.;=k�k(T�׭������ې�֟�ɾ�P������U���<xP=���T���}2:���+WU�t���tr�<bߴ��V��&=��)�xP=���@_S>;�Eu�ea�:�I��p5of.��w��l��|�^�y謝r�s�)[U�C�e�厎����.Y���9L��]���v�e�݅j���i�x�oJ̆��2��h�巳""���Wu�҃�����G;؀S�_v�ڜ��=�%J�Y]vdNݜ!Z.[{�2f��ĪtO�����b��R�`g��Z���Q�ִ���}���Z���䳱Ve��gd[w����ф�W�ټ�n�]v�{��ԉZuq]�Pu�ᕚ��V҇4���}�Z�u�ss�av���j�)��QtC �T�mο6�◪�!=�a�Q|���m��}�ќ0T?n-�F��[���to�.�)ِ��aT�����Ź�F�F�NpZ�\.m>�5�\rU��)rdԝ1=g5�8����M	���qwE�y���E�V��q��gf��'Pv�ザ�j��EB��e�հ[��ʂ�vKޑ��M,�Ϳ>ΫśU���b�_t��c��7�þ�yPX�����`>w�14.O�-f��\���]�)�%�ǽ7s��o]���L`�8o/���>\ַ��a������bAez�U�&���;�\-D�qǒę\�^>@h$��FL�|��������� ��gk�����D%3���r6�2;z�5�oK�wݖ`|f��!4�[zF����S��#Q9�v]�Z�8CѼ����f�t�qL�r��� �C��ZӠ
�£彋�[����7�����|>}��jܞ}����=��]I�'`�찲������T��_NÄP,X�R�Ql�7��պx�pv6�7����a�W�D;6*�~�հ3H%�]�VVО.�q��nwO(H���'��[�zgn1Y�0��b��W��^⏦�]�_^Ӹ���rO3���y�*�{��Wo�W`sL�����O��S��[/�y�*{6_^��9,�U��坞e�\H�nz(�޾���ڃo6��������.��k�8��S�^l���>�ԉO��֍�ܓ�l*D+�p��\�
�{�qKk�T[ɺӁ:
��\^Z�����@�$��U����GY�����΍V5���{��Ϥ������h㑼�l7j.���y�l%����jx�k��2��K∳3�u?z�¦��k9�M�,9��tBo������D!�۰�7P
K�׼p�:۳��?r�~ή��U�]�YķYwX1ڝ��䮞AW6���%��c�g�������	�E�7nLVf!ƻku#d1ˁ�V��ZͫױU��f����>���sEwkͮ2m]i��`����Dڞ�̺�&�Z��g���g����jeh�qwp)�����ky�r���g3��Y�r��qj��1�J/,�βK�3ǈ�N��@��Va{������z����5[*��d �6$�BJ<ۮ4�s2ܝ�<�Ӎ5��f�=ݭ� ��X-DދVn8v�l�B����ZN�8;�1'ҝ��a�&�����(��o�M*c�ͳY�[1���jл8޾0y�QΞ�����YŶ�]��}>�r)���f�qqU�q��'�*WXO��?h���ǥ�-{sb���j�a��S��z��v�v���q]]r��\��
���u:#%�r_��[K2�8��w�'��m
�
�#�r|�����`�C�+������tP>["�E���{q׋��<o��g�'�C�|[���׺��é�������A��eSw�HB�H�jeW^0���&�wf�&��6woi�YL�m�2��4�"�����p�ϭ���Ղ�yݽShI�Nse�ݶBC�f�4�ݺY�A�<����*X�΀Wb���\u�K��3�,�<�eq���z=-��>�5�_D{����tr9��(��F��9�+z�)�*ٗ�|n{��8y�^�W�+ٽ��%��X|�V�M�<%�h����.a)�r��{z��:�9U�.��e���R*7�E�!a��$>�Zx*��y
>�v�7!ͪ�l������W:��m�A�"���RA�[�P��m-�%g�4�\grf���_��ˬBpb����n]�/P���Z��tZUz�#6�#�p{�;�}��C�g# �fV��#}����JsP�N��w��LJ�}��� N�x��cf���~�q�'�@�~�N�ɿ[Ổ�0hW�hA���0􉉓���ȼ)��!�Raw�1U�u�Y��w�̘�T�ձ�;m���4F�S��ߨȊٙ��8|���ɡ}N#�L$�]qk�X|\�� �8�����\.�dC��J�g���c��a�ď�j��wި�q#�ԉd�G';�g��{B]T���Z�ї�� ��C��V���V"jX�ǫR�����5��XH��=�(b��/��G�����w��f�}�puƔ�-��&v�6xt�z�i�|W�3:Q�{�n�U�i$pG��EZw�����F�����Iw�ig)N���W�}U<ۏ��y�J�G���[f�|�p�!����N�P��w�cΚW�:�n�%�=�8uŗ{U�U.k;�A�q�c'��#ۢ���(�`.5��K�w�H�ᵾݨ; �M����Il����S�D-�#`�5�S�>�C���+&ܤѿ�g�����̭53¸�C�?�za�_^��Jَ��'����B=r�m����ӽt�I�*�z;o{Ӑ���c��<��H"�C���ϧ���Z��i�\�:s��33L�w���Ë+7N���O%��+�)=I�����HĔ\]�C�@������Z�ԟ�S9>P�\S]�o�Y�NS��0c�+�F�:���d�y�i.�-q�uV���ª_4=>���koFVG�����-'UK3��v)t��a��wb<'���u鴶�G���W1�K6*�q�Ei�`bd����.sg�Y`�ķ���%xم��	�﫾��f�i�B��)c#x㜯��5�b�j�B�͖5/}��c�`�e�],�,l���a�[`	�fW�R��a�6�\{]�
9t:,�A�*�ty[�0��U��c�޳�A�tV)�2��ЫY����;^�u�.,�����w��k,�jl]�CgU�
fvs֘�T�\6��'>�6�s������K��LG3��O,#®ً�Y+5,(���V��Zt��9��]�A�jL��s��z��y����u��z��lv42�[�k t*��|�s���)b�w���EڤҜ��K�;@a�-Vձg���A��2D�aMW�^cn���ԧ�ё��[h����÷:Z�9j� ��t�@Ah��Zkф��p�n� @3���\[S�4� Ilwfu�J�����r�X�H���2�F+.0��z����[�=gI�۱�^`
^jQ��˩v�nP���t<�v��s�j��&ح�	R�lB��Y�Sx�$�8��4��㤣�a[v4���D��K&�ѽ�U�s��Q�'�ծ��nỸ�=G��w
��!���3Ƣ�K�.r_��+6u4.pd����;h�o(�i�hN�HM]�1ҧur�٢�Y8������}(>5ҕ���4$֟:M讻���3%J����E��cͩ�sx�Мʓ\v�����^X�3��	'!KM[�F��_oL�>��ͦ]@J��G�P��<=(f�k���YF��n�I�9p[wZ^qo-�ۡ(&>���,����S��.W$؝x��=AE��2�y�"]�6SX��������oc��N��IT���ƻ�΋�W
��!���2/@uрm*u3�Ѧr���኶a��+3i��l3��.=wv���\���϶�p�Ȗ�˹c�8�P�!w��]��(yd�r�>N�X�t�Ѓ��
Z�j�N=�ޏ�y��su�1]:x)��EԄq�\�H�����={HU���GN��iP��w^�e�хE�!��r�lM����:s٬ui���j�b���cB�6e:�5wv��;p�h���gZ����P��1�h�5�tvޚ� Ì��������[̠����o%��X��"z��]RF�جѫ�����������)���ʵn�Y�U��JX�	Ytv��ջ�o�t_H�.��gq���oVt*��#|_�k�9���v0���ࠎ"V���<�%
�߷(֩]6�;��7��/�TS,��f���2�+wD���q��av�v�֚N�s���VC2��e;�2�Bn�o�A�.�'�/w���X��eյOj6�fn�ל�h�e�V*�R�)����<7�����O�6���P@)>K�..���8�vd�"X{�M��4�T�Q|��/��3&i��v��-A��E�F��i�v���r��X[�/]Z�$'�[x��$��G�e��m5��%�vvCj�V��J�]����qγ�S:����W=�cb%3aY8;�#t� ���I5���>�SIA%-5JP�QT�d�EDӑ�I@UUPPД�R�PL��QQP�CIKU-%LP�Y��QUPR4R��DICI35]FD՘�TSDP��QV�5���DDR4R��&kZMTY�T�T�DFYTT噘@L��fffa�fYIa�ICNFCI�1ՙ6F-Ra6XQEY.Y�Y�M�a��M���XkYL�N�o���E���5��U�JL'wO@��r�htt5I�б����v8�t�[��6�0qj)F�-���y�N��Q(������3�Bo��<+UU�÷h<�ۗ �q���9�E�(|p��޳/�����[k˥b�o.lDZ��6ŝ�RehnA��xUB3}��et��o�L��(<���L�h�=UiLw�֢���M�|*�o�.jc�J�]�fF�4�#B��R'TތZ4NKH�x����+���ϳ��x�N�x���o_!��B�\92���t��z����y�`�tovx��kell.��<!�dK�EV�k�V����凴2��;J�/�L�&r\g���0��k�_gzw�fW�C�.���*��
��m�f*�ض�<�|�4�wT#R�+q<X�k��޳�\\ׄ�A�~dm2���_�c8楗:ك��^�Ԗ�
����9��*�i���ŀæ\�x.]w:�B�N=V�C�\ǇOH��σ0]?SD�^ׇ*�uq~�P�e��iO.#��ok��"捻�&�Ϫ�̅:�=�gD�}�/�	bm����+���L���� aOg���襛(V��G
�^.]Q�ios&�vQ	7��>}�L�c�9s�K�%+��в���yW�O-z3�|7H�v�2�{�h��rZ���#�qn��wr+\����vn��t��i��򠗩Ճ3�嫦_�aY׭]�s��UU����}n��!B�Ftd��A�6��6=�|����q��.�.���Zǔc���Ոi�I+�7�r\�(\j���j��p*:0��xÎ�Z6#�7R���n�73kB��2���e��(2�u{5ؤ��B*Ğ��Z��Y:n 3t��Yu���p��s1��XWWc�X*g�Mxlx��}��扱�
Jr�֥��[�����~�yݬ����FǪ��6v}��g��s�HMe3(gmZ�v���d	�LcH.��=��a^�"�u�T���]����XX��o��Z�_�G�3���Tê�y�>yp����O.1�6����cˍ��5Z8�Z�8g=Tb�eTLS��꣮�z�P�軨;����M��J�&nz4�+Ftd�l�j؍��j�©��0i����������]����7�xO�h`>-���$���vJ�Ա�ݱ��Xp.���(�Iג8������\EUpg����M�-��ъ�@�v)8�:�E�m�2�B��W�iE{�ՊJ��vg�j��j'(�Ns�+wc8h�3�vBA�b��A2%�>m�Mbׅ�|��vD��s�@1�֠xE򑹮ou�X��ؼ�@�p<�f�>r�m�4u�8�v]��!�M]��:��;z�HE/����!MMBW�4�I��3�/$���=�J�ʕE��Q�o�t,h����.���#a�_�*ĳ1�=����Z�J%��K�O}J��J��:Y&]!��{,���K�/��X���,юaT��t8��5,p������F��=g����n�ϯ�����m=���<>����]��]���/���&qY7�:D������e}� ,�Ğ4/;E�e�옉�ljߔ�!��_�D�m�\6`�����F��K����9�(.�����c,���>!�^�a�ޮ[V5wee<� ��a��mhr�ԧ�Bfe���蚋i�$.V��3U�˃�!�S�S(p�B�5׏�k�J�C�����$h'���ht��Vu��R�t���'�������^]7Vx_�3/��Y� >�`^�[O��<&���	�@��z�^�}Z�aw�����/h[^�{z���{�EO)#�}kC���
7�?"%��oK$VOo�x���Q�͠:����J���j&V��{���{�S���­�g;-U�
5�z%s/F��Hֹ3 3�Y��\ �GB�{{~���#,0SX�ȳ�'M�R��T�Q\��@�[6�z�:��>��)l����	5��ޮ|b�Ԓۆ�|�sc���t�T�2Iۺ�W�UU^]�h���Y�z>�7�E�'jd�<�;�)�/�W
�ǚlY���G8֋��:�o4����(�W�HŤ1�C����j��wr�<��v:ѣ��]X̼Ƃ�T(���ZK��r��}R#�0�yuŮua���z�.�@
�ٔ��Of�o5�YՑf��0AZ)Yt�g�%�S;AUa������UN{\ǃ�����z<�WjyM�,{�u�䳅\�F��t���p6<�a�fl֓��ܶ���^,�/F%>(g�𧪣ʢ�Ҭ�	�	q�9��C�5�t7pY(��G$���G&\Z;r5y��s5Ҙ�7�a���q���J�bP����b���k!$�U��9ĪA�m�G�i�ӆ��ʄz���[�f�0��@cf���s�����V�^�IO��qz��/�����՟sV,oyL;S���g̋�s��d����nEڟw{WY�܆���K�yh몇��K��aíM��O.�+�w|�KU�����"07#��n��P:�M��p�����[K�PX��R��l��5���o�V���ͅ[}���,�6���$�jj�Z�'�kG<�a�����ZO��(���\q���d�̇)G҆�-�۷��i��&�  ��>��+ˁ�L��ҝz��Y��9K��4�7-L<%�'Pm�J�3OF�"�u�3MI�ʭ�|�;J�!�^F���]��o@�f��N�<���$Ň;_F�q��S2R/r{ŉ��Puޥ�N�y��#zji�<6�`ϯ��͕�ˁ�;���e�٥�ky>�`�.&�ؙP9!�vלh������ẞ�Z��\�Gc�������Z�4oAc}�y��VE�ߍ��>e��i�=&�CڝaN�c٘��T�<lz�>�'�Y���a��Wb4ⶄŝ���T�����ū�p�3���W�1ٯG���)��¬��������>���&d|<���;�݈U���c�=ǜ��I�������P������ܯڰR�B�t9X��Vˀ�e
�q��`�;Ǧz,�y��}�����P�NX�7�������.nQ����[jxR��e�C=o�gt�%M�^�mУ�
�D��+��,'��N�J�½�_1�[�x\���}ݢ�J�a̳���M�Q�(El��G+�1D]�/:�(��@�4
C��=��9or:m�]G�Č�e]�:k�Y�W\&_U�9�9����xր�V������ٜ�6�=Xl��ْ�.�-C�E),峽�A]βf�7�W��V�����#� �Y�����~�|&�!9Y&1PSp�q�Bk��Pdp��cy��`�[��6��r]��b�u#�S<ׅ̿����Tq���i�o���g��r�ɋ��ݧQ��0泘�m��{�"�&�_K�������̿SJX�qO:~]���e��6�꼌j�v�t���Z�K��H������~^3��a+��J�=;.��>j8n�z��!��V�w���y�T��6+��#Z�~^�-3�.)���=WZ;l��]�'�Q�8u'�Y����vu�����섮ާ���0��/��T����.���1!̕���d����V�~�E�G+e�>�f*f�SW��P��c�;H�U
[��^<�����g#�[��X�"�,��Rfo����e({z]%�
D�6�5�wz>Z���j��x��=E"v�W����˴�������ҵ�x]V�|D�V<��� �oZ>�R/�]vYmsy�G�� C�6�Js�<ֿٗX��5XR��mYJE�m1�I��$�/��Q���)�=[Nm���ܨ�`'�Y͸�:7�ޥ\�������ԃѾ�D�-�rJ�f�7���ʧ�s-�_:Ϣ�"���
f0�m��w�˛<đ�7�`�O�ܼk8]Z]�]�ɍ��/[ƫg˝'����\rz���6����cm��m\n�y���b1����1y ���cU��!��@Mv��݃�f^փ���xo�>��gFx'+d��#r"��ݞ{Z;�zl�ȪۗIv��
���}��u��^ �A���D��=�qs����cVX��Xpa�-6�=��r����Q�RXI.���z� p�l�c��9	��X'gZO).�N:�u	�����;C���h�fߍMpG���1ML��P�LF*_�>�՗�ol2���!E��N=�Po)+:�G���RІ�Q.�]�xR�/���g¥<F&E�z�V�9�7,y����i�@8U�ַ�q�\�5C���
߇
��{�ʕo8����x���;�ܺ7�n\D��^�[|��˷�r_aV zf��2 �o�"C
Q�k.t:��q�iу�^W�N�y[�%ވLLU�s�g�!a`��x.$�Z��=�Ζ�%������-T��UB%+#�י���mh�ݕ�S�������\�93�O)�w=�~��#m jf7U�c�7�>T)�Jv��l�D���3��(�er��B������T�lM���>U�N�k�<�Ģ�Ĝ����2�Sq�ܝW�qcp�l�ܤ�̝�G�H���{WI<��F�p:�vN'>���U}��gr����{X��Z���Fً�E&�f��՝��+�/�+�r��s�J�c7ug�K�FY C����NM�����6�>��Y/-��
UL�<%<̿$"z����ى��y_e�+ ����`8)�o����~���&+�]:C6��؋ڋRN��+,�f�K��^��W�Ҭo\���ķ�wYKŚ�3�f���O7�:��J+�'	}�ʋo`Z��U�@<�Ɵ}�mA���k�5�c���e�ݢ�������w���^��ڢo���Wz��%d���S>ڨ�ZC2�s^����uSe�c�mehݩyϫv��t����WÇ���+Z�S�T�{�Y���\�W+0�:Y/k����t������%8v|�f�v<+�+-ό�+G��__S�jD�K�vo��X�Q��9r���]ҌsM�F>�V9�3H���j���EVz7�''�h1j�f��[������	�4����pN55�G�E�J��6�m-Ή�w��[\��2눣wȃ��z���+E��n�} �O9�/���a�5uc'�ܮ8ʳw��t�SVl @�81����J�٥��*|�S�m)��ͦ;�ӄ����A>9b��+6���:|5�N ��8����ۨ�wE�9t�d�$�c����OVo(;��Du������3Փ?b�結����sҘ��a���3`\'R�u��I��0�^.T˞\�fw14�[Hu�R��]M���X���1n��F1�O-�a*��f�8��d���3{(�R�kdU�k4:XY��֍2��t�L�P���eIǍe���wU��[.6�.�zf��"Һ��߅�=����`�Sz��������I)^
'ݹ���n�̝�٦"嘸d#s3�WLߩWg�lu�Q�C����]ϙ֨�OZ�qo�2M�8)�>
vĪ"ב�=»/�ދ�au�V";�|�Z"��^���.�q���z[�ͅ��.�NEf�/�T���Q�4��ѯACKw��ޝ����:��0�L=��d��򋉿be@0�6O2��yƂ8�s�eX�u�tl��p%�ͬ�4ŝ�a綶��:�D^��[I���rU�J��7�U�^���Ꮖ�T��Ĭ�zˆ�YG��c\3�jA���:o>j�F�IT^�Y��c�;�����ǡ���0^��Ȥ;&@jH���̢�g�q���̟]�++�K�6�a��p���Znr�8�ܴwsh���mf�1�N4���O�@�W������Mk������˖=Z�@�jŜ�؍�|4�=����舢WcL�t��&>��WN�u�3��Ճ�kQcn��l�*�������xl�p���5xoM�z��!�Q�qYčN�d�}K��L.�w#Ag�Τv���r�)�g{%X���Y�����3��[A��P�(x�޷���av[ܠ��B��ꭹw���,��PZ�R_��ݹF��+)۸"xt�b !a>��|����;�lx���_\��s;��W5Hϊ�IB��#�|V|C���:-_�zρqsE�A�*`�6��n�ڹ��ӹ�7�v��I�'�*�/9���PeU���3O3[��Y��Z; Xn�[�"�i�]�Wb���s��	��ť��N��P�e�SJX�qn���%���EK7�xl�5)��l�S�������u�f%��"�C\�ԭ�5�Y�2�g�edvqI�ujj��T�pq߷�U�⦙����2/\�y�*��#���:������tƁ�t�&5����;e횝�p�L\g����~��8j�tUg�Zf[�$v1c�&�Rz/�F8�Y���as�T(*jb�'�ú��٩�`����6�G$����:��S��YlMKb�'��h�]/K͵R�OY&�:W��u�b�+X�;z�F�pdgX�S���}��9��.nۇ\����S��.�'�q�QV��]�n z^|��yA�c&a�p9��-���{�y���G*���H*7(;G�#f����ݧf+���r�u�����]�u"\:i�p���WB]���ې��dHu^�@q���W/b�W��c�Ԓ�ӣ��.�lsmuѕ���1��'u�7�r=?��u+���R�������8{&`��:�<���u�%R��]��Yt;���g3���d-8�T�:��b�Ԍ�̈́���[� q���`��M+���́�̶�h���qG�՚x�5�t�꽜v��&�p�cT%O�#�j�sk��B�]B�kfL�;��hL咢[nlbC"ۉ���Gkwa,����V,6�	;�O�+��m�Ʃy؞F�W�� fu�/a�h
�GPu�,�=�6a��R^�(Ck��Y Z�v�6u�+��˚�Űv�5;b�겺d1i��m�9�O��^G��.��uc�8�t�]����o��P���jH)oV��c��5�؆A}:&�X��3�
}M�l�\n� ���J>6��V����}��5��@J�*�Cm��ˉ�N�)��n�SW�(-��Ïn��"�i���y�+�]�n(j���@���G��(��G��(m���_n�ZO�S:�]�{7�W��;�x�ٽ�(�u�s�vZ�S�.�7����­[�S���N�����7_Bc%Xꗷ�9�)�;�|��Vi�t��$#qNr)z����uԏ_5��j�BA���Ǹ���l�x˗}]t7��;N�bs�ۉ�9js�+Ii�`[�0�՗���\��Vrr��ڹ�����k�ϙ:���Ŗ�(CŏDյ���w�a���΍vK���A�$�/;z��8��	�� �TVkh�N\j���\A[�j[�!�u�577��p��%�f��
�A����`��V�ٻ��U�(��H"�w���t��]9��n��v�튢!\�2��W������\V�;.�N09;:̚�H}�r�h9:��0U��E��Y4�
-5���j̤��]������^�yX.z�)b�̘� �u��Yá��d��A���5�s�	2�<1�#]"�uàw@0�"����rEc��8���S�>X�Z�mh��0 6�n��B����؈I�_�YxyX<��u�*xi�.����aS4��[�=�$��f��j��=V�4RDa���:��`�]�p=�9h���M�����EDk-����k����'7M�k�89	C��J�3�{s�\4Y��?x���y��4����D�H��Dk32�L�*��)�2lĠ�+3���2���
�P�Ha�f%�f����Y�d�a�f5Z�&�XfE4e�fQY���U�Y�F�P�fa�8a��e��k#(��ɌȌ�*h�3#��� ,�,'2#p�,�,��1��
���3Z�dVY�UdTeVa���efcYc�akZ��XDف��1�9��0�cf3S�RaA�$����M�0�)2232�2������$�̫2�0�b�����a�QQY�e��QT�E�E��T��ݺc-����	xz���p��+����MO
f0a��`v�m6���m9w��P�J0��(i�ݫ�+���m]����y[�pjDN̂7��!��þ�Z�{�6xR\�"���z#�DYy�N�����ğD�1(s΀�(!�p� �8mm�y�L�qAl�$a���Q�5[���l�-�n����/�r1���xG��ʸV��8;j�>C|�f�Ut#�/
s���yq*��H���X:V��ɗX��j��a��Jڿ��R+���Ah��\w����^`0�����ѐq����5Z8�5�#�G=Tbϣ(b�i�l�*�{@,>���wke(ި�j������k�ў	��1�[���ߧ��?T0i�SՈ�l0arv�ksԵ&y)�(_P�����2W�9�C���Xjw.��`��_�={�ݙ�ǯ����f�V�N�e?0�T$��l��F(g!8-�p��3.�F4�y���ǘ�������LtEh���c��2�WY�|��^&�Zr�_T7K��Y�J�ߕB�P_
����X~RІ�	D�	v��J��];]cÈ/�i>��NXY�Ɍ�@/8hm��+�uϩY�R[Ǩb;3�g�T��&p�}�@�%[hǆ�cJ�Z�c��@�h^^��;����87�Ŝ��U-.4���_R1kV,����woU�u�R�tZ1:Μ��fo>�̓��}_�6{�(�;��Jm��L�|��3]B����t8�&�y� $=2��ylIV��Hg�5�zI~����N�$�+cV��o���]���/�RI0��VM�t�8����\�F�]�z��X�]>B���P���{��t�u�R�hYjIN���xX!ъcFwdKȉT6�; ��g�^q$y�>%�µ�v��6�-�!��O�y<����"{s�H��L��Q��;������˧�𴉺�Dm����I�\5�,s�Nv�9��f㥆�6��Ē��E%uOط���$h7�+g�&��(}U�z˥����vxJ��ɢ�V��=R�v�ŧ�/hK�vin"Xj@N% 9�7�b�s�[0�O�<+�0f��u©���S��:Qg)Fq����)��Pw�?#�<���:Y"�^,�Y��5�YxV���������祭%^N�V����G��#��5ӎSK�ɖ�v�:x�uƍl�=:��s{}�y��vò''�a3�� ���}�-!�v9�]=�Bҹ��a�)z��'6�R�Y�9�mE,{^�<��7��R�f�a�
��E��}����jW4!��4d�2-}�R��Q0�w,(����"�V;�Y�]����tB��}D��,�&j��þ�Y[��멖������Iv<�=�s{�_v�����a':`���z�
��b�B��|���z��%Z����q�N�V5�F�#���e��({�*p�7��n}�&	A���m�J^z���z�ĉK�� rw��h�9Prh��٨��G�0N55�D!��MƆ�&�ƺ�E�6��:^��m�a��v�v��ˍO��=U���]YF\k�'�y��N�M{����aiH6%4��'+fJ����y��0�F��&)/���aq��΍ڑ�y��1u��V�H#�g˩�w� ��OV�Za�����:�y=��S���T�a����M>��K�Tgr�}�M+��k�PL��ϐٕk��Z:{�w��e��=޴׺L�&!��2a�E�>oL���B��u�Y�w��[�{o�����C�q K\x���w*��4��:*�c�a��r�l���Hk+RMi��=`e{S'���1��Gf��<�:o d�UC\�,r�h�pS�|0�˻":�lOp�ċӏ�T̨�.����bƕ��U��6�(+$W�������	D��Az��۬�W���6K�w���5��݈�R|���MwT��V�E���>]̼�v<�K���t݋*�ug)%@����M�����9��*�Eu'N�.���ٵ�	�F*ow�+>Y`�
z���d����R���hΪ�y�]�c�EmAKǲVZ�,y�"��m�ƥ�Ņc���;��c���2�ղ���M��fL`���q�سHY۶mm˃᮴�ނ��c�iqcλ�N�.M{�z0�Hp��ߺ(v�S�٣n�l��c�#��'�J���"}���Ūƭ1a�1Y[؏oM�ƶ�	��2�w���=z�J��=e����M�e7�SU���rE�|b�u'��QXf\F��)�F�Wf��k�`�av3���_�`����C��gL���xp[r��D���q�bcl3,S��	�f�<]r��7(����t���y�<Q�,Ճ*]B���	���D,'����|�
�q|PA�X6��j�P��ј��\��(r���<.�����|�~Z1�j�>���洊�J�d�1� L���cH�!��&�e_Hx�Ȏ��*<<�6:%[_��L�,�< ��N#��5=�5pIL�S익{[�W[,�s2��w	�yԾ=�Q��Y78ŋv�m�y�Wa�S��a<`|+#[]������|�n=���h�����lF+	<�spU��鉳��3hC��"��Vs�t>3������D�s[x�������7ܫrv 0�lN�C�w@�&�a:��B���iK�uҿ�c͒������8��!z�u���a�=.����~Bx!7(@Et5�_�+g��)��V+�T���k#��7���3Җ��/��ǹ��Zp�Gã��K� �*����j#i�#Ů�3���Q��ux�99�Z�%�rK%�c��m�$�D=�{�k˙�:D��RN�n�o>�i��mԗ+eU�<���"]o/��{A�!��nY�w�-Uso��6�<`9�&e�K�,o�g��N�=��,sۀmS�V��T�\gf����'$��0�[W�K�}�˃k��j�+	Ou��:�؃8+*y3�vմAb���輺8w3U����zr���"׎��1+��֟���6�u��+���mA�Ym]G[Z�U[��xopW-�EAE��ϧ���cFA�yq�9�G�zc��Q�^{��p)/<���oG���"��w�dPe����~Zp���dw�/��:u�ZWzV��33�j�a-J��h��'�تb�M��dyP+�"4�d//�tB����q1 �|tr,>�S`�B��c'S��>��kЧ�5�����)Aq���Bn�f�W��QF�>��'"=]M�Fk�Tf�n��۲�*��!p4g[���P=���x�~> 7�gF���)���k=ᄿ��S�]A���HBst�,g�����K������]���7(��U���8>���U��Iq��&��BM�ql�tb�tÇ�ˠ�\��5L����NN�ˎ�L�Y�P鞹aE`%�v/WU��J���e��4������R,���qu���⤩���]�qV�N���Θ�t
Z�Q.��Sqt�&yf#ț���,L����r�D�p�O�4f��r��{wP#���QD�G��F�s�=���]��YBzQ���Z��y�Wc��o$�\/�X��������=ɗ�1����'�2�(>V�Ж=׺���p�߂��B�9�9%:fz�vs���D�9���}}WY|+L�V$�IK���GR��gk��~\���A��X)��y�WaY9��r�=���'{;�N�G,�^ok�gˮ���(�/|��1yh��ᬱc��y��>��GAv�tx�y�^>i�����`r��K�3�>k.���'��J㛗l��x��)���]vd�2�pi_
z�¾f��s.��V^�A�t�Y�ٶq�(��$��S4���c�_��rBG�)�y�U�[���lR��=��enu�0R՜;j�+��O\���3(�����^7iR��w�-��Z���P�d�9R��Pwr뎊5��H\���+�Л7�.~;�E_��ī	��6�I��Q9`I��}2���ؔL�ksM��}�G�'}۵����8`��X}Jh]��Ptc�ȉi�[��/lQϹ����O;m`ų<Z��D�c'y9����b�L{���������L�{��O�'&l��d����j	qX�P$��^B�Bxa9<�&%�X���ۭ�2csʘS#��k����ݜ\�2�q���\U�v�j����A�;4�vM�Za&�]q~]��e�\��V��?=�ll]�P�b~����ɂ��J�g�y�/躂z�ča�c|�K�W{6�o���!2֊����u��Ʀ�Ȅ;���e4=��C��8X��ވ���(�u=:�R�ߨ�bqJ:5������O��S�X��aи��!�]���cx�#�DtW���~�T�J��L��d���~�Y�ޔġ����bwD�%�wF�5����TM�M�+��8��b��#ɴ�1�L73����p�����1F�We2�P�K?g����	3z�Ŝytw�3"u���/9��5ìuu��@���'����׽�Y��n&*�GJ�۫�.1�V!�o (�UO0C(���l�"7s�t4�!�l7tOp�[�@6���{�Ցұbn�Ӥ��\�������5�Ͻ�����Pn�}��\I��UC�EG�'�W3Y�CO�^��e�3'i7��&�pfy�-΋3����k�<W������H���qw�z�.��l!�%�	؝s{�]��z��q��ܶfEw��k���B-O��Hc���d�i���-�/���_H�a����@��:�����%��"a�:���>�d:��[e����B�I���<Q�T�qw���;h���7��V}�VX.�-,��^6aC�s}#�jWj��������=Q�V)z�y��]�SEj~�`s�hj������=��b�d��\��'M�:��fq�|L`f!P3�%�ͬ�H]���G��>�u��i�9U��a����=]����<�
��ފ����S�V=+#����*�x��v�v;<R�q�\k�6���{�L�o�����Oҷ��3:����V{�.�f������׫o1��g��*_���'F�x��ɍ6�1I�7�[0q�k�g��m��X<��g)f����)[�fW��p-u���0ՙi�B�@(�7 ��݃�������z�~�ۯ^+8bP*� LÑ��:�pw�zu��bOY��*y��z����Kmub��5��z�kB��̷[b\��\"�{$���N�yJR�%ֆ��v�&8��E�.2Wu�݂�
Uu�&�9B�l3.��P�	�}�޷�ll.�{����y����/t��:a^����-?
T
;1/i�;>�D�|�
�q9x4PPʡt)�Su����7I���e���t���ϒZ=>i
֗h,Wx��|����[�������o$��P�7M2���{'���N�z-���T{v��eB+j�d�ē7馵�gm�֮N��g��v>Ȳ��*ܝ�¹|�D�z����KZ[�L���˔�a^�ݙk�����"�k����wzY�\�x��rZ3��yQ0#����k^Nr�]�I>��yX5��9 ��3�8�5\<3�;�p�.}���Odح/���U;M���@���<�u�o�O#����boVD}�Ձ�Vx{�;ڞUo�Պf΋�cUm��mb�l�;����˯ZC�0�r�]��T��"�%@9oK�À���Ꮻ~�$������0aV]d��"Ƅ8������������-9U�Y�&����|��,�I��\�\����r�fb�ףr����Y
޳�C���Cu�Cȴ{N�Xfe���2����z��}7��j����Q
�o��]*:+��6�zz,��/��*�J�7��>fGK)s�]\�,v�R_c��4?U5��{�{��7�DNٮ
�3.�;>(WX#�:�xk]���n��(S{Xp�3c�� M�+`�L�Ұt�����پ�V|��F,<e��^F�Ώ�?pe*�T��~��	��_їD%�lh8�2cˍ��j�qkVT�Sϰ։#w��&};�~#;��{���R�^��WU@x�Ac=|_���i'����#r���Do�����k}~�z�s��0i��1�u��eel��o�.j$�qp�=�OJx��,�7�Q����q��|N�q�޿����*�L��>3䖏J~`=> 1���x���ڵʙB������MK��	ƙ֯�������v̥����*��G�<�4�c�����6a��X��&N�~�':�q�ެ�U�!���hǎ��=�ƏV�(N4�ޞC�I�pJ�2�*��qX
�i�`�/�i͔�ު=6�Y`�}�+.˾f<ط���̥�
:_��3�]S$�S�5k����|��n���/�*�����>n�]`�*?a�ǔ�6��Ƕ�45[ѩ�h�͍��K��D;����k�P:%�j���[��wh̕5n�Z��i\����wj1��UF���U��ü�����]�:]�����H͒Ћ���3Qat�a!��˾s�M;scwv�����Zs����p%wvȝ�v)4oKf��Xr:��x5�}����g�z�]*1m�䌳� mC�Y®��YYK�xҙ�2�uΝ�&��wK��Y�g5�us�G8���iq�:z�Mm*}{w����n�yVE�]thhp6�V^l��)P�%m�E��}�WF�KN�����]�k� "�}������.9ӗ�O4Ƀy!�6��`��:y��;�ȥ6\)�c<s,�`�7�����U��`��գ��":��'#��.[K96�u���zs��~���;����q4.7�J
�nw2(,i�딓�X��G��Z�]��vo�]��� �3@���ؕ+����Z��1ӰW��(l�w��:.�v<�����B���V���q���DV��A�w[da�{���ε;��:(n�t 7�ӹ���{8d�Z�S໪��f��V�c�����ϵ�haen�WJ��w�]U�M�>�W��2�g�9��;U��!�����ܐr[cE
ܵ*."\6F�%5S���[�v��ys0'��:`7�h9��ͮ�YvB�<�o�87�d��9������nn��7�V�gv�[�s��T����wh�B�	�B�k��e#pfh���̘&C�q�Ǔ�z�h�2�&�s��M�i-���os-�18]n�2�FV�p���P5�	D��$��Ô�M�O9��f��q�1���S�Zƥ{v�X�_ �VǴ��N�}�-b�×����؂f�
u��X%��jlp͗�sn��v�Ι(��x�a�g;%m��8A��Չl�{;�E���Z��7P����\T��N�N	ݭ�{�O�dmp�D+0�ӕn��MU�|��X��g�hR��]> ��Z�on�NB-��Q��V<�;�Vf���;� ��2���.xۃ��Q���څG\��k6R�v�]µl�r.ʗ�fi����Z���fcg!���]ʌZ2WS:8U������a�?��䠾M��E��d�#/�P��s,��͈\�
r��w�ܽ�/����4��Y�j�vީ1i�yK��'F
���%�֠G�d��Ruh�tњre�WKm�v��ؓ�D���ˤܡ�8i��n������u�<���b�<kesP��_r����v�m5����V|"�s�6�!҅â���ã�J�Z+u����ec6�t %l8�PtI�w�H��&���nL���Fd�d��*�����dϬTۮ����@ 2ަ��}��[6t�nЙ�Ew��6oC@�k�F�r.s�7�����8�G;m��4���2�k9'�t�nrT��m9�yp� 
Q�~?�ɂ-̣Yac�U1DUfc����TPA�Ee�EFE5�NE1QS��f5�3Y�ca5FYE%�TXeU4�Y�U�h�`A���fQf�Y�dQ�fU�5Yf4�Y1��eeFCDY4�&��'QYDLE��-4QM�e����f�FXKFf9��LTU���3\!ɳ(2(�2���*����a�0j�2̧&��,̉��#
31�D�46�"����$���(0�#2d�'%�b��J�k1��i�%���"���3
L��a��' ɳ0�irX詈��dZ���C�Mk5Y�Y�e�Md�UFfX�Y��1&N@VNM�i5~�@G�B �_I���.�y\�k��C4�iS��I,�]f䜮����G�d��{�:��nq��!�L��!#�����=�WT��3(��s\���Y��?��)h�8��h;��G�1�:������	�3�z$�,%4"�|#<���΂ݡ���I[��7T��Vgk��w��j���y<t��E�a5������0����1Z=%���0\1]R];��T�"��u�b�8�qA���]���㚽�ݫWw�&[����̆����$h6$��������%dߩ�ܻBHEc�i��w+toN� �����N�`��3&��7҉�=V/>7ըLc"�'s0v콈��ew���f[�V�>�.-Ŗ��]�o\q�"Z�I������D�pp���~e��t���a��˧��tO��ZsƜ�녍�����3ã���ɖ�vT����ϫ���Hm�889\(^,�b�P͢j�ٛ�tŝ�p0h�컎Rb��b�Y�����{��^�����7�t����mז�5���V2�`.��*������$;4me�Э�O�����2��
ͿS��A��`���v01�T�����]@�W��Uэ���.<�x��`>9�+�2)^��>���8�v-���ݧ��o��b�w+MM��CK�ݠ5�w�3����m`�XυN�WX��Z�tm��գ;M��{Β6�u=��[	e.��R�8_��/x�p�Jf�}u�O*<�c�]����x���/ԦN�.i���u��Ʀ���w��eq�t*��j<�b�9^�3[y���60{��`��f�ce�0�';���S]d{t\TQ���td	������{��-�b�Ċ�-��ع�7��{��_�r63Q�'ɊC�5:�]�{9K�mۦln�H��!ŞH</�yu6�����fs��ڙ����ު����H�����Rb�xN��.$�ڨy�
	�B���Y讎��X`x j�§�wݗ���;���\N5YӐ]31@�Lɇy�����ZV*W~p���K�q�gQ�޽du�i��66g��wz��\/"��p(e����<,O�t��'�wԫ�����r9�`�j��4A��{�	B�
���C��z�W��C�݈`��ԗ�	��Ū�Z�Pge�N��1��;lfֈ'5��n����6�VL�s�5#�u�dnV�3��i�V���L��n\O��w�|Ej~�`s�h�y�Z�J������N�eI}i2�9;���ʉ�=b�.�I,��1���dk�: ���r�Ω7X��{6���"��#��Ѳ�(vZ}8<��p��Va۠�Y��F�g5YԱ������2�,�WJ�gr���ew�92�<�{V6��G��C�`wVM-GWӃ��@�q�8ІfiY��{6��L����5e(�����XɗR_��Y���=��8+iz���^��>�V�k�C��dѲ�QCb������x^=�I��/$�z���Da������F�VИƝ���u�'��Ճ=kYbP�Hp�l���xx�}�t�!����Ս�c6�����I�5����.�e�����Y鳲Bnq�� �z��_Og�i���Bި�e��;�o����q��޵�������;#[�vߩ�S2e�����K�H��Mz�k���*��<e���O����m����{,��;/8��gpg�\v�0��g�zE�	c���Z=B��]���=U�h�{��c��r;��S�-gu,��1O90�W�b��=��i4 S=���/j�y	Ъ���v�<X�Vۨ]�����:�Zav�u"ۺ�KA-�]�U2��'>��=��'=LF�L�r��ˮS��<d�9-�B~�a(t5�W��J~Z]ѿ+�&nd�g8���i{|{<��I���8�tQ.{�yr��N:f�^uf����f���{QHӖ�B��,*�:j�ut���Vm������X��s�9)wXu��,�br��z׷F����%�c�����S�[e!A�'r�_R;�Nn��3��궢:h��p�x�N��g)�7���57�
6Ƙ��uf��퍘�i�ůT� C��>��:Ү�,<��硉��᪘��VxP���Gmy�o�{8֔4����E`�gԏ�Hpܫ�+��[.��f*g�����]ҭ6��rs���G�(�"]T<�U� D� ���2YWʞ=�e���i�N�����y7��}Io�PP9a�a��Z�Dp�#lh���}���/�ϕpw���#�g9S��ܮz��*�f��/���U�I��+J�Q�|6o�U�|Y����rwFQ.u>�*$Q���q�V7�sC�FF3Q�;�i`��κЃV��Ħ��{=�; ��m?b�%-u��xR��}BP���?�>�u�:2r�N5lF��5�Z�&��ޚT�/�M�T0i���z8�T:��
}A�c˚�+�	�#u�e��(��X^՜��҆�,��J]r�i(̪J��I��~`'��P��7�Y���F6=|���S��� Pm�b��=��;�y7*p��h3�H��R�mr<�p�딹\K4����-�m��K���.�*�yn�����ֹe�����u�)J���
�����Z�z�t^:�ź+ys���v)�[9S\�uA����1�A8�:�}:g��
+	r[f}KSA��T���aB�z{��=�y���ܑ�����L��v�':�k��<T
Z�J%��ڣ��1z]�y����#��8v.'���Y���o���B�|j�k�j:��4d2�~�:�MX�@�ޥJ�\z����LJvƧ5���62��k�������:�\�O 4=̛�D�3�B+��׺��p�Х�И�� ٻuݴ���F'ϺU��:�[s�	^wO�x�$/���-.���}�l;�r��ܕ��&�5�ZD��o*�g4��.:n���\�&��O�/��|��2���M.�,`N�J|��)����|�:ovv�~�뤯�P�����$h7�+L�������9�d���7!�}���
�/O��k.�_4�7��x{��I�҉�=V/ 龭Bt�[BI�R5(��[����QS8K8'y��*�xYj{��iW�plc����<���v_����t�%Qº�������4�V�(�4nc��H+	�,��ů�j�kn�0L���h�Z�E�ǶK+�5�]��]��S�u4��:���ڨ�A����Z�F�~�!����F�5{�
���ˬ�G@9o���-��v[l.��Yz�����`� �վ�ڿ��2`��BǶ�3�m1�C�����tX��Y�xv�~�|��W�QW��-���Zw����&&O'~����/Ph;���n���x⬣rϗ�3��ݢ�pS7�ձ�:V��Z4\F�l˳X����sf{��po���S~���K�Ę=u�Sua�rެ�8�����?o��,���K-E+��n��,�d�s�lo_����R>�N%��α;��=��N55�D!�~�45q������1wr���]�iʀ>�W �ع�Iuz�]��/��x;�תv�G����s7�եj��1��niG��`����DtWr�?S�J��3pl�0��9���d�iռ�y[����.nz�N�\I�:y8�]H5+�����z���]+u�R�[�S79Ol�Y[��a��[��d�0�͠_��&��C�z�d_ �̭��W�a�/)���9�#l�x�}C�ؠ�Rг��<�%��&�9H��T�.�~�N�77�����Aԇ��	aT�S��̪%ތ���L(`&}���qڙ�`ؘ9(�udq���Ų��vw3/ީ+d�*��s�����^��hoF��;T�B��rb�8�O���%�L��W���.n�i�bO���"rE����{Vr��XKV�k{W���I��joV}O.�]ø2��=P�O�5뤅�5�@Շ��I�����\�I����L���d�3��C̪h�
|��P÷���!�ڦwk���0�i�s�35H0\FE<��o}v��;l��5X�۾�Y�Y`�pSԩ�����Vw�"�9w��,ޫl�E%y#zj��j�u��}��i>+���M?m0�um[$;Y�ٸbrNP�	�f����0=yƁ&03�@�ؖ;6��!q1�^,g�C��kvN��͙�9�kת�u��/x���0'��{�ەY���(�K*�+�����i��,�X�Q��:��˾�2��#n�{���(1��>Wj�3�O�;�dҡ.��x�>����HO����޺#32\V�M̝6�4�#r�[0c���J��	���^kY�ʱ�Cz�%�y+z�U�.�H�!��P��[.��i���N�(y9c���M��<�j��Ĕt�v��{�A��)��SE*E�b�XLĨysMxc�,�/�=i��bϕ*+F+q�y�ػ�b��%(�vy�jς��8��(��^���2��Ó7ʆwHD_Z�^d��ř�wʗ:����r���:���^�
��E�M��T�`B�P|�++"�cw�����j�$t�x�Ss�9�]ǉBt����Ok�þ����`>�Z=)�+Z]�X!��v��,��;���J�~��#�x�0�Rb
��>3Q��dʓ�H�e3� Y�<�ˮ�;[�νV�s�1�ᔄ	�nV YfL��|'�����av��Ԉv�z����t'\_���ay�Z��Bn-~5�*�k�`�D�ʫP���<<�d��0���X}�5f�^\��z{m��j��Q�>���qq>��y�f�W'cg�S3�S} �cP���,�/V+uo���!��#��}�ZU�e��jyW�/��k�⻚��V�Ƅ�q���\�W�t�H<.�Yd:+ah����t�9[.��k1S4�Yo���9�[�h������SН�|�`�V]d��"Ƅ8�] �8�X<h��ŭjΐ���	��ݒ�RY�PRKr�֥��W���|������U�;�n��7�M�T(���~XwDq���+BH�=oD����kQ�:��͇�f����{��x���a��'�fy�%�h�����l��wۮћ�+��=�<����#|�4��Yś�=��±���PɌ�-W�g	��^��ȫ9��lL';�M��[���T�R��:X%erPSs����/EN�A�W<�ԗuI]��p��?Y>�P��7��scA�&����vs�V�'��]&��Tޮ�j	QX��ڨşeTb�/��=K�]
�S��t����]���x�Q8�515#��p��t}Z�[aw��0��ڬǣ�z�����T(g���!9�N������m�EH4��sy�W�������r*�L.8���O�OW��Au���w:����i�w���^�u@"���rެ�i��u������d�;fR��DV��n����}nh�omAU���1И�1�.�N�~��C�N5�Ց������\e{��Β�[Y�=�2�.~����\�b)��1.��qX
�i������yU�\���Cj֬{����>�����D:D�OWz��������HN���y��F��.�I�=�\eջxq���m�q����9̀;�޴(8��h;��{��.w�+n+	�6��.�L�-Ƀ���L�\��g�����#�)rVS#�_��uT�u�-8�M��y��l
�z���.K&�l1<ɳpkm�K;m%xf7Ԩa�Q"��:�e��e�U�k9K]ӭt����qw����K�9�xSw���L�*	˯1�k��A���u�]|tn1�T'�K���\�5�nL�trģ��N��<�=3N]�[;�k��]�Clӭ�a�9���kC�&�����Δ�b�J�*��Y�F�6���ZO,h�E����C�����4�JX�I���]L�aD���n�0(�K�� �T51vȫW��fR�J��y��a3&Áp���r�TY�t�˭kh�����q[����b�MӤ3j�#N�'�9jytZV�@Q�q�<��;/�����F>F����C$�!-�1} �lJg2e_�ڠΌ[i�g�d^���z��A�!����􇫵��=M����^4?�ܴ ��yzD��ᄹ�����Z�u����е[��踦�V�/e���ZV=�ܭ�i��鱨a>qX�g˖9 wks�]�Н�ʷ�
���q�� .2�5��,	��`8���ǰ?o��e�x�)e��M_k-r5}yϴs'���T��W4���R%��Ͱ�'�A�O:��C�b�e)�y�*κ�K���;�5Z��(i����Tz���4�C76x�o.40bS�y𧪯���c�o�&;���s{m)��Oz����r�4�Ŧ��䍜���+ ���o�����/�XV]��-����.sX�_@���k�)wV�v���R ��B��}۵��i0�x�0�[S�ܕ��S�ë!�����k�+���F�^���h�XtV���vU�ģU�!���84kB�{�V�SR4��`���j�e���N�3���,=[�܆��%��Q�vh�@�nS����պ�p�co;�=2Rr�����+�q���v�!��j�aS5���T铥N(�v��
Қ���@7���&��EGݸ�,�hw19V����ںE�胠�zYޏ5�uP�M�w��ȃ
�Y���rݫ��M�	ᵺFȠr50�e<s�ska�?�!3��Q�����Wf�z;�2�%8r�A��]΃���� ��� c��u4����N�-3t89�!j�\����}F!u�ZܛSP����롸�����e� �\[��w�)��uo8�\�)�hM�s�w_>ۑ��΃���N�Ԉ�q�Ӹ.���HhG������خ�̘؄�3�fmҷ�n��Y�
�;���h� �������Fk%+u�\�ZxP�KvA����A��s���:j�m�J�����(�[u�U	Dj䈺J�"r��	��I]��Y������d�II$���;B�'�c�-+3ؠ5�����h�¨7�c3��W���&�B��2��v�����xc7����wd�Z�Ov�
�C���P��
t�#��4�Z�c9��i� �Xu��y*d�WR^_e���wlIf��q3�(g�t�)V������ *BL�4ޗ� �ln��'N��\�l�}W\���)�Ým3�Z��0�U�T��W^e<��D�wv9sF��-��):ڙ_�����K���Zu�Բ�N|m�����s����è�
Ѣ��-]����Yֵƫ�� ������o0X�vFV-�!,7�Z�V^��`�t2vqhQ�y�.t�-�֐;4(�B���:�wi����N�a%���]x����Z�Y)�6E��)�r�t���aZ�=\�;y8QL�QYG:��
WU���q��ow����K��i��/	��ko�X��V�ė0�a����ѻ;�_U�<�����ar2VmBlF��қ�%K���3��,7j`�|mo+�Zx���r�J��}3��I]�ES��{Fŷ*�#}�+�i�V>j�\� �Ѣ����ϒ�Υ�i��P���l]P��;�PB��j�".6dd���r�9R��,��>w/l�&9 ��25Hg�tyZZy���w}8(�<�%��e-�0���O�г���wBZ��/g���ˌ�X�5a*wv)�N�;d�y�ԓq6�9x'q���l��d|x�R�Q4�Gx^-\&�ݜ�����yo��9ڠ���;z�v̎��������gq��V�a�&FAY�a�0F�P�Ѭ�3�2
�8M�R�dkh+-CC�#NQ�DčjȢ��Y�SYd�aE4CMUXD͖d�C�KFDE%�fXUC��fd��YPTK���JVY�dc�E�e�aT��U9	C�Y���Q,ATӒS�RRQ�FI�Bd4�P�6a�Vf3Q#K�d#E-I�abE4���`�3��C��a��E3R9S�d�+��RTKE�%K���ѕ8�!�NB�cfR�AECT�A��fM!faRRSfdSU�T�d�9fRٕFYY���e�fd4Y�IH�.I�c���XBd�d&NIII��Fd�$ANffC�d5IEENYeFFf9������y��a+sh�̧OrR��ޔ�����|H�bd�]]�'w�ok��R�έB�T��#�'ë�vw]��� �"RR�Q�s�Yemq��K��#��r�w��|�9A�k 1q9�`O���y����s�k0݃�;#C�w��<4
����5�e]ǰ�~��qFpu�����j�Qz���]��jyy�V��C��IC�mȫ�A�u0[�.9w��j:�K�^��;�e\Ň�2��B�7�`Zu!L�5���y�q�S��m�%��X7 �TTк԰��yM��yp����BZ�|'���f.Rn�`���"r����8�v�DG"}�G�7�_֦��*_4=(�,qSV��V��a�w+�;Z���p��w��߾X��C^��n�ً��;l����7�[�ͅ���̱+3������%�{����a�5������&�'����/��cR9�a�K��x���`��^���m�Y����t�ٝ�>bg�e᷊�\&%��Y:;76�L�ўW�Y�����/y��1�4����}���(v��F�TP�
�������X�v5���f���cӎ^r��q8E�����>;rC����4�Ҿ�ta{�XP�;���um��#�)�<.c�|-��{�ƴu��`�i����}�v
�P�����v*c�@�5*�!��p���`lL��d�kp/��X�B��uI����_�c���}xg�wdo�;�����Wj���vi��ѷ��y#�9�ď�޲jȍq,B�����a�1�I̝6�4�#q����>�P]0��+,ޝ����N�b��f}��~Ԏ���+ !}Z��9Ԃ��;�o����q�\�&�,6)L���L?��[�����[���]�L��m��T8���֙�P���d�J-�Y�[D��^�{]T�+�U!K��ƾΝl�����<�#�C�$%����Sk3����js�`^'����mO�h򷏽g���N+�!��c�]�����g��A3 ��	��Kj�Onf�������q!�B.�2���3��]γ��@'R!ͻ�prip����C8;�x���Z%��A�x����q��OlB����4s�O�;\f'����ޯ>U�M�����@�zj%
OW{�B�����ܖ���ؾ��p���_�l���b����=����gAo��Q�º+4����M�A��u��5�l��;�u��y��ޏU>��y?`;3_jO��v[	]nG�����:4w�<�ӓ���`!¶;��gT���=�)@���AT;U���IJ6�oe��.oE�d�4�ˉ�n��wV�	|���4���v)d�vB��8ۋ/i�9�ؔq�d#_wu�sb����^��ƽ$\���[���ۮ�����PT����Zy�J컊�~;HE'v�jt�'@`�n�>U�Y/:��*g] ��=���boZ�Gw�{[i��T�8()��6�5�gJ<�DN�Y�G��(^�[�q2�ypF9RM�~���(2����>�q��^� M��_�6�Ns��0֣����z�ܻ�較�J=toş+"/ňʖ��fՅM�C�����ѐc\n�.�s�o�k'�z�i6r힀f�eh���)ʴ/��/:���z�P�*ܸ�7���gD]�	^T%>���y�X�77����j��,��j��J��0�Sԩ|�WPp��}�m�g�{��Ls$#�J�h�VL�C��b���9x�ǶQ�1uM�U`�&��3������#(tt���9)�Op�΍Ᵽ3Pp-�ϧgZ�1�rh@�;� =�,Y$w����x�.]��W4���{ᎉv��/�P��xN5�՟G��2��|�{:�V�q��;ztg��2��A���e�9e��x�Վ��	t;@*,Q7D�T4�ocof��U�wF�s�ɾ�r�l���ؐ�fի�^�)��V��AeE�>ί�M㯯:̾�1����< ĥ��V����oV��\��3�\:��7#٫�Ι՘�W����Қ�xE��e.%����c���sD��g��=��c������ɼ�{2EB��=��R���z�]O$ħlj�W���#c;��d��V���s[�J}Է'���Ge�\�鸬�i~g8�W��u�|��:�1���������<.#���7L�^<,��1�	�\�zf�T�uM��6�
F�njx��;��jɼ��f���X�,swCt.v�����K�+�4K�"6�^Z)V�'#vF�=�=K�ި��U�4K�<<_��`��$h7�+�=�05�IBL�`��ti3�}G(��n��o13���^�TV���J���a�L�c��
pgL<�J���4�9Uh�[�����v+)�ܻ��kF,�=�贫�F�8���������j�2�ЄP\�ۺ�\Y����֚�i�����sƜ�넫8�T���w[�6�V��o=5�s'���ζ�OS;�P����B���aʭB�IT�%�/^۸󾽼�g�P1M�%�Tں-T�uˌfn��b�Q��oa�MN(~��˲2��3�Fe��@�3�[�_�R���g�V�M7.�����T�:w_d��0��q���Q��CDڱû���7���ϲ�R��w;�;ڔa�k�	��ַ$�6^u��������-&=�ܷ�=�=;�jRꢱ����e�z^�����y��G�ZY&�]q~�߃�\����L�b:t��7e����av�<�sٕ��
����p_S�c��K�ZO�8R�T/>�V9�7Pv�b�.�)>�]��u�(x��l�������3���{���\h`�J|P�N��+u��KOc�;�quv�P��Hb���%�;H�j�]��|������Y�Z�ʢl=�7m[Q|u_��kl8�Q�'ɊC���j"�NeH���(T��0Wn{bo6<o�����d5�o� �C \=��)۷+}7�KW��y9���u@�K��P�^������{޺~�X~�҃�L�:�����h��\�:q�31`�Lˣ|ޙ������T_��,��#כ���~�=s�e�]�K�v)�Y�<�^Ew�-p2�#B�'�<��^{����&�u/;5�x�㣮S~�L<%Y��Q�t�e�0��H�]#`�B�2��nUT5Q��Wp9Y���5��k	ķ�$l5C��R�F"3^�/�6j�����Yf�-��^����R��6 ������}g���g`s�����F�8�A��(cc���t�k|NX��)�G73�n�:��h.�ڑK�I�u=�sԷv��^VC�m�>G�q��x:���U��RU�1S�m͍���]���Ɖ�rC��]���y@Ǆ�5�_ji���e��O��L=�M�ľ�ۈ��'z���ٗ��q7�l�����@��={�CP{+��᷉3�Y��;ۉ�;���O��,������ނƮ����/��[��P�|�h�B����������b��m�6s�'oE�ڵ#'Cri��v#Lb���ƙPo�bU�Lv�xC�)g�s���m�3B�.��1]H�{���fӉ{}h3I�7!��������|3�LM\��e�c�
���e�vk�,*��V��V(0B��>��^�˧s�<p�9�����9�8���J��sy���p�˛�a�f��
��C��)�&bU��5��'�խ��k;��w��y��r��o�{8�( a�`�T�6
���ª��H��.�)�%�n�ݶ6G/{\�>�"<�/�~����xNLN5ő�;��Oy5��"Ŕ�E`|�
�+1�Q�^fv�	Bɻ�Cʼ�j�o�v*���x�����xn4 4����y��ׄ��49�/s �F��[�{yK�MB��4�sL�壻�^1�������P>������͚��q�-�|/�S��4�a�Q�\K�v�e�hɫ���`g��Zz���tj�g��:��@����0ˊ�f71!*�������ʵ;{&#5b�{���	T=���ҩR��.'��F���;�v�.�N���J�/��9]޹�o�!���R�
\�9Y���f6������s�{B&��|4����N��Զ�T�fOHu��d�w �^�
��#��}�\n�M厷G��=���^Z&����ֽ�0�L	m��(eq��� ��
"�V3ީC]�;c���3�;,��]ϜU�[;E�;�T��"��T�=$�tٞ����]b��t{�*.�c�Q��|�Kʾoed�V�	W��/:�.�[A����'��֒Z`#��j3�TI��D�/go���;������L�*h��m2���W��$Xl��<�6|!���g�k�,z/���){뽋�F��cD�_�G�7�AF]���4d<��f�V!n�)8��)W �V�U��T�<���]yJ���LdPX�_\mR�7��4A��U��A�W�y�\ݥ�Dv���jwX����[U�y�K�)V#{\�kz�q��L)L;�}s� ��]��\"w6�#Z}�����]F-mLO�Ut�/�����+o�x�X8�Y��Ղ���9H�u����4�s�5Y2��L!_������]5[�V�U=6Y�6�ُG�ՙ�`mU��˶��Q̩��8Rq֧:�3r�+D.���c"y���Ա�,{M+�'ݨ�s�>3䖏i{<�u�o�+��@;��&$�\9}0�Nެ�q�u��3�\��'��*�D>p[X��qj՘]嬡�'Bw�a�i#x�<^�o'`�	Bs��ƻz��Aə�^�׷�����CĜI�>K�x�Mpf�\�b�,��t��~Y�����2Gv��5�wf`Eh��Z�{<��ꛙtu��4�8^���w��L�}]S�����eS�5��>��9���ڬ��Y%��jH����" _
�(�x�Ы�My�ۙ�e�4�mn/{�}&�exMv���(�@r��^L�>2�*3
F�R�du/�ҭ�����u8�����Mۧ���;��S���+���Q���X��*`�a�d�[�F�[���}��`�_��o���/|�?�5�\qA*�'D0��+����蒖)=v �0fyeW�ɞE���6���b��{O[�Z�g_X�,rc�E�\{��v�&<w�oOr��ZOj�t���!�Q!�������ڡ��˙���9c�Dw;;sB�Q�=�flTV�gYÛC���+{6���0D{I���ǳ��ې�*�S��3��s��u����yh��o.�	��̹~h��%XLƉ�2HSqv���.~[�2���Y�0֚ه���&\�wb�b��U�g��8j�1&}��?r�{��%�h�3fC��^̟'`F;ۊ݇%9�^&O�]'<i�n�J�8�U�L�%� ��=�y��m�hZo�2q��,`��W
�4سC6���`o�}��5Rd����P�ut՞��`�b��t^��{�p:��c��;����^X0:�XO�V2á��i���1����7�D�P-�9+C$�ˮ/��� \��"'���=�d��z�D}|}���.���K��x�qV�=��8���R%��αS���MuVOa��4u�|�t�SxQ~�^fTC�q���I�*=����s%K����x��^���ص�ZD䣡��R�MePNhH@h���.!���_�.�z��V1�3w��`��B�yQ��]�J<V݆�F���!�ϰ��cQ�u*E��8�d���߬QC�b�8���j�7dW<�m#�y
��$2���6�r\n_R(��ť�%L�dWq�W�yeѽ��SӁ��et�'U�[J�z-v���a>���`5Â�os�u����Y��U���T��$ғ��Z��A;�J�dM���v��4��Y�ޏOR�[<00�r6=lFd�O&��z�Ri]T<�b΋Cl*פ���C��W	�#����Z��i�]�gN<�f,3Lɇy��`��̌�"d5OL��\�.i��-�^  ����z�@�B��gZ�՟S˅�Wp�A��f���zYq��y3V�M��1�i׼�뎏\o�]����C
��J=��)�����b[��w3��</�u�Q�u�ر���H��uH0o)��^����F�z!�2�l�Բnn*��,
z�:Q;J��H�^��m�T�d�*����I�~:줆G|�[�ӻq�=�c^��x��wy�.&�e@1HCg�������vv�C�!קaFՎ�ܱ�F�`����km@}����z<��^����6��(v�Ϟ�呑�Z�=)�%�K�RU2}E����W�Y�� ��Wb4��&cw�-�l��t�>Qr�6*b]�V?Q=X��_�{4m���� ɻjnՎ�c6��ii3]W���UQ�˪*�9D(W��8�v��ЈQ��Μ:tT�
�v���Ŷ���.s�w+@i��P�se�o@F�j.�>
���4�)[��v^_< �uvw>E��SG ��n�Z���j0�5�sj8j��B�kA��M6;uw��t���Qw{X2�����l��b����[� ��*]ԟ&�X5����m�[muAiلǢ�Z��:j�͍5f�ʻE�Ʌ�6�V�]��;g{&��Ӭ��Hj`+�l�4v��sܵt����-b+��a%3�tWo(^���.�b�Ma�ێ���$5�����p��vZ\�S�zX�m�G-m�ʘ����ѭ\D��ib����}j�*$��t��1p�j�8=�(@]e�0��o���8�2���I��u�[�R�s8#e�Z^�&�V	&J�2d�5@���H�J���Anb�(ܮ0:WW 䭵cW�o(�������Q���D�k�]?zN���Om�Г�������b�h�6�ӳ��ء��������˾��h��k�zv�\�C"��o�m�r�jj*�t!b�G���w���H`�5�YaK����2��4��Q�,.�i^��y��m�|��Y��L��K�!眣�y�K����[���JU��Q2�Yl�e,V���wK/�2U�)�
��a-�5���67�n���痝W���xǧp�y�C=헛T���p���f��nv�1���Z���rb`�l�Q�۬���^�=x���hvV7O�� �����	2�`82^���ʖbh7N��KeÛ�f�R8����Υ|j�CNE@�BK2�J m�|U��2;ζs1"_6�p�7]U���$�Y�Gzf��yk[�H� 1�Lq�c]XE�gj�E
�[�ݳ�}���}��סp���ud�}����4�����!-��Y�����U�ʂ�ʃ���^��;�O^�3c��
��teud��æ똷����xROq�ZR#�چ^��D'ncyn�R+meϭ�CvW.�t�Һ\��.��ק	s��$�pI\^AYM^�V�$�������Qv���r��{p˽��/���'��炛����B���ކ�E]z�H�|��Dm��7E�v� ���^��w�!En۝�K�:3�'pQ���ܹ�Uf����ӫ���p��6���vv\c�v@��8v+��ɂ�I�d,�/�9��Y�^vg+b�!®�kBMU^�g`�ݬ�lrX�m�H�צ����m�ۛ���\���l*��*j �fތN*ܬ$��l5W�\g�S����v$�r��3v�d�J����w%!]y]]��*k�bi��P�@�2�t�E�h�n>��C4k�s�0mޘ�-o��w#Xras*q���s����l�h-u����t(���ǽ5�%!��ʼ�V�U�&wg,�(�{:_A!XO��]| �KHUfS��(a!f4.IEd�99.1NY-d�I����K��U9@�DY(VJeC���4�@ҙ�!��T9d�P��999!����INT�	IM��K��8M�5!�AE DS@U��9eA���Ffd4��%��JPБ�aK�44�NCC�R�NFT�D@�ӖA�a9A@R�VAFCFJ���Ya-FNT�D�fd�f`Q��QFfd�CC��dd�E4VIf�E��%EIE�A��YE9!��d.�C@Q�ffa�CF��2Q4�f-�&I�ѐ�儣FTRdd.Y��,CA2Y9-K�VE@UUDRQFY%�N@�V�~ϳ�����"�gF8M�n�L���CF�2�M��2�-O���Xx�o}�3ypp��I�f�7gqi��H���+/���6jQ���|N��5�k�y�vk�,,Eo��4`��Lͮ1xm�gHN=׈�6���<���N+�
}ke[�;jg���w«mO
T8��
���c	���vU�����V�Ւe�8_�}LN�>z+�S�P��g�z@c��ª���~�86������E�U�U������غ�pNyI��\<��w���;�.Oo��fVȻ�L7�V�f�JL�uQ�T;�_��L����{��γ��Iԏ�{�Y���5�v�7�K͊���}A�-)R��:��T��
�C>u�pC��A��@Y��{�C;�Y�{��&�O}�*�% ���B��(�:=զ�����x�� A�li]r�vN�n��Q�k��w,f��=d
[�t��N�����pu<�J�Av*xjf��~��}���S�<sv�r���]C~�L0|��ȸS#k[���H2w�9r�����W��6}��W�l𤯝B$�`��P��0���a���e�} Ev�+�D��X՛�䜕�阽�f<%Ġ�:�i��%K,����F���}�{Ә��;U�F��o�-�Y���X�.����*���K�ν��ή
���\t3�S��R]��K�b�
u�N��tsGd�`�K��Y�nݨ�X�wX�:��^��g6H��`w�%�e��5�.���Kr�Խ�J:�L���,q[��7��8��;GOC�X��A"�%���P����m\ZG�ΖJx�E�=oJ������ɭO]I�Fu��K���{�:�Ô|�S%q��-<۔��О�1^T=�r������-"7�����U=��q�?)���!|��9p�OP�*x�J�9�d�&�R=퓫��nf����Zp6=��*��m�y��C�4c���[K��m윌E��Rs0v8U��lg��R�n"��O;[8��l{v>���KD���w�ۻ˿[�1��͍~=`T[� Y�	1���9}0�:x�	ƙֳ�:lS���'}I��|���U�5��[V���:��4�F��A����a���Nt&�3i�;���;�g��ԧTF��W�h���3�U��.��TL�Jd{��a� gC��V�U���̭��DwK�����z�#�'�
ޭ��E���_	��IW�h�o3��n̉��h�������˙���c:p֪�f�VN%,T�iv2��t��
�^�� � ���=�l\�L�X	�١C�Z�L�i�-���Qt8�N�&Ջ�΀݆�#��t`f��n�n�;1�8���[P�F�u��9k�䳥v_q���,�y'<��$C3<���~g{ B�4/M�ٕ+t:1�[�/3V��}�r�:��Ѡ�Cؼ�O.���}/��D�$��~/��Z�����9�}�£}�hAkU�CL�Y�<�"�}%Y��	�>�O"�>�nf^vb���Nf��o�#�!�kE&��,k������f���Q#A�%a	.�u���\��oR}6���:=�=e�-�K�e��<˪�������qj��w�h��3B�Ww�k.��-4k�]b���Jg6�"��t�bҙY��u��\�`r�_f�������9�~�ۺ�^,�Y�y�h�^m��~4�*��	H]�e<��/Xu=�3P�9\�ɖ�`P��9i���5S-<&�)x�*V�A����Ra��U��>��/�˸b�s&5K
e����+o��1�.�������.��5Ml��t�	�����NA������:���z�.����Ǫ��|.,l��2�.���������K��|�)=4^�x���2����m�X��Ҏ�3���ܻ;ft)���;S��Ү̅�0Н.��������bkNB�s�����u�����b�	Փ%trš(��ή����t�H|Y�R1��.x>�oW�jV:�/l�As�N.��n�`fqG&f�z��ٕ��>�!����h(x�!��3v�h���n1S����%�s�U���A��Ō|)�kn���5��	q�!��v7º�)���S����S�i��Nvo`)�Q���7��3�}tt���ط)4l����F;�湸:q��?.鏥�1;I��;ӣ�p�a��N�{����	̩�6��\��moWlÞxi�(."��ֆ̫�vm`�3����*y2�s�����O��.��n����HĬT�/ª����R�gZ�ԟ�w5.�(K\��/�;��Rw�i��"+#꤆o�].Z<�7��X88hY��a�|6ǡ��i��5�ѵ3W,�Jj��Q�q�)�>
v�ݑ�b6,h[�j���2��9>���W%�eZ�ڎ-+��T�:���qKg����URfH�[Sr�E�.���+o�gG�J�����7[�
� \T@�۲2/DZ�����2�Ǟ��u6�����u����zn��z���'dİaԄ��O��>�:��3o �a++O:��÷wծX�ãǜ��}�r`m�;q�9��w6�ɵ�z9�5�J�'ݷ��qkz�?m]�)�a[s��Y��'M��DKB��:��~�9����Գ�]��<+U;4(^m�5e(u�^�/�9|��r�.KXt���YҸ:�O^�o��˩a�4�S�62�?S�p{�J��6��f�b����n�fѽ[(�^\���M���{k׷֬�?,P�+���c�f�r�M �&H�TjVV�|���ܺ�z�
�77�c���y�v|b�j�[hXN�!�,VK`�6��֕8�"q��Ż�iGS��[�7��n�Ƈ:ާr��b��`Fi��«mO
UZ)��P��5���{�o���I@��~�@b�c�S��^:S( 芄�Z��bߗ�z��̛�v�==Ј�A����if����sP���������G���J��F���������MaozR��R*��nO�PVU�F���徵t8W.��Nt~�Yg(xs0m�k��<%�}7;�����D�]�6"���A3-3-iN�w���2}��M9�\ƶ�n^�N��V��+tV�\��ZN=�Fmv,�M�H���V}}l��zd� �D�x`TnX����z���j�x��e��A��-=sS;��[�ǳ��Cf�e�|p���ְ˺M��Vm�|�j��3�t�n�(��G�.�|�w&K��{�Έ,�-���B���*�*P`f	��"��3.e�=Z.7��9�HĽ8��N����B�)�gF��O�cL;�	���)}�GAt��IV��\0��wG8�.޾�ud᜗u�1����n��CqV:���L0U���iH���VPL��:s9n�1[C`��	�WU�k𤯝B$�`�yp���fz邫.��Q�M���n�*������(z�/���B�ޗI^�,+����%�(�y�GΦ�Yz�߷���i>��}Vl;����W��tg�jܝ���y�&�[ G.W�r���)��}Ej��2^�P֟���}Ba��b�Q+��Qq�^&6�Gc�}G%+>�M�/ם'V.ظ� �l����yq�8�h�j�k=Wʆ*&)�lߍ�
d��Y/g"������3�8]zG�LWZ3��-�!��̗��<zl�@&<s=l��f�����s)W�׃�.1]qՊ��2zS�'&z}r���"*�I�B�-m/w�}����l��^fi��M�Լ�Ofw<
��{���}�ii���ʍ�G��U��v^J�EB���죹����Ł�˨r�ޚ[�Ra@D�g�p0.ɽoC���ѐ� Vܛ�l��|{���B�9�-��+Eu�Z��0=m�0�G����/��w�z�����u�9����3�`�6����9(f�����]<��f�5T����,;�F�ƃ�ю�v�v��Q��&8��;M������ٸA��D�4��~�Ox]KL��3`d�j_ :ݥ�cJ����=���o����,��s�;�A�bv]�w@���I�S�Tu�<<D0ߝ7L�I�m�_�{�g;{Oݬi�6.�Iȇ���*�!�7�`s�I��!r�4(�=��f�����۬��p�Х���%bqK[}��C��/�'���K����X�
n�9��[V��������D/%?���y��狼:�5uL�9d�7:&m��gmn��7U����#����I��,k����i�a7jN���6�A����v�8�[��,Zm����'�WQ�.����R\)|ˇ�y���h[������.?^+�x��<&�7 ?fE0�:.�#æ]b����R���.��~Bڱ��>5T�Y}�D��=uJ�]�$=��w��j�i���3�c ����tS�"IkzV-���I���}|G�:�
X����YԴk��!Pٓ�o
�Q�5\���]7�6�<$��ĵ��D;��'�}��7���0<�:K%�˵ȣZ�E��^�6��ٓ����3�({:c����C�碬��7�]s��ng2��K �1Q�zXȃ�a��9m/d�g�C�L��[\���2���zp��^I�97���E)~*�Y۵ �N�Qq�p��s&70�KT��������mB744]��xa�
T'=V�t1j�\�OW�D��r����_ú_E��q�,Ｑc����k�ǧN�,z��I�F)ޕ����H���R%�����L�Yꣾ}��l+�<��)�u�׷�Ƈ��C�h���l>��u�f��2.��|%�, ^�J|PȉƦ��(6�$a�ƸK�w�D3U/i��NY��;7<^�>����f+mVl���}ܪ���F���Y�:|F��сn�]3y9kj���t+�ϒ!�ּڜ������	m�u�y=�@�7PY�/JGzcZ��:ڂ�ԩ@�./}Aq������;6��u��D�u�8򙘰|�X��C2�W��!�q�rW��k��U�ϳ��>&��fU���V�!�.@�/NN)��w��,�Q`U;.����<�����s�YX֩<f_#�X�g_�y���z�ޕ�w�3��&6`����S�Q��q5�/��_V�wt���s�-p:�vN�� G�BG1�ޜ�������ZJ./@���z�.��԰��Z�Ք��x5.WBm�o����Ӽˁ��XV(l�I�k��u��S��Ѕ���uU[�ǃ��9W�z�4ԑo��L�H2�n��1�X���#ڥ��0�{n�Ԣ޸��@�\���g���1Sq�[��`�pS��N�f�8R�è�U�r�hŷP�dK�;�S����QΜ�[hX�v	��������^,��<N��ח"�30C'm������+V��Z~��2�@���n*_S�~�XϨL�^�<�r\�d\�E�K�}�ZF�^ff��V�_1�1���p��c�#��չ���M�f��ح�1�g\�꾧�W����Z��	3����3����%��#¡k�n�&6����g���l�g��|]�S�[x�Q�D+�dwV�P��spi�ܯڳ�[hXN���*�l9�Aʻwde���y���e�t�� �}keiv�싛�De3�U��(qԢ�_'Quxf��r�t�Y�8)�sfW;⺥�;����k�,G��2���6dÍX����mcu�e<S9X�-x�Uʖ��{4ˎ�5r�ۼYU���ڽ��� �r��;D�2YI��`5��9I ̊�y*[�C�bs��ӥ �:�t+�Vl��h�<R�ﮓ�`'\���ҙA�[z��6��֯Ԝ�^Ǵqs��NB�_��>��qT�O����7����'<�W�-{U��p82�r���ە�`��P.�gŞkE&e�ݗ�T;�Zu�+!���/�?\�[���C:T��Υ��/�%�m��k�,̫,p���G�ʗ:���E��gy��ʥ�*�����K2�eT�G�ɖ������"�-J��ط�+������у���|���� �Mi��VϡM3:3�����1���d��S�X��j��j���Z����n�O27�Y�^��KU��_�νy�ՂAV:��L�`�*3r,!d�y�ci��Q���AB�=U���u����b�o�1�(��t�n�h�5�}�|�j��y⺥���h
ax1�p� �80,to;�����m���)�I")>��JQ��>�;�u�;\���l>����JU��^��ڸ��a��<J�IS' �e�)-����M�Eغp�Hp�a�n�X�agm��AW����Ess��e��0@m��.)�r��,����.��e��y��Rk޾��Ff���Y�ءD���ti���Z��tC{�2x���/���'��B3�n��\�Ԋ.�u�7]�*��+m+j�I+W��4�Uȸ3UNab�������땚gG}ۆ'}ı�&���U���R=�R�9��r��n����b�� 4���+;�<��s\9�5�%8�V���gL�ͷd�:��+u�P��23i�yd{�Ke-�@goU�Fq�fjA����9�2QiN�f�CZ��fes6A�Syͨ�)�\n͹
��t��
6u*�]xwx�:Pb�s 7��q�x)R�����8$�_�6�wgiE<�-�Fn�Y�J��]u�͔�� �B�!��� :��7�G�m,�љ���K����z���Ev��Š��i�xg(D�E��$c���mu�<M0��^��Œ�S\���e�#��3w"���#��I{:5Q%��x�q[�&�b,^R��-�zj܍깧z�4�$�[�5mv�f�<����O�-5l,�*_c�n�y�zD� ��lc�] h����I�f�
aj*Iqw���q��X��t����:�*�M1��P)s�J�.���o���8C)*[0��vP�ѻt H�����ۇ��q{V�c�7�≠;�-��0�]��4g@�V;���jܠ#�p�wT�tಸk�5�O*]�F�q�m4�u��������I�4��#2H��B �bۢ.����:�ޭxu�=;��r\;���_,=����L4��w(TOz�&�][��}b��K+��ԗ/3��*���ѡ��+W횣8i��S�FәY�TR<�F#�Y����з�Y��Iw)��`
����ʹ�h �H��9p3���-�.�WG�����8�u�V�MȞ�8��l~�Np�:$m��KLm�M���֑	�2fp SJ����Y��p���r۽C�(�B#S��n���uR�(�/K�9�<�7t7.�:{˅Zud]۫�y�[�^]�ş�tps��M�n�	r���U�{s7g�8ɺ�Y���ූ�2mKs6�}�tc���Py�֮�%�w�������`��R��ˣu�5c�4JCuh��GlR�)V�2���z�)������l��EN�L��{u���B��Zգ��0P��/u�a��u}&�9��bz������{l�1X���Wg&sxW<�:�;�]��r�ø4S�aN�d��� ��[C�̮Ք,�l6y8�Dp��ZX�%�<�9��Ѝ^��������>�T�3y&�m��Շ&�W��w,�^%���Q�}*ږ���/�E+���K���D�|�+u��.�jg�_a����/�~�R`C�'�2As����M�����$=*��^�Vfs�����;����j�L�,���r ���� hrɠ(�$Ȋ��*�!+&�r�,��
�Ɉ��ri�
(�"��i3,ʪ��" &h�rF%(i)����S!0��,��JL������*h�(hJ,�0̚���"2rbJ�2rbbJbL������� p�$�3"��"�����h�����(�"���*�������0�i�#%��2*������
j$�0�*X��+$2(���j���rJ"J)� ����*3 �r%��
�(j��� ����L'
�3hL�JZ�+,(�i"
*� 2j���������*��L�J2 �
�Jh()l�"� �b
P��rJJ��J�3
�'!r�0���X�)r(p�2��
����f*i�L��\�����Jhh2��*h

Jr&�����hi�X���@Pe��ZZM����)H:��.�]ڧV0��=Uw�	�.���m�Z�p��8�pJ4�=���׶����ZfN��R9�fN���ꤎ��_9\o����]b�����XF �5dz���͹NuvP�o�t�ojm'g��/FAǗ���h�v��1jAUz*X���*!�[�W{���Y��!��\a��Z3� '(_�V�e*#2u��#�M�l��@�l�tި�Gn돒�SA��1.#��+����O���.\?b�_�P��ƞVu��y����^��s�`|g������yql�u�9	��Y8�:�Ҋ��?]�oۻG}��4x���',ŉ���4\���F�:�:%�����!�[E�s�H����7��+ �U��-l$N�In'�U��JL�(,t���ǈ)8`�4�B�{�r�<H�3�·��b;��ˡ��5�6<�*�TxΊ�F�kuA�޵].M�ۗ��,j�z��l;t̞���W+���Y`:�D �pͩ�äuiD7Ll��D����B���G*c����ud�L�^D<,a�E�`<�F����vA�zZ(��cW�/@U�
]�3{��^��� c)1t}�Qs|��ő��o=c�:�c�5+��<�]D(��]��V�g�n��S��3uy^�8���o`V�.��7��P��q���%[\T�_ic�j��n=�g�跨�c ����6�P��\��`�w�c0�<��0����w�WkĒ<������.5ox���z��d�����ϖ�D����s�Fl˞��LU(+
��K���}��e�8A��mc�T��Q�-yh��\)2��>y�R��jT4����|]��ǹ�Y�H� '��J'.L��u�Lb�+�L�໇�!m.$:�.���m��h�+�uh�޷E�h��̭�<��c:b�<������$�d�a���
��Z��|1Q�Ǻ�4��I��l�(p�u�X_^Ft8�����L��{[������M\��BY�]Nۮ����S6Z�;�|V���ۄMԧ'l����� �cfv��2}]Z&˸��nA�eh`ˮ��Y�	;[3�Q#��q4��=/��"����qe��Bь�.x�h*z��S���*�\"\>�2�u�E{�Ϲ?��	�5�}����)�x��"�R���n�������
��ӳ�-���
�jd��-�C��SUD�m谳@�U��TQ6	vD��2�p����TK�i���vr�� J���mŨݚ���
��k?G��e���)g��qeX�7��t;�,����t�Uc�u:�cs;�R�-��s���3z�hw=�����6cVU)�}i�h`�|P���5��^L�/�¸	q�H�^��/7�ynS=ݗ�#����˫�:���g���;�rP�^�L��]=��ŹI�u�cx���[YOٺ��3xџ ��ki
R���mwJ�ޝ<�v:����q��͡Fm"����
R��{���3{(䚉C�x
	�Wƃ#g�>]C�k]a���j�yg���YY=����9��kK�<�a���Ô�IE��T=c�	uu�a��M�O�8��T%��鋣��]b�V���	U�)�Jt�}&�g��:<����CBː��M�!.7�s�2�mU�|������OQࡇlK�":�lh;k �ڥ��a��%f<���R3W�נ����b��s`��P}�]�o���	�k�P�M�,ͩ�e����|Qn';��O�>ն���`��9�
�s�l��zx�6�:����]wP���ts9�6�CٵV�^K�g�km@u�#:
y���d\���"z��C
�,��}U`w!�=K2�ʳ[ԟMMM�䨲���M��#�G��R34����!Kr,��}JG����Œ�6>Q�ٿ`��#�j�h���x�\K]�S1�5ؘ|(���%�w�@"'�I�׏9�޲������Ew���h���c����R�Q�cҲ>v���d�nA�x���o>F60�Ic�-��	�;dL8�w�)�l�@yէfWZ��`_U&G��k���9�E��Tk⮐��]�������q#s��-�8յե�v�'�C=6vr�n`)�}0�Gf<���0L^7��r��t�\�B�J�`�;�
}ke[�;T[ܢ.3L�[Je��1�7rv�Fd-]�BЄ8y+;-��,�:����}4W��&P@��ll��}�|e�kq��Ԗ�G�Nq�/���������:�M�>6NyI�¸x@]�sNv$7���/�]�Q:E�3�z�2�����C�yb��ϸ��w<
�M)�wg-��^m�<˾��P�v�u"(L��oW%��]\b	�i��\G��v�q֎{���3;S��t��j�K�UL�tw����S��`B\�C�ԫ�]�|(Wpḭ#z��u�E� zm�+J��V\�D�gg�U���)�gF��l�[���+�O	�T����"H���x�b�+FЎ$~��������v] ����V�	��9�;�6�q�$
�pJ: �<���Z_C3za�;�eE[즉�o8��h�c��:���X],)ٲ<Y�wݬ��΍�`�-C]Z�usMˏom�����+�$)uB����s�V��~�01{�����DEv�`�U��P�n��YDL�����Z�훏�p����Ԧxm�u�V�uIy�H�[�»©��:�GH�W/u�)	!�}���9�>��bD缀�P��kG�I��`[����W��,+���ѝƷ����<�B�� д=�����6� \;T�}.*�U�C���|0L�`ө8��e��6������'Mh&w���lJ�P֟���g�&7��V�ඬ��U��&��e�����=7�y����;������}�L���Xw�׃l��kxYy�=��*�r;�8��}CH�[��|Fr��z��}]s�NJ�lFҢ3%���zl�T�,6Ae�n���4ju�S
d�LWL8�8�Ɋ����D󵳁�anX����x	|`�dr�됿Sٽ~}�B5�b7��)�zY7�sˋecN'Jr9O� L(��q��釳��P�FJ~tx���7KSZ=������d��@,v*�6�+�uI��5J���*����qb\�����<f�u:�]�5�|$����=��/dK���V��cKn�H��f�K�C@��ٕ
��
8���;�	�X���T~��s\^f�Ywٍ�X��X�I�c�Wsܭ�ht���h�ؖT�o7���8P�(xM57�z�3)t%�p6�j~���R�*&�S�w@�ˡ�u�u�fs�k#��,����_,Ӣ"[V'e��N��e���ڦ
9*���V�D���1�9��Y׵(?S��������9]�e��,��Y2a�j��%�F#���g���wWsÆ�~���7㢣�S�ؔ�[�F�ڸΜ�L�^<,]�[;��S�W�Wzzot�eX�J}T��VghCp�ƺv�f{՞���b��7L�@�������'�毞���S�V�Z멙��Di.���N���ōqx�U�5�>��WTNѻ�A�W��|�Gy��#����6�Od��a✺�`�Jɸ�:�T�a��@�ʫҘX���ŧ�/hK��P�ũӊ@�:5p�5Fa��n)��l`����@Oc��z���6pO��k���MfV̘�`Ec:b�糦�z���\'�K����e���:��j��b�P{:��������l�Ϫ:nuq�wSE	+ғ�o���5�K[���HZ� %h�7���:=�oT�˞���K��I�y��VV�1S:og �Т�QE4�
�Yz��!�ȝwM[�T�-���F!A;,���5�p�	�y"����5CԪ�؁����gm�im��a1Lj����;v���
/�wI��MD���i�o�A^�}���MA���I0N��z����b�����v6�������Z���kG���F�,�{�H�G||��y�t��ov;~�,��^$r�N�����c�T�_>��v{:TM7^�R�#����J�!o��SC�q���#);�Ug���}��o�x�|�����e��'؈۸��O����km��*Č7��\	<CA�RJ�uc^���͎֨���[}3x����<\l�9K�(oy��-[��Vҭ(mL݃����T�+K$ǰ.���w�&z����:�y��,���8��"d��L�0#�i���_���"M5�A2*��dl�L��a�i�S�g.�6e_��"��y�N�}�X������sE����ċKjW��܊���a��>�G4�rҔ���^�y�����LuJ��P��\$͢k>�ĵ壜��v��=,9'��`&��V��z��W;O�|g�W]�[�Ɛ�@y�8�::.H�3B�Be�4A�7/���5le/l$�t*����)uV�"yv$:�E�"���7Do;��Y�sv�ѓ��nKʻ}6�%1�7B�J:IA�:oҁ�;�׽�l���E�t,�ߚ9��V�,8*�(a�UDC�:�l^�]���]Q����@Y�y-v�TƄ�5�}�R"��1S~�)̓l(	�-�΀�6(0�T���zvIE�S��Ŵ��D���lm�_��s�2_���i��$����7=��ŝ],�7= ��ʔ2[�r�̪�M�&`�R.rr��f���f��ְ�ނ¿9�Kv�ը�n+���]D$8@���P��k��Yp{�S�����F5�7⮺�A7��<]X�ܸ��/W=�b�//��p�3����g�A]n���]Ƭ{��R]^��3�{u�j���C��|8�6H܆��cT�k��܋��U,�0ia`z*�RЯw���YX+<��s2�阶�1:���.�0��b�=.�3�p�՗�Qۗ�B�;�bwt؏����2!֢W��5�~&.uC��Y8W���,1�dWWnҽ��a�8;�0{��䤸>1%�Ѥ+Z]���=fԅ=��Bs�s�[TL�0��ϟ�
8��iTe��v�}�N�.�ra�j��`�:�cÖy{��ݠP�E��V��K��*[�K���Z��M�8j���8��8����r&2P���)vS�IF�=K��^�EO��sAӼ��\�ċ4,'v7�K�4�H���K��{ٞvw�0�'n+%�E�JE�)��j�m]�b*���S��� #�-G�a�cs�'{����[N5����xs7:�6����x'\b	���jz��6���3lV�JvJ���Lg��a�'qY�.Įk��ߍ�WZ`�BX�a+��J���w�S2U]H���[b�#7���3ҷQr��p�y��Zpz\���O(��=d
U�GA���G[��o�>��pM̩��^u��Þ�n�u�Ȯެ�U�sj{��9Ə��9�7�a��k���j�C�&w�Fxk���Z��%^zR%�/
���P�9G�
��	r��b��o7��H��h�y[D�Hŏ���h�%��ŮH;��f�;��&�ռ��S��.፣�,xI�3 �
re�t6n�l6�M@e�K�����C���ڪ����n�_;���*b�m��c�&nƮڬ����ؕ�CZk��+jP(mώ��8g��|/v�����N�(:o3�@�~�ѐ}�.7g�b���LL�j��W!x��f��^4��[V��O������[���@EC���j�DR:W�*ÑܺS��3kV]v�;bg��E@W#�{�=�u�ӝ�k��ݾ1��ͬ��ӟYW���'^Q���*�uč�&	�!��B0�&�9{�/D�{:ݮ9��QoN�'_P{��Q�wY�j�P�*/�F�ٝ����-[�����o��(�S�r�ǡu*L��Kx��\0��5t�WPp��b����g�oV�/qn�F]K��6�q�X�u�p�78b��>�HItꄛ���^���)�Iȵy��r��7�t��[���4δ$Xs��MY:Nٔ�1������/q!�|���Ь�WE5�շ��\�,�-�od,(Nt&�3jv*Դ!��.�K�?"�tk��
��y)�f`����ve�Z#+��<,"�f� ]/MP��P�8V�D�k�ϚXb�����\�r�W�W(���bS��G���#`�v�Ny��&VL�-� GGLocr	�\��x�MB@ü�4�t������e;cV����a�q�9�t�������8��ZsY�J��;}�����$��X�du+3�����z�mi<�襌�b�����:��!O_u����J�du�1u��}%������c�ōuQx�U�5�>���[���h�w�ݍ� �kh��
R���/H-����a�O�������Z�67�l�������Rb�G���*�j4&>��V���V��X���h��
�+ }u,Y�i����W*�����1�p�j���.Z�CGrn�1`��)䜟/�9F��f:��oӨ]�fL$�ewuCF�$�\�.��� &���o`LoϗwD6���kҷ�0�Vi|��3`�L��'���ۉ�z��hN5��|��BP�hK��o:�
-���� �a���Ŝ4�l�a�}���2�e���B/��76�xH�#�æ�@�8�B��|2LE(���o%�[�w�zf�ckD�M��<��VU�o� [�����R�)wC]۹�Z[ z��#rýL��XR��F|&��s'( ��:�(�7B��o"��54tޮz�`�� k�����lZM�]FN��B��5�n�jDҟ��v�f�!��5�p���A)��m�����ո%�Dݜ=��
��fNUy��]£�ݶ��LP��2���gv���Ê���V����l��0 ޗ5`L(Mkf�`֊5�#͔z��J��˔:ڤƞ�ʘ��4���vy�B�q��J��V�/�'Kb~�2m.���ɖ��q޺1
ޠ�q�1Aշ4��T]�x��Ք1�C���#W*����_t�JG;KM����3#xpub6��'�[8��sP�"s[1,�G{r��U��P�A�Xm���wt
�{��;�+ �]sE��Y����/�m�
�u+�f�ǚGb�đ�kMm��Pilk�����qЬ]׼6�h��Ү��Rw��)]���a�]��6�xrv�������
��e8�m��,3���R�����r�Gx\X �s:����*һ�tr���㩕��q�����yV�b%d�\�GԨ1c�K;p^��([���.��P��������n}p�Df�]|�̳u�m��_teJ�41Iv��s\z!,q0�8*�� �ݗ�㹖;)Eʬ�z��ʰ�ʄ��v9�o��ej皭m�@R[�ʹ\7���5
U��7l�I�o�au�w5������j4��e�����5V��*�U�&�Uɹ7�rK����1�ل	͘v�+-e�:�������R;�C�nub��]A棢qj���$>���f�W.Y�lF��R�t�]o%�*��p:����j�m�_S|aw�|�$8� ���V.��rA{(�gzr4ؗ�N�)u��u]#��4-|]�Փ4u���gH�S��Z��60�Eʹ%�v� ��1nl��4��b�{��J��>Efl��5��g.Lnٚ�`���?�&���]��.���v��H�6zVr�gN@�]�@�xL�D���5��%��T�]u����u�����v�]��k�5���km��_:����}v��L�QT҅4�6`�e@PQCE�(��M	K�AALH�d�	@�BP�䉅T9&HC�S�C�eTPR�����4D9YdY�eE%�FL�Vf$@e�fH��E%5DEK1TDђ9	ILH�U4-,CAA��E	�BTYdĶX@�R�R��TUSM%�(EQ4f#Tҙd4�M5D�ESTR�T��@H��eB�T� P4	HRU1R��EM4�J4���4�f-UHR9&MLQE%�#HRRPR4�(R�B��{�]��t6��Urm�)R�r��z�L�:�/,����WA��5$�1A۽�L�|�[�;�;Ն��s9`of��=�Z�4�"���P'@F����S�+�"D�oQ�.�yh�>o�@��Xkϙ���tq�2�ק-@=�tU���o�Cm�L����&_�Ʋ����]Jg6<����vFV�]�ל��c7��U0ʳl�〼��u}�̭��@F�:b�糦�\��íC��Sٷ�z�������6�S�YS��Yi��}����-��-�X1�E����w�U��n�X�Py��ÞB�IIxg�����Lo�%Y�]O�n
�������=��y%r�K,���_!�{,�(��2���*�7�M9���.2�@�l���t�d�g�87�G7�WS�C���s���N̤m�O�=��S���)5�P$��s�jəy��\��u��9��[�!���)�x����{J�Î�w����=���c�87��3K&t�8����rq���G�ϕbF\k���������'B8K���1N�f�Sr5��<\ln��������S�l�t���|�R�L��ǒ�F��-���&��eѳ�N�z�VEwWH_�>\�z4��h���+Yx����R�㋹�7���Ct�H�]M�Rvҧ�G���1�<��y6������`w��t��6v���f���g���b]*L�.^m�<�b\6q�Rb��/|��SV���wa�ֈ'Iw a�-��q/Er9����>��lκ�\K�eC�x
	�__\�g�::�vj�k�e�cƐj�w㣆�߹ntY�X�Y�+o�&��u��S���)�����
_���K �=�����^�3���l��	�vF�-p2�#B���RB�iX�\]�C�2y������������-3�X�Q���=��[Zs�_#ࡇl	wbRdTf�]�o4��l����S�۹�:tbG��oG���c�/ܾ����s`���_��[ �6���L����S}wU�;�&`�e�u(vm`�̿{}�gڶ�͔)/st���6Z���}R�3�c�"���6�����jǦ�:��+�U3�ߕ<z=Vj�c�sՔ5NgЭe16G��0â<�/���(v�,�6�8y`���9����h~ _cM{��k8�Ҏn��/��F㦄x�t�;ɏ�έ>f�Z���	����[�,yܙILÔ[E<��ٖPpq�2�kZ��T$;L��ql3g[�0f�"�Km�J���^�bqu*��7��<ud�=�֪V���h����>���g��^���!MV@i7��#!���s.���U}:Q5�)����r䒘u9ݽ�2�q��v��Y���g��A�+�>�f'.�h���
�o�c��Ȼ�T�X�R�����z�^k�̝��<�4S���:���� �ԭ�c"y�`MS����ᡄ'�����s��L+�Tv
���J�"�
u���<����?�:��rެ�k��Һ�i�R�W����z���a���t�K��Ė�F��'��[��.�}����B�p�I�~�"�$�Vrgv^�4A}�q�2iɗRX�9��3@�vZC��OT���߫ǭ�gC�nq [��"ϑ�ʷ'`0�m�":����ɥ��u� ��=N��K#�Gg^���׺�:e�]�����a�\��[G�<�d�<��p��`EG3\��OWM�G�,㬉9�
�~)��L�q�vLO+�vz^*i��J����%y����@�27]ld?�R����=KU�����^CP��Ζ�ޗǎ��S��H*��9�v�iL:�ER��ֲ��W̛0eyZ.��d-�3�_�2WK^:���JEsP����.�*t[^v��x��S��R(�y�hA�1{Ek	��rB�t4a�X5{P���C�Ԁ�P�:U��r�E�+t?ml���	�?h&lY��Kn�wV	�vf�\��lW)K���N%S4��/�(�f�h���s�o.&�
ɤ���C(��u���d���z�z���tk�}��'ҵPPCL���	Ӂg���y�L���nQ��0"��v�X�3hx)���(��Ϸ�a~���>��Yk���*�1�̡M�1u[Qe=��M�a�/�:4M�"�+`�ͭ�·M��1e=5�a@;;.�`ű���S�8���[>铓�mX�i��O9E�bh�1�.7g!:�ŭY��1z���J/K�W�`�U���ٸ�yv��TX���T��G��ұ����ú���]�:�Ԋ����\���P~�=.��L�%�	��W��]A�||eRb�M�r%��3k#R��8���_M�Y�Ǵ�,8
U78b��4�	���
�� #�BJ�s�*/���ga�:���ܚ�5d�L�XdZw�݄ե�v/WU���4\�_�i&ڍ��S<fo�V����Pod<�A����g��̤!Թ.��Oԫ�^�\��WsHQ��:�I"�l��Fc�_ �}�ϟ�</���tu��4�8��x�{1U& 84�L�S�I�ț�q��)���PP��>�u�]�X`�9pLt��R����]���h+�/z�4�YkGHWN����Y�NjoL�6J	�Z�Z{gF�euK�,�Z�Xyw��.���5!�/�VA]�.f�5�klwNV�u<�QQ��T��N�HN�X�<=o9����K�9~�3C�_{梂N���&�D��x�:,���5{�������n�{ݴ�[��u��(���sk_f�9yG���l��(�irX*�J��Ca�r�Ѩ37�?KRu'�8j'j���N������H�FC7��z��J>���|��Z��I��6��Nv��s���p�jf��x��meq�ř���H�t9SW�g�&��&
�Y7N�m�]�#9v����3N�DQѽ:"��pq�	�|�� o��@�D�2�&5�X���<CS\V���k&�w6�<��Tu�v�Z}�-C�a[�lq�d�3��^�d���𣑼�=��w��ܤ�ʠsd����y��_���݆|1e�<3�l^��~��L��yht裪����F�v��{�1�G�ZЃ���="b�xg�ؼ�것���[�x��jz���t����/@�Oz���Y�[�L�
q`�b债�~�r~"Z��P^��ag}X��d)g+�0e�8g� 2b)�G��K���\���U�5��c��������e�a��{�q�-|Z	�L�">bl{x ��m���@��w i�y���;������D��/:5�N�(�<@{���uƅ�M�U�����H�YngB94�Y�؞�j{��&+�9�}�]�6t���YjxS�*��F���m�ٌv6+IIH���d�"�>0����	��J�!��hxƆ����5@����H�{0wq-�������SiL�*a��@w���>(d>�VGP­#!�N�vJ�;=��*���8�*�C�
w�^:�nl�0ؘ��-�r��!�L�\+����[gs�ޜsݴx�,�0)I�e3��C�����T����ښ���o��d��<<B���#�眖u���}޿	޺�r�Fʇ��ȡ|h;lʺ:�̬O����M5�$u��G�[�����rϦT�e����$�C��J�J��(T=~�K���ya�(��һ4:d�*s6�*��K�3B���jxXnz�!�4�\]�<���&�=;��ބ_��A9�|�q+�|p]w�="||<1��+�r�(p��n0��q���>������7���s��"�T������'�
�8��;k�}���i���yk�sr����eq�i,��Uj|�L��4�$�/��[�y.������ j4�5���uf�Z���L��n�������wqY\/8��NS`Ԃj�0�u+.��8m�������3�;���	��>�f����ӻl���	�>1�H�[<��#�ţ��K+�SEj~��7�:������{]��1�eȦ�>㯌���N偁��&�30Cޠg`!�kb.P�ua�*�Pk�r<��}��	DU^_�޿s����&x]�^�[��E٧�s�j�����#��'��^]���i���[�.���qd�1��؍8��0c&Ow)�e�V��}jϰ,"�&F-�t�ߧ���[�ݐN�&���m՚O#�t���$ny����յհ]h���\�3P�S�鑼�Xy���gص�(4��=[��Φb��f'R�;��q���쭏l.�f�7u]�S�gX��co�3:����-w�*E���j%~\�X�x:����z�r�'=�$1d�3̈́�}�>����^�Ș"ԡ��UW�uDu�T��tO��ENM�J�ɪ4�^Q�i]����؃�Z��q�=;���E�"Ŕ�E�������*�kE�&����.���}kj�u�OP~��~~�η4Twbv.���3¾/e��=���@��ȫ�*Ѹ/=�ʡ���ܠ�o�X�U��z>��Tg�Q�7#�e���e,�-(�Z.��.�X��c-����j7&�3C�7;�CP�ls��?�v��u�@(t����m%�a-fK�'or��\�I��I!���.ZG):��h��{��v��_�zgby,IΔ��|����Czf9
�'g�r-NaOU�8�3�a:��U{�~�r��
]�5[\��7
�O6&�����^Ӫ���ڵ��R�C+z�Զ�
��Vj�y�L��V��jT�����νzv�@���R����Z��u�pXۿR+�ͮ鎿\��mu]6���ѽ�j�ɸq���lcwO�㣍Jӆ"��]⸂]�R�_%=�6�y��^-=�r��\ڋN��^l�_<�g�kҸ�\���%u9�'ew5J,�,.#2����T�Zeh>�^zv�5�4v\=�ǝ;&ݸv>9~��U��sFmA�s<���&��en�=�V��p����ܬ�]�7�0�-/]O6r§�'i��������y��fǣ����3F�M��wI�C�M���m�c��=��y[�>�j,�b��_���g|2���]w�ԺZ!����2���+���O9lv��0�E�P;���(d;,/���-+q�U�mS�i�I�m�c-^�X;���Ë�Bc�OH��յ|RىҵK�a�:�KֻM�h��+�e�/ZL�vww,j�����Gţ8·���
IȽ[�F8��xl�*�_[��6_=飤<����oOۄ����>�z��d�p8v\OR��wN8�ɖw�\5��Mf�l�����y��:/_@O��ν3��S�xQ�|}�4�����7�-�N��[ �xqB�Gz�=��뇦v���;NZFpz�^v9TXP��hw_'��߇%ً���U~vٷ{SEYË����~|�����Fx�{ևJ�.��-��Qv%���U��}Nxc6�� G��8���W���8W�oU�-��E���� ���E��|S8w�1��I|<%͵<%�d��Y�A=�t��y����l�[L{���7�(����_SJ�����K6�)2�q�Jܪ�u��^�&i��[ԣ6K��f������r�	-�p=6:�'�3j�|3(Z)�^!*^�O.h��x�a���L�::#�br�'��ke��6^p�>ṟIy���|(c�4X�����j��LS���wp�fU�
�k�4@�M]���oSW�w;ӻ6҄[����$g&C��}{5�	��Y՚�EeqPSs��[�2�N㭸7J���]TP5�o�4�E�,�S��z7���E�e���7�E���u\���#��̫�� �
��^_�G7��V{�YյJ/m9���&����}��5����<�h'���{R)���d�K�����:���U�Y��`{��[�N�d�o+����Ai��9��i���Gz�V
��/�Gs�}lI3OC܂�=�L�ua�ݹJ����Mn[}�^e�^���{�\+p�x+�i�f�:ǐRc�u�Q�x	������O�x�
���-�{8�Z��,��:�+c�-1^<��*BO�'�C��%�&*�Øk�w��.���3��u��SGc$c��9Qj�N�,��Om�m�����X,��-u}]jw��s0lٟ
�级���ך�זI33��]3���碲��q=�]ů�諭������pW��W�(* � ����D��* �� ����D��
�+��W�@* ��Qv�
�
�+�Q�D� * ��@TA_��
��W� ��� ����1AY&SY�,�>�K߀rYc��=�ݐ?���`�� �)T� ��*� B (Q (R��R���D����騔E��T�*���9�;dDI
�T��URQT%T)@�'6�� G]m�#8.7um�;u�iũʷN���7;�ųڻ\N �@N 'i��pT����gwv�5�ܕm��s2�ܪvn�]���:�]u�@�*J(p@        ��W6�-l�Ju�	h���(֘�)B��t���3Fu�J��#�	%H��+Ll�
�*�r��"T6��0��j�m�%+6Kj���R8�҃	6Ĩ�ZUi�Q��6��X�lP���;�&�2�MU�m��6�����J��� ��5�m$D�f�+Qj����mjh� �K��E6��4Dl��LƉZj�5���RI��TH�b�hi*[224��@Mng\s;Fnv�lp    M�b�P�  �  O�)(M0@hdɠdLsFLL LFi�#ɀFO��U4hM1M2d`	�i��101��&$Ҁ�(F�L�OSj'�z�L�d�������-�7��~I�-wp�4Ǘ;��l�-��&�I$ '��%	3$	 ?0I1	� �$�đ���4�x������8�*I�! ��RD�:�X!�2E	�m�����֦A��O������B@ s}.5e���X��Z��A�zd(R�������%�����kpݗw���y����&��4� �K�R��6�S�CE=�J;[yͼ������݊�R�VV[!�����J�w��U����%�*���]jvV
2�{�q�6���Ĕ4Z(��:�
ͱcs[/z�SyX���&�h�@Ԫ��5mH��S,��U#*�Rޏ��j�5-��<�����y\n�n���H�aYg�l���Ἐ,Q^�Ӫ�0ԑ��%ܺcV�.��h^�6�yb���V��-S�\�S:���6���W$��s v��*���	��e��5O�!����I@s5}yX��F�t��}ʮ�9;��f�{]��@T�u*#�@�	Dq����9L�d]a[��y��n�nfS�uf�M�e��N��϶�4��6�W���b@U��>Ŋj�*�ZΨf�c��ŸU5t2�٢��91��f `t^]��z)�M�Tԥzl��ZA��vh�ˏ4j��c*m��l(F��T�͊��B���Yo@ܭ.���r��1i��[��t��V�	��V��7nLi�#s$w��A�����1����q'F74!O-cձ�Q��C�N�y�wY��2��J6+���U�B%Ll�B���y�G6�+Z��-gHH�(�f�=�r,��w«L0L�ѯZ�l�7$��'�B ɶֶM����(^ۻ�&a��ԋO)ۨ+t�`-����a����Ǌ�f^%ima�Ӗ�H�7x�j�4n�9��G��vuf=Z�U�辺y��7c�yfc�b�X�������
k��^��⣕%�MV�@7�	�C/j`�+q�IM9 �MQ�.0D �[*	�g˽�Ul���+j�SB�Jm�f�o��6��c�AY�g��hK��|�{w���/�;Zu�/o�"�g!�PaE�y���K.1��&͢�2ܼ�e�CM}��x>gE�/Dwn�sV�B�.�Z�]�-C��H0V�7��t�8�ɖC��m)t�en�,Q5A�Q볻|8$q-(=婾��bYy�vU�H��@� ��х�̂�$lI���n��Ym�P֊-�.�nn[I_ǳ����=�ڬ����|tJ����(�2�T��h���:lݦk.բ1>��E�Xg
�.v�O@���$N[vҔТ7�� :�Lٳ�3/%^�y�Z4RCRȫ�Kj���v�7>d���Y{��Õ�2	Vf�Zw	lCna�9����5j�B�����+�чjVe�7j'&��b�!:�F�ݏ��+a`��U�V�m|�W���5eɰj 7���Z��B�W�S�c
��,�킄�܌ұ]�4�����7�VR�`�f���ݱjIB�����*�2��
�(jZDރ��ot�fb˳3j,���em��mSa�[�#-�k5��!ϲm��Kj�r;�z72��`�.�@�T'n��� �ݬ=�ڝybB�Y9����ބ��y5��yz[�[����[��ԅQf����c�$8��m鵘�GwRp�wb�ݻpA��'
��7��^h����̗��ҷְ���]aIQ�9X�����z�օ���Ԣd��t���2�nn��
|�*wB�وЬ�ܘ�HG@3^�ڰe���j�2ļY��ˠ���:�5.ݧ�@-����5��6�Ӯ�+���tR�khǌe�@Ԗ�aR,TT�Z���[�-��I����*��Yf�z��On�|�כ2�VL�da��m=?q!p�����m�����w���^i�REN�M�cv�c*�q��]�l����fǭ�1��i˶�S׆�t��̷vv�޾��t6QE�:^�,"��4�m��v�\QJ�ʛJ�nj�k��G�5�HӸ��"��B�a����YgV���D,���Ԯiu(Z�@�~�L���Y�B0�=��C(��wi+��m<I��g+*�h�bM��$��f-� �� �Y�wv�J��R�ś��e-�*4	�8sF��v�y��F�i�88��%���ʧ�)]I�h�B���V�U�W�{�C^�7�:�t-V�v���J�r^�q	 �ˡ��y��«@�ȓ7[6�[x*`In^�yW W�4��[N��"ܩ�o%���i!B*`�ԫ�	z�w�ːa����Z�5z�G��խ��[LG0 l�TĖC�Dd�������Ksf�`j�vU��۬�
g��O �D�:�c��߭�X�����sN�ʽ1T�0���+rżUv�^��:u�TPx�q\&S����mM�
z����1�(�j�LXT��2
;��u�3�$��-�*���M��x�'�Ҭ�7j���k5Q^��/u��ʴ�^��GAV뻧z͚�r�����y�Z��)��{�6���3-�׶R,4���a�H�,�"�t�oU$3R���dѳ
�6,���Th+cq����f�8���+��ޅ���BY��r��9�Q��*�~���q���Y۲[����7cU]B��]nDY}wG�.�C��4���f�Ok�af��!U��E �ahnf��~4E�乆ł�:�p�c���7��RX�M5ϳ�_5���=w��]g:�$]�,ӦU�u]�����nlX��CU­V�4�o,͉��z2�8���v�-_@E2�h�SeҖ�{qG.�^S$��(����Jӥ������N�>���[��z��E�m_#xqU����v]E`�O����j�ö@-R����H��ߥU��?�jlH���;�6�>>��挟q�w��ْ�)mّ���� vd '�c�Gj0f�q�{lK��e��U��68`)��U���0N]��܏��@~�&i�0N�6� I	�tW;�W��Le�+��O����,*��u/j���gq�y���+a<��v���A��=
�2F,�6�^�]��M���ט�e�y�6��W!�<j��l�p?*E㲃��۝}{j����͘���m�޿Xڇ���(��u�s���jy|��qJ��f���{�+��j��t�Pۺ��*M���Yj�d��vP�m���fL��.#�3��Wy;s]r
L{Eٸ�o	E�t��9��b�w6���Yi�%t�2�����3�ȍ�YLU��d�]����ݰ2C�8]Ɠ�d{��+:�k�N���=Ck��3�[�څ���ܠ7���&�&~�dX�)�;�u^��� -��l�l�����#wv�t�d,�㺄-�AK݄X��d����7�P�Y7�V���-WWum6�Ɯ���5�.�L�KS [�vA�١wӰZ��Q%Ķ^�; W�RC ��u�4+2��t��n1"��r��qM�*�݅�L;�wROa���ҟQ�Z�9YF��F��+x�\'v��N�Ƶ0��,٬�Mv��Ge�e��M�������/u�����wʌ����O4_�e�����*Eۓ^���ʑ�VGq�
��h-ˀAxg�F��N�L��g9M��s�bfE��a���a(���ۨ�b��*d�m7��/�^gJ�w=��{!�1�)�o�-%B�n��ׄ3�3�7ȥ7
���t6�i���i-�Xl��˼y��J��ۏt�T�v��x�N�/��oDFr��I��Ѽ�X�i�pW^���欐�P���m�ڑ��p�9`�u�i��9���q[4���H�ioyN���Wh����p����KvVnh�!KOt"��d�סY]M�*\z���'a�L]@���3�L٪�e!�t�
��:���Ï*����Jj�v�9D�u��N�ut����()�C��wcC8�ABn#r�b�ź�MN)m>��ޮ���� W��q<�`u�4c����ִ@{���t�M#��0V��b���s�i�U9�&R�b��X�����fۡv(��\|6ld )Iױq�Ѐ���	3d�1{��@�B0M�$��ݴ���$B{��Pà��o2%"V�h���Xy�ӧPc���݁Y��mu�'8GX�l�Y.ݥ���1P�y]i5\�)�-������Z����y�68d�HԷ�v
Wl�۩����4�L�x�]B$��.ӑe���u
|�U�N�L�VF9]ڈ�>h�����We��l�:v�/l=.WG�ŷ�����t+^�N�v׋L4��ݣo:�+iw�se�[Z�a�6w�$,��ǚ�:؆=�`����)uDs�S��Nf���n��Ĕ�ݙ$�,�b�:�X2D���i��w-����� �.���*��*�C�a_d���,�4��{��:4�����/��B\v�8v��Wk;X�xR�������D"��N\�Lb=B��j]��YO;#5a#y��'�A;�1:Ь�:v[�/��Ѷ6����G��\2V�T6w`�;:PD2���p���Y���e���"����r������t����#B�1v�մ9�3��	�G5�k��FXں�_Uʍ��7��.N�i-P[��щ�ݵ�R]��tq��u���.�kf��7;x�;$
�.L$��7Z8z���MH�6�98�$��ܺ:�������K���{���R�opla]\�f��b:����]r���N-j^X	��0ć.yt�S�,b��nR�}.G�n��`��I1�:4+r/9,'�9��Z9S�@�o"꽦3����������WP 3x�>�s��se�N�@��9�������2�|_w�����E��U��Ir��b����or[c�K����ΖrؤQV��Ê�n5��=v!�1�t�^����L&�\gu^������R����P� ��\��d��嶬v0��yV�xc^�ݖ�U����^�7*�	����7λ�2�B��hcx㖳Wl��N!�z�)�8��KҀ�o1-��Ƌ=5M[z�ݫg_v"/X]YtD���0��f�v	(��p�G�b7��Фp��P��QN��)Q�����a�{���9fʇ��=�Y�Xfz�'(�yJ>E�ݲ� ��z,�6���WԲ���Ec�lVZ�%���v��r�kk�+-)3F�ӗ��(H�r��I �$F����$�I$�I$�I$�I$�I$�I$�I$�I$�H��ǹ(���2�T��+�wQ	Ү�2��	�`{��>@�f$���b�٫�N4�4R�G�˳�GWڱQ�j����]Ƅ�i
R��U���ӝ܀<u�+TvM	\M�1��)��֞�#2F��V�C7#x���+`�c����GfvW2\nK�3�n�,@�2��W<�M�M@�|ں��%�q^�a����G�ø���H��mu�vh�X�e�nт��g)Hoq��ǬNՀ�]�*���l��oKE#v�8R�\�t�[�ݥ%�]����ǘ������38�e���<�khD�s�(Ʒ�w���z�������:S8�,��s^P4��֚����M�"�v�uY��1V���}�K啻��E���fÙ�#a�6zO�}ߧ�9��__=����I  �g�	>o�	�I����I 	���o���~��O�[��ӑ�yXw���b����1��[�!�!N��9Pb�U����T+5Œ�)���[�U+!���U�ͪ�W��Ҵ��o��k{N ]�o}vȱ��dԚ�f]K:h���\gD�"��)"��뜽�<��wa�zQ�M٘��ih^<R�Z�e���]���X�[��]�m�SU��\u'��D��ˆV��2���I�x9:����q���
ޛ#=.:��}SAe��o5�;�"t�L�~Q	k�8.uu��Y���XM�E�E�cؕ����N�ظ���>�蔈��7��I4��> �9֮ꀋ�q_dTzm�$y�հ�:�ѳ�Hr���;V��"*��
#o�{2�mp)��e-��36��&�#���,��e�c*X�(�D�#gVi�.���C�`I��B��+�sC�%���j��(e�%Y�\�P�է�YV�ޝ��C���ǒ�%�[��gEu�:�T�[�ZT��hmΩ�]���.��#vE^L{�+�ST:��7�/�ҭD�(�O��oFk�L�:+3�)Czv�����4����x	3o"Μ;__mD����̑l�np��t��7ί�����:��+%p^=�Z�I}jw}��T�)�0�u�}��[qی���@iQ輥Sm��j����
O����x�R����9�����(_Wonqa�(ӺN[�G�OX��N�)f����{v�j2=qnU�\�����~ℋ{h�
�8�rY�	��5��tF ��
�o$�n�7R�s��N�'����e��(
��<��>�����묰,>f������Z��e9/�	�q�W�$'#��q�q\"Y��wW�v�a���/ӝ���'b�"qݨ��9��!�Xq�����x��wEeg=cHG�'�`ҍ�=�\��ZiC�\wP֚����]G|�\e^w�u'���K�S�HD_2!ͮ�ȝ�	��-��wk��j�����`�M��y��aM
�C$�pi��";P6B�>�}b1,�W��ޏ.�r�5'#C�㓜��JC��8v�oh��ѽ�FWut�;+j�bVof�\��3#U���Z7�q��_R�==W�Q"�MЅ�rg'8Յ��Sk�=�����f��Z���O��N(��h����iWf�U��nbT����D�8Ws� ʩ��컦Y���]niީ�`}v�E���G��7��U��������yt��rP嚳%�r�ʻwX�~��룯Y�}be�}\g-��7w'浘q�@�j�j����w2���wh�d��܀sB0����&���+9�Z�+p_;��mu��U%���ʅ,��+҃ˊ���^]쭙z@v�a"�#N�=4�ط[M�78`h+*^��|�T��
iŷ2��c�����)V�jl����o`m�,}������o���G���M��#��(�e��K���T�B�[�{�;��3��h�������R�Hu��0͙K0�[��T��)�-i
��厓N%o�������M��n�۽���ܒ�*b�7]�ϲ#����h��E
��9A� r�ʭh��d���W�r1� *� ��%!|A���Ǥ�C�e�VRx朡�+����j��FU�� 7&o�C'�c;��mv�E���ˁ%�B�]�t(�%
�|�6���n�f�M�t]C�{��۽ZiR�΢���`��:��J�Y(�y[�nj*�c��,���v0)�|n̠��Xk��H���i �p��!����@�t�c�*�y;'7!����&����X�9�7fEE���e���b�X*�ͦ�L�ʾ�ݷ)*]�@0nʹis+�s��C����j�9ے��Dk(CG�Zϔ��cFIք�a�W�����n��BA,�5c0X�i����9`�*|�ޱ���*�c�Ttht.,�������o\ӖUP���'l��j����'h
ou��5.}�,�0��Fna˔/M"D���V�h��7vT�	Y�����uŃE���f`�{��wf�p��V�򘀥��#(1�شAD٘hr��Vk(��4l@җ��Z��u����C��s���p�.�m��jI����z_ƍf����T��n���K�"�J��<Ņn®w��+r*�o� 5ٝhǯq$��_PQ�C���t۷Z�:�]���y]:=Y*���Q{�̑�ˮE)�đK����:.ȓ�d��ĩ�!��G#&��,˃*��A�єh�#�y!�z�bC����4]���e��%0g>����wM�굣2���<�mˡ� Í�˯5i
��k�����C��t;E���x��;�����(�h�� (J;[��Uo	�BJ�@z�u��%#&n��tqVh{�xI�X�R��4�'P�tp��
��j��`�鈄�C�3&{-��ʗ��0�b!|mT�P9[��5�_wqfLw�oiiT�U{705z�p$����cʂ+)���)�ku�f�VV�<�9M��k��Ag+\F��U�JS<(vgL�ј3���pT�e�O���%�;U^Ǯ���Y�����c:�ۧjq����m�̟B��=�o���qbw�����RƮmj�6��hڶ�ot:*Yn�?�Fn&@��p�X�['r�G�̺laʖ��x���V�3/%�<p�Y���z	fS%uu�4H�XΘ6^c;[��|���D��AY������pO{a�g�x׽����q۝��S8�W=���b�J0eNb��v��#!���F��=���k�Q�[Ͷ��N�Oj.��F���-j�+{[q=HV^T�:.ҧ�`ʼ���[�`J9��V��w�j�R��^�q*;'*�_nD+���h\�P]K-ȞV-7ˮ*��z�u��N)�����K*�ą���n^;��Y�qC!G�U#g1��8����]�5�uͦ9�	W-+��E�鬺���$�7�[��W*�vs[�Qm�H���5ei�r�H�H���񻿢�U��(�ڴD|��E�.���S-��Å�͹eT���,����:�;������*[AE(�0��DJ�v�1j"ʀ��r�F&3��G\TˋM2c4*��Zcu�e��c:�բ2,�-s\�b�[6�R��8�L[�0���L���r���T��%�YQT�q��ýXiΩ��	��&���SI�S��fY1�L��6̥A��,��&1A�K�T�Z��a�U�Kq�,��d˂�
-[.-1k�ف�E��b��Y\9p�"`qi�V)�Q\�7
�"����N���>o��֓��߳�|l��]L�m%sfg4�c�C ������P��'���˟���3��_;��g��ΘÞ�f^�E��Z��^:5�缾{����I�o�����k˔On�y}Lw�l��Yڠ�p<،��6��R�"�z�u�᧾�;�Y��o����)�7�/�{j��%ퟻƨ��I��RV�ׯǉ�7�N���ӯ)�)�)��1V&`Bg8FBiЫ�}ۿd��b�f�>:.�K��x.<v�p!wa���y��g���ι�s::v��7x�x���7ef�^'ѫ�u���X�`Ӏ��+w?37�`��9�z����^�P����d╨(�q�N�N�`��aYJIH	!ߥ�W½XP��
�x���+Ce����1`�h�Jc�r��<���z~�Ss|��.l�f���UM<*]yU[�g��t�u�y�^�Ywp�q�{�8{|O]�����zcSǾ_|�]�̾�p�7 �<�ez���_��j�za�dhɈɩ��[�(��O�	r�ˆ=�:|f;�A���!�[p'˅p���Q�"{�C
j'�;-�ͧ��0*}:=MW�t�0�����A�0�#���z�n���.sO��O||��]��|@�pu�^�MoV�6����1A�!W��-��3%ېEr�X��eM�w;d����%i/��m��u^�6�_Lɝx&��G�ȁ�;��1�&���ff껿"�Ga
��F�+�5���}5�7�ryn�ѩqO^{MY�8|��Z �+[�����4w˴:��̛x�)�wÛ��(q�0����ڄTơ������׫bՃ1uY�)�@Eh�ab�.g���m�p��x��r����.C�Ҧ5�5�v�q��*!ϊU����nu��"$���7�S�#.��LA�;�u��!���B�P`� ���;����o�3/[S�+�ɡ����<�1��W��|hR�Y�' �b^cג�7j��ц��n乶�QԳWC�z��H��<,l�%Q�y��qȸ滯50�qˆn�x�M�l�����jz}�tDd����s��m��e�w/{�/��|Qу|ɝr�'�f/�W����0z������fs�
o;�\��g������d�'���R�X83l�ۖ8�7})�W[o��2�3�l�o\��j�2{M���\�����^>�dÚ�0kxX��=�䐖Y����'���4�}OS�2�0�<O<μ������^{����^�g�8�;Ki�y�,��]x���8Ü����zN���3��k�"�l�w��J�i� �ج��4��|M�jL�)��m�e�i�8��;�f9x�޺ߝ�������T`��tܹ3����τP�e�ܽ��}�{G0���s�c�S��>�|)�v�ƅGL��LB.�P���y���l֎���IZw�o�0 ��xO�������U���~��x�@1�gB1D|*�h����k�']�/5S��l���p�>�C�r`���ͽx&	g���;��I���
3H0����;���=�reό��*�4��=&0GR6ȍ��P����ǝ���z�<���_��9�cW�-"��5��æ�zSu�^k��9��g%p�:e��`_����̤����'��.�V�ܧt/z�=L�{N��1玱|����w����|b��\����h�|{fr����W��x���)���PԼ���o��]ם�����i��)�����f�}�/���7�ÎˇI���Ɉɍ��W�U�خ��̴��¸1TD+�6~���}�Ǉ��|������P@�`"�j���\���:eoa��G��e�4׭M��1۔�{��s�y�i��28��f�@�T�����Fޗ�rp֏��@�֊V`�*���[�v{ݎ�+�h�X��z7bs�l�fl�LVt�z�W�Z�j"�a��2cqf�;)۳~�_�⿽tF+��R�O���헃�}r8B��z".�70$0��2���׺'�T�����걬]s�F:�ݧ��ﭴ��I��.}�70f3 \����1�ۂ�t�6�Cư���[5�G�X��X��7R�_����7�M�9z�ݕ����Z�o�g}��:k�w�u�{Lj�r�������ף�ݱJ�u��t[�.�@�y\z�v)�8W�Ț��b��R�U�pB���F�ƫ�΄!�G�M{X���C���}���f��8Kfꆘ�n�mZ�{�i���]Qn�ӔM,�B��y�B�r�x'6���S�x�ޡ�OM�˴SN�N�������5�:z��<9|g�{w�q���٧s��[�������A��
�����6]-������D^8��򜝞�=錞��*���6"5�W^�E�띘��+��Tp\f�<�!H���(����\+4ح��i�z��xx�m��*jؠ����n�|1��u��-��Q�
zm��S
F�.F�D�o�3hGK#e\���n�T�K����ߩ� ���^T������A�����×��jVe3��?:���z�Խ���(F_o�n�j\Cz�[�WqIwȗ6Л0�Bd3����u[ݞv���Ä;����63�C�y��C80X�*~>??!��W�d���R����ouM�]��S.;M<M��/��Ȏλ��UX��K�AX)>�b�5�\;�G��Y�W��>:#��o��{�s�N[�c6e<9O�=}z���[�4�p}�Z�|
��
�7i秘����e��pr�+���>�����μ,1��_xT]�7v����ɇB=3S���)0��^��3��5�^�p�h�>cS���h�ߝwxׄ��̝'ú�+W(��� ��X������^xY[��t�9z�*Uܝ�)�*r��,$V!��r����d�ߖ�FUЩ���錈�ˌA�|)CPc?m��|)�Çњ��Ikd��n"���3v�u:�Zo�X�����i��t��CG)��~��^�|������y���l0�v��4�=}L*x�s�9��~˺�^Y����!t>B�%�Er�ݴ{[̚k�uqE*��_�k��4>�k���W�o9_��RF����uAJ��/Ƭ|�3�;C����/�:<5��*�5`񬜫|o[�3���S���u�<L3>�y�yp����A����ݟF���_�뵶���/ln��!�#&�eX�E�X�9��7��pۨ�.+�.��VVDkn�in(ح�1j�r��I�[�Ɏ��yr�f٬✛�P6���\';{����0m�kav����Nk�B�gt�ɧ�R�a/kG[̉��B�$a��� ��ୱ�{X�5Y.kvc�5Ի�[�Ҙ��9!�]g����fF/(�4t���Ḗ}�c:A5W	x�c��_ʭ��K��;����i����BT=����޶�G�$�NG`xe�����ՊU�B����7Q��n�^�1�;�B��B�ץ��K�D�v�/��#w�I��Y�i����T_�fl�ӈc��H��}���D���J<-��QlVj�d�M��~]�^sw�e�4!4���eF5�u\Nv�D��8o&�6V�7���Mgj�E=���][�c�C9Nv>M��R��SI2x���c0f��X_<�I�s�rV���AR�e9lϞ@�3�P��N����yҷ0f�X�ۭv"����+2�@�o��yQ����2�m��zr�bH��o��'�%����5R N�+D�fr}	��q���5�y�k|�}j�C_�n��+D-��%\�b˄Ep�DAs����a01JƔˇ%2�0ѥ�1��Q1A�R�j��Ჵ����L�mJ#�*aÁX��lj,��f-�Ja+�&+�Uڈ��[�a��0Z��ִD]YqJR�J&�L�\4�Q�Y�W5DKJ�q�V��8��D*۬�1�0"[Kf���*(��\�E����0�*�*\R���qkNOn�{̯~��m�׷ˋ�1�7����9J�����}�6�}�����'�}��"1B5��"�P�����ϭ*���l���ُ�8�b8>���/��lӾߟ)��)m^���p=߷����>3/5O���n�'SNPޮPǷ^]�}	� c*���+�e��֏�(��ӕ�M[�|�1
���C�k���;Q[���I��3�C�|�9��/��Z�/�7׻t�ei��������Ä�2���^��"���x񞳛���O�;|�}|���U���F�=i�]��h6�f�^{y�׻󔵫�L����bE�&s�e��$��n.������ث��r��ݗ fc@P�k�v�M9b,�cIGe��?&����8�uƪP����i�힗y����y��Tۯ,5�4�������zuO�.Y�[C�];��s�rs�֏{�5øo��(z��M���߸2����ox�=�^��������C�L���~�߹ֵ�z����1�x������Ƣ�M,����J��OS���i���<+�J�.{�3�:1��)��f���Y�ic�B�e���>�������Wg�M|��~4͊U�T�����ʔ��*J�`���� ���"8�ʪﾾ�_�\�wQS_Y/mn���7�tvAH��#�t�"��oI�+3�	I�#���;�O5v�ٷ�(i�A<�z������G#\�����0^�4*�(W��ު�v`��˫�S��@�!Ϲ��N���!��-wU/K��������S�^F9��^c��b3x#FoO���<Og[ǜ���=L>�NX���x�}�|-���v�����O1O	��p���ЃS�V
�򪂻Ɨ1;51;1�[0���'n,�;)Ǜ��yC���Nbe��y���(;�r���Wa����:?�P����pg�]���=�}�pӸ������b�̶��|8f�_�֔^�^q;f���2����ٳJ3R���G��iџT�)�*���nߣ���iˮl汛�]󾚮p�WW_:~6 ��[�,zуR\�%�Ϻnc ��xO��)�Wz}����C����/���t�9p3,=���}��}�ξ>���e�q�=v��Lbr�
�} s��1r�{�F �*LÕ>V`e�ޒ��7"|T9�����N�C�`���σ���'S�ŏ.�h�0�󴺡����8a�����P1X8Td
c��Y~��F;I�g�˫����)\{ӆ�L�Í۶�f�
�iT��Vڐ�f�o��7���G�<��F#��G`%dX�4��=FkoD��#�(����I1��t���x�O7��{�x�-˦�1NO-��kT����ѫ?�]�~E��6���O<PUT`�����#�Y�T�g]'S�u��n�k�e�כٜ>�Y�sM�����6�5ۮ�f3�u��Vwc��醰`�(
�����r<��=��їˏ)�,�ｾ']"�����7��.f��}�q�f�,V
����Q�3o��O�T��������=�_��3�c^�ٟl\yp�g[�Vo^�U���Pk���ѩXvX�FV��;���3mu�{��S�D�l-(N� ��u9i���kɋ�mO�}_|��7�?�51뚚�=O��Α� ˽٭���s�`�u��4�g\��]+Njl���'�����Z�OO�����;0�V����6�P��m����|*
�MyS�z;���b�CGŜB��4�C#��|y�z�߻��=��K����~�H��͚�p�����c;�Z�����*����"���A�k� ��S�LDd�ٹ7&}${X�XV�g���W�y��Ƿ�k���0�E*i|�tQVڃ>3R�&�rg�I��4czP�0Zu~��o5��F���ӓ���Nv��4�!�gf!�0���)`�ܚN���At὏�o�_}Tw�k�xi�T�|�p�ܺ<��O��X������ڲ��}�k�����}��S*_������>b�T��&�_3�/Y�i����s�=.��^��	�#A>U�������i��]O���v�M[=r���7�5�wk�o1OU���Α��¥
����]1�X�ԄmW2ҭ>yʀ�uj�|�%�R���b�����@����G'�8v���5���;z����8��_u����K8�9|p�4�l��omj���<�op�N����:5=�W�e��ށW��J��A�Z�I���
�U�+�I&�#{���@��7�t�߭�x��8�L<�;i���{��y�{ڝp�L��������Į�8���f��j;UB�^��+D9"6\��Ef�7���]/�@Ulx}��S�<z�{z�]s�y�s����Wo��>3ƹr��±��ǝWH.�*�F��H�=1�s�s���v����b2h�5��C&&cf*}#��,N`?J\�/�hW>Ӽ�a��h��L|��m��n�����g�Hp�}�8a�>��ƥ�޹�ka�4�VtT�~<)�w��Ŏ�U�q�5�D���v��܎�s.�b@��3Mv�j�N��5���R�مV3&���U=���q�	$����{�|~ �`��n3~?��{i�c�������l�g��'��r#��CF_*O���
�Q���C�A���g�z�r�|N�Ã=�q�;�=N�������߲vn&�"��y%�')�ǎm<M����]��P�x���:g���}6�qա&�-5�W(+��8�;o�˞���I��D��F+�U1P��ڠ�{�u�jq���G� �L@��7��/�G]���UJ�* �b5b�0}��U=:�["�fJxj�yU��yV;( A(Ч���b":Y+d]�`�ҷN;�[�0���L���ם,�V�#��vZ��)�6�!w1ڰ�rK�{ޏzoo}�t���L_ʽQ���S��f��ǝw�g�Y�l��3���t�ѓ1U8�D��?z��˄8��b���r�꿽t�;|�̻�ȚT���_|����q�Vo^`�t�fo�ֽ/9��K�z�
�J�=S�>��o�) C���E����na�$A�M8U���i���l��ݘt��V��x|ߚ���� qE
���+'Y�J��n�aY�%L��a ���,�)<a�f
C1����z�R��aE�_|��g^x)�f
AdX���$�(T���>\0�§P+�ve�C<��
²m� �3���AM�!�a�e�Χ>y�h�H,0�gsH)[M@QfJ�d넂�P2c�a� ��L%H,�
�'YS�o�H,r� ���1�	4ӊ�U[�[v��	���zj��lb������Y2��ˏ��恬,V�qĐ�aX�Q��-du�eL�ssv���<QsJwI��h��V�N��@Y[��bm#qm�V�\�:��:�Lu�R�3P7��ꏕ�	��nm+*e;zV���ct� �j�E7o;�틣��i!:*�)7�3o�'x�����dQ.9�j�����]�`�ե�RZ�:���J��Iv8�땦9W.�m�Xs�d�Z(vpr����qսT䓫��md�X��GB�N�,m�x�6e��q�g%�̋NMɗwrKCv��j��$��:)ҝ=�)>Mj4{cP�c3gT2��z�b}�&`if-��v\,l,Z0ӆŭ���F4��'	"�[�rr�wՌ�V«7Z�*�>G6�|�PDbS9E����Ա��F����.���k��ΎZ�g057.��\���B�����J�y��nP�L����jc��6�K����`�]��Zh�^��(��F�*Vc}��@R(-��s:���6��%��c鑘ZȒ�b2H���H"9C&��᮸;��8ݎ��aCu{�J�]�s~ϟ���yS.?N2�O�T\(�R�m�ZR�)FֵTk��ժ��,*%�����p��*���\*UE��F�D���T��V�e*�*b�TSV��Ek,A`�b	P*hņ�%]S	�QV`�������)�Ա[lTQET>�}�9o>�y��מw���1�'x�j�5FR�:�������%���E�z>$�
)�gl�T
�Sh ��
�Xi�H/�J� �P3�� �c�'sa�"��P3r]���s�s��h
)��6�)��:°��0�P��ܤ6���$��%H,4³�Mb�R
S`�E ��g^]�|�H(J�Xi�L	 �Ö&PRg�&Xx� u*AdX�C0�P�q$aS� ��*{=Ǘ����a�XT=�	���
)�e�7i�(H,�|� �k�a��Ps�0�2x�2T��i����es�����%H(
,�eO� �a� ��p�R
{�S�g���+&~Y���R����g�&�/Ϛ���ι8�AO(�R�8���H) �(�<jm�0�Ay큆T6��
�a �/ơ��6�S>|8��>o��<fY+���
ͲT��SI*)> T��R3��AH.Y4�@QfY*a���O��Oy˞p�~w���0��Èa �����f!��Aa�
�*AaXT
�2�R�0AH,�a����=��d����^�����P��4���H(|���0�<B�a+֠(�u�;�
T��i�a �)iE7�������|��a�OP*wL0�
�qHT������)6��`H(J���
�偄���E%B�ٖ`{׿+���&nV�����L5֝�'��U!��s�r��R��T��
���)�w�s{�D�������Xi�a� ��%H,�V����:��R8�S}�a�V|Mf�))��%E ���a ��T�Î��o���:�H)iP_0��H)�bì+G�	<B�ͤQa�:����Aa����Aa����<׼���ݞI�T�Hj�
AaXg��XjO��Sl���AH/��<aPٺL e+"�E��r������s����H)ߔ$*Ad�*A@QL�T�f�*i�a]0*AH-�ɄR
a��"AH��>w�����Hyl4����AH.-��(�ĕ<g�0ɣ�a ��p°�����QC)*u�Y��ό� ��
��#�����M���Sĕ�L�T��R
zΦR
EiPƤ�3	��E�0��Re
��=���oyϚ����
,6§�
�X|�q�3i���sHTu��*O�)�Va�R�Z��TR
x���n�w[�֠q+�*e�a*A@Qd�ل��R- ��4�	��T���q�OP*i���O+>i�q��ߛ���{'�<a_�*
A@�%x�QH.(
IR-�ܡ����n
�c4&��0׶H,<L�fXu�H7O��ϙכ;�i%H,�¢��*i�<��AgY*Aa��d��d��%E �P+-H)�3�e ��%@�VD$���s}|Ɵ>o{q��g1��F��+��Em����9�,oC�6��s���Uf��n�]Ȯ�N:q�	�� ��ι�'Ă�a����H)1���
�<��OP��L��Xl�6�R
¤͆
AH) �P+2{����yH)>!Xa��`u��� �Sߖ�H,�2�z��P�۔���� ��m�M VL���s�oÝ��y�y C��6��RN�=I8�L�Hl͇���ה��0�$0y����i!��
q�a��H,8°�
���0��*A�!P�J�k"�Y�6�3��,���L
� T=��|�;���i�����6�&&�	|�_�F|8W
�Z��]˺F�qR��"�(����d&v�	x:���Yr�Mp�ゐ�+�A�o�ױ��#@b�;5�5Y���,RR�1��j4pع�;3*0@@�|#���mC�80�w���>4mpB�4k�1CKzU�l��^w����sR`���L7�*��Zfkk ��9ݶ��⒆*����[��V��oB�.�qG�ވ�G�>�~��?��K����Dj���:��>&��qv̲�x�1�.l�yK��u�9��z�8`����:���in�km3�bX0�$"/m\\p�9��4T��l��,��k��������PD>vwO�h������b7���`0ׇ�3�`�����u4�2y��멷Hx�^`�� ��疰!^��n���i��u�L�11c�Ct=�B� �xN����9���+���̸c�ߘ���9K�s���ju��0`�0q:�tL��۔�7��zy+��R��pS�1�N��j{�ސ|㖬 C�p�U	�5;��*ZL�/y�G3�U}����{��z��3�#&(���}^�ޡ%�}�O�����z��{�:&�Ӝ��j�s�]E��*|��}P����SZ$d�>r�'���:c���C� �A|�&���E���u@��31y����!�\��ui��tQ�x�!�o�F�����Z��u�y��m�D�:ﭫS�����3g�j:���� f�a��s���݋:M�e�N�h$�Ĩ�Q�*��v2�p5�*����X� ��b�J��rl�侈�DD�[��|B��~3{��k�V_�E1���h]P�X�9��;P��i�#d��n�T�M~+"[8bL�UA��ގ0O{��Zz���{�����G�ԭ�u%�g\^v���0QY�4��jĈ��v��͚�.�s�+�y\╰��mAaSҷ.r�����Q�y�^���MD�ay��߉�R9�*��'�œAo�z��U�W:�w�Y�n�(�G�T_*@����5����F	ꏦ���u�fӡ��K5ڡ�oJoo�*�͞��:��������Kn��'�-��l�~!��$�6xB��Z.�}�v�"�Z�蟜(�Pʞ0�29�.F�-Gv,
ӳD���)���$�6�Z ���ٛfh�W<cZ�Z��,��U���J�Ԟ(���[n�����-����t�=[Ķ'����g>��Ws'^�82vn�qa�(��"#��Z���NA?t�џ���R��\����/3IxP9����	3|��-H�(�*��<)%	�d�k�f�؃��4B��zPx�*,�k��6�8y��av$#+���' �$ͼp�X�on�ww�3�=jL9{���]M�#� ��%�#��u�z�.��`���9hg��V���$)�P�)P�⺶��gG�v�seCs0����3$l4r�<��z"#��͸�u�Xcr���Q�!T�	�Dٔ�ڬ�{/�����e�k~+����v��ŭs}�`-7i/8�x���x+wP�6�iD�}�����{"�m9n��f��R���ްd�\�ťgi�֥ Ů&+!'�3q��ةjIy�Q�1��G3.�!�����}.-��%��]��\Z��F�3�7�"F�����q<ފ���]��X��ʚ!r�]��pQ���K�E}��zn6�>��š���7����A����YM�N공�	�k���Aշ�I�\�
�j�g�L+�N\ѵ�7e\����^�o��qK*Ȏ]����N-��x;�%�(��7j�L{��8g��姅c��j�!�o��3�F�m[xpKK�#L�x`��@"*ۨ=�8��?���^t�c�ZV�~+^����ݱ��͹15V���P4��ۇ�B���F �m���b�jY�t�
	���_ٟ�t[67�t��H�v;ܳ��u,Q$n*�7*'��|��y��T/z�h��Kn��mkQTX�'qe&fV�H��8�AS��m�j����x¨�D��li�b�7��iw�Ab�[sG7�g�b�.�9��.X�z�p,S�v��,�Z�
�Tiut� ��Eyw��r�����u�ۘ�띴�NX�>q��_j��
͇(X��6�0���.^5"�M��_*�����e��*�/k�+ G}�G*��.yD�y�����
}Ǧ@��b��F.��;�8:y�2d"��^FDw[�+;Y��u��Wi�N�{{�*ԗ���62����:��d=׹Bc�#f%��:�%҇`� �~�w.������oY��#%�g�S�3���
,Hv ��7t�&X��l�n��	��1W�i��f6oǹ ����lF�Z����G�K뺽j�����L�����ye�N�H����;+fN��H�Ǥ�X��%/3d�6J�ea��	��Ch��\�#쵲t���Z�>rK�M]��R�P.�dQR��).�YZ�[%��,�*,cR���8��T�-T
�YpR�[mkb��ڪ3��0T�,Ch��4�DDX�D\�sj��DV�"a�`E&[PF ��K[EV���A.����z<��7W]��!�����t�D�E~�"=��i7�=���ř��k��+&�)=S'���8�u�����ag�_�TH�*+2�~�>	�1�o�|*e�땮/+P�;���EZ��[|1�S�r�<\[�T9~)�mn2z6�׫EMv*�|�K�ԗϻ�B���}~�5��>ӳ�_�(}EVK��)�]B/��y���F�WJPo��7y���R�5���qN��DǹG����w���oE�r��a�R�_J�EE�j7=�!���/��{���e��OّE�n�.����]V����X��\nf��ӿQ�M��,r���L�+�]8�N]��vu;�Mĭi�J=o��k"V�ڪ�>��U��S��*gZL���ў�N�tZ9`3�F���[l��Z/+���2�Xh=]�噃c@/
�g(ā�ļغԂ�'��y5��a].����Lm:��GW^���q YF��-���U&�.I������������OD�>;܏{�>sd' �o�Y���F���9�*��
���K�wqF,޵鈋9D*|��<0�e���'��b"�pyD��1�)�ք�A<w4��[[�}�4��3�����j�W-�	��RoXCI"�d¬d���[�[���5��D��{������~��th���]^���	�V�V^�%��1�W�i�J���
e�h�Y�ʲ�@�Q�g�:���t-�� ��g���qυ�1�v��5vkh���|$����� %yP�0�z������>�����9�k%�f͞G:��4�R�0�;7��;7� �͘�qP��yO)3s���p�{"g��@��'Vj #S��N
t{.�=����b��TW�]��E�m{��9甋V��̎�ޛ��p�VGM��h�"�$o;J��W�-*��Uݔ�=)��5�
���^K��MI������U}_}0��~Ѵ����ƈuv\�{��&s�#r`A�$XW8�7M��ѭ;�a����D#�*���.�Ƒpx�P���G@:�:��{�	;|O����g�����ε���<�b5�q�U�}-��%Bq[ڻ5�7$�ⲭ���T�!8��N�챈��
��{Z�p�ռ�h��m���/��I�2u�V�(^uP�,�弴 ��7�%qB��_y|�<��=舁��6�����C�@J��w�W4g�Kuo<˅�Q�m'�gn�6��z� :Vx-Op5��4�����a^���N#g03���p_+C��CN�W�F} ��ȕ��^�vv� �1��彊(�{��5�=xb��7�x��_�2�*�V��{a8v{8�F�l ���m�=Qp�}����ex$X�^U��!��l>��˖��4ݨ���"�,7�CFn�3.�t�s4b*���%�?��U}���Ͼ��)j�tvK1W�|�K��a�ܐ0���j¥��9�L�G�ݮ��Ik�VJ��\(iRGjGC�w���7sf�ӀsĲ�*�y�xW��!W�-�.�a�}���[	��\T�U�G�������(P�jI�F���X��9�d��v��7�h��L��D*;����w��31&�tG5fY��=0��ǐ��&wZ�F6u:-0� ��$�_}��1�6��r�g�Q�.�+�Un[2�wjڠ�{E��(��~��ʆVn��Xm�umu,�㛦ֈ�\�����ni�`ۑUr�����+��(D���0(h_�������6���@�.�K�9W*i(t�^*�y�u��+�x��ܫ=$C�SQ��i�Ƹ^!���x��t���"�Z�������d�_�[L
U}�� b�}Z�-֟M|K��-m&ި��kɚ����}�S⧽Y� ��g�����`�� q?��l$�\=Z�޾�칌|⑾	�=��+;����f/G1����Ɏ
���_��)/j��w�蠱氏y9X�-=p�&U؝b���k�L1&+��{|�Vu��,V�ESR�4
=Y��k1���y�f
a0h��m�y�Ezn�5�@v��O`�[��u�ˁ@Ua��y�2d��$Yw�R�"�˩�UƷ�ɂ�iV�G����%���/����t�F�N�%�x��r��3����W.���(n���
��Ȟ2r��WM):���x��B��B{�2{�{�Sϋ��z�T�ˎ�S�� ��S̘�w�c>��n�v��wwN��,��}��J�3�B?lɷ�i�W�T�9���.���f���̫�$C\#�c/�=�rɶo��Z[P�sD�� 5��ZX`Tdwڱ-t�{ze��aL)h��G�
�>븭�Ԑ�X,�.M[��5,T6�ø��ӧ�oz�82Ѭ���:���̫R�\d:�G���.��Y��gU�-�yD8���NЬ��o�0�CW���̫m��g^Xn�F�C��$_d��m󗄳�F�^�)�$
*�#���;1#�vFۧ�bBS3x��a�쭼c{��պUa�m<�Y���|Adh)�6�)��Ε&;(5R����_Nw��}{�����+Em4x�
׃*�"M_ڈ���]�F�y5p�!�|��3oq��KP�[y�^�ZnJ9G��Gw��vV��AxL�^��:ԍ�mJf�O/�VD_v>.���q�i'�v���U�v0�iP�v�-�;�"%ށ9�T�9@��/>@��r��z4�v,�#�=�D{������u-�`3�,��E��|��gW}n�!��M�tu�P�����I�"��]�<�Gfv�B��p��'���A�"�m�7wDZ�0��G��G,J{]��ԓ|�:u�I"�/is�q^��;�º��T7�RjĈ�Xs��&NG%ou�/�~��,QR*�k�ڢ�[�0,ݦ-TUR�ҶՅd�����J��
�ƌ���Dc�miL�&���ˁ��PR��Ky�D�*�	+kZP��lie��%��+U��*��[n��ZĴ,�l���D��(2ЩR�-J-�ҏn��E�����j��a��/#��ÎpM��E��:���fH�qA,�75�\��qJ��ʺɁT�q��3�cE��`U�TZ}x=��P���_���FCI_��#�i�v�z����b5Ѫ���=�Xȼ�j�tA���DX��]��e���<�x���%��,�J05m���tc�x�oD_�Ю[b�n���r^�
�\e����$��<:����2L�c�w���Q���lR
��Ss��.�vyT�J�W6g���z=�ZۂD.��\�K��`"���+���g�����8�~��t;{�1�3��⤞�*>���&4s�e�q�A�ns�(��B.�E#|���]G	|�����m�C��f#�(���X����&,8�a��o=������(T��=z\ωڼ�Uʒ�wU� �}N�((+;�ƍ`���X	`�����v�[ᗉ֞_������i<�%Q��N܁��
�{�����DI߾��_�����7�vr�0mn��%R�T,�S\�zYkb�ݮk-�|�}���Hg6jQ�6njJ����W.���f �d��j�w>t������i,�0 �a^�|;1���%�H�a�^<ak��[C�y!m�L���;�
c8��318sa���=�,�u�Y��m
'$�)�������h�
��Sl�^kbmq�͒�_��wj���7�yq�1�N�PR�����*�s��{����G���~B�U���;�9�g5lO1�2���.t�ݞZ��c���Ү}�^>��;���r��W5pN���dy��v�nVK����頪�R8�U�[��~�����
�`�ƕ�p`#��v�5�u�7�����Ϡz�ߣʌ3���v'�qTBb��|_�l�_AW^r�xޗ�:Ң<Qv���1։�	��>�b�]֭ͱ\�y��ÄݪI���+���c������>���O�~{����/(��_�7��a��3����Wۦ���Y�
+[�'y�T�Fr�%��Ͻ����1�<��W� �#^�>E��]]�l��P��3�S8{8��g&9wf�f��O�n���(�gi�Mk�v���-F�ifr�{R6(h�u~=j��"]o���v�$7���� {�g�~;K�P�<��r�,��'vl���ff0M�BjO���%�w��n�~�9��jЙ|�!�Z/O�y���lC�2��]h!�|O_��|E���X�.��� ox��(S�9JJ��Ι\fj���pxdKڮc�����w=I��{�v�z*�}-�!X�g���T*ň�NNP�K��O7~�fe��M�E��Ɂ;)r�G��<ǅ���{N�*Ӽ�Z��^>�J�,�rZ����ǎl3���p�W?ȃ_>q��� ?ξ�}Sh.͊��j����5�,�����΁��?o�gow���5��O�-�Xk�����2
Ȉ5�j���,���|�y�Bո<jb�J�3	Ѯ�=}������ƳF�921�y��^{�7Hvk�e�$:��h,�q�9�[h�8%]��3��� }u:(z��8��Id��ܨ@M,\6�������>�V�x��,0����Ϟ���¿��i|8��;���nn /��)~�ۜ\�}�)������}��ל�vZ��=a1{�uOZ��>֗Wc���A�kQ+�O8���8k��$}ٸ�w���2����)覲Ѯ�� ���cC�V�z�n���P��]���$�6s�Bp�|uk�`o��nX��y�Sх͈���6���k��O�8��ݲ(�]���B���<�� ^��o�	��w�n�\��<Qo���Z��ї5�	�|tvo����g7F��p��uY��Bν뵹���y�����]Ö���@#�֗���$�20{�85�v�,o9ڗ	�;��O"�*�ѷy|k�GJ��5F�cil"��nUݿ{r��at��)v�֫����^̱�~>�lw"�:쁠�r�6��u�}g��K���|�٘`1O���l��?C�De{�Q�h���T��R���s���a�iAx�㪁��uu�C~�'#N9�W�օ^42��v����+X��:����p��~΀���^�};w��P��u�2�z�s��RħBk!٬�e��w����D��ǵ�|��W�yl3�s���+����bc�ߔ�^��.Vc]����t����t���16#b��wU��D,=Q�t�E`�ν���uֺ%rtsS�-��j�^�J�]ǵ��+;ܭ>8i��Pv�f���.���h������wP���9ֽ��	dL�e���DJU��V�<JZ _Sz������nZ�8c7������]Lo�,$�m, ͹:5�:��K=}8��&�g,�jr}$�@��BC7b�t�5�XL�t���Z�W�֚��6��l�YѢ��Pa%�z*]e�� �Qַm����@�0�Ƕ�ݧ��/�RiD�ٵ�llp�2����o�8�څj92Vl.�* VJ3.�(d�mg
z&��:F�-nV�71_4�c��=j�dP�s��������~��ao���������n�#��
�Q{�MF��'	J�=���k"�1�f��g^b	ؖ��1�����@��<������u�Wt���m���=�:Q&e�Q]��8�u��evVa�m�7b��ܧ�gi�5�\�}�4�|�)w��"W3r��t["۽�F��9�
����nV(].��)��`���5ՕyVD)l��Ǘ�����D��ѴJ*T+V�ciAZ�ҕ�*)Z��KV�m��mō�"(��Af
R�X���H"U��a�QH�#Z%e�V,�jT�5���u�E��m*��������

����-�%C�_9��ݽ��ys�G��o^7�g#�%NG.>H��rO�x|������c)<��Gu��/�9��o3��1��ys�K�=7x�.d�fn�ϑ����+����ԡ�b�����9(��զ�M��t�d�p'~�l<Jt��=@K?c �;�>a͙2��b�j���y�������=J�UזQ�R��|���M��8�>�o�(j�{d�ׇ.���u]�5�;bv pLtz���3*������R����
.~�����~�^�ʹ7���6΄��v�+g���4oMgcjs�Z�ң�)戺h<�](��)�~�=91�塜7�ʦ�8����*>�4�p��W���1q̸�]/�&���ͧ-ѼtuYހ�o�6��U�X��W3��}�irG��U.�Pj�<sk����P!������:#clK��v�W5��4Yz/�y.�q�{zרZ�	����5�gTO*�L���I?U[A������#'�Xs�<mn��IuE��,��E�x�އ��� �}�,L���g��{U���ݚI�+:�����a�l�gE��^�g)d����r��qݖ�������H�8oN��p�n���//�Z5�����5��p(�+�6�=����4V�x.��Q�M����E���"(������ݻ��V�����M=�:�NB-��t����\f(�78#|y���9��	��.�K���^;��Y���W�Nل-k)mN�lo��.�Nޔ(�qn'�[��u�[�8��1�q[���F���z���1-�k.�u��b������x��ǳ@���vOb���{ճc��O&��s�!~$�S74u>�k��[���������_a��ڐ�s�J�<�2(C�s��{�5mht�f�x3�0���Fn�pe��T�׽�S��3�mO�:l��QZ��$�܇Y�A#]�/>�c���|�5G��bF���u�վJ�U��]O.���W����x�.������T̓D��2�a���9Lv���^��v�T�<�����;Ec�Κ�k1����
�g!�/�)��2�����cnFN�S�{/�Σ�;�M�����(d��g�W�{]�u��:$�bJ֞�H#ђ䟪�/z�AN�p��%vpbv�"�t:��^�.,D!y��q�y9�fz�!Qi���3�:%��\�=�B�B��	{��S��-W6���B�U��2��9W}yNy���g_Tq���e ɥ*R*�(N=��q��S��m���՝G�V��>�}6�1�N�b����4#��W���ՍT�yU̺�^]QD9�+{E���5������L�r�^Aִ�_Duw&�_��	��o!�5�t��^��ݳ�쥝o��/�4�-^��wW��v0*����=�M�f���N��o޼��7�I����\g���2���]~d,�$�44q??k�Cr�ߗr:�����Tl�?b����_�]�l�hy�XG��;w��<���'������yp��.�up9���q��K���.�뵅��^�EM0}�}�wXِ"�ʹjX9t�Ũ\��At��*]��Y��돳��3��u��Zpn��z<����>[��Ml"Ϫ:��z��;�L�Q1{n�b�� ��M�ԥB��[����G���f��֪%<2�)�m���X���&*p=��ʤ_nZb(��D�П&"c$��/	�4�;�
��4yեׂ/^�/�]wI�vj�9�~�*��_Y+�۔��MߗSk�0w����$�ͼ{[JNy������8ݬ���E~z�)ӿ��ow٢o`)���ގhF؊�+����A�&��w��GC����T��&��+���޷�S�a��v �z��@�tئ�7�Z1z��,��|P�Wc�oc^^�j@�Vs*���ժx����`󇕳��}��fy?x�ɱ�~�_�a���NxHB��9���~J�.�U�]�<�n*T�=*���KM����wՌ��͕K��=�
�w�?G�Ze��`N��������)/��h�#[��C�Cͫ��3ݺrD��)�(f�<�L�ԷY�<Ì��~g��%�ʖ��V��NC=�m��:�^>��\�_�f}����E�t�'�  s�|52����m�+/�T�tv&�kxQp���qV�a��Y��I�+FOU�Fh�+OP|,oPOK�ק(n%��@�������7.����O���Ϋ�E�d^gH��ݸM��7~��.���Efe����%J��lo�J�7-�O
M�L�u�Co5��kH�H�\:�pPvmw8Ә{;;�k�����H���#��dW�:[�+�o�H�鳎�fS��0����0���l�\uņ�2K��:��*z���*���GDjU�Ŋ�ߋKǸF�řV[�5y����0@&E|w�j��ޥS/V�x
�WD^���Y�p��+3N�2��9�91.�5#x5�S���ړ;�+���( ���4M��S�c饈j�$:>�4-�ױ�[*�EH���Qu�q'��uGx�E�u:��v.�חe�Fڵo/��NgQd%H�S��e�sb4-�ã�K���qm����Mn�b��vJvc���L]��]�f�odu:����+5(�K�h�O0WK!k���4&<U�.ͷ[��XJ�jV-m�
�X�/r�;�'n��P93����O\�.��$*���������w�I�w��U��dP���f�8(���	�3y�0��������C-aYYKh�UJ���t�p�FU�R(����UZ��b��KJ�����YZ�D�+P(��-��B���Y�EqiW6T�-�TPDmiVJ�Qe�nDeJ�H�\8a��q�����J�����MQDU��ͱ���0v̡{�G����Y�#)I?�_UUU���?=���y�oQ�vk�ÜY�ŮLd�'��%�p�C*���]�F��ـ"�U�'0E�Hrl�z�K7Mu��o��p×�t��J�����v)�5��ƃ�dv�"Z'�*j��ܷ����z���U[�����9�����Mޭ����o�{b`�^�� ̫�'T�VMy%�"��xYzj��F�R���d�r4�[7ڡMQ��ZWވ�D�}��{(zL��� �(�Qku�Núb[����N�q?f�b��d�tZqҟ�}R��:���J�ڽjT�mB�x��Y���8� ���e%���r�ʀ����$T����;���G�q�-�M��G�.�~% �9���#{*#i+���=���^�������vNA΋͡�*"�t�x	.��[n&�*N�F#e;��BLϟ�_���`}�/�p|�Q�	,����ӹqm�.xJ��t-r�	�(t�:�3�1Uq�9h�kY���4��԰
���{*�I�s���\͋�w�o���1[�x2�r�+w!mHPU�#�h^a+�Zٖ��{xy������R�g�y�wϵE���.�#$=�@Uw��Y�E8���W,�t,H�uA7M�+��H! �WRvp�k�(���"G����n�W�Q_@y�:��OU�}ö`d�^�n�]�Q��&��;�����&�۾ѭ+8�a��jT�9��U��j[�X�i�k�)�vOj��/�T �B��$�W[�Mt�i�y!�|m�K�|\K���F���l�8�u#��+;\I�}�p9O�����r��Y�E�����Ym@Ә���N�w`�u�IY׾=�m]Jz�d�O��6�J��Tg-i5X��;�ګ��Q����~��n�w��+?V�u�����u��,��(��v��P�/iǪ��9��/rХ�MM;��j��7��{{�l�ʹom��!�Uz��c�>x��3ʐ8S��[.�:��bm�]���b.d��3T�ֶ�%�ævLg��D��ulJ��B�;����O��Ʈ��`�Y�L�6���A$z��tj�r���I�(o5аT�����~�/]Fs���>fI��^��թ��ȏq�C�/��x����q,��*y�d!B��Q4�}�a��xQ֌������4ei�#9��!��-�*�V��w��y&�|/�1����Y�|9	Us] ��5r3{*f����$R��3j����qŽ��y`Z�V�!3�]�3����YY�*�ڴ��	�]M��}j�{��Ǒ7���7�=�Ҡ!�FR'�/�B���SU�����A�Ҳ��o]E���]�3L,el_���|�e�㵠]k[YTEo�D��U��N�!lYJwJJ�t3 �>��#$�~ٰ
�B��$5�����lֳ�ʚ��'}�<��kUK�ȼ��6�֘���t�g�^�v�2���|�VZ�kb��p�`���*Y�9�spܮ	d��_up��!
�א� ��r�9�6hҥ$��ҹM����_���ވ��T�u��U1q&����]gТ��2mE���Kde*���w�G�߫��ʍ���#�W#f����`<'�&�x�_�4Q̰ "�~�	�BѨ�>Co�W�8<�SP�^	�=���J�.�4�9=6J8�{}�Ku`r�,�'fo4=z�zW�R��</��V�D?h���}JQ�Μ=6	��"H��e������v�j�qru��Ia��%�>��5ϛo�%�Q��p�X���P�k�F׎���w�:O��s���U��ِm(�g�j�6,B"�b۬(�*�E�ݶ+�"OVU��ގhF�34u�`.s��0��R�n���^`1� ᖺ����,���uvt�.(���uE��dcpoOw+���«�v������m�1�t��^�Fڐe��9>���y�T��z:!o�fu��o=P�Ó�{��	�����o_z"w6�]�������ͨ�4?V�Rch��x�,���PJe{��7��W
����@��f(�M�=۾y/\v:o��+�q����i�Λȸ͞	�������y���_���36�=J��MLj��r�����z%R.��m3p�_0��^�sN�Q��^��~Y�0܅����Uc������u���W�v�b��oj�2���tb����0�-�΄����n�Z�hٶ�A�n�k���{M�{��d����9>*�]�\��p�`���IL��"�30���Yjp�klΰؑ���H����C	�CT�|���v�zw�h��0N�����6:��(v>9Ԩ�����{\󳡴Ӓ�o-�=���М<��;ok]\B�� 5	�C��0m�6[��yzZ\�۫��W����)mf�G\�(���AJn�p#`�S$�ڐv�o���A�r]_ �j���Ц�Y'�ck U�5���:u&����w�9R��
�J���Y�`�2��Z�c<��{��3�G8��v��k���K�<�Y��<1���c`�u�::}��o>�٫�\9�l,v���%��q�
���7�ݍ�kO��e�@tM]ԍ8ՍW�Q�Bjƙu ��[-9w,��u���Ւ7G�,���ՕYƴ��!�ͺ����҉ff�0�)�C\���9��x�l'�i�|d���2u�'�8�7m�IV�f�,�����r)�K�[ cp�~g�]ښf�Dbĭ��	�pZ�[j��E�a��*`B�1��\g&p�[_s�3(���nS*)mY0�h��bًm0�\6W
�\P�E�Ë�q0�%m,V(�)�q�G�k9S,nn1[ŸF��X��U�.����X%��,iUe�1KDb5a�&1J� ��T�.LEi���X�5�e4DU0ҶU��K[��Am�QqI@E5���+[�S6Yi\5QZ�L1�0`"#�2�10�*��QE��"J����b��nY1�`*�0��jX6�E� �����=��q�K3��S�7N�Ø�_��z ��s��+@�w��p1��3�t��@n#����9mգȉ��>�/N�T7��t��OV���G�Gt0��R�����K)�yR�`sޖ�<|�
8r�ʖj�_����
����^��4��]c��QY]2�{^G�^/���Ǧ��:D"�z�r���f����.�tϾ�p�˖s�Rw�ƹv���d��I�뜦���ۦ�4�y�"��235A���<�����ʗ?G���vR�
����:%�%�7pȅD�q�]�� ��<��xV�h��3o���=��k�kbB�S��3a����큥=*W��b��۞��� �xZ5A��� �w���R��6#�5'u��$4B}�ޓۿ-����w��I�6��V�f2���I�7��Q�QK��P��:o�)��9�)�X.�GX�/74��*�T+�E�tZۗ���+=Śޛ}%j��0%%q�m�)s��������~ڦZU�g;��(��lfiO�y{/+�����^9z5�V=F�\��@���5��Pe�m�L߻.�^����N� Cو����4ơ�B���Z7�P+r(��W�ȉ\�7y�i|]]�9��Υ���dmUp�е�Vs��:k�I�PhE���ٽ�9���vz�� p�F���c�ᴗoA����=������x؜k,�l
�q\q}�:r�YT��Շt���D�����<f3��8k��
���.��l�4�:Cݐ��q�4�m��C����N��sr�l�������HO�iä�;�<�ڇ���j�=� IO����{�˽nJX�A��')�o���n	�I|#=.L�sȣ�Ar�gF��|PU��Yzgji_L����q�:`��[xp����t%��	��<6z��#�țw�{g��83��@�,�ќj!Q�MJ.���]j��R���Lc(Sz����u�2�cʚ�q�
�O���S���'��i.���gp��JV��п?t����UY�4���Q�	��	H�vN�ս~�~�,L[eˇ����j>��m�;�����n$��vR'wCŵ�Q{}�;�R+M��O�����%��(�WC�/X����S���s�
ɿ'1����a�vc����%�Y*b�?�_y_T�5Щ��,�F����W�rS'�|92FW�Bt#E����ß�"��&E�w�l2ߚl)�K�r�,E3�\^@=v"�[zwD���t�|��N-bn|&$�1�4S ��**YT'���Z������21�K�y��Ք�����Vk��!�C���7ҥ��>�oQU�Fnb�v�ru�ì�g�I���n�����|���K��JP�=:����q�0���||:z�Y'n�t.^i��+[|5b��R�� J�M�p}��z���|�(^����n0f���x�<�7�d�m{Ǝ��=wW�ͷ�i�}��kz�(R���:�^nBݭ����O$ȫ��4q���,�����Y �d��J�#�����e�N��[b.�K|��2/2{{��mz�X�{l���Ջ��,I6���Ar�}iM���ߒ*�m�mj����lQ�yOBc�8�ñ�+㒷A�5n������[���/sg�)a.�L��u�/X
y���w޻�����E��ʩz��J�XR0�~u��UkW�]�N��ĕ聴lM[��e���ɣBΦ}j�*!޻eӇ-�yXiճq�p�jq�����(�;C#{wqE"�]5�|�[>߼��]�-��R郦g�/�Y���*5���ph�r�G�ю^WiU��v����U�C0�JG�9Gq��bi�E�������I._'︿@�Ә���l�ldX�ء�7�Qݨ���{�� g�%=\�Ô��W����\�nm��.:�q�p��l.�v��̦>�yfw�֩3���m1���W%S��Ջ��i/
4��=�/yM�k+��p��iV�w�n�.e�CVHod�*F�z��$;.�����Ϲ
�
�KK[��۪��.��K'c��&�d�>��dwX�|e���	w��h���^kɛEŤ9)n|�Ax8M��!XEtM����Me����G��o��H�ޒ�w&������u)�/b1T��+;�p�o�
 �w>b�/ֺ��c�2(��p#JW�oL� V��σ����P��eiV9��K���ּ�n���uE��\���	t�i��Qp���Zyd�{p`�y��u��e%�	���gVV-�N�B���-�+���OWz��[�>��֔Cy|�x�Kݙ�s+,��[�;��]Sr�'��m��c� m��W9/jHU;�kU�6�Za��R��P(�g���+C\��o�T;�)�	:F�i:�ۧ�-�=XV6�f�x�P�(]�����HDnJ����!�v�V��O��O���ݳt�v_zEP�T��1��޸�\��Z�]��@��˅�,�׊iK���;�>>I=��}�l��Ŏ����B\�0���r��KF��(7��c��N�C�ݾ�\��1�!h�Q�r�G)��VƐ��{��˗{��fF
�.�e:�V�3���,�r|�Dpvܘ��R7ze�8�ɣ��۝]�������\�[�8/������cO5p[�Yjܫ��hU��D9s7��A��.B`W�s)ogp,�k��K:�&�W?�a2�C�Yr�>L~%& U�
o(x�ڑ�U/pC��P�2ތ=)��oÅ�4N�И�c�ۢw�m�e� �D!|��qU�$�۫�2�d��[�.��D�+i�a��m��{ꝝ�����nJT*� �*�m1�P��k0V�,�U8fՑQX#%el���EEE�X���:�ADŅTDTEE+Ukf��Ua��M	qkib��[Kj�*ŌQDT��(�*���ÅD�UAVV���F,qCN*�!2�0b�UWV\%`(��(J#n����TQA���J�Zʓ6���U`J�b�s�_=ys�|�׋��yv��S-+���)�W� cP9��L���ӽ϶%��i�T���=XŎ������x//O1��F=�H���L4g�t`�ST*j:�o*k�����Ot�֝����mܻ+<��{�ܓ��#[v�S���^^ث�V��5,�~�NmkOGy�{2o��h�z�+��X[�f4�>O��gZ���̑ڃAM5��>>���!�MzT}��ǭ�WaY�+
�SF��az^���A���Y� ib��UԜt��,��f�ڹ�B�,�co�h�J�=���W]m�{V�7	}��bԖM̜E=��8~�Ilr}"��ҵ�c�����]Ʈ>�S��w��f��zK< ��f0/.�(D�	w�xm��د6�Uej���	�Ƕժ��&vX���\����j]o�*̃�t֐D�fzݺ���o9�����X�-�r���1�gx�����Ou'-P�3�d��驲���l�֓��V����)> =�RL0�f�.U�'��Ŗs���q�{mb�f.�W���ql��I��/�9\����<�iOɘqn�֔�\�s
\22�&��|K��C"�Aʤ�G�Z`&^U\�;ڋ'V`���䜌����dS��mv�����w*k�YqDEu>r�L��ۃ�qh��l���7�D����qC[�O*�ݘ�N�bD�&J�Ѕ����Iޑ�V`as4� �f�e� ���3סg$�
�՗�=���3vg�#��Ey�]�T�Q)�&�t�=�b�^l��M�RA�lh���}�.�]k��r��7]؎Y�&���x��N��ڋ�;Z�-o1tR��Y�u<t��c<�<
M�W�|9s��{�Nغ��c	�]wW��:5�����5(N��S�
�+~���#e�e�Q�%��{]�k�eJR�1�^ԫ��d��R=�@l�]�^�Z��6r:۶R֬��W뺩��4���f��j��ӽ�~H�M��~�"�Xz��]D�Yo�鶯FI����RܽDSu
`�;���o��m����bRs�4�%���B{2��r	���F��nw��^��T#6�oH�D5�����R�=��ΖY�gW�F�Pל$�]1�:62v�I�C�n@Ac�<d�u0���D����(9fɻT��15�W)�[���\��2���S��d�uwyn�D��X`��OBaKx��p�.l芗����'8�˻���{Q�� U���)��=QDZ�ؽ��a��\x�L����x���(��k��q9t�U�P��N�t�éi��ڋo���F^v�t���=�IKF�|��*�!ҏ7~��tN(��A��3R�FH����&�j�#�^�4��1i�w��Ԫ��:�PM��^0NFGV�Z�p�Kٌ��/\�P���i��f�,{N�B���Z�q����I�+�aNs��c���]E)�Hp�"O#��:������Q�/k�^�)�tm�(B9�9C��U�Rr�d�o��L��-,Cպ��bq��|U��L9�nMg�^�����7�_��I/��ڢH�=|vxV^@BE�"���ݛ!S��lʓ1"˻LV�3ɰ�C`ٺME�I��6��m����/S�ʪ���=�#s}=�n	�i����<;}����e�@�J�iq-�g�UE�]%8�B�{�f<Vo�=��j��Ԁq�^�Ks\:���]W�.n[�dxu�+��W6j��o/r�k	��j�ڴ0��KP}�$�k�0>|y<��^���l�̣��p��S	����{��_����]�kB=\�s��t;��1 W�[17oI�Ģ`4{ڀ���0��Y^�~���7{�/�W�n�g:rxe�y���������jXU:�*Vw�v�or�mq�J�����<n��z�U�N����ZRly��nm!u�o�K�֙w�A�h=P.x�>���>��4�0Vy�VL�Ǳ�G�kJ]Խ�Q�8y�+T�nn�W�P�4��1�CN��{�~�g}��1�4thJdv���-��a>�G}����ٲC4P2���kmG7!N{ۊ����S٪f&�5(��]B��xѮ0gA�N��\��w����e�y'�W��(��n�ւ��ۃ�扱*N*�s����n���K�8���@#��E�(M��˗���ն��+��^!v�=�,��yhF���D^E����m��ڍh��OV���k��r��Ļ�:N��8���K�BS�B�[
�Kg&��(I;z��hn��2Qyۘ�<����1���$�wY0T�ݐ�� ��U7�%��u��˚WH^�P9)�J������[��c�J�^\�K�T'.3d)��Q�:9�n\�7'�Y�S�P�7.e;�F�R��7{#�a�̙PEyu��[y�*�ި;�����!Q}S�;Y�#n�fd:Uv��i- ��jn�u�f1F�����5�U�= ����bV��*�R�&,p��r[W��*�D��Ki�G�׷ǰ�l��wh��1�H���e�{�_��R�������YI��h*���˃lj��,��j�B���E�#��+,k[�-`�7�Q��VzY���vC�xmg:5�"�����z��.m��,_vdD#�M/,S��ܰWe��~]��{�8���9"ø�$�R���v�����{z��h���w���ԃ���X
�ق�<���5���YO��O"��dG���3��o%�4��f��2����q!m��R��ȒHS��:vC�E�y�KX�����Œ�T�Z
��"|�2o��w�D<�mmc�*�ADE����b���-�"1t�rR¸������J�Z�h�h��"(*
9�P�3���1����)Z"R����ͫ.Z �.����D#�
�A��j(1�������Q**Ȣ��L2*Ẳ��X�5Et��DuC8mQ&qLR��Ҳ,Q��D�5�c#YQdPB$CLW���p��R���B�J=�ݘR�&a��ؠ��w@g�~�����!������÷%��i�yŖN蹵���J9�X�����z�u�H읕��)����])�O��/rک�}���sS�\oQ�V}~�?p���gz�((���Vz���)Of��s�2��Gzc��w1�Q�>!�_@�'>-��_����H��9�����g/�<���{_ag
R;�'u��MGK��#u(݌l��i��,�3L���b��F�+0�o���8}i���m]��g��X=Ex (ǫ��[0���eqR8h�;Ńyծ�d��gs"��е��Zv2��o�� ��;ɿ@�Z���m�g���W%�Q�9�1a}c+����r=m�#�t�tuj�ɉ����|��g��q�!�w:�eC����j��
Z���!��IP�@���T�}2%w�ubH0#��ZoG�fU�ˠ0�n[hJ�o�i�[SN����P�Sb{n@;���9���nU��W��� eBع��C��@��b88J����O]2�Е^�d���rt�]��0��n�^��ş!i6����x���a�9ot��}#7�*��}�nWE4;�;�uY(!���0P쯷��\�xs~K�:�r��<>޺�y4}閂�py�spЋ��\�Sr"bouGi=��_R�t�����y�/D�L<��٫���j��\�-�!#6\O*�L���I���	=�mc�喬�b���=����I���O!�I��چ�
VO!7x��z
�g+y�{f4)��޿W��������&�A����&S��铨U� �>������"[�
��7^IynF:>}JҚ9��E�$���Q>��WU���zv���8:i�w�~F��V����ɡ�5��p����T�tć]�wN�W%��(&���������l$f]x��!d�|���)��#�z׵��;���x�-zޑM[��2�¡���:��!���x�6�u���(,��T7�Ņ�n����w�٭:�S|w�~�<��7Bv0Ӟ��^R�]������&������mJ�S5]_%:T��~*��HTo�U���M���
n��>�\���h��^����̅;�TIO���o���=|��G݇y�ٛ�ǉwzԵ"�x�m�gv ��xX(�*���R�`��%r����S�ޮ�=������S�_���i~]�g6�mT5����&��#�e���%�'�|�>@���J�
��{�$���ŵ=�VɎ+��
�[����a�Er}ʱ���7���;��龹*�:�i��u6���t���"�%��d�; �h^X���AV�t'`A��.�Ʒ|����$�P�}�nX^���~��E<�x�\(>g^�\j"l���p�����daAD���jZ��c�����!�p_~�S��ɺ͆R�8fGhf�i`(<��YG���0�����X�O�ܑ�>q(�4Ow)���3Ǫ�f��|ol�7�4�:���GfS��k�ℕ	W�~|`�o����w�ܯ,�Y�9"���]���q�Ћ�SG���x�.\�V�z����"ފ5����C�q�,���`r�3�z��{���7ˍ����z�MM�&urɟ��/]>�q��K�>-Q�)��6�3�z�y�W�y�(���GATf�`H�|��M��y�1�_<?!�H�Mq5b�`���-��\}�|`��3^*
�j�ڬtRw{t����*4�kAl.>
�G�u毎7=�s����;x�A�g��۶�ø��ֽ �PU:vP��΄��^k�����|�x��x��`�/����7������%E���Q@n<��@čV�1�;)��u2����s�G���AH��hL���re�p�����q�$�~ D;4�"Ј|�6zCX�m�l��!1�-��#�j�X�b"�W��"5F��|�}��{�0`��f�4���p��cY����}����u�/�\"�]�LF��>I�;�>[Z�h�+Dư|�Q�������PVc�=���ӳz!h�b4|�a��|C����X�Oڢ�2����5b�^�ʐ���������Κ8)i�゗�
��Ŵ������5B�ۗǮ]�w�wvk�v����;�νt����g�f��`f�5o�b����rb׫�A,�d��z�Ӄ��^��
%�� �A��rM��Fe^K�.�:4�|K�n@�2����g�V�|�P��A��.�}�{H�>�t�u=��c��x�)���7��������\(!U�,�Ѻ?p�Pc&:s�6�jH�9��^z�t����pTJ���ՠVq�CY�4i�K�!��n�u�{��$"���^�Æ��\B��G�cN�٩0���"#�ώ��@!��a��f��͵���Z�ѼtX��!U�9xE��v*
�.�Y���f��x�
b
�Q�s�K��}�ưz�3g���˧o�����������j~jV�*��� ?��d���_�%�I	 	��vм�P�
��4�w��`Όw�:ܰ?�BBa d��*<�ChX{�vP���L�B��C�������l��O����ֿ���d��1ߞ��\M�Z�28?e�Nߧx��~�7���}�H��>zjs\3� � ��{�;�����(h��	$ '��'BI 	�~��`����r~�~? ��I�d������!����F����@����B@w���7�����T�&9�D?G�L!���/��MH�O�]� ��8V7"�����롐�X�X�	 ��z��k��f����0 $!������XN��u��������5'ס�\��$$ '��6��q��'�>��1�?�&!���Y�_��䇇��d���F��~��!O���������	 ?Lg��O�l>���?�~��e4b���4��P(l��~�����~3�C���������wԟ���~_�����rB@}��A����P�����p?�	��""Ԅ0��$$ '��I�I���I�O� k���!��æ�HO���o�Đ76}�F1�L
w��'��ɫ&��~i����䉭V�����71&�O����>5����#P$���~��������$$ &�~������@�R���P�����x~����&O�����6?����~P?��~Ϗ���?�����3��$$ '�~�_o�!�������B@~y?������I?����Y�}I��������2H�O�?�LA�0��������9�7��x�������7;�}ƾ��&����O��������q�>�0�~�J�g����Tn�>�����P��h��I ?�O�c������������I ?>���l3����i6��,�k�����B)'��P=���6�.�p� �� �