BZh91AY&SY�����_�@q����� ����bR��            ��%B�"��H�R� �J�I@E��R"��H��P�	)T�JR�ET( E
*A��V�h {h����RDum*��%
�!$�UIT*	��AIEP"J�I%*��	4�lJ)IUUU F�l��J�RS `�*����D*�OyE��RACrF�A@z4H �QJAB�E"�H�� �V��
��
��P�����Ғ�4P<��4jSR���R��j��cB��b�r��Z�\��m��q��J6�-����\.�[`Tȶ6ԉ�y�)I! ���U$��=Ҁ��JR�$���S�4��1���B�%AަԕI%w�C�ARg�s�*�Rq�z=%*R�w�缩UE*N��"�PU�����**���5� �QB�@���(��{�T�AQ�/=ꂒ���W�xPT�8{�=R��y^8�U%J��<�J�*��O=�R�R�=Oy�y�y^w�R�TG=��=RT*I��J��E*�!R�BﾕV�7_	A*%���ި���v�/��	Sz�{�R�J��y�JT�Q;��z%;�y��*�Q^����!U'�^�Ϫ�>��d㯜�+�T��P�D*�$�R�J��*� ���J��B��Ȕ�"_/k�k��R�u{�PT�ަ꒪T���R�IS�Ox=J�h��Oy�R�J��R�zP�J��ÝJU*��z��)HET��Ux��� ���aJU)N�7JQ)JW:���EB�N�Ψ**�[�J��U��:��kTJ�	R���IB�3���ӶIU�MԔ�UUn���UUAE
���G��/�ﾾ�Ҫ�\�^�i�p(��wU(���g  wU�U*��Q�T�:��(p��WA���
u wT'f�D���RT�|��d �G��5M�;��hj�-p����(���� ӷG4 ��
 �+:P7v
�};� �
�(�%T)
RH%E  ���(�;�b��-�p��wH Ծ�����΀QKqn�A��(
�ԝ�@�@�� %D�*T*�)N��H�� �}��bn�UAد���� 
���M��mJ]�=� *�ޖ�:j�ΌJ�c�:4��  B�P� �  �<	�T�(     �4bJRT�!��`	�� <RT��L  i� 5O��*T 4�  � $�IH�*�L� &��	��&L�j��$�d�AM��O$4���	��������&���%�@�������%�ӡ�]��{����^���C�[�mη�QE�����DAS�
������QEW�@���C��_��ݪ�"�+�,�I?�TQ_T�QQ@��>�����dIJ��p��I¦.��A�(a�L N0�p��I´�9�"N0�p��¦�(L*p�8T�'
�HD�Q��S7
�E�)8S<�S3� �*�p�S
<'
�@�P��C�f8D�(a�S�L \(�p��K�-)�.0�8T��B�'
�@�T�$�S�
A�+�xNaG�	¦.p�8P�%¦g	
@�T�$�S�
8@�*a�S��"\*ap���L s��
�D�T��W
8@�*a�p���\ �(�p��K�$�[J�D�T�$�S7
�A�.!�C�C�
8A�+8\"s� Np�p��	.0�!8P�®g
F�S��L#�a^g
E�P��C�
D�*`D�T��S7
8D�*N�G��7
�D�*a8A�xA�*a�S��#�&8A�(��@�,�C�\(ap�.0�8P�9Ô���S�L \(ap��K�$#8T�¦'
�@�P��Ss�-)0��$�S�
�D�(a�Sa�N.0�8T�%¦'8P�8T�$�G�
�D�(a��p��n0�8W�
Fp��n��	J��L#8W�
�p��K�p��P��L"N0��(��(3�E0� �*�� g
���@p��PI�9�A@�(��n���B�D�(�¨8Ep��A�QG(����TnU�3�p��8ERp��VV�A\ 8QG
\*)�g
 � K�U0��Ey 8D�EL �8P"�*��A��(#�T.T� ��0�%�ARp��p�p���(��n�"3�a�p��D �p���*8S�Pp���E"#p�.T�(��TnA�3�Q) 0�0���*��PnT�3�@p�ª�@Y¨ZTG*\(�U'
 � �@p��T �"p��@'
��B�UC"��(\*iD��D"�\(
a EY�TW(�Qp��&'
6�Q�*�
(�Y��Q@� .P8A �T � ��@C�7
ZP����
��XI�EV�Q��p�-¢�DRp�4�)Pp�-�*��nU�*�� p�� ª�*(a �PC��Bp���
EFp�!�Dn0� ��@C
�(�a Bp��E�
�0��*�A� �
��¡�®g
A�HQ��S7
g
�E�T� �C��*a�L�J@���K� N0�p��g
F�P�$�C
�@�(a�C���+�p��g
8@�W��"\(ap���aS�"\(ap��9
� N0�p�'
�@�P��S%g
�@�W	8P���K�9Ï8T�¸D�(a�S3�"p�0��$�S7
8D�*a�S-(��G�"\(ap����
< \*ap���L"N�)�Np��	n"N�p��*ap��[�L"����"Np�p��np�8P0�\*C�+�p�p��¦.0�0�p��In"N҆.��S�(a!p��%�
��p��������C�@�J�f��R��<D$��DUܡ(���!7�iE�����:�fD�8�d�-9/MKiӃZ�
�u�������Bu��^-�O�����+�Y2�����Pf��dU�J�RDq��<0���-�w��j�e����u�d��I�5opQb���&������n�+GMm'�u	�i�Z.���MU�kL�ًlE����p��Kn�B2��x���h;�V�����j�����yJcn!b��ے��L-�F�6ێ��=���TF��DM�ML�� 9 (��r���Z^ �v+��ʣ����YKl�� 5Ǝ����qu�J��r��|�C���0��3�l��d�a�G:�A�爽gCb�!3����V�[.�A�o/E#F���Svj��PS�k$���rZ�Ӧ�W��ų�aݸ(�<�>	����an�]eZ�^��6� ��C��Ax+#�@�]G���p���ImÕ݋C33e#�-�vS�5M�v͠Em	J*v����c8�P�LzZ��F�wu`�Y�`��*�RL*���N�U�nh!�6�goR�m� �:�n��.��t=C{.A
Ӛ$z���ꏋٝn\����e� ӣ,޽���ODE-����x��*��lO[���
�n�h�����hZu휗s%n-�l6Q��[b�u��Ef��H�.ڢ^���ٺ��9�2^Ag0֋n]fD�$��yw��j��sAͅ,��,�2��6Q�$���i��YX�eid�r�X9If`A��2��:�Yh�4��n�E�L�rF�5�n�ҏf����Xz3�9VڧHL���(�#7C44�&,������U��1�����L�L�opͤ<�Yd]9v�)���m��d�)�=ŁA�n���:̨�qc��ۈ�ܘ�YW"���L�
M>+7u�)�r�rɷ3(tcD�5�N�әY��̸F�pM�K^�䕹W�f�ZS�b3e]ѣh�R�Y%�94
�tޚPۧH��v�3K��{���4�r P�WK4��@�6�J���[2DP�ՂB6�GF�B�.�m.7��5�E3z�nU�w�G$�CP�[9�mha+	�V&�3N��8�V�+�ma��>ve�Mݺ��ӻh�"P�hEVI \���7�D����2ʙkvMWW6��y{������̬V�c�I�ݭ�T�iP�����������I#�;lS^n�B�;ڲ�����F���M�X)�U�����4r�PP���kP�y�XS�ZpiX�V���N�W���9Ϧ[�8�F���lچ�Sh��:�΍x�(��v*�8Ԉ
QZ�,���V� 7j45��,k���RGZʻnYX�J����l#�*:-	��h��a]�Hem���ݢ���75�w��`��n���l�;ʕf#d�Xe�����uÁ�Eb�V�)�%��^��.��q�XN��}2����8��o�˭@��T����d��t6�<!��d����䕢�VT���Oq�ꆜLdk���f5��B��x馛��kL����SEW�6Ii3���&ұ�=aY$���M�<7��M�Q�e�EР�1
�,Q����m�i��ʏo%߁k@ZےmL�tm��
d
h�ΠY݇;[�^+��5�`х�t�O��Ih�A�����xoA�Xd�u0���{f�V$�2<zh�F���r��@7�a!�3n�1�Rݷ��u�v�hXt�U3W��Ԑ�"�i4N�n�Qe �ٷ�r�0��;��i���#j��x%�;��7tm���2�Y[P�<I�E�3ZФ���]Y�d��YfWohD#G��Է2����̼݂n�-3�����oE%�,�u�6�p�N�n^�9��ʤ�[E�z)̇+>���'.U�,���PnU �P��j�<^lݻ짼��*�֕��xa�v�;����Jh�2��eS!�O�l���ģ���#Vݧ��n�7x�h	@t�l=n]
��u3[�0YƢҐ�3x��ŇXyK*�w,�f���M^�J��;���Shƥ����44�;V)Z��(n�鼴�n��orWJYˣ#yZ�y��ɷ�Ai�eı\[�4�8�5vN�un2� ����炊7��� �"w���A�#&��6���Y4n6�񴵤F]1rU�I�
��V��tt7�mL�O*1A�Ge�O,��bS���b�]�l%̲���-ֹ.;�C7V=ݻ�QZШ��q$�L��ef*TVܦ�\,�we�	]X�L���+0[gN���06�Ǖ��6�	������X���oD��5���i2�!�Sq���d�(�e�T�)�f;X��Z�ZP�6����ۄb�#/t=�3]�ۆ��������&H��R��aBoiK����z�p��p�Kzn�p�x$��m'��[N�����t�7��`�>�Z�F����CF�(���ݎ�Â�,���Eq*̬͢���"���6иCY
z���V�!eCZ.�8�{���.�KklSx���nj㺙���wt�Z8��Q��.%b���ݔ���Wa��u����O$�E��ؗdkx.e֚F�ɴ�Z�Tm9Fj!�iS�RxooY���SX�m[b��t�BF�Z����bl��E�����eIK᮰�ub�����X�M_#`Tl6�6��`ű	
p�5�
�	٠br�[���v�wY`�Ĩ���ԭ�u[�/*T�l�e6(犁]hd����&���^]��т�f<��lq4��eBkRթ�V޺ �P�m�SڃHx]]�hAB�4�7�R�wf��V�fe:�e��k%$a*Q|j��~��2*��$ᛳ�[�"�)W<����&�rC�U�ud��x�1��aUʉ�PO�B米�rf�Z��/p++6�1F�Q�]�4���]%2-��=^{�**��u�S�.�-.<-Q+l��]5z�8Kyx7�Hf�j��mf��[F��H�*����-�2��qK�k�
�'mL�2��!rRMÇF��O2tn�D>$(��0M����LTtR�Rqk�i�n��ڛxej�f�nE2g�vu^�;�!�����T���^�L��,�˦��F���S����oJ���8�Māfx�q�Ɋ�)3ū>ћ�9�5�iX�<9xN#�K��Ӂc��6���֔q�łQ��l̺.�yC2�F��0Ri��vu�07�榐�R��Ĭ�� ݑC鵕5�!�]���T�A�[1�cwi���K�:Ln�nd�o^ݳJÖ��s�S�Ƹ�lX+0��o�`�MTr|C:��ϔ%X��$�rִ����f�[�nS%�@��B��K��n�HAv�;R�{��b(޺j"0PX�W�iݪGhH���a��HY�W��8ln����ִ5��J��
-��)�Cq't���1�朐�U&�9�9xjP H����NaG��,�����[�]l�����V��j��3Tn�Ui`_b��%[e�`
+��P��++���a 	�k4;v2܅���Ǯ�Y�ۨlKj�͐��f�jCِ�gl��J�M�;�3�aN�N���`-��H�j�%��NRK�ɵt�c���^�<Mբ�\�-V��q�n�}DmM�$��0Ym������v���b��Z�ͩY0�Z��h��"�e�(�r
Y%���5ZP.R$@�)�å9�.��=x�Bj�z�ݣD<.��/Y�S8�Xɮ�ˎ��yS"ˇH�@�"��Z�7���3b����*�z�dJ<�ViC��$l��`��/�2�#�TV� �X��	�^���˩��f�ve&���ZSv����mV�*]���ui��4�ٳGim��W��&��S*�-�ʙA�3:B���t)V'Y� 	�츦���엘�j��[u���	y�M@0��U�r6�db��;�j���4�s7 ��\�J�0N��Rm`l��-Yl�2�(R'w�V	(?���#��X-�.���]"�U�YV˽u��yW5�0S U�>���К3(b��VZ�i8nBh��-ˊ�0�C^��'o��jS̬��:����m@� �IM�n�h�U��`��\�{���2С6K�Sh **(���j���WI� �"��Mƚ�x�&��ֲ2�5���u��)2Z�d:����z+�,��e*�v�u�(�4	�4K�*9��<Ӎj��ǰ��Ţ\"�o
�vM
�C�K43m�-�!���K�au>��^����
���iV
��[z�\3�xxuK��[���]���L�G6�+�3Sˈ�9h�f��7&(֙eL�b��)d�-�^�Vi�l��t'gH;Y����El����`+X)�h���`��0��eˈA�Q���0��#+hV9�!$5�j51�13����ɸ͖���7�rn���Vhɍ�Ź�T�%,l���,$MV�{�Z�+P��f���q���)y貀�M��B!@T���V����v2M�+�f�CX�c�(ժ�R���fF��A�6���C�wQұ�֌y�[ݥ�6��5�Ϯ��b���u�ӵ$�z4-����Ѝ7A��X��.�ef�[���wd�v�5�dB� ���1�����P!<wq�a*��&��`^�1=�B�iH��7b`�e�[zh��7i�ʹ�5c����%�(�+h�x�W���6�,�K������T�ųCH��PX�pm�-ǞcAm�Kt�"�6A�1�I:��j�i�J�dj�2�w��:�5]�6��y 7KM�ҥkDeg�U84���#�(M��Z%l���T�9v��N�a4+SB;�Shf^� �,�����I}�*����J^��᠎��aY�L�e�EnaQ�Һhw*��J�65�s2�@��xj�n:P9Gwc�g0�WC���oq�+6�qS61ѳ�An��ᬠ�v�%b�n[��Q�Ꭵ��ڗ�.��5�yn�9Z�$�l�*Y��A�엫r%����mQҲ��=z���]�XvBE�N�5�p�ƥ�)�7��tTt^���/�-~�+JaP���g�ww󐪒:[�9�Ee��2��T0��ɗ`A8aUv�\Tk) /�pт�ś�*�	���x�Ϊ�ٗ���rL�1{0l+\:):7��F�6,������{ZX����� :�������J��mŠV|��
��e^�8�cli�V�bv!�P�tۂ��jS/"�f��I�A,jC� �D���N򣕲
� B����ܵ�F3nmb�YXvԎ��I�e,��v��vKQ�Z[��6��x��hIf=t��h[����t7 ��C(�y�3�\�{�{;�z�qf컑�M1w,�A:Ś�QUf���]��V�t�N�4NFN�3엂�qk�o�Yx�TZUY����� �0%�dt��0x-+r*�8��
�F�P�,�T*�RZkC�����,�NSx���U�
F�*^8��ȍmJRW�N�e$[��.n�l͌�
l�Z!���Kr��v�f֬�$��*�Pu{t��Bjr1fó��9e$Ȳ+��ځ*�T-B�Z
Xc*��J��F� u�Nb���!�vٛZ��ED�T�{i�
^[(b�Z!jkx�S�� Ū=.�F�f�+lU����jV��MjݺT���>Ȫ�՚�tuɵ��<R��咬���y���}e�* nV��a��ml+Z,X�֬7P�iV��N0�66d���v�4�nXLZ�ҎG�R�u��s~�k+,k)��4TZ+Z��ڲ��V�����%@� ��Q�e��ti�kV���]e]��{/d6�������e�1��SiE�Z�q�{�P�bQQ�wx�614�7���ù1�d4�s�ۙ�f\ܛ�n���T-�{{��&aj��J��+Ҳ1S���w���#�SNGJ%A]
���h�P���b���0������2ϴk4�Ǻ ��ϴfoS���fC�.��>������/H�Hp"��-��όa����@`Sm��t�/��E��k�{,�lh�)�!Hg/a�RY-,��NP#w�4�Rh��dp���L�0,�(�렗u[[����ޡ���]�?]�W�����|i�ѠY.���p7��H��E2�nJ��(G,օ�CIA�qh�y���5b$65w���@��[t2�Cfqe����,�Ց��ʁ���I#@x��8��3�v݀(�@��B�B ���T0VE�p{����:ɰ*�VR� Yi�Y�.�w�딸�B�p�b�<8[9g��@ E@�"Hoj	˫DkQX��6�PV����^�t+�	&�#l�	8a��Y%�9Z���+4�f�-����wr^Q�o)3A�/@�-]'p`\���uT��Þ�W��Y[:o;4���%��C[s�:�s#y1ؿ��ܯ���0��ѠlӺY���5RF��b��6��>,��tqa)Ձ���P+��V
%+H{K;R�]dS�}0�PP�`'GF3Lz��|���X���x�8��m�4 �6���"l��в�z���Z(�#�*ZD�$`m���!a
ѷ��;�˪B� Wu0X�5��8�zk�u���ެ���
���7�����Dh�+��}Z��B�v�S* 6neɔʥ�Ut�@R̒=��6\p!�o�
"]�P�$U��5i�Va�<�m�EJ���$	w_Af�4I�W<k� ��ZN�`�F#c�$�V,�� �7wY7D]g�������oG��@����?��@���ݝ��{=�ˌ����x�>���:9-�}0C@�gE��N{;��jY�-�bq��[W��lJ�O�,k�<�w���p�h�h�Fzj=�:�Q���X3Zo��w#����7	�N ��JF�2�����g����4��;)�C�.�^"�
�σvVvv��%���Y���saypդ���1=�Q�9�z�I7�|��3w}���yu�D�i�%Ho�����	�xLI��wl�o��f;����y�K=���u(s{�@��N�Tp\�b\Wo�1Lt�4�_j㥝��k�ݎة�+jf���i�0^��.���|q�J}�K�͊]\�,mc1\�:`�z�.8ud�w���ה��*|uش��+;#U2����#�{-��6k
[�)L�J�{-ɄVgY<��̥"�M<�5|o����Td*=�`�W}���|�K�n��5,�\ySq'τJ#Y�hB�a�M���K�
�w��֜��P�˫�Khvëv���g'B�5�&��!�6VФ�ݘ7��W�h5�=F���=�˸7��]V^��Щ���I���t�u��7�/AwϪa���v�H��'�Z:�f�E�mG4�x��Ɠ������9u����L�ߕ %�u���ª)CK6�4�s��j�#���R��6/zrv1	ǝ�R9X-������`��x7�����lg���ö�-*�n�>9�B��gkݫꮪÝ��ba��kP�k5P��B?DKG�5w5rD�]�����#��9���e��Y�Ŵyp�!�����n���<	����X��롸+�(.�ܬs@�y�ͭܩ�>{��T����s��i:����k�a�kn�9��Luy�r*Th������`;���Е�6�[im�����,wh��uz"D5�(�*�go��s����R�͙�T�Z��/.����7�����ڂ���e\��6�$Ѵ'	��]zNmƋ��Ae��ͫwI�8�X$�,�q������]jjD��܁Kbj�N]� ���R�O�Y(��6{l�S���������
�>VG	�p�An�D܇ۄ&2��"�>�{��B��tB��<k��>�Q��U�*�Q�;ޗд��v�+
x%h�sIia��K��s0��V<*��n*ᝰY�^4Q~�+�٥}"y����������B��9p��+hh���%�7��Ev�r�e���a�o�we�]]�VF�r�����+2f�C���

�JM��gIv�e��6Vd�>ѣ�N������K��u.�J�t��d�5��@o(9A�)m��^�M �յ�1a̮���*���;��E�D�W��t���C��|B�7���쐊�X�CB��=��{�E�/-�{wut���2������;+�T�rN�É�+��v�m[n��sq�UsWŎ;����9��=�vGp�;�w���X����Ϩ�.��3�Ǝݸ����D�C7�3��A������T�t���z	��n���P�w>���إ-��e2�fTLYP��4W��l�7�澪p�0��;�.E1�K�Y�Ms�����f��%����M��^�}�����tD����dgn�[��r�0�}���B�ϗ������&���w�|ia��U�}��X��r�g2�R^����N�ݤ/9g8A�J��YG����v�ͦ4�4��Qd-�`�|;0gV�Ʃ���-w3W�@�jӻ��]�mq6�+Qk���{�Pi���nM:�S;���j�g����"rG������99owoP�y{����>�3T�0ni�$���y�';mQ�MV����� �4��e�o�x�U��,a~2J�3q!܃�czm����kGQ�j$�4k�>�cb6�lQj��
�t\J|��K�"=�jB��j;OB��0�O�9�xt�&e]����p�"��*�k��._
;�7Ux躈�Ģ�e�]_+5�u�8�2�xa���.�=� ��aoB���M��)D�W��q1��^�o	�
8�m��Kʷ���f�q�ɐ���1��Z�h�SO���}��`�+�i˅a�ua[�׽�P���1ѼQ�W�W9e�)�j�����<���r*�=�Z��[m7YXo^\MԾ㍚����j�r�1T;���]���$�]�l���S�:w��Hh����{���2�d���׼Ď�,
��h-Y-��W��)�/'Uݏ�f۩ۺ������(Z��G�����o��#ɟ^bh�<76�.,�ݎ�p�JYQ�is5g��3~��Nt2b�����io K�8�p�]M�8�^�O�e��Z�jdh"W6���S)�sz����.xܻ�u����q_����#��yM�gu8�n���;sZ��N�L����Ν�L[Z��!������1s�j�MmB*�q1̴�"�37�����[Pԙؑ�[j��Чj%/���<��MRd,�y��;�v6�g��K��q�e�z�f�i�����׊����yP�����[�ْ�����z���2V�>2�T
�ʷ[�u�v�;74�֫�'H�q�β�:UwX�3o}�*�sP>5��q����-kWS���ͩ��a�˳������G��q�����t;`oy*ݚ,N0�g\u��fݣ&���6�ro ���؅Σ���]t��8��Z��Ms� �5SV��uΆk�NnK����'�]Wh�GSɃWlU|�0��n:.۸.�N��QV�T�]��u]��ծ�*B���]>�ζ�h�	0��'PIӕܳ��΍�bc�yI^b���:)�*���[Y&�s�m���'��8qKS��9�*l��D�_^kY�tGv�J�H�[��[C�����nv�
w\�P�+�̮��(]yT>x	����օ]��o���&>|9^6�̽5}ٻ8J�c��������(Uܣ�e�}d0K1�b�bjJͼ&<��Op0������-'�KCB�W[�Oԡ�l�շ�otuXY�+8 #0b9�t��#/���y������v(r�ۑ�tH�˳\�7ْKO��l�׵d^�M��fؐ�U�2��*e��H�@]�]�B[���"�¬�k�h�Kq�x����f��m����1��5:�yMk�.��{R��6u.ؖ� 6�M��ru�MZ��I�����e��ˋuh�E�A�҈.�4��\,��K���\��5�������| 9J�u3�i��9P�C���7�9����^u�op>J[o�vً��WD�2�78��np��۽�r��3��r�9p�62#ki�A����ZE�zn8+q�e^�v��]pm��٩�*{�+��I�h�gp�3gIl_v:2�#�xt}{t�]�q򧅌.74XI�&N�]�XOW��S�2N��۫]u7��m��x�aP���)��ȃgmŎ�32�V�0�彛��\;bv���Ieq��Pؔ�4�k�V�c�I��h��&�h����to��)d]wX��O�ΦTs�_E�.[��ZJ�N��v���XaOp�U�����lip��b�##S�s��`��s\�,tч�"��N�owP���T&�v8���uϲ��
d�	ӝY��fn�\��^�)E�<�&w5�9ǐ�G�mZ��/t�,Qe�̶�(���tN��;]1�%3�|�<�3��=ֳ�����V�o*����]�h�ݲ^v�,�`����a�l���Jb��'�;���E�\3U��J���z*�d�*����OE�5	��@g��DS��WJk6#��<���SQ0�\:=�cT��}qܷ��"�c�1��:ou�-��,좏C�ۏem�J4�"�׷��<�m�A;�-w�Z���*P�8�z��(��e���!%�uˍh�{*��D#u��OS;F�Cm>�Cx���͌�23�*ƭ�RV��o�_Q�
7��-�w��DN�IX�o�B�|�B���
M�~ ���#5� �R���:�T�&�]�mou=�p�x���)�X��\�*��_RG1q靅f5Ȯ�o{6���Uo[u�8�j���Tv���;���R�}�ҝ�Tl�.��1S�z��Z�_+�.]��b�7f��Q�]�v�ór�8�HF�:2�#��HJ�6�j�T;�V���&;y#O�l�dU��*]1�=�R�b�7p�^w�<
����Ճg�mTz� 3�#�Ԓh��Od}ѡzMm#�gd�[�@��؁n��.{�کw݉�ݦ�Jd'���T\-����j��u\����Ɖu��:ș&b���e��8����8f��\ʹ)˾;[�b��:��C�Ń�ճ]L�([��n�c:87ێmݚY,� �ٴ�}Rg8�n�l¨M�ɴ��&�,�v�4k���R�	�!ՙ����j;�m�%���;��*��XO3��
��hcΧ)u�bỦ��L��A����&�;���w��鷈LӍ:J��x��P��6v�:n^�=�a����J1S�*k]Gy2��5�2�F�Չ�ʳC����&c�Nft�W���ge��ٹ�%��=Qݲ�L�NNƥ�Z��e^���ɥ��ֹ���V�/z��ʻX>�ɳ`�we%��&�UÞi�����@�)K���t���ǩ�.n�a��H
�
#.�0���֏of��,�8�]�s#�}I��C;`�+������EG��5�X��B�ol:Y�gt���u-f1���A��c��mʙ3>yC�ޫ_��.��]��乓�H�Y���;�A�:Qź��c��GK����������2QǰR�ŀ&<Tڱ���S]���'~��y��^D�RC����o�ҴT�I���ߙ������诔ۥg`��R�r��g4h-�ي��zF��cw��]�;K��^,3s��:��a=���q�/�`o7 8��$�8	���*Ҋd� ���z�-�G��:��V�4
����-\sMɸ�nJ������m\�q�ũ[k�e�K��l�ؠ�L�ݷ5�חR�|y{�>qD�������e�YA7,
s4uO�`f�-q��%׳�ٱNFb=�YLF�h7e��z��/w�_;ź����]{��{��w^_�V��&&Έ��,������f���'+�GO\�mX��w�ыV��\(}��Ʃ�ń����K��ڧ��B����n�|d|GI9w.�L���_#L��}4�SM�=��9�,[J���ˬ��;v2AǳC�T�V0��gCԭ�۾�r�����͹�I��l鉮�-�+s
l�Q�f!6�L�j��ИkS���B�����&Z�m_Q(<�����ڏv�H�G,�����@#}رɂ�Y��T�������.Ƀ]^���}V�tybl�4.��{�O5�0�ݏ��r������l�}ײ�%��\��.ߴ�i��Yj����<�Nq��r,�R��^��nڴ2I`n�:]*�4{@�>�[�;2U�7��U�ҷk��$�ΜU�v����L �Hldby'�}q^ �J��a�(5}:3���ޤ���"Gu�7�l�pd����
�j�m�Z����[Zר�p=�UlA����U�a/qC�t56�u�������ѧxӔ��q{&��r���C�J��̫9�]�����'ek���x���%ɼz��J�/���v�Y�5G��F]Br,L={8k��0(��IZNX۾���[}ۜ�fd������[�Z��n+�g\V�EX�� �[xEg�4�uoǫ��f�٨�d��t$Y*��������#��2����U�]&�x��<[�r̔��V�U�7Ϣ���t���뚕��ʘ��9�B�5�6�����,�M*���k��r˜��PtZ�����BT�7WP��;�l�3u!x~�Kus�{�ON��ٵ���9�8��d[���/���]��|���à|�� :h����Z�q�3
]G�� r��7:�f�ŝ�[�N�zl`+����T���X�Wy�t�gq�����+��wwt�S��}�nun���>�{�j��uФ����x��N��X!����$j��Ȕ�E�4/ܚ�U:U:U�պ�r2����T{p��<�;�P�(�cE���Z��-`/�6���r���"I��	� ��J�GN즦�HՁ�/*,޻��7�? �$���~mw�y�J�l E%��,2IM��|�(�d�ƴ����	&�e���r
�I�MQ�umQ���c�IǑ�{pc9H&�T��^G03�ٙ� ��V��gKN��D!:b���h�j��h��+&��L-�[@u���z�^l�G+�* @ҫ�@\ <���m�qE�;����A�.�hR�����Hã�c2�>���׃���d�h�ر`�yݒ��t�[<%mۧa�z �R�tӲGL�I�hV�L"�G!�LR,����7q� �AX�:^��MJA4J��N�b��@AQ ��Cj 2����YvV^	g��oaI(M*;]� EL�voCC�شh15M�a�z. t*�4vm;��}'xQ �\5�(ŗ>�B�\�P$�@T�"���&�,Y�%��kE<ʈyl�(�D�F�q�瑜t��Kd�H�a����r�!�E^�]�AeX[��5�A��Q,/M�-b��Xp�i4�֡�42��d�uj��E�l��u��(K�IT֖������� Q�>��EQ����~�=�o�� ��?���H|ߓ���9������ή��M��b����L�{���rQ�_,��zf�\/wj�C.ΞH먹��$�iB�V�p���{�N�ި�`4��'LȺ1\�*��w�P�zq`P�ӽ�u�OT|�v��{�J�1,ǚ�ܙ4t�7��i��w�xm��+W�6a�ʮ4��ù�A�;Nر���`-٩[]��yӋ��k O$��D/êeC;{^J�$��8�9Zp\(�����æ:*ؐf����l��TN������-šcy����-��1���n��t��ڛ�������UUX]J��K�w,�7�V�$`�HtM[��Svv�//��;V�9���X�XU�p�9ҡژR<4�)b�V^���'D��"
p��hp޷P�!�g ^][ìc"��]#Y2�3 ��[/����Y]�Km6��W`��N�C���mH��X@����&��v䒮:���;�<V7���(V��_/�xƑܩ���&j^IzGd�
+�{�m�Y��'1pє: ep\�]�H����޻��RN �.�)�
1����Q��aB�An� ̻�*O�-yi���M-a��{�qr�h\��̙Ɔ����ܞ����C�����۩�:u�]u��[�u�]u�Ѯ��X뮺놺�ɮ��u�]8ON��]u�]a��]u�]}���f�뮺릱�k������}>��n��:�	���뮺�ө��k���d�^��	����:��{u�_f��u��뮺�5��u�Mu�uӓ]x뮺��[��뎦��u�����kvf���O{��B�ɘ��7u	B�C�ifV��ճ]�O��F�\I���'k'���w�H]��׻�ɛ�
��ڕ��OD�^e��D6���}����0���'�YLgvc�{���=t:��1��7��j��t��[��Դ5�	����m.z��Y��;v�؁�������D�lux�p�u�s����­X�VI�%8Z��-�B��2!(t�!����U���-��+d�aiu��:]8��b�|�t��+�e���z�ӗG�yf�p�[���Y��K�9�&�z�e$�(��l��,.��B��}K����:�=Р��|�A��f�ٖj����A��i��B�B�ʊ�u��)}��f�Jlb�Q�/ss12mU�Bz��:�P��K6���V�(�v�!�fS-���]�RӴ�0�aսyY7f L�(tŇ���*WRhV:�������`\�,�x/�`]�Ζм�W��d[-�+���c���&�_eZВ5�v	���!�_XUآ�=�u*�U`�n�V��;#a��A{��b�4��6���6��;�<WL�ˀ�J1���@����+&���]��Iv�k���٢��F�ER�`�G�v���:��%`�fl�ﾢ���=g~�o�zk���=���k��i=��ֺd�_N����u�]z5׷��k����뮾�]uӄ�]u����])u�]=�u㮰�]u�׷�������뮾�]u��뮞����Xk����k��i#��]u��5�^�R:�	��d�]u�צ��&�뮝�^�:��u�]z5׷��Y�����kuғ]u�g2���`SE�jD���r�����ѓ4�A��}Z��\sD����^4{3��.OWm.�I�=�B�=������җl\�{mKZC��U��S��掰^���2gq=��W��8�-;&����K2��,� zNV6�����(�
�\v�Y�U̳E�X�c���+��/gfa�.��Ƅ:��Yݍ�"�PV��BWZ���T�]�~���G�Z����bJ�)[X�7Φ��ZC/��m�4��C-��t�q�\�I�{ CQ��!��ܔs	�^!�oS�<e���X�69� Z'`Duax� �)�K��E�,Uu�[�7~�a�t�;ز�Vsf�T:m��U"��˦�A���k,$,�4Ʈ�ډ�v�����e�o� ���x�^���T�jk��ʎ��VK��Vb������݇�d���F��-�k2�Y��a�Zƒ�{��r
����֥:M�L*�t>�m�+	�n����)��"�.u{q���KD��Z5�/7�|�^���9�r��z�c�
����p)]���X>$�V�>�p����ؗZ!�+k��k7C�$���n��ҟ���~�F����`��ۘ>���F�p"�Ah��M4�M4�M4�M4�M;4��i��i�F�SM4�L4�M4�hA`� �AX �F�0�M:4Қi��a��i��M4�L4�M4�hi��i���4ӆ�iM4�M4ӣCM4�M4�M44�M4 � �AAh �(A`#+�i��KC�t`5p�&����c��E���-7�B�8v�y���mp�s��n�v*HPʌ���˖H��"]����_P�Iһ��_^6���������Q�ˑ-S�a�ܫX>�۷Y��H�:����,���_6`4��2�v��V]*��$cF� \;�\�������;�sC�w�F��{i$.�&�@���e�S�yU�����k�|4�)����0�]��r������"��?[c��n*��d��5��Q[v7&>��#J{�k6Pj���F��Fu�ej¸�~�(�x�ĈW�p���:�^VQ>�ť#6R������jW\��*�����gh�ˀ6����i]��GB�y��ǼM�v�s:.���0恙�ckYrV*5ϙ��3x���UA��p��jQ�c�U��w�������쇝��k��j��hHq�l��;��9����
�um	x�}�l'�f\!"���9�:Vh��]S�r�^��V�-ӣ�c�q��M��*sD:�mm�Pk�[MJ<��{�7�83L)(���t��3,[� x.��>�˵H�*Z��A�� H���E5���8l�Y��F���B��,f�2�#u�Z��	������.(t���*ܳJ<�E�qry[`�$si���(6:M�:R�>�R
�&�.���p��| |%�P�,�5/������x�H�Ä�8p"�A'�Ni��M4��M)��i��thi��i��i���i��i�F�SMAh �(AA4h��F�AAF�"�Az4�M0�M)��i��i�4�Ni��i��M)��i��ti���M4�M:4�i��i��i4�M:��zi;tBh"�s̮,�XGW8+�!�sirovդ�»�ot�u,���[Ԑ�z��es�W�q\K�SC�׍Ԣm���5�==��x�̎*��SO�ʺWIS!%�����	�,3�b!�5�hTFk��6h�mr��U�-���)����F����[ty�[^�+�ڑ��ҭklŘSa����4����1A42��k�5]�ڐpA��%��ۡ�B�a�8U�:2��|��[��Sԙ(.B�R��P9���$q�Զ�����X{�{GNN6��"��ugE�[��Ӳ:z��Ήӕe�b����(#p�ٗ�!�d��x�'0u�/����`�K\�����������Ӽw5.ǲʳ�[�,��<�
|Z�D�"�ގ��)�_l�4�4��T��x�d]�[M#��!�[�
�)�>���dF��|�2�
��|u��I��[)�A�׫r��+�@�4�n8O�Z4��$zY��ʊ7�%����Tw�9�}�֢��<�k#�i�97�z�M�jr�OEp��[9�
Li�����-\bD4���>��ϡw�I��Hy���M��~�xd)QNcU����j�'�bI�u�	�u��Ѷ�W��1��w���*�N֨���5H=d�:��s�ZUR���,U�];��������l����/���TN�D�|�*AF�3:R���3�:�v6Y�k�2��Qtш8���h�
)g8�,e�ʱ]|�ӹ�S��J9��j�ݒ�1v6Ǟgsݒ���)��Z�[2�u�O,�����=꣠�|�8c�Xt���ktPl}��
���4�}��2R�i1��P�K�
t;~W��1jvoE%*hh��8��]�ۯT��=o�U��ޣW�iaPicU��aU(7�G�;ܹȟK7��ū%�Z���(6Z�!��Tj���L�}Ȋ�j���@���w�结�u��� 1�s"���b��v��P�ݢƷx���):��Zs}�7{�ş�v�z��̭��s�~d��iJ�R������R*�d��!��[����[t�I݂�Bj?m5u����s&W�^oT��4�fU�����GYUx]�t���Z���E�U[�ڐ�^d�vrZf�E�Ш<CO�@2�i4佧bl�m�4�5�=T�@7e�Ô-�7���>��0�<m7��y���)=�AP����N�F������6��.7W�BZޒ\cr���7��屫��R�VŦ���U��*z�S���.�N˗������T���1�jU.�]�j���ا�k�2��)=��;-㽿,���~�Wn����A�C;t#˱��#�=1GJ�ЬR9w]\^f���YO�mA\p�|P8UqȅʐaVk4�i}W�e�LOZ8�$:�=�ƥ_�l�V;��[���Q[�4Cn��Q[p�.@5X�b��\�d$U�p�蛽v��ei�*���BA�vu^��&(:��Z��47w7��6߽Z6�^1QaA6�[մFih�`f:"�:�,�<|ԙvi���/�����<�n���pW��K�r�n4۬����k�T��C|���>�V�A��Z�Z;m�n�Cv�Q���\"���]+�����e��x�_
4���\�s���c�.n�-4L�ר�t�T ݝոb3���=��JϜĠ�l�|�����6!]���������'�ޱ!���/Gh�5�:�����؈��̅�ᗦ�(�ı��A��6�:�����{qQ~�4�x2-�d5�M��W�G��;��'��.|�v�m-mi�LFų,��*ǥ��A^=�;r�6��FCN���?`��dzƵ*%�6��)��Vgb�͙����J&%Y��N�$&�ͼ9��5��ܮtT�DV��mlk5y%Wb�@փ����nڝxMK�$��+�g&OL��z�Sw[wvYG�kgq�2���|V�t��%8!xZЂ	��[���� �q���ě��tt�J�w��wS����Tj�I՝Qa��}ֺ��=%�&{F7�%x<�W�N޽}�;�=C��GbِeM��� t�v��o6���Q w�Ҷ��"3L+�+���,�@n�or�,��P��R���+7�Mwrmk�Em[n蜸��j/��s��2���_��mR����ǫs-�R-�(�oph�\p�����d�+�Z�6k�bQ��B,�_�N�K�-�+���ʗS�*�����t�&uQ�}cOT�Q<��DX����?fQ�uf�v�Ef@�[�r�r�r3_^hKoES�{hVi�]���%��$;����GG�>�UWj�I���P�]\hKE��L{��.�7�Wa;�&�n�-��}	y�����Օej��=uw��I�E���ff`�����rZ6B�n�;Gk��k��(�[�z^Ͷ��vT���j��(��O�"V���K��F�u�Pa���F��ԩ��)3��
�m�k͖Wc׷���,m"�v�AGǑoyΦ.�=���"�՜s�-t
WmZ���VQ���PA>�9�<�K�Y☮��p��s�X{)���/�Z4��.�"O.���K�a��K�W��ս���p[e�u�ƫ��:N�y]�&�w�ܽh�åj���%n=�=vE���%]lK1벎�,�>���0i2W1��;n	R�t�.��+6����U���K����MX�tC$�n���y�M���t �c8��=��L�y�'�N�'�n�9�9�D%ز���z�A�M���Ǩ3����ś��2����W}`˒���u(%_U�E*�R�#I��jm��9��l�\���P�b��r�5�o�W3Ҹ���*+P7�wI8u��N��]�D}�D��(��3o��8��Y�:�<�DhW�@�򘍼iH��hq���l���㊍���(�v@3xa J����V�Xv
�n����2�#��� ����mբ�,����/r����$�ΊD4�[��N;�h�/��4���p��s��S�fL���Ǆ*��=��� lP�s��t�)i��ڠn5^B�&ͤB���
+% ��y�4Eb��>`�[��]�3qM�5�%`;�C9�IM֬$��� ���k��8�N:͝%v�y��:��Q�P]��\���'����D�"b��s���(��d����Ȕ�-����G�МH��#�Z��V
�438G�d�̆6�� �N�疡���!��}wx\�j`;����ɾ��ݤf��f�P���3�e����j2%�m�nLt+�[%�j�40u<F����\����3��z�x1%u��!��z�*ir�IkVĈ���z�d����A�������C��ր����'LH���(��E�3x����*��������L���S�42�k.Ǜ�s�l����xY�Y�2�gX�9M�	� �!��+%�=�h�1�k�gV�5v�i�4i	F�.\�m�Ok��[x�2y�H��V�E0�)�vl���fօTf>J��_�}p.K�b���V�ZMC,�1�\�Lf�>b�p]ݺ���0Z�a�J���(p�;����0�����{^��֚oWi��Lo.�n,<�*&m�;�ǒF�yŸ��H�<ۆ�e�r�&�ԭ����[9�Vc�mZ�Nܡ��������.;���Ŕ[��ca|���j^� ^<,�:�umr����ɺ�J�6�]�zL�Q"^�1�UHxo��K��,���2yL�Bt�F���w���\�,o�^A��`Y���+D��޻ �6p��Y�f*�K��H���j�4�,
nB�M�8.��5��Wpba	h��������\%i�´M�S2nA���÷Ěb	�`��[�A�x�o!c&�}��/0�q�T��7�������0S"�����B����t��EG"�3iЫS��7�T�5l�����EY��+��־4T�ګ�()Z�B�w��X��H�O�V���Ҕh
�d�$�!z=�]���/��"(���!�ߟ�����+�����Ͽ�~s��N篿����W��E��܉�Q��ғ�&�"������t1Ǽ߸jQd	|5d*b��F�0��!�ܝ�L����Evk���m!��w�WfI��<O��V[�����d���r��pX�Kr7�6��6Ƚ�dH%�N|[�������U�f���V�L�&�kԧ�}��4��FӢP�'�XPVvk�:�^)�79'��:��Iݗ�7w��'�cJ+�5������v����v�i�ƞ���*���z�,�Zq�J[�ʺ����Y�s��62��Iۀjq��B��E�#6��tR���� �}��wl\�l59�(�w�*ͼ~�+y)3m�di�QWK��>p���ۻ�[�k9ݓG�N�!f��ᆖ��>��ґ��:	Z��"�/#;*�'js��g�z�'MRg�1E@�bݮ���ז����U�7M��kɸ	=8^f,-T�9ܰ����*���s���U�8^r���]���}��գ{Wg*n�y�MT��Y՚[��&]��,�Xų�N������k�=��p���[�uǪ��*�ZÜ��,�'u�IS�����]��疮L�K�a��ܹiT�I����q��K��䩬��o�g)ۧ�j�k�$�(u`��5ԡY�L��T��ѭܵ0ȝ���=)��=���\��r�U�"�1�0��� ��y�4�O�\#� ���AҤ
 �A,�ҁ����H�=PrU#YE�
Rڹuk\D�)!�5ܹ��E<�i��i� ���b��7w'8��]0PdH0�h�|�؊����B�2L�[��}o���������ӭ{7ae����,�`���d�H�C$$Z���,� F�뮾�zzzzzz{:f��ƒ$�G�����a�"wq~usb5�pB�$%�(�HB�a���::::::;:4��Z_%dc8�9B����wD�^]���z�m�����Gp99���w..:p�k�wvw[�n�}{�����M�cp�ŵ�Ȥ�1�C���,X�C����><���|��o/�w��7\�r/!�+�ۮ�r��ܣ�j��u�ˮ�o3�ڢ�)�8m�����r�u${���r�s�m���ws���6�{��.�s������\�wrN����r���c���뻧]λ�㮜�kr�[��eN�t��$S�,�p�K,�y*�R���9ڗ4��%�4�}u�r�jQ�{�[۝�I{���u��n�5�u�.n��l����8r�ë}笲��vĞ���+$��ݲ��\�����t��5��.�Ҽ�.\�xY"�67��]�7s���){�P˦���8d7���]^q�]Q0���%幽w;�����X����{F�7"H���H�������k���ޯ9HJI'��)�2�����6�S�\
�o#��C�y�=�Q�Gs\�v�X���vr�ǻ shVW^^�9���]Ck�M�ͱ[a�<�0��Yh4B#T��g��Ff��B�ʛ'�~R,��g$�{��fˉ�u���r[�#����}���us�:�^E�L����h��}�n��s��[@ǰ����"�}��D��t��"~�����ϯ������#G� Z�O����i_bC�f��D��ψW�E>�u-��.���j~W�+a�g��t�E�fpou�rV{9��J�*���k���k�^��mY^pYQ�	�ģ��f�����~Kzl����F����lp]b�zn�n�ӧȑSk9�)}��(�qv�	�T���s|'ޝxg�y��{�c|��$,g��W�oVw,����h�����U�n{5�Fg��}��{r )�ExV_½�*�<$�S��{�	��*Mq�GS����D�~U�!�G���^}*߽+��׵��F����:�άy�u�oԫ'o9X�j6hK�&ugS 7Q��Z��Qom�.+��n+��}�<�����m�cQ�6�tiJ���r?�x��*w'V����x>���4�7�9a���U��L�&oC�.��+Es�'���o0P���np8l����up�����VM{L��~�~�W����oy6�g��S��b����Y�}1����%a�ĻаU�[ڡh��^��s����"�
���p?�uv"E�Yh�> �`xV����	�%Sr�]f���O<�����J�>�1?���Ib��3g���{�g�(^VwoQW��9�,�Z8�cv�����*��o���� �ؒ����=^�2ׅ��+	U��B�^�O!���d�u�J���4q@ρ��V#�<rke��3:3�3i�+�����n�����}�������^�I�˔�����^�(�0n��u��)�ǳ7��MLd���k�~~�����h�ȩ�=k=����:�v/�(h5h���^�p��C�?}�T�¾�y>�q��o���j�.Ȃg��מ�)y�rs��g�QϷ�H�b>�����Z}�u�RR�rm�R�`*2�t��Y��Z�P\:�<��L����&v��ӷFڌ ��*5)����-n���U��:���jN��?-�/���o/��i��
��wq;�iհ��1���e.�j�^`$�W�o%�Ck��t�߭���+��*�Z��<|g���RM���ʳq�~���i��O�=�{�������!�2}WW�<�f�f�!ʕ�]��a�j^�U�Ϳ�B/䲮T�k�b�B�9�=���ۛ'���n`��k�55�>ꇺ�[k�vk����%OT����Y�oo�zw���vf�����ݦ.d�s�����~͕���;O<3(G�U:�g��>Tn��}�ʌ2f�(�+�D��"�a����x�l��������.�غuN���^��>���:�/{��>�R������wt��ΏJ�b��gɧ��o����y�o�O��z���֒�W�x���K]�����#a-B���D�����o��S��>w��0_ʼ}K�*�K;N���y�����W5�W��C$�{����5�S�e&����|�5�xե�Ewfeq8;�w��-ՓKol�=�T�qL��2���&�u1�T�ܡ�"�f�K|kz`^�ؗ�o�jbݭ4ps�݅�ű{!��yS���[����G?c�^�0V��m�[��A�Ve��]B�Q#�%q����E���+�ʴ�M-��Ss��K�:)��� rsw\,�	�Ux3��Ѵ��p`v���`���wj�,3��&w`�~��sSЌ\�{�r�����my�=~����v�����5�x��(,�@+1y(�+���F�����RX�8RŔ��ݪ�ە��0�;{��wxl>t��v�ʹ^5��\	�[�y��ͥ�%�u�9p�W
�������yk�3?*���ZC�A��%y��,M�y�E
���׻��A ��d��R�T��~+�*oh�~~��_T�O�U+�W���p��m%���>RG��kƳ{�پwg�[A��^�W��/�S�+�I��n󸡹k��<�f"����O�7U�דE��N�כ��iI�>��|��a=�]�-Λ�����U�]��G�y�ɴ!���[�9@M��ᥛ���Y�G�%���{�w<�q��*�2oNy��z���	�Ls/V'�Oub�W,��4�ŧV�k(�,MEM�P�����.KS63���{�6�Ѣ��.w �;�1����6V����T.w>�#ܻ[��nqV���[h�7i�KA7���B�S�ۛ��mKX,�vAoA���5M���EFKA�ս�N�ϊ�`(*��뇥zŽ�]�D��f�p�������V�݀?m����������V��~�
g�"���wM�����g|m$�M*^7�4�_q0vDZ��/^ȱcS�!�j��j �]�Dz�`����P�g$R��c9��jF���k�g˅b=�>�U֫�Յ���0:���wr�����yar^��+v�E��:r�)��n��X�cU����Ջ���]S>���[��O���%{-e"��^�{��[��[Ҽ��V�S~5ǖ
J��$_���i)(����]��������^&�q��9��<�b@��Rۢq3�{�$�Ψ��G��G T|7z��6�^��L��}?� �ZI/����G�}ݿ

ō�+��#��Ib��c�)�ힳ�<�cΛݞ�/��g޼Y��E�xz����N�P��n+;Z�<�̶y9R����S��(��z�n}e����or}&Ժ�A}D}B���!X�IߨϲN˂���Ё�+��1��WՑ��/t���`�A=��raB�@��=$�v�{�)���Wq�mB�a�g1p�ͭ�بS�g����q�P�{�.���*��R�|
&�\g��Q?g���z� ��ZG�G-��{�Ο�aBp-�n�iɲr�;޳Z���g�wqߣ�ѻ)3+U�{���<��m�"+ʛ���A�=k�.�dҎ�x��	�UQ ����s�DXI�g�ҥa���/����0<�z��~Ń�r"��}��=(��T�^U^:��q�.�j�s��X%��ڳ�[W�֯��^�bI�g��k��]7=R�gp�;���96��ΧӁ���7�Y!R�f��h�}JD@��<��o{�xu*��<��V�L��Wo��K#[1M�Ϲgb�^��?C�ƕ��U��7��#PĔ��z����^��a��n�1?{n��*YEe�x�؅�ϧ���@�����&���nOd@ R��k�υ���[�A	bFkT�=^�
�S��gz��<�1�ig��ϳ�����AP+��+����|�M޽6��8Tx�f��[Z���L�������Y�b���	K¤7kkQ�A%�[�����ْ@{�#��x�����'v�E�[��O���̻-���'|.i�:�����
cޡ��vl<���_W/ݱ���fĠ��VT��7��{	��B}�=&J��������W�̟n�`��&����l
J�`5��:u��fqh�o��|v'��4�+7�EfO��7%X�`����&���]w�y��-��F�۵�t;<+�u����k�f�׻�~>��Fǳ�]�ǟ��Wy������Lz�*�~Ϩ�PΥc;>S�r}�-
I�1۷��=�fn�;���ɦg��ho�
�o��~~*��E����_�}m*xv��;|��Դ�ה%1�z|�	�ݟ�v�s/�c�ױ��=V{<��{��ӵ�u�ŏCuE�8�7����@O���}ڷ+֧7Qnw�=s&P��-�ok�۞�j������V��@TB��G�:�t#SW��b3m�I�n�!A1��y��ӄY:�VvWm��(�x
�*�գ�Z�,�gYO������a!�:��jv<�yI{�3��Y��QvQHwg��ЯR�2���ܥ|~<����~S(�^H9���.��f�$Y��/��u��#��72&R%]˻{(I@-{�oeL����r�Q�,�WݬƟM�uHy�c���ܱж�O�h��`�'����{��i+�Xf�����}Sv��p�vU�sU��l����;r<w�?���IW7<f�i�v)E��3dk����j��+h0݊-�W���9�#:������G���Id�"���x���үx�Y�{����=o�x���$�����=��c*�$���Tß?n�S���Ƶ���wҹn��h��}���^B��n�idͿj��U��q�͝�9=����u�Vo���=#�$cQ6UڐV�gum&ܶ�W���z��q��wKν(L�!U�����e-Q]r-Lx�5��V��>�ן'R���M�[�=A>�FA���,M�y���l�Q��j繿0'�@�K��`$e���7�&���˯^V_�Y��.������B!bbЖ�q�������gc�B�h1ʵ�+A�FT�Թ���v;-�맽�^V!5c`�r���};:�`��Wt�<�3ہc\�ԇ/X��eG���q�h}Y!��.S�+���<��^d�wR��t��5ŷMR(VXB��AnP�l�UU4�.}���$���ޔ0�5��l#鯔ā�N�t��,���p��W4���S���M��6Z=꾜>ݝ�������{�ǿE�١����U��W�񬳦�!�Fe���'o�;C:Չ�=�A��������P����޺��/��O�}�yTF��a�[���gzp/.��}�+����3��4}�ԜRcڇ�B�U�شx*&�w>�镒�T��j���g�R N��*7=�*�x[�B�n������e��a.����x��>Ձ	���3�V��1h/��.�Df*�c��Ѱ�����3��j�����޸���X������yo�����C��hy(g�Y��c�4����da佊�b�`��S�"o���0V�eH�\W`�+w�áY�#�/��oN:����ә�u�J��yUK�����F�զ��W���g����L��i�d9A��c}�c�{2%^�AT��/w�E8N}u��D�o=���ڇHq��t���[�U�/O3@ � ��� M ]��B�P	v�SU�����	Vڜ�9��m��V��!YV���eL����ʋ���f�&�6��*Ν��5|,�~����!�2}�����KlRW�D�yg�G��c��ii5�t<>�1t����0��<�K)�}�������(�x��;9����ο\�]��;=�@z}�w�=�7o��3\Y������̵�%�EC{����b����{�(�%.�6�W�W�H� k�5��n?M�}��*��;��;y�/;��ٵ?y�(��r���G�7v��rz�o� �5W�*g��eڊN�\�כ�8�I+�O^Tf�~n�#��6 ���b�#����)����Y���`{���#o/�������ErӼ��iY��x|GW��V�8"=��^�س�o��HU�<|1����n�ee{��ЛO>����j�F���ٹe��w��z:;��]���N���fXy�Oa�˧~�7�=�"A��n΍0�r�T>o_��<������>���7Y���#ǛQ5��.�뙶�͝A�jݑ�1PG�_�]R�W>�j�����@E
͵�����ɋ�T�	d����ua��_%%)�ъ-}BN[��S}H�GN���V������|B����v��f������t#=ʴ�f˩��X���ʲ/�]��w��e�̞h�*��+o�;�f�pm2�_V[<�Upi�9Oҧ9�[�w*`�J��nq2�(ȳ���%=�N�ٺ̙+K�}!V����vY��+p�»9z�Ӓ��/�r������xh�X��"�U:�	�]ו�K��y���0�t����a�OM��7Vi��v�;�|��0j<+)�*�Z�
�Z]���@��]L�*�JR�k�1��ǌܨ!��^��Δ�P�;'.��C��U��*}8/>�f�x��y\CWz��8�B������j��<��a݈����{Tc_mc���!��C��O*>�s������]
��䭳5+Әq�[Y{=ʕ�m��m���uz�����˓���@��2�.�MA�S{��Q��{�:k,�|�\�DB3����7�A��c�!�ǃ3;�̩�-0"D#��h�zY޶|2������iw���ww�6h�a��h��H�s�e9W���D,7KR��"���f*����9�{BJx���a=,��L����f�j���zv査�,*μ���;Y�A�;f��\��*�:��tAD�9y��7�)k!�klSU��v3_��S�
R���,�.����=r�sާ�*,��5Ы|%�y��6"{Y�]8j�z+R��BL�W��]F�ؼm���:=kmӮy����'�OBGC��ω���7�V��@�S��s��M\[���n����@�݆��Q&�Osܲ;������ok��]���A<K��v��\�^�<�o"9�}��Eء5�p2R��#.系95M���K�h=x�=�ΐ
ej���/(/�t�8��B�1slR��A}(AJ��Q���y��5Օ֗�S��if�d�X��J>+g.��DM����\�%5�t_v��4��'r$غ�x��(G��[�.]����r��E�6�f����ӑ9�v�2��t�q�ʵ��P�v݋ݸ���x%^Y%�ժ���&�r���e*�C��uJTR��
3����kᕀaC��K4�!iM�tWZ-s��I���Fb��t��x��4�kŚy;���]#C̫>��>��\+9h�(�"��<�V��)�;H.Vn�i���3Ӗ�#Α�u�~܇+G`��d$Wp�̽�[��ś��u�SN�͡����؍�/*�m|H � �~'�~-�t&��ܒ�������'�.#�����i&Y"V��o�o��t����v�����>G�W�ǅ���IB{���� <�+��>+�cnZ�`�o׷��|||{{zzzzzz{4��y-�	 ����\!:wwHK�n\������$~�Ǆ�A<,xx`�bŋ,XѠ��$��l!��v���w�����%��2�������I�E<$xxx`�bŋ,h�~�#|��F#~u�!IL�&�����wtSwW D�߻W�1r�EI{����湈���s�s��	�3Awv�]0.�z�s�i/����E%�\�L_�q�7<�
��dM�E���^WH�4;���e4�WҸ[���sro�-&_N��v$�(�N�_= i�Y9\�+�ʓ�$�!��sW&�9�\(����}U�[�e�+bs�å<�4^v�C*��[}NFK�ch�B*z�iv����I�}E�̥;/�"7DU��>��@� w�I7�$�J�}�Ne~��}�p[@�`�����X��zY�
_b_C[V�JwRܞ�U�HF�8̺��]�}��?<�xa����|.sd{�H�À^wZ���σ�����r�"�{�(DG�Z=>J1���(H���2�,?3?p��5N�{>��=��/��f�b�vB���:�Lv���	�_*�L 
���)�w�8= Q^�hn���,.�:x��dz�m��([����U
%
ڽ�W�cbe�� X��;�����7�6����3I�N�����*j��;v0TL/&�s�֘U|`6��#T�S���z��h�w�=�&6 �=JұHL+�PF2��]8���t{����W�1�ɜ5^���ϲ�ܭ	��`�ָ�I��G�j^ i��NF�h���~poŀ>#Fиu�b�~bI���ff����nTˆ�()_@���Ծ��*Yŝ\�tp W�˩��+���R����@��~P'��ޣ���ܧæ����I�k�!�}�fS�{d�}�J��O�� #"L�JÜ���#HEő�9"��N��{�'��x��W �OO�X�j����St�Մ���G=��w�^C�-&��Ҟn�jt��k'#Zo��J������żr�p�wA���Ih���u�E�Κy��va��'M��b�;�}"](�N�S֚�O�t?}+��}>�M�3VV�>� \]K�nqJ��!4�¸PG_�<ֵ��o��sA���ۨ�D����=��o�	r˹�F>�����|�{t�� @.²�x�����یY�E�{0��|>2%&O��A��1Y��=�������G����Jn�(�T�Aj�/t�#t��� 1S����)�תǯzӟ��F�P�
�������J���7��w^�.{�Y����O�+�<(��7�R�}8;�$9����UO���"8:�#�M����N*�X�����]��(�� �5��2������8�H�.�c�5>���|ܥ᾵3����'�}�Ecy_�K�s�,ೕr�-<���%�"4* RyO^���={^�q�F]�*�����v�c�HQἠ��[��a��_�`e��/Τ��W>\��3���ꣴ8Y�E��r��*����d�X�͏��z���5u ~�p���tNG��ڛ�]"#�|�t7�ׯj��K�>B�V?���/�+W|5W���P��zb���#�l�Ady}F�n��7��}�au� �5hVV(�����pBϒ�Y����⪍>�T%h�]:Jf���hDMZ�n��1٨QO�uvU�_��~�^#�|)����F�bթ�w-�b��5���֮ЍwD�ń�nY�ٕ�i��Fsk�J3���Tti��ט�p���ҡZ� ��#E��)z��z����a�
2s׿���箻�&��L�YA> <~���>?=w 
�.��� ��Q�� 8_34��i���g�^F���ͮ��3�t� 0���ﲝ�N�?8
�{>~�'��z������|3ϣǽ�@q��m/�Nv%7㆗�}� ܱ�v|0OV��DϽ?TN��AV:@˞rp�齑G�x>Ұ	�l�b�������z�J��}��S������Gj7�9���O�ꄨ��!ء����]�#�u���b^�v�������
�����S��4�3Q�j�nw��@	�.��.��&~��q�����i�z�l節ȳ�.�W�m]�/@y�x��P�j� _k�������TpƩK�"���8ޫ������X(���VCs��i(Y�]���*̪�aFߥ?(���;	�(���s�_sI[[�5{��s�c�d壟�>x�r�D�K�����d��W�>L�C�+=�3ٍ�S�u@+����(�y�g��@����:<�"��4����B'�E"~�':|Fq�<�����r��{�ẝ�&���.��_:�H&��SW�b}��`����r�%�ܢ�λ��Q�w~c�����W]��y�w�/�p�}��8��t^h7��l��]�87��D݈M�;p(y��8ܺ�˞���]�s���˥�I��ǬI°�	7@�+xN�����8�l�z_Kcnp�ҋ�V*��TA������_�/�A�ξ��U=< $�J��.�yw�� `�c���!')��`���#��#�����$�GeeN����|%����X���7�[�(5��wKÇ{����x��wA}@���=����̾>0d2�2�zeo� �h>?�z�;��~�&B��
3���j]?1��-�h�][ s�L����R��>�9�}XoGw�K��\�����H�6��oٟ}�E��J�p���a�w�2"�F�ڟ���'ɏ���s�SJi3$
(�<�� �C޿��T����gV�����5m��L�vw7�0 �Y90Q��>���n�\}5YG�1J�G�
,r� -��9��@ ���T��ލ�q%
�HY���q���� K��"=�O�I����rE�ޞ � e}%��� ǘuN�������&�_0>1���_b�ҤV9�|-�3)�f�>X�@�����@$V�O�tn��v�0�;3k����Z��8 \������)�{ȿ�+5 8��r`�]&�����[�yBç�)�o�>��N���\���|�h�H����t�T��] *O�3��EcU�[�=�XV��,.���g������Okݵ
�Kws��Y���~�:���ީ+�x&`���:.�{)o����k�\)�h��znu�Y���ʲz���9kziW��bqG{�R�n5].��'[ͽs�2Kϣ����Ҕ)J),�����s���|ψ>Zdz�o�v�x��Ń.��ySFH�=oP�D{5�ǱWl��b���FM�VY���ꚧR�U02[�	!f}��P>x�?ܑ:�H@2NR�T��Ue_��./k���S�����MO�+_�
�Zxh
4D�R"
�_1NB��/�⢖]��#"=]�E���&���|���Y���A�nr7d}�4섍�i|��/lc��CG�쩛��9��`��� - ��88i�T!Y�2�X�k�
#_g�j���x=��X'���(#�/]�ޤ�cr.;n�e.�>+�0�\~ �k�yOо�S������@D7�j�"���d��FV�z��	��'�>��?G})���8s��\�B�ꏧ���DטƮg�6o(���N^O���_�$�����`�qV++���)E$�����Q��r��>�L�!2An���?;�>��
�Z����}4��0,��T�/���)��T}T}�*d#9x��3]�V�ǉ�ڹ�L}�G� ��s��u;BdaUpR��������-Y��
+�J��@�?��uN����I��/p�D��A� ��BȾ��*h2���u�%�¹9e(o�����~�j#ٙpu��8!��6�]�g98�w1K]�_a��c��u�M��l���<�t�Jųkbu�P��\��s��o�G{O��J��T����+Z4�iJ"���=u�>ow#��ܠ/������ ���#\����7����@}#���H!YM}DX�VԲ�"�+}=��۾iiJ1��a}b�g�k�� 5`�K��� Ծ�K�?8�UN���`|��a�,���XJ�1ٷ5X��7� .�� i|��t@c����_x[B_���|��;#e��<�o�v��!{
T�@�<ח��V?p ^�O|�?H�9#��ayJ�P��"��B�fH��j�o<�cb��n"U�f�����q�O��<Ԁ�Ѻ�r��/Cq��ȇ���ꆸ�D�kl�\��Y�}�cv���_�V$���ڀ7�;�xOz>�Q��}S?�)
� �'�PBz>1�t�U��1[3�|ɟc���j5p�ǫ��^�zu��@P���Ӕ��G�~آ ]A�@@�$�5k'��oo6���}��PTp�����W\���{����=������ �'%D����Tz`����fi��1��b�3��0,s�k��?����G��u`�4�ª`�uڞ�|���b9�G�J�f�T�B�>Q��W@�87X0�=0Ѓܤ58�ؼ@���L;�'Qe�"}����Sݧ$ܹy ��TmY���R�|�W12-��͑s8�T��]��Z�
�x����KԺF�P����p%��7� ;u�z�μ��8�9�-��y�I֡�p/֘|x��[�n�$����9s �BE��(�	�
N)�$&U&%Q�D"�� i�h�� �)J�JTB@A~��� T]s��m�㥋	��(����Ń���ϕ��(��� MU�}	����O�=��>u:�����(d8���@��?�t�<5�25_x%��Mw\P3�w�qG��:F��|��X�l1Aw#��/=�d�]��b��Ӑ�r`}��9} w��o�3M�B�aJ~�p�7����G�/n��t�"�8>���e�w������%��� �~�����>�!���S���["�z�w����f�N�zNn!eB`}�K��E1a������r�CC��Zhkn����Z���gוq�U[�ۘ�����/��'�E���X�p�B��Ϛ��u�1Y�#6:{>]B����ӝ]x��d߂ �FFy��Μ��W�a�("E������=�c�TR��Ȱ~�|����ý��4����-Jn��D�y��˪��Ȏ�8_:�5�����Ww�3�im� c��^zŵ�0/[��p�����]o�^��K"94��+P���i�ާ4���q����l(!l��r��v鲤iN�	�ꏣ������;
.g���/������+iR�{Q��S�:�V�Y�4���8o
xVDM�u�SRsfV�7�%���y��ߍ<ܝw�c�J&5��������Q��iuk�:��u|�|��)�<��q���������]�G_.������z�ߠ��5��kEJR�4��@�@$Gߝ�]w��\����@!zB���a����Et�9��НV�Jt��紣���Z����W����X��I����*S�ر!�?��L�r��=Q1�q�5�Fzg��������j]k�"��`迷�S����s�	CG�O�M�-�x�0y��M���9�s=�ގ��Z��zMxb�	T���h.�ƚW�b��<��CQʈ��yN�s�Z�5��0>���mG�ͬ��P&xy��`zã��Ⱥ��/�b9���>���ܶ����p����fmA�Tr���~�=�������W��nl~}��ge�����k�$UI&~d��}�s)�(��6t���a	�����]"ZE^;�鎩��� �?}��XG�-zF�+��|5x�A����?vR�f�Dǒ��v:��Vcco*q{���6� i�)��wj�Jf��(�������1���m�J���P�o�;r��m{��"���F`��HWC�j[t��ኂ��+�#1����W�+I�B���V�I*>�q^�h\�FU�S��Uc^Ã��Y4��{�EC��v�j�hU�T�V[Qr"���i�`o-�Spcۻ�Y���M)�:G��P�*v��7X��b��Cj�nNL�(���gc�,G8Ls����*�Dfڐj&���s��հ��D>5�-kU���
R�U�������KϘ|S��G����?E�rӖ�j�β�8=Zdd��9ϺE#kT��O~g�ν���Y�*}���6�c���e�q��Rڢ��d��O������p�w>��^�-y#�)���C#���(t$(��Ų�9�z��� ��5��R`����מQ�q���àO0�}	{�:N!aEr洋:+;�7Jx�pk��OZ��o���s�ԭ�O|>�����{��f����7�_Z�lÃ|���Y��o��5��sC�=Z��i���֩�J3�/�v,uv=�c�F@ �a�
{�!� �ǡ�\�w��z��g��(|�AQ8|u�}�V�>�[��`F����P^���x����^��6f!^�|�7u�ֲ����,e���aAӒ4RQ�+���s�י+�p�l���6���|�kNT�k~��!���RQA_���7�g��aS�ukG�y���j�>�k8
pW�G��D=0!(��h�ݜ^���n���P���=��}B�7���Q���ϯ1�1s�7�V�c��w��o�J����ؽ>��GP��+�����������R��|�C�Q�xV|���+�=�.������`^�K:����k�M�rt�L�!#q��=z���/��z�g�
{~� ��P,aJ�����$Q����g���c�L�H�Ui�3{5�L{1"T��U�_��_r��~S����=��=��7��V���SB5�z��ｒ�X-Q]l	I�(!E����כ���}��p����Ix�z�L��z��C7���/��&Ѕ�Jy�D��wk���E�_v�
�������Qzw�ܘ�z�xh-���uS
ASPԦ��1a�X3vϣ�K���F"���|����^fָ����w֚�s� ���1�6��j���s��_JN�Ơw�66��'..��M�Kq�0}8|�����1f�� 5`�5�Hx<mL���r@UNߌ���X��zg+ݫ����o�#OF��~G���9}!x>9 Cߏ���?+�t3�5�s4�w�ww��t����9e�#;^@&C��}�06,�C	3X��rf�3����<镪�u���\��?k�Jj�+:�O�Ju�H���4��D	�X�2�C\wΧ�¢ �7w7��U�1;%�t.��1�;c�W���򊞏���"d)]$,�|~����	\RޯGOe��Iu.�\�Þ��2�*�ᴤ�����(+�v�����vz�r�Az���Ol�Y�����ۻ>� ���u����+�^VL՛��Z8
e���u
"=rZ��;�eP�!9���|
7F\�_-ޭ�7F�^����(nJ��^��0lS���A���;Z�N��.�g����4�� �v���p"N���f���s�S%WCI���Ҝ;0�J�9��%�7F�\����!����:j�&moqott����-���J"RO���Om��k| ���oxh�zpi�AZ��l�pZ�#���-��oH ۳0+����j��^C\yѵ;c�5p��q+�e�D�E�X5���́Zt�]���G9���oxWK�*nm$:��FVK�jn� &w$�Y�4f�"N��Co�Y����b����m���%wxrJ�\+q�×��s��ob�}��,@�%��K��w��_gW�,oV����2�-9�7gfY �ۏ���t�����ٔ�(&�ht�\|�f��/(�0�	����tS�_�e'l㽜��K0��7�TyZhq��e1�Fc�L:9�]���0�̥u��7�u���Sf���N�p|��f`��W���u�����y���ᖦ|���&�k�z�;o;'C/���nTY.�����oPx��v>�k���4!)9[
Z�1�R.����"@ �!E�钎��dD5A#a����Z�o�s���Њ�wo� 7A)Ʈ��f��# _���[^��
٣�	R�F�w*�RD^b;�V�]=8�[����D��HqW��<T,9 ��S���4���^һ��#�LMݩhd��m(`���b��o�BE��詉Ƕ=�Ut�8�m�؝�poU*���.�B-5R����+j	�ݮ<%\'�t;��̌��v�!I���bw.�:�j����]yW� ���}�n��3�����	ֵ��IU��ce�;����#���p�d���/5DR�u����Y}�R��7�dק�M<�C։˗e�Hn�L�h$��6�p�$��ml�w"A.r	�lk��n�n\2qُ,��ac�N��
�*;��Z�ݙk���7%��r�A���:�p�m�<�\�|������01̋y]�yR��Ż{P���-^����깡���v����������up�0��F�Λ� $�V�n�'3�Fh�)=w�^t��C%�Rq��mk2Q�����b�>̡���:�+eq
eq��+e+en&q�~�������䮍�g���mN��n��G6V��g5G��W��.ނb��}2ӽ%:���픑W��l��]�xh��7�G�G6�tw�����=gu72�^FR��b�ߧ$�@��]7/�l���T2�6�cBr3EU!mR0 D�*U($�[u��Q i ��N�s�*��GH�R��4iv��&�Z�-��Ƕ^Z�RF
4l!�Tx>�Ȓ���O�ߓoy�X�9,d(J/�M�<x�x��󷷷��������Ӿ�=�H$�IE��I`��*P@�u�]<'�o;{{{{{{||��Ǒbb�s���2]��
h��6�PE���]����E����٧G�gggggggg��ޤ�&�)H)�:Fb�qFD2~5��ro5)��i�G�ggggggg����D���P~:A&��	IF$5Ε�(�Б���]�^[��>7"�p�
+���|[���b�9�wuwv$���=���21%r�4g��!C(�9���"����}+ȯ�l�+��;cF6M�g/9'+c"��8��\,Igήh���d�8nk�SF�9t0s�*P��t�^�]c��Y���F8KO*p�"ի��AuN�����1I.�dT�6��\;]�����*G�i"��N��&H�B���)���a�ɞ�ʁ_�E��V Aֈ6 ȃ
Q�XR�|>D �}25+�lzxW�($RIX���T�N��(���o���ث`�C�����/���_e	��ʴ2C���On�z��� P��ُ��j�G�����.A��@¢��Va�!7��8�g���F��g�PH=L�������W�w[�)\��h�4<��gk�)����i�[R	����T�w�g�Sքf\�U�2$�v)���)��r��/��y��{_������߫ܮ���T�v�>8g������jǘ�b��;[O\s�Ty{���Ɵō���F|V9�����yHGՈ�������,�Q�I�@�5y����sN�=�+|}��&�V��� ���G�n��OG��
p?P�X�Ώ����YR�̝����Ϩ�B#���Mt��R��8��O�U�AT��~x1ӳG��+��;^'�ݕ}u�w�I�Tf�.�P�Nv xd�j�)�x~cϣ��nkd�z�z:e�RUU��U��Y2ݡ=�5sy�J6+#�9�w��wO�-I~��,��E�]�C^�^f�x�o�`L*�D�mQ�)D����BN����<[���6�G�#,?[�N��e�sc���zq�ɻ��]�:��9���VE��T�n�����|���ڰy*�7Z�FEgq����0>h,qvpJ;��5\@�O�c���|:��+ޯ�M֖*)A��b���Ȁ�*��/�]u�<���֝���\�Pޙ��q��3���9��Rd@�c���{�����pe\i������d�������.xY��Lx���>ȝD���R_$u�=����~�����u�b��r�\+�M�8���4�3Pum�)��&�Tf�ET�N�=�::%ږ�g��Y�oѱ��a�3��̺T��R7Jx�g�͘Wn��t^=�fU�>��Mfx�zA�/�����8�����zV�R0m��t��N��������w�kz����>S�=��4 $+����|р��Tib��F��\-��~傃���׽��dp�[�+�X���P�9�S�%_��l�X!P�(!�����X�R��s���ȖK�N��	�s����O� *�/
�Y��ߎ��ұ��z���	�꫟��ߟE)!G�;��A��Eݱڳ�c��Ӿp0=a�Yڷ`�����?5�,��lQ2,
�Nr�6r0o��},��]-eigѳ��</JA�R�}[��fV�Qni�j��Q�#E+��͕�u�h ���ע�m晨8����
�_�F\�܏n����j+���K����
�G�V��h���v��w���la��Kӎ���=���w_Ͼ�﫪��Z ִA)J(�T,BA�K�����;�|����v�z9���mn�)�r(�v�]���@��׽�I�Jq���Fz�<~�|�V���!g�!G]9kg�J�B�Я�8�h=Q��e�}W�#�����o�S3��u���f�����-��T�h�(Eh�G)�ax�X�r���V����zU9�ҽX�x̞��Y��=*�'AV�8������E�tW(�'
/�{�"����B	�M�������l����.�*>��7�����s�)�M��2x�'{�'���֡*�,#��cN׮�x��	����C�L.c��Ϗ[~Hq�R��r���B�3��9*7c�фH&7+x.؞��(k��Zr��;M
^q̋U�}u��yW*7�(?Y�Y�-I�;ww�{Ό��U*�ޟ�Y����)��?.���7��7AOM
����ŝp6"�6�FCͫ΃j���0��R��a>�:�h.Ų�O�c�:�9�??��.����3s�G]�v*�~�QT'�c� \�F@ ��?�P���>u�`�P�927��S!��nfe�7 �Z�;�eZ{�8�h��%R�K�z�X�[�;[�MB@�3��<�,y@�{��1�_�7Ob��"{5��yLSC��}����Q6g���/�M�kN��j��\lu�Y�1fu�ߣ������w�zߥ^� ����k@R��)@Ps�����⳧x���s2�^쌟���t7�&~�[��2`G�!��&vq�P��(,r��±��ujo��uB��ܦ(5��؀#�ֽ=�k�Bp�vV|�M!#���)^El�GW�Tļ�{�W�A�I���H�{O>�[�Үn�أ�7��S�����a�߭�d'�=A��-�����倳S*��0<.��3�j��%�W��<_�u3����trɓ�;���e%�9g���ԋ}[�uE���ILPz`���,+w��|�vulw5 ڙ��wx��!�>A�Q��{���al	��ϹE��m����!*Lx����#�&�
����Gy���Qx�Ȩ%�g�x�q�*؅����dg�ݩ���~^�<??Wٹ[��n�����7�ZC��y# \t�t�
ASP�2�w��[X3w�цv%���.f�Sz߆z�v��s;���^M)�0;���"��h�T�Ъ������hn����LYY��n�缯�3-o�]�k�y�5-P�tl�xGV=J�7�Z:�%'ݲCI��T��Iؽ����K-5��[7�^��v���S�Tm��g�&�<���h�mͬΉ;Qu�Җ�a�R�I��R���#�2#���q!�y��l�Ϡ��V�;�]Go���ݓ�̖�E�쓏)e��Q�vL�z.���w���!���e�ɜ�a������֢��
P �aJ�� 2 ������W>|�oӕ��t0BW�"r��i��w�?+'��`p�/����|u�;i �K�ل_�2�ބn�k�s;�^M}����uj��P0~�1c�U�&D�,E�O�e�	B
=��D����l��\߰eZ���'��a�}H�V*�	�2����2T�TQ
��>=�,wټ�n�\e����˵���7b��(\t�[3���uv��Ds����R-X��d�FTߒgHy���f!I2�z={�$ف���J7@��c��ۿ�����wbtez�������	p_��L5f~�:�,�^�pi���>��� �K�.���#�����^��3���ǌ���+�x�C�DЧ����,8o>f	3~~y�i���W��%�Ԡ�JZ=��eL_K�����x:�<����!'��6)iMw,I�(uI���o�{}�>ǝ2I��`O���m���"�78'�G���ד�X8%��b}=J���&�����7��:X����a�[��i0�R>�= ����g���@����}��^����yOԧEX3���usz�>Y��wj����x`�ڻ���J�k���+kQ��*���[w�m1�g���Į���a�*����զ@�e.����crr����G$���JiL����}u��vu빹��7טna�@=�B?f��kP�	R��)@lPT������w�߫�ٿ���-��܁95��6��н,O�.������>��Ge/�dۮzGk`�nS�P�,��.o��PEj�'���ا�P9�C��N�<~x1�뺭�.�mZ��ؽ�/z��N�l�j>�Zq�~t���#>�
�������Rd�A��G���<�N?� �i͈ݿ^@��辟�,� ў�ϒ��xsB[�P������K���:�>�M	��X;�l��)c�DԦE�8jϱ\0������P�����7a1��
���nt'Y	K�h(|f�w˯�����L`��������4nY�2��"<���]��d'��_6��j�n|��k��TjdG�+ʐ��u���ԺH��*]�Xr[���})���S����3��F��:�~�t�1��[����o#�JX~���'�PT�Z.�G�j�#^ʵ�
4�2Ї���+3=�)S�.�r���F}f<e/_��X���O	ZP7��h�]r*4�1��l/81��yno�Y��\��oc�R��'�*K]ޡ��W���}[su:y`��j��)9B�mr�t�w�wnL/�DZ�&v�:��u��ݩ�÷͉V{Z5z�>\Q}vN�=Ę�,G66�����̫C��{�j�C��h�X�l!J"��ID ���~w���ߞ��lg�e���+�U�K��uS�t/���
24y�ӥ��A7v�v+7M�����XX�.#�XوY�j�թ*f���H�(���$�y��a�S}-D��r�Nz�M�j-�(Ts0\�\����{�5%H";���\�E����$�d�_ol������D`~�?X�m@7x���}����X��c>,�Gh������{����ۨ�ps�*
�A���Jv�����[��t��,���e�}:��bX���=�9��y&��O��U��9����r魜rSQ`P���Oо�>�g�~���{Ǩ�yW�3���٘[�>��P�������b�Z)M&bUX��G���2���e�Zg-x�.�y�DW���t��6�[��;pe5=�	�Zd�^�I@ Q9^��o��H��ٽ��ǯ�;R���^��_���)����9���O"*
 ���-fC�H�^�Twg�����<c0r�g�7рT��6YE쎏���@�s����W����'�/�F��r�#��Xm��&M+���)ɲ��=W�>�~��$bl~>$�2�C�/7'3Ko��;��י�������x)wDn-`

�� �*����ѯB�K��S���9��}�3e^ø�[qi�:����fq�����7�j�Y�_W��Ez����kPB���JUR�EEQ=�������|��_/�'�i:�D<�aP"�0��W="�y�؊�F�_V�/�Sfs����R��fr�>~��3�r9�2<��r������
д�?.�H�Yށ3ҼaҲ�bo��bkڊy�Pg�֓��W���oH�R:�:��R`m����F���.ŭ3}���W�;�]ו��Q�g����?,f|�����tUo�tF}�w�bHC�W	*e�Ќ�k��9�Y�W�\o>rxD���B�SΑ�5do,���Z���B}�"����5�^����E���^_�݊��Q����Sq��t�t�����o[����iG���]��,�������"�J��8.���7����g(�L���т|���K�8Y�q]�\�]Տ��^��nk�|�*��a��k�rf)G�\}5;3���;�m�5/qL[�*^/ nn_���R7ӎ|��E�AT�dp�*���G�zP������f�b�d ��v5�l����z�jD���v{������X/"�Y��������(.��U-��>~�\��n�i2�"��#\�u�O{�MA��]P^g ��)Y�8�Fr�J���{�p�>a�g6�Rnfޚ�ڂ,]��h��\��{��޼Qj�N�����@�xWQ�{��m*͝Fɑ�`YɧK6�(�92�EG�ա����-P\��'9�%�0�U?MDJր-)A,DR�-� Ȣ2��'�L�_mNI����?%e�O|3�P8�ۙ���ҭ�P�4���
��z۴��R$���Tm�Nq��y��� ��������{��T���4�/"vu7y��n}s��s��t�Sݫ�}}�R�V��Ǡ?�!T>!���J��2f\5%U[����@a�ڞ�3��}y�ϥ��h�S2�5��_�y
2��CZG�����djC6:;���rvc��ܟ.�.z���w� ����G�ߑ��tC9�|��TJ�� @�]s2q\�)+��o0���0҃S��_Q|��9u\Al|C��|9�G�P��q�y�.,���?L�0�0˽���{`�l�`��
�������!��~SH�lf����V7w�y_b�hz�b�J�v-�ˡgdi���B}�5G}�1�0.F:K��B�9��A��5��;�/�B�:Ch3����l���j8��aa���zVƑ��~��f��Mm��kn�"��n�\��ϋ�??�����E��%��
����9����������"B.7琺�$�h�p
�
�ãE��	��Kv��ӭ6��or�_*l5�*��K����b�7�h�v���b�q�N(uA����>W@K]���Դ'vy��K�	�����i\��"!�&�M���a�F�g���d��y����/W���=�y� M~�J�#Z"���B@BF@�* ؠ�*���"��u������l��s�#^����T*�iE���i������$����3s�6�otS���c:h�mȺ�
t�T���[ӟ���f�-4�鏗-��{M,����Ǌ��9����^|=���t��FǓ��r��?`8E}!��ǘ�/8���m����G8����lA=���Ź>�*B�M!07��gͫ{��fFD�R�Wq=��'��<^T��g��>��UJH��.٩�(ǵ�,5�������ϛ9�4}TG��5�W�yG92[������AwьXi�I������_b�oA�[�Ǧ���C�Xv.�s�T�������� �ӣ�����TS��~c���3�@�49���In��s/!=k��U<���:���|���>�r�\"2����E��$-���w�o6�:�Q�y���3T}��!�b�&�~�yU	�3c�ef�]^3�Ee���,��!z}������x���J:��V��R�
ɍ�ߊ�����h8������͜��O��X�| �b����Q��{�Y�ݣ۬{�a�d�=ٝZ�'������U;�]�\{+k����Y��m�R�r�1����زs�5�k&\z�H=��9i{�d�/�һ�:^�m+��X��vu��y*J��p#�&NMT�
t{��U�tf���P�kW�9̮1��s.��o:�JdwK����^���p�F]<T��Ԇl�}]Y�f;/y�POr�x^�3��밷N�v�ɜ�w�	��{kC{g^���L&cM��+�:�ݓ�yj���_6q�����ٞ[n��;DP�M�HD�2 �U�[�Ek
й�ԩ�����T�u̬쮜�����K�x�_����~ݨv"5[��/B���U(�P5�6��}�cN������}M:�>Օ���\�I�viu�]�;L�*��%�v��U˶[��W(O�I����T��"���+7=�5;(���v��ĸ+�y ��oF���9�����Ϊ�-!�, �֕F�w�MD�
'-�~ՑBcYVjNخ�Z��5�.�f=�8᫋y�}�ԫ�ά=����\���u��:x��	о�eQ�x6ɚ\1�5
�=9S��l�8�Y�\��+�*�l��K�]4⩍�rg�۽����@p�.��6�K�+�k&�I���\fudӰ���0;�>/D�Ǫ�9��v�~b;C�]�U@Y���+D��|/V,�|a�v9t�,����V��[���rt͓�C��w�7v�8�W\�il�o��[X�
�&Sܦ���^ԥ�����ڏs[�[a��7R��mO{"�����u���6��X34���2C���o���*�U��x�m��lV��4���%������N�iX�k�YV�ʴX�_�r��6�Z�$LR@WT���C�L��-�.κţ�-.�:�����fޛ��b2��ۣ�R�m�]���u񝢲Yژ�79�t�b��Y�]����t��:��M@�ڝ�p�(=s��L߷,z����r[׵f����m�NcT�f���_ V+Al�W:B���Y�y�{�#�WW�6��L�bdj�ݔ&ڀ��'��	ܭ��[�m���e�J':�������@IU�K�-���WJ՜5��Rk=��)��v�t��w�,�76ts��_i��xCʵ������h�� C}ՙRTkD>R�*vN۱��$t`���=V��4��i�|Cp4{�#�I�B��(^sr鷜���ZΖ ��puՇ����.˧�І�,�]t9�XU�k���O��2��_^q�쑊���|�u��k��fɥ�u�M�.���k*�΁&^����驷�d��D�-��e��l��x(0Ƣ�V��W9�Q���Wm�������(�K��;Za�}7F��9<��\
�������׷����������'%�~��E`�&�n�)��xD�˺����{�y�{~o���������������w����I#����f��6��{�AIV<�8a��i�����������?/�{ĦX�lȣ�+�r�f@�$I���
p�OF�ic�0`����� ���I���.AHQ��� <��ė�����(�@���Ă���/�v}�eƄ\�b>�	%SC0��5� ���E�nl�R�/��߯{}8�ID��}����}��۲ �fgu�l2	�;�>u�O��I$�����o���JC�q_�{}��$!��>�RxoxJ��s�o�6�W!�ר�k:�o.ڹ]uJ��A)�dr�d�.�~34���t3\у��Ep �R?MkZ"ҕ@�B@� }�D�ď��v���u�?�A�QR�'?e˃z�Y�}�`m��[m���(Xʟ� w7�E����^a#�W�fd;u>���Q�m�{��7�zq`��k����
x�k�8�R��Wk{`>����~{[��ԇj�&9�-G؁}�Y ��0����~�eq/�+�*���ڦ�S^��n�U���z��c^V��/�T���_h��=0V���ת^�z<��=�X�z�=]��-�u�f�g�g�z��>�T7�FO�#Lc�� �^�%a`\D�v�g��.��W]�[����O}��G>Wo�V���;=%	�q�"�Ccb���n<���c��<{$��>��T���r菽�$!4亶7V{���ϱx_�9&y�eU���M��w��7�1%��6�S��尦����٫^�+c�}'Wu1������r�;g2��u�����Zu�j�AO,Y���6�o�l�4z1���|x�>�}2�޽�Y�y؏1�����E�Z�(*�1E����)�#Tr��C+5:I�Do�_���d����ud���Y�h�ц��};^
5�vM9ty_K�Јмܣ7���i��vx�4tT�����܂�����`owm�r��v�r=�m���'Iޡ�ݯܨ_q�r�k1�(���5����/����{R#Ϲ�yw����z�U5�#�$k[HR��0�E,I		�D�����]��9�|��?c4����aB~vDc�1���zv.>Ȩ�RQ���r�r`fڝ����۪�������R���x��3��Q���):pK>�<�.�H���U$�]����~��X��_!<�S��&�~�g/�@���]�.����\�!6��"�ށ��_�7�ηkR����f
�%�O�?�y�����"���+`t_���j�.#�/-�~k!�Gd�[�b1_��:��ᯩy��4-ܖ8s������u�q������R8j�}s���"��[�9��f��<}xt��Xk�Ę�al�#��ه��Eyu}H�u���Ī�Q�3�:{�����<^3�:�Ɵ��޶4��_N�	������ �W��&�͝��(��ֳ���u1wEÿ������)N\���X{p2F��{" PѬm�5u��&D���Oա���d�u1f��C���,�w����%H;�,X3�&]�/.�˾QR<�ӻ�^��H.��H���!yJ������t���
���oѡ����{4`x�z��w�'3��/Gqv7 �x���6��R�g�u�� �PC��:3n>�:���T�jy�dw����e3K��J˩��ݡ%��J�e8c�'34�VMFquŀl�%����ë���� 7�rRq��!֭`�]з|�Y��,=����ӱA#���h��0�HR�b$� �H�H�>d�:��{>|��
{�ե�ي	�k��ZC���'μ����򕎆/_G�4�޽��/�������y����|e�b�K�ܵ�n
~2��@�e�=�aM)���
�{>�Y��ax�b������0iZ�,��K��Z����L��?�:��<��/(��W%<<|[����ۈ���?`=c%p>�rF����!]d_(���6��(�߮�N&/�۝jskp����??���Y�s?X������0�����)�i�= �u
LJ~R�1ꛏ��)�M��JK����;"�ت̀�^�{�j�20��ju7y��o�p5�U�=α�Z��*+�%RP5_�� �D���lv���z�y��֦��C�)�*��e�8�u�p�7��d?��ůVԬ5��APؖ��B���7�̅����ǁگ�nc��|`O��,�(t���y�g�הǗ��"����ڱs?���@��V�����1�X�W1{�aԐ��1������D�}���rB��
8c�o�`F����9�#��K�$�}��b���W�������R���0�L���ы3O�D�ٮR��ʭ�{�t�C�P�h��y7�)��-�qc�oOm+��s�R6M㹮I#��=�����Il�Hh�W:=�Ј�%/;=vg=��}�H=�M��$BAcZ�JPZR�6�	 /����5�OwD#dLL%?���o;�M�5"�����{���,y4��E!t.)!"���[Y}��@�!](k�����|�x���^1�}HOc����Q���[��7Z��D'�����_y!Ҹ ���Wy"yw�8j|�v���d�5��%��#h�z�ﾹ���V���4r��$4l@n0@�^4~��FB�߆���¥>�n���i��G�*�ną��1jNʌ
�uC�bd`zU(s7Զ�1Ǻw�vuc}U=��Q/>�K�z�`Ji�J�QTjE��)��/ՄV&%��h��Qϝ�w�&����,)e$M{msV{�E}��{=֔�t�,����F���'������],*s=腘3F�XG�V�s�����7���܌բ؅	�h��@|L���s������绂䷆hO˹RLh���R$C�RD�L�s��ؿ���:��X���C����E��u{O����+���"a5�>�	@xs����4�.4@�-u�KA�P�o�'|��a�5��,���ờ�L�HYNi}Ƀ���u��0Sܖ�N,�b�����,j���]⇹:���m�h6�y%�l\�O�!JÒR'�C��I�R�Z��:�hؗ��=Y�j[��)�N�/��kvo]�����#$~�Zа$XҴ�H	
J� ȁ 'Y�7<�������y"|�D�\Y�R�J��}��-@",;��~��~�y�ͻ�[O�A��ܔzڣΪ��J�M�xt{�A��tE��E􍏬� ё˸�������/ogM�UN�ͮ�w���.���m��Ua�~lb�l�=Zg>��L�lCv�鹝���mVi�����\!O�48V� ����1�d���(���fh(��͎����� ��Q�j����/`mAM�k�VX����L�.�|}�c]�nn=۷�u:P�.~��g�?nO{���U��N�014��j��BC����"a�/O��M#;�(��{��Nׯ����+��#��p��#M65JO�@����7�Zo���������ܜ��{���g%qd�cK����r�0/��0�KgX!h�L�¾@k�i�jd����'�
���ۀ�Iv	&�ӥP������F}��*Hs�@Q�~ z�.���x�=��\�}3�sh�u�<D���Gm};�=�3��(�'$?1�Cܸ�g!�g�����]{���3�z�~���o�����9��pj�拹6��גQt[-���w�}��gk��/�/r��*v���fw}7�u�o�'��|w��{�z���d����.�[��pΊ�T������٨�R��H�)KI Y�P�����V�ߞ[�`�0��'����"Ϣ��"iIr��3�5B>Ѕq�Dz�@�V;�Qt�S�99��O�����gg%p������B�
iI�*ݘoڠȭ~Ց6�\��V�T\V{zҖE�)��c���GǾ�r��MGؠ�A��
u�sUA�	�LJ���Q�j<:�xeۼP������B�-� T������P��a���E��~�D(㻛OX�*��{Ƣ�s{?%�`�������X�,g�b5�N}��_TFF�Ɔl)d'���3�Ρ��T�κ<:��U[��8%�cz���Ӱ��m�&=Zrf!29Ufm^�7�.��Et�>�t��Aҳ�nއ�09M\=���d,���nK����Ę�r}\�;�Np�AHٕ�����6������V���x��K�{ y��+�V��ǵ��L�ם#c�=߭��HL6C�GR����q?d
���䆎��b�c/��j@���/�uyK�j�)���!c�g�ФC3�?.�p�g|��wLU)�<t��{�ӝ<`mf��F�N����ΠV�`��I���N�V:��f���
t��Rۮ��l|d-Tj�^��s�~�S�z��	��eX�iW�E3_n����gJq�9��^���Bhf����m����vG
��G=a����(HG镑I#Z-)T��*�
Ȅ�I# �g;���۷��1QC���Ǌ X��<U85ׅ�R�O*�v���L�4&�"����!�D�{m���yyzQ���H��oظ�ݎ*�N�IN����a�1�_:!���1;��i7����٠xp���s�G��4NR�6��^t�����>ү����U���t����}�W���ױ��h(� O}��O��(�zsʡY�a'DNP��t5?��4��W�+s��R���Y+��|�輅|*c�)x`��߃���V{��w�l���>���937��u3�6_�蠯��ʅ%}C��m�Lpa�X�OfY��ܲ�=8�z�A�c+�5��,,H��zſ�#��>�4_��
�<�j�L��1��\O���{˵�c}��g{�Aw~��F��O?���sz��ލT�,�Dx�z�,�|��TWF���9bL�'jK�m"�h�#	��"X�c�K�Y��#0נ7�ng�<P�*��f��l�@�kޗm����^ϓ<3�-sӗ �h�0y��A��ڠu����;�H)MC�T���!O�<K[4�~���,Wzٗ!͵�l)e�C���V|yJ:��פJ.J�W���Ft5EV��o����ױN3��s���y�v֣c5g�'GP�Gw
��^Ыu���c�7�i�3�Z�g�3�����9�ܷ�r��{#�t�+0MqcU�{�=�5��4�@��`����}���]���~�۽�i������a���˧cz�4�2f\7/��w���� �x��T�@=�����Q��5�66��#m�]?k��?�`>�Cz��9����u��=S\��SG�{��B�x�RQ��͌X�1�}U�8r��^�y��S�2n�������X9Ȃ��뉼=s�NN[n��P��`g����-�Du��QCq�V[Y�nq`ơ���\������~�����ѻ�zf�j��T�tL����SS>{�wݑ�o5߳�5+5�L<:�}|�?sA�� �|�'M6;��W��Q����ۛ�<��z�W����6��S{_S�\%�A�� P��xD�z�4y��`BX��؀�Ƒr�=k�̩�6��x�]UG i���Vǣn~�Hh�g� _�+��q�����0��^�����}�q�*��;�N�}#rD�x��#ޗ��ixו�ĚlV�1|R�RB����N�x�P���Ǣ����} J��#��E����U1���B=��YS�������pS�g�z����`�w��7*�)ʺAث�ӻE�!��#�{�q�羬�����*�h�2��W�m[�07:]އP<-���k����8���MnR�@�ᾫ��n�(���<����&ø��m\�A��fBL��f������N��\����;3��s���?�Z�ܩuծK��(��m�P�tV_\z=9�#����KRkP��S�&~W��.�8��F>^�J%E��^ھF9�a{�͈=z�ɔX�P���A����|�M�`z�z�|i��*1��pڀ�X���3�[��ij3�kv{��(�-0�}B�8B��R�$
h#�s6-�nz5u1(�e}�|�zo:V����R���>����B*���0OB�P~T�0�Tr�ƚ�]p2�fQ�<�LNd�;�8�R�;��+ŧ�6�D���"��@{20��.��TW��t��d]|����J@����b���EV�0C��z3�0ʯUU�I�~�t�~l��炾��9�����b}W���R����ѧ_�Р!�W�R�#y��X���$�tj�>]���V:�h���0j�r����x��FsKne]X)����k����91{�e�SpԶf���YT!�W�K�
��@�؞��.��p;�����J�{R8j���裄��	G����ն�8�[5nN��<1{�wǐYF����y]`����=3ӡ!l�� 68��W�}S�f~U��B��t��i�\B�69�ʥ�Uꪬ,��
vԠ%BZ��D�K9����ӚY��KH��f��2e7Yv�����| 4|q�Cv��P�;��KŠg�̝ɋ�Er�o���y��M9r^Ǌ�h�ԻmSS�䃨ow8\�yY��d��޽����}��K~�z~�,H֭)R��(�EH��"2�����9��󤟏��>�诧��c�B��Ǥ:p��
��O�s������W�&6���tn��񁏾��7k�1#o�>�?yQ�K�@ܨ�Hm�ku+��`ʉ��<���|���*Ov�E�] �uT�v�8
=[�h!z�g�*��X.��|�F�E��_����w��++��p]���K*��R)R���l`��5�U0{+~�9X�����^��	UG;��e�fΧ�0�]%COG ���(���DHf]ޛ�B�s|��gZ�HI�r�a��p��[��vZ���,����	��1���O����^��L��I�u�`�v���X�����U��������JϢ������Z��
t��܄]��wW�/CU(9sy"wVhN�D�� ���:q��+ݗ��=�!d`tD�>��1�T���ʎ�1�8�3��C��lb��(�����1J7�J���ߟnWюw�`��J�M&bUmt����6_���1��8#���wP�vؾ��S����x�*��c�͸�i��gջ,}> >���{�ͮe���zhd���EGvKw��a� �R,�]�H_Ŭ��*�ց���S;��vHo�-v�oN��җfa��^���n�\k4��T��ct��l���;a�+�˰��F��=���3���fUA��:�BSh�+���n=�ع����7��h����l�.;��!vRS={���23�3�7�� '�g���E4�ǋY2���),]���̹���sx�� �JE}�goK����I�j�]���m	�VP_��C�/�ޤ�Y6t����A���x��a�}K�`.Ѳ��;;�7�!-��)ǔj^w5��[��P(&=�Ւ^����lT�y�u�6o-����V�I�_gyq75��Z�N��s�*f
��MM�*xz�ۜY���v�+r�f�ݣ89����t㾭���ΰ�x{q1�͡I�B��|��^'z�rk�«�R��НS_>�5�6>7�R�]|�R�%�`u�qPen�����̺���I�(z��"v��������W��V�;y�*���� �ל)��p/z;E��H&j���fN鷂���~�����u��Uh0�Z�Φ�씜��cpă��7;t&Y]j��/$��C�u>
�
&擮W�k�r�ҧ��tK;v����.������˹Y.�V1<�����M岮�)V����h�4�{��j��^����N��0G��SܱF�D��B�=�cg*Z9�����Q쓞��RR{��8�D�(�w�Vs�Ԉ����gN9EW�i��Xn�>;[L:PU�'f�;���OT��s-:�D��Z� ����::�����Hz�����JX;v�\�'|M��wK8U�V-ۋ
��x>��y��+�rY�Z�.�v\�,�:qk#I��  Vn[���1>R"��b�
/1����c""	`���O��>�B����� �zI�����S�ٲ���J}�n�O�o*�V�t��k��v�{;������y���Z��2���e90h&������Ջ�sA+�O]y���>{�;��{�^�:뺔�H�G_=�2�ut�]��q�Z]�����8�)=P���Ǖ"=r���ZxJhfm�S��ȲهY���P�"�x�K� ���4�D��P�:*=w�F� 57Ir]S��+.�T���۲i�m j�9�9:�9�o9�8���f6�+i���Y�.T�@Eq��Ԡ��z̚.�=w	e�E���p��;w�1a�oE�Wgmt[ޣ�r�^�yK��h4u�&Q}@��\�T�vc�P"���D�]2��V�]r�5��u&�>}ֵ�Oii�l�qsA�`i��5��C�[�b����c��n���,*�!r*�X�i�͢U�L�R���QKV�a� �e�����H
 S��d��E��b�K�ٗ@�}L;˒X�畳t�X6�n����f�3>h*�a`����&T�2���!$��8FWۏ���^ޟ����������|�H��2$ �(ߝ��U�QGӁJZ㏧]u�������������j	64X���E���4�M4ӳ�ó�������O6�jH<�4)
J:n�Ƀ�f�_���~_�gG�gggggg�����T�r�N�t�&בF��ݺTn�9��������nt�o{�Gһ �`��5����d��[��뻷�˜�]�k�^G9�n�b߿{�"�\1�ݼ���[�^m��]/+�5�c+�)��7O��6�ˮ�L5�Wz�Օ������k��r����t��ny\�]��owQDm9��������{r�G�!�޶&����lξfJ�~��wPj�+{N�m�r�>�M�L���5a��dxJ�ɳ���;�
<芁�ZG� 
)*+e�!$Iʸ���A7nۮ���k��
$���#*|���ӼݤR�����l͋��%>۠�ޚiW���vܹUwN�_^Ļ�ϋ�s,�7Y+8���:������/���@7�u��^צý>�S��b��i�G�z��? �ɺ�镖T������ix�H�M)/�1��a�Ɇ8�V��L\g�'���`93����%P���iW�9�SZ����(XͪZdr}�,���~�Ds������+]�gޙ6yN�w^��g�Kpn��تs]}Ы>O2� �93_q���U�(�^&�o*!����=�����}��t��_�s���ظw]�nF}�[3�'ﭵr�y:���(@�C�;L��oy1��(�;�/�\4-G���\K��� AAl��O�=� �ϹY�J��gN��b�
�y��v�M�����;Ö5y�P5��>�����\��S%%LM�yeja�>�r�oo{�Y���:%V�\+{j~�
A�]���IO�qμ��=���HY�5�뼼o��'~-{�s�<e�	#ߖ
B	���������/���\77[������ٻ[>heҀ��}h:�;ᦡ�)��fi��vY4E}wS0���:WR�H��{��-ج)�>����s`غYhxQW�zJ���X����zu�d��T�FE�:�Ӥ���U��}.*U��"k��D3j*�g��H�Y;l�����|��}V��R��! Ȓ! ��7Ώ�<}�����O�7;����,Eϴ1����D\W*�����6�+tmT���Gj.�1�OX��j�[Bϔ��e�U`I���`ev>���9�pt�O<�F��r�[R�2�p�D�m}w򭀖nN|��}6VPbTC��T)#�c%��v������9���}�i=SF�?L�C�X��������[O���uR
FWL^s�/�/N�fy��֨���T�j���ՙ���Q,�4$K��1K�GO�f�lv����tc��7�,јzZ���ꚵ.۱��mG:\n���_�1�(�,SZ_.	��[N��x��t���B�p)��jg�.ōς�p��617f�w�*����9�AC�j����=�x���Q���;ƘW�:|Ѻ��䚝U�K>�`����בpL��|>��{])�&����d��Z�N�&��H��fr�\�`�h�j��T���2��i��^�ԡO�]h�������nv<1u��5�D;>��ό������':7�'#W�Tv����=Юj�}����e��>���!���du�aw+s��կh�<��&�7O=Zh�*�v�X����sZ2���8���=�z0o�������Y�t\1���T����r�����=yY��ʐj]��]��Y���΀ ��PT~�B��IaJ���z��x|���;�������+��H�ǂ�'�5@i/>�"�^�=!liū�����#=2,�e7�������=o]�THȈ20 P4�*�z�y]'W�����/^�pw��a�M� ����6��^:���@yXH<����WӞSZ�Dgno�I<rW��+X��O��X��w2H�q�?o�kJ|����hN�?**�H�FZ��wy�;���qW��[�
�(��	<��x��i��5���ᛇ�ғ����H,����ZɾO�~�����M�MU�b"H-��ptC�S��U���bm";rJ��	�y	�}K�/[��W3��0U��C���`Y~���Lao(U)2kd3�y�n��y9W��7J�Y=�u�.؃����hy�U�9���88sfՆj�OTTx��fQ^�F�E��i0k��h�T��Ji̷�b���H�J��+�,l�j>�ˍ�IH6韤s�f�{�Q��l�����;�#S�5�%�}:��	N�Unmoɽ��}�MB�-�}?�?S�@�g�F�ͥ5ԃ��t'O���!��w�������=�(0n	L�N��Ԩ�}c/��w�s�d�)q��'��ɽX�15ǫ	;��o�=����g	�{9ؾN�L��{�1�]�K����;�!_T#�tU���Y�!
R��Ad��~������2Ǹ��^�R����-��j�v�|Z�ă	�f�)�7+OV�����T^g��j�؞��x��4yY��r�� f�������rb��˝���j_��<h(�����7�~�-0R���B����ΪI����z�:jl&;�O��>b6v��U���R���0zL1�u[~E������ߏ�u�Y��������\rsU��]Q0�}�=��w�=ٴ��2<�^8�ُE	�� Tp��)?�����	
������A��:^���S�9���T~3�ᵒ1zF���t'IN�909�F2�ްB�C���_Ͻ{���VбOa��3��0X�O�F��h*��YPbW�CT�
tD�h�І�/�����+��=��a?�<!�ߩmd��)O�Οg�O�7��;�� ^T�{p�{��gG���j��e�*���Ay�Z�=DE;5��U�2"E��9��(F�٭����^��������6����')��-����D��:}�D)�&F�0�����graxK��6�''�DMxCΩL^(:õuw���+�]%_�%�pw�4�cV�7�E�+=�p����rH�0��\�N\�Ք�3��
�n��<ޡ؞U�2Yfgh."`�9s3V�[1-쎈����&�t�v�x�-��bjr��w&��詵�Yv���Իl��}�|� ��	 H�{�{�'_���V��CJv=ҽ<��C�ig�{^�q��m�,PS���x.�`�U���;�\�!��*��K��X�����}0I���Goρ��2E�t{SyE=r}cK����֌TU�w�=�a��x4���<�g����P��?<���ӻ(/�[뫍Jd���x�_\�r�
i�(5!�w�����:�0��~4��%�;p1�\��X�y�A�3Y���3xy`�Η�QF�?'N�UC�H"�qϬu�R�����mP�|g�Ȭ�y�=�R��w��"������b?ǘ�o��S��V��������^�ݵ�^y�:����ɀ��P�t��ײo�FſA�e)���*A#�����a�>�}*���偞���T��ߺT��s"�Ҭԕ8��	��jS�U&<�b�WP���pn��-�N�\lzu�'zN�� G�è�r�]zE�7�t���5�B�	�&s���������%?���]��" }�d�^�Y��01���C3˜�:�P�`���x��-��nm�}1�H���7Ͻ
�b��(�z�a�_)�x��5.�;�O�_fT$��Ew2�Wi허�Rr�57od��fX���Z�U�j
��[:�[��B��V��-I���v͏�xƖ8�W@�D%i� �(�P��e�Y�Nt��RI�zz���u�O����
ZRd������HU�L
��?���8��E+��ӭ���	�u�+�c�t�8��Zy^�sh��^K��Z�yr��6L|Ag�s��k	�z��8lߔ�.WS�q�X�o��w>���g0j�@����m�'L�����v�B���� ��$�.)��Y�W�[�������4��y�n%�0*,wSs�*,+�O�Y���_bP�Bڄ��KMs���Q�Nb �U�X3{7_gԥ��[[���X�[��o����u"[�S�E(0-A]]U�yz)N]��L�hj?�4+�k\����j��Ǽ[��U;�4����������W�Sg*��+h㺼��ҁ�·X��hHش��=�c����+`%�s*��-P��U�
'�Ǔ��7��LAo&k��ߘ���;9ݩ���6"P��-�2*c���;o:�Ð��%r}Y�>�Ξ/�Uh�梳)����o>�Wz�Κ+�ʤ���'�*a��7��s`��^0���5�z��3��hFk��{�I���񢲛��5ӯ��Ws4�����308�de���)Q���c����{������]~�ށz�%��wi��L���8gV�B�������+{����E�v�ȩYk�+sWV��QI��իlW6��k��Ρn�<�\�-ۧ�X�Ғb�9)>��7�n���:��>���֖B��R�B|�.[�>^~et�T�3��qǍJ����)�����0`F��@Q�@(-Q\f�E<<��w������,I�wRĝ�.s9\���u%*�%㛁��;7�.�*��9�D6{y��yl:��iďFk���I�Upr��D�L��caT�tL�?;�譝+�k|�;�K�r^v�H�8���=/b�׎�bb��0q��;*�_r��w_��Z����p�'~�,ɶ=�"(ve�`� ���D�a։��L٭U,_G�0y�u��Ir]9KŘ���o�}��/��~9��Dn�;D�A���������W�U���:|���O�v�7�DD�p8�j�0~R�l��XBe蟴C(�`ţb\�7뜲����0���]HPI��:z��<
�S�S,�5$F"+�9�T}�c�;Z�S�9�Y�Qu,$TR\a��H��/e������7��)Հ��_CEFU�bp	���9��b�>��s�K�C̅�G�s��\eA�G�>�L��XԔ�i16��&%ʼظ��*�<	lWZ2>8̝s5���~�w�;������C'z�)pw=V��Џ��߱�^��F�����B�|n�����]|7��kA\Nu�K�j��Yc�U�f�E���}oIתqUf%�\vꮊ��x���|SV�o_0�nn��f_��4�5�B��D�:�����ϔ�N�@?���\I�������騱��b��R�,#H{j"N�־]>ت^�(7\�Hk���h�8�B�`l�#�mT9k؁+�19�BOU�I�+'Y�w���b�5�$��:J<*���5D\��Sϥ�v-�x`d`]���4Up~?{��˳<E����{�+�Pܖ7�]%,HB�ێ����%:���*M�r�9½~�~���lK>�r��G��=���i���>\~e��v!���AcǬ_���}��7�D)����N|=W�I�J3����gvj��$��kܣL1�)z'6R��oU�T�Ud5/��Ț��}+�󥴟�<Ä�.�@ɓ�5�R�JZ>w��I�3P��U�8���ke󝫗�G��O���TF�=5���\�*ee�A�6ڴHϏHt�z��.�E�Pk})�Hܵń��m�����{��O!8D�煘�)i�av O@kǔ���f��=�U�b�c\	� x�F�*F�s�})ʏ�2)�@a�F������~�̰�'�G�<!T��Ԅ;�y��}����(T_x�&`s����g\����w{ݙ��i�n9����0������i%�V�ܙ������\瘗V�k�sd�K�̵ �iwi�^M���aj����%X[:���Ļ���e��=13M7r$"E������0�!~���[��<���R�vIa�f^<*�@h��zG����G�6�ʚ{\�x7�\�f��ӹ^��̞�"R������`*�	�y1����A��+lC'�*7�U	����Oڟ��GmP+ɪ{i���!W��T긨k�E	yg�G*>��Sv���&i�hgݪo��،��~/_np�]V�+�}�oF`�ݡ�¡3���(�4y����O�3���{���'+��\<>u�4L�?*jc�=��J��<6����-Wڠ���(p]Hg��G@�1#�vw��V��5u��.��],B_?{n��O{��,�ʕ�q,e�):��&����l�nzŽ(��yQK�H��~�c�|�0#t'`�����S��1���z�.������~�[�=�*(�,k��|ě��S�O��� �A�͡��UnV����8��{��~kE�s�Uw�k�`�N�W�v��(�)P�����Wb|O*�c��[��8ݷ/����#�VM��J3%��Y�����5UC�
a�@�����z��������k�SV�Y��V�̛}�8�}θN+&ګ����}�i�-굩�Go@��G�����*J��|��}���P�������?8�Ne�fw˗v�P0vU��H�k�.*�3X����m�������ÜCa֒�Ig�}��<7��}@�|��V��л�_U1��ʁ�埔K��^f�*�ʌdp�����r�~Z�ʬ��[p��GW�����1�/=b�Z4Ԍ.�S���rbӥ
{c�i�Ƀ=�,�X�p��E쉿B�㇫�7�;#���0�Q��ql��n��⹿�чXy�Ώ8���*Zɩj��w^�����,#8o�]��C�.���di���:�RU�9��4�p*�6zƔh�����D.��AC�X��(h��4Mҁ��W<�`�il��}�F�Kc�ݼ;��Ai`����k	������#��S��q�7/	lyw��#��`̑3��<���;s�s�A�@m��i p^!�]�C��cԪ�Q_V����#�B���刿��D0b���wŏ@��Y���R�7-m�U���p;w�w/n���+�#��V_N\��v�_�l����j��g�_� �[�S��
�n�tx�ߩw�I�gyw|�7վw����9�&f�T�fW��m�3Y���`i�R���=޸	��go!;C���2͉�.�X�8�ق�x��k$�#
��A�����j�U�}wr�rmN��q�U��(�Z��;����rk+��<���.��)��f��vܕ�p�6��ڗ�e�6���x��J�k��H�{�/������+}�cC;��H��f�=���w��宲�eЦu�4T�P�I�����/�E�\�Bu�\�镳(����epky�x8�7��֚�OZ�R��L�:=W����=ܴ��+�J�6��"��<�IA��qN�����u�^,<cCp�K�"����sT�-�]��J޵�/�KWFS���a�&�N���n�w2�S�Wy������Hl޼Z,��mbd�W�b���}�^r(���`����wn�R?\�1�A�5�iLv[(7g��Ô�]Obs��KF��m��}�S�N��x5ۯ:NK�H�'��}��]+i��O{��y-�7$=��p�T�*R-��&X\���w���1ܩm�8n:]� x9����5��k�TD�g7��ܕ{)${�z1G�q�w�T��8HNp���+b�Wr�+����f,M��X삩V��R�5z���;��j8��:
�c��6b���h�+�tVq ���;�,�����r���̂:�G�{�]��Җ�ޭ�a�-:�S&���O�̊r�P��I���J�OMZy�'rګq�v�h	�.#�J,�Z��uͧ�x�D�`S^G�)��';�Ax��R�\��]Z���M�ÅԠ�/�]X��'�J�C�9�`=��}|u�N�f��n���Ư�F�4�;�v��.����)���� $E���T���Ī�tc�!�䱏�被J#Ҋ���M�^mt��P�V;��2l¸^���j��є+[���1z��6[�7��b��/��M�"�/�5ϸ՛V*��뻹�O%d��t-��a�H*x�$ݱsVq�v���&��s�թ��T�0��s�{{�J����
iT�t+�1S�@5���O���rX�"3��j̴ﱦi��a�n�r��W/M���9n�GY|��+s/��R�Q#������5�w��WQ���!Զ`d��%"8�o�c[�^�ߒ��s�8����7X��u=C#���0�O�L����)J�\s�2h��cu�Y.�F5P��{�'�I��u+��WF�(--ҳg�Щ+����Pe��7r�x��"n*���"����l{p���B�ɋ�˨����N����:���ۛcM�g8�z�8&���s�%m�V:ռ�]V-]!����W�^�\�Zih�Vg{������-�I��Bk�yۤ����y�g���`������#v����a�����;���l]�0NS8��$d$'p�"�>�O��^ޝ;gooooo�����,	;�'FB�̆濝ƨ�W���t޻=�o���������������l�"�	d�?�^|oz럝�z|yN�R �B�Gp�Ç(D !��+��LIQ���,ܰ�� �
{4�ti�������������4��r'����=e�"X{��9[�9�؜��^��侻�����b�gv����5s��i6��x�y^o/(�sw:2Q�����wn��������e�%�s��}\���\�.�l��gK�ͯ�ힺ߮�.kǺ~���}���|�����o}���u <�/*Р(W��b��b�-�=۲<�w�m[{�^�ˣ6���t{m醲�H�w�\u�;.�b�`�t�P����:j�`{����AJ�˷��g٫�Ϝ{X��XC~�yW��\}<�ևt{�]�hz��җ�t<3Ϣ��{�����[���J��yr�f���{ӟl��4�	�J�1[�b%�myO�ld}QӆB�3�����b�՝�w�n�P����w�L�I�j�TW(�|�%�9?!S��W"A3㾙���T�����FTΩnl*�r��S��}�X�F!L�{npC�' �&v{���\\Y^���z�W�����Qý>�8Mt�?Ǎʙs����Ձ�0	�k�#k�ײn1�*��ՙ���
���p����Ǧ���E�:�ߺ�\s�4��%��cOEO����s��.�8|q'k�����=e��|�=V��E�;F�fi�x.Nxqt}p^>�w�#.���&�! �,(C�|{U��D3��1">�=���RO�{����Mu�����^/�o*������t��c�="@-j�����ʄp~:����A���^��ݴ~�(��3��xo���xh ����H�����z:){�X;�J^SBٜGN����'l�"f�7�k����K�)����nwyS.u'�\�D:ɇr�u��I��vB:"pV��ǔ���5�*�*`��-ݍ�xԇ���e^�%n�w�'�c(�	J�9�n�U�a�)�_oh�^�H�{w���S����}�/��
��A��O�=�ڶ�faX�%�O�O��=�zۑ��Sy8�q��-��Q��R��x�QJ}a���z�{%z�YG�a�ߩ]ch/z���k�3��g�T��*�H��V��Æ�Ʋs���D��ѓW{{>Q:��`v���2�(5B�?p��&Ur�����x���B/yiR�a�FK+P���:)�3*7T�O��IX�ptCȰ"�Br�u7z׼��K��7���M�@4z��Ͻ�T��t���Q\�a)���FX��:FAn=C��MBZmǱY#�y�W����Ch��oǼ-:����l��u�= ��*��a�����|,9�~-�,������l��Պ_�&mOt�uS�t�p�k��w���lg�{���R�	TS�Z���5w��ꋚ��FzG�>c���MנX��qу��%:��t�7�ˤ�gW�� e���yrj}�'�/{��dY��Q�܅<�����Εb�+xᨐ�'lb�S���L��`���j��7�u�S�1�P/v�A?��]��p��g�Nl����#`��􋵻�֤u����I�ӓ�M��ﴚ��*�(�އ�S1"�c���պ2��u�4�y�T/�h�4h���v�v�r�;����`�sm�o-H��7��n��cx��>��^�CG)N�����}�l��YjN��%mc*�*uh�)x��X��3�x�0!G=I׮��y�ns�#��NZ��c�{5@�����)*Jc�pCݎZ�3i�;u��'�6���OvNS���nu5Vۏ�hN�&U�us"� �٨��C�ڠ���uyW�x���?L��s�kh,5�~k��+x�@�o��i�� ��(���Rx�x+9x��]ơv��ֱZ�bF/�#r�Z�0��}
��8-zRu�v7�t`X�9��<'jI�\j�U�O1.�:������7���쿘]��D�����{����J�~J��+�>�*3�yuF��-<2�}��]�J<������։�[� =�W����'ˣb����u�]����"�p�c0'Av�Er���~�<<��x-�Gܨ��ˣ�U�"^z(`s��zm��q"s��k	�4��8��`o�������3�lW1�ח��k�{�Z���}��!kD�y�P�>�ϧ��q�_J�1��E�N��|ke�P��2��HU^Nw_�O=�VV<)��3�"��`ذ˰�V.�־����A`��">�s�^	���Ѫ����F��
�k�T�赫Zw.�,�/�f���4���G��k��Xo���4�g��gOs�Q�Vo�y�Q��^fkqy�V���_v]uS�]X�ûo��p}|�)�s��v� ��׊E�[�ST��̷R�+n몿|>� �?==���k�oA_���h��A����������׾c�����9�}`��n^T�G^����4�#0|5Y�!��t}�X����B�qUv�{��N�eZ����Ow���H����Qu�@�/"�V�+�J�Bb�yw��	c�E�g�r�/@��/�É�+�iyv����Ŝ18>�C9������)�-UC�A�1Q�|C�lB��r�87K�����]_�J~����a�(V	5�\/-�|fEd%�?����V�����%�􋮔VT���c-�^K��V��1�
��ŝ6�~4�5%N90Jr-ãJ��s_EŮ�<�eP�����xN><g���G�;�8�C��k��0�{�'7�Z﫞V�9��v�Ǻ��:]q���&�R�I�ZD�#��(/�mC�]"{�6��9AU���� }�ִs��U	[�w�a����>�����{ó�"GU�!d}P(xk��$N.4�7J �rzC烵/Ink�quEQ~�/)׺���PMȵ����L+ Ј�M�bݪ���W>r�坰�2Rq;�p���.�zy��&���+�FX��J0�MŏU�em17��¨8���j�8��T�dص&�6�fwq��\�8��ˎ��MK��-���%jܮ8�Mv�޾��%�R-kY�=':vZ��e� �*Z�TF���A����C�m?�1���g���_\p��6;������H��A�Ŧ��:E��Ck}�M��9����d�()�X���'6E��ް��c��e�	`��cr��e]�]vH�5X+N���fJ�4p�����r���ٳ�G���7�R{a�v�@�N9������d���1�7T��p�*u��!��#ʵQ�����[8���!19>�?R��uwFkY��7H@��.���9V䭑�%&(!E�Aw�Lp2��eL��|#��_�G	MW�s�"�:��B6��^)+|#HZ�-�@U�� R%p���_PpECcڠu�חo���Z�U�������mRBSPԐ����[X2C����3�r�*�p<��|ks�gi�V.r�G{��aq���@��ɜ��
p��UV�jvA�}㽌�+�`�r����-O��f{"�E��~�̓�E<#�Y�}q[r��0��f�&��0Q�)��gS�ב]��r�6�݉�
�OE�h�����pjP��hS��	���dԵ4Uk��~����4�Z�S}��&GQ�\�-K�r� �p�BmI���7��K���}�z��>�ܮī���r!O�R�3���
R~��^����z��>̽�h�������:ۼ��K�qL]��K���I�3��G�[�d�\��n�|;��?� �	��\����;�����">���}�Þ@�"BZ{��NH��Z�c����ư�W�n3��ji{˼� ��?,4Q�~-��bG����v�sj+ �.S](���y�x�ɐ9�����k4�N���� S�c���A�8D��>]�������'!���Y�!�v1�1 =����}��/��:?
Y�m�H�`@��|�4����w
���3e��s
}cU�_�zӐtB7�0�����Q�| H�z�N�k��>�_���ry��;xW�����;t+X4�����֎��{��54�V�>��(XO$0�x�`���KRk��}s�&����^����$DX�^}��}J��2��3��.��6(X��<��:=�_E?�&⋻�[O�tAҗ�����p�z�D�Yb/}z~�(���R^�����U�UK�2}�H�]87�sۇ�h��lU��:k���Ogv�8R��iO��*e��+��yޘ�[߸�l��6J�]�u
�K��y�bw�����si�����\H��l�s�fQ'Þ�����<kX�˺��Gթ�PTߓ����=B��#������N}sfN��z��xM)6aE��(��e�����y���3��7�G9��VwumF.�sҪ��*[r�L�u�w���A �9��X������C��^]xC��EÜS�HB�ҩ����xc>��γ��'�5�.'t�OLV���yз���ڶ���EM��Υ��nJ��(��9t����
m��O����C0��ظ���t~@T�|�G���@�����M	٩�Q0�c{l��3���6}#�e趱+��ZÝ�S�R3�*��rc4��L�F�Ey���3��5�������.�3�L���7&8!Ԡ5�����\v��uH�f:}V���*l�CS���6��f��_:Н(M��}uB�]S�K���&:�t�	pU��[������3QJq�����ˑ�
����4�a���!ǀ����(��Y�2��wu�:hr3�+7�:Di�B�O:��yz'�H�l>�	�S����}u�oӕ&�=E{�ޕ3��6QB��oc*�xb��@j!���W�g�<#W��|
��\���[^��y�?}�U���4�1��*���(�*o`������kK�b4�>����;�w���9��p�Κ���*LR��>��{�o<��;���y�b��O�� =�ek �7u=�A�=�5=��y��f��3]a�C��� sԖ>�<��o�����:J��fnM�C�%7o:v��_5�n��V�0�m�cy�Y�h݂l����pi�}�¨�A�=||����k��mZ���s�hrfu�+�(I�a��_�����s��c����^���Å�/�`Q#2����N��>Ф�؜�rE�M�8?�D���Б\j�*�y�d�o�83o7atb�R8�&~�vc�v�����������G�;�����u�;�
~�q.:s�+a7�x��I��D�;�j|Ȯ���l_ȫ�t�	?{,�N�t��/"Ȯ�fLgNup�E�g�ok����y����3����g�ٿb�a�w���Y2pΛ��f�s��r��t�Ħ`ɟ�����rj*���9��c�����^ʈ����P�}�n� �����G��*��ڑ����'�(�]�r!�;9���w��S����zt�q1�v��)��!V�:>��OqN�aP���9Wڂc����Ӿ6Y�`����q<y�Ac���}U�Ƶˁ��/��d/3`�GeFJ�k���P�[�M]GU^�<E	�ؤ{>�,DT)��8�F�F���{$���}JU3j�ÁQ�{�b�Q7*��S�%�q`�nZ�Ŭ���|��PH^�O�S�@�5˼w�����J7�����VP�vv'�5���n�(���-j�|@�8ك���V��.��2�A-�yu��4�v7��u\�d�@;��:̌ve��A~���{��E>
�|_��T<���<0�R��Q���{����s�S��r.!V�6�������Jn���r�P��C���wl&0<#`c�Av�H�:b�3�N�;.�K���m�7��}�Ώ��?M��`_փ��g�_�5�֫�.0:'-O��0�h]�o��%NN���ǐ���hJ��N U��u�����	@`��}�����v�dzꫳ��W��� 2��]��	�Ӷ9y���o����:�U�A�)_����a���g��5���C�����P����h���>��H��Y��+���������wC����ޕ(��
�ڗN\��-��7��jϛ�`j֋��fn�O��}�;���l�yv��n�Jv1�aV��N��>z�qя�{��4���,���>���5w��C�}�s�~�^��y�5C��B˰��R��:#�Q��ؒ�H��Bw,-��_�ȇ�Jy�}i���sJ<��D�Ø����������K�֛W_�%f��<q��=N&��<�0��@:�K�s�����ι�G�M�%'�ry��i	�f�J����5!J��
+�/:��Co�1v��tX�竪���\Ļ�g�"g;L�L�hwA���0��zlm�j����W�c	_���%�� � ��{[�ݡƿc�Y�����*�噰������-Y�%r�T�!0�n^�h���.��]=g_�F���z�!zm�_^��k�
�ܝN�ѱ8X�c�ޱ��k\-���g��ZPhn�s>���ٴPIXX,w�<!��8S�A��KB�Y(9޳28ڶ�S����>�`�݉���ÓS}�7L���p
�Ɂv"�/|k�?�����.�@�S�g�:{��V� ��������m9�Gy���'h�[�$F��B�+Þ�kk�KL�������oV����3�oZ�����u�i�$M��ră�ɥf�"GP��6*Z�.���ʥR���|F���D��7Q��k4T�{?�D�x���
x,�oz��T�ֳٜ�O�xy�Nb�Ǭk��>�2'HR����[�i|�LJ��!}1�X�6ַ8ۓ@�=�KHY����gL5�ڙ:�H�++#�x��H�Q@���ciB<�`y�\��5e<�?�� �ep���s��Rև�ޱ��N�ƭNS"L/�� ��� ���q��\;o"�2��Ž�Ud�DQ�T���L�3�U�	Y�i8����V�v]Y�0�e��n>��.��5q�}�q�Z��'q�o��B"�����.�I�9Av'Z�Nt|��\�Y��[�*|�n�}|0�2��WCk�B"�i����t室Mt��'���*v��+�L��{���׵Ս�@+�`����j*Wrn�M
��4{ynД�F��U�F՜�j����:�~{��+����,�a����bˣ�\�*i��#7���Wĸ:�$�R�U-���fs��p蔦�²�ѩ��Z��FWv�6�;g�i[�Xw5n`�e�v�7��y&��}`ߛ�j�n�$�j��]DN��	@܋/n��g)n�*vX�v��+��XԦV\Xwoi��[K3t.�&3v-�2�+t&!6�t���FӠt7���<�/�2�p�[��U����Th����kB�
�ʜ��JB@����vw�ۭ��c�,�F���8ќ�Ha�Y�y[J�U��B�{�iY�&�(QW���GRab�U��X`�H�Z��J�@1�m�gb�p���ޡDi�0)Gg>	�pѳ�@��m�5�/��eP�(�.�M-(�I��� ��-��S��w����fj��0���y�8˰:���R���]�7�z��m=y�l�m]hC�\Ԯ�ށ��O�ϻ��@=:����UI�w]o�l�j�X��6R�è�6�������ۻ8ZZ:#"+31!����;��}W�sY��Ԛ6=ʷ;�oM�
����v��j�dھ�����V�Nʋp�2���-@��\�>�Si����2�G:��Z�}�ʽ!��\n=�͎^��z�{d\Cw��=nVr�m��h�V��G{�u,콢/k�óu%#4{%��2��q�4«z��|֫�ٺ�G�k�$"P�՗��1T�sh��)����+v�_<DM53_9t\��]�h_9�&�Y;$[ju��qU��^�8�@�)���V�w��I&����v�]^�Nh�<rec#��Wv)��개!��­��Q~�V� ��Ҡ��D��)�ӱUq���҅-i�J�4c�8K�nc��x�u5�������^ܶ���׀ܽQlabs���3[�''B��C�QJ�*TX�O��z�3W��&<�9�0իӆ��7�-s�y�)�w�h�AU���J�6�9�u��Jz����*�]�HD]έ�Ů����Gq�Ao-C�s;�|qa	�M�L�&��L}�qK��mep�&��8+/Z�S�;3��;ɇ����_U�Xa��W\��l�5�x��ۺ3���	G9>Yt�;���Sѷ�����I����������;�B��/.��jy���H ��E��Ex2�E����H��K6B��6��\=&����F�� j���$*:���ʆ�R0�t�S@��C�y�R�5i�Q�Up�\�	��y�2��I������%�wD��y�k�9ڸ!i�6	�[KC��>�ON����?������[�����=unI]��n&'��v���^�{{{|;goooo������Yl�Ko��,����+-�+�KI		��i���������O*�"BKS�Y�b�ܺk�\�/uӞ��p�fb
 ��Ç�8p��}q�(��..vK����]ݵ̘��;����y�n�k����ow�W����}wPg�����Bcr-��u���\����esy�W����:��κ.|sЋ�K�ܷ5^}j�5>n'u���׺�=.�;ql���wt��0N��]7w.ݻ{���v��7��˝F�4\�鋓�I�|��_]�HX"��7\���\	D"�(�Qf�v�EƼ���fu'�]��Q���=��J��@�u@+�=ڏ �q��v�8!��R�@bhZ�V�R� Ы�k�o���2��~�~1��-)K��z��=�d� �a�ž��hSk�U����_���4 [����B�|���`|7ڰZ���aۈ�O�T��H�͗�����l}�ѮZ��'c�������8=� ��k�P/�g�q*��2�p}v|<�5RR3�T�o)D{� ��$�b�#�R�������91$iz&�I�A=Ξ��+���p}o�i����p�_U��y�l�+�	u�+�DsY⭕��o�y�K�]{p�4Aq�piʁʣ��5/ح-�<
�>~x1ӳFO+��'`c탃����Uf��=G��ۢ~�a�J��t�����P޵��	J��)5a_�M(Pf+g�]�1����1�N����c��}V&�ٰe)CܣE��b���!�֮�"��R���� �Q`F���j&�3?H ��G�gC��y^��楖�E�L����>��	��M��(vc���Oyv�<z�1~�D꟒��j����E�Mh=�xں�"їwu��K���w��GO�t��6��j����(L���x;�ѣ�vǹ��o9�8��nbhh���zuv�v��.�@ǒ�K|ne`�C�ډ����ON�g�������v��h����W>C%n�@��9yբƶ�g'�#�'v�\��/}<h{mE�:8���ӱNz�b�o_e�o��]�	8Oڵ�%� �!2����ι0�y�
������ŗ�Y2�>�����n.;ئ/�w���I�p��Tt@_9x(��ڭؒU�\�����+g���2�����xc�e}*D�ǍH�;�#�%����!��L}��^jGf��[�yf��y�X!��A����2��b�h�ƭ,�WI���j҃�YR|)|����T0�j�x��-�����c�ƽִ5�����	H�T�F-xf��6=��
��|�Ry�;߿}���F	���g"��n��Wx_`kD����ܕ"b���T�w}���<>�|�{X�F�X��M����4�.���a����>�q[�Ƈe��d�O�Ŧ3��ߝ���n8e�	W�h���m��w�}�|j�U:>�K���~�ٻ��{�Ѵv�:�'���T���>��s���96�\{��ې��"?ryX��]�T�;:�f��U�+�	I�SezB����}��.�K�E|��$�@���7"�C����� �gAֺwZogX|�`sZ�Ώ+����0�)ݨŤ�l�vw�sv}�>��O����@�_"�s�ծ!���֫�m��N�	��\=�ɐw>N>^����J��F���w�L͘�8��m6KZ�߯�8���2}���]���_N�T�:%gW�FǴ-�aP�h�=�[N�>�,k�7
9D�����{]�5��y�Ҹy����צ�}�p��~M+��%'��*�D�\L��N���ф�\`�1�R�T�آz����Sٱ��JQ<Eg/\d����t���M��>�q�@Ɉ��+�+�y=mҁ~SQ.�R���r�R���>�]��CҁM�@du������~��ѵ1�k����\����A�bf�]|,�vD���A�w���G��t~�~�|T�v�Қ������A�{ǆ�$&-
��ƿ.eͦ���}�}���K{>�Jƍ������H��w��3�_ˆ��_)�Ҝ��*L�H�vd�^ iJ�^��{"Σ�P�����Sa��]�h��s=������v!�����������e{]��2&�Q}���7ӻ�J<M�_a�
<ň:��|n�����x�l��=�*j�g���{�x��A �@�~���;�Q���pB@��3��@�z+}k6��/���?19��v}�E�N`93��YjWp�(P��`���;���k���l��T�׾:�G�B)"od8�����/�OX�~=����v�)�K��� n��}�ƽL�`Y#�J��a.����-��&�M4:��ۼ��_:���ʴx���?�����^���Bnܵ^~�|v]��}�z��n������5|�)��\Y��M_Jk�8
x���9����EO�FI�����En��c�)�!�/y}�n0�M���]�-y!�:B��V.��5v�ۣ�(Wk&~��P}�GP��������>�^φ��j��\��3�s��O���@�~���4����ͯ��b;`:x�Au��&��ԊS��wn��r��ư�4�'��h��ٳ���oۧ{���k��먖gp�k�+&�jy���s�����sl�IyO���ܡ�WE��.���#+�ڻ{�t�g&�����N�$���Yg�I�p_=�A��ʋ�����A�^2#���W���i�b�\ኜ�\�*�sr��sv�u�`H�D2��I�N$Y��f��/��A��XK7���㲈e%�'"����?'�3��=��A[!؜�_ݑ>�P��e���y)�[��pã2>B���u���~�*A;�y���s-P��+ć��®q�]�K�g�}�������1?�zm�=H��<��ODǥT��g'q�#�{P�t��(��LKŔ�x<=8qx� }��9���7�=~�J��D��}�%��5��xvLX�Ӣi��kS(h�k��+{�sC�=K;�r�hW.�/���p��U#n� �C�|�y�{�ǐ��S�9��s�w(�py��c��B����_���^>�ftۓ|��Ë�����m��SӬq]�-�F1�VU�Q
�$���;��5\p)�^�+�s�e?wI��MZԾȕ��1�4H��}K=��r͔��؇�&���9�
��6v."g�X������rӍBr1�f��o{��y�����8�yh�����0`���e�Ņ<�cHg	@+( ��$��������te_< �#���1���5�}8ivL�-�F�L1�1��8"�/�K;�;eE�tN2)J����26�_�߾ ��(M�=Y�F:+#�?G����%X�/.W�n[������9��s)/d���Y��zs�ކR`��W��fW��p����C��4w�ʄ\z-\�%���ɥ��O��+��/�2����@�F�#���nIT��u��)79��Շ`h�^�t�O<h3X��d��+�Ѿ�������\�w�.����6O�����gŗ�Y*��u��])�.����[��]^
��#�g��y|G�a��ܒ�s���s���������^Vu��	�B��|�z6N<ψA(p��P����9�M�}Yݬ�'�Q�������V��JV=�+l��=K�<|v;�<��;�15���o�F�
6d�"3�J����W�T0�����1�_�܏x��u�جi�[�"4Wew���4��8��ѕ�ro�^P������y�5dA�":��~���EӼV�o]>&�l�vk�[��{�*�v7�l�Hl�����S�����3b!�|^��>��/C���<�E9�('�\B�2:��V���ծ�LjA@�ܽ�Sh�J�L�էz
̍��XH� �A~N�Wd�DA`��,
��os���Ռ��yD'>۶��uG{(�PyKRe�Q����;���߭�O�X,=�S�*�c;���sǇ�@���*�����-{C��Z�x��UkEq�}��^y��K:���/%fƀ��������� ���q��<��d���=�Eh�����ֆ�u�������U���y�O�{;{^l�5��� ��*��}���6�Ц���f�J�)�B�L�ݯ���2����4>q|��Y� ��}HU=�c��{�"�ͫ�[�e侭��a��ٽ���}�1���~��T0z��`g=ԯ��5�t���O���7뼯m��Fk[���Âw�"���a>廙�e�a�o����e���}Js	1vN��M1Y��Io��`j�G8�ٴ�K��?D:��Ô�ET��N���2�i]w-<k]���$�#����:i�.�l�1����D��Y2`�֣�[r�g9���)lVbo;.�L%�V�x��R����z���WI握-�fV芉a.�[M�}�/�]O�����B�}ޝ9�+��{����ߺR��j�p{��}P߮�+�G5�W}�_�����p\����=x[?�Kc�^{F�Y��q��.�u�CMO��K�D�!d���I��y���s~�5;�4�F�1�%�`�F{`vy�׊�����P�z����4m�5~䊅�zD?Mn��;�����/h��R`y��d���L��i�-��Nm��PV�]q��S/�l����ZK�r6X�ޥ$
9X�u�45�CVޱ9KR��[�^���^yD+ �:�oa,k]�׷�,,�`D*����xEta�}��|�/�����0���?�v
��=�O�g%^ac�}�$������s��%�G�6 Bxb��2���Ό�[��Y�b&rf�Y���&0�1�X���������m_�i)���Ɉ���jg����;ʈ�ʨ�c�s2P����:L�ӉwZu3sTa�����z��}���F����!܌v����.)SjT᭚��W��+Z��\���".&7���'�e$n=F��|B(3_*�h�M�;�j�Y�F��Yn�D�ˈ�$�`��e
��?� ��u�>g<l	����W�V�'���W`�o�x�l�/��"~�t�{����[�Ho�8�v�R:���;>��X���������6�]a~���v��y;ޡȌu�n>��'H��'�f��/�2-��FǏ��d��g+�����ڤ�,�_�YF��y�j�O[��*j�=u�g;*���J�0/�{�`❌}ư����t����E�]�����_%#S��Pu��xr��?O۸q؞��y��������ȧ�S�u�˷�;�/�#i���?P=θP~�[Y�p=K��"O����~�"��t��1�և����!Ă���ڻi���N��flo�(5{�8�͸��4�!���=��'a�4�c��}Q:P��Bi� ef���C0�p��ko�3�p�~�EX�J��9`���~0+iq<W�cys��������w��ڍMإ(`��L�'/���OU+�y{_iGZ�x�p�������a�
�7{6�D�H=_A��a0����22
�|�rs�Rm�Ӧ4�=o�x!Wݛ�d���z��;����k�Z��X�&v<E�fR����vs���@���n�������������O͜P6�-20�����v�
�V����&��]�"DL	�ϛ����ͤ���	T�`l�}8�h�������lz{\>hh�~��mxm���C��^>wa�ఋ�K��{o�.����8��lHA�:[t�a�M��쏽�!���%u��=5ý���r�(���v:Ƕ�C3$R�ꏃ���=wa��Ю�3�h�/q1�h�S�=3i��G��\��G����cX��Y5Ai�����4Vf�e�(��-��u�����O��5��A��z�Y��P�߽^�Ys��/ˏ=�š�1:X��@q�;Z�J3X�c|J�q��04C�-\��w5��{Q�6D�-�����S��b/3�OY*��}��eK�38ه�eي^��|�pˀ}�J�s�v���\�����IR�WT��6�;�&K�-�F���^�1VJ�5�Y�.i����]���=Jh�\Rgw/��+����l�}(� �P����j��B�QX�S��)�y\�A�u]���:J�㨖b��]Y��L�v��4f�B^Y�D7�,�� �Q�k5�9���{m�����YB����7|�2^q�ݔ��e��Nd+z�h+���q��+XA]�mc�����8�+J�����yzN��C�E�y�Ld����F���,�]�m��s5*}C�J��hHs���%k�Ҷ��̍��=���$�k}ڠ#�({¯�� ,�%bߗT	^ӆj�Eؑ�_`ۺ��
׷]w1��*<�3-��\�m۩F�q��W��|4U�{���<�ޓ���8,�У��FKt��8 '�W�;�v�f��ꎬ;��TU����m ���9՚	��XhB�9ls):�T����r
3)�i��:�P��BY}�{�ޔK��1�Vwj�t��,Q�Y����QL3lgL*d��K������!�s�l˜������V[QP�Kch$(��V}����s��um�"F��;gY'��Ůk��]h��1j�:b's�$��}�*�@�SV�ˇ5^���)�]�q�ݍ��Ud	j�ܡ �;��c���f�슔�ޘk^Q+3��.�vy:�IV�T�4�Պ������1�ɝ�6��2VÆKgr�7,X˵4��:�aN:�k�Y��]���i�a�+�����O�]AwČ~C6�@Rzֆ���j.�;�Z�oKʙ��fR2g7�%h�\r��k��$�ش,H xM�9b��f�O��}x��١<o�����;lu!�;����dc1K��t���Y�Q�|ţ ���&���Xr��=w��8����a��s.SOs.�J���ظ�"�L쾊�=;v���G,W�-����ѷ��o��/UK1:Ӽ@�=;�;��q��|�EB,څ�:4(�z��1k�.��8�M�v�+X��"��bڸ֎ԼKb�(���3�����(L�V�V�̺��n.S�kE �CcRp�M����nfW�	hG�b�}.p�Ό���Q
CkWwf@G[0:R\�݄�.�
juyh��SG��g^c�K�8]�slP2aM����K�/Pc��gN0�[�}�i<t�G�����ö �Yf�qo,��e�<H�$
:י��_Δ�N�}G�	��gR�x�E��miGue�݂�Ɣ%@A���π�s��wM:wY���g:.�v�	YP���mOYFe�������DMv�P��;�:�c�>��wÛ��{&WJ��.d�݋nظ�uA�+�U��kWKH�D��K�;U��C/lc-�[�Ћ�l�}��������	 �ᱫyM�2������E�wY[v�Ǐ&�3TF���$��	��)�)��ݾ���S���t[��Ð�<}��|u����׷�����|������R�8rI$��9t���u滺�Gv��Nq���J���k����ooooo�oooo��� O-��!e���^s����K�g���es���E��.��;�ws��ׅ �8p���8 �� @����3$���䯟7�����wGN��D0�B���8xa��i�������������Xyi	#%��<�&(z[�Ww;�DV���w2���ϧ�����J��#�]�f^u�ss����2r�9���	\���4�����׾���\�wGwtQ;��h������9Ӏ�V��{�w�׺/>w{�t����E��LQ}7���;�7wn�'w+�ޛԗ9}�>�_Ca)��r7u�;�D0\� B0;����ۜ��ws9�"�Wu�:�w]�OU�'��&�4����B\�P�t�s���+���HR�AH���j���lPc��o%{���k�^Jm�j��Guf��0ʙ7kX�h�NH��f&�^��F� {���� ���g�eg���\G�E��C6N���E��5�/���>����d�L��hC�K�����v����s�kl��y�ϖ�D]����T&�����x߉-�_����O�I9���Nb��NQ��˿�~��ay��9����M��)�K�#%5��՛ݟH�ɡ�G��(��ءl�ӓ'aYYY��KF�ăA�*�5ԡ��f���9�U�7mg�
K��U�[E�V}��Io��c�&��(l���}^�<;W��>��=�_��}Aq�)w�m��V��9�1=w���$ ����x̈�H�^L�����.13ݨr��!����|��=�J�޸̪wR׬U�W�<��뙀#WGJ����w�>d?����~!�'�;�s�{�ʬ�~�<܋I$������_���==kv�R5�+��q|m��4ם-"��;�m��M�7L ��~\�^�E�M:/9m6!���"��V>�rO-�HJ��\��7J�e�G�vb��#˪�p�g
����>�;*��3�Ԣ/�zk�J�BT֏}{}�p���}��::Bl�\'fՈ�|q*=�U8�iU�~�|~ ��]�{�`���';}F�a�ǀIQ_q�Η�=��a���>�^�s���{vu;Z��}�<�(xJ��u����粕�u�a]7�>|��2mc�Q��鷊u� ����w�UǪ��gX���2��'�y�6���nvM�����3�I]��k"~>�e������*�qX*��⭷q�'�=�v�G/��Z)�2n�|����9���Q��.��Bn�_L_��گp�����|�>�x7�����i\�(�������2"�nH��~N���L5���<�8J�m.�xa���\�	�|��y�S]�
�'�:bCW6�ekw�g;�V=�`£�;��6�3�{||�r�􊟩q�%ߪ%	cd������.��gF�1I�7 S�����ۗ��ל���Mf㾬�c��ָ��k*B��h����7����wS1H[y8�nI4��uv�f�����W�!n��
?Q���x�N�B<���ލ�Ӄ
?(\��SGm<<�D��aޥ"��#����3���1���c.H�yw�����gG��LD��kT�H �SD�}�a�Pmo�����B� ��j������C1 u�B=�c	%�6��׷z�
�i^����R��W��G�s�y~�<��X~J>a���S0#��,��o%`p��X�������+ǅ�)�����g���(,*�MRc�f׳*��˯~����Q5�����0-؍��}�S�Pҍ��p�"S�����C��i�Lj�3�c���d�[�[����C�@���UBh�x��D�ٝ�yVWS��oz�r+����G��{�]�=�p�!���|�GU=��5~���<ᮼl�0�3��u��s�zϭ�0hF�a�J�.cq;9~��K�؂��Ο��ۈ9t��[U3����L`����|��#����Y}s���{p�I��*���^2�{�`S���"�,o/��
�+9N�F+����9F��4y�\T���]���t�wA���"s.�Ҳ�h�1
��#��u��_d�����u:�2��_n�A;�5=�R��D�%mAX5ur�=[C�F�E&�e5��vv����"وbw&}:k�����2��SL��v��bޕɗ���@�r5S��[Yˍ�x���-�xxxP�B��ѫ��Xc�&h���~FjO=E��5m}���&L���uǬee�>�mzO�[�����8���S��'�!�ts�-���ʏ�;�}6;�O�H-'Vu�A�v
3_.��*��<�V�s�wD�﫶�4I&�͊�����k��^�͡C�E _��Ʌ��4*��C�p{?cƵ>�9����_?���{kT|WJ������� ���s�3���T�0����=S�n3��r��=�`��i��2�U�yӭ{�z��Q�$��}���(p�!_G@KX���}��C��^�EF�O�x���Y�ب��fZ������g�ʻȔ���ئ�	Т��Lhjr��sժ�ΏV���\�����Zy���`��cd6��5��a�S�d a��ODUD<�}�E��lͫl���w+�����U�~�Eu�._�Ƞj.4B&�!N���Hy
W:���3�ʚ�`�[�5]��Ew.{��#�o�=�|z���5{�5v�2^��Ʋ�[�Y���ܡd`�f��6�&*乑��Fe�ovR��JW֒ˈj�c�U٪���|(��cɬ��3�*�Z3�u'��lNF�}b�h�S�HW(��Cl�Z#�����f�Eg�=]���+J���PN��]}�f�fA�M�L�q��ؾO�vb�!TZ�����L� F��!ݛUM�G�Q��ŗ�Y*��۪�Fc5���vR��͎n�Ď�Ǻ���&pQ�_@��Jw�֗T�T+��w���ɏ{�kc"f=_v���X�}}�]�$!Ƅ�:����!�Oyo�d�/	h#Y�U�OQ�տh_`�dF�82���%�<��ɨxR](��v�
��������}�A�KE.f�`zn[����lK����+��.�$|~��s�=yx+���M�A��������Uo��#٧�����}>cߦ�E��~_�~:��s��kޕ��U��I{G4y�w(�z���+�Y�W�����v�
�@_��4�ʲb�DMVw���G$�1F�wW������V��FP�;���@�]���Ҳ*E��X��t�<<�`?�I� E�A���үq.�}۟J���6�qS�7����0����}�D��\	�M�3g>dp�[[DC:>=������|>("-a>
����k���v3q���iY:�Ά��Z�����w�2��c�p�G�sx/����׾�������mx.ݱ���6%��թ���swzY�zB��5^���E���¾T��r�#'����j�'���=v���|��j6��51XS��Zo~�R=�5����V�Oi�Z�7F8�����7��>�$�M�݂�t4�*6#�u�˶�3k_��{��k�[R��!<��|�FO��"~�����Vu�Ӹk�Ú�{=��L�Y�ǳωw�Aj�tp�@~��b��'}�7Y}{���Mvή$��Jlb�Gq���������������;qT;Y�x���Ι+��u>-��2��y*�}n{���r�M�M��m<#V��#��0۱<�G{��z>���k�쮣�tA\n��s8m��?,�f{/��q�h�s�6c�_pWb�u��2m������8��7��oy�b���=��DEX�٤֔�ZZ�כ'�u����s��~�uj��*3�ror�t��9�̫˘��u7>�}�s�T��P�:�(�Lu:,Hh�*?j���}��� ���ݚ���9&s���1G�f���X���+�v��p&�8�i=��4��~�ֻ�E�����C�;��	��w�z>�@/�'\\�����Hu�K�����v�Z_�^�X����3h p�c	-��m`�7���OZ~�3\���|�$GH�Қ��'>^��U�f7�]]�목�������Şc{s높��;�����^�=��i�eYC%ػD�+�i�͚�[��X{ೢU�|2�h2��0���_#�X��F�.6F��b�G�+�3ϴҝ)W
u�G�_;����G�O���3�3w4/�2}q�ź�Z�ϣ�^I��@�R�n[N�=���-�3H���1�f)��X�:mT��L���ϴ�y�|žٲ����[����oc���,�Ǟ͗����Pӽܾ3�`�%��>Lg��5��~�A���������y� ��)n�kQ8�Uŋ!�#�E�X5��M��]1칁�|����v:�/V�Ö1�s�4w�BS67c��*r�C�r�w����F��Ύ���}�Yv�'��ͬ�7%���;��l#�d��m��V퇶���9�<Ju ?���;7�$�旯���e�+|�LV��_���&�>��Y�Rʽ��"o�-�U	�UY9��'s�7I�~�iLH��ip���q�w��Y�1@ܡ+�g�E;����}ż^+_e������s(USo�N!:�3��7�va���]v⧠Or�y�|Q8�L�|�^�ҋU���U�m|<m�8#��|�7��5�_E������Ku����N��nO�?=b�dOp�#y�V+.��'��xpQm����<�o�Jw=�6%��Բ���[��� WJ\1X9
�Q,*?_Q����6n�ULn������61���5�DP����l���]��E�g���(�Xl�ݿ��{�.�zߚ=�m���n�:=t�� yIfS�X��d`N��Y��lm�[���~�Q���l��u������+���ڛ�!8�gb^�Ǐj���}2�]�����oh��R�����8}��=kx����@v��Q�<7}V��W��u��Ѯ$�82Q�8����u��7z�9�ڢt����.�H/,���>��xxP�Z6������g��.���P{CE(��m��;�GQ�3�����g����X�[~��Q狷|�m^lHat}NVئ��#v�S����8{U�(�ֻ���,��Z)�w֪�ݟy��/���c[{m�K���0�x>Z��/9�G�[(z�~��~�޺��`[~����<d��H �پjo�ϪAD#O�m���\��	��e��l��j�����x}�����6=*����x,R�ϮX%Tw�U�;x5�Xd���${՞���G�z���l��'�,�T�YT݊F���oo)9H�e��gu�}�wU�0w��e}�B�p�`�D{�p�+�G�s�_3u���9$�����������#�{7�<X��E�1P�DL���վ���~�,�����H��]^=�|�b�~�#�u1dZ���\�}�7|���s�2*sn�J�c/��}}e���]b���L�Xٷ������q�Y4w�d}]B�/��3����,�s����}p�=Z�_x����9�՝���z�^5�}:��%�2}�R)Е:4軍�Q�ݢH9�|@?A�EǶ���^�ַ��B,���&�֖
��ϔJ"<H�Z+���̬�$���<�&���>�^9~��2�|7�o�5!(£S{Nb3ڜ�G\�<����9�7�ª�U3��8+2�oz��e}��!/��@8�b��I��*ce��q���I$�ڥ<eO�G�&�]�2z�^q���#���1���8-��X<C��'�m���<���!ȍ��5S�PU�ꃏ�E��/_�>Y}�8�}���O��۹W+Fo�|>aL�C�x=�Ǒ���b���Kt����AX�L�I�i����������+׳�xg�9v��B���C�YP�B��m��M9�K��o�Z�$+�F�.�Z�A�#2U�	�-�}���a��
�;����Pʶ��D:�uN�����Z�{���f��p�Ro}Q"!��}Qy���'����`�P�&n\\�qg̡����a}�2���٦���5�l]"df|���^�&ȶ�M�#�8�*}��V��{��%�*������\�=wݕe:��Q���|6]u�7�fd\B2b�oK����Q[��6M5�v�Խ��8;�s�Gjbݜ�%׼��\�Q�֝�.��E��������)FN����;�t��n���:�k�
t��yY2)�֩S
��Ӳ�	Ѵ�nu���n�#Z��$�S���IL��˙�.�]׮����N�VٗY������!k�̑��c���F+;մz��V�6Z����m�o��Q�ZZ����ǧ9ޅ���á2Q�֨��t���O�Ǣ�;oMy�)J� "0�������a�zw)\������J�cUu��k�w͌AR��/9��\�,V�B�Μ�3ֈ��3��i�c(��%:��MN��V̜zN���-U�\\ԂCzD��)|(�wN�\mm��D4���Q�H���R�7�z����ި��KMa����ᡫ< ��jܠ�c��3;��,�*7.���\Ժ�h +Vo���3(0�.*��dL��o�̽��Q�7�,�}�*�;��P{�h�\����*�<ӧ�U-���FL�gV瀈7l�n-�;��I�J��բ���n��ls/���(W,�SqCV��1�}�j�w1���Z�CH�-�kk�i��R�w'P�]k��JU�E�O/.�>��BF�A1��׺��R���� �����z�q��r����X�v�o��ޗ���Dթ"ta�˫�츩��aK]ӕ.叫z��Wؚ��ټ��w}�NK�Li0%�����0
�f�Z9N���*��+7�y,��δc�.]-���=��k��Rs�ЏzBkD��L<�w\�*�<9�i�pnޮ����>��#����u��da��Q��;�����]�>_�F�k	I ������M��h%��b;��e�2���n+��\��j��4�}ƺS�1��	�[R�vh�w�=+X��o<��)Ұ���o �P}�d�Dq1�����5��z6�O��8��$9}4�7��Z.<'\B�v.�|�5����W�9W`V���+/8MM=un5m<��ںk�e�w�p����>U��MqOX�ҠK�n�0P�3�v+(���/��٨�7�b�p�v�GH�wi	��@��ܪa�0*U0,pdd�m�ιd诓ƶ��%Bh�}]�I����:Gt6QI��8��T.����pZ�}���K�3.�Y��y�k�(d��,ɂ����
Bjۼ(�Q9}B����f'�VU�Cd=�9���g/ի'�ӕw�y���"�����vrն�z�m�S5�T���X"
���ĢBR>�FeU� �LP�� ��4,�2�if�eP)���b(�Pd��7�I!F�v@��A �h�ԆT�`,($U�,�<	DQT�:%��߯�tt��qγwwv�wt�nr�rw��A�]�����v�Ӣ\�;��/7���^>8���������t��~>5��<����ciK-�����Z��!nҾ�z�d�ns	78&D��ww:�6�����7��Mzzzzz}�==:����({K����b���rc����E.݊�̺e�a�����$���/.�"�ܑ3�B�xxxxhC���mH�]�i%���p�&Y7s����|�cy�!\�;��wr�K������ܸ" @���#����B ��_�]ΗIws.#��r뷗ӛ����I.��^0���\{��{�8��剜����bM�'����F�t�t�$�깓;�&�û�a��wq�s�o��|�s!�Lw'wA΄g.K�M"8�\Lr�����]�]�L����u�g�\�P�����t��s�wa��4wII�w]׽\^��wE�"���0�)������\��9ӻ�)B�rI�������wq��뛻�����u�n�b"�tl��;�L�Bd�u��t�3Nk��}��ܹ4�s��]q؈l�p�,�s�0�wQ4A,�Z7�S��U�+��w�e��gt��n�0�R�8W12��ڏ^*Vď�&R@<��2�ΊI�.�i�څ:$QL�T	=���� �f�-�R^���8Da���*�Sm%�A�������^���J�0vN{	Cj��-�4�?*�������7�虘��_�!��J�2�g�+�ע0�%�G�i����
��'<��>��ʧ�]m����{���n�}�c'6�{Hy�Ѧ/��Ձ<�;�<8���|�ފ����cD��ym%���'����X<��=����I�٧)�2��{k�8�'r��18�v�D�bXf���U�X+��Ѳ3���m��ۘ��z�R�z�28"zO��Ќ�,B�#������bɺ� C����W>��uv�]�~���e��xf���L�z�lP
���y1'��݌�Qأs�޼�$�Z9b�r��=�-���ZX�6�B��w�4��嚫��-GvOLp�ݻ����̪Ex%j����-|)y}�>�Ƌ���?%������i;�T�X�L��2d�J4��B��&\����Ou+YN�ኘ�� ����G����~��#��\�Ԗ��\C�b�ۡj\�\"���!7����˔��P͙�Lu������.҈���U~�|>(P�����*>�]��9C=�����~�ЁES/�ݷ�9n/N�����=���f��/�Uc6&�p�Hp�{���Z޿�u#�ҍ?G����.�Oz�vg��04ӵ'inK�ߝ��BPu~�=���v�<�f�C#��mw�����M����P�zk��ú�}K2U��0Vmc�cO.�G]�P�v�y�\V2�9��<}L��#zW���n�{�Q�Ã4�͊�����]��o�)�L�>g�AO�c��gV���<=�/.���ɋ�H���0}�=�E�.�Sw��fj���pT_|�sAÃ�SӞ"|�1�+�_���H�B�G�#��[�����h]#Y[���D�9���Zh��c�`�ﳾ�A��W�ص���OTI���}g8�앧�ЎV�A��k�؍�[��V���deu�x��\85bW8�je�
�z�cޝ�,��rr�^3�eݻ����W	����f�]�
�Xݪ�4d���*�=��D�mfj\sm��;u=���:ި�2%�:ڍS��ثrA�J�H�Գ�&
�Iy$��w�蛨���_xxxxP�@{�t��yi^7��3�X��9p(���Z<D�aT�;���p�}b���vq��{ٮsp׹.m
����z��Y/y�D���T��0�92�C��^Н��C�{;ǩ���������k)ΪF���k����[E�}OB��k��� �fQ��xz���W����++�\��}5u;��f�>9*��ӡȝ~]�k��ȫ��{_h� \�Z���V1�m~{(��������<�S�|��j�Թ�V��Ʈ}l�<��Oo�}��ДCj��2j��z���ہ���KE6�QY�w_{%����M���܎>�9WNO�|��N�7L*�@����J�/枎�M��=��;��s���ŗ;]��3�+�hQ*莡��;�8�oYx8�+@��kRnb��ޮ���S^�B��Q�C=J�o��A�����#�X��/�R`v�z���D���F�����è=���a��l���.��/�����/�U�2|~�<��Uf���<:��;zv%��{[�۱��֔�6[���Z�2f�ũ��m�	�<V'��)�.�����DL�nK��ˎ~]y�6͌�G��'Rv)yd>H�et�ll+��E<��;x^�s���$��=��$!>���#ݰ���׹ࢌ=�#�%������#p�:Q\w��c�l��7�p�bG�qٯP���F�z�I�)=�<=�	@Zf��g!�便b@�V�l�P�th��������l/u��ӂ�U�$^��KBW��P}a#�E�͝凰�S\�tsۂ�Vw0VkX<=?f���`4�8�x��FK��)���=������X%Ġ���N7uygY�?q^ӓ�.��eI��m�U	_��5��j	%���ɡ�	Ϙn����Rvn�z�T_��
��q�zz��+�}�₿��:=9��co%_\Hc�k�w�i��}�����/.6�<+��y���4�韩�X]��r��d����&f+�"�����fZ��e�
��0N���r��ie��2������U{����;xK	����
��=J������)�r�9wn.n�j�Y�p��S���bG�ʝ�7�z���eh/e3�ú
�"��Y�3qu%��he���`a�s9o/8a�8I���~ @^ח��f3� �D��6���+9�B���k)9���y�4�S�T�V]'�p��Ff`�l��Op��:�\i��uW{�ۆ�;�w��|Q����n^��+{�p����f���_aQ��_�F���"��Ә�;d�uYW�q�F��f����GZ���ֿC.*ꮬ|�K�{Ε��L���d��HsPo�>��:��B؉��e���E
�De��s�ʵ��U���Vg�57��J�嬫����D�
���>�7�}k8a#�[H��j�{��O�&�[v������[�ԯ��\�������z����ڎ~���{�V�G����rOn�7�e?��f��=�>���'�Hz���3��{������V�6��Fo=��8�0�\	C|��±� ��������}�ʼ�$����ݿ�'�I�S�u��+�Ws�M��&�m����pl�\g�
���8�1"*��=��8�a�]94,urk��y��@�F��$56
��
�D%�u�9H�-�=�/���t��^L��yŽ����3�#�hq�_W�[��?��� �s�'PZJ����
��|(b��>Q,L��jCS�6�[�L6������<*&<�|���ņ�
�;��ܫ�Ƃ%�8T�x����>��}���/
_Gj�}N�r�}��4�im�G����xf�_����#�ȕ�$� 82F�<ϛ[����~��X�ZQz��Ӣ�t�{ۇ!��~�b�����D��Y~z2��|U��ͻ��o�-�4f��-�+���ls�W�()r�����_�@���������|˛՜�ϐ?^�y~���O6�d���{�~���$<�z����ܤs}�uG����J�z��2�&dX��qxY�@�~�׫}ܫ���W7��z�KZ3ҭ���M����k���2c������K��>�[�5lv�LF�%����]u�������X�O�F�����%��d�&z�.g�*��˦E��XY`Æ�|�7���gWL�훭���ٻ����uD}�Ŧ�A�x�<�K:��L��Q�|X��c�`�z⭵m�k��Ko:Iګݵ٘�	OU��nV��!��(����e�N�V��5iHp��~�V���p��?]��z#�k�eX��W�=�3�T�1�՛p:�M_nx)ޣc�2Ǟ�bGp���c��W]����]L�*�d�o�v��g��{݇4�b�P^�_ՇI��>�����ޟ��}Itv�p���m�^�B6s�>>���VU�"U�te.2���v"d�&�R��94�$�?[}y���z��k�q�VQ��+����*��3~�����"{%��|.bQsx�i��5~�srr����ua	����w���ٞ�,ê��N�X+6�g���:g�xF5��fz�B�U9�8<�ٌ^;����Pߒ���^��w^]cE� �~�?_��]��F���= ������;C*�+�=Ѣ�P8Z�����+$�w��[�x����@���%+�xړ������/"C
��X(N/�|;|��e��;7ʹ$�(�eJ����k��M#���y����IƷ�G˴(yeѿI/��T�dޭaD:�o+��C�y]@�z����X=w{���Ԙ\����5�ެ[�e֤��MrQmիC�r�`����B���|�5�=�w��}���J%���(��z���0n}^�~�o�OE���_������r�hΰ��w
T���6[(m����N�P�a-���sb�1i}s�o�ݰ)�T�g`2�U>Lt�	nܻ��n{K�NS�O��(7��T�?H|� ��L��V�����n�LM��Mg�>��%.2��I�xu�~�|}T��8�I5�>���{|��=�����I��U���E���E���}�3���=��6��{�5<s�}�?W�L�z��>(�{��C������p0rc�~�df/k4�?�$a�r���|�#{����z��԰BTemxHx�=��Jr���b�#����D,��7�Ũ���~�C�ʧу�o��4`p�|�;̐�{�h�!>�O�k�lZ����yKf���?L�vi���((����B���� "�X��]3&wP����;��<�A5ז�W{��!e�����o;Qm��PQ�ٗdZ��i 	����&�hݵ�$�̃6��yc��JZ�.8�*<y�f[��gQU�F�����{㘐�pIIR�PT  ��n9"�i2$����B�
�<�����}��*
��a���ro�1*�+b<c�Lh7��ߎ�]��1�d����@��W!|�q�f篖���Џ��~���V�vXS�<�~��D��~ZJs��m���Ÿ���Ͻ>�~��W�\@�1��z�1�Vq�
��k>(qy���S����k>�}a���䧞�=S~1�eRgyiW&�Ê�zW�C��9�A_ة�*�o~��B�6�$U^��&�x��Gf�r��q'�����
�_)�X+)��U�����r�%א}{�d������'�lF�J
s�����£�^�ۋ�b�i�o9��4�qd���Eo�{�9�Q�#w}�o0|cN�C8򽨼N�s�O&	�1�T��zxߟ��1 ��e���}j��>��M(%�}����v��sI_W3c[���^x��/5{� � R��	��2~� 㕃4}��s|j1��l���L: ��7�ڴ@g4�_vc*޳��!�w��I�Y����n�tǴzPN��Hz���)׳+v�w۽�A]w:���=�Uy%Y�����8�T��̌�ѳ#h��S��-09�U5����A��n/M|��;�g�炩T��-����j�jr��42�fϴ�Mfg��=�������������
��j9�v�O}CvFw;{��ύ�R�0O_ò8'>b�	�V(=�!X�`���q^��;�_���R�w������4��1!��j%���T��gN��^+ ���1��P���?\3���8:�Ё2ĪK�����{�PEq4�C�v���[�Y��14�����^ed�Tk�ށ,V*f���Y�� D @%|�Lfj�N��m2݌6�KZez;ݬz��t�_=��{=���y������О�C��گ����L+�=���������w�G�ߐ����}"���G������_}�<o�dO�M%=%��Ɏ�x�t���v��k>���{v�=����{q�/�ޯ}^\?Lh9�#��O՚��s;�d�k^�W��G��n��;����n�^��-WT( y�o��i.��4]�D�ȸ]��ߣ���}X1J�qŖ�yӝ�:Sv`�O��q8k��N}��';
�$��{�����7]�	*g/��Q�7��n���{:��C3�ǫ=%M�"s�󒌙W	��8�K0��e��x*ʢ�%{,�=�n���k�I4��a�s�Q��`gq��Rڕ��A�V���{���͌�_���k|EA٧׊�;A��❦��cgl�yW��v ��*�m�9_9n@u��FI�9��a�U�#����V�V��rX'm�1�kU�f��ڈ��B
Nhr�Y�v�����J$�h\M��l���g[��[� I��^%�ug�K$ෝ7�OL� �\[�,j��:F�m�5>�V��.�+�<�*q�{�vu}�4���xw�x�c;A[VlGo�O���fK�ux�ҳǡ�i�1�1�bj��j���: /m����C[ʙ����RX�hIKwQ�hwgX��0���c��°ֵ��k�݇��'r vѽ3���uS�=ɭ�s61��3��t��ڄZ3���ޏ�w5�;eC\����h[����\��7��k�$OS[��b���:��Xw��(����w�����WQl�^���;���hr"��Q�!cls���Nĥ���yŮ4E#��oN�ʽ5�(���)8���L�3Q��� y=��]�N��⣝D�ܸ�v�A���%�\�rue����ǯ	8�:&��v;��>t�\��in<��htQ���oE�W;zj �����I���B�Em�,�շ�&���1^܀i��m��]Ue��4�yՂ��
�@��"3@{adՈ�aa�	$Ƈ�Y��?3^��==.�^��ef�I��Tr�$ަbRdG�`��X�{Y�����\{(vv÷0��U��p2$2�L�)�Yҥ蓦l�n�P��=o�?A�t�Ʀk"��!R��n��!f��&q�o��@o�5r���O�$�|W7eO.���l��7�6��Yx9G]��d��un��wq�r]�51b"B���Tv̙S@,&v�74*v�������7��w:u���<7+��
��%�m]K�z�E��5��xV�\�RF�Ӳ�Z�|�u`׊���fU��O�ZF���w���SL�d'�/���ҭ�'Tr��r����׹V9	,�]��ݸM�Q��:�\�O ���)����RJu�i[Ħ���N��&�1cgv6�M"���j�
W�b�x������#��ϴ�w)<���	��?ꏗp�l�`�.�O-��d`���Wb�
}dֶؘ��,oq�*�4n��qѕW(eq�9�p1�K6���je����y��Dt��w#������t�V��h���T���6.�����v�5�&��ƂX�T�N���p��Z��'�;�ΜZK_|^]����<��m��8>&�"z����zt�f�I�qZ++[:�ũ
��(���I �I$�A'���$1�����B�D���L ��L"D$#�Ò�XƼq���{zzzzz~==:���2�"BC�JJXY��ܝܗu�n���$�� ȆK�����t)�C)l������`���O�^������ӯ�~y!�
I뤈3"�v	!�bQ�3�܂���`F�_����ttttt{<:<<<�BB@`y�Er�$�np���3Bow&Lu�b0��}<D ���0!�<<<<<4!�B�)$	|q{���w1�A.�K9qܗ.ۻ�Gs�;�ݿ�]tџ?;Đ����?W��%���қ���Hf�@�:����:2�rQd_���EJ�k�~���1H�!�S^�pp����+��M0�{�����F�d�c�˜�s�]��H�we4��� wn����ٔ9���ޜ�wur�������˗���4K��&;�wqsE��WӅ�ۇ%ˊLX6�{N��٠IB0�@�B�bw	Qf���y�h<�f篈���x��oR�ɾ7��轸>�6�w��ԩ���'�a�s��j����|(P�^O�������7������ۿWz�>�d衊>����C�~��q�n�n�W��Q��q�ޙ��߮l�\�|�G�xz6���w\���z�%ﳽ��B�ӡu��d����q����OoW+�"�N@����ڵkp�[;�?@}�[��6}��V~�\��dN�g>����Nk'�a�Vfq��T]4s6��� �y+'��h���ݯ���rǴa�l�ٽ�gb/T<>�Sq��^z�"!�EvK������/;�_!�� �����$�����O������؎k��_��.�����<'��4D��9漻ҋt�j��D���D߸q�R�z����@��+��*��r���}G�8r�F�鋼7������N=�ϚG�O�q_�+�r(ϗ�X/#�WY�U��֏}���`k�Y�D�þwd7SZ�o�3�n�rM��]�	�s9կS��
J/5�h�yyD6�
�0��;r�/��ͅjC�N/��IpѾ�������;'
u;ڶ��_=,ܞ���O���$�v��/�z��A�-�nL����z�:��-����s���:�Y�I ����¨P�#�;�Ω5�4yU#9<Ȁ4:���F�����n��m?$sJ^R��hE�i{�����w�ͮ�{.�7 ߄�Y���=75��P����Q[��xx.?T��Qט"=+{�����E���U�X(W� ?0���i���*F��Mv�uE���yf��|d���I�z�B�G��h�N�H�:sF>��ͳ]�~�bpʯxo�=ko/P��>ѹ��KEhSMbmؔVgӺ�w�].���ףk]MS�gt�i��dq;b�y�o��e��O~3j�(oeS4`u�U_���ɮ����N��� ��JfP��,+{�b=���9Q�s����"G���~Ĕ��z��ً���!��h}���؍/�<��^��*v�z{ҽ��$M�2��q��m`���?w�K�I��넺�i@���Fݮ$|�`E�a��-�[�n:�j����L9�j�����LS��Ye�T�
�,Y��zs��ߟ]�5��jmv�1��*�]uUr�}�"5j :�Ҏ�QP�d�/^z�.�����u�8�\�#�&�����+��\ͮ�j�N���p�&�3ˣ��s�R��y�P;6��K�%əs%9s��d��1�B�Z��%/I=">��ؘ��4�v��|�$�|���+�1�E�h>��r�w�����OLo_����C�4$5R;([+y��Y�9��Ӈ�y���{��jk�F /�O��hi���s����V� '��w�Ӭ��Wk4x�{��Y璾f�M�?p��E=^�ּ=�ܞ]Qfe�����1F��ŚаQ��xgB���J�-���G����pvv��Uy�}�p���{��a�׬4�f���
��0�I��z}�l����{Oq�{Y��}��ɿw��+{��l�,m�ED�@=��qt��#���=5�!�z��=�H����w���ϭv�mFv����K��詉���o6'���m}���3ϯ� ��T� U�ڋ�ZH�v��]�9��F����[Q�B�&��Mz��oJ4����l�ھ����{z^:ꇚg5Q�J�\52�(��E�w�}Z	�a|����|�s�����X��p}V�|mн.���Xga �Ž*)�C�J�Q9Ҹ,���Lޭ�7�Jkoa��g�~��Ȧ�âCR]Qe}��>��r>މ*����޵Sف�{���S������ϲ�x\ڽ�y�j��y珦�B�1[_w����zfՇ���}
:�c��쫧���|�i�#��ݦtϾ��o��}���-°��LLL����'�$ֆ�eAUE��\��.D�ؤs�O��_���䵕q��!{��5�|��ͨCG���T��;^wT���-��VU4R���WG*�G�r�g���r��!�����]�T�����y�������g�	���V����8�p̗�����M�������Q�o����K�;��I�k�����1�ǼxY�pD��S��
���Щ�׹����;+Z?��|�ӌ
�{?W�.*#�|�:�M����uP����E�u>���^�#�d���\�}yf�|�oZ��o~_^WoY7�/�+O�8Z=�^�"�Z١�Z�ӌ����@9�0�p��yi-�Y�V8D�09�.�6v�+B�Q�E9���@{��7���7-�r7��P<�}u� 7��s���<���P��ǚr	�$���^yQ���-Y��[`��� /�|~?A��w�����-�cQ�̗��D�?�icY�k��
{�U^�c�z� A��{�x���_��`�F������^^�̠��paY�T�;iG<�=��I�κ{�����g%��CkE-����g��P}�{%ژ)47�"���6ݼ�g3�۶<�]��A8_f
i<�U��4#m繊�vDw��!w���t��K\�ō��d���r]�-�Z}�}���=��3����M^��V�`��R0�E�X8�#��ζ��S�3�ڷ����p�~��|)�`C��|�wXX�����u\��	Pr�f�%�k�O7�9�\=���@|3R�o et@s�V)���w{w?��~�Û�,{(��zכ��$w������"���b����8�]'���V�]`����S��ߏ��0m?���Z�C�G���ӻMe����8w81[�4�����Jո-N=��n��� ��.����mOa����P��֛���J*Zꅫ��;����c����c����w���	*3��Ro}�x��X�B���K�V�Y�<* ¹"cvѩ����{�?%?a����G����Wh�_���D��=�!�U��I'ݯ�lPj�-�o�A�U�G�9�$�{�~�(@���~��=����d�}���{Y!�I��]탱~�_`J��T(ς�a�e_��]�tU���Sg��u8:߬!�SI��7���p�Xo~Br2LE��\y(��=�g::7`Rb��U0��	�jm�_����DչW1�'�4����#�k�[����ꚏG�Ժ6
�T��2��{rz�wV�չr�W�9ש�}��w�6��l�9���ށ�� ������;j��s�ao�`}ǋ�S���Fa�scl�����M,4U"�{��7�y ���'D�m�s���;،��އ�<$E�RI\�?5��i6�q�;����������r��Fr�:����6�� �;�l�����y֨��� �]�!̤�+�v��j�NDi�I2*t��Ɍ��`��ݪ��&���JhWnl�I��u��ӭ�=��Ց	d������+'r� ��	[��,�t�f���{X��<[ym<��6f���
��4�T:��t�++&�È*#�g6��tJ	U�I3��Y�R�����l�߿y�r�8l�z9*�ete����o��}�q��^��;��T�{&�:���Dz}���j��ػ��a?h��w}}��ϡ�z�oy�Ľ`iJlbƓ$��]������j4&���QQ��寗w�M��� �X7����uN�s���7I�{��W�ۨ�y��oã�,���L�%_ܹ�O䶩�8>��r�u�Ϡ˺�%�O#��{��A�xW���"��,����9�{��s�2��/a��Y5f�=c�!�" `ǐ�|&��� 'X2��'��~�o}�Cuڹ��t��Z[��q}v#��/�uD��p�SM��o}�<<����|�;1�Y���thXZ)�R�e{w�3���7&�İ�U1���~��xo�d��|�i#ˍ{���o�g5�b�q`z��e����~x�2�g�O���{���;��۰R6�($n��WA膨m�;fcf��f��=��C��]��1P�ٕ�aw����Ƹ�ZUY��v7�4O{;�I�5���]�ν���N#7���n�Ԟe��-�#����z���3��F��g��'hn���T������?iʟmθ��`��]{(O{;kx�`ҁ��~���^�V�y��ܫ���;�~����`��.����m���=�A���L��"uxM���[qD�;�Ltv!��w�iz�GۂR��(/�LQR��D����)�ǯ3�|��9�V�ʩ��Vh��k�)��
��H*��Ǔ��r�e�tC�Fǽ���Y�f�E<~�q�.�/�������&��Y��7�S?s���f�J�o[*���q[�ֻt{_p�9��MD��.�Uc���Ǫ,���J�X�Fι�~§�8��ұ�A���]bz��CsDg��O[zQ�9Z��ޯ��A��z)%:�3�W՚�M��kYz�*���*�^t.�'��h��8��}~s�O�k�qoɚ+�ٚ�{x��Ϊ>;�
����&�C�Ϩw�W�'��������IM%���P��]�>D�vnf�]{pPW���֩s�� e��k-�2���)7Mш�ٗ�|�|ﬥ��*��SUv�[��*��t��Q[��n���
�=�^�=u��%��������ݯ��Y ����@��/j��+��,o���h����^1#��A���Ф;��9�0Ng�<��k���ؗ�A7�;8��xY��'������k���7qf}�����˵H��_��wj��4T$}'�������������-��e���G/�=�m?
#|���E���?5�!��C7��
w�������]{Sf[	w)c%��	�[F���n���X����A�7���B�{���Ʈt��o���C�����d�m]�u��<��s���cך�ã�l�̞�{Y��[�v�h�×���vǣ�*dD���\)����!<�H��%m&�)����o�z��+�`C6�o����/ˮ�a])M�>攩9&�yc�!�Z&Ô��p��i�vh(1޺�_4�M�Z qYܬ�_��)��
�;��Ǹ�~_>SK:>���2��>oM�OFU����S�k��������lp�5��,��bnq�.撪�AJ�\�9I��P�w���i�m�$�T��$6IIyA"�D�}D��)ӯ l�w[��$��<  *�eP��٘c�'��\�m�l;��.!ԵV���Wp�+���-���[ٳ�,RbǷ0n� t�K�ݓg+V	0}�y��L#p0��|v����#��B�ț޲荅����E�o�E�J�`������4�G1?0���3a��z� �菧;��G\-�z*��J3��BPu0x�p��m��%���ljYS>{J��n�ˌ��kǟ�崼/DH�g��勸�Fӧ���#�!�8��Нxnܝ��ꄯ�cg�g�`��X'�x-��WԽ���#��@��Z��6t�s�|�n�}�-S����Ʒ�j�ݗG�o�
���V��~w�]N߰�6I��pz�Ԃ�C�/���x{#����XT-ٹ�[;=1c4����QT`z�c����BT<4��v&��l�������2�t��%s����\�t�>�CɎ檻�}�w�{H�id�
��|��G���ƻx+	a�
��|�h�z�	T�Y���?����~����Q[�` �������  �;�������=���[�,�d�ii��M%�-6Դ�e��1�m��kLl�Ҵզf"jҥI���ږ��-*��-��ֲ�[R�-i�ڙ�5ib�m-+l�Kjd�Mm1��m��5iiV�[L�M)+ih��kLb%���KU2�5��&MZX�Ui��[iQ6Ա֙4��KFf�������kLd��KKZc%5�b%Vc5�ZU��m-)mLl�R���)��6j�&)���k1���ٵ�I-��-��[f6m���֚�i�1�kf6m����j�KYim��M�ZU�l�������RKYik-6��)[1��V��ҶZj�J�iU-5�Ҭ���KYik+MYi�����VZme�Yim���<�>����$Q �e �A$�QV�@ �P	@ �	 2�T$ �A$ZU���j�i����کi����j�{կj�KKj�i�����R�[U--����T��U--���P�J���H�T�֪���R�mU-5j���T������W��ת���T�MZZmR�U-+R�Z�����������HA )��[iiV������D���P�8	�	$A �ZV��V�٫KKZcf�1�ڻ�]���m�f��Ll��ҵ*%����Ɖ�KKZcD���}/���?O����" �� 
F'�����Wο�������O����������������	Oؖ�����{���E�g���C���~� WޱE������� 1�S�E���~��C���(���_���?�� ���N��?�?�N������)'���V��kI�K5����Z*�ٵK6��Z��Rʴ�m�6�m)Z�ZҳV�ښ[R��K5i�Zj��ԫK6���jSZ�j�m�ieZm5�m���V��Զ�֚͵%�*V��5i�mSi�KMjZ�ږmSeTԵ���ҚԦ�%�*��l�K*�-���J�je�)V�����i�Ij��%Y���Zŵ��f��5���-X�͖�[����P� DD4��[\�V�V�j�6�jѵ�*��ZJ�b֍j-�%��5ZJ�ٵF��%�6mSRڍ�l�ԴUT�p����/����  
2((����
�� ��:����~��H�� �t����QEh~�����}��tП��`�8��������0�_�(����CS�����'pEE�Q_�C� ���iD^}�<�EE����J��'����@�п��>���~8 �EV~�?�������+��I �����������?H >�'����!��EW���~���(�������CD��ÿ�p���;O��?/�xv�D���="(���{� ����@���~@��K��7��(������O�B" ������O�~��q�?�b��L���q��V� � ���fO� �w���յY��56�6�mm�*�*�ʉH�m�+Z�ٴ�Z5�j���խ� ��i�6Q�U�kU"���Գe&���"ƚ���Mm�ٱ�k	kiX�����f�	W�:��k)�m�9�-��m��d�ц�lbm���&l�A�J�ƙ��%����m��6Vf��h���F��m��lجUU�{��Z�7QK�Z&f6n��v؆�j6ڕSTҫ5�m��f���[kF��	m�Zٱ�`��5��SZ�eT��%WH�mV�ڍib�͉��;�ƚ]w+}��  x���.�4]����{޷N,ݯOm����v�n�n�v�r��a�^�v���ޝ��G��븺�m�
���nJWY�5��N�gnպ���=׽��^�%Ef��Yjkk5�b�� �nB�CB�w���B�ؑCC��}��xz(P�B�{���nϯ�J۶�=�P{j�����i�fiҽ���j�ǭ{X�oqg�ͼ���iר;�շ���V�=Zf����U�(��f�k*�b��]d�� ��_.¶`.��z�{u�խ��N��k��쮽�'�6�m*h�m�{ON��m�<�Sݴ����w[Z����WCW�wu��.����5����W��`��M�KSQ6�T�X���-� n��Mt �N�qQ�l��s�v�{:�ݶv�eP=����������z�4�K
 wgrw=4�z�r�b5l͡Y{j�)_  [�hУ�Э6�;vWU�}�^����u��(�*ptu]�f��۱v��*�\����6FT�:m�M2�ڕ�w]�,�USj�e�|  ����v�[�EWB��k��W��p�P�����t�����Ӷ�CZ�ӱ��-w��UzttS���TP׼���h��[��Z��Z�h�[�  \��n���� P�i�  "�h ��  ]�8  �ہ�A@7;\ 
�t� ŀ  �vi��X���l�Rfv::�� ��  ՞�  �� nf�P q�  ng  �5� 3N��48�} o<����]kU���&�Z�m����*��  �� ���]�  ������� �n�  6�g  up  �8  ��
 h�;�4 �nb��(�wr]�V�5V��$[�  w^z( �,( ۭ� :  �+���` Q�F  �Շ@ d� �Bd�� �S�)JT ���ђR�   OɈJRTb0 �b)�CIJT   Dޠ4�T3"`�BRBx��� ����O��~�_iL���H��oZvq��Ec�N���n=Vk��6CG�o3y��o{�n�����_�EUE?� ����A�1DVUTS�����g7/����)�fּ�ٶ����n���փ���/Z�i<I��P�̔���5�ƈ�j[7ESL%�E�W�#e�ܺ�1x$:d�Vآr��4��7��Nn\�d��f��Zh6j^�c a<���R���v2���5�13��.�L#C#�+hfh��7��M8�6� ���O j�ջ�.�f����rS����)�-G�b�����TteXW�O*��tv�m����*{��:�䭔��r�EFղ��B隗���4hc�KU�ܘ���0�##�0K;H6%31��#�v��Ol%������U���"��z/�3��W,[' ��w�O���F��(�gpVRV�B�P�[��	%�KT0[��
ݤ�<f����x&Ju;��iJr �=�M͘�ӻ2�w��8������c�R��K���Kn	���i��ʂ�m�G�b��qNe`z7v���4Z�6E2jX&,V`t�<��Hּ��k1Yxc"�����7�2��{���ͣyWaQ��N] �i�	pf�&�܌f'��b��!BG�)ܭv�9ek2�VEh�+c�{���6�x��6�;p�C)�iQ�gAH�+� �t�B�����f�V����6������{j��o��H���bQz/o4ij�L��S�)�m=��J٨��M�v�&ԌU�t-M!i�+j1�B�k5��0]t��{��4�Ml`ۙ����1;8�7a��In�ܕ$�@�P�6^QL��r�E�%�AL&R�e�\�^���yJˤ&Zp\��J��4�2�2u:���ڟ=�a�(�l�RV��15�@����޽�Qcm��5#�KAfX˷{�5.��v�6vʋQ�4���V�
����d���
�Z�T��ԜN�a��Z�*P@�:9�U"�:�N+)^ �K�3];c&����XN<�v6�6����H��?�����ě�2�<ؐj� MX�m�FA�:^B&&�8��K�_D.�V��sVbU7E�V=Y�T�M(5�e^���ǐ��P�N=[d�s�05�̙`�Z�2�#�&�]��2�h�M o�m�Ay���q2������ʸ�8@�d��KSF�B���/"O"HV�`�hXߜ8�j��P,ܧ[��LR��G+c0�����=�$0I��ËU�V#[1�L�L���5B�ґ�k�p���Ug�ΦٽP���*,�"�t7, �#s5�lFm���Ӎ��$rݩtԧM�s*
ʴf�h3$Yb֭�o쥶��V*(.��cB��ժ�-�AZw���Z������25�-�H�qքV�'P
�S f��*�0c�p3�tL���
�ɔ��
����c�J��^:E�ݍ&��|���e���XTM��z��3R�[�A��C��i[![�C䩘�n�:���+q3x]:DMk��@Z�tN T�+v����Ь8^�!�X1�:��q��r�^����e\�OMY׻�اA⎛%[��E
,��;����n�����C������hbr0�Ō(��bmZ�b�/�ј���t��T�X�
R�D��6�؁t����wS�(M��,��jA�AA�t�p*�]���7��;w���(V�F��:F�@��^���Q�y"�YYR�N����8#�wX�*G��EP���&f� �>�-�*i.�B�R"X���V9p�{nc�,f
�6̖+E��65�(�7 �x����@��`O.d�`3�0D�y���hc��]e
���Xm�aS�d���Hc)�R�[{��k#6�pB��3M0U^�uՐ��n]�Me��u*n�n�Df=Pd��8��CpM���ys\
�`Zdr��v�w��e
��X�Ky�U�Zͻ���.J�9qD�^+ �7b���3b�r(��#d3x�Fkvk��L�8˸w�W��:JC5G��7��µ摌���1m6�qK�A �RO<�W���/5Ro+M��u���!b�_��
�@ɲH7n�Mǩe*�x�ǭ�lظ�E*�-�M*�.��c�PӤ��ov0dt/c�ז`D��K�ŷ����8x�=�B���3�LqB]fF^G�5��H�*�04*��A����3\��'��fNJ5v�<��"[��$/�)D���T�iVn��ncg#52�wfR��+2�.Х�S(ee6�Bh�.�J�P��ں۽�f���b{���p��L�6��mX�6Kɖ�7N�hP��k���e�U��L���!�P�rB�²���4��J��U2d��`v�?�6&,l�۵W(�ӛ
`��D�ci�0����_�fe�y�>���m���9%
�5�%B�n�n�6�Q!`1ľ��%Xu��^eێ
B�ɛ�h �k*�D��m��;��A���/N7�Of0E&ѽ�5U�=):dR�j���#��ᩡ���#X�M�&���QmZ�%F���D�ܗq�Idң���f\[�}�wm7�c�pk�b���:m����DX�G�L˛y���i�B,�K���s+1:uxF�T!Y[M�C�2d��A��+f@Z$I�Ȉ5�oL+0n�,m��ӡj� �)��<�Bl��W�]4����]��R�ڳb�z9X���5�`T���"�R�N�7�˭�5�K�*%CM�Y�k/	Xeɂ$ݬ�x�f�=�z�:�q#	�Y�T��h�D�6�X&Asl��v�2Ы�yp�NW�;yc%La��E+�%�j*�ճ�ve�ͭc6�)�Cr��fP��E�#(Lg&Q���[J��7Q�K��e"��m��94����B� Q�ږ�'�+JB�r�[�o��m�ַX��U �R��Xwx᫭1�>y�֌��X��dL�B�#��2�u��ek�T~��f̶�XB�g��AQZ�O~d� T�8^͆[2�!�xk,YЂ��,�q�-[��Kn,�ʴ��ӎn$ͪi�6�8l�K�W�ILuo
�Z���ڂ�єv��%�4�����i���rB�J3"Q
ܕ.c�������a��]���ȅ�;�T(�:�FRVtF�Rv��f�3�;gq���%m�)],u+&��l+򙚬Qb���^�$�˺����լ*2$+���*����ܰ�RX��V�H�[��r���#a`�6�܇	QUƮBsj�TC`��Âl`�b�q]�]�֔��(C؅)�%���M��j]嬤���:��e&�m�-Ь��]��r�7l�NG���@�5��g0��J�]I
���ނ�)V[����W$8��軒 7+3+� q�G�%�Q���d�3�1��3�ȗ�L�9E�4p�%
D��&]�1eb�l���6U�ۼJ`�%9WV�Y�w6Զuj��ۦ� �9I�,�T��{��+�M��K�ql�e��Ւ�Cx�wML�E ���]T�J�R�4��dF����h�㊚�j]2�!G[���9�HE�5,26���!+X���P֬���^c������r�[�	��ሒ�0V$�cS.����n�M�5�����g�4ܛyy/E됗N;tJJ7�Yr��,���8�ͻ��i��h���N��uI�UE�uw�I�:DE�,E4�h�8v=�i�Y6�7�JR�w�.#���'J�snh�)	Q[�"�J	�2���˛$tN�d��+�P�"+�N���nV�8�V�h�*�WY�=�7�� �#8�㧅B�۬� ���B�5�f!w6��U*���
E8�YE�wVv�M�Yd��qL��X&��7h�"�-\��Ce^C�����N�7p]3 E�e�.��Ð]�ov4�0�Q�a�t�Xb0�^��h�eJ�y3�[�u�M2�[BM���sA�=VX����X%5�4f�;��z�B鱆ةa���-��v$T.m*�)�3(�b�m��cL��0�Ltʱ���9���@�h�Nr�hTڱ�.]�i�\`2�5�0f�����1�)���oksS�w��m�u
xGَMmE,\�6頕L�t�H�ne+�fnh����H,�)\_S�9��𮾬E���2��ڧ� �Lح�K�*V��H�e]d��1nI�j !��6K4�x��3u� u�r��U�9lZ�iM�����r�Lr��+v����e��*��+�!��gE�3!�S���o\�ن�ók#�y�1�
,w&�6K�k��2���j��>�񷆖��U	��r�2@n�i���e���v�6�\�Z����M|��s ��kvS�CܳM�����u�f��D�,�Ǖuj�����ÏbS5[��Zb�G������v�cW����3re^����"�H�q���e��t*�A���q��jiq��6�$��b��
9���e<�&���3 ��� ���p^L�w��x��	�%УyGrƵV�ˆ��)M!�V=H��bR�Q�IFv2P�v�Ja�x7P��T�fEk0L m����L�m��*��y��2�;6�S�,)
�K�ڽ_�[�����8��K9h������lW�0�.�Ţ�s��S�ll�7F�q����u�܎�e��ݶZ�:*�)��j��6Y���b{��ʕt�1U�������|K���mQkb˲ӄ��,�
����&��雴¹�E�T���x�l��"1،y[��a�� ���ȭ5[��jB��O롔3oD 㲩mb���z����|U���5��d�?r�`ƌ�uvS�)�� 2����)���h��ǏaY�#kLFj�h`�i�����T��f�[v�e騋r^Fkn�2���&�l�vc�~�&��:�5��po�v���aOi��6�t�Y�ULypE�,
Z5Q���"�y6:ؙ�#�ұ� K)�w#�n1���jeՐ̤���K#2�{���̤J�hh42��R�������lJ�n<�����if�ţqm4��Ii:���� l��t�����GVV\#$2���x`2�4�[ڑ%�l�عN���lWI^�XFj�V�02�dys���n[�J:d���e��t�ި1,wm��p�4p�8�c���J��VufeA�ߞc#[�yH��2�VֻqY�u���P*�C��櫴��kHշ,�yp�a��P��p`2]$���J,e�0�L#���,�m�Vm(!+h�Mf'#��Ĵ�{�e��M�W1��gi�Gw�Y� 8ۗ���ͽ�p3r)d=�t ���YF��ȷ���A�[���aĊ�[,"��$�ێ;.a���KK���'XjVIL��,x$�g1�Q���WY)*BK{.[��c3F��\NIY�;�y%D>t��0kjL42gٲL�]��i1)$�7K��RӬ�?�(�h�)X�7(h;���YXlH�ɳpRVX��I@<��1�q�ݐ��RAZ��a�VL�6�W�+K�vN�S�!�R�&րVٿ�nU�B�	�Ïkr*l�o�0C������ً3#�����c*��nm����i���SrZp���@hke�k7û��mn�e�(h�pF���\�"s#�=+m,[�,�"�>J�^T6��gj0.�����X*L�SnAm3�5�G*�f��~*�q*�Hq�S�r�(4̆
��XX��\�3r��@'F��@�B峣5�\nܖs�a�{XY
�͛�0:��E�-���ک��v��O.�J���4�.;�
G� �Z�n�޻N�J�Ա��V�V��7�HL��[��.L<-�VXɌ#wΈUi�Lh��3Cː�֚�sd	�U�u%\uf���S\Ѧ�,Z�s_�VY������Xtkg7��-к+n��$��`��u 	�n��F@q3�>���ں4����3\���^�M�E<wWI����8�B�MD���L��Y�n�u�h�Ŋ�jYZ�Y�3JIpSWgriT�2�j`QMQ� ӏ\��V݆~��ۭɢ���1:�qŢl:h��Ӻ "R�U�#-3D��J��}(,�t����>8r������I9��?��6�L�K�����0��R�ami�6D��N�hX����j�ǂni;rf*&*�f���Ty�"���F���]=�9��:�f,Z٣U/�a�R��Ճ5�	i�FIM�2\t(�k!���0n��]3����bt<d�� �u\t#�*p�b�C��n�����:��f��6��-�1c�V�XGrC�ո��l�W���*(\�nc��*�7N�ɏF�Q�Cp�ux�1a�k)�<��o\�ۈe@���7{1����$�$G���,J,��X��,8��Z
�xI#fx�� Q����d�f%���F�� ۩L@����a�[)��w�(G����iS���/ ���B�P���:�$ȶ�F�JrQ���
U���>L�*�֖�-��[��l;�(^ޣLѫ�bH��i���Ù17���s-�����<�T���\�pE����EC�9%�Kʗ.�������4��(S3n̕`&���	�6�,��U�J�E�"v([�q�<�����̈́K�&�5�a#[!ɉړ(4[�x+t�z�9m��
K[j�٫�nm��M^�ٓy���;i����y�q"r"4|�V@�{�q�I�I,0�,C�#�l��P�ke�YP+��;�v+)Mw��;̘2��Z�5���H���洓���X���5������ڏVZ
�&���N�*ZO�lj�jȡ,�q1f�d���nZԪ2B�j+�iQ�q�ՙ#� .uS)�,��(�-��r*��v�z�pbx��&^Q���6��QqU�l+4�ejj��D�����L�nb�?�΢��3�tﹾz42�{��9��%���c���]<�z����W[}F��wl��]Dm��������|�)C��ٛҚ�Kr��*��we����b�;�l5-�:��m6��>�Qs=�ۨ�B��mwP�9ql��IT+�lּ e��	�%��s���y}A����L���H�z��-|�B��P��C��A��G P��r����nb/�J	�;��F�{�p���u��sg��y]j�*�����obt0�뺊P�V{:L�>ˮ.r�8rOZ)8J↤��sE;-N�	��휌gp���%��환����d��1�7�3�Ճu����J�%s3��I��7�S�v8�a)0/�PcWԡ��Z�H!����U[���� ))�r9F�������K�Z�c�c�|�bjտ;>�:΂�4�EOc��oc����&�̼Cz�	�O�k�ؚ���\2�>g�8�=�@+e�95��v)�ŵDt�^zt|���r���V�fU�k��%r�n�luj�hSif�}���d��ǐGY�{q�w6M 5Ia�V0Öf��3���>�]Җ�V�ӱܞɂ�qt�vq�#OU�[�v�I�c�9d��؞�}��c��룩5���S���!���k������޺C�;���J5�#A�o�H�Qɝ4\�Ȕ�YB��\ȅtȭ�2n�%N�hϜ�̼\��G�\6L±U�+x�z���wN���O��/��\�g9��lY=B:��-��Q�{�S�k쎻�]�wu�|0<��&�1xyE�I�7vTz��l��t_W5�����81;+��@�э�U-���vXI,���Β�+p��A��l��MD��Mf5r���+������n��@]|	�W]k�7�-�Ҹ��\�";{�Ptb�A�N���X���բ�u�m>�E��|5MܢBǗ��#}ҝ�۠w�4̻�.�c$��5n�8�i��zuLtܧE=%Yb�V)��Y�g�Zܮ�sc�򤵳<��.�umMr�a��t>�%ӏ9j��ٙFV9����sQx,��Yj�N56*p32}I[Yv���˳�L�HP&�L�d�L��W���6F-A�fLal�J���-.%�B7�L�*Q9�˨��]_R�q���y.�Ƥ8��8�V�L�ՙ&ۨ*L�%�C˨�ڔ�ɫO�V�/���ݝᒹ;'y��Ѣ"=�����1kY��o.s��Զ�u�J������o�+�Q���S�Y�;�î�yԬ��eK��ֻ��qQ�i�gV5A�;�M(v��Z_�IG'��v��UN�O��H[��\!�5E� �|6b�"�WJl��1�4D��GF@/K1Z��pF��et��d��%ƻ*g���k{���:�YV���1� t�����g��ظ�:d�W�8n汓9[��wT�"��lP�vȖ���n�����hǘ��6iױgX����(��ݵSR���j�ʶ��Y1����}R_8���k���xL�٘��kuД�'��9Wb�)΋Ap�:ʕl�w!���cf)d�Q[�$X�`Y��/��i��wXܵG:��	XD��g^1Ά�R�:�K@֔۬�U�j��t�g�)u*.�m���u��O5XǮ�����nE�:.�`�FC��X�9S�řt�>Cv1�Ϋ}�ms-Ne��/y1��3x�1Y��n�$����1����M������jXKM�vP��7h��'냍0��7�A:�QXgu�����{�O0w�F�f�X2J�sU��k/9?�ĥR����Q-�F�Ū|JYD>,du�u[fe_\�3���Ojϫ��AL�{ggu����r��f��d]�s�{�U��vͩݜ��#����O>��2`�HEV��Y��S��0_iT�V�7��eY���eI������ţn��{3�G�GS#eg�[���]�z|(��+㳮�l��n��J"2D\
��2v�S��S���-lɂ^�Ա�7�����a���W�3�9vK9�ͣo2W �ԩ=�e.=�E�q?��d\h���@��d��jSE� O[�x��,�OI���C�ٛ��[�orM9�xO�[-�����h����s�q#gE�ެĘZX} U{��;��L�M��}˯U(�D�<.�m���.��sɋ(c�P7@�a.m���6�%��xZ{���XS]br�Zn�:�Uj�[��J>�)>0o}ęR!��+VY[6A����WY���)F!E0f�Z�X�]*���أ;y�I��a�qv�;o4�ߧ˫h�Ja��4��"�~���*?"���y^7m�s���`M�.��m���I�N����VE�)Vc�Ò�����B��n��ʘjR�g�ڷ�q/��4 -��3L��,�n�%�ל(G���]v�h��#һ����7�S��1�;��6�s����I�9�d�OQ��u��dd�Z�s�I�ʚ4Ԧ��:�I�p���ݛP9	M�*S+�,��8+TGX����`HJ��$ySi�]Q^wixeIv��;��u�N���a�X���S!T[�V�����eֺS�'[�V�i0�J)LU�Ɉܰ�;�׽���9�eZ�%�"���ᎴP=�87�B�de�5J8�M�Q.A3ZiAL��C��6/fe*[�,|۸s�B�j�/]�fu}��!���+�*�o��$�&;��kwv��t���V�ʒ���;��sZ{V=l����݆&��v�D�������`��	ެ�H�b���z���+�+�]��]���֯����L8fOZ�1�~�m�u�c��;��%�����_,I���[�R��L��O��:��9S"�G� 't�O�f^ز!*��m�+�ew:ֱV�8�u�Ieߋ�%j̣.Dr���sv^�A���%��E��+��+{+/> �x1�w��L�6s�v��w�YO�taVb���x;r���RyW^Fo����U�.�	O�¹�¦�5��;Л<uw	���x;&�������;��ˊ	��{���\r�ϳ�&�}�Z���_S���Ӛ�"�W>qC�yl��v��m�-�͝�V���4����<36�7�ܻ�NM�ދ�K�-�9�v�B�3�+/�����.(��w��r��.��xð�*�[��
]���tf\�m:�k�̵�YG7z�n��3�H�5��.����T����
�rҾ��}_1�����!���F)ev����_)�n�rK% ^����Ͱ�N�ZmfU�<��u�JTb_u��|�n�
@���J���v�ʢ���`=�a��\@S�E�P�]��(�r]������1r��I�o���vH�n��Q�9n���J�G;;��� ��9w�;�*���xmٮ�V㷭�.����� �<d�&��kxcKƅ/��T�%}E�y���IR���^V
��w�mY"pi�O����#�4�[&>��\}%����Z��E@�Xj��Jh3��_N2v"�Q��pƶ�c��$h�鵆b�=;*>�>v�o;C�:�YR�Ԯu��v��Y,;����$0�8BΑPtpWu�b�rA�|n���������T�1*��hkƯ�[q���
�q��6�5�EV�JGfJ�G�n�p�U��J�ەq4i"V��YK�Zw<{:��S�]��`�@�6�n��ׁ�tI���Jt&��"rҩZyL�!m>�Q�g7�u��� \����C��7�	��ǌLf�}�3\�û]պÇmҰ�F^�eh{�+��!U��2��[�Xjk/P���u
�[EN�W.cLg�/���۸b���s��ۖ���\�Ǝ�z�^�:Ŗ/	�� /V	]�ͷנb��D��{ӗ ��s�ax^��aK�*�g���nW�q�B�5H��Ͱ2N���:��oo�L� ;�޳Y*jf5��WR�X�ݕ��Ʌ_U�'y8kː�}A�@��o%@_*���ͣw�m8������<˛��K�*�2��!��͏}�yD8 ��i�.�\�ξ�1)k?;��l�W%+s�)
�[�t�GK-���X�ҫ��+oN��c+�J�4vd������ݺ��X�mj6J��G��{i�S�r��W.��f���z4��'�f��-yA�j
u��������a��=���ͻ�f�㰜��ǈ%��˿�����Ht������^�z���M��3:��
yJ;E�k	4����
�!�W�t+���	y��d;�j*-Pe4�c�t�1I�zG�C�&���<B-�ʤ_T����X\�q�5�n������kf.�ݙV���md������
+�SΗ�|�g>��IFp�]R���Ļ��3&��<�n���9����.�Et|eK�]�;`6�JxEcKD��}���
�ăx��&�V�w:�e]���emE��
�Zas�c}Ue�#ƣ��m�l�%��};o�	��	�����mɲ�R����t���+��Ğ*C����]��B��8�V��g����%�3�݅$vY]�*ubQ�E��D5Y*��7k.	�j:��ɒ��2&pG7���۷�:��Ӟ*Bj�S����ا.�8�Y�����,q��q����5�4�d���*����КS*U�N>���2�Y����9}��VQ]�L��$x�*.֣�q��<+�{g�w��ʗF�N�����<�uwݹ�0����s����n�]P5t`}LV�i��L..n����w�%q��9l�Z�Ce-�-��L�nF�=�.�%qi	Z�2�$�[��9�Z��'*��j������˓e-�����`w9��ײ�|�e�. V��F(�QBg����P��*�C\gf�#�ȷ��v;��%�����+z���ƯXM�W���k��Ӝ���Y�ݵk��t���J��6���j�ڷ���)ʹ�qk�w(̲a��Ŵ����֥���u���o�Y^��V�E�=,V�O�Ѻ*�]��8��j·���+A��@f�{��ݭX0�0̧�P/�
�ҍ�u���4Kn��Sb純��BXDԃ���Wue�5*�b�t_�������#0��I:��b�i���ރY�N=�D��v�G� ie�LЬ6�r��4'j�'ns�t�b�xf��)@�l��m�u��@u�eS��brwE7y���O�r�j�ϩ9�I�m()�=��2W�=���21f+�l��K���@ƾ��]�(��w�i������"I1^>��n�3���f�=շٮR�{�1(�Hx���l�M�\�����:�z�w/w�iR���N�Ŵ버�{�8Kù��˸�G��l��1_m%��]�m�9�)�̙3��߆��}�C��e�i���*<�K� |x�̭7m04ȅJ��W^�m���g�����p݇A�o-3���u��s�����u?F����b�.�j��)��9��������e�Wg&�'ap̽����/G}�>��g9ӷ�텏j� h�
&�:�M"��ԚO<����vN��e�e0E)���lTB�)U�:�3��V�`1m�cܭm��� ���o���}9�������&�
W�H�Pm1Yr��V�wTV7N����9��n��FW;�v���a}Pf�[EjQ ��A�͆X��s� ���x�Ǣ!s�`:󡤍!q�*�M�J�.�a��{5�����.u�n�i��"u�,N��ڎ���f�HD�K QOvQ)��]�8���9��ue	rr�}�,���gSkN�&KJ�n��Ү���˹��������r��݀�����7��ݤ&��!4��H�n}��'�b��w�I0������Wc��O��3�MSOiMSQ�n��c��un�Tܾ����������E��`�iX����zW�H�%�;��])eͮBp8K��K�S�O$��Io��d՛I��)p²�
c��n1�&.��b�ml=�KҔr3'3+&s�-���Pΰ���ܷ�ܾ�ܵ���a]&q�����-��V}�X��n[���?�p�1[ںJ�-c(���9f�W�\�ɤbJ��bC�τ��mƎ�jE5�Uwd�8LI���vQX)�z��֐=���3�TN�F���$�=Y=�j��Z�9u��ՐtU�2B�Ԭl#v���؜ɀ���A��}&��z��0m��y[�;��L_Z��	QF���U�k�K��!]9��FwG(�mNӆc��Ggv^:OB���Gࡒkv�;2��NZ����g�/2`�R[����ʹQk��5}��Kk��/Yo+���{)M�:<·��Ek�h�]g	��]���w���m-0�9�<cwu���ZYWom$/*��G|K��,w��s+6�ө�b�^��]�厗+B�c�g=�0�ɽt�h�)�7��ysh�Yۦ�}ҍ�"��'N��]u$t2�q˴5¸_G&�s�i?+MT.��q��Ӵ�UϻLr�"�;��a[h��Y�:�V)�v���z;㥬��.��:�C{(c��Lq�ɚ&�Yc�#�л�2�mI�<�yz�:"/��ɚ�;�W\�*T�����7]����ɺ��RJg{���5^w0*PGY*�7��ځe5ܗ�w�t��J]�YR����͗�.�@�;%�ћ=4Lf���̓r�.�L<C�xȦV��p�b��e��Y3��QwP�����k�Lu��%9�o�mU�$�I��;*��#|A��q���o��\�Wk6�\ϓ��L�vs����jW����Dtn\��$4��K;0Kd�.A����R�=h�K}�]_v1IWr��Fe�'��� ��k�/���[X�V�e=k�N������$��w�{�qj���Z�;V�'"y���]��sQ���M1��j���4�D�Ŀ�����""��{��~��ͯ�޷������4?ej�^��.�d�r'M��#R� �$E���gJ��T������q�0��	�l�wWr����kb����B��++9�y��:vǯஈ���>�hM��"n��zi��Փ�
�bȎ�<�w/\�9��8�ͮwQV��*ޚN�G�3.���y|ۙZw7E�$)��켭�[ѸDq�=���;�M!Tw�M��fH-�ӜBc|)8�Z���Z�jk�A	�b�U�%劺�h㒣 �`}��OR�cTs2�f�؊�p���t;��e,�b�#QQO�˽$DJ�PV�[C�-��W[ٜ�Mj��	��\ot��.[���6�<�ڢ��o�,2�d�9����:�-:k�w7�ťGi<���^�o��M�u���s�k3��S�5����	`��+�����^lq�.`GWm���Ƹ�J�b[:��޾z�ƥ�:��MW�eе�E�f*�0��n��>�J�נT�買�]����[���+��-͕�XQ�:1s��j7YNwb,�_{��*jW�1l���r�.��}]�w3�$��.e
t��8X��5c�S�W)�:m�z�s	Hb�t��"�&��erސ)�{岸�.�Ể���C�R����u�ǭ5��n����}r�R���\s�"	���A��SOZ9���ݠ;���|�X��{�esչ3zB*�]��Ct5:��G����.g'����'E\p��ie�U�
_و��u�Y���99�-E�i�-�{�� �������%yƬ���ԩ9q�s��9�//L��@^��=Į�wͷ�h;*e�F��e*lJ�$���ӳtQfXs�77!|�X�xQ������^�)�2b=d[�8��*�9.�b�ްt�g9C;��m(d���DomT��/���e�]f�PB�@4k1'QX��C97#�gqD۵���SS��V�JZ�ǋ�<��.��-f-T1���FrH�u�޹���Y$��x�%�
���'>H�Y���PԻ%�^���ھ�S���1G`�Yۼ|+%�Il,oe-����4�d�L��Keg]2�����cr�ފ��\O�� ���m؉��e���I��s|Jmvwj�������=��x�*�YY��t��4�<�L.��D�mI��_t�˒!t�C�jN���&Ԭ\��\��"��`9x����T�]3�ێ%0;5TTЗ�o2S܁X]9��[��^ò�1wC��فݽ�O�&��ɑM�����dQ<@f�s���� �r{el���vJۖO��2�\����I��R94��e�_)��}�ؗ�-_b7Y��u�p�o)G���Y���/@�t��]���ZZ���|�:�WYYI�V�!�����f�鬮�����I��VwAK�:��eW: `r'b��7�Xm�Ua�j���إԏ�VPD��%F�X�rԭ<�NY����pKH�*5��8ku���8ip����f27+&��=�� $	���FSk��aC���źwB�9։��r2�8�r�������3y6h�6�L��1�i�c�T�Buec��d�;�+{�눎�N�YX:C(D�_-|{�,C��ӷW=����	bֺ%Z�)C1n�P_5ү��b��"
n)��֎+�����ПRˬ/.r��L�k���x��Vo�nO�N3�gj������=�r�*K��l!���V��l�/�M)A�C{vs��X����7&�'-jN����Z��j����A�;E��b�nh�`�_]e�\u�4�:�qnB�>&��oi��ov�Z�H]�\�m�QOnH&oC)V���Ag�=c5u߭�든v�!�j�}n��dڐu����A��@�G[s'[/�pK�]M."���Z+rt���
��km ���c�[}v�(�5l�4���$鷓,3w�]��[=�Mj�)�tM�p�)r��=��D���KS[�nQ��՝/Oih��]��0� ��+���2;6�lZ�.v؅@�c	�!x9�ԣ�>X�e٫���q��ø�8wd��s�꺳{���-��{H3g��&�MK=\�_b��n�Y��	N��F�^��}�����jIw�BI!�ud=V#uG�VeI���=�.���Ů��+>wm�Ze��3d׆q��Dm���fJL���&��{�X�����0�Wz�l��=E�TaTXy�sW�/�Y(ښ���m�49<��c�8!,�M�յ`�&���!�^�!��P�ˉ��.6��[חkn�H^�׽�2����;�ܜ���y�Ę�\U'-��"b�9�kK&�ͼ�#�Cz��F"�:�a�Y:��	0���dpY����Yy�o���5ʦ'u{��2�-�Xx�Z�۾��>J��ʛ���Zi�Ês���t ��۵ݖ$����C\�[q�f�2N��FY�v�����N���U=�6��:�~�5n]�P��\ǭ���22���r�@�����4�l �3���'�5��V.,�#5����@��b�v]�o�_E[�}���5��܋8��Pts�;$�+�u*��,튱Vl�=���vjZ����Z-?�]�٨r�R����{�^�څ�FrSSU��C�|�Ըi�>nPM��-R�G�$��F��b�3�p'6���{n��Q��r��mgD��hX��%ݝY ,<'��EDK1u6�5,s�fL�ݶ��Ut�ջ���� �iΖL10~g.��ѧH���ۗ��ࢌ��}��E�E�]³��]/�u�U����RR�/W+���umv�6H���%�wP+F���a��J�`sX��CQ��n�GS�{j���2�Zd�X�MVN!I2j���Ŷo��;w�о��݇�1�b��e���ɲa�K�p�!DX��{*G7eb݁��s��i���Th��ܜb�]�-�2ã��Ze�ݽ���3�囉=
ĥ�	�ue�e��8i���
l](r�\r��ǖ�ӳ;]	l<�é��M]�����6�v����wx��L�ʱq�.Ш��q�������KV�=���]�3v��J}O{��`�Q�m.�K������$R�U����7s`֓�Z�<����cl=��`�֭�xm��s�3 :��VR|6X����*3Zl���z�2>hC�;r.��@*7 ��2�,��=is�#pP;l��M�X&d�z9�֣�!������'�]�H�X6S,�a�8ZhS���JWKy��v-|�q}׮W]�����)�k��]�k�n�NB�e��7[\Dʇ��k�ե��nT$�MQC�8�5���	T�&��hv�d0�r�*���U����t6�9��M��,S��z�)L������Lʺ��z�&���a렻+��l�1���s����&Rq��Ǭ���C�n��c޻��RK�𫴯���e�F�!F�Q�����6�C���Ζ�JE���1ħ�˽n�%�
��u]#Κ��ai��y*�ݤ�o>&�u��fdm��go^�H�cN��t[\��L雧 �uh����L�jq��0^����z��\�tU���h��X���u���\��v_8��Pgwf�E�r��$.7�O��fޔ�AH(lïWoq��+:|
�YC��zųx�k���A�o�5
Ѥn�`���_:.���;c���-T|*�Y���O'�zݪT{���'O��h����[sp:>7I����/E'ԻEE�T�`r��$rG؎�b���[OVe�������z���Z���.Ux�u���k:f�����n�w+��K��8�D�jvm��Zʷ
e�i�{%�F�U����+��6T���-9��+�$͕�A]���a�㝸陋'������JQ����ֱӫ"�Fu��%�n�G,�Mi�6f���!�@2�]&>IǊ���5�㝱��ҍLR�6hm�U�(WSzu>1G�U^2p� �0�`���K�x��_d�v��.��P���Wb��$̵�Z`��NI��^Ć}:Yu2�#q>��;��n�zv��wi.1nP
��.h�e-��]r�b�3�XyԷ�1���ts㯖��Nj�R�����u(h�9'c�)wi#��e��'�m7����Ιs�������ev�E�Kq�i��M�ܾ�:��[���s(H﫬��B��:�#�f'K^@�d|�C�նj�j���dU�q��i�]�鵲�d��vtY}I��'7�ޚW���Nk�Uo!�ܡ����v0�cG�T7-�J�����V�h��&�1,�Lq)�������)���y�����Z�Q��+(f�"���@�k�g*P�V��b�	Y�uۋV51N�g�:��Mn֕o[��
ߞ�T��!�m�ƃ�0Æ��&4��L6	U�,wj��hŹFK�p4`�����7{�r�z�� �w�\i	3B��KƳo5���%�(vԑ�5^tu�"�&�	}��8�8N�YX�w�&.v've%�� X�m�{��VY���Y>��S�]�x�zv7{�����9���%c:nP2-ΔU�Z^N�-�u�M��B��Ck<ѦF�M�V�<��zM�ٚ��ֺu����ڗe7�_Xv�bԡ�����pkFe�%e'Md�l�*��S��q�:���]lJG�ạ�8ṦI�����[
�jYa�E�ݧ�֪�˰���3�*?�u�u��V�=�Y1+��|�R��xiͼV�	��R�.����0܊���qL����4��k�q�̬��d+���c�A��4vj�Le�k �Ϻ��/��#����]�Vۡ��:&���$N�!�4�v���<�y5,L�Q*�p!���	ϰ\��'ܒ�U�+�@�L��CB�`W}1�恨)a��P�Z��j֡m��d�n�������V|�s9UҬ*����.o����i�S��S°���t�6�v��[�ȒA�9�
�/�#h(��uB�X�ʮ�Nm����z*����x��W��u����ZQm 2���K(�����l�&H+_δM�K��ڐ���#���d����:��`k:�8�`��j�E��J��;�pJ��ܭl�˻�:�|���V�nv�n���4,�S���Ȏ��aզ8$B���Z�=���[+���olv-j`�m�ԸY����ӧ�nENԓ���}�ʉ�`+��Iڶ5�bjG�F�������� 	܈��X�e����w����}�7k;O#�̒!9jTWOe�Ѻ���+]�}d�������KɹK{*�[��"\m�#���c4���ݸ,<l
\��l�kuW\�f3�:PGz��m��M,�vɉu���L����������qws�{O���J��øk��E����niq��Oy��%���/UG�8��l��j�^qjޜ���/7.M�l^؛�;^��|��fA�n]!�q��}1�w�4��'oJm���"��)qI�V�铻�R�5���q�/p:���̧D�2�(`�NV�O����5`>�y=W�c�5��Գi���e2��E�k��f)�n�e�id�X):�WHjp�V����%Ϯ�@gu�G*�4�����f�@3"��aN��P/���R�L�����{X�ڙ YϨiٯ�c6��*m�xj.*R�o0�7�r�a�ꂯ+�>�\A��et�H�͗�K���ѮҬ@�ǂ��]����L%���7}���]�Jf]l��xRo����E���#Q�u���d��T��_�+��|ծ�bm��b5�_.Z�Ц{�"�7�:��gJd�W.]ۻ��I��S�ht�E��+c3[ʻ�ؾn���8*:��|:��*Z��2�	H��zPpK�҃x���1��쇥��8jj�NAZf�W\'Ftp��e*]�1�dk���kV^H�9���;AQ���=��̍�m�ϛd�&2�k[���]�l����4QyN�ل����qV�^1]��&�FP�vm*.t�Y�2��:�Zjf���.�I�lRj�Өӣ[\'�jrl��C])����*�S�4��t��Y������8[9�|�Qզ�* �z��2#)RG����=`aU�A�t�4BV�_1M��i�e�VP��'�P��.�t�}Ҷ�U�;&��^]���ޠ�u&m��B������;�_[��;o{q�:/A��ѓI����ܜ�0��Ң%u���{O�Y�ǉIqt�H>�P����i����PͬR��xw��Cc~"gtw�_G��!�q�jz(��Y��r�k%쥓Z()@��������'�R�,�{����w�t����彀u3q� T���.2���Q�=���=�N}KnN�mS�q�S�+h����Θܡ�c��Lʵp8{�^n�]E��e;eoe�ޖQ�h_������P��I���f�+�^�;`�9\�d�:�p2�]@�C7dJ�ɤ�	� z<F4��Q��]�%��� ���F,vn�e@�VN(���$B��*�6��.��³v�Gq\��˰N�z�G9g9�R�9� �R���ur�b��]�'��Xt��,�,��|�7#=N��MfK�mri�a �4Ы������
Yk郔9�ӊ^���$������ �]����;U�f''!�G��Fp9΄ʙwR�S���6��+��+A.�[*����h@��+��M��4��bw=����VU�q@ξ���9��y�QK���vބ��.�Č����8Z�u�*�QT�s���ӧ5����� �QR�\/lq������Z��˙L`b������\�:�F�5�v]���nIm껫�֌cd�q`uv$+.$�z�yQJC��FeC*��7���o7����өv�c�i=��=&
�.=P��I�p�6m=�:�꼏����<"l�v2�]晔���c����i[l��q��q�'��o�S�@�	G�L�:AW�&�;�:U�ZS���c�֚�l4�іGNm̈́Z�w0�+oﻩ�h��ݞ����/0����V5*
3�*s{���:�>5hN���+��E�1��f]�Qp�ƶWVD&��ї���D5#��7���]�D�l�fmv���Rџ���u2+��QLS/�.�xhw+�b����]*b⧜M��j�F��
Q�|�!F4�Hy�(g٪��哓��W��Sm_U�{s��֚C!��Hm������A�nf"#�R��\"sf�:�j��(����F�����O8 D��z�M�SS���e��Px��`6t�([/;*"��S�P,0�hX���6�T>���t�ʥM��(c������*��F���r�Jb+�vC��	X�r�4n��D=76�:��[!xھ��TN�c��5�d}�(�čl���%K�y ������(.��P��$\�{�s���НyHq!��m��O�,t<z�@{�)�*�S�hG�B��/U���IR��`tb���f�%��b�d���$�3r���/��yM�H>B�K+����/ogm���� �"�p�o!�^v1&���t=�giкr7��
�*ZJz�P���i)���-)��Z�P��Qi����(ii��

(6�D�F���Nڂ*))��������(����;d�$h(����Jm�D�AEhҔ�SPDP6�S��j�"! �:"j5�(
)i�"��
��R��������)��JV&��gEE-U#���:*&�@���SK@R�� D�Dұ:�Q:d4�٧KC�1!T�A5U�S1�KM%#�EREM. 4�%�ADAKTҍPRR�BS�HD1!HP%�HR��P%#AQR���H��^�]��w����θ.s|@\����=UαY�*\V&;ד��rc]ĩz'N��⮸��K�I];k"x*��[s;~�*�'W.�Um�f���k��qHeR5�Z���U�nVS�� 8dc���V�|6(��
�,�Fi`>�d�D��PrpvR�l�#����]-���V�Z�eoA�#���}���(p��w���˶�5�Z>(K���>W�N��S̵�s�(���m�ʕz���j�\ӯk��5{%����/�p5��چ:��|�N��o�wxag�\�N-�^��ÙU�]k=�Մ���z��aVF�w���.9�����L��wN�p��c�Iڅ����k�^ξ_SO d:�L�;��M�����Mh��K09݆��"��]�\hY<�����'�E)u�ڠ�_�1'��\����b;�R���ʔK͝[�sU���̯JK*_m��@�t�{�<�����H,�s��h[j��=��Ls�p�|�9�J��s�(���b��I�t�{Us�]��Y��.�l!=��68uf��y�nk�ؗ���#��_1����B��e�������aԾ�
`֖�@#2e"c~�1)5ad�Np���wҙ� G�֟�Mtt����Z�q����ƒ��+&h���1��*h������rζ���o�*.�7���i9��/lm�;�SW-��k{�6�`t��]��s;#�6</���a�u�w]�yO�4X\��Gb9���,}��!XyRͨ r�ʥI�K�ȺȷI� ���"o�hc!�W���N�����tتs��-� �w.tT������d@ި���u�1����]�PB	>���"b�Xd܋Y���=5�015�޳i��f���ܥiR��4�]D����g�׫���P�*�'xY�p�VP��Zԃ|�5ktq� p�c �n�p���W���OW��o0..Ll�!��i;3�8n5
�Y�=�}�W֥2d��p��Q1�+6�S��c��?rǗ��i\�aX��~V�1l�ts*�Lܯo������L�S2���),�+J!j�x�c��xw���{o���kx��e�iS���Tq8:�^�R�]b��0����p�mΙ�{uQ��;��)�	��7�tӳ\��H�z�@�`�_9���A�	1Ƭ�� ޯv����;e�9���at|�UE����v�*�	�����̖<����D1\�m���I�� �f�*��0�"yQ1�*P�y%>�R��l<Ycc��h<����;St�л�^�Xcƾ�ה��� ���H%y�.�<ؙ[���&ټ��lh��9���Ƕn�Γi�WS�2�;C��6� w)�Da��%f>���K��9<�r��\s��u�Z�:�d��w�Q��e/$��20���g���{[�B�� ,u��w_0��1�7u����U�"xGA-4�ަE�޸j]���8��Ԡ!�w1�c�x�~:��.�¾��ύy�w�]����1�A���niŜMB��B�Ezt:��S�jhE}]1������gSU^����#5��(���p��욃8�7���'��x�4d�k�&����0_9h����c��w;����Cݽ�'M|�f���6�*S�u���S̪?h߯��J�Qà���D)a�����K/q�`�Gqq�`���M&��� ���#�n��>�
�U��eGmAͪ h���M��Y���tBd<�7Q�f�K(I(TuI]6H~h����L��Ͻ&Zl� M�iM�?5����a>]l&c�0��d��� �n��:�"�۲;X���3���$��pJt�i<+�iU�x��c#�\�hӈI;"�Nb5�U�tl�]r���#sռ�[PT~��Cmݾ޼�+�l�ܸ�rZqY���Oq� %;`5H6�rf�k�ML9�hKp�<.l���Z����wlx�7�I��9v��v�2��ٳ����W Vh����r��u�[���*c��Y�/�vi�n�-�x��Η|��'�:v���ҽ���[���뿐��wt!2�7,P���|Jnh4%���N�hya1�U#�^������^ǘ�`p�iVo��>�1���ⲅ�u����J��p9Z��Х�N�E*g���8=QmWb���1L,��.�=|=��w~�x�+��ċsT���(C�:�'r=���eA�]jǰ��:Q,-�H��� 7�c�3T�R�D8��y���g}��Λ�����
([�k��mN��	Ƣ�Bz���9cJ�b�ι����ύq���lc���)��=��j`��d�w��L[Q���<B;�&��� �R�p��{"�p|_	t� ��mI�l��cv��� Cn�vPة��C�L�:1���\L1����͙�!�)�ٞ,�R��[};~VsE���n!>�n7��i#t���5����X�����w<��)PV�^�c�H���N��nJ� ع����C�V��.�\��pQ��*А��]ȹa�me�cXâ�7w��u��[���u������;��z�Sv��F�r����X����^�=Bf-��c\A:[Bҧuڀ=OR�
�R2�:���}���-�7�<����fFMQ�����(E�ťd�\]v%*w3S3�����9	��ݑ���ߛ�E|��*�@�J`	 k��oRٖ�p��塑0Dn�8����i�`�M���ݳ"�6��Ef���7[^c
ۇRs�lޚ�8e�1�p����A���Ɍd�u�Kt�'�ޔ�ag*b�k��w��x��D��axP9�{M'X�u�dE@�s�JY-|̰9��Fh��cݻ�8�zW��DS�U��vP6=�������x;U�U®�=	��,�s�#�I�7"�g�UÇ�����cn��a��*U���>V:ꟛf�3�)����-{o������b������r�����uC.Qɛ�0�@�6�X��k��+o9�1w��������6oQ�w�#�W�>�j����sW3�ꘕ�6��lޖL`�;w&��ޫn���^-n�p��q�Ow�F��}�H
�ֲϡ�TEru���VȎw�k)��c�޲�x���fu��H2x] �C�G���B����/���A���f�N��:!���`��5�IY��#�J�wK�5Y�7%)��u��~�@
�y5J��2<ݞ���.���M�r�����Z��Ղ�ՖN\���������ٙCy�Y*dW'=5#,K���k}�J�)^�z��Z��%]qΜȳ���O����y�.�[��kiq��t�@��*a�U)`zS���� ]9�{ֵ=�n5����꘣%��:�HBr��e�=�.W2��Q�i0$8z|�K3��擻T�3��LB�w:�]�P)U�.O�;�n�3�LiW\:NɊG�'��.�qS#�1�;�p:�!Ѩ>�!qc�К����s����2�>�B�.m�����Ȁ���FW�z�����M�}�����WM*�u'/�Z�#��i댘�����Yݣ0�0��gsw[�1� � I�O��B&/�h�WW�[<1�]Ľu�gc�8�Q>�q=�۬���tx�=�,yW�ؘ[Q�u�T|�V�<��-�̉4�,%�]�����:8q/��=J_��4Eh�&��"�~e�[��.�#*��g'��6��{�w���%�-T�lL1���'���6���W���g/�;�+�F�-9��N�U{Z��ʾ��lBR�2m�@s��D����ͮǅ�T�Yh�F��&�ֆ�'T��K�ʶ��n��X��k޺S�n�/6*!w�ٗ��'����C�d��'i6�ܶm�Z�#�/�j�0��+���w-���9֬]y7�l�$߯�	�k��P�
��nCW�ZB8mR���R�ŝ�r�ř��wk�l�w���aU�㧟$��_ю~d�r��&̍�0�R���n�%��q=���g���5�`_"�ҧ/G��X����T���70��n�X�{,��3/bf�-�af��F^F��/���ÕC*�n���ʿnT1W����g���>s7ԙ�S���my{�t��*�f/�vпW-'vʮ�<~���V3��P �z]v��"�c#cg;YNL���t��r����8/<�u�Ƀ-.���Rߛ�i�Lor�ȕX�)w2u�I�� h��e���e����<(1�JQgB�_.�rļ.�N�����N@��v��H(^NS+>w_e|`z\�q`��XG-��7+�֯b�h�	������9jhB�,}�C�3 ���CЦ�ٷ<����cuP�$�w ����xq��SW�3Ý%x$),Xq�Z1c�λg1�Y�K�q����o���g�W��qXUC�ب��D��=�Z�B���W�>��w�3��U��ց����[��Y�z��5zR볿޹���Y�]Q���xΫ��Z��s49���Ś�˸�۹��d�oS,�$��[�NI�'J�gYa����i���٭���0��i]P^t(;�V�R2�vpJ�9t��*^vh=:vc;V;�c���7��)�%9�s�� }$�T��>���i�Q���Sw�[��uN�o���M�NH��`����:�4x"x:���(���V���_v3$��+�2U���5t�U	u�i�p�4�]� ��0��I[��f9u[11�Q��-3Ya�L!"��b~���rB�<*LW�'d\'1���nMふ�$�m^0儚9�����~�т�b�e١�V:����wB#��{��
^r�;(,S8d�����W�5`���uP�^�8>���t�
�:�����Xcy�����2�4)��sݛ݊�W����}��:�v")S>&*��-���j�_Y���$�V��un��
�E��s�w3��%�jX�1̱9��f������S�L�O��ʭ<���&��5׃��=�_z(���G��b&;\,�S\�%�g����]f��1xcGY6o"&b�t.���5����Z��q3��zXg�u\�U���`�L�<c1��
>�8'N�\�<b�.á� oc͊%�e�R�0f�a�{�l�HU�P�>���q��}��̏� w�	���(�8R�uu�ޝ�r���k���\�3v%���i��y.��8�μ�7C��ى�h͹'*�}�$����\cB�,Wnmv�VgK��j����Q�.��0t�������
���Zr����p}u�!n�QX/�Hu=U�k������3�ڃ)]�9�>Զ� �kw�#\L1�N�>��;�\Z�N�n���ہ�鞜BF�s�@zc�(�q��c�Ȳ��pK8¬���V�M��}�	�w�_Д�cn1�M�>�ۄ��v6rJD�z"O"C�{�X�B�A|�)۞S�{:��K��늳,�Sv����m�Z6ݰE.�!�v�����n֋A�CQ�P`�Xr��BȉN�1���u*�yQ�y��%|N�)c��;54z�&����@K&���c.���~����2�@�D����mR&�Q6��^�-e/qZ��$Gu�"t95V���%_v��;\�I*d�8����VH<�{���<���"+@����w*�C��Z��tz.��N�p��-u{��;�D��ok��V��fb�9`iy�dY��t�0�
����K�0���>ĭ��қ�m���e2rK���j뢮���s���kr�:7[�N3�M��Ue=�we
t߲�/��N��g�mK�Z�H�5�������{\�![�[ܬ�O�B���w�:����t? �jݼ:d:�i�{ԥ��6ӽ�:�a��p
N.��]�%պ�\�d �]8!_'w�:���Voy����%w�
�U�g����O��1��V��r�uc<�|K9Z�3�S��xb�q\ι�'��h�nbܢ���k��\���lȪhгE���CVH��.P���k��ݕ��V��~1��,���Y[n[�qU�S5C�sFǾ�F���<'j<2���s�C����+�W�,l:{�P�G�T�!��ͬ���=�^�H�8J��8*:?�������^���P6�cQ�y*Bh�e.SO唄uĺ�k�Y^\�e�}Q�h:C����v�jy�G�ج3�f����|����:��1n�1�+/���]F.(�I��^�\��3:q��5�Y���n������hM-v��5%��4���&����q��Д�A۠~��=�Y�5�$t�L��O@��3ʥ?J(1a�=v���#Oa���uC]��pn���ά�aWN�����'�a &�>���W9�!*]\#��܄���[Eb9�YP�t�4V�!��\��Y�sk_w������ml=�Vg_3q�:a"�_V�C�h�ZVwJC���x5��}Q�W����M�w��V��ԤQaB��{:��{G��O�[�����7dۗ];m�%Z������Yc@f��2Lٔ�Y�#���3.�Y;�fR=��h{ީ7�/f����OLv��V=�!o�9S��a�W��
�0�f�9>eƤ�#d�������PG9q�ݦ�R�l�1�*`��aVU�C�������̾S)���(41�-��8#�+�;s���i&�_J�Xu���9N61�������o҂*��]� ���/���c����a����R_�,�}�`b}���;���}���+���.wWH\w�
�w_I:�&�1Ժ�N'S2�gm���P�#��\���ce>g�u�9[�0�6]�,�B����5�E�U��
mlgVՌɸh����V��Wnk��j�]j�2t��xa{�) ���Y���'h�$u"�'�Kj�uE�G��Z��wT9+`��sq�b��޾G�7�is�Q�,����t�-v�+�ۢ��jRw�)Nܓ6�����׏i�3��.�z.ẍ�S����YX_u��s���E�>��ٴ��`�P3�Z�I�n���ҧh�X��Y���Y�m����c�l�Ý�\�N�[�|�pϙ�Ӏ%@�=v��/2ZӘ�
����z?�sD�j����|mY�4k���Z��+��oj��Y��T��ҙE..�g'�4�0�^��²���jlh�߅���j`c�>��k��_
�w�i"'T]��˾�]J��e�3�pR�+R\��D;u˱�0�캾/k98j.�Q�,�t8͔l�uդ�Y��뻏F�,�̧�.� v�3]`��ɏKRZSk*��q���k&��HR�=�u�+�KM�q�Óg>P��np��-n�����
�u�)�[;3�1��՝R�x�JH����6��aM�ت�U�5����\�G�<9�8=���:}���=�ep�v��'F[s:-`���N�b�Ȣz�U\l$w����er�3hnd�=]��_sJ����v�A]Y�U��|i�Y�e��Z-α8�V�q.죜�t��r�ܛ���.M�]4�^w %��y�J�������Z塞����0�:GR�G�]yLV�v�9���-�w3t��ٔ�{��^y��l�S�{���,7�e�Ec#f멦����GH�{�L뎛�2�-C�є�d��S$�X��`j�!��u�bHͣ:\����*�/���� �mK֋$<��S���z�P��ض��u�s/sv�7-������U�(F�LO�0����Ҹ(��N;u���a��9��t��M���v�m.�쵽����Æ� �m@y.���;����r�-����7�o{��#V"�9§a�ә[3z����W�(
)i
h��J�B"��(h���)����"V��� (�	E���4�-QTCT�IB�R�14K�H�i4����HJ%#MP�-)IM+H�ACK@U����(U1$U)C�ZE4&�MM%RH�AT%EIM1D�4�,ED%N�@�QQ@�E+2�DHL�@RR-4R����
SBPP�3N�E4UE%R�Bm�ih
R )��
�
iB�*�$i*�� >�>�9�3�szv^uY�f)s���u`�w�;[y}�EɁ�Έˌ�U4N�B�Y	���XB���+5i���n�N�ӥҼ�W�}@|�}�d�{��*�����(4{!�y��-:}���@h��N��Ǟe����>��ʏ�w�~�r�����)�������_g�t���v+8}��Ǽ�ڬO/=�0`��#�������/#�y�Bu?��>����}���y�\K���4��ʀև��r��K�0�z����;��r���w'#�?���}�U��Y�ף�\����""�}�{�:�9/%���=��ܻ��v��i�]ͮ�� ���={����&�A��=G�}����Y亥�r~s��HRtsy��a�0~�B�F����wWT�}}�#�"���?d9=��<����I��%R|�����!�<�y��9�����x���4�;��p��4��_2==���u/�uC��@y�R;u>�lD�y~_�����#�|��/sʐ������o��9�����I��?��%>I��=��'������z�h��9'��^��N�_��>@u_����>O?e�XG#�����K��Q��|�r9��z"��#���B]��J9S�]�w/��]>a�:�K�r�����u�k�_��|��p�|�}���}��Д�߼^�]u>���<�<��^������z�5K����}��`���>�=������u�r����������Or~ۗ�?A�K�}����c�y������������4�.�~��ϒ>����/�>�4�>r����̤�ss{�T��b>����yLu?%�/?�ϧ�:O�>T�?}��?G�:�~���O��A���p�� �<�s��!*��X�P��C��;���]�sPF�I�����l��x�j�{M=�$���
�{���C��hu�θ�{����u��ޟ�~@w����z���v~����������9���A�o�Y��\���S�!)�z�c�:���}y_r�,[��Ƨ1���@F�����:�-:����ѥ��:~O~��_����J��w����B_��������t��o#��/W'�w�������/!�}������>���%F-���≛i!����|V0U���T4%w]�珮��8���/�2�^戯]G�:��F�����:잜sӰ*C���i)$�5�۠۔g!��ۜ�i�o��Y�*d}M�o�O���������B��f�y�Ҧ���S��q�����"EB�vu~���_���&��z��]e��:����w/[.��?~��!���~��>K����t{'#�G/�{�:�#�9G^��>BP~�Þq��;���4�A�#��@����ι�2���>�����u�������9��N��g��:y�K��#󮸇p�]���|�^��q|�?�?q4yp����J%�	�!��1�7�l���.��$�}��oz�����'��%���9�h>w�����^����4�N�����#G��:���'ǭ�A�;�쿏�y����F���t�Ο����� ����>�U������������ЩJ��c~3K���xv��1�y��C���߼��}������$�|�C��(
(;�'�n�/�������4}�O�e�{~��h���w�_h�����~���[x��~5+g/�B��[���>������}�>�<�@h����|���A����\O���i�~'��>|���u�i��^F��B���y�<����Ä�H����$B���Ǻ3�ޫ����ĝ��+ާY~b>�>�}#��G�F����׽��<���}�_�45�y/7��u?e������~�r4�G�2u�	��?c��^\�	��y��
w�~�G�}� }���:j���@O�����9'�4��nC�<�A����r}������9���>�w��}����{Ρ��h��9��r9y��'�Ѥ���>^��(�5V+�>�#�F:�`i��1�����<����]���?e��%�t�.�l�F�/�������>܇���9���?Cλ�I�z�BW�<����9>� ��yE����P����VMO�t�v�Td.t�!���4z��=O}e�y>��BS�͞w����y��/ʟ�������=����y���5�^�w�G�J`�~y��:�i��{��e��:�H�l��ҫ�g��8�p��O�c��@JC����_0u=K���xz�c�r;��m�:����O�����BQ�����O�rO�̜�����?������]��|��/ <�;{��������q�S�X���f��AH���K�>Ԁ ʐ�ph��"�y6]n�6��,v��Js�;e�V�P���3�ٹ&us�T��+��yـk\/+��>dPLc>4��g
�ym�1��eFB�6Q=g�,΀bѽb�W�}��XW�r�Nioﾫ$}?|��i|���9�?%��=_�W�=�O�uO�`�1ԝI�O��9�����۟p�}���}y��?��%>_C�O��O��~g�'�4?��Z�<�e�^�+P�+�N�7�����B=������w/�cI�u�I���/ >�� ���!������=�u����?����C��x~����?��9�ne�<��C��=܃G�9�	������^�[�T�)w��Y��c��ѡ�9!������䜟��}���KEO���w�Kܿ�>u��{���7����������x?c�%Q�}�����pr��>�ʟ�w�� �D���#�ؠ��t$73�A��}���}����(��T�����G>�5�K͗��:��pz�e�/����]Ƅ��{Ρ���e�Ǉ�x��=����9�q�J��>����q����{��}!�C��>�"94���<�y���O�>ls��K�c_~c�z���?��F�˝���p:�������|��K��s���9'�j�}���#�����W�W&���_��+��f>�>b#zjD��9	G��9���~I�rO�ܜ�4�ps��:�������I�{w/$�|�A���_�?�|��!�o�����>��t�����:v��>�~��ԁVs�@�}�������q���~}�ϵ!C��\��y����|�nq?ZNO��~g�ܜ�I�����%R�G�c�9	y�������y��\:���ߙy��xv q�� {}�733���o�#H��Tzy�}/�p�A�|�9�e�O�>���4h�_�/{ù~@y�{��jB�߭����/Q�2_7S��/w��|���]�tl��4%P�*��˙�ƎTc�/�Wz�f9>K�޾t&���NG�����a)�yם'#�G >���}�^I����s`����>��K������_3伀��é��si
�y�����K1��Vi�l���y��!�|D`�ݏ��%:�r�����5T�����~�??��}��u�?`�c�����OS�����*O�i;��=��%�?��q�>^���i(���z9��Dq�h��I*��6:��q7��)��^�4���V���ٜ�V�e��,��j��
*�-?�f�
|O��b�vs��N��Tj)�ȝ��;E?�Gf�\��.�jm�sodT���Ż��mh�,�����:�j$�^�c6�U���fd6։p�yw��#�켟����A���z7 ����9��X��~[	z�C>r՜X5�d���ɾ�)$��d���S��zTEĈ�4���]3�ia���oY\�~�/��euX�/3�;��8N8fxYD`�t��
���d>7Tv*__j�]#^�U®�p��똽zwF�N�rs�iU���sr������4йu���ʣ���Q6o=�R�@|5ƻ��T��vUF9�ݕ��wzs�΀to
 F���}&�hC�������y��ɵ�[[�?q/�.��S�N���Yח��zb�8�g>�Tĭj�*�޺�t�վ�NE~�)�e��'��ᐚ���`��D��~u~�'r5�cj�36>q��2��XJ+�|vs2��+��P,7�����7\.�z��B�u����g=?�{�(nܥܜR���tU�d�����LJ)믻��r�����9��'����:�3�uO��1xK��{1�ZrQ+�6�ǖu�[U��l<�#��u�F�5��c[t:٪4&�#g�v�v6<=�vװS�]�Z��#NC�]�Hcڂ�u`�}�\��Gj����L�f�!��yy��c��DeL�\7דY���Ͳz���
M9Z�4�&WcFc���櫔���A%��V�lԺ�5�j�I�pem��pRW��E��8:w���V��_�興'4���n`��>�2��G9d�!��	�&b�t��ϥe�%��`$��]�9���@y�}�=��B�Bo��EL�F�GBF��-v��5%��G�g|��b�*m��gD��ɤJ`*
��n�m.�fH!�6�:|򘸊��f�Z���J`�z�#��i댞a\�j� .sl:�c���S�z*VZZ}�J NtT\ GT�N�
d�b�_E���03�%�|�|�!�o$ٻ�*L�ޫ��p*��P��eC����;TM1��u�b�8[V�8����L���"������l�0a.��z����J����H��q��L���{�wo#]w|��^nw�=��wʡ�Pۮ�8#�uL��,��M��6tմ�sM��o������:����>g����s�!w.�(����W� 4R�1�RҦlf�3�)�իRp��r�{။���C��\M}ח!'wF.1�̚n\��y��k4t����W;�0�}^4�u��]A�ס�.��O��Zpϧ/M����$����[V<���,�y[g�,#�@:��CU�oC����ghT�͠�����9j�7xT�B`�f\�/�׮'<��������0�t��p^�sݗ��u�p���X }})Ṡ����[��M�C�4�3Tλ�y��ui|��pe�6~��7jj�}�+=�DD@��nS��ѕ���ǁ�[����f�j�d5�k�X��k��ي��
�pш�`��.�P>�O^���E��6�U�n升I���~4l��R˫rrñ���3u�s4� f�!�30�-��{Z)������\a0GUwЪ�x�{"��,��=n)��R���h�p Os�e�U������Ul�Ux�5�KmМ�j������bؙa\TΩ�� p��u��H�(^�g�5hB��:t[��r��>|��E+>��⠎�B�:J8-ԾS���(�,|�9�n��W[7ή)ld�uGtj�Xm�+{�G�����h����Ү%��r>+4�p^-�~��k��ܩ�kվ��ǆ����p�e�G)3`�@T)i}��n�a���.���r�˔���\!qe>;�'@of �sA	���� �t>`��L/�w�B�v��l�hg���&5����.�9gD$CɰvvFۺ�_$�*:���x3&�(6���b�������q��Q�NQf�D�V1W]���b\�Bl�:8貨���^�Bզ���͊���ۏ�u�8.�*A�q2>1r��;n.��R�x�C�k:�Aq����]]�V�L�
��9:��_Zn�yw�krUƝ�7��p_�����5z�zf�6zi�=<.��a�aR]m.c�\�%g��_7V̌k�,���M�z�K���Y�L��aՊ�S	��>��b�}��:�Q�04�%�qlt�k��F��rm�_U�ɭ��(�q|� *�w�u����Ҿ�P:��B����_1��܈<�R����%J�ۮG�d���v O}�}����h|L����~>1��
�?�6�<)Ͷ���	�׻��}����8���y9��ZY=@�|F�����3�N�b���֎w�BÏ�%��]H(%���b��T��ʱ��T����@z7��pj��i�Q�W9��8'���tR'M������Ms d	gY�n��?'�LG~�Ԍ�Nߟ.�X7�8$l�l_���M��)�����d��N��]R�V�N��є�*qX�2̞x]l�p�tK7"�wTA�.��(K2 �س!ꁪ�
�S̱�3�ݹ�bxv���S}��S��գg�,��٨g}�<��6S�v�ϐݩ�r$��[ܖ�M]�J�^�1a"/l�LH=+ޫ�䍻�^r��{>̷�=9�F�d�^��q�C	��6�6e�u�k��Z���	�ϳ'j<Y�����m�u�D�t��n�o8*��ƲI��4���f�aR�+.Ps�!=��YY�6�gO��"">k'��L�RZ5A�/�c�;o�U�½
�][��%��l���e>�3�K��@�Vv�=������Ӑ�K1����R�//�cg$�R �5x�tT	ʻ-���bh|Ŏgn.h&mZ늸2�a��L0��k�#j-�#.բ��gA��Q��4�f�)�NӤ� &�� t'0 G3�:-3δ<���9�s*ۨ9Z��y�{��2]��{��lz�J�r�#�6`[4.)L1���~K䝠�|�,��=��U�}��+/PGc�������(#�DwXP�H��/�y��[|<�9�p�}�AT7Ο��|�
�����[�]S�gJ%?��`sȢ# ����漌�P�7Fc�K��m��Ŕ�i|[Ț���d^,N��Q�-Yhg%W&�
�`a}�3Cn�0&:a��<��:)�9��L�Du���\��0�)�F�vcEGvT4�V�@T_х #y!�v�Q�
����]�Бi��3:�)���n��_K�q+I�q�l�/�?�V�װөޥ�2��x_LU��0ގ���Ď�5׭ë[ھO��@��:�;�ǂb��y^���\K��)�K�7�j����YN�ۢ�
�/�Y#m&@ޫ�\L�S�õ��~��k/�y>9+�sC����/���;'m���f5�ȩ��v�T>�Ȯ����"#�u1J_4v,?��cp�%�Ε����c�\��W��폷�N���
�L�,]fS]��vή�Q�=�{Ƙ�.�uƀ����<-�ӿ.���.��@C��݊�Y|δ�[���g�!����s��mRQ`���;��^9�HC�n����d�GQG��NOc�xH@URy�y=�c�U�@���L�o��~˄�H�;F��
�OV�ۧ7�6�)��"&��>5�L,��:d��D0��;�����[p]t��fL�(V�v�k����8y���P�BQxr0��:����,�.4���ɫ�4ˬ����%6!z�-�]ޞȧ�n�� ������ILI1��_MB��|��G�]GC������\u�'����k�L��׏Pt��
�� *:��yT
W<���˦}����
�Lf.o!7���ß�Wq7]��J~����" 5u�a4ǳ>\�e9���`�Z�܂48}��'�����ɺ�.[Ȣ`�8@O�'�먶r���u�u֭�n��$Ɨǡg�8�4��;�
�a�ʞfF!�����r*s%f[�P1��w�*��ݻ�)Tԗ����Հ1������s�a�a'{���]@t:��������>�y���h��R�[��9<���޹ۚ����W�W�l΁��p̫=~�O�/��-J��P���@u��.�wl�M��������ܙN	�u�����\|�Bѽ+MGs�}˨���2d�n��ր��9����xV3��)� �/|mh�<,*\���{�������I�Q�G�Kn\��} f��l&��<�y��<tp�5� �r�_xpJ8�^3�hXB�>�bqYp�n�k��8��������5yr�}Y;P2~�s+��Ƃv�<s�0�L��N��Z�uVftpi�p����x�b�f��������c2��VI{_W�s��5
���U(��)�v-
���@	��������p��ӑ	�p���C���\a0By�j��L5=S'�g����%|�W�z�t .#y�2�û�������wW�Ul�:�4��gUCe��k��8a�,]@��n�]]>@@�*𕜨o���7\�2�)��lD�=|�\��$�E�c^�gݫE.*��
��J8>�z�Ѕc]1����q�ٻ9'�;)�/aU�+��&ȗ����dX_Ew˻����nuNu:� m��*�)P���;-*Kޖ#��@�^],8�tWU��kH�e��Lt���j)P=	1���k��=�NM0��uEWF�6�ם4Sw�Q��R�ݝ��&�ޜwm��yЩbX�f��<�.Jg����Q���ve������;�v�1�gc&k]+��e���s�x;td���TZk�4�L��ʛD�������ɱ%ѴkR�b��j6�z����
}ll�:ɗ:3���b)mul�o���L�s(^q����}���7��$����-M�-��)]p�Ѩ�\:�|nJX����lr�fG�]�A��-�1�3���	`}���4����F�p8�o&��V�xV��W)� �j�B�Q��N�Day]1��P�T�amW���o�3�u���7t��J]E��M��q^�i�nM�Xۧi���x7c�M�\�.�G¸���T�����N1V�Djjp�}�l�l8���Vj�n`�[�Y�w�(ɵݵ�R�U�
v�gb����.&�G�Hf����P7�v��$����Mǚ2�.��S��N�wD�ƩJ}X툧>y#@]g,#�e�]JZܽ�#)���Z��a��X�pIǪev!iԇ0T���()�p\]\�Ԕ�������Hڼ����!�a�9)���^�ٯݝܾz]�ұ�\v	��e�z�Is�wҠ64�f�z>������JK u7z�F��yj�͝y��٧^��:f��,R� 2�����r�%����}QF]f�0-�G;s*�R�P*�u6���WQ�����%fve�2���r}�<�d4�q�۠�f4n�N}�U;.�q�2��a�z�b���@z�Qq:�x9���2�T��Xjˢ��X�E[������"��5e���=������:�.T�i�{#�A��E�����;+O>n�iF4T������˰�T�ĕ!�j���*%F�$�s����_J�ݧpR�ػ��W6��f1*ν5�XL���]8]%Į�R��$�#(Y���E�)Ak#=Rz��tlk�Y�l�C�؄T���vz�gAYf��n��Qn���(Q��<�C�[��8��rH�Yn�5͗�N	W�پ��;����]��m:v�=yզ���H��&Q5�%�Lsk�� 
1�g�J�h�؜ѶqV3+�axؔ�\�r��\��a�oS�2�%:Wb���e�����=�Or�'D��(:��^��U���=Ɏ��nMrL��wC,g"��t�{�s-��kV1мBL�ud���m�L�b�G�!s"�N�̶�1�YvX{Ya6M������K�o
���m�Ρ�ާX��c�["-���YW/:��X���ۛ���Ju0���ge<±L�jv6��֊m�0oYf1sL鳻nr)�'R��k�wWg\�A�Jî�=}Jì5�S�2���)͙��144�$LBU	C@P�QEIGS�)�
JJ(bj%)

��(t:
��

J"�((j&�(����)(JV��(*���JH���
�) І�)�H���@h�


B������F���ER%P�4QF�th(���֊���h�*����(Zj��i&J
��mUs	��"F����!@��!T5J�4SA@rG����@ĔM-,IH�R4�t�E�b*����`��4��}�v�򦷷7�]�v��.,��Q�(�u�� �G����ʚ������w�U.�3˾���Rob�t��L��v��W�U�}N]-��z���7�=6�Sy��O,�K���;D��d�0O:��b���)�����_�L���R0�1�gn��>�vԣr�1�$�@R)w̬8�fJ�s;�o]��+�=yK*��TG�z뼀p�o������ͯ+� ��KT�of�L�ȫ��G������p&�]���t��3�9�`)�#9�X�������ũ��sJE�r�Ù.	�������/�a�aT%����8C�d��� �!�Y�	�7L~��=�Q
�";�mX(�!�.>��!#�d�\��κ#�qm˹0n6�E�\�{��YK���k��	}����k��\���ኲz��X�5��g�{�w.��
�B�', �?X��*t�z�0��N���\���=�g������۝S׼�Xh�.9:�]j��dF�к�=��|o�P����EfԎ��=j՗a��W����o��߹:���1;�~�f�z��S�pîU�R���^hM�-���N{MU��y�uqPu�#7ռ,؁�h�3��C�G��J���9�+����j����A�T;,��9>�?]�*�f�`cz���j彫��5��\�SrU��N=�۴���146�Ց�'���}�y����S@�toGf�>l<����R=ĳ�.�o��NV��B��{���5�����#k`*c�E���������e��D_��]�`t�ǥ�w�.j�����b�=���ɚm�u���n޳�D���w�u�𿟓�re�11�z�ӎg�����:e�����;�_������i�]��p��h
��Т��m/B��T�Nx�͉��7V�x{6��N�dk��2�����Mʺ��Q�G�=F~�[t"p��S��o������d��E�Q�j�����cq�c�C�%���M�Z��e0h+�y99;�D�J�GRf�
L�����W:��(��0���ڇ��e���N���n��l*�j]��n��Œ����Ps<"�B�?_:��%�l�+ea�NcDo'�3w�w3��^�X�.r���]���� T�@��3ژ�|�����~U�N�C{N�sTt��'!ٚ�mR,��	K��>:z��l";����GG�3�i<\=uT���^/i~V�+ꎳ>�r)�\��o�@e�JNY}���PmPJ��q������0�����˻��ݓ��-v2*�o�J���N�9�٘���6��vt�0��W�ghl@���S��ۡ�:hغ�Ժ4��	dҗ��y�Oh*��>�">��.�0�K��wnF��9��7\K`�5�`(n��Irx�#mT�Ѡ*�p�R"x=�R'�鍗u#u]1��\�Sr��� )cn���
��&0~�=UR�"��({0��<�僥��i��3���;0]M�3P�
�����Fүf�����{��N:c�b�O���TOV�`YVo
����n��sF#��y�MJg:�w�Ne��Ϋ�A-���L`8oOQ��?�����c�\y�Ù�<3x�=���f�q<�[���G�z&$�޹�V6�`�@7�W+��Vg}JX# Kϱa��;��:z����d�W��Y�N��7�+�Ƶ�H�5)��<0c����,���ʘ	��;��k.@X�W "�c Lo*���1r농kk�ƶ�v\�'�IH�ی�f�u˾ll���!"�lel��:d��D0�ӸL�jXΉ[|/�j4$����k�,Og�����L�����dp���#s��e�Y����Qˮ'�MN<�q�4:ٛ���5�[�S�Pى�t�s�[T��A:>DT�/-���c�$ƕg;-�[��ú>e_M��B��r����U��q���U	�ݥ���$�X��-�ǪAX`�kRtb��;�f:�\����yH��Los �n���q�s7��}�}�}��s���ͽ=pJ?����t	<Ҙ����n)*�Ҕ��.3�O�̙��m�c�����C��P�;�,ڂ x�� ��Ϧ�!�pHۋ�̔����T+���p�xcN�����x�
�?Ss��D�� 4#��7D֏\���{�E<$�Y[5ۜ�e]�����5hdA{\�d ���y`���'wV8-4iTH��.]!���t�޳g��LH��;�~A�_i�W	T2i7\��0E�,	n�)�3r�s_./FMP�wQ�O.{P��0�[��G�T��:*"�)L�6��9ÜZޭ%0L�]�����+@��Lr�tmALAa|�L?��lMw^\,����{?91Y�ȇ�Q}K��'�g+��_+̔�@O��6���B�_Q�C��<i̾��XAc��f䚸̑��Բ��ڭ��"��0�ۆ�(W�^\��Y;~�f�za����k��yNL{o�%)��}u\#,�7ʟ9��4 鷺�^�ĕ���:7]
>����q�cw��x��ge%.4�4�*�B��~�}����e<'�\���uA d�H��*�\Q�-l�&���/���c `��ƻ�bYrJݹ�ӝ_6K/tm�]�r۝ci��¡p�3Y}R��;��[n�%�*�M���W���5�Mŗ��������{o���A�:�V&��1ʪ��ja�}9	�p�[�?���i�q��.���t�2���GWbs��]�U~��鿙��]��  ���\�:��c��1��BhN���s�#��v�g0:N���a<k�D�n�Z<��U��3��%g* �2�NS)��Q9�55}�/y�����<_�˅/qc��#
�꒎�ק,��1]c|�>��B�^�/9�{�W�p��`#�ڸ}�X�Fل6�O2���m*��%�^w��~޽v�]<��MvV	�R�J%��3�X�p�'n���F>�f6��
�ݞҟr���O%;�z�/�Q{n*�+�e>;����1���BS��) B�Lu�nԫ#{$~�����0�����.R)�膎���&�u4"r�����7p�h��,��Rw� "�G�TIZX��ư�0��h�c�0��d�9���nꦧR7u���q�����B�TB�$GK�?�*�A�8L4������q]r<�ֿA�5��Ys��
a�%[�?$�Y-}zmF�9W0�]$��(�5�&�����r�������k{�-Q��]�����y}pzr��Y���*��p��2g��Qm=W1���!ԈZ�u+��nr��G��[f������7��e^�2{x�Ye������N��� *�}gX��(ywت}~�:5�e���
{�3k1���癳��U!��s4ܰ�F~�P�e@�������t{=cCԷM%zΡ�22�啂:�gZ0M�7��p��f���;7	��h]H��K'���Kλ��^�i�n��^���.g��������Zxk��!��T��G�vh�����6%(�����Ļ�w�@�M�_ps���c�&�۪�S��ҹZ�0K:�d7w�!}�#/D�ϗ�G������n��h�K.}w�/���Wmˬz^Qw�.j��)�B�ۆ:z��K���E8�������ᬪ~�.��Q�.҆E9��E�ttcX��0f�����:� c�e��w)��u��*�u��Y�*#�B����K�����B�Y��oxbL�X=���dn�dk��2��t�������S�p8J4�#��	%��i8j���bx������LF>�t)=>X���탆�k����.�ށ���wl�r�d�G_���ֹ��_{]>�s��]��f�ɫ�s�7� �9+>�Fj�������\����_''�
m�^˺�op�F;����=�r�^��ftSz�*uu	g6��+�7�N�=�]_fr�{s��0	f\��c�J5;��}}�D
�yk�j�� ��I� h��h�j(�L�_;����a��>� F�j��^��98�jq�9ݹ�q�w��}qD��*�9��Zf/�hy-�f0�Zn�'~5��c��Y��^2T��:9uN]��u͵��� ;y����r�����0 6{U���a�9qI���vY-������?]+⼋����P�T��"��4�0>�;�8l�/�;�('�r�\�~��q-��֢��a�c��T�<�/�5V|ŗ��SZ��=��f$|�1�_eC�����Rlp`��K�df�4TU�ͳ~���5�j59�Ҵ�p��ώ�x7�g�>G>n�%脓��˝ ��F ���J�O=��ԭ�i�G�S�!e���(#�}��s/|\��ƽ>�^q��]f`{�u���;�.
�V#ꜫ�i��,7>��[���<"¯ے�法�Y}OԥIz�lI��MC�9�x�Vz�ݙ�|i��.��@7�������\|��%Dx�Z��ښ�*����`������;dl����Y8	�[nǘ�ThCB�h�PI�G;��WpVnԝ�������F�Q��JV�_'�;/W0�R$D�/]�ܛI��A���j��,Q�x�hÔ�Mc�u��=ΣnR��]���UUU��TL�7��r��z�q����5��]>�+��:���(�,Q���m��';DmZ��3�	^ݨ��p ����w�� ��ʹ���yLG\��q����ݍ��������7��g���,˯�Lb5:"�e�Ý2lh�Zw	����cr%m���K���#yov(�$X�z�`��XBE]��ADxN;	b;�r��Ӛ~cZ޴�wp�ɶ�;{�ͻd��"����ǄW�(�P��w*D��]��ܸx`�Q�:�'�G�:�#+�krO!�]b��Na�|7*Y��9W�x�O>�����.]�j�I�p�,��r�Ah��	�q/]D��J~l�gQ�G�Bj<1��@��*�q;+ǩ��s�������a|���n��V�*�f$!Q� \zDv@�6!�v���&x�Ԩ�|s6���}��_�T2Ss��``�����Se<��7@�睊!2p�IW�W��/�����_�zV���+���T%)�&�tz��/���+�'بU�;d�
�Qk�ʗ{�,n��X�=%������wR������$|͞�r
E��\��n\PEڣk�:[�5���iL�|��Fs��v��=ۥ��z�k�s���}���r���u������0ˀ:�����AI�G$�1�y6�-]������?z�f$��LX�ը3�YC������z�A��~�q�J��h�m��]8�p��Φ��K������ۆ��UV�o�����ƽ	u�u2�f>��MGNdm�Þ�Y�$`�+nϝ"ل7Q!CW�(�qd�a��]�[
���?n]\�i�����|����ǉ��P��2�|���4 �{����e����eWa{M��u�Qe�����>��*�GBf�pg��ۯuʘ�Ӑ���s���Q�CLc˳��t��[�"X�]�F�W:\�H�{H�@�Pw�s,������횋��l�>*酱ޕ/��{�束ͳ��Z:��q8��]�Aр2�
�J;H8-�\�+SB��S�W����]w�
^7N"tW�`�\%	NR���p.�x�;��^�J��yX��pt�a`3���|�?t@�0��4$c�3��z��O��%tuJYtv.3��$��h�n���%��C;pX�p�N���F>���}��P�E÷hS�P"��4�X��<�!�®|�J��wݤ�=�{���k+;����&�¨7
"'N:rl�X��e�����(3���Xͷ.��1�D�t0�z�\�g��Dܸ�4�I���z��P��Ƿ�C�h����$��{k�#HJ:�;�s��}�}�}e���=��&��3q/���Rr�2�j����q�`�sA	���Vl�d�T�Ҥ��>�~)�
�ά�L.4����R�#��tCG��o�ݑ�X��0���5��X�`��~�œ�>فlS���ih�l�i>�%���.c�1P��(��7k6j(�OU�Vwl:�*�fE��"c�H]p5�k�x!\%�ϰ���x!����kڗS���jL?��;,�9��w�U��l�ꥮF_�/���4�k�K���`�|-^��΂m���)��T}!i+�!��r���|2�Tt�b�z~V�*���x�rp&zPS��#�v��ц�����Z�3W��y޴)W�b�J��2ءX^�V��Q�u�zd��{�s�a#PTg�o��C�P��!��uLOd~�f�Z���e���D\��r������L���Ń�O�l��뢪y��Ӛs��|fzk̀�]�qŘ��r��F����YŎ��Y������v`��=,3�:��������9F��6����Z��+Sٛ�����f%f�r�iR ^;ҷ�"[�����l���ǔ�v\J��+�.��GC�_Z�9|��[�c�R�ӌ{]�5��;������"�ӫʖ���oY��ڙ�'�;'�ʰЖ����C����Y��e5o�hT�c�������ހr��o#��H����jnUK�k:�S�i��z��^>?l]f�}���:�"J|h�V�Z3�[_ l_EC����n�vB-����]#�n�!N�����-C'���]*٥�f�@�7��9�d�ђ�T���X�����4���Q�Ӂu����^��C��'��.Q�v
:�oqr@I��Jm�Z#�:�V�R�:� �m�F�e:�����y��;LUjŖ�dR��G��oRjA˕;�g���D8t`�@e�v\��ys�X���&PÕ��m�ֹ�o����A�J��+坊�Mۦ�[Z�1NcX��VL� ����[�i���X�e%���Q���cڔ���b:̇�T{���u%�˵v���$����Խ���ήe�T����\�`�CPn �r.�"R莇}YRwjW_�5Q	Z�c������;F��j��8f,��\��;F�pԓ8E,�5�HK�����C%��[�jS�	�|���JE�j��w�!B}G:�;��κ�{x�av��y�R}\���v�D��z�rXۜ�Ef�iu2:�H�����AU��f�W��
7����吭ȫp�E�+�&�s�!�͉�6�_E�ًn���o�e�7��IiUrEOw��vW3�W*M���L�W0���]�qwɆ�"'W��-1j�7�ϸ���R�{��Vr�vv�k!�I�����������)����*-�h'�#������[V�V�:�
4�P�]F
��>͵�.�˖�rv�G�u�8�ڵڮӹ�'�BL\a�{\}WV��\*t��U�9ӣ��з�� 0�[@v���SJ��Y�,�Lq����J�]~�� ���*������l�v�28�*`r�s:��3`P�6�g=��W�z��k�&��[`e�u��B��;H�q�QU�3���ҫh4�&�;3�V���d�iq�E�%��9�5`����T5-R��UqO��Y0��gj��a���V͗9���D�Ws��)��cup��،H<��=�����F��7K�B��tWZD$݁�;Q�V�u-Wss:u�{0u�tiZ�";�н��9g_wEt�1+xk��vK�s-N�Y/��n�f�<�=C��([[��S�����fn�Y�d:�$�q7z�{.���u���\iέ���Ysu�o���oWS��\�G-Q���"Z�5٢뷪(_t��T4�r��*ɋ�ٝ��+��<n�'X8�^I$
�x{K�ɵ��N:����\����{��79䬉��1�嘰�y���]/�9�%J�xڒ���NP������%��\.����]������߀�4�l%#@QN��AK���"RP�KB���SBR�7Y3%%ADC�@�M��QLM<��JPH�4SE4$CMRP#KH�P�%ͥy+���(f�
9��еJ�P�Aˑ���-PRQ�HQTE%R�@ECl����� J] �JZ
����#Hj��&��6�IU@ 1PP%%�'� (F��Ѡ���E%���t:
Z
���)�����4s8y+F�j�ֵ�)����U|EU��P��g7���^��wE�n*Z�wa�#��U$�u��F�8�K!��s��}{IN!E�A˷��`��BA'6�K�W�UW�7ܭ��_���4ۅ�
���p�?[
�R*7����<.���rb�Y�� 6×��&z�w:����X��S=�ӯ��V���eN��3�lx��<F���{yo\\,/�"
��+C�B��.Wl�p5��p�^4��'�U�U.�t	�����iU���'y/�{�R>��=�⒣KSۇ���p�����]��7.��g:��M�p�9>��.��$�IT��yΩ]���Z�4���й3���Z��7d�u]����!A/��N���Xm+�S����mn"*�����ϴW�i��t�$���]?�9�ԭyaqRgm�ù.��Ë�N�o���_a��Ȩ�隄Y�!th���r��^�9N&9w@ΆU�����*�.r���Q����1�*f~���0�z͜�n��75Lީ��욌Y;�%'�&Cn5��NT>Wm�����E�!��ԗ�#��}�l��5�,�����ɯ
��ॗ�_V��(�(�>��̀Jb_˻�s�w�����ŏ�e�8��۝7�ّ�x��m���҅�q�V�,�4U�V��݂�np��0!3xSV��D"�޼dV����DDh�v��$��·*�=�]��ŵՊ�'[k\9��`�+��n<a���՗V�P
�[�سU����P����@�9�T�>{��6����/(AS&��ХW���zu��K�pǞ*>�r��UW�MΦ��/.��ݘuwL����e�i�s�x���×�H�<������:�+;�����en-V9ŕ��t��Խ}��u�<�kg�*�eAW���F9��
cV�j��I9�U��>����'����|�>�q��>[�wH8K�����{*_9W���A��*9l-���+7�	������X�Vh�������fd��2�r�=�/�ґ?v4���,֚����hS��z;\c�ۂ��R��v�U{��f���S�Fo�1r�u�Z�d}�3j������i�0����[PL(�6t�[�!`pYj����qX�{:-���NG;9��z��|H<+��h��jXM8�W�`T;M��T*Q�{F�P��o�\�V�Aܯ&����K�iP� |�X�昩�Ї��Zg�8��t�^͆v0���N�:�������}���y;Z���mn��۾GnB}��7��MCrB���ö�E��	^tI�f��b۰�~�ҒiC�I�`���E9�!��s�7U)�l�����v�@�]5�2ؾҒ�y7��vÿ��Ꝍ{�v�ۮc�r�i�!�|:�
�5/�j1d�����vL+�[�I©I���ɛ!��m%�ں���v�f�Z��2�{��u#�s�ov�3Vl�Ui����6�)i�Ѽ|,��:E����"^eJǵ�N���7{Ԉ������?�ջ�/��sNx�E�VV�qOb�g(5�-��b���.3+R�Z��c�׵��L��'�Yg:�Sy�/�fg�iU�&��K��̩�ʈ���1��c�jg�Z���<�y�O �:NtN�r��+�Ys�b���n~U}*r�C���do>ldyw�����������3�YE����ӷ���i��+5i�ʊYxL,�Ǭ֕��]�K��f�ؾ� 4�%
����9Xm�7olB��#��Y���ci�|kZ�]��`��8Tȇ;]��_>\J��	YhN�8���+@q�3�DR'J�nrU̧v�
�7��7�p�n�]��]��\����H��]�}g�U�v�>��+R-M��;=����\�k;s�����Y��ke�W�_H<��=�2�N�:+�e�D�u���]+X�v�5v�cM=���Wp�\�;�����7�%�w!	Ld[���2�a�ǩTj��q�2ih���%ܦ�q�j��@��YP�#?fCoI[���j!J��q�Q����)�݀&p�����uv�hZ�P����'��f;q"��_v���r��Q����YY̸�㖃��7�iʨ���mO�_˷�t=\Ҫ�:��/�ln�l�z����l;�+��n��E�v�+\�D�ɬL�7V�BG~Oɓ �c�z�A��v��0�Q�:��b�z�ڀV����[�n�������ގ�^rI������>�Ȫ�ᚈmƻ��|2&>�:1ov}��[˂<�ʻz�iϳw*�%�B�#{;A���L���c6\�O�	l���<%�`_L]��P� ���3r�c��f�{&�A�����>ǌ`o7��I]�WV�U⮻qu(ug�*L�el�Gp���f�2'���*����_J>���2��&:S&�n�]��|�j�U�GS9�4,��Tz��(O�ۃ|8?|1ʓ2���8��|�o:�e����Y���M9\����c��R����/�3(��f#g2'�3�F�>w\��_`ZR����έ_f�iwz��Yٳ��et/�;�{y[�������N��K�eMA���u]���[�����ũ��q�W���]X��<��y�����u�y���{~������Bz�/�79��|�����]p?ܻ;���.n ����㓂h��^V�aK��w���}n��*�F�V�m��A����h��A�7�%:��*S:�=�|��=�|�ȣ
b~����7�uͫܬ���.��c~�U%>�s�We�-k�;c:����l�ec���v���uRW�u�S4��`o>���o��V�>���E����z�:Ld�yV]FoW/���p�+qΒfZ��9tV���2��:�8�]��*˭X�Bc��Y��� Cb_j�\�غwF*ּp.�ٝ�r����W�Z�b�4����t��b!��,�Z����¹WY�n(�Y��ﾈ�Qi7Mެ��#mn7�*�Q.��S%W|�~���f�V���]�fs-굕��;���ahHZ���At���B��s!+Z0��f�}̸�y8��w_%�i���2�]�Y�
Y���{r�+��e�A�Q-d�b��kc��Qi0i���*��woU�� Jh r�b�k��n�T+��[��±����饩:�Z�����s�+6__.������2�xm�}��'G*���*x�5'y˗�*��d��\���O���1�:��ľ��1焈�n�����__A2P��z�83�z�%%���]��O��k�������A"���{{��~W����mNwQ�@Js�}\Lv>-8�/_by���������b[#-�!Wd��Z�O(�{r�WR��'�tc��Q�˛�v�ٛj�}wi��6���Y=�"{]R�k�}z6dز�s��x�Kh�!����cW$�'��V�qh�,Z�R
�n�}�Y��$��)�q��hnN�u�5Wǯ�V�x�볠*.���
Q d	w_Im�������S���Ժ�ٖc��Ι��j����֯}�G�#�s����s���w\����Qʡl�p5�_c���4�&�at�:.���U-V�}[˷�9���˺�:~;�Q'������H��i���e�T�^9P�^X]��-�m=
�聸UD.��4$����2y�<�zl6�r�U9��-N���-k�5�m��Btݍ���a�3��x�5ҫ@�e�Y��U���J+���ې�觌�G���r/���
f�A�����ű���h[}�jM+5�0Wɼ��4�6�4ۇTk��/�r��R8-��oTֺJ۽�	���_%��&�;�;aͺ�k�����W���qӋ�ªҢ��k�����۬*��]�dQ/5�sv]\����-�ލVC�1qԎĭ��̸�O&��Z�c"*/��.gn+/�j�v{̷��n�59P�Y�L@�����y��yh��Nܜ�[)�=�<��!�����2Wu ��fJ�@�*,u�r���xs�߽g�?d���'^��<��ǘ���kpa���::�������x���u��u7,�X�\�5͙CR���Aj��w<t��q��v��W�����k�{�s�=�6{�ʵȽsQn�ۆ�Z�*�����U��W�8:�7��'d�c�X2��n�/k�����9>w�Y�ǹP����R������)��$Zf�`<Us���:1Fv>w������w.��)�n��z��ZWW=�.§ �s"T>�Q�1D����	���g2�Y�ۉ4r#�'�I����O>^|�ϖ	����C�lY{�1N�n;Ut̻o��y��4���������K�x���I�˪���Y���d�i~V�<�N����qCYc���{pU򍲶 ��$7!9=��"���\��9<�N�K)O9�X�1��|/a:n��J�p����:ґ�ү���?���J����ҕ�ac��N3j�)�Y��`B����sy/��_��E��p��wU��쀶c�u"�L���P�s wQ���u���m���\�Rh��p��u�#PO^���ͯ&zezR�T��sX��{�U�+����b�ݬ�YB�U�K��H�f�]	~rov�98o��\�����Y>��jB9s&��u��t�<纭٩+*���kfM��/�ǫrK��Q�+?}��DkTE���p��2�:��ARt��m���Q+^\��S����mh��0�G��[X���B<ð���k�Y����h-s�J잹��앛C��3�/g>\��=�z�tEWwx;�\k��&Ԏ��A��Ӂ�n���E�czډ3nS�μ��x��J����Fr�|2&9��[�SIs4��v����Y�ʷ�Ǜ���k'9�\9�t��r9t4*XG~'/ ��;��y������m�J��yίk�%ޤ�ќ|cmՋ'��4�8ӏ۹ʼoaxfTtf,���*'�3�F�c掅8ր����F��Î�����y���w�\���¡��<�C%e�2Ҷ����������/OU�\���骪{���ctr`�Zo��K�܏��kKQ���q.7hd���b�sr�=_K���I����8ʧ�
�/D�!��]0hg��Mr��<�����8��j*��L�o΋����߀ڵW�7�����O	ٍ.�(s����ꗹC�Ik�ػ��C31+y�Qj�������E57����6�U�wK������# _v�9o'�W;yJ�G�Gʕ×�'9���<�N*���Ke(�����4��'��Wˠ���-�[kI��RO,w���C����W������m�8{�O�>���yPmv.W]��}e/��;���}%:��5�_lr!��o�dC��y��Nm�jg�	���0ca/��L,/o���R m���iS������[�'�*߆:����<��tB���M��1�x��Qs}�b�Um8������J�e�w�8�o#K�ig�]�t�D�Z�P��¹��5�j^��71��%�{��q���-�f��>*���e0rK�9��[�R�MF,��׊㒣i0y��GF=%R�T�� ��n'k�gKPgS�и����/s��DOf�v�mGuZI�&o3"��Z�v�
[ݡ��늽������W�NU~�_A�����*���h�ٯ"��b��@�Z<�C.v�����&������A["k��7�Jv���C:���Wl�ZN⇬mb5��ٵ4a���t.�]E��r:�5t����9=�[���C��nL=u���
�J7�Zq�%]w{�f�֐��Ov&�L1PGH9�����3`�-�j��-7a�-��iC)[���M��̛�N����j��	v��5�CJ�V#j��A}��ѩ�6ep2l]8F�ft�t�r��-zk�FT�͚Eu�8ove��e��]�˸�4�rz�5��eH�8����t+m �\V���Ij
��Z1˩���n�T�Ak�<��#�7[\�B�9}z��zϞ!S��-�@�t����[.ΈS��,�7h$J6k��k��[ĝ�P���բ��&����K
��B� T3{�Lud�yX�6���MR] -�uͬ�×r�c�ܑ߮����r�Yj�#�4s�KB f�5�d!�P'���beb�ϳ�\]o)��{r|���|��Lq�X���v�����6�M̡��X(�=6y��ₙt���K�$��j��lY���<�<��ҩ"/��$�p�)nEt�6
ܘ棑$ͨ]�ƣN>$='����s�d=\��ĩ�BZ���4�^���s�F�X�'1
VY������7e<�w/"3j��E�)7{��n��'_n�u��u>w�>��0�������N�yDN��9;�lm��C��;Ao(eu.�� �t8�>mޣ��l��{��J�=&�-�k��ɉ]��;q�[��
Y-1[l���t0^�^�ol�E��]�����C0c=��R�/����{v9�5��;�hmCS�g"9���d��;�H�����lL�iG���sM����	���?ڽ��%5��s�α�Y=�f�X}E�m�ܤQZboP�qe�;�2�4��d�k�Pj���\�����䌔�5w�k�9��'aᝨ���O s���s�PV�\f���7\��}��Ge�';p��)����0���5�vj:7V�m��YK$��.D�6�ڛ��F���sq%V�QG�.��h�!�$��MW��2R�ta��eK:�Hg�
��e���e]4��o�:�PW;��9ד_`�=�D�	S��[}p3yE��s�AI������z�c�g֦��Y������//a��kQ�:*s�5;`e��u��#���f�y8(`��q�Y�V�7�1垽�L
|�^T;�6��.�"�u�]ê�b�:�$���3V,��q���wu`�@�q��d�������Mu�T��c"��'�i*�-��V��l�Q	 K�5�2�;��F�27���Z�q�f�� ���}�CƶV��ڱ'h60�8�d����m���!��p#R�k���ެ��YVz�0�iT�]�1dK3@˝/�&���wv�J*��~]�D���ԇ�PU-4J��E)���AE#�u@��N�B�Bi��
ZV�ѥ�H�h@�PV��!O%�4-<�j-!�O!t���^G"����P�J���'�:T��'Z�4�IABrA�(e4�l[)M&��ġ�JRj�#Q!�t�˪
e&�	ʑ�*�hZ
JZC�
M�)(SBh��t��9h9��:)��CZ4-�Ҽ��EP�r�ʇA@i(����SAHihh��h"MM	h\5TEU_V�5�X����2[���۫ڊ��Vm���G�Sggt�Qec۝��t���*P�lD ���b����Ⱦ�ү���">58Q�U�����b���s�Yތ{U�w�/X��f*���*Q���m����ù�X�آ~�|�����P�wn1c{Vo!`�
�x�N^V==:��k����_A4ulށKiũz���w��'j�t���C�8��r�pB���;������T�_o.ns�i�}�iWj���j�-S5	>���v��컊�:K���C���W���F8oe��B0���z�ޤ�Uo��>��m�� ���zr��!>�ґ*D��;ЦL^dev2zQ���po/=��Ol�n��U��د�p��K��ۙ�p!8V��[�'���5
[���������黈����Sag^L�]�~�-'=FouE���d�x��v���=�OʇT��nC.Ϊw3g�(�:���M�췿d�`7��жb�J�I�a淁�
M�>�/�/.��"��S��T+�pBׁ�䰓,wֱQtxtW�c�\ܱ��Ǒ���fI��Lwמ�\�V�Yn��'s@T{����`��[+�Y���v^]r�X]�.�,�}կ$����r��,/"��*$^�v�K�h���vb��ε:�\ϊ����c{*V�XNb�J����M�t��.z�j�Fc�b�0������t|?�#����%��}�7XO.��ᦨHP-��v{�V�����Mƻ#\L\u#�+p;��S��ٜwW�r\��<w;ڻf��'SK9m�͆�
##X��Zځ��+���w08�N^�ҁ�R�v�kڈ��W����j�#���Ue?c,���ߖW�z�&�?>�y��x�vĬ_v�Q{\��2�\$��k�{\�cs���Έ���:�tw��9Fz��1��Bg�������u*���Jz����8���r�Bꋯwrܛ�����S��	�P9��K���:�	�/��8���WK-b���r��}r�v��OV���U���!�D�\�'��#��%U�\�ec�1Г�M>/�z�ݫ��Q�@ΞzV���X�nf���繽 ����4Ջ�5���v ���ڻgs(<���X�r8���l�r�7��U�!�j�:��m�6�b[,�ǩ�ǻ=c��+S3WR]�g]��,72��<�l�;5-��{'syWw[8P����{q5��H<z�d�S7;׋�.����Ml���W�������ݽe���Bi�|���T.=J�.μ���sҋfa��Q%�I�w�S��p�㇝�e'M���7�+eLf$���Vo��pv���.���oK��R��[�N/+FoX��3���S�6��$�}�c���uѦh%=P�c�u_�ZX�.j�I�}]t�]�f��˥�>pWГP��RGH]P#H��V���|ʅ4�-����/�5;�un��|�x¿�����\|UB::�Q��y��#�;��V^�pʾ��1���ܺ�$�l8������}`��C�r��Kf��&�o����&�d�k�q�Q���mƴ��q��=���Ä�	��z�d/f,转W����j-�:g9����@���g�9��є�=BN/�}+T^s��]
e⋑p��L�5��t�Ȏ��K)�8��)�n��uf��6��3���hw%.�"���[r���׳��k���V{U���x,Fr�s��H��d��^�ҕ]���z�1RB��i��p�uf}��fڝ�VU���[ Q0S�Kn)�ؖe��
$���Y��kY.�ky5Q=���ǹQ�[8�.��Fb��ʞ����T��_Z-k�*�3S����)z�#�[�=����u�H9W����ѝc'k�cv�뽽ۦ�1mB������𮔜\+��y���-�;��H9l̝S�؇���ZNzUN��/�W-j\;O�\���{��AR��U��M��K�`p��{R_TD��P�R�����-S�.�4�z�5�����%g*�p7
����@\�K>��*S;S�|�ݾA��ï����77�瓨ʏ�[��o�nP��?�;��iW�%:��6��s:�H�bc��9�ˤ�q���5�k�m̮L�u�������{.mL'.hb�=lKT���ۭq}��KJ��sV�}��7��ǉ=���[����/m/D�2�]�����IMG�}��.�Ғ}͗��8�&�+�.��Y����4��tea����7eꎻ�Á���5p��4R�����a��R'Y0�&� 2*\��DV����V�:)9'�[���<hb���L�����fR���8a��G 	�q��q�\z]2.�js���0^���21ٖ��nZ��DMH�u��&���9t�Jܚ��;��K���5�.5��dF���l�E��˳+s���W���F%�=��.�'�b��x�)=����&���f#����	σ���{�U�tT5C��st���黩�\u���C!#�۹[�RګJ�j�s��ϵ�������%�WҰb��bt��6.�2{�T.�W�qSެ�S���ؗ&Z�$Ty��ݯQp٬Xuv�L�����P���c�q
e������Z��ۈX3	�wk	ND��IRՌbʉ���R_aq?v.-8�R��By�����"�|���ؠ��d󊰰m\�����qъ7��-�}V4	,�Y�aR�B]ܕVۇ���Kg�+�邺`D>ȕ���{���ڏb�iN`q����=:_��燶.q�g�����fB}:�+�����C�*g�lUlp<}�yځ⧽��yd��p�L�I^�Y����s�h2���J�ON��^��մۼ1��R��O!EBn�z�WV�ɑg�&�us7��:�h3Wb�⤠�R��w����$�ֺ˧[̙�D{9s?����ar��g�D31/}�ˌp�4�*i�ª ����t�cS3g[yh�T2��SۮxQN��z�dk�ڷ�*!:n�����
��3�:�qÁ��j$fؐ���[|���ac���E<g+�T�!���Z�덇��T��잔WjFŸj��%��-wp�i[�M+5�wat�7C���g�n(���o�:2��k-Q�[#�_@���ԭ̰��}�%̥Wx#�N���o%��7�)�X1�7�_�dKt�'���'K��;�=�݈*k&���INno��$��Mƻ#\L\GR;B��ve��}=�D`��.��.m]WK�[�4�!'SK9��h�80�~�sXɵ&�������³�s^��-�/mk�5��Gn�j����,U,��W��/C���x��u��u}+Wjw�ϔ��$�޹g�5�~�-�U�|11w!t}d^8���1z���7��F���*v��.�=H}�`��*#o=��[Q�Uv�ftUt$��h�}�����غ+�)���"��,"�6��e��Ӓ+�3�k�:�ӏ�b��c{�r��Q�l���I�;aή�}�~p�a����+X�S�<=S==+��Ss���w5n�$�i�{��}���7]V�j��/A"�=j���ya������7{���7��*n\;筌t�\K�ۆ�Sէ��wQ�_/��{�IZ�Vמ�z�)�p�����o���z�_=�����˸P	g���c9׃����}�et�O�U��gy\E)J�kwoCYx��&��|�nR���n����Ğy���f@�P�i	dI�r���)��8koy���o��%�[���~O�k�y�+p��9;��L�]J��{5��ac�Jr{e�3�o�3i�z;�cc:eN7!������"z�n�vn�Zx��EF^�O���v�.���O =�����C�C��OD�]��te�h�9:Z���/�4�|��(u�2�9GE�i��=n�#uy��X��e��;�Ӵ�*�v'��Y��ְ�kl����8�t*g����-�J�/1�N����#63�a�Z��x��%m��o�׸ن�WK��y3+�WQ���y�
p��fQ �p�ê8�p�3�tW^tf�(�s�NQX{RF�.�f\����;x>]'~I0�q�����u/��?ʚ�䛃�̜c.~<�.Zɨŝ���%Fӆy��̚zh��GL�{���C�����}R�*V=�յ���:�Z��C
�P�]RC����B��k"����_���"s|�-��@9�H�5K��w(�q�Y�{/}�g-xfTD39�X��3�뺽�]�4�OQM�Op��?�{]��p�Ǽ�w\k��W;�,�U��$�֞a��j���@J=��.&;
���#�:=����ƶz��t�"�����k��k�[��(et߆K��b�sr�=Q/����yM��)_*񳽜yG�v�y�FE@�4}ꊖ�Q��F8o1���xN�qBj�6��b�Վ[����:`��IJ���__4���h�2����/:�ƩfځWZ�8N�MPAe;�Ui�o-V��+x��t[ � ��{k0-G���:��{\k��M��ñZV�����&n��;��w�k�:���� ���ݐGKC�m���ޏj=+1P��>�r��K�HAuK�}/nr��^X]ܣ��Z��|7
_rߎ��`4��&	Q�3Ae	;>��o�גK�^zrƷ^7��|꒸�p:�_r�BP�65b.��l%�&�zy�h[��O.�<��-+�sV�'�)�9_K�iL�]��3��f��A�"Hy.���r��3zj^�X]1}�RM+�_ű�&�+����m��2�3��B�|Fm}�`��k�[�Q�w��9��pˍhJ35����a�ȫJr}����Ѫ����;%��KS�g�f�#{eWz�R����u&�$���y�}��U�2�.1�^^�^Ȫ�z�9�Nr�~λ)G)���bi�������z��[P6�����e*���	9_�zE��3~�c��}b���&�򗸜k_c�z��W���ˍc2������-�7�;���Q���j%`��QX��]��7�2շ�f�n�n�amqs'���9�WR�f����Z`���%�-RJ�c�� aݾ�e-V����]��{*dl��W/�%q��]7q�ǋ6&����8W#ݘ����������5q�M�}V<!>n.��:�j�r�:�L���pZ˅�-8�w0��nr�[Q�Gb�-8��K�����G4�[��Nc�y�-��kw��`�<�_�+��_q�N���Sۊ]Q�o�m��]�wz��ySϕo���P:e�Y�__T��;�(Ȟ~�����=fvI�U�hF8o-����+���U�\L��|�$��V9_k��!�Q���+�t��m�k���=���*۸�T.Iߒ%eut�+^�=So�W�M���w��Y5����]��3j�N[����Z.�݈t
���\��4��	����l-�zuJ��'�*3�ס�n+n&ݲ�}�r�HU�5��KE��n�iT�J��lY��d��C���q��u蟓<�8�F(oz#�w����Ґ��x���u*&�E��E���w�6ð��23<B�Sk����7�-�V����WS'P�&��G>]��[���Vl�)7� R=��\�R眩�}#�.�aun�����\!�m�9�n�zؖ���.|!e�*%,&�m ��w۵�Γײ��%�K�Ϊ�*VZd�|��SM&�[��w���w5ҭH�����o����eXt�eԡ�/��z��V+z���N�Ӹ�ڠ�:�=0�2��9��i��0^ðvd2�6���jDGX�٤��اb�<�0��
ڂ�>�(e6P`�V3,����9��9�'�P��㻴t�+���p4��G{�qw++�n����O����H�)Fp��Rx��i�4�/'Y��$:K0l����èp ,�6���`^����)E4<�b	0��˜�n�{��I�m�TD�֩��"�����	�3�Tv�$��vdo��r�(�,�2.߅��J�c:졗��VY4��f˔���h4�Y��ʞޛ^�����B�;�C��#�x�<!�Q�]�nYV����/�6�b:�&Uӧ�ւ%'��5=&>k9ص5h��y<A]�{���Ou�WFdQ�-]:J�!�ٴ�Ĳr�H���bC���I��3[\�������5�y��{��u9�ޕ����$�1��{{�1qw����Wb�/;M��T��Ŏ���̲�ko#�\�0�XXjq�V�O�޷��!ɜ�H�R*�,s鈑ϹZ�n1��2�sݷ����&j��}��i8�j��k��7��d�������Rm���F��丷��V����ͦ�Ƽ��+Kq7n����Y	놏RT�gu�U�p:�7�#��z%8/&ܶ�ڗ�(���_�dA���)ٓ$�>k%��˓��{g:v+#)�nԖ����R�N� ޻���>7Q�	){��B}&	�r��)Xw��㯌ܧ�듬�Ю��IF pu�h�Ɠ\�#h'*.|�W'�f�4��F7'�h���ĲP�k��m�իTvV�*��Km�H���]̭����▲����>����p�)����V[���8v
uN ���/��TytK�U�5͡����w+�QX��;�fo�9U� Y=|A���OD��}"|��XyF�5��b�q]]�����ڸB�=�9\z�)�IU�
�u֫���ͽ��$�S)�űb�7��(�sr�����v�X87�WK6������T�BpQx�\��d��{7��֝��Zr�� l#u�t����ӣ��*�o��)������Gpt�14坺�\��@��w}�g��7.�~%�q@w59`�T�F�:�m_ ,C{���PfC�&�ˋc.[���xm�olk�9�[�K �B�i��ϫ*����Q��ܢ8kw�ݝYȞ���M�wǌ� u:��^W;��N�Hım��A.�R��];�Rk+@r���.�z%f�W[N�eZ8��6��.�7s^��t.�%�0�k�7[�W��^�A��8�[��b�/����}��Q@|	M)ZLE���CN���444֫l���]!��it��К��ևBk@�KN�J꒴RP�S�"P�Z4h9:H�CBh����HPhM��<��JhC�6 Ĝ�((tPP��h��@Uɫju���ak�h

xF�Q�N�v�kG$4����P5�t����ѭ9�Ҙ���T��LA������KJ@�-�aJ[XБ%+@�i�&�
PP�F5�[cE��tJbUR�N��@������}����61�X:|�F2#0�-�Y��]M��=��u��n:��wE�W{m3\��0z�!J�mum�Z��[@���Wܚ�}˨��<��w�Y�c��Ka��L)���-n:;]�g��Q����i9����6�kF��o��"��<9+A���3��^^}/�Fj�٥����TE�Go�����a�7�C�mN���}P3D���V��S���v5'ϳn�'y:���7��,���֗�fE��`�|U���nr���
3��w��7��JmFϹ�{�|�6���d�}�o+�ft6j�����#�W�Q�isw�֥��1ϛ�:O��n�x���i�_P;��#Z����:��7�W�q�WlQ1}4���c���Ml�P	��b�}w�k���G�q���^��D�U=��JV5��z�z�i�|����ic����O�w �Ӆ�t��0;�DIJ��;��Ҕ��n8yU���������`�0���U�޽��G�8�����(���X᭹�_�`c�柗BI�����@�ڼp<� a͛�@Ү��c��u۷�;�f�-�3x�Αŏ��|;.�1NP��NS݉r�:ŁL��%��β��Ǖ�]���a�s���R��N������W��RvJ$4�J��{5��o�Z-S��8��kݚ9�ާ'��6��P����u��������z�-��®�S%m䨞�<�7/_�盶sZσ��le:�5�R}�}��M�U'em�ڱ�b����oWQx9y��a�j <a\q-�(3�G��\.d�T/��'^�u��/Q�֯�mo����i$ÿ�q��"[s���9;���dM��W�L�1;=�y�罯�Tj-8f�q��M�9�o/%��t��U;C"cP���e���V<�ջ�kb9:뿷D�f~�G^o+��R����S�3��t�}Q1W�o+�X1��=m��R�>E�a�:�M�}�~���9g��{r�=�g.�eA�L�Ss�ə�[9���v���+�Mc������^wF;��X3+�1`����O7�����]�����i%�����ٷ~�͟7ޯT�fъ�U"[�F���8�vKY�V�d�::{.,w��C2�e
���:Pʝ��M��w��{�������;m���"������'W8f�� ��[Ve����B^B�7���=k���n�V��t��X��8��1��5k�y�kw���+q����]�:�zz�%B�/�b���\������n�$���qOG=:�GS�v�n˞���yTI}R��җn��p�=��|N޴�p�kSZ�GR��Wp��p6+��TH��AګҔ�nQU9��5���f���{x��E�[p]�e/�(;w	�4�e�`X�9�b�K��g\�鯺_g,kTk����8�R�p5�-1�#m�Zu����;���J6a�-=���{�r�b��B}��3�.��S%N��N乺�9Ҧ�)˾��a,������U$Ҹe�w������c������n����%:KG��
�"G��o�]���sJIs����pdf�bh(�Qք�=���+u��\}��,v�=�R��n�uK�Zr�٫�:0�N��@њ���.G%=��Ɋ	�B���ي�kŏ�9�.����j�/�I��ߘ�=��=�����hʒop6퍇;�c�K�DNO���٢��tGF�|��w(��q�;,� sBNM.��}NL=�}Ү\k�u�r=�����5��NS�q=H�
[P��y��rzh��H��N��Ifsq�W;ڜ.�W����\9�j�Bs���f�5������d�h��pf@C��ҧR�6m^'{4�>�/o�w�9g��7xr���{u�������%�<�Z��74��Ĭ]�+4K���o�w�N=b�s#^_8��q�g��1�hI�T�c���ꟻ
��|�Խ|M��5�Nj���y�/�W�����%;롲����c=Q�ަqv�����%N��~�G�֪��O\W��] ꨒ����}Qn��nX�KʽIevJ���c7|�s*��yG�*�q�e(���NĎ�0���M۱�:�
���}q]"~�I޸k.1����*۱�UB��u��b�Fo�R瑘p3�����;V�QN�����-�ʄ�:�`[ب�.qT��%�@a�Q\tfu�en\��kG�PC�v�D�N��%{6l�k.7��`��:]�/lx���曵]ƍ���Tt�[6�+�MD��z__���,_����:N����Wns��h�䐂�̌����b���C�X���p�<&h�]���*��7$��w�}:�!����酻�J+����{��nu�I���3N��W���%�*��5��a��پҒif<��Hi�=yU�t�V%��K!e��p��9�*B����#S騕��:�î� ۘ�`�J�(ʕ<�wN��\6�;f�vCr{�]B4{|� K����:����>6�<�V����i$���k���&5�D�#���kU�%��6�n��c���ܪ�6j"��}�j�'SP�Ú�m��js\Q�,ꛭ���� Jѭq�!����=��KǷ�j��\r��\9�<r��OFms�\��X�s_Ԫ����Fbߦ�T�Q���s�2�N8|�uÏ���7�ҽ�t羝�W�Ꮆ	�OM�T��G9 h�e��g��35=���{�7���z��N�,�U��R�W��z��#��-��E��\�u�Yc�F��3c6�c|�=K;(J*��abS�f\�k&�r.����0����_�T�N�XL��Ci��7��})�j�2ۓ�����X-b����U�(뎎��s�WR�������2_VV6���թ�%�u���eBȭ�q;˛���v�v����C�`��l���٘q���u��-a	����1F�};�4����B�O�]�w*�����![%<������H|JԩJW����z�z�&��t��!�>�7�׬�����*��rw�Ȅ��j),5
S�h5�(���i��q�vY\������kE��M�©}�`�	D��_�+k��{&#Vh��(�)�C��֗)3s�{��՚��o%-q��D�bs����]��+�ϒ���3���b�s�pT&�T:�4T�_t����-l\8�ۃ->�<�i�s�r���).i2�;����j!U��ԡu�+|�f��cFz'K�'Y�S`U��$�l8��E٢��;�����KP�S��C�-��O&�d����G%F�ӆF���:l��ΘҒ��J�C<��?sʾ,fɮ�vQ�*�-�	n��?]�F�g)�ҎU,�D�˺�L���9���5�G]y�6��$�o���k��N�����]A=[��w؀�T��v� �#���ɝX��b�:�Z�������qޜ%��oT�j���o:��W��}�x�ڍ��n��HۇS��;��	�-�cp��:�͆���:E��ſM����8��:Z9
i<��]���s�2��'����^ǽl���>��4�7�­Q�m��D��5}��{�"���,|�L�/_7;��{\��d9�Zͩ%�an��8������]Q���b�]-8�<��Sݿ���ܕ�ޝ�ox��ã��X;�,��W����/�(�\ܺ��64��'%d������V.��Kg���+�r�����e+�Ë�����ܹ�,>{B^����@�9��.��'�_+�TB�:�}��g�Y�����|͗\/�)�n�5�e����˃[�w�o��v��«��u�_�/P�e��Ʋ����]�6ܝʝH�)]��Z�q�P�uI[:<��50���{vL��k�F�;��5v��]��=tInaU&�o��k�&.�=ۑ�D�y���yZ#2wz��W/]����DLfˑ�i$� ;}۶u��8��������x���~�����y�n#9�!ns�s�_.��I���!�q��N��)��b�6$%�6�c�nZL^�Op8���D�e��o� �KWPe�|J�aY�������Jחt�iU	4�������%V�pG�ߓ9�W��J�L�a��.��7+rq;�)D%�S
e�l�Ź�ڤ��t�c���VCr�B�x>χX[���N+�Tfb�]�Z�ܳq�Su���u��5��p�C�q1Ԍtk����L�&w�h�t��Q�;}S��J}�M{a'[k\9�j�o!�U�L\\���������Y_D����f��){�Ƶ�Y�Ǵ�Y�W�(�C �mo-�p�f�`fuD�ډx2�TMc�p�^���o�w����wM�|l��c���xr�c�=j��5kxM�Ԫg@���ԭ���duؗ3��\Yz���z��K��=ؤ�bc=h�yGK�ь�A3Jf�a����xtn�.�wkI�_�k���2!,�6hۮ�B�N��'�+A����Ϻ����է�
�Īq�z�̹%'8�;���շ9lY�r��,��*e��C���R�|����Z�D"�KI+2q�k�в���"��@�5[�
�K�[Z�����}�mjz���EG��y��j��I{׮��7tu�1���p��&�_���=��l��4�c�<�(SDQ+gT��bn��q3���R&;z�Q���ߏ?y�2W�V-�hg�SswC=�8��́,�Б���z�d�)O9�Z�\fվ���cK�Va��Ž��u׎x=1T�u�_�Ծz^P�y<��������O���RT��Y����9]T����|Ԉ��Qk��-��+R�%��z H�KdW,]�nƞ@{����S�~N�!Ϊ!�Э�Ek�2�ʎ����=���ֶ�]��\��M�lS�ȟ��)S3�.��T�9��MP�in�t�$̹�X�w����i$����o���K}N�|wD�=������ZJ����b�9N<˖�j/�uZI��,p桷j�<�f��q��tr0h*^��W��lh&��}{ �;��r�}�EG��\��^�:�V\���㗔�ѨD��
�(�`	�|����*t��R]�%�"��5�8�jm���d����5t�5�%�)���s�.�C��#��+Op�
�j8��t����*%c�Օ�IG){p�Óp{�S���=��RC��yM��d�-��m��J���ju��١�~k% n���j�]˝�z�ǳ�L��H�����w^�n罃,��iI�fe��*���rP�{Z%8E�����u[�y��a���u��J�Kմ7�s �Q��c��q�ϛ��u۶�*����V;�e��.���w�9U������_OBꁒ��(��i�����_Ǧ�-�=���o[�/^��ߩhwX<�$��m)J�kwqCX�<I�W��j�3r�{���b�v�_�p��-;��q%*�=��,4�<M�c����e(/,.��ծI�v7
��ӯ�����J���S��C�Ӥ�wK���nu�����'�m���R������a�t��וTT(�Y$��k���t��Wq[�@e�ֈ8̣faAmjZ]��4��y0jᇲ��t�v�{��z�S4rʸre��K˛š�;��Wk�P 䫷���)�dƍ�m*}��2��B�]O����fآ {�
��;W[����;���2���%��.����Z,��B�;�an�@�e2&P�k{#4���V8�vp��5]6��C�XyYrړC��GK�� ��gm�]��J���t�2�9�7;�Z�{���W���)!!����P�V�9���7F�*`�&*���j�m��>I��3^QqV�{r�m]t��o9���*����+�"Эwfo$�����dV����썹���x�IP��B�uĬʹ�vʅ��N��E :\{@3%b��L�:�{*�.�IsgG`�{AlS����e�D�u�Չ{���IC�CEc�ʋ��� ��J���YXv�Q\��ݰObJ���b�.���b�\�u;�`�j�v����+\��Y3Jk�1���V���2��;��
�9�M�[�2+:�-;��:.+o�OJ`�g�vh�m^���|Ma�������뜅�+uW_%�VJ�r��΋���(uL=m�	sc���V�������S�2}��}j�ֆ.�c��w%*�'�ԙx��	��nWL�6�YZ�v����7�|��si���!�ĉ���Ss8��J�S�yDda��{��G)��P��VV�O�՚�5�����ץ�ͼ�LLzDg2Gj��V��>��-�jC)����q��N��&,�0�:��Į�G>j�lm�uu���"��4������
Jc�QH�1f�+�;9M����|�Wod����v*��­I`�s%k��ݞ�7Iҗ�/,��c*��>�Nv�&�
��fs�-h�}���)Vj3r'9�:���ӹ����r<C+��$�V�:U���.��(H2U�qV2���+�빜.wp�5��N\�M9�˯���۫9�e��1��w���׫��yg��������Q�ݼʾ�\��i��z>��Jn��ڝ��t�4��,u�Ң�\I���Z�r��U7���b��>̂�d��[�S*S2�u�բ�8�W>CA׋2��]h\���+}׸Rxg[+)qH��Y�.=�:�I)F��k�Aیggwvv�G��+�2� ��ZH���Y�V���)��M�WQe�|�L� W��Y���wj�Z��I�F���L���Ds�b�o{��\Ⱘ�\պt�9�2�_B;��.]��[�hBjvT/Fk�	�9B�d�ұ:�v8 ��V�s�T�^%P��C�u�!+��Q�M+֕5����4qڔ�lT�{X+����Ľ�_ڀ�cTV-e��O�ӫ���J�L�{i��t�kO5�V���z�54�12������ovA�̅ 3"P����;`/sJ�Ʒtd�j�SC��c���r`�uhI����]����W�>"����A�4�5�i]c`�ƚ4P�E�
��M:4.���1$lh(�i(b���i4h�6)*$T��ڗN���1kKCBiF�E���5����)(����ӡ�-CTPiJP��КД�ilm��6)�WN�l:�P�j���
����@��i�ti6�A��PPP-�l���6�M:R՝i���*�����f�4i-�QZ�m��!McfڃJSHPDDSE	���%�D�Jh%%h
$M��|��w���~务=K�ʐ���!�ޜ�d���Uך�[��e�Ɏ�]��<jk�V�3���>����˸ֹ�1�rڥ��������|��p�kY�
��ʗL�Bΐ�J��'U�-X&�"�k��p3zj^�\@}1}�R\��/����:��Tn6��W�Unt�N�b�q�f�SV���]�X���U˨��&�.5��0�yk���͹���0�
��;�ڀ�J���,��^;��o�S=>.R�7m�L�dwf�*D\�hȞc�-��]�����SN���֬z���	��7g�k���t��s�3��H�ј�鷃)�sV��{1��w�-�7W���S/-'�w��q�[9p�3�yE�tF�:�om<��%��q=;_J�ڢ���S<�Խ|������/>s'<z�cks��`��xX}��|=��Z�T���z�΁���_ܧm��i��񘷜�������O(a����[�qV;��Qg���|�mP�Y��@V'Kޚ�D�k����3댙��0;^�Gk���.���`6�\�u��T6�Rv�s�J�8*U��V�a��W�n�61⣷�KfbaU"%~��z(3�ؚY3#7����&\+�ӎ��Gr��ge܇@�}R���U�A�l�6��Pv�!F��2���ك�����W? ߾�l!�>�Bߟ]EQ!�FUC��>F�	��,9���7�o�ۜ��*�����#�ۑ��~S��u��� ���.�r�%TD�1ʡ�-�e��#�b�`�7Y-qD4}��M�����>/K�H���|=7����Â`�Ay��5���^s��S3�(O�;CFB}�h�w�i��z����ه��|j��.9�G����ǀ��:`�|zW���-�p�_z����_�l?R�n=���#(���y���Bwt��Z�J"�������q�����pL5��C����"}:���=������}A��}8�_�%��FIh�$dK���/���C�ԍC�>�]��fcw��C�����:�޺8��[��ց_{�~�s~���3�l��_N�ߪ_�њ�ULԷ/*�aO7Ԧ��ϡ�ۆ������2o�{�{ :���GF��:nX�����Ӊv����h�ڏ:=Oԅ_ٵ�7	^\y�Ui���Ez���<�R3cʎ�q�ĥ��O���Ǚ���<XD��\d���R���e k���k#��aQ��d"k�^�}�����d�Wa�Z�m���j�dD�>>��E�x�Z�n�n���>��u|��a���U֔�U����m�m�/���cy�p��xn��m�vrn�]�Owb�Kk��M{N�gI͌�C��V�:�dk����׌��}|,O���國Wz]ο)����ǉݳ1�BwL;��q�t�]l{�^gՀ�����6�iSU�HT��N��9X;W)N���{���ٷ#qΓ�pf>U����q��U��`�Q��@����К�:�2��#ʩ��{'�%�.7κ�Ϯp�4�g �T+��T����3�f�r��'�uFzd�^.Sz��g�T^���~ˇ�ʣw����s���E�$��aT	���qW���r%xv��Y1��<��Mx��w���x�
��~++��ݐ]j6�Wf� �;i�y	>;���Po�0���z����I�cc�I�}nh��<���1��:������nM��3�q�7�k��^�>��$�3�H)(�l�(/sǚ(9~��>G��þ��4"�±�%����W��^����GzmO�}��[�*J�U�	�Ʊ{�&��X��w�2Qu��+������[;^�W���p��#o�wlW�2}=� 9����~��p7�/�� Lz֑�Z��y͡Z�9E��X�2U�ƧP�BX�I׫\b,�r���%������=p��"�	Y�3���g�ր�^�&]�$�k����~�ϥ�u��&H���;x� ����-
D��������q�m�x�.m�J:��6lAȝ����FP��y_i��F��"����w����#�;��:}ՠ�?z��U��˪%��T��� �?R�n��4fE� ��#�����F.5�W�/�ȟ��>��@����H�s�5
d�������p�Q41ǣz13^��'��t�i������C��ܘm�������:��� l���ܺr��
�F�m����.���P�a��koFDW��j�ͦ:�+�7�
���n=���0xݓUnj�2�fz�{c*A��d���;��w��ݟo[/:��ϓ��x��N�ߏD�YK�:�y]N�3^�uXSӉ�
�":|N�8<�ݘss�+�/I�k���8�x4x@�߇L�����KC�S���=U^�r��x���	[��el�GÛ2����wYU�b��{�Od�{%wWo��	F�P<���2�@_:�w���IM���>ڞ	Û2�F���!2#�7�ǽ�\ט~��QB����7��`+�G/Z��;��J�wެF���(��K�����h��=bk�����g���h�E9��4<�]@�=L{�����!��{˿L/�]v��q��.Q6z_tڀ!̄��N��`cU�LW$��op��+�&]v%E�{>��nSs�5��̬"�#ڝ	7.�_f���x���9o�u�܍��_b{�C���<��;�Y��mS�L��jxT�/&�BCRw�w�M{^�#C�<.>�ʦ."�R7U>	廠�������q��캲o�j��B{W�_�]��Z�}>�A�d�=�(���@�>U��-���Ax�yQ/|�.��9R;_I������~\}I���}@{�yI��~�Ӳ[ ����a�!�b�5sN�}{o]������Q^�W�#�\���4��g�dm��٫�z��"����$�`����\�l�1��|j�pn}M�~���#�p���\���ߌ��K=���u��q�٫�z��de�|���Ӟ�܈�b��!�~g��ώN������ղ[���2��ER޹�Jd�$.���F赳W�ǩr��M]�mω�F�*gKG6����pͼ��X�������pO���!񿏲���n��+��zk����긮\ٟ�C�G�S���'��t��~�������p*��Q �|o�;8�z�M���G�[��(�5�2�v���{Y���n'�q��Q�����H�993O���0�-����#ӥɞƊ���1�C�u s�"��N��� �
m��r�|�q�h�H�y�|�!�"�u���d�YeV�Y��н	��]]��k���"R��R�jwqc�iRL�}s��T@Wp`e�ð�4Qf>�JĤuDH��[8T���湭�d��:���C+�g#6_�u*���S^�ߢ��o��%g���n>��s�t�?���~c��@�"]D��)j^���çF��S�t\E9D���{�Ꭹ{ 9�o�(���]��c��lӞ���Y���x+�V�x�;�fP��Y5�Y˴��Z�/�^~��<�
}��S��v�xs��}���Ϯ��8JWa�=P�+�H����fG��r !��oݗ�����g��9�s�w�և�d��-���TQ%�Ѩ�*���2̞Μ�3�¶tT��	U����>c��aϵ�������9��ׇg���x:vK�r�%�G��m%R��*פu��e����~;��}_�ȵ��M��~��'������}���g��t�m�>�X���Ϩh�#r�#���0�>�}_��RU�7�hh������W��\��wl��[01�N��Ks���4Οz	�@� l��5����/_O�0�ӽlv��K������u�P1����-w9��D��S�������D@j�H&
�u�����0�b��~t��韭��;T 8du�g��$W��g6�U�x:�����jM��|Pi���Ma&���)9c@�9��ٸZ����`�!�g��s�ºa���i�ɽ���Y3X䩍������7h�/7T��r�Y|k��86�[�؝����\�BT���^�Ks�w�'=ӡ7��.'�쉸uU�FIh�$dK���/���P�v�W/�v��[-��G{��Q��(xK c�u�W�w�m��f*ϑ��D������)h�O�sWM)�Y�67��yQ����ъ_��q���@uCo�*8EB�T�|%Fc���>�&-��r_�_�W8�ke
�����7�1�>�W��zX=?�~�a�RS+�J�}i��{*�;:;�̜��ѳ�w�+N��:N�ٴ��3��1�׻#5������j���p=}�����d�yf���8{mΞ��a��a�Ee{�ӝn[ U��c���&>�%c�"�����uJ}�F�Ζ{vWL��t#�uآX]#�K@1`/v�x�z�3�nf���:�S,k�����п�κ�ȹ�Pۉ����T+��R:���y���C�m���2��{ =>���F�@�N���~�\?�W��vy�1q�:��%tL��/{��#N��ѳ��2Inc�WH^���׋������������W�ǻ�F�J�L�^b������o�I�H��[N�k|+�sf�Qxpo}[�*�/b[�2�2#Z)׳	�5�y4��o!P�+�3V�����h�{/�Q��]��k�rܦ����3s�n�o�,)&sv4��8o��.���wi��Ԛ�Pj>YS���V%�M�{�A�t@>��EO���i�[��[�c�#��7"7�<z���{���
+Հ��rWs�0�;j|o�Q'�x	"EA��d��!��-���^��={�>��Jf����^�������p�~��Dڟ��@�-���U�a�^뉭���P�׫�R��������{ӣI�zdg��v�_��Q��̀<树�7<��'�{��s�Go�],��_}����~��zgx��{g��^�q��uD����� ���w���ݍ>��-('�*M��= �Ƣ1q�vڿI�~�"|r=3�'�� ���Hp�}$Ԇ�̘��j+�!��%ߵ~!?��
��qC)zV�����Hm�wF~�%?O�w��بʙE9�"�f��`{;�hv�x��RW��.��+W��ތ�>�W�f��U�:�������[p�2_�+3�y$=������.d��*�d��;���6r��?���xA�b�����k���ڞwv�Ź���8܆k����2:<�v=+o�8������U�������1ߴ��$�g�tԩ���ye�f��Hd'J\���Sq��.��ﷺg�y[��ަ�x���a��T���{h���خ��6j�ǝ����%)ؓ�e����FV�>��&A�Me@{�KM��Xw7��u�}�Xmof��&h;�H;]13ʭ=���{���<�_�C��i-χx�X�Ƿ��{�['s�:�%�8�|�i�׺7K]��}}�b>�<�f�g��TyC���C�Wx���K!Vq��>ڞ	Ûq퍗��t��i�R��i�맾�~�,eԺ:.���i��k��K������^�Q����0cbcd�MO����ܸ�9G�E�%�̡��𸩟#qNC*�l��u tb�S��~*�[ ���v�3}>�ʞ{�_sW�<v����]x�YD�Fc��T���Fd�'�� w�x3]�_�ع׵�;Ո%�U�4w�tC�z���^RmK7�K���@��Pn"�P^"'��}����y���]��;O
D5;���甑��w���[ r�O!��P�>��<�ڱ��{��#مQ��z��W�;H�;��?H�מ��������z�pB/sޅE��o����C���g�⠁���_[���:��c#ӽ~gO����T��~2&�tx��Ν�f
�l��ѿ.IވO�����N{�pQ��;��~dz|���N���fT�xb�����,�`8"i3�n�{3W}r��F�]C��N�;��o���2N�m�t���t����N�|�i뽸�Ǭ��`ǈ���6��y8 _gp�E���!�ݧ2��u ���=xP�|ݍS�L��ޤ�qp=���o��*M)��=f*_W���j�e�W˕��j�EF�j7��Wջ�^�������x��@w�*�*�'z����}���NQ~;W�JSE�z�������3^U���=�����Q�_���f���CnD)�*�����};��_������I�3$�\5F�|�j�f�Ѫ_������~�E��Q�T�:�H�}�Gfn�|
5'�d����nU���{c�����T��J�t�l���\<�M{Lc~�^;�	����o���ӄ?�O�]f]ea��5ͮ߇��^��_��(����������,�uK�!ׯ�V��a*S�Ǐ��������z���~�nm�9���;��X��&��9��M0�@��W��yRbT��ٹ��Vc��s/�xn�}	�!{��H�Y�R�0�ў�w�z�����l��Y����X5��1EV��g�w�5�=�+և���?>�
�$��%�_UA�:�j7r�lf9G�@�z[>��d���{o�x�s��������yh<�;%۔	*�g�Q���{�����J:��4~�ܬ�f���9m�Yu��K��xbBh|D��)'��6��d�!��7��n���ol	��R��b+4�F]l�r�+z���p��r�j �ڗ�˰m51d�֌���U
�F�8�t}%f◔�c����q��8^�8M�mBiMw�hy�iݐ�Lްx����6y6�-ɽ]����m7�L�����ۚ��\���h�����\�t�\�ra�ͩ�9�1uIՙ/b[S�jN�a�z;��b�G;�&ˬ�ԩ�N����.	���Y8�Y�
N<w��H
�s�@�m�;�/�
��'�*�#Ò)��*_Mn���x�˧�v'�ٔ"5ڰ;���8���H�=�:8iuc��J��l�.i��
���db���y�Z�[����],����ޜ�Rᖚ��{��<�W�gD���7��e�-�]GWČ��Үن�s��9ձ�7M�k}���*{5=#�q��h��FF��)Y]�$�զ��=u�($�ʋyBMex윭��{w�z�6�*���R�]>8���@)�e3�,���v���s�/�5�ݹK���w{���W]��2D:�e���������r�\�N�
����Q�w���I7;�^�DoCMv�t�.eE��7G����
ǁ�m���g�^���Y���@�6벧'"{�d&>]A��<�w��d݊ݦ2r��<��򕹫���:�7C&
u��~�^�z�Q/9�{�Lj*ot�!G7��	�`R͈n�\:�}/j"�]l�R��xqfwo���Q�<��>���)��HrH:��|�g)��m)9�_L��+t��R@��&���#��S*�Ο27h�\K��-�lu]wJ�m�ӑ�޼��>���=��+�Ǥ��M	ˋ��o��`H6�QT����]� 1,]b�
�}R%Y�;�n��!��|Pn4�Y|�]`Γ��g
7��z-v&��O_;{�=�mi�m6�e�&�O0:�j����s�oV�i_3�A(�8�v;ה
B�����"�Ϗ�*Vc2ms�ym=lf�ڇh���ţ+r�	v���(�� ��n�hx���)�C���;]M�ۛ��Ĥ���\k�n���⽧8k}�^�zb73Z��?���Vʋ%X�)�Lo��FT�ʕ5�yx_L9���[udx�ԥ��2��6���;�����)c함�me١�EM�w�#|e��x���9����W�[/_\ػ�5s��j�Q�Sx�Ε��=b�һ�:n����a����>���ݓ-�*=�,=�Ǻ�ٗor���䇹�;.P(�t}g�h��E�)�)u�)�B����SW��Qv�����Y�u45��+6�:��#f�rC&���ΦU���8�_f��/������l7�B������m�W[��o;�:�0]<xl��)Md��c�l��ؼ7����{Wػ�rbu�˻��w�������̆�5Am��ED(%P�ɢ���())-:�Ei-�h�&�h4`���R55PkKUA��V�)tSDKF�T�,Q؍�STQDE%QU&�[:J�����+m�:*�"�:�i�*��j�)���(&j����(�����B�C����h*�b��Y���:�6ƚmf�*f��H���LTTT�:L[f��)�-m�QQT�S�MT1UUE�&�PTS�QT��AMlb�����Z"�bj�%�1LAm����5Qm�b��33�h�+!�5�9��A��ͻs �%!`��q�]qn���T�ޚ5g=kl�Wom�Rgy��M�*sYR�d0(��G9(^fmuk�-�)�>W~���OR�ȶ���>w�9�'����3����ߏ�����O"}E�'�(�.�c�Uz�������\T��J�&�Ӵ4d'޶�x�:�޸;^���Q~��h�1[밯�����4ɞ>P@L:����^SY�,uF/_�W�����c��j��Y��#O�\�G�ȟ{]��w�rfYߑ� p�+��n����0�F.���{*&N�G�V��.�x=Ux�dN�oޭ��_�&��zfђZ7zH����2��ӯ<,�����Od���w��Ͼ��G��~���@��׀��z�����"|�F��7Q��Y�蹟nxOS����oO��w-��&���F9~&O��|�:���GF��;W�2Dy��y����ߤo�N�����
�i�J������d>�W����p[���2���3	�6��Z�Mw�2��t�a����芟i�q�I��C�3��1�'^�~�ޚ���ͣޑ����J}��z=���w�z\?�o(�~�-��Z�C��l�3�{�~
;ϼ���3��Va�@�ߤV��Mß>�����mw7��R���������p��׳x�"�$V�;a�D��;��c��nu��kX���e6���(����U��.��-�M<֎�&�.��v��Yݛ�Cb�h;�k� �\rJf�c�}�*kӑ�4;�}�k��yR3~s��٘xG�Û�ô_�M-�t=����;Wܽ4��w���ʽK�d:���/m�{�]EQ�P͉���_u���
�	_�٫q]�9 揢��o�;.�����x��u	��y\wdy�1{�t�2ԒV퓜����p��r',���wS:�%�����^��<}�������dAu��}�.���}�:���1��5��jH>�3�O��X��T���s�[�o���z=Lno�x��Y�Sy�=5�s��=凳��l�1ށ�RͲ�.��0
D���[72��|����A��ilw��{�{.r|�^^���1�M�_�=�����:�1�$�@Q�^*�����
ް�_�g�&���sr��]�����?N�%{}R6�wlU��G�C 9 q��p9��Q~�=]����g��@�l�.5�o���L�x���Z�?z��U���.��-T�����[s�����Ms,F_Ru>�px�b�P����M�����o��|h�׉�^�?���x(J�q��٤-T��4s�<ޥ+*�	��KϦ
����m�
kھ�6[��p2-t�t�O���"�|���Zb@ˬs�.ử'q��e��{{����ԛ�ǐIEawx��rt�����m6�w�D�x�s(�3�	�"�W'�G�rDl���a���4'�a��zk��CmUQ�m�̗���=��%�����t#�蘮�Dm�I��\Ǻļ1Q-m�}��3i��J�������w�+ޖ�{˃]���x9�G�P�ȭ7ތ��|J�0�D�w^��qE��g�����%�����~�5ʷv}����w�x��Þ��ޚ�yr}>'``�#2a�ey�Z�p�³};����ڲp������Z�2!�W���n��w��%do�4_���ulL�%U��prSHz��� ��*�2%ٗ��\{$���:����K!z��NmOYx+^����{υr���:�U�S��7��`+�k��ּ|�����Z���{��C��m֛�o���}�cя���>����ʀg�S>FY���C���*1G��e������+=�6��L�E:ap��1�����,�J�1�k�*���H̟���a̦t�q��߮��j�)F�����r=�G������PjmK,"K�1�,��^�}�S���Q���XlY���fY�4���$z�Wa��t([���Ũ2�/��h�F�-�ۛi���,ќ��Ώy�e促͂+͔o�͖S�wOKůp�J�
�E�n5C�Xg��)��U��x�pbM�����fї˭���d<��;���K�:��ND/H�ȍ��7�Dm�]�{"N�v� ������'��'�r>u|�Y�uz�K��2=Ǖ���t�#����;�4�{�Fz���9�Y�tWM�ζ}N��<$�@R�|���|j!oW��ُ�h��{I���\�"���`�&�	�o�e�����	0
jh]9�ρ�U��;�W��}���*�']����]��#�"n���V�%��(�(�`��Q��M(�c˕���E���ꑻe��oW�y���7���4
�x]��t���2>ʊ�պs�/�k�Ȓ�x�����7���\�YHy�W&�������4��#�Cn|�ĪC�pvp3�/G;��7�`ou��zt�"��\r;��{k*=���ސ=E���b{=��tvf���kі�yeE��,�1��)A\VRqR��7�+��:���S^��'�^���V~�}����{񉨻OE)��vG�x���X[���늜�����],�����T��2z��,�[s��Feȉ��S��].�S�䶖D1m���t9Ǉ9f㘯���|�ަI�n�}��ù�[��+�<��}9RŔQ>u��5n��-�\�b|6����x�u��=�s��e����M�e�<��.�\��X���6���&����
�]t�.�j�����u�1��C:N���yB|��Zn���X��N;�z��\�P�~;Q��sU���=�}ʫ���ׇq�{i��>�G"���fza�z�� 4�Yίm*~��v�rd�r�귽A��J����^���)�)�!�"^����,��IF��Ѩ�*��r����n���A�������F�Ux8�O����<}���~S�z�xqwH8Ӓ[r�%/W��V����]�(�����3�T�r-��/�{O����[���W/	��Ȩ��fE�/gW0��p��Tg���
P4nb�e��%^:v���>��v;�4�=��Ll�sT�W��/g�o�z�َ�����p@N�2H-�(��)������ឯ;bVՃS�稪���V���~As��}��\N��߮*�MK7�T	��z���|}�a��x ��EEH�}0��3Ozws�8{�%��Ͻ>�O��G�~����K����2KDq#>���$ҳ#�ؤ�/ 7�@���U��j5#P�W�6��@�#Ƽ �C�b=�p��3�)�#S�6d�c�xd�WQR��=�'oB��b��`��:�>�U�X_+꾛3\n����M��ȹ�
R=�'�q�+�`%v\�Y]���S`��F[��o4���ͱ.Tu�{�U�c�q�=9���6R�wn�R��zũ���3�S�̧�N �|�x�θ�#�@�u�1��m1RR9G����x���F9~&O��|��m�Q�3�BeО���;��{��&v}��cӁ\EJӢ}��]�O��W��Ui���7�z\���Ҽ����P��nM���,�P2c��և'�plS�'se^�Xa�u��[��l@��/���s�=�H���|,_��s����=�s7Y^�t�Aۅ���e��/Vް�W����u���=�^�<��ӞSC��k��vm���Γ���yL9��2\\����,��W_zS��{��\���Y�K�d|�;�u�i�������K�%����tA�پ�Q�{e�ҍ/C�R�f��#A�p�tG'K���~<⼮;���_{�t�=�ί����Z�=S�S$�D�
��qS-L\S���>��y�^��P���~��+��ݞ�8�ǧAͱ���xo������f� ���0E���H]T�9ϭ���ǂ�G���f���)���:/؆ε��>����՞1��R����:H�<[;S(/cǚ(;c��C�A/��i1�3����]���c{��UΫ�euWs
�H��7/����'sj���A��Ar��]�)d�����=��Z+�y��u�]�x�:mwV�<mԭ��U�gS�蘶E�x�b�8�b����ܒ��'Ο\��>��v�B�i����'�?}W�V�z���� t�W�<��>,	����J�U1�n/V>g���}v���ؗ\J��^ב�~�MǷ�#o�v�_�T}7�<�{=.u���@�^z(��g�go�&\fD7�l����}ՠ�z��U_�\K�%��*�6֡�fΛB�w���̐ �}��%��� ��ơ�6��_��>>&�/�h��M\�D�9悥��������}.{ƅ�zV���^��I�Wtb�~�$xv|��p&��װNj�=���ꍊ�*6@�s�=a��'�b�����k6Xބ��1]� �Z��=
�	#���=��L����y���FT�Q>%Pɇ�wL>�V���e���b�Ӄ=}���OC����Ȅ��z��^z�9��zhW���y�GO���F���;te�븶�^���T�Ԡz���NB�~7֯�U{Iϛ��?%�_o���2�~���`��@��>o�$�Z=�������ɝ;QH�n6g�*!o�ǲL����?eGw:�5/�]<u�~��(̻�U���8�=̜��b5�^Ǘf���6��%��k�0;;�6��wOa-���t%P�]GNn���<��T��L�+�lr���D��Н:jΗ�r�υZpVwV-+�h�p�j� � );������vۺT;NR�>�Sw��\�;�Ԡ��QӷT��%���:-�ܮ�� �]@����=t�T�����I������>��}�F.5��G,�)Y�2�x�$��!�cf��w Z�j��"g=�Oq���ER��ֆ�z�+"�H{���a��W���#QU1u2�����6��3ƍ��f;V7��r~C�T�X?7�w} {W��Ǹ�r�C���eX1�,�T<��}G�9�p��GM%Cۇ�T��k�q6�ߴ���<���ߺH��w���t��9U*�m���1+��z�>�<;�x�*���W���C�i�x�/�a�}���������}���y�پ��u��}`����}Q2G����~<@/�.��RF=��l���l_.�dbx�����w?�߾�w�E�1�TH����?-r���\�A_�+a�X�oX-z����{�SX��g8���2{�뉸f}&�L���'��}>��E���ǽ^�q���^=�1d��Ȕ��n��=��\&���#�|{"��*=�wT�=��|G�c"_V�̏wh�s���@
�*�5����ɐA���u{��}*�Ncv�r3
�u�������)Q �ڒ�+�7�Mmdv�	T�-͗�V��K�v�z*ԄAf���OR��[ri4���;�4:�D�Lt�J�7���x؍�s�u�@87����_�ί�V�[���&椨���~��>�f�ߐہJ|J�t>!\k������s5Ӫ�
��J��J��Gt�����4�U�|����g����X�޳.њj�oTv�H�u+3�s���T��ӣ�������:n#6W��Z�nL�t7�㑾��U~s�]��L��9��C߷����N~3�!�gng�U����*r�����'mu0*/|�<���2O-��QqO�������O���*��Ds�F.#}�uŌ'3b���O�b�kM�9���m�3�Wi�t	�~�R�:��p#�^�d�T��u��}�o�]"�J�Cu�F�u4��G%-�-��j���۷��zU; o�NW�4�=�ǖW�Ϣ^�Ϯ�˔IF��]�+��/!�+׽��*��-���7��w��V�G��}P�����ò^ZN�n�~�������z'��t	=�x	�G_�2�1T��9�X���q�'��q�����P��?��2L�^7�<�z�=zW�N����<�(�|�Ē�v��	�t�	��#��T�P��fV�����8�S��je᫬������䧳
B��L�)C���]�l��!{ӑ��	��is�}3 ��։v���r��q�:O<�T�v�6wQū8��R�����W_f�m:�b��f�W���=�]��dmc���ֶ)�g������|��y�S�n	�X-�*J��X������V���JC���r�MZ[~��:C}�R�o���~���_Φ���D���~+��n(�>�����w�G�cX'�b�YW��jY!�����"}�=:<M�z��_�$��L�2KF����F,pOu��R`�礿�M�Q���#P�~���@��׀�s�o��߁�s~��wce�g׭m�qET�W-mzt�6=�Z*�|�ѿ��5��x���c��d�{ޠ;���ފ������vML�C:�L��M�.E;B����ߢ�ׅ\f��q	^\<o�|cz+�A��u{5�L�����!� ߾�]���7|J��F·�T�N��s���f���s�f|�vc��^v���U.��{��/N�ό���~��-���|n�r�m��-_��^��^q�c&�{U�{�)y�=�J�2W�A�N��>FF�Ǔ��ݛr7!Γ�;9|����J���G�oM/,��S���##x���|��ȸU�^#W�yK�O_/m�{�]Ed\�(mGз8\�_�:q�x|�V[��T�t�(�@��*�3�]+�ڼ���](�,�co�$��A\+���X��:ZJ�ABTݻt#�� r��^N�zgcR�1�ȃ�����l�:	���2���:�[-�-�}��c��)����b�a�􊽉�JK:�\t�}Z��z�됉L��6[��ƶ�Ԧ�F�	;WvѠ�HN:�sQ�w%,p&�^汮��k.7�œ�G�9�n��n���M�t!p&�X�v[ ^wG�T���@�Nb�O��f�H�]��-b.�[�>GP���Ժ徽w��>P��X�Z#lq7�"Y��ס=r1�v��o{i��uJ�S\��f�S(�Hj�����#�Gfޔ��Kqn�Kn>����s���\;d��t��aQ��:Q!c�8�Wy2�`�@#Z�Z�j��I8��\t�[��g=�l���'�>�6Ӥ��fD�4+e: �n�f�@��f�70(ev!g�;�{�]v[Dju�T�aLv��IH�|nn>�A�q޺\9��(��tXt���ړ�v�&�v�vń��镜����c3fAK�f�H�P�9�&���������O��t��6a�fG�.��Y\3�]�H�����/ b=���Y}�xB�- 6���5�����jt�f�&&�}}�����pR�kv�,��lP�cy[�&��]ڻ+Y3�ܵ�$l�r� ��) b�b���*�{:,�9���ܭ�;MXܐ��)51��.qqށ\j�Чi�bkhgV�d	����m�A6v���I.�����7*�z1�x�g">[(��l�7��Y������ij����F�k�B�t���y�����yw���}J��z�'08A�uԋ�(�|!7a� }Z�tN'w��1����a� �k��»Y5��e��³kg*�n��*�y�R�3��� ׋N�<��sq�5��}b������l�C��LU�Gu-�n۾���"x`�*�qL�>�L���iAj���W2&��ޝ�h��^�X������=��Ŷ��Q-kߴX�$�nf����.�n5V�������\�V��˒�*��-���j��j"��ݱ�=�>n����`��w�O-��1�tvmu�)�+h���v:��#�M�x�I*dD�"���^�S˱X/�*�W��RgS��v]sZ�K��hO�^w"�R��;��J��հ<�zh��T�c���7�b�r�$�v)�Q���V󚦻�b��������D�}���}��1�����幦N�t�S�����R����/mX��.�ʋ�*U'�*T)m�`v3c0��4qB[i>�I$��;�Liw� ��Fc���C���y���=|�L}�Wm�2qy��mI�5�|�=��qsxC���@[���֣���by�'TGn��'p�@��uvv$wo�G
��	A��:/)�'���۳�ŕ��(���'�,/y�R��-���ꉋ#3�ݾ����S�1T�IEZMUkVڥ�5��
+Fh���mD�hŋ1�U;�Y�+Y���e��0E�j����6ƈ��������Yњ��(b�ѩ�J�������&j�"���"h��lLţT�;b��kZ#d���&	�IN�**)�m��5�
*��cc5k-EPDE%PD�0AQ4EֳDMkUQ�����*����DF�1�����5�LAm�l�cV�UkK����Z1LDh�E�Q�TQF�EDTle�mETL�[f��U6�QU1hpQZ44Q�E;fJ �RUDl�m15SQ-IISE$�U���AU@  �@��(��)�t�[���'��U��guD�핛������Y�eEM�);,��jL/0��vƍu���e��]��s���>�~U���
G�Ϡ+�
�N���}��ey\wdy�1�U~�=b����G��w�%[�O�A`��눩�)������Mx���7������?K�[��B����L�MWc����~�����6�W�H+��<��X��HL�'=�[������S�=�ͼ����r��/Pg��Q�o��vԳ2�.�3�H)�gb�P^HdRY�}
��Uz{3�()�X=�y��ޡ��=H6�~��vL��"uc�LAn��%aH�����e��*��\q{�'�5�g��y~�J�o�F߮트������ҵ3�^��;�7�u�!�7�>Fl�>�}�f@�|j1q�v߭��s��G�pC��@��U~5M��ꋑ�G�|v�}������l�y�T�:7~5��C���~�o��O�G�s��PѐM���[���Ɗ;��/��Gꖹ�rD{���������K���w��pڻ�4!)ؐ��<�y�j��'��P9Ø���d
�r����}	��koF}N}��e�3������8Η��ۺq��RZ����k� �X�]g�<I	�q{�V�����l�x�S^T��v�НZ.��8��f����GA�e�r.��b��� &c6�8�o���F�-�E�����:��O�e�>R�	|�iۃ]��_iS���J�w��y]м��zg�> �G�Ei��ѕ �t��_�}	�0�[�ʳ��d���$n7;;��_�
�|���q�ylg��{�>���=V���G�]HO���@8<�������8M����w�^�T���^���t��:�x9�����x�w��%o��w���v� L�y�c<�_1���9���t;���x�k&\
��w�SO��׫�V���%��ʟ��Ӱ�sބ��ϣ�9�,d-��I�3�]O�踧#�n ���p+��x���%��&gwk*��Q����e��j�!z�����r,�)Y�2�ē�z)�e\�[�VVI�dNd_z���Z��^uz �z=L{=�~+"�H{��F:!��׍I]��5U1u2�v*:���K�3�*1j����	���<�߿^�D����P��c�r"^RmK,"K�3
�Uȁ��j#ըM��E~7S<�}m���:w�+�yο���甑��~�;%�zo���N�I����m׀S�:�~���~+"��j��n��C9ⴧ�z��z��~��u�_���U�#�l� ����PlBqj�Wu!����JQ����%���7����܅�39��Uïm�o�F�ʾ�u,9�Vb���;��ջҷM�v��c�L�<9pI����H�e����ڤ����dA�]����h1C.]�}���<�J���ꚫ�t鴻}zj��<|��]D�!����|㋧�_K��c���-ƅ�E�O��z��|�>�;��J��Eĺ�ʒC]@�W�и�=����u�z�¶�=K5�����N/�.�X��:,� �wļ�ꌁ^���n�I��2CW���F赳K�Ϫ���9>�ާW�a�!s�mUP�m׉�G���:��P+�'�����Tz{�6蚺��*}��*�D�V}_���mG���W�jjK���q�_���fho�ʀ����jK�E;lo�1-�2v�E����>_�g���s�_ν�i��K�H���]1=����9�ܹfR�C����&�ǦW�:#��8VW��T�'Ni^+:��rg�c��R�[ۨ�I˅���RS�Bo�~��7�s��������@���(�S��],��,�	Uw�P+�r� ��$�����V��~�	gz���f�q�gI�f��������.���S5�]�~ܑ7Y��K�w+�E����Rg�O���������hY)w�aᨃ=P֟wʿI��[@�B�\T��8��j��'r�i�۩)T}w����v��U�(P�o����gs��Ki恏��,��hv�oWzq5+�%9Y[M�<��tˎ��$�������u;8��Y\���qC0��`�ނ�VuHI�zMU�?����
*����S�3z=���Uꎵ���̲��A����{�[�c�}Hxj�^����,��IG2�Bޯ#��T_���pN.y��2����P/��L<�ޯa��no���z�xqwH?u�����=��ۼ}uւw&��Id��%P�[���Rf���״��#���㸅/R��Q��K;�d9����g���c+"N�f��:3�L@R����I/�b��	�N��n�Ssƕ���ۙ��}�z\��>��z���z�ه��S�n	�����^SP����C۾͑W�%;��=�^��N�����J�o�'O��Q[�f��	��]F�y�#VI����S��3�ϝ��0ףd�������D� ztx�~�h>�dM˪���������ؙ����ǣP�F�G���tn(����{ǣ�H�;���������}�ցQ�߁�Y�Eߡ؂'�t����IT'4�?�K��w�_�gG���{n|���c��d�{ޠ;�Vr������t#�Яc��WM�*l��u����ԭ:.�ׅ^m>7�W���Y�Gu=��~��sMmM2͞I
Y��]Ό�lCZ���8�=雕���:�h�S�/gm�d�u �f�uBn��m,��S3�o�����Ka��Y�3Z�;�6��{���$�C���\q_R�����L]'�fq1��wA*Ѹ8y�©ǫ6toE����Һ��ۼ�iG�}� ��t6�<��7��d�WkC�����I�ͤ=�1)D���)���R�V����}�������"7�^3���/�͹ӑ|N��f<���Z�C3!���
�5��������o��w��sж�����ϝW�A�N��9�4;���m�H��Iݳ0���G��E��f����hmx��/E*�2%p�`
ZՑp�ԼFC���)ߡ�i��h_��]E_ν$���45�W ��Dϰ��t�����y���
��
��x���e��Y�y\wj�@�xg�����Tg/GKͿ`�>���jI*�|@���|�.�����׋���7����:z./Dϋ��=���m�褮g�ը�C�\i��$FxE�*P誟'9恅����q�R������=�=^�����Σ�ߌ?@�f�D�`�H�����Dߟ��O��;�ӊ�t}!*]x$y׽z3��2��CO^z�:m��q��mO�`����NTŬ���Izģ��zK����X�\Mæ�/k���W'=�#;�]��L�N�}�X�/���ɉEXō�Mb��\�q��)G�����=�]s4�j����ލ�K��}�V������JV��8]���W;�V�s�vS�����i�t&L�|�I3e��yݣp�`KL�n7&m���@ۼ��O�1�P�[>�\�o
�q��9z�b彞 mO�$#'ޮ�|}�&��|߭��s��Y�V�o޽M)@�pL#��H)e��s��Q�K�'��T���$�{ԅI|pf�/Ƣ1q�vڿI���'�� �u[�l��7�Wn߻��>H���ՠT5V��}&�S$5
hd���ZkKñ��!�=�)>�g�(�;�2�H��tc�.~�&ߧ�;��lW� R�rz(���0Z���S�i���q>�pn��z�b}�n�{��ruT=��=3q�O�=~y��ѕ �O�Q�h��4���e��=�����o��Å�^[�W���P��3�a�NG�4<��C��rU�W^�=M���7J�`zGl�z+)#t^��q~+��WᎪ���Bu�s��W���o�d͖�6�}5[Q{���|��d��N��n&^��G���M��Q���p*!o�Ǳ���!׫�Tމ6gj��{��'g�b=���{�|n7�5�2�ڎ��K���k�:-�ܮ��_�]�����O�/s6r���!3��,C�^+Ԫ7{�z����>�G,�)\c(�ē�e��N
��>��;1���)�hA8R�2��V-��P�u.� f�;��fI��r���m�����t���Z�8�o�KI���A�uk���/��l��,+k� үWIU�
�¥湂S]�1�Wq��ή��Y{l���F�v�8f��ѫ��QR�KH����I*��A�	\_b�L{�����R�.����^9eU|f<�A�LR�O��p�9�N��*��*���>�t<��o�|�����\?[�K�A�ö��%�}��Nۺ㼬\�'>��3��ϸ�L��r�ۉ�t��r�y�f�����6�����6~30Ǻhe��������99MI�'��P#Ų���j��n��p�����;���+��RMRȭ��U�,��������"�&@��
��x�Q���ȗ�l��y#��oسs�M��r�>�>��n����W���uE��RCW@��^SB��x�|��x�隸)�1��)��H�}�W����GşN��������lϤҙ!��=f*_W��El_�b�b�Fvt�G�׾��+#��UA�>%��|{ ;���w�ӓ� �|f)��b�e�w{
sU��Nu-9E#�q�M.�߆Bn�M�?P����q�346��m��P= {}+�j��l�c̞��q���\E*�2=��{��|n3�n|������.3�LOL]Z��#��_��__j�ה�K��$��n��U zu� =�=��'oW.�7�����7�QBwMS�>�X�p{��Ý��7z-�ﯦaҵ��ڇN�;�zqͺ����p�|x:����[O���#3��ă��W,�f�2���֩�9�W��3��=Gfn��`�G%���+�n��:o6W�u*��M{LV����ŉ�s���y5Q�E��ޏ޾������㳤�F·qS�tJ?�ͅ����7�=���c�YԺN����1�:�������XK;����n��:N����|��d֙��A�lxQ�T����qmx��H
���R߮�T����xw������r,�)��PӣEy1,.̝�V�K��J����<���]Q�/zk}�ǔ����/m~}t�W��ų9%G*��ԏ��Ϣ$�A��dQ�#q\;�a�ý^þ#���}p��"=n�;kѕ���l�`��L�����N�h�I]<����sS�L�[ub_:��ޑ�����'(G�[��{�"y�����=��+��}Y��ӢY�p@N��0�k�|�Ē�e)��~�Ⱥ��U˥��h�>����=q������v�<ڟ �{�[ +�i�����J�(^k��]��X�bW��ϝ0�;��k�.&����t߮�qW������ p��-(��/F@q��'/�Ĉ��9\
���{���\��������*�i�4`Ħ�֩,乩��M!#����%�^.�(��%�h�����Bήԑo|y���s���邔�u�#p5��q�;6��9�{5�D�>��X�Ys���Ɂ���$�O�#��a��d��<\�/�ӣ��?z���_�&�]W�OD�[�x�������F�)�>��MeC�i����{ҁ�� ;�h��1t��o}�^���=@��}32��ϥ�h��~;F��5�ۇ�U3��'r��뚽����g{xc���Cm*8E)��M��:<l{b���~	�^�ܚ�v�R��s���v	�{���]����^�g��=p�t6�<��7�Ĩ�h����N�s��E#�7^�rY2D��ԉK�����}�u���}�ӟo��g�}|,_��mΜ��������a���B蛝�蜆l��L�J���`�_��U��}X)|��yM���.=ٷ#qΓ��ٮ���&�}r�<����A�Q��Zd6J聵�|��!O�x�3ᯧ��H%�=FKq���{��j��@�n�о:��%3�<P���[9���;�L�q�-�f�ޣGչ��*�Gcݾ�󮒆Z�J��XPO�S>S�Ny�׋���~�=�]�b��%�C7V�Js���ʽ�~����-J�;��,���æ��V�E�E_F��s����C:�(�%����;|��A"���"����\m��x�Q聲\�a��B==3v�b�nf�0��ƎSu�SJ�¯���fY��5�ѭ]��S߇��/Jeg޷q�ϋ�F�J�L�֤��� y:*U!qU>Nq�`~�s��d;�g�ɮ������77�<zߝǻ��d@�f�D�_�$��-w�.����w�M7Cۇ�2ǻ-{4H��?^��3ϽCO_��@�~�TyDڟ�q;���*�ߓ�.�/c�����@Q��*����Q=����:���q7�Q~������;�� �?ߦ5#��?�����#���\���0L>8��>o���9��,��A�B6=�bw��O�������?C��5q=TO�©?���s�HU�R��܀_�b�P�W�7cB��6@��qw�~r�r��='���"\9�=����S$5pX,��	�XiF��G�9L(�a1P�Tt�Nnx���	�Q����;��2<��+�'��>���W��ހ����K)葞��\ں��-�:һ��7���=3~���w�c�X�./����^�#���ß����U�F+�J������Ϸ�Æu]0�ϴ��ޡ�W��zsޚw�!��	�5���4�zk�H��+s�4R�|oo*/������
��.Fu����AX8���C��R�ϱ藦g\޿�e�S��s	�M>�z�����g��.�OhV��6h%���$��[��d%Y���h�C��ѹ�I�e��D��s��L*��.e,!�7����\����ǎ�-�I�H���B����t��\ x�����7�v�zѴ�Y��96:��#�N٘��8�b��T���:�x��)�l����Q��aۡ�.��l�ټ�l��}�о���w�gTs��R��\5��$���kG�<Ř����c�j�4�&��(~x�h�z�V�'\�s�s�EEA�Zw�^��
n#:�-4͹�R��QţlU��MZNq�p'^�WL�ذc�f�U�-��|�w�V�+q�#��e;�֡F�������is���z���y-t2֢(�!��7n�۽zn��y�i�q�q�r�&gv��9C���]we^M�V֒�7i7�䚊V�� Ux�-���jmb�f4�LUtv�@�EJ�L%F��&"97�zi�i��^�%˥����Z쎋K�e�
$ɀ�D� �9�$�6G�Jcژ��Vk�6����׎�N��ʖ�F�k��������(���8H�ü��}�bI�"�"���˔�YY
�4�w��{ge�skY���WS��17p�V�����X�.@y�Y���eru^�s��\���*N��j�k�e�<J��ޢ]�a��['K��f�Vp/�G�1�(�ڇk�=��K㬝8�.R��z$�'HCϹ�!a���|@�A�f�So��,�KrsqZ�,�nsys�c�%϶����eXF��:»\�������M���N"��n�g����-c}�<����ۼ��Y��08/ZwT��k�	�rN㛙����<���dK�j\�����4�6Z^�0�	Iإ8�=��r�S���i��h۹n�+�
f�L
�s��<x�������ؘ��M�#K`�Zuw\�j���Sq���a��6s�$b��^P87���ק`��i�6��ų;+�5��8jq�7ŷb��<��^�`��jF�f�0o�"�z���qQ���J-�h�7�!yVZ�S[o�Qv�7��-�&����Ol�W���mr+�l�\6��6�}r�s���m�H�6x��ЧF[�2�����B�����FfZ���[D7��� 9�@�����}�մ]Z�Љ.`k��u:�/(j�� ���L�|��	�����A2=���0���C�����6� ���K�Rj�`�:�Th,a���w
ǝ.5c`N��9�N>�D@�����s�������IJS�tx��'ne�c�e!1��l�39���t��rô�����(��C@MR�tr�w�_%z���6�����n�c���o�w��EG{EAQ͜�ƒ��*����kET�14�cm����*�KURm��l�%QS��6ŰDU)UD�J�EkE;h���� ��
���������kU�52P[)�5HDkQē���KmmX��(����h�Z��D�IQ4�UM%TEIU�1��-��L�T1DU��ADPZ��d�$�"KmLK1TADTPDEDƱ�l�i��j��Z*��������
(*��������j��
h��B����M ET�ĔU:B�t�F��-	��
 �{=�tfS��jNó LGH���{���]��oKr ��Yo���e��;]Rv9sFҗH��+;ٜ̈���r��~d��xf���Q��e$n(�'M���q�j���	�����*~o�S�S�{�c?�o�r��}&���1��el�ΝN��`�t;�ʮ7Ex�n6e�[�Q���zs����f�Le{��:n�S5s�e���	bw�n���ja8sR��������~C�l�U�үk���:[�(U����^���;��=j�=��c|��g	H/�,]L�Vg��`��u����k:�u���M�7� V(�1�������!�q���^9eUD�#�~c������w��q��X�L�n*��y������^�3�����qȗ����R��﯑[lx�엶���^3 y�vQ���S(/���o�N��!zG��o�q��*#L�͑U�[�'o���k����{B���>�R ^���L@n�G�et\�|n��*�Ӵ�As�+�ر����NmiY;���E{}�#m][5q�P>7�u t70/�_���_F.����Is]3�J�.��W�a�m�g�}=����������U$5@�:b^SBY��=�r�k�r8nM��/*m�Z��orx�P��@���T/��n��RU��G�'ɥ��۔�m:#�UrP>|̋n�/�i?�Gc���Uy��cd��}�ت�sV�����u>����/{`�@�(����.u�,�����;V�ÿS�MW���g�x�hz� W����n�I��L���'��o�7��|5�W��k��UE��\l�z�+#��m]и��x�g���q�W�.�*�'��7n|�i������X���_~M����v�j�����ϓurq�@���z�0de[�`����E�B�!�6N���|vp;�V鿨�>�wK�q�{p�!?]�}��M�$v��$�"�d����y	�}��ܛ�����}r|��Ⲽ6�^���͕�J��VGG�G��n�'��*�/]��$◎�g�{���>��s�t���;;q3�*�:�NQ�t��:k�oպ,ƙ�}Pg��y��`{���ez�/�ׯ�VǽV�V���m���'v�3+�>E���=ޚT�d�_���Jsz�s�Ϣ����P�ց���̦u;������H��p��e<k��P{M"��e9ʞ瞌��.�.)�#R��T<k�;�N��5��c�"�hxvD��+f�GS����Q�\8�-;nC��,�$�hʨ���7E�L�|�����^Ñ���������{�ϥZ�$ʮ�.�:X?n�f?��5��Dv^�nP���)��-Z�)�O�ɪ(�I��z�v��`Ӷ����Ŝ_��b��50��<U֕�B�n>�1�����'|��85ϩ��$�����<�)�a��Ś��]�U-�dƔ�
�If��Y���N��,;'��J��G�C�[�ڟRf���״��^�~C��zr�����T����������W��������	��XR��|���L���Ba�A���/ם���=�|��C{�|\w�i��=냷�fmO�� &pdvjr��U~@9��s���H�^t��^��;c=;��l?R�o����TS�2ʄD�8ʘ�pO�P{=�
n���Tn����ZېÈo���O���&�~�h>�dO��>�z�ȡּs�.֏��}�$�7���_S�!��ɇ�#P�~�~���	�|�,eί=��}U�y�I����Y��W�S��/�l���z=�v4�5��y	��;~��K&�L���z=�Ϊ��2}��P��~Tp�Saʛ�r�\NIZpm=�
��i��7!]H��5~�6��]�m����5����7�� ��H�)6f����U&����O��>��/wk����C����s��L;��bu���ޠ�9������G��s�����ǖW�����i�jF~��W�r��CIG/+Y�3ygYF��F�8� T��8�(v~ߏ�U{ޞ{J�x�z�m.���/$��	Q���gܻ>��#&�t6��`�Eۻ�Hosz9��Ww����fl\e���粊��ۭە�Y�Wm��m�R�]����N�/2���#��>7Nt��[ U��c���)ϻ����q�׵�~�ۑ����M1��SGP���z���1�G�a�eV��+�� W�Z�/�^��1�xw�������HB�B�d�U��BͶǽ�]E�����9z�_��d8G��������t�}^���B�����|�;Й~�j�{m����IC"ԒQ,,�L�rO�Ĳ��k��%��c30����j�i�>�P����ޗ���=�ͣϥq�r-IT�$"ĕ(S���۩ɸ��w�%E�Ԉr����4������1�����\?;�v|]g�z;&Yc�,G�z���������������n�x/d[y�Eç�ѐ���V�ޡ��=H6�~��@��Os�X��B�f��{�~*�f: ~�.K�U�a�^�rՠ���#�ӣIQ�QYw�v���F������{����L��D" �G��p6��τ��Q��C��m�������b�~����#2��Ў��>��L׍2K
Ijn	 �?RT�:7"~8��:~G
�V~��S�ޮ�嫿s >��_n�A#�(���j�|/'{��{�zE:�e֏9���I��n^�:��D�oڰ[[�>.�������u{;��ź{'v�R�rM�ȑ��� b�n�e��jd�����b�!.�]k�6�#���r�]Փ����?_~'��<O�́��_����!����K��>+P�2E��.\ؘ���z�_y3�\�ڪ��Q��~�@�dQ�_yQ�B�rz��>����=�]u�:=oZQ&}����j�|6�]��ϒ���1���������<��ދ�z|J1�oԽZX��fs3�-��'`��Ez�M���wu1����'U�8��<j�=V��?M\�z���f3"}�ѳ��U됽��v�Dn�9��E�:mt�ε~��Js��7��A��V^�9��)�;�S�	�}���'��w�:t;#�謪�qEx�n6e��[�q�"\�^�x9�7�Tik\@�]��nϗ����Ӛ���;%�%_�~gE�?!��a����ˬU1~�}R&���5����p*����ޮ����z�\o�]#�g	J�� �a�n׈X�&�F�.�}�VEzG�4<���
��=���VDW�ps��|����,�J�6V����'٥9�_�l���gY��A<yty������{���L{J����>����>}�d҈���HF�3Q�յ8�aں]6�"����܂[����a�4u=��EsCq䁄s��6�� ��دR�)�L,]u�w��b��2��.�:��}�-�@�:n��ͳ��;����o�VD����k�I�o2�������ϟ'_���Fc�O�*�qF[7�L��r�ۉ��;���zG��}��=�2�?,�vEx��������;��g��{��X:vK�� �O!��_Kee�����*�;Hϭǘbo�7~����T-�篊G��4����F߮���z�pB,�:�7P(����� ߠ�S�]{7(Uw��_�c���,�{I~�AΊ�ߌ��M�D�t���;�&��*�'�����1G���~�
���!�6���*>.�|K������m���I�MU�e�b�+<=�0��B�_#��UE-�����.VC����-�����4
�x]�Qo�U�9{U�`�/s��L��Fi�
��>�����zk����Ȅ�\����G�~�����MZ;�e��]���ьm���[ �����w^��t^�q�/Jν�x�����7�ʱMy�I͹�<ϵ���޶'�#i=����cgC��+�d�'����z��o�{]r�vq���oz����2��s}U�+?~���NxΜ���go�Ðvǲ�^��O�gɲ�vX%z�e�{��8�6��x�/uӋ_S�J��/*`؅$�/�F��K��f�Ak����v[	[�{��\?�9Ƶ�7կ��F��Qo9�^�.u���nr�eZ�����̎z]�X\��u��;3m��ednl}��6:�v%ǵ%�'<��{��|ꗲ:���؏z�%�޾F/}�u�!�'v�33���?]�٭����pj�J}l��S\n�@j��k��^~��3��;�����>�Go�/�`G�؜�_Fr����a�}���rQ�#�w�5���zi��<�����Ӟ�1�ɇ��ǳ�:�+�{{����Q��ѯ���Q�#q\;�a��W���G���y�S��@�x�8�)��6�O��>�A�çd����Op<��L�1u>��}mՉBn6f6o��}��,�ߟ}�G����G�\g�����d@��,ۂux	�)@�>nbL{��O��w��Qw����Mt�"�V��^�4'����w�i���������S�8 &.�P��:3D�ծ�~J���t��Չ�O�0�;��o�Ը��o�'MǮ�qNL�'ֽ�]�U��,z��2�y�6�$& ���n����V.�[~v�z}H�d@���7ޭŜ�^u.�)M��_�^oR���n�1}�P�8�C�q��m����H@���*�Ps�+�!�y��37�sx���5��VbI��Ό���bX�Mp#k���?j��Dco:���eѫ(f��nKŬwm���b�s/����{���ko��T8���=���>�W\��#�7{�ju[��.�9�'vs�DV񔵩�q1�+0!��ڸbG� ��xցP�[���f)L�)������qR�v������T7�B��~Q/���*̫^�>���%���T6�ʎJl9Sf厱����ӡ{W���D��UE��]rM�[ϙ�5yp�?]�~����� ���t6���7|J��X�����y%�Q�to�ε4pz�|N��Q�x�N���Azs}5�=��=�ʜ/���瞏{X���I����焭1��VWq�s�����|��!�z��N��9yM%;�����8��������#��/}��wl�<5*�]eV����*6XakVE¯R��;�k�!�)3<=Ҭ�������k�!��v��{�]Ed\�(i.�D�u����y���
5���H=����}rVF.���_y��]G2�^W�{l/s���E�$�XX&x;��)��r��5lv^`|x�W�6�}L�U�o]i�~��N�ھ.��Ҹ�9jH*��ȱ�wx��=��(�����P�`�T��r-MM�>�xh�!�cs����q�ϋ��dږXD�'�;T*�Ƥ��gI�>��vs�����,��y{U�]i�z�E��_��.�mg��B��EV}�ciĚ�Q�s홃��U�Y���yEvz���+��*J.[u���r�t٧�λ�'pS�h�]��R�뻑���-�ާ�w���؜WC�aU�:�+ڝ���ďA����L��M�	���d/uy���z�=H/��;��+�z�/�o�f��}�+���̈	���<�=+�T|{��m�X�A{^G����)�x7�'�{ֻ��ψ�G��
�US�d�5�3�n��_f@�|j#�7�l��\MF����ʛOj���e����Z�߯@��U~5r�b�U%��$�ԅ\T�:7>����*c*cށK������y+���z|��7�|������H�s�5�Hj�����~;��+�ﲼz.7��o�Ƭ�}ޢ=pڻ����7�?O�w�:���*6@�r��Q���� ����ĮW'�_��~���J]+M\}���j���%��!̨�z|��ȭ7�ʐUoQ��lp��XS��Ū���随�P��vU.M�G�?�ɞ\g^��W���q�禽W�M}O����w{���g�۹#3��� �h��v��VW�����+�񽮯��L�L���ڇY�5sԳW���)�{�����5����N���`���M��l{*��|�~'�'�%U/6<�7ٛ�u��M��z^��R�-Ьg�	��5sr�ZFӰ~��>�
\}S�:����i��7�S�xI[k���>�
��{Fn�%]=緃�]��^[��7N��;��pُ�m�ɫzlb��5w7~�!qE�ث��md�\�O�S�Vfk�����:�w��{nȅ��w��C�:t�/�qS�:=��yl��6���*�Y^g�% �}P7�N׏�؏]?��qݑ�^�����9p���,dl�HW[gޞ��9�J'PxΏTϙ����l�����
�ǯ±���ȯR������^9zv�v�9�1�����}D���DO��#uR�y.�{׃#}��H��Ǹ���<n]{m��V�g*���,��>6 �L7FX��(/������N��!zG�����R���9�`.>��6���=�:vKd ����=-��\�|U{�+{״Ƀ^�[��w^�~�>��|u�z��z���ճ^��><��Y u���҅M��OD��Y������=UOo��щW�lÏNu�G��=�냷��YRHk���o�N8��B�[�g���&���_�|F.��W��G��ώ|};�^|=Q�*#޿\M�3�1��s���z�TU���	�P[f�)��g�S�U�Se��빴;�y���ny_��>��DE� ����DE� ���DW�D_�DE� �����"+��DW������_�DE|DEp�"+�DE�A�QDW��_�DE�A�!DW��"+���e5��D#p=�!�?���}�����nUPP)UP*%T��P�BAIHEIP���RB���J���(�Q@�T�B%T�U
��
  � 6JQI*�"�@�P��E*�
�*%T�J!(�H
�$��A��
kM�U	��h���&Ƣѥ@lXdl`S��(RB���')'`�@1 �   �  ��  q� 7Z��!5�B�T��J�H���J�B9�TP�fJ��[`BلH�@�L���R���T�U�j6�
l[�i"��X�d�����
)�k)Ji
)D�n�@V!����iLCI+m��Z�$�h�HҔm�h�LkiF����QB�W w��6�4��R�Y�[j��mBR1��5��U���Պ -2���*�ّ*� 3����CA�6����JIXM(6�SIV��P��@��R�(UPp njaZ0�"�j֫3Pф�l`R"��Mjm*�P�P������[�k	$�di��f�آ���6�	��U*���I,��(!��U��i�*�"��DU��$ (   h�Q*z��@�h��
R�R 2h��M �I & &�bF��z��hf�$��R�M 4      sLL�4a0LM0	�C`F&�A��RF &L 4�`�	���u+��<���<���zէ^Xg�b��i�DH�Vg��Ȳ���%�`� �"���O��Kȉ 1H�5��:~2��g���⍅$T�*$n�D�h���5�$�@m���A�QPaRH�:GN\m�F?^�Gk��$H9$՚����N��9Ѯ�KΛ3��Ξ�Q�����������0�����<	�}����	������̙��Tҍ���<��#"!T.%eԘL5t uy�*�������R���zQ�A���-� �J̧H��r�Tg)�ݼ��t�L%Z����1�ܭV=w�*��r��d�{6�8vj��يeR_a 楙g�)�N�������a��{Հ�Ɩ��b�	N���*��R�U������ӘEӺU�����8%�Y�Bw�{B��2˙�b���Z7A�[��b�	]�t�^�M�j[��8e��7�E|F)�j��m-b��EZ.�D�D��6m������dgr�<Q\V�#ʹϭG�.�x�m�������iۭtN��w��V闰A��3t�:u�u�M�� �i4S���H��U�'w�*���K0�jK�b�X2��+4P�r���퐷j�&��p�f]��P�Q��S�vܭ,�bH��W�w�?�����{m:�������Hiⰻ����wW{�Y�Gi�����W�f&P��֢��ֺp�v��+iԫ�Fcƅ�{�rY�d�vnY�V��`���%SVV���.���`�q�FR�[n�q�+ю%�[WTh�a���ܩ�nݔ��F�8�٠��)I���DnQ[q(�ȵ`����4���X�Ly54eC����P�6��x��X1�K	�դwY3�:o0W��*��ɚ�;�;�kq�!��Vf���j� St�+9o��j:����}�W|��z�v(�$7���Bش�{W%bjŐ��l�j�I!�o���u��r爋�E$�U�+ZN��}YXm�+���϶�hd@�U�X�.�M*�kFf}���F��4�<+u���+�d��}N���MB����l�k�lm^�л.�`�L����I��ռ2�mQ��'{A���8�]zb��ֳ��X�8+1t/q���e.ބ�vR6ۏv��͙�ʤ�s7i�ƫ�#U<U$�{Y���&�ǋ^��b�r#T3
vk	`�3n�T7yZ�$M���̘��:	a�j(49U�PF�q�V��QM̷6`y��q��P�*�4fcݬ��ҍ0a{�(Vi���Z%ZrٍXV:;�� $���PG��Q�A;�\�0�Kj6h��h+��UnGG[���Y�b��� Uޮ�v���tQE����Ϗ^��d�)�@�c{hn&{����v� �̈m�siV�E��l�h�,:γJ���*��M�x��{j�V[=�Y�\ˡj��e�O0�e�/dc2�4��p�r��%<��Z�=xb�*A�[x�[o�]�ú�Y�*]��	k�����&G��o%���cA��VM�nŬ��ݶ.��DHX�[�Z��˳@�/&�UIV%#[�����VN8�j�Eb��n�i���NY��YB��hU4�CLr��f��}���oA�b��V��+��Ü�VG�ڍ�M<���uk�
����3T�[��Ϋ9+A�m*dZ(MAQ"�.Μ���Dn�<0�� 7�,�d���ʮ���r����t�,���f�љ��cP4�l�/�ٲ�$��7�V�/*��o��|U��U�l*Y;1b�Z�Y���5gB���w �u��^�k.���\l��݁J�c�����j�;��Sa�w�;$ů�]۳�9mxl颱E���h[�ޣhգ�ie�Fݪ�B�B�*!�*fb�v�0TobB��[5�FP�9������m�vF8��Y*������V,#0U射��ߍ�s6+4��inE4��'�&'H�I�]3/lЕ��D(������-O�ñ�,��gy�׸�(iCj[�h`��ݝE�d��w��22D&���Ze���#�.bcJ��CIh:�����?c�M��д�mq���O2�-� pe��}�Y^�������|<���y��v�.�T������TЖ�2�a�{F���B�Ya���9J�;��,gP�F�����������Zz�u��x��6������$��G���@˷qfhz(��qμ�������ר���X�)Q�LO��VL�w�ax�X�I� u� `���&�*�5����*�XRڀ�R�$�4�m^VԢ%Pw-n=�s��l�P���ZP�!A7X��RC�T�V#�Elhb[�ĥ^�R;۽�ݚ2Û�L��"�kTm4�Y1�Z��U���h��p�TM��[{�Yu�#�X���[�u��]��O^�=�EY`QCK���u��Z�`�'�ܙC)��#��5�"A���w��.��
���*�V�:���V�+kҮZY,�Fn��-��ۢ/1��U�"��,3����i�MJ��Z�����̙R�udt�7T�`'*he��v��&�]���z/o�4�KC�w.���b�qD�޷���k f�)�)Vi��d���0ob��O&C
ӧJ4M���ۆ�uP�e� k��F��`�p��3":����;�����X��"d��lWT+K2�8Wy�]E�hJ��7�i+n�A)1ѣ��9�7���J�krڠ�kO��R��*ڣ���|���ib�LJj�"�[h�:�^�+"���Ӥ���ۻ�h��y�R��q����#���c���h���	Ϲj
�U�l��xr��m!�$�kiH���g{-
 �}�.٥]�-b��@��z�o|��v8�7��^������؋
�4ؖ&�@�ݑ@�F�Yh�[�3tP�*�6+�j*1)x*E����P��Zn�lm+OV`�f���Q[���ܻͧ�N̊eVS�iw.n�?�ނ픺��T7ps)�lU��Lm�e9̗���"��ݽe� �[9W����7v0q�6+5c��QJ7�հ�^+�˚���&��l!����r��R���r����Jma���ҙn�Yoz2���{V�LuJUf��vSɣo�D��5fo���*i�E�޾b��]�H��h�mR��U����7n�����i=���Bsl"�Z�sq�LO�U��[� ������:���MU�}������W��⥗���3*kR����
t��0�%�*�3e��]&E�:h2�+.1R+�k&�z�R�2���U�	��������me;f�.5ˁżQ�/k���ז�3�F֮�F���٭�RJ��U���+O3}dg�.����gC3�2�-ͬ[����jL��S4��v-�;�y�D��re^�5�y>Wo)���fI�*�ؾ��I_!�Sh���X�v
��W���Xm�ȬUˢ{W�ؙ��i��x����a�aM'���]���Ɋ?eX��<��b�NڤS�u��DfH^��1!@����OGu�gۏ��c8�$e��`
JČH5۵w�2MT-^�S��S�����)��#2�X����D�һ0��[����Z�/+yq-u۲��b��׵d�MRr;32�:��9�7Mp���օ�x�VB�0�tP#&G�ջB��*ƕ�%u�dZvR��=��]��(1i�Ɵ��W]�9[��5��W����tf.c�h��N��K�`6�;I�%��I\������m\��,H��0<!��.���1Q@�F��F]XW��5�I��Y��$�e0��*`R�l�1���[�Q���ra�Z�gU�M����
����m�i�qc)���.4	?3R�(MJ�hJ^��o(���z�+Q�T�	�#(=��������S�u�9sYL6W]���8��y�F�����uJ�����G��:�A�����e)EWY�T����&�=�"�Xx�A(�-|k����ҙ��p��Ÿ \j��v9�*-<�W0�n�0Nr���j@:�_�+���*i&j�b�D�Ak7S��!�fE�w�G6(\�wz���9]G�e�JK�.��}�%�������S#<&��{�
!vN��wg��ao�>!\o}.�7�;E�'�d��F ��u��#uzOAYf<��gi �=�E�uP��9�׍]bS+�=�1���[��8VsSw�x�=�{�v�c���
�K:�[��]��q��J�f����AB̨��Ӆ�Y���.4�y�E��s�"M�"�eh�����t�R|�e<F�SSz:�u[�E׌�Z
�L=@�[���qH�q��`���a9J�� �v�L���:m�WP�.:����R7\��,T���r/�'����yb׎�R�Sr��tX��*�V�5�bY�����R�k;6Ԥ+VB��ݺ[LԹ��`cIsE�{h�J�;w�b��6�7Ɩ\E�
gG-�4���M������_wi��W#�S��ù}*��u�͚`Cy���>�f�ŵn��JED}�Yzjkz�%��?l��x�ټGt�!�p*7���c�N¦��`���1o6��\������FL�K��j�>��n_k���[�AG�:�mj��5��R�	1�5n���]��7lJ���W/�|������ԭ굕%8���蘺V	@p͹wV� ��u�����76-����@ՍS��6���2a�:��u4�Uީy.0�@m����{���2C ��.�u���E��E{\�]�|��s�1J��`�@#[���͘�_P�wof�
�MG/��i�.�V�G�/zcl�u�)�mA-, �N�6��wX����7���&�Mi���Z|*p�X�Z*��<9��KC3hn6^$��gu]�F�J^�
��Gq�Q�.�����"�R��ݎ�@䫷G]fnL-�y�B��u��[C��X�d�m��V�1�0��,�uę��R��`�
�ٻ.0�2�P� ���݆�f(l��Yh�c�3���{E^u�۬�Gn��pm�Woz_BA���֐r�5�3E����T��˥t���yz�,��0���*��+YV)U�@�[�-��iG%��x(�;Ў�]��;q���ʸsn�wB q��\�(���2��:�\��Y��� ��.OS�rl���
��J$;���s�(� V՚�9]�"����(f]��E꒘���`ӝo9�rNmw\�Ǥ%u�%�L�.����؁X�J.��ͬ�Gd ����wq0�Q`�o�l��u�vVP�/�؀�E��\s&b��YK��޾����"n^�3r�Fֹ����]6=�ó "������l`�l嗧v���ˮ%�d�yC�"�k�ç�0��j��o�8�[AVR֌6�b5�+(Q��_D�U��9v0���od��Q}b�h���
�/on�2黗o_�v��)�f����`ղ�r�p�\��3�P��h�*��f��s�����+DOV��3��Qu��:�`!f���V�;mSY�-dOn_M�ә�8pf4O$�kS�F7M��Gdr��".�2;ioXW,�.Vs�)��3Vw
;B^�]�P)�/*4�&�#ݎ�J����V��7_&���݉�(��ս��(em�P��녗c��컺9o++���Ԝ�ߺ�*kE;��;��!Y�w7��U�#R��k}���� ��Ȩ�\�%�ZUU�2��2fև"�2��Ǹ�ؒj�Wb�Owt���#�NI��w���q�����5\���D$
V�0�A�}��+B<ݠ��է4C&���îm��K�e��:�ٙtJ2v�ɝ�h0􉡏�Z��;������p �8Ȕ+h��:!���4�v\��Ʒ.�9]ۙ��$�EV��S�M[ju@]4N[%����Í�t��P�=�vPxy3��tD�j�i����Z�;,=�)�N��7H�Om�,^��,����\:���.�s^L�r0ip ,�;Wx��rN�s�=kJV�vY�U��|�;����H�Z̦Uu8��O����dT7�JdJ�4�$AҸ�<
#f�
5u�&���.�A}�v9|ͨ]��TW-�@����黱q`AcS`�}}3��z.�g��2�!z� ��|p9z�����û5Z���J� \�۲���,��4ox�!�e��B�5�����o�8��y�r&IX�U�_vǙ"��"��hâqj֌9K1�{וiĮ�<�كf�J4f�IӅ��n�9X��)�9E�΋�Ck���Ԯ�M)R���6�YB��n�7�.�����7p;�4���l�2�e
����杹;+�����x�A�;I��'`�ܑ��,�m��a�|�	�\�1cku-��o���eB�:�#�ڸ��;`&�+�a-�2���nk���}ӬCtb��w���RCQ��8__uUq����z�J���pa\s�i���@�˻wB��R�9I��K���o�K�u�G��aj�^U�i�9���]� ����J��JZڷ*�^P�3�R5��u\˧6.��7ب��e���|��\�/#쳝LkJ�ft��$���3��h�{�O[���������WR�������}x��ط�Fl)e$,*�<��Í������ ��eof�F	([�k|���R}���K%�V<ĩ,(d}d�wi�So�w1֥iP�aF����vlQ�/����9DKBk4cW}W�f����Tق���`*ݽ֐��Lq��i]x��l4���
��޽z�6��n�˔x8rm9�W�d�{d��Yf-���hG(ї�X�#tŅPV�����!���52I+���+�;���f�T�ZD!�-;U�ڔ�Dv��)"ŗ�f�c�r$�ڻ8\h�Z���FWQ�K�T���ފ?A��{�S嵃vf\�p��޽�ꊹD3bB����+���zo��6.X��k��,����HE�8sgMfG��l���@��p��i�
3o��1��19ٓ,1�@=�f��Vkd��2�3&<u5V�`0Έ���y�ow$"y�j����R��7U��kB�"��C��;\���`}%&G,mnax��kz���1E
���@��-	�:�<�Z��e�i�x����y�)k&-�ve�X�U�g�gL��`h���AEV���v9l���h���THA��1̩���1pӻ|,���ڕ֐��t�Y2:�-h��ݸ�G|w�<���DW�%2V�y��Űd9,�V:5lt��ok��ilⷆ��+��{4JJ�zK�c�8���QJ�(͎$�9$�I$�I$�I$�I/2t��u�q˺rF��^c�1QL�]=��\�$nS�LNK(����l��ܬμ��Y�'rz�|�[WiYsMl�6�:嬾;V��]����D|�Wj[��l�\�Qa��!����و�5��o�(��6$vh�s0Q�PV��֘V�%}��!i�hNu�.�]Ϭg��R�����yF����jB⛛,��ы7�_Nl9�6����r9O���XԱd<�2�'[���8`�{k֪��5�Ȕnp�����*9��\������_s�ر�,kx8)gZ=r�Ś�F�*=��W�VAaY�lJ�|	���@�&�;ў�1��+�5�r�-�N=S�WP`�8�:&	�,c�w���������g���n׵���Է���"��}1I$���t�:ѯVʪ�O`�H�������w�7������Jq*��t���H��,_V��%u�SA�����]T�n2q{7(.SK�sfT�7�dN}�j���s�~�h���g."�������2t�y��BKLa�:���Й�C*��
ɖ9��!�Ek����^��b�n7յ{[��`Q� ���#(|���1"/�����pN��ɓz��i�v5b�eJ��U�sא��.nu=�]�a�R��i$�jo�F�)Z����D�Q�Uu��pU�#����58���f���r��U����{w�$NF���^�a�������r<�^#�x�\ڹg���isb�/s����R��i����$�ں���P响p�|��8�ֽuu#��:=/zK�*9Oӳæ*�j�:e�8���m,���tH�)��^��˭h�G��w�o�n���^��1C�>M��g��NS8n���.�[��ng3B�g�+Ŕ�D��#��.�wTw+.��1�F�DC�� �J��v�1&w^J��P���[{H(ծޥ�e��8�h j�V�q��VM�4D���2>ړ�wS��k�#�f�`�F�����T1���0K�㯧���_�h���g�����!�aJ�.��m�����L���o��훦�C;���a!Y�IS�|f�H�0v.´��;,��{¤��2��2)�)�Xa�EÛ�H��lv�t��R��g��ة�j�Q��N�2��hDblͱj��ylr�Q��MQ�&U�p�@�;	����8�n�T����yw�&�����cBiRѤS0���{��V�n8�lGK4<�r�\���RCi�lYա\�T����uw�$�73H�Z�4���,m�|�k��*���nb8��l�/�}ʵ��W���=�'�1�"�45��a����O.�R��M����BX;�Q�7�星U�K��A��s
Z�qs����C��>ꐋᏜZ�3G��8TЏ�ݾ���E�ʬ��k�^��v�:�i-\�-���iZcsqor�v��ݸ�^�&N��|��e���3��c������w-YI����n�N�7z2`/����x��|(R#U�>���E�3�Uц���e��D���6m�S,��-X�zx��i��ޑ��Y܊ڣ#TA�4h�I.b�2�(���Zɢ��]�*X�9ˮ|�PYQ�eU�Z&���]��Wm�a���
��
�`�n��9|�j�����Wr��]1�D&ee�@�a\�#�̊)��y
���GtC��as����]�"��K���q	C��&!x����{7���
��}dO��J�Qg�l��&�u�쮼vU��$�Ҝ�U���p=]��SsE��ʮ�SsA��RnQ��Of�]��=�,U�Ԝ����M9���M�u�u������		1ަlJ��F�Y.� wKW�IO����x��{�T���5�Z��vUf�C�]b�	ڱ�bm���@gK�u�[w|9r��y���\e`s���:f�ͳ�j�Z3K��ە��\b��_�&9W`�j��u��7Θ�'�a޻�i�,o3��#��\MH|_u��7r�p�p8x
Y��1���_=`��Dd��"��0��U�8�B#�Jet��c����b���p\��Q�]�C^+Ɋ�Q0���)�YK�v��y��Ggh�#+]q��t�}҅<8�#L�btzl:��d5��8,�l�R�N3���T��3�aj�.Dw�E�����r�0�*5�uN�_9I7!֥v�%a�+�٦�-��v5����@��/M����oL]Q���7��7�[\��	�@����/�u���\_${/+�AV��U�� �4�ǹ9&�-��/GVEX��s(�����WA�,�k(P�B	��rԿ��#�[f�J�6@R�o 8�{(qެ��
�w%i��U2j1U��=��5�>;4�W���9��]��4��W�;]F��ڼH7�J캋���qu�0NG-�@�=h��Xq�z	�;n�	��Ly��n�a�0��RVQ.���O�[�(U]�-h��
M������l�7�g6��[�e=�ݨ75��el�Q-*��,����a��Z�#��[J���jQ�+�,�^s6�"�j!X��p�Y5��.��:�';�y_@��\�N��Wv�$ˏY/�C��nt��H���ܛ���B���ax.�z;$^<>�w�^u�H-I��b�W{a��#t�*[J����$vf�o�U��2�v�c �Y�q.�Tf�s�<]��v���>\(>ޖ/,�R���۪�u/�]Ӏ�[Na�Ԋ��:����#b���+��J����B���|]e��\`�2������6#pE�k�ͪ�Ղ6]]P���7�7{�6xK�v���9|�1�4��+�w*� Uk"�{�6�r����i>2u�[��3oaM2�VAd�|0�_���d9B��0�hn8e�s*ެ�h���nf\s��3�d��R��sv��]��k�,�mte}ԁ����[�)�K<�f�N���pP�;��!mn��,�ؗc���><�h&T���*�[��E���u K�ZΩZ���<��U/U̻{c�5֓���E�=��rv�æl�����Ȯ�Ҙ.���լ�RE�����0��,����vw=���{[M�o�YOgf�st���"�lX+%��Y�7�k���>s8X�ά��06�84Pͼ�Muol�[M�gJ��E�1�"�2_b��:L�R���[V.'")c��CE0��ed%u&W-N�}��t��p��#70���g�T�[VkaA�r���Ԡ*����x�ה�.�)�I�Q4�l�Kz!�\-�Cch����9�_e�֜\��>�Olk�l���i+�:t��|j��Y|Kjdk{4����P#v,�G��6���0g�u�^;�\wH��v�X�g7\��a �%��@oo]���������f����W�S�/��XjZ��ncK��F*]H�]pי���u:��)̾匚x
�Ŗ�@3k7-��l\R{��+� k0��^���a��6��1T����w�o(�FjG��;˳g(Y�tWX�.Ch�}����2��n��>��t�J���ʐ\�\�ߵܣ�fmgE>V�[�"�4%R�8��]�Ya�{��@^q����U��)��W���^�6v�1ls�7�1���? V�*�0�H�/ࡥ�\�s�7]>�l�̵��X蓶��+k��W%��H��}V�g(�q���s�rs��:�T�m����c$�wqoE�0����D���,g}�і�7��Ʈ�4X[�0�Q�YVл��bvuէ
�J�k��-,�Y劲Kl܁���MOh�I�:�֊��V�[��k�&������e�"}|5W&_��z;k�t�����!(�,���z�M��`�vU���ݻB��]��a*�d��,�
<I7[������+A�#���
g�҉I�"���r�D�P!rPʔ�>v�'�։Č�tZ�3f+��Yz6�Z�c�h�+e�Z)��O�L�F܊m@h��L����:=�L��r�0�}p��U��nLfM/�֗xr�Y���K����MĲFa|t�b���=ϋx�R��x]����Ẍ́�s|�̬	#�f5��aQ$N3��kI�;]G���੻��0w$@2�+��v�����y�kK޵������~	�$$$ E�_��� #~� ~6~%/�k�_˿Ͽ�o+���Sh�B�������`���I\�t��qڡ�7/�>]zә׹N��OS�s5����r�^
�"����2����)Ꝯ�^Z4��'�A�o ��Ř��{n�,������5�`��G���9\4Ȩ^wMOD\��0�y|�rh`���ˤ@��.V���vn�F��soz"n���P\�˱&�62�N�2',U'2·x"+1m�]*ޚ��'!u��l�Eڥp_�����W�������҆n�Ye&�3R��_m����b�r����z�X��-/AB��Ͱe�d� ��j!��.�&�:J�a��uy�����H�>�&̸����2�QV����wD��BSau+�s0�4�krfE���f�M*�&3���Y��FT*
\����*F�G�	QAdPY�&��EAB(���J"!��,��,�R�UYiH�`�T
ʓ��'M`�DF"ȰQdFDb�@Y"�J���@ĕ%VX��X)aXM2�.+
ŋHc1����)`)XETB�0��Tu�<��9|��hw>r���0x�v�>R�2���EϾ�6�i������+*�$�����=�H_�w���5�%�[�^�܍d��e�B�����!l4���W�];9�u��&
b�Y�f��C �:�D�dG�{�K�ՙ���8���ַ�!�N;=�{��Z���*���Pt���ZW>v�h��*y�&�˳2��/̞nw/uX���9�<D.��
�dPv�u��!�ݍZP�X��ų�<ƾ����]������L�_2���M�NIAP������W���M�#�׭��pz�l�����A˘�.�Sp����T����;��k��ĊNה9����}�֦$�����/F���:���{]���������\QTm3�WʼpC]S1bpA�Θ�\^�N+�Qz)�n*hY3Gs7E�ru��+$'RN��p��xjĆ�^��sf�y���Vn��5{�HQ��p�Nt�lNp�u��/3"Q<��u��8���c*O�{ �	�d����e���UD=<���}^�pv�i=�'�].��r�?^��������]g� *��,���GU�EJG/.^�d���G1̝�w/w����9��cgw6�k��,���tY�N�\���j	��O\(�6�0:1<s����e�ƭՍ��D�n��B��ў%&zM�*/E]T<=q�:c���#���R�M�����u�^C�*5����Y}v_����t^�t��:n�;$�5���8~�V�j,ӽW3�j��m�"M�p"����o#���ׁ8�Ɏ+�&\J�t:�_#Q}�s��'�2�'Vy���y���יV��4&o��,�o`)�h��R���>�uS7�j�OR�-Z1����2��0����d���r�xPTr0t�������JM���B�t8���e&`�#{V�O+E��2�ԂO��۞}�mQ@��KD�>��l��x�r���Ȣ��,G�g�r)��lk~,��B��ά>�������ӓ�*q<� ��P*pv^ES�n�tQ/�-
*f�|�Ua{p�>�n��]K.��f�Aԧ
�K��{w���I|
�\��7O�X��=�ﶹM/�6 <Cq�x�ʋC�Q%�V���n:��u���iL�^�#^
s}��[��?I�iz�_s��_Z��ؤ��Ay~��4I���z=�ޠ�x�p)��elt���f���:yK`�d.�6�tƤcXm0=C2��L���Z�+� B��+��:�(զn����dfk1� �� �R� _w��=�.�c�C��f^$�jr;��=��~���O��<d8F�+���z��6)_�ί)o��Z�1��Q�՗�k�Ii/)���ENf�˭��s)�sl�܄n\WUv4w&�>ql���:��.k$��y�]ڜPqdpu���"*�0fz���/���[x�.� �Q���p|���6	Q�J���u�����Z��\�^��)̤��e�YU;��2;������8Ҽ��'�b����j���%;V����\��E�kRi�9�+���7F��w�ޮ�(���B��F~۷_oF�gX�~���_�]n�j{k[��Γڍu�9:	�Q���5�q�\t�=m�5�F"���J�129⪎�ڻP}��qT~����t���ӆ}������L=5wh���\��������pJ=˟3�#�}��\�'������O�\��h'0�[C���~�k��̸�%�E��:�z28S���İ_���G}Xa����T���r%��ڰj���>�cıd�����I���+�ܿ�2ռS���:�`�G���@�]9�k��䃙���D#����JN���D�0Z����F=��囬��z6�$����F+ta�q3��&0��ŀ���W�q7��>B���rhL:�\WVr�/�C�f�.�l<3��WT6�$w:B��F�Ŭ���bw'J]���T�V"Mk�}�Sk7�yҘ��lR�p�Pޯq���fl�5�D�N��7Cr������ �.��W�^����4_�a>O��F���T��k;�t*>2��x�̖����{��S��sw��[�H���K��)Ŧ�WnXy���TD�'}�ǈrmv*?A�P_���`&����t��3�k����������Kl���mv�YŮY{27�	���C�Z%��4=����uy3|vy
�O�~��8�f�҃:n1
��Y��F�|ݬj������4�N��ͻ��u۵�����N��=��Lrv�ú�/)��11��ǁ5��-I����4�u�3w:׵ 4���	�f��Sî�����!�#�A��х��N]Z7�'��'��u�ю�Y4/<q�u��Ǡ�cw��� �^�i�/d4�����o���8��Z�eh����1/��~rƦ�l��r�_bk����7��劇[,�z�L��Ʀ2e��$��w�����cݞ2��0;tĹ�T��/���c�c��jXo�g�L��}a�E䮲��h���Kʭ�ԟv��H)�1z�6}��C�W�m�P�3���d.R�Ύ��f�ݭ�R���$�>��:��њj<'q������^;�x& �����cw��$_K�Eb�/�sGr���l\���E����mNdz��GH�M�(�^�b6e�Yc�K�`!���~h��m�"њ����_*ł�[��]`�:J"Y�u� ܽYx�gZ7�i�e���v�/!�1�2�U���
�zl1�#9��~G�d:�z<�D#�*���u�_0��O��'-�W��kza�j�q-3qEB.z���R@�Nnn���\��/�ˌ��g��kgU]�J5w�Z�²�x���D�8-�d�E�WvkE��ksB�X�z8�-b�%
��K����E�ݠ��g�D<|��jz83�J�
��Ա���9�Z�7\,���\ޭ�F�ۙ�v����W�lF�UH�dֿv�n�^�|���;��zh��J������|������mu����vM������XaJNeز_r�wz�|y>�{�갉���d`e�̵��q��C�iX��m*�
���R���Ǚ�o-�/�;�,dt�`R�G!��T�g�ڠHʎ��+U����.�
���.e�c��QAZ6�(:᧗��6�S��\bu���X]=2�<F�m���]F'B� k������`�U�HR��gN���э[Πsgm#wb�JӤy��Κ�gY霕���i(S�B9w�;��&�M�zr�*�����;]-�-�v�$d�EfK3u��E1���Y�u/-�0-�]�������� �Nv�V���Z�]ۡ��$4G�move��,uȎI��Ha����X���k�K5K�<���0��2�r��t�:Eq:5U쒷Qj��~���	7Hۚ��?�^�b��ݘ��j�fּ��	\)d���G����ʕ���d�q���$�u?�6�)�00� ��-�����D�r�R�f�-V,�hۡ��Pg7Zs��·�N��Vt�6T�wv!���ᫌ�����L�-�I �NI.�̼�w!Gkr��e)6�F�-Ï��i�i�C�l�	���f8�6Mҗk쇠u1Й����6pL���ܜ�;#��o%���4�\ʖU�"S�`퍇�/�Y�MG�)7B��(VJ��2K-�z���Ua�nL�o�5�c�+s;i�v(L�X�lk��`�K pf=˸�%倰�8��]���27r�Ϭ�Yb."ó��}e�;u���W�y�|r[�&�?:@�*I����b��
��,+
őB�*LaY&!�h�`VH""B�	
���"ɍ@Y4�ɉX�Q���V���
(���@1�&!���diY��X*���E���m$P(i���C�7�?Zg?g���Jr�����=<̥��֞י��S�9M�d~��D���h:w�����':1F��U��đ$j%[�W�h��C�ױj�v�����c{�����:�ޙ����.�����:��0�vUe���V�V�VD�U)���tČ�i���"J6���hm�4��σ�"yĲ��܂��Ԡ���S��Ն��3oӏ�+�z��uje�Z5�t�=�W}��P�A��*�f�3ЬC������+�B�d��Ou�a�tS'��*Tn�>!��mͻ@壭�����t�W2��pj��O�wU�
=\���u�;�D�ٵ��=ʋ/
S�[��%&;�䬯�g�݃˃�s����f�<_�Ggx�]Y�놳9|b����7�R�;���lU��XU%�.�`%�Mݧ��d=�י�k�WYw�����_M�6Vk�z'y�
�pn닒�ͭ�Q�~@ް�;��-!�ϼ��=�r���AC�Yp�H���By�b։�.1�T�^�)&d�����nGɽ�QF����J<G�kί$kG��{�v�2h�P�@� �}x��[�!Ж�����;;ܽ6�Kg�I�O��Q�-�~�v	���C+�qon:5�M�ik:��5����ٷ���5?��T���y?�_Tt�7�n���4����M���0ĔĖ/�ÿ4=�фb�R��G9�QC����TU<�1�;r]a�:����,󏈥�yi�ѻ�w�W���z�*Yћ�}��R�<כd�.���qޭ����y��_]o6ɬq�z���;4UYz�:�ی�ˍ�3܊Y��f�0��m��Y��]��N���{K�|�uT�7��ފ���hf�Ƽ�Ȗ�/�t���h>��u��h�nQ��=~&���^��x#�C`w��tJ�n���m�h�I�<I���q�7d�j�2�~�|k�l��O,|)J1sރ8q�w ��7�BI���r^������?�ԝ�0��Y'̚�;fs�	�!�%d;a�P큖�<f��I��}�������t�>��=@���a�;a=d���'�,'��&��� ì�hx�vô��}}��3~������>�Vg�!�6��C�Cl�2|ã�l'��!X!6�����I8�C[�BuΎs�}׽wߞ��$�$���C�p��=M0� u�!Ě{a�����	����$� �M��{ٿ�}o�9�VI�d��z�Y<a6�XOP:N��R�$�L��I���J�!6��>��u�_{����2ΐ�!�'2��I�N���<d�5�;N0����R�C:�
q�zz��ﮭϷ�s�v�4�s��Y���L9Ld���I;d��)=d�P�d1t�9���|׺�}��~������$��z�
t�2`|��	��AI�N%B@��o�d� �XO�i��ޮ�p�����}!�C��q	�O�LBu� qq�T�q�8�I����6�{�m�^kW�ky�|���>�ԝ��Xt�>gۤ�'L�	��2����I�!�Y!|��	�1&�N�,�6����/����_�;f�C��S�Q*u�%��N��x��!����~��1��sJ��+�d�S��8,���)�M}�����$=��}��~�!����	�i���H'��!��V�?�!�Co���g,1�i���!��]o�k�� x��N�d�&���2M=2N$��x�4ʜd��̇��!>d4��'�:��w��{|s�o~�$N���&�O6�z�8���	;`i��'L����&�=d��$:�{��5מ����N0�� z�l���OXOy`q'O��d��x�$�!�6��,Zz�<C���y��>�߾�H|P�`g��I�CGVC�O�k�|�<��OMu�I:vɴ!�xs��CL� �8}�o�}�����
��2�Y+$�|���|ɴ:d=d����&�<@���(̙Ն�'l�׿z���5�����C�q��i$�KI;I�kvL@6��C�C�OuHa���I�&06���=���g;�|�	;Ld�$>��x�=C��(����P���!�tjöM�!�L{B�=a0��_w��ў�k������:��=q ��r�̓�>a'�����>`h��M��,��L����z������~�{�&���!��0�@�,I<d=Cl���$�h��M�T�'O����_O�2��w?�۱��j&�5<���@�U���
;7j����A���Yx�N�]����I��aB3�]a�t2�EA㜹~}�{ލ�Ӥ��#�=�0~C� �2$u��m�w����6�m��I���M�!��>����k���>��w&�4��Ї�1�$�!=d<��T�>I��Ci7`��I�AI��r�B�^gF��[���=�����ɦOP3�Iĝ=�!6�bH�4�2?0��6�*{�>B`m�������w��_o���� ���j�K�l�;d遅��$���$*t�0����!����C�8�����_h����sf�!��I'>��a�d��d���I�I�L�B'ILM3_Y;C���ΎW^�����oϤ��@�8wN�!��>@�M�4��'|���i�$���g�����$9�\>���]w�_o���>@铴6���	�OP���wO�C^�<d�OP����'L����i�0<�^f�/g�������v�s�L���ud=`,�P���H0��|��\�6��M�z�4�y���:ϼ�۝����8�0�3�%`[@;C�h��&�z�X����6�NY�$����'�'[�M=��{�9����~}�7�!�>��2Cl�I�큅���XC�x�Xd6��7Ր����D}𽒝��_���T�tϯ�b�'N��
���,�g�0l���D~��X~>��G�{lm�Z����J�n��-vH+(鋤�i�?�}��Wԟ [��$��$���O�v2OG�Y$0d�!�$���;I�m��KCi9Ch2m��|�s�}�����8@����i1�����	�8ɭ�m�gY��M��ߖ�R�<I���:9���7��׼�|�4�P��x�'V�&r���5�O�&�@+'��vC�&����|�z��}���0���s����v���d�35C�O�3��O�VHxwN!6���O�YBz��*d�Iw�ߝ�|���I�d�Մ��a;d�>d�C�+�'h�o�̓�+k�����h|�t���{����}��}������15�!����z�L�Кd�>C�2N���=�ֽ���}�(i��� �'�Y't��0�x��RO;N��z�i~HX'�;`
�vy����7�9)��!����0�<�SU�$ռ��i�>e��]�ߝ(���v�F�;#p��6����ӭ�M�;��>}��fp�U�e�T���D�e�Ʈi���2p[.9������[�N��B6u��x��~1�U�{l��N4P�s��ףj�*�HIK��Ͻ�z(ES����3s���7��1���F\6��h)�����e+�W�g�F�3޿���üw�㔷>ܡ?#U�4��`ν�����士�6(�mZ3�Fi�F/f�ж���߅M"c>C*�Y9
�>����-�4�GB�0�״�qs"c2�cEϵ䞅���(�=�a�I$��0Tp�j�y��/��A���8!��hmR��}��u�^_z�%sTn]�0,뇰�C���k8-;1���3��>�TQ�q�Z��,S�� �u�)��!�f�T≩wW�װWp��ǈ�%��'?�U}_}Tr2Ԇ�o���q?YL<����0����|2�ɔ��[C��`���W�X�d��HR��CL�F+�0��S�˼éH��9��U>�s�=�tL��._m`Y�7:������|�ͽ�t� ޖ�{�R����,��>R^��[��. ���0��+S�8�٫�N3Zl�O(��:�Y�
��ˤ�>����(\xZ�^+x�B����։7�׵��U�+�d���_uz���h�!�<��n���8�z%3]sF�s���$"{I�5W*�X�T.7�jSCbo���K�w�����l�W	%�i��
T����J��k�7?��}�A=gIe�:�ۋ�=,��Ր�9tR�5#��|��)��{{�v�0��<�{�u�!�𛆕)ؘ�U<h�W��C������R��c�77�k����3���2i��I�dx6�7�'��믄&��>[C���Uj���2��t���u��H�<4�	�mF��QSz-�2yk5�luC��j�"烌��ek+���iS\���u�K�7c��m�-�{�������C�y���~
�`���o���R�l	�uu�\�X�c�E��w�%�߰��uu�MrgnGn���C�ޘ�L��ͰҴʓ�.�սT��V�;b�ԝ �j��aYW�'��[;�1x�og�TS�*�\���D�K[[e�6����^�}�SPC���Fwl�Z�53s2��Q,�OϏi��6�Y�I��R	�v`M�G���t]-��f����:����wL�	%Ck�J�+'.ś���ǛF�c��.1�K�N�]��})�j&6��Z�߂{ʯ�-�c�	s�+��+�Lʾ��y���'�E�ǎ��Թ�{����o\�����5u�4�]��Ga��z�L���Q�{�d�u�.�4�n`]J��1뫨���'=G:��T�*�+����7�<7`-�G{�� �H��Z�^�gKlҨ���'���̈́X`h�u��fO�gN�=z��:0٩��y2r��E|%�ά��&�e�����;w�w�\�0ET��:ȱ
�^�s��U:}�2�k�L�)��rK̩M�[]�p�2�Ei���:��D͉`�A'��܉Mf1�% �}�9��Y�h�7]�H�r���I��,QE�����ueh*^L�b��R��(�˦e[K��Է1^���]����bXc�R��7"��WO��
�Mf@�3�8�8H��f,�f\��u�b�-NY����p��[r�ֱG\�r+��w�관�׷�ÔNf�t�^�vӂb;6�Pc"NOPH�Q��r&e��m��Â}g�*Ê^�v�*�g�:�t�S1��~��"�_�~&��O~����c+C�GT�B.��C�HMZJ��	�cf�b(T%I�J��ɬ����E*]k��+�Z��E�IS���
�t���=:dή'L&���VH�J����YP*�i!P��R�6�钤�aQb�(�,Xt�����4ԭdS�!� b,DE�dY(��<��_���[��{���ձ�բ��ı��5���1��*4��K��z#��V��+�?��Y�W�z訜�ǟ����,w���eP����5�v�z��f��Ɵ]�,�]]��<�iS��e��4������zy��[W�W�\�ɶE;pI�;J���#4�I�|6^e=�{/�x�(�xM�����=t_-�I��#��o�1Mڜ\%C"8���!ThC7;�=NX��Y�SΝh�������x����64;w����y�)I��O2b����	��u���K ������tk�a��
����3q��N�D�{�x/�8h�]�Y��k��x/�����5�����1Bd�����ﾤ�k�5q���'4�ܯMS�$T�-��u:���t��z��E)���G\ե�a����g�Q�1K;���|���c%Z�h��ˊʬ�Wi���#�ZW������}3F��OgVD-F�⨜]��U���x%��>����kp��������U�>4(F����Ҩga�O4�M>���B>h[�}��q�z�]�/z(�z�j#��zz*�ή��
������BЁ�X�B+��i*=II�b֊7�T�X;[r���q�^���Q�Vȷ�~fc ��y��HXV���ۈ��}�H�dIt렑H��}U���T��Y�Wt�����h9�zA�Un�^��{���3,�p���;���{�Jl���5U�lRt��NM/<��#GW�u�zD���ڎfn���rG8�#�x��f0��|Q,���XV��r��)̎�\�p��(1-@��|����v'W��h�C�^��RN*W�N��Ow�ی�@W��X�-n��"&�nE ����:�ѯyxLM�C�lM�ۖ����v��35L?�8�T!Mg�oS�.ʣP����5g�3Gk9S3�6�Q�	i�gi9b�^
�K�	��Z�ޥ�5,r�?�U}��Ur�H�������Ot���s��bqco��n�;*-<��j�Oe'���ڱ�X�r���m��d���Yg|�� a9�Quv/69.�@U�-��!�Bkס�kD
k�M���z�3�	BW�?hl���M�0B"�Ӟy�$��o1������	*S���7я���B���� 7����qҗ&��)�먵;Q�D�t\_E��i�vsT� �
��mu�%N��~���yAct�Ȯ�j��R*d�%��>0�A�F�N����V>��ʼa��f�/�k�G74���Z[�s��T�G����M�q*'�>�M��!S��y���#0�NTtkq<�\hV�>���o��(�/�e5Y�����S;��.�}�ڌ�@��YF7����[��n���˛a*xk7�8�i�7P�w�__&��U���R���1�y븱cT�(�|����L�@�E��=�|
�܌��=�,1Jv5ѿ�{�y'������a�q:�tyZ����C���o�U�ؚ"��?v��Ʌ��{b�XZ(���e� �:y[5&��s��{�M�s�gJ�)�seӺ�Č�D����Ѻ��:n���"=W��$bz�s�w*��D���s2, �aU�[����+4�Z�a(y|�)^R�t�堦�x�&M���l���]��h3[c1��������MeM,�Ӟ$�H�nP�a��=8֦Kx��i�΂F�O+��k��O;����j��s�S�7��C%_{\�Ѻ"����5��i��6דAU��Y�w�hYG7k�%Q������{��Y�������S��3G]��Zc㕞�0C�:����-X�XyfќM=��Dݥ:�7��*�R��1��3ex��êU�a�WޏG��]|I_V���7��<��!��FjE����������Mh�5��|\V��0�r�o?V�:�/M�;n��[x�D�w=~�����p��XL�0��MV�3��dQ=�
�-Af���F/�w��J?{��,ђh�Oa��,"Q�Y�;���NJ��CUc���{�J�|���E����g������O%4�ٱ$�PT��9�6���/(,�:�"�VO:�w�(��U�K:���l7O«����-NF޽0�uY���X��zwy����U���,����W�nv�ڛ��+��5�ePɹ'mR�q%������.R.����W�N�雌Aщ����>;�6�C�2��S�0-��v��SX�����N�5�E�ڬښV�u�d����7���V`���徃`'�����łV$o��������]����F7�W��*���W��K�6��'=��xh=u����}Fr��]
<�K���v��	��}֌������L��j�=��B�w��"�e�<��q{�}�o��;�kZ�?<��Pƪ��[-g�����;w���{R-�ۥV7^n@�w�H��0du�Yy����2)i�ۧw�BF��l��,������t�C�C�0"���!�@̵�-����m�װ�V�2Y���a	އv� <���t�mw���*l'o.��:E�(�������;�mtw����N)\���k�Ȯ���P�J��Ǔ��+�s2���I��vt��hh}<[��[�8UL�R�YL�+�
��h�J?� О�t�oP��j��-g��7u����7���{
�<h�v-�'5B�D��W;�un�i�͡�>�>�B��qt�ƈ'r�WQ��h�X�_j�;����Wo:��dW����H�BWo9J��Wo��r��r~����YM���ږQ][fo皫K�ḛ���kfx������b���f��3����&����:���B�;.'6)ȡ[G���n~\]�W��+����ϳ�O���v��G�f�SU;��)�D�0��J��� jv�Q�+U���ݡhQwU-v�- 1la��� ͢�cW��r�t_5^e�gc����Y{������g.ܡ�:�U���O��./`8�m��D2��DF�ao�P�c��|*�_m��V�5��2�×Av3e궋��E�Յ��q��SeX����wķ���#æ<ӵf�<���UbK�K�#YA9�Z�a�Ø9J����P��P|��2���u��r�D/�2E ���F���Z��'UM��v�d�p�]��Wt@�ԾZ��T�F݇jҁvB5U��R�﷥Y�f���U��qf^ɗ��m�KL�k��m�ۖ�0v�qV_'Ғ+:\i��cq�{1]�R���/���'�p�Z�UO�,��ի��+���*sU���
����aY�^�.�J.Z/�^vNx�K5V�<��oh�!�A[���u�ero����=���zY�iJ�];o��*w1�8e�C��u��ݚ;��4Z����M���1|/�,��{��j��)��9E]K#��=���L^u;ȕ�a��%���5ᑡ�Q%�eY�6����rP{-ܼc{O��U���ɮ�yK���w����dM�"G:c'���V>�M�v]m���6Y���Ռ���'Wn�(��X9E�N����Q˺O�%n�%����l��c�X��!T{������5��H��Rok��Vk9ہ���/s:qGM^1	�����r'�r��yw�ڟLXLݒ���ФS*=Σ���V-��T�`% �q�NN�Ttg[��I��!+d˫��.U==�W_XqV-q[��/��\��{3�%����/,	�O7���Ԗm#��%�����n�"
�fֹ�/Lo�7:�������1��N6��R��Y�J��vm�fs=vob;�:��`�\a+{��G�AE�'�1��̤q$PQIz���e�R,��dQ���W�b1"���jt�*��V�Da1�����J�*�B�e�Kh6�)U�%J����kR�ՙ�*c
�J�+R���9�Y�0qX,*LeLd�`��\edPY.Y*��ũU����c ��T��Vc+YXJ�:̐�+'I*Ed�	�Z�Qea#�~#�-�)<�E^?�B��{�e���d-���v�Yܝz�l�������}�"�O�(.�K|��(��j�^9Ֆ��f�I�Ō��M���qp{i�Ʀov��d+R�?~~bL.&l���5�fx/5�9���n1K^�5� �Z���c�=4��A�ؽNm"���*6�#����3~ ��=��"�H��v!�Ƹ%��w;p�^�HY�:3|j2|3:�a�g�OD�L����]g<#�~�F������9�+�R�j�Za�IW�����W�z�U�hl��e�h�#��6*ݧך��/���Ϡ��x�:��-=Z���k�%'fV{�K��;�Ɛ�9j�k�N�hW/�v�N�=0_X�!:H]�IW[�4��OM���M���yl���K���7P��bf`K�9�Y�<���6l�N��d)�JDI?P��w7��-8a�YDt��ǈӠ���)��u�|BXj�9��4��dY��~>(��4�_i&_CgZM��wT�����*#�ԁ�c�a�l1���q�P�]j^��w�YgN�-/��t ��MI- �1��qԳ��n��=Pi�9i�F0��z�0R�Q�dTm)�i����)odNI��"mq\T?�DO-2�9JZ/&%���������w�����2�إ�Ex���H.c!w�7��1��7o�̭��\A��.nrm�fg��tԴnwxTC�>��v�W���zt���Q����Jo����-�,u��h9�$KŃ��W0��Ʊn�N���_�=��^��0�oR�eb0fMq�l9u�y}����zv��$�@��镲ɯG�u�ʑ��^�:�Gl��b*M�qj�v�.���ޏye����*~��
�hW�a%���6v��de�Eg�c��j��s�V2aF_�D�`��8;!���2KZ�ws��y\f�ȃ4t�7��E��ֈ:����d��Y�>��S�E�`��=xf�,�8�CN߮_��)���X]=4Ĵˤ�C��Z�[Q�}ˍ�A%�X7e�{��V~�<�R��rϚ�>>(�!��8�Ӯ�S�950�R ���DS����[Q#O���,{��ڋ#)(��z�ľ�Qi�<P��Ly��ΥW�ݚa�aYc�;�����v$�_q^]=�f	�c���f�|#��cǉ�d� �k��e�}���b����q��pټ~˫�����y����9�:����l��f�n��&��m�u)ZR��ۡxk�Tw��D��~�G���R;�O�*j,E�S
�ǣ�q�H��9������ە���!��-2�4GD8���i%\tͧ��'��ϻ�v�a�y)k��0���<���ø51|�|EZ�@�B*V���R9Z���8�Hq�g�g	��EOy���{��#%O�wy�VMĉ G;V�*�L���j������l9RѨ�4�R#K�`��(�5�D�׷=	�+>��NR
Д��c`���a�;&u�)�ږ��D�	�ġ���ܵ�󽿇��Φ��b�ۅ�$��GbH:D��k{�	X���G9q�~�ޗ�I���ﳦ�s�Hy�'b�(��m^�����R�~�VY��-��a�zo9@�^u|��8��P���
�{�m�]gi�z�n��a���$)Z���|�ɛ�b.TD[�������|2�}��ּ��&_�a�7�ɠb~�=Sկ�W�_�dQӞ^>#�(�7I�cK������ՇO����w̃���Np^8Fכ�uLax���wo9�P۾�m+�^`� �>?i6���0��t{5=��XQ��6G�1��B�Q����9)������k�J� DO�
�ڮ2�6F��tzy�x���̓��r�y�ڡԧ(��R�>~I�l�[��H��[�/>r^�A�H3��ɸ�Q^��<"o�"G;3�J�y��yNe�3�s�_>0zޝ:zf�}�2ҁ!�Wy.������85�F��c������vG�a�L���+��uO�����ۦf�*ȼ�wiF.��I��#�,ŭ�ۓ�0k��8�/�Y�ذ0����4!�pd�l��A��}�Ut��&��;?�1�G�YC7k��w����;Xl�n]n�Fx�GM�F޶r����g�t�P�z�&�U�k3�MKB%�c�ڰÄ������:��-=�	�����w�,_s�d�/�)�!�r�	&M�C�o��w���X���&np�����95h,b�H�CE�u�w֖�108F�Z=��4eH�0e�$��GJ�ʶ=ܬ���1�G]1�P���l=G�Mc�'��5�\�i��Α�ĝ>�UУ�.kI=@�|x��m���5u^����x��~O\p�&a�zT��{�ٳ�ܴ�j�ϼ�B�eҠ����"yi��ydQO�HF�#�1�TYu4��t��l݀Л�ׇ�+��7�+H�Ƕӹ"�K�P����j�z�Qei��d���I����4@��w�kn��o��P��O�[�����"=���x%z����c�"�t�?6a�!c�X�}^�p�X���L�fs����}�� V�HNX}k@;�	8z��o;�yѭVY$o�k��4x�?^mt�
s���d^�an�8��'��L�/��*zfm�z�l�j�+�Q���[�U�c��H��C)�l��x��6�.ؽ�^{z�R{*��#�5���(�q!W��4T������'�@��<s���Ն}���9\��ݙ��a�!�_����ei?e��e���#1����fLU9�d�8�3�6�"�|`�e�Cy{3t�GƥAL��z����Qv�C���Q�~u���뷂�; �C��n�+����A�36Xf��'�!R[͚�"W��A5�Is��?I��2 ����
|��<h$7LO9z�{]��HG�iz���E�7��^N-4G�Ԋ��ng]��y���.>$�&/��z^.5m���!������uo����(�\ǎ�Z�P%f���6_���Ӈ��m�O��)hT��1c}�S5�M��4y��Ax����f<��{W*A>�dd�����:I��N�d�\Jnf{@���!E-tT���g���t�W�vgs^�^hX�������X�~xf.�#�����as�)�/җby^��a��}x���#:t�&�w����9n�v�\a���+W�>?qb_a���Sڸ��4�[�^e�{�����wޡWjXZZI�}�9���}N_J�ȣ7CО;��L�K�5|r;�r�����萊8��'��)��)hJ]�m-6w����T<nö֥S!Ȏ�31,A���K�y�g#�<!��	���6�ƙp��La ��iʂB�Q����Ze�%�S}�H�;ۓLI+5�${�:�����3p`ogom�{,8���uj��-iIa�_[@���ӭ0R��μ�H�ADx��c��<bг��UA��=2h�L�]ZL�"yҟL�`h\^!�y��7��z��y���a�Gx�yV��	�@�>4F�����1*��{�m��EZ��q���a�f�P��-	�;�Ѯ [�(�^��8D?&�!�XpKp�C�e:>�b�
��0�9��mǦ���z*�0���e�᧟$q\
�c+�tl���u��V��P+�l)���t���n�ܬ�u�����睊m�=*��ǋ�8�.-?|���
6z��g�������M���&�TCЈ3�E��^��WuL�0�/y��	f�ߨj���f�z��W�~DÉ��se����!��&��4���a�_:�dX��9�o���ｘ|�|����\X���j9�DUW�F�h�7��܉����͜Hj�@^��!�;����whxZ�(/����TE+;����L��>��1>��	TWT6��!����]��k�N����/��R�?+�x|x��(�C_�<Ej�p�P�V��(��
:
T0[u�fK�.D������D��Vw������/
��r,q��i�:{�$A���;ك��+"���ᔕ�;������C,c�|���t��B�Tߺ�Ϋ}�AF-����1l��nj���W�a�p� yz�$m�β3�ͳ�f�9����૙��E���2�׺Sb��G{xCַT�De�M��GoQx����SbI�	�vh5���gY	�9k$f
n9V���Tw=��eA��*�gچ3�ʸ����!�Vbh�y��u�������Z3fq��W��j�դ��`���s��&�lP���܃.7��u�ґ=�O,�ˢU�]4��,�6�2K��o/2lǋ0���,VH���Z��2�I��}�q��Q��&e���L��W3�cbB��(��+lQ�,+4��Lf�L�]B�]oc�NSI��]%7�:w��Ҳ��6-�Wc;��;���O�=]�n��۷X����J�60Z���aضwr�Җ��Y=͝G&�D]L�<_6`�f��(��̺۝���C�Ik)�\�A��#�O�ڻj��<�"Wnp��s�U啡SnJ��K��j����8��-�t���&>��ًxl����#a���+ua�`YX�fA9!�8�W�7huoP���/�.4`��u�N��:�9��Ս�&��K'Y���v%�z�ON�ĵ�|eR��Z�;6�8.6��qdn���,N��e�3��E`t�(������v�9�B��V��&W2�͔��
�P�w(u���q�;�OL��ޥql��#�^a=+q`s�6��=M�W\����'ď�$�{��Ad�J�UJ�m�9�kYRc*(��Ր�&�gl0@�m+mm���f*UTQĩl�&0�j[T1
�\Vd�s.Z���,1��%c�b��.9��1YP*��X���2f6V��XdH:��QIneE.d2`�fZ�"�1�bG)1
�r�
��c��eLq*bAB-b%L�kF�X�*e
�/��� 6BD ��xG�W��oTtp�J�r�a�l}	�7����*�E,I�~�����V�ON��(F}�
�TA�_�Ť&�˵9�F_U�ogQ��r8Y�d�>��|E�i- �c�ǻs7޼�B!:�!�\|p���aG�D���޼U1��c�����
k������."��~X��!�͜t��uo���=��p�ÕL��V�vwO�[�H�L��C���w~�i5]!�H����1q�P�*=V��)_#��/݄�K����|ǎ�?^�-�\���=:@H�.�W�kێ�F�I����԰�2�.}W0��kzm�yY�^�i�3e���A$������گ�����SD�ࡈ�LL��^A����E{��m��O�Ll��f9��ZOݝ^�eC*2�|$:7Z\�,��2�,s $
�i��{��K�ٛXHѼy\� (�_���P���ha��mz׊�l��>�,�I�8����n��S �a�X��@t���;���z��Xg��]��F��4E�x|�����?e��e��������e��>�g�E�Єc093lu�ANC ���?�
�|�SK�I�d~��%��ؖ��r���u��l����*3LG3�ΑӰ��ra��]y�=<$-�3�ӎ�3)ȍCƶ�����3ۚ���g<�Rh����\�yi/Y#H'5
5I��{�4K�/�µٜ"��E�
cxL�
Trw�>�fk���({�Jd�5��M�#0S/�C��k���	���W_�d�!���u娅�l�m+�������^�a�EY�'m{��m��$q�SjF+rPc�S)�&irj��r��'���q)?�_RZW����V]o,�Q?�)�֜���8wJ
����UmfnA����Zk�菓V����qo����&�e2"i���S�ew����1�ϯ4
)!������^J���&Z��C��������_qe7���C�����ۨ�(�ӡ>8}�;H!hJS���Ӈ=��W�+�݅k�z$A�;kM;���Y����W爍�w{Y���-8F�n��B���x:j��kxQM�7c�X��#�ύ�����;�;���O;eUv�Ϳ{l;B���D�P��]�l�Ia�U���;��*%���)�0����2�xv���/Mٕ^��&a��r:��Ǹ��Wp���u��o�$<;+������šl2�������+Ϸ�e�"ӽ�(������O &HM����lQϺ���F�-۫����gH_��ͧ�k��D3�k���'�yJ�	z��|~�q�!�1�;z��,�>;-؈?!��BG��c�gyw^{U�O��cF�����:騽���rz2�^(�8�yE"�F<�c9��x��- P��𲍟mZ��������ֆ���)�ֽ�H��7���9�xD�X<�'ZM��v�ɕ3ce��k
^&zU�=�3#�d�#��"���W��Li�-9�h��2Y,W���]��^g��,�&׏�1n<��&���a�����OhzU���b�!ۯ�m���Hg�9M��]2�g�Ƒ�*�y�OxwgV��R�F��a���[�G}�����m��G�N��[]���n$��&��Ν������<�����(��Lse��?�bs�>�b��+"� ��?����0>�^>�pߧ'd���"9���p�2�Һ�]]2�%,zw�Dƺ��;�4�����ǈ45���!�M���k��k&�fb�Ș�W�G�2�#Os��Z��6Oa$��>-!6�n�O��1 {��dN�md�,�9y}�#�Q��h�l�Kz\��� H��1լ���F*\`Ƀ3�P�ǭa�!����:�9&��U�یoS�<!�>:x�-�Ԥq}C�y�=���x��;�.֐N�G� ��f�os�{o�~h�;ӆ^�=LD���9WT���]1�͘o��ǱC����l vf��s, ��.�j�ظ��ׂ(z��eoHNTO>��N��W��hQi`��K�W6�k*􅆕�\;�r�㮝aI��0H���X�ħ��0����l:�ش����U��i/\<l�TYiyi��Ǝ U��=�7��\hќ�=�i��&,v|�G	6c�'Mg�ǯ������FZ�^{�H��&���ݳl��=�
�P�~���jԪ�_[��ߌ�7Bސg)<��V.��<�ik�)�Oŧ|��@=Xy�m���:�����6��3�e��x��Z�[Q�k���33�e���mi�a���g���жy���]Yw��4Fj�|��N"ϊKb�z��Ô��7Q)j`��훀#&f6T�lGQ���3zk�g�E=ei4p9z�(뫥A�Ȅ��տ/�����Z�����_��J�tl]��έPģ��Ѩ���z+d�52f��%�+vr�)0Qs�	:H�_�{��+�Kwҳ���z�Ϟ�v�_�4]V��HG�|�>C��Qb����^�F�K�Q�%#��9�q  6m���FI7!��^"|�#��S�,��d��bG�k%8��gJ�O+#)6<�kI-e����?Vg��5�#����qB,@�:�K�:M^L�UKj��Z��xXdV,8x��K#��X�z��^ �dQ�d��*@=w��tNG��G'�J���^:0�H�R~�*�{suB:��s��#��p�!�������6KK�Ε�đő∷�N;;H!hJS��8�_��߭ښ�~x*_X�d^Q�IP�-����sMDC_�
�a�O'1���CVO[�1�����,�%�E�"�y�#�	=B��͗�;fj�m�"���X����/zs��h�9S�l�?}E�Sq���ن�S�j�] ���#�.+���|2�����4#t����������d�܉��-��U+��g�_��v,hcZCZ�xn��ɐN/L+�כϒ�ꘔ�24�L�=�OkcO,�Fs2�y~��-���O�"y�Q��=0Xe����㜧���@�5N��W��`� �]8�4�:����յ��J,�Z�谡k��n�A��)d�3P�*���#6OC���3q1��]��ɦ�Ӟi��<w ��z�VL�o�0�!1X#��Ɨ�q�R�_����0��jy�_�3۵�ƭi�2�. =��j����{[`�5l�0{D����#��g�1Fh�(������<M"Y|%o7�^W˥�U��Rn0fX'�����Ti]�嗨ۮ�}$�)��ϓ�e��}�Ԍm]�~��_�wj���>3%�v���M�zl:ӆ������i!�y���F!�ܰ��q��Ar�cA؉��6_���M����b��~��^�<�2��nU�n�����L ����$f�r�ڻ�6��[���;b�s�B,��:l9\6nvG����`:9�Ž{7,*3)iت���my�XF�1�ar�\�}������v�+�'�X~_:��~^<a��hk�Ϗ�u���]��[�v+,%���j����TfةSR��Z�[G<��c�,94.�cڎ�ʒ+J�b��|�z�=f��0�|^����þ�>#&���kω���ʢX>먹g�s�=f=�)��[������\bm3��1O�iORXgv�u�9���~w�Ǧ\��T�%.h!bK��d�Y�������>�CTT�Z�>��{~�o*M�^,��>�,v�*���h8t����jR���YV&��{���)�="~��Y.��q&��D;���HjX=����LH���&��`M[�$Y�C�.=5��i�W��r�u>�H��g 6��#�˘� �j�һ��n��V���p���5E���-55�A���NЕa2�w{�_	sN�3kj��(���������&'�n.��bқ^�G+yhxVw> �`�#�g��O��[���<�ç����4��z-5='�E�A�X���ԏ�Hg��(.|O�@�Ҧ�ɸu�wѱ��GBl��W����3�W���e �f��T������A�tn��Y�:^6#YSv�֬,f7����TeM�³dõ����"�#Z5�m.���З��;�;fq�yM&z�,θ\͒«O��xYHu��6E���ݼ
������Kǚ/�=�t��֪q��� ��9#�9呷D)B3�M�L���fL�N�Vj�w2�9U�o�V��P(����M�C\���z���J��i��"ù2�;��3��[C]�Z�x���sܩ��F������J�t��rn����S�X�XE�M��.L{G�tRgS�7���4�����L� ��w�L��%��+Aq�ZU*�.���Yzv덐���Н��&5o�j��w�A*�t����ΰ�l�W1�oS;^�1Rt8ݨZ�o��N��ہ�s�%¨�i��ܛC��p&R�Sf���v����ņjz�6f��l�ãs��W�����-�=Rn4�b��VS�� �˥̸��o�`�Z{��(;a�!�#]�mQ8��+�v�*�^	��<�f��R-DU�I�����!Ӟ�9ٛ"���n�v����އm�\�"�k���!*@jm����0����K˼�꥚��/�B@����nQ��P��Vf}�6�`��陴��y����V����e��k	q�9`�ں.sֲv��u��� �w��.������c2t[��5����{AvKrBDrێHܝ�g�f�V)kM��7��%faD�߬��]�q
?V�0���1�5�,)�
 ��
�a2�4j�l-r[�*E��B�&�*��
�bQZ�q�J�Q�,�B�bTQa��8�C)q���
�m-,h�-h��(��n511&1�f%��,Lj�Z6���L�ֲ�ui[3�dƫ�U����۫r7-N�\�B�B���.��V�3�U�����6֡P��c������ƣ��.�-u�LZ6KD�Źl�5h�L�ʋi��r�8%J������|��*�b_���B|����O8hĭ4J�]�r�-H�Ox�I�2�'���ψ�9K�I��#��5�<���)gU��E���_a.��}��R��ו4/�с��:骽��dfh�ĵD��v����}��T�y���^�$�y��4��		�H�M!����#�@�4��n��$�z�
���5�Hb&n4D�r!O� �{y=��xI�C��z�jޔk�����D� ��%#W^��*�qrZfWO���5b-��07�e�R��\IH�Ӽ��e$z��Jq!�g���2S/�Gvp���ɻ����6�D8����-�6�婂�c]�D(|�)��QC�1�EZ�L��8~#�Xi��MY��'f�u���uM ���X�BO�]�|sy�B�ڊ�n�ɣ���nNč��t�`ǹ9ǔ�۬�';&��r�h��UNaG#�_�c��7Y��Ј������^�="O:�����\�s%��L��/9�mk���`<F�@��ܳ۽����#��9p��㴴��BȔ��mA]9B�,�_����6p�,�$@��嶴ծ����i����%N������h�W�ic��XG��w&K(oU��-<��-5"\�EZ��3#�t�܉ޙCjV^u&G�t�=�
L����f	��Ȱ�8L��mwt���q{��!�l�C���c��5�g����ւ9i�,맦��<ǧ�:t\����t�]@�7��r�v�+�I-�<�ʹt���q��x�%�w&��A���q�^��a�?7)�sj3g�gv�&Զ3%�^�o��d�X�����6n�H��Ea���.T�T����"ܭ�ܻv.��vlZ�vUL}���&V��)&��D<SȘGy�g�R����Ze�{sJM�90�ع�"�u�,Fh�ML�b6'��{{[-��.l�)���U7~ʈifڋ���s��͌H�b"`np�3����j�6���V=챆�{�ӟp�C�!ߟ�"��Pf��3�GVk}��?m�� �H8��Z���w�x#Hf�7��gwz�J^����)��M��e��=l��-��b���G:˅�H�c��(�ߢ�f��՛x��O}��k���z%^�/3反b�_7�o���lCт1(t��[b�p8n�;RSuw�78$���0�6���c�E`�v�f�(s!�n��+�J\�*���G��6�K_��5��Nߢ�6�F���!j'�#���@��L���z�GJ�*I��hk���
�n�_a��Z���I�jRCU����(nmU�Ҹ%������%�_CgDOS�ϕ|2�0oykeC�8��13�g�&c�&��p\3�ZD�î��ϕ���i�fB!G���'W���=��½���K5�e�r�rcX2Ҙ�t�l�49k��ԥ~����������NVnD�+�x{�LѺ��Ij�V����';M���y!].x�rۦ1���[K%�D�仼�`^ؾ��jY��s`\Dt�b4�9����w��+�_<<@T.�l�TYiz��^6)a�O/Uy�\g�\�7����t�gZ�*�"��-��^���S�6�����-�5�o�����P�S��GM@�]��ć2os!��㇓Nc������|�&�����7�<6].�^�0�Y���$����Ð{�0FZ��f5�30�`NAm��[ݤ���)�f�?->��r���u�ŝ3��ݙr��9O{s:p��͞�������J�j-;<�������}�����XX#�|G�Ce�6�ei���鉦�b�<��T I!Kc�3[]>���4b��0cq��u,jg*`F���L��yX|��N"Z�xn/�]�>���'�mq8p:��/C��!���2P��S04�5��;K���Է<�1F��9"��<t�<p��(i�/�|�����!ش�T�!���!���\ǎ�Z�}�s��^����ˑ��o��;A+��<P_��+F�N�컲�ـ*�iw=ަ���7��$� m�7���g	fG��`nS͚̒O�|�8Iy&�}���k��ѓ"z�[2�>+n����Tg̑b�����Օ�N�$<]�2��Df�x��8�9�5W��B���gNE��i-"��
�Xy�Nl|L����.z��G�C�qڷ}���[ٸ��_�')l���G����.��j;�e���Cc�[����D�=��5��0Rǘ��x�[�$��Q��gnr!E����(��p�;t��,�He�m�{8:Vx�ti�Zm�P��"����B��`�%�I��O�_,B�Ok��3�9LW��^��;;W��0ңg�{g.5�L���|t�%f�$�;\�Җg���S���d�"3���rzۑ���Yn�}���Oww{�]�Y�I������^)�Pȃ�(�r���֜�"�;�r�a;��}��ݦ�G�e�E{��"���|��.��w~�{��^��_���q�
d?.=�OccOQZT�C<�wx�}�����ޚ?X�y���:k��ɕ���g?y+���.�arlg��0N�WI���/;{j"�Z���&�;ج۹�Oeo�������yŰ�<�~��"jhw�SȘⳚ.���mWWL�T��-��Gsg&���nFW�������JZ@�un�oz���9�Q�԰���H�L�}����������+3�p�x� `@��O���]*��#U)��f:U��e"�h�q�4H�=�Y�	��e1��=,f���7��ᨰ������.�`��gWX�hyG�&������^��,
IY�ÈoM�=��b�w}�����i�T��I⾏{��q(���&�a���&XQ:���Di��<�{��5w���w���R�xl�l,6I�@)�ѹ ^��X}�G;h�*]�B$<{�񳮸D!�����b;��<|O,8)i�Z��c|��#v���`�^�T�{�t�.Ac̝.[?*+�q���#`�h.�۹䍝#���K	�4 �5Kܾ�k�`�����]W�ݹ�E����I��Ϛ���j:ıт%�s��eˣ�VtX�J[�<A8t���,%�}.����~����&��|)�/���uPli�ְ����t���7{�;;�|t�L�R��x�5���,r[�%91��*�"�&��彺����d��<�)� 
�@F��	H������2,tm�0%!�9�q�3vG6V�P�]��Y]��=����b�3�'�\��׈�k�,�[b[ǐoL��g��C����[�@=[�����2��}�^e�ݞ6s3�:�}f���A=c��s���;-��RtdDV�Y�I��~9U��R�z�����x||e��;P��Q8����~��Rf�m
^$��?����#-1֪�1��A#6�l��^��)��F��=��Jzv
cKהt�{���gU���ϫ���}�B!$Lƈ8��k�) �T�_E�`���'��۪ۙ� pݙ�,,�9�|Fܹ��.�="�ڥ���U^�>f���<=ό�8J���ìha�����e��?"�X7��$5	��5iH�>Ed]E�'n��3
��p^�J3�|`Ҭ��Z�)��!7뭝�fK�:�HC�,t!9�{��VJ+kf�����OL6�EB"8t�F� �����י�.�8�aЃ��7e��4���fk$+ZCΥ�K���u�%���@�*kE>b��0�)Ȍ�ӽ&s�շ���:\psV�q|�����(�s:I0j�RS��ۚI�{���R���?��M459�lB��`�����/�u�hA���/�Jq!�g��4FVu��z�{w �Ԅ4I�ӧb��@8��ic�����H/iqD�Ok���I�**5�QkL�ױ�&��t�u:I�۵�Oŉ�H���Dx��؆�n(��������kEˑ31�Ә�53Wԧ&������{A����7�j��ޫ
:�YB���-������0wl�o�BK�w���կ>��h@fV��ĸАfu�޻&R�|�Z�%�ʲG�Πn���ص��k��}m�2��CK>��z䩑e�&8����9�oS��B`�-i�,n��.l�����՚)��ɷ���k��}��]c���w���p�S����L�rj�;(��'�t������N��Y˒��$E�W�3X�n.��Tr��+3u	9bn����K��J���dح�";��n���zv����� �1��2q*�i#s����{�XbG.�M�+�N�ǫcVJT+Y�[�t�]Y/���&�(F����Չ��9���45�@[�ui:��\
��!����ݶ.�i���Y��kk<QŷgȯZa�]�S-�`k�³.t�΍}���/u6�n�\�d�.5w^�l&[�+�`���(���{���묃G��(���e�h��� ����E9���0[,�Z ��r�򑡎��\�PX������[�T���Z{�N+�fZ��ppe·K!ڽ��R�`�aP�km�zj����� �dbk]��!��91�F<:�p����Q6�TS��{a��`��1��-nį���N��J�uj�<4b�:}#��wb���XEޭÇ{O���j�g4�Q�\�GUJ���m�f�ce��n�b.��-�ݹmT͔(��IΏ6"ї4[�4S��,�R��k#�I��ȸ���1�NI#rwV.�ز��xB�1Wol� 6�2v�-.���k_f�Q+��fA1�Ե�)JV�Ƹ��k�
��ب��ѧv�TU�uq�z�cn%q1�)m�c-n��լ��V�ee�7.K,�]Z��p�j[]6G.�Fdn\S-kQk%-T�����ĳ�\0��ڔ�Z[h%Kӎf�ծ4VZ-EKm��Rް�^�Y�j-��([� �KA�nX��Z�ֈ�V���&(�n\T�J,�C32b3!D��YPR�����5���T�4�Mam�ܪj�(�9�[jZP�M�Z+�^��v�k�}��/����q��d�C�=
�%��n*�m0����u��f��G∧l�9���0R��u�ܭ�h�^�c��8|��h�E$�Z����3Z�c��K�*�^#fr,x1�(]7�j��$#�i�6�웹��b�$U����_A�.5/�sޜ`���8X��ݻǄ��\FT˰��Me	��B1@�Q��g�6;sq�|O��IY�/�4^�8�5�2��FS�Mpư��LT�P p�����7�sM���zq��=+�^��2�{�$>�jH����^�"�#���9S��f|o��۬L�aJ�'��j��=)����Xe�z��{/|�F��c��'�63�.�G�Ѵ<S�!�~���˕!>�����^ ^0�/u�E3y���'��
ڊ�o��Ӷ�h�$�Q>�~H�_um��Zy�� ���t����Wq�~��tgv���Äiء�!;�7��S�+T���=�ц�ԕW}�q����
>!vn�[��6��Ӑš�S��5K�H���:i�-%���c�_>*��#Ϝ�g�W������K�C���#W��Li�&&�;���,ա�_:��Gj�x�dQ:���ŀ�/b&�ݻ�G��S|��w��XEw;8
6p���z��}����W:���O�V\u�i��� �TT�3�gS�w���l� ��'��
Z|j�ː�*k����z���4�D��A\��Ķ<~UA</ˏ�[3JǕ�u�֟#�F&����&6"�d��u̍ѻG�n��Uu�;��bX������k䋬9g<�qC�kٽm(Ş{4MXl���͂�Z�#����3���y��v9[u!�ӟϾ���-�4���?��Z���δ���2#����ޣ����B-�A�
bg���N�p�'�5��j'=r����p��9�%�!�Ǘ�O͍<x�!������ھ�CJ8l�&a�zS��y���<A�lm�����k���M�km����ݽφ�k�/Ѵoa]�9L�D��vFF��[���9�]�^�ڮ�n�F��GL���l��%�Pz��Ƶ,۽���p�û|g��P��F�0���c^�
�w^�v�Zx:@�O.5�u�_�(�)�e$H;B3/��,l�j�;DW+5~��A��u��.|,B�;"��3�Mv���Y��.��8�7fwx��69� %ɏzQA�B�=gV��O�W<H��9�ԏ�W�Wǻs���_��:ٳ�<|z-;�Ɨ�{#&�����Uo�te>��C�S�$*��(/='V�Jxoi���^���u��}��DՇN#2����p��
oM��Q֎���4.���ǈ�p���?;CC<p�����ݩ<�ј�ж?k�P>c�3g���R�����{[:ǲ�Q�ÚЧl��F��KC�D>�cF�W{�B�Y�_!�������!K����'�^�yΤ4�':��Tf�)�˳1s�b��S6��� w��gaӨ������
�'uR&�������N�Y�g^�K�s����/n���%�'�*Y)�����C��^OQ����Y����p�-c�K"]d;۱�e�΅4풢'qAf_L��kfKe�b��4xnŮQ���諭��Q�>N�ä3��<p�O���(�P���$�aEiFb���e��vEF�z�8��}:u�uRb�n� a�MmY������dW�B�v�c�q}��u�y��5��ӣ>(�;��������C�ާ&x�z������y]0�T��!��<_�
�ɡ�N�ӧ.���k�~����R��l��gM�6������ Ջ��t��f�6��#$F�WI�=1��La���:v[\ r��J
^/��F�������8�$��V�\�zev�r��C؉֬���(L��L�^�W[{I}|�k�
����z�D��k�q�Qˌߜu�����Z��Wr)�7
�r7�c��pu��S�������,��)�A̙�C ��+��9!�a� �Ԩ9Fc���������e�livV���68��K�j�������A�i���v�}AQ�2���s� i1���:��1���p���x�&�>s�N"t��<s��gOKl��X����!�N���B����g�w�	�=>�6��W2K�Ǵ���`�0��G��Š��8j��^��z˹��.Z�������R�2�/E0:�j���zR{}����>�a��ט- BΚ|t����?�<n���������x`姪�+�5bP$0����²�2��y�i��q�u��Wl� �H�����k���l7;=�q�6�X?Y�/{�<�x�^�(��t�	�Xl�?.�߽�x�Z�����`��.M'�m,[y�TF�]jE����	b�\��w�Т�se\w;a�t"N����)�������UW�S8F�n�$k�`/�����R�B����a�5N���*���gN�ðy�|x�Xa��x<�N���y9��\�r��ي�A�A�d閅y|�5�Ǎ��M�}z����(�ŇO�!�A��H�Y��`ƫ�1�+��mz�GNȕ0��D���&���#���*�6��y2�LOg0��.�X��G�4t���}���{�w�B��!����"!e�ZC�.HiGt{؝̩wՄ#��1�ϏNye\��ޣ"��à�p�%}<[�w[�X>�c���D"yi��]:=<��D̮y������C�2}�x��칄D�"yl�2����ǆ3�̒� ��;8pܬ�,�v�b3sa�R�4�gs�:�Z9�n#�t�tŀ���f��*g���r�2��#��� "{�������ǵC�����}d�-+�z��w�}��k����Lsb�i�c�5 �"�0�iq�^����99�K�.&�9������Dq��q�g�.\�����e#8���EZ�s3S�L���H�m(��PO2z���XX9���~��ʥ����m�#��l'��tM{�Hg��uSXRںq�o�C,$秏���YD�չ$.�:�K֝��O�OβOG����f�1�찯+N�59��DL���S�P�^*m?��%E v�<oVn�cB�&�'t���*�R��͌�z+�[�6T΂��jD6f�yy4(�>���+`a[]6DÓ�}_U��)q��_И�����Qhф]���;)�x4��p^ʏ�P��'�^�̞�_A��z�/R����0y+U�����Q��+=Ө��t��ü�@�sXı�c��	��{C�1�ϖ׮���P彧ބ�}2Oj�Z�>���mx�8��bq�[&�j��pǾg��"K����v�M�^2"�+M��}F(���p�}��c-{ki���M\%�'8��gعq��f�3y�v=.�ryy�?n�(���u_�)V9���x�e�ҫv���2�ƶC-��*�w�kVѐ��wJ�gS��l��h����pH�=����oվ�	����;��ZKF$ֺ.�r������n8��cu2v%�j�+u���ݩ��"��m�.K���;x�)�^�ؒ��p��f��Jpc�pP���1��:�K�Rk���M_��sOnOmS��|���,�M��dt�Q���%s�ل�|�7WK!�l(�}�F�g{�DYHeo���C[�W�
���K͜�ԃo�Te���g!�|!�su_�{��5�O5j�����Ȩ`���MD�QحB.��m�S�R��kwi|�>��_uM�{};�r�O"�5�����/��G�أ7d�˫G�F���OV*��8��kv��4%`�ӝVh�S�"ڥoz.�%yy��(]�=�uQ��x�M1� 5�N%���=X��znh�z��2m���~���B�*��+�/�Ub|�U�9�3���4�uTҌ��D�լάJI��V�,u�|�8� �]@�+�:�ڙ�e�
@��qv���5�ܫ��Q!3�)pn1U����iZ���ј��6V
s"�pymz��0��,���[\z��̖[��;F�p���L;�m*N̵��\�;!��7m�t��hҷf>�|ma��e��ìڜOn=�f��JpP��$O4U�� �"��m��*ߣ�ͺ:�u;7~3�I=9e�=88�G�h\��U�kk,r�C���m�|�vP��mSuv9�4��t v���]o�e��2䠖
�84Hج�&-�c�ȱ��f�D���7���o)�L����� In�u姴\ކ+�l>6l�feք�B��-���BX��8�0Z�Y�5�+��n��=|�ps��kږ�6~�z���wKk5���9Z��!�
�R5��T��U�b���bb�����/��ފ���*QSQ.�4"�[tV����t��:#}gx�"��io	GD��x��s(E�S�3$���(#�j�3%�z���3H�N19$�͝j�&~���9Ԏ��ɱ�5-0^�4%v'{�=��7�TX��Y�
�KT���������c]�b��efQ�ƍ�[X���U�EYYR���ujj�QQbi�M �]`Q�QE���U�&$�ѵm�YZ=0�.�r��A�D���b`��˂#m�iQPX�F�mF6ю5`,�4¢�E�Z�%chA���[+R�DA��*,���P颫N������DT�
9IP�
+&�Qc��-Jֳ6��`�PFE��d�,ښIUum�b��\����L��#mPU�c��MR��E�a�}��´v�2M#K��[��K1q�N˖�QnT0܈�RO
�fC��>�f���1gx^� z`G���R��4�7݋�E�B�]w����/:�x����D֋�ד���8��+uw���c]�;B&�I,�S��pZ!��_Y�-1��#~�W����$�eiW����ہ����ؽK�;u�K�FI���Vu�i8�hɋ�CIQ��U��f���s)&K��}�����u�g�/ae���L)�T:�y�ߕ7��LZ�:�~D���Q�%hF�=���B.�B�'8�y�����:��R�c csҥK�{�U�39�ZrG��oe�QL�y|�Q��-�Wpo��]��<�Ar��1O8�]�E��uw\)�v�i��:1�R���{t�Ude\&�Z;=T�e����fU�+��ȸ�xb��Q�ۨ��f�x��F�{V�v���{Ů�/x�(Q��G�zG
=�v{cV���Oy�w�S���W��Zt1c^�>Q3��^�c`=w�Z�ܾ�o�=���t���]��n�d��{�r⻴9yg~���B�W�.��L晸�j'�H�V����hY����}����[P��{�hO�����y#f��
�
�;�Q>[M�Φb�ݽ���Kvkd9�BI�(���<p��ӽi����7F�%��Cŕ�O�_W��F�Vti(��Ғ;�#`���˛�2Lë���ӭq[3�l��9M�Y]�WUٷcoIN���ŰأiE��V��MO�v�v&���9_���ep���P�]C�0���r=5�5@��^�;J���˥Ѝ���KU�͇
�,�#H��������Z�}ɗ��^ �a�D�s5e��������	�a��E��撯Δ���`��,��ɻ��MϢ�����9��vu��)JV�F�b���\�����8dP�f��r�J1�iԵ�k:�aJy�a���i){���Xp׾��лd�,��~9>���[Ya>�B�՜Ǭ�Yn�O6��V[�z���B�!nK��R�YU|�p�c�Y�!��˝��T�Ɂ^���N~\]��hE�&�7�����.+�^y��]g�؛\�������H�A�Ӡ�㜉�)gzg_�=����v�q$�lЌ1���l"�rI�A�k{��:�.�����ψ�Q&xӔ;z�G�W�K^�Y��������Ԅ6�y�V��*^tFЛb�6a�O���8��4]����M'���]��
wWIW	O3(��5�r�aE���,������a�oۑ�&��r ���׻w����E5V��G�
]��<����v��o,;��1��W;3E�T��l��KC�S%�ǮT��ީo����ɝ�f���<�>+�/��a||��s.�e�F{�M�8��9^8C5���v���|q���tS�XY�����<�i�����e��`��6or)v�i_i��Th�#��g-�7�yI�+�	M�;�s�����E�LI�-G�I�{sv��kː/C.we�L�Ҟ�Rp6�vY"�b���1Ö�LAʀ&�p��
z�}�U.��F���Lp}X���r��ܪ��x!HhP�Z��Ѣ��t�?���T��ht�}2�.֣�n���40�x��wu��PF�Z�iQ���z�dC����A�s(�ɔ�,H�>�V7)t��N�v�h�֪(���R|�B��i��v����]�V=MT2�"�]���(<�Ȣ��q�Y��s�Wq�zs9ū�q^7PU��h�noUC̭&0ɳZ��ֲ������7�U���O�>���p��`�ㆻt�u��]g�
�.Kd�N���V�̩���pC���ٷ�F���e����k�ʳ��"�Z�����i�T��N�K5Pل
e&��2z:�y��,�݀LX0��|�;}��a�����K2ы���ٿ{�>C�F�\��5Z�Z�d\�F\S5'*�hF�7�>� Րz�0�v��Mg,N#^`o灌��%�lR�5��Ȝ�%ͱ0)D�Z��#�T�/�1�7��78�Aa[�������9<B���n�Sb�s��7\f�v�l��u��^=�/94�F�MU�~�6��l�[��k:5�[�EB��w}�Y8��W�D�3�$8���u]A�F���Ɏ���>�z1�S��n�2#Pt���;X*z�]Ԇ�9���ut�m�+:4�Vӕ�zr{X�i�׮h��z�ﳆ�d,Fg����{�\Z����.�F���v��6��&[�o�#X��;�\)V����j6�L�H���R���d�k�u,�Ҷ��쁎�6�\l�1C����z��}�̹��<B���XH�|k��Z��p��嘵[��PF��qAMh�v�Ps%���Kyܸ���C��\�����WP l�u��f�R���X	���m�6Y�LTX�OFB���5��a�>�����:�ڬ�h���re�\�[A ��F1����e�nq�:�˘^�y���0b�a����
�f]nor���C2W��Ʌh�Kz�1��|B��k�!�]AF���mn�ӡ��q�V��q�0�j�vx�{�Y�
tUKTd[�aꋴ�z5�Tĺy�<�_oc��N�uz�:��u�����ϸCW��٧g���4���q&Ͻ�s�G���RDz��L���`�QX#��q�jP�^���V���K�b^���`���BC����'n��ٕ��������E�FF4[wH�z3Q���Z����01�5MTf���-q1�J��V�Ǟox�ŵD?f
��X`��qÈ� �x���HR7Yս�����u�N�,���o��u����'Ľ��S��D\%u�[l������%���]*����[�8��˕�&�"Ȅ�`�Mq��$"��-���et�vzڇd�4K1.�;Ɍ5wh����<����#���b��~��Nk��̼��,���ﻷQ�8H�2֎��MU�򺎑ctEʪ�ZT�*�e		�d9�N��g�
��~���1ND�*08�U6��d�)5Uּ�%ɽD�[�����bj7rMOjQ,�I�&[)��/�9�ӫ���d��l�����q|yLUQ�{�E�B�К5:��T#�:��Ue���(�(hS��ҋ���2�7�q�}������x-e����<=�˥&�Ke�=P��^;�4*�=>T�*=��D�J�1�7.,��t���`h�Q<o*����%�6N&���V�O�����7�TY
�a+O%\l�z�����*�1���'�<����J2�����8��clPs��-���HzV��m�Oz�w+�Fmn�9mkL[竃w&k�t,,����8-W��+(p�4m��[�.�l���$�{z��yf�ѫn'ʖ8&���c�\��X[�'r˦Bn��n��Ytސ���`�F�>y�x5�鴹h�Fn4����U7�{,܌W�5;s�@��K78D�gz^�ѻ�F�\v�ѫ�"�n���s�.�s����+n���h��4�!D�p���݋�3d���X�f�n_u�#l˱Ӝ6tA��2�uL!/{hr|9Lꗽ+���^2r]��ۗ}��&�9�*��J�<��ˈ���Npmv�K9h�2��R�apٓ6e�8;MXܱ�d��pq��@"�8\�6�dثG��C�
7��n�<�� ��J��������@?IX�Ԭ�Z���ciR�Y%��4�,��f-����UX*�CI\`T�%L-��-R�L�2�uJ1+
�Q4�dX�� �cY�Z ��EPXiz�iTTAX��ȺJ��PQa1�dQ�b� �&P��*�
�X���+J�FV�T\I�QPUQb�(,"������WL�C��,PQ�T�)m�$XVQ�]y~�מu����j��F��6:�b����7(�IS�S]^��2�e�JE��l&���=�!�Ӟkx�ȗ{�[�
�$�_��c�Ms"�kE�{x��:�1�3\�ρҷk�^��)D4:��f�o*����-�Cټ�q�S���zv�c�W����iFo(����X�5I��v�h�גnT�)��u����Bǳ��θ�\^����7G�f����
[ĳ\9��jY���~4��+1	S��*t���Tt�!�W���6f��1��M���Ų�wU�ر��~��=�Kĝx�IW�+�B>5n@v��v7�e:�$Ih�����F:�H�f���F���5W�Q��g�-K�� n+
n�Ù!���Q̠���b�`���+���|l�^ޣ⟊sO
��׿5�-g�?daH��C16�F�o���;L�-$�*ڨ U*�z�ΕG!�Dot̮��ʐD�C_���Ql�q�^R�-d=����,D���
��YׄU��z]�3-0=�z��Pޣ[�{�6��@:.�ɶO1���?G��5�o��f�Oٍ�N��M�}���G8 QT�C_imL�ט�ɩb��{[���%�D"-�����i�hx��s�ɫ{�K9&����"��rX�"�esi����~[W�y��یRP��V��O�i�_�t�ei/�NQ=�+�=�ꘑ)����	|���Y�z*'r�ʁ6C�Đ��t�뽧�%djg:�y}�u$��Uo�H�Q�s��L��g�{^�q6�q�^��5��F��|}��fX��r���:�sXD����$���Wq��F�cz�ސz�y�F EU�)�����C�m�K+�J�Es�2���-�q[���K��#&0�4pI���\Vόȗ9Z�䥍Ԕ�ܣL�v���suχ2�9^��-4�1�����o|�o8��s�DT�`(�{^���ڞ��.��]��&.��z���@B�bhw�{73�qQb�1�^�j�/�F��gd�k��s�g�	�3�<#߼x9�T��0����[bw��eh5�x�眂����1ȭ�/]���n�C#V���xa��ŷ�}S;q�s &Mn��eeŻ��GwK#��?^�X^�ͣ�S쾫��n'႕��i�Oˢt��G����Ef��t�47\��B����f�}���!Z����#�L�4���32ƹqb �-7���lڋ�INw7r��t���p�]���|�D����Q�-��/u/0�w\lw�fDK.n7��w�FS��"���w��:���-Se3�~w1y7��Bv�5����MW}��P�I��$ꣲ\#1���wlN���1��.�gT5�bx���T��|�C�K����B��q�F\�����׭�z��m�\���_k1�������ky�yܸ�	�!y��j7���T����5N�kʯ�����g��ë����n��]a���]-yQ��焣�k>��5Su�c.U����|�&���b�3�3u8Md��=��{�ڮr�>�:�C�k��y\��sG3	A&=\���^�E��jӱխi]g*y�1yx���y��7(���}��i~\��ʈOx�|��Zߚۘ,���֦G��\�^U�W��n�'��
�<s�����pbE�i��4�X�������k�������a�gw�Lك����q�'@_K�o.�}}���Q)��7��;y��+×R}�_w3���qk!�lußq�Af�{�����.��50�r�����@<{�Z×�gNA:�7���L���ফ;^��Ӣ�a��8�y#�
�/K|�]�<iM�h7Y�`$+{�a�@鳦XS���p�[�:ѧ��iW��������}�X���{�Wd�s�.'�r�>o�yom�v}Z�% ӊ"�Fyx��^-��ߢ��i�5��h��W���޲3�������o�	Dl�0��n�<7���`jź�w�Q��9*�D�C�|����)��vY�U�w����2�c ��:�x��������QA�Q>��6c���7�Rqq$fr[ ��a��DO��:e�ѝS�e��Y����UI�H��_()���({��t�e�{w}{�e�os�k7�9���)�[��S�K�rr�)0Bs�6Zcnz�{�W2zoB`��ލk�擹j�/ �;���tgl��֣d��Ҡ1N��0:,�]�N�g�#�g�����Zg�5}�	I�z���u�=y�y�Y�U8_�AѦ�9q4�r���ҫ��m��2,�wY�|=�;W�<Wo2�۲�뭜f�uq�����|ra,�홠�1�G��-���j{;v��UP�dY�Dj�3Y���WI��.��u�	���8t���J�oo��i�Э���h(���Z�$`M9[�\-Y�R\o��gA�T�Q� I,�lmE�2K&���ٽ?jk����d�<Յ���k���,I����f���R �t���^��˚Q�OSz/��&�T�c'�#fz&�D9��p�K2�7���a����*lX�����T�)V�G���>hGne{z��t�Åo©�nvw3Wl��"�����gg����u��ѽYb���V�ylzD�B���5�^�!O:���t犯b:�nhɊs�y�+&�
��2Lȝl�\�͉�����b.�O9�����M\�<��bu�s�����	R�|l�g��i��X��� ǯ�׵��C��e+������gL�궙%�u_q�Χ��|��<��OR�л�Q�GL���i��>�g_���P��վ���ˍ��+V��-��n7�c,�1�j>��>!�$g�x���'JGg�}s̎y��ו�V�.7��6JI���o�߆��Bc��Zs��S�6MK�e�z1uw��w�<gtc��rf������y�?;�}���lv�z���+D�.�n��8��7�����Ĭ�ǅ�[�������'A����i����b�Ư��:H�U��V���6i͘�l�{�+r��ؔzFl�;q��w��:�Lj�X5��A�;Cg���"�;�X�6�������`�G^�!tw����-�絡��zs5t=��6枛�#����<-/�N�+�tީ!��_�-f�J�&U�UWI����2���:�C���PWܮ��o�Bj��ĕ�SqT�>9}u6[���� ù8��	��ﯥ05�9�I��n�;}YA�6\ٽ�v��`�);�wz�CX���u�F7��r��u���ݬ`�WA�FZ{�+��G|e�/Q�8mnB����Ҫq���90ER�w��G*Ͳ��C{#��QI9��^��e��튄���-kI]�ɻQYZ�����6ɮ�X�冤K��;��f����]9�n4*ev����2W!��s7��(�&�,Z�Fu:�q}Uj�U��3FP��q�ǳw6.fT}����C��ϑ��ݪ�_fL�pt�q�Dд���Q�K�Y�{XEO�����u��E��t�4(���ӭ�L����n��ȋ�aR=G�~��<����h��iAwuʺI-�+sw���݈�����WNs�(a�6I����2����K�XH�yEL(.�U�K���Rf�X���չi �Z�N���.ܧr�&Vv��.y��f���W[#L"W��痲]'滏Y$Ȥ�ԍ��Ij�m�V@j姹����vv�	Ws��g%���EM�DUȌTV*�E�bȪ�!� �ȥk���TC��k ��#�X娨��t�,t��Q�"������cSC��4���eX"�&��Y'MN�P�\q�m"�X(��S3&0�H���b
(EZʘ�*��.����#E��*�VP:`%AV
(,QA�T"����X�J���(���AG�~h���xw���PKQ�f�"�)���hc�2����$��R)��^e��L�,�Վ#�g���D�ݜ,nn�o[�#�-P�4x|aa�)J"T.<�ެ�]6��5��q)��Յ.�����*�9���o5�:��o�yl�D��uL���B��[c��4ϻb��*��p���b���J~~�sA%�=��{*�=���nGvf2�p핈��G��G������:�&�]��7���gnV@F�dA�s��Y��b������=��\̷��v����,�7��5^"2$�ѷ���y=� OQw�yJU�㸺ɤuw������ŧ�u����к}�Y�H�-��f����<���M��Y��qq�N=z�m�Ov5�&�7�ȟ/lM7��ř�
�;�����õ^첸���5����&���!]�~/b*,�ď���$MI�������3T%��}PR8A�v��'�w.jH:�@4`�GE�j�OUvg^6�W�u=��Wtۺ��1��h��LF\�a3N���V'h����=�!��8k&&�E��w7�.7��w���3q�i]:@į�E�͓ٳ{1� 
Ef52�����ŕ�].�6���ڬ,����`r�h�����N��{�U���j��"�]�<qO1[a?W�q�D~�:"�����i ����eh5�Á�=i�pq7x�7�1��g��kϴ?3H��m��M�A���]�2��y��u����׽��dh��{��@9�������%�<��y�x�h���lƯY��\�y�y4�Ǻ�I�C���@wl�̄\�o|#eG'�t�0��\	����dن�N�\c��_
�*�W&j�n�62m��c�Ej�Q�z��zN�|���`�z*
�R�����[�\�`<L|�33eʀ(p�&fh�ջ馶��^q�/�6�t�\�y1�e�p���2pՍ�wn��D���%�at�`Gc�Tk�9AE���������T�lo�kH���N�=j�
�55�z��X��|)�w̢N�B�S!������3�5��<�xMߐ�W	����(��6+KҞ��'kϴ�][bl�?=.�d]�Po��:۹WX��T��:�n&�->*���Z��j�)^:��3^��u��Lv�gZ���{G$�k�^�O8i�@���Ꞩ���_�@S��#�JȮu��g'd	 �k;�nH�ͼ��n'͢w�{0�ڶ!^u��q�i>`��q0��R0�o���dB�ڹ�uť!�=���}-�6�FF_`��V�|�+|�s�p;�:^;�=˰�0�{y�'�yc��M�[χO5#ZP..9բag����:���-R��č�O�9�X3W`��{*�tհa^��V�\����=T��L"=كCX���y#�1����WM��`қ�*��#
�L]^[�
׽uY��(�]�rk�]�C;YղL��p����e�"^u%�,��o^6'CD#ׄmfj;��n�!-C�{�d����i�3ĸ���꺝�\+��0�㣙�>�8{�=�h��[�i*�@<'�'��0�~�QY�Bh{�o=Ɛ�?(-�Sc!>��so-��<��t$j��xO!�e�{s+�>�4'�xgB��L���յH�j�/��=S��eM6��5d���&�zۥ��o���N�v��w`F���z��[ ��OrIG@�TLiZI�]ځ�P8y�P���{��ޛ����{������k8*��;�2�`�Z�%kqE38�M�K<�z8/c��_����f6�ɼEF�vA\�����5�H��$���;�n*�y�F:,�=Um^!=hb�|�+�6I[�P���]U�7@U(�bu���dm(��+&,Tb7�V�u2��[~��~���:���T��X�7�o@��Qh1Ui#����Y��of뭳�
.AO�޽�F��W&��W	�%�[��
���!{|����p���k��N��w6)X}N)��|q^e�k��GTa����նtWM^6�-xEj��-dE�4w2�9���{s/G�a��v��D��/�dz�9a��dv4�
�Ƭ�bC���+%�&z�f9�y�q����g	��k����[Ì�k��e��� ݥz��+Y�B3��q��^+�r�Qn��CH��s�Zw�s0uFu��闙�����9YӴ�,n&雦WW�{+�Xi��gp&7խ)����9��|��<����N��S��h������%��7��b��7A1��X�h��"�ص�R�s���-F��X�����n�In����b�E���l��Z��'*��'�ܛ�"�ʉN�
=�ˍ� d��μ���oQ][�C�_��.�� +��6���
�6'��m����е6�:�O.@m8��$���k|8曍b���5]/:t��6K��M����������U�j�&^�^�lf���6e���r���HH�ֈ�0R�_u\ἶE�1�F�g9�2�lΚ`K���w�tD<V{H�Jj��\7D��z�������<ON�Z\��O^�n\�D��m����8��D6��fg-1s���r:����ʡ�O0�D�E�������{�)��p��L-�.OW�ڀ"p��=�w�AEM�#�ˁ�8L3�	r�fp�1}r�o�`�C�͛�G-�F���us��5�q̕{qƦ���:�P�aR��6_E��LݔO�>\�5[p�2�$�R�F����@�u=�{��rjݫ�/���h�ѕ��n/�MíwWבJ���.�r������fʶLq{]�V=;*���#�Z/�o�f'l�$�֞�Q%M�T���4�\���9p�)�=%��.�BkZ���Gvƚ�D���˷�����sq%�6����Jry_v�g�R��b�cD;cV_�G�����s��$��V��b���B@~�턑 <�Qd�Ia���*)S#�,��b�ey|�-VV��=�&95�&��! P� ��HHBH���f���'GQ^�
�š�JeH��#8��6ʘe-[�!�c��m[��ԉ�IU���j��+qՖ���l��f�Q�YJ^e&,NX(��J/�ƌ��4�;,g�y}��,�e5l��rg�,*�5�&x�03�	 ?�5���W��U��JI�v@��*L�@~P�U�����khڱ�����'�<V~�ni�����9�N�q�IVvyD���H���s��RR�6c"�g�R.�1v=�H�\�e��A��QZ��Y���o�"��_)%�qs���RQ�m���ȦR���'��BHH '��tY�I����c�:�D�$H#»0L$�QX�U!�$���&ՙ�-r�<�=3`���b~�^�H���FJ�URYő�ǋ{���{��-zT����Rbo=�f��N���?sc�����o��g�e�ٻ�*X@cޖ�����󑹓��;y���}T�e�˦�ZE���v����˧��X�	1'�v���q}�Ns/�����$H�RQZr��%y��SF�&�ԧ�,5���eKZF�I$��$��B}dSQX��'}ZUYWj{R��i�SF1bF�!挛�H�#!�zQURk�WE�Q�h��V`-&+I�f)#�����<�5�Z�Q��V����Vh��%"�L����R^��F���%ʯ��c(�$�s��w�9H�"@Vy��~�$�p��êR|�n���|Q�Mc�szpE��6��W��J.��ul;f�u��"_�:$a��4�>ϵi$K��C�p	U�Yd�R4���D����L���]�8|ƣ���N~�i�g.܏W�zўCE�R�O_;0T�%��{r�>>A��Sm��֣��t�m����f���wa�n�D�~��rFQ�lg˔U����F�z�,��Q��7쪎��(ڳ>���F(���#�dtQ*��*I�/<�Ǐj�GMy�7	������t���Rd�L���ɑ�2�,�IP�;��M�)��R�#�)�Y#���M�&s���"�(H2�4t 