BZh91AY&SY�qR_�py����߰����aV}�N�  �*��((t � @�   4��´0�*��vd�5�)	-��E�A�v�gg;[MQ�h�ȋwNͶ*��� �  XE�`�0@� >       >�      �v    �[c���w�ݭ�]���s{u�9ۃ�r�Ǖw�onn>�6����w���j
�E����4������x�۞琐��=}>M}i��es�v���8�Xy �ep>���`  ����2}����sZzn�ct6��|}��/��=iOy��h�n�
�8�����#n����@
+�)>���m]��Q�;����S=�
�����׫�!ېu44�w
��tn�8{`�[�(�` �|��y����ŝ��u�l�:{x��;�5;��m�������ɼ�r� �@��;m�dc�::��e�������{'��^n��;��U�vB� <E�� �^
�{��vv�wwh;�=���j.�s]�ܸۋq^���`�� �Q�{�twb�s����72ۭ��h�w�n����q\�r�]� r�z�  �V�+�ٰ��2�v���u.���w�C6��<r�0 w@��ٮZ��qIv07�5܌�9yyt��t뢕�H|�                 �JU(*             "�jz�)Hڍh��M0��F�L�HI*�d�`&C��h�	���QJ��0 &      *j� �)�SBb���OH� �j�Q�H�J�#ѥ3D�M~��4�= �4Ѡ*���J�F	�	�d�� ���o��\�[��NsW9��MB~'WAV�)���ITI�#�����%除��T �w�?�� @4�a���`������y�s�_��?�������|?���]>�\��/y����%l:M���a�6��_�\��*~�쨊��?!����d�������E�>������'�~_�?���1���@�\Ԗ���V��_���9�̥bƮ��j�6��+�B�B�S[˅b����_�_���[K-1Nz�b�Y!\)�J)@�T,�E�����m��)!?H�����bw�d�
%	��b��Z�I�k=~i��T�T%b�7��e���j=j�^-�,�M�D"y�G�6,�n1R�	��Pb�T�1X�(�Be�PS��^~'��V!�"ԣ�� ��V���3�\�b�Lp!_�!R*�Rh�&����i�Ȟq��8�(�!`��6�5~B�c�b����.<#��I�.D1�q��%��c���B[P��,1�����!4k�h�B�xB;�bhCV�
��E9B5���rD1
p!b<!��x�Ǎp!NˋP%F8�ŊU$*��h�T�G�Z=Z��@�B��!Y..)��
}֥BD1
o���ňW���B���H�!T�@�jU$S�(F��.G����.��S�z�v�)b1�;�m�!�t8;�w;�-Z�t�[r�
��>c�)E�@�^�R���D!�Tڔ"]��#^)�-�6J�l��!��2���{�ВH�G��E�B�\!r��s(B:�r�s����'m���x�	��Xݢ!b��Qy)G&���q�G6�n�G�n6��lD<V؎b�:D:R=P�P�5�y�6jS�Z6�r�m��?4sh�=׻��q��ԱkW�~W�^B��m!���^��c��Q����F�����X�/�fc���An �dF�#�����=I����������bQ�
q��'�sS�t�}om�s�v�7-�zs�y)���Sȗ�W�mʣI��x<[�FSy1۴ۅ�-�n<x��L�Β	�+�|���p�%s��R*Y
��'-D���D�p�o|jnИ���\,\,V�V�P��s(ZRy*�O9X'�L��i�Q*-(�LOP���O}��&�4�X��^�Ӫ�a�����R�Z����R����OڱJb�l	�
W=w	��$�5�߃���/�MYf�ۅ0ShW����;�sn֦chZ6�Mhۧ)��P�F�U��j��]#|��g��J��������bdc~�Λ��R(!6��.C��;�j��5�b�ҳ��G�b�n��b|�
#ܡ1w�	�\&��~)��B�
�P�)G�X�F��x�lU���j9�&b|4������6��K�Bx�U�Z&�i��(�-B���څ	�Q��t�2�2�Ҿ��#Dq�ھF��R��t�!Jb�`�)1
�N{%?
-�1J1�.O��Z�����DVx�F����y
�H�Q�X�X�P�ZP��#؅bŦ.�@��˔J�-bb�SL\���W�|�@��Ą%P&!f	�O��r�����'�Z��(R!b��"�
}"�HB�B�#�0�fDw1Q���uQ�8�=�
�O��'jQM?r!1\�&�.Bbg���D���MQ��kq!u����X'�����	���r�~�
lLLB=��,L�i����V���pb·R<*������j�[�5>Y�P�Z�T��)V؜!�!0�|ňX,Q��x�b�B=��6�^�U�D>X:P6��
Kb�k"؅B�C������`�M
[�iڍ��<�p�p��cjWz(�#"�Yi�	R=���'h\��#�dC�
y�(�)�l�P�jy�1`���ad&�d��Yb�\�Er���"&�^6!� �^�Z��*)9[	��NV���*&*9F�+V�.���Z�P�b�1R�[��q,Qd8W��a�2�&1Sv����!�����W�g���c˅Qٌ�mC�!ʵ�Ά,Q�HZD;R�b�B97(V:P��&�dC!*)G��D�1J�PعP�̆!�K!����!��"�Wd?؆)��t��#�bkGj#�LBݦ�P�b���R�6+B�p�\C�[Bh���~�t���M���v�-��Bӡ�!�V�	�$�(G�+D���%
���rD1���X�]>\�
�¤�b-�HR�b�'h�+T�(ED1
Q�B���Cb�U2�C�(T؄FC�!�nzTJ�DC��b�-lB���יI��Y�:z�f��k��"��b�!�b�HO֐�>b�!�&��r�8B�t���#\!�J%4�-K�F�؇j-ǋ�r��8X�+�H��#]�b�`C�!��X�ɴ)G1B>B �-l\�Hx�ة
1���Q%��E��R�,C�bZ-^��M�mG�	�$k�?R�z&؋e�f�1�o!�����K�S�"c�z�d��M�b�
�P,Vt<V��V�&؄��1�������?;~�6Tm#�G��s�=�{���z��l�"6UCu�DC6a�*��!ݦ��eT6��fl;�wC����+n�+N��������}����aɰ�.Q��C�M���ɆmC���v���t��*-���Csq��޻]�Ç��L
,U�����vZ�ᔐ��EZ�i�̻T�uO�N���c�k9����>�{6+��_��㘢i��sq[�T��M��-G3�י�US���*��T9F3Y{]㠇P��:W.��0���3��ob����z��fҎ9Ţ��s�y�!�;d8W,Y��1f���oƱGL8���x[����2a��v�3^����C�z�e��\C݆��ɴ�����L��L2���3Y�i���.��Ҹr6�e@����b�B�zK�R���h�q�ؚ��\�b���<!NK��!L�yǅp�R��P�� ��E1	��B���Q�]��Z��1
�p)�P���x�������t��N8V��B���F8�)(El9Q,B��h�T�<�Z'\zQ�q�T�b��!q�9J��H�!B-�1Q�B��ňW���B���
Q�B�s�E�P�LB�k����)\�
��5��T�T���b��"�V��ն8�xGC��·��^����h�q
|#��#�Z�`�j���i�%ڔ�)�+s�+��8�Ji$<x=�zJ��e>�B}�*!
��y�!�qjU�Gs�]�Wp�:r�SB�0B�w�ة
�p.ZS�Z�ȁO���jgL@�koV�ڬm�[b!��s�\�	�C��"�F�>F�@�l��h�G;�,��m��n�;�B�{����+�,TЭ�cY��C����1�c������~�sڍ���|�3Eۈ-����S�\Y�(�&�r����	q����&�X�9�n�O-��s9޻k�lU.%��P̈́��ri�N_�����h�w����sz�O2��*�.�������r������NS2��_䢿����;���~��ौ�H2d��[��	K��R��
=زκ�]j֍Y�����E���a	�BX��}���춱Mǵ�xD�$��$�l(��L�wY75=X��PNO�7�+{,���v��u/��N�\F��Ak�jv"I}#|�}~����OS��'?X���V󱦶,:�|��g���U��8���PB�d[���n���U�rx�ۇ�}�rvb�.+F�5��G�P�?j>�/F�vNĽ�%���~���潧G�3��=�C~��]����38���r�"S�w�g��G+���:w�y��g�ʎ����C��j�����fo_�]���l��&�{�[�oe$�����,�!�*a(ۅ0��^��s�U5�z�T�yTl�<��� �xߩ�inL��3sW�w�ڵ����d帶����]����~��t�>�~���Uλ�ޓl�H�vGg������"ʌ�o^$Z~�~ڝOv���>Q'�ǒr����d�ST����)��M9�Vު(����My��?~�|�E��2̍��[�Q$j�Sq�i�S�&��<Y�Uf~��ZtN�ġ=	�U���~�G�����hI�Ӻ�����ȁ�����LGpW(��\�̗���z�<z���#���u�y�����3�����^l�Ǖ>�E�����3��4�1�V��T�(>��˯��-��WB݁�W���t���9v�2���Ӹ�����]�t�6�7[���/uDbɷ�����[�v�t���O#ޮ���2��9h���������Y*>~���oG9c�>S�+�Wt�c����5.����3ї̻��Y�Ud�¤��E��W��Mj�UI4���v�<m�Q���Qv�R:z�<�\�d���=!���s�MMK�wo#�?�D�j���棨#�jJ$��T��w��..�/*�i�%�p��ë�-Gd�m���So��<r��8���)�5��ӆ�w
�U�m�����q��]IqyE�������a�SQD�n-��#�{�ջ�7����><�p~D&�H!�#�.�A��l��:C�3���
�!V3�HD�1�	�vT��r�4�'r���?<J��s>YVE��1fu/�{̮�q�z�ꉍ��簴�s��K]�Pc��^ѹ`{t�>�WQV�ƾYQ�<7�'�|��c��b=<I��G�_�*ʱ!���i��&Yt6=�%q��kɜC��z973Q��ap�^dX�������Ժ���	�����E9
�Rr>��uL�{�������M�a3n������s
��̬�cp�r=�u��u�{��Gj'?�\E�<$�§Q��ՠŃ���� }�qJy��Un�nna�zK�������:���!�uf�=<McU�d��;櫛��W	*�k�lob6KK�ƫ��h�őobفRE\F=���#J0N��|��Þd�5F�cj2�'|0��,�dY��yp�*;�b����YD>�61UgQ����x��#6�}*�0Iٽ���5L��Ҋ���;k+�N$�յ�^�u;��$Q��˫�{Yγz����yg�E�FǝY�z��;��F����4[J�,�d�	Z������|�C�Ou��}Gߩ��=���i.=���e��\Y��{_-��YW�׋�J�vWһ(��q5�����̱�폟#&�n}��o��Sv��s��
���k{�t:��=r��x�S���Pd���K������}5>��}��L�~����d�#=��8��sG�\d"[��*F����5���K۩\����W���]Y��!5b:��ĳ��#c�k}G{Қo����̺�2�l�Չ`%�rR��y^���-[���5+q��7^�,ϧ8��ޏ7��se9��ϩ��9����qյ�n:���f|��:C���.i��J��B��a��/椩($=��+���9d��[�Ϩ�o��ۥ����E�H�_��a:������,���U${����r~�=X��z����췺;����=�<���K<�D��+�*\X����_(�����s��J����[��j�Ƴ��\�ϟ�v��ɬ���,�eXm+�{��Y���roX��B�9K��GP���CTV�p��1�9b��w$�����zT�bԐaD�nB�O�ռ����˭c\��\��6Jeb�J�Q������#*NJ�����v��2T�%�&��%��/�ti5�%�S���|O���ά��$��ŉw��Zs�h�����I��$n5ʋy+�qĸ��u&�gn�=i�+����W%vV�qJ���)�vükR�PʸrڹV�z� �6���F�M�r��{��ݓ�����wz,�騇��=��UG0�S��Jj:�H���s�j2��duY�f��>pwK��x?A��,�89��Y�uL�'G՟�y�j9�QygeQ�oJ�Cb�Ԯ��9)аۼ!�Y����F�Pϸ[���4���C4����ZM{E�%vK5c��^��|�ŋ/`X�ǀ�=�۾Y�p�G�^��Lơ�p�[��<K;ەeXE�	bLYX��D���mbŚ�]e�rdBֵ+r�*J�%�n�b���Za��V��db��te�9�j���?��M��kP��M�v?@gG��ze���6g=3�����X[�}Vn�dH��H=Y�,��q�qcY4_<��g�aϷ���O������8kqo6w{6��&�Oc�WaX��{G�%;Q�~Y����(q��G�����N��3z�y�FT6�h�I�.�8����ݤ���K,d&Z_R����G���s��ӆ������,���h���/��h��|��N�^��^1���:Q�#�Z����k�s�ۮٲ��\�}����-y�k����E���H�6�q��*��;PSq,��),c�"/�<��<H�����y�kEjB�C5r��u*񪞀֡�%�8��#!.�6���}��F῾3��C���L�J�<4�d�C�G�rɛjJ>�}����k��&���Z�W��K8���q�����X��h���5�:�i�7�{�>�y+%0z��tw$/x~���H����U�����]����'��wH��*J�,���ֵ!�&ԞF�F{�\xU�Y���n�/r��N$;���-:���F.su3��1#����ؚsl�g�y%��]�o��cY���ɞ��/r���j�7q�����+������+��5y3D���!�x����R��x�՟����W�[_�#�������e�')̹g'k��6����7���Ħ��y�nmd򎝪�Os�7�|�l��z�`�˧('"8�P�(�%K�؜��Cڸ{l:+���2�9s�7��dw����uw_w��V�蜊lz������ox[�{��s|H�q>���G{l罺n���c�3�����ֵR�s�~�c���V�՝d��[ͫO�W�_�����珶+�}�NV���i?��G�y�2C�z�U��|�뢝�#�{��j��p�u��}U*g��<�n!�N>�n�NT�5\˹N��M���������ͻ�~�^��5����^_n���o���%'��4�:\�o5�+�G<j]���-�}��ot��
ޝ��T�:$���'w�rݚ{jU�j0��ʇ�d�^��^�';�N��Q�5l+M���q��7�:��&�y���ԆL\���uM���\8�	&����_g_V�⽚���p�5;�FUu�q{IÉ��N���_���7����:�s��[�޽���v�d_F\G�2�oq�n㹮����Ѿ�t�\��'d�ԕ���3U�d�3��9x�h�jnC��В�!�b��S�����z�M7���e��Y�`�eB�q�q:�c�	T��*�$d�m�LJQ��	U$b�����]Ia�	`דZ�����[cv��[ND<CMU(�j6d�1#"İHi�������Hj�Z�Ul�i6�lp�B	!��J$.,i|�,׍gj�Y�J#lN��V��EP�J����ź�\�Y�IQ#�Zc�)ȳu���D
��i.-JA��B��8Q��V26�=�p�f�$�k9׺�,a��R�	HQ�ڤ1+q�����P��YPH�ID�+BI�	E+��vLb2��Un!")5� �A�=V���	�b���DZ�숑���؋q�v՚�{����8�i��-bM������lYr?�ő��#���VBJ�ǣkl�<��Y/�+��)8A��L%v�j*� oKx.T��"�"x�p��e��I��$�Ӯd%ɐbYH<peQ%��y�=y��$}�KQ�8�"Vv>��$6mi�d�>N���i(�q�홍!_&���n�eu'h�{d�m&-�"Xrו\G4ٛ��qĶ��q-�P��W+K$��7TG�,U�ڋ�f�j�tݵ�*"�Ԅ��Q�$�FI&D4&��Y���׹נ��n8��"�Y��H5FŹU�D��܄�$�-IEYm���*�֨�謉�	Ke�奤�o�Z$��-rcr����2f�PD:��U�ج��*�'SDM$��0�i��+
}eHJ�!,m����k���<��I�I`4}D�kI�>3����"0��3qD5���~�a����Ū�0���g��֕q 
I��f�FǕyfE���ʝo�7y�U'W�Z*��5EnB��7�z�έP��LAX)Y�ڒ ���n B�w �C|��w$K��'��@���]�*%�V�)!��73Ԩ��b��Tr�Z"jN�djz!�� �:������U�ں$P�����+9��Y�/^{�rۨ}�D��S� ����j`�Fr���k�S{��X��?��Vk��(("w��О�~6(?����$?��������}��k��Fϕ���E3��>߷���7�?��!�    p�  p�  @ �$@� p�  @  B  4  ,P �  � h@ X  X@�  h�  ��C @  �@  ���~m[^��G��i��yMm�XK��ղ�ը�a��6�3VPd"2Qj��b��\��,�y��     0  �  8`  X H `0  �    0 0	 � �`  Ѐ �  h@ �H ` �  ��P� X X �P � �	  �/��I��BP�~I����j��ۅ�rf�͔h���n\�m��-��6YcV���Cj�"�P
�1���e���3��z�@  �  �@     � �P� ��  �`    X H `�  � 0 � p��( ��� 4@ �4  B  4  B �+��{��:QE��ȀȤH�TۓVn[�jfV��&���Y��ֶ�M���TrI4�
 �I6��m���~�� � �
�  ` P`  � �  `  `�
 ,@ �  ` @  �@   A  ` P`� 8@D@   `     � �ʡ[y�$��z�)c�q�5�Z��H�$J�� ��.^06�
���r6���)O3�X�[c�lScc�97&��u2���:�1NL�)���'-�)�����6܊j��l�?G���7��m�h��������g<z~���no�}��8}�����_�6��-�����ȤDDq�ڐ��"#h��Dymi�!R�!N��2�(�#(��6�:�#μ�:��<��DG�qR"0��""<���H�h�"6��")�Fі�m�Q�<B)�yDDIU�!mG�De�muii�aF�J��R��6Ra�S��:�6�#�[R�Dm�G��F�m��!B_�7����������~�iH��D��uZ�2ڒd[*�ԛ��QVƕB�V�2�5(ȑl��厲ơe��DFʡ�<u8�+�[��)p��m[TTq!�Q��^B�CD��V1Y-���*,NJ�)�Q:�I"29,�(L��m�24�Pe�1�+���J�UF��k�K��ؒ��GE��J(@r"?�mFN؉Q�14��YSwbM�"�IR�7v��E$OrJ:���p�l���G�A�F��qڱ��&�
�v�X�YEIR�bO
�ؤ�
�5Q:�,�ĨǒB"�%p�إC��
���D��f<B�C���+��ml#Ev2̄m�+����P�d%$�em�KP�tq��!ז�M!�T%l�#���dR��Yj�,��)J[r�0�U��2QFLC�AY(�ڬx�Q�+���6&4�q5TUܢ��R6�$%-�eB�m5B�DQn�4��ܙ́��1
5$b�SDs ��*Q����2���)z�ۢ�XA8'
+��ڌ�":()Kpb�N� �$�b ;m�-�E�����Qj�E"��2�64�XTZ���!T�Q�bCd����"��X�(�A1	b%�kYl���Uҗ �ȓ��*�:��D!�T �(�"�3t�#Diar�1�Q�d�dth���R��c(���h[�e2Fƣe�:51�ʯ6�F��l�2�NGcHDEr�F����"
���kv��2�\��Д�@�HYmE�l��� �nb�",�R���FJ+�P��TL�B)),$��c#X\�6B)���&[H�E�b�
Z�Ҥ$�Yp���㨨�(�L�!!G"���E�5	aHvB�ő��Ʒe�ZZ�DX�!��;KX�%E����حM�D�5�"Ne�i(�.ѵq�z��'�*V5Q\ �-v��D��ceޛ���C��r��ATJ��!e�Et�W(�Bt�pB*�Y��<bGQ11���$�I c�lt-$$+#T!P�,HI��܈�
�����I�*n���E"����\�����S,E�'�Ĳe�V�aJ!A��G��c�:QU�bJ�����,lp&
0ı�n�Z2Q ,��G
��B����V�8	c�
�T�E��,l�����F�|P�ƙk>��=Be��e��Q�:\���x�x�A��7�H�֥i��-�'1
����4&�J1H�\�s"nZ��M���Ec�P�\��R��荦�[VYeH;�AF<d����L<b�q5�)@�[K���F!�pH��ah�G��M�h1@�B9F�q'�d�j��1��",D+�RG2d�,C �!e�RA�R�eEMwe��ѐl��M.�葨V�HI�Zw�.l3LC����:�%��B��dq���jKdh���J5����.&H�ň���i$WqX�Bhq��rX�(�r��6FZ�r4�v�liB���:���-Ȋ��+,H��T�5��뒹$U�X7Z��D�j�ڢMc�J�V?����j�W �Z���N�(�Ҫ����]K6���T	忶�Ťġ��Z�F�I4+d�mQ�+S�cx�96̲��������v=�u�&����Nؒ�X�u�\��eVdE��5�$�#N	ب�,��X�M�Z�$NH�U\Yeǖ
2(B�+N�Ȫtm9+�J%e�Wk,M��N�
�����PV�*vWQY%�C#j��G"r(�IP�:�&X�c��U��J��%U�"V��+Cq	&��u8�		�REm ���j�-�+QH�X�Ʊ�F5!-E� Q�*�IF4���E��.�ܴO,R%lybu��v��Ҳ�8�mGD�?n�٤��[UL��ȥM��q��NBW]�v̍5|7��!�(Y%u��U"%�bJ(�hqB�V��,�D�&*2:T�m1�쑨�)K(�,$�;S�AEXB!)Rx��.	h�ؚ���162�L�v7T�Ci�������F��V�F����C�
���ҖWjq�^'#*EO#m����jTrj��8�Nڋ,�%J9/wMi�L5	���h�E,��A�ԝ����i��I�
�䲫]c(�ov���[2a��e*�,�UE1T�r)$j�vB؅	�j�h�Z6�r���}}ߡ��0  *����Iyy �@  UUQ�^��^ �� 4  �����y{� �� UUG����I}��|��R���[KZ8��2�#.�Ǆt��|�}�t���,ʖEZ��,F2c-cn�L�(�(�ڨ�Ih��X֌ѡ���r!�Z�n㪎֣(G��N��;�2*�Un�#ĕ&%Q]��d�YF�Z(Z1g�2&đ��Dh֛�V��(�-0��%��!E$l��D������k��J�\��D�#Y(�I�!�F�B�"��Qa�ɫ6Tʢ�Mҡ���ǋ �To&J�0�A"�����D�U�1�P�x��(�un�Ku��4x�&k�$��8Т
�FA�(,�d(�&R���� ��|f�]�2)d',R��q������P�h�n���H�kE�I�G�$�X�(�(9i�Pc��diW]�9�VM�R��Tb�T���CI��,��c¹R�Tڃl���]I6��HRv%���F!��Q�V��Z��V��j$i֝�7#�4��&Ӕ�ԒJ�υ��Խy*�_�g��t���:��Fx���U�y�6���x���S���U/�����<�=w��#Ɛ�iǺ�x��������8��8��=l���=8���=5��C=�|�Nw?o��zrau����G���>xT������dޔ�Zdu_�ӢMc�p�b�Lk��e4ݶ���p���L�|w�_�gT��͙"��ǃ��e�	*&d�kӂ.f�����8g���TYUv���Y�t�d�c�ݻ���:s��|f������U��}f�댛i����|h�\el�O���"#̣�˨��t����B��`��RI$|S{
2����Qd da�ܴ9�4h�@����ッ�����ѣ��f�Oi��Xe����Hhӑ��228�NK����eC�X� [��de6e��^��G�2}�Nj�K�ό�A��CEs\<$R���b��
�d7)�.GO�鱣n�`����)�Yu�Zy�qF�FG�#�}ڇ9�5�X�"�2�j@�W�J`Mcz�I �qTD��H�4 p��q66����x4�iF��vS��A��:d�ò�Km�o��={:)���-%�-��ڥ+_;�u�,j���V-�7��%�:����4>	s x9�%��$�˦C�a�IToZ�aa�<=��(4L��=	ޙ��Qѳ�z�*Q$�9\�2Hh�&��4�e][�^�DÁш��!<[���4�0�<�q�=^ƻ��I)�=�I��'�,C/�3��D8�u&��EUJd��G�.�`f$ky�6A|Mk��mi!�_�B�t'�M�����fT���,M��M�{�:Ӏ����i
�MB��a�@���'S���!`���r�9N�)���=,�>����ыy7*j�}��&rIv6[a
)�u�Z��"<�<�:�<GN�ѳd�!#�i���s���%�[���x�CGWaz<YN���]UZ��H�<Iv���r�U��M\��I$������M����U�V�]�����3�;��NO
�<_����ui�Q��+*�嘅�g�l.���w�Z��ر��L�)O_GU1����d��މΎl��ɪ��	���/%�3��O�mR��t���Wـ�P��HI��"��n;-c��d�#A���c�6�롷!�enH����~�C���E:x�����Q$�x[5!CO�Z�:poD��ɬ�o�rJ��HH�o6}��)�n�4i��浵l��9�(!���IJ�N�3�7�y���pʮ�4nX���CC�N����0ٗYF�DqG�E:�<�\B{E�_��5��㻺�`�9�I$���N���5�ӷF���lɃCFt�m�GdP��̯b�sb%�!�IZ�᪺ٳ��(�ew������?tj"d\nEc���Î���'5q^q�f�w�v��ޓ�$���5	�I<���4ih2[��Gif+G��]HBNZR�_W~�'SH�̼�Ȏ"#��8uyN��5�J�cZS\�$�,DI"r����^������<`�����Ju�Q	5q�[t(x�|i�̃X��D����B���~�æp�d��l���*WR�t���uO�Ӷ���9��l��_�f����B3ù�Й�!�9��O#�d9���eI-3�#�٦���c�؋���l1�8�sj�%��w'E���.bX�x�>�b��^L2�q��F��"<�#�Q�댦��u_H�:Ҳ�j(�%e�I$�_o�1�w�����AƵZ*;�x�.�#fX���������4Y�WK+t6�qP���D�ZU��&(x����`a(����oC���B���b�!1f�<i���qB��豕$����i"�c�K�n7i��EL�*L��+a�!���ˍ:�8��#���y�:�,sk���Mԭ���!�Hhta��7^�qA>�"$�,@�|S���8��d֕FL@Жb�V�UN5R)Kmn�9Ǫ#V�RI$x������n�t��r�]t)���R�U�c����j�1�W��9�<�NA���uz���p]GN�"#��E�C�YJ���Zr���fy���u!|�q=Zs���vqB{�PCl�nt�.���0����y�^\�}-y�W���w�e��L�2`
�ѣ�&a��䐼�$�:r������徒J0Ѷ��Oh0��Υ3����?���d�T�$.y�!e���
����U556E�`�sx�	/�w��g����s��iL���F�Z�DG���Ç��!�e���^d����|��jI$��i2�4I�<}����]9`Pj��̛��wrF�]ջ:��hy�tiႊ�O�	�w/.��F��L�S	h4àwZ3���ӣ�k�G�tn6W���I$�ʲ�1�ϳi��6i�u;4⎝4a���e��Fb>)�R<�fv��͜ �kbVֈY��%��C�x�#��uM�ZS
�ثb�b�j��Ū�j�c�b��[�e�^*��V�/V��V���ob�ձ�6��[�ۖ���'�nI�;IwZZ�����*յ2�iV���Z�[Wܵc�WUj�>��-N#F�c�F��F�V�-XU�-�+���g
�Z��-l-�-V�U�*�u�����b��[bեZ�����RыU�S�cJZ��V�jiKVեZ��▫W�&jص[�Z�x�Ÿ�
��x�c+b�b�b��[x��Z�O-�*յ[l4�:O��L>&�d��A'ĩ������ԝ�nݹ��S��.������j��-��UŶ�֯+�y�W\f�j�c�b��[U�ůlqlZ��UZ��KF�-�=qӒ�K�������I����H���B�Q'M秽
���U|���]����ļ�M����;���ݐG�Ƨ�"�q��9��t���a1�H�8ا޵,�]�#����dF��9���]��/������\gP�w��Wg;ݦ�_����6.�}.���m<׷I�����}�R���}b�4ήV���$B.f6�T�)��]�~��+�ک<�:�'�즩�q�w�f�uL-�-}��~�&�V�Xʻ��.=/�^�\v����  �}UU������������  p�&f~���s����� � ��>^����{���  �&fO����r�y��y���kZ-��t�8]�K$EEEA h�b�}S�����g��2��>1�� [ ����D������T=�Z�BM5��P6"�5D�Hvb�|S@LC��]��}�4@���8�N�������r���dn]��P���l���c�!�&��!��V�j`0G�(�����,C5��'Z6A��pY��@Bvdm�3��>�Fȗ���`p��������%$�Ʌ�Xn#��>�WĠ��� R�xD!���Z�0��}�_Q�T�l��4��q�yo"�-N��4�~�3TՍ�l=h���$J+uZ���	C�; U��N,�	
���GH}]a��-�-��Y�I�6|<rZ�A��hIgUa����`m���Q���Q$
�K�FM l�FHe����d$(�d:�8A6xr���,��œd����t02Bv�� ���}�'<E���:ߚ;VQv_�$
 �D�\K"��p}fX�L���[�d
H0~D;]!f7J��t�� <ÌG�|Ù��)Ӓ�0#�&h�f�8`�ո��#ȷ^R���9�r3�=f�7�����4���q��%�l�ym�4TC)�H��&=h��pZ��$L/�J$��F�I��fee�[#�^Ho}3�TTT�����H��l|�Xʿ�FXU��������G|}�<#��PG1����t�P��E��;�}7��%t�霉�{��#;��*���\���֩��-���{��w���t�\k[t�{Bkm 酼�.F�$�'���$�ȇ���`��&�����߰r�)\��>�pa���6�� ,`h+�QE��.�>�2B��a�،���A����sLe�ro�3��^��]�2f`��=���ީݶ�Ӯ-$��(v1h�m�EA>h�t<Ѫ��#��Jo�F�=`l����6>C�b�;�A�����'~{�V��
�Q������B��
Y�qs�M�F&�!�t��a#M {ٵ��L��YO�mO<��(����"<�#������G�tD8]�b�j��J���QQQPH�R��<�6YA�	�`�"��� �Y�X�ƙ�T���7M�@�ܑ���0j��·��M@� BH�e�M���pq�4@3��L6J9�QVdA�w~���!A$D1��B�.cG� �J^L�(adM��L�J>���n�"c���I�_��O�!�\rf��u�ɨW� ��%p!e�[����䁰�|��JR�C ��X0�ჱ��F��Whݘ؄<4�0�@〠6�C�@�A�@��7�oH�ө�S��ގb:t��/̭m�?8��"#��Z(�f�g������H&C�EEEA!G;�4���%||D6ꁡ���J��&�R�:@�b�Ly�����Bm�P��ca�)a��P d��Q�0�]J����F,l�٨2���X¤9�0�$>�p�y	��O�g�C�
�s���;�,-.������ml�"X�s[o=-O��X>�I���A�����{sf�a���0NC�-�a�rE�Ê2�kf��D1 tA��,�H|�{��{#�=T�m޳$u�����E��#u��,����q�<|I
NqQ��x��q�G��!�=�1�}��8���Q���o���"<��:�yh�̺�3����x�N9��,�����QQPH�u�=C�$�ߪ�������bbN��KMR঎�-0Z\��B�g��l��k�2� ɷ�:*i����<R��Ym"{���>Q)x� ��%t)0@��~i*c���`<4O�:��1N6�v@5�������0�|äC�,aqzA*&�(Ό�eA1Y���L�  � B�sݚX�J(;�{�a߉��	����ۺJ�d�vXt���|:(�t��`	 i�Xh�a�%Ta6�.C��ɳ!��ɀ�9!������=�qE�=2z7�t���ONm}GMc�+qM���[Ϳ?8��"#��Z0��J�&s�P�y�]BF��rXDmbĈZ�L���h�?'9yJ]g9�T�J�P�a�7�v�=M��)d��*��y-��Te�&��z�ب�$}���RN�̮����/�%9�l.k:$��o�����{�&s�ڟ���T�Vΐ�T��8S���g([	�hŽ,���޺���wy�V����!Ƶwf��O1SfoK�����xy�_?�\�HYAeK��nd�h��Ɔ̑�Q懄��!����K��QÃc ё��WFh<:).�A��D a8�0�f#�'��,\1~}@�y� tα
�t��(o�IP�<>���l�G�w����a�˳:����X>����,r��#�}�=!�7�]�`��t��m�_��٘Ą�c�� �错הEaL�(���KM��P�L�F]-�3ɞɼ5�K-�z<�O�����S�X$��}^,��CL�E�9��%�1h�Ai8�SUf�z���C#E,c �" ���ҌP����3�C���U�L}�8��^e����"<��:�yh�δT����ƭ�:Ѭ̘ڵu$�쇺���AD�3�ϲ�mF��v���YP,�ս۝�J<0/$d	�5�m6�p;���@��&�@� �⇇0���8�̙r`J �$��992���w˱ѡ,�h�668,`d�cm)E���B)B@���Z�n�����B8�sq"C����?bX3�����2Ǜ�W�T�:<@�F�����X�qda��R�di胢��q�K���� X@�9���|J�.`��F2L=x4;e�GR��2�6���"<��:�y��5��m{���P��������p+���Ö����@�@���%����x�!��?T|�p��䡅���� p7��0X���\8��<�w���{�M�~��w�����n�烰�C���<1r�aC���ɜo�N�4e�0��b8�� j���-�o��H�8��	���o%��f�!�w��sU��o�cx�ᮿ!��G�1�v��61��)Ƥ(8@���G{ɖ�W�j`=�[�eBPd���W'�2e�F7M��C�'�2�v@(���J�ÆM�6ڜ~e������"<��:�g��x�3�y��ce��m��&��a�"���������ufotC�RT2�ւC����ˉ�� �i� ���a�'�Ş �<�V;F��c}I���������e�����F���{Y�uf1�0�,Z���0x���Յ��2�26&tfy��Y����0vu�#
�@H��P(;�4t.�&M2C�],kYe�i���0 ::�����h�A��j3�3�3a!+G�A~!9>u	�I׃��A0Am�e������(v��0�,4�P����^��W�f3;�Fd���+�b�Ⱟ��S�0��kc�qq�����ڰ���lE[8�b׊�-�-V��o�-T�-V��Vū�b�i���*�h�ϕ�y��+���O�Wª|);'oW8�InӴ��k÷Û÷7i�v�����-X���Z�[QKRԍ��ah�я�^U�TU��q�mQl6�:Ɩ�*�j�Vͪ�bԵZ�QV�U�ՅR�V�0Ū�x�Z�_[�Z���؊ql[U�j�6��ڭ�U0�*�ū�Y[8[�WV�ձ�[�aVU�[���U��՘�EZ�KW���x�Wf�$�k	�,��>%���'�?K�Wj�������'kڸ��N�s�'kv�.ׄ�=kxv�ej�W�y�WX��Z�Qm�Ū�Ū�^j�V�-�U�TU�я����۞��t�S�;'��Uީڔ���R�T�S�~+�W�s�g3S���l��§eb�$���ƫ{Ҝ�9F�����ȎtQi�;w�����;dGu���&O��Q�N�|5��U)&����ٻ����o��q޽�Ӧ������zr�����9F��?}}��)�B�!)�&pұ�_�����%n�SϏ�����WwNZuK4c� oj����3��j���ԉ���/�
�ȇ�7=�O�>����6�d<3x|���.g��BY����}���E?B�V;�k�ʭ��MJ<�{G;��(���!9:���[�N
ٜR����8��י�D��ŚV&�.�����ѕ�d�n��.2��/�������[�[�[�꽏����YP��z���'�{��������ԇ�P�S�c�Y
]��7�ˇo�e���D�\��r��)eR�,I�T��nʔ�Ɏ�5N�����l�+U&������KT�V2��O�Kt�H�+.V�\Mjz֢*�.�sSMh�����IP�IYIa"�G�5��ٿ��j�&A�>J)��3F��TF��K�3�[joob��e��WQ����<�k�����>_}�  ��>K��������}��p�&fO���������}��|p�&fO�������d�������L�9����<��e�^y���Dyuy����H�ln�
�]cB�i��g7ې�������L���r:h�OH'JUh�nU*X�!$�7m��1;S�P�)AA�<�qr��M@�&'Zu�5��#��B�\�Z"�U�R�u,C�ʈ�h�B����"N4�V�Y.WGT�Et��jT��Ɗ"����E���iT$�&*(��A$�q�v��<���+�(�HQ�E4�1�Ʉ6��\��HpY��IA��R)_f��FQ��:A��Lpe��P���`����*M�(�B��r�m��UJ���Mi�n'T����F�I�T����G�,R@�����#�IR��W�\�+5�"j�N:��bu;��j�Q�b�e��ʔn�n���Q�k��G��J��J�A�-��(�A�X�u��+�	2������@�e�0���#��i���$sE�_N��ݑ,�J}>�K����}����`�B�ֳb�c�o���X��u�C�ۆ���Ҽ���4ZB����%%��~�E�~ߧĈb��n'�Cv�3�i�+L�c�����.3:SP2@![!&^�z^���a�i�F��Z6U�=�t�a�b4��e��<0R���v��<��[N���r�Nu����϶#�RV(��NB����5
�Fd09���^L�a�%���@����65A-�8`�:�o����L'q%��N�&Gèd
 ��⣤mIAm����{�����tF���������n�N�>��_3M����`���dv<`x��8�/��F��Θ���}�&�:�Q�Y~~m�n"#Ȉ������~'���e�mЗ�N,cR�Q��w�ow���ldA��þs��;\ lԒ�U���Y�T���G���O�����G7���4Ӛ�s�K��cl���ۂ#q������$$�Qbg�,,4��e��li�l,0@85Z~6�m�CǱ��Ad$�-��39L�tgG�� aDutmS��+44�|I�+�_p�1�8���0���f�;�a���'Z+����q����IA��M;�Kw�pk���c�h9��fʡ�$���!FTӬ������DG��QO<#�㧑�=g+�=�Q�����jBC =M��;�#�1��e?~�;$��ItΙ���ܜ��:d����?��<ј=i�Á0���d�1�� vP��[����e�����cₐɫ Q�G�Ќ�/��j��ɭ���+�w�vy��c�l>HC0=X��$�Hdٱ�����d!D6��0�E.���g�m�9蹄�Ə��h[d
`S�Q�T���M�F(8�'LY	(~���{}/��O�ɤ�&�u�#Y!_Q�GŎ��+�����#D,��f��$r;��֡Q&(w�IPx�#E��t��ĖX�s�ZR�e�Q�����D8p��!����60�d- ԑקc�1�����*R@?)낦Up�	���7WM5V@�PM�|�d�L:#�d�HJ��O٬Ƴ?҇�UXQ{�HS$.T�*�ez��Ï2j�0!�ZpL��W5����1��BHM�ae	�0��&X.;���8B�$,+/�J�#�4@�)���6T��.�'���\��k파�lm�!x���x��&3�g��Ht��! �D1�������!��.��!���0胝�9o4bV�u'�!I4>"��������ӣ�4A��CM���D4Q�#lp��P�t�6Y�(��ߜZ#Ȉ먧�S�u�_�n�M7H�ʎ���>c���k&A�j��y�Dc��AF;��qn�x%���
!D$E�R�27MLV"$;��q4�MÆ�&�|�?3�6ҳ?6<5}����,�s���n*t�gһG}ں��[J��)u��Ը[�][�ڵN��"���k|n���yR���S꾢-�q��ur؇wKH:�4������j�V�����7�����v|I���MoMr�,�}��PA�M�����BG�Q�s�trբ(�C�M�Z�:B#;�7$74`�h
 �v�x�,���u��4N��l���d���J��S0nm����|�ѣ�x�ɣ��!��VH��l�I��0���H�'r{L�O�����
>� .�KS0��E�!
��@�D'��)�uHv�I�%���e5�(�C���p@�L3�v�TxCc�6:^lj����Q!�����Cd���|u�"hc"2���@�?�����3�7)�M�(pA�SD3��h#GN�%e�Ǔ�+�UZ<����S�`��î2�+[o��-�Du�S�)պ�*�k*c�޷sq�c�H�B����[m��#i��v@0���J1����'3fY�4[��@��O�RF����EŞ?���g �pq!FrR�#p��U[�H���ֆh��%9���jJp=4���sN��nӓ��q͸��1�bHB����=��	�7�?.��%ձ>��J��?�ʘ�]c��G��4;�Xxa��ս�ap8@,����g��
;�eŎ�>�TA�A�G�L�0���g��hqLr�(˱���X����VF8�Y���SFy�Tt��㬼��m��Ţ<���!Ӥ8|q���^�ڻ�[3�q�c�H~�b���V��y���,�F�dp���s�'4;2�1��4b��Ӏ���,H��;��d4�q�Y� �J����w�8iĒF�)���˲�� w?8>��Y*Y�VF�$�i$�p��њi^��nx��t��[<Q�7�́Wѷ���҄��`b!��ݸo��j��3#lK�P�:A��r��|4�|>i��D(�0>v%x�j���c�#�mS�;qI�&�*7>rv�y����1������ƺXV�J.�ٗ�
j�� ���h��mX�˵��U�T����6�,#�#/#k~qh�"#���yN����0�s&�"JAj-TDWyTM4�M4�p����bKm�1�g0	\ 
�C��,G�l�"�9G����w?y7q1c��a	��۽]1��c.ˇ���A�Y�i�X4p�7f1�ȅ�pB��8KoF�/��.HN�|0��J+{��4��z��m:���44�8X�Q͡���>r`<@'	�6]���yy	7[ J���n�����M�m*���ё�@���Ln������C�JH`貍�7H@��Y!V�EzKlw6`��1��,0����L�K j�r�be�<h�|�~�}�`��m2���?2�Ϳ?8�G��QO<�V֞�E.�:�К��Rp�;t:7Y˝�tӭc54u7f��64��=I89a��u1[T �J���v{WMC�P�Z�yk���ojɎ���q���s���=N��b���oO��5��'��6:�\��\��Y�l*P%9ox9;Y��U!n��QK+.鹚��V�ґX�!ĺ�Qp�s!��:am��w;��u�[�d^w�O���#��V�'���j�3�����hR�� {�@�oۂ㒰H<!��9�44�����'���ܵ���`�5�QG>y���U���8	�8WL	���oi���5��g�kE�P��H�ʬ��0�(q��Ð$r���\���PW��u�)��P�\�:��1z@� a�������5U!xd~z4ߝ66�����	0\C�oO	S����bL��)�c2�8 �~gߏ�dh�U�յ飅Ժ1�0c!��*���c�EX���\7<>>q���H0{M�h�A�,��E���x`-��e��&�y������yu��uZ�|۰�i�Wu4�H1Œ\���ɸ�1�`$��u�}��o6��^���Hv�!b�J�6AףI�:4�c��yiqp@�R6A����D��9C�d���A�cTQ��^�#)�#��<6QDh�/$��80t�i�c����h@�#�Ϝ��S�CZy&G-l4@�zO��a}uT����Z��E�,��kF�a$��,�s�3!�]|a<@�}��.�El%s�茊�2��r��.K�b��� �z��0\�%V�����	�$0���$cJjx

l��,wrM0iXW֢�Ӭ4�>Ҷ�8�L�|L�S⏊!^'������|O*�hŶ�jRص[+f�j�صZb�H�U�����0ښU�U�Zv]�-ړ�v�ږ�;L*Եi_Y�>��Z�R�իR��^Wߕ�~U*?0�~~c��0�ahŪ)j��E-Ql"�Z��ϕ�4�)V�[[�q�U��jE_U�U�ՅZ�U�ū+c��Z��*�jE���-[q�V�jqV�VԶ��
��Ɩũ��k�ylں�m�/��j�2�-x�-�U*�j�Z��>یZ��q�*���e�U�*�X���V���aJ�Wn%�ߕ��I�no58�㖪U��iV�)j�E��+W*����E:�Z���m�*�Kb׊�ٵZ���LU�*�h���8���t���-;.�ӕǣ�ԝ��R��S�qOʥeG��c\���+2�#&��T.��̷e��7�m�l_GI��_m;m[��F^�W��©�hf�q-f^En�E�nي����8�>���2z�r��Y.�TFfmTr޵��4�M�d�s��"c��k.6��u��K��
ƀ�Z�̖ڎ阞��\[��x���u�]Ҝ{Xgel��g�Ԟ��3�o��_����\���*Iwww-ws32|��������||���f~�������� �|���f~������� �N˫���9�|x��y��y��mkqkG��QO<�X�o5�b�XM4�M~��k�M�m��s��t�F6X������d�[ ��	8k(�X� �Zph�Ph����܇[��h���2H���`��b|U�Z B�T}I(pP졣���;��+f�}��NN>�.s�R��o)T���"ʬ)���e�����$#��İ'_4YD �!�-�#
�̪�[�Q� `����m�fHxo�$�x$ }�BC	�#���tr%���2�NrD�P�,Gt�X�B<,�\F �ϳ���RS�Y�ct �}`|�,?t�f�@����"b2b.F\�RCm������f��Ϳ?8��Ȉ먧�S�wR@XK�s#�1����~s��=���xw[�Q�c�1�QI,�hax�)����6į�vC��_P�P�6�0��fT��
%���8۪J��'z�0:g� �^성ߊ3ѣDg�(���䘄g� �vŔ��a���@����OJ�\x�Ns����?p���@!��1���i�!Ё�`E���7*�#�4	 ��X����j�h���%R�x7�"C���W�/Ǆ��R���C
�*�5 �B�8G$r���C�� Y2�nUC �x����`H�$�r�65�dHђ�K�i�������E#N4�<��ߜZ��Du�S�)�;�e�~�}�����ղSzj��ɐGx�jntѭ�#���ۖ��5��� �WY9]v\M�V2�%��T�̙w3�f��+BA�k��f��{=9�~���E�LTl�މ�D�y�/fn̇z��\��5p�J�P��j+5u�Z�Ψ[6��Y��֊�Nx>9E���f���� Γ�?t�}�=��V�ֈIGB0�6i�o��:�Cm6�y@�
�1�RY�����J���CD	�=��*��~
{nF�0/�'��!!�8��M���b�oͲ����=~�ߒ��a)�'i����g�
iJ����nc���p�U�0�"�a��(0��@[�QǃTC1a��O�Ɛ-���\G�Y��G�5
m:v��ۃ�.�8j%5H���>>x� �/g�7,X�cm-o����2�S׳�2��:�2d1���F�<|跧G���2}��l�*[�/�4����Z�DG]E<�o�QU�c�U|�EEhHJ����)i��&��L4mrR���}�ᐆ^[�<�k�)DG���,�iۣ�"d,�n8*�G�Zl��H�@:A�+������,`�!��0D6�+?T�r�����䥄*�n�,,j��}_7�\�h�Ą4���Ye�F\���(�B�	�mJؔW�Hb�"d+@X��0��i
!���S�%��Or8sM�+�N��h�p��Ƥ�nL�'�N�:SD�~�a%���x}�-)�~q�帷�V����N���'w>[������������$.�rV����t�S�?�P�8�`~l2C��Ն̗�e�yY6�J~c�4��S�~�c~ݑ,�á����	�����p6J�A
4Cod_H˦���������+*�T����Z�X	T;^I�a��vYx�����Κ��o\<=�7�w��'�#	�7C�ɉ2�5��m����.�9�B������:�X��K��gK�ˤ��᱇x`�x4��!9z�c�>9С��X�g��>��󌣍?-���^<x�ӧM�:C�l䚆��r�qU6� O��TTV�����A�� HX��O�G$G<�I���������҃�%��u�he�j��R��תI3;�7���Ɔ` �h֣����*���e����;��צ��c�-f�	:�͐��wml�<B�D5Q�!�Y�S�D$\�h�#���:���2���m�r��,�<<ft���&3��!��2�hlce�h`����e�?���h)ɷc����Z~�%L8-���4<n��V��������Me����>,�KG��ַ��QO<�\���y���}8�/	�I����/3#����D�Lㄸ�6HD�i7���Yv9�Be���F�eɣ�������}�������ޕ���}��K��"�-���R>��zs�ӝֶ�m:�j�9�Ӿ;Ntu���;^��2qw�綮Eέɹ�Ꞟ����/"8��o]�綜���[M��i�j�-�:4���%HV=���~$	1c��â>��
g8f�˗�h@�<�p�3�񀷇a$��}���z��@��hn��B=pm�[xْ��_��H{]#�Te�v]eoީ6>�	���㷮]U�Ӡ��Q_C�jGL����Đ�Ҙr�4��u�^��hh���vP`��X~0���(��ܒ�)���!�%46��뒖Ĉӂ|���R	���k:��.|��C����<�=Ƈ�Z0!��=e����v]�ܻ�}_M�����Җ�/̶�8��V���G]E<�o��q��b��f��[o���BXٯ�QQQZJ�������LTP���S&@�Ɯ�!m>v8#����6C��FN_Y(�W[p�o�pj3f�I\�&�@�>B��/_�����x��m��`��O�q4ш��fk3~a�'�Ɨ>&����/OHI���sy��I�����>��C{/!�j0����ta���D<�����BI1����[B��aF�2T�ˑ��� ��M��F_�m�n??:���:t�G���ۺ�����5�*�7n}�EEEhH}��|ՙxbd�fb�Ie����#�M���B�A��c�{v��d!��,zS�oTyK.��C���U���V����S�&�A�q/���uM�9��@�|���:�L���礙[E#Z��ge�c�����L(k��ސL�����!\2X����K�M�zՒT�%5
��۳�C#�P�6��G�C#��0�\?�RU06�4s�ȥy3�bv�2�l(�����U	E�r;M�hi�L%���(! ��'
ho���C�?�ѳL-�V�2��?8���kyh��u�8��J���ȶ��V�% ��$o����['��**+BB8Y��
�´l3Uo]p7X&[ B&�b[�����d��Ũ ؖMl 1bhU��X��42E"\8.����}�3��o�d�ɧ|�nn�d#A��`j)���!�i�FBprgG���3h(���u��e�2e���!���Q$(��$2[���&h|����u���g��?�s�#&���G^�!�kBa��V��uaf�B�yzѮpt��捈Q�d��eM+��0�0ڭN+�a�m�_i�-T�<�Vo�f�j��f׊�[�U��հ�صZ�����׊�y���X�U��6��W�)d�T�KvNԻS����	�]8�L��$(���|C��Ɗ>!�l��V����V�F[Z1j�Z���[�)lEZ1�u�4�*�j�fՋW�b�kb��qKU*Զ��?4�����۬~W�~���j�-���֮)Ű��qV��J�V��W�����uX�Z�V�o-�V�m�l[Z�V��V��b�j�1j��ul8�V��[V���66C�Y>,i�1!� ��Iv�]���ݩ=T�^j�R�t���M�ե-\U���ej�X�>W�ǘ���Kb�b�l/5l[lZ��uy��E���V��ʫc��K��;'d�U�;S��d�K���!��Y>��}�_���Ϧ�Y��1ji]��ѣ����#���|�[jZ�q���'Y��-7����_.�5��ͦ��:���ʯ��ߴ�
�z�Uꉼ繝��5�����m�]xԛ���ۜ)3w����ᦡr=�!��8T�;�F���O&�c5���R�Mf�hm���S��n���[^���o~�β�'-�m�;v�XXs>g�j�\�OK�;��CmA�oᒃ);���N��qU��ה�3�߸S��gi�}���p��pT��߆](���c5n�"r�2��A��v�.�;yb��`�ro2�J�ٝ���U�����m��WD�Ȼ�<��ډ��|P~D|�4�n��O�?��|xG��~�������[5��:�����d�t���$UAk�^��#z1W��U!�QD��+2!��H�I;��PH����u�GZv�;�TWP���m�-JIU�IKk��BNIY�%�ʉ�R��qӓSm���V�����  ~}���������}`@ ��������� � �`}uU��wuww�X�����{���T.\�̶��-n�kyh��u�8�Dm�!9ch�Ɠ�!��[��;m��aJ�j������ڱ�1�'a Ӱ������,N��\�h����I
�RHl#%��tW
VB5\�n28���-
XB�尪Q�!F�촱�A�Gj��d�^Q0���
Rd	���ɖ���&A�\�$��R�`�f	�E�#�Tv1:�i`�Ȳ�cC �,@�F:Uj�y]�4<)FBZR�"<e���A�Ȅ2�82R)��)��eq!����T�(PI��8�!\�[F0ju,,��J*�v%+NV�u��(�i2(�Ƞ�IF���[m�iVAF�"���[��A[��T�vA���$�LQȄ�x�`�#�����R�Bֱ���ڱ��,E�"r[q�+i��U�Q�ՊJ�i!�Є��bQ�+���#I�KmK\����E?sh���	�==}͗Y���Y?9�]лZ֐�~�v{�l%y�b]���� ���C��}��)<R�s{���������c�t���|���IHk������>ص�ou����R���(��)��������tS4(��ْK%�A�a�9x9�;�G#�,!8��S�2S��]5�etJÜD4�'͗^[0KQ�=r�T�7����$�V��ph�c3�)'d��4B-{o
(*Q�[��o3fJq� �O��f(��TtX��Y05n�d�?{LM�0�W�N�J�_B��M�cg�|u� W�����>�8�,4�Ke�����ַ���]S��JUW���L5Z�S���A��L��]EEEhHX�lh�9*��X�nO�,��>)�M<yT�e��6�f��JR�1Za�}��z68��9HP豁D=��@�wbCa݌����<��?����y����xq���v��Bܮ���%ݲ��R����ģ�+4I����/Bl����`�&��/��0C��866�Bh��h;i�������87��M3�֨���q���2��i�[G��V���G]:�s=���j��JS�i$��э��6�b!V�j���I�����ɔ?��a��]��}G���oL>�ΰ|�6C��
g*�O�:8$!�q��`�c���\4�`�6C�Y^��r���S�Rc����K�wKͺp�H����l����M}���a���ȧ�}ǌ��u��]}pO>O�z���o���eo�g�ۭ�d68K%t溈#���`�B?��	!���A�������<9ڬ:�,#�?2ۨ���ַ�������bL��|��lq�*3Q�J**+BBʳ��:I�ٲ_HIa�k'7����?�$���x�!��%N�c�&��"l�������dp��:p��4!F�6h�4;�L�B��+��H��.�����*�R�qW��X����ߌ����p�d�&}YJ:��������������2L�J-�p�B:����$+F�PQ�?8~𦕄��i��m�
S�ig�q��kn��}����n��N��+qn?-խh�G]:�T��;��Fl�<=�t���N���or��҇e�e���8�Rh��!�ޝ���M�&����T�v�ءm�Y�}�"���$62_��O}�����{��.s��<��M��q���~��e�QcOi�x��&s�r'�zu�c͕*�����DUL>Q���,-o.��'�+���?n�	FΡX&C6vG����}%�O���J�a�`~�A���=ɣSC�/I!������Q�b%��HBD8i�(_�Ĳ�\;�Ǜ40(��$��Ɔ�((��o��Ѣ�&f|Q���p�XQ͒�4[��6�1���$�Ir���I0���!hز\|WjW	��B2��F���]�S꤯�EV#v���q�>ѓ�̰��Hˮ?8��V���t�q�f����Q唎*�#dXDT~���UEU%��G�8�<hv�r�c��$��+�u��5z�j�t�M�0@�&�C.�v�CƜ�B8C9�&��3x�ioD�Y��Q��B���i�փ�NN�vp&��Â�43b�S���j�����C��p����4G��	��@S�N6,�!Of��#�ή$�s�3rA)���<��E�����]S��q�e��"a$KE�{����	�"+2��`k$��
Hr��0y�޵���n�$64�e�,�rB2O�����J�v,��s��V�F�p;~��DUJrGy9��2�������>4t6}'Ð�.GG^䲬0WI٥�>]���7?�!� �� �GIO���:Q��f���8x��p�-�/NGEhh�:`��٪�l�F�?��3�@�∥:S��m��W�V����]:�Vq�Ƴ32�n�w5�����А�&V�Q	���s�}�!c��p<:#GD��S~�~�i�tC�/g��muie�+�ڜD8��#9��&{4���,!�>6|�[�w���"��z
~�� �D!{< <���Mn6�$�b5���
�!�?����d-����J��1���u���5�Q46�פ�����'P��aD>p��}Ӗ���[�#|H�0hj�k�M������)�Γ��E��Jq��i�~u�խh���Ӣ8x�!`�赸������ȃiN��q���Å��g�w�Æ�:��z�����n)ݻ�+S ��U\L��mS{���4=3�(���	g���ޗ��9�c_DO�H���(O����C���E��Ju���n�/M�q�w��iN�G�M�ow�S���9�k�~��N/в�P�U�]�^��m4�"72�o�w�w�QR�	\�h���d���o�6u������TG��-��.JS�i�K�Λ�f��W(��P��=a�pr�ަM��W��,��W���OVd�|[ÁD:��S����r<��?8O&� a�3�L8"&n3��?����~��{ʊB&"&�k��/K��{zÆ]�>��C�Ş%��C������X	��1K۠��+4N�iO�6�4�O�q���V���t�Ä8&�d-�ҽ�T�V�z��qc)��3���**+BA,�!����f�u�C��Ñ��<��s�?9����rv�.�\�HI�����
û����eE`a&�!a�@�Fr;x?tv%��B��.}Fh��i�ɳ�t6L�B�@4m��ɟ��>�b?u{�m�Ĭ$w""��D���HD��w�3�x���>ud�����ᠢ0���$'F��qahQ�L��gE����C�&m3.����Ub��??}]}�1�\am��]i柚q���#h��":��(aH��#�"<���8�6�GЄ!DF�Q�e�R#h�#��:�#Σ,#��8�#��#�#θ��[�ym-��j��(DR#,�6�"2�"<�#H�4�6�2����i�GL�H��"8�Z2�[�qm-�^eF�F*���G��ґL0��2��4�:㮺ۨ���iDF��q�DGS��6�B�����a��u����~8��lǎ�lÇvӊ2q�{��~���H�<�����64��y���K���3j���+�d��4]���K�~��#���1G8��S����9B�=��U�ī:�(��\�����9�'wi:$�=F��*���s��=��e�;g^G'�yT�Vl�Ϲ���U��WE�^��]v�\�g��QѱTI8��Yv�6O�<�َ��"�jbfr�t,@�_�U�wwuww�X�_]W����}�}@ }u_Wwwu�}�  X_U}+ܹ5�4�O4��uպ����u�8&��������**+BB��ޖIE1T�鈁�x[�-2�#7��B���A��0�A�����ǜ��'�\���u���בO}Ƴ�b7����S�Z��I�]��ˤ*�ڒ͢sX��G^'r!��Ē`�S\���N��9�|X��2���V����F<�(�:ӯX����\��8��%�O|���և�:�����8�C��8�#l8��q���]~ukZ-o:�:3�ӫ62�;5UQR5���2�SV�c�g�ZJ֯g��**+BC*�Ƨ6�O׭&�e­��	7�ǝa��A�y�F:�ӑ2Cf�����%)��Mٶ�Z�O��(H�i	)f��f��joT���3��t��>�GÃ�x�C6H��>p���B��6��I���M��*H�<�������q��d6�d��<h���n>8���{���˪&V�{F��%d6C&޶�'�v6�pp���6C�!̜68x3yoϰ�|�����Sl8�m8�ȷ~ukZ-h뮩�b�����g.�6,��\�`ۻ5�8�S�Ad-(��Kŷwco�K��6�G�dJ׍�,�T��V�ʛ�M~�����$7��xzC2{}M}�e�T����79Q���I��כ���㜿d��}��v�k2�r�J��fE�acj���˽�]ֹvl7z���1�S����Ak3��'b��PF)�~o�
���ٓͿ|6�8Pp�u�0r��J���N�p�;��@˧�Nm�k�Cf���f�􄳅�4�rƍ+�~����z��5�����T���Hl#Mƞ��$��۱�#"M3£ޛ0;筆O&��x4Ӏ���8h4l׎��d�4ۛ�J�)���ⵔ���]�٢S�.���ˁ��8,�(�Lwzc�������y�y���<�]~ukZ-h뮩�i�v���H������� h��2�Ov=�@��B���V��p�9!	&Ci�ޛ
8�IojKs.M����N}=�4��:FC��V�7k���p:s�@6t6Pm	;�i�����Ua�܍�yJ�*�����ҿ^Y�����3�~����r/�8�?`�}_q��wM�B~��d��$:9�x�0m��8T�ϝ�Q28����d��`~z60C4d��:��խh�����XqO��
��V�RQf4z9��-��*�>֑QQZ7�%�e�xX�!�ql���C%���=>�O��a����҈A����7����?����Ģ͒L�M�e�%y��q��_h��p�8a�Lߦw[q�)�ڴ|38>� p�|FS��ˣÜ: i2<0}�2^C:��󓵊�tI$l��!����}�>���,����&�S�-��F��[��:���u�T�:���		��L�IL�s!U���**+B`~>����u¡�_� ˻����;<�����H�;t�Y+����<�~e��y���y�?nxCǕ�e�2Ǝ���+oy��ﻴ��M���v8�$tC/G�h0�H�4�Ϳb��y��'ܫ����������1품��:gs��@��p�Gp8<��Q����B��!	4h}��&���GK��fr)��}�*>��}�p�
i���N�����:���u�T�)�إgGEvЂ�z;Ť��]�����sy�����]�8��S�w�u(��G����G%�1�[Z��э�QZ�bz���﹣�u��8l̽}����]^�d�������5T*����^��}��F�{��v���*z���pb�X����y������|M�ɋ��[�6��23�F^)��猎���I6�a��9��#wb5�ux���]�]]�y�����-��?0,:L�������G��΂��g���dx:]�!�HP%�㐲�MEP,J�e����_l���q�<}��>�!����f��d��tg��L�Co�$L�cϭۑ��u��c�C��C�W�:7y#�9�vS��7>%d.s�<��t��ʬV.���Z�a��[u�[�?:���u�T�9��諭��§q�c�R�E����F�n��|��><T��9Z)2���#���!��F�/����$.�'����L�$K8x,�+�r���Ӝ8Wg'9xǔtH�����^6�ϲ��W�?s���!�>c�ç��]J��灃n�}�$(�*t�3����3��Jc?���_��~r�٨�MO�4����l��'
N�ǭ���ڪ��h�A���64��6�!�����!!��S�:�[u���պ�ִZ��]ќ4�ʯ6��{���z���x2���@��-uEm%"�˧��N�<���<����X�����3��<T#܍8"%��|:|p�3D��e ���4D29+xG��D~HE(��T�$(ۻb��|���$sCP�;�Ç��a��u��WZpSцL����ѡ$����?g3ri�2��!x��_ҡ�A��/@�:�
7��Sa�}\���,99�m1eσs���8\����	��MQ~ᶇ;,�0��-���:��Z�kG]tGFp�����q׎[dU6��&K~�EEEhO�xxu���]�%���$J�r5�Q���u5߿i^����8��I$��F4�h������ޝ��zl�/X0����ϼ^��(����;:ON=}�'��8t[�!��Ιq��l�~�4��O��Æ]FF}�tJ*��N̛o�,��xSmt�1�x��f�[/c^~��ʨ�U�\���{o��nO�?w�t�o�ˮ0��m��j��M#*B")DDGQ���Di"<���q[F�aB��!��#H�4Dm�qGQ�Q�0�#��:�""<�:�")G�F�o-o2�֥��F��*#(�#͢4��H�/3*��)�"":��")DGF^G�ie�Q�aF*��B�#*Z�el����ֶ�q�qh�:��"6�#��"":�VѶXB�!y)��ƻL]�g5�~\��;�Y'���b׫8��m~O�V\�p�7] !�}���%�����;���j�{��4�s��弚#NI�Ҝ׉A�KJ�Qd�P�"���*!����*�"�����֛��1<Z­��jV*|J��~��z���V��T��噜��o��}Y���:��MLy�Vo�V���5�"6hv��J�پ]�%��|�N�����w;��/up����9��oĴ@��א�̚=-c�ۋZ)϶b�5&�\E�up��b�MLr�mҩ�s6�A�������ļ���?c�k�������U�k�WW����=ϿR�{�²GTJ�RH�dR��HZ�SqTՕ7L��m��Hb��r�����b!��v!�e�2ԅ�Gc�2Ĕm;�b�:��4A��h�!"i�cD��b�Q��Nb�iW��|�kK��
 ,
�ʯ�www_w�P@�U�W������}  %W�_Owwwg}� X�_]})r��(\�J�ʗ._-[�ykE�u�:Ì磌��f�F��씌�&�\����X��IUWU��YRU�G(��d\j�����D�۰��9�Ti<b��h�Q�B""�#�ӑU��rR��e%CNV�%!`�\��Lo�Qɔ�dk�	Tn������G�b-0�L��2$�u��J�c�!̤n��K�L!���I�
I�Xբ��!<�h�xB`ܬ@��(�w	(Z)' ���E,��i�&A�b´GD�)���eP@�.'���,-�I�$`�Bhp$�Bh�,�T[�V��*M"ʆ䑎J<���]l�*�DX�K�q6Z�T�آ$YG[�*Ցܨj�1Y]�M��d����Q��%kbx�n��4�u)��J�RUQ���Q�i��"X�i��V�$[�2W��c�8�U�Yh�k*mB�ZV����o2H�a���QQQZX%�P���Z�܎�����Z�r�\էJy��H�N!F嵯in%)��OR�t�l��Z�:SZ�����Rb-@��q����K�j~���=��=ēx(�j�V�He�例�譕�T��.	e��g�~�BO�!�g���IS&�;����Zy���O����:W�����s.�u=�����7Tԩ�W8~#vs�T�P�Cg�oU<P���!e�9�'�d!&�48�	��2>-ɉ�/ݨ���8Ό|MHA��CIA+/�-��d���]N0v^�;����t,����ˬz�ٷT�m�������[�Z-h㮩�R��X���|gxgZ��fD��W�|� ٽY�~EEEhOV�[5Ye;����I�#�w��eUB�%S)�8����\*4X��6l���	<3��˝|`qn\�:5��n��G������>Ol릺<0K�Ҫ����h��$&�>�cX!�E8p�)2㐒�=:8>����v) �ne�	��B1�pw⃧YǇ�̵��3�I��x?�f�Ec}�9q��E*����8�X~q�ߚ~~~u�ռ��֎:�a�[�W��wUU�ؓ��**+Bp��$�]~�+����<t<:l4��s]k�Y��HB7E�2Y��G���Ae�c?b�S��tc6=I$�q���Yicy������O�x�!��8�M������z�4y��6+B��:"���L�����`w������p����Om�Ő���E�N�̒���0m�����o�Af�`�F�2l�տ:���Z�kGuN��8O��6�̊[5m��lԾ�����'��3���\��������������
�ʩd,��\�~�8ǌG	J��
=ܙ��&���������j�N>oF'"P�����d4e�?I��c�� Q��hفА�d�!��p�#���YC�Y�US������S���O�T=�g�F�qO0��m���n�ռ������ќ?���K�w%��������KH��d)�j�4���2z��,� )�Hc\�����+Y &�Y-X����R2��͍�QZ��������=%�o-?��l�w���߉Q{\�<^'�M<��׻ύ7��;���A���>z�E�%#�X���á]�ʶ�E�62c�p�
����*��M�vۺ�1Ta��7���Me�qj�(���V��.�B2p��8�Ό����Hs���(����;>3�@A�H~�r�8;��xP���&J>Ԫ�<$��GU+Vz�ļ3F�C��*QZ�a���f���Zd�>zwe����af��ٳ������(!�ě�>����c�<V�d�<~3-rH�q�yb#k|+�n2La�����$'GY�w��a�}��8Ҟa��uƝE���֋Z8�u�c�}_n���_f�Q \"�J**+Bt���L;�����V��;gP�I'{�����j�o�]{�K���uʢ/�Ӳ����}$&�2�0 xlD�e*�| �'�\lp2��_�]�S�I�&8:6�5�W����})+@��3�kdQ-�b��Ϗ4���p�M9�����5P��'�&?G������V*��Ƙ�aFM��6d��r�h8o��-����5������SL?<ˎ4��:���Z�kGuN���~�V2���,�m�9�vn'˴��O��<s�a!<~��TV�9rT�u�8�	M����N���n��<$�af�����>HC�,��x���i!]������<}�����a��G"��Ǳ�������D�f	锃ц���t>H#�L?gC�7�]$Ѷm�Lg4v�&Mn�U9s7
-tG�L>ӊFq�q��n�8���Z�6p�	�4�|���	�[,K����**+Bz��P:&�kO�(t��Ζ�>�:�x�+�g?������m��M�߿����H͒�uE��m���~�BR�1�����}�� ��"���`,m:��0�"�n덍/��T��ٶ~��w�|ۇL�s_~`�+�1M%Q����aC�k�0!�-<=:6��g�PS�2��o:��oCn��kE��{^qO�8�V�N�:��֋Z8��g>��w�,����D�vKm6CD9u+�.���M�qS���5X�%�cj��q�u�*��uԻlh�h�R�,�n"�Ւ7��̵��}�����&�MN^�<���o�'#�~s�C�D�!�m"����
R�WVE��W�����Q"�U,\V�Qם�&�n�UKV���)W��=ʋ���X�Grkn�ӂ�k���[%LD߱5+6�����)�]�C�o���Up�f(�qE�ǧL�r��Q��G���-�F�dl�GL��e�h��>��h�&̅?45����tQ0~xp����5Tԩo_�����k��36�Nf�R0����:��e�y�w6�Q�CT�����XIv1�˫��W]��J�ՐΈ�"��I<�s��e�uy��6�c�C�J!e8Z�iտ:��֋Z8�u�>R�j�.K��n]�y�TTU(��M�t�����}�,$�˞�+��`�}���� l!Cs�U�����`�����C�]aI��5o�v["�KT�m�+��d���9ag�CoT����¸Pp� �Hu���#hIB�%q�̄��äg�[c��	�����>�P#���!Ҧ~r�]
���T�m�}ϩ_���[i�y�eכii����""#ȧT�E"#H��#��"<�6�l��!eB"0Ìʨ�2�F�GeWQ�yG�O6�#(�""#Σ�����4�Du�V�ֶ���ַH�G�DiF��XDR�H��"#��<�L)H��#�"<�#n#��4ˌ��0��U}��!�6a�0�)��u��qŭh��YkR֏6�#��"":�6����!B"��5�����Yr���q[_c�O�Tj����2⤠�,�Uu��w]��Yjp��u���rI�+�����T�6��U~�Q��DN��WmӤ��(�~�=���W�η�y?��7�T�"��y��z��_����-��2������ܛ���=e����Y�s��'�M~U*"����-�M��G��]U���s:�vU^��FgF)J'"U�H����e��} `%U}_Gwwwg}��P�U�}��ݝ�� @UW��.������  �	*��x<�c��/4��-խǖ�||x�ӄ8;'qEEEh����a,%�KD�������_a�(f�׹=g�4�>����z�$Ș�}���>�h���c���|�n�^���� �b��t�,�K��]�O|t`�|9t�h85��(�!o��{�=�3�4i�9��
�>�%�v����{�\�vW[&ʔe�]`6��$�r��(jٛ����;~��\
s��Q�c��(ӎ�-խǖ�Z�ǝQ��9���0��\�e��ħ��EUTURm�$t=N����C��!6�>�>�p�>�3��I�L8tt��:�q��O �I�c�L���JI*�@���zҘICXD���Ml6�pl9�M��|k��DM(��ʙ����qq��G�O������>r���Ô��w�p0��5OB9�:9yw��۪���Te��~G_��Z-h�Ω�8��;U��T�`�XD�,.���HE�&��u�`��,�p�Z\|C�HjPz�ojЍ�T���A�X�Qe�#3&Ye��oh���S]�M�(��5=���v�U�Ř\.���M��v}�N9�m��J�;�u�+�4Qͧ:�lN�Z�MM��F��S9��������sb���[�J>��8����xY��Y�o;8i��\��w�Z��$��O��s���ɓ�f�p�*�6]'G�?C0Ϊ44w�%<)�f_�B���u�ޟ{��HA�|���#"bq�
	ˁ�����4�-��RL���>��N�q�;(�jHZ��Z*�i���>������q�^~��a�g�[�-�A���i��GN0r댼Wаߞ0�D��4�WY~i�~GV��Z�kG^:#����<�Q�Q��Qj""b��u�����}���+�}^>�����ߏYp�|��S#!�������}�O��o���äm_l�����|/ӷ���x@$K�W�Ѡ�$|<~ǧ��U�G<c���$��bŤ�L1�È�'���+���|�p���ҏ���v��0���$,���*�Q�=t��:�+m�4Ce`�2�-�GV��Z�kG^uN��-c"i1)!#��clm���m��	[#���E�C�r�)�4�5����li2bM��(��K�����27�:ͺ0��7	��+&��=��>��!�bN;d�����<�u���_k�#�����Z��~��붝�24Q�ÇuUUC��3���r���Yc�gI��j�I���ö�=����`:Q��4��[�?:���Z�kG^uN��߷?!�^E�dF$���n������
J��6�`NV��\pg��z>s$���>l�Y���i����B�x�K	בb�{�|{���2�ZPǡ�IN��;4�6X���	��l{T�ώ�e`x��!_�Xo��DE:���9mp	6����E���Blx�r`�`{O49�^���a�>6�>��h��4A���X&K>0u���V����kG^yN��c�i�
.~�Ƅ�sJ�d�t��qx:#X�\���\ڟ&��#R㜲ܒ�e�ı[���w�O"����]�V.�Q�������U_U,��7ѷ\�z�����]:stD!��J=�]�Wհ��}[�>$=�3�����:�ǔ�yԨP�z1N�F)׺����/\�J�(��T�&����NRd����Y9�f��Mh0�ř�������V�>��w��}��!�Z6�����kY�j��_YXX|v|��ܨHB4��x(��!���ro$	!��f�BI(�����cP����6���eF|/�����"�	BIdn䛫djI �3!����B��^��Й:t��N�/[�a���6�2�:��έo-բ֎�xGG�}����E��c����6�Eh�VU�*�Y��x�Xr������rT���_����| L�&'E�w%���hC�k�����ƻ�6,x9aϠa�$�
(�����],�]�$�4T6�R�cY�Y>��I"�Z�[,��0�����������l8��߈W�i�tގR�x}�Xa����X�˭<�����[�E��<#��#��ކE��(��h��ޣMܑ��!M��EEEh�r�i�$�$YL�s�^N�x�1��i��Z|8�v����%��Oz6�>t�[4m��	���]i�E-��47�ѓM&�f�.T����>g�+���x�~x�>��S.2tc��do�Q�?Wf���o��0��z�V*�Ee����~g���l���HJ~P|l���2�O��-�強�Z:��pvG�Au+Re�ud���**-$B��M�����0��u��2Y���S�zc�[^R�`ڐy;����R���v�l���ϋ�
ƾ�w�܎�Hf0� �p9 vI���$d*�4O�<}�<�6[��;,�Í��O|Jc�II$��w��C��C�Х�(!��a�0�Hϕm:�m<ҖDR"#h��#�!��Dy�yǜGm��!BDFe�F��FDqG��yu�k��2�":��:���"0��!�DDy��akik[kZ�!�mF��i��R"#h��#�!FF�uyGG�i��F�aT���!�)�B0�2�Dm�GZq�q�q�"��ֶ����V�"#���6�B� $/�k���-������
�Ý��6����k7�=9y�vA��WP���p�t������ֻ�����|��)N*�%�D�k��ʪ�9S���X��q\�!9*R�u�f�]Qçg��?�>k$!۟����},)�N�?��g�/�tf����Ijf����NK�R�-��=/+���r�Ĝ��E�yT_�+��DL:F���}�Qvyv��i���k��<��-$�3�BJ�����E~�.�U���6z�wK��X���/�����C�<-�ù���t�)�	e���:n�Xm4��p|��n^���w�n��y�>r5(�������D��-���|=��kE�>n�����}��R���L���	���qw1M���R>t�����;o;_	�m��98�����Ѿ�E!{7�����wF샿�a�iD�ϓ��d�-����+��M�^[�i
��B�z�]5�%R4B8��R"6YR�#i@���D��nT(F�,�,c�Ȫ�"��*R�GS��R֤m���U˯���d��:�gբl�$N�*�t���v�*%:��~��پ�~7��� �
 *�������߾� 0	 *���wwwv�� �HUU_|������ @
�����rk�)\�r��yn�o-Ţ֎��q���a?GV5������w+��Q�,���%PǤ,���#��+H;)+EIȥh�Y,��HZ�'1�������"CH�,v�X�:!-{��q�Lu2,��G\Dc�c�P�nd�MZB�ԡeX����*(�"�AI�)hJ(���H;#��ʪ-L�U�ܔ���7 �1�EK2�d��EGjE,b����D��$��(�J�1��(FA"���"�E�)�f"�CM��[QL���)��d�2�$�%DF71
I$)1V�wZ;
"Q�Q��.I�ҪcV��R����NѭRT,��IHFңlE�k)iZ�#q�VUM�u�4W��\Ȓ��m ���!D�c[�cH��(A*���$ ����k��(R5(ݔvҠn���h��
�Q����R�R�J��A���hr2񺗗#���s-p�oh����TY��1C�*QX�3s�tu}R����`�r�5^2�B���j�+Rv�_R8xH�4�9�h�=��!�܇-F���{�����T�=���ul'n�y�H�|_�{��:?���/i�*�e���
wS��S��輅����NWC+�n�s��Y���p�g��p����XHCS���:v}	0��c���(ܝd=*I����
����/�	���"��L�̲�|f�������tt�|x�����3�ޑ���aÅqUyު�"c�C���2��*�T:W����$��U�r�XO5$��O,��߻ t3��u��>�_r��'�����y��Dyn�-帴Z�מS�2�i�Ռf�Y�W�0�UZ-��q-��F0���R{[8�,:b�F�Rvo����5S�9]�|Gc�&k��A��^�Q��I$*���po�+Yl��m���xx5��\>�h�`�2�M}�^oη�;�{wa�L�qW�Xٹ��2�-<$�Ӑ��y���~�I�������Á�G0f�Xo�0d�_		����:�1����}��Sm������-խ帴Z�מS�2���J��w�����-�!F��A�k�			(J��
�Ң�%HB�{;�Hks��v�t::d~�!�#c���Op�P?|�P�=Q	��ɳ�$:e���q�"$%L���&*^�I_�c*Y����ļ=-&�͍�@�>������߼���I�$�y�I���'>䌇�Cbd/Ъ�>}��c��!C��(�ƉC�Y}��#>l6��|a�`r|(���ncA���̿2�H�������-h�Ǆx�1g�B�ɤ�&�V��8p�BBBD�z<~���@��g���k��Pe�!-��cyQ�[
Ř^�zT��C��|���<x�=2��C�s]��j)���~+Q��z��|�Ǆ�<����W�j�V�:쐝6�t�}���`����
���6�>����@�����9��{<h��d�<�z�4�/̣K~Du�o-n"֎���!�!�޹I�dZLCGKM5n���Tǘsn(1��uQ�bᴤ�M���5�,#�bQ'q���Q��&	����å���O-B��Q�/����ʋ�X�nwY�sR�>PGO�]����i��)ߍ�M7���|�ڞV����:: ��핦N��d�������«�U ��>w��x���1��n��:~!i���Pl7�P|ctIa�����3��b�xЧC�Ü��Xߎf�r;ޭ(�Qd�-e~��a��������[���I��0!�ဳ��r�/���h>>sˬ�H"XYi�Dę$��h��|�'�L��Q���۩'Ãa��D4�-��H�����Z�E�y�<p�6v\�$�ȧ�Sa�l��VBBBX<��!�i�MLΜV�l:}	���+��o��v7�14�Z0��]�^ٲt=\��O�!���hod_>�H`y��VSF�I	���6Y�X�M�����<Y�m��^�UM����|q�*p������"@;
��dH�� �VJ����`hi��� ۑ��	C�p���$��#)vk6�;:����h�g6`�è���Z�E�y�<�)u�T��JA�Q45VDK��!!,�Iߋ�#���l�y�R�sS��$�����5d�����h:{�m8���������p��ʏi�����(6=�-����3�C��?�j�h�d��]˗A��sOG����޳�ƙn_���_�e�l�釚dbh�Q*���r8~�y�e�r�~9Q�+�70Lb�ܻ�C���'��4T�1���4h�
el���y�n#��Z�E�y�<�.�����Li�1���ղ�<А���fN����i�'�r�>�N���3�B����r4��,d[YW�߂o�^��ަW�xJ�[��2�X�ڔ?V~���A�u�C��IL�P��!��F��(9��>q��s.\N	{����&&�C������Ǳ��g�ۇ��ۃ"�ə���t\B�``�"�B�W�r8x�A�E6��t�Jyl�˭#�q����kG^yO8ʾ�c�����8�ճ��!�S��XQH41�S����s�Pb���q��lLĸ���8D�Q��4�[V�8��2kM��~_{p��T�R�Ug۫�못�����\^�v��v-�&]�ؔb�K2�����O$��Ump��tڔ�
���of���ܝ�;*b6��R���O�&���iĻ�[�:{��*.�p�����[��s��	e�tp�Μ�C���|�����F���l8j���tl>�Ί���f��!�.�ct�IV[	}�F�:IW	��<���Vx~�Q�(~���dr.^�����H7�<���A�4�����n�����2[����:`�mə"}�W��q�<�.2�KG��o-m�֎��q�7]©LSX��HHH�l��oBCYtd�#��x�xQC�)��>�L������%�5��,�����!�9�e[�{D$7r�I�&�t|�,,���|�v5�fC�C#�;u��C��z9�rl�X�Y��<H@�-{Ntm�����Z
�b�7��v|8hyO��֬�c�6��ǻӰ���F�Ï#ki���FT�DR"#h��#�!F�Dy�y�u�mS*B�!����L�*�H�#h�8�ʯ#�<�#��<�8�<��"<�:���#H��#���E:��#h��"�o6�-����[*BȤDF�GB#H�#��<����6����l��0�#
O�WЎ)��!F7U�m�G]q��Dya��"6����qkE�㍭�XB�!���B+����Zv��q��֎'7jm9�uHj�~���/{�7z�E�;��龚���D_��=jL���[�{���kj�B^���F�)U"]��|��k)jڝ��j�^���^Y]�.���n^�k*_.S.���K�����}*����.\��.���/)e�Ȉ��K���.�z�+'�U9�+:��/wJ����w�;e,�GNܭ;-ƻ������b���?{3/����  UU.�����  UU%�����|� 4  ����wwww}�0  *���.yO<�̼��-ŭo-m"֎�<#�~��!!!,.c'�J[Ik�n��<K�CFR�}����<P~�=1��J�?%�e��#��K����:o�P�48���?��}��I:Ƥ�%d+��ZF�,Iu�t���9��$$>���-��	��T��&C���}$�p��ֳ�uVYN�����$�_��rm�tKB���H	��[��'^��IV����^�B\�	>���o��T�l���y帵�孤Z�מS�2�1��Wꪪ�9񏾧��l,~6GcY=1���Y��D��u5�������իW7��SM�`({ю�I��}dɯ���=��e9Δ>��Cv�|;tmv�`n�!?ݞ�٧����HN:�n
h6a��CQ>��|br����?2[j~y���K~~qk[�Z-ţ�<��e�޹�gxg���<8+�S�I���R�����"�X��#��3�(���d�Du�1H�]�#7�$��C�i�J�*�YETi�4]ԜEVTE+������m��V���
�^:Q�AOln��%�/���v����:�����ǣ�H�^Y^����
��A������1�Q5��e��&�dk��Tf�ȅ{9}���B߇Ҏ�����ߨ���;Q(�G��*˘ӳ!��3T��0:��P��d�d�}C�a$!��ω��΄̲��ʞ~()�dr��4P�˞ǈ<w��۴�ZM4��zm_1-cp+f�K��[�?z��.��m�'�$	�Bm���������d���RȲv7�ѭ��Ó��Cs�fy�/��0a�i�n�����k�i���ɒ͙[O??8�����מSβ����[�3W/*�s7SX���$�HKs�����D$-3|3?��4k�1���~&�\�7HSec*����ͥ�vI4���I���B�I,tB�ѸQ����Ԍ$&��wभ�l`|d��Wv�,#��߼�9�� i���H[���vӁ�ٵ!��O�,&��	"3/��$�#��*�����ކZS.��/4���Z���x����N�����D�%DX\`2Fڒ��$�Ho��D���$��]��4��<����t���R�w����ɒ�>��f�;�h����	E��1w�FF@�4<(}�)�vI�A�j�F���_wټv�&�㥇kVrB���σgO߰�baZ�Hi���ٚ1/��w��t�E�#t��E��R�(y�:,:t�~$��{�s����}[2l��4��ŭo-h����u��:���U#ˍ��}I$B-��P�q�qpϏ�x��+�K����o�њ��KD5Rh��~��y��iu�׼��+fFܬ�:�ɒY⍴��&�9x>y�����B�m�'HԮ�9�s�
�e�j]ܗ&��Y]�����T;tW���0����I�#�c�`�*T�AӮ���;�8R�)$F�2�i�,K��f}��Dx�<e֝Dqk[�Z-Ǯ�Ω�y�#~��j�}1�4�F�� �n��[����^���� �,n�f�%f��0���)ZcM�P\�%�&q9��ޒI!��ߺo����կ]��9�n�+��l��n��z.���n��&.���4���`A�Q	��Q
�}���l�&!E�"f�]Ifc�l�v^�B6��#r3T,��� ��Zώf@k!��v�8�~�̝ ��h�ޜ�9�,����:((~�d��^%wN�nHpx�_�J�`���S.��ׇ�YM�C�\�?x��ٺLD�w��:]d��_��_��Ŝ����#��R9n����g�7u��Ђ�d,�>,aO�>~2��:�8��L����6ʜq�Yu���Ţ�[�������Dt���
�ҲC�$��2�bl��^�rl��O_C#񖣢����,��ߜ�bK�I����c����Vxx���C68���鉗{ᵄx�&�[و�a�?0����X�<��|}S�8��(�ѧ�$#	�ّ��0h�=��i^~�9���HJ:Q2Y�/4��q�E���y�:�/9� ��QcRH�z�Hf\�	3J�Y�V��I$}��l��pf���c:���r诸�٩43��Xd~r�3��II��63o?������~�୚�k䐲�8�]f�p�ѩ2��8�)
���2a;�ყ�'_(�d�s勞xz��C�^����Gr@�%�L����1�F�HB+G���P���%텖HG�#;!&�N��ŵ������/4��Ţ<���:|t�,U�]$�IwN�$�A�:GC�4d�4<��S�2�~3��Z%JHB��dw�'�����Vj�&�հJ����FMG�2P�I	$d�N�8<�˓��Y�i���wy���!�f���$e�lr�l�惶��Ƿ�FQ����0e�NƜ���UǶ�~�Ͽ��2�R��UJUQ����?�}����m?��\+��S��d�4�B��#����[��߱i)�-��""B( m�����ۦoZh���"-��DZ)Mi��KM���E1i�-4Am�4�S�&��Kh�Dť�E��&nh����1m4B�D�Mh�"h�" ��i� �:�D�4��4�MI!�E��4���"h���&s�6u��D�KKE�M4��M��-Z-"Zm4Z-&�-$�i%��IbIh$�Y&�&�Zm$�d�j-1E�DKC�'ZI$�m$�K$�I�E�x��&�Ii%�im,M��M"ZId�I&֒I	$�I&�6��I�$�I&�6��I!$�Id�I!$��I��mi$��ZI%��h�I,�I&�&�m%�I���Y,�m	$�$�K�%����M"M$�I�M��BI$$�Ki4�K%�I�K%�$�I	$��M"ZY$�i$��M$�X�m4�4��d�ii��K$��M"X�m	%��$�$�K&֒ZIih�i4�KI&�L�-,�&�4�M$��i���ZZ-����%�4���D�X�I����KM���Z[DI-6�D��h�I���4M-,�I6�YK$�ȚI���4���4I����H�և܉-5mi"�KMM�ZIh�id�id�,�K$��&�I��--"$��iE�� ���ȱ�d��D�&�I4�--"$���"KE���di��F��1m�FF��m�Y��3�4i��6F�#Y�F�f�b4�i��t�4�l�f�3F��6F��M�W�Û���iiac�����#LF�F�#[h�Ѭ#CF���٣Y���5�F����6�6F��FѴ���ۆ��A�#X��b44km�M��kf�m�@�3#[4k24�4l�6�F�dh���F�����kfF��#X����4��F�h�b5�26��LF�4�i�i�5�Ѧ�4�XѦ��m؍lѣh�Ѭ��4mY�&hY� ��l��B�h[4#hi���-�����Bd#B�B�[:�%$Hh4&�-�1d&��d&d#d�3&��Fɠ�C&�4�i�M0�ٓe�4�5���MM6�[l�lM�d�l�CMf&�CMfMm���M3M6M��5��4��CM6�L�XM3M�m5�M6�XMm�L�FM4d�e�5�M�XM14�i���FM��4[[d�[d�i��k2hɲ�hɬ&��2k	�&��bhɲm4�kdѹ�n&�h�q��MSe��F�M&��i��Y6ys8�hM&��i4�I��d�i��I�4�Mbi6I��M	��Mi�i��d��4�i�i��Bi4�&�&�i4&�I�5���M4M4�k&�i4&�d�I�5�I�4�I��"i��Y5���M&��l��i4�D�Mm4�I�aM�i4�I��MM4M4�&��Md�M&��i���i��Md�hD��"h�E�dYD"D�#-�DE�h�h�BȚ$Z,���ɢE�"hM��-DBE��D�!h�DYh�,��Ț$-�:�DHZ-�FDHZ-	�hZ2Ț4�dM-��&��4YBE�,��dZ,��BіDА�kF�$Z"CZ$-�"�!h�h�֋"h�&�!4B&��rl�&��4H�Z"�hDH�-��Z��BhY��"�i�D�h�hZ"2E�Ј�hZ-�$-����M
5�X�h�kh�h�F�7]q���pi�MhMM�i�CMhM�	�$&�Ѧ����4	�4i�MMh�Z&���4&�D��i�4i�Mh�F�,x��8hօ��дkFZ5�Z4�֍h�6Z"kKAi�DZb"i4�DZH��Dť��I��h�D�[n�;�����o�<���z�4������P?�� �2H��(I ����q�~����Ӛ�^�F��>����m��G?����x���ŀ
��5�|��8����g��?����9_����4g�C�_P������������c�Ͽ�kC�-�?o����q�1���������#��ˇ��~�a���o�lf?�8���~�|��>�y~�>���ߴ�7������|�a�������|�_���������^�lo�g�[�>�T�n��:�=Y�~<�A���|���`��9�?���))?��^"-4�~��:��?j����L!���~vS�.B@?~��q���� �_�,�ET.�iQTɦ3m���ܶl|5�� IE�E�EM��P$t����
��]��)����+	�����S�ލ�� ��Hle	1�7�9	f�lZ��j3f(Hm��#li������O� �~���_�8y鼿� �d����C��[�����'�|���?���χ���2}`��~�Ѻ�w��h�m����7D,��Xխ�x������#�q���!�{OTt����2�'�O������{�'M�G���羷��~K�z�^�6�d ���_�#<���G�������޻zl?��,|��f�l����m����~�_�?���X��S@G������K�c���ͷ�8ɱ�6#f�:�%
 ��+_�HO��x���<��l�}P6َaKO����2�D���iE`h%%��SG�����
����m�����L�8���f�������K�g����?��'�~��k�P���ZS�،��������?�?��߯������~�%���]g\7��O��_��N~];�������oɑS��?y�?�?��������P ?Q�c>[�e����������jj+)Jeb��2��ը�MYZ�YZ���55jڵjիVV�Z�jը��+SV���e�ڵjjjԬ�Z�Z�Z�QE�ejQME�[Vj�+j5mJ�YB��Օ���ڊV�Sj(+�
V(+�



5b�X��V+��B���b�X�V(Պ�b�X�V)X�V+�jj�b�X�V+j�b�X�Vڕ�F�Je�(Օ������R������eeb��J�QYY[VՔVԬ��E2��J+f�R��e�VQ[R�e(R�(R�++jV����)B�)MYJ�5m�++++++++)������++(VVP�����eeeeՕ��Օ��ճV+�
2��ej���Օ��Z��b�����Z��ej�j�Օ��S+eej�
��ejյj+(VP�L�[SS+P�VV�իjP����[QX��(VSQYZ���++(��eeej���Օ��V����YZ��ej�Պ�VVՔVQYEj�jյjڵeb�ՔVQ���+jV��Vթ��Vի��jڲ������VV���R�MZ���V���Ej�Z����
�b�P�P�V�+ڱX�V+Ք�6��6��)���b�MYB�b�MMX���L�AY�m[++b�E2�X�իj5eb���b�V�ղ�2�2�QZ���mL�P���V��[(SP��m[j�YB��+5mYYMZ�Q�QM[(VVj���MM�+j�e��jիSQEP�YEj�(յիR�իVj(V�Ԭ����(����B�lSSV��+SV++e1F���
�SVP�SPVV+��AX�PSjb�V+j�m[(+eb�X�Q�+��b�X�Q�������b�[+V+emX���+��b�Z�V+��l��J+Sjڅ55e��Z��J(ԭEe�S++VիjԬQB�ڊ����+j+SP��E2�ՊԢ��jj��Ee�VSV��SP�[V��[SSVVQB����P�2��+j)�P����������VV��+j���eemYB����jښ���mYYL���VP�V���YE5f���������
+(QAAXPP�f�V���Vm[j�څ2�X�V��ej�j+e�B���L�L���VՕ�e52����

ڶ�PV�V+b���(�Պ�b�X�V+�b�X�V+j+��b�YX�V+���b�X�VVՊ�b�X�V+�5b�ԭJ5mJe�(Օ��P�e)��J�+(�R�(R�+(QYYEmYEe�)�՚��(��R��mJ�ڲ��)��J�J(�j��ڕ���+jP�
V�VP������������Y[VVVV��+++������������VVVVP���[l��+SR��(�JjSS)YJ�)���s��ɽ�߇�ϐ6��c������zg����k�y�������L���c�TS���&c�+c��Ku�0��������_����a|%?Ք��p�A��}�&T6�����m���zy��ZϹ�{�o�yKj�������?����O�?����H��9�!ZA�|~y�ڧ������(@P�b?��	f@�3�����l֟�%w����O������?k��#��������?�*�20���I���ܑN$�@