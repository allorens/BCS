BZh91AY&SY�k-�/߀@qg���#� ����b@�h    ���Dh֛m�hJ)��Z�X�45��+M���l@�4jA� �J��)���`PQ�4i��Md��Fj�tjI]Z�fƑ)KX�k�5[Q�[)@��fhI���Z�Z�mK6�C6eVڢP���,5$�Uh�E/�t�klH� ��Tl���R�dj֚,��J�֚��R�md�2*e��&Ͷ��5��I�M�5��4Km�-�mFl�iZj����bn�zUZ���&�   �c}E��F�Wm]�k�MS��B)*wi]��Y�W]�ѣ)b.�l�p�*Ci�i���ݘR���=�[Z��
I%�l    6yl  {]�ڀ5����p��:��\.��m��u,�(r[�� ���pUR��w9� 4kB��8� ��sܢ�ƶ��l���	TZ��   ���x6 ���z�i�4�������w�j�
S���  ���CѪ�m��zPm/u���  �kǀ: ^��ڭI�6�E��jjQ��   �c�*@QW�<�]��oN��(
P=����A]O]^� �w���J��^���Р�� 
�@Y�]Ҕ$\���J$�H�ժ�5^ t<P������P�Ζ�PR�;����ʰ�P�r1Х()n��(
��u@i�Rn��� ���)�'L��Y���A66�2�� ����^r`:P�wS�
P�\)B�6�p����7P�Ke�((PT�7
 �F�:j�uM��҃��b�Pl٦cf�*���O na� ��NB@;� �C��� Tn:�� �� 4S����;Q��t� 6�;� �P#Ȫ͵*m�"�m��Z�ux h�z`���84 F �3 P�t )Ƭ �Aۭp(;v��h��d�ѶmkM�����2$$� hx 6�p �f�n�� Q��w@����TP�  ]u� �7 ��v�� ���)�f�[�KRґk� u� nkq��-��� �thP��P N�t�[� 8�@8�� n�p: }�    ��IQ!��2�*���0�`�	� Oi��(�  �� "x�
J�� h     �O��%J�`20	� �d�R	�jz2��M=L�Ę��M=��BbJP�%	��4�h  C,�sOL�gu��Ӯf�u�[J�_i^j�C�'���v���Q��.���N�7g����������Y@EO�@@U��WB`�_�q>���>�����U_~_�Е?�T E}���?����i��0'��̉��	��	�?s"}a�g� u�:ȟ����P�{`N�'Y�a��YS���� ��z�?��(��:ʝ`N��X���T�u���u�3
u�:ʝaN��YS����|e�'XS�)��"u�zȝe�'XOl�X����e�Y���P� zn�'XS�!���e�'Y���D�u���'X���:�e��Y�	���W����x`��XS���"u���u�:�a|3�P̡�� u�:�dN��:�dN�'Y�
u�:��aN��Y_,`N�'XS���D���eN�XG����)�� ��z�=`_l��Q���������/X �!��:�Y��� �(u�S��U0��`>���QG2�=ezȈ��A�
��Q���Y^� ��"�UG���Y��=dE:��u����S�TzȪu����Q��XN� =aU:ʠ��A���"� �*�A���dT|�*>�P���
�����US���X��=`zX���`zʝaN��Y�)�D�
u�:��a:ș�:�`N��Y���D�u�� u�zȜd��YS��T�嗬	�P�u�:��C���P�u�-0����Y���83�v���q>�M�����}̢s]��=W�yD���iC�6�3��+i�bLЉ���P�f^�d+�@�[�4��*����l�,+T��k#F�]���U �ȵ���F����2=V�W�h�`��,�qݣ�CX�U�YX�n�
�0�'ZӬfi�TعM�Ӷ�EACT8��U�zëW��;f�F��y%k���$�Cl�@������o�%����E��,��q��L�r���kD�pZi����(�ےm���x����.����h2܂�/f���u�.Ec�J�M��Y�Q�6JBҧ�0V��[ѧ��Z��S��"��=�ͻ�a����&�SC��2,v�'c{qo'̞��<���]�����e��, �&�
��ص��9c.*�)]Ͱ�ӹ�E,K,n5��� ��eK��y��=�\&��u(��g2�K٠L2�4C�!`�ʐ*���R����GlcK����o3+)�fi��@iI��0��=�p����E��:B�ZH'Z{u�J�>�=�䍤`Y����©R��
О�3J�2R��-@ða�<�N�%BY�Kp�du�w˅v��h���GI�1�q��mo��B��vwiՍ�P�X�]`��[����6�M��Mc�K�/����c���jVwQ����6kKp=�{��k�X�cB]�U[�}��Xg�Z4RX32j]�v]�]v�z��m�`j`�2� �ɰjcz�2X�u�����G�iKk�vؙji��ҵ��Gu�]�Ҽ�a��r��j��^ZI1�t2^�3��s�ة[Z���A{a@%%XB;yGum���[04K�`��S3R�ڿX���ƭa˥���G�"������Gpf��R��5�m�e�5�LU�sM	KKSE�)�8pdݭ�Ml��8��j��ܨ�RyG1b{u�r^���%(dT6�֔&̏d/qQjH��0*�`�jػ�)e�]w��.v�����D��<�hՠL*�{-f�l�`=e�[.��X�m��A��ܫ:%K	��v�����Stcb�C�e��M'X�m:�(�a̵����TĘ��{L)d�Mf��H�:5f��S0����X���=�������W��V��ki�$�N1Tͣ��&Z��H�R�y��&�Z;L�&��w���ef
չ+�Ab�X4EM���_5>���v�[@p:�rk֯��KR9퀣�p��M��-��J�а%[D��41F͡�SX�z�lH�![��[ �1�pD��x��{�����l��_+�Ӧu
6�O�T�>�{�:z;�ư��iU��t�����ZY�*��p8�p�r�z�0Y[�5��\�w\KW÷O�^�e���h<��0)��[�0G�SåM��A��	4��Ҭ�ٴ֕.�hV�eZEb���VҺ�j����,��7d×D���v̰���B2J�,��y�RO��{��N��m�^,֊�Ǝ*���qS�����Y�`&���z;�!&'�GY.Q�"�6��)j2kO#,�@���̙Y&n�lMY��հ�Xp kF��K4��ZR=���cA3uh�K�i�c���Ǜ�FH�AT��g(���On���f�q{��Ջ�YHV�U�WnyM��S���"̲�e�.F@0 *�F˥1k"��5V�f\��nU`�����ڎ���m�f�)ݖ���A+lmݼa�	�����ae�lC*OTŲ��#��H��0����M��l<��s�آf�dR�sЀ�i.҅
��+�m.ѵ�e,�d`��2%�X��̽�S�IP����{k>E��-��-�[l�@�Y���$����\UX��F����
x�g*ś;p�F��
I��[�b��[Vv�#R��d8�S�eP*9V)�V�%x)���o1f`R�V�T^�����s2I�E�,��)᭢4���n�n�v�e�J.#�O�j$����M'�FЬy� ��2Z	ҵ6��]
��t֕J*O6�Ly����/-1e��b��JPd��s*^ ] ��N ���� )�j$�,Ҿm�0���s�ݜ�4��Y�95+�ț��.�Iv���ٌ����F$�'u�����$�Ÿvh�&�l���b����1-ч��4K����:ݻ&�@cT+���b�;
!��[LY���[��j��G�J�BV����7x���q�|��e,[@#k�7˴����b�㻎Q"�+�j���ͼ
��|�'�)���Yf�r>a-��XEi�6�CVG�;#i�vc��2U3lM�wU��lf�m7��b]�oh���P�7kF�X��S �źf���^����cs*�bνU���m*�MF&ګ�7dS)����ֹ4(��v��4d���B^!f[,l�1<{/���7�*�m�ɍ(OA�4-^<��9�oFX��*c%+�,%��ҽ�+���jH�vP�ۼN�i��̢��`����a8�a*�,yx�7b���T��!p��)l٘�R�++h���woJ:K���ȒV�e�(�Y�E����=�(�Zkq��wXK�T�B|r1�֣�<���.��J������Q��<�7Et삫f����AcCi��⥗�M�.�;��Z7z��E�V����n�j�)d��,�b]��ը ��)u��c4�qIC*���3��K�*��[���ط��n�B�L�5��]����tT�d��Nd�����b�̗I��&�N������7B�*�:��8Q�3�w�O(\��\t#�:)Lٰ�h�kr]1M��R[����p0GA�Q��b.�uڲ��Ow�[�̂��.K��0�&��+4�0�������h೪�s(&y�C��*|u aA�TE݋Т�Xk;�:V�S�eJp˳�M�J\Ǘ�M��diQ=O� ��L�[�&�l7�޽���wZ{hѲ��[��
b([ww˺Q�#e8��qf��WFV��顪%�����9�b�B�5Z��U���q�W�����WE�n�'YN*g �U�q�Ҧ��12�i����*@��oXǃ7�Cn�륻1�S^��6V�{Y�*�Jo���&fW���l2����p�N;fb��I��44��S�Ѭ����ܚ���,�Tسt���a�yR����71��� ��x�vr�,b���v\U�-�z�
��-ҹ�Y��@~e��sZ.�S-��U�G��v6��V�ko��0�Fc�)�t��Ak�W2����1��x�pG4֬��[NM���6#�	�l��`<�m�#`[f�3ql�� 
ՙ�5�*5i�}��|�iu�;Z,�0F�Ҍ����O2���f��ޠ͛�a;׺ ��l��*�Y�����*:l<Nv�2	��WM)��D�kƙ���-[yN�@X���-�9m6�Ubpdڳ�C+p`v�b��ĵ�iӟ�4m9Y���!��,,�1^�*�D���d�wn0��$M��^�5�����0BWHҦ���썺sj����(��
�iZ�L\�1�v������D�"���ٗ��kNK�gM�pw�x\�X����)�'	�R����2ڇ��x��uB��&�/��z�q{�>��S/i^���(�]5��7� �݅1�BE�d�С��F-Ҹ6ix���NKv��;%��"�0�m,:U�;�l�ږ�;ܖ3bf�l�
p�$� ,[ݺ�N��Al�~�V$�J�DQ��1����Kg1���$�f'5$]o�m3�y����OV�<v�K����OA�M���L�2�D�3��qY���#رͭj��0CV�����Xo3O��+#M֫CskmPh��N�Z���`�����\��˺H�w���H���nߣ��j�x�lI̶���G �k����4=�[hf԰���F����*���f[�)�=���8�n��Vt�#�C6k6�v�J+bX�Gw,Id��qXxCG,� �Lh�Lh:�ֺ����sg��R�O&����C�D�ָ�]���Cʧy��T� G���˹/k�V���.�*!M�[@[�i�,�(���x0`^k1��M*K�i�l�R9b����{�66�j^��*Q״I���r�"&V�fb ��,��[�u��쫢ԧ��F̹WB�[fD��(d������Ձ�%���YՕ�C`^��R2	z5߲�nÒ����tD]��$�ngs�ޖ�`�C!RH!�)= A�i�H���D���k?
U�JCt�(D!���m[9�M��yn��pH�ͧ�*�Qij�	��@�;Wژ�J��n2M���CK%����L�K*�������0k9j�S�q�]���cJ�m-5��dcr��b�w�Z�].f��A��\�X]�V�j�EhA;�D9E�ӱ�����F�G3-A k�pAA�Z��D�)̤9.9�S������1'`Vv�V�F��b��m�u��T���&.���頜��f�Ǒ�����e̓)PQ�ZA�Q�V�Mɔ�f�jifw�,�&(cT0�ĭ*'����r�VK��"���V44Sլ���R�64W�;E�՚�m��
%w=�\w�@�� ef�|V�.�$Xvެ{����hܘ6ein�U��c�VFŵ�1iʞeђ�hVɗ�IcqCIT�EL�{[{+]� eҼ���-S��"���쭻��������J�:��,�a���	�nhY����[�X��qӷ3.����t����Dr�&n<6v�"�CQ'3vB+5[{�V_➤%	�����i�ȣ��t��L��5�*���h&/-��XEGkv�h�̸U��cZ)Ӂ���̸�����כ�.Y�X�����ޡ��qB19�'h�5粏K��
�+��KH;;5���.f�v)�G-һR�M�Qu$ř�%#̂���V�حU�^(�Eiz�R�߁Ƽ@�y7i�+ů5_���:�J]�B�O��x���g.[CX�Ճ{u�.ж�$X�$<6�^4���C}fz[Y=���8���B�2���kS
��q��j�c�+&1�P���B��ů�9Y�)�76�)�5�$�87jb.����Þ�	w���oU5�n�P^ٗN�[��$�	a`��<z��N�)V�8��c���%Yyj�ї6[ZɉLҍ�d����$n�r��sj��Iyn�+׻z-�MӦ�f�vū������݊�����$5�������Y� ��K�|iKS]�cpʕ�9.��ԣ�R<� iS �3kK+^b�Ʋ�[�ȫ66�ZF�$+��DDMTnK��6��ۿm5�d{��m6M<ɥ�����1cuz֊ Q�71��۩o4��fQN�������@�U1�2R!�S����;���32�r��NR�WU��^��N�~g^�Ȇ�]\�k!ص'�+hbl��"F1����6�&�tߒZ�YB�IX�˚�WqXORp�/c̣�Xc2+�Bi��-�Cٱ��pȃ�$#kf�ǁ�b�YV����1uh�6{{��r�O��^�ĝ����j2�thQ�y�b��n2�W��M�72�,��v/�e</���$�Qe�6��n_4.��{tY�Ճ@�QZ4�62n=Y�^�58vnʛY3�F$.�m�Z�3RX����0sdq�ܭح�n��ƪ�vy7CQ`�;KiF�F%,̹KCI5�B�l���V�;s	�g;X6���ff�P�ѽ44��+\������'�63�C�-KqJ�m�]����7j3���[�0$h4ݍL�fL�� cҶX�C1�U2�q���ۛ��c����5��GRic'i�Av��9@jzw���V�4QC+]G���m��4%]Br�#Y�x��� F�l�CG]���ۧ�omz�r�x�̭P��v�'YF�v9� p�]���X��ݼ1�����T��+(Җ��Y��:�@�P�wL�
ә��JҬ� ֪]b	z�c�T�F�amo��O$V��6�IUN0D�H�'�{Zm�e�[����lLaX����#��T�*�Ң׌��Ѫ�MA�AA��a�A
L��É�ܳ�w0���ܐ� 3-�(7���ywY
�57^�̤����Ew��	��Gx0�G,��te�Y�hbNf4�s &�wVF�{;v)Gdj�yS49{�����e�K�$�6@Ee^�%@[��4�b��lz��M�!'�J�ј7���y��y����-�J`g�(���=ǯ7�&s��+�
�"4j�N��Λ��u@���J��"n޻� ��WE�$�lx��v�W��r��I�Qf
�V�,7������6�jPJؕa�S&V�@<���A��I��z`�hH��+nZ֋��9�-XHh�z�h�"�Y���'z��5�Q��;Z��I5G��d�:�yJӕ�U��.Es,�#�V45'�Cv�F���mcN��\����N�QE,�AM�HK��4�(�z�	u6��Uy�惣3C4����/H�8��!�aY�ݟ�Z�H�	&ի!���D�/	���k�r����xv�۾���g�}Zv ��-�FBPd�;�ŭ&%_P������{��L� !@�i�� b  ���lbI(�6Ww[udbp��흶�AhD,
��bI+X)i�KA��'j�_'�R<��D,���i.�����[Fc�tC���|T7)Rz[:�����C�$�t�[�e��`.�L��m�K�8���9֑�]C�43K�Isv��披Uh��! �q�Xv��,���B�� LD�	d��g(�O�!d�:�'4�B#H��1�B�u	��,4t�A�Ȟ����ʕ}�l�0���Hb��h�$kzz�ʫ���K���LÍ�� ��K���
Ư�S������I$�I$�I$�IPC:9V��fb�)\N��<T`V\���h5.�7��Y�H�wv��؛Υ�I��u˴S�L��.� �HQuz���X��q�	{�A��`9]G6�,=����M ��޽�e��}j���)��}}l��*�v&�]u����R�2��m�mi�:�S����*�M���O5FE��6P�X(������Ymt�T��+f��76�I'mc�0��)�m�-X�4�ʑ�e�r�=�1��I��p�z�z'���H��7rc��.���/��P�&�*$���-}l�������o��o4~��2\���ƪ�Έ���K�[�N�(���>�6�j<!���/ ���5�Xnî�q�4��ݘ�&' r�\�3)��f҄�2���)6����N��y�ݗ�e;���ɤ�uecKy��307w9⊒2���״�zűe�C1zV��U��9:P���Ka�+�/f���1{н��p��7�
��S�ym\.a�꼝c9�q�R8���%k�A+-=�M�-%�H*޴\�l���@Ñ��G�.��W[��&o�G1��oƒ�i�ػ
���m�Y@�P���yi-aVD�8�iɕxz�m�ɡme�MfVkHа��ls�6H�'.I!�F�Nʲu�xg�VBгJ�5	7.��H�9�e���aJ^��}��S5̀݉v<��5����0)Ժ�d��Φ���w4�13&q���G|��ʧ�׬���umN��n���𡮝_J2�[V��wk)�ׅ��k�2��Fv)��^����o��Gk�4��i�-�)b�јҧ�t�R�̛!Y\��0��l���:��'8�M*[�'�k�V���Z��w:t�P\�+n�J�N�*�u&r��蔐Mg $ö�û��ђj	�r��49��"����S	`]��w�"�"j	�ti�dBLw׸^]���;e��+8�Z�R�Epsv�p4�*ս�ܖ�m��;��3)�ʂ�v4�|f��.� �oV�q���� �ٙ���Ԩ5��c0c����w�ܚ	b\������	�/�w]8+;6�s�a엘�i׵�
`�}}�.��k���L��GO:�db��+5�*j�����B39c�6]2N�3���ޭXL썳D��7N��Mh@d��	v��56���Ք��-]}V���МY���%�=D�b�T��QŹ�����ڂ[�Q:��W��svCb^&lkv"�7zҚ��K�����I����v4��K2ǞZ-�Y�D,hS��YF��s2fWm�����!��l��g/�n�ܫ�$��!��B���d�t�`#;��{�f�1a��$�m�a����"-v]��w ������"��yb'�^��y�)��b�7k��ڣ�ul���'��٫�(�E_ܞ��O䒱j�*;��gon�f	�3%��h��k���!�%��3��\.>C7,��*wp���g���`b1����	�3W8n�Yu���E�Ԏ-�����x.��@��$���H�XH�"s�����m����c9'c`��Ͷ��\��gf8;��˩(��êe��~�e��-�a��/&���W3��M6�U�X�Y�9�lT��iK}X]p��nd�+�z8��(HU�\l�Vo5"B����b]����윙w��]�튊�u���5���� �7��	X�2���'��66�uI�-�7�(dM�ET�tẐf\��Y�Ү�[��{W���p�FV�	�3Vk�̩ݓ�9Wmf+�6��;�d�E.c�s���6-e�����a��Å�W��A��(_3Jӈ�p�0}����f3:�:
�ͦ���nY;��(YE;tt;\���
�N���̦�t���X��y��F�<C/�z8O\�.�`�r̬|^ ���9ˬ��|��;Y��f}o��Գ2ޔ3�i����� 7���)́u`L;�$�x�s��|1qw��U�iV���U�5��)�ql�ْm
&�U��6�e���&p[�����s-]B)���az��Ve`�b�9�q���%R��R3X��]�֨#��זM��2��R�i��Ȯ�ޒ�R��-J�^�4$�a;(f�#�ɦW�]�{�EL�YX�C�9Elx�C�Y�GI�Z���U�2��PV��q.I��1�`ax�k����׏bˇvf���(,�o�LJ�;eQ�����^�3\�y-q���N�q�(+A�e��v�N)����̅u�N���%�rw/U���ت,���Md,��B׉���j�%$2Օ�fH�l���Zߟw{���!o�[85�r��Τ�4�6�Q�<�8��)�|���*59�R|���l��n��w�T��o&J{"�6M���0Pe������anv�����X����r}���Ey��:�N�\XٵT��w-��:'�	,#�4���B�0p����y����b�af�i*\�AX�j�5+�q�V���;z�^'A�� �k��P�R��\/+5���@5�$7�E��LY�g3y��L�冁����kNh.*w�+�(�	u�#��A�dR��YPS��4��͞K��a�W�/I�6+$��k�����keL��ŗϵ�
�|�м(:�A�p/���eU��%;�(�=�9X1�6Yff�i.�cCe����%�:��$�[����^҇&.�w;e���!��66Sp�cj�NGK�gR�K�!�s:aT/[�n��!U����J��jooyF����.&Ӱ�������KjZ�l��xVc��y��Qr��+�oi(ޙ�"��l=�i�Y��Vn��s� u��IO�QD��(EtQ������.Hv`.����T��0�{H����9�E���/V�n	"�D�g:k����$w.]|�eOZiX�YF�vM�Bgbs���Q]AZz;*����
]@�+��c�X��6��7��\����w��ԕ̌p�e̡OFfP)�r��Wg����7�	�&��T=�tǶqT&�t�5PYٴA62�M�z�[�%K̹ޮ�i7ڥ�vS��,6�wgi���bA��Q4�7��f�%�ս_p�mt�:����He����gZ��
WeG��@j�`�s��Qb�)�����;IC'>����;]2�ڕ�X���ͣ%ؐu�v��lL�*��!�N̾��Ub{����r�j.xzT7����-��̏;��8�䐭���Z�.�Y�vy.;�zѹx��m3�5QV�7���@���Ž܁m�6;��������|���]fMC�%�Ȳ�HB�Qk�o8�2����t��9�۫�é`^k(|/+ݨ���[kU��B�y�\Ķp��4^�kqn靪�t��2Cx�L�3���c�ؒ��q�v�zތ2O��n�9.n\1t�j��@�]ސ�sd�AV6i4��7�w64����j�mN�|�S�Zy8�uv�HӬ	_c�X^��<H5�l�uf6=B�H]9��:d�M��$�Zl����O�х@ocN�mr<V�0��Z�S�e�s�7x�ZmV����[@�*�U�q��#�����먺�©YCc�B���8�-}cL��b�:��2�zo�f�V�͎��e�D�p����᷺.1�\��:Vp�8Ç��Vx�A��V���6i�5�v�by�8�m
�}��m;\���3Y�Dqnm�ѓq�ݗ6��Ex6f:c�X��RTQU:��sL�o�2I}�vm�D�3,�C��S��G��V�w�Vr��U^��Ju���>�
Jiy��*�y�9*�n���KnӺ_3Ǘ��/��%MȻ�@a�Y$v^w5�M�����B*��at�d}Ha:!�T2�ѷ�� ��ZKv��܇F����4ZV�(�B4&س{�%�� �l��d����^�E��ox#�U�ʗh�L�]�)܉�C����ٗ�����aF�
�_E�]X����7PU�m+0�4;�4��]lYz�t���� �=ޮ��Z&�vF����@Ӡ������x�&e�;"G�j\���&3zˏN2N�Ji�ڐ�
��M���m;}���@�MM��]�ow^����!����Um�9����{�*I��g:C������[�V�	�a�o;
H�]g1�\��n����ddյ]uX<�3�A�g8nBf�H���L틛7��L�mAAe&�݇�a�d#L�S^�0�M��Mo�K���:{y�ft���r�.�zݫsq���)_;�f������o鋖"%jЗ
�ʔ�5=á��b��E���X�7�TJ��.��%�X᥃s3V>�a�Xl�����3��-sf��s���h�,yF:�����gSDd�#�P6��+�;��|��"&����f�1�W�M�����Ѥ���I]50W�����w��oj+ZXnr��%��]�����U�!�;��2�4ԉ��'B�I�˓2�3�N�������m��J)]ұ�֋b���7�{��ks6��хt��[�-u�YDcSڍt�؈����pӰ�wC��(OhƖ	6�^s�a��7&�]���{Y�6��ܸ�s;��S���tȔc�B��pJ+*cs]��+Qܽ�
[)��G@N�<����e��uzN�e�;ia�՞ޛ�u؇2tQ�mn(����c\�@p���GRR�K_#e��cT��Ns�[*JC3���j��J�v�d�D�3�jݦ���.<�8�"��K��:�5M��$ڏ:k$F�j��y����uoR�uV�Uj�un��[�5E۴9u�V-ݠ�>�c}��k���Uc&�H��Sz�V��@�Q:�#�ޡ���۰R�W��l�qYf�U���,WQQr�:]66�Xk(���!����y�YG �&3�F���m�������J�@���C
	���%�,,3P���:�r���P�3���n�%��8VR�3�s�v��ײ���hU��h?C^�/p�a�����K⫪��Pn��w���!��#�A:�*޷�����\{c�C��W��; ӽӶ���,�F��CM>B�(�]�u)�v)b� xl�+8����8ukձ���Ͳ�u�m��y�#�����m����e�,l���(�죖����Oh,��&��)����✹:�s)���
/Uq�G9�%���n<ţ�GHV~,c��3WX{%�|p�۔/���A����r���;�X�rC#̜-qK^�A��0��Z4��Gx�&[�w�Cbh�������N�����e�&�8+������{�J����-���/��P#�vW3���+=6t��)JhwK�*�L��ؗ��
׺D��r��5��>�w��a+�xt��y�SP�}tu&��YR�C�4�Lv�*��dڬ�)�n�U�~�L�hL�;�y�S���D�`���®�Ɖ��5u���[������1{��,t����.�g���g���h�]`�Cr������(�� o��(=���GH�X�6��k�[���}N�����a�{^♻t��'Rm$9�}0�c�aT��f���m_]�9W��5-�tcw�%�i*�yȹB��qpG���v����]����#Q�j�@3;;$�4�C�Ò��@ZB9��NY=��hN�ë�͗`���T �;��c}GV�a�r�-Q��P��ڻv3�e[���N,l\Ю5�v_+$*�%Ƈ2�j���&T�AU��府� =�d�tt���i��i�C���z���c:v(�r�`��jK��2v�u}���$hh8l�@�:��v�e)wOE#�`���o��i�f�Ol �Ab�ZX�,�]C�P��޸P��d��quI�\����)-&S�m�|��h'�[��a���ߟf�0jX�6��9z:��ýҨ�������ŀc�{)�[ �}���:h�VL��^m볷z� r�F���(�6L\��,ۧ.]<�tƫ4�!mf1��nX,�8��'cT��K��
J�ȴMW4A�l����.�']c�=�����t�_NN9�>{u�\UՊ*�n-u��`�G��'G���Ȓv�閃N��8���������oz%��Z�`��A��骺�͆�u�Ƣ�N�*31��D���n�eU��0ۖ9M�T�e��*�\2f�m�����7-��2.�e��8�t,�A����ƈ�X�}R�ʹw��Uo/K���1�0��8�/M�/^�r���a�������2ٴ���y�.���dd�í#�̧��A����B�cx��̶�g�ׯʑ�f'�D�W���\-�ڌm.�v�\ѯL'�p.��J��N�e�w��}��v��d�Y�p[)��1��	R�l�sx�H�VS���^��zS(^��vm롽l�ӎ����k@���R�Uy�I(V.�7����H����˧��D&=�d�1R`�M��0b/�[�d�C�a'&�%[C��d��p`��������dF�"j�ˎ�a��g;)M��)�1�r�5"��d���u�㛽�	A3{+��ww�q����H�}��}�������K��;'��NI�}B�{�B���=���])��r���>`�$_R0���O��'Ϟ��%��y��̏��Bz��m��>�O�ri��3�+��T�RQ�D^l�*���� �6ap'�ߍ�'�� �"�?O�F��┃]
���)fEgY���J�V�e�&���a�.'�ġ��v�r�kc����CR�ΜO(��us�^V=���9J^'�mt9��� ��zw{%9;�v�-C�6��ͪ��2�Ylb�טK��k�lc\���ȳQSR9ػq�	hC���l\�-
	Ѱ���M�r�7��*Wr�y]��tc=�\�+
.>Y���
���t\�ț��@͛u�A�EfvWb����D�n����h�7\���.�{{�)���֤Q��I���z�E�F�l]w�;�HOZ1��hb�
��:̖�r��U��y2��d^�E�[�j��)�l^�	�Lc����%ǖٲ�ͭ�_�Y�|���5)����*�;w��[�v����pojUyʵ��DsnY�b�)��u��B��r�k�aǇ̆ɦ����i��vd�N�Â=37kvݱY���l� ⮚(M�0�3�m*}���:���gs�}��_>f؈h3[+��<�����Szȩm{R�uwz.Ӌv̶�X�cɴ�B�	�QH�hcy�B��B.��Gj/��Gt�o�c�I0xALVͮ��zyl͇L�g��	��oT[�6��qt�t�
����nn�;�'M����]�-Y��,��el0/�rS9�Z �]C+���ދ����-J&�S�|v۰s}���<�4�WǗ'�LV.y�e�5�e �H�*W��n��[���%>�.���r��4������D��Y��X��:iI��Y�"�T�D��bJ�u̉dI�&����ؖee�jw�Y_-�����{s��h�ʃq�Y6�
T|����,�=b�0o>w���+l1���씚��c�w����p%N_g:У�l�(�"Y���j��%�Krޥ��_��V��9�4\)�g8�*h-Q�(d�`��w�tZTj��\jګ��e��Z��1���3�t��J`�i�ҕ�u�$xa��Q8L��h��I�K���'1f#�dUc�������J�6D���ܖQ
Pu�L�-n,����r��M��+�@����۹�'#����V[�
�rZ�]w�r�U��;��4�f���u���Dp�o1c��EvJ����o
��omq<@�wbzp{5�U�	��ڭyu��oIq]M�f�V��x,�|��&��q��b-���Ly'>�Z�XL���F�TwQ5'�b�ӹ��QVV�8�]u̺:��Ed�K��k��r�m�6ԃt+AZl���v����4��ew��y]ͻ>L�0I�;/y��w�.�C2oPV����kG_l�o��'n����S�mZC����(�U�.O�q�s�������ԭ8b��R�����c�,��s�A�$T�|igN#�c.�\�'$G�棑oh�dέ�[����T[��l8��g��t��Ww����P����uĺ�nQ�GQ@������t���v )��U7u��g�c<�W�|�JViao�;-��Tr�ޘc�kQ���Ct\L�Q���J�yY4Ą��z�戺aVlksl5%�z��e���=�FAV�vl��Ho�r(�yb983^�&���F�U[ˊnͨ �X�a��$f9�a�y���J�Z�OJ�-w9֥��-ns�>�L�#U��c��P�G���������wE尦���k�"u��\��*S�v�\�f���Ŗ��Nꫂ2X�[�7����xBD@-퇄�@5�T2�Uw�5j�.�pdpڝ�ڔ�F�b�78��E�{ n�lܚ�v�a��Z2��{}ղ��4�����r �Ͱz�m��R�j�R2� �)��0�^Xc�2��:����iH�q�X�Վ���tfܕ00�]��У��޺W�~n���;pXW�h"�FN��!�F�ń�LD�h�i���KD�����	���`*招���ۯs��Z d���95;ȝ�܌B^c�EZ�JA���	N3Q
*�]f@�K��$��%8�'�R"�0��sv�l�f���]���Υ��mRu��>��t"\�.�7���WQY�!�z�,�3��;������oek���rp��6v��0B&�n���!�X��d���R����^c�t���
��WS{�]H����6c�vN��V1�ղnL8`�<om`^$I[0
]���f�����$uYKH��z�n�tv�tS.�$�VRL]X�A��w�^��o1Kā���Ç�'��LPCۻY*酄>�J!�L�\E�����ݦ����Ƞg�͒R��Cz2f��;����4����5ǃ�V�W,g9���Lͳ�B�{g�n"&�92/�\ö�N}�5�4v���+l*���{M��1ٮ,<Q��D��]I�-�Ĵl8u����
�I�"��/�]:] �Su1��&=�,+X�1Ի:2��\�,s�r�x���:3Y2\�U��m֊�td�(-dۚʆ�
���R�7e���u^m�n��&r��Uw�;ʽ�M����}�q�]���{^+Y-@���f��]*[�/sI u[��b����h,�J�:.Vc!��6#���Q���������<}�0���L�}��edf��t:a��wĕn���xVb�]G�v���	ܹ�n��A��_����s^ܹ��������Nn*�e��؝h<��{:cP�Y�3�O���ls/��ڳه�#	���G����z�ꚰǝCUcat#�݃ge*��t�
� ��Y�F�\��Vh��94e*�i8�;�C����YK�%MьQt��n-eI�>�P�ྛ��8�n�p�:p���X�m��[v�!�@�8l�{�1gI�2kSՐ$h1V̶�%�m�|̬)��u/%ޞ�X:�Mm��q���)O��Xy�\\ň�h�í����.�m|��:��t~�%=��v��Ԋ}X�<i��D��1����7Yt���L� �]6��:Vc`�"ɜ��bSct􋫚(Akz�mL6�����[M� 8���3�`�x�4�!**P�Q�{VUʎmmf����O(8\�7L��'�})���q��EՅ��֕�j�D�M�LP�����3h̦����w:XkF�X"2U�9��1�]i��&������g/�"��
p�&Nd]\bޘ95�����EV�!��������>9��]-0Nh<�.���VmF�Pf,�n=��z�����ɡ���>u�* ��u�	�Ɂ���2v��N��f��܆l��OU,��8�c��}V�%�w|�`�ӭ���%�,�h��(-k
��GY��J�U�K��AsC�����v^�[���Tfҗb]d����N���'qL�e;��W���qj�m\2Wp�T�<G3V�/�}�"�yf���B���t q���8n�VD��zj�s�+�vʖ�ک�M7&�OcZn�����}�'�*�O��Vv�*��yS��ﶸb�b�+m��N��\-��T"��EX�b"'w9>�!E���z��|�uR]bݜh9-0��[Tv�=@:��x����L+F�IK^Zu7��Ы�87�,ֵ]��-���lm�n�c�|
�ZCek{�CR5k6d��&(9��6�5�,5R#����P�a�}׉�Z�Ft��N���}O�+�V�dA}��f�M�ק�:y�,e�Ī�_CY�{�$��u�6s{��d|�9�V�':�X��i�xN���vm[��\T�kյ윞s���<�%,���+y�˰YB����-Ǵ67j)Ґ#Ww�Me��I3 N�K��g��Os�F������v����Z�	er:l���a�;��$9�_sy���ZY�Pn2�1��{	� +�q���u�}Z�Q�5E�Y�X&��&��$�c8"rI�7����j�n���CJ��G��F7q80R�naz�4K����zu���f^ݰK��lvRfE�VZcU507F)�v�eC���.@�QT6f��b��x8L֦N������8V`ӫ4u�ݖt ��S���ۂgb�Û4f� ewĺ/Ckc��D�c)��Kw�E�n��ջ/`�X�L�p��d�I���hHGK��N=�z��� I����jه�51���4 ���ɗ��N1�܋V֬$X�K�d=�j	�Ӌb�7�-\x:�{Q$���F
gD��L/Z��:�P�r̎c�ϴqhb.���MA
��ղ<�+�"/���-)��n�>��ǅ6��%��7p)�9VMh2��M�/^���q����U�ܭ�-���26�����7�#s��O�1Yz��l`+vA+{����C�,�/�\q^7o�c��Gȧ�^�ǔ�gӀ�櫱�xܱ6�}k��F���	v�u�}&�Td�A�x��(��Yt��c<���H9]�:U>��g)���fR�2��i��gu������W\�DXԧ^��C�Z;��=h�%&:-�4���6��dM�»�`���7�����}|�3\Y�;�IK�s_]s�#a�ݙ2�r�c+Fa��W,D���m�:�֣]��� �k�����)"W-��o���g%�@7[*��n�Qh�w����y�F��CrT���e��s{\L�إ�S��R��X�+cW�+{y�"C�e�8Ŝ�k �^��_Q�w�q�9M���9��V��s�o�܉ۋ���Qf�b�W;��_�c�wb��O5�v�^�4wSpl=ʐoMk�(�I���r��':�\�k�H���4�5�62]�E ��yG�z;uF:�qW(Fj�*ٖv��y�r>�r����(о�p��{Qe>�[��G|y�q��W:��&l62��hR�'��Ԫ�`��6���I����'�j���x��q2�E�L0�;c�7�є�w[`�ow�VOt^ :-^T���V�imԤ���w�����0���l���A+�!��U��V�iN:ɺc�#�ق�%,��(fr�٨#�h�G��Q<�%�-F���NTȶ;:�=s6�E��Jo�����V��l�:�]5,	 �E�u�c�Ow>�qk�õ_F�\${�XΝi�ñˊW����Gt�I�9����+�:���]�qw2�啷��s �Sj��D���k,�$�&s�y�U@�N&�ν��`�};W�g�=A
CˌI�ǋW[K8�#j���o��F��Su}�ɜ�rݲei�ђ��Y�����>�4�ʏ�p��`��骰�]�iY4N������7ڞ�����|�^�3S'�.��MPB���V�l(�M�){t!8���HMI�'*�U��]M��^����T�Bn�A�҈�Uj�7/���ǜ��S���3^�a�G%]�d��*�B:�:�[�3_V����f�ʏ%l�j6�B^�\(`�y+V`I3�`$�ܻìO�ۄ枷5�*�&��δ-/ew��S���P���f�Q��
ݏX�����*�=��u�x뻘�ۤQ#�E������1Yki�7v�6���V�q�
�һ��Er�gB9�ő.X�e��9>A衼�Wg;=ٶ�x��#ѝ�6AM��
K}�{$����ldF��K���o�j�tT���b���O��Cv�,I ��k�u�^c�[��b���`Ιz���:�|�Q������G.���o����h���o+��ե�#��)�2�f�������zd`5�TQJدR� �y5ܵ`huљb�{�":����	��kg#o{aպ�|��J���{P�
����E:�����#o� ��yƅ[��Fnv��/��K�8�J��7 ��ѝ����B�+�Z���"�S��!k��K%�c��/���4��<�9��3,����q51��t��]@;�.�l�K��V�:%�᧓U_�������k�.�.��0��U��u��9Ԁ_Z�:{���{�2����jfnS]��=$It20n &���g}N�T���v]��|�V>E�\j��E�)��̑�P�]���rʒG�N5
�0+2�%�wv2�'V;,�����]Q��H N>W���k)�7Ov��P���m';t �U�����3`V�ͫ���ż{�y�vl���ݳFok-'vsČ;�l�̀T�u���*���k��R�U9T���pUh슀�w"�T^S�.o��^=���j�Fog�S�wOY�v!uz���&C�Һd�v�ħJ�Y�;��G*j���!���%7�E�?)�ӰzR���f�����WI�%��R)�����Z�$)ݒ�>�B�pCL�:�e�\�0?�0�W���2�VX̽j=(�1��[h'��h=։(��6�g8���k���
�3jڦ�N�.Ԛ�.2�B�@&u� M���y�f�N�ʕ]k�ا��س�ΌnX��`��h3���y��Sbⱑ�[������q�VR8\z�j��uuN�,&���I^���]e=Z�!����1[��y̳J(2L�+5���M�_���sl~�LKb�gc���`7��"��v���Sn�_nQ�T����\�Q5���*G.c/b4�{�]�W�)7��ܽ�y��*u|���T1]�봵(�k�1h�*��`u+~���7��w��P�,6��4�W����;آ1�47��:]e1K,��]���t+HΌ����97gf�T1�ʥ�'"�މ���N����)5����
���ot�ڢ��̰튉uq��9h�n�k��,c8�ǠP�jP��X(n>c,U�y��Iݙ�E r�7g��}�K���8�4ss������~�_������|?_.|�_���z�[�����[G�`uG
,����N@�6I_�"0K��4���tەNW�#�%#�*��&��	�e����9$,������)����D��=��۟w���桨�2s�sc8�8�ө��X#l�ӊ���%u٤%�u�+#��[CX*�[Hnjo^�a��ݫ�Ƣ�|EI���wo*�FO�no@e��;�b��wq+q�[��]3�YӼ\��x��3m��+��ٖޗ/LQ~ycc��z��;-L�����g)��ɀ���ds7F���.Ң���*�	��+[f�&���'F�3�0�Z��[͑��ԓ`ƴ�q�8� ��O��5�jT����kc��.�qq���p8�҅���	f��68u�ɕ6��!��*T�2�w
\`o_J�f!b���@0Ȏ���-�����w���`���ַ�kjZ�:\G��l�b��՝���OmX�����^�{�)A"�����6�b;9�����Tk����ob�s�ծ��nc�t��!/���m�����b��ۮ�@�ڦ��M�)Z��9�/N��rY8r��ilv�챬lh���D�d�������\��P��ѵq�1�C��{-�+�����.�6j��RJ%� ���[�_Q��g���A[� �Ҏ< ڻ��	عR�,f�&���/��zf$]w�ҡ&�:���'S�5#������!	��k�m���j��x+���E��z�vi����-���	뼚;�t�vZ  J�0D~5U1��-#@�B�ER$3%�	(F�R	 ah��r6�QG r����B䑷��)�2�!��H4#�F���i'B@�U*��T
�AIdQt�U	��?8-����E��$2���!F-8�E��m��8dI�[`�ى$$j~i� �l4TR5�$%� A��R"j��$���}ڂ�J��b�lD��i��b��l�EA>#QTTUS2�A�nm�`�i�*
	(����$�(�X���*b
`�� �b&h�Y�h����"�
" ֤ր�����jb��Z"���*���"��ff(�`��4M��EV��UDUSATѱF-�h�UTS%�S%M�Q4D�QDEL�E4���T�S5UT3U�&�ͪ����4@L�ESD1TQF�&(bj&�&��*��&�*�������(�	jm�QF�"�)(���3�R�L�3%4�A��QkZ��A1DE1UV�"h"�fi�������*""+Nj"��"��H"�*���j������*�����65K�MEk&����"�j�"$����U�APEPD�D�8��3L4�M�����V �O���h]Y+���*z��\e0�דl��[^��uA��S��W�Z�ŕó�[Gsz'R̽!��xr��[�{��yP�G����D��-"�"�Tq�Q"8�0��
D��DB��	� ��^�(�֧�k�%��������s��\�:
�jH���z���"��<�w#[������gu�vhU���dl��7C��6d�z-��<t9M|`Ṵ����7�$��0x@�����Gn���<e�!�Tp�l�1uǟ���ݾȫ�@��Eϣ��m�H����ls�&}����}����)��Ɨ���Zj��C�h^���^�~�o�/�H�����JC�3[=�~>��>5��%+B菽^�����_���x��eoR�s�6j��/=gcEu�{��y�@0��-e]?��Dv��+78y�*Ⱦ��By�="�UI����){������N��j��,�˫S���x�W���.ov��{�kƶU�4�2�D������|ޡ���q��//d��&o�)�����-c�����
��G�m���b���
G��ҡ�0����l��	W�mz����[Y��j���Gr���f����䦿�������Wm���F���\��LԨu�S*���z��q��<�*}��w+�OE�v�<���e:��L�]��Z��0]��EL)!��O�6��*�KU�]5�)R�ތ)\l����5fr��Ͻ�ՠ��LG�t��v��/����Y���k/�p���W��g՞v�%)*VH��oQ3U�~��ͯR&ѹ����6w����ɳ��Z�N�w���6F�f�WG^^��X�wv��d��/��m�Tp΀�s�le�NFU�MѐOcM�1y�*,�g7p�'i�={,D���A�4H3dЌ����[����w��^�s���N���}ꝕb*�F�!�춐`�0�s-�����]�U�=]�Uxm1(�:�������\�1�`S�KwÞ�#�����h� �5A��Z�̍g)��4?1��.{VHX��h�\��1�=�px��&A�������O��/�u�<L|���Jȷ'�Wp�C!����ՙ� 
�m���3=�E�y���s��d�S��BU���u� ��i�%^��X�-���+ƈs�������c��m���U�>��'��o'`.
��Y%�̑%�=,�d�M̽�)r��:����8�eb�SguF~�o?dôt��s�	�/��%��6i~��羺K>������T�9�:[^Gg��o�����k����y�X.�H��O.�v=K�6�쩐�2_��0Г��g�F��:/ Kl{�l�d�|��+�m�������9�)z�m��\}=��ԣVm��rȉ	�'��̽��}����x���S�^��0�y���h(�W����ts��_�J^�گM9q����n�)S��[׾�>c�c.�$�8�g8�/}@jC)ˉ�yl4�D�<�7`�8���:�W��'߼����9�j�r�͏��P4��~�{�O��R�u��@D5�M7�KS%�=�ga����U�����6I�5y����]3��������<�@�G���Z{o���N�	�=���wP���z:�tU����r[]�����~RWY���Wܫ�g��������Oc7�_h�q?�֬�:�/��
�w�S�[KJ-Ʉ�N�<�����^�hҧ�wJ����y�{+���Ԧ�)Dww1���,q�gu��Xz!�b�{���4�P����ݡ;��R�A�F	=L۹����Q�8R�.�����!���R�N�P~��A��'��&��;w;4歯�9��Z. k�w��b��Oу�_��ث���e��b:�ki'��'O���-��m�4����3� ���k�:n'��� 9!�9-�<2��n�&ۏ�l��s=���'Y�Y�XE��>k��v��8\ ��JyT�<~}>3�d�OX���c,�#[=ޡ�>�O!�^e��o��y!)���mC�l^;G�+���jvkL{��W���n`��z(����h�>[\�;A��9���fR
�k�d.�|W�LY����>��wڦ�L�wʥ'�I��n�͌{�z榉|8�îI���$��#�M{o�UT��#6Cm�������|szL����n����+�&�1{�|[�挞�����x��ݕ޶���l��]��[g�*-�ʱq˂E<�2ƻzd�u��(%��WK(�]�/��$3_�hۛ��`z/����s.�۹��/����t�ڮ_�4z;��Ge�W�N�j��޳��X��٬%�2��������&:}5ݴW�V.���`{ٴ:��^��������s#�k��{�n�>��pUd�.uI��T�u����s�9��k[6�O,:��4�&� {ѷ]�(d���{l��n3��;����_t�$��y��Q�����j�����|���;�Ͻ�[��tT�t�I<'�{49n}^#��#]z��K~���za���^D�<[9�Y�tW����Q��S��g�S��>�8����ώ�,�K��.��(�֟T���~��@����k�d2hA����P�����Vs����\\�+Y��v:���b|�����:4��9��'���q�פ?�;I:OP��Qp���
$�]�m�F�@݂Nom�OR��~w<lɺأ���g��U��^��eJ�����ۼ����N�V5U�e�A��L��z='�{^L����v1'�������ޅ;|��:��7{�I]�t�7WA�4sxo�K_K�Y��|�ql"�b�0����0v��_o,#0��Dkq�r�����W�z��of5��,��ƃ��B0���E�W[�&�A2�2aY7�h�DԔ.����R.d��Ә�Kˋ�C��/~�熫f���w�K��cdy��q�.����S�Ƴr(A꠫|Q/�C['�%2����Fۚk(��z������!8p���r}�9ճ�h9>�Ӵ	�����{�7��m�/�1L}��K����p�a�Y��/h��'���q��D}7M`�OJ�l瞮�O-�)�rw��Zu,�'�T�S��O6����*Ǜz�iʊA:�F�O�ω�>U��4��n�. �[Yͺ~��e3�������]��>K����*F:��Aq��/� @�y�0Nw�[5���m�.�a}!���~~�y��`�|��;�Ƕ&/�;���׽����ւ���[�����z+�I�z��Pe���?T��2u�<�Ř[�`b���nW���/��+�IΣ�h_A�.�����V#n�N�j�ͳ�h�#�8���Ǔ���ۣ܃�<i^��^X�'.q�f%�P������G�����9�/�S1�u"�E��v�V��z��֬VЭW[��%����f��0v�ţs.�I��zP���Zw���4��Un�tퟭ�~����ר��^R�����VNJ{���<��F)r{d3z���U۠'i��T��0L�ѯP,q�ƌl&��n�g4��$�9<�SI<j���ә�@��9�����Lh����;�5S�f�N����l�{���{��>�mbl�'C}hm���o�EG�ו�}�u�
�]h>b3&8f^�g���z�i�ǺN�����-�+վ��߄�lZ�=�/S�<�����=���7��ۏD��X�7g��9gx�t�{1�� �BF�oz#�%�fEBN��hr��W�q��W�!����w�h�Mq[t�ƥ1)˥�Տ>gz�z�.l����K`"�_���>y�~�^N<S�VS5o��bW�#p!9Yv'd/�o:�}��t���E�M��ӗ�E�Rd�[�j�S�?q'�U�x-V.!��F������l֜"�
���/$�wx�M`M��J�q�uf��<e�g`�P�0�����5~�Ϯ�[t�k��0.��-�L�͑]I�i�ŎU��2�o1�v�#� �w�/M� ��z�p��
��ۏD���j���ev9 
S�z���w���
{[�AT�2�S�7�伎�����Skݘ�s���.�W�9���W@x$ףo+�۷u��Gl��՘�u�N}��Ư6]��K�#b�g%���"�Q뙩�Ǫ$��w��D�Ƃt��I5�H�X$���y{�Yn祧�Ǭa��Fl���b+qR���^��^�#���2(�'��*�%��jE�ϵ�_��y������5�:3LJ�o�k�L�=v�vi�շ^s��3���x��ӷ(�_ȍ��6��5��^���M�秷C�q9����Xٺ��x	��ؑO��S7�@��lO�d���ƞ{�ܹ����A�(�8���F��F.��vЕ�rT�����d��
��~�|%n�m��q/}~y�1�jݼ������9�uG�a������i0��I�����fӻR�x�|A�ڣ�Vs	ˏeȾ�
r��h{8�0��{7�0+�U�c]F����s�p80q��N���Y8�U������[�4�DJ����ʂ��W�u)պ:�����7\GL��ۥQ4���uӋ�t��6:����B�H�%�VZ�v�Zb��i�,�r���0;w���������S���}�=�����|�Uw�otɜ�6�zX^����ϭv���sx[�-;ۑi�;=��h׳��}��n�y瑤�[ܭ~O��'�Z�#�<@>kp2#��v�a=���ߜ�R��02x�{:B�&/M���e�R¯U�{\k���N.�̔.�k.�����xc�,�G�C� ~�J��*+�u�Ϻ{v�J����F����e���g�݌t�'�H����I��Oӏ�{�+��vI���+3G\���q��K�W�n�R}��P5O�Oz�7�8R�A��+U�
9�n�)N��=9��e#�b���~'����)�˸��jI=m�f�z�_�6�;tP- �Op̮�';X��Q�Y�H9dף#u����6_�jO]7�ݳ�B����k�5]�Dsf�Sa���-�E
V�^]5ۦ8j�u�om����֧aG�57�$�ͭ��0o�d�|��%i��/g�E����f��]c;k�Q��[,�;�U|_I"T`)|H�}�����{��i��=�+R��X�s�M\]&Kv��8fWqۏ�)9E~����\~�{| m��6�z����fa�6�3K�����&t�qp���v��/��eh��W���:�u�헝R�4�r�m��<��p~�-�g���e��@�q�'g�8l���m[S<3���Ƙ#	x�kǤ�ւ��~����D}��t�GB�sȮ�{�h�~J����6/;�>^�zC^p?���_�?wg�sZI�K�S����E��/��b�w�=0��oپ��W��g�LYG�Y��+Y����z��W¼������o��G���4ɨsN����8��ƽ!�{�����?:v>o@q�<��w��ht<;��Ua�1=�Fg{�F�.������c5QuC�ڹ��h��z��_P�^�˼i|vl�T�)i�^�'�;�d���׳���^C���ςg��z�=}=~��z���~�_�����{�}������T�no�7�hj��f��9�Y���ZX����(`�@�O�zQ���J���XLDwu��r�(��h����a�\䬧��w�#������P݋bTzY��h�x	�y���BCmJ�A�a�K�=��X�we�,�ܧ�SRr(�nH���o&�̔n���Bޭ�}].�+�7���w��[[�N	*Z�b��8�J��R����9��RA2_kj��;�Q�<n�3h�v*R�u[�dӽcU������Hid�n�A*�t�p�FA�9f���cM�r<%b����w�^��R��	��2�����R� �N#y3;��n�uB�(��r�ᤍ��=U���%I˪:�@f��V֎�ǃW�F�E8�*��P���Uo%�6j@���+-�s�c�It	v�B��e���"+�V���|o�� ,�H2�(��>"�����y�"o/S6<2�tv��J�u�l]Bk�oF����}OywF�-�\�^w�YdL�/�@ޔ�B` b	��>d�W c��yR�qʹ7K�,%ԟq�fR�$+�v����(�9Y��X�=���Cm��N�ve�Ą�ke-cb���������@���N�HZ3�����-!B�pʔUo=F� r���\�v����+��Z�3��=��֡���۬��1���{��0�b��G�#v�N��҄��L�_>-�p���[��ʽ#r�N��ȴ^�u��ݴ���k���!r�P�t �]Y����J��Y�B�~����}������\��7��l��+�^��C/'=;2�p�dV��\0٦�W{�ߡ�"����u�\�O3�F�H��$9Vk1�;�}C4<�V�>:�3&�Uǵofx-c���,ɮ��rlX�,L�}V�aǴk����|�����g`�U��2
��74�����'u%_Moz�o9�c%Z,n���-�ίZϻLsX���sC<�&����G����͇�'��-����y}Jq��*��.T�r"�YP�!�BV
�7���+��LLD[����õP�Ɓ�N\[��+����+���(���f�m��u�e�qQ����خlYɦ۾��X��ʻǰ��r每��A �pg\uoO�P:K�)8���.�Z6V`�8���ٻ�o�\jgg~@�
��iq/�ȓ������ {w�[���s����0��P�ΰ���������\��Z�'@"�h��N��mM�}}N��5:䵫Q���6�6�k �vE��dj:=��a1&��ƪ:�o#�����/w��cb8�j��v�<|���;�M0�	3�n�T�)1��.f
�yG�~�5f���{�����(7fPÓ"O]��)��MmXyJ� t���\�ct��r�Ǘ[�N٣q�ںα��.��	f*�p���
sub����EMUL4Q1RM4U�Q�9��b	�*(��kb�FJb�)���"""����a�b%&���`�bf�b**��j�*����#Z�����ESUPPD�S�lj�	 ����*h"��(�"*�b)�/|�j���)���&��hb ��	��&"vƱ1��4D%DT�LUA$EUE���Ji����b&�ib�	���j"�q1QMQT�Q4�ULED�A4E5DE�A��PUE$O�s�ب&
���*�1��1���*�j�H��5�عh��X�(-:�9r���"*	�d�TS%EUSl���h��r��[��P7,i�Q�����;��MA<y�U�lm�,V�b)�Ni.Z6�dڍi���9�\4S#V�Y�并B�mV�Ebfj�1M<��X�y��k!����s-�夎&p��a؞p�Ej���Qh+h�ha+�b��'Z��EF#U�Y2lh��p�Dm�`�TC��l͜hŪ��Z"�>q0r�����Q`�V�n���߻X2���63�uFH�;R5ys���s�l)}Rә�ͥ%UƓ�o��K�<H��R,��մ��}�5^ގ>��7��{��MzJ�s/z��A���0v�rC�p>'��)�ck�#Ն����b��U�?��5S��_����|`j��_�;�~��sW��&u�a�,��R]����p]t<���qm�Bػ���N���ֆubK!�FFS��T�y�rf�RR͝�PeAd��\�"����[��.ｽT|yl�z�o��)��a�y��O
UX�+���"[zr-�uE�˃�kv��%uX�O���}�E�~3�(�f=zޭ�[����0D�� }�d�y�&f��5񋕤�Q�c�Y:���rq4�:J},�D�I����|njgO����aD�f���/H8n�'T��h��l6�g����-�j�%�|���H�T4����{�l�=W���[���'��������0����o��v
Gd�q#��|�E'(t	\���5\	���(����Wn���gwfw^���@�A�t!6И��#ry���S>�	�����)���H=�1N�Ѫi�7��os�)d�L$i��,"�/'ֱG8}xeϝW Su���x>q��)��c�m��@�|�g��;5�1��J���P�Kq�lx7#��<f�Vo�,pa3�������3ucyZ[�+c� ]�Q�������I�9B05w5��c�2�hҚ�0e ��r]\��-�:��3:��͡/7�w,Z����t�!m���y²��<�GVE~��Br��G�ޡ��P�tf���6n"$��7�S�������\ͺ����{��1�+��P���$N�75)&7ߓ��]Q;P����E��]z�'��c�^/�U��O���uƇ��_��_2h\Q���|���a��I��f�}��ž�9lנj�������pl�i�{�y�����3tŸ[��^ÿ�&���t�*��\/A���g�|#Yہr��+_��K�l[�\��B+��j������Z�.h;+B������+O�����R�.�>!�ߚ�a|��=��g�:��.��S��:x��7�5�e4%p��;�s�>f ����M�5���6�dS��?��1A��<ܿ>��OP��Tn��lή����/�rHq�����5��A��f�?V1e|�*I��0?�S�@f=7��HY�XV��z�o�p_x�|)|%EcRQ���� ��)�A#X�F;�j#������~?!��%zGn�٫��|�����ӽ:�5z2=tG��=�1I�%"Q���5y\[N�\:oO���¿g�o�ivl��2� ��hެ�g��n.4V����[�N_Xilh�i�{��X�ӹ���0�+%�ם��\9�^�x����9�u	/f��E�PwAe����3D�k�w�,je��Y��u]c��F=fL�X�/�&'p4�{��+��)�Q��|� �c�����o��"�0�V>�*x�BB1�
Y���=�.�������&I�lD�W�W�TS�oL�:xl���&ې����6�,�h��5;{E#Y���2��.�w:a��ԩ2� @LS��&���V�}�9��Su7n���A9�/�w�xaB[͹ `fA� 9	�8#�=�Yv��gmg�K�2����U�+-�r�e�0���z^F��G�x�X
����_�r��ˏ��$���Y�w�ÔY�.Տ҃ƙ,$�ye�7)<�Rc�e�jxwfܟB��R��ᢽ���~��cu���܇5۠�+��l���w�J�¼����?O�8SFJ:��E{M
Z����Brs�l�\-���X�����@P�p��n��еaD�q���~*	{k��H[Bu�2�A���dwn�V���P8�<�Br�m��˲��Ú�:�a?Mk�wh����oN�4�\s�Txf�����*ke�7�Q{���z�`<h����ߏ��fT���,�u_��⻇��Q�Vc�Ds�����f��x%2� �cC�[9yח�����CY��S���O�_���!����{�K����&MV�(&n�8R�*Wx��d��N����뾛ae� ����v�;�173e��Hִ����;u���n��v�}��b�δ�hp;u�xH�^C ���6%�P��:�N;sm�ݳ��2��j]�o_ �����q�u�/.��l�H�,�PHx�.��z	@A�v6�wC��ƶ3��e��4a��(��dٖ����^��݌i��<5� �O�`���|�.�,��u֢?�W&�~Ѭ����>=V�H?a�;�Z�Xg�0��%��o)����ր����p���xj�l���<ئ���	�1��Ά,6~g`��g+��njJ�;XF|*
NF͞zU��X�;oo]�����b�L�J�,|<����e~����>�y��	LoC�|������5�63-��SOhr���-^�U�9�^��xO^��x���<� �S'��+��W���r��u��X���,Q^C�ʷE�'C^X��)󊎉�^g�n,���2r ��}���ٙ]�St�G�T�9�5,֑*�ey�.�Z5(����i�`;�u9j��50qu&�7���qf�B8E����3��B�����W�O�t�1i���]&��N%Án�970�YE�3�������ݔ��0rŤB�lė[�S�QӴ.�*��Z��R�Gs��oR��ew�M!ⲡ0�I��d��X��6��Rt�d��&r�Hjt�z,�Fk��뺮����ǆ|a�>� ~ �10����]��C�X�oP��Xm[�W�dga��e!e�=X%��%ۋi�4�P'7uK�]�� D�eԹ?~�~�%��_���*A1��z}`�0��u����U��-l�J�aD��pOQ��	j���]-x+L�#o�� - +�f��E�~��3��~/b��>;���:}�d�3�5�褛���h~�u�P/
�l �ӯC����f:Xgc �h���c���I� �g=�+E١�^�Ƴ�����HGz�4��gHfRrQ~���!�Ĉh���D[�u�v2:%�,3��;^����=��6?&�ӷ��p�"L�{5�|��a��P��F�D=D$��b�)�cb*�دu��o����eóS����h��ϼ�s�W���3~��f�e0T9e(r���y�y�}F,K���o�gݟL_yKL��S�҂�Ϗ��*���[�6ڒ�l�M��!��:���|����[Od�Y�����X�ȧg�-�7��V0F�;=gD�uJj5�r���ۣ��v�@kZ�(2j�Xf�ܣ:=�V�o����(#zi�2�@$o����갆
]ws�:�А�r���N+�K$���er�&���|`(s�:y�=�ă������laA�a�բ�l�L�H,v�ϡ�c�N����j��ǉfu��u�J`wamHݧ��cf�5˞��5��	�{��:��aڴF�\�����v{m��қ��]����8�lwr�=�4E���atҭQK�g��>�ku�^`���`>�+��9�r�|{]����'��
e�9�Ks��b�	��Ğ������^|��M���X�Kg-΍{������BRͭ�]R;%�)�;��O�"���n��Z�MV��� О�	��p��U�;#9�*�f�7�"���AЄ�Bc�l�O5��a��&�p	zO��U}���ea�}f��Gk(�j=�V: �y
�3>��?i��G�Lk�!�r�N�߫���c]�����p�ʟ)>�_*��H-�{˹p?aC��5�D?��H�B�y쟍uP�tތi���a�L�j9�+vƠZTX֌$��::���50�/��H���(x.!��@o��iN�9}ڕ��z?���u�P���K�Jo,��x������j/��:�;w;�4�~�&��n=�Y���>��f��� 2}��A���I��pZ�V���զ+����,���y�n��	;B�:����/��A�v�\��&9��#Y+���Ƕ(E4]�ñoz�gD^w0�@�v=ܩ� ���:=o={"]�����DL$�&�����s����d�����Ϙ�~�oKA��ư�C�:k�i���[�f�^&h�vwV�<#u�+.j`�:�&gM�]��wGI[��o�Q �%ɼt0���d�����V1��w�(�����8��Z����_:���* ;KQb�q^Y9v�z��z�`�x�^�����KR��x�Ϻ�B��5����B������a�k�L�H�ƴ��}Y J�_���Ǵ(>�X)���n_�6�-�����ظ.u=�C��2`)+��3���8ʆ@�t���V�`����e��љ��)����x<dT�V5�!>��A9�K*K���c�C*.ۆko.��O/��-k����}E.<�a��;�ʹ�>���(2��1G��*�J���`)�90����ӇbWo;^ʈyJ9�="A�,�Ba'm�v��	���$�����F����P�ߚ��n�컹ap[�21���hT:q��i�:Añ��r���Θi�>L�7�B��՜��A5��5�0'%Ɓ�A�/A�-��@A��!�O�&���L�Ğ�ef3���"������b���搴����sW;73���+/��ڠk��  �/������r�~��y��{$����^Yz��O)Ac�%�$���܇ǟ8|moR6"om�l�3M������5[Q\��ȣ���.�TX:ΞeE]s	/v��t*�����;���9���e�o]�T�(Mi�">
�ni�賊6^��4�<�3e��{4�2�/���#���ǒ����Iq���x��_�}nr�G*<��N�q�pf·sk�
8p�t�uMf�[3�w\ې��6��ܨk&�8wD�E]=h��Ž� ���&��j�P�!�|��`�ֿ@PX�T�m�;MI�c�wy�J���ʎo�{m���S�S�p�E�;��s	?���6�����f[^�Ú�u*��֠3Է}�#�cC�u[��}mv6Oэ����RP1����g3�B������omu�ʄ����t'��ï�p�Q���C��\��9ۺ��f]��C��B���ڢO��$��,?��V錶Ľ�p[;��d�&c}Jڹ4�#2,���t�C�Pi�e��zd��y�π���1�[�0��(�u��ްv�!����Qx���cH̄��W� �K$!�Ϛ���l=C��r��O���6��f'c��4 ����.=mE�1��NT��jR�� ��H��%G\;z�ͦ��G�����u�8��*o��C��zg��c`�M~��Ҷq��NԷ0�D���2&�vw�3mLd�U~��k�8?Q���t������::�@ �Ʉ���		�ex��ا��[c-.�k��i�ш�[�൭y<J~���L�����z��	��=!Ųd��	�Bp+��
S
S�S"g���Н� �2�ndv��PY�K�9
G)C�[B-�+�E�si�kD�߯:e'�d��fq��ş�0Ğ2�������؜�ۄ��G�,���28�U�7�%!�a2u�7����jT�:&.E4_=E����s�������a� �< � ��j�J�u���}}.~ �K$���RF��q�w0�i�f�.�����-ʇ�U�v�~�.�0��^��� iݒa�vEL,#R���eKMCuNY�6�(��d��K(�ۊ;�	n���B��`&�����P��⮗�1i��rą�����&�SU�좁z�B:����&֨B5��������.�X�QoKW�Gs�J�*+b�q���N��m�܆k�-�� �r�"5�{��:��SL�����R�[�^4T�SP�hd��:��zo�Mے��T������;\��t�%~�=�>�4u�G�r]���*���F�[�h�ζ�ޮoi��\�3��o�rb9�\3���0��E����]�:���&��u��W���Ъ����f���d��Y�9!�a�x�zb�`��g�$q��'��^�L��� �H�೜O�W�d=�����"d3x�E�v;�HrC�4��i�[�Xʻ��3Wv(ē��Q��Y�`��KJ	���|��^=���#73M{�KA,��yy��F��v���7�����[��+����{�W��������g*�N��1d���
�L�Y�%�F^��c��<��k��~^|zѩu�P[;E��6����B�v8��T�k�c\���$�=�4^��ɲ�ޘ�*���Ǐ׃�W�"�H"~�M
�HBP4�-5	 �I�	$�羆�{����H/[�/�)i��vHo������-��?N[����}���Y��bze؅3�V�ݹ����4�E0�'�C�����V��>���\zx)�`����A�7���ro�빮�ğ(HO6Z2�/7��a�O`J3�(�f=[ռ�|w���%���3�	���wyB�aQ���h:�n�A�O1�A�	�1,��bY%MvGc�W��t�On�oA��X0��`>��vm���OcH"@��A�%:O�J\M7���˒ Rkk����JJ,�{��'�{�Q)G�C5��ۓ pc=��dq��I>I����-?���z[]钢ϚEooa,���z|��l;!������;7'��������Z4�s��'u���xt������������u.�a'�?O�E�2�F��r9ĈؖM�k깦��Z�Py����`��f�}���}b�Nsy��1��c8�1.��u����0>b]ِ���+�~�R��K�3Q>�+����AU�}Г��M�X
�z<j��<��zھx�ȳ�}�O����/��_Ǐ^�z�����}��}>�O��~^ysϿ?x�X[3ϨM8�WZ�ph�ֹE5#y���n3H��Γ�tr�����Ю�-V��>W���(ʴ�Ҋޜ<3��#�1�iMcYƯ�0�+d��f�8]�C�軦�83fY���@����Iiֺ�R����Ɩ�r��J�'DZ��^J޼q����x��L�v�h�.hѦ�� lIr�:�Ft\��\�7Q'ُcO�ș��Hz�l�\��k�ς�]�֬�i����+������@q���Y�1L<Bͬ���|��n�a�*�M�{�`�\�����a���$��js{Om773,Rǲi��������s�~����{A�~�k�#������Go�iD�諾5�Ԝ�`���֋��$�gZc���2���ykgi!�hb�a�U�):�3|��To9A��(Lf��"��%�45W�rQ)��/�S���Ds��3���Xn�lY����A���tR�t*sڇ^qm�8y�L#6'��FCN���6p."�>�����Z@w�E.�$��d��4�ά��9�i@�p�e�0g0/�5@�x+��*�3�(Eu�n{�g��|���Ћ����t99uo���������Nz�h~���ɮ���4J6f�~!�xvk����0�)��b`�����l�Y+�Y���D���q��V,�3b9�dv��n�~G��7�q~��։XseÙ�;�J�N'@p�/��[u��e^!���us���/�Ӂkv��,Ç!n^	? ������ ���j\��Ϣ���b��޴�Y(�'���6�9P���g���x�M��r���U��p"�}0�-'2�)��ۑ�8�W��ؒ����Z�9^�i٘��u�вq� �8i��q���hD��&������gti�����L�@elmOd�ub|���y���0�ݔK ��l|){@�:�g��rCʯf�E[I,���_l�Į8��6LK��']*v�]s�~�p�+�߷��n�-xɇ�+[Ҙ�y#��'�Ԙ]�vmw�s`�K�e��f�EX�.j�S����/r]��C�"��t��[Mu�i[ .WZ��˙�s��[h���r���eL�Q��4:mdۏ����L�bưLg3n�g���#u)�UgD#;aQ�
�M��U�6�}�#0oq��-�����˷�xΡO�Ǌ`�[eӴ�FA���t{7p��5�[�wTZ�N���вw/���e4�p$6�I�N�uf��ǫ��s9v��dXLvy
�v����c�<Z^��EMk��
v�&��1�H���n�q_[��(\-�gtfF^f�����c���v�[8���>����Ѽ���ӳ��$:�im��t��.�I�"�eЉ��s�J�oQ��t.>܁�xi�T��,qk�Yb���| �-!T2�����.��xt��H�G�
�4=��8�U��V1��N#��6��cV�Z5kV6H�NvsE��Iͨ���%6�ư�UF�������,lDELF1����0�MQF6����ƴC3EQTDD�RU�SLEV�\�Q3K�D�5����QV�DV-4�4�D���c��h����b��)�j
ba���bh"�r�[*.lPQUUMM���h"��
jH+�s-j���(�b�.`5SU5AIUQQr4�ƪ媢����E��"#cETL�0R�si�)(��(����Z"(�����*(ш*�m1��U5L�!ԑ3R�L�DTD�P�ET�5E4APTPT1$AT�UD�L�5Q��FJ�9.I)
b)����H"
J����"�*��"�����H�&�Z�)� ��`�$*��h���
�����y߇���z׍p-B�$0���^���o��8��Z����29�� �{{Zw	W%C��`]������혱-v���F�\GY� ��z�]࣐XI ��`��jS��%
n5I�A�	a0�8���< �����Vbi��xSm3�&�X1:����}��~��M��x�Z�8������j��z�;sx�g�ں���V�m����A���-��t؞�����i��rQqź%���v�LW0l6�fuf$A����D��57��/z��坮¿Ij��-s}R5��wW�s�;��P&@����ڽ���V>�j�h�ñ;C�c��v����6�hl&>2��o�����S��wA��I��e���(�b��u��f���e�g�r2�<��|iO\�M��ȧx	�!���p�ܓf�G,���MO�x��G@�u�+�V6H8�0��,����<nus+��;Ń�k2�&u�T�_¬#�V�S�鬐��r+����^��b�]X�_��eE���y��H;>���K9b9	��y��#�i��T9����1I�V1*�U�p;��f���Qn�R�T\?[�>zD&�(2�p�;g�%��)���L�و��`��_wFv��Yk��_?n�X�Ws������k�����~$F��m�x�s�5�ą���4D*��%�N<nkk_K-X���}��Üi�<.f�K���Dl���8xS��F���0��󇽻��BT�[���S���%��y;��@��V�ܢSӌ�]e�j�Pޗ�d�9���J/d���������e�htNh3����W��~�� x{���S�LY�곍�y<˯��):\dp�;�0�AƑB~�s��e�x��qщ5�s؅4��T4�r���6Ⱥ�7���h��A.+�+?>�U+J�3����Sqc�OW`�������)T��vS	7~��L���)),kܶ���<;�F�>=�5��k���%^>౻͍n�.�TW8�ȣ����@��E��<ʕN��^�>�cX�cB�Rm�Z�à�0g���t���sL	�{�G6�i�j�J���y����/�S�0r���!黛dRk����6�܈�C��<O�<?��h69�6'9��v[^�Ø�RM�~�C%e���f�Ĭ�A(v���[��1�������D�yZ�4��쌟�����1���]��9)�C��V�0�Q%ډ�c�D̻'D[�@�r�.���24F{e��u�/�ok-^�v�r�� f��wS0�{A�=� ��� �O�t�O��U�467m���3���Ӄ������(��q1�'�f��M���9�Hxn� �%���r5�\e�m G�y巩���P��������#VL�v;e[%�c��j�G�LS��T̂��%���+M�
*mm��Q-�z|����&+u����������"`Trw![���`%��+�$��m�;����Ah,��]��<[�O|x��ǟ�(~�P
Dc���_>�:�X L��S>L(Xt\H����*���*Zڽ�HZ�atR�{Tl�P�d�)�c/6����"�/\�C�tW�x᱂?�|����?}bmCƇAl�V��U)��b1M��A0MU=�B�b����e�YE�s��2��^{�J�6T'&~���4v>����D5�x���2�&�B*��l�=[���-kE0����m磁����3�^�x�w�t��}�G��
r�x�O�$Lu\��FS�p����s�ߪe�Ku#[�����O�~]$���v49�F{"����	�Y 9�W������rۣs�n�fPp�a0��1t>>�vb��Bn�����:�P�*������PX��јn����1{�iռ�<��q.���:mi���6���58��^��v	Te���jr�a��.s�r��_c�[��}롼������A��y~<�4k�mM6�%��:n2@�L�f,�k��s-�e�d�eA/t��4��̦n�N�]:
��'����h����?z��qz���b`t�'~��ڝn��ҿ�֗�]*f�׸��7�]�=�GƵ.6(w'�q����o�͙FC��X������a���>��,5�9:��Q^Y�jy3{d`�M]2uZ��%l���3�1v� MD�A�{n�Q^}{��� B����{�z���0�u;T��{f�Y�I���m����^����v�v
9�%�Jug[���0~��M'����;�k�V�uCs�n�f��_����C�^h4��Nh�b�P��sn�9���z}Ţ�*�`� ���� ���7�mt������0v��$9!���c�w��K�ݼ�bk�˅?�
"��tK<x���������{d��=�g�F�f�i��%��ٖ�g�$D]ݩ:��l!�w��/%�W)i�'�J�>0χ��<�����ό����g��K㫞Û�L�v��f��Pe^Y6�5��|ش��O�AI<Y�~�T�>�j�κ���}x��[�Iy#Gu疰��y��)�єɫ��{��
�=�V�o����x �d�3k񋈜0$"q�XE� e����@C���!8��%�t�K#�F�]�v>5{gNێ�Z2Z�0.׋#s2�L��r�]]�(	��H�ivA��?D�I˼'D.�L�#I��k]��=.�V�BL��c��e���6= �5�JY��,����L8�wQ��������=*��6C��i̓���7�:�������;�byoʲ�u��i�����[6�W�+�W��)��C{�t>�۽c���;~7Uv��.�����j6�!K�S����T�\o�m&jT����-�.��6�+^�e��m�`�=s>z��~�|������ �B
�#��sO�N�]w��K�>Z�1�|�1V�LK�}���"�BG�Ȅ�^��l�a������
��0Vk��d��X�/�辔)�1/j�����s��#���Brg�OubC餱uF[�!SR�s]��0��k(~I�!�;G�H��j��]��p!�����,�:y1{�2&ߑ��k��Mֻ픟��\8��=��K6W�-ݛdl0c��i�p�r��{_��2�	�y�'�OC��j��Z!D��Ʋ��q1��쨮j��=������l4m�l��y��W0.ڔ0g�� �:b���_}��kݱ�B8��StK8��	��uc!Ctp����-@��q���Ds;F�&9ف������hE^��"vd˶-�ؽ�j��w,.�z̻k%��4��ǡ�6�k�"]�|gE�6����Ggiy��:�]0����m�j���Ꮧ��i�+��v�
�d�#.�㑭���®�N��!�Lpݗ��*���M�+z�k.��}F�b��gAA�0�&��Pd�[>���T@�t��>���0�@��1�xX3)��!,��Ul�qK؆%�����qۻ�U��jN�2����yS��2�J�];�L�NJ��I`J��)n��x:��]X:]K��~��Z�t�@��D����%*��)�����k�$�.�&T�s�3���>���B� �
+�����}����#E!|��!��TM���m�����]��	eA.�g/��ӂ�f���m'>ǣ�u|�ϼ�(`��9��`�:ɪ2=�A�=�1IՌJ�&���ܹ�uB��X�|7�]��,a̼�'�Eê��3���Pe���	;O�%ۄ�Jnj~��9��Y�Ky�n��X�n\�����&Er�E8���ȶ�C�� �ƟC�H�!�ʀ�j�N��m����Ȍ�]1�a�C�*L���[t�N���/N�o'r�i0B~�F;�a���b�M�F!"^��1]���vT��LS"�s�e��m�\���Ϟp�θ,R��`Ic��:�m��X�`�t!�mǆ���F�i0���]����l%%��i� �٧�U�K��J��\�msni�ݤ��55����@M���Q\��e%���U���U��`wy�]ۦ���{B��������ǹ�x3���X>�4��Ƽ:�smv��(��:�~��\�EC�>�ʤ��Q�-|+L��ò���|Нj��z�d5��@|NhN˲��Xs0����W���k3�4&�v ��$�Ӗ�������,�Ή\��y�Kݫ�ym�A
~����K!�ow�)rͨ�R#V���߲�{�`j���X� ���,��O�GG�^pp�=���$�iu*� ���T����#+\�G�dy�z�����_�?�@DPf {U�vR%��c�������v��P��c<���^��D�y�|AKi�pխpcv���vMp�z��_��,�V�Qa�Iv�,���3�{���W�Q&��@�o�2�ۺ>_}�i��:��{aY78�wK0����C�Pi����p=2Ή��0�ׯ����m�;5d�@���LfI/2��M�v1�2	�������Z���G�ks�o���ғ�#�`�������l��q��4��Z�2a���T��xaP*s�b`sK�x3#5yht��t/W*�p���uk
�9��3�[pL|cA�3��a��j,X��剋�?^:B����pu�R%�D��(���uV*�����v`�	ಿF>�j�0�"oY�|hʫx�B�>����KPr��6x��Ғ�5F|�[�]�}Ǆ�-��$8�ӵ����j�+���~h�qc��`C�פwo��u�<Kbu��L�$i0nz��s	⦝�;]�텛��s��Ya���!0\�.�G7cH�]�[��;"���J.�s�2���7g�z�{���|}�+y��h�j�6X���R��m������k��^�h�x�;�R�9[�yS��e�kZ��I��Yxt@S~�KA�1o���祏X9F�����̷3�ۿ5��h�_@��.֯�˫9հ�(�&���;2t�w!�����Ϯx���~�x���'�JT�U��T
]��w������{�����O󇖎����B`&��4(��P�ʮ��1i��Ъ6���w�˫�A�o*lEOC���K�:�������k:��tuM'��:rEu]4�v��粳��Ogm*�^F59�
�w=�Oܫ��Om�>H�������WV��[��M����I���a�u[��8��W=����{��7P͹�l��ØO���$3Oi�5��Q=6}�.�}ɋ�!
���ˌ�Lm<u>߸ϧ^�L�5�f5�b�;0�<"N��r��W�5!��C�|/cj?Pݐͳ��E��^=$= �b�t=1m��ԭ�g�L�I�{��!��`���A�Ĉ�6^��5��h6x��ci�uzIHpE�i�z�d.xY͍v�ޕ��ů�[���¼Ś�c��g��X7�M�e5�/%�4c�A��\���q'�9KH�������z�xh5B�.,���bȽ������+��U�f����G�v�L�c�ʼ�m�j	������1��t�w�� c`?yW�?OUY��Qa�x��I�6V���j��D+䧽���Dӎ	D�
��j^A���ۋ��ߍj���u�fg�& A�~.���7,����V�͙lG����5P�ޕ�sn�����Ê�^�Z�'Iޭ�x�;�p9[ԟeIJ�j��h9�W��{��=�{�JE�F�)QiQ
 |��=��oxv�Q�B�OyOy�'�5�u���(�����k�7eԝE��'���Α�/;a�OҌ�
���z��[�z��v�����-���6�;5ci�|�!�%�H�CΝ�EF*���t �W�Ĳ�HĲ"Q���������3mSO�;�R���vxt�y	�Y�N͔&"�H"@��A�%:O��N�t�e�ǟ�S�X���E����-O�p�<�3[L%,�SOd�=�o�������4�T���홇�0v!�2j|�H���0�c�?�p0�`��Ȅ�Bc�n�sIv��1���	D���Vb�1�2�T��1�g�H%�'���a'�?H=�+X>���[�b�6ƾW��5�T>������2��k��B/ԍeIGs�,g�%ݣ�>�ha!���-��з��;E�[r;2�C���ڡ\��jE1rfڳ�R~kZd�Ҩ�kǧvl}8�p�1�UW����L ��:��vNK�o�;�����Q)�P/�^�����Esi�9��B�!�U��d?�4!��d0n���ŤC�azP���M�^J!=�3���=����|>�@�+�]y�1^O������L�f�+k�o���r;}k69�ZyL����჻Bˮ!A���lw`���D*
���MwaR:�:e��]��,�����r�fVޚ�ڠYE�"�y��7�*}�o��e���j}c�)nW�<���������
@X�ZP
X$ ���UfhP(Ti�R��������y~{����k�TV2n鴽�q s�<������mG�kw��M�׿n��m�Z�*�cv5\���U8��T'q>Z"��<�­�.�0>��p�-"&:�7Q�7P�f�8�}W�KQ���{����3��e�f�����IN2\��M�5��y����*4([�ɚ�L��Wю٪��=Ƶ����W_�b��� ⋠ŗ��A�1l�3gV@�t�nm[R7��[[kgv��������c'��5������<�f�!>��� ��@�It�;��]3���T7���t��ʢ�ոf��@��Jq������Y5�\�:!�{b���V��y�伆��Bvt��cC~���\|)�ۗ�������t�^Pe���vۇn��M�dh@�Bґ}�Z�T��Rێ����a#BՉ
�qv#�Od[B�t�zA�`C�L9�[=��74���?sn'w�;@o���I5�&E�&)7H��q�L���O6=pA��T��c��o9V�-�s([��%���5=�%=ȺL`sO����Msӿ3����|��>^�/g�����{���w��������~�65p�i1��"�V��G��CSC܊� ����x�s���v�����k����l�W#�棹o�So%����fm�9����J�V����ف�^)�44��Z5�5_�)��L-Rn��B)2���}��ެ����{�[����+3Y[+o�AO�U�c{�n������+f^Xq�7�O_RR�6�I��,���B=�ٻs3 �@��X�$p>y��c(׍n��z���ل&f��uh��498].<�����\k7�܂Ṽ�}kmy���'��6s��+	3�%$�؜.�.{h�i���Yyb֘2�谫�}��h�nP��G$��뷑�H�B�um\7����`/�f��J=�"ce�2`3�ݷ�h�X��B�t��ωN*ş\���׷܅��=b����,l$�z1��ɜ���|��Q�܃kZ��	x)mc�]�YR�M�/�Zzr%�n���u-����k����le���M�+^4��k��	c+oz�J��wq���hӗ�b�=��U_(��pR��E�d6Цf�{�-q�u��7z��[�sF�\Ae���9�Ϟ���Z�gK���K�ޤF��i�� �/�U��J��rIM�.�f�|��K�mI ��d9]�%�:�2�p�S�7؆Z9�w^�Tc���pJ�R�bM��dԉ�9�3���켅���s���� ҝ��Bm�;�7�\U-"�`{�h%g��^eiT�B�u���=��M��wr��2]��ʼN�t�LP��,U�\J��h��ٶ�zA�!��i�w�M(4�J��䂙w9����Z�Rӣl�[�Gp����Mu���~�܃u<�6!+O�Ǚ��Z��a*��{�M���}�K�t�	C9:6���O(��T�,Ydiu�:��D�NS��Xz�g����*�[�	���]��\����m��A6���'6Cܝ��JsA����I�EG�2�^�������{��=��93]%p���qY��F�f
�����4sI�z��yIh}���ؒģ�N�{�:�b�� .���4��9��<���4�Zze�1�ѻƠ����x>�A�G�Q��J��2tPӈ�6q�^�{����!���+(�C�4ʱ��e�ٵ�|��2Jp9t����ݨ�v�V3��mn�8��VS���B��mJҘY鶽�ˤ��_�ǳ�h�L�K���+RӜ��rN������`�%a�OG���ZŁ�B�x5q�iK�޽-\�Cl�/�7QQΖ���E'Z��G]k"�[�]0ŧ�()�òإηTO�
!n���BO)t��Bm��r<�I=��Yt�
�_%_�ĺ�� (�{d�k3z�m��F�����Ⱦ�i�Wb�r{lP���x��[�gT�y����}ʹj�%Bp�y��֦;WAr{�Ov�����/�vԷћ�}�1\�+D�A���翿}���椉��)*����J(���l�%ئ"*
��)�i�$��*�����$�&j���(�����gDMUD�EKSMTU$TQCR�D�EDp�IQ3QIT�P�U͒��f
�JI�"f�"���hX����(`�PPD�SDQ2CTR�IIAAAMD4L1,@M3QLUD�UUD�UDCCTP�ECCBMQ4RDT�%Q��H�f����b��=�ĕ�EDPSCSS0PTEBR��5I%P�UQTM:KEht��!ERm���*����*f�i"���b(��f)��
&!�)�щ
	�� ���)�!�b�`��&��)(bӈ�d��A ??����1e_�����&�~}t�kMt���-��{��7���~;�ۆ���+���˥�YX��}^��珧=��z����x���BЩ�J� P�I(�@�M"
4�(H�H�����y�[��7�!�k�:��B~ΣB��L'�9+�Z�ܤ�'ܶ��:��<����}{�ʻ�i��ň����LdDܞ��W:�j�Y/Q*y���cT��Jh���$U�k�c�A���@��-=O����uA�hv���%k��z��_3K����7�&�|=��+7>�Б=�&�4��C��J���ϗ�l����kݟZLu�S�mȞ� _8L��r=@ߓ�ֽ�0�4�j[��`�/@��r`Gz!�p�4B`��f�rwz�9z����N> K6�6;�z��N���^&Y�=��UKW����@�r���.��m���!��<�[���!DK�y/l(l��q�;���n�Px��;�$=���O.�i["6?t��y�wh\2�g>�(`����q��)=�E��^�cH�Hxj��K$!Z�3T�JWS�wg��Tw?��n���htS>L+�lqQW4^b�9�f����>�JЮ�zw�*��,Ȕ�˕Э���ދa����:��`|�#��϶a����<���Q"ըW*Z���� ����@�9��Ygi�AV�z���#���v�`�僸���T��� s;L�[>���X[�'���7�0�\�gq�½�	�����l��1K��׸�ᝢa�I�e�d��t���-��ϻ�~����ԡHI4����*�"R	%%*�R�J�H�!H�"x�{���)�T���
��h�L�)����.�zw_iᮞ��[01��N$��R-�z��A�{����ơT/'�6ٍd�D�6^%:���y�:*Eo�g1����	����c�c�ʫ���a=s��<j`�M#��#�׻�u��K$�s�.�F�
�|�]Qn�	���.~��f��_5��,.d�o�=ʄ^�v4�U�F��a�Ԣ�<S%a�5N��W_Y]�+~�ߙ�W�SAQ`��ӳ�Sp��R%#���S��n'���eX�\�SٞY��0XחO5Ƈ�D����s!|t���	������:���k��7�%�~��۱a�P��V�ը�u6��s�Y���z܀�<�k�?�í~�$��.ǛY&n��p�v�ֺٜjb��Z'�s߂PK�:��5P͚���`0n:�LY̼߮�O�{ܾ���f=h�-�:���eRc~OO�8ϧ]�D�s�f%�}2�"�T�C{�&��可���|1á�;]��}�d���6�s��x����D�	���-�� �M(gf�#�����u'���yBx5�-d�o�_�l��ǔ�z�gX밊.�n�z,���T�d�y�}Sw�xs��L\R�+$���t� �t�%��B���ñ̠`/92�ڷyE ��o{�y�t��]����sU1xx�� �3 �"ʉ$�4��4�H҄�>�n��Is�}x�>�g6s�X�*�C�6�a���|�z_���P����^�]��&�;�$=F��!�#��彯o�ɆC�E���a���-,�9l�a�=�Fk���9��|�m\���OϚ��0�JFS\���R]��E|�����
b���|�3�ǔ�:��qU�U�΄:���DS My+f�eT;&�&�����O�ǬxT:E;�����a	� Ž��f)ݙѧyv����.�y��%6XFPd԰�'�Fu�x�f=oV�^��)u���Z��VkQ�P�x]���N� ��U��1�8�8ĲOi�W�(�k�^n�ueL=V3����r��?|��R��������+�5�a5�$''�۞��D�U��y���,UU�2M����Q_������'X�s��dف��-�1����.�O�$É��U
�0�z�9�twL�����N:Q�v7H�Kk�sP&0�x>G�e�[!b6�����lض�,2�E����w��-T�LC rt�a3�����.O#�g�[
�??���kX��ǲ`�����U5Y3A:.0h����v�"�.���rM���Z�����:Ǽ(�}w�%��hض��I��$��)�Z�T::S�0ŏ7�B�A����S /x�����7�y��݁���v�{��m���i7����;-�y�$+����3���߿�?P�C$Ҩ!J!IP@4J$�P4->����0 uv1D�9��E��A�kװj曯��5�EⅩ���R��g=X�:LK��������I�qfn+�ż-�e��d�tȞtf�0Mc]��I���L�zU��f��Ѹ��{�oP�*�D��d,.!�/���Fy}J����i�j��S�^5���=>�;�_�hK�WX�k-nʹ|�1��*�;F�������xƅ�rnu�;k�C�s�J_j"b~��/]�z�u�}��`�h��b��p�-�/a�@��Ds;@�����X��6�k%'�
�3��m�2�m�e����i|9�!#4]�ñm�Ѓ��W)i�Xi|G4[�|뻩[s�|�{y{,wy���)T�m�gt�)C6緤�j�S��W�v�|kO\�o��)��#kD���,�y���!��[y��,�6�-BB}��A�PJ�CPH�3�ŲƉbZ����5"o����SV"���h�DS��s�Xڜ���vOB�	e�<֢H�90�q��+��{���{*��x�%�C�;X�:ɨFB箈A�=��x�/T
*7~5mm+W�pZ3��$�yw �N2����:|�~�^�͈���^5� �� �Yy���Èqƹ$�-�F��ˉ���*׀g.�^䲊$�LGf��<丛�=����RS\����l�V�E�E���^��=�c����6;{W�����)iRJV��%��a�ox��I�FM��5>��B�),%�.�Ʈ��uo��"z<��5ИI�}�.�w��KUC�^S�Ml��0��:$���#B�ʢ�]�8�Gd[B����a�FO?c��9}M�_�3����0��e2�^b�@���@������F�	\:@�O��|{fb����᠖B�}�&�; K���vT��dת�Z�e��n�t�=:A��x��G��w6r�r�������w=N�)<P�4(��L*��\��jy���:��43�u��ۜ�����">M"^�X�������ӝs��f�I�`�E�:��k`��~Τ��ܱ���/'��\���\0g�A��C���T�m��B�N5��׌�ʭb��1i��ntn���{�����*9���:��aߧ�0��f#_���9�f�W8^���C�p���f�GR�m?Mk�vv�5-�yŗ�^�9�"]���1�}'+�P�48��l"�y�6�|�f�3qud�1��E�q�.�Lߝ�=2�t=1���_�~#���|ѳ_����6ѣ���:�ɻa��'��_k�_���x�dGv9�/�7��*J���*Mï�V$��
�#F�f��ϿL���_���Wp�~C�H�UgP��ٚ6�?��X����������d���]Q�eY���:i�Ó�e�w_���P�����(&F��
"����}����
�;��t9��%���bs���{2,���	I@A�].Ԏ�Ԛ�.e[�Bƽ=�Sb򉷆4g:�B,�ga�)>�7�1�nƴ��$<7c�\�=��r�Ym��ܽ��ȃ�hC��5�S����tS>,*ä�b�h���xk�L�l�_|`�-D��|6���]�Z�T-]
V����8�}sڡC�6l5��W�9��h?�ct��4wZƞ��nd�	M��L��.���.���zǫxi�����,v(�C�<[��k]:����z`^	����6��	LK<'\��5B*�ߣg1�_q�;�W�Ԙ[���k{2�D��t��mdC�L�c@#�ϰwL���$�k����Pr�ވM�N�Q���|��e��N�y��|GܰE�{���`�=�E��F�WZ/g\�۰���v�����L5x�=nZ���=��N�?�Tc�ӳ�+���[�r���Ӫ&;v�ˤb���r����|��h+����s/����z{c�_�}�o�N/a	ng����*]F�۠m���O�)J�_|�S2�--�a�2f���`�CLgP��H����X{��3��u��gg
�3�{,<�oɲ�C�� ��oB�C�3y�{VT*5�4ڵ,�}n���(�O{��ٙ��tբ�ŗr	S�7�=p� ���X���}����y��R�X�D�8L�[�Wm�*��Z������\>�8�*An ��i�s�(��L�v��(�Y3�#okʦ���Ml�J�a@���a(%�¸�n�k��a�����MYcö�6p5)z�!�"���FC��׷:m��ʤ�3��h�>�z��P;��ygs�����k�����x�gmJ5�p��^}:�_e�?p��!��l�����C�I	��LY�`Z�&�w�zc�g��l=����_&�Y!���o��}/�<�����c�:�!�uv����[ͱ��a�k��_\�
5%�[�v"���$xBKO��,�l���^=��~����lVp�\/��2r4�4;%04�W}<�P^K�W)i���>0χ����
y��~��ٽ��zܪ���܈����jf�eTɶ	���z6q=z��@t�w�:r:(�V��C0wV�%���o� ��\�Vy��D���(2jXf�¿vFc�`��d���f�k��m�ݍ�Er�x�^/���H��� F��C�yO6��A8��Ⱥ]����u�Q�y�ƹ�m>�g3��ٲ���S�RF��Ā2�G+�k{���`�}7*|B��n�V�?ygq��_�5�C��N���N?R{Bh���5B�ǈ��`��ٝ����՜��6GD�+����sGt�ɬ.̢�]�D���}���������<��,�|�@�.�X�"3��e|��i8<�A�D��#�| �����S���Հ�����i�}���õE=��E7RF�[X���ȸuC�� �5�����vK�G��T�p��'2��-\ti�p�R�����`�)-�a���l>��?�9�^�t	�Q�r�63+�b��y�]S>9	�^�1i�`�����r1,0��-����Ù�&|V[����P��)�m/c�曯�W5�EⅩ���w=y�3�qxwl�j��9���Y�l�a���H\�0r^}���U
�VjE1�7��k���M�XW>����٣8���?0��;�<H����x�>��h���'�s�a�I(�è�e�Bƌ���m�_v
�=|�ke�'�����:3����LZ�>��eC'��4���`�1�veFWif~�Q�
.��P��LW5�1�W��w9���v�����X��(ͺU��"��A�BZy4:�2#|L�v�<iص0]��tE��sͼdK�Co�z($��<�#� ��}Cw]�wץ�f�W=�z�JҤ��ǜ���0��;���ҭ���%��X:3�i6��P�S}y{θ&�,Dj들p�	b{|���%����T++��O=�
"\�ɚ�)u0V��d�'5�V�c�p��/�0o{�f���I�2!�������7�8�n�������+zIv�%8�5r2�6}؞�/8𱜺ܔrq[o��;�6�k0��_#[�Uϫ�۱X؝ ㅘA�W��B|�3��LF�be�r��f�XǭS_8�r랝��:O�BO"1�D܂oӑXڜ����ݷ�����<V�����-�r��z��Ƭ�����J�|��a�!��f�4�h<rl�M���
��̡��Ⱦl����y\Ruc�JĪ,)�\[`ꋀW�1��-��Pe��a'oI�ن��,K�5Ν~�^'h�қ���EzS$�D�Z��DJ��[�Y�c��	F6�X��sH��}ܬ�'���.��C�k�u˶��Θn�R�p/1Vt�OIq�o�gם��*l;�C������ބG3�	��C�Gd	e�f{*Jz�L�"�	��PMw��vjm��g�љab�C�ny���ӧzg�`��88:��7s��ul��Q�\��,ܤ���YF�%Q��U���N �{�6q�v�$g�?n5� ���^=�|�/�z���1'\^yǩ�Z7ٔ��팸������$��l��/E�뮾���0��*��ْ��ok�R�Xe�����f�����������{��1��U?����ٻ*�"�e��)X���8Eɤ�-��;j6$��9 �����k[⓽;��9�|*�5��d����{��޾��k��ퟩ���_y]i���Zhr��A��i�����_��G6�ba<�ݴvT�'n��n��/tJ��x�2�����J�a>;Bv���,	t�_�0�+�_Y_L{��uތ�2ܻ2K�;[�Dq��r]��m&��@ߓ�ֽ�0�;DԷ5��U�`�OA"��W�|��֎<_Z����]����
��ʖd]X�n�Q�¼D�j&Y�= L˱���
��١�Y�]� �+;�CF��<���C�}���¶nq��a�2,����I��C?��!�5�o_l�����T:&�=_��V��|�d��uN�Y�VtfA!���1`���V6��5��s�rF�Hךn2�7g�.]s�?h���t`@�����Ʈi"ߙȮŔζga���:���^���Z�����ޜ"~��P�E1�0`��}(��T��u�y��<�Ώ�#����Ft�xO����Ф��H��u�cռ50��Y�-��9�����Q�L��h{�G\����<�����ߦ���S�P�U�F�c����^�/w����{�}��W���������G�������o�q�ʾ�7����)]�(a;w�l�ui�Qވ��C����b��Jɔ��zr˂�d�iQL1`ܦ�W*��4�0��s�mӛ��&Xb҈Z6-Ɋm�Dnr7�:�R�Ͷ^���Y��A\@��I��ͨ�^gLrލchي����仳uoF�\μ���gcv�IVMJW�pb�v��[�\�PUp���k���R�;����we�O*c3�3�N383tW3�2�ws]�9V�ٖb�%�	w<,Ί�K�py|�E/�1�,�E͊�ՔE�7HT�����V���Ьl��}rQ�Z��9N;��W]���މ{)�{�Qx��f-@pT�#N|�"�Jk�v�A���\u��͉x*�wᑉW�ϸ���&�r-ǃI������)n�u*4&�'<��a��3���0]GWV,Ǒ�d��Yv9P�7,�{\yJڽj�F�[�\�ڝ%��'oƻ6��fw֭�a ����$�8�9�ۘ�����diz�D��@n+Q�B��6`�=�;uRz^̱}#E�@=�u���3Eofgi�iXc�0�^L�1m��U]�
e���:�U;ۉ	�y������bO���Y�ߕ32�A�ݫGQ��KÔ]K=N����I�N���`՗��=��L�魖;L�]%Z�Iz9����;+C��aU���	�&2��ua.)U�x����jw>���<5)�����ǅ��Gz�t�TM�f��f�M5����E�D`�C2�]qf"���FwR%=���7�����������^h��c�u��W�W+f�@�C��8~��y�ևxDM��>��f�7ko�73-r�'đ螼nb��{\tZKuA�or�Vh�x۾����ss^�;z�P�����u��uQQ�=��`u�1�w{Zљ5��,@{Q�����*4g	�p���y����4���d�c-��-��d�oYS�`S��<31�1��a*+=�^��p���d��k���,j$ei8_kK �vAr�0�>tbw�m�w]�ўr6a��d��
���P���M!xB��<�56�q�������1Wuj�2v^�v��R4A�m�@v��ְb�թ�vR{!�Gp�ګ�ת� �-�C�`j��oE��M�n�0�$-���A�i�;�$c\��S�vK\oy�����}L\8v͡#w-�n0X��r��3H�8��s�.�nJx�T6%@��y�"b+�T�]���3s��p�a�f�Z��䣋)�t�\u|@]���Sd��������_K�y�K��X���U�>��ve�S@W���C��g�Mu��U��F�:��/�'��	ŗ���4-���s[�螄m�r��{�9go! 'ՠ
�x53�U	E�]R4�S�LUF��--!MT%$B���PPR�I!AE!T�KBPh4 Q#I�SQEM-%S0���!4RQICEE+JQQ2Ĵ�TP�CKK�GEPĉACHU44�P�R�E-4�O�#�R�	I1-TR5TP�'�M%T4��\�A@P�TIKAC��>����z��D���͘�-7�)U��q,�X�iX�O4�hۋt�7�%:�^��]N�(�i���=���*�Z�+d"��k�x���t�Ԃ��A�;� �0GP���Q��a@�H�$"� �1�(���ޝ7��u���A�\�x���9w�	-��] �^��;�3�0v�锝ax�I�7E2C�'�T��ʁ1���tz89��E�S�8Owʵi��' o�}ʢ�=a�}]���;"��Ź�/�i�?^�:��Jq�y<Su����u9jw����N͍����L���4$�C��5Z;rsq�N��R��Qi���yt�~d�<�ڨ�Q�4����$����ۇ�3�ي��un�MoK�S�P:���*��z�w:�R;��@�-.���#Xs���&���F���w� ���>S�ji�t�jd�N0D��{  ��uO�j��;���6=Y��UR�UnkW;1Cz�=��u�vNZ@��m���F���Oo�0�կd̖��Gu3�Y�OX�o*}�����w�;�X%~��
4B/>��|/~چOջ!�g�Q~���/g<9սϪ/SA��_X����Q^������v�1.�C����ĩ�����D�b0*Yf�_i���Ѻ���T"�"���_E��lEC�dK<y-->C ���N|��i�l� 4���Է�N�V�������ܰ���9����?W�E�֗�lf�����v�7P����G��{��wh$�"�!�DHXN�dͣ[�6�����fW`rV��V�V�NV݋O&������)�f����ԩ\�L�ѓ��]��3�<�l3$p-�����}Ƈ6nf��KC�e(r�ވ�f|�yKL���?i�_�"�u�� �a����ӓ4�d�}%��g�i�o�ʂɶ	����l�z�oF`��~�]Ka�?0!�K���m��\zz�V0J5���Bk=1e�i=�Q�`��̙�����C��vZ-֪]�o	����
N�1�5l��7:	���;�K��q|�7F�6�^�v~�ߩ��8a=?�<�ĥ1���y�#��N��c�*���E�����j����5Oz�DJr�������#�y�ϑp�G�f�t��v_�ڂ�eܞ�z���.�l�|���*H;J�r�)�J���Ľ����솋a!�hm��ՙ�[ޝб���^|�2����0�Bn��LZ~Y�R	zT��f�I�ݵ.�{#_i^wa����G|F�(�>Ajg�[)ý��s]�2��Z����~��X�9�[4�s�*���Od�wo�1��"��$�y�o�����_?���B	�kX��ɷ���윣~K�:#�[��ю=�Nj�p()�R���2��������$ny��}�N�U��#W�b$�X5#����)�(짂��N�X01��֐����Qsj���[,��࡝���R�h:�Q&_!�ʾ�:@��������-Y�V�S�'��i˺�`ZD���`�.�D����\��i�j�Ja�v,N�tɭQ�����1G���5Ӡ�O��ʫ���X�����J�����>1�9�����_{�����ä�Z:gu��K�Š&�����XHqEM�/�Ɩ�I}O�Y�kZ��	�ĪF�7�A���B(4]����8�wC�|�x46D����U��E%U��Cp��2��l�_�b�i�wO�2�3F����N2^�e�m�=OY�uz�	{�D��V�����``��?���g�RS�;7kqBA�0���Pi�+�\N��xT3�ޥl�l�*�@�r��N�癰:�pf*!;c�َ��/��m�Μ2f�ld�[����[h%Ռ�Q��Ƭ��sn��(ޟXy.2�1<�#T�&�'�g�F��˫�we}S�'��L����n��):��P�r���]qm��r�k�?H�ޏtf�����u|���,�ݯ����vB{$�3s�I��Jue�U��6q��E�*���b����w����M|3"ә?Z��G'�b��t�%o�ǍJ����|4k���^�n��q�l��2V��8�nﾸ��j}:�R6+�[M���L'1��M�u��o)��:R��ԴqzLCs*ec�Gk*�eQyyr`�fܻ\�h���}˘���̺_��.*����n]�6�D6wQ��x	����.2	g�9T`S�k��H�k���yd�:����p�5>�)��3l���l�t�	خ�:�_Wk����x���xf�B����Ag/.3^}Cw=xK�~��B���RavJ��E��!�ue��LF#��ҽS|���"#�$Oۍb� ���B�� &���<�|j�Yv&�o���9%�gǳ��\R��I�ΎeG��XI{����1��lmn��d��8�nUY~���p���-�{dQJ%k����+�=�*M=��Q�'�hN�5~�8?��G4��L��Z��i�7`ǯ�?(e���^��n��m�u*�����;N�5-�G�az�3���4��\-�q��^��!���?0guN�*Y�uc�Y�|w(���$�^&Y�=2�hUي�"h�S.m=�wM�@�t����A@��C�$_���0���C�w��oA��B��U@�Z��Q�@�Ӑ�[�xc[��g�E���ߪ���۵�ƿxG�y�Q)t6\�����f�(.os����a��lo��/\��(��	�o��gO�8�1���Y��d�2�����ثF�VX��;�oVVv���Y��f�VwEc":ݳ�\!�M&�9ϩ��J@4ҙ����F�[���䦼�w���/^B.�p��9�5,�3S4)�}�<�ޥ�Y!
�k�>���Mc�2PޛgO�Ia��軚.�ת������O�o:8urƒ�Ե��-{�2�WB��%GPT7�.:>����=�?yX�q�h9�c���5�:FfL?u��]�)�ѐ�,2%?J;B�>��{��xi���M����a6�+^��dQm c�����DH��;�W�����ħIA`��*��xMG@�S0e赡O=������q����-N��\���R8�c����ݙ%��,X�K�q�YB��=]��۷T5��W0���)�������' �GܨE�zv'�;+���%�C�v��q��Ƕ�Jec^$��џ�ϩx��7����<��|]	7<%!�q��W;�offAK�(qG�������0�ܜK��|��2mcMn����k�t�q��}a�[b����N0,t��Uz���u*�w?ycg� ���Ċ�:����d�;/j���b�X����SM�����J1�����%���4���6ǜ{aV戛 ~����k�>��0_,�DKްDy���W�5��'B�>��"�MkA�wjX���c����!Κ흃�$�7�b���-T	�61�H$omd���A�/p��u�[�������ٸx��Sn�D��L�?����ۼ,�ߝ����k����v�M>�����l�T��~����u�;a�9�;F��$^�ᯋ�U�nB}^v;�g�48y�Ƈ��jj�+چO�7d3od"�rb���8��eꗳf����B�y(�H:"طPwc�ވ� ��4>
,���t�BŞ�Tj����3�����*�Һ	@ =�R3�E��kt�V8W�x�C���g��r���le]���E���z�ui��L�C�K^K(!^�%�<�M���Zfj�n�����*����{������[K �- FFS��z��͵jJ�� ȅ�lPH��3g�J�Ci�S{��'ۗ�p| �z�����}�)&0!mK�\zz�V0J��W���Jl���ɖ��JZ�<SET,5�Y�N��`��c׭��9���
<7 ��& $w�A#sW�� �6%aҁ�����mx���2Վ�)�7(�k����9Y_*6����d9�NT�ac�onB��.�1��Ut�V��N�S��b%:]YrF�[\vO5>Eê����ki��j����/�������@�2C\st���w'J�b��8R�����.��M���f�{��G��)T�=�T��Fq�$$��O�B9޷W�Ψ�[ҡ�d녖�n�Bs�[���9VJ��8��^E�:�	E*��{0<�E�c
z:�6���� �uk�W/k����͗`��L8�)? b)9X�Uy-�aM����}l3�l����f�r�[���8h^mMk��ܒ�\�n9	�^�1i�`e ��*w���0�5Rd�yvީVV[v�tgAPa�|\���8�ؖ\�:�i���U�w�2��j�CYK�J	w������fd�@�h����J��,s�c����Vb�rdO:�R)��5�BO������5l&zYM�k�_=#{��w,�C��ٺGC ��<��y�ק����ȥ��lّ�Z+(�4��P��?1�'cӫƫ�K���!ݺ�������lZ}����	�5�L]h[�[ץ��gmTv�pm9�aC�@;^&+����-@����ɔ�>(��Fx-�W6���<��9[(��}�mH�*��A�������.ŧ�pt=�x8h�y!�=^-f�ȚYo�]�"CF��c蘂�:�m�wO�2�3EoI.�E����c�޺�v��V��������>R��z
J=��L���B�=F5����W_�cՍ�zrd����~5S��t
���5-���ݡ��͜����X��*)�Xh��h�˫4����u[��o5fu�S
g3����P��^�m�����v�d!E)�;K��L��+��!}]�K���ŋ�kQz�kMwS�W�f���=W����鮀�}�Ůy�&s�ho��g�f{kX�gNZ]�X�2`|�k1Q�˃�x���!�Z|6粛�����j��l��	��	e@%ՅW�b�YN��[���]���g��#�Q�N���\q�A
��g�520K�12���,2$�%QaM^rq�uEê� ��(��N����}��,ܦ/��v"Gd���	�T������Q�j�QN-�-�ȶ������U������I�P�#��p�!�e;r���nt�Hԩ2,�1Cbڋ��P1�s�����l�>T�?��;�A��.�R�#ZD:	�	��<���34�egUCO�T�z�#6Ⱥz�C#�U���]�F2����s��%�r�+/��ڑ�=�S���Wxظ���T&�2ƺ��e�dg9�Ք���ܢ�iIcC�Ӱ��ٷ���`/�@�����9}�,��$�}~�_�!\�q�3�ΞeVְ��v���V��3�i��O�)`�o�l����q�*��hT-Z�Z��\�T�З����'��s�0_�z�.����RC�˿�j�Me��3�u��X�~�)9�z�WxL^$Y�A��,�V
9]�1�g�p�1����J�.�,l�¤�9e�_nu�>{bW-���glZ��p���71��=/)|����N*�/]C�����t�R��[˺a�US��4�v����`omĻEU��3}�Y�Zu�8v�>pZ�R�m?M��ݣ7�Է5�0��[YM�i��m+;�<�3���@r0��m��T�$��a.�w$��q�.�L�~�As��O9#ì�{�#��;>�b��?j�xyCC�(S�P�s���D�����J��(����V�E£{�_I@�җK���-�<S�p�`�������O2�oL�0�L�>�[M�J�kH�\����t�K$!\��z�F��WL\:��L���}��8��tC\�VFY��M�B�5�\�z鱯�FBױ�e^�t)%'?{zq����s^ئw�Hs�[�v���hV�ȉ�i��������KsP~"Se�!2XdJ~R���#=�	pP��4K�����´�<2O��[Iq)��HH��;�P�Jce�S�	I`�*�SϬe���.���d�=��	����[Bt��L��h�1�G��̮t���Q��n2R�Mn�j��E7QF�
�\��s	����3d�&��L�^�`$J�@�xg�|B�Y�-E��%�Ro��+Wfqjw=
�eF�J��o^�kG��J3�����wo�qPYGԷ��,Ҧ����S�;��h��WM�LNwך�����Q��{3���ؗ"el��0�Ϋ�9"��:p7#�\�p�\�AO_M����[f�l���2'~��EL/�J.�s�2�-5�u9j�mx�P͍1�t��y�ݲ�_WCv!-4Х`�(qT,��z�Z~kAb��ߛ������՟��%����2��Pw+΋S!F��SIՃS�9"�S���w:�WC��di/N*�9�[�7i5�7�A�E��`c�:��ji���je�J�aD���E�(%�S�5��#	�۫��ok�nC��>lA���qwf�M~��m���\eRci�����S-j]u�W�ֽ��S%�nK2�
>���<<���?��SVyXL��u��|�Hݔ7ii�{�����s���Ή��z@9��Z�V c=��k���F��)^�b�8{�j��E���-��ʃ}#v����A!� ��H�<�Z�5�k��8S��~0��='au-&K�k�۽cM2�Ʋ�'b��wH���T�;$�4�W�Iwy�s�vOKk�9EVz�O���{{�W���g���Jj�����T�y�ɛmH,��eTɶ	�#����/_������{���w�������w���{}===���
�hD��xPe:�I6���%��
��պ�=x�˂������d�|�&ؗ��9��s1�+3�۬�|�Hf���0n��#��h(��F1�5M�,�u�W���jX�9rE��+p���pB�����%��ɭd���ewm�Lqf'����jDkh(���+�k`���ہ�_ C�r=2��׋y#�(o�'Xna���9�oe�3.��rGa-v'���I��Z@��ui�:Â� ��j8VZ��yp
�[��D��r����`�,tC�a_OzCO��e`W�vEf��r�YC&9�|������ӗ�-m��]Ƿ�E�
�S3�+r��W��c\�A�v
ȕ�<�7'BB��&��f����E�1�zx
&�`8v�9�V��ɹ�tAM�Uu�j�#�cꭽ����m�ޡ�n�i&�8�u�B�W[�s��W]�CU�KBҩ4��/;va��4
��ϵ>�ao��^WY �_[y`���̶>Rf��yo��J�&���(6��ۙ�C� �y,Zr�0��2ZU:\���n�f��@':��33w4�AEg	x�}\,� 2���m<�n���d{v�x�|���9�oi�|$"�@�92��>5v�*jZ��,�^;V�p�����&J���3�n�8:�z���
̾��5�rv,�R��m
��/�Lf��}m�"��r��:��*\o*]E�6��M�k�[��ΰF��Ww|�f�˓2�w��繳��+{֭�o1��F�K=��OW���gAU�ss���z�h5g���+om��E����ݷK ̃#�AR�.].�\5�xI�n��t]��n���e�t�7@	f����5b����S��3*
�qڝ�v�4�L{z����d�2e�k��4�Ԏ.f�Y]�q�&������ʶv���w"T�������oد�P-�{�%@�Pr������P���s���0�(3{��3���lv���G�bs(ޓ/0>N����Wnvn`�Z���(�U֬k�'Pu��d�3��1)��y�놅SD/C��6���+uD��������F��e��.����J�gep��!�~�ʖ�ڏP����i^��.�&v^pcn��oMK�C�(4��UT�,�A��]F�L�i౦��C��8�9:$��';�	u�Ee�P�.��ҵ�,��vX폺�Mʒ7|mN�6�N�V����-%l�;^߫>S�(��)�}-}:IRZa�5�� V���h�d�&J�aŊv�d'���)����n=�Z�-yA;�ZƵ��]�kFʕ�P ]G�6�Z�%{ڙ]W`����\�'v��\_�z$Yqu�"�_6[��.ҡ��*ɋ���b�>���z�5�H�:vof��U����}A���;�w]�n�"(W�4�
D%#AJ5��t�G��B���4�R�����i�i:ց;�@J%- ���3�
9�%�5HEJR-	�BSMSB�s���	)h�)�e\A�IIKJ3' ��B��:kĎ��h�
���(䩡�"���"�Nl���h�9��iu��$$(j�
i,��>]��{�~x�^�4MՕj���Za�u�^�u�i�9<��c*9�v��Kqo6ҽ�����5���1�1�nҺ�>�>��;�|{}j���o`K��-�2N���S6�"'b�#��M���;��Wa`��{��}��Ҷu�wFc׭��վ;�
N�" F��EF*��^0r1�Kv(g��P+� ��t��ebQ��a�Ň���V�C>Oț��#��عhS1u�͋:�A���Bޕ�^s�'.��)�$i5���j�p���S`,��0��5�jk�sѬa�����d���:}�&H�i'.����5��L9�^�#ϷL]
E��Uqc�u��X/Dy�t�s6�G4��S"�6��LZ~Y�R	z��麼iɃ(�"��/]֥��$l:C��8}xeσ�曬�\�`��Bԍeq�owL�Lx+��0��Y�U��-d6~�/^C�Br��z��W%`Ԋb�͵u���Jn6w��k������Ȯ�oW�s��3n\[�6���ǂ�.�B3��TS<���Wr>���|�j!��}���� i�L'z~���?W?N;��:�G��
�	����<v1��-���ܛj��0F �s�S$��Tu5Dx��K{���E��m���:�}Xu��m�ʓ7fet�;h`�39+��k�['�;Td!�[��U�����еq)������s��e�o�Kە�n.�d��"������:�޷��߷-Tx��nRpHNf�P��׉���Z�{�9��&��ڧqY�Vg���v@!��"&:�mH�+�Cs�;��P&h�P�.ŧ�`��DYt"�Q�?v����6ךw�~����/��h!�lZ} L$�-����fY�h�7��d��l�_�7�҇ޘx��˾2��t�?~�a��I���1>���"�Us��ݬi��BA�d�ti�O8R��
6vw��'���ʃs!�g�R�8��0�@cW�T�<�L���b�+�OWl'RU^F�\��+�<�+]cqr9���֠K*�]X�F;��j�3 �]z�Iq��5Øήw���f����i�x��&��I��C,{���U
P���չ8�T\:��qnw��0�+�AΨ������f�&�,]�!ۆvJnj~��=��N��BՉTS��8���,R$޻6��ɹ\C^�^
Kz="	ƯK�L9��]�4�Θi�I�g	�Kˊ��f�s.v4����"����_��L�7��X��>]_���bYP�5 vT��>q�u~�9E�Kt<��`��j�nj�Z�غ��7#����t}��1?]ڔ��vi�'e����xqk�*��a���p�O�;����҅;����x$�ΐ�v��R���xLʴvɈvԏ��0n4��=3��ȝ*�E�I��[ ��#��53)�$|&���+� �8�>ߔC�ʒ�@��>��=ʢ�.��P�]��P��U��~n�m��ǵ9�R��)���j�'�	IcC��"|�D�%�� ���_�6>=�\3K&�A��g��P�;5m� :�����i*�
:y�*�a���Z�=�x��}n��b��nmf_4���v[�x@ضU� ���T-'��;���{*	{k��HhN�{������j�]�����	�6���uBv]�׻h���@�~����њ	�ng�u��.g�֫��o�ww�j�@����`xy��|E(���fT�B#�Y��H���Iv}l�i���aUrx��TwY���f2�ئ]�B��sW��`|<�г��1ӳ��u3��ӪN8Y�6{y��tμ$d$���H���'[.x��9���2�.'љ)=�<�h%A��`�3�B�WoL�ތi2	���B9i��t�L\:����H�����Uo��{6;c]���{4^�TcWX��kj�R��Z��*:��oN0���s��坍���HLt/!�NT\�'9�z/糥5�=a���JidV����i=Ω'6�e��^h�� s$���u"��̧�u$��r��A���J+Wn���S�xd�p�Cۇe4w2���� �����*�JEZwx���Nҡ!F�{��n�zN�o63�8Gg.g^B[N���^i.�βV�K���"�l���PY^6->zQ���`���Qn%V���7Z�t��ᦞ���ҜI|�	��ñO5?!)�g���w`S2)���x��؞��4���+ېW�&b�ڶ~�<�RĜY�$3�`�}���v��mwu�Wmw��fѻ}I�YC�Yp(�aA�+�7M��V��2q/���E�z�Ք|�e	�v*&�:�筐�ZiC�Ȥ酣R��g�\��7�r��p��=4 ����S]7����E��joۃ�>�1m�*l�*���{/I��g��L?5'� ��ƔJ�����l���;�2�!1��4�Y�����~%Q��Q��o��w=,�͙��=M�i�����5��v������_j�ښm+����*�OJ׿%����Ó��FD�I�1��w*cuր�g�P��&>��掯�x�ٍ��Շ�)��Ѹº:iNƩ�ڊG/�U�$�zu�#ުv����dA�� p0���཈y���6���<����g��\�K�p����\�E3Ԗ�je��S��?B`�(op�t $?NH��d���M.��~�v֘�NUW;�DJz����I�[B��h0&½�7%����f5��fΖ����Q�	�K�z+D���f��2�k4�r��E��RD?�}���]�������IrC�����lZ��!��D�����o4�%�q��x�QU�no2�6.~W��Fk��&�a���l�C�"=�ӱm������+T�� ق��r�]����C�lsL=����^=��ui��L�]�XK(!^�%�Z�m:y�6�;
�2�C�Z�Z׬Bid����suS��nL�Pԕ3m�2�*Y6�5M�4Υ��)���=������K|�_˧Sֽ[£"��`qm�輈���yV��߸�ߌ����J�%�|������5��6���{�gXQ��z��x/^��x(8"X\� V�#���y�v|o��z��¹�r��Q,��������՞����i?�y��9���4����̻��[M������<��]'�&f��t�d����~�ٶ�>EîT�;l�����t70mL�B�;˨��Gl�'$É�I>I�W��9����ۧY��N��k;��y��F0����9m���ۓ�I�S6�9/I��oxO�{��ɞ����x�J x�0|޺ɳ�l�{Ui˜S�.��\o�ex�~fN�����M���	�� X�/s7N���U�����Q��y~.!|��6gfV"�P��B�	U��rSz�<��g��%tsqQS5h�������K� ��Q����z ��~q�3�[���v�e�;#�G�J>R���])����q���^c�]�����j80zЦ�}/���:~�?k�j�]��˽C��s�5"��gd��f���vQ�z��RԆ�)�_��6�j���U,�[�ͳ����@!���v�E��w����7��f�����-X%0��x�Z�ǧ���OW��:�G��d4.)]��@r.�i:1A��s;w��x�1~�w�?P;I86��Š�b���r��`��B�7����p�����1񐉎��9N�*�5l��&-8E�5���,Mv8j�
�2�yL�qk��Â}r�Oz���h.9��+}"�m�H~�H��������$n�,�����߻>����茵������_�
I�bd!������W^�cn��3�l�a��\����w�Tpp��A�PK%�%�f�?n1e|��IX�``|�Y��غ���7,|1�-p�BJa�X�L ����4�&T�V3�^���{Q��p�'�>onI�Z&i��UM���z{���p�M�poiۭ��S����u��^\�����Vd[�7(��*���b���V��B����^d�jK��vn\ ��Um��FG�2~�Z����n��h�8]%0��{�t�V7��Ҙ*l+���t7{ ��)��='<U.�ڱX�p���s{z�
�?�u�ؘq&$��4-���;�Ox�ʿs�.��:!j�JĪ,)��[gT\:R���XH�Ō��u��8�9[��Լ&v܇n;%75 �	�{1�X(еr���Y�:�%�^>����������ٍ�����2ݹv���L4�R���LW��H�
dEI�|�i��n��u`A�/A�-ᄁ�<��4�;��L9����@C,�튈�DR�໧�Mws�[�h�d]g���Z^�=5ʒ�D��C�P�r��s��݄Yw�(��{אER�I��j!s�u���m),k�Ӱ� ٷ����l�tܱ�nc�Y�l����M��δOr�n���~�j�Y�bN��T�,��Ua]i��i�V�cP ���uN<D?W{z�,|;�k662~e)��u">����%k�-е�����؝e���?��10���ݢ�P�`������G�����;.�hv�a�@�T�?Mk��ӱ�39AJ��t�m-�B�q�W���"O��O�����8��ʖd�_t�t��Qo��cB���Ke�2UĽ�ѹDp�Vf}�\˕y��wF7��\�Q�S%��K;.�w��ʻ3�y�{fN\.����t�F1J�ʋ/d��_�,��6��
Q#��qهnR4�/�5i��:��]=�2{:�3�]��PU%΃0����"���tD7άl��ב(��Ӝ�t����Cj�~1hT}���+�j�?���y"�VF:�de=M��W�i��Q᜙��xCT�C�J�NC��ʆ����π��ˎ����^�kYyHݩn����|����׶��ә��P��	d�;�O�m寍����0(���RGo�w���tXվ�q����DfMc�TcR�9R��5)_��ں�%G\=oN0WE��y�1�[�'����SW����G;H[8�\�KsW���،ȅ��'��4���B3�[��F�v�޻#P=;�X�o"���1m)ėȿ@Homx��),�D&=�E򈋖�V�y�,ƞ�ݮ[��0֯B*�����e�'�o��[&H=�'����^^�jusS����g�L/r�E�x�K$�tS"�����y����ց �6LB`��n�s+7)������c�3ZD��0��]0�jQu��e^Zj��S���^<���6�
GeA��{0��ɚ��^��a�D����*znE���.��^N%�	�y�m#jo�5s���/M�!:0�ټ��l����=��o?^�H�mU�;���O��,�_un3j�|��V�����kl�RC�v^]+Z�xl�;2rC�X㹼¦�9v;k/l)��U�Z��E�µ���׮�Rk��{uhV��:����e�L��FwY����U��@G��-"�n���Yu�T�Եm�rTa������sư͊|q[.#Y,�n�h���1��î� !�p�01���f�T�Q�8���0�OJמ�'�m͒���(��#o��Oܳ̕mvB�+���X3�a|�Xh��Ǎǡ��l���2*�"a���sK�c�b�§�J}:�	��;p�tņv3���
�(SVy{���W��(���H?H�MOKzC2�;%���^�H�v����lZ�X�c��1aO����T.�	��6���m��Ec����xX	��F�ci�	@� �M;I}��f��U�l�S�7_�q�ێ�?�׌���!�z��ǳ�#[�������e+ܤ��v���2o8���n�l=�q|<��g�P�K4>?�R����s�DSjJY�2�.�R{�y�E�T.�/�'M�C�G���Af��ъ�?������Ŵ�ȋ�OR��	_�b��X}�hP�����ݮ���Pd�Jx]õ]�2���k����\l{�����g�>��"��[x1'F��9�uk&��%��S9��ZlC;/��`쀐5�m=F����X��}t�n���ca^�I�ѯ����QFMxI��f�\�¹�Sp$�z9�7p��F��4S���b0Xʻ�'v���tp�!_+u��{�ܾO����>9Qf.�q��K$��FT��kw�{l`?���J���f*���}�+����	�f�&-�Oc ���A�%:O��Ju~�S(�$m65Ԇv~��mz�N����g�ݕy��=�+� ��b�!\�u	�Od�#�L8��4��s���%p[E�1G1��oz����+t_GR�v���z`����:�h	���<�^Ω��M�������q(Q�Uug�܅c�׀P�0������>��r9ñ��7����l�9��O�m+C��m�^��v������Rq���D��>3��;�������\���"7�R������^�v�&Uc]�)9kZdگ����Nh
�'sY�?�]�s��NSv9�[ϗø�|�J���T-Z�L:�Ʋ׾=>��~�b�A��B�v3lYۊ���wk�9fp�J�Vl��l�e�>�i��@�$��s4½Š�LW5x�r�t��Y��e�R�y8w	<3�"�� �`���ԍd���sώ�	�.�8˱n�|��/w�������{���w�����|G�����ܬ�;��:U!|%��L�kL"�������]P걢]qtF^�/�-� ��}���ڝ&�-gdea��G�7 ���������O���u�ɢ����\Q�d�6���`�ܬ�Kx�m��u�A��UV�g3��ĸ�T'F�+L�=��Y� ��#]�"|�:i�1/G#�E��i�/-�P�� A�/���Wf��(�2�V<jb���t����te;��ڝ�A�vG�k�y�ǵ/IH�
ƛ3�u�r��;5��v����ȃ�����{�I4���>�D΄.��P�����wK8�壵�K�W�`̔�-u�����Ng�ǏP��ce^kz2�)Gd׬��5nuw0��6
���҇Z�[�P�O'�V��"o��5�ʺjz�Z��a�\V�fl�\� 2���u�R�%Sfq��{q���S��l�:-s�xr����θ�ni,��-��Hd�3{pq���K����5�:�\8wtl.���M�;J-�o�%�Ž;K����P
T�ݕԞ����r���B��W�
ޢ�U��jN<렅
�#���nQv��Kk�*#�w�%��C� z,T�8�;�3��c��H�{	A�`�u��n��r�(e+�%�i�,�±�;Ш���/�����@T�r��Fɪ�hIٻQ']g`@�vbt������v!q�Nb��]��ⵌ�og,E�N���5m��ܾX"Sj��{�y�kz�Ȃ ��:�w�k�j����9����c�gi��r�x�+�?:O'���OŚ_��1&u����~g�9��i���l�	f��4��e$�.Y;f�@ٚ 4{l��`x��|{^���+��y�SF�-�R�v��$Ķ�"����t�%�5ޘkN������J��Mֳ�u����t�p�&o<�#Y�Q�î������3D�4�H�	�2��w4d�q���1�;6!�Ÿt������[n�	�ƱE��L]�h�S�Y�R� ��.-jF�K�a�_omT&�V�Rĭ�R]ɀ{hb���w����
���lJ'p�M��̝��%RqZ��Q(w��˜���9�1d�FWQx,��&�\�z&S�X��3(v���PP��k0�:���ϟ��������i��x�4��i�R��dؿ��_v����͖�;d�z����X����<X���i�oQ/^n+}�н�5K�7ݼ�T��	f�cxp��Y���Λ�Z$�1Tօ�D!ȅi���y�&hV���A[4OdN��;;�&�p�W+:E���ڸ3G_\I�hJ:v�U�΁y't\����� �����ck��>ōoh�,�I��$�%^r�.�;/���ߞ�ޖ8�}ԝ[��h@�E$�"��k�[n�m���
��c��"/�X�H�U�&r%ܕ���Y�n��g��o`g��~���D�C95�|��9x�}�>}�AMSB|�!�t��%#Ƞ�5K����s�<�TR�R���s�4hДP1*�8�4J���@U-RD�CJQ�HRRh]�-ӣG-P@:rt�d����j�����(���� bW�� NCIA��r�\�E@����K�HhEB:M	N��!4�$�)���4P�@4R��x��Vy��([1�b@�m�Y�8$>��.��{��y�/x꥔��1�k����;[}ɋT�-����e��ֳcuf��XrG�L�v�) ���'�9&$���Q1(�I��H������S� ���S�g#ۺI�"�(��HXw�_�KO�`�x�E�)��_`�v����fY�h���m�j�fj��\JWܫ��Jm�2S�0��ԟ��6�hl�w�ϐ�`��Ⱦz���э���Sx��dU6O'�2�Q�8�vBX��BFq��l�*���=;�.2�BN�[/���f���ᔹ_=0B'$%s�X���!>��A9�K$�m�Lv>5��sB�3k��os��G,�{�Y��)
@��q�Ā]���|u���2�C��i:��P�r��X[XU�����a��ێ���S��¶TC�}gR!7�k�u);Ud�p�vG�75�Bd��"S��˻��=��v<+���9��r��FN0��m
�t���~�!���n#���Fw��&S0��M4��A��-+�u
`/S)�Eq�n�z�o'ېA�C���1���!�&�d3�����2�U�R�Z�J���Sl���x�K�ӑ:��~g�}�A���t�e��9�8��N�,YO+�F�#��I�Z��Y�I��RX��v�٣r�ckz<�Z��JF}�L��~tg2W�'�R#=Z��Oz�٧���9�2��M ��^�+���X�=��!;^�n�+�A���Y~b��j�#�䡓��n��¼D��<x�z^��V-Ъ�G��!�k~]
�Gj6��4	�J�\��.u�o;�����^�_�^k2�Zz���V��f�qG�fTX,��TUְ��}j�=�~1�ӢC!��/*�WF��<ŵ��ƇT�m�2)r��-qŌ.r���_����	R���E��ok�́{�F�	1�3��-0S���w�Kni�k w�$��GY���x�7�'n�3̗1�|�h��$�0���!�M��fI���Y��������}��;��`�1%ؘf6�	�v�ly�3��k˽&`M�Dip$C�|a���u�z�="�f�1���ƾTi���^(oH$:N>w�������Ϩk��<Ĕv�p|��g/��7�w~у�H*�|�Uj�{v1�ِ�xn� �y,��F��.2�7C�:�{~����U*�s��\ΐ�a�����K̽���NT��jR��0�*���J�%G\<5�
���#y�	c_S���u�,�8Bli�0�|!��<�^[:�_�jX� �D���L��z�1ze�q6���z�{m�@	[�.��u�z���{gh Ŵ�8��B`$'ݕ�{� ��F�,Ɩr����]�S�h��,�^���_�(�$�E�'#P�ܨj�N��WJ����+Ev�IwL���:(�.�U��F�P��q��d��n!��������b���i��,�:�}����vN����γ{N�sw��,��G^�=�}�>֏�x��iI`��B�b��}Ǆ�,�x����(*��>D�ѭ�B���������@�3��e'E�'I�)� �����=��z�֏H0͖,��7rݼ�W��c�v.a��5�q�z;(��<�L4#R���d��7p1����������E�魽�W������l�o��K�܇�*��iC��eWC�9���PXחJ��YtA}����ЩVp��!�N@{�������T!ƽ�4�������w�*�=Q��FXgt\�����U^l�ֻ��s�1�zp���:�tz:�����j��ˡ*����6�U-������t��IG�{
�A��m�s�s��ls	��P���;���Bl⇫x{UR��9����j����:�xǣA3<�w%�ы^�%�5���O�����gQN+�r����z��$�\��m�_�����֟\���wX�c#�]��U��J^�mtg7>p<� ��'�$ͧ���Vx�d���;���	�e�,ƌq��z���^���4���Gw{y���@�vF����0�]� �A#�Qh.��G��oe��g��t�C�~���L�aI�3�:�|Q�.���[n�]�As#*�ٝB��3��{��C)�yi'�k�@��﷚�C
��K9Uuf��P�������N���]���xĳ�M,�:gj`~��ǳ���sP��L�G'XK( sY��Ƅ����þ��N�זM��y���yg�X����&�Nn�}<��3m^ԕ3iE�������I�݈l7!Jq�2�r�-?{��WH�|$[�!�߄Tzz�V0JޫH�\��9�u;�f޴�l/i"5�#��2ډO�J3�(�ǡoV�^�o������%��"yT]�������1�!f�*0�5 �'^'K�X�F�]���Ʈ{gO"��ώf��-9Q7b�X��q��(�v�>ب,�@#;$���Jt�D�V�^uiMmprKMH]:�[�FE��)�A�kO((����ц�%{(�Qg��d�����4�㘤�`�)vf�F�Sb65fsS�:w�0�S�屼���~��`A�x?�����Ƽ����ϱ|z.�ge��.��q��e_��s�/W�3L �B��=(�rg�ܸud��q,�in�j
-���ӎ��j��jԍe^J;��`�Ļ�lc;5�_�?s�;'���7��b}4������.�;��I�+2^�Y�M7ū*V���uЦgu7��,A������7mE�vb+�h��$����0h�c��}գ.��(���-�R�Y��f�<�P�RFk&º�G�n��&b�y1�A�Z�q�A-ҭ>��̊�Jn�
춴vl6�QD���߶���*�����-ai�oV�|ja�/b�٠cp�}a�]b6\�f&��;<���i�u/Jn=R)r�L:�x�Z�8������9e�`Hﺝa�(���/)>���xW:�0dp�0Ali1OR6>�i��a+�S��
Z��ss�+�؋��3
cD^�<��� ��q�� �,���3���ʐ�+����r#,���ӫ�cԯ��ю���A�>?��B���������-�M$��؜����v6��S�:V6�}���r�����r�v �5���6�v6�5���R7q�4�Ȓ��D���Խ+��m7�Hq]�C*�Ԍ��{6ʇ@�t���@X1�YC�*��6�MŐ�M�aݪ�X<T�9���>7�еYR]X�_����s�Ǫ4�#6q�]t(�m���9d��S�%Ĉx�c��[Dd.~w!��'LW�*�O0�JtA5R�X�V�E�,�E��[=��ޅY�'l�8H���M%�+��=���~�E�ɳ�^5ԣH}ݕe�m5����LlTMjk���&��t�*�lrZ���]��$U�̑�|;/�U���`-�ȋ�ԩ쬰�-kJ��}����9 �|�#Ǌ�����:J��z:�v3��z�?:{�$pv�k���GN\���Կg�5��&��]0��V_��#^���.U�j߽�g������~3S;�A<�Xn�I�ƅ�z���	0"1���?P�s�s�0�I�����u�����Ԫ��O�&)�u��2�xN�sӸmx󇦄,t-��ʅ{rO<��<X��Y/ش6B�-���o��
������Oa(,iq�a>O�ێ��Q�q�7+.,�gf�[f��65/DȽzv):�����d�,(,��U�g��*�Z���xbr[M�խ�V�p�8`�A��X:ap�7Vԍe]��aՀ�V��OJ�)�zl}W�@��wS����oL��rd�����4ו��s8?��69����fn\�5{
T�X�(o2Yp���[���/�UӒ�1j[��/���s&C3������]c*�������|�WR�]Ll�rf�=�+�PF$�Q2�u虑>:"��@�r��yw@���_cv�`�m���W�v���5�o�l
U��7�u�E�� ��ǀ�i[N�S�v8f^��TڿV����ڿ-�'�,G7"��ͣ���^[s�9�x�q��dCh�.C�.ـ��Ү]���*�})7P���l��IW'7&�_m��V�T�S]K�+��gһ{�g{t#l[yZ�B�����	<(�L3o`Be�V;;���������o8�	���µ�[�����~���T>�$!C��4���LԘ��N��j��u_�Н�輳ňL#�:.&.�̸��ʖ��JB׼0�*�t6®��-��k����,��N��sy���,-0���峌��԰��Bk�n&p�(�)�vͶ�a5��6�ʅsܮ����M�c�f
VQx<���!�Ǽ ��2U��h�Q[�
�1��j�
@��K����۹L�M4�H��߳B�w������8���w��}?H�t����dx����N�nx
+tM�����u�`���/i�6���Mx�7�s��0nnHө�z�2gOw3�8}�7m���1��Z���q>�Z��up(�MZ�3D_0�ݽ��3Z��s���--���0Y�c�m3�mG���=��^���~�m�LN^Y���� 9�mt�`�����`��lΪ2��Ϯ�^Q��}Y^h�t�L�f)B�N���IŌv����^4��!u�m�M�����=RR�9҆�l����T����ƪ��M���9I�ij����[�k���]���eך>�XV�=�e�:WWq
�۝��س����/�wt�L��g����>�x���?D��T�2/%>�����0b=�,.�/OЮ�U.A�i�˞��>�Ô7���c�а:Av<Y��6�~����eMO��/d�uq������4Z�l���|!r�*�1�롩�z\���W�Ѫ�v,9+���֥\�w+{��Q�<T6rL�n�k�ay�$H$O5>;:��9�0���ǸJJ)Ԏ�r
��+�������9܌t�=��4�V�Ŝ�4;$X�}�����q�?4YŎ��	��Hצzz��^��I�����Lܦ%��;��� ��T�Ƒ�jE�(�j��0�{1�g�5>̇��zѣ��5GB'<��T���'�i�ɹ�4+�QW�e�Z��n�����.y�{���P*��)RFUB�;Uz�Ӝhܝ��v�mj���v$��PU��p�����"Ζ��*"�<��$Z<��= �2	dX�p��׫}��h�͛�T��}���!��DE���F�)��r㥘��/ֹ]t��"=Ձa�1-�ìf�Ъ=�6�	{�A!���}|{�^�V���k��n�n���h��U���� �ڵ�������Ҽ�'fr%ٻ�\ӏ��*���A���D3�����=Nq\-���pQ�չϝҒ���E�d�q����v�=9�{#��^�\�f<m��ӗe�7mz���Q�[M���/f�Λ�eO��T����'ݲ���\���F�F�?y�
w�uJ�6+��d�Zs�:� �$��]ڱ��n�d��`�eOJ���ם՝]Ú�37�
Isr{��Rͳ&V�����ySb���-]wz���wxjHnC�����#p�.Wŋ�{��A�l���i5�`��Gjѫw��`؏����va5�dv�q��*��ޥ�FcY�	���x��6N_OPe�mӀ���uz�Vp�9e�'�7mCI5�/}F��נ�lR�h:(�u���p���𔍊�Z:�+;���[4�ƢFrV�!r"R"4�@喫Ȱ��C��Dh�zEZv����p�?�M�*>~�=��r����m;��5v�a�<ҕeζtz�A�v'�=�I�S��<x9������g�d�]C)�EY��v�Ua���bه�1�p�j7o6��50;�G�����ȯ���۩����굝�O:t�v�WA=2�"��um�5���sgOQ:��̸��:�%U��p��Y��цw��8�v��{�p���Z�^3[�J�x�2/RW���"��A.�=Ms�����f�T5�z[��;ަXň�n�5-�u�G9
�ܑ�lɖ��M���Ƿ���{z�/����L� z�.a!o�m��4�t�:�`o*���Z	�������.x�y���[����t����m�^�g^�;A�qxٺ����4j63���:IXn�R��ϛg_��9^����u8`q�7QsFO=�>0�P�2T���J�Ҹ޺S��@;=,1�M�Ӵ=�^e��/3�`F+���:Dg��9�h]U㋢h�T�@P��)���͓�����Cnǥ������>t�����I�F0��r���T��)j�$�(ڍjl���Y켆�Sb��}˫'�Wi��Y�Y>=>O�ޟ��~�_������~����z�|�]}����6(���3D�;��As�A󡛦GX���6�����+K+�7OU��7Aʂ���F�����-��d{�D�Ur
���뀻���ヒ���v�����n�6B4(Qđ��O-f�V
�c�4��e:�7��0V��4�����g:���[�GF�ݓ���%�N�wTz� �h��X�c�vI�����6ի���ʫgQ�z�Fgi������"�7���B�
�ݮSMbs3��ͱL�&��׎�mĤ�T�Y2�A7ؚ��fm��N�+K��˥Yɘ���H���m��Ͳ���w�2��bʗ��cs�i�X����V�!ʣ�e0�{3v�Ç��_�뷪�D׆R����'L)Q�9Y��;5p�ti���6Վ��;~�JמF6F������^��:�_�j�ؕU���A]9��OGe����׳�]eaG&��\Qs����)���q�� �t
����c��{4���)�\���ىf�x�"e��VU`������le��G��No��5j�䘃=������������y����F���gKd�:�p�
;��46t�j�ɸ�n�e���flKy ,���{�O��`�l�ɔpC����`Q�WR�ڽ2q���n슱��wٽ9�����fR"c��a���8�i�J#��7�%�',�n�{����*�ܦ�ww�����'򮣙��B��UACV1��hѧ��4���_g�מ�o��C۵����h���2��[�5O͹M[�����~;:E:aX�+�ɒ�W����%sZ�
�@��(m�)A��;��b��&"�5ėͩ�]����ef+=MU�ި�������qk٢�bo&��{\�R�O.ō#h쟫(@�^�Iw,:�,�\�py�N+������yј�4�EL�`����0Un.v�������l���7��X.�MRKVEV��$̑�����A!:���Cs{��=�����-ʥj�����1#�dI#�'�T}��b3C�R[Օ��{��<:N��1i�Jnw�WЮ��cu������D�f��9M��7.>�r��a�Qx*��i�bR
��ǖ�v*n#	�E��Z�u������w�
��l��>����y�f�u-�nK�4�$�W�H�Mm%t�pFc��#Z��.�F����mV�Z��Wx�V�}N���k�]������4F��/l�xԵ�0�`��EZs�Y���.����əD�[��*c��eV�ʆ6��ׄe��fѧ4�ou�<*,�**�36�4k*��LƦ;�٩ţ��i�(��'Ǉ�7�!��{㲴x���ݐ������g̸5vk�U$��7/KÚ2rTZp������Z�s^��&��ٛޒ�����N(� x�Ҕ��Қs*m���SK�A�Jj��4��*S���Ms hh��(J Ҝ��4�JR�@�
GE�t{�#�s4:@�HD��	AJ�!�r�!@4�GE.��Ё���˒&�4��Z��6�
�<Js`9��i%ABPhJ�QADK���:�)�k@�ѥ��������GꐍN�ť��n.�/�瓎����f��B̍=�P���2s�f3��r�0�M�{F��W\�/::���ʛ��ӆ����X��91C�+���t�ks0-㳸ۗW���do_'(c;�s�a�a�8|�e�o��5&�Q�te�ֈ7�=2rA�<��H&#�WN�s#���1.�P�t�����d�lu<e*�M�W���3-�{�x�A<��P5��j������"g.o)�A�L�ȍ��L��^�9���ă��]!"}��\�����9�V��S6�ݑG��2�b����^�����Ċ�g�'}�H��ש����'�Έ#Nǭ��@\H����y�8J�J��੽��x���������(��J��*�#�@ۺ�s`U��n�\� �/�śwc��:{0hQx�<�!ҮX��L"O$|!T�w>�ei��:��6�6�%��M�h9o�7�E_[p��S�)+�*[&|O�]�t�<��ף���A�I!~ۺ���g(il��>�̝��~>fw[@�۰�w����M�� �|������yfDm������J�����4"��b�+y��Nqᆵy��sӃ�wp�k� 	�Y;|�;���% �ooW@�ou[o`�[�������׹��0��-�AG[(�/ݞIE!� )���v�͡}�94;��=qg̚���p"C �@�[��M�>�����T�vU��*�:�o�{WZ�Z��XI��*N��
�@~�0Sf~��~ڣ�c��h��̵�k_ٝR���u���]&�v����z�ٝL�HO{�"&�6��n��!�ڠ���$:vD�ڭ��F�����q�q��b3�o<�n��c��<:҄�k�qZ�at�ś�3|	�;B�Hm��g��ߝ���}���-q@�?���d�5�٪����B~r�2c5t��<��[ �t��By�s1�J<A0��K�F��,Ď�D��\mxs�Әm=��BR�9��r+��%QהoݷtC��o>�}��cexNb=�a�t�t.A�)w��R�tS��k�W��H�=0}>]ٶ^T�/�[��s�N�W}F89�����|�i&�-�0���wi��v��9Õx�Fev�(8K��Фp�n�Z�H�W5���<��9:�о�a��f��w�W+3���֜��ާy�g�Iڐ�4�u�'��@���U�.Jf��׻���K{��MUC��@<$
:	2��q�6��-���XD��;9������!a���T��J�\�sI�M?"{ٗ���{vh�E1���
���|$h���^�3絳>}@�0��2�L���3��&��<�����v�N�g��!NLyn�p��e����%R4̺u����m����]�3���\��N !l��ಛVns�BI[����CNQ���z햂k6kE�j�	� 6cǶ��!p��������W�/r��|�/~�|T�T�Xe���#�T���Am9݊��/�������ZS:}��gb}\����V4`�mq�3lv������y�r;A�ddΞ�'L��J|�t�PP�LĽ�Ss]�Hw6g�B^�fX"pt߱�pү+����Ǻ�A��yH�A�=5�N��>��
����:��֦�&pB[F�pϝ{�{��\ɗ�>�W6���3�w���A���M蘏X��/.��`�iA"�vClK
�i�t�ۥ�I�;m���Ө]�x�x��x���nͭ�٣��&�ě�e˴�������A�y�|�!O�Dv"G2ӇM����guŲ�ݯ�Pۆ��َ��duQ��4s8�f
<Ь��:�����^hU�̺��1���)"G;>$�du1�d3�b�xK�����<<���Sd�]Λ�����w��$H�DF�n�&���3��`���\�4�M���V�~v�V15ery���fX/RC݄��b	ċ�R1[�5���z`���6��ok F��Z���`F���evdQR�%�ˢȄ�;��D�������u���Lジ�(�Z;�y�W^�A�t��ٱ���ٚ`��駚bhPE�$#o�m���A��k��<��1պ�m'���*3�v��u=�E��H\�]nSKU�C(ӡ7����m�!�c�7��V�(�##45S����zVB}���L�QM���`�I�jMȖ�.��7ĕ�A�s1lև'T�w���X�.z|��n??�+��}�}}vD���#nX���Gk�p���Ր�Ox\F�-��k69f�:T�R�9s��o���ø_d�俬�OA��a��,dz������ ��7�t���ρ���s�E_<����"Z����8.�Av]�3�ؕP9]5&��%�'yӛ�v�X�{Þ����j��|r]-ꍒ�MY����\���G�>v �unmEc��wZK2=����a�6�k�+�'�W�M*�ؖ�W�0�]���7�5Dqޥj��#���G47��1@{ex��b��$DI�槹%���J��~��i��wFϻ Xc��ρ|b��k�3E=�c��d�3@���D�	$�+�m������T(�ƪw����v�A��J�M��p�2��/��B$�y͉`:y��dO���=�2����ρB��/�s٭Ϗ���5;������珖{gv_#~���{�2Yk�^�}@A({�1ח8�Z�>�,�k�IU3���PM��j�y�('��ݟ���.?)���Nb���̄��.�����*���E@��/��E[�F�0��맍e�� ��p�߉�f˕'m�1�E$�ј��bP��/1�Jx΂�k��["�݊�
�}��縤�4_Nl�#Md���yj�\��gB�0��T��t�6V���j�z3�}u���:��Ia���n�%�ճ�md]�y��i��5,ލ���F�@�:�Z]'��EU۹L�i�����N��踜���u�W�<6`��"���t�����d�<U���/���R;�K�NtUs��!�a��yƊ����#��u��/cvy+F�W�)tu,�|�<������:�'Z������I:�s��A8n$F��ΓG���iiܮ�̈�:��8����gyff�ԂDΒ�!�u�
����l�lWr�W�%EYl7�x�Տ��/4p����k�`��d7���{{)� �U˰��SL���n���Iڣ!���K8��S��S��|G�h:� =z�i��xX;K��1��;��[<�syF�|v�0w�O�}yR���«lPA3:m���5D��jɺ�rӍe	������5\��y�NYJ�x�4!,n��|>���)����x�g�$�1�mk5tŽ����Z�E�Iu/h��6��k�IY��×V���:Pڗ/E�����I̝Õ�3n�(��n	���
w�����0a\;O�����m�v#ź7�o�tl��<bP��y�#�;p�#�3㳎�0��K���T]�jOz�����k��������q���t�F९/א��C�B��O�>�::��Z�깫�ԋ5�\��`o9<R��n%�Uҝ�s9,�:  �5R,�N�d�X��+q���)+�d�)	�@��U�6m,�ee�
�7n�5՘�ԣn�ls��Y6��#y��PS�p_�Ob�s2�\���5���s�^&��G8A��
�#Ǆ�:g��t����R��x�x���O�ϗ�G�@�c]��uo�V��:t*D"����ڑ�r[nb*.�Omęk��e笻���+�
�4�sq�t�t�-���e[�i�#;S(��J��ϷY�^��f�{p�<i�L��]@�21��B�9�mO>�\ݙ��g���yl~��������A��K��H��-q}t%$Lم�ʇ�`�t�%�]�5�!��^`��B��kܫ�}�����kǯv���U�S"n�1��[�ƥ�Es2j]����.���
L���f��'V)Υ��/� F�{�/"m%4ei�1odx�O�J�n��� 5�:,h���9��w$ ��t���O���t���E%ݫ�s绶�|xd��w�{U����zXMÒgft��Th�ʯw$�t�HԌ�{��W�N!�V�}#��BFOd��J����{�)�g&��Bo8t�oWT����G�́�؍F�yoi� �]�����f����7���m�_�����Z���y��h\�J�7��}\���@aux��[�}�L��k�D��ܤZ�2:���g@���>]C;��]�Q���i����N̯�ؒ���P/�G��88n�l[�����FS��\�F��xA�~�(����]W�.,�:�2U�)p��Y�Ě�w���w����W���N(#T�z&����E�W���� �P��쒻��#1���mR�;� �
�`��>N��R&M���X[3��ꋛ�~s)E�{���[�PO���,V�������a)"[����R���۩ثP�Z=9�7T�:	cw��L�|dP�O��2�VvL��UMI���҉��,�������]<>���7a�;��jѡ�y�Wx�U����f��:��k:p�3�UG�:%�Z��A��Ky���fAs�C�1]��c(�t����,�w�*\�)���[����y�)D�J�"���E��>�0;��|�$&~u����,^��>�g��7G�p����C�d��`m�5�^:�=+��\���;=�bm�&k�Fښ.��v��n�ýdXD��к:��xv$�v�D�Q���.뚚�l�s�r�:�i��\�3����l?.4#��2s���'�RV[	X��޻)<uw^���!^�Kl!����vOj�����8B��]y|.c���I�}�] �ӆ�?�K��9t�H,렽�7�.�׺�j��n�i���J�:���9CLgs�Æ����[�^�T�Q[��a�6��wG�σj���㻲�p�zk���o]tw�WKA��su�����&^��'-��B���[��Yf�;��Ë��f��	��ӑ�ܺ��<��\-�՜�t�
F���S.s}�Z�Ǉ@�6j���t6U��D�&ws.�R��տO��j���#mq&$u�LG`��6�֌`�}�jG��K]�ZO���:���o�txf[G�{�$7���i���3oT�����<�t�:!1礤F��_�v3	=g��VŠz�������ՙ#�^��~�[�3F<�����rjf;.=Ԙ�Vjӛ�fby��>��p^
�I.���-M�9�jUh��/��#v���Z��};oh1���t<y�PT#�v�ENz��2���
ɷ@M�#�9�����20�lF�!=��7 ��:O%BU^s����~y|n�����WE�p����Q"�b6��t��:\�L��W�XYB��|=?*`�O�w>��t�aC�|�8-�G��n㮝�F�MR���Mض�{���+����ϸ���2m�§�/p[�E����hO��������������{���w������}�����kg�s%�^X��)dߕ��]�ԇ�(1���hu������5v�d1ȖK�l��R>`����mG,�;Z3qV@)��s�0�:�ڽ{��YD�VL��(s49��e�F�g�p�YC���T�k�e<�:�vh�Z�����<���q���Ή����������ze�=�*''��d7[K3ukT��ݜ5�}�d460:�2��+�zbI��5��b���
�a��:r
��1��v��:�+�Dۼoj�x�[�<t�������K�'.'��$���xc���Z�g��U�N�L��z;�J�  �IlJ��W|�Zý�+;�
[���G��R����Qx�0��KJ��_.%{%΃�A�Q��4u�Jc�t8*�h��NF�"5:ݍW*T�թ�ՙi[�K÷6e�#���H�f;�#Ԓ��J�ˁ3E�o)��\��Q�sǸ�ׄ@7&�!���2�S�q��ŧ�[��(uiՔ��d�6��B:�nQH����z��./"��#����7�lB��43��T�#k-8��9���u;̌�j��N���EZ�u�;#-�wIh%ŕp@d������/���s��99� �is���&�_g�tC[S�7K�^'f��4N��I�����]�ڠ�����lnV�:�t���]0�.d����S�ǲ��f����sV�	Pɲ�\���@_�!�z5.L�%~��Oc(P�n��Ô������\����
(��ְ!��_E����&�p`����&6!�ҐGn��:6���&�P ��ۮÄG-E����r�����п�KM�\t����i��d�˯k L{AYW�F�U��	f��tNq�<���Zd�X�5MM9w�Kݗ.4�:P5��x,�j�ݻ�e��Z�%6q^	����6D&�b"f�Lj`�o�9�W��N�L����:�v�WD�v���]��C��^�+���m��u��aBFy��G@���c�1Ŷ�s��DS��\f҂�s�r��:�<���i�-0���7r�ma�"i+L����t�lΰ���k�t0�)х�+"1��IU���Y'Bk��Ą�S�8�p��oz(i�]�o3��sL&r��o*
R���2p>�z��wFkt�ʋ��Eɛ眔�Fh���5��x������moG���vG��:�����>I0D945��Û`���K������>����z�]��Zސ��p���*n^�%y�S��R��b�iH�J\��ܯv���}��2��V2t�16x�a������7�_rx�L�����PBN��c�`\��r�F���Oyi���u9*��o��׫9x����p�TITޚ���2�R7�N��$��;,��b� $^�r��Z��r4Rt&R����ߏ����~��)��M	KE&�B�hJ)�%�\�m�hkIJV�i�� 
!m��ҺJ
CA��4�-V!Д�iJJGQ U�P�4h&����(;d����5E���#�t�P4����4��4�!��KQPST�`6�L�@TD�E��jF��6v�(�JC���b)����RRհj��T%1�h*��Q)�aۜ4��9G3����l%-l��M5MT�[	�	 	�?/�:Y%��|�-�XqF�D��A�P���ψg��E��F�"�'|��6�Dpĸ[��ٝ�$ŭ�jX�����i�:��Y��e��JK�R�!��S����M���18���<�I*(!L�H�6Z2'!j;+���ރ6g9�sô
�����Q:�v�f��+���~Ȃ�u6�V57D*���zX�B�''I�|�ٝGQ���t7���8��g�y�pJ��k�U2�{�zC�Z�ܖ�D��T��y)�7ڕ=z�0Y��V��~[�w8i#.�T��ܝΣ^0�y��o)��1�v�\O3=�jn|��-�·�Q�>S`��׈F�'$,��[dv#ź0o>x����ې�t�tf���t��Y�C]���³��v�����`¼����܇�F��AF�c�R�m�n:]�kB�<�����*��(�p��ɶ�}�8�����ey
�E�)� d��W»\�c���w��F=Y�c�3�r����[?W��u#�>͵7L��/i�@{��GH�k_��7��:+V��N�PE*��'���_dlMQw��w��;n�F�௕�7k�me�Nu�OG���ODs&�c紶�+sO��0c/Y���7��/��y2����ʙQe��gq��^e�R>�#���E�R�ۂ�ݼ�(\o&`R��J�*|���7p�98���m�����}O�7�\0u���8@ժ@{[:�C�����5�ζ"�p.��פ�s�V�E[@2�ީtT�7�G0mH�=]�����j/�=�:�M'������*��IO�7�� �R<4�2��t��e6�/¸� ��Ȏ����s�2I�,O�d�<��8d6c��A��-�燥��p'������� m�ק]44�[(���z텝����ݥ�z��b�i��X����C�1������g�kbErJ(%�>Ս�&�I�m*i��ϳ��8�o������w0;�lΪ�4h�ʮ�+�3^���5q�q=�@��q�,2G�F(v[���^��H�]����x�[�U�ۧ��m:+�Xu�*8ǖH�A�7�����k �Ga��]�X`�r��{[���q���̪�����A�t3�h�q�;:��g�����
�[���U��׵��ڷ<8˱~�[]`�����ć�.�`H��g��y	����Wp��j��n;�Ϻ��~
��0�4����̒�4�)f��CwZr%W��n�l^*m���h��ڊ�;�w@��ձ��s2�Ω�5�:ưS<���� �p����%��=Lq��)kEG]{��^F��L��6Ϟ.������A�w9!(�4�G-�^1n���^a3�j����@"�Mv{�]fVY$u� �]�B��Y%�w�@fD[�3�we���?�+��ߗ����M��ǋq�,��m�a��>I���7ݣ��fr�C�e��wd\w�vz�<��w"��cf-��N��Uh���Cp�}�H�ή4L�yUx�gD�M3�'"�BC�D��4����VcDp��f��%�0����jF庞̑y77��R�λ�$�؞Ʋsp'�Hu�����H�:I[t�q&\�4'���\ъ�ε�n�	D�Gn�`)U�^�\�z���i}�m�b3�E9��g[����Nz4#���=�g�݉U]�4�z=-��ɧ���ȪGߩ��!,� 8��0��f鹖���9�՛=+�gszi����&���ޟ���g����gwZ�YJso��W��Vjr��i������OU�Yn�r�tyf��`��B��u�)�(��u��V�j�}$Ϧ�u&8�l������2Ux͙9�\-F��ƃ��!�l��F�v̫��\�kʷd{,�lͦ�
���]��k�]�����o����~/abt���̴v���n��h�pF���V�ey����ñ��v�ϒ6��k�d����p�6����y��]=�q�X�-3�62B9�6��	�4�ׄ�v
��Z��wtO3p�N��3��9c�
���o�à�h�Ñ"�Rl�^9��,��]gBv=�/�$��/��rl�0���f�𼾜݌�C��ևZ�;�N�^9���΍ ���y4�����k�܂WT;��������uXzw/��e�uSWb�)-���oZ��s;,�
z�˭��-U��Θ��F���L��I�S�xv�ji�մz}��.��+���IQVWy�a'���FN�OF�o���aƪ�����3���!SvB��5�S��M�q�˜�-�����X���G���_T�%�c�]8����5Ӯ钗G�A��'�(�s��
a29-"ub̆_4k��r��@�K��+$��z�Q��a��@*K-ևغCrK���I�P�Tm/J��?�;��E�OS�{�ޒ�K�KÒ0Tu��Ǻ#�.�%Х��3C���mh/N��־��緯����ө�pEC����Q�P:����U���8���X��0�{6��1��s�Gu��m���d�ճ��U󫜸�z��jv��c���^N��e:������`��W�^=[w���^/�\rp�Z=_�r��fң�j����X^|N��b<&�8�d7�k[o]
w��Ii�/�prC�2������Y�䶒&�����"����_a�1�)�zڐ�l� D���'������[͆�o)��HlN�Dk�"3.�X���������8s9��b��+7n�#źl=�sJnl��;�����N
+�6�@C�Y՛8��|��`s�]KC�&�5K���'�W���Ւ��x�?A�G����b-J��&Ч{no���쾔�V9]&���7����{���&n^�u9\�]64����X��zUt���z�Zbn����@+l,(L�J�ۚ�C9?@��m�iRd��v�R̹��#�v�H��O4v
26)�FC:�u?$�7Z-p����l�g9��컭=�=Mo�����F�X��E�����}������l��[����qr�-I�xf{�!�P�Sչ'����H�n�o�7��J��X��k\����e����S�&��
l����NB���\'����gX�n�H����0|f���g(B����R��u�*��I��1gV�*�TfrU���I�<�{������z�N[�S��nظ:|���(�����u��֍ad���ג*�8}r�K��k�HC�jOJ�9� ����34^�w�P�x�Io��m� �]@�2ُ��/�o�]�ul̷8FVW?e��n{Fr�/`�YA��_4Kz�+�f�`���yP��#s,A�w�)K�Wm�c]���D9O�ewD�gb��[�g��܀��7�E�(��W��,�lo�У�o����gg�;q��^;ŧ�GP�V�(��L�˹�9V����B�I���1`�OA>��\'+�Vfd#WK�{ҕi;�8r��u+�-�w� EvevG�����}�q���h<r.PN�Bop������˙�x�27/�	�%�=7�X�>�����߫�ԓ&����tͽո���.(w6}ܐWB�[���ͣ68o0(�Od�T`�j��4]<�T�ݚ]9�5[�ecݒ3d6����7b;�NR]�k����� �_\;�X��qL�'�g�:��j���@�ԩ�O}��wг����gǣ���� ���=,q��1�������.f�3���	�B������1�d?q#BD@���*|�u�`�����86�^�"���b֧Ϙ�L��ˏ^�:��A�U�1U"�\㺺k�����:���s=-ag��P�n�M��ȽI\3��&��6
�6y�2t����7��F �cI늉s�� �,A�~j���в!���k�Ɋv�ճ�R��b�.G] x�6dׄU@�gD�	�tB�.�}����om#��[�L�[Vg_{����b-�8a2�Uh'���,_��s)-ż���d7ة���#D�'��+C��=U�@`��gp�w���C9CI��J��Vk�m�KscR��V�P?�V�^q����V;������z����z��v�� ��ݸ���2�}�QF�^���<j�,#r�H�Ή�2-���mU��Ỹ�o�І�F�o��%mҧ�q�k4V�{��c]�=�;�v4Ztz`���+����*��\o]!-o}��n�ێ��ս����Pa$#��wB��3݉O]���;4�O�F�����w�HP�� �V�l�Tٽ�T:�$i��ǳx�'@Z�Q^U�>7���͏0�o������OT6�U#��9�뀮���T,�{V�=Ԕ����:���4sH6���yx��5\Ӝ�`��.2�n��:�M�'4d��6{6��ȓN1��g����H��d�>#7�D(
�d��ك#mq�	�$H&2g�6��u��".[9=����[� �8'��+U�y��;�@������}�-L��>m\(��mZ�5���B�!��P!�V2�j����v�˟�����ȶB� ��
SP��93]�"��xp{��Ig�mL��/���сm�%v��cy�K����+lW��s�֛�IS��v���v�CS��u�<�v� v5��v�	�;�Ԑ���T����9E��g�#�Y�������kv��ʺ�51ӭu�Οv49<O#4�k�X:)�a�P�A&�����:����y@�|�w����-;�)�*R�k�X.í�΅@溋4��uj1sQ7�7�s��(fb���z���A�=��uꃥ�h�§qK��!��3?��m�ӄH�] 7 �L#D���%T�����!�7,�(�~��i�&��pR"���F��q�)_���Sv��\����=c2��n�_f$�}>k�S��������l�u�q��"e���#.3�zwj�!ʑV�*B����X�����c�����b��>������
M_���Kd0��a���W��F2����ϛ�"qXg�U�����{��^E��:���� ���l#ݭ�uK�NЀ���@����U��b���|�#Q�$�Z�E�R=�'f5c�WK�����h��T���cu�-ˆ���v��h�K�f��n���i���;ܯe}�>�]wh��n�g�����D��sEC��5���|��m��G�_�䤏܂��������N�ꮙM�G�,ISJ�tȷȣ�L���.��g�p�d����8"��ۛ���l7�ҧw��.b��wy��l���D���g5��sHA��˯�{��u��90�Q�}؛��g��Vu��1���=����Gtx`F<���ħ�s�K=�N�kVKo�p�uč����`�#b��!�p�!=3��6��Tr���o#e�W��{��] �Ib�E������jŝF�#'m�L^�l�[��s�jz�yP�ף69!"� �E#m���v�6d�Z��v�H���}��A\X=w*,����Y^E��ܱz�ř�۷f�M�Y.ｽv�B����H�bH��ժ^֍@������e,�b�hv���0�ʃ�'n�S��w�;01��L��"������~?����������~�_�����������`���ǵ�"e�jb�{BȌ䕳�r��]��:�]]�79���d�����hՃ�7�;���4��ڦ����!f�22n�ջ�y�lT�:R�Q�:Y50�I:Ð��m�.,�U�]�lS`{�pZ������>����)9x�7�`tQ�um�-84`
#Z�Gz�`͎'�[ܭ7C �ݏu��=s*�e>W�i�a�%,3fK�PV��_[���9��η��q��$n&l'�k���	��&����F�v�������0s*$���4�#5�u�]����oܩ�Yfmp��wտJ��0��»�!��N���:M�v���U6#VU�خ(���y��G2lsp�A�����Hi�@��fo`";�Ѻ�E�G����S��;�����m[Ƒ���F�w�3�f�zEM��S��u�;Os��V���x����;���\��]���A��9ʝ2���"ˣPg@McۘK����j	��MA%���:R�̌���p��WL�.���ږ��X�κ���'}�������#�.�b4�8G�ռj�u���`J|�E`=a�; �o�̗�n�*�\
8�%��s����fÇ�0�kݷ�7f��'��ݙ8oZ��t��@��0��Ύ��Zv���1><U��^50X���+�S`Y��O*J��<�����wP�\v���>Z�A����D�K�ч�e$��11Ʈ=�Vv}ΟPwWck%5�}�6lYT�d�V8u	xӘ4��m1��;`����x�B�X`� 2tW�5��sPW}�N��)u�YޞM�ko;2IS*J+W륇���9�?�ߚ�SO���Y4���"��Vצ[�˸�\�D�m����*y񩎳��J�<Z�X���웜]*Ym�!՞��������q|��9�'��c��gj��:R�ϳ��RB��*n=�9RɅS���,�j#���vZ2����ODI��w�1��+dXfT�9Y�A���6�!����~@Ch:rލ�����l��8�ӭe51�Np#�׵z�!{�Ip`l���0���Yr���5��ݼ�\���h���Y�d2��w��Ң���X�b�k�f;[;0�2tzN��]f�n��Sպ���.c˕�|s1�W�-�E��=<2�x���7�냥����(f �Ù����
*rͺ��}�}[9�ip��ƸZsl��������jPv�{�<"�-�M��xKW�J�>ڛ8n��o��t4�[E_i�4�T�W\�)��d�@(H
�^n���[.���T=�"�D.�K��pT�ü`�N>���{W���D��v�X�)S�V�w4VK��3�3n�����;"ĕ�*\��,�ŵ[����%ƚ�����wf5�d�kU���&9/7�u�6�	9��/��r��͝�R�]yĞ���r͛�����c� 
��h
���bR���"��&�9�Mr��9k��T�"�-$EPB�I��U$T���LDD5����������nc9�G'�AAIփT�s����l���4�#E4UD5UM1D4��!D�S���"�M1/-W'EDU���V�� �]�Uͨ(���kZ�X�UE5@�MPQUT�1CQ�#�Ĵ�6���(�������\�QMͪ���b�A��"j(��)�b�j9b���"��m��\�6� �$.Z&�b�j��H�����:H�j.F(��$&(�*")��)"J���j����!��	�*�F��?�z���������>�Y�m�V85�|��x�Z�?j*�)OV�̔�ʻ��δ�ن��K-��m֕~<�P��/+h8������pތ�16hs�4O�)�ESuX�S�� �� ��s$;��N鎦㯒$�����_�
C��m�$��l�����f�)�}!��;؁L�3&4qӶ�6�SD��`2�9�Gl��;fX#
��lnQ�n-�c���}��<�j��]]5=C�L���\���]Ϝ"Ax̎g�s]��ڛ���C�5�����6gWA�\ܑܖmS�'�����uw^輻��FX�`�[|�oG���Q����*"5�p�O�DeU����Es���uT�vH�om��6��๻/J�`uVfoEnMl1�i�/p��'�l.-�I���>4:���;P��gV�mlI��B������n!�*��i]Í�1�}��d�h9�ji���K��nQ��U�����޳B��v	���ot�e���H���<�����v|�J����&���J=Y}�������D�T�?l�:�|�Hg]¶�mk엓Xh|��9��F�#O"��C�h������n�/"���˃�x�/L"& w��@�F�G.��p�[�\��W1���P�[E^=E-�{O��u.��)L��\�a�/�۝��V�qng����Q��F�j�. �H��zl�0e���+����|�&�N�u=�����I�`؉�ꌋ�.ʞ�7�ڞ<Nߪo���|��R>�R�#� ����5,�+�Y��0�uI��\GT<�K����G]p��&|]t	Dك�yU��WU�M��vj�a�ɸ���y���QB~S�z�z����ћԑ��$S3���)�A��}�bl��^n#�]Q'y�I�E؄�p��ۮ��HSt�qЋ��۞vڲ��}��lb�9�����u#q�Gd��ܣo�h��\l�3��c���v�z9�Z�|�zCq�����uz@�3�ؕ[Q�᧰y�e��+��=G��9�Sm��0�u/?H`\0���^ٔ�RP2DN���'e�=�'*�UjO�����!����<�}��jK*;�?u}9$8{��U���yL�t,��2�Y~�LY�4��T��|#M�����0�׭��X���:�>�8��5e��3*I�y�+���7c+��]7����!�d�u�V�T;9���];���KRv�c�(���*Ԏ���������	},L��
R�ᱪ��5T�����2�R�B�=�k��R������������6s_7K�pL����{er2���	�sK�wF��8n����6Ԛ�;��O0l>!�B���>_X��o#0f��&H�H8֗]�1�4^h�����O�
�@S�� ΋0&�ãٖՑ1��ׯj�v.+ޭ��W>��>�g����߭'����za��\�ԋ�ozE��'�϶�Dg��i�ԁ�O�g��$+��i؋�̓|'V�3v�y,�(*S~	��i�ԋ�s;-��_�`���}u`�Ӛ� ��d�P;���HW@IPXeT#�v�uv�!�c.��B5�0gH-g�nM�rDX;HnAitt�J;1�kȺ�.};�IǼ:5ۻ������u1�4�ZDc��lDm��),���lґ�e�-¹Y�ɍ��4�l��v�- ���K@�3�a�P�����}���[*�αP5�ĩ��i�E�*x�+���%й�$_��dn�Z�����z�y���J=��;#��2�d�@^�`nEI^r1�XWHi_v�;�=}��p��WlM-/:O���z�����Ek��~�?y�n��r��s>�'����Da�U�U�JY���|}N� ��ak��k�K��;Ta��4ʣ��מ�:��djM�Ś���/�+CH��#}�՟�w+f�^
��U��NgH�#�Qy������0�FN�V\��~��Wa�-�ٝ=����rZ�3<�����D3׮KG��q�m'��0C�1���#[rF�R�	��^]F��"huv�q��u��w�j� -��6��gG3���fFHY#p�����4CZE=M���3���<�g��'�6}�/��6���"�ZT�e6����k��XB9?q��t�W�v3QO��%���w����\�Y��6K���&/)_����s�L���G��N�9<�c�\�ݨ�Z�a?i)k�g8���u���Mǟ��u��x��-j�0v^��]5���c	 ��և�ٱ�����K��������-���L�re��&L�u�!sD1�}��[v������1;��2�\w0:C3<{Yx���EQ�?On=���� �F�Gԩ�q�2�&����SG���qA\��ܨ�^��Q+Ƞ�HP�yH	��=~~K��ʸ����T��հ�KE��t�E�j8����{\bK%	N�3����R[<���E�?m�BUo��u^8xl�I�s�4	T�"���]:�/�O�
:�\<mJ��ƾY��Ź��RVܸ�m�O.�p�f;��Z��dͨ��W\�6�l��y�= GۏA����T׉����c�9׷�m��*fO:���8��\�t7�Ѳ��jz�ئz��rJ:�3�/oԭ����s�§Z;��3t0<ˎ�j�F����n8�7����ˇ��ٓ�M�)7b�m0|�3`��pQ���W�&�Y�V0���N��X<�'I��k6���A9奌�l�Z�ԥ�i��S��졪�����#o2��9�B�i.�
}t�7\.�G��tޑ�qZ[�gUZ�?-횽��ݧ�����ش` �ڣ���n�⳥W^���l�f3����
mY��uP���#'h6�|�m;S����5��+���K˲=	���8�P/>�WŏI��zC�b�)�lFO_n^Z��w�5���\�����gLp���d�hE<�{1�8�˲k{���a7���]�#�>�	�tU�7Ne����BK�b{��5�a8tE�a͘}��dVZ���ȉ��G���h�j.�.�#oQ��;�d��cld�Y�7:�x@����gK8�h%Ca���+����"���S��[s���&�'����T�	i�늉s>�Ν�.=Y��u�s�--��§����2��Q����+�u ٓPyU̐M[�[FL�����h^r��j0Vy3�D�/q�i�iH�xJ�*\���#�tT	��c�N�=*Opk�w�(�3P�!�B���G����(�$H�5���#x�I\�+Ɗ1ͼ�tō�xE���q���7�f>A�㔜6A�W���TDp�;ww�����_!F��wX�+��)y�:�Y�.2BB�r��� ����j/x��Z�%��]v�ގҮY�;V(1��p��4�԰'�uZ��|��!>'�l�3�yy��Z��� �W���#clʡ�����*c2lmկy��]��������K샳��0���v]fxd��#}�CI�{��J��5�.׻��y}?|�Cp�#Qc[���e���a�q�n�7M���n�NEr�9T;�*�ܢ�nɽ���-��y�kY�叓�Tu�5���_ �c�n��2̌���U$����'�QUǤm���ͩ�1��Q��ՃA��!3�9�0ط�r��H��~��1�ϳ����]��dX�9����U�41�02� %v/G��&H�ʺ��M2��0��m�_����FF�p ��g�Ƌ0�To�9h�������H���ws�r#O	�r �|:*����d2г��"�\Ӎ�&����]3:4weT���^#��5��O&�o�]���P�?+��k�b��}!f�:`́}�:�qћDS�܎��C⡘�w,�}�eΰ�7ƙ�Ω�Y��L��g�:��,���uG"ʵ�0R���]��SD��z�(�\�e'-�Q�h���/"Ǯ��(�]Ɇ�È�c�v�ꇠ�%;x�癨gg-#7�c��j1��9�w�l �en)R]�6ڑsNR�޺xyjoF].���c�%�����[�ɪ2#ݤ+��%�z�5=*3�Z	h�\`6/��O0�����^�g�Y7!�5aظrK�ʡ���x��	�ͻc'��ur�-�m�����<� �2}	G[|R��֖�Mvf#��j����;&I�����N�����S����*����A�#�7<�뭜����J�T���R?����b��)ǐC��O*��Q}�����Fq��+6o�Χ�Y\�j�L�Rn�����큵�T�i��Gq���\�m�	��Ȟ��j�^iay�ɵМ������v���5����z�*�p��lΪ�SwQ�K�&��sm�.��^��m�}�MH�����s�8׶<5���vE֯G�������X�l�2�re��h��fU�9�,�{P;A��Ժ��x�Z��-eH��~�dL�Z���귮";��.CE�a��P$1Uӆ��4�`0,fuwg)�Z�� ��ٴ�.�.���1|:Z�e��
E��l�<d�]y�Ϸa��(��qnH+l��_���� t���g9��:�b��Y��I˝˫~��3�O��oP?L���;�{Evu}vq��0#Ti&�u��k�c��g�;�G{��9�$q�9ӭׂ��b��錡]���R��
l�f�>��������=��wD<��2�	����V$��ț�a�H���r+a� :YŅ�p�D�OOP܌\��+�3�i5�e�]6�Y�����9��t�e�PW�0�d)�hE�N�gBd�I�fnc:j�m$���Zf\K��T����Z�So^���[S��������獋,H�r��U�FS���X���[8�SU�cz�Z%���L��0�y���Z��A�e�C�	�J��R�[R�9�b���j������!�D�@�[.���wIHs�q!�L�J�`�=��st��q�2�=*�{�}���+2>�5�`�ϳT�������LEA��a�x5� ^쾝z;k]r�V0�|�%�C'��"�:}7���0���E��etP�}�[J�88V�(�w�X�͇���3��oc�#	��F�����ut�d�����9�������6�)i��d�&W"�q��5��-Mk��jӣ�sA7*F���An����:jz�=kbHy}�-.��۵l����V�彫��k�3a��u�b5t-�n]��#b�Bi�gq���x�8�7�f���F^��!�lʱ^��������>��p:���������=�~�I�푲:�t��DS@h��u�Z{Fl,��^R�ǎ�Wݤ�ʯqc�	��_�f��b8^o[�s�[t�оq�gfz���i��]B���q�8_D��=�K�~�J����0۵S/Y�g���Kq������r�lU�ctǳ,��w��i��ȇ;��Xwq�f��5e��}��/)�c�v�	���˯p��:������:��f`D �&ȟvi�3���5>�P}s�kK�ͧ_-=U\%$rU eڀ�"�S���d��QD?�"� ?у#��=O���9	FeY�fU�`Y�f� �VB�VeY�f�FdY�	�f��fE�`Y�f�e�	�d$Y�fE�VeY�fE�FdY�d Y�	�fE�`Y�f�Ve	VdY�f�`Y�f�VeY	e�	�fQ� �`Y�f $$Y�f� �`Y�f&E�e�fU�dY�fQ� � �V`Y�f�VeY�f�V`Y�a���d ���2��ȳ�2�ȳ(̋0,� ǈE.`T�¡*pe d@`a@dPeDu�Xr��0 �2��0 �0"0"0�2 2hU\0��>!⪰ʪ�( C  C
 C*����0�2���p 0��Ȁª�  C*���2��ʪ� s!� 0 2��� ʪ�  L�*̋2�:0,ȳ̫2�ȳ (̫�<�"�0,��*� L0,��ç̋2�ʳ̋2��3̀����pc���� ��B*�@u���xl��pd_����ֽ�><CT�O�,L��g3��I���p�s�GB( ��r_����+��$(�*�������@�NI�ޟ���� U��Gי��M!e�-֖/�x	} ��C@�$Dz̙"�� �"�!@"! ��!H��I  D��������2 �
�*��!  B��  �*�(H ʪ�  I(��$� #����'�������"���@�P
Р߼?@���o�~���2
�з�j� � �H8iR����'M�S�<�ISh� ��9��T�?�9���@@_�C�H~�?o� UPW���<�� ��N]) ��j3m0�H=a-uJ=| ��PV�c���C�����
�
���Ĕ���٠to7�-xsH�v�J��ه��� ��j8\�B!7�3I����A�7��K��|�{��"����A���I�?�<��������O�_�ET��� ���*������ն���I	�����)��O,����l�8(���1 M�>�T�H�!DD�J���H� �J���*$�TE
*�����U E �!)JT�)IED�T�(�IU(�	S�$�Sm$�DE*��P��" �B��B�PHQ��T��ER�EB��$�!�Q-�R��AEQ% �)T�@��@�E
IR��IU*�EIJ�J���
� % J*���F��<    �}��5�u������5����h��]�%r����mIRq+�&b�+�6��5v�Q�N�.����Bښ�Ӧ�l�6[m��J����D &�   n3����h����
����7�vƴ�k��#�V{9����lkM��l(P�{����֚v�vU�ֶ�Wq�4�R壒î�Cv�2b��;�݃�[�݊��;�ΩQJ	TT���%TU�  ;�6���J�Z݋m5F��f���mB�T�:��m��ͪuM m��t]�m+H��4ֆ�MR�U4��s6�J���-�ZRkZ��JR]5@�;j��W�  s{4�S���[	T�mܧ)����:TᴢA��]�SZ��J)c�9u��Ψ��@�Xhj�b�l u�!��ԩJ%%T�D �7� 3�U�=`w.u֪���� �U�;�u\M��)U.C����K����q��ݪtL��]ڀ��4 9�)J�B�� �*Ro q�U��X
*��j��e�&ֵ]��gUԨJ튇L�:n��AuTdږֵ�أ�Sb�pQ*����������x pUt�6�zkAÌ((����ViLt(�Gqʎ�iV9�i҄��  F�C���P��UB	>�U""�	� �| �+z���݇: r8����  k��� 3� :T�;� ��9��ӝV ��݅��XJ"��!)T�D� ;�  �FM ��
 
;�j  �:H(92�u�;�[�k�  Te�� tpk��7S�� ��JRh)(JU�  ����[��۶���(  @4
�0�Pp  љX� �:4d�  3H� ���&2�T� ��F�Oh�JJT ���z��i�@ �JT�@� �@eIU4��4i���)fUJ  &�S��=����Y�'&����q��S�V�M�s�}V���g�WA�������ܻE���mZ�~�m������m�[o���j�����j��[mm���?����������V��i�v����CNH�n��6��i����g�V鈍����/9[�U�D��V� �l��֜�e�d��=�V#$�a@S���l�XAN��68NiZH�#����DU��aЙJ�pڭ3�0^9ojR�ژ/)��,u��5�x�s�+	4!�J����]kF"� U4�R3~5�Z>u��2�!�Y��$"�GvⴤzՍ;m�'w�VIj�먭$�{�e��Ģ�[�!6�i������՚��v���e[��1$(�T~�f�e�;�mG[1���b���،��Uu%�����RN3B��gv�&.i�A��6㷃&��X6
��8m�;jcN����t�s`�>��ĥ8�v�Z-:��Ց5E��J��@'!�[u�z��N\���
��#0�k�dP����,ʽƵRj:eT�V7::d�6n�z�P��]u������V�yj�кJ�nk��#�������Ʊ)�9�v��6�k�M"����V�
pV���f2��N��Ćʫ�0@�ȱ��E֍F�ΛU���(oسq�-��}��Ѹ�xU
����x�T\zNYݬ[2�udi. �F=f���u�U���Â�RP㧖�cc&%&d�^X�$�,�
��S�:��]7!Ta	�j�-���`��y��ݹs��T�n)�e���X���(+�J�T��Z����:S�֌��2�I圶�n��&��7���Ț2��0�u�6h�%�ܡj�X�۟h`%eTCD��
y ʍ'� �@;���kx amJ�SR��3!řn�]ը�SZ�Sp
jm�Փ	I�LL����F��y�c�)Gx��B?m(�K��-C��nѴE�Ok5�RR�Ha�;ge駶�m�*ST�[n��XaXʒ�*���'ISs7h��e\�`!��U��Uum˔��e����e���f��mcv*����ad�lM����m8	�{�b�Z���u�3�a ���+Jj����6DB�֣K�+� `V�4��*.����r,�r5�pX��qҔ
-�w�GlёZչbX�˷1T�6�7�q�x��ik�\�#x�Rݼ�/X�Og��Х4�q��Lͤ���i]6����iք,`�V��c�a�{%��%�q�j��1�ة&�m�w��M"���;V�=���`�c�N�4ꍹobu��l<��=�h���eD@6���7��Rڻ�C�v�-�ܥ�2��E�ȷr�ͫ��yN�Q�`ۡ.�� �RJb�����.�B`�v~��L��=�{�K���4"�ڲ��q����λ���6)���5	�j�ǓX�Z,�#P���[{Y�%fᘨ�j�Vʑ\� F�*�^�Z?\!Sx4\���Uw�淲�Z��5[Yp�Wj)Z!VVPu�vu+ɸVJ3	X�YKR;H��Lmf-.�mn�����)⹵d�"O�;T^��
���fyJVC�J7R6��PY�:p�-]��Uw�"�
��U�X��쿯&��p�:G�,G"�`����x#oJ�b��؍��J)�Y�jD�]�+P;�bB�]�	�+F�,�O+���.�Gkqh:�\�e��b�@4G���ҩ���4�VM]�oѭ�$X'i�� ��#�t��ık	|wԨ�crc�h]�J[D�";�z#�$�[h��%�WtA ����wM��*�X�f�$�6@O�nl�@M��n�%�nݏ��Qӫ��6���w�fb7s7*�S�4t�Z.���E		�֛͜K �vK�)�:-0Kfa�L�dH�Aw�ͺz����ݱ*[E�M+��[,�V���{��@�n5D�7D��c�@^CY��A��Itj`
��]�"�ݣ�[rQ�X�b��{N�+�N�!t--t񇴚�湊�|�!��e�4ha���ɴ�_ ��[��p�B�1�����.�`�j���l|$YHM�@0nZ�)B���'��En ���;��&<+*�*9����ha��+���֣��@ì�Bh�]�#U�۸��Rk�l$v�+�g"�e�{W���n\["�-V�R9B%E�1�Ug/-R��yug⊼�iB��n�ٕkV�uP�H�ӹ7NM�G&��b�Vfʏn(*!.RL\�N�7G�.S��e)i�� �i�"�Q�`��f��S�写�T	X��C�v��u�X�Û�ޤH�y��4t�)�3w7��`�7]�#�.8�!��$�X�i�rP8oF���F豮<ۭ�A�p�{�V����Ү#z�p�͗��)���ą]J��$���x�i�;R�3+ᆂ�7���I� ��5� 9V��������)�WT�(Tee��j�h[X�:�ҷ@�9h�2�mF�
hD3,��+���4���5cqX���b3ne1��J������/S*MʐV��i�tibvF�Y�LR��wJD}�򖺙Ad�Ɠ{�kbc�T����C��
*��A�,��X66���aݼ�m�6e��Q&-�DWd�@��Tؽ��BfV��+�E�h��X�G0�+�o��I��4��1k¶�Kۢ��0j�tO� �6#HJ6iبU�`K��n���(����Z7C��ٶڃk7Z�2bu���R�@"��r	&RS�R����CM�{LBU�k"�v�⛿M0fS�1��x�P���h�z^i��;t�$1+Ӯ^AA �^�yt�3�f	W*��N�8�#f��-W-^5�bl�md���٤�cQʷ���N�Edn3z�<xf�����5@�ucD٬�(+a��H&/LVU���R))�=�W�#+����$����دǉ�[�0P���3so(d�2VK�f���#�
�SV�;��-*�򌛈<Ahr�q����[Tuf�ӆQ������Ɓ�6��V4A����L��Z�s!b)�6ުN��m^:�į!1�Z�Sp� e��m㫙����/0K���H vc[B,)�*��k!�Io/�( ��ǌZ
�05֑��	SLGk� [.�Ew�� �Ѧ��do*x/d��#.<���D`�),mC��d�:n�}�UgJm�r�x̓l�N��bˣ"�us/hP�;��Q8�i�n�A��vM6�#oS�˪֛��E���*B����-� �� ��{�J�ʋI��ڭCk&��{
�[,�.�%���F��k&�Uf�oB^a��fM8���M��.����q2.c����w��Q4�!�L<�!���٬��H�&4��:v-�i�Y�A�%�8�:���̭b'���q
4�[����bD���B�%K���������&���Vb�
�A0R�z��wR\Q1̔m ,?�&ݪCf�;��ۺp�I�;j];�v��1����HxT�X��mީX���T\֩����VV�-���/^���,���R)$����L���NRd8� ie��1"ݕ��F�3/�j9�W6T�R��tU�8�Š3f�KF�Kj��c�ʫ�� ���DEK�twz��F��I�CZ�u��Q��tP&����U�3���J��
0��S�W2,�3j�P��mԎ��.Z�ij�Ҧ�A)��s]T�Gm:�od�,���
ՁPq��tUR#�⼘"�Kϣ�$[��f����[��'�+5nRε�QQZ�Ф�%���o#'
�B,%@�g1)��� �EOhTX��k��H[�Qe`�ƭ�.a;spD$$X3�Hd�kk3P���c�w ��
Kx�L�[�E�vh�M-��-���☫
$��ur��4dv���ٯU�n�J���0�
��wue�������֮���e�@R�*^[b�wu�Q�nɩ1�Ӊ��ۢ`*V�E�q����`�ʞݗ�r�lR�i'�)!m�v6kp53V�3!�%>�jY�ubU�ٲ؁C��B)��ڨ�kr��`9�VYN�,�՘0����F�i��u�t1��  �6M���]d9*Z@��\o\:���Fobh��f����û�`ÑK^SZ�N�Wk[��w�r�'�m�T4�C�bJf�E��@w�Pe�ʼ5a][c K�� 歂�T�ft&C��`oR{�N櫂��8oa���X���W��\ܻ����ST]J :A
:�ǻq�ʊPtrP#>�Y��(6|v�����A˕��^��CV���~�ࡍl�*	�J�S.��4f�ֹ6Ի���Ԭ[�փf�S'D��i
�U��������(ѥ�^ư;J�R�4�3�+%��0�2Ssk.�f�a�wD5�$�l,'#�XE��nPB]%2:�ۋser� 	��	�!ҳ����Sm��i�Z!��ï~*2����!�ż��h��SH,nf
�0]hR�`ݲ�[�*T/]e�㻼�kB��<�^7a9b�� W1�f� �v�ݡAf+��YN�(-�hn|���cO®�B���k;�(�̽�F��2"�b�&G3�n����]m�g���T)�r��zq:R�L�����9�6��*�z�����3���:�X�{��Pv���AelhV�������L�`��u�	P|iU�J[Mct��3��%��eo�U�q�/-$ؠA����4������5hjcدJy&��-a�[�zr��LP˵.���gso	D�Dj��ZC��+�g"(n�EQy�*ש�׭�m�f9�X�Q�kQJ`��C���3b�ͨ��A���0_ٔicF�Cl�Ϟ�9I13.���u�N���a2wD-3P��{)Z�%����Ei]����6æ{MZ.l����mT���୤ihSq��m�B��G#����tj*��]�8��OsἍ5L������P�Tږ�m�iKSIT�60����[��l����	���.����[m��Db�"��Т�1aҭF'�5�����e�w�7C��˭�������2��-f���Q%`����)��+MҖ�-���fad����%�g@Á���7����t���0-�d��fm]d�/-��VD�#jif��1R��$B̒�.��8�w{WPh �j��sQ'l
�k�L�6lytM�+����vv�m��n, YM��/R5�X6�9cq�ն��� ۊno�:6hM�՛Y�ڇ,9r�T��{O键Z���h���XW��W+f��ct�ax	�U�O72JQᤕ�d-3�ǋcwt����`��&��9�n��:�u�n�#�S�P;F�mb`���(�	�8��EF����,���Yb�[-���{����)��H�V���L��h�����z0�tZ��t�V�sI)�u�rWSm��7"���b�niЅ�W�A0��k^�Υl����ok!��T��jM�`�e�%Rur�Ӕ
%ض�X�2��32�r�(vq��V)�'Fn�J�`��w�m�rI�5b��˺�"�n�D�1XF9�U�y�=��H�ɥ��J`o6��ٰ 6Xqd�q(d�*ްE����;�ז�j��l�Vee��6�S$��(��qg+&E,�Ҙ�&\����S�k>��X�6�+���L�
��ɨ����q&r��f��<Fq��qa��2�gZC%�:���v6�%��,V8�+S@�*;VZ�!�7��B�\T��B�	 �*�^�m��Eai8�t��@P���>��dE����S�u+wB[RP�Y�(��*
U�Cw�VoC�˵ �F�#Ђ�Z���L`�
�&�MX�Y����V�f��_�2BW���iC����*0�F�,\9`��{���D�w$�B�*����Y�@�N^i��ا�w�η��8�����l!�,��Q%Qa�6�ub�N���Z��&�z�^�)f��LT�'�%�L>��&ix&��T���X `3�ӳ#Klɺ�ݰA{p�!�f�B�8ٹ����=�u
`�L��!�3NZ�~3H��A����f��ˈŝ
��&�3]�E{��5yD"Ru՛��u��4;-
:�L��6���@Xwq�Q;��a�Zщ�W�t|�2�6v�l���ǆ��4(ʛV۴�NC��m��u�q�j6 ��n�B4Q4��B�����+PV*9l*�Ȧ�qV��nk��fl×A����#+U2��p��\���I�ܺj�� !f]���5����ө��c�wR�ʸn�%�}���yor�ǈ����6�1f3J����z[̥/pJ�Ĳ�BT��x��L��5W�kidyI]�Hn��ZЄ��2����K��.=�����w��S����EC�$��[�Z[9�$��p�=��qeƫnн�$�t5,r�A2��F�Ր��#����I["��XF�{�1�K�&lY�0��-
l⨢����,ڻƒ�Za�U9@�p�a�L�tJ�SS�򀫃$��LP�D�!S+Sزf�'t��R{�0f^U��}6d�ʣaV�[II{N^���j֐�0�j�ia`�-�V^��d*@���[�A��Z� zQ����Br�!��B���ʃ�ظ�{V&�����u�M�}�Z��\�	�m^9�j1�q]^�R�*Vk�6ؗA��+k1��]��N�yZv��.t�)�a�
�6�Ӵɉ̤Mc �%f�9[�ޣ�Z�w���X&`GK�zը����ăl�˼9��>��
�����m��)(�|1�ҘA�[�V��9x��n\��:�h�&d޹rˁ\x���3ǳ0а���b�2JyAm:��8���u ��fx�Wu��`����v�ǻ֜[ϸtZy�L��&iܗ�{:�Dܕ��6m�h�7���[����J���'{�3�Xx��v�W��9����;��.�Q{K���'���Շ��wa��@m��e��^n�^�%æS�#���ڔ��>��H��E�H7�e4�����_'�^Q�k\�\f�w&m�ms۔������鸚���#}�W,y�a��W6��,�r��X�]˶�#�U�-��ì#X�<8��Ȭӻj�yX�,膜:jF�^Jy�O��1S�J�F��i��ӏqe�A`r��!��K���\�و�u�:m��:bV��Xn�P�[V�ef\9��ˎ��=�{jfY��Q��4��;����$M5�N@-�C�8���<U��ԇw:a�j+�b@N��0sR���ZX1�g.ө`nՑ�����a�<],�m���wqG��@���v:��P'��>�r�M$�Z4����ٰ���{�/��&
w*}qjT��kN�o�tC��[FÐ+���,!�z,�[��2�����Z塧AE�%hu��}�/����\�;ked]-3��L�@>u#ݓVI;YZ�,�Z��c�LMmLI ���:/�����t5+-]�7�w5�KJI��+�6ep�}5]cl]�0n-�gw;�U�5Ӄ�-�;)%������R�]2�����i6��#��\'"�	8r���<�آS,gt���5�Y�S9��7t��N��UށYԇb�(�!��� ��qK=H��{�b��W�H5�iQ^�(��;�Z�,���^&�t*�6���/��N�u�y]�iq��uIwYO��5�p�t���E
������vj�c_T�T���N�����]w�L�y�TL��@}������ij��^߫\]���W��0�.Q��Uv��%�Nm㛨40:�7�k�{�a����]k� �W\F��mW^�Yq	�u:Ԯzd�ӆ1�̐H�s#t���}û�n`$�G�R����N��w4��1:��#��g���K����U	�� )ۂ¹����t[�'7vr:%��cTJ�Gk ��ھ�0�;�	�܌,e�M����a���F�4u���X�z����4�X�ڈ��+]��"$��,�:�Nr[+�*�jH���Ʋ�a`�ˌ޻"F"�����m����.ʷ��o���;��x_�����e���v�]Q�T�k�������֧�{�	�	/U�kX%R�p:n�c�%��:��F�qt��<�9}B����V����Pèo�1������]$�D�ν�p�g���înKan0��y��T�7M3!s�<jk3�r�t�o�ܬ��7*���3�V	�N6���3������w�Wk.�^��(�o�7���������R-�����;����������"Q�%)�m#[9l��P�R[ת�q���gEW�nM��k#T�X�fPc�w���Squر>ʒP�V±Wbu���m��Tf����3{�=xq�upG�\%��W���߽�6����ҋ�:��dٿ��r��]�S[�2��h��4���BHw���^�/��Ֆ�e���}�E}��O�VE��=�}
�]K�]֑I@u!�`�y,��ȸVӚM�c6h�j������}(P]n�v�X��u-�5�|�:��*>�`D���0ȩ\
�p\\p��˜�hخ8�}W���ΎK���:vᮼ��)�	d���;|K���_S�^"?-7�u�~��[7Nt�֏`��9��U��"�Dok�tM�*��x�F�]�J��=�ݤy5���r� �T������*.���y����7�����+�N.��b�����b.�6౜�e�s��:����G���6��gPwh�(�˨�=�ϯ.D1c�WQ�芦��a�7��`6~��	c�b�I���bؚ*�k�Z�Ddh�,��8 ��*�����ܰ*���'\^�WWx[�1�^=G��C��:r��ط{�q��Pi)�Q�����t Ұ����i�� ~J/:�Zz�Y%G��7UkK��y�,�:Wr�XK�l�m���ce��m�oZ�g��y|�VD�d�ڧP��fR��\dCݜ��SϧlQ$by�G�G���ܩ]��CS�_-J�e�Ա۽�`娋ܮ��;��2��r��ת=��A���+���Է�J�<޷bI�>w3�]ū�.z����z��6밽pg+��Z��|92�<5�����o���E7�%�n
��G;Q�j}���YͫV7� �g;-�ړ��k�{����j�ƅ�>��D؅�&o�ξ��F���"���.޷W�����ܮڴU�s�Gl�Y�0���=�u�-�+4��x���w�q�Wg�Es�
��v2���q6�����o�EP�Uۖ8���[��2���PA�㷄����6��؆]�`��i-��Ț�4�_���.T���eX��.��C�1$���9SL��w(nq��v�� ��R��C����p���a��:,�m��{�&��t��4���}����iGO[Qm��W oPv�d�kl��e �'<�)��E$���:r�>�*\������@�t�v�4�u����|	ATy�̗#���
���jb�:���Jhx���hWvj�9�b��:݋��9_pgH9�"��n���nK�w�A^T��jB�ҋV^]�洭�}T)E��2�c,˕g�����;|m����,C�$�J�5}��|�r�o�[pћHѫwN�������:��Y �t�J��Y�bH>ϯ)�����ĎV^b����u
���9��G�W	u��wϞ��tTKohW%�e�M0�vo2w��G��\��Lέ�a�ĵ��ش�\���q�7�(���D�ȕwq��D�C���� ���F�gh����жjƕ���G ���k�"�����I;�,���9�\#�m]�ܜp���+��z�L<}�u墽�[��PÞ�T=VwX̾�S@�cCm^�mYNv�yM�������f4�!����e[��)>G��6������n�>�F��k���x^���y3�:pȡ����cs�PN��_�VcMtgJ!�h��Y�`�X&[��&���S�z���<:�7�/�I��47fT��z�gg�A�l��Ha2eiP�����.s/�LVuj%�YW�-c�N�kxU��Z���
�v�a�-:]P�hW���������;��f�lgmӏE5P� f5l��2���ƭb��4N�ݛ��rʥ�U}Ĉ�m��<����j��5����:)�{]�����XQb"(:[R�9�Oޕ#�Ҵ�˼�+�-�P��kr��/P��W%./�jT1mtTV����R��49<	���:7HS�����b��\�#{U�wM^����/��3�u�}$Y�%)�2V�}+�au�m�\gS'�t��L��|��B�ٺ�$Y�G�d�peH_n�+XH���m���4�����Y��B�)[8�+�������qs'��XCu>a򹖡^@��8J��yEfݘ�j'9�L;�3d�ܡ�-f�Ku�*5��K��ƣ1Uڌ���<�]��ء\��tۭ�Mt�Y1|�蜐����S~G���G�u�%��]�
'��L
�l8;��e�{q`J]Jĭ��7W\4y���+�E�t�jHd{x���Lr��*���x�=�Y<�)f^>y����u��;A��k8�;����Z�aN ����C�����V]i��@�RP��D�_;=,�nVh�T�5�b�㓪��yu�E5�_,[�I�GvEpΊ��<��S��ڻ�ݐ�������|ORY��[*�J�8�U�q*�y�����ښ�KN8��b��}���-{|l&�FB�&E��|x�T�{}v3^�!۳>�]�ֻU��F��[ዯ�Յ>,:@
��aWx��m���ݡv(�U&Z0�L[��K��r���V������Z5���;�.:��K�E"p���K}��y��ڤ$���ZJ;&*�:�e.�Xvr0'B�m	ZeC\1i�����ڹ�k���a�2wR��;W��X:���o�^���pxPG�<f�/k"Ƀ���V�^�n���n`�T�V�סKܹ��&��+�����)Z=�5���e��z�&К����i��b��
����F�[k��M6��+9t��h��o�Η����Xy��gZ�n�Y$jfK�\A� �^���v
o5��r9ېe���tܨ��{��K��\:&���l.L��q�b�hj�So�n�fH�b+��m|����&
�f3�Ȏ���V]�e�S�7���xN9:�o$��w���jI��ͫ��_k�,dm��-W�w�z��>�)<hcasE&ZSS�ݔ)p���Lm����'�.Y:/�.d���]�L�n'�w��E��h�ԇ��+kh� �\rD�ulթy���Ҏi��aY�Z Z{za�n�P�����Q��$����J�5��_ܳ�CP)��:9�����k޻yۇ̒��`QVر.�Ҽ1bf��9F�{�O!Cs���=���x4����T�bڒ�k�3���r��ǿ{��:�uI�FԶ��[xP��!�}̧����P��w֋7��:����y�])Y�fD�c�p����/39h�5�-m=	�C�4!7%��7��BV5�ha�]���*�,�H�� P�E������^�Si֋�mG��u�[���2����B9uom
k�������(�Y��ۆk�XK���o��F^��;������0�#����H���pͥ-�� �����jn>v�-�q���.K%M7�)���)JWFg3��һL��i���"*"5.�{t$����-AF:Z����r�Z�;�B�I�8�m����}g	)�喙̧t��&d6�:��Z,�%�.�%ȕ��;3�T�^�RȾ�f�&��m�����:�\+�ܹ�n>��E��:�2���,=�j��4�$��b;WY҄�� X.�÷��!8�3�]��86-(�ݩL����q�"�V�������r��Xa�
i��v�k��a\;�r�t��P��G��>z�)�U�ִe*;���z��GYD�k^!��!�ȿ�h�@��|�Xa�8�\�
��	cM�����ל�KibK��Ӵ��%n\[�l��qԹH��[��e]��&���v�YC��y����bO-�d}���9��C,�-��9�>�'
����7�n#�����fհU5Z�2��4yWV��#j�j�Gwfhb�c�`�o�����8�#<hgmq�z�^���;ڶM-
��A���5,A2.�x\z���;;�ݮ�e�>ݻ�ŧ�P��eb��7]z,�|�����m,�aos�7z��M7;/x����H��-�����Ԕ�.H��A4���n$�����t�P�D�щ�=��!�3��v��fN͜�k��9ݷw����7m��g���|��ݶ7`�ڀac, �=��`���}2�������f.���8�j|�T|è�,�z5)T,:���K�J3��J�Z�C�ԋ����#h`�N��*L[��6b��sor�:�4���f�wuu2B�n�{�Cwqc�Z��L!W\3e8�&��Ǟ�*Nj΋V�pr� ���}е.2r�(��õ+u[�����)����2���]}"U�R�2 7@�Ե�0:�X��}��r�5����A#�}1��!�՜����Of�J������r�
���(u��ێ_Z���O~t%a	��D�4�얥�n�Ar����.zjﻍ�q���+.���gW58�gT2����w1)U�|�Ju�Y�$�����w��Dvv.�p�����k "*$Y�%�ۧ-F�"��n3n�Gf��T۸���Ro{}I�֑9�*�3��ܶ�.E"���f����90�s>��9�%N���������p1�ۈ���0%�o(�	m)V*v�k�[��s2���ci��h�;3!�yz�z�E"	V��Յ�j�ZiL���ǝr��0���\�WE׬�a��v�5���Q�3s����O�>vVQ�Ge�ʵ��913f*w�k�e��^�)1w!}�Ҧ�ů��U0S��˺�A�46hzj��3I�!�����j�¦��fan�����v뚳���X9U�}2���n���u
�L��N�)'b=���1nc#)<z�IWg�+�0%V�e��j��5��"u������U�� �y�':���la�k��`���8�{�`fg�uh�/��	9ҸDt�.4A47���&kh�(��{s��zn�bA��㫫n�Š�������oN���*E�ت��C6w�k��y9��5m��U�so����LEkꃅ\��R�/\���%x_3- ����I�,f�P�D��53^TA���s^��,���{�lY��`�T�鐹E�N��neoG�;�"]��p��s_n���A�`̨:��!a�[-M,b�n$ܻ,�8��\8җ��5�@����rI>��Ӱs۾�ܨx�v7�;����Ld͠d�T���Pub��
J��3&b$�EmvIs�3�.���+��H�\�)�OmoGYef��C(�0U �Ӵ������{o[�W��-�g�֬�N+rj��m���/(�7������h�>I�wu�ѥ�dB�Nh�6�'���w8�.���7d㔜�j�5��o��z���G{=�YO;{�wڝ�r��v�)�EY��og�']L;�;x�w2����Q�c��b���@���篸���wm�%wuin>�0�Cy���o��g��f���ӷ����s�C�6����YNo3R����x{���=����x{��
�+�(�-���:V9��**�EZ��H���7��������nv�vz��h�b�Z-�F�
mA6K{z��.�FQ�k]&�L^c�&�Q��5+�ơz�����4�L	Ǭr;���
�>�!���f]���� �j�@r�8�j�J�,�յInl2�0����l��lU�)<�c;�.+7�a��j�5��W,���+j0����_gT԰C�&���a`s����]Gk�����t����!ֳP$�FZ
��ĸR[�9Y�m����Z��ږ�+Uo�Ci�+m�
�^�U��;�N�˲u���J�\*.���(Q��uy�wX:,od\V%�bY�x����NG��"D���N�=��7u�:�W+OguKlҨu�K�<F�v�}�'���J��T�@�tM��3,V�m���z�u��!���M��n�ʅ��S��t�}�Ҷ�>�o\Ⱬ�˜)v7"t;�wVҭ�4��{\u�IV�Ͳ�ﵫ�W�P���J�Y+kJ�y�O�s�M��EbPB�T~��|�CS�������T�)�))�q�}�M��7w�Y�6�Zh�BOjQ>C!҄+\9�-��u���b��W]���8-����w�F�#e�ۜ�:��3�r&��+�\F;���4^v,����9œx
����Y&�qȻ�iG�o)efMN�ƶm��tzz���75���t�����]1��hed6�ܧF��ݥ*A��.��A-"t�,��59dH=�C�Հ�4$�Un��\�e�N��޿��kK��2��h[�i(��Mw��ًA�I�|�Un�Ǌ껷�M�tӣi���f�;�]��,E�͊��S��V1��ʊ՚6{�}�G���[�_8���3t��Y�J���겆v��m+�p.��[�ŕ�v��g�;u��o�yWn-=�+��ĹJ]����v�}�q�я�D���ͬ��©�n=�A|�>+�]��[��U�rV���Sk�㼝[{YF������z�, X�%u�	�+/$�ŢL�������QT����.�٫�W��m��R�6�w1��<���b�p�2��}2�]�����(O ��A�;]5;���yA�9��vI�u�L�v����Q!�Ιt����l��Ǜ�T�n�ϹH�k�Y`hi�s��׫�5_����5	yu�f�Ŕ�+�i�� &�,hBv]3܂��u|M�BeW@7^�3gۦk� �[�C!�H��Ӻj�/e ��'q2��7�.���\ZW!|o&��9��#�]@�������-!����ʵ�`Ce.��cu�� %K��/m���E��<�t��̽;3-�r�u]`}{���[]i' ��mS�6Zx���kw]2�TŎ�tamB2��p���x;:��f�"fR����c
�W\^n��Y��N���6���t�'���͘�<\WV�޵{o:�R�ϵvތ;K
(�S)��W`��֕vAF�i��;�ۜ��c�o1tg8���n��T�U�˴(<�B�KЀ`Zrjh�i�ׁXV�e@���4�v%n�j�mn�ǖ�*wB���IZ��ls;�e)���ateb�IJyЗ1�fa]�}���hr| �[sF�[��k�*p����;mi�T���ޛk+�Z�L�.��q�r�|�;����+�)F��F�r�A�٢(����#���J'�䚣�T��Wq��m9���h��9�gsQ��"�wD�˺��:�c +��U,��
�p=&�X�-U�m>/W+TugR��R�9F��8����sV��2���;�2Sb��\%v�Z�����{�9C�C�X���E.I�[�Yײ�gOJ;mڢ�������[
W<��O7��� �aLA�
9�ܵ�߯yn�ʺ�\/����@��E��OR�N5�,�\�i����Z����=�E05��i����'�L��p��ӵV=+���
�8���H�&������K��>ŊRc�,������Wԅ�Gy0Zw�uMQ��y�Kxgu����}�#�N$)-}nJѿZ/��v�V�ܬ�DK"�۬�#�`��M�өQ��b��NN��x�<tp��}t>�3�7t�Y�ہ:��pӠ_$�)�%�#VY��α8�&��.���J�f,�ĕ��Z�|�\�y�%�����������ݐG��b_u��Ί�Bi�MwVZ.�˄]:9�� �8!ҳ��'02@�����TwC�Ϯ�pmm'j���h��k�a���[�;�Ig�tv��8��E��{+V-�+N��8n����آG:�t�VmJG�#v���$s��PR�5}��j.,�O�]ٵ0�f�,Z���Uu�{���&(*cЏu�	��6Q�6Ã�`{Z���ӂ�ӏP�D�t����o\6uhn��@:�{2�y2sJ���ͺ9��ũ%J�Mv�PUn^d��4��V� ���v���D��c�F(*�0�$��wo�6rSkx����"�N7s��Xʃ��ݝ������:�\���ќ�PP�b�4Q��v�Z��[��k������c�f�n���W�`Yj̼4����_d��/9Z!%3��`��tuq��@�5rh�[����5`�T9�7��� �)U���ծ�õo�]}R�vg^5�A�ʝ����tmk����ۭl����К����L1�(��-޻z��0j��S�K�X�.M���R�Q��$��h�ced����0&+g}���b��g!�V���Ԩ|���6WT�Ы(B�ky�yfgQ9׳��w��Ws�в�/�b�^�̈�}�d�VK�8<��>�*��gV9�}�wu�p5x��$���od�{-���Q������5��G�pv�Z�4����6�y���u��*�:E;{h9}��^��h�����f7Dw�mk�-]��`Z�7��tQ��M�=z:��&�)t��
4��p`Z��E�U��9g2�}�4B�o��n�|�Ҕ�;�D�h/�V9V�WR}jN̥t)Ѯ��l�{LV��m�r�a"J�lq�F�nweX�rܥv��$���iӕ4�� Ӝz,��Z����,b��kJ}Kow��KA�o;n�SV:Q��W�!�*�fſ�f�y�]��V�D���e�C����n'���2�gr�-r�O�C�ȶ�.�{��-�k�����3VIZ�&�`Y{,���2�[3]f`�P��e[�s̀Cb��Ug[��`�](�=-�.�m��X�i�^7ֲ���@R��e��1��DbnZ��=F�I}N,� ��;(��%TaL��M't6�4v�N�󽥯���:ݼOW����_]<�C[>���5Ԟ�d^�1*��T����g(�n�P�v�n�Ѱ���e���F:�+き-�a�j^f�.Sje3n���Û
�ggm�|-�uU�4��NT9n뼬P���ۗ�.�t�_{�v~Q������_L&l���n��q��;�[]gEA�}��C�L.:�����p4T�|��V�C��
�ixq��Vf!o]��#c0����� �s�_��:z�	@�Օ��$�`'L��6����ʻ3��Y[�Z˜d��;&�w�]�]�R(ݘ1�7��<�/����L�R��mذ���S�����b��Yӓ[M7|�k���.�'+��gaM��1��v�ͩ)^W�˘2r�!�1)J�a$ͦ�q�HV���p񡘣���A��R�r��J}0�Dc�T{w��R���լ��(/�%Yu�֫w}ի
7��i��IvwrfF�ҪHt{�6̮V: `M�]�A:������T��tp�'���̘[$mu�8�6���+�葭	*����X-�۽�ˊ�佳�hd���R���K!RJaVb;��K#9�)�[I�ƶހwe�`^p'��Ҕ�
�Q0n��r=�&����ŽWj�jF�ۣrt�+.w�h%���ҽ]�[����\��-�����5�X 9x)@���7���vB��,OR�[+8�0��>խ���w\����sib�l��L[��ҦP�JA��y��p@�ͣ�Y�����oHC�z�]OwE�.:o��/I<�ą���Wr��j�t�}�t���r�6�`�F���
��&���,pN�m��)ϋAgX��\��lI�i��{J�(���
(�6���csN��Wt�N<��̉�����I�gQ4Uv��"-ː9�cXq�Q(֝�����7]��ا��]}�{p��9u�pA'K@�!�\���Tr�t���mLs6�6�p\X�.m���ٓ���ݭ�٢Y(�j��v�Du���z-k�`2�v���|�
���QP���3�{��'z���A{�\���wB�:�r�6~b�g&��ro7H�2�}i�k5�:����^Tz�22{����jGa���:fkk�	�ј�o_]���e���fU���)5XVM���f�>�/���p�c�7jdƳ�LӲ����]W��4�2h�M��!I�>�Z�n�N4�,)�ff*䍪@$9��w�O&�*t��̴�ik�m�Ym��B�n����e��n���%Hk�V7M�g��)f6qMyՖ��	���7b�4��͜��k�o���X��܎R�jȐ���ۢ�t륌q:��Wr��!ݬ�t(���7�2)�^w>9+;�� �ǁ���D���s3Q�=�����sgN�#g��Z�YΦJc��ֲ3���]���SN1��;t
�U�ᒜKa��v_�R�Y;q`8	X{��v����m$����ʍ$�o�Y����`6��Py�7��jֶ����ۼx6ܭ@���#�\c���'6�[b̩��^kA3����Kfm���j�(Ț�ڸ����kk��R�A0��jRs@�2bf��Ϲ�o����Ɗ����#�4s/q}c�& ��'�l�61�������k�n�1Z�U,Z��[��Y��BA-21V�ЁfȮ@�S�t-�6/1�nݛ܂rN���>͐@��/b2�8�Z���x���I�v�_3���/���Z���,�%2�1�ͧ�+���S���<�+���:;�;��C�4rt"������V������&�Jδk^	���b�����k���j0�q�[���@Lw�D��AWS[ȹ6m�7ln�v-�r亱3�	@�E_')����'���
O�IC������n[u�8r����Q�e<�F��ܾ7ĸ�L���i�V2�eV�t���.6�;H�b��wY�o7��n�ejIp��q����W��j�)aC�D�.���7�A(ζt��x32�ހEx����k(������
:+FRgP��h�k%�-�Ui��m<���)�.mif��!'F�ְ��T����x�� �����ٽV)���C�jq���we)����+v�g
A�//�nQ��!�\0�9���Z0<��*�X̘�)m�۰��t�Բ�����W�];#ݪ��=l�)i�ҵ����}WCEX����a����X�7��)5��Ç;��+Xzk���O%r��T�(��e}�2��7KbR0���S-`�4�@�l{�e��T ���Vu�F̺1�3z�F`놮��,�k�e�,uEB����:�Q{a�Q-6�d*��{rƅ/�%q.[N����p�N^�qakk�b�LӔh�����lT�c��1kU�R�᳓1tʽ���S]�vC�أ�q���\1oVU���-�Z0��d����\2�_P|yạè�ڏxj�y����9;F¡e7N�A��΄Y\�iX��#m�Y�dx�sD�X�J���GwHssw~���Q��{u%>�j\��dy��*���Ыg�ݨ4�i��fl�%1}�^cX���d�:g22j�N��/�TP�Z�+X!&�Z���:q��5tr��R�W��z�r�ڑj�<|s++��D_*�a
H��:.w>�j�n��ਭ���ȗ��a���{�HR��oq�9��Z�e=���;x��b��B.�vb"�3J��J��8.��@/��˪;D���t�X�H1ZZs3tܦ�,�6�}hq�^��ٳÝr��]L�Ρ�\W��'��A`�z6��60�@�=��b}vVe�*��~|9@MҘcYٔ/�BŹ}��O+�q�n��67A]rc�dG[856���
��|8,�~�%Lڬ�܎�4j��,a�5ʒ�j�������=��c�+��qmh<��&���c�	@���{��xJ��]���hYݣuFҖ�T�l:Χ ;�,ź������,4$�w��S�l�k���_R��U0�ۡ�ݵ���=I֬��t{�<u�\�f�Mq�;{\������]}�6�J'����������Vy�[k.m[�����F�FŦ����k:9Ʀ��Tzi���)���]��sT���W� 秭�,���r�Yn��^uY"��X�G�K���uX�U�ŉ���6|���Q-\Q��C�4�f��N�-�-���*a-G�]�l��i�T�R�����K�;��a��1��i��}�	+lӗ\�=k���ĚU�k�}��V<��0�@�gެ�p<�LM�P7і���˧շJ�j�D�4RTYF�nv<� l]c�:U�zT��@*���#�P��u�f���-w͗5�$)��Y�pj������SF&]����F��+MA�Gi��&�FXr\"�lq|�ʮ��5M���97@�M=�؍nG���#
�g�=6����憾o"���7Ive�a�y >�T�Xq@����	H�3�y���8��Jݛ�Z�h�����%�.�Y��M7��0�:��Xj�W^�]�OV���9g�{�����������=�Ц�{)t��;�x�����n���Cq̭H�1Xs���g����h�s.��mќu��ܤ�8�0��e���ih����,�����:s�GF���=�<Y]�3Z�a=��/nК�`��:"N.u��x�z�߰��n&ڮ�u
�ډV8Xs+.�����]�̽�p��!�`���KD��Bfn�x`�XMZD!-��mwmr���ϘW:䧡6�־���+�{:����y�]�N���V�^ �^(���>k�8K9	��õ�aH�.�hhq��s	Ia��_n��RI�x�*,���hu�/����o:-+�F�۸�0�U�#�w҅a�=�=�݂�D��P�xZ=j��:�]ڲ�^\��k�_n
��u��VС����')��oFX�R�oD�1�6����L��t2aJ�������^�M��^)ӖZ�����X��qWJ�Ly�[��آg�vf���zF7ѵ&��Ԍ��v�Ɂm��t�*q���w�A�'��t��e�nSΨ\���0����%rw+f��X��i���ғ�������:C���S�6u�2�nT�zPN�m#��2�TG#|Ň��7��f�a�ݍ_)ܕ
��UŲ����w��Jܻ
]	�B�b���� [�%��C)\�Q	*Îi?��]2�躠��ݒ.�l�1�צ��
QS����nc��x�К6ȁAF�H��� 5�G6�Tk��D���Fŉ#^w9����m�᷋���I���+���6"���
�A�:�W,f`)5$HPQ���3�I��K��!Q��1�\��t�Q㠅�� �"E1�n�� �$$xݥْd�4gv���$�K�����fh!y�a��x���v�ڻ�x���^wV#1��t�wtX���n��A &&r�@b�q%�1��DI;���ID�$II1,���C4x�x�y݃B%F��H�a�t�H�QL'8�1�����Ir�1��%�JW���e�@��I$R�۔$d�f0P�d�np���2f^wd���!�ur��<t��T`.n&7���0wo-�ֻ;Nu+���ኡ�wwƤ�@o$Gk���������7j���F	o��QW��W���m
��.�{��}�y܁M*"�ǎ�e���P�R
�WZ��#R�\�h����� h]��Sj ˳ݱ+�Q�ͯ��}C�~W��6�����+i��U�ep[��gFr�g�HL-�}����X��u�&ĮU�Z�l��J?�����}�,����qX��C.��wW���~��="�����N�W�3M".���H�!C�9ɿ��}�R+��x�L�Oh�����3�DW��� �NÀY�w��\og;�E���:m���a��S���R�~�=��!�i���)�04X� �����I;�9��ʟf����E��V�������w��~�$��������l�{��LP�Jyܸ"��2��ݑ/׵'uz�RcE���i	��N�;ŕ��{K:�
���u�7��O+1�w1�c���:���l�� ��:ߩc�dҭ<	8�����_4�ׄz�q(ŸN���nݠ��%D�}o��������k��&�W�7�p0<�V��TƟO+5x�ۀN+A���Յ�gr^��|Y�5��1)�-\������>{��:�o��q��:њRv���5p����]N>7�}eN���p�: ���&f@&ego.N�{V�<4]�oP\[/8�l�ʝyO'k��9Χ�CE�hX��B.��g9�q�^��o{~A�ёa�v��s�Ҭ�>�B�����Mz5@v\��)ܓz����XLF��s�3�19���-���oJ���w~z�OY���ywn�oy��<T!��������������X1�ɪPʞ$?22(��S�!̉�,w���XN\Cx�M A�:���bem:7])�J�⽭c�K�j�����B''/ �����dd��+O���GWñXw�U�8�iZx\4���oiAw�{�PJt��Uny�&�ۨ�x���d�!����;��?){ ���Ԟ��zoor�{��P�ֻ�'v��|ɦP��VQw�a���]3��\'+]�(O���GE��7�֒,nˇ{5/�S���i���?�����8�.�e�νנ���p�PϦXHS;���V
P�DP�t\�3��23��]Wd����X���� Y�&�~��[��?�Ua�K�N�"8 ����Uw��q���v
������j9�VjN��X7T���ݪq��Dm`��R��i����#K}���cts����U�>]��1!�z��z�!�ft��ӄn^�ޱ�'�'�%��]Nu��󧍞Vtn�J�\�c�7J��������'݈����	�O��G'-��bȧW`�*d^�����o�藫�ω�q.�����)�#b�@h�;,B�9��Ur�{-�j����S+���°_�~uZLQ�ȓJ����KJi{Up���G9�PE,�ޫBg��!�����<\C/�岳�����^���x�$�ڊү��0]�+ɡ�4R��_elR�Pkڝ���r�ל�Gi�a��}QP:'j�����"�B��Tp�l�ɋ;!q���K��`���u���8z�\t,�b��@��Z맊�.o�'�G�)B%*�l�̬�U�O�O	n�E����N�iڃ]��6�,�U`��$��%|��^UN&��S�����`�+��$��8�ϵ�������5��7/*�Of&�j/�v��۾�f�S$�6k��h
��Ӄ6�%��: 1:��2�۲nuqp��O�ɶ�t�D��5�WM�"���0fcU�������TWLؚ������h��b+H�^�v_�9�F�y9]�h`����5�ڃ<7f�R������j�;�\�΀�9Y�.�@��2���Z��bV�c����1��u�z�LS4>�Y�����p�UvSg�Ͱ�f*��<Aӑb�m�Ĥ¥�S�'{bՋA]DҺ��Dh���{ua����`�z=�GNd�[�N�$�K7���X��6��]�`��eFu��/�]ЎDtΥ(kT�}bW�����\g)k��5EL�I��d���>�s�n�T���!��qa���:�_f�˘��'D�o�У�|����0�ƅ;:M�`������q�4��+?)��S<}j���衼��+���^�� �!�>�n�����z'���vd�!X���$�Ģ�(q���k:!��fg0v����,��h�?t�w���
pՇ[�lܤ�[	}�ɒ4�ؐO��k�.�Qz��K���a��P�)� �M���/7ʳ�Ȩ8}½�{}�t�HZ���ٝQ���ນ��=�X�aU���T�\%)�R���1[���mdq���*GR�ˇ$]�L���Q�4�����1�>��U�w��X��/��zfK�Sy����|��;���ܨW�,��*���T+f�+m]�́E����n���YR�΁���hI��d&9ю�*����K�ʠY:�Pښ<q�
��]�jw��G�gt7è-��;y襹mS��	��v�k�Ԧ���!��3wBx�p�]�XCg7�6�e:i��*&�� 7�l���������s0_%�e����ʞř7�[�
"¯�^��\�̫<��U��#��ޑ����<��<��qs��B�4��	��͇2v��@��s��N� Em�O�����T�AYu��Ƽ\��Yp�x��1WGd�m���Y"�6�N0S3����}�3~�X��k;�-K�A"c�e�G�P\�G�ݴ��J�(� �J��%J�)L�]�>uHBa�yru�D�ΰ"{1��૕�Wt�hkW0�'���D�
	�t�j/|72pf�V�Ȩ�\0���>=n��ӕ�mXݰ�V���j�N�/�`��R-�	���s Ǫ�� ����9�x}:Y=P|��ɸ�s�g
������L9����6�nK}T��q���U���0<���[���:҂�V���g����G�{[�s��N��j�w���H���x�_m���T��4��<�݂�^�gPWp�b��R˫��{�mk7آ�J�������J"��X`�NÁ���n�7�����:b�c}9�8���ʤw��I(�X
���Ϛ����p�;�}ޟ	���{~l\r�*v���-P�X��M�C��y��evL"��^B������]���<�ҫ�l۫ޛQT6Q�[�WN�[g����ܟ7�����U������f�$��3Q9����Փ�4TʼU�D:�pl���Tp&��4B]� �}�pE֯GFY�л���<Op?PvABt�N`w_�[?��$m��Y����!�jXĺ���T�Q�NW�v�LeܲN�y�2���6����,"Hٛ|Ȉ!�<��Y�+sK|�c�	����6�[����������.P���M.5�ŭ*J�u�^��kn�>���\�i\J+
#�Zڎ��l; =���Hȃ&�����teulߌ�{���U��s����Z�#���g�Ð�*RQv�6�g�v�f&�����,1";�����T��bu�G�R��
��ڕn��TNV\TP�sg_70f�O�DY��>�D�"D�c�GC���cU�&�C.Q"��J�T'�bP�4�ӭ����� �:�$k�d�[.�WJG�W��h��́���k�M�0E��n҃�����W�9.EJ�����ί��a�[�l��}����Ʀp3{�����_�5@ţ̙<u�5Q\E�V*��Z)�����y��͋�YJ�2��lv�Sv-l��Jv3�V�[L��^X�o�o*9�3����q[��)-���v��rV�n� �!`i�nc�.��o�TH�b��hBwWt�shq�;�FlZ�I|͝�9j=Ώ'8�[3y�Z�����VG�j��K�����G�I�ϩ�Zkگ,,���ϙ([� ��l�zʇ+M�@:xZs_/v�otq�ʝDl(f�\�I7eC�l�d8���}�+�?o�������]�7$GgJ���щ�35wӥ�Q;�|��srCӰQ�9~ε7�R�Q��u̎L�qÐ�)UѼ)b��g���ǽ������s!U�Y�?�5`��'5��;�������x�O�,4`T�R���T�c�+�Ո�g�踗Yec��?7�=U^�煘L��K7ۧ�n�Ўd�Dד�e�󎇤f0�tM�ܛr$�=*�X9nz;�<=�s����3��%PH��ו�.�.!��ۖ��Sw�/L��`5JL��"��K�.զ��뛺ȇ�.�;<΋좍�R*�N<��[��6�>�8ϝV�����j�ǅd�e5P4Y%�X;��91�uTĩJ�HR�]��
^������$	�JA��l۰�U���(�x.�!��i6	�̄��ｲ�^���_q^��HG~7L�s�(����X�g0�L�Qge��+��Y��'h���-���5�\��9�2F��'(��P����f�r�\oi0
�u�h`��oT��T��=��MS�9r�Wv����W�՝ֻ��8+7���I�]�wxRݤ���p����[ʐ���7FmNU����bz{z�6�`�S<'��'�@��|;�����+tI��b���ڬ����}�a�S�Ϙ�����@l�s��l6�,9�T�+������D&zm�βv�6Ȕ�����~���C4��vڒ���&��Qư
�$Tq��~31�n@Ho*�b���,ޗ�;���\�B�ӸjPޗ���F�Ƥ�iѣ���h`x�e1:y+�+���T�N��j�hk5k�_������gI��6�&c�[r�	$�7�-�;��b�]Y��7�S�Oo�$>����9��\����B����S��*�uS���y{ϐ�4iW�����TƦ��Vx�.x��[�s)]+Pw�2��_T/ҷ���[��V�fa��㪤����N���W��Lz���v��8�/c�ʎ��[���\���ǉ��VJ�L�v��z�ڿu��o�VFErp�*.u�K�Ȝ�;�l#���s*����T.�%D$4�p(r�˃����W��3�`��,O֥t�oH��^Z���R�E4�a��^v��5!X�w��`+��R�U����A���*\��]�C[X�,�b�������ĮA���ٛ>f_�-Gwt�ۭ]�x�%�J`��[�S�[J�!*�]3��\t�Ӡ��o:��9��+{�M�W�ھ}��Zyΰ�+�=EA�
�SK�5����pu���×�r���:�j���0l�׏i��1��{��k����T~�(�|'�-�(�{�Ou�p�d!�HQ�p��1xd�SP�t����%nG�����ĕ�|>!N�H��v6��ob�׆%�A۸t.����%�х��/k�����wHڳ�x9W�?��kSƶ��6��b��Eab������Ù;Ny9�^x�c/�i��`��8�	t`[�8CnK�5�r����*<�������)�dd�H�s#"��*W�y�ܑ�j��P�T^�6��n�;�Q>�b$L�ޚ���GA[��m%��F9j�91�������Ū:D�Wj�f�r'A�:�L�V'|EzNÓUr����P�Z���>��2]���+6����J����
�#�"��EX|�Z|N?�;�T{U�׊�W�a@���)����b�s૗s���R&�JҀ+�R�¸zhB��}V>�7��;�l��A�[��G��d�u��4�DF.���7h���W��u��t-��'�)�	�ǝ��l��{����5����X�h*w��`u#zv��X{yL�-�Hf���3�E�#��Z�K	��w7����4�\�P�@l�jk:�Vr{d`ѧ��+�vH���ɲҋ���b[�Uc�Ӑ7��Ӊ�B���e%�qzV����+B1p�B�ݽd]١�vf��ܞlާ\��wJg��{�
���+YZ7�Q�X��5���j�*^;����r\]��>���r��������J#q��NÁ�\�=����wȋ�Z� �ؒ"��6��]Ԣ����k�
�<�ٟ5�	���ޝⅴ��,:��S�'$�^�R؏��n�̦.3r�M�e��f~�1���,N����;�6�}Qg���W�rč���P�	�&��W[�\|�x^ҷ��H]�\I�BO3O�H|j6��.nl�5��.u�۽�UV\�oJ�Ɵ8ya�ȹi�i����iV��%�W�W>԰�Eh�J�-v뭙�I�]04��Q�45+|p5%��#`(�}AGx�E_��5��8�1���I���7Yzջ}�s6!�V�}�V3��x�g��Z�k�o��ҍ��n���t�1�n���UgJ��Td�XH�9:�s>�;�']-���oJ�nwI���ȹ)T~�����2�RXU�!��^��E��o5&��u��%*6*�_^�IV�#�I�
�������MC�]�(��̽�M`;�ŋz�{�k戁��.�Wiy���6t�9�O�C�'N��!b�����әչZJ�����E�b�����Y�d-bVE�r�,u���v�Ju��y���
4�V}��Pwd�{�p[��*��Qp�6I�n.��m�}�hj@�Ю}�>�|kk����=���M�[3���b�)']�0Zt�o-��#�c�˹vB���ۇsD�Kb��F茡*^����.�;�gGK��WL3sz�5*����_+�VvO�u�e���@֭���u�R��6,Ay%K|�T�iE���\���6�`w�8���r����''X.�	v��kE;��
B�!ږ9���'��+:o� X�jEۢ'N<��ˊ��Ĩ��,���@�`NT�|�:]d�[4��`^���R��8Eؑj�&YY�kx��:h,�rq[�`B�s��֪۸�mkt%xV�jp�j�`��	ΗE׃��ϕ���'r�e�\�ZN.��ܳ�WqO)(<�� �L�]h�4ӂ��/��b�5��;����j����V��o]$��l��/p��h��"E���J�v��4��;$��|�qėR�qf�ݭ�ά��#��v�!:�Б�ܫkjm5,���wd�jNge��4d�F7���3��6.Kͣ���9qځ7�d��4��:0i�8wH�������\6Zj.�ُ�NP�M�O�-��Z]m֥Aq���"�B�'.M�Qw]J�5����n��T��������f�F�h�jk�t#���wC�\��Ƹ�^�����W���c���]x��^+���7]�7@��B�
6������N��b��mp�b�N���i�����
ym��wBpU�}v k:&ڮ�h
#'{}]n_.ƻOVn��W�L�-w��sd��~�Sj���b�76��wZ��>��9��t+in�`u��aX��[Z���v�;��Uq�<��u���.h�PC;x)\�[ʽV�M���;T�s�1��F-�@f�����5�>���3;��J�j�5���F�u���a�����X ��O�g�ӕ�ҷ����8����9��m��<ө�`U�D����ۘ�~���Y[egM�t�̭(gn�:��+e!�7&T�����z����Ȧ�j�Բn!�$���p��"�v�}����`IBu��V\y�uu@����Uӛ�قX�K2VP�r��%Ζ��Q�Ŕ�����;2�-��e-�9�Łn�,e��t_N�mM��{S ��J�G�®��s;�E�,���9�3�P_AJop�5�\��<�6=���Y�߃Z�4hU�x�%z�4�Ah��NuӤ��J��S��N��7(�hZl*�[b{��|��85r��w�)�ř� D DDZ.WPLN��&D��h%D�a��i"��bB�$i�$�4B���`2����鱈��D��m�\"�%s�\�
FHѤ"��QIf��/�J521��2�A(��II�ɑ�^whAa#��
1$�4D2�	��%(�
	���
�ř��	��	"JB��Őc�@P2H�\�0�;��&C&��LIwtd�D�$���
1)n�0�ĉ
	� ����g.�D2R2��%C)��û�.��u�E$��#E�Hh�D�If4-� ���R�cb@�P!wp�#	�%��6��I6����
C���34p�)ӛ��̘�m���x�i����I����u�va�8��Z�c�ǫ��РN�8-odb����VS];e������z������k��x��|�x���^-��������E����ţ�t�>��=p�
���@Q����d��C�{9�Dzc�0 ����y�G�{�&��:g���d�Gk��q�!}"<��y�-�W?[x��}��ݯm�ۻ���������{��<�}x��h�j-��W���~���Z��z���׵�okſ/�W���5��W���<�Z�G�gnY��XV���_�ʎ����#������V>/x��߾}^���y�����{[깹�w>wT[�\���:����zW��^��oJ�<xѧ���ܷ��x���5�j5����W���d sV��>]F��f�ľ�P���x��{^>�}�W��W�xߟ�>����Z~|���{[�sW�Ϟz��}W�Ǧ�>��Ms\�__+�[���ͽ������żo[��->w��W����6���к��tZ��\{3���Y�q��>�n[��﷯��������~���]�|��ވ��2�G�xhO��~>+ţ�_�}z؊��W����z��������������������y뇶 �Q\�"9������\e$�3�/ͻ�Q~�ŧ�_�}��C�r����������r����^���^wO�@�}�MH8G��}��߽�������z���7�|�߾W��#��21+�/ �]�����XQC�w�Z�߽~/�^ץ���~_z�7��^/�~�W�W���������^->u�{�������{��+��ͻ���~{T� y�<c�6;~��=� `au^��>B"G� ����tvgW�D��Ox�>�ү���F���ۖ�/���~���ֽ�F�7��zW���[�^7�x�+�������Ѿ+��=�u��+��o�[��[��ו��[�^?��
�0 px�0,)��w�i�l������|>��}" ��Y1� ��p��K��G��+u���@"��lz�6濿���_����m�r�[ǋ+�;Ư�ߏ���^���������XB"G�sN�B�M��C�#w���^��߃b+�|W��}�W�������>�����^6�������[���w���6���W�Z��7��W���soW�~�K񷧍�mߛ��|W���^�t( ��"cocv�ܚ��F�%��U/g����t���N^�;
�J��*������<��������A��\����E�9�Z��V�]BM��v��jTF���B��j/-����dE�l�`�S{�[H%�cSr�e��8���O�u�Y�u"�6z�q)�j~�G��(��YG����h��������x��|���okE�~o��꽷���j���ܾ�����x��~���}_Z�|_���/��Z+��/;�~�Ư_���W,x��x��Ͽ^��1suu������ǁ�xǔ'�8��ywo�W�\����o�������۟��)H���ju�8 ���d{#� ����(����c>'�洞��o]����6�}c�#�b ��\�Wη��o���^��ޕ|\�5�w�_���-�{�~�W��o�����xE���}Cc�=� 
�s��׽�xǶ=���d_yǦ�s�ٙ���]y�F�i
<F��G�$G��\�~��o�<{��^����o�˺���|W�{�������ם�i�7/^w�Ž�[x�W���,oｷ�:�����#�=�c_�<���B�s��*��Z+؝��1T����>����T���}m��Z��}����s�������^��\�^����{�ֹ�7��׮����W����wu�<c��}m�EyI�.=��#�����	��t-n~���~�Ab�T��ȑ����>B�}Jܺ���xD?�z�ǃ�&=���ս\��}m���U~�m�m�u���[~-��n_��ׯ�Z�^��z^�x��[�^9zm⯏��4nm�������~��3F2�t�}�_
�"G����C�5�@��x��3�*<��� `<�\�Z7�����~7����>�����徫���^U����������5�W��{����|m��+�u�so��{�����Eؗ��!佫w�M�����Q�W��mʾ����6�noM��<��Q��=1��)���{�`{_P$x�V������ޗ�G���ƾ�Ƽ{W���}�ޕ_���v�����W���,�,7�o��M+P�H���"D!��;o?�G�Z7�F�޷�x��������sy���^�������~���� ���s�� y�1?���Dz��:��'#��Ԫ�>���
�(*r���#��Q�x��������m�y�����/�5���/KF�����^_��W�E��_V��5�W�{�y�>�ֿ����}\߭��e��>��|�Auݱ�O�;�j���OR�4Y�zc�U�C��o�Kf�ؒ�<EnZ�p)�	�j��p.�c>W�|\>���s헧\��G�:Ь��J'R:[6�C�3G��W���v�V��YҔ5��n�����ꓹ	J�n�3�ȀgQ/�<��ܱ���~��	�=�K����M�}_H-�ەx�x����{m��������5�^��^-�x�W��}�~u�o�}o�y��W��|~^���}o��=�Sꈏ�l A�
GIv�]����nl#
���&����@���^z��__��-���KC�m���߿=[�^֞w���;_��߭�o��y6񹽵��z���w����;�r�ؑD1>1��O����P�y�	��ʫR~�GG�G�	�𺚏(�p&<&>+���}yW������⽭>��޾Uz��>�鏣ޘ�̏�k>��0}��������������z��o��9�E���$}�8l���%��g5���������DA>�LP� }}��L�����-E_��B~��
b�+Z�龶��|~_�{����
���<��Ͻ^7���_���*��Wּ_����˖��6�� t �	����y"~߲��\��%$���11��	�}�}��.X���k�_7��7u�߭�[��{��o_{���z��|W�;<���]���{o�ܫ�����F���������ָoϿ|������7��?ߟ��qn���@���{#aE�M���G�;���򿗋E�w���7�x׶�k��~��v->u���W�^�ͽ����=��K���ƿ+ߞ{W-�޵j�@�@�#��~�{����{�b�s-��w���T���"�}����������������|��Ƣ�[������_�k���wk���x����5���^w��؋��x���X��Q�8p=0���yC xDz~>����J���:َ<ۼ���[��}R� |%�{��������*H�=鈏txg��/j�\�6�x���_ͽ���ߗίk��[�zm����~w���ݷ������o����w_��[p���ÿb�f$Jz����G��GӦ"G�>����ǁ�tm�C�@���@ʯ������x�������V��_���|��׮��������o�^�7��>�z���o���ν7���sQ�������?��~��𞸫�Y׻��۬Q�"��>ܷ��^��4n[�~��o���k�� ��@P& CZ��Dx�4S��~+꾯����������_ﾼ����\׿�|��kO]o��_z������ �0����5����ؘ�ޫb�P���̋��剁2,M=C�ei�s��UQ�Y�Nj�A~�W�un!D����$@�Zh��eObW�6�&��TMJX.���M:���a1��meX�`����Urug�&��]��)���YV���8t㕽=�׶�^>6����^���h�W�x�U��u�����zom��~y���m���_��[��U�{o�>�z�E�[�������U�:�/��ןV��k���iݠ��>�"G�!�b�����˷�b#�_��{Z����W����~uxޛ��o�������o�;_������+ţ���/�����^7���ϝ6�om��. ��{��T{���?�W�b$�@鍟?A�f��Jt���?[x���}�|�zo��ݷ�����9h����z�:����m½_ݯ��W���w�k���k���_V�/kF�z���׵���xׯ�׃}[�潯���k@F ��SOm�)���^������ߪ�.o����[{��鷋~��깹�|�U���=-�\���Ͻ��y�U�r�.���<hѹ_���W�ƿ����j-�~��:�-��s/�}}k"4D�����NUhܕ�+ݯ��~����~+�x���W��|��V�~�������+������|������������\�/�M�~o��kڹh�{��<���[�\����z^��o��.�7@�'#ިpDU�c�_}YN��Z�s���G�Dx�쏼(�� #�=k߭�o�x���������}k������_DG�} �މUPC�&q8�k���紘��F�pOǶP��g��{ ��>����S�}RT"r�u(��`q�];	s��sQ�a\Nl엙��M�]!VL��T�a��(�@|TP��>����,� �oN�B�w�º�4.�9)�3;k�V^�S��0�{��n5�C�{���M��u����*��N���׭r�c��� \"v����WO����o�U�>��8H�`����t��*���k8T�ڛ�M����V�ж��e��*�|��[�8Q�V�r��.��̖��!i��ڼ:����^�BqկX�����%]N�[H��`h���Nư(s�����Ԡt�tN����@p]�Q|�>cW+�%����76nu!|�9^OBl�7�a`�t����,=������[����������n�����w59�-��l�29��Dt_��B5	���Xut�V��=�kn8Y5ǬN�fj��(-&�K��NM�v���֎�.6y^*�g7^4g�!�t��sU��>�O)Y�/�*u.F�gX�����$�|G*�3B!i1@��S���X�ttg�����*6��VGF`��i{.��W�+��qx�<`q� %���A�=G ���<�V�6
��R����!��w�V�fW���(�FB&�ۭ��;DGP����[N���H��\���yV�<ĲO}�oi���P����h)	@�<�R�<Q>�A��q�Ff�Y��)�qԊSu��RGq�/T�<�׸&��Z�dɿ��07���u��%b�8���͝���ӽ�W��]�!,*�����ep��Mxj���:�!k�2h[� �{g-��N7��a��e��Г55&p��U�vV<+�`����j}��zbbËS�5:�!+-�:0�lAv���쮡��1:������I���S��;Y��gwdB�p]������w���bdT*�r��&�R�c]n����$�(�xZ�yg�3V^���j^+�.���,T���*�J���B����E2��dj�ìCI6o���&�b��9辺��ڹ�?<N�<����肎A��u���n:
�+Y����zr�sŽA0��+ռ��Orb��}H=�\N`5��s���:Iw���*VK�]���^�╈ ��"�{+�C��xk��]O,�>S
ߙ�:.%�YX�}e�y`������n.�H�^q�@�/�e�W�Yd�jy��ϼ:Q��̕�Z��*r$���;��<�^���Zt۷���X�Og�	�ו�K�ˈe�ܶT�^���C���dg�޵%�0n����[�A�V�CEp�k��l��S;���Zp��L9!Y��6�����F�G̭�QW��A�I�+�T� a�Ӫ�%*K�$\�Cª*@��ќ�rrO_�98z�q�p�T�+���G��2�)V�9�}�U�v���q�wS�Uf�K�Ën���Ga�1���'�N��8�=�}A���kw��Yp����LF�>5����9����;Y�۾�f�I+LIPx>�īn�3��Ay�_�Lͧ��5Յr
�t&��k�8�� ��2�'��jk;q���R_
��YgCP��Byo��^���^睦^��M�r��RY���*Su�S�Ke*A��_Ns�m�=�ݼCޙ��ΡWT���g@���]������I�d�`��BG`+�Fol؍�#i��&�nGC�s8�y
�"��D�n�����%g��B*A4��������<wOoJ�as��|jH�i٣~N@תlh1e�
sE��)��B�s�d��G������i��V'���8]�h��H���g�\p��^N��h�b^���	u�+?���/��-Wl�,���vf��>��n6:�%��_�^��SI�;;-�p/��C2�\\5��Tt���NT�f�wh+��4��&�Q]�%Sw;#�#x�X͵n3�f��i�5]�ب��p6i���ھ~���x���ʾ*)�u\d��G�� M�V	SI�N��[j���8��U���9Y��z
�=���.M8{�X����l	�'rg��FF��(R�Ω��.���10<�9��s�f0X<T�[��r���ixSY�q��`���8�����y��Gjp�2)q�N��YW��ݶ�����+_	M-�c�z�A[��oer��G��8ލ��H^r��C���-�oQk�Vkv�McF��J}*� �|�;[�Y��{^�\��s�����ji�x�7�W1H32�x��g��i|�{�b�`ZS��K��Ӛ��!V�������Z��y����9��x�n�jH��?{�{�W4��ꢭlg:/�c������7;(�88�J�>C�z�i"�4�^;���(�h8]gМ�-���ai�1��U^U��1�j"O z���Ɓ��]��eu��_x��x�&�I.;�$8�<�@�8��'�>H��+�s��{��pq:Q�_����WW��e���/�]]�Jv��R8�Ȧ�	ۛO��1���Y���IN���#e�5�������/�Pq���v_m��(�-Yet�_GH6P���5﫠���R׮����$sl�$�95W+��ԡ�֮a��3#uc���M��0l���"^y�q�Q������3M��(J��8+d8�c�%��+ɵ��d��Źz9tԞ�� 8RR�¸zhd��m���Ǚn�R�=�7r��$.գzr��"�ԤlU�P�VN`r>�,}o��J�ؕύp��}͒��~�����{�_yҏ��z�I�oJg��zm1Z��w`��zx+.1��J�Ӌ�XǞW��w~�}��K�o"j���%�������{�}�Nblؖ3����w�ճ>%7�s��,ǯs�.�����v���ŵ����E�L�굏����Ag~��NηV��]���ai�T+��ݠ���� �|���̚�pp��$e�H���u9G��=��gR��n5��	t�8%�#�@�NT:s���l^����[�Y�@Hh���L�}T�0��&�����G/@�Ka+�򅨃d���n�}�ߛ��Y�m�	:�|o�
�q<gT�%�t�3�6�m��Ō��Q�Ǚ1O'R���b]t8ܜ�MFw-� cpO���Ȩ|��0��6���.!]�Y���>p���	�Z�ӕ�� �"x�$�`'l�g�fOo>�jE`WZ���\=��C���hMgu�+�EaP0G���ㅓ|x����V���'���w�.�(����D���f�)-��z�� �z2/oA��lt]��
�VlևJ�$�J|#bIӰ �� 1�H�9:�s����룠��2�i���x NL���λ�����ϥ�����y�Q��p#CP�LM��5t�[Z[�<A��oU��9t���؋��AduA�F��12��=-�%�=�-b�;Q����UA״��Aθ� .��P:8��iX��Xy:�VXb�����,ګ�j;I�4:�1���Uv+�fwa5.�*����s�-C�q����&��7/f�,cR�l���q��ׯr��wh�罆q��y�h�����h��o�f��v�+��b�Q���IV��� �Ƭ��)֮'��;Ŏ�J��\qn�i�*�̿?����w��^��_��˨���M�@�_#T4Ev<��ji�W�q䮥��g�%�ܳs~܈}�q�!a�WC�����s�Mr�Ic��/D�8mr	g(�C"�6_�,��"FB���er�$^�zf�߻}L�	�K��hJG�wo��liף��\*��9�(��|�a
�Y^c~��XEC�v}{�X�	xgtx��\6��;�q��E���4潯bi>���B����5��v�]�=0��ֵwz槽|N�#@|�ȿ�f;��xT�S��z*o�藫��>'E�І��kiݽu��G+�:UL�)�ge�V	e�MO2�^_�(|Ff�����VN�A�wp*d,�c�]ް��(&�Й�Ol��H&;��_u��R��p��{ԕ��⽂�]�]y�cx�h�4���0w���*�zy�����2��:�8��Ҍ~c.�2��޸��ЈWY�ꛓ�� :û!s!y7k�YU�Z}\ѻ�_")R��3_r�]p�Y{�&\�JXӷ�9"*A1�Kdۚt\Uм�rm�6pJ-�{�yw*�qk�Pҧ4h��J�X\�oP�)��_f�9>�S�e�Ad<F,�@�$^9znT���f��ؗa��u�p�,PE+X7x��d�����#8�js��g��Y�s�b %V���^0�ᴯ��cSD�nS��1��`�aUNÍ�;z�b�Ov,<Y�'��Y	�5f��0�wM��ΐ���؁�5�3���e� ��=&�5ۅ��P�j�sf���/�^eK�L�˶��V'�	\j�����q=���w����6��'7���y����q�㼨7:�SӚ5�غ��nR�ŗ�:�wa�e��L�*e4Dn�Gct�=�z�Z]
��7D�(�AA��Fﶦ�ݨX��k`�����[Ǥ�βxT�!'(�l<�qFr����p� ɵ�*h�t�fK�1n��Z3�y��,L��2����z�b�	ˡ���7��Gt�efF)n'�f*�x�vk�p8/��4��K�}���5Gx�Нi8�[V�p����\���50�^3�3�+{TTX-����:/R_<o^�I��{��T@Ai�n�kE3�"���7"v>=�m%w`FP,Y�y�J\�r�&��;ÕIj�fpWe$�c�{r�aO[7�
]GR����wP�u�7k��x�2���5����r����Q��Gl0e\�Z���2:��Y��B��3�xx���,T}n���c�9I���K���H�o6zB�_6�j"(K7݌Ǵ�V}��>�	Br!��<@�X9R��/R��#��S�j�u�-�����:˻��M-+��\Et7�`d��"�Q��<�ҖN=����)��[�㗃T��"�+����1-�U��gy��u��^#�TŸ�n�233��wZ�4e�wnXm��l k]a�cαB�J��;,�1�6@
�F�)�|r�w�o���X;��.�ǲe�
ie�'G�'�5��.�'q���.(��>���ׁ֥u���N��T�}��9>{o/Z�ljĲU g8��[�V>4y.���1<�i|����xL��ÔT�,]绵<1�3���c=��+fزs����a[nC�y��6�W�VEgV�Mu}I�p��k[��p�����k�L���]�rs/�)�y��B��"�܀l��h��L:�Eb��u�����DH��;�l��;�m�Oxb��鱵�f8����Pnp4�������+2���	lx5�ק�l��״�Q�%Ƴ�7�|c��t�tZ�8V�K�չ��\B���e�%Ԫ'e�E����^���Ʋ�JV��DX*�(,R���wѨ�~Ջy�,F�b��8[;���v�=��F���X(P @��B'wR�C&eN��D�����FB0%d�P���2LT$(�ː# K9�遜�S�쒈��ݑ$�2�wn��L$� Ww2XD͐�	�D0�&�& �4�E�D�Q43b��a�S)���a�II(�ED�2��C"R�s�ID$���#w\�H������P��S&a�]2A1BX	7v萤JS(I\�iY�t��1���IfL�	��
l���R�쒘�e�QA!�T��IBCH$$0%�B\�F"�fl\�P���
���Xv����Rڴ���m���s��J��.�B$6��oP���K*4�P���Z{�å\ۛ���&�J���{�{±��K��������v��+B��N��
��TqV��5K۾�ZZ7���|���W�+���}nSDc�8zt;�J���(�>�!�
U��e_E=���]]w�"Z��$ɳ�����M�v:�|s��K�D^}^o�W$y= 4����М��.�>�D4�e���xlWT>,{��o�9H�nE���w�� �%q�z���N�JR�Z�^��b�� �1=+���Lߣzֺ����6�Z:��q�)M�ٵr/+�%fa�d��ٸ,���#4��ч���;4P;�n�sY7uq�����FF�4�40P�xd�Y=B2}�<�E����_?a�pp�Y�}�V��E��]�#qR�W��TMl��k1�4������γ��/��-Wl����Ὃ�{kR�ͯ[Z�w��n%�"��Y*,'T�_�:�edL.���XQ9Pn9� ��UZo�1;K��>Ԕ+����7�q�4�EX�^��/'Ozɦ�ˍ�W@��s���1t:\ ���pV<o)�J���:r���q��c��j`�+m��L��ὖ�-��-�G�������Y��"�z��;�J�B�\���;|"�H�7����36�ˌ$Y)�k�`�6�7�n.y��v��t�N�}Z�9[�6v.���ٝ�����Y�� e.���J�(t�83�;o���'��%T���z�]4�d�1�����o�;O�Ѿ�q�OJ��{/i]~�	e^g�s=�=!l�ѓ<^�"�zy�RGTD�I�'.�KQ^�����"��5@��*.��:TI.	�P����f�^�ʫ�ݯ'���q�P��U����vT�Z�˙��f ���"�[� 5Z6���"3R�/=
����j�*b7��f�!�X�Qm���bnv:(�:8��~����=š���;��ÿW`�~����j��RY�L,<1��U^T �=^鈇��"6��2�p�A��u����n��.��ST%	���s!�i�� u<w1��xd��)l=�q������S�v60��b����^��ʁ�g��;%;l�+e"��F@z��Z���Q�0[�:���:&۪fb��,�
��i �[46#o���V���iw݈�Z]YL.�"rw4���i)��b��=+��&��Am�t�"���i�5�����M���V�)i��>|��ʆ��';�/��]����P���4�$���˧� j���m��Bi+�3+�5Ӹ�Z��,N�>ҥ\��\���X�?�3f/zc�/���a�F�fn+}/H���b��^��zmnL���k*�f���������v"�S�f:?UPmS%�f\G<`dD�TE-<N:�P�2��ӥ��Q
��y�`dD�����P�c���Z�یMUɸ�@��0�qʱax�'�N��`�UwG͗��[��F�o��uen�T�U��H%�09�C�[6f=2��$>��xB��&;��g�r�,WR�x�t�{iס�������U�� �)��/Ju��C Vȸ6\"E�P��&���C&�:�En5��K�a��6.�j��:���l��T��,W{M��q�(��ٮvM��7^�����ʦ���*�p
R�x��Y�;N�mj���:���~uM��J��m=��q�2��=��ĢpW3��*�vΗ:v-�{U�O,����G�Yh����OhyN.zgNW���c(�N��̦#���sY�񪫕J{����r4���9xP��,=��%�q�9[~H��*DyPz�\;z=}��/��I�z!��C��Y.�D#P�����8=�<��u-o&j[��apw�/\{�����TP=�Ɏi�N����Km�7���=;Fn����jqQ�@�w=���{+^f2uux��|�7��_l�W�ސH��"��8O�՗�K��v�q�5z��o��,�V�-��נ:�V
���ﾏ��c-fN��"��vǠ��<��flF�G��c8)��[=	c��U�[�v熽�G`�>�RQRQ���wP3�-&/�g���g`P��F��i���KC=<�7'ޭ3�F�;��z�OY�D#>��"t�5��4��~pM���2N�q��Ej��l��Ȝcz���i�Q�]"C�p���lE��0!��<��Ʌ�tg1@��%�lu3J�;(�Ny�J�↴j2��4��z� �|c�t�I���>��S>�C�N��sr�P��PN�*HH����7����T,<ɣͺ�灚��X�fm�c�	��\T���be7H������z��??��O	x����yag'v���|������3�R{�P��c�^��}�2�0y�@�]̸��UV8W��oy�53J�ŏ8���I��{=i���[a�:�!k�Fߜk�CcI�����O��a�����ׯ���k���x�7%�={��%':�目d_��Fi�}^��u1w҉݂� �^�tB��q3<���l���4�1d�_5����g[�S����MK��f`�^p�=�7�\36L�[�d���7�^�O�j�[��ஏ8V�h\h	fb�ѓW+:C�;�9�Pf�өZ5D�
��:%ѣ�.j._u-Uvf*��O.��~����f=jړ�\?|��'m�S{�Mw�xT�VU�,s��gN�(�z1�I���ZM.��g���f�Q^u����=U]���(�Y:��/��/���������*��N��PJI�ܒ��nI"A<:��u2�bⷨ�b����P�-��Ev�1�3;+%���cq]߼�_�
5�t�r��
¦v���(�"`���Ǖ�7!rV��ٞ���1]я�G�����g��
�O�:�}@��[�|�/Ztuຜ�X�T��j��L9R�"�O)�0>����A��H��(Џ�d!
U��8�*�J �M�]w6�,�(9�{��>�7-�������I^{ �9��d��q��D(,S.����j}�u�`ʬ�q��V�O��{�N�8�@l㝬�m���E�V��W�)a!l������~��@<W��q�͈ނ6�]nM�#�8��q��{ԥ���{9�;C��d�C�Dp�Ո�ȩRLTZ=�^��6:0�ţ^�-m*x;�`Oِ-�Y�c�xSV�Fkv���|�(�]D�Jo}ךH��{���(�5P\�Q�[�2�..q�m,��Uo;�-oT��p⍩.��F�|<�帎u:��-+����;�i�ԣZf	ԫ3euGN�[��}������LƷM6bc�(��@��h`�l�2MqD���>���ub+��2�ş��E�{_wY^�T;g}�Bλ�	�) ��q�W3
'E��a��0����c���g���o[����2��S��٫Z�ťT�^'P̢��l��:��{
'+�n9���r�|����g�C�\�����-����A����r��jY�9B��ɕ�zV���:$�*g��fm�ƀ�}G����]��ɐ$_5a�e2�tF#�W��� ����':R犾.U�b�{'��2ź	}��Fŗ�{U�\L.�)�.��-∋�C�uM��ca$rJ�x���,8!ݨ3��<$�#"s�qC\�#R5�Ed_v'�����C��@�ܶ{)�CX�^��D@��F��p���=Y�I�MFa���v�S��m��m��bC��u�ۿ{Q`����u��<�x3�aO�͇X��%ר5�k��t枞�W`�t^�W�T��jK#o�h��x��m��*�N��M�0��+wH���	[�P~'*�{º�}�n�Z�gVW;6%I�P0�r��,)����lfmnY�t��r��8��<
���X]B>�D_a]��it)��)��s�;R]:2s�j���.�V�Ӝ�Et6���H��V��K�V��� � U�-����3��
GG�9jj3J�Չ�2�ۙ;Ny9��~�Z�6��N�3��`��#p�j@��O]R�B���b�t8^�W�]S��b�s�4µ��0�r����#`?6�N�UH�"J8��&&O>��j���#.���lJ2Oes�bm�;��[��l9����Z�|7�J�7�T��`���v�r��w
^����;ז�f7�juG?&�aE�z��%L��ˈ�`dD�:�(���(��{���!%؉R;깳��=��w0�JB���Om�jjJ��!E��ix;W�x}���"�sz0����{2l�G'���﵏a�٭���|R<��B�nZN�Nju���e%rB�d�L���T�N�ɵ��"����#`tH7*:�>f��竩q<s�ҙ��n�`�H�4�k+�oq�,��%�ˏ�+�6�F��(��B�1����9G�$�2r�u(��k��c�+�#�r���o	�u��PE��n)�8�8��EW���eB� <2?�G��ʼ5t[��d���=t�X�A6�oK�u������n���AL"Z�{^����V���Y:�D!����y(���_�Զ��W����-WTU���ka�Yt8�z;��[����k�[��k��[]�]wQ����霤)����	츿U}�W�|��9f��}�o���SN��T�����;��L�kL�����ȮZ��tf7�ҩ��,
j��U�e"a�ֳ�nW��WJ���/�o�"�N�Em���M�y��9��c��#x���ij�#�=84��Ǵ5���4Ń~��>�d�Rd���$��' Cv���x�[08�ø�MJ�Ie��#`(�e"�3"/W�i��靄��9q�
���@���<�؍���-��p
n�a��q��HM	�7�2�j�	D�I�g��=g�2$�{���^d-&(��S�@WX�Tc3׆�N"�l*ӷoW�V�~n������ϧȈFG���i|��Y�aU���z�����͚�]�ɫQ�r�,224u��	�AduA�E�==�8��Y|��Mfq�%��7�R��J��kF���B&�IV��� h�1�:g��9���u�ʫ�%���|���}`����9G8�+����5@��̚<ۨ�zj���HۻM�<�qce"�R�1����R��P���ٯ�͒w[IL��^�:2�g��H6/�Ǥ��#�fy�>�(/]�13kb�2'��]]1�y���[�ƾ��
��Pr���9N��E���z��i%H"���Qa�bz���΃�3�#���}�x{����G}VrG�I�#N����+r!���}e<�ci�F�Ww��X��F�B-�g�}�,���X^�x�A�1���"��X�F�f��XMgً��_�K��U!s�S��-E�dt?-��0kuB�u���\_��NJ'v�����ԇ��or*�ݶ��f���mT����8�9Z��q�ps���=�i��7�rɩ�der�>�t{�2�N�}=A��}��/s3��_ �{����$p�����碥o��6�pp3|ً!1P����m�&�z��4�
T�3����+%�M��}�<�8V�7tFS옛��"��%p�f��٪#�MD�UD��'"}���T)k�+�����xf�b[���8nx.L���H��>�u�zg�v�B��q��/�����m��>T�>^��$X��`μ��H�܏>�t�3�Dq��.�[�>G�#D�D���wIs*A�:�j�HhnO;�x�b���.%J�W�|t!��ή��%<I��[�66c�Eq;�eT���ڽ)�k�|:<[E+)��h;[����7�B��0��爝�\�P�]�י��i����h�ٺg����J�;��R=�F�~Tʶ1a���d���v�����2��[�񢯷r�{��.X�ΝF�M3�mχ���V���R���Hh��B�tb}BxKv:-�����G~{ �y�	�G�R�מ~ע�q�p޼�a՚؈����(7��|V�O��\k��N�8�@l㝬�ۭ���-I
1j��Ü�tL١t�7�IZs�`�l�
Ҹ�n��S7�ނ6�]nM��tq�W#�]�تT�\�FN��V]5Ď0�cV��
��BE�jVj�3;�6�T�9� ��׻��0M�7U�6�5�40ivd�Q=Q��.ȡ+�d_�=6D-ܰԼ�B.k{��&�c�]�b����X��)�n\A49��kʘ:Y<,���|NLj��n�T��i�{�i��]t�z� #+%��*�����\T:�Q^���6��n���y���tq��q��	�RF�L����S+6ո�0�W��t���:��l�|>��]����J#=U��O�zG���;o�d����_5a��4�d���p���7)��wVshU��cmk7�X��K��������͉��{U�b\J���{���fk���B�2�tW���,y�_Rw�����klR��J	%�ֹѬ�'\*�������4���̍����.6WY�I���6��]vի�)��#��%L��V�	\���s�ƛ���T�����5&G/C��W�*�w���gh^��)E����jc[���4�M�����ns�`�
��x+�������K	�d|�=�ޫ}�i㶪�F�f�G�x`�DP�F� �u+1j7y���v���[�%wi��g�֪J��f�nǐJ�u�\'g<��e�*�4Cl>J5	��x&;X�]��V�-%�]�x�:V駕Ǧ�9A��N9�WG�P�Lue���AZ�j���K�J7��VHcQ�W�h=����<�n}����T������n�_K=6�k�0����E�n^�YQ�[��	ZF�N��2���-��ޑ�S����{����Vet1� ���5K���6���a�/@us�wp�W����r��&P����a���ޒ62��,}��G�+X�����d�Ճ$�}�9>�ڶ) ʼMT�+9NR�d��41�(S�Ƶk�kHbb�v�1Η�YS��s��mZkhj���ˏ��T�#�"aD�V �ճ�%5U�n�͵��ݼ:�f�J���)UT��`N�;�&�t2��=yW�8�c��K/�5�%ڙO/�`;�D���R5�n��QݛV��2�{"غ��|������R�u_��f��]��m�,:�ob�2h�'��u�Z]3�pk��5��v$�s�L�e��􁯣�w-���Ѷݬ�xv�+��ui击�)�;E�1�ʴm�'!h��N���p�,E��������i���k-z���S��Kj�)IL�j���v8�^t�|�V\���n��XF�� �^�����vޡ�q�N�k2�r�v�Ȗ9H�c���o^f���6�>:"�]����]����Z(up\ᩖ�$3,�[r�H%�w�����/c��z6X��Ȳb�&�
����n��L� ά�(A]�}�w7W˻Tʂyyr"�(<�)*�Ȭ�VN��]�I�G�ru��m������i޴:��!VlgvI�����\�+���\͹�S�.�ʏ\>�ڼj�.-�yt�.�ܡ�ܡ)��`;�(V��i�-�hj�i��(���T���� �)b�b�K��V�0 ]Vk�af�����=��
�Z�c�v#�0V�6���b�B	�9Y��
��,�j�mK���ʤ!q�\��m�܊bf���q<�or��t�\�[��Q���fJ��P��v�k�j<�7q���r��id�H��y�I[�N���EVΝ��/U��s���x��+z��s>��]kVE�+���F��;�Iy%��
G�&�_��.R��[��gF7�,WD�-�AnV:Be+ZkpM���s�ַx�&Wmq�wz7�f��R4G�P��L�H6iP%1&���dI H�I�'wH�R�$H�BI��$
��%�h"�M�(��@�"BT�����R��BIݸ�6�LA�$�hXBAI�Q�D�c��1�1���Lcc2�FD�D���I�&&))�"Q��4���I� Ņ(�urƒ ��$B0Q�����)4̉3��b�BF�2Lh�R.�4�扄��3�����R"�)@� �,0��n\ ���qJP�"˻��n�H�E��+��I�*	#!�E����"}@UT| U@\�V��fx���օ���TUg�s���m�����K���&m`Ч�`�Q�M���1b��,��̝ҭ.����M\�P���
���4{*zm���"ƛ�[�������ixS����v/�6���0$.�s�9q��
��*B/�����s���R��cɘ=*6�C�� ���}�q�����{�é���۽��$8��Ql7~znnv:�o�p�����*!���o��E�Nt=]4�{j�n����j��,��х��>��|���B2g��+7]�xI��e}� ]$h:a���X��8�&�M�����C�Ӂ9�zBm�y_5��^i|DݓS�֙z�"��t�s�:�ǅ]��utqN� ��ڎ��<1�irf��~鑐)7Bu̳1�L�kʧʣd��}5֨8�F\18�0�*�{�0+e�I--B�'��m�P�TYbc%8�R�N��G J������������up��{��Ϊ�[�S�u�����8q�}�%L���q��`dD�:��'k�f��f<̮Μ�B�oR;BLh{�yR��n�p(j{n15W&�QA�q^{�8 ������Ty=�y�a�<:K�#���L��-�_�v�!��أۗoS2F���b�������'9}c��5��lǗ0汣�6�2����ޤb���=��&���j��vP����j��1G��,�w{c�V�d[}��hȣ���U�+ftE�S���x{�׸"�n[�̒{�A���q�+�tΗ���#!ٸ~	;�:��9,5į3M
���u�}eIg:�����W]K��~��#r��i:{�S=���T���2����e"�{-٢�~�C�Qg8�U���f�yV9G�GG��}J �S�W���$�ǽ;��8��:J���8�75���{yS����̠d(� >*(U�a9a#�wo$��ɵ�&�%��#�$N�3I;�y/x�����Z���kL���O����POdKSs����)x�^/����U�YH���u)�yN�.�nzq��#B�k�>`���}��0����0\��Ƅl!��.����4��˯d�x�^��o�7���˼�=�[;Pd֌��Z���K�xG�������9椲��
��Ȫ�u6/����Yq�ɴz��Ӱ C�O ���Pb�?O��~����6-�A~�`���lк7.�i�1�_�3�R��O���$:�}�4�*�ّ��VS��J��֒]�i��m�o'L�u]��N�}�����`��8AY։o*����y�Γ�j�I^�cF�nJK6"m�����GV�Y���2��G-5��Z9��V��>��;چ�d�t��L��h5y���ǲ�T5s�N�u���x{��|Vra�ٹ����c�Jj�~f����t��z�-2���q��@��tP6t+�gM���Ja_ne�P����X1�C�V��D���My�[~x�Mx�����Cs�i��29�Oo�Ǆ�y��Q��H��J�↴hm�T4u�^F�E� #��sx�z�Ǥf׻7�J+h�8OޠFitu|��;5[���\lr}~���̚;{�qN�4:��� ��Qm�����L�����/�^�`�|������O�k�3�}�q�\�^)�*���%�r���l�y"]]�Vr��W�^@ڪ�������{˧����
�s~��&���t�juB�u��uqQ�^T�iD����0�k����6hV,���g�Z���pt�Υ���K�Fs��2,s��Ӏk������҉�b��[ئ4���{|���#5}�Xi,d�	0�"@�J�!"{�@��IN��{][z��@t�.{xc	D���Cp��.��[>~o�z���^��x��jy�����g�k ��f��&&9�9�����3z�/K�z0;��߱�n�۬��}�Ad�f�nvWc��Bo,1N�ڝ΀�5�#��%�Ȅ��a��]`4A�DF�n\���"4$��p�y��|)�j=ǥ��4��9�f��N��.�n7�\��ީ�34woB��C6�:��{���kyQ� �I��~��6�M]Q:9�KF��U�*�Eyk�-�.	��8��k��fud�%	����_�JE`���`�� qأ���A�Ep�|+��-{�u6���p���Oe�֎V��}n=a�:Q��Gkͫ��3�P:'�Y'�����LG�޷�ۛ0�L㣁^梺�@�*�z:Y)�^�"4�?�_i�ڈ�x`0�z�e�T>�͂Z�Ey���\�uf�+���4C Ө��!�k=
��C�~��t_��>;�N�q6�1��T�ffI�8�˛���ͱ�0k��h�F>���l����Ǘuz���G�@l㝬�f�m������{c�5�v�j| �L��o�R�� �芉���w��,S�M�#�xny�n�w�+WV+��+�z�y���C�C
��o�v˕x ��k4����s{e:}l�Jt���d�i٣a9]�+�/E(�}��.ȩ]C#{_�b�S��y7��RA����Ǉ�:�w��U"9�))@���ы� �D��������-b�'�V��.f�V�{�ɝMI:��$��]�	}}n"�e��<MA����t;��da���h`���J��YMԶ���|8��K_o=�Y�b�(�p��VkA�V�PH$�+��h�Y���Iꃪ���r�-�ip,Uq�� �s�M�����C���H}n�Z՞�ݻ�����\|6}�Hbi
R	@2��8c9V|�{xz�\�C{P֭�3 \_��������j��ޫ�s�Ub�1��鸵�D��'���.�N�f�=>V:;oio�x�%T����
��,��q��{�o!*�H��|\�
�gw?��o��)�Vo��q.�_kK�؅��x�ǄOՂL�^�ڶ	���kh�T.�)�:l�z��f�N�~Ӑt��T]t��\U�����8J	�<�ٚ�-�!�|U��s�y��gP�]a��(.ʔlYcɐ��EF��8{ef�<K�b.�M#=�3���*���w���W��W�>�J,(Dt�!�� ���*�Ko��U�I�����<��W`�b���j]��dc�{F����᡼���R��j������Y>� �$p��"���걚}ˮ&�e�jf�2E�۳6��j>��\8��)%�#�e�A�l�k�TD�u}t�xuԫ�P.�-�Fgu[�og�*���SS$9y��s 5�n���M���5���Q�ɕ����f�B�:=6�ă�)�F��-��k��д���mm4 �z.�E�a�3É���E��*��hV)J��	��îU�@\O:��@�qw����6<�}���x{�=Pܼ�;�}�Q��̌�M��ꙘD�p*�*��'�MGR�ſQ���-��m�}W�|��8g�����m���Q�/���.�����@J��v��Lj�9��ˬ�<�<
S�EX�Ƶs,3�}A%L��f|��VyQ4�8p6�YV���FOOsV�B���c��UZ�ޖ�p��喇.��a 4wǴzhx��H�6�\����E6O�����f�)��+eqh�)���$���QM1c͛�KM֩�V$���b�"l�瘍
�vGE�����9�-��)�W�����Κ��LD�׼ƮT��6�������w�.Xqn	�S.�N�ӣ#�q��f�;��e�n0K����{�2��(��
��>]㚗z$1=�T)�'19<;�aBE�Lؔ��-�zWn�{��wE8�m�UUh�Qͺ�׹N��k�����	��=@YJ)f���b_=�{�2*]#�����z}�г)Ν\C����wY��0V���Z�\:&�!�wL�3\���yh�i�.r�0`��������h]���Z�-@>�vP�cpG�J#�u����V\ް�e��4�h�Y��+*(�Qo��imv�k�>���?xxx	��&�k,�C��`�/�uU�R�io/o,=o�c�N�8�%���;�ͥQP�Dl!�*Rv+�JNjOZ]N�)΄���Ls���-�HLu���#���IJ�w��Gh���{v��{��Y{=\��c:��q���S��t���Ĭ����+v�5��=��9�1>�m$�����<gh9fQ�#����ݷ�<��o���!�Y4'{��ŋ�r}�_Cqj5�����k�̏u�T���hE�b��'��	��WܝkGk×2��i�5�F���
�x��Xu󎙫6�+�D%�G\��&����X�kS֚��sd�)>&-n_(B����w����Y�B���cӚ۶���5d廾��R���c��l3m��yU�ָ�k�3ys].�e��=�6�l��)��7kX�q�����w�f�Xq��K��b�4��uwh�����s-������o����`z�,���<&����<ӓ/4����4�>}7��6CeWf���l��y�J<��˄�G�#7�6��E昖���������j��vz3�ɺ���j_X�Ƶ��:�ǕAU��Q��\F��	�"�]Ko��#��[�P��39�[Nx�x��u�z���Vm�;Q-ΦY�����;��̃��"�t����6}�	�J#�(�%_m���)�-teF!����G2��au]����R�Ө5b5�^��W����[!*�$���07�ߥ��y�/l�z�FϏ1��_�|�����dk�|#�O+����;�UW_�m��%��[��zTF�@�*�{6��[G���8���?+܊���F�m���w�`�K�Y��(lƠ6~=NĮ�o�x݄s����f�uЯN�����i冱�}�-�b)h��v��YF��;gnk�Y�-��`W֞���u��}��lW�3�K�D�ۺ��cej�L�՝����S�P@)lP�\� ��C�ɥ`3z�Ce�c�:s�o4����Pi��2zNp��<�Q�7f�I��B�z�+��xnul��ƊY��Wj�˘��P��g���s$�2���k�_��<��5�ˬ���}c��W��p���1�-�ujw8;3�v��J���Y�G`��S��=�S�و�%����i�+F~�;hOu�����{O*�f��~^�����q�]w�qnX#Ѿ�����V*'ܣg�1�~+\צ�mJ��5шq���Z�r�������I��lk�#�uى�g�kC��ڦ��&��P�mB��M�ݹImX�[Z��N�L#@6�o;�׆'\s����m7�����u �1+0�׻��ch���<��q��WdvI�{�����935rq�FK ��m�Wz���p����.�,�.�^��/E�~�U�L�{��� �������;!�>&/3Qr��x7��.n���6����eYǾn�ETk��l.�mp[Oʍ��&�9�熫(sӪ)���p�ٶՐ��}rh�>cE�(�"���n{Q��r�J�],��������7��"����E}d*���vҶX�����
�]:��z����m�v�t�%�r�[NqN�D��b{�}�@�?r�,z:��}ID��q<��:���9]oV���x�<ԶS@ 䃫�L9�պi��l��	;�ϟ��0t�q_}"���ԵgdܱQS�9W�ik|������ �T�Ꝩ�co/������{��#mTSS�WQX��fh�`'�ﻝ��I`�P�Kzk�z��keVز>۵=[���\UBq�|s�����g�^I��5%~�Y����W�HM��.�I�93Z�C9�7�r��
G{�K�Kb�jk�*E�
W�[�	˓��� ��S�+�7�c;�M�����F� ���U���͡�T�x�$�b9�͞U�|v�\Հ��w�q�qc�z��kIв�	��T�-�W��R�6�k���A>�I'�cZ��^��Ls��b��.c����r<V�_�ڰ7V���߂j�z���:�-��e�Z��!^�}��s,��6��mb���Z{���ń���:�����h���]��-����2�M��Y9�-���n������'mHҞ���j]	o�jz���!`�u{���#�cɨ
̤m���#�ó&�n4K!Clj5Jj��_EOԩ���v[�d¥)��cWL�%��;�b@���\��pɯ�&]�,3b�l�-R5��t`���b$Գ���a;�5����o�����p��w̚��^�ح�,+n.g8�J��sƏ-y�ם�>r��R�\�Օ*�'���a
=���˳�V9��أ�}*T�uzec��;i�!��w9K�%f�V]�|�k#�LN�N���n�Q*�u�Y癴"1���{.���_�M�te<���w�����ٍЏ�fᆻ�<lq0kt5�+t,Ur���aκI���2��-���KN�ָ��SFM��X(��7|(-���Ꮃs'�ά�ث�����2ܺsoE@��&ZK.���mDq꣕'J.���ޅaڏ�ItzO4��iT��I� >�VY��t�c�v9���b;��V޶-�U�F����:�[��T�w��ϔzc���_´�Ty�yY�[�����J�ȥ���@ďKϦ[�u|�RB��!�m��P����/]>�hỦ�n�N퓘y�/�<��{n��on'>����ְ
�h��W�s���8*��3DMk�ZJ�:պ<z��v�՚#�ykK9��R���X2��3��v0gU�u;2�Xu7(<�%�{�Њ�"���V8�-%mB������n�)�B�{(�7��R��:)Be�܁�&�}m��������s�VO��Մ*9���t𫽫��Y2��f���4���ڋt^�%*y�ځ�;�vv�j��-��k�Ae�'��ʻ�O,�
�����,e�.jJ]�]��ѹ�V����Jm��;�184M���
-�[uu�G���S�m�lC}���̣�f�M�+Urwۯ��.>�.䱟k;Su���R�4�ז-Ռ��+8�3jVnҥP*)	fL���J�or��.���SܩQ�ŗ�ߌ�Me�Qw7�dJE�j�n�iu����]���`;�reN.�E��>��[���җ�X��[��fںeʉ������י���^��n��:A$���X�:e�6��w�n�����V��<�1%��ғ5EA�O��K���J��)ե�@U��;pvw�Zo1Y��z_=Z%*ĮG=ui{w���:�F��k����+�u�4dy4�ZE���m�}����;�e7l���,n�3�,Ό�h�[��uv�
����R�#m�k��ӹaBr]�����d���1�س�w}�Y��G�L웪���c(��[�R/e���1�2�lwU���])�R�#����J��Wv]b;�+��Is�!ݗ�n��jl5���$S�)��z7{�}���Xw�ԫ��G�t,��V/*�V�Pt-8)R7�(�\�E����<�Rԗ�� D���#,��d�G$0%3a��ԣ��cb1F�fF1��"�%�"
���DV3��j5$lЋ(5�*(�L�Q�"�Ww`(�b�$kIFьs�#	E�J��"�Ph��1���h�3(������X�H�ň5F��	MDVd$�JL��lh�ݹ3M��T� ��Ő��5p�CPX�+	�D}����Q�,�C�:v��c9i/djJ岕KC��]�֯zGW���i7���J�f�eM��CQ�R��V�5�Z�JG��U}^l��oy�������z��xk���h*�z��
c1`���<cۻ"��E$ϙ���� �y-xrC-��*Sp]���6��z��g9E�:����+�n'�>�A���7��
/�f�����t�ٚ��u�*���{��Sc83&�x�/|d@�9���%b6z�(՚��o�՗{Q�R��8if��뷣}T��.�|;���$��:�*�Z�X��X���~ǱYM�^�d��̺������oz�Tt�P2`��x��9#�{����l_��\D�Yz��p�]_>�ko�am�����*;���Y^�I+{3S���/V�Ø���s���e���}�ٶ�^��=���uj���1l��R	
R���%�l#�X�t6�f�n �lW��r�R��=�XB�������M}y�����C�M+e�;gSoGv���L�Ż�߹&9Y�lհF��qm�8n�P���Y��V��/(u��nV���k��>H�i��ܨh��e���X��w���dk�n�=�ND�t�i�(�\yWK�T3o��V^fk��D��F�;�th�m���CY���S�tk�'�Zow?UWʟ���r"��K�`.��+��nU��,\}�ڍBKB�zk�����4ޞ�=�k�����n��%V��y���թ��3�׵=l6�T��1*��x�ݘ4o3�_�cZ�y�xb}�:b��;u�����~����N��#�F!2ufE�^����L3m��yU��ㅮ��Z��5��F	�Y3����q-p��3UFz������&5��Q�1�R�7CfdѲWL���R9'���������EiN�H����z����6�׽�����s�����Tߨ{/I�'�5ӗ�qn��H�"�(��7%��Ti��fr�t�v�uդbQ.,��l�q����ư��Jno7]nļ�K�)&��c����}YF�z�FϏ9�����'Tٽ���눵B�!]z�}�P�a��6����{l�z�F�@�|�H���IZ��^��������ޢ"¯���0��eo�z��J�����:B�V�
:C���K7 f!`�7�ե�S���t�R�r�1e���Z�"vf��.���I�u��!�ӎ�8{��N�F����LT� 7-��t����\���V����J���7�B�^��%�,��6u�f�+��w��tgvjK��]�sC��>�ƞ+��Kza�zƻ<Fu}AJSRS�~����p|�����O���ؿF�Y���>0����OrԛK(d8���Ú1	�$�S��:�y �Kb�W<�Bίb㜚O����`���MȦފ�d#��)P��S�<�3G�yV6��_�3�Q�W�_�o��8��,�57���4��������f�=K�����*���mje�}F��8�65�G�5ى�"-j숲5gZ�ݭ�Y��f�r������~��զm��w(k�y��
��G@�Av%O�.SO�ZN��e	篰w=�nV;�}c�u��Q�B�vc��^�{H;^�T{��T&�W����N�y�/!\�/3i���ʟY`�Ƃ����)�|�w�%��F��0ߓc���q�vZ�i#��*�4rtL;!�zT3)��=�R�JZ�o@�|�˘�P���k��g�A��J�ūZ�^t�ԧiym��؀简���s�5���_D(b��JF{<��C;�U����c�X��zO}~ѝ�Q�J2�zg�ef1�*�_�L��%��	����^ʆ�o��=(fϗ��Ձ���̀�7��Ia�hZQ��[�䛂�Εٷ���!��\�T8�75;V�9/��+���l�p��Cq�!�m�R���dCύ=Z�;{�	��{ὖ^�WP���+T�ѭ��o/���k�L�N��[��R'�ۗ=�]�C��?��I����K�W�.��������IJ�K���J9`����y��$�jJ�Vu�|hs6��{S��d]]�q�ۀ63�[q��FϤχ�������(\���T@��w�e��l��l�{`���ԓ;�M����S�	P�T.�Vq׊$�
�n[�KsȷX��%�[/��8�8����(��o��1=s�}x�A؃�+C{l����w�z�9�.���Y/z���5'�\䩨\>62j�۝��F�#�ɵYL9�o]#�%Շ��a		�2��H��V%K7�ɹ��r����A��aWm�C�4�b'X�R!m^I�S��aW�:����T^��듻�^����׵����y$����E�T����CW�:�Uoyę���t�ݯG\���'9�X�[Z��	�4-0�Yb*��غ���+�Y�ѻ��g����=�f�y-���|�=��3i������Vw�ͼ�����<��C��k��f#n�,��
�C�_i���e	^����]:�5�o�r{]�}ih��2 ��o��NH�o�v�Wj��1�󐜴���M�v����i�ͯ����ZHz�l��ƶ��b���u�u'������	,wd1�_$͌����}�~΍��b�9[�v`����5�S������Ĺ���	X���n)�7���W!f��UQ�~*ʕ+��޶�Ul�y�'��v��oe`+;�Q�h�;v��V�v$TW�n�)\���m
;�`�z��+ٷ�o������]QDm^Dݾ"'x�Ak�%�Y���}�W8���ҼS6'L{ݪ�V����enߒB�L�I����1�ȢU�K��Z���s�Eմ��W��� �)f����Cl�֊���]Ͳ�J:��X��u�"�W��{δ��Z�Ĺui���5����ݬ۟��Z�ՠ�(����}m����r�6�����
��ʚ����u�շ�˵s(�4�:�>0�^��vѝ^x�S��EB��r�3|HP�}u�M+��Ѯ%�|．uO�I3z����v��f�q��q6�x��!��UB�V�F�-l��縎*��o.���Z>�= t��F'���^�&�MB�h�qӴ�ǱM};ە��kGhr�N(��L�s����94"rs!?#�U��U"gܣD&:�eɮyKylD�H��NL��T�N��箍��kͱ��3�5���G[��كr(ٍ�����7w
���{Z���0�Ѝ��k�t5�H�\ŭ鉥��D��3�6O���Cﳚ߲y�o��������LkY���U*�u�:�7���O���P��}ޠ�}i0cx9Z?)Ո��/Q�޵c�f��B�G��q�jX��<+�y�vo��|��{޼�)�
cz�ȳk�y��S�A̍��h���qu��{���vRw��ۘ�n�ςwۇ�9B���qve՛��Fq�\�GZЁC�eޥo|VQ3����.��W�^��Z�R[�Wώ݄Fr����F��7���Խֲ�7�y���:��v��C����#�,�*�����6/��+;q�ҴL���-�fw-|��;�8�Uȃ�Y�A���ی�n�:[�=����f�ᅉ��m��1���{g+Ԣ6A�0uP���
��:�����Й�"ߛ�[�0հn�w�Ǣ*޻yC�Xp�#Ƅ�}��{���ثlq���օ޸����Ol�U����s���}��.ceVh�hH�owT����^.������>���+���o��
�Qg��볇\Tl��)�@�Kb�o5�:�'ƀ-��6�$;#�H��;�q��D$�PR̄aH�����(F�x�b�F�J�)���1F7��ƹyT*n�+�!�	%���D�F��f�w�3zhھ��ݹ:о��Dܭ~K�i>f�}���,�R;Py�u�S�����\�S�¬cqV7{6�R�11ѽ���RLvRo{8�[T�F���<6��@Ȭ��������R��>��"[O#��W�^(��\ s�qm�	u�� 1˺�V�@�$�G.�0u����v���WY�LGb�Q̡9t.j+GVg>`Ku�S,����JKj�s��t�49'A65ߑ�>����i�����nw{5�9�J���72��{V7V׵V+�'F�0�6�m{�T�:�m��e��ܞM�3TL0�:}�^��R�(O-}�����mK���=��^�N#�Ӵ��=Jŉ�z�r���g��.��V�)�/;��Rgپo�0ZZϺ�6ƻO���۟ߋu��kX���b�T�����j9F�����4���!�<�f�^��s)��K�ɬ��6�ig�-s�.��`3.��MoT�F�:7_���0��p����gD�y�<����L�����z5��5�������	X�t�-��n�6�X�Ϭۭw�Hz��f2���rE�+��p͔�Gu������ϧ�<�n텝��e��<�D�7�ؽ��.��3iTT9�(��P"*��]uC�)i����d�k�ˡ���9;E`�\�g�%�#�8X(u�j��on���R��'*6���k��lt���α���!�u�[j��q��*��ӳ��
�U˕c. z���+��K~㧓q������b��/��M�v��!9N�ƌ��4բ]��o�����a)�Vs�7*-h�t�W��G}����U��*�On���*�F$���!z��Q�#
G{�|\B[�,$(�b�aW��>��H�����K�m�ҶoR���Sl� ��H�=���O'��
:���dY�d��-�㚗5l��l�a�#�B�w]��c3x�@�Z�wG7�2��MM���O�}E$�c]�nT��Mp�����^�*���:#ؐS�g��}�����Dt�x����XOF��k�9�LZڌ��/2�9�*s�t;/l�4����r����y��зL���s�z�E���Fݝ�c+�*�7Z�9u�ьM׷)8E��ֹ��x��7�.�r��t�q���j��B��S�*���/��H�i�*Sq��u�Y��*�3#�[�]FZ�F�Q�Ȕ�N�iؤ�֙Qڻf��^���!� �tD#&�N��I����M�0X~��my	=�c����]b�=Rq��ŌZ3ûi8�!7*_dYN:��@�ᠻ�Vp͑ ���_a۠uYR�J�<��;��j-tՆ{9��\�����立�j�6��r��"5�g0IA�B�䙹�HZ������Dﳣ6v�;v*s��1�g����݅B3���P�A+����an�y�E(G��K&x,�`gu�m�y{��~�w�>ӝC��9��p���T����b�����������W����F�@�#	;o5��y�x��\����ȶ%m���������[`�U���>�;�V
�YpGAIW>*����5�kk�[�@��~K�}���)TT+=�N>���Q��W9�����-��K0s�b}��N+;o�(<ggAusҒ�{��rd�����Ϧ6	�us�G.9���p�%�=�~��a�%����OEhϑg�
T#`��h	��V;��h���=+Wp(�\�S�0l��P�2Ƶ�{ܭ�U���89�߰�=�Q��Q4S�Ps�i���S�ǅ�-�$Ƨ����<����+V �Wp恃a[c��W\�72;�Զ�s��Q�ucI:K��\�J�3C����:U�^�w|���Y5���t{5��*Z@�N@���lڹE�*���$�_�a,&��n��]�%���bT��e
���3��w*��@�T긺���	�l��i�{%E2.(���B��u���J���F�������|vW)}�1�;G7;4�q�D=�;jl5��q;UN�-�N-�8��.n������[����P#���e�u53�k;��f�=R�6��F����auwD��|�;&�o=�"Z�M�pXM3�,WF����[�&�w�q��pu|�,A���U�̡�Qֻs�i��c��J̵������b���/�8_<p��  U���I���h�RZ���% ��Ըq�컮��e�R=5z�p�;���%���}����Pj[Z���Ͱ�o
����%�F�j�z�ol��X,��8��7W�e܉W%�zI�Q�6)���p+N�=qY�&ͮ	���m��D//V�JVɲ�g�̃��w�.aDWvpǡGʭk
���d��:2��Js�;摶sz%�;�Yx��OJ}d��VR@�*��Xl��k]k�%�-5i��2�+ko��u�ٝ�X�.i,b�V�0e>wE�g����eΧ� 8��fܗG�=&|w�lm��;�04��(C���;�і^�Y�Y�����6�v?C[��y�1�VŜ �x�MgWY;�g����̱��,D�pl]0���o�����5�ltfd,��|���c�_F�+72�U�Mӎ]@������L�"	}�º��r�ۮ�Q̛} �7:��=���2��t;(3��lW]����7E�u�d�3~ok�q5�[���"tՋ�E��\y�3Z�h�wm�1�N�M�Xf�we]ܾ�2�O��x�Z8�*�u����7���1qL�Y�E�BF�2yc�b�����;��>wf@t�W�ޒ�O����0�@Y��d�#�N�!N�n���B�:�B�#n�ot�G��٭�nZ@�X�����j,E�ŕX$,V��C����>H��4�)1E�tWK%�J����w��T�w(�̺�wl�`��7+�ġ��iM9�mS =�F�.�l��c4ih�F����WH!W�V���+6A����L�q�}��q�:�$8`9�Y�
C�c��ioG�]N��vz�� R�Cm)Y�7�H�]o��N�q+ uZ�v�Q�HU�V{=\��d�7��lsT�	�m/�:ӭsU�nN��v����]���㝡B"X*���>j��e]`�T����K��i�9�K �Z��}��M�U_�.ڳ�hG|]yz���hb`d�� �jFIu��%v*
�Č3o�e+��k+���f�+*r��	u� `"� +��Q&��%�i4TIb�Q�m�m����DF�*���wj�ۦ�K\�m���:�&5E�6�<��Q��;����� ����Rm��Z�����U㕯��EDh�TJ6ѴF��*-��4lmb��1͵�A1X�W1�4�I\���ۥEnr�ۦ�V�r�X�rەx�^9Qb������>�t�#��o3L��w���Gp��.��o����#��^WƱ&Є���m�U�Nๅ���\��1ZJ�S/\+s����9Ou�;�Kk���MQ���M��h�V�1<���kj����|D��q�t����U~�[Z���ba���#i��vk���(�1�+�n�=o5�WWUԂ�Ĭ��c4n�[��ڗ�&5��:�<���g�Vz��533WGљE)�f3ow�VF_���i�R��N��������ĝ��(b^����H3�Js��ꛜ�%8�4�&5�5V�OM�|��&_��������Q��WÎUXޡ.z��wD�sw�'f�k��Ud�zuBi�t�?K��y�{g*�FϏ9����iѷ����F�q��=�9���B�.��ZW,�7��v��8P�Z�-��s��g.���["��=Ȯo��Y��MOEh@��ـ�s��fj�\�S��#tH���u�U)a�Zymc\�/{�������c�eLM.�[d	G��p���q�y2��	[� �3#�*�:̘M��V��]�j�΍el�n���'���_h�M b�^�b�\�܋6����r�M����FT��O`��O��Er��v�3��W���	X�S��V5g| 毻K���ϔ���@B[�fBΡ���s��
vO�>`���K�!�<g(9F@F���qE-��������`��.\��[	<L�oy[7��܆�ِ�.��ذ
}0����f߶��ֳ��,���*{ѭs<}��+��GpA�x̗�R������J>�6���������K�����a5ٌۑ�Vn x7	D\�?��s�2�8���um��X��д�-�:�(=w�9=\;�P���g/���^����y-����mM�K�L��"Ve�S�豦�wA��SH+���KK���V���W���T��y�\�1Y��r^E�޵��GW�|������߇�}�nA�Ζ����9p�w5f�vz9���O�
��`�q�{�3�m-!OY(q���[�|�^�խ��g��� E��>��E��ҼB�"�!�N��nm`��I�x�u#70(c��7�� ��Q�6PO��&�g-ӕ����N���P�zNL��ݑ��%kU���^j)u�Re�呞��w]Ʒ����]v]v.8�%g#ir�%�*v��u�C�aN(rMٯo��gF�y���Ω-�����&����`��Vԕ�'PHk�p�0����/�(��
������QF�h��J�U'�첵Z�5��c�e���L�Nbrh-j]@����[`�k�1��xG��=����OX�]�f���_ER)�k��\*W϶�amZ�ꎞ�6c~Z;��2wu�
GZ��8����Tŝ����@��`3o�<���*!p�wH�Nݩsְ;������g��I���]#4;���f�,�;�M����#��ۗ�*|�y�����۲���1g>R����R�>��8�8���ֈ��]%������T�I\p���e�X���r�7yb�9m�Aa��+h��]�U�o3��xh�~��9ى�dA[P���9�n������hޏ����I�%�����Uڶ6��n���dF�Bs#�38[�7�\���fYJH�}kٵz�]�ހYGa�>ٮ�+ǼK9h4�M�G���]�۳k�� �ܮ��1�ʽC�4l�o!��ڱN�0N����ۮr�ۛs�4�_�lkQs�����#/�^eb��ko5'�*=��)�=Zw��K1���f��;~oj�9�����[���=q,��q��#�Ľ���g���07)8E���u��B�7CTf1缫 D�?I��×=|���'\e��'-�eJn��u�c^�{�E�(�=ΰzuG*����j�����F�A��_$͉I��M�r����n�Vm�R����y�,�^���7GQ��~����[�r�z�f.K��Q��*{,h&)�Aϗ��d,분�X�B�Nt��r��w�����s��hc凭�i� oz�Tt��B��:�t��IA�+:��7�R��Ύ����ak�Y��U#��b�5ԑ���k�ڵ�w4?C�4#�v�;��Ɓo�+kS�Π�e*�֍�Ꜹ˕GzF7��P���6�h�Cn��MN�ꭨ�����#�c�u=]A�z\yAJ~�,=�W��Y����L˾��S��ْ�A�%R�ҡB�����^���s\/+T�tv�zCB~^��T�$�j�ea�#��F���:���e�Ԃ��Go���"ء�fs��ҶoV���2wV��I�oaǪ�5ǎ��#~]# Փs��8_o�NW&�eu]1�%F�slA���9�A%�P���=� �Ss��[��F��G��z�V�<�&�9�CL��A�]�T�u}��\7�e�9��!�(�V��i��=u�q���MIW�%�ƻ������U�~�'&z�=w�r�^����Fp4}X��?7��tuؘf��yT5�GI�[�ڊX֒����z��\Sm&"*�s��n�@nV;j_X�Ƶ�cGIS3�A��S5�{���Z����j3(�3	��%de�!���/b��Nq��uC��*cb��u�z��h���\��BnP���T�S͛�4�O�R��R�}{��)���g�C^�8jy�o}qm9a�	s��/n���DM�9q�YZ����+�*��\6�<̾b���c�EʷN��sB0�����,��oB�1�Q�j2�eRΟ]����cS�G}zf����S��6�!���[\�9�Sz���ܜ.��O��r��ξ��f$&��9�=InvT4S�[�u7��;�YIM�
���o]{ӫ=>S!o��o(Ob����?<�щ�].��-�lڞ�~�����k�cKq^��m��i����{���=���vv�,�m����P"-�I]Bv��Ou�&��CYoa�6��U��C�F!\�ճ��ߗLv���ۢ��wz:躖��-<����K�A6����u,,h���ޜ�)hL+�y�P"��s�ir�K� ��}��&���=�[j��z�=���<�dW?���m@�J�3O���3)��)�̜6����V��X܊m�p#
zR��ȁ)J&�8���7�-�W�X��ۜS��A�t}��8W�R:��ov��w��u���wzM���5��I��&ž೹�(�ٍ���L����m��χ4�b�z~me)����ѧ�\%�O����L�7���O���u�+T�^��gsF"�{R=s��M�X�䵁-�U�����)��ԳήT�tᳪ���\c�fT�%,nS����W����m�.Խu�Vxoy٫4��/#��X��n���D<�rq��m)}�v5Bt���ܖ�O!s�/�������9�Z������yX#+.��o�L'y�Z}<��Ey�R�}fvե��e	��/}��ʛ��7�Fԋ�[ª����\�/x�t6��T*�u����@~��v��:F�qW1=�廵'm9;�^�H�I�)�R������i	���I�z`����.]$U�u<�Н���;����$�/M��Wn�iL�U�ֆT�����)֎C���)mNtwX�ڳ�;�ױ�.�"�:��״�x�]�f�Gm��>;ʁ�t������ϥ��K���	l�U)�%������M=�oxLw(����c�����W=.S��\���Y�kVXNװ��o�J[����
9��wh�y<޵V����g\����?&3��8��B���ˎ|
�FY��$:[��!���[ �{�ne���A봚��{�w��g���-\�����+ $��ܨ�(�4
�.�/���t��|��ŗqZ�М�v� &k]}׬�==��Y��	�̙uu��i\-[����ed�[���˶�SI�j�7����r���>y���}
�a!P�V��h��T*Xm������p��8g(3C[�f&��a�*8�zU}\����N��<����M�:ѫ�Nn^�"rs!0��V�>U\��bz����m<�Ҝ��7��Ō�=���E��N�窍mm�v��?x�V�o�ny$�̬����ȶ��W�~k��.��w������m�a�����x���o��m�^�i1Np�s��J�<�3}��䶋��ֵ�oc�
h�7�j��!j]Z��3f`�H���*JQ���$e��j,7��'Y�%KlM�C���:�V&}�]N���݂GGb��V�{lud��7{��5�اo[U�ѳSR��sv�M���Vv�S��
�uK��N�j��f��ÈU��]��⹸$r��c&��~̗7��NT���3xshLt1b�b����۬O��DZ��I���m�������{�u"]���!mծ�ɑ%��l��t�<WK����]pHaŧW#6�f�����H�mj�:�v0���u�;l�R���`A�O�pP$�u=~~S�C�Jw��R�&y��R�-ж�m��i����2�]��]Se���-@�����u-�G�V1;Q���[����!e����Vs�>V��!>�w��"�տE���]~�N�oM�ZX�c�Π��Z� �ي
&���p7�#������[��k1������F���3�ה#�<�U��\	�p/�G8��6s�����	���U�M�t=xY�ʛ��yT*n�;S�8���]�>F6D�g��˲$����y�E��}m\��ܸ�'��o��x�#�J�Q���0N^�w�(�J�x{��8$�T�t����kͱ�E�(�1Z��P��'ܲ�iV�O�n�	��_�V�Z���E�#47��7�%�#F��0��)��d� �n��<�!.�.���=sۻJ`Q�Y�:Yb#aɷ��@1S����ܫS�5��&��%fo�U��
��W�\|y��n�9ђ�7uy�V��"c���V'н����F��Ǽm��j��ǅ�!�С��RVF+�p.�X3tUr����^y����S��X�}x�j����{[)q�o�A�ȶetѫΌ��Eڡ6��'�2�s�e����W���ꖞV�!�x=Y��3�;��L��.��{���=m���C������7�b5����n0K�����<��ˌ�q�@r�w��v:���[|��y�\�F�!h�c
^Pi7n��V��Y״s�2/�8+��q�]w����-:[����	��+����a������e��nҳ�����Z�L��2��'O�uW��P����89��a�A�=r��-��\d�����b��c�oDl��"F4�t]xKzh��0M�hF�Ko��Z�!'&�?s��y�+�R���=���s���b�x����������Uf�/[qO�;�3��(�F���펪�����T=�G���Ɠ����6��gl�F�l��)�yɲlO���	;�֍� G+9u��o��8K���4˾Eî���ǀ"��m3���4�|�.�9��)��],L�z�oN��=Me��kiϜ\z�u�wDn�N��L�ҡY/�/yT/��Kv+�3�\�I�)��!��;K�S���@��'X���ܤ�FF��3Z[*�!אJ� 4:�_u$�M�wta	�b>�Hd΢����ϰk5��j����h
AC.]1�g]�\RB�	��]}V;V�C�TV��<��J���[xv��u�ħ�`���r��vt�u�(�0J��x�:�Bt�Kjb���2�W���C���Vj5��u���|yQߐ��4�
o�$��tr]g���%���ZV�s�"Ғ�St����ޕt"v:1U��Cta��sC7n�8.���VL�n���5ܷ46�r��kN�]�
H��W�Df�	Q�J�1(����,v�0#;�RW��Ŕm�=�t����_	�!�-���i0^����j�.�(΅���Y�`a�6���<0Xs2�c�p�W�e���[�kE1@���.�[�)�J�K�@0��ܷ`]��4p��ώo3+��j+30
�:V,C�C�hwx5u���H�ʹzE��9@q�g=�/��
�^�p�V�>7�vT廗1s.���}"Ve[��Q��˥p��m.��J��XFX�'cu2h�6i��BV"�奙e>]ĝ��]���v&��b�;� V��*в��bС�T�;S
=d���{Z�I]���2Bb}S�KlK@O�ګ�<Ub�M��\3������aT<e\�`�;\�ko����t�$����C�ޓ���HG�u��$J|�h{}X�ۼp�P�2�GY3��ά��S�K�FYcz(��`q�#��ӻ�2�YƟ�vk|��w�s\0L������U�:h��ׇ����bV��Bv�f�Y��p�0��M+
�Ku��%*�Am�Ƃ�y����5���x�5jf�����]���WM�]���h.PLFt'�,Y�wE㕵�8ugTz��r��EvC}�9�����-o^��ub�x��u��J��`���m�ܮ�t�VR�l9��d����Vb͊�ŦN\x���97=f��):�v
��}���t)1�<`c:�ޒbM -��N�`��1��q��iͥO�98�F��D�\o_h�36�-�v&'��=�h�q9N�LܼI޼t��5r�'���N�@fIV[v�lFg`o��9)�»/�,��d&n�;7:��=N����Asz;	�ܧ�kOUؔ\��,�iQu�(�邩49��
|]�gu�4W`5��;I����}ع�]�[-�`�p�K�{����1�<3/�F;(R�8�xsm.�`��5kS׉�]� Qm�՘�ݾ�][$ͱR^��[»�+�� Ǝ��Y�Z����jl�p��=v7���g{ڽ�5��j*5�&*y��ot�*,h���*�lTm�nU���4[cQ�Ҩ�bѴh��cWM�5�Y�\�Pk��5�Z���76��kr��A�ب�%x��6ƍsQT��h�6���ʍ��᫐m\�諻����^-��gv7,j5��cW.k��͝���y����qFwQ˥��\�W+sm͎��g����=��w�%�N��KRG���v�ݸ�}������[�@+�W��Q�cyd0��p�r�':�$��ϣws
�����s�j7�9�~]��mN�q��/�}��6�]�(Ғ��g�4����O7��Y��a��ո8�Oz6�\�6���v1J�&r���v7,G�Ћ�:"��ܞ�4����:�t�Q�rlcBJ�<2.��9LVݘ�-��������O=?6��<����o5��3J�q[�҅Q�cK	��o*���t��J/�����9��-�nw9�g�⌝k��f���YU�ѳʣ/��:+ԝy�U�F�sׁ���jE�Fo$����ya��f����ͧH�p�����b�V�.����Z���%ʡ%��Co�p�n���7�C^nMɳ�=Ѻ���HHi�m�]�b`��[U*r�P}~���I��7֫�M��~r{sR|NI}�l�7��Z��>��S���	_�g�YJ%d˘c�Wdnnݡ�TYV��g�a`��`�k��śq__�A+�x�<i���c���*��٨訮k�k���r���2±9���H�]dh��8�-����n$P�WЪv�c��d�&R���}xgwۧ�#�e�Q��q����C�(S[��ٽ��3.#$�A�t����Ý}�ς0v����o=�ݴ��U�85��p��[�#�A� a�T���.*Ge�-��ȷ=�!��چ���ڷ�ART"����AC��ս�XV�ױf?j��Ox�~��HT��BS�@��V�S�3��
�]3�ݕR���;�q!W5�񁽺*v�����s�SI�j�7��:���"�6�L��Ԗ8��|64�f��\�p�<��_;�c���}�����\[Z�!�vk��3���F�\��nU��ʣ�@-��3�w{g5
�l��P�5�����`�w�w%nP7�)eNSW��Vv��i,�R��_gXMQ�����hκ1cF���w�:eh�
��4�#{t�$�Ք���s�10�n6���f����m�S5Ha�%�[2�賓�76�(J�g���mI7��;MV��H��4vؚĕ�;W�o���r.��OZ�ݶ�7V2oG�GLŜ�/n�+�|�ba�+����Z�M�U���W�4t���SVj�����mG#��I9��n)'t��N��U���NBs������Խ�cZ����c��O+rS}#��U�Nɫ���v�R�Fd�YBO8��O��v
�����*�[.%f��ö���B�1�-ǓG�UB���Ss��z+�tgu��2�2b��xX6L���O�o��Vv�N:aT�AΡ.v����p����|�YS�i�����m����{(���F��0ROfMW�gt�ݬ)wu�s5�B���n������->�{#�:}�#FD��{&ʪy����W����+�[���<��$ѵN7�CT�Po�ߍ��+L]��sox�(��\Y�U�ܝ�tTgw_�ӯ��-<��5��3��62oLU
���(7�n�[�ꊎ��t�����j�9��O�o��.�ٵ�iJW�]��|;�'&ky�϶3����H�wL8�{`��W3�r�^s��G]{Od��A\�X�z*��.�45Y8�f+j���[h��6	�����:?X�^3Y�i�SȦ6��U�ͭ��,h���$���>[�i/iNu��X�MU�7;5st�(ū{k�^��\9*�+77�T=,'ͅ���f���O&����F;�N�*�wZ8���	/F+Fx��v�dG7;�eSF*�ZO17�f�gb[���3M�����pJ�9FϠ��/�(f�����oR7#�}�G��{CSi����&�c]��vb���ko�D��G~���=nM�p2w��~�[^�X�s֘E�#,EU�s����]Q.��6�g"=^��7��[�E��<��ڗ׈�kj�E�9n���tX�k�c���e�	�C|�IΔ��$�Tdz���^1�JR�ݏ�y߼y����'3F��ioÎU��A�0�@Ui���̳˗5�5;]��	����M�K������l����+�\.�x�ڈ�Iet��v�����|0�Յ8��n�7ל�<�z_:�BV��f^�|�3W�:������PZ�W���a�m�^^�w���t^�0j\����U�T��qU�E�����*�c�ݳyr�巀#����;��ʒ���xskc'FfY���0�)�n�����N�·+��n��R�����ȵ����`6�=P�ӆ6��u5M�O���z��-MO/V��K+ ��b)���_�6Z_�O÷�;��k���m彆��D�:��Z��Rr�|��dB�{�f��*:G(��
*�줰R�e�6f�Z�/-ݝS[�b�T.���v_�eB��q��Cw壣r3���}�ϥ���[&����h�s�}����9FQ������H1:j(�̻An��0!�Y���Cv�)�a�Ԝe�l��2�Wn�#M\߷��P�C@�齥�=�*�f���\���g+��D�+�42vXಫ{y�����GOT�6�sSk������t�Q�I�:�U@�Fx__`���Tdh�h��s��q� ���n^Nsڿn��jz�;�&Յܯ�k�w14w��c]��UxbG8�ksї�����5�wn�q?�Wb���:�~�SS��ͫ�W���/�+��1�Bv�w��XC�t��Zw�.��)ڂ�q�h��������KO8��5ɛ��*f�D��cľ��K"�s;�u�	k�����O�Go���	�n���PHn����%���4�qhU����,�h�szM=:��G��Y�Y���0N��fY�vgovk��y�m����j�g�����ߛ�)�^�C���9�ݥ˻�*����[�79@I�y�e��j�]m�m��R�8�����
b��܋���ʄ���_��7˙�I�r�:孡�^�����ū���/���7���Ts^Z�uwA�]C��i��ekPX�7}�ZH�y�7��g(R����o�ŝC�x�xXu~��4�Lwk�U�)1�/o/}~����Q�9Dl!B$�mJ�A�ا��R[�����y��΍jOl>����[B��hov�����g�������4a�}dsO�V;[���X�`�3���)^��avLb	V�U��7$G����o5��Y؟d7ܢ�����HM��Ŝ�����l�a��i�fQ�#���� �٭��p#�����M( $GY��b�
4�>g�t_��^mm3}�^�:�]�0��E�Nr��� 7t��gү9_uv1t�Ҧ���|�����w�ۧ���cL]|�Lq�	��K���ۇ��Za�#G^��e_%-G�:��7��LU
��=D�k;[�1C��X:Jֶ+��\�R�c�wwU�ȯ�G6x2�g�%�6!k�����N���a��И���x�jx�a�#A���5�8�lr���녹6"��{������{��C�n�����omԁ�IF+�3�+"s�H��ڞC���$P�8�G�g40����mbo���zi�;��&�[q������fD-r���������x��Lt�u��'��O)�s�in]�c�S�G�:�dk����g���Ot#d"?�Q����Na�/�a*�a\W�麕X{:��<ձ�T�Q���̏A'<�C��vF�>ℳ��ۍL��]e�����2J�x� ;��I71�f���YF�Y})��S��l�%Z;�WΜ��r��/Yek���7�:�OZ���ٛ-�εȿ��
��M�<��u�QO�7}/�i�8.Ԓv�g���Q>尷3r�m�=�To���qS8�/��@����/}��L����lꦮxϴ�q�+�<��2ö#_�f�N��L��=��O��y�7�M�L�T��� ����ו���Ppn���<�1滗�,�U�2�<8��:�n�9�g�su�E�-*�g�%��`|����TkEb|�qxkX���N�e�i�Sq���w�T'r�]>'��O�I�їY��ٻ��� ���`3�J�Go�E���z���σ�3�=���j��Z�� �kq�����U�J-$�2����G'�����%�7�.Zw��e4yz:3F��\�k����GM�����T����qQ�P&
U���efB5��>���x�v|Z�Fo�C6��U[��r��놓p�ԍ�T�ҙ*j8���䉈��A������32�D�UW��f}*'��5m;H�oKe���mށn|��)�W5);$b���;G��f�1��uϟ�J�Ӄq���>5p�[��|K)��%��+�6��qGg��i�'�<�p���-s74\{\�
���4'�{�F�-6���O����4�ѸN\~F� �Œ���r�����ժ&f�ђ[:J����1_J��T��졝��I�и�t�E�/������^��Z��B�`�q�*A��D�L-��c��fⴽ��4^��<����V�}Yy�w�hx\w:��;�:[��깑{(�����̨S�|v�V�e� ����^zA���T'���qf����q�� �-��ڮ{�b��$9��^�T����� L�RM��!�<]zC�lW��pM�7����}�![�$��_����ɩ��X[u�j|�l70l)tأ��׳��J0�4��f����o
���uU��󯭂�^�5Q��}�A��������0<B�����7ެ��
o���_�3�Odʁ^��)�J��:�z!�q���Q��3���';����W��]��������&Pۊ������Dd��
��T�`��}�YMX��:�E���dU}����s�k��t���(z�t�$�9��+�]XX�G}���峳{=�I�y���qtU�7�7.eev��d�=S=��n���w�Gx6�ˬ4�������A����Dv�H<=��tu�.J4�$� �b$��;�M���v��uǴ_�-�kuV��Viĸ����KS��KΙ�UH+��� >��	��=�C���,���Y��7V3��>���n���s>g��G��<w#�g!L��@{̼u}������{ȇJ�=���8���)�F=�m�r!��m���uL�o��=��\.�P��Q*��\�&$��B��U��#,7�Db[LpEmQ>D�U��u-�7��J*Rd�%0�!:��2��S���Ƿ���Kqa�/�%�����κ����@wK"��kT��v�븹3ʝ�7�]����a�����.���hS)�\�R��N�X��0R�6�ݥ��N�5;���.�Ҩ�I܁3\	���m:7^��7���W!���EO���
k�gޮk�NO��9���I��(�e�?-��Ml-y߄*C^����ǳ(�2���Í�Uɸ�7@)�n�_�G*ƿL��,��|�����N�L/qﱯn{���Wg]�����ˎ�BN�' 9+��\%���zf���F��p�@ӎjj*�Dc�����^�O����J�e�S�t���ڸ~�4�ǚqZ��wpz���4�H͑/g�K��PH:+�s�`�xs�[�|w�g�H��gR�<ס��;`�u�������tY�<����vMd��x��0��Y���9�a����^��f� ��i_{��2%'L��W��I�����t���|�wLn�7���;*t�d�o�ax�����j����/!�'���wvz�1Ul��)��r�����h��r�:j$�5z�\Q��q�7�Q���e�L�P�[Uƺx}�2���閥���h�l��'r��wux~���:�8�W�s�ڤt��,:�r��hҎ��4�r���S����V�U�a�]�����sQdY�8_�������YY]�q*ۮ��͙�d�4�$�A�V��v�v]=���c
��.��RԹ�y�׉P�{h�w��m�T����7����d&��o�s&=�a��4��y�;�[�,KYԮ�j�!e���f�d����a���u^0��a|!���`KQ��k���X*(,RYS�S��Y'.=wY�f"�..��U�KfJ�v-�9��'�wY|)Ҧ��������mu��"�^�[�f�����܃H`;*UCV4�i�ͬ����1�;��NGs ]ڲ`��?�ω��F�v�ͨ��[�e�j��p�&Ra�
:�rM5;UP�0i�M���Ћgg39���mfU�D�:	��[t/���oE��f�:�mn���`kÙ״��+��o�����H���itJ�o���z!��q-:�udn��1	�k��Ӄx��/V� ;��@J�]����V>����p;E�qNْ���0w�T��u�o��sg&�#2�Τ�'�z	;��Q߷�ٷ���m�N���b5\�y�P��B�ۼ�� {!��
���v����OtSX��FG���3}��|�e^<�O(ΝjD$h��>붇u�I��ق��Z��\-��f6����P�C���p2�iq�ьd�x	��Y�7��]�Xh���%J�Q��9F������kz�&�J�8������o2�Lq���L'��[���[f��\��y -8TWܮ��d�!F>]�{�������cG7��#�\�F,�z��]*gV�wi��K�Y3x7�r��$]=�؇VTCҕ;]�Ԇ4e��G/&_F���B♺.oX0u�'Ad����Wi+� �;�2Q8Qn�/��Yg3x�r�M#ͬ����ǙiN�BV�1
젆�Õ��[�+��}oo5V �N�!rc��*�/;����|�cxE:&I���*�)�ci�1
fl8\�kz�[j�"򺴾w�^���f�
��.������F�"xhB�JS��!��Έ^���-3{8��� ; �w�{�Ig_�U��k�k#��h���ı��ì��WH�q�B;x��;i���L�J�"&����*92�#���to^^Y���a�9�9S�%[X��5�t �[2�W
���޵r��v����uŌ�Չwmn)K��}W$�� ��/2@H�a���C���7�ݬ�7;��D�Y��2��������Fhyl%[���4��&�ٴ�H���oY���uum�j�T��Uǭ�ܔ�hV���Ngjrb3�*�+�f�){�j�ɇ:f��;�e�����O�j.\�\\� ނ�8p+%��7�N�z�vbƷ�r'�2��FQv�5e�j|�F��M^r5]�1Nt�����ł�Dy@ |
��.��ss\��\��;Ź�.r��*Lkr���':�ع�Ж-�<\�b�\�ۅ�^6׋ъ7M;����mx�(��طxᴚ�k�<wtDk�Ex�#oӭ�����yݯ�%�\�7��<F�v.j���מv�mr��ێ��3�\����*�x�^9;�N�9E�������V�IcXڼj��˕̗+��<x��W(ч]\ر��e�p�y��t�#26-wq�z��?��^��ߞ��z^[.#@ن�Cc��(�� ����NS~�R<ƨ���Jv��=K/�K(c4���{�s������;�L�����(�%V&�+z|�K+O��Gn#Ϯ�H���X�2T���d�9��Q�چ�3�G��1��C�S�\Su�n[�<�;\r5�����F�$�q�ɛ�g8��hd[���:j:��%�@��O�S��:ჾ�ա�>�CUE>�(�+%���gc�hs�����J�i(�*���;Gѷ+��F�U�b�HЫ�1�Ӷ}ٵ[~����m�>��K`�"u�Z�;��S.g��òD�+iѿ��q������m*Yw��w���ԸZ\s�Q��[�m��_��i�5��T�3��D��}�����2���N֎�WM�?
qJ�;g˥鸍O.j�OG��&M�۠5��[������^:�܃���+ܿ�۽�WU�ư���T��m�ٴ����[���bqNM��.ۆ�,���62`|<��7ڣ7\�4�L�h�=1ݟ��^�t��ݤ���<�>�{�N��Yw�KeY���ۜ�7G(HI�j��^eٳ\V����]��6+Ƶo�7*��Fu�Fy�c�|V;�f�_X�	�9�}��s�;�ZK�gm�D�r]��dm�ڥ�*��@s䟎�̱Z%ۺ~�K�p�S;�t~��2[��]ܽ�G��I���D����x���,��{H��ya�:�h���,�^GS�D�I�p_pW{��yǟ%ۓ�Xw��O8���mU���ו���R=aK'v�����Pw�ʭ7S/�V�Yf�ь���J����ۛD9s�I�E*�sͺ�X�j,S�z��Ĩ�]�3����F���3C�$�W���@H�ˀ��M�S̽�w������^���}��-;�~C��q�4��L��3�b�]�k���`��e��r��E5p��>�3V�(q��>c���r33O|f��$pqBOO3�ޢ��IU��N������J91�1�7���OG0.�8���1rY�(���,�E��u1/��h�Zu�^��^'��mP����wD�Iw�>tp��TN�(�p#>Td1u�ƞe{����E�,uq�َR����GU�q%g_}O��u�Ix�Fl:�&�L�5�SQ��h75}Vu�-��cg��{ڽ������j1|f3c����ϴ�r�`6۽�ϙ�I+�A�H�gd
c:n�ݫ���ݫ=s^� �N
q]K����-��ƣn�rm�|K,�2_D#X|��#4Y�ʨ��ez~��k}�����6�e�	:��)��Q�-؋F/��V�Wt�*3c�%A��٨�|��}���7j5ݹ�-�Ҽ7o��yխS�%
�]kR�}gip1��j�642�AE)�j�;�8GZ�V��]�;��+ �ܮv]��B~gW�U2�At�o����~��Zn:!�}w&9�F�Br�k~��]�dS�zv3�cz����7>�i�'�FH]q/-mdmk����q�9��C�;�B���:}�7GV�񎡢�ٗ	΀v�`�q�*A��Y=_L-�9�:\��X^��cG��s6������U�ɮQ��s�Gd����̯F;�:[��Ϻ�R=q����dfL)�zN:\�St1���7s���/�Rٸܵlz]W�N{�CZ����:-\����̙^/5�*=R+|n�s��~��օ��U��Z'��o�����2��Z;ͫ��s��xo�8�u���o{9��p�3��2����Q�qR�>�%݅[�L�S�l�������}�l��UnJ���6a�z�Op(_|�BI|gT�z1�x]0Eǜ:c��ڍ�48:����x5��)��g�c��x�Yd��0��3Ԅ��r��_���ٱ^u���X��e��
�U��+���!�h=>�N���rx�I�3
�}P��٦��\��1K8KY2�$�ʚ��0;������3P wvZ�}vD��r$�dgp%X�i��:���&���C�m���>���Wi�0�i�}�W}� ���6 5]�:���%t���t?�c�u�;�t�ǳ�q��䆗k��T`��,jl�	p�;�Zs����q7)���jKS��{D-7�F\*��d�t�MD��t�>���%;���2��V��<�U���O�&��,�g��r0��R<̣<H<Eeh����o���*�2�z�������l�����.��N�1�s�C��߿mcVxO��T���M�"r�Y��D�
d��uL>���D�I��B��U��|�����	u�����ϗ��\uZ�ٮ:���'Q�:zb}eI��L�;�1R���J���ԃ֪C=.�O������OfV��� ۑ��Ĥ
�e`�߮ _/��P��G��k�����v��:�y�
"n⟞�7��ɧN-���MUɿ'@)�����r�k��9,���|���\��/�M�=n&'*�R��3��])H�9Ҵ�W�;bw|}��O�Ld%��q�dϯ��6���r�M
����뫪�AG	ש������)�����(��i�k+]P=��f�R3�:�03x��v�j
������Y���b��M[8%5��9gR��z*S�
�u���`�fA��K$�9�R���C��9kjK�\=���<�i��R�ۻ��ٮ�����嗍���9a su>}sqW3Z2�����%Ĭ;+t�m�6���@6�m�����M
��ɱ�0�,���o�WGL[��Wm����ݽ��U�����Y��?m������/�T�������@���+�XD����Ebv�3��E�tp�VYU;�ilݮ�].=�w\7O���y�S���'�����B�u\n�P	R��-���_��Qu�hBqǝ���S��ҫBnp>�T���:H�x�T,ǵ��+�k��i�<�┨�k������c���c�O��MS�V���l��'MqcS��j�d�{�ޥ�Sv��{Q�%��]RQT�X�ԭ���,�>{%����o��+d&�q(��w�>�!�$Ӱd��Ut	<�Ɣ�U>fR��[�<�;\r5���OY����/	�%����1���� wa�ȥ�E��js�q����mZ��˦�
�����ױ��>����s��^:����JFJ5�*����m���!�P��1	�������p���P��\�]q/��M��@v�%�v�;$LJ�t[qR�f�~W��{�ѓC����n㑸֍F�.�&�u��C4���`�����N��3)�����������f*ջ��1���[��Wv��{�|(A���fYȜ�@���M�b�z_#�����絘�6q<�G�Źթ�'��u�9dwb۴�9���@�u��q�~��T��VBZDz��[�#�#��l�zv�s���꘺�'3��z[�yKn.�jvt���z���[�~���Y���߹��>:�+��2d��hL��Kuu;�C�ѝ=�y��zxu���늞Â���+.�\.N�v'����.�/w�<�"G����s*<�p��=���ᕁ]KÂ�+�i;�iq�w����şPG���s��z��`�3gu`��;�v|V��<f�W~�د?�o���j3� �O0��v��E���C��{�[����\oﶔX�ʘ�Y9�<d<5���&t�o*��32zǣ�k���Rv�\'@ɫ"�zy)>��G�g�*���wѝ9'h�x{&W�:ޟj��g)��)GV㊞�Ft�ŝ�\atɶ��{��+���7���T{g�pr���e����v�y���%��2�b�U��Z�����y�e��7-������[�0(�rǣ��v9��se�i�F��H;Fx	qB⧫���(�RUbo�N���9C�~�!�^�[�6|ojTgf���6ὸ�م�.O�,��P �*OwO���K����FD�����|�\�+0]N���{et*~���cٔf��wB��~5��[ǝ���h �m���=��7��H������K�������"�ɍSPz���o���]��eY�FD���Wlv�����Žx���ph����f�����u񨺷���h��>;��N�R�W�(�
��Iy��C�v��"FIF���y&�\O��7��IO��D)�>;��p�m�pꐚ�2T�GR"�v{È���8���'\u�?�y��Fq��ƣy:H�3�-���`-��5ϙ��2J�f+;��i��[��r�}A�H�C���W]K��ϸ�f���k�ɸn_Ϝ�2_�F���8��aW�����	�uD�Ξ��3X��,�42������=��D7�;����=��6$MlA�n]؜�9��{��ǡ��&��v�zam���+��N)xo2PŪ��|�+p�`Kt;k9��OEEM:���NXy߅�ו �d�|=0����s�9]+K�M8��צ�=�xep��CG��\��>>��̬u`���_�~���Q9ÿT���/ڔg����ZG�L�ݸݣ$��󧑸�m�`���u��]>�|v�4�Ծ�p3�f9X�w2�L�ױ�ꛖx���FϦp�Tβx��P+������Q>���{�ڸ��s��_G�����3K�F<���Zɴ�GZ�X��E��j�|�^2+�V�w�����H�Wg`�oi�[����/k��T�����r��ǖ�Ű�5׈��\�㳸eGRCr��-v�W�1L\]
��z�
;xH�ܪ�q��2�-��$!T�of)+"�WC����&\|Iӗ<=��.O�}*���L�:�`�)�
�t�Ꜹ��=�(c���:=�,f|�Q�3�l�Z�.2�x�����V���4FL�c=�FH`:S}�K��yꤏz)�ރ>����Y@h0��$��;S�k�6&�D]r�>��;�|n�R��w�ю%����Cۆ���>�q��(���P'���_C�]d��)�5����ťW\�k�;]UL�ʉq-[�������:�e���d�t�I��k��ʩ�(T�:���Ǡ1n��6_�h{�SڇKw�}g���NFx�G��4���:������	C�N���:eTOQ-փce2�`S�oW�Jv��}}���3�g�K�B�����~쎉����T��"jU��d�(j�:<;����.G�0���Y{	w@�Ny�\)��^���r�N#.OB�b{�}_Q�+�oc��w��i����+�=���*N#�x��6���2���n0�GJ'�|p�P�/�t��,|�>�O���eNHsgI|8��}+Z6����7�zXvE�:�[U�#�ϓr�m�yբ ҧ٧.��n����U�=8��z/[~67U���	�w�6�s�S}���N�9����E�纨-rVP��:��r�������sBS���Of5���9݄���?��ƺ	��&����N�R�00�G*��ʐk�OP>Nw�I���¡�i��]�3~~�p�VN�\s�V���Go�;�>��&��奞�iY3�����UǔN[y[򻸛r
#Np2pl�x{+�i:}�������M<1�i�k+>�w�So�[�d��k4�Q�~�,W���rr�Xu'��}G��~'=�H
��^�=�?0n����T蹽�.F�>iՌ�j��W3��'����u�6iP���I��\��]w�E��d?����g�����{\/���A�ݿ��Pgj�N���u���oX��ɯ��b�Q3���a�W�Ցk'R�w,>P�N��+zm�2}�:Z=�ٿ�����C��Ͻ�5}U�G?��3V�@(��w�]<>�!����p�O���7����(�����z�����5ְu�2��uq2��辺(�SBu*x\>��Ӄ��Xϕ���a��FcNt�󈿫�\`�J��&O366R({�WXϩ��7�����k��7��1�f{�2	.m]š].�n%�N�/�3��݆Zp�	���9)��W��c<����,�e�l��Կx'r��yѽ�J��i���3�.�t��ڂ�[��,��9��.��v��:x�/ǹ.w����7oJUr���}�:rx�j;�GcM��檙���}�@� �Kd����w�����W��s����^���~���nD']��<w��Ө�	G�D��0y���ە���-�`��gm�*qݽ�3�q9��#���=]q-���ߛu�\C�S.g�	�쐕���~z6��\��G4��l��Ѩ���[�pۮ�,����ғ5҉ѷ�웮�SK�m���k��8���m`��RGl�;�i��P�5w&��)�L����ЍP�Y�.�f�����}3J�d�1�H�ѱ�Ó�>�Ÿͥ��_�<?������}'�@�oI��h��z|�7ޯQ|^�(����2�+��xp\Er�'}�H;ܻ��O��!L�l�X�|��/�	�k8�t5J�u`���.͟���� ��ew�lW�j��O���r�o���M��D�Q��H������c��ޣ-�3Ϧ���ו���R=t�s.��/��R���)��f$f���"�gx��a� �%D:�J�Q��IN�{|3���ܲxe}�>ľR�0o�b6lvS���?��9����+hɇ��N�7��Y���RD7@	�ټ��\�啽��k�g,ni��WSE'�1����]aݧ�=|ƅY�Nb�8�u���}�s�i�qr�"�����P�ۦl��L$':���G�Y��������8D���~��XMv�A��0�Afʕ�,w>�@��x��"��79����g)��QXkK�{Ͳ,N�۰��/h���`��#U8M����1 ���r�%:��E�
��*m�
�V%�ugK����ek�f���W��ml؞S��Bws�a�ӫ� ᤮s�]o;n����pʥ�s����̻�e�!�Ō���FE��Y�7�=�y2�bm����������rbפ�� v��	�*���M��	u&��,X}����$5�>Zَ7��݊��T����
��5��	��=�/P��3����37��&�YV+�����d�`�i^��/�<�\��эҲ�������8/����-�<ݸeo>�����Oj���	��S��a����]p;�߭��wS�|D��Ka�l�p�ź�»%I����š]�l��3��[C�*���[霗e���u'R;�����3����^�=G)�D+���A����R��gZ��Օ�>��������9�74��t�J�v��Wt��EA�A"�y�u>�)9��N�D[�;5H�d��׶ֲ��7e�'�r�/,�;>oFq�6i>���혒ʭ9���z�"̛�D�J�4����E�U.�� �)�ݻ��Gv�C��^*�M�����\7��r���K1��T���<���h��2���\��8+����g͡�Z�Cնw/6�'{�s�]�^�����r#e��`f)؟&�^���
��)�(#�7�Ul�*X���X�V������"*��2�a;�>�ս/���1�T��et�U.�I=:X��2N��RJ���-&vӵ�4IZ��_:$V'.��'�tm]f����.�:��_m��>�86QW����\�55�J��!_	J�������y`c�Y2�Tx�l�!��jooo5y�u�M�!�2�Ո�R��ܣy��dZ��XC��R��7�M��W�-G׹\����W���E��.��L�i��R��w۝&�Μ���]:���Y�]���6�6Q�(������.㺵�PԧH�r�Q��s�gT��6�eKEW<�G�ە"H��z�q����<_i����i����K��O�G�MG��
�)�����);����XS��_�Z�E��۳`�as:gS�6�j��SR��H:�i9�9w98���@U��8�#T�t�v(�#��:��7�v}�n���;!��.����H-��[�&��]J���wW	l�c��׈�Ix7۠ Udz���ڲc&���ی���~z�߿��������cA���WK�J�3�-ss�ኢ
;����t�r�;\�b�*��nncλx�.sF�lI��W"-r5Æ�nwN�+���h��Ix�$^4;�����Z�6���tɍͷ1�chԄ\ۗ6�2󶹷<^,b��ѷ9f�lQ\�E��WK�v���d�Q�*5:TA�E��b6f����2�$*n���(�
d��ݮA����]�uQ��F,�M6,h���K�4�ۦ��(�7��^7�����x�$w]��U�d
�ۅ#�+�L9��T�4%[��]��t�YgL���[�҄�7�Eu\͡Eɒ�vR�K�uU��� e���H��6Q�p�t�h�/)�$y�O�3_���v��uv��Lz�D����I�?IA�nI.�x*�L�rK錊�@����-X=tx}�g�{'�BT`]�߂��7}����;�#P���7�� �A��T�s>��QF��J�MƧlh�m��q-���l���5 ��y��nW}|�(�x��$�@L@=Ċ9=�>�wQ.7V�3ּ�\�b�eؐ�^����h��>:�:'�*U
�\�j8��%*�u�W��&�F�̭�o:�9Ӝ�Ǵ�O�$��áO��܆놓oH�uHM)����)Ȑ�f���K}�kon��A����qY��g�ƣy:H�3�-����6�@�>fy>�f|�
y���[�+�5>�4��J�U�R�s�2��{£Z�rz!�|K>�3���
����x�}���wF��+�76�q��30����(�42+ʻM�Jµ�	�}w&o��Խa�͝�o�QC}�h�99�5��d����[ُD�����OM�3ik��)��T\I�l���ה��&a5�ާG
���ސ}˵־�vi���vZ�Տ)S��0�Lx�%��xb�``�(c�#��c��U��n���F̼%�t�23�V\��`��Q.�m�;u�_*�u�sR�ppZ�͉���yn���o.�|{��>ݮ��8^�5wB��t�e�sy���5�H:Y=��lNa��9�3�[�7�/u>\j��>�����cZ�|}��fW��7�X����h��l+���o��o������\9�<�)V�u2�>Ζ��m[�US�}��mOv*�;B楟���������YD�g�~���q3�#N��V�R'��e@�sWʦ�,��:�{�WӖ��9O<�W�k�\>z~2��%~�p��&=BgG_�.��J���d���*�7�%I���3�s�S^����tt���|���7|�8�{}S����}peP3�����UTk�
���w0�]g�����nqT�~�u�<�6{�N�>��e��8��&A�C�S=�b�꭮�p�����ߊ���ߩo�C����x1�h�C�!��ݠ��}::���Q�z���9˃.��o'_8]Gke�8�4��E��,�S{q7-[�椵;�B�o:�e���V�ʐ�����Jw�zN�����0̹<�����g�^�V3�����n%��,�g��'#[�r3;�m���Ks��j>�V�]�+�>�#��+>%�Z�u������=�]v�
�9=Nr0�C��䐵�zh��9m�H�M��n0�;�
{�f��[��l�=�f�Z.���s�I��+��+�I���n�S"����A�,�� �:͠MRg'�H�XwR��/���S0x�qU��"~��A�)�3 )�7����S��{�>�H߬/<�������Ύ��N������FF)��I�����}4/�\��#,;��do�'fu��}��z�P��}R��qӪ�>���%x:��Aӡ4�'�D�_X��"��}F�Y-t��n¥N3��'+��a�ڼMKCumH���	*d�}�_�����r}҉�->��Q��{�^��������n���x���p��ڞ�MUɸ�t���`i~G*�Ƽ��Y=5��^�y���������˟q]Y��%�\s��Zor���N:ɿ;�8����w)�t����ˋ�ˆ���Ӫ���N�Ə�������c/��ZN�}�)�m*��*i�|ӊ�S��;��;hzv7Y��xۃ����Fٟ��99q2��ÁdT�����Nz3�Q�k��wY��&~%_	�]���U7o���i�<�����}|����:l"�ݰd<�"~E�+�Xn*��S���$\<�U61hv�W��x�����}�;��z�p�>Ok�w�t�d���axѝ�L�2;�����c7��E7[G�\)<�F�ő�g8t����vu8:u5
c�i9ъh�ȶ2e��+�˚�L�}W���BA륋{��W�Χ�P�t,�6:Z��7���][ɚI]�fi�T���݉�M�r|�[:�xh��^>�BfpK�L��W�=�w��sv�VE��Jw!��k����h���H˹@ ���c�X���I�0�>�~��c$���n��^����C/��}>�j��O�G/���2�c��`B��wI��$��`��<��WS)K�%���z��/�eaOd��� Cv�����a���x����ҠP,������(��φ�EF+�f[�[�+���	��ܤ^g��4��R0����N\:�aX�(���@� 0��O5>_8;я����4����QՅذ�^����!���+ʢp�Sђ�,�N���WXb��p���N{3��n���ᚍW��#E�&�C�\K�3�ۜ_����e��3�F�s�k��~YF��C��h�WJ�����F�n9u�7�n��f�Z�3�t�̵,���)��zF������Zl��TJ��W^����wJ�z�\?Bj�M�O2d�ͺ]�
��*���7���-�iUg��q��&�Ɲ���s�*{	Ŵ��ٴ������'w�5tP���0R/�������:����yR�B�� ����Śsw��,�˽��c���gG��[�WSu��U�@����Z=��=����N����@f�C�qR�a}o�w+܅R��uL{;m<gs��$���b�l����9u�tr�W.�ή���l�	�@;p���K�>7Y=_L.�XԼ8/��ZN�v�~�k�o��x��`���C�m>�z1��`����*7���id���s}YOL��KTdP�1�ouM��+@�T�Gҩޣ-�3���_����E�d�3!���4bLu]��ط����:�n�[%f�q��1�T������ڜ��o��NIػ�j}t���Yv�X9o	��L��0�]U��e@h���+���d�y��-�6W���mB~�T�M\8�X�w�]��rx?������&t+�����R��ѥ���2�و�2-���Ox�Q��g>��g����H:
~�_.�������qIU�������S�N5�}�:b��h}���J9�6���3�a_�����=QP�=Ċ�9=�>:O�{�U���=�׃�VO�O�Wo��q)��沚=���y<'�U*�q�Q�@}Fa@G�=q��L�r�cv-�^��,�h��1�>Oj%�-��3r��s�	p�ԍ�T�ҙ*g��7�G(�[��]�,A'SW7L�Dr����.Yp�A�@�^m`�x�V0�)\}�쨄��Nl�hwM�q���4n޻�Mc@&/�[׫�V��]�WG��Lռ�xK�����[N@��!Q�Q��tgT֌��gp��`l�=$�_�Fq��c7������Kg"�`7��-݅u99��~{�?//fh�J~��$�������1-�
���o�e3p��F��u�6ܾ%��5�@O�6�P�s��F�
�$Wvh��;���R�Y�>S�ow�i�\����s]qo��ߧ�~�j*��&f�E2�c�j2*6_�����n�+��2�S�~ZU���W�u�8��ܺ�]�h�N��:
f�`�����^T����fl	�!�߉�q�H��\+��[��w��S����4^���j����3=�V߿c�t��ϱx�����4��3߷�;�Z)uC��R�u2��9�2����:��I�|�sS���=z�:7����ߎ<�X��ۍh�V�'\t�8r�ex�p,��V9��}2�{��}��')Ρ�NN/
j���[�g�i�o�����-,��#�"^D��k�8%�?r�ɔ^l�n�f��Ό�;e���RM�
��wM��֢݁(geN���K����gJ2��V����_Kx���o�����=��W����ICt�Ҭ��F�����o eh�R��z���T�@] ��΄���ͥ����R�$!�մݢ��<噵����Zҙ{�j̮����,�u�<�}�.ԧc�kzιRS�n�P�ח3�÷{��\�������:c=�t��S��g�b�;}S��N���P��_��&����!:V���=�b��j���\�b;��������{7h=&Ύ�rx�qD��hgIy�nd�m�wݛs�q�}Q뮚h�UPY��\KV�KS��B�q��F_ʩ9K8܂���M�M;&\l�����O�*`����*��}�'�q-�q��=�!9y��F��lz��uC�7d�nk�L�ƺ���)V�����b�ᾈ��#�'зK��^���NL��\t��-��͈uLȥ2Q������DĞ}4/�W3��:�$ׯ��7y�)��,�^����Qng+��d
T�&��*Nؙ�pv�z%m:=9w.sl;".�����t9�l�S�bꐃ���E����,|��P��A��N�!i����q���}~��[�)Wa�Ed��F���j{l&��������KC�C_�A����>�g�eo�$�xo+����u��?puݞ��e��U�~'��1:ɿ;�9�3�%5��}�/v9�(��v<�!��J'[���U*�[wq4��0�:�d7�C4p��#��Y��ǍI���v�@z�z>�l��Fu�`��=Cf�B��Sl��� �y��_ǝxWK/Q�W椲�k�u��)a�fL��Je]i�
"��.z<+���L����Jp2p+�SuԴ�>�ݔ��*�Ҧ��zD�5��)
��:�=4�*�:�~��l�3�qŜ�%��'����p_�=_���@f'�1�S���g׻=�ty��q��R~@�S�G��X��Y�=W3��Q9�d<��.,
ɭ,[õ���2��d�_0<�B5�Ty;�dJN�.�#�)W����\geN���0�f�p3/#vg��f��z��ޭ��S7j�k�j�u�║}��N��0׾�|�D��Wo�FZ�������f��o��I���4e�l���VʀQ����^���C/�u�\E5Lnj�	�P��ʻ��.����R<	:O�uB���R�=}tQ�J�MƥoK�YXf�¨��\�L��g-�#�m��A�V�6� >���$t�3p6R({�3�n�ND���]7^\'u�δf.����v��k���㸜�uH±rQ�� wQ�)l�pvy��n�Y=%��;,�K�罶�Jj��m���i7��q:n:���d�Q`CuČ��n��vG��2����Y�v|�-�����0��f�M��s���
�O{7�m>$����k/k�[y���A�=�p]i��x��WyP�t�c�=�������z���>���CS�Z�5j�!%���C��C+�;��k�)��7׃�����W㜊�&1tb�H�|��<����M�ۭ���ҙs=� ��Z^F׸z��bV���.I�]Fx���ݸL�h�o.�'��\�3L���UR��;��{)�o3r�L���fgx��z|*%m`���s;g��+M�yp�������2x� �ܛ�����h�c�C5B��L���gf�>��Y=���b�5�L�K���~��ZRz_��!0�0È�qJM��.�n�·�6r#K'�ƽ�޻���ó��D�Y�����O(�q�6�k��y:}��bt5�ϵՃ��{�yS��4�ݳ!}Q9�=�,[��
n���]Ӯ����.*v��u�y*c�S�F[�g�Mak��s"�҉�mщ��{<�f�V�Ԩ�#zc&�p�:�ｦ����&�ŉR����CO�%Z;��o������
�+����iܞ�@p�IhGj䴬=Cþ�>��ϛ%���N�e:�^�������Ů�2�g����;�$�*z&z��}1:�:�Յﴺ`�����#����g�ڕ3�bs;8�mGz�t|�1O*�2��#�����Go������.]�苭�㴾�S�Y�N��[���A�L)��ۭN�A���:�7���+���zo������ҍ�V��r��Lʝ�ZKS��Y�3��OD�b�x�㮚�}�3�5��7���e1 �(\T�s>���Q3�t��U��4�ݶ�����B^>�4zHg��v�m\=�3
�'�I�2���{���"�ʑ��'޼�=s�<�bvy^	Zw��e4{!�<�z':t�E�f�0#�3S���s���;z��-^����u���|^`U���-��f��ħF�:��e	���R.=~�5�Wxg�Jʖ��#I-V�ceqy��g�\j6�;H��3�-��s���R�\��>_�F{^�������)�W5?�H�ҝp����F�)���F���绒�#x��;��7�O����L撼�`�$z8��Ff9���S�и�*�7��Z^`�kϮ��X�N����ܘ�M;4n�Z����$�Nǌ-�/�*"We��V@��m�K|m�7]W�	:���S-�͎~�c_�A϶Y=C�i^\L]O��%�om����so8ǧ�<\WOi}��ƍ��1�5T���N�2�������'Kh^}�[W��IQ�NU��/�r$ۛ��ų�m���-�8�]�|�MA8�*�]�}+/ma}�q�3_roM��k���T:�U� �`��ψ��{�!4$�i^K�|^e�������h�������V�No��Տ�A�=�RA��&��|�NLfW.@�v�B_X	
ݎ�WI���*��,��>�(X�l�����j[��eNb�:�k�F��N��R���c�Ӟ��X�6m��e�:��Է��d��(��t�y�]��ClJ�C��knp��+`� ��Whn2k�QwU�*;��p�ܗƵIurˣĈ���q{�n�w$@C}�Ѩ�[�]L9y��[cAv�Y F�mt��M��S[]�3��_@P�1�}��G&��r���W��n��wV@������)xέ˻��S���<��z��왶�`����&|��ț��>�\3����<�t�c-�g�*��Z�M�=<LU�@�Ń,vo�J�Ýԫ�#1�hP6�>�R���U�.б��GN��I\���Ӱ��޽��!Arws���U�M�����������9gV�)�5eWB�����2��c�5}��jf��*���x硊Ip�q���"f}hp�i�`�"k�=�ie�۟sIa��R33�K/9<[���Q%�#���3g>�Х*���n�9���2Z°�ԶEo� ">��o�]��u�x�⻷�<��oD5J��)����:�h5q���Ld���N��^��C���2濺�k�{]=e�:b�n�����3�v:��vaYƥ�Np��� #�ǖk@(N�k�Nي`a��M�b��%`'��{u'�m�|�ܾ�50rwx��L�%�E�m���O�YpM���O
D�\��sTa�!]�6��J�8ޤ��G()ץ�����$j��Ŭ�x^��Oe�V�he �n.�	�:$�l��Uv�"��8��o*����u�S�W�Ilj�v��An�*g7o��O�Y�>ո��/��&p�8R�R끣�tvu����Kl3��IIB1o*֪�Ӛ
�7(ӕ�5��vnX���^X��QQ{�����N�kz�>���ۣ���t��c�F��1��b�p)�a4��]�����p+�$���b��7ac{��|�/��jە�|�v]8�+T�p�K�楱C�N��:���J.EjV��n�aku������[W]��΍U�n��-sT+�(]�;B�����Kj_:���-i%3Xlv>wӬ���M{�&�g�J�����w]$�i\��j�Xv8-��N�Ź�����o�8e7���Ħ�z����#:�6.��`df�C���к�dd�moV9ٕw���h�]M���A�ج���N�8sK�Ϊ�կ:�f'�_"��[W��U�=eP}x�	f��Yԙ�������X�>I�F�k)Ջ��e�q�fYNeNހn��b�Ծ������#_��k�cW*怱PFJ����)���69�&��r�X��;���(�I�L���\��E�`��WFwWHр�E�T� #st�ōE�cg:�RF F��#��ݵȶ3hơ)(79b�PE˻nF��F �&�(�ɯ�b$�&�� E�s��H�"2#EC"1FfH������&��b�F�����n�1��䥤�lb���0Ȏ�"�AhĆ�':�Q���1��&�#c����H���D�!��QF6��"��p�œ!5�M�2Z �&afW�d�X(�N��ZCb����\(�*�P�P  }�E���$�\S.\W;&63���@s${�����h����+3X��P�N�sGTU�9P���]�s
��_s{�������K�G#gv�X�����zN��/�c:ձ�U<'�5Q��ULNQ4ts�35��*,K��ܛ������^��V���d��L��*�L�I�7[��+��f �`~��J�5��xo�8.9�×(z�Ύ��tp	RN������v�uo]���(�T��e&P.��ʚ�ݎ�Y�S��~P\X���z�_T�]#^{�GwngU���c�B١���8t�z��{�u���3�1�s<r,�N�	�XΘ��2�>��z����*g������b:u���Z9��m�A�6tv��<g Ca��ٮm�OQ�߹��_i'>�H9��+��.�Tz)����j�5%��D=����#4w!��fG����ӱ����]B�9�����0n�Ez1U�����Ku�zϙ�=��Ѵ9eSpP$�Fg!�F1��ͫ���fQ ��8�D�"~��A�)�3��q��j�a�1��f����Sު����}Z��3�M��'\�2%�J��'�M[���7�A�NH���&���dwP(���!��ͳ�YV�s��������Ǜ�
�[z�z�ۉp�s�]:t�Go.ޝ�3-�ZSw;pp���
+��H��܈֚��Yf-�M��Fm��(�hV�K���f�J��3&��:���]���%���B�.�+�۾��hk�.�6��aC��Y�9������h��	��'��2�"{��$��U�˘�B]?�8���~�d���a�U!����E�$����2���FV �߮ ]W/��l>͉mfD����zx%��l���[[X�k���M���=�=�j�M�y:M�l/ЎU�W�������5EH.�=�t�A��w�0�VJ���t�;��I�iq��L�l�X{���';�=��z'�������>����>�:�N>�=�R����;��lv۱������gP��dU�VwV^�	�U釼�����ךX�f�}>�c�a����pI��O�ȵ��Jb�θ>�����^�� ��~`�:�{�Ռ�k��W3�8�s,�/P�� ӓ�>�Y~�d�{wK��<E�k��a�{��2=�$��[;�J�n�'���;*t�d�a�^!���{۞��4�t��ⶫ�Ӑ�B:�R�;�8�P]*�!�"}Z3$��(�C��7	I5�r9ܲK5y3���/��ʀQ�Z��z�x}�2�B{'8����]�����c���]�4s7�o^(�h
�K��`��קw�;�����j�+���ऋ[�oH��AjKn�mҚ�ϥ��H�	f�x�c��V��3 J!H䂮�W ��=5�u�Ne�"�q��*�Ӽ]$ӌ��w����
r���M�l��b�h�����c�� ��]Dt�Iډ��T+��JX���F�����ڕ�>�1�N��%�zH6Y���'NZڎ�m`�<z �@GfT���|��T��d�z��)��cj˱.^�<�;\r5�����N9�ah�(�A����R�"�Î�M�5��y{��+���O |7ܫF�ڴ<��hn7]�����N�P%��Ʈ���j-o�['�GW�2b��\��Lb�w�h��j��C�\K�387��-��K�����vڃ��j�o�3���&{iѸ���o��	�h�g-�%%:
l� k�����w�b���swI�/�7u�f��:*�Dq��[X*����G�Ҵާ�ɫ�>tЖ��ڜ�E{��CC�&KOh^f�Ti~�50����ς�����Ŷ��6��|�
(X��]�ک΋���8KV�Q*K��\����l�d�Y�����R���齺�����꛹�\N?�S�r��j�z=���+5Ճ��;�b�_�|o
'0�q^R�Ml?�{�ԩ��z�rͿR]t���Z[g�eƮ9��&33A�J,�A6�S�+���N��(�����"��yh]���u�<+��G�geY��=��6'�[��3M�ٵn1.H�����g^N�u>���&ͳ;��>b�U�8�7���ks���F<�V�qR���@��VǥS�Fr�e54=�u�p���H�f��9�7�p�WF߉���o�A�P��U�������˨��{��L^䯒U��;mJ�����Μ���e��>��\�<2�e���v���W��T���
�d�S̽��sxf�[��/cs�t���Λ�����^�����$�DL�ug��?)s�.o���p�<��앪�5[��X:�����gTSW��i�;�<nԐv�� >(z�����~yte���*��a�
��>/�[V&�lh���{%����D�0���QŒxf�Q���K�j�͇[O�He�͟r��r��Zu�Ҹ��>:�҉�aӠ�.K6*��21�f���.�\�6Y��l�>���+0*���D���{��ϩ�܆놓<u#U~���E
?~;��37O�_L���� jk�*H�J�+�̄j3��.5��EC����]����>g��~/bTh/Am;�-O��I+�|jR#I9�]�u.:7�L����]��Q�s�j���vب`���o}�Bs�PvZ<')���	e�
�x*�˩B�`�{�ۇ&Q�^��<O8b��tk�]�;��ۛ�t.T��R㳼/fl7���hM7�,�y�`���W�)`D���g�Wf��|8]!�(j����ݝ��S�_���Qng-	�
m8#����6=�Y�u�]��yy�"LT�ye�z׉4֗�����LsN�N\~�j2*6_��_qD�x�܁/�+��*�+f���Y�W)��~"����e��w�$��y9
e��9��(8ו �d�=�&�^^����r�뫪��	|a�*�7]/K��4_ۗ�ǚ�|}��fW�߁�ߦ�7���N�^;�]�fj����������P����L�'�Δ���lzUS�|�F.��كs8}�����]X�5�9���}�rNX�`���������:d�d��*�����|�/��;�c'v�(��._�x��x��W��{�\��'\��3��*]��R��裘{%����xopޏUyP��n����ޥ���Z��3��M�d��q�x�9��a�{0�燽�u=\k�4�t�<����9`��Lg���z�p}�>���7Q'b��oPJ�d_m�u�ʕ��[����;X$��[u���b;�w��c�h��o������դ^ю6�{m隸0������V�H��$Me!���Ϫdp�@�
��|�u}�.�0͡Zq�鵚�R����=o2��ǘ��ɬ�[G@v�lbW��#�N�\�g$ݜ���0��%��X �u�V��'RWfb2�[�j�B%��{<34�o	��FKE�]��;���i"���n)����?jKS�����E��7�\!8�{�⣭b�3��6K�� .��(	��0n�E{X�>���n"[�����V���b�#�}.��-�z��p摚�2
5�G�tD�)V�p6S(f}Nq�X���=�:s�)�����K�eeop��i���Cn�v�S2)L�zL%�h�9��|=��q+ͬ��5||�O6g������	u��/���s8�^��2*U_q�'lL�<̗/��w�3�:n�V�vQ�y�%*�3�&���w��b�O��ZJ�/�3,~F� �O� ��z��q��\����p���;��V�a�Ւ��ݨX{S�cК��~N�Sm�K�{�Iq4ja�ܨ�kҪυ>eH4�� �=7'å�xϊ���t�7�n^\w�'w�>����(��~��]#E�6K�;�97��q�dϯeƏ��8�V�����0���T���}ߖL��l�y�q��V6ⵕ������ךm�F|o�99q,~�8�S�8?4{(z~ț� �a�q\�k�����3#�Փ>YJ�`�_)�V�9C*޹)�DHa�Y��)�=�����v*ǘޱ�	y����'r���n@�1�h�4�L����9�-e��J ��n;�7�ov&��L����gK^Z���]��J�5��wr��rp'~�q�*@Vy�C�U'�S�G��uc7��x����7�Ne��^�x���)�R�7����a���= .��H
�+LȔ�0]JG]*�}	�p��ʝ>�y<���<�Y��h���83�*�OL�͵@%�B:�R�/��ԧs��a�E;���
�EMw�'){�ư2���s#��tԔ�A��We�*G~�j��ᮞF9�t�^l���9���f�Mʨ�O'�_u8���t+��d�P$�}2���
IJX�뢍��X��>'�U�"K�m�z�¨�~��d����G|��`4�/��x���@|
�t�3p6R(��wTO��t���
E��]��ܧ|0z!�v��ѮF����r�R0�\�j:��8�\`��#��O#tOOZ���˖��û�=ڴ=�9������鸇N�i(��W�Vy�dڿf4(����bx��J���|^�1��1w�h��j��\K�3��pۭ��NK��T�Y7R�x�������'藴��t�;~���3��߹u�7��^?s�~Fb3�Ȭ��#}��Ef��qu���u��.b�De,�B�f'X�pL��ᇺ+�zmp�ü����csr���!��S�K�l���o+W�N��yp<@��0%�7�����Ճɽ�nv�Į���T8�r�$�j�]+�x- V4k �뮓5(�e3g�¢V�
�����oJ�j{p�8��TW�*�[�����\�ÜL���5��̝0�N�}<6�|�S�p]b�b�Fw�5?U�Tb��*�֟�^X����c؜S�yˀv�n���xg���z�zau�2�*��>I���s���޾�{�a���wvx%�w��5O���k��O�lq��g�n i� ������G���oWUԸ�ĭ0���v���Fu�g��=*��2��<�j�f�F��r�j�����k��A�v�k��s.��Z��&t詗�+�q��1�T����b��ܻI����������w��přL~���;qs��J��t���ղ�4}��p���&�Z�,T�ks}Y�ԃE�Ǳ�\$W�������l�N�$����΅$��ȭT
����zu�o��+��%]z堰l�_�^7-��SW��9w�x�Z��@@|P2/s��m�9��~������z�7�X�N��σ�1�s��p�f��<k�$��z���*��s1���g�q��tw �|sm���S6yEIOb�2ޫU'c�tr����B���n�	B��\�48��Y���5��7�����]��$~Ywqʄ��0N�\���`�/��Zm�iξ��ھ�B�.��=���o���|s�@@/���iϣ��K��D��i�CYM��p����J�T����jg���H���ls�MS<_�D��t	��ZM���VB���뉹o�����:�O�'��3��}U/Y���n�r-��MGL��� Jj �"e*�cJ����g�\j7���б�%_@S���%�Ux�<r|�mށq|̢I\D��A�"bS�uԸ���)�F�|�Vvd�{���[y֤�_�'Ȕ��*�$W���31��ׅD��h+��(�f������һ���i\���ܘ���f��r�k�5��d���0��|�ƺ�1�un�W<�6��J]x':{�J��w�$��_���m�`���5�d������edM­��I�:c:�������Q�lhܯS5T��r���c�.�WE�z�����
z�T�2��@>	��P���>7S+	���L�iS����2�j+.����zF�K�����=��+F�j�8rY_Q��yZZQ=��=X��g�~��cJŠ�wo��� b)?�m�C����vf���Kz���h��U��e�X�G�|M߇��q�r��_�o��y���O��I��RP��*w
&�i��f��4�G�*l��d��u����`�]R�AݻNH�\Ol6�攒���Ժ�^��94�3�Nq�j�{����
���È	�^���~����|^���C��T�{��º��)9�_х��Re��M���K�3|�8�}��N���}Iq��{ݻ��Z�Z6{��OS>f�UW����9`��Lg���K�xϴ�v����7��%��8sϙ;OĞfbѯ��/�2ѱ]t
�RYp�c<7薎y���A��W�U+���Y:���c��_#ėFa@��;���f����nZ���5%���o�gO�v��ό��?b�G�!Yi��
��`�=Q� }5P��6R+�b���I�����fuP���U@ �߽�5_�~�}3�{Kdx��p摚�2
5�G��tD�)V�ce2�w�u��� ����we�8�������#s�C��%�Q9�:�d"J>��a+D
ј _P���wV	�G����U��q�,;{�F�]l!�/����%pu�*��2���'9�ꨮ9��	�n{]�./��9��n�R�	Pt5��qi���2^�|?}�z����V����խ��5�ڵ���m��m�m��m���mZ���mZ����V���m��m����V����խ����j�����j����mZ�v�mZ�~V�j�����j���m�խ��-�խ��m�խ���m�[o�m�խ���mZ��1AY&SY����ـ`P��3'� bDW�w�*�"�Uh�$J%P�Z�D��T��	�R��@�I
��J%@)T���(�
�J��P
�T�U6��
v���C�����FIB%*�*���֖���k�����Eze큣U
��ӽ`�A
��[l��A{}u*�"����H��R�A�%RUu��YaDA)%D&�� I��u�T�R��BB�������TB*�o��mU�UTT�^�u��  ׽5��ν^���ޢ��s^���oZY���-��΍kwlp�����u���5�R��w[Uv{u:���5ƖQu�-Ӱh:�j��E[h��
�R���  W��b��zovi�w:���������|  ���  P���=��h���n4 z4hGB�u� Q�::3R�:(��� 9��F�(�Ea�UU*"��JU*)S�  cE|�R�çn�cp�9�%�j*ت;>��@P�t���j������ٰ��h��[�nݯq���zЧR��TCѠ*��T/�  �}�����;��2�0��X�)N획�Ύ�,;;`�Nݥ�/j�+�E��%&����n;��\���ņ�{��ݢ] WqQ�T�+�X����T�   �����l���\僚ֲ���뜫�n��w��{u�t�=g�Uc���wݜ�Κ�K֧z�ܪ� 3��p�N��]���F]P"ػ�ש��[��(����J���픓�  Z{Z�mW���t���thi �v����V]��9l���K��u�m�w����7�wOTw9k\4讝Wn�r�;�u�b�M�t���RH^�����U�%"��  �w��M�s���+�ݝtn��X%�N�E�Ը�J
ݶ���c���{�#QV�=�g��.�`Nղ�[�b�O/z���]���ܶ�Vۭ4��̄��z(�ڪ�_  3=�e�(�Z��s*��zq�kݥ��Y�@�*kWrr]������íN��8u*�s�4J���c���ͻ:k�m����SY�z���**�
QR�� �揣��[v��v�ݯ�]�KU�T�:u��)�z�N�#<3JV��]�S�kwwmN�ӥis:ofּ��{Ã���޽��\�
��uÒ�B��M&̻*>  _S�m��J�͛}9:��r�]�7]-��봝�L�me��U�\�mۻZ���Ҕ����ݚ��c�zH�������P�jwk,������ "��I�T�   ��1%)I�� )���JhA�)� �����@��4�U2�  ���E@��������K�t�����gA��t+G%\ķ�����������:��TA]��QWB��b* ��TA_�
ʢ�y��,����Vu�������ޑ);m��31��wY�f�X+["��U2��en��ӐZ���Zh���iwr�
r`Uh�T���-cKiM�RN��RBWef����H�v;�n�2�ĥ@s/QD�ja�/T�yBc�J
W�	�{6Ѡ�1iY���5���؍�{eQr�G J��09�y��1�q-�(!��l)����k���G�1��h���_͖[� UfU��lY�ى��>�Q+qk��"�f��t�m��,�;�Pı+�c�UwL��^�)<�耳y.�kb�Jz�2�`"��5n0ʭ58���0��V`�22F�1Rj�P�3�Nl9Ku�ulӳPl7I]���O/$����E�E����*Di�t�O1�j��ًp�e�"u6�P��/r��Mw�|�eZJ�K�j��Nѷ�(�N�حg�.�����ar(#��M3E��SH��cG7^c��n�*�36�î�ä깉l�n0�-S�ncGoS�P����)�F������
��V@U��wVN��;��ia�3)�NQz�H!6(�I�!�{�7D��G�����JutB��C�y2M[Xi"�e�C>1k���{��D�ܬi�Ө�� D�h�����|�Ղ��2bZ�\`�Kp-�4S�cK��*�4X�eec�!RB�t0�͌z��"�-wh�w���3#�5�*��5"ZG4�5�6�D��
�2җ&��vME<�5���1��TQ`w[Sw$�M)7j�$դr��n&4��G�X���^���,�IYH�Ʉ-�jq=���R)�M�9���k��
I[��Z����G��D�*kv`(��4$�7�Mޭ�of�3s$f�/`�dU�x��Ŷ"�v5BV��1v*:Hb�֦�טsv�D<�8N�!�71�%�//77K(��^>ݱ@�R�#��R��c
�[�h��2]��Z� ګ�R�^�^�r^ؽ�Q���q�Jf!X������R�ST�umm�*�G��&���(р��gY�(]^��r��j���\4k&#����p�n���6�:5U�zaۺ���ט���,��Ս��Η��M9�P ��~r�����ЍY!�#��ZEM��c&�m[�HW�AZ�a�U�&%x]2�K!v��jbX��@���Ax��p
���mj�u�nfMn�uh��Pf�&f-��*�H��K2n-rm�*F�!h��W���ݨk�/*;p_����mi.�ctd�,�8 ӧ�܎�� �c/���l�	q��K-����2fjt�8e�Բ�eJu(���m�q�<���N�%��Je�+M$U=mc��0C5���T��&��2���YI��G7a��**٥�+5j�اr+w���Ӳ�����+P� t�!��Y�m �̓]ʙq��j�sk.�����Y��[j�F�,����5��i\"�m��Փ2�T��VDy�U@CAd/]<���(��M�h���B]�Yd�&��8.�P�,G0;�L;�F��NἽ���E��*�0�x�S�Z�jܡQ���-4s(�����9���ۗ�Zye�3	gw5p�0ح�L)�z��̛B�S�z�e�Y%8U6�3t
�xkM�݅��d*���E�ݪ�K-�eL�Kr�L-��T�j!����um���RV�ThDl���%�5f�֖���`k�(6[7�r�Bmn0-M�L��YS��n���u8j�E��q�PMY��(%���3m܆��m`��ƂB�Y���@�d��,�Nm_�fL�L���TĄF��CBD.h�P���M�)۽A��zAZ��Bm���hɮ�Jj��/�B��5m���/"�P�i�շ)���iɚ�[F%S+v��:�9X��C����&i�$R��6��t�<�5u���,�J��)왷1cZm ͍z�;f�Gs
���o�+o+)�I��>[tUhŨn�[2g�V�-A(�(�ˬU�[).[��M]J[�*
)��l�yW�P6b����k0�4b�����d��g�ݷDlȍźTȖH��м�����C.�E�,�Wz$��P݀��9x-��b\)"�o۴����]��5%�M]��rU�4�ݪeӽڻ�>���S����識��V��7.ࡲ�a�Um�rč���-B��Z!��r��Ou:*��Dٺ<�V{{i
dV�ܦ"��ׂ�\
��#V�ve�N�e��YIy{�t�����1��l%J�y�&��T�oF�Hz�6���b�xa�nN�~Kk���l��*˗�B��1ފ�l*�Bdb�,���q;��Lp�e˸�5D��6d[�$�N��b4n���)�X ���i��.�G�QL�!��
�W7k2�f�q�;�w��u)"�
qSwF�\b�z���{��lnVbu�A�!4�dR��ͺgR��,��2AZ4U�&)-�B^�f�Q��n<�`An��陖�]lr�hR��toMB�U�V�X����Pթt��9>K �EJ6��v��� ���xq����WiT�M�9ou�@ނ4���ٙ���G�n��aȯcG�[�v�h��fP�.ʭK*�VA;Yr��*��1A�[c5TšT AxV��Yw7YjJr�[�Y��2����ȬX�R:µ�^M�zq�8�k�d�Y-əs�����4�$F����x6�-��%In!�˺�6����O)9,L��a�naWB�8�+L��Շ�laL�.���S��hŲ�<�50ұ6޸��� D3�T2�'B�-V,��]����B%�l�]�1��Uz&�gd��P:��S�̹�뙭�ԛS� �̗!�wJ�݀�N-�c��v��@|j�Ӛ6�v��I�z�s�ȓ���H�X�3pH�o����	J�V��U��,�F�Y���P�&�Q�Zp�����A��_ٗ�aָ>ǂaMmn��ʕus�ŨLe Yn�P鼎����v�ul#B��hf�8b$�c�BP��bГ巚��=b���Gi"ë���Sv�3]H6�q���֌����*WV�l\�y%��/m5�iڊ�o/rѭ5�!f�2��, �t�ʻ�f◘i�V�+e�7�^�4&�MϤ̲s"��5s.P
�m�	�˲e�,��N�j�p�!",�)��Z2�ATU�7��85 4�(d�G�ۋeMx���[��Z)Le�Q��t�Ŗj+�/Qm��MՍ�n꣱En���#y�f-ŀVi������"�}-PtNKIX��m��'waNf@-�v����u�xұ�V��'�Hv�+8�ٌ5���XxT!>�X�q�b��j#�0r��*���U�d�Gt+*Y��/�U�)�m��������d
�һ�O%藂�����N�D�P�K[�Hi��t�
���ӟ^&i[��E0-D����.��0ӵ�٧��d�CN��*ŗF�K�`Ƙy-4Pl�(��'����C%�%��Քڹ�U�Z�fB��֌ͽ�&fb�)���۳�����s�2�MU��`�/[��g�[���A�F���b����(��ț&'������<�.;�͙!-"���@iS,��:�
'� -u���RZva[n3dE
ߖ�I��Zan�2��	��YA�̽��!̴�j�z}���yTe�X�v��7��R�G5PA������At��e��Ac���]�P��N��a�NmB p����e�+t�pnkjb���z�i�V�N�C^5/ �9��&?��!�-[�a�Q��D$�V��2�#շZ�רI�Ev�iպ�CN^��1]\(t��+U�����1f��	�,S���wj�;��@���	Q����&�ձ�m\�N�w`\+j�Mƛ�&��B���]i8�+Sv50&oJ��ӔMSy��6�p�n�׍�U�!A�d�~Z>4a:�u��D�񀜢���ٻ�Sh�mAv�j��c֙mLtޗ�sE(�)��ur��ģV�^���V�M.%zstm�C-�0-5K+�pl��UM��J�Ibl|c`�%��Z)ņ �C���Z^7[S(օ4��쎖N圚  ��h	e�
h`�r]���v��-�	3-�72��'6�����r�J�a����N�ܵN�������c#�O&��϶��<;C6��kt�F���)�7��[I]$*�R��wkVlі��9��n�:V�Q�W����k�a�Ե�q<m�F�N
Z$�ƪ�����n�ɢ�3+n��q`z�6��0S*�4�2�n��;�Z3�,���q�l�
TE����ʕ���4^�&��ĥ�n�R4���7n�̚�`!��Ę������ғǁҔ��l����#X�"�j*.���a��d��ď)�!y�*9eQu��H�e����۫G���Pc u��Cv��a�܈��`�ɷqj�v�)h�!*�L��i(�h�ک���,Vݜ`�}�n�����s�e�D�)�R<rm6�G6�'u��A(	un�QQ̫@��0եKl�U3�S�m�����S�4]Ekjn�n�W��aͬ���{#���"��[����*���Ȣ6�á�#�xkv�2b������`�t���4��1�u�+�6�pH��Z�i��k#ڷ�ˀ��6]m�{�����˙w7j<f��;neM
#C$�r���n����W�fZ���m��0�&��2�]��̓i\I�0�6E�]�V[l��j�*�c�u3���M�1�q��8ZЂy�[�����jda+Sh�����;���%�ԡ�����Y����w�N���W�R@c&h%,j�^�Dp��&Pt �ݘv�v�%b��k�eJ[��$��tD���N�u����z-F�tER��8�Ɔk�wӶnB�X`����v�,G6Vb�!�\B�n�*��˫��{�0��&����&� ��ًi�V�fbR^^��G�Y{�h�ۡ6��E����M9��CH�e[�ۛ�Z�
��y7)��`A�lǘHZy�i�^VK��tm��SFު�!]����Y��Z�ij�4C���8�K����QSv,�i�n�W��*+L���N�D��X���bAE[Pʵ�n8�����DiC1�+1݈���/jmb�M��[ف9����\�`M�f�Q��[jem�:{n7o4e10E���ٕt/skր�9�FdH[�N���*,���h�f1nۄ��Tq�C��u�f޳�e�.A`�᳼eN7���vf[�1-"��ji�M��5����N(���a׎�O���ܫ׹50�-�^�CV%��T���M;�*��&l�f�$1�*���^�^�͘���D�]E�v�*���_V`[t�E�_N���{v,��}e�Fޔռ!�%���՜u��Z9v�3m�On+%@%'Rn2��uvq�����zV(hd��H��ː�u�&X{Q&��Ŧ .����|rT��Y���R�ɕ�5K%�Ux�PF����t�5�a�.� 
՟.�c�������3n�*�YV��tJmc�/L��%��D�@P�B�!��ʲ�P߳��)"�vRg1biC��d�.��Y��ۤñ�7��c�u��R=1 �ܛFЊhո�l�S��=ծ�:tZL�?n�h�v�p������b�C]<8����w,���]��Ш�T���S˩��[�Vչ��nX�'e��wO�"fX%��0�+���A�1k��6��%�iϱ��r�(��nL�l�Y�[��1��Q34KC5���w�f�즢X��՚�k��HM��m��deڧI:���ᬧEm'W��c$�m�Q�K��x�"�e�����I�ei�M
֮ǭ����q����[gZcV�Cc�$���TYUԇ-��\Ɋ��N�V�[�ùi��b����޼�xW¦���q[Z-]�M��lZ���iOw��9E�uou�hn	�wp�	�v��Dz蹹�,)-��%��ը~XidA!5D�<��E�I@JO/1Qe<8��"�]$�p�*툯�NC)�ʺXܖ񚴇#5A@�*�ҀC&�f�R;
�.ɫ&E-T]ͻy����CD�նC*X6��tv5Gr���n��*��� Ѵ��RQV�/o��!Ԡ(�	Ӗ(|�ǁLf�
ZP՛�V'�3`�AtD:S���;�+`�{��I,��ٻ�2;�Іcj�Y&�� �Y�XI�3tИ�G�mC{v�ԨDS�v�`6R��
�Hi��j��72��b	�9+infm�.U�EcWB�'�m�
�]+���,L��L�0�f�J���ՙ5<��b�ڥ�!{��%+.�Ti�㽠�%on���Z�sn�*��#3j0U�t�9��4l��r���S%��	�sVZ!��7��pb��-����[���>��K$Mɗ)��$j9 2^B��łʖz1 KD�Ț���d�^:NcCp����n��Kq�%�w��fedX@��.*'i��ݬ��Df@J��vŽ�V�72�.��E���Lf=�M��yw��IQ�=.$�앤a&�Fk�A��d�`�',*���U�m�I�Ѩ��t5醆:W���̵�Cr2^\4��b���ڎh��76\C�i�mj��76�8���|%^�۫�5�V]���j��n��`I�.d+�b��˴8�u��=Y�7��Iێlv�H�)V6��CCl�,�4P� �+wea�Pe-�t�U�0��/s���9��i�^ל:�Ց��x�q;W��$��Tį�B뼅���0?:�uf�ޯMZ�;��F#=ko�U����#�����0fl]��u�����a� %�ǹ��-�M�Uy���oM4qR���9Rk�A�]�u��\mL6*c�3�K�;p��FR;˸u3On�b��k��e��Ե����R��ج���n��_rYܬk�MS:.l	����@ʸ\�cyi�2Ĳ��k�8�k]`F^ID�/�vm:q�҇�̀�%�VĵR����ƪ�����Ѝ�h�e�pb�q;�z����n{P��V_��c�Q�6��2�n������w�_b�V��ǧ�wo(s�V���S���^k��]�$�uo>7ҏnPͧC�B�(t�΁*���3�ʚ)��NW|E��x�Ψ�(3��n���
�vK��Q��pZp-eMV�����U$�n5W ����v��{�N֪9R� ��s��E*�JK�%#�_�"��븣³�a�.�Ĝ�yp����G���'��h|�e���U��-��О���V�:���"�r�L��V���c���ۻ|�.��X�� ��v,�/k��V�`+
�����I@J�Z�+x^XΏh��e�ݽ�\��'�;zs���4X괳
[P�����NE� �R]���'���Їkv�s;+hr�2�_#Y��ዥ�菴B)��چ�ܒ��-˳+E��˴=��\��ʕ����e7�����#h�.*�i���!��d�2������!��ն�a�;"��)�\V�wQљ��b���W�k�N���K}n�y��5Ozz�٤z�]hZb�(1u$ŕ���^��v,�Mb���.fQxEK@v�tS*M�[�Q��'�P�%n�7��6a��ɨ����>f����A��85��6�c����k��i�K[ԙ[WP[ۗR(�;>��&k��#��p����En+�̬P��ųG|�Z-��:��Y#J�u�n��}8�Pb�-�3�E^ܽk���wU�9�;Y�����|�b�.��aě�[��;'E>�]\�*��أ��&�Z�ՌЭ$��c�hk����O&r��WۙW�&�$h�̫tC��4�b��A�\�R=���5����-AU��E�wZ�27��(E�6h�^�R�L�V�=�D���
�+�������W�[���_k�]��������Ƙ��ɜp	ܴ�][ДM$79K
}m�f�;;�iS�4ιW;�OݸU��I���5l(P8���͊�ټ�[h�d�{J�Huw�>������n��VJ#��e�Y)['3c��t��We-���4�]�rĉ��Z�����V���ۚC���A�c�b��/^ZF�� � ��䣬&إM�{�o,�6�Ү��i./�{N�vs��,>��pff��Z�A䤸������-	W/v��"mTw]���@8�G��v؇�����&:�{��ν�y�!ok}8@*#�zì�e��A�jf� �tn8�΍��k؟SGJ��Qm��(�Y���,'����e�N��F\�w&�Y�\�eꡍ�1K!r;D�*m&����C�ږ�}2s��|Q�oZ:����������cq¥`u���ױ�e�,��K=���\�ڵ��}j��O1@��d�Г���q�ה�EL�D/���%�(�ϳ[�����WC�ݫ**�3q̬n���t��/4��b�)`|R]&��	H�4�e����m5��2�*/rv�����}NmM�CSD��|�#���s�m�sheG	.���9�ʑ���&��|!}��ۛç�ӏ7�:�ٍ�*�lj[�gRk�VY0M|����CEU��jP��ܙi,w���+�5nL˷�§�2J�W�:t͇�,\�h�.��.r��';w֫S�n=;�eH���GE�n���3ye;U)�R���1dٺ�Ϣ�o���Wj�=ي'�Xv�����ors� ��I�׸�l�|�Z�ڙ�6a ,n����PHK=˦�LM�Z򰇏!�Ծֈ�����t����*�Ju��l��li��qmN�1\�o��2"�Y	�=e�\o;m*�3C,���tm��.�jvH��g�^u�^Ý�M	�&lU����"��i}(^^��;�<��z��|1q��fm��#�#�f��.�1��8�s���x�N��Z�2��;?*GM�\�%�rq�.�#���B���e��v����5`F�b Oz7��Ï�
t�����dJ��\-�\�b���S���8�׏P����Sd�5ě}{K�]|B����j�'��9�k��3�f�Y޽U�Ej�+'��!�W{I6N�s��R]{�l�V৷\j�Wֲ��M�٥w[,0�����j�C��B;X9K���W�X��k�sD��ҹkW����۾�"뒑9rb���|�>�˒���2]a�=���+��j4�
a��x+M�v���Hauھ�)���Ȣ����k;SR�C�㳔{��K��:��}#nu�ϳ	�����SdgP|os(���_��l�.'���ѭ;�(>*�y����H���)�GJ�;"�W�󗯦s7���t0���x�:h�4�8�-�*u�+���K��:F��C�1�"�&�n��U�������H</֩o6�g{e޺E�1X���Ɏ�ǒ�Zd��o��E�%�AAr�u�3tGq�/hb®�L��i�]*�����2L��B���t��W��6N�ox�	��c��d;sR�xN}�Wk�;#�{k��-�&��mn��-wu�J����Gx�u1�|®��+*bɷM�ǔ��kq���� d�쑳u������������)�ִ���� �h��\�s�]�	�N$�3q�ަKUj�ZѼ1+�C�ɦݒ�јٰ�Sѷ0��-��'n���M�_c�}���=�9n�s&`X�`^i\��Պ��v��8vX�<��T ��|� M����s�p]q�j��sn\��K:!	ɽ>;$ ^�P��h9���K��
�E��Q��!��P��cis�	o���ii�w\�Ǎ��*]k�Mn���%v�ۍ(9U��o`烓�܋DH7p�*��E�u��:��W��k���\���W��>��oP��d�xݚ�H���a�����t:��VY����%cW����bIz�@�U��Y����6�Ӭ�ǐ�ͬ�oa2�����]�:�7+3%Y���6�eO�<c�P��ܶĨ�.�Ǹ;�;�9v�A���w5u�kIu�:m�#.���k�U�eu'�-�啭��]%����1=/��z�Z��-m��h+kpk��ݏu��+xP�����_k�O���l��Ζg�K�z0q�OWJY�+ȗ�t�&�Bې Kf	�*���qc��,)�e�T{��/�wF�g#�cb7Yhm��(�58�{N��Zu��,Rlk]ڗ՛j��邍ftLX��v
� Q�kϲA7��p[��m����o��zr�r�\(�KW��ͭ;}m_�-�n*9�j��W��D�y��5�P��*�Omt0M逛=[��ñi��ש�o�Q�P�s7���m�B��i?�[586g�n�u�4���U�}��%�R97�ܝ�a�)gC�q�!����p�.\�6*Ցu����\��;�>�����ƴ��Dz�o�<J�Юj�ٚ���t����\���,`@=�l7�f�z��n�V���`V5[����x��B�)V^��3ӳ�%�F;$7�w5`��h�WQ�TyӺ�.��������w9�.�VW�=������[��l|��}����#k#Vjob�Z�0��>{!R�z��޺��u8�k5r��u�+9qTrqV7���E�{�o��%y�(�ޚ�<��G��E��\F|��n嵥;�緓ve8^�k^�ϗW@\��ʒ*Odu�����On,�0y�P�%aU�dgNB�#��7��ha�*���Ԍp����VE*�rػY�}��I<]/Wm�6�BQ�������u��R��n�M���}��w�RA2^0/���,�kF�'-�ۨ����Ã2��GS���O�E@y_�cG���r��0���פW"m���t�7�X���xQɁ3�z��m6�V�zT�Z���C�i ��%]�����͸�pR�
,r��9>\�'mAAί;k{ �\������SI����K2�tI��6�����:�y���7��N�E����S������	χ`Y%k|Nk�w��(}|ۋS:h����r�GD5��s&e�;O�Q�v+������w�u:}s.ƊO��!W{A ���!z^�0�v���ؔFb�Z�]�Y6�v������5�.���]��bn-��O�j-��QF�x��X�u)�%�U�44j�}�+��� 4ޠ�5�����6�ַ���\Sw�S�>O糗ce@�{��;;�8Eγ�hI6��B]���0�M��;��G�Yt��:�u�Y)mJ$
i�����ì��x��96�é1���4��+���<;:���Y;+���5J���I֗�������ڗW��'�ไl��xk[��O��9f�+�LF^vQ�G(#]M�g�꺍�:+]j�I9�Շ�61�ّ��i�3;�^fc��N&�e�=	�O�S�����j��;��)W2z���S�O`�X�[ǳ��ke���~sN27(U�\i\�����P�����T{9�N:�yx��f�(d)p�7���z�'\ɑ�f�&X�Wc����������s�R�/�������-d]�j��9���ǎ�O9p*rz���ڻ�MO���
��Y�v��l5�5�:�z��4�:�&��a�>b��yY&�̪�5�c�x.U9f�Uؑ��=�9
��l���E�w۝�V�$r:Y��k���P
�1*AWMWcWe:���Oszf�w����B���L�(13Ou���%����s��ۯ���Y}�ڸ��݃�G��
�옫��7۩ܞ�v�*&j�ݐ)}����V^R#�6���7���ժ��Y��6^|F�_�gTQ�������n��M�.s7`�ڎM��5k�ol޴;q�^s|+W)��2�JC����p�f7W�Vp�g��}����Z{�I�{�w���P��f��ƽ�~���i1��؏��j9a���+��3t��0\����K:%QJ������#b�[�"��$:mֆ�u;��s���]�7�R�	�Һ����0g@�swti���50��,|
Ӈ�]$�ox)f��Y�k	�]C�b�'���F�>倧BFb�(qg�Udi������(H��Rpk�58��2�>ѫ�^8��teM͏����tQi�9�>[����x�達j-�M'Ý�ZFb�{*G��b���oo"&�]k����{���&VV)��9�Қ�kWTٙ��;#)�'p�5�"ɿ�B�*uݴηժN�(�kL�ڑ���R�v8eF;@i&x(	5��d[ܜ�0���v���p��>��)�X�rո���1Zۄ�>��[$�n˳�v�C��cY��-S��uI���\�Q鹬��,�n��.N��,]'4�Ǿ���E�qc���\��oT��y�9�������J��a����N(���S�@����g���V^��S�k�{��7Y�2l7g=�j;l���c�H4�v�����6�iJn^[����feѡ�i��9��.��M����Em��I��S͹�η�e�Q��6�%Ȃ�|�3��i�G4_>�CI�%�V��C-���a��x{�t�|~�A�m��P��}N�	���\׳M�+�v��,H�T��2�%�q���V��3�%C���jV�	�;b}���wM�O6�R��z�����S�8�uFGFK����[ٗ�W6[;��K��.NG�����U���6T��um�\�3+\R�f3�;��L�V��-�L�RݸzZ���q�w\ck�t��:5����2N7�79a�U�q嫰��-ӱt=�o{��v�`tD��0�׬�4+oc��Ѽ�E�UOwzfM���C��E�jͧ�P�N)X}D�%]�
%a��v�vb�u����t0�;�kфJ�.`35���S�혘�,��{��������w*{lU�Q�is}+9k���7��`�c���C�6������]+�V"�6��5罹��V�1��ߕ�
�r���>Qj�S�~8���zi5ʹ�ꙮ+�Z��\~�=B�ŸRPG��=���	�ևX�ݖQW���-9Tz��2��JЪ�gpDw3�^����>��'�XFқM��2��.����)O�����ǣa&��<K��;��o�>��k)"�{[��Iq������<��6[�)�N�mn�V6s��Q1l�t�����!������F+��� �Tkm�hײl��� �|���^�;n��M[hv]�O\���C]���_���W�	���Ď�{P5�@���Ӧ�ck�r�\쭛m�ǐR�����җ)����]|�1Kn^̸�3T=%��`M�� ����_c����ޮ�FU���p���J�=NY���4�u�I�H�MV$)����Y�(�
{P�����
����+h�!v�^R\�<@mm���f�gq��Au��/pn%��&�3�Y@b/u�8�k����U�}ϔA��dEp�j-�֙�]�U�tn	f��n�;}�P�\�!C�N�GE�9�;���
p��c�G�U����c+�ct�Z�i���k�^�<�xjh�O�{EI�]D�≯�m�Q&�vIӼ��{�߿� (��"�
��민�}}��- ۺ�^�`
F9��Y���B��
��2:Y�����hԑ�$����yC\���z�u}��5��'�;v��쎴���dJ#���P�0jc+7�Sas��
k���]q?��e2�f6�� ����{X���N�n���B�-��"k�ԫʻP�=x�۫�ڪ�J�-i� ���癫/�dTV��M�Q'����
�8����(ڈ�٭�.��Wvn:\�e�6޽T���|Ы��ZԱ�Z�'�ml�(� 9u3�_Y�����q�R7dO����˔���<V��w����mf)�TZ\OK�չ�����+��@�K��N�ko]��%-��l0�� /S�܌A6�����5e�r���]��Y<T�)'�y�/.���6!]p= �Ȳ��ZVH�S�<�)*Ƃ�	Ӗ�X��p[A��A�r�a�%����hT�����&���ti���4����; ���/��˪
˛�#��Z��w�j�3+1ȹՈ-��9Bu5��g�tvGH_tk�"�s�B�h7J�����i-^�9��5��{|���� q�;��g�����mP4������Vt�dif"Ņ����`�7�*]mR���%I5�g8�>�.�	E�f� ���ve.�2^���:��j�eY�1zٲr��	��u��H/���f���v]�ba�9\�3n c�ʢj쫕Αck�;#Ki��"�������k�mv>'EGC�	��R�Zf��9�)�O��Ꝥ�*��8�z*�ػ�����8�2�\��q���U��}.�s�`)O5�=ռ��<=8Cs ��0("�r�@��N�ң��^�a� �O4j�|mK�z7�	�L�ڷR��� �;h���ZO�f�5u&�DXs]��#_+Ɂw9O{Wf�]$��
��_\Q���4�}ڍt�okywP̬w��ݝ$s�^nf)կD�Nr�༦�V��0�V��흸3+�J�;�4@�ms����t,\�z�s��NHe��ք5�`q�wys&`�m;OS���{j��#;%����%ku�4�<�#k��r����m����ݥ�Ч�v�(^X�z�\���1�5�~T��fr׭,��V�kd�ܬ���9���Ǚ����1EF;8D�1S@�۳���we�HZ<�gh��5�kQ���LXn ,(
�°}w2h+�<Sz�v�]X��7�m����Gv�ѯ��Ù�э�����wq�XҤ:��"eM����5w6iP]���a�Ĵ�R��N�\��
�y �J�L�����bZR�[��)0�p=ˬǵԥ%�� ��]�o�5g�p	�`e��nu./ZwwE;NJ�Qc ������U��[5�z3)�Iò�m�6W;�C�������.NΔ������\�"Y+���:�+�����d�\��;z�t-\A;�|�G݀w23$R����k�a�YB�C:�*%�`X2oY&s,SU���F�7��X�y�D��L�j�}�WaF_O�=Ϡ2���2����܂��!P}��\t���]k�ٳ��Rʛ5e\�B�"�	�X"C)�:��p��J�߬-a��Nws�WS����}��nSB���Ž-�r�nS_U3*;F�&+h̷�xn��2�AJ��
����9�^�s�B�F=y[i�mU���WGVM�:����K��8J]�	��sʥֺr�j��`t�Lh|���^Q�� '�_h8��PS3e5 �w����[�1F�vWn�ˬ���K��KC�V�����4��z�u0bӫ��z�]�V �rP�����&[�++1�׳��qf��'fca�[_YK��Űy5e�ӫ�KMk�Ȳ���,���Yw�	��{�"ot�-��t�.�X�D�&S �\BoVQڙ��o �.v@.���1-ȕ�O�H���F��:L�uwW+�: m�CY�mgKp����i�N
7v��;(]9��BTi	�[[m]�Mn��B��R��Ӽ]�d�]:w���rYn�.��` >�P�Y����ѻ� 4�׹y3z�+|z�u8P��\x��:ZF_b�@���>�y��,W[Ä9ޅF���Σ�  fѩsh`r�T�Կ�z��k���B��w������Q`�*�|�����Z;mSx�#�6����a@�,��,1B����I�㘺�g��q�sdKRdV�FB
|��E�8�I��Ѻ�2��T���:���@�si�H�SV0���
ÄQܴVؾ��nc�A�'�f���T�����Xg|~肦}�k.:=m�e�C3T+P�NΕ�y�:�.hI���*�Y��E$�"�˙a�z��y�]�����e�)"H.6��&f� "^gPWc�u���ѪDn/��Ĵ=b�������޽�X&jym�'݃Dܘn>���_$��rP�6������7��웫�]$ͮ��h.%�����M�=vL;[۝����e4]L�Z]�8�!�j9���ju-��WY�wgd���F� �iR�Y@T������Y��o�3e0[��S��5m���G<�"��J�J�Wc�gAM4ڜ���2w��p�K:Pm�+�������'���֯�+�iR��߬Ffu�{���m�s�Ы��d{��m�Z��.^��?h��sf*�����hBeu4b��YA>��fR.]��J�f�p���-�y��xt�i�5snޙ;nε��)R�����|U�`���F�7|���*V�5��ş]Ƃ�far�m�����7���H����e�d	F�h�,<�	�L]ӧgW�]p��m�B]�vyG�n�h2y�����8.W+�ŏ����������[6��E)��[&VL�]1(M�����n�N?����b(�r�٘��p
4�w=�A���f�+6)���b�H�hf'��4B!�Mҡ���f^]1����M̖�����:tf]�s]�nť�.��s7�7Cm(r���"��^Q=L�������dB����^?���SP�*�4�Uq�w��Ux%�3�a�^�I�5�JԗS�
]��\=tp�[���I5@v���GJ�����eA�����ԕ�K��5Xւ\Ҥo��{�&���J�����ѲW�af
�m:�v+�aN�N����I�{��|����	�C�\*���ǭ����BU�c�t+ ݙ;J��Lҩ�s%[=ps<n��ti
�k*C��H�睝MGgN>�1:��FY��K�����\7^D>}�ub;!ޏ%DU�4��3-˺XTE��|�&t�����d�aR]*�[8),�s�Vfl��� ;�uz��������SMX)�:��ރ9�����v��8�72�wQ�h����jN1}����q7��4��e�룐]���xF(�ώr�}W��}j�[t�*�7�z�*�ND�iu$�w��	ά�HQ��2�R�g>��>�[��,s��+jֺo�ǂ��ާaݫ��S�/`�ɑ��vs!�M�N�
f�{6�)J���Wh�Yu�5)ز��#�%�$��Î�(�͈m�M�+�7����ɀ*��;��ݕnb�7t�u� 4�ʩ[u������ZP]���d+IǓ��(ީ��0]ʛB�ۥJ�T�N��h/Sױ]�Ud�W ׂ����|���ʻ����G��A���2n>�j�;q�5�ue��u�L�(>�G��]*�b��ab	��[*7,�Q4-��-X\&�lBw��y��&���$�@�7�Z^V,��2�WZ���E�kꇍܲ�x	���VnV��\��2��6���|+>��BJ�o	��"vT�S�;�[i���5|�-Z�5�,oi�K-�9�Jy�[��$4x�mF,�1�v^Bhӣ�]�]��wX��ӹ�,�3!ThgQ�]��ީ��`7� ޶�Lp|�<����prO�9�i�����;y��YA.�J��WU�D���13�2����e@B�w+q.�Q˧O7OKHٜ�k.s͗:�6ƺ"���ΐre�w��TH��c�޵O��bN��&���ԅ0:�Q�WC{i��|��e�cs[W{Z�&�jS�R�.���[A_P!E]7�.�n�,�]r��}q0@�qM��U��4�� ڞgu���+���r�5��#CJJy̑1�X�-޹��N�&�5��K��Z���NS��y5����W�cB�v�Ք� ��9���i���nn��N��b�ŋ��;9j���&�x[����q��oKH��/��F���rU��R�c*��J7��U7�CO#��^���T�N��.�g;-��MVe&�;��Q��
!��AY�r�3mK�&S��ٯ���x	3J���ceA��ϑ���&�)�|:�ek�p�S:+^rK�<ݢ,3G���Z������ p� ���rӿ���r��a�R�� �hfH�˺�-���ם�&Ʋ���QtŔ�a�6���<�k4&1҆k���'�"�Rֹ��s����\�zu�3f�#��Rv���}v9wQ;���NUwa}xPOxU�/��T����q����K���YG�h� Z�d`�����ˇ���;\*>lz8j��&���(�ݥ���gvV�g���b3^'�c�dm�,��b���`�붛��ֆ����8�<�e�M\1�%{1V-��7��,ښ#
���NW��'V#�hn^q����١�#@��6euh���YI�����;��t�v��l"�۬k��y�F>��?����9�Xԭ�{�6]����6q���Vl5�R��a��`��鋺B�ĕv�Zؠ��жv��fu�v����^�v�LU�5��P$��	�O,����eھ�u��q��ݗ�vgB�ƀZ��U���9¹*LnG�g��"��x_Q�m/�=E�˔�6zs����3��]�b���[o�/�2v:*��b�;Ŏn�Zh޴��4�	�)Ș4Q]�:�ݵ!d���S�����=ɚ
�C�!��3����>��w�� V�l�5�Z8oe�Ա3HnT��s��d����X��o�
t�В�A�Z��2�S:�}��/��:�]X�`�Z��n�4$u��w�v��^��cu�'$��o-�e�q���\�93�:�b�⊖*��'o�����8��k(se<c�3[�Y��5�t&�)�����~}Y��ٓ8�nJ�SBb�V�o�
�Y���S,�u��]f��2��`��n!3^@�
 -��
��w:�Aa: ��Y�7�vm����m�����\�c��{(��6��ё��
TXkCԋ�ٷ�e�o�v�u�wZ�WD����E���B��r7Ǹ��|�o7.ޠ��f�JlU�e�e�r�+���c��ɤ�OOat�Of��wQ@U+.�Ώ�-�,4��F��P����L�b��ƻ���m����q�Mm���/rtu�������oq0�dKnY����������M�ӝ��՜�	%����� �(�A��q�r�.�{e�<��'�4"�-��'�����&�;&��=HV�� �%��Nŵ��ˆ�ۧK���FkEo�r��H�������7Jɧ'L��T�Ah�w(�����f�C+$�O�q�(�&c��8A���T�i�BȞ!}ֳ)6�wǒ�pS���F��3"J��u�-���S���i���Ldtb�  ᓎ
&�(MG�^%\&v�=�;	�m��"�|�D61\�FNV�,gU�@ED��o.�F�ˮ��5��t��*F�=��EԮ��N��q��W�xډQ��V$���������]�| �AJ��]�;�w�R�Ou!���9�9-��	��re���Ӟ�{��{.��4c�s5��T6�'B�r�8���mLS��u�I��X:�U�r�Τ�����O0K�D #J��X[�����f�)ԝԻ��M�Ndd� a6̛�绍]�P��_wוb��nq-��&CK2jyEPp�w�;��EH�s2��f.F��b�xV1Ҷ[Z��$9Z��ӂɫ[�ŤwU�zS]�u�u�S���D8�ԉi��Z�8��W������g	 !�[��0Viy�]O��#ݔ�_dYO��/L��A7�>]��9H\�,����m��%t����t��#�Z��z��VU�\P����l���d�v��w���������vj����[o0+BRf;�YmɎXp>8�U����%�mm^�|�l�]>2��l�8Ǖ����Uð�TL�z��c?\Q )��*�cy����|Aud�Җ�pE]MK��e�������+`W��)��xf.��b��,R4.���`X��n�nja�n�h�+m�Z��X��4{�GR���䶷���W�D�y�L��Z0L �N^S-eD�Ů�5�x�O,� �7���<#�n�m��'V�ɛ�dk3%�Z��/�$�$@]��]{����H����/�JXw�Aӡ�U�f���3���+K=��Y�G=��V�c�;`�L�3Hې�%w ���l�*	�TL��8V�Ú0���p�Y��6JT�%w��]�Ð]֦(,-�z��м�ژ+��Ȟ��qW4[�V޸U�>����ʑ��X���M��v�@����S˳A�89;*�.�N�V��R�{�'m;�傘Pwtُ�i�"�H��Q��[�]֝x�l����%�
?��-sw��k��G��hz����X�R9nKÍçm��ފ�.m�Kti�Fk�1Y�_l��WJ�� �Kg8������s(��|�^\��5�}���W�}�}��'G�n������wv�qT��Y{�N,�s���x�����e�g��W�p���^��k����B1Kv�dv�M�[*�y�����c2��0������;SJ�s�-�nV�Z2��̵I�@kS��u{��K���V^)�y�z�+�Q��P�����a�*me�L9�m#�68�}����rhn�Zu�쩹n�?�А����W,Jd���Z��ͤ͸���8�*�X5T�G9.e���ɓ�~66�������2��~��'@�Y�WÊ)�ݡ�S����]1|�=<@4Ɣ�X�6��\�|��[ٸif�9��E��WeI{b�h�XQ��.{�N����T�ۜ��_=��u-�R�q�D�ٟ{RM{H��Z�4W��X���yj���E+,�%�:4��Ӳ��f����[���W�'s����JvV�Z:3C��U;��v�QV�#vlg�[Z蹲Y��\{��t���-Z���_2X�W�e9���XKb��0,}��e[՚{,+a�l��K����0��Y���7�wxD�3�.�v��b�7&gTYV6�\�쵮4�#N9�6kBܑ�t*a�u�p��s�؊S�Qq������_,�x�r�c��R�b�І^U��; �]"õ��N
�@T|����BW!0�딖3ݸz�UrZ]�ƯR:w�VVV��1B*�(�+31���� ������&�"k32�2*���,̳,�1�0+	2� �����s���0�3
�3
	��*�̣"��2"��
0,2(�22L��0��&"�2�³�«2��1�p��&��0�33	�,
3����,s#�,B��"�+0�3(�
`�2�2ʲ0�H�33,���"	���i��3 ����̫2*r�(�s2f�0���Ț2"�,̌�&��"�0,2
�s)�33(�� �3,�22*h�#�3*��ċ"�&*�',��l̪*���2&�0�*(�*�1��1�,3&�j��(�,2(�32�3#�*�r�3
�330�� �	�Ț
�"B��2Ȭ2̲�0���"p�"��y�׿���|��nh����uul嚷x�d;�����x��viu��i��8 ��C-����AfҾ9�/~�w�G��V��k��mX��N���������*�U7r�]�ol���_��ӊ�l���<w���!�8�X�~�&;��,R�P����_�!�L��ǭe,&��i�{�����j�=����^V�"&T�<�L� /H����b�^l�������}֟���4��qVd:�)*��g����訞�<�����o@�I�.I�L�D��g�7�U�3����C^uX��d��/�.��;ܝ�m�'z���S�8�����nkK!{�v�c=�X��"�GC�y��L��o�$�|<�ُO�	�G�U��N^os�\gX]�z��e-�gN&_�x�5�l[��p�5�~��\�{V��ƞx�{���u_Gb"-�>\�&UH��y�`��s�w�����Y9�Y���(kʩv1���n!#K����h:�Bs婉�nfz�C��;Ӛ�q�SϾYᕁ�jR���X�N���/7cV�2�C�L�t+lK�:�E��^�!w8���^z�o��]V��1�8����m������I�lb���뒧�_H�ٗ��C��<�V0��*�C����jEЇ-Y]>6�BMQ�3I����/_=�U��8�؆,�V[�ƒ�Wkɜ��%��L�j��{P8�����{x���[Qh	Ʌ^����Ӷ�7�Eg5az�p�0�R���2�A�<x�T'ݨ�Ͳ Aθ&=��VF�Ž��͋��70���C6Ļ�t}E�G�
u!ߒN�$Wz��M���C4��z�*��2{��UglɆ
�T�u§��T�:U� x8M&�H9����e��Ch\���8�.cx��<ޮ�N�c�ʵ/��X����
�Q#B������տh�f��{;;jLx��c�g(Og�TQ�̚Y��ƣ���U��j����E@r(8���;+�i뷼�_���VL�2�A:~�߹Sb<D|�9�6����{���Gᆢ�A�ה�h�hu=��A (�v`*��ye%O��w!�C)�s(�%�4��)>+���� �����o:�։�!���#h1]�}e�������8u�q�em�A*g�M���8�{��{�����LΡ�s�
�%�p���S3���<�?�v4x�=�+9�N��Y𞜉*��TS��N_��}],iƗ��֍�M@^g�K^��h����Һ���v������1��=�T��ýJ*/��\�Y��;� *c9�=��)fIvM'a����X5w+��t�5Oe�b��R�*�ž�ORՂ���j�I���-2V�C:�1�u]ݕ�:��#v2rFnW
y��2�ݙۨ��NX�c�����a�=[�Oǆ�r�G�	� �y� �Nb{EÚXx�%��.�����#���zU�aL�!���W�$=�G�p!���F����+�lF�o��W{[#��]cD��h<��9�qV�X�������ƶW��ﭩ�����b��hז����i������B��EWo�o�&V���At�
��x���X�_���ŏ���m�q��`����LW�ւ�}�e�Wz9Ww�/ .�� ��eK���*�2���e�yF��2�"���'W����	
Ҿ'	��Uq��y���Ss-qݚ�W���N$eNS�>��DQz.�>��@c>�i���0���9��|�ϡ�k��g��+jX�~2�˞0�କ9o<��	ư'R颦Y�n�o�K��nxy��B������]]tUX�1���K���j�W���e�����.���h���y_)����<3�,��@*��w��
�<�x�U��ꖳM; E�,}��B�>�ܯ���Ǽ�SLK>iM��]W��M�2����^���ԣ��{stj���t�2x��0����2�\�VӲ�e�3u�QwrU8.��OLŬ^C�S�m�[yS�J�7��*3�s)�a.�P�
�a���K1����8���������yo���*���},�W�lWYB���W��r��y��#��i� б�eyd��q���ȏ���M2��%�J��k���K�V���(����'��O%�{]��=�ҵ����"M8`p]����+�S�KBa�y� }C*u�I�#R��+h9�ʂ�oR����d��{�s +�u9V����O-Tb�hz]��7����4.�,w�nyd4��U����3��]�o�xF�i�IXjuC'��-�/Ӡ�|���։U�-���+�%%��*�����X=�����e@En	�xi�O޴m���qg����1BǆRVY�;��\0�<�T���R&�n��1e�ק�拉	�n���%�s��9S���6*³e����C)r�\�i;�Tf�^�)�����L0U�2�Ŕؗ<`�g|eg��ʼF�Qg�g�¢W{�R���%������m��!3��O���2z�N�g�ԧj�Y�D,zг���uV��X��X���*�(Y-T��Y������\ȍ� ����0�pm�\�"�9�s�RTun�ڎC��pxH�͘`[r��`��v&rEu�Ua�@��A���`N�n�R��W�ιo�ټq�r6��\t+ۖpwu��Z^�غ�
�� ԗr���%=�T�"/��h���_8�8��i	�ݐ��F�A��*�sD�W/��ª{�o�	Lފ��/��_��a�Oq;��E��}b����>������8�<���]B�z���r.�o.���g�I��9/�u�[�ϸ��VMv�rb�4��s}��s{�\�oeW[�ϥ�6���H��H����
� ���pJ�ï���������Z2 ���Ӯ�bI�/�&xO��U��R��������5s�}e��v7����	"���J@���Mݬ�Ys��x���fz�Q��n 2:�e�U�B���6��r�:C�Op�;��y�V�';�8�J�ʟ[�yO;���D���[|�w��G�ړ�:����z�j-��vΎ󽊃�ڟG�*�V��^��|��������ꇌŜXa+�;P�Cry4z�ԡ�_>u'>픃��4j϶����M��k�{ybP?l6�)�c.���Jn�<y�Y��:�e�{��65�%��A�'�8��ņ N/&ֽ�����s�5���Ӭ}��^y������y<x���6�����Q���y�v[�+��V_��Q�6�����a}���R~��O��-˙޳�������'�=��w��\��v�2��\Y�:s�^�s�/&���׺ܔ9ۑ��:�����cŎ�r�ڄ���z�.t�&I��OZ�!e��9�wp�>y
c�EG��;���A*xOmb���{肒M��]���wt�=�'ʊt<]�Q:�\�G�t�>�׃I��eL|���ٛ{W)og��뎻D5�����5�k���{q][�v�^z7����3.\��Ι������7��;��K��T��|�Q[��Jw�.<}0�,Y½ғ��?9��r�ަ���)<ҍoxp޻��U�Ȇ�j���и/y褆�u�F����?1�#��vS1nIROP��*x;�;j�������;��#�4p��>����M��l>�ԵX6��p�*�G��O�AN�Fp�v�U�ހ(��-rh]Cm���Y߆�owV>֗�aiN�l�e��hCA�hQ�����yÏ?I�]`)��� ��^S��
Ԏ���׺� m��	_f�OU�S�F���f��%O������ю��ǧ��R��wZx�����N��%��3O?^U�����I^́7&Z���ݒ�	ZՁ*��M�K�)�.��e�	�mL��X�J��]����h�C|ߺZ{�۳_'��9C��:_9�:Vߕ��1���N�x�w�xF���۽)��Y��uJ�}���8É�oOj��_K���w���7~kN���}GG���^��R��"����y2n�����9N+T<����I�?V�+��J��Q�vt���%e늋�0h�ݳd�����8o�S��Vy,��6�h�����N��P������λ��EN�NO<��$����wl��y�X�gŏ*�����s��Ձ��Y�_e��b��e��	X�pT�$s�}A�����M6�(m�	ǭ��WDnVE3��Y� �@]�1�1��׺Ȃ8��u�n�hKW��j	���U� cu�rL��8���Z��x�b�H*3O,w�/f0���W9W�K�ۤ�I�Z�lN{�l�:�w����\=���U��C�Y�ݓ�u"�vєڝ]L�rΛ�u�]>�z�l=gMdֻ�9�N� �7��63�:����94��U��U}|��?g���zp4׵��9�y�?
���_c�>Sl��.W;~2���������w�i�꾶�����|z�c������F�_���4�T�h�� _?���h��"���U�z�9�O=�<unWH���*�M���t�q�ھ���澓��ˡ��y���Wd�ѷ��p��'&��-�5�YE�%�u_J�=��>�����)�[���p[U {I���յ��ʎ��B�&���=���B�:����\�ۗmʥ�.��à�g=������E�ݾOY)ױ���_by����(�xv�B��-���t��i��i�d<�?VD�1�]N�)0c���%E�_bv��?-��ꎧY[�8��n�P9[��ᔷe.r,��+�뫎���04�g)V�:��{��u妯㰕������\�t��Υ��2�	ŋ1�|M��Ч#���	G���S�td��L<���߃�%��1b�c/N�Z�B�F�.�}D��*<��B�m�u��)�y�ʭ��{{�b���G��~�vۨخ}_K\���ﲥU���^��
�9�}�:�@򢽘y
�{�������{N[�O�*u'��2�\T\O�y�8�m��(K���O����J7R�t����h�[G�C���S󊋝1�=��p����ϊZ&��1�3s��N��h�ρ��[���wmI�&�B\�;^�j �쎮䞹ܭ��~��úz����O5���Ty��{�o���ϬS{�o���f���Qly ~�m����Q��]�a��[��}�JMW1���kw��o%*��..�xӱ[�<��Ohh�OW(Bݼ{��3�Ώ_��<���s:佻��T݊Z�
W��{<�_{8n
4�=��_�K:��u���������I<����<%e�����{␞�Lu���|�	���bސj6�Uq�n�=*�mr���|��}�Ҟ����A[���4�N�U� +�T:d��BO��֫WV��Z��y(I_�rh��w�(ڷR��}�^���b�Bp�Au�j�<Zrp}�:(��FW0=Z��,�v�/og`�;ۮ�\��Wm9�[��P׫�݁�Β�~��Vr<&�{qyNV�o�ܻʬ������ V�����iߐ�ʂp�G��s��ƺ[�>U$���^Uy�8V�o˫�#�_	��.���/���ҽ�^����vz/��*��?�ޛk��'������v���}��+�籅Y<�eI�U�b�g����E�v�Yt��J\��1;}Ƕ�Rz�l��rG/6��#�����ïN/)3nq��fsqL���N��=�z��UY���������=z;c?'�~mt��M��_�
S���NN�	+�����:P� 7�|���p�̾�k���uC�4}mQ;�뮻�@p�=YY�w�����)��Qw��fs~��ڢ|�����b�w��0�x��jf��%�K�f��:���:Bwt�L���EG{�x^)s4�j�Kuqx(Mq�8��2G�Uv��pCJ�ge����a�\]��@7JkF��2fСX���6�^Z�I�o4�@��&��s{3�C�Õ�h�<v���g��ZyMI��ѳ��iyw�p ����y��B�"���氵E&��,�d[gV6����$,��=R�����2/�ΫtW�櫃{�+(B���٥%j�ӳ!WC2]�#��^g>n�������qqɀ4�u��\~���f�u5+�0]�m��<"v�|ǰY�_�,W����k �L}��Zsu	-�1��,�/Ty���2��l��8�k����uw[�<f�36�i��[��Q@Ax�4�o�q�-���=���UaԊ��̿�з+3�����EU�o�E�܅V8/eo­�]j��S��38�xB��+B�M(jIN@q��Q�7�SyR�h!�p7�2VΐS���,]�u53���u�HRŁҏi�8�]�o*�SX���h�W���^�*%yt�����2�t��H��/���N�z<�n�wB����ţ ́����y:0ww:��{���S�GoH�wڸ-�z�T�4z�&�]%;��M���c�D}4��U9�j�w`�f�2�}��T�/��f����0-�ɻw]��K�)���s9�k��\����Z�8#�"H�����5W���\��,V�m��R��o^i��{�AnG�{� ڙ�YrgLP+��
Se��Ukd���b��&%>S��
61��+h�br6��mf��sr�{G@�Y��=Z�\�����T��ǁ�]Km��=Rũ);[��t�]�g���M���;�(��v^墱.���R��Zy|�@iKǉs�ME��m�F�y��9s��F��A`�2oI{�_&2�'%���6.����C>;jL�?F�Mv�J�I�n����n�ǯNck�ٝ�u�eSWvΧE�S�|�����u]t�a��x�^�{�ۮP|��[����-NYi��\�T��ݯ����s����U�݃���t
�C����ӛ�F6��:��6�*X�u>zv�S�R�z����ǧ��t��`��r�q*�h��vp� ��(���k�7,Q]������cT]� ��-J̅�G!�y�l���-�V�ז$U��;��nK\{v=�OJ�-0+#\VZ]��ޞ����J���_rR�޷Fd����!�w�U0f��������Z�8&&T��KL�f.�Kw��+`��lu�|�%��LUc��B>�B���څum^�0�"�u6������D=�Ҹ;de�LuN�d-���-�\�Q'f%{��on���5�wz�Kr�
J� )�%o�֭��s{:f�|ČG�B\9|#\-7|l��<��ch�I�,���̭���(�x2�u�����_`:ۡ�How�����{�}�VXٙf�نM�dU3��D�FX`Y�QeQM�EQ4A�dEVfQ�e�XT�c�e$3UYa8FE4�f4QUL�TASAT�aD�fA�f3DAI�eRœ�e�`e���U�T�adQ�d�eE9cME�ٕ�a0MfcdUfUMSI�9�4і9�I��NSTMS���FXS�fPU�`Q@A�6`�Y`VXM�dTVe��f5YcID�LUS��fD�&U��a�4��TTń�U���EU��ffa���e��fQfAU�UUSE4�U�DD�D�9DE�1LADffTRDf8UD�AV`eE�Y�6eI�KDY�Y�NYM���Qed@�=Os�9�r�#�Զ�ۻ�o<QΏ2Ss(b ���
|L��� ��/F�.�!���%��c�{P[�o'@���;���4=����A�l~�s�d��D6�����>��k��w����=��M�r��k�|�:5��<W5��q���.X�^�z5�yO�g]�^�K�}�Ϝ�Z�p��<�/uu�n5�"�������4�n����P=�=9{t���I��%�v3�)���yNAU�C=8sdwsյ��)�@k0�־��Y�c�{\��������eε����<�'t^O����&�KQ�@3��G�ɬ�SfN�iZ����xU�)�7�V��앓@�C�H�')� ��G��u}�Z�v{&tU�%'��|��M�����nU1�>�7�vո5}�S��_X�� ��Iͧ�Jv�+���ݬ��庝eS�Mr��c�*s�7מ�q��"V�g#<�2{+�#x��H�yoݚ���R��r/��������{ƕ�7r	E4(�*]�O�Y1ݘ�zb':X�ԕv��xW�-���I7x{�:j����c�)�x��b�2y�	��X�����V��b3/�f��-� U�0��:���E�tz�� !Ë��1����c��d�!�X�[�h�y��;y�x�k�UپU���H�Q�vt���U��0�U��n��4���9��n��>ޝ"����;}�b+~x��y����|�z۩(s��&9ȸ�}�?c�oz������ڣ�h��@�
F��o��Z/�x�r�;*!:9��Ӈ�4�(m�	 >~Y~c�w�C��J�z�^�Fp����OC��ny̕�y����4�^��=�[�p@��zED�W���~ʦq�N�^ֶ��6���}y�^E���,^��C�`k�.�O/5�9��;}�>�}efO2:乞�K%���اޚ��]r� �ϑ�.�o�~}�l���<{����D_��Je��"�^��v��g��U��p3ˡ�q�ՉI�/��S:�*{�eKQ�6�@}Z��S*_� ?>n����Y��H����Զ��K�,KP��{�x�zẒu����3)>t<7p����p������<����������QY��79���zQRa�lF��N�q
��Ut�9\Bӛ':�]a�,��`.��#,�2;W�:�o-o�-;.Rk��])�� ��y�6�@�[NW���5	7��~4 ^^��g�h���fL�}r,^O{�fWt��n:T�=��OS	�4�-͝+��ճ䯕<m{9\�*��=�SM
��B�w^�ܑ�񽑏^N�*�Պ����;]������zv�~�����*\Pf����gzfE[�A���k��M~�H?e�!y�Ƌ��w����Ÿ��[��ō�羟'�ܧ��x[T}s��9>�����^���-��]�g׮"�y\c�8�o�^~_%xS>�*�;}��y���<���[�����:@z9`q�,M���(H(KW=ع>��6�����E��k�v/�WZ��z$�}4I�`�Ku�Ƅ����e��E�w߼����6��ۡ����k�y��|��a�w���/�X���̾���f6��<�X���ۋ\[J�7�*�UbmO$���wv�y��7�s���|ws����˝�@b�s��
��ځ[0��E�%m �e.�me�>md���|d�\��R;��S+��G_�b=�oNZ��]�f��rq��oyg�oc������;�g�\_渿&�G�G��n%�^��\����q���*��/*g$�6E-�����1��ʾ�Z�~��'����9���2Lb�c����-���j�'���
��Z#�!U6�w3$=u�U�8��[�nuO�g��Ӭ�:��vܓ�_�I��_����	W�u1;�c'���b��j��ٹ���4�w�URdy��t0yw�V�u3�n��q�X��G��M\U�U���}���������w)���w��.�����{����%r2O���vl����^���}���\:�􎣝�GR�!�7��ܾ�I��Д>K��Z?J�O��˩]����`nW���O��SǾ�܇�w�����:�_{�_�y�>>ם�cr�9��}� ��z9+��~h仂��0;�p�9��Д>���?+�z��.]���G��y'!z��g\��g�ϻֹ�^}�?}������}��O�x}��R�'��u��:��V��{��}��r
G�7��q�?�O��g �1��_Ozװ���<�I�}�q�w���^�pζs�/���ν�=^K�d�H��w��;����=��������%��p^���zyJ�=�oG%�dG|��9/����!ܾK��y����,��{2�E��Sz���s���-N�-���K$�U,']6HS㜡��me��Ie�Ζr�O�R��:�][x��*Cnt�k���btW�f�s���� IgY�&�1�͓jw���>�2����$�%ј�����O���w�;�P�_$;��!Ծ�5�{;���X�W���u��y�>�Y�w/G�i}�r�2{����:5�<��{����K��:�=�F���Q�^�j�}�V>�����d����ц���H~Op~���z��~��������pR�}��r^AK��hrù��ߺp�Oz;�=�=���^������;�/��-?}�W������{�G�>_K�~�K�.�u��=��f���M�ӬS��.�a�_`�t�����������������?p�����������r��r8w�)��'7�/�y'�֞I��w/��Ҿ^��δ���:5֗!��NK���f!��qְԯ�n>����g:����:�o�{���}�����y+��{��FHu�t�n^{��ϴ�K�?�Gװ�^���4����^���w>��:�d���b�>�v�?A��
Oxh{.�V����y��z}UV��b�U��}��Ԟƥyy��%����w/;�縇��7޽���z����9n��v��u/:��I��=���ߺ�������}���u��(u� �~�����ON��yI�b����}//e;w��=���ߴ�_dw��z���懓ԿI�ï�����3vy�|���u�{��^wނ�����P=���y/�`C�~�����?={��]�F��nL���w��䯢
��~C�>���o��������2=��w�^w������0}���4��Z�y/\�AJ������pܙ/ђ���9/߰����_c�~�=�%���ҕ�=I��ٮ~�������?�y�^y}�w}��R9?��w���ݛ���>�vs�L����O[���ΰԯ!��z\����nL���b�_e��:��n��ތѾ�y����@��(y�	�3Z�ډ�;�Âx�	�ڞ���kY^�����c��V����I��}�s
(�R-k���Q��6s��4R)�����*Wo5W�u˘	1��G��ו���Y8)0�;4�����_5c�1��m�W�˓ղ������ϵ���?_K�A�=ޔ��Ԟ�����=��rNH�9�C�(Ow�%��
~�	C�;���w�w���]�>�����|9�~��石�>�\6w�|_�>_G�7/ҟ��Ow��'!��C��/ ����FI�����_�ޞC�(N��>C�}���`�>G�[��W߇�_fC��/s���~�ֺ�<��.Z����-'w��:u���w���'R�S�uޏ#����t��Ի��h_ ��AJ�zw��q��o��ܾ�I��~��﷝��u�^޼�=��{}ןy�>��^=���w/�b��>��{�G��z����g��x�I���z=���<����/�u/ �L��B�����_�`�ȝk˙��B�O9�5�kθw/��N}��M���>szC�~�����>Hy�K�w#��O��r�FG�9&�|i?C�!U[���
���
�q�Wd˽zb���W������������F�߸���r�_o!��4��>\�%���~�_�n�b�O�y�r�FG���AT}���00xW�7q�o���!�
�i2��2zw��<����rz��f�wr?o��$��_���W�?b伐����C���գ�>�
Yu��=�?~�)8���+��?`n
}fA�~����49'%�d���	���7��b���ގK��~�ǟZW��z�Z]��z5֟�������O�	����^�w��d���y��?K���������ҿ]�I�w!ӿt9'%����y�;��q��}������^�����
���럷%��{-�����%|����>���2�I��=���22G�w���/�Z�I�w�)����]���<��S to�y{_}+ﮇ�(=�x�ٖ�Y�^B��M��5�Y���x�]ܳ�_��̉3S>����N\6�3���e]����*�X���L�q���#�Ó�0_SK'v�nِrފ�������ٵ�J��ñ�N0�-u0�p=�룂V~)]�I�=J*l���3���x���:�u�~�@u~��?G~�?O����2W��o�� �t{��d;����w/#�F+�;��`}?�w=}�A����/]�1U^S>�g�~�����C�=���u��_{�:��^=�__KܽC��4��K�?��w�~���}�w�}ir
G��K����ܿGF�Gp��{��X����L���\���>��{��}翺�ܻ��p�����n�~�ԾH�w�h�I�o9��u/����z�u/\�AB�����d.�sp�FK�������߿]���^g���|�|������.K�y�'��w'9愯e����^\����;��v��<��9��?C����{/:����¾ڙu��|M�:D�����7֢�{Ρ�{��{��w~��b?Hk�t^K�y�sBV��N�}��rroI�]��4~�pP�s�L�p�U�����|��_�¦[%u�E�t����g���W�{�'${��wP5��d��u%ܧ�]�;���w���C�����k��9�ǓJ��K�����fW���6s����~<���Z������2��)<��~�������+��t��]������^�#��:�r�����z�p����:��v��\����>�}���t~���y�>�^��ޠ�r9�4y/ѐ;�=C�|����hJOe�yּ��w�����=^K�<5��^�G]�u�KU�������j����J�gW����'��s�4/p{'G7��R>O^oO!��\�Op�_}��|�K�����^Kט>Y/��:u��y/QӬ���c�+O(vn�[7z����O{��7#������
^��h`�A]��@�Iѭ��u+���ޞC��N����~��í� =�۽���|��y����q����u��ם��s�uա�_\��L\/NK����()�`��&+��'������W>V�]�~����v�����o�3ez`R���� *��@R��p@6tvW2 WyzzvCW˫^�ur�ڽ�Һ$q�p�WògNO�*�H����e�}�=���7���e��n����L�e�?�`rs���O����������4�n^FF��w'$���r:�ܝ��<�~b=�7/%�����W�ퟻ�5���gz׷����uϾ;���pr_$;���u'�q5�y����~����br
G�Z���N���d;�q��1��3xr�Wrp޴r^y�����o�k���|�~�￭}߽�Ww��;�K�_n�]hra?f'���$�Aֱ���f�}���9#����Mù�����y/<���L��_k���˝��{����޶wu+ܜ3�v��{���~�ZL��o��$��by.���'�r�F�R?C���'#���E��^���}T�V��Z��F�� ���N_e��}����;׷��^�����{��|�H�=���hr��o��&��>�%���	���Ѡ���}P}3g��q{nw�?=x����^G�?O�i7.��;kA仗��7�����[��z������^���#�u/N�����o�� �tWb����(��/���
��_��c��޸P�/��ъ�&��o���o�M��1O�kF�{����u/�=}��!��<:旑ԿI�;:��C�δ��ל��g9����s����mr
��p�?NC�X��]�ï؎��}��J�=>�JW�������ܝ����9+���K�=���4��p����۔�;P+�#���~�'~�=�����|�����d.��Ð�9/�X;��y~�?b;��?~���^K�<���/Pu�~����+�¾����C�����9d���8�/աM	��4���=��<��zy֏Ҽ��}�r2G���Z_��?:�ܾ���Ԝ�r������ܞw*������*���W���ݡn[��f*��.�GfU�֧Q|�4�mm��G��]�0�3,�	�6�ZH��O�mw��;����U �)P�t^
Z�7yҧ.+�A�G*m����v�G�����<���־	�ǂ<��d�h��tF�t�}���gm�Ӗ�,���UUW��S���+Z���|E�3��H�:7�K�)��r�'�sBP�/��Z?J�N��K�r���-/;�?�ܯWq��'R�S�j��K����5?ߟZ����_A_A_~����c�w}�H�&A׻��)\�����w!Ѿh<�p�9o�Д>���4�%����w+���=�K�����畏�uk��6�\��t��A_}�W�WRnG�]��z��9�q#�������9�ÐR=��o��q�=���>NA��i%�_g����n��+Ԃ?�?�[�����}Z,}����_�b=ۗ���'�>F磼��㯴{=K��5�/�r^A[?{�{��sx�?J�>����w�3p��k�]Ի�-W�?��dy?WI���P}�<;�^é|���,����Z�=�K�t�J�?��9 }޲��
_��������t���y�z��.ϻ�p���>�ٯz�ܿ�dx������:旒�]:�K��!�����;������tk��&G�7+�ޭ%��y����G~u~���M��WNկ���i��_X��}_���7��N�ގK��{��=���~�K�.�֗$�R���y&���)�~�qְԯ�r:?`n
G���{�>�{�x^��}�}�og�k���!ǽ�r��r:7��y'�{���^Iٽi�[�r����_�֗r?GF���>�Py9.懷1`仍���Ǉ��מw��>�~��^��W�>��7�}��˸�wK�p<y���y';���y/P����=��ϭ#��^�u��_c��\��M��,���]o|��|��������A�����b����%}���'ѩ_�u��~���0;��y���=���׷��/R�u��p��|л����w��\:�o�܉P����Y�̩��g�.z�d�J��^X�՝ h�oc���E���J��{��g�w[�-�÷�����WbQ6����g��9��HGL�=O.������EG��/��ڱ�A5o9��Xo��jBdO2�X�����~�u���l��}��2GR������}�%����>�p�=:0_��~z��1]���}//%=w��=�����<���9n^��C���~�������go��k�_h��p�������9ނ���և �u�n������;���F#�}��{��]�N��nL���sxrW�py�[ߛ�V��<�>�d����������3u�h�������/�Oaδ �^�w��w������2_�%�w�~����Gr����y.��׶��{�g#�,��l���}� �}��zc�r}��9��9+�Xj]��9��j_ �f��9��s��y[�K���ۓ%���b�_e��<���~�a}���?q�|��}Z*���������«�sJV��N��u�\���ÒrGQ��i��Bo����)��������p��.u�������}/��\鸙���V�W�}�UQ}���
�⛗�������ɸ|~�H}=K�;��rW#$�y���������Bo����2O~愡����\��ܵկV�n5܏�����C����U5|B��i:��q�NJ�yw�Ի��<�K�;������]�m���9'G���)\��{��w)�?w{���U�~���M���5����L}X>�E�~�`y����_|�K�p�/#$z�������<����M��~�G�Լ���׺_��^Av~����.���_�fc>�_�3�F����X)�������]�Js�h;���{7�y/��}߿��C��,�������r��X�W���NI�:��~�pP�w���3;��/wWI<���X�c�*��Gp�oG'�^���z9.��{<���~��Ǯi$|��.K�gx?Y/�7N�O'������|��=E/;#�x-�Բ�pfHٺ��k�r�Z�9���l#��E�W�0ۨWi�*��V.9��B�۹�����A$��F��Ӗh��I�*�"�!����qb"���ꍃ"����(���0�B��ɉv�vi����]��:�K7k�9ww{�%ɏ�(��*��*N���	G�q�_K�a)�'H��qj���kEِ���)va;��͐�+��8Ne>w˥<
��-+
�F�q$P����g
��jf��o�PU��擇���59��W'Ǎ�v����*D_n�=�p���E������T�Ï�T��y�+���޽�68��(Ng6��r����3��r��WTV�	��#�.�g]��)֍���NJkz��7K�E�=�\:��5��) 7h��8�hR�g%��xVd��֙������B�룼�����K篍e=@p)bv�)+S$Nܶ�R[SiӬT�P��?r��3a�S����$U�z1�����"X%�֭;-]v&K@l���ܗ:��]\�ѯ-r�����)վ��s1�[�&��1ԡ�w�����g5�1g˷�H�.�n���c�3+U�'nWb6��9qJ���2��]�Ķ^�lF��nj��{n��֮���-�1�V8 d�xb��ǘw�wWb|�9�)�z�F&7����:�T��?��A�+��+8j�g\)�{�;��
�W�!����{�37T��.���Α�yV���%'}�WIw&�2H���:=56X�{�'<�eө���_V��󴳧7���u��`�Ys�D��Y;����:t�ԇ8k+�JL��p�%,ðZ{.��߅�E!AW.ʫ���6�s2�:��F�������5����=ܓL{fn�q�K��C���v�(t�)����B�%*"�jTK�v���!)]�uA�+9ݝ�V�U�Eq*�
��G�׵ح��k��dGi\�.�r<<9]��w2Ű�]"c��
7�GY]αoaQ�;S2s�}gmŊ��du:�v���l�B�Ѯ"O!2���i�5�6���|�JNˡ�'���ò�k�B��N������bj������4���m�Ց]tCb.��Zch9B�o{Uq[�ֺ��u���%g-2gD�='r���H�n>op��z�f(10M�nr7f���f�f[��tw��%��8lg��+�e�w����)�ێP�_o*sK\϶�!OU۷\���K��n�[;�����A���4��<�M��8�F-ʈ���ew*쥋�em�|#n�K����R��C5�6���##ct�1�[J���m�ר���@�#��mei�2�'�p��S��xg^P��o&���bQ�o���Ǉ{��kD��ػ�
e��;uȱ�s+�i�Xi(����C�)>���f��m0lu�7b`�ZU��M���v3_�#���Q�C�T�j�*�"��"*���&j�j��#1ʩ��)�'�*
�1��1�j(��j�*rlr��1��ʠ�3*&(�h*��*����h���c#(�̚�2fs0(��	ƪ���Ī�������)32�"*��J�)�&��&��&ʋ0�����*JB���
������,j�bj���)��# 2JR ��j�0�2�(�K3*&�!�X��f��"Z�	�,�$��rh�������`�)������j"�$ʚ���j2��(���� ̰²r,�b�)J�&�0̨�+0�*�̱�,��`���*�*�1��j�`�331�h�#, *�\���(���L�%�
#
�&�&��0Ƭ�� ��f���2#*r))�32���
�����(�b���j�*JiJj�b�'%�!�'������2�h31��)���1)��,���0�ʀ���������v'u;��6��C���w{W�R��8>�c�l�R�qr��j�q��W�	@.��}$q����z�����}��w�}3���h
��ߜh��~���7�!�^FN��w ����#�9��r]�H��kp���|��.�|�5֗%��=���;��x����o?-���sǍ��}X>C���ԯpru�P������y!��9&��d�o�	������د$�7������9��|��������{�/��_�V�5��~�No�����A�d�C��'�j_�#!|����J�s_i7.�$:ߺ�������y;Ǟ�?������{��q�T5).������~��A_~[u�
������~�>�!����K��XjG�w~��B�u����~b��փ�w// ���S xkγ�7����m��g�0}���_~κ�����K���(��uc��k�����ɠ]w+6�[��$z�ӻ�������K~����P#]J_�����X����ɚ����ָ��*����s�>����1n}$]y�Ȕ�w�@k%?f��_xs���--,v[O���ԫ��ʖ��m�UH/kä�	b;��ӆ�>��ٚ�'�nv�E��$�_-^��)����!�J@���88�:�����':�ǵ�+�N�D�{o-N^���m˿�r�gA]�f�5�Io��h��3������*��{�)�����㫼>���vUdI��W��)����f����
��p�$uM�W@�ڏ-��CC:Jv_pKe��吲����l�\����ԕ5{S�_�wZ:�i����]�M�K3���{��  >�:x�wh~*ev^�\ן��YW<�t�I~|�/;pj�O.A������h�M�y�s�����NA>�� ��bu��u���!�ǹ ��=�>��p��ܝ�ΝS3�uޒc�� ��,�M(r���Ε
���,�J}�O>����/�%e^����1�¬�v��O۸�=��w�����3�252��T�{T ����!h�<oA��"�y�?g�9�#	WM�:dSq�Z�ӂ�J|./���3�u���Wx6󊋝;�|ߕ�,���q��Wb����QtTP����z�����r����Ix�VNCb�9,�����t���j?X]]a��� �����p<�ڂ��^{p�ݭ�e��1��|�I��\��T�z��n����\�l���rWn�Sщ�������R���;�ѩ�x���Չo��\�p��[r@wp�n�JȘ��z��5C�����u$S6����7�>qM��_�<�����o����wu!O�C Ӧ��1̨��]��u����=ΒV��N�(�h0{����_L��˷�;ʏ�u����Y��l�����_U}��U~�<乞}���ٹ�k���v���L�)^)U7|t߳�6�����w&��ޡ�R��]���~x6x���/s��=��o=�m��^�M�j�[��eu��
��Z�wZ���:��ͮŖ��Nt��^����s
c�9]��I6#0u�Dú�Ŋr�[����{Os��F���duHgH}�����zWJ��V�vk�ڙe�՗"}��ɾ�TI�~S7o�j��tЫ\�t�'<�g�+o�/E]�{iq7Į<���J�M^�y�����N[�����y=�/�y��=�E�\�/+Μ1�+m�s٧�^���K��磣��q{�0<������ҏ�en�߽����|��ؗ�_��).��]�pqA�!�a�Q�U��h�������`d����T�5���0���H2e���^�҅��x��`p�x��"X'�iÕ�uf�vV�SrǕ9Q2ż���:�
�pcu��o6��������+�su��HN_�W!�%�\B�]mQ�L�5��."_2�+]1?8r���B,k�`U�	ل��wt拓���M�i?����bAO�v�Qs�Pr{*o{��E���j�.��J��F�c��\��{���hpLSs�S3��N���Clx:��F��ׂݜs2��gNk�9{qQ��{�o�	s;bs�u8=U׾�n�fp<���f�L��P
���Ps<�*��L��zw]<�ş'\��`�])�ۃv{%�r�@�>~!�<�l��+\>JI�>��.>�{�eĳ6R�]yS9*yN�F�X��<�{kak��:,z�i�u�=���5~Sֽ�L��$]Y�S�e;hZ���Z����{&�h��j��_Ken�w�{#�m�T����Tˋ�k��Ue��r�2L��u��d��>�f7�.��R'NS�mWJ��oH��
��kkX�˜����^�v��Z��#��=����w@1��qҧ<� ��g��u���y����U��gq�)C����mM^۩��Mq�R�k�V�v�1�O'&���	}t�%�퐜��0ђo��q�����;�u[e%������2�����:�Z��WOv�ۑ�0�	�z�Xelׁrf��������뽇�Δ��շgy�}���TfybwT���n�O�uk�/`�bŤ��?O6���J�E�؈�^TF��|˪����Wf�=��R�Vzf��9-O�ǻ&{y�ڥ;��<��>��@�^�G�������.ݮ	D��Vwe5^�NuQqfs�s���)�*�2���KZ�������)�����D��}]� ��q��9�t����px��jn%�;v��6���ؽ�r�&C+l8:�������t�oN�p��V�=�f�mnY��ΉO�����A���֮_lm=zh�2m���z��x&�xr���<�u��;��:}}|��~a9�m��PZ�3�9$����%^�b���Ɨ�0mӱG����s����[3�潷�?x����λ�7>���36M䢒e��9'��GxAty��}v-�On�o��O�9����G��6�kr�˄?�*��n�c������9�^,Q�`����S[�q��|4�WǬ�#F�����E��]ѱJvn��f`�H�I��9�vO9VH����pr�z쎣���
ٔ�����ꯪ�_������=�����cS����<�Z�1/�REןTȗ�2��.��$�0�޽l��{���j�o��Z�V���d�CorA{J������L���	M��^��-���5ګf�j��)��vG#��gjԷmz�.��8w�ǥg�]Y)��� �[S��U�k3���']����/3 �_�66ϷبO�{�GOB��Z�k��sʹ�K�����_�;w-I���F�|�W����y��P�o{�S��et��/E�`ƾ��_��Ս����ʏ/����fs6��y����,-���9^U�_Oc��9ܾ�ت���nQ�Vlٲ�[Ckw���^�c��۔s�S�苋�<�v�?n�$qZ���'G�I��j�4�0�/��Q�x=��7�X�oJ�@fv��X7�nt�[i[���� �¯�G�]gQx:W����Ӻ��B��-��]������N�X+h��ڶ��w�H�ŷƦ���j��gy�[śZt��;�/FeA=�.7�h�4=�Ŕ����7��ɂ�S;Q#�4HjZX���n�Ŕ��M�뮒��=fK���A!����#�=�+�%�˶ng�ﾯ���l�@μŌ{q�,�˚��c�4zڢv/�WZ��{뚱�)\�r1������S&�g{��j�m�PC�~�D�|a�4R�����[��=�ｓnpU7�o��	s7��7�>���Cmأ[��V���CK�8�u��"���o׏�(�˥��[�1�7ѩ�x�H����<]:Tm/Vn�{w��Ir���*(8Y�|k��pi���^v;^U]�g{�"떦��.���&!Tw�7b��r�kX��j�������V�O����;�oV������;a�[�l��.��yL�4�X�����[>��P���fi�9�ή�ךA/'��f�I]�I��O�]T@0��Fr�H�l��I�&Mr�iu�~]|�F�s=��w�ߤN�9OB�^�j� ��ڙ�d83<�c�z��4�ֿn����\�o�:��Bߣ�T瞌��o�ұ|��M���c�X+�(Rk� ���a�u�a�ԗ�Iġ�դ��3׺��}��EH�Z<PX��w�ڋ��B���:��10�ڸ��5e��u����4�����j�Ur�De���
�}	w0��ü��W�q΅�I8]М(^�q��������W�U�ܔ������[�~�5eb�=q߽n��EZ�y|�0�'��T��|����}�N�8<�>�Z�x�a�$_���ڝe_�Jϯr*�/=�R]��FN��h�fX�rv�?kZs�{�ڪ; �R��'t�x<ޕ'��5c�������|w=v6wm���.�&5��|U�(��gR�`.r�]��ݧ�U�n�O\t���M�q\��ׄ~��p)ó�)R�W�8�����d�_S���D��xK��Lfs~��ڪ�|�r.�M2��G���y绘U��d_\�_l'�&��p�;b�9�T��O:���ɪx�s����@<�/����<|�����?e3�=���y.��yXN1)[�F�y-�^�L�5�%]|��K�pw��r��n@/���Ē�ӱ��l���I�K~�c�z�ީK�_1\���y��Iu�+=b�/|<lu�6Z���[����t��~�J#Y^��xǾ��ﻗ���S���ᮡoc�U��젖h�MЁ�i�V���ҩA��}0�����΅Z�3gJ�=ؤ��r����V�Gr��=�'�'ύ�*+v�-v�Ƈ�A4��1~��������������cןK^������E/~�;�W�ާH�)�����]ܙ��v���6��44��O	.u��Ϥ��rj�e��4��/u�[�5/}|�z|s���W�z��K��r�:T�=�ҽ�u�u�?���_��m�ݾ]�,�S/��t��'�wr�]��.��tn�F��۾�աoFؼ�����Ջ�k]l�VT�:=-�����m�WM����\r�"��z�it�Z�r��{�i�t�=͞Akڣ�J�ث��5I��o����	ǭ�oN7�������iw�yg�u�*kI�z�ǐwu�^�'\Ι��7��:<G���ޚ����/��ˊ��xD���$Y���|�̡ѰOp݆1.���t��pw�\E�3�~���/?S�}Ց^)���{��[G��:�����߄��{G{�}�o�f��n<&���Ȓ��z�t��2.�Z�*9.����\�%:�pKѲ��;NuQ�-m��X��w%������YاU�dyZ�[�칪�[E���Wf�,�XI	��4�!]:�=|�/r����ǹLT�y;�����
Gt��M��ﾪ����n�s/����>TP۪*���:���G�	��SD!�t�w�a���Jf�1\���}4MQdnU�l��k���G���0�d̩�ڳ�%7`�{VϹ���js��j!��ح���a��u�;Tu��v��-��ԟ�d+u��q��ǜ��'<W$W�L��;hQ�ul��WQÛb��<w��gJ�R\���G.y�K^�f-ʒ.���]l��䩗Os���ǽ�P�t�;ܽoo6�թWo9��p��I�h4��S�Δ��N��ɼ��v _	��햪����{��݀\r5��5�̡�dk��B�}�u7ö��׮��� w�2���,O��f��6T"�w�H��հJ���;��+�6VF�/�5���U�������W];N{Km{��f%>]���h�(mV8§1�ϺVߗ����Wg���(r����Mf<���|M�h�҅=�ӑ�3OaƩ���Wa�Oi�4�1�׋_g��N^���u+wV��(�[xµ�:T������.\z�1�Ӷjf*��T�dGh_�n�>�Ԯm���ݝ����f���Y��4��w׽�.���I�U�vK]֠��'c�ȝ�$�liV.C��P"�>U�����>]L�b®���b#��,�E�Ց���Js�]&E������y|�yE��p5�wX�$�Vk�P7�O�.���+��9�:q�<w\w�ܼˊ��S��8���N��+RyU�pjłH��4QyY�q�[�K�P��4><�!��荝QVP{�>�'D͆��<��E�5V�o%��ͤV�@�ZUs%�i9�k�am�#Ny�F����ǲhJU�-Z8��]+�p��J�v�b�3{l��Q#zGo2���w��7����rs�q�:0�-OGVs��-����Vn�����Ks��S�íp�٠^���u"��y�����Ǻ"��(��=MgĹ��ξ	)��Gl>��33�j�5;��r[��P�(��%u �j�5��,eJ� &wU����"Ջg,4�u�[�]ף����G �]aU�ݏ��؊��7�&B����n�:w`c�7��Y�ЙAl,B�v���e�?o�=�]i�˶/����#�	t(ы����Z�F���D�Cnt}�~hԮ�b�W�[Y"�d}�
�i9�+WgH���P��R\�'�.�3�7`p<�hU��T�+�|v�R�B�,7��J��gV=��>�zl��E����S{�NVq�z�WP����w��D���7����9t��İgX�؃2�T9U�ԖwOJ�X�ۊ���Մ)�C���S}�:���/$�⍢z���'���]��W6���9��M�Cm��3$ +��Kj�����2���C�B����B^o������FZ� ���Sy�N;��Ԯж�
�E�'��I�Ν,��&�	QM���#>_G��ݼ�{�b�#i�=�!\��w|��t,iU�:&��㯖RKo3s)vK�&o=�y�=�h�SĔt���&�bw\
��-+6���3�IfУ���L�#��əi]
�����=��̗{ڙU�їY��-��]ί�j������Nܩ���.�zWv��ռ�T��y���n��o���UcX;��L��L7�7ǔ1��g��}q�I�H�[�ٹ[F q<gX��,ICy�E��΂Q!�
F�3B��u�-P��ڷ�Θ�=rM�O�����+S'a���M<*�au�i��߳@�Z-̙��v!�n�v�.�u-5�r�b-�Q�7��dt�@��y[����P-��tz��ev�PY�G��u+;`l��u���	]�K�Y�+����7��;Pǚ��w��n0km'p��햦U�8V+6���}�.b��������B����0�R&$bJ\� j*�r�����(��

�B�0��(�*""��*��� �
l�R�(2r����",�����,�
�h�*��**h��ʜ!��,ŧ0��
2h�
�i� ��Ȳ¢@���("�����2�+3*��p��"����2+"��L*� ���qh(h�������0���Ƞ���\���)�
B�"	c �j�@�� �ʢ��rk%��*���JJZi&b����̘�� �j

�,j
 �2�(�H�h���%��)(*��b�����j����l�Ă��H������)������Z���"
g1p�*����j�j��r��2�
31�i�H�2���������$�,Zh ����)J���i��J�,�h)j�())*��b��j��
Z�ÿ;�z׾��j0�3��v��s�B�K���o	�K;���1�'��ǌ@�p��o4�y��#sj��Fb�:�l���W�W�T�/	&�ݽ�����s�yJʽ�ܬ��)�۹ѿ;ٶ/hp���F�]n�I�ܕ�t���N����Y{�Qqf|�c#�W�����P{*"��[��uw>��|�=~�G�#</�N��.��3��q:�U�?Y�ۭ�B���ٮN�/?/������� ��t�+��
��]���)�vIcwt�G�#gM��r�t<#_�������N���J�`�}%v5��w#�.�M�T��c�5ט��b:�P�w����Ѹw��&�ם����c��l��7�ϩM��R���X�.&3��G:)�]&��������<�gϽ�ѯ�{�,�$�`K~ݹ�/�o�0�)�����SDy�5�s���7*���{�E�dOgw�`�{_��^Ծ���J���8�.��]��}9Ań�u��E�qQ��U��1�j/^L��se���d�,L&3�nn�ڻ��"�_Ws���[9zR̡͌n@:���W�3qP�D�����E�� �ʅ�O�v� ���;і^Z�mF�4�L���J���_ w��_}UT_�ys�F�r]���}�.�s6�Tv��<�g��^�r�<U@��������s�������K�b��I]��M����� ôn/
+�p"C�����>�~~R���zw<�w�rR'K�)��Y歮��+u��K�U�C��%�;/k=X��E�ݻ��Nnm{z
C�p�L����SytU�����Ͻ�<�y�3=��e��u:ϟz*�\�=�i�3sE!\�ï&?s㑩�E�Z~Z���^�얹<\�6Akn�sDW��eK�79c��plr�.t{�{�{�o>��ċ�Rr��{g��9�ɶ|{粨��5ǹ��o��Eu�-�>���JȮ����ث�Z�Ǔ,�T��'R���*z�.t�&t��e�4P۠����Ư6p�r��ow������p=��nt�g7��ڪ�}޳�1M��Ziw�`�/��o��YٳW9ZJ��ִae�B��2���Y�D	U�G��6�fU�s����WI9umq�8���;HP��W�¼�r����WA5Ȑᴒ4wH�Y��'V)�r�B��v�4����g7x.Ww����*��MK�):��������ܻ������<6���D�Ur�l*{�o�p���ز��NF�Y���*�Z^�ۃ۽�1�����*�k��;���S���[��Ҽ\r�i�-﷜��~ƒ��W$iL�;�}ϼk���]�6f�{���Oyh��;��uO��W�ǝ�"�ɜ��wM
:�G�*4��߻�e��s��v����yןK^����*H��)�S)�@�8v�7�w5�v�y��o^�z{�9@�4��5w>��&G�T6�$��������:l�����[�E�ب�-}Wߓ�k��ݕJt�E�~h�ze�E�^�n�x��%x�x2/�je����Y����S;�������73�s��Dp���REi=��Uy}�W��U��NeK��wQ�j�t��ЗP��sj*��d�o:Yͅ_9�Ft���ث�3X^�U�T}�����o��W>N��Y�r�0YDٗ�<�)��[b�/���4[��*/-�����'-ڟ,V�!4�*�U�JJ��:܊J�a��sw8����t��iWf<�wO�\8WL�^۫�x��*�yϙ�];��8�py��2��()��';2��������ͦ��������Թ�YU{��y�q�=�v=�^����lU;��=�m�W�y����7��|�dz0zz�N�:=���b!��Tu���I���9���3������GK��p'�*.)�q��9�ߨ�/�E��G��q�P��_�����*�z$Q��>�l��T�݅7c9wً�W1�Uj�^/��֮_*<�u"���r��v��xe=�
R�KU�{1�,o��ۡ���z�}��y�g��ǫ��s�_{��o1�4׵��9�x�J��v(�V9�g�%޵{7{��]wkζ9��~N˦|��w9I��Ŷ�Sv(�n�"utt�/�����!�
׫�o϶z)�
�����O5=�v�V�����x�1�>-�=�;�R��חj����j]��KQ�Cod��5�8摶
sZa�<;Y�Af�K�����§���W���F\ʋO�\�X�خ�7���(��g�aY�/�&����q�,���(��+"o�2e>/��T+��7S'Ȱ�@��MNע,-��Z}I����]��������NO�b�_�꧕-�����ej���M*ݕU;�;wZ
��V�}�#�nߓ�S|;+�R��{ �Y^��K�ܜ�9:�Vc~�g��u����=W���u�9OB�^vfW`ƫk�[�WPA�T�J&��\��'�x�f����|�S�}�P��1���[~^����!^��z��] �=��6ƫ�ٞQ���>RSr��uK����A�����+����s_����5:���Y_^�Eō�)ҕeI�y�Κ����������g����T}����B:UY����!�ث���U=�$㫝���\����(N�X�6��iѭA��ޞ��@��/�29���s���%Tў��ap���!^�pKv�eȓ�~;��vmzmt�j)se�:ݎڛnCP��wn.6�er����+yr�j�r���T�i�V�j+��'Y/#Ky`B�(� -vx�A�	+�N�ԋ-m��O5�`��ݱ,lRK�.k;�WN���-�s{K��}V��D�5�c�B[i;<L�u���6���Ŝ���t�U}��}^�ͽ�r�s_�?��F7���p�S7�����UD5ys�d�w��u��z���x*R���zE񮖺���ϟ{ϣS��b��y׾�wl���]�Oޥ��/V��"�o>�Q�������ʅ�c�����d�������}���[���R%������=,�Mxv}?0b�mʢFL����'���@1{���vؒy����ʖ��X�e�����D����9;w.<��=܃�����u<$��!N�*Apu ��HA��,��?v����qkeӿw<��:D/�Zpz���Wr�}��Q%Ul�(ȓ��t�0
bPX�O+����̒-����6vm�X,hC<L*��3������r�����T���&߼V`��5m��ٮ�_Z}���J�Fϧ*�4<i��c�s�!c~�匁��r|n0ߝ���W);�3�
�k9����ߢ�^{n�BFx�qV��2�p�]^����{�\��.��n����6b��-�+��-�4��J7�~�k��i-��L�*�=�{;d�6�]3BO9Z� klY������TJTP"=-c�S23���Sj�J��������\%%-���Q��8gf��8�K��_�����'�6[�X���~��P��sxF�K�ʌ�δl�:l^&x�e2�Tjm��-�V��cwhJ�M�oS�ژ|=���j
�U(��*��]\N#7�$����Ύ%6�߼0�u��]:
��ag)��*����a��F4��ڽ^��o�~'},�9sk�^�if6�GҮ����g� ~P �� 3I���jc1s/c
����B�㭷�V��wuQ��FO�@3d��@i����H<��$N˩������J��l��jP�;`��Y��ژ�s6%��CiY<*�x����m˞0���y�so���??>�����1��8�`N]4UL�"�$EN�T��A=�����}���yޔ$��7�[�lνU����h�T�~��$X���<���y�,�du@:�|��2N.���ׯz��y����>��%�N�B��s�i�"�X�~O���3�,�=�;�k�\IN�oS�z��>Kr,VU3�����2UUT��O�
U�$��ӗSIyei��^B���Z�tl��{���k*=\�,|����իv�XtZ��o#y0۳}��_;�3'u�>\�!�úr-��yQm�1C�z�#An�JN]�A��T��2��be�����N�#F�a&V��ƥ�݇oM���r�-�͍�-u#��������b�;ë��L�?}v�+��G��墑< �n�CŎ݈���U&c����S���;zt�7�=��ȹ��WC�MB���7_�V�6|&јL#ـw���W����]znx��(,�B�P�Wc�=�*-� ��J2���|@���z}�͚�[J��/:��[�4�����@���.I��vk�t��s;S���ZԠB���z_�n檃=�塓�Vݱ�h}nd'T{�\�y�z3k�l�1��u�{S��.8�(.��>[|�����3���7�j4�}�^�H�>�vU����X�)A��R��U��^�Qp�9������d=1ʻ�0.A{|cSՊ����k�%a�`.��
������� =�&U�����i~���K=�Z���sY�(��}��u��g�Ь�]#l��z%�C�.;��L������7N&UгsJ���w�)����KY�jT��ő���d�P�J"�Q�d��v����%��K��l��5<�E��}��3L�dr��ŋ� �S�+��[I"���@j��y�+�pO.������Z��� ��;��2��]�4e��1W{{���������=���H
�.�h�;�Wb�,GV�gl�{Gu�<z���4�9�k�� �Yqi�h<��U�isx&������CJ.�}[?�U}U��[Ws�f1��	��9�=S0��_voe!l��N_'���.�لnJ�;�d>+���n��8q��7p��89-�v�h{�^YˊP�r�;7�Pi<�|Yݯ;ٱ����*�x�w�C�t`��ੳO�q�JfZ��´��\�V<�t�'ekιG1��WطL�O	~$�Mq'���R��:w��+�E���g�=�ә7���^����>�*;���*�'��W�-�-r��ST�^[�:'ב������_v�:�%kW��/��m2Hi�j�!\� Uβ���{M�^��U��ۡLrjӑ�MOV��N��J}�2��R�L��'*ޓ�� �F��B���*;��۹�l&w�>w���֝{����w�kl��<4��7�2d8��Ớ�[q�_o�K-��6�/{��q�"{�W��7��𔓻�4[�Y���e����ؚ�Γ9�a����������t�}v��zt��~�+Ur�
���3JdeR��!�ɉ�\HVw"G!�O�ۣ�/E���U��罜6$Q���)��>j����i�����g�X�d��X0I�9��2��WL��U�3�כ�R�F��*S���Y<ml=�He����VU���g5l�Q��)vmL���:A���1�;=�x�K9Z픋���1���������HQ����ͮ��%���QӣI�v�褨�^6��{��t3�C���7W�z) �v팗ۘ'��~4㹻n�m�*ȃ͋P�F��\UӡS�v^sT\�v�7��n��'*ڜ`��*h�ϻ��������F�wvVz��������
�[���N���Ȉ)O[��񬧡W�zB0>ah�%�Pq����s}�����"U���]���W+��,Rfa�L0L}r�dk7t������]y��Ɩ�y]�u�)P<$&�q�&U4���|�����00���˵���}�>�$}�|����@�t�44q0�_[>��"��d̚��R����Y��-�S�9��yw�$�དL9T
wN�P�`�9g��1ݷ	�;g=�l-_�e�v{u��Y����Tߪ^d�ڇ���qU1A�,6� Q�vxUe鉹r����^ܻ���1v���73�âr�n�<�Iy?B�� 0mq�U1!4,�J��['�]u���</��2��E�V#����lQ�q�D� �̺Kl啵���p�dUj���.����ci��c��Y��}��N$hS�گ�=��jΫ�<7̆aŃ1�(Y=�K�H:�ˑ^��f���N��7G�D�Gn+��|�S�:]�Ȁ��flKs�l��伸�l��y-��.���6�y9�Ϧ����5,�|o�h�%ݛ��h��wL�h`��"����W@Ӆ�9q��60��S�476�v0*DTW�q��P�Ͷ.�i�LY�\���y��XM���^W[�$��7H�W׶��O71g+��!;*I�)�V�S��jU���<���EֹS����8-��=J���̻u��v����+�������N6��u���b���
Z"0��ۗع�;���W5Ѱ'3x;�ymK_vR��X���1��TV�ܻ��ZȲ0��ӎ�*��S��N����C(��r��)2�.���{G�j�P���1��Ks�#���xK�L��S�(��Ywη�#�J)b�t���ms�9�js�]S&�wx��D:r0o��y��dEj@��\��or�3ٚ�˞�4�̺|;u��/y��+t������ݞ1QȺSu�fv�1���v�i�T	�ݶus��*ZI�Ʒ`X��9�+f�!�pmf!2g��������)�^y4P캙;���/E0�գF�%�;�I ��a�8AI<=(��4u�77o8FVNO|߫خ9��ޢ�L��Foz'\���m�K��Sw�E����n��K��5w�������N��.�s��'#�k��Q��]���K�L�B��a��w;m}��i�tb���]/��9*��f'p;xM���o�*,�P��T��W�b��R򠩻Rf��S�U�r�,vcF������e�_�S{�� v�cӟk��w:��껤&�s��u}
�d%S=Z��u-��+�ޭ�Z����3�w��Z��r�2T�;4;-ѭ!v��v������֣��X�}=���pٜ�%_4�n�W'u��eB���ܯ��R�U���>�-��َ��XY�Br4�ΘE����Skj7@��*ܱ>�Wee���e�xc�Fh��@)�PJ�D^p��
�6�6��77�a;H��֫������\��1g�v �kC��}9�oZ��N��ػ�v\*�s]h�{�R�fEG���R�]������`�V�(e�an�R���knL7�n�����SEZ�2��,R\�q����[@�)��hu�'R����9C�ʥC1��P�Di{��a��=|+�^�n:�-9�j��j�΢�Z����{Ow�<2�,т�/����rVZZ4� 7��
=}O�^=�!pu��l�=��B�˺;��\Id�Ha����v���w��h�_j&(h(��e?C�E$K�EI��P�YC@ST��e�NfaaP4�9�5HS��4�Y9RR�e�a�ER��P$UE30��R41eFTRD%.AM+ACAEHR����U�$�JTH�a�M��%9fSCY dU4�P!A�A1�KHP1 SICMM-�%RcXE!T�-fd�PQYd儶b�	AT�P6YNC��PUf��Qf	��іKLM1 S��4VK�Ԕ�EMT��1#T�ESE%!QM5K@D�d�4�14UQYd��C�SPU3,T44�EY���EAT�TKKBSERR�QCM�DATTBRSLEYaT��MR�O�}e��|�ߛvU���AVsX$j�-֚�H���0��!C��r�������C�����)��I�LU�h��]���߱�mC�_}�?�(sW��
�sN	﫹t>�72�+�t6������4f*V�6(M��u���欢��+E��ؘU^��x1��`}�q9�R�6���c��|�4;�){�o+e�:�pδl�W*�4<i����r���7V2=���7�ȫ].����s�n�����2 ++yg0UWz�;���vg���^u����1��Gf�G ��&�9�E�t�y�|=V�ϋ��8���^�TeUgZyM���b�q3�_��9�� �(���龱�u�
���ПW�0��q��mL> ~/Ѩ+}J(<2��U�-ez�1����/�ڎ��%)��l ��W�#Ǎ���t>]�
���ePp�{�PW PN�a-�GX��2��l�UGJK�)]�w,�?( T�Ȑ�f��Q�s�]I\�gg�x���W@�g�8�*����'�������yJ$[R,G�N|#F��93�fK��?Vw^�:��x2Q����8[�5����'�t9��R�΢�xJ���9wz8���d�v�7�RNk�cm�w��3J�/fy��]QϠ�%����V��S�(�h���q[SG�67�S�L����p�����wb���5RK�ʇ�so1��͢�h,��ngT�w�1[M�XԲ��I]i!�񰶅lƁ���YRܜ���U}�H��燮�j�)���)�]�����t�S,���F�X�PUS��;��f��r�����=��:bUg4�����ڭ�����)eL�<���� W�-��-�Y��~-R���edeSʣ�xL�ek�E��:Q�"�^}/Ҷ�`R��"�8�S�g4�ǝ��L�x� ��J��z����|x1�L�O�
U�$�����g���:e��v�l�3ׄ�IA�k���'Ay Eb7o*���>���=V�!"[ݑ���-T'm�[A}�O��d1�Fa0����1z��!��!��Y���b�v�{�|�7��Vv��6@p��K����#�u����S����y���<�q�z�D7���Nh�H�+�]!���b�t"C�L�?�Z��l[�֕ᒧ��ǫ^qy{z_[��ҫ�q��J���a�媽`�󉓟M�c�j�����D2o	]w��s���(��q̻cIUX�XҔ2��
��z�Ö�m${ǆV���3[ʋ��[�킺�|��B�����
�m�u��ݖv"�����`�M鸸+9���+�>5�g^�����:*�M�E^q�D�Oz�*b�j�YQ�C9�s(��>W��[����#s�ɮ��HI���֯,��L���]��eq��&{W���^�������^R�*��q0�)��d"S�P ��;�S8�Rξ��ޒm<��E6tJX�{*�>.�`���6ϢX=P��`]�D�
Bx!�*:�^���qi�����t[���14�:hxc�'�5�w��wN̤(񫻹��=S{D��N�������<6����:Q��Z#]y�43G�8+�Ύ��#�n�z|�7^��
l���sφ�b{�;�y���|����X�SȎ
!`QW��of�s}��Ls���f�
�e?�����sNr[ǫ �>���\R����IK_�<�>˷UO��0�K�q��?�׃��j���o�,Z)�~+i�f^z�M=���сۯۆ�b>FT�]4�̐�,�Ӥ��u�
���a��U�v���❯9�>M<iJf��r�2��x�5�.�E�%�m�c�C|n0>`��I:���޹���K��-2�AoH�z�݊c��јz��CrMYC]�KV�����qmkH&��ř�ʹlã+��#|��]HJ�5&�w��'�i;������='�
zF�Wm5�:���o��Z~��ȵ@gw|;�jN�{шjTlo7�w��I n���ydY{�z�b��jK7xd:���%���A�A��'����������.��a�fr���Y��2��P����ʾd�� ��V��S�/G1������Ux��fe�^�3�p����>�r��}�2��s���̨��.�^n�N;���o��AP*���Tgȱ�{ۙ��HJ�
�nR�e=���r�g!3ʇϝ��S��Mnic��d��Ua�kΏ�m?���y�t&�e/-�ʥ��#Ǔ�����9�˷A͞r���/��9��G��*�ΊC�x���V�Z���h�u��[��Ga15vn57VL\2R���|H�՞U�r�P�^����ɖ]z�J���c�|!���_[S�ˬ�}����#��� �q#g̞�mҏ����q.���w�'õd�jS���_ܖ�,}�HM�db��aU׽Q��[�/4]K�%�UGjCa$'�J��M��ȸf��}1��C[�6�ב\��h=�K��_��J�.����$J���4�ݍ&��k'����+�����`I�|��Q��6Te������K�a�^�Y�.R9�����H&�>�RTr��a-�@�	�{���}˨wu�ZP�z/C�rP�� ��q�(�Zq�z�bS���Ѷ�I��JSq�2�|D�=�eFn8f�*cVs�|D	�ʖ;/�����w�_���i\��GkCF�m��L�N�i8���"��&Lʚ��[���Ǯn!��?�N���R�nh�d88{$�ད!F�vQ��G(O�.OS6��T�^:�-:���:�2�Ʃ����v�þ*B�Hr����*�X�)n͉x�4�;W�p5=�<��>-JJ�*�9H}S�3�S�Q
K�i�v�H.�ى<>a��4
l�\y�y�/r�����e[�a����הIl�=_6��WӬB�f�ĎV��r����˽	��H|E͉�^��x=��Q��X�w�Ѯ�W��m�����i=��z�g'�L�mJ�Z6c"���*���s�<ɛ�bR�$B�)>3�`�=[�@Ϫ;�gyb��)�����<H�q_��ʭ9]AH�J��WG.E�S]���'|:�婈60myǄez]e���X��^�0O�c��x6-��:q��O+�ް�~�]%³�F�1jbe�0�z����wy���`��@~g�0fXZ�L��,ˢ���95@��S��U�hӬT�z�=��m:{G�V:u`�p�����s���wo�N`�r5����m�G}�iYY��u��{�/뼳W��:1�J�w�l���������}q(�����yf�?���;�͎_�y�',��`��V�t��s�k�
�qA�q?����DVUң���zop/ݠв�	�f�z9Ww�\�9 ����9Ol�j,(��m�����郿w���(=5��aUD�<��tEh��a�!#']O��Y'�o��h:{������]Q��0OhXy�X�aQ:OPD�3.�<.���p���1��޳6�p�>��y���V93�z��G�KF�$E[C�/��d����7�^��c����G=][]|��|1�ܼ6���+��2�<�̞@@�o�y���3���cl<K�� %
���q�e��.�����}�H�i��`x�,F	*D�{9���[��T�>�c��c{�M6O�ITe�>��sA���L�OХZ,���yzzv&���>8&w�g���h����a0�߮������Z��һ��.L��5��wq�%�3��[AS�<]WF�"8emBוK���'�Uk��vl��G;s+����y�&�{�;n�.j[�{fg[D�=�*�F�9#خla���ەFd��}{g9�f��y�ʕ34�O�ZLA��v�&^��*����Ǜej7��nl�F�"\Y����z�gm�Ǣ��x��@�c6]I��1����sޞ�T���zr ��0��d o���򧖪c�#�0���{"�����b��m�f���,�Ƈ�Ͻ�l�"�g((�ΝdTE�����꼼������r�J�J�^纮J��w�ϒu,�#>��c��v^���C��8�3r��꫃�2�:�9[�sL��\1vz���.��p�4�R�S��R��U8r�̯x�X���! G*�|�en��P�X�VJ0T
���&�`.sS�^�窠=�$4ֹ��>ܵ[�=�wB�y���'��Ӈ�Rƫ�x�(V��$z��Uވ��t/�[���N��l7 ds��g�k�vT��ܛllb��}2�EY�H�]0��x�[$������w�g���׆4���lM�N�"�U��m�����"GmD���Ca������6dt���W +��\�C�1�p�=9\�{)��w��9lt�#��g.��\a�gs�D燛��L�x׀�%"ڕ����sNKx�`�>���e&��`�o�-�Wg�m-�\]:�l70W3�fRy����ݢL37���h_kr���{��&��h�����5��g���]�K�:� �RTL.����]a�f)�b��;shV]��&s/0����{�"/O���eoq��V0��[�y��=n�}ԯz�K2�#A}���t�q���m�t�橂{ҷ�^Y[=��^+ײ>9i�+L��vB�������4���O5������d@_����c9�^jܵ�[h;��g�X��S)1ު�V6��
��F�j��/��.�Ew ҧ����S�ݙ��o�;MxO��y{�	�.KL���z�݊avt�m\��0��&Y���A���=>J2=s6�nج��J��UL��*r��9� �������՝�v?Tj0M/+_n_i�,fKP�׸kEZN}�R���Ax��>g|��Pcٲ�y��/-�@�a\/���w�x{>���*��e�<3n�E�}�x�fN��,{�O����W�<W��e�]�����|�_�`��i�d���.��ܫ�˥*�R���k'5�g�/x�&�d��
cEYK���'�Q�n����k��i�/G�O���8�12���Ў��;ѵ�����g�exp*sƅ���ߣ�Z��U�D�w�=��Nb]��us����Y�_����<n'�c�ra�x8evVrs$Gd���]N3-EO�S�p+��X��܎o�4���gP�#,T� Y�L�a�j��s��M[W�jz�ި�������3j��A����6�WVN޽\�=��5�+�W1�D���8ʥ��V����qW�M�ϻ˃ϯ6����>,E��=�[�>���cP��������U֪;���fMD@�m�c��Gm3����	�քg8��_eׄ�0\�a
��!$���v+U^��xR�x��0���$���F?l�lx߶���pT�/�Z��E��d:U@�p�G��ӛR����{�W���6�ci^M��_1ۚƇ��	�|"2������Hк�<L
�[>��"��d�r]�{;�v�]�=�r���a{�3G	
�hR�$�]u�B���9Vg���۶�`3������]�OV5	�lq�����K̮�nC¤7�uLPnO *� �%�R�/V�e��ߟZ���i�$f�Q*�*�ܤ>�u�s*s�!Iy?B�� �]���VKǦ��}�4{"�$1��[�4�}�}�(�!��ɘ��%^{�YO��X֨wӻ��V0�)�1�ۙ��N�:�`V�c��I{P�F��d� ,H9�ܯ}�r⨉���ˍ8m��A��O���qc��~�כ\��Ip�˺���Eޜvܗ��c�֋<ew<JƄ�e䝪둭��]NŅ�-�IثY1:���V�x����9YjL�-�e�u='t�s��F�w�D%;�����|��ܚ��5���vNV��=hh��r�:N �|6ԯG��pc�}0Y4�h�y�=��#��?�߽&�ur��"=G�	���s� )�޷���Y�V޺��do��fE�A��6_�O���{�������|���������s���|r;���6�M����2m���6/��$���g�2��\+p]��Z�ʥ��]�po����PV��`��E=���H�]���VZ�ǫ0&:%��K�
��U��Ao��)��*�Pq���g�n��uvj�q�闻�&��J��V���0ͻЙʫ��2�@]v\ w�����5����`�]���G9و�Hup���<{��+�n��0*;p2�(�u�ސ�K��گ��t�1xf�4�d�������*�]j�b�,�'�
�f���B�j�D��-[��~��,���54��낲m���yk8=X���t�z"ܑ��
�����/f�Vo�'v�y�Q�����˳̪����yZ)Sq��r\��c3������3eR���LM�:�S%�T��R�;M�&@e��Q��
��iS㓨.mg	MH��V��b�O~�wzb/,Β���ls+zs���u��'�.^�w��"t�< |SW���+8�m�w��B��&�[��=�-J*2��O����*q{ٖ����+}�h�s�c��qb�8'M �+&^�B�H�	c��˘:�е)��~+e��s��Ô�<e[��5L%&�|��v+�В�6Vo]olb���C���WgQ� ��z����n�F�̻�b��!^h�	��O�?[��h�ST�)��9���5+iLZ�9w��u�z��g���%�֗Ǫ�I�Tj�]ܺQ'»Z&؇��yw4l4�,��anv0�6�7[�V�_q���+llU��ov�(���Xf��.존�p���Ύ��v�����Y��b]R�G�� +���q����V���i��vU�Y��	'SO3�%�VV��<��X�$:�Gϯ�\��X7�FJ��;k��4WU�6܊e��E#�v=ᬨ9�.�]Ei���Њ�Z\�t��r���4�F�5�Kr�Lۢ9VY���l���>��R��,�l�V�we7$�A�j|�)��
艷���t>$_f�ͣę�6v�9\��z�iZ�.fn>��(�;�,η[��`
�K��D�+���|��(nhN����j厙6K���*T*i���Jws������y���Y����ڹ�����͒��$�5`o�:ծ�T�t��g,���s��7R�X���DJ�4��x�mwul����Gv��Q��-:{�<_ct���]B�e�˨�fm7�Q�Vn��n������^^]�Z���Z��gz�>�G���;���].v�ʘ�;˖6��>�y�=�f̑+3G��Ъ8q�̵k:Ch�v�a^��U��X�%�l6J�ƛ�v�I]#۹J��O>�u��}q=�-GN���u3�Jn���:�W��F��!��f,�usuom��ス�Y�q�:��将�;#�dZ�����<����2��jJ�}�=t��]'V�n�s#�����O����.>r��N;�y���
�]�+5�&f-���6^����x��0����y@�I�5��.W��.�fr����h�]�S���;�f�s��ތP{MP�R�.i+�A�[��\-��=������D_gq�دiD;j�U�a\Inu��r�iՎ�ҷ�8�>.�λ8��[!ʖ�`��G]�z��!�w^�nf9�:rv�(���X���[$}�$��.Y�Y�f%xJα�紺��avXFW5\�f��ݵ3�>�3���\�9��7Id�����b�hO0`�=�rtVi[��w:�^YWJ�:��FSj���6�`w3�{��毶	�6Й��|�,�j+9���:k-v::������]y�4PNXDTU4QE!HQDde��QLA505Q-P�DQ5M5@EIAM4RUUCCEU%�+YIE��ED@U@LU!T�Q�HDĔ1C@R��B�S2�@PSBdP���9�%5BP�HUHdfcY.IKY&QA�a%Q�4�MK99U%4�Y��L�	IH�5LSIA1D�Kf�T�4��I0���U4�f!�ILD�%4E,HPU%TQCIHU4�ESR�T�@RPPPD̔�E4QMY8@SM!T����TKFXQ3DE45A΀*-^KXY���3�m�.��(E*9{ٌ��Ѱ������ۮ�q�畵��oB�u����䓄��K�jsդ P�;��]N+6O(��*9����i�ZrK�]⻮��&������{kjf+��!o��]%��h�/�xu�kd���W��c�]��;B��L�n��Ć�z����w�fY�<I,��j'Ax%Dz�B�؅�t2�Y�;�%>���L�m'C>�ȭ��}O���G[Gе�R��y�av�w��&�=��^�wDAU�`;��	�`��v�W��,(�l�c���]�W�3+���7��f���o���>]t���Z�U^q�&��E�ח�A�)M��Ď�3$�j�<9�
c|��-��CJ��2��-����-U�s�`�U�'k�g	/�1�Z�jC�p�9��tU�e�'Y[w�����)C)��Gn�=UnfW�#�A���߲\�Q��lO8��;�UhB����X$%����U�FS�P hr�ӧ�^o�m����>��*y���CN���Q�B�R�Ѷ|N3���OSR��k�I�~������:��C��up�n�1a�f7��gZ��ڱLG׉M�߱w�S۞Z.߅^e[2��5�d����2g(���ٿWV"�O����r���u��Hή
�������̂Xж]������<\�����&�J]�؛���LT�llb��}2�TU�4��]1�����޹������Ǔ�6}I1�}��K�`�ꝄESʴR髸�is,�Q"8V�v����~��{��Pp�L\�vU��2��b{�;����R�쾧-�����c+)gK��ܕſY%b�:�!P5�5���\�L�}�o��>��49��#d��&��#/5X�Q��}�zׇ2hO���-&#9���ז�]�u�nz%�ۏ�V��O�{ݫ��y�+�(=+NWK�j�F#�OU�_<Ds$2K04�J�]t�b�m�IV�kq�Y�񕥆�TX�~�&;����p�[�ʺ�Y&��b�/�'S�6s:���su�k��2��z��/7l	>�� d�� �d��*h\^�+���s��x�r��F3��/��s��7lVwED�y�&`t�oIΈy6o����'_M	�ܻC��x��t�k��ˋ�����}O�p�S�I��)Q^s �k_�^YӳLE&�c1G������X�t��+UY佯��2�k줨e�Cc�>������tZ,��Rt��z�%��LHN�xu��?
�'���H��.8��ƅ�v�ީ����|�	Y���{���e���]�˰6��V$����|����miC&|m�C�^�c�Ԡ����N�
#F繨�:wdBQ�[�ܱ��0�n�3O���iо��+N�M��՜UdL!�S"r5�
�+�F��&��x���R$+1�5���*i�OY�UH�s�l�Y�
E{)pՊSW%�SO���{�h,uɔ�12�����ӎ����}~Dx*tn<%<�1;\¹=���^��S�.����F�Pgh�ʫ��UmN0{����x7;<�n�)S��̃�;=���{]�H�e݆A��\��_�	T��3&� A͸2���Yo�dyY����wLO^Rf]��}�I׾:�4)ԇ~II���7F�d\3Nчo:�{�Gk����ٻ�^$eCQ�ʐ*b�B�SH�����J����X�Mr4RA\������-�v^{{:�2�
{�xg�"c,��EU2;�i��&G��h�=���W��5�s}���=z���Kն�^Նd7N�\�n��6B�V�(ޅ�w ��Y�]˙r�'�Ė��e���p�雉�+\�ZZM�r�L+
��k��+���c`��s)���҅+�zY`��nQ����Yq	#��m�,<�w��z��\�e��+	��J�!B�<�G�7#��t�q�u�9k瞔�!�'(�ūX{��p5<�0d�i>j��*�nC��B����ܩ�g�9'�e�n���|�S���Y�ŉS��r��u�rsTGIy8.ؐ6�h-3��zd�^�y�>�Hxt�c*��~jS����0u����ٔIR\t��*L��<䋤/�r�>�Xg��D�S���� R~�bc=�`|xr0Vm]��wh�8ԩ�[U-��/��Z:,��qS>mJ�Z6e�3H�#�U�Զ�c�Bs�қ�ztO���G�<<"�s T�����Gz-f�?	��8Z7��0�׎KI5�����p��ݾ���Lm�7��PJ���0�P����������s��b0Z���'���3$zߏ��%��Ү�%WʼV*���]C+�k3>Z��V����f�+Ѩ+Cw�k}G�C���߻�`���*�-	�w��`ԠA}�Hp�n"�7���=�y��V�{s�p9eO1q�5�ī�E���|L=�m{���uUX�*���5�Dv6���U����鹾5t�WZ��N�1�f����
��(��g����ĩ�kB�-#�|=�|e۟wT�Y�^,��H�uc�$fQ=)j�hQQ�]������*]�H;5�!�{-FOg)�����m��ǝ�ܙln�g�}F%��8*�����T0�l��������͎�O�CP�$1��u=�Ɖ]u��"ON�0A�Pz��]j�b� �z�|N� K/GDy�$�s��y�����v��Ϫ�ꂽ�*��Z�c�<4��L�(I{�����̼�n+�x�xT�2�A��^��"�|Pʭ�����E^�Lf	E�kwg�V�qwm9\���@�* ?
��|j�Y��x|�	U����M?}�����A
w{
���ƛ|ݗߝmKV��
���.��	B�Z�_����c������خ�ֳw-�C�j���Z}�`8������fY��Z$���j'Ax$��=>�if�/�};w{��wG	�Ȓ��"N�IdV�p�>x�t��G�}����F����cb����Bo���L��s�"
�s )�F@T������쳆�r{����}bo�U��^�ز��:�*���Y��op�}N��-jP#�4G	��6�� 93&�/∴n+gG���{��vWV�s�r���F�G]��sR�W���ݗ��]U�<6�Q�{%�O@�s��bArw���nA���/�3c��/�E���D2�N@��ո��],֮��������-�_^m�+�\��er�/;�C�!�<���h,��I^*������nI\g�����`�U�'s�=��pW�S��#�Wf�b�����pR��FϢY�'�p�\���PWit k�:���-�OM����:���V���2�y�h�
�EZ'�-ނ�ƀ�]W!�����`��.:r�=U�	���qe?3�ꆻ�B|�_�3��V
ZZ6ϢX=y��R��~�ϖv<�ϨJ���HǢ�'*o�Btv&�I��D�Z���ּ���i����%�F+��tK_����P��C����y�����Z�ʪ�y���!��e���y���V�6���AQ:)��Es)D��_<d�����jW}1��U�-x�]�&�o��W�[n�(�	����ev��g�P��C��H�~��pr[Ǵ���T����]��ܭ�w���	#�>�Y�|��U���,U��Oӛn��MW����i�w�^�~C�1��j�
r+g�,�S�x���"�\L��������I�"��z��ZE����%�_Q�IS�Z�ҁ���a�]5���9����tǋO(>�g����5��Z븹���U�fu���xIa�5�-ܪ��w^�^�M���y���*�mN�o��32�}�W\/�X�j5��d�O244�<��i�n�U+�˓�b����w0c�Dw���	�B�fZ�|5˨�P��[2����j��Kʁ�R���U��gO${���("�^�P1�[��DL�x yP�d��[�z*�]�i����E{�7ֺ� ����rϼ^ng�k)�nج��D�<��ʅA|�[�s"p�Z��f����|��[~~ l(X��ן؇�d��/���w<��r�E�<4��9z��]{���e��a�!Z��߽�X�#�!
ղ+�Ԭ�c-uxͻ�4[�ق�BV8ߴ��Y�c�毅JǴ�ݭ2]M������pc��k���m5�ǥ��ՠu���KG;}[�g�D�\�l�|�xL��!^��Q�Y�����K�9=���%C�`��w�f�Kޞ|��Q>y��r���:$')jbe[������jw[�}3�*�� e����|�^\�ߜ��ŋ��զU�#J�]2iЬ�"�2�E��^�"�ڜ`�qW�M���ý2/��Ə�g.^�O}c�Y!�pBv�4C���|a=��lԯ
�ԣl��[�W{���L��UB/YB����PVn����VWK�|3U�`Y�fIuo��LN崬Wn�9���qȒ>�}�; w���ӭ��<}ԓ��v'��RLR�N���eX�=uʘzZt��ָ�S7���_6���MU��Aĕ������><�;��(Z�v���:���⛦�>I�~��ҁhO`���Z=>i
ֵ�>�R��Sۅ^>��ɭO�Y�+;fL>�k�����]ji(����×E��A�뾆��W5ffy�}v�\�J����ߙ��=�<1K�q h���u��BꙄ��Q�Ý�V�k�țr�Ǐ9m�u�د	R��o��<��pp�I��{"xp*��t(U�������{)˯<j��3��N��{��&�Y��כ�^f��3sP��"+��D�~xo���f�M��`X��v`+���%O��w!���s�ԇ�C�C�s8�ǖ��a��ٿ1�6���B��Y��C����ǌ���I3�/��	X^�'7>��b��&gP��v���1(2������_��3�����烚�
�!ŭ|Rq���h>(yza'z����T�*r�Γ�8��Ġ�~��2��L����$ǻ!�<����x��F	[�Oǆ�Yܲ8`��`S� ���m�Ŭ�����.}�E�����]�>*[�6�
㸬�9���x�xњ;+_k+zEW]���xc���<qyԑ:�>̛�2*!^|4DQF
�Ee:�m�Z�ﵷ51�.&Ю_i{�1&�q���j�uq�z���֍9�����U{�l��5��[�m����y����S*�FB��	W��J.<2��<#>�����Ăuph.v,�o�y>�
��a�8-�~�3늴�T�v�C�ka��S/��PU�Ù����{�\d�5ܽ=��nފ^����T��K��w��}p �wHp�����؋W2+-q�sd�������0T�+_���&���Y��XI-�?0�� �=�W���{#����2���UdN���:�5��q���(�&BY��<��KS=~��9�u,E���d[�ɫ���f�R\�up�|n������g��1d�z�Z�'\;ы}��$\{ap"���'�+�S�}(f����Y��kK���e���e��W��f%'�d=�Y�h���h��g�9�k�c>i���/T�Z�'<��)⒅Ţ�זO���e�)��,��S���A�? B�(s8�3����z��>s�޻���l��<�Zc��`�r��L
W��H���x�%�?pj����`���\�쭛�ׅf�ʦ?vtw�M	
�����Q�;@�Yi��o����T�Ն���r�����[�k��q���$8��M�k=c���)�y|_!s�86�Tm�g26�����t�EYYǫIw0'��9Vor1��L�_6G�õ,|�U�b����f�jw����0ų�sҷ�C+D�����3,SĒÈ�a�j��/�+{Q��q�s]��=���h3�+�"M8`}P��eIdV�T������,*�3��|���i�1;gbܭi���^b��u,���>�s *��dT�[ t g�媜���	$z��ݏ�74���������m�f�|�t�V�(���0L/I���X.�笽��'��@����)�����:O�Y�5��WE���ǔ��e�W�w�+ڻ�w�{��3��Pwo�������0�Ҷ�%Ud�^��
Z]ɹW�^�|��=�v/O���J�q�w�~�U������]��g˖�0/\1�fV���{��n��� e����1M>��<���L�*
�9VV-9�Q�}A>��}wӃ��@���l��E�NT�9T6�ڌ^�ɗe^#ơ9���:�Ĳo<Kq�.�O�z�Uf�LJP၆N��pM�����h��[��aU�7���#yV�'jG���vn�(��}-�t���m�}��9]	N:״,._'o�%-�\��$�-:�J<.�D&(�6���U ��ڮ�q��ܔ��;R;�ɸ�켮�����D�D�2]��d1����̭�w�&�LǮ�n�a���[|o�q���I���Qٛ�	k��v��ѹ�[��cX����[��^vv���6-�r�;�o�`EsYX�n�xƛRI��+�;��zN��)��/����.=̹��}��u�p,y��Р��7��.Vܮ3a�����A��v�/hC�EX�0���ۘ��]�}�[c���|nJ'E���������$�7jm�`��:s���	�bjoz]��4���c�5;ٳ˄��vd>�c�IM��	�d��2
ݱ7k7��F�[=��<�R5c6e�g���QVi���V�T#���5��/p��gl��˵-T.YS^��ו(�.��=�ˤ�uǙ1hĉ͹X�V𸅬Ag`P�X�SF��p}��+s���k6��Y�]u�VD�t�G��,��L��i����l��dk���<nX��}a��Go!T�'�@���-��c{�N��(��m:�u	mе�u�j�<c�@9Յ���m ��x2��k-��UF�}i���`zɔ.+��&l���q{y	I���)o���}�Syŗx��.�h�ʚ�T{%6�J���*�:본�|�hL�t�-�b�,
�+&�y�U+�}�[��Ƴba˝�o��з`�f����f�xlUʾ���M��	�δXkgW-�p�>�Γ�ڄwJ�O$H��,f����N�2C����(������Y�N���3!0҂�+"����Ȝ�v�s�E�ɨy�6�P��-SD���[�d&n�e��̋��֥�(�0��p���4�-edʱ�Q<�5uu�6��2�u�j��!��wC����}g0�̚�|O_��Ȏ���υ��^z���3p�<�J������=o*��8CC�r38�����AC����c�8NZF���Wn�66����p��Y��]=0��͉��fͮ������gDwv�L�+i3-��n���ڥ�e�2<,c�Y��S��_
Cs%��J��Tuϛ�v�tn�;��2KO'N��F�V���.	Q`\]�s���>b�i��H�u������[��Q3+�:%&n�<X9Z�b<�ÖukS9�Mt[�,�`����q�v�WgV�^Q�}8�WX�#�w��e�����P;���H��D+�Ƹuu�l�{6���]s����*�W
ԧp��wd���� �5��`���oS�Y���y>���k�;���KG�է;�g%�u�gv���ʗ)�c�
���s"�����h]�{ 2`�Pث�ræ�l�/b�j�s9�w���umn�#{y�*��D�y��^�]��������"�(��*�&
F��
�����i����V���h����	��,���(J�b
H��������	�*)*���J
�
i����(*����%�a��������**��$��*���b�(�$����(�%""	���
)*����������b*�"�������r�� (���*�
����2�3\�*�R��)�(��b�Z�( �(r2k3��bL�	*�(�b�(
��g$2��f�����(����(k �(hi��(#10��fZZ���"*��2Ȣ �)�!_@P|(���]uǏ�	�<���ś*�;l���i�GS;h��`��۶�\T)d �;��)��|Cn���c8U��k���Ƴ�U£��D�̪Q*�猚�X���D��!��7ۚf��混ޚ#�ۘ��oc��8K�f��|h��e����W]�<�ۓ�$�n�������=~hK��,�C�˰��e.�D����|�o�P�t�7�n�Jц�s/&���mcw��&5�TX�`n^q�K�j�F#��t��hs$2K05���2ZV����%��>#�yQ��2�g>��
Lt5,��e�Je]F��J�z���R��������?��������4��9[��DL�^�@{Hf5�a��iK�y������A�T�0e�g|��_f���v�fwL�|Ԇ�UB��e�ͫ��_?s;Ѷ/7��I����B���^d{m��	�[|3䗵x�����S%pJ�3W1�~��6�Fu���b��|%�����]Q�+�|��c3�A6��.����w�J��u�P�/E-r�{>{1��M�����iз5A�[�\>�v���=]��gB���P�u�Nҥ��ѤI�1KWl��m6A�-2���9k��^���}��E_E���9+�1�y�ă���ڮJ���a� k�D[����yH���/��w��a�f8�*L���V湝�8�g[��^kK���
�1��!#�q��	���xN9ڬX��&!�'�C,�N�,d�|��Z̶�Ӥ��
��g����@}���+g�
f��+�-	C�C�����[��ޮ����w7mM�5�X�g3����.�\���i���)�����>A@����*��L3������=E�^�	�U���?wv����2�៪��dhuG�?D��XEC˂�N��76�J=�6�=���zGL��W�K�ٯ}8*���8h�R�htq!�:=�I��H�*�w�1��Z�z�)u��39�eT��}P�3�8*b���M#��*��.��DٻB
�'g6���>�{Yi�'�g�j���	��{"�|���.$h_�x�B�.�v��Fި�;ӌ;X�R���֡3&�+FT�,���|�gd���"xr��M�h�E�s��ǥgk�*}�/�UVu��ulr���0d؋5�G<7�Ew��qRˬ��>f�V��
I��Ru�R	��`�?Y��Y��ͤ��_{����a�ʎe�����+�p�R���}�}�e�E��uwi`[4�E��c��ƞJ��4��r�t�r\,6ӺĘ7��jY���|.�]��w�}v	qO.�hv %�ͤE ��v���t;y���]�ͥ��:H{B�jgk˧�V�̗���h�r��=}f+�ޝ7�ۊ���JA�1�Y�r9e���m����8u�S8D�NV�M��d��V�j�+Ŋ1��C)��c�
�%?Y��`�����1ߏ�9�X7����ѣ���;�$�tu�N�r�Œ���C�s<6�YG�R�L�GZv��a����Or�j���b�5g#�ܲ8`��`U=PNe���Kx�%U�`�ϛ���F�d�n���Y�9�mW�
��Q��7�	^\�&
���U�X�=�����]����9��M���b�M��q��]nW
�����ka���12ژ|ɣj�^��B��5tޅ]���qA[�E��,+�Bc��c>�xa.���J�`U�x�qWl��8�N	ͷ�������$��i��|#0o+�+���l��и�]N��G˾W4Xo������c�;��{f�3�L�bz{c
��PL�Wt4��d9Wփ��=��'u(��W=����v���r�Hv\R0GHL75��u^|e>7W&����b��>Gێ�r�� �
�s�A��[|�;��Β08�nMS}��[��_
��Ҏ���%���h�]��W%�歕�R���+ '!�t�uz�8C8j	r��Ik��!ёE�6��3mɆ��87ʝ��Â�4�3�p��\`�z��� ��}�Vv�v�o)v�A�g{ywf�;(�.rj�r���Y��X�j)��K�zu��<��p{y�.�>��ˉ��Ot9\�����t8T�d�a�\��r,e4���}+{b�t<$}�u�Gy�#L��0���fiS|�̞@A g��.�po�!������^�����M.��磙Y�״�4��6R���J�10)QGBY=WlWYB�۬�s�!e�u~n>l���q�F9UL��J�g�#��xFn`R���IN#]��Q:�5�}�V�-��Fͽ~xD�$^�%�Pu�&�0>���,��
����T���$���q�tːw�ig���~���e�pmq�0�wDAU�`S����ʶ U����m"L`߳�9�Z�v:��m�p��������U��巸g�����@��8��P{����~�׽Y�;,
�,YPnط��I^).�nxөy%p��a���^����t����w��*%zjd�5�$>1>���+,�n�;�|/����v��g4��/�n���ۈb{����&����3���.�]�hĖk�z�,Y�#�Dem��5���I]$���7�1lu�3h2n�����,�V>�]�����L��=���)��8P��S0:N�����\�����c!;5&e��y�.���]C'!��]�Ӏ�o���mT�\J�8x�U��;�~���XUf�]��e.X�Ẍ��n�s����J��=�l@F�_ye6%��4��>�<�n^#
­��9~�cKp�{����V_P��n1�	ʚ���*�LܛlF���O���|��n+;�u�;�4����u�
�-Y�׉Jaa��'��$��Z go�ǶiGmI�����[�lg�l��d@�,_�a0Wa"��UF��sg���~ѯ+�E�I�^,Mm��cJ���r��d�G	`�����h��=f��1�n���VʚJ=�J�_���wrz컊
�zJ�gX\4ho�m.�e��՝�5۾������U�k���l{��,Z07/8�%�5c*e�3(�j���G{�A�����*8��������jU%^��k���q�#9(�I��K��Pɗ*�WP���U�9��rOzu���=D�X�!�z�߽��i��5o��DHP��Ci�2���/x[��YV��#��=ޔ�\;XW����촬4;���y֖)�R��#��x�}��~�~�;�WkW��)��p�7j�=�.�}u
�ߥ�.v5}'�dJ+��:ف&ޓ���,;�3+n��:�q t��a*�kkjB������ƍ��.�^jw�.�Y��	�`��zH���f{Ʋ�)��>�\*J�w҉w��(*�c���ڙ��sp]TZ'���� `a��cֲ|��*��w<��-���=�&�_5�9���&W�R���J ǎ��5V^D!@�]+�C�+�E����x�)D}�n���7O}�����P�ފZ�*�ؙ.�/a�}�:ۚ�Ϸ׶i��<�b����wӴ�o���>x������!r��
�Uy����s������¹ڬ���nȻ,�y�WV|)*<+��K��a����-jbe��=���jw^5�Oʮ"fe��z��I\��$=/ȏ��j6�k��B������g/CU[S�=b���x7�K�w�q���PoOe;�oG�(�����xzRXϧȪ�N�R�Ty�J��a�ų�G!U������*�.������W��'@�3�Y8HI<%�+q#K��8`���Y�'��n���^��39�Y�|n����å�\<(��|>B��`bMes���V1W���l�E�Ǯ�Sy�VWB�,�C�c��P\*��4콮r''wi�M���1�%Z��Hl[����)oB)��3k��/2��$�+���Gj_Xf+I9YW�+�X��c�Xe��w`�ZH:ݶen���o����yԘ�T�C��T�k�9��*��b�x�"+�@�u^�4u\�G���ƒ{q����ћ' 1uK�.&9��6�^���2����KBR���_4r{;�^��w.b��B�;�B|.h.���ЙSb<D|�9���3�i��V0�W%f��bI��#r�^�p� V7g�V\<�����qRN��G�O ������g�y��bF�T)>>pZB=�<�|�¾���yT��^8ps	%�����yW��l�Z�|8��$�X��]B9a����@hS��8f�]`V!����N�~�s�ݬ,y5W5�i����i��N|�����R�N�'�E���M�;���#ˎ�[�tO-����N�&<������8`�q eS� �s��>�{ƴ��'��`����Z�sO��2R���P��V��)�^8l`߼���={�C�ټg�%�[|)j�w��i��>�9`�[{�>�LzU%~2/:��:�K큾����ԭh��n�.�Y��uFV��:�n��1o�s��~]��1���zfힺ��_4��zl@��=�gIB���׋1�݂!�v.r�+3�_t=�+����;o��1��S�,S)̗��5%ؐ���l:W�]�F�U����������f��^i�!�4�ލA[�^S��^��O�,g�/%�R���P;Õ��F�����S���_v�K�X��i��׊��+A@���,�����/x_G~�'��{�豧�{�	^�p �z��S�0���je3��U�pW���HV�N!V����&]��/}�}|�Ӛ֎ �qrBe[R'SMF��G�W�S�ub:M��H5�S����,Y��\��x*Ī&�*'�̳|&R���SO�^�+ޜ���yk8N�ש��������>�{�֑,S� K�/�}i�ս���)YС�=��ȑ�]�N�������-�o`��5���=���<�@-�@B�>Tj�³x�y��=�*�i�2�c��-4���[k4�y���$������\
`�/�Y*�خ������O�Y[��WNb�[1���8�t9�Y2���FT�Q�ϜU8̣̲M���ܰ�;��"o���Q��h�r����� ��d��8`yP��HH�P�,x��%Ns��n�p����`/i�	}���v���v*f�I�������XSN49Y��Eԫ}Ev�R�G{\{U�%*�t%�e��b�L�XW\lf۩�N��s�\+��l�rkR��Z"�	��w�Xp�w��z���Z�w<ܛ��u8�>흭KQ��%0������g�k�Yu,�nx��� �Q�5ʶ ��p֟z��I���Ul�^�"kp�^�z��U���߰�`�=ZԠCS�;p���b��ft�w++dp��v����J�ۯ	X�*�L���^W�4�=���sORq��R��6ےǚ��3�hx/��2W��7/��3�X�H�|KG%]�d��S��|����=�koO5�:��S�*�̯x�Y*�5q�ǫ�x�RH�������h���AA-���NQ�Y��`�4t[#^��^��j��pB:� �����W���)��ٽ�˼�Ai�ߏR�ڂ��N1�	ɪ
T\��������<��m_h,_r7o\���d
�x�.�B�� ��%(p��%�'����c½��z�d�Ż�̾��s!P�&Y���h2�)�+�J%\{��!��|��V(�|;��S׺y��4{d�X7=n+]�|&�p�=`��ل x@(W8�~��C�Ս{M�ג*Iw�-q��ں�i���t�f��X��k�W����Z]��z��i�$mP�����2� �)W�a�x�����Ε���nA��~�FmnN�=����I�������	Gn��痋.k�nJ3�������P�nՌ����z�[՚�h�p�)����<�� ioӿS���>���e'3+����C9ل��b3]�H���M�n?��1$~����y����=m�J��V�tV�\R�UKR��0!���Nc-%/
�+'Og��{z��R���wû�@G]�Ì�ȱ@��)1ވO*�@�?)~w��up�ű��I�ظJ���%*�/q�ս�DL��W_Яq�n�m��n��Z�9ϊ�
��h���@��Qu_x�/��������!�.���Z��9�텪۱���F}�ǈ؞(uQս'+�aH���X�	gj������j#�E�Y��v� ���/�&�J��R�}4�LB��Pe���z��~	�d7��u�$Sɪh�[��+��{�����R��)W���M�[$K9Z6�Ҭn-Dv9��v
���-�\�}�/m���3ؘUXt(E��HC���g�$+������~�{��I�Tt�=S�z�[[-�3	�$AV�:����C|t8NU-LL����EOM?�y��Q�f
�D��[���GyEy���ġ��ч���S��T�W\�n�Ѝ�#�W*y�Sm�{���*њ^��WL�T�&y����/3o�΄P5yj�]G�t@<���j:�f�����±K�0n��\�Ag]�:q�O����iov��[8�0V۝Sї&��4��͡��&��W'd{��e4�x%5S�� �	4�qp<�
m
���,�tv���pP���1�ef��2�opUrf�}Fw�u|(U�����G��ou�~TgpeJ�Z��!��]'��(��u�>an�S�(����F �A��K!�NC�rp���V���;�5�ܥWO[O ~P҂[]kX�]��T����z���tw��LXJ�U�S'U��Z$v���x�*+����K�9����kUu����	���v�ł,�v��z~]t*��g���2��)l�7z~um�u�_�%rH�(�^�w-��1�b��,�k�Kޮ�K��G0a���7;���P�s$��ݵ�@泷�)9��p��n�퉡���yj��˿�Ttʋv�Gbze̜�5I�%�yg3[��/kbʻ��Έ��ҫfA3z�O22����b�Qf�*棣�t�g��W;��,�6�ܖN�f�i�*��׷�;]t����o��C-�e��=J�)C3��K��+38);�Bh*Òs�k����Ru�9]�Q���վ��{:@m���Ȫ��2��)��r�3ݝj��̟\�SYx��Z��]n��<G*�6<b�dA��׮�or�N�8��j��!�8���:��3��w��[֝Y�c8�&r��5m`8���aDI�k:���[�iS�Z{M�s����[2�7f��!�$zﺴ�b�}Ju�Y��Z��;��Mxv���Pˮ�'db/�v,79�j��X mX.�P��Q�U���3�&<�x{�`�;�}�:��<˽����r��6p�Պ`:S��d�*��]6�����xEoJ�|1g�R��ͅSs��Y�K���CD�']T��z�vF�j61�pr�D�Q}��t��9�F� K���M�D���}Y}rV�����^5a��X=̀2�-��w2X�f��3w6�Ҧ�A�PZ�>�a�E�A<e'�{��%^�̛�.L@�#���.�`��A���Ι)��._-}�Z9fl��r�6_iKq<1��3�q9�r`}0��H���d���jC����G���mkI��M�����S�oT�E@�Y8��w���G����+\�*�H����6������wk�7��V#�V&��2gD�}��V�w\{��O;�Go2�qm@yT�{�k+;�pi�V�.=	�Ʈ�V�Bj�nt�3ǰ�+��F���%��`JZ��#�a��[��;7W�=�XND������%�2��ui��X��gD�4S8�[IM���( �I�E�IIA�HMS25TT�BQ9�AIBRTM�&E!U4�M5J�PĔ��UISFf)C��P�UA@Y`%	ALA��PQ���KBP��UBdc)DAN�3%Dœ��aE0Df8FF2�DT98NH�@P�ST��bR�TfA��Tda�d�4�9	�UYbE�E.E%	JUU+@S��4�9d�RPD%%R��TLM)9�Kf8C1IKT�	E
d	a�TAE�R�e9���4�aA��^H���Ȅ�.�j��O+��*�H�0�f�)F���b��b+& �]3]Kmd�f��r�skm[�
o���I��m#����}3�/�ag�E�H�5⮝
�%���9z:���C���p���%3�y�r�1�X��m;z:(���8��XϢ*�S�uuʏ3	h����j��p���~e�h��m�󸹚��u�1ê�ZG�P:=�Z<�p���>�"�}��5=e�P��:7�"��1����s9�S��)}���:Gq�[���#�jJ�_��.��9!3�T�k)ߓ�{*����8��EUBK)VϦI�>����M	�0����*�؊�ɓ2j��C���W'������38!�If���/�N�t����xP�D(P;ԡ>E�v��~~P�2lE�ʎ*��y�:��h��c�o6��e１�(o�d�����*�g�!��R�����3H�ack���gm��Vԕ�iQ�3[I������$ ϟ��a��+�,lW�Km����^2�d�X祽��ҵ��gt�$�`��&c���z�����xN��`�p�	��ܾ��ǱdQ� ��(za�P��o�X�`��XxWj�lm�q�9K6S} :�u����0��,+���\ �\���T�l�ve"�����|:޳cp�f�X:����]K1M��c�ϐ{�mb���30+�Lr�Q{�ӹc��WPy�wl�����cթ=C�g��Y'��R��T�/��gI�F��J�cOa�CQ����c����v�Xe֭�.�yO6��c p�;\�ۀ
�s��3Ɵ��zb��/<�2G��m��r���GǙ#4����gÆ�!�f��*�z�zQ�,W=՝���f�l��,���[b�a������x���.�r�U��Cj~>�C7V.J�D���Y��K�|80�_�PV��^�h(q6���0���*~8d�2��Z__a��ՃKh�͎���K�L��Dg�6_�P©JzJ<NR�,!�M��~�=�'���"��hx-�;Ĉ��{f�S���*�84�HV��rX4Vɽ������guq+I�c�U��b��Ԅ��p��96Ȋzvu^ e>7W�t�7�Pޠ�&�%���N��0���Cb����eN�2������SQM>�z��N�;�y��5����5��痢tg�/hSn�*�Y��
�'��WW\�.E����;��ygir<��x��޶`]�P��:��z�Ӥe�BVC�"Hb <gD3�޵on٭]S�ީQԽ���d]�b��.�s�\���h���Q����$���OGi��gÒqd0���u:��]�P��u����&/�)��S�%��8�-�^�j災�\*Uc���{$S�L���W; �>i��VoOF��r�TO^_>q�,�-��ryZ��NW�����.UՉ�J��F�#��亃D�
��W2o]���jM���������9s:��e?B�hʒ�;N]M3(�>��I��۠�ϻ^���_.#�e_���xg�Q�3��PݖI����А�^���!J�w�5���n�-���D��Fx��|=�J��Yy�[UǄÝ�u��wQ�/�`��{��3;�G=���X �l�a���,(�l�h�j��I���I�o�֙��m��2%w=h�����X���#�ϴ��<�u=�U��exmD1�&oL�ty���X��*z{���MCu��%:��TQW��2����&|������b�t��}�q�۾N/lW��Dw'x��;7gu>��X�w�gP�<*S�T��s2�,���;���y+BE��4a���[/}C��܈�2�Uc@]R��z�@^�+�qe6%�PӇ��<�i�����esZ�M?n�O�K2� ɖۿz�a����E�@1���:�R��8T:b" ����h�2�W�J�*9��a�ˣ9�������Wh�M�t�_�y+���]G��dr�t�.8���v5Y+��ۙ��U%�B��@�<��m,��N��(��}Uea��߭AH;�К�!3P��ؙ�I����Lc��*��y'm����Ko�e^#Ƒ�u�]e��u�))C���%�0OuN�!Պ�K���$�o�)�i��Ӆ�b$v�H�A�=�<)�*q_V{2��s��K�D�����;�4�����©�yHb������;*b#����u��!��\�y�u����N9���ơ��[��e~�|y��hp���ϡ�<��;7�e.��"�|�&�}7�V`�����׷X�A}�§��ͷ�Ϫ,Z3�ܼ��0ҫԳLrk؎'��7����'=z�	�Y�}pE�%*�TU�@l8���Ф�z��G�[�0�'kϯ��`�t	gfm	�F.�B�z�%U��%/r�cϬ<�޲#�x n��`�'����+��x��E�#��]��<�/���UY|ue%!����=�v�e��l��l��[������%yy��A�NU�'+�QB��#="e�3ǽ��7�:&#O,�ZoZ���"C�:�@7Rĵ]�����s�ON_T����މV�w��k���6��R��͞#R�c��{:�0�/��E��lF���pN�ys���v���V�]��]�\yu^pCH^�L�P1���H^�\�IӽfH����t�F�]׉��**��JP�cOLO^xh�Z:�[�30ī*�y.u�߇[�xǖ¯{s������O��U�{1���{�<tjۃ��{aZ���Sx�}���4�jVk�ˮ�����ؠ������!�r�R$+�w#�t�e��n7�1t�w{ϛ7z�4�>dӠ��|�.��La��M��12����������yi�o���6�*�����;�M�5ߑ	�}Vu_u�}t�Q�B)C;E�˻T��`ޘ�Ζ7۠�v�%xd�^��í_�:�iJ��[��`\y�˦Nd��؎�So�D�%�b�8T�lGqs5��nL�8Q�,�	���f�G�5��2<��S���v+K]�tqӟF�>��圄>7qׇ
����vagr��䋮�ԏ�v����>r�)�{��id3i�]]Lt�pOO=�l�g�6,N�O�l]è���J�o�Q��4.%�Tz�yulE�L��MPV���}\�pb2���1����:�������S�s��#=����:V|nPs�ϭ�i�_pYH���c�2d+�n*ܱ����U<�gݦJ�/�T����ʀ�x�L�)��S&sU/��E�f�3��9al�j�&�[V\��̝]\֬
�b+���j���D�gA��^{M]
�!B�ԡ>�.���<�&U�6"�dqV�rl��޵kσ�睚ޏ=�:i��¤7�t��T����<	[IS���HJ�WS�yt/:�)�m�[�8����������I����ʣ����)�Y�r9VXخI�1.��Gv'�8��+���:<�03��t�$�`�"]AӖ����h��(������|6,�U�A��
�=����#t�O���'���x�K������ګ��Z���h���髇��(���4<k�����x����<<"�0�z��t����a�Ks��#Q�ϭñL��k
3���"��|]ϼn�f�=W�և���[yW3Q�HzMs��E�`���=�m/,�ϸ��E6�Tؼ�k�w��X_��
U�7�\��
�ATi��/9<����jϭ����S0=>����b���b�;),gҩ/&�]��:iz�7q�G띘�`��A��%�]���s22ߋ�7�X���A@�l��=��o�������r=��@7!y�z_^i���W+���תjOR2�7{�^4~r��m��:�-)��y�O���ё�X>�؀���7�����*e?8r��m;�՜�N�T���:=]��!���0��z>ޗ��Ի��V�fJsw��ι���`P���B_X����C`�=��N�����I��jo�9��̬=${�:�9�,���I���7���[R'S�"I��c�f���e�	����%f����ˤ;�P�D�`������,g�E4��ꂽ�Ȁ�8�|h��Pb��w~��Âf����#]١�
t �0ѭ�U��c>i��_�Y\�aƽK��we���UI����E<T�auO  U0X�; ���~!���ؿ\fq�y&���P�y��ˊ��KY����ZrK�yz��=W�,���`7��:L�;�!{�:5��`�fU
�^Fs�}a��:�&S�)V��,���*�s��(� �=��o���{�ne�4��\�*����}�D���%|0<�Rt3�,����:��S�E���{z�N�0�F��[$�=��.����n�*qK��+N�C7|�/;����'s�}n�=��yĞ�D	tt��}�lF��ie�G�W���w��x���]�D���fiH�rIVF��QاS܁�;z��R�1�\�m�u����[���,�Y��VD?xb�Y�{K�{P����i^]�!F*�iWZ�:��jJ��
�U6��{X��$�9*��.��Ȼ4P����H�r�w�Z�Lcs{��hh>�s�?���+�y�
V��Ac��L��Ip�KsƝ�5a+�����5|���I��i�KK�b}���n++:.%����J�u�v�xf#�XI��ļ��5���o�_�w>N��d��B��N�S�*�̯{��d��5q�z�w��w���D��;���ŷ�&���z
��U�F=\ >��&[���{��GB����뵷X����t�ӵ��U¬�����`�	�y܄��T���(PKj��^�=j	���C�-�T�n�m�M��0�`��WYj��lʤ��OE�5J�N �]��F\�����B������_8�H�Q"8*:.PTO
j�8�{2�����eq�v�6ݒVm����&�Ri3�s>ʫ�L�Nϩ�#BhX�ȡ����G�0�	���w�]���@/vv�%q�xOu���K���S[U�+a�u���4hj{b���]7��7��dĥt6�t�mҩ���~�%��h���*�X�E�K�f�#�������P�|��]Ɉ��Vv��:�=�E���)ƟM�,Q;E���\ݲ1�.��й8_�ֺ/\=�>K�n]�P���{׳���2D㷼7ۂ�T�;�Y`m���@�p�dA'b�;[i˳�����}W�ɋ7���p�+j���4-�"��bPr�T]�Ì�ʋ�P��=~]��^�^��mF���\�О��J���j���K<"Ԡ�^��4�����"#q'�wN۷����v�J�
�5V�.f�D%l&��tW�m-���8�~��x���ك$�4S���ާ��){��N|�}�b�ӕoIϺ 5,0��4�؞����2�����Q�d�s2t|�g+��1�gg'd_��&�����iΘ���
B�oyf}}�>O�S�w��F�\w�$�|<�f=>��r��xe��/���ad�L;CUj�Z�V${Z�ٽ�*]�Ω��#��~V���O+adw��D�yr�]��]��j�{[�A��<���s��ѼH���i�]z�Xp���M��VW���l�	�_Y|�'*V�r8v�f_�tU4�}��}{Y9A�,���$b!�y}�(������z�i�gOk���N�A�[qw8���^_M��ח��׈�
���eޣ5§�H=W���Z����P��΀���VKq���L����4��޶����d��7v�W�t��[rƧ�YJ%{��C�z�ǎ�+O���Ӧ��7��Y&�]��t1l�ޥ�J�
�p��z���a5��}�qT�@$���Nr4�L�ʕg�߄%}6�0��p�s�w3^�p����N"�htq _(��6�?P=��y3�����Ɯ���$�r�ب��FS5��>��aSϲa����pT�*�]k�B	�V����{^��<�"��,���]"�i���r��ϡ��U=;Pվ��a�f�[�y�F,�Vg7��Z�!����4=L�}@CÝ���W��}�°O+pf�x7�����j��x�{/�����K���Vz�b�Q��
�J�_h.�瞄ʰ&�#+qgaqt��K/vE�s�VK-��W�xT�􎪘�ܪ�@0� vxe�3s+��5o>����h�X�s��{�5�g2��D*�/!�����A����dXb�p�ۛ@4�<�k^9~C�l.������ǎ7�D�U%�EI��g�Xg�)��1(=|{4C��-5���MF͗�Vh�1TjY�nx=<92��$��)QR*t���37n_�����Κ��}R7�u�g�P���s�Lprסc��c#Ǉ�Z� g�]�ߝ�N�ϓ�⮭fU�Oo��Ȃ���jb����yB����Ƭ���V�^Q*t��b%�z��N,��s�睄U���]Ң�k���Y�v��9��6����JY���zl��|E�Rm�
��-��:��:ء[��6���8�@�;̈!����3��G�L�0���:���S�2��/M!�2�ƛ���4f^	1�n=�����uw�X
�>��#34̊�؃�v�y�Jc�`�k<�6���+.�QwM����Uޭ�[�]�����8%;m,nӪ�ٹ���˥Fz+j�,��q�u�#�&p����.eel�ծvn�ɤ�o^�^o˶���RX�gy�nK3K�b����]9]��G�L3oz�U���|�x�}�qbb�R�u���Y�iU��W���<��A��H,�f�[��.��c���lO���.K�ň��{I�s"��n^��Y�ɡJ|�F5]Ap"�#�l��4�;z��_Q˫�4>ki><�}�`}��0oag7%w�:)+v�)O&�#��xi�*N��ae�2�I�㤵v�\ܧ՘��h�<E�X�'"��/3��+ڒ+����,w<:�Ր����#e�O8�օS�F��I,��u�U-V��D�ma���lZ�T
S7��]�W�5(����plpzu�Ę�{�ӯ;Ú2P)U�Af �%��Yfzm�/�k����*f�����\2W�:��5�x�q����'!�`ފ�B��qQbp)��'�]�a{1�Lk�����}-ޕ�p�r�*(�\r'([W*���<RXCMέ��T�a=�L����H;H����u$�q�O.��z>�����o�3�Q�#��[�l(<�K�J����+��#�nT�y�up��P��g؀�R�7�r����W�Y)픧]%i YJ�=���q�t�Np*��^{M�.u�$�X���&������l��3by��}�n�P���ה�eE�9��]��W��F5�.��8�|z�_w`<X�&,�x0�y�>�G��3}�>�X��g,�7�j����y �{+f'|w��N�u]�n;V7m'5���q!�d�.�ӱpծe�4��Q']��� ��ܮ����V��-��R��R�Wl�ڽKn��Tفݝ�T`��aj�88uH��_6�*��2ș�h��'�	���eF�lE؜�hf��w�C�U��#�'�&s|{_m���KT�ᏺ��L��jw�5��v+��f��w��i:�aɕƌ7�y���B8�jzKV��vJ�*�0Q���d+��O5��M\z�k��)YrEi��Y�x7�G�p� ����]:�p�Ȗ�naI7�U���+�T�(�p��d�Vl��=�[�d�����Aܝpn⻶�5J�����5���$*��';-f�"���mi8ҫ̈1���{P[���bNd��un<f�h�e<�-C��3��
�2\����	�2�����(2��L��*2p�����(
"�3i���)��j�'"�����2h���j 	�������hk$2�����b�
,�,���,��3*�)�*�������c++ �ʄ¤i2̧*��1�Ɍ�"i�%����\� ���rrih�k�i�11�����)�ʃ*2L�K1H����)
(��'3
�Z�p�����Ĥ̱�+!��J(��$��*�2
/�4���>�U��э,�k�x�ג�}�髃�+�hHz��a�A�|KV�y��2f�lU��/�!"��^�v�<�x�t:�(�Eӱ]�: �[q����ئW��(�e3�W��)��d=���^��a�U�X�r.�累4x)��(xg���������ͽ�`�f�D��J^u��u½t��o�������?+ɭR0����'�i��>Z��mL>�`zs�F�����`83����FL"�m�k���f{[�VA��)7���b���a����[��{�'��0{]b�+��AA\�f�^�=�zd��ʹQ���ēڥ]���Hl{fP�51����]&i�ŲWZvu��	�D���t!�'I�����<˰ݵ!#>�.��M�Rdw�{�&�g�WΝ���y�uv�ͤ���I�K��*��S'�X'a�f�<V�c�i��PW�*�>y���v�voq�ܵ�
F�'.�*�Y��hU��]��F��.E�7��k��ۥEy<���~�.޾��[�����Rs���"�+�<�̞@A gu�Ш:A��W��86�ڞ�;�]V���vqzf	�c{"��(��C��0��z�U0YCs��{M�C�:VOf��r��.�ۊ�4B([�=��䴟W�u��&�j�MF)���v�#n�u' ���0ͽ��$���H�*I������0�KZ:vr��23ۜOL���O}���3k:5����xy{t��j��fPJm�v_hnj��E1O�
���x���O�g2�:�,�N��>�]�C�kG�y�ؖ3�:���En�%�ja����B��!��q���(8`y
N�h�=��=�p�ߟ�g�E]�P��u�b$�f���K�E�U�*�oR�1�=�������}�d)�o6}�Ā2�׸��:� _t�<�媗��#�0����g���{���a�Ɩ�'F秥uv5'�p0__���	�����	X��]�%�n��~�l�^bέ���OQ�=���#)��W�ʆP�^q2r��Ɏ�C�v�xf#�emAv3�)}�/1��ğp^;.�d����)C��
����9}��H�����l��y�;Zq���u�R��*Ǫ-lJ�C)j�\��u\�eS�� �'}n,��b�o�(�VgZ�y���5�r�7���J3��+�[*ϑ�_�n��p��	u5A[��,�{������:�ץC|���pY�z/�3��
�:���Y�Y��V�Js�+���W�J{A��uة�%�6�&�A�˓��j�����j�ϔ��:�w(�qC�\��u���8�X����o�t�q��q�۩R�K��<z^2��æ�����<fBi�خ"��b���V�xZ�BʙBp"X9�*[��'�_t��<���>�5����^�8ʙdr���|t\�
`
�E�0����C����3�ldN_u�z����J����[���1�UD,�f��~�Ƣ�y3~��4J4kDTv�r����;�e�߇Gt��簨`�}3+�����z=���6�ʼ��[�\3;��Td��C�E���
�4筸�Ϫ,Z)������c�ܿJ��6EJ�陕u"�C�!��n�k��v��� 6e��}(�+@7[/����VR��P�*x�����_�#z�'��|߆ީ��oݨt^nɹi�.��'g�`u旈���g��d�[�3�u�v*�5:�a���Ĥ5��%0�ӈǾ�;�&Ϫ�_
ݓ�D�.��,:�[�s���E.#="e����>����9�(k���3���3:����0����ΗJ�ux�@x=�PO3ň��=�,�Iϯe.��_��u^3�'ʮ�<���нQފ_V�J��&K������Ӑ�*ٹ��N���M[���e�8�Jc��#�KՂrМ��lG���TUl�T�nP]�Kf���d�^K���S����o.f��o�N��[��oF�h���؆�b���Vm��֡��s2lK�� �]�q�v!�5173�}ӊ���۳8=.�H~Ֆx��8eV�	���D�_^	�H��]+��}=�3�Y�q�>)�稉�%�:.-f�����*��,W�����t<48H{=�ڼm�(��};��_(yuH�Tj��Ͻ��M�5���G���Y�i��ZZ��Ez�+���Zˇ�������b�d�bu�8����yxw��)FF����䱟Y��9r����}�9;���S�uu����Ol��D끙|�9���c�^���Á�TW;\��|��J9O�&TD�}|��P���a_O>ɇ�C\�eN
��y�V�y��<'����?�JČ(��)U�C�]"�ƐyM*~5�N���چ�<��Wk�
-F}�s�s}�R:�������Hн<L��[*�؋��d̚��R��j9���(lI�?d�>��N�=�7Sf��\�n��=�B;!B�z�'Ⱦ.�A1�����>2e���{���70�^}u��4w������Ep{jy ªF���UYp���a\��z곭wq͈��)Hz�]#���n�%�J�;�����j�<|�.�ͮu�rC����xw�j�H:�A�Zi
�-�ytH}(��Z� �j� *��
�q���m3}��q�*�$opr��l�c���T��{r�}ÌW�͗o���镾et>�u�s#�D*��~��H-��]A�bB��d!��b���JG�sώZ�*Y�#�R��Jj���3�eW�\W�f:NXg���fM�W�=�:�}����|�_p�Z6rW *
���[���]��xr0wK$��J��S���l��`ѱ�~s�_����3e�+q&2������Ӫ<�YC�qz7\��=�i� ���^�9�:;�{�2j�*oɰg�e��5�⬦wo�Ph�0R�!{�3��4Jٗ��y�|=S�QxM��8���#W�Se{����mSb�q+��)��~��OzǕ��>�ف����pKhc5�eb��ʶ�U3ӕ������O��a�x=���o
z�Qz���J�|���"
vOZ���w+��"q���_�P���n�A ��zd�Jս��O��Qd�v��<Qu]���Hl��a_C���ϰϐ~��o���<��5ʮ�i��|L����7��(�ymHH�L=6Ȟ��԰Y���\�\b��,�ЮҳZ<)�s�N�t�Z�2�űК��^]�O��,q��w���^gj�Ќe����!�uu��eʡ�{	�$jK�p�w]�V�8���,��]t���Mf���DIw�:����T��vŘ�Y;l�I��GCg}��}�*`��lV��x�@�m���[E�r牽�}�n�SF�{Τ�_�z+g��S<���q���h��djic�:O32��p��.j����q{8䶏,��Uz�A�~���*�����d�x�O&3'�*�,�v@l���y	<�n�Z�3��}̠��/Lϧ���פv}
�`H���r��L
S�xf̶��gr�J>b�L'�wu��޿���03����e?B�h�,�������cwä�8ygo��9RZ$��5�mD�Z��.�j>�z� ����L��eXC׏���ǔ$R��r]tn�b$�ͣ�-yh�J�e8����]K$h�T7'@��w{��Ҡ毈2�;pƛ k�lЁ�yj�rvʶ���=�����-�	3�״��%�3��@����g��/)[G�kR��<"�/�����������If�(���,+��}e�iֹ�k�Y�̨/O#)��W��e9l��|7L'� S�f���ק>j;�����x�뺀k���ڪi�4S ̢�4�]�X��J���["��l��Z&s�q}��fGB.��#{�:��v���{Dm���y1cn<�/�:�N�\x�@]u�mY���X�m���n�Y:7qP5�C��S�����˶��D���w��V�|em󻂖�)�z�ß[���%dj�oM��OgG����ϻ}]ˢ���H]"�[߮�&���+�h�d!��@��&}n,���{��.�eO9q�Ƥ;��_:ȣ>.�h�ţl�W��Aqu��n3��''Q��X�K�#N^�ݻ7�>f��cj1{�#u^#Ƒ�����EVz7�+0�{�z,[�C>}+�^&}�_�>�"��Z ��w�_��{l�� E����+�%b���Z���;vk���Q*ܷ1��7}��"=�)����[���Y$B�����L�OO.�]"0���t��y�d�/�Ђc��>�P�c�v����^�7ø>]�����h\�0�WlFr�W[�<�t���Jg�-��|F^�Ys��ޜs;2C�;Y�ҕs��[Ȏ%�.P5wmv�����*�b2��藴��R4�9r�oF�rxpn;�����e]F��Y�_�������{�12!��w+�x�鶷&�Q�y`�6�>*�]雌r��ft��Q����B�r�;b�h%�b�:�#�^��1jsC��yrޣn<��}�Y^���� 웼5U�r��U'wT�����ItT��I�P���d��z�3�wI��c}s~Ƀv]I�`��>�V���\�cD<�x pd�[�!�=	��]N��}e���t\�.sm���Ǒ����C�I�L�W�y!��B���ʷ��WD�����Fzh���2F���<#��6ݍV챰��߂[�!�n�ewEZNk�����d���cNt�40��v��=�u��q���I�P+������d�/g���=�Gz)k����ٌ��nL��w��[���#Nid���c���vk���/>�~���á21yh��.^�60M�f\��Ǘn��g��/'K�v��lL~Zv��E��u)H[�^���Ǌ9��_E�����&&��3�Q�zk>�j>�������Y�iu�B�sܽ��Y�2˯P�^�PϞ��U�bs�\U�M��ު^\^"8*:.	�&��޳�c7����u�J�����b�ن��;��\�.f�8]{rf1���`w�NN'<_�w]��,Э���u/�Pe��:p�9�h��3��9|l|s�WtAC��!��}-PS���8;mc�/-�z9�퉗;f9�BƝ�p���u2b�}:�孪g�(�J�[�{g�ۧ����yev⠩T{1[\�×J�����*'�:�n�T .BS$����v�G��W��P��-7+.����7U����yS0��Y��õtX��ƐyTҧ�X��͸ �C�`<��� �Iy�]�x1z�8��@р
����<L��[�bv[&?[�7{J}j�����y�ћ����	��p^ȞS�t(V�a6|]���ըSf��{Sy��2��N���f��8�_���h�3sP��#>��ʞ@0� k'��]t&]]��y�斁�j%R^�T�Ӭ3�U�!T����)>>�ZY.���Ą�B�br���->��G�4�{.���x����!��D�R\W�f:�z�� i����ҽx��h��xp���)@�r�o���-v|�m?"#\�'�����xl�kz��ļ�!P'k�%{�C�s<7��}�K3YTz�TLpN[��[���T�OZ^�RC�\Ǻ��gVǠ��v\�_��)��,��Nx���Ѕ�K�g�M��&����Y�<-�]pM]FC�ʼ��j�L��99m7oʲ�(���m�ח�׫���X�oE�s�]�sJ�̜e�H�ǖ`7uj=xI�&뮔޶y����2-՛'?<�f ��H⬩1!j�mj�Q�@M����S6��.YrY��o(9�u�$2�9]�pU��,��gGU��<���H�)�@�V����M�*��|F(B��]M)��9��M^:�ޫ3�U¯�'C8��+*��&[S��f�*����J/��~�{3�����y�L�r,���w�`K<x�4���WW]���_w��}M|�.%�]q=>��{W�X��wzԑ�i�Xl_��0����	� ;�Wz�l����5=���g���$c���2��
���5wCM��d'���f�<�>��$d�u<_{,c.�(pJ�o=����#'ٺ��z����X��f����H��^'a�N�|���z���\�������޳6�諾�B�o8�uS��ÿ���z"1�a���4����k��`]1j�׼��ti���G�TQM>��{�KU������^�y1�S�T�`I��Y��8���s»���%
��F�����Tg�c�)���-f�p����SI�Fy=�����������X��ȶ��U��U
cn�a�ϐg2�:�&S�)V��;~չ:�z;u���m�����IN#]��N��K�ƣ�g����I}W��;��l���ej��Vv]���MĮu��Iۢ6 Hj�Tu�`�Qk�"TsxKH���u��̽�W�p�����` �r�v%=w�	�3{������� �D9|�7�hZM@���d��2����� 2�T�ue��;�4�پ�0�8� J;9}������S���Î��^��b�e��Ú���V�3�����=�Q_r�����vg5`G˃�V9`U��k��\�=��&�{�%w]c�J��_+��;U����c[����5����7r�:F̹BjQ�/Yϯ�^�K-e�]��#V>�O,(�z�n�|Vrm���b�{�mh�y[�K0���s�x�&�v�;���I˾��W�p6�Ϋ(��v��ꏷI�i���bR�<�\��`�(���-�
�`��]�ūU��9v2*�O1�,�3	�4�x���ᡝ��Ze����e~e������=~�!n��f]Ϭh�-�Wڱ�m�nB�߮�h�2-7|7 D=5o�����Nӹ��@򦈢�i�sY�N�rip��m�x��κ ��y��˳l�����s��aǵ�	wA+̵�t�Ue ���I6�u�ݭp#[�j���h[A�/VT�A��;�b�(�)��{�^<��Tm�)Sw��U�i�Ά�Q9�)��T��W�q_ZӶE�Kk�hC@�O�=W�"S<����<��ܽ��w-�QC/��d�u���ݪN��}y$+%YMi:��M��AY]\>���;�:�ҍ��\�fgo�5
۔�!����G�c���c�L���v��`�}ں��
hQ��ʺ�U�b�u��Wï����rV��o=��lt�fKɕm�Ov��p�\��+����O����b׿~G(mi�GN
�W5Ԧ'��΋h�z��Ӕ�f��ݚ�P�/ 嵖�GCo��jG5��̾�ս1
Y�O
�tR9�tO�p�U���A��f�\d�u}����]�'K�k�g�X���t%�^f9ܻ'd㡽oW;����R�T�}2�"{N����˵�H��Z����
���q�\/��	w��< SRͼ�6%�wz����h���.�ث&�s�oåf�ݩ$/X6��u���bdogP&t������I����Z.\¤V�զN|����;�;�"�٘*Q�C���1�.�)�q,b�p��N��o$[�r� ���d���I�Q�<�sV���1*�[�T�I&Ε)�9�䊦����ۺC����tx:f�2����\9y�۶��T��/��&��^�t;�*N˱k.Ph�N��8�
�4aO������ܳ��1��mK�jA��1�����ձ�ևλ�.��h��;|7�$�\9>�\֯>�]�0ɦ��}K�\V���G+vw�5��û�r}3op��1.ȭ������:^t��0�F�����K2;k�N5r^�������Y[{z�ce���יy﹣Ϻ����`Y��Q��Y�AT�eFA���feE�d9�d�RU�e�e�-�&N�X�e��VeS�eY8A�cTd&FQ�d�U�fd��X�TS�FI���PіfYX�9YF4QTS�d��FT�fcL�-��a�d�5���d�Vc��fYfeR�Q��Y��faS��FYd�44�Q�4�e�Ud9�)�F1�F@Ӆ�S�D��FAFIe�3C�Y��E�FfDTQT�fE�3VX�1%5��e����T�NXf&Yd��QNFY�`e�Qd�aUS�fc�f9CNY.f��U�Ddٔ�f�a�fQXFY��VFae�e�k3X���>���������e�BgVu���R,G�_^sn�LI餉lܹ�͔պ�fq}��_l]|��F/y�n��#c�x��:+�#��T�x:���/���ۮ
�R�pv���s(K_�o������gޜ�+�s )�F@r� oK�媙�Gƞ}]W�1D/i?->Zl�f�>�˱s�"����[~�����(����*"�N�@U�Y^X�;*����h��3n�N�mt�m���I�K��=��ݎ��-����R�^�>�P�U�'�-�޸4@�+)���Ұ}kԶA�W�&�=a'����t\R�|����A-��o���f|z&��r��K��n�)����ȭ��!uH�����i��`���Q����� ,Ei�_�z�B�;�c$/ݧ!ӂ�4�pPtX�1:/�\);�К�,ػ�`�[i�	�#���+�AH��S8�5uh�KY�jS>E��i��=�"�����Ur4μ�{˕��
����`�-����D��� ~�����H�Ɲx�9�J�ڻ^3%f����]	���%S*�c'(n&��v�甆){޷c\�G
��R^]ߧ��X���+[	}1�n�K���k�K�f��x����ˬ�|�K�VG�v��`�N��ߵa�*jQO�!O2���^�xmuK�n���Z��nHu�0�ۘrJ��(@��3Q�r�*��=����b��p]v`�d��#�g �$S;�]� ���#��ѮQ�4�)�K'̿:;��Oo;�����NRs����ދ�� �+�����L$�#&�
{�<��9���Y��b�dʛF�J��9�E�m<>�b�i���쮌�[Ȏ%����S~��Ȁ��:ժ��N���_�[�;��g�&;�2��u�2�2�����W�_Y��Pv�*�l���fg�닯��f�P����헂��d��#%��ب ��J��e�<W���Ղ5�q�\�3�w�D1�C��u�ܰNw�*�*b��.�f������S.�}-�zn�I���KԬE}fgp��/j�u]�����w�@��pU�r����g�Ƚ�2l��)矸�3SC`���Q�=�>�[���"��2���S\�X�3#o�d>��gT��-�}�K�~�6����E�z��Z�f�}��}}h{V�
��L��萈��gc�����}q�W�i��~��~�/ᓥ�:.-f�?-9Zt�}g�%TX��)ۦ=�����L��$�B;��_�tye��N5�X	���Ι�v�sTP*6����R�kWwu\����ՠ.qV0o9�K*��;��3Gb����K��h��v��u>x�ݻ0��e����K��8���
Y ��m��5y��Ga�q�4�G-gJ����T=U�wp�Ćlj���w;mM�4呂S�j�w�6N�V:��cΞSk��Ř�@�4t2��\��b*���X:o;nގ�24
���,��8b����^���6UߑyVn��r��}��%=�9U7�|�>w3^��.��xn�ٺ�Qn���3�!cԠ^�>!��C$�K�T��uE�4�ѣ�]7�K^c6^7���/d��1i��z��
��T�:Gz���ʺ,EX�+�?�~Nm����«��E}��	�ݞ�.g��@�U.$h]i�eTz�yUulE�L�����Eх{�Ӻ=�Z�)�[~X6\Z9���38/}�<9AP��
�N��yP�'[Lvi�o'p���t�����e�i�k�K������xT��J�@1�0��^��3��b�מ��P&�K�Ct�1��F����`ׄ������AhuCP{4�Z99�f���/��`$@�L$A�^��ax���)�L�J�K���1��J�.r�ǫ�S�z:��Ғ�	����*+~5��s��� L�+OF9�Ǣ���U��+���=�O��ٔ�I�Squ��2�_建cB�up�uX�Z��8����ZWd�ĭQ�ݙ.���.�=�4D2����wк�v�og\����E�����ip��h���@�pb:�?.�X����|����������,y~�4W3�|N�4�ĠxN�`{Mix�c~X���k��T�U㡯N�urm�"'�U�`|�@9������U6��UVS;�~ʃg�1�×��#?C��C����'x?U��ߪ�x�Aw�\�3����v�j��/Ww��Yq�N$�^ç�g�:�u�AVWT.�8%3Ӟ�A[�Qxxo
98���^�ŗ�%�f�D����%�OU��`�t;ĳ5�}nfA�JVU��?R,�ַr�U��*�T�<E��qĖ�/ .���Dw;�3�^A[�F��޾�6��E�!�==���A3M}wCH&CﯭA���D��jB@�o�5ms���}:_��o#O�dy�x������f��H?+'I���DV����~�cn=i߯���A\���o<)/L"�c�����t�U2���4*�
t%	�P��3�mo.ѓ�N�=]��ֆ�W&����{S����=���6ݷ��\�trǗ<}�=�wc'�<��Dͭ��3���N�>��	�f�wIi�y4ʓ9Kߚ�c��+Lݮft#U��ѥo+�`ꊷ�\\��̀�9ffa�ͅ�Z��5.%��qf�Fz�뚪�ȱ�4���7-W
Rs��{$S�zy1�S�;}������8��#�>�[��x� J�\$Tj�Û��g|d��V�KY�����$����!^��Ai�p�tTNu]�,a�RU~�HϺYd��خ����l9����w��7�\/�5,�n�@�q9��m�wL<%w�fX2�	h��5�s���]K���g�z��F͜�X���Õ+Z�$Ϩo��2���IdV�NX�j�}xJү�wu§�gc��p,��=^���+��;� ��� �wQ��l ������U2����Ϻ�|gt���i�#i��r���g_{ګ!�-�a��ph+�jP!yǄe	��9�D_Աex �	�о��L]���c.0m��W�J��_Ksƥ�u�Y�z���ʆP�U�'=<���K<�xe[4��1����b=��VY�Wq�߮�4�}qJ�wpR��A�|:���*��H���s��}�8p��6L�8��;;�T��-tJǡ<p��T���F�<��2,$�>wZ�B*~��`�n��ߝy��htsNt�KZ���k��}6��]�nm@����M��6	���ԩ��}���H���Q4o�BH�D�7�[#:룍�]��)�76*Y��Ӄ"*��&fJ��u.�|ֹ���֪�]��:��xB:���a�0�A��UY�3*��W�n�F���
�>���[t�=�Lۂ���S��ɶ��/x��.��xң�����T6�,�zA���y�2w���fϒt8`a��E�7Ӱ��yV�2��]�υ�re�2�ل@��7۳C���=�8�,���TH�ͻ���2]���};�Os�B����p[��!�/���=��9�Z[�#�bγ@��Q�\��i��1���^��Ҟ�Ö�YĨX>o��rIRUnkYCT˱�ne)^�hs&K�tX���
�4筺�A���{S.;7s���}ٚ��<����[>�x�Lz)f�;������\�k��j�Yt�Eݖ$oz5���W��Qb����jY�S.
�L��$oQd�˓����cn��\.���#g���jT�/w��
t�L��H-��K�6*<���:I�Q���r�q�~��Ӗ|���U7�4����w����D�����A9V������QW�J�#�E�eMc"���xXE;B���>���O{�����m�P�q&1��5�P�@�����_<c��7j�z�i�h<�qiZw6��9v�:���z�p�����9�g���𻥻�ah�5 ���:_f���#9���C|�;���8���}'�#{��{��i�,fdY���tC	΁;e�W@���x�\����3U,f�V��V��(Vȯ�9�d}e�I�x{�c���o$��^ڱ��N����0�w�L��ʘv�ڥh�X�t����ʸ�:��ژ��2�:������@;���׃d�
�y�uc'K�t\Z̶��N��l"�z�R-W�3n-�r�[�ڬ>��B����s���%x��NU-LL�3�������k'(8呃��Z�vJ��n�d�G�ΑCO��C}MAO(�2|8I��8����yxw��{Dc����Hv��ξ�[͈�����z"��`!�]P��a���f�z�5*�����y�,W�)뜟LO^R`'�C8��t�x�Ih�i
ө�u��f�T�0��V��ﴶ���@�c�3w쵙���*T੊U���:Gx��4�ʦ�?�{C��P�{]�7]��&˂;\����#*�.$h^�&PTz�yul@7�������9J�@�}|i�>���쎯���X���[�õ�P��8d��쾮�{��Y$�w��X"���8�Zy�)M�u:��9�vg
��up��R͈�dA�(P]:l����z9T��
�%N^�ŭH�.>���Lm���d'��p�7ֳ��<��eY&g��x*١B��J1^�N��4����E���e���)f	��4㊵��y�;���<<$+�Ϧ(6e�����B_��dn_N��T%�.��FC<��m�R�7bt�k�H����������?jm��t��7^�=�3"��G����yKm���܄9��(�����>3�f��}��^���B}��V}"B������ѳ�Z��+�V��:�y,v|tr01�^i��`�v4���W5zI��J����A}N_��}U�����g�gڀ�4��ʥʤ�ݻ3�c/�%�wW=�קD��<<&��;������z�;���XQ�*��w\����Qg�ܧ%�\�
����o�C���P'z=*�x�CW{�����U�&�6�D+����V�qGe��ާ]��ڭ+AW�t2���+)jbe[S�����F��#��<g����뾔��=WaXw�1�3��K�	OR�N���0���.�r�J�r`ό,�LWb_;n�1o[� �bE�آkp��V^sVӺ��+n�ɷ���t�r:+ݤy������w�I'}��2��Pɔ��{�l���sUC�Z�Ԕ��#��DW{CYܝǫZ7�ME@h����)��3�}�U=�[�R>��㗷�����m<��|��m�\*�a�:�E����}I-� /�\ /��C`��r���8w����3���Fa�52����­g(&i��aD�>�1�����ӐT}6ݸ�s�Ɩ��<��x��")��c=������.��%��v�ctup�'){;^w�|�#�"�i��gT�C�^��9��颦Y��F�\��Z�^�xO�0��nsY��b�	�1��uu�b�`v�x�K������I�3VH���l/	otO[cG���{�i��ox	�u��
���p��*��=�TS+\6�i�Ct���.|y�n{wT瀒t�fz��4o�_��3��J��+���Lnl+�{c�Oof�K����a�n�.�0�<�Q��G�E����`R�-\&�����]J��!���.�S�+�n�m�[�����Ȓ��ۡ�%�[A9c�;��;D����'Y��>Q���)v����\�����[���j}�V��� /��`���-T쳆�}U�t����m���l��;�MOý�t��`�L�16j��z�2�"V�Gt9�&'Eи֮~�yy�׭S���o���ͨ���T4k����}��	��Z�$�ס�ev��WG��-q�go6BэY}k���굹**��nS���t������8M�CQv�5*��U��m�fխJ*����;�J���G��{s�>�m��9{-]r��yߑ�(��#��Y}�ז��9P��&N�I��߻����q�
{����B��+,�j�i�K�I�eh�wpR��A�|:`1��*e�������[0�s�)���AB��E�%aw�����%)^���hlZښ����>~T��S��OX��=4��t/O����at�e}g�̫����ו��N�o��{r�gpͥ5c��Bn)A�c��6�����ʭ#ƕQ�`Q�.�&�}1�����u�)-���OE�6r"9�Z ��w��.e��2E�FK�'n�o����@v��N�h�\ʥ��猜����v�{�R��z��33�e���n������	�`]s�Tƍpj�Y��}�9-��t
s�πPF��~�z��	�n�>��e�α����j&��OY��{�h�cG�-��G�y���Q�"�
����
��ED�W�(����ED�Њ�+��TA_�(����TA_�QQʊ�+�WTA^�W�(����ED�
* ��QQҊ�+�����(����1AY&SY6�� ʨ_�rYc��=�ݐ?���a_��  
P(	@�R�
 !   �J@�U+�� J"PT��B���DPS��QIPJ����UQR�	*U@�J����J��.��� 㡈UJJ)lCJ� u� ���h
� wg �R�� ۻ���\�AѢF�-�6Tʂ�ff��44t 4�IAX .�p  'w    0   f  �]���N�)ͅ�21��:wwf�Y��Q�@8w:tuj��TkM3�D1P�'fB���ȶai�*�1%*\�҅A)T��"i�U��+ZT�5TD�Q
�p�U\�"������ɬ���kM�4iT)T� ��l�DE�I"ٶͥ����U&�ͳm����j��QW c�!�Z�mʨ��h�J50�h֛Y��mLB� ��M�F!�IS-T")[2��keCR���ԂZD+�#���lb�kl0����0�T���\�    "c!�)*@h�M�h��"���)hM �14�bhɉ�	���0 �`�0��~%I)��hh   �  9�&& &#4���d�#�H��1'���##@��c$��ߩ~��g�����~�8Խ]�p�zJ�zkE�� Is��	�됐 I��IBMI$�!���$�O�I�$o�������hl?ќ���j@�D��#$@�����$P�!$����������G۟wː� f�.n��?57>ֿ�)����)D_�N��g�G�B;�_�R����/+i ��,�<�q=�k�ޠ�m_Km��O+�7M�f`E�M�7�C*Q�tۼٕu3
y����3Uv���ۍ<VT�ې����c7l+EnY6��Ag6�d����U�f��l4����ڭ�Ȣ��v�Qm�zG��5˟f��k�O6��r�7A��6��¨'�7��f�u�SJ�2��dT�a�TPy2n���U0�2A��7�)�'4b��x���"1�Wn����6�Hܼ��:�aXbm�d<	;�N��GU�̋ܚE�"����nm���$^�F�.㛫J!�C:��J��5��F�'��hY��68k,=1���4t9���ɹ��
l�jy�M�e��敊������2���2�J��E�fZ�eM3sv���,�E��6����@�![�hyW��ͻ��V�'oA��y�"6���f��[�2B]c�Y�	;/X�CI�a7�.�:���&i2�G3/R���Z�A-׺�U�0'W"
�HU�'M��������V�ֲfP["kA���cLY�WlQVdʺ�)ϳV,nL5`�����oK[���&`2ʼ�f���Y-Y�h������&�@̍�趱+Ԇ���1W�v-uTެ��2Xr�Z�D[+h�ś{��(�k�М��/&����A��e:��tm��Q5J��4�\��V�%5u��ٯ
��T����+26�ެ�&=��
���/,��KAU��K�����ɴ`�5����Z���E�y$�]��b����bpѤ�n�Wۊ�h�����X�P�w�%j��]�R�Q��j�1YBX����7X�8��e,�4ZcP�T�V�����b'�5��n���;�kpaK	�Rp�WoML�Ub��R�[5�fnE��r�𻵯k�6�-�Kb:�j�UK�i�A�F�t�c�˞�˴�H�j�j��C��_5��Yf��hZ�,2��wzj��y�N`�̧Z���rY�Ǜ��)���=4Uo]��0��x����o�oZi�B��+<K Iڦ)/7M�X�s�ۡM�8���Ø�4�a�֭R�Q�X���K�c'��
��i�E��V����8n�q�wK�؍��h��U�G*	e�hk��U�*���WSa�U�fե���N�I�6NT��������i�B��w������f�/,�����r�H�����']�;G�3#�y3j���vn�|å@Yt��2s/p�ҁ�֝�u�cG,`׺.�̈́Ji�ˣ.���Dnӥa�*�=��Cj)�b�Tݶ��	�ڥr��1���]��H,���tڂ��[0�6�nfU%]��y
�p�)����ң�6'w���j�і�@�Vk��<8�:�W��������$�!z���E#�]}�ܓ1����J�]��I��'B���a� �^C��cs)Unغ	���P���J��n��%"�P�l.��]J�!�k6��"�������2-�g9�ݸ����#q��kw�V����ĭ4��Zǋ6j2e��C�1x$��Aw{f��F�n^���C�r�H4�	�JX���R,�#ʢ��չZ5f\Wv�FjK��m<Ӧ��I��H����%-��Bj�n���fVJ{C(^o]L�tM�)[z̽ȴ�D�
�s-+^�
v�f�4���߉t�w�,���3`n��+VҧX��x�w�7E�Z��%�hޑ�!���K���,M���1i9�zC���I42�[�9ue�1��P�|Hf�	p#���	r�k��֧ʷwe��+-9����.)r5��gZ[���J�6�9��<�yyoP�B�]oq֚޵e<�]]W�,"���V�"+(�/l�34^n�����D**˥NM�wF^H��24E�J�Z/r;�P�Bњ�[V�S��ĭ�^��4�+8IJ��Q�{��<x�uUmh�%V�����Cc�׷TV�B�Jn�8��I�a�D�8S�h��۽՘�7M5u{c�C���pƇ4�<xq�T\w4���9����Q��5;
��-\��H�cQ�9z �t�#�iȜ���M1ʃ4��unX�V-]���l]�'.��VQ�K)1���/��f���k9Q��7��X+�:��[0^�o�8&����PԌ�[��1/�![e�b�:B��-�x��xP��Y��ȄvRܔs�o+g*ޭ�^��RY�l@��B�S�,���re40n w�gF���"�h��M�b��5�[���5NT��X�Ӥ�y:C���*�Y��ì�h�Q�4/4�Q!FG�-�r���[�S�خ�bD�8ۻ��t
S*�����m�q���D���H���5�J��vP��vU`��R�|��A$�D�L_-������1�P�J%5GJ��,�Olڳ���T��f<e�X���w1M�!��r��mXЪR���5�lR�H�Y��B#j��@�5�$(m�(����B�a�{�$�Ǘ�HG���3A�@������s�����|�U��>R����f��ȃ��ê�EMX�5c�ΧWF�]�1觵S7�z�2%��V�u"�ј�7Z3�Cn�yy4��7�l�����VR�)�d[.LS+�yYr�#�]٥GOV�F�k�'IZ�čخ��m����ܖ�.A^�j��������� �+S��C>Dn^7��0�mӦ�ukB(���V��ڮ��ȦC3�:E�,h�(�V�ea�S��ȻT-U��h��ل��S
if.w3wv�����H���Y6�܏9a��Xv��!F�l`˗f��]&)�ʭP���y���X���0�.�2�����]��Pfm,Q*���p馘k~���ǆ�=���S7������LkX��̸(CF��Ve5Vn��m̻�b�L�\6��*�]9�H�v��۳�յOTہ�c�elX+I�R��O2*�nQVV����+�xŗ�V��ևYyt�솄˻+�F��l�;U�5�2}WJ�t1f4�LuiVܭl�T%�ҘX�,m�Oi��^�2G�U�a���m���Q����8D��;�I�nUk4C��1Nn��t oXʭ)֍�5e�v�� �䧹x�ֵ=�������U*EW�f^]�&�i���Lջ��E/����5NԢQ3�h��"�X%zU��N`���ÓK���Ⱆ�Aa�����+X�:Mۺ��]���n�ܳ,�
їn�ޣ#�ￏ�����C���t��S�"}'�������>>���.\̹Ɋ�����| �1Hn�%l��eT1��*=(	E:�*\KVL�Q��\Q"j�''�U4�y�p.��B�ٖs4:�Й��CNz��	&^�u�6���k�ٿ����{\U|p�Es���K�����!��0�4.�&��Y�:FO�QB_^��N��pJ�b�P�zA�0���p�*�fcn�ǹ�PbWUk�N}B7���Wkhd�����$�Vz,�Lˬ@��Jp�/Ki%�2]2��G@�f����P�n�0�l{<���Q't�K��o"����E�o�):Q�j[��
�����G4�T���k���=S�e�;I�J3o`�k+�L;�]�i.�$o��K�L�f�[W��)�ow�����.�G~�yu|���$��s�u]���;� �jVvi���c��e�Ic�K�h��Lw^,��l5`�3�����Գ��]-�ή�$CV^�*��^e�х,��T׽�2B52PW��e�F�����}qK�9X�ÚB����ڷ����4�<z����@౫�N['-�_mÔ�o+�vf�v����dp�!�k\��M���ds/)ڣA[��}�JR]�7��F��>���k��؃�I٫d�[Y�U>7�;���ES���W$	��M9���n�K�,���Ghv2k��)�2�̽���.����ɛb���X�4 �����kj)	7�eM�Ih�vN{�4S���֊ޜ����j,yB����
�9J�#�n\�<��ʲⓉ<�^9��ȏ��_*�<%��r�\�N��f�
(:��3K�B��^�}�T�-���5��r���*&�O���vAp������,@����Ky@�I9��nܮ�,��1֬�I���Π�'�ne����+o^��=��BMp�������I�J*�[�������t�1 �S-5�{O��]�1[Ǫ����1&T��{8>��X�r{0*�v�����T7S4k�ӫD���|�Ǜ��d���T.=�O���w7��#JZ�~Œ��w�=���h�:��Q�6�y$lE	��-Fl9�ۓ艡cF�RD;s�/�Y�ss��Y�l��0سŉ���T�̆�޼wڲ}��ɻM�U����ݗ�t�-�:��W\'oa�
�rv
ݫh��Zk#qU��	Qܫ����n�+�Gj�>�:%��݇n�\�IJó~�7Xl.�6�u�{��i��wrn�h��V<C���a�jݾ٪���s�h;�mn����t�%D�NGo7	�P��U��r�s;�ۙ(Tմ�W=�9�� QܤE�U�X��ajK���V�ƥ��8nq&�H�{��g~Ωx�u�9V�z�]�q���^��M�ոiv�e�Ss���:/�jq,V����v�l3a����)�o5:��na�v�Ά"f��N@�M侲ݓ��L�nhm��0�՛wD�t�� ��g+���)[!���k\�i7&��:�yj�z�ˤ�ԣo+p�I�1�F��j�nHQo0�]V`�(�d�Z�v��
>�r��u2���V,�uE엺�wU,�,i�8���W���$=�g6�'JN�zꪷq����B�#Xx�u�S�uIݘ�TN�jp(�`��k>d��8f�ȨoZ&�odVC{�;��R-*��UC��oDŝU�0��rn�j]n��b2
)g\c(���6��H��M��8pp�z��%"]��|=���x� ��{�m�/��C�s����8K���m�m;��2:���ʭ
��7]��qԊ�<�o#��,t���m,]
TK����)O_Wfɥ�M�������:bp�LY����it(�̴��FRk���?�;�[��C:�t��-��	"�D�έ`v��q�4f��	1N���m+%�5��F�q��U��6�㾌_n�^�N�U�3�x�Օ�����w9��ZK�*���wS���{*Pm嘴��v15G-ќyp�nSw.��:����P��v9�u�����L�On��2�����Ud��ol5�u����c7tl��
�μ�6,S���ݜB���4ic�z�����Rń�U�*���Y.�O�J�꾾�(���/n�:xMNV�D5e��G6��R��6y��F[ӍʦFb[�&�Y3
"e<WI�FH.�L̏ivu/)�:�5p�U�� �����iˣ�c�-Z:�=����[5�mp���DN� 	�\��7��2r8�m�����;�y�� �wr��K;�ok�Y-�w@��Τ�*yfm�#�2�uv�N���T������ĵ�c�݁��Ӥމ�8�S;yь��lk�rm��Vьu�/Q��U9��Q�:�_e��J"�oVWu`�`'a@ڍ�%��Ð����b��+�d��_�n`��U4���xT=Ó�,e��:��W�]:�t߁ �%�H����f,yovb.�!����|���0D�ge��>�w�oJ����	pdՂʒ��(��7q�AiR���YG4q3�k�6\e��	mjR�M���S�`P��^Ԡ���>��.Ü��W��*�۶[}��&�Z�B#���ڕ(/*K&cr#�v}i�P��=�]v�~ۖR�Vu�7L��M9�Y����Y�*��.n�5�VC����[,�9�O9Ta*�O�:4�Yo���L��1M���}Fd��=:��w+X��{]&LMP�x�A�-��(�2荫��1wb�h�8%�\�8l��g�ԕ�8��:��W��LMR%m�0�:/�
�]ٰnW;՜[��Y�em���f�!�N��eNE��0�.�p�3�G2��s�^�{���xmeW��6՜�ȗѱ��}����_]ka��\�����ݍ�7s*f�iw	Q�Y�&�I��]���g�l�;�͞��=�tb��p��r	��iI�#2e;��R��#"��V��Q�ϫ��7݈eu�Ox̖��2Uc�{�ޗ��b:�jooN��鹹CM����z�]tɑY���:ݘ�M�Fܙ�(��R����/��9$�I$�I$�I$�I$�I$�I$�Hb�H�J9#�Ę��;B�1M%7;a3��/�3V��xďC��Y*�o]>��&�����-k1��<1�ݠ��Pe�5���"$ˮtB{��1�j:;��n��KҏV�oh�{Ʒ����ֺ⣻�A(GS����˰���	wٓ~�����Xv�5�R�vk�d3J�麤�H��=s{y�����Ggo�������D�!$��������y�w�BIO�;��>�:?Hvd�����?o�d%?���M~Կ���ov*�	�;���[�:q%��zO�MB$�
u��n�5�G�#�����n�oe�n��Ap�lCZ3�o�M팬5����������h0Y���nlѩ9�2�C@}R�,ݳ*�i;h�2� k��txj�k��D��^]�(����⶷^�i`.�B���F2D5e޻:�s���!�˯��AA��K����Ni�{�D��R���(����HYa��w#�֪z�N���a�9�pE�f�è������)�KmˍJ�FMs�*�u����9&l���ޔk(V\�kk��:��];���D��k��I'N�w��D���T!j��yX��ɴﬨbȬf*�`�U��?v�8�uIT&���s>���f&M�<{�BP��P#�Jř1*���U�؊$�N��eLj����z־�.MiȄ����<ԅe#h�kv�'qWN��r�n����X���R��A���.j�p4T��T�#�t�C�yQ.��{}��=rޕ�їA��N�0�;����4Ӈ�B�i��Av�CJ�u����8y�d��e�]����V	��5�nݬͳ�W*腠vț�W�e�n�9���9����|�������ʌV�8�g(eb��݌ۓW`�/ev�7�O\�A�s
'��#�U�����$��^��V,�d_�y��JVY�x��%�r��D����u7����䮙���mea�Oj�D��F�W���_*�e&��ɲu�QV��RƂwnᏥ�kw���
�oJ�Sr�%�K�i�K�0��!|��`1��o>���նA�bzU	S%�5����Yv����]�<�xYݥ�a�[XGp���p��s�n�aϥ�����U�7�B��;���MU��5�*�4�����̘F��1�.�S���o8`��]VX�	����r#��r��4��w	�8tZ�8�ᛧ��p�`(�]%Y����l�l�B$3��9�0�<�4���{��&K5��mځ�OUBIQ�A6����2�rp4k*��f<�vr���9�EV�&��n�F�_uQwM�c*d�7Է���M�Y��hR�-f��[I��z���פ�b�&�\uS�y�#F�Uvg\�ݡ9��.���&�ȥ�&�d�-\V"��_
����.�q���s&�����ʬ��6���L62�5V���Į�Ѕ�/7e��˹��zȿ����D��-,P�n�ڡ���Ɠ(��G�e�9�l4���]��օ��ƍ6�b^�z�����j�1qTw���O��tv��Aؤ]#q�.(M�j5��B�˶~�v�\�7@)o�V($w�Z�>�⻢���̲�6��24���n�F��s�,*z�+%]���_q^�rjy}���f(-��4��L׆�L�n�Z)V�e\�1��7f���x�(�������Ѣ�MvC�J�{����ە �r3rp�D3q��j�|��nF,W��2H�rij�c�"�-�.�L�S�:� �Q
�"��r4&�N��u��I�oh�M:�R�8Ͷw5����	����.�Mc��{�����Fa^�68�Rm�=\��f����
����R����V�7!V�TЮ�N�ݷ*�b����`A��%����'W�-P�5�λ�"�N-���ioe^9f����N�=��`!6$X�Λg�2�l���S��P���6�_+3�5�R�&�W�n��r�|Upξmn���s�r�d�-�GK�h<�n�m�6�hGf,��Y%�i��9cA5I|�ү�k���EWQ����OϬsdgayV[P0a�6�:*����|���M�$�n���Tx���GM�!}j�m�Gw�e%�-r՛��A:������i23v�]9��d�Xd��F�uU]�t]VT�^(\���T�цM�]ZV��lR�
�A�}f�n���fT��@woN}x��5�fR��)����7n�)�AW��.۾�1��
������	,ͫ�����H�F�5�Oy5��;rnsA�Ԣe_V�`�C�	�S�LV*�U����GR�tԏ���rУD�_<ڨ�3[OQ�Uw\��-��M�Е��l��w+�ue��̷����˓�-�P�8�c'P���BRLw��Ǖ{a�|�XW�wlT�Q�	�+�����0��ͭ
#�|"ϻm����6;�2�ƭ�d+�5�x��'�sq��W��LoN�)��('ҙ�QDX�X���Ѹe_8+��`�8�LMWc'1����3o���b#��lR���Sv�q��ֹ-��a�x��:��k�Y�Vk�f6΄b�U
��V�����b���61u�=}
�(+�|�H{DS�]]s{+�=���n=�MK�gai��V8�$"�T���y�b�E}�o������MG:�/z�i�z#f�)t�D�0-$.��2ѡpU��eK��><�[�
�[�� ضi�׀��*��;	e�M-X/{l�/��eʹJ������������}:82g܏*��gR�,�R���_)YNC�$��(>��wW5c0O�X{!;H��ɳ�C��};��Wectsm�H^>r���txO�	ϕ�>�-,ʋsI�`aQ&������N�mEֶ4q�����V2�v��p�=!2c˷�Q|ژ2����ڷeX��A�4���[����LZ73v���9KZ��M���8#��n�K�����`<�)�5G�x,޾{Yt.ڭѢ��SB��N�Gἃ���@ܘ��X��'���0D�zz�U��wX�F��j��v��WY`ԭcN�j־:-�Sz�Umm�4�����-�/FK�,�Jμ��N�����6�v���^RnޛzV�Z�a�N�E��%n���l#�7\�k{��_6���.0oL�J����!�+J�J�3���@9�RBX�O���C�Wun7�wY2v�@]w.d)��wIF�AӲe,V!A�s�f��^�q�ce�콹d������#� ��W-!�.�6V���p��v�%�v�-dfT��4k��:����z���(�k7�JR,���	Ws���Y�,�/�)/奥��х����J=s�5{�ݠ{u�gD�335s-���uc�����z�g:l]4��`��kX��u8��֧�J@����/��/�<ܾf�DS%��!����6/8R89,���R���A�J�O�3/�}� @�"
ȿ���:�'�XG���S�d������Y����TDa����b%��������n�K��m�U&��{�c�U��)�n"*i�Hw���CG2�`����˚z�m�0���;��fNWY��Y/���E>�E;Nf�|��wV�7ݑ����9�UIX�:�Y�2�f*�USb
.��f���[۴�:6�SJ�`�-6�-p5���)�y�v�U5�|��>�O[��W�Ji��QLm^։����I�T�4�
�r�L6;�I:����7m)yP�ҳ�&���_mY�j��z�x�|t�� ���k�%1��Sue�J]��X�\�M2��7Y�+vj=����/��~�$� *%TRT#����1��@�%Me3ŕ��;�4�ՙl�j�*���W()�+k*�)�1���cr��B�MI��-��P*�Ui��Ęͷ-e-Ն���l�Ţ���\�i�+�f� ,�J��²�3�Ҭ���L*E�J�UB�
�X
d�1�)Z�Q]R\[�S)Y#l�U�q�l�
�SAq��[�s������͗�zE$5��hgjW4�
�샖:_9��ʠy���k�k𡢜��2X#��k��Z�G�a\���`��]���o��mr��=ڍ�s�[���0�;�'���7�gk�^�{�3�hékL%;�s\�qb�D'��A5� 4��i����n����6��g���#Ƽfq��|B�=���Q�fc�Ci�L�nc�^M���L���Em��u`�⸎\K�1���j���.��-��Ա�[ˮh��G�b�C|0�����Y��,ݫ�0��/%r7[:��B�|ܜ2N��\
2�Ìk=9��>~�,1�g�!�ͻ�N^]�Ux*�����u�[��ײ:��O������#x�R��y��ip���'Qn��#/�e�r�v�f�aYv����oF�O	֭F�{���H�����dS�h"ܭ.�Ӕ�`�d?3��o\%���ݾ�(����R �0���	Z4��E]u4��ڗxZ�7�c��ᰂ�z2@��m
ž;[۾"Ij��js�cv9�^gs���㓒�f�� %Lݧ��!d��c��%�3��S�I����u�>���ghCX4y������`]qEv���jޘ�����M���̥@w������ދ��绅1
s�v�Qsy�U�^.w.5�mQ���-!y���K���I��U�!�ZZ���=c�%�f����=��9B�ZWp�
������\��z)��{��V�� ЖO�h��SE�²�]�g��Pa�f�'�n�ʮ��꒲�B9`��0��LVr�H��x:��~��פ�4�JEz{���#5���s�b]���8���8U�v2�m�>7�P:�{��G���b٘�7V7�d�1����W�i1���W�x��S��[�-�ꕼ��uD1�Ӟ��ԁ��r���D�/+z�N�����*o�#30K�Ө�w���s�2߻�U|�$T��7e����Pge0���U�.�y,����-���ӏ2*{ƷY��񶄽ux��;"��R2]X�kr
b]���<7Y���}k���;�h�����3s�{tkp-k}�w;/|�㷤�n%�Q��,��[��!�5
���<T���1x]b�M��dq�-5>Xq�M�����3��[�Y�ra�����۳c��Q�-:�'һ�`�,��Y��(��_s��!f���H��?i���/�?6�v��錜�^m�Ž�nݫ�}g�p���Nȇ��ş��ת��gڃ6@���T�CHC�(|���Y=L՗�G&×>�JI������4�!Ix����q�����0���*���6��}q���9|��׫�]P�g�b#�|��?`#Jm���U�M�4-�g1��ls9ɬ����,���u�1s���b�@ۧY%쑺K4�dR*-�ac�Ue�&���N4���I�O�'�c��B;P&�C.�zf��x������O̱�<X_��k���%gid��ʱ�X����)����_&�*���҂�	ha{V��/�t��œ�k�S�m�#�B!���X�G�	�i�Μ4CL����f���LQg��}v��zl�X��4e�����?���ve/�h�E�����C�TDnvN�4D�8���(r�*y��<a�����e�{��C"���Δ���H�������i�}YW�;�0�=��� h�[�X)!��n:1���pS�J/R��s�RSbiߝ�t�-�cZfZ��,sӶ�k�r˺� ��Q�R,����w
� Zƭ���W*.>i~_U�ӆ��"� �Z�~�j��8��y��}9a��Hm
��U�f�#�³�����ڿ^S_t_dZ_�B�G�1���2��s����_r�����|�A����!ŏ/�I�=*�rz���|�!�r��a�ӗa���l�>#��<w�~�H��d>���:�r������B��l�/��#
�W*?>�o���]Q��L ig�a[ɘ5��s���i���o��G��	��<C�x?j��,�MĞ��U�H�T�m*9�� c^/ʎr����z+#���W~ř��/����ӧ̩�65�iV	���9& ]��|�j�.	zJ`��8��\R�)e��.Xs{��}���B�mz��Tѓ���y�	�ox�فT*ɸ��05Q��Ge�C����:��U���gy�b���B�޴4��t�#"㼉���=�����9�4붡��0��Ȑj'+�Ue9tv�����2Ǭ;�>#M#&����G1���۽���4�/���B��aE�.ЯCw���^�<G��򴾞_#��OOQ�<r�[����>0�(����(;���s�����<F���찼Ɵ�4E������t�}���!-�{7]�1g@ ��n,�q�e���^
�ۚމԜHk|�ީו���gTZ�u S��N]�ȸ��T�^��i�t���F��N��7khgؾO��y�C� ��<{��{�a�w}ݤ�Y���/�><\agy���5v�o\�ې��)�!&4+�2 ��uYQ�0ކ	�h,`	�L,�dQ�Đ=Z�=��}M^��n����׈wy�1�B(�i �Y���έ���}��z!�S���YF0ٲ4��ߑn�����>��<j4���7�=��"�
?_����G7�z8�8$���=�cE�.��ſ��YRoWN�q�l$��A���r��e'�FM��B����B�����O�T�Tg®�E������$�H��NI΋*�GJ��r9A�c C�5�����oL�ٗ�J�j��:������x��C��y�^���vrk�da�~��kPu��Y��s�*����@�Vg���� ��R<��Z�G��T<<�A�IY����8)}�q�]���"7���ͬ":`=��[c�Y��#L�Z�=��@���-$���\�."ځ>k��t𱼰��/�T~�A/��,/��~8<�է~G��a=~�>#
�!ya�J@9--�_��8q��4�8B*���yi�1�}ޮ���k����#�š�J> alii�~� z*����Gr�ai�T�v&=��{���u���ޟ6<�w��ϣ�Ð�oƫT��h�iM�d��ҮK�w	�s��7���9�(UA��ڭ�$�)�j�=�5�^|�d#D��wM��+R��u=�72=��3ْK] 9oQI2�K=x`z�l�^�`��t]��sz;�qQ�Ť�Vܱr+�kbw>��ǌ>�YDk�p�O&P�Ono��d��2�.e���N�\۸�omicA�[ǝ��ڍ���ڽ�X�r��Q^�����naY��1-�x��l?:٣	���J�W>8t.W����y9��է���tk=t.�6|as�ۨ������ow����e%]6Q)�v��̲�CYs��t��Q�,�5�0Z�n�\�r�V��7d�3���W�;X?/�/Ƽ��k�~I~]�f��5�̮9G�a�0�%r��̨��X�3�>c0���孽��7��T-� q�.�n�(�<��[G���N^`@1Bm;wr���L�hFk^�J��wa�<��H��,�'�ow��3�"1_pN��;�<冽r��n���I�-�1wR�|�kmet���f�
�n+7�tk����n��m��۬�Sz�����'u�30� ��to��'�d@�f0b��sc�׿mnы���%��������T{�N�����U�֑�N7z娹��Z���E��A�����K��re�E�$�ɰw�_;{��8�\o~���{�7�*
Tk �j0�LJ �1%A��bʀ�*M7+��GPX[JZ]P̠�T��-�іȲ�m�G-TCX*Ņ�b���d�YRT��kE�6�
�A�p1m�,S2�F�"ʭ`��E��J�Z�Lˌ���L�LXԨ��V�Q��Q����Ԭ��,��WMp��b5
�q�p��)E��Ř�\�Eb��.�Țb�k*"T�+%���ȱb�9�������`(U���6�V]�D���U��I��̒�T��8)I�Xi�x�R_��}�C���>����
_2���/�;�I��ʺ�<<��Ӈl鳻�g�a�z���rr^7��:�.OԝGe{'�違�^sUm�h���	��ȣ����F��Ժ�Q6Hx֑w�#��o�8O����O�ˈ��3�����q����T����.!ŤbCk�`x��_�����0�����x�t?��C��NX��k��[��LGO��-׼�z�t�J�5
sF.��V�߼Я�Y@B!�y]���u��]���a�y���Y�i�͜Yf�I�������:�Oo�3��z�@��7���T�{�mc���h9R�� ]v�ՌN��JN.ݍ�|lۣɷ��%��T�l�-�o��;���M����4l���a���B����8~&͐�?��(5�r���j���i񸰒7��_5�$��@�lbF��y{��L�#�6��?���~Ts�{y��3km�����.?YP�b_W������?:��ۗ��(�!�T~f�8��!��J�V��̒����K�<x�t������ڠ��J�Z� �},!����_x���ׂ����0i��l������t�!����9W��^�`�<x�I}��gM�"���D��\�7O$&W�6�R��o8��K�(�S<룥�[��YR4����v�ˎ�/�6T�%C�'���ܝ�9]���3+���]1��A�q��~"ˎ��=�ۭ�҈��Äq�~���E��bj���]��q���ӝ��x���f�1x��+{��u�0��64��Hg���P�������o�݇>vǂTX����/�
ra�B�Jb��n�a��V>�\���L!���9������_-�3޷Yw���~6���!	#9i���? =��[�Ƣ׾��Ɵ}�� a�1
6 �w󾺫(ȜV_��r��Q����h�D��V��N��ć{��S���hitÇ�=�w{�ˣ���aW�j�F�5a0v�]սه8���@�X�:�>��<�m󑪄w5�n���^'w�;��#z/��+`�=
x��!m:>:E��u�n��&;���w9���G�m�:>�=�"!���I��O���l:��;_[�J�1j��+��T��B��!����ϣ��80��ܬ��C"��@�|BHC^�W���GZp�)
 l���=#�C"�S�Rm���ۛ�ϐ'j��In-,r���Az���5Ӳ�����	�:��H
�Byo��\~��z���"r� ?x�$������2:������9�0�x�g�����|ψX���廨s�C���5L��Hn�/�iV@���e�
�gM�������e���C=�"�x_�e�o����Z�C�a;}��)#+���ڳHI=/�}���C��<GՄ&��A}��}�{fv��9*�8�t�#�m�p��x���ׂ��ٕGǈg$v�<�!�<��_y�ɞ~7C�2��e�>?q�E�������4�1Q�~C�����yZ48j���!c�|��;DО}Y�Q�8�\E���4�� ���$���3���^m^��D�����E����� H���	��u��b���!ڞ,,���2�@�8h٢2���N�8��RDS���Α���l�?���~x3��~�.�h_<���f�^��XzA�J@�ؕ��S�{�����1s/���wf�#[v_;a��6醚g�Z=�ɓ�*�����0����ԾgM��W'c�K=�Vw�����t�������=3�W��w3�Ixr��4�����yZC½�.���l�3�����h9iw�m}GH{�{|�#���g�H�`�l�K�Ѳ0�j,f^�\����Z~a*:Cz�E�G~�!B�*���3�����3D�ޫs3+��\D��@ܶ5��޺��#��.t�ٛn�yQ.e�<�3���@{����YF��F�����ˇ{VOZ6x���Z���* Y�8��׮��X�7C%<�s*���vQ�S���1��$a~��X���ܕ~ ��v�wLN=L�ڜ>��;���>�`�����`���W_̊�/�
v��?S9u�;7y~�oA�#��ń8��;�_W��ךj���m�8G� �>6ns���"����8G�����Օ�E�~��I�i|�fN�!�A�J�{	}�m��dj@Q
��p7���q�d��|·~�S)g�	yr�_���h��=��}y�7��vk���ܾ�_7H��3��|s��p�����Q���
-@�ٷ학�4�1��Ǘ�����4�hKLv�K@<Y�t�{�b��Eؖ��/�״��P���v������j�J�aF��E�t�5���*�SO����~�ܜo��ӝ}�L�drӈ.�Pݮ���{C� �*������k��K��Ar��?Ǧ�yIk췞���ā�B�������?cBϏ~��xgV�����{�az��Bkc���G�!}�K�{s�,(�o�:Y����,�![�aZ@� ����Z�w/�Hm��^X���>0+%�We�r�3y�o�j�5;��۪|DH��g��Q��᫨7��K���0��������:��,���E
���]�L}�+�|G��⬊�O����J�uX?Yǯ��0���A���r��=�q�G�\i���1HQ`�����,�A �֩x|�%q\�<�1���ƨ<傶��;Z2�w�jӆ�+J�qG��7Ƌ��ɭ��[�1����/g����#=���G�J��|��H����� �-ns�QOV�tO (��ǒ:��t��!q[<���A읛s<~x�ZD?q$����Ǐg�v;�0N�C���?���0r�"��3��B����xy�����?C�Ī�u_U�?���4,��/P�4�Մ"�k�;��_x�<��,�k��8���� 0�4���w�
�4D��5Q[�cb`�sn����Z�sD�3�a`��Ee�>4~��|�~YG��T̹vP�����a��*!dH.BƬ!��ɹ�2����+D�h�|�{���Hagju	u�2��a�y��#��D���:���94��CI-�,�5W~| ��{t���j�?�������x���><���x+q���?q�8�7��ő�"!;E�(��U�~��	#O�vg����o.=��[�)�ˆ�'O[��֟��G��ʚ	��Ǘ����-�[�\6f�ۿmmw���(�8�����/�E����^s��^zƟ0�WN���9s���:�G�7Vx�?O!��>"���¹]60�hc�v����1�OAL�"@x�wg��:�n=��5�	DU�����h�p��E�(dŧT˷�(��6w�G:i�0��B��d���f�~C�zp�Z+F�M+��x�����lgM1��WSg_`�mJ�؈,����.�4�.|�zƥ�w[��,�[	[�2o��H^ν5ل�<���"��W�8k�U���l����;P��vK��#�:0���t���}�Bqm�B,Ť��4�c%]�*t��lG� ���!"me�u�t7�P�7��� wϸ�NwO��ӫhʺw�q1,�5[�a͌�
�zmc%�2Vܪ�J2��5R�t�n4Tpt�YJA�B���#�J[8���ɼ�n�&��kSx���1{ظR�L)�q7a�m��:t���Vz�f�!YۀHR;�Wr��%:��eS�;Oe��	N�nEy�]Q��B��+����A��\��F�c�J�8�U�:�:/O����d�[M���ܵ�9�Y��F�,K}SQ�����x`�]pRN�L�^9\x2�R�A�u�n�4�γ�>��x�3s�)��E������v(��7�t��k]�-}xy���(�
��7wq�RQ�]53��x�"k�����v���%NހA3��,RZ�GHM<���gM��lWn�E��3X4��:�}d`g�;�ޣWꛒ`3����$a�N�H-�[�AR}�&���������R��	�\)k�}1�,Ʃp�S`Ì�t �66POxvܳ��kpL�H�䋔�e���ɮ������{�|~�������T+�I�mN�`i��i�+*ê�,�I�Z�F���l*V�)hU2����T5h������`������H�����E���5d�]Y�&�d�$Dl�
��V��X���R[HUj"2�3Y�)
 �i:IE��µ���bJ���`�*E��Q�$�(�"�UACM�-�%b(�����z{���/:�uz��̍1�e����'�jg�ff-?������/ʉ���ԧ*���SS�_����z��,�����2(���ӕB~U�t\Ţ�ݣS�teuD'^ѫ��D��b_S��fQ��ݾ�~�ƌ?_��0ٲ��(�!�g�(�y��כ맳o�¢�P�\a4�Y;e��1�Hp�AH)�
������Y;=���!��W�H)��|㬽��2�y�|���R'�ˌa�B��옐Rk�����:aR���bOoL4�P�9�Isۈp��߾�+ךߝ��2�^�
Ö��q�����T�ő`t��sHV�gᴂ�]�x����2VN�Rs�H=�*=�5�v�s�8߻�¤�C
!Qa�
Ɍ��[�(�*h@��
°�
/���)!�� �HVo�m���������Z�7���8`r��T��寇v$(h���6�H(v��(���&$3�L�zɌ9M��$���PS�9�8��ǝy�� ��M ]�=�a�
����Ă��0�R
M�C<e@�_)
åB�`T���1E&N�c����>���k��f[ClW�$Km�K�q���1�>5�*��%����赊�6ҩ%3�)Q�6������
z�pj9�=�{��I���c�5^�b|{g,4�P�4��YE$���φK�=@�0�;��H(���������B�������]��SIԨ%@Q}�8eC�� �&e��VmI� ��E��+�l1 �m��(�L8.a�Y�y�<u������*A@�5���!^P�uH,������*)�μ�$���OL;aP��
3Yb����&�y��u�<IR
w�8��La�
�R
A@S�ӄ
�Y�J� ^l1�0�
���bAH/F��4�AgL���T�����CyHV+=q �a�EN�1�,+&�RXp�r¤8IR,�P�J�YR:dߚ�D+Vy����~k�9�Rz�@UP:J�X�������Y�i ��Ҡ(�N�SH �d�Xr²k�1'�T��u��=���� �Æ<@�����h�Vf�)�������@Q|N�1 ���u@��a�� �C�
�AI�:����s�y瞥{H,-}�t�Æ1�;��Y9�Y�z��4o0�՞2bzΘbAa�
�P:�0S�
�u����g��y�ݻ�޽��:a�
�PĂ�D�,���v2vʆ�#�!Xt��`i �5�Ğ!PSh�,+XT���\ٶ��9�ݾY}�]��<�T��TP�%H)�0�&n��6º`y����PT�!R�ԃ�!^�t�Si�I�G�>������b�H�p����ާ��K�\��d���j�֩߁s�(	,��۞!jfS΢ީ	�<L�pp�O�u�7�]� �ߜ��M$OS�
A�0�,8aX|0�;B��Ö ���
Î&�H/l��$��Ł��.�����[�޹�Nr�x���a�偿.$-x`T��L<q ��;La�
�R
$��L*$��2�H<��&HM����<޹�<��gt��6 h��t��r�Շi*,�j���nu�s<I�!m ��NP*A�/�0�@�T�<IR�C���"�Y�6�uHVg��� ��`*��n���w�1 �:jA��ی+:LH)ٔ@�*�&��
C��+0��
��+XT���y�R
A�}���z�}�̢�Xi�H/�=C
�0*As��R41&0�<�N(bA`k�� ���8�P�Kh&0�/=sםo�|�;�H)C���J�X�(x���͜�cXT�����2T���PĂ��p�T�a�+��H(f�ߜ{����{��=0+'l����ˤ�i
�3�C�a�;B�i� ��H)ى�a�
�`��J���$4��/7��w�w���:�gt�a��(i!�5�Ă�Uû
uaۤ��Msf�v��jA@�*AH,�2�K���߾ﮯs�,��0�AI���dĂ�^�bA@�*A�t��bAzN�,�H)2{C��RZA�B��F�D}��A�"�������C��}7集�*=�:��Wי�{[�h�ĉ�m����R
��i���m��f 5�y�� �|'� (�2s�����n��c�
�P1*	*���ACĕ��T�՞3���p z� �]i�h�k~�Ʒ�IQL@� ���B��y`T��@�l�*J�Y<��H;�(åB��tI�����������Ӽ�7�:�Ă�}�!�a��wd�<IR
�IR
Af�/4�C���$=���$ժAH)�'�$�u�r��߶��|�vE�,��O=�
)���(�凬Ă�gV咱a�
�Rr�H(
,�8a�&{C4Y4wtæ �k~o8��u��p9H(z�E��i�!Ͱ;�搬4�̧( ��@Qdᕁ�RZA���0� ��J������������ACi+��l�|�a�
�|PĂ��PS�
���Ă�%H�HV'٧�`i�񒢘�R��<�^y�>�VbA�!Xp�T�y�AI��9��PqN���Ƿ�,�B4�M�!�����IU�h?/������랪C���\�0,@����a�e����� ��g<��B�G��2/�S����s��s�v�\g��!�i>Z �\nm�ti��i���j�;�T+xU�lwD��לW����������u�����,���o��o�ߔ�z��i9o��p�g�����W
>Ç�L�/�+@x�w��V�7^��o�+ �Frt��/�Vɣ�y}�)��R����G�µG�p�������!��U���E�g���c@�l�$���5�'��{��!W�ν�=�q{�8�'@M:q({��얲rf��u���0�/���x��^�D0��������O�Ҩ�b��}Ϙ�ū,�C,����%8��߮��d�8�W���iҴ��C�޶�E%`�W׫fҧ���:�m��H���x1�q���qֹ�[�D�,��$x���+��j�˃7p�,[,+��6��#.� � ���W��4i��di�f����|�;D�
�?��z�]n]jN�&Dx���F(�ܞ^�K�[�<�#M�/}4��E��X�K�Ot�y�;S����9|jw�r_/i���ݜ�B�O۶�����Ś��,�
hi�W9]p��$��h��j��WT�eI�C���@E��1)����D!��^1�%G����{���;+ˠ=�33v��Z�P��mq��9<�z�/J#;��n��uxĹ�md�H���QMZC+1߯<�{���#�R��z�Q~���.�}%w����p.�/B�yA��
�2��#������8j%�f-�z�8Ҋ2fwhQ4n��{x��G�ҳ�5T�g�?mE��c����^�&'�Y���;v����F�-aDv���Ȇr�!x���)�q����3W��?x���.&8��B+/�=�>��=u�>��G�x��	ה�H�b:;eͣ�©S��������`�C�k���'ud��x2<ӵ܅�?A�V����G���}
ӳ�zH�d2;P��yi����F����]��H��l�D8B���HQia��H��K�-�h�K���&"F�?v�vmOtɽ^��G���HZGˈQ܁�_�13/C�\�)o.#�V؃�jE�՞���&v��ܛ�����M㕩�ַ.�q��饢�GnB)���G��uI����~�X@��~�<(՘P�S�6�U�TC�	�qӧ�K����R׼�j�����N��1�v�CO(�7J�Q�>2���];��Sc�(��
PQ�xº�ˇ�S�i�qx���0�t�#�m�p��U�\�z�����O��"��yF�ͩ��k�����p2�LE�W��ND�.�&�S-%�4�9��¨wq��"�Q��"�W;�����6Gb��V~��U�־��D��;g����L�^�H��P��L"��O�Y�	r�]6��<��&�su4o/o;�ƦQ��Y0�4�3�
ﭦ�	�&��:�pb:��`��y��0�!o����r�*r�噺r��/&�N~/���˔�{2�h��G�"��H�_�t�t��}�}�^~�*��W�0E�h�~�L:l�>`xx٩�s�>�s
�%�_��<�����E��N��{佻N��e������5�Ny�,]���1�o64�@*1��]2t���K:w�^g�fo�h�� �GyyϜ��*62�L�um���}R��lѡ�����k�/�<T_j�'�+�4x�L�P@�d"͗��bCm}>k�Jr���q��7���:Y��-�(��U���_��2�X 9/�/��$��l�q�0D\�V�_!#z�0I�d��L5�Qb�/�p�o�w!c���;�}y�j�N�c�\ݽyv3��ίe�F��
#:��/z�;�~vT8p�W���9Y0:�dO�r\1h�ry�s���+�Q����?GƸ|��z���>��W]Q�#��[�<D~?,"��C�b���e�W�0��r�
A����xx:�ѱ�Oz��"�:����#�24����1/��Jd�g�*��p#DipZ�zo�5 ��,�+/�e�yK�����0o�B�����m�ʑ�b|�\@Z�6s�r\UD��l9��
#N_�������$���D=�li���5�����������[�/pJ�8~�~;�ז]ΐP���>ʋ=�i=�>�?4iS[n�yҌGm��eg0�G>��&nQ�4��*߃�K.R������YF�5}�ڷA�&vA��K���ym�̜�S�P�3\(L���2��lH↻�GV��W�f��He�|j�n��χdΠ�`�����3���"N�F���	�T�9��$\�8�w�U}!�����ʢz�pUc#�_U���'9����YK�y��)���M�] nK��k��}$�g}�L&�D����6��b�"ԯ��w��ۡ���� ������k'zul;c�w����W��ѷ�gB-ۧ&�Т�����O2r��Lv�CI+�$�x����䣽ީ��r[ǪL�J��R���fdjwE"��&n�n,*��!>��^"��]<6�B����j�j�w1j���48��sng>/�Ŋ��Fa��%%Y��X���"���d��I���N��Y|8({;����X���I�����Fj�q��W���oR�R)R�8�KqV6�"D�e3��c1 �u���(�Mԡ?���-��N��זCN͝gN0b���,��S���c4���p�A��`�i|i;�6qe�]�uf]�0=lMp��Ň��rgt�SYB�6�@�S ����a�&^$\rB�NW�;���StkR�w~�����V�����H(RЩiH*����0X��TEQb�B(�N��i�$����1�@U�,P�D�D`i��L**ŀ�b��"�b(0�aRX�@X����id�Y�bEPYQ���Q`�� ,XXdR,�,�Ȫ)�(�Pc���k:� 	�O�,6�r~��H�2�,���ltb� g�=�z ��'�cg�>�B(������/s��y7��ְx�f���^��(�t�L�̸���]θ�{���vug�����w����i�r�μ��b�����qZh�>�� #H~�pBw���Q�	?C�\����5�<�b�E�=�����~�����"�_Ζ�Fr�c�7���7y��Tj+8��~���8��/���p���&oK,j�0�?Ye� �4���O���fX�
zY�,�"�2c�O����i�=��iWoc�m��r�NyNC$σW�ՙ^���i_�MaVjձ�����H�3b;2b�ݷ��{���*�Wt��'O.�s�j�&�-H�e8��#A�&��W�}_U,3��K����8�V��s�OZ�o�Ȭ�:���gH��yL<�>=��O#:����M;�J����G�C#���/��"Ft���Vg�������@�'ަ-#�HQ�=|<���Z���BϏ�F���_��$���������(﵍<ED<��Uha�i��EFWx#�m]z��+ ��z�P��7V�j��K���
�"�_a^_'�1HX1����^�B�w��p�W/���H�S��/�x�C9���/K���4ΐ:���Μ�d(���C�b���U�+{B��}n���X�ˈ��&FGlٺ��N��VNk�;)f��Db�e��N@��i�/��B.t�U�W��]�;G�����zQ�ZX?E��/�ݞ����x�;�M�Q�Qu�YT`�:D"�HQ�\ە�6(o��r�|�l�^�#Ծ����M_�GY����<���C�<0���s�!�Y�.9��o��v&'�_�r�Y�ö�yx5z{?W�yt�^�gǎ ���)���kdk�2Y:.d��&�9�X�aC?x��.��O+%?������
�
��@��N���5U;���P�V\�<�.�Ƕk�s�z����zwa��O$,� �j��D鿼����_r�u]x�A�z|��3V�
��W�H]ӹ��#�ʶ��hb�e]�ۓ,�J����ڹE�.iܞ�=�X��[��Dz#ހq6����|i�\U\��A���T��2s�b��|tW����#�x���?��{6i����W^Y?{P�,����`�g�i���_�yَ�J#��2St���hi ��O7�]�4��?� ���x� W�&&:b��U�.H��˅1���Y��'+��l�ȑ�&}6�'Z�s)�U
D�[�Sηr���_��yՕ�>�8Y@����-�����~N��~�#�.���{��a��`���+7^-�/GUxn����X��NB�ҏ��I�öYF��,{泚�9�3��2��r/�S���	�'�n�z#��wnp��rKN��ՕY� ��Ze�SW����g������1�_0�#�DNׇ�Ԁ4���f����5}lpz��.��x�;q���8�;³=�4y}A�C����e�<��A����zuvQ�x��5)�8~�%�)><~k�L��R�݈xr��#�"�^΂����o>��XL��L�])���=��ΛI��f�G�;�q}�K�	����+/�+"��<�������H�\a�sPF�,׷�E����_�8qp�'�0�5`��i~_v! ��
엾��]�5��=H C�f4y�Gő�^��M����x�޽��V�V�����g�����:�#w|��E�y����n4<6�oB��׭0Zޠ���x��W�UUA��i�e�/n�׆v��^q�o�箹|�N|�7����l����!�-/����{��y{!��ۂ}k������Y@��٫��z����b�`��yK�~������T>�g�A���̀(��7Z~�8��Nr�׌(��W���Ӯ��D,���]�Ǖ���"�|�S��Jަ��D ��@�?s�"F�{ݳ1+<<���#V�,�ȅ$y*b���mG�yU{E{E��
���~���O����B��bT�лG]t��Hʃ丈Gj�`����~"z��~�nz̃O2�W��䥺�e?W{�3�LK>�4 D��.�p`֕�k��R	:��rS�/_9�N��U��_Z3�n࿨��?���ps����C�f�����~��/�	�?B(�~����!h_���~����}�Li�/�?���<DJb�Mx��<tlw�m��;�W��WU�)�]��k���/�ȒΤ�^��;h��C)4wO�m9��t����7�����m�j�H�@���q��+f#o�,��[txP!��=��)�y���Cs���lL�`�5OCawH|޲ow�[Spk��ǻ���%f[���xO���i�a�*ݩW;�̝w4a�u�X��]Fҫ�nN�9Lf�]ϢC!��UUU�tq����ο3Ks�յ��"��o}�/�Pc�Dr���>Q�<�g���] ��do�]:���=C�x�e�꠫"hT%�!���)h�d,�G�in_K@ltv�)��0�����:��]�uCv��&�f�����=e�R�s�&�p�F�$�A���^~��u����
���q��<n�{UE�޹CM{��j{�0v]�N��q7de��}��^��ڮ�D��9d�<�>�e���ʏ�V*��z��K���/�ZZ,`�W>C�\��ZQ���_Ul$����]f���k��	�g�r��/J�y8вrSŻ��5�wSx�ߌL�'d���e�����	���ǰAE���/c���+����}����ܸ�� knz�����5�e_�幫�L~F,�TݨFn@��D�S����+�~��=�I�*��*O,�ݐ���
>�H��a�<ob4�C[��>�.���M�f/��a-PU����ո�_�_]����{+�=
����R'9�s�Ը�8�.ν��[�n,2��,h\������׈������ޡ{gN��a�cD�=rq�Է5��Pg��������0�׫8N
��j��Ǒ��chլ4�,k�q�4�� R�����[+�-^¤w<y�h��"혝��0Ot����L��3�����=G*ǳ�T^��B�>�k�ә!�K�۝�wW�g~�Kk�5(w3k��	�0��UQ=��8�������=��3W^w4��M1i�3%��5n��CE��'�i�;��Z���ݖ�8�j(`=�*1h�P�����2{����Ή�� )ya��k+���@�Vv��K�yJ��i��X�R�.�B;K�=�YJ�Y��<p��Y'F����9�Kz�+�i�
����Dx*�F52��4\��\ԅc��`tO`��؞�F��Js��k���pW4�r�{i��;p!�x��2��HCv��W7{gI��:�6_wG��Z%)R��7�����ok��a�ppe��`��e;v��kҁ��TH㰶���\׃�ʉ�s{���&q\/��}��Vow){݇�RFv�P}�]:2�|r����n��iи�:ީ����0��`ՅAxt<���镫v�.���� "b���M��Kݛ[�t�,�j��\{�r�\:z�
|�Ea��[��96%�e)X^L̇V(����h�s&��N9��5Ω�f��yCW.�Y��������H�jC�6dt�a���;!-5����7q'n�޸n����J��,�]'Z�q�s��M�k�Syq}��5�uu4^���z��$7E�B�R�����y��n���g�o��o��=$�b�j�˚�v�I�f�
�����hܑCGe[��:�rfiH䙙�:�;��J��s����ͨ#�~!E�Y�
 *� �X�D�E����
 ��*�đE������i��
�fX���1 Q ���,REX��Hc!R*�QE �@XŒbVa]3�()�
²
���(��%�H���f5��}�Z��vj����<]Agzu�E��^i�W�}}�2~�&���ݩ���l�zxQ���m�2:�q��:��(��Tʒ>��+te,Irǥ�����F���gg��[��z��E��U�ϵq��r�=Z'��h�)n�_U�6�o1�LVTY�N��dɩ�Y�[�u<�����C\'�n�	��o�ե�4o��i5�ZF�eM^��Kei��nb� �t��;Ӱhv�y*���钑�|ov@����X42࡬U�7�;���r�W' Q�-�s�\%�64�e�:�Z���3�}U���9_���N�ɯq�}qn����F��m�ǫL�RTgPæOC/��.�<��qn'&�4�+���v{��Y^�Y��Li-%f�R1Z�����LkI��b�Iᶞ�u��Q�w3Ȁs���0y�]B�3R��v�Ī�7�إ[Cn�Mn��ǡ�(���N*������,<ޝ�^����0w�}�"ۧXj��K�;ç��З4���*�1E.�7�xt�Ee������ʋ�]Žv�)NJ�
�	\�Xƿ�}�v�B�G���A����U4*����֑*��7��f���Q�=��muh�E�������z��P�¦�A�%�N�3l�3�˾ט���X����aj�7�q��r�_v�~:}u�7af���&q_ۂ@Ѓ��a�K�bz���Q��Y�ޙϚ��ָR+�Ύ��e����M�mӷ�No�*��OS�3��9���m\�K8�������1&o'�Hpe�߈uz ۭ9��A�s�޴���5[k\�Pن��Z�o��oq���S�w��)	�~���)�6��}H��=����#��l�c�8l�����Cr$l�p��zszZ�㣇f�=jQ.�yy�D����a9���zHU]��Z=�I��m���
������Q�C�����Ü'Z�4���6�%j�*eq�I@�z�-���J:�L��s��f��=���g �(���[ׯ�����L��C��H�v�E{s�ޭ� �"*�/��U��Ls��$��*S+n����j���k2���l�� *X��N��DH�삧�3����a^nt�~��������O�:6�s9�^ B�U�5�l�~ߞG�>N����Ϳ�B��q�}]��%�@n.':pwA�r�����z����z�o�Gv�(�K�W�4iguum���Ϲo7[ڻ���zP�U,�u�xX����P����2�:4�]s&�%r�$�Q�j�>�2�C���-�2j��;{�����×��{å"mK싖� ����v��]�.�b����N�g:�����\����Nݰ�˾cC���e�kw��� ��$;o5"���x�	B�#����%��v�ٜ��ﯙ|q����+��$Ţ�0^پ�(E�=��\��_8#ۥ��z�^�^A+�w����v/P����{	�:]f���⻠[�=h���ǉv�ùa�mc;E����oF�N��[�Z nm$�ł�g���jvD]$�N^�KM�mג �#%�GMI�3Q/h8-�`�}�n:�3y��m�������/�Pc�*�q��|��,_b7�*]̒d���8강�u1|Z}r-�E���Y��=�1�S>�s!�%����R�}�jzW���WO�H]v��j<G�\���NR�]-d�51�����Ew_��{s��бoo��)���b֥x�q�بQ%�5���13� �Q��*`�M���B�M+Q>6�Z�9���a�sg5\���=Gk��5#K��i��$��v��j�Y�B��y3�漪��UZ��'���;���=#�;�-�Sۍ���۰�}�zB��u�ד�p���+�,sH�Ы���բn@�,yR7s�v-��ISES��~���]{Å�{�I5�&4.;�$9*[�p���p�;�A��h�~5�^���a��������e����#�a�̥��NbÜ3��^ں�iк�o&���S2"rI�R�$ؤIp��L�Gz��I���5Z��*g���4c�����;�0�)�-��k�9�\u�TvW��Sb�6��N��Qfk��]z)����m�MF+u̵�4��1Aث+��kd��^H�6ϥ����5|E����y˷Շ�鍣��'s2���:Y.E�1K�=���̾ {����Ha�����#��/�4���]�c>��zm�3��/�q�����h2����}���M�,�7���7��ġ��u62���MO�.�|m���$�O�ŌL��&�O�NҊ�"��W-B�V6=������8#��;�}�pL��~�ҹwk�,����.����Wc����9���i�0��3������c�1}�)���&��y�,
vW;�����\�-��9���Mz;��7ntC��Hy"7���_�� w��L���o��r.7s#�����+��.)�Q�e��DB��ҕ��o��brW\�v��e����1�j�7�E�:O՞Ŷ����k�!��b��u�=L�T���%U�g��Z[9,�(��7u��rk�SVa�}|����9����T�R���#hB����k/����=5���5�����B2b��*�<é����-C�R�oa�nb���������SX�W�c�*�Ε���{p6�ߢ��;�"W�'o����7:g\CM�lumj�ea�P{����ɶލ&-$�*#)kb���X��Z7;�şmD/m"޲����t�\�_`S��P*9[���<�����<g�b��ǒSz��rALA{�/yQףq�ń*i౜��d3EL�Lź��S�xS����%B�EF�Gۯ8�x9�%���v�jX��.�Ь�Afhp]�:Q������]�w�֫�Kz��\������E�M�g�dy�3vo�nl��u�[����ie�B��K�s�O!�N[�r������������/+71�!WE�9�
�U�Z5yv���̥N���c��r\wZ�7.��y��v��o ������[ګ����0��Pb�fbH�d�X�Lİf�j��(�r�ꉷ�x��-[�ihs;]U���A��;��`W:ƫ�g2�ho�0:6��wJ[�N��'l���mm�8�R���9�Ë'M�+r;�'I�լ���^xr+O�FU�t׋�S)�*�,��F�y{ܷ&�^h���I��E��Q�0��q�Z&p`��l����o����֥j��{p!���H�O��2^�D�:n��Gk�T�����sJ+�-�CN�U��T�(,�W��9\��w���x�D��%-AYDn�j)�^z�0c*G$J����{���9(�d:?o�R�)',�R
ER(DH�B(��8`cU"�QH�
c
�b�������j���0�AE�D{jE"���Ab���H����"�ȰX��C#�H����2")Y
�U\K�(�����}�u�׾��5���|���^�\z��fW��>�U8\��+�K�_�>��<0���^y�n�p��>�T�q{I���ܑ�� �7ڥ1A�+�gk�5�	HԷ0a�q�O:ȕLu�WT�F;g����c�j
X"c�u�b:�ݰLQ�C;|�#/r�����H�l��K�32�u(�qn(-���x�w�����ޓ�8(W�s��5׷8��q�T.���ʽ\rIcR^c��:lToe\5׵Ԫn���ܿ{y!����R܄�Y�4F!�m���I�׳��7*�F3�jv�ʷ+��`��udnY�/��f��h��o�h���b>�\=�yя���7ǂ"�5������x57��̾�1�^o��uȩlU�S������s���^�x+ l<Uo^�c҄�5�`� *�&p���]�-���ٕ�V�̢,��^���ITw�{���늞�ZN��b�<�4���*��{�&Q�W�%G���GK�o�-�|��Q��~YS�Nf\nm�Cp��)JډڞS-�-<׵�:s��eK���7k�f�K��ޱ[�L�gf��!�=WZ��fwU$wo~�uc-�W��*eH�t�O����8�7�^�J�?z�W�,S��:�Y^�"���8���9,��SB�{�M���h�w��M�M�kj�>��7�E�1ˊݿ��p��{�(�ҩO6��V��hֺ�si��.+s�u��RӏS嫕��
N��Ҫx��5/\\L_q��^�3�\qm2�ҹj�+���6��l�
6��ս���5�����h�����SW�;pޓ�4��D�w���YV�]�3sF9/Nv��]n�ۆJ�aiV�I����j������_=2PO? �o��r�����pE����qn��+��k����/M♡ǩ�c�f�{n+9ws�gqHk���#[�t�ǥDap�\7Z��"WG���bW���Iཌ�-{�t���>.�gH�j:�%G���~��^E6=��rCA���eo��d������ټ��
�
����f�*/)�X��m�N��J�C�W�W��4�yN�,I���j�@�ם�n0�����fB���5�'�P�Q3�Vb�{br�zFd��:.n�E�T�����l�}�\�w7?L�K`��m+��\�r���Q7���+8W�v7�u���z��Xd�	n�;P�*/mG�/՞������)���
���#$�w��lq'��}+4���@�'Y�ȶ�d��Z���g�7�4��(D���7G�ޏ)Q��/{s���侭���諮YsEY��f�T<���J㠅�O&�z��ZSfAGօq�@�)��x��u%�tk����Ś6��@�ISRx ��xNo\7�6�+9(к�&T�74��%]b�0̆i��h���Hl9o���'5gҟ��K-$��	���q>��kyo���׹�H��*�*�*,-&/hu��mQ7s�e�뚡ݕo�g��ʓӞ�q�fT�#�a�K�y��p�43�*{�m�,v#x-�}ܮ��j�W���g�U��oH{�io��+d�7W��������F�F����[�wd]Ç���ls�"�q��i�S9����g6g��O/>���yZ�,�g�>~�y��k��������mn��';H�F�l3�o�<��.��u��{ܕ�y	���P�1����(;�~��[������g#Cmr�B#�^�Y11��HuBI�L{��W�퍏:�kz��"�����R��IԼ�S�t�"�V�=� �~��n�=���g�v�2I<�;8��3���Z�u���S ��x�˗{��c��f����!�\�'j��g� ȷ���aؖ������ĶGC��\R<s��z8�<!b,�f�Ƕ����	���+�\��ٰR�p;�j��:��)+TEnrr�#��R�lB�q��ͻ"d�:����naq~������u��?�ǉ�\+�s�N)
>}~�W<#v���1�8�uC��kJ�{�����!n���r����s
2[���W�r�m]��JP�v�1g܂��3(�x۸a���VOg���|s=�a�Ǩ���jڝ\�Ӣ�,�4�gM�e
�N�޴�ۂ�jϵΜ��QlX͚�ν�Z�{PkU.t9+�uMy�faZi�h��"�O*d1N�7X�����#��QQ�x�\�8[�[c{
��/#
j���{H�hna�fc����n��f�k��u7��"(���\ۻ',�������N�-����:��mztW�Em�{��g(�M�W�9w���l �M��o�a��Qg��9,'����z"��ټ(5�3`pg�F�V�6;�<�*�ŗ$G<���U���ƦRH��6b��ح1is��N�J�x!#�1q�^��P�͸�:�%��^�����#�Ef�K��k��/do4�=笭o�voO��΅�m�z�Z=2�ɱVu�N=Ī�g���ڳ�����Q콅��yɈjɈ����/gꯪ�3�n�?s���~����H����c�L���~�����5�y<�O{#q�Z�+�$�����m�ا+���u�d򸭚��J��:����2R�I\xJ>G'�������΂�y�"�/5��w"v9�c��=e��0�3��@澞�?J=`#p�+z��<��,ާF�f�'Ɖa��?6�C��3��Z�c���Yߍ	,ex�$[��i#;U��f�݄:�l&x��{+k�{�p�v�4���gz$w�>�\������UA�
�n�
�9-z^�g�{:#˺��]�h˻�;%f���U�\�0*�a���V����JkBZ��ͱϕEI���Jlx����"@⇯�;��N�wX�++�+��"��[����|)��g�c�K�&��	�%}bs�Q��]�xd��>`
���PѮ�Z�e]�\��H�W���"��n�I4[U>@rx�,��D4�;����5�[ۋ����Q����e]���tШ��#�}>P��`�t��*����r�Dr�|�5gr����=5&Y齘�h*�Cy5�6�c2�=�q�UڣµJً$ھU���ke%Ɣ#/.�b���"����w��N8�Κ^w5r�=�g!��[�7b=X��*�[�w�j��i�9����e�e3]��E�)�*��`#�Z��\�m4��L��*Wc�����).�e^.���ٝ@�˳f�]�a�wX���뵪�<�ş�wh�t���/�R��l�)��	��a�E:4�n���bZ0�
Nϱ���\���$8�+���V�d<5t�j�A1�>�*̘��l]�(�(W\W�`�����B%�Ohq<R9;��Yȳ��Ղn����"�9h��`�PTH���(��X�V0Eb$�V��PQ`*˫	�
���,���Nr�鐭H��E�+EJԖ�l�hE�H�V�keAB��AH�%b�b2.5D�(�G��8���#�xN�w2�Z1�L���p��R��l�}�G��������۵�qv��_B���� f#�pg�%�W�0��7���ϓ�k�;�F�L�2��q�eH�bM�,�tkl��`���+��y�t���QU��X�ἴ��_y��R�SOk�C}.��]c��'a|�����G[���Dx��X:�_��o�
n{�Z$y��$�N䞉�m�S��W��~ߺS���j�ݰ޽f��.i�|�=����*v���Wn��	��0�l��Y�)��Ip� ��B�/�zK�</2���'�rg��2���WޏE�����T�alռ���M�LI��lY(*���Ѣ��e7%jٺs;��7v���J�5�5�){9ea.��-�ͥ�+Z.�<��QAl�uڽ�)o��eu��r���q���]�V��b>�=��7�<5;���x�zr�"7�u�'k�/ʢ���/�i������#�؆}i�F-;�/b+9�Ř:E�'�6��fA�zTuU��!�N���y�R�b�p�*���(�޼&f�.3_��[�}�c�^W�(re�����n6�+�ž�}��{Ҍ��#���<�+TR&�=z���Ρf��L��k�c��,��]j�P��'7�
�j}�.ꖞ,[Y��5���.���k��O�S�z�*4#Yw�W:�ȧ�i������u�X���E�e��7����W�q�K��v��P�n�͡���Y��.��W�{P��\�>������2ۼ�;;H�&�070�Yz+�ТaQ�u�����=�m���T��3�*�WN��.�Ş��t#:[�\U'�u�h>}��့�Bkt�N�@�|^���?z{�/�g���>��b�o�1����r�݌��R{(�w'#/"�N��5���<׵7��H�]�;��ݾ��<���͝�P?g�>tÂ���M�j뎋�8��,�,5
��yt^Д�_!!P��*޻�u���`�|����x��(�t�^��W�$�Ǩw�/e3�1�uJ��F��H��M*���%cҭ���}�}J��ʋ��Y����IW��%e��R`).y�ڞl�ϝ�w�f���/}ַ�pӘw����  ���Ŧ&�3�o�����NP��L���=�*U����mf�N����;�ѕT���h_0�\���p�m��z�o�����l�j Q	��*aL�'���<}
�q�'�urk@09ԄÁU݃*�-g\lW6W.{2"�b��(j�`͛��'����m���ݰ#�6��Y�R���C��K��#������{}�)F��Y�#�S����q��!B����n�qB-��:s{b�;	��uU��p�@���� �$���{h��e�h'�Í�3���[l�����J��͑��TCح5:(nqv��f١�ȅ�J��&L��b�y���Z�c�<����\�I�^�7R�v�v�T��m��[�=	nM���Ll���Eu;�)ൌjq[x����VW��떷q9{��fݦue�>����홹���6��(ۊ�AQA#�묧��A�M�7��z�� �ei���a�Rg�?h5��N�F�ɶw<��'!=�v�oKO�s�oU
�!+a��Ie8��BnE�;x�	ɘ�q�[��;�)wH�!gk/氏dܣ��^2�%��ɲ۞9}f�d��޹�Q��2�;�Y�ߡW֘䞬��|w���ǒs1��r
��k{jY��b~�P*ei�P8��!ɋ̧��y�Kn��9�<K�-�Y�$M��%��R�!p��Kͫ}u��A�½���5��=����^�Kͬ�9�
��ϋ�uQZ��6J�ҙ6����WV������݊��ieK4Q�t�Bmc���[T{��u]��L��3��}$VQ�\o�
��F�R(�Q$\�(������2N?�=����qĨr�y���D�AUl[ج짶�uE�ɼ���'�φ�r���P��[0���C� ��{�U��r��÷V�=��1�{q7w�L��ѽ���Yyݠ<wZz�=Қ���ؐ��k^���ʇ,�o��]^�+P�-}aC_���M�����Z���R�a�X������aa�%�3��W��$�q:��M�^89�|s&$G#����w&閲'��� �(�.Wf\h��M
�m�F�ٷR�{ �10��10���T_z�"eS�9��׆Zuf��Pq/;����6��G!��z�N��1)��y�EY\�%���?Br�VwBu�]ط��k����*U�$X�]`7�$� ;+T>�{��svo(r8��J�t/������׋j��O,���D;{RA���Jk��Tq���B�����N�[W�H�Yc��-�I���I�Sg�۵+���yLW,�kO]rt�����/����K��ArNMP'rPh\�Q�|�M��LsIf���֨xB��=S��2�h|_9�V_$j�^e���2k�n;h�y8����v��9]�M��16�S����;Q��ƙ�M�ػ3nffL��t�*�*Օ�uyQ�ل��܍KD.`�UHu�o4�lʮ��vw�y�f�t��!N�f�xV�c3�!֕�n�a��v���f2m_yj��at��h����b�85�P5c����^��U$U�Ue�3����Vi��������y�*я�q���ٽ�{�^MAWu(�i�v���(#|�u��4*6e}J�+$<��:���UzV�Xn����>8�;��A���Tj��Q�ǂ�*��0��à�u�*o�3ܒWD����p#�ʓaX��5�X-m7&�W�y{.I��$�e;����}Ո�6���hCT���.ŉ�T޾�u��,�Ĝ�u���b�s�8u�as�"q���z��2O\6{l8e{yl>V�M����o��	�i~A���.����9ݘKW����nŬ s]A%=�Bػ�7��X�%�X��o(r[��`ˁ�:���z���Yz�f������yW6��; jI�*������Y�9��C�C6=Za�(C�cC���e�5lN�/si����r�T�t�Ys8�GPZ9n�f�{�o�۳ΆЫڕ|6����Hm�yB�f�׳1�n���;�Xp��Ꭾ3,��r�*�r�(����e���s`U3tl���9]|�u��Lk���,�+bq�yRj{*�ٻ]�^}Z�I&ƫ�,թ�wY&��*k����5�Y������@��6�hZ�[���V?�;�@֬P)�9!��b��*��C��Fۭ�f$���7]Q�2,��"�rwEDlܙ㪫�˱����uR�~k���
D`��(�gIF
�A�QUM5�E`�)����-TTAb�:B�b�*-�1��Db��e��*�����DՕե���A�G-A�d���*��UL��)kA��h�԰Eg�EfkplVe�\��G3+�Z�+�S+�,��QD�Yyv<h�h�p�yC�ۇs��^"�Z�u�6J�!gl���&���Jj��Vt�O�GŏV��q�3C�לN-���IM�]L4l��|(U�j���z�L1�&9���� Y%2�
�NR�--nt�{SW��O:)#�l�y-m3IF3H��4+9��2���#�{d'�g�v�>8-��>�y�a��q+�\�vк��Pl��$^�mY��z��髵��RU�:�H~N����{���@,���C&_on�t�SP�V.=z`'i�����
�Wk�v0F�m����C�:�X����ޗ�dJf�'���s�z^�3�{3	��X�o.
���Sk+��]p��y�`�9�ü4:�ʍ�W�p�N��ʿ���[��g*��8��3N�G��ᵭ�J�֬y�VvUn��C�y�7N2\��ٰ���+��w�jI��nR���U�'zi��f�~K0F��I�.o�;źz��R۝�{��DO}p�y~"�lx3��K��L$��]�]������y�|<B ��	�����ƫ�1gi־�ő�t;�#�|⍫T��$48��=��ҟw��/W��jZ�9E���yk�{dw*�Ԅ��ȅ)��.St�Χ��ϫٽq��r
*a�}�֍6�v�[}r�	Hm G�PY�׼�&�`im&�a=bN��cֺK�jy�y<ͫ�x{s�����\|�+b��X���y�\�D��n{q�dgq��%����&�Yq���k�ו?L7O��T|V�2<�Wܩ�$v�;�p��Y��v9��RY��(K��^N@�ҳϸӔx��^���J�wԖ��"��Y=������c�C�C���r���x//N�=^�#��O�-�������mh�9p*��s��jf5�{T��O$.�Ʌ/��:T�nv]h�%��70`Kf�^cX���<㖣��s<p�C�wYs�Guhl����ͮ�0bY�� ��
�1C3���V����\�������=��}�[���ytm�ÐQ�jEV��2�J��	��!�Ŧm�� ���$����.Ӎ�^��߆{͌�n�����[��9(�{�K���1�*<Ѕ�\t^L��A�<ú��=Ok���n����Q<oԕ=0�jj���|�:MWs9���u_�����%L� Up>�j�tջyڜ��U��j��P�g�u�Ð���q�qk.�x��
����������+�2�+Qu^�lce���f)~���}��L�{.�^���4�5�<���Y��bЖ^�^^J��c�ѤO���?,�+r��+o�R^�|I��s�*
8��ج��ov��ۚs\�%�
jr�+�,�T^���G��@]~��6�_|C���ݺ�z"�����[�tg�%��EQ�����J�b�!���1{x�un�S��E.��a2�GM�ۜZ�ვ*&�R�gXFrU?����m��X��\��T%<��W��k+��������²^��]Qy�GH=kώ���!����|\Ĭ��#�r�3Y7+ʅw��U�U�����آ���XGAp	�ga&��C/6S�h^YNN��A{��������N�S[�d��/^���y� �6o-ş�Td��{\l�+�v�jN�p�48��GI�tf�Or}$���v�I�o3�����9ȵm���[��v���{b�Q�Nً-���ݧ����o�ὔ-Bz��"�ˎ�L(e�Y�\1]p/�B��r�J���>+3;t>]�2�*T�ﳐ;�O84�ǍР�c*�c5��j,�@����O>����EK�S��7�gD;*��j�_>��EN�'ugj�T*�k1�)0d��#�zm�A���������/e�r%~��j����;��89#/�ne��e�ȭ�r!.+`)��y���>P��fL�ɭU�5F��k��+�_��õ|sa�]��GNb��Tv���zkgf򚓜�-�Î�q�.�:�Z��o���� D��ke��)�]W盹]��G�^$��2�n�{�ͤ��H�4z�+��mM&���ߋX*��h�O&��\s�E�o|�W����s櫵�ı�OF�:�uii��'�;�v���6x|��g�.#�jWK�t;�s�­�y���a!�}6ѳ�G��)A��q�}џn��?zfx�PE�Ź]լ+x��4��e *�S��y�^��	c���p�p�����`h��j&�[^��HE��a�g&45�b7;��-,au��Y�ɕN8��C����8�҉�q�ٓ �WE�^�+���m����'9����̋�z%�k�f�g�d�9�XQ��YI���m^��ͯB��mOz��t1��"έ��g�2����-<ӧE}��%r�x����wf�2�+��xy�S�6v]�۰1��d�Ms|��]��Dl?T@�5�'cg5
ɩ�CV�^v��{{xN ���v��ΐ�Y�1Nޣu��f�5�9��I��K},���u���|r����]y��~{���Ǖ�¡ S:�]����F��A#9\]U�T|w����{6�bK5ro��qv����7��`�f������,��wv;�w_������i܁5:�5r`�Phs�=�n��<o��^Q��]xy#�Ҋ�7Ξ�2Y��f���vg3���ڝ��U�n%�ӵ��c�-K�M���e_`j븕c훖#ip���|�ʌ�i�}�V�N�j̊���lZ+��2.�o)��u��\�Z�Q1	���r�X���wQ���;��[[���\�{;}�h�׊�6��o��@:���E(����H�rB�ҽ$e��oNu(q;�'�
�ӫ\�Y=�tG�{���t;}�+u�L�ܭ��k���C�V��[�B�f�����ׁ����e-Mf�~����^��m�d�S>�<n��T;��X�������!����Z�Rrv4!\z%��=X�wWe�D3$3��p���>����쥀s�U�\�_��+�SP�:����XUy�{o�63�S�c�6:�Y|t^���N(�ժ�p=˟_[U[�R�f�ÖU<�H8ټ��
b��E-;�;�79N\��/)�٤a�^��U�zA6 �b�;뗙�3�I������Hnp�:�^���vN����!����{���o`*�vT%� p� �竑},���h-:t������+wl��ӝݸ���j^��s'��zr�=֦������n8r$�U�u�y�1+�˲�[U��sF�+��:\&9�3P�7��"*��׶��2�roW�����es��b�@' �	��E�k1�J���j+l�*��a�CKJ"�5�X�2�

%���(�YPX��Xj�:�$U��B�F�+V��\ԫ+R����īe�V�����d�P[KmD����I�"c-e��+���0�X�M3Muh
l�B��uس���iK�v{��U��Ms�79��U���s��U�	{i�]y:o�zg����W�������H�xU<{o��ޣo��sw�E��n��qy،O�oa�f�:��y�;�
��h�\j�{����;�Ԥ��t�c�����e��7�)o\�s��Pk�']�F���7]���5��d	���yF�ˌ�DU���5E�&��B��G��bv[�@��لu��u�z;2�V��J�K���L��^j��;�g]h�P�q�YЪL4[Q�7���Q�APwhUSg j�Lh�1p�늠X)�I�ަ�`�}{1ƣ!���|z�b��L���V�\,נ����e�>���|J�}��lyЮ"�{m�m;֭��Ӿں�*2�p]0�[oX�_�������"�Q�!F��!ы�U��}�#v��nX���|r�ZǱ��Q�d��Q��8U�Ha�K�罣���z���*�^�/0B�W__��Y4�7FIv<Ƒ,������֊�y ��N�E\׌\d[=iԉ�͌ͤ�1	C7�����	��fHd{�cJ�q��S+�"�����/���ty���T�\�\��@�xQI�g0](1P�gkB���0QXĴ��6s��&S��'8�/4��V�e�A�DQ��7�[�A�j��yŹ�ռ:s��1�{��E�U�����Q�t�i����*{i�9V�sZ�U��{*3�ύԗ�F��"�F�^�tn��5y�v����Ξ�R�1�7�{��n��;)�iY�.�(Y���Ac��u36����FeE�8�-6�RG寮5�c٭���Օ�S���O��y\;���G*���S��}E���E˞��oS
y�l)h+�x���R�c��1��1n�P-������B�u�[�S�;����J췙����_��0�ʋ��[�1^.��D�=�p}�}=��fi�8��Cv7t;�}��'l��V��0)[t|�#7�h{�tا�����[�W�a�[=y�N��S�-(�#F�30�i\Vh4VYMǌ|=�G���g����G#��7�g-��q��c�LW �.�^��o�>����t�e�8�an��P���+�6!@ܬ�������9�ߤ��~�D���k�����[���+��x���ў�����t5E���^z��FIs^s1j��E�u� ����#&��ı�l�A�2�W���\cݽy��K�~�*���E�,q��[x�l��s1���,�����>۠�BS�oc\P��kU˯����~��u���=�k)��	,`��9��i=�L��W_pY�
ᤒ�Z8��L���[n*2 �7:qo��6u�[F��kzc3i7�Q��!��p������4��h���� �"�8S��R����p`���'Y�#W>Ξב"w,���uk�`���^�����Q��wk%f�m��Mu�Q�x�Ð��wHj�\vhNQ�il���])�f]p��J�c^�~tf����6^�t6���{&�r�7Ǹl(ǮT��->�ŐVP��Ц��R�Uw��BU)�;9�nS��5��-�T�L�o�:��u�5��[�g(8j�7�]��z�!r���w�5�����h��Z� (�N��X�rɁ+�a�M�������m�8S��+���[<�f *+Z��v�nAP��Q�dռ��;��y����=��6�w���P�\@����x�%��*;���v��;7y���ɯ�O�'�'uh��V�����,v�ū�0.��gw3M�srʿnx�k�5yQ)�z��q�S�E�\�m�=;!휼���Xtr@���G>���]W<�#rK�Qv��B8���[��&݅���
[���cS����P8���:6e����ݣ��!�{�x��|�bg����(D�(�ƹ����/VoC��⻭�L��j�r컄�7���:c�	�y�\���n/}ew&3ʰ!�U�t$�&Q�J����g+�eY�8�C�g�˸u�܆=���\�na��oҎ��;/��=�㱎7D�D\�����L-}���9>ȏ�	�(ͱ��v��+>��>�c�1,r��f��/Ou�Z�\hL+V�sWt��M=��&6���<pNc�n�^�a�=9�x����O����#�&��a���.�:��w)^j>p�49�L~u
W��|M���g8t�9��*Vm��y(l��S=mi�F軩���/���</2ai<k��?f��Ўdb莵z
�]��u�Kk_g�,��vqsá�::��ett~��.��oO�sƬ`P��9�G������3�Ξқ�O�]�B�_���v�zG��?u��3׏ր�����hv%�A�d ��N�+堷�GI��7���Y��{{�_Mgg�vR�:a� iя�;���ҭ����^[犄�O�t�_���h��ʍWM��$��%+՞|��~�����]�v�w�^�eyq��0��%�kJ��k��ڃ]��N�<[����.�)�ŷ/f�+��1M�ˍG�	��V�Xz=X�K|u��ӛhu�W!���s�E���`ҟ���+��~9��Y��zJy=wh�٪����z�S/�W��R.uF�ԍFM*��^�2�۫R2h�%\5��!���*$��4q2��;��]��E�����\8��x��"�tܨ�Tf-�F�K7y�@EZ문2n��4Y[�eX����宴��p�U!����-b� �t)a��V�y��=�-�g��K6���.��oQ����
����媕� k/KG>�K���F4kBs��#}QÂ��^��kC�-���\s���<`�>�b����m>Ivf�TC�������[s\���F���]��E36��\����X��to��Q���,�Ӫ6)�fS+('5v%�ݴ�6�ѳ��N-ԵnН�jY�N���l��ٻ)�3;s�M�q����9�����K2S�2t��5�&����$�C[:��n�Sj�I���+v��u�D�\:t�D�V��v�N��|�kJ4�u����}��FcB*n,���|Nȟ�N��ml�kQ����e���a���]:v'�u,�� ��+*�P����ۙ�s��4zh���2�7.6iê_3rWD���ڏ�P���v�\��";���T�����hv���^�R�2*�hˏI�+���Νk��J	w&U��uc��z�K�i�tH���K7�t�>썈�Ʋ�i�����2s[���{�]o\���g5(��b�PP�VQ*x橥t�iq�b�,�4¢�-��VH[��@W)Xi���YIGL�J�iR�Ȳ�B)��ePa�M$+�V��0�
ʙZ
W��(�*,�XQI�d�%Y�.U�1P��]2T4ʊV+Q�^s�u����x��q���Ü�G��eI�{Ӥ|����=�@U�8�B��"��d��؊/��WL}ȫCG�L��򜙘�=�[(m�"�D�QM������B$Sھ�L��v0��T~~�vV3a$�,a�~�R^��c.ѭ1��T!8'�M����¹�ޓ��;<|��u�[�yL�u���>���l*�W]gE����^�^z��5�����5%\�OKojx��Հ���ʕ̲Y�S��:�*9}��o�q}%^��KfR�u�3)� m�N@��	� u�js����ߘ���;�7�+�}Nk�㞏wg�(��q`��Iʝ\u��ج�^�Y� ��H�󫵃��Ldq��`���p�z�eTK���y��T%�;���9A�/�!�V�=]�s���� ��>j���p�T�w���k�4H��Y|'���L�1��x���e�Jj�w;
�$�>���5a�2�&��V�Hl=ޜ��ڿ{��Ж�5�b6OU��� ��Q{/uMX��(ex��k��B���0�)��'�{��B�ݭk�|�rQ�+��K�m��vz�@�.���8oX�[g�H�;Ql6��Fl�-�ܭ�(�5�.{�m�L���Q��(���Z+H�슼�~� �f������ݻ�II�B�
��{N3��*��L�]3{�r��i��	c�Aw�����o~}�yV[�;�cS%O�M�&�h�5G�^y@Ύ��Vk�ǯ�0��ʹ��^�ܩ+�=�O���̳�\rch����ɣ��*
r����uvC�^�!����ec���ds�Z�'��=�a~���籆=@�ͤf�5���ݔ��c�D�Tc�gZmυ-�$KlGS=9\�}��c��[]9�7�[Bqf��,Î�°����cc|��}w)�&�f�s�u�Ok�	�x�)����ڼ���(�x�x��ʇ��9M^�ǔ�Z��#���wò��N� I��҇��6��i�K��ݮ��a��+��Q��t߹���׷������c"<���/.Lv˞�[n�u�����,�o'.l����]y9��z���!?�)��ޙ�����l�6���}�w��-p53����
SGl�ޥ,ʊ�^�����]{=��#&�mK���)���r�~�p���Ʀo��a�B�ȫ;��p$ڇr�����+iU�� ���S)?��KI�Ƕ�m#%�=��2�m���+[S&�.�h�q�]o54x�W��oJhB�����.��:ˬ]�D�\X�&�wLӋQ��]V�ufNG��,wMRMF����K5<�zu͊un5~��*�%��EE�`�I�k�k��un"���Y��̽W��Q�/1�vn��X),.�оds��{�����چ��D�T�㷉���<�]g���UI������w�ל|�_�nh�٠9��y7Jש�@I�qeNG�3x����/�W��؃���bymQ�i=�r��{.�4޾ֽ=�y����V*�Ojzb��r���z��f��qR-��K�qEIWv2I�<a�\�Zީks$���(���\3\� ��{E`Ö����(�}V�.���(W���|I�o�sQ�	Z+��GeF���.�֗�9h%c#��:�^o�o��f7/��_X����m{��T?'w���0D|5f�(�?!����aV��"��ؘm�sU�貘�gm�;{�73���1̦�S�S��k�68F�k�m�{�N��w׽�eY�ɂ�V9��N��ax�>���������Qiq��mÂ��Cǘ��[]�/�a�5��r����oB�*&���u�i9|j�ٌ��6m坆�.�ȾJ��jk���f��1j�z�e�Rڷ���+�������:>?���`�Ҵ�s@mN����q����$>�T+w��'J�=���xE��rc*�Csռ����!B7G��q\��ˌ[�0�$����]5ݰ�\���� �6�m]��S�"����!f/*7�r�h�,zj���U��a�rv-�|rv�����э�p
�WBb�,n�`�g��W�mIW��{�:�1T&u;ڢ��,]�d�k�,%����؜�f�%��09�f�4�a�@JA��D����^�׾,����!�N�w�8��nxhLt�ACZ��.��<LZ��K̛�G��^�{Y�a�6G5��iἛq���\�W!�� sL��j�8�ϊk65�ǏZ�����e���G�b�-��2l�6D+#͑�+X���ӞA$�W����4�b�z>VYʼ}��A�(��Ko�����G���fXQ^R#�؞�=� �k�y�\�vˉg�`@H4�}2�-�-\~�(��ʼ�J��Z�Q��kQ�y�3�����. x�s/N�5��U�Tx�x+�
��X��cE��̤=	*�v�zF����;���̽���E[IC��I�J�^�i׋�z���{����>y7��,��ts�ȋp��j�싶��xl�8���q�3m�����B{��!N/~9�ݣ����p�2t�6�,�R����v���������w��͉��/yN(��u�i������O������� I�??��O���grz	��x�,` �Y�������CLa���l� @���
!a�g��:��6%��C�B I�4�/��Nߟ�_���'��9���w!��:>�i�Nӣ�Y���Î�^�GGa��;��=� I�)<��������!C�p	?�2v�O�C�XE���{�������r~�0O��8�\���G�l>�C�)�~A$������r
��ɜ�b>߽1����	7#ԟ�/��X��Ĉq��I�>��b<�?���	?���@�G�=��Y~m�N>�~���C�t�	��L.�/,���������-��!��p��A��O���ω�D���E��'��C��g�I?��7����p)�����A���A�!�|gV>��?8|q��?�����/��6�:%�����~��\�a������pG�/�?�������#� @�����g�E���q:�6`�'��DD�!`?h~!$���?�"}.�zOšd�pv~��h?pvtn������6H I���b���2`���'D��a!1�vM���}S����쉽֥��<H�2N8��`��~�M�V����$���>���� ���� I��|����O���I������{�|��g��|��d����D�V?_�ϑ�@����������|�����C���@�O��M|�<�_̄���@�O�O�h7�ɇ�23�����D����	����M�8CrG���ѐD0��7��P?(w�Ϩw���?O�>���Ӊ�a�7�n@�O����!��>�9�~�60�?eO�����.��ߣ�6�P��l���	��Oݟ�?_� }/�~����>`$}�}'�O�a�k���)8�x'BM�}�['��I����(~Hw��rE8P� $D