BZh91AY&SY,ӭ��g_�@qg���#� ?���bI>�        x �R� � �  P   ��   
   �    
   �
 �T���t�F�3,�֤M1Q+mR%���Z�jY���DV��m-e�5���ZLhKk6��L�l֣-hƶ�a�ʶ����Z� ���J����Z�1-��,�Z�֖�e�e�ћ
�+B6������Q�Um��6�Pմd����d�l���4��Mf�%�gLژ-``�   ��U4Hj6���:(��m�D(I�kG%U�� �SUWh�$�wV5]Z�h*�Uj�Wm(l�R�$٪m�Y4mX*��  wҊ(Oqܵ@42L()K�˕ҀR�����T�s�F�)J��]T�n�J R�h����E
wu�h�ĶE�V�ͩ��   ���)@I:���)�qΥ��J\q�T$(+t;�R��I�ox=(HQ�I�������k� ^#��y��(:���w������kf%[6&�k6�4�  1<=(J�V��t�4	'�+�PUD/T��J�EGW�<z��m�w��PT�-�EK�m��w��m����:OW�x��^K@��$Z��V� �� OPUu�=�4��=S��#���z����
Q��� uJ9���{��+����=@
U;x^{ݥJ���:�Ey�ց��f����M[D���  �t�A����Ҁ�j��hJts� ��J	�wB��R���(P�c���;U��)�4�k��UA[���Y����Vjٔ��RZ�x  oP�m�Ӛ
 �X0A��k�hP�`�@���:�@;�\�s�ܡ�s�p (�0 �]�`��kH��U�$*�  �� �\�
�vp��Ƭ t�w�7g  7v�ՠ n9� WMݎ P3I�P ���-V�)��6f6��6�x   nw��7;WP �g]P�P ;N�  �ت k� f� �qn ����P\U+I�"�i��k,�F��   3�� ��Z �� 
���84(�0 ���: �k�PZu�P 6]8��ƀ��  @ � j`�J�&&`i�&#��)JR��#	��M4�a1���Ԥ�P �h   ��$�IF     4H�4F�<�A	�M�驣�2=i%H��J��     ۷�=�i\�y�t�������W
_b��	��
Z/�	[A[�*Z�+y�#	]~�Q^�AVT@T�@Eڈ���M]W��8�_����!�PAEa�J"",LQɇ;a�f�q���$<$?���H�����!����!�^����	zK�^�$>� :Jt��= :K�������'H�t��IzK��%�I��:a�/I�=%���H���#�C�I����H�%>� :@t���_�LH�� :@t��	������I^���	�G�����!���/Hz@t��/IzK������ :K�� :C�^������H�H�$:@t�����$:B|$:Bt��!��������C��I�$:Ht�����!:Ht��!������C��IN������!:B|!:K�C��I�}!�!���C��Iz@t��/��!�C����IN�=%:Ht�%:JxJt���G�'K�!���IO�xH����:J���S�/C�'H��'H�%�!�C��HzK�����$:K�C��^�� :Bt��%:Jt��Bt���S�'�:H��	��)�S��H|!� t��	��'N��$�=$zJ��	�S���H�N�=!:Ht��	��I:BD)���E:@��QN��t�S��$P�'HU:J�����HQ:J� ��= @:@��N�'�P�t��(�%D�H)�@��t�G��?	C��=  :J t��@���t�O	@�(�ID:B)�U��p���%�*'IP�BIQ:H�DN�}$�"IA:@	�N���:@��� |%@�(�H:H	�P�t�C���%G��
t�� � P� 'H:J��@N��t�C�*%Q�
�I:B	�T��p�C��%� 'IP�B�HD:B�@��}$D� 'H@:J��Q��}%�
 �"/�AN��t��$�*IA�!�N�"�B�QN�
t�W�*!A�IC�zH	�D:@)��
t�� =!���I1)�G��HN�� :K���X��H�������IzHt����Iz@t��!����HN�������=%�@t���H�����OH:Hb�'I� :@����H:A$:Ht��!���%:Ht��H�!:Jt���!�C�����!:K�C��HOI��$:G��$:Ht��)�^!:Ht����Ht����!�^�$:Jt��$�������#�������*��AT�uʡ��Ǜ�N���� �6���������RH�N�T���p;:�20�h����*B)e͡����ˬ�זN_ ~�M�c������K�b�Ϣ�H��q�('�?�Gv�l��ZD"���QͽʽS�����|l�Ce�y���\����a�G
��Ze��>�"���٭�^^��w���l���<�����s���1���t��[���gf�4�A�d;�c�J![yv2�-���c��h6�
��́��Q�P�a��p8�&kv��<�Dǚ2'�ht���֐�3Po�b�j7���	,*R1mUǗ�cA7xP���q0F�S[sy��%a��nΙ�|�L�8�X7IR�����b(�:�V�jk_���ܲ�a��e�%����3KM�2�Y��۴�� 6�nv���pB��C:�ag^G��(CYA�wsk�a�Wt���m������FD���S�Y�^w��	<�.:�TN2�X�����5�H�7�͘�)�|�ܦ�Omg������3Lv���n	}U;\�l|K�܇h��J��u�6�ou�a�1'���W*���1)����<&�r�n�
/�<Gf�7��Z,
32#:^!9�Z�(��&CE\�q
"u�.,gy��;5�/A�����˼De�������;�*<6�a�'f(o���ق�ꅹv��t�+a�2v�n�rdΥ}���]��s�)�׆9i�|���7��e.b��`I�6�ͅmt�c�7wR_<��q��ݤa�T-"�X���w{�v�tB�h���h7+<&l���t&�P��"d;n�K�,��g<AӾ\hVe~�z��(g��Θ��:+�0�up�;���ԵnD����s���s{$��;�e5��2בŜQ���up�q�5��ݟK�k�Ȭo�����%�-��:�p%���w:,���ta��_�����^���;�	��}�f�
W"�^Lvl�عʤ��ۜ��Vr��n�����UF��T�
c��mX�@sU9�]�)'P�4��+�4޻��bJ�N��]��޳�����'���E� J���U�i�kΏBȈ�+�E<�v��O�ˣ:�.̰#YXָ́��P� 8	���h��^pa˜�6���^+�z�2���O+u#I6ڎ*�u��Bu[�ץ�#Y�ed",6q̴�m���V	��dJ�cM=����K��&�
g �
AmW�����w7��Syq�\��mc���¾j��V�$�oJ&nM`�Ҳ���
m�2�̴L�n�� �y��y��okH {ǍS�����Sˡ��M孩t�ܑ�����΅@�᝛/1�H�9v�����.^(��x���I�^oB֝<rݕ�i7yo1j��[Nvn����gv��޽��Fm��v���"���̲��a���,y;P�����H��,ǫ�r�\o���#6N%j�g}���sx�Q�y�,�v�/79^�v�<��a�t���4�4��ٸ)��sR5sMEG��k�Y�.:j$Jc����5l�����ke�/E�u�������bP�кg6��7�
If�wh�Â�����x�1W���q��ex[h��K��47+<eS�[���s6q=�tҺ;'÷ ��𝣚��;	ɤ�@ɸ��Q�40塙���!(�sx�ި���8�h%k:!+�J��o2�,�ӏ�>zCG�'�X2�w_���46u!�u�S�?�ק{;�D�v�9"��,��o	��r\Uq��+�;�+�F�e�&��M�^J�0\s�9��PMcpo�gr�nZ*�����!/W�B��v<2��P���;�-�5�WR�U�!#���V&�Y7)��F�cIs�BV`�՛٠É���{p�
ܨglƎ4{��W�w�=�n��=��
��<#���gh�܉qdۋ���B@g]E�yNBeR�̻�K�i"��w
 U���k�fM�:�Hf���V���ݧ�j��
0��V�ϑ:	�`� �{yc�p�hre�5��|۹���9g�o�M֭��C!�Tq�h�1�=yE����v�� .�$��y(圦�ń���]X�o`l|�Y�<9:ξeCs�a�����֧d#B��j�K�A�
�Q����b����ٯ6ˉ��7��]���Z8qgL88��G_�#�N�f�H��me'�Bۂ+{6m���X���1��ٸHO�m5؉��Z� ���x>���7@�����Ҷ������8Mwq��5��rOo���L��V7�$%�V��M����N��[�%`�ys�q-u[�Z���v?��5�R�8�T�����ov�e/#�2>�ݣ|��b��$ ��0޻7V3��D�c
���R�J �ۖNɓ4�)z\z��%W7W($'���2u Z��^k���y�A�W\���SM�v�At���cv��Z�8�o���c�
��{2��Lܱ�X�`�1F�'�Ԥ�D�R��[V�d�q!�vt=©Rkԋ�F^C�i��='}`�]�=�R	��a�N�{R�Kl(����&���TR{YK��&&$Wӽ��T#�'�������"��*U��8� �l�ݕ+�ސ�v�x�:=L=D�{sn
/n�V�׵�j�v�Q�y0V��A����������(�c���[n��<�
h��V(�5��wy0��l�]�ƌ�2K[Ǒ��כ�b��of��j}��g,qt41;�l������K�ŭ*�upc�$:Ź���s�5ɕ3w&�>�)�M�Ԗ����gE�p�N˫�mY�7	·&Y0o'�����η���X�%<�o)�R���幎��ˋ.��h�f�r��a�����[K]��Aꨫ�޸C�; ����S���㈜s�y�h� xXV�Қs��Hŵ1��Ѥ���,�,�gȲ���ǵ��}Ӱnv%:gd�oM�qt� �3L�-�"/Pݕ��z��l�{�M�t���<���$����.�eM��Q�sֺ�屾�
��ݻ��_<�od���Y�I�~ںP�/~.�:��.<�p<�Ã����m.Aq� .�}gz���d\7�v�x��3svn��Ds=�&qZ����u��SslӻHL���On^�Z�kv(6Zj�"��Gd �!���ǖ'�L���r�����7 �y�i�v���}������X�t�Xª���:�G\�I�w�;`�yKٹ����j�f�W���.]3$���c5���& �ێ7���Yfm:�5�O6VXu�/E�T���h������xh��To.�om����y���w'��v�������Rm��X���Gk2�w4;��ouN͓O-��K��D��,�Ku+�N��Q��2�&�P�FP��.]#�_m��g(���fŌL%s���,��檴�ާ�1|�ˑ�k�Rq���.c�i�ټW;u�ь]fm#,��m�e:�ݨ=g7�����)3H ��۸`�˷$��v�tL.��I-�jt���a��Ƭoi`��m$wn�@��ts�[GvІj���#s��콋���V���'���m EK�E�(ML���e醂3���������n:�Ν7D����<�-;I��2�b�udtyE��nl}�95i��Ȳw9z	�gf��%�,�B$��R�s��u�`�K���E䱣��s�f�P5���R�'���4�_+��(姱l��{֒�9��{�1��1&��1g>!oe��Kn�]ǥ�o2XIŇ�_.x#���+�*�R^T��w��L�+��9�d��HUy�c\Nʻ��b�FT�
e��vL�orN�ā�	�/��6Œ��GG*F5��J	�b�F��<��d)��q��ǰb�a��Ԗ"&�Q�;�Uz�D�6i[����z��0=�S�{���ktg.{�5�L��a�P�X&���&�j���?��4@t�-��^���Z�.%p�X:���Z,9^M��
6�o*��GdS��>��X6��E��r�2��7`�����͜�]��H�W�����RA5��<!r��J���:���m�`��W9�%�f���`�����@��E7R�u1;-�f]����6��6��4ר���g�O8�c#uLX��D�!��Dp�����z�ov8�-&�/��K���>�Y�\��� .�M{�&FoQ��5(tɼk�'�L����QP�F�<$��������5�cy
2��Y��H��I9�c�)$��(�mMP.�2�N�頢{w��!:ƞ�!TEH�;���Gݜ*��K���y��sY�����ʵ]㣟-ʪ<�]��q�^Q�+�1Rc����/ Y�k�5p<9^>��VOs�i�u7���`���S����E�A߹�N���Z�b�,���f��X@!��ߋ�ٵ�Y|��a�����OU��r�zο�r'7_k����R{Qn��V:Vt�K���n�*`�υ��y��nEӎU���k�o8U2��p����6s5q{��]G5��tr���an�,�i��5�C ��=F�7��K�s��nl�:��$w��ڗ�heN��lPhV���&��q�(U�'�>Ӥ���^o.]:��w(RI�YՁ��L70������1��Y"�����Ɖ��X	���(�Be)&M��sF��A%X���k�nC>��˕�>���{���gLL4V�k�G\j��}��c:1���{��G@���Ρ�.�]�z���1Os
8D�{���)��c��Gλ����u����[�=g�@TS�����]����R-�uG^0��K�Xi(��3�}������� ]6�ɜ-�/��$t����S	pz��;)pcb��E�x�>]���w��@���&]+rt|˺�kUn��E�m��J� �(��k������j�U����J����uv��WU��^�YK��hd�ul]�\9VX���'���0���ذ����\<��d@�܋~�]�g<x-����	�k�GS�1:��N.��ؖ��w�nL�Ʈ�гi�Զ&H��Va巰cRd@�Y�p�6�v��	3r�E���Ϸt̿.u�ǚ��Ǹ�/w&��n�\s��z��.�hY��֨�`:�wF��=J�$�}\'�^��<�Z�y�(�� �n���}�`����>n�+ݥ�Z&�+kBŮ�-4`PS�Iã��1�]�r�M�ܫ.�,`�߻D�'��&�^��vS�n�i�T{�[�^�v�i�v�2W{e^�v�t� �FAy�K�6^a[��AK�]���(,8����D���m"��xH%v��
�<�k8�3�d�ow��B���q@���E3�tA�օ�h80�	�|� �j��B"B�����Z5ض\{�]ʓ�r��֎{:��L�)�xr͌b#��ֻؔ�v�W�<����ko�q>�YL,���͡%�d<�[�ֱ���e"�ŋ�%7�
�A�z�YMmf�v&���Tj9��lo��Qy;� +��/���ۭ�p�5\���u���� �b<{e�;�b+N�UNص�9�i�6���@>(�\����S�w<ۚ�gA�^�ƧN��>Ӊ��nqr���t�0����zv;��3y�e�p���쇰c���3�����E�������Y�I�9�|�v"n68y^���uo;�;��yS^S�@5���-��:N��7\��i������"�c2�t&�+媨wr9װh:ʛwz�M#���vӕ�#9�緻jS��y�DE�s{&ǩ���q`��֖wHZjů�L��*�ï�3Bǈi����t<�M6ybլ##9N�q6�1�[��#`��rB�{���
rӃ���*������:�跸Vt�;57�,*X4.HΓ
��^5��^�ަ8�q޷"�.z��`�H�Y��z^@֋l��Q���Ovp�5"J��o@����p�^�vHm��}�դⷕ�������l��&�JM����&Td��ß	u3�� L��hC7;A���u����tܓX��avMz���wx8����,[��Q�����7�.;My.���v�7�����G�9oҰ���&@��VRR���7��J���׎̈�N8ZX ��eUe8-<�����9f�L�Y�n6Q4��F��a�8Q��I��,��:CE ����(  �S6i� À�&�ÎN\��l0��w묀['X�@h#� �:�iғ'�ٌc�1�룤�ȳǉ����F���@X)q|���׬�����j��;C!Ç�q�ͳ-cӱ����d�d�B"Xg�XIo��%l��>����!��v��E�4Y%�Q�,��� ��C�)���¡��$�׌���� p�z^ �1A�V�:8��$��82�,
$�pѐ;���<6@��47`�ց��$@Mb��kƁ��Q�d��H�-6ӵj�a�O �E�� ���)i��f�ή�4��	�  � d柀��,�.sHAa舆QFʗ��	���l���h�N�7�GOƫ�hq����D�������0��o���P~��ܫ>�۬��nn��'wE��kpq�q_;}}l�/n��6!����.��v�`]�VX8�����hR�z8u���@��f�8���]�/W��l�r�l�V�S�n� G/�ݾ������ ��k���v\�0�3����������=�K%d����
���ٰ���[t�E"����̻��h�*��Cս���H�|e�}*���[��\�q"�.��!;��'�kV���
�@�N���{�1��v�ȽdM/T�{ b��q�9�s����ܧTjq�T��V�o5Y݁�nqb�h�ԕ����Φ�ъbv25�f���&z�uU�B��L|;3��\>;��ŉO��x��n�H��u/X�
�ق�m#E>�9w�Ŷ�׾����>���8^��	���6yZN��aX{Ef|}����7O��m��{���V�����Օ���Z2�>��5��TY��GS"2�m��6�U�XˣT��j��HP�/s���Ev+)6�ʚ��۪5n޺�m�=�����0ӗ�3��C e<nuP�O�;�+��׉7�{�a��x.�;Ⱦ'o;���)�bn㶰�tzP��3�Ik����
�Vi� �'v�X
}��;i̋]���(8�S����Қ�}h5�_<��M����W�
`�MAZ�tOq�Qu�	�u�s��xr^ۭ����^:�K=�<��J:�ŏj>xD���4aS�뜧�$Q�ְ�u�����U^�����3{cw��{*��OC&V��i�7�)��h�j(S�4K��j���޳�FJ�{lWtԴRQ-�c��{�:1��P�s&��H+�T��Ӻui���f�}�U�f�^t
�`SWkٷ�C�.͕�W���/$�6[��]>���H�S��c'rs��i�,J|:t���h�r���ۮ;E���g���p/lb׍�:�	��P�:6�wy�/1� -!�]k�=����4��I����_;r���ɥ�7R����wogf�І�+LuZ�}7�X4��&�oU������l����G��?{�zY}-:ß
�|�9����V�د��d�si�H�_Fz��'nW�pw�kcC{�"pu[�^;ʍ@P+G������V���h;�ݤwr{���v�y�fbf�)��k��n͸�qg�V�@�֨�p�����K��e�XJ�P���=D(�-��ng�t�R����5�2L���N�����E�hQ�|��9�g�'�$��h����+�݊e�B��'*�u&����"���@�{��9-K��KOl�|��r�H�-�+s:��k�����Ew#�|!���:�x��w�a+~U,Y��L����[�n�s��1���6],)��=�~�?o]��:��x����z�nk>�Q*��|�B� �����ͅrwBr�+o������ˣ#��t��;d�F���e>�B���*�������%��]���QS<R ���B=����z!��W�s��X�\,
�_nz�_��<Z�qguN8J"Aܾ�7h'b�hb2�N���U��+�}��5ZEV_t᝻F�e!Yy�76���7P���������Ρ�u�'P�n�dy������n��J�s�vjpt{,m�ƗP�/zoB>�R��r�$�[��W6r�v2NV+]Ǵb[[t7%m��X�^�uH���)2∋M�g�UXUɌ,N���+�� ��]��V�d��AQH�]�q׮���X�v�:�;9���A-���k~�Lt��8�e����w��n�z!Cˬ���T��zIT��ǲ�YL�)/��>�	��A�����W�y���!B���D2������co�c�|�L�@E�33�����=����l����nJy_.�~���s���w>ڃ�����Gq��μY�|#�>��ygp��z!���d��mۦ�A;y��ݷ�q�y*'��%\wH��o�U�AJ���r��`��3��ʳ�$h뽩D=������ɥ�g��A��|��E�v(����wn�$�hHN���|�Y�2t���թ���Bu�w��^AS��׎m��8�7�SC�����.���E@��SI���iu��l�O�/p��'-��GMk�|��^S�3t�xF���!N�����<};��XtO���׋��!�]�wQ�]�=���7Z��x	�ꢄt0e@C��U��<7O'�g<���"�B�Y�{E���RFr���d�TVu��x3i�7���8��Jpo*�*#�m]=
�g7���Xr:!�o�T���d��x��xdn������+z��ʩ��5�%}�$dL��n���ۚc�)�?n^�P�-��o�G�t�Bw>d��KH����*d��L�J�wc��M��9٪d���.H ���>��^.-��O*�v��`��`>����`��ܱ�����:z/��[�W9�G�RZ����]dR�Ί�)l�e�A�8!o�Ľt]°>����0ơ��7x�1Z����4���=��y�=ꞹ}��F��f���X�$6E�;Z�[���/o0�ֺ��S�՜z[�(E�R̭�I�o��̙U�l�DkIY?l��Ȅm��o��t����3�5^��,�X|�^��=���?���'E��t��p���=�^��I�U�w���7��f����;;�~3��N�<r���TCby.��|���X<=ގ���hf�\;-C7%v�7|k���82�.����n��<UŅ�t�Kbnoz�]�����s6�3%=���qo�tiaZ���0��\�WY�hG�TP,�N�]ꎚ�9zIV�P���x��.���(���|n>���*x-�UR잽r�+�t���j�=��(����H��=��cz��o%�+_wNAX������ouR-���o���k�U��75J�yMD+�d��}�1�ɥn\rU���}�8=Jޅ2|����{�y��5i��o9#�'�1)�6�������廧��[�n�{޷�빛D>C����]���tC�]cH��R�w7|0H���ib�;��+wm�T�-2R�m��TU���)]�6YCy�Z-7�Pە}I�Q��QO�;ǝˊq}h���9ص��v!����-j�
�tiGG��<1�;���_Z���t�b;A� �]w][��a:�+8v��Dp�Ż}���I��]�ad)�޾���:�0�ج=�͞8��s�]�d�`���[��qe=Kw%�5Rz��t�ܔ0�X�B��x]�R;LN'_0ŸRG*ڮ���\���tj��eQ�ݣ�� ��{�{hH7ڱ�͞�5h�QK����b�g�^3��	3I�i��V+9���%�u�^	܁�I�3�
�W�M̾�t���	��Rs8��w#p�K�٦̉u�J�w-DL��#y���㎰�鷪쁐�BC{v���{�%Ec�E`����t2��Mk������S�I�{���t�YRu�-a�%�0I�Dߖ��,�;�o��9���[���e}x��Ap��gA�MҮ�-�	q��8��u]lg�;4t�5Cw���=�˛D���l9M��&A�T��,�����+76��'�Õ���Va�;�:�I�J]tToU�Uݮ[���n�n��'����{����'��Cޒ3�����w �Rڬ�1K#�{�^<�Բ�:� ���4�7�繡�we٬����J%E���vOY#�v���er��z�4�S�ɚ/Us�\��dd�2.&q�G[ݺ	�ͬ�Ѣ�"o�r<'p[��cu��^��z���y:4��d5�ݞ���uؐ)1�]�Yϔ�l����h���r�l��B~z3����=S��.�&����KV�94u�MI������˃N%�k�3}�g���68<K���ͺog��=r�9	j�q�$��
�ѣaO^�}-]��r��w���<�������٤Ɋ�˭��Y���NSb��H�Z��}4�6
� �v�p�9�s�D��{����M�M�	vh~ћV��dj���Hb'9�K�x6�.ꪂ��ݻu+;�S�~��a�΂�fTm�0�d�;H�_��-a��:"У�̙]�O�����㝪��9�Fx
�jͶu��<p�;{S���?o�\�J��ޯK4Ro�������P�Nq�����/6_v:�*�T�E�r	O�[��4�i�ic�Փ*��;��8��{��J���9�J��}S�����ܹ�V�d���uK�Z�dJ�;��
ޣ���ӆ%��C/,��5{*T�]Q����-w?dppg���m��M�WF�Z��F޽X�۾�-l��7؟E�m��Րv�n�'�(�
�0T��� {G��	�����~�SW	�Q�D��yQ��q�Y������VjDR��$kd��թ�ޢӱԝM�n�h	\�ڬ�m��O^� b���L��̀s�Gid��*���m�e�
<�����)�܈�u�l��u�U�0�xGB=�u<���#��,秧4�'M/�u�.'��nN���es&�7EF�o:���w��伃2g"C��=i�j�6A:U�O�Ժ�+_{���))d�=��
7lj��I�֜^E�kq��o�b�+�l+�a{E�����,��n%��$n�0͎ϙ��<r�6��x��;E QV�ʊe�wa����.�I�uH����e87bXF��Ւ�ȕl�[�Y+j(b��n�;���I�.��ꚪ3�T���Hۋ/zN2�;Ђyu^�p�j�{���p��m�QvM�s�|��ى��������2��DsXA�3�ҊS0-�|��l+m�=��?Q�Ԗ]f�Y%�vZ���-_�KZ��M���;��0����A�Z���9{ٲ�.��/+f���!��~+f��}�r�*ح��_Q\ԛ��Wh����!��u�LU��4R����(���>�w�ĸS���+U��jPh������R��jďuxǭ���s��Y�WC�r��T�~[W���݁Lz�yvj+�m~%�K͙ȏL+cw:WE�� �=UP��,p����*��Evg��$��N���z�[>W�ݺ��Gװ#��uw3sv��'m|Į����a�U.�>T0�k/�@�okO=A�ϱ4�,\i[Ό��4*�{-�xs��l<QA�\��!����yEvPj��A�:}@�7flkW�vW��=���\�@%MᏫ4�l��xby�](X���z�o���|����r������߶��5
�v����G�_���=�|����/|!|\J�n�Ag��|y�-�c���|6�聣��<�=�0_:�t$t�K7��	ڔN�������x��OB�U�:vDz��Nr�C�;�9�md�yC�M�Y�_E���8OQ�̠n`I`�w��G[L0���h(�7V���dĕ���MOZ�#�����|De�sƦ�w�xn�5q��Zݲy�c��v�Ȉ��u��k҆`�.�l�P��)���w�al�;3��L��rwyb*��DQ����v[/���&q'A*]v?�N��4�αd�
e��|0Mʽ�����$�q��p��o^���,�A���3]8�ݼ�w�S8��U�V���u���$NE�$q�
�舷o��M�����g��i'k��ʧ��l��t����2���+�n��P���^�۵�uCM���4*��i!�NJ��q�`�9���`��T��5��kS���'Ҡx���_4U3��B#S�Y��jV�h����e2���4ӵ�X���9�c��
�gc��,�J��[���9�V��QTX��5ֳ�;� V�y�M]��+P��k˵#E6�qow]1K��3Nd7�/�b��+
;����*vhWlNF�}�+��nC<�~����WAMY���"Ԧ��?4��|O���*���	S�r��̭��9��]A��Xk��QJJQ�]�k��5N̜���Ŏ�ly2i���mwE"�Tw�s6������#��ۻ�d �3AV��'�o�i��]�y;���sjr�(�Oe3��;޻�q�uX���\�ް�]��n��xC�yb�pcm�Kf�ҋbʚ~C���mM^	����=ԙ�{:�!9(O;�CsMl�H����q�d�kw�;���YP��JFtn]*�A�Y3��7$�*��Q�٩��;�;h���3B��j�W46��=6���(�x�+��[yv�0�vw$o�D EE ?N_W'��ʧNp�W�ۊ3��%��[�o�Ȕ!F��%�d]�K���X��\�,���Ygq�&i���]���z����.H��)k�A#pZM��cj�n�32tԹ�o7X0��o#���H�k��P��9Q��Lc�ב��q�Q���c����~�Խ��
O!|<om��7�>@���*վK;e��	z#�O8J���pa�����5.E$:��AF��RM�9f7Q�X�����<F�]T�3�G:n��@TF3%���@���L�bH)"7�Ɯ�C�w	]�2G$ʔ�DE$`� 4�-$j���H*>T�TQUn��I���"D)�O�[!� ��ɻ-S$9#Ě�D&�0��Bam�R'.��D&)�D(�14!	F�:dFQI�����Ȇ&�.�WlIb��F	BS>��	�&/�P$�FMvĲ��
M2�H'
�"�JBM�n,�[6�!��� ti��?�\t,6A�����"�L�]�%��F,vU�t�Ķ׫����0h�rB�v��!�kn�[H�(6�!��A"��%	dT�P��UO�pB�a,�th�e�l1SE(�7O�
�L6ST�Q��(��1�N��&�0��k�d�$�I@�D�,��h��*��Um;!��"D�!B��T`���fG �n�IH�:�)$S�8Y"		Ln��-AH���)�����#
�bD�������.��t� E��Z�v6�!>�?se�巖s��[����/���xDRŧkaZZ���O^^w�����Ev�O�2��wT;�5������/듚h�5��ZІ���ue��e��)�糫{1>ߋ��q����QR��Ү��X�k����8��������K�� Ӯ��ߺ�Y�ǲ& cZ*�9Fs�Y��C�x�$<��CG�kgW��wxp.�Ů��=�;�}�}��L��p=�����}��L�h��R��;JJ#[f�[�r�{{Ӳ�خS�����V+�0]M�޲�*J/aS�߀O��X�]��W޳x��:b��e�ڰ�r�2C�g>��n3�41:��;�Y3��M���kJ���1˨ǆ�q}(���}�lW	�̗�:0E����E��[�PO=�:|�ם�1Eޞ�g�n� iJ�Q��xJ�i�i5:�~�{���������&���'#,+�0�Nz�
�{��:s��M���/*��\l�nN�kc���hv-}g#�4A�"�΂���EF��Nќ�O�b�[��L;�R"��sd��-�̣3����]xd�>~���*>gb�`�����p��9�,ɑQ��pj�rF��0N�wټV�/�s�z����]�3��C���Yw}�X��	�`����R�+ˮ��[7���y�7�W\�N�v�ރD1 � � �AA!AD � � �A �4A �rὸ��J�v!�v����%�Qk��^ܡ����<veƻ٩5FP'w�6#���+�1F�aiD4.넧�)I�8���zT\��j��n�!3W�ҳi�����~�-�L�3_og��H�L�,�zG"<��/=��W�x�p��G�-NR��2oY��R�o�wKmZꎶ�e�َ�
S*�:Ea�����z�-2��k�|��7��60�X��}�c����l����f[��_>�OPqݛ1g��j�_���u�v݇�N�v]�Fw��0��,���JQ4�L[x��ު�E��S.p�8��ƪ�C1�������!i�>O���vL'��&9Tc{�O��ű	1�d��=��m�5�7��i�b��X�ـ|��}���8���I�ۥ�EOF3�{$X��+djl��v=�FU��k�E��q,��0^�k�-"Y�oF�T/i�̸s�l:�zޕ�
�����z���f�'���[ >-����1S� =�-8/��R��'Β퍄+Q���r��8�x�� t�^v�vQ-�;76ef�`�UL�_8�vꁌv��$}��'�ݙ�%w��ڇ1ó�[������;OL��nk���(i���Z>�CV��,���M����$з���h=��s~�x:��fA�Mꭨ�0`��� ��AA � ���@AA � ��AAA�,:���9�sV����pd�Swq|NW�//U��֓p�b���y�Ho�2�ɑr��aj-��Iy�71��έs�ᔸ��1��-�	<:x�RǑm�/��>�w����s^��{s�ޛ�_��7��[���!�Ҽ�7;j����N�{|�0E.�f{�qxZ���P���P�늷���ޘ0\Ձak$��Pu%���T{9�m����)b��#�5�g5�M�]v��n3�^�9��|�3:�S�Qܛ\�E��Ԏ۽��v+l����YJJ9γCn�M��իWPu�*�Nb��0>s���
~�+���/x��R\R6JY}��#e�E'<����8�K��4?�jdq�����#�������߬pp�d����6f�x�:����S]b���2�k�Ԡ�d�>�p�Y��P;r闫���RӸ��RM{��g�����Zv��m����k�9ޮeZ7�݈u]<y�20�3�B�Ӣ�{Y��~e��0��J�f�<鮭>\Tѱ�T��̽ˇX˔rE�,t\:��߹?=SG�{"齝���8��o�c��bQ�����5j^>�w؋��ѻ�Azd�$��-�7�*����0>��V�1xH����	�ۯ*��5d�����:���g�,q=���7��f����V�=�c���œ{R�K�ڽ�p��A@ � ��AA ��� " � B(AA1 B)J�B�}l�F��|>��#��-s��Dkع�}ϫ��w'���\&!�%z+/�.a���0t��`�9Ni]�D΀�V:��-��}1U��,^�*t��>,{��:�T;+S}���X`hX��}(�u���;�c�w���ԴՕ�Ȝ�mW�_�]� �ٛT�r36UYS���U�ۚ��aGwک���71G%Q�Z	����C.�ϸ�ج�@���cv��-��}Ӝ�ٍcyF�/C���)��"[c��ĸk}��_;��䓆�\��V�\0n�\
��V��rF�F�^gC]��aK$��h��W��ܤ,����F��Y�V{\p��n4�=����݈8s�8�_:{��7ˈ�����s�jIW�28�;����8�����4���Re꽟]�M��v{�״a��w��ə�I���nؼqd=˙/�J9����-��O�w��u���׊d�k�?i�5�D�gf1�\�xX�P����p����컣�^4�T��c���"`D��o����N���k[�_�'���S�e��K��u�=Uoۯ����r�"�ց F:�#�5�8,T��6��K
���:^X��L`�j�]*��M��-S7��\
�_p8�?�(�N�7�o��c���4����NM�5MۗثO�u��.��Ԝ<��YHL9q� C�A � � � AA� � �Ab �8A�q̇�;)�n���D�g�<S!�&-�g�t�󍫮��/���L����4���;	�Lx��2߻=���"G56�9qa�4�����s܎x�	O��}�r�Κ��x'����oC��.�͵��+��}N�0K��Mp�!Y��\��U�u׻U��99O5�;{��=N�qSw���x��}p�������w
�+љ�a��H>��GA��Yynh�i'���R��#:o����/��s�w�vf�;΋}r��/����.�F �;W�#��7����Ò��uf�ոxu��N��tY�"������k��u<4u^eq;҈�L�s	޹\\h��hcb�@��ܦ/�eB��R��긴�/�}}�aڽj�3T��Rk{��=3$޵ч]F�9�d��X��Hp��� ѧeSkSu��qL�}�~��m�ttc��Inke���x���	��Y��΃�����9-�ب��g3>W���r�n�|jou�g7���7s�(y^ᢛ�l�������w��<�rB5�J;�7��g���Cuq��gH��ܚ���5|�g�y��k�x��z�diͦ:»�,I^��'�[��
q�5;�!����;�I������D�y�]�偎PK0G����ix�`nB(1a�CCAh� �Ab �8A �� � �DA �0AA� ���|$�%�x.�V:.o	4b��sѝӷ[hoQ˸��������Ǉ{�gDg9y�r	�g+�g?\�ci?/.jS�=�U����0ۂű%�uݲ�4�Z17p�T��ҜE��ځ�UVSB�o$��{����%~Mͅ���T���75�����|��
����J��P/v��K�xu^G����]N�d��V���v����(1Vh���9[5��Iu��*gr��8�[�u�������dQ#*-�;1O���Yj:˗G������,X�s�+o
��_u���S�{�f�.&oQ��O��r���w�8VQO��x�g.
�̠h,cG�����E�w9���񻕼��۝��P�U�#0nGt(U���p�	z�m'OY�ŏ7�վ�[��U���Yn�w,�_pI�����U���w�;S�PN���l�(�]�'c�c֟qZo��1�k��-dҲO�F��wH�+�+x����,��oop>F�>�2��acS�g�(Tˬf�s�������Z�b^�=&ĕ������H9��4���6���xSF�����e�%��+,�xr��/�.S��|��ЬV�->�͕�ޟ�s�T�v�
�U,�2*��f�+O�����w�+�	}�1.9���wP�fi�Z�6����w����E����p�AA� �A �4A ��AA �AA� �@.�ǫ���Ť��s�=H��7�+�ȑ.Aw��}�ٸ	�T�u�k�W���+�K��w&��y{48hKW���Jĸ�ot�����ܕ{���p�A�|1#cn�H㪇9��s>���}���̮��_iL�Κ�عji�o/Bo!�k���Ϸ�'x��B\(q����h36Tٶb�&��e�؇�;���o7Ս���,���v�[2Ql2:�����p�[��XHƋ�(]�|�s����;q�y�e,�mɪ��ٞ#<�氮�lή�������+���c�K'��k���c�gxvU�/]/é�<�%1�V�}��9��]â�7Bf�`5#��@�������F�ۺ����l��u��wlwv�;�7�F��G)�̅�JA#�'�eS��Ą�ܭf�c	�)v�K��wYn��N֢��n.���]9̀sx���$���+�V���Xٯ7�[�v��{;b��h��V���O��[ږ���v��$��"}�܇1V��]A�ԫ�ݳ�;x�\�垠�qEk�b�k�WP�����Gl�-�i?�<Y%#*#������`6 1�odUc0����(�4��6]��r�d��S����k�hYt<2��w�nςS�t{*�BA�c~U����hi�.�Ç�ӟ}�Vɋ�ݯjAi�����2��c�A@�A �0AAb�(AA!AA �A��Pǂ�^Q�̪���<-;@����ܮ�s�w�݄���ɔ��U��{#����w��c��4�$؅}ۑQ��N!��Mcf�\_-Bž�\��%�խ�tÆ}T�!5�����D�^؇'ommt�C/�0�z�x���Ro;sBg�vj��;=�푵v��u��{�U����xzw�@kpx]��=��y^VXP�[E�>₦j�3���I��dr�4��t���W��
'`y�D�H��-�]�9;�j�n$w����f��s�xv�U��f���gS���us���,��ϥ�ǻ*��w���B��c�1��F�J�ot��=ⴽ��E�+u����LR�� ݻ[n��YNT8Y���(�\���a{���{���i����W�+:�X�_{���/�n�f�om��.�h3�aIe��m����"��ґ������=��u���D�m���+���|κZ�'6�fN�vgv[���z��_12d]�1.v�I�+p�^��I���5Yl�K��x�m!�vF�,�[˺[��λA���ʯ��&�e䮾 -�� �gu�x#��x��"��f�K�����K���Fxne�x�΍�Yvj:I�h~
X�!N�/�ϙ��>q7r���I���:��u��R��T�����q����e,C`�h�w�YW��]}S�sNUnӮt���C[g�(A� � ���AA� �Abŋ � ���AAAB aޥ�c�5ɚƍ���RN��nU�
"��(�ܣ�
�/,v-��r�)�At^2�1���f(��ge� �ꋳk�u}��;ndX��	��� �Z\9�\koQ����ˉ��X��P=�@J����ʃ��s!��l��싚��t w�^e�=����z��tJ��E0��P��#��_;�����t�=V��wp%���roǪN\�g3�zn�(��l+�̮�����y�3�-�8l�,=2�[��-�)�_W�3RLNW*����p�W6�PS��|A�D��W�Ucjû鎑�,�ld����Ut�jZ��9����	��Y�:��
\*��1��r��z!(�ShR�r�WI<ȉ�3i;9c�\Nt�WOu�a�95���ʥ�; ��q�z�+��Q�w�$,�Se�b,}��1��eVl��N�e�;a��]�N�s�7h+ l\����ٽ���mz����Ӡ���eʽ6����A����F@�#ԯ������^����n���ɗ}�K�a��HG/=>�����hk�W\����b~<��R����	�>�� �Z����:p2q]J�������l�t�M��(R����]rZ��U����bUY�5�����s6oM�M�~L�:̟���̫�u�΍���VS�`���Hcveaz��f$Y3�����X�ieꫩ�����w�ڪ��t?��� �h�Y����C�M���&�Jnh-f5y]ڊ�R�a��f��=��w�b4MJg�X9�ub�7��G=n,���;z�Դ6�s쭕��Y[1�*ge�BHj����޴m�`��f�_*��d�l�MoK�8�4�OveWڟJ�1�d\:�Z����ʥ��c�������t�;�ުY��)+3��<�U��r���$����D{��Vq<$\��P��Vp�m�w|���*19��U̺|;f� �o}Q�^��g"�x�~}�F��N����5,ަi������ZR�͡�M�M�4��N��75e�m�3|���7L]�>��� �鼽oN�m+ѡ�¥4�6���Y��5�qS�NG9�:��(�^Li {�Qe�,~q<�$���mw�ʃ�L��d��"S�l�шs��}��y׆��c�}'�VѓI�(R��{bj��]_#�l��/^w��f�#%WbAژ�g��ػ>��L�)���LJ�(t0��FƖ��+���,���<M��:�[����T�q��R;���^��qIA��F�1�z3��Ѻ�p6	 ���P���=�m;O"�����:I�)�z�v����|��;�������»���������&k��R	r�i4��A�N���?����r��7�U��v��A��s��Q��W������i�v���bf%�8�sQ7��P�j2���uR�U1�h�]b*��U�����]��]&�9zR�z�9%�h�w��������W=/�����l�F9yឮ/F���U���u�/�oxhYپ����n�\vL�-�����g}��קn�#+c��#���r-�۲;7y���1Z�Z���b��o��U��p��f
4F�F��c�yY�Wي��gPT�=uSd<���n���r�ڲx�C��ʛ�W5%1nc��{,�N��{�Y��(��ZDWΜ�݊�zP,bc[rx���Ǟ�=���7�Ї�J���ow�~;����R�q����\k.�a�b8�@u&:���vw�����F\��ldWr�����G����Z`��32]
 ��m��TM�8'pY�E=�8�3�9�ݴ��TN��������������������^��|-�7\����fPue�}��<�./,f#ro��f���`ޞvz�$,��y��cc�����|'�$u8~5��õ�\�f;T��6�w���5wx���]pgl��G��b��/r	���1t-o*�Z�{�d��qn����Ww�j�-�`�J4�����L!Fɍ�K�E����@��+�0A��.6"a��h£�BCM��%�>o�>m|�����EAEEE;Y�LQ5�PűX*�X֘�*�mQAF�[D���NX��QAm�65��c�#�A�����UE�4UTDU�bY�=�|>�ON<(#��UM�#T���ch)�+cE�h�V4[gmTQ�1UÇ9�ƹ�*�<(��6�H#Z(�jb�*�<�|���EÉ���O�>���9r�EUc&��Z�h���*�F*�a���J�cU�Ç<����j�0UPUA��m4�>N �<�V����W���Q�/y�OOOO^^�i�(�&(��f�׊�S��o(��)��E���6��/�>>_̞+�I��Z��xyT���i��ӧO^}�}�I����C�Sd熯-���bڜTӋ7�7��2���c��Ȗ �@yC�m�U:e[g�lyo��N�8����e�<�cv��D&�o/<���)�m��u�&��xy���E�����X|���y>U	��hյF�mQy�y��3�����h����m��	�(Ӝ&i��
?+�|�L-�~�U���K�g�z�!m�WN�Rܖ�n�Nf��г["�'d��`��.ڠ�������m���u�g�E�a�#,4a�#f(Y(@�~�۝�׳�����X����8���L�&�#�Opm���?M=�r�yB��+��[{�����2��������A��L�m�I�gn�v�\K��ޚ�%�K�L�12z'ȭ�7~�"+xQ��9���|8� �mg��ު�n����8���/�m�7�_�8��5�,>��I���p�u��V��,Ēc ���)xt��;�$lA��3o�}4��:M^e���h#g���$l8��L�X)X�
��w��Z�ݫ�r��D�d��^%�� WQ��)�����]��Pf��->�z�5Kލ��-����LE�'����]�����%k/|7<pT1勇�o���A�f�PF����.,�����z3̋t-�m,����yS�m�@f��Â�=4�Am�<ÿyh�x��y�㍺��CF�V��UG�{��z���v�r���vD��y�����.[2���]�NYñ*K�y��)���q̌�֛���<
)�k{��a
j�4�\L��T"���0o'q�^�xk��Ly��A�3B���zwN�-����bQf㋒ѿhn���+�xx&|��Ģ��k�<ﻅh�
��7ւ,�&�cS����a��'h����DǇ�o�6����,Gw#�¼ǳ)�5�����A���A����Clp���Q�8<5�T�c:,x��jm��0���9�3,��=��"}���O�.��&q���{S���ݹes���R��)���L��d=�t���q�i�q����e���9Ś����OC�S�'rb7x��{��IڳZ!��'-����xpv�Hi�'�� �K�Y�ᗃ;��xZj���S��s��x���L��/�R�qܞ�l����j���Sa�w���6b�z�p��~�o^h�FH����~�.������M�Ol�����8�$a�y�����/fh�5�aG-�Y�4K�O�l������N��9r#õ#U��u���wZ�ے��R��KFflӖi�[}6����yx�0,oO-���=�Լ2xt�N\�B�,�R:Q.��,�^���wG��i��+�p �mgU>�r��L�Ě`�p.Ǵk�<��"�%fĻ"�n[���R�ڞz/'y����W�<ؗ7�/L���sGܲw���*�A��j�{�>X<z^{�z_پ^>�l��)������� ~�ap�w�O
%
�����kc�o�@m�{¾#0���Tc��ɗ�凵mk�a���a�w��z���g����&Ȣ0
�'��v�R,
v��PtD����	����k�9�Ib��9���1ʜ�Mrh�T�����h����^ư�6w�x�4"��`��>~���,9*�1��]�c��׷�jcڎ�X$06_��=���$;��	�0{��?Ji����54�z��k��k�t�9,�@[�Q�5;W�d����lϩ�Ϲ�Ͼ��J��������z��g?w�a\=�vҝ����鼵�g�1 �qfN�V�՝�M�'
���=�p�c���dթ�d����Z����=0`�,%��������?\z�r�K��z�͞꧎���t���c�Vot�WN%�����9wa�wRރ� �='��ҹ�6i�s�j�]�Eʩ�ތ{�|�����>��ᢼ=���}�lq�y��Oc�V�}�b�̳�+sxqd{�����Y�.z��]<�7z���^,�Y#����ݒGӬ-�3�	� F���u����=F��P}�ۧ8��v#/�z*k6�,��>������3�FV���'��-��t$�v��^��}6��b��w@�i����>�>��=������]���/�WU�^Ԃ�߇��ǡ��N��ϼ<�˃=6g�o��rx�>6r�a���QsS<[_����I�������m�ִP󿁃�ļ������yfz�fj^���̡�, vȼ�O]�!���v(k���VmZ�~�.Q��6�o��l�.'�B��l�������Cl{|�3���\ǀv��Gf������,��\uea����9"����D��ϥ�pH��;ßkri�n��t��Ի����S����rxU��s�ٜ��G�ٱ�Ɗ��q��������q���kǱ��4���.���+A�[V.�J�BT	�YC!t���wh~ŻqLGk75?XĪ��r}�Jj��R�Q��Wb�
�M0"�B����<��� �a���]X�%��w^�b{��A[]3�d�:��I�>��<4F_ާ�.yw^�5�#Lϕ��ht��=���H!ݬ�c�r�Y�0[���GLh#����b$��A������D]�{�XP���	`t�R���K���݋�������՞�z}��M����x��o[j������1�gg*�+8���A�o��=B:O{�ћsB��ҜU7������}��'t �p3,������i$��1�kv>[�m����;Η�JFj�aR�G_���b�"}s�=�v�i���W{�S�����Z�����b+�w-�@��8�O�ċ�z�p��݂Om�,A�dȜ$���i���vv�ں%��<>����$~�'ް� v���Got�T=Ij;�Fd�9�=��i���l�:�C}�]-���@�~�^>w�6L�`�`I	X��(�8ޱ��[�\��쳓_\�n���R�좆�:�GbKxt�豶�j�{Q��)�CFKU���W���bٷv��F�N�<�Q'�%I�d5i�G��6d������:1T�&`��ubs���	,�P�O#�|�ON�Ǯ�T��=����՞��{L�R(�JA?^X����L�&�D��3E��^�ݓ{ t��s�;b�h4j73���w��z�^�jɾFr�����m�����U}[�ໜ�^{1��F�,ʞ_P��^X/Ys�y �ޚ<^'��_]��4����vW�ͫ���`bQzQ��u�%á�.��ڤ�x,�#$�:����;j8�����Ho�g���x[�o6{i��s��A;[�?�~�n��VM��]���%�a�A� �.
c[���:�f^ۗRͮ�_k)-7�q{�ݏ���g��^������5Ҩ�V1ù��}Yg����^_ǻ&�[�]~~�Qx �=<�;W��C|�WOo�E�JoV��C����ϻ�k.ۃ��C�������I�Vk$9v"����̧*l>9��y+"�d�Er��/��t<��~}�䷬�͟i;{�>�;�SU��Ƌ��޻yw@�G#���Yb> �;Kr��J�� �3}�-
�}zy۝����hGi��vמ>�\ؙ����]�x_�xh�,�}�oR��{`�/�A�����hn��R�vؘ+�S^��=F�d�6�X��5mb\�r ���/UmF��D���*ă�'��8��Mxa&I������Z�̌�X�Ά�m�<t����j'�M���#A�7h�W=7�^�xKo�&�I�+�n�Ll��2jT��}@W�ʬ���`\5I5�^Y��^�g��t���=Aǹ��g����{�j 0���~�s�2H��Ǒz_y��Ygֲ����{<2��u-�W�{A�#�e����Zwm=Ю�r/l�U�{�Q���&ތ�/�ං����dAN���YF����^�)���sΎ�;���B��ǏE�`E�ئ��0Q����k��>wY�p��rٻ����M{�G��ʋ����Гk4�����ռ����z�n7Q�o�e�zu�ѫ>�8u$+�a}[[��s��*-�����m�T�0����T�����r�]��c�����'���պ�z�ѹ�W�$�lt�ѯ���p�:fA�\t(��=�Ơ�RZ��R�G��8�:�B�x-�}�E_zo�P�a��$�1ʗ����Wy.;�p�~�/o#��6�؍���e�����M$Gv���0Ow�^��&��W��yS��G�����Ձޗ�e�]�5��3q��d�2j��T?	c16/'^4jN���E��{����H_�����d��?�7]�6���ν�WG�� ɸ2N�@��w.R�@� xz��.�O�踆���^��=wĵm�.t�{ݐ�A�/���OP~����@^�d� ǩ�]����X�=d�`�X�:4��"n��q��|αR���$��y�K�q��bu�AD�A���x�{����z��$Iܲ]d��"n}��ã/��a\=�*!��Y�o�nw���uP�b<��hzWKŻ��::Xx�S�t4�yA�ɦ�]��&F��庫`	�h͢�w'�б�C*K��ky�
6v�ȸKo�;;J�����yݟ��Չ/��=[Ît�	�'K�{�\����Ԑ%$	%Y��38��jݨ5S��%�w�����t�PJm�c���V��r�����w���V=1����c����?`�`�	���@��� �K���������1Pws���R�cx�O�c�v}��Z�u�.��Zȕd��B��jy�Ǽ�l�v�A�n�~��/�ñ/�P/�G�*�m#��iN}�<���X*e����\M]�螓v��,P��h6���te��n�[fw	����O��,kޛ��?Q�\��ѯxT_FM� �u��v�}}�DV�Y��,0N�������d�J��'*�=8B�μ�~�]$1��?���ht������jB7aa�Ͻ�����H}g�Hπ^^�x[���p�	6�x%g��������9���.�^>�x'��= �Y�w��Q�[��D��g� A�y��}�ۘ�⬂ي����s �;]�u��kNl���"��],�ۗ=�5�ﯣ'�%���=��᪌����I3�}&���y3Y]Ӗ��j��0ɲ��˷Y���#�y
(�⼅�:+�Ś[�C��;2���D~���Iu^�@=A�X��!�>80���2�DK아%�ل\"��hī�>ġ6,RoX�&'Oi���5���(W��)}��w{�t�-G�w5{1������7�D1��,,��6�ι�97w��Mn�SQ�};���S�Y��Ș�[8�N	"߁�����;��uyf�#�uĽ���Ƚ�3�I:&_�1��������#�����e�8y���{®<7�����_��O=��O$ɂ��7��\�Y�"n�$������^1�_OP�湁v�o���I愲�tZ��ch�oQ�z��{���C%���/��L�(�d���f�{�6�E3˹�3��O>ֹ%�*�зC�9t=�On�زo��.,�G��m�OVk�{�Z���vKV'�Է�6+��!т��O���s� �ކ���d���]n^ߥTi��;X'��	0WX��L������M��OVmjX�F��ŸG!Ŏ��=#h7@�gs��xH�� ����j�6"]����(�o�X:<�\�������l�;�����ֵVT���א�۩w�����c[�P߻��A���h�ls*��&�QN�e�JT�,2�;[����Ջ5qھ�Ryww��S9�r`�]�0���SI�'�~,��t���,�krfNc��ypڕ�	%>�-���Ehܽ}upzԪ�/t��ں5��l::��i\1xV(�� �2�|{e��+�����}Dl)�)Z�鎋���j*�s
YZ���z�4�I��lfk%�� ���s�8ulw&H�s�U޽n�$��ݷ�L2�I���JD�v�x�1V��iX���Q��2䲗�f�F�̝Օ�V�P��8�Y�i�B�$U}M�͵.	%�yw��m=q���=���8��n�~�x�n�l���}�uK	�u�q��$���٭3�Sc[��8�Cn�F)�2=ٻ�1{��zaX���#Vz�������y�7+�y�� �w��ҝ9D�7Eo�HwR�)�����ZN�W����h��	��c�XymȍЛ���9�s�Y��qJ���Qz4uёl�&�eAP�s���A�)zv�ا�,~��@y����ǷI�0�J�*o9Wa�q�E�$�I9�Z���kb���;���qɶ¤d�;��f���U2������=�^��Qލ(=ݡ��N��v���᳻~|MQ]!��k�{�V;��}�e�[�(�������ԥ+@$@D�4��4�v���B�����";6��`Z6�}��Y��٩z���4�	Y��y��l�P]Z��[��<��Ӎ1�X�<��Fzz����|�ۧ5��D�}	Ž��Gۙk`�����q�I]��ڨ7�-�Ěm�+_V��{�[)�1�J��c5T�qL�|�ŀ�U�󇈷��٘�s�?{c5wn���,���3��R;W�u��1��0G!v�kyR^�u�U��ǰX��E������Z�=X2fE���Y|��H캼>��L�ܹ{X̔�`��s�Vz�i����N?�����A�8:'���aHt���R4`}�&���;X�"�K�E�D�Cel�.�]�鵠���oy�&�9���w1���.̆\�£U�k\���q����v�wh#�N�7��-�L��0C[�>!���l���;g�J<:`��Q5�f�(MW1Vk;5���=e�.-xZ���[ò���']2;)�jI|/��ߍl<s��]L=�v�N+�Ѳd�DƦeٸw�#�!Ν��=<���+�$���\��{��{�?'�}��m�@��LUPˆZ?\��ܑ֔�,�Y��5v�0�$]�1�gg��\|�����������i���L_	1��	��w�S���t�oV���a�����Nk��+��[�U�յ�s���.?Y��V�ff���G���("�6�E���8���F�yk�W�*���~|4�Q���5y;�4����~��?����q:�;��^Fj�9�l:H�#&����#N��>�8�J咨�� ���o0h*��`���1j������b��lx|===8r
� �m����~��0h�&��4DSPTMQ���ӧ�M4D�EI�qPSCE�����=��TUE5��zzp�T�Q��<|�������b&"*" ��44�x}>���9ILD�EQAUS5MDT�Er0}�5�c����ÉȤ"f���h���w>�T��A��)���(�zzzzp�%PQLEv�Jt鈈���a4U4�S�T�AMLTkTđ	UIA5>˘��cTzA���*���Ͻ��{�y���ʾwv]��\�[Qs*�m��ڸ��L������y�q����*�;9�f�|π���͓�}^��}��z����M3�5P5!�!�� �$�4���9	��W�,�Z<���s�/1��}�X0��F�?�H�b���'rHokp�i�(��
W !�9�9�i�m�"]���O����A�L��R�=3����"�	S��W����~�m�vPc^��NO�m����"M�څ�(���ȹոٴ��V2$����aּ����)�0K%��;��t����m("{�����}&���X���.�Ǳ'��v�oV�^��;ǐPH#����!�.x �U3��EA�����'շ�ΡpK�'��(FQ��/�k�X�g���y�"��''
��k�z�*�y=jv�D�$��?���)�r�	��
d������O�p�dɾ�Sf&��̚���� Yz7%�cF0i�ѣ:Y�G#a�{��$�g�ŨV1�j�W0�Larxۏ�qa���Wze�y�?�C��#�#̄&�<n�^�jO`S���M��2[�r�NW6�_r���.��SX0��/;|���Zc��DA��]��>z#��,C�-z���n�ګ�E��\t����Rgr|$��1&KD�#v�)�g�]��M۔1hه������y��G��������Y�`'�s��h�2��M��Βw�5fq׫RLfŌ��+���	*���EmS�@^Bu�W�뎱�����m園極�c5 <u�Vk#`�i�V�'�� �6�Յ0|5��.��q�щ��ꂏ~v��� �_.�U��Оｌ����<�/2c�f YL22<���k՞x埪��[BǾ��}������Hw��g(Yqj`��/�^��T#�z�g��~ɢ��4+CQ*/P�j�Wu&�����]����$:�=z]��}}�mg5$��s4¸���*(�b)�iXwh�yי�K�:�u�����ZDL,ss0[�0>�{��f��q�o"�x.�;,��[�Cb��[|�Ţ=c�"a�Hq�/0��M��r<]�P��%�l���6��/���.漢CQ0��-�ߕr����P4�0y�����·l��Uϫ�ٵ�\^�^9.��ck�nt���BK��py�1�q�!�F}���ٶX���=;�,'�!'�sLH�U�m>%ִ����Hv��*ڑ���:��A܅�%�z���v?��*.��fta�۪�rn��mͭ}�[!E��2%�����{u���e�c�Ruc�JĪ,5y\[N�\:RzdXfl��?������,��հQ���\�?�'S���̍��°�OP�󣱖+���t�hq�^V��i��,�HF���G�ft�&僵���t�����m�(�S�k�Y�ZT��������z���"[�_t.'���.�m��4g�T�$�J������G�<��1l�8t�m�?����At&	v�{>f�#�KsS�&I��"S���j�QN.� �̶	����D[��UŴ���cz��q0�2�[�5��z�|M*,���8NX+��l%�j{��hm�fZK3�.�@�f�Qa֑��k����#���1��v1
�3�t��ԕ���/QÆ�:����ru�pH��T�6�Msם���C��� �kϡ�n�K�(�n�a�D�g=�_+7xEfY�K	K%s�U���4�*|}_{i��I]�����^�ۡ�Ѻ�u=ժ�|����!���^yҕ"���`E����P��̦�J����O��N�5�d���
���z.�W��k
����6t8��q`d��8���@�%�m	����	�� ���8<��z������#��+�ό`,Njb���P͢Ú�;R�StN>�iܒ��"�6Է�>C�+b�Z`c�W�}�D�1��-�)7����u[�ͳ۔XW����ۇ�Iۍ��t�s7+�@.�c�D̻z� tN1��l��/�/��և�_�S�(����S���{���ݱ�gzk;J��,H99���g����6���-�Y�+��t����kq���S��V^�|JvԻ�j�[ď]N�(�,��7�#���^G.�qVQ��"���[ǀ(/6u��ȟ_)�k!�M�}���^؉�ϟe�� jm�ÒHk����⻤"�Nm�g��(�e^16��8�=�@�����O�~����Uꘚ�o3�k6��,������xl�#��X��A/��{_R�C����*gݮ��,��Z���w6@�����p&.��TcR�����w��Ȭ����0�d�~1�;���<�W��̵���z�϶�%�9loX�0�D8�y��J�j[������o#� �Ф����� \U�#V��8l�k:q��cռ55���0)�5y8��Shq7���#�O5t!>M�c�;ʮ�l�<׳3Ә^�{�v��s ���2o����{oc���(L By��խ��������E�����������^%�u�B)��&�������Z_�<��|G߹|�d�k�'|��.�����n��*���y�N�_*�_�tS*����`Ӛv���E���J�m���^O��]��'�����d	'%C��fga��_Y����a��w�l���,vs-<�iw��a�`DskTH�ot<'X:��-@��J�sj;�M�tC�+)��pN�?k~x &k=��Ә�S��zrՊ�3��Nr,TiS�9%�q��Y|��^�����I��Bu�zR��������<��\[�_����2<�at\=4ǅ_S�W��m�wX�<I
��{+qk��ko�ɽ�j��x v5�����x*�����|�p[�(����pȼ��%�vd�2�5�(�˞�������Ģg���5��+���{O�������a�@A��)������ e�i³yO���b���m鎳�+"���-�y6��=�_X��K1/��p��぀������<&+�K�mf�D�Ż�Lb������' 3sr8�Yx���Š�1^tE1n���=�.����j���򖌌�~X,�U�������E)�^�c��A��uki&�$@"A&����[�]�˿��{��^�\��H���r����<7��>K�=ݡ��X�`��4vu����B�IB DEi����C�.����:��L�(S��0����ǔ�r�����rTͶvPc睊��
�n��Z3��Z��!��ݠk���I��t�����:/ Eǧ�J�`��ExU�Fk�+7��F>�;����g�&�h�'�]9��$�XGx�:8��.PW���[���_��qۗ��зŵ�v���hB���NQ�d��3L�Q��q���L�,�(<�4r����s7�+�&J���-�tOڻv��V�u��sI����T?˼E�o^�A��#��\g(����l6���u�=���Q]g6��cBQ�#�h��y����U���أ��B�Lα��$f��n_dͷ4��d �k���NI�vjS�Y8`��A�%:`����V�E2����e��1��>�î喺9�;wk��w�0���[�F)f���7���8&�Yk�yNR�t�T���� � �oϥu}���t�ؼ����d���pC&�f�y�E�S'!7K�(������Iay<��/�Өu?����	�a��s�0�`.C�B�F��f}�;��0�^�k����mI�O���5_�ψ��ćh��(/�4>�g�b��?.��D���`���W5��&��k@ʬk��Kű�oG֧ʢ!���˻6�oR�HA���K��S���������t%ۘ:����f$�^/�_�G�{����-��A�=�	wX��F�����:^B����1�(}lO^�f�E��)`�H	�i�{�`v��j�~姏�澟3f9���&��A �+���h!�d�"�J�7遌����;pЂbK�v���X��i^��Ր���p�R� �Z�CT��[ �|GE�9����!��^�v}2���Գ��
j����q�<��$�ƣ[�9t�o9�ɽo��W��{��U���p�Dt�sGu�5�J#���du���yć���'8�d��{b�&�\�^��ْ�u��2��B�P��ep�Tnew����=��m�k{�u�v�e���N�ra��
4�&+� �Xk�k|=.�El��d-N6��&]��Z���)��E;�1'�� ڴ�X%\�\}^Lq����,ӸD^+e�Q�
��+�J3�P͖~�1�8|"�%�5��ߕm��\a�ܸ�˼���UO,F@�C**�S��[��	���˂��g���C*.ۀ͝6��h�T^-C�X�-X�.:����N��P���A���ܢ��FD�	P[[X�u����4v��+�7�s�&����xS����b~���rs���;)����,��1bi:��P�{b̫�L�!�<�{S���!D��ȦvE��� �4�t��o��e����6�M*�@�Ze��]Ft��l�Uw2֚L�W=q�@���4n/�F����pƸ|���� �`C�M����sl�ќ��7�3'�C!j���QL��� k/B�A���vlg��=� �k�}C{����5a;TfA���=u����������,*�J疳Q�x%�#�$(��dy��6@}�&�|d,��|���1���G7��_`�V0�Ė���G2�)V���c4|�a8~�:����e��Y���=*�fdA�[���#�igD�q�!e�;�e&���.x��3z:"bͬ*�s�-�����jd�+]Z�,4�[���U�]�ÿ�t-+};1=e��[÷�o��|�U{��ջ��{w�rӝ����0�D�]WD�r7���C�- @P�T������^=��/2��%�J�`�Ij�n�)D�ŷ�cp�gj���ú�Y�g��pڟՓ�/d���ڕ �	�u�>�^��@��'Yt_pB��v���ږ.�O���s ȗx �v4:!����"?|���	�Ϩн���;�T�6���#$��R�j�c��}�3>v:��@�r�Þ]�(��>C�|`7Ki��}f�1Z*:Փ�ϲ�����q9��� $?� ��˴��e]i�V�J��Pb�N#�����s��g`(�A�:�Տ�l��l�$<6��#��K$+Ț�[�l1p�G{Nt�15�]��+/�;�'m�|�ଊ5�Qw4�e���hۮ�޳�Fs�t@V��xG�=!�6ۋOThl]V~WpN�X|Lz����L��|�Ɯ%�H�ϟ�F<6�y��M�8�L�g/a�/E�A9���tvл�ס�L-���ڡ� cS�/쩀����أ������x�-a�:nT�m�kj�x�u`�LeH���}��6%=�}`�!��{,B`�4%UU�{��6/c`[WŶ}Yy��
�mɘz��"q�O���g��'��?_������P޷����i�h���T'r2�7WD�vnLy��&�"���j��K�Y�f�ޣ�<���8<.��v�Q�
�+l�{�I�� =������u`��^�L�N�<2`�.x�2H�aߖ��)[_ʶ��Cȝ��������v��h��[�eC	�B_Cy,h�;)C��.�r�E��tz�V.�� l*�5 ���������d��vH��i���GL��`&�Oa�D�q=�*���O~J�a��՗ͱ�}F/0,�%{�@}��<|ɻC��0#[�bS�����;B�	��Q��oofșԦ�gӄ�Av�ñg!���4�{���:9�a����ϫj�Y���a62a���蛬u=�ݧy��%�+���z����]:
�!�/�VGW���_f���a3��}w_}��n����t��ϤTj�ӯ\c�8i��B}C��GӘ%cA0������{��8ˎ�&�<;���P�+I5)������^���$��1^��-���z%ޕO6�zer�4Q�ۭ�C�#��B �K�����@�v��`�C�"��f�Y�z�&l&�.،\�N���%�������Za�z�o�67hkO�s��+�K�,���g�_�dQuc��w�������eFv���D����jw�K
m5y���.eU�U��{�&
5���0P�2D�VVͦ�;��̀�A�G��AO� �ݜ�b�� w���7_2U�=\�h\Y1eH��+"���7���&D�6�E�5i@L�<�]��%�~ miK=~�������g8ـj�Ņ�����Y����NW���S7������\�K���\�i^Fq�j&�����z�=[���x[G�:/��\zz��Y�4��J'*6�s���K��P���D�u�҃&�F|E��Uӌ({�b�Ui�U�ؓ�|�Lu�����s����MZ�����+ѝ\���(�I�$f����i5[Dv>5{gO"�FC�b������٘�Ĭv��X�9�b4}m����> �d�����_+�|1�X�S*�F�z���ͷ������a�ծy�EߖC����E��f�M��#�L8��4�&�I������@�0�(F���0-\���/���n�S�а~;Q�9/g����0�r{��m���F�b9��^�i��U�V�)	:��;��`$�
��e��}k�s�>��Z��n`�d�0�,��.�S����^/�,��0���/��c_��E�xQ�t�B�R4C��:̗O5T����9k���R$S������Rr،y4���S#5�ݛu�1���{��4�Bb�8��Ѻ�� ���m��F���ty�u>�1�2Lݵ����r*I@��{��D��[�V�VuLϯj���_�#��?�7��^+�U� ��쿕��YZǇ���u�������S"��m��u���D���I:���-�/��D�V`�GY��ZY��܁%�um\�ʹ�ګ�j���>����Ѧ�n���4��������ۣ֞��p��S�:N[W�MP9���-
2�wկnc�*����A�b���Aª�TM�
P+m䐳���� �w��V��pxwR��{8��E��і�{�����M�O���Z4c�����b�KnI�k�r,�z1��a�)��Ĩ-���uy"���L�
i^@ f�Rd����1��Z�U4\��Ut�B�w����	..�8kR9�Q=Σǰ���[�<ѡ,f�b�<₄���b�SO:��)��U�l���Y�i}��r�������.�;�%-���6��{Y���GG�Ma��k��Ǉ���N���쪘Ob�2^ �BE>k�l��>;/���y�/�h1��v���eݕ w^z}ڣr;�0��W���*��H��2��D�z�s���7�P7���w�;�ċFG���h�M�̡��I�ơ�]:�����kq�/uh>�0V�̋��5YXw�7'hT��U��i_0rJ"e����	�0�U�S$<���Hz���q�;�J��uT]���9������s��7p��{�d�p1u�Ŕ"�Vӌ=��Z��[�AL%1n���󊻗�	��Y�Ᵹ6��6��13���TG;CN�U�/��:u�2�W%L��a�Yj����M�aG��x
�%gb�	�e<�Vӵ,�ė���#.gmt�ps��6����[��7+�ʧ�L-������f�Px�!�w�Sov��������d�9���l��|7������`�:|�af�vpk������5(Dkfs�J�&�l��Mi��m�d�x� ��iK]_�r<,U	��F�/+i�os����z���q�gI�$��H��.*��B�mt�n���5!܂i�(G����N5�������!��〉ٺ�*v��/q3���H3��э�����p�υ\]���T�˹7V^GSm��m�nNw�U���\{���!ëۗ�c3�\���A��%����5�`���eQ���s��u�
ݝ��ʋogu.-��D��ػn��o�����
�˦6ٷz1F=��9p�1ҡkt�y�i�b����؝� �֫��i/pL���fs�4�ֶL��6DoS����كE���nl�(X�I՛f9Ui�[|e�̒b��#�����������!�,�'
P�Ф�R�`#NG���h_�$�`ƭ(�&��,�
-�F�5�ȒB�Ɗ������@�q��iQj�pG>m�/���~��5T��)�W����U41-MTR�UQ�OO����1��^HbB���24U��T��	Lxxt�Ӈ׎���#���"�$"Jl'��R�T��6("�������MU5G-jZb���IO#R7�-�Ʃ������Ӄʨ~ΚhZh���Ӣ`��b"i
"(�)
�������y%4�4�݊
��`))��N��WA�c�ÇJ}�@RSICKQRbQG�b�)���Z��4�T�y�A�OON	�* ���b�"F�F�������Z
-�IKtKQ@������������$�4�Q�o|ʢ"j$��4�F��Q.�ET�QLM4�gK^ZP����k���S
QLV���<��ϛ���Ƨ�zʯ���WX&��r.����I�d�|1⽋��pB����p�l����<(�юk�s"�*L������c�"�� ��^�s���"Q�����'�z�_{�%��^5���V��c�}����!۲|���T:�q�鵽�?~�aL`U�yP���E�P���-��~Nf�Q#���y��3�(K8�S�zu�8��V��	�������g�V�}01��n�m~�2#I�.�$�~�nY��h��]���xR����`?��Ô����$�|e����:�L[e9����J�W��-|�.{^xOv��҇3�%8�7#��}kO�ʖ����c������Ǉ<��qwTK�3C=^��Z�#6ӆ�#V��0Ppq�nd�dQ�g�fͲ��l��sӿ��K�ԲU5�O6�;!F:��L".-ݹ�k�'�5��ז@�T�V���{lQp�+G;^ʙ�����z=]�)��zE@����q�&$�O�N�g�\�΃+t(�
�jR�J�
e�ʰ�ú>���4U�����)�BnH���������>?����#��oY<0vJnf�L������6x��/x>S����`��Q..�r� P;8ѕ�W��m}�A��O�͘����rǅ���_�`E��Z.���{ңx<���o3:vN�E�{ת�3?L����a�Ƴ3qW��7}�[��$_)�\]�>d�%[��)�B۬RG[r+�\���1�f�߸��K�-�&�P��t����]-9���g��� �g��u��9���"���A?���RYi�7c��x`k��_��Ý�/����	�_����7��-VL�/aRS��d]cع�n��\�����[W�p��t�Zb�U��קwz)@i�@Kκ�hУ`�&r<�Y��O6
�Ƒچø��|}�`��C��s�a� �������]w��0k6I��I`E��e7J��%=��V�����eե�ȢGc�7��A��B�`�J��� �c^�ٸdR�u��Z�T���Z�z���E�Gc�)�7$�B��'ƹXKӘ!p��j�L,�z�d��^�a�]�P�mC�0���Ec����)�b �S������3k��x׹���`�A�"Lp�	���!���a2~�|�����8]�՗�í��6�F�
(�U�h�U{�#=���uX4~U�$��3�3��Rnݩ�ޝ���z^��(�,U�v��Ȳ�^z*<��H:��:M���	�~�4�(��
�g�W�(e�B��q"3$��{Ǧ�^ǲ��ȂC�v9��R&��.����ܒ~_�=�?H�d~�z�!�>�\�����wQr�N��soS�) u�ğ��ϭ�7Π�R����l��}��䀜d:�-j�����r�)�n�=�e���uZ��M�(FA���=w6諦'&v�W7�xҒ�I���| y��z���v�Ӕ-���8���/~��j���E@�~H��eТ��x�k-v(��m�����%�Mv�U����^(��3��k
��?)�q�����DEܑ�87O����	��S�_*���QE����9���4=���gq�'�/����-�6�)s �F6�<;��S؉*����u���b�"ɱ��*����\A�䳙�S,9�Wg����hxgw�B�>�q�,5��B��^%�u�s�2��-,��鿖ZL.Ȧ��rU迾�݂�1Q�5�K�ot�4�T;(��<�L9O�s���U��ۋ�r܍��GW+���Yw�E�-|�c���О>=T���l�(qUeWC�b��$�G�$x��י����|�����cu�����ŵ���v�Iu]RX:rE!WS�S�l�=4J���n�1��C.�O_c`^��a>��|�}��g�d�2�M��:����29�u�e�6�ܹ���K�(8�/t��|n��h�!ts�x.������+�+���?��Z��C�9�<�Fo��v����:e�\Y=���r [c�#�]�۷j���H�g�z�������@�.�F(j7���
��q�A���e�[v������!��cL�}zgs���jA����(�붎wK�9;��� ~ �6���B�3��;܇6��ci���3�ס�9��KK�,3��tg1qֻ�vб/Nwm�ӝ��i�|�[လ��'�.�'�yW���8�zA�ū�C���l1��sT���n���������qG¥9~L�:[�s&�;p�C�OL5�>�$np�\'n޳�0B��]3r�^��!4���Y��'�4^=����6p�4vB`N�a������>�u�]��K��� �_Ӓ
�זR�3p:/���|�1��_8�>X/^��g�Ի�M+��fd�Gp��,؀Fx2X����Gh=ٴ��V�3a� ��Z'�f#K�dzy���d�p푱7��w��`;R��HD��m�2�&�h�'�+�88��C�<T.xh!|�J�ezз_j����
/_x��HP@�t��y��N+ܢY'�$f�X�i��`��W�{gO7���C_	�.��W��ݤT
ǂ�֦9��� ���#�����)ͮ�L�#K��*s��o&*FJ܉<-'�~X�P��9�0?���98E���dq�&Q�E'*^�ߔ���4�^�#oB��em�ˤ�M@fN^�s:�C�O;F����·QRdA��"C�_3�P|�ʻ��B�J�4��⽻ԟ-�\]������1R�ǌM]ܪuʽ�G\R�ۚc\~Y�Cz�W��6��u9r��D����IA�,�� S0��H$7�`��xI��!�I�����<Û9�����{a@ ��"�}�Tpk�{<�^�uL3�3]�i�A�����.�1z��)�./#�#4�I���m���=1�B�ګ��fz�f�9�b�DN⦴5*��)c*F�����W�l?&���
!��k�L.��R�AZ�4��m���l������G���Kʽ"��t�c]�IN[&ލ)��|n���"wQ�4/?B�vO�~þ��k�j
hj�B��<3k�{pе~1%�P/�^��WA�sh/�ԧ:cF	fꌻ��GT�"�'kU�09g�!1i����̟0^����I�LbXqg��p�T��!���͕��[��{��p�:��(��|s�ض��p\_��A���s�Bm}6�����䞖��ܮ#�������}�\\9KOհD�� ��o�k��Q��s1+�ާ�G����Hn�3�^C���`�V�[ ��z#gM|�����D�`I�xE�1���Ys���eSV����e�X�g.���� ũnJV�c8��ӌ����Py�M^������&��i��2U���:�c�V�f�,���D��j�>��<�j@];�q�(!�i �L��� ���P�I��>�\^��oK���4����fl��J�<�$�f�|�
�oz�Hh��'��{���|�>���~wؿ��$��! .z�!)�ġ?��iwl�L0Ud��eE[P�'�vOK K*K�Y��H�Ƶd�zi��U/OpʛWo;Z�|^�������m1%�WN�g�\���A�=�QI��4)F�a�DPP�;�������L4:����)�����SI�E�p��)���$�gs#^����귙L9�k�,�*��[�S�v_���x`k��^�[	�uH����f��FF҆@�U��8LR�)9Q!���>�:]�>;� @A�v!?n�l�jn�����R5�v��ꆞʔ����"�����N��N���
���^���_��ff{'˾ζ�(�@�����a�����*��~�4+l�&G%s�W�ܤ�T1]�O�7w_5�0�L2�ko�k�;��˧�%��k�M��^u�uK���U�9��J��ok��;�/��pv�Vq��|�a�H/�$P<�P-<`@_�צ�O��q�Y~��s�^���lƲ����ƍ~kd�\��_�I��ȏ3!��@@|Naٖe�����3�K����n|S���׼�a26e�̭z��9G�7�Wj��q��Q<n�F��cl_+�r���ʳj���iL�>���O8�g}x��;�w�ի����}��[Bg�u�4iR�L�W��ˎ�L*��x������/~���=���?�%"!X7�7��=�<=+2���jB{����Z�w�3k�z��C���x�+��"Lp0C���~G��uR�0�t=F�� 繁���f2�LIza�uΓh�����~��0��Q'��&�3����O�Ǐ���D�x������N�P��`�|�� �~�Pi��H:"�WD���[m��A/$u�3*
���}��g�6�5xfF4�B!᫲�J�!�^nh���6����iiUR������;)�~�a}�u�,�U���쪖���H\��0�+��p��D]o�g8��JH-��^ޛmT���c��8p������mM͝f;�K�99[S�M�1�!��/##�PXhR{�X���1��i흣��i	ė���HA�t�U5�M��a�"��htUJj ��Yx��L%P����={_q�=z��0�7xŻK�x��v��74䨐��L�	�
"	��5��I�x�K$�=�ʒ4�S�پqa�&�;Sn5�ժ����yw�b��_�p7�}�ρ� �,?�����u�L��E�	��~�l���ӱ�y�؏����()ޗ�龳�VU
B��]Q����ň�=zv�ĦnY��6��qEaca	�T�s�G(W:`q��dH����9ek]	��N�?<�d�	^�SiN���n{�>�@b�]*�!�4�b�ٵt걽��rKo���P?��,H1 *��7��{���J�H4(���p���MfƘ�D�pT�@:����jO*������3j#y��0�0�4��jL9j.%�;b�F�����sL`�n�LIu]RX�t��ȍ�y4��%-~���{�7���r�t�/�j�w=ydi�O���:�ã���ֿC�e�/d�3���MYg	�9�DO(bّ`Ӱ��:���إ�n��k�N0���t�"K��P_+���oF��B�S��7oJ���OO�9O�_8�6��f%�3���8;�u�ͫ᛺bF���ѯ�K1y�fHf�7(���������+���-�l�<�3gg[7k2#53\��e��5�D���%�.�Πj}&������@��G���ƻ��1�!�
z�E��dEC��D��HTh���8s�U�����?��%���o�Sp����7��?Y�pp�|�Un���-3�S������<�����ݵ�[v�!�i^N>-��B3 +d�����e4�q�j�Gh=fͧ��V�t�w�`qm��:cmS��ּ9�W�5�o�N躧)��#}�.���<�זw<A��ms�F�v�Nf�F�������6;	Ƴ��}B�&�	�	~A;Z �e�}xh���0����ט�y�<IV�O�핳t�7S&l��Pj�����Ӽ���Z�����_c�I�+F"6B�X�A3m�yp��<��}����Q"U" b"PbD"bTM������������ϭ����~��&l��I�%6��(3��4�Į�`y�dhǼxOV���)�\�-��ގ��f��$Z��f =�!�<��`P,r�eo~H�2�e5tGh��%���ܵ�"����X��i8<�O9ȟ�B?���1ᝓܨ?D�I��"S��S$�'p�U�X���f�����4~{��(2\^�������Y��81��f
Gd�q#��$�1�ֻrvS�:���NWR2�]̫^�2�]Gk�sP&0�>G�e��@A�"m	����Qt�]�)[�;�ܸ��أ̽jl�{��������=���İ�@~����|����zy#���y�W�úFfFU�=t�����[����P��)1���Q���v��v��(!�8u��uHݯg�ﳴ}�H�[͇�v1���k��%9k�d���R��cbE�2���d��u���K�c��C�y'���C�y��nt���k��pе`ĖE�Yk����I���!?kN8b�I�����W����?��P�e���0��}F��/kՖ]/��ŰZ-���N��i��i�b�/�m>�d��A�?����{ʞ�y��O�{c�}�o����7��ߣ�j_-�E��P��(�g�\�ͥ�,��� ��?�E��
�I#�hʕ�W6��c�y�/_�տ��0x�M𫓽_�	�M]ٖVڙ,F�UUԧ|��*�w�{�|����=��?�(1 � �
�
B�BJ }��}?{�??��Y�>�_c�<xR���a �re=�/����8�K�7h6����F4�U�w���W�I�B���{�?�������~\]'���D��^�|S_|�n��'�ue�Ϯ�{�[�2�|z~c2��oI2!試A�r2�����=�oZ���״6�59s�t�l�э���Us���ڬi�	rnb�m�Fq���8ʲ����A�v�LZ���aӻ�`P6G�y1�L܂o**���S�Y�A=,�,�%լ��-m]��� ��/g3kxC���_�����>!�}��C+�s��t��X�>��A�=�N�1&�O5�gf+�o��ƚI��A_ϥ�F�vL=5��g�"z<����Nװ��d�7`s������EZ��2'��m�.�RF��
��q�l$vE�*���Dkg��ChI���k��M9��gtS5)D7�&�&X^b�sȤ�\h��/A�-�K��!#����f�?^Yon�P%�L	�,�	n��P�;*Jz�3l��c�qv���dto������� Qrƪ�A�L(g����k�v���'Z��ק���|,�F�VR�-q��v����~�:j�3��OP�ōR"3��n��O��z�v���;8𩳤Wu��w�Uj���m�TvS�MZ��^d���\��o�+�;lT�;����}��Cw9����,y2-�f_A���ۜ&e��۪X�$.���22)li�������VQ�;�e����Ջ���{�I�ڕ�$�_��G0N��72H
a'^�Y����\a����
��[ӊ(�K�+��O�Ɨ̋��b�5I��yڴ`\���>�-JSt��V�p<Rj_C��YtmgaS9��{ʘ+^���o�\2�(�!*������6�d���k&��0�/��!��~4��g5m<�Q9�y���߭�.��N]��S:�,�9QUJ�.�P��v�u���/{�9�Md�u[W�yh�.
S���{a�9M���O�1�� �P�#tt:}gN"U�MB�g��e���]ڷa�ۛ��o�y�|�:㻪�� �\�SZ�8q+{d�x�Wjq�ZtUD=�G��u���u��9��sg\�V�dEk�!��>��O&�'7i��$6>���ޔב����e(�SO���>G4`<�8V[L�����������om�G9CW���d[��ܬʔ�W˱R��˱��κ��*�2�:ټ͉���ޱ�s��y����H��k�{(���|{�,�J#~�#G%�A7(�~`�%�C�!ä��ʟ���=Pr)������fS�V�d�E�)E,@���6(��;W�{���ꑛ��x����ʠ'�HMz1o���՝3*��s���mn\���=2̎�8��h��#���������y�Q2k�8�(�7#�is:�U��\(�'��[C4�}�2m`��LPD.�]Zgi��-��7z�l�r�uQ�n�D�43����<��*��T�1��o���I��ܤ���Ύf�/wES�lPＹv��_�{�$��U!�1��ǻ	�N����1�e07t��E�{�{�����E�%���p{;�r�����,$(gU�bU��V�żl�v�2���{kX�@Й��e�^�/7��wu���qJd���{^��"[p�=y�\B�˧�*�D6��5�/�J�91��E�3�A�foUQ*����t�}���Q�/�7'7�a%aǙU����q��N��@�����iݦK?Aԝ�Fۦ%����+o8��������~�"Ԇ��_v#�j���U�ݩhb�^�ʮZ���m�i8�7}9�,��h��sH�z�8>K�����L(ݭ̪� �h�t0PW)ט�@I�Ĕ�׃r�X�g0%�+�ߝV�\�����Ҿ�Y�)�j�Q�ҫ���n�n�2wLs�����>�#������!�hmd��=�����%PǇ�����r~È���F�V�ҔҔ.�5JGN8H�'�ҔTE#���	��h#a���Ç���H��~�WP#~�4D����(��O�癥��m����8��h���4��ˣ-AAM#BPG��������D��E4�iJ��8�=<===8#�	�)*��h�4�RQB�p��ÇE!E�$E%S/��JRI<8p�������T'^�%1URS@�R�?�MP4P^�9�$�)�h� d���Q5Z1����u�Lf#G���{��(M4���׶(F`�~wU��S�X��d�1�l�`�+�=��7�&��Ձl���@>�?�* �H�Q*$J�H�
��������?��������$�/)��Q�D�n��uA/<c�� �j;���6�E�2�N#��*��R�LcӇ�>d�~�	�xh�Y�hY���a��E���e-�,ƿ6d[Vh��|%ϴ�v.:i�~���G4��x@P�И�;���'g��E�0��ݶ̉�Y�V�	s����O����A.�9��!��'5>�e�,�7*&����߰�ց,�l-��T�~�׾P�>�j[��@���g2dK�{���hf��c[^9�V<���ji�0��.�v[Ͳ;r�
�1%��a���%
�jC�c"���z��C:�	�h�,�isn��p}��jj�(:v~���#1_'}�z�!��r2킋��N�gM:w��3��s���|-�tj~B<�C�R�Tj�1�2	C���]M�C���a��щP ���FOu7�^eQ��f.���cC�`_j�%yH���2�P�leJ�3��Mݓ����4�n���ApޖDh�������1����1��n�;q�4�1�F��[n��K�O��ۼ:���}�4����O��wT�7W�m.gl��.��sGe��5M�P^�;�{�/y�r� �0�	�H;��ku�E���,�˫��g07�/�[z&G��?ӝ��2/E�=~�v��^P��`��r��n�7��������� @�"@�B!@�U�Q"S�����������~h�m��:�`�	�ya��Oa^���{�yV*��L��S�>Byb�����yP����V��/_W�c������VħV
��5)*��E[���xO@YD��?�����q�:�h~ �ጇ?h|�0�;�}��e'Xx�I�y�)�D�L-�3�'nn�k���L\ּ��;���C�<���ze0E�c��H��;08��]�E��Qu��L�1�mA�j��89���9Y׍$.�ݖ>2t���dc�ӳ�(��P�5�J��ɇ���y�pࠎ�Z��&K���F�[��w�w@~��y�sh���1��+������r�_R9�z��v��Ԩ�ը�u6��w��@����r�B5�{�����槷��u��k���0�F/�\�\¼���~����_>3�P����]�xr1{;���<��n���h�Z����r��l�+4�8���(!�����f4b�;?<]���N]v�ʬ�N�2�pr�O�r��l��9���ϸ'�yg���%+<O�ϘM��9��=��-�/se�k#��}�"n�$�:���!�I�َU�eE�rK��f��w{t�^nx�X:��ʤeL����c��{�h*g��U=��q���W�;]v�L�a΂�<.k{�eK��S3/]\H�!߫k�϶���Z/�IbU�F!�TbX� �D���Xs�ekV�3ԅM����d��,$h|.'�*l���:V;�7O�k;Oty�U4��v6.�]h��]�ϡ��CH��o�P꽒%��r���� j��&e��v��/����Q��N���~�y"{�3A�a�e(r����G���fƨS�����|q��^���N�4���P`��9�xVj�c��m��K6i�A���W�;A�6m=cռ*��"�A��-1��퐣����c@mW�Or�oܥM^�f�ܮ�a^���1�ޭ�p��D�ز�R3�'ڗ�����;�}��>ϫ� �'�%�{�Fi�#)���obTfW�Z�Ň�VW��(>C/���#��"�H"Gd�z~�`�'��N���5]�^5�&��	o�L�t�G�ϲq���G��a?1�0���v��~��>�vO4:��o�� ����ڧ�Z�R��8�].��(�X�"���9����������8���yJn���,���%�����"�kV:��0Ҳt�r�O�H%���u@����4[,m��ߵ|��X��/��v�ˍ��$���I3!7�T��S��=�:M_}�9�]'�X^gߵ��:�\v�|�N~R1��F�a�{ڽ���8P�Ե�l6�����j��������J�](��J�e2:�˛�k!��a���+nbY�������>�}�
H�V!�U"EH�0oi��y-��K��<6�3�-�ګ���e�����Tw:lw�%ݹ�wR��Iͫ������l@'�����2']W��Sut�c]�JN[�O&��`n`n�t`������)�8p�i_S ��i�}�:�cΩY7}B��Ė^.�5��
��߽I��DP`G����f����}��_��|�Qh\S��x��#����Π��{�G�*f�<a(���ڵ�Z��EsP��kƇ���TX>~1��/\��J��ksT�x��NW&��A�����%4]���h/Bq �/Q���k`�?��!�����L%�������/��jgn��׵1l���g�J����TY���4`ľ_~�-?V�I\5J���E-v��ձ�2�!h`�` =űZ#.�|�鶑f)d ��VJa#8�ý�sMt&7e�:��J�[9l���)���$�k�k1Q%��^S�;�"B�n�A=���du��<���y�*�}�R�V~�]V�+���.�~C0G9|��}����?b�e��������i�{u�}Wϴ,�Gk5��Z���˾��S��"�7ǫN�pݜ�.��[����:	��-HޡVA�@[�{&��ħY�����l����N��؟�4|D�e�{|y�S���RG�����{:��s]������(� B� ��
,@��w�����������~c��=��0S.���{�.U�3�Вހ��]	�����f>ݬ���wm���X����!��4��4-Z�*�OJ"�e�C�JzQ���yc�?���)�å�K����fA��0�;�Re��&u�/"��� �6]�)ᅍ��M�f-7d�O`��,�Թ�.m�1�3GeIOW�m�u��i��#h��?�֞[V�HZt������vL�kg�,g�^p������7[ׄ����Q�F��N(@j%s�Y�I璞>�l�8��u�ߟ�̏�&�y�f�������D�^��Ό��*ju��䨰�7}:/x�lL�_[o2������y]-5��ZA��O Laƶ`�5�k����r�4y�^�"ypu�n��\$��_�G0;"5��;�����<��lsO�>'%<�l��A�*�W4>g���˵H'��k_��Fq�mbz��^�9�"]�p0f�5�Ȍ�[��vְ�]�x�Ρٻ]v�l�۔�q`9�/��×}̻Ls���_8�����ޭ���yW�"���݆��$^mK]�S՜0.�����v�l�!�����1�fIg7�<��X�]r�8�szpf����j�˰�6o?/Vq�1^�
���'���W�)�;�NI�z���؝}I�������-�qmɛ�'w�PO� }�|>1*�B���"H��� 0a��{Ж!�$���# I��u|�����{�H1�'C�C�*<��>�L��᧻a���� �����ܴϨk�>bO�ϐ�Ţ��<�=R�+����"�U�q�v�;5�3�i�0���?������(U'�x�!����S�]yU-m��b����ٗ���Gc��82YR$�=�6)�C�?m�4�K
A�k@0G�\�g�}E̿%W��������U,���M���Be^Xh���5�B��׬z���{gh�-�V�AN�Ю�%����K�8�_W�4���`sbS+�x�tT	���B�FM����Q����8�مZ���k\�!��5������GcAðϳ�e'XĲ`�ct��IL%��1[6+��kft�wU.ȹ�b5���"!0%�K����!uɇ�y.� 9T��!<{pd���[a�~�V��~��Ԏ�甼hlQm�0�Z����	�Ln�vl�(qY�3�x��b?Z��w�N��ﵯ��w��=�T+���pN%�;`>��G�:m0��������w���LVBl���I��mQ�W�\�����n�9+�<Myv���!�2�"8�LYG�wQ���U���l���ƃ�7]S�2�TvWW9h��f;����p�e���筤�]�^��u�n
���Kζ&R�7\r��)@X?�e�UG�H�*�����/�����}�����H���0��ƖP�I�"�P�X�C9P�<W� ��1�zG@G?��d��&k�,�7L`Q/�LKr���Z������S��)���<�\�v=0~ΐ��8=&�!�q�-n�����t�/"��H��B⇳�+�T�9L�O�cюE�3�^=R͓����b{j���*C;T�fZ �DpL�ѯ��K�}͙̀��E��Ǥ�{�G1ኋ�M榅 �dh�ʸE75m�v3�.�1a^��\O�T��ؗ�t���$P��nՐ��Ͼ�}Z��{o���޸x!�q5[@�����2%�����2H��I��L]ਐ�k
�×�6��m3EvO�A,��r��o&���L�P��5���~�%��XN����3u=l����5>�zьG%,�rnWÏ{��l��Ui�]%�&��<*��_}z�ëّ�A!$0�G�P��q��顎_	�� ŕ�4����{�&���F��W~e7�^�6�_�u&8y��"� ��V=���>�j�qU�i�|IM5�a�i���3����$�QwNlӨEReނ��{ڗi>#%K3���Q��~|�Z��.&w��3P/��N��1��oq��K��L�&]2�+��wm��Ś)ɽ)���`�qx+�Ձ�Z�߯y.g�G��a�%���e�/Xɺk����ĳ�� �%D"!Q�@�%Q�T]��ｯ;��?����5�����J�A�>sȜ��+� ��d�z~�N���b�;��e��cD�s�B-"���Ed�������aoX�@�`KL-�m��H@4�!&ұ�]+
"����xc��p�Q�O��Rr��E*����1����}ƋaT	����?9X�'K��y��D�jpֽ�:ԞΙ��^;)��Ǥ���������Ao�<(�r|��?�۫?c�����f�3�}�S��Wp�(�W�H�P�Tw=��q���ۙs�Ȗ�����ݯW���<0B�k׿C�~52'|��"������ғ��b2mK������r���UWҲvoQ��b(�^ȷve=��7vmt\�K��H�4-Y�,:�x�Z�\!x,4
,�M^o#�Ɉ�}��-�)�?pE���!�qO��x4��9�C�3��3���|R�i��Kqg>�Ʈ���s������τ��񃏫~<	!�6�gh������#����lj�����d]L��!�Pv�W��������c���{��	����Oٰ���st�4�'����r������T5YT�8ڜ��'r.�"���^)5��%-�=G3d瘾Sϝ,u���]֐�&�pt�\��=�I�o/������V��9u��Kg��Y��{��/�Փ<7/��M�i��X���q�������~k�8s����Q?���(H# �(� �@�>X���6�C�g��{�	�l�����n�P��K�x��A�v�~"9�=��xG۝��|�ǒ��Hd)�	
���<�ڞ�*�}]�6֝ ���sQY(5$g�-�zl�`��WG�e-�.��^���2NX)=}צ雐NK���m�'Ƴ��s&V�<�T�ʯz�ai^�խ�tv>6K�9�z$9�1���P�r3�~4��˫�y} 7�4����j�>8\��[ί�J�QaMK�q��.PA�E-���	yڪ���t�n���#35�T�MN`�Of"S��������
qx ͑������A��_Oz�%��,��Û�&&�@B_C)�-��7gD7t�L�����h�A\h��/A�-�z6�>��[)�Yw�3^0D�z�РA��F���˰�6�T��c��"�ֵ�gi�\��N��i��<��];�|y؆^��n��oi�yVХ~i0���\��f�'��s�Y���g��~љӂ����td|&�c���PAe�t��Y�OR�Q�f��:�]c���+�ۧl<�\f�Dkc9Y��X�㸩�%��kOɑ��nu��Oz,��/4�W돯yJӀ�"�&��D
D��Z�h�?�d��F�Պ�S�l)�RsEV͖7������}��/�+ǜ/�oQ�x��W����#��ҥ�����s�kް�ow=�����
b� ���A�T9��?����>��|��G1���'�}j��8>�y����&/5�5g
���W=}����bV���W;*I{k���x-ԭ�%�AU��ΫՈ����ey��=<����%�	�c�j�j�J������;N�nm ��\�r`C�qjz�v�ܔ�f�wolH�!����ߦ�9��f��E�,�����v:���x�-n��eU�tFrf�)���<��N"��N�	���#�n�0�{����i%@A��MvA\���Y1ъ"v��zb��6�ʆ�f�_h!\Ln�OwP��ׯm�2�nB��`u@nJ���&2#��V%��Ek��R��N���*Ƈ�,�B�p������F�w	��J�+�ݾ��#1c[/.2;���e^Yt(�Ty�4X�t�	���5�L��&Ɵ`�-GQp�,��5���5j]nG2띬���Bl�B�d�ȕ"
��2��s^�=[�M=��&�5�Y�!f?.��0f�X�l����j`�n}��Bk�K1�	��N���,W��X���� �� d*��V��?s��h�Z-uc�[���K{��݈$P�j�
���Y7tqeʽ[�i�b���5g9�I�g=�KS�j��&(�.ϖ?�m�L��,��L�'u�����Dd��.B�d�Ze��R�X��%�hM�e��E�����Z�Йc.)Ӭ���(�;4(�p]+���I�4�;�������8{@�ɽ{-Sa��`F�|�� uV��Wy$5hM���?�F��Q׋-�svZ{սT-��v�ʒeV�8��G��P�yIWˬ�G-�Ak�����>mj���/;8�]9�k�G2�0�Y�^
�RB����ԩ&6狯$�=�J�[��a��YW	m���nlAבN�

��[}w{ɗgm.f��/� �N�׸���~�������z�ZOS_�p6��ZRS��|�;����.�v�/{`�k���N]�}�F)L��UE��,��{���rK�{p=����U�_I�[|.nCXcC����,ݒ�nmvc�̼|�g���^\�'�o����x�ڣl3B:OjIc��Ⱦ���Eg�i�Vcx�;���I�Q|EØ6�\C�hǪ����|�Fy�ul���\������<ɶ���}�$�X\۱��6����l��O(��S|��w^�=+#��=����c��Rs�葸u��t)��VR}�QwCk�Y�ko`�nc5����_.�Rm˳�;�;C{��G�2e$��j������\����?7eO��j��0���K�@�naLb?\<y���a\��:w��,����t����^��(A��*�� �IRO�F���Vzvɝ|�����X;�ZB�힚މ������i�����mV?�y�y��|w=U���-�2��ozd�,`1w4b�����[X�>4$�����q�>Q����iG�_��������w��\6]��˞�w۳ݰ�~Linn���/VK��e�uJ��~ӱ�d�J�5�=_/wA<����ll��CM��d7�V�I`���w#�Y{��"�Sf��G7#����7ݚ�^��'���h�t0-�1�,�e���׷nm��47Q���W>����}@�����j����T�eA�NT{�V�xe&��a�w��G���R� o6��9y�/��M|���2�N��婷v�K�Y՚�^�W�F
�b��C@ɜ:(3b���vֻ�f;.C��*�.���YQ�W��B:�x�ues�e�Ҍ�m��;R��hW�.��z֘xuЙ�����-ڙA%���}۟sb����՘�,�רe�݃%�f5��[��s��lM�P �K�vE]J���]g���.]E�r�$MM��:�$	�i����Oꉌ�A_s��h/&���^gK�h�Ӛ��]0n�\2�K�H�$�+񦜯�9hC����"��Y$�"D�!aa�:�ш�M���dmB�N��I��4��0�I��cB�����u�"J)J��h(*�(j�F�J"H����z}?�0Q�LT��QT%S@A4�g�O�M?�0y���))b��((i�zz}>��*ZZX���(��4!{�T4U/����������aMRSE���S:�II^�B��`���|:p��iB�H�4�͐���Y��BhO�Ç�~�P4�@PDAE4ɉ��R�k͟Lzzzp��(����S����H�kEB�T!^���zp�}���()4�'��0��DUQJ��D�O��L�	ETN�AT�;`h
��a1|�2���Y6����Z�o;�-��Q�@����ݰ����=�W74[w����j��#mo�%u���v;3|�7�����<���?��"�@�@�H,B$H�J�}6yDQ)�8s���8��^���;�al��{ـBy�hv�wL��ĲN��*��������{�P�e2���2�taqK.<���Ǒ7�����F����`��(�ώp�.�5b;U�sh� o�Vڿ�����E�w9KĐuXJ�������:nɀ��Oa�F�P��|�Z��۳�ËKMt=�"���~n^]&��x0��p0�X�:hj8F�� �ʭy�@��ǚF��V�,�>��\�5.[B�Ȫ2���u7�t;����^�<�@p��a����)��W�V*��d��b�u�LKv��s[#q��zSb���r+���_�l���V���g}�':����Y%Om[���vA�/H����òt���g�m��ޛc`ʤ��OO�=�}:��1��\��~n�(�(���v��������O��)���55g�����f@NN��~/�󢪗L����ٖ���=��$.g�{�׎�Oۡ���?g8�A�������6^���_u�v�xt��~��H�ʲ��@�yP��$�t�_E����~ǆ{B	zjl&�C�bq�vo���R~�Z#,�}̭^tk�o��#�5[��O��x�H�
�Z�]y7^�g���8�����[+�wr��о��S��p���|G�x�B�;t�ʾCd:]
�R�����%�ޑ*��[[�yFغN�HԦsu\q	�Gpky��l�z���ʟ����"D"""D"@bD�x=� �f��䙟�Ք�j��;���;%04
l��(.����<��Hזx���+O@3���=�d,O��Gd:�}{��U����{�5%L�ge0f4�q�j ���f�ױ��i;��Ed��0�M��V�t��1����1��U���	Xڊ�q�4"�&�bS���`�E��韆��t��E�_@���!@�"X\��`��[�� �W(�I�v<־�*���[�/�i�J��K�Y�E|��`��*��b���-U1��	O�$�ƯaF��f
hAWvD�Bԗ�tD�]"�$e57�j�p�G�@0-�Д�m	��c�x̊^��꼬�q���1��ʇ���|1��n�J��0�cן#Cy�X$;{�������\��2�y��2��\>&�=s��Ja��&�~/I�Wa���)M0���9͓"A(n�ސ!�C>�+��?�n���yQ������Qx�jCu@���6�]�>.��[�s��W����W���靇߳�}�B�P4~]�M_Pꃅ�ϥ���~2��朽xxm6`��d�1]ݜTC��ko0���l�vP��+�&ƥ.x{&���ۛtuhJKt���8�����6^��ժPwS�>Y[��U�V)�g;����6z�<ޛo�)̚�Yf=���r�ճ�F��(;����.���IA��(}��+�( 
�"D�D��ϗ��~r�&�{�;2�;�v{a�8A�� ���;���Dud�	�����Ǭg���<�݋�F&4�r��t�ϫ�UsH/� ��t���Pи�����C�F~[�o23^�T��G�c�~��a�_�g��-�,����K5Yhn���;>��v���lY,�Vn��]��9�_mM=C�n+v�k�n*@���C��ϧ�Ļ�?h��tx�{���Ι��S;�N�����Dtc<>���Nlnϣٗ�"����T[ ܺ���=FP\��z#)c�g���s7�E<r���o�4<����q���{>��?�L={T$P[��Yf^�lM�Y��.vyCV¶u{8ʲ��;�+jyu�	��M�E[P�!?1~���~��Or���q�"P<�ĺF�P�|=|U���`YI��[���.�~C|�Y3�U�ۈY0a��U�!��mat�6��Z�T�,)�z��T\:��|)���oO���"��2�g�ᘦsn���K����! ��sS�&I�)Մ�VQN.���a#�-�tcz8Y��_����U\ԆA�ݑV�L��v�Ν�KJ]�4��k�f��]��]5�]��+:��3gJM/�! =উH��Vm�c�q�-�j�����WN�6ẽ�î�%Ơ�{��)�(_Q��f�o�`����O� D	J�+�f`����Xܱ�࢛�}��a�m��fD3��p8��;,�x��y�Ճ��4�Q|2c['C��7u^��:��z�p"1�����%��CH�)�S"�0s�e<�8;�7�O�p��'�B�*$�fW��r�.+�e��Tx�QO�t�w�i0�%s�`7�F.�ʾ�s�ؓ���e^GjHO���>6�!��D�^����4,�	��'(�;|��M�.a�-ʋ]�M*��t��������y�}�nzY���=��OU_u�F�hf�S�-�8���@�'�m	����'[���`�8?���j)N�-ӷݢ�3��r��6������jR,�&��r�i�j[�� Z�y���ݜ�hj��%����˪�iзt(h�#�swV���f\�e�dܢ�/\a��׉�vt$�Z/�0��a�M�k;�t���חB%�������E�?{;������ޒ	�ur�o�Po1�g���z��P��P�~�`�����ؿ0��.^*5|��<ɯ����h��,-��lv"J�rӼiEInZ�k*��&V21s�m_M߻Y�R��z/��}$}ox�`˦qݢsb��fM�tw����ܴ�ԑ���T/B�q�gc��v]�nh�����i�.>u;�{{l\$�ͳOM���ǆ	�����rG�A��Ͽ�����"� �bT�P�*=ۯ�^Pqq�wj�#a�Y&*�!���O�2�7C�:�tX�� ����w5�0Ti�"������-���)�L�52�#!s�t+��G�=m�ap���ĳ�Bmc���N��Sw���;d9�P��;ڬNԷ7���׼d$���B�ڮ�}�x��O���5zr���z1d�kO����DE�O�01	�����f�!2��)ե%�jRU@*�&�#�`����.DA�{7i�i/���{�[C��C����?n�K��X�~�Y.�a�Y]3oo}:ҭz�A�\�wʆ�,A�NO��GܨDCwc@��ݔa�Lvi��'�7�vѹ5ݗQ��T_[C���bX׬�;*�/	���g��N�|{c��|wX꜆���[�s0�k�ʮUJ������9c��iC��n%�l���CM�Չ��\J�/I��������B��&$�R�,Qӵ��<J���Z��Sa]�\6���8x��ٚt����3;��`P�.=��}���c^ڒ�Ș�	�Z��	x�)�����|>i��k���-�^ڷ�<oW.ū<�}�������%`!�� �G�S�v:�r��'ƽ�
DI�븓��y��6�f���y���|�:�b�>�!��⌸X׫�����f�?<�w������}��ߞ�w���IeX�b "U�B$�Oߝ�����B����!�8���Eݛ]6�vm����e~�T��~��ƽT�ݬ!9�w�tU����f���g�����{��]���Hf��E�:�>��|�3+63bas7/d��b�?�����>��O��x��hY�#����xk�I_��^���^���w�!�{!�tC�: I�l�[�F�T?W�%�<��C�F��^y�����������Rӯ<�R�ӻ����%04�PB�Iw7�&���V�կ,񽩜� �J���}�l����6Lde:�����{ӥ*f�;(1aK#&��~3�h<���~�o/��n��UB�c۩���RO�X���b�O�����F�TW��(�x����su�f��nm�����ul�c1�9��������߄Hh)B7k���
by�\�
�;f��.l�@Y]V�%*�n�}�+�$ǐ#~oț����@��i�s�	�#a�.s��+�b峝&��JE6P	Mm~��;"��?�@0-�0%L��Jn)����L�����W}����Wh�g��?6{�뺛����{q0D��/a__{&^>�nO_(���sn5�iz�S��C���痕@���]�yjPro�^���.-ٓ� A�L}F���h��E�_g9�t�s�7�s?π��R �b ��R x0ox3y]�O>�QX�5���g��q�ԩ�Bc�m�)W��a�@�������0��D��׽���,'��SgrD��Q��YK������i�R�=4��(f����u������>!�(sӟ��� i��WW���B��es�Y��C�����u��[�Ƨ)��{��`4�H�vS2�0s�0��ȝu]R)��Xנ���,�
5�2�	Lz��p��fx�a��W߫g��ek���A�H�;��غ/B_[$7���Bӊ�<6�����h��6��~f�M��d�u�����h��h��P?���?yya�~�=��55�t;�����dh�R����
�&�w��5;���;?,�udtD�!Wү������=�Hvջ!��v�D��.��]��Q2]������ڄ-3�O(���2���x��pZDL"��ּ�F��2�DoA�b
��r�v��e���]�Ž9�C�j�@[ͻc�8 ����0���U�\�T/%�-A!��!���	ۉV:1��ݻUF��uIM�@�ևL>�}����U��9�[��;�_�l�'�	�l���g��Ŋی~D%��o��X�q�e���Q��p�%Ϸe�}����{�̂��-�j�QD��hg\N���+�߻���?-��}���@RĬHTBD�D�Ї�>���=��D�}���r�܅僸h�a�_r�5x1���A�c)��?Um!2�O�����|d�	�d	eIuk=>� ��V�N�����\����TȐ��'�}�+)ٟZ \��+z�!�=�P�Z2%t��Ǯ-��.E?xA�k]�OOvK8�e�+w'75d�!K����'�SsS�&I��N��p6��)��l�	܋hWv��Bm��j����E�{����[Pqp�H��n#s�H�I�g	�C���NW
���j7f�Y��}s�)�T��[�	̊��G��S���@���ǰ�6��RS�yd]M�Ta�R�m?U5rۤ3��}|`���+�$�T_��F��TI�}��B���&h�A���gX�험q�w���yd\�S�PX�\jO�xH>ƱO�!�������*��_v��#�����Y˃���)Z�ʀ���q�O��񣇹RH ��#S&��}f��]��Kt8�(����:��\�
�^��hN�3�����ȸ�G�(��鯋N�vj֫�sV�݆���o�}%�#"Jf䟣{������Ǆ �0��U�p��}o<��Q@3�F�ِ�+xbf��;�_����OP ���~^j���X'���I����#�N�{�k�����I���j���K���j�O/�~�>}�^y��>D���"D��D�JĴ� �>����������s�ϥ�f�!К}�<óy\�W0-ڔ�S�ֽ�s�}���J�#lz�~e���Ӧ%��^�ɼMz��P�y��K��yk��a�'��f������������9��9�o�|�ˇ���c�\$=�T	�r	��0�,�E���o�g޿۴Hy�l�k'��c*4d�8���T|}�����<3�"�>���ˁ����Y��Kݽ2����j� ˘���Y��U���Ghxj�:W�&�0zk�C��S�)��1�_|�l(^XV(eQ�w[���dκ��9}0��yH\�]D,��Ru��l�	��T9זt�Wp��t��U��9a`jj���.'^F�k%bv��r��q��W�������{�;�1UCK��i�~�,���Kb����4�K[�DX]^!��O4��%6�Q)�Ғ�4���N��M���h8A HJ��y,aT9Y^PT!j���+�'�ƀD��^�wL��6α��pi���Ό�~�&�2��tTSu�_K��Т�Y�T���r�Z�je@i�35���ohw��aC��l�Zy޷�����O�� D�^�[e$�ӠL��N�������R�t5�7�V�յ2��A"	��'���8ԗ[N��쎵��ѭ����^�p�`�lmv6���ċ�Tv,j�Y=;��<>�PO5,����������O�	J�,HĤ@�3xxD�Ą��5l?�Q}a~�R���L�t��6噃k۽4 ��a�Bm�4SG���k�{��k[�B��0�8����'���8.it�~j	�,{X[ !��t���*���د>?{;��YG3���Xڞa�ڲPk�%Te�Z�e	H�~ sIzp�$��"Z�fQ{�\�(;�(Ia�tz:�0���h��L���a^�R��r���^]���
��iT+gUzf}�(�������@5��?��U��K�9j�e�����T:�Ƨ��i�� z��U���� �1��=Ы�L�@�G�kG;����6��d����]L�ZlU�M�����ey�푷+���i��;(oF��pzin��ۯ�70���p��д�t��^&�u^o��s���e>;X��Gt"�x��=�S3ҁ���S]�K�1��8dC�T�A�f��q�9nǯKսv��h̾�h��,y,��R]���~���ON��4ΐ��>+ۉ�m�(gB�#�X+hR�����ʿ�f�祥�4�)����C��(p��6�EA���O�#
	`�ӳ�5�[M��չ\��Z����7�c)�e�	���zn�b�U���v#:���rز�C����𝿼��_n����v�d>�2��Ƴ�2����VKĹY%;�ݭu��+n�U�n���M����Z�1�gvT�y���ܲ,I5_=���`�ή�����i%c��n�������=y��*�ec��i�ɥy:s���Y�eӂ쉙���.�N��q��i�ӂ+N�&�`��A�<ޙ&�6\�{Q;uFL��m�wwʡgfe��z����O�[Rf��oB�:
���/}
E�̔B�&�`�{���m̜�y�M���MR���E����T�5ϼ.xt�n���=�-m�穷��ʼ�'�{�>�gP�Y|�B31tZ�����w*d�OWi�y��7��YC����W?^icn�݂�ɑ��]15X4�$]����-��]���!МxL����Ked���E��&�j�+A�ްk�6s�p�l�Od^./�ٯ�v��t�����#RP;�b#�.�={�W�.�UrO�<�l���w�<{yb���t,���WI�=;ٲ��t>���*�W� Gfr�/E�fr0�	Qu.�@�ްl^sk۲w���+���\���x\>	(�v<.���S�'��9yS�e��6�<�_c:�ܭ3�i�B	{+JS$��q
32�{ٻ�|G�E���g4��o��#��s+sp�{��U���Tu���=Oy�`�g.��ٱ��K�T��o,d݈����b�V�l�ö�ql������RLlX�{IL^ޙ��+��;���ѕ�~���Y�E�|�n�o3�M�y�P�YA�w�!R�MG_v����YxV�cG3(�ދ7��0�j��\�ϒJ��K��]7�V�Q�z����z5���	&^�r�BYj�W:����8R�ܧ�,�څz"u�����ضm_�s����#/<�	���n��3��M�,�#ˆ���f�6$#1̰�ԉN-��GS�S1�!k�%_nS=�\�(\�k`���L!�ݙ@З����Z�%������j݊���Y�a���FIŜy3ڰŒd���o	��*�^�<�l/V���)����]��2+v�4�����Ԯ��̉vT����`6E��Q���W���7���K�y^^&P� ���Y�<@x�^�X��p��7��ǟL���^�� v۔�VAܪ�y�:60��ywo������7u)���r�̽��-r=�R`��m��q����	���n7�y���s���D�p�����/�%$��_A]*�k����+ӝ�>}|�:]Y5`L��_"��T������{��^έ�WMAI0�}l��O��� � ��"�R��`t4�>�8p9�ei()*�)
i�(h��((4�"��*�xp�Ç8�RU55)E^Ơ�c͈��h֨(������DCE4Q]�	IC4O6�)�i�iH�:|:t�Ð[. ��
�5j(�F�*
+���4ġ�4zzp��Ǝ��V�HU%@Q�eׄ��4!�E,�AC�t���Ç��i14�D	KJD��ĚMA�MG8p���VLTZ4:�Ӣ�N��:)(�4���RE�\zzzzp�<��(��� yv��3AT��S��Ӥ(�����)*��/!�
)-����������>���=�_>����z�ɠq'��@"�	��I�\gcE��^^f��-�b|���z�5d�>�gt�]��v~����0�`����&$�~���߿ϟ���;)�����zE;Ǭ8��Ƚ�ǥ�[w*+��%6߸Π�F����U�u�VM���z;�u��[ռ�vgA@���LL@$<�vGTb�f�xL��Qvj4p��\$b[S�bYF�)�i��VW�
V���|W�7b?��J�[�Rfn�K34��P��`�O`�JuiH�T4���vH����� ���ڲ#cvm�ڼn[٦�
�L�C�k�2�6F�q=ԩ'�b`7H�
Һ�+�=�ʿ�ܮ4����/ϝzE�;�-`��}�Ƅ���"S���i��3!I�:��ӕ�1��!o<��W���Λf��\���0���0�a(֟C������D�p�T*��\�fe�ձ�33��WձHnl�;+i��/{� C$^�(���6ܣ_�a������j�	{E��_�g�7.��y<�}0=uз��%� ��?����C�E���ے��*�"]a�6v�=s�qs����[���T�4�����]�>	�?���t�Г�{(g-����nb:�};&�t)rrrwVZn��s�U����1��]�U��G�ԏ~��߽�^��ne�₉ �	ԙ��'h�2N�m�a����-d����,>�ze�e�m����wa[.�*n���NVN]ٱ_2��௨P+�3x0o7vo h�Q�e��ms6z��픜O�L(rhx��i~�,Z��re�������k��{t��{J?�b x��7遬��a���hP&$�P�.ŧ����x*�2�7D�ƪ��،�$� Q���A|g�k�a��ʮ;hNov}2��oA.�Rj�f蹍u/}��%�v�'a;*}kOC^m�P!��>B-�^�2/����W���H�	g�ԶM����B�����4��Hj�!�b�g� �t���B��'�v��"�-L
z��&�#xoH��W�� �'���A9YYh��V���q�1P�\3Z
͈��w[�3eKZ
�q�'��9w���5��zЃ,{�2�hХ`J�aM@�N5{����{��}%C�C^�x&�`��`�x+���0u�od!=�����2O`�Ju~		D�[ΡJ�l���_���%Ȏk�&~Uk��N7�C�@.�p�C+�l�pi��;�Re���s@��lj�A�Bu��)&o����}��{�<0�����?w��s�d	e]���ݕ%<���kzT�Ǵ7�o�-�-E��������ER���;[z�ޭ�NC1&�tu[C��
+"�+�3��}�{5ms{�#�D
3����>�R-�0�[:��6ɩ���	�� g��OK_���bT�m�ݱG;���ׯ7�2U�%�P%�#�2`G�o`�oxe��U$ך�Ǖ{C��������kߤ�/A"���<��e�^�M݆D�]��m�؄i�ir���XZ���U����,H\i�?|�A�5��B��l|w�߻�}tbՍc{�+T���|Y�mmGd�|T�Z��S~�Z��kA������(
������ے;�v�e�ɞ9��N4F��N�ݜ�и���(zW=����J�a(x.�\�/�1܊�̘�n�;����Of�d@pw^គ�I���n�y�nĤqm��\�Nׇ��!�l6E�]ٔ�{z����u�oa�H����x�e�\Ǚ�y�͒7�bK���Wu	����O�͎o���N_*�c��au�Y_)�5���<'��S�
��bo۴���kR�̽\�k�ƞĳ��F�L&��V���D�X�	����T�B~v��y��sB�)_��WU�K4^�����Ѱ0&ǆC:1�fF���; ��Y!
Dך�%�t=C�|5�����2LdB������w/�A�p�vMc�P%^�5��k��eAg�nT�p��6�}scUق���V0���M]+�|�P���Q�;8}+U���/��QR�j�sT�}5;CK ���Dߝ@c��p�C�c9<�H��xP�(�vwqD�l<�n�k��Բ�giW��ԥ�䚪[H9u5��b=R�)��D�p{607�xxJ��]��,A�<69����(�J�jXw	���,5�:���%
��_��
K�I���R�2(�\	k�����׬7b�b����Q)�=�����ƫ^��,%�nȥ�ټz�����Sۼ	�l��b`$��� ���~��(��+tp�G_POܞ�E2�#I��E����'���k���kԿW��C��#{s}�.�kq�T<�]0�ʥX���H��jw��Ђ�a��60\�%�J��}���K\8�(,4(�;J�O�)�~/I�w��Ƃ�0�ԜKGlӷ�e�٠<����i	�l���������	MB�����YB���ը�Q^J�s�No=M��4V��ݷ"��x���@`���ֿTķ�W��S*�OV0��+��PKܺ��|���WxY�uwD5M��&��D3r��`0jC� �^�������uc,�T;yR��3��ե�v*;��v�%��נW�q��P�ʁG�k���~�$t�'�s�~�:<'�0�a�ƩHU�[����"XK.���r�W�b�`�4����/Oj��(�r��
UçA��L��:Y"1�9��n�k:־���]�8�+X��lVdںŢ#�<�+�ef�h���%��v����¬˓��
�7}J��~g�6�8��7��ht{U���|�L}�/�8��Ds3+ݬȬ��ۃT�\�[�w���3��ૼX����yh��n��ؙN�3<�������A
e�tN5/,SЗ�z7�^�f_S8x��,
W!�.�}y��\Ѭ�����1��D4(��T�O�����W����X�|��卑�׊�`�a�R�'����̩�'\.�2�ߥK�P�ez��0!��K^D\zf�o*+�F�%6���6�΅TQ�I̬4�u�+���ӌ(��fR~���(}<
���# l}�v�Q���;k�L������]��(��	xd��H�2�F�?��S����{gOMn�$	�;5��]2芼f�[v��jv�|$! ������	�=��Js~JE2�$i5��d��d\:��\ʆ?7d��,�6̈o���2�U�S�yT?`g��OuI˺b���R��W0�b��S�,>G]�s���Z�w�/�΅G0��D��r�F��O��S>�,����������,ó�ۊ�};�8e	y��i窥,�B�yԮ�S�򤣑u�\}9�B��8pwR:��R6w��}��T){Lt��ש��1L�ĳY}�o�ӯo�74����g��F.��9Y�ޭ.w��d�"+�O����;��*��bC!����uV�OZr�c���� �at;!���Lx��������"H�+�0f����95�Hx���՜9�l�0��!'���gwi�ų��2��=�t�jdN������B��jwe�ّ���56�j��/Z��
*�h�O��ʔ����t��g揗�UQ����CQݵ�1z�r�<�����w�~��i�/״;5�P��`�؜J�5�C�Р��a�[K(rڞ��_/zG��I��'�ɠ��+��~�-@���2y���C�Ț������EM{Wh����\
z�ė� a�.���#��X8֗*���y�H��-ܾς#���VW�a�c��渘L;KZs����f�*�}$��mR�F����/����@d))v�}k+������E�bA�xC
ݟ���Uϫm
��C�P����Y�ϲ��<�/#2˄BFC_�l�.ql��/N��1b��F����\63��U���~��v�y�H�O�`�y�p*�]Z�@�c�1P�\3_�
�gsX4�u%�cy���{;Â�z#w���*�e�G.�"1�Cc���vc/me�v�)�yے^b�]��1�E'
���)"@�9�Ģ̘+�� ��iSjl���`�[4�,��s-ZE�R@�Wa����V�gV�P��.�ʲL,�ʨ�L��	��)��C���K��}��;#�`�q�$�/r�l�N�.�Р���Θ�F�+����pv֞���:��2�)C�s�iP*>^�R.���; �6��Bd���t�H2h(p�l^�x����G!N�X/Ra�k�8ސ��ΐq0�2�V�7���*�,/2K �6��rb6ڪ�K�:����|>�u
���*	]�D�b"1�E�I��1��/@�hjekz����Ȃ6��l�z�l��y���tӫZF׉��0n3Kb3c�0e�R�%�^F)�y���[�"���%��J疯Y�I��ET0�wq]����7̛r��w�W,31��ޜ"y�\�29 vN��⨰�]<�n�k	�{m0u�l*�2�����k0[�W�����!6З1�z�е~��qD��\��'��OG0��:�xɅFf̗�>�}�4|22U�����,/Ŀ��y�fW"���j픬���j�:�#a�&�*�PՎ�5��t
/C���@O ���	���?|�9��TXTW=.��*9��cO��\˩nJʼ�J�H4g"�9�u�JNK]�]���]E�ӽ}����jݯ_S�|�U���]�m^Z���yp�sxJUs��X��ʾI�m~�I�\p"g��tj�ߛ������x�b�b�kY��J��z�'�^�����=%�Jf��÷E��{�p5�rW�r�|<���Z�탰��G���F��^.���z���⻠�C�	���o�3����g�ftHf��Yq���n����Y+��l)�^����f1��2]����������橫��+�~���5Xׇ��e��e�L��\=�Jd�	T/hcOq�����1���*N�z͛`��_*`tm�pL�A��.N�+���-�A1�c��FpiZ�Y+��a><���0#内';O<��k��X��س���Ve&H�vV��a��oCc<��ux���<��Bj��a:�XJ��{���p���u���-^RU�7�Z�Ξ|)��$8-��ʘ	<�4+9�*h6�j����=���$7�O��d���U�&��)����D&]�tc��wʓйMbpַZB9�wE)�X�r��cƱu���A�a|��
���2Ϳ���]67��YfϢ8k��A�4w�Vߎ҇t��1i��%�.�AkN)�Ix�^�7{z����7l�xVu2U+�Ʃ�aLrM�S�.�<�J����3#�1�n}K���2�S�;@�~��]��ZR��Z�H�uL珘����He�i�·�.����+gٕ�sM����y���
�gB�=e�&W;fL�l�� �e�iC���_0�dͬ�Y�ӭ N�0�Ք.�*��zֹ?�?J}C�{�w��{��N��{;��#z��=��Xs���ֿP��ų"YgOV0�w)\�fr���L�]�1B���Cg�򸾕�A� ��d-����s�{'W�r�e���Ͼ�=�q�9��|+�� q���{��¹��A�ˮ<�}?s���'�����Zs���}������ߒNU0�zG���n
��Y<g�e`r�E��߳���J�	�f���B����[����z4=|��%=�|mT7h6��`�#�\Z�	5[E?�b+��� in�����fq�pWr
���8\�tܞ��[�m`n�!�n��f�XK( E��N�"��x�������0�Z�Դ�^��M->!@k`���.���^������c��v�{�{ڈV��6�m�����
�C�́^:����ez���EV������)��TW�2��d�\i�ح3�{�p�[���=Qb�XK�XQ1���Z~VI����7L8E����P#���u!����|8�u�3��z�yt9��e[����[νHlA�q��+�����RQ]2�ad�};o/|��$�{���/��]�f�Tǜ�gs����z)0�;��E沰����dx"[�����n��W���M�����Z�[�5
��!�	��9�	�r�d���j�d��T���ۄ(�|w�	 �c��{����tw4�D���`��0vI��B:S$�D��Ԩ[+�&��T<س�p�Nnqv���N��<�&��/!�E�^X: �x�,�C*�f�rzwJ����b:���H�T��h����\qGU���TZ>{?'�c���ahz>]b��n@��a�[�I�Z~Yqk*8��@VK��&4��BY
\�:��4ù��l!��ׇ!L��g8{{~�Nc����,M1�o�2�s��	l�e^J;���ǊJVQ�o��+k�ǽ_��?-�\��M�g�f�w� ��eV^�C�3I�_�;�'���F��H�8H3�i�o"&(�u}T�d�M<�_�H6bK�Ʋױ�z�v �s�/��:�;l��9�n�d��Z��qiyHt��&����7>e�c�a'��4Ó89��[�i��Ѥ;�l�p�xJ���y=�o�4 ��Re=�c�oֻ�HM*�7h6���K�~.��� {�
:�N�$+�w,���$=U1s+V�'N54�d]���F���w�\�7�O:�U �̓zA��Y|�]U�r xAeݴ�p�|/5-}z��n�U1�8rٝX�K�9�Z�^��#�}Y��M��O��'�i�4	}�
��;��{�ZPުb�3}R��1K�v�U���w��:u<��6�n��`3o�ӹ�Yj�k�nb�o��u�w*Ě�LڈlC�v��T���{��Y������&G��p��V��#�d=������i�4����p��x2a�0�s-m����#OԼ�k�㽡����q�ww!���W��-�>�g�5����d�Q7�Kf�ēz���ݤu��=��¯�M��z�>�WE����GL��pn�`��*еInۦj�2�T��G�^H�N��l�\�?6�L����n���f��q���o`�$P ���������#�k[��ɘ��B�a̻��K0��6�ZV뚻P^�/r U��j#�9{m��F`��Fi����&\���uV}֞[�Q䭚�;��>yK4���1�Y���M�?n!�$$D=��w�t�ಝ���Z�a��nR���f���E^1�ʭ�o��	p��쭘ޚ�2�SW������~�FOo�|����s0�Wh�LZ��G7��'�2�)�X�H��z�͵��nqA���8�N����;��e���l_f��+�	+����䙴�+Ut���s3��^VqMޯ�`�	#�>4��>�������1�F	��n��oќ�"�=J�6��F�8E���}b�V[�aa��M����������������m�`��,ʬ��P�TZs��q����Wo��UX��4J;�d��RD9T;Twt{����/4�A�Z�b/=��d����m�|���w9fM��8]1^ŵ
�*֕[�&�k+;B�E���ل]�J�6�Ϋ�Ӟ������V���N!��z!�lwx.��I���d���) �:1�u���ꪐ:��rr1j�؏zt��F��,��6*}���)o}�ӳ��딾� �m[��G�6�&��z6��Cճ�]Ѽ�C���'S���CBMk��T���y�t�ҝ���y�=@��QJWb��`̭(b����@����}ymj���V0d��l��٭C;�S��ӿvY�"dPu�͙��a{�o?Nb�q���j�f�LO6���l�ժ���f,��]�֣���o�B�����-� 2nl�m��E��-�_�[����о�٭&hU;ю�pjţ��5c>V9�#� �9�[t�&�T��T�Ѣ<��gK÷���f�p�q�y�)\�%�e�o��a
�fٴ��z ��E��&���}�lW2Aхu6���ڬ��nh�3c��#�ٷO�ᓲ�7��hI�'� ����MF�2#.	���m7F�����(bnD����!F���e��Q"�!@$*$h0���HU�B�Ɋ��=��R�%/�B�E&�!�hc?ӧ�����Q_$�AG��M�<&�֖�#^l�1���F��:i�zp��ƹ	@RZ�D�h)4�t�>	�<�kk44�J�A�8}8p�Pr)���m��M�D:t흳C���
R�4Ç8W"�)E#�ĺ�kjɢ�b)���PS�A�J1Ç8�6ҚTѥ�&�]���J��A��u����8p�qy����h��hti��D��h5���"���%鏇����M��A_�^`ą�R�:6(4!�49���������44��ATŢڑ���+E4SMR4���Sk%:5��V�h��JKT��ݾC�m�||k�THW��4�֎ԅ�;p�7�A;.�ϸu�M|���lնa�Fݞ4"��3j�4i���Σ���+{3,�jH��F)�0�E���x��h�],h���!���qtj�C����`�?������+Q���ݟf_H��xVl;9u��t���]��4�OP�A�'��z�m��l�̊6#G���'��S�<��smWK˫���xm�(�(vB�@���FCpΛe�0-�9iw�tH�!�{��&!�f�ij��]��K�*��	�����cW(���vOAd	d�N3�1� ��V#���mkb�b�7vOޕ���v@�HZ"K�j�<���d����X��P�Z2%t�p��)�Ǯq�M�T�^�|'r�߉����,�<���]L$�7�8H����2O`�Ju~H�Vg�-�(�N����Ǉ��h�a?v;/�:a��V_��#^�[	�`ѝ#��L)EQˢ�S��5wxoD�w2�I<�נ8���ώ�~xa9�!�t�`��N��7q׾�#��T�,�0ٍZ���C*ʜ׿QL��ހ�>���\�� u4������r���W^ud���?��Ύv���Y(b��\��f�'������0���c�=�C~�
c�����7��)M��yx7&4_^D7ў�ͪ,d"��(�;�
F�"�l�h�dW\�&��7�J���|��wG6E����Y�I��|��X�xU�SvF��]s�2v+;p�͔���#g:��`��w9�T�n�/u�7����0�%�s%��cq�����_�T��;'\]�*�
��̦�J���guW+CC�uk˹8hӰ��U{j�W;����-�?0�8PX���R�h�z�'��b�|���Q���Pű�
�w���=��Ak+{wZ�#�Ά�4��y��油�j���ֿ�0ĵ�=M9��l���4����4
�t���&4?�a7���'��l�����Uq�2xOr�j��8ñעfD�M�X�}��חx@���^��=���u��a�6���ϲ���$f+*�c�pLw��0{ތ��T5;L�[��<DG��/���r�?}}��
$���!��U�*�ʍ�v������/����8}=A�d_�������5��+o�gȯ�`48�#��^��	꽡��@R<��F�A��]@�:��/��_7F
�U���&v��}SC�)��,}	���ϳ�Ơ�Vܱ@�M�`&Sܜ��NQ��SQZ�;�����K�r�u�j�3)~����6'�1 ����;�b�|Β!F>�W.�|�Fm����<����l/<�w-Pu��c3����.��Gs�����ʾZfŻ">���en��|�rS�Ǽ1�����'�i[��%�+�����H�.��	�Vj�����سc��4�n��?�O�U�P�0y�y� �裡o*�Az��v?�Q`�AR+c6�^�=����{ų��Q�& 2N���8X&�4۞]���.؊�^�L�N��,�ߗE2�$tZ`���1�������]�UV�On��r���ؖ��-i�
 �.�8���X�ʆ.���ܵ;��~���QUӘ��6]����`�1�L���J�v�8qOL��1���t�lt>��a���L;J/��:lo��8�U��~AW�1��L���L<'T'g�sW�VP��2�j$k���]lq\e�ޔ&u@m��q̀����!å�G��6�*pLKj���nŲ�<�~0��DA��ӡ��먙�f�[΀]��إL�צ�6C#�O��9��g�`�~��Wu����g�������:�l[&�W�Ƨ�����~m;R� s�gn�lm��x�E��R�u�ؙ���M�m��w�L4ˡ.���lۄ�e���hr���ڕ�I(U1�YD��m
D��SU��7m�A��LNX���n�m��X��{���YM!HIT4��-�Y���5M�؈뮸�+zx�w>U'�ۿ�s�L��r��o`��G�QoX��5���#�k���j�l�G���q؞C���k`�m�`f8&5]-cƪ�,X�:�38)�̦�{���{��~�E�P���6��>���O��Rb� �������t�1�3S����\K>��H�-0D3$�/V�wgۙ}B+zK��B�����+�� 2�9�0�'T��[���`�
������|�#��u볿}�-�_X�'��A)ǂ�m�a�yt��'�A�6m>53��.�aŵ�Eޟ�p��k��M�}mt��1MA�����V��:�c���òxN�Ű �7zw�x�-��������Aߦ!"^�o۔��sV��=k�`P��@���HN(r�d����ebQ�I���=�����xzo>vku{�n�u�<{^q�T�-��萄�J��2O`�JuiH�IP���Fnj�jE����[o4����|C#��!���z�e�}���K0S�&Ou*I˺b���R�������$VLNCM�$0,���Q��ь"��@��^���>ܑ%��a�vAe.��D?a֋�鬻z����Z��H�U��6��0����t_��|�Ƽ9�?j�6�~���t�'�9F�eFn��'��<�@['�(Z��C�Q���b]�������5��/�F�=���C�G��R�޶8��]C����C�Mz�j5�krQ/�Sn�<�zU���`���n޶�Y�V�{Z���Ӛj!��7jQ����u@؋+ �vV���-�]��f���#G_�I�o
�jo/Tuo��]���p�[�p�b?K�^������N��|`�}]S�����ƻ=)8�k��̨����@lK�4{�8!���i�npr	na�ӝ�l:�;k�z_�'s�Z�Xqg�X�@�����H������;j���#o�����7���A�@�a��,񁯏�T_�ϓ{�6�e'�~�aC�@66���./��]ЅI�=�������q$��#��![�8L��A��p��LIz��XL�j��9�\�å;KU9wn�|�r����B�����k|>n|�<[f:���'Y��>�$���D�j����@�e�|_Z����6�ke��
ށwa��a�Ň�b���V-��2N�v��{�u{��F!B������0KtM�]vQ��A�xGDU���!�DU�옩������ԯW��l��Ϸ-�2��bzW$�W��;yTb�'@H��4F@t!H��j1t�X!g$�#*�U)�z%���e�]�zF�vJ5�[�Y���M7��d$ 
���RV^�KA��U��Ǿ�A���.���CNB��
�OT���v:�l�e�tM����T*x���ܮ�)iB��.[�`ѯ���^���=�|�J����i�A�찆��}��b�&��S}0η�i�졽x�U�<'f�Z�R����������˻�/�|6�|�#r�O�2�2�.D��p��Ѻ�iݣtU�ǒ����뒾~�q�6V��3�xc_}�?Z�s`�;K�ʳ�]6w�\��%ׁ�*���~mK3c�&PF����ߒ�J�T�f���[{�˳wTS�������§���>�I��yԨg���i>
�zp�z��$����ں�F��M����R�0���\�ap��z>����̾g�v����
���+��ؤ�K��X�aˎwJF�9:�%���9Ol��q�틐i� �hM#zb�
�o�WjF���_E��"����7������Tk�E�280ސŧ�,�e�6��'e��&/79��kG[_Tx��︱��1�WH�q��΁m�k�M	��μٮ6_n%<���2�7W$�$��5�/�G�0� 7�	"�?w����B��H�7��(��F�������9��ˀU��,�/9�Ӝz�T�Z7Y��F�+=��4��]��8�o�`��9��V�t�����74�2l�=\PU[�gy�1�*��6�C�T�r#��ϾȝҖAC,Dغ�=q�E
iUyC1�γ�"A���m�q�׼:o%��_���L2���
k�s�Pf��w���ͥ>t�ps��*c�E�N����#Օ�d�͍�p�PF�<,��թ>=�
��TdSR���o;��jtl)J��3�>;W Tә�[:�dܹ"a��mY�)�AH����ᵙ�J�����0N�N�JJ�O�7��i�uXH��S�م����j�:_s.��z��Ғ,�H�R������t��u=���d�_�:x�M[�}�=����k� {�M4x�n�7���*z/�2x�fY��w�]4 �X��u�v�*���mloI��"O\5C�S�ޤG@��޸�nOb
���ڲ�����	�z���x�]X�z׀�"?���i��:��y�޸�S�+a�F~��'~���c�����D* ���ǃ���:q��Yn%�pbk���憭��6�B2�jWf����^�)�,�v�)�����YE��[���{�_F�6����\�Mxx�v���P�q�b�xoT⭾���-�Y�χ��c�����?j]�1�S��3u��dm�t�F<��Q�n5������~hV���+�~s�=��������ZgNsFh=��n�����80aP\�ȁ�i�w��~���;ѽ�{:�e��62�GuVƭ��m"����f��"Ҝ���|�č���<����ȏ�Q�k�;�~�F}�:_� ���/�t�E\�̻���h�Nۃ?3�z~7t)]�ܖ����+�Z�_�ڃ!qc��A���3����\�հ�_��LeZ�-�$?v�`�iͤ��:�3i�Q�z�"�Q#/W>���r��U���f\n��� �)�$-%�]J���@�d�sb�Ն*yظyd�__=�+}޼;!Ԋ���K��m@��)J�3���m��u�c;.�ex��)�����)�9�5�Sz8v��6�}C�	%J��U���k��>�g�,yGۧ�Oi1T/;�9|�!�UvN7G������ޗ�GX�T�qK�Y=�����ω܄E����P�W.�Y8�Zr�5hÛy�寷+�{�J�A=܉YzwD<�-�*�͙D����5l��m���.�v������D��8ˌ%�p���s<E��5�g�O�S��H@�Nhm���=�)+�:�ƎKw�f[�{����x�>�Q�ޢp�f<��r�`��6�϶�˫��x�1����������A�����?�ͧ!��[��r7������o1��#j�]:���+2��3"��"�%U��
��4ݵ��\�j����*�>^�a�@��&Uu�ʮ��t�zJ�S��-���W3�C��U�{���4Y������ŵf�=�^v;$f�Md�mNU+�9S�������y!z�5� V��ĺ�}�C�9ݤ��]��
�j�}�l�������C>�l
��vG$�n�}��&y������w��7��ԑ_����I��E��;P�ċ�t��4��ZxeB!���5�r��^%k��� B�Z����6!3\���6ZG����D�+�W�|�C�Ay+)ۮ�r`��Ĭ����l�������h˟��c$C��g�3ʟM�2��4�����P�|~�����^��ED�i�t�};�].��k!�.�n�o�c�57��}Πҥ�o3#gs�.|tk�ݚ����g��ﯼ�<�{m�h��M��]qep��t��B�/k$j�n�gW�)=��Mc993w�ƌ��bO�gd�Bé3�W�b�q+hvM�Z���b��n�δ��G;y�m�H<�0Eÿ@Yl�8�u�W(	:�%����Qyi�l��f��l����$t���d'5��6�h���%�<��B�'�n��:�e�{��q/p����2$Z���B�V��M*%�q�n�%��V���8��̒HyR�l��5S��z�v���;��_s�͘�f��]�d��Pv��\�^�+�Ը�>㿠�N��_�׶�ɏU�G�����hX[Fb����)�+��(�i�� �:N�h��|�no<�.w��4��/̎��J�J�;*���-V�Gr��{���vFa�x�����]L�q��j�0��z��E�NXܞղ=@~� �ӵ�Dđ�vl����R��S�>s�Ħ0cJi�ݪ-ۼnaɵs3�I,�f��;�I��+��6����y�&�e,�5ul�LseZzo��y��#gh�*Iv�6�2݉v�;�A�C������F	�M-\�7G#ŏa���Щ�$�a��o�no��r��Ue
����j���f�����s��G��oUs�=r�w<Mxei0������s���j���]�L��K$LN�<�sya<�F;�ziRFꯤu�Y���`�]j���o�V�������o�����3�\��4v�;���^Д5�m'&�q��wT㬳]G�cf[n����U�|N�2�=*Z��Ϟ䝣k:k��c;<,z�޶�A�-{���;��������\YAj��Gw�����eZܨ�V���A�y�Sa��B7���<��[��b��FJ���)p��A���M�w���]2���)�O=���u<ؑ�7�F���/����Z����픳h6b�TM�m{_4��[�K��H���@<ōK��TFZ��2����rn�h-Y����,�nv�{.�����>�9��b>�LjG�v�w��Kd�to�;�V�vܶ��aqVE0\.��Ne�Q�ّ������J��/u{7����Q�T�[Un�!*]��li��i�R@�Lѡ�:`e]l���+�f���4޸��pU͗��_@�����+��+��n�8t!�|g]k�t�ץ%�L��ga��
j���;I�иA�*u"�i���Z��5����@������{&��'d���J������(Q�W����F��qI<!�^�.�_pi{��p���Z�IqB��y���ݭˍ�.ܴ����_ `�_�3��m��f�U�_��T-뜳��[Bw���]��`�qk��47��y���=$��5�Y�M�JioY�R��cZ[�M;�<;�<uPͼ7�!ۃ�ʵ�VqU]s��
�:ַs]�\�I��>�"uc��=�����zC�Ώ�m;v�z��8����r�����m��0��<�����ߕ=|7j�VQ]�܋b����3����gX�DU#j��=h����V���{Qi��B�ѵ~�N�y�.�Wfs��=5��}07�{�4t�����"��0�Rߛ��Y$�b�qѣn??z��^:
s��諸����ꍻjB��-�۬��"}��q�y��M�'Î;nQ���׽!z�zF�y��>�w�]]s�.{؉�+C�X�#{ۜ}8^鞶Ҧ{L�E�˂��V�}��\gJ�ތg3�����F�_A�]�F\���Q�U�.�WM�s=2��{ۉq��6T��ۛ|��[�ؤ�ܝVL��:�/ߟ=����_�&�?#U�;d"�����@R�!�i���=8p*�!@���'̍j�Ɋ��F�:]��it�(�!K�)6��5�==8zp���m�`�ډ���:�4��}��>K�lPU.�F�m��f�#����Áʶ�X��i����&���K^J�6���h4��zp�����IJ!��M��+E�^�>|���UJU�h������ӇQAJu$�QJDP�(/ph�h4���(+@[5���Qk.���-��:t����S�6J4�M:��TŤ�@D1	l�Z�Q��j�Ǉ�����

�Q��5Qm�[FC��b<�F��ĺ4��~Z(��C��)����Ӈ���
-SA���)��ր�ETԚ�Q��:q3����JѤ+�)Ļm!�hv�:)���E�� �*�Q�_W|�ڍ-ww��
2��9�����=�s���fن����}s��ֵ�fJ�i�,�$����;�!-�~�oe%Z�^��>�,G��St��ho0�A�
�Uw"��`����sn�u�)�Is�Fb�-c��b�F�����x@|Ĭ0.6��誎�ZC�����u�*�2g�9^& v��4�:��9�+Yȡ�-O_v����(����c2���>�H�J~�Lj���g>X�m��V)�]�6r�lJ���y|</櫹:�e���/�����	=ɶ�Sq��ef��t��EE<{!��9G�I���x~�VZ�VYC��42���ow�'�ؘ>7�u�f�C*���8C���e���,!5FA��x��ݦ[��}�J������;W 
P�E[8@�,�"	YcVVf蚊}�1C4��E�,�%����N9F�T����W;L�i�u�3��'u�\��nod�	Qf[h�m���ԒL��d�7�S���ӤOvT�j���P׌j�~�\�sw�r������t�B{��s��=����LѠ�xM�PD�1��4ͷ��T�h��<%�U0S���Lz�4���H���E��땻��$��lu����5��	|�i��[�iվ�����~|U�s�����B�a�[x�Y}��܏ŁH3|1v��Ǌ�v�}�U<��hz�ɮ<���� �B6V�oI���[d�ї�[��U(}�����r|��`��N����~U�O�$G�nb}����W��S'���9�P��A���L4@�d����j (�L��9�4c{��m{ae׉+��LM�Ja�yI���0#�8�ˍ�Ǵ����t���j7ޞ΅�د�ǎ�:CnsCU?z�.�f����(ܼ
�����bt��>�'���n�ލ�v��OhS�U�z�����C�c� BL��1)�;/�q"x��&��ƞ[o��Ϡ��s��J}�Ndd2���v亢�}�P�%��^�w_�bTA b.�`�pv�)Aw"�����.w%��D��� �bg�����l��9;��t�M��{�/.�Ռ���ݏ��/�I�x6����N��n�e�#쓥��łB��{7N1����'�ۭ�釮"�+�
Sr�y��k�df�8�:5zp�0�jH�/tQ��g�u掝�3��fK+J��D��p á�`J��_%����!��E�g�͸��	�_�m*(�[�Su���3�z��XF�Ut��d\6OomZ�j�P���\�N��҃ ���ݑsO�	"�ҸOw�4wc;7�X�"�-�Dwjk[�����@$e:���{OPm�1����#��nqfT���� ,�P!>�8H�]!�%���%R�ؙ��ِ���i�Ѓ�ėˍ�~��y��H7�)��p�	�j*�StnV5�А���7Y��\�"Hc��}ݫ��#1�m�C�A[���շ�~�:ŗ+6������;4U.I�mo�d��T�@~��-��wua��{�;��i^w]t�\\v���:��(⻗c�.϶ֆmVwH���_s�+�����THG��2�Ly���9T7��z����
�$�ќe�7Z��������%1�,���=�������B�g	�@��N�n�Z��l�>������q�k5Mj{;�|n�v��=�f�|]�G���{�(2;s�����(��W�K�-��Wξ�=h��+���BH�=M3T�tX/��j��#�M�(���%��5KF����Y�YWmvb��e���UNf^F� ��;3{:�s�����(�!����~�\,�ӓ�ĺ�_eNt�33f��SnE�n6Z5�����2���ÚF��꺄rJ�F܆���T�d��Í(OtP!�t�7)�%���F�ԃ� ����
�V���kf��V�P�Go	f}��7��3-<�������c�ڮ�v��g�,L����E^Zw��yՇd:m����Yq�f�#�dqY��
���U��,�c�;|���5��;��ƙ�G��1�-��A�S�^��/�����ޡwssk��D=N�gߍ�+�惿,�tF.F�{
/ݕl�2;x���7/�Sъwj�駉�p��Pm��4m�X�^�kx�j'�[.]���J|c�6J�˸T;vFW�B�OO����j:m
ﲰ�t��'woB��%c�T��ϛ+d5S��d�g����_#�[�SF�7H9j;_�5h�
�VS���r�}�:�]��ʦ���D�5ڭ8�����;s$�q/w[V�N��'���~�wraY�N�Ӆ�N�njbo��v�3�#|��/shj:���:�.-���at�2�67����ft;M��^��a���hxڎ�O�rU2��jX��L����u�oF�uV�vuM�eZ#0�!Y����@e��c���Ԫ�ky��i*�]�(�K��vd32z��hnQ&��k�K��2\]�t ��ȋ]����-��n��$M����W,�r@f�p�#")�������0e=B��zK9�q�	<K���_?�}���>�n��h�pF�8�2P���}Z�v��_��/Z(�~��z�k�;6��Y�#[���ZSO����q2�4݋�e��[�3ŐZ��:)@ź��N�V⩪J��c��ۇ���EZ��2��p�D�$�R&��ȩ{[��tsu�3������I�@��Y�=% D��^>6a��gt#d�'�˹m�ǭ��m�d+ik�׶�uxx�	Q�UQ1մ��Q[��[��rN�tD�YK��b�{�z�\Z^#@ŝr�H!>�-e�'L�Q�7�=>�Ȕ)�����iU�|��xN	-�żqR�}�]b��d�������{=�xP��Q���Mm��*��.�'v�2�
������I��)���|����m^=]�����Vu��g �e���ر%o�m������Y��Þ��]��xZ2�)듵s�sV�7&�R����d�ޮj`6��H^9�!��V<8H�Ib<����6�2���[<zj��TRמR�0Of�ݯ�ar�:`����<;�$Y��L��
���9�B�XƂ�wk�w�{ [8�b�秂�bO �'W)Ey�Jy�5�f�X��bgy��;����M�<Ԃ���շ�N'6�,�m���/G35��lp蜔�$�����;Z!�w�7�� ��Ow���c��h�#{%�#��'�E/ ��6�5�lv������8[�L��̍�-6��|���;#�mw%��SR��0cJ}�o��v��x�kk�SM=�{FX� n�6���]y�^�8x�`t�=�_,����p%y������\����t��룳�w�AAVe#ݽv�!�а'��U�,�{`(W��{�T�Q�Bҋ5o�:���f<���˴t�Nw�Oo��ލ�❱:�nե(�}�	�K~�ɧ0�I���7'1$ri���*(���c�q�U��[i�f0�k?�Vl
�e������]�ǲ�m|��s��y��]��`>��-��j���7-*�a.����l��Ege������v��x����r�wW7$�E[�47 M2�7m�{V����k�Ĩ��{�h����%�s�!;U#T���NK]1���y��3V���3��m�\,��ú�}t�6Y��mc�^8֞��eL�s;d=��)|�[������aJ�R9��N�nS�C�Χ�OW��2$@�pJ�
�"WX�A�t�!��)I#	��_?[�C������q�i[��h
G��H�S	� v.��	�i�����9��Z�wiь�;�v���P����kL�h�?�T�s��LN�{�5e>Z�����_I��&@'WQ8XO��<k�A�!d��È���C�*�K���_G3{�]�Mي��{o���&}��X>{�����̇}Q.�g\�=s�e~q�J�!,�Ն$]�`q]�"s��q��:�_��\�/vZ�ת�֦�ŹQ���ʲ��4�|n�,��K|��A��V]S8�u��і��m�bx���"��U��:�S@��[0Y��0R�n�
� ��55<�\.s�u�M���͊q�*)8Rd�9#k���+�QEw.����m������0��f��3��W@|;1g�*���po%>��b��
U֦���N��P3KݛǬ ��<��.����O@��6BQ��_V��{��{�-�<�s���H������n��@6�B"_�0
ӓؗv�A0�hc���Qś��%�̺F(�h�Pc�h�q�;:���w(�����{5�]��-o�Ci0H&7q�L�:(���d3����3>�r�g���ܣ}m�����fY���Ǆ{8>��^��.1g�M��k,�8m��_��p�vUz*�Eeǯ�^�#���Д�:��������y�4�%Q�����(1�q�!��H�Xt�Q�3g�d�N���2mJ`��-�z5�6%�a���ї��Ҟ�kn-G�Լ�D�i�Rn��Q�f�Зp��a
A����F�#�Y(�?�p_���j�_�"��"p�����%E7/�7Q�nԽ��=wW7a�_
{y��k-d�|'="�L��B���d�&,ͣ�����Y��<ϳ���Y�^�VH�X��^k
�>w��e��1 ��b�_��9�wU�c'��5ANN�j�=y#��i�<�����+*�n�U#F�c�Ӏ�Xs���	AS����n�̏H�	!qCw����w�Yvo*�j{�k:�F�{$��R�-�_Pk���e9�l=lk6U���݃�8����f-J�/�rS�Ķ%>�Ͳzz�rZ����B�e�n�ˇ-�c��OY��ؕU��"�%_~�'m	�����[���\��~K�� ��kr��Q�g�;*�x���P�!����4�j����t���%���l�L�a����W�Wu!Q�t�eƝs���Ov�va��J�����h��Kto�h�pF�y�)6V�5򛇩,�ǚ��Q����5?�=8�{ vz�zǰ�8x�>V�hK���$�§�(iW#�&��h�4����Ѧ(��E-q�8ޅ�g��g3�����|(g��,�+ԟs��T�����.nái;���#�����K
f46��Hg`]}����D:i[B�jZ]h�ĎoU�0WbŬ�V�p��7;�6o�l��������p2�Lh&@��$�pA����'5��ƚSu�θd�6o�H����үEZ47l6�[n���H�K�>K�8��ϳ#��1�tPKHh�~�ؿQ�Y��%Bl[I�܌�C��[��ܽ}�v�������QOYw�=��9o�O����y�2S�̕^0dVX�mb�Yy-mY�ge��G�˱{×!]��/)z�\��:����Y��R�O[W�;�^m�f>�sGZJ��Q�@;W�4�/�.�+"6[�l���G7�TR�F�p����R5B�l�P�*��Cu��2���W�M�.u����o5�HU�C$@nN:؈��=Ғ,�p[&I���Q���DΜ��-�=��gx�=�j*s�0Ol�u���<��ʑ[4Z��M�Xj�f�ř��I9�9��ɶ�70e��p^������ {��қ��LO����놟oxD����s��nE�Ɠ����P��3&	81bQs���WդwH+��l�1��qu��C�m��"�W��H��,t�\���J�	���p]n�����y�t�����Ym�>�W��z��˝��+0xg����h��m�E%�c�r󶽏����q���sg���aO�����ˤ�U����Ϛk�qA���O
l<<֚|��5�W�I�����Y/T�6�!bW�]z�Q
�\�$x=Eva�U���t˥tĢ,Q���c���,�`+��y��)x?H.��R����^����ݷr�s����sfP�Y�ӡ]�6�������"g);F)"\�X;h��ź�MY��x�O\����҂�U�p�OsX�Ts5E�0/�]˾�۾����ܙ���,��h-�&;�����jO���C. �8	�<#8a��<=�mԦ��]�H]��_Q�*���]�d�3F�⼔����Ɯ��m�Tt*�z_u�27F��ݕ��k�24�C�^�ɝ�V=˽S>m��W��
�[��B��؏��e��k}�����p=��v,�m<�Oo[� S��HӜ���k֡�D���������PS��z9q�&J�V��]��*���؋��9&���dFʆwn�m�8�g F4�:�h ]�_w�䋉��{㪶&նla�w��cp���N$�]N���Uo�/N���i���R�w��4]B��sOu���M�Ιݘ�	x+S��r�t31Ռ�(T� *��v�!������2a�c�og�d�9	��Ӗj�;G����aӓ�I��aj�V5�Sp�Ҍ5�>6�ӂw���ڻ�d������J��`0��=��<�q�L���_{b�o��<�p����㼎���d]��$�;�ȫʠ��"��I��%�`��A�NU�g�PF{;&�D�;>�����w^��yx%�a�I8����P��mZ�˳�^>�
Ox$���1w��r��Wd;����d��}�=7|�u��N'����ԾV��C�w��[I:�:�7q��`rh�8Wu�\#&�Z�WMX��k7e������h���au��6�on�f)WV�������̒� �kG[�M�
ٚ4h�f�i��γ���]b��'T%bm��a>��\Ŝ!��R�𜹞�R���J�C��Ξ+4-̝�n9�K.l{b[�2P����_�̵�d�3��Z3��=]w՗�R%�6f8�!��]�A��9�l�d%M6gV=�������ok`����Cs�R=꾾55#1MǙ��`��}!�,X���?J3�����ӹ���C��&�3T�cG��ΨNX��~��U��^R�Zu�$��/�<����s�z�{�q�Mf�^��+�^Nh;8;��N�az�S�E\�ٕ��xB�t;�o�G �[�6s(�5�KY��7��.��fN��]�u@Z�Y�bH�A�+?�fL �I�D�	RisTe�p/�Ƙ�*P�c���(�@�Z~"@�5Ш�,��j&��Y�d��E��摏8��
F�a�Ba�Că�i��j��S���h�b�����UCA�F*�ͪ�"�*&�h�lG���??nUS%ӪY�V���QE1Θ�A���Dk!\�4�8p��.El�Q�c����ڴ�l%�EF�UD��E���6j�k��5!�����#���y�
�]5lRDD��I��TE������j"/'1�ӧN*xX-�
4�Th6�v-�Ţ���F	�J(
)�����yLS\Ԛ)6�i�AC��[km��b�j ��-�3��i���j�	�OOON�i����**"Ū��h���EAE��yh|�H�l`)ǧ��Ӄ��㍢��bJ(�1U�<�
�2Q�4�iӭ4D[�b"(5�4��li1������*�)�d�R^��b�ɚ�(�QN�Ѡ-`��-�uE<TM7��4F���D�Q�u�j)��7�h�EU��������J�^gU�s�5�CwP��?j� sr��#�$P��ӽ�M��<3��z�&�)�7ǌ��)�	�̖፰}�~���}�S��pP��h��g�견�eqzH�Gst����kn���a7��)���HxcjYU䑉�.b�]&8���r�I��ˢ��]v�y���r�7�ވ�&`	�����MD+�7C)>�a����ڈ����4�#�t8¦Z��=Иo�|Y^�S�OG�Ȫ��/}n�[��=k*tP���0�(m�b��6(n�hk��4�.��Y�)QJ����#*
½Ӵ�5�����K0f�s�e�W3���_\���C�\�y�{��Ba�&�ې}B�:Z��W'���ES�9�m��لQ�y��(д��/޸-t�b��KX�|Z���.��,eo�����e	p8��v��l�&T�^������TG[6V�Q��E��UU����b�,)T4�����2}�������{�Y�˷��+�[y����WGqS����Z�	�^tM�+I����[�A����C[��w,�����*�9�P�S�r�!?�D�I �9~P��V��N�Ӹ��]��lg˞TA�WS�ې�gǺ����<,kބ��mp
%JU�I�Q��	�kÜ����`a��(B���j���CjW)J�^��\�hn�hw~�wV9�{�]٪�M[8��`�t!7��L�mH�?l�����2y�$�U�EUy������D�{�:A��́ºЅ�Z��yZ��0 �g��dm��=��9�M�duu�|ُ�Ab�9a�e�ͩ��.cg�8��aDfA�ׯm%4\�>����=���E`���Kc�ӏ�9����1H�b��TϪ��0�IEܻ�-{Oq;8r����)�c`b<��#�����U�����.�Uw��ҩ�-�L���=L�V@�al p�L�q���nFY�ϧy�}[5��n��S�޽����*/hN�	���m�׃�I�d�G��U3I��mN>Ʈ�m��v�23h���+G@V���N�;������{�Cz�}]�Qpk�rr*�Ĩ���r����H�f�ˬ9�y]\01y�e/)�^��*S4OyQiK?��Hy�*�e_!��5��V⹕�qwS�:=J>���i�6���]w#����Q�L�,�!*x�����F}�}���;�;�K7���=#y��[��^�c��{�$&0dfTJx�o�C���t��s�_<��D���4�@��=9�vn�s�J�y����H1E({�5��yW���^�C��o%�k��>h�5��emg��V�2Z�B��xXJ��L�
��׶��9�N�� ��6}�:�8�=Rqa� ����E_����0�,�� �w喎�.a�s�~�X�QTV�(xG��L����;y=4�L��
�%�zh�z(��l�;y�xfeĞdR��Ip1ƫϔ�k��T;2��qq��YvƳ�]T�4��B��(3��/a#c�$�s�K����T�[R�=N`ι�Q�g�a�b�χ�G��*�ax뒫L�6d��C�&��7	��������_B�r��S���v%<,�y�_}>���^�T �Zg�N��`ز,]L��r��%�@��ȓV)��E�3��t"X���s�Q*k����.�rju�d��K6�5)|�vu��z�\U����L�ļ�����v�"3KR�[��P���u,c7�Y�����,���{����g�<�z�e�a��l��@D
�I9�-�����:w:���O7>�^ZyE	[��t�}�Fo�8b�#����R���X�.�|	��+1������O�u(]�dl�7F���gohCQ����rz豾�1���{WP�H��O|7�����;�/�D{�4AK8Q=-h����z0��H�$b�18F�D�7B�n���<X�/�,7E_X��m�ʻȌ�f�NP��q�?��Ψ�U�[�s-�w�H�c����&�������P�pTy~�L�$!���MO^^{0�{��s����i�~� �T��ɧ6E*��ż�qC�J<�r^���ҝ��m����Ź�3*A9���PAPtJ���/)H��3�΅��������"��4j�-Z���Փ�+��
�iR���ڹ���Bܶ*����򒼋C΃w�M��hyh"�b�d~#ց��L�u#��;z��T��t�����ˮۥ)˱A���x!<N
�^[LI���4)�!m�`��,����%]~�=.�|
p��xMs����6ޫ�2Q�����v�y}�	*Q"�D	P�>�T���=��g���N����E�e��G)S��QT�5���\����De=�a.��G���p	n"�b/o�����%@-�=�ǎSK\>F�4�����}� 6S��85�N6�G �(�ǻd���l4
e;�Y	ۯ�r�y��d�����M���� ��d��m�AQz\>ͭS�vq�����s�=�&���5\_��v��
�`[oã``5��ڳ�oQ��z98��j�F'԰��wg��O�0t��"Zݝ97���k��z�Hӝ�����#fT����;��(��P��1s��[K�݃}%ͫ��%��0��8%H�����
.:�>,�o)�y���z}59�b�M���a�,���)	Pڰ��g!\�3\{,�H�FQ~�۝*2�;7d�2���Ca�z�f	��ƻ�X0³@E����l1��f����� sik��ve�=$\{c�.=�5�K�}/�Fk���֪�sbq5�h+4HȳD��S�-���������6��59l*8�R�&��Ml�鵳w`��VmmFu�Ҫ��:J�C�u���-`�e����4�=�����'��Q����փ�WO�-��e�&ʫ�uuQ��gڊ��绢�Q��Z�-H���c��a}A����Ɋ��l?�ܩ�*��RC:���6�u��${YK���Y{W|r���^��4>b�Fi�t!Y까�D-��Pd���%�����HC�Z���8��ҭ���Mk�gt
� 9JN���A�`�͊��&��&Hvwj�j�Ul���V��p�ظ��U����}z�E���}�$p��Ay�J�K����S��l���]3�GY`��-��-�a��Vq.�2R�9��l�'WQ8d6c���:������`����2�)�`�n�}�T�4�p�]6����svc;T���!K��̪��>�q�����
�"OI�@v�W-��(+u��M����C�{��{��-�<������\�Q�"{��y,sN�}/\z��
ynz�`��c��q0�>���U��.���o�{����՞Ж$�X���z�(Jy�ַ�q��>R�
'uK��[�u�[Y�����K�� ��FbCr�Bi���?�;�
�2�g䘭tvEo%Ի�5��FLCt�6�H��"nR�;L<�f��a�FA��ܾ�5c�5r~��&��bc�7iޡy]B�'�m��D<x��.�����E$sK�U:��;[��<x���Lvx�I�2:��Ch�`I�*J��{�u�<��0m��K��tj�� ��Q��{�c�kCDAY��uYk7%�N4Q����+Dm��y�s;s/��#|Q8��V�<�.�m���ˇWɚ_dg���-CݥB*�}Yq|H��#��Z��"����n6wi�V�3�g��k ��=T�	�=@d�jK�k���x0Μ���v2GsH��Ociꊉs��v���foD,�	��Q��Q�� �P�<Ox���ˡ�I���k����3O�ny���E��G%��Tumh�q�7V����d���ox�'��t}��\Z�u���v���EzzC��rwx!ZM�2v�n"b֔�
׋�?#.����F�E�ir[K��e��[��3v͚���^�`Fb���z�M�:�j�ْ�,� y.O�OV�x �Du�κIYt���$��4�6 [�lZ���7?V����~|�r���dfXSlZ�ۮQ�s����K��V�����.�;!N���d�������O���G{eq��T�v�oouRV	#۫c|,���K$>	�G���b]L,�x/�ɑ9P��nj�w�6'$��3�w�O�3�6{e���z�T���¡=�;��o9�''�(�<�t�7�I�g��l�0q��������r���-�/s��1=��
ނ�rj�{�X���6z��k�9��ËN[&T���N,l����:�.2�7V��S@��N׳���a#��]^��ݵ?kgUn�p�X�E�u{bQv.2�4	�>��$���W8��IZo{Y�m�!d*�d
�P��ktk��mcw�1���.U��Kp?�#V�0�B�UO�����i�F]�F�'���|�K���g~�k��-;~�&���=�Y3}ļOx��>�$�*�����5:u�s/{%9X�
��o ��VңEn�ys �T�WIV1Q{�m�r����C%]��Q\�l���]a�� �
ӄ�"�1?F	"��e����7�""�A�s] s˙���i
M4�&��^c���4g-?v��=���l�{�VJ��OH����=ܛ쇼K/�mh���v�
��<{:y,�����2
�i��\ә�gB��m�@ƥ&v��s��v��lÙ�!캃't�{�X1�,��=L��ڹ��0���Te���v�]MجRL�2
��uL��Djm �덎Ar};�$���F��3v������h�n�dU7M5
㒐�BR��"=����RH��,�]�b7�K]�7q!�r��]���m85��೭�u�x؁�Wf��'���a��8lv$5�Xn�!f���[`5?�A��>�n�vv�¤�]9��%ǯ@���{��r�=&y�=������!X��Kn�y�Y�w��A�w�#�WPœ=ˢh�rt�y���A�����s�w9k���ʹ�ެd�i1@�D����K��+]u�3����⽶fn�)��T�p��̛<RD����*�����?� u��Pǜ�2
WgWi7�֙^.U�����Q��ደ\3F�3�b�9wrا5��O��U����|�qŦ����)��E�H�
���b2���R::��ܗP(���^�!̵��j��&�Z�&���8R����1�xO�j�2�/�P�[<��e�7�}:<Pr���|wٯ����6��L�Gy�F�}�"�ˠ��%�b�q[Y�K��f5�X�g�t�tQ�C]��w`G�M���]��T��f�v&��FWjt	���,o�t`�dtS�;/y�
�}+|�����ST�gW7�uEU�t�F��R��o+5X�쐅`��r5��Mݿ��8wH8www�>���DkD(X/}z�:�!��TQ���6�I����وwƛ���-u}�]���,A�n8F�()�Zr���ɺ����g������̛�~�
��uȃ�j�=��#P+^([�h�1/�1Qy6�~�C����4#2��}��M[8�\'�`������%~�S���B��ʺ�U�b[��;+2�WL��%�^���K�e��S]��v"]/b �]�	��lֻ�	ٷ���#�s��f���E���,�;(X��}Z�V��Sӳ���(�L	/xݗk�<�}���n^g��� ��mN傫u[�c��ys<iY=@�>֙��#X��3K
��[�>�ڄ�Է�X�$�{��|�#��Rt��hp��&[��R]����Z ��	�55�%v���%�<�8���5pĽ�6�j�����M���q��cz냭��B��δԖ��9�6�م��n;�4��c�L$�4)2��j�AW+U�W�n��/e��V16���7�l��˩9Y6�Z��6��M��	��¹᯽7�v�������s[����|Nón�"�_���{.6)��	]L��6��������3��ϐlH�=XiW[�Tt�S�tF�Gkvأ�&�u#�����m^t���M��q�h�NK������r�.�`�����2���^Ne��Dy:��.�;6��Ǖ·�\����9�%����V�R�U�ځ�t�w�dx �
�*_*�4�,v����t�	���6>ݫ��2�p�5��~K��H{V�<�����5)/
w{H�z<�K1\���G{ȍ��-!�9��g@�ɐ�r�wk�w/�3q�⹬Rzn��'�f>��%��5f��܇r��e�e»iv�7,�{y�#>ĽV�'oz-#�nW��d�����3K]8pmO�&f#}̚�u�e͋:lک�B.�$h�397��=�|h�/��i���m�h��b�u�[M7�.M��WD��G^���y�w�[r���7��R��nn��.cc}����%nQ㯕â�!Ղñ��M��nWEig7I>�UQ�x�#�Ӥ��$��ȳ]X΢�Œ*����X(dO_R�<�3ڑ�� 4cد�����N�f��JfgR�cr�f.t5��v�΅���ѵ�{<A˃���D��^3��K�:��������6��z%�Z�LB�B�7��)��̱����'&:�ViV�>]�ݝQ�j��䂶3X}p��0'�Q�<P�d|fX��k��ic�yo^�̩�"}������,f�QUܽ����MX�x ^�=y���"6�.�t�������/�1����mzs���j��汭Y}�t�%�6N�<pS�h�7���ؔ����b篪+/�y�x�������:S/n)75S�7�b?Gh}3[�9e�&�%�����c!.��y�Rz;u�X�cw6��%��e!M��]�0=+�9F	����b\����zv�եZ*kM�	��O7�K:)��f��;�m2�P��J�5����0-���� ��{�6�^؊1�l��:=�sK<��j����N����e��'r�_J˄^0�Ꜳ��|Ջ3U�`���X�\M=f[W�t��{�{�}|�oN��V跓5ԟL��k"VRe�u".�륽S��.���)�4-$I$	)@$IJ+C����&65kK0ml�M1����:q�u]�mA1����J�� ������cgSUQ>�͚���h�)1������ƫj���m�������AUT�`�%F���j*�F�f��4c�8r���(�����&�4jI��l�d�6Դ�b�h*��F�F�IynZ��=>��y�ƈ����M��E:ME�&*m�1I�YΫTF���j���3�8p�#�\k�UDEKk&�1E[j��bh�f�����b��4Q�QN====8r#�7�4�Q�N�����t�3E@E�4����V&��&q��zzp�W"���}ƪ"�u���ֱm��";�Ly�5ETM��`�z}==8r*"���jn�E7���8&qDǚ���b�6�e�l0�bѪ4b�����-��f���j�������EQ��E�0Eh�~A��j��~y�i��q�j���n��G\5�pU�CI��f]u̤�Y�|�;/����-���ZR3�^o���{�\�k����Ρ���%R���vv8�W�K�!��!��i�߮�f*ryi��kS��В�uƛd�'WP'�c�܆u�N�j����*3gH��(љ1�r�m'ݲT�\�2�𵭓�(��cKY�^�}�X�9N/��9W�
�Z`�]�{���ϫ���O��QI�a=d���#{��}پ�I���蟅���2>�x�F)�5�:;+y!7�%_4v	���j�n���1���$m0�`�< ��XB9p2�.���!����9=NzȢ'��wk�q��쁗��|�|Â���#� �*tfD�y���{O�P��_�R�S.�S�X6�Mg���9��3�P{.h��ؼ����~�Bj��7����o7$�x���=,ra�p�P¬�D������D�a�y�hftxf_<�VF�ffg����FD@�Ur�1������x�;Y�R{swj�vVq��+�)�>�#PX�n#b��NQ|V�3*�VӉɍgi���`'X�{}q�#s�8��\(x�?,�u5QyZ%�|�����v�Ϗ)�vJ���wU-�re��,����v��!�趧����Z���k�W3Yv���q0�L�x\��+�3;��f���+(ϵU��k�]����{r:��z��-�f�����-�	����ۄփ&Ԫ+��F�������@�I*)�-{h���e�Xyy���ۺ�2��$+��_I��Tv�}�Oǅ[@@��!�eX�7|�it��9/D_��gg�]$����~3�t�r�A�K��x��^T��j�X��8�.�(�#��O�a#|�%�R��I��q��Ě���]:��G��W9�p����U��Wn�����������C>�^Wͳ�wO{+�.+�����wZR���:�l�{�{a[n�����rv�׉�T��1��Ü0YN�\�)���Z�6�s�o"7(�9U��k�EJݟ+��a��A���e��h�4�{����UҦ������W
��a:j�x�I�78�k�N�zE�uV��>Ğ#eޞ`+U�"S�}�RW��׶�� u���kes���:�-��U}�6�Wbޫ�56ϴ�+�῟d�6�]����]�u;ꜺpN�'��C�i�`=KL8@{�8[/N��� =^��[�+�0rI����(��dl��������F*:f����љ��!7�b��uP�<��#@'�׹*7�pv,;.f�gl)e�{�d�5@j"Cz�3�*�����(����&x��s���Ю9�Ue`��@���A��t3��u%��6=�m��g�p]]Q�L���2��%��EF��O��%0�!��	�t��r�=�{�6��{DY��t����E�ε�1O g���)+縫L��l׵l�q�t�l�a�"r����sJ*��H+��%`��;Y)�?���T��?u�����a���{>��r��gy%BѱIO^��in�{��Ug��,��(K%�H"��t�����âa�ظr�B5�y+��,�#���/s��Ɯ�YW��������!(lDm��\��Ɇ�x���5�^I��j<��;8qK��	_xh�NP��)iD��.L�b&�^�x���y�T���f��*��42<�".�5m��q**^k��\��s�^pܯW���<��V�f������}*�[��N�_hm�O �����=T���b�����'�r~�;>'��?_O�������< .�Ю�m�sk�7t�g`�ᑸ���+��V1���v�I6d1m�qQ�p��p�=Ss�9O*��֧����/��飮D���Ѹؘl���3^z����;����XVKX��v������wd]>4�/&��5ꥏw˝匃pj�L��%�*ڥ7}C�.��s��7S�O�.�yOgu��d�r��G8C�8�d@ˁ���]�}
��ŻQ�O�+<��G�7U_g����(t���g9��#��h@W,�W�J��h������'�8�]L��쑽�'�Cn�1>;�"ΩC=O	inQWS�'.M���U����\4s�7���"N��b��ڇ������&�����F��lŶvC�t{*8^TP��瑚I��G�@�Z ��;bnAs]��PW�kGʚ�]�D�s����r�����;W��h���ף�l��|����`�O6W�i�Ѝ�Rv��+��������6�Cv�"�(U���vm���/����25\����(��{��O�<8S���J��;���I��{��y ��P�·W�0�?���ہ�!ֆ��s^3i�b�v=����m\��iM��z
�#~w.�����CQ�YP�Uw5P�C<�[��6�+��'2}sN�Pn
�M��d��";�֮���f��m���94��4j^Jz�#)�F�r5[��g��',*|�̸�&�f.���PRI��&��I7�Ue$UP��{LtW,�5z�V�u��뗀_��}�^t���q�C�5Ɨ��:1��j{��)�qO�x�ݒ3�
 }���n����*k�.An���� 53Gi�׵������k��r7�D-����N�s��UM���^��ގ�$F�I��k���C0l�Q�Ϣ1O�i��o���,n��f\��72Ks���(I^�*��6�g�� ��
9��~�,���A����B,������eb�H���k�����=�+&��P&�E�����2�J6����$M�іe��s�ko�Q`�HaI<�2!D}T(�*��$�yj�Ad�9�;�g|]�b�z%�w�%�jB˱�/5��j�E�u5��̥�5m�Z��b�V��2�>���gL�D=s����l9��?�'��?��P~�����	��ͩ���(�q���v%Ų��g�w�:��bC��k��,Z3���gg���pD�g�lL��ktlvY�����d�`��~jȔ��T�~ﹼ���w�2�@"�</2)�#��t��(��sW2v*b��D�1𕶫b�N�ρDH�Ϙ�ÚYq�D�;�-��ug�v�%=tlAZ�0�	�"�����)�hOc�<�S�&l�@�,�r�ޔ]wm�ʺ����A�jU�ƽ���3�΂��H�l�;��>mm_"խƳJ��-�+�Hɾa:��U�ד�4�Mq��}6tp�rĥ��ptX����-�r��^���j��%];�4��-Z�x�<���Eک�P�(��(���݂��+�)k��`�h�0�oɼ��b�S��؇%��Qt�r��۰��Y;��'T׮�t��j��ߨ�W>�$��
j�F�1�>�wwL\�3�V�X�\�J�r�w�e�b���ć��J�5�}�8���<�^�Nj`�ew<��}�9+s��J!�.�iю&�G���i$���1���j�Rc�FC���#clʡ�^=�%i�5�����]��G��ʣ�)�a�ӱ��iYV�AP����f:����B��{:�t�|��V��y�I���:����m�$�Pˍ���ΖBNv���@�����8q���r�[��n<5���O��ry����n��.�ф0���ozQsH���W+�A穻B�am{7*y�+�w!���EsX)��w����������~���%\�GF�)�]�Z-c|Z7;`%l�/��}��&�
�����E��@��|�s=��ѣ��wQV�n��c��û�Um���_�H�o5�ʾ܈�X.4Mk���3�Y���Wf�gN�F�݉��=���$w"�PHke"|{�M�f�Vc5,����&\;��k�Eq�v��t�^@��%�,zj��`-Jص�F�pa��&�wNK�'���#ouEL:e�饔%�;�ʰ�k��Bg챵-��K�<#�1�|�B���:'Ur���W@�ӈ�uR�-j�Y�dD�����|��;!�y���&��:R�(r����y_[�ßAUFU(�v����ׂT-A���X�Ĳ�i+y%Bє��m:��G�Ն��A]����
IߪR�
�pB�9$eD.�'�p��\��X8k�z/���2{�_aJ
{��M�S,M�n"2@���lDm�kƾ�^��TغY�$p�@��4zt�+�#[{�~�S�05���"�S�";�;L�K]��qt���wM��+�"��T����|�kp��8k��Ja�{w���vm+�jEឣ����4H�GU�J����kle�6�=�q����B��`�Dr����9:	F&�Y��O��P�����n��4V��ˣ����R�Il|�-��#fT�m�w%�Q5	ݺ6�h���1�����7Gё�2��o9СŃ�~��x:Չ�-��a,�..��P��g��Y��̵��~��{ڜ��{���d��-�O=D��5W��-*�Y~��k���A �?1T�"�D\�C_w;����c�Mf�$�n{�3"�B#�O�bx�<2N6��5h�%TLk��s]�(��N�N�ܪ�8�~��~�=0X�)�Z;�B-�fmsp�&8����a��_��a���\�c�ݒ7�gôWt����wz�� �1�r�.�r�ƨ�%�;9��f��X37-<�XDW��F�h�Z��s���;`FV���uèIѕ��7�,�=�\���&��$r-��*؅�P��� ~٫߸+
H;�v���\p��k�T�G/I��ćZ�Waٙ�:�n~̙���t��zb+(Ϯ��S`YB����d��d�D`LA��r�ux���^1�Z/���8���D��>�����Gp]�Md-ŷx�-��5����#b*��<1
䌪�fF���p�����\�v�5��:���w�^���K����s��ĪT�T\�p�0�O����TMV�b���\��0n^�	N�<�)X�\F��;�P����F4Q/����L��݅�zDBN�N3���lѤ��ޞ/ͱ���W�5%m���u�X�ͻ�x���.d��� � 0}� *�'�uwm�KfZ�`I���iY��g����հ���e���F����O��]��3���1Y� �Ԅ ��:�ݕ/�Ю|<$yН��!��tc��m<�T�\�̷1�f���c��ْ�D#۫an�}� ��E����>��(�f��o��9��s�gV�r6�`4DUp����m�א��y��\o���g5���4u�DY�=��
�'OQ�1%S�6�8���_@pQ���QK��Pc[Xx�F5X��]@���=��pvH͐۾��|a�42X�Mp���ϹzFt��h�.���"Dnd�t�%�����vC���":n�)S`�{�k�'�錋g3��յ�@n�쳅�ki�;��.��T�`oj�����6��St�/��%)y�k3����C�jxgZ��-����o8�H����;��[g^�f��|瀅{�hE�i�Y|=E��������(N�D� �"A��rd{��r��'$�^c�ҭnÁ������VRz�
+/`����A���=�ɛ������%��"�(/�"@��UL�@ $"(@�� (@��*�@
�P��? ���"�! � �  @  @� @��eM	  @ *� H��"�	  �  	 � "�� 7�  B� @�- P��P��%�4� ( l��"	� �a(�  ��% (��!@J@(J!� ��� ��
@�< ���P �HP��� �UB���U�� ((%(�M�4�J�
�� ,
 ��}��/��T����
��0�Օ����M����c����3���L��NgˀNo��-�p2��V�K����DQ[J

+�� u�C�8�|C�2wX�
+�i����i2 ��װ/x�O�	�i���w
 ��*0���C� P�Ъ� 	B 	J B�" ���A�� �  � " � 	� "P � �@ �D � 	�  �  � $� %� %%  P �UBXVRU��	H@��V@%a�ddU�f  H �`@�d`	 �dXBU��b V �bU�$FU�V@!U��
U�E`!��`���f�� ( � � �1�`<5�bq�܅G��s�P"
+��&d�fT'E��,n�X*b�*(���91g�/�DWW�� ,w�t������j�(��N�rPf�&�0�2q�\J[���r�
+��7���w"�
+sxm%!���כϼ'}�ϸu0�mBJ(�)Р���8>s�|�#pĚ�<�{l�׎����[*� ���;�͘�:���Xa��AEw��	3u���
+(����Q�3d:��1AY&SYkY�^4ـpP��3'� bF{�>@P !QER�@P%J�
�@  P U���)I*���@R�	"E ��'f��%!TUJ��RUP�E*��JB@���T�Q[���H�T���UBUH#�
�P$�H��ݪR�������
I(��)J��IA"��)u�PED�j�( ��%J���*�*�EI�P��UWZ**���  	���텶���[���b)wu�WUZSj��L�$!ʲ�w�lƻ�4펜��[6��J-Bˬ�\�%�fT�R��ۭr��t����RA)x   ��!�dhP���lP�T:ƋbEއؐ�CСB�i�Ua�P�w����Ӯ�q��Jv����j�l+e`���Uv���i��m��-�݁u�WdU*P�RPJ��   ��T=�p�eT)�v���I����9݁vu��4f���Cr��*�e�.;r��\�[v���q���۵�-m%n������띝�ԩTC��U@���  һMj������	;eۦut7[S��kcn��V��Y����T�3+*JSFU�D�Ӷ[�'m.1�R�RB�J��QR��2�|   �eE�jk뒶e�0EU]j:�[��V���(��U\�� �m˂�V�`��CV*��@P*� %U
�C�  �j�`�d�%�Y/��@��F֔)U����٪UїTL���zױ�ړ�0l�Ѧ�B$4U�H �R�B��   ��+eu�U}�:�E��P**z�]�%Z�[f�@�:\: P;�` ��`P: �:
Pt0:)F��I$�
����*��   !�(�Z  �` (P�  @���,� �0  I� �� 3)�U���$B""�kR�$Q/   �s�  ��U� t  6۫�� ���� vK ���  ��( ��r��]� �%*� Q$IJ_  3��4Z0�Mj�N� �  c t .�  7B�h:����� ��S�T�F�di�M��
RUA� U?��M5U� )� ��@  Sh�*H� h�eH������f����~^~H��~Y�k�?7��K�Y.m�hA#�jvϪ���3�=�F/ <<=�Vu�>�cm�������v0�����co�1�v�6������<���$?Ѳ�;taCFԷ�n�o%X�bVX�� �76������_�f��@�E�8�- �׆�sqК�n��2�pE��y�Q'f܄a:����q�H��qe���4��U��{ �7xU�B�իSQf;����S]�G17�[�㆘׶�V���a�I�0�h�/SY�.��Ӧ�bʂ�*���;�5c�Sʩm&i�"��;���X�ikE�����`�Zɗ%�[�2oDa���W�*om�Ѡچj�̄�W*�hӛ[O�2� �X�塚k����
d�U�Vl��K�5m�,���P̢PQ^ԺyJ��a&�$8�����n2�j�A���v��Ö�d�fk1XA^+��6��Ն�-Z�^���������l$�4��,n�h��[W���%�pn^7[�RfABKB� �ѭ�z�%�]
�b1����� Rl3sl��	Ռ=q�r���C�e-v7V�`{M\��6t����y�!�Tͩ��m���wd�N6���L1QU֕0�sv� �Ŵ��K���N�w�7yO2��ڳbUw6���j����[����[�	VRY+q�m��u� �U���sWj��ߡ��c�ӫW.�(��w��m�vV��[��/Z���%a٣%��31����d�!��5�C&�wX�!�$o6��%��#��ѧ�/���ؽ��,�@�tBlÁ+�
v2�'�m��-mͽSvV+��ȪB�l��pէz�3�K5�ϖwlv�p�7�sh�lQ�u���"h��^�Z�+tp�e���֑g#������ON<c>}[�ls(v�H4]�k(uڬn��0��7���N�.����Օ�.��wEV5a�@?�*{���uoRX>g�vw�lX�R����eJ�9��G��&�V���A�-e�����0�.�0nm,�N�*d4�S�$C�n��.8p:�uc���p:X�tR�?Z]��:��O��VH�\J�v�J�U��f|��r1p�b�X:,�n�P�5܊���tS���	a�X�(=9���ھy|�v�A�-]k�d�%$�;�F�1���X�,�r�M�3E��T,R4]�@�w�������������Yk�8�;�a��ͼå�a�.WA�qb�DO�V%YZj�=tj��uݍ�)R�l��M�\�
�I���M����ȁ3u%4��le2��,��u	T��r]`u������Sq�!7��"�Ș`7k����ϲ�9�P*]`̤1ݪ�P�B�b�a�����:[j���t67�>rM������;��+7,!uܚr�F�l�z7Z� m ��dOj��0�4�˘�ѳ�&Ͱ�.�ƣf'n�4�amA�na-����j]&o-#>�)�e�5)�N[fE�n�I74�E���T8���x/^�e%E�[%��bm	�ie^�Ӂ�4l�v������T�C���I�[�w�U�yQ�ڰR��B�Ի�AG��8���j�d�ڸ��i�ՠB;�7��j���;@-Y�N�9�NJ���5���b��ǀ�d䐌�X��Ggn��ٲ���T�F[������2��{+����M��]�3��e
�y74��1�L*�e��Ii�h�� L9���l�ˢ�>�*�*�V0=2D�ͬ���P2s@�
�ͣF�3*5�D�]#M��/iS�já��emj�kn�2�K�ϓKݣ�O9.���0��Р�wǫ�÷�cU��m��JF����Yɣ�.vhc�v���syvV^��&�PSB�����,w�
���tsŌ#��������T�
�Ӫ����z��u�e���/3%��Pʓ#�5�U�vw��mm24��|������(����25^�2Y��%���gὧ��[������6[n��<���-#����,�wr�o��Y]�\��l��ˇ+(�����Z nƯ��bΜ_Cim�So�F�b𐝍�Q�̢
���6��䴺�WD�<�gZ�yd[�����Vm��Z`��P���&Bظ������r��;�Ǘ�U�7L"��
�dQL#$[�;�Z��N}7[ f)N��p�ڎ�`K.SiA @m���Ij�:�m�#�R�s4�mfh�WejI>�&�i�t[�u_-�e��(���V\C �$[���a���.�+��e>]4�u�:(A3ȼAY�����g���r�n��t}��1�i���6�X� �wJ�*,�oQ��F�4%x�/)��r���o�lw�n��1ij�R������[F�T�بq����"��=�A7���[z)2��^�������R��ۗonn��г.[7)�L-���U�kFz�Z9J�ڇji�6�ZȠ/J�d�^ݨHSO$�J��]���*ё^�Yˡ�i�kF��=�ku�s]�=U��T)P���l*v���NaW����sp+*�葩-n�拫GCBGk�WtՊװ��f�,�,e	��u�,2��w-�N�O�f�Bl0r�-M��ӷ�'Y.dէ�Y�H�ݬ
��(=Q�b`[z�=f�.v�|Ƽ�8���C�r��4�iT�X`щ<@e��9�������\�Ք��Yv .���!�CBBؠ&Y�&]iqe�DR����kl����ͻ���}���m�Ab�S�
"��{��J�[�5D��ߙܤ�c��H6Т�az���m�h����[)��n��B�<(,wO�]�����m%W����c1R�P��rP�0)�3 �R����fZ�b�7Lmh[w��x�+��ӵ{35*nX���f	��.��M��ʹ�P��2F��b��2���#`c-��a������.���%����kr�Z~��;s1��T�s�L+$#Fjݹ�G�]�z�謰4�.�,��ѭy�/��P\HLdcm��kei��_ig&���k���e�g���ͭ�kAS7K"0.����;�eq��u6�� `�L�S̎���X��v��eb&�;���	5��b��$o+4^���t�f�545�`4�nQ��jpP��^3u��Z1��n��Pn5h^*W��-͛�n�X��3<{[t���nZ��%ආ�q
���Vl�����������o ̫`�3���CŁ��bx)3y��;Bl�a �0��5�]��N�m;��+v��ƝG�*8-�MY��������9Y���#��[�Jb[�1A{�T�{*d��Ju�ж�M
�p=9�Z(�wu&���d��1[qK�Lnc3]
x�Y�U�t��,�jȡ��M�Ӯ�0�6@.�?ESsMXY� �i,�njPج�����k��U���3F��j˽
H^�Ɖ;��SK���so^4uha!�m�bԫWIiR�$�����c�����]���tt����	j��b ��Sij����hlZ!F����Xѹ	�pDڵLbҞ��QZ�5���RhyYu��˥�t޳ �kqmFl��˧����`�P���H�1fb��	��9w0=TNU���Ι34��8�m�&�y�F��Y�䴕+�O��v�"�a�D��w[q�co t�+�AX�g[B��ۉ-X��m����I�1{�u(2�)��[���65V�,S�Wc}�J6Q�R6\Җ�S���?MU�I5�[xw~>B�	��u��:��i�M�!G3V~����Ť
6�7v�س뛎4�U9G+@��̭����]uzsVOk���$V�-�-/I���fD�&������bA��r�H�,e-�Qּ;-X���k��n�X�5輠�ּ�ͫ�H�ޛZn)-4+0���V@kӂ*�ͷKU+f���m�T�1�9�m!�ŭ�ͬa<�[T_a�O@��YW��ӣ��3cK.� ���`Qkq�[l��4��*$;U�by�0���9�hڕv��VpG���^;�V�g�e������OEg����m��tot�	�G"�s��ƍX��*3$.K���k_�c�%mf�7� ݪ�I��t��A+	�v�I�R]e�c!����hL��5�I�̷�"XjΗt�]"-,�S�� ���`QS+I6�fc�6��ob�hl����͗k,�-���,U+7(SdRx��Y��mP�M�T�^��.n�,1���r��0�׷b��&��.�������sn����jl�����yQn�k����X�(��V.�2�^��b��JXh�q��˙-�H3����9�t��7M/����J�9�F�Gn�7���Yk�|�in������h�y[e=�d�-�܊�e6k%�8�Qϱ-�a4��Kj��!z��n�F�j����ސ:,	�F�rw2�&����-����B��i%�6�2�{�� �z��G�[�j##B�[����%ҧz�����KcX$����K�N�Z��#Գj�x��-�p�f�:F��N
�JW���g$�q��h�x���YRc{-����G�rh�Q�R�U���N9d�H����x޻�V�
�{�v�lB�����V[�
��on\ϱ=#S�X;���0����ܾ�0f�.��3F�A�݃�ϓ���{%��	٪N^Yu2�݁�� �-�/i������:/��c[촘ϯ�m�#:�����zF�O�yA�G	�x�,��z�����`Ċ�t.�2�C�Xçu�i��ݜG&c¡J����↮���l�� ���3r�v�P��Ǒ1V��shh���y��t��-�DV|�m`�jm���/\����ɘ��t��zkE�n��oKN,LՏ��\$o~[2�kES�������O�`{Ƀ{oR�hࣦb���b{6T Y�H�5�\��%�L�����r��n�/v�d��m u��uWm����- s���ZǪ���c��6��/Bۙa�� ��P��+,�#V Y(�K.����ں�Ļ�"�IaE�7��i�<k�%��]$N���η���V�T�Qt�{h��d�$���)�-�K�b�(o-�6��P�B���?�-�f�G��l#}�w	J�p|Ͷ7xq�yV�����9�"iP�B@)���6�*t�4�ge.�%=}����awd^6���yZ���d�8$��x��K֞�Ќ1�80�Wj�Y˛)B�˥Xf�F)n�+th����m�	���s�7A�w�NQ�ud�d+�k)�x3A��15R�i2�鎮E ���_f�(�.�2�d�X�]��n�/v�*	r�����N$�$Q���[��F���8�Ɏ]�2i��$N�iK2Qga-R7�dR\"�{�33l��׈�T��٠"�N����
cTX����R�َ�oV.�]��)����u���iAR��
�,6�����b;X.�Y����һ�5{�4Nf������1��7oZܰ��G� c��op����#q#|I)jgu��Wī��x2�u����|E�"�^�ŀ틫�k^��e��D(�L��e5&�ܸr�ER�Z�i�D�l"�0e+Z��@�{b�� N]%W)�X�ot-T�܎�˚kAף@]��2c�t$s^��Ҡ��ۀ��؝�p�L��f�ugXm��D�[�vJ� �b�u=�7R�W���Ch�� Z����j� ze��<�jL�*%���Sx��Z��s��u�@����Ӷ��W���>y��3H�E�������2��Uq#�%��h�$(lͫ�le;.�Q�5+�Z��1�w6X�)q
n�P��LW�vR����}�PIn�&��N��Ǻ�Z��1a�t2`ِ�,��Q�0�O��X��yb�%-{�,�n������qn�I,�ucMǨ���;����+`2���n%u/Xe��c)ʵj�!�z����c-�;���E��{spL���"JgJ�����tQ{W�&���(h�,���Y�7kQcx�tP�:�=<�V�|�夫q̽Y�eҥc�S�~���r�:�ʆ̢^���
Rj2�e;�r����j����Y�⎑Y�Y&Eҩi:�C1�v��[{�a��N���	V���W�
�ޢ(�;烝�$��r�/�X��;��4�j�GHen>�ʃW9R��t���^f��*h5Y�d&0"IR�]Ku�V�BL�s|���2@�}l�u��5��G(��'&�޷Gr�b7�VhڳZM���H���+Z��P)���l��M��Qf�*bWp�m�E�+3�&b�J.m����ٿ`)�� 0���dZ3Q�[�զ�ɭRb�6�;�)!�f��է1�� !�{�k���l��7nH!Wt�6���6aY���o#n��|+3⤇XU$��k4=ԋ���-gN�Hbe�/.�+���0����RF���3����3^�� �����ח�:�y+ue������Y�d�w���Q�)��Ʊ�h��wzk���Ҥ��#�vhT�E�KB��!V�c��d���u�V�=���J������j�7KA1D5��3��JVw*GCsM��pX��${[�2��Y[5���r#��CV$*4AW��m�k4`�̡���N���V<��t/鄉����	+m0^1���ެ%��WjU��eJkMew����*&^M�"�&,�+�/JW�)>���͒]f��P�h�7%��oe��65Qz��1]��eL��ʀ�P�-M�b �W	U6�L�YԖn�e��IB2ĨPU���×BnZI�T1����B=�WI�$M�\�d�*Ij%�ӊ�4���j�U�c2!N����H��ݵ����Y��ܽ�p��N�x�׳\h����R$H�5-�,�B�ѷ�m^ӭk�Ė�)�=v%٦�3�U����˽5��F�X���C@V��%]Ԗ<__9���_�r��3$�ာUG;n�������KǑ\9�q8j��E�|�HS�e�Gk�8$��,�m��r��jҝ�(>0�����pQ�/j�)�-J�IvHwZa��﬌����
˳�z� �6�<�Ky��.҄��Dw�P�4d8/�����W6��֙�CI��33SV^d���;VoE�2pc2��X�$+�I��T̶�.��r8K}F�I:�`)j�)�������|�`l
[7*o
,�#3��g��WE��y�	0�Me�Ý�bQq�o� q�s]���e����l|������l���x�Yw�u���6l�jJzv�0��]���`�Z����]Yx��زč2We��e�;�+�(���y�'ʽܮ-^��#+qGhݷ��ͤ��]�2�P%o��wu�>���}�a�\=vh�@i:Ju:� ��y�;Qw�Ӹ%-��<����d2���nE�j��w C\���S�Pq�p$�K�G�8�E�nV��Aui�w]S��T�8Ӿ�������c�'��� ��%��5	� �0���f�]���D�����p��KI�HcS����['v�y�,6����T�5�R�Ǘ��͉SÐw�G��wP�F����u)od��:S��5&wη47����g&&��]$)r'�MwJ��S��X� `(u�B�)tj��F1����D\ww�� 滬���g�Ǵ��٫2��GA嚛��'�[�q�4ԯ-�ޚ��{�4]��#^�����wsx^%؉��FZ�},���8e�S��f��� �ҷl�L��k[��N���U�V:�Zn��eĒ�+�MuE���*�luZ�((iuv8,Jr��-p�el�m����]n���Y�-�Di ���o*ґ�wv󊻭kk�j�r�er�!�>L�^s����ɽ�n�����y[I��h��>df��@�iZ���!�p���E��s�,P5���b82��ʙ>:��eGBֈ��p\O�Rn�a�Wz�H=�3��
�оt5�WcT��t
q`-Em���fh0,�·�um�;BP��6�o abp��Q�Ł��
����\5�t�gR�)�dX7$9]��jhc�xe����3Vt4��r��,mu���՟������u�Z�p|;q���^Y��v��:�gwg�A7���'�!��n̊��ʡK]��V��[*�
%e[����ֶ�ۢ����n�t$.e�E!��DtxX	1�p>U���Xb����-�?�xR:��w�oq7ՆP�����%�6>�r��W*����`i�1S*=ɖ�y#��&�Y����ݽwâ5x�����?<��ru���T�f{/ ��3o+�C���QoM�e��u���
r��2ۻ�dx ��l}��Ë��'vWv�_`&�,Rx𞙻�o:9��:\]jG)��;�� 8�!|+x���Zaf�����`��9�#z%<�8���Wu>S�T�f���v�ˋ��rs�B�W|�1zEJ���E���(������9��Z��A4r:�E�v�:�Fn�7��u�m�����pz6� �a�-[s$s�aR��D�㕚�u�s6�0k)4&h�ov�kZhVH�m\���J�d<ru��"	a�Blyw��� >�\+Duwr��hw:՛nB�dvZ�d"R�ӯxK{�4�]9�&w\_m���0�sv;�z�Dii��83;��bB�oT۲���77.�F�6]���j�)�ӕ����L�i�ۣ�^�ݰ�$����L`EU����&����4A͙
���NL�
�L�9\��0�|����sý�.���ǎ�׌)���W�|�ڮ�X䲺dl�nVL[�Q�EF,�eu��߶6��jN��+������}cv�&mZR��;ՙ²\*����*�J<kCF�dËa�ѣ���I�Gh�����Z���Y��Fr�kEZ<Gi%������R�d����fv�(G�K��+��X-u��֮1݉!S0����Ê��V��d�m������j�W�gZ_	��Β�)+.�M�F=!��Y{���P2�x7��#A�sC��t��V=��؋ʮ�{@��jkp��q8�a�����Qvj����8I��9���e�h,��v��3A�5�ۅ:i���S'�'W#	�5���_	���I�ذ�1쮾�D7�\<��+bJ�:�6����_!��Ԗ�|ν�5d8�T�ow빙b�(p��Y�X�����(	�fc;�F,<��O���='$G*�+}��3���[����-R�:c��GIS�Ե
v�+j�b���r���l7Et/M�c���Ӡ3�^T9�!6�)��sH�RXo�) ��ݐ��oB��!�����d=��Xe�^n��频��gEZ�W]�Xq'xɧ�Q[=J�`D'f�+G/���:Ȼab{}��G$���
wۺj��O�U���8TMX�7�Y	�.���Ej|u��L
�F�A
]��ۮ�l�X�����a��8��̟L�-E�V�ȵ�{�[�/�Y2W(c�YǼ��|�j����s~46�qP!"ř*yK�ye�N��Zf��z!�^Tc}�Qk2�2I��=�´��Ϋ�ݫ�n�����}s���:���c�0]m�� ����ek䩶\}��w"�ٟٚ+�]RnKܡ{u2���`vB͎���po>��r}�ꙇ�yP�I\��c������/L��\=f�B��m��:��ΚZx��U(�ͮyW2�'H�������׵�s�W��[J>M|s�x�� ����bj����u���:�IZ���cٴa4�`rݳ���X.�j;��N+T�r�m9K��?v��ب��p/-J�LTp,����ұ��h���r���k�R�О=�9mdWL�N��u�_�*��Z�Mr�iu�-��!�u2$p>��LS"�i�g�늜�������ef7n��H��b6���Ygx>��4B���U
[���oXS������/����T�N�m��[m4�<�ed[�7p��@RZ��f��T�po��*dbL��Hr$;/I�h>K�-��z:�A�ܬ�bŚ��V�Qi�J������M�uua^w��@�ILtn���ÐL�pߞ$=��X��K��3u�\J�������[ŏ(bI�)�yy���+����4�<����\$����FFҼ�綬� ����]ݴFs7ąĞkk>µ:<��sVt�nN��`���Y�8�ѵj�C��R�r������n���U	Z���=�ۥ6��,R!X�V�m�(�ɷ̑�G9o ��R��{j���(�A�nu;��xM��P2e�-Q�TL�*V���/��y@y�x��������Fb�=�e�]���[T��]n�<�m��=У/^V�K��7�.T��k�Jk��ϩ ڻ�Hv�j}�����WESw�xq��{ë�P��(�a�2��]�{>L4��Jj���e����Y��ܖ��d;C_^�y�Ό��;-�����{���\���+)\7��ǻ(�ٙ7�35*8'o�I��E��[�sj��V�\t��+����̥-���y�V%�ܢt;b:�EHL�
�-],"ۻ���S�͛Xn0��f�[ѵ��G�ɱ�R3F�#Y�!*wAǬu_T���ݛ�nVhN��۠Ug�i��
g�U#��6�]�15��a�v��)*e�s�,���\C�0��'�k�t������} \�{�	k5�W@n��$P��{2!���4n�k$�1l��匣�܂�/�=7ڍ�.ئ�m޹Y�m�y`��j�u��}f��-�8���f.n��w4Fe����|d����(l�MJ�u���{|��f�O�Ǵ]�
�,��v���G�n�<�w���'WIS�YX;%��(jdt��F����X	�Y��_��;�	G��ګ=m��Ԣ[���kr���˧���|av�Qh$��.[��kw��	Ƶ��z�����9��^;'-P}�X��(���g�f�]�ZzZ��ū&��wYWaJ�9�C�E���*�4�d�Qr���K}M9�u��s���_XǓ�t��֓����w�;�r�5���\�Q2�������Gq�w`m�7>S6Ŭ��j�Ҙ��t�ײf<
�fc:#����/g7B�����Hwo4Z�g$r�1)��[\.g%hDά�.����>�i�GVv�4�C�TJ��Suf��.���]�1���L4;2���.�����Zȫ�Ů����t\��X�< ���7��of�RˊMFP.Kƃz�(V�.�v���-��Rs�]NA[���5�Ԥ�����0n=Y��@��Tܻp�t�܋���K�i�tw���$��J�̙�|�T.k�y3�k
|�r�h��X�Tk:Y�B��r)4LZv��+}�m-�C�ۋ%�-p�Na��q�7�0e<�.�i�����W�0ҩ�B��VP�n�|���wn,���7�e區K�����xԲa���R�Ҭ�	�Ra��+J;ζ��O{G<��\og�\.t�yQ���N�Wh��h��ҥȡR�����C��O����VP�4�0i9Tݭe<'Mr�ʎU�CJ�U�ZL�$ۀ��Kɍ��'��f �����n���u�Wk�]��nZ���[4W*MH�3丽�a`����@oO���p����"�.t�Qa\:��6s�M`��@�����D��JF�[��t��hėY�׹Y��NL}�8HGn�& �WP��j�]�3�e/�=�^]��Uް�J�s�yb/&�
R�U��V:�w=A��MD3����'��Z�>�\#h�[��}��ή��\z�q����3���*��#�7�&T�G�0���:�+1ݝ|52�4����'c OO,n��1>L#k���*"��7��9�8lʹ�D��6���d=ݼ��s��OWJ��3zK�eZx�`vOI����vH�c]9S@�Kk6�g��6r���zT.��B���D��wa܆
�ÜЮ�t_[�2�̙O��>NWQ̨�:�e�������8r��-V�1]k*�	��uo*�v�[5�JF����D�;wSVa�8�Z{�f��R�Wō�;�݊W�x�!�����̣NΚ����8I���Wsn�pƣ�s0�B�
%F�W!�.�'j�c�.�������&�Y�$3J� esxh�sybF����}\��e
�� =��	�����$c�&�F���*fv��^ T�J#�#|i��p�V*Й��Բ��P�ۗ�5LR���!�/I�}��]ɀ�ս��eI�oD��2b�ҭ�����M��f�ѷ�Vc�E�y�FTܫ�T�-����|�� T�#��M:$[�Q��7m����)Ú����7�;V����Y��v��2�,:���$;�Ioe�Ip��Y��+��ݍtʡF��8�p;J���������m{�����%�p�F�u(������=���Ʉ*�}b����Q��8������0�&���D�#���)+cX"�:�G��h�6�l"�V���:ƛ�լ���k�c�K��޷[�h\�>�"}�����6�|�J�
upw���4�K�s�=�&���V��~�C0e%��S=4՞��Z/!�ǯ�H��w�@Ϣ휡.�����
Q���Kd��5o;:�͇K�V�Z����bx.��6X�ee[�-�[�ô�v���G���n�Fu��j��T7�0�Re�U3��7D4GQ�.�םdJD��Ω�#�k9i�8+I1��w �M��8Z*����kq�e�8�ۭ��n�x�:�'!�klWF��r�ڗk���.�,��]v�=�S��$�#`��".�O.� v� �����[��0�Ɣ�o�e��Y�6��}��fТ��I�ڕt��W�z�Ћ�JԂ�6T.��wd����M�E.��<�Jp-��#f�������;���li����H�0�a�ܻ3���w�j��oX�-T���dH]�@U�#shZ6㘒E��[+3u��Y����{�%�Gr�������s;SWab�`�:k����g�1��H��U��qMS |�V�8��fac�sJ�V��3&��t�n=	��E*7�CMS����΄���h�T��Z�(R������z�v����9Kji�HВii�u���70�9�H����y��SP��2풍� ��û���:�cd�"%��١0m;ƽV�k��]�ugq4�wG9�!V��BvCǤxIHڨ��l����ʌ��aٰ#�n�Y�RWj<E�0��Չ�5��r�6(�}s�\�x�K�����W���(Nf.\3���N���Rw(d��aIh�cF`����"��Vͣ#���s0ڡS����}���@ё��g]	�-j�놓T���c{>�+6T�+���
�j�g�&Y��|9!є���X��U�B�tS͡��.L��hgq!�G�*���'j���20���	{�����u�+(J`�G�H�Y��Et�3�����7Xoq,4�X�6�Akv+����;��}/h�� ��}]g�8�J���Cf����tK}U�v�3-�9�e��I�TU��3M�Wu]�P�΃�P[�f-D��B���[��[oM��̦.��єne�KD�L�d�]`�7o�->r��I����cH.��3��a�W	�&�B��^P�r�=R	��ПS	��)J!�Z�F�/,Ks�;"w�'L�ND5��w(�N^f�\��u��r	2֒T�{�E�%(Ps�9�R9�Z�諭�ﾯ�?������{Lv8����F��Vkt�o�t:�m].�љܕw0�p���4��>�ݗ�ֽQR���� �.��CYu7\��r^m>lm5�����[lΚ�o������Xj*9� /pv����m�[�ms"^��X�m�uqA\�Zӟ#� ->��e���o�s9xWN9*rs��̹u�`��+�xn7 ��q'���XV�K�Q&��v����
�r��wD�%6��]b�?���v!���s)`��E�yG��b°�������U��C�2�w^�*;���fQ�IS$}kI3}�R�#�yKs�30���JR�Y�qѺ7๕oe�M�;;@��i��<�>��5\��}"�|�+��LZ4�Nܭ&�{S�A�g��'sP��P���C��B�q���_b��h#�h3� Ƥ� s�h��1m�|��K�c[z�>�%�/�*d<Fh{���ףY�8$Z�u*Z&�庯pÃY�Ǹ v���Ү-��u|�@��{�A��^��]Qj�OpED� �CC1��'�^��tbv�W!�|
�49i6tDK����Ҷ�H�}
foYm�n��ŕK8#z��Y��t��n�sd�l���c��k��7��.�-Va�˧Pӑ#�Լ�.J��Lv��YcSOs#�f��&K��J�����K�Y��4�xB{J�u�*�rﶦ��fm�2q.��5��E�k��U�6a7D�B�i�KO2�����"4b��]�d���@�mvF���5���Rn�좁�6���Ҵ3i�Y�3����{�a�!�vy�J�8u^�M�l�.��B�	?d��R�U�c���soO^â]�^<p��Ŷ�	�b\ ��<���Z�ad�����T�t��<�u惴���:z�_^��رg\n-�����,��ڱ\����]p�`F��,�\�C����
r�)v�����`�S�&e���)�=�Rx�GTH\K�:�Vfv�����Γa�6ݕ�OU=�!t[��8R�QІ�^m�IZ:
��9��+f��*�PX��c�6[OqC-4��%v���o�T��;�Qw7u�B�;���bj��͝6��w���Vc�E��5����I��ڇ#��<Y����VvP�&Nr��V$fQt@�:w�r��Z/laS���_Gf_ߦq��&Oj)ύp�7Gz�+ښ+/�[F�ȕ�P�u�٫�5�XH7Q�®�l�CS��3m)�Q���W�%�����6օWF�\p6��M˴{�rma����~�9�h�t����̦sF�	��yEM�
;{;��9i�o��;��ݢ���:�[9F�M�qk���7�^}ֺ�H�b���'ʱ�*����"�}|F��5|{�M4�O��Y�7��cˌ��]j/���'���l�ͫ�LN�Zo:�F�t!��n��n�F:%+E^��^S���H��H7�t�G.�ۣ7��S��,��Yg��C�we��o��p)���f�4��̳ui<]�ҫ�-3J��6�w��jmh�Ӕ`�_q����F�U.��'n��W�M�ƛtŉ�MУǝB�N!<۶����J��`�=w�=�d�h��}��2f�c��4�/5��j��Jnm�t����C����}��z��AL�]7\��[�!�"�Y�q�ѷ�>Z�%Ŵ��Wmލ�ȌS�����1����G4�i�gZ9V����ɔ�8�*�]6=��z��q
:���w-�?7t�u��/1�V�'Z��tu�lV�m����>�VC=�]����o\��,��Z�-ٵY�0�u�tt+k7.�[B�E):s�<�'�6adˬ�a���a�GJ�����+-g��,ݥ��æ�*z{��Up���(�7}���P��݆^��Χn�2���ZF�3�X妶�<',�E�v#�����8��`&��Cc�	��'kjV�*�u��W6Qb����lZ�XhU�Zm��t'wr�k.em�k��3`�i��/-.�ԡ,0�.������r���*����
y���#��9:�5�v���C�<S{��Uv�6)�c�ps���Yw����o4���[ 9[`P9d��v-��e�Lp�N�u�̝�f����k�v�*�U>�[$������R�ls7f��c��P@<�j�y��D���n��)Pk*j��]d0R9���L�����5:l�}[{϶�%®�U������6`����Wq��]%X
�/�VI/��,�����oN�%(��9˷gP�C���Q����ܝ�M=�w-2�Zv�����b�KdVmںYC��u-�U��k
��Hq�a�C��.�s����M��Β̻�*�W۸�a�\��"�i��qPZw�{����#d&�F��S?g-Y�QOw:����,�B�TE;RGKuƶ�Uۮ���[������>q��@�����0pc���s�Sx���9�g]ne�w&��7�|�'Z��[��u�����M�}K�����6l�k2u���P#D�K�N5v�`�l��Z\uw:�g���� Ԫ���P�nu^G+Dj��ec������ޓdCX@wh��]�b�T�,�v���p��r!��5�c�e��nD���4�آ3T����S����tW>�aҥ����ӛ��s���[��*y*s��m�|r�2�]��i\@tl^5�l�o�	�ѣ�pU�U��B�v�z]�4u!�
��zfņ+_hV��Ӫ���R�9K�����i�Gr�������ۜ,Ŗ(�-�up嫝� �i�hJ��]ݼ��m�Q�9���p���嚗��b��%u�YW+�c*��SHN��^2)��n��(�a\�f-[�����:���!�fM�J�MRス�����^��:t>����;|W_t%ޢ+(��k�)G\�P2�v��b�[G.��[� ?$o9��{�z2-��0)ܵ+zV5���[`�w�2�	�70Ѣ�b��W++bvE����V�ޭ�G�����2�l���r�j�g'��:2�����݅�m��=6I7K ��_Y�;�"�QY �,��X7k��qv�ѬjN��uf
Qm^m�@����Gv�M�W[߇_n F��I܁�fӚz����7X�Ǫ�T�EXY�,ҽqлfT�-3;Ψ��3���gd����_^��F��8튇���z\Ń���yb_Yɔ)̍�L��Dg+�z�/Ǎ��S���NJ+��o4�XNS��0��S�*
��Ձ�P��b��mL/����;��r��x20H���<{QS�ٷ���)���{/-)��f�Z�d�VU��pz�r��p=���˘��͍�Z�m�ϙ��(.w
3
Y�7e�tu���'
�8̺;�"1fZ9��fLM���P�c{u��$�ld)�u���N�кv!R��=��&�p)��Z!���vA\kV8'J�F�mK�CL, :���j��f�ݠ���Y�(n-���U�5c��V���P�9��v���Je!z0]�]��5AU����Zq��s�ۥ��@_M|w(Y��tĦ��M���-M��]Y�%4C��nR���T�7tJz��i<y�!
�ޭ��#Σ��7��;((RN����̋M��hʒ�%$�ni��� ׼����wũ4�eu[VJֵ����wĹ�qڕ9�' d���b�W2_s =�.�@ǖ5]�1X�����Ec�\ê��cu��ڥ3
��-��)�AY����8vՌn���cN��Wz'a�L�ـ�����3d:�Q�0ov�5ZЄp���y�,�jU�m���Z{�n,n��P$A�;�;+Mm��.�]!�ڲ<^TUfS$����Uٝ*�)�"��V��t8A��b.l��
�j����M�]��W'=��fd*�2���j�ڊ"�E{qo)vE�՗>=3��!�F|��
�S�u��tw^e�zw��ؚ���@�@��9�e�̳�7�+d�9�^��V�%�t⻷wy�5�b����RA����N���Օn���b�!��e�1J�"�%-x@-c]݊���s�D;z���w"0BCN�z"k�䌭��m�.�i����2��0�ޤ�N-�oe�rtr��|9��`o����$@�z1�c^��%7/Lp�"��Ad+)��wx��V���r�cȌ�Y�����Ï�;nfjڦ1
$�7*�LL�����{-YWv^bD�7-���ƔDr��+��y]j���d������oRZ!KSդ=#L�ii�e4� �[ʥ�����ʇ:�f���v��F*e��@刅]��5��8�¦���d�,o[�w�Մg|:�ǖG�?����/Z(��y�%���K�P;�d�\����7b33���|.�4�*�k���=-��L�wGB.�Q�t�s%_Tf�v�ԁpX��'��r�fn����� Lg�m٬ʙ�W����{�Y�[��>��v˷eѢdS����C���J�X��(�S�1�B��{���u��'eVB�h�3m^?�*X �;�/3��A��\��73�	ש����]��n���㻑�n��i6q3b�^KU�.�ʭ�#w�v�Y�toJ����VA����:]���F�t�賎V	$�S��}�������X��XK���������c�9��U��:���oU�4\J�0	\F���+�q��`��ֲ��ہ�۵Y�e>C����s�f�*c\xW]�v�Yk���;'��BWMg���d)�Y�w�zKcy�m�����;��ӟ=��\���v�$*v�����u��W�Ʃjǜ�p�րE��rւDv�y{���	��^�e��u�\�Td�S[|.,J�f��Pzm˾��!ƕ�x�	IԼ͛��}� PẺ9N�X����D9�CzJޥ��Z���&�'6vj{1�6�ͭ���L�����\�!}�ɝ�k�V�wCbੁ,�Z_`�Wy�7X�p����7�(��!�s�@a�[�=^Ի�>�y�9y��of]�;s�G������B��R��ޕ�(u>��SAL^v1ҴmFRXn���ʬ-M*���.{8�Ok�����WM}&o=Һ�
,*�l��*2D�t���B%f�}����蝡f�#{X�3�N�f��Vٮ9
{�R����x�����cT��geMhv����Ys4a��M�up3�@���nȕ�>s�i��r
���{��{1U]��T�wP�w+�c(]]t��]Ziy۬K���äe��a�zN@(�}�N]�M�gn��'�ݾ\�7�_hM���I����W��'�4��{vy8=�c	|ļx/��n��Nc��.I�
U*+�P�z+�U��^�_]�4\��g:ӽz�
&���/4Kd��oK�n�;fZ�1cV.��� �aps<mv�O��!G���.tړ��������6s�j�T$�n��'4NC�ܮ<��H�˵�Z"�gʂ��IԕĚ����-��P��,՝C姨�2tiY��.`�5��Э>nb�� ��E����3ye2��r�i��`K[I���MaRL����ɓ���P�Wg���Bp�7� �U8=�wg��%�G!o�5�è�����7������VX�`<��B�
�
�.�U[z��8
|幍�f֋y����j\P�]�ƌ���;���D�I��x/Uq̌���m��l�Ja�:nd:m+ef��4�g|���h��kmiJ�7,�X�ucK�6�Gj��°]��%6�켊6
�0��x��^�w.�T����
��@Ys���b�\�b#D���Q��:,$����豏 :��M�q=�iu�P��L�p����tC%�����{�N=��q�՛Equ�M����[�3J�/(<[m�i�o^�8e9���Μ	���}e+=�ӵZE�v,��z���]�&�o����l��P.
�)&_S�� ��p �4{zE����X���U�I[N���d�u�%3Fj�8��S$gI{%���ɏ*�1��Ap�X�Dˮ�;s^ڢ�j:���Z�[���;|H��ۮ�Fz���.6eLgr��-��m�����oMq�N,�S(
�▞2���U�YÖ*�s*�s���	3'z����e�2�]p
v�b�w�3yD��+ui�E&���_�	���2<�wΊ�ک:�Fb$֓v��#�D��g<}nlUu.��灝qf^�%f�{6��AdjQ��.�����˭��V���BGUn2�V��N(�����'$݊G�l��4�y\�ʎk/��o~�	�j7��*.|tg#z�wS�nب�P�%��>ܤi��3J5b��Ƴ��A���9G�.Z��Y�:WP�3�wF^_;�T˕��S[S����_f�U1��hy.�x;������E���ns]}gI�T�l�t��!Ļ�%̙�-"�� [��M:k���/��+��r�5ʲ*�^+'�έ�b�=]C]�M1�7N���$c�t.e6�͍�5�������%]�#nG�,w>��F�.�f�B5�w�ѱ`Z��'|4+�F�B�!�2M��({U����[���=��' :���������L\q��9��QX�i�ڂ �:�7NΫZi�����iLm+9ˇ�R�����gwF
[��^�Tͺ�sz5ff1�h�j�,�|�b�IqwO)X,�����ŕ�e�`}lD��F�Z��R�$2e��cӶ&L��N�p
��{a줏	+n���j����>�Θ�?,�Vj�Ԯi�)��.u[G*�-N�ѵf�'����VA��r�4���HX���:^�PE٬]t�.��}��m���<�]
�W*��)Ė.4A}W���rM� iu�++���c��R��ċ\�P�wOp�oU.�fv�_������{�{c)5w1I��D�I���w��k7����{J�C2��z�q��--7Jΰ%_97#Yw;���������j��͚xn3Z��Z��oK<���-(�S,�����3��ֽ$�C&Y�����p��^M���"uv:;�4���R�zc��z�����m&�Y�Sq�լ��5a�g�9����}���|;t)�$A� ��i��vmlq�b�N��	��d�y:Y�GLb	j�{�l����x��;�%@&�>O>�z�ڙv��Sl��FpGV�ڋ���`���&�ڮ�Ţ��e��9��{om��1���c_;��M G(��E�Y�����6�'�LV8�ʌ������$Q+��7�t��dj�7Zæ�ˤ�iЈo��W:g͗�]fs�Ř_�jMf<�뛍�-Q��q��]-�},�*Ӻ�D�N�bV��cL̧\\��L�(��QW�+M��u8�ӬPL��7��p6��$q70/�C{�K೶����M�M��{��T����-�\��V�r5�NiݗR�6L��N(k?���xV7�~K0\>E�Qs�mP{��7L�����7]�� �`%�V��5㨩t��/��/k�R�7ۚ���}�45�ns�u�Э��ɫڼ*l^u[��,��5�m��W}9��)��CR�{�D�I�d�u)b.���>u��|��i�8<I*��#��ʊ�ȶ��J�W�9'-�Ux�ĳT�Eș�9EE9**�dDDEʪ���9dDAAxۑ(�BQ�Q\���\̹�#�E�Tr
��9ȣ�YUDr��*"(9�ˁP�\�U���DPQʃĄTr*9AEQܴ.��2�K*���yKP�L��U]:�UQA��2H9U9)I(�B��� �-H��r���Dr"� ���(�DU�9BBʵ.�EV�*(��J����q9�ZE�&DW.r�
IATQD����I�Q�.Er(�+#���V��D�2�"�UDr#�eU�p�.����J�d�~�
&� A
}�W�&Kٴ��W=[�\��9C]:��[f���D��j����}�)��K�Ƴ��fm���l"��=��ˏK���2]��U}�&��g��p�5�ӗ+En�u�wkA�'8O���,�0�{�yg��/ig/@ÊM_�Y�N�� ��E�:����v�q�Pm\PV�\6AG�]����;z��y���[<+'��H&�bW(ׅhF/�_sQ�\���FN�q%�-�k�We�vEt�c6����zG&'c{˝����h".���H�!C���@��)er��S�ݻG�D��r��qz�ꕁjg�SQ�>/(��rTʻ'x��u�Jc���g�+��}ݎ��i����ϋ��B� ������z�gS�����}��c5m�x��vyf=[SE��R�>���ƽ��!,�uT80�Lb<��yNn��,u�q;w�ؔ	���^a�42TXI������k�]a��B�n�~y��ļgE��y�;Ly0��������N7WB�A�B��N�ʈ�u�������gI�|��<�16��|�5��c��b�[ボ�/�>Q�-�����^�ƾ� h��:���[��9�y*ӆ�9*u��9�=qK�B`�[�sy�ghw6�����TR+�u�8�8�[
��2��\��(��� T���
{�qZ��.�iH�f:pv�3��	8�0p�}ئ��#(vu�<�x�G�R�Z�_S��d�[�\�ƹ���x��!��|���9M׌6z.7��H�1�VK�e ꂀ�E�G�Do7�3�b�Y�[�{�.vLQ=�s �.��:3�ڿ\;�q���lcv�i�s6$�l�rXY�<�xB.��Q:H�KU�l
#a��q���29>��n�"�H��k�!w���x'^H/w�� S��M�x�����1>����W���杖�Ԥ���Wq�)���{ �T����PǠ��o�z�%�w�:��ö���[�����3�*���Y�׀�w���&)�M	���鋚�t�WF�
t< �����R^�:���ǎS��V��9Mw� ��D`}>r^"q��(/L�"#��6�'�0���y����M`�e�Zr)ۭ$^l�w�n_*}�:�5�?�r�"P��]�]ץ?��ԣg���mq$ְg�"a~�M J����j"+ێ���;�*|�`jj9�]{ԝ<"�&d�S���V3��HГ�-'2[e�}���(�â�x���� *��M~u��������{w�D����ÙY�2�X�(��*r�7YV��%�DVX̠%-P|y`�%&:���j��͸p��d)�K|�,�t�<V���#�f[㈾b�2ew5���c��&u$�{�*�]�ݒ�ٜDN�2-=�_e48@/S�ti��Ŧ.JϚ;��;�OǝʽX�6|N��u�V:�����U�#
��� 7'՝�,�.�[ykn�4Mx��u����a�
(gNIر{$� �~��p��թ����1�q��}�y%C��:������6ܶV;w�DV����<j�H8 @عO{�}S}|w�^z���G�W�z���S	��ޞcTZ�#����<Uc>�B�Q;��Zv��+sw��w���WB��>=!��t%�%�*\dX��5�aC���Ø�Qw.�o�Q�/ݥ�>��(�xk��)V�`�eb��E��%J�W쇼�T��h�7�x�1��f��R"2�UJd��q��D� CJ�\Y��.��o�̢��G�V@��H�9�e�zr3�/+ �n�"ĺ����ִ{T�hC�tQ��^���pq��IO^�cO6��tm9��6�y
�"��&+��4��t5��C���!���5�9vX5�|=�=��~�ta��2F���6�5�*+eْk�'��[ɔI��!�﮳E8k����{�����e��e�vޣቅwVC�-{�]1&�9��U�m(;g�3�S4��'3R�V�f�Β.f�8� �% \���S�]\`WD���ԃN�8c3�ۼ�ʧ�h���gk�5n�.���^xeui}Fƽ��9R�l���Wt/�L�(	9�# ��0]囇��z���j��T-V�0�וٰ:�@}�޷�ʹqc�S�k]C4�f�U�Hk:L�z��*CV��H{�hVB&��n6�u�щ# \`�͍��px�5ܪ�[���,fҀ��]D姞�k�]l�|b��0\�t�g|ju���9k�ij;��M�gj��U�P�Ms,��Tj=~M_��ίL�|���p�A/���vb�gAV���n_Vl�;x�Tj� 츅cM;Ө�8�G��7l'z��9M@p;�@��Op�؁g�p����QرS=�6�B+l�5�K�Db\^^�ۯG��i	��U�:ι�Cy얮ov��Z}P����A��>in�>��T����g��2��Bۜ�{j	�ia�����%޴X����d\�k��%W��>!_��G�ݗbY�QZ}E*x{���+�ma|�g^)��!1����>��o�h0�|���<���ә��i���U&<�]Q'Y/�8���t�ٙ�Fiӑ����	�f��J���\h�c8TK�,����u���U�n�+�^�/�՗^2=�P�S����Ճ]}�&H۟j�@�+��r�vWw�)���Z�+88��+�#C1=�s&	I��9cMo��W=�=���=�^�zk��Y�$�[Da�T�}	W�#&���׳��C��_1n�Q���5����t��VOqe��	����x�+�<]sDV���P�_b��>�p{�չ�D]sADVLp���xp�?{7��(�j�8H�J|�B���5�!d7ҕ�[�Z]�rl7X��"�'aɡEqC��;��8��}A%L���ſ`�Ԧٔ,�(�eO,|n��Umx�8�ClϏ�Ӫ]�0�5�i�K�·}����T����[��~��; X�KXX�b��?����ѵ]�Kzbsi\�iӣD���l�o�����-������J�D��0�o���_H�*���9�؉k\�9��J/˥�c�����zE�b���]�띌�Apl֔H� �*1�
DYP8AI��[/���~�t}B%�I�K�G�׬�{�
���nN3*|��X� �c3@�P�[�F��Vm`B���������4>���ю���G�"ԍ�͙����:+6y@��:���.E��
��\+�q켬���6	>O���S�ug;I&Up7L8���c�RN
N��e���
�����1�*��2M���^m�h���;Ț����t��J�Q���ݬ�6Y��G���0�E�tr�A�ٍ�'�{�����3tgzg��(����� ��ƶ�D$:fd�b�nxճ�͸9S�[=Mr^�X���ݟo���eLm��$�<�U����� ���L�w=�:���zu��Z9Q��;�aҧ�V_BD��v�TD�PW�Gڋ��qy���	�}�(�J�Bi%kN�XW�~�kn8YSh�r
4���TF�hb��t�i��\�&��Y���3����ёc��H�y;-x}o�7\+��+�󹲲N�w��,�d�c�H�����ok���ڿX�eƧ;��7`��G޻y�n�q��Q����"0ϙ���"��06��A+�`��rj�g��L�t���Vlh�Q)�e�y�M1z�	�"x�q��%m:6(�;]��5#Cj9���H4�y;�籊gEI��|��y��\��NK�T���G��q���hO�1�yY�
rܩ�뜌�㹹^a�Bb��L�6������U	*�Uq�ͮ�xA�~ލ�L�-\	*��r�v�^��+*�
���Cpb��*�6�^�ì�-V��@~�6��+lP��"�כ�������oo;�]am��Y�Wcv�'L��(3���2v�L_��n��=��y��v�6-Mf�V�-�7n:`<�W;7'1��f1)E�k���Vm���S#��޼��$�����J;`7{f��p������.���Fx4e�ڗ����|��@����0xM����j{��\�+T�0�m���]��Q`i�wl��C�%FA��7���lr��F�wP~�/k�Z 5�[%k�O<�ﺮF�����B����:QU�E.�;aT�����Z��8V�ƷRǼ)zy'�t�
�_�}��m���y]�$�Y=>K���������5^��ze��!du#3-4y�	�#8Q4�e��NtVd��Ҹ?�U��T�I�N�0�:�����Sx�s;o9o;����l��X��XU(6
�G��[<���ڑ|Tt�Y �
����[Vb��ٮC��bg)ō��JU�1;�ۏX�(� ��v�VaU���k�����2>�x)�4�~+@T�!�GʻL�/.��1ޕ.2,s�h��1�U��ca�R�*T�.q\(8^m�Y(��B �I�O2��tV'�&�; ��C2����[��s�]#{+	W�˧%E���u�T�/J��S�I��F곊��M�W A"I#ݻ�M��y����3[�2���y���>��ޛu`��v|�f��cևe]᭖ڳ��v$'�}�MƤ�
�q�׽Ld5p�I>�E�%4�H,�s���|�G���- 5����0�����SqZV��CWgk�k�^�&p� 6p���`&�b��qL������&�?��C�9(��KVl�[�_�����wJä�om*;�4BD�^���!�Tp��o�J�(��P�Mg7;e(b\������Wl�6;�w�=$W�N̛n@�p�X�6]�'�Un���7:Z\���De�=�2,K�����U��;��E�9�	ˈ��8 ˪P�EB����c w�S�r����Y�L#.���Y�g��Ü�+߆�,���_vm�¬a~�Lb�>��0�F�X�e�xʣ�땯qк����N��{�'��e��<�^	;�{g�v���'-<��^�"��l���Y�M�\{�~C��F�܊9�*�'Ϧ���N�����I�e��Q��j��γ�����rp剕�����xW=16@�{���������-�pRΪ�OT�x`�1�甔���Ŗ�X� ����
����jʳCN�����/�V�U� cd���r�̢��ΨzD-w�I��S�ۏq���wz5�s�n��`�z���eu>�&�]*Sa��^en��P�j=p��fl����M"W
h��%��*�t�R"�͂�|�g:�����\+,?P+�Ē�fӨEdl�5�]�"� �����g��C�';8bY�qK�b�1�Zg����q���'t�l�Ws��s���Viz��g+�XM���r�� /� �^3%X�O�X�,��ᱹ3�<¨ρ��*e#�;.ĳ~����0I�
m�%��<ox��7v����u�Ϫ����7��O:� �N���T�n�����ڕg�c��;��KܳXv}T����2�ߊ���s6��f2�բ�$�[Da�I�!�Q��Ĝ�V�6b��8�@�Ӑ�ƀ����)�d`�{)d\M�9~�v�Ņ2QtZ���]r`_��k0�ӫ�x���Gr��d8��.���˩j�8"�d_�����Q1]|��JjU~�<���*K��\Oa$�93��Υƥs.T��J�/�74V�h��<�Mίn7;�A�߾���UZ|N?�C��yB���ӂ�q�B�]�-�슘`;�3�:��7}�;R�����x�>ڡɋg�uZ�N�~�"�o�0̉qh�Y�J���D�mM�,�Ht�`��w{�d��@o�s!�{ҝ�Y��Cr��S�L�OY*�B��z�	㽼�Lr�΋))R�ڸ��S0�ȖU�EI���+&�㓤��C�쬹NR�.����&�1��EXiv����g&P�9�&P�W�]!���D:7E@��:L�!�����G>��+`a�?.$���t���Oޔ��vڿ_��zE�b���PY��uƠ0������aOf�W��k�kED�r��9G�"t�s�TGư8�:�`"o�o�U�v%z�̷��צ�H ����-h�uv�6�G��N���`xJ8Szh"}����]y�Gqa×�`�'�9�]KsP����;�</-,,x��������-/'0;�V߮��=�˻�u���L�4>>�$%��|+|��=ۑ!l�&�|���+������F���8���l�[Ư�L%��:V�8Yc�Ȱ�S���4u�6M*〓��T=���pe���������C#�ϪA�P���+|y�e���F?[�
/�Ͳ��r
4�����j��!�����f0=C�}���l�7^0���Z�#��Y.=�ꂀ�c�x]�^mǥ�ե��5F@��HV����Z4��耯%F�;�ǀ�-����n8�1����E��4���oXm �h���#!-���<={X郅aԣ��u��.�Q=�WtJQ���v�)3i�@����}�gz�:�5/��`fq��&��w�P�'" z�.�����P�e�0�e�b�v�U�m�mq�E0m&^����Bk�	͎�XP��鈁�Wgd;iL�0�.���P[Nq:E��<��a�9�$}�th�&e��������
k�vY���w��hՋB���A
=g�I�D5œ!���+�ïS��;�[�ZX9��59М#�%s���8,�[�je_E����!>�:^R3 �!��N�ٗ�� ֔q� ���|�w�^<���ot���rKD�*�}Ƀy�2�=�b��A�!��t#�H����[zi	7Jw4�z��Wװu���Й�gR�-�"7D�I*7�<��V�������ll���x8{���R���9ܡe�hh�o6�8o�� �@m}ҟٝ�
�jD��ζo�C�N�^Q�i'n�j6�meje��F�%��_-G
��tD�W�)�t�8X�~-�����,v�:�H��Е��I	y\�>'x�&�S�j�
"��r�mJ�
Ϻ#�Q�K�o%��4w jQ/�<��Z�;�u�`�`�Bӭzt�l���~��p�9�e��(i�6�լF�+V;�*�U�WY8,�k�$�������&�i�:�e��M5'Z6���Nrp�;���8� �yJ�3��eX���K�#Ek�S(ԭށ��ol�1S� �\툖̬[�V �8Ɍ�ef^�/V�k�������[��n�T]���=�,���H\6�Gs^d��#uN�Fݔ-�P�id$�<�+]d�:�K#�<r���p
���做�&�=�Q�)r���m�=i
�)��� f�3�yQ���jَ���:��[���������W�p���$��������ͫ��K��]�
�H�U|/2��k�b��B%�PN��m�I��LP���u���lf=��잣X�V�dކ)Vu����s�n���Cm�u���>��Y��%���xY[]a���i�o�YX��7eE��%�p|��4p��"��mc*��~��ǚv�i�L�>�M�ݽ�^��傸d#�7t��GA�MV=�q+���N��V�(̴4�9�6����ܲ�@o��X���s]�U�Ni��BnwuaI�����zҭb阨d��ĥ�\��\�wY������I�K��,�=��"�Ԏg:�ˌ=� �/V�ι�{�,�d*3#&>��A��ub��]��j���I�i��}̩�=��5�-�~�.���6�n�D�s���顖��Vza]3��Zμ��#V����|��L�V�g%Ӽ�k1�n�g0ҽ�i�zۮ�͚�U�Y�{��wF�3l�a�9��e���nY�+��4����h�o���:��T�Y�U�t8/��x�C���B��T�iPR�$�jZ�4,P�DW9W&D'J��J��p��&J���J��C3�EAêF �'B
���rU9t���(�"�0�D��.DDPr�R���Vi�j�A�$E5�DTE�gI�L�4X�IQ�TFvE�s��(�*Q
+�QE��F%RBW��(-L�*���/+#�yH�$�h� ���9Lpl��]YgT$�"E�EΣ#*�
4�r���r�����Q�+������!jVg�&Tr�V���fF�Pr�0����r�E�!V̑ZԊ*&p�X�*+�hf�L�T*�A�vTp�Y�!em"��˜����2�H�)Vp�QT�6Q
��CG<(*MV*�*����q�8�V�g,��@���@&�s;�+������x�H!x+j�e���
��Ҝ�wM�.�n#1�TR��/w"�`�$����r�N6��!b���=-���|L.㏩��n�c��8�U;lq$�&����N���tt�;q8�^�Q��n�F�!��T�v��n# \d8���TG�=� �`ZW��#�=� G��}�'.,�ח]��V����t�������I�!?��Nw����v��j�ïxS�awI�F���+�M��8����F'y���i�nӉ�n��O�8��v���|� �G�V
�<���w/ϻx�?}�����~A���'N�v��y�v���-�o���7�N���~k�&����<���#��g�t�x���p�6㴛��8��G�+�q�'�\�<l�7�]�����Ou���٭�g�#� 8�� �.�Q� (����y���aW��΃��!8<�s�ޡ��۷Ǟ�oS��?>�u��nА���t�-��M�u��0�q�� �}""���w�(c����+ܛ]~���ﾜt���_N�׶����\7󾽦��|��m;���w���[�|L.���<��㏏�q0���6QC��;���mז˧t�'����۴�c������1��]�nl�W#:�{���ށ*N�pzQ�&c�t��� x��#�׎��'�p<C��ۉ�C���c��!>�|��}����κ���>&y��6������(� �p�o�o�U�YG��{��q����b}?��}q�t��q����S�8��|9��0��q�\~�����q2����C�s�w�k�����v��'N����ہM�ys���a������p|��T�{�}�d���%I�à\(ب����&=Q��==��?�v���������k�o���ޡ�q�?��aw�|w=w�t�Uߺ��t��n���#z���H�����|E��l9V�E��lL `���G�P&�>��s)�����u��޷�ݠ~HO�����v��ӏ���[t�+�gq�޻�~B�|��ӼM��9;�;L.��>�q�p�	�V�^�2/�lX�׿w}��vQC�~C��?����eӽ~����N;w��n���n{󿷿y�0�z�~��޸���;�p>+�v������ۧ��v��p��t�ۉ�A�x��} ���Xn%䅝��mS7����k��I��N�f+���η#�..�k�{�ihG羯�،o��$�M}c�3���<�%P90Ʌ!�4��)[��=�)�훃H���Y�<��;�`�Fƾ�ۈ�KBN�
��Ll̛�:2��Qe[�I�ggި�x�����l8�#�'��Ѻx�ݟ|��&߻�o:���Þrt�8�~M�8���`�ާ�8�'�~p����|�e���pvxeDL�����Ѻ,�d}C᷿���}7���8>�)�|@>��1�(����O�P=P�{�H����/:����7�ݻ�����S���
=�8�e�t�m�Z�u���I�����
z�!!ױ���q8��g-��8�u�p��v�n!'a��7O�ߓ�?wv�I���o�<�����I|�yζ�Ӿ�N�~����~��G��~�S8�z]y1�4��9�É�<M�{�����M���v�S���_����P�n�?��ܺL>[.��^>&��v�q���w�m��o���sv�]���}���� xE�ӝYj��9�3�Ѹ�s�z�#��8���t����;�O}��o�O�n'>o��c���/lt��1;�}�����t��~�:v��<r�X�y�����o�w����o�r����<��6�D��b>�>�>��?tC����t���8����}�L������z�v��#���o����'�׼�#n'~GIӷy���v��q7��|9p�v�~����]�^�c*����=�$D�������0��ӡ��
�(���Ҩ	�����w�y���޻�8����7�$ޡ'�{�:��8�}O��1�ԜI㸝>;q7����������|�]��{]�y�����"�}���;���]�Go;�i�X����qݟ���I�w���߽�;�bw����N:wI����~q�v�Hqw����D Dh�?P��Y��"u��v�O��3I����c�
�*=�0>Hc{�nyc���I���w�s�o�q0�u�G�n��]�|�ǉ�z���O�z��!?�߿wô�'�=�ݧ}�y>�'�qP*�^�>��Z蚊���s6��\��=�H�D�����������;\��n;��'�ھ�I�ߓ󏘺����L)��z��돨q����c� �/������> z����F�{#ި� 1��}�I��{���g���O�U�j���V�,�G�wP���wG�dt��A�`6ȹ+'da��s��I��t8�����OOr�q%r���!F�J$Г*�]�/k�O��{��9�at��t��	���Z��e��|�y��t�S{���A�N�<�����v���?�O���Nv�!�����8��`�o��>��+�#�C�q>r?��N��~wo��޻�8>��_0Ղ���Q0ԃ��t=����Ȯ��VE1��(`|7��{� ���.��O_�n&�~�:C���m�9������������&�����t�;���z��o����`�o�0�#���q鿆�M���1 ν)����~��鹨�ǃ�1���8�y��:We:��ޏ�|L>�}<﮷n������N=����-��>{����S�|����� |��>;q]�����=N���^;�������u���CBIk��� cc� L	��7�q��ۤ����s�;w[~'H}���w�����L*����:M��w��#���ۼOq?;��|ߓ����?��� �����YΘXo7l��g.ߦ<�x�ǅ@�����/��w�c��;���V�v�oP���N�{N��[�:I�ǞF�p:wn�z�����|p�];Og�9�=N�z�W|���ާ��?;�J{�����Վ)wI��X	�;#r�5������G��{�\����q0�{��]ۺw�q���+�	7�����oP�\���۴w��t���v㏗|�!�i|��8v��$�����m�|w���t�7ޮ<���e� E@���;������o�����7��x��w�|C�щ�?uc�ӎ;��~[����|w{�I�]�S���8�|��q�t�q����|;L.��n{�`��@)5A�T���:�����*�������7�8���:��n+��|���$��o��c�I���w���v�7�۷����N������'}@q�;TQ�Ӕ©���4:�T�eGnײT_y�}��H���λ�����q��;�ލ�|L.�>u׽bO�~C���w���s���c�	2�'g�}�o�I�]�w����ۉ�O��Ӻv�N��aC�;	�[����y�#,o��{1G�|G�C�G�׷��n뉿��8��D"@�@P& Z�Z#�ǔ���b��q0�s|C��;�x���xJ����=�v�y�|;������(ԯW���w����z���f��b��P�N�k�A���U��<�c	���]��S�Dը%H�?�:Gc��5}:���N.��;�iMGF�U���}�VԬwӢ�6�e>)
��9Ϩ��9�sw�V�I�H&��A�r�o)rxgҫH�vm��)�����c���n;��C�8�_,vQ��&�A�s��o�ӻv���x�޺w���p�&��o���[��S;�������/#}��7��w�����}D��Bg��P��/���^��������vQ����v���0�o���t��I��C�[��0��,|(��o�q0����ױ�C��ny����ݟp;@�$�����u��;I�B~^�}���� D^S����U�`��l�Ny�w�������-�/�n��ڭ�>�R�]۵G� ���aT:?X�o9��둉�'�������wל?8�?��C�>�������I��X��#D|�<����:�\���/���o<Iޟ������n�M���A�N״����7�I;<����ӻv��Hz����t����&�8�tp���d�a���u�^K���w7ޓ��o�YڊE�������wz}���g���Y=�J�>Į����ot�=a��r�kN{����|Oޖ�m*�yL��rbu�}T'NE���>�K�naט�yМ�Z�$�`��rT�P����m(��`q�f�9��9�FR6�,����z����ڭ@�i̩��D]�2Lǃ��N�����8	����޿���rF5Wfێ������Y����w�M�<������e���Ϯ$���t۹[�]{��K��ϔ�5� P��-�[�z߅l�z<2�\���C$XI������k�fJ|,s�fK^u9�����ġ���>���\rC�f&84R
4��m\Gz5��-�X��cл���'�k�K��X��� ��&x	���J1@.���c��1ϔ{�f\�t7����n�rݮm))��]�Y��|:ʻ���(�B
5�T]=9��X�a�,:�C]h�|Lp�I�x[��A�;.��xkVE��*gO��Y��5^I[ボ�/�xi�o�(�\�,E�F%`.�V��h��^�� A�tB-�n}}uI�n|x���厗�cOX;����ݱ��R��D:�'��t+�	� {�T��'VϽ����U�G�.��+��Y}�����u�Y��y�:K�O���1���48����,&��]F�Dl<�4�@�G
��i������F�b7���3����2E�.5��lAt�N�Y8�q��b|%m:7Eq]���!Z��ï<�ϮLk�~��u!	T)5�V���T�.8Ł=U�������,���~:\Bs�ǵ{,��T�v��Ҹ�Oo�U1K%2h��#_P�b�ڪt�W Ζ��C�������Zݫ��8�rV`�������޼��u\B}>ri�����ج������Sw؞���h_�vPU����WZ�$^l�q�jo�S��P��*l�"��k+*�@��(�����1��n�Y$���*fd���5�diِr��g<�+{�t)n�ys�z�v��T �M�E��]�����Y��.�?�g������E�V��{2VWR3�42�^��k`�o�kv]�ˣdݭ����n��X��$��$u�߱x�l[tb��K�߽�xNWJj�������^�Z�lOye���S���O�{{q�x��mM�o���hIU���B����5�Ox�ם݌�F�U�W+�#�!���1`:t%�c�O�`1�+��d�����U���֯b~��+%n���s����N��@�1��K,�G�z���=vU{�puz�ꘉ4�߮�y�1z�tJz���F1=u3�GS��7اݐ�����J������m������=����z�}��A�W ��x?��tmT�S�Y"�q:q����Faq댙�'+oN5Uv�BP+&V3�p�x�'_�WCt��v�U�:^���!6o���|$����kM��,�)��o��A�A;vFIf���2�*Y���{��[d֛�*�҂�2�1s�_WXq`���w��Gc���'��H�� �WB�}���{,E4r�i|�O\p���1�ܺo8��}�Ӥ�3p(�������upx)�TP֏jZ�?|�Fߌͻ�oϘ˺��%�[w2��g��z5�e�Y�rw1н��tim��u��h���Q�����f�Z�[�G稰����R{r��B��
wrQ�X닻$bﺶ�ڋ��1��{���D���7R�r�܍-��}o�.���`�)��č�]n��9,��K�B��|���}���7�K�x��u�dY����Z��<6�n���dzW������%�0u��zk#:^��5�:��,���I�B����4�k��/Yr�Wn��	]ޑ�wg���V�y�~��a@b^���]w�Vy���q�U��?�Y�^�͞;�Z(��[�|�E8�hh��]ת��ǋ�yS�w�!�#B�q2ꁃ�e�
�e4]hC$�W8�U��uR=�B��F�ݾ��/I�T�4p����ЮA�����
��u�μ����r1��S6j[%�����β�qQ��j��9�q����״_Ffnbe�=Qm��廧Ny,�_y������ʈW���7�QPUJGP5�n�h����]�~�F��&�c+��T+En������ixV.C�h�ǻ=�ߢ1.=#*��2�`�Ʊ�!_�G��$&��q�hw�+_	�I�ݞ���^�zo�B�3>5n�hU���;, n*����uhÂ���B��e�-ެ�s0�;* �| ��^ߗ��ǟ��
��@�*.����N���n��U��Q[���i��A�����4��h7��F�Lar��n-��Β���+�C)aB�O�}T~�z��9�.����D-���M���X"䢣�+L�>#�+���Y΅��̜^έ^Ze+>g�7.�3�x�!i�}F6ӻ�6Ju���<	�X��Y�i�S׆�¦�����I�K�����1h[p���q\H"��+��L���O]�ׇw�`�2�@��������ݳ�*�C�p���qn�v��uTF�{o,��%���8_�"����j��Re���V
��˭mQgjZ�*\�VT'�m�=�IM@�&�σ����+��;U�>lӤpy�i��_q��!�8i`nھ^)mϳtgL�O�f�%�\F��\D���N��0��yB�un��d����A�n7PܚJ�H����}��]��8���iy
j2�]�D��OW��i��p�W,/g�qM����[Eq�)��)��V9;�9�΢���m��q|^���t5=�C�-N��}���9�7./].'��L��j���Ɋ�SUAg|�^Hz�ok����i����M��������4.P��n�L㾇|��YdO:�F�X������$u��ͮcU����3('�H��{��O�Y���R������-�ƚ�Or��Gr��d!7��`��<d��9����3�ֹ��Oa�{ȟ��2��޺O�����<<H���2r�����i�77 �{��/�����_�
�՝��|w4�OJ �N��m?S�<je�Xg�\½���Y�/��c�U7���r��_����w3_�����6�#�׷M��ѽ�<{�Y)Y�@�����py$�$���z��&�-�7Рdb&)��<��:��z?���*��N_#�.���~tUw�6��N��<�6B��������r��_��l�t�����аA�bc�N!Ҳ}���r���ы4�-�����ڐxЎ�Q)*zxs�e��?p�S�+���O{�w�ZVtoq�%������B�t	�΃wO�S<���Ɓl�dX��:9�i�AP�c�-ɯ���6�c��oEl��GK� f��S�1�H��ճ��o�V�.���~^���&���j�7<�7�(�±f޳��"�0!p:H�<�ߨ���뫞�u��d%-W �Ọ�+/��/u[��D���A7[r����h����D%����U=�Z�8%n�KAZ`ӧe�!÷[A;;��Q����ݖ;;tK���k�Ѻk.Qf���`�7&�7̅�)G�F�:�n�Eq�N�	;q��vn-GA!͗w�X��k��cIo	 ��F+��*	+v=��%�z�d��d_J��2J��C�}�,W�6����u[�폣�����Jt�R `��L�7Z�%�w���Ӄ!0:�RV�7ï�{��b��9G{��߬6�b�JdѴ�Ds�uQ��,�9�����P�p9��K�I�`�p(F�¯T�P�������儓���),<�"u��=&�u�K�V�5\�wqz{L�DGH����FB���gZ�$X͕��7,r��B�j��(��$�1l�m� �^3~����2{N+y��߽VNT=�匞������l կv�.��7��V����2�����F55��O��f+K'15>4n-��������+<���8�P&00����S	Ч��SS�8s��gN����2��*᭚��q|�Eg_8�G7��E0)Uq��@hƖ!D2�c��/����Xs³=θm^�G���E�ɘ����;��Y�IP�*6I}#��D�C��
��TB=�������t�N���p��ۿW�yg���υ-� �:�\&z�/�wN��$TMN�{Xr�z���B�7.:��W��>0�}��������CV<?l����`�9���4�L�tO]:ʡ2���Tuڰ�7��4U�_7���O�w"�]�w�PۻX��Ԭ;=�u�VU�+7�~�7�s���c*�+�
-e���iq9��%�ɫ4��\w���6��TE$+p��5i��7Z+�[�Y��b�o�r��<�l:-�=dJ�9Ɏ�&uv��������vβ4˴wN�QP 3m�_P��(�p�c��4�Pܽ���F�Nt�"���ۼ���j�D6؉�.�[N�Wa;���{���Ѻ�Ag���5���?Z]�:��k��Y��>%��1�	[f����'�	�w:���c�A��s�����Mh��t���n!���^ԏ/p	�v�(�wv���2/o����׫�JyK4�����Q�b���I�K���v��4I��y����Y����V�����[���B�7�i��­�AY�;+�ږҁi[�h�뇞Z�4�ݔα�b�]L�fScR�T�����]i+U4v��zT�VnZ��Ъ�١w����Ln|YR�:�W�*��V�lHVVe$Kd-�J�o��s6�Y�C���3J�ֱ��t�,�}���7:��+�؎;�/�����=��]C�ٻe �O�f�@$�l�*޵��8Ts�]4�#W�L�k
״�^|��|Q�G�k�����p_�o��M<�J�q2m�̱�T����*0op��&�!��µ%C���2<�����^�t�y��vЊL)�3��Jq���:ւ��K��!ۻ��|g4�I^Y'��j�a����UyB��Q�sa��p
gP�Seǫ�;i>�{������)�Wz���a��_#�����.o:���o2Ʋ�vK���͜��"a�G\�Z�*�+�*��>61�N�]+�6��ͬ�������Zt�d,��KN*�@rn��*:)*�`�b��l�[B捵�m�%w��ү��P�}.NH%��ԙ��q馰}-��gTc}�QM�l6�ԧ��9H�y�u�K��af:ܰ��6zJ�B���Z��o9Ĩ䔔�V�q�/���;Jc_�t_)h���eSCb�j�_]�ԛ�����zd��ĻA$�x����4��d��b\g:}��O_t���璻&=;x�
��4�Y� �t���:c6�G����a�׼X 1ZSG��FSò*;y���j�qY���¶1�
:�V��KH�Ώ�.��X�r�9�������傸im钗v9Ĉ/G�8���gr��a�uv���,I^ov�2gm�
�F.T��^�r���&��K4iu��B1b��;��+/)�l�G�����8p�
ؕՌԧ,�x�La��#�]rμ�ZIEn$F���sf"�u�p�Bѕ��*����"�b����g/Lb�[�ze�U�h^�f.��Wx^H����ФH��l�e�$����\�PUyNDE\�R�UU:x��"ҌɔyB��G9Ú`ys�8*�ҭZe&���#7G��dQVG,�Ԥ�T�(�J�3��l��8�$"�ũ�31
S.�t�aAp�rąY)��g�-Cq���������I���P��i,$$�9	�r�ԮVFU&A�"3�EG$��%q�ĆHar)0�I)��((��T�p��*��\Np�ʹq�$�EA��K�eH��<���QIәf��㧉�Lr�s�iE]d$���V(�����RʋnrIg�"LT��ҳP����NF�K�u4�9�jY5K$̒dZir
5S)KZ*)\Ua���L�Ҡ(���+Y ��t%Yjԫ,�Ua$�Du3+KT��N�*�,�5$�	�f�t�"�r��"��ZE�Y,�B��}��O5��jl�%)'S0�\k�DYw��.��J���/r�{�Q�@=l]O�ݜ��4�e�Ţn��YgtO���
����KB"4���av���.+�$��\�t�<k����z>�Ю���|\�/$(����^O���_�;)�5��������a�%��xoI���xL����w��:�j�;�O	Jt����]�����VS��룉�~T��x'\��Ʈ�U�1p ʛP�t�޹�z�,������0�ƽ\�$p����yY�����%��(�T@ٍ)�г{�u{e%��t�DA���(Izr3�Lߴ�#yu:<����˛d��"#m���O���tG-��c(��d.7��c�8�#��;��÷=$PI;2V>"�9R�kqx�߱;��e�s�O��D�>'_���C�ԥ���\�eϭWn��x�w����fon�ԵF �1/W��.�ʫ<�}k���vPY�漮��<!o�;��㐵�9`ue��,V�Y����ʋ��k�f����;6�Q@u�H���}�#�2���.@Vm��u�=�Ea`ԅ"��y�ݾ���X�q��J��sCD<>��V6�����'��B�F_V�`��o�\���!���lT��"���.�RT�i������m�G���],g6��t��܃X��aᵚ�2�1ᠵ����u���^���`��n<�wJ5z�5T�p\%r�0��_u!y�Ed�*P���Ћ���<
�Q�Z[SFQ�YU�$�%d	�}a�
���H��w�W�5Y�6j�`Ф�d7�{�ʽ4Ǫj6l��%���͉�|ǵ<vT��Yǁ��>㣅��^��*s���@����/NA�^��A��|
��4�)��8��L{���M�u�7[�5���R&���:��C�HM4���!�+��U��in��p�_3�b�V��x'�@��w���$8�s���=6]t!D��I) dy�
*��UF`�I������K�;߼��O���W�T��0��s�o�~�I��	�� jT���3a���ϰ���!��}��z��&�M�L��0�q�y9�^���]:�d�0�w$�F��,�չ���ڙ$5^�S=�8�ƱutvJv��R8��0��:e�v���(-�]U�;�x�<��u�[XH�#����^A��Y|��c�.zy�����ހ9���\�Y��	����9t+��:�"d.�m�#�ȡ�iM\=*�[����G���mv�R�ZhZ��ۆVY�ȞV����i�t�Գum�F��	W9����y� �e�������{|��y��<�c��A˕8�=25+
��V�s�0at%�+��3L�U�)'v���G	�S���;(T�⧋1sB���< ;w�ָ�k�3�mO�&���C��=�N@�ǉ�
dz*���
��L[�]�1����a
��s�qͪ�7��bRr�4���!��`�K'�A�Ҁ/5�s$>Xf��6s��٨��q�����+]VoH79��4U�$.���u�099Y}��cr��Pʛ��g~}U��e�ǘ��{=����^YA�+�Z�؞��x� �����IA���H�6kȲFQ
Dd�+�� ,�4�K��׬��
�(^��U�b3\'�<�`g�Nٯ@�PD�uw�k6�_
�����/�X�3 �P�&[�J�K��Pw �[�=�T��w^�6�WE���`Yd��N�P��X�����>�=f� ��Q�}�ꁵCDX1@b�n{C�p9��8Ε����6�ΒtГ̊��(�T�ƻN���}���$o��v����6C��g�w^Ϲ�L��g_$u:�FW�>��I�|� �g:�M/�cTt��X^�/�~��ˍj�>����ߗv������4�Zߢ]x��i����<�^h���in�?d�N��\���(&ܗ��Vҫi�"l�@��q)�T�4-ͨ����6.�Au��^�ZPe�&�뷳N�uo)Й.�'�An>Y��������sz������ov�z��q�J����bJ}`u�&s��x�g��y�C���͸���{�i�t}UG�'�Dl3j���$W�����*N�:9jmK�;�ώn��fr����~n���n��b�3��0!uD� 󞣞�6O4�����t �&%)���6)��F�"EË�My7[r�����>\h�!�N�4H66�V�ssڋۃ*���`.�8��5q�P��%Z
�T�/�1`t�t�MߘY�p$s\��'�+#=�{~��Ȭ<�ѱ�+����a�BaaL�<u�:���vVO>>U�7öKi'�j�y3k1�mm��.����n���光;�F��&�������~Fң��W��F�3�4�yWm���X�^���	����q�<)�Y/��gV'T)�{Ҳ���1���|m��J۶�ʬ:N`?u	r5�;�<,���ka95�	�o�s �͠��2���ʟ9��w�>�e�L]���ݰd,4U��ګ�*x�ӵl:�'�ui�@�6�M��n��-y�g���}:>����Wt/�lcAM�N����N駍�e��?n�ڼۓs�E�ݑ�I�us8���el�� ��]�2��vͨ,�MjY;j�$?�q2�x����d��nnZ��73��־�����+l�v���� fo�X"C���c�1}N�d�s�}6碷�h�Ո�'D��Gڵz�n����BIn�,T:ze��6��ĲɮS̾w^q�����������d�}�z��ȓ@`���M/t�j�H�SR�
!���ek������WN�䄠z���E�3�
4�q�� |+�:�^H��t4�������,wf��e��%I`���v�j����}qP(�O`2�$A�$:>U�el����[��n�X&6�&���h��1�l��8k�۰�ђY�G���D��I[]�2� ����˔ū�Gm�tc}Byӱ�~=�Zs#�h�|�xUĞ�i q��=ի<��w��EY~J��=��}x�C�LƱq�W'I�@l�yY�w�/�Ub��ٵ����=ݒ���xT��,DA��@�%i���)��č�]n��#�8��d���_3N�]�mu�:�9b�9�M2b��A�Fd7b:�+Ҥ8��;��+M����g�d�Ǖ�f�޵k���#�.���Wv��-m��X��3V��'�ua��;́�����ZY�d�Hv�-�N�Q<u����0�o.Rm��#�8�f�M�2���,��{E�����#�ܠ^���,;Z�u���| ���#��(£y���/��w.�J{�M��Xd�1}
��.̓Љ���.�+�5�|s�ږ��o��J���{0֣�1u�E���y9qhs�$k��5����d��wO���0��6[�P�]r�����j��.��W.,r�p-o��~4�+Y�ySdhS���;��I^rn���y�Ȼ��Vz�>񅪱V;Ke��q�a�49S��Ʈ��۝�TD��-�|��/�y��k�p׉�h��;�ZbO"Q� u����e��(g��u��]b�1��Vv�%	�j���!��r6nR^�_i>Fŗ�N���M#zu2�&�F�<�x[k���>J����唔���p�^����
���WX��=Nɕ������u�N�ߢ�
���l� �`���(.ʔj@��g�Z�Jin�Y���x�OT�{��x�*~�۸a��^�$8��Ql'~zT��!D���J�>K�N�R���Y]���Y��;�.ĳ~����T��9�_��o�h���]��'�d 4��l|�T���p��t�%1�JD�\+	��Ӯ�U5Y�Z���������R�ywP�;�Ka'�	�1�4w�gk�:�m.���a
� Gu�ω��v���R<�N�\Fs�p��!<�!���A�6��SXp���VyqM-1S?'�&6G�;�U\.8)5bne�q�!�i����n�aڙ��Jv�k��]|Z���Y2��aU��#�� �:)�G��|흞�}|�Ldr��@�C�����`�M�F�=��	�$x���+X�BG}��O�x\Ҽ:|{Oٞx��#@z2=���Egۥ����a �h�p��|�;h˓�"d%b'���py�=���|c��W�g�=<�dwl��Q��#���?R�J�(^눐�#�'DXa܊
e�A�Xs�5�'3�Z܉�C�����ܽhy.��cȀ�G)@a^4<��N��qSw0��,Wf�}���.n��RI�ͥh�]D�x~��w��g�]!^��w����u��G�����V+@g�xZ��/	l}���]�z����C�/�̫'z�A�׊��v�t�i'K=��|]q�88��k��V:�r��&�Eְ8l_	%�+ee�#O��x�W�;�b5�p�́L��9ƀ�eW+�x:��(�`x?VU��Ȑ��3�b��9��D3X*~����[�������,�4�_6� ���b�с��B�ͯOԭq#%����٦�6ywWf�1I}�
���)κ��5�D���U�V��hy+lC�a��X{zE�:�Q��$=,����l�H:'&Gm������{��h�m#��LtG��{-�O=�=��{t�y]���vY)_���#`-��	�V͇g6����8�zu�l¢���5`�P�X��1��s��8�zg	Y~�&{m
�1e��5%�0�j~ww0�;^�#Y�iAF��]��]=;p�c���J�nzV_B��4�X���i�[i�o]�&�g�'Z\�v��iq��Tt��+���"��0��$�63t�_{&����=���M��,s��8
��΃_���FR���8,O���P�'�=�{z���v���i�%ǲ��#��� �ό���c��D�����/�mM���2�,N�~�o���_����q61�M�4ϔG��t�T��Yi�����g()^�.z�t�ᴰ�n�#�7�_AJ������%X �|<kn��F�}A��7�?`�坳��tR;W�~Q^ԍ��&��A^�� 0_�b����O��s�VA�u,�9��:����a_�a�^��7��+��'��mP���S&���Ds�OƸ�*9��Xf�;���5:�R�Lkz�؝L<T�S���^֪���h������Ѓ�꡸��y��V���vo�A��u��8��e�J'dm�o}oթ�4�h���C��b���g/@��P��O�Trl{0�a��_88d��������_W���M�;��"�2�q�*C��'��6���qg&�d�*!|�1[�#��雱{J��Ŕw�����U��[މ
�xr+�V�,fʇz�K&�'�!hy��r��3�}�W^�1Ƨ����,A+nڳ>ä�J+�@ݐ��=+�)q���M^���{aAO�m�Dn99g`��O�����8���hM>&��Z���"���w�;ժ{&o�J���D�!DF�غ�_S��,��&��_��tg�)2����k�����;NY`ʠ�R6:��aP8Q+zu��!��Dfr��3 �n�f��F0TZ7'a��$H%���i{UO�sӾ_k��>��]�[��_��U(��J�?R|�{jiq�G��� 㢸@�WIk�2N�M?C�׽A�1��P�I��Q,k��\y���FC�G95a�x)�d	���N�+�T�!�*�5-5�r��������`�:'X��q0Yqq��SD`�1�l�᠝�Y,�gq���e�
�~�l�\F���|�5��Y���]m>����7Uԉ�^go�m�}�ʳ���|��(X�*X��s��J�e�8��|��M���k��9�|���b����G{-:��m΍�w;.eq�
W���sN����t�{� �O�SO��U�}U�;&_�����v�f��X�X����+)��:��lc��]Jd��O6�o&�Bo8��� q� Gnփ����Dw�.5��$p����yY�w����\�زiv<�{�� 2d����L@��	��RV���4�fƞ$mˇ�'��ׯ<����C<\)t�:�<��v�O��7E*�J�:\���[9]MlX߷/׉Z�Hy��K����!�j�&ې5؅BƗFI������Ђ�����r���z��F�X�5ݷ���=w�ʪ��@)��(	5�T�Ѡ]����݁f��7��k"�/c�oآ�{�7�Q�LKWG{}i��*Wg��r���X�ySdhS���>=v�=/��%5λc"��u�ѿ��2/�S7�}n0A���*p8]D����&����7d^VY���Y�Do��l�'к>V:;o����#VM����O||N3����b�W2&^�:V���简�7�ۇd�ow�%I�񮠶F�0�@�#1fdջ*v�+�o�(h�X|2��c�:hwieq��Em��1m�b#��J�9H�R�8��{�v{�{]����ֻq8��ci�\�w
���s�y@��������΋+>�э�d��ǣ�u�RGk ��;R���Ě;2C`8R��4]�5IW}�d��&��w;�[���-r�ӖX�2�5O�f�U�cRN�s�Q�|Π��vL�X/���F�۰Tb���*ң;�^�ݕ���U)�O���2)�^�I����wW�g�fCx��ҠY�\H��O�\Z��Y��q��vs �H},�^nwFe�u�#�G�Qr��q���/MM[A(������,�(��ޭe�Wz��AO�:v���eY�1���m�&m��v��u�/�)sR7(L��ެ�(�u�l�k��Gl�CM_L�S�Q��(tD��{M漳���KfD�:�:�)
�=�	řV�4�7սO���@�c���9��c�=3em^laܤ�9JAјξd�Ns���l�YM�V*b;aA}q	ج_y����C�>��&��M����hF,�Y��֨�^�i���;55�s�}Z��7m�Co@��J�Ic��yR��ΣÙ&
ÐK�²QLOZ����+����E3M�B�Һ2�¢"�lY�ض��B����enB^�|3��(��R�p��n��Q��n��	Xz�i��&mԴ��Ak��nm�X(�	-����za&`��
�b����̡�S����7DV��j๸.�*�p�j��'v����wr���"�a�W^b�Jm�SnWv�]Z括Ka�/�42�e*�Mb�<�lo`Mq����C���{{J�mq���d���(�v�&�`��W٢�u�0t�oy����6��|��������/Gz2K;�J��!��:qT�vL�9�p}��Pw����SR��h�,�dn��:��`Y.a��\,v�q6UqIH.gk��GN�j�%4'����l�'��:��)�#3����K��у-g<�:$6�ɮ-m;$�,m7"��Ы��X�u��af�Gi�qmu��@����%��Vz�h��u�,���m�+�w؍4r��y�:{��".���9*��j{ KXޒ���7ױ%��]��Z�S4(3�q\��&���� 4�̲ ��#�\�麵ve�ցD:a�A&Od��s]]t̬�(QѮ�XT��՝�6b=�NvH֦�dU7_v���CV��ڏ��;��;��������b���â�4=ȯ��w�k�8��SqշX;+n�2�α�1JoL�к�}�E�)eU�쇧��$W��x_nf��(�Mc's���a�����]�G[�)k�����YkYn��'<2�Vu��/y�|�6�W�L�%��2Ԍj��)�꛵�n�M�5���<�抷���,��-�SOR��Z�v�*A׽���8u\�H�}��#-���a�c�-O���P�p��b!GBhYf�B��P�H��D����I2$���t �$�V������3D���)4�V�êIΜ��ETETb�E��&�J�2�4�dQVf�QF$��N�V5TˊF�J�-3��uB��V�H�Rå��(�˒��REE�3Ihd��9Vde,�U�H�6(�RT�j��'U�!dGJ�ZF	r�Ȣ��QuLR*ԍJ,"��"6�J�0��LْVA��N�B��3dF%D�T��U�&'EsEZfu�E\��#$����C��T�̸Z�h�I��Z(�%���$ՙtP"�K:DDf�9H�L)9T�̖Ua%TZj� �V�b�E$t�4:a��	EӡG39"Y���]*�D����JaFZ�]|����.��cwB3�ȶ�$ݬ�t��^��d�IL���������-kv���l�ºtݲn��ē��}_}��S�u�>�틱��1^�����S�����W�Xx"|*��yi�G�פG�#Z�ȭw�a��u����`��_AvT�vD@�>L�+_	�>w6�Sk����j�׆�P���5S���in�3�ć�brw�«������y$��{.hHL�TN��bFdK��2�ݚ�B��ݑg�&�;�s��u���1��ߘ����r2:+�����L� bh�r��N^y���j���t��p�� m�l�6xe<o/{����b"�e�RR�#��9���^���qያ��Jv��Q���T�V�h�9�_)�{H�b�7]�yѹO�x�9#��DV���7ژ\k�?�o�T"�0u�q��=QIK̥	�>�/v�8�Ֆp�h��7.��#�	Wtl�G�Ͻ�4JtyP;玜l��gr"X���֪a�{3�T�x!ˈ�+�!:GN����\�ի�,[*C��t�:/,8;�ZK���� !Q��zMYV~��UT5x=��9�k��p���$��I�M�Fw͹;�F;},�0m8����uaz���\�'�� �aT�5��ͻ�����;ՏP,��;�|�bw���W���M�;y���I�J�|9�S̬���lv����g����>����~�����s��k��>|h��b��M��/�G�ۓqP9���w��;��7�x�77���IW#���3���Q����q�:�q<szS63�_�)���]�N�ׄ���S���^�	i��wbz�c4ב�{J$e1�!g�NQ��,���J#_Rɬ�R�����P��2����n��Ӝ-� S)��]]�yR�UמKњr�eqx���	wĥ+�7}66"ۮ�:�y���=�w^�6��omO�J]�>��f�,lvé�hԎn��E/�	ҫdѓ!����ּ{�LW���ѭ�}ݵW�I�W|��4�n��$�~�|`������m*�ˋ��=��X�a�,:T�M��ZJE�{(\5��fq6j�eK6I�%�!�u���cTt���a?wOi�s�3'�����;���QB=��/:ㅕ6��>�}�@�$�gA��ҟX�L空�҇�V"��eN6�tv�6j<�v��s��ג��^�p��#���5�P@�a!���qi���<�a�id�I}��&�x/���p�D�ӏ]�v�2������^\����L+�3=��ڙ�hf�;ĕ���wY���۲T�6�Y�J?3��e75NFXV�ہ�2�;�ə��!7;nG��l��4.B�tV�,BR&/r/�D�������1f�q�BZ�����qт[V���N����<(�>�D#<`B�:H�5�]����֦)��Ӫ��n[4���7�W �t�AMrU�J�p�F4�f��4��p�Z]�Z_��9��lQ|v����5#CR���M�Ax!ӈ�����T��c���\6ḿ�p���EIL�Ҹ߂Ooͩ��fv>��l@������#��ܻ�����$�U��\)�������a�_��Y͂*yAq�=be�w��,[]��g2���>Ri��w�z��hT"��AU�uF�fƾXM_���#tﷲgx;������`����y5��_u�,A�%&�J��7f��X�<�4$w��Oy�c���&�) 7=�_G��Z��V�}_z�%V���5�Ȧ5N�����>��I����l��3:��B���]f:\��^{�����v���<w�12x��`:�y�'EĲ�8�m��:�W����(�Y;�S̾ח������(����=�ն��ߊ�Fr(yQH[�ټQk��J)�vپ��r��ؕ����za��4����Ɩ��\vIl�̂�d��b�;w��*v(m��Rr��WG�ms�}�&wgmn�(�d#.��Ȏ�6L�|_+�W���"^Zh�w|7�3���LD�G��,^�Z�k/��c�����ˢR��:�Y�q�����N�c6R)ӯg)�G@(譓hʈ�(�&z�6�])�US��*��"�6j�x�s�<K��zư�F`.!��������T�0���� }T��a��G�8��]Lg�դWH]폑�;9v����<0^��]b�
��욁�^�EiF����ب:@D����Eb}bl:v:,���u:��o��DeED������!{�+�й�ۜT��" F�[B���^�N�8������ۈ/w&���Ջ��ޫ�D�X�Jd��%��0�������S64�#k×[��:`���g�{������1���;�Ҋ�;B1�ek���5ڴ���S��5��wu�z�?ZڔӃ��5�+ᮄ�Q��;��pʸB�M0g�f�Ҕ��XR����[I̫aKM��7�g�
�1P����i�f��7���7LFb��c7
Ǚ��u����Y�/t������'-8�2@�y,ΰ뫢q�&�G�VL���� 	��5�Oa1bV.�Ƥ��q�gb��z�xGL��Ή�\�Ƭʷ	�=@Uu�]GC�N]��h���� ��u&�t�o�������wӹM�6֜ϥnS���7���[�^�Z×���ڣ^ǥ��P���X�sdw}�U����+#+�=���e�_'�cTv�*]���\�%�y~��X=,����uh��'����>v�������9���K�\��Ŷ�t@���OVA��簚���*̧F�w^������)A��^W���,{�SY*x�,��[k ڼH��Bf�u"�}+���'V�
Ρ��g^Cqh5m6��<��u9�
c&���չe˟���7�+Xu].��R��-�a��ri�7��T.���r��^>R�v����BK}�%쥦w��[c[o���7��[��u-���o��.6|��|W��Z�u�O���B��/���y[&r1]sq�L�΋aU)��.��K`'�ò>�w�g� �u�H�J�V�X�H\;Hۼ;
c>|�Z����#aL$w��(�"﹖;&���.��Q�̀_�Lm=��^S`��[��}F�=7�7��������ty(gJ=r�(��R]d�Z�=\�+�ǲ龕Ek�5;�w0ܚ�v>C; �K��������x�v����W�ms�{�I�ʗLב�=0��lG>���.H�Ot�T0`3�T�=�n{X����t��j�7��v�\;�kȳ� ��gj�|�Huj�l�7�ћ�o&����Tc�V�[}3����65؅bS�<�_E�.�>�Vߧ5�o�$EN�H�_��3k��ک���4c]�Sx�.��^�^��{�Ǘ�"�Մ��!���z���2��']kXr�AǤ_u�:ws.��jU���}�T��5�}�Fb6쾊Т��.~�����\V�����{{_�t�5^}����,�Y3�i�~��R��D������_�V����{u���ӚLA2r��j����s�9�����z�]*���?;n���n�o:���N;�A���05���Cij��
ci��6Z�������v�_��{`���.zиL���5�_K�F��'Zw��@SU��c�s��d�j-<>ct��N�#�8"��)��XG���oטL�c0i0�7k����?s�o��]���:<cYduv��Q-��s�l�j��s�cW]\�og�[v��8DA�X0o���xz��V���<g�R��;��<�I}[HC�z[��Ycm�'xu)y���6q�'�ec�g���p��b6��	)W���i=�3���+צ[�4e{Ȱ}�Zg�ʋ�q���.O�?d���H�1�ܮ�y�.�e�1]�oEo_k�%�Ս�Z�����)�%b.{{%�z����l*>U��=�.V��/V{�
��݊ی�.��aH�.�9�ON`�[:���j�0�;��8�@b㼚J�v;P����7��1�Th���|�[��.��F�=�jV����jGR�<}�61�as:����/G<Ux�Q>u�k�yW��A[�^�Oj��x�6�u��lމܣ;���t�>�8�r�X�Ѯ�3u�xb}�:DZ����aX�f1�|;t�p�ǌ�
�_�|��^� u����7C\tŮ����
�7"g�i'mFL���&�Al^{��V��^�n���\�X������݆鮨B�
����t{Լ�}��N�A�m���j�Z�f�Ja*	l���X��ݨ��$��餼�!=��Y5���Y���id։ֽِ���p���Q��PW.Ю ��0��d�Z�{�{�֭`9<�t��Q�ykU{V����w�r�'���c��B�}x�C�(�o=��e�9nW0^E�j2�;L��O_!�͊^/�<0f�~�ݳ�z�$�ݣ�v�&h�xD�b1	�]K��k���'�b�D���c��S�^T���.��	s>�A���:��szbB�;]�`�"�蘹+>��!��E�]Ԗ�?U�7<�ʊ���w��2�w5��^�;iY���л-��˽�Momϫ �(�[�'vm# Jʁ깋�1k�,�s����|�^0�X�דOmM��������� �[�[XD8��s"�[�~wE���)<�9���-�o�):n�\e{NU�,��io�����بo�w�>4�����O6��Ǩe�>�T�!�Y�SAy営��˫m��<<��U9��)!]'���׎r}�����fU�q��^��5�;w�oۉI�������O��܇��"n ^�u��N��<�	���z�;Kg�;@*�@N~ȷK2VQQ�P�}��[0ٓr�Y�.�2S\m^O�gzL�c��C����P���/UJ޸�Zz��8�Z~���<Z=����u������5��#��`'�7Y��{�Ǌ1����׀�W�����&��7Oz�R�*�%���V�M��k�@�Y�MNYv�8{�:�W,w%�9��w?v�uy���$�Slk�!J_w�
��*�y��jX��cW�J�8x���-������'SAch&������/_��{��nx�D�h�Rz��.�2�\�O�b�/W��zj<�jӽ���GGS9��p��v�[��U��u�%\]�u�\�/7���4�&)�u6����\&N��_y�7\.��?uDMϫ�:����bUr��rF�//4�˷�+��دy.�����ḤA�_��ʉA��3�"�����,�.��F��ץ��H�搞;�CWz���*�oVQZ
�p�%�'���+g-T]a\��7�o��=��R�2'"3���17O�{�9
W�LsKt���۾2̧r�`D�Mv�U)�+������v�w�V���a]�T2<���b���%��W��n�e�Ur�u	���ض��.1�{nԻaf̱H#sze�Lj�k��n]��Q�ٷK��[* ��� �<)K���π��Ru첖)�����7��'�=49�f�-��VJn��_/?��ED$Gk�'�uIz%(�jO/�klb-�.����[�w�G��~�u�x��`Eß/oO�G{w,c�e>=��.=�6�:���
n�3�Q]������Asi�����X��˹c\�� 8��P����/�a����N��"�n2��eD,H��y���ms�ŵ�f�Ǯ�udc�����}�;QA;�3H��q��l���*��%k�y�,G<���C5*Ԍ��h4�;�ư�b�=��険L�s��-��༡r�QJ�b��x�6�h,nSc�ٌ�̆��
�rKx���������:�|NC�}o��:oy�	cAF��p��<|�m-���]SǺ��^��aP=��J��w�W��*��0��($�2��wut���;q�mL�,ٖ�u�M���U�wB0��\YM̂�5rkЋ�Yc:�]���e]vnZc���U>��r�
n6k9�
*�Uf�nr��kf$��s�S6om�ۥ�*��+n�Ӹ~��҃L5�J4�X�Hh�S`�L����V�f�MZ�oQ�mʝ�V4J r�4SW����O7����{V��I���f�
<�e�뮥'@D/���CzI��k�<G@їF���'Y��G9�.;	r���2�f����Q}]�gf^ݍ�l*���P�y6�[�FF��=�����Go6���9p֧��vd�"Az(�I��ܭ-�����!�{��"���\��q+�C)��9�rޜ��(i���2���h���mS�#r��!��	]�3�'�����G{wW���,N�ǵ��u����-+�fު`;��ǻ˹���Yg)jYL��;s���Re�m@&Co�jۻ<Sr'J���t�L��s����]�||u<�������g%vNz�L��wZ{�l؀�Rȡ�m֛7+�T:d��9Kr�{|�nb��v�^캝t��%��L�9�ɕ��6�M�X�P�(�3ӈct�kw��I��@%&wRv����\��"�j��mG��vvݷd�厞l��,���k��w�s�K�9����+��Ǚ�#Ws����4�Ӌm�v�[\6�ἕ��!�U*uv��;$���{�W���'���}i#u�Ⱦ��j�֋�����ҥ� Ų���̋���Ln��M0,�������QGX�:�n^���8݋o`�C��ǗH۩j�뙇�./Q ��oE*97L�3h�,�+�tW)4�&�,{{�3��!�^tշ���-Eb��<�ǧJ�(���g+7��-��.8������Şx$��o,���ᕏ�9)����z���Q��/��:I4�Ar�>Ϝ�߀�k�̴�+s���:8�2��`Z�s%�9�d��� �� ��ge���3T�LX�OQ<C�l�J���H���#Uwmv'R�=(����
բ�]�J�J�7;��oY�e��KYLr_���ۏ���d�{��v:b�՛W���n��oX�ͤ�ih�h	�{M<;g����u��Z��o!.�F�`˹8�>�C�h��^-\a�z�u�8JB7W"���*�R�W��K)*W�ӝ�=����,N�aM�f�P(Y5�õ�y!p�=�4Xid3Sǖ��G��W�Fb��Mo /M��Q��W��
��F3�s`�)�葆4fT��"��'���W�u�X�T��.�Š>7��\�oM���oR�����9ָ���#r��tF9H�.��w��D���\~<��뻒;�����7�d�EdgK19_ cs�v������쩖�V�嘘�w2���@hI���,�'$��Z�R�6���]#��dEr�f�#-B��$bʊ�#3	D$ژE�a�D*���$R"�5 �4ӆ-T��dd�$JiRg#,�.��Qe��s��FZQERVA�)-"��U!eAa���T��M��YQ&Ra�r"UMC(6m��uGJ�"D+��Y��P��e��r���E$$UR͔*hJPZ�r*5:+H�Y�&��ABf�TP�B%��%2�HR�\�*��9("�Ӥ�*[12H�H̒�bQb�L0�E4�,Ӗdk�0�fr��ՐY$DDZ�q*��B�%QI�h�U�E��+�i��0�NI�.$$Qi�u"$
M0�QbQ	,��H�Ur�Ef��$%D�0D�$�j�)2�iG)"�D�B�pĉ!*%4�評!�jRHt�,�(�E)I%�\�L�S�ȡº����e<�#�c�\v%5��i�C�R��G]���0��ySw����w .���,�kJ�4���{�����|�W��MV��4�4�Nw��Tk]�1�~4����	�V�f�j��tƥ�D�?9���p��N��9`w��FEs{մT�6�0�n�ʖ>��$_.��|�c���n���,�����]N�=�F��5;^��T&x�V#Z�-�r�����v[���V��	k�h����V�l��>��������l7L>��Uq�.�wC��,�x̕|ר�Vx>���v�%��H괎�L�3��<�/<����ꮓ�[
�>[e�w�S�7��{�+������Ed㥬�lJS����6�}���m[>	�B�w���lv.H���g����*�S�euO�}�+kp'�m�P�'�v����4gy=�o�����co�(��x�ÓJ�=n�;QI�.� ) 屑5:����Mʕ���5����LoP���YYJ�O�6V��ݮ:vt��9ހv���"�v(gN!���������ZrV�bi����m0�l
��e�U�m�wZ��U���N���3GP=��1�7�������� ��>y���E����ף ���lE'�N?l����c�5oK�������q���Z��|�5Go��������̡o��YPN�cw��T_���J1p�TF����A\�r�Rםޞi���z���bm~�Uy:���)�sCyT5�k����fs���UJ^\��:~o�oi��n}�΅�_��o���^���OǺ�8�!���U�\��"�G�9��_���E�z͖��-�D�����Vױ���3]�c�7�c��x��;��nv����Bˠ��X�t�s� �ĤdN�3�^Z��v�i9���e�H㲊�w�	s9(>��PS�$k�Y�/��{S���I!�I
�3�8����~߯��>�t���UW�}^�k}�G�(r����*1�6�_����[]�z�b6|>�˲6g�����ĕ�Bo�ٱ}�u���6�w�څg�B�30^zQ;�8k��^D��v-��%fm{��.W?��<��PM�aQ�P�vlE�#��( �����o>�]Z0v��g^�ٖ3����^M�v���:$�Z��{��:��N�<q�*�uWNڷX���0�^0���{~Sj�c��#Iw��c6k���qc/v��+s�]R��)<��,amz�FRt��%lT+��X������r�<����G>���������e�<Re�"
S[ �|f�,�\s�[ߟ�>���f�߼��ƻ�=%�5�:733����j�9Yoѹ�۽.���.0�#`���;����_W3�bN�pi:��J������C�.�J�#���s��J��4r^���n�W�m�.o*�PɞAn�_���I�6ư�btb}�6D-�G�̬ӥ���r_�[=U�ȍP�P&wU��ʶ�chs��f:+wB�u���R�m.�)[C�'n�V,��ʌ�]��Z��yJt�<y�L�
gr
Q�I��%�^]}����uY3�{i�6C��ە�zb���c����)�⋲Z�v�n�5-�L����G�ᬺ���<�e��^7����GL��p_��u�]4��
��o.SoҐ� <'Iu{F��Ė^t�ĞJ���STwGK�c ��e�v��#м���*�ӨiC�����̀�s�5��N���+��&�@w��n}Bu���B������_wo$�;�<�����Zp�W�\@��Y=�D=��9�"P���om(�O����5Dׇ�[I�,T���!<t!�}i,b��Չn�{�jߦ&��_{�z
��d717�o��=�)���̊�Jٺ�de�z����Q:��ԕմ��������a��ki4�:�=�ݑs���c/g	��(b�.���j$�ۢ�R�I���ku��Z�aQ����f�,��P��ެ�'m�\)^ޟ��7r�������w�&���u^Go�f�����ؼ�m�PuJ��S�ސC"����gY9F~�o�F*�c�ޚ�/�qm�R;��䅨�H��٣w+��٪ �R�Jg�{7�l����Gi�ɫ��õ	���{ 
����{�5�<�ҧ|A��w5���Ix�|!2[}��S����<x�;{I����x�2��gT]��0ޠj��]�ݏd<�v��H�{�}}��L�;��H��J �*�6��3�����Jf������fn��2��dɑUxJ� ���+u$��ڷ���SB^��o:�K\�Iølk�V�rR72�g���B]ס�9��� ���S��m��x,nWn����Bҧb���>�f[�}�\�ԝ���b����(	X��uZ�F͙0���w�Mߎ���M�f.��p׆��\t���}R�P�[@��ƶ��M��������}&�NR��b}�����tt�',���=���_���C��^�DG�Sw��8ZNrB�2�����ˁ5�z�z+�E���k�s���1	ˢ�K�����1���3ؽd�}��`��V�}�+{{S:���\�֫q\�������N�@���)��X�H.����W{'������9ʯaklԺ$��L��q��i��b���d���%�|�I�2t�r��/j�a�ٱ`G�ptu��^`ML�
��\��[���gW�_��|���VnaD���>�6���Nz(M������3�nD�v�#�DD&(n�׉���Gn���+�K�S�U��/rV)�9����ݝEC��U؉�k�O~����x��|�g<��k�g��������b�`Cz��)���k.U�����E�c��Ӡ�����X͡l\��t�A�~��Z݄H��O�����Gj��݉�z�V��	��n2�.�U�n{gT�G5͇�e>ބ�����>-m�ݎ+���^���;Q���k7�xQ�^�{��w�����"�����A$���s��W��������>�Y7QN3q�FąJ$u#� ���V��j!ʎ.��N�����ˀ{��w��e.Q-65�ؐ5ى�>����r2HE�����f��^/oz����q�駡'SKr�7��ٍq��DW��W�I4�w�y5�E���#N�_`�{Cr�߹K�XsO(�;��5~�� �pAX��Gw޸U���u蕑����\��e�_'�cTu����ѥVؕ��W�w��8.)5J�.�/�b�6<��(]�2�3k��X4��r�1�#�<�~�gݒ�wOTk�f��9w(���1o��Vq�ɵ��Yl!�����Ʋ��z]�Ԭjìv�WQmC�Ȱ{z�<�<���`,�5�y����q˝]�D��mY�]���0��{���b̠�������_O�ҵ竉L_�cŶ�?�_��m�y�&�W�O�[n�qG��}�t�xy�Y�~��æ�®ݰ�*�ò�AV#Q��nQ��9�w��Ry�?Yn*�.�m�s�8)���UV�l���$:C.����}��R�O��1&����Jyio,a��am��
o��*-ŕ�b�bMyt��"hq}�%���Eץ-4I�0�!�-�o�&�]�5	9��|'�αQ�?k�*q^�P�ǖ�Vb�(��μ<�!�]�w���w�0�G����D4�(O��؛@������8<�#���G����7ܐ�J�j8���Gm�ٯ��z�M�_u���u�{)1IOo?gq��|Ոo���à��Uˊ������'l�*+�.�[���{>�)�ӂ�t�/]��u�M=Q�(Uƕ��s���=Nݷ�,kι�ޗ�V���.h�2��z�󃽮�42)�:���[���"vy�l�;:�R���w�P�pe�s�-XF����L�D�5��S��;�wt ��fTk�����d�;=�{������Ky�ԋ����Iñ�lk�
��=�{NZ�.��8�#� ��gly{�nݿC�9ٗ<�j�m{��6�h,a�&ƻ��g�Dk��:�{��ֲ�Ǿ��J�<�
�E�2��S��*&�H»���t�m1=�g����th�[ڱ��L��� �z����zX[��'�/*jy��c�;^�]#X9��}��j+���O�پi�]�ޱ/��Z��.f)/�{�b{���0�`�o�+���<�x�{�{��F
�����)-����Ŗ1*�[w�M�w��NgR��;���V��o�w�K���qC7����S|��vJA4����v��<e҈�;�9ܗմ�U媕�o/�o1��,f̜�����g�t��%֞��\T)lF�^|�J�O�3Ωw2�;�����jh�Pe�$��ܴ�Q9ЅɮjJ��Ͻ}4tꚡ}���Ra��E�гfv���qTMnG��=,g�u^��ֆxW�M�׆ٱS�%�8�����X�a'#��«[��9�[�Ħ��g;�.�+UYX��x�&�7��׼�\�]v�t������S#���kL��<�g��>r�WǾ�n��<�փ�OX)�_){����^�,���x�f��m��RW
{��a-���j0[��roX�X����u�ҿC�[���[q��f�0���E�ob�l��]V�r�ن;���-P�.;C�J�7����x(�d�O:M@畢�b��u����{\Е�47y�G7�s���b�fʺwc+4����*��*%�h�V#nJܚ O<�՛�����䥺H��t�-�q��D����9��d*���t=<�m�]~N_gz����uɌ��_���yz���+{Ǘ�r��V#�&w��U���Be���>������j\�E��p�s|��z����u�{�:��&߮�w�$��>��!�0'��l�Ӗ�+�z%�e�چ[��S/b�lc��!�e���qL����U�ݝ��V:T�p�g��;���c�<��Q����r���%Ʈ��+��y��������Qo��8x~դ�[�-ku��<�)Y�����#���xY�,!ʷ�+9�����3z#��xզ�prG�­���Ʉ���?��2�*�I������N��+�)�X�BE�讗�Ü[�&��v8�.���ѵJ�ҹLn��
�R���w A�,�m Ո�xF7˛�"]�ٗ*q�O4�l�o���~��I
�3����]�lF���e�bt���*�!+y��C�s�UM�V�I-~t��]�u�U�>+ϑ���e�Yx��_.�x�s�E��}o���M=����� -��(Up��:�j½l���d\1so�貖� ����]�X͡o�('M�\;��ؠh��ؚ�<�������nl���WP���o��[�O28[q���"����[�����,��5r�Eb�/���xS��U�/{�g�y�_P¡e�&%�B�{���iS�Һ�`��Jۼ���<^^ܘ-JK�#�б�5fn���1�;���*�OR;Py��Z��K&E�:�Ⱥ7\�+9�AKiL�d����ͭ4��].ڌ��ޛY��Z�&��wY�Q��׌�o%���{�۹S2�[�%ܗb����!�]��}{�� B�`(l��=C+�lJ�����7ˉt�wd�F[b��T��vw1x���d�[��dm^��w�KPK!�EY���uti��T%�f*�h���۹R[�3R�x��ݐ��V������b숅�PI{�1�������AG�e&+��EX;F3|�X��)Y[{�6\��3�JT��-�K]pޡM'��Ν�[N�-ǓW\�oSt��*a��vw5� �������]������u���h'z:�&�ȩ;Rm��t�Ǆʮ+uH w[w����ͳ{�·���2t!4�_p�uב��im���Y ��.�(�pa���l���L �	U���R%�c���8e�����e,�W���+]巋\��]KK��Y��m��+i��:G>Wv3B��h�B [���e��� �<s+��4�;�s�>��T��oY�sq-��b�f�����4(�֛�±�Ѿ�����*�%�� �p�l���ȯ{��_�����t�u{)z�4��Z{&#nrU�q�7:��qW
�1�dEg= �������i�2���I����,!lV�n��j����{��*�꾈!���3g�<�yr��lJ�oNR&�<�G={���/%f���[�dG��\T�tv���u*h�);y���vT����P���Dj�8�6@��CfȻuۨ�U5n�̬�-��c:��f�ޔ͇�\�[�ktT<�F{o�lLh�D�TF�����]�cŲ�C�ۏf��MtE�A��Z](vv\
����w��V�jr�Ձ�\�V�9K��m���8�o*�w^�����0;��Âj��T��D8Ŋ���D�n�u�*��U�h�P֝%U�=�����kj�D����-8���!s�yP�ʳ wa�[�M���v��G�qI����.����i���=赙MKf��.Eu�����g�MC�Cy[5=�u!CY��n8�=����`V�ʍ!���M�:u\�8��=U�<	�:m�]Kl-��r%Gc�7Z�f�^�G�d����N����wq�D����v΁D�+����[���o� �6Y8�u���n�n�~����C�������XcS�9c�c�7^�Ր�zQ0�	iۮx.`��YX�v�_<�,Rh���.]oCor���ެӫ��u�Ԩ��kwZҙ�*e������E,ٛ��Q#q�AX�����f���J/����R�҂֠��:(TW�F5�uva,aK��9H�^ݒcR��v���lA,
���w	��J}R�����i�m�
 ���輢�E�ޭ�{I�� ���H��L>;����ʗԝ]����k��.�vl�n��.�v!F�؄�i<xaf�+-EQ�B��2MYQa&T��&��\�J�s$�Rr�H�*U���̕m"�YQ��:������*���Tl�*Q*Q9T�$����YЭDŝf����!j�
�F�&���H����-"�"�����9SDӲMM��.hH���-.$i#�QW)MgV�(�Ue��"�9L����F�X�,�����8eaTkhrbZ�Tb�B���-�\��-2*��A3	#3.RGHY���Z�$+�]DC�)T�Qi��ɚȣA:�[J;PIQS�31Nҩ!�aEĒ"(���MDeqP��jW�U�Q��&aSB�C�AmH��PQU�(F$�`P>|;��%z$�A�Z�ܑ��%�v��q �t�=f���ח����9��z8�?��ط�s����! ��͊��=U��Z��.i*�#;�vts}3��q-���
ߗ�^�klE�_��~�$����I�K���yٽ�m'3�XÚ	�v��[㖽o�J�Л��r�֥����=B^eu=}�y�ʷ~�/�kh<���b��	����4�0lWI�'ݡ�+"�˝mL���'�"t��.Gt��d��D���d�A�~3W���Y����j���/�G��.�<�˓b���~/�<�d�VA�}x�o���=�6Vd�ǥ��Lquk�,+�I~���!9�<#�,����s��\�0�$\�������\�e^�8�t;�-���<�7��*�lF���Q�"F�7)k�[���BN:ڧ*ժW���a���-��{aM�٠�r)9�[IB�ֳb���x#�В�_]^��I�0�����Ӱ����U�S�o��m�XS4�𫒪��k�l��Â�������;۞9m���v)z�j$9W���S ݓM�n>*Ⱦq%.�]XQ5ε�峜F^�Ǖ{]Bk��a�3O���*-o,�f콙�V�g�����X�`�u9�yx^�_����I��*6�W|"�ϗ���D$�%��vR���r����q� �C=�|�^�\'�:+���g��2]��Or��+�`S���N�f��&��v�1sQ�Ɉw�w���tʈX:au�'�L�ԝ9
�_,Z�b5\1j�J�7X��k�5~��õ
�;�O&*��n�OT��a�g����=���;[��^�JI�P��b�N�n�of�ҸLD5<�t��ı�F\���_�,��k����M,a�lc=��`�|�v��n9�}@���z�����v/"��#�=�Sw���Lmq���Y��짦F˾��o'|9ٽq�'��B���d��\+��o)���v���뺉�c&V�ƾA��?ٴ��O�OV{��$4l&�
ؙ������L��Mo	o�'���Z��u������� ��L�ͮ�}Y༵7�ە�z�HzT<z�de�5w͐��V�Z��ي���7XzH�<�t�s���� �Gq���y]���ڲ�ن9���/��;^�wH���n!��n։p�"����EYΏt)Aŝ9�s�!Jf��s�a������BT�<�U���s�.��*X<C����%��"�C�����//�eVF�ڸ���N(�~7s�)ק��i��Ѳ��q^���;o��=��Z�#M�J��Vk4gm�����+b6|Z�<�K�H�J�-��o/�5�����m�2�S~��!��]�Y>�rO;&I�&X��Z�Ƶn��}�Ӫf�<���)�b �n�"�J���wD��e���{u@�;BR�����-�r���bی�T��.�����3�u<,�:�������*�ݷ�b}�[J�!ޭ���U�R����b��ٕ�f�O\��}���m�lP��q�9�+�w��;r
;���\�1��βD��UaE����>/\ԭɯn����6��핰J�!E]<ݹX��p�p�o�]��Z����Gz���ME�7��ŷ�K��zVV����Y�;1>ȭ�ڿm5Bz�/�\~��3L���T��h1�%��^�.�J��y~ѩ/q^���/'[); ��X��3k"g��	L�z��AO��W�J���$���uɢ�.�K�t�)֖�3����k�j��$�|��yN�[w��w��4lk�B��vbyGO�ևO�e.�*t�-���`�=WY���9TZ�;`4�-a�y�[��f�k����fA�����j�(V����E�)h�6i�K�k��9�=�UF�b������)�͈O�J]R�6��kj'�2�J�<�3<mS�1�|���wn��
�H��u�8���<���]ȇμ&�(D�b1�ѽ/��u���s�c�g�����9�_y,u��hW��@s�;��ٴ�W¨��o
I¡���evSQ��˴�>�$b��!�gqj�G��%�m P�}5\���k���y0�<<ⅰ�Zm��I�7�YT)]��y��^�_�s�o1k�׆���r��F�ooXk1��Ol�lT,[ׄo�;Rn����3��]��Gې��;��x�`�3h[��N��-t틩��;7�wE�Ş�������w�49�P:�PR���2���jy¶����W<�h��mܝ���/�eErݓ���Ai;��̜�p�?0�-�Mgc}M^��ux��Ru�Wp� ��|1(���F��JD�Y�*n�O�B�<�A�@��*9��⺀3�/�m�py�S�]�R�u�w $���V��1�v��Gg�˦Rء]��ǅ}NzD:�/�ʍ�X��}�ݧ��ndPm��,�F����M�[�b�?W뱿i=��qOK���3�AgJKB�q��z�O�\r��P6�b�t���ī�{YS\j����6�g7�	��b�������N�ˑ[uqқ��z�yPj.o�{���	�v��k�7sf]��n%MtE1	�xFb���O_f���o�{�]y?[7�y�V�@�C{�=��g��0w�f��Z<��"���y�fx�>l��oW^q�ٰB�;75�^���]R��q�@�����8b��]�,��-��>��Ϻ��U�%��(�Z�VU��q�
�Aޡ.p��S�_��w���eJd]�yk�WU��V��ΦqW^"��Ӕ��ZMcj�m���jG��N`l3�]��q�u���,Ug�`LCZ�:	n]�@��!=,N����y	B��S�k��C���j��V6��%���aX�	��wK�x+:�s�������:ol*�����qo���A�/PZ{{�W;�[�ǝ�|��S�_��\%�m��}`{���qvJ�w����5
��s�Wv��������)V�W�-����+�,�=�B�N���=������j�$cb��@�ʤ���EД��I�a����b�M=ͩ��z� bb�FRt��.�oI@�p����ā�D��d��gaK�V��Ot�эJ�K=��y�o)|U�mZ�q��K��;W�"��
Jt���i\;Գ�dRn2�^~<i�bR�B��FnZ�3O�j����-��\v�sA���;P���"���+�dEY����ngy�fu�z/�j���4;S�jE�o�RN�Ь:ә���[����K��1���Յ�e�<�ŝ��mT�a�ۦn�l��oX���e#�%]@�pj"��]�V�RX.�.�5�vc{w[�����iv͹l@u�N�T���*�ǻ&�8r��̥r,�H�<�eK�a<��f�N�m��v�O!��q�KkgWKܾOX�V/�ԓ�W��;k}m�r�n��P/8)�"��-պg������Xk��}U�'�E�2��6b=��]r�{GZ2'����|S����MB�ywS��Խn���&v���Z�j�ָ3o�����I�ظj~����5�>����m;F���2�H��|��~�a.Z��y��^�dT^��>~D�p���n�}��G9E��0	�̵�ۈ:L5.����Nm	��P����@t�n1�}`:���y�d=9�"0�g�Ǜ�W'}�o׊v�_.� ����an+ع��m�1U7ZHO+]H�V�!(�{7�Y�� �<�I}B�J��N�g�T���B��3��-0�ȝ�3R�t�ߔ�+��!lFϊ*���T��8G	yW���:�ì����Xk����[e�v"�/oa@�w��r�vi�[El=Cˏ�P����K|a���vc6ۋ�꒸�R;��[��#8P�R��t��=,var3: cVZ���2�g�o#��ZO(��2��cqܡ(X:��W�N�g+r:fs6n.	_-�]P��l�]s�#����P�kO�k1�nfv��p���P���DM�LDA|z建pz��4L]J��o�HrD�=g���j �ό�� ��u�8'�m�W��<��@��Xu�)k�N��R��=�^
�N��v����u�KB�\$N��E^����U�Cŕx��4���� �sR�&�7y׵#���Nȼ
Hyi���lֺ��l��P��+�*'�� �Ul\GN�����k�ۼ�G�� �h�s����8�M�a�k�9GH�[B�����^��x5Stx�A��u��w�Tc�w�s��P�^��uʌ^7�n�ދ���] �u����"�q�6 �Y4��/o�X�>��nUQ�4����L�7�b�{#�
�z�}U�˪�#�j	-�^�'��N��S^���]����Z��cn;���a�6sJq�#%hq�=����f�7���v�dL\���?Xī�l����_R�^���W�� �y;i���S�}��w5px^<��a��È��k9͘c� )��x�|V%yf
�vFqO1G��1��h�l4]<��݄��V'��P�Hd�ҋЩ�Ӽޔ��cw�r��3U��ej����+��^�`����B�)��1C�'"?xO1���m�Tv���<�j�I}�����s�͈:��y�rS��P��	���=�7��*�b6J`Ј�+�ʔ"[�Z�Z�/�����ؤ�ױ7��5��-���*۸�Fj�(K��cC�jR]q�x������t%-4
O9�Z��3k��2�>:��$��k�7��:�q���|
B[�WBՉ�펵�������"6p�ݫ-mtȼ��=<}���o� `�`�دGn��8W����-zI�������{�m�y2)7��t�#
}��6>�������&�dt��������	��p�ð��T�}Ԏנ�N�R����SϪvuK܂��k%�f�����M6ƻ�buщ�k�@��5J�w�P�Eg�z���,���A�괓�Vl�sr�S����F��WV��\K�0�����FWi�53ĊS��=�̷�<t�p/lu3[�!@v�V�0N�;.-�˫k�:�_͉4������E��_*zPX%ܳp�H����� ̷g8��w3V��N#�
�Լ���0;���Ф\��U���K����^���?*��[�^�aL[�.�!�F��n���7^�|��ݜ��b{��գβ��G���oJֽ��*��i��ok�QQ�}����ל�s<.�臯���[ᾗꁷ��.���)�3�������{u��}�1=S�|xa��'� ڼN"b�����v�#ΟK�ͥ��<1_��q@r���7��]���;ˎ��ג���]�wMh��Q�V�,�.�EcL�x[���	���ڛ�CNu�5�MMb�<q҈��<��yԞ�T�XV�^��n�0�4�(Q�V�;9WY����L�޸�R؎��ӫrF>c��"˓��0lz=���/z�.���`�v���P����6|��O����G�3ѵ$�*���4�L1rX��÷ؘ�v�ar�#
G{zA�Kc [���S=�`�(�ɛU�Ug-`�\�U���U^J�WC�Ր��|Y�StK�سF�
�"�5�2�6�G.`�:7Y�ky����r�����X��܅�9�*I�❢�Hh���@r�.������;�x$�3�\v��J2�ެ&i�Kۻ�U�&!��|����h�H�C���:��E��t�W��\���ݴ��Nb����=;���m���-��'�ڙ�ԣ�j+����.�Eb{ ӗS�D�u��[sg�2��:��m朜(^8~1% �0m`��ս�{�i.͓�@��u9�Cai�������S��&8����;��˫̕h��f��I8)����;����͕����m���ۃbcTOd��$Y�t���<����wA��E�}Egu]v d�l����G+%����	.Q�0N|��@;�}�Y���R��[l��-G{��]���X�^��b���g�dRx�Y�2 �.��h�ɻ4����G��n�sWDA@�ɧ�`�q�"&:V�[���9t�6˝FX��41bN�x��8�*ɼv݌�ň�8��K�F[�F�U��}Q^	W�(wl��wk9g<"ֱ��:�����ևj���x*��\��S55n��X��A�P.v�O\��WTWMꉩ[�Yo]kծnuK5��Ch�ej8�z��i�i����|Cu�2՗��M�[oOeQ�������Lm�9�z]`V:�g��S6�-!�u�a��^�:����W��Y4�X�70JJ�HJ�8G�+%d�f�/�̀���t�bmU�2��<%�C9$��y�Y�F)R��Q���h.O�hU��L��ޔ��G���ֽ�|u����]��7�+ \���v}e�����79-<��I�T���6���]�Ҳ�ճ�Rt,(cE�lWvݹ�����5�P�Ե�9ܛ�����W o`���Ty����[����Yb�u�.����봹��L�r�uê�a�n1���G2βtoe,FmI����]�_
�7�eu��i�:��R ���Z*I�,�j��B�]r@<i���[�]Ĕ��(��N���4)ګz�hH�|;-���|8�q�dˬs�eM�G�]�;1�V�;`��z�������tٙ�����X�3���%�q��f�ϫ�p��$X�I6G��ٮ���y���g�:ҧ��C'�K7'A/2j�L��ݕ����ߢ��2��.��v�<tޘ��ö]HK�Z̓=��5o�-�7v���6b���P��p�sV:TlL���a|e�h*Sw���xruւ��[Wt��Ŧ��},M���=hE�B�k�.����R�ť��0n�.�FM�͢&Qݜ���xrJ�YOeЫ�E�a�����k.�Ҕ0�\��xq��\�[{0+/�(�ޙ��3�G�TW��wb�Gݥ���ڳ�p���_;��_���)� ���5i*	��L���S!#	3��Tf�DdY'Nd�EvQIЪ
�9�����$KXW(��(��
εZV�*5	$�EFl��"�9!�PQdiˑIP���VD$�UAq�DU�%e�\,0��Rt�H
�UD�9ʢ�;"�\�Q̑D�E�*Ùr"�E��ˑU�"�9AT�0��N�®S(�U&�h�U�G
	E��T'*�r�Q$�
�Er��")6f	'iĨĥZEʈ��(��5��p�+��dvG+F�u�TE*(�$�sR���R��9Dv�ʂ4��*�S"��B���\��Ȩ�)R�2�G4�#0�*ȫ���djA�Q�(�fQ��9Q̓�5
��-�\�H��tȃ�U�j��&\��eW3.�����G��������n�ataE�N�\�3K ���	���M)���7���
�k�]w-�V���WN��Jb3����j�u~��CwX)�jA��%��5�t�ގ��@>��}��|r/��ۙ!|i\��w�wo�NToj뀖�|��
Q��%gr�WT'3:[]�hF��e��R{n}�ʳ���g;�p�CD�/{�8]O,'r�����ƺ�܂�2��ɫŽ��6�yw`v'���oy�����}�+L�����9��f$s��b*=����E�S������}C�\a��|�o�m��.���9���͗u��Ok|���^k[k�`a�Н��ԧ�Bak[�ς�{~��5�������֡�맮��!�­�+0j��}�0�L��;P���S<�c�]b{�e��wY�̟ �r���zM}��ϣS�	�ʉa��!7ˢ��|�e{��=�$u��6��Y��7�M��ӱ��]ȃ������j���㗞��l
Hu�����H5H��.����٢@����A]-AըV�w����Jf�a��Ty��f�Vy�ش��wmcr�s"��v�+Fmŉ*��R�.�'^��JU�n�OJ��\kXYo�݉i|c��B�-"_����4�i���#�(�W�>���
؍�yϠ�%�m R�)���])x��Iꝣ�UE�t�49[<�#d��ʄ���F�v.�m���&�!ҧ��'r�6�ް��0��o���b�`^ސP��1�tf�3���v����d\8{�a�'`K|a������fж�(T���`���]Z�o�L�K}F�́�i���k��V!޽��W�޳f���5%������0f��c%��c`��١+^t%ظ�M+�o�ձHiȺ�\�\��o����Q�eC=������V��+rkۼ�jGF��3^�˜��dA�Ek۫�ĩ~�R�ҕW.�|q��cb=���Z�����ߡ|����~�)��_�7`~�rQC�=vb}�8Z���LW`Ggvg�h��\R�w����a']kXsA�h{�=��R���T�T{1v�
���N�ȳjh�հ�˩V��y�8�iǧjIW��D��'ˌQ�fN��>�S8���7�%AM.��3)em���wc_��t�>��)��R-1u�fƘ�b������[��]�B3�e�d�9}�>C�VS+�!V��s\P4H�������+EOO����^��9���;Or�ps*���{Fڼi2�O+��Q>:<��a�ԧ�~7|�9����|��;�p �'J�+ԙ�@��S���ߜ�ѧ��zث2���=��3�L�=MO$�˷�+�.M���b���8���l�dx�V�_.���Ʒ��fR��rŴ�<~B�Qq���\��v�9��b���hV�l�{��Z���2�w�)�k�V���X��t�in*�k-6��t��\��U���C4��/6.^���8{f1�ڧ*�)*5����5��-�&�¦��9f��,T69��>c�_z��[�����H�1Eץ-4
O/�5�5�҃���g8�
3��FO[�Ͼ+�X����}"���0�6g�v{�ݚ��<k�uq����U9^��n`�Hz�W��l�@��qx�F�����hR���s7xͰ[*��en��^��-jY9Y�h�Q�[�����Au9�B��[u`"hWB7F](Y�5>0���ϳ�;�,���rt��F`P[���={�>�Պ�j}R�\��s��w��Naqc�n���+;�V:�tj�C���z��gb�j�9X�����E�4�����^d��f�Y���/����-;ԩ�=Տ��.r��hC��6%R�}1u����;p�A��w�'��ַ��N���{�6�e�I�כc]��raC���#Y����9iq�~���m�v^Ky4/�uZ�����9�`��U�^��w�M�=����s�iz�9~��V<����[�z�E�i?.�xxS��▂w�ݬ=-�v�F˾�����y����;bz��G�d6�����fq��喊�]U.��O��5Gkms�<�g���0ާ���x[�"���L������L�q�֮��u���/��;r��Y��B<�����]�T�:X�C�
qC�7?!9�<#,�2�|A~�Q��C-w��Ȃ��%��	p�-X��V �XM���?+���&n��{h0���j���1'x�h#�\�.7���>�EL���	���.�D��Ou�Evh�C��a���ջ�UX���:�\����{�5㲩�ɴ��6�k��o��k�b�̜IY��u�z����i�3���3�k���Wbv�U����������Ꮻ�ڿJ�n7˻�@�l7|1��!h�yܻ�K,��P���R�o��B�-�� �a�%.���E��<hdf3S��S4t
��1���/|���p����
Г��J��k'&�}lJS�6����
��!x�m�T�F��=��!����o-�1OYŜT8Kn�/�ػ��iX�z�y�I�����l5
e�$^]A�Ny.�ZGwK��C\1q��?�ݧ��g����K���G�)���8T�\cF����vY�=N)�%ؙ��'|`��G(�ɫ���\�.�	)d�O���uojs����׽�Wmp���<uR�Y; ���_�*V�a����=�M�<�-���}�=�TWo����fu��HM�`ip���~�������0���a�������]W�j�n����|b�iq�\o��w�k���
�'������`���c�NԖ#�c{s�q�X(Y�Ag�7v��O����X�\=�z�MYT�w���rǒM����^κL�h�·qέ�nA[&�j9E60D굍tR^��K�r�ܢ��w��Z���T{�`�&(�e4�F�B�'|>;K&����W�
8�P9����o��ş�Oy�ܾ�~U4�ǣ���Sꨜ½��ϑ���NV��W���E^��GWc�P��}G���N{���}�c�
���8��ucwϯ8���?o���yj�y�/2�v=չ�M��0�wl��h��Y5��*��R�=��u>~`�;����09������n�!]��/��.3��M�d�_�ax��
\���@%�T^�-�
��f6�x���yo6��_�g��]�w��Su�m̌��N���ў�We��@�T⼦a�N�I�ȗ���W���������^{�}>v���ʽ|�%#���2����[�H��̋�gW�,��=�������S�V&�R����2��!�>�Z�/��hG*�rg:X�e��?�¾�t#�\��C�޺l�)��7-���dx�y�����Q�̥N`]�~�1�N��e�@}F@ـZ�"����GC�����-�C�_���N�I���ہi�5^Z��n[n�m�(��D�'I��y�Ѻ+K�}ơ,]r0o'��j����Qxo~"�_�Sͧc�-{���ٸ���cym�v�t�e�I۬@��v���FYsw:�����g!�n�+w��Koͼ�Y#t�'�X�vr����ћ��fQ
��C��@����n���BBR��kA�J���	��Z,r!>Ph�3�iKn|˷蛅2�z����&VӣqV��ݸ�qn�ݹ�MT�]�}��\s�vڣi��_�:`~�*��@�tڙ�fe3g�¢V�
��J�4�@�cT�B�/9EQ�����\%�to��l�)�|P��s'�#��҆����t�f��n<>��R�࿫r��d�;����y'w�=\S�p�P�����:�ٚGs_�2��-���6�)�ѓ�mOa�q֫I�}�H;��w�Ǿ�O}\�s��X�KF��˔����Zo�S�"��9A��-�S�f�`9�� ���aL��LDJ�8\��q]��Œg<:O綷թ���:6�F��%�U�]k��;o-xl�Z����M��H��_V}�@�!���)9�]>��p�s��yӒv�Y<2�ex�ڎ��UƳ{ϴ�t�N�⎳�@�,��v1�&��/s���y�\n���/N���$�D��&j��wv������c��ه�K��N�/it����L�uWT,p����G�eXO<��R���{Ҹ��|=Re�XQgv��I!�<�ެ������ Y�+̄oJE6�t�˩7J�F����e��ϯw��^E��j:��h�3wU+�%�A
T�ŝ�%.�;}8n-�7n,�}��3E$����z�%rXn�k�Ǵ���f����A�:�����U��n�R�JhN�'lh�P��AMT<�ng���x�N�K�1��t�:Ite �(�K��먗t��H������h���eGg��=e�Y�{�q����>��" oW�a@��i6O3��L���Kߠ���~�/�8:1��.���<������R��h�n<��ꐜ�2T��@��.H�J��Z_��cj������ӎ'K�n��m�E>����Su�K�fQ$��J�Hsu��Jpc6b�ߺ�W9�W��:��<��8��f��tS/�e>d�&��Sl���\��G3����#�ߐܝg-�u�c���*''��qJ{_ݴ��s���]ы䝚7ܸ�Tz=�ɷ_����|}8�����x�>�Ln��{���R���)����I�P�:��K�l�U�c��ۺ�������{�O*A��D�L-��c�)�a�+Kލ�cE���ت�tY�隟efP{�4��iV��Ay4d��A}��H��J'*�L�̨S�|w�5+	�ky�������8�� ?mK�Z��ɰ"a� �܎�c�>Q�k3����{EN��]����e��{��U�=�W_�r��ڛ��h~��o��ԗah����J�ҾS&V���d�k<�Pޛu)��mt7���E���PV*ջM�׳�(_B�+�k��=g��T��G*c�����v�{E¹��^�\���WTT׶��Su�>��o�MaoI��K�Q�}p��k�d��{��a,�U�ha�&v/��:w���:�~�=q����hy���S�pY�C�|rPxU�o�s,C�l����;�aw�m )�צ3]V���yv��4ha=��W�Ζ.�_�!��|���P��t��dd��WW�e^	~��+]�J��Y�|�e��Ğ�d?�=H_�3�on�^�yz�/in�l]vy�2�������t�*��@v�v���z�1D���$�!���V�b~3c�z�����ÿozFˉN�>��5;�t���G��a@�y���P��}�eR$O�}�k.�r/mc8�*�q���\K�]Ǌ�g��'#ߛ�2�գ7
dk��<n4Ϸu׽��p����:�6�C����7��w�;H�w���ĸ���˧v̎�\q�� C�\ꛇ��幬�rH�p6�!�����9�2¸��#n9u�����Y�>D��ƽ(����t��Z�Cn�!���W�2j�K�YJ���Z���s�p1^�BR�v^��8���kl���׺�F+��v�:��>�4�x)^eݱ�ÈVT
��v�K�v���������&Q��k�-O����[=�]�)l�T�z�_�L~��l܂�a��'|b�m:7Wd�l��uHa��t:yA��׽~�5��͛g�VM���k�W����������T��9G���T,=�eL�: 2E�[���q���9��������@:����ই�5��,��|�9>
�f/�������w'k��u�S)���v�Xy���G<��ѷ�HV�=���o6X<G���1�s;��ܹ]�`���[�zN�Df�f�r��2���'̬��q;p���g��O�.>u43���Ŭ�̝��	��@d�w�O�࿍u"s�v��<��ǾU\���u�������]8/�gt%+\O��~�*Q��d�ِ��..�kM�iP�2��W������������]���c����N����y�S��{��/vaz)�q��� ��mPaR����f jߊf:�sP�����ֿa����c}+���]�#n.t����5z�]|}�����ٮގ������@�_f������c���F;��}�1�n�(JP�A'j&P���g�G�ȵ�w�V���p��7&h��,N���.uE�p��
�cBU�R��d�5l;:�j�1�{d�q!cE͖��j�G�}}�7�ߥ�
m��8��@�eK�٠�*�-9׹+��Ӫ1K�+�%�JgJxRqŽjo���%'���.�'����Ҹ�*�+�[j����h��j�]�u��S͋��C�:c9/vZ��# -�6��Xك��Εl+�&5'��ݬ������k:	\^�����$��ܚ71�y|��w'O���3k��А*�r�����gc��������(P��Ağs�a�i�s��z�p=����f�������*��U��-��·������٬q�*'Pd�a�:$��!ܑc��p(�.�����;�_q�Ka6��أ�v޺<a�E
$jʳ��/�|^�3d.�Y�MmƳ�V)������z*�;���<��Y�2��D�0*�*jht������;YVu���z��"������.4f��Q��	�5�w]��r2a�{��s�FK�F���d�}�d.��{1;���(���W's��O{�mJX��x#�{U�kKe��e�&�W�jPw�q9�;쀋|��&�-C��b[Q&�F�;��w�k+`��y�����i3`鲻"(��wXL]8Q��+�����2�pHλ�³gCA==�  �3|P���i�˂��v�q ;,�z��o^�kl6��LmR|+���n�mgw\эc���'2������YU+GdX��Č���$���ϒ��u�]ݚ���(m�-][ֺ�Z
���#������q�ś�C@l�0�]&Ԕ{'5��K�4�R[J�t��^�}��1����t�� =�X�hڻ����el�9P}S$���w@1o5�̸�-�)��k
�*�M_��l�/U��^�M�Uv��y��3�:��彙����P����g�Z���!*�wAwa���,�&)
�/��զe���l���F0i�(�P
��\��R�j��=
��W���Dŝ��lGfPK2݃{���X��Y�����4(�}�^ͧ�jWo�*wu����)��Ro�D����/�$NnwH�ʻZ�T\�&�����v��*b�'3����+h�\Q�Ӱ꙼��VtG�����
�	eL[��C�=NQUpB�|��3��
ا��Ju���ky�4��l$}[������{,Z�R��	qWv�;)Y�.�া��d�ä
L�tŎ�C�&�W��X��Y6O�j��V�f4q\���I�amk�p�C���LW�hR��յ�i���kq^cϡ���r�@]���Z�����r���)�K;Z����`]'[tf�kUIb'��4���R]mN�ʰ[�s�9i��&�ή�w�������[-��d�{�ʵk���7f�MV�qV�C�J\S1Ij���m�E�o�u��.�w�Ύ�"��GC�Y�:���PE�GL*�hDEI�p���@E\���(�,��N�Ȋ�� ��ʓ�UU2̮QDP���(2(��3���"	����"��""�������A9���DFI&QfDh�VE�+C$��(� ęʪ+�UW �I\�Zt*PH�D8r�Y��"��T��s2*
�U(�B#�UE�r���+��I�@el������s�QEDgH��PB4K��*�KYr��\֐Er'&�4��Tr���\#�QW9E]X�L�H��U�� � ��P/+qШ�#�9\��ȉ�Yq*��쨹�*�+�Uӡ˜�B̨�x�I5�TQW"�PTY�Z�TU�16k@�*���N�I�PEUp�fDs��Dp�#'9(�Dp��*r��2Uѡ�4�Hg*""���o뺺�%dQ�5�h.}�F���V�&��Z��"��f�d|�q��m��lk�ȧ"�8�j#����^��ƙI�b<Hs�6?T���u�vi��Y�����T��F��>�rۏ>�[��̿} �V0z`��W���[)wd0.A�"΂��燣�t��E7\&���r�k�k��o�7psۯ'�DrDMbV���\��c�tӂ�@P� {6�������m��TϏ���c�{�=�:�����+��╻��FJ5�@]P'I��u�n����ơ+�C�����_�X��X�H��=�_�Ŵ�p̈́N�� �v�je���������O�9�b�wO���c�����3��k}N�jt�:`~
�W��.�O%�QKߌ���큠�cV�񻩕r��Y�Z��h����o���UG�d�MM��P����2k��1��S�����f������;�XpJ�B��e-7����$��B����%@�N�E�M�3���PmԾ�}��/�IU��+��^�Z�'se��~z9S�G�k��S��V�zŏNP /IZ�o���L+*�p,��ڟ�Na�>��M*�s�v� g�S�>�tI��jf��V!�Tl+%ߦh�	+�J���s�,_,o:&�|�u�{y�
1�T�9fBj6ڹ�c��̹���̬a����q��r�׭l�¥e����	|���z},m�&���-�[��=o\B"�^$�����c�%�`��6�C�����\�g�U���}���ީ�����g~/��z�����ފh���?#[��[�u]D� ^{(���7'!�F��&��s�pﳧ$��r��2�j�G9P�鮛}�/k�d�e��@�}��p�tɿ�O2�!��3�w���k<�q����v&oc�o>8m�
�v��Ԇ13���L똽�BT�sAw�]0o΃+���yڸ{�׸ѫ�
���6ig?y��v���eqc�=\/n�ҟDZUbn1;cG�ä3��#���h�&-:�鬾�螃�=��y�^��,�:I�2����$T)t��u�+�#bRw��s�	M9�S~�����)ƪw�x�;w�IexP4�ZM�<�{��������j籷W��л׸�Eˉ9�hr��)���7De�;�&��SQ� �j�&%*�n�~��O}�ğ\-�V�<��=o�Gq��|j7�����il����n��V��)�P���J��'���0q�>��ܔC�y�
���=�R8��g-�E�/�g�ϙ/�@U���#��=A����)���>V�7�9�F���f����ճ}keL��]h�ΤD�K0i��2&3���U!z�P\bkՍ����u,�T�_Esz�Տ�w[���ZZ�Y�\���)I� A��<�̠OGg���m'��y)�Ϗ'f��+Q3d��7�f�N����f��N{_ݴ��w:!������'f��r�k�{f-G*�u7����[�t*]��d8��2KNŘ��/�+�]��ԥ��Rq�w���wt*;.r0�n��۞�,mK�l��	��ו �d�Y��su�:�7r��Ϸ���Y����;��纯Τ]��uR��ɠ�%<�w2-FJ' x&p�T+��>6x����b�[��;v��z�E��h�n_[UT��G*c��j�'o�y��}'�X>>%Y�/�t�ύA�}:�N��S7��x�*��\?D��Q>�\�{ɫ��s��xo�8?���O/,O��t棧�T	��R���>�����­�qʹ���6uWTfx��i5�f~}�w^Fx�*r�o�e~�<��vx��2Ǩ҅���{j�+A��av��(t�Z�=�u����f������=ޝyu�o�׸���T�CI:&x�ROq�ۺb��t!dYɞ�|P���=���St�y�-�:m�h=>�^��䢆�xP6� �x�s_e�~�<6S�C�7�����Y�A#��;�7�=��Z�=�0Lv��;��.j�����9R���_q��Ͷє���%2ܟ�A�	��;�7�sOu���a0�T��E7�+����2�
0���n$� I4޿�([ݮmI}`!len>=f��9�?V��[��n"[����CS�� ��y��	ݰ��U
@�B�9p;]���.�m���ahi�yVR}q6��q�S���NF�7deӫFmL��g]|x/b�������.d��Z������+��b����S��{I\�p��9Y՜��iG���^WA�<�yFC�&N�I�6�#�MR�g=�XW��m�.��y�c!�z�	y�����4��?���t�+�'��3��T��F�울��W!�c��]Z��Q��fWmϹ���tٛH��偮E����
�D�@2/�+k0�(�9U��S��2j��^Mk�sq�w����WF�c�_��K��Mk��s�����g'�^���vX�]��>��s���R=�4��]G>N�� :/�<+{��o>�`��%���3���^矇�@r���S�+Iù���ܾ�~�T���⹕���v��4��D��G����в���,�g3;ڱ���x�����d�WS�8,�S';e��ކ�;��
�8����q��G�����+�ꇥ@/+��|4�pPh�띣!˯��*]�wɵ=0]fDH�G�������{������f&�)ӝ���K&WR�v�$�Q�+i
�p�@���[�7����Qi�5�a��5�	�9I�$��%��{׈�]�������/P��	�9� �2P�W���kҌ�I�F��f�eMz����#އu�t���q��:n,�{� �/�;P���϶� �b�~7"jP���3�.%�C^�vE�b�nw>~�z�7ҽ|.eHۋ�$�<��[�ϰ<��fUQ�N�ޯd�e��=t��]�/it��!��:��\;T���^��d�tw7T�Ck���3����*=T�l���O�������ei�c���y���^e�5r��@�c��wX�;��l���x�t�4JxuԦz)��7-���dx�q#ט�G4JՈ���߭���X ʄzO����F@r
[$Y<�}��(u�wÇ�[V�����/��M�u��{oNS���n�~n��N�r��}�@]P'I���u�n(�/8L%7��ә�{a��=�"܋�n�c�[�%� 9�D���N�R�s5���d�����rB�w�����>�w�2벇q���4:�o�Ѷ�p.�>�
�*�tڙ�qE/~<GlY!��F���ͤ6Z��s���E��a���&��L�A�]8��m�R_(�;w��:�9V�ײ�|?nz��ݞ���e��po�Ynf�$�eėfoSw�-����f!m�XeYg�LdL(d��hm�K�v� ��n���_�e�������Wgp�vK��S�'Q���zw��6��<ɣ�	�\)�y/�%�CܽF�K���-v��R�
�:�l�+��8%�[����꺄���!k�to璠N�9��zc�}=K�ξU���������2���za�����ꗇ�Z�'se��w�ǹS�E�w�㖰�\dv�uo~g|�\[��޽C�
ňOi�K8��c�D	�0����U��m (�o^�/W�m[٣���*��>j�9X�\$s�崢�2�1���d<4~T�Ui�3d�I�c��L��N�Z �}DoS�nN;����MW�s��gNI�,�%Y9�z۬s�WF\*���>��ۋqJ��ù���]1�&�O2��BgS���kև��N�0�,��j5���$ۉ�
��u2�b��t%M�)�ׅR�ʂ=��ܶ{�;Wg��v�Gw�<�m�� ]��/�x��v�� �(\T�p����Ji)�;��5Ô=~LI�V�/[�[g#���ڮ���0��Q�t��Pq 2�N�޺�w��H}i�<�8��F�F�*0ѡ�QxM:��aM9�\�:m��N�� ۹'��{fP��E|Mp�BN�,�dlN�.Xo8>�4�Y�ԧ��������4\iO�#w7�iS��X�n��a�������o�R�QEݪ�e�#���l�+w@kB�D�SM�S4w�ge4{5�þs���v�����D�`�ZM����v�SL����}���~�wK}�+���Bu�I����N�	D�9� �@�o`!�$��UO�Wg�l��R;�3P���1���}ϴ�p���w�_��ٛS$�޺h�lE�y�T6V2��[/���sk�\EKӃ=e3b�Q�����ĳ2_�*��{�2:���;���{d��\�r	��:�*\�4/�s�j�ii��tC���_ܓ�F����`E���kI2^{V����A��G��K�$�Nǌ-�/�*We��_�o��Cn;��-�vj�L��Y�W����쑵/��;|�+_�A��܁��9�;~�Y���/y>�5�lY8�w��=u���[��Ƕ�hy���k��/�U�[>�=��{�#�(���3ps*����Z�p��s)�"M�>=�Qq�}l{�UOI�*c���bs�{E��I��p�b=���W'e݁x���sE�,t�gA��O�@�s��3��}�h�j�w�����6�a{��La<6��yE��'�`'�es�|.�'y/���ʺ�;F�kj���A����"ɧ��W��'�=ݖ<�;��5�9����ᨇwr.��v��WziT��㱎��&��x'S���7pkT.f,�H�S#0M�d�ϳ@nf΁�0��y�6{���t_�::K��*��%�@Ϸ�Q@�!]$v��&���%wy��m�'לc;�:v,�{�B�:P�_�T^�3A�av�|4�x��~�R����[�g�R}�d5_�K�ʚ�]s(��0L���!$����)F]�N�9UF�U�o����z'R�;�����c��H<*ntr�rQ�GI=_�`��]�v�xe��ɮ��=���븝7��M���>�r��:i���#.�a��|J���7��"ϝH�[KЂ�xlڼ)f:1L ��oU������u�{��)�����їv��6@��f�pfw����@�����a��|
g���q���up�D�i��*�>��
K]�����~��؟�7��y'����"?�>�H�'�Ї_eH�}�ւ����Λ��ͬw7H�7���U�I۸���fA�1蕴��]���G���\�]}��=��b���m���2_�9`k�Q`d'w�������E}+k0����k�f��5c_Ma��5�����}yc��v�zz�ƓWB�fesWL#Ol:��z�An.B�[�p��6��W[2�� �U��f�����*wv�u����5	����u�լ��:ʋx�[G�ܓ�7���C�y��%X�r�eE����d;Γ0��O�ˍ�.yl6���B�@:����ই��H9�K'��`���jϕ�wY݇˰�1�:�7s�_�zV�ʺ�������@:7.���{���Ϭk�IRS�{4e�o�g�Y˂��oᓃ��Le�u��t�6S7��Ъi�rq\�}U�`\办*��o}=9�-Wp������g��g����eP2p+���p	��O����}�cʫ��gR�C�a37���Źy�q�iy�yDӎ��O���/��8pҠFJb}������׶�b�m�����g/ s�t��S�0�|�W�ʝ7e��A�^4gjӪ㭸�(�ˎ�������s��mP����"��s���0������p�*F�\�'MI�g�o�[��2�3��׾�q�(ϸ۹����]���O2~Q�ᾟC�Lo�z�/d����"��G�3��j�I��&uG_�2������=�Jޟk�����!����o�^N�b��efIx��q���`�.O_Ҟ��]&}M�	�������{����-#�����ш����G��r^�P�ߣ�������������[X�؝k�̋�4]"���Qt��O:�ZL�d̜��INU��ᛏ�Zc3��:��*��^=Qs[���v�/�*u���.�҄-	��X���	5;`ro$ۿ���/±Z��a{��(� 7��AKd��y����P宸h�`t��� ;�����#��>�a�s��ks�M�P|];wh�F����1q<�h�QZ^f�m�סǤQ���@>��Ӯ'_�}#E��V��uĸf�'Su�N�Q.g����i"W��ģ�&<%�VzO��^x��=�*�m�3z��ۄ��m��0�^�U k�S::;���.�w��x����N
����Dv��q����Wto�Y<ɣi�_��R�nFڮ�&���������L���<7O����8.���Vm>69^Xx]�|'�2�u�o�9��{~���/�O=��7��|Y(ao�kaة�NŅn���oS��=�~{�ǖ.�RG��}�=ꚝp�Nu�i��z�
�
ňOi��ɘ�ͩ�9��z��*pv7wo���"=�Ϸ��w���= _���L��\}ʟ9Y�\$p|��X�ʘ��݂�?*�ӫmQ�|�׺���V쭯e5�����%�7�s�"��srq�F��Bj�w���S�z�~%F��e���n�`�̓��Eg�H�=�H��T'G41v{_�[�Z�u-�y�b������� �$v2.;"�y���lCմ�v@o�E���X�s��Y;�U�tO�>��X�j���nD�!z���af�7��1��5�M7�y|�ı޲`o!Bn�=�.�k���vk���2���v5Վ�_$hx��[�6��'��gL0��"oxS�G:Ҭ��M�e�oou�7����e�y�]�T���Vj��`��J?d��E.��ru)U\I���K9Tr��]�U�5Y�koUf<�,�c
��Jպt�T�f[�R� K�1Ӫ��n��aӷ�P��J�r���{/#\��H�J�{u}㎳β%d|V��9g6�{�n��f�5�]tw�. ��-�m�fn�OT�8�sf�w�KY�/JIΧh����'
gZC8�b0�AaWJ��HN��y�ͤn��ۍ���� �]����Q4����Z)]�J�p��m7g�wƃ�*5%XӺ�}h56�����c:ĒKI�*�Ǫ���onp tՁ6	��W@{�t��g��jY�e�X�{F�b����\mm��x�,�s��f��.	ݫz�_62�e�ٴun�w�sԗC�����
�}��i�*�ZbfU�5��ZpT��*r����ݩ��NN	7�t��۽ϊ���j��0�9M�u�˫�	�-����E�m.����Y�`����\*\�=����ȃ�Nk'���8EuY�>4��v��͔�ŋ'f�7��"���t����-�O���6f��h�7:'dbjJ�E���k4-z�N6/��m��\�mj�P�)�CY[�f�v�@�sMD�T" ��s-�7��䄶S4�]whk; ��h��z�8�tY&b.��[O9K);��7cYY�+�Q��'-K��`���r"��c@(��D❊�ґ���N[k1�R�-�`�����F�ޗZU��nn�x�j��Ȟ��}e�<��� ��\��0ѽ=5f�m�Y�K9B����VF�(,и�v*tS��"�r�#�Z"��3W\�ҥj��Y�m�ݭ�,P`�u�	��(u;e�4�T���Gċ�#�j:� ͷsw5�:\�P�(�N�v0D���;W�����о�R��ө��+i�,�j#q�|3y}�d`qquu��٬����!;}J�i��@��eⳐ��e���oFuA٣��5o.3�p�d�Tq6��� #���7{S�Z��U��~X�4
'��xV��j�i�l0F>���.�4�ut^<�!`��c��i���w#m0vQ��G�S������]@�뵌�7p�ϷJ��O^�\il͒f�G�N�]w�d'b̽/p�ghWe�+Q������l]�G/�2�̴s��In���֫B
�!-�9ܳ&.�.IY*��#Up�U���`�l��w�*�۩l�2����V*k:�K��=��ؘ�iһ&��9�U.\���P�
УD@Q��"��\�� �"�,��습���O�x��DU��jQ�DF��p�BrQ\��ª�j�a2�*"�(��TZ)�]%�RD� �Y�TA&��6�A�Ȏx���Z���.Y���9��Ts��.juk9EvQ��&�:��-D˕\죤������.r�\��<���N3�Ep��"�DDʍ�"̨�\*�՗<w."������r(���eETFK.UG ��8F�Ep�9�$!D�Es�QEW�TUQr�9xȪ�(�T�T.D�+�U��"�Ȉ�"��EG(�TDQEATQ� �$�B�E*G#�\��L�l
� ��І���q�9B�"����H��L���nV	�u����Z����AA��=�XWԨ�f
����f[N�v���?������ꙸۗ#�ˀ�:d�)�^�?\&{��7|�yn�Mr��T�8�o%ߵo��4Z�J��BgC����JD��27�
�Ǖ{�n[<����ӓnv�Y:��r螃�-8���7�F��H;_@L��T�p�ۺt�м��^'lh��,��Q#���#}�=��3�y�P����M��zJ5�'�@X=Ċ��.�����@l���|1����W#	��x<�SG�5�÷�\���?If�z�3
�R�%�>7��z�>>�ᜏvzo:-��v�q��7��Ė��q^��q:Ѥߛ�2��p�J� ��w
�νq�h����:�7 ��q�|o����#�.}������ɻ�/�ul�l��z/ӑ�Y<���I�#I���\T�83�e3x��m��tm9|K!�d�տ#��ډ���ƿw��2i�+�s��pfa���:�	g�k#����tC���1��'>����/����gs�������;_�����d��z�d��"~�(K[{N~��^?+|N'!˧��Q�����Z��({/�]H��G;�N��֪=�:����J�ŀe ��Ӭ������F�P����+:��+�c�~�Ab��zhd�[����3N �l��iQ�)t{צs�}C��t��f����V]r��R����T�ήמ�:z�'�=�w��D���ݵT��R�9`N�?E
��k%��=1�0�m:�3S�n+4�<<M����E̦;eV�G���cE�_��}ʩ�Z�3JU�[)��빑}������7��On.���gmd�a�:U�٩xNv�f�r���B�����T�59]D���h�s�>��u��O�����P�ՠ����x�8W���<��gҠW����S\�'!��<��ݶ �1���n};����.��M�g��'\L��3��*]T��<P�U����P/��kk2'3ݛ7�8�3�>���e���;�b�3��MOp(\�S/����"��i�m�מ���X�3���vm�����7-�P�=���5�,�x��C�猪qu2����&fpUf�b����~�Q���_�����[����}��Z� ��W��F��OQ�P���x�����b��Y���Fw��븖n�ۉ�J�s����O�I���~����W�;8ݻ8op�݌s."O#r�@l�j���>���N����g��'#ߛ�3_:s�"hp�����5_��J�rk��[�׋���7��9�ɼ�-��E"�z�;�3��	GD�(��CV9����퍵u�L��z��3���9l���YNf��@a�{�e>f���\�z�jU�'�]2��s�D�>Y��a�6O�m܎^�*�2h�S7�n�����L��)�|
g��eq���ý��c�}�������[�
��H��f�/�K�W.����GT����'�M�:�{����]r6��йӏR�J��,�;�VY�%C���TW���L��;����+�i�����B���is��!q���ݩڪT�~X�ǀ����WJ'j �_�
c�e��F��g}3��.�	k���ʸ�\-7�r�a�5G�:����4�4=z�rGK'�a�(�<�!����Ưq���F�R��q�+J����7�~�^�N�� :)�������\/k���[O���Y[W���L���Q��c�Nq^�2��i:sJen_\5&^��u�"�m�Z���
�����ؙQ:�?^33�g����N\L���Nu>����W�s��H��=׭��[b�ZNFg�-�ʚ�82�4�sC3au�~�S��,��2TOȸ�3�A�QC^���%���~DV���V���-yv�s�!�6y���;�p��Ν��'���z�sWJk�j�v��is���o�&244�O��Ȱ�_�s��K�%f	�rGK��O�����̾�wr���3��K��o�n���"��̻׮�
R�!�XZI�L驻� m��ro��2��,p$n:+���(]`�ۙ7'�''Q�ɦ�҅f�y �����v�u{'����^��A���#��S���އw����+���!vT���$�M�����G2����{u�.�G�(γ�\	Gc�������9��c�o�Җ1M֎��F-���n.���k�,ϸ��l�$�. 5#쩖�_]T��8ҷ�ѮC+O��Gs��͝�e*���{&�WO����v8�pv���>���(	�<����]&}�p��n�`ż��ɵ��k==�m�L��"�Hþn���R1�d�_t7�� 8	l������8�H/��T�~q����A�BÉ�VǾ/�lnBu�O��>2��Ox����N���W���t�^Y�U���O�y[�z�i��}�.95hzuĿ>�M� ];�D���2(^Tz:o��2�4��tk���Q�9[�	�H�j]N�6�~��\)�3�T����}��PG�D�ywk뙰�̽7�����WR��7����ˇ�����̚6��5�ǐ]
������E.��k���L�c�NJp�;��8.)e1W쥦���	'U�0����S|�`_X���$<��o4�`��p�����-/9���n��I�<�p@��a�[�/�II���7]��S�'����ӿm��Be,�vA���O7�����������3�	�yan\zh%��Ըb�H�NN�3C��U����-*�m�Yŭ�����B�l���k���E��?;�7��ύ�id�@���X�KÂ�V������95R����_���~:��=]s��	ŕ�C;ީ�iD�߁��;�=���ߕ]�G�"����
�ݵH�4
ko��}lzS��ʟ9YU���}���=�뎖Ne����͊� f|����>�Nﮜy�J��5-ށ����GK�jK�u�}��p�S���������.[+�
���ӏ�ф���ʨw���ܸ��\1�&��/s���y�\n���5��L��e�h��[�-�x�$��$�L�� L�WS/�/mP�7��^H)���h�zoo��_��|wյ���;�Qؽ��@H/��OW�n�ҟ/*�^����f��}�ᛙ���ՄgC�3�c���&��6�>��#���2��{��r�M�~q}O��ӻdd��;ӥD��1 ���c�SG����s���N�����j!z�3
���B��3G4S�7�ґ.	�;�3P��b}q%��z��N�i7�茿�ݡ(��s�����\�d�l^Q�0ЃkZ��@�F�"��<{s���OV�*�.�����t*���b��l�+��:x���Z=5��;4	;o�æ��U�2CIJ���Ԙ<�����9Į��/p�c}��p�fmܺ���5gǀ��;�w{� �� �\�^�ơq��c7�N�!���E�`7	��=6!�V�]�B7�հy�E��/&I�_:��7d���]JӃ=�S7�.5|��N_�U�D����^h�[���}���'��`=�D���g�s���S�Ж{Ʋ;ii��tC��L��۝S��s���:��?f�4m�p5�*�F�FI�d�FH}b'� ������5p�n��	�+U��Y�}1�C�n]�h�N���A��r�����(Tk�H5�K'j�;`������Y��\�W��Y_�����������/�ǣ�S��f���VO,����(�y �tE3�������x=�L'^���Ԭ'����_[UT��G*c��������{Eܻ�|�-��vs3}��}'�ޔ���P\�W^��d�'��J�Q�j���S\�'!��=�y�P��7wk{�WDʌ�׈૙�̛7ԗ���Z:|��pJ/�~�^��U��^���Z�� �ӷ����m,�yGA�n�=��V;�?�Y5mO�ĥ`��Z|#K�~C�ՙ��e��{t�;�[�e�;	}}������wU��/vK�E�c��;s�Ӭ"�5�OuK��ފ���!�/��`�K����H�ӡ �k�Q��i�x7o�R;���O���!1�bä�듭Ψ��tO�n�{g��G)�O;�޾�;yނ�.q�m�/:c<�6{���)�q��ީF��'A�Ϡ�R���Ķy��7���:�V�y��/in�{Kg=��	�O�z�/��B:I���|}�#=�gw|��qp��G�������J7��Mĥo����}�:i���#�a��n�/����wl���|�@����;�溰��)>���N���*q�ҙ9�OV�9��y�����6��[W�n:d= i쉐%:�L�����7�b��ޔ�#2���8��g;����q�S�gp�m��wlȸS%�F��Ϧ�����c���y����cT�zo�;�[�w�\	mYs�J�u�P������'�L���N��[.����zڕ��o�S>�ٮ����)���׭\�/���JY-@r���	�����N���X}����'�j�vP��>Ƈ{�yÈ��p�裨�_����yl6���,t�N�_�����T�d��&e��{�wj$ۀP|n ��+���qr��;�a�U�v���k���]!Z�yD�y�wV)ߏ{R��"��E.�����c����N�GM%�U�te��Q}aZ����yTǍ�P5e�Q�����}��&�/g�hla4w]amf��9�B������ue��!W�]��Z�o�m�5�'8�ʈ���7�a�Kd���0g�o�>�:0�Srǻ����4�sյ�*�za�j[K�������^��a��=Wq;o�曈g�ύ�g'/�?P�����pY����i Q������F������������U�{���j��s:tY;��!�D����+d��
�T�)�ͅg9���ZG��\u>~`�|�=�����Xյ<n�ĥ~C��mۤ�s��rUtv�9��n-�*�7���/an��y���L>����W���ʑ�����nٵ1=ݜ_c�M�&���v�n��;E@�w�J��4�x}�C+1�7���cM.�]�.����xw�~q �;P�A'j&x}0��L�1{uS�⻪Ĵ���rZ_O������V��,���4��W}�u�_��(҂�@G�iO���Su�k�:�D,
f���u��3��f݄=�U�\k��n#���wv�(�Q�� oW�@r
[$\ϧΖ�*$�X�P9��Wt��ٶ�D��G��m�ϓ��n<���t��M�%�"�:Lz>��4����2��=�{N`{d"�!95rr��Kɳ��66�V|�`?2�㬝�3�2���Ô��(��j�+tR�6��׆��l��R�9�noTӗd�b�:���{q*�����m����zr�D��xҘ*���	/-=�۴�go����-Q�E#��j��ޑ��T���q/�ς%7>e��M��3ꢷr9}R-��7��k�t�kд���"~��Tn(��ˎf�$j5.�G�m��0�^ �w\�MTι�{��@]�x�6�X�3�n ��T��%3�9����ˇ��L�вy�G3��-&��E�z��S}��`n8�zԿL�0�N|}(m��G�Jӱ~�����|lr���瓵\X���WB�����8���U��,D�yf�4�������2�+�xp_Z�'Wx����u�o�-���~y�{�Z�k��hNZ��b�ީ�<3,�r�>�
�{���e��̞���2���5��s�m�*3˭�B�w���T��jhn���\/���G����Q��s~v\:�Q�G.�q4\�>��$�'zR v.�7��7'!�F��}	����\}��Y�y�.#��,3�{��v��۪���)�q��(C�K��wܥ3�
�:��v�Qj��_>螃j}��9b:'�Q'Z\?0��O�_�T��azo�SC�)@�ם3��|k�9p�4{$o�/NvSfP�7Ws�ːR�`�zeӶ��v��_���<f���V��{���۳׳�*A�WQ
7{(m��̴pq�vwEOTV�(�ěE�W��.��;��d�V�r)�䫝TN+���썕f�L�snɮ�c
O�=%SH6��������{�d�����*�;�Q�� �D@O�℞�wN���/Y�%i��5%��5��D�B��[=�!��t�M\=�U�a�zJ4��z��b�$?cC����(��ܗ��%�w��v�h�q);���4{#];q�\N�����j7��k��U�dC�b�=������^$үx�>7����:}�����s��F�~n�ˊwhN5p=�0zjO�\>y)n>*_�@��$�V�`�/�&�ƣo���#il���3J��r9��^9�����нޫ��8�ڶf��(WT��6vH�N�U�JӃ=e3x��m�˭�9����1A����K����p�Q�zO�vSH�_uʝ�Ls�����h]9�5q���i#��uME���{�g���<��Ziْ�p1�U��eْk�(��k�^�9][肰L^E��I^^�@�ʿ�[��ZF�Fe1���1�;���Sp��'y�H�s �d�v��;W@�M�[�9�ٸo�ጞ��Tw
��C������T��!k��[ʰ�gОՋ붅��~���҂�ƛ�ww�^�-��L/0�U���lAK��*GRo4͛{�P��
uÅ�)T7Ըg&hR!�t�2J72������AO��"Q��c���N����1�tl�u���2p�x"��;�ʍ�7�Mܣ�l��xT�^�V�K��w�P��J�$< ��thhk+e�9�������J(釧�Y{v�Gu�qC�ZG
̦N�g%|�8�)�ᛮ�j�ɲ3I�[�KD��F^��%�9�32����c!-��+�guDѼ����{VtXň�Yr��A������[>u;�b�-�yi��V=1Ս���h4�3�[T�𓣊)7(���]I�K�7��P�����	ז+[���mnQ�Y[���EJ�Z�c�w��)][Qbc��M){Ox����b�/K�*��E�� ��۳{�etʲWp��n��LE��F��=V]#�9��� ����T����r�T��q�=o��[w���3b�Iݲ2#[��z�0��.���\���r��՗c��U�q�j��v�z([�N��uB��v9:��s-^po��2>���;��̝�.�h:�jp��N��S�ͼ��Eգ
T�[J�тZRX
�I�k��|���ۏ��t��X&��Vh��Z��_U�
�(s�{1`ʟ]�c�}�ʴ���hF�Ǽ�{���7N��oY5w�N���G[m����i����(!� ��T��x�x1Z%�a���]�zfl#@��ϝq��ɘt�^��^��x��t[A��S*3�\��<!5�8l�E�
�����e��N��9}X��wY6�};��f���u)�8�rdaigJnj�F[�&�mC���{�2��b����ܭ�]+`�.K�	����9� qi��ieNi˼ر��2�\�d':��qo��b��� ���3@uH�<�՞�9SU^���o/$��C��C�j��h��*5��'5�3eP��՚�Е�W0��"���gb�hv��M��3%�e��� v��<�Stҥ�w>�+tٰCZ[��K�b���w�j>3aɕv)uf�s�3Ș�M�7\�طx��Ȱ5W��V��x��':p�<i�_#]f�}aHʛ��J�7}Z��@�"ٕ���	��kDv��
�e�JQ�r�\�rs��+��ʋ���8C��=!ӛ�wN��J���W[����7O7�OA}�!�a��vK�vgVյ)��44% �tC�V ���zeW-U�=����%[�Դ���vHWR���r��bL��o���[�k)D��|V��Ŗ!Ma��6g�m���,[{K>��ն�������ltvܩ>�[�K���.��1��4�T�k�䯔N��d��_Be�ǇkE���=�"�����>ޮ��,��F��,�ф5��r�h�=̰���y��w'}�P 
9Q (9p����&E�R,����
����)�G"�(���Ur�G"9�+�.DW
��E��o��ANQ�H��*(�*����Q�Ad�p*��j�U.UW*�Tr"+�QW"*�gd\"*e®4�AE��P��*9\�9H����dr�����r쫔E�UEQr*�
�+�QF�TUG9\���a��\���9G(��*9UȢ��(��\�nA
�(��8E�.Aˑ3�T\��D�"�UQE��EE�p�PQr����k�UAG.UQ�(*("�99@���rr�*��WL+���"����TPDTs�E$\B�
�ud��b��W�XH��]"Z���+�B=�r=����L������n�n�o,��{y��}��4���6;���!���?٘?���^�.��_%x���L�n_[
f^���js殢w�*Ϧ�u��O�u�O<F�ۈS���=�%�u�6jy���������Ms,�57�ˍƮ}Kݶ5��w\w{���~��̟d��tw�]iP}>��8G+��)�����+[4�Y;ǁ;���_\n�������qY=��=Q Δ.�_�>>��o��,p��1ǣ�O��P��t��C����1��R���N��f".J��
�{���6�:��wu�yz�-ׇ}�%��� �ӷq��)C�%�u�M���s�����դ�pf:�uF�-�߻�q,�%�R���5;��@->}$yP�N���׶'ܪm����C�����!)�q ��4��뉿�;�>���'�ц�g�i�_�X�$1�_�YqJ��S �]i��d!*�nL�����b���������>����ϝه��|�;��Bn���;�d_�d��H]�6��<�h\R�gS�����^&����M$Ӣ��x+&�>+�ѽ�!�h�5��Zp)��Br��T>^�~!�㕞��x= �wŻ�GqF�.��C �%e��`?R�tkxX��%	v�ȋ�\Sk3��ʽ�3�Y.�w��� �}ә����)c�����l1�����y4�]&����R����P[�,���%z��
N��Z2����]bw�:��[��v�W��}���wVxKT]욿��q�\�.�	)d�e��q�+���T}҉�������o~v����?e
��Nz���X����c��WF�X�V��4�4=P8�ǲ�3
����5�zo����/'��Ӈ'å�x�����oJ�n_�'U�����u�;q������H݃/�s����E�Ϯ6X<j�����_��c:�i8v#6S7��]r�Κ�����/�4�?�5Er+]����y�ٿf}��œ�㡋�V�_?�8�����n�-��r����デU��1�j=�:��j��s8PE��~2��;�!�jp��r���֑; {��`W��|�|킝�g��n�Cy\/;*tݖOvz{e��./����b��×v8^.�F�̳�n�K�6�0�[�/�S���?S�W3�z�tsy4�ut#���M�]�:�U$�rw�D�te��@�o���.�F9��c�o��{��"�_�>d�Ď����5�b�����L)��#�&��FmMq^c�s�nd�haΨC��J�z�$����"Y�u�z/ڛ�a1�<��%m	���5�y�R�2�o(U��<�zT�Of�I��{XVq����5�����7�2�υ���z�}�p�䭕��N6�z;�d���$�(���L�1�3<r����Jޙ޲�ƥ����fv�b��ߺe�8��!�>�[2��E@{�&O@����;�I�1P������inR�C�?u���ǭ|�;\u��n�㪤ah��k�����}�D=��_����6��X�^m�}Աl����뇮�p-�A|_��܄�t�7P|v"����FJ<�/�R�7�\7�1Q0��z���+=ơ�]r0r}\n���D���9v���������g��{g�uu��#t�$?���O�>ݸ�o�H�j]N�|ۮÖ ��Dؠc�$����c�����<�3R�(��2�+{^����^�+y���Cj���Y���{1O�%�Eǳh~�z�_�MGL#�G҆�s��b�c���������5;�F2o!��;�+��q�1u��C����%@�N�G>��g���z��X��������"V�ˢ��I��vzwZ%5�¿m߃���-t9Ͼ{4'.^��O��'0�[ώ�}\/�Ƀ~�s��M�ι/�+���sٛ~wV�N@@X��'�^� ѩ�#̭W���G��H�ł��r"���-�Yoa d&B���)]�_v�u�{B#'k.�X���gu0Q�3hW]{�rC�t�>x�U��m"Vm��]g���{�Ov9�R�f�:�s�v� Tg�[�U;�}ʟ9X�X�>��\2�d_��ƺ�i�Vy${_�e�C��Ua�5)�ށ�������\ܜ��F��|������h�,��F�u�Ro�6����$�(�%��;Q������_х�&��/oh-����3)�h�q߆�X����q~�;'�邏���^��_L\m����4:-��Q99n5g�+�۰_��=������Ц��=�Q�� �A��EOW
�c^�^��0�z�4���gKUӷ�B��ݱ��k�Hg�v�5p���U�a���H�'���щ�����;�x�x����!�T�l�!��%�}I{D�������Cߝp8n�p��g
�g{`�7w�8�݌@�fc�O�r��%���0��b}q7�{�����r�MǛ�2�ay%�\�.���}�tߟ	l�٨d �@�U��Z]������N�>���[;>�b�a���w٘垣kAy���'�ٛ�L��}RWM��"e:�W�JӃ=e3���,4H��#�g��5�P�:.����T{�nYT�lYhM6�*�6���L�V-5���q�0$3]�_-�|��X���Qݡ�6R��4��$6 �6�q���L-H���U��7�h�;X���)�
Q�A�sD�Z�k��D��V�LO�p{�q���%\���W��4��\�ٳ3�uxTJ�f�Ӟ�^����Y�T�s�9IN�ǟq�l������vd�7.�Q����<9��lK���.`�u󹝎���3σ��/_���Ua����X�:�NX��$g��Rd�v�����Z���s�=�%��)�a��z_g��Ƌ�r�lr�zV9�yVl��B{���D�}\�K�]�;��=�G8��r��l��2�ϥ��5+	��S+r���ʪ���T�53y��R�,�˶��{be����!j��}q��×�%�q^��$�'���P+������w����S%tg��mvT��:NQ�:�Tn�w�n0ߦps'��(z�Ύ��G��A��U	\* �^X��TJ�1�������G|��7|��1y�S��{���t��z.{�j.�z���MN*�KV\u�*4�k������|�6{��=Fo�-��TY�N�w�"����d����^$�\,.�x\EL�7wLR����!{Kw���[9�@Y�	�O�z�*�w�O\J�+މ�*�߻����C7��\v����|�fM�h4��j�o`NjnTP|���PyR�9�D|Q����
X_����I�<�P׆��)�z�$�Gӓ��5KR�D�㏩�{K��3ݥ�(��X@��Ź|�!��F�7��l��3;�������l�(��f�0��H���q,�Ԗ�Mĥo��jw���A��Ip*6���n�n�sQ;��C����Q
@�_I@HJ�T�w\�\{�O�&�Ӿ�i[�
��[�^�b��2�ϑz�a�7Dz\�2��2
= i��J��S<=�����K�+=j��^"�q���f<��i��p��7pr�ݳ"��G��� mG>�L-��.ļ����]�͛�q�~U#6#�[��!��y�Q�	۸���&at�اk`Z���y�;ۊ�Ô�h��yd��m0�R�_��]д�2_���q�);��ߎ�J�����A����D�C�g=Q_N�fQH�_��i��yly�WF�X�W��4�6��x+Z�M���oE�����4�� �=#��N��e������7�~�\�V�&��D�=>��G�f��`mڜ���>/&}{,5����'��S�+Iñ���4�`vq=�{��5x��ǟ�SKLy�̬�}w���y���|�ᰏ�go�?G�6v���������~F�]/gmuu���u�5�7���sN�C�9%��{�<�D�"���el��T�&����[3��+�M�8ͦΪ�Cφ�K��t��p�.C�i�`��c��J�D�`�ب���u+d�4T�4&�dq�.�c[��5;|ov�gf�WƉN�Qx��ǝR�c��{���s*t�E��~2rމ�_���ꥐ��ǘr)�D��=(�r�_�O��9�l������^vT阥�ˇ����W�����D�83�L?EuW��t^��A��-��78���Ϋ����ǍeNkn��>"߇��F��$騒ѯ��T+��/��ʁ(�%wѥ�Ì�W�X�x�z/9>�?��=��K�/��:��P(���A'I@X}P���3n�x�WuX���FB ���~�a,ø���/:C+O��GoϮ�6���(�( oTA������	�O~㞟d�^.�i���n�`�r�k�F�v����UH����@x�a�exG�s��\r+;O�ϥI {2m�̡�]p��Kj�����:�&���7N�����F{�i3�is��w�X��'����ZVz8�%x��4_&�D�p̈́N����[����+�粒��WA�̋�8��-�����t}EiʽێgR3��[�i��\��>��cٮ���o�,qZ�O���M���w�i]���q�I���>��Ny�kƠ^G5P'�\|d���k=�s�rk�q��)���J7]x�ڻ��v�Fҩ��3�ե�orm��ĵ�Dm�H�PkV�.�c�=��v4�kx)
&�����.���7n����Z2�^�a�a�k��^�q�]���sˇ�����.�y\͞}~���jжg]Q~��&��n��耪��6_�Mt�=4}(m�>�{���m{�{ejɁ�9j�v�ź���߮5�U�8�E��v��7���K'��G��=^q�T<�~�͞�{ӝ������D�ͮ��~{�=�z!k��|�hNZ��`T'���d�H&�k�0{�q&�s�[0�Ҵ�ƺ��v� W���ǡU;�}��U���}���_|)��3�'f�m�س{\�~�N`0�����Ϧp�L���) ;Q�S�nK��{"�{A]]�N��w/���Q��o����[�d���%F��灞����;��,G���p�L�|A�]���6���s�f�eK�;�u�[����Y�.3�$��$�}3��:��cv�	S|/^u�T�� ��h��x��_�;H�*�Cr��C�p�Ц����F��t�nʊ�k��ci���xs��:}���\bvƏk�Hg��Go����|Uy�~��(�����)<F���᜽����Њ����s���-�s��.��j@��g��[s�Ha�w&[���FlV�D�'��3��V��&56��h5������B̽�����щ�YUr��";u�4��G��^��sɖ͹B����1��U��[E˙���-2���7!���ik�oWf~�~��ڧ�޺�W��H��'x=�)�ٮ���~N���o���3,o�ћ�=��QiT��%��@�z�8�.7���ۧ���+)�����W�tl�w���n����n�M���� ] �ҭ�A|~��h�֍�����7�?|�^��u��{gK�9���`7��.%ճ7�)�P��+���9�^���{L�i,��ɥ�EŌ>��-�fw����{v���Y_>d�^�M"GQS��f9�M�J�f���	�.ś�V6kc�;�$i�V�\�������&ۗ\)���vd���酾��5��M�f�9��]�Q�)���+Ʒ�HouU�5'wB�:��9`N󸑮�A,#�^�����*}��l)��s+���u���7���~�9L�=��f��XU���}P�k��:��z��#�哔�"3&ܽ<jV���sմÅUOI���x{Zyy���［�Qt;�/Tt�?\ѵ����8pz��`������5<���9*���NN��Ks1��f��V�w������F��|Q�\�$;�z�����D��=�y�;�*�(^��5}k/:��͚��轍��p2��8��pS���"�8�L�����5�M+_"X�y�1�9���{%���7�b�(�y Ȣh6� �.�W�T�y�Mh�s�s��j�w]{J���J���ȗ���Z:S_��=��Ԕ1]@U��³��l�;:��oV���t���c�׬�����?��q���ۇ�]��ss��<L�w�^�l�kх�\b�Lbr����D)�q��2�LD�Q��������|̋F��J.�Z7�t�<yp?}{�%���@-�����s����k��;�M/8'KI@�_T+������%�Kj$�O���CS��@�o:.Ϛ�;�������#.�a��)��I@HJ�T�v�Յ�S�R95&�y���xy�nc�:��ϑ�8܌;qn�ˊuh��)�Q�Og� 9	V�`�x{����zK݊]8�K�m1��[��3{I\�i����ّjd�J��C�ĊW���������4��۟*sAҕ�<̠�\�������ʂ�ȕ����QX������V#�<�<�8�Ov|��9��ߨ��K�>Ԯaņ�)%L�����B�?xx���{��<����cmc�m��0���C�m���1���co���cm�a��6��1��cmc�m�`�co�1���co����`1���1��n0���0����(+$�k4�L��'�0
 ��d��H��z*��HG֣f*��;5UE	�R	UK�$H*���$�bH��IN����[b���*�F$*�gvl��n�������vۺ��M�,��1����۳]�s��kM���wn��s�]�ۦ��{��hө�����tZ��v]w7Z۬��j����k�یXY��c���}�]�T˦�ۻr.Z�YF�'n��u���v-���ݻ�m�ef�Ѭ�n�UݧWvww]�sK:�ۮ���v;n���m��b���m.�vNڻs��۲n�f��K��v��]yڮ��\��  �ǧѴ��ޯ:뮀�-os]���]�z(����oU�kU�=޽u� l�뻗m������w��q��ox�5z�Zv��ݷn�]�]�kn�Y���۪��k_  �>��C�C�ֳ�ۺ3�h�ݠ�ƀ�����  ��|��>�(���G�F:4� ����q�    ���x�4h��tQ@g�ϼt} h�o��44�m_T�v�ƽ���\��  ��5�\ͻV����\vե��������0uͻ���j��U��֜4=k�;�q�)�u�n��G������v�iu�nʮ]ͳ�ٺUw�  {�[��u};�J�[v� ��m��Vj�����z�{j���C�K/m��R��νízWlz�8�T׭������GKvf/v��ݜ��vݫ���uu+��  �j_O��.����k�5�y�tt���uN]{֛��wn�X�㠶�V�S��[[J�{���]+Ҷ��^��C��)ݭ���F�{z׭k����f]]�o|   _{�}�U�n�{Թ�[`zP�w44��u{q�OZ�-����ݺ��G{̧�zu�{��<����i��uiF��TZ�w�֏C����އ��v΄=�&���ۮ�m�-�
�;wv��  ��j���kt���w��P�=��ޝ�Rץu��w{�p=�c���r��t:���қ��<w�xh=;��V���{����+����鮻�^�뜮�vYի;Asum;m�r�  ����^���z��`ˮ��]��Wu�.����)v��y�z���hk��xt�/p*�A��]�] n�.���z��F�:�N������[o{���s4�3��ۻ&��  ���h飷wk���Ge޼��]�V^m� �]�uն�ҏwZqХu�i�m۶�ѭ;���pӭ���m
9V�]�{ǎ�퀪/w�k��ZΧgN�wnّ�6����  �O|4P�g��{v�;���^4J��95�V^����ku�\��W����y{m�hDz��v�6W+s��;��g��վ 5O�Lʤ��!����S�0���=F  5Oi��T�� ɑ�S�A)U4��E=��e*���  M%OCJj!�)������@�s���f~89ŗ3N:�O��M/����[�����k�hB����B�$! ����IO�$ I?�	!H�B!!����ſ������5S��m�f�[@^�R�oP���%��2�ovKR�"����e\/~���v�\����dQ�+8��t����4�ސ����1
��;f 
B�LM3F� u�;&;!v�Z� b)�2n+�pZs\b*�^;��4������l�Cy@�[v+Ef�FZa �	�z3<�Y��+z��V�u���<D�rLV.�[^�7v��X�D#k(��ҁ�a�1@�����k�TwZj�`�#(E��e+.�u���H����TR�T�5p4Y;>�T��.� dzv�/mi9/i[t�Z�$�t�մ�6n�B �����`'J�n�y����HS�0wy�W��ӗx�%�ɚ�z�5���[�n����ʹv����J!��S崱U�W�L��
�mi��y�)V���cp�Ң��B^e��I�%�#ݹ�q���"ڛ��j�3jF��$��m���eIFV]�m��z�YF���P�(\�oa�M�&�VE/+v����J7X��wRVż��x�+@[%`�v^I�g֒қ�p�ضL�����%��C�se-q`�i�Q��lk=XK?J9xS�����A�3j	RJ���,�Xi%^S����A��쐗�Mh���0sg��"��:.�R
�Ғ&LO+p���]�z�]�J�Yʁ��B���uS ������oE�]5c#����N��(�� '�.���Q_ K8�z0fˤ�kS��7(�n�S�3IO䝠�
�����4��6�n�i�s浡���QAЄ�%��$�.�*��)������ t��'����-G�����3167�4Ռ��Zѓ��1�a8�f�)Q��ۧS^=J'F�l��C���+X(�j2���teH�gZ���JV!,��)Y$�v��:i^i-�hC�t����SN��c,8S���j�YZ����mh@n����n�t��nřt�`2��B	g��2ŐB�^�$)�h�h!q+p��5"�3l0�sX �*@����2���n�6 ���ڂ��H�v�l�e`�%�u��pKٴU����x.lX�T5�חyIE����6.Tu� ��jRҷ-7n֍.���\��2�۫��*2P QD],����݂�T+T��Q�x*R�(���5�[�̛��Z7D�1�:U�b�0m�CB�X�kn�֘5ʵ�̚��kیV��鰒;2J�8[�̴�2�׳�4+�X�
D�N^%ߤ��F::m����Xu��(��f��j��*C�h�����<xNaYh�jQ5��x�# @�ʬ�bB�3v���-�p��ܫfXa��쿮Jx6�H;*�VV��ea"&%�m�D
 �9.H���|W*�-e�Ҷ�tͫ��6�R/{|��Ao,��U�:�	^��m�`	�0
�v$���I��EE%��l�;VL��6V%v-	�����1Dh���I����D��lF��Wk)�QJb8c�w/qBuKr̗q�ٗ� j]Az���� ��XjCel7��V0]f`��Gom�u���ЗxHkcMD�Wzb�L�pI08um��[ {�o-+P�z*2X��!�����
 �W��4cB�z/r�ɛ��߆��x�܂D�Qh��=���F�n�x��۬Z.���m����n�M��҃35��DY�Ӥ�YE4��/M�NZ$�v�ѹ*��9f��g����2��`�̵)��/8����w!�����)��К,Ҭ/��WV��v��ht�lZ���72P�L���"�˼�&qT(��n���(2���9Z3m���㫋��z����	�Id
�O B�ʻ�H� �1���b��ې,8�a�&3Wc@e%I��b����~n�Ţ�̬��8�E��>tkkZ���Ej������J̷wFkXV.�
:�{g2��Օx���(m0Ɇ��^'���g;Z�(��y�ʺ�(68����Ex+4^��ʣ%+e+�>���n�&&qT�ح�i�y��âҠ=ĉD�ۻ��[�ouE{����^K��D�`"��2�F躺x(@��v�f�W�"�e<y`���`Q��"������)�B+��|
��t$9d\պ3m��ι�Vܩ��Ca���E=ut�-� $��[Vr��hXN8�����ƍKN��W��Eј�ǚ]�n�#�-L��t�M�:[AXʔ�86Y��~��D.�qM!#�hބ�ْ7d������r�+���	�15��*�N����ДVj�U2Z+S�V;q:�و!��B]d���ud,ư&p��t�wYp�Ne�Ej��#�0X�V]'ͷXu��l�Z�!r�J�YS+��TX�;�t��Bx�8�$լZsB��^�#�e7��{"��1՛����jZ%^Y��9�[|䂻X|��]R�(�e�2h5�����nRa�YH�4ۡ�i��*�d���ˠr��m8q<P% ��iC0{S5�n3#��Y�bT�2�l,�5Z.r��wu,f��v�)�z��FΛ��i����XP���(�n����R\�4� �*;�7Lv[�Q2�VB-\���R����mY#���(-ۨov�$���J�܌ԥ�k'j���Ed��.�Hn��&ê�b$�^�Ŧ�7�aı�U����K�.���o���2�%�:i�˥��6�֙I3a���+hU�N#fhF�]�������L�X-�h�6.ҥu��a���J��F�\�#���K�Q�ѱPB¥�
9N��XJ�#U�B3+�N�kp!w��aAĨ��CsU���ƻ�*��VJ���lmJ3p���R��̦����f������v��h:��L@��)�\-��q�;��]�#w[@��)ܤ�͐�f,k2��j7�/&���CVE;�cebӗ[%��j��U{����yP�e�լ4�`̖��LM�%i�j�pU���l��7v���J��l`�g^�I�J0�-��4��n�\��c`��]�@��髓
�Y�q�2ц�eF.�G���V�e�k+�3hJ�&R�"�WP!o"qfҐ�V�>%i� ʃi
TؑHkUt��G+t�j��W�m���f���n��`��*� �+���u�{��y��zcsfwjU�M;�@Z�R�S9��Uz~�l%K�Aln�� �7\�F�-�X���r{J�o�V�`��-�t�;�f�d�[�0R��n��)ԬU��<��Z�}	���*Xw�K,�:��9�k4���$���1�Yf�-n#sI��!���r�iL���/C&�1I��4�L
��03v�z*�:I:0�1�9�v(�opnBO$ٙ�[���Y���Ė���`�t��iJ�8^�N ����.Q3&�p-2���/&�
���5齁T�\ 鹵$jb{u�7�r�ǵq ��V��5��wJ�U [J�1�ʁ9�q��4���5�*y��LO%�m��mdD�<T�����p��R�½��Tr�a�n]��W��LZ
�OPS<B́�FÔf�ɖ��U��&C�)�͢�c�E��JW�n̔q%f;{*�.^V�����vÒf�:���SX�w����݃w��Ђd.@��HS�*�L��T;m�{��V�w��ئ�-�� ��G���j��u��툷�e\��d{V��o�'ZS{�r�#]�T�b�3�##�H�b�6��lY-�T]@R�������MU�5���Z�C4,T�ѭ�W�Z��][��b̩��
J��
���m�.ŕ,~���v�An۵y@`�	�HL6)=��L�ē���fSF��r�"r���xԭ���EL�	v��D���B�Όm��u(��eo®�����D'���n�X��G(��!`ֳ��x*��,k�T h�a;L+����b�0����m��M��6N��Z�� �fi.��ʅb��+2d�87V<�:�C:�^���O��˺ț�ۚ�eA�#v��j�b=ͭ	c�wM�O%�a�N������cq�N�b��VT2��3��4�Es:Lg�;��n<�+�T��������hXAS%d[�k4
5�&�N�CJ�r��J�
�P4d�5 �_;��X�Hm�۔dOH���k�ԻSJ��1��,��d�����	��j�<�j���o-B�Pń�֌��Q�JbEQf�@�K�
�=�����[��n��J@cD�ۇ^����Gxo����hM7fn��]U��V䣎��c���*Ŗ�QA5͆"�Xŭ�e�if�Ьt�Ҳ�\gI��R��X�($���bG��mI1F�f��vU��:t�`�M�ޅyŬ�7����S���:��|&ma���e�܂LM�P�� ����-V�L-�l駆ȩ�#�Qj�SȮ�%���KE���F�t�i2����s2�e�P���Y�P�sL��@�*� �A��a�ڨsH�)�d�x��I�3��͘�w��&
&��ZG,
��b`+�R���/Cvfnִ��:F���̴V��z�0��CFm;;O-Ku��cj'y���L��Jko`n5^l�ٻ��v�M�2a�Wn�(�mRIiӿ:kv��e��ĴV�]M|�5S][�J�GN�,V hau�r����1A�+"��&�ʕ��ЙF���M��;z�MR�>Pm:�a5jR������4��R����4�4�[A,D�2��-f*:َ�NQ���횽5�j*���7�����<���U�$pʍ9@�{L�������md�z7y6Ém
�<�1T�25L:]�I�J�5t���Ǳ�A�}���h^@�"7eb�,,Yv�1Y�b�jlʓa�
9�V���+b�����q���i-��q4"�:A_�n�XNZ�Ջ�N��٨͐ǻt��n���o�I}��7P��vV���Ǝ�K>T��5�:��SK&F0��uX+i$$U�J�tZǖ�㠒;��P�Ԫ�؆���"Y��ڷRS��,�e-GE�]�`V�u��"���."rS�[Y��Xz�����ϳvhF�C�� *me��&'VrY�T���q�A�Kv�*�����w�WH"�+4�cof�5"qZ�[�[�*�-���UjDA�Q�5��e*�, "����v�5�u,�`�i�K5 �%��]�I��&�C&�T8��`Te�(˖�n�BӲi��w��d5{LYt6�XB�4eC���e�`��N!��&��	���BZ#%Y����c7
�- �/^
��\���VnU�o/
���^�u �\�]iqw������?�QT5e��El��z�Q���uh8B��a���f��eҫQ�|��ZK�d1[@"����$�lf�&&H9��K�;{K.���U>�~��V�|�z2SQG 	fEa��Շ��l�R�ڽ+x�^�U�GOsR�x�+�ҽn�f�K(�{Ad�FX%�V�ߋ4��ös1kة��]�J�*������y���!��1:�������z�n�$śn�-��Gf����R�tCUvm�Pf=M�j��+^ϞE��������$�lH�I5F���
�l�OcR�R�s4�:����L�0����+�!4�-��3@���r�ɶ�ء��V�k�1����+ N���82���b�k-Y�I^
��b��!ӷ+f���mmd�F��0�g@�4�2f"�[i�k]�1�[���VXX�Sr҂���ԮGR�80��r52�jl hT�0n�B��JY���B+J銽;�b �T n&J;�s`SҰޡ��c��Z�F�)�f��8���(�-�ţf�����{)���6��΢�l��!���,b�t�+��e�C^�A{���b�ؖ�&�h-��ތ%h4$y�]��)��4U����R�p���(	j`���F*�K@n
@��R�l&�T�e��v,��j0��VP�l%+*�M��7���d��(
�:i[R2�mC2;sf���MP�V&�NA��.1Oe=��n%�ulFr��$y�Mb�f��kߠbK���7!�Bȗ�TJy�q�8�cY��S2��:͠7NW���D4&-eS �-��31�������:�ʁ�2�l��ܘfH��L5*��P�H1��t4nX�
1,^fQ? ~ ���5@R0F�B�z���劆{A���
��㬎��p*�lӡCZr]���wX�ٛ��ZػT�Z�ô7iQ�.��z򮓫d�k@��y@D.ުIR��I�E�V�x�aš�őB0���b�� ���d"����d�N�в�k&���fh5NVd�c,��Hd���
��q"�U��	I1E����,L���o`qg���a��9>��*0�@��wD�Z4E��SE���cy��ʉ��S�O1�X@up���*�`ϖf\�+Tnj����Z�f;�ɱ�b=�*IIP��N�̱.%Y��Z4u6ZP߬�F�ѹu��Bn9q�ɲ� �ϞA(榵��5b�d��`x�M�sh��.a�L'��Ux�z]�?$+lc��8�����w��Q�#X�QWݢ�#@Ð�Cq]Ɏ��p��½��*Щ*^[v�᭐�Q�)�[Qդ�n�"��J�jT���[Gu�Z˙G.*'whPX�r$.Y{�]d�tc8��������nջ��I���yW��j��m+�̴�͛�J��Z&�?�p��m>�F]�����R.��!B�QT.;C˓�����ը�K�8��&p�l=��.Vn㏮��Z7`��T���o���oCGz�Vqťp��Q���.�xN��.�A՛��;����B[�EU��+�}jd6K���q���Υ�y���uxw����`H#�E? 5n�;Eõ�ꅫʵ��"�x�[��gN�+��IAu���um��]�p�h�&XņE�@�c �=o���o6U�L���!Ċ�U+j��~՜�[�1�xz�d:nd���[W�a��5�Q<�T]B�ٝRĮ�F��;:�iiw[��9��`�S[�n$�R��\Y6Q�Y�kuG��dD�J���su>��{�Ĕ���,�j�b��p��[�u]��;l:}�/ga�\�2^e��m��B[��;��w|���Qd������^��w�m�g�y�K�+�,�̛���vʨ��1+6�Ų�}b�k�U�9�V����#Ov��t&6cܼ����[R��*��xw�ɠ�O�ܛ2�Z�$Ku�:�x:����n�y�т�.�`sE�q�����A��E�p͂\'+�i�q,;U���r9؋2e���l9eE\�Qf�s�qkp?�C/Ywpm{oǰ�{�t�6�D5/7��|�qU��}b�n������0g.U�*cS�����6j�R<$�G��a?J+�@�ыqut�#����\�
y���[=]ϲ�H����jP���V�8���Y��]F�"�h}zܒM�W�2]a�_9>#4ͷ(p�մe�իTk����Ȕ�� ����B��Vd����Q]G,f��n�t�۩w�&�Lu�5���WaWK�[`�3������yW�D1)����푖:VA�ū�n༫��0H��&u|��M����R��	s�UU���o-��!�˦s:��Y�j9O�fm�j�8)=F��s�e�����i�o�#���p�67�jڭ�Q'�w�o>{"�� ���8H���^�n�<(���O#���i�\���ܽ���*���hl��`�m���#l���o����v���8�W1p&j7N#�� ���M�yC��3������Y�M��v��y6��S*= �h�ŝ�
����y��Xs��;q�ʵj;���eʺ��8e�qrk\�2�6��k]��bM��X�j�f���P���;-�t�A�s�!X}�j>e��H�ˬV��lJ5̨_H��a��մ��k��j�@��fH�q_7�׷\��un��K7�j��*�q���A7Z,�WJU�j��/h�UJ���h��R�$f�f��V'a�KҲ�,��tE��m�q �fU�C�g`��'�+ٶ���]��9��d0�VXx��r�]&� ��ܣ����+�8˝�C�ܱ8
o�u���i��Y�YR]�GXz�*��*�k�A�c�X�
���M���dJT5o3T�DP�:���>z�I�#��.U�J��S/�ս��^K�j'FG4��L�J=�f=5�}�cz��o(��Fm�
`��xyD����B��:�C�R7���E���kL����l5 ��/J��R��c{m@�]L(�ok�pr��\�5��{񄽱�jH���NaCCC���Q�������ַb�w'=?+�K+���ŉ��C:b:]�5�7S����R�ݗmL�&���f>˫쇅��MvCF���xUt����`������K�8�ӳ��k@]ʲ�ʥQ�L}c���уt�'��XJF�,u"��[�1��z��F�C#�o��m��]�se�d������8�3wʱ��y80R�˥�M�ۺ�
���H������K��QT$��r�����Ɩ��A�,��$Y#�+����fK�5����j�3��%Kek��P=��T8%��R�%��@��v��m֐Q�y0�0>��A���s7]'�8��l&/�D�u�V}�Ol�
�E+Nq����2h]��+�@+Im�\Ut�#t��H"�d�3��>���M��֐� �ԻL۽d��Z�L1����}�C��L"�h���ɋoRf1�z	����;�\և$	پeC��"����;j��(�,w�5g��A���0+��1�I�Xq�gvZ�H
�$oE��y^�����a��	���F^�x��Z�Éқ�l���F<��N1W�A�7fzhb�:�LKp4ֱ]7d� ��p������3y]]�3�2�t4<�b��j��������e-o.};Dy/Q$�}�ث��d������\ZA-]��[;}S�����6�l�iC��yEJ�3�vf����
E\[���B3MƖ:@$N�]r�;�����S���DХY\_ZO���6ܷ.��4��E��a��rY����f+�d�rf�n�|9���)?==��d��w�Zg���x.�z��p��"���(�+�����i���"�0������φ�:��E����;"�o�v�2
o�[g`C#�k�Dљ �V�V���,ղ`����Z�A���Wq.��[X���BɷX��OC�A�{2-���a%�1�jnM_y|}�(f�A��(l-"�;�]�}� �%�`���^��#� �ދ����;���k�x#+��q�[����$�1��t2�4��	�&D��I(\��I'� ]*fg+��d��4k��hN���ud�]�c5Y�����]r�ĵe`!1�/皆)��x�묫��X}��I%��R�� ͺ�)Xa!On�o4%o8�!X5��c[�3���/�n����\�*��%�̥�+q��g[��	�h>ƇAw��Wo\G�ՀNLv6:L�Y���7l{�g�0X>�����b`�Q��f���(\y>�`r�^|red2��֔��u�YC�Z�1��͸Y�r��h�L�k'Y���L#��h.�r?o�w�xz\����X~)��b�}�k0�Qʳ�v��B�6[�ʏ���B�"��y��Mh�ofѼ�U��:26�^ȵ?�J�X:��^mᙺh:7݇H��_A`I�S���n(�o:�O{8*V�g/k��7�n���{Qkl��(���a�ٛ:;�cQq�'3��b\��F�l��z�ٌ��ˆ!I�M��X�mG�W),������ԡ}����Ǎ-Ys�uvJ�"\	u;K\B��[��"��縩�s-a��Ǔ)s�W*��U�_45c��0mh3��\N��WiȮPn?�o):�aV��p�L��9Ԏ�.�s����Af�#E��nLA0٩�
\L�'�Ȩ�l�Sy�B����9�x�������k\YgFr����+��ܓ�;��'��9G�բJ7�^�q+$N���ZV35K�$��Qu��^mIX�ŚV>�Qb��F�����xMK�:�/��}�K;pK]s��	��^B-yZ�]{j;�X�WaUa�ݻ7�:�j�,yjh�]7����'vTZ�ګ���ge��{5��n{Mzm�C~���'o?t^+�����H�=�R���Y���]di��5%�D(:u,�i���J��N���c�oU���KH�Jwa�Wb{��Z����{�����+��ewD 5��{�3��+A�z^<�<��,��m��ݗ���K�g	V"�}���|{���Ψrr�	��]y�vs��
3���E�P���K[���+��l���ЬnV�E�2��,w�ʙ�����s1�~q�����&���ԴƧ�����=g�7lug:�S�]c���c�H�u5�6° �����RXS�����/(˘�c)�dwn6!k�I��1���d`�pt��t�l���Ks�:��GJ\[w7��c�3
ɕӍ��o��Y*89�V.� ��uibŢ:�P�	��7{gw����c����Z�ȕ	���w����2���UbΚ��0oR��T ̩n���-EAm��� � ��X�BK��C,z�*�[׳�O!X00Y�:v��'�;Ԕ�$��1SY�^�!�p>�5�f>��]��бsrb���;���_s�xlò��n4p&�JeI,�g.��\�nT���ne�WX�qW�,D����]��=L%���kd�$�r�v�}m�ėxu��������١�6w��`�]0��7m�(�D��K{�:��v��ω�u�qS�w�A�3����ˑ$��r��6�| oTwN��y2����;���7ɟ��q���բ��Z�o1!��|q7�2�����岡;��)G] ګ��}�Y)��v�!�E����+�7r�Z�����bs��`Yח�S�2�s����(���:�=-��O^�B��qV���������M3|v$���x<�tP=Ƶ4�e�s������r�}y�X��X)��D5�V�t+F�+z(^Ҋ�P���d�<�X �s����W�7�V�]���^�Ç5�a~~�@��}�Ur�d$��y"��z7S��*R�]m4����I7�s��KU�v�B��*V(ۭs
������P2���AH��^��4�Aȳ3�A\Xn�A�$Ѥ3O�t^����ٲ��^�0���4f��v�̽�;�8�b�ΡmCkrnq�1�;���6��PA&2����7��H��P�4ڭ�{�nku�-��M��}@v5#q��"���n�_��H<��g8�� ����_.�ޱ�M�M���1]�Ce��"�9�)yK�t��,�OfZu�W����<��j�M*��x�E�k��u�Q��kM��h�f�DT����H�-놈I��i�i1��c�$�� �����Kw�gu���i}`�����g�U�����L8�0Fj.��rѾ��Y:�%1;�4�fF�j+S�8,����ⲷSͫ<��/��R�����q�pň ��:Br�9�0;U��s��u�ꙉ�<C�"X\���|�r*�\��%���K��i2F�l��5���k1n��#עN;��\��Vf.�̊��XKF3�R�B��)��7@9��w�+����7l\��e���He,���d�4Rt!PD����2Wm�Hq�Rr���*��Yu���:���|�����;��4N�#�YL���8��Rj󬽀C�f�DS�����H��1��8k��VZH@�[���������Q�����<<D [�1RjzZi)hvT���imu���+���#opv�,ˍE��IcZu�p⏅s�za��X�Y���ǧT��!s��]��.TU�y1[`p:�Ý��%J&��
�(R��Sv����S�Zj���|άA%S��`'av��4�늃�\�\��}K;d�a�	�7�u�B�S���
^�s��5NXTG	i2�`�ԩm�޵Mwv�ccPJPJ��%��V.ɽE��J9���p�s�	�h��)}�E�L%��s�t�\j�ٕw�HS�]޻�Q)&�x���VҜ[���^Q�,:��WU�.���f�Q,6M#8�x���b�\�7�T`���X���n�Ek��f`�m5:2�f`k�����l�.�
�G��T6X!�Y�
�*ѝ�t�;��o
���@�y�����Od�n�{�}���.����B�v���.q��R�
��_�I�F��;�ѽ��d��{���â9ho���'J�q&z+s��Ok�*��u����7X8\��p`Jo�L�Ɲf[$�F��:Mj�:����/�ԧT�}��)[�TW&�6!�b�y9l����i4ɫ'5#�é1�L�,N	V�B���	��o�L㓢Պ��V<�����e�������Mrӗ��)���OOv��-G�c'�
���I2�#os�F�U�FӴޣ�B��O�����3I�@I����`el�-Kf	|K�:6k��1���Z��Ђ��)���6N@l�����A����8���,J��.�o�,j�	6�	�8K���+GC�y\��Z�f�D�	�膨��s4d;f�[���z�VhX����e��\��56Z���͏�����[g1*���s��y�zVR4����Gb��6�O:���'lP,��W����E�y��s+����y�X\z�4\����ҷ�,
p�{��-4�NKZ�^�앝]�"u�!(�Է_kF��S=���,����w�s�6��#W�uG3���+���D<�[��x�l!yg�uqzi�ĭ��,����C�����w5a�\Zܒ�����(
r���UM�Y��ё���ӗ�z�%t��Pe -�D>ŝPF��<�&L���F�еy�ā�N�}Kp1=03�{$���(q�q�L��
�FEˎ��jP��ʓ/R3^w�6/fW.����"���wN��5�$�.-H#JCƖ���Է�,:�5�KX�'ْXb��ɾg��q^�ب�ؖu�z�Άۻ���z'Qq�-�g<qD*+w`���-��6�^��Y#�6^exʂ�:�u��[X��z�����.Qįr�(���kue��mfm���Fٜy7Ң�r*�>�xm`fP�}b���,ӥ	wB�q����bΔt�ȃ`�ۯLķ�B��0N�\�,���oL�:�9 k.!%�P�}�iE�U���l�.�37�ۓu�b,iL�W�y��F�X/6�S�|�]���\4;��m��m��-�m�Ռ{�4�:K}���y�Q\��ы�.�F�륰���S���;�D�=֬8ߦ혪f�V^2v'�)�E����ە�k�X�k' ���\��|��[l)�a�� V���mï!�� M;w�l�ֽ�~�u�l��H@$$?�	!�����ń�G?/�k�k�]�1橝["��)�/ �f�Ta����.�V�y��kg�����Ƃ��J1̭�-�$��!g�ܒD㳷�|RfL�hڂE�$���b�:�+g����h���Fh��O`9�$����II�X�ΘF�X�d�0�8H�W�>��#rV=GqJ�4�*�7�]�y��|�쪒O�@l�uj����>y;fNf�@�
��Q:����Y{`殌�H�΢� �����{�#���S��}cWy�m �r�i�^���X�kEo/#�n�=����+T��v_mY������*���N]I]])v��q�m���ϕ��r\ىu��f�o]7-ݱr���}uN=�a�t�n]K�ݝz��x�w49o�'o�%��ī�w��2�k���^2QaD��E����]M@F�W����) �v;��۴RB��D9=���Yd�X���i���ғk�[ڵc3�+L�K����V���
4&�V�U�F���yBR����vL��H�q6s�`ȃΒn���Eb* �։�A���> 8\�g�k}ːg�qrKm�K��3n�M�+V�lˈc�޷�ifړ������'�f������bp��"��:_-*'�eŔxs:1I���������YE������'��qʕ�X�]52���4�$���a՜"�Rͧ�Zȸ�qN�+!��<��fA����N�ה-l�ۏ/DB�b�p8���[;,��Wv	l���"��{�<�Yn���V��gN���k2��$o�S+`�;���M��3eG��	y�a2�9$`3ј�sY�xBચ�OQ}-��}��b^k��`��7J�]C/Y��puwu��J�=]������q�_d��:��}ھ���D��ٕ|�MqpoPv��Ν0���۹"�j��y�}�1��ϕ݁���D�z�*ebzH5-	yz�o]��u�<� f��ygY[��tc27Q"�o�f.]���8-�Gl�+�}l�U��y�B24f=��t1�ʶAgW�-��sI��<��� t��h���P6�Z�n�iqՕ)�J֋����-���S�����S�.��i��"����լ�҂�;c��xm>w)y~�5AƤ���k�����c�Y���:#�NUU�,t7�&���`��.��ɕ�2k+���B�f��}���y-b⁅8�b>z�UpK�mo��t�r=˽:؞s��=��T΂�X���F����8a��i�ǚ����'LU��E)ǛH�X,�c(��+2�Zo����}Ǳ�\�5%�̌�</�|3�\6O[���-����.>�i66����o���Q���o�X�0��j��S����v:f.�k�j��::�u7I6�ǬSj{���GE�
��r-�P�u���Z=��ͯ��X��=�M�g��@��l�.��K�����;avj���NFԠ���]p����C٢�2.�R��5ao���F��GFS��OJ�+J���۰��cSU��E�'ax�{����x:��1���<x����@fYV�;��WQ��u4C
�@�c7O�R�R*�y]fb�v;�L�'����ۮ�߀r푦��Glê7oI�W#�J�we��m�ܳ՜Ck��T��v�5�%���]����M$� l�HbiK�����Zjƭ=�-��.h����nĎr�P���[Qˇ!��4��e���s��i<)r��VPK7�_�ҁƛ�{K�o�wbqk#Ʋz��y�]�=���@U��.��L�t���Dapu�è�l��7Q�r��X��M��U �f�3gW'��ӓ��Nbǂ�%B�*J�l:ޢu���s�
}W��+κ|᫈lx�mgќ�{G Mm��Ea&�I��ssH]7V8{C�ؐ���
#݋1����{�w�JR*\�r��a���r��h��#�V�U����
~>K(��9FG���9xX�UԳY�|Gd-R�F�ם�N�����,ˋ�(��`�e-#gXY�����[ԉ
m�^��ֶ�t�n�U�2B�VZ�s�r=�Af��
$�q[��Ψ����&��{�hx3�e��^r5������ߡ���&�g���nir����=Xh'���ٲ��k�ڼ���ӏ8��-��>�&2���m��"�QN:��Z9��0)��՞��c���O�1LĦ�d������wlJ��7O7�M��&��كW�Q�� GK�,�O���~\����30S�+����u�啁萍�ᙗ�SW�BTH�lӾ���\��2$��[`��V?��%�OOo93v����	j�����,T��m�&�Y+�un�o-Ů���m4iuX����t;�.�ܝѣ�(���P��R8�1�vݾ��G���]*�@����lmƟ��h�LZ��gr{6-���|�{f�n�q�ޮ��E��KϕJV�}�#�i�����ҤIk��m�̞T]a���j^(Sظ�/.�h6��^�ݙ$������W2:���A$-ZXT��3R=Y�6՜uEb�R��8������Pߕo<�1tlm
t��z��s���r�ĵE�kY�����V:�����Gpu��&��&�w'q	qWf��:
��%�ۈ^Z�$p,��VR%�T2����'���;;j��.��a�o�x��Sz+-���kga��&�p�>̭W��y}�&��RA���lKWN��$K~GiO�����YwDV���N
ky�L��X�3ʾF�}.��f<�(ڜ{9�U����з�$P>�f�NU\�����{V��
·��ǯ ���t�ԁ�ԓ�����ُ�}��ha���S�n������^��q{���=�G���>=3\�[[v�����i�J���ź�N���X�	�7�B��I�3��̙�A[%v�J��I�K��P��m(h��h�}gf�s{�\��4�!kլza���t!RF���v����$��0r��UNOVu
bNɾ`����Ao�]R�����o��M��]��._6�V�+8�x n���w{��R*�ʽ��+��y�]����R����,W���yxo5S���E:<���o[�f.�%��n���a��0��I�\Gt�ɮa��c�@�Hn$�ŀ��p#z�눫#I͔J���i��ԲO��9��GF���;���*��90��~�̦ƚr�+8������!=H�B��\@ym�X�,��e�Y�v�B���e��n���.Zai���"R���s�`!?[ؤ�ht�v�9�(_o�V���:�T�h�wh��RL#�n�+�ܥ����*���R���.�:R�T-�!��+��i�Ӂ�M�{�ǜ �κD(|H�2Z�_<���k��6Q3�5d�n�� o������G��@C`��P�Sf𼕭hJ"�G�Us}:sHEt1p�/.�������M]qut�X��G�杰��D`&oձ�͵]Wk�<�t�*'i�J�`�x���f���w|q�AK���ݨ�@��.��/����T�VQ*�oE`Լ��^�I����3��{��t2�9G����6JTF�A�xA}��Z,*Μ[���p�@�|��� B������mV5)s�����Q��m����g);���w��䱍�E�365���0����B�v�.��0�U��T����8B��K���uS�f7՛����,���q��XY)vK�|r3-A6�����b%��*dК:��WfrǇ�-���Ż�>��#w�Ӿ�z�4�T�$+���bf�e֞���)��2�_H��i�V��k�}�z�7uD�=�vb�V����idG�$VQ�`u�ͪ�zF��]s��!o`2z�U�>TQ(�l�}]��2G�]k˻��(�����Ԫ@���^m�;�13�o1.w&,�N�VE�ݬ{w�8�2�ŭH���͝��fb�\K/9�,���v�0�X���[�B�4V٬�d�.25V�M8���d���&��c�JѪ���%��O2�4�	�\t����}���0tVݴ��zK��m˵��XX�B-5LQ`Z��^���Εqb6[�}ՀhՎ\힃� ��v���y���{�"�4�}�Dt`��KmۤT�9ֳ"��|�}�e_$��g���amR���&���P�a��m�a�2�n��=����Q��|�F�G���++\��|\�{ԫ�]�u��TW�ƏLt�.˻����a�ˢ9 ��ϫJ��n����((�A:�Iw�u���9�^O�����Յ�p�׻��%2k��M�+.,N�\v(�l]�Z�� 4�%Xt�S0�j�S�E����弔x��]����2�3Y���Q����AL�B�m2u`��X���7X�/��wF�Bm�Qѣ_(�%���ha��J��м�V�cf)Yy�$����m�H-�nc�U���,�I���/�����P�|Y��&/+V�!q�Ab:���L$��X�[�v�@p�����+��� ɂ��3���\��{Z=�;�W�`��=��M4Q�U��~������۞���ss�𛸟�k\���:zV�33�3�,n����"{m��w	����� ��Vt�X��Yk/'PJ��2��l�Ȓ�e�3�`�n���
�Į<BnrT�I�{:�r�k-��KGWLu���u.K�_D2b���x��{_��=�����mY۽�n�}�S�\�q�~�5��U�&���&Z�t��Ov�	t5�D���+B�W�/�-�r���Q�2M�g���W��6�T�����t!�$E�v[�g��B��\'�5ܳr�����vlB��Jcĵ�n�Mù�Ru���]�vْ�ŀ� �w�T�n�^�i�ͷ ���%+�dg�D(�ؙm�b�u)}�iK�欽&c�����.y�9N����%y˛�wnQ����
���;-��Qv�V�C��r��M!���7�G�q�'7���+�j�$'�c��9�r�ذ�N��xۼcqF�Z�SX�1@P3�K�}u���$�D\���Vʖ\��XD�5�Q�.��E*��`87��eg�fuǍ�}��SU+BS.�R��<n�\:wy�{�#�:�N�9�GۖM��\Ի�09z�|o�M�wK�gE3#�T�8�dP��T�	\��k���9�RI����v ���2��P�L^1/�ZOu�6�T3m^�jR�X�yM.���VB�z1qv{z�b�.e�.��	�ą�ŉ��O���g!
�ե�?<�rު*�-���ծ6/Ve�K�絒�(�w����SH�j��l����S��SH�,v�f�����)'���g@�	��.0�S�"NM�7�f6�s�����	^���t�˽��iM�\�p���V+5ghЄ}�B�K���7�5�������m`n�1���]qu�`�D$��GE%�k��0�"���)�
�Q��}}���IU�e	ז��W��13�c�(�`�!�R�/QQG��4g2�i�(���x��*fd���������W�����9x�F�\��xn5��=�7G���B��fU�dPS�l�|�'L
�}H��e�A��L��LV�_5̢*�6�G��rg���{��Ou��F>�w��$��0z>
?cFvhR��bpL�&�8����pL��,�[� \�FP��n�<"��9�����(�|�]��;�M��y�d�㘍3U(�e�%�t�o���S;��I�)J���X8�����g�:�2�7L3Leۨ��hM]�f\	yǾ�>��Y�Rׇ�N�V7`���krn�����9��Yi��fq��ɸ�Uo��2�2�P�7orWL� �����ܒ�҄�0z��ʞի{����f5s�7�k	X����ڵ˄Ȳ�CKX�.�[���Z��nMG��_(�3�<n��"�ۭ���3~N�������Y-[�����+m�v�X�L�ՉMUŖw0`���V���}f=W���*DnĜqZ���	^)�Ne[��anqso�'�!�PK�l�����1�)����`2�6J������f�]InA�� dNUz����d�>}�kv�PL�n
q��� �f���{P���U)}����´օ%=W����'-r���t5K[��ԨjVR�gxR�L��/j���<w92�\����#�2;�V;m=���N�`����I����yW���Ю�bwׇ#=0�j�tٲ�܍�����u���7�5�Wb!=��V�ʵS�.׮�z���Hp�HT�'$6u����SǛP���x4�y�-Ρ�x�NX:��vA�f}CZ�����
C0]�:	[im��u�qf �-h��ᵔ8�
�E9sjԲ�����5&�څe+R�+�qs��\@����x��\����]-�Ő��Ą�.��QR��}�
��6n��n�X����/
�	�f�
���Rrԓ�e]�]���|�Hd��HЮ��걦u�c���]�yj*�&d�c>,>��1���=>6�B�2<�H��ӏ\��j�v����!ٕs���	N��[�(�3�ys^�d�9���ޕHY�O�4b��h����	�2��6:�r�W]4�Z��#5��Da� �+�)��$�ڻ����P 5�6�`	gC���Q�]HS�屑S=9s��[
g'vj@J�ah��n�+uf�?m�q���^L����\�	�TΤ5R"��R����>���}��3�=�����י�D�鞔�wj��owءM��8`/ҕs1ɴEt���L��إ`�LٚMلq�kW]�����i�]B�ru(�
����h;��;$��wA��+�d��膃��ؚl�b_<��5A�֣�Qt):#�S��"��W;*�>���gv�.>�{��JI�(�rя2���2Y�xo׮�ijY����=cź+5u���/��0�t�R��$��ЫIҶ�y@IK-�,�gw{յ�S��-U��{�-�
�c���u$�@��Z��v�Nx�v�H��v�E;`��[ϙi^d/0&,^��Qb�Ӽ�a�X�\Tζs�,�%�H��S��bm{xr���w��!�raPR
�m������a�����]](L 69�R�MK�e��M�u��S*-�n��aN�7�{a~O���PQ�,��\���)5��v������j�B��!�\0ղ����N��й.��)�e��םHR��scu&�,���P���"���Y����	��<��k�F�Q_�qm:OF�������e�i�\5;�f!��KV7���#hU��1���w[�eg(N���@n�u6j�B����0p�ԣ9g�h�t��'e��J�Oc�e���؞pѩ�x8�y��� :颫[��qIu�p1�ɯp[)��m�w;^�F���$�I|�J�V�JZ��QF�Edb��J��TV�
��m(�j��PUE*,�Kb�"�)U����+Z��ƵDPA�����(�*(�ZQ��jUj���EZ�IZZ�[KB���2Ҫ��b�ZX(�[j%j�B��ZUF�X���%�Z�m����U�R�����,UPADm�h6��B���5+bTZ[U�ګR��V",�ъ�l�iF�TX�cj�X�E���B��P��T�(�*PDF*#-,Q��B�J2#V�+b�[Q�
+ZQ��[V(�EiF����+XR�B���
�b%V�h6ʊ�lAE�mD�V�jTQU��aX�Uk�Qkke����-Q�D���b����E��Kb���@R���B�,K��Z�����DF
*�2�X~H$?%�����ٶϽL?k��-�F�2=&�T��a}�̫l7����V��<�ͥ�$�Ro���󦦟C�tЕ��?t�w�c���6o�z������b�X�cD_vZ��k�=`U3����	��V 2��K�� ���n�\[�<�X�L�!)x�ʄX�(Kyi!_k5�j�K�<==���B�����e��a`C��]��{eцZ����1��D�Ϡ��p�iJʢ��^�z����༣���w�4�*�;s�׵h�3zR.�$j�-0d)�/.S�_�;I��W`Z���M9h�
���%��P���-3B�^E�u؆�c��Ab�feh�]`o��8���	��C�=8�w�1�O�:�P��
�2���c~�Z��\�F���΃�vRC$+��I�Gu�V�1��ap`K�޼��
�����+��Pܷ*�s����촏��p��4уr�����3 r�ǷC�3�l]���ӧR����|�FO_ٷ�Y���![�ČL��*��ZdK�0;��}�KP�6\�*�_�x���uVԈ��<�=k�{��hXN�W�U�\>��)��V�e�w9C�Rǌ�O�slC�O�}��2B��^�U(����$�p���,t�~v'S��d�zMN=:�ה�6����	����,X�3F:zd�_�)��|����U{�=��Z�8q<\h�9����6q�u��`f��7s=���2X�ļ|��t�mC�=�we��2^����%�d�}�â�v�2�mL�C��b�Z�V<��	��6�����:^ᢻ�sm�{{�Ъ�Ug]��j���t��xī����
�l�,�ST��za���C���d�O�?����s�lz�&:����+	�=���ߨ&f:��^��#K����x�Ӆ�T"��?��ߌ�72��bqj��$IT��94����֫�K_�&�`������	�K��l�8�[����ΰ�𞙜s�z�,x.P ���_��
+;P��n��Ak�^JR�
��)��w\�9Cͅ3<{�S��9�ˇ}:��𩫦zs����&� �$(�iV)H���>^ҙѝKVg���� �e�����Ϧ�TշOՋ��s>������:�!����jS<5���{Ԣ�7�
KoDO��U^-�S����_w������t��%#�L��>~��4�LX����Ϥ�������IK��p�zǹq��t���X�r�ĕ�/-W�w?R��CBt3���j�c�l�K*�Or5i;ޤ5��4_F�ul��6t�u�GÀ�D�f�����$�<�rg1�ϭ���[�%��=c6]�����#�,5;�g����$��n���r��߈�cC���4��60ŕ�^-im>sDl��1u8�dֵ�&�F.��V�g��:�����j��$��O[ҽҺ�SkƚЇ�gVš=��"p�qy������:�p�?Y>�˼pu^ǃ�(l���<Fo�{�DuǞ�F8�]�rM�%����=��Ĳ+ߪX�e�E_�;t��w1o�u�V�����r���?WK�lm���e%y��^�`'�Bح��ᷮw6�~�.����/ý��j��� =���k��=4پҙ��[.�B�8T��G�ܟl��c�束s�0���z�-�
�P:u�L�q�f�;5���Q��+�?����&��s���[������u��V��8��r�x�d��X�=�	W7�e��v�=���
��9��2R|F�b|c��W���=��~�'6Ü����6��ot\N^)ҧ�	��zn�KvB��K�ZV�푧s�#��/<F�!���|��Q������T�I�`�Y엫Y^�y�nb����+/���vZ��O��k-A��wZM����pw�	KD�/x؎�c�3n��S����ݎ�鉞�t��v)�)x�R��`!�O7#�p�F,K����gt�X��gO������0;��(k:it�����\�@ӽ�<��ִ��'����@��g��{$5�rM���A�+Y쿓�W�ܥFpN�6�\8}���;Y���>�����hs����{�����Ӹn�׶�+˹Ԣ�1轮p���}.�o=�3>ވ�{��F$/�������o�K+�˺y,|j��Am�˕~��ySw��X�c���	F���RV�_yr��j�Q���8���]mg�=��q^4章�g_�(nZ�j9"�#��elJF�U���Ɓ[�P�u��C��3�^�x�mu�g�-%t܂Jΐ�<��rY�/{�}7��m�J��Њ�=�߭�Ux�򰟽.�������m����;�I�w'�Y�ҝ�号kʷ�����&�w��j��ﳅ1���#7���tƤ����zl����#^�]d|[���04k+sB�ǚT+];;a ���fC
=S�m�˪m�ƽ�ٹ���#��i��9`�Z���Ωqh�f��_gPZ^;��<J�~��
�+��N�+�B����iִQq�D�w;ǯ~������w0֬���킩�k����s�6���@s��'P�=�A���f��{&�rl�{Ӣ~�8d�/��;�
հ�{��1��.��u�	s��Wl���7�`�s\Ʉ�.�hz�f��:����a��Q��XtB��G\#���;�� ^>C�\����Tx�y��m��w.�f2Y�w��dDg3��\��(��ix�b�s��6�s�w ���׹u�K�zx�.K�ɒ�)�۲�t��]+��\��j�w�:����2����{��|��	%�Rf����e� �w:wc������m�J{C/������jw�dy�ć�k�uV>�j`��W�87�n�Oa>�� S}W\����vf� �:��W�	�7�f���'�9�������94K/�8U��O;�;��Ŧ6�F;:�v�]���AZ�W.�i�:�/z�^f�_:��Cڍi�Eg��wk�l��>�*�m]�t}Ӷ��|��z�q�ޡ�a���0V��S��v�S�e�W��g^�d��%`�B�,At�D�[���]��ˋw��������p�5e�����dOk�ժ�zu%�����[L2��
I��Z�L��StΚl��nV�蛯UIӧ�>~��%�y���^�C��V-�G��w������9�j}o7�O���[�<5\�׾^�k�-�v��^p>���ˑ�/u�Q���3/��(=���r�K�����;jO{��`㘷l�&��St�����]ƅ��D��f޹a��5'�xO{���×װF;��vy�g�:�z���]1�/�>bC�	������ݟjZIBT���zw�!ݓ�'u���Y�F��KZ����ZF����TGu�ڞ���&��띪=��7_����=E�u�s�?��ޯQ�)�Fe���ɾ���{f�9��	��y#�نDG3��2�{�w_�+��I�8�_��/�n|^?w��ns͗+��L�$��	Щ�M��Sӝ���Y��Q���ۅ�_rٜ�R����������X�ΰ�1�^��%�~8��V"@N԰qߊ����J;�t_j�%Hq�_M�hL�� p3���$'P�ٝ�"�X�i*oNupzgH�q}nn�T�ݘяV|���v���=�#;�P,�3%�bw��J�:�`���H�cZ��+�6�<'aӁ9Ԟ�<z������N��#��y�x��%�,��.�($/�^*��ϼ׹�+8lt{<��Q�����{^���77j�L�8e{�6����6�h�A>�g� #�^R���ދշ������F����b��ӟF}C�S����W�9�$���S����M��좞��H��8�>��\�/~�ys�<��˙+�|�i�Tս&���w����e��T����������s�N�ժ��c<���)2:O�CYn�+��l�Ԍ��/�R������U�i��<�[����^�>���^Bz�e
ίA�:\�����+���\�<���`<߰I&�\��Xr�i�k����c�4n������]�3���]'L���fܘ�+<4��]O]k�#;�Y�^�ET�i�a��p�Y����:��u�TϼW�ՌJe�$\������8%�8{�P��үA�EV����y��=|��+{`���pS��s�-ul�y`<������ݗ�䩽�Wg$�vs�&���\�^���`+�>�yf���P1 �p�P��$�� &��~��[��[d69L:�<����p@N����]]k�� ^9��J�󬹽��;N�����r�R��OZz}�Dr���������~�|��s��N\��{�nG/��[�_�n;�~Ĳ�}xdT�w1����m	�s��b��=�I�玽���`�/k&K�0;�ZΚ]:�S��_K�!W��Y�	�M��h���흳^.<2���$��,J�Z�e����ɢ?Wz�y��:������z���9���)�����|�<�%��ѡ���Y}�{��b��;+eש�{�foDi�
�H��_�����1=`����o�9�W,t��-��io�X�d����[;4l��0^Hz��,����]j7���{�"�����d��p��g�n�i�0�U�x��ݑwe��Ofn&S�.�vE�ͻ�����SUz4�"A"&�Hn�n�9���lksE5���)Icj��˘Mf͎��.���3���%$�e��:Q�tk�I�+z(+�=�L)5�B��UY��Mb�dT��K��̸H*s�j�_G+
�뼛�b�ܽ��S=�P�Y��(�a|e>Ng�x�g����Y��s�3!�R��t����n����x}^�azY~3��n@���+�{y�[��%`~�̱�店8���I'o���
��������;��l��Δ��e�´t>��~r�u:g�I�O{s�=5��s*��*T�ƳO��i��3�uK	k�*���7�$�M2����}��n�{ɜ;�tقQ��}݊_ҏP:tP;��ةL��iM��ޯWk�H�n�K�K�����N9�ʃrL��f�Ds:0r��B��������&z?}Z|��U���ym\���o���]Ɇ\��Κ\���*/�^����J���}�\�~�L���3jJ�w�%�StFgJ� �˵��tN{<��e&|�7i���z{�'q�ޒW�
��,I��pȁ��*�����Xٹ�E�����H���*�=�u0�=���VT�/^�~��:hw�E�j<�C�u�`�,* �]�e�%e=��VL��@����E���10\�ȝ�󆋂\��M'Բg��/�zvr��ǅ��C���U�ox?|Lf\����_�ϽǮ��Ks#�)����"��ڋlt�U(���r���m�(p�9���>�;y��Ϲ������RŠ���qy��W�~�-eC�����ۂ=[�g��ͤ���*d\�F�ɻ���gA~��0wpU�zp����k^4���j��~�.����6�����{��[i=������}�{��c+��Ş��2ݴSu%Jc�����t��9�_�[����~��^��/��I��0��D�7չ�����^N���]�񯯥�L_y���r�K�l�s�Gޕ��3ިx���w��h�ެ6yXg3M0���86l=r�N���l��(JTQJ4|H��s���W�Ϊ���^�a-�Lu�����uU���KI�E�݌9�_ӏ��cf�x��_��t���Z��uizc}��а]�Zx;Ce���[�Jc��g\�(,\T���C{�G�e�	k�*9|�5+�f�d�����K�3xvBH@C����`M���NB���cU�6�p�A#7%��g�v	�I��Ej�}�p����p�A�;�w�k�*��MN%7�/8Ӂ8�X]]��!�Zn)��X�Zb�6�G���,Ѡ�Xl5xUi�s�t`:Ҭ�gS�5���v�L��/M�E�y���(�7�Iic���j#q���rƗ&�$�׽z�u#��r�kN�S��`vq��������eEp\9V�۷�\S��I�O6W(
�{�+&�������J��Y{��D]5⺀��J�Ƴ4�j��c�VeX���J�4N������Ȫ��%9�{G�e�f�PkB�U�����`qfYn�Ka�@6 ��[����y��[����Skՙu��cRJ�|e��0�G��a�3��W�reD���P�;s�.͹�n�6La�Q��a�E.�\��n���]�q����GX�Cfcb�pϒ(�Y��,B+��k�f6!^P�p���Y����
Հ�j��,⾃��_'�^.+a)�;EetG�Wz۷i�L��t����<�Wv���M�1!(fu���)���>��w�M��̡um����!��k��vW��W[���K�����1�}����-���r��f�\=���(�dN�U�'�-*�7jMJ�۹����gt��e�D�-�:wx�d?�RbT��׺�CBC}�6U��c����q$����}��ג�]����ϋ<���]ܱ�:kJ��9tWx�tv�硝�HI�E�^yr�I~�n㔣��oU�o�m�P�m6��cC���d�C��f�&=�
���w'Z)���b�-L�&g��!��5}��mm�d7$���
e�l��Xf)X�"�iܫ�<̉���N�غ-��c�*hp�6����K{f�Qj4�U�l�#DH�����а��0t�+�y(������F��zzf�䅩C��D�Gt2�웝�bɚ<Ot�󒣎m`E[�]
'aJ�����iм��R�3%Zzڽ�g@�!w+�c�����0���j}��׺$���8�O���@��axDMR��B𨺫����d2��z�vy��>�[�d���6��J��=�5꫐��c�����|�̫^��|hj�Y��Wgvn8�X���{tr�W�鬩6vj��=F���|x���,�z�gVԵ�N4n�|Æ�˦�q޺��,��AZ�:�4�z٧J:{������ά���pb��4s�����f��s����J�sGa�p˳YP�4��w�H�#w:Mp�^B���wrV�ڡ��|*���v7g�e�c�-�w�S��@��+6Y�Dݵ��ww����3�ݵ((��YhU��b�++kB����VE�iQQ��-�D�T�R�""�b[(�b�V�R�*(Z�Q���-�" �QQAX�F�VeQE`���*1�Z"��Z�`�E��"�@��aR)D)��[h���AAE��أ[[���DV�VA��kD*T��`�l�6±UEU��AImdX��R�PUPX*"1b0R��"����"�����EU��P�X�b1QQb�b�J�Pb��""��,X����#X���
���*1+*(��b���ŀ*��+��EeB(Ā�E"1Uk
�""�*�1D`��
��h�UEX����*�Q(��-+QuWuWv/2�vb�TGB�(�6S���#'�6��{_�Mn�}�,���ǎ���tn�䎖�l��R�\���VOF���6i���s�/�l|����v�����u��[��Y�@낞��VH[��]����5L��
7���ٲ���Փ7��Gw�����nW�77h��b���`b���F�����o�)}�+�8�o�l���ħ-�Og���vU�e>�頹�}p��峜�j^v/ن��t���S窟z�'ջ�U�o	_k:h':�S������pr�V�c/���9
�g꽮�2�h�m�.�������=�t�+�{aӅ{rP� ��������ؼ�rU��r�b3�wN�a�cD����O��.�a�y��腟V��j�{�瑧�*��bĞzs��]N�np��.YPzg:�^rza�*�Y�yr��7��c���'�Ky���v�Ů��+Ǘm�^�6j;[��p�X��5��t/�"=���=;��P 
���}+�l�qFm��\�&�!�%���5`c����T�E�,�w�d����5�[Ԑk)r�׮o�3O���ײ�ܦ��#2Lٚ�l�����͟�[��>�Ǡ䚬�������p�mZO�謰hJ㙽�3MZ,�:�!y_�OtF��*l��S~�j�7Ɓ��Oƅ�|�;d6����UZ�h�|���!�������D�v��k�k��Zr�Ws�M�:�����=�7�R����k��M���N�Y�����mS�Nw�P�z��+�Ù���'N.?g�Ϳ���Y�N�X;���۲y�I��{�$����b��������V櫎s����0��VV{S��MBV�5EΛ�����y�IÏ�m\�䪻���s3ˎh�J��;n���;����`:!s:(�S�^CA�-��lM	��ĭ�jt��^�}�z��ח��]�$��|O=`W{6_l��ɼ�tq��;�n3χi���+$��d�S�d�:ON���ph9���\�]�=�x��8XG���R��+���$�B:'F��z�'3Z��=�lv*��&�<4�ڕm���+�WQc��nW{���8$'u�9sU�vj1�kx�\�^��3�dx����R�\oH[��*m�_l�Ab�\�u���0,����%9��&���yu,�IL��-���o]����;vf{�+����kF��#�e1r�����[���&�p�;@^���K�|���үrf�|�]#$/Ǽߨ���P��3ZǸ�]/A�rX��2�S�~����7����׆9�V}D78f����Lf�ݳ�d��y=���Z��7ƫL³�V�+�OXŤf�Z�r�H������^�߼ܚ���@��W��pM7�nd�7btl�� ���m�aԿgH��I���ws��=�N����35���q��3�]��/B�𱝲�9Թ�vw�I��ƍ^�y�Ҭ���Nh�Vx۟,�[>­�g��QO�~ڃ�[�r��N�@�;�ֽ��Ve�e���%���l��bOM3��6k[���g�҈`^�I�6�����3N����~���s��ֹ�~n��[+ƈxV~�6���D�b���}ˌ]�퀸�aJ}��7ZIf��ʬ�J��)��ɗ��g�<t��ͯ�|L��W�^��쑗����wˈ�xa跍i�[���z��_SZ��+��4/2̴��K�U"êp��\�&t�w��s��o��u@�{3� }{0��D.g~�<�pt˞�^������Ξ���ё*״��o���]�&r�C��K�j���ԙ�$�����cT�.����ry��3��N���佬�.���;"o�_%�nڼ�Xw�d���u_¦��e^�ك��eG����g��?~���F��T������*�W�[�qY�p��w�r��{�|����XOw�d�*I��IRq���Ru��N?�~��@�<g��N�q���Wl�C^���&'Xk��ğ���O�(��?>οO�]�[̽1w�y���~�aP���:{���5�0��8�\�$�XN���M�`~2���2z�t~�6�i|I��l<;��:��n�bV<���ܿe﹗�w߷w�?}�i=a?'~�2q���d*d�+��=d�9�?2N0ެ��$��E���7�8��OS��d�@a�G�GЏ����W�?=U*���w�o����M���gM��h���$��s�:ɴ�{��N$��;�!Rz���rI�OM��W�I���>�u+��}f{��������h���������7��V0�Sl�ɶI����'P_>�|�P�����9�:�ĨN�g�>I�*;܁�'̚>�|�u^����O�8���ӏ�]������;���e�a?:d�t�XN����m	��'�y�O��'P_'��OP��'SL��y9�d�T&��u��}I�<�2|����n����Oߜc��X���.�����H#���@:7v��-*��
�r[Y�0�=6�)�zYP��ذ7��X�ϡ��rEdq�L#Ki�w�W�Tyat:od�f`�M�|��-�F��B�=�À�!�nj���� p=�疲"$ݾ��\�]�5+1�����>�a>_{�������a8���O���'������,�$�+?CT:��OƷ��8�ɩ��O��'R���'uß�u4�=g����N?0����_�_�~�u̹������|��'�OwI�[�:��'ϟ��+'���=jO�8�Bz��:��a6§�8��3҇Y:������I�T�>��I�?w^s3Z������f��nkf�o��i�C���N>���d�O_�9�=�'RO���Xm�������B��2q=�Ld�!���C�,&�����N�`r����~w�}y����{ٳ^o�R|�l��ϲB�|��y�]��a���xɶN�O�6}�?I����*M�?Z2�|�'��!�N&���>C���5��n��6���~�}�Z�]�Ld�zg�d�+P�� q��P�wy!Y:��k�m��Ě;́�2y���6ɯ���VI��Y*M�=g�� ����?=��.���uo��۾@��8���8���jÉ��u�o��}d</0<d�'}����0:��ݼd��&���|�'�4���'L�>XN�޽9�s��������߻o7��s7�IPP�3�+'Xt���N�S
I��OƬ7l���kxd��!�y��'z�s�:��	��so<a����?2z�K��.^Mw�]<��e��}����}@��B�IPP�<IY=J�ٔ��M�XXN2|��a֤�g��6��:����O�!{g�M0������}���k7��}��6���O|�߷��4��y���|ɩ���$�Ւ�a<��aY>J�Rq���Og�	�O��凭a6�鯲B�������Ӿv���{��߾��>�p�	���~�u�l�1��<@��r̞��]�Hu�5�a��u&��IR��}x²m�S,�d�����g���]��{^��Ppf�?:�-ŅZ�t�0I�WA���&��͎��P�shS⽝�N��)��V)Y+LF�D��w���x$����`�l<+9�z�b9����ˆ�s{G�_>��C�%Y��J'r2'Z��r��Z=��gya\�ʊt��s�q��n�<�=�`��v˚�y;A[�󼿾���C�=�$+��a����I�X~�0����\�M$�
CS��T8��;�B��'�5��IĚ��_,����O��U~Ї�l��wߚ>�����#�<N��d����O��aԞ�����:����Y&%a��a�I��gRq!�{�Ԝd�+;�!Rz������߯��/~~p%�~��؟�����^�}4��"�Ǭ�M�d�>��?2u���'Y?$�5`x�̜b��$������I���u�iY���8ϴ�~l�w�����~rN���&�� ��N�翤�d׾d���jn�x��L�q���M0�Ì&��~d�N���2O��'|>��OP��O̓���>z�w��ss�>���~�G�}��d��'�9�6ɶMoϿBz��{��4���2�x�&�����ԩ�ՇXq��kfC�N �jy���:~�� ��АvZ��R�~�������q�����I�}�8�Ϭ'���u�o�=�r̟$��wܒ�z��{I�Y?0����'SFY�I�T�i|! ����ֿe��/���}���w2k�y�I�<�Rq���ϰ'us�f�N�wN�q���s�a��Ou�I�I��y�VO��|���N3Yd=g�N#��=�����^w��G9�n���;��|��w��������'�4y�"ì�J��T���rwvI�^a�N>����M>���|�'H~�e}�?~�w�9�������x{&�����VORq�2���:�2��u�_�u?2M�3y2q+^���'_P���!Y:��]�߬&2k�é6���|��Ͼ��]|�j���A�,Z��6v�w�	Y'����%a�C�i�'�,?���u4e1��N&�P�?$�u��u����8���>�Y:>������>���?a��;}2�14"�"h�Wvf���,.���z�]�0��Y��ޠL�]O��nPD�����x�	�`;F�9Ց���,k�$B:$�Ye]Yg���i4k�O	��/��6wΞ��^���~��z;�'s&�_PN��u�j8Ad`:���'qo�~�� ��'�?'��M��'�s�Ь�i�~�*
��*O�R~�M��'SXY&�q?j�����5���'_S��(?,�����+��Ч]~�ߏ�8��I�{ϝ�x��'�<�:�d�&����f�5;�E�u��T'���VO��~��q�iF��d}\�}��FY�sT3|���ߩ)#������M�$;}��I�<3�i�����8ɦ�y;ܓ��O�~|;��d�g|�
I�59���I2}x��|���P6ì�?�<�����3)ǧ|��s�~�|޺I������M���`q&?2x�����I��<�I�I����l=`y��V�z����2k��	�}����>G�~=ɾ�NbW=T��������4�����y`t�O:ɷ�c	�M��P��'Y:�����&�j{�?I1���N��$��c'Rw�
��z��N�T��{���?g�߿��?�׻;�=��z~d���a++	��"ɷ��Ru�>���:��C�j��Y4��<=�@�:����I1��ϲu�$��o�u��)w�<>�7��y���;<�aP���T=��,<d�u��h��_,���$Y=|@��d�|MN��'ڧ��&�q'���=M2u���ΰ�B��������L�y���:_�k}�AI1;��|�ĨM�Oq��<7� ������I�M��ua8ϒ)4���6e�'�S�?$���~�4�?}��!_�*������}�p���d��m������7�:��|�ygRq����rx�l�}d��p�m�[�|�:ɣ�0����'S̡��}O������mb̮���喿O�}�?oY��v��Oڧ����N���6��/�kq'Xh��:�d��ɾ��N2���d�'��6s���|�s̒�z���'�d�����_��.VS�k���\�$
�6��%$��p��5���������iq�q�bvY�Z���ɿk��d�F���
ǖ����"���yPԬ���+�O:wc��ʛ���V i��(����ǁ��s<7���RQ�}�����1��$>O8�ɔ8�u�?j�lY'�d�'�o �2u*y���:�S���i��7�:ɿl'��ì�d��}������ﴮs�~'����(yd�a��ﹽ�߽%d��(u��������N3Yf�M�S��:��g�2u*C^o ��'��=�N0���]�N��s0�'}����]]���s�\�����{�W�q���7�I�I���a*M�?[��|Èk,����ї'�G�����C�8����2
N�w�w쐬�a�ˡۇ����M��������̓�/�|��Y6�߻�I�Mߟ���l�Y+�=-��Y>Aa����u'�.0�I��Ld�n�8�������۽�f=޾~�wϮ��m�����B�m��N2~d�`;d�'����q6��u��&��?d��	���� ��-!�d�jad�a�r�Z�.���޾5�����=���ޅLa>gṡ>��<��N2m��s |�~��;I�'�Oܤ�6ɦ�f���M2w��V�}��*
&��+'�Y;�������y���]������T��q;��m�Y�T6�I����6�߬��y�XI����'�'��z�ğ {��M2|��x�$:�I5���,��{�;�׿sW�k����?o��n��	߮�T�eI�(I�M������3��:�I����I�̝C|��'�p3�i�Y'<��ɶ�w�N��OPY�歾]��{�����o�y�}	�����䟷���I3�ĕ&�Y?L��'̝:?XN |��,��'Y8����'�7=�'LN��i��I8����n��ϵ��{����M�x�!ٿ��z��s��|ɩ�0��:�A�2J����vE�~X�Rq��O_Χ�l���ğ�6������'�{����k�g�k�{�������y��m��_tЩŤdY&r�d�[�5>㜎e��[���$y�ٙE���i�2�"6'��Ǥ˸�o��`�"HjR⍮s���)Sh�014t��6�W�y��r������.l�͹�=#��}���V��:f�ӓ�,?��1+��$�	�7�~d���T8��V�0�I�'���$���]2N}dY;�fP�i<}O?Xi��~�y�%�?����[����z���D}|��}�>M2m�z�|¡��è,���p�&�X�q'��}�a
��O{�N�oVJ�s{��>�}��o�jJ��~f~�����V�~����|����z�~�=g�O�u'��́�i��/ۤ���9�:��z�y�d�T&���ԛI�*w��O�5���}�� Y�mV��DS5Oo窩��Í��M�r�x��I�������I�'�[��i��P<�Y'�u��/ߩ'�u�ܝM2O��ϰ�'�;������_-ćh���������瘟��̞~�0�0;�'�I����YY�M%gY'�Y�����C8���7�|�:��}�	ĝC\����I�7��ߓ�xO�1C����]��ɞ�\>��v}�8��M�I�k�'X$����IY<`~�'�I�'��'������q��
��C�,�?|`u��,�7�Q�#�~DF}G˙���`!�qήf��Bi'v}��d�a��a�N�����d�O_�9�=�'RO�3Y%a�AC�VO�qr�z��8�+$��!�	�|�S7���Z'�Ûބ�g~��BV}���M����HVN�����i'Xx^d��d�'�v��l���~��'��T�H{-�Y>b���>A���"�Y�W1�=?0��
?}� Ya�c$��wl�J���0<@�'~���
��5�6��bMw��i<d���Bm�d����+$�k��J�i�s�}>s\���矼��fyوVOXt���&�XY'�6��VO̓m��q�yCL�d�=���:y���OY?2x� ��Oi�i'�'���֎_����:�����E�f�x�������8��v����Q~rq�Y
M�V�w^}ҋ�����.����\�;�� e���K�{��^�7���WǪ��K��w:�ƻ;��N�3Oi����Zȭ�ft�f7C3�Zк�5�IA.sY��}B������=�T&��VO�X~���M��&�u=5a�d�g��m��̇���N$����N�|�k�ͼd���|z�($�T�Wy��싯�}��>����N&�4o���uu��(Lޤ��%d����M��'>Oua֤�g�o!�����:�=x���\��������V�w�������A���z���a:�2|ř��z�����$�9�IR��'VO��xe':ɿ���a8��x�ְ�A�����Wf~b�
�m�����}�E��?�����0�i�d�;Ld�O9��*�=Af�ܐ�2jwX~d�I��d�*I�^0��|@�e���2w�;��og~�0��{���=����01�՚~d�y=�HWi4�S߳�����a�a?&�ܚI���{��q��w��I�N~�N$�VK�$��_�����g�;��;������&�:e��N���y?X|��CL�����R{����'P��y�I�X~9�Ad���ru'R��ORq��<�0�I�O?w�|z�~յ�~��{}�^~����}�-}�$��;dXx�ɴ�Xq�x��0���C�S��&�q����=f�8����'�u��7�PY&'���M�d5�׊?�a�r�wg�lR���g︄~�� |ɯ����l���]0�OCv�Ԛf����u5冘q��j���N��O=�$�2q���z�}�k��t��{�vg�?o�ӌ�ht���'R��}���>~I�X2|ɳ~}����	댚d�VOR~g�,�$�*i�Xq����q�纻�>���������\��s���@��̀ ��B>�9��?$�!���Y9�����u���~I>d�'ϝ�$���z�ֲc!�YY���Y�I�T�6���W��K-��G�tl�8�jyAÆ�q#L�ߡ*�jV�B̼��4�gT-D�F͋d�%[�{ej��{H�vgH+E �jk/Y�/�:��9��� �Gs���;r�����\�����@ >��VX�Z赁,Z��i�����U-��%����];�w"d�O�%9����%awz�S(ڥ�d4���З7\SNV�0�ee�.n�R��x�e!�l�__7m�r��<��㜺���i�������J��n��l�b�؝�:D�s%�0�C)�����l��ܮ�0,��|bX)�k��2�eK�f�ҫ�)tO�k���W)M�%	�ʌp7�v�18��
�e�K[{�wGT�.�V�r�m�:�wVBd��g�Clu�k�k-�:�
Z�e_i3��D�L�iƝ;����j�u�0Pv3�D���Z8��+����\[T��SߤJ�D\�R��^�}��]�u�D�7������d}q���N�3<"pRʜ!S��)��y��z+%`3�����@�pe�{x.��U��f�ry!�"�Q��7&s��]��X�t�Y�}�:�
�Çs��?>�1ڼrO{�]Z/c�W[��sq�η{:[��LA1Ǯ$�}��l�&gf�����)#��%�N��fI!|-��*��n;�֢>'/�Β�,��k��K�h�jñ�CA��rw&\Ǵ�u��s���� o��$��aS>�K�d{��Ҕ��#�p
�э�s5woSl��ʄj���ިZ�Tŉ*ǜ�T��S�=vY�'N��kkSǞ�7�"�V����kɠVN��&\Y8�h���P�����_�u��:p;�����\��1�g�3)C�%FFO
^�V�	�c�s�(T-e� ��FF>|�^(��HWC��S���-hRMT.�fN.��9-�
�E����r�j�J;w!�I;�j얫���-�8_*��g��w���
j��K��
E5�o4�4M#H�ɥ��lvMDo��)�a�4Z#�}��n���f8O`��51��,:�R�g�2��U���$��Yը�s)-4ܓo8�}VC�.���@�˝�Պ*N��d���ja9��5��~^�8Q����}��œH�,PT�t�jU�l�&�*y��<�b���o_G�����d�v=X�:��
�جxp�H�RW���q����E�V��Y]{�U��_�`5�.
��PtOZ��d���\`eJ��ۜ�|s��=��Q�>�/`'��}+�'�e�O�;� Y�v\����Ct
m��j�n`�D���D��*�6�a�u�k1�} �����s������+�<��/Dj�:�s-���_'�w�l��癍�Smm��U�D�we�C�}�u�%�Nj�Lmz1���;�A����Ls��{&�H��n<r\��"檾�˰��-`T�VB�*
�R�Q�#hV��Qb#��`�����Q�%dF,QIm
�+AER#mR,PF)R�*�(ȪER*>��J��fĬ�@m#.%��`��PQV��.Z
#l�b�+&%b���b��&!b
EX�,TH��%aV �A�Jʂʅk%DD�h���Db0c"��*�2Հ�R���b����Ȩ�ATQ� �"�YQ�P�TUFFZ6UPX,EaYX��7,�#Y�%QEUAV,+l�F,-��Z�`��T�E`�ZA\�cZ ���E��H�,UƢ�2*�Q�+"�"(��*ȸ�QX,Q�(�%QA���5�i�������&�ݗ�xջ�(�ϕ��Eb8���wm%��p�U��nP�B0��U&X�T9�2�����OL��O��Aw�{����k�
�����Ğ��k���d�Vh���:��~ì�	�xu���'��Πu��=w��u�|�3̒�x��n��Y?$�=����������~����3�N%k$�3��m$��ء�N�`jy�"Ì�J�s�!P:���'wd�a�N�q��i�''{��8�q�������y����������+����u&�RAD}���S.C�~��(\����?5����Y��������e�G��Ί;!3�L�B{��=��^���K��~���LV��{*�2��{,��!}���Z���ߗM?f�9��.����̉�ϥ�z9�*\w}3�Ğ��B���y�Z���1`���^��'�^���^>�.gbw����I/j\�
`n�ϵ� ��'�:�������
Lۨ*J�4���0oM�T|ew�+��X�3	����S�S*s�x��fY�as�}C/�{�W}�h��#��/�xx/M�vg�՘�=Y�:�	�j�V�<��#�.|��Z�홛��	v�����}<��'N�n�#K���Ƶ�h�su��a.�TX��[f��3�Ç�e��+@�H���N��Щ\	�_	V1dx���\%&�{�a�d����=�I*�9u{oz�Z}B�����Ǣf ����C{3�D�������"0�����k�_��ڳ%)��T������0����w�h�'��W�lٌ_��0�
��x�}OԳ�W��ε��LU���%�Վ�r�m�����k&�����7�x��{�L~:B���ʱ[��p��{��sxe��{|3ײ�r�u/��3s�n������;�]֚��o�\{�i��}�vxоV���k�6ܷR���I�W�$k:F����*����:�N+7A��Z�q�}l!Z7�6��S����7�S%��twl�I~O�|�ۃN� ����A޾l��z���[֣#F�gm-����Ü����s�u�W3�v�~�@N��dSO��:�a�^8�x��jf{��}��(\�u/z�HX0��#�р랩V�������U�t��\=���zEPǮ�v�sL�s#������3�L�~wK������-�\o\;����
�J��1Eŉ����X�$��L�o�$!�R�i�.����Lk��Od�)��t%;p̧��#���.���}�2�>�n7�+��@��SUk]���V�kx�-+{��0���
N ��ﯾ]�_���/o�s����u}�p�<��z�t��/k�d�x~�d��k��|*YFt���t��B����3��� ]w��rYٕ��Z^A�c�@�yS*mإ-�P�0������:��u���QS��ө疼�;\,s=�&�ʖ�\;()�V1G4���#����c܏��3'?wwr1�ua�b����3�wN�a�{^8:/���k�|��;/�>�u�+��oN/�O&�$�����_a�E�Y����V�]�<��n,ͼ��~�0{=�E������?u�䊮&�;�2b�s6c��^����>_;]O���R�������{6l��c�{�S2���)�/��{y%c��^Q�ϋ��u��}��n׻��Y�t�cP�=��c�@���6Nڙ�Õ�4�z����xF �w�&m?�^����&�����p��|����w)*Y�;wc��{Y/2�[�qL�JN�6���V��(��:�$�!��w\��3l�\�b޳z}���e(óB���)�Z��uw]�X���Cx�����߹8Nw&ecP����}��<���Ǚ�����߹G�$o{�z��n��\��c��=R�W��מ�Η���}�}�9��7|\{�z�-�Gx�d'{2�f�Ulm$�̟8+���́�'�M2�MQ�_1�������^���A��R�St��0P����/�m͞]�J��s<y���"��YW�eg�u�}�1%���9j����B����E�-��B{�]\���]r�=�i�K��'�(�$�ǧ��`I�,	d!��-�#��B��d��������:�{#ׯyӼ��h�Y��{��ب?<%�頦��l���>�ՎSc܎�m�p^]�c�.1d�`rM�q�:�]o��n܃�_P��;$mj�u+P��L�����hs�Ôŉx_�PwO�}O���J@��c�S�].y쮔.�y�'��*##�c�}L�ί��EY>�Ew��x���=��>�^j�� �ydIR���>�����ե�Yږ;��lS'	�u��]���w�PY��dJ�2�^�T':��gNɲ��&xH�mE�#��MG�]��d��m
P���t孵y)���P�z������=�=�{��	�|��G�ߞʹw3{e�����>�JG}��A�{&��	�����"�i��4��G&|v�����}tud�:�,��x��ߞ��Q��~�Q��oT:B��~�7݂�]L}*���<�0o��o���m�u/�>���η���}^�9%4��We���o4���2�*cxgHy��sG��I
�=�aϏۃ�H�I�O`}�Vxۋ*_˝l/�C��fߦOzx�����*�s(f^�eH�2r������+Q|;��<�,ҕ�/u��}����;Ä�u������a�g���t�p[_]*Z� s9�v�9M�]P��Ւ��ޛa����*Y����T����of��9���oW׵�]�pn�W�KVk���Q�}h���w�>>�ީ2A,���Ϫ��k���.��W��t���6j1��o��s.�kM�(;�C7��f���ua 4�kv!@4���Y��Zy,̥�}ڐ�f�����Q�����m��Q���{�|[T�J�K�b��xK
�$�+{�����{�;��|>���ܐ��8��2����zgW��?�^ԹZ���f�#��l`̅xl�:L��j}SkU�^y��ٟ)q��6J�$����m��[ҷFOY*2��ub��z<���(r<S=�o��8*�t���83^w���+D���Q��[)�Np���o�r9���p����t���e���~�e��A�5�2��^���wr-^�{#�[����m���v�y�����l���8�ܷ��y�z)�gm;i���݀{)�vM����3c!���&�x���|��	ƞ(*ߕ��M��V�W�}�Ə^�0m����gH�^�N�or�<E}��h�"u�SW���]��5������m�ԯ}�w��6Q·�]�"�4}���z՛��&qL������z�׳�{բ!|khB�Cc�Ӛ��6��,Ysa��*���q��vi н��I���UƝ!5��|%a��i(>�{�W�t�_p��\�l�|����7Hc鋋�j���FU�gN̽�`�g��#�
R��YNPw�]H�q��:��tk�?�����UΒ��c��o�#\�>�f���:��N�^�)��އqj�ël{�Lzzw�� �=�l��>����gXP:tQ��$�{ӷ��U�}!9����>��7�q�s��z���l���tI����U�E}��ou���]�3�b)\�گG�{O��L3�͂���W�V�ؤ���q��_�s���{Ao;s�:tͩ+���V������
r��o�h׻.�?^�]8���}�g9��tB�����s�cg��>��т�ۖ�%{���W���w�v���j����+��wt���^�w'at�C��-GdM{���FR�:�?e�̞\$#x��k<ќ���b���X�PwO�����No`A�s_�->��d{�<b�G<+�*�8\�zpF}^����6�{��3��ΗW;o ˰JN����[	Gt8H�6�{)����÷igS8�-k��K��D��%��+���n�M�e���Y<�v�W�Gn��R����V�gh��nm�8\�usi�ayiu�3�X!��c��\���.O�������ұ���Z����+y���8�>���^����Pc#j�&�y�|�[8_�r����Gfl{�ޮ������x{rp!�n(Ы�e�����1��-�����R��{2�M�>xz�־�40���ޖު�U���+j���^�y�>H�os�j���J���j�r1�7� bߤd��	�����Ƥ�Q�	���M�eӮ�^�޽�x�,�'�?��c�ѣ�uh�S�o8Fm����逸�=mɍ���:%*U�M�R�=nq�gB䰔�*W_˛7����g|.MQ�_1�2�=s+�z���wU��ONO����:(�v:����G������4��.��}���ݪ�ϻ�5�o*���}��S�|\ϋ~U�u[���I�3�צ玽��ف�{y3�����8x���:x\/ē�z�fP>��/l�8F�@P5�R���gySO�n��n����mؓHj�'���w�!0r�v�v1ǆ��fl[����Ӝqa�������S9������O�P�x����>��	:u*�w|SÎHq�S�o����p�\��3������}_V��9���	�����)y����{�&ؕa��W�Κ>�L�c� �,uϮ���Nh�������ޗ%ǆWzB�I=%�vNן;W�65zQ�o�YpNx�ɼ�d�[�Y����h�9Lh����}��wP��PN�����v/-���g({�nza*�7�oDy�
��>���`����?u���İ��X~�ʿ#�8�;��qyE�4��ຳSՅ����\�����yS����B{(�:=+�����\I��s�#������̓��c7=�ݺ�n�����?!�{��1;s����U�3����店��v'��*3�����%y���Ke����^����N�t3�/\�R���I��,�^ͽ�|c�f�K�r���p�X^�kz�����ٿ��IӾjO1�.���ݼ�D
<:�د[��ڱ>kR0����{|�	�V2d{�Ӏl��S��=��0[���-��6�ػ'JX�4�4�Ȏj�ԖЩ�SB�r�R�p��<FV�s���osmZ�L�����)λ�/)�r~��}�kO=�6":���`��>>v����u:��7�����%�a��[�?Gϕ�ӝS�n����ه�G��}������G�uoE$�{&��|^��'sy��قG�,��D!��\#xN�y�xt���A��?��vf�]�,��оYS�8x�;�1��/{.�N�zp��{��U�^S�\|�L���U�k�{�p�;���$��v�	XO�=��G�ڏ�e|g��J>����^��y�����+��J�|��~��>5�����c�Z��g�]����*�k^P�#U��;���0��g^;�-���*�[Tiœ2������	Ȇ+0��^�f,
_{E߀}94�z���m��$/Ǡ�K~�7����]yb[�6o?>�SޙU�^��������T9�[�ރ����_a��}�Z�%���J�s��BssFj$P�7�r:5��ip�t�$5&�ɩ-��Y�R�$�\�.|�Lᓨ�}WL�hn��^)����he�Tn��'2f���N�LdY1��,Ck��'��m߇�$`��k���mׂO/���W�D�(�B���=-ɯ�����ϩ��7���gp孝�Ee��8雄�wD_<eһꅠද��.�밎�eჅ��p���.�N� ���1��9��8;��&�<)�{�ȭqK�]Let��Pu�tr�������:|�x�Pmt68Iے��:�[��^��Bk[�=��(J,��ª��7�^e6WX|�L�S����/���s�Y��G1J
<�í֭��/z�&�\�Sxje�9W]|��2O���qȞ�4D�w%=��+�)��w\4�Ց_;��f�P�Xh�m�g4#��h{�6뷱˹V��t�<�p��\O��gj����*�>�)���#�Mqҍ1`B�{ga�Y]��I_�h}���Î�V�GYm�o�SoBU�
�A�-G�.�N�M��O͙o�:�]K��6@�`Z���i�$Ag&��k�8:�u�{^gOj��H�9ڦpْ�Gi4Q���`�c��r��?C�9	�w�wd���ɬmW�xЪMҴ���]GT�9gf(Y�wJ|�X�,�s���k��0v��%������~]uqFۢ6�N���4���[B�Ny,ĳ4�3[D�uck���;�s;9�v[���[�jGlU���wYv�l�t4�[\�qP*}�+Y��y�;]��tqT�A�k�ݤ#���w��ew7�T��j��GR��Pr��&v�|�}md7�vM���ٶr��]�L��)�Ip��X�kv�FL�6�i4�v�����b'�5�m
�`�Z�wDn�R�U[^��HEj����{���3Ү��mX�0���%��ǝ���q�.�O;jSO<T��� @_	�vh[�� X�]J�#��@b��H����Plk$W������B�,��i��"U�LQ�r���3泼kk��v�qNa�����t�A)١�f�����d�9�j5��Ҽ�{�.A>
��L5s|����E!�X�R�r��Sc���8Q��
=�ѣxݹ�;r�ܼ�ި��pKת�0,n����"9���ݺ�8@�yr.�q8�튭��ge�<�a1��&t(\���Q�,�Ă�k��H�O	�?���R��;$iם�����mB7�+R����C����[+E�[� ��у��Pw�(�V�R���Y�rm�\�Fϓ�m,X2R���[�(�b��8 r�N�så�ut��!��IɗX{�k�i	B�Н��Pp��1�ҹ���f�\����H;�NEʲo���FzǵK�]f��9(��"��V(* �J�TQF"�PU���$X"�R#�AA��R#Ī�,QDQTSVD@D�TdGY`+R��*�AbȌ�+U�E��*�QY�(��EYf[ ���IX�((�AdUTX
)b�DAV
bU,X+��,�b��m
�`�*��*"�QA�c"1TTQZ�PV)R�b�,P�V*E� �� �"�b1Q�!�*�*��1b9h��DU���X

*&%TĶ�AdD[h,b��F"��6�[eU���`T10F�F
**&Z��"�1Ƥ�ATUAa��*�DX�b�cS2���Ab�
�(� P P��J�:-��^�U+:wGw;�:Ke�[�E�Y�	��m��Q�)��M��vO���kVj���yhGWJ����諭����U����"���j���^4竊���-w��.?c�>�����|-��ok���}nW��lg�d�+���t�������kټ�T��N��^L�|�[�-8M���:�)�W���p��店C ��Û�Z4Rƣ�}�Fg��>UG�EY����,.�B�/�C�3�f/f�\k)�B��K)�V��ǁ�=�o{pI�qY�:u��:K�鍍Q=�"s3��Գ���d�{�9���Γ`s{g�q�N�vw�:w�Y�L�<�y�w�N����Ԣ��S�߻�	�U�5�1��c^��HB�
�[�f��f
�8%�2+���eU�~]�9�d�R3b�+k��P��jm�3}t�����y���J����7o8��:tͯexM��A�1�����@7*���-�gI���nB���s�#�cg��>�Z?*-���*����lA�+���P%뮫�!��@�+�\��mʔ������G�4����Z�誻^�]%��D�!��\�'ݺ!Sگ�5���=n����k9�
v��A�E�7jA���T�-O�bn_e��ߪ�����U�nG۾V���N#�t�*M�3�����U�{C��/q>�e,HO[S��'Ko����!�M�2��phۥޕ��`�H�u���j{V@.��W{b5�:�-����ӾÍzC+	�.zVjm�<4��|��ץ}w�3��ۛ�s�I�d�ӂ3�7w��5^��z�j�r�7�+S4&�ZGپ�ߖ�+~��1�������s���Pnl�+����<�,.��˿������ײ��.�ö�Q=��VG���)���o$�N���.u�\$����M��������^��[v�_�G�&�����0��P�ʒ�I��ʁ]&��{6����p��-Ԗ(�$o{�g����i�si�$+�3%��q���]��t3�����4��|\yg��ܟy
_�����9�o�oԑ,���Q�s�jvI�T���L�wV�/!�W��]����^���Z\hpQ�O{���a4�ᗟ^��l<��a�����u�78V-�xz����]��XT�Vv��Jui��w�����y����5���zow��� yF��mĞ��Y�����J��sf���4�&����u��{7OW�C�%���[G}��k��������l���~�L��;g�+ӎg�SrL�q���A������J�t�O'f���"��F������=��<�����	<%�d!���n:z��z�ۙ��Ν�����;W�����n [�9+�*M�V��Κ9�;�pY��t��	��'����뿽�IQ�2��!�M�q�^��#���+���\><9o��+<�rXr��x#��Y����'Wu�`�"3�����Q��|ݷ3�f�F�{�5x�!	��u~���8�5���*񧷳�+x}�Q^/V��:<�x݄�6T�z��q�C�z^׼�^���/3f?��D�Q���Cqݠ�K[��H�.]dH[��ٵ�5�T�&R�ú+_$L�1xf:H`��q*]Wa�q���k��Bw+o�YǏ��.]֦�1q�RԥZ�\o��Q�U�WALTyiǢ��X�L����2��
g:�uG��\�7˧<�:8�٧ݲ���I-�)?O�������Dom'��:�g�~��籛�6��mB��.4��.{t��X>-:q���a��U�p���nXu/�#u��4��|l������?q�*�N9׺�l�n�����h�^s��{|n{����u�bmJZ�r3�(9U�43���:T���nڜ�K�������AYG�]��!~��S�飴���[]%��N�|ٰęGR�1���+�����s�`����<�]��a��Q�;Kz�JⅢ�Ud9Vw��K���<���t�es����jG��[��tQr��h��	M65L�f7�x�>�Es��Zx�|`�Y��p�H¾� �Wb��{�*�0�U%��b��W3�=�\/I��<�x��C~�^���]�������7��ܑ�+)�D{�Di'��<o�]� �X����9�)z?�%��d�<}u���k"{�r.����eC�YK�׵R쪱D����k,�{9�us�Ly�ZC{o8�L��S��Ի��b�-�}D�{�J�c�����yү�Τb�2���Ձ��eJ�X^��gD��������z��߾����ã�M�5�Q�}��?b�wI!��q���2�����A٥0C�<��w�|�/"�8����v��<�~G�}���lvA��Sţ�r%����~�>:u����S��GF�
V�!�$L��Գ���+ F�������f�دw��	�:���E���W�<�q��$�
��c9�՟t�t���8p�>���n(Bk�yr�_Y�w_�]a���0��-e�3���u�_8,ny�ig�k�q�Xow��l�t
؇NS/�!���X��J?Ki�0s�y�C����E�b_�˲=���P�'��m[�&���K��.ӽ>�[�W��b�^9Hئ��)�4/EB��-.%����u��sñ|�+���U�>�gú��J���J�r���0�$}Hb���B�����W��И39wM��b�Z����;��:�,Ob�9u�l�ۥG�Hy�� 0{�q�(׊�rF���!�z-Jǝ�	��6ST%���q�������pN��!����i�v0/X�<��y41M��%��x7�Id�0^S�ʡ��xXܳ�I�F�=�,�]��n�;��
C+��y;*���ݕ|��M��4����=�Ԝ:a��^IV�ϝwʔ���������yåʼ竵ԗAr����������r�i�_��K�����(q���N���ѰY��lP�8k�c��x
w;�;qz�WJO��#��şPL��Ϊ�j�}�(p���l��-M�{V�߫{t?g�yA�D�aݠhM-7��e�
f_�M)c�4����s4�z���{Ns�ݜ��z�x��ٜo��f��C�@��Z��K����*�5�b���f��ks�y�'1�ػ0v|]F��(oQ˗���H�d
7��-���i�o���^y	ޞv�l�z���=��Jȃ�2�
gþ�!�eم�H����f�~�ns�{!�����n�2�xc����IXr�9���$��䖎��w
��ܤ���wbo9��V�}�H�����x_���P�ޖM���[�8��֤6�c�\��.�e�j���X�[��@�k(�T��b�(������Ə���a��Kao��W�� >�����'L�'۾��s[��gX���a��Y�"���uCF3�.c��=g�q�ܿ2���&�-	׋6��ٹ�v�L��K+bRNC�jv�ZsT2��/�Z���)��J�N���$V��,�p1���y�;=����L��[���@�$-ʶ��Z�.��wa;[%�:-b��C4�Wkk}#�f��������t��7�� |�,�HÀ��7߾�/m٨��Y�<���c�yCLO�c�^����U���N44x�����hX��ǚy�l����Z|��*��c�X'�x�i�/*�Ԗww�\��%�����:D�z([p>�b���N�C�Wb`D�;ޞ�Ԃ���OZ�90�~[2�oQ���y+7
�f`,��	>΢[)�Qw�N�3�峀z
�Q�9+�������w�×_�*Q8N��å"�t~lq�"G��ByMH��;������
t�o��h`v�~�i�ˮ���v��0Uqx�&t}N\�fT#+�Jk"஬�=*Y�}ݹ�Y�����.�}�֍����x	o)�(t��̼.X�ݹ�M�{��s�~P-��תX��;��,������0��D�$�#Oj��T�'wod�ލ�m6f�*z�%��p�hC�S_\�(l�z���y�~�ƣ���tR.��}��Z�_jTD>�4:�������ɓ��]����X��ڼܖ�N��y�/s$<�������Ӈ�q�Cܓy�p.B6���V�W�\�VdƕД4G$�=�YF:�ww��q�Rt1�٭H�F��3E�\��C�(i����'np-rwH6��(Yݸ�X.3��9l�u>�g�-����c	�_ow� ��|�\ҷV��I(�/�WVP�
�D��j,87��W�P��Si���V	�}o���ן~���ґ<�/�.��a��LWR��*����A[�v�x?���
���:�������߳�ɩ��<�$�t�XoP����7�)��������]\y�v#�2G���=ˠL�o�G{=Џ:����[�^�n�j�2R�}�v�>��Y�;�S��!>λ}km1ۖ6,.��{-��M�g�j<�px:�ma�[��G�u���.������q��ִ�۰��s0j�{� k�����v�<��c�a�G�W}��[���8T�{K�"�q��[L��ܼ9S���q*�o�Jr�8˽������/5s��+-b�4�j���S;�0k�q#�i?S!�������[�jN��&u/T<�g����VZ�-i�͑Ԛ(l��L���#��vrho�{��qy6b.��cL8��|��Lt����v�6��iq�H�k����D�K�CR<ow)%�cL� ������ʳ���%S+f���q��
��� �~��ǄH�6" ���{�����9��]�&�e�J��PW��N��H� ��Q��z�I�9�2�lZrm����s�0�}�</�������5�o�fa��^�zg%�Vf��L7�Nx(��[ޯ	2���Y�,�4�ȏz�s,��M�]�꽒$��� ��C�l�LPN�1�Xg=D*��n�u��M���rN[��د�c�S�s��$ԢVT1�"������u�z�_��p�S�2��w+�Su��ü]���m�X�)%t�x.���]^�Rؼ\Z�}S.\��0��&5q�}���m���)���P�A	疒5���N�˪���¥�8�M�yrK~�w(�sOf����L�.��pHi�9(C�"!��	��N��kc��2�<�'��NL�1p��շ��wW��0R���jȔ�;􆞥�����,�6��ў���/�Y�a{Ӆ��[�;�3O���B(��rXAb�9�bgV�N��ۇ�Y!�++5����E �hC�B�^�f�m�3�o�q@|9�o���������o/��v^�e�3�M��j�����oD���������c�독��m��"=u�9˲4X����3�.	ƦU�5��T��6]'o����R����C�Av�_&�*�x�e�YI�� xf���k��*��:S���cMx�S}x�T8}��0?Uk��E'�w,ă��J�t��_Y7�ڭ���xqMB��j�\�F̩J.��ྼ�cj��LC��7ۻ�ﾯ���Ү��q�:q�_�s�d��A혎�Z�Ŕ��,�/�Ռ�VX>:\I�%OOn�A��:0\ݚy����u�a�v��l��[�������m������t9]�ك�鉰s�)vh^`Ͻ��k+K2���R������{�WH��q�3*�ԂlU]�oR�����=n��$4�+�3�K1D�h���f'/��h{�w��>��i��ߵЁ��k�X3�>/u,F��g�U���
�l�,�SW��Qd}tx|��i�E4Vꬮ���W����ddv����xY\dX(&e�we���?!�<�6��{׆��^������Ź��8F��T#���w�yLD��u2�L��)�/�4�O-�q��8�Tg ��G����������ޟc��o�O[ş��%]jWK���3ו��ޮ�ζ�i3��8���^�B�c_�����b�5�{���9 �>G��p�x�˙H��,V
�:�X틥 �5���fo<lIY~]�^�՝%v�˳?F}��G�R�,-��r���u��B��KF���D��6��o7b��6����R�S���
u�0�r}RJ��_
[ٷ)I��ŕn��aJ}چ[�>�yh���}��tb����M�d}ˤ�t��}�=��7���R�u������Lp�x�����#�$����Q��*tt��7���N�3�5F�����ɍ��]�gpR�	.��D-m��.��������?�iǗ`8s�z&�HVn�ǌ>�O׉�;;��G���}/p-Bk�C���@[������2�ޞ���ZJt�;���D#"��𘀅k}Ea5r�uK�}c-��/6�ʸ�V&��<�X=�Iek��Tg2��<L�h|n�mtVnv-Kق��O�j/�+{ٌ+�{�����#v{�<�Wt��,K���Ɯ�#kd�&1A��� ���M���#H;�#6��w�p��0���&�Q�u�o>�76��;9FӴ.,T���6�i\��h��`C�!�f��vhZ�#k�0����Ӫ2{}m8��u#��-�����eLzS�Rz�D���j6:��J�1oѧ��.�[xS��ƹ���!��˝��+����1�I�z�󼷹�Q�Uu%d&�B��"�.������'�}�*٩��F@���.�p[�&Nd��w�%����k�����Ք8cv
��0�&��;�nK��̢�����%���rr�������+]�Q��X(JEP����R[�@��#JŅlZ]�f��P&wD��VHQr�r{��fR��j�M�
!g�����>�ɵ�����uї��V)G�J�����r!qv�A��ٮ����J��s<1J�Z+�m띆�ww��	k������@�ch�D.6���`��	f���iiJ4@39�I�X�q�*#N�S�,C��� i]�B�giS��0k�y[�|�6���5��mfF��̽�o�6�vJҨ���󵑁e�Xf���%cN�sW;�Z;�y�V�{����v�Q�Z}|�;v�E-tR�-iD+~�C���.Կ���u�x��A�n���Q���R�f]����7����s�:��t�� �5u�k�Q���^�L��
Y����//O��Z*gy�0���b�t�m�۾�[��	�Iw��QՃn�cЧ[$�c�Mbr�;5�Щ������%+#cB��b�:�'$CNqns�C�}��\G|���M�$�f��vktv�{г*���m�l���;h	��'� r�M֑������c�2�{�.�Lvčbu®
��}ܠ�|tP����J6������;8��-hO��δ�F��BG%�Ы�gJ��(W�8��=+"��S�}��'.m��6�J��N7g ���cY�f�YN=�yY�j^�wІ^v�-.j�3oV��b���R��s�y���j��wݜ��э��a;i�p~z�>�|HI@$�'�GV"	����E��YmQc��TPH��U@Uq%QKB�,q��ȤPX"�Q�YH�(���f5UH�DTYZ[(*墨�,Eb��2(*�1Q-�����*�E
�H�,Tm��AE�ŎZ�G
���
*�EPD��e�AAA �[9jcPc�R"*�E�E%�c�ư�b̶֕E�c���lF
1F2�Qb�`�)m"��b*�2�#�c�b�ZcD��b��R)P�m�-Z�X��L3kc��h�-X+���m��DX)im�T�[�D\n\ʦR���K������W.�10s(��.XTEb���dDb�L�s,G�eJ�(�̹��ms0bdF�����V���f8�3)��V?MQA���S%cx�䎄)���
5�'�}����\h��A>�V�h���Ws�O��M!�4��s`��}��6��{�� ��^��=0�$^/�Xg]`�e��|Z�3�邒��B*�s1��RkF	-?=kݥ��<ޥ�Rǫ-9+�
��5�^^�c�c>9�.���X�X`���m���z1�;:'�o#��do���>���4�*�>LpT�zYx�z��'�:�̠�����
������đ|�oJ��3kƚЇ���9�f���[�"�dҪ0��dS�T�=��ѱY���x@�������v�v�������i_w^�Y��w<k�&9k�z%��T����O8��{� �z�y1�n[3>ws�5Փe�7���uO��E�7y�����br����
������\��)OɈ��{��!^''U\�ن��uΓ�Lϟ�ge%��-)���{K�5���(��'P�\������4��_��с��|�HQ-Kb\��W��v^S�86
�&�0����7w��=�A?Q�s}'+��:�*m	�9gOĖ���lQ���N�9N\�_oN�^�>;$ý��.N:��=c�LB��q�3�$���K{+r�ӱɑV�
�T)K�Y��岸��*�7�H��F���LUr��2�V^S뙑�Ō�n�d��Nb�T���M������㜦=V���z�&!W��)l�
;�)�6J�������U�w��u����ǴO~�&�5g�{�x��ힴ{�@�,��K��(P����{��/�o��Ӝ4j|0K�b����u�C�s���>�����z��1�4Mt�$y�OⳲUV\]�D������C��;��c�]^!�]@�{<C;���Ͻ��׫��Kh��1>�r�������GR�C;@d6��kV`���TɁ�˱�	)Z�;jp��ױ�4Ow�������ðW]%o�f/-�\5�b�}z��79�$�0�}�z}i�r]���\�U~��]*�N`@�4��� K.���������w���n�*a/1������*��j��h���$߹o�ק�lٮ����\�\�9�S�"l��;7�t��
�<�"�Z}P:�<G"�z�}�����p�����'^���h�Ѿ��t��Z}Xu���A�v!Ͻ���ۡ��=��ɻl�(t����5s���J)�ݻ��C����D�a.�/;d���� ͻ'R�{T��s���R�<t蕸��Z-A��f�<��E�����,���y�c��ʝ�Cس!��Y�}I�9`R9Ϭ)N�R c0����<��7.��ɸ��Zt�S�[�"}fZ8w��[��y�#�l:;_\!��{�/�n�z W����.����?}_}�WƤF8y׮�1P~�e��X�O������D��鄜m�3�x%�ʷ೔��ყ�ej�v�H��n�~֋+ჰm+O�L���	Ď��*D���� ��6��yy���I�<'�� �L̬��Z�A��'�T6`���ݕ�؎v��V3�d���H/�&����\�%�0�s��߇AZ�|:z�x%�,�\k���Px�iR���Ɵ��������Ɩ�,�w�0�ld炌��� \zt�"�K4I����~N��~��+X�q��COX]H;��1A8;WO�9�!}K�;7i���*���ec�ž���>ۤIK�I�֊	�@_��X�C�^����E~XR2Z(z�xp��-��^y�B�ܭŝ~#�@�}Α�S�]�C���k�l\\Z���_�	�O���7z�x������BZ�r�B.X�-夅ഖ�h�߆�xk�)��j�KQ�����=ioT�E�S/>�mrz�Bl�"	�/�w��|���ܯnf�oW�M:uu�����y��f*U{�����T��oz���:�$��̏�p�*̹ۧr] 7:uso7sK�y}
�ʸ�X�\��%��[�J���r
��h�,�಑Oo>Pf�,�sR�S5�&�iu9�{��諭�e�3߽���n������K�iɂ�ۍY����Q>j�lGxF+{���k����<4�ߪ}Kj�2��uqy��;zX��*��0D�ϖ��t��ƌa����^;�����药=U�`�f�n��^��u�[�,k�m/R�ף�=d�QL�3�X������{,�X�W_ڪ��^3�L��]xȌ��nbm����_O��#��p��d���ܰL�ӀjԮ,�����xg
��vx$��{̜�t}�m���a�t���.wU��Ֆ�����[h#tB&�I~����x��H�+�i��D��;�8=¸���T�����u������Q���t-���-[��w�ꮎ$�n�*E�+�k��_���h��NP�	�懄�C݀N��f���f�#����Sǖȓ��1:Q �.,U�`��:�����YȦ��Es��ϋ;�!�YS�����9��fx�:<,�������+:G������	�c�x)�~Cynmh0鿾�����M�v��*��;)=�I�%���J�^�o,H���^qW>asj^>t��ܶ<ϥ�|�̜OnJ��E���a�Fo��%\�{̌�J܃��5W�z���[}2�TZ�ˬ�ќ1���fL��m�9a���V
n�1�+[��p���O��}����IѬ^��n����ZxS��&�v���4�ɗ�P�e�4��v�Ҕ��������{����{OS�����u�M�w��z�,�/%��-�XKGx�T�k�r�>MWRٲ�m�yi(`�;�C��������b�$U�w��ᒗ��Y�����{=k�&d�!9y������sQ�&o� �+"�˷��CVtb��2��ﾩ��j)��������t2)
B�e�G���mSˀ��M���T�ug�00��:��!3�ok���;HY�|��@#ΦP/������Ԙ��U��J��D�����̀�m����N����<������@�US�1��﯈y̻LV�U.&8*v�����=S��L�n�����wvW�p�.O_��uܳ�α3}k�kڳ*X�x��p�6'cZ�iTZ2H���5I�c�<0n[3>u۳�?q~�{M���p�;?7y���΋��b�Ԧ3���awk>Pe�W���x�P`ܶf;��K0�&&���_o��c�¹y�j��64������=��F�X��ޥ�����pv(�Eue�Ч�;�G=����܀�@��Yri׹�Ή����X#��]&kbm8��r�+b��5m�[��d=�4���nu��/�J�6�w`��wt1�r�?Y�^ow����ֽ*G�/�w��W�LP�W�P�0}�E��;��n�d>��z(a�y�ξ��f�q�����w�ILWy0�~�Y薛k*���rɾ
o�-��J ��w�Q���U�Vw{]�_������rȱ����KR֗*/iW_���N�H��Byi�d���uX�v������~��
�:��*rχOƂM-�����V��s<��+��~z�O>���1G��>ۿi�3�����s�j��Z=�v�#A��53����<���}~�bW&��=}i��.j�
z��e��~��}=-�d�f��L.�'�㭇:qC>��P>��1kkȓ>#��B��c8ЖWՋ��w����]����s�29Ά)����;�������e�B�#���V��v�Ca�m�Y�A�
�01*���5G�s�o��$%+�J� !W�4�����ZI`�H�,�quL��>�g��Lm�s� ��]�ٱY����>�Q|p��l��dK�˰�i&xCk�E�\V����;�n�[�xr��f)�Mˀw`h����Ś�y�m4�"�$�
�o��MT��
LA��O�9�Z��{nھ��e)'T�o9�WH�^�@�wa��S�����s��Q���j�+3��:�'�"�Y���(�\!�Ju>7���?}��WެNK�!T��w/�6�	��ЍbCL�q�>��U��w�y�n-�C=m7�^C����fv�/!u�{+ا�踫}p/c�{�^��,���SV�N�e��c��y��/��Vc�-0V�{��idu*gi���l=���7m���#h�O���?[����7��h��1�����&x�d}���q`vX��4ȚW�n��Z���R�-�e��o���6\_Q��*�6Z��+�R债��Oi{��/�v�u��ڈR����ű��)�q��;7i�@a�=W%ue�VF�\]#l�R砺��*{K�H�91�e���mw�a��b�҃z���'��6��ˌ���Yk����6GRh��Bu�>�u�\�v��r23CC,�_R����Fd��	���z
ְt���]��3`���ÇZ��_�	�`��	�wb`���K5afo��&��k{+����؋7�������)�\���0wR��\Y �/�u �K~E���֮����,�ZOJ�u�dg'�W��]],؎'�I��������I�V��X&�)}��Z�N��	���B�W�u_���@#����;,�I;z{o�iu~��mF+U¹K�fHu�W���{&!��7ܩ��V�F�Of��pW��V�:-�i�Zo=���}�7՞������n��?�K�9K�����`�����q鵁:�ܽ�<�1]I;|����sу�p�����\sس�~�@��#�&�w������^��Qޮ��itrr}�AC����:�}�P���B,K%�������Lw��t=��3��]��o_�ͷ����]��F0�(^}*�&����pJ�ʢ!��Мb��C1�}s����xZ��|J��X`Q���6�[܍Y�-0d)�.�O��E����"�=�v{8�zɝ�~�����	jZ��U���b���c�,W��13�:�s�bF��Jɶ��9yZC�{P��	�..��z��C����}���[�������9��'��'0����0* ����;Mj8rb�J��?����Wx�o�z0��ҝ&]?s�����dn}�m�2l�ܴ	��Y�ק�J�GH� �T.�YR-%-v.9�\�	��E�<����f`w3����`�.wV���ܬ�p�l��>�q�Xyi�!pr�F^��y:thH��q��*�V����t��P��.x��2-f���5���s�B*Yjm́���+`+���r�k7�SZ��3a���MR3��%8�ƴ�|����j�:.r�x^Ͳ��k^|�H��No��c19����������Ps���iCW�8�1���Kǌꧩ��c� ����p무YĬT1��tP�#zw`�Hs��.U�S �A��C�����1E�M�a��(p��BqC4q�~�[��W���%{��N�+ơ���#`�2,�����뮶���g"��%�#�-��c���ο��ç�w.��Ԍ(�9�� ����켧a�O-ͨ��z/���P�Q�zjY���<n��Yi���l�D�H�Z��^P�f&��v&N�3���z{�̙to��F)���u�M�w����x�E�D���V�����_f���K<My��ӭO�h��䡼���rƿ)��������ȯQ�P�K�Y$�[V�?ez��=X���l#~:���i^��G�炌����z�!�:3�:��7�tw��1�[�ό�H���X�ˬ��}����R��ޘ)+r�a��.���Bה�u�Z�?{^_��0*�Ը���o�Ba�}�
����&;1V3�3|�#8N&)7�S���4fԗ�M5!����>����F'�E�p]��K�.�޷�~�o�m���J�/�z�B`�L����Lu֓���k�(v|k�ާ$�����@�جHΎ�"�q�4�o�h�U�K��bC`���M�2�#�L���}?����}n��b�gp�_۶7�:�Z�iyv��8�>���4�*�)1�S��xS9���>�[Ɵ������܌��a��i��������d��6�j�Ї��L�K{w=~��qVڿw���)�K��p�����^î�5����7TkN�{�i��j����ډˍ���Ǵ���ற�"���><v(3r٘�ŧ�5Փe�7�/N���Wk��jj�[����`Li8�b\0���*W9����s2�oS��e�n�zet�J���TF����q�������Ih�����{K�SP���C�eV'�H�;||	����(dvޭa��E��Uʾ	jZ�-Lt��Z:|���K��H����:? p���{����ґ��
ϥ�>�9`��a�TGZZ%�L�N�z�u��|���_��\0K�/�	�{eɹ�Y��<��(]���G�ݠE��k�����5_�4����C]�R�)���ʇ��#��e�=-�g��	������W^�*�1����9�;���Ps��Gz�.|�'��j��v�{�/���	�=����5�krk�C^��D�`~v���O�/:��'���ҦE�S:���!)PY�����Nr׼ �Σɏ	��wn^�L�-Qc�1���=ڲ�{[Vde�5���y��f���4-��i�����B�1���]Ja�6��(�4l2B"J6&w��x�������˸��"j�pj�^p�8-�9#�	����>�3���3������o6���j��J��h�J,��9�7��p5��ؗ1ٰ?nl�j��V��0u�5�W\hjnzj���z�cI�YBOs�%,�p^��yp[z<*�iY���nIҵ���њ	T��>yh.��G����w1�{\]mQ�l�w\��E��p �;���,���W��!A�����[�x�
n:�u�Ļ�P����7�Y�>�R�e�W Y�腋}'%�u+6�ݮ&__	���#���
�m�[4%�u<��5iL��X��2=�3�9�k�ȍ���Z/�݀E��ʕ`�I��Ĝ۩R��=��"m���2�T��~i�!9�m�Ǧr撈�׼��I�Cz	2#,� u���G���(e��:����T䰺yǁ�]�I��7��r���-��r���ˮf(��Q,N�s�o\SjG�V6q{<3s�L�ܷۋL�0Hݓ^ٯ�ڄ��a�л�iX=,N���)
0>��+<d�h�5����W��n�Oiy�Ed�S�aT�{ӬY1����4��9	n�s���=��sJ�J.o�J��Ϩ3��D�:e���u1��R�VN��칛�ޞ��^�2��&u�/�qIp&���.5���u�΅�wt�^.ɃT���]��-�C.�s+3���ش!�+����R�_���樌p���g�b�Y}�Z'�����:���:����X��� 뾧��C����B]�^8�����n��K�� ت"�>��H�`��*5���O��{e�G���Eqx`�:�q��pg@�1�(�)����R�7��ڻj:œk2;[cr�t�i��xN�K]�oj�,Z����b�+U�e�u�(����1H���W i�(�qk�خB8"T���\�%��9e�G�vy����|,:7zc'��r�1V�ݨ���^��A�7t�SiŇS�|:��/Q������伊Z,hL�hu1[�e�T:�.u�{4�-��2*�5gf	���xۜ��ǝ���j�L�C'�5�����=T��Sn�*�ݝ�SIqތ�L�j���"\q_�R���G���r�4Cx�ћ�7�c+���ahZ�j|i���J�i�R��i-�/Um���xRd�nϬ�f2�]��)���y����� �0�;��N�+�+��xcJZ�Qk��M�`�}/�'awo	�^r8cC�:�Ƹ6�z��׍��� ����5����E���6���s3
�`��EƊ�SE2ܷ+��J`������!TL���c��+Q�X�f�h�U����1�+r��X���eH���F
�*V)�������kiV�,�U\Je�TC3%�*��1��E#�Qna�ebe����,�QJ�#\f(9T̢����*+n8�9�)T������"+Z�jEQ��V��mh[�	���bJ���Uư�Ĭٌ*�����l�Ɗc�0UY2�3�j\E��1Lˀ���1�̘�q�0\�m��YF��
���dX-��j
9km
�-T��E��\��h��%`�-�8�(��2�*am�-"�m(T؈V�+1�q�-�\���LH�dQj��q��TEDDb�FՈʕ�Ve�k-(b��R���,E)���ˉXc�$el�e*�RѢ̭���[`�B�("~H 	$
vs)s��׾oX�9��}>�rhv��и�n�T/-�)c�ҭεt����'cܷ�m嗖rD��Tz�:����꯾���)�d� �"M!��B��8������҅EW�Z����!�~�S�<�8�����V��9Abӥ���)�K���GR�C;��~͵�3�ˀ{}��%��/�O=ˤ�PFiߤ��Vs�9g�C`L��D�Ģ�+���G�jh�٠#[<�o1�D�I�V��V�{�`ȑ�K��]���I3*�B��KMn�]Y��+5�4������n��x�wWb��tU��a5aЍbB� ��tN�6ٳ]6�YA)���\��P�.�M�p�E
�=Kqh����\���p��},���q_��s��\[�t��>��X�yW�۰�{+q1�cb�e��n�=ݕm���z�d>~���E�w�A\�En1 ,k��u+*�ِ}�\DT]�7z�t��6�z֩�r��s2�OLX3LaY��D�z�`.s��;�	1�7���z�h�n�=�{��mX�λ�|a�=W%wՖ�}�&�(��mS4d��뙝�peM��rp�uK%{~�t|FM�*i�δ䭺�Vp�ܹΗH�]���>8[3�/[����3�t��v-e�Z�$���-\�Ytݚ�[2G��,{�t�Gx��o���ӕ�̔��*P�ʉ�4��]���.��}_ULt�����g����X&�"�u;�U&��kڰ�L̬��(3�:���ɫv�ATT��ҰĄ�s[�}��J��C7�N�e䱦Nv>Z:
ֳ����QgAS޵�ƧA}r5����!�F��wc�;iv�,���&��Ʋώ8�W�Y����^��;-'�
[�s����QDϤ���\a��C�!��C�LPN�]���].���J��R���kx�[�d�~��a�t���.J��f4�dz��v�X�}ʲ����{;&�ޅ��{��y�r�Y���breLY/��σ��hs�y$�.�]�����םң��l菷�*�j�bֲ�\/�]���%���JF��B����u�Z�;4��bn�yy)�0�QL5�+�lR�e�_*�'>���rP�nU�P���K�y���o_�cs�
^��|.��_�"���3>�+�F�ᖘ7!��`�d�X���	��t�^�G� �N#"#C�����}����"WOV�o˼z��f�oW�b3�A��a���v,
���2�N�����M"��:YLA N?>��<LR�yK�5���1*�$�굇�:�c�u�y��;�ÐӢ�':����:�������OlGEh2�@�C���}ٴ�YYư_5�e*���`T��W��o��K��jίû	ӷ��A�0�G��g�0�u��}~Tֲ=W8;��)���Dֵ��lu)�f��g@�� ��q�L���J?Ki�V=.>����4(���6�uzL��V{[������˲5�FP�n�T���:��Ԫ.��F����(l�^�_I��OPcըU�<��Kn���þ,=C�s��%C��e���5qn��A�Q�o<�$��(r�B�u�s�)���g;�� �X��5���=�]<+yۥ����a#��䱞����:��W�F(�n#3�<��hR�f���ʯ�a��W3�E��y�-X\GHt�x�Ih����:���YȦ�	Ԣ��K6q�H����w,��=YF�E�=�"Ƽ6;��i�<,���,���N�� �W
{�`ݱ�srwUd����P�M}s{<o�c�׭xD��D�*�894�]L�)�l8�߽^l�=�@wҿ|&��߅9�D�V|nK�7��X"�"\�A�����ֱo��5z9�/{�60<թ���H�N�ye�� ��2>��� >x>-�����M]��`FJX�t�`ʵ�.Ɲ�];�tPH+���1燐k�E�7W��f�m���ۯNsJ����}����;���=����^���HRx���
f_�\�61��C9c_���=�u1i�^��\�w*f�6�����k����i�8?���LM!a�a���<_J���IY~2����ͩ�=V�������g��r����4�du�Y�u�Z��;�՛�H���YJ�S��Z��u^I���x�\� r��s.�x�)ȑd3���3f�ﶆڅ��!���B�:|sޓ���.��{�����^kR����ܻ��yL�'څ�ʥ�8����W��w�y�������#��4��V��$X����}w,�6�i�z��ͦ��}�W�i�OuI�xǌ�~V;k����0{�����6t�c�f����:��{�i�{���ylY�ŷoMY�WE�)��yb|*�><v(6����Z|��*UHY^��|�V�F������l,�c�%��K�	sԩ=�]A�C�X����fB���UY~�	/��.]���Aɘw�'�B7 �7��m+O),����J~`*{K�5�
�*�QV�F������4��r����]pzQ��E�ԗw����lEJ�m�a�PikZ˫�,��\����+,(�ڤ�;X��i���4O�Bw*
�DN�m�8mr8� Ru��0��^b�P�O
��5s��n_e�� >�x`����)mbh{·~�z�6
�E��@򠖥�.TZ+�b��e��-��X%���w�Bk{v�F�C���g|2N�7��T���*#�$��m-�/t��!�{Փ+���?Wq�.��T�<�ʄd�e�2m�V\�<����g��v���n��$����b���bN.ϨP޿�_Zg>��pC���w�ƺ���^^1U^F^�SQF��ʉ`M���;�����z�@��R$�#��Pq^q����ut2O�iB�����=t)��=G8S����=U����;8�ub���H�J\���GR��gk!��6֬��qf/K�fS�U�͔��^xl�����t�xd�',C-$�$^.�\E]S=aY�P�˿?:)=������8���-\{��(�0�2�"D`;%/+yv}޴�<ġ�-㮚p�}Z���;:��$nxT�r��z�,ޗEX}0���F���4�=9�b`�Z���y6�O�]�NY�1��J��/"�TZ=��P�ZW��oc�r/�t�E�hGَ��`�#�)����Z�>���Y�|��幔�]��y�~�������k"�Y��G��;�At����ʩ̐t�c���� �}���F�k\����o����³�q"o�ݫh�4�ggD���p�s�jTEKN�z/����|؋�m�r��X��|}u�0@��5�¶�ݮ�H�#�U3��gýGg����=�+����u���}��c;�K���N��_�^��TΥc%Cx��9��qc�+�<��6s��GnwpU<_=�Sҡ�;UׯF�*!K����e.X��|*Dz�ŧ0dZ����m�{Ϭ�&u�/�����0Ȟ����ҵ��MO�"=�VB�fzot ��������@����X&�"�N�<�I�',������'����������藣'��t�b�A�x��V=��F�W��^s�P}W�'v217�$0�O���mII��a.!���X.�ϫ�4�j��ݖL,d炎L�k%*Ǌ��Uj��Ħ�+��������a�Q>��\�<a�qw��A�t<���1-]7�����n,]-�;��e���>sU�) |��]S1�"���.=6��`3�cޚ��Z~��R�/�'j��S���1d�>~�t�%b�B��<�(������IT�)s[8����3,��lih�|. =ף�r�ܰ������m�:4��5�x)�W�W��:�\6W<�ete�u�\���U���*-m�`yT1�T�w*ڻX-��ތ��<&��%���V�ĺ����I�J���C'$�=��kW������}�v>�~�Y�A;���.���Zʙp�|e�;�BZ�r�B.X�-夅}��%�ȧ'6�_��ҏ�V]Ϯ���Vj�-��tf)��ʶ��!���!�H�v��a�<6_���8�g�)���-�7�J;s��৿f��l=�՜2�B������g��4o��Xń,:�!�<C�:G�Y�;)���-kml��?�Ab��׽ƪe�)�Q����"5t�KBM�W�p���u^�C���7�d��P�;X��z�ɶ�;��X����I[L���y���>�0�i���Mc�]��&+��2м����Z�	pԎJ���i���m}�zf.��{q�0M�;����Y3�N}�R����q:c)_����=BG�tG�Zz�nU���`ܶfs0�J�0&˝տd�u]#w��~O��TPA��T��������Z����K���e�+K1�NP�2�������"9ϙ�\�I����R�>��ф�\f���0R��]1C��D�yъ)��,�L��z���S�J4 7��^��ovt�VPg���n�n��$d�� ����}̮�1�4g�����1Z��I�1�3���t��*�0��a��Ŏ��8G�Z�Z��%�YrDGvʿ�kv9��e�ij���qt}.*r���g�ǔ\�/���'��Ҩg>����o��﹚�ٌ��x�6��#`��Y�Uq��_d���χ�
��!���i��{
vדS��D3����?����ZG6��>Txy�lr��^�՞���f����;�՗ݵ�xз��7n�Yi�v��H�%��&��k����e��}=��3x,[�p/}��y�p'���~�3���Ϗ�3��	�x��D�(D��s����ѕz%�Nb�����v
^SJ cw\�s�5��/���;U~��/=���qw�Gm���Q��+�^�fd�ZR2.���>W�4��R՘7�
2+�>�v�u�Ċ~���y�A�F�xu���i#���C�l-�<Gn�G���$��n\U�J�_:y���7s89�kF%���]ß?R�:�h���~~�Lpv����?2���wx��ǹq��t���X�(0dY��1-W�������G�KT�Fn����j�fԳ�pϯk�q��o">�e��	���H����+�G]�;:����(k���ꮥ�3%�Y�y�=��CN����s�y}�}ti RWA���p̡V�+�`�rx�|G@ր#J�Kȳv�x���R�Vu`ޢ�z�f,"]	w�ˤ�d�l�$�.k�qྪѻ��]s0ұ�l��NhR�[��ZX�8&�,�~��Z���"��u�ò��u�8�<G&����m:~�O���T��P��y�����2��.
����@���l �ؠ��fc������;8�l�槍?bW��+��[u=�]�y�;�l՗�Um��UC�X
��P`�΢�>�!��x1��O՜�����W�;���Pý�=���Y��J�ʭ6�UWR���I�ٞ54ze��n3��u�����Barޯl=�X�tJ��0��t����KG��ݙ�km���9G���G�x��.��+�����5wO�8��Z
ۮ=ӪVVw��m$�y9J��ӵ
r��=p�{e�,d���	�y�K��h����:]1����ъ��\"C�S �C�����n��=p�Х�"���Y���ߖ
�t�kFϛ��+���|�Ϣ�"a���49�$�#����.a�{3��*�5?���}�l�i1w���Kj����z8���	^wO�W�"�%��
�_¸b��b8Z�KUF�_d�<�̺,�N-�-+.�׃��G	��
�������n�����*�<6rS>K`U�������\MY��g[�P��v�K�g$P��CeH��۶�9����B��9b����<WŭԘ2�0򻶘� �h��rn��B^���N�%]u����Ƀ�wc�>������L̤��":���K).ec�\����l(�;�k6�S^��k��wI[P��v��)�nJ^N����I3c��T��	��#�)^�>�9G\cMZ�e3�ڦ,�z]`>�MXt#D܆�'�'a^0%�絣L���? h[�T��엑͡mz�Z�E�[�ѷ��8"�z�ǬV�rX�C�uՏ�+�u�m�u��Uᒒ�~�nxӢ�k��8��T���?_z��p��b0�qp/��?�M�%>�l�&t��Za�g��D�U�S:�E�}��ܮ"WGG�5����W�g8(��g�k�pp^�[bW)��n��nq�W�v2�c�Q{V:�v���ޗL�62k��)���d�n����<��x�"zo��:ȣ0�X)qh�>Y���	���{����7�O�\}lW4�|<�H�	��S�O|�I�=��^Նbf`���*�i�畇�l���!җ�*`�����KP�I،��4Á9��h�R�+��9�ǂ��}^+(L���q:��ݷ�#X2X�,�Ѩ�F�k��E�B�7�=��r��Qu���U�����i�T�L��\�^û�����c�q��ԅ����:/U��uqK��z-�YF���,[0;��'�_m�\���8n#�F�x��+���:�aW��Z�A�:ả�kmGG2��q"�L�Y��c�����,��\�����.��<Q�A��^�:�ƱP$V%>c�o3���_@i�L��؏WDiAvJ:�,��q��o&��>�tC@�C�Y�>Ui#�P5�aZ�64br��V�b;�95˃/�t�=��je,��n����eԺ1J7�9
;������c�|�Z��p}	#+IsF�Ck�vb��eA�V7��S�����)m4*vA!���K��x����hf��pgi�YQ��i��be�<`�[�le����yQF��]�%nX���V�3���Y"�1������`�C⏴�Aα�.7�ĮѺ��8 �
���ٴ������ �,Z���xd!��V���qcz\Ғ��%l�,P�M��Vw�:m������:'��%���n��s�tKgl��0�X�%oV(��WwY�lP�B�W]+���l9��q'���l���&�C��hWb�f��'����r��o> o��t!��+��+���sب��ђ��I�j��θ��+���\#��e�L��]�q$���~9�#��z�v�l.�O���9&:��U��N��i,�0�X�覦���I۬�/��g��Y%��U�����|2.�5��vc�:p�%u�WB�aK$�w
�Vӑ!S�/4P��O����Ԡ*&�U�4�-���C[�`�ymĶ�-��i�/W�Ƴ'4�p�m�	�h��nlU�t����a�4=q���ݙ[�xC�b�
��ł���gb�7��!0la}Ċ��[���n�W�@�U)K���v��:+F�o�U�"m$�tQk���i�2`bv�P�f�X1z,�*�]f��n�T�nȭ����֣5��#xcWxd7�
ݽOh������W+��'pv+�ʋ�p�6ya}�2���9/c��>��Sy�MYE�3��rz�==�N�:V>]�j���u�{��}�ci�g�R�:�.=�z��V,x:e���C�v�t<>���e�ӂ�-�!�w G��B���n_V	ne�\u��,�t�ƪȷ�>�K�<�T̒���p�ʭ3��X��X�����~~.[ێĻ8��Cf�B���aH�f#��?��0Ðl���2F����֪O�Y@�;T>�D��Z�Q�y�WO)���,�̝�����e6�����V�-�C��v"�'X:�P�t�*���lͼU��voU�dɓS/�
+e�BRȫkʩlcB���FV��i+��1�3�cR��Q*�LE�,+�����YL��e��-��P�
KmI��b�%AXɂ��+%���11�(b�V[�q�kS)`���X,�J-B�e��*�)�2��Qj)���R���AJ�T��K�V
)��*jb��G-�T�5f6�2Yb�X(T1�%E+m�V �(\b����j��R��aeB��\E�TU*E�����Тc��1�p`VVB�-aDJ1��dʱ`�*V#m���9V��[J˔
�%�Qrظ������c2�LC0��VD��++*\sT+�2��`V�HT�R��KLȥE��Z����̊�eA���	Y�U�Ĭ1"֢�AE�,��
�VB�lQd�XJ1b�`c
�%ЩR�C`�P�kQI���Ԫ���Y�E� T-�LC-*UH�1r�b���*�;�{X�K�E���Ch#ز^��\�![;q����oc,�P{����UZ���q�m�������`R�vZ�j�gb�k��׿	y*���]� G5R�w�sƖXY��Ʌ���Q�v�uSf���U��~�����A�*�t�"�},�.%�����R?�	�	�o�A��wJ��9γ�ں�ͦV��Y�GMWP��c}~�*����~�k(K�.��c�X�Ǵry�{�L��s�g�@=�m������4��^�|�t�}њy���/_n6h��GU�J�M9��9,���L�N���������lﾔ%�ʄ\�BX-$��|������d���u��5ژk��Gb�y�J>��e[D�S�=���d��G�W�c��I�Wy��]�#w��Ց��zkm�C/׍zuq��R��#Vs�-0k�:�2?N�gl���Feޥu���!�֑y�!�N��ظG��r��"��ڀ=.�ԏ�s�]*#$��J�W�_>/:�t�t��C�#����+��Ϯ.�7��9�N`mxn��l�+�׵p07\E��Acq�Ɩ	��@���/}f�ǂ����ͬ�W���,�T�Ä����J��O�X:x����u�R�ݴ�
0�w�k�oZ��|}ME�2�� �{��}m��Pbz:�{�*,�+^H�W^�k^^�\>1�������U��b��h͐��ṹI�Z��}v��.B��8\�{�G7{e�|D���:�r>�3�#p=��6L�[=]�ν�L07��;-�=��S˲���V�¬�s�-.%�n[3��w�,=C>�.wV���Y�V�뚵6'*JOq{�V�)m�`.��ϫD��&Zu��n�r�Υ�5�ZZ�cf�FV^�ߟ�������{²�f��3ꭵ0R��_����D�ΌP�ȿ[��gX�*-<���0�v�C�q�����e�Vd�\���"�U\f�#�
�l���5ق3�p�=ɜ��Mt���>�8;�3�1c����uK��H�W
	��վa��U���/����a�C�Up׫�Q��h0�o{<o��5�P�K��$K�h��KA+��2qI��oy���.}B����x���.N^�7�ό&g����d^N~>���9�R]����=E4�(� ��ʉCc��0s�5�/�+�����X�ر�'��ץ��a{�n�f$�6Rү�N.���>^ҙ��Z���F䬈7g=B�4�i>�پ��Acq�k�6��[�3��4z����Ԏa�+%(�N�i=v���C;3��� $b���G�,L��k����&�G�5j{�&zUq��+�ȞVuH0�!��6���l9�9X#o�>���,K��B��u��aC�^m�?�[��_�r�B�¶H��5>g����u�όuy���w�dOӎ,(��o=u��l��Z0	-72��b��H�@�ؽ�..�?*WUн��w6�[x���Cmq��t��(V�,0nJ�Z�����gw��<��v��:#���B��{����k��¬��n(|7�y��e��MX{p�/�=oJ�J�Y��k�Xn(�3a�w��I�M��T�ϵz,]C���ڳ�mH�7�x`���c�l�Ǳ�g��6.`7��zya�D�[J��&6|�񒗝aq�
Oi��(h�V5�ܗ���1\�b�5eR��ݏ�=�ڛ��뗧uxM5���/ ��Q(u+��_
�Z�ѵ�L-�4��Q��^l?"z�<hK�-w���𬔘pn�aq�Ih�~`X�¹������Bk���L�8�{J+2u	��oV��j�ƃʠyW�jZ�WU��ۊ���{�+{�n[�-Jq#�`�<�M�e��Y(o,9����*��t��Z%�O��	;�fkŅ�C{��/Y��ޛu�e�Yj��B�����X��m�*wdg!�Ѣ�:~�j��Q��꼵s��X|<�IT�<�5#'W�;9�u���XΕE|�a��˱:�F�P��"i�}u-�+7),Ũ�t�R���S��ܲ�=-�+�_�~pc��r/rx���O\#��e�/&�5g�{�x炅�
�cyŜ]���ɾ�z���]�~�h8N)�(s����8)�����fP���m���]*J�N;���篹��P>~�s OȘna�k�"M���(8�/+��9-�hN�Sp��z�L�5���x[�A���1O�2����W����~	�H�J\��T��_3��t�W���JwD�{-501�*_0!����v<s拉k��',�*i%��"���墒u�R۷�����ysQA/��R�foK����˶���R�a�z�LޅScZȥ�S6�G���%�=Mׂ�]�����37��L&�ЍbCL�t�}OڮP��VU�Z�-�<	䤎){Ս��QG�b3h[X=��Sˢ���h������ʍ��˝�ԗpXO��X��n�J��j�2R\/ҭ�Ln�O�-�ǆ半�
�u�e���}��U�҃��@"Y-�Vz��ߠw�Z���}�gRȡ�1�d�]3�-�K��iN*�ޭ�d�9�����Zi]����8!��enSHH%_)o��<��tNF��)��pbrs;ui�=�P��kLDVېf����f�oE5��u;�i�.��Tft$�⬦�ǻ�������k��kuY3g�ݩ�Z�٥��r'�9W��n�ve6Biz�{� ~����:&]�6�^ �ɵ���7��Q������yv^�#��`wK�����Nm�3�x'���x��xd�7 �����)�MX�'3K'yc��I<�'>�l�L�N$s�T�g�nn�`����hxN5�Xf&c������1��:���ֹ48�J]*���--��T3gZ2�`O�����3�=��b�M�	]��9�S��f	v�'��|��"9��v;+�4��XY��L"]z#����G�s;��8�{��I��y�؋2�'�)r6
�����ԃ�]1�|:l�[:b����37��sj�"�z��u��<�س��p�H|�.J�S1�5�Z�g�3.����,�ا�o��9x^��tv%i���O/CHO����L<-C�#��3��TY3�W�I���]�/�	꽾��x��2�~ ˶w�JփQB6X�)���i����X^s�^Vc`
��o<�\ZO�����3�{�vVk�3��b*h�
�"��x�[s%{�Sf�+��`uӔ�VF�\��o����*�o�:�v�]�R�[�����3S&��1v_gP��J���������8n롐J�%S&�w�) h�@��T�M��ƚ�\~�.k\�7�D�r�WECE�����4,�λ�/%�Rl��)�|�R��HV�^m-��ӎ7v��uq�y���VNz+����V�i��o+�k�&�o��o���6��h�el\�y���7�p�NOx�&{�t������,U�9�3:�������A�C7�+���<�G]�����G����huj��wS����|���-J f�676������Vd�S+����N!'U�ū�#�ͻ�G}��D}�zc�Dy���&w-yn�^��&v�x��^6�W�x���q�K�]���*��g
�����O��f:�g����&ʛ�x߷��;#�N�b'nWw�ի���6cf�������0B��9��X+K2�ws�>�����}��T�T�mH�ӿSp��＞���e���ĽJ"���S:�\�J���h�8/|�RW[`���t���h�5lL�	���ol��g�Vf��\���E����TGGϺ3�`�sȳ}�+�k������|\�lB�?P���f��#
7N@�̿��᳝�خ?^yN�	��K�
��/�=�N���>��Ƹ����-�.L�K��z�}���{���e���y;[=�{�f���-�nzCS)k��w7��X����]�M����?<2��w�*ּ���0�9��"R�l�Wo/S�Q�����*"�מ�2m�x�B�9<��~�xf��S�Z愵{(�,K�zMW{������:�x1^�K���^P�.��iK�l�&�Zݮ���Ϗ�3�̧inœ�x�E��t��ks�5�W�T�A��gԹ��B��ʉCx��!�����L�K^#�Q���u�/w�s�Vu�dy�����(0g��G�z�]���S:3�j��O�q�������'M��[��hڮ������"��G�y��Q�:�c���>�����U=m4�o%aʄU����)5�$�t�˸s��K�g�D����S��B�s�חx\��ƹ�h�7�괕�h�tA�[�����*���":�Cӳ��һ��O@��p׌U0���v���s��V=���'�}wt}�gXT���H�.�c�qm�����^�.v���^՘*X�x��<vԋs�������6t���}��ɳ}B<̎�:>�j�`�v8�Y�tW�T���XdP�l�b��\b��&QBP���Z�fc��!���҇�Q�>n^a��vY�q5;�ނ�z�']�P�nԐ���9992�	
cSv�(�ptd�7�[�r���k	75l���,2?6J
�ŷM�Ί8�6��WG�B�KϦ�tmG��|���6	N{MV�m�fʘ�f|�3VM�ڕ��)�}⨷U��U�c �|`�c����OGNsh�����m�ڰ�fCﺥ�P���=��*���J�KM5�UWzD�+��%X��v�7{��. :���WbQX2u	��z��P�,�*��IjZְ��>��SΪ�4����*�2�ىԉ@��&�2�N���Ã�T僧���%{�c�:݋��NR|F��%���O*���i���FeCFU?m߶���6�yN*��%����a�Gx�<k�n��y�@�,��\��B�;��L���FeC�4����r�w=ay�IC~�����e��~���@/�� *��ѥ]��\�ј~�����[��2a^��'��ԧ�҅En��`��-�}=���/���<i)r��t����y�a{ A��g6��F���=kV`�ȰTɁ�T0��R��%	���*)%@t�_��#6��r���~]'�w6�=�c�j����I�Ɲ�T�|��]�pIH�"X�˺�(��C�����{<h�B��7��z�l���mŤ#m7�*^�����ɍXj��Ѯ�9K�,��f>������W�]��0M��ٝɜԉNcK�WB� J=E�ٔ3wW^�#��%\��>�2gP���*uhy��垱ç��+�k�d���I:g��\���v!�^�g����7��O��Z�F��2N�R�y�B���X���'Y>�f�{h�'Ɯ�~4��Ӥi��;3꼵8{<��;����A�!�~�pR��E��5hԚ��p�O��s���z�@A��1�+���`����C����X&cỔ�4hu�����ZW�JK�`d�V	�||0noy75&k���uV�gݔ�c>۰��s0o���OK��tL�hmҼ�971_�y���Q�z���ݬ�M���y�I��L�w/��Kz��EڮJ��X�ڇ.���wmOpo`�"ڟR�S)�*��`��9�*D�	���v	6����/�]b[��qN�ޙ�ذ�Yj!kM~䟅*2���2Ұ<�C7ӱy,i��6��#7=�0&���6�ۮƣb���H�T��h-.!�G5�]��\�Vf�{*L��{[�w����g��gv�
8V���AL���p	f��)r6
�	q~��R)Wf)��T^yAzL��{b��Z��ڙ݂��}��K�q%���ˉmj��M����3Z�U���vYg'U���&4�$��Rg8�%��a/%�RC�^�Ře�θe����3�>b��v#ǲ�N��/2�Pl�w6������2sw(�Ú�ؠ�%��[��W,룦�����?{q_9K���cHn'�{7�/��w/.I���p"qA��~1�bu�������)j��S�-KJ`���@���G=½[���gB"���W���7>�@y��v.����.�bUq�����P��{�_��gm����(d�I
3M+����zǫ5s�K����2�/��`���O�ˋy�l���(9d�hR�����3G� ���y0����'O�W����J]�.Q�R�^Q��F��׶X�g�=�	��2��s�C֝#�Y��pu'��1�	�-f�왭�o^�!n�%���W�1��bgVt�t��ۇ 8F}G�P�T�:��j�n����~�-�/1��r=���a�5춓�Z�%�էoj�V��� ��kCM_��ޕI�Vו��q�C�����{J�6+p=��6L�S�ݎ�R��Νg�7���
a*���$n	~�85e�ğۖ���f��,=C�ټ2�*;�X�?zu�)S�O��*��9�ř1�TѥV��fZ4����n�-�ƪ��*ڷ��/��Տ*�Dc��{b�,�+h���wVN����f��KZ3)�;b�D$�%��;�7ɖ���yCkR� ��.�"xdc8hS�74��X�Ŏ�%}'d�ſ����C�X#t�՚�Po���ך�8����N��TA��H�6��\5����f��|�;Yރַ���;�A�^%t�e��H譫�ܱBT{��l�����Q@vp�`�(��oѾ��h\�m�+ȵ����W#��;�2㨭qBj�z!�'IX���N��Ac��+E�b��}���Sur�+��X�K[�o����Sh18-�"���ȃ�(�n5d+�*�b����9k+���{��g�Ő(S\���.�z��P�S��]��c̣������&��P7�=�;�w\b}����\2ض9��Vi��.�*�n�I��T������m�u���l�1�������;�ې�+	8 �ub��
}#	��C��)�.'c�ٓ��i�wjh����^�05�0��4Z�����]K��7�Wk<:���0����l��SBA��������ʛ��")�_M�����L _BB�����J���#�`�sv(ݬ�r\���]9j�*����r�aѹ�I�KQ]w���^i��7\�������b�N*��`�$��q�[kZ���N�)�{����@�k���I���cwf;q�e4WVF`̲�t���ֻ�WHA��@̻$j�k��b�h�NV_=3�˞Ȯ��`Ӷzp�Ȳ�3�I�*�vK�##�h%�w/&#��n��u+�ct��v[h�b�u��*ms�D�i�&%Qd�s�)���ъ���l��c�P�����+�3��2o]�@r��/w��V�Û�i���F�3LB{]��+�jYՃ��6b��h�*L�]��2�M[�0ɵ����`vb�{� n��ӷ�[{�>�_��BGi[�\��ܝr���qsd��q���շ��/XY�zC�tg5�)D�n��ʶTFz���$�\R{��C���N;�p���[ ��	��:�
0������
-pc�+Z�.Y���2gne�իp�[F�	vX�#̯��zR�����6;f�It�LUr�Fn��ϧ����]@�@ҳ�psG�j�V�	�[��h�e�A�)\ƪ�'>��h��0<]C��f*z1y��:��w[jfjjo��a��溡�2v�܌;1��B�����c:Xp�S�X����iTĉ�J��wZ{�6�b�{;�1�̻��Q,43M�7�d6�͐��Q��*TkU� �h��E�'*:���}�w��3��Ky�1(���mŜ��k��&��T�[˃]*�-r=�V��F2��f7�Q-�X����� V �Z& b
�2��CbLeaXVR�(,�ʁm"����+%eI+F$m��aP�d���"�RT"�"J�%j,��m����(�A�����j*��l��R��+R)m�`6�Q�Z�Y
�D��!Z0�
 T�E�i+(���-@�+YUbȡDX֔kX��H�J�X,���dR��X�*ҥA@X��P�J�,�`���YF(,��aU�Q )FȱE�P�
J�$�KlQe`���-��Em�Y
�R(V��H�F�T��%T%dR�(TՀ,m��`(�2z`ŏtB��sw���|o��d�ҧ�ʷδ=6��?*hyǛ$1�qV�3s�;,�]s�x��-.DhG
�+����lk�o��ym-�C��0B��K���e�+K3W�K���{��̏aU�=�X`��8�z�g�!�Yh�aq�3>��S>�qP�����.��u�K�����T��x�jx�,�P�r���8��`��2ʲ�ߗR�l�E����Býtwo7d'3|Q>�V YƦ�|'R��>�Ǘ:��LVh��HӐ��
/�l�W�"I�:�2�;�2���0:�skA��[���~�ױB.(��1�w���*�e^��sqU>���@mJ� ���R����]�]9�eo(0\�����H{ޗ���z����e�w��#@�0t5�].k��3�TJ��!�P�3<z�Z���J\ML�קN卞�yi��+�i�>ߪf�P`
?g#��{�\n�K�����tÜ<��⋉������Ue��dC�]���$5gF;beه�h�;,캢�%J��dɼ|��i�Y���v�Mf邒�*V�`ȓ7[�������L>�1�ש�I�� ���rڑ�%�����X\#D���y^�����&��O��̲�:m������'���M5&1��Ľ�i��h��%�C��ٍ+�`^i���m|���3�ަ��S�X���;��7h�\��|� ��K.����ԙ:�f�QQ����h���c��z����6�9�.���Ab��W����I����'V�p�vz\��`��f{�N���P�v�����#èi���[�ۄ�I�zP��+}�����<�<�t��<ք:��{*[��ь������Z�����I��%��]�7�Gv�i�����\?E�4��5e�])CV��Ƞ/���a�����ۮ�$kw����.u�b�ŗ��˄o��Ӻ�����V^Um��P�W�P�i�b���n�>=;�5���{�b���|�fC�oW���͹�^�@�u��=>K�u
k˴�7����x�۵0?=`*}K@j&2�=��'P��~\6
�cA�̫a6+��d`t���?U���Y�J��*��w"G>�(O)��'xV{)�mu0C�5�2������y��zD3ID�-��*����g)˚���=�ɗ�M�j�^X�qn�'2q�K�=���rݪ��iv��#��@���q.jg�(s����9M���=p�<��K�S̜��M����O�&��'���)_{G�l]��Jx�h�5wCo�9u �p:�x�@����ufv/Oyク4��'�/o.��j����:9SHu��*N����~�P(�p���/4̼}-�8�FhulN�p��#�p��\�%��[٩7ױ_J�^�ͻb���̿[�!��<�@*�D@�/�A���A�ƞ���}Ә�v�oG����P���QC}���*�{!ßK�rx�5җ%uL��ᡰf<��S�N�g{ͫ�HaV{���m.%.X|�8$�k��',�*�I#V[��
�^f���|�����U�3��E0{�rÀo;����]�pIH�"X��W/�g�k;�MK�Z6���؁?%���3A�qp����3��4��:�^�#�D��Ob�=P�t�Qc���0n�>��uE�
���(�O�m��������/O)��,��HTع��[���s���|�Om�,Y^�QZ���K��U��N�7\"�V3)���۰Vv�Z�m����p-6�[Jo��ިxhzpx:�ma��xdK�[v�w����{�@;=��賘z=/d��E���m�q:�c��4�OK��k�_�XB�hfL~������O��y1����c�j�S���0��n���^	���a}~�xF7��\�\$%E���r
�1�\�I,j\�c��7㹽��<�<+t-ɨiT�B'��-x`�to�\��*1d=}~/Uz���e����lJ������5�c����d8x,��z�	���u�g�n2�On���ܴ���
�������M�S�M@�W+�iா*�5��9�*D����v	�M��[v_9��~8���5���!���Z�Mo�:�E�P6Y䟘�f�v#7Mfe��죣�?t6���G[�'.�{����]���x���X.�g��X.��[�KS��P�jHd�|_��N�Y��s�G&V���AL��h��K4K�r>��0��8��D�W�?H]��R�VL�^�:�OV�ZE[��Y��£��l2��Y~�Ѡ���:M�6}�,sb��I>GZ�"���Ǧ��������W�T�(�ʘ�����^ad��G-X��ɼ���C�J�T.�]��@��o�l^.-k*e�Īg�	K���ϸ��ݳEn���t,W��Q�[��Y��7K��9�~�ab��)�?'ۗ�<G��.x�v��Vd��Woy�Wyv�Q�%��4`�q�e�iG`_y�ܮ���~����x�Y���6+9�7!��`�d颋9��Q�H���L�Ƭ<�09�}�����������u�K�i��,.f.z1�&�.�P���Չ�4M��G�F�Xls�x3��[�<�}�m�Y�����h���F�@���	F�.gr�{��eFc��Ԧs�r���J�[���'V�9"��Q�\�Y�F�o!�zX�AB�y�`�3:�Y>>�T<���G��v6�g7}�����w�Z����ͻ�7+֠<:�,�X�f4�mk\��j�{�pյ.�n7Cwڽ��UO3i�}������e�b�m�^����9TG�=��7�2M۽X�۶��䏕���2��jԯ�
ZEڄy]F�3�Y`��q'�;���o��k��k�E��x%l6�{L�#�.y;��/��Eh�s�g���jt9 �Z%�s�)����[W�P}���T���6�be�C�WylͶvVZ,�ˍq�U��
T8���9H+��&�ܓK1�w�`jr��\КP͛=�YVS:��"���u��r�idrAo���˪#l
�̬��j��Ld}�p���>�8���=��%f#Z0:=�{/����V ���k(..�;��S���|�-ͭ2���qW��gB��o�V#+�b��z+��龪zH����5KA���yB���Җ;di��[����fs�:wֹ��׮�=h�����3��(��ʥ;'U��['9��.�V���&L��<u)�u�r�j�5}��]Yl�3�>Z3�|��2��Sn�,�gPB	�K���w_˒&��&��d4�ۺ�wJ����~�t�(d��m��qSrH<é���'���c���޷��M�!��+��vP�{J���0s�5�F�Spl;]篮���ӣ�mx��Gˇr^`% ��pT�x��iux�s>�b�>F�=/z#��.�v(���?v�xHjΌP÷2�Á��4Y��3��ZÕ���ۣO9^�3s�xk��oK�|�B*��`䔚џIh���,z�_-��}"8|o;n��ᘻ�×�fo�CmC�z]%o����W�{ؠ���Sw��"��ug{�WcՖ���a���q1�;^����E֪����}��
����y���K���4�T��ݐ��b�Ї��pLY�{Do�oG��M&}�zfl��^C�Z�����њ�[��9����7TkN��v9��U�~^����28�v�����dV��c�ބ繚��\z;��O�P�Y6\#.���~��?�c��c>'�	ig���B��(c��d���#���(xΣɬ���+�d>��[�衇{�0B7)@�n"�<��Og�( e��'u��o
W��v��oZfud]I<�2h�M\��}��Y�a��W`�t.�(r��Mh��S.�B,s���ݼ�5*&{B���N��Lt��n]��w����yaM��̠ZK�3@]�G
J1o��T .��U����	��'9�\Ҋ�2u	�-���Cܲ,h>Z�)K��Goľn��u�=R��̥\]J�ө3킄�ɴ����*!9���FOf�*�a����_(ߍ��*#� �KA�آ+�ۧi��O.O\#�,�/�t����y�c��Z������|=p�U�D[�JP,��K��(P�c/�2���9(c;�{�z�.}Mړ��D��w����?zϧ��,�s�D�ba�k� �Z;_ƕw�ŞH���G뿗<��쥛�hl�g�`	��'y�;�п)�o}s�	�t�%z�!o��q:Z�O;�˭��
N��"�4'�m�u{�B��2`~2�xȕ,%���P����T�E�#NH'�>�����ϫ��I3��Y�S>�Z�7��W�P��v��"0�md�\݁�㼼�uCު��=f� k=��"j^V���ѿs�����y��ջ~{�Q<���=yZ��@���'^�m�f�h�'�9�sƝ}1S�.+�ƾ�Wu�p��e��[V�V�+br�Z�"���CB��U܇XJ�w�+������D&�����#ӗ;4Ro��\91}�N�So��s���7����v��%6�E��/-�vmVYs`�x��j|�Dԏr��3s�c��!��b��&(�&�"�PJ�'c�:�/����6;	��*�n�6����'�3�ב��ጩ7z(3����Ƙ7+�p�ܱ�ap-6�ig�v���6�˖���[�y}��!+�8:���~Q��s�|���;1��\D�aŕ�k��l�}��.�t�9Ʉգٔ��%�b����
��:ҬvM_
�w�v�3�Շ���^0ȻQ����֪�O�~}���hr��+x�j���]�/�����>jD�n��2����<��������wi�}C�S��3��Yk����6GRv*0]�x�&ZV<�C4�KO��{g����H�7lB�s��t�`��E��o�ƸK�v��J��}Z	7�؂��!��� �ݶ��w��k��W�wRѳ:�9dg���ν��!�w[� ���CM@��vtW��u�Q����%֝�ͧ�g�0�@����P���͡S�62kʖ%W��z��w���k�f��Sק�W�T�(�ʘ�};�^��B����V+��x����fc�{	f�j���7y�u-�1����ֽ��^⌷`aI������AW]w;5p=�Y�b����E͙�s��#;���fGCU�q��r���� HgbT��^�d�l�T�xk��A�
z@�H�kO.���#4{ȍ%��xs�߆�T����qqkYS.�.��˾��i��/'r��ֱ�^��D�@s��*�It�h�M�m���e^��^rW��������[�x�~������'9�z�J�ʢ!����]�t��r��QZ|M�+�l9J���{��;t����{��9�6$4�,���XC��!�x��4xm��B��,�W���N��"�`�y�Z�C���K�,U�9�3:�<GM�͸E�e�������ۭw8��="��Edl�V�Eqћw���Ýq��,n�Y>
�
ׅu'��aȞ_�Ds���j5��-�K�ǥ��Á��x��c��#��ی����д+ٙ��J>�_��w��g�:��Ԫ$|Ep	��_]Ƴ����<���}�lɛ�w�cҽg"Р�͐�c���ؚ��Sv�J���_�M\YKm��/	PMg��L;�}����x����z���a�k���{��Y�Ƹ���mL�C��x�RSW*�:��2��T"��ѿ�W3481��`��ڷ{[�ӥ���gB�n�Tb}�ͽ�����9W�� x]�����)ɩ�;ׂ�:�Ĳ��& �M�C��c��؝`�j���>�B���wzR�n�~�z-K��鸌,�P�����ol��g�Vd�\�P�������S����Mi�S��0�!����A��yt�Q^G�G>,�,ϼŎ��o)�e]O;��D���a�I�69@�#��ş
	�`c�-:ߝe���x�'?i���f.?m��ۉ˫�Gx�<+�n�"Xwh���l.�^P�e����v�Ӂ<���Ng!��zsD~g��k
Kib�~��]�Q�M�P ��֥b�5�&{FTJ�r
)uk��zrޓ��r���{`]���.�->�ȯQ˗��Y3맰���14��xE�L"1�/o�z�}3���'pϳԵfo<lIY~2����0��.�8�hG`�,u+Ű��^g�{;�9�x�z���3z�W�))��.�;���ђZ:e�Bz6'#�^�y���V�ȑdi�Y��/j�ݡ��ޕIs�,a�xԫ?{ؠ��x����r�ޣU����L>w��#���=�b��ʥ�LpT�z�e�E֪���o�
 8�����F��-��ҭF^�3lg}��V��ڽ�U>]�Q��`7&;ۈa؍K����0�䐮#e��f�)���bU��Eno��;*��0�"xlw!�������-j�o�q�ŜwH��d��-���b6���Cm�J�(�j���)X�L\2lu�
��=��.��0�������gc�*��T"�˚el���Q�tlUʲ��4�wn:R�^��J�NیS)�b�]3��x.3R�w�;׼ҫ�����
6�j&���޿c�#�1�)�Ay��#X��̾���(��˷f�UЙˊ�s�k+8���-�z���;V�d�!�_9훥J"y,oy�_W3L��Z�N_	s�8M��%�L=�Wו�,W�ʦ���$�ӳ��� ���#���h��kuaͮ.�rsY�M�n�ip���u��)T�&~N�°�Щ*�:���X`h��}Fj�#�[[c5T��X�8�	���o�<̕�uE�9W�7�]��Bno'̷�z�3�B�lugGuc=�R�p��/�7cHv%q(T4�%m�Rd��u-b�T�O�j�T^ox����<;�%F����ˢ�a���n�hn@��td!GF�����32�i�Pp��)]o��Z�����q�vo�
�fh�C�=��ap�ˬ�ɍ^��ه���w��t�v�N���jV�r�:�FT���0m��N_Q�t'Oqe6zVf�vLڙb9v^VrR%���W�a�$��pj���ʹ�'����W2�Zq��}7�us�}t�㹛�n�7����͵�Venp���2/�c�+Y"��a�V�����˄��O:���ʷ�XL�5�r^���z�m[D����o9�v�[�9`�׽wKF�������Ś��
len&��1XR��9.vR��yۗx�Lĩ�:�����-����E�3س�\��[����۝�]Y� �F��]5嚒k@ɔ5���\v��"}�|�p�}3[�X8>H��,G�u׆�N�d��S��W���n��{"�d����r�L�Ɨ�]�E9v��f���#�ԋj�!�l<�3FˈI�i��aZP&��t����������5��)m9����)��=�����]_K�.�|�8'o��+a�sʹ,�M�x�u7� �x�Z�S����R�+��Xǫ��D��X��V`����=څ짼�q�5��|-���{X�.-�mZgz�=ѭ
�E�/fѶg����'b
����qf.�܇d5�l���Vo#�q�r�>j�EϳK�X�Cm��un���7���#ت�)�մfz��Tc�dQ�Z�%�ރ��՘W%Ԗq��E���pnwp�E�r11cYZ�q��>�!H�C��yzp�ѻ�Y1ƻ���B��z�5��}��/�o��c�?���H'︄Q��R�T��J��H� �%�jV,�jōJ���A���R����--2�A��V*"�J$Y#ZJ�*)PU�ATm�R��0�UmYE ��"�(���AER����Ub�lX�#
��K
�µ�Kd�P�Ƞ��k%E�� �H��AAX"VV,�AQX�d�(V*��AJ5#mDH�"0DX��,�`���E��)R�eB�b0ը�m��)QE	D[V��U��ѵU"�-)D`�Q���*�Ũ*ʅJ��QDB�"(����H�J�X)R�J��V�K@Z
���Ȍ1"֤EE �Ŷ��Ȳ�UU���TQbZ)�u��ǔ�5?��t��5���_���%�4�p��=�ON�%AH��%I��O;�rŝMq�.�r�m���i�k��wt�Ȭ~���3+Қ�g�q�2/:����t4c>����"���g;�Ӊ�N|X�n�\����89���^oi���d�j�����m����s�5^Xd{m���3<T�^7�7١ca�\=u��w1i�B�d�p��^>�٦��ۦ����̕m��������{�$�Α��h�V��ΣN�qw��d>��z(a��L�ϫ��\t1kr��<��u{sԥᇉ�q�$��rɡ|*o:�l�{J+N���^�E�5-I�	ӎ�R/i	Kٕm�k^�e�*���e�;�#�!1p�H�'xVm��7����d۷a��3�V��~6Dq%��u-�`�\^
9������>�[��~Hm^Xo2�Vf�ҥ��\۝�����cg����"�dh4�52�v_Zf{�{�ZO`���q�IS�a���[�=��s�e�z[��	�g1O"a����t�4_vgeg#�!���nUm6�Pg��X���{��<�x��J��߮xA�)xg�"��{5y��wf���� ��{�"�qoc��$��;��cazgX�
�r5���(W��j�U��N��&�t�C-=m�f�fb˽М�^�����Szk�(4��FMsp�.4��Z���[��
�ǫz��=���������M�N��>���`�6�&ZԿU2:��D;C��6�����ŕ2`~2�x����	(M^~��S;;#;]ޅ�+t,9i%+܈�2���M.���zΘ&o4Oa|�`�����&��~���ؿB7Ȋ�ɇ����l���h�˥��*�˸�_�7���h�����K�q:�;����su��j������|���:���l�J�Ye��R�y�s=�x�����<���^���50��ҧϮF�{#�/�gK$P���;MZ56�Z�ݬ�k��� +h�KކTO��{T4Ͻ����卋p-7�/�?W�޹�������[�{0�nkz��Ɲ��&�S���S1+3}����A�nË���DҘ���v�]����v8��	�R�L qϒ��ūu9��{K�"_= Lk��;��y�oV�l�Xzte��b#�h�T�:ȣ0�X)q#l�.z��5��>aH��p��-ӯ7�N5X�u1�9WM��8�ޯ<��t�-4�GRw�*3��-&������ƴ��];�r�+��x\Iлt�x),�����Rmj��3��p�l��m���a��S�fH���p"U]|,�/�����!�&�ݾ����]�����>#fS|+�T�I5�P#���U��:�ك� {M{"�Ts�]v��,��mà��h�]�ہ<��^@6b.��cL8���@������R,�+A���$G41ݿK�Ó��o��&f��>���i����L99أ�L��T�3ϧ�rY�h9K���������W��I�<g� ̰� ��珏��Sx���+�4z�n�ʱ���}�_��'<�G�x�ん䁝ԢIC"�	�|P~�M�	�3]o�=zq��5xd��Q#�%����.ނx�ig��
�����$��ޏ����f|x���A����j��|;�*{vq��*ϧ�Cm0r�B,K%��M,ഗ���|߆�xk�U�;>�~>�j��c|�g�/I�^9k��K�h��COQ�;r��m�4%��1�I�BF0�{���3�g�s�R��>�#0oL��F��2�Ć��7���k�؇�XW~�,�ԯ�o����^������>	�B(���X����13�#�t���/�r%����s{��)�!��Z/��Fm�3�o�q@|:�,>���{1��b�:O�l�|�ZCn%�gm���M5.ĻJ��ʃK0�
4z�;xr3�{0��BT��`��|��i�:���P	��o]�1�M��cv-��jQn�v��[O�5�<-�J]���;ǽ�WqYݫ6�*m���6��f���\�z�KԜf�e��y�����L��֏��t�X���8p>"�Ȏ�x����X�M�S-�:���8�Ӎ��� ~Y >3]�a��݊�dyP��_�¬�|t����2���J�~K�=2�{�Ϻ�0��z�6\��P�VZ8|����������wU<l��|OH�)vh^`�g���n�r��:�<f�~Z�!�t�'���[jG%��^�iܬ�4|�䆑+���&��1E�qm���sA�4=�3e�e����ې�UC2�`a{�y
fD��h��:�u�Vr)�өEc쏲����1C��_���muL&��ڭ�bzldn�F$x{�Ȳ�f^;�Ӡ�u��֘x̜����=8�g�^��o��լ�5j��"X�ť��.�^P�e�4�:dx���<~�����Y���+|���m߆9���'��Ϣ�"\�A
԰R�(S=eD��w�C��ݺt�UF&<�te{q�W!>ݖ5�)����ŧ��9r���	g>	!t�����^��W��0�{[Yod��=��������Q[T�S/�k��6��1���YLrW�D^����V��)��{5��P�Ҍ�.ۥW3�4WtѴ���\�L�ks��&�9��";6i"��f�:�P1���[���و�J}�K�D�z���h<��ڵ�Bһ��)j��VD��oT�Q��0�̻0�~4�p/�4na9��*����p�����jS>oz��������P���c$�֌�KGJU�[�d��I�<�O
�SXg�wF��F��fm�~�j�z]$�
�X`�������+>�]��<���`cY��5֍�ia���s��T�z->#GP�6�Vt����g@�����9컺�s�����mx�Z����'�8�+j��"n�l�����ב����+7]{O�����6t�{#�M��{�\54�ƛ�Y����m17��p���ꟼݼ��#��^ x�&3��f`ws�|�/V	����Ӻ���v
��2�o������K��si���:�Q:����̇ê[��Pýr�#�Xq����G͖�:OM3�Γ�qĖ�^@[�^ :���Wb>"N���L����[ע1сꃖ4&
�yW�j[�E�\^r��D����ɴ��O�l�Y��oO|���+���ļ�����Q}'5�I�u�89�P/Vo7/3�G������3Y�WAœTk�>�>�ۊ���HAI��5���gY4��q�{qt8Ue�Y)VU���C:�k�K�Z2���,�쨯�%
xy�*8����)�|�يH7:Y���݆�PLz���<TGI����DW��v��N\��Ӷ�Po-��ǝ��'�����Kɷ�Yc'<���=h�@�F�A.kҕ*�/o9Ku:��)�~����x������ï~RƐ�<�==-�g���s SȘe�O4�>��ԫ3�ؽ��|�8�L�Y�ѕ�u`�t���	�y�t/�E-z�Od8pT�kx�>���S7s�]���VD|KK¶������y����uv,���a�%+^0��1�Y.�������Pl���$��#��^Z):K�����^���t�0����ÆC�F�����>�s�ҫ���Un�M&�� K�
yX�\}��е~�g�����G�v�̞ ��O�M΢���{w��eF��!�I��O����^A�[�i����
�{ԋ8�7�S~��zs��Do�踫�F�ǈ����Y��=~5�֭�^�B!/��q[��9�>�Xu���A�v!������e�����Ϧ���ߪ<x��\�l�.���*V��:w�~�=��3ujylF�w���>��`������7�k��*�L��r�9��6���ٻ��z��7��o���5�1\�Pt�rk��ws��*Z�.�Z����.�t6��4�N�-����:��L%æn�wǳ;�5��}�W�"\0�S��2��� ��aŁ���M(�����#�ו����<�+׮灺���e��X�e/,�`/������G�9�L�������G��Z���7y�ʴ�cS���ڽ�X�t�g�iՊ^��+FS�'8&/�f��GV��m�R�xD�ف��M��ƞ�x�ଵ�Z�A��������b�R~3=}�E'��� �U���=FX�cL9�s����1���H��q��\C�X��ڲy��#����R��v
�Zl�=�d� ���[ޫ��p�[�p�a���o^Ǚ�
��Wo��ֺ�w�tǫ�:PN��3��&�tK3i�~�=|��6�ᙋ;�ž��[f�@В�%uLưPL��4�Ǧ����ꞽ8����nz�N���qqDV_��A�ۧ^�tf���F��r����V�_>/x/�xt'�"a��s��I��>WϼzTϹ	J��B,K%���B��ZK\�yϛ��/p�<�6�E���&��˟������,;��}ٍhGN�
k쾲��El�:�WaR����W&녵՗���#q�f�֝���[�n�\�L���������m��dqsC�k�cYYZ�7Ø�{{'�&�(.�6R}-��Rh��S|ד֖�N�t^1B�ʶ��=G0��*����hK�]�b��^Ӛ����+��tjo�a^�jk�#0oL�=�՜��L
~K��E/�Gz����>8�_,��N����g��)^���y��]�g���%���W�1���L���<w�`f��q�ݏ�?y,ͻ�An��7��/��LK������s�"�Ac^�ik�m���u�-�4�'�������2�[!������c�����q���������f��kn!�+��8ë�>dwms(O�ɝ�b�]3�N�J��ii��Wq��e�l���E�(p��KrBsy��%�\{�ݟN���e���2T=ȭ�μ>����L/7��ٝ� ��zt����u`0{�qk+K2�����c�k��{�WH���q����J9I�fl��"I��r�"�������ъ,�����'/��h{�f2϶�(O>]�ϗH��i<�Dj
��)";º�+9��'R������p����`�g��*���dw���|E�3$�+4�5z[/|�^�ds��S�,��Ǚ#�%���u�M�u�3zz���5�Ɗ�)p�%q���s5�뢰Mރ
3�����8<w4������2�\����d-Vr�8�/��:�.�:ݵp�R�u7p�n�rН#��\\YA31���r~�;�y^�~g�ȼ����z3�����;�"�/��ce%�.�<ZZ��e��)���7�4�Sί�D����M�����Za����3�̧k����V������S�k|8�����Kž�=� ;�Q]���|�x�{�����y.�/0�E�F|5�Ү�$���qvm�-ͷ6�bw��V=�����j�ޘ(ܕ�z�!�2�u���&�Օ��No,KίX�����Z:;ZC�r�Ky������I[��f0pII��0�4D:�J�fW�g�.ȱ���h���A\:תT<36������t���(�o��g�Q����fd��i�Ӱay�u�gҫP��U,��ݯC����n�a>�OJ�T��6��9eW��KVLl=yQ�!
4ƠhL�{����;�
���x���Ŵ �A������1�h��N�g�C�R:��ײ�J���뤯�T����ǻ�|덝���z�ӵ6���͔@���;�P
_t��@�8�+E1@ k��Tyտ'/�fq	��WYQ�����*��0r���s2�ß/Q��EGo[n�dV����h�<���<OwL�V�4�.�=-�YKo�e$R�n�D)�D�l��>�tT��Һ͕���b�7-����Z|�/V	���.^��馴�}X���fq�W����/�w�Uz�JKF1B� ��u������}v��\�i��a�ײ#�5V9�~��əLW�"�JK�Zf}rɫ�P�c:�l��E���$[�u&�O�K�'7�{}	(Qc�xҩ*Q8Nq�SZ:U?͎<��F�'��9�t�%���%����<+>t':���o,��a�TG	4��-�`�\^�i��*M�}��b�y�~z��ei>�d�79�>��<l��ze#�;��Y���ʒ1Q�]��z	M60mA��L��%�^�O\:�)cH�9��}=-�g���s�D�r7ͷ�L��[�/=�� 
���j��;+���;���
�v��|�k�;)��/�;������@���rI2:��gr������;TɁ�˱㾮��:���b��k�v��C-$���*WWT�Z��*��0f�D������72��:`�v�R"k6���H?<���n�qPb�Н��m��3�}��M���9ӉuvK�eG{��3/V�[:��=���7H|��eq�`�U�����Cs�S�['N_+��r���z��@�N4�+�E"^�TI�	۬�V�V��p3U�H�5��q�h/VQ�:4l�G���:�]1�� ɘj�e���n5+E
J���u�	 R�U�%v}������Y0��9�97�l��$;-��4�,6��Cj�5P�lb��1饽����geАZ��^�����C���y���@�w�dw��;A"�Z�m}/,��Ԝ����s-���dz3dkX�C"冲��z·J��L�\G�{�����n��'S�.?e��Ҫ�Kc�v�up=�2]�v'��W8�19�h|6QJ��c� �m<
AC��X�=��Wr)i}��;C$�D���켙������N5ck���yx�ƢԺ��]W�2V$z	�2�n��@���Z�ˬ$t��h�tO;���t�C��1�e3wa��X�g	{�\�l�A��Cdi���t�:i�e8xg0���7�Y����f>@�dc�a�.Z��l�$��cΩ^tERS�qcF�ݲ���ͱ���4���A淆��l�q�qME]Z�f\D�ew+ow����u�� ���:*�,.j����k�߹��m�+mU��Rw��������W�u2z?*�U�G=�D�$�վ��j$����,g�.�(=��͹�-�`��
-���oMN�z��X�Ȼ�fvb�����˭Ԃ-��0]�,�G�K�q��]��V��q.S�˱;1�z(�F����޹f��yiv����k����7{-����(�M�`��1�z��JE�
��+U)^�n��9.�z�������8��h���-��H��Q��r-��3���.[�hVwVH��3���v%&(�3r�W2����8��3(>���C�냓nNA��}��0�0*wӳ���y���{0�n��S�'yiJ`�M���Ն�ӴT�E*���e�J�w��ef���ضgmĳn��N�Q0iRA�ٲ��ܫ6�J��!3��n�^��(���y}�|�K�A���Ƀ�ɳ����:"5+�9�Д��8X����<=�,=����z��]���̣j��^s���gϩ���8���!Θ�^)�J�KT�3y�L�y�X��b�XtTs^���&Ԯ�# �PɔQ`����5X����JyE�&K�T���Y�7��+�[���e������*��n�C]X��f)�A�:��\�g�Eԋl�î�lמ��X��e$dqmp�U3/��1�3���f���MҨv�.뻵Ԙ�;���'%XM�w�<������_�D���T�*DAJ�FJ�E���j��iD�jQQ[klY(�`�%b�Z��*�ml��ER���YU*Q[l+�DX�1E,�aR��ZE�Ҕ�J�E���AE���(��X���*Ui
�eHƲ�T��e��[J
*���%b���DZ�D+
�TQF�TFڊ�m�DDkTb �bF�FER�H���"�mhR��
�����lF��+-R��Am�(��P�-�
"*��[Eb*�m�R,m*��Em�*QDm����AAUEEb���,Vm���`���%J+*�0b1U�`��*"��k*�-h�X�[kAF,�-�Q�Dj�E�*#ؖ�-��kX�*�`g߾�>��Ͻ��/pYO}��?q�9�ɞ7���������亖��%�l�Έ�޻ԛ��U���cɹ}��^ۓ:Y�]ZYC�o"*�?��l��7]+m�x=��-yh���e�\<m�O;�i��`��
�9�: ��IX5���&B�'@�D��U��w�y��o�h_�0����n߮�L���ڼ��Ρ|�{+ا�]`>���0��$�K$P���8;���ޡ��zd��5�]'������{i鬘�p�C�yg��ߜ��ܦwx}P��~�zvN��Rk�2Z��ͺ���ڱ&u-�%Ccf@v�۰���f�4�a��� v=-Ғw�א��3������AZ���ZV��ɾ
Dt;�	8�3<��[.����|j����i�~Pd]��$��Yk�BkԽje;�e0o�q#�R��9r�l�z7�kr/y��Jo["�N�<�I�'��&&}>���XZh3`���R���Vp�f�μ�s�}�OG(�7-��>J1L͝h�>�cL%η������輗h�Ƹ�n�K^�uV�2��!Ĉq]��0
�-6Y���a�'<pL��W���}2�f�n	6w�ކ�����5B���Xn"���()�2�Ϣx>�{�@@�_��u�������>�E9��5������S70�z/�Bf���m5&�8�7Yɹ>z��ˈ0us��X1ʺx�Xd�}+q3�6viZ���ˬ�}��&
������=!�M��?	4�8�� ���U��|��o�
�~ATY.��L/3	�~XW�K<����۫�7���Hr�%b���
	�|Pe���c��}�G��md��m�	�������PPx̄VY�9�g�mq�:ho4��\�9��j���ZM��%���S��pU���sq9�F���>�S1�D%/ �P��	a夅}��%b�h��mK��b��ר�9߲w31�$<`����ta��|e[D����p;"d�;�w�����-�����\�g6�ī��(��<w[��m`?=�՜Z`�S�[����Y��{d�����fh����>4��/*R���V�߳%�^�]�f���>��w��c����}��5�v���w�Z�Wȧ�| �<��!��x^���b^��yÝq�s%%^{{�,���<�Gvh����*�a�מ��<����K��K���p>"\x=�)��F�,��^΃��n���vF����3�l�v���8K��8U�o�y�N�ߴ�+棰�7�*	k���=���q=׽�r�!��˽rDM�ع�v�̮�ݴ$�R��I'\j0s���}�]j���+2��W$N�ە(�B�p3���2�Idf�2���$���Rk�$��V�+�fI�VZ+�]�dYs�뽅�e�Y�r�w�Ǯf�KPɲ�uo�*�}~�|^�Qh���R��Ӗ|�k��:$��P�(p"��`��*���,;��:�<pN�p}����f�r�x��+5/<�H�?@���-,��*��(u��D�ъ.qm��	�懧燽\���	� ��'��[�L�5����\dYU\fuDr�l�,�SW��Qd}toȡ���f�G�����T��E�E��c�R�'H�ǋ�h&f:���v�-������5Wv�w�f,��`^c�v����� �lD���_rih6��h&f���.����^�ӽ9��fM�*�s˽4A����M����Ϣ�"D#:Ԯ�5��^~4�3���ܝr|6�L�J$��3����fx��u1i*�=r��Wd��	#�j���Y��ʨ̸���������v+�L�Υ�3y�"��z�*��(a���U�l��J�v|`�B+�h�g�C���2X��|_f�R$�g��x�V��<�Tս���z[:�8|�Q}kV��^�2\�L�y"�L���[ߔ�����&�EXʳ3��ۺf��$��%�������5�V��*�e<���%���q140���V^���`�!�;��:Wvx�{�͓2���joe��H�Em�:,sJ����:o�l�KޢF�������x��5h�^y"E�,�y��������XV�[YﻍJ�����#��o�}֍�ia���eNסf��|�Ļ�v.Λ����܏!����j�{p�.O[Һ-���7)b�Z��ʖ8��#u��J_��2�7Ir�u)I�Ԫw��g�m٪��"ϛ�l{����W)�4�K���!rLV�NuT�Zr��V2�W�타�ؠ��l��b��z�l�F����A?9�v�+�z�������ؖ3�.L�����u��8�;�����ޡ-3瞔���C�-+�|xӺ^�ͳ��EV�kUq�(�_
��:�l��(�����r[����~|���ꡐ��լ!��,h<��:�����
U�Ԫ/E;�#w��=*��3tk�^�c���#׎w�`�':���[�:x�x��9�� w�����唼���N+�w9����Lϫ��W���=���&��b��ޖ�|9���F�l���e)M��<{��B�$;{Vs�rcW�O�gSb��uL�۞���TL��.���J��+fsC0h�ҐM�;��.n�t���ؒ���a��G�����k{����TKm�x�< �%�U�gw2J�����dd>9��;��	o���ѥ-�[z�� *H �!=���S���M��৮z��Xs��g��ߖxO[9�)�L=/_mO*�>��OH�œ n�'�c�B���ƃ��|�:�'y�;�п,J���D���<~���������,ye��]!WJ\�L�����l;;��r�'S&WZH�꣫�Rn�OI����gu+^9؜�`�ne$��"��T�"�f/���� ��~�.F��r�q�Z�N���]%5i���`씈�6$���� �] <�q5.k/��,f�mmש׌��ŀoK��K&��,Hi�z"s�*��޵��H%W�m�v��B���<->"�z��+h����e{�����h�����[�K���Q�X�i,=�s�9�c��|D�����V�LJ�eŐ�^GY�z�YS���e�����2.�ĥ�3}�[�~���V�ƿ�=l��tz�|7+��6�8�K��xp�z��1�+ƑN�GA��[c��l�{tm ����>�ZU�o���0���ݱ wᗇ��DF��#�yTT��bmjҭ�=���U��{��cB��A�I�c^5 ��z��{q&��r��З�F\�v�G�%���B��f)�葽�Yo���m��횰�2��-X��]�ZZ{�q=݉ںy�^E���ý�t�ĽkoK;%�Ǘ�DŹ���0ȻW��,n
�X��^��S)��.���V۴�U�[�^�z���YM#=��K&�"é�'�U&���=��3�WK�:Pg��O(��ͻ3i�{ y�ج�y1�.�,�����*��d��9��o�kY���v�8�˸��k����K#�H�Ջwc�W<if�,��لÓ��=2��R-�3/�o$UM�;����߼#����$�tǫ�ךz��[u�g=Do�����|�����r0�G�p<Xߕ�) |��+�f5�PL�ו�B\��C���بK/�S�jLE����ߠp�Yg�<A�*���P5Α䮝B��P%��B�����<ܠ�`��ap��4���2�P�%�ʄ\�B[�I
�rV)����d��{4�ffj�S�az���8<�vV}�wFj�ʶ��=G>P÷*���B{��һs����t��L4�����w�]�+/בxN�#0o<�=�՜��L
~KGK'tgfc��+�d�_��g*�ziY�@x�P{73���b�os�R
_x���-{�w�м�z��3:�1�3�I	u�̙MD�uS]k�ޮsC���=����&�355�}��G��mm wn�".g��]�T����ĕWu5:�]=��[�7��X�3S�Cn�Rg���)���-kmޖ9,��^r�%`�^J�f8O���y�b�Vp��adǢ| �<�o��/����_�����U��1��un'���=Y����1��ȖM�k����ۇ��k��[N�+�q�u�I(�3�ﵬ���^r�{�6�q[s2�{��̡6K�O���R��tjԮ,��]�G���0b�ܯ4���qB�*�nU��g�Y�l�w3�����l��Z2T=��֋Vju���XҨ6�4.�}��$�B(r�B�u�pp�Z��̰��(|�X�Ϧ�z�D�d=K<�����uGi�GL	���
���C��(u�j%yъ)��<��'/���t�1fg����C�1�E���}��3
��ߗR�l�D��6����Y�g"����Qig]>��[�r���ݭ�|s�(æE�=�#]��;��Ӥ{��Ŵ2�;�Ӡ�WsrZ�s��k��޶Rba�|�垹n�h�rw�z��b�Aڽ�H���@�&��k���fIF][��'i�f�R�ⶲ���q����U%Y��f_A��z�ч��=5:x1)�%0���%���<� `?n2�PS�����0�7,Ӈ�`�������c|���Vâ��E�'�싃�7`;�nŃ��qP�y��D�i>E���!���+���ˮ�LA���^�V|^;�9'�� A�CZ�
�.{vkԹ�l�j���x��)�e4��n��9�̻���k��9r�ܗ�K"�F���o���M�8�d����*�9��\MG��)Eq��.ޯ}!�:�`��V�w���,_����6�"�V�G�Z�w2X��|d���K�/
^C��="B�x���4F��o?�Mh�-2꡿�ѳ�
������]b�góٜs<쇣_�6Wt�OS��J�͞���c^KDt�X�p�~��3�}�?�*��W�1�jͧ�=�c1qù�Fu2���ڄ�&Wx��uN�5�D!�ځp�w%����q��L��Zse+��>@w�}Iq۔���Qx1�Wg��Wg=�F��VK���XuW��"ۧ��AU�)�Ք!�l��n[3�ŧ�B�M��^y�T�]��\�d��>���?�0&:*�OT:����}|(0l�-E���-���g��MA]�d@�[F^�7/�W�`�qg:)�l"�y�b����Ï0�����.j�{N[�&k�b�&2�՘3�ȑ�e�	�v&��R'CIv�.���-'8���s\#������s��%ތ_6�i�i�0��lb_���G�V�ڕ'��M���4\�j�T$�"[*�8y���V��'Fݥ-�MC�(0�?.�l=�"ƃH^KRֱjc�ȭ)����F��puG3�'��!5��M#��OR3�N��X^�[�:x�x��4�KA��),C�3�F��^�`x��w�];L�.j�S���Y2�ɹ�Y�Ny�fK�z��whRΕaOd.��#�$��Cz���9M���=p��,is̳2V�:-kɲ��_{K��Ȟ��}%"M|G��B��8��+�����aK��*O���=��<7��N��7��+;r~������y�E��%�µ+�*��bժn��!L8��=nw/S�Y:>xb����Vɥz�o��rϦ
���I*�H�,��qb��4}n������A��w��|�䙀y�axe����6$��<�>�ZK�j� <%�Ӕ�Yǥt���=�<�#��T> �O}�.�},���F��!�I��<��� �	u�b���*�Y]>O���Ox�^��ŏ'���Z{ovj�J�`+M����ޛ(K�q�X���r�U�#�L`���d�7\�CY�s�M�zD����Qt��@@w)��:��M��z�8t��v^�ԣ��l�)6m�P���l��nm�=��P�ZW>��<G>�ԺQ!��=L9�j=Vj�&�m���}�(l�Q����90��^m�g �V�cn����Z|�4�i2��������O���Kv��,��s����2%�	u<���/"�^���x�3^޻g�4=���S����sQ+���s�z41P]�-tJǡ�����{G� t��'���*�ڽ��7��$Ϻ闁ܼ�OɃ��\�=²�+i�>�=N���nȫV�E��J[��@����Y��E:���M���i�W�0�U.C��;!��Wf�v�I1�N
T6e���e�~b���;�(i��Nv>Z:
ְ�t]5!��/;8U���\�=�t��@m.!�G5�c�W<ii����	��Nf���Ì���z�ݥ��W�n�m���3�f����ȃ� �k�u�v.Á���4�^�V�o��~ib�e�Ֆ�i�e�Y|%sF����?;���g�\>�/���;H@����$�ā$ I?�H@�XB����$�����$��	!I�`IO��$���$ I?䄐�$�$�	' IKH@�y IO���$�	'��$ I?�	!I�IO�BH@��	!I�	!I���e5��]P���!����}������p ������������*to�>���}���F�D��/+�RT�HCZ����+CZցR׵�lk�u��
H$wn�R�JQVXx>�(P��A
����      �~�!*UCF	�!��&M` �d�*IF �� �0��F �HMU   2    E4i�4ѥ���546��4�@�� M2L�joQ��(�G�4z�~������i�HB��`��t?5&K�Q�UD(	w�2&
(���w?��|??���.�o�a�O�`�E��Bn�$0�����f�$!ީB�n�j1P��1�7�~cw�q��Ä-B�g?��ͦ��)����i����i��m��tۖ�m�ۖۦ�tۖ�nۆ�nۆ�m�m��nm�t�n�r�n�r�m��m�m�m�m�m�m�m�m�m�m�m�m�6�n�p�n�n[n�m�n[n[n�p�n�-��a��m�'��>�33f9m�m�m�m�m�m�m�m�m�m�M�m��a��m������6�۶��i��m�[m��m��m��m6ۦܶ�m2�m��m��e��M��m6�ݶۦܶ�x'�G�K4�.���~���7���fyczz���p��f��C,%J~>J��������|��>7Ob�����
��n��H�&�2�_@Pr�E�L��V];�8�nчX�b&�c�eT*��qsn"�S�b�3j�3�1��S���MA����N�.�<9D*n��8�j���7��*l7bj�Rmdbu91�^R�&�iLe�ui\�ER�9�B������*Dr����a��7����VRf��Hĥ�DX-�r�ش,�ST8����yb�p�"�1���"���A8�Q��̨r��U77ouNZ�(ome�R�F��B j�\%�F@PhI�#I�57LT�
t�&@��
U�p����Dmj��b�E����	6v�vP+eF)7�Cp�Pa�5&}��Q1���bDЄ0�Q�q�,�bB&�1��%SL���eb&�d�$rNma�m��!'$�`�-V��ڤ�"1۪���͘q��P�DV�/d'���ǲ�Hu�	D1b�T��EȤ�֣�5����~X�%n�8��v���1K3<i�W_��X���y>��:�I�W���#"���UE�\別K�K&r4#"#ۛ˺�n�L��צj������`��E��Ց�ksZ��D��
[��[�Y�m�׍J�Z�±�g���8�dk�s�;M�3%�D7�gn�"$7f&rh魻A��6�ۤv5�t�b2�ʤ�e�+�lvH��ݟ=�%�]ƺ�q7t0+Y�$�D\��	EW��-pn�#U*��V��<W�ͷ��jâ���ݬy8��E'�Ƣ�*U7m&��s�7\!���YhF��z�����f�-Lq�&q�[��Rю��z��ը��}�"!��X�+�[Z����vtdaPU�&�󘸳�E��{A�y=Vt7�N]�8ƙ�1� +�!�!i�P��R_��������  ,f   	 �X�>5#�Ԅ��Q�D#rTD��UC� �   ����(   'ءU��ʫ�o3*32c#3����R�5��  
 � �� �� `)S4�J̫D��*@�B(������]  H X�30 �@ wL�l����ʨ�
��
���e�:7�#�SW   �@�C���@ �IYg�&Z��.0A(K	2�a"�q�\m�*V��L�����̼�y�@ �� @8 H	G6�$Af����Į�� ��dggFwI���� , $ a�u  �` (dVUd�u��څ�T%��l&ΚE��d)�V`  0P ( ww  �@333�s2`�ce�Q`�Ҷ�f�T�:L��"FR(�7[��i�"�O��}d%�R[(�$a
�w�A�Cc��� Ě
 �h�q�K
I$i
i�dE�J�z(�9>4�֡>W[����/���JR;�%�M3�4��8�o��=�x�'W�(I&/���w���m��%	$ŏ�nn��(I*|�$�|>�����BC �B@�8�7�ˬ��㴗���p$�G�=��]qv�
߼F-���W�UVo����W�b�U�F�h
�0���{���ҩΕSڼZ2W�H�~�2�.0�@��-��+ib`-Ij�mXT<��kbT75��wޱ��(4��$��*,b7q7�cQ,�Mlݢ��5�,�Kw�R�	 Z%���"�F`�aL��!�+xugBs�tx�Hoi0��V�(s��D7ሖ����4ku���t�Zj,n+���	0iA�s"Z0<ؒ:�j
�Y�Y�iP�D�f�k�έ��Ǯ�͘Խ�}�IL'lyu�gVY�M^N�m�n�[��)9���<��[f�����$��j���_�M��gv(`�B�Uwd]6a�,�:�s��l*���8��E��_n����o��xzl���U��F�sY�6�����4�o+�\�u��Z����rN�^�)V\iv�If*�!�3�5��E^W%g|�R�3gf�e���1Ni���Ūd`�eRJKtx�3|���	�Ցӽ��Q��-�y�a�i�Z�5�Ѩ�g���������� iJJ~p�T �(I*����� JJ���$��>���~�X[��+U��8(hhuZD��.��2Q�+��,f#<.����կ)��� 4xϠ~��>�`�Y1���N{ϝ�g�s�׍�B��X��M�y�(*Us����p��x�#���-�|u�t�Hr��I���Ս�B�}��_�������	z�љ�ȪGi��Yx��{j�>�Gda����и/;=� e,H{�ká̫\r�3���{�ц�3㖮�d3�Ŵ{��8��j�8*.�s�))�z�A��o^l�ժk�M��$Y��q/!����v��	����_h�k}���ͪ}pя�ݢ�B�Y'���❃O�ǏXs�y�V��ݰ�1��5o�L�T(�N@������gn$�3PHDK�<�M*]��6���.�AF�Xx�Q�^�sE�+$3{nw�*tu�>0OCUX��߹ 0�&zj��ӄ�&��	�_�A�ʡ~r�Ěq�#~��Z $ ����W���.[���&�\)�L;���g�"@��쀸��&"�v�&-��9$�B��K���,B��\;����[���:YdJVf܅ks[ۆ;��1��F�ы�4�8[Eʕ�ֵ���ֵ�ʕ��%@|�$�| JJ� %	%C���l��Ȳ �1� �fg��W~E�Ja�|�(D+��"��TR!E)IQ�(�
�k�N5�
��ޓF���vl�νzt.�� t{\{��R��	l�x��e�Bt��]�"t�v*擙���'&���<6�2�^���u���b��W����=�3�L�5�wGɗU|��F�R��n���׌��6H�\�-B�E�ï 8�����i#T�[<����!���31�X��c�'ޑ�~��N��3�'�e���gV�
�L��F������X����c�){<������8�����>�m�x}F��I�5���;>�X�����+}�:n�� ��$��I#�4�r�d1f3ߢj2�dI�q�6�U�΄M����������*�A:p�c�Xz�ߞ����άHŞVQ�Q�bM�u�M���=>�w� t�{�	2�t��l�{���T��&���0G�3=:7��e~���O���Y� ���q]�Jcl��T�����ׅ�ܞGM��s|���u�X�)�r@WB�Z��ɕ��{���BY�>J�A(I*�%	%C�$��$�%	$�I*???}c�dIuY[]<�(��EVJ��Ù�\��B��"���<lv_T�Bo��@ѻ=�/�<8���}"�r��Kbw��NyC�CԬ�[�������>,�j ������(�d�s1�Hf=���[>ߞ4��N1���J�}��u] +T�����R=��^��4ODlo��������ֲ�1ێ��M;��W��Jaz	�蝁u	�[cn=^�^%F%֔|��}꘏���z>�6��*�| w���8�p��OӋ+�����l�˪CF5�T0ܭ���d�W:�����U�������1�^>����X�O��6e���xE����L�<9�]��.�	h�`��u��zq���u�(q7�X>9]����+���f!؟�ud���WfԚ���G�}���ý�;�X���C�ɁsҜg����� ��S��ô}�(��1�Q%d����t��Q9����� ]vH���3r�M�5e��,���"�IÛ��#�e	���Ѫ)������R �r$�n��"�|b�L{��y��kZj BX���u��ټ��X�9�~W�jI+I$�	$�I$�I$�I$�I�������9x��M���b[���P��\�V?[]��2�I���;0�ފ���0�=�]��v_�� "�����<y+��U��q]���6\]��U�H��E�v�}7Q�k/����� ms[��;������@�Zx�Uy���Ȟ�'���?uzr�]� fw�
�;����W��Q9� %t�Nt3[HDP�OLg����zCHݼ��d��
���&�������ݹu���>9�㖼m�c��,�9m��ډ�Ũ)�z f����X\����wM�d������u�ʂ�jd9������ܔ&׸O�5^� &��_@O$A��2]i20��Q�d	>ZU;�W��1���.z&� ��`~t��O�`H�s��Y�)}C�M�O'�I�_ׁ���(WR,�I��< Ǘ����<M�j��*����~�5#ҫ̙�ʾ��c.�L�%껨DI�c5����I�xGB�h',���>�����\���yN��T�\�c�+�9��pmnb7-��e�Ɖ�`�\���i\���*�� �X���Q%̼��o$�I$�I$�I$�I$�I$�I/����hD���g߂X��Yڗ��@�ތ��Vs40�Uv )��d�~����v��Zw8cr��e�\���ai&��S"�+�xo�W�wו�~�~�MA��۽��E��g�˷������ULfj"nn�Qэ���;$�5l
 7j'7�k����^������M�j&Z7S�r.0� �g�}nޔ��75�Z"�7Q�2�����u8;n����d����͟N)��nV�l�R(��^���Ep�n�4���
t��'�eOi���W�u�󭉧�A%�I m�L|泵���Ŏ���ks8��S�Erw�G����&W��;H�Ro�Z�!	�����no\��[�ʫ㚋�Mlq�l��Ne{ޠJ�x������N��� w���j�5�kN�^���'�~>��f���Z| �*�ǢL_�dA
w��3+t��.0͡W�u$�*T���*�E�-k&"$"�,���)�%�b
(�0�q-z���Cl�E�{i$��o6��[wy��r֭$�I$�I$�I$�I$�I$�V���QU313'y����O��Ml`��Y����%s��%�_�t�:�5�^>�W��Jx���7���λi�Hp�-b-�J$�6�4������_4js9��mE:�}�*3��]�t�+���>~��O�d�Il�jKd7�v��ymvуS8�ƋǕs�+������Mb{���F�����@�0BS/����//�'k���3}�/|��>�|����tď�M}��� � ��<��01�;�Oz;v{Cҙ�Qs��Yl���3K M�c�p}�n�~��:�lmR�T�w9;�<�\ �%�
u�zY��;�DF��=n+D<D�1�5� �λ�R��}�}��)Mfx��^ŋǮ�-�-����Q-��"@�zn� �⺧/��g{L!'z��laG2�z	ކ�:��6�=4}[z _{�M�cu)zز�&{�8�(58��sV>� hV#<Ll�s~�(3-^5�f"�w+9.�P;Q�M�Fά"��WXᴎ��y�n+�U����.��*I$�T�ZJ��(I* �$��JJ�%	%C���`_����~O��ء:��Z���f�+:��A��[�c���Kr�����[{q"3k���Ẇ�J� ���6YI���J|��rW�Q�ދ�/d�γ�lV��o��c��{����}K��3�ou��l�<�V�;3��oF��-+�]@ޚ����6x>�=:+�N}�4_�\��=L�8���9On%	�-Л��qZ��z���2Y'��'O!�ο/���8N��Q�T?��J����~�L��qt��ǵ/Ò�Ƅ�1���|wG�`��]��4�m�nB�=-PM�<�-���B�"�7�=�(��m{Y{
�q�s�f��/�5�w^H���g�y��x�33�>{��A�q#��mT��ɂe���7��c�H�HR��T��V%P�Ȫ��(F6	+RS����$�DA\UT��L����6���2"�a�4ۈ2�$�a�>Ed��C_	T�UQꦪJ�P�I$���P�T�������/�ء&d��%A��͙��_�$h?�=����CC�9����n�tl��s��2Q�_�)^c=���5�:חl���t�!2�7���f������vI�qE���z��Ѿ�CFD���������9_���6�ic���9�!Qby�0��s�*��
�R2$ש�l)k����]\�Gk�x��E'��y���w�Gw3Y{&���b����Vou�\]�����g���dU�6��r��ʦ7Ff��^b���ȅQ�/���L-�b�b���V�H�m9W����Y[�c1�Ăe�LD�����6�7Ճ��_��Pݎ��ʙf=�܃2����q�w��鏯�_�9�"��V�mP�Bǚ����[�Mn�{�m�L;8h��eH�yL�*&'Er��%�֭�Y���m�Z�]�ôEh+�/��ﶾ�(I*JJ�����$�%	%IBI$�U�rN/�^��w7Zuued5)7*
�G����z}���C��v1l����&���c3xQڷ��E
�$���2�\z�s���փ����%���B��!
����kB�N�2{jvRڧ>x����>���MϢ�5�F������]�؄�ˣSFg1�}Ҍ�j�k����s���Əw�����|U����|}��O"ni��OVA�G�/A����!Y`ɉI]-o����j�c�rQ��v���z{+s�Qت�!���j �u�.�3]��u���A����3R���s��ㆮ��$���}��jѥ����)!�.af-����}{�N��_�T���<Y`���qU�`�ŵjԶ�aX$��0�~�Bw�0��B�1Ib�����Z��e�)�6]!cE��դ�ߜ&�5��.JȲq�3��``��012�U� ��%d	�W�P�s��h�;j�D!�V��QeE(��(�KhYEQTR���QJ)E�X[F�1YE�YEEQe��Yd)EJ,��)E�YE(��(R�(�)E�UQJ)E)[$�k��L��5�t����L_2��7U�"s�/�"��%f���u�Z$J�Ũ�ػ�^M��ݎ��]wߙɏ��y�����}Ubm&�O��%5у�Di����H�s3:��0�,s�o,[Xݽ��Jɓ��jV�WBl��"e�q��i�Lz�d]��Rɺ�H+󅐶����t�����d����E�j:i�v48����'�y<�If��y�%���"I�O�#��'��X�(�պ�,���S���Š2k�<�B��BB]	�C!=������t �y�I1��o5�}~ӻ�m���_��1�V�9��>YO�!
��ى�X�ۛFFՋ�4�ZC�CH�BB�]2M*)�0�	jDq3��[)�12��ч+#1�W���Yf��m�i��5tk�C�bF���J�F(��\�XJQ�|��Ïq<\�^�~���?"5�3U��z�lG��&�R��Cb�az��z����f��}���8�'�+�ɤ�02*��k Cb�s$s*c�O17�S�e�CƻSn�29ædd�8�|���/6����o=��6y�?i�;���v�v��7}����8px<�$��q�'�QR�����JS��;u\MNU_�0:}g��0Y�H��[$��+'��$��OċR��vG��-�;�r��nʋ���I�U$Īp���D6M���Rرd�31��$���em��!�,MX�T�����n4oɞug8Xٖ�a*?��\$�M�T�A���L�������F�8J[���qlI$I.��:f��q3A��T	�c����ѭ�,)ӹ�.:N����>��jڛ��߹<C`��%��Ӏt.e�y=�L����	�vq���S�Ě�D�@��<����.=ǁ"*����^W��J�_�1�����8ş$I �O~�g��/��C�N���~���v��w�e�T|���7�p��7B��z�ZeVK��_'_�C�7����>{�a�0N
Z����爯�v��beɣ�[z�{λ"I^5�b5غb�F^U0hu��njXqS�s
�oq��kН��S��	�2�p�l��Ū4C�V}�U����9�c�Ĳ� z�=�PO8�2�S�����9܌�=]�	>������ju7��	���T$�fP�4��)y��!����nH�㙨WN��rE8P�0��!