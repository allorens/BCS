BZh91AY&SY�o�ֵ߀`q���#� ?���b@�� 7�                        �            )B�PH()!@PH���� @T�
�*ER��@R@��B�� IDJ�$E*P�PPT��NZP�� Q 	QJ*��R�DPP$	*@
 (��$�J�%QD�J�P�$��T(��B�V`� R>   1� PE
1P�� ��!E[ hQ�
V����P j�
� ( )J %%)$�   3]*(U*�U*�2��(V�0 )�eP�T)�SR��@Z��
�3UD��Lj�( 4�(�3%R��*�H��   �(U(�i-@�PR���@l� J�I���!�P�P�Z� dY� T�`4R�R��B��QR�E)**���  nP
���@@m����0�@�SQJ����P&�P�	�` ���(�PJA@	��RW   ;�j)TP$� R�fS(�*����¨�1B�he*�mXU
�b�H�`P�M*(��
T�"��   c
*�]�XEB�R1� U�0(PP��R�,�� �3
 ����  ��T
(YS 
�)J	 �Q�  u ��;(���M�XP0@�6�`Q@�V�(�V�@( �° 
UUTL
*�
H	$��  ;UUJ�F��T[T�ZUU*�	��%U`��*�j&UY�R��R�5
��3)�URJ�T��J���T"�  ۬T�(���T"M$��ĵP�"�e���UZ�UQ*��-��%S*�"� ��J(
UA!�)@)!R�U%8  ��J���h�Q&j�hU��@����S �
�cSJ@d�T�UcKUQB�lUUJ�x�    S�	�T�P 4   h S����Tڇ� Fi�!�i�L� `�  O��IR� �    &�"&j��z�e6#P����jzj	OԤ�T��54@�  �i���[������_�����!D�IL�5i<R�v����\�o�;���:�~ν�B}�@��QB�"x7�C��e��������>�wJ�B�����=���c���U��H!������{���X��ʏ}�s���XUvX�XG��W["_(qd�,QŒ8���
��P��+�Ŋ8�N,�\YC�*8�K�:�qaMY)Őq`��\X���S�(�;)U9�
��".v*E����E8�J�J�Չ�T��*.,�W+�*)qe��Hqd�u�*��*#�$�qaD�ȜX��$qb�N,\YJ��*�ȫ�qaXS� ��}Y����{&r9X$Yo��(~z�+�n���f�F��Z�O�V^3��j��\��׆�"��_�h�o:I���,�w7�7n�7ӷ%��Cȋ��'^�C�f���6�38�݉�����;+�\���8"��z5U���sJQ��q��A�v!{�o"��#�FU	7v^��<����vQ�l�Z;�n����D�MBOľ]���:C�B�uM�(v�s���OZkVlΆgf��7�W^Ȩ����;&,J=��.�X7��-��5H��Z����;;d��<���9!R��T�5=�&ǀ�
�Gj����C���.G[������pn�N���a��3mz�m�F���+*`=�1h��ɇT\�y5��n]��ի��Xw�M�}�SӇS1dZ��NӺlռ�z�}Z	5����f�������9��Onȡ�ɹqdK�5����Y�[�c6���fu�W#��s�9Jq�ފ��P�pq]�&g7�QX���r�!���n,V;V_��G'^.9�s�^]㶻���#�5є���^l�S�L�{2օʽ���kB�	��	�&v7�8;�WO0φaW��Ѭ:�$n��l���\@���V�u�"����1tɻ��7CM�,���PF��%u��Q,���,�N׎�8���gm�9�]�)
ؔ�Q�����Mwi��c��ȱ�|U�z;������׀��>ח6MM�ћ5Ѳ��*'�=n�p�	�{v˒��7��\��p+����j��/��M���V~t�ػ����5������81>!��镍.LشLV��	w.��(u�=�)�e��R�>D3��[��>#R���C���S�[
�8\�	_�-��Ypd��pN�e�MȞ��B5c����&=������C�����m��{����Q��#ӷavW@fݒB�g�WM�wv��f��Ȋ�C�@�o؆��{9�0�އ'Nͽ��!bq�ʑj^�Z�����$�P0Y�6�_�3�Έv����ji� L|�5ݷ�kBZ���[��`���B�]B������&�j�Jj�w�ku�����(��e�+�H�n���wO�H7$��Sv��^�}�:>�̩ۛ �\\w��Aۚ�UDh��L��T
1�X�q��vw�,ዖ�!�˦t��ވ.�Aq��3�#q�7{]��eN�:�f��z�Q����V$�J�vI���G�##�V�|�n�j�sl�<�t��Ν�*���n7���c8g#{���V�S��9OG���_�-�w�/ZrCrb��n�C���:[�4Γ�>s$�7f���V����I�L�Φ#jeX܈�β��n�;��wu��n�	A�s�ǅ���0��3]�#����ޞA5�2f餞��E=V�K��9h}�Qد��;Jר����[;� ;6���e�G:��:�VM:��vN���y�K�t6������ѝ���E����+qND"�8)ǧ ��C�gC��#�J���['dD�W	!ǕZmG��pȊ|�)�S.�\4MV.4B��#��pp��E�2��y�ڡ�]�LA�� ���/a웸#��3L����招�upT�d��#ېa�c��F�;O6l���c�fp���Ni}�r�x�K�d���`OD=�y�p�v�7퍄u2�ݥ���OS�x]t=��n���v3{;i�q9�%��96�M��=�Yư����A�D��bjS܈�#N�jHv	�ܽ�U�:R�S;z�]�͙�:�ٺo6��rd{�jV'�j��b�ؖ���=w�F��,���<�f��N��wh�����]۸�J�fȪ��,�h����S��а:ɜ5��aՓ8�n�hn�p��g'yk�Ĳ��t2�·FH=����z��Q���7�(��OoU*�njf�͋gǓ��i=�[h�Vb\e�S�<�ü���S�40�q�]��<"��Z�����G��v.���;>�XtYr�Uu	��zv�f�&�rbǥ�<��E���rqP�ӒqM���35��I���5]=�i�mi�2uXov�<��B��l���#�1Sj�1�sk���_g'ݐ��gmW	�¸�[E���;�𸬛B��K:�.�`n����� ,t�u��!-���f��!\g�!�d8q���e$+�b��b88k�E�e�@qr�¡���ثY;w����	�����{�g=�դF��h���qW���Z[�t�\&n�6�Z't ���3C� 5k/
C9�s�G*��$f��77y;�ZX�"�h��p��{m�ٽ���;���u+��*,y&�Q���aN�o9ǩ���FFGd�$��ThC��[+�i��K ��]fMP���.��R��V(�7(k��>{3p��eY�����'f�9ŀ`hݍ��@=L��pr��*61��w;�Sg1��a���
�T�N��˫8h�5M��`�4�JӸ!E��k������OLh������L�L���ӹJHt7Y\����>�R'M9{5��	鷳kc���<\��b��슀��i6��(XЍ�$rb��ΩR�xu��;��n��mĈ�wg�wNލI	�OYՓ7�q�.��A.�Ѕ�0;�٭���`��J�4�
&*:a �3T��G�$�r�z�Rs]���+9փ�� D��=��Cu.�委��k�Ɨ����s�)�i�*O&�u��k�zX��3�
����3t�Y��@CY����8�#"2�+u�՘��HfU�l�ޙ���z��^J��y3r3�QÈ0\�^$:k��U�f�i��4�n�&BQ�SN0Zk��۫B$��;�u�󓽣P5����\z�����ގ�B�r_N]'72-�g�b��N#�v��f����Z���ݤ�Hb�`����yf���q7Ԙ���ڸ��b3�͹W���6d)�B�;�w���^�t�q�Q��,:�,����(Cx��fЄ;���I�2`u�Y˻(o,a��܆S�:��!w��=�o��ŷ{_=|f�?	��/`�Q�1t���S�s�~������蝻V����5��q�Z�e�^\�)C�P���g�wx�9���Gqc�欰򝜲�Xj���H{H���W]��}��8�q���	>��cX� {��Y;�"́�91�_u����]b���	�>��x����R4�O�1��Ԙ"z��f��Y(�nYX���G��}'N��9�����k3&�YsUCk�D�t92��B��
H��+���^�s�g:t��}����8�'�����$zլ���������?:<��M]
�!��\]�kB٭6��ˈ]��nrQ�;�`�N��n�������
�Bd������hI�e�Έg>"��,T�=��ƧH�GCخ����v��6�+���s�����-�����κֹ��ƹFk�	k��v@��/�c��O��D���|���]�7S���3�X��b�Fi�Q!"�թ��j�����U_!n���<V��]�{0ooL��2a�D�ȴ�7�n>v��,�r4��H��] ���w��yf��׻PԸ���=�����F8�"n�=���;-������ ���le9_M�v43�t^��� X���{��#œ$�0�xp*��<[�⣡&e��5*v�|hP��'h���>Z:`K_�l���BB��5VΝM] ;K�9O_*���1@D��*z�Di�߹�rv�B�C��jX��dH%y�gQ ��4��ٱs���Iۿ�gi����0r;k�oZ�kb}d��<�ϯ>\Y~V�kY6N���zxotn#�Z�qq�6�ὐޞDvAP���!�ᕜ�`&��^��՛�a�
���At��VqԬy���ңТ룷%dX3iu�z��� mٛ�+��!|EHy'k0�&Q��9�BY�+.�:N�k�ww5�������ɃsRzP3#ӀH~�ɾ+����ւ(�^���+ݝ����#�R��x��Ǟ�o˖s��Zv��Ӎ���glѰ��_/v45pd��%�w��x5و;�����nǳv��8q��.����A�	�E��B5�^,-S�c���ع�[��_mʷl,��W������m�p��ˑܰ�q�6p�OY�(�L$!Y
��u9D�F�s&��$w�-�ݦ�5j��\�"��-�s^����#�7�\5����f#�c�d��7J�7]�ʇt�yW��;�y�gkŜVv�.��Y�2��AE����t����hph�v+p���/�%t�vQZ_i����/���ik'Si�31y&2`�)�h��e�Z8��x�&o.��f��	�y`��r)���
Є�n^�m�`� `,��@�Z�宀z��q�L��F����Bu�-\O^)�t͓���943�/��-�'i��L<:�4���!�	����2lY�gB��~]��*��u;�=v^l�q��n��#׶��ص6�)ݠ��7)W��ő��ץ젎gY O�ކ9$	�'j�t�A쬨q	ܤc^I�oh��Rd��Qn-�޳|WO�z�)���4�PL� 
kԩ\0�fN�`X�n�/{7�2wA�+�]���������Q����i�c;f���Z2�b��d,�˰��ȹ]y�s���'�N�ɐv��6V��;�^��Nn���n#ݻ le��@Z�Y�����!�A˟h��Ȩ#�N_3��-� ����A/�Ã��j"n������Ѓ�)&��6�ez5E׶�γ&<:�Ӭ�H���iH{�`L�{��9��2VB֔�8խ���s�ak�C>�w�۽�w!B>iӃ7�T0�;ur�Aeǖ�Ih7�t�Vm�0����nn��S�w�:F���{g(�j�>��\�`O�7�I�}N�"��1E���M���D�q ��R�W8�v�|a<�xpt����~lœ��݉���XP{wP��e璬����M�t����!��ٱ4��� �HgN����믙���]^��|�����Q�u�	)Z�KC8wcf�H��R�F,�vW��v)F�P�0�(���e�C�r�a�3��Jk]sGRq�ѭ���x�Bg�s������L|H5�-�"\�E*g!�ė�ݺs@׏=1��ݼ����Ĕ3�$�06�W$��	�ݖ�T�s�·\a��"���*3\]�f���s����;/3��s�U3T	2c���ϒ�ڝH�05Λ�r�2�}�{
�0���օY���ᝥ�o)�)�kR��,#MYd�=��]�=P	�U8���N�F�M�@3O-{�M���⦘�;wH�E��we{A}��H��t\Nh����C��������tsDۄ�K�1�Cѻ����0
�(���PӉ����;%�^7�D�)E�cb����~Vɯ���t������h8����u��ݦr��}�{�O�|fDj���:��fwh}�V��5\����:K��5�����;�R3Vp�s5vZ��?��Nʆ�E�eK`�cc �w�����`ֺᏒ��v-u)�5cٽ��Ψu��Փ�� ���A�A���0Q����ĵ�nu�.\�	�$����7�h�ǫvT�0�ܱ���f�]�;-�ۖ1�(��v�- ��E�a[��myy]���lb�����L�}��&�.d� ք�I��΃;AV��jC�B����GCv(�ګ���T�u�o^�m�x�c�ѝyq�;CĆ�$��p�K�f�5�+�XU\���Ε�D�y�"M���v�G9��[�56������	��yq戍)�m�Щʖh�)[���;76ُ.·Q�f���۷�$v��zBh��G�ɒ�����b��Q��/��ksE�>����jKK�8�j��Ö�V�����/Cyz��͐��&o6d��n=��]����;Zo{�%,�8�)QJ�����}rW[����kۛȼE���)A�Їh8˷�7g4�(-�H�����A2 ޘ�C�tM�EEʵǙl�)�RduV�V�c[�nԻR��S��im�������&s����5��pD��0��8b��u��1�,�vC�Dz���r4��>�X ��K���J2#���tBb���:��IX�����y^���Q�u��)��Y�*�{�j�4ӽC���t�Wtū�`}W˛�]����(���h��񁷬�l�ۜ(r�"�Fo\�l��!E���N'h���|���w3�p�J���w��7Jawsu&�UI�L�l�>ƺ|(-"�
Â���[{�އ�8��.��]7��&����	.��1-á�"s9�kΘF�,�öFƻ���[�������Á�.Sin��i��H-��Ł����N-�#�X�/u��Fv7J؆oB�-��Y�*:�k��T=�*�w9b_>�J���>���5�:�ֶ�H�ů������<���'׎�p�!�"'e췪�mm.�e��l40�-��'��t�7n��S���'T8
�B���D�t
{MG�����+S�k&�W����ؘVkg"��f�v�R;�y�ʁz�ڙ�8�%*��%�,�wWar<ԁӬ]�"RK9�4&BWsaU��$Q�����ٍ�}���'��ֿw���Χ��i���	�s���ЀP�7r��F65��ԕ���)��:�k3*�]܇��Q�j�J5Ck;	YuDaR����i��N�u12]�Q)槚-5��W7��j�xh�w��v�2'O�52�cݾ(�n���<���^^�m*Sy�)��q�e�ui�E�����4�8��4�dҽ��:�ܵ����X"�Z�̹m)N븪h�T2����0�MK��$��_�@8cs'���ے�p/-0앥9y�0HߝQ�"�&n7)iz #����j���L�l�~A)���=ہ�+�"M�]۩���'gM�Tނ=�o��}�w{'M��:[�8�'�,�z�j�@��_o�h�V�2%C�ߝ�,ܽ�AD���R��^�6ܥ�:����rh_;�9�g�\�Ƽ�E���+q�w�֫�mç��k�+��	r{d��|����(��8�w�[�P�o��v#m�&����z��K�{���!G;��)n�"wU������ҽ4�K�M�j��X�߲ȍVS�7����<�޷�zk>�ȼ��S'�`�<%��A��x�n+�P�	��/f�E���y7���Bn�6.�soL^��\X}�x{��|�y;㦎���4f��������\@�Mrj�9�틆p�92�SA�����=�'6B�˰\�A�Ge���]ث19�̫(���^pଖܷ�L�7ݷ��7.^������X���ֶ���#;`�C�0�Uu-ӤŸ̲n	�bWY�N��$�r���3��'�.�l�*�^n����7;Ƞ�N��v�^TY+B��7˞[JL��1�nJe&����>0�,ذ��>���vJ'x�|=V�}�9���@�(Џ��g���{���3������Lװ�I�Z������!lV�0��1nHZoU2`D��@\��X�o�������$��l�j$- �|�����v����7;D���[Y�����1RCF�L�yN��l噛(��S�ݡ�
 55�D�+ػ��Vsm�ż sG���]�=���&#��7�s;2�jڏ}
�WI�@���ݾ���4@�`�a�i�)����:B��s�/��Qm�L����SZ�W��^m����\i��_�\<����&�bnl�4���Dx3�	����;�ѻ�^x��;���G�GA;�J�'���S�|�/h 4g��r�u��y(���^y��X�ٜ�ri��݇Y�ؓlo�WO9V����XYs���?@74��욆84���f�)�7�Zi�\�N'˥�,�FN��]�`�-^͸%�J�G�B�O7�t�ݏ�wp��-�� �p�.�8�7���#D
.��w��}�0^k�F���=�<\/��,e.`wEGG��\�G;��H��馤�����!"E��vf���[�[n.��%a,wZ����:���ʛ[y�2c�TM��A�r�����un,��p�3����&H��{�-+#XM��2M���r�*��/��Ʉ���w$��w���z�F�����`�[�&�&IAΫ��O��$L;�CW�1�R����~����{���A��i�<`�0e�	~�A���2�⌙ז%����A�6K��>H��&L�4�������)e��}��f:���O]��J�gZ��f`�ŉX{hC�^����;��;==#3���8e�7bz������ё����/�r`������8Q6�ټ7�i�t�a1n�^��;2d}8�B֋*׿X77�y\��{[O�^z�l�����M�
tX�K�3W��T�5,U^�!L�r��ؖS����5�z��,I�0��t��gn���Ʒ7Ϧ�x��=�������v��L c^��1�|������cZƉ��t|��RA�'�IR�E�����Z�q�щg����1��X�o������k~F׃f����\as���d��wgIx\P-�V�1�]�#��#|�/�
rD���r��x8b��`�W�G�p�6`�
��3����W�>�X������cY�`�7�q��(�p�UP�������<O^!���o���xH���Ȓ�#^xz��u͠���}����9��8
�X�hn���=824:��=�����t�p���7;���K��Q8�K�Av����*r�ۿX3� ��#�r���Y3���o3�s�����!�czg�(����N��U�.�Yw�0��d���F�ET� ��_�Yp2�'����{���ȞC�&��-�|9>�p��7���O�5�ʾf�G��`۾��4c%�}���xe�2gi��Ǿ�}��9ڤ�˺8#ŕ�{����>9��4Һ�S�g�Nʇ>�ye�Ć?x��5���?n䙟�D���@YL`���lKy��n�0��Ǳ�z;d�Y�'0	�Ê�-AU���*l���黊��c9<�ۈJ�W��+;X�%�P�r��F�9e�J���eUάro��_��YQ�@�zE�YwH�T�w,r�����TұY46R	Wbt��l�r�&lԬ@�����{��|#4,�Yژg���p�(+57VV�+<˩��ڼpaw��4�n�7м}�A��ǋ�#ii�sD�����J���8�~>v�q��#��V���F򛲭qj�h8:w�j��G��S���/l��Hœ��.{�%{�t�t;�i �9
�o-U�I�H�o�YqN#H�M�59�.	��1~m<����nza^/"���f�m��D�b򠋳[9p�p���޸/2tE����3��&2^�ݫ�I�s�(��K�k���OVo���Qpc���F�N��5�|9�������d����	�OOۡ!���<��)<�WcΝ e�^�����8\�=�&p:�V�m���/r���1�23C�͝��.��������:ن<��F\H�/Zo �*�ŁF�V�T�iQbVCGOh��=�����p#�,�w6�mS��,\�Q��L��[)1�}-?y��!VB��.�XI$��m�E�����;G��_��w���� �6�B�$��|['��a����`ﷳ��:�x��,7��3����E�8�r#�0sVY�}}�O�7��՚�eUI�X�[� �E�\+��U���BJ�bؤCȘ׌+�t�����B�02�7�4�w�`���.�Kr��2�y�}5��X3�� ʜ}�9��>���}�<�͇�[��� bȳf1*1�Υ%ɬ�uU"Y��8���ҟmq����pk��;s�AB�=$�N,ٞ�b��d��Z����r_Y�� ��T�Ҽ^�3�d;}`��k4��{�)ly�QYF��OZ��8y)6��kv:���Ut�:y�Q�dg���=�y���mC��n���i >��a�]��A�	�E�zfN����@W�+~X�M��X�O�l��o��ꬴ��i�P�ʻ0�����sW��XYt0Aw{7���a3�2e\ƛG7O����I�>js�+p��.l#=�^���f׃��}4͕z��C"�czc�W5�S�Fr�ѥp怕>\���+R��:-?.׸��������
�M��F��\V��	y.E��k��������ޭL/�) ��p5SA�\���?{6d�L�Gok��}���C ����%3Dy���Od;��1/��^>�g��4<��o����i��Ŷ&<�H�����8/���q-��䜬��X��<��ܙ�?��=q�}�w9[���,��m"�e� Ӝ ^�<�m�1y�p(�Ŏ���/�k��kS�y'����`����gw�ax���m�ݔr���bX��w�Z��!(@E+���-Q.�Yӎ�� �-(OXpD��q���o��|͸֍���T�s�qg({�v�m�ٺm��{����%�M[��Fh�vo ߉rz�9���/N>ɻ��@���LwO//r���6"�Z�[��G��_C�B�zS1�l4��\��=��^+�yx.��t����c*�q���9t�!M�J�y�+l�e�&1��ꭩ�b��i���g;�R�~θ�
Hc�=<�<�Z�7ܙ�F��
��織�❫��KXbY�T�bs"�Э�yUt[{ώ�*�������#$Tq�b��t	�"7SKN5/n�UJ�Ԕ��Ei;�����
\��8������yECj˄l^�p6mU�7��V�<B���9h^D�ɣ,�v�2��z).t��$_$�o<��BU]S������n'�J�$������8��{⇆t���M���Q
K}pp=޲��A/?K�:}�]}sN��C�����]#y78�b��J`�l:���|�R[�L�c�;�zw���9�����ꆚ����\�Jdޘ������y�%��ڏ{
ឌ>�������!S���&mM:�76���O��v'o��s�\��[��tk���^�h�"��jP7$�^'��]�=��<�0�~Z#�c �'1ۢ�t<���].&��B�P)�����ᾊEϺ���C��K^�D9�w�=�V.X�����ٱ�|"������PM�m��yٽ��-n�5����ڴ�'|�V{BÃ�.�s���lOx�{�ho4"<��&�ϒg�Z l��D��S4����羶�R��(��5��7���OF�n����yt疼�{Z�s���臞�4z�R�[�q�z�S��NÓNw�y�Y�}����(��p]9�=���M	q��q�r��	��ѧ=��Ը��w{�y����]��X4	�SsV�K%���p��[��v�X��z��/�5�z��R3����M�o�v�Ge�.k��ro*)����Y/�n�7��N�#�J���V��ya�Ԡ�6.�<�Ѭ[f%\�(�V��8/*nX˝�ow.�7p��T�>7��Oq#�S���`ó�Z��K!��.N^�֦��kt�^P~r�1�z%N�pù1p���&�ɵl����ߋY�H<;�^��W��m�p��LY��+x��Y2j�t�+�x�ۻ� ���b=ݫ
�������{{�\AV)ɉ����3-d8.[��Ӹ��8�P#5������:�W���K�F�:��S�vnn����̊ʁ�r��V5��~���~�P|,����v͏�|@�j��e�Wj}2�U�I�z�īnnٛ�t��aa�Us���^��F^�r���pzť�~�ٔc��gMn�t��X�(é
�n�c\��M���G�έ�6�[xM6��� �h���oY#�zx���S�%�=Z�,پ]Ҽ]���{���ntm2�<����|/�Py��.l�:���m�us�6����
2�͇����y4����(Fc�]7c�RI �简ǖ�$[�d��y�x2����H�|}jۥ�J<��N�Iw�Q�R����
j�6By�2���!��rM;�4k%9ILY�6⤚s҂lUZqT�D�Y�ui��P��W�����X���ӸC�ǻ�`��Ӟ	�/d$��cq�^���K3�w�j;�xEu�B�I�2�6Q;L�$8�QJ611�^�=3��sŷw�}t�߸��3��'�oc��wq��<>~~�*�7��ݦ�r�7���J�}	��a:�7^�
N���d�;�/)�r�Z�Qct�y��.uI��v{�\���M^>�~�D�؝2��C���.Y�jR��ZÎӝ�I�Xvo%�;P��H'ְ&E�t�'t��t�f*bD��Qpoq�p6�.2ݶj�b�bm�}��:�?O��rs����s.8n���g'�ݺF�Æ�q�g+pn����`i̗�����pa�{�F{��7IEc��zGS�zyʻ<7/<���	m"�D�ڽ���ҵ��v��R;X�A���kA����i9<w� �ƳG���]��h���ͽ����w��c��)�&z$�~w�*q�Er��
�@�;��&���i(��2��=�_Y���{�@���?SRf�C��+<'}f�����w�o]: �7��[�p����p&9O)��x�/�<�kt�� ��i���2�K��VNK��I�մ &s��ܾ�{��{��伦E�<��'
ea�P��y�h,h]Ɉv�T�c5�˝�d��h�ۆE����/�vk�~�1�!��{{��>e�l�6f�9�*	i"���I��l:���1��x�,VVF��rj4��7ʋx"3u�nnS;�}'�g���~x2�3��$���{<2!V{,�m�C��-�Iؑ�m+n0���p*9��rjE���R��øt�t�[ܭ,lw��S�z$f읰}��[�uJ�4>>���c��tU�\�rz|�a�U�::�e�3��	�7�)�_���p���r�4uw����:T^��90�t��2�T���EX�@~���1yXw�_���@���v�}�G}��v��,��6��=��l��.�d�.�މr{$���)�O��s�N�V&���{.��=��,�-��V�Q�-8��y�=�^�A_/Lun�2f���P۲N�7%�v��f+�w������^�g���|�e���	�HL;�D(l$f��ʍ���ى�FP�j�]2�ՂY�8&��j�k�L�DG1���o�4[Z`�Q^Za࢒rg����ݗh�f�Ǯwr#�
�l�_{�w`�3�=��?h���H�w{}�m�����N��m���#\�=��w�u�B/f͞��Km�Y�k1�[�M��Sn&DNi�ˉe���8��6��N�=%�i����&v�~9��Q+'��m�V��Wb�q��e�u�k�:��A�o0�;/��XiԹ���6���-cP���U��M^����*M"��Y����;�д�^�(p�0g����\c�(����U�iC�MT���ch�\��
�8��g�|R�@B#�"/�xQ<Zc�Tj�3�(�c��_b���5�}����}�������ڤ�n�㻧(���U$�����[���^�/.[�����cg��u_�L>�,ag��j��N���(n�t�᳔����-/
�����3;��ˑzy��Nv���a��O�E����Ѽ�m���oˋ����݊R����QE�X�t\9���q!�</N[��p�;Y[Y�{�Q��=P�{hݯ/5��p2�m�;q��J�E����뻦@�>���7��r��X�>�HwL@�%"��Q�·�Xf s��<�:`k��=P��왪�����Ż�����}ݫ���V^ظyg��t6��p0�'�ox�"w�o��]�{l����w2��Hˍ	ݨ�ʖ�0�[/ .⡌�I�k=��p�S�ݙ��_H��y
��o��=k÷2����;���b�b]]`�.i�q%d3����S�C�����m��N�a���A�[8t^Й]�zIL�;ze�|0�<��yA��_(rz��أ��c.�:;=�$�w&���%=�\��L�QxM���-kZ�@�GϺX�����Y�끱���gm;��N�^�lL��(B���;��7�5̽���^��8��1?(�Ѧ� _�����͌�4#�V�1�J5��X}��v\{�~��o�����]���:#�Q��2pݡ�-l;\W*��wW���o�/��ɤ.f�+U���n�Z�F�_��xg��8��mu��#`�\�	>�@g�p�O#���nk�J'���A��#��O=��tfo_$n%{:cndXH�'0��U���w��!�i;��C.�W�Ƥt��q/~x�)�WX�=Pӱ��ٰ�ٲ�;���
3�A�Ysǵm�t 
8����(Ԃ�؍���w�l[�e�n�=�<��T(ەu;W�%��{:�W��}��a�+���[Eْݗ��|M>8xn{���F�K؎3���3�R�Y�X��<�fS�{���)ڵ]�.��|-���$cXi0?*#�������Ȩ-t�ՠ�דx�ӱ7��S�jnf�0��1f�������E�.$�ҕMPKv!�����
#{�����~]����4��y���8opÖX�N�i�Y���]�Y��3
^��$z�vQ��1��re����H���˳;x�>O������8У���x�L��BYe�:��lSť�/���B>�T��:s�i/Wn�Y���w��&�pY��ZOH¯$����������2��݅�.�)�1OS�v�Vyćr}���FMy�\9����;�� �,�q3��}2�Mj	Q�>��u>�׷Z����gm����sFw�c��:�.x�ԙE H�:J�x����z*�x�&4Й&%iz�/�)c{Dߌz6s�x�'���n�WSN�V�T��4�]9��N�e -��FlUl�2�c�t�{�Wd��9T�I����q��=L�;�[E�hâN��mm�F����i譩��j����@��Gx��joY�9�n����뼼3Z+�枽=�]I61U�`��ر:�n��'��w�f�\3�|m ��/zi�>Ow&�_`X.C��8O{�{��/yn�Z��UſD���:B��#C;�3�@p5�*Zo'��x,\3���[�7���ㅫ���{���NK���D*�im鑆3Le�����K��m��kg]��&+b��2��$dʌq�V��9����y�^ޝO��Xۦ�������#��#,�܃��_�Y��<j�����uL�l�<���e�5�*X���?�B�u�`E�ƁV��sV�@�&��W��{+uU��y�ӗ ���'�n�-�b`TJШ>�N�Al^��	�	egg��IS}�3ۈv,�uZ܍�=�tX�B
e�j".��3:f3�2�dK8AUf�{j4�ξ�GcbSۉ,���[q[>���#^�D^>�g���әe�ֈ$����Zn����l��������[�Mb����w�^1g��ϻ=7p���˂��X||�<oR�����1o�Ǘ��̎*���^=�3�a�Y�w�9n)�"}����T�'����rْ{���\��c�D^�19� Y�N�ciAK�H?[}���'$�eL��w'��� �����|����؀�����ͫ�pX�qe,;+��:.�CS��h0m�e�/K
�t�7�DCR�M:�i�ª�B�i�n�[�����WJ܍yz�>�ބϩ�S�1�Vk�M(���2VN�u������t{!�������YGۃ�s����N�ҿ2o��hWҡ�Ȍ�uE&�te��Z�⬘W��׼�"�����ekSXo�9�;���[4/.�{��
z&̛y;���9��9�%���=>���;�p�;ڹ�=|sɿ��d3���VnG7-z.�ޚ1n����	�NG�d�N�zq�R�oM�2��ʋ�v�/����M��[{�+-�9����n]�g�s��ǅ?xz1��ok���+����ƞ���|,���/aǧ+5�r���k^��oyB^7w�����|̾�f#79�����tY8@%���5�|���[�9o��~͋)	�ŎM�wR�6+�`pL2�Ơ�)l�X��qMMF^��������3r�`�O�'������N�Y[��{�r�\�6V\}˲�U,{�ַ�^�Lm!{N����gH��~�!�OB�����|�x�i�f�n�g�KЗة݀�a��᫯��|U�׽�Jg�����5z;�[؍86D���Fv����$��/^
��]#���6�J[KJ����bN͞�|i�;�H�.{�=zwa@=O!��R^]�DX3bFE�i]���w�:;.�0����G�7�`��&:k����Ä�M�y�5}u��r�f�\����b�>G6����7i�TJ24k�R�F��-ӆ��M5����ž�����U��OM���>Ҹ�_:��ʡK#�~��b+t�u�W�;�����=x
B������N�o���E˾^l6<J��x��2bsx���ʂ#�s!��j�����yR��pMj�TrR��/)�1	B0�-كݝG?_�Ҿ���>����Q�/�E�z�OO`�z��ɬ�7��I���^�2]}(�cSzo	���zf�F�[���Rh�	}�{���w��Zd��{��X������^bC�v�󼳨Ѻ0�'O{NVg�[=�iĆ�'�H�N�zw�^�X��};W��^+U`(lL�{�ۋ�}�G���IgRD�{؛YJg�<q^��wJ�.yA,5\��=�`	���죅b�"̛pN�d�cM7�:NYy.�E��u�;�7�/b��bf�`���չ�X~?]��w{��+��țY3M�����a�j���Y���P͔��� �hw3O�9���u��><.H�TGH}�xo�����ۑ���5�6�<8.�
�Vt�n���Eۏ��h����u�C��݂[�(Fzj��z��dgGz��g�2��Kj>�^/\�1oX�^�^��4f��c=݇����L-�t���1�Svt�Z";���^�[�Z8Tʷi8^ܬ33v��K�Kgw��։��w���k<�Mʆ)�z�^��E�s���=�{}h�短,��i�������4��Q�B.87��.O�cV�B��D��s����E㓞�#뎟)�4��O"�QVԹݸ��y�śQ���z��8��/y�$�o��H�Mg���2p���%k�ق&�*0\Sx�*u��Ш�و�^xU/=��ׄ���4F��}�^;��(s�����3�б'�"�\۠G�%�F�����P����}�-+
'�u�3{�. \R��6)8ͼ�j��sNۋ�����`����J�Ɋɲ��M�l5YKE��3�"�P���s~�-������:gS{����K����{7���8�#k�(]��ˠYԚu���)ڍ	�;p	�B�2 ּ����{Z��U�*/)����B�v�b�l�]|ѾՃ�r{�=�	ov�#�L����s�ZY�<Wg�ys�Ӟ�|�~>�g�,~��l}��#}AGn��K]\ۺ���J��$�Ê��S��`����[wPsS��N�^�GZ�X��eI[Zk	��P 7�Z��WC��� ���&�=A��s{tc��\�{�iK��5-$x��O)Mّ)=�$NQ��f�A��6q���%����v���:�a�-�{;u��m�N������ѣ�tta�c�h��q{�-ד� v��ڴ��^6oG�{�E�Ռ�&����
k|�*R�AY�Fi�v��ѹ�z<����p<	m���_�<��hP�����Ŭ��+�v�T����TIK�ơ��h�S��l,M�s��x]��$��;���#�� �i�n������R� .v�V�,��N2^����a<�ˣ�e��;����＄q��'�wo�ޠF t��;�)�i�������/(F!;!�(�o��/Zh��u���ִjgXN(S�����{��(F��!��/GY^�ʑ��h,_e�󢑯'������v�1�[5q���1٭DZ,E;������8.Œ%C�_�ϩ4�CAM����Kƹ7���K	��P�隃�e����M���u��Ψq�H49����w���9=�،�L~����aB+������E<�a*�B��ȗX&-&��`�[�{���ș�Om��[�����=�0��)�{�Z��>2rN��K��O!; H�(�;�D�8� ��wn�Fì�,�a:e:k'T��^�����I�UZ�ɒ�1ZҎ��F]����EyG������B�P�o�^���=�NFqu�;�+��YƮ��l��ru���rV��n��!�&�5����hX���:;h]S�|��O�W5>>�_���Z�v8�kX/;#��
{���;��G��J�����zGz�g�'��j�T�{�Wx��Z����`e$C7w([��`�.���훬�vmA�Oc%:��r�`��m�b)���[:>Ώ́ ~�]��y�S��`S�5�տ�U� &���gwk��ÕXhc_��6gM���S���[c7gCz�Ԍ5+o�o2 9�����Jt���n�vׯ�����N�ؕX�ΗϽ��$��Ts 鶞��s�oc^�C��.9��"�����:A,��t�����?iM\QI���: �c2�h�DTR����G��Է4����L���ۘ^�i�����{d��:eF'�9��n�������oOw�-�^��U��o�Í],Q��W=�=�/�w�
Z�b��DC�#*����`5a-�R�o��,�6�.L�B��e����Mqp&HZPq�ء4�7P�NQ�RE�	�7�E%Wkf����xu�=��E|[�h6u�+ݖxqk�����#����2k��û�M���ģ�Q�w�XM�&��8�냯rNUƒ^B��3Y�r��o3&C��zF�Pe˻9G�<�D��ק����$;������q���U��:�����"6�t��ybp�I��a�WX��ÆF�4��y�	�4�����z���${�!`�������
��9g^�H�Z�����P��i�ŕ0j�A�b�R�HQrŲ�3��cj���0v���VĒ�r���ۛBq������-�V+5TG<��!]r��^)�5^ܓ�#OmP�U9�N�S��q��w����2��aw���t���V"�2��H�5�ୢH@U�0�S'ޞ���=w�!�7�Fݢ�锝/�ypcټ�w
��Y�l��~�v����n��gwՇ\����oM�Fon��4U[��X����{��>�Oq�Ru B�藶�;���7�SɅNmg<�>"<�x6��N�g k�Ww��Z�,�)�ҧZbfjT(S�pcʉf)^H�]��*������3|Z�L'/Z=�$�5ts,�v3X��m��s9�Q�;.�{�v�.��#���X�6)��u��o��^�����|�c��iv��I��燴;#L(���`�y5�7�.2����x2D{��+�3|��Ŕb� ���rFk�u���I[�D��p��{�p�~�L��P�f��[��L�,��֓"\;�=���ܳ�r�g�u�y��D0�/�2v���Ԉ�T�������fkvĦ��i=̭���M;�b�7/a�B�P�.��@��RY���<��5'���b�O����{۹=���8hE�L�ٶ�ek�ޛssH�|��H�}�&L&g�kS&"�Eտx����z��$a+v�����ĳ:	�&]Ňޫv��f�xm�Q"��'�G!��e?v{�.$�b~UOe��Vq�,Es�����>'=���l6�7�2�>���b�__z�z88�<i�74����W�������|{NA�|NsE�\�c�a~�݃�C�^�)��lR�u���(Qj�K��}g�����' �O��P��8
m�\�Џ������%Sp��AN�#A
�4�K��N'w�G=�����ei��[�C#�l=���Nϐ�Ku�uy�z�C�`�w���&sa��յ�;[������ldܙ�l~67�����M��]�r.��|N<�������_3;����4���>��u����Ɨ�(�7@{�5��e8��J-������|�z�I���}�@������:�=Hta#�}�x��ywM�&��.b�=a���[rcl5{ڷ��O>�#49{X�Qgx�_�"�g��_��ۻ�g�>���8$�I��h�Fz��$[[�@Gx�*�R�S�s��W�ʝ���&>�⦙�[�7sTi��Eo/ vF�8m�6E2{O����Y������i�L>�jKܼL$�Œ�}���l�2f���Cc2�#����iNӬQ9�sE5�xc^<�/q����C�u�]E���7���&R�r�L�h����xM�z����Ǿ��x8�ti݃s:�Hʉʱ��1H���m>νu�K�.����os�ח-�3����!{+�������?��x/+���7���^5�Z��Νv���n;3�~�9鏽}7�9,���.�G�7��}���x͍L������Q�uͧ��k�<���u5��d�n	�b�v����{v@�W��jg�MzQ^�Qo��v{	���m�tzՊ�-�=���]��M�_�j1�b~i�7��ť��t*uU9(�����k�A���}�}�,3]"�Ç:!�W9.]�pF��Pe�$�N�U�	i
s|F�G���_�Of��b��#�&��(/��D�2.U[m0�[$��Ǽrlچt�4���ē�:'oQi'��᲍X�y��,���q=\=���ӽ��P8��a�{�̞���.��3n���ñ})E>���Pb�������)�>�=���}$�wBy�[Ngyʑ�9�¯48C���|�վ��=A��x��6e��������wl��z�܍4��w��e��k�㹨�e!��9���{�=p3���w�y�8!?O}�Z���Y�T.�׽�����Ӵ`ښ;�x��/:#t��gf3���rp�-��>��+��S��2{oc�n�B�r�n��4c���υ�rI��u(u����E�7��w@�X�0&i���F�{��;�פ���1�=��>���*p}�7��DHj�wuV��k�3�p;�
lR;	�Y�f�LV�vZ��e�H�Q��p�E�H�;'ch�`��1k{X�05��g�k�S~T�8�g:N۷��e�����8��s�_4�<Ѷ[v�4Qm�ȧ!�q�5�m���#4cn�6ݜ�˽���M�[n���I[ZN��������T�"�ɚY���I���n��n��N�rtr�;[q$�6����&�ac6�e���k;a�v=kB�[MX�m(K�k�Bt��=5x�&�i:�vdp�ke��������ۤ#����XYm�#��E惇##r��f��oo�Y˽�N�t ����5���X��|�|ϳgf
I;��P֚����������֑Ç��洞՝�9�w��i�f֝+��r����\^կ-���Ȝs�n�c�d��(H��p��Z�m��
=��Fݻ�2)+��28'�Q�q'<��rPBM�8��V��	��ŷy�yݶ�5��ɘ0]s��@��A�/���O2��;9���{�49��i����V�vn�5s��o�:��Y��|��>k�����,N��)d�D+b�PG�E��p�p��mNAB�����pt:��C&�7��ʉ���na���P�ᴧ����Ȏ��|��4N��t9��\��m��.��
{��] M�8�A��o��C�P���wewv�Dr̰��K���"��b�m@����t�Dێ�g�3��v��ί�{W`Oy������N�w����:�'v�A�Qp�OrB�����sS6����j���ƹƂ]��A�}�m�.�CX�*LmttQ�,�h����ʵ��I�L�;��/mw���3{�g�o-|�.���b��70��/s��s@Y	��p����$�S�,w�1�������F�]{�dpՐ�b��JO}Y�c�wR���r�T�I�oD�g ����u���.��/����&��&{d%�o�0���`�g�-�}�9X�݆a�A�Ya�}�y/m���H�Xs/e�� ��k&��;p����f���}!��ɧ���1�6�a�i�[�� ~t�D���Շ�|�~�����ƺfŐv��k�X�n�_�\���f�cˡ�2݇S��6�
T���^s)
��c,���{���,�S�v�x��x�'�79��X���"	�qsNcF��Ӑ��۽� ��`8[�7w�<�Ļ�s�� �w��.�"��Q����U�N��}�Ƴ�}��zsulƙ�[棺'�>��<����9�g �k�y��յ��bI_5tD�~�_lٟI"㝧T%�b*����X,�kj���,h��g���]�3����w18�1�R�wU�f]r%�nD��ɨq��'+A^K��>�o �ҥ�%q�	�i'f���'7�6�Dh���]�t8qC����7S�؝ǲ$RZ� �,�wwgm��� b��͚�|f�7ݟ!.�/J��Py�]���%.��v�2�،�yWR\�ϳk��*��8]
�]��Sg,���wt���d.�t���U�r���*ǑŬ��ȉo�͋o�)�
���;�9�W#j=��Jcݚ:+��o��F�X���3q��g��܋@��:g���y���C�=��e7���>�19�\�h@��Y8�|��&uuUᮤQ���r�yR��jZ�ov�aV���zf\�\����3ED8��p6�!��w��Z|+��"��w@[D�G��(��իR��SY/�`���7]
�ݵ�$x���Gא�+��Fs6�N�O�v��ATQASvH[�6�U�ǎ��+���{K[N���� ���c9k��>[0�}.w��j�r���b�T��6����{�1��k:F��%ό)�q����'r¸>sU4f������uyt*�/%��ZA{���K�X�4�����ޡ"�v'lȺ-溘�[���>x�jP��ҁhPH)��x_V͞9ʫ={�1YV�k����z:)CWϗ���$tV'��tb�?�9���OK��v�F��ÓP!_@���s7����И���{X�z�4�,�����w	�B�<�s��b�w'8��{�^�[j��o���!	�@�YC�O��T��)#���W0�X�T���m�CS�"�C�^ڹ�gY?(���d��7sy�mW�tÓ�>9�s~�����흗ڏ�Y���p��9�-T���]A�EӹZ�[��it˥�#+7�%5A<�a(+c��;#z�s�?4@ͧ�ltv�����8�]�	�&-�%Z�,_}]݊�p�O;��=��|�8��,���5p��2�\U���wV�[r����j��B�!	�[ZRW�t��R+�w�E�]��%�k��trNKWtd	}o���E_w(�϶c���Ւ��c�ʭO���R���f(��8吱��o����Y�z���E.qH����i�\�˾��y�)W0:9m8Kg=x1�=���8������8q�x�����͎��9��1_#&�
��W�rx�7P{�z�ۛ��z�0��j]��w���8%��Oݻ#P�����Q+��^I׷={��ʸNC���|�ou*�ܖ;��#��ȇ�-��"���;_2����E��tX�qϵdr�e�{��Xxotm�ϭ�*�^�7=���ⷛ���?%`	��\�F���ff�9P�t��T��1vNPs��#mt#�����Ϊ����3��@�)�1�+6��N���p��c�wF�0�QX�QT�,5
�/l��ط�e�%k��6�7�(�L�M|tm{:�䖫*��h�a�M������C��O�$�F��g+�%HRAx]+��P�A_	vYy]Ƭ�����C��q��4ޞc䢀�W���p�� wd��
�tsN'!ڛ�b7�e3���w�X�3N����Rk��|�����%���T�+W	�Z�Eg�PpqF6���P4*J�_pGٕ{[���F�A]Ş�q�c�fT.6�D��#t�I��Hp��6�o�-����!�bͥ=���y���La��ެ��\��������2&�$/����kJ�:R��%Rn�s��
M_1��G��c�`d"+�D�\1u�"m�G*�w_wN�f*5oT�Z�k�{&oGV<�n;bPy#ha�Qp�$���\:��+n,�aVT��6V�^'���[����s��y�K>k�(��PCd����R���0s��`�"$cVLى�*�g���������wz&6''Q0h��H+.@��X�(�Bf��ܪ��@U��Ǐbd-)�zEԋ�&�ʭ&L��b��q���q-.a	�E):�V���C���MF���!��otĲ`��:�o	�t�ˬ�ʗ�o-|�r�Y�1Lɿ����0��)i͑˔��g�#�>y���l��>u��u�rY5dCم�7�Z�uN�qk���e@A���U�ԑX��m�ݹ|�p�ld�^�(��3�7�vM����"�� ��p��+�vc�j]��J���2��vq-��%�*юv/	c��	��Uۅn���4P���أ�2��f1�ؗj棡�������R��G>����]�s~����	UH]Ǽ*�h�d�;6�U3&8�_"e�0�Fޢ�s<I+��ϻ�F.s7�{�,����z��=!%S�j9�7�e����z��*��%���h\Tힽ��6���{sk�Έ݅��+�s�etv�O����dME�6�nE�ZE��Hr
�rS7��a�z�`��Ķ��ȃ5�uyJ��Z����������8���+��d��A���&|M�M���X�}����oA���O`���i����{{�{.{�D���v*�ctk۬�v�n[DS{���]��k�"�d�tb�P��KX�[��3�v����'��IR�\���f�,pD�^��J��]Nh�:��W�*o�U����������$mvB���q��P��"���m��-*��|1�dGlu+;�DK�|c�-cA�*2�����v�U�s0�\��gtdW���A�!��y�Zk�֬��Z��b��n�Y(0]�)�U{#����F�-�X1j<�C�Y�p=gwk'>wv!s��8t���)Ӑ�b�Fk��Kj9<�Y���7Oq��<V!D����Ӭq�C)Z�ܮ�}�Wc�6�l���������#����5.�D����:h����q�[Xv>�j��,�V>Ȩ5��s����&���/��:�8ds�e��g��.�a �C��-�u�:a^�+��I����
�p��,����jޝ˃�"`.̟E�>Z<��3������\xtT]�x� Sэ��H��>�;/����%W���%]����9Ր��ç7�٪����F�N�8гe��e,���i�6�n2�#U2*�Xȕyd�� ES��{�6��턡\2^�oFwGldsumF�Q���t\����5�q��.`�$p�FRF!`Z���'��5�F>	��Bs#.���Ĳ��_7�Ў��Y$GVG@����#3q#ZGw@�!TM�;v�4�/WP:���=k&���l����{OR�EF���`u���G7�1 �SԗdP�̬�=B� �lOqBp^E^��w�S���$����>�qm(,��IyJ+e�͚+/"^�;�6µ{�.-^(��]&ٌ���Ғ���+����˨���7���wJѠ��5�Y[�.	���B\\B�⳻�K��
�����A���ZX�j��$����8�,pٮ{��Vw_:����x*�ŭւַv7{�|]g�R��]�/��Kcj��5�ޒ̨ܫ뫚H�'L��n��1y3����V]6e�ݛ������ow/@N�
��~J���nr�8��}�F����D�����Х2ti���ۨϼ��t��a>j�Ͱ{��s3"�2�V*.Դ���a5�n�̛�)��z�>�ެD��;���cUMU}B�e��cl�,�}�{�_7���ι��d��WLr����������uo,�����	vv۰s�[0~�R�#Մ<Z.p +��'v�Fw+e����o��-�ov���{	�Kuz�+v�(�����c��s϶��YdC-d3��'��
[�fT��ll17w���m8M�}�*����g٧В����f��UI�mD�6��@r�bj��F5��5'���`;�����D%��f���`�1�{@��Q����9�#yVS$C���w�X���:������i�ľ��:;#�tg˜\i��{]�,��!�ц(�p�<D;荶5���Ѫ�ܙ�o�Ǳ�ԕ�WN¼�8�Out�+�7K]��F���%�ݸH�6��v����gl_#���;՟apj���>�W<�|�9ի�r4���HR�P�2���R�7dM������OFV9(�"�W��=��G�[��������N��j��g ��겮��4�[�9/r噊lP�<i���&X��Nꀁ�2�E����Xi�L���uf��h��S�*%!Cs��-�*9�K�쬍�����.:M�-5�\�� 2 �&�2n��>�q����{;��������=HwU���t�Q��.ʡ��$p����k�\2�v�ݬ�U�2x4�4�u�oc�wϹV<��5n���6����xF�I;(@���<���w{�m��Vg��S�>o>�Բd��fN*ޢ;��I3%#������9��}�ϙgu>u�.��{����8�z��F����ow�!5 �R #����W�������.���x�9=k��lSL��[&;��t>�(T$-�w����o������l�PH⍥��u3�9�K%C���;���9����cj �0|^��[-� �������7�{º��t��!��v�4"G�	��'\],W=������j�h�Me�ܸ��V�墲�q�7S��ݞ�bkJ�z>K�S<�!9� oj;��}��O���������-E���	E�NB��ֵ�,Un��F+�P�M�s)�(U��|��9��&{^����_{غwP�۝ށ������ ǻ�
�a@�]��1	�a�g���Ӿ�"-�R�癇}������{�����c��2�{C@]em��fKݔ��A����ݓ���1d�a���y�V������2�����Q�C(t�S��~wԠ�� �n�*��8}�ih�K��m[��w=<=����#�k-�����(�μJ錃���|�cn�I�,��,�6=��M\<�|y�E�g��<�)����7��W�
`�g}�q,� �FsR��}����<�zRT�G��^�����wjkhv��Ӏ���3 񰫄��,{�i�p{7���$�>��a�oV�{�}/^��7'a�}>k})$�|�;�x��{ڳ��j��ϣ� ��g��R�1����<���y�u]��
k�Vi�8�]���%�/4{����v'vۚMh�;���w=��zK1�Vy��f=f�j�x��Z}�+Nڡ��]Ş�}ϵ-:Om}=��	��N���/��)�0�
�/Z��P�F�`F�����xs�#��S���	d�uև�)��횏t�����ByI���u��|ޑ�$=n~4sg[q�/vŇv�����{��7�j����3a�M�2i��t2���1�ax�{+������z��zkcV�Vn�F�b�H{�=˚����м<n�yO-��lXWR�Ţf�����yM��^�Є/r�ÉX����R�׻nq� '��d's�>�Ƚ�*ٞ��������u ���Z=�m4��ׄkԭÕ/���e.�6v!Kq��9
��hy$�Eع��g�]Xow�Э�;wd���C��\���1z=�����[���-_{y���g��";[��~�����jiB���2xS���e�%D�>��i� ���Y���JqW`Y��]�W�q囬հɼu+0�I�^�h���&v��}���'_j�Nspa[�y�N�ud�ȶ17�sVm�'X1-Z��B���M<�q4�阒�ɰnKc(Mr�p ���ޯ��&M��Vo3��lT�C�_lZϭ}=��O�|���M\���Q̶��2��7�b�X�鸽'���B��A�a�lo�*zĺ�����3y:��ؽ��:��r��;��us�����u�ؼ����)3z��u��Z8��]��s��qI���S���2��&ҙ�.���.t�bt��J8g&�h��� U6+&��n�)�.���Ƀ��]�;�пw��)�U��"��j�v�@�J��񿩽��N���VAO[������d�V�f��*,\	�,�pvk0d��I��`�պ�-jM��|��سЀ 9��@ ����>�uk�N�g������_���}���kSfk̶�I�G����+j�yy�=�ڳ��'���m�$;:�;�y������c�����{�fo=�{[���:=�����xmo=�Y���{j}��m+kC�<���՟R>�3�N�m�{؛���4n��dRyfe����o���ͭ������I����e��+���Q��'���$f6,��3�k{^���/kǱY��g�Q<�畞�b����ͳ�u����}��6�E�1��m�9m��m{Z$��Iyby[��X����y��������{j{[��[v�_o{N��i��������"�;�_m�g��;�ޙ��h�܋Ò��}�#̧[9m��kE/���ۄ�;"��;�<"6��f���tNS�B�w�B���	ZҴs�K��;m�搎���."�����	_3�y&�^�ݼ�NN���dm�#&�0�'�y�vq��b�>i2�3Ěp�iY�%m��=f3�G�0;���}}�˓�{�Ȁf�����Ø�
9C���v��unנ97�R�6�Hb�i\�|ч��fv隹��{�f�C��Zˬ�zS���L��@�9�by�{aP��}.w�m{ff���;��Α �ͬf3�dT�^�x��2�Y��}��V����8�鯅׫�2љZ7�ڬ���F��m1��^��[��;�t�����;]�L�^FǍឱ�,��#"p����p�;ة�����~���xʁz���(�=p9ЏC���K��,.�x��(��#�<&�?\U �6;�A|��^~[���,<�ŻkvCs,i��6p&����ո�wG��n0�����F#�v�f����\��Ly2���{�p��s�o�i�ς��^k�p�T�㾝�tX>��~q_e΃��� x�v�≇�9�Qu��ɀ�K�޷m�6�~hZ���������Ԭ�*��(���}]����S���T<;^�G�S)q�R6�4����.�Ю���$a^=�[;^���1x��z�	�Pq�RP�+jj��\vv���
Z2�U�����^�w�U�%������=l���R�툷��b�Ǖ��G��&�n:4�;B�VK�5�L���O��p[�6p����ʝ<_쵇J�͙����ٽgR[�F�����?5��}�9�8�f�����;�w)R�S���G�|t�Eu��rE��̈́|NGXSd����
��{��g���|^t.EZ�R�ק�	>�({ej��K+:8=��̨����`G�`H@��D��TI��94u�`��^j�阹~>{�]8b�=8���)M�Z=��]bLu�~�z�owy�>�y�oq��}eNCG��<�����9�U�x�sjp��Q�H��.^���Wח�hw\v�(��1�zW�]���G[�n+�����D8�ԩ"��7OgD�Mު���{v���;�$�@��)�^_z���+��|H�L��<�T�<��&�x���+��r�v%w]O�Q��czo�^����N��bvO�骹����>�R�rbjh�zg��G'��R>��ΈQm���mW�ߤlz�H�,��d���P��}�;� 75)E��=��S�����9���(3��e�m�D�M�l)�E��$�" ���1�1��O/!-{;���b.o�_z�X�J�c�X�㜦�x��ҁQ�<���w^��/�el/9꩙"�V�J$���P'��w<����u�]|8\:Mr����D���Xf����%3�a"2���sCr�cے�&FcQ;N,�\���H`��O�`1[�u���P���72����
Uz1L�Z�V�	N*5@��UGFf�>��֏7�
Jt����TF	-���p����3.0���7c
v�V�K�R��x�~Mb-�ǣz��k�?a��Z�]�E}�:!�z�!�U1_o[���	��k<��F��,I�!?Fe{��vǄOW�����CG�Ha��A��tG�Eϗm̏G\!�z�u^���5�F�z_i���/�##���Cl-��P,I�<h�����#�����V��k7=��&����_Z�'n��񘰽�ټ	҅5�>"�f����'Mv:���Y�z�c&��n���aEx��Eb�Xş)��g'J�?ut;w[�`;8��D�8rMׂŦcUon���;������G_]��ڬcf_���S�7)�e"8�WE�C��ި�)H�6�%�e��b�z6�b�QH�z3�'Q����_�m@赭�Y���|�D^�������T��B�{xz�.CGAP�x"�����������}I��G����8m�%�{6�н�<�~�̹��'�F�G�M!�"�D�Sl����DnD=����y�q)�g�Cb���!�CD���yU�7�h���z��Α�Y���P���2���0�;�h�0k�9vl#=ԛO�I���$��l�,��;��N��MC:�Z8R���L�	&K��{h�5f��b���1��^����f=���6��7�nC�O�p����+�"�18��c۹V��,{�#��|���2�]�ws��=+��-�0ץ�m�Pc���Ϭ���.�n&v2lV�++���t���[ft?@lDPU�^#�3+�
ۨ��r�-�!�ް-`n�loW��	O����}�ćn��0�K�E
����{�[୺�����q��A�~t)�5)~�s����s��T�iV��U����A�a�E|���Hl_z�B(w�tqb\|�yש��B��q����_����{��j�-��}^���2����ȠC�%�}qRf�z$ ������sv�o�V��W��oj����6[�7
�j�;9�Y̩f��v(#Eߦ<�x�U��]�֓��Ӌ��y�
v;�����l��h�q��=W1�XS�U�#L�A��z��ȷ�ٸ|���(�����u�P�o�ZŶ䋼N�M���ςr�[�rz/�EmwV��\+I��<�5�ޘ���1^�9,N±�V�U9F�[c3�	ړa�{���w��}X3Ta&�}��.�I��Y0��������)D���=�d��Nї=<��6�þ���}��g7%f<��=�ՙ(bA�?u�R�	{�M�W�n��oː�/���W#w�̂��f�A�&0���)�S�M)S��:e��;��
'3[s�)f��+�
�o���[�6���-� ��C�<����^�ښ�}T���������H	�[�Gz|F��k�-���ט�t����T A��H,G����b7�ȼ�1��R�����E��-n���LB�gW�w���X}��N0�)��H24KG�kN�]�깷�#����^^ޚ���&9�ץ#�!Oԁ����c�����Q`v	0��&CD��+�\v�R존n��v���?U�|�}�4�B[��M�-�a�!�+�Q���6f������Z�~&U�����pXb\TRv*�r9�9���q�E�ݮ�&��8����H!f�^�W71���xʰ���n��{�X*�>�Pd`���)qB���)�̿��7	��2�r�D�
,)wPqת�x s�]��]��7��W���2�u'�E���}>����S���
ٿ����E��j[���zw3������s�]p�1��r��@����xe|L�Ñ�P��{�X	���ሁ6V�[lP�:=�n,t��������y�5n3>��GE�g�p����m50�z;��ڴ
Ǒ/���b��~Y���o���r�2��M�qw�|���.�1;�T��g{�w\ͧw�J��{�5dg�t�幼�aA�W���5�;qu.1N�^�{��꘍C�U���}�������w�\"�	[78�qb\��57�f�|�)�
�\�~�X�i���'`s^�P�R���.��
f�y�:/}��H��9�6.��t�_�g�zHf���{v��	1KU���!E-������t�e?q�j��P:6����cxi$��U�*]}G�ُ|��\W	q�6�u����h�Z�cq�w��y�/��]��.-�֙~�hs����yp&�]@���@s�a#d�>;Y5�u�~�n�;���~O�Ey{^ї�C�Q���&��6LH;B� �����ƺ��{*UI��k��ůb�ѱ�ӿF`�I��R�x�_��*#o�&#����K��Ik@׮�Z�dS�kK�0ʰ��ǎi��;N%����)�3������G���,34��O=�Vk���~�������q��g�j�z��l��CUp|�sj/�xaq{G-�T�y���ρ!ј24O����zW��t7�wX�4�[���c0��8�q�I?b���So{�O�ܮH�z^��=chQ2�4d�PWM���vﻝ���Q�.���w�A��=���}�
M�<��F�F��6Y{�v��>�,�x�j�����r9�ץ%����th�rc�ֿ���D��\#d���	S5��:�c����ɺJg���u�;��+c�^�5����g"���sB�;s�:4J�b�5�.�#�>����o��j���\N������o�a�{Bɟ U1?z�������W��=������~S���a��/�ňp�J�j����v�dhq�g������~��i&����ﲁ=w��!��y��&.׆���ߢ���Ų�6�"�7��:��}�rU���q�I�!��)��f���'D1L14���s|b����Q	��L��)�[�B��S���������p��sT]y�v��]��|���(Kg�]De��l����;��~��M2��݌xlx��P�u�����Qވ��1�3bo����h!B�_�[Pڔ!�I�#@�*���n�4�' yĬ����|_mO���]��h��%a`��#�3�zCA���u�AdW�{�D����9���ީ��|(���jn/����l-��W3�x��E�|hIB;�}���r��纅ƿp��ӱ��@��O����fӞ�]�!���N� �vVx�gd���:3�g5���s���\�+�W���4���N������|��|�`;Y��VFy��}}���R�9�o�f��U8��}��[�f���4)�W2�:��p�9��㓺u*���a����jgf�hY����Go#���=��o�bn�gu�8]Yp�lh�(dL����a�A�s��vS�M�`�oC'�����g��Q��v���?�c!�����!ʇ}t:6�U�x枑�!u>8��F}NR#X�qL�'12_�:�&tG���U+�����f�=G�[S���a-n���Y���]��R��5�л�)o�:��ɟ7p:��pAT�Q3�H3��p'&����[F����e�3���<����t�Uv(��q��!x��+�rpQؒK
E-�j�m�@�f�{��I���U���n������8����r��,O��
��Q2u����ٔ�Y�"Ƣ'�{�G�q��wl*"�F��Ņ�b�o��j��;e�I��8�f��l�|}����B�M{�{"G���{׌��贅m�d^���[>�����Q�o:�!:�!����� ���%�����]M�w�pg���z<$�|6�Z3��xbܗ:�ў�!�G�Ǎx�V��f��5�f��{�`��%ZkE\�1�9�|$�����P�:�����wΌ�F	*��~���G��^*��ŉm�̟W�oN��7��Ѐ�Il	!~��VOK�@��vnr2�lV���`R�Zy޵�k׮ꂯ�&vYy���\��|ǜ!�Oks�n-������,S��p2�k��z�VO}�ȝ"T*�E��^�v�s2�+%x����8w��A�r���A��c��c`�9 �"Ƥ�'�9�8]��ᮩ2���6_��°ڷ��q�̩�j�M���L��ן��g72�m&�~��ŵ�z�obD�^�&�t�.5t�~��+�깎���Fđ]���Mkٜ�W�}���=��\6.bW�ĸV:�8W��X��m�"��N�J�z=/��ҔT��1��c�� ��M����A�?)�������^|�����Z��g'jM�Oqw�٠��H�̧��P���7��H�68�Gl�$1=T��zD�=�5���j2 �����Ƽ����O���p�gf��9�g,��(����
rJD� �O#BLiqC�1�-�� �S�!�@���{jVE���:v�z�����i�(��eD;S�*R" Ήh�N��b�~��=u�r�q�W������*�hDmw�����	��)��h�����4O�������^qᓡz�:iW���>�T! 7o��)l�5�0�:0���#��׻1�j���w�U����L0�����l�\�^]n>��w6�No(1�9N3�V!,��u��K�U\����WP�Qz�����7�Rq�� s6%�JilиytƩ1ZM�^cD���5_��0�Z.j�K��y��j*�k0ڷ��F+�B�j`E+4y��xg���E�<ȜZܕD��K�sd��um�S�����%1�� �E.���&������l*�f+MA�⡆\z���)�̿��7��l�]�NvFE.�І�8�/W�����K��my�7�]�&G�N���~�����{}���r1v?%�U���݈O�u���pSU��]>�7�Q��,23�&�?^����1u������>�qC��G��z,t��Fa�����q�3�>��Y���d�XG<��R}�ݓzQ�L�1b*\�D�7�K��:f�l�L�/�=�{ݾ�"��;�RG��t4������>a���b2S�S�[F��NH����f�Sؑ\�k�uX��TO���Df�,7j���	j��DQ��dLN@��B~��ڞ�mz-Z�cq�_�=k �V�}�kn��׎c������a�\	����>��g��F�NO��6]K�9f�����J>��e�h͕�n�du9Oq���9��N��,t�_@=ƾ����ULA�S�>�]��
�}t.��_�0oSeF �R�y��S̨��ӄ�w�t�C���ɞ����˱��hO��gű턄U�/�S=��y��}&{K��������; l Ya䷙��A&�kN��eT�Z����AN��-�bdDͼ�`(����uԛ#;���kܨ_�y�nt�������FK��9A�����2/u[����o%�E�����V)���3�=U���5w�x���e�q[�w��������Ulo f�ѐ��������MDR�u1��wT���j�K��3��_8�f�l�F^�2��u&�{*AUr�RChR�+rw��^�w�/��Ӧ�EG�L��,L�u���}|�[�x�'�e�'HWj��C��J�����B��iS�M�|������5[1�74��x��Ë�L�g���"o�-N%w�نP�0*c�bb��҈��z�fkcxL���K�ˡ_8�Dje{�H1WV�()�y��4������us�=B�U֗^��0�#�~��$����{#����N�ܨ�h��V�.��G̒����xrĪ�)��,��j��-^�M��75������9Ƚo@f��f�RZ�K�����M�g�;�20^��|�zl��������H��3�S��x��>Lc��{�篓Ú�ҁA五���&�j��n��E [�]ŵM���V��x��w��jO�xx�D��0	����'W�r�轒{��Wl� �M)�5t�g�!�\E�{�&�����,UF�Ӳ[v�;Bg���w��߽�^�(��|U�,sC���}�\������v�ձku������n)��	�;����;T0<U�tn�\Z��&�!�>]��*g���{}l7j �ʇ�]����>ϝΠ�ԽS�,b��B�oA���{����OޒU`xV\s�"|�5{4��ֹu6H��b�����\r���ޯT�m�y��x&�����Q�w��Wo�gg]�y/u�f�
zzI�e.�˧��Q�L>�����=����=��{���)�=��u2��#�:���2���a����>��#/\<�T���ϵo"��7�\�,2�6d�ٳNٮl粵�-��������1��4}g��N���@n�<:}z[;�w��F��c��ps��!b�wp�q�p�4�}��N4�h �'
sS�˙ݍ�z����p�7�;�9�}��$��ws7�a���5�d:�3G-"��;�#���P�6M�8[�Ɲ��Bw��b�:v�ﵕ)�چ�B�r���gC�embg+>��%�a���|��d����г���lΉ[�V��:�5Jn�Bs�n�ǒu=����o=;G�/Vȭ��v���>�N(F^��E�EQ�r7�[�K�TV	��0�U�t1^�E�SJ����/5��I54�Ԍ��)�p���l�_.�:����b��[5��!<����K2ɛ��Eg�'�\�0�9�]S
��z�X��ǿ?������\�i3~�]����,+;��#�ڈ8)^ּ�{[�=�׶��QQ��ܓ��g��P��[,�̢D�b���v�C��s��8�������;���.:&Y�iĂq99'H�,�;�c�f�A�pu��OMgk�����ȶ���%�v�r9<�:N<��9#��^[v�7�yZGyd�3�qӗJ$'�J��B�Ĝ{۷������#�؄�&�<��9!I�OlQ�K�� �$"�[�$��8�����,��kmby��8D�39ųn[om���u�(9ɵ�z`䓧H�Μ�=�I����։��ydq������#�Q��� w��9K﷜�H'83t�k/�nO}��w|����ݻ�"�::"R��pf��2{}���<Q~�ަ���x��v����tX��,�!Ǧ��./%��+9i�{��,Tb;�ك�P�*L:���Q�j�D}p��S����&,�o�a��c4�u�
v�K�����E��`?uc�y���_��ˍ��.��Q�� ��.W�\j9�\�=-V-��Hj�����Vt��>�s=��ӄ߄*���$0<f�.O��=WOJ����u��-����c�<D�=	{]v�gtw����Ip�g�l���L�D���'����l�}�^�¼;��ٕ��;j�rg�Y��~:>��H���Yu/�OD�j�W�}͏��W�,�
ES�2�	�P�5Ҳ��"��Z|�����^	��=�0B��(a�Sa�^��/�#�Y�l���=y��i�Ӫ��S^����#ݵ�Ƅ�;�c��f�N�� -����T&��B���z��J*6�p�f��/�ml�7�lt��\\n7�,w�aŉ��<K��ܦ�x�b��ޘ�,B�q%ڿ	y,-��;��K�d����FUD`�ُo��
�q�c�\6p��[�<=��WVM��N�}��c1�v�����q+�uz>��!>���"�ڔ!���0�P�*���WD�k1]��*}��uW�h;7�J��1#;�Zl\ޫ�	�E�B��7�f~g�T�2'�c�������t؁u�����^ێ�*�i�Æ�� �n/m�BH0���cԿ]���|�X�`��^G��'��K����2��_������J��A���=W>���F��*��	����cO��������\���O��:�t�~���W��5�*�h�dtS�hm��|j���<`G��`����
�)��v�z�Ŵ"��4�n�b�-���T��Z�Sf���B����Xf����:gc}隢%�v��oz=�ꈀ�' �:�s|^+��Y�ZFg'j��������)�1��]s����B/7Л������0Hr�_�t:6�j���zG`���G#;���V�{//���f{��=���w`��p�)8�%����V6�!��ځ�-n��Ei�z��{�����4�"�:�P�e#�
�B��� ��%��2k�qeO�^�߽�<�w6S�����~��q	��P2�jU���U1KD�+�ȋ�G>�D�E }Ǻ�z�~3�U�汚�~�|r�ʄ�?{ӈ��	a�E��1K�r���0��uz=�z.���V=�H�c͉�W^��>��sNF}�/M��l��zXf�~��5_F���Y	�����3*,x����4�MR9���'�I���&m��-tD�v%��i��:��d��w�D���������s����xz���/5@�����ۍ��wu%u[�]�5I��h�S�6��㋸�Do9}��� �kۥ�R����0�aB�~��>u{�ϫ�������	�0���^��/@̮�Y𭺌�΃Ӌe�o�B��§�dԾ��ܿ=�7���/���
*nN�8��^*(z�W�;Ϫcat�N<>��*�*(�T�[~��Ʈ,�F4v �d���=�rta�����@�I7+���a�5jFw��;�ۺ�y��h�<{zT[v3'���N���9�ȠC�-��u_m��SQ�uO5���/�`�ǜH�^w�}�T�~Fj/�q��m�p,��w�Q&VI�2P��}Gj3�x��$s��&r�}r�+b�5�rw:m�W�4_��7
��s�QQ�~��X������u��B,��<�z(	bTu��P�-��Xے.�;�7�^�g�2�n��ނ�tw�x��i/,7l�]	�uFu�w>�?9�TlP�����Z/���ն3'jO��:G1V������w���c��	�^��l#��D�=?X �=`m�Ƽ��E�ܩ�Ҿ�풶^���]���1��y��.-���A��1��) �@�ä��hI�.>ܽ�����6���ϯc풽{t��n�[�w�ϥP�6[�g��D��q�4d�!�00�Lf�p3h\j���$bfͤ��Mi���Z[&v���Uz�܉S�=�O�k�v��=�RK�=��e�5e��PT`�P�D#���5�͘PR���yW$l6��"$����|�e������ty��~�g���}n���W���g�WeD+S�*R" �P'(�9Y�>��vQySxZ>W0���C�M�!Oԁ����`r�����Q}�L)��+�:��~|9�v�X`����#�N�������V!V���%-��!�i\�:g�c��*�-�ij�=�����xf�=x���S��Ϻ�4��]n:;��D���ݰsA�O��|�].���cT�Ay��o�a������99�(��j�k�~�Z�`�]�;��r���#]n钘�a#��j%1��E����{k��*̾�D��q�E{�"�\y�ڼ}�0������?�͈\ЧJX���,SU�����EY�|0���#Þ^��Q���ݯop5i���lw��ʺ7�Xd_)�l�ɺ�yM[��3�>��Y�q�6u{/��n�%��u��1\��A
�\o�i��&Yk��ȫ����4�@���Z}�Z	���՞���גW��b2(Ju�6�;�m��9"���l�4�d]�gD�U�==���̞�$��v�Fn�8�M���r�Ea��\v�@��oc�ugb�潫�pŃ��5�+�`����Y����v���e��x�D��fC����f��!�M��v������������"��%���ҽ�\ɕx�[p�~�DD����n�Oј��O�;�6�㾁>����%�mJ��ȧ]��s]>{=�i��<�8j�@��&/=�}%��q��46��o��M�W����E	(q�a�y"zpqΌ��ω�Ǔ}�����k7}�y�Fl?P�tl'=�����F��;��HU ����>�7^(�tvU�=����U
��]�j��3�6T`z�a�y_Hwu�8LF���tsj-:_��ڹj��o��0oI�eq�1���B��9������ͪ��)��X��U�h���Wd�>#��b=R2�'���P� �Nƣ�a��m�BM@|ǚ��2�^��Ƹ_Onu5�*-�����c�=WOJ����#��V┄7�7�tVnz��+ő۾uf�Q
))RE-���Xe^Тd0Dč=ut�}S��V-��2���a�O�g����%눛�$b�u�b/�j�dz-�q�2�hY2<�`�X�#�p��}�9i���fV>����W׸�׉����qm���o��b|����c������O�f���ج�g2i��ZWLf0��?d	m�q�!�����2���;������������!ܗo���&|m���^��GJ�_
{)ەP] 6P9Pҹ�)��*��nK���s��d�[@��2��h�ԃUB��6�a�ޓs��*��v��}�}g{G �mY����Dz,q��wN@�������`�a��e�m�EB�����Gen�1J�����W+�rۏd��#+�H�܋�F,w�a�ϥ�:e�~89M���n�5�O�Z1����vi�َ�w3�lYw��2(K��ʨ�[1��c��8违ߧޢ<o�����z�����a�<��;�
v��v��ӑ.��P@�2K`���?w����v� G�����g��PQ0�[���d8O8дm�V	��6O��
�h�1>�3�+_i�vr(�נ�'�cN�Fï|}q��{ns:�X�d4_�2:(=����ھ5`L�4>��c��TVg�C���XairpC��i�+��Y�[n��O�ůe6o-;P�?m�
fI�.�#�ǟ:w���
��int���(��#���L����7��XŁM-#3�������lA���/�RXLM7c�Ed�a~�!��v ����¿��tolB�4�G`��O���a����P�ۗoV��iC��Z"�X+�E�W�R p?DO�l�T��U��C��P:>�,��Ś�;۽;Pf^M�m .�U���2³1��L9���
�m^n��g"D�ͻu焢ͩ��ϱ�sG�3CZ��=2gTe�����}po�^?"�<��}8�{�>���w��f�����^���]�f�������Vb� �ܝ�!~����Q��u�/s�w�u{ �7Q���H�6�*�
'��+aE�`U�4��xUN���)�h���o�D:}jFQ�J���U1KD�+# ��$�
EUt]5�����o���5�^���1K�ofb��z��~nC�I�/	�v:k���r}�p9~�ؗ^��~�����"aȪ%�������ӑ����ݖ��������ߨ1c��������3F�����v�FI�+�A�T���޼E�etb�����!����;��2��}��ޞ>�c1��ޯ@��7%�,z��W�J��H�1`k���V�GA�y�E�Λ0=�M��=9���sht;�ų��lf.��~7�b���#���@��6%�:�l��[S6�vk=݇3��G%*J�`�4���ŉm�������n0��>�]�{�tV�>Kul{q��T��^�(w��[�M����6_A�M�(��,ʖay�����g=�xg�p+�,]De��q��(B��(S��ɯ���p�h�8�·��\�X���Qq����9s��R>о�� ��Y+g{WmZ�+�<	�����j��[���w}�sC�s�[�LY�!��.kNw+�5�".x�ˣ��fh�V�L�]7.Z�3C[�Ԧ�A@ҬX�2Z�S�v�U�6+Ef����b��=xY�-: ��������  W�37�������H� �q:�z(	�*:�]	nP��NH��'}&�63���mq���Ք�4ۜi��'�Δ�Ȣ���	������u}^۱�c�}��`.�"g�S�Z��[��Ey�ۮ䱮yx����� ��C�,����A{��uq���|���7/D+׋z�&��69�N���|q�H�x�E����S�
��@�8t�,O#Ll#�n�s58w�7��W{���)�5&!ic���S�9�:��8tr��]s�N0�)�.\�5c��v����1�~5�T�:Ͼ�e^���;���?R B��7�-p�)AgН�����uo�v�x#	��&G�'���"��[�#��>�߾��B���&Җ��Ć+3�:��}p|��]��۽Ncc����雓�����\L1⢤�6P�Ӌ�.��v���C�\V\]��}�s����&�~;_UE(��3|k�5pOEE�����߮���xR�;��VV�D��v�'�#�d����<s�kk��k��*̿�dρ�7���W��)�\�י��Ȝ��(2����S
N_WE}&Iݗ�a�TF���ǲ;�9��i����������3����6>9Js�7|C=�a�''�;�m�&;�yw%�\4�'������TZ2�Sm�6<px_q�!�Yp��/����Ӏ#?����mw=�2/�ԇ�v�7��o1.3R�!��ul���z����a�2���>�;�﫨���"Jjkw�|����?�����.��m.|��L�ȱ�P���ɺ�yM[�'p�T�j�=�J�_���Ww;��E��9q��1�T���EH��R�c�i�ς��^�>Y�e���J�q��[�=?z/�9�6,����!LFAnb7�n�C��`:^�$P޷m���vG:i��Wl׻�x�0�Oi@����l�~;_�$0��?'Җ[�l؜���u�N�������_w5S����%q�u6h$l>f�X��M�P�>��g� ��@,˪��K^�m��}�s��Fl�O���=�{���F�N{��ω���M�Ӱ`O�t�#��O+�%]��S���=V�Ę�ݫ�l�WB�Z�~���M��K��g�ܹ�>V*�W���8/N�� ��)�vx2!����l�cJg���*�sNX�;N����k�Ş~�9������5��ck�
A�%I��v�*����u�Cq�W�;�����3�[^<u���������76���������E�
����c}'����}��W�Y�u|��>�|�XN�Q�M���)����B�.���A�leh+�(�6Y�֘�ىy���7/��GI�N�Ck#�~Z��
PjC���D}��}��$��c�[��o57���ʍ��0gpEt�TWޫ��xu��ou������&�Sf������^�a:�b�n�4T��qk��hQ3�LO�2z.j[,��"ra�cK<�ލ /	ޡ����3z7�#�C����g�k�B�#�H��w�3㵫s�ޕ�@��q�X������F�K`���8��LE���o�^��.;�_���;���Xa���)ڝӐV�mV��_���;��a�~�P��^�,�u�5D�Nƨ3USۭn��:G!��IXDBE�	�\nEͣޭ�'���L�Ǒ�Z�����n�g���iQq�S^�}�鍞B�{�rJ��>%G̩��Rً�}F8W{=.Q�!��vH�}�j��X��^�5��m�ǟS��̝�@��ӑ.��P@�0IlCjP�+�i�=�xz.�Dׯ?�/ٽ>k���ߝLV�V��#!�x8дl7�����1�00h�1>�.���.��i�Z�p㫍E�c�b��#]�p������5��鞃�G��bƌU�����dȿw�~�F�'���TF_5���o����6��M�1.Μ�p�����Zuz�mcZn��{�$�hŦ�{<..�ڑ���^ j8�\������Ε.����o��9��Mf��� �=q}M�Ԇmö��>��"����\Og9��o��Fi�V��'%7d��9J$���t!�Y�c�<��>�YӅa�A�����\Q*��Kt7'������Y��bM�wm{;ݚ�k>�ԙ���P�E-N5<
Y�W���űi���y����Js��=���lU��-��4��(jg��I��KߎfI���w� m8x����{��r�v��<n-���N�gh�,:�a£�s(���\�}�֥�7�"I�5�����S�����Xa^\�Ċ�����ګa�Y{��@scr1JU�qLj6�VP�n·2q��s��UbtFF+�a�m=��R��ɼ�w����J�� ��Q{,	��bj��ieʚ�=�b���y�eE������(�.�ہ�g3Z��z��G}�8O\7��d���K���{�� 9�;�d'͂�;�;<<��)�{2�׉S��{�:玓�B%_u����	L�B��i�U�7�^�~ߞޅ�����yA�N�;hC��{�~��:&8�� �Bu���|<��P36Yȝ�E�^���T0e�e^�s�ލOɤ�3��4����3���=�ޞ?����'�+�Nx�^je��#h���Z�QXr�c*�c|��%�O`h�������c�J׺xU��
���^@n��ڰ���+��*qV�����*)e���$`*bV:�j!�I޷�=���š�u���N,Z!�e�{<b�J��n�Β�����	z�����87������3��ʟ�7�o;C+�j�������MZ�fhFNE��e+R�ŉ��b�7�����1/�O��� ��#�դ$��"l:t�t.NV��(l -<�MJ)Y�X�ys��	D�j�2����M�=��MU��� �`���O;{�UH5T�����,�x2.���ރs�ic����Y���x��^	�>�3��[��<�z����5=������O�W_�b/�Um�w�������<8��J��߷<���ߘp���Yή��|�of��Ó7�oJr���y!Z��t���*JZ�ժӻ͝�i�h�ȩ`��l���r��C�ș�1]ʲ���PɄd��:'���%n��������,���&�Jy��/%�ت�H�{����_��4{��ƚ�2�����v�f���y�K�'�7}7��CD=xh2I4ۃ�j��8J�9i1-�Jc1�u9�E����}�\Jޣ.�=���<!Ia��Ow12���W��!�s��������Z<��7�hLYCC���^��.��іu�X��W��x�� ���1�(|�9����9�<�܈9�{۶��$��C�q)%	{n��NgZ�{h�%$����ܼԜ�Ҋ	k�$����ґ�g6���'��DDp ����$�Q����s���9ٝm�w��mʹ���@L���bH���Z@�V��8�r:'J��y��j[h���!��,���|��;��S��2�r�R�[n"r{VFբ�$��m�on�k�n%'�+-!C��G��o{q�q$���ݙi��疠�ݸ��C�&�$��{XҴe��)������#̒m�[kY���À���Om��p)	A/k,�:���j�Y���\G\Y�b{d�bIC��pI�c����S�7����9�j<�ټ{Xw�eܑ..[מ�ǭ+��G��#*L�dV���;�x�c�r�x.r���^O#j?��������g�o���jK��\�)VP��m���O�Ņ���v-Bƺ����8���KNV5���I�urt�������B�F����YBҎ��PϽ�1��ϴ쳻2���$��0T7)�yLz1gb
��Q1>�R�@;2�� ˡѽ���sOH��wrMzg0��pe�^���P��H����a�R �Acg����U���{G����]���>Ķ��/�9���m� ��ג_�u{m�B��y�GAP�&h!R� �lEi1�.q���z�vcn�/�b;���	M#	LB��US��9
��MuǑmv�'=��5I���<؜�ri@��������N f��$�܆"��1K�D�`�=wy~��rm߂��-��\�����"�!8ȹ���To��|_�ݖ����a����;�q@��]���7�l�v/�������$����`������ws�iV�FE��A��[t9_W���U�i��y�Dy��z#:U- ��z��*����%Ǣ�*TP�H�1c]l6B��@���u�=BP��Vۨ
L���ɥ
v���{Wp��,@��f�s���Ĥ���\W���C���:�;V�����B]�|}�}ǭ.�>�*-��B��"����	p���r���[E@�{�g�M0Lض��b�l-ks1|]���:�}��8m��嵫��,VǱ��L�>��un�7�b����S"�>��<v����^��������w�_�]:X�)�Zr�8_Kn����>Ӿ2���6��XL<���ٛ��tNhaqrq��"�1�����yW�ުl�#5���n�ոJè�uҭ�l�=��]g���u���~��#�2�>7�\�
��
v�nM}�6ˀ�KE����P�f�b��J���=^][=�s�S�z,#L��7�
b='���t+[���䋼N�L�ɨ����z7V�cCO
ѭ���+�o����Eel��~��ŉ�;{uh�S�&�e�.�:d���=��޶-��ԛ��{��ݎ��E�ߑ��� �bz�?I��^�kce��J���^��梓�;�.��r��.Ԩ����nJD�älW7�ӉWG�����}E�&,�����w�����n}z��J���Uк�!#b-W�+�{k�����C��D0�H3�	h�ީ�uu�"���_w���OԁH�~�7�>��[�&�2�dL[ډ*w�w�6�q�0`a͹S<D��	[���,��5�$Ŋ�9N���(�l������5Xށm�
��s�n5 a3�&�*�0roc[����T�R�
pm�6�@7
Z�S�5d���0�]eJ�7Oifַ5b}}��}I�u�7�n�
?`�C����t"+�n�����[�V!V����l{v-�\Ey�>J�ח��ņ�s�F���.�5~BTT1��]NCg �Ӌ�.��{��IN�EX]W�M{��%)�m��Α �mc7ư�lL%�N}���sp��KWn����a"��w�����VE�N�7�b���ŀ���~��7�xe�'�C}�\��q;4%��^S���ae*��Ⴖ�Xl��7��JX�cul�5^�.�x��(�i�����]vΘ�M.Gsw��R:����T��A�|����)�l�M�Ö�ŗ��P�,Eg����}��CÐx�a9CeF�(�{�R�>�HC@�R�c�i�ς��^	���_5#�W����Oѳ���oH��tXӒU�:x@��)��T�����\!����9"o�]M.|Di������c3H�}��sh��еom@�O�����@����(K��������Rʻy׽�o��+�M��2��S��q!"�|�����]@��@U�F�!���_���VQ>���'3:��3>¬��(��}�燡�H�R��7�d|e�t*Nk��T�Szzr��6�T�����i	�{���Ktd�؋lq�靳��z}݋]�����'����3��7�#�K�G�BFd�%���"菢>��l�[d�)��Q�ᗓ�B��c�\�{=�~7
}���ٶ|NG#D��K��D)����������swN�k�0�����x��¿�+�foSeF=T��<��;������T�_�y���s�b-�s��$0[4$��Z6\��ڬcϜӁ�h���v|�}*|���f�� X�����_<���SF)M_����AtUt�e�Rߞ�D)��e%;��f1�/n����1A���ڋ����8	��%A�*��0�!Ͻ�LlQ�<*����)ڌ�r�cj�+ n����!�EID�68�W�(�1?h���p+L�t�A��(L��b���\����d��ԑ�	ס��9�1C�3c�a�chY>K�S�n�W{y橃�la��NVG#뼯�i��R�"���/�x�v#��3[a�5×/{l4	���c �l�28t�W���;��:�Pm
ټ���;�XfߤT+��)�L�T@:|��S���٣:v���q0B
F`2��ع�b��VË�K�c�X���ӂ����7��ї����b�3X����U`�sW���t�ar�.X�7�#�A�=��ON�PWZ��vn�Rc,j'+ki��ժ7v�SU�����z+������ݞf���9ޛ���23[�ɍÐ��޽|��n�z	�'7��  
����w�e_>��mط�����迺�$��'�g���T�f}-�����x��5���:������w�FB%G��2�&�c�)�dfNנW��ȗuz>�O������o���,�Vg��+^玌!�u1_o[���p�4-�OW��O��#�V���l&�E{��J����';}tF�Ȩv��c:���d4_��s�]Yyf���(�H�ҽů0��]AE�A؞=4�#��\�+ W��Ӂ]�*|f,/e6ot�8��?�mGVWa���������2LD��'ƾ ���鐣���7��
�c2�E�u�<�u��������j2�e�8��|p�?i ����v;A���ᇹV�����UC���S�i��9�N�nR9NR"�X+�E�W�� ��A�����>eϼ:C*S�����{˦��9�O=v�8���>������n�[�f�G�I<q����.3/wC��v�>�ff��+vb7���SHťQ�Q<�f<�NB������VR�,����Yh�anH�Q�l�J����(K{ݏ���}�f����rz���"c��Ǯ{;b�.�f���h��轖�վ {ЯT�>��ľ�f����u3�
��7�E�q�dv-�E}��Oe�|�oˢ�ӷ��/t9�m]��#~s�2�V�9����G�D}��i$�|)��j�E�!��VF��>��s���${ӈ-��jwS>��d�z5D�:��������f=�D`��A��E]{���ӑ�_��l�^��7�ꛛUNu׺�����҅����C'p�_�S�]��pg�鋁�Ta�tuy|9>Ź"z1�0�'#@���G��d��ŀ���a��-7KH>��Tܕcf��b\z(
�����c�^G�ta@��.ז��WJ���
q���~v-��lf/>�4�Pp�G�~4~�b�����-e9]���Ͷ�BH��;��c�R�X���S:p_�۱�Ә}�|e��q3�z]�?j����^���>C����W����3P�~�7
�V�R�L]lSw'�;��v^v��!��<o�ؠ�G���B��(S��rk��\j��z>��/K����ʿVs�={��)�j������H�2A��Ø�EO	q��]
��Ŭm�2^�����&��{�:���~��o���	��=��V�u���ѱ�`O	��۫G����r���=�nO�,�.��Bo�ZG��d������n����C��~������?x����Y�������1����4���z��<�3�x3�/Tb�2�{��G{Λ=��k8f����P�-6���9Al�9��;��ܩi�#6�}G�6���K�n��@�������&ߥ���������8;fbA����?AȎço��'����Q��W	b�q��:w�/�S��G,��
�cݨ�#p
�T Ec�bb�S��W�Z�;�,�zk�0ʊ������r�ۅ���J~���jz9����iV�B�$oNZGy��z �Qx�����Ө��eX�"6��SG��H		޿ ���١��bi�^������;EԼ�wD�`����^GG\��iP��o���������ң �{�Z+ݻ�^�bG
I\�|��?Pٛ��=5@bTTW�zTU��6z�鵏���Z�V�������t������M��p��a��}�X�D٘����	�a���EA Jbo<�����w>�[s޶�#p-�!�:���w�^g�Ve�&��r��{keVK��.�3C�����hz�_^��`'�V���ĸ�	S��7V�SU�O�W�6ש�q�q�w{�촇v��>-�!#��5��6�ޑ�����/�Xd_)�l�M�Á�۫���{�&��h�� }�dkU4��N&�TP�%L��V��v�3)���u������C�fI�yx�w���  j�����X^�-�=�s
�V��1+A���5b7%��r��t��n�J)�M+��:�el'n6�:tY[*�`[����M~�>�""!�N&WY�3���2�}� �q��.7�*����p��ý+����[6����QϨ!�l��!i���W/��o�H���:}9%����S�R�Dm��\!��0��5��dDTt�6�g��Z�ү"˛e?4-X{jE��#`�~;�����
�g�RbB�=gޭ�mow��z�G?�ע�ϻULP�.:JF�晠�������J����<��[c}�[7q��`��=������j��U�v�ؼR�����ãa9�6�9aM�h�'׎�ML����������c$w������b���+�p�R�Fg���Q�U,7�xg��$�Y;� �?�o��d��g�����ml��=C��'��to�c�����8p�a铗ӵ��g/�9�i��z���~νs�鈯��]K�w1h=~B\(�T�j9�0�XZ�DO[>�b"#����^>�B`Cup|ؠ�3J5�\XG"G�?h��������U�����f)r��5y��T+c��f��[�nm���!�5*H��N#|k�B�����´ج���MЬ�Q�'&���:�73�`��x��2w3m��U>���͇�5RA�{.L
����Mft�r�Ss�X������Ƃe�;ir����J���?E����F��cx���oKת����aY�ҩ�
+��>N���+�����]����0�����ԏݸe��o>�N+��ԑ��!��j�Pñ��M�I�.�t�uL��.U���$�r+�p2�+#�����lߣȶ��b_����mW�ͬ�k���k��l�����#�>��mN���h6�l�E��,3��-�C.��0��}v򎮎>�23R�A`!=�追s�]��"a��&�q�6�_���qO����h�j+r�8y4�������;�{7��z�[ϩځq=�z,u�UK��A�(J��S�"��h�F�ͥu�㯴�s1���Î%Cg��e�ɻ��v��NנW��ȗ�����t��1�v�i=ȳ({�*=2�Olqʗ�]��zݸ~�p�4-�PGg8�e���'&��Dg�L���y��ݰ��ŉ�0�=��Al-�P�/;���t٬*�h����OQ�����S�dI˭X����i}F��>,} >9%�6:��Y�X��m�`b��b�^�l�{{z�3�̛U���{�9�<��W0)&"{�|h��ڀTq!�#����W���4��1�z$:� Z]�!U�Y��U�ݩ!�\�WE��p5cįZ2�S�	�vv�i�˅�&�@e=ٗ� �����[+����8ˇ�C�^]�BX���$�q��,�ۺR,���4���R��x��)}�=�]���}�R�M���k��ٻ�t2ga���U�h�Tf��}�G�u<(�N0�)~ɏ��:}�<5Ldz����i �v:�����GF��}]�ED�D��6Ƌ�^��������r���r��X+���J��@<'�4�T���3u�Vo��tkȠ��?]D>����a`��z_����n�X}#̨�xB������^ţ��n��P���bn����!�������	M#����*��D�*���S�;�[y���c�܆�E٢g�Ȥ����>��k+a�}�q}���6�q蜤�u�b�`28ysf���z���NC��X~��" ���S������9���۲�3k��]ڝڱ���W������.
<����t��rX����H�["��޼E�̮�W���8�B���;��l���Ξ7�F�]ӟ=�!���Zn��{z�����]Y�bn=<*T`h�{�IU����]�e�(��Cq;U:X�ϹPp����[8)���������U�������%���]���S���x8������P�:��ĸ]
i����݌>����"6*dl�`^��\��̮�/,�vÛd��CzX�;
����F�X�g���\PQ���ٍ����j:(r��~[l:�[�xI���ރ�H	��+O�K5�D�]݋���lX8��T,����������ɷ|�e���{i`{��Dq�N��K��dZ�"ne�(��ڊ�
E�����w�{����	����<���j'��~�?t?"G�?V*�.~@<�V-A���VOz�{]�r���.�>�#v�#>��{��Л\=�j.��Y�������5�o�/7�Z�!V�6M	c2��
��`�v�M��)ַql"�j@�z�t��[U�0:˽a�y���R.����oYއU���Ҧ�mf�4T��9b�l��c܍ËV�r(��H���76-��E�����s�C�cU�}ϩ��$Wl���Q�;9l���v�}��^X���ep���4�5i@�w�����c�7��n9M"+��rZ)坻�}w�o�h��z/6ϭ�]�Ǘ6uM3�'Uk�*bf��"3Z%��w�����Ӂ���.�|��c'�x���q{w^�a�����;�������[�k��}�~gSd���G�����こ�G�W��0<"���#&=^����f?@���`�ۤQ2��������@p���r	:���e�7�D�{w�2�>�v�_>D�o�l+�V����{F�ף�;��}��������ʲ&}3��q#��.vJ�l:/,��azd�x_�׾6���s��U���}`9뷱���	��騭*�Ѫ%}�
n�kx�f�%����ǎ:#��Z}��M�"��Rw�N*�����u���
۷�[,�ՎV�ܦ?''��+.�N���'�փw����"
hx����ݾh�^;��h]��xX8p�`?x��Zp���;35��JU(�*��bq��Nr,=���"��;M(0����i
�(|s�-j�p�d>�
��s�1���8�o����Mq�r�nE���q54^�M4n�1.�l�W2�D��'i�\�4�H���G6���DPyIe #'+bd�y	��dc���-��T��AjB�]d�]�k�d�uF�CNw��5�}�����h|���'�⽧\>��9�p�狄�e>�{|�:^��2g�݁��e��l�r��90?o1���b#��7U�0�4��E^���^�v��l��z�h0u��cM���<n�I7.�c�<r'|Kנw��mDae|���W�E�(��Rr7*n?�K�Po{�4d�Y�2��n���z���}�����]��V�K�Fu���P	@���5Ŋݙto@�un�POוT=��-qvw{(����f-��;-�y�X�n����!u1P0YG$��� �tTW�Q9�QW�c]�5M�HW�cO>����o�i�B�Q��'9?w��˼��%c�#��J;^C�wZ-B��FB{��9�,�S�;
X��i`�L)�h��0`�!��4��<����҂(ᵒVi,�H�E:rpIE�o������ݮH<�8C��@�C�9:	#�:��r�^^�"+����;�����������f�dg�y��v[��w�������KS��;η#{Q�۬��̨(o���k���ޛU�����+5O{��ϑ���cm�]��q�A��VQ^gkV�v�$!Yg<���'~!�G���{�4�S����s��N�+N����nБ�8�G_��n����_>zB|���[���{x��Cm$�ɴ(\nO-� Btt]f�DyY$�}����>M�A{���p[c��:N��鵗�j��/dյ�̂��K��[l���T=����^N����קe��;��z���'}����vv�ED&���D@?��z<�'���1�\��U
���+��ٱ�sK�Z���*�v�1T
��\ܶ�l��	�{R<3x	�5�?a�?}�g�g�90�|F6�}����UdTq�����DԄ�މ/*���M����f�-[�j4��~�}��;V�y�{�vF�VeJ64�:b=S*��P��lP�azܜ�L��	����6k;/ʻf��+����c�s)�*/�Di�3����K�{���Gc{RV�p(n�;�ˉ��x�w>�)���M�N3щʅa�9=Ȣ��Ё?����wz��뼉��[��:����=�1���#_z�K~��� �c����h���,1=1�<9�1��y�pp4|ړ��z���c��g]��x;���zy�H�jTs��#�9 �OŚs�d�ı�����S>�b0��28KF����ꘄi{<�=��>��[쿬R}��j��O7���}z���8�f���Ȉ,9tKF��M��}�0ʿ�hDmw����)��>��h���EV����v�hB������&�E��&|:h�Dy�X�uϸ�	���=�u��Շ5lI�}����a���GF�fnO_���TL_�zTU��6~>J��}��`Pd��C�c���X;+�������N��J6酲.���j��&��n�K��'j���b�<�zl��ML��r]�y(W�3q��@��{���EzW�w�pp����Ƒ{s��Y�ZI���u
�����ּ�cm�9m�Cِ?G�G�
6�I�Ѻ* /�e{����E�k����p��a��l�>�Xf+�5F	託�OJئ�:��'�P����O�vO2��I��:�޸�Ŵ�;�^�^�l{k��*̿r�[.r�w�]U�~J���Ē�#�:q��^���
w��+f��b\f��1,cul��z�G�5�������[�}��0�F���𚀽qT��A�;��Xdh�5�>����Mz�\ϯ�մ�����:n�f|&w��|r
5�Ƞ�Ɠ(�{�EK����PB�Ը��Y��UU˭��UعG\�9��˚E���\&�8��;����/��!LFEKu2�!n8�A�۬�.�M����e�N}﹘�T�ƻV��Sl��"�=�����6_O\	�	����N�[Y�6灉�w�ŒZ�q����lya�����\t�	N3�Ą���ճP%��	ۂ]�ja����4�{w����r№&a����\wj����M����zۭ��,�֯yǋf2ߺ�\]Z���LIp`~����� ��Ra�V:�_�иV+�foSeF=T��
���K�?�����'�H�JU�P�m�g�!a��hO��H��������vD�[*�<���4�Ƙ�mC��ދ�iV�B��\;Caͼ�����3S9���ZLdZ�a�������7��Ĺ؜Z��p��6(;ٹZ༛����蜧�M�>�����e��9�k����ۨ��b�~�G@�#RcKF��8�ڬc���t]:�]�J�oR�fO@!��8�������u랗�_bLut�����	p�>'c5L���z�E��MU��+�zX)��CUpbC���_�����G"x��E����z�L~�l],c�6F�~n<�z���HQ�v�i�gR�7X�[u�jT�Ah�F��W�Тs��e�����w���''�C�=��exuף��wW��b�����#�C�I�v3�
���Pʍ93���[�5o�26���gtN)����=Gtg��5zgc�[X^�!��ߩ������^dbY���n�3�ɤ�K4�ζ��G�	�l�jwN@~���l�E��a����r��x�3D�9sc��W7���^�\d�����=��\�y" ��e|0M"�r.w�v�>�ª��j�_����:�ɯ��Z����-�e�*��jŇ��E���/�����UDa�ު˺����>�Vyx_Lb�,�F���*i�����d_};^�]�ȗc���FagS�����SoA[90�٪�u-Yn�Q��}�^|��E$>���:���D�|��	�NѮ��ʵ�&�މ<��d���7'��达��ݿ�sN�ā�X��n�ӗ	&N�4���G��OK��q[m���Ǵh�e�[�N�ʶމwVM:�b����\~�����!X-mw�9�G���t�#�;�a���U6�c��d8O>�BѰ�+>��Q�
�;P���)%�ޮ�sf`!�'�BK�T�߂�ם�gT�kR���Ǫ�ȫF�*�(��#��gk�=�/�\˃ƀ �'���IB;����V+��Xہx��=�9�Ȏ�\�en�Wq}f�iC���ƈ��"�'ƈ>���T�q��\��+��P��~���<y�Ioyo��o=�-���~��w�/`8�cÎgH�F�\��R�I\�a���\�g�M����֬cf_����nR9�9D)P��G*��D�ٸ�zH����vϛ]���G�]D-����>\݇�U�~����n�=#ASD/\�\fm��5��7�}�;q�%�= �.��?��!2�9o�@߂SH�S�w�US�&9��C�y��ֿZp�����4�Q(2&Ɖ�5u6Ϡg�Y[{���N f��$�ǭ�"�Ub������,Ci��}���f���Ȉ#�H��19��N��wl*�_��&���R���&�3W�&�����;�KT,��#��ݓ?x)�(vr�ۓN����g���������Q�tx=5m��%]׆��eWrz����us^����3�^����\�˯��}�47 �v1f��8�M:&%���������L��2sU�G�����ˍ���׵PG��f?7<8����_�C'p���9%��2<%@���Ez���]�1s����}��޻����\��u5�N��;~��Xݮ �N@�5�`��K��Y7��͗���*"��\b���{�bܞ����q��r����l�>��}�VnLZ��Yb<�$	�b!� �S���������5w��#��~�b��"�/���n�1�ܜ��������n����g	��'�9qR8#c�#s��ڤ��Fj$��s��z�nn�پ��t�w�E�ը����R����O��z�.�}s��lP�/[�`�?iE���9���R��:��"����u�jzʋ2#M �Ø��q^�^�zxmz}g|Ϻ<A�9�J�>�~�b����"��+���r�X}NOC�$[ �@��`�o�3��/L�ՋҶ+���T�j��_�j��Ғ��nݎ�a�Fq��g��M^=�b��(z^¨��]˻�7|�L@��~ �v��\j����\���jR9d}����.e�z������"��\������jI0���h#8a:�D�ՒP���^)�LҤ9u���n�n&g1�k�t�j��9�Z�*#�s��� �,l]��lT(ǵ6�D�@����GJo�
�k��f���Р)�v.�m����td���4����'�G�G���D%ˁ���1[��Ș�P�)��Ͼ�\P�LF���ud5.�%z��J����{J3t��S�۝MC�ʈV�h����t�z���>�enșJ�u03��}Y�j��Ǜ�x/}8ą�|�B��aW�4K�X�|��ӯ#�uϸ���
�˕}�����!	�v�l�K`���!�i\�i~��7'��bTTPcҢ'�(�z�w8�"̓���3�g��v��>{��ݮ�%z\�'�_:D���g�q�34��p�L;��Y�n���ٝ��a��F.�^�����g�f�7q�i�x� 8o��C�^e��O�ۦ���{�]ە�םý�tϘt,��2$`-�z��;��l�ռ�8���qcul�#�z6���o$��-�>=��{��9�xgNG��)"�*`?\U����B��;��,2,{�JFIY��,ǝs�{e�۫�-S������/�Af������4�G�EK��w���O�B4�$��vo��R���3��2�_t.�ݸ�;�Ѡ�rK����1��Q�����d�[#w�7	��k.�NM�R9������-Z�"�ŁF�Eg\�߼ �>މg���t*��wx}��z����3�����"�\���v/V�5FÓ��Ń�k\�%�DD���6E$T�iC��.��pA�S�M���] K�#���y��=X��L��NH��v���M���еa���6���v�M�7&��zD��'MD8�ӑ]#�qĽ��3�B9{.s��IH�<�f�FƧC���p&EFk��y^X�w:o{i���;�gc�8��0����q���3ʚ2�#a����y�x)n�{�׽��d�R4L1�p`Hc�:q�&�}v/����µ��@�<����T�z��d�7za�:[cm�z�w5����~뺈���1�X@�	@�4$Ɩ���1�lv�۳92�������q�y�2�&;���j���j�S}�=��_u�1�:`F��4��Q^�R��[��� �Lm��ͱVAi�n �6y��X.���腂���6(=Lҍ���� G��<f�a�a-�{����z�k�`z���இBx;�G[�n+u����D8h�#�-��M�S��;N.������k���,��`���3ss�^0��\a���$v�ާ��;�{�%���[�{/J��f��ď5�߲Y�e.��9�'s��ţ5]ߎ��=Glߢ����,C��Y�����DFD�?��C~�ނ3��4/����y{ޜ���f/�je�8�՛_yy5��}�{�d5h-^�Q�)�(���sC�Ӭ� �ͱX(l
��[�F��c7�-6uTM<qnܯ���=�����"�ȹ-{��<�����	˭�.M��Z����聗��Vgv:fX���z�k��"���ɑ�H�xKf��t��w�D7��y�"���ˌn�m�wp̜��OC���f��7װo�=��\�c�Xr2��4���"��Of�\����˃LV��_����!��)�^=v-�jŇ��E��^f�+���u��e������Aצi�<�_z�!C�J:/�\6p4��݌x)�da��"�^�W�e������2�;��n����ŉد���6��wޣGyLǆ��p���>����X��J��rO�A(�U�+�U®czD�O����_]��Ȩv��Pκl��!�Ī�����o9�v��B��F������<`G��>5%�7��eb��1G׶�Z�ܐzcW��Uc�����f����t�[[s��b;����F��9p�77Ż�1��W4��I^�W��}�_�}��8+S��e�
���v/�di ��P�v:#"a��^��ݚ��E|,�ܡ��k����;>����nR9�DsX+���J�"�ى�F�91�	>�0⓴f���{�=q賟�v��h�|��\�6$��&T����a���m��o�-���ɦx�z��i���x���?|��?{M�g�&7�s�Y�j��{j� �W�8��8�F��Ca�e!JE�ͭ�D؊�*�d+�&�?D}G�4�̓�(A��L��m�ȸ-���Qlvہ�akv}5��7Q�wP��H�7�7u�]Oj��k����;�D��6A�%@�3�=��!��&^Dr;������X�F��C�9�z�Z�9�.�/=s�ļ��Y4�eU���QG��xn�0!`�>���œc���[;"mzOw��� �`iF�dh��n�3
�8���r*��Q��N��~ݰ�M�W6��G�ˮ:ϯ�x�Zӈ�a�K�~�Ł�_�Y;����9%�8<%@��Ȭ�k���U�m>̫�|S��V�FE�7���b��b�7k�6�z��*�n��m�_�$xY9�ǝ�Cb�GI�3�U��V�GE���8�)�ź�k`��Ti��C�)�oB~z��7ݯp�0�A�9ȦE0}`EHlX�_�E����p��-9pR����H����!�z�N�go�ދ�&�"e�|L�/[�"� ��މW߲���̢��
��]�Uqxq?6q���+m[�`��ʖoAؠ�G�p�!Xb�2�ʋ�����*,�(N׭�O�=���01 �����=���h�9�h�ΰ�?�=q}�
���Գ.E]���6�g��2KR��>ɽ���Jv��}���3k`�(1xڪ��&�p1��J�j�hI���q��n�˺C�	>_�����Z�n��� \{菾�;��K�1����>�e@Ʈ�/�f�[�s`)�*/�Di�ĀØ�E}<%��Ő�b���{׾}��e�ƿX��mI��I���z*}NOE�EV�w O�V8|N��D�h>�c�vǦ�Q��ĸj��Z��E�[c=��IO��]ӡ�y�Fq�p��ƌ�S0���f���a���?Y�W�W��E��;��^���H圏ΔZ��}�d7)��&)+�ht�!��jLiq�1���VC�N�,�����W6]��n��w?�Ņ�[�b6 �JDA�:%�C�7�Q��q7%j�]>\���˕�k`��)�s� o�ą������6���&aq"fX�Df���[�#��7��y
�ߵ�_�_���b?Pݿ@�&�R�-�k�c����l�����bTT'=��P��T��]�O��`��|rĵB;l*u8����'=.��a��g�z�`��o���_�V޺��X�}�$��lK���碮�^����}\o��VE�M�F��b�u�-��b&@��
a���me���H���@,^�Z1s��]��|��SZ�����:/�.a�p�Eg��>����b���fHpq��û�Mf����a���o5U� IfP"�N�(L��C������G�u~�6�Q"���FxO:��W.(`9���f(�I�k�Y���×������[���i�`��Aߵ���O�o�~yzh�W�!1�~1��[����;/q��G��bQ�[y��j6�؛�f�jɣ�u��廢��U�r��k����	�0v	����a����w�톙<����"1�|yy{ޝ�����ݞ��^@�rf�f}�,#d�Ϙr�66��V����6^�ў�/.��\��OMSW{*&{gTn�Q)�iJt��v��1��4�ѷ�D��wrS�<���V��M�ť��uUD�um��w��bC�*ϰ�xiN_m(q6��(�6� ��w÷E+�"�an���A��f�g��
M�^�.����л�>kfl�:�w�����>�z	g�7/Cܱ��ptfߓ{dkt{:N��}�I����[�m�����t�R����y6O?}�I1�
�=FU��8'u�{Ӟ��-J�w7ۨ���a=!ࡀ��/�b��=�������(�R�'��9ؘ��z�B��3���(/���ᖬ?+'��{���Y�=�$և� �x���"�e���w���gjl�)Kknai W�{����{���Iw����{}�r��v�S���/CqhA��nƎt�P^���O/s�O����|!�@˾K&�� S�8.֣�7��2��V����g���Q�	t�F����S����X���49�%y�����ۛ��%�z��^3w��i��kEE�1����A07���z�}�����$���lE����w��3���w�<ջ���h�$|���9�b�
�����{�؂�H�|^v��;u3Th���0�3JA�m�5+[�2P��/3%���8�P�:%M޺ʐZǛ��!�h\*1r`~8��=���4ޑ�3nт��r@we`�uf���	9��]�,I��̕��ⴭ{��{�3u1��3������{S�tI<���Ȋx�m��ܤx��(cU��WL��L�W;�i����?Ww�ᡫ�&Xxx��:�x�M�r��xb/�sOw-�wE��+Լ0̾��W���j>㺟zg�{��mQ��d0RM���W����e6"���Q`*�p	�.�^�8*�*�����[t��6��>[�<����-j61�;l��\Qc�ۆ��U���:���ըgNvC�`�V�L��J���<4gV�Ӧ��܅�2ۘ*(ULX�b��������3�v\�k�q��Gܽ��hƗxG��S���c�	��s�,�sNSw:����o�2�{BQ���j�Xf�����oi��	����;����=p�U��P�8��xG�؇J�ݘVF���2�A(,�O�@ҹ�FTL}�3�=����I""�`�ADN�{uy������+˾y�q�"wG�{wD��[i9���yg{iﷺ+{w����e����S۬�;�.8�����+NN���w���w�^�c^���,�m��]���k��g�>�Nyh"}��>o�o4G��o�����OkN��>�;���Ȟn��n�/q^w���9����^�ﶂ�3�j���o����}��
$+��� ��M���h����y�vV�w|��ö�^�Z��K�88,��<��;�ϓh[wlo���M{h#����l�w����v���+#������/^ڕǝ��}�pM�2�}�^sn��	��5�{{�]����f�D������}��ͣ����_Kf6�,�"�"�f��g�YMZ�[�Ͳ���^۠	��n����zO5�ZC��:"Aol�}�x�l���ݴ��i������{�a�E�XB�t�7��)�/1J��ng5�

[b�ܤUK���L b�!^:Y٢6ܶ�x(c�b���qX&j�Ǚ�]�G� ��3��9�.ۮ�kM�Y��u&~�#"pf�����ϩ��o �������K����D�څ�ڲ�<;���|]7^�k��9fY���d0�z�&�?l�G�����س�r}���Cv���}9��q?MF��7W5n3&w���pY��d"���1���nu�+����ŗ|�q��c�N�7�4�f�Z�B�[n�dd﫢<nK��?
b27F>������k{��iϺ\Bc�HC���K���t��T�)�O�Z{Wa|�|�~�R�_A�>:��X+�f��Kc��b~��bTu��HG_mz-��f;�f�S��q!"�|��R'_#޺c;ځo�����9�蘳1��ǭ�]t2+�|pu��;>�wўRј?H�tn�.�e�^�M���xӪ�!ޓvt��wL3��]���]����"Ǽ��;�Z���^�#���s��<7�<���wQ����6`A�(D�ih�u�q�-�_Ew����U+�~,o?�Ӂ����%���
S}�`?uc������G�A��
��Cq]��
���hzbI8���
Ӯ@�v�a8Z��g�S*=�:��/�^�*@��l-��R}�1�ʊʋ{�V��S��y��6��AE�"���q���/�l3+��9$�t��F��8=�Vn�{�U��� �Cȡ��Ú�CC3a�?����Ea8��f��s�z�V�X<��!(x��4iF���	������r�#�7�r�҅׃�a�������~��О�Ƃ�u���3�C�J��h��Q軟`-v2��:U_m�����*.o�~�����{�X�?7�\A#�f�<��X�D���2���쓺O"��M�T��JG��5�z�вg�ȪO�O�9Y�3�6k���ފ�g9�����u9z�5ЏC�\"�%^�~��;�248�3�H��-�}�;� ?}w�y�G���E]G��^�vc�7��{,q�ǲ�6�T+��Ox�=F��"de��^��,ݜ�q�rC>��I�[�nz�O��:e�~89M�޺�;P.-��/+n�`Y���a�wnA��c�<�w�f�9����*V����P�S��2᳟4�ϓv1�;l�����'��
��z߲�����91A	�PZPڔ!��Q�"��*���n�58M�doUs1�1Ad>'�U�҇;V�/A����1�03G�JO����� ��&�u�t٨��n�����^���<�L\f�@�#j�l��X�*ڮU�n�Xk��UP,䅛�+�،���sjj����vKx���nlBՏ�{a�<������v��&�ù��{�s��wOb� y�d��!���Q�D�b^��٤O{�� ��� 
+}��ֶ��ߪ=�?3!E ��k�h��<h}!�(Gq�4�Я�-(�a�H�Yz|�u�v��)���a��|�
�[s�fI��ޓ�@��ڀ\u}2r:)�#=���AUכ�={��Y[YB��o�N��]�<��E���|p� q ��=n��㯳�UԻ��]���*�.\;렣o�Xǁ�= v��l�n%��X���V:�5�I\n׫۾:�=؄��GT_�G��!n��jE�n������gVǽ�='<��N@�aa>	^���^z��,9tK�?d�o�OxnTCe��Du���)�cE{��K3�6���k�	o��;A�^��dhkrk�
Eh>G�]M��7; ;� OUNC��g8�2��-^hޛ23^�2ӡ�	�b)�S��;�3
���"�18���z�77�:�׮��狫��3^QQȯ��ůK�~���W�VN�q}S�]��� �e�ʧ�Cڀk��=�&=�Q�9�C�Q c��������[,C������q��zeM�P2ע�ob5��6*L\���bMĉT�fxü7�<��d�{sN�w��h���K��O����,c܄x���tpʠ�����f:���Xw�s[�f�^�F!�XOҦǭ�`�o����ka2�@;
���N�%��uɗt�63U]���[&?G�}�!WpZ����ѱC�OE}�\b���x+n���X��ʃ�x݋g)��g^�yS�Uh�[S���on�wKXn*�ó�b~6r	@��R����,S���/�~.�R��k1k�evҞ;Ϡd?����>�x�Ӿ3����f�Ƅ����HA���C=�Td��C��3d�ji�GZ�:�fj/��.m[�o����wAؚ
b<K���u��#���bj�kܽ�9�'��nMsh��h��P�=W1�S�TY"4� �H,:��y���	����|
$�q��܏O�<����䋰1;�+�����B�����H+H>�؇�.��oz=��N�pX.7ji�W^��֭���)+���.�[��l?H�7�݅G�t���yա��H,U�#A� 9�H+O^�\kλQ�ܺ�C�~U�M���z�Z\6)�s�=�TF��9 ��P��H,G$Ɨ꘍��VC��ۄ='6T4j#���!�������u�x�J���]��)�)�
A�ѯTޝGîa�H���z�6� �!�fiH�S9��,�$���)F�K�Wi�ι8)T����"���f�*������͸t��p 
s�uj���:&��d�3bX�[�F���#bE���V�v��cۛ5kp�7���;GM�6��H(J�Ę�l G��;_�{��;�*��������6�SR�7
,v	0����
� h>DWމ��t�F]l�����y��6�̦�Kv�ɴ��lĆ+��P����7'���;ur�T�p�Fn�����9:���c'������\�^]n:/��w6��v��.�����pz�n)�}��Z��e��f��;8)QB���+�]�����s�{�2s�z'�X���)ʼS���6ZC�uk!�ΊBï�V�瑵Vb�D�)����`�{��P�S�h��UYO�=�giw�Ő��ę\�z3���O�o�7�Q����a��xM@~�Cފe\t\��K8��,,��Kw�}�4��Cgup�SV�2g|}8�j�"��s4�G��$�U1ڨ:���3:;������(/S�c�i��#,���	�N.�v8NI|~t����0"r��k=L?L���d�׹�����\���m���O�hZ��� Ņ��}V̨@lɽ�?<��+�/��'��0Tn����NE"��������	y�	 @��.��6��7�CT�'��܄r�Un�sj�U{�^hm�}� ���xt���
:���}�+
r⧲sX������v��n2/Q�ĻL���{j�f�Q5w�&q����zh�h��$n�./>�ߑW
�0�?�n���8�ܹg[�����GȜ���ճ����"y�=��P�;$�vg�����q���g��%K=SX�vp	��M��E��ͳ�r:&'�`����������a��]���H�@ͯng`�ʹ-qE#�.�e3�����]�+DxW���#�l�vL�=�rLih�]��=�FvM��SW{��O=j�6e�������W׹Jo����bLut������ʦ5ډ����]������h�\�=kU�ֶ�!��>lP{a9��<0�F~l�^���`��bBrHЧ��Z{Eu�{�#M��Q7�J���!Eq��q��4��X֖8O�ϫ�+ZۋUq�Qs(�b��W�=�,W��Glͧ}�!�^Y#����^�lkrϲv'�ޣ��c�a�{B��DM�'�$T�d4|.��ٿC��08����r��`z���6�D(�ߩ��گA����w���q�p"=�[>���ȥ*Up樇�U��{��s7�.b��E�r�;K�$8V�^�G��xz�$��$D0��ǹ�����i�:��O�r��_퇭}��:?�y�{�6�x��ݮt��D�3@�?go�_L����?,���o��唎�v����zg����Dvx�9�^ǆ���}f/*b`��V:.Ð�,!7:q0%֘�u[�f�L+�D�«b8��±q4v�����_���Ŏ�l(���<K���6�z�W:v�TX{��u��*�/L�\-��ھwMoo��}�Ĩ�~�u��T�1o��
�S��2᳀��Zn�����!��
^Ý���z(�	g)[��V:�H���*J`���>�0�p�S���p���	���:B�}�w�/u�z���,&���XW�������?hb}%z�]�ȨkΦ5�w�;0O�U����y�t��O]d&_�2:)�46�[WƬL�4>�`�ƾ��wsl��J"'l�s� �v�b������^�b������>3��ٴ�BMm�
��&#�O�}P���U�OE�4�T��3��f�Nz:p���M����٨��'j�ut;Ǘ�+�sؾ8A�#������]vWw�i����'�q�@Hr���toyP�ÚzG`�����G$g���~��#�[}����e�i��N1r h?D0�F	ȫu�����s�U�m�E{b�9/���ߍggk���w
t�#h����B��
A�\ɪ���D6^}�QK}j ��]-ә���7�x��u��1�f#[Nct	�>�HoW�(��H7�e�wr���%�m�Vc��b*[�P�*D�˦snL�b�Ĥ�R���>N�|�� чs|`4M�Ӫ��j�dR����u�]���3������};Y��^
�%�u$��b�5�-͍@��b���Q�Ҫ�����W�2
5��&XR*�Qg�7/}F`,���(��l�Tt�����G��
������܆"�U1AxNC��Xf숂<�������L>:k��ŅN����ՙY���w8�F=������a�o���_�Y;��I�/�Aڸ?t���{ݞ�7�gC���B�z����h
ۨȱ��=8�X�a��-`n�l	޿@�&�׉ݠ�3e����5����>F��*2�QC�"�ƹ�m}w�qѝ,
q�	Pp�cv-�<��㱙-m�s����a0�}�o���W�rO�9ȦE k�"�6/�!�y�E��N�va����vŻ�����r�6ۧŉi������;�,���f�Ƅ�����3ނ�wZ�8�(X�Dڽ�oo�7{���ڧ��3���Vڷ���"�̩f��aTD��>+:�C|��#j*����]w��b9��
w޷&�Λe�Ʈ�/��.z�c��*4#L��+F�gL����v��y���6��}t+}b�|�ܑv1;�6��ϓ�
�S��2(��8&i��:�tp�Wnz�r�dc\�$ Ʉ"����>�~�����"}�D��O�����m�E�bѡ7���[��q��:&��ax�<5���Ɩ+N*A�Mn37.L��T��r�H���ޔ"~�O�<w��d�v�P�}������[�L�O�"q�bv��/G���_�V����&���yn�q�Ⱦ��3N����}��[�9Le�g�A��P:~�Azz�۫�}T���{��yѹ�s�q>�$��o���{�=�����)�PT A���1\o��Q�]��L�C+iW�$VFH׾:������&!K���U�x��U�k��6 ��R"8"h���֝F�od�}����k��WY9�z�D:ԑ���@�BB������Qc�I�]4L�
���s*{X����=��`kɫ�Ǩ�M+�v��!)l�%�0�:0�_l���Hzs�[1�
=r��eS���z/ӓ���]NBg�ޛ\��twk���N���1|��N�,,����-�ۮ�ϋk�5pOEE��������}����;��̡�=��:S�j5bK��Ur�=�P� �����q��xe��O���Z>�O���
w��ٿ��	ȅ4}�;g�ގ|3'7C��5�qc�fZ���.�x��xe��#;�j����z+�����~��WY���.ñ,=�w�f��J��ךz9�S����p�l��:{W�������zy�b��L�V�w�2K�V��2�:=�{-��?��b�4�������1h��v[��԰f� ��\&�{5 �E�*͝s�lY�l2+N�����{rs7� R�OC����7W)�q�&w��|r4,�2()q�-ǌ��~]��{u��Ƥ�S�*z���ޥ���e�⦙z�T.�q�w'�G�Ӓ^�4�j���L�}�f����S�@JU��!	l�B�9"���g�M���hZ�ځ�U�`����n���Vfv��YS���@��<���.6�ۮ��mz-Z�b�̈́��=J�=Q�����_���{��F���U�K���'�@s�E	(q6���οU�`�w�(z�Ww��*��#J0���~����=���9jl����@c�*��5&��Y��FguU
�cT��������aӿF`�I��R�xW��Dz�p����@�	���j�4b=^���=�J�/�0ʰ��ǟ9��B������)��G���I���`D�Y�yӏ�2��H��f���3���:�u�3ֵX=am�BM@|�NmC�\oM�tx���_�v�>����}%�.+�t��WP�o;�G��qMͣ	LB�����<&6��9�0bq�����hV�ݘa�Ǎ\�UQ3���y��N�	��I�8j'W*P�{*�/k$c�t�\�J�����yh��ޅn�Z�բ��ȞC���.fI�z)�uC.S�Z�9إ�b�O����t��>j,
�E%Yer^=�O���������.־��]�N���;��z�j���K;�j���5���p�j�K���v盀� k�$[7����w��nzP��Õ����5Ҟ����ݦkӉ+J̸�N�ZoVU�*5k )j���(��8,�j�ݾ
?u��ǵ@��!J�ﻼ��^1q{�ǹ]o�I�5�E�y?y�aZ�\[���ae,�]�wo�������3�5��pnN�ǧ>�S43V8��E���lN�dc�'^:�>'F\\�N<���7޽<���=1�f^����,�\�ET�n�71(`(be�e�F.�`�K oU�^�����$�@ZWg�����F�.�W���-�e׸���5` -:���`�$��
����DP&�~fy���,�]�N}ױ�����$Ҹ����(�����uՑ�s9�Ӛ2���x���)�	�^�ӆsr�8�$�V/9.q�=���4T!@�*�jB����q����C�e�z�/9�M�ǚ������1��z�9����/y��5ÛsEB+����k�K�|N�8���@ܘ������i�L��'.ս�x�~��c����i��oy���Q	�d9����3� �͑햷�;�k�r�.n�h��nd�����D�s�M�a�.�CO�w��.�X�G9�_N��y���+�[�Fnr�q��b�6���<�L,�᥎`�$����y�c%��X��<�a���������ǇM��X�a[�$ `"щ������zzxmX��߼�PY�}(�Ia��Ȯ��X�S���f�8���ui���]�\AE��$�������d�C���f^�o�HJ/��j��%{�r���\���Z���OM� 0�t=I\J��!��Ɨ���q�"gl���(�b�n��Bb�q�S��RJ��{"j[�Y��ס��o�L��f	�z�V����g�ag����ώ�І�"�zW.��"����s�>���D|�yf~��̰���������=�s�D
�����^[P��P�64�ݹ[Pٗ[�!RکsXmS�Sq���m��{���3������X�zw��4G���z<E�ۆݒ� �}��������<�T��y�[�f��hm]�2��S�S�F��9E��S����tl��`ʹp�໧������^�{���ud����x%��NzWW�|K��W5����ḵW6�^-�	Ek�)2�[J�����-k2��*bg2��k$�٥)Ⰲ�xL�``��S[���x��.��q�j0�'(����e�S�q�,a�;n� �)&v��91"��k#�o{����������� ��A �(y�u�Yh�Ԏ�;�6-,F[�m�L�����֞[ǽ�g72�Y�� ����ݍ�n8�9~}���F���.H5a�kim8�Xf��kG�B�me�ngmZ�����qm�Ν�Dm�9"H�ǽ�l�f�2�s��󷭅�m��r-��N���9�����y��L�3���۰	˖�d9��Sv�aC�JA[ZH��i�YvyVP^�(�љv�Ye���ݳf�f�mY��t�mĉ;��nm�:g_��m�5����Nv�m�-��M��]��R��t$��ٍ�I��Sn;-;C�=�=��mY�fMn�+I{^��gY)��r̢�����s��7׬�2�ݼ��z�/be��.�)��Q��JQsT�݇�ʭ�XԅZ�u��'��(A
�jl\��;/r�02����n��U�`�z�2�CLh�џ����u��+������'�}�yM�`%�;��B���%D�����o�5�VȢ|R w�9Y]�}|�[�3�6���i%��<}�������8��LE��z��C�H�,�'#��kl�mv�y���K��Џ�)���ڰ�}[?ȱ�,3�����*��^�G��e��$Dy�t�2���.���~���)�4��(����Qb}/����pr�e�z�[�JF���K��tqÎ|���K�6�>G޳5y��r�#.*[1{�1z�tX��FYi����פ����{�}=��Ī�
�ND���}?PB}%�EmJ���@F@s�s���}>;�Q"�u"�/x4گV���+K,��k�Q�w����$1�}%{�B�["���!�>�&�Y����9oa7�>�n����A�46���=�}�����ww�ھ�����7/������x����*|f/����N�+�������'�>������P\.��ί�Arc�B>|���5Ǻ�-��<�.j9;"����A���U������s�\0՜��j�%WF%i�.�26]C��J�`W{�e�ɍ��i�?nሞ�?��"�]tO^��I=r�3S���,�k��w�֬�9L��aJ�W���7HRJjM�~�_��gޭ����ô�x����ځcWC���
��v:,��G�ABD��4��{sv��v1���(!���tm��c4������P��wTZ�L�J*���^)���f�<�0�'k� �?D��� ��`m�C�� tZ��,��z]�B�\EM��g��mlw(����6/�G���*��D���.�����l���}�קn!a�kܽk�������75�,%Q��*���h��c�dk�4L��f(�՛���1�1Ֆ�}{>�:p���FgZ�X��qG�8����r�i4��G����p�������g[!�o�%��L�U������BZ�4Ҷ����a��C5Ed��9%�Լn��4�����r���s�ĸ����{׌�̮�Y�m�dX�t�[,Cǔ)kv��v6��0u����m����~Sr^���OG��K���,k���V�GmO���#�}���aZq�@�>#���4tk��X�][��o��A�ANE|Ȥ�����_�Ew�t}��ԅ�NF���n�&������;�˳2�Vl�Q�)�؃!d�f*�����-HU�YMZ^������p��������:]� Xy/a���Xq�#����ea�`�ͩی���r(��ϰ�.~�{8ӟ���z��=�Q9�E����A!wa�1`5���U�ct�8�-;�O��;�Y�>&��a�sDT����U��B��U��_f�ft1��w������
�l�3p��ո�qs*Y����{)!�3K<U{��v��{M��c�(C��
K���e�]R����W��saOYQ`�x��Gq`�����$�p
B=�ѕ2��~�p����k}b������^�g��
�}NOE!y^���vk��=�q�5�n��q诧��v��-T��\� �����i���Ug�/��Cr��c|_�Fi��hwH!��n}�� �=m�Ƽ�;y�.��ȏX���/h�c��,s��Y��R�������P��ä#�Liq^����]�m��u����_���;P�s�w>J����-vTB�8"d�R"8th��s1hMNY�����W�����W�B#h�4{>�?R�BB�#_{�M��xT£$�3G�s�gN�Y����4/@a��EuZ�2�������X�[��M�-�a�!�i\�ta�,��iM�+��Xו�7����x �j�5�y�^R#+1P��Rm^[���$`O�����feV(�9ɞ�+pra�&͹(���bt�ጽ�\ G�N�o@����g�����S�>�qs��`:��g�E5s��FN=��oEF��Ը\�}��*�F�R�' �;3[:�n�&;��?����(��<\T���ѿ��tX��"l/S��'�W�j5$���v��>��d��k�5�b��Pg����r⮽^½w_W��ǵ�q7�S	�?8�̻����.��գ��F��^��i/X6=���*̿u&|Ȝ�^�W��)��n38�C[�U}yg=�|,���U���݈O����C��[8)��]>���(���d0�z����p{�k�������2R޽B7��'�y�:�ޙa���;<�������gMߡК�fЪ����^y�'F��)���M�-G(�k�*\���A��R�t�2لe��иW�n�d`����#��CId���|�������N?��d9�ȯ�����m�vр���rEo[�π*m��ƅ���	^Q��>��νy�;=��d0�}�<~;�	�B~�P�~�q+>G�W/]��zU֑��3��4�#����o�h���U���l�����'���`��[SP��_��F.^0繸~���[L�N��y�~����s�l3�r:&'�`��:f�{�I�y86�x2}�֟E8�����W��R�-y��ិ�eD�ݝ�4�a��q��lKk8��!W�4��M�GRw]ӗ���Xޏw�q+<�n����1bm��iŤNK��lK<�غ��[G�z��4pF�CH�ru�bD9��d�ʭ���Jh6��$�Hai-��j�^Wxuиw�~���l�Ǫ��W��Dz����
�n��s�V�9��kc�a�$Ŗ���0�����8p�a�ĺ��ϩM�Z=��]bLvu3�bdO�S����/�3���"��*:�\o�aZ���!g��\ؐ����v��]=R��+]	����(ET_ƮL�%���R��R�������Ƈ�}��7X�^�2_���e�Q�~}^W���p��!���o�M�.��?0D�nr77=��{�X�8��b]�yX����w��g=�Q���6���sRcp�c7ưʱ�,�
EPb}jr�5�����J���Wz�3m|������ňq�������^�c�2=NF~�&��L;E�[��]�}��,eJ���w��5q�7��v0-�~"ao���{G���IN�pw����+7���k3s#��\\n��1ޝ�҇L��)�^�ż�Ll�Rx�y�Y4�7o�w+n���Н��S�-����8Y�8��\6x��p:u��ƙGg˯�5����	��"2��+*�45�.f�����tI�ެ���_��I3w: M\0L��V���ſ�ܽ�zwft��d���I��n������L�7F���̹Qq�YVb�&s����o2�VM�E@<�S;g��:H��n�[{u�Ŵ�yi�A�ou@�����J��G��'�BK`��mJ�F:'�����\?^�������9>�P�G
�;�ad�y�����'�b}g��A
��J��U9����J��\�ݗ>�{s�X#���ǪGE|�-��W>�<o�Ćh�B�sR2�����=�b�H��sl��b� ہx�������҅5�s�������YTN�^n��LϷ|��*!��c�o��~��,SKH���>��X����>�=u�޷�;��<�z�w�W�{��_�D:C�Ê�]R:7{U�x枑������!v��ϒ��0m��jE8��s�C�{l_�p�H���,l�P�|ʰ6�!�m(���%�)M�I��=�~�:�ܦ"��wP��}#��GJ��oD�2j�ǽ�Q�M���6�����k}�Q���Q	��P2�%1�r��Z����D�
EV��%-�{�!�Ml� N�l���Bc�z}�;� O���{�$|܆"�U1AxNC���0�l��|:!��c��S���Nnj�'t7g|Q�q\��N;�����*����I��������7�G��Ȱ��ssB_�IɈ�(u�3T��[1��^��k%p�{#v�:�媞1Z���Q�unK�� �N�]Y�>��}��Ow'�6;���%^A9QB��֜P��z+UG�p��D]�i��/��-�1�PE��A�����
���;�m�8�t=Y#׭��7���F���O@���E���{�̮�Xm�d^���[,C�~�k�Nm䵰���.���kut��;���2��퍛�(J�G����Eq�s�ڭ����%ǐ���MGz&�=�WBN����r=����B)w�f|��M��xf*�A���9��EHlX�_�B�Oyֹ�"E��U{�o�n�\r�nX����2�:p_�ӱ�'��w�Y�����	-����LqM@��kh�J|�vW����ñW����Fj/�f�Xm[�`��s,�h;��1�i�r���h:<!Dk����ܡމ
��&��H���q^�������ڗ&2$����]t�����Y[��#=�2c�X*;>렡X[��m�"�:�<�����X�\�xE������t��I�h�&~� ���bQ�S�v:���y��W�^�NԝJ��E5۹��Y�w$�[������E�s�p�'�*�O�!�ǰm�Ƽv�!�����V��a�>�b�v��r���*�k}��ػ���Z4�k��ȫ�p�>���/k@�s�F|#�^��3�>��w/�*Ӓ9��7t9�z�:?g0<����>�7��{��[_��Kc�5H�$�ٜ;
*N6�@����Qw��k�ބG�떙�&?D$�ql�n�x�C��1�)�PT A:A���5&4���9��4�/�*��M]�s��>]7	�N� �Q�S��_r�迗eD$lA����
Aq�7���-M��Q��a��*�G��W����ަ�gЧ�@�Y�����M�arؿ�����^�����	�^�_z�ߑ�\��~	X��^��Z�Ć(5�r��8���=G˓��T׶}�9~��G	訶=**�r=F���[�:������L{s*������bZ�=u��ņ9�$��||�1Zj��z*).(]z��UH��@��T��Oq�7�W ��k����|�9��;�^���k��mc6<o�Bɟ2'��C����1��Y]B�-�~��װ1No�hK���!��ulফ�/�vMh�}BMQ���IsZ���T$u�׫kp5i�P���w��}:e�E�SP�ςn�}M[�τ���/�Ae7�(W��L����ݷ����_�4�G�*\w���\w�i�ρSL��B�_ͻq���94�#��g$����'���d�}|3Z+ϑʞ�W���y�,�fVi�ƑVaaY�q`A�3��c+2��4M�!�(v�tM�lE2�UM^�-ƅ0�IVѝrK�,b�5A�M��Zz��@\a<;�x{L�N�c�q��pǚf�KŦ���O���u��ꈸ�̉��̣���l�d�!}�n�>*m��ŷ!�u3[�'�Vޮ���*�;P[��6���	�0~�������m�tZ8��f��ܑ�����:��ϣd��D���3C�M@�.�z�O�*�碤��l���+����4��=[���kM�Fy�FW��6	�q�ω��Sd��Ӱ`1�,�{�Ny���_VC0�g�����{���شR�U+�foSeF|�R�x��C���_�g	��ف��[��<�>��՛5��0��4$�+���q���<sN\)�{�.��r��B��~�~���9��N�]��;{�3��?h;X�
='cQ޹�z��`��l�����ޯߍL���z���Φ���B���0gD��EG�����:�ȗO�{��F����o�aZ�C�~�1�b:�)RB�m��+�$��&'FOE�Ke��GaGGq��wUUٕ[�R�>�s��^���)��Cc���Dٕ�Ox)���n�����*�\�zv��µ��t�:��ˊ(���^���<X��#1��$4ܹ� �S.���aL]�J}4�yFf�����rsN���w����15Z �yka��J�s��j�[��NP5l�\�j�dʚ��&����w�;wKCw�c\��ZIN89�^���U�Ty�`���8�ߩ���z�k���25���%��(���>[V`z7��סT�[A5�Ƚ�a��[,3?H��y�]lѕ{Z�z�V&C�C�ǲ|��y#�늤+��5`O�WË/��k>V��7FBY�=�j�wz|{)���]V]^A��~r�TKcr8{q���b$��gýǵs'Jm��ڮRWg���_�ޑAIlf�?�!>T8�^�Ln�<��|�����Kȿ'�q�A�]gs���+G�0Ǥ��'8�lha^ �O��ӫ!t�{Y���.�������_����;X�o��bTx�Q�S���3�{=����'�d
nt'ܻ����Wy=^�R5O��{�����K�_q�y�y�ڬ�aOz��;{�Xw�=k+�ӭ�U��[��7V'�4B�y�,vO�7���m.��V�y�y�~$Pc��}�� b���=6j�1iLh��Kxr������8�&è$[�I�F��bp`*
�n�oV�r��;"Aݕ2�{���>G;�&�2���g|rR���O�nj����Iw`O ���Jy�Q���_�$=:�xˋ���T���s��<ϺW!r�N�yhs��˼�n�/]7~[�u�����>DϮ�6˳�]��������2�zv2�Oo�7�NW����KxՅ�9e;����E7w�w6<p4%{9ݹ����_?&��֠��p�;��R[�'��zl���O�y�ܞ'fk��5�H9m��zIGv5�+�{�EJ�B��X��\�lbCR����v�B�6���x^���/H�+0��ńG�훕=�&u�ޯ���pӻ�K��O��^�s�D�.�b��P��fŭ��j��ɷ-<���dnMJ��l(�m8w�8�g��ֿM'�殾TX2�؝�#E�׭�	"�	�y� 3��>!�7tMh)���_gM^^Y3�/����9�k�W�f)���|��r\�օQ��\Ɋ�B���U\y��#w��� y�CHކ>��~�L`Y�#����?S���TCA��Z�G(��˻�L��$=9�����ױ&]gv����AÑ� ��z�.<|���'��j}3b��;���J��;	K=����}�
�wf�e+��ԝZ�ID���8 ���|���᱄��=���<"�/��_��W,bFV����D�=��[ԈJً�����Պ�c:ƨ��p�O�������vwHv×r���@D�������Ở�t���7��x#�����pJ�O
^��w�X�mkE����Z=>��wTn���i��c�o����I{t��܆��6{������\<��a����y���3���M�G�3NΞ���ӤCFV|��(Ff��6E%h�jt�;l	RV܄2b�	�0�0+��bb�Rb�u��.Ì�������Qlԑe^!�C�{���Č:��;��!�-6�<2-7�Dh�L�G��/f]T3;3�2�Ix�K���܉�T��ůM�y{l���ݰ�q�?]��}�W�#��3������\-�y�E�~Dj��Lq�l�Dv>s�k���.�R���+Ҹ��5�~ӎ�GO�`$��wib�1J�.- �ǽ�����`,�S�u��\|�w�7w6f�дػ������a�3��w�!j�2���]t�RtwT��+s1|�By1WvVD˺ݪ]�oe���j�o6�7$��^���L��b�8�)��\��%sJ���ߩ=u�����:��R���a>ة�C:�W_�ޔ�R۲��[Ho%�MmF-���I~�R��+3��O�{��UoZV$ĽC���=�s�;Ę=oiޛN�4hVFicŧ�����+1Ce(� KwD;t7D9�R�*������=�'����� ���2 -G_���n|y=۫��\X�v�[������?�����n�u���$w��n����aM��getvYhY�PX֭ͦ�ki:��N�J����l�N�y�ė�`R۲�,��i�e`nݕ��!(%���k[]���ά�8�9�Z]"���k,d�'mX6��m�x�,���d�mg6�䲽�G��Z���B陵�gvg���7l�.,賸����vw6�������aYgr۳�2�΋���Y��k"��ې�v]sn㍵[n��:��fUfR�+:��VV]��)�]Y�Cn�GY�ZN0�˶l9+.ˌ���B���4��,�פi�Z�N;��f�N���0Κ�ۨ�ٖ�3sH�g��Gy���+1�u�n*�Ў%>�  �A1 }/=��'r<�M�YF���D�T�vX����񨧐��H�/�m��qm:�>����6�Yj�~Ty�٤O{�7-������ؿ
�%c�X�=�hP~cz~#�W�O���s��yu/�ʪ��E�rʽؐ�RSԵ���/)�ؼg��9	7C[>��Z΅�H�g;�
H,�N𾡫
��a�wf��{Y!����Y�y���^�p�#��ܐ��lP#+��t�CI�6�U\%�$�cN���#����g�n�
���\�>>��8�fqP�k��v�VS�dЇ��d�x��ڹ��kos�;Ҩ�k_tu�f:��Ƕn�Խ�~�*ˠ6���F	R2z�//{�ͳBY��Ai���J���x�;�-ng�ʲ�#'��C��brv*�D��`IR��C��,.c��|�z3�i���Y��"G?Y[x������I�:����=�m�e��i���;s���/õ�G�/�[�Oә¥_j����u�@����ǃ�"��;J��v�엠���h�9clV�ɽ��[:�T��.�B�D*�3{�GnJ�;z+)\�+�����n�}�Q�%�GyF�{ȟL�
�J����7�b�3\@�q�ԡ����^	Bm%���gGFE�k��Z
��Z�}{I<[O8ҧ�:=7.��O_2�R��I��6�z�0����-�+^f���@vZ��*�RwX�y�8�,|9�w����0�Ǖ��z��'ubKW��5���zw.�v�Y�Y)e{���o��g�&*��C뉅�O!f/VFέNόK��^�dߏ�)^|��|�WV�PY�h}�ʥ��8sQ�|c���ҡuY��ʘ��~yA��)k�׻���]A{�b:yE�D����x�ǽ���6iy`���q��k�B�@�H/Wܘ��kA���M�v�^C��Dj1���C�}4��uf��;��nl$�l1;7a�����Г��;�U�7��㱕q��X�R����6��w|���1]$��w;���sx�~>�qp��N��+���?`���Jg��ӻ=]����5#�ԋ�Z�ug�s�s����E���hw;S��E�)98���٧��X�e��n5F��Ӯ�H����D˭��4�ڞ�;S	mP��9�ܹs���WQ��:d��p���St���8��y�U:�B��,�����Ah:�f��{c �ʪT)a-iv�zr����k��^��۬�.���9��N��a�'�[��8{2���i��N���0�[T��]���z������x=��܏x�<��o���'A����S^�#=�XN�Svt��Z�2U�\yj�^�Oq8���횎���DL��w�	�.�2�ϣ�+Nլ;�*�W�R<�[_S>�����E�@���W�\}ބ���g��m���cTq��j7����f�n�GV>/��3�M/�����吱��dgn�}yV
��{Wwv����],5o�{�����sK���<�+�w�рz�K4����X3�ߙkt>u���ٽ���k�mJ����d��h���ݸ�c�p#���L���v�)^��o�?@nC�ځ��I6��S�f���'Ԍ����<�t��G����{�˹�7ԥ5bƼ�\sZ��� �37��x1&�Sc)��ÐA���h ���9|�;MfUb���QW��ZH���J�+'�kb��F�96�]mi��s]#�I���M�c�֦Y��̄P�����Nw���mڄ����ԋ{�6�t,i ���kD{۱*�?tt�=��\G�G��}�g�{�6�u�vexi_z�f��p�K��7E��z`�� x5b�Ǉֹ���~���Δ�#+�h�9(r�	�H���XcC
dhΚ���>]�x��O��.bY�➍ -ǽ	9��[���]o��
����S
�L�~߷�����?x_���PՓͅ�y�_7�7���c���v�{����0G��
U.��'=�u{��s��?_y��o}�����fQTm%۹]��SGP�!�#��*���<�ϛ�u�����5��4M��[�Y6���������겫��?H].P��%�ᾎ�<�f*G]�Ǵ�<��0?6=����������C��{lf��@��^[�2}�~כ՟�xp�Ώ��[��OU�|���P���h�1�ѓϮ�YcX˼���1�y�͉�8�H���+���!)�o���;z��Z�'��}��.)�l�tk�p{�fwY��ky�;�����͗��;�J��"�{��.8׎���=��986T-�@$Z�����Uͼ�Ǘq.�NPr��\�q��IZ�qom�s݈������[����z���٠ƍ����4�I2�����
H;TXj�U5`*���7v1>5��n�>��/ 	��e���`*���&��D^I�w�|Z�c����ʿ=뿷�;ƂN�y�����5&�[ד���r����{j���� o@mf���m���]���P2� xt�C(��\�|3���J�.��(,oH#�W�?@Ǟ"���ꗑ~/�m+���4+����;X!J�#����M��w4Ҿ�ݒ��w�ۋt\4ɂ��'n=��!����k�\+��s8�˝�7�k�	܋PGF������Y��?{؁����b�H���a�F�廩��n�>�MDt;���1�W���v��lc
���$6��9���V��6=��i�<����O�i���b}7_{[{��n� >#�g���Y���3A��f���4uY|�d��]�͡��'R�����:��< ɞ�שÚ'���JJ�w.�����Fż4�0of����y�&�W�N��̹���ܜ=Y���5ڭu�-�
X���ޙm��N�	��N�IN^�@���l�AC��6���W�OWz�s������C$��庽�l����e�����yN���w��{&���!���R,�7i���P��x�C�M�ϼ8�렾\�w-{w� d"+�'��'�p�z�l@k�2��{��Sz�q����bw9V�6�~�U���� �r�l��T��7�p��?HC$�_�h*�.��f��xմ�%�.�٭�3/;bk/o�wN�m]��6D!= �{[V9��vҸ�}[�;ʋ�*�Bm^������yP|�W�Qcp����ڮ��э��2�}u���5V�;���Ɩn��Kv�<�Y �� �9}���~p�K�+kkNp>xwV�l���{��ϭ�	e��|��2��:MH��iǟ��Wlz�l�E'@m��[E��'��a>���;�%�n<�{]T�2�߂֤t~�nj�k�Íͺ&ks!�\:��v�A��ɛ7�ȭ�:�cK;�d�rap��ʏ)�БH�)U�wcՒ����S{�a7�/�yx]��}�44�����]�)�e޳k+%�'�ZF�(h��t�I�q��F̜�r�l����k0�[�G�ށ4�ɧ�Au{�7��p�ԅ��^�UT��b�0�Unڟp����؏H�����,����՚�w�{�	6-���9w���J����( ��6_� ��2�{��c���nH��Y��tL���p�6}�`+�Մ���DM�4VmA��!��2�d�u�}>�����z�3Z��s��1��
���k�^�t2���$Gw�<3�ϋo`V���n�|w��?XI�mJ�]����f�H�&���,���^���3��	o����7�q�ia;�M�ɺv%�ED���%#��KV��uu�xz� ���2�P�i���A�kx�5�Ғ�DЙQ� ��/781g�g/!?��.ݤDe�CQB �6��:�Bu�BZ��tg��WYt�^$:'��X�8�;��G�v�a1�>(=����}�i����.r���Zab�
1�G�aC����S�8��1�� �e��7�V]���RB0�2*�5� ��f)A��fI�y)�Ws��nF
�U%e�+3FĂBK��I4(^j7+�vco�&Tj���,*˝�δ+`1�m�/-s��{�w��܎� ���{NWGz��}����lЯ]�|��3�/�v����|�`?:��z����9�@=��HQ��=ۏu�3w»���	m}�Z��ڰ�z��כ�J���Zێ���ǋX��|��4�0)}_G��7$kU�;���+v��������^��:t8��`��M��l{#�C��>��XjrV���R��g,G5,ح�q�PI��z��=����-�X�?t���G�R2i�\ز�L]�);wٛ>���5���%ޚJ�w��d-��^1�3��%ݞ�~�ff{�Y:sp���d�A!�bn/�\aq�3��O>Y>�5�Թ�VW��.��-��KEU�����aw�y�C����M��!M��hp���A�����w���]�w���{�~��	c���e�fU݈W޹�;����LiGno(�3c6�ަFP���3�g�+��
�qD���"�}����^�W�aw6����Yd�qo#Yn�K�b	�n3��[��3|��;����;�%*n�!���
kSJ����땮p(.m-�eƛ�Wx���h��M'r�˞���g��Ae���qT�ny��>��Ǆ�}�  l�(��kW��t׳���U�B���\��"[�+��{<*خ�cK�v���[՟C��7n�%q�~�.�ޠ���n�̙���������v�m�v����}�i)��y�M�7H<�]�(3�B~�w��qDÅ���������3}M����,������;5�Ŗ-O���|x=����F�����IX
����7x�-����Em�ю�q�s����2�v�׽���s�O.W�\��Yj�����;��]�'rsv%ή�=���M��+ގ�@u�;�o\�	����*vX#]�s���8���Lj�|��7��5c�X� w���P��$n+�3=oqJ����Q4���Jj������޶�ȵ{xЯP	OR��,�LpP���O!��`���N]�����Y�<�@��{�z9P�:�|tv�#zby���5\ ����fth
��qsw��H:c&l�V�F_gbuff�m�4@��:�-C9	�կ�{uQ�A���Uv�z�m�қ�3le�d�Z1Sa�!Ո�)!������������]��9R�W)3�ի
�U�,M��j&�����G(h^��X�mf��;2�+�!A����.�X��^�H���4�Sd#�m�>�0���:�,xfi�>k�/z)p�vc*��2l�U��Mw8c7:�l��0%?`n}>�������^�7C���.�/���+�^�Z�������)mA��
��z��}j�3=Q1����rс�"��0���n�v%�]��ޡ�eWאC.fP�7�S5���z�sm��>�!C������-rI�ӭ������b�����8��{ܐ�ݿBA�ń��K����[��P[k�5������l��c�):�}���>����a�Gdq��,f�RzV�u�K"�l��u����ޙ_j����d@�����msKrV��k~�A{�c#&",Ϻ'���7zV�eџ���q$_��ݩ���X�ᑇ]A�A��a��a����w�تW�������TL�{�+�ا���㙗���8�r\j(���9v)ƶȼӖS�Yױ��Nl=��2~�7��-��v$�"��1�7�C.��۸�r��9y�`H(�Zf�Hʨ�h�"��!L)�Q���
s��^"3�R�V�N�:�q�W)A������<��C��L��r�r�J�"\�[�X9af6�રp�W�<�1 �[����ļ���2���:e8'
�&�3��%����."���F�V�e�,�E��Cu�W�X5Q����`ŸϮk(�*�kͤ�\7�8w���@�ia�����X��@� \��)� dkiCSv\�Ƶ� ��8$Ȝ����d��D��0s�4Of�&k�u[19�j�M�Q�J���&���l)�HF�3��6����A�|�k2%����]�%O����ˁv���G�����[-�g�z�kЊ�����O�2n�^O�e��S]�
{wn��䚱�G|��R��({u�o��`9��8ԝ��q�5fE�c�GǸ ǘ��w1�&��Qg&'�U�)��Խ3ݗ���0�c$����1OҴ�ՉF)�����!eT�#!�j.�1kF7u��VL���3d��k
;�O��ّ� �=a1�[j�ڽ�# d�Ĝ�Y��%�E$��=�U��ف�3��>��i:����%��b2�WU	H���ƈ�0�7Hq7a�E�H7D�U�F8ǋ%��a��O *KO�y��1��P6���s��(��Y�2��#�A���Ssw�w�L(g��+u�J���%]����u	<� �I��yr�D�N�5��׋G��}�%	4��������}W�N�N���=����	��1l8�gc)J���]ˉ��}�����j��n�6����:�hڕf2���S��<;����v#�b.�\�,���1�~�<���n������I� ��cd��ї9����,Ln�}	_}���{�h��Io�O�QO^}����ޞ����b��alIb�p҆�����cm=`9z�-܊rV�5YQfM�<�/���ؚ)��݋w|�r�[��ң��-
����������֑-�{���1:�syhktd�v�>��k��,��w����$:�cb��OPv q���6���K5ak'�ţ���}��{��\��{�U�갫5-�7ۄ�!X���Ǆ�P:���n�vMae- LD	��f⾸7]��o^U�;L�3�w@�wuL��L7O�z-f�����=��o�N�ǆ{{	soj]�I�cY8��U�Ѽ�4&����^�Y��t\d�˲h�z�dрu��;`eE�0���5n�Ê�+V�M�����e:���R����5+/��{Є9s���&�]�h^�V�Uy�N7.-��ݷ���o�����|���~5�2;��Ye�Ee�+9+����9�n�-����ovv����-��w%�o1�8&S��6��2�e�`f��
��2�JJ��l�]�m-3vv��i�+�΋,��e�8;�N,0����ݪ�/kO6ڋ,�mm���q�e��ٗDu�vY�$���ui[4F\X'Y�i$u�6��٪;���u��Y\u�n�.α.ʶn�,�ȸ�Ӓ�,��[wM�6��XvVG�tX�Ӂ����;2�#���gv�م�Ega���֔I�n�8��$�΋�ח�h��[[l��H��Sn4vƶӣ;�kei��L�K;t��ΊD��k�k�=�=�ۣ�'�Y�����tDD]�hOĐD3I�{(�z��=�5��ޫ˨,�.�ዡ�i�]bO�v�UDI�q簍�D�זz���>���z�S�,5.*����I)����A�3��?-��:D��{�&�j�u��Zmw��-�q��z�on��^n��Kuc�Ր;`S���h�_i�پY�$���v6�/|��>����*����7��྅3��fp����F.\X�9�B8�o��s؞Xu�a�}o>�ּH�y.�>t4ى��q"F�	_�5�X6����mw����otq�o��0�r�n����o�
m��Q�ķS��*�/��p���U)���7��v��sх�lG.��n���_l���0��YR����R\M)��.��M_����oyKA��������yn�l�ڂ0t��������x��f�?gr
�������c����aZ����n:V]mE;¯,���f�ٟM�\}��+ɯ�ӵ�����um1o)�yvd�7�,ߟ�=��ܟve�A'Øq3�ӻ)@C��]zo����8���=�E�j�G�z�w��w/r�e�q��s�Q�H�V�CpwXb�r�>�/w���ع�BOr��{����ɏ^c؟���8^�饘I�-�����[7{T(ܓ�nw#U�:5�����C�/�;M���|=�,'c�7&鵚$xϋ��)f��vi�/���½�&��"*Pʉi��ž��E��o�U�$�җ�{}���j�n�Ρe֢�2Alj�0����k��Ԥ<���7�:���*\�i�^����*��Cd �J���z�y&�iհ��|���~�M�����u=Gk��twد���א��pKl�Q�g��;��9��f���g>4������r���ʝ]ף�����jg{��3�@���t���c�Z�+�{���uW|��j5�{S�=QU��V�n{�Gz�S����?1��!�3������O/(+ng0LWvI�����~��o>oa<�c��5�t{��\G����.wkuY�M4N���O�����6��9OE?u�r:`��#��4���G��q��z| p쬵�*���vD-9�E��&\�aA�[og.s2v*ɤ͕�:�4>Z�z�l�pZ��Ǒ�;��@*;��;Ob(�p�qZ�04<�v���% f�3��".�$E�*��rj��P�T���Y7:ڄ��ơA��$�73���~^�sa�B�	�iZ-P鲨z`�����Ƭ]��ד׃��������o��o$)�B�tP�o�|l�������q���7Ue�鄂�М��s��U�� �W�a_��:�}���V[��eX�Ek/�n7l��W�M@�;����7W�J�|_��a���� $�EU׹Eo>����+�ٕ�U�_Z�`)截B�۞h��}�T3�>b1�iy<pl���]�{;o��~��U�y�t�(e��9I�̏
��������9���M��-������>�C�����PW^��va�"p]�J�>2����8������꿠��pu�'�i7ˣע��E��X]w}��=�b�P�(v���w�;�y��n|��,_=GF�q51�qk�}�[���fQ�z`a��B�T���+���wc�@,����] 5��*?u�9�����^>��S[#�{�}���$aS��5pI2#,VXx�1���ϷN��׮�'Y�pk&��wU�[H�)��H��st��j�������n�0����ɕ�p�tL��&�۩_{����:%�٢�Xq�r6�ܦ��f���m�u��L�ޏO��`-�ϕ����yL��{��*�N��o���f�0�)_����^�)��yck��@ !�07�����-ߦ��,��=����ul�L/D��ww[�M*j�*���
oo��FM������z���C�b�w�|�����W� ЯRS�^=X!H
c�Ǡ��9wӻ�{<=^�)��4��m���6{���gFwG}up�k� _��P�z&Ύ8�ݽ�Jb��uP{$T�Ńk5���t��b���
�����{�V���3�A/�;)<؋5��{H�Lz�G�u�X��3N�Lyb^�TJ嗵>Ү,&;��Z
�r�>M�p!�w��s�;�G�A�w����܌��^&P|s{�/'�����+o���}�ePڂy��9c���&}b��{K�G����7b}=ZXy��C�`K�o��{}�VA��w�c����8�K+�;!���Z�8Oo�=���zeÛ��8@����E��~��S6�q�մ	�y������Gv�(�GV�����G� ��vTe#V{yg,s��0�������ï{�;�t�_�˥��i�����kưC���[UU��qP.ֲVomy�8�¾����>`q���{�����D
����q37�
d�n���A�C^���(<����T7���m�ʱ���vE�|y,+�;V�/{�ad��_h��$�X�A/Aj���I�貇�;�_��ZƯv7{�GI��O��0Ǭ�mmsV�Rْ�h�'�;�7��Ym�V�U�7�����?S^�!ll�Θd�ި�:��m�B�Ss^{ʹ5o,�.8����#�.͈�K!q�����G����+���QuIFyvǪ�8����_R�)^w�.}m�t�V`ަRd�-3T�Nf;��u9�v|����νC}[]�ׯ���}m��{^�ܚ�Ug{4���	���X��C$0��NMo�}�W��s�}�g�tv�^�{qK��2����Z�K��-P��t�	X���/��uf�n��ų'��Iɛg��\��Fz��n!��}i�؞p����?Q��x��{�a�W��zp�0lc(b��0���}��4�d�8���CƼsr2�����}$��C�A٢WD�1�`��qOӫ.5����yZ+�����!)Zk@0��ߢ;ˣa����<6z�0�4�Ec{�֪�'p[�*g�J��-����G��0�����=���f�ً�Ҥ�ȇ��q��.��E��[�f{5�{�_�\-cm���㬫,e����4cz��A�ڴ�S��⡳@c��y{�f�'��t-�Eu�����\�۞��zZ�-ھ�멣�p���-z�;5
���w|���Tv̉svaBo��+�zz�Hu�{�Q�vh����5}>��y��&y�yǔl�n�2M�%t��zz�_��m�w����2ˠuO��-�����[�u����Ȧ�\����k���|��k������{�h@��+�K׾�z  �����už�㳈��;|�JT��{��;Ki�|�9�U����u�=�����|pJF1��t�w���׃��-Ο�<����y���c���q3~�o�=O-!k ҡ37�-�#h*8.޳o�5�	�ݩ��$�e>O=*��B�b�h18ql
���F�"Q�G�eV���Q�ħz-vQ=ˬX�MT�l�eՙ/e������^�T��{W�v���nɽm�� _�Y�wg��ޑ}��H�~бR���;��w�9q�G�@����mV��ԭXS�w�����e�������"���������vc���z�C��<�Q���}&���Φ3���⍢װ�:yu�b:{��R2V�Ϋ��O��bx.c�=��Q�E�i.�Sxa� ��E�b��h�>ZOdwN!<��S�p�-ދ>�x7�~��o
H'_���Z��eP��NG���7Ϋ�:GWr�B�x{�F����<x|�Y8������
WD��5*���;3w��lw��B��1�§1,W���}^m�����1j��%=<��99v�ےu���hG���z�6N��^�ڽ/��\����+��è���w�m�}�eU�,<�S����5]g1ԗ�6��E���KoS���#{��x�+�J�v��4^^A��C�0x�(�Q|/|g/lܻ�ow'G�R��"�Ͷ)j��,ʣ�:�Y]��N�ɾ�+po���Č�Oxv�Ș~\��h������	�ӼF;�=��=O��/Q���6�B�qN�W��1-�~�S؞[�kS�//p��9�o ���PS��`i�gr��
rY�m8�=�b���>�����RW`�z��{��Ͱ�n�:���������a�������)�ܚ�ԃU��S����[�v�yb�wq��cO���l���Nי��no���`_X�Y��.}��$���=�6�kf�Q�(7�P�閽�1�>�����T.q������w������k�����?�R������_�w.�{a�q�]�L�s\�cs��i卮����� o@MG��f1븛�5M�xJn��ߟ���|���!kԻ������
@�hPz��U�*2�y�2��Rwa_Tgr�d��������М�u|��V!u]�L�������T42��&��m��{9�Õ �W�S3�����J�gPMl'��>�s]�P;*�8���H��E�8�˳�%PS'gq��[���/F��d��.������
�EY2�/{ E�[}Ƴt��K�O�E�P�^VU���� ,T�h�;W�)S��.,~������ۤZ78�G�Ѫ��W5���{�}��:����I E�	�6�ɕǳM>&w��o�v�^_tX�xL�
X:l�(�2�7u��]�ƚ�Yx|7Y���n/ X�c޼>�`+�:��+W8ͷ�.����,�6N�����bm�w\��9g�j��<�����n�x7ފ�t2��ڃ�ۃ��n�Wj��O�u�s��[R>=�ô�UiR�+��=��*�^�����\���G}����l�<CݞC��G�2ՎI�ӵ_,ʘٿ4�j�o��O>�5�Ǽr��r&�<��xnr�����m�hѸ���Q�5�M���:7�H���:���ގ�5��R�v��\�QwѠ�k[�i��'�;����B(FKl R��F��w+f�w�ўIV���u�ڦ0�C��S�U�L�ќU�f�����țjuŎ����,Y�s�Af�[���Z����jɪw�&�\���o!EE=ԀX�N8REȆi����x y�5%mv1r�T�*���jl̆��IH�'�D_	U�(ڝGr��_/�����C���ڌ���.p�WP��J,�xiZ"�IP�87-^9��F�P�������2�
ȣyd��a6h$c�c?Lw!U��S�+��s�m+�w�@,��f��8�.{:֋�Y��g�1�ߧ�k�G�0|�A�G{����㕂߰�N����w�6��{s��ݱ��!H��
45d�<G�A=)�s��z�����F�K����)�E����!��y`7�<>x�w���
���5��+�<���I��M�l1!�|g�-�͞��>aL�1e�g�G��=P��v��Ve>�j��z�۾`�&�?1\�D�[�El�G��2}}��3�1|����_^}w.�i�����+V����W�nV��tL��,t2���vMC��4N8�{����;�w����d5Ғg�w{SK����{Օgj�
'��Ǉf�G���f��9ܪ�ެ��'�;�I%J�r�>̭x]�"B~�����KO�1��"C4p�����^4��g�G�{�vun���38.~��>���� �z�i�vN�Ȭ��HJF^k��;=�~m��Ǹkц�����q:������.�����p�3s0�3�b LS�˪rL�o2�*7T�M�N��O|�Д��d�	�^�Lb�P���4�0n�:�J��&���pB�1R���k��tN��Ș�cW��Y���S)i������
ڎ� �^[��[�zA!�/y�Jݹ�5��|+��34^Qe��C�{{�;��u�{�3_/f�Lgeg�Ym�l�XF��|34y�O'Ȣ��v��۫�Ǹ��5��Gٹh�{5�;T^�K�X5�탽CRǅZ4	7(jTY[@룉����'*,���s���!�MÙ$����X&�����<��%���N�qrΕ`g�M��R����=�{�Y9u�җ�ɵL�Ϛ'�����qzvo9���np�ɷy�������}޼s|]j�ͩ���><|=��|�`k��Y}y|��5��
�s���:7��d��W�{�7��ȅ*��n�df�{[��=��X+����F^i��Q�W0���s2V��6R,M j�A���:��Gon�g�kzo�k=l�N����~C�-�+��z�{<����2�M��{�p=��ш�l�ؗ���'`5^���׆��[����K�-��$ۼ�J�N p�\؈q:���o��m��^p��٩=�\E�G�w� l�{����'����#���R� K5uW�\� ����e�To[�Һ��l&�.���X�E65��{R���J<B�vn��.�������9����^�y���=��7��x4�&�6�jgm�ݫ^�3_A�sU�i�Ő�5�Sz^>$�v��vK������ Q�E*���V����|�cD7���V ���h����9�(¥Uo빴��ʒ�hOBEP�ݺ�L�j%:��Pu���*/ڏ��=�����\�f^�{�`�Sf+D��fe[��c^�61��-��7uI�D�`:��$�ɪr�3^��B�L�VQH��y=cp#�9�D����:�^cR/1�:Jm	 \F���<X�).D��X>�~��I;�,S���q"s-�����2V)	Y��aKW�n�s���yMJS�9P̥�]��tZ7G	,��	���|I���
���I���z�U��#<7�7!�aK)^Nvi֬����s���ǫ0u����q};E�
��$8*ZH��7w�m�5..���Z�~�T�1"|ZZU[:/&x�w����a)����%�]k-�e��Y�f�_h�Su��%��.�ṹ�Xs����Nsڸ.Ui5�5d���CS��)�j�P�n0)tƄ���͘�р��-aO-��x��ޘ����}������3�#p��.U �}�5;x��S�"&���f��:�F���AЦ�+�y�����s)�ݶ�:�Jй�b�v�k��k�3ښ3'�ל�� ��8���M�$8��b�nΜ����,Q#�]���6�ә���ɶ:���:�[����<,,ٳm��$���[n�nqI��R���6�8���X��М]'.̶�nY������Vu���{޻3������k�Z�v^|����_{+r�n(	��E�J�وD�:�mkn����b���"�G	-���v�Cf��ƍe�}���,�m�;m&�6��ܷqo��D�/k'r�$�C��³I���:mzQzS��.tNN6�u�@�/k��G5��}����[��{W�:��vVy�{X�7�N�Kk&5��i�r#��[���0����2$��,o�䞶1À� |�Xt�o�佡}����K�=6v�7M%�U&��Qf�!Med��^O�$��11CMA3��naN=/��_5nv.�	i֛Էu=��|^B��y~�m�vw8e�Q�B�:�Q󄕫Ǹ��aw����g�p�{�>��f����v-���e�I�%��(�p��6�mp��}�d��p%m<�W�Q�[Nj��}6��H��z��C�W/�`���7]�3���cg��Y��ٱ�o�Q���qw�D���L;9m���<���ͪ�}J��_��檆�ȟ
w�zAx�/���S{v=[p6w����)k]#���j�BI{ba�yzW�Lw����5�{���|���X��GAA�+uS~�N�Yݪj�3��<�������a�e{��u�s�h�}!��
�%�F=SN��-�y��[�����?Z�oE|�N�FB�j�鲨S�7[�����U��p�SC'�=v��*��?<7�.���[�
��B�����j�ꕲ=齫� ��[Rj,E�ׅ�#`����3��m�1w�ֱ`�#�頯2��'sH��.��G�#X�A���_z<.�d涩�Fc��S����Bt-�Ni*g1EV�r�����+cB�[�+^lJf�R��ܴf�a��§�Hͽ�Y;�Ȱ3N���o�Ͼ(�ɡ�1�ENcY�_gl������5�B+E�X��o]3y������^ǓP#�����:����5��3Ϳ"C�}{���h����vGg{�������O�%?X��4���8�����/JunNP��6%��_*iyJ�\�ޓ�6��&���ZC��mlW۶�^�4dJ>�_��;���Х��7l��O����,;�-���Գ�E/o.���ر��͖� ��m4��-��iP��P�aZ�k�<45j�%�{�~p�#�?=����R��o�����;���Z��qZ��y�.�׻Ξ�]-��cf��ꦭVWX��#辻�^%�4��IHW�ٱ��G3^�Lk2n`���)~|a�?q���֮%�-�Ԗu���+��0�c�s/wC�C���7�@�m��ღns�����ݝ���>�z�4��~i\��r�Ʒȼ"�B{a�'�+^�Լ4�uV<C5��ĬeV���o*�`��)�dJ)3�w[����'�pPL��f0�+����Y:���.�ۊGf�Ŕ�k�
�ʙ�/�93�5R�����8X�Ŕ�(]�^n�!k��.�x)�@5c�+��d��և���{RX���8lV�:���]akj�>�<j����:�sK�%*�̽���ݢ-Ё��P��9���n��=;��)CBAe����E����e1.�/;�cA�]0¡�x����w�{�L��|y�ݻ��+�\�PI^#M�s�XS,yQ�������YU�i���U��Y�~S���C�h,J�K��/��tّ���s�^����F��˽�)�e^��T��zn�������*�F=�3k�d��{2E����=�:%+�l�ѫS_O�}�<��ۿ��w~c#������X6���`N��DSoa��xǀ���}@qa��-\>��+��]�e���'�$S�La~=�[p����E��n�!	s�oSo	�ML���0Q����z˩Q<Gh�|�I�u��T�>z�}���g-��Oe'1�G�l���z{��׽�r���y��}��
���4�' �K�V��x�M��wo)fV�Sq��Dk�A�����|+(�'��Lr��%���7��Fj���ލ��������w:�e�Z �.~-=������v�4/�O�w���Y����w����Ŭ���o�A��ß����D�r��K����}咟y��� M*���[�p�������p�-�M�� �S�=�������ܚ/<����<�YʃUhס��V{9����T ���N~!�ٝ~T�������ջ走Ewɨ���2tΈ�;�X��w��P}�����_�3�����]P�����n޸=�����wX��#z4tRO�;�{A�Z��r��ֳ_[��^>�B����#�Z-P�t��a���O1ކw;:;io�M_�Ū�Ør���M�ئ×�m��b�����T����F�V�+���u��xvYw�aVm��k�{5��n�~b�5�6V�8%F10��We	��T�����6�K^1�U~rOsG��;q*�����yf�����ٵr�5��"�&d�4 ?u��wè"�~�t�5�����M��Jy,-Z��e���C�ǋ%��B��n�ݗ�o�x|�1�fɣ��/e�Q]�ZF8qzn�eW����9_jlWc
�X߽��8���Z\h�7 ��n7l�m�����}>���S��l�����G��C�5�o/u��7-n���d���Xw X�~���;5��ץ��"L����/�3�ka���n�}>{3]���"Bb��D����*R�7T�m�����A����J��2��NՆ�݊B�����f�
�4Nm��h�F�G�Wòw��z[CV�k�%ϭw����ޅ��~Q�K���3۶+���,.�C���K��́zۛJ�<�u����y@�8����r#�}�T�~�F� ���j�t���Ϊ����[=_�x�ք��6�a��U��s���t>Y�Z�Z���]�;�xVx�<��b�,ӌ!���r}���n�Y1�~��*�;���d<fx�i��uWgBw�^m�j�}��A/�5��O ���9��ѵ�p�WT���>t�_K�|�v�v��uR���on'��B��0��˨�'D���\��\6v/S�،��E)�	��KN�J��0��H�-��V��^0،�Y�(J����!Ι)�����+M�������Au���#�w��>^�e��P$��Q�������N����Y��-���X���a�3�Զ�'�)jX��o�ݞ^%�V,�6�����\)�t�2�Z���ex�2�[�/!���r���̡�EM7cf��n�{>�HShr��E�%/;{�i���T-{�����4G��jM�ZU��|�^m�94����뜽��Y��p���.#N�k��uA���܌����w�ENt7Ӛ��k�O �֦Xdw�ǣ�z��FR쟮h�����)�Ϯf��`����y���g��3��;�M,R�J�v�ޡ�fG�q���r���{���Am�B%h��'q�)���&�$��1��p*b�����+��K�^�����C�Ob�햖qm��K��&Dt\,ֵ�����Ǻ��	~f�A{f�۞K-���K�M���M���8p�x��j���g�L�y���p$�i�O^��3/	�?R�Bl<W�C�/�
�˼6��O�v���N� N-�F��+6Ͱ��<;���L���&� �E�Pv�3��[X��Zr'v�����=?����Щ�3���}�����r��wuo<k0�cuϟG���A����w��x�ݟqԶl�Q����k۫�o���|h��}���9�̟�}�b��U�Rw�A�nv�̝CXz�-��<0���oױ�K>�՟=��`7��D�$��xT\�X�o������ JU��v�|�G�k�	w[ϩ�_5c��|
U��M�z�uә�g����(	a3�gr���N=W������
D\#u~���xou�'��Ӣ a��P5��A����缩
���ZOe��_]goh�K�}�]_k��t�"�S�O�ְwF�q�5|�&k']�8oU���ag�W&�����Κ=C:
g�1MM��&=�	���H���4�.�6�����`���
��m�}�fF��jȿ�W�Ef[���cy�E�8Q�ܩ�����M��p��*�˙g�\�u9'9v�=ɇz��d�{w8bܪK�Β�<=�f�:2k�vu�3P[On��Vdq��Rvq�.�W���w��@��u��^�T��@�ʧ�=�a ��dþ�����p�������o�(g��ʲ�,\��q�d��jz:�� _����[����0���o��_`3Y>�����5�%��{�F�׳�pj����^���|;<�w�W=E�߭eW��m����ޤ�u�Mxz��v���y��X����=B%��'��Tg����^S��s�����+ʺ�\�m��,� ����y,q�y�צ���jD�S�\�B�dyW'��i��iS�mv���۽�;��̓�?k�{~}�[c���U��ּ�4�3�D��ciʺ��y���{۾1��ßL�mgu�ڶ�E��P�,��o�1���^k�ِf�� 'o`U������V7���=��ʍ"�[�v��p�OrN4�9�c+��פֿ,r��h��o�ݩ{e^������?L@iqs�G-�~si��ۯ����^M�����.r��22��� �\���I$!��'D8�{d������oYb툱�m�\���W�Lz�6�ـ�s�;�}��}pE}�n"��=�dR�A�:z�V��Tf��8A������z�	O.���F���t�S�L�y\{sZ���3�M훕_��V���>�iҴ$��Z-Pb�a�����Ǣ���f���gގgb���R�o���M���ß��3�x[��=^���q=�Wpć�?o7T-F��o/Ϙx���#��o&�������"���3�F�3��h��o�!��7m`����NV����J�SN(���D�'�y�V�˞� �J�kc��wlaÚ��j};_o0�ѹP����a���7���j����k��ʲ�X�ù'���<f��;s5��>�{���w�i<��	�w/���+^B���
tU\ٹ���yKe�������_<U�v�K��rv�n��vQz�M��r�(�qY.�sy^����;(mnC}� ���m��ܫs�q���#c��t|P����~d������3W����ϔ������t>V^>���|����Q}.-'|z����P� �J}:*��jSqR�L�)�J̄�Nn��n�cԘ�AlP����(2��à�����s�ԝ9{Y�JA�mש�4��d0�>\:�zU�f��6��#Ԏx���Mn���=m[;[��z�s��a��Pճ�O�Ueu��U��� *-p��c�`�M*�c~{��>�G�9_)�w��czD��[U������-I�W�o}�����,��[]�.����{lz��=��CzA	�.}��ɇ#�71em�uK���ߺ��byylw7�+���]b:G}��t�O��>ץ-�]���ƺB�^[K�u�[���l7�\c�|�'�ip�焜�ad��ꘆ2�����6��H�����9�..�Y��S�<����k!>��&�>q��2�lߚ��>� ho$-�A�p�<�cy�y�n!x���{"���S!�Ts����|��TNZ�m�F�����xu�
�h VR����q��Z��~�|�u�~_o%�K�!��)!��U�]$3����֮v���e��U��,��,VN;��J��.���-쨬�Z�-[s���e���� � 2��A�P2ʪ���-�YaX, � e���,��2��m[lZ�,�e�2��UVY@� 2�Y@� 2�j��-���aY�e�2�Y@� 2�Y�[lV� � e��,�e�2�Y�P2�+-iZ�L���U�RU��,��o��%T��IQ�RX����K���;>^7�ӿ��~��_�W��-^�5}������W�Z���w���s�z]��B�y����_��Z��?��^��NWmzb��k��>�!������C�Փ�������[?�[L��y�y����C,��U��*��J�J�,J�0P��B��U�YIUVJ����)X�J����bU[���5^__���̢̢̤Ϣ�.'�s1���n�s�y����B�v�����V܍���x�ߛ.wZ��{��>WY�^��[
늠�j��xY_{��Ũ!��t�*�&M<>����M�i٦?�_.U�ڷ�������;l�k��?o!���kS����=W��쭺ux�������jC˥�!�mչ�2�g��^4�X�����d�Ŏ�&WN�hB�;5��:<kɴ���gW�OR�����gs�$!g�����O�ɩ�_�b��L��L�b�Ψ� � ���fO� Ď7�_>�UB�(�I"AJ*)
�D 
�*JU*�D)JP�D%"��EJB�R�*	�E@�%R�R�J*�%EkR��J��ʃC[i&ؑ�->���*�d
)l2����r�R��P�6�J��J��J*��	���@͛m���Z�Uզ��%lĪS,QR��5�U%J��Ѧ�4(!PB)
�B$E(�h��h�R�(��JQ�(U���*T��   .�imT�۳�Ce��N�.��]��0�u���&�#�v�wh�ж�r�m��w*�����۶�7wJ�t�s��WM-U�I[��n�7
TJ�����T����  wnOa�"�R�H�/=��TJ�BDQ'{�w��(P��dD���:����2U�(l����V�mR�#���U�R�quv�R�ݻl��m�n�t��Nj�6jܦnuݱ��5�ٕT���WZ�+��ڤo   �m�䪻��hg*튩W.�t�6��r)�i�7u�'q�n˻]kJg�t��]ƥ�M
�]�,��V�*�Z�ҹݴ�[M�N���wj]ή�2TEZhv*B�TT��   {*={mu�mn��m.�kt�.�]��N�mћ]۬�Wmu�lnun��3�\�j���[�]�N�tf�ܳ��s�v�j�Ur�h6��:w*�Dv�I�Z��RIR��   ��h�{]Κ+AwQ�f��GN�¨�ڋVTGE�V�MQ�XV�g9]�5Ar�:��2jtaC���$�����R��UPH�  ��V��κ��[�mÊ��6�f�gI�TN��w4k&��ƗE��5֪�f��A� �U��P�;a QUH�  wx�p0�C9V�mR������f�X��ۭVզ��k�ن�l49����n��]K+� tPRw2;j )B�  �B����c@ �t� ��.  ��  a`: 	�� n�4 ;���C��(�i�Ԫ%I+c$����Sk�  ������ 4 ڷl@ �T��Z�@��t :�wA@��
��5�˸:j�&�T���9J�����h�hҋx  �<4�OTwR� �1ӹ@��r�:
 �S�  ��
 ��w' :P������n��܌ tx)�4JU#@24Ѧ�S�0���@h�0��I�   E?��  ��RT�� ѐ$�T&T  ��ȴ�]�F�`�  ���C��9��T��!�E��ҲW��P��<���������3����m����6m�ݰl���6��lk���=�}��)��
P��٣V��>�p*�M���vݑ(xI�Tr���m��nRҫT5��Uv2�nU�W�aOE���.�g 1�����gJa�fR͙�r�۩i0�C���:�+V�G�m��e%��6��`̖1%��ڍ�;n�M��L��g(*�B�ݧ�k�E1�-^Ҹ�[E*%	B��)PՇZH�f ��:R�i���K\Y�nV�Y�X�Z=wI�|l�����ۡ����
&r����x�5V�Yw	.�\%k�Ђ��XN��>�&4�I��.�be0n��QQl��>��Ja��zʃcH��t�H���'Cj�����1"bo9f\Kf�%�gwM�u�Z>/u�ś������ZdM=u�8�ELS��3�xv/E=؎��{�u��:��C�V(�b�XFi�"q�H�a0v�n�m�^d�j�9�]�m��{���
��2kj*S��#�kwL5e֠��D���j#y�^�$�'n�y�h��`�,�d�mı�J�4A���؛��t�^�lک6�����e� �L���q�"�[�l!y��^��40�Q	�y��"��22[����Ƶ��;W�$�iÖ�Ad�v�ݥ,�E���r��fS-���b&3[1�Q[dZ�vi�!,��W�m�t�b���q�y\e��kK�}y� ��M��1}��VV�HL�*\FKwM��7�M�%�1�w6�L��*ݽ��B���qdn�T��l�	�S�o1�B����x�]4���R��bm�W�Sf�T�V�� ��,��u���L�&�q��جQcu��ܫ�Z������e�WH]���m
�MM`U[O.��@�m��6�Uk��ˬ�5Sh��hӴ2d� �d�r$��E]�J+1a'sN�MDE��X:���*��ʎ3��I-�v��iV���x�%-����;�ɓi�,+��	�ji�m�e�H�]�tHx�Պ�Hb�*��A��@�x˦�7RS83n�,���$;�ma�Tv��Ռ�ǭ=e)�s��B��l��.fӁJ�D��]�O5����]ܘ��1,�iܶ��/^l�.AJn��H3�V
ƭ�ͷD�����Xik��n�_�Ph���X2	��t�BЕ�l�-d*������������U��h?��P�!�lU��&�ȷ3*D�%�l��Q���[(�n�6��R�A6��g���e�r,�H�ċD�;q0�b�F�&=y{�*۠���da�2�Z	e���i]�m�`LvlC���sq�{�\6&n�*TM��]��2�0���<��H�W�4�4˳[+̻�N8�ۼ��[E��KG)e�t�w�.�8�^�5-坨�pổ��>gV\6�+mn_Ҕ����&�^йyE���Kj,��r^�)��u���Oa׳Y�s2'��7[��`*<۬���h�Z��1�JѪ���PZ�ڬ��IH�z��L6���h��S%�'�d^�x����9�V6�1�#z�Ŕ�w�fHv��J��G�W�i�J���XU���Q�1������fe��N�d����N<	6v�f ���]mml��`��i�a�ÁX��qc�B�uv�[J;4�n�ԦZ0b����[�m
�ڟAB�6�j��Uz�%6��f��U\�P�������rɤ��6�i�J�����az�V�I�h���E�ҕ����әgqAK19NVc�6y��k�Mm��XXp�ݬ�4�V���p���Qj��ƷQ�&)nRxYv-�n+ׂ�6��'<���*���%	�RZnݴ໱��^�PDg��2��E�gN�݃�!�Q�r���9�2��j��&�0c�#S��Z	�7o�z�M[J�m��n��M�O",�5�Z%@ӧ������f�N��&lƣT"?6��2���=�ҏ��M#.h��`���>n�i�MR{�Py˻*�obF0�7]l�q�8S���
IcY�dx��yd]e����a�E��t��{5�b��'� ��9�P�Ѵ}�����vѠ�;�-V%)�!N��rb(���ks�2�R��zpKI��f�l�6�"�!kl�Ӊ)���-�EUf��������6�c�N�%�6�]Y%�V��Vb�Me�M��SN� �t*&)*�j�{�ѧM�Gm�ɡ���*n�AS@����eYox#&
���Ջ2d�I����+.ȵQ�:�+W��9���A�F�H�F�Ux��2J��A�z�*�Ym
ґp�A����ZY�PƋ�z*�jB�k^
N�iPx"��H֫�7j�c�Akd���߭�z-M��7d6�oi�X�8��tˑ6��^�aSoe��R�$�Sk0���
ώR{h^��ӕ��Qf]ʷm���CR�Y�ӐѨ���N�e���P�rE�7��R3`�S�u���c(E*j	U�E���&ݸl�v�� �T.���Z��h6��l72��h��-a��Ӧ�U�
2��_֨9P̌���0^۷7%1<��Y4Xƚ�X��ѣ7*'��Z�)�a�Of�Q��kn�lJ	�j^�y�D32c�jf��2��'U�]�ux]�cDU1Ki8�D5�wid6`z�����̴с-J�䁍� �(�a�O)+sM*++�a�]���a-ٻ���:��
�!�i��4<waڕiV�Owm�5<��m����w��@eјw����r]��nP����x�֖l�w'�@�2���a�h� ��]��X�m���X��R�������zؘ�i�q�����7l銡��Hj���y�#e��`b$kW)#2��H�+x�m���?�:�	�)W�(��
���i�fQ�-�KJ�P�s#�I�ɪ����R��U��ޖb�p�{+" ^[ʔ+��R���'�7I�rHh���	�kT)�u����B��E�'bX��wx��e3�4>�V���T	Ù��lgV6���ʴRIf������-�ŗKM쿣���=ͬ�AS
`KXV��[q� V��ܦ�v��7r��e04=��1���V�]'����Qqˌ��u���4Yg�p��+�.wd�MdXU��&$���nM�L�޵�*1\X-��1�.�څXf6Q.m����W���ȾX��2�w5,S�w�GQ�sYyx$r�ז�E y�h�J��晴�q�D[0�R���q�r��^
�[�e�aJ�x���U@l�p�C5m�-:LM�c-�ŤG���Rq��;-��A	Pd�n���ʂ�?���(�6YI��6�9J�.�,-�-�-AB�T�n��"{s^��gJ���5h�����
fꆒ��j�;K2�V��F=`���GGٻ�wN���ۘE�L\���m,se���X��a:I3t�v%���,�z�ѰɭST��Yx�P��Z&#��V�&�;��d��B���%(�B�+[`e�4H���o1쵫LZ.R�1�t�y�4��K)Z��+C˳L�2���j��hSCqU�����M�ȴ)�d��l�Ve�3
E�]��{V�`�������-�8�חm6���J�� 4���ё6l����Z��`�(K*�Pa�s6TG�+7TM
�խ*K��trm�:�ъR)d��QHF�[3	j*"�{��ϓa3*��C�ױG6��{�mU�q�XM'�Kg4�QQn�LkN<5t(@����Q��������V�J"�՚kl�hbt+B��#�۽#o	�s0��M��5<�gF���@.	�1EI���Y/Y-ޭ)]��F+�t���M�Z�^	)����5,��hŻwj5.M�qZ{%Z7kuB޼n�B��
C�kN��L��q浻��V<�Ӷј�2/S#"w���N�o�X�ysI� Vd�ͅ��]蕯��=k�t�մ2���e�v����n�%+V؈�[��M��ie��uP�[HlH����+ �4�П����17���Su�K�q&�c��kp[�&���g\����Shk�KOCE8C�ByP���j���cd�� �m;�3BN�9���|��킞ͣN`!�+k�A`�Y��7d8�'��ʼ����f�^k¤ˇv觪���2fZzu�6��|��[S*$�9�K5�}H�[���ޝ�����*�)�
�՚�W�pJ�V�c1�I�Dm�π����n��3*�gtQc���5H���:2��3pҰ�n����)V:P](n��X`�[�z��w�CXś�4dI���X��g���w�cx��S��I]�%E5Zܦ�Q�٣*�Fʦf��L�е]5HSy��;� ��Yy�;ݸۀ��� b�=X����� �5<�p+Ꜫ�g�eTU1�9T�:��M��F1�G.&&.�3b����ѹ��lIz��6:�kIU+**�wL�����L�O�6�+�:��b�ҭ[N���m���L\X��h�X�ݽ�%L��G%��L1�{Y�> �ͦuYV��D\�(u���g��e�Tl�kݴ��Zw̺��Cfrӛ��E���m��e��]"�7[S���TKN�c��N��k�YTZP)��kEɔIܬ()� D���%�FDJܢ�Q[�Z�@�kYt��q�&!��Қ��a�b��󆷀�E����3
h����[om;h�`�k��.�Vs��k^pV��6n�hf;$�+Rj\��0���f]���7JR�]�0e:3$L)d�{x�^���9��yC
��t���5sfRMïbm�m���dT5t&������*�*r�a�;AVA�6ٔv��b���$̇n���$�
I��*v�����ٌ��Ӛ^чq4��w��8�˘:���\�y��uA^���xUa�L�`V�7t��b�:�3l0��V�X��jM��S���ť���EQ�V�L��Nn����[��ܭ��/��3�P�W��jŚ%��6U����h������v��eըvm'1mc�t�+7�j�dɧFE%���h�ܷm�b�-�j#3v�r�ˌ̼D]�KV�.��Z�#�5���M���2ĭz2�5���e�������3/r�w��n��D!�{��y�+��B�D[�\$-�`����o)� �|�(h[��Rm����Y]��)d*웼j�&bIX�u]�a��-X���E�ٔiZ2�cۧ���(��#l]Y(���8t�tMӷ�X����y5�0j�tn�R$�&i̳��i�\ YnM"�F�	�hꝱ�H�vs"�]h�ˬ�J7���liqQ��f%z�)M0Tz�F��-��f2fn���hi�P
��6�Rd5���������Z�ۨ#�l�fR�!PJ�� �L_5����#�Zn��sBL��j�^�F�Ѝ�i][���n�ׁ�9�b֡m��U��5��2��SqS�k3i��"�P
�76�Vd�Z�D�3�@z6�R�p�ƞ�6�l�3��`�m��cP���Z凥k�8��0�����iS*�ۨ�h���
Vl]�%Y�**82�홋^���f�耚yN�[�X̤�Ѥ}��� �R��b�,9Ww�lv����*y�h.U�/V��e��Dq� �6�90�0TY��ƞV�:"��-���'h�(Ѥ��Cf�Tٱ�Ǆ�����>�+L���7�Dı԰n�Ld?�kBy)��e,�n�V\����aYS"��I+��X��"����%q#��3�dӋ��Q��˳M[/��B$݉�w���l�ݰu�4[T���#.�*YLC��Y�*��
9��������f����kh�����^L�N6mn*ܒ��p)���`��o-�!1T͑����J�=�9�+�LK�@�{�6��o�(l �Z�4
�,k��)3V�[@P�*\B��ԫp�8�l��D�F Z�h�b{���]�[��.�0;jZ#)��ݴ����P;��e��ܺ���m��ѣ+��V�B��Z�����F�*6�|��.f�̑�M�X2�<�`�tV]3z��F��[D�1��+�(�e�2�����i줨�J�@7)��nM���,�g�S"��*�ͬ�Vʕ�Jzڔ\Y,��n'�&�z� b�0Q�U3�VQ��2���
[�%��x�D�	�%	J��v�Av+1 ��v�])5��⬁(�Z�E5���{ܖz��y�0EnD�Cm:-��Z�q�3j�� ��V��z6Y/�sTx�A���n	w���e=N+&O�U�Rm)��CE���!�z�2`7(��v���"�5x�$-⥵-��)������+��#�իGf��l$��)�f�,Cj��D
��zغ:��8+��P������mc��KF��Ӫ�9��n�M�����u�l܎�'-#c�e4ت�H��u�yXީ7q�^��%Ge"�T�*0 S!���i�cD�Yj̲ռ5�^+	*ENM�a1KѶt6#hwq@̍���ަ�Q��֘ka�C*M+4���P�{�˺��V�;G_K�?�gFX̖�^f��� 
�e���k1�˭Ke�2��/�jL�z�1��R;��G"��Ա�,h�.� 9�o&��/E#���yK�F�5W�S�)^+[
�v6�CCn�Xfjt���6(n񸔖���cV�.Dh��j{���X˵qdۼ;��&�[ �-���`�[X���!`�#��ݷ`h��1F��լ�e�+*��WQGbY��,�keJP|qգ(�Tz-�G,��s��s/�s��m�H[��z��5�1�4������.�Gic2E��nW����s��5�lvl�w�&cL�ܶHGwd������Wق[�D�_U�A:3�R�5�rF�����/�C���+7r"���P޷�����o���K�9��D})m�S@]h��+d�����&bż�dvs����9ȅ�a�]dY��dA4��z���FR��3l���y����Cta9�b|�����쮴}����u��Iyշ[]�k�ي7�7/N����=hkV�L'��˄�a���KY�N^��iyӐ�yvO��z�J�Aè`�5��!���^Ͱ�-me���X�8Yκ��]���]�Hvd��'
l�N��Z����9��q(�o{"�7wGs���ѱ�c����	�M�E:�B�-���z�-�q�7�p��Or��i�ϻs�S����<�����9W9U�
&��ovR�2�.��r�"Ɛ���uMF%J�-جU !��\v�V�!|��V+����ם� L익ԥ]��fb}�phc؟�Vz�5��AZ4Ҿ�h,����]�F�0\8v���J�v��2�*p�������\c�a͉dXZ1h0�5��R;B&ɧf��]Y6U��z�IAb+/�<�2��6U+��
D���橉{�se�i}��������=�m.�=���6'�l3E�tDw
[E��Oz�bW��iC��[�9p��p)QI���YN��t��"��NQY��:}\
X8m�u��㍺k��(,���Ώ�����3;��0�a�qvT�*��`{ƴ+{/l֟2(�������d$|�����~�ټP�[44`J�85ć�N���Ž�������6�S���fq�;`�KRU7�zv�ZҹR�t������Z�Y�u0�����]�/�Y ���*����j�a6@O$2q��vs h�qᛵԙ�����\��uk��BE앺�`5<��p2o���
�	��eb4�s��{�z��fU�@sR[���bi�'ŝ��V�|�dݸ�W�|��ӹI���wT-�����ɗ�;{�ÝJQ���� X�*"�7S�r��K�i�ܴ��^o�D��9�U%yn��=n�c��/��&m��8kyԬGg�e����r�V������2q��*g&�{n�ۢb]u�F�����q�pƢ\7I�
Dk{Nv���ݝ: ~���Ѵa˽{�c�t�t>�9��%�]:��V-yMX�q�*���Q�\����%n�T�� v@�6��.P�lk��}Ʉm������%��7�Y��v�]�u��5����l��9e�Y$|)�lr{���s6��ݒ]d�I"FC:ֱ�4W �ge{�[@""�K4zIMa�S�n�JQX�0c/���ɹVj��ǮX�ĭ�t�"��t8iٮ�λW��:�:!���E��f�Y#_7�C���f����J��QV��ym�a��V�U��;�� �� ����l������:�I�F��ʽ�[���!�ޕjPN��v�w����l��&�nJ�����r򻀠���H\Ш�8���7�9T��Բ���л���V­u��ʍ��b(�k�1a�Õ����O:�8�"�{F�ǺhU����!���K��O�X�����(!w��07���e��$m]��g8_},l���2m��u5����6EIgu���Y���F���lT�iktX�@����;�`��ԧIeIt9�i��'u'o3U��D�el���#F�V)�n�����74%`V�u u�l(��X{��j��98c6)�N�f���X7�O���Cd�}�`O��mlټq�'X��r�曹�Qbv�s#���H�N��	��|o����1ݻwyī��p]N�#�I����]�q�W���p�q���d�p���˺�Y�pw*��3����BQ���U��e����2Y[M�xU�{@�w;l���rn���\�zBUv	��q��)�|(��@k�S���rL�߰��E���]�W����Y:�f�=�}���Ѱ�8���yf�J��n�F�ٲ�u.���Puu'�K\���nb�,���w�����u�:��ʌ�����9/k���qdFd֊9kJ�.�1:l��"4�4%x��2�l�;��9���2qÈvhW&��g҆5W�Qq�u�0MVjMʋLE(�1�Ǹ��g{k��k��6`�u��Б <�R�mc4@�uٻ��:<��l;��H����$C�L�ԯp#\�wn�
f��y���K�Q�+&��іqRyx������V�Y��9L���:�b5��T��Wk�P,�N��-�%J������l����ɮt�N\��dt@��0�ky�)ۋ6Gr���7o#;ɪ�hn����}V�«����ю�uVt�ɘd����@^�ܘ�Y�2�&�����{l��cEe�6�tjt%e*�T�n���s�w��'�z�y\�K�[^���{x�S���ր��h�_�[ �q9�v��{���tf٠�������\/8;�Xs`ms`miP
1c�:a�sNc��BZN;|8=���eږr
|SfR��&��w>F����{`��æ�;��C��oZ��f�^���̭��}�����u�'r��z�&P��N�M�|�M����9#'lKy�ƥ�iu�O1�ӠD$��i�����hfV�Ҕ�SI\�I�z���ޔ�	�˒��W�g����3�,��	�����t�vEj�4M�j˜��[\������swj
kD}IGՔ7z�f��R{�T���ޓC�H;<��؎l?2�r=#_�l�D�:�LY��8N�e���Q��
Z�J9p��m�UƁi�}�)4p�ب�
�kq�M��j�t���P��p+��o(���I�[+����8oS�َ,�ئpz��Yјv] ���yW�^��)�b��	)e^��ie$b�h�I:���|�i����ˤ��.���1:�V�,�.U��m��H<C2B�jaƉ��v�bvf�9(v�'�	VX��n�[�'�+��c�ɛ��q̠:q�\�'h6�of�9ݶ�mJ��u�����y��・hV�Ů,����b�W�d[G�e�c�P����=�D�3�W����ܷd�@`+T�j=�\��5;��rE�2(lK���:��y^���H����n��ø��Ƶ�/jnWo*�2���a�:�g	��u5���[b<d��|*��vʘ$] :���r^!nl9b\������|f�pl�3}OB�ʴ�,,B�U��Պ�����us�fX�������{�Ko��Z2��̌X���	���ھ��H����݅_n��s��p����E3B�1j��;�d�T�ɝ�[Ϋ��u�޾'����$�zL���8�J�+�A*(T�
���	OT��Z2e���[H�ޙѳ�r�/2u�d
�F��	x'�Kz�YD�N�	M ֫��n��ҷ��^�qf��d��t�{ä���63��ݪ��wYm��޹u�t����tJP��KkZ�P#M��}K�{ϤNnb� �՘�� ��V��դ��]�'K0h֥^s�����x�շƲ�+��;S�e��dB�̨�snc�w�Z-=Y��/lH�d:�q]���Ʒ�Z8�f$�I�O;N1�����§l\'�(e�m���]���y��nh=i��՜x�L�:��Ss;��C]�Ƴ%���¨�i4T�׹�j�RqAvE�2Ç^6�I�v��Օ'U��n�}6�:i���x���!r�4:�1	��-]f�vO�I�̖��z*�Y�Fr���U�% :u;��)�{M'�/� 6�$f�V!�	��.CfVL���mmߵ�|���]A�9ܟ�v��E��pu�L��;}�ҕ��7�
��:��x�<X�u�J���zU�1�T��]Y��`�n�IS��{��nʷ|��J<Բ6p�0$����&��6���w�=���������JA�L�.�1X�Y*�D�Y5�>�/�v�	QQ�W��X3xD���yT�Ye�/z����u��t����َ����
��T�S}/T/��wԖl���"�z�o_}�XOT/yn"�Kmo�WT����[���J��}Q}woۭ�����V�3�	9ar��C�__׊N�t��8�ʻ��;c�˱�ҼwxɮS9Qww�p��u�`���cv����<�ˀop��� x'7tn���������]�6�;�-�ެ�N����=�R`�c�ȂH��'�]}.=@L��fk���ٴ97�na�T�r�\�q̳g��Nqqm�9�� �����tO��z�ڥ�I[w�k���J�8��]\*�n*'3�ڡݐˑ�"�jk���>K>B��J+k]J����Q˓�|1��S��"د�oP�t��i�&w��%̑��-
W��p���eZԺ�����*D��w8s���o!��ɍ�-^�~�;Cn�W$JY���Y\�0�U��6u-`��H���PV��LqGr�9�i�����\;ZhS; zt�6i��:�k6ڼom*Ў^"�f��z�9�f���/��q�u�^��M��'s�qNZ,������+nK։���gb��E����\�Z�B��m�L^T��k���F�T�U'�v��X��gGlu�gVҾ����C���+m|.e"s����JL���-�uB���pl��k8��)ڬ�E��� � �;� "��ؐ�(����$�Lֻ�����m4,�2�(V\˃���D����#}�;�^٧jXb�vV�Xz��2�4���YF�E����+�)���[:\+��}�f��i��h����K�̸^��)=���p�3(�����%*��Xں�5���XuU���A�]9Ɯ�.���2o����i�*���kU�v�]k���.���wiYun�# ��H�L�t�G=c�#]��R�aڇ���Jz���C���zo!��n��3�C-���GC�P%��o���k�R�w噰`����>ⴽ�DՃ ���w�DZ��틽�yA�}8�y+XV��Z�!�]�"�/FPp��xe�Ւ���ќ\շ:���c�Z�Ɗ�4tj���N�֦p!I�α,�=�iePT�v�*)�}5�aAm:t��ّJۼJ 0U^!C��7!tʐe��Wut�:��y/�M�ө�ˏ7��E3����)�}��a�/\����y�8��P\Ű�[����j6�J��|���o�u�R��Ђnf��o��Ĺj��J�	.�v�����ČSx���5n^�u�/����tˇkiy�=A�a�-��&��$=X ��,Ox���x�& {X�*\9W.��HSzF��zfn�v��];���� ٵcV9�E�)�ttd�B�>ћ�Y=W�h�^Ԥ�ؓ}���[�V���׽n�޾[D�ʺ��M�r_Sח�gz�7ˑ���^��|vE�d���:r;k�.N�ݒΛK��6��S�x�I�T)�b���dx[�K�4R���L��A�xJU�����)�,�ޱt벍Eh�ͫĚȫBU�goti��_:z��K�7b�j�z�<.�o:���[BZ�Ō�C�ܦp�T�U�=���%�Z^�c-]���NebCn��8�����Y���y���8�J_��������B(����|�r^��Y�,U���dK�󻥳ܡڌjW:�=�;Ou�+{��=�Z-���U��=�e�g�;4f#ڂ:#[�Y}�)pV��;};�����}�;����lf�A
���;�f+�+k����'�j�ͧ�o��z��/�M�ga%�傮QB�E/U�R��`���Xm�	m�-�;�{:�\zXˮ�I>��ǰR˜ܩK�j�^pp�d�M�p�jr���%�*q�����]n�4`n�ϣ閁��Om�e�u7r)A	o7y,m%��k*n��n�ӄV����*k��UN��)뛊���6T��঳eۚ))�M�e$e��b�5��\�#}�тU��y��H�s��p����$f�r��tmKI3�PT2�}.>����J��{�k�Y ����B���C�W�u��od�H�Ϧл�u�����7�Hu8lږ���e���Wb��l`�F&�q����ŏ��X�]�8���*
����rg=��He���7\��a��u�N�僳'L����y'tۏ��
�V�v�����7;�o�8�I�YdA!�ծ��7�jX�7(���;���T=��9K����1���z���'�5�y�P�\�.]<u�~����%��Go��S�Je�����v�n�2� ˩@M��#��Ȍ�}��rՆ(a�{w�j���H�s�Ff&N0Y���T�k����!mJ9aK���E�ү����&A���pT�ŵ���]aʺ�ʖ��Ogu�����y��L��E�o�IC��5G}N�=����t�n�4�^��KxW-����b�
$�q�[��@�zi���]f6h�2��v ��o�f�i8T}�}c�fc=V��a��Q�p��GjE����:Ε���"4' �|���qb��ܷ�_rĞd8�r����K"Uٵ���a|����6sTs�*��K�b��u�Bt�bKU+����}�r�0�"�K��I%���]��n�7���[@fu�a!�5<���h��&�qn�}]g��6p�к�`Ӹ$K�@�b]�<��\�"�\�ul��5vq�9q��x���8;LH�"s�ֳ,n,]����ߔ��*�D;�p�˼��y�g2"��#'K��L�쳄��苝I0��{���DV%"�(���
��z���{�{����������������L�¯�D��������s. c/��tJ�{i���R��o��uL�ŋ��n�U��x���ֺ�=��@��\ɱ��\[6w�Pws�c$V.&$��tto��x-�eIW�n.=u;4�lbWi�M�@�(�j�]2�<����U�ɤr�5*�A�B̠�C�u@h^k�B�ID�1۴�86�rmAg�wC#)D�T��jWB5	�N3���t�nm����__f�8��&����[�l`zxA�i�����{Bԕ��C��F�I��h�:��y��X�.΃,�Ü�7����cK�h�gx�A1xp�6�5�,S����b�W�j��ٺ�C�'��`��P�KV�rve�^�Z��Yv��e �T��]�<�$˪���E�w�Ϥa3'Y�qT���)�vL��K>7�2[\^�( �cb���z����,fՃ0�H_S����e󷴚
oSa�ѕo-���Ҷ�,kr믯��X�ͷSU 7��������$�ٝq�r�A�ȶ�w�tJ��R�� ��6v�d�0)ż�vc�pg`��}׍a�����ss7�-Y3�j�6��,B���l>L�,[��0���c�w�ȉ����T6
#W����E���p��j��Be䮼}y5�ܨ 5��+��wu$�5���q����d�ɚ	���(�r������R.=P�����~6�t���e�u���f�؝���Ns�u�"n�B�	g7C�Ih
��^��+�3��)�]{Y�������mN��=B6d�(��=��$<���Η�&�OT�®u������;A�:c6	��m�ְr��������ef�C-gMf.	Y��+�B��Vq#���c�.���ubS%9v"�
��A؛��\�:'*�C��A��{7rGwV(%b�Fgw��h�ٸ�o� lNl�gb��8�&�*6
ji,�۸����8���k\��	� 'qɿZ�6�W��A�\��+Eˑ��t�Ţ.q���S�|icB���$7i5������ǫ"��[O�;��(k�I�grD�-�sU2O��6�ɧ3Z<�]����F�T��44el�N�a;��'�@݋����{�\�
���.%���>�v_:�e$� �q���M)f� }�_b����"�	��9�Dw��	�#8PP��+�٭��guE�VӡO�����2�-M���� �"�ήWd���CZ>�껣s����6��]F�����Z��!T�m2�&kukI{w7v��������Z*˙M��ԛ+=Wl�����G�e��2������E@�}&�˱";�e0���L�%����VB��{y�V���vp�֣�FX�T�
 +Xe
�=z�U��L��8S	�l\*�&x��q��[�+)q=P���uԌ}����v�����y���u.��5�@t�kE.�X���a����@i����汭[�3���tX5��o��y}�U�eu=�HU�{b%3R�j��E���m���ޢw��$��(�v�˩�Ej��^S�<�M���և� �s%�iJ�jK8'w�N!V��o.��
�z���t4T��	h�8��y���"*ʻ.��T��w�*��PL�A�kjac�L�݇n�Do��Wm[���/6���n�CnopTڜC�R6�\g,�>wܕ���W)�GAޜ �rn
�'jR�k_n�;gCQe���c��F��@��N;z�s�+U�')z���Yx�@o�|~����im8a]�[N�v�q���N����lsi�Y2�f��"��%GE�V&,K�WS�jt�H��}K^@��F�˘y/x�x�
���
w�׃�p�sP�G+��^/��b���Xr�8h�fS�Ӻip����V�/Yʸ�6C���1�ne�G�r��fV� ^�Kj�.T�L�����q��"f�|�[��`�f�=�Iݬ�73Z�COfJ���n�eW���]���H����5��+�>�=�9���!��ne����n%� �q&���Z�g]�\(��%��kF���:��|�nnA!��� LFe�����U�xyzh��dwm�W<݊S�u:�|mt�fr�9ԫͲ���{���3ۥaTmB��:p��Ѽ(s��q*��
�3|�o(,,o��-��N����ԃ%��N�bA��%8/(f�`�z�U������٫�R+m��f
C+$+q�;�P����a�QV�8:��[�x�,�f�
9KV�՚7d��1j�+�0��Cb�0�^V��caU����`��SEN̰h$311C��wM[��^�	F�N�����u�����}n�'K폑�q�uh���ܳ�è��l[b:ژ��/�5�4�|{kl��WL;�ub/�m���N���bG��ݙ�DAD-E}`�����g�mB����V6�mGh�2u��0	S�X�����Fj�&�JT=\�׺N�{�I˻#�5���J���	Z�u7m
y��N�"�<K1ZMf���>�8��r�Q�P8��u�!G^nI݈%.��.bCz�,��V���.�O][y��_2�e��#�ن��׭�Rp,u��Z��ws�Tb;o�ѧ�`�#)�Hg��d�e^s��R��w���(���L���/� ���H��#W�i���]\`���Fmd���;Vj�2A�7 JVoJê��Zk���H��ˢ��w�;�ڌ(��)�N�Uۥa>�$ᓛͺ�lo�yK�L�amᾹ �
]4�W�rn�]da�l����bZA�����Z�ԘӒeRw��%M��jJ�Ծ��.�X�"��i�0Kd��kp�C,+$��&-���y���eKu"�(C�@IF�Xe%fQ�ĩ��4O�lXJ����Y���X*���l(./K��!Gd��l_�6��� 2�a�Z2��Bm�E�k��:Z����V{��B�\��')t�f��K� �m�}��Y�e*�]�� �כ��WJ�y�3��҅�Mڮ Q�|����Z�-�U�*܌ְ���s�nd�r�4�̻6!̾�Dm��Wn��+e
X���Qhwf+F&�m;�\�,���Mp�[�R��Pk96�l�Z@Z(4�0S,7�Q�MO�4f�)B�!guԸ��՛��x��WM�b����8�r��h��kb��*nG���q�����r͔���dj�^ �g]����q�aK�6��Z�Ls2M�����4��w;�X8-�t&aU���Z7��X��Z��6`v�n����!�v� ~�}}}N@�����2�[��v�vc*PUt��2���V�F���G��K}�$ز��n�34�2Ǝ�p&�q����ԲZt�U��7@*�#��N�r�t�jeZpѿ��Wt�Λ�cB�՘ �u�A�uK���e����,�X���B�"���B����
j�E�i��-�V�0��r:p��ڙs�+ ��QV��ΨSZes\y�Fm��:}�"U�����ܧY73-�]�R��]�ʛ;��l��6��k�M�}�Y�ll�<�3ed�:��	���]q=A�΀�%z�m��v����7-9%�EdJp�c�Jc�I��A�(�}.���œza4]�ЫcYZ�M�OQ,��p�|
��ƙ��2��EH�K/c��E�ց��>.A�=Hr*�(���6ڀGI���ٖ��3�/��\�2�piL�J�Y�/a�M㒆B����亏�yc��˷m��;;��N1*�o�J��v�3��g�5�s;n�I� V����.�V��)�v�=�Ҷ�gu��!�jY�
l��֡jif�`eE e�v�u��ȼ�)�2�*�L��<.K%DK�퍚(��ݶ���vt&���]]����}�XhQջc�#tkq9��r�B�wF�֚Rgom�iu5��p�����D���bɸ�D�hs��\�Ӵq��6�ޮ��*����s<��i��^s �/�=�B^kr���e6�$�R�����f%+�v���'z����;6Ц����_oJ��vp=�B� �yI���y9����Y��\&�ܘ�"i��>����}q��Q:m�e�9@B�����8+��\mH�9�h�U������jt�v1��5�W�vr�,n9��-�"+�Ew�&Չ�Ϥ��wz�̮��l�R��0y�$�Qi���q��@�7A��^���Q|�-*����O�@��#I����Q��z�@���)����Rg3�����i�Iv0������̬�3t��I׶�rr��=]�'l��NG��Gy,���u&(s	Ѽ�6*J�I�R����>{w����
p!��H��R��1⭺Ce�j7/!94lq�Ѹ���{)�:�[��HN�Ә�,)n::����'�#Hj�]`8��ufǮv�]HT��9^�K�U�o[���@�&��?RXt| [�J�J��5��[E��$;5���kNu�ΧI,�9����;v��קX�Xu��H-uׄnP�܍.�74[�΢Y���~��%�븮���w+��.m�@r�j����ևqU�L��)�;)]�8:¹*�[��s0���Epޣ�i��}��Bc)	�^l1l�����H�C��>
K��#���fc�:��^-���Wn]audh�iXMD{.������s9V�o�J�nڴj��{�[��2�~�}{��
>�\��:��u���n����D:֕��A\Ǻ檓v��������T�w�'65\��0ŽC�nS���v�����(r��1O��h�Sz�3b��w��mVP�d�ͷ�鋈�4.��W7Y[�C�QWqu��ĭp���>�.�P��i����{3��Ng�j��-'���9Z��Օ7��A�6<��m�5�użV�@Y]V�V��:qw��o��(xu�B��̥[˺�X��s��f1Ɂe	��SuE�[�Qt�lÖa�%I5�gl2��I�+Eu�����9\��U«	5��I�O��Sz���{�ڑ�e���l���}i�Y�2�'<�ݯ��p����*<B BuZ��,K�=Ӳ���R2�ɬ�¥�����$��5%�5uלx|N�J(S��W�ɹ;X@�e�������qc:�m,��m�ݠV��f+Y��E��h#ڴ7Cq�Z�j���g-�-�{p[KzVfQn�]!��&�Wr�∑�h(�ɮ��9I��J|z�*�1n��Zլ��ÊT���D�wzs2f�q|-�ظ8~��y��-�	��B��tִ���6L��NL#^�r�1��mP�����f ���>�y�Oy�HmLW��)��}�Z���I��/f[�v3x�հ&�k4��r��E�@�pg�Qm<�f��-�x)�:'�Pv�Xu�����;���R��&�A#'wm@�yPK/'j�&*�8H̨ݚ3��$�9���v��G���6�>�WYY����qWz��N��BML�;��(���,�Kwkq}c/u=}Z���Moe�T�폮��)�4m$o�@������#�a1ɧ�3���Z�i���Rü5R�����A	n�l�3����,� ��'m�r��r�ɪ��;9�p�ܗS1j����N�r��-^�]KV-�}��K;����j�"�Nf@~;-S���h����5i���ќ���mw��h����_k:�E�R&e�'r����/@�C����h���;���	=%����yv]Kw	�@�V%.�<y{ZVV,��+�P��M�6������T�d�ya��5����̩�X!�ig39�T�v�Y�ne��)") s����Z����]]5S�6���1Jqw�d��6����º)un�;� �H�}z�z2N!�&=�M�j������0d����N���!p#[�X�N�Y��)�hH�q��R�غ�3"�7N�]�ɵ�K�+t�݁q���W���O���{x�u���b�D�f�SV��lC4WpBSѯ0.�Y��e���u�z(�R���=����`,�hu��o*e\�x�fd'�B��6�R��ܰTn�n}�#ZG�u�uB����g�c{�fN��B8p�>[b�Ð�ǉ=�������K�,���i�9�b"���'�cR� 0�v��d�%��-q�}!�ڎ��Q
���-�he6�jT�����:��0�H)ڭ	��:�Wq�)^*�R�L8ұ}��%��.ꃷsٱ�"sLw[�S�縯��1�گ�m�R����%�A.�,���մ+��m-��;D�yu�����'��]\ٚV�v=y�wY!n�<jM�X3���]�I4���*��62ՑN��v{VAemi�AHw�����%�t�q,�*��\媝���-��Ź9nv��Rq/^��d\�8=���H&2�7�"���p�m����
���1s�Z�s�޸����]�A��F���WQ��H;���b�N��6ޢ'�%kf���ܧj<ĸv�:�}���[�B�gQbvA�Z(˹V�X��b�wn�ة�[��Naީp�Q�v�]��^��]��+�Z����b]�\a�@5Av�ܹ�o6v̹��T{z&�g%J>�3^Cm�.2'rȢLuuAŐ�5rV=!�e)@�����w1[L�zAtɦ fʠ�5�20D��
����'-Z8�ԭ�CC�s=�ѝ�)����J�ӨCB�V7A����̛�>BqF��rPVj�yN�rWTFn r亠�Xz"l`ڈ-�Iwu�h��+�-t�}϶�c��9�R�:u��״����4� �]1{��?@�׌O
H����~on��_5��R4��}�u�J�m$3����+R�rH��y����o�J�{������z=�5�yK���6
���Rn+��l��zT���	]S��s�׍�Ԣ�؃*C�j,��!�fd�w;�b䨁�����f���I�4�ל+���ȣ�����`��;���+o��k�GS�R���ӌcJv�X�fF�㫄��a0�Tk�s��^>H�	Z��;�ESl� ����ܲ�tv���sTӬ��s��i.� ���G]�k���u� �d"8�wS
���#��ACpQ�x��$�[ً���]n��,��cc�=��A��r6�KڒX���W�I�{"4yԨ6ʏ+f�e��#]��gmV~U����s�l&j�?����5� ������]$s7z�z�&�Zj[SN�W��)ݡc0����ϟ]gV�;(C֝�u.�@I�ڼ;����]�W_;'�f*��:�u2�W[˪�r	ku�md2pl°u�mj�-K��������aX��	Lf�b��}��3��R�w0E]r�޻1��2�:��ۮ��u��.�[�Z�3�%�b�ލW#�����+�n����`k$ᕓj�.���Catog@WWd(N[�����k��%L	��vɡ	]��؇�����$�%n�T�cru�G+RT޺9�Sk5�6-u=�%�}����B�����rV�v�^%Vu�'9S��VCPg#gv�S{I�m�O&�˻�A> @$���l�]p�����*���z���Ԓ��]��QP�-U ��Ȕ�����0���DP��QAEU+rp�]ҕ��R" �]#h\�k�q%U*�1WP(��QE�d�$�g.ʽ�r�s�a����I2"�ԺIAJ#��s�&�;���qݑ*��9ˇ��Ne����Ae97*r���^"�BS2-QP�����玞!&T8�E^���=-�!��w=Ζs�̡-"+A�n��]�Whr��(�n��wu��'"����]s
�d9�ť9%�5�!S��h�d�����ԉ0�ѻ�{�L��.��3*�ETD�ۺ�%f)�:,*/D��"+$�CL�tT�'3�ab�4�U
�Uk7qt��)$�WL��H,��Oi��f��Г
��j�9E��$�]!�((����䜓,��/tu0���rCԋ΅d�s��E��z&�	�l�k��Y/�-٣���{Æ�� fʷ�3\���W�Js`��RJ�ŉ�S��ɧs#�P��l;��������7j|�P�	A���F�t)��2i�t�6M+em����vpu�'��p1�~W��@��_�mA����U��msXг�(��R�P��l�q4��<����K�>�z\_�R�HR��֕�5¼��υ����͏��
��;��O�~�r=�z�3��W}3�^�ˊ��B����*���_@���`�L�U��u��R���54����9|�/���+æ-��>�2L0Q��C��]�n��M�yjG�s�4,���Lϧ.k�OI,ѳƟF��W���Y~u>�TF&�H�wUۣ��N��秩^�D���'w����F6��m��y���-�%j����h����q��6���u�.��|-�йU�p�w�+�α��=5R�yQN5���B��A��:B�ތLρwY#5�K�9uvJ��je%�C$v�&���ƞ@\��l�����w��ea&vj�h|�X|3�)�|aO@EQZ��<c�3lo(-k��Fd��$�j8޽긘�,�"`���@庘*0D0�K6���˰��y��굎;<�ݢ�����jه����̮ׯFmc0�w��Nc��D�fl���2�����wHǬNQ-�],]��i�O�U`u	f�A���Ruu)�:>k��
�����ӓ�\5���TtF�aj�;�nv��U۷�]f;�G�!ܑ���ь�#^t��bW�Ӝ�L� �@��M1�{����p�3�I���'a��z�]�C����+j��`[״	�:��6t��x��r���.������{q �gO���6^����F��ҫj[6�{��51��Fv�Csp:�W%��]}��W"�,���Q��0�F������񗓓{�3�i�pŸ�^u���2�!���$R����*LZ�`P�M��y�Tt�IP�lL���E�T�//)Isތ����0�4���N:��}Tпj����6yDpt*�@y��^�V���̏�S5y-�kՙ^���QN��&\򧶥uWLs|~cɓ�`�YU73��2���C@ޑ�q#0F�E��dgiS3یÛAαV��"�j�����C5A�|C>��U6w,���mHMϦ6�a��$�I�S���\r��/;�/+�En0\F�-DA�ՃSR�hY��طB�/���Ӌ�����KR֥�na��R����q⌮`��t��r3G�27���bXy�� L��4^�q=���s�칧�Ku�q�R�Ӭ;ũ�Zթ�u�frX�٫���5 5��>]s3�����dN���vt�Ӛ�~ޙ�]6]�q�`ॣ�����m{P��R�m@��$���(�]�e�˫��X�F�@y��.v~s�l�cf:j���	9iQ:<�X:Udo�p�~=T�����..k6�-��^�\���Xx]�_����F-6Bբ\"��Md�ut<Nb>i�,U�,�nں�y3 �kq��ukS.~��m��SW�"*c�SlEѼm<��I�j�`
��.$sꩾ�������o:L�R�97�B25���u�0��j����{^���t����5
ԃ�
&nq*����y�BhGu4�Oj�(m��S!���{�[��OKH&\F��[�%�q���
�b���!���g�1�v$�Qy��;ڠ_^s�ŜU�	�wTW8�uI	���&��$	R�-"�����ϱ���ls�㚹�U�(d��Ҩ>��q��\�[�& q."�C
��o�T�Ak�|l�ocooA��QR4��j�؅y�<T��ܴ� ޲(8n�5�73[N� c���X^\3��Qש|�L��x-�S4h� �EGS;�����u��l'�6&�o;h�Y1r5-��P9��	�v�H�<*fz�M�7�J�fJ+z.�%�/�}Yum�7)A���j���থ�ӛ���'�!��D�'�[���ӫ����73Sy�Z��~~��Ant�7:Կd9#:���o���k�q^�L���9�G���Tɽ�����Ŗ@OZʒ�c�3ڐ_C�u���UqxM��*Wg��ץ�aj���'�7݊#H>�H*̍
vt�t���A����'�r�ҳw��3�>������fO$����=T��ڡΤE������\U!g�B�,�r�F@5���"{z�������V^W~���XM���׶��b�k�Շ��7).�_lY�	G��E��OwB�<�����e*ͦfU��`�ʓFD;)��xF� �`�	�ְv˻wd4���]w�����:o�P�4f"FOK,gD��t���8���cT;=/�U���h,�f���|�ӵm֠N�,D�*��!Q�������&�|�"fKg%늇9c3+bC|�Q����\�8�vj�!�r_���ع$���NL6���P�U+�zSs��ǜi�QOs�O(�nu�=�mi�3�T�����MZFb�O��ɠ+���X���ѓ�����C(kYf��6��gy-,��=�hBլ|+!�xږ�H�^Ԯ�	�|�<)��=�����gr���k���qu(.7�0&�S��A��o(Ť�y�oW`ԮK,�C�4V��#4��h�r
�gK%�ۋ���SX#�E��y8w��H�ҍOD��DPai�Ҍn|Rˤ�GL�]ʋيjۖ�30�i��ógN؇�܅�X���Q�RÙj�Bރ��o��fR�j�
�3��,K�Z�`m9r�G�ѧ�#^�Os�˒�V��>�H���Z�pEu�s/�Dߨ%S�]f���Q�q�;_OoC.n_���,9�{�uX�h�Is��w~�(]d�c.1~9G:kb�r/$27]q���Ju���22�J��*N�����d}7����^x�\Qܞ�ţj\�k��i�wh��;=�t9oE(#xn�V�zI�p2W�=�2g����#�*�v�n<��C�f�����]��v-^�ua6}�Tؿ��_�򪇁�Bd�~j�+�>Ә���ER�M!r�=�=t�V�Cr�<�T�+�{�Y:�c뉦v�2w�39�aд3a3sݜs�xkF�/'��Og���z��79J���4��oF�˛��sV��*qZw��%��
�ۢ��B��'%EV���n��;��������Ř���p�-I���q���M�v��ۖ�S�:_jO(k}��{z������9:���Nf���!��9�T�ɴ���I��ە��A��5_g�KZ�t���R�1���̃s��3�����������T.K�yG���:��0�)�-��3��`K�U��R��No7��:�r�-�6K���[Xw��Z'< `\����t�EH@��w������+�ݷ���|Vj�D�p��V\F;��\3��/���ii�I�x	���l|)ȑo�"��9�=bjj�hp�I���Wj��<�U�^g$Wmh%-0d�V�OY�S04�2We��ٰ��[�ˤ)�
�>����ퟨ��NM��k�}�C�>E�\+Xh�66'�d�����py�Dq�9E�#Yی��t��k==9ڸ�v��Bg���K����+�[�{n�{�+G�a���'t,HP�;*��=�����'���j��{#akM�X���8u.ދ&z���8����č#�P뤇��^��bsZ���`�u��w�;�ut*{wg��=<I�MQ�0�-<O��u|��ɂ7����v�y��3M���v�Yš���b�Ũ�J�s��:D�����W����{,m��=�SB�Q��](�E�bU�uy��ʀxT�DW�#(�/r��yL�M���7��aQ$�t��@�}�8+���ۋ�����FѮ�K �O9���vH^sT�U-�x�l���T�EA��F-�Ru-ٙ.����;ʃ�7L�քw&>��_
<>qnԜ�l�5^\,Iݡ��G:������a�*̬4�M�!���z�"�3�MGJ���P��z�$��C\���2�vl�e��Hڽ$���Z��Ş}4�� �R�+��]�� v,	3�]nS$ϲ�G�AαW�gX��ũa����ع�8O1,��Z�}64$��s!U�Y�?��m�4C�C�8)�����q3�Zb�ge�γ�	iw�=o!�#%Y�VE�#���8�1�I�������﨤bTas��N��UY����s�����-�+δL-9i�΂X9�Ĉbކof8��Z���������ѡ�"��a�L69C�m�::v�@�{�������OQ[�S�+��3"�f�n\�T@�����8t��̡��xU��U�S�-��Za�qb���$�+@@��!5*�2�#��?M2tC�6k�z���`���:i��{��N�u�EJ훐Ĥ՟��I���J�Q�N���e�m	��4����v�X��sN�ɦw8�fQ������3����P����w�h&Dq�4e ��~�3=Z���*�D�.\/�+�e�g�1ԋ�c9YȺk��6�CշK U�� \������A�g��{��N��t�o�l���ni�
��1,��7ct�q赜Ӽ;Ӷ^�\�5�Ƥ��K"�����*�
\�P��';�e�6�B{GH�6���{���!��]Gr�.���s�&\Q
=�N�0�$BS�D����T���9�4V��lSb�w�F����|��Ņ�\�8�Z��(
 o[�,n�{s�Ø�j��Q��Ó7�p���\ȗp�Ѓ�$���E?�w�<�MgVǷwލ����S	_�9)�[�ld��)��8���p�ޑ����6�2�!AZ$]tK���r��>�;���8䜀nhY�أ��l�Gc6��pk��:�� �ws7B�����RX	�Ru鋑��g�B�U�&����]���-"��|�Fˮ�Ю�v�\�xK�Ͳ�2`��N?45{콓w�َ��cЪ?����Ʉ��E�\�{6�����H �GN�88
�*��s9�c���k9�o�+�ԅ�Э]�sb�Gw'5j��@�}v~�K�Ӏ�-E�t����kO�����N���S��#��2�xZEwfӰ=�X����_�g#�B�*��Ԏ]^�	���*�ټ�Č�����2'�V����H7��_x./�O[��b�B�O'��-hn�8��[�ƛš�]r#���0�vPZ�w$�̜�vMn|9L����ZJM�;y��"�i�V�6�L�.Yw�4]�L�2~����N���K�1�J���}�q�L!��s�R���ڏ(�f�l�.�&�|�"fKg%Ƹ�s�ę���*���s�էw�C�0sq�6hp1�����L���X��)����v(���@l��5ٱGN�<#E���P�nC��ϊ��@pI��4�s4BAQh��r�{�6�����3��WuN{��C�џ'S1��&�:(Q���LW�O�D���$vn���uuo+i��Q|���/6t�}]�XJ�sV@�$s��|�Z��-�tj���Rܻ�soC�su���q��ck�q�B��u���]nT�mXc �@+����2	VYƓ�����t ����k�	�=
��6�=�y���<h�1�}��<��$�Ng����I2휭�u���jid���G��r��Vm@�S5�Z����&g�����d���3򈛕��K3��㇯���^5��h>�PXn=��$9�=����6�csE�bH����|-�Ԭ���:+�/,�8:��Xn1�,u%T��l���d�aa���i��k��m��Sy7S�ʚ&�t3-e�O\1��19l��JM�zd��'u�.q��{ԕ�lڭW.�΅������"Q�d���Icل(�)#;��V��I=.J���8]DU�cʡ��n<�n
�
לkՇ���{�㳀�S��C�� u.:L�'��P��2o��ER�����8�<B�n�g��y��xj��7v>���3ۍc��es�b�����<�����VN*t���˱�5n�@�穛�5�Թ'��� �ǘ��i��l�ƺ���V�-\=�ݛ������_Q񼨌X)|�t��c�a�zM���Y�󻟯`Le�=eE:{��'�1��~�����۲�ln|�:��Ĝ9�#�,�<j��O�R��r�;��E�����4{cvv��9yx��J�����J��$�K�T=���H�=�9Hz�͞L��y�T��ɉ�7]���]�����ג����Z	<f����K�w�z����-o
q��_�I�1�?Q��������s�p��Y F�g];�X�9���]���t��H�[�-��7�:tߣ�׫ǫ#�>�ď��%�LLRسF�Z+�Z�.�8k���_�-&_��s�p�U���A@`D־�P�B�t��`]0��l[�J �)�`�����!����.\�&���\�oةA7ޛ��b/���%^��� YT��QQb���{u�s+���4&��Xh�mn��x�*T���9�=����jƮW�k��i�!Әw:��ǵ����d�ձ,㦲�h؃e��Y��&�V��K:�M�\���O����qh-c��2E��Z�%E¹��`��d�����޳ϯ��mǔ/�7�V9��u��n�L�fT��Rr�*��L����ټ���+��h�uyK��ȕ k9�i�so/l���LyOR��B�v����#'�us���wk��2/@����=���sݬ�le��]�,�so������	(5��܉c��xܞ��-dl7�եg
����7���ᵌ���͡��9�P��Ǚ:�˺�7����@��G9� ��mKy�I����Ǐ׺Ճ��E;엍�`��{nei��k�
"��)Ck-�vik/jf��\ޗ�c1��q�Ge�wO��ml.ui� ���kL���}�mM�������Y�o+(��� j��;�De�����^m�/���R�*Չ�L`e��'�gqJ#4��q�=��
�CO-w�4��7)2���׼�L:�ʻJf����;�7suYe<���Щ�櫁Sh���i[)+��E���z4��x����
2���ٻ���U��S8pƲ��Wq���F滔�=9����;@�6/&��HPgN���9�zR�$�s��s�S�l��1{9J�������GC�K��c5�{Vut�ǩuM{��Y40$��1)��{:Gʉ�77Hy��ѯJF���F\b�q�D��.V��fu#;V�"��u���e
�}�.R���a}���$겛���*ʼ������x�����34��vr�S��y�#�+�0U��&2kogqu�ț[X����~����uzS<�n]n���8gw*X���g��̪x�L�ܠف+�\��a��&����{��lRr:���E�J��Y3f���e��|�.��س���f4&�����t�ݷ�[��W�7z���GC��9��-�����q�&fu ���@�n���l��QY�]D+nKYt΂�ܳ��x��H�����;�[]V�m��B��x#!�ז����o/�,��[A1�Vo�2]��lvh�8���,�q�vNƚ-_`s�󽲶A&opȚ���;]a#��*�5t5��S�<�H��@�1I���Wt��i0�9��En�:_ �x��kz�ҭs�7��6o�3]��ד�4��v����V=̥M���k���#�;�`^���'#�V9�@����s��Lk-t�yԓ�����>R�E/ir̨�Pc��Y�wDO]�0�iRD:�KJB�-�%&YJVaEG�r(/(�EJ��랡�[tJ��rwp(�<D5R������P�B�&2�R��1,H�sҏ6�b��2�s���rS�9�m
"�0�Lأ���Y���ʍr)���9����Z\�Q�rj�k��wg)�	S(9(�m�ʢ#�T܂�D���AAZ�EF��;�Mu�U�Y�0rp�
�2�����'P�)�`mI�#D�PJ��"#��{I*���A� ���4;4(��QA(�D�F�(äRK��D���h�k:�j
���]Ցʍ@������A*�U�;���djdfm<<��S.DZ	��B�*��yJ�Td$T�N:�DT�d���h`QT�)
�x�"/7oC�/i�s~ۗR�o��Oz������'K����K����`�֞;��7Mh�}:͊*o�G!m�A��l<F���n��2���xs�I��lx~!ɅS���"��P��4F'~~����ۓ��/zZ�3��I$3�/���@I��1��#�" �}>�>���u�M��f<M`ŏu;=�w~�1mۓ�7���M�	����O�|���j������	�I8S}g.���������d���������Ǆ���ro�`�}O�9=���>��I�O�#��O�s�/�轿����W��Da��|�����xv�o;����]���~M����7�'N׺}}��ސ�x�`�����y�-���8\>s���~Nw���<+�q�w������Z }�	�jP���f!(��gC�}>��(�?=�'��_�}>��q���	�!8>z��>F��'>�����'��>?������oHN�/�nNM��|�&�;|O	?�܀�>W9��TQ�x>����0����|~9ӽ;I�?��]�����W��������7�/6��N�����|���S�8�������ra|��E��}���cުC�I�/� (����>�A�b��P� ��a�D|T��9��uX� =�N׸?Q�	��~q�»�� "�D}�0}��DX� Qgނ9P����7�'����1;���~}��>���?}��o)���}w����O�$z5��R߄�}q}�����|'s��1?����ǔ��9G�����9=���pxL*�<W?�?����=<��2�On܇�wp}I�ݮ���{��7�'N׿��<8ߐ��{��{�}$V23I�z�����g\>{r�� <`��t	>��"=�i�����$� O�׾"Ȣ��hz�N��;����X�<&}C�����P�U����?���o[�px���<G�"@��>��ks�'�Q�g��e�q}]z1}$z��� "�ہ�'���A�Lx��qq������q���O_,zw�{v�z}�ޭ�;���y�M���o�_ףŃþ��y�z<;�yL	�>t��Q�D>Uv�k�#W��6�oݰ��	>� �4�@��nπ�1;�_���v��ogϽ�;��n�㽟���aT��|�G�����_����;x=^��zv�󿝯1���z�H�^��@G�����}X���4��˗�sP��Br9����3Ƹ�C���zbH�e��	�įf3:��}q�>�Z��o���Yo:�«��L<�PzM��`��T��@͋���Ǒ+n�l9��2q������oUI71�ŵcջ�)�`��p�*��޲�����}��{�"H?&�ޣ÷��˽�����S
o�����yw�k��t��r~M�9���`�����'���?!�0��������4�@"<L�ނ���y�^T}����?޽��zq;N�C���[� 4���#��ٹs�z#�@O���}� ���$qdzϬr�Ͻ�K�����N��kϳ�����돱ޝ�L)����7���7!���<�� ~I����7��oF9��>����@�<���~����;HR�m�ӽ;N��ސ�������6�\P�W��gv|/]��M;�ɽ��q��bw&�y��.��S���='��C�y(?'�x����Q�'��7�۷'!�w>/z9a���<	�>���2��i],F���*�:��FO_h��ޢO��ӏ��}�'�����{q���<����v��G�1ɤ'�~q�<}�N��_ ��۟���z��;I������t}��{v�7��<;�|q��7�tQ
��·�t}o/j��H�'�F#��@D
#��+��H�>@��`���?��/������xw�k�����oHN��}���bM���xpM�7�9�÷ }~���p�v�y?���=��*>�\K�ɝ]<,�>|�*��Ȃ��tG��� |}\���<	��)�Y���@��,w�$y�������x����O��(�8DH��"��2G����xAG�� �d59���fOl���k_z�G�Ť���Q�y	͑@��|�����ȏ .[{w;�ߝ���]��޷ߟ���N���|�ǇxNL/��x���zqτ9[��7�=�����_N
�{��}�����B����Y��~���G�A_ ��!H��w��<��������{���㷕w����c�yO���w���ߐ��o��z�zL)��?~���"�|�>�y%�q�$�ȇ��C�\;�ϝ���i�y�(����>�#���c��<�õ�y���ߓ�r}q���]�>8��=��L)��~G����w�G���|5�D�����z��${�>o��qk�9[2f�/Շ	�P��\�u��\�y@��'}�ʵF;�I4w����vFVb�Z7ax��s��D�����y�.��/���e[���|{���Y�v%���|��KQ_,j��Kܓ������լ1	�7w"]��2�!F�ie��c�6��������|xE���괏�${�����2>�	�;H�<�ߠ��;Hx=����\xq+�?�ro���8�]�1;���'�=��������;����Q�$�i� ->��1��}՘�DnB�x9C�@�>{rϽd��g���A#�#�Fw�(�O���"���S����xw���~O�:w�Oq�7�.��w-`�}w�����	�<�EM�s�_�&��V����Y��|Np^.w�S�s�O����(z����y8*����o.��M��nN<F'z�m���}���I�S�z�cǨ���!C�=;r����|�?$����]�'�����3m�ߧ�{���'ۏ�G��7�x�?]��{�O����o5���xC�~�xt�&�����~v��Ͻ�7��s�;]��\�}O�9>;������]�=��xOH|C��*��6���eh���Q��`�Q;�Vϸ$��>���x@���8�Q�-�ۓ~B}^x��ߩ��ߋ}CÃ�}��~���.�����.N����������]��nM�?'!���F��߷>�n�����뛅����G�����yC�90������ÿ!�=�r���{g)��o�w������@B>��|(�h�|d�b���I��P��G����<��>�{�,�O�����l�,���?q�9щ��껬���:w�{��i��~߿w�p)�;��8��{�N��<���9�ۧ}q��9��xL*좜Q�>!��X���yw��n~�}��)��?[q�����ʣ��x��~=y9?Q�$���r}��=�#�t)���i���y@�O���}�㷄܄�;��)�\
o�X9�����O��N�m�����>����C�t}|9w�i$zr^��Oٗ���ɸ��_x���i���:��Hg�����#��I3��"� �,G@�O�#ȳ�����($��?~����;˿��<y��nM�>';�����l(s��|��[��ʪ8��}�����l�)�����>\.I��wxM�>'8��S� ${HdA�k��hx#�@��=D?!�90�:��n�~w�9/��=!8������ѽ'��yO/�n@ۡ�>��f�U� q�d�]�/f�'Ts-n����)�䫺���W9	}�B;s����P� f[�9��.�>�e$ �uc9��u�0�Z�ĭ�JհuZ'VDг����N�W�����P�/
��]�*t�j��9^�<z��FI�'g�_����o�çxC�
������7! r_���ü�O�����GoΝ���=${��{����$�G���9�=����~M����9�X]����,ˌ��~���gs���ݶ���I>�#�'�<>o�m�;����Aw$�O���	h{G�42�F�y|��w���m��}v�w�}���'�o�>�>��"=�_9���$�@}ݚ�[}���o�ӻ�5��6}�"-{�yt{þ�U�����P��t�'`��r�v�,ro�;�B�x�N��|"�@��aG�>�2�C>C 2|�c�ߓO�	��<��I�����ߨuCIK'�/�=l��I���8�}��>�Z�z���H|���" ��$�~Bp{o����yw�i4�O8\.����~NNq�%r��S� ��0�M����������>�T��}���h�Ҭ��	���z~��z~������}#�I>@G�7#�@�<!���ȲϽ���(�#�����'1{�zC�
���<����z�������Ҡ}Hv��'˷&������N~�uw=���wޣ�$�G��C��@V���Ǹ�i���D�����s�^���<�v��Ǐ�����X;��G��G��r�(�w�v�������}�T��toHt�}�ӯi{,�~hު���*~��w���@�I?!������o��x���޲ ��	� �>������]���������C�iӵ����˿;J��ɽ|������ݏ>��#>�)%�3�ܚ϶��9�$I� ��o����xC����ە�i�q�Aɇ���|v��>O?8�v���ݹ�}Cçk�8�_�o�N���<���w�i?��\o��Ӆ��0�ޘAz�)��	E"�=�/�A���A�de/I'�=�a�p���<�f�T�\��W��Y�|b��$��<��#5�ͼ����}�:��	yk}�}�gy�R���p���"�z���7�.U�h�`M�jOd3�u��R��qVߟa�ݝw�$��O91�J�]��؀ݑ��ޥx:�����v�:0�;Y�9�oo�m�]�]�¹�2^&�qtM�*�*�����������	�b�[&�FL"7va�TƇy�1�C�M�aQsQ�45�w�z24|��3�_7��.�x6	���'R\��� 7�\m�����U_L��OS�3@<�r榳�J�bXz2~�´�K�

�bz G��2��7�$guG�Wv��)�
����Rc�ZN�����lt��r~=��=��4=�kF�i��Bo���k��3�3
���'8�F��ȍ�[��t������6��{Nw�%醳H��y݅��5��w�HV��9z=�N|H�,&��=flU��WYӶPkvZ�N����`Z��Y��,$Xq,�isTM�N��2:
�j@Y��8���Hq���׌ֶ�h�tW�.#�L��7#�H}ӥu��$ᦨ�NW��"e1p:�+��n�]75��4��$��2���S��ѩ6���>�'z�]Q��RJ�k`�1�M��'mr�|�nL8�7(²�}���(l�U��ĝ��>���zL��8@�y��XV���/OgC�|�Ea����`\� u�4ӝHW�!���4x׆��<�4�w�2�jz���7`n�=��I�F`*u`m.o���+C�]�����W�������uf�ѹ~)�ǡ���iX�[b�!�+D�*
�t4xr\ne�t�>�o%K��ww*Y�2(�31JY�Ɏ���2�;v�Wwv2WD�g�`MY;٧�����4��� o�{����kqL@��~*�Q2;�¯rY'F_H�)Ʊ.���u|l�et�D��)��u��rc0�e���A��n򊮲Ϲ����>I�� ��9US���e32�s=h]z*������)�碥lX��M�ր�ǵ���y����*��{�7Hp��	�S+��s����ϫ�EfO:�0�l]T�I��;)�4������B�sT�\m��9WUS����eȿ��a�L69|���b�o]��l�W�{=�SQ��A�x	@���1}�iDT�F�n~�pʜσ�Cp����8j�����O,���V�.׸��SIl�d�+w���yR#��o:L�*s�-����s,����vW����6��4�R��jR�iL�)�Ĩ��v�{OF�lDږ��=]�>Z�WT�3f���
e|3�3�R��PL��a�D�#���	�¦�n!ט��q�^��ĳ:�<�Df�zO�92���a���$[G&J��*��,��y�z ȭKdt�L���Z��'�L�#����2�m���7�5{�����[�G}�!*�'����䲍����;H<A���i+c�ðmg<�؃N�I�;��X��I8����]�E3��-��l���z�����$�(M�Ѩ�=c�9��?���JZӚ��g�9�1�9���)1g4���zV��4��\�Xsd�q."	�'��\89N��{�P6�(�.�\�W�4��k��(=������:4�!!$�P�n�5���f�T�����{'�z�\(��	�B����4�_l��<}�wY?)ԝٕ��K���]��M綣@rW�[?�����\O�
��h�jAC�u���w��پQ����8��b�ˍ�T��NN�b�au�H,�hU�&X0o�9��Rw=ǒ�Q����|�t�͍��	SB�6����WDh���9�1G3�#X�T���FS�|LN�������k匝t]V+
c�&�� �omq.#yr\�mey�mlV) ��,��`�cL���q���U��8b&��L���Q���:Itr>��`uK�5��;{��=��#���;a�^���۩u%�3EF&k�aq�,��[�|M1��9��{�܋m�)rZ��5�赨o�=�T�O��������\1���G�R�9uD1�M׺P��j�Mȴ���H���9��s �DQb�*�P��HG$h��8m��(;9kj��M�B9YK��:�	L4/7Cs.�]���p�ǝS�#��Y�72-��	<�D;���u�a/xbH}$ܺA���<�CЎ*gn�xW^^��s]�L����8�}$����ؔ,:%-[������L�*[O�gfcT�i5tp[x��MWEhpF!�̻W��<�U���W��Q���-�l{a4H���eY�:Ws������p29����$ޭ�΄W�8�	�㸟"Ft6D�tP��UH�8!앭\�vv�u됨�z��ǎ�24����gN�>��/�V.j����Ut����:��'a���E٫F_�y�L#s��X��Fs�s��9lt���ܩ�ڰ�ilCz�3����o.(^�=���9�dj�q������?��FU��iO�_G�Ĺ�6B �l����Y�k�ݳ�u��q;��IO�"4���P^*\����Õ�y~WL]i�y���5��q���S��d\�*Sr_,01�~W��@��Y������hVcw��ñ٪��!]6ʣd���k�W�$��+׃�dϱ;��A�s��y�$��0)�m��Ȣ�����a�\u��p��L^u���UC��>L�c�{�����1�����*�]B}��;��*�bV��T̓A5��5��Bz���a��!o�L[�v�̧t��c��n#��tv��a�s����Ү7�eί���L׏չ�תS�J":�{�����k,���ˏF����SFT�5)�jf��N���������]�vd�[�_�ą��zŖ�.W��\}�L���38�0�.!��7� N!9�����#�u�cG��,5���&��;S3;sX�K�xѳ�)��(5u�<f��r����c�.�~�fg^[Xg��>�W�/�*�X�/'0;��8e|�<̾��Su�W}??�kLZ�n�a�sl��;���q�.�.$�#|n���g��y��qoU!�!�C���k���z/����;��q��Ŝ�I�I`]�$�x�X��Y�s���l��Y5�\Õ�Ó4u+|3�K�}��:~��
o�

|�*4d��e�z���	P��8c�i�����1Ck��g9_WO�@]�M�󩵛�ql8l�����D9y�{&�C���s���궈��B�'v����+�
�zzr�W�gNr,2��
�f6���]R���.00����	-���;*��i��cÛ�c������q�=.7�ۜ�7-!G���qd�s��ͣ�1ؼ�&���m��y���E̽�����<���8��v|��ۻ�rS$̩��(m/�٘BՓ��m%��r���=dR��#20rj��:���6�͌&S����V5�����͌]��ruD��#N��+�XV�}��x	���{��b�'?{�y�����t-}ӥu��Ĝ4�sN�'�@��,@0�،�w���m�x	��O��7��cH��R�������j��B�fg�|��Lp� `��b>e,O���+�a�z����gc{�}z��Ѩل�'�8��������Ι|񬁧��N�g_n[N�f�E.�.@�X�T�z͉U���S����xME�9b�+��Owf�y��ՕF����|�}sFL�똵CK2�{�v�Q�bL�WCr�$>X4�i�������r�E�l�Qús��9Ĝ�c.<��BJ�\N`5���?�Z�җ���b�<�A�q��u���,�·���P��eo4zc��8.�o� ��R��jK�a�]�l�~x���>�t��C�tuи�ʰ`�W0�~y9�u��mKʢ��V�7�wޙN���G��N��0:z ���%S����+Y�l�r89��鰲��E�!�i9Yy�)޹�bd-R'!�i4
d3#c���WPf�jv�������&���o��ܘz��);�:8��Ȫ���z����ڦ:��vK��7X����;ȟT�zӤ���{���±�u�n�U�ڒ�!�"ZA�.��z��	9�Ok�׷n�W)gW7L8WK��u�q�7�y�6R���Tol�5���Ι�;]9�Z4��R���ϙt23 Y'*dJ�d�Vz����ciν+�"�әY��٨���E���ж@���T�b�PqB��#�2��d`�%�Uh�7b�V�J냺*"n�C7��f�=ˉ\+�q{�+tv�e��B/3PDF�����5��������J��[��J���lB��f����#��:]��Īȸ�'�%ּ0͢�v=�0��]y������W�e��:�.�g<��a��f��U���mgR1P\��iWK_004�Z��J۹��8��X��3�-{�akc*��p�I��Cٴ�i.*@���o����w�5�Z.�=�|J9�h�h�$���R��+<��ko-�r=T�
����&��]��9�4��qRaF�ۯ���������G �0���k�,n��Ϟ��ɗ2]��IR:w���.gN�<r!�N칖�F�sGjRɇ��u_/�f`�o������I��g��[��gF�����VZr�]��7OU{S�uR!v�����vT�u]��3�����g�1y���_5�n�¶Joh:�"ڄp�ctbI����uu>�j���0�4��*�/�ZR�k&��v���<Ҡ�7\;.�+Q�nDt(�_n����hRr�C��(�"�%wwJ8v��j�Į^��FuN�0Yg���w��WVeҎ�V`䛱�߭�7x�6�2��>�K͏�َ����\�����ˣ����*�ڄ�������-n�9_-���<n��qv��ga��x�$��]�l7;y�G����v^p���ooQ��kk���aL�X�u1��6%���-���e�}F+�{b,�7���
LS'�es,���h��k�&�n�;*3�}�,� (����а�[��w��)J�?v�F⫥&^Z/�#c���㥙:T@���Wt�Ạ́�J��o�6Q�.��'�%i�sB�5
n�Cf�����&^�g���eڳ�����w��#'���e!}Nh�{���F;v�%Ss�dځ5r�HT�iM�/L�2\���Zr�94��N\��:��9��7zaD�j�.8o���ak�ub�ղ��jιN��Ehgsk�mi
���a��dáfi��H��[A�$l�+&���xMFVD�����;j�D�v�@2	Ք���QXz��N�4XI��誝��K�WF̿�[br�}(#M��R��ʺ�-�{x�G���KK���55�s�Q��a�mlq�+�'�9�q��b��r�p�c��� ��L�v����1�v�����nn��F��&�O��ub�eõ��[��t-��V4��\���aԇ�M$R#P,�[�Iy�W���;��[1�@�$� �9	\��W��9r�Z�4�*,�xqt.r�"iY��(��5ZE��<!�R$�+	��G��z�C��\������
�D�y��l�	Yh���w%̼�ʊsww	�8�Q�vy�DVd9�҈Q��iVE�lYEg*�X�Ds�u�j���aG�NF��@��4�5OqwS�-����RG\�"�7WZ2�G�eBG��t�f���ܣa:�'wvz\�<us���t]K3Ds"]�Ȑ��
�8��qn8�NV��Y�y&^����SΞI�5��4ڥ���EJڱs���3�&^���ιYh��\,Sww1�P��S�t�PӮK�UH�2�ܓ�Į�.r�6��璴�K*�A�j�������n:ܑX�xd�/�|�=x�݂�8>�SP�|�E�BGun�0�Ӎ�V�HO��GG�gP��-R梫p��v"�s\ɩS��������9טh�W�
�A��E5�2F���N���;�HMJ��쎗�zz�1�ڨ�}Jz��A��nw9Zrնs�RhҾ�ҭK�!�5	����I-�$�&Oeq�Z�y�E�oz���(��'�4�N��c�É?@���,č�[�Q,���!��nV#��9��quko��
��	��aoI��e!��L60<9"�h��`_T�15,�av��w7��u�����V�"���ơ�҆H׵ҟ!�qatW%���{Ac��1�Nb�Iۍ�KMUK�(T��أb/�q�V�x� �*{ҏP��4 �Iء[=ieۅ�g
ƋoWu8ND���R������Hu �쌝�J/A�s?t�apT:�M&�1���q�1�}��r[=��������=HWG��c��g� ��:���,���d2�ֲzX��מ��u��������p�V.!�#���Gye�]��yf�����z����#ZE��>T/+k���_D>�sLs��p��#8��AF���Z:vv^BVo7#\JOv�v�̠���V	M(��&q��C[�n��GM��<c4g.ͯx��Z��Ǟ��+��X��z,N�v��S��t�+LV>��Bٽ�b����
VGU�fƆ.��d�qg����sVP�/��\�U���Q�������آ=�R~�Ƈ�1��Xt7'�|U`��&��w�%`ɶ��|��Cb�[Q����F�OwW��p���]Di���������-V@�fU��9��*��i1�N̚�YZ���in7��(`����	��R��P�H*13@�."FT��f�l��f�p��5�zt���F�L�������~QZ���0�
@�����U���#z��H~�i���i�wv�䢮��Jcvu��*��3+m:�b��ôj��Iʏjd�� #p��_������B�%}�Ÿ�Y��<�P��^*���9A���*R����'ai�#Z=4������VZ�cj����<�9�9��urִH��6~tP��s��(�l4]����r�e�ճQ]��X��d_��C͞�	��8�40:��'9�s{έ�ğr��@tp�B����M�h�P��&�ӑ�-���:4�$k���k4zN�q���ڳݷv�� ���� �	�����f6Бsz]ChE �Y���3�ȑ��g�q�|�y_}�(�����k8H��轔���\C�7������Yh���i�{�
���]�Ico���&7��߻��n���}��D0j��3m�"�z���fN�!�x��;9�Y+�b=�Q�U��W7��"�,�۶oM/�$�e�5_UUTSW�=_��sF�g�ݘ�ny.�G�bE_ ��H��`x`�]{2���4ͅ���h��r;v�"q���sR��%�}N.�;�3�z��{c��y��xm��\�1G��2���#��h���n�q��L?�b��oH79�>�\�T�9����^�=]J�v.>��|)�;�����:Ѩw�*s;��x��W�9N�P���k�`�B�Фgrem�mC��Ptx���vеc�n����]xnK&}����c���
�W3���p{����I�<�M�0�R���5\*읢���<�s��	Bǀ e��8�����F�6*t���2[�}�9�yma��>�~bQ8+��$CjF�Y.����Xry� �Y������
�%���G�܍�EĜ/�wƦ3���I"ݴ��[��
/�ơPS<��Lr��њ>r���&Qs����
��������\{��숤��ɏ�ɭ��8מ@\�r�&$cuڬoA冼-{M�<��e�Q� �*�.�x�-�-&K'�FP�q��T�c�c8[�{D�x����u���T�6WG�u�c�[�֝i"�$�.�g$<xX��ѡS�Qm���޸\�Pf.��ÐS�s���R��КKk�'�6]cYcn�ux���w��"#�޾�ˬ�J�w�!�L���OW1W��\-'X�l�F 6:ry_KՆ�y4�j6�����9q�G�#D%��Nbx����3Q�O�t�җ���{0Tgf3W9�+���ķ�B�/V�u0In�bBo�h0�K�~�u���33\��� ������L�]��-)�ɐ��C#��y�+!��J]���]�ӌ`��!��!����SQ�T:�O�A��<� �+���T�\O�ȭq@-�m�n�^r���/���oc�R�����F*LZ�`P�M��nɕ�N���Pݸ��.�5�bQ�WD����S��^/k���ؤc�5ʻ�O
�{�1���+�&��u���TGGB��a�9��PUc�U��{`i<��f�k[��?�bҬn�}���ؑw�\r%L,|~cɞꈥ��vW��v�Q�bL�W���c�Q��dv�l�"�f^n�r�1�WBg��j��ܯ���7�RvD+�h�N([Y*�l�iX%�
7{P�Y��ŝ,)��I�!�!z�db�Bd��=H�}k�܊�9���A������7\�B��U�5fR�8U�� G���>�ѫ;���F�*�LN��V�B|���ȝǚ^Ҏ��1��z��3c��=���xrż����Q��08����a��z��o9�6V@ৣ����GM�ެ���]�S�]��f�8���㩞@0�<��v�]{��F���4Üc�"�.m���=�ty��9i���zdo�pń��Z���2�\2���lr��T�Pb�|��r9C{�p �6`0`�p|�pc{��ݵ�tT�gzz�;���ÌgѸ�13(g[�v��w�W  �45rKd�wz �A���/a�;�E�e�k<�I�<�p����:��Rp�k5	���C$�U�\�hLne�m��2pm�j}��l���4�1ڭ�aĸr�%�JԎ��
�>ܞ�?u�'=3�k���.]j3S���R�L�F����s����*�` �AXV̹��ǚ�u��W�����ץ6����6��5��P�^�J�>��q��)����v��|��҄���h����@�Gf�Źdզ^!Oa����Ѧax���72��T��cP������ZR��^�Ý�ݝ� `�{bV͐6e��ڵ@n����ۙ_/��fj�	��76���{/
�����{�Ϣ��������Xu��V����r-Q��T/��u�釺�TV�y�j���=�m�<H����/��\���&��C����I�ҡ-�[&��J"���y.{�@㓉���:i���n��3�̨���m�q����6���� a�}�-WCx��hg�!AH^Y�yd�]]�Z�+&��c�-��7����<^��u��ƐUY�ЫL����L��ܝ�g�2HϷ::�W%�S��z��;�q�����&U�����mY�����c�P&�yჵJ�ӆ�����r��h�X������~
a��8��V��ngyrYgۏ�W�Z�7�O�n߽E�ޱi�j��\5����q/t�]c~��|e�φ�2��ڇ0yW0�Z��mܲ�_lw'7���P�)���o�m�X퐡���4f#%�i�Κ-v�"t\f�%,3�6�V��1*|Oe��!��X�T��*u{sW�F@^|��f����k���iZ�G�k9�QST>��#�/8@�t/�����iB���P8t�߅}/�N�傪�A��;䋄�^2p3���v�������H�V7��B�Ix�_l��Ϝ��-�3�6�f��p�m�&"��ښؖ�X�3:q�y,>9	�Y\%�ښe`&�Q-g�H�g ����M:7,�z�ԏ`Yh�*]�-ۛ&3�P\`��[ΛK
�Mp�B��;[�}vq�f&ehK*=s��T�����E�ݐr�X�L�\n�ُ��L������$�G���d#m=y4sU�_:�աT9��LƖț���<��]�V�3�;b
"<8#���j��(|�C5<�Ӛ!�w!a*��@0U��਩ח���5cHƂ��Pg��� �<�$hB�ؓ[NGeq�X}j��YZa��Զ%�g.�vX�v���\�Ѓ�0L���O�@ޠcm���g���(oJ{ii�Z�d�<'T�v�*\�5�m�%×�Ċ$��ZYeAx�.��E��y��]iT���v�����m:�[���l��beIN�·��ܘ�c鮦S�oq�]oQ�N1r+��«�I���t�loܪ6w�[���\����r�|:�N��^ޘ�{�mF[�7�z\Ig��`���Z����U���DoRc8��B����|�<��=��wrZ�B�rGwV�V��p�0c�\�.��5l�!j�J����O���������3;�=*gg�i��2*5}��Gv�oP�_\�*hw!@f�Lȝ��V�'��.'*�I�A�e�����l������.#cal5"��ֈ��e�׹�,�3�)h����C�p͌�3f�2+k�U0T���}�רޚb(�>㵩LS����,ϮGqH:a����(�S�{V�i��KYZ�\��=d͜���-B�9�����T�sfN�	3&��>�v��.����~l���[�8q��.q�����le���/'(i��D��06��j��sq�'���Y���S��p���^���+��zpN{_1�3�P����*BQ0�#�/F��]�w��y�������n��ybyř4�j��Ri2k���5�dqx��ǌM=J�bXz2~��X��S��Ŷ��GSR4�Jm: �+��K$�s�cyEb�׫�&s����� .�΄���9��䯰�Z�|�tu����_:�1���@a�!t�x�ķ�^��H�����p��c�g19���N���{r�N�T;�+Rr�jS���1!_W3�f��9�zWNc�vm��s(�v�r��C��8g_:f�t��4ZR8�gΝA2�#��՜z�̍�s��ZgM��3��0K��tȸ�c�%^�=�����R��J�=<I�A�&<��R��(v
$���כ�w��~�QFڔ�����V��Y*��z�_ez�m��9�C�fg��:MV-������TvM�u�1�a��v���.�{������+$<a�e�'�L��6��wR����TeXO'�Wkq�dAZ�-��B���_NַE�$�/lhm��Ԟ�(Zw���KK��\�]k�"@����آ�:x%�kp֮�B�xx  �v�vnS[4)%-�W��>ʝ����{\f��8��;�}v�v�v��wNz*�i�)��4��Q����ad�v��C������VZC�Q�m9ԅ^C=s8\�������[J,MI��Wc���T����0ܙ#z�-P��̥�]��@�H��:�����n4�*���L���ƚ�5�N��|*s����٩��@n�¡`�j������a�^��'�0����Tޑ��ܓ�I����iwG��P��SC�E��^�]�K�f�|��l}�@�@u�)wn�먆��fe\ �%:�yv��q��F���*���E�����Z��r&�Ut�E� "�(�Vʽ�Y�*�cV��2�Xs,<���m5��伻��nΨٿ/P�c�!j�=���� �!�ɝ��~w4���3N�^�҂u��=����.����t�\KY>|�v�Q\��4��%�R���uS��P�{�I�/v�)�l^�|L��#8:��&�8�f��y�c:���*ԇ.C�V|;aC$諞gw���^�w�1���[W*ވ��i��Q�����0�N�-'����c�1� Q�ǞH�V^={��X�;��<�ي�6��+w_�d�`�6	A��N����\��r���jn=��,F<�mT8�j�K��X���`��B��1��E0\b���� Dž���7����D�1��I����i��U��?��"�|�R:��?,x��qG��j�a޹�h��%�t����xB#5O�i�H��ڰ�,��z���sd�F�
�A�ݹ����=Qvt=O0�nH,�hJ|���ڳ{��>TsJ#^�J�N���]�nV�w���O=�mCŗWW��V�r|��(�[�C]�V�׌�x���kޔ{���N�f�im�]�Ѭ��Q�{ʫ=9�b�(����ǲA]H+{"�Î�8�aL��u�6���#]�u^�M�T�q.#i������ e�'�Z��Af�i���-�����w]f�G�箺'�ٯ�ӛ�K�����A��~b*u������o�涷���s�|��������)��Y��|�'g�����~h_�Y��������~�Z��eo�lb����a�hHK�HN,�7U����MY�T��g�������b��Z#P��/��9�j/��a�߮��j�� ��!���l��R�j\�q~Y�K�Uoϒ��Ƨ���<v����.�4»~3��T�af�A,l7ػn�:@>D��fKq*C�A�\��hI���r��(���Ʊ�1_c�����6��bӅ�Q5nt�sX�k�<D�'ffSi˃xf�ҖRѴ�W�̃��Tt�ռ�6Р��XtwI�F;�s����uq��t����1®K/i`����\.�M�0d��\<�'�2X%s���ƺ�ܖ/SR]&�=h�\յ�+K?4�����}��im�ȟ����_h����RO3*Ԑ�����7��j�����;1�s��[��Q�}����=8��p�Z�/����A�Wk�E��m��6��಑�brN��K�A��E�roeNٟL;�۫n���{R���P�p�-Xlm�/t�B4W1�(�gc�I�f�Ǭ�jokŅ���'VA��dItuy�+�
�p��J�GЎ�>��=}.ı�qݜyf�i2`��	�l�X�V5kq�}&�mVj4a�a����8���0�]���E��+ALie��5���vͽ������A�ju�=�֍�>��K
4�ᭇZ�;]O��x޹\$�S�δ�}L�C�a�d�x$�p�*e�yp��l
T�*V��;�umZ�[n��I�ܽ�8�������w:���h�q⹳�q":��I�"B��/w ���N9]A��t��|���f�8�ok`νT�$��d�8�P6��+n�&&����6�;��"v�lo.��,�4��W��˸���Dui�6ir�c���|�˙��l����\�C:��V>��=˯�^F�P-W��;=�#q�`�ɣ�$R����rWa�� �Ċ���<;�)���_%o`�l��)ͭ����WBk���J�cꂊ5��Yb���/���e�Hk���u!9�WP�+���K�[7�9��%��E�1Ý�WYQ@C�fUР���\��ګ� N��Xos/��C�����B(�\(>�B����7j\��������8h��]a[����m��v9����,�I»�h=�Ii��[��h�yk���_V*4C�X�LYj��ۄ��# �]m���	�1���++�&\T2C6�0�.�B�iC��%��Fp)J)������&/������B<BǑd]�e�����9��#Ϡ$EA��o*���cM艁�L�X����u~{P�)�8-^��	M�"Wۘp�{WtT]r���h{4��N�ӊ 9�k���EC�J�VDY��ђ�[P��Y��N�j��ЗQ��kS�k�.��Om
�4PW�躺[f��+�.����'�%��Zr�*����of���T��)��ǧ'���}��\f���1�]כF��*�Cu�,���{�`D�tc�����0b����&X����zX��V�ؼ�o^�i�j�|N��{���}�1�S��!�^�ԫ��L�y!��M�v�چ[,�B�Ai{���i��3�,���J�ݸ^�s�����we�'���8������r�*�	i9��-WW���Tz.z�:�'<�C�<;���u\�/C��Ҋ��,�:ꅷG/p�5<5��Q���st�\B��Y��Q����k���n�E9J��8*Q�y薢�QH�JH�7\��t�2���-]ȭ0۞z]4�<�t̵�(�wn�\���j���Yz빻O:����Α�Hң��ji��ܢ�����U(�I��Q��;�.m�1Y�ԋ3;1+X�k��G.9�Q5��s,R�(�05M"�E�=���Z�=s��].'U*�R�Y���P4a�
)��U̲�f�H!Q��RfT]&T�j�!���9��#B���%M3��j�5- ��D�h+K�i�R�*j$��)Cf��B����b�"az"�A@�IHA���3a�D2G'./f��Ў����g3W��iuv�����l�nWWa�ut�mNU�\�*a�cJB�l����<&�N�>�G GGX��w�U��=�"�jHdv���Q��	q����]�7�_C�ON�Sq��ճ�dS<E�ܶ��Om�Ejj!�� H�υ
����M!�6���ZwOS�T��2C�����8�t�ϫ݉B��B#���O=�x��n�~�Z��λ�yC��L���y�☲��H�[��]��GG�y	�f�:3hofwnG���5�J�ր�����
cm7�&�o���uW���qX}���zzs8g5Ϗ�������fD{B:�D9F!��&E�3T��z{"���p�'�{���Ig_�h�>:��>�Fr\P�N�qk�t1�}Fx��8�9QV1���yuY�a��bQ�����6s���B�N�|�0��q8�%[��[f���ȝ�Xn��c�fa��1��g��;]#Ɓ|k�,�.��<���b����"�0��ul�:��.�t9��N�c��z�^m:�[��Ѳ.q��%:s:,6GJ���#�>���uwT���I+�<�ted^���X5(߷D�.mě�f�ѫ��m:��u�'�e�s��z��x��ێ����v�Ǘ�A^(��V�6�B��n��LY�ٶ�U��q�46����p���F묱xg]�S�"���{��xz&���֋����g\2{���{�YD:����ozI�q`�/b��)����vݵ9��k."�!�
���n<�(#֌;����C���fW���R�r/�9����k�R�k����uƜ�CB��8�B����Q+�cW%{�ɡ�v�s;n����E��G���dt*j�Ϧ�퍛�$_\�*�@���5�L>
I�7������5�:��I�]"�I��N�V�n�W���Yn�ـ��{T��`����ڹ�x�g�܇e59��5$g�3e�<��z�~��&�su�𹎸d��܊��Gm�,NҬպ׉+��w���Y�#�_��t�TT��U�,��ѳ�v�$!����ՑP��hT
J��������Ip���4��CjYh��Ó5����R��c6���Y�3�0״�V:�	KN�TV��Љ�)���b�4RC��i:�.���K���K��i/A�g%����NP�u���	j��'vB�F!���8�V㓦��e�+:`��+�;R���:J��vp�A�8-4;w^!��[�Cf�l���l����W[ ���v��	/ymr��s��ݱ{��Aɸ��إ����Z���$ԱW������j�5N��6a�{�x{�e�W:}\��V��K:n:���9o�u.�
�\�����Ka0*����}moG��Nj[�a���{,5#=�N��6t��Ɗ �Y2~V�(��0��l�FK]���5���rp�xŸr��j9��׸��d��$a�)��K.fvm��ՒUV[�������x�^��~_3K���g�a�Rw�J�=������s�G���P�����O�ii-�vN����˹?1Z���mp�< �Y��c�`���v�إ׺��d�P9�>��(ŎDW��܎�cad�_�zʳ+����h�/@�Vh�:��Dm�*�c���n�Wu�ǔf�ʹ_db�T�}_�?��ՙ��̅}�ٮ��FQCʭ��8�+�I������#/��̘�f�ƱX��!�S�67+�f�� ٳY!���>]Ԝ��$=�߶���eDo$�x��LV���r�rO���7�aw���VT������=�7pW�C�_�]���}n�"!�8�g�08�]�S�9@
�+-{F �A"���b|%�����O��շX�6��d��۹�WP�[�ԫm��M�ێ����h&/r7Ҧ�\�[�.,|{jqGfV��3A�k���V�Lf���k��K�P�ܺ%�/��g�m�77��g1����4�;k-�x�x�|�έp��S��cՑP�ׅl$�|N�0��Y�U6sB�g��0��0Q���|~�J���bf]��z�������i�ZpQ��� 㢸@�WKYc��}��1�=�{NF��z�]ՒF��^e3�c��<N�ײpQ\�&Hӣĝ�+�_�䀪���ɓ=c�i�Y~�,QC�;X�<���[}�������87�]l_v6L�B'3�v�K�w��Ӭ�vh��W�L�����S�3�}�!wHӡ:�՘N�J�j �޼���,эd��*y�wk��	��.�� ��X����Df�{���[Y�u��H����5��o�v�rg�D(脛T�>j��J|���ڳnG0�w�F���[!ة[�%Ӝ����[7}LS�:����'� ����ٳ"����.�װ�����^�3Cq=�V�,J}]&�䝊� gPh�](��Z1{,��������� N�=y;ۛ#��N�l�}R�1�y��}U&���'��q�#U��hk����q�OR�k#=��0�s�P��֫V���R�77@�H�a��:l#o0m�AL��,M!�L�@1OuT�J�v�E�����f�R����EW(�8u���,g)�b�h��F������b���Er�ڱS�kI��n��ъ���,ۂ�@������1٬�[w4��jèdv�m9ٌ�Nv9�.�,�b�h?1:�Tî�Ī�*-���F�Uh�l�7lN�q�f�U�[��e^M��H���Bg�F��;;�V+-.����,~�uQ��lӢz���tN����4�� ����m��.J�2��jDpq?_�E���������J����l%��XL8<ဲ8�(B����u��خ��	#��Ze_T�[`)�3(9�BmQV���Gl�Ԃ�"�%p���g�i+&{���J�V�s�nVhg��Z�\��t��vz_H<#ۘj� H��Ȧ���w;��}�z/6)K��%Y7c�QWs#������������h��;F�j�"�q=m�5�n�{7)��i(�(�Gya2T�N�ڡ��/�pރ�ez�fV��|D뙝y�ͧ4/y��N���x�Kd8$�D�\a8D�A�����W�|�EDq�E��mX�]kti�2h�כ��y������F�tKQ�Ey�ul��F=�n|gء�d[C5<�Ӌv��l�w�t�׶��Wמ��J�Wv��j��� ���s� �W��hӸt��Ҳ��?8�[,�T6K�8h�g�����s1�إ45���	��%�ulI�d�vN��Y��_&4�s����]�L�ʎ;i�E�7I�]k2�u���Yά_�<��U_<�Q�yʮ���[	���2`�U�"P��:��Fv���9����J}�n�s{uN�K7�c�}�k�7���r�����t�G�4��㠕o�[f��G��=VK�y*[�!Q�]�քP{,�v�G���y�<�X=N�zM��F��GR��՚+ipM�i�j�rp8���ê��m@g"�(21�O�s��F�����}��s�)��#y�s2�N�D������>�F���	έղ�\�p0ϲ�w��\��*��Jw�W՚;{�Kj�B���;Q�C0�gE�<QK�Їzs;��x��Z|�m��q H���[�P�L����O���ɼRТ��!K���B���$������Kr�sjv�2��(Ø���k-��ݿlޡ>���L�j��0�]z=+�3p� �a�DE��A�x1;p�j�.If���&�N����t�rˮ;�`�w����G�v���x�gs6wr�E����I��p���O;���xmn�<.c��OK��)pn�����FsA����5 �7���O�~����"A]@�?j-�T����׶��J�?s{��Q,
�l�6�'r���ȭ�^E�Ԑ6�%iI��r��s��9�����K�� ��3�}g}]��v��2+9�f�o�رO�a۬�s��63u�S�9Y���χ����s�V��D���� 0~��?
G㦇Bu� �������_�/q�_P�A@˗�`�4����N����8�D�g;�R�P�T���K,D2GlcjY^(t0���+|3{����5�*%��{ٯ6�f0�mw�{NH������Ej���<�&��Q^��Py3��<>��w�b�<�k��?g��f���k�[@.>�A��Ռ"wd.�`#]���x��Ű�����˼W�at��q���VG�N�T;�+Rc����ߊ%��]�L��M��7׻V�j��C��YDt��@ƫ�[@�3�|��ZB�-)�ɟ:t ����4Ī��m��]�W��N����j[6�q�f�r:�����~ `P{ԧ�x�n�ٹ8��W�a? Gq~�vL�����w�o����wdt:�-�k;MYV����c+MBJ�\u:6�}��c[g�Һܜ�/F��۳�#��{*kb�(NWhC���5��cB�V�b�P�0,��j�V�	hu`�}�I.�06J�i#�����9މ�I��{����ٗ��^c��p���ؼ�Y��Sְp@-���o���T���v�
z>��V9�N���W�Q���y�m�"޷�B��t��6b5��̑3���y��D�He�p'����h�`�냧@�%NU��M:㲆��d;�,�sFN�DR�bi7c�I�OFo�>p�*T¹.,S�ٻOU��W�,���_H�A�圢��w��{����ʧ�BE<^��o?gz�^%�����tz����@(�䝘I�+{z��u�*��^�s�Tɕ]������5b��K�u� � ��<V�뎷vG��̫��\��d>M]f��xc���͠_��
�/V�Ц(��<�4���A,27�V�50��˥f�&���kaub�m�b�嶟.寫��Db�XB�2��2|�pu��~&um	��54\��.��Q��e1�{���3�K7~�k$>t;l(�^�d�05rKJd����������=��~mZ䇫R����/mS��&o�T�&��g��pm��
(¹�s�޿����Q�T��)s��_F���V���i�1�;o��W����N��	���L��kNڋD�Ǟg<[n*t�{bĴK"<Y�	�¨b���И�zk���C��lH�|X�mU�$Sa��Z�U��{w�U!z5�N6��O}:5��5ot�[�����x��&�p��]6f�t�Q��®}���%���yK�(խ�&jz�G�X�t�6e�O4&H2�Mܽ��eN��\p.S8Q�]���f�O��  Lgvm��j�����ɟtQRKZ�)���*S�V�6��)��R���7�}4��U璜Qӣ�&W��!�'���\�$��C
��o��a����yf���+�\�J�7^�G�ƟFm-�K]�Jc��B\Ƞۨ�w��D�<N��Z�P>����ϯ<�G��vk� �^�YN3^��mZL�X�Q����U���)y�FĀGn��q������
��ϳy��6�>��u��Ƙ�uHl�^��4�s�|��l�}6ш��E[�[8{S��}
��	�IV%^2mh���ӱ�{���??Y�G�P�|ʎ����}K��W�j����ʜϩʳ�g/}��&���j����'PVl���Ls����6�e�i�*���1���nm�����{ola����+��j�=�r�l��!=�=]γ2��:ʼͨn��M��y����T����=��jv��4�kD���P��f\�`w����l��̾�m)�\�'�۞��F ��oŊ�d���ɓ��[8��ʌ彇���i۳��9gv2�ΨY�+�ݽ�tv��΄|I0��+0Xs�*�����f�=;�Bҩ�p�A݌�ѳQ�{����G���+�v��1�u+�박*[ˌp�\c��������t����f�<؂�ɮBw����x<��w`�������2��s�(7�݊���3Fx8� ���=��|kn�Nm=�}�.�����ʼ�������R��w���j;�v���;��k⢃q�ni�-��#�N뫫�st��v]���j5Q�	�8R���Ҝ��w#��7y��,�;��٧'^�ݧ��2�u��r[��&��l��d�9���Xԩ�紹5��Ul$�����Z)Иb�6bD���5�l�*��������K[W���x�h�p��n5�6�>]Sy�y��7��Iʨ�zbr��Z�o�+��y�G�'�]�C�RV�珑K�|fw w+�{�)c�X�T�����7l���xoE�����tZ�pʙ���z��d3@�WMEvm���>���(Ҝ�i������%�9G/��8$��윜�;6�b�W�+�-bʻ#�Z�u8�������hfA)v�M*�Y���-Q�5�V�i����1��VY�dݔaV���ў�fm�:���2��I����;����5Gl� b�q��^�4,d�v[��	J5���&c��l��u�V��ZA�fA��w�k%�.�K�m����ͅC��hX�η+� h��+�;����zB�wgE�h���F�u)�W7.r��e��]�.�s��I�X�c�p���[��e�u�0t5�6Nw��u�J�W��Шj�v��u1ڽ��Y����S� �O�Z�&^�iz��u���[=yP�P�a��O8���=7J!�^[�vYѾ{%ܽ��t2�nI�@ʷ�ˢ���ܰ���s�;t�\��=S*«Y�Y܎[�H�\�Bl�&�b��X_Zs�A�NSb�Gw���ӱSȎ�u	��#m��O,>�*�r�]^��z�u[�v���Ĝݕ��h�Y���Lӛ�8�<)\q�����}'@�ʙ��0�YP+��L@���p��ٗHְ�(�Y�<���玢z�+��vtM�P�}zݖY�{�Y�1U�l�T�hݡ���@e�q4��~�bB�u9�o+�T��uϬW�oqpFk�`7��H?�K�U����[�����U`�[�bܹ��1�������@� �� ����k��A6��Q�DðD��K0^�ݎ�@Y�&�a�]���ɶ� �T�>�2��2��f�����lN;���ؘ]� �a�NX�f�w#yO6�h[�wN��A�0Ǭ��R�ٖ�d������um�I���Va���2g<�N�*o�so^pD�m	���F@��l��)�r��򽫣�b2[� �w���+wGIWy>H�}��95�Keg4����w*�w0��a��W��^F�o6�-�?p���m��k6Z=OZ�p�\�WU��WF�j�v���VŽV��լIō��K�p�
0=�ni�$5��v]A��R7�,����`��`9!����JL�/.�`g(bMB��R�U�[�+�%G/+7��q�n���NE�X�kp^�y�{]1, �ޛ�W_˿��4X��q�D�N��F�䠝/@/��+���B�r@R�<� S�*T�����J�#�ɣ)hCE_݁:.u\7�&��������H�����?��Jsh�&�IY��>�z&������q�q9]�(�	R�cx�N1������M_D�۽+�6b�s���"N�f(�a��=��xT(�9��Z�5�/�1�m��6'"j�;��_%Nc�t	f���T��w�x���cՅ�e{q��f˦�s]wgen�el��]�h|�j8��_�	����,��q��o�rR�@�ib:�F:��J����^��S����^��U]hF�B�D�I'Q2K����PQ�а���3-
S���ȩA9U��3P���"�&TY�E\N��T:��!�EаJڂ��X�QI&Euad�B�T�iʩR9	��ap�f	�b�$���:�*��u�qN���I���D��+JUD�K2���J*�sJ�MR��\̌B�!C"�憴�mBD�(*�$e��5��Q�DT�I!�f��Ά�`Zd���fE*jr�̃E����'4"(J��S�m*��A�P��$ՙ eҐ�'XUIN��
YUF&hʨ�ӡX��숪�Xey�&AD�%�D��D"�"Ȋ�NZ��e�
g*�,��fE�U&���0�

Y���9(k��QT�31"���"�D��
|:��P��Z��2b�0���8��5ɻ:��2�20�M���t�n�w�D�Y��tLj�Q��r����D�ȸ��� T5u���͊UV����sX��1���Y�S�~��Nb0*�f[�Wo(����g�%��{�VR>��\��8�:�Ûn��S�(���Ҧ�aF��՘�j����\�\҆�q�Z|��<��-���{Q�2t�Xn3��*���Ӻ�M�x-��Z�E�d��x�K��ܛ\��������8c��{�K9ڬ:ٝ�T�GM:\@Z�q�����x��+���ܓ��u]��=Y�n�*7o�S� ���' &=�FK}OHg�Y����SY�S���)oA�Ǻ;��|H�ה�&N��v�L#��p$���^\�i̙5��㪈O��c]��4����$�T/��9���Us�t�ky�Nb�ا�R���Z��6�˽{���rq��yq���=P�����p���nTή���nB�ޝ��R�K��jO�\m��I�Ì<�Ϋ
���Uq���Z���6�Q8��3�+��r3�}�$���]wi���
Z��`ҝ�uՔ⺼�i���u���WX�M�R��R"���ɜ<��b���ͦ��t�1=�$�}L�?�j�i�N����pO�U_UDS<��ێ�YC��T���O]\qKiri�)s�	��w,��]��/v�_8�d�P��
}>;Q�O2n5�w˖�v묡�2,�/�*ءխ>���*��s�[q��D�r���Zb]������Oc姕��r�;���޴C��F��g��s�3a�Tb�f#����'1��b;V\s��͊�����<�n3W��|�����d>#N]Ts�x����mo�o2�R}�ߪ��y���G��w
��	���Gv�oS{�F*;����糧p�����z�.0'�Y�[����77���Q���-�3����Xe��Q{c	r��q;���h��CW��܅t2���On����o�:��w���R�܁Τj1��((T��A��ʦ����sj�������� nR�d�~�v��+�1�0�����6�eޞqIa����E�42=��o�iƟ�^(�׎\"��,��Ђ��(wnj�fs�bx�x�f�Mrb3˖�wS]��43��7�Tkr���Ւ�P�aK�R�V���1��
�j̕ɊV�Y̻�ĳ`[��Q��}VUƦ�ʜ9]�v4�h����gwB�<�ϲ�S�|��'H�6v�����efg,�r���kHf{R���vF��/��.�)��i�w|���I:��2�����ގk1�O�@o���o�ݛ�|�2�-n�'��w�I�I����%�5��]���M���Ȯ�[y�/l�[#$��꫉YJ�B���14��vGƓ꿸���&N(�]�xh�l2q�<���o�����94�k8��:9hö���D^9p�M�v�\��|h���ۍ��Δ`k8)�(�6�k�4�t��+uK�\�]�4��q�kӬڸ����£	����0�ګ���oq��6_�OmZO~?M��Ny�5�����~���=#)m=9*�\6-޽�j�8��;]�Tg+K�����;F��i{<z#���Z��$���K�Ȧ����E���F]b�8�����lP����cܩhЎ�u��J� i[�;c� �]sJ^w:b��_o=]v�C�]̗]ٜ��|���T�ִmI٫�i�g[�J۲}Y3�W3�hٯ���Y���9C��h̊l$\w������;��-vP6�ш�?�+������.�u���]G�u�isάj����0!�)���u�'��/>�����q�q�V�:U����g��NL�K���b��{�z^�;�^u�YJ�/�Vw��17B,�w[�y�'�+hu>*��e_��P��m���l�#�����n�s{֛��W2Xީ����vEqˈ��ㅧ���P�����*r�쮽s*��𞀘@��1�%p��~e�	<�p��P�ن64��ylg^a���Vi���;}�BNoBJ֝�_Vc��iw`6_ZrK{�n�����q�a���HTp�_wg�Ȁ���j�Mp��:m�ʵ]�Ұ���۸��O��՜�U�j5���V�r�B�5�
#��H�ݥg#gU���ޝ1˚�o����J�p!�g/����� $
���b"�;�@��E���Һ���Pi�����V�O{t�C��G��4��_V�P�y�����'����-t���y�Z���|GYέy��okW�5�����d��۪����-�ݭ�+*gn3F���{�zg-���9�.��]DE�%YMer�δo���q-ƻ�X�I]��^������"Q�\ Vd��_]=��<���էS�ڪ�A�TN�l���������{�w+�E�g�y�ر��Oz{��z֞砪�rkǠf^I�p���X;�S��W�~��|A]~��-.ڡ���M�o~�b�T;�g�y��k �X�Wf.5S���/�oS�Khp&����/C���:�+~{_�\�;\v[�j����Ŷ�ݸ���v�%+w��B�x<�����Rsڕ>��v�&�%N8��>b�no�[ۄcg�.{,��)+�(�u���7ծ�������f��%��������;o�^)K��U}kVW��_*���k���L�@�Q94�qjT�`k+)�0	�|�]��B//N����~�e�S���Ӌ��s���̖q���ml�%+�FZx��Gl�n�.���J�v��벻�kyt��4Po�D���Cr���@��z�z�*~JԶX�k�vOsޢ7/�C��v�T�EԸ\H=��G�������¹ԟ
|�`�.�f�����h�]��z�;�#jU��χ���Bb[�|j��g#�/1�{����k�
[�;��	��-���Y�4�>�%�P�NVk\w�>��}�������C��$�/��*gB�u��c^�̗-�8y�oZ����PμO2[sl1���!w;�{�����;}�+`��瑐��Z�!朝M+��]˵=9ݮ��D�[�R�v��+C{=Q#�6n ��W�-��ɗ�t�΂�8�CRo���}��}}��2\Op���(�p�f�<ɡs��@=y��*wD���@�RE'�ƭs��	�֚�27��N���[vu�t�'ժ �l����8١�O��Oڍ��&z�k�\j��=�����Vz>��/AK+#g:{�3}Ԭt39�+��i���ik���_��Y�`:�Y4�n���F�c�,��'����h�Ո�x�g�����v�%�P���T�VV7��tk˷���N%��W�֢�;Y,e"O0��lr���/	�IN��]uv���m!z�W#�P�L\�]\o�n�wPv�{poH��[4:�.�֓:�e$[w��^)���r�F�$����'����� �28�W!f}_UW����;m~��{�0�먕��ð����<���>��t�n���\��Z��R�!��Ő�z����<�E�μs�yZx�]R����Y9�^Ż�coԔ�5^=�k�5�2���]���5mXN�R>ڬ<r�<z�\�p�O\hnL[���o���k{������!Hu�ǹ�R��WFr��N�ҥ}v�U����p�\c��!4��h������j����E�T]��xO��r�KHe��`$󝵫\f��M��U�8�ESӛ������d�w���-��毾C{����E�okN�l}T�n�nw�j���5 t5Q����A>w�S<����t�M��$����.�8�s�=vg�Z�j;�7`�Bi>���/Mo{�\� �	k�z)���gO�s���w�˿�\H
�S���� �6�^�f^zl�&&����w^����°ک�%i὚"]ϴ)���Aw�Wv}�V"%4M�����O$��4-����ӯ�ґZ+(��;r���o�Ť	�lQRm+�N<n�2؈oM�[�,Z�ٌb�ءtL�f�f,+����{�Ң��R�� �m%���W9}�	' �6�]¸���S��&Mf��Yl�t��3Uq�FwcҞ��:ͫI�X�Rhc��-���x�o+��$w�+�-�JX�*oOD�Y�u;=?W�H�׹�m����o4��F	4y�
�U�ԗ1����;F>����A���Ӣ5��ym���14��[�r0�����Y�9�a��زY��k�<+����	є����e���sr�g9��Hax|Bڞ����-��۽�4�'�ۇZ9�y�iB�������ͳ�g�6k���Y��qw��ݢ��o��S}��8�	�ң��Q��`nmCwɷ��٭J,S�;vfJ��Z�"��T9T�g�5��:�"�*�7��X�ov�%�����_&�j�G;<��e�9��_(?F���!�e�	5ݗ������NN��۰i�gx+b���&����,�
����D��d�엽Y;�q<�W���d�������h�m]��>�#�+-b���z;E�[����Y�\�b�GR��[�_!��w{/)򋱙\���<�FP��7��&��9�Y�#qm�s�_UW��<Is���P���ӆ>T��3��>����e%�N�7�"�Nb��U8������nX|/$w���Ga�v<�G�-�T]�i�
RV�67���/�g�9�=vy�������w%2�L��cAn���S���٫\���#�NN��@�=^=L��~pмbӵm)۪����ޓ�Y����q��;�-����C|h�N]�q�,�.�5a��>�q�C�����b=��ώs{�y�f��Oj���uRoO��W�l�*q}ѭ��v'��D��9|k^�����[��#hP�3=l�s�(�̌�<�ѽ�� ��J���@4�|n܁V���5��y7n���{�o�1�y�*��!:��c/*9س�0�Ņ�lҙ����p/�^H�c�P��E������g�Bgv���\�BWM���m�R�t�4D�V�ע����`�B�F����k
j�u��u�����hވ�Q�7w#g8�Mu{���[���}vI�)¦N]�XYS]�Hͤ"�fk�3]\	(O�EY��=�]�C�V�o"���䃵gT���}����u7}��qNDKL�v��P���O��G��e�����4�xA���'��-�b�#V�Xg�q�;����f��T%s���ܓ��iQXo�%z���<�I&��5�k7&����\���Q#��N��\���MlQ�n-k3e�Y��V8톲�}l���;�SܦsB���GJNh�ʓ��/6�y�y������G�oo\5�����^R���N���<��wF�Q�Wv�Y���WX|5%����_Q��e���S�'��Y��t���7(��8aB�zsXy�}k�L���16��͗��Ҹ�w�rݖ���{]�����ϰ�VL��8N�E{%�e���ӛ�&�ķ���gG>��o,�Y|�8kw�N�b����	���������>S�(]�w|�7]����>�g��}A�NQ�g �N�O2j�y窤��`�fÆ��Үu��/h�ei�K�v�6���x�ۍ�w;H�SVN��n+���w�X/��_6J���r�F���4���̼Y����a46�W`j[;X��C�����R����4�T�f���5^�o!�c2a8֋ɂ�D��6o�|m�_`�igf1U<#A�|�u��+ʼ�44W�ѧr��FD�7W]y�"��ut�8\c{�U�sl�+������#O ��q�sp^T�%�aS�r�q-�a�B���Ϟ
�4��eS7̽�sj�X�+M��B2f�:�F�y��Q1�JM5�W^J逢����f�R�-��5�$uC�\J���$��)n�����U,����}��}u;/��Qb�!HYgl��TН/)�[�ТlN\�u�cI�m��m����:�����"'p��m�II��!A�ɬ^�b�<���y��*������=yo馐Ks�n�Z�.��2M��JD���3�	�Օ���=�޵��߶w ����}θc�n��:��D��Aס|��̻N��\�FR�PE¡���!,�>�-���ũV.
���
גؓ��\�	��i��
 ��}�5Y����=b�_B�v�'<��ю�U+�Ի����1Vb���|�i*�ri��W��m��9�Z3��1P�X8�I�6���i�V��I�ﻕ�4cCgIy���*��bebyӤ�`܉=;����.��k3�X������f'�βԺ�S�6�n�X��4�)��F%YYX(��9p���2�z_i�I�V��,f��n�'.��맚�8J��1��I.˩�1N�WM9��N�N ԰�b�gX�w��h/�������F=��v���Հ�3��� В[�SPo-u��y�B��ϻhN��2�R�ũ��`rN1�+yE��]���Z;^^켍Kwƣ���T�W_Yj˨�U�f��Pa޳��@�R r����;{�Y�k鵺)�R���凙��&;2ޛюژ�_t��75��;avhaΧ��ݮ9��; ���z�ov`0�[�]�1�r�5���E���s��]�=[$�5�9��4^�yǥ֭��
��������&�$H݃�.gH y���wb��F�nN�j�l��*�������V-�ש%�1sT
��ُ�65�L�W*
����ή0I���B�,뢭�=\��=���eu��jl�5lݩ��CU�Ú�ޡ�����H:�ň0�Z�X�S�%�Օ�w6A�_ �<w�W,�Ձ��fԳ`�k�g7�#Z���bN����+�(#��$�6�_"j��giIS#w��J���"r*�y_f(fɹ�M��`�S�0K
�T,�g���SزK$f�1�K��;cG��U����@�L�e�f��'Yp�Eemݔ�˻�����k5f�kA�)���,7Z��ong`|q��Ѳ���#aea�OX���m�R��Pf.���z�,��*�6�
zNd�,�Ӳ*��gId��Q��yVF�B�J,�qT��RE�eE�����L���J�6�5+D/t��
��R�J���P�L.��UJ�8�B�:�',�.'H���#A0�H�Y�e����IEh\�)�Y	D�gGG(u5)�M(E �EX+��nd�����%Y�#�E�\v�R�3$L��.Q(�B��T��H�Ddr��4)9e�t"�J�VU�Q4�+*�*���U�$CD�0�֔EYY��D�r!9M#6X-[S�dr��:I*�BDdʢ�(�E
��*��8�AL�g.PPP\Ԛ�>�>�	����� ^ڗs�j�3����VEu(����ܧy�F����a���zOU����s�%�N|��V�n�s��Kh�Y��f[����V~ո��j�9	��Ɯk�5�)�Ze�3w5W��9��������5��Q�i3�������F"��Z��Q\��/'��_eBM�Q��W�{��/�+�sSQ��|�����>��G2�m�����p�1���޶�����zs�V��&��\v���|�U=c��#�%%�/':v 3O�� �OZW�m�<p���r�"q�_>`]��Ls*�,om��M�/�8��5��w��J��+��4�F4�idw^$M5doZA9ÕW�1�\�/����n����le)�χ:��%�`v����\�fe8���]�p��&�:O8���
��wʞT�tZד��d9x��W�]��Uf��\5j1���{`�O�����ӏ���d<ٜ��w1q�%kHf��BO9�Z�\f�{8��<�����`��9C��"�m�w�w"�gMe���mp�#n��5��%N��j��񭻭:��y=�<�T�sǧ*Z��w��th=@΢�mt-�����P�Fj`7ANǓ��0ᲅ�i�[W�3���R"d�/��xO<�]q����r� o��L"����Cx������n4Bs�j������TL7{v{�ƣ�������-嚦:yu�O<�]�Sy�X��<���)�{��gpꣃ�r֓�fe5�ԓܩRWWz���E������p�F���Ό&�]˷.���R���H�9Ľ�ur���Qu|��w\�\aOj�rҹ�-�rn5��IuՒ���q^��\��8�uWP1v�F���3^뢶f�б¢�X�Ӈ�	����3��W"/+�}G�U�4g�55s��zw��T��ӧ��Z�.{3;���M`&�V^��C�]�1�r�����ECW����,����4Y�V��}��r.��,C�!�0����!g��9�;ʿ˴a�3pX�r����!�{�%��JثO�\*��լO�Tu�E��n�J����V���ee�,�αp����,�붌I�1dl$C���s\w]�3� 5c�S,���P�ػrT�]^4B�m�c.¨J
V�D�Ng�7�ܚ��DA�[g&ݕ�AM���]ǈS�]Gu��l/���9s5�V䕶�/�$�j.��j�3��ﾢs{=��{vw�qg�iCW��D�r~�����{h��¾�������|+��w��r�8gK��cM*�P�c�Q��6��M�L�ב�$r1X`���O���l��r`��[�j�p�����|;���^1��b�V�k��͍���1��2v �'`���-���]<^�%��UV.h�4���}���}�H�nC���7ݰ�-�M��%^�!8k��}�|u2;���Ľ5�_zI�uۖ�^Oq��j���cˎX�"�2�l�+^g:�Ǘ֥���!�V�u�J�޵��$�6�3��`�4��}���P������R�����{Ӧ9sW�K��ڕn�u��,	�N�k��֣qVP��UHH�����WRڸ\�փ0�1�9v�֫��M7iŵ�o�K�{�/ju����h�6�=�xi>z�ˣ�eu�AoL_V�"���ίm�"��k���V��s4�cYY��4�� ����ҵ
,N�)�j���s�^����}�R���Z��T��ŮS�#y��Y��[��r��w3�+��Tܒ�Y�����:�BP��w�j-�Sx���Sa7�-wӆ٧`P<nn}}w��uW�^ee{9£��p�׆u#�v�i����^�{�F�-���&��Y���ƅ�F��&z�k�]ol=���4��Q�D��6`�Y�|ۉ�[�ro��yN�j{�ϡU=i�|���EOh�O�#��7�3�✤��߮-�(���1����z뷨8���N���PXb�U��3՜��Kv�_�w>]A���;C]8�>b�G�����a�)�y��-�OW��7sЯ�{cJ��H�cO�ҡ(�K�7"�c.7v;�����E�K'˴uU��|��{5��^�3��'�Pt�]�ܱ=ta
.?uf��ب�L��zs윯�׷2�'#Ʌ���Mnݓ"p��Dh�k�g�9y�"8��4~Ԟ޸ko-1�m���;���H=�c���nx���}�v�9e��^�p4�i�q���o���v|�I�g=�$ʛ�#Ύ5�wK{]I�z��%�y)�+��� �EՓ <�p��K� IO_�7��"-1��.���'뜵<X���S�ǻY�;l�,3��bՈZ��j*�8w,X� �<��W-��<%�mo���cA����>���׽q�W.��DP7��n�z��ѿwT 7�tsY�!�V���r�^�{���)1��;�;�f����r��AodO�^�3k�[ӧ�H�[�x�0�_&��mݣ'���܋r�g��7 (L<譖�*&�l�
��-�}Wy����D���E�i��_Pt��{Y�>�v�*y�Ч�V�}F���gC�̎�x�����H����gS���Hǵ��i���f�듹�e"��c�ҹ��:ͫI�Z�ּC���b�C��!0^�ޝ�x����[�߭'b"�oKejf7��O�k��m�2Vk����w�mP��b�s�b*�s�V���1�eR>�=��ᚲ��QK�rg-o'tX	�f%�^v�zҾ�W����y���J�D
��A.{q���||�1�<��_��u=��xY~����=�����#�V-'3/�,h��y _Vӊ������O7i��]�O�Y�J	kZvhttKJ��n8����5��'uR�x+�&Sj��wJ��=��<r�ѧ\�b�k:�2�����vGF��9r�@Vq�Y�=J��,XTe�ٌ���/=�D#�x	�i�u8�̍�̎�Ӎ����;O�vc;׶0�3�9��-�#�^�&�鲟T~�?-e^��ۆ��o�On��O7.��e�����n��z禽�K�QF�ѩ���e��i���jE���h#rE�r��:�L���/BJ֐�7���_���R�q���J���Ѹ�0����P���;ݱ��-l��dB؟l� �3:nf���j��g��䯺��dV�H~��$w�Iʱ�{�,���e���^�Gok���j%�Ij�B�O34��ٻ�+�:/J����*����TM�q庥4�NH׽���W�A(����*G: �$�َ�U�i���8�wQX�^��rҹ�-�	' �n5ڡut`�� s�.�3f%�,Ve�=s��2��Y�N�j�f�8UeX�ۘk�G���ף��R�Fa��0q$0�����ޕ���	��S�X�vXB��m��5�iHb%�(Z	��l7uqA�u.U�5K�\��4�+�x���>/&�s섧+�X8{%]������7Z��'y3j1�{�1M/��>�at��Rs�щs�;7;��i��y�/ÕU�{V�߆y#Szz/��=kO�oS̰2u�3s|�|o�:�w�z�'������\��j��1wΊ��`��MNX��C���89;\��v��v�0��_4F^Wy1�swS�H�Q����=\p��Z�k��c����-W76�&k����hJ��%�;<^�f��i{ܳz3������(��ӆ�q�nLr���OUvb;(l-鑺�'�j+�+�����+��k1��m(K�YY-�Z���6�3um�飝����{l�!�S;P��i��ą����y�N�8Ds!��|��}���,gB��{`�'c���	�{X������*|���ܷ��6��i�7\%m�8Z~�ӈ%�&z��PBRr��Z�Nv3�:�B*n�_ˎ��"�������krr!�=p��wfx#�6bF��;�1��9
�՚\��ͅ�d@���źZ�k�����P��IhL�
�̀D)� �6m���������
�w�����Gs��.v�Ku���.IR�:@"F�C�����;z�q�Uj�#��1u����H�b[���`��fKܟ�o,�7��iC:҉y�~�j����g�S�B���}[�(���Z1*G���q\�l�ޝ?r�"[��z�{�`�l��wk��j�djSQ���k��
[W�փ��]'��V�N����g�M�2cv-7b"yN��w�s�o'�u'΍��~��& 7_h�^)"���8X�Q��k����v&���jvX����M���~�ƻ.���{d5>���{Oۆ��/�Z��_�lig1�u���v߲AcW0-�d��f��s����/�o5��yڪz�:��i�Ou��U�E���93ݥ�;|�:��`U����/��Q_e�v���g�bU�V)i����"�-��H�u��;q4�����1q�si�=��>�a���'5���Z�0�,��T�!]D�F4�GJ��'Y[ٙ2M'�V�u�S���(���!���V(�\�i�:�GB�_ʇ ��q��P0��O4�	|С�cL�CXY��W����ڷ�y�P��}%D��un�8*R)ы��0�(n��9�ҬmV��+�}S~S2j�[�t�=\�v�rv��l �˚c���Z�}kB��+�����p��d�.b�Ԇߒ�檝����k��R�܁΢G#��-3�7�J��<z𨹬��������_>��}��;Z�������.���\$���8�:��!�Y���p�!|Mv�0�'W1����{����㯬0�D�Ѳ��Zu�̾���V֭q�ܓ�kj�s���y����u|���I?��R[;<���oZ�����׹|���ôS��-�a���x��ZN�7�8R���{ס�r�NtV:o�*s)�U�{�wX3|S3�t 9kY�7 �^�yѰ��B"��ַ����W���Y�����o��Qi���\�k�	��3�5S]������� �qoj�-\��hыI�0��v��"yO�nUwWVT�X^aZ��#�\K�b)=ۈ���k��Y���X�V�9��QR���~[k�<��(���ؐM�;�C15�]:<�<�<z����K��kN�T�xdE��3�7�R��bg]J˵
]>yy'oq���tq8Zf])g�3lEº�<���Δ���B�t��B�)8۬V́Q�}�)ȱ����cK�����;�2*��hg�57���}����C\�=��AZ�:����2??.� h��9�6AߩKKj�촺���̪����.Zi�B_�x���;�	*�O9=�ݭ�^||AߧZZ8קL5���r�)�{�m����;G�$f�(9x��y��g�[�׵{c/W�͒�gWO�{e���g���%G��F'����i��۶�/le)�ذf5�=����f���V8�	�J��[��UƆ�ۆ��M���On �gz�a���jۭ@�L�ʠ�J�cMu;���(����k�����]]�O0^�o9q��Mm��ېd�{Y;0��)�ڸZC4ރ�I�T2*�P���o�g\l��}�/'�� ��'a���%�20sY�oL�)��y��qmٰ�bW*�r�f�6:�Ga��)7���ٕ������1{����b9��ra���ZiݵNcY{���H��V�f��D���&Yj�݆:���w�0��)�T/-m��\�$�y֜�zZÖ�g�H<y�� �n[k�I}��8��.�=]ir�wZ@9*�ھU�Ui��dmt� �*!����嶹�x��0��Ώ(ݰ�j��]�VC}�n�$*I�;3a�7z��wYST곗ιL��W�4e�ǖ�g�Pm�����'�T����,K�n�Ža�HB�5��ʒ�Wܒ�l9�d����r�T\����s�
L+�Σ�*7������hmu��r�e�nqX�f<<P�Whћѻ=���Y�`X��e���������e'�8������a��)]"�
�5�b8s�\l�����IV;���t;T��2��v;��0((�R�X�(�C%m��Tz�nY��oKYXW:f�P1V�Е�0TYƶ�n`��={���,�L�Q�T�[��7�8i;�_	�n�5n���
���:�f���ϱ���p��]�?g-�]k�Z����%)K`Vf��d��gt=n������j�ww�ryY�L���v5�M�mM,]|d�[&�D���Sݾ�q�:`2�y^	����@�rQ�8oYc%�'�X�q���25k0�-o�>�Y�3�Z�ԕ�M��d��ثSi�]Rjŗ�����q��*��;e�.	��H�@K���)ȼ\�R�0V�ܱ�c����W�͑fI ��\L�FLTw,�g7b���� �L���-d+�9�H5Y��}��q�ff-��d�.���{��䦧��_u>߲���s��Z�`�Q�Kum7��Ee�_QS�zi�2�Aڏ[��h�(_R��Ċ�o}�1�uq�CY�y�Rj��A�&b��ݼh��l3^���b��s��:8�'%��>����t��\92&Z���E�t�.��qL�W��{�Y�z�e����������}��˛B�|Q;F�z��"N�u����8����R:aA�+��'$:+�|�X�<�"oW%�7t.�z�r{�@��V�
������4<Mu8dfe��Ƀ0V�!�'�{jq�h����밷�۫S]:���O1aR�)��p�ַf'�-r����T�ќ�J���u�WNh���X��^
dh����tZ$�������r�b�T�^*=�^�{X�[�Y#���t��m	~ش�+��o�~��GU>��z]�`�N��ү�S���+���B��U���u��A�;��Fq叕���R+�7ٱ}�^��4��6Vf+��H,�C����dx��N��J�"���\����w�&V'r�������*ŏn�uv�t���e�B����pi���#��n7�.n�(>/eqݤwPv���Ն%e@����3Wv����7��3MK�O_)h-�%�q�<��m��V^�98�<0�|�����T4�"�,���*��	�Ą���r�D����)�,�.Fl����.�4�TQt�$�f�%X�$fQ���:U��$20�E�Z�#5�L�G*ΖaZ�#b�9g
A5fejQ	!!�)iĨg�a�j�p)�%Z�p�S�IY�ȣ�&�˘�BL��J��5
#�F�R���Åˊ�6Pb�)��"Hĩ$�Ւ�P�����B�U���S��8琝��ʥw�-Y\��TNC�s���T%��s�5d�UTGbZ���@�*�L�M���t�DeEU*��	%T2��v�|��Ծ쾌3Pdva��6c]X]�>�T�8�nqmOI��W3zw;���ouѴݝ�Z�-��ћ�r4 3�+Kj���oW(�%og�7�=��M%�[�w:�¤/����N+6ohG6�^۾�[��R���� ���N��s��K�T�
�B���]�����;8���Wr"q�(ī���z�0��p�i\�o�$����k�6�օ�q��ݽioe���t\V��c��ς�ڪ{�xi?=��)'U����Y,����V��6j;� :����4�A��Q�u헽��}s��|���ϩ��t�3}M�C����0qM��1V�o��KbGgOvN� �%�3vs�s����U<c!>j�0���!|��>���}�l��׎3�[˫�QӔc��x�[����,qm���FnD��^H�ʫ��K���3��wQ!3�����\N>3��.nS)�̸��.,2�y�ص+���U�OOq�"F���*��U�ni��̩��\���,=�f����Z�S�0-Mlb������f5������K�l�9�8M�r��]r�#����v�8�#��g�*糯�/T�sx[�%��Ñ���M���gZ{�����VJ�J>�4�u��t���ˊw5ww�B�k93������>�����\f���ț�o����X��S�����'>r�E��7V{4���.�fl�c1�a��6����9���N�a����'ɝ�2�����[��`�+�ۉ{���<����n@p܀d�G|��ǪDm5���g�j��7oN�������V�q8�nN:C�{+3t��`�wӽ�޹��L�o�\��Y�owJi/�޵��$�6���L՚x	���^��;e�;u��Ϩ��s�A�zt�˚�o���6��+�m�����\U���N5������C΋����\��Z��F:�nsq4�9�]����{������Tz��fF��7�2r��p�m�Ƨv�YY����ѣ*?&�Z5������z��[{\ ��%��vJ$���y��z���o=;���ɞ�Z��[�]�j�f1K�x�:���˷��Ƀ����_��5n޷悻�̵ն@x�l-�tP^�H���7����!��wpS2�m833�eD�)_q6��ͮ�F;�%DU�Av�v��2Z[�u�D��kC:\}��m�.hkA�VE�9R���y�䴺j<���\��Ƀh\�r�QZɍʒ�V_IF.E.r�ȷ}Kg;53���p���ƾ_>#N^9�o��0;Ύ�<��l�Ky9������9�����*���[�������n5�dٻ}n�����a����5�v�5s�*->aiɠ��x�!�˶��ժ7z&�K���=���팥/�+��j1��1�BL��{�fgj�+�6r��2qK���;}�:w��mʬ��o@+_�'j���3�sHOv�j5����u$Η@o/7���\���T��)���yC�65k'{3�d8���i��e�1�=�p��c��-��%لΩή��Y��w����ʁ�'���$���2�7��S���QRQ��ѻo���8i��%�K9���f�y�{�D�hYx�EaiGϼ�Z�nwz���5����7 �AodH�{�~����B&��K��!�[�X�k�͒�{�M��	Jtw��]<�wHMI"λ�5�l�A(���6�v[������U�'���d\�{���7:��nc��3�̔�;�"Z��}���Z��h��
�z��_5:
6��À�c��gV��E�9=�W�����̎t 9kY�)����y�(U
6R�1}��vG�{�k9-�QM�������
��r$&A���X�}ȼ*��ԝH�-�_˖��<m������cF��N�n7p�����s5=�@N?�u�|7�2��_f�?k6�&z�k�]=����ͧ%r�Gk�ZK�9Ƹ�D���U�M��hg���Ԭ��ۆ��*|"w$���\�=|1�ky�����}<A�]ih�����:��v��m�t,&��X�e�.��T����z���w�֖�8�_�LX�+n�;��t� Ƶ��<�V���9nϵs5=�^B�����v��L�/��u�������*��l�Qm���g�{c~��!#
�cW{��f�N��Lw���r�-9:]]�Epo-6����c�lf�������˻��ʦ�H)@�ǜ�`q��A�{�zY�Z@Z��L�d��Ox�Ch� u������o�gV3x����-��S��5L�q�]��/�ޝ�A9�YmP�ܚɸ��VsZ=��v�r���V���Rw+y�v���X���i�s:�Ž���D��5�靡�%r:k��u�G�Q����p�FR�]�U�Woc��9זhm�cy@)nL��'K��&0$��}M�*�@ˇ�i���MoA���o;���{M@p�A���� '��ױorY�S��k��q�{}�f�%�<;�P�nX}�{�ߺ�v���2��0a@p%�Lӽ�b+���,�psk��<�W.��wrф��	�d������)��r8���Yx�T�X�_�T���N��]��p˗�+�{��'e�=�wnoW�	[;�����@���\��Ar���,�|h�Iȧ˸�}KI� ���iu�L���;�ܥۻI�,קQ���	Xz�w=}�W��]<�
�c6:�x����9�E<ˎ+�c�
�M	샘5Yy�X�з�m��S녮u��Ʋ5�w�S�7���-�#�
56����v���!!��sЖ��y*"�x�{�>�4�
5[�!�uK�ѫ�����ru�LS6ҬQBK���\edX(G�n����䲭�g�_kn�&޳�iTznh�����os���Dg��SF��GxZʜD7A�k@�ܾ�:�7}Ao�v�~�<�U<c暡~7��,�9̯F�����8K}I�k~���0�5x��3·���k��S�CkJ:/;q���H/w.�|���s���cuJ���q�<���e=��������S�Fy{��X>��-�飍[�Q��*��YW����yFY��X���ik~���8��������ןFD�N�V�ɍ���I�����@e�W}�8��4{�5e�b���-0�{`�'`k'cɄkTX��v��;؟�/;������	<�p�ㅝo�*H��ʟzdF�,���B��}��u������E��}�*�jqxܗ���KW��罽�#���g۳��{&4&��Y��wK����c��.���ٶaW���٨	/����h�NȁϨ�{�mwvi����G������=�$��Eҵ��p���zN����^�P}H�����NVoS�/+-ܹ{EI��K�m�2�[�9v��؃�P�;m=�dsk&��^=�O*����ehaΉ����7�c_�T�Cg;��H����������)�`gp,k�sz=ܪ�&x�i�`8hF��V���@�yՔ�WD.Mh��8lc�w�:���>�4~I9w�cG"k��}!i�w_]-l�V3.9��d}pz��7�E���Iq��?Bn5��β'��M�T��e㼗z���Q�.��_m�\�7����N���u�liwU�ž�oA���7չG��;~��I7�����l�L���������k�W"t�a��wz�뭴��nس�0�U9������`�b.�z�oqc���+���Q\��:��jC{A�}io���ۑk5y�(���"<R��;b)Lf�=}�q���n������*_�'U������pU)�wJ����̍�̮x���e�u�;X{AS;C��5J�˶����ņ�qƕ+���+QW����WϷ����s�Pn�Ϥl�cE`
�w����� :�jf����e��l[�}u��3<ZY�v�aɍ�WS>줾�x��Z���횛�f��:��7/;w�9E��H<�A��9Jap(�R��D��r�#+���Oq�ϯ�Gs�-M��5Cӫ�U̗�D���|��~e�?jOo\5���|�t̠��%�a�YȪ�Tw\I��_s��DOsBJ��v��!��G��,$��9~�����k^����ɻ53��j:�2v ~݀����#�ov��K�✓ܬe5�߫q�����ޘ�ݓ�st��<�K'd{G�+��p��fђ(7�{����^�Go{��h�i�=L��B<������(�l�zά�-�"Y�`ժ|ym.MC�:a.tb}.���1�*@Wܧo]��}]=M�N����B�B/�x��a�.Z~\��6�I�)�֍+c�Re�l��I��������-���q��ޞˈ�zb5�V�<�íN�E��ڵ\����9º���x�lM�?Nb"�e��t��jgp��QF$Ĝ퓖��hvlH�yϒ}C:2��1Na�"s�U���Er��d�߳�A��PV���ՠjFQ:/	7:>���]����b�|���).\���M�{J+Á�s*�V ���=�;���7l�H��X����wa|e;�q���
��.L_1.���n��+��Mt:Vo'|(te�]\mr@�i�k`<c��;�wmس�su/�X#�iـ���ʆثc��ji����[�ò{���\�Ot��^B���<���;p�CIf�gs;�B�U�\5q��18ܘ�܇i��۷���Nb���$TʞW�H״diA�����ۆ�o��8=�D�J��O���r���z��g�v�(��5���(����b�d����ko��{�2�?&O��e)� �{x������>�۠�	t	G�0�W,}���8�6{���p��2���'`?v�ax��E�=�G�L
v��=$��o�>7�r��/��a�3c�����^�O2���R���O˰���^��%�9�[ɥr�[�y�a��HA��2�)�R����U���B�4�U�KuJi�N�\��]˷/U5�aaѕv#K�On��sY�Fʣ�)��djH��	[}�@E�w^^?��ǲ����\G���{���2�+S*�C�_q
��u�D��η:����u-�mn��h���)໐!���=�t���9y��W1fgN����U�y�,�ϢCG�뫥��
[W��r��Y�8��]-���&ѐ�5۸�^N��Y��F����.��˩�22T�-�t��H�}�k�-��6�~���A�3�`��G%���Y��f6�a1�]K�(�v�Mz�vCu��������f|Ug�W\G�̘��e��i��FR���j.�N�L��{�y��;��h`5�F.�x\Fu��c4}��5����&+?�^��+�댙��T�W��f�_r7ʗ��ꭜ3����D卜�YaV@�s'�^Y��ez�#Ʊ��~w	n���*g۽?����a��V��v�a��#�y�৏��u3��t�U�;�����A�9~c�7��u���=�/������
�Gga�a��"��W<j�F�[3-��޻�y���Q�<#o�������}�^Cq��|�=v���VzJ�4��X`"��?
F��Dx��G��7^�<i�rҠ�W��z��vC>ћ�n�̽	��O]+�I9�)8�B�X�9�Ί1wr�),q�opDY[�mV�r2�����V��`�y�{���64f��ňM�կ�t]Ýhp�N��R�=��:ț�uEV�R���4mrھ�V��оtH��������5��t�f*t�u��7Xs"Wf�l]$���"�� ʽB�Vk��%���pG�]+���ӐǛt��N�;�Ƶ�bn+�R%��[��U�|��T���G������rE9v;{[��w�����ۋj��}Ϝ����	�u��ı�6vaz�B�%���4��hjZ'� v�0�=@P�7y=h�+1�18,�j��`�7D2Pr���d�K_)���w�e:��\Q�(m�ώ����)G0�T�ԇ|-��C�6~���,8U��9�����qQ$�L{�>ʾM����j��[�����\G7n����d��gv�_�Ӽ[�0�x�Ԑ6/N�ܢ�5�blX�KfWw_~�Y����ۛRJ{��e*J�'-�qi�a.�mΉYՃ.�"I�RP�ޠA%���Cu�)���je(�H*��=сJJ�boQ;�!n�q�\��[���㻴���qk���pQy�V�i���[�u��Fؕ�e��]�� _(Y�8qQt�˨���B��u���]|-_>i OR�*��G��bWo'�f�-Qx�y�h�{�;���K\�T�'Pj�C�N��é�2Q�b�aY��Y�[��x*]��+��7�A�w\�PAXrQ��.uˇb2¬hA��w�r����-Y�\��\D�:J ۢ!ˌ�]fbW:WM(�oS����3�u�z����iKKhuG6�s��Z�M�	yO+�����vo
:���N4aMe��m�w@;8���[�3�G@n*�H�!1ȸs�ʤl�%�:iv�įozT���`n�/aQץ��
uX��Ф�fr��!ӑ�{(��d,r�`���6���x�����+o0{Q��;:qR��K��f���	����5�wʣޮ:�5%�����J�ٯ�뤗b��bb�QEc��H���f�ࢭeJ��v*巛�E���8���,[�hۆ��Mt�C)S�ښ/�r�Tk�t�.�jE9EVbu���4�kZ^N��:gu�=T�p4_Kچ�w_\�/�Իk�ތy2Y}\��"���{�/���/�b�7����Ǹ�R�1�+1Mf��4\[.��_'/n!���5�2�ik]�f��ԧ<F*�f�H��`+�ֱ���8W�W'^�p�Ϸe�Z�u�;�:o�va�Nށz#�3���8D^Դ�̒�f�Ǘ�[���j�깡@{���)Yƞ���a��ι}k���1\=h��ߤ�sFv��P.�v^Q�[F��R�·�f�. �wЅ�����s��ܙ��]Č���9�����9�ь%T1�=Sַ
2ͧ��=�3���^�������=�ޑ�8Xt�R�()�9�M3��%���	͗U�,�$!�Et���
���9�r��t&�圡;.	5X�iїaT%F,-hjr�B���e��I\�i#"�����[e2(쨙WdL���r��*8�M�8VeP������,�L�J�S8QQ˴�dTX�PU�9]��iEE˺��A@Z�XP��fQeAT')�I�
�E��UTwP����.ʈ.�J�V��WYTE�2��$*
�&�Hl!0�+Z��EU�^�\;��]`���&�"ePP�Q�#��)VE�r����S�g(�=Ĉ�ɎE�Q�Nvs�FHD'B��a�J@ �AE�kY�b/[Y��ƈ���qm�톶���z�R�m˼�4@�o���9���w1[�nΫ5{����ͱ��Tr�x�����Vy�8��x_��pn"��h^��?�}R�g��S	ȹf�Έ���<�~��Q鞯@�5Y�!��|��!���I����!z��87ި����K��y�w��j�ڭq�j��q
�����wл��u�1|�t���*r)�ۜο0/�:P8��o�)f�ߵΠXt�+�!Arj��*)x�-]4=����r�=;��^�>œ׾[�gx�ߺ}#�=��g�GƉ�t�A3��ϊ��Tۑ1������lq�:�z��W��;��ܳE,��z=ˁ����6E�l�G�������g&��ԃ�IO��\�M�{9�mya���Y� ��z׼8��z����{����ˠ���'�rx{*���^��®����;�����tb�W�{�.�[5�:}��ܫ�;M�|��Ќ}���9W�d���?O++�;͙�-�A���ç@Qa�zv�|*��'a[(�����k#Ӑ��g�~~%x<~^<���<���}�U��J���BXk�p`nب~�|%'na��ok�x�����;�O��L�yz�.z�f�U��.2)���n��v��ج�K����9K\t�k�oz� lml+\���t�Q��R��u�����+�od�*�oV,:j����������HT�`Ļ��Q��XZ/'N�*oCn� �3.>���vc��Z�jsz\�d���m���z��쮓��Z/��!��F-'�|3>s]��g W^�����C�3>�3���9��P���O�d;G������V�J������Ek�=ya�x�빣�o��b��B!D��y��c���߽��^(�uU�����7��C؏]{t�.�ڱt�r-��&�¸�%s�	�.3r󇏴f����27����w�|��TI�¸2�׮ǎ�[|�xȡ����bZ��n�9�ׅ���7��zs�/�}��c��{�}N����JYx��m�~��^���T	��
s1)z�s��u����#��Rf��y^ϱ.�鱧�L��q���_a�GŇ﹙�����
�n���H��_E6x���a���c3J�(Ez��WT�3f���Mz�9a�����_��	���*�*q3-���&�x�:��f���NsV��ʚ���F����Rc�!?[c�T��{�~g&K�b���@l,[s��l�����i��~�+��(���T�.#�Ɏm� Ǡ{�g}���:.��w�����*�9���۲���3�fj���ͳ1������u�(�M#����y�uJ��I�S؅z��������l��鳷���I
�Mo�˼4s�!�=�d�<i]c�C��^k��5�C�"���-r�h�f��\!jR�����}Ϸy�G�JV+�`���|T�(k�q�yݑ߬P����=�7�Л����n�&����C����p
0C��5ˎ�G[+��������\���	�f�LY����{*�zY��j&k���'^�q����@��"��t"�H������w�~�{ҍ�C�)tX�\�;�hd>�^c���ܣ'��7@drY��d�Qs�����M;�E�m1����=��|�3;�Gҙ'����vz{#���мT�h۬�!߲�e�����m1�:�2w�=�]��{�1�k�'����w^c��^w	b9��VP�/}�F��6׎��+�T|4?U9�T���Y�����gγ��e���#�/��7�O�g޵q�c%TՌ���wO9]�<5�w�$q�g����Y>"㭚b�xܼ�>�7�g��ӯ�i� �����Y�:�t_�-��a�/���f�E��}\�S�o.LΝ�K��g{��a�\�7�֨&����^������n}�>��1 �P�jG�/��B�`V�P��,V���N����=�F3���o��[�.k�آ�E�54%ر��Ύ Ү�)�̨���+���_W��%��k�Tm����ةp#:�WE�\��׮�q]�d�O���%q<�R���6�N��k(��Sޮ�5�v��޳�hmQԵ�3r��a/�Z=^���^�hϗ�����3;��ʄ�d�W,*s3>T�7ʹ�Y���ۼ�+9��9�b���c��!z��*�޴�Y�?ml����X�
�BT�G��01�:{�r0���5\ʑ|+�9�#P{�Q�?[b0{:��>�w�ɜ.�f����-�/=���^�*t}SB;�<DՖ|���l��9�r�=&��C��v<�m��{�/T,[uoP�c"]:���^Ϣi`����3�_��s�z��K�ʍ��Fx�ݾ5]���|g�#�U~�zg���&f��jAT�����a�Z��u������s��,����9>�w��"�-��6�~��,�'^���푒�X�0�����ղ|+1�ؼO�>V=��C�7�O�2|��TϏS�v���Y�ެ��NF������x�tb�W��C���_�����.��y֮=��h�~�����+o�����{���E���ǧ�yФ=	�ѷ�W��.�]�9cg |d�3���3)���Y�:��^�!�+��R:��ܡ��k��Ql�r�1x���;C%O�kb�|�d,�\;{>�;g}��΂̴�i�6�x�vSw2)oq���0����(����:l�\w%�⏄'�n�Qn�¬EB�0�v��^�N�����v�/�O��[y�&�hl�褕�bZ��3ѹ�G< �[Xg��O���+O	[?9�/ ?{��J��H�ه�Z���:�|�cԣ{�My��m�xvG�����`�a�V*�.o�����}��_����Z���g��ʫ��Dp�X��q^������z�O����]������`R0���&�S뗑y�]\RoH^��\WW�j}^���T�{s��̾�ϧ�����`#� *�>�'�*,��|�9�g�O����>cӐ��xx���n��!z�����Ky�bu�a�'YU���G�;qᚋ�o\��=�R��H��M�9����I��޴�`y�\5��GG$�I����g��'|��
��>�U
�2�����P��g�n�]*�+R�)�ۛ����#L�3����ξ;f�����ف��2�QB��5��K��h{T0}>�dЌ��'\�o��n�$��#�T����p{���aצ�U#S-S�H�^�Q�a}~#;�c7��h�!��T�➏B��Џ������TH���d��fw��K�*`t����-~�{�%~�����<F���gcl�R�R=�F�m���n��4���`gxs�.��*c��!]F��GyQ[Sǈ���Ol�z��z�^�<���Z{z����pmJ��h]�N�;W�^�_��4^*�+y��� �4��2��V!��X�4��c�V�{�� ��%�·?9=�c�C��	�}Ng�<���yݑx�f]����<����T8�Lw!o�d_<���_!���)w;Y=Ɨ���!���/����'�#!�����츮�#�ӂ�{��y�}���1�+����r�v�]�D��.���.}q�k#�꽷��9�R|�zhs�̷uo3��]�{�^�f���+�k�W%�^
} �b��q`R���������x���WL]�9{���t`�d��;r3�u��~7=ìt�{hR���P�F�[w�j[�������{5u�R���Lfzg���L�����wKޡ�����h����ά���]0<��xޛ邆Eg��{�վ6}���C��
z�}���^:^���q���~�ʳ�aue�����z}7��3s:�x�*� =�\j�i�,&�|��Q<}�7�>ћ����f=�a��˙4�T��ay�h�����ę<���?
S5!���ۿN>�^��7��zr;���Of�v	���bQ��ٿJ��w�U��n�D��(�Ao�{��c��O�>���6iMq�C��p/){�z�%,L�w��ĨZ�{�R�!��3W1��V#�Q��Z�E��J�޵ǒfv�uy��Z9P�a��9Y2��gݥӫ��{�5�»�ovq�¶�������R u�c���Z�z9�6��3Czg�f��lc4�"�L�B�wgTi����{>����lGxΎ���ŘWt0�ĤEx�l��K���`��Y�����_�SW7�����NS�3���ǧ�����\R *{��Blq�A�mW�o�d�Q�Ƿ��G���{��s���O��ȁ�#�>��.EǙɓ�b�ʘ�'W��{33cѫ<�$�yV{4JMb*O�Y�F|�?�rc�W�-����χ�fw��L�:��2}�L��w����i���DUt��U�k<{��m��/����{�숸��b���f��vǪ�c�����Wv}�=~�rßX�3��T>��`spyu��t������7.u�z�)~��io�`��R,�3�J5���L�_�9&Lk�X.40<br�������H���p���sU�]�:��b��N}�O�}�����e�w�h\��s!Uߋ����7��aO���N�5����M�����4�2x��yJ�d�w���/:ϼ���v��z�� �`���U㖽y���=x�GI����`��I�^W�Gx0.ט��p�B9¢#bO[~�:k�����W�x�X�#�,껗�ϖ���i�@u�U<k����ݏ���#X7���RJ4�"�B�u��أZ�-�w���V���o���rͪM]m�Yb�|p�}]]+s0b�3K�������� ����5X�	[Y���l�/�c��R��~����VR�15]*��>�Q}lϝp�L��>�p�~��ëS��R����p���ؕ�F�V^���^�Xd�A�W΁Z|&��E���0��e��x�D�ݫ��UZ1M{J�K�uT9���9�a�_1��4��a���f|��}�J>��f�ط���L�\�'ud�)3��w���Ǿ3/��ϸ�:| �*M��V͟�w�;�v3})R�gGz��B����t��F/i�~���q�Bp�%ʸ�aS�����t�	��3\�f�{�_n��L���#�{��/}�=q^��%��Z��{�NQb�'��g�yۇ�s����*�Hc��1К��="�4=;���[�&9?�8������V��DW�ة��N|�}�0�����r=�iA�#Ŕ��A��?%k��o�
Y{�'o�䭑8,.[�M�������e���EĺuT ��5P�X����F�OAP�s݆R?T�Ub��Ύ��"����L�g«���/�$Ƿ�*\r[>�v�}r$d�7f�{|bK���L��Vʼn��k�x��
 �-_(�o�B�[��R��b��w�N�'m3[�dR�s{F��jcI��3������1�bh�N�^1(��W��
�a(�M]����W�v���N�hsGTU:ޔ0�e,�ˑdj��8�Q�^�8�;>���o�HO|fY�~�Mp��dƼ5 �0=��*���P��6�Օ�oH�_X�Fz(�ތ�t����;M�OBd����ϊ��a���Y�ެ��ừ(��٘N^�^7���8{�ճ띭������4b�~��^��&9��1Y���C(2w;������Ӽ*�@`��Np���wNX���V|6��/+�̺� �KU'�8�x;�k˰�v��F�p����g�֪�_%�AGjf����aOI?u���x{�t�O���O�U�9�V�G�D�j*G��_�3JwG<Fv�qV*�.o���{>�����z�kZ+����L��Ou�����X��W�7>~>�,�]���EY�]uHm� �~��=�3��ޙj��|^+6=Ю�!�,ˊ�v���!������ۑ����ߙ��}VzUȴ�����U����t��ۏ����2b%x��~S�5���0Cg�<�S��g��:����D.���=��
�sQ�g*���H�p&W��M}��s��y}JJ���HD��Z+�]2*7���(4̹\����P�t�b�ϏG��É��J�/Mc���ށf�W�`8��f�b����I�u�c��ӱX�%�*�O"Ԣ,��é�GXg���Oe/ �h	�[Z^-��]��2&5��S����b�R�K�IcF%��yf�ߥ�x���x�*P�e"<D�o�O^c��>V�N{�N�d���7��q>o��~>����~f�a
z�MCw\TR�DZ�h{�S7��9��U[�[uN����.�=7�nr�P��d��<2f��u!��:�;�v�z�X�����K����DP���Lq�j��_y�����.g�=�L�y3�O�jAT��7r��.�̀�p����5U��z�$�Y�����c���\/�����"��ˠ���'�r�v���qt�{�e5�]�
��K��+�U��Z��pu;?@{o.B~�B1��������b_�YM{�+;��Ez)u] �V��f"r����=Q3,6����͞?V�;��O��7�A��]�X�ؑv���)��F���+�k�튇����G��H�ZG�ĸT�������pk��\��3����^>��gX��3�:;+��{h����1��U��i����(ᣑ�k��fe��>�����,��P~���v�O;��ά��t���:;�g�G��ǀuu�Ժ]�pޘ8Vd���Ԋ"E�Gn2i�Ldww���ńX��-ؕnZ�j�].^.�9���N��X�ƿ�=�ʵRK��]!j��h��'w�����l�N:��rr=�.�<J����;�S��[�K���\���F:˨��j�w���:��u��V��ڡV�.��2�mMΊ�ؑ���tg4����45`nα�f�Wo]������6�h-��ZŔf`��ч(�.ָo��\�Z�󭥦7��U�
����B�k��Ӈ�\��wi�l����nƼ��S����Ny�q���",��AF��ihbS4]�î��g�b_�0p$�.�g�Z�R,�&c4.��5{(f-��} ʷ][���E���GD��/*a_�E��e��9$���!M�ł�Q�F�i�]�����;��u.������|�Fѻ�gc@< VS0���hUܛ�k��0슞c�ϻ�n�t�nT,n��~u��7�Im��z���z��
�2�⫓���O*驴mrJ����7*�{$���V�t���hOr�X#�����\�q�d�ɂ�]Lv�[>Axn�HNA)/��p
 ���b>��Ⲑ	Rvf���qG��f���̮sI���`yX�0W] q*,�	;&�[`�m�l��m�*�qd�uz�95�]�N��U�n�ۂ�:h6�f�](�4�Mڪ�t7�8vQ��F�t�8+\Ou��z:�@�eC�4gY�J�w��b9��vm���� v4�Ҳ�����6eC�MVY��h]�Mf�χQ�g7��R��"M��s$�h�T��eo&��+t�}H���CD�خ����&�J�Y|�=q�D�sn��N=��mysΥW[��Ԗ��]q��PT�V6iR{@�vՙP�M�1[2�]�P�qi�����hl����:�[�_^g5�4p�m�=l�tj�C��ӡ��md�}��y�W���V�[�ő&���@¯�k��XEn��3s ��:��V�E�j_V�h������v�3��.�o&#ա;i*��+d�+-��5V�k�]���m�vo%,j�IJ�j����@c.κ)4�5D������U��9m��jb�7����&�wҚ9Y}v*�8;���OH���i2m��I�P��Rw7�櫮L +p�t�yA.�$r�)5>�s2�:�/qX��T�)�̕"(-n��ڔr������R6���.�@~�Zgd���h��[ �j������:���C���q�z�EYxܻ�emv)�u}�r�/c�<��U�rP$��5{�%�7�f��U4�u7;c�yN���a���봾�5�ʱ�N�k��-�p��xC��z�G:�w�ήzgd@;"Ѯ�������w8fg-!SIV;OWp���N�X���s��莺�Z1�z���ǒ��(�ͺ�-���Vz����Xmw+ܚ�֕�m�@�������]���cw1t�}M�� �	�����9r�$���BHC�`��ál��&BIE�PE��(�#���r�Q�]��
�UEEG�KU*����+��+�l�"*�����,(������)\�+�v�*�Z��	�MH���((�A+ΔQ3��t��̨.\���Jdp�Z�ZQ���n�N�դ蜈����*
�y�����-B1�t�p��*��AV�F�zйT�Jue�*" �䖧j)�\�
��Tw6y[(���yzma�W�w9xI*�(�D�**&zh�
9
�Z!U�E2����D\����^�Pnq&\s
�g��B9PD:�	2!��p�p��U�j;����rC�4��z����;�{�k)�TEy9�TW

aH�J����.ʪ�N	�s�zG�	��s���B����I%r��qDIT� ���Y�p�[)US�ND�[[�Cn�ruk��������-Ӿe;�v�p,+(��2}�i�#���q��T'3�.�Rv�F?�g����t��D���޻��h���c�����\{�x���VzUWt�|=��V̷��]��z�K3Hǯ��r���z��|<}�|'��3���d���_]d�����kj�ym�,�A܋���;`S�����[s𿽱��~��}���4	T�D����c��>]��euT6=��C��W­��jRD��Lx���46#���jz|�kNEߓ�R\���n��dv#�������::���f��A�ĥ�+�EDSg�4�A��N}�S������>��`�!>�9�;s>��P�zx�ޡ8|}qEUN�$L�3�K��e}��x��sVg��t��m� �a�žRc�?[c {�H����\y��0�حK֧s�x^��WZ�N��z���%9{�I�V[F|�?'5�ڿo���x�﷤=��fF��{����ܟ�A����^���J��L�N~�r/�^�Q�;� {��닃�Ew�Z��5h�CةD����c��P`#9P��9�˯����_�����n2�[�!7A�lܗu3��˞�����I��y%�j�f�w��8�複Q��Y��x+_Tz.�lc/�c%��.��s�3���_,	cU{��m�&!�T��"�_b�q�����t:v��f1$n��1]գ��ggt�ov����EDJ3��t9v�/���n��ߢ|k�������$Ɉ׆�_����n�wG׺:=��"oh��݆yq����r�p�s����W��5�,T��59m07lT/ _��ѕsk��=�A+�\�U��9��Q��0��!s3's��8�>�Uk��Y�g������VP�GIJ6�(+V�o_����U�#C�Uv	��8N�������~��^Ǯ��^f;�7V�8�ou��X�H��{�eM�n�u^�1��t�����GS�K��q;���~�=&�n�ש(����\� ��;�S0ԝ��s�`�,u�V+���'�\u�L[���9���ZЬ�xa]���ՋT�D�C���?x/cھ| ��H_���ϕ9Ϻ�G�y/h`�]��7WI���EMW����.L�5�_NGz+�n}�3/�����E_�;���C�"M�Rj���V����t=
��x��+��>�\U�7~ы�|��T�h^T'%ʉ!S�M�*����U���7=��3;U�u3QY�)��~`�!q��*��Hg��x.�Ǥ\{�Ngs�_35c�T!z��M�Qe��F���Cc��u!�ao���EȠ�3�P�q�@/�l�{�Q����S�1,���.,������^t5��E<�,�*Yk�rd�]}F�����73it�A�!B�/qMm���3t��%rMgz&t�r�g���ٖ�[c`:���p���u��/��Lu�	���=�~���5Cʴ�>΄�p[��^93�|*s�T���n:��|��]=��>��r�=��pw\;ڽ�3���Izǆ|=Y�=��D�uT�: ��K/��dm��Fu�Q��~��yg�w�H�>��ٛm�
�xzg|��L�T�Rr[ �ک}r'Z��;��.��w�s٫���]{Îo_������-��7��(ɍxjA�i����a¦��gĒ�\���wG׺1]y!�r�p�����&O��}�3�>�a���Y��|nzDj8v�vg���z��Azt�ez]��l��_��i���\{����?R�p9���j�ֳqo������~9��X-~��n�ӆV˺',l�(�
���N/,�̫�C�o&�����tk�����;����rG8Fz�jv�S�?H�
n#���d�ϙH LMײ�^����w(;���r'�k����;�=�ڨ��5��˅C�`W+�M���j<f@�)5q!�n൳�wo<�{6	lS'�.����;8�o�y��{	�ퟯЊ��:��iA�wy�|kGZR$qfě\�"kj$5Y�F�z�w9ٲ5�.�ɭ�&C�p��N�e�9r1��urɧ���R�H�yCc�:́s�X0����W����ٙk'�w0�4{�&��{�q��|��j}=�VzO˰�԰��h��ԗ?b�u{��葕ѷE��󻇈x�F}���������}=�g�Ft6пm{�y�]l=�����%����T����1���>������X�O��2��sӋK��{���¾�]@�+�!�O9G8􍐐S�.����I��z��y/�~E<����}���c�ΧG_��<K~U	��%��#P��������ױkVG:���zAv���W^�S�k���οK��ΠXT�)�PC�!�5�@^�#�ϰ�x�r4X�Ns�k�eMy�[��0��ޱ;7�޷9����>���̪F�t ='�<�	�90KR��I�C+��3у�dy]/8����o��tBl�G����&rk�hH�];�^ܮ�����P>ZŇY&�u��1�(}K�?a�{Ȓ=��.��x����i�� /�}�Iom��S�7*��u�|.��ϫ%q�p����sG�z5�\<�O�hE�wf��觵��m����m�����d�W�DeM��Z��}��/QY�k']7�p@�cmY��&����q�k��Ǜ^ATU�ki����ѹǙ��f5�>8�U�6w%1��1cn�Z�����p}Z�a��'j��y2�$��=p���s��5wY�W�3���rh��T?���ꅪ�BՎ��xl�P��ϻ2:b{�\����RJ,z.}��zv=�W��#s]zrax�z��z�g�)���ǩ���]9�����ny_���~:�d?���:{���,��~�~��m_V�q���WMU��>��^�Bh9�Q:}3'���"���x�<��Od<=9��mv��y������3ܫ�ϾX��}����Ka���	��{��\{�g�\mV�{��f~�]t�>��s�G�Q'Z_���ؒ���.;���>��=S��E(��U�����ݏj���j�p�A��C��p)�ԏ 犯J�TÇlܘ���zWA���ױ��j�~3������Ko���D
�!����l@�3���#��t�{�!����}y�{��3U��#������g>OO�[�zN-�} Ҏ�#h�-R��>
>!}<�Q=�{�U׎�u,�Y]�`{�uK�۾9��W�"�]ט�?��ޡ8|L ���ǿ�%*���ʎ���en�Hk�qT/�#Y���;���S����˩�3>���x�v���Y9U�.���)7tV��B��u.�+u�O���&):]�.�GC)��8����	�U��:�crW������k���:ڲ{+z7�U�:�-�\����"��7Ƽ�݆r�I���m�������.EǙɖ�7�׌���ij����W��eM}�!p6�՗���V[-��ܤ�_ɫ����)s#�ؼ�M���^bN���;�9�����䐕��P"=s�r-V�\��>�s��mxǱG�&����<�ֺ�}�2��G�%�.=��N��GOҡ'�-���@�ք�3r�߆�>�7;�-y���7~ħ���N{]�J��L<�J5�~&k�#�$λ���E�}�5�!���[��)%���?���Z��_�a���o[���l�S��C�J����{(Ʌ�59���j��e�Mdו���F.G��<wr�	�������K��o��?^u�j3�l��裰�,����gi��ApR0g���X��d��x'����~���^=u�uz�I���ڹ�9��s��X8��9�~�`d��6�����q�}b:�O�/��fU���@&:=�s�~:�u(�����L�xE_�5"�j�J���3��Eps}d��.�� z�P�=�z䁀 �:�7����O'��3����b���T��LO�w�k��9��-�K&��,�m� }�o.�z��B�0�۶lț���t�3{rT[��|�L�]v�YӇ�G�oV�%r��u���Z��O^�V�涕�q"w�9r��N��9��>�~�xs�Y����,n\ƪ�&��
���Q��Y�"a��ϕw���*��W#�3����E{�w�2���z=WP�� ��1�ȹ��U��wם��dO�{K�ۯ1����W��{�*⛿h�����3/��{�%�}Ӵ,�_���ú����+$���wO�W�C�wli�|�EW�i	b���[=z%��0�gI�m��|�xM��GUH`�(
j>��$vE����#P{��O�؅|��
3��yg_�t�[�\6c:�*J��q �7s�M��
��Exv�N}���g����׽�]DxJ���=���c���|�_�,���%��� ��,���ׂ�ry�/3+óe5��^\\���b}7�+�-��
=���{���?Y�0;dC�B1�W��eE��J����+��q����6N�e��o�ȸ{�2���~��WFLk�R7�<�"|,�آ�?��g@%\����6o�㟸y�^�v�\\r����g�V{��q`Hs��"��D�Ѧ�܏��);@9�oJ��*gph:F�1�W��ZuSG��<�ګv�(	�,���|��(�[�}�z��O_wY{Ws����1�H7`�2��n��QL��S��;���b�j�>@_��՞�OE�3N(X&��仕�U_����u����N�˸���F��S�εq�f��zUOB�S'Po�o�]����wq[q��?�����T���[.蜱����\��j����{��8�
�H����;��Dq�nFzα���Gv{h���fPP*_jf���Z�t7����<�}�9���紐I{��&�~���/ò�=�TT^٬�P�+�82 R�
�οu��mi���q�dZ�f|�'�w0�}�&������Ͻv���J=�����B����H�jfI��q�U� X�<+��]�>X`0��O��=���������קb�F��=��s)U�����������ѥ$K&|{���IK�U��_�Q�n��xO��]��?z���1��J5��ߥ�s��ul;*�jC�����y8����ͽ�ߗR�4l\du7�I$w�_��#��-oA��.�_�l{�:;ި��X������̄�����~�hu͞b��3a�ӾK�ʜ��nr��ӏպ���zDKP���C�-H_��X������gm���OzJ7�N�)�ۢ�"�G�X����A�*�MzN^Y|���JOE�x�ܶ��'3��n��pm�n����g	0���NTü�"���WXR�m�#�%2��V3
��B�<w}W��9N��L�O�VƉ�j�>�l�������u��2��N�����@�����`_���*�g��3N؃|��%Q�>�yW�sD���l��]zv�u����0~o����g�=�L�yC9;K���xV��Z��Wȯ�>K�K-Q�E�����咬�\9�yCD�^:���Yb�9GN��Vww��I�L���w%�eP0�'��S�>��ƽ�g����ӛ��͘u��t����5G���,�X�j�BϽ� Ƈ��^��NTt`�B��<]p��|~�;���}U�C�9�Wq�3��K�Wx>9�^ɲ�*���aA����4������^h�}����Qr7>]~����~��|}"����FwGvWNz�`fzr=���?+�V�q8��}��xø=�|&������̜~^ʜwKޡ��?��ި���;�tj��0��G��D�'B�ڭus�3���*���1��f��F،7�#޼�������﫣���V�	9u�%��=��S��M!p����p��ѯ	Te��4����4�³NN���Q��%�U���cr�~nĲx-j�ϲ$E�T�Z�_X��)0J��jX,t�;q��.�ʅ>�Y0��\�dz�L]Zq(���iO��Q�0q��n1��]�/����Q뮉A�}4038hD��ɡ�#J�9�˴uW�����K�x�Ƣ�O����Њ�
8�|��s�i���a�cG Q���'*�>�>�\t��O�W�w·iS�v��&�'�(�Ao�1��
<��d��ϜzT4�*S�;��j�+g��f�)�^�y_r�����Q��mx�-L�~s�d�����%�V�A��y������&r��+���R��;a����	�U�%lh=H�����o�;�>��>mKn��M񦇷b1�[�&:�O��χ���=����9�{�]�=��>Yۈ�����qO��
�_�q�>���Ѷ:q�~�Rc����� ����3Y�_i�݁c�R����u�uU&!:����z�LU��9��>�q��Ȍ�&|��/B��"��%vD&�E�^��d3�=��P���Kg��vя�	������$JY��[�(٠��Os&��7븷�2�vC�3]깩ȍxjN���C���Þ�5��+��pF��>���O�>޿O��o/Ӊ��z�=�5���2aynZu񔶗p5�h�����@�·��ϳ�(����һ&s^�^��H5R�{@�����n�mm%��A�@ԫ�Z�@����Ʌ-�|���nm|#C�􃑝�º�TĲ�K�\K��{��l=��ڮ���V*f+��1d�%�lL��ݫj��`����n��ڙKQ��'@(�"�Ļ�	&;�����̋ס�g&6��g$bY����&Ƶ�EY!�%Xf�M�I�;�A����(&qE��yX�iv��̓�k�h��ao��7�7�E��ֺ�D��[Ӗ����Ա]���H�\nR�uy��<�.
S�ֳp�.����,�Z�Rkz�ߘD�r��T�l��,����9���u^��x��
�PL�G��T�e�.���&�qO��$��ֻ��T��J|��:���4xo�qr�d�ea�y�k[��PҨ�����gV�S]�����{oZ�\��l�pp��nR}|�ݣb��^�� �P��h�0�4��f,aٺf�W9;O�.�ٴ!�-�$�.��U\�z�=�Ǚ�^�V�;\I�,�M��5ή�ޜ;���q�?f��y'+U���r,���׻V�P�:������=��Ng/��	�A9���t���0��N���l���([:#�����Ɩt�-��cZe㮊!nD�d�b�^I��s���3o���0���q��J�;yN�M=������o7]'jK"%���o�r��.�,Q��4B>.�_�˹^�p�9G���q�fs��Go��p.�o�A:��K��&�Ѻu��ٝ�!9?����*j��(Ŋ���H;z�#�����gM��J.�2�����$�����q���nZC�eG��Q�cu8yJ� st(�9�t����.
���Ǣ@��p���7u>����k�Lюo,sD�y%��M>Mq�j��r�k��j]�ez{R����Q����x�ݰ�8-�iT�-��j,TBh�i�˶�kb���a�3�����D˝Aڅv��:{����I�A�J[�ݨ�Q�(u	h�G`���VJA��ޫ���Y�v)QVD��7�ڲ�\�v��oK֛�['R$;���o�nBJk�fЫk:	��C���~���ղ���auf��]9r+O���Z��zfsS'R�ׇ���X�jm�P���YS�:�� ��V�m�1�p��p۪��\t_df��om�ΣtMI-M���C�f��6m���(g�$t�n2;:�˗+)s���7}�15��5��{6��=�u�osS�`���Ǻ@��3�7�	�s�Εt0g^��0m�E��[����ẙ��G��wos	_�7d�{jP�oxҏ�B�X��'�,���w�U��ƻ�Ty/����j�;Tyڪݿ��޽G�������5j�.�Ů7���w�I�۽�����(�I L9�W
t]J��y';/*�M���W �먕&QNu��i$DQJ�����"���*�0�:9bW/R���:ȯ2��L��;O':v�$Zl9�J'"<�T��ҝ�)�'ZY!AZۺ�<�G �
�����:TAI��]���"� Ԩ3RKR�%4"(�\u"�-���7Z�(J"PJ�h�U]�\���@���u���"���E8���<�#37S��\'M����iҊ(���;�Qp��d���]vTr�Nu��e�HTEUr�]�Ȃ�q�M��eP���E���N�y��2�E�s�G9Q���^T�\���R��I�Sa��J�y�J8�NT%7=�<���E�Լ���ر�
��!n�t*rk*s��4�,+���y�DTs�*�Gp�CYD]��{����L��8��"�p.��t��]h�/z�sN�<�f��������������ku܌�E�_^M��c��i}��	�V)~A-�1o��s�1uzO۞W�ϙ'����#Q���4��c�m/;i��t/ЩHѷ`�!���4�Bp8��qs�f�����هr<W�	�蝅��=�\��[��\�K�0�|��/�t��CR��>u��2���W���.�b�];��]V�l�r=��^r=t�;��s�B/n�}��\?0V�	[����߿ �M�][���ђs�>�������8�6;�G�Ƕ�c�p2��
�H��ۯ��{}�i�]7��sˬ��b�n�\����g>�E{�r7�e��������FJ:D��Z	�m�������_���|UuEx��]?����늺n����vo���~T';7ح�Ӻv�k�}��T�yQ����J<>D��"h��ZS�s�l�b��\U�{֐��<���ӋkVo�|�0�����(��9E��Ԏ	��FD6vF�^�LW �Ti�/c�3:��8��wj�j�Uf;�=o�`z�@��1�ձR�ՠ�7q<D�p���Exw3��@mlX/��'
�.]�������p�oG�NT,�u���)ք�q���f�㡱�1�X�膐���e����^%�Z���>��ulܝ�yY�u�[:[�36��E��(!�/U��ζr���� ��v^%#{k�E.��'^�wY����0�ȍQ-�8��9�B]bz�m_�/��+=X�y�=��|�%� ��hvi�k�u��t��]�)h�ȏ+���qS�D�}�$�J��ޯL��������U0:��yg���y���^���G��­g�w]&8�o\l���8ߍ�o|fY����ں2�5�Lz�{ʵ�V��$Mz�{k@fFOp����tb�hy�U���lr�����UI鞝�N3�}c�o��7B���̟�X�HBl)jv�X�>��|���8εq�����Ӻ��������X�������0�����sB��U��'�?���{��6p(�����wœ��6r��3]�=s>����L�x�_�x�1����7�F{h��03)@�}���j�oj�tY��tb�S^�=�,̵^����p���FG��ñ�S�1�E}{f�_���.ͱ}�b|��z/��B����,�.:�f[Ȟ������X��u��~>�,�ڟOdU��S�[�މ{ܯoʵ}S��)���q�_�tYņ�0��<}�#��O��#}p�V˸�8 G�m;�`Q�+룴��kr蔳�V���-m�4�]�)܆Gi�r,���<�&���ږ����}�Qb�ޮ�|�l�d\�Ƣ��s�l�.
�ms)�'S��z���4&@�V�djn��VE�vX��Gv>k�Cݯ[�J�ǃ,����!���tqۉ��Ͻ,�2��|RD��R���)N>�^���ߴ[��/s=^y{�����Ӛ�F����j�m�r�QM0I�炎0���ˍ����emö�h91��fgR��i���[nvr�[C~�T��x���X�qt.�G��&��}Be6������!���JK���#g����EL���|�{������(�w&[[J}s5�s^���9������\��5����i�ۜ�{��VK��&Yf�O)��t��3|Wr>�3�"�ؖ��{��liP����:�W�-��H�G������/<�4����Z��#^�Eր���ġs�V>��Ͳ�8����~ۏd{�쎿��X�����������z6?}���_*��ͯ��鰮9m_����N���W\�{�Tqkb�z�������|BϽ��u��.�Xϴ0=!���}D�F��R�������ˮ���Cg��;n�}9�g�=;�J�{�nk�4�0���l�37��FF��&c������'gv�]��}��s�`l\��۫ŉ�+��ݍS�[n����$U��S���<����j�ϒyr��}��uQ�ke��s8�K�1+�L���K���+'m�1�-5�h��qƐ!��|�d�N�_cDC�Qb���f��7z�Y�4F�(�� ��ϡu��;�W��gǼ)��Ôy����]9몛�>;u�]��;K>ԯ�W�r#l{��c�m���DN�L�?/]JwKޡ�Q�iyWO�g|%ܾ��;����\�{'��(z�.�v�*����0�:�vE�Ӊ��f]���	������7���ｼV��kN�$f|�3�ظXh
�["!�@/>�'Ɯ��i�}�r�W�c��_Oj�uu�ՏT��R�`L6;��w������t$q�Nf�y7hׅ>��w�h=�ͯu{�^����W;�ro��~���G��Ϸ�X�~w�W��n��I9G&,�Pɯ��U?u����k�N�|����}f+�����f���{9�|���q�R0e�Wtj������yw�ܟI�r�LNׅ9����6(`�!o����,S�!�����.=��Ȉp:ߌ�u$�{_�וP�w"e�C�5M������B�|��Z~��@�gx̥�iH�<�(���y�#мrd���Lh4ر�&���(�cg[�/ܤ��x�[��&/�N���-���o�vά����ZjK]�J�UXJ����Ձ8���_;8S�ÙK[�2v�R4�mwkU|����X�"��y�Vr���O����Ds���ZγV��oo�|
6�7zf��-d|�s�.=��y��h�xt�<��CA�*d���Z��{����|�/�=Y�=��LӢ�T�տ
�^�W"�w�ʍ�_s�UV�RX�/׹���Ϟ��BS|I�dP��^��:����� ���>ٯ`����"LW�V���Tvj� ���p9�}=}뼗-��)K���rL�xjA����n:�z-��M�MF>Ez1z&���>�ъ��yoܯ���l�z'�>�zO?u���Q�E�?N��^��q��m��=R�����7Lz�_�Ȁi�3���.#���r'�ꭇ�΂&������E���k�`�����J��\uzF���TV���߁��φӉ1���2�K,sFks7ַ��oD����m��v}��,G8ʭ���6�*�ᚮ�q�}c�>��h�m/I�~ ��*c
�L�t�E�����/ñڸ��g��ѶW�ሑ\��^�����bz��Y��<��*;�e��>�7�<};��}�iO�A�	vB�0f���{�;�!��w�|=�.o�Qt��)�0��=����W�77�e��[�pʺ��:��|�V��>��Ԝ�C_�8�:s��R0T	�q��>ޙ!�4��E?)kek	���X�_A��xu��#K\"�	�4�L�tZȶ4� n�;���{�pm�Clwcme��"�bXS�	����٩Z�E�?@{;W��S��v��k5�\�8ssw����3��D���x�a��q^�늿�����>u�7�e�Q��4'����#�o�k��	�C'%�H�<~U3-Q�u3_Ϥ_�)����2����HX������D������h�÷^��S���~�(UR?8
Q�5M��p���u��F�z���G�I�S%i��<���؏g_������?2X�?*��W �7Br,��2���������QNs;i��4��k��{ܬO\&���}�G���`<�ȗN�f�T���1�֫e�W{e/H6�_����YG=����}��O����ٛ���ȟW�{�;ə~5R3�r������
2/��g$w�z��D��b��K�h��w�=��Ͻ�l�{�2Ϳ_���-tze3��w�u��5�2�
k�����Y^�Ӻ;�hy�U�������QAz_�_w���)�צY�κ��<�'�Įb�?�6�:X=*���e�~�t�٩�W�ެJ&�٢�����J��ȿF{�4^�;�+���W_��b�j[u_�Q*��%~7b!���a*������V����=���������A�XzCY��-,��' nJw��`�%���SG��<��;&[���A�GP����d}V�=OK]�_u�>�p*��VNU'-��[����eo�A�=B��RUӚ��6T��s�=38���Fzα���>�#=uZ�3�x�`󨫕 �rSU~��X�txM*�j2��1��
���_�dzϼ;!�S�2WI�;h�y�ސ�z��o�-��=ʽ`m�B�E#�:��]L���w0�G�bq��V����}�>�q�:�(�>^��n�׻Q>��uR���-@�a�u��]T���>�W�(�T�{c%k�ߙ�����y��f�����]<v���.��������G ���GYlzrY��_��6=�z����sݦ�x�[�o�Gp��F���������iTSR�'�!G�N�(j���Ӯ�<o]�Ù��73su���W�ɺ~�;)����::��x��%�P@A�̥>�/��*��>$r�~�������k�(n��xWJ��zԩȯyۜ����������00��0���^#|�t^����[��f��4����Q�^A��c���zm?;s��(g���`\y�L���ù���>����L���3����5}��1]68�5p�/���m���H�sC�w+*oKS��TP/e��n����6�pF�d��+@	2�lUå�P�]�qk$^�����I��� mBK��z���rvJ�H9��]�`GR]He���Ε���O1�"�@�>�Ϋp��/5�;"��[`�X����q����}G��)������4�Q�L�*���s�X��oM/!�Z5{>�͝�mn�X�U]v��zG�*^���x���]ɎʠaT0���=/z��ӝm_������bX�5����\,��v�>�W���f��<p�����^��ӕ_ӧe��z��8��aś}�����;E����s�ۼ�N&|�ӱ�J�~Tf�=W�ߎa�^HT�ɏ٢U޽G�u-H���M-�[ဣ�7[����~�^��Ǽy����]%��N�����Ye��3�X��+�L��`4a�[w� ~���̜~^ʜ�t���1��G��0�j�k[Ƶ~�ct��x�@p6s�[9�B����:���x/�x̻���zr��s��w3۝��N�Y}�p�Y��\wg�Ԝ��7n�j����t��'Ɯ��	�;�FxW�}��@6�&�,���h��^3>ѐ�^�Y���{�U�1v
B�Б�S��A�=0Ź�33�\*�ާ6�u�z��Xk���7�~���;���w�,k�0�A���&���N�;�k����Ѽ��%3Ok�{KJ�\� m��&�����L���J���Y�S��8��ѧ��ѯ{'q�t^�ĩ6J�p���wLA;Q�@�.�S[����{kor�;���1�c�I�Sa�v�\r�bnt��X�]D�Δ�[�����Y���3��uSq�^~�}f+��gI��oײ���9��3��Ԥ`0�0��(�d;�]�{ެޣ�Ǿ�1)�f��x��^w�`�!p������,S.��j~=< ��s!�Ӕ���o׷�~"jP/�~H��
'�G�Gt�T5G5�`�#Z��̍��m�>�^�_��Z�j-k����m��,<�Y#͜�?C�b����4�I���T+-���)�3��C�ǰ�ɮY����"}�+��W���g���E�T��0*�z��X�x\������z�^U��z)���}���_�x����숸m���ޯD������X�
��&�E����1�S5�>8#�V/<������x�{�M˖�I�D=�i?UMo|�I�wU!�2��^'���fj��!�����݉u��Q�_<��_4�e�q2|�|���V{�&�mc��y�ye�E���%{w�C�}���6FJb��tr��O�ы��\gZ�K��g��{����2*���-vP>�j���m��{'�YC.:�#F�x'�e��xl@4���q=;K��aE'��N�=q��g�|;%j/��a9�����rw�9�r�'�nP�I��x���V��N	n�u�T�:�|�t8�-�ˊ�]�+M�îM:z��Y��}�p����!��������^��wl���)
͸��.[��~7o1������O��%Wð{*�mz����+����Lߎ��\���~c)�:���F�g��{�3.�w��-2�=#Ɵ��v�;��q9�kE�`y\
s�+_Y^2|�է{���,9�+%���KQ=�r�4x�D�8���?x,�YS��| ��4�k�x��m��,�o,N{{@���R�5^.�,��������{9������̾�~�>�+�3d��)~oR#�ȟT�n�� <bC��E��Yr�����qWMߴb�O�sV6_?F�\��m���w�k�x����t�@Il��O�&L����)������/���=\v��w�I�������|6=��P��Qb��p��qM��q���B�}�&}�+ەY�o�z�oݣ�iO�B%ޖ����.<�0�b�ª�pCw�J7�ے�
;`�o܍�yW完����G�z}q�V'�5~�9�V<2 z���Qq;�S(9ꏳ/!�#��v�i�oE㉧bV"��˦��|��~�t��0d6��ˉ�I�<����[�����`��������l���`���l6���6m����cm��`����������o�`�1���l�[����`�1��C����0l���`���l6����cm�̓`���`�1����
�2�����  �����?���>�������;w��*� ABQ�@�RB��)IU EPPPH$���@&�zz��U
�JQ@PH���R ���� T�*���U$�P
�
�"�]�B��ED��BJE	PA��RQED�D�T�� H�P$BD��:ª�	  	�H�LF���U���mU6��M�T�b��b��Y�(�P�JEH )�  ���iY�%(l����e��h�.��>����E)���2������`覚)Jn8ҁJP(XUѥ	�$%ٔ�I�  �$]�jж�l�k4m�հ�!P�Sc*֨���ZS�M�P͵��

�J��)8  r���FP��ՠ!��� ��
��Uk!A�hba�J�T2UTHEHP  e�U"F�Zԋ�Р�6�Tm��j�5f��m�[h#���UT�c	�)CZ�kmUUK)6b�(�I@R�� �u�Ԫ�V`&�m�jF�FH��J�ŭ�ي��"�V��RMB�h�[F�EUM�$�DA�)+� -\*��ZҤ�ZRͪ�k	m��Uh5X�٤��
�Q�E*�L64īb��
֭���)*��
EJ� j��3Ҡ�X��Mk���E��Q*�aj�U�Ml�)@�����Fj�JC�J�UTR�6��	� vٕUT�-J�U���L*�`�JJS	XU��b��f�0FJ�UiZm�E���R�5QEU�Ak8 ��!��K[l�`��Km�hP͵Z3ch�
*�0i����V��ʄ(@ 
  b&�RT�0�� ` 4фS�)H� 1     HИ�ИM1
z��j=��4�i=4�T� JT��LL&�a0 4`��=T�SS�I�H6�  40���EBaT�L&M010 �e�=�L�v�v�=v�e]�!$�<��Z5$1��}�(������Pv(� �/UA� R��|�?R�s\�
�`-��߷3��;���{��e����+p�X��*F@��(� [��w^���{��ALP�Q�C"����1��2���()�2( �V��-�=�3���ff�"""MQAD�Q  �uEPCT@5AE]P�� ��V���	 ���@�$ ��$!'����B�]u�]{��I%�$�đI$����;!�o�^.�=y�Ay��Cg����FyyU����"��A#<f��`����`�Uj�*�#HV�P��p�P�0��ݥW��r�,G�ؔk씗�E)�������J��2i��P*RФ77��3T�w��c��Wb�F�����wj*����m���,��o>Ӝ_�di�u��s��U��)�K���t�U٥����6��_��Q;Vt��Y��E��v��M4,<�31�#wc�XM4��֤��6����
�	%UQ�oMm�[ʍ�0��l�\��ne3��.���m���g4���M-5L<����Pڿ�DM�Y�]���B��\AL5媹Y�2Z�7u�e�w�n���ʇu�j���e��giX���Ck:�$iV]�g!3*�7w~T�{sp�B�����+��\��;,@Av��T��6�+����V�4�[�d�H1B�r�`{����T����y��G*�{qW���:��yMEw<=�xHM<�;���m��V�CK7l��ѭ�ĺW,`��/�2�9l��lݹAШjm��Ĵ8�\uf�򔙙&Fe�e-�R%Y�p��B�YGHxi��,v�A��u�.�)�x��yT�EU�mh]<�Y�{�YY��7E!pmP˚r���<�*f��ae[�fd�,NhkSWCV,;�8�T����6���.քP��m��A,AN���ŗ�uE�tFK���V��v��vd�$aVQ�n�1zX�e�藦�j�e�����LU�l@��+�'u�lR�����lD��sv�ĦL�{�"U��wr=!g2'�lեj�$��V��m�b����6�::�Xܣ֎YV�<��{M�6�7�7j���*	������F�B�9Na;UA$��U�rm4Y�W��fU-˹`�j���a�J�G^al�9�h��W��-Ӵ�zա������������vH�t�",���w�V�Y	=�jn}qt]]=�J]���j�f	u�[M=�)�*3�[�㗴�ǖICh��#���ė<�q��w;t�X_9�]���^��,���M�����b�u[1���u�'w�l�˯��]:wCn��#r���۰�t�2q\��Vj��c���{�WW6V���ͫnB���V��k]|ԑ<,�j��.�+8��r	>��l��i��a�k��mo��#~�C�"ي�յ�V��u2�T/q�������5]]5P��35�����Sh<�b`��A�e�P�0���ś+Y"�6jP۰���7�@Q�5|9���wy� ���Mg:b�v�-��MM��&�Հ���Zt,�Y��iilM���ڷϓ�������|8����xE&5��)]����q�ճ�޽]�kH}���U��H��'sG[����щ[[w���b'aQ-��U�˗[ج�4e�QhS��c�T���/*��WO#,)��k!�MHU�ۆ��8�h�-m4��hL`�".���wJv�9Z)�VK�����i4;�w����m�ج�@�%�[��85���c;���+d'0��n��5���8t`zj[ز:"��e ����Z���gNd�oO�K�C�9-��|2��h�%m�{2�,A�)��Uoj<&tV��X,������N��+_0c�K�s-ٽȻ`��M�:�Hg���vŰ��Gx���t��>Z��}cp�����e�4��[�|[�v�,�JE���B�^�h�&���$C��<W��̺�͚����Sַ4��C�2n5E#t�ۚ���{mE)�"�*�5��IQ�Y�3df�9g��[L#{\�D�Ė+:�q1��J���.��n��AJ�d��ʫ���{{;�H��w_,ygp�R�����oX�ev봊�Gz��u��F�e�ڱ�h]b�{���OFY����S���qd����ʢ�a��D�0Y��,�1C��ЉՐ��h5y�ilR�F�uut$�:��賻/U�j!�(�u�	/qE������:�a5�֣�`�՜�,ov����_^u���%��/B,^r�i�ZoM���^=4;�ҩp�Z�H��opjyu�+�r�,7�x�u�V�gq�������CF�5�#3׏e'��jR��44��t��b:��i�4�Y��v��[V��׹Blf������.��1S�;������С>���&��A�u$v1�F6�āie��6���cBb�q�$��wheGZ��:x�G�uI��cQ ��[��'X�3�kB��	F���#)�W��m:�5���YѨ�zHbN�vʽ;o��xj�� ������{w��B���[\�60�������%�f�`
�W[��&�w�ǆ�Z�1ն�S�g�X��8�L����ɗ��µU۾٧�1�������{uQ��tm[K
F�vn��^W$vRD�ۚ�0�c6���)x~y��Pt�3U�r�ѢG�V��{��(��҆���nSTl�"jĚ�jQ���l�w�[
蝼��1�M]
�0�V����lf��VR1��j73[g��V����j�M����U��T�� FX�9
��[��pm`��֦M�I���&��ul��7���(������Kq����\`{�;x��'��s\^��$rءeej��c�P:�ݔN�=��m�e�dmrѱwlP;u󼒴�"��`���e,�;�%3ьИ����mb;Y�&5^��c�����3[j���k��m�܂�'��H;�Q0�|�2��Xs^J�-D�]6-��!��6�e-�ݡRZE�)])v��X�T6�HZ�j��E���e�@������Y����{�|�W�ԉ�v,*Ȍ��,�ͬE�e�p� ��)�NV�w����h*(��Q#n��X���y�F#��Ǌ*p�	��� �,�X1c���u.Ÿ���N�&�8��,��Sv/�E���P�;4�u�\������w]=ڊB���ͭ�ح�tb.nT#pfn�<�͠1��oP1��Ǖ��h��&�0��%�;���Ҭ�u�bLZ����svѫ�xԲ������r��)���N� o�ٰӮ�ݼ-,�"�4M��&Ҵ�٩b��{t���A�i��]�N��)Co+�z-��F�ۻ����I�n�ʵ���]v����݄d��`�Sώ&���Rͥ����z�zӁ�:�ǩ�7��f��8�8��>��u�[�ۥi�2�Y��ݫۺW��x,]o���4 ���7�5����O�����f�n8�k��f�X�Mb����åPu�|�l4-��n���j�MF��.���]�,�ν��Q�f�i��֪/l;�l���xq=�ŃkC�j�T���Ϡ��mXd]��U�qA�rJ�Qb3-K+Z�&t��,�XN�2�Xh��$f�aJb3�a@Ƃj���!TUT%��]9"�P*I���h�&���p9�D�XGk7u^�����MR��-��E`)��z��=ŉf�\�(X�,��h��׎��T2�3��Rz�k;1�{�Ɂ$�`�Ո*i2��v.�=:f��_<X����=O4p"�6-Z�L�E,ܹ��,^���eY�`��J�Fv���iYւ�a�|�}z9�Ŕ+E�@l�n��,�Vu�L���4qRm�Żv석o$O0�ݲ��+|��h�U��hz���l7�'�N7��yu�ұ�t�)j�o�y��oF�*�u}a�l_3�� 1�
��2�iFѳ��L.��:�4�2bz���yxM)��:���w#�D����N��`W[\s+jh���U^`�[���t`���M�ϴ�GE.��{��͢E���y�{�Z���NY�D��c!v]k��uq�ƶ�u��5�lݣW34<��JAG7-�w*\�N�F-`��R�Bw�{FTK*�sD��\�5P�ЩR�L9Ts0�B9�M~�.���l�[<_v,X@�lqGI�͵@�=�kuLG�F�Gͬ�Y�c�tw+h�6��t�:4�O7)ڦ�յHᑝ�:���dijigBwYo QABV�������z�(�W�d2���:�bVf'D�:���J���5�F�T����B)JB#6�W���R�2r�n�{z.��n��w��wA.���F*�z\ʡS2���L��ŵ�
�������8�X5�-OkW|�m0�
�O���j����XB���m�d��u���TEGd�����z6��mR�QM�J�o2�E��eu݃:����Ǽ����Q���F�8�R�d^�
A�*�)Fhwwq���>8z��j�E:�sH{���.Eҫ����\�.�c��#n�u��T�rMX�8nԥ�e�+L�]3)$�ٸ";�D�0�f� 2�5�!�����@L]��)iH�Vm#M#e�������B�{�Ng=�3-̠]d��ڶ�^Cn2�׻V����J'.`yz��d]-�#���[�K8jX��u�a� @ku�|�K,5w��W
�P���� �Y�VU1R��x�e[m��g~zJ=�	�kZ�.����m�v]�ˡ��k	�c��+����Nfn�p�Wb�S�wF��n����(�Iq�Z�7[F�צ�±�-����.�,/� ��y��k�o7��b�9a��$ca�������jZQ�S�:4���Å"��L�5��;×Y:2���t�ѯh��Ίǯ���U�Q�'l�uZckJ@�Z/n�ePܲ-n�.4J-�CZu���o����̙Q��Jǚ��+U�E�YL7@`$[1,.μ�Kú�[��u�:��2�oe�;�l��[�pV*m�G3s3$�hV	i��f�轪[R(��B"�e^,!(fm����L���`�K=tn�˽���(�aދ{���Y��/\څ�*1Cm��g��9�k6�o3*��F���F1�]��eV��xF+[�Cc���J:)o���A$��s,fĉ�Uj豯(7�7��3x5yQ7ooq��K2�&vnҴ���9n'�Fhkld�bǛg/`���\ ��8�J�f�s\˩M��tl�:j��Ֆ�6��a������:,�(�������%(��W U���a�F�ȯ.�a�k��+��1g|
�]��Ӭd�z�o���V���Hwm�ӱ)T��dN��V��"��G,��E��|RTE�����X�BEu(!���0�Y���h{�ЬĂH�聎�n��m�gR��"�&�k���u���˯�{8�V��b0]벑�\٤���s�W&�7������m�I˵T���gs��SZ�&kgw',�¹�E8S�y�{`�b�}��э�=iR�G���v���X��U3�G�g��VD�4R�ܪ�c��6�cUՅÅ�j��gv�+Fi���ޡs��qD��v�=a��F��b���5oS`=͏JSR��꒷-��f��[ܶ�,m;�c���om���p�m֗�\�^��=о�n��6�޺xx ��������3���m6��Y�cA�n�м��u����j��3�6�z��hk��}���dP蓊h�W�[m������1R��������A��FՅ.TY������
�YZ]���6i�`� w���t�R�tl	&&6v��M��¡Yy�u"���W�#�yw�'̱��PU���k��f37p$��>�N%��w>��ɹ��#[�+���lת|��q���=��*���IX�z�w���%�K�][�Z�(N��k/��4mkG�{��j�`�Cőa� ҔF�[R��e���p�5�A�UK$pz]�jeŷڻAY���'8�h�y���:�.r�j��pM�u�B�n�s�7Q�[Ȱ;�P]�FtJX�,|nr�]�(;-��s9�f3C���T�%
��R$l%x�V�Oo B��sjIYYr�Pqg��<5J�K�ܣ{�T�s&V�;v��]`�s�N��^)��Q]G�3p1����}h�>Z/�N&�ό�S�����Ձcک.�1��<u�����[�[gR��Ü�FD��5;��M��N����K��G�4P�����2�#U7��05�*��K9��	�0E��<��%�޼=��7��'e�ހ��VTn���!�wWZ*�:��qi"@���3���9qs}Q����b���J˭y��IĞpT`���
��EZ�3��|��"e�(ڛ�x}�79h"��^��nV��d��c;95����(�1�m�9�v^_�@k�y�q�Ν�%�˴���*�P�VCQNY�o%�0�[�G���mf�C���=��x�z��<	7)|�4��a��}/uL+ؠw�w��S c�\ݓ&=���Թ �̷ܰ�dD�,<eM�&��f���ˈ��+8�(%�{�8.��!��Y��|����Ռ2�^�ç=�����CL�GV9U�Z��e��4u��f,
�at��{��Id������ak�0r�u��v���D��F)���`���M�Y������@I<�9B�,�e�e�$ͣ/.����s���0�/3gC5A�7�Z+�`��1�V1yi���W5��#���ծ�.��ӄIF�j�2QHA��tm>���.��z�gYP�xv<'!�8Q�����v��8���FHmD%�Z����T�b=Suo��?*�F�tLV�� d,*R��]�0� uWE�_��E3��N�po8��.���fgl�,��6�X+9����m�W�
L^	�{��m�<o��1������G/]�y�\�/�̠�}�R��m��dR��gT���Z�,9}�3&@n�R����xI�w%X�A���ЮR�Y[�\M+���e}.Q��N�Jۂq��"�v�4f�2��+|��7
�vv��
(�<T��?^���0�vy��A�gf����ȝSo�-�%׈e�d%2x�tg��fm�k1ՙ��ݦ*�뱢�+q�L���8�є7�D��45.*β/o&�ghH���DW[Iq�ڃ+JtN�c��v�9W���S�zuz� ���2��I뉽�w�|�Ͷ��0���`�wٙ*B�k!��,G�-�.r��[5n3�!��ͺ)�
���c���ly{���C�3Hy�'dX�&�c��e�g�6�
=�u�}Q��>Զ�I�sVps�;4�	j|j�Q�̎zw�q�=ӽ���4��1M8e�P�+Iyg+/2}ƺ��:�!�۽�̆���·L��d���� ����C�Z�|�۲3i;V�DqQ�ĳ��n��%����-�8���$C�7ɭ;[o"ȹ;ɻ��w.ÙVwtƈ\�|У�܃}��KAA�z�3z�9�6��t(W5g��T�0tw]٬�E����@�w-u���<A��)t��Ҝ��|�f�<�r��4w�2�,�P���Th�}B��,�SD�4�3�C/r<|7M�*ƺ7�+fJFXl�ڹ_e�;�1�� t����<����˒�$���[�p��y]CW��'�V�M�y6f.��R	;��J��QN�IFž��dg	�.�����O�[2�Ieq @32�y�'{��K�r�23�\su�P)��:�`k�' �������m%���Df,fSS5]�kw7�l; �J[ġ�a�lW1𻛼XW�y�W�Ԯ+IN�5�=��υ�s���n�Q��r�1�>�"9}�F
�c��W74d0�1b��fTR0,��{�� X����kI��]���UP�o���V��Cg�?��0ҥ�\�Vd�o��n�hh=��Y0�Ka�c��UC�s"_b6j��h��e���`����uvP�(͡6
�s xT#*����B��#��(�Z��g8䦵���*��2/�XFu���M�Y�
�6�C1&k�n��_��ǭ�!�f	�ܦ��3;u���F��;I�l�q��u�g��P9n�m�!���b��O��v��zW&Fޱ$�1��-5���]��Y!��a�A�������Z��_fQﶀ
�3V��)g?�\�J�9��M3��;y1˰�|V�Ҕ��B�ʢ�oL��T�p����=X��u��u��2�������D9���ɛ���9rü��ݨ��6꫁�A2<[4����v`um̈�&O`ِ=�J�r�,���Њ�H��q�X�w��QX��]�5\{�o:�`��Z���we��L�#_!ZX=e�Vq��,^����#�ǜ�Fw0��s�.���K��܉hu�Z�)<����,	�/b�p�Oj}{�U�}p��s��8�u�Y��sh���AjY7�s�۪�����O&�ƾR��S�����z��K�&ȯ�-��}��8�2�SS)N%�.����#��껊���gN��6���w���Q��]��woQ��F�n�r��Yf|��)�,�i�Z�ԍ��Ghdy*�^W48��wC��_Θ�l�%�פ��x�n���w�!{��w��ˉ��잖���\L'�9���U��`��V�b�`�1n�M�S_�$���/
�i8v�C�W�:�q�),�]��;��i,n<o���G���su���݂l^>�Y̪�+ha��z��t�G� V3/�N��5�S��Sp��F��V�e��=7r`�]*%[܏d����Kb�Um�	l\�3d���z:�p�n����/es�h�p��B��o�f�����}��!&��v��q�g�MLm������w|9';�.�)�Z�p���c�=�r������J�X=�:�v�XE͛Zے����.^�I�L��ʤ.��ĭt94b��3tT�fK8��v�7^J%�^��\����;Jz�-,�ۇf��]�ո�ffC���=s�ō�.��m�_-PV��r��&��q����I$�ǔqb�Z\�/��>��W<����MGnM���B���uٜ[:j�=�W���5����u�&�VNAE7�����.=3/��n���V�)�^�h�Œ]�RN����7��S:\Of���s���5�4�ف������C�s�v�_.Y��.�
mE�{x+Tfc�=;���Z�gm��6"3��EK�:`��Ɂ�����:�P��0k�qiMwD�S���k���z��{w}n��kV�A���Nk��I�Aȵ��S�1��P�N�s@��ὣKZ�y'q���u�^�9%n��`w���aV��v�
��RAS�&Pm� 2�C�h�$�bͬ���=
�y�əSP�IwwrTZ��OLwΎU�?vJ�`"�u+�m�2���
�Ȝ����<rl��k�2�U:<�����p�;b���9�ܦ6�%Gf��3Z�<��a��O3���eȴ�L�v%\1�tb!��׭�dug -���d�C�K��e
�V��vٗs�)1}j��t3j��j�8�4�R��C�~��:~��,0����Di\��������,c��/10�;V0V�I6a�L�,p��6�C�#��d�+[����<�r���T��ؘ��C��le1�]��j���Hw;�U&�q���͒�<�i���[�(�.G2kgJ�%s�L�9��V���v�"�x�ﻕ	��^�%�Ǆ"q�o�iVE�5�n��[KsUH���ڷ�Nm�P�QU�\}w.ĳs�-M��;mn ������ù�{���۾m.���Q��z���9Ve�"��;���X&����tG�X�1�F.�p!�2ٳ[���w@;�e�jh���O 8K[[e�S.��/T��N՚z (>���L�,pt��X���k���y�M3����1t��`{�5����+�(�RZU}��3�(2^�9�r���:�]1v�r
����h�^�I,�G��ok�P֧���]ABᆬ+�f+Kz�D6�tڒe]p+i��-
ĜY�.����u;Sާ�t��Q�kΡo�&&S�=��j��-�ͮ\}WJ�WH����/F
��jp�o�a��X���$鋱�#��(�Y�ᜌ
��h�T+�ܻ�����*)�7������5Gnj��9P��d�<�ԳE|�v&4]�a48�㒗uÁ�ݝ�^Э�$,���S�*�3�˅�R����W�7�=(M�ώ�t8�gOlΔ�զm��S�&n]6^�e���Z���|�ћ��/���a�F�x���۵i����&�_f��p�ˏ4��(L���.:F�w�s�uWQT�@Wh��M�Ul��(����x��G5$��Yf
�W�1^�ZC�t���#�̤�\����D���٧l���_45����Egff�X�k���Cs삜��M�h3Nd����,��orp��n�D^��-�٪hШ��v���t�q��l2�X�`96�@   ��ėfVX��VJ ����噆 ��&�4�*B�@9��UM�A�G��3�w���g�F�Ɋ�e蒉QUWYI����j�n<˖���n_f��U�F��8ްyӎ̦Li!�_R{��6���i�b@ k���R�z�<:5^���]����v�ʵK���S�3  JU�@��{�a����������'�[Z�p�w
��6�^���h3J>Vn�#���(H�3�5D΂-�[Y��δB�3�;[������8i����d/�c����U�aޙ�<�9V�u��Ş�7:܂�7�F����Z�	��4��)���,����Ƒ�ݮ챒���Zي��e�BIM�0�v�f�ᶩM�QU�[��A�*.E���ޗ8#�5��P�ﹺer��Cnmd���{�ω�U�*�ڗ��uD#=�Z�u�o����{(c���sX���'n��^����%�m#ۑ�� ��{[A��>#S۠�9�鵻x�ܡy�U�5��y�����G�1�ސ�6،��i����[���NwHs\&����Խ�wҜBfX�	Vl�O3�#	�Tށ�G�oy��	���{n Y�rs�G�Z[��a�Cp�c.�)nKpV[��6�3;D��1a�Š����μ��l*"٧̌ȗ��no��y�J�v\����Z�Z �`�a\Y�S��?�-�v#��z��ZE[�������V����r;�x�>���B˼3W����9;tR�,��x"ps��o�˒��;��سBw�ܠ���:Y�S����Pb�e�{zD�#��M�1>��N�Z�9S������Y�4��y��l�\�1%ZÀ�Ѐ�pN@uoh�-��F��W�X��Q�����6����ݲ-�Y����a���v��łoZ-�r�m��cy��9�9e�Y�0j���ω�XK����N�h̪xʃ#��bwx1j&�Bk��K4L�{Z�f�_\��&]�lb ����cy�X��{���p=qv^�7Y/h����$�H����1d�.����:���er��CF\���%C�3��볛���v��M&m���zɵ&M�:j�"3-d�&A%�2�SW����P��y<O�=�Z܀�;Q��أ�wݽH�R�N�ceY��ZxV(�9y�g��z:����������Z�(�T�1��[5kEn�L͋�޾�d���EqJ�S$<r]yo��Ig_	(ԙX
�ڤA����q�;0����e�;��r:5���z�;��$ٿ�7]��!�ݳS& ݪuwtDTj=�dc�k�H�\��a���k�=u����o*�)�i15�]+wDy��*��y�m]S��u�mu��`��mr��w�� �+ac ���[
ޏ�F���u�62㛴{������k>���u��[7�s������:�A�/t٦wd�KrL��ȵl7+br{r�t�}b]&ᚁ͟u��d�3�r���iL�2���9D�1}f��+� Y�Z���fK�{�c�f��k��,��:�фv{��F	[9Z��HVvu08gǥ�S��B�� �.eM�ܕ��RG��pܽɍq��ੈ��XT#��ǋ����ձ��G톦�2S����>-*�v�X�͓9���+�0^+��_˷d��|殮��$��'�45��9;�Y�ۉ�C��N	S�&�6/4/�C˺+dom���g4gVЍL��/s���QaD)Rk�.�1��q�����m]MZ~�2���c��+�f�<��r�0��r��.�#(��[{&�l�vN_q�V������]��̶�H{���N!��V-�G1Ƶ�m:|�.3�;n�(Һ4��˕��m�O�^N��Z^�Nd��R��K_d���; k��%����d}n]�zj�*���Y�*�2Ŀ��/dέ���Jq��+�"n�l���d�1�k���Xޣ���n)����|*�9�`�6�ޮ��"^�룍v��Vᓖ}��]���0���gT�jդKN�L=T�uF�W>䅧m�B���sy�Q�_0%�ig%Y��/\�u҇s���Һ����U�p��+&)Z�s�]�Z���©�v�����\����
��b2&!-Vջ��Pd�܉\�+��q�%q���V�q%4�-�4��\bM�e�E,ە;���Mwi�:�j�W�iREp�@�g1�7��NGi���Z���^��x*���(f��\���b�h�<�m��=D���Zݝ����(���4P9YV��`����V��w41nIF����� �
��:4w }Ƞ�z&�ၮܭT��&�7O���f3�OR�W/���.��*×|���=�j���˟���������{�p�B)�f�(ݥʔ�;��K������Z�l�[\�q;�rE��w:�bt
\��j�Ɯ���*��Z�vayV��+C#X1R�]�a9XfQ�t�D��waݾ�V ���Vm'��'6Vj�ń�Gm��P��	N���\���%>oz�������>Uaݍ���u2��f,��&c��W{Y����XSr`�}2�nWVF���e����i��GY�Y-����$Ѽ��G8�\�8��;mٗw���o�d]1���U�*��w�+���3��\Q��F�j�Zs.��f��2��<3��ھc�9*�;#IޡA��LХ�wL�9��e9���6ЩX��9Y�p�	x��ų+]���t��kJ�S�k��:8݃X�s��e���ܾ���V9P�6��z���cp�m�')I��w��\�e5@\�Zc�
���p5i��c�dR���Ps����S��U<ޫ/IF|Y����B،V#�4��.TJլ�h��d[F7��[#�{B�Z�:�v)4�ʇt�fӕt�t����=eY���o��a�,��ӓx*O;h���1��)r����C�f0����V�oM5OD�I�n���]�/�Zma����9�5sCB�5u���D7l�
x{+�Y0tx�0���v�z�R�4���CY�#��pQӘ,:���jc�+c�޺�7O��R�ñ*okoJeX=�E=�s6�=����I����:�����ﮒ��}z�b�b��'����+�(Zr�-�A9��G5ԣJ�6�������|�;�\[-��wE5�^G)9��qᶢ��r�)�����T8,ν�}+\���J�L�	��8l�|P"n`��4ᇍ����Y���RʖF�x]�[�P;7pp�X+'�MN.��-ܫ� �aVX��œ�C3�3�kݺ��Η�<��J��w.DqV�=��Ś�$�US�W�KM��{�k��&.�**��SP�4�����خa�Q,:W���Z7�9텴�q��2��v7�B_M-��q���˺�DI��Tw_$��0���z�9�;/�Q���\{:�2�(�=���,={q=�tPv��N��,�-4��!�ۙT)âaj΄쇜]��SmN�I��/,"���	ފ�u�q2��ﮧ>�k�)��%�V�k��Q
ej�zdf�����j�Z�ۥ�櫢��%�+��6h
W,�e���'.�tr�u2n�ky)�W�c�*�nY]�;�BCǵeNFݮ]�MKI⪗1�Zq�EZ��<��=��S�k7s��	ُ6�^��7Fz%췠=W�{T�ˤ�|F>8�m\ԯ:�p:a˴:��N��0�1������b�pƴ�8�Փ��yΨ9!rȈފ�[��o�![sZ�iVU櫮l]�E�4a]/��2<7�J�x�u������䮒�T��RЁ�^���ޥ�+Kn�8'���
�5��4Vʎ�&�H�P��&NY�|�*y���E�M����G��l�%�nr�|x�n���C'��g8Ȭ�V�ռ�u�2T�=�B|&��W�1�S�b���GUp8ҧ�ݣ9Lh���c�F{���'*���u��k�r�'��}Y���*L,��A��"���W�u�]0ܮw0)`Ш��K ��+I�c��
�R���w�����*��c!O�m�w�#G���^��b�UYo&�	n�L��C15ҷ)菭}l=�"q�9yC!��i葋J�3 yZ��Y�pu���|�9��j��F�N�Y�X�Ժ���Dj|��Xڻi���p/�����}�@8��w�{�D�s��#�	Ќ;��͹� �̨�&s]��^.���&����4��x�G�/(.��
�v��@�K�S���\�P@�*�QSq�X7��j�[�uW-�p�`���s�[2��%:�f����;��U�����`�£�J�N��w�U�N���t�B+�-��ҁ
�Ӎeds�e��!==��5��S;v��8�\�fVp]�ؽK��Z����q�����c�f��}�a$�v���*�X:0�͡m��R{��x�ҋ����:��������g��2k�7����\}�H�ꔖ�k��Un�)\5B���C��E��ٹ�oT$U	4�7R`G���ō�j��.lN��GN���۰�W@���L��!��y7�ͺ8,�Gʤ�i���`����]�KPK�����I��7WBTz��6ޫܰ6��N)��V���Ot��y�}4N2�oqM+�������*�%P��Ҷ^��Ys��%�K����p8,ܻZrq�(���5���zvM�fP�i�{��#0���!WVdܮ���n�R��)r���E�]�m�Q(�rr�GU���z�S�Q��TV��9���X�5Pa�-"�)���ѽ,<6�a組l�p=��w8�̅񽂚�ǐ�o����nf�6�"�s:����r��ۚ5�+f��R�W�m���e�ٵ�"p�6m9ż�垫�L��)��!�1�N��٬�],�p���h/�u��Gn�+��]5f@vX��jZW�m�=m�V2P�U|m�T	�՚���l;Qs�O�9Ӟ)���y�J��z�K
��ՕmH�� t(hN��M$�Ec6�b����L�S�_n���v��8�7H{z�p��#�5զ����2�H(,n��L9��-�d���JҐ�J��tK��0]��g�+��V�|3�빎���BV�l*Z�XY㙊�=�{��F.,�9d�K繲QMv�9�`�{]��Ͼ����|>E"�Y=��-�M2מ�1"$�2��W@�Z ��ﰈC0�Ν(����^&���Z�C��1��(���� Q�PY�E�{���w0�c�i�g�2��;K릅d��5�w��u�\��I�KGqn�ش�M��],�9�������<N�i�e�e&fc��*���>��P�r�W��heo�5�W�[n.�n����+\�tz���ȏS�AxqP����*�,�}��u�2�i��t�2Ǭ�hm[�*48n#���1z��Q�f���e�˧�Fwh��N���0!,�}���;*�{l�B�XHnn]JgH=x����9	�Su�5Ul�+㡖)�����G�2�����#n7��5YS"�C�ϭJ�=}�ؼxe��[8 ���*��oP]H�),ܥ\�ᛇj�Yh��;���E�#e ��|�	{d	$�+�}�V�C��u�|�zS�a���	���c]�ت��*A�G�Ɣ؁�3zDJVU�G3J\����;�̀��1=9�Qu��] �(�ʹ/U�m�K-Ǚocv+�%҅�&m���W,˯��J�a�Jjڪ��Q+�ج�P�*((]MZ��V(�j�Km�(Y���R����p��e���������*E�mb%v%++X��F���Yv����PEW�\Qs5�
J�VQPu�Y���,T�9F ��cVZ���۩`�+[�j���EEQR��b�����C5�(�D�����U�e�
�#5���T��Ŵ*�����EUG6�v\6Җ�ը�(*[m+%J�����,X����T�PJ�-�R�Zآ$H�ڦlb�	�TE
�U�j)G2� ��D�3PX����eJ�Z�KG[-��(�Z�亭op�qo��z��_����w�n�1�(�ͽ��q�Ytr�ǩwC��z�]���;J\� h°�)s2���W���ջ�G���t�_T�p�[S}��7�~֠Њ�0-�ƩUt����
�H1����U:���7j��_r<�_e,����M �Uᎋ�w���麈n���G��Z�T�%ߪP����s�+i�]2!����*��	�W�R�<㨪뗼n����*3��&�]�[�Z�աwW���^�+.4����)IFؔ�P����NW�V��}4�y\�4NT��O*.s�un+ʼ""�{q=e�t�{�-UC�@Pw+~��eg�.�7�ix����3{��M��.�S�sbbr��&���n��ۋ�����roY�㡻��s���?@K$��lF�&��wP����`�ܔ3[w�hm�.�U�wQ,P1��Gu��W��=�+��n�b�^���T����1����nn����T�_m�S�{�7�veEe�r9G��ݨ ��Fl�����T��쨶#^u�k�*x�孤2쨺{�8}5/_L����.���2z����I��������\���u���w����_�҉�N�c7�W�}������45��ˬ�K������f�K������
�Ҙ�M����I�����z�y��z�!oO��ǔT������%l�fi��qb#}�B��-n%�N+�!3_��-�79�q\���@]�ޮ)��e��LwEnrUT�xQ���5��%GhR�{��۞.
����Ejt��+̷[2=�E�8��Ms����ǧ�DXU���wX8�{+��M$�����/*Wa��s冶b;���^^�d (�Wӹ����L���ۮ�8�,�a�`� ������i.�@��� gj�:o�t��j8�rTǝ��=��ƣiC���v紭]��ʱ�y�o�U*�[B���/�s�1ekO�h��or-ٍ�sP��,<(�A8��7�Ow�[�y��&�{n��Ҹ��{{���CM�ur/�����n8�t��'n[�u	�Р&��	95'����������N�F�����������b�VfW�4B0u���j��8y���_Zژ��w�s^_�\-���i7����^ �/
2מ�t�(��7���NƬ|Р���2Y�3�h9�fӉ�.�Զ�ni)��:���X:Zs�elƻ�&S��f�c�k}₱��w|�<ߧ�����g7`�<;S�2�3��iz�Z�����FYٷ��O-��Ѱ�p���Ë�D�h��#�.i���Q(�F���!�(��T�Y��:W��PY��=4�٤�������J���S�oN2K�H3�y�=��mH��r|9u�2\�o�+��c˱OÄ�u�U�64̮��L�S�(�Dz���y����P�x�Vw�M�4��3�j�{�)��!'��O�x	��s<��Z�Ѻz���}yDW
\If�.X:p��`��P����C�`���+ކ���Y�;N��@��:������۫y�~r,E��>LxCOǕX��Vh����.�
\�K{Y$P/���,y��C����[�@-���w��9��"�6�o���mn�E�+�rj�m6�Uf�\�q�֦���H�uP��7|ӟY��1!��Y=�)JQ����>��gOe���	˵a���f�Wa��pl����
���/g]@�6�t��N0��R*�[L��1�����qY��P�i+��(/��M͹z�{�Ȼek��ϗ���;F����'s{��S����\�,l���Ӻ��_T[2�"�k�ٻ�n+E��"���������t�䗊����Q�$+Ƕw�����ң5��\�M�(��U��Y��!^.�܂���%^�Q*>�?^O����o!�ϸ`��`ʳz>!õ:��ؖ���<fD�o�h%��N��}]=\�̝�n��GR���$�F��������#P�"����-Tf�0�9�.w56��0�Qn�K1�F 9��]:P:����:���@��{\4�w���O��ݛMW������a?�Ù��W5���tGP�ߞ�z�D�tE��u��(D�q]�r�,�+%���݂����/+�;�Y��l8�#qR[�c�)Է�2�����։�ґ�ڏPB��pę�b@ԣ���� ���������X�'R���*{O����|��'�?V�A��@I�BK��zz7���M�~v|��	o��~������'�k����x�Ç;ѭP�����I��8��Ĩ�j+��o^F���@�r�;��w�ދ�p3�e��q��P<S���V�Ԟ��ﷷ��j��.���R�;�����yGv��=��ϩ����F|Gs�UyuA�N�/���/��?<�g<�i��������b��Q c�GyTv��F��R��3�*Qv�F��zk:��W��j��CV+$��E���҅���z��`��*Ov�DC��c�=۬J�i�G��B�ׇvvV�5��a�]lo��B^Z�什�VI��6�Vr��d��`�҆b���0�4�y(q7��y%���)�݈w(���Yn�nd�n���'1��i�ױ7��c7���[�ې�t��~�6j��=Ll��}ǯҘ����`E�oAu��⺂�	�]/#������P�{�#׭�kw��Ҫ�&ʙ}�z�g�y5���5���3aG"��9��X+2��gh��s�p�:���c(h�]az�����_�e�2�v/U��6���O����V�[˄S���V��6<^[���\Z�9���oR����ۋz�.��; �^���ԉ��l�f�k5�뉅�e�6�y��:�ѓ->���ʹVqcA�Dv;\���ogW�;��Y^���S�v�\�̭���S$���hl]}8{�Y{�P�p*
���e�z����=�8v9���(��#mѳ��֘"Z����[S˭ÓVlx�FV�ވ��02�;���-�f�4�\�6Ԝ6�����Y��:�ϗ�����<�a���Tٴ�[2bs²f߆����~�3(7�q5�U�K�7S�l+_/g�f�TzC�`W/�;�	�;�%�m������Ls�ݑ��Ɲ��������ڎ ��N�B8�;S�.o}Y3}~7�
m�b�C�$�$~��S�Er�~}YT��#����Py��3{�Z�+���l����c�B�3�C�Gow��X��x��2:&�tTw\.���8ᶽ���������1^�ޕ�EՅ"W����)�_h7�h��hj��'A�A�l�'Vbዞ׌�Њ��-gj��qns�j��n�:�9���2�Չv��%
�k3o{R�T��0�D:�-��K8�rv�O���	�Ot�n�ml�h���2�9�֎53v�~�C�N��Q��홷�(&F�.:��m�h�����٪�Jic̷�8�ҍ8�I='��X]�Z�;��Es/��2|��}�C��uУU�L�kZԅ�O@܀q;�����E~�Rx���ʹ
<�����6v��\rk__=�T��A[�BoF��&�x.v�:f��S*�3��4�u� QtB�-�7t�y���nt��N�����)؎�-gn�yj�܎g1z��B�w�+ƫ)���7w�l'^��Ʃ��(�\�W���W����J�e�[C��Ń�S�����5[/*žʁq���}�
��\(�����tهW���׍���ƞK4=ꑻUsܨ7�������x�݈�u�n�*)T[�^�R��fZ��8I�1�:
	ga��[KWb�DK�����i�yǍ�Ƿ-�PIDf�!7���ZS�+E�B)��\��Ѿ�qq�dP����m<��H�T���>�"���joln��5Y�<b�_J�W���u�:�F3D)��� �ɩ����Vߝ<o������^�<i�M�xb���e�>�Gz��e*��f���ǲ��-����s��:��+7*�V�غ{M:��b����ڰ`��	�)��=�T������u��V�ס���uRPaT,����W#8�9W�.�8�_9ؽg{��1&�7���z����`�:�<��ҭ��M�#��3X+�^nz�~Ѿԓ����Պ�qGw��>�U����.�����{��>��y���r�D���w�z蜠�0�[��އ:�ںh&�W!`�EEp]��(N��������0(��Z�1Mr���Ա9�_#ws	���ٶA3nε��W��I{V����L0��� ��a̠d��e��{���Î��8��W��*�v=�w�����k�8��V����ֻ0v%S	�J}�3#+kV��zwt����W�:��2�h��=�b��bW76�Z�̤�<W04�5ޓ�*����f	A�7��ٳ{��fm��2�mT�`���捪�7u�!��G��:9u�䵄���)P5���-��;�8��ʝD���q�j�5I����M����Ǥ���v�OX:�ֲ��n�p��¼<D�.����Wv$������3��,g���m�f���ށ�׮C�M��6�]��o&�5���q�����VRHs�s���z�Xn�x��KU ĉx���{pM��d��6P����]��i�ɫw�����h\d�t�l��O����Ss���8�U�zK�Uw!�s7�1�NY��-25�귷ɂʘ����m/|?��>
��Q��Y�괁$~o
�d��w`�;v�g7�R��y¤'��\k�X��dB����g�I��
�[���t��m�^�;��,������ۊ��6�%4�ࡣ�[fb�wx���\���tIA�/�% u<��]ލaJ�[��B�n�s���f�kIcݶ��嬈>�v�F	�*��ɮ����Lce����.@�mĲ��I���H�|!t�)�v�ڕ���Q�kf�g(7XՎh�º���V1k��h��M���(�l<���њ��XGN�Nӧ�(�ȝD"�4Nw�n�Գ)����MZ����K�e��u��=ui`�+:��phrtw0V�W��ڰE�=b��/vd*vх�e�t����+�6l�?�����x[����r���
&�����2�9"�ei�E\��s�����Nv�4����Z��['i`�z�G_ar�L;v�8��:;��*�\03E��wgn�tXk�2�_d�#����]�՟LϞ�� *&J�GZ�ҥJm�2"��F������+K�-�Q5)��MJDEE��UT[f�R�Z�J�V��)�
*��AA�ڨ�"�D�ʗc)�U�E�%cim)��mh��U��UUEEE"�1�եD�,Q�����2�ԩ*6.��[4Gm�*���5����*�5��J��ʠ�UUKKl��楶�X���Vҵ�+��i]f�֭֮---�������2�l밴j�6ڔR*֖m�]p�8���mA�sfmj���kb�ֻ-ԥ������[hUV�U��m��R�mp֎t�
�+A�RщV��LZ-���l-��UMh��ۢ�f���*-��Q$�Š[)���E���h�{��ɷJ,��	�����m��'B��1#�5��0����za�[�2z����k=<5�һ���\�t�*�?�'�,5Tx]@�R��ut��V�CY�n���9��3�)�ҹ|{�\\G1�Q���NC�ޘ�֯�Ǿ��������B�R�Saө������� 0aK�"��-vT�K�a��MTطլm�n�,.�����Y�ӭ��\���������z���uL�%<bSDRQw�ψ^� 5��X����)0�+�*�z�$��2��{���9�N���E�Q�w;�vU2z�ދUTj�6�e�a�R�|R�R
uz+�Ѻʀ�*++�bi��ӎ��e��f�����`~�O��p�hJ���#�I�Rӻ�)�KAy���%>��X�v���.��2��^V5(��⫂�B�_K`a�;�NFTNŤI�7x�fPy�ˎkhM��rr�nqʸm3n'8"�&�\���������^��oq��zWU�W��}I���>�"(�p�\s�y��Ց{&j���s���������+7��>���mm@�Agc�1k�ej�ɑ��n�l2�*�9ǉ��<����e�jC�O;�}���I�sU�]����i�,��g�9-\�w�錁)u ��ׇ�b��w�x���f+��w����!�T��ܹF��a���b^UO;[Mi�UO�,�m�6E��/ۄ�?n~ȞJ�| ��}Z��(f�¸��eI~;[�IPS|amN칱˥.R-������u],ŏU���=Άt��!���q~��nL�r����d��2��~VS]�hZ0�oU�׺y���EV�_���.�`*�Q�-��ck�]�4`ѹC����Ndm�r�m^3� ������ZB)�8�wD�]c���!��n����	�U��EA��ƅ���� �Z��ʘ�����i7�`S=Xxbu��S9N�GB��wƵRǊ?<q�)�[���z�Zq��~�5bpW��עk�-���p{ ��ϕ�	�:����߯�D��Cf����ϖ�r��`u��K����Uٛy�����������>����k�V=`�rSKe���(�Oν.�75�m����}.����.AF����DV�*o���5�ڡ�sn���Ճ;�g��sY��[,�O+���	-*3�n�W9O��czt�@�E�=����|����&؇c~9�}ޢ9�jګ�O5^��l�u���G;������u�m�27�a%곏}.��*��!���GXM��lv�g��o"yEN���v�t�������T�j�qp���!N^Nc����ǡSفL���-��z:L�����
����!$�4B��3�Q��P��νR�
��݊v�u'�=5OZ{�w�U��l����Γ�v2f;��NkuWA�bz�$��Kzu1l�.v72~�:�����~]@?k��MYW~�ؖ�K��Fo����T��������,�����^����E��M�h���W9ا[�'Ssj<7����|2򡅩��J9P�'i���
����5=��+�Vk��J.ڛ۪�N��[���$^�i��s���M<�+L�bjb�r�]�X��|�㟡:C�8������|�	Ͼ��'�;eC�hL��7I'������݆�?G����������>���r�=gR�8N��'VN����I�����0���z��T=�O�>�{tG��z#g���W�	��>��O�d�k+���G�	ZF��b����ɸ���������tG��5l��h�e����^�ٔ8�/�7E�J��0�J��B-��GKn�#F�J9͝g��}�d���p���6�B�����ư��ē�V�Y'IY���	��̝��|���|ÿ�'i<C�|�}�\������c�U�|���2���F�{�����Hx�8Ğ08�Rx�I��9O�[<H
i�PY&8���OPY9��'̩���'�9���m��wǿy�^n=8d�0�ӦO^XO��$��VOO_�q���C�T'hq>�'�'&���9C�I�=d�+���>w~����|��}��\�L��NYS�����S��I�N���I�>I��'���O�hO�C�TOl������3�yLC�1�Ҋ}}�}�se�Ч��S�O�X�<d��ud<Bc�|��O�����xPY?O,I�c�4'��,���~��>���}�����~����}���O�l;N'�&��'�N�z�}�N�����I�7t%ϣ܄{�1��W��LǢ/g*��������W��PP�3�+'H,>-$�'l��$�'���'���Y>zd9�=I?!�C��w��^�;g�L�|>J���O)Ǽ��T�臇ވ�b�P��dY?%d���'l��?5$���LuOY'��9Ԃ�G���������S�Sg���{�">�f<��	�yB|�L��Ad�!ל�+$ǔ�d�+'�z�ާXOsa��D�L����v���%9{�;yE�,>��>d����O�9���N�Y�!��yŀx��,�*I���¤RdD"��-J��� �;������{�}W�򫍍�t�y�
L:,ٛ��[�mb�F�ᮏ'E�T�zD�M����p"������E1�]��\%c��-1]P8Wl,q�W���f����E�7���f7��N�ē�>��/l��)���I��2OS���t*2~Ag�)<�d�ĝ�}i+$����d���7���%_�[_of�;���1�\��"<�ފ�������C��IR��|��=I�
C���2~J�ć�9I���8b=
�|��ܽ��������O�z=�l=d�<�>О���'�;`p��p�8C���IS�i�'�'�Dd���0'�7o9�^NV�������<�I�'>Y�I�,'�����ԇ�&8�I�	�NO�C2v��叾����~? ,�~^�¯�W_�����?2t����p~a�'l�y`~I4�x$9I��'i��	��H'���C�N,2OP8>�t���������L��~��������B"�̏���z��	���z��'o䟹�?$��1'�Ni<j������'IS��|V�~��n��?z/́�}�@}Ր���Vq�	�O��x�������	��oRN�9���$��q�>`tǦ}S��\���?f�v)ў�v����y�;��!�$�q}C�Oz��̞�g?��7vy��<a�{@���4���N|�x�6���{��5�&�if��&g�0'��|�{�}�1D$�ِ��v���OR�9I��<a�VC�Cwg�P�����N�,�s���jKZ�yIr�'�G��}�b=��ql�O�,0ZC�;d�953 x�j�����a�'l�P��O����9���ُyO��;�3EꚎ��v5�!^�o���soj[;ʸ��m�cѢ���&nr�FT+�p���~��r�Z�2L�ی��)�k1,ĒLˏ}�^I������_�=�����bRt.>��s@�UN���?g���t�Ƕ$�;�J�pyg�T�����O>J2N�<N��� KC�}����+2�]}����^����c��y���'�}�~I2M��	_N��;�<C�(O����V��<NLXC�߹���'�������}�_{y�]{!˒',��h|kԓ�t�	���=NL�� ̛�0)'�q�:J�`����|���P<a��)��_*�7�i}F��{g�}z#�wH/,��ϙ'o�T	�O�z����I�?wBz�L�qAd{����W����#�s׿��~�䕓0��t���|XO�ä��8�^���E�����I��p��I��bǶb&|�""�ޭi����W��wع�����8I��bVVC�"����ē�q݁�z���/I'�|�v����$��o, �zǬ� �=�����B7�Ns}�����D?}�>����2q�8�;��x�O?RO�P;B<��C�Cqa�Ĝ}`r�!8���
D��E�c�1�]�ꘉ�l��d�v��I���~I�'iXtyHz��'���8���@7���öI��O��1��yL{�#]��現�G�ZNP^N��S�w֞$�����:I�'�N���O̜O��'������}Bv����L�<�x��o���}u�u��:a>➧�2�~CĜ}A|?R�74�8d����i�OYYOh2~$����$��1'�Y<m��z�3b���4��9K�~tlmi��S�`�Z]W	����;��Q��l&�Pv��<��bPo4q��ِκ��x'����Mu�٫�s6��c]��ɠ�b �T�G�:y�]:�����ѦfΉ-�,�m��H4�*M���/��eW���2��$.��� �s���|�'�	�Xx��Hw�2}��t}�=I;$�H|�����{�s�}������'���"����)��=`
n�>AI7�z����;I�'�S���2Ø��>��}��G��S��q;�v~����y�$��2�;d���Hn�:J����I�x��I�&a�
I�x��V?$���=��x��~s��xi�?`[��ܢ�\�����=����RO^�9<���P��%d������z��V��ְ�8d����˯����W*��tń���?}����\g�YP�'�'��y����ڲNY?Oi��i�Ho��
��-$)�s�}1d{���9�v	���>a��������a�'�l�%��I��$�[�>0���;�<a*pwa?'��,��J���S�+'���>/ 1~�g�o���#�<g�ُ�{�>�>����psB}͐X�L:��&��<}B�4�'�L��'���=b>����=x����X�𘉘�|ǽ3�T��O;N����q9��Y'���C���$��¤�]?��	��ϼ�.}�x��2�:�[��K���}�8@�|i*T�O״�'l���z��'Ć��'�8�R�!�6x�=a��'��u�?{�|������>|���(C��*2r�ϧt'�~d��t�qd�RO�N��?jOO���^(g��2�<����|���7q��$V��;ڛ�u�(gi�7;����,�*]m����� ��s
g��W{_�	��zp�~�=d4��򰮡��)6\w]���}MnH�Xu��+G:n	��Ǎ
$CeK��9���jc�]��^���2J��@��y�3'����?2s�!�O̜�'�<��P�O��8��\�~�;d:��B�|�q��7��U}r�=��D\�ϡ�s~H
�x��*i�x�����$�$����$���,�j}�<���}=�e֞�>߹V蹏O��}�$2t��O�tw`t�2xÞ�'H|��� ��z��T'3�t��䝲�״�M����y��s�<���_������/�Y�!�~a=02N�����	��L� t��2v��u@:C�8�ϘL��=d�*����{tG��H2�������E�{�u�����ְ���'��g̓�����	��̝��|���|ÿ�'i<C�}1S�{'̾�+�?����B��O���u�;I?uI��$<w�bO�Rx�I�')��g�O���o�>g��L��1S�|&5ּDJ?\�V����<I��i�$��|���	���$���x�|��C�2�;C�C�̟'f���8懨,������y�G]n8����q�?%`}�'�<I�*s:��n���$�v��$���=yd��$��	�!�hrʀol��������s��_{�V}�T�\��FO�!?sC�OR�8:�>d��d<Bp�=2P�ށ��	ׅ ����:M��C������>��~��O�,>-��2v��z��ᇉ�'����'��c���E�����[H��&{�E�-_����W_� ���+�C&��h�הe[��>AP�}���cY�8��.��gs9�[�~�ɛ@Rz[�X޾����"9�^g.�.��w�\�#���QQJ�T���˒����G�g�9��_ŗY\l�ՙ�Kܙ���P��**��].���٫r&:���t)����z�~B���ǁ�xl�3U��M���k��]�a}��P�T�OM����9����;��ܦ�"�|a�N��H�j����2!)��L6 ����oV�'��s��O�u�|��O�cH[�c�������%��F:����"/R�i�׹�l�Jn�K'��M*�*�_]��UW�I#���F���k�gh��vm������g���H��]a͎����M��;:��-W@�d�zϦ��#��Y�Ec�xH��]l������Tg$�<��`�]7�L���DW}"#��~��`��q��Ī۷��{5���HN�]]I���e�zL!7���o1Yb=��xݕՊ[�Ky
�TT��a+��6�PICk��.�2�[u'�l�e��������q���j�з|г��w^�����=Z8V��I�S2���#t7uz�ȅ����
�l�T2m��k��x,3�E�����D��*���_sD
��oE��s����u��n�5��]Zj�I*�fvE�B���P����q��]��[z]]�V�iL�������9�,�#��6�&q�Fۊ��v�r�9�� ���S�=骽���$�zF�pJ��{R-��+��bw��
�q7��ӮV6���Z㵂\ɚm�1䛱���vi@�^h�S�h�$��oJܺ��[��tz��R�>��Ԇ��*�GYi�QW_|�p�uPAޓ���f��L�ך��{8*�.e��;tv,v%��rf�Ӽ�;m��ctA��+z�w]�-���[5�,ڷ3��o7N�0���:{@+�3w��(hf#�]�uq�8��6�aߺ�<�R���Nj1���Ejp'�c���KNV�xV��;µ-ȹ,�4_4�챎�0{�����~ب�����x��?\~�8<v't��sub�f`��}��.��8�2k�P˸�KNN���K�R'���`�թ-��������`�ʈu��Q@6��6�:��,��o>�ž���X���g���c��o#�[Yɵ��J��޶n������`C��������l���S�և)WiW�+�J�:�Ӱ�/������P0j���'2���b�u�pT�Ղ��*�� �-��(��r��Ȣ��M����b7�D6�38Ќ^�'E�Sj�Gz���:�aY�k�2K���s��q *K4�z�d�-f�,!r�44�q�H�Än؄�� ��K~�8�T볨+*�Us�e�w֑�:��mq�a|4��SfY��+�5�1mɀ]̫��W���Q��:�!��xL��چ�3�j���i�5�ZK��j[�;��U1⹹�_�G;��� 3���]+�A�nK�u6�nn�/�L�.0����{c2���Re��a�<X���<��L㙕��j��3syן����@]�� ��D AZX1Um����ʹf���m�KGYn5s�֍��k6,���Z��fM[�T���(��d��Z����Rڙ�U2a&�[M��emJ*�W.M���aG]t�e���)V,֭�%��ef�]cJ���\5��ݲ1���R�ZV��F �5ŵU�J���T��mfv�d��3ElQ1��Kj���[mJf���fJf���Ժ�QF6�:�����1��*�Db����X�52��(��UTE*�lQ\�b�m�(�Z+Z�U+uBĮL9*":��m��Tkm��g1a�iB�ָ�1*Y[���m��Uu�4fs�[f�Q��lsD��4��m-V�j9�ڹs��a2G%qm�W�i�o����/+=�S�v�˭UB�#qWi�q�qİN'V_:���8]^�j6Ӊu�}U�r>~��ܿ��5V��ǚ;;�d}�Ҿ��GB����i���=���d��܇��%=��uhv
�r/�yx)�<m�[���)�G�~���8L^E�%.橀�l?'
t���LLtO53��M�w�$i�W�B�i���jq�f:,i�Ԩ1<�ޭ��'6zCE�|�e*qV<��Ts���k-_I~�rvS��-��9=ӹ��Cj��W���q�c�C�|C�Sկ7�X4[��(�K]�]m��g��ȧ��",WV.o�p��o�f�":.�SWt��1�v���!�}�'���Us;e<�"���z>���X����3�ʣ�wp�fΫ��R7Y� ݲ2.��-��S�9�ۧ0m	�9���OT��d��v~��4��7h�Y~ࢤ����w�d��d�{��F�E��U}��^��T�?��������)�����'��p�<���^�Vߙ��X~;G��:2�4���0W^5�Q;��(1Tҍ���<X<!����,�Q��)�����׍:����=��tb�g%4��\<�����f^e^w�f]
��`�o�Dg.B�7��ܕ�BLN���s�)�#0�t����9��g��嚓m�M���or�;���<X��5�Py��k�6Y��ݭt�T����lOv����۱�����O����sv�[���p/ܘ������Ҹ����5[ͮ���7]�[��g�U	���f��-���"��V?W/�g�q_���Xۃ���j~ȄƉ���Xx=-�Tkj\�a��G�^�'��'=��e��zD�W��7����ȂWp$z�`��z�F�9ϕ�������6"P���{VU�_�ވ���������w��o��T�W��)�*M�2�s޳�}�B0a�� [���)v�Q��<�PBMP���u�2��Yw�%�˿{2?Ej="+���6zMrϞ�ka�Q v���W�^�z�C�X4�5�ה=�h��1�wߩ�����<���\+�Ӛu��E+�ܭ�z�^n��L:$^����Yh��[�"
	�*�0\����Uv�7m9���ڽ2����j�dr%�}ާG>Hm_����*�]��m)w+��׊&���`��}����F�L^�اi�oB:�C�v��Ir�B��n��e�#��4㢽@�����Ͽ~�l�M���_���vާl�+�:��� u��[��ݨyZ�f�gI�v��n�Ӯ&̓��i+T�B��O���͙�]���=���[��t�BVx	�*+|O�}�}U#{9�wu?�4�}��c}�9�#.t�.u�ȹ�1���N���V�7F�ے%���}����掭�h3�S��	��O{��([�G��M���.�j����x��VW�}�[�P@��W�y�����0Â�S�ť}��j{�6�\�t�9�`F���i㗶�i���V�Ҽ��ȷ����_��C�7�aYs�֊ �bF]+�x��S��������P��wOL�{�ٹ��ƩUt�\=����4R����y%�׼�V,���i^@�W^�b*Uxz;�\o_ʏ"��7gj�僤5R��L����
J�O_�@�y�[��\r�j����S8�R�^��/@�%-o%��d�2����^�1��D�G��6��7S*�0'�ٛ(htq�*��j��=��	�*ƾ��v⒴�3���_W����Zy'�u�Y�x�CB�LU"��#�o�����/x{ ��ϕ�]���h�mՍH�$���^�=�Ci�;�x�ٯ��/����=��^@K���+��:>S4/6���Q����(�V!�ݾ�Xoe���+�ܛ�cx��.[C��g&�6��x�3�&V��|��ͽQ���k`�3ڌ׭�S�4�f���pV�;������F�
ni��=L�շN�O5P��/��
טؘ�=Of���G�Ae�.|�t��Z�>�W藃A㐆6�s��ծ[8ϖ�d��M� ���8�'z��%�目_p�x1�̻��E�����QfM����d�(�[���/��4�+�������\(�Ygx�u��'M\.p7�����>��N�BU�A{slQ�Ig�{��@���'_��~�l�fz��x��J���L���sݫs�ց"\};~*z(��=���q^�b�9�y&�3}�"|����\���JC�Lh��dU�K��Mͨq�#�{S7��{�o���֙�fx�Mk�����>r���
����ϫ��x���-M���^[����{ͫy+��}e���*UC=]�5�WXVrk	p�K�V�o��� h�i�8�\~�X��&8����� l���Eb�{9)�X�-�l�6�Ų�m�7g~�pX��<O�i�x�&�Eè�s�\�z/7�]&'`>����9����}��X����Y�K�u��i�����^-�4�Ґ��U��W.����r��?N.Lܡp�M�u1IΝd���XU���U��	����]E`7"����FZS��^r�=�z$�n�I�������w-{nx�@�Y�5Q�|���Dǈ��i�՟s�:��Z�\V��ōs3$��ʍp�rm:������%���.�fR�Z
�}���Q�FL>���1�c|�{if��l`C�D�(v�U�<f˩�=j;��q��m��������T��\�ky\�>3 kPy���Ca-��ew�������Iǝ�*��dwN̦g��躜In���#�c����¹B���5)v�?b��mncS��;��>��w<:j���1si{�� x�(c���i�L��oD�E�QM<��vU?�7�m_,RW�[S{��3����f܏9�t�-C}�T��ãj�3���\����H�i�Q=b��k���9ˮٖ�nwI/��k�q��`l���;/����MI����}��rk�唵o�G�#ª�Zn�Nޅ�Q�4�vʨ�E��NR����b�0P��������z�[fSθ6L]����[��.�o��=��~x��	�E3��V�7
���j�ar� ��}��b�$�y��#��4㢡���+����]ŷDvEfˋ}'{�[��:6��8�O��#�/^_�})��ü4&>�Y�^WB���3̌�X��r��%�dy��hy�|@O{HW��Uy˖L,�1�"V���G����b�������]���4��h��{\ƽ�oRu
�b[�ZYt������Х��.3g{&��d}3���\�P5-2]��1�9Z�U]����oJQ�M�C��H	`��'N�3:aN����"�a�e^X���=�f󈕝Wȷ��vl+��e�N$l�3���j^�lE��5}���W�Dz=ikp�<�����7�6�:F��wOIF�5�gb<+��x�ѫggb��Wӧ�u���ITȤ�EH�y��$�8�=�D�{
�5�xz;�\o��"�|�s���K't��KP���@���?9���gp��-�����;}���zF�=��D�hx��	A����Z���"F�mbپ��b��3ɫ��/"o[E��ݲj���
w��uf=�X"���\[����:y<I�4Ȩ4B�u�oq~��:ټ�Ҽ����N`}��6��=\'�(i=/�
����yfj.+�*�<M\�t[4LM�q~:�E�SX�����V�*~ЫF}}���q������+~�5UbK�u&!y��_W@�U�Y��8���5�wq�e��|��x4����U؎+���)�:�� �Jz�� �{�4v
ɾ�Z��[��z=�'�&�Z�h��jY�`@�P^�9��ָ�5S���Y�N.��ru��yKq�tW���w�W��j���L����3S����z$�+ݏ"[�aA�sM�}�}_;B6��/��o�)�ݦa)nxKޗs���UcFLk9*�F���ĕ
���!��M-��,
\%9&��^7�����}�����ݡ~�]��Y9�Z'�^�8J��HA�z���C����p�w>u�j���&���]1���qZ�}؉3-������z���C6�,'���2�$s�|���HqNlH�j��{<�r��:�����!��˻���:"����B�J�Kf�8�&i�wx�=o� "�SPN�fT��������mR�Ֆ����/CO��>.��],�Ʉ�u��`RR֎����/.i�h,��Ż2���p��m,�T���|�j�{�~�u]W[�EYt��ː�cr<Í=9qԬfc/+D�*u���*ţʭfp�t�7І4��d ��s�Ʈu��R>T�pjMe�[�u�W�B��X�[{+/��wu.G��ʍ���7W�XO�("��/��1g�y"��l�X���=�Iw��W+A� ]�@\��9����̾ff=���&���Ex�0B8zI�%d@Ay�Ac]!*������i�� :�֋6@X¾)�чn�w��g���v����}Ja�0�,�d��ی�E<V{x���4q e=gF�	pJ�%NaV��![f����t�/i��X~��>��k��gB�{4�[�Z���*����X�`��=��ˎ�����f��ٷ(
���FE�}Z[����lVU��y���X�m�ʈX4��@�ͱ�#ϞS(^b��yQ���n�X�
C0��D���l
m�T=�F�����W�$�:��7��M��m�\+I���E��u�ٍRJ��WY�f�!��B�ޥ����[��Zje]�4���Δ�츍�n<���0Ix6�����+��n�34��b��I��9w�p�p��=Prnup�9��8�Ȧt�7''*��օP{/y�y5�53W�m*4�-$]�_�yB�H���X�,�;l�c�b�m��R�u�r*���&�Eh��KDq��
��C�q��3�"���ѹ�^���+U������O��E��Xu͎u�̂���s���X����[a��zNf:��`V)u�]�]l�6���Ϡ9�+�^��hVWI��wQ����{���RX�$��C��W
 sk�//7�z;��tsn���Þs=�
0[���iu�wa���y�3�*���K��"�l����#޽Y{��-h�77{*t�Xt��=�-���������6nt#p���X�τ��[��ntl'zJ��۾�����H!|MK+Z"�V�uv٢��)�Lͬ��n�ȬETTR��j��m�����[Z���GS**�L�2W-�(�(��K���Tj�h�5Ĭ��2mJҥf�iYQJ��b6���TYmba.v(�LZ���ݰ""*g&�iKn�1��h�nM����j�[V�U�ժ��f�֢����V�6�Y��͵V�Trdأmh�m�-�L�"��l��f���\ͩ�Q
��
ai��stKf�+(��n.t�kEXQ�.ȋ2e���(��ճa�������շjjks�ȵ�7�ը��sQ���m����-UZWSR�⋒��E�UŵF�D͎��.�]]FQJ[m5��Z���l���V戭j�l�K��rж�jݭTΊ檈�WZ�m��eaDj6�Z�ŕ&$��{��v~���':��mJ�DV�v�\�U�G��.��멀O����w��1>��Q ���ꪯ��	Q�q�s����z:S>nm��%�ufa�+@�����ԝ���X;G�1��L�^��侨|N{��׫��R9�y?��%Véˑob��u���B�dh��[|.��}�yz4L��'{�{�\�-FWR�ڍuƇET$�;����7��	��u�����qK�@���;�k�@ɪZ��\� Nh��w���98���~�/G�<���%t�"�Wk�R���3S��3eq����x�g1;(�aCz
+�7^��X������7��^�ǔ��^�μ.��n{�R��	c������-�<y�K����Sa^G���v����A�v�l�{�q��Y�}�`�ʪ�AS�6�v��<�w�q�Q%�*�ç&��r��څ���sf>r�M�J#�nXs6�L�,�tȇ��Q�y������ ��}_}�}���)��7L����/UG	��;'�08�����.zqM4��;ȧ����кUF����*�q�`/���M"�T��m���{1N���wnw���^��
���]�s�k��8���l؉21��ԩE�z$^����Q7�]�[ԛ������D�U"���Uv�p6ӛf��۳�5�Nś�qv-��ڹ�ƍ�*6�0����]�n�\�Ř��lV�7r�on������9����=w[��u��x��U⻦�3=&����ˮM:!��Ⱦs��{�Cwm��ds�uˍ:r��W͡d����<S���V��f�k�_/߶�J5��Oy�ܸ��!�qo^X�m>����oqF��˴��g=�*=��"f^VXܽZ�#);�`j9;;��1������S4�ѣ�5v.��/�6�:(s�+x�aU��IpIq��UU��Uǹ���m��l���u�{�ɷ�W���j���I5�N����q��teD����ns��Z�[��j�Ms��Sst3��>��0<Ԩ1:��y>��˨YDeG��ӽ�6�7��I�\f:������U�d�{�R��N+,�vOf��T�b�|f����l�����5�X&��b*�{���W;��qZ����*@�n��wϖ2�)�-�&kvEBj�tlwJ�y�I�� �Թ���G�5��o$�T�J�w��"�6�6�غ���&���GL��q�6�d���;�HJ5����W�y��7b,ڨء,�#o�������!Y��8ҽ%n���O�.��v#��~�q�ٷ��A�.<�]�>#n� �p�i���I��2}�Ͳ�Ci��]e�v��D�-tu�.iH�(�6§��dϫ꯾�rS�{q1���w����'�T'O -��v����3������Y��]LzWQkٽE�t3��4�w�+�J:`��<����gjȽOU�Q�4��~�^�G���y��vf�DV��.oܛ�3,��{-�U�{���@^E�Uxv��1�A��=���t⒝����o͔x(^.�u�nK�3ںhޑ½�>`A���-V���sA�o$�'�..'�I�i5WQ��h�u�z[�q��S���xi�ڠ��kkG˟&p\�W�F��t��푢/;��B��yJt?	b�k�����u�M��V�91G��*F�~���� ��~LܙUhc
Ȫ����t��d4a�g �3� �v),�V[��{yZ]@E��C�D�+�K�����n�n%etr�\xF��N��:5��Am*+��#S��   �;s{��p͟�@���N3��]P=t3�w9j��;ŵ�=s}ޖ�s\OV��p�{�@r(p���q��(h2���=sz�G�����ӆ����&��k�tC���W�`{H�ԕ���~�#)���7�bb�M�6�5���	�-*���*��m�K��	�ķ]� �����:)biY�g��:3*����.�CS���%//E��e�=+)��|qtd=}���)�0C�ܵ7�����x��"�B�������M�Y��݋����l�M���G�ny�X�5{/짘�f��䘬n��犸i��o-o�����-�d
��>��>ҍH�O��H@��%����/��9���+�Ǧ������ʜ^4		n>��P\4��)��V^�p����s[RqGiQ�N���F��@
%m�%55	������Rq�\�}ᇨ=����/���%��o]��?fs��?OY��q��{^Z�U+�P<�+�yRa���]n���0=�z3^xG3ʵ�
���������=�6_���1Q��[<���k%�c5ڄ���^,��	�����T�3�;2�����Yv��R��u2��4wJ��Շ��T�Q�J�Z��e�*��ޫJ/CR���纭h�=]�
��5��X1�u������]��%���z�W�y2]���k;��=���N7#�;𷵶U��n.��T��FRi%������ڡI�L��bSγd�7���Dn�����Ď����"Ã,^��S/��.�"�8e]�_�1���MI岁����yM������L��~C0Sڝ +ᣬޗ����j�<��|�[5Yt�XB(JU|�R��z#ވ׻�����V��}4�����=�����=��{�4��v��{6�8�n�7O�ͻ<QJDr�;��Y��a��a�Sz��%�m���`��n7z�֬��2��eP|i�NN�OE��yա��V5�;uժ�u8�Q��Z�u�]&�]E�w�����6n��Ş�ӆc}�\�L��-w����'މ���nv����]�T��γ5��&�B�Wm���\�Z���nd8_M}u��y���w���^�s��j�E?�1��exp�J��U	�1��pڿ��Mo�3w�(�k�&����=>�+�*3ڭ�G9�Ws�7p����쑆ڡO6^��\�U���6tT>��2mY�I�a:/fʅQ���6�6Z}�,�h�&��}]b�l�fEmP3�itZvW4h<܉�"3�����DV��o'F��S�����o��*5x:T��(�O�e����+�>��J>7�oh�u�1���Tlg7�f�Z�276�MG;*��=�}<i�/���{�P�Y���e����$F_:k�L*��nA�ؖ�����ǋ�=[]�g���}	��U��wt����՞�[���ҋ+���@�F�T�R�[�
3��>n���Φ��Mb�
3�ˉ���Y3�v��oE�� ��b�_A����Me=�ڜН��4櫲�Uw^�:�v �P^��sf1�l"�7��Yb����@XuC�WκܝY��?��h~��׻^=XvVY6i��,u.�%p9M*ͥbP�Y��p}ܹ�aep�s��y�F�]��N�W�稺���B͖��z*�HY��c�un4s������FZ�7�U}�W�[�����y��}��<ZZq&���,�.W�%y��H؛��6�QΕ���yI�'�Ϫ���Kb|��i��]B;<iى�>"�ҡۻr���o�sŗ�1��%���S~;)�W�Nr��S*����K�pJ{���4���f���C�ƒB{K��>���"��3,�y�xv>����zE��ԷM;Cô�b4թ�e��J��k�(Ŝǻ�@n^n�OI6��Z�	��	�ז�7K�Zx�ed�6��+�i�GO/2nvoU�.�8}���*�W��:��1���+pqs��˙����b��;1��f܅7�����_��Q750����^����f�$`�|#_.N̚rc�ሞ?e*J��a���9W�y�=������4j>�(~����բ���M8�QY��-�SC��e�/ �˲�.}�m��t�27Vr�H����u��Q���VN7i��J9؂�7Pse�33n�
�Tq��z#��X�7��+$G�N�FB'ʋ���s^��=1`�]"ʝ���1r��u��mv�R��&_�0�E�j�Fz�7�8/i�Z�#ACd�u�ݘ��莬���Jh�s\]E��f�/��@�����O6{�֙�4��);��)��A8��<������O��k֠��U<GN2[o�Z��䌫�Ú�Cm�FF�
�x�����=3�-	A�b�7�>��Ɍ��Ì�'�M�}�#��
􄑍
_�T�^�f`�F�r~���uYe9�O��K�=.�`�v���3"n�w{R�>OQ�R�|U0"a-1106 N��OJ��r=!V�����m^]Ͼ�c�_&-�zx�=�Z�\ruBC�1�ȸ!K3L�ՊUh�{�mY�}���F�y}C���rA7K�b��9:��:�G _���_���d��?*Dn�o5->:kb��c��3�oz��8�·�j����6����h��@8{;Ml��,���0��(ׯF�Pt�ypaʴ9�.h���wnŕ��ڕò�+�y*Ð2(7�^0�n�%���$9��#QwQ�������#(�������6M9���'*���C�1VvS���R�_jxd�
�pe���r���w��PN��>���a�e�a2茈^�UtF�U��\��<����Q	@�Ճ�gp���r��Z�����۾]�����Rv*z�}ܴ^��٩m�G_	F{��^^ukY"��"%���R�ʉ�]Par�C�k���n�QU�5��7���+h]�͙��pk
�ÛC�U�P�y��q�w�yY�1���	�BԳ��;36T�{��Lօl��k�]*wK�{���xW�{�1���C��+c.~�����uP׆|��S����XQ���NvwP04�
��ōV�]t�'lwx9K��+3�ۛ�@�L@�v��Fh8�mx{/ky�1f�*]�m�cI�3%%.]��u��0�l�&�c��
�@����o�M���[���L�@UW#��g]���U��Ap�5��7�Y��Ae�%��o	�]����,�ҥ���S�R74V��_/�zۭ8�W_�
��W���˽cq _e�=�ǹu��v�O6����D��M�-JZ��2h;d.�[�	��w�L/M���&���I��Ec�\2�_MX_i#�\��ހ��b�9"亪�s�#x�/�%��[�K�����-���[��Wf�*��0�/���:��L{t��.�5�d΃y�{��:R�&����V4��;�;���fn+�<8�$��^^��yK&kM�D��I��C��ڐ�0���gC-���%�k@1��S6j��[���u+���vμ���խ{��l>����C��wwp�m�tU�
Ь�uWxGI ՚��D���D*�W>T��@[.�'p+"��:Q���t�y2���Ȋs�i��2۱�e[%����"Ӛ��B��J�9����XymL������͵�iOe^��������D�me�^n��3�l�[��DEBڒ�F�A4�IF��Z-�n��l�5R�7b��Zf��͛kM�WmqmiQڻ(���Y��&]L�\���T-��غm��h�Z�SV�5�em�*�[u6[��Z�ڗ[��D��KL.�R�i�.����W�-��,kL��k�Kv���F�7]���۵ۘm���4�*Z;l�lb�+K����ZQ����n�T�+ڙ��0*Z:�h�-�ET͵V굷�-vԫ(V�r]jU��)+
��T�ZRѺۗ�j�p���-�n�Һ���m�1�P�b�����Rҕ3�&�C(����Q��v�QԮ���M��kkK����-�dK-���h�ݝf��]#Z� �4e��mr鶸�ZZ�E��$&�|�q�~_��<5��^C�S��f���v���w���=�|C�5�j��.���� ��{{�����5�Z�Q��Z� �9�J% ��N�s�^���9����d�~FKx\��!+�/x0�X�W�9}t�1�۾�f�Ԛ��9�VE��6e4=4��H\`�W�q���Gs��`�2������ȾV_�.�O�mE���?D�R���]��U�wrrF��n�&����E�����s�XX���ט�Ι핼��^�����D�MD��u�g������������D�E�wI�U	�^:��b��D�'�p11t��/���^�1�OZ��3CxG�i}<��w]��;�F�Qx�þ�Kx��úU��C4b~.৲�<�X.2�ى�� P���zQf���:�X���'-�B�9��U��;�L
�h"��g	$�1~}����Լ׎��㥙�~?�9��V�U5�^���쵆��"AUP�|�T��#l��(�]znoapV)�}�Aq��7��V%:�웺e�Q۸�E	QN�u�ڎ��q��T�������}U�Uqa�H|I��3���n�r~��ig"V����p-,>�1���yGh%�5��P�R���װ����������:��E�Ēqf|������*�#1�Y"E�&1�[~LoS��b�s�J๼:�UU�5��bQ��&�<P��G�r�z�M�f�=x�c'[��
��m��-��Ē��h�>ZC��s�.����z5k���,���w3W�7.�:a���h��ԣ��,E)d��Ρ<.�7��s�8$:ʁ�	�H��5x��pdJ!��N��J���uZ���3�{5ptz*]
��.��bD�Ʈ.�z��u
ob�7KP�q"o���f�o�ޔ�����Ĺ<hbgD�+�//g���2x�f͚"�yFE5�׽�#^�ڧ�$/T���k���,�I�Up9�59���7�^eV�����{��Ｔ�\�M��m��,N�2Xwh�25;�V<�ŏ]�^� �a�y��@Rz��0���,c�0���Xbذwң=�V�:��lڊ�v�r�?�U_W����5���,E�1?�g��_����#hx�����ppg��q{�.I�����8��t���Y�D��z���fs�� ��Ȩmky57��}�u!O5���ַ�\XM��E�#���Rx�T�ÓѩQ�;G�`RЋ�γ��:
�C��li�O�U�$+C����Kd�|�W��|�}w��11��ڸ��M�6;(pr����3)Z>(Y ��c-��RZ|e�7���8�xF��v��v��[)KTDNp&x�.a|�6=I�2�k���I���_ef��W;L�re����ѡ��������L�0�9˅PR�>�]o+�[�g+�x�.���f-!��0�4��+�|}(I�F�k���Pt����
�7�.��+Kze7y]��}�K��(֟~6F/וY<��$����#�K ��p�V�y���&B�Al�%�f
��&�m�aCW(f�w�a�e.3H|4륃L�w_`뎦�ؠ����Ӳ�]��_^N�Q�����興�5�y��Vf?EVқ��{�ģ\���}�O,�0b1�U^��*�V-kR�(	��Ƈ&)�.h��l�pa?���u/Y��Z�kz^�{�w!�0�X��<�j��ԏ�b��\X��9;c�U_b�b���ۏʹ�Q>k��T}-ᖟ+Y-��q�e��#+ �u�OX'f1�V��^�L��g:?K��GH�L@�ؗW1j��v����Tt݇�g�&y�v!Cj�Fz�åuTK�4Fbq��+��4�7�X1�0;M��*Xҥ��K{�c��e�?���o*6�6/<m�y컽�T��i�"a�x�&"�[Vz\�{NP;j<�Q�ޱW���Hh�uy��;�M�h�;�$9$E��W��v.zr���G^h˪<�]��\`�d�޴tB���5��͛	�A�ظ���>���,,�Q��3��4�=9���4���
��V�O��|�ww���� i��חO��vC�Q��)2��6J�*o$��W�7�(K�bKX�)�SqU��W�InF�S�_UUW�H��z�����˝��յ��m�_ܵ/�ǧ�.>�O��i��9�N�7_�G��I8a�?n���o�����se�X#��D��$�Y�(7�����yj�wR��K����am�1�'��KZx��H`�H�X�>� ��OW*��h�UC����NC�\��N� �/����'TlY��cb�����8��@���_.9Z�I�B�:����m�̛])�����mߘ��#��H���v���(yW��_�9�!���،���;�U�,�3<���,;�1�(A���.vop�ar��F��w��z�5Xfv�iec9Yb��ډ�[j ��v����^��w�y��**�˯7Q�]�؛zc0Z<p���LsvƉ�����7cTtG�oA����o���Y������3"�T����~2�����>�џ?<�����ec5����nT���tev��UI�xq��V����[ۭ0����\��nm��vҔi����]2���o�.�|���k�1-�Il��ڎ-W����D
��i�T}�	/x11�i�?�Ɍצc���N�v���й�|�����V��k��B���l��3&��t��0�F���4�y��usJe�Ɇd�(0���J�u
�@N��.�[����k�C�q	Z�4.8Y�I���d��YT�f��7���wے�ޑT-�6&{�P嶸�Z��#�����by�Y�o���xwS�}��n�2�Eǃ1����}p.O3�J�9�VY7V��g�{��$��ZBjiaעʓ����*`�SM�b�s�8������������LdpO�1�Rcfl_�o��#�US��5�E�ڷ��ٹP�8���9�+ �*e��8O�jv��P�bP�I�o&N�.�"���x�4E��d�k.#���%�+WJC��-:���?�?{��_&�-x;M������|'��kg2`�=k���Myk���{�� jsz�f��޼3�+U+8֡K*��q6z�-e�V���-�%E˷s!_$'M�u�H�ʯ���w����M��"�o�N��"`��L��S��j�ڼ�1s�b�;�;�Q�#�/�1o�E��P�+>Ĩk�
u&G�ݴ�onw�.։����1.O��)��0�^�%]�<v�l��:vU�ga���Q"�^..7*����Q�vi{���d���;7�>o�U�9�±�Y��ԜT|b�e{�=M�Q�̘���y��%�O��i托���σ�=>rx���R)�U*���1\S�0��˭v�k,fX=�Le�ԇ�_b�9q�oH�����Dkw�ʷ��\Q���wǀ�
]�/��/i���}����������v�t�%�P�1o�L)0r�83���K��Ә�
r9����&rqx��ǹi5���|P�A|q!.~�_%���om3Bs����<a��6���X�x��l���l����ZCmB�����:����<6Y��(g^<���jd���Iv�3,V3#5"�Co�5 ��^�A�(ֺށM�*C�DNފ�vRI�߽�{����ēʨ��rcʈ�)��Ґ>";D; �آ6\�Q����ٳsxӣ�jؙ0��j#���0��\��bdx����in��]���T^��0����̍%t������ɀVU��7If�N����#��'�x�[�B����jDi�nd��#����ݣ��r���T�xt���%�>5�A�t��Z��eu���l����X:pA�vc����G�E^@�����Ɓ�^8�:#n��v�V6�wv��fC��N���Fͱ~b3����rb����6!��|��� �s�1[8o� {�*���IQ����nr<��Ƚ�P&��=R�n	����(vyݯ:C�a �xzzb���[��i��r oD�K�yХ�uS^�a��mV�ȡ�UC���к4�L��7]��(wy+��U�f_()�;-k��ix��s2��^s��fZTJff��`�L��u���*0�V�����7����˝�4�������ϩ��0c�۬�]��g��{�����M՛?�FD�Xzs4�CJ�ȹs\]E��f�/�K�5_gn�CF��w�gJ����B�B���c�K��{NP;�Pa�O,��U��j���Q�8P
S y�Y>op���Tt؞zi�V,'�Z4}����k���cB�H�h�{y�+q�+�1!��R�OQ�W^�Uy��݁��
0m00!i(�� ����f
�VT�{}q�4U�-y޻�C>	3�q�}���Pt9��s�`>J5��r��'���S�������5c'���c#C�9+�`�
r�H�#=UO�紺��}1&�^Q���B�񜍧\���`�n��Ʈ6J���@�ٻ��g g�E���k51���>,W0�c�b�*�U��7���Ó�U��;�c�w/�Y"C1��1_yW��̟��~�b��@Q��s;3c�C���֢�E.R�\�Z�bD�s@��j&���٧�(\��9piN�IoO���͂R�-Neh�M�G�>AE��(�FS� N_W�UX����v�f��Wt�*��e�B�,>����.vW����.���9ۣ���L��as2'��=�X�e��V�x�<��^`]e�(�����߹�3r�0�����n����}�˞[D��a��~{L�}�I�Ti.b�="�~\�-�ٯ�Y��r�b�j����aȽ�O���s
�^	q%��c��O����=:v';p�t�8��7��cY9#`r���k�<����K/aû"��f"�Qz���U���ڐ��u�d{��PH1�م���OAԽ��i9'-�Ǹ�,��yu��Rb�W�^���;:�L�a"p�j��(/� Ta����|��D\�<vks�+1��Bf�
嶠�J��?q��ӕ/�b\>��[܍�A��vzibX�~����\YJ��gf�ל��wȣ{��OO��I�V~�l���_	g��G:%�|�q}N���^[� �}�����'�"����;��BK�ݢ��N��Ȳ�o]T����
�Ar8��&˩.�u�8�䮽�v�#���k_U��[9��LK.�G�V�*�Ņf�lz�V����f�D��b�.s�]Ü�;f�W�T�톖�d��A�$�V�i�.�	�
��%�m������yY�{f�j̲�Nfd�ށy����:�V������j�ಧ*�.�}7VMvտ�*��4���|��&��
���j��S̠���1C��̀� g%\��v��vQ���w׫!��ۮ)��r�m�Iq7���]V�ӣ�Q9ì�k(W9��0�!����ԭP�g4s��FVr�����q�"(�����nWU;���g'��F;�;��.у���4�Ol�Uږ�ܗn5�+�i����Z���kC��z��o���'�ˮ>eA�g"�W���tH�Y�o�r9C�gUY�����t���xo8Z6^S��Jv�v��]ڸ�1�&k5���sq�����ۮ�����ғ�8!?Taы
~��V�*�V(�=�Hg;��j�7�uŉ:��v����UDu�Aq�C�rӫ��fWwrju�&�8�L����Q=}\���n&�7�y���p��<�C�]��
�j4����ĩ�f)��j�u�b(4�����;�z:hM���Z��j����u�eZ��{1�U��X,\�v�.R<��k���vTK�%B-�k�̡�y���4T	+���4yY�5��*�?�U�3�o�n������=��-)��|�V��u�2\��R�R��%���i.=�:�����>.���
)G�{|]�����m����g��b\�k.Q)t�o�v!MoZ*>{����ξZZ˱�N�"�积E'{y�d�gd����:p �(_�W��غ�o����껦4�6��ET��:a�q���Eb��z�i����j�AADʋV\a�"Jz�sL�\s�Va!t����ND76�YJB������wW�Ʋ�К��5��ڐ�F�U���û������OȲ�˗qL[�u�,�R�iUK7eڕ-�-ej�\�T�]L�\%��j[e�6��kn��ErR�&e���[��W\�L1�nL�EEKs�ն�\�ch�2%�8B�V��S(��e�6�b���Qfr��+k����a-����
��*6�v�ʹmm�hf�iV���J敢�[�4eUJ櫙Sl���bʮ5���˶U��j��6ں��Jm�W��F)-��*�F���G93H�Ҫ�J�((���5*QZ���L��;Q��Y��հ��	�Ԫ����Z\%����MLĵ�j�6�3
�G7R�Ah�ё[eVT��jX�Z(���2Tը�ڬ�����I�y�e�w��G�Oxh�ZO.rujc��\�`���Y�+�����r�t�M�Ŗ�IpI4'�U��[��y�C��:I'����qsō��]����5�ʱۍ��˓KZ�k'���+��С[�rI}�QP�,<F�:}�[J%�ڼ��f{�k�9��ߌ޳C�c֠�|z$��4x��4�r�2�~v1#9��L�`�=]��{u���"�Ѫ�� �q<�����|V�v^u[���T��qL����L�?t�c���(����ܯ`o�ԝ`��vaЇ;$���f0�H��\\1���X�
WX�t���~7r��
���\v~!�.N4>�Ί���*%������JU��:���JȇN#�U4zs�Q!~S��DtX���uQpGIb�v�5���ǭ�"��|r׫e�u*Q��=�&�1;�̙�rYYX�k5}6�/�E$�ج������04��D��z�?O߫[�ڒ�Gղ��H'e�1��f]�G:O�����Oc�QjzlN;+��T����X��c�Nwy���W�`�9�Rx:ͽN���%d��ٚP��/��|TO�}U_Vk�tBZ#�c)�z}��:��3��2�P�=5�:w����#��mU�ȫqU��� 7r��P�d�Օ�~΂�_��*�:FքTӛ*����A�?��C($D,��������O������1٣^V$6VfpH�a���:O��Ե$�h,h^�v��&SN1�!�rܻ�����>���>'h��̆* �HY��#�C�@��"V�M��[z�r��95`�(�v����h�%�ǒ���=y]��r�=���Y&��H��y��lb�5�&F�v�����H=������2�ާE��;i�H�a4->Ct��t/�R#L�%����<��ۻ��
Qx5�`�CJ�5���I��k��7K�U��u�%�׾�{�t�KC}�mF���3��W�'/�7��������;2�	���Ӆq*�Н>�ܺ:4�O(t����塋R�R��╭����:�D+R��:�J�h�Z�M���Ȥħm��u��NsKkxlAr��e�N�Ͼ���UL����_�aÑxلB�CP�5��[�A�5��ф+WS7��rf2Wu0.!��t�=;;X\�h�S���[������O*�׷׻\�i���L�TgRR!k9���Ys��s�<"zb�Jq0/Xů����;9�&2z_"g�3}�ηFP���T}*%����c���7D1�$�FD��\�f��4�}�s����6nr���1^
�Og7�'���#�3�A���^RXN��\��[���#��/=��Z�_v�u�>�[\�<}���# g�G��=/�7��xS<�M�\��W�08Xػ֎�
��H��
�	#�nq �ﷶ�����ݸL�(�-��-�թx����<��ۛN��v�t�OE�C䙤��7�G��l��1�X��I��Q�=H��(����֦&�ïn0�֦��m�#���c5*�Ʃmn��ζob�:v�0�kg�7YZ�k�2U�R������@��j�xё�@Q+��)��H?����	1�=�5n�wǩj^9�+.��aB����@��j�q��	��3wOW���ָ�<sVTq�$]y񃑵\��/s�Ҹе�)��osm�<��P��䉈�(�|�B:�+ϋ�a$��(LfگiGz�k���.1�ߡ;4�ʰ%�>{ɪU�-���o���ޤ�Tˬ� �U�s`nqz.�.������M�~�2�w�Z��/޹ڃ�7`�x2]y��>�.fa+/$l!�r��_�&��2�k�gm;�ڬ~3R�,�7e����t�FMv�bm��~Bλi6e,����f�{��R�q�\�>��f�Ef�x�������i��k-�w7^���"2(_
�fL7V�Q5�,kǦ����<U��]>�^Ťd��ݴs����֟W�,��͝¿����Y��DGV��P�`1�����VJ�xJKfPT~;H���\vd�"�/!���� ʅ�&:P�M��
rou��tڲ�{0��R���Ǽbɨcwաt7�J�$���}_WӘ>N?hy�I`�+O�\��I$Ą�|v�zz�:�Z�<��:���ҳ]�MLmc�m�`>�%hv`Ѕ����H����õfU<i��St0�,�s�)��l'53z����C[@��: ����f�2%�: Bܺ�SQl��ڌ.`�>��)S�l��1��2����Ìi��,���~�B7��ce?1[!LoR�%�3���W*���.6gP|z+��J7�%���F�6zn�/���7m�\����]VM�N�u�:�:�K�H�>ZC��(Ï�2�u��v�u]��G�5y']�`���$Yq0p^���^¯6{���ާ�Ͼ�ZÅ�e$�N��D���9�ƠιCbQ
ꪢe̪��{�,D�{'��q�ڰD<���0$�bW�O︌�|}z��v�ȾK?v�f� �r����>�V���"�b���-�(�ݗ��;�vw�e_;��e8]��3(�l���ƛҸ�2	R�L�v��:��YV���m02l��POo�#sN?�����0�[���h^��-D�}�x�Y'�L�'+����`5��.�Bn�u���;���2l٢(
��O��"���g��+#�!��<���ny�<�^S;VѴ�\e���z]*n\�Ӓ)���؝���;���s�}]M�I�Vrw�7��6t=c���JjE��Eed>�T�9�v%���q�SG���Q�!ؤ^ł�K��w{������6<�S�i����Z�,��=����f����q�y�����޵�4�@��[�&��t3���K��s�Nr/�n���v���yiJl̩�")2��S~#g�i`"�_��sX�;緗U)Ewf�f{��U��k���\PbӍ gsL��4��;&:�C�ʪ��ISM,�H��^>=ˢg�8���ۭ r�Ĺ��}y��wE��=ɌQ�@��(�ǌ�*�y�S��p�+�U�ݎݺnV!A�o5��z}Xdt���v�t)\s��J��Н&*3��u����(G9'm;�W	U�H�}qZ��FcϷ:2�;�ή�n]��k�a�B����pb���4��a0]87�`�k�^�n�R��N�O`>�2ȅ7
}�V��W1Ӽ�'�s��ָ�E���9�IS����{(�-t���=�s���g{��:YDz��Cت��%/6'��QW�&�t0���l��],nл�r�{�U����a�Ce���5�z����+&_������90rm#�4�yi��9�sƱ�}��J�����;+-����ս�GNj6�{["^��B�s�6L*.nPvǚ����*���:�s��x���mil^�.��T�s0�Ch����rֹ[qTժ\�$F|1lP+`���Bw�Ư�*d��E˚�.���s���� �>N�ל�<��A���4Ƒ��:|��<;K�����_71��}�f��*�N �v�l��4�UF�]h�r��9rH��gLf����V��J�����4yE~��1��^r�,qrU����Kb����MI����\��ٺ��1��Ĝ�\��з�ٜ�����zb�����,��<�1��Ȩ�R�4��{��j7FN>�7���!X؂���=���ɰ���� e�s�]�Y46��L۠�=(��V��Z��ŧ�n�r�[�u�{����Ña�$�F��oy��Pt9�#�0A�Oq�����Z�3�8 �x:���;,������8�k���KU��>�t/�m]��a�$x�"3�ZU���rA��*k�N���1��ڨՎ��T�����4U�ߺ��E�5��� ��� 	�=%wta��VR��z��Pzl����Y���L�If�[G�Y"C2���+u�e�;�n���]!0L�p`gT8�h��.#��J˚VE�|cfP�v,�1j�&p,m5d����Cm�*��y�cm��'��=�q�N��D��'m<Z�����X�����
Pv!�Q7|5����j�a�R������zh��de
f�R�]����ݱj�s6�It@k�p���0 ���4���Q�㸋�n!���ڋ���%�os��ܿ�2��k�G�^�Q����~[D�s8y>d��m�9�;;�w2|O��oH��a����.�M�.Q="/3��I&�^n�k�!ִ��a�^Q.$��&!��->K�cl�N0�ݽĵ9�������H�ޑɱ.�9���_5�ҽ	�ě�9�'�B�"�Z�U��5y�4mu��ZB�J$c㨭</y�Y�����n�𧺑�CԨ鿧�� �ٚ����'�����ݿo(���Nʫ=AHaN�*b�@"�d�*��`��"�t�gVzf�����,t�o�L:`�?Z���-����A�Ov��Y���z�}p�݌q�E�ƢIDa�!4'�>���쯂|D�K,pWZ�;��o{Ɲ3VŇ�u�:��� =�{�")ɍ���s���e�����y.C��ht�8��A��g_�Hv��iC��,�ٚ-ݪ������߳y�F�����%{p�t������5��.���	�8V� ��-��bXQ��8#�u%���-�U����ox9
� �D�|��m�k�{�M��۾��!Ӿ�q
'ʇ/��䈠tj����2�:xE��2��nguZT+�� 0���y��;�0{��:|e��U�����vw�kyb���9���/��U��9�Tk/@���k��}o_Y߽�`�CE=0%��	i����
��sS< �+��4Gm	WO�N^���U9Ix_d��(ѣ�T��,�$W����mD�Ʌ	ɰ�Vg-D�T�&)�c��b�;�ZY��B*>1c������<�k�h���^ٙ��y��Q[Ξ�r�·�z9<` if4F�b�y�}���Ojq�YؓH��6fٍQ��y�b��xE��.�Z�w^���9� O-%N�p@/b.^/���:��o:
�b!՟��3�}I�2wb�C|-����Q,�If����8�\U���.�Ĭ�'NG/6mK�Tn0lp�k.�����ѕ�%�k���j1S^��sU��X�ݨ%dԏ�db�wx]�4�)u�`B������z9��i�j��2���$��"zcھ�x�2dy��'Q��lN���a_f=�wg]�d2��؂���o �4�M���2�� 6k�H�"�R���0�$K�.�]�LbDݕ��v�0x.�rr��w�(�����z�ݹi�Qo*mֲND4ѰF�싆��]Y��_tS<��[
IwLW���!�9���m!|V�z�V�:j�[��e]%�e�*��B+�>B�B�zM��왏AVt͠�H�]E�dnj���
HnV}�_�guU����ؕ�@f�R볖�9�|�Y�56,�c�ݙA��|f�]�A��Vs���)�g4��vE�oW^�ȝ'�!R{�Ŕѵ�u��Wuj9�&MЧPtC��kj���Ž���u0�.�N��0�ե�2a�ZG�ogl2�4J�!B���ݴ�������J�휫����0��O9I�z�0VL]'^�T�6�u��K���i�Æ����-#҉L�6`5ح�K���Q���%��=�ڒo-��rkJn���7{(b�e(R�0=0�������}���ץW�zr�6�}��r�91F�,U͉�Vd�{:k�p��2�v�2,�7d��˖�f�].�4bwa��5�IC~��V�u�ʦ�f������F�(��LGx�����w����C�S����j�+#ʹ�K���X5��9�k ���b��g(�3s�����8l��7$����{}��oCgG�]�b���%2�i�3u�1<=�/���]As��cT*����ʰƅu��P�{ZS�5���^iv*��_v����Ԭ��u@�].�D�T��Lp-:v:}�m��t]���F`�˦I�� ����IѺU�j���Z�GlQ���Z95}�H)�ش�����8铭�X��Τ6��$],�T�'+сA�%��K�,+m�4CP��nP��EPPك�{-�6���f�"�.�6�_q�1u��d�\�����޿��+.���UP�B�X������U�FjQ&���)X(T��Q�J֥�F[b��5Q[hԣ�
ʕ�P��bUl�QQ+X"2�Uh���6�bmj*
�EѪĥTmY`�*�0��1h�U�Um�-X��,�b�PR�ҫ%��-�*V�Ym���mF���ش��T)h�«mmmP�T������ű-U��6����V�����QEKej��m)iX��j(V��!Y[j��+�+D[-�*V�ea[j��b���EQ��H�mQeZ��J�RT�����	���h�X�u:��).�����C�|՝ڏ	��)o�������u��%�2wf����ݮ��V$������/<5����<Cn�^e���n��l9��39'�Ra0��S����N�����<��U��s�q~�ݙ�G�}�2�h�;DD�=)`x���e�Y7�w�dP1��C�>ŧ�ϩ3�aѵ`n�X*��W�v,n�w:5y8��Ȃ���㚠hS����4��!6�/*�S��8�;�y�G@�e�*�N,R��9N�>a4͹�V�}����s�}�����Ƀ;S"��V���X����N$��H�Zm�_m��sٻ�F\��H�
"���YJ�������ƪ��0���N�ԭ�g�cB{���Zmxl��S��h3�}�a���=�\�K}W��GThR���[<�r�,>�f�?�eO���/���_3�7�  ��
�3X(W4)�V�X��9��h�W���D�ޥ�6 �H;�A��]�XA��T�Z�8�U��E�3Uv��<���	:�rU�ג�u�(����7��R�w%����e17��f+8�"3��E�X@9�2yU�Lџ9S4�A���{BahR�&s���.阙��̒�^��Ρg��"�� H�"�w�ƅ���C'�/�<��s��{g7U��]�����=�g�>��L}L���� |gO��<�-�������R�� ����Q���Pu��u+�uA8ō~D�����?F�>op�pG�͗�c���^<���,)1L�釣R��V6 ��=䎟!���|��u�y�l�$. yz+?~��ɥFv`$�L�:
G�V:�\��L�xz��`�$�Ii��׻�q2bLL%Ot+��svI�����ba�#8m�=*��׬d��am�gK<Gjt��k��[�%e���G<6�!�Y$!x��;5����m?���yx����`���~�^c�j�m�����x�Ǔ0�9�	�	����f�tVvv�/niГ�.�6Gr�Y >Y+����L���I�C�6D�UvH���Tm�Z�s�d��k�{,��YPuq�E���:|�b
:�+Ϗ!��:���+�P t�$OD�h��tK�X���H���[ì�d�6������I7G��X��OpA^�����U��e�+"þ1���Q%�����X(E߀NώRz�Z���Bv׉"���*�Yb��[�J���ވ����}`E]�;�%Su=�Оzc3iH�r4߅�Yӿs���߫=�p�=���<��o=�/\�ǄhŇ�9��T�
�N"�1��[��k���In�0�j�K_YOf2�V��F��<V}�ӭ_���7�z|����`OK�u3uU��ඃ����F�fL��G��=hl��kBK�Z
$aS�l��|�|���8aP� 1�C��?��0*>Ѕ�͟��aE�M��Nƿ����k�5�o�8]�"�Zj4�^iFpF�Ƃ�"(��7>��{m췬j�)ҽ��e	9*U	z�wa�AY�����ΝB� �-k8C-%s�54�һz��Wj��f�iS�
C
V2�.��4nvn��š�&��+E��/s�ei G��`����0�Õ��7�{iq�]'��3H�C�ʝ~�uJ�Z_��/�d�$�E����
iȎ��qZ3k�u�Iv���S1�P�w��c��u�ȇr`�B�����P3v^.�-�͛��|#w�=U
m�S�q�
򲦕�`J�����H��V�]��}n�8zc:��u=\]�w4E��:�����~y���#�4�� 4F�.jM�S��N,���]�仵T�X+�A��c	?ܱ��!��>'�:����H����"s��_q���m+f�qf�����e�t����rq��������]:�}��4}7'�����H�Fū��w�(�+��%D�^�6|��os��'���{}o��z���6+�� kR�u��^dW�:�����M@*C�i�-��8��2Vu��>�:m^Ԝ@�	�ٚy���$®Jsk�╍
�C
��Rb֒n���P�1��zAT��_Oŕ�2�u&a�ʷ���9W���o��t��1Ě8{51�f�{�8c�= uNj&#�z�����W��j�`l�{�D��Z���{*:���q�V����g{'N�wYפ*ψGLgT�97��h9n0�u�Ljó�.k8�c3�u��j�w/}�9��i�����đ�e�F�u����m9�&��Xq��sSuT}X�ʹi�9�e�a�y�#C�c�nM�åB��|����~C�v�/�����Z^F��Kȝ=��AO=��[�yӜ҇y��I4�3���4&X���h�.oٷ/j�����.<��7�Ҙ%�a�9���^a�c`b�fT��ט�r����L9VK���;N�/D8�"����7x��>~_�#xa�el�7	A���#�&�\��w`x��4'p����ͱ�%f��Xx֦[ݲy-���<��f��̬&d�Ѝ��U%�Yz���&Y���+-ڊJأ��R����Է�yC�K)@�j�����9���Q�1?y���ʤT��/�V�'(���6oAV*!����4G�Ӷ��o�k-�K�����qK��l��S��f�E^;��^C'�׭�NF�n��.&���j��C��=;5����L�=�2�@��V�������8\��>�uY��dH/gqB�=3�Fʂ�sݜ�}<���: �R�xD�Ń�6�Nv��ʖ�2���������
S���Q���3�⨏�$h"�w�Ư�*��ܼ|]#�hy�T��w-he��������Tj�c�L*e�E"���:|�9�^�2���c	�懷��|�M�bVW��J��9��Ka�a�f7�Ra��v�ܭn��T;ex�;JR��:G�gp`p"�$�
��P�?w㿄_��{�;Ƨ�[��
{�u�]�S��"��goA4D%Q�d(-�{6a75�׼ӆ����\����S�U��6n�7���J��Ǡ����%s�x���M(�)��\s�d��.��ʝ�s'a��
�M(ψְi X��r̙���\Jς�ô~=)��-"I�KM{���<�ȁ�_������#u���${V[z})�/)Yw�;(&,b���ظ<�v��%Gڴ��H��#1,)<�H4�^|x�W\�c�g���D�8ϋ�M�ʿwT���<�eA�/���X?dM�>j}�(�ö����$�K�� ���mS��H�6�s�P�O���鬑�� 7rq����f�a*b��%�{B�h=��$:.��ZG�����������u�������;��� �\�|��'1�y�h�������^ɳ�mX^;ZY�>�*v.0䪆�2{[�=Q��%u�s�*�v����s�X�r�>B�}sHq�$�+�������eiO����_W+W(v\�^Z9J�5����v_F�:�k�qɟ�{�?v���)�R�����-����q�MF��vBd'�Z�q
K �e��r�r�-�bjgŇ�֟���.�bv.;�W�IL�n�
&�-��Yط>�w74��}�?R��d����h����0����}}]��ގc'�a%���Vx����b~2�1֨!������AbI�eQ�d�u�
�e�&hm()i��,=�V�F�!s���$��~��-:|�4	;��������S�)��� ѹٸ��qS݂+]�cm������o����KO���Tæ}^`�:{�	��9bn�j���"����s�'1�̢x�Mg0�8��Ŏ�Yr̮kge��Ǖ�ȹ��9�ʱ~A�M+��\�>H� �=ӥVOg�����I���F����!�vN4٩Ⱦ0�*
qY 6��^{����ZQ���Al�H�x�y'_w4E���d�r�j^3��_��h#j�4��V�Cٹ$��O�=�hZ�he������a�˼3��-@78�o���Mu>�&���b��ah�����춮���%7/l�{rQQT���Z�������&Z��(�H�")H@a�sZ)�S��j�K��2�pp﫷7�j�ӃbQXǥ��J�O�CK�"�CִyS�gyL�s��L��b��Y����Z��>�r�Oyx��\�p��A��ͬTȶ���nsd\^�᣷�gݙ<t�4n�T����* �ceN��Wx�W�)���Q1\9�+s�:��J���TܹWv�et\�z�����v`u	�a�],=3\7�؇�:��߈�e8���o��Y:���26q����ű�`->��q��q�V��:ǃt�˗�����7dO�f�cU�)٫����[�c&h�39Y�bZ��{�L!�~>�k%қ�������#�$F���S������n%�v��y���\�x��{�j��M�d�cc�kȂ8�Yر���zT�'����VX�:C���Z����A3�+*�Iy��T���7�,�y��5[���M<��ˮQP�X�0��S�L;��]���ަ:L'��s��<���k%�⥧ |;?fw�mjq�4'?��.)�K�/+KOrwSos_9	�\��Ez�Dg��#�	ٿ`GO�]892����er�U.+ފ(�1���4I !s̞��� ��XNr�
�i��l���V/\L�ʿwa�c�H1�/L���BOJ���t��C�3n[4�s���Y컾ކ��#��-l��KB�(�鯈>��R���1 L�_F��U�j[𩉘�����ŧ��(Y�l��Q�)zݞ�/������������ :FK@�o�	��x�ǭx���f����ة���C��{�*5RM�+$Â���[>�#�ϲ�y*��<��՜W<vfU�z,����]�h �U�I�=|�ܙ`�Of]i{%�:�ܖb�IVu5��e߳޳���jC�JT	�S�/BaF�.����f菫���'����<l�����B�������lS�v54%j�W.��V�⬣�us0���ݽ����dJ](j����z:��"�{SEC؁!'��Ҕ�.�D���"�������+ڝ��3!�R���7.+|�%�1�[m�Mƥ��� ��ya�g�eg3˷z�8�m޽�#�z�õ��i�B����M1�i z��p*bo
�V��j�����z�NI>�z�[�
��}ܖ;&�+Pհ�k�x��yr�U�Z�,TD���w�DF�z�4�#V�'r��R.ty+�H�tz�4Ft'~t,,2uݮT�{A����j�{C���d�F����Fn�����y��f�4�NqоZ"�eP�p�R*�s �0�FՃHE;VS��̈�̭�{A`b�i'{��e>�l�ɱH3��u]�=�pm����ۦ���|"V��gU�$n�!\2���p#{"�뚡]�M�1�M2e�����*���g� 7.�g=�{[n��t�`�;1�����UK#��]V,\KwJ�lj�}$Z��ԯ��9��s��V�)nخ���:�՛*����8�ձJ$xeǘ�_)
�KDxu�j\�ߝ'CE�z��K��c�×�_��K�/k��V\�����87��N�ܬ��b6:�o�Z:N���U��U�$n�]I�ivr#Z�ܘ���N.�Q^����3�S�*��r=h��J-û�vfJ��^]�Xh�n��H�:�k���M6�t[��M�y��2I�0�����9-#�z�Rނ�V�ϗ!mZG���:�U���{�W���at�*��3��+��ir"`���r�ۇ��r�6S	�v�Ƕb�Q-nw��j�V�a�Ϟf�4Cθ[s���U��1��I��2L�%W�&�
�ݛ���MMӺ���n+�S}ۆ�W����U|@�Ñ�-��띹YڳVE�|��������s�Xϒ�*#y���7t��;&�J�a�t��CÙYsn��0�l����,"*kqZ��r��p�&�9�/�5=�1N��`�U�&�ͪ�Q�R;���ے�%sJ�(%ږ2v�B �/fܾ�)�V�4.e���S�\�2i�&��j`�ќ3u�3�� ����7��W��^]1E�eAAd*�����**֫Um�D�+
R��H�TkV(֊4���2���D*Q�-���D��h��jV("V[DJ4b���KjZ,Q[J	m
���Ԗ�X(���ŭ��Z��AbT�m�bԕA���kJ(�����ŵ,+KjVJ��K(��iB�+J�YR��ȖԩF-b�iPKIj4RVTQe[km-aR����*6"�h)Z�����P�U,Z�X��Q��)h[e�V�����jժ���D��-PXєR6�"2��(TY-QT�)XF��h°m�*�+e�J��Q��\��\��A[~w,��T$��N�,�+�W �>b+�:�0N�oL��O6q� 
)�g>�y`-�������Â�qTGP4����5�^�*8��̻ �귎��>C�ނ��j�=4Yޞ�O��,tl�i�">�>J�ś5��j,.Y���ٱo
���{NP3��b��L[E�.>��^-�V>'_o:5�b�ː�aK�V:i���;�U}�Ԏ��h�����^�=�t��č��l�$2 uz+����ɥ���D�D�Y=���=�[H<����Pa����AOH�f��.oƵ�+~d]�<y� ϼ���ױ0�����ƁҨ0�8�$�h�0ܪ��ϼ��nW�:����	�HY�aH��li�\t��Y�{n�hT�����E�:|zAi~6+_] �c��X?\L5��O�!8��xw:��7Ԫ��5�ͱ L��ڥi��.v]�X��fb����+�R���
Q�*_��zv���mev���r�A]h�D�FI�2�2� �M�e9VШK�3�z�6���X�d��%c���d�
�jQ&���%u����� ��"������]J��Yl̞P`gT(�h��:]�V\����wr�����u�э����\��&a�p{�,e�$���+��5�#���y<��¥Q��˗=� 3ヤ�Yb.ʝ���P�FM;�n�Wl_խp�u��!T���˟J���?�ũsHqD�MLZS�}uG;�Ntۋ;Cr��>���b1�����*�.$�x1W��d�g뻯k��5����/�y1�����ּt���O��ݴs��:u��{,���w�;��+!0�&�X}�P�Ń�Cf'����{yq$0����`��ə�8ZvU�\��P�?rFhm*:nz����B}Z�DO#u/ݾ�(_{��I�O#��Y��ό�>"��N:8h/��x.��wy�]��/Z�N��|G�X}c=L:k��g��c��uݟFM�ႍ�5V�� j�k֫d/�G�Km��y���;��Z3:.�t��8�g���6���i� T���u6v��:Ϋ��X�3n$KC��6u�78�s�������[SN˯w��C��^xg!�}%�$���Rqbx��ͳ;��b	,�RP�����5�ʱp���W�+�!PO�ۂ�#y�_v�F�%��Bj09SI�ڞ�r�3q��
�eMB� ��E�rz��<�6te�;0j �LԪ�(A�(9Sy�J% &.'x\�~v��4�N_	����z+�\��K�|^�U��6�˱��2u�<"~��ߞ���D71����T=<C�!��@D=ya���m��j�D��P��}b��C0���:{��l�8В��k��p����D������ɍΦ�nӞ�F�E���O�����Lk��OR���;}mt}�n��dxRw��R�.=���8�+ۗ��5?P��}���qS�Y��jycė�,=3\�/K�;5�<M�v�����l�pG���}O0�̽�w�b�������*| �:��wY����1|�m�6d�/M�U�D�jT(��^��o���)�C�I��
��.!��5��;��a��+�Q*=?5y�����ʎ��\o)q�jv��OU.��XZo4W���6�Ρ'�+[���w\�l����v<9�y���#�oO�kG!��b�iqDt��l��(�E�<���Ŗ�ͧ��9���~�\���M���y/#e$Ld�Q"G'=74M����9b�?|�o����/X��ŧ@�%亮�NE9}z�Uc6N�`x�S�x��-i�;�Rg�7�1��8�`���v�����ǋ�d��2&d��NrDU�6���'X���������Dy��I°�_F�n��0F��0��|!�8~���﷫1��n�L;�+��Ԇ6F�K��֟A��IS����;-UI���V���Zi^��W�C�b-��!ү���y'2�$3�Y�Ѝz�z� `�Bc�2�`�%����0�>�Y��o!��ք5;HGF
�I4�G���Wj��J�o�mjX��h��.����U��FgU�
�Z����|�f7����$��a�N@�v���x��^8�������>�Sw��23v��m���;�����խ�
TC�a�l�U���O�d�Yr���6j�[΅�ہ倁s�<]&o��.F���dI{;��=3���F��Z��Խ��r�S����1`�@6\�M�Ҙ�Х�'U 8�!�j�I�f/D?c��B&��;B�PZ�#A�}<o�&�0�f_���;9ŦE�ήb�xk����l��͞DGL_��
�L�ů�7G� 3�9������ޙ�pc�C���=0+h�R���fu��+/w�a�� Ls�/��G�R����C�O���B�UEg~lt5�W����!;$l�.V�+�0$2!��U���{t}2iF E����WY~�Y1$�bXbק�AO��="�I��7��{�����M�[-� ��<]�
�M��ю�9\TF�aq��&���WL��q�͗� �:�;��m�E�h�CY��Qqe�x���dC`.y�`�������\��j';�[��e�1�`����r���=)�/,d��an�#2�n�^�c6�zro�΍��P��d���Mi�li��G��ܺͽ���M�L������� ���65q�Pq�R4~țZ|�o��KP;<�i�4������ i�>ͪQ7�m��f��9V�M]��/���H����1�r+�/��`��s`lpx"�z;8Y���o'�>�j�bqy�T�T���A��Gg����=!�u}�i�N�����$�=CY>>;j�^Y�@�h?�����tC�5�<�XSn)��B��p����6\�
��ϼ�O��B��s�m�<Zoz�1�-���9�˚�{��3#��L�,C^W�\Is��U��t��֧D�\8�c"nzX�;x��e�s���ï�>�"uf�o���WJ��5&gR"�n�dK��� �!�ٚDV3f�n.�;կ�<uV��Q�qE.���Kk�Xף�̜����}I��+���3]���[7���)�O{�y>嶀�5��A|�I�g^���k&��%Ňt�������W�Ђ��6c��Vޥ�������=<��E�H�6��������n^��u|��pv_@��94�Đ5�pN�Xd)�,��eL}�c��-�Y�˗��Gl�y��m�ȝI��I�bkۭ��A�]�������bx�Ÿ���.�	'����a��3&�%g2���9��힓N��T�!n��7�)�ʰ��Ϋ��Ƀ�8�)u��4����R!�	�b�K��lq*Znq����;��,��o �&�PSL�ǦX��B�9���H����g�ל�I��Ls�.k����*O�U�s~�"simZ��\�ԋ��!�1�\2���&j�S��2��6�?��%y���ix�D�=/���[~�rl�,f(k�8���\�e.���w�}%e��t�"=��J\�>y�WZ� ��X�e�����Д�+�UB�ڌ2W݇���y��l���Z�6�f�
��۷���BR���bD�ݣ}��W����,_�d��Lq���~Yj �����j8����r�Vk���̗�TTY�b���ah��㶅�6h�9�~^F���u�`I�;*,�7ْ�}0�J9N�/wP����G8�}r�]���С-���^����S��G�x�������c�ʝ�|�P��f��J��\��3R�)��*>�����_?y*ؙ�}��<��M S����T�{��*/L��q���'�+_�������E��D���o�(�$4ߋ��*�3�i����$F�� �u��AC{ޜ�G��p�l�wZr�{i�X�l�Br<�(i���/�k}��Y��Pƽ�H�K�R\x��3{c9���z��1f�6�Z�f]��;��SMx%�z����4��z�#i#�Ů:gs�L�G�-����a��Ź�$���L֬ǾRc������~Z* ��Z}����2�Ge� ��͠�)φm��.��c33EҘ�5qLtᧃv{f�bn�D��&�2h[�u-����"\G2%PYr�s�f&G�����C�3������"���7�Tأ��j��!|�B������7�t�T���,L��8��g`�ui�B��08GiYH���"0��Kp]J������eLd��3��²�ww���t�O`$U��K�U��E!�1��hL
q݃�+jZ�7mjwEqZzk��k�Q��0�w��h�_�-~6s)��C$�I��̿o�'���5ʆ ���*&�,\�p"�o��~H�/O �B�7���|�OUܸ�3�{lLܫòj�3��r6�`�dI{;�弣;�z�X��M��]��Ӓ�5n}s�,���bv��ʖM��OP�w�����}Xǭ
��f+�y��x��x�DuiD E�紐����ٙ��z��e�^0����5�
>�^�&��e��͞��4�Qk]N�:��^���h��5�_����ðU��=�V�0�WN�~5�q8��J�W�H�ݲv�5��j�ӗ��Q�Q&"8�x�Ո͞�.�`�Q��M���\�5�!��S���;�j��zk֠�˅Q��t��%UՇ�rփ��clX]$��6��� #��AKK�N�س�0+}.����9��}٬��������}]!��@���|�^��:zD��y}��e�pjh$Ƅ���O���ҟO��bL�oJ��d9�������j��7`x��,�c�/$�Y���?%�)Y��*�׵����.��&5�u����P����d��B�aP5��H4���/y�h^�V��U\���:���T�TW�������0{�b0��qx�N�뤕����*`�>�
\[0 >l�i*'!"���C��3��ėf��y�D�D�|C1�x\��yW��D��a;�8KÁ�]�*�3du^�k'k�Vrj:ʥ��1*��S��C-�*;=О�>����+(�?��Y>�e�)�.n!��=ݼ[��0��g��3t_q@i|�)��*=����O!˳|u_%k	u)��<YgR������v� ڶ�e��0L���'��^�7I,��y�t���aИ��ګ���z�u��Û2����������`0m�x��2�I��bU�YB<U�OO؄�DwZ�ft̰�O>#j�֛r]I���cy�Wg�5mOjZܫ����(��K��\�7ʥJ&����;-����1su�RX@�a�*�2r95���I��֦5�φVZoUq �u���Y�Bz�eJ��b�����C�̘_v���� 4c�c��T"�a���l�r��H�W�I[�̮ќh����-}e~lg�u�9� �2�^ie��K۫Ν{W	�w��Q�7�����w9�]��;T�,��F�t�{6�6;��M#�0r�ďI*v�I�S;G�h:t$��n!�V;�v��\Gf�	�gx�w�8����@h�Ϻp����ǣV[#��W�m��oldv���AiɊ2����o�in>��]6�%�����]Yo�d���s��ڟ^G�]���HəX=�� a����S6b�Lߑ�G��(D���%�h�c���x*��u9�bQ�=�Ξq3����9W �۵ᵓ��F�(��1[���ԇ<\�sP�.��W��qk{aپ.�A��b��r�Y�N��P�g���9��vs$鐃y�@�q�9��Nu�

�2TB�f6�.lW�Z:��yCï�q�g.��.L�m������]��Y���r�$@l����'��z�gu�y�r�W&�-V3�;��bRܼ\��W��ǯ^�ZN=�H(������O7�>��ۗ���d�M�^��y���=�lKW�~d6�.7��$Q�0��B�d�\�Z���F��Jf�v������c�a4�l���ڽJ`'7+q09ݧC����9{-��l��0��cg�{R9{y�o���K\�hU�j�ٍ��3Ji�mUI�rC|��������0���zG��8p��Sx��k7�=L�*�t!��آ�M[�d�� j�Ca���d�yVtS�s��$��v���y�E"��P*UAE��XV+(�
X�Q��,��%J�@�V���5�bҵ���k]E�Q������*��#e�j1�$��V4j%`��+�l�R�A*4�Q�E--J�:�4[��Z��ղ��Z�1�j�#,TEV����J�Ym,�F���F(-j�V"���GYTjQ��T��Z�ؖU�����iU�բ�X(�XTJUX����
�5�m-���V
�*��4Qfb%Bչ5�:��-*U���.lE�#��)A�B�BH�H#�8N���h�c�����l�QJ�D �%�]$�،r��x]l�ø�0L�S`�w/���j�9Ij�UU	"e>��}�ͻc׬�/�mE��8��\�T����Y�1�k�Su�Q�^ZՉ�=1���VW�/d�0�1��+�q��S��y�R#����m���Z��^>>�~"�F!`l|f�a�yk򹯴�/�����|%��4><��X�9����3��F�5�)���ws=���O�z��%Ňt��Ó/v�s��� ��8�����=j������� ����z}Bz�����=9O*0*��uD[�f�{;aٚ����D�-,����;)�.5�eN0�*�&������>oQ���J�����mND�H�������S�.���sQ5��jY|��aTasy�
}���a|��}вX�%|E�Ż3�*����pX��~���;)>#5B��eX�?|6m���ɍ��+쮞Y=T��)�J~�n��ج;g�T�it3�5ec���v��W�՚p;�V�����\9c4t�d�:�ݗ�+��Pf��m��ǴfF��:��A��$�����"&e�0�e��t��6ܘ�M/�7�$�#
K�G�r�����p�b��v�9�Zu�5��e�i'�h�.zC��Q� �y
'�yqb�Nl92����?o�o�}H���T^��ˈ��J?1s_�!���"A�K��O�kbY1�L�4zfk��N��j���Z�%y���!�\f���ת���1S�H���p���Z��1��C���FVP�"�u{�m�#Ӥ�Z�����P�����vd���FNI�s���m��[Zs[n�!��򛯌��#�!�~�H*��.=s}h㠶��8.b����)<�f��RqQ��eMa<}���cėKO�\7�؋������v*6p�;cc�Ԋ%G�����U����`T�Dt�)tx�~|����z�o�P>�w����zA���NcLg�I�ᕯ�[o��%�ӥZ�k��t��r�f��s���f�׶�h��-W4��B*�L6����?`�@&��y��SN!�9wΤŻj����\���}eC
�RN���Zvq,IJ|�;���B�5�~=�,��vt^�بr�A��\G@�X[�ݙ<s2v^�s�&/Ϗ��v���~�\���M���0[!�w�vMU�M�X�;P0��\�H�>8������P���v�P�������.!24T�и���cg�z�!��k��L�>��m�vZ�iᾗPaҺc���(�@9ܦ	M ��S�F���
���������a�b���H{J��-|}û׿7.]�����d����/�!�Ó"}�_��X�r���5��_t��NI^�;}�y���&�?{��}(ז��}��q�,���6~�Xp_�).�g�z�1t�)iL~3�Uys�
���m.6���E�S�� �v�S��-
��SZ1�V�x0��1���w+��_yQ����,-;���4����v�r�p�{��r��[I�-����=띫7	���y����AŗIփo�6���'0a�<�]��J�JY}ʤ��rGo5���o�u�V[�#�z)��7��r�~�eܿ�ʻ��;��n<��#j�`�ȅ��w��V��pg��n���+$E�9���Ue9�@9��D���d�����0y��*���
Su�ͮ1�!�U�2(CDÛJK��W\�aP�w�Oe�{�oF�X>�zP�m)h9s�]E�|ns���O�$B��qu�����y��LЄ*x�ĜZ�=.Sҥ�zj-A�����=-h���7Rz��FU�|6w��UR�@�ZN�9�c��S���ñA�}�	�����MI��zȰ;��d�GE�W�֟Z&V�b%C!�{Pj�����g����L���3�I&#�D�=.��R�){zb�#S��$B绝Yxֳ��Ķςj���ba_���|�f�Ai輗���2��w�ɖ/�˒�.`�ډ���B�K��B��s$�Դ�k�?;�Zs���ڡ��퇀�ƴ�=�^� �u���x!�&��Ӽ�<��K{���-؏ ��S�]=!�ʎ[{D�Wt|^���Ó�����+���떌D�]*��@_^Af�z���ZQ�7���v��	�3�W��8��.��F8�)%<�mmunv�M#���uP�y:��ٵJ&�"�A�N�j�Z�r������=5�!g�5�M�%��y+�I������E*�]���m� ���T��:Z��b����M���r�`"fo��i��J�'M$���V�4��f�Ły�g�����Ol�ok�N�NCÓ��FMGkv%����>�^Ɏc��#�����Xjә��m�Ҁ�-p������Y��㾾�"�Gf����K�:�n���ŝ�&zp�q�V�G����&��=�Ǘ��#�&YÝ�|�N��ge�Ďz��`KN�&j�&�t�"�93�#�Ax"�޹�ݽkE��,���b^5���V���:��#��u���'��ݯ��c�D+X��%��jk�<�����t�6�kN&���O*���AQ���j-���,�I�NqRu(� ��tɴ�@�3�NL�k��aj�*��ү�܎2�5+��p��<t���V��T8!�3��XKyr+���q������(��q��������7,W?1R��2��l����������#���)�[Ԫ���;�X��*`�>�%"��=5HÒ�L�L���.��z��4�`���A������A�[`���
r*��\�Ҹ.{�c ��B�q����)�i�%�kVG<Xz�'KN��d;'���㪡%����璠pq
๥d$��G��Ӧd|Yf�A��R:�x���x]�bl����X�f�<ˡV���d�k.$��֠~b�/�."����|���2N	D��D�.��f�)ʅf��ȱ~��W�1y~t�9n���\�~��yz=��P��O�x
.�7/ ���eeC����p6�v�q��fwKYG3���I�Z��)���9z��]��,ٳG�n��;$w������R�G�ۢu�%]/�����(�v�Y���K-]h����ic	5�/@}�	>f�
R�V�r�n�Wm�b��V���t���j�9�ZRvS��I���I�(�x���ǖ����˓��������zAT��fuC;��;t��҂w�-$�?a�Υ����
�O����M�1U9�S���I3��~x�Y���G�X�ߏÍ�"�c����f��}�~� �����5�=0뺣��F �r}>riY|a�1��'��gC��.r޶^y�������s�hܷ�U��b�2���wf�U�˨W���RFbJ���H�c���"��1եO �r�ӕ�frOQ��o�{4��ZFj�	q��!�N�(/<�N�E�_0���f�>��2�˗�hūy<�J\*"'8x�.aqM,t�Ri�Zl�.2�qM��9F2��iѴpp��Pc�� ^�G��>~=A��	��2h����I�h��*o�s���m��Xظ��?���AG���I�F���P�mJ��&�.���m����R�HtY/� tA�;����ΟZU0�d�.2T¦��;�b����u�S��.$uX
���7]X�闖�8�'�vrU*Sɚ�&�.n���9Kb��z�+�y��!��"v֍!��"4�%�GO�X~�����޹)�ݽ>�W�Ma&6qD[Z��jㅕ*o�؄���9���;�kf�
��Z�U:r��ȶbd� �9ۉ�X�qk���.��nk��oou��|"��Z�s�]��ի#�VWFg����kJŃc q�vj6���"|��I��ϱiϦ8f+=�ڣ�箺Q�U�jZ�;1��T�p����ce���g�����O}-À�I�};1ź���v.ru�U9���窷A���x��_��q@��~�f�v׶�����x�,��˲q�����"�ᾬ�ȣ���x�I�g��!���T�5h��+x��LE��[���7�OMZ�.t����n�Gdo<mY��m#ዏrIq�F�ԻJ�<v���k�yا��]
�Y5��;�6� CDǓ^�}B���0��d5���U��K3/�w�fu_�Y�!U�Sa�8E1^�u�2�m3#���73��pc�Y�a�y���;*t�\�_Ce��I.�i�pR��β���0��=�Mi�sg���Ԩ���̳�,��߷����}�ւ ��/�.K���Pa����Ҟ�D��@���%E�G�,_���c^�هq�]s�!}�y&�X��ǧUV~��ٽ���g �ō���`.zR�}-
��n�O�0��ZR���Ϸ��D��ޖ�~�x�V^#i�?��������f�=���:��s�w�?4�o<
xK�1�*s�T1��w	c}i�����8�k�㱚^l^2�j9�z��d���mIƶ�>�Y"|a��K���U�+�J��
�
;��{�w=^U �f.4��u��'���z��<������OX3~��Tv5�����D�3�d%=�ݩ�U�VX�pmk4��({bz^d�FGH�=z����Ȍ�r�٩Q~Ò麌���OCݨ�
rl��d��y���GY������̊c� �����A,g�v,�f�o"i�u�u�V�5�ڶ�t�ghu�R�{3V'+�l�T�Yc�Ү32�.e��vQ�b��V.�+�a%���81��؉���j.N��'�xq�ڮ��a����~��^>3���[Ta���d]b���O[�eG�y��*9�xK�����ɦ����V<���;V��m4B�p[WC7E��ܷ�M���M�ɮ.fnzR�сɞ�����d̾y����V*��Z��	ZQ,0{]O_�=*��+;���A�Kx�{��u��n�Ӹ���x���gKH���L< ���ANk�A}�OA۫�Ԫ�,�XD��,Jvt��������m!�8t�y��la~�W���4u��P�<^����E���B#��#�G=���<_e-W�]FN<���6�&+x~yq�1gjY;�H�=$/v��'�����1h9p��c����CU��z��W�	]�Gg��ୃ��vN���կ���1�(��0��/0�x�[�CN�}�݂+5b��7ω��5�靲���5�k�d$v$�Z���Z:o�;7�s�[ѢI�+�3kp��!���v�\�6���Wλ���Q������h+�V�CF��X�,K.��d`b��Ob���3-�A���7�ܬ\8?���Fl3y��Ӳt�	��|�`��c*�a�J�3��0Z��fb����&�S������ �Re讏�#x�w#	.���$F,��-���C;A۬��Λ�0,��*�N��k��m�0�c:��1g+���H؃�Ky���4ӌC|S*_Z���Sz#��Kf��IDf��@�/M�P�g��������y��q&����(t��8�uܞ��<{�ڻ[V:�u�-���ݪ��ԋ������Qni�9�����B֮�jnL+P朙.F��d&���ȆU���{yoٓP<	Ӝ��&`���L>VB��d�ot��ǆ�����23�K�L���a�XqU\+U+e=)3�(3��c�^3���7v��*=�pf,��ݟ4��tv
��5����c�9u%�߈�dod�S��j��$�{�խ��`%���/`���=&قQz;@����W�~�:��@�h���Z��gP�B��68bm�*r����ئ���}%n��5ƓJ��v�WA�6-�h��Һ�-��z�si�;�)�v�u��a��/�%qcua�K���:��D\��h�"����y��;�A�d9���p#)*gq�fܸ���N�5��Y8��bO9n�'5qbd�j��Fn�93S`����"�sÓ�H4&�Y7J۪�ʋ��&���Cs�f:vf�]O(�֩sP3�ͫ���м���%cy�^�U����o,}�F�Xo�v�Qi�y���j�Dc�2�o�Ӕ0�:C{��\gܨ=�Z�N�3��3�(P�r�z�C��A�� f�mS=ղ�X��(ɼ���+(�J�ZnTz*z���<��\3cFr�R�7�j�ed[*9@�Ғ�xjS2��e���Iw,*�1j���x���NֻȝF�(�M��'�7z�SF�-��O�!{5�i��:6��t9��Ǟ'�m����[V/�ZT\��4��l�Lɒ�mF�ɓZ[���Ն�)�C0m
\�U�	��c9�
2�5����e�����[R�YR�TR�ڪ����UD���V+S3%61�Yvì��Z��5�֓"�YP��m�lR���ȴb6-l\��"�m��E�[j!R�]h�!m�h�4j�me�Q�K-*("8�s��mmDZ�l,�J�����X�Uv�։Pڢ(�cZ�T��.L�ie��J �0cZ��*Q����iD��f��V��"d��Z�L�]iY_���NS���㑗��c���׸t[-��r˙Zgi��?s�P���%�J|�LCxD��������ٮt���e����]O574!�b����xo�2�2�L���Qq�d�r¨����w<lJ��YCS[�]/�5�&2U�'W���v�s��0���.&�xҫ ��9��5I����sP��T$�յ��8U�=;ޞ��rVR�4�l�SƢ��k9)O�7+xLewS]<�"��S׼�om[6z��]^3�\ԙ��	�"�/��h��V�e���z4crm�O����V�x���u.�g���U��w"���=`k�Z�;�~�o:�J��~'�9�\C	��jź
���p15���D�vLoՇ_g����TfV�����tt��e��U��p"�d-��Z�0q���e�|p�})j�,ˣJ�TWs�[ �b��gq:�O��q>������vsyΖ�LxiV��j��t^Xt��i�8�ݩ.	&�$��brn]�{f1^�s9hAնO)�yl8"����m��=�~�I�����{�[�=�ւ��� �U5�l��R�\8B�t�^��=�B�}��)숨K�/*�?��]Y�
��3�;3ɑ�73�	/�gIU�]:��Q�+%��:Ol�JO��r����p6sk9=̓�x��upg��;�U���z���%a>���ӢnvwЉ��jL�wӘݥz&�(j��5��ϵ$�O>�?d3�*��S�^ٔ�T����u2W6̺Kc�?,E�C�a�����O���7������p]ɮX��NS�7��A��n��m�����W&/v2xԫ�f�l��!<b�X���ͪ��xHQ`!�W^D�!Y�ա9W�f����cuI%���nP(K&M¥t��:��&���>X, KU���^ާAjq��^1隐��/��|cER��v��@�}���܍�o9�ܲ�,�t���^�U�ҫ7ᕝ�Og3�	��}�g��WF�.�ZLʒ��3�s��)ɭ���;gWB�]\�-p��*��u8�@6bzF�s<�Ş����y��o��5�D_��߸BW����;g��wދ9�{���1���R��6�7�j6�HT���N����o�W���8��b�H�s���j����w�m���F�nZ��˱��X�u�mQ��q[:j�v`�I�P�S��yL���wk=�۾��G�LK$��EV�z�.��]H-U3mV;Y�����L㝫��u]]Et˝@�8v����ur�����\W�;��mf]^e��n����KIέ�`��`��Ĥ��%K��hm�F\�!��<�9J��!kV9[�9!Ǜ�}�ө5q8ajU�S�ŉ^d�폮*����3���w��S+6{z��䖠LK=�+�,��vUQ�6�7�hD}S����ݹ.�����u�3�~ò�:�0M{-���7[K�OXG����wF<^���\>N��R��f���V�N���9��	�RՔͧ�+��qOi�B���O��&�٧�/8m�7y[�j�~���EE�7�xo{Cxr�*��j����Z^�.�u#~�g�J�S���cՠ������6�w��p��{��g=�5';|�;�ͽ���O�x��A��Q~]�u}R�S���ȳ~sC0
Ex������瀣3��45�Yu�\��9�ޒ��� �^�v��# Ħ�@�j�����H�c��w�W��������?n�c���j�=j�mԧ�V�jv�^�oj�]�Y�a��xsz3��F3Zh��(��@t��$!'4e�e���	
�;�ngDLu��
�6�w<
c�ܿ]0��g�����VF�|�Y����nn1�w��I����i��>Bx�	���֫�����r^�4>y��ᯩ�>����Y�*����"���W��^<��騘�;�Ξ�{+�k ��r9����Ĵ�=T꫶����Qz�+˥d�r¨�����|:�� Xڒ�y7x/2��ghө�蜴�ǳq�0��:��F'�5=;(&=s�T��j�*�^�_��s��3y�)��/��<M���vTM�|���GF-`�S�pC�ٽ��֋�r�-k�����Q��g�N]�[����<����������t;�K����	�w(�	������ݳ|^e������:hp�|O8�(+��9�����X��`�mt�X�A����ɪ�w�b�l�+X�)-��[ڍu˚��_r{�D�侉��R̸�*��TGar��s1�WS��\��X(�Ȫ!�S���3�ҙsզ��\��脛O�w�
Π�w}=A����~^�v�]�c����~�ia8�.�r_J��$+��C��+U��j5���iXų:u��6��7vsU`�D{���sv!�bi�'���|�;Lf:o��q�N���q�b6�7e���Ҵ�W�Z�_-1��2u�ȧ�P,NoR]Y�
��3�;9�ɚz�F�+�?���5���͞;V���F5a�=^����Ce'��6pD�;��v�t�K�,�κ��\��� íoU�7��1�#rS�6����Գ�c�(3Rh�K��N�׻��6j���U��,5����7{@�%�+o	��8�3g$�S�X/U<����#rPj�;e+�����ӦH�[p�Z���ެ�1�	\�](�#שC��������x_hV��Ǽ��.���y��k�r;�\�	�/f�{Z��W���Bt�i�߮ry�p���s������[�b��ޖ��%5e����l�lJ�k��;�����w��Ԃ�-�9����b�b8������V�Q�}ټŒ#�.�8�U��{�Cv�d���4��_^s��y��1�v���`�'{��������TN�ĵ��\.kDH�5#u�ʽ��w��pdG�����ɍoް�<4S+ψ��o�
���/m+q3�^C�a��]V6s��=�\��q�@����]*�벲�=~������L�}�	�6��yrp�C�������N���V�s'=�h��H�U�v�=Eַ*�'�9�5�Ũ�jD�V<�WW�xݺحT�cyo�Q��s����2���ngL&#���Rע�K2�5����p9(�o��vjY�N���*9���U�r���93E�"��ت޶�ΪW�����q��5&�g����T�ޞ>���"�adEB\�٣k;�.����6�-�G_C�C57<�n�*.VxoV�L˃s��w:�{S]X��j���޷J��£�ꉪg�$`��6�``��à��{��-N�Ԝ3���D/'c*�n�9���{k,T�=J/bq��T�^6���Lޜc�tmEgf�9����9�UW��j柴�Rk.]Ɇ�A֢�9�YƢu�8�����l��������J�C3��d�)�N�zU������>�.0�i�7�+�w{�d�ã��"'v�H�f���t�Gxs����5(5���0��ͻS��&$�N͝sЄG���3[�B:Ͻ����e�m�ue���m�f����î��wD�D��v��"��6�Y��~��	��/˝A*���]nC��	�z2�O�:��vY�=�ei{I�|��G)m�^4���'"���Y�XWQj���o�T!Qa�/Yٴ�g��؞�$�꧷XU���}��W��01�'�s��aON��/Kǐ��������s�c==ޘ����9��7�uG��1������N?���|��N���Vs�V�<�����6�-�e�z󕗃�s����ȼ�t�Bi:��D��oYTt��ƬG\怉�\�
[}�}���kU�V�Gx=y��A��a�M�3��|�Z��1EŢ�+:��H��Z�k��*l����{"+b��	�<��5sv�^�·�	�>��Aٷ1n`�e��A`B�s�^���G��nut�.�)����ޤ����t�4������1.�t�Zꍣ�Wi���r�>�;Q�
y�سx�0���am�M�� �O��Ĉ�踡u<�r浊;����Ǚp�qF�Q�q�7b��yD*��k��ݝ�w�b:��mn_�C���9 �`�}O_h��[6���(<��9�cW��ڧ�̂6�7�����\�f�� ';Z����ñӶ���^j�6_w���6m���%�3�;d�wQ|<_�Z�g��;7����N�j�<>��*�����;�9���ڛ������K�o�Z!`��Y%�X&��m�;�`P���y�����M,�HHHd���O/H�:�MAu'ى��h�,ر�d���"\L+�K��֤磞/�=��iB KJ@��
��k *U
�@-)@�$![���Dw\�p�ڕ�TQb���Q"��mEE�,{�EY;��%�'��(��c(}qԤ����UC�Rդ���G�]�H�(����R	!��@f��M�_��a�3-����pR��}��-������(3.샤�Uɕ3�W�2ik���K����D)�a�uͰŠ��QO�M^ӯG��c�	�O`-�J��)���p��(�>HE	�l=@q?9w`:����o}�].O���3?����t��C�9��VQ�⊢�d���봟���yȐ�B���<�)�ʦ'Q�K�&M��vS�T�|X�D����~UE�3.�4^^\�X1@�1���B$�5�Ƕ�قC���X,
TTE!���q�>���R��8�N(0$		 ������9�d�H�ňB�4ؠ�4(�)V
�^vl�#p�ǆ m�~�����EDSh�B!��"��UH�F2F��v���=:��sxc��I�^�Z�{��s��&��/ֆ�?P�]�=R�����>�
}IV�N���F�H�� TR�h�Y^�v"}��i���pQ�Ch��E�Ԇ�)`��S�t�v�;^A�ɯ�8��A��X�!�,n@�q=!��=��G�E���S� �,k9�9�7^faxd!x4�~��	A�$� 
��!`䊢�|C�~�H�����8(M倸3<�����\�(٘b�,`��&����n-$H���V
7,��h�
����,F������q���u�k&�!UC����n�H��ni�-�(О��9��q�;����B"�(���죨�<�q�p�EQE*�GP�� �{��4N�Mq�t~���}��m���/!�WB|x��K�O1��iu?�,N������5�Q;����,��?l�ϴIq���TQNG{���	��I�SBo��L�>�UR��8C&��`>�f�v���V�7	��ch���Bc�FD#d���\�e��:��������ݘi�1��3ͼ�w�ӌ�z=�-z��1���{$�pt��TQK�� �]P�,p8H�\i�b�C2n!D'�0k���BAӞ���r0(�f^%�X��TI��:�jo��UDS� z�>�,����P)�!�{�GQ�kսUQ�ǘ:���q�hb�=48�� ��m!�Vﰝ�y���#*
D�'�Ѱ�+�9P���H�
��	�