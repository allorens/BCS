BZh91AY&SY��K�b߀`q����� ����b,           �                                   4  #>�}
�!��o�x   �@       �(` h
 P                 3�t�U)�R�E	��Q@*��
���T*�%*�)UJ�R*�(��T����*J�
�|zR�h  t���*R�BP�(|��oaʅwgH��w�:A1
Щ�P��J�ݝR�ݝ�ꄍ� q�Q*� Z�H�����    ��$� %*��^�5���y�
{5Rx�}'���W-6 n�ǰ� =}@ ;�/Q<�d3�w@���@�{��` | � NǏ�J@��B�	I	%RE2d��\�K�`:y����`;���X �w��8 6c��0��K����ǌ{� ;�}Ԡ� �|�� ���   m>��J *������� q��J�� Hy����|�����b� n�!+�@�9� �s��c��@   �})T ��R�)H�@�d�T� c����yz{ <�@ �T)8 l� )�1� v;�� /y�*� a� ݁�   *�� X@<v>@������ 4-
�{��ܤ����2��n��     kϥ)@ �TP�T�(T	U�Vc @��: d c+��r �����4���`H���0 �� �΄( �|)IH ,���!wp��(� � ���M(��`��R��wc��;�@�����   �/�JR� `��I(� �R�:b)_ n� ��`�`��{�GuJQp���2 n��o{�Ж!0lt �8   *��QJ �� ���n�RG -c�`��Y�42 ��*W �݇=�{�7XCs < |Q$P   U  �A0�J@      O�4��J   d� ��U$2R�      4�*I�USj@4    �JAԨh 20#M  �&�5$�Ҟ)��ȍC4�#a4O����?���~O� 
p<��78�e+�����[~�EV!�K��*
��AO�D�_�����"�Q_��N���h�����G���a���w�����?EV�ԒI>�����,�G�'�E|������U�0@��U�@��F� �1E�(�@-�L� �WLm���U�*6�Fث�[[b+lm�-�E� ��F�(� #[`�lEm���Q�
��Fؠ�Rؤb�[`�[b+lUm��l�b�S [b�[[`[[b�[)��A-���(�T��m�c ��m�lb[��Ŧ�-�lb��h`��4�-�lm�m��lKb[���%�����L`S�Ķ%�-�l
m��&��[b[�Ķ�-�lb[2ؔ��6Ķ�-�lKb[`F�K`[���%���-�lM0�%0m�lK`[���%���l`[���l�ؔĶ�m�l`�)�l`i�lb[�6����6���Ķ�-�lb[m`��Ķ%�m�lKe����-�lcLm��[�:b�ضŶ%�#`�ؖ��%�m�l-��Ŷ�-�lK`�m%�t���-�lKb[�lb�lKb[ؖĶSؖ������m�lbi��)�l`�ؖĶ%�m��0-�lK`[؅�-�l�$b[�6���m�lt�`�ض��F-�-�lKa�%�i�l`�ض��m�lK`��l��lZb�ؖ��%�-�2ؖ������-�lKc�Ħ%�-�lKb[�Ķ�0m�lK`[�Ķ%�-�clKb[�6��%�-�lKe1��4���-�lKb[�i��)�lKb[�Ķ%��`S���%2ؖ��ؖ�A6��%�-�l[`�Lm�Lb��6Ķ�m�l�$b[ؖ��%�m�l0�1m�l`[ؖ��i�l
b[ؖĶ%�-�l1�-1-�lb[���i��i�l[b[ؖ��%�-���`�ؖĶ%�-��[�6Ķ-�-�lb[�[��%�-�lKb[�ı�l`�ض��%�-����ؖĶ6��%�-�la[���%��%�-�lKcl`XĶ%���-�l`[ؖ���`i�lb[ؖĶ�m���b[�6���-�lm��Ķ6Ķ�-�lm�l#-�lK`[��ؖ���-�la[����-��-�lb[���4��*�S `�l t���K`l@m����!� ����� � ���"�Kb�L�
�0� 6��*[b#lDm����*��-�A�6�� �[`lm�[H�R؀�`#lE-���A�"��� �� ��ب`lm���6�F�!LQ� 6�Lm��T-���T� 6��"��؊i���T�(6�� � `�1B؈�1�
6�Fت[[b�lE)�lTm����� b�lm���A� 6�F؈[�m���Q�
��Rؠ�b�l@m��B��lm�����[b�lm��@-�0F��]0A�*6�F�
�B� F 6�Rت�[`+lQm�-��"[�@� ��F؀�آ�[`����Q������w?|���o '_��kٳ�^Ԭ�ov�^�+L-�a��4@�"����7����엃bŅ��s޼��D�7J� ���>�Bwq(-��ޖi���8m(�=�QEۧnn�w�~�N�5�&tvn�g�+�k�Ѹ��8�rݛ>.����F���Xy7ƧJ��4fߎ�i����a���-x�!���R��H;^��'Sˮ�ҡ��-=.��:wN< |�mX�
��U�\�;��@�yx䊣����K�D�`�FM(s�C%���%��X�hvv���Lɼ�.���/3tB��6foN��-� 
Xg3��ٜ���V��9!wrjYN��u�-����$�8�#H�uD8��w9�g����h����Ł�&LО�V�NtK�0t6���/w�vl�s��}���)v+�bd���c���9�!�0�usN�F�A��r:Xm�#�$4�q�����v*ɏw��p�h�j9~�̮��z�ۘ'-�%�!��9���;��#��j����;/q|��]��z��X���\s;�@܃������Q�<4�9��ٓNʎ�f�46�Z�<��'f��:Dx�%.uT<�5�Q�Ⱦ ���k���{w|�*3p�[�)�ad�7oG;4ʒ��ؔ*�E*&3�����;`q�j4�-�<���:��ʩb�8'����X&�Z[FI_`s!E�P�M']/�q����4�]G�v�q��`�g���87;Q���#nEX�]����w^�p2�G�f�ŵ�ٜD���j�;��N��AX��;Fw"��7�
O��]��M^����;�=���]���8��'n>ZޙW���Ŗ�`��=�w��:+L�r%�5��;GL�f.7VΆ�ɼ����$.�K�7zۈ��ו�ïoqc:\k/[!�]�|�=�<+N�M�:Mf���Flܧ��q�t�w#9�CIN޼�G�K�����F��_rz;����\qN{G��m[���N��w����2}�lB�J^S��2�����я����nnL|t:�>	O|UQE;k^-�@��3ET0y�Jc��۶���ڻy��R�&��X;����;^�ƶ3��L�T�7!�9�-ˠnW�'�j�G�wx9D/䜜҇͹;nh�U������w�ځ��4|�\��BW�<�E*�Xnѷ�1i͢k"D��A3�L;�#�(����Wt��/|
��:�MD��&2��DH� ���;Ho@����&���0޹;��7t`�ЇG�'�ு �.�w;u��}�/����;��r�� 3㗳[��^��I�_�Lߺ���	��Zl=q�Zׇ���Q}���ܣnH2�߫`rkZ����;<z4F]7�٭�f��=̐!nq�����3N9.L��wu{2�;��\�Kn@GT�v'���]S��zq��q�9�wf�F+��ˇ��u&ć�.�wX��>r��/ ��;�e�0k�Ů��ǖ{�7��q����8�;��X�y�-ԃ��fŻ�Y=�˝xoB�0j�A���6�S����&�7k|��xg'M͓��/{h�������FI͛���z>{�Bi�>���O''�v�qMjc's����W�84,�]�lޱv��/wVX�0�۳�ʞn�H�e{��ᡍ��¸�rnvH΍t'%��6j��nJ67��[yo\WnE�,�WH�H}���ϐЙǅ�M��ս���$�®*��ِ�ό��Q&�[w[a���lԾ@�����|��á&��o`�0p�ǃ��ϱw8������Q�X�x�����r������Ϟ�ٿH��+�	&��wT<G,8�60ϦGf��Y���5�wn��o�V�\GL�n�8�qcQs�8�y�gM���pb����
T�e3��h3��Th���w^��^<K��7���]ܙ�l�(m"��1��:U{4F	��Gt��3�P\��V��KU&lК/��M�l�9�K#�n�� �n���5vv��v�G�t�P`�Áٹn���p�zA6]s�:��9F2;��8N���8f���滝�:�%��jvn�g=ǌ,�p�;�=�0r[sc��,6s7
iA�u�����0Hd۸�*_�0Kv��2F����mʄAv�u�nd��u^�g�h�t^��@+.��<����'T�˻w2N �`�ii`��΀^�;Mb�0�p5;+�-��,,�-k4B�m��="M߮n,�-Ѧ�}�<�o��3����]ӛvܺ�y�Lg2?��Ca����\=�"&�eqa_Y�r��[Nh�x�L=WyN]8(
���.M�{���4M� ֠��5E��OUgpgh�(���@]����7�os}vԌ��:l�AQ��Z�]�鹣���Hm/{�Wc����^4uu�u�]�.��q1x=���XŧJ�v�Q<�Uڰv�L��ku���	�a���{*ے���׵c+Z5��T�m���(�rr�CsI�)�ݝ�Cy�է���p��7��M�b�mO)�թE�Hځ�Ժ�K��Zz7;��֛������V���.��	�ӈ�/c�Hy8X�<��0��ZY�v-Z�@`j�m@�G��u���vZY9�V�76q�Az����-�p�!p����ݹ�+}��-hL�YMi�@�͈�ހl��D.�5��wsT����n$qô=8��Qq,�{UlS��e��M�,<9�Q����M�'T����b�q��h�l����-�`�`U	��勤��y�=�2���a�XB2�Tn�|�4���ގ�L��T���ju�8���f=ff��rת�:�3�y�3D��q�c�;�+�WnI��:���fD@ɱ��,9s�f�*�#� *����^.ݝ��v�׫D�)�ss@�:�f�
�3l�ʞ##�Ks��X��ۧ5�H.��W�����ٝ���}{��$�)�`��ڹ�5���;{G���`;ז�l��ǋ7%5�#p��Z�Ihp�;~��UT�k�Tuu��ڷx�s����)i�b:�J�c�h��.����^��s�a1�wWϬ�(Q��?_��{�`ɝ8��ِj2=�Q!��yýp���D��;�Jn؏!.��p�͌c�#:M��.wm_�m��7��b�Պ�d��/k.��g:����r����{��f�3�X�s��_]���7��:��'����4:G#�r��vU�v������n��Z��2����uv�|��9W�4I����̠�@������<�%���� �7׷�8sf]�/l��w6�������SpM݋J{�`S)���2�N�]���&�qK+I��x H��Z�NI���GH㳌{s���K�s�H��]�GY�M�`��;j|�Z�=�&�F��2hS���5Ւ�W��-��7E�t����4��6���x+z�6@w��n;��r#A�C,�s����vJ+���u�nn+h���i��`Deye{����eQ�嗊�^nIg�=�Q
i�;"��@�������ڳu>�`�ш(#��oC���u�wi�5��oe��@;&��-��N�lc�E�iL��q;ǥZ�`�����N�s�U���|��0����"�Z8�E����h�+4��{8�w%��Ɖ*U���S�LN�=qc�{��y����dvrU]�#n�)�㏹sC�:u�_[�&�ۻ�P[\p�( ��[f�VIӮ]pam;kҴvF(S%��(:�%vW�q�� ��UhQu��{���u�*�^�x��#���`��3A�C&>�� ��p�ޞ���}�5����}g�$�E����0�� N�l�̍�{8��s[i���g^*�q�+`�X#:��̈́ �U��8��:��V����N�Y�!ثJ=��M�W5���3��32s� ��3s�-4"��2�l�01�Ώ�@Jd¶�DB�����;����Ϲz����/.\&u���x����/{����$��e�,�_|���v2�T�LrUL.��̣uDtMq�G���kmKA	�h��3�]�bP������f>�<WK��7����kR-�T���N�5gh�8Pd�a�㭺iWϮ����G����,�[��pѬu�i�.i��d1/�=ڻ;���<�wJ"��'x
E_k:��3�)���ٓ5%�ZK����l7xF�k'e�dc6��N{O�}���>���!���H
�Z���t�B�+��5o	�x�u>:����V�.hrrP���3��,|V�ܤ�0B.٢���GIݷ&�qU��ĺ���i��t��=í�725�֓�5�9��f�,��p��� �rn9ڂxh˷����{tq��7r��<�mɜIl��e[�#�����IWpT�9�MTj���0�
}62~q=���s{��8 :栌Z�����D�ƈ��|���gN�Y�pk�-���s�]���xM����r�ɼ������.xNJW������È�Z6n/s�1�K~6�1/V�Ii)v���1��>il�tu���o{����Ah��8��f<8\�&���;Ǡ���_�7���.��Nh�M(�� �>=�(cN�m�����x^�W�d����u1#��{��RY�P���a8�����M3t�7Iǽ_-a��!�d��A�C&����� --�8l�6	���{r��3�n�ķ��6m���o�[ƚش���V���
Ķ���{���TZū;�7��0�*ӗ�y�%9U]��+�N�SrnDێ�t�e1��يYA�*�V��q%�3�I��M��.�������3f�X��h9�4-�;�&�ܩ�e�Y坿q��Ғ��Z����c��������C�we�{������8����5 :���M��� �`���Gjob"��B6p�[S��9vd&���ݠ����}ƼZ�.�[]��so��+�l8���;��	��@@f�ʙݫ_Ǯvw8�����pn��uwڮ;-�0Do�&B9�1�lS{,���gvE��ޢ�5ۡ�b�[\���1���F(k��a޸�b&����WM]X�`Z��[�m�f+���� ωY���.{������e�j�u���(]�7u��k�P�fږh�!�	-<;Foc��J4����3h�fǃ�;ظ����en�c)t�����d��ׁ�y:q�}�NsIm`�o �=�u�^T������69�̗�T�MÜ���:%��ݶb�#Q�Dג�JƗ|�lf���W>ky��8����!���4ign��v>&>@�͜�d���=���V1��F�����[��&e�3�	P�	�,F5עtεܕV�os�-���hQ�;��n�+f�ra�g��ͺ���kt����B�D��������t�r��mٿm�c:�P]Q�p��^G���-7(�U�;t�$���*m��gOP��p�Gn��v���ոRZ���Ų��욐[�[�2�d˔���bɋs�Xs���:@���J�rZ�M4F�$���˸���V��
�&&�=�rӢ���r�ӎ��q�� +/.����Ek��a���5�ֶ`/gN$M�n�:�G�amѶg@V���!�M��ҋ��c*�z#���=�\����T�kI��2����y����4�<������a�!��<nF$�X�YF�m�FXN����I~/.�(�zeEo�	s��{���jˤ��w��|z������,e9DD�[w�v����G�m�t�\�{GDG�vط����;�}�퓻|�ʹ�7�^��<>�����f^/����+��E��V�?O]:���$��ŗC���-�c���;��:V��vǎb�9NG��[x���ޝ}��=���d�o��{w��f���<b6��\1o��3i�0�NZ7E�;�a:M����i`U�B��k���_����4�Ӭ���>#F%�Ke�� NQ�r9?CN3��0?S<k�Y�����#��@��Q�YyӉݾ빣R!�I'Ɠ�˽���W�G�oe{��]�l�q�*(����jy=|�%�%ޞͤ]���{�E�,�F\���7Nx�������Q>P���?��LR.���u�\���3�Bo�n]i�ޓ߫^,�w���7��m7ܴ�q�����+eO�o�x�c/���k�w�A�s۞<�O�y�r�@�����L}��@�D3"���W�����o���i͵��,�G��]��}4GO~��f�{�����q�G;F汐�L�ZY�X|)O�M
]=K��������6�����A�Y�K3����ùw�yA��/'�0�� 图D/; �^�>\�!ͷY~�m�x��x�V�՞���=amiF����2���Ms}�l���iм��I�r1M[�^��ҋ��p/U��"c��w��獫=<wak1"tb��$�j@Uhp=�}�L4�����l0�\�^��)i���̚Oqd"_O�盉螰0����q�W�����Eo�2#��͘�])Nퟏ��H=��V`���x�	�2�}��R��LLoxw�2-�le��Y����A��;�NE㛾�Lӎ��կ��O��jkq�bN��x{��G�����9���"h��儖x�e�-d饃ӌ�~�3��S��Qor���Y0�.ꊩ"�k<�)uSt.�ز1w	��O�x�:�Kk¬�Tǡ��='��?�~O�"���[ߔ�}��S	�`}��H	"���"��!��#QQEj"�QFET'bM���	0@��E	FDdAV@I�Av��l80 ;`EE$DI P���TY $�$`P��S �`ˀ0�6�$6�@0N�&� ����SL
`'�lS aM��0
�* H���+ ��m�� l���i1�b ���(�* � �"� "� ��* �� �2�$�)"�(�TQd����@YV��H"�����UJ�_]֊�'>׹��z�G>#qaI�j�u1�x�kh1�I3#v��u�n��ߌ�צ�d
d���F
��!
S���	nl�^�ɃF��8xxb�D���8�O&A<G7K�ͅ�L:(C�b��&2��@@��ň2�,�|IY�=�O4�zs4%+c�˱mږ���c��:�W�XBq��XF$������g�줏N� �8�?��0h������S�� 
/?NY&��2��p�A��1����۸�Q��'>?LG�3�����t�g�1� �0�q@C���0͂>|�F���f�b��m|Ժք)f����Jtǐ|�oĊua�X������@��`��.gnf�����x'��>>>=���RV���	�]��ż�)_V8؄�ɘ+�����t��NW�X�Ñs{d� 6�lAi��m�k'��,U�R�0a%M6��.r'��|�;ޤ#�13ݗQa��8Ct�̢��Y�m0w}�W�u�FT�H�N�$�P�H�X�¾�H�HZ�:��BbU���m�4�O~�Z���8��FjD aKe�Nа4��#`4WI�!�2xI��U�׊3�Ls�G�VKH���`��ne���M� �M+(^L���O	��~z�>�����i��@G������>�}����������T����}�����/��/���y��T�k_��/e _uM�y:d�n/@W�����s�������-�=����[ �{8��<���k��u�)0��w*ga��89���|ރ�m��ݦj�k�E.�0B��rK7ʟ-���&��H����!�g��$���� {��������P���.�1.ۯ3>{��.�Vg�}��J��4͝�$���a�d���Ǿk���6���w��˺-]~������fq�f��|x��Lo�������{'<�_t�=�����=p�ǈ�x�F��{�y���>�=�s�<��o��� ����K�ط@>Ӕ�7�o=������qA�"�⻼���V��w��E�KX�A�������w,�W9��R<�V�/k�w6�4�����*�������B�`Ԧ_o�`i>�4yg}���TV�Мw}E��?�y�m��#g����7�Y�.r~0y{��S��Mg�]�vr�P@��r���c/	8Q���<zv�ڷ5���,[�Uջ��f/`<皀U�8�x��;=V{�|7O �Is�/P�Ho1,����{5=1{ݷ��m��{^���Y
\��D�gl^󻔯͛|��h��l���*�o�9>O���}~�q돭��8�8�q�q�q��q�qǮ1�q�|q�8�:q�q��c�8�8�1�q�q�4�<qƝ��6�8��q�q�8�8�\q�q�q��q��v�ۧn8�>8�8�8�q�q�z��y���5/}��Wuz�1�ޡ�x`}h>��w�|��t�-��`��Z�DRO�|��p�`��-X�������g�7�=�0��S�H�����y�vX�o �eyy�+���z6�r��x?g��R�E�~>�|2.��������w<O��|i;����[��y�`�&5o�tF�%C����s�3%��t��wj�/&�{�p�������?��j�.y-շ��v�|=�zj�#qO��O*P�!��/u��1�۽�3i+�!ޥ\[���Y|������g*D��ǹxGw_���LL�縮@���۬ʏ�'N�m3���Dz��/=8�F��-�h=%cw�ˑ;O�އ����xC/%�@��p.��L��ŏZP��9��U���qW�͒0���<w�僙�V�)���`�k�=gy�6�ԏG�*��h���C�i��N;�y����yoybs�ܛkJ��.��W5"2��{��`Wf��7\Z���ee�k���֎������O,kt��ᕑ��㪓�xe�j|�\��M���v�^�z�����{a��,;���Ƕ�>��|n�ɔs\ǆ5���n��탹��=�Fz�*�N�=�`��/.ɟa�b�|����=�D�yAt�k���y�x�n�x�ǯq�q�q�qێ88��q�qƜq�qǎ8�8�q�q�v�8ێ8�q�|pq�q�q�q�qǎ8ӎ8�;q�m�q��t�8��t�8㏎8㎜q����nݸ��q�q�q�qێ8�q�|q|�^X�W�����H��~��Do�����q%C����OaJ��-y&���h���װ糰ݓwuw}ݞ�����Yֲ�c[��u��>�e�� ./(X�m��3}�Q�����{z{%;��܍ox_(rIC�*�N�	ys�� i��xC�n�bb��f'�����;��F���m�{�x���3��uCI��s���j���O��&kOr^����^=�:Ǐ�9�>�I��}�Y~G�y�{=���b�2�o��}��{��g���7ؙeeo�;�ϸ�K�������wz�M�{o��}��.v}�M�(B�ۦ�4�s&�}������x�h��7s;o��(����:9縥�y�Aj�`�E�]��r�/����i'l���T�;�]�����C��5"�E��\~^x�����}H����y� ���=����$��9P� ��~�G|<\�v�������}g�R�=y�P���֯g�θ��{6�/T_��u�
���N�}��v6���+�x�J���p�.���OF}���g��*�7o��� wݷ%~C{i���Y�ڑ�u�vg��͕�q��.��������\�n{���2o��o���ֶ�ǭ�q��88�8㏎8�q�v�8ێ8㍸�8��i�q�qۃ�8�8��i�q���6�4�8�<q�8�8�=pq�q�x�8�8�q��q�qێ8�n8�8�������ێ8��q�q�q�N8�8��>���������~��=�����ő�YД�
��+�v#r�2B3���ٓ��KĶ�w���~y����xO��4r�E���=3�V@�q�Bt��~d,�Γ6A��;�ay��8��(|&!�)'c:����N�9V�'\�����ͭ�s�|�`՛��Ͻt�:Ytc�i#O��Pw܉�<�as���#��;�g4�W��7̼���74`�C�����x-�=��V��xüf����w�|[�33��c� ���L� !�_F�OL���P��[
�-�4��@����=�Mk������=�Br�q��X�Z��U��C(p�������!.�o�?(������^Og���v{��]��Ç>��/sT��s����^?g=�F\[�J��{���ޝ�d��j��X��~�T�@��`(<e�ɗ�0�EdΠ���L�����<>��wR��D
NjI�^�p�D{�� ���W:�b���vh7����~��j��ϳ�C�:�G ՘(W����{Yd�U�?J��^�ag��?ٸ{k��z��K��J�~9�m(��9�s�64w���ze��vё���V���\�ٓ��ib�a � �hwy���Ȱ���J3��WS�����&z-J���ct@�ծɜ�@uz��wټ+�L��Ǐ��>=q�n8�q�q�4�8�8���8�>8㎜q�m�q�n8�q�qǮ8ێ8�qӎ8�;q�m�qӎ8�>8�q�q��8�8�8��8�8�<qƜq�q����>>>>8�=pq�q�q�q�q�x�8�	ɛ���uu�9s��;5�_%v�ǂ���^�{���Q�����7�fg��܈_(1>Lq�|�=�&oJ�<o������P���}�]�&.�"c}������.�#���\;ݨ��X�H��|�4d��v�2Ќ�v�8��qý�rO�k���ݲ�{~�1�H�狓7�F������/�T����UK�}�\�Tz=��Q�b��uW���;�bG�5cd}�1cʶ]�zsa����3�&���}���ž=����,�����չ���f�6d����:�)5�Տ*�ީ�������rad��Ps?9���=�q.���f���נ�6�u��:g�(G,9�5��Cޮ���7�@;�<2}�f1��x�r�pc������>��w�T��5�Vr���Z֍�ӄ�9��<�_Ovr[��G��k�hB�C8^�I�χdھ�<@:�����n���7vC�i4C���P�f|7���xa�;N^@ET�l!��8E�0�(3�L�-|�g�#�:��G�{�$�cȊki�l7Y���2�7��+�cU J�,�4np���hӭ��MI��/]���}����=�����ƽ2�p�+�v�<�����ہ��&?.$2��ow{���M���y��r�����o�����p�\4'� �.���}��IfÞ���l^�ϲ	�<8�L�[�mbs�S���T�2q�Պ��l��| `��/^�7(��e�7ݎg�J/*D�O��3��M���0�&�ـ<;[�B��(�UĽ��7��?a��Y�yjB4��۩r��M���˨��2tbs	��F��z{�>9VtÆo���Y������ا�կgu)��� r�%[B���,��0U�o�-���c���E;u�Z�)����B0�~��'�^�{�����S6�c��^��"eý�J�r��(u�F�Kܯ`Y<�b����^^!�|O�W19��U˞�Y~���c����a����<6�OW���7����I0�OR��zN��ٯC����o��*�Wt�;[dq�Wf�Ͼ��P!fD*�{x-gڶ�M���������D�:�1��ɚ�������K��y�'�����||e��ܖΑsw�������ѡ=�7ȏw}� R���ǯ�o>2�;B��ו��&�L���ǲ,��^1��P\��wKY�"��h��cu�yw�;��w2Xzm�UF��q�o�TToG苖MK�>����&�ov�v��3˼^+�{b����3ܧ�t5�zn�<[l\d1��7�:ߪ���� ]l�<1��mŃ�T�^���O
͋%mL��/��� B��-g��ov����}�xx]�Ƴ�<��� ����',�7�|��^��ἶ��o'�������=N�+�����{ú�`��P{tu�s�bn�{^�<&��n�(�dbkN [��	���{y�ハf�1����;K>��s���v�{�B�3;���Un!�o[�7�}�\���4����D���qO�U2�%.ncU� �<5E���������:Zd�����&k���G�s�7���m�ї��	ܬM8'��:u�P=��wq�k'�`{����S�@8&{k�k�Q��A���S��}J��Y�����\���w�r�6'�%ċ�Z���uf�j(���Y���}i���{gy>��_����	��}�+��{�<۱��}�αg�:����W���پ{���j�B��^��=���s؄�j�Zֱ����<L��摙yC������Oaw�}�_�y�gk.���j��ig�s�g^�C-�����Mwt2=9�)�b��E�9�`�3i��'�>8A�b����{@u�������^ŋR+du	b�w^�PC�a޸(N&s2���:gu�>��L�'ـ}�d�z`�>�}(�6/q����y�FF��;}��kV�xo�ݜ|5��O�����J��M�v-��8��=�I�s�}�i5˚��w�Q����&��z��C��!�����5�Z��ڋY�\q��w�*�/f�5{�鼾B������q��)�+�ۏ��s�R���
��#�}�#��]�/bɽR��Ɏ����f��h��o_f�G;W٘�g�'.���O���j�`�%�}ē6�6���ma���=�8���>��=�d��{Ľ}6���Y��뷻�F�݄�]n�1�����O�D�;T��7��	�ñj�C�=O�|�A�COzv��#�_����S��e�����[^�o>w�`�1�2����S��]�O��/�ܗ��ibm�Zgq�_g��<{$�燃^-$���9�󳽑�������=3(Y�����ûZ&4����b���s�z0���=�%3{t�{�,;��ȏ{� �LK�x�r'Ž����?z��W���ܽMyQŚ�{з��±36��Ɂ͞l'"T�d��({�}}Fe����-ί����WS����
��7��P�\.I,�ū�sb��$���ZpZ {{[��S;�\jS���,G�ʎ���tK�fAeպ�~��/�ϗ$�yO>-�E扃�O|=5{������a�z���*��>�&���,�P��Rwo#��?y՝+C<���^=K@��{��L��㒿�k�QqӔ`>xD�a����z�}�^]}f�=��[��_�z�=va��S�qվ�0x���9e�狌�����v	H�9�Z�WS�O;���oLc=f��w}9����"�A��?'����Pbb�}p��|�.��xB��7f������Y;t��K���i��d��-��<T�aO9�wQD�Sɟs�]�n������ �����R4�O{�&{�2�����i���1���}E�\x�����u;��h�q���^�w���T:czqߞ���ٔ�{W�x�>�;6�����6y�+�˥���<�8w�Af�v��j���wP}����m��a��d\����/�N������_��.���é5����3};�ߧy�8{�_P3U��	�+���D1�Voڢ��zʬ�R��}�?��2n�o�<�W�q2X2 ��Y&��Y�O�h�>������x?p����=���>,�����ٕh���{���B׵��}��Ol�:_M`����A��fv���'�\�Y���A�4��xsu���g�����7aگ7�'���t����=ag�Ǐ^]���^���qU���Q��I�=�#���N��b�ժ�rh!�#k<wy&��R���@��=���K���'��>�sL�[��s�I�=f{)�s�oj��q��(���{*b�}��Y�̔K{��x"$�76�q3�ύ�\Jzm;5���A��gK9�㏀/�g�a>���xcuMm:�4�{
�F����CXkzEv>&�b�(o��������e��r� x�=��Vw٦S�g�<���̬��!^�׆i~��Y7"~�g�y��L�s�&�V4�O��S��jw��=l�Ɏ��z�h�qZ����\��ܢ�G�����d���Y�����Q�IǲE��Z/[�M�%r�������y&����=R_{�X>�����H�W��T-�������s��oӶyf�/˜��wG�V'�)��6u����������=k�:��e��}��Ɇ�YSjw��G��׺�Pv\���Gr��u_R�m��o���-��:gy�n�N�5���h_[�W��юy��8��M�p��ғ���kGh�
�E���y�J�z�������P����$��N���4m�L=�{��R��<(�;�:zWG��oq��w�I����z���Q���uZ�?a�=y��
�үg/{O�u�Q�2�Ӿ^���ɜ������E�H��/�~_��?�Q�o��u��j�-��\���W�5/����<KSW!q�ue�Mdnk���y�K)?����}z���`،U�
`�J)��"@P��7�WWg�z秞yO�ͅXU���K4i�pʴ���v��PŁv
ACql�h�l�0MrjG:��,�	��  ��6�%�
[te ku�X��UAŘ���e�� �v-,�.g�&q�Yf�t�v6-�Di.�\�0��E��Bl����;q�1r���պ���c`0��a���6ul[�bL�3J�.�u��
jW1,ً�����rYl��f-M4%������Q�JV�h-
�uD���e��0�V1�����k�R\���J�c\�deY�7��{�-vd�e����\K-�[-]����I�u��[�Q+���n�&�L]SK`�3G�fuF&��t���E��:3�v�� �A��s�P���[��If΅+D�`��棖��j���lYk0r��c5m��F�֜B����ѡ�hg1�Yb��h(�vlZF�M/cJ�I�,H$�]a��J�J�%�1��KwDҍ�5\ˌf�C�b��\�M+"Z��RX�t�:e�P�p��b���r��ŵ�m�$k�v���U�$+����m]�Lۭ�x#�a��j�Z�KH�f̄ �RLb�[�����1��^���ݰ�[��-%v�0]MؗGp�͊�!5k��A�1�0�ť��ae��WX��n��d�F]31XZ��kS8�������DilTt���B�qt���!Hrk2�W#i�u�#����]� �Xm
�+�63c]lo[�Z���npg,��k���2f���\+��48n��VhL:�`Pؕ8¸�dU�{;k`�,��m^��J�D��հ���It�0B�D��g�vfb�<JKf��)+��X��8�'Y�fIaf]2�mP�M��Zc =�hc,��z��Y�6ٶ�0^Hؖ6V��5�1�j��Y�4��eLc	��qY��fB��,����Ii��5Dڳm�q����5֛"��X���Ü:��V�;Jh"�c��&�����+)\��Ҧ	T�&B�!sqv���!�va0qZ�.��	h��2�%M�Ҙ͚��PvR.01k\X��Cj]W���=��!�*m�K6�ck�c��S!n���q���[s�v�L�I�7nkmN���B��&���Z=�3�!M�A�\�W�bQH�u�h�j���[��6��sf��l6s�Rk���Т�Jͬ�I`.��]��.Џl�%�Ě:]ma�q��uy�L�6�M�j��3�)�q+\��Eb#{�x�+YI�Z�ˁ�D��W1��Y�Y�4l�2��M�ir��6��v��:d��	�� �lihh2�L�+XrF8���;&������f&��V��\��m�4uZ�Y�b]�T�&,,��4��H�͈٥ k�{lR3``kK,�V�+�f��L��J�:��W1^iMP��5��q�*�ɊK�eI���ј�rMma5d5��!��фi�tG��]�Z�M���*4H;7�͡3+f�KvH7@�ː�2��7Z!-���8�z�G`c�XCP�hJ�e��� �]��c�յ0��#���u��[�Kj,5�n��B,��Y0��Y�(�F˥m�Gmke;lwZ�XU���҅3����d�F\��cGu��n�4�)sx�j�궓f�k���ga9�(�V\���M��Li���豳Q(��C�9���S�b�[Fkrـ��m��%��A��n�A�6�1��r�Ү\�X]�ծ�p���Jhm��ť#F#5�`����3�&��䍄JD�]���b7�IZ;#X�	P�Ό����$��m&��ԌGf�Cn��)��:��U�,XmSD����h�P�(��Hn�4��fԠ[^K,�����Ą���,��30�i�Fkt�{]4x�h2Ve	qscBhk&�f
�m��xV�eGpޭ���ָ�A#�]�f	��(�j�ڦ�U��:h��wW5ZZJ3R�,f�"ˡ���X�n�h4�5M�4�cH1��m��X����3L/;%u5����]����7;u�Y+*���Zr�R�鳳�N�S"1c�mڃ�/0�ْl�4�xX2�k���n&�b�b�e��*WB�kں�	��E��a���
ƀ���{Z.���j&�qR�&�eY�����m[���:��s	��ֈc[b]�[B�5&�6�;h�f2�tn��˜�m��Ĩ�0Wp�U�X
&�e�-�V<�`[R���@�e�`"M�r�5��-�Z�!m�.��;+�����T5L��,3�m�EJ�ã6�)�2��Kq�H�:�a�af{S$��H�t3w3ephܘI�RXWBPw9�][���Fs�B˥&u��ǲd�⎻F	0�ҔZ-��ڱ�8�ݚ!��붘�8��������f׈G�ĵ���JsڨM,`���u�v�YRd!o��з.��Y�j�1�Ԕ!b�bZ,Z:����ҩi)T6�Zh�*b�-L@V�qHD[c��A�,�n�6{)��e�(]�^��#�5��8��5kv��	�hS�4��5�v$b��aH���ʦݭ��1����-��R@���UY�Y�kFͮي㖽R0��eSm]���V�X��i`�݈A�kY^4{-�C&�e���!kj,JK#�Q5t5��Vb:e���͗K��5��Q	Q�m&�#��ˋ��b]�E�2��ԅ�P�t��
\\�-��Ɗ]j �5-��t����U,C�6��+,5���1���6@�٬�6�h�Ձ�$#j��Un�%F���fg�t%�.�V����(my1n���vu�%j�b��5�g��ط�mj-���+,5��%k.�b9&�a�4.��G���C��v1+s�6kRG���K��q!ŗ��e�	�!K.4�K�`t4B�����-(NTn����3l�k,j$ثqu��Q�qc���8�0�:,����#�E��en��)iN\���B��������7:;Y��	�pY,k�F����n�4uM�si�]�i)���]-�	�P�A�m�2LձB�];m�!mx(�$�6]�ɺ���	�8��t	�bT�^�F�β6���st%�Hꊁu5��kl��!���@+i��aC[�Gem��cKD8�v��T�%�ǖ����)�؍����VS��	)�d�t\�R�H��[{k�H�FJٖ��三t�L �^���l�#\�l�]��ۥ+7kunq)��՗E�tl	��f���T&�-	���ŨKc+ep�`���h�� �ݠ��fG�TF�e����H�9#��%8�݋(����I�:����X��Z�9i�nf��B��K���&�%�,����S�����`@�HA5�]N���&exk�MDb��Ll�0�s��*lY��
�5F�J�ңv�1.�J�	r�]*1��m
�=hG��H�Hn&[���]�n��;j֚U���T�.Q����[,&��M�l�5�� `�m29ڬ�һe\- ���-)��]�F�/:f�ڰH��ųR����L`�Ŕã�Ʃ�,ژ����' �D��rl�������YsQIBe���X�kr��]�
J�CE�����X3�����kB�xca��f6��Ǭ��ڇj�1sI�%�Ik.K���fRi�u�V��%dlj��ţ3�F�$J�X��l�a�K��ۜZ&�$�C�M�4li(ECca�,,�i,1�v�Q�ᖍ�Z�ꨚ9�@�k�T��hV��X��%�`� m�(m-�q��i�f�f���ArZ�S������v�@�!+��%����en#D�f- �A˪�k��+���ۖш���[H.P챲�[fn �����z��Yv�t�*ld���92:�6ڰaV K��0�1�lRg,��D�\�gHK^h�Q�Q��-�u
���[�%6�8�bPL�0.ɮpg�#kfn��9BҴT�����A�Z�u��1���mŽ��j��L�p	K�r@�c
��r̽�M�4
��xR;��XhJ�b20��30�2���F�[-Q����n�&�X��X`�ʠ����<v���LқhRUp�d���i
-�pԶ4K��e��!J�!Qf�)j��4j]c��eʽje�f��H�ي�]!*.��k�䫰K�iM
Tn��5Q�ub[���s�5�.����7$qb]�\ICdi���0�f��@ت�0l�۶Z��J��e�iWfQ2��UUT3e��̹b��c1O��>>��[BRj�]5Ϋ�֌<P�e<n�ך [<{Kb#a�!d�y��F`v�-ѻ
<4�G�[璞P��:�No�Gma�|w��l�aW��5�
 ��E��;�,���+vŏ�2魾*M�ޑ7�-��� m�lx��f�Y}y�@JBS$J�PDU\���
#����Uʢ-M5�B�z��Z�Y�f����}�7������㏎<x�!�%,dUJ�'')2�UJ'"�dU��^��'6m�¢-�ox������q��<x�h�� (�CPK�W��i��"��M�E\9�}��Q��ǯ�1�Ǯ8㏎<x�K�H��P��	:���ye�:�i*�X�o^�Z��rMB�"B��qw/#���تR���BT͔��#$��^�z��q��q�����g��JNj��e��
�Y�<8�2��p"��U� �PT$XL)�N]���CF!��ڹ�t�۸�9Ls�y�-���96�a�.�kEe�c2]��t�;j�
:�B����a�3i�g��rH��@�E�j�5����&���C���:��::�lww<©
{{���aI�I�a�S^�k�:�fT�k+Q,�v���$��(ZЬ*r//S0.�P�FNy+J���¼�L��C�x�u��O�rr�Gq���v��*��ŕ����� ��48\s*;�Ϟ�HyҧD���$�U� �"�Ȉ��*(�"����%�EDȠ.\I:_v�IaA�*���(�E��JI��@�(z�Y���W����3���@�K�e��
=t#y���pQ�����A�l��\]	a`Ѣ#�u���Yke��֮��BdST��д�0Yn�XS5hn�3&f�GG��������]+A{$T�gf!\�V���3+��79	�\�5f�SZ-ԌEIRm�H̩r�nY�ۀ������;E;e�X�i`��c���VK�z\���4n�J�_;��h�K0���c���+W�!��Z9��\�%�RV�\��ST2L��/YDi�rԡ1�V5���\@�-���\�T�h�KΔ�#0�:l0�*�tIG+sS�E��#��j��XDЌ!f�me�!��$�$o9��Xచ�ĶИ�*T�Eseњ�I�k`�XBl2�mv��r�:ܰ�Ti,ű��� V���u���ۥ�`P�n0�(Mr�)nЍ5G�tA�r���6���\�Xvb6*�f�89��xyHP�G	�C&D���,�w:9D�J�vp&lK-e��46a�V���Zv�SHK��̚Ý����i� Z�k�� &��"�X�V������<Q�T$-��l��*�pcP�-̦�q l5�IoJ��7j�Y�i��b���7\
��Ś�n��	��R���-Ƶ���f��4݋4l�:��Mͳ6(&hMb�JcVikj�qH]�[W�mmUZ�e���[c��;L��i���@���˧�Ǟ-���1,M65i�-�Mv�ٶi�&��n4�pԔs��-�֥W!*����n�����h�Z���Z�����-.)�%cva��R�v�������n��M�6�Hh�Ń�o�e�k�C.Ί�DCGYYB�v�
�c	tb��\ﳺ^���>y=�[Z�B�M-�7fs�KK���w^�P�(���B�y������\/L�(��ۮ^���1��Z�cF#
,�(�-P�שYB��JEa�	x�e*��r��]C�v���E^!�	V��l�����eHV`�J��0DZA���J	P��cJ��-(R%B
�R��ߟ��_�'P� |1\a�A���A �����k���8|{0��!{�B�m�ÁX�ɖ�T����3��}�u�C�L�&͌��35�����҆W��<ߒ�ex�q��L�u�-��ҡ���	�G��[$J���I��hk����B!�N�&��m�@1�w�{�YY�y7,	`}�ْ	b������EV����r�=�$���d:�}
��{n�X��v��U�d����� ��1;�jC�d���+A��PG�_��C��W�2�H�u�x�`���� �f�o#�D@/d_��M�����Ll��t3��,	��oETm����/ٔs/$H$���o5ɸp��N���w�u�X�{t�Fb"gpo���eQ�=�;���1�{�!Ɲ�p�o��R���{',���g��]M���5Y�i�&gЖC�C5\�� H_��{���9%>#��{ޥS�X�ͣ�O-,� ���3�7{���>xU��!{d帀I#=� ������$p`H6�U���!ËvY�y��:����4��׼�>y"�o�5����zÉ��)7�ǌO��z��6�ݦ{yvy�n8�a�F�p �/gdNԘ����L&>J�H��U^��0��f4.@��iT� mE�ȵıQ�Ѫ��P�4;�*����ē�yِy>�xc�#n �e܉'[]��5�I����}���=���������	����AUN�e2;���y�5�נ�<N��AM4fH��rr 0y�Ό�y���:SS�,M����o�s��~�;O�S�cK��ѣ�{B~��gzx��N�t�xb,]-E��B�q��曃	�M����2�(�#[N�F��s�0$	��N��ٰ�d�\p\��q�h�S������bSk"Vy�I�NL�$K^F��O�X�UY:�;�M��l	c#&j�d �k�0+�ک��T�,��LL�4�|�eN�H$����[����W��C��Ym��R[������T�-r������\c,������>��U�������[�P77�%��	D���%��Dk�L�*FO��i��<�L�P��CC��Vk� 1�f{_FeD�3	30�u��I���52ML�uژ��Z��KC�	p���N��5�I��0~���?_,`��j� �}�Q��D<���Nn��M5�<ׁ�@0M����i�����QxA��>��㗿<`���+��8�����=�]���CʌI%�NX+O�F�Ӏ5v��v����5m�w����U��ǗG�ڕ�l|33�&��%���V)ckM�|lS0{�}k����|��k�p!�&�r
$z�I�>�cW�5�m6� ���^��o�w���G �+e���P��YjhJ��r�׈���S�>R������V�[=�׿R$�x�]�� ��}0sw%�!Lܚ&�$	�&�&��#[�4��<B)�ǽ�y"��g����ﻶ��Ie�i�$l{5�:�^*D�y��r���B�{�����G�')�#5�@P�H���N���@� wT�Ĭx�?)�=����c�L��/3�Z�ı ��Y2&��_sN�1H{��d�;�˼A �O�[�p� $�ӂY Hdܴ驣26� �1ld��f��qU�-5pϏ�3*k`אwʝɾ���o�:.��\=�Q����Ǻ�w��ڷA�^�ŶP��차>��߫�\������9�gFQF��8����6> �X�5��o�/�ġ$�i,l��H�J��]0�AIm�3U��e s�ԭ��_��/�9��,�SHJ�nU�T ���)�n&"�2���m���Bc5���t���Cj��p��m(11����L�U�\���2�ƴN%���lM`�66e�W%��J��bmuA��biqcDn�ё�-�*��e��PqVb�r0P&Y��Ɍ�#��qd������+���gB4�ZEkmeF��^i�ZK���"{��<AL�WK�$���v 8��qG�>���	~6�3Ć� x��������rdޟz��ٶ�i܌��|%��B�ّ �9���.c�R"�En^<�S@9}��D ��Na�{�/S�ZO�ȉ�����)f�b�4����
l�k����n���kS��� �I#r���,�f��M嘟nUf;Dx�_�-��m����'=x1�dI�k1���T"b�j1�
���b�����E��78	bN����R��u4�B���
�1Z����[M���x� a��]^�ǀ� N㽑�g*�K�R�rn�5{j��S��-�Y��u���0�I����Y��D�옆4�J�Qch�9�qs��g����}����w�͈�~8��=Q���F�;}5�@������y��s2��N���T��c��u�$�݁ا�[�9�@�7�PW��z�p�� [�ṃU�`���hd�yL �Ym��p�H3s�i��L@�	��^|�@*	��5�Qz��/f魒.��5��"���ĝ���^���A�}�N5S=6DGQOT2�}{$�@b�k�z�ʷ���*��d��!�B9O�<���k'��I|'�5���q9�jTM����h@4B/�%�M�%��ȓ�.��D��w��q ������D�Ă����X���=I�מ�N�;��,������gI��%�>u^O�s|�I>�q�����V,����ݑ%�Nej{BB�a�x��ڣc�̂�G���sU�w�T#��7��z��w����;����)g����xgc�EAi�l�e�0��'�sތ�4���*mh�"`a������ �`������Q��3�;�E��Iȧ�X�%Y� mYZ��bv[��kg��DD�%WXf@7�ٜ!�z[�)b�A ����H�ݸq�D���/^�w1E_�j$��x
��m��dd!�\@��3ds��q���ݝ�mdf���J"�
@>�x$m�q�9��H>��}��ޝ���I�{"���pz6�%c��ߩ*~�:6�}P	X�x�Ai��Z � H ,�Aj���⿽��#e�v��� ˠ`����	�
 $	��`�$��ĂX*ݞ��h;j��Qם�j�]b�B�PaǼ_e�����s��چ4��,f��I'3`��EdV<Ml�,�q�>œ¥�����}���v2�z�����p�VvH����L��7�f�]�1^�{�Y�0A-:�`歴l��r��&$4�3$���1�[�Tz6��meY*��,�ݬ�ݖx�\2r�p���3��%���mS��$����(���Pdl���h��(c���ٳv`M7����Lu�>g3��$f�iD�M<4�р@�)��촜B��)D:w!E4KPYZ�I����͕S^����(:A5��� ��{� ƼU���>��3�'N���nK[�
��.R�F�y ��ِIḿ���k�0�D�&�-�}��T��E��D�I��C>�0�1��a����ii�-X����xNTB�4ce��H:k���d��M�)g�3{2	��0�j��5�)�Ʀ�TCM>�U��>d^@�K��ck�q�⴦���=��jb�]�8~7�ؽ�j�{7ἱ
 �\ы D�����I}fk<��|,�p*�Ho2��\�wI�Hjx���c�rA�cXMoh�+R����F��\ěTQ�d�&5	��m�� P�����NΛ��5��9�j
\ѥ�Лm�j-�P\i���p]A���Ұ���i(�u��
��f4�&n�[�h���1�,���$�CL1��5A(�ṇl�0*�(����V��TEqe� p�6r���B�Ƭ�,�merPIcpj�`Bi�Yf�U4D�,l�A$�F�^%�A��bAy:�Z�w!೶��!�r�+=�=D��e!5%�� ZjX��!á'L�M�����25�ۥ�ŧ2��$eMy$d�����_�_sH�2ꎷ�^���P���(�I�C�|q�`!㐄1 ��LD�#Dz�� H� %���{Ib�����b=��w3*��Ƃ�tz��	7� ���Pd6}��J���$;�%�ކ�a:�E#]�T�A1���v�l��yN5�S�F�b�"NN̴���{}tIbuAw�x��h�3sK�2i�r,�mn�13Tc1���T6l����}�L��Y����3!�[�e����ñ&�)��ܕ�@m�Uk!;�Q8����Q�d�����ߺ�Y0FE˳�f؂���K�7���3ҩ�(	�F��e���,
_�{�'���W���j+W���`�~�ĵ~ ��{Ps'6d�s���^��o�E{| �w�5S�x�R�A �fȐAԪ�����s��%�YS�P�j��3�Xd/�Z�&;o��9�7焍j	�JY �2ֆ�q�ҽ'VV�s�g����r�Ű�)�ng?�?��@	&o`i�N{լk2����� a��}� >��L����?,;}��ǉ ����jU�]�g�hk4fb]^���tAYn�����G�'�_���u�M�C�=�4'Y v}q,I�k�t=���5xJ��	������<1��@�^[��"�G�Ϙ3F;�x)�y=�2�ޘɐI#3a��jx�y.%�x����q��7��yﺸr�$i�F"����W�穅~,������V�\,>�;���W��z{i�|�N'���Xn8���`ݏy����{{O��wޣ���q��3��g����;~M{m���ju�6���i��d��M���,����h�F��V����o��7-Ʌr��5��Û3_�M�5���}U^b�%���M]��_:�>�}H�g�b���w�Sr�xzt��l���ާN�x{�c���W�!��]YJ��p�
t��v�p��^�B��wP�}F{D ��Yi>�y��-mA�-�L7���W������^�K>E�j������I�8�/��V��:O�?L����{����3��U�sl%�4�=<�U��w�cf?�p��Jq�a�����緔��|�������mo��oT�>H�a�����3����/-��tr��o���'�}�^�}�o@F���w���bާ�3��w12L���s�����o�tvo�5��HM>���#�����)��}��2�<��;���|��n����kӛ�}�l��[��8���{�/vl��y���{�b~�_��_���-�v�/Mͤn[���x���v㾒�Nq2a�>�S��ኸ�8�X���P#;sN-�RHmG�;t9��	®{�wp�=��\�{�h�2�����Q	�yn^Ƽ7ۏ� ��r5��\X���:�6z?w��쾀k=�J6Lۢ�����&���/���(E%!i��%����!:nt1���O�X�����}�[� һ����>�߇_x�A���L���Wϗ>30�(�����^�&���L�o��q����8��ǎ��	FFI5*L�`�ȦDf�EP@s�ȲF@�Ԅ��ׯ�=}=q����~o����k��Y�%��9r':QDUA\)��t*�jвBHI�1��ׯ^������������ǎ�E�a		$cQ���EG*+�Ve�U�T�M���Js��"}�w^��>>�q������Ǐ� BH�%B���wZqE:E���C5�DQEV�@�&bHWH�iq`�'{�
es�L�B��بQ��T]&�?Xz,�)2�Qd���P*����2��Qp��qP
������er� �E�SĜ��.\x�.��_�H�*�
.PQ�i7��U��tev�|eUI�.TW"���YA@N�(�A.�L�*���T	�E2�"���I��$ΑG8E2 *����;�H��W�s�9�M�z�U���T����Y��RDE��D%�&lw<o`�P �"�6����[��!wEm�6�ae� �����{�Dtʉ�5>e�ȟ5�Qi�2�.���}�7d���Z�,@�,!ݯŚ�A)�6s�
�ei��	���'f�sߗi�QI�O{���c��;$yΡ�C {`���0C�\q`<�H�@*'�r�	lZ�h��CtGB,$�E�C��x���$L_���קu���w7���y�n�L�;U(`�ԶYKGFh	��\���i��5S�������}��!�o^̀y�
��eB��ϛ��!P"PA+����&�A&���6��U|���G�*j0u4#:`1,��/`��V8����l��S�"51r��C"zgVwTO��u�\�o漈n)"xiD�}��8�C��w��גcЄ�:p^_^��dk $��~,��+�z��*!@��!��@�D0�Qf	[F=��O��÷�M���'����j���T5��C��Y��T�|��qjJ�Dz��_n��$�df�tC�91�Ć� ";��@����7=�qE�QcC�;����Ӄ�$7	&;�~�&=2bgb��O��n,�Q��; �A���=��]|}��e������|v��nxa�s�d�q�Fs<��a4/;]��W��k��X�`F���<`���eT$S�v��AF*�T՗�>����s[�H� ��;���O @uۯ{��VE!���>�O�Fs怶 ā�V���Y�O�����k�A����⹂|�J�L�4���P�ep�B6�a���ʗ:�cW>b�z|=}/E֙~�䨗�|���RAd��m�T�	P��B��5��Ț`�>OgϞ�o^�H�C����RE$Hk�y!��/	k,�xF/ ��r1*���"y����k�/Z�eO�9�2&��[�u��J����w*%�4ME(�3�o�!��&�54Djg���w_(��(y����A�.<-�"��@B�"��u䴙b&��@�-C�+���m��6㥸���������s�������bI�Ę��}�����a$���\���ǈaA�4�PPxx.+�0�� `�=�����m�0A&`Hm���\���	���T)����`KQ "Ȏ��������C��k~y\����%@�����nD�m�tC�91!�LX"7�)3P,(�@��@���_-��7��7�&ך�D	# �
�׻�{�H����"�ͻb��(��-�=�XD�$F�&�;�z��< z=�UȎ�:�G��_�{����w=���ip"ׁ�@�����>�4�vqSu�0���?i�L���A�'�q՘dM�UW[�s��F?�M`���4C�%��s�'��i�ۭ6*�]�����6�m�
U(65ыfB�MfM��ZKa�x�A��̔�.�ԓG�3Gm��Wk(\]�٪�e�F8��$���,�6�B���lS$`�j���`�vpl�1M�fۖ�f1�Ŏ�Ȥ����K��g0&Y�T�%�
�6֎�uh��r;du��4C��<	�5�]\7F��<�QX�kZ.���A��м�B���3�
 '/40�>#X��\"�	n4��j9�t��y��Q`�tt�D4���!�ރ�vz�0�\���ul
�Tj!P�y��)|!�F����rC5w��i����	�Q7�˴ܨ-J|��2�7~j�9��d���QI�JeC���=�<��� �����q���P*-E��=ߵ����L`�JǛ��+.K�.˭p{�ƓP�U�PxD�-*	P*'��p�"X�!�aQ��ƚ��;�=G^��u�*	A*)!�k̤<�%����$����EC�0E |��Z�K�N�~tp� 6�"�!��(���RD�5����;"T���|����+y2�4��y ��¡���)�=�oO�����FG��k(���C	(�Tm�01ޓlO�~�N3S�$�[<:g��QXFJ�@4�LXYF���v2ȵ�X:��>���,$�D ��j�<OP��%�s�n��Tέ%�-����`F�+���@pMx�.ԃ*( �;�9!�B
��Ć���[H
<�P;�]*���m�Ad4Ŝ����q҈a%�}�ڦ� �u&�]J@.ʃ��.�H�'���+�.���P�����t]��T)�V�����툍O�o��h�So9�۸�B��Y��.~��&�t'��]�w����"��T�����ۅp����� �i>1��3�JAq�yw�ו�|n�o������3����D�Ly��SL����H
�g�q�$c�9wv1"+�.��!�(%z�dH	�\�7���x�D�izP�w8ˡ<���']�FD��%p�蘁	�{�:�9���Ō�6�D�*�No1adx0H����"@K���RN���=+fa$��j��,��Hj�Č"��@B����GI$�=\��{�A96���f�Q�0� 	 ��L�P����
���Þ�N'�WsJX�}��,?�$� ��,ԫ�c�@гm֢�-uV�,X����-,�����������Sj�_��E��|0e$)�,�ʩ���{�8=�fX��C��=D�|�26�Ƭ�NHw��&(��|�g�^���{��M�f�k�x�0�L��� H��b��:�x�B�2p�u�B����м	`�d@wxF=@�2�E��du�;�?���$�
�nt'�Y�a�~�u�ߨ3�{&���-ǯ�y����O=4����b�f���_{Ӫp�c��h���~�<5�t����@�S���j�h��Ƃ���~���|�	 �cL�E$���@U-B�����c4J鰺���݀��#�H��[�.��*��{y��8N�鬮���K�dI�0�����+���O"왷�@Il)���#���ѵl���w2<^e��t��_*�H���F�ע��z˻��V�+��[v��V��gV�eH�4�
@�G\G�B��fPEvgjFQ�8����$Io��4%6�D�j�TL��~�f��rS�r�i�'�T)&���6p� �<:5v)�x��
Y��1{�Bu�� ����Hy��3���I��k���מ�_xWEy>070Ԣ�WNN����PY-`���I���d
�׉	 ��H������ y��W>0L��tU�)�IgtI��KlO�& ;�%��z(���k�G�0�)%8���,�g ��ؓ!$�d�q�{t���:�5��멤�n����F�\�Ibi7�$���,cO��.�?����7�༨�D�"Bǅ��~���e�Y΂v1Z�u:��ߟ��u�d_�+"��1"n� �?DJI"}�@� &�Q9`�fXH+��w<yN�	+܉ �kg�;���,%lV�����	Qtv}D�I ��%�K�.�!ӡ�6�.�Xn�IB�䰙�Mj�6�8��Y}��ϓ���n�s%8���I�,��n�JD�H��ڱ��n�.��`<@^|m��^oS:t�z��gw����$TD'<�O�"d�[�w�{Nc3Ws��P�,�l���d$@&��L�d�����+)Ӓ,3T��):�C3N���I��"Y$I����d�N֯TܿmA�4 ��o���lw&�^�#��&e��u�8E8���c�d�Ou՛��a�f�	���x&�I ��D�I�Av�r����#� IM��$�1T�ף�Б1��(�v��"d�$�{���޽���ݗ��A�bL��@.b˳ S	E2LƵ딛Qכ�ǹ�,V�ʝOn���E<F�ڬ�0s��ĭ��oٱ
ex��1UO2��k�AEN���>�Տ�S^a{��������[z���M7�y!�o�7]��C�頩"F�F�hB�iT�#"�!�8xp�Yw��p.�6h)�Xͳ���˅�f�M���6�[�"ؒ�33cA�Yh��\�b[+�ĽpG,��lF�E�L�mVjJ۝�n��K0��B�1�SX��K�Ё��C9�Ύ�c�L�F�Sp�v����pQ�h&�h�jdn�@�o6��]pVS+�����i	^4F������ƚ8B3/l�r[D#�w�����y�27�]K7R��]��G�"��V�Y@ɲ?'���Ի�}��߯�c*�2���wt�wG�E2⼋��j^�`����$��
Ao�Dm�>�	p�'��Ju롞i-1�M�j`�b�sǒJ�:N���wd�g�\���G�ig�����>Y�w�ؔ$L�9�/���1"��������ع�`��]R�$�Z��fW��-��*��ךl������ܿ*y�l��y�V�3:�	G�̉I4�]�%W�D�ws��Nt@��u,�Y�lI�)Uc\"�BE@1F�]O���ZI�cDf����>5�*7c �}�s��@g$�=ę�����?�SR$�3�wT|d���h�,I��	B� �-���S��X��R牭�P��`�+5��mk���ٛ	�"��.���ۉ3)6;�Y���RN���_<vqa(i�zߍ4�)wEqeT���x���p���LTw�- �J#�G���}^1x�~������ET��x��پ��we�'�{��=�3|��r�zM�6��uH��w����߹U����ϸ��H�cM(ֵ�Z��HCl�˂�Hg��J�H�މ�T�I�����I'47�Z3�]��=�}{D�����E$�.�̔���zIDׯ�IWRFO�7�\g�Ƞ��z�B� 7y�͹�W��(���O]Q;Rf�����F ��;�W�ݰ��,�W}d�����?<q.;9nJO���@T�C:I�2��/2n�6I}&��e��=T� �d�zԖ�
������_�U�6���[�����:-��P�-�vs��VD������w��Dw�`�B�z�9�U�-\�\Myh�X��Ѯdj�3X��N�ڗG[gϞ��p�q	rc@<�u>U ��A/o<IdRH$���H�\9�6s�i�|���2����gD�d�����P/T@�����}H�gX�������@M��^�x�$KP(�R%W�_U��E<oV�q��	= ��'�x.��DG�Os̄�%$�r�I�	%�����N���}�f�9i��ɞ�)����}|��\��^o��sx��}�;+���Ϯ�4��̬�t^��i9\��0-�-�փHgZ6-h�`�\m��� a_*�� �{��%�;CD:��P�ٓc�t��B�x���1A/���m�9bɒIO��|��I.x�@:I �DW)g�yVBk�M���/3�:]=e ��iNQI��B���B�"R�*�SF=DG��]y����&ޘ֠	J�꜠�;��b�I�vc�ĠA���}��y���[.��r�Vl��j��RUIj�n�	S�\�C�1��#B�w3��f^9$�lyh�֩� �I7lW*-@��&���Sv��v=ʔA%����͂��s�S�(C��I�y�����A�$�k|���e�i�`�2� 󤱝�&��RH��".#ܤ�C8
�Fџ>�oE�ݗ��%��삁O ��yzT6Je�qOI �v����q��^�8d�d��~�a� �����ҦQI%�ʅ.
���.�B uЛ֯6�5/`e$L+�-MN�'wt�cت��4@����Ro��7���u=�^��Yj�����w���hӋ#v����q��os�����	O���t���
���H�;(�T�N���Wҁ�G�V�kִ �،��`ʒAc�  ��2xc�.��(Q^�K���4��â���Hwg��j�(p�B�ϒT��4�zg \.��UH�[���e�a���tl0�\'p]�!�]��Ҧ�vH�.yf:
�fe�r�36b����¹'�
5�(x�"@D�@�׫���d�k�Q^ͼ�B�X6���R%� r޵Us��ޑ��т!D'�)�R����Y��XE��yW�JL� �ثUIs$��Q �%Uz���E�eu��G�k�S�!��a)��Pp)���~�tH	)��6��O���@A2�,���I$��$���!��@�b�.R��@�	�z6�U�hI ���)��.��^j�$-�'��������	�]q���-k�6�'tZ#�it�.�I��T���\)�� ��_<�L2\��}�! �Is�.iPS30���n4F$�ڪU/U��O�� mZ������3ރ��fɝ���_xg�S%���B2L���7�F͑��ї��ޝ�gs�edqA���&� `=5\W��)cܴ�nr�i�/� �os��I�0i}x��y��73D��hlo�o���U�<�ry%}�����Z�~��U�G�mv�@�+�9uL8�x���{�Q=�]��ω>�C:o�}�����}�/������m�r��{�ur<�1@jv�|���kZ}w����"�6t�0�9���:�Q���@����4���&u�*�k���}��x(�o��#�X;���n��/v�yp+�@ͳ��/yj|'C|5�����/�5X�Zn!{��5�>ݚ�,�k{��Ě�=�o�R�4t���N�3�HdȤ8̡��c_Fx��5O}�}�o=��������سs}��D��;A�7E��r*��n���yk�/���K���L�&��|�x���{w�Y0��t�#|'��M��ҟ:��,�����ã�0��z=�{^��^�6'�th�8Ԟ޺u'B��T��:�B��}��R��}���%�����<]}�1�|��b�/On��»^�C���x;��L�nM#�[�9ة�'��*֙!X��-+�h[��:{���]<Ab6LWC��a�D{w�h���� k����^k;}E�3�����MΒd��EDhs�j����q��5`�{}vQ8*���S��z�>�o�Cs:�ue��^/y�&S������XbpC�84Z���HQ�mތTx��J4`�9H�B"Az|���$-���in��-O+�[<���2O~��V3d's�N��fA0v�3�Ck,����i�0c�!ޘC~-����j�E��#�)K�<�x��x��w߾�.�M9Up��6;�(���29d���kH꜉�� �o{�}޾�8��������׎�D��!�*�
���$��UǤ���9Ȋ"
�4��_w��{߻�<z�>���z������!P�dAr$�AeQ���P$d�$$�����^=�z�8��ׯ^�u�RBTJd�$�Q�r2����!	"H�HB��u�ׯ���Ǯ8�<}z��VI!	$�B��˲�hlJ�eGN)�QL�z�����d�Tɔ\#�*�jh�'$#�T�DU�)2N��D�ZDE�AI��'N�#�$%UL�<WD��&��9Re�vS�wN�F���ȟ�(=Yp�p�k �� ���RBgi��EW�FHqR"� ���L(*��'(��Q(*����4�"�G(���<O/�8�;�u?!���vq�,{	�F�V�b*ō�ҵ@dB��i�����d*[R]S[�$,Θ�ΪR�Rݤ����p�m�6ve���^��a��ZH�"ʔ�KKGG":��KX݇���te��h���i�؄�b��j'&�3ei��]�w-.��ѹe����R�I��˳I��.��Ȏ�<f�sq����6��F$�DXe-�֖��W`s3Y�Z-�v�v�j���b�.H]-�g�)�ڸ��#���U���6�-�[�U�)v�l�W��Mf �TY�J�W�b^�Z,���1)H1��6]���M�VhC��y���-y)m��(KYF�J�W	Q��H[�A�]ei�YLA�t.�\L-�k/j��n�:�-^�JBR�۴a����׉�ڰ5��J�:rm#4&�E�ō�[-'�i,S/f��/V0@���嶠��v�˻X���-2�-⮇n�m�Qf5�HG�q��Ћ �P��[lͅ)K4��0�eW�J=Az�%]�6鰚���FӐ�5Tҙ�M���:�kb�.(���m+Z�x�DDH2Ő���3�GF��
�ٵ��j6��Km\��.[`W���CJ�sm�ǋ6Wd��{�Ӂ�(��qR%�"�6R�� k�34�雙s�c�%C0�fkEv�mx&V<��l�a�X�`�L@�P՘1!4�.��صqy����ڱe��m�Ѓs��SmB!Pz�G%����MM��e ��Q��%S=tَΆ	��Plun��oiM���v�4[lԙ5���T3X�]���TK�g]Kb�1�vv��+n�.#	C`61-Sk@�(�y�;eݘmriuY)�1�U���M/^ܫ���ܚ槡��B0Yq��c[e�w�� �|�v���\y�§'�6�~��iu� gZ��k[lbq����������ߨ��(Bցc%��M�{Z��6�F#�m�E��I�
��-�ЕN���[I`���V	���b�c�nj�夬̶���F�,n[vHS=tF4�(k`1��B�\�Ɨ�T���	n��B�75q1h!�u��B�٢L�"�B�&��Ѧ��4��i����hU�Z12�����5�.���y��˶���Vs��m��Ye��,sk񝹶�� ��K�9�������� K�;TN����ؐ��dP��UL�����b��Le���H
$�e �:_eJHu@/��)�%�	V���$�����U��{3<���I r�D��׾P�Q@[��G���^�/E,����IzE�X���U�`r�F��<� e$��u�`!�3��yܲ /Z�R��m��ܐu��W�c :8���n]_�Y}Na$��] I ���I���z������w�Vm2G���򉖪��7�BD8�0�^��$�=u�~u�B����v޹�Ii)0[��e%�Ur��F�{9�[������b��`���P�G[�r)R��,�-66s�V�ZB���h�XH�����bqE�+�;�ǐ%�E�I{�LI��W *�4͊9j;��'����W�.��G��0�I���������
��k���*��!�{\���D�yC/����<��`�����/�����1��-�s��36��?�Ζ�Y�<��-��a�j�nD�R	~������I� 3�m�-4TA�PB����+���n�����4�V�2��|�R ���K��nk'��d�[k�������r��ƗgD��ǲ� �	u!
ޢ=�+���Tɝ�rȿ���+]ܲ�R�AۯH^���	��:^%�/}��b.�q��I%2�fQ ��3ʨ$�os��uo��)$���� ���$���P�z���G�_Ɂ���.3]BY��G&R,��Ej�K'u��B[s�y�ڟh��p�.$;�������cV�=�MMMiFh�vq#f�2]F�E�ڌ|�s`�q.a@���D����D�w-�����*<�du�Zz~>�I�j���NEC�:-'ګ�����F�sSo�,�N� �$�q�TM �d6�d�!$�Z�����Lg�h�H	Ca��lA	�C��k�Jy����t�UƼeAҗ{�,ǋHEea6:5_䰩�h|��'�>�T�U�g����Y���o��k�QV��Q�
7����ɺ�e��~ 
8 w�F�e63�Ll����iP����2*���G��)�d{�B��߾�2�oi��p� ���S�}3b=�t�]�|�M RI$����%,�O��l�A�`���,�:O/�	ʙz�V�ݓ����̳�$����у�DY��^��T]�>Ű�a@[;��~3)���?��9�Ǐ0$�L����PC.��Zk�Җ��Ba�$�G����8�Lq�Ki����$Y�׉I+gp��� H@,�݌w���2�LG�I4fWx�d$��(���q+,n��]ύJL�c�z:jp�4�G����	$��$�N�Pp��e.��e(��+�HL@����9�
ql�C�@"@��a)2I*y7�����Cwnj����$�^T�B$����!��ZN�!;�r�wiF�{9���6��|w�$@=�I K$��,�I$�c��`ԍ��q1Ry�}>����v��O�;|�yy��w^G������k)�������xZ�����k��뜪7DՓ�� $~�Tj;.�:��� �X1�kclH!"*���I��}U}{!+���
e �R~9��9� {	�]uo�'��3�����ѷs^4H��� �I0[��U����9��^���)��UC�KsvW\�V�A�զ�jV�Qv�Rc8�s��mj����Vl�����.tE�Éa�,�<�H$�]yZR@*d�8�x�ڪ	E\��9Г��0����2@7��O�"e&�$��j8�N��1d��+���InF\<��W7�x���"�/fH�d$�v�yB�$C���t�eLtZ������7�
d�LX0����!/c����@;;kDf���'|�s]L����� J(.gK��UI
�$�C�]��0vs' �Y�.z�Ⱦ��K��:{|0@��&�GyU$@=��C�q��f�Ȳb��`�A�lA	���7��)�@I4�׉J�Of��t=?Nj@CNC�iI�%[�+�.�,gm�4��S��:Z����o���ўv;
�*��Ll5���;7=��<���	�	��z�f�,?�ׁ�� I8.	PAr��[���;�Ø��{���kX�ZѰ�v�׷׶�U.j��Iu��d8������&�%��k.\d��%r�k�1t(���4h�re��J�����k��%��ƫr6�*�%4Mq���f��	c���-!M0������f�m��p�v���eT�pL=���MIJ؋��Ĳ�.�����
�F�d@l9��Bmn�Vl�$v�U��a�]s0�7lD)�k��D��F٭��8�LV�6�0�@#�4�i�����Q	ɇ�
�	�8��;�	%���z����I Z'�6J�ت�G�Iܰ�c�$�ǿ*����<��A�<�nߪީ� ���D���WCѶ�� ��D�Iv�I�H���֣B�&3�x�}�S �q|����8�Y��z�I�	��w�kĤ���D%����ٌ|:�J`�q�UHd����$�N���HD
�z�N<��w�L�[��&�i�W�H�]���1�`���-�H)��^*��a�zE�js'g1a&���I֡Mr�jUڞ�	�x&�~�z�� �ׯRA$���dg�����������@��Z�p�H��!���[�z�
��"˯�2����~S�Ivq�������S=$L�޼O� 9ߌN#:r�Ml�F�K�L���r�+ى2�e���b�O^	�8̤�ힽ�<K˒����u�sZ���o�����ʨ�O�=���u��=<����w��5�Q}9V��Eϑ�n�)���B�l&��/��u��n�����ߎH�L�Ը��xkZ�
~�Ei��B�h )��* �H�2
�A]޽�ĕ��$�I����ǒ$
��Y����_]����4q�<��p��39�}o@P	��}��B@K���m`P����W��ݝ��f$�JYúe�[�`���$�ȼGRN�C�Œz_��r�B1��d��!�N�ą9 ���3!$3����Fh��n�2F�D���I�
0 D�;O0�BI �K�����E¿nѩ�*9	!�|->�A������x4$~g�I�싥T��r��^m�<O�E/'g�0�' ��F�q�(���^ΈP�f��׈K�Z��������Cy<�'2��I$�M�h[S�y��%���	���-:�����O���QY%���>��s��)4v������%�3��Hf�Ģ�	�%vř��H���R()g���}�1��'�WY�	 }�`�;�O��s�T�I%��ji"������sN��=WCd��������w�y��<}�_v��V���
^���咸W��n=�w7eAo/DeE��O%�����<I)����w�F�0:�N��:э&�@ZӶ�S �\m�@�I	��������iԯc�i�) ����� �m��u�
s'�]�<�����u��a 	�~2% Z��	��z��m4D$6z&ugc:WM`2^d���[S��ڎ���%�M�~^�y�J[ܶgD���:]���aL�8m�I�=�^H���zU*K=��%ޭA � Rt����:0�a�hl�n�6�b<,Դ��`v"�R�����,�@/��pn<`�D��u3�NI$;�$�!"��C*=+�9���!2��3(�X�\�)!������N�����%$��l��_�D�g>�JL��t]��X�I�<��w�� �T��|��}���or�U��3��bIu��xcAN���&�����{�`�Y R	u�Ą�$K7�[��Je��JH$=�5592Kw�I ȍ�ν&!��q ����c����K��-��,�*���I�M��$��$Qp�㏻D��o����pT?������=$�5O��]G�ą��DqNY�m�^T��	�����>�T�c'�^5q�p�Y~ٽ�o{�
�>�S��� �4Р�M*�4�+PD�DYY �6�C���߽�<�7����|�P`���"�뷙d�D�o�d�����^J�N ���T��;��1��K��Y�dqM�xr�b��(�p��Z����f�儻rll�t�4�1��6��a�M�.����>C���eֲ}�Ci��	�
����<L3��Ƞ���3!)~��kf2�\{�5��T)y�.gt�-�U�^�`�@/��ފ3(�E{+l�j����S�R�I�"ϙ�&R%�f@E$��d�~�Z)(l*�� �
�3��$0��G	��$�=ֻN<��[8]�K��L��	2����S��&ǀ���ǽ�G.�t$`Շ���[=�3��Ͳ@$�I{#��vw��[�s�j3xxG����dI��Ko[�0���q��}�2���.�~y׿q��Y �TI,�S��]���&Y$����T|����7�B�?�^g��(2˳�x�F?U��ը����r��b��~�j��5�<z�Wᔿi����%�5���ɉa��zo�����c�T��X���a����*ƚD*21��&0�@i ���Cly���/�Z95�6�+��b����@9�gSM��n��c\��kqR#����a�eƚ�u���w2����c4��\��9�av0��TfaJ�X�"�����L1��M�JFÔH�:�MP�T ��8�n����M���L洆��B5hWC�l�а��4Xd�F�"VSb��vUe$�Z��v�e��֑+����&�I�b9�Z0�5�X��`��|���Pbw̷��S:.�g��4�L����-P�Y���a�R�w�޺�3���u�`�p��Ã��KUVlI-�A�у}pڞ5��9$C�di�d$Z��z�U���;�zt�a1��,�HWJ� D��9�s�6})$Ybϊ�hE �7��x�4h������D�U�g��Խ  $�k�cФ���80!QAF.��/CFM	7�:&��L���z��Ky�@^��q���>P��eI�d�x�5���}�D� ZاU��1PD�d��P��X���/�0��Y:I��m���<�Z�{(|�J5�Ukvm�2�$��ZkG	�5�\�[-��fl6�C���c���4���($�/_�|�G�}w�D�켧��^�^}�  �{�.��R'�y.ȅ��1*v�jeS��O�@� ��R��Z}�4��7�gk��{G�zw[�g����9%p���;�`�J=_�b��32��Iu��X��0~�0��@H`k!���gZ'�Zm&2�6�2��k\ϭ�m|��y�ݵ��; W��=��k�T���p��*	�b��79e�1'�}$c$fΡ��t<�^���1o�kR ��N��� D�@���/�xbP��k��z��� �ӻdF8Fw����y�Ɠ�8H�݆|p�"�<��12d�l���{C��x�Ec�c� &�y�Y0����б����]�C�������[L�Ke��t$-��j�Is�d1�P��	uW����!���Gp0r�a���މ0P���-̖n�\,�UZ���mR��䳱�Dgv̱!g��Aq ��(��-2N���;�8��l�]��$	�.d2����s_W;����H��-�aӹPbgU\�i!��r$����A���2�~\����r^�n�n���^+l�nF�	�ޓ�r��z{���+.i����+Ͻ�agŎ|^������˧��jY���p�В1�9�_{������f!��%[�}����&��L���0ޣ�͙��n����N=��ntY��|�� 7[���Q��	�0����{�G��w������A�N��Ӹu���p@E�����J��=�0ͷQ��7���j��}�ۛ}�x����lm!�|n����a�e�Í?=��ӣݥ�{O��n��.�O��!������(-�b/n_[q>^�۳gZ�Q��?\@����^3�8n���pE�h�- |�����)�U��у.$8���_w��/�=�;��x�i假���9������@��~��������-ߎ^25x�>`�.т�(���J{��ç���I]�O-Jgq&o��I��2m�=}%�gK}��H���=���u�O��}T��m͛o���}��-�%��x�i�5�f����:W��j݃ n���s}�C���*a������Wֳo����>�t�_8L�Ք�X�ri������u�	���N�7\��>2��Eʽ���S�c��*o���'w}7��J�͆�� ZM{���Y���8�T�x*���T�a��YW��s)�� ��hH�R� ��D.��Tn&�EG _y��.��O+�:MG�e;k@��*�ٗ���H#)39������� ^�YY"Gݸyr~&�OO�&>}|~q�/ӊ�s4k�B=��o��A���\�S.QQp�I#�HB<�$HF@1�돯����q�?�z�v�����S�\�{Bv\���.W/�Q�I!$V�ׯ�����q�y�w��}ׂ��8�%L�T.O"ʹʂ'�ˑG"9TU�IN8������q�>�z�y�?_ÕgNQr�]�\� .��eGe2�+�#�6������q�<}z�Ձ �R2iU��EE��Q3�L�Q�\�\(����dW�(�UDEUTr9r��L*�(�A��*�A(�$�NI�~D��(G.(�r��ECӈE\#�\������*�$�L��"z��w��!F�p������9!�PJ���Eu�\�+.=D�bAW �)�Q�Q��G
�i��1δm�6h�8�q�Ci VEX$@�����OYQ����igvt@/���6�h�	'eQ@y��VzD�+|�z��d�;$k�a��l�b�گ�"3ݶ�����2d�<̰�pQ+g�H@���e]����
�<Mk��r^ �b#fA �����A�{�	 ���툐��P���Qq����[B��#ذ.�4&�����ca3�Zױj��C�y����� y�a4�H�{�A�0o19�)��Z�ā�i�(��ڂ|,P��<P_Ur�
%�gw`7Q0���$)�'h
ۙܐ9��	��6��^�%��ǭ{	0T���6A�@"Ǽ�r A�y�or��t�5����)�#y�H�	��aB*@�U����rՠ�@��D�I�b�@)���v�Mm)9F:�1��n�;�I�L9�H���zz���+�htX;|����\V��n��jw[a���Ͷ��UO�c�7=����2��ǐ��}A��?���s�����Zp���0��ZL��S)���&S`]�v�D� �R��P�>��t�d��	'eQQ�Ҷ�� ����Z�^��PpO<JlX�Fl�d�{�ڤ�Ap<ЛOl�>ea���[�I݅?m���<��(�xrs��mVR)Lk�4�k؍[���e�.����8�J	��K��r$�@>�]#�C��dK]���Y)]�`�{%����[�Ԃ@��J��C�x�q���'ٿLt�	 �2\˒�R@�L���$	�؞zbl�d;H�,A'
;������h&\��<�0 ^vULoVh'3n�rĊ�ɐ@0�<��r��\x�a��z�$�6\�L�v&A ��M:��-ך8�/j��
V<�'Pbl�E�%�$f�d	�Yy���Z�5Cǔ�@9ד$���2}�c�G/1������FCʗ��2�5���%�$Հ^<���9m�d��� �>�S/�q���'{{AΚ`��5|s�p.�љ��m$=�[��U}B��O~=�z�������Y�U����7�F4�:֝�Qֱ�֍�`P�(e��\�7zG�޺~yxx�X��w��k�O5�d��XX%[�.sNĸ�բ��S[pCe2��5��A��e3.��pö�*d��eؘ"L�lY�\�K
ŗ��%��SMt
�	c��Zb�]B���Z�Y���`c+��=a�Ȍ�a3�3]L�(��H]���c�&��Q���d�1�v�*�p��֪i\�"AXV��M4�mt)70v4m%���u��)�6�SM��ʋg�����R���EG�߅�Q�X����� �̘ ��^e�5�vM�los���r9�S� ��\0:�&�1a�rs��{5�7:L��o�nC�H�ܾ�(&H���a$���Ft=�����%������X���Fh65��i�y�K&H3��A �w��m.W0��A���Aa�= H��|,�!�DxS�Vx�Dz�� ���I�H�G��d@#9��8^��j3Kc�-g��@KD4m[��Ax$������	 ���}�nn��w���y�m�n̐2u�$@�U�N�¸�͝˟2H$���ѕ"��.Ɋ�R�M�ِ��C9e�v�2�8���}Ͽ���>��S�����L��[N��d�%�"׮R�f��:����XKA]�L������J+���Ra�`�$U���N�,�Z��������������?�x��Z�>��������=A�;=�3 ���ϱ�O�|/W���{�xP�#�P����<{�\.�����v�o����"�L;���e0�[`S��@ε��aq���`�yw��q�>4�מ��$�ןTI��̶�~��ы��P��x&=@�-�z �d��(�$��"_����Q&;�9����Hl�\��l�������y��f ExZ�pzN��ys�Z��惈J����߭�s��c'=
�p�\=<Qe�M��{�<w�M����U)���S�{���"�~�����v��I��CK�&ꁱ��G��]!�{ݱ$�86���X/�s,��<���:@��:��Jǣ�L_L��'�#�qj�K��ֱ�b�U��P6oS6;L��h.����$1��G�dFyM�xd�Nvt�i��Y���)^��羐I�@K,6z����Nb�uw��������n<��o;L�e��� �l�H$��\>)���ö���@���tQvO%GimK���}a�E��&#o?��f�ݹP?��Ԟ����F\ٳ����g=ۍ&;}�)��[t�%O�p������s�ɥ�^|�P��ߎ3��4�u�c.u�b]hi�2�/ϧIbw�~@H%��g� �D��V���"�Lxy�g��.�&N��A)_K9`I��%�bã��L�
���cs�F�F�$�$����	(�woX�t��d�6��23�G�u^F��]1^R@$�v��$�G_�F�l�^�|���в��B߇Q����L��8� ܬ�����ѳ:��Oc� ��n��t�C�������E��� � ���j�)	�!�F֩OB���� kdt� �rA��|��O����#�1���T���l��"Kb�}�2��)=����p;����, Tt*C!р��
���� �E܈iL@%�*�x�"��؈���L@C�"A ���i95c]]��IEQ�]{ă����&�ZB'ՙ KA$���T<�w)�߫�����ڼ��z����r�7/d��9^iW7��-�w�8w�CI[�v������}���vﺹL�]R;��b���ǊY�����x�l���N։�u��րӲ�˰�ce�3ڀL���'�/���ú�^	��>v�$�b��=K��2]9�#s�sQ�`z��%�g�� �� ��av��W��R�g��%ܞ\�yO,j.&3�H7F�m������J��kK�I֘�:'�sK&��I� M�� $hyw������Ѻ=�9@P0ɔ�8z�\-�#�9��"��/��\��C{&z7�S�&�=q�M2`�_�4���@;7��l��*�_�~�y]�IO�LWmL4��~�,q�)���צlo��꽃 ��܉��� �x�F�ã9�+���ɯ4�xz c!��2	>��y��$���;InPqt=,@Ly�dMt{�(�C�IE������d_@�b�6��7"���m�'�uP'��@P.�v�OX�ٺ�8�O��˧��q�z��f�e\]�	َ�;��xy+������[�N*zծ��uo�7��,{�l���~G�{=`@��k�_�4f�]~|�H�f���0��;�@��~���k@i���D��le�� wH;�	M�z�[/](Ʀ"ᔺ����r�aM6
Ifɨ��`������\35��l���u3d�՛��.��.�pc`9��^a����4M���]4a5��+0��3-D���#�Mv�4`GK��Ԙ3)�0�C9�T�sNw6�Ur�i+p$W,ch��nK��#p�rE���Z�hͭٸ�ଵ�4��d�6oҁR�1�i�jn5��ip�9�a��P�=����r���c��߫d	�k�oTAj޾y���]}
�����o��}��/�4������A�}�q��&.ϧ�n�9��]�!���$�2A��t�HDb�++S�a!�f̘io*��ɇ1���!+�}� &H�#�o/_ޢ�^���EvG��A-�ޙV�A\�`����J.��Q���<���	 ϩ�!S%�������Pi$��7W> ��|�m�:��
�Ω� �`�Yu�P�YOTm�d����$��7�Iiw�2Ӟq������~6��U�%(�2�3Q7ea��p8� �]Xe��׊�[�Kf`T��m/�����Iv�0�n�UKܲ$o����[I��'_^�'�'k�>�Y�:���'�˅����<+�o�j�S����V���QQAC���#�/և��T3���,���~J��J�{��n�?"���h�^˰=�/�#�Zٷ�ƛ�7�3�w�F�� -�ε�-h1!��
a"�~{�ϑ ����얐�~�޹� x�i'�{5]>����#���w����""G5�eL�0��L�,KE�n�[t�a�%�k��Ơ�'��[)57��axL9��[ �����K���Fv�$4�f, D�H��b;y�q�=���[lHzܑ"�yf�D!�${���-${�v\���]�X)����VcĝdȞ|��N��K�a����
�7�A>��`�h�k1X*�Y�%�rdi�6��L �^ՙ����2�u�'�z}�"A'=~�&�G9����^5W��>j���2[,�zoYi%�@*.��S���h����s�{��2B[��!�ޙ%���)bMUoh~��KXD>q�.�#��X�N�� ������Y�+�y.�#`��6��vA���_{r�jգ����j�v{C��<nm�u��K��g���͵{�v��ׯy��G^����|T���`�ֶŭl��ZM�\�(��@��#�37��%7�G�T	Ru��x%ôG��랙C�we���4P�5 ;$	�9��C�,V_t����O=��G�|Uoy�f��!7M@J�1���\�A�K{`�H|��^>/�4{���X���jI ��D����Z�گ@D
$a���At�� �l4��fk*Κ���ke�2e��va~���on��x �Ts���2Gγ�䃾ސ�ۈʽ3��6䡜�܉�܏<�K�[�l�Δ(�Hּo�N��xǻJ�s�6ɥ���	�����ɖ$ۊ��M=��eD�L@*$V�R�,�$��_D�$�W3�E����O{d�5�;�e�-�}"D3֝��(
�1����uޱYt�y-H�����E��Ίb^����'>��]�/?������({����*ȫ�bG!���,N\{(���N>�|H�{����w���XM]�������������F-k�:֓��6SePD����~}}v)zN���p]�*��t�&��}�鄷ٓs+y���y�LGb�$���`A�M,��ӗX���A��{TS�%@|-!��-XZ�"Rdsvسs���(�Pn�O=Yo�wܰ��P�#�V?b��I<���I��1����qk&�bX�i���pAa0�A��~����<%��������Y��t�"Wo9𨉧�3�=�O���'P�Mcs{��,H=u�$b��Ep�O�MX����8�d�bA'}]E[-%� bQ"�.�3�����A'g�2I;�Ԝ	��Di��I۽]T)��$��娹P�bŀo}Q �>�!ˌ�LC��&.D�D|�KKc'��)<
ff�;�1{9�n$�T�B3�׻�����>��sh���K�r��>��>x�<\Ӏf��h���A�W�ރ�;���^����s��z{go�nB��>�"��{]�sM�i����.�b�����qɳ=�y�2��]�t�?2�����������P���c���u\91�U�ƵӼ�;r�V�{�x�Y��l���J���nY�V5b}%�)�{#�y���g�]�%�l�����w�sֽ;��a8u�&�k���䷘��. �B��C�$�-�����O �Y�{}�������~���D9R鞉l��ûS�PMs���;<_g��-3��.�U�ң�ͳ���G��f����7��T��/�w�ٸ������2�(7y�z�Ц�� ��J��ǔ:x��'v�������>�#D=�rgn�l�ݞ�+l-%��Xq����d�z��O7�]��7�7X��^�?g�i\��?M�#q���|��GY�<�{��s���Jo���'�b�+�B��Sw����n[��5�m�~���x��٫��Y��{ݡ�[��![J�L�+��'�����ǻ�9AV/d����%n}�����w-\���g�\��G�����)�W�~w��'C�޾|yg</|��n��٣�=��^;{���z%}��Ӑ�������=�d���1�l,F�@�ށ�}a����m�Rs�x�1�*4\>g�㛐��~o'��k ��kPp�3��c�F@�ds���/Tc	�⴬gQb�:��rG~�(g�N�e��p�@b\ ��D,}��xN� �1�pr���#Ah�O�<G�rz��ɸJ[�z��P'��_��2j�	�܀0ӄ�H0���y�=����W.]�+��L��n%r��8}R���
x�����<z�8�׏ǯ]y�U��L��(��/���ߎ?G�(���t�)$$�����q�q�q��ׯ]x.z�G��0;x���U\��t�PA�Uȇ���ׯ��8�^>�z�[@� �r��DQEaׯ^���1�8�=x���e�H���(.W9L֔E�e��ȉ��;j�S(�*��.TE>��EPQr���\�\(�QfE�p���EȈ�*9TQ=R"������H�gg�
"�+�����(���9G'R(���L���U�(��EAUȋ�ª���<l�~��Wم�l�c<��H�����%�+��65k���i3�q(8C��l��9�l��iL���h���:��l��2�ۛF\�ms�k2�t�*����Q�Ʋ�+ i�t��M��X٫p2�J!���k��0�DĮ,�ՠ��e����͵SB,���ۈf�crᵄ�d] �M�6`�f����H�^"�r�m �k��))�7/m��5�o$`�T�����T`�6�
��1V5�*�l�ԷEZ�]f֐�&bښX�۳�"b�O�C_'�i/fCe��݋�da��$�͸̺�)y�g$ٱ��������m7\�[
o'���ư��]�`�d�k�d:jL�hh�@&:�r�p�D�^ֱ�8��J�*�VX�����롔�����1X1cPu�F��h۬�6�[-z��DlSU�V��R<4��`�DV�h�Z�]�8#�KasBb���-�᮵�尚�f�j1 F���#�F��m�֒��E���4Cf�m0��,���֔����7\�434�g\��(�l
͙�܈�q�k�E�R�Z�L6,�tv�A��F�nH�uD����JSb%��'�J¼��S-!d��B:يi2V2�I�2��m3FуKaPr�L�t�(1Ú��nb�c[�A�6wU%��M�,]af�gh�;���X�aэ�m�a�2!�&n�x��ɣ���	�-81^6�4mR�s�KI�f�󚎹��j	�ZV�k�q0�A��\ZBb�L�#R��F�s�M�-����ғ2�qp�"��*�tvV�a5kZVdb3e���խ����tE�Y�x��[,e��E(����Ӟ�y��9��"O[Ɉ�k|P͔��D�@��p���UYs�\���\ɋ�=e�c3�5��Q�$Ƈ�k�y��.��'��lK�m .ε���쉗 ������t=��f�0;՛cBPJ�F4��!BQŨG�x%��,�5bD6�м��qf���.�����2�	��\��up��й뉇q�Vh[2ݹ��Fep��+KA�66��ThBiP��a��l����	H3n���`��C&cX�ˬه	V���Kwnv][���؍�ZM�*i��#dA���7�'�."�ce�Þ�k%��2Ų�
٦�s
�f�,�;���=��ܘrDG����&A`A���I�;_�I��u��e.9�7,M�O<x,A�*�U{���(�E���[�K쐩��%�g?E=gv��ޞ�N#c��᪻a�*�%Ǽ9�:��i�(��R@@b����)��S�r,I���	LS&Hr%�Q���8P���Ω�|��Vk���[3ޖfS$S!�ͩ�H���ѳG��������R�K.%� bQTx���M��%�-4/x�ue>S':��1�}�=��,m��ls��J��%�Y���ef�a�-�X�3f�UEn�r$�WYlK���Ҵ��Ŀ9��i �2�̴H'o�d�H_(�r��.�S�$�k˥Jb�mߊ�N�(����ɐM�#����U���~�m �}���g��
�&uZ-d�My�;D�v�;l�g���~�^A��Y~��w-���.q�h5wfN'�˽��ޏ��;��h�:ыZ���o��~�������BA=}-#�ѫ�Գ�s2[�>���9 �s"�c�	�� �m�zwkG�m� ���2Ē�s�o'n�W�^@%����Oi��ר'�֬���%�]��L��ʭZ=�>/Y/eF�$;W�o�?����E��St�{=�r9_@�tw���"��D�@���L�d��BȒG��Y��s%�5��ab�R+K�%�VX:�Jݑ ��*��D'%�$���C��@����w���$��ĒA9N�{�L��p�N�W�2	;ݑ,Ks?_E�9P	�R��В������^���<�8v�id�l�@;Փ)��XÒZH���D��Y��� �Cb�d�	c���F��z�R1��!z�j��Ѻ��	m�c�ܰI;����~�nh(��:�O�����}�Ѥ�r��u��c�L8pj��RK��K�2`�d�#�bZ��G(��"��?|��Z��&Y 	vK���H�:Ic��+C�b
�10�J�Eܯb=a�kLH>޸�M��2D�3OE;)����Z��Ċh�S,j%u�8r�b.���MH�	���	��:$x�CϺBiD�����lP�ފ ��f\����i�ũ/�B@6A��I�K��e�Sh�5m�ʴub
	���|�;��q�'n�X�̭�s�2A ��G���A鞑�iM�˶�	��+��In��!��D�z����^s�!LNtKiNO��2,����<��+g|��Ǔ�/��˘ޤ�4nq�\�uA1���y�L�@&��� L�w�{������>��G>w��	�:d�f�x��+:���QB�Et��Y���8c*S��u"@�שD�H��9�>�@Ȁ�A�UJ�w��L�^s���<��-/]]�(�n�~F������yGӬ<�cњW^���3Z���9�Z�S�0#0^ڈ��$��7�K�x
K�/����%`wtI�3Y�K(S�n��D� �r���7y@�� �D'�^"l]����a%��)]�:in"���*ۡ��L��%�@H�?L�v�Ç." ������;��(��L����L	��ιПl�0>]ԃּУz<e���ZϠ��xP�z��ޙ%��7\��*t�Þȭd�Ec P�[�:d=E�qǑ���Aj����(�Tg�)���o��A �L�UԬBҾ���1�p,K{:'i��tA�h��|�u@1���$d���z�|'�q��fj\Έ}��<�"�˴�b�Ϙ��^z�G�?��%��A,T_��0�x(�wީ� �"=� O��5�_�6�����x$��$��L��ӱ�	�����HGZɲN�#VU/$ڠEnx\�z{zȫ���p~�k�}���R��@Ft���ʻ��ۛ�/Wk�;�n1�ψ��2�7��I�]J�x�<yi��N�q���G��Q�m�[�B�AK1m.���l{K�4Cc�[��E�3`�	�2��!K���	R�Ij�1�n4�p;9�Ҙ�
��#Y4��B�D�E&��`P6�ڗ�f���L�[e�tv�v�0�ܙ&*˩�v��Ku.a����9�֎V.�ڪ)h�����.�<�H�1pZ�L��0n%�4;�4���`Q-70�6)EU�gV-L&�-�%����)�my�|�>I@�,!=����f�n�~���|�ȀS ���I,Lo�d1���j/v�z�	b@ͽ�k�*��`�." ���lu=��H�V�5���Q���� H1��$�^�I��8l^�g���%�29�wN�8���H&;�H$a��s�<c�Bȕ,S�}H$��ED"�WWd-&!ȇ�Tf�:�aY|������	����-i��8���=�>��f�@��zfX�>n��P<z��$�d���]*�e)v^,KV�L�K�W"I�oz$��*]�D�o�},�"�N��XG��*GF�K�3]�X�-�]�ܓ\T��Mܫ%��Pt���_�c��W��}�	��qx�M"
gG��$�Nz|���{"@�JY _c�����{Jֲ%�xO"�1�즒
�'��4����C�g�_�S�m�����'���=�-�[��Zy������M�{;���dמ'��Z�N}t|��� ,X�Ǟ�<Q ���j���!o\��H��$�I;��cf,K��C�	B��P%�2V˳r��Ko�69OX�I5y�H ��D�d���U��.��'zȁ}s���9�S�ְ1�+e�؉$s���IbF{�q˛zs����˪�w?���%]\��A�?�$��d�E��?��3Y`z�bA,H5�I=��	�Ui���(� �r���첋3���7f���1&1�J��r!��݇-�u��|N�×�Lp�vke��9�7ޖ�2��"Sd��vT�K��bd�$	 ߺ`N�{�gwD��=�:&�X��j�$�s��AL��<A�׽2D)�Q}�C.c�)��R�E�	��F>�H$glILQ��.M�c]8z��R]��NԻ8`[݅���6�=���������:_���K�Ѯ�x�ذm�:2k݆�^�����{8}��#��F1���3W��j���G�Q���~5P��Y9q�$y��S��P���-� Jd�vL�H;���^�x��1�g[���d��>�Hd	��:q\��	�c:�ܐ$�����޻���MD7�Q>ܙ�L�	&��Ꙉңѱ2OԆRƣJ߳U�u����0̭��#v�-Θ�1�8ؚ0�0"qCO��ϵ���a�~�����ă���26�ܐ��=/���"n����z�6�7��j���^�N�����D^��4�_V���\�)WCƽ��,I V�$��a��(�t��(&�z�}�{:<�Cz�΄���/��mH�A7�p�a�����9mP��F�\[M y��,[}ޙ"�U,d�A/^���f<up]a�~�LI0��!�c{��Q[ފ[u��gxǽA���yx�q��ɍ�dF`3�y_n��h־Ox��b~�}���&\>}���ky��jy�;�r�EQ����z��1��|�I�El� ��j�!ˈ��TVuL�O!垐&_[��:��������s��Ac��j�4���~Vbx.��JZK��i���k���A䉦hf�u�e�2��<��X0Y�Q
F{�!'w���s?��,i��,ZS�=�qLtLow���G6@���?��^���Tп�e�[�]Y"x�
����zdL2]�3,}��L_�"AbO�=*�������'ﴜaҁK�x��I &C����^d^�ƻ�W�}����t(�tH:�~+z��P���6����;����t_�R�,� �]]�����;����o���2r��ݝgtaʈ/m�o$����g�=��Di�����������E7葌���|��>�i�w*C(з�y꪿q�Y�,��.A0�L�����wI͖U>�݂nE�ks_�^=�1����jSׇ��w��	�T��F�;��� � Bp���p	���L��5�4���U(��`F1�}��r~T��69f�#f�3��UmL��	]�k��R:(.��j�UCK��X�Nm���{l=E��Dv�*�Z�:��sL��@D�D�-n5�S0��t�����@y��Xc��lL�1��5��(�C՚\&��fF��3��]m[�Q��[6�%&�� �jU�����`ь��  q6���(���]�[Ky+�[�^��j�s6	c&�\�o�����&4T!��ʁ,EFd��I�����s��r!��Ϻ$�h��C�N�	ӏy���$�E��^�u��a�n��Z� ��$��ޙ=���k|)n���ϩ�lj~�U���b��G�!	���l���y��O���d��� $�:7cX�������t<'*A/z��znW	��s�d�/+dIbI���[���,�F�&ߵ���I+h��N��
.�U�=2�X�w]L�ӛ�<���}m�A���5"|ɩ��(Q �_�o����S�OQ��j��f�PGgJD�4��X&V��L���ӯ ��D�z���<'�~�\�OH�E�>�ؐK���� ��{��7�Ҁ$糤	`g��}�`�" ���_mD׉ �^�!��^���������BL_�����U��~+c���I��ڳ�Eu>׾d�k�}�R>]^r�x^����^1��O�,��X,X�b�e�&�@�DL�������L��$��1�뢡z�z���uh�.�qT�T� S$z��$�@$�Nn����@ �.��X�vD�N��D��y9\��q	�M�ީ%ɻ��S���&R�H�w�&p���}#�>�����1B��"V�pa�x�
c�Y�7E�K�җ��r�O`��f:$�a�퍖	��"ZY��P�"�f(�0��H��I<v�<QsD�L�u���0$#��e��ؔ��jir�:������� ��N��BN�#��m�"��]A'_�<�Q���w���t����u�y2w|@�w�Y�w��GTdI��(�l5;�s,@$�~�L�]"���ף#C��gd��1�Y�q �<G`�I�%�$&�	�M���	y��L����}��j-��]4D��F�7�#����b'�z{�rY��tN;�k�6vΑ�]	��V��<vx+���f^ۏ���Un�R?Oaf��<�}gOj��<�^@ |z����W����hW:��S�5���FZ0\�����^��hzw��������'-���WG��]�h�';̓ꏆ���g�<�K7{�N�o��.��ϳ��.��a�O��r�y�{ܚ��e�ۮ3��{�F���<#�w�ΙÓ��xX��������������O.н��2Q+���x��V��S�9�u�ɯ�Wנ��=����ٝ�闉u.!g��OC5r	z%�9���v�������`��	�Ywӵ��+�����)g����7毽���%�ی(������cޙ{��"��ߒ���ż��A�=�Z3b�
��@��-�V}������]���4!_M��zO]ů]��7�n6D?y�r�YnH=u[�	� �+ w}����J��ҋ+y�>x|'^�پ�|N�t��v���������C�e�@��8�>W���o��6�m#4��G�^��=NoO
��f�N7/{'x=z��X6gv�{���\���6���G�$�nn���W۾���w{;,S� �]wz;P��:���P��>9��Y�����8����,��Ύ+�˱.�`�>f}>(�	�{w�l�|/}ҽ���x�� �'��*x���-.a4y�QD+AI�sm����p�N�빱���?>���hwB��vS:x�
�t�+N�$)�Ts���AU�L.ф�$�0�$	#�q�o^<c���qǯ>�n�	#H�U�+��"��"�~�o�5B2C���^<|x��8�^�}z�ð*$�HBr	A(��RA��ީ$*�	N>8���ƞ��8���׭��i�d���`Ip�H$���#-����׏}q�q�׏�]6��"e�H~mH�"�U:ҹWT���h��n{#��Q2���A�2
�eL�9p��L�P�M!f�������PS����3�dQS#�y��y��C.�"Ѭ��d�̙VI��
�"�]!:AADDL��K6V�8'*��(.\�	$�N1#1��e���ϝ�Ļ	8��,H���O��"�w7a��}�}���zI}�,�I�J:�I$w��0{˳��c9��2Ӳ�uH���m\���O�b�u`�Gz�1� /ۜ�#�;hY�j}w[�����$��yb@%�}�%�8=u�l�(�D8w��;�\���u4�&�P��T&D%0m^�.�z���ߛ�a�ȟsI�3��I"��3l�}c{hv�!��>��M�SEjJ�f��*��'x��5�@�+ELn���&�9� �^Y��5�$�o����-�	4ۆ�x9q	����L��zP!gl	b����i���Ih�]�,K�ޙ*:F�$�@A	�b��{�O�r�&M�K�C8�����5��A-+���}��.�{�L��t��-�-��� ����f?l3j����wy~����Ծ���𤯇�qiq�_f�h���3p }������Y�(:�c�g�Bќi��y ��$��䟁xE<$�}o�Q �L�����cڏ�����H'z�H�N��P����C�x&�H�/�4�Db��kF����ۓDf[cF��]HM۰�٬,W�o������O#���p�I�̉ �$oo�H1>6���1Yl[<_��H�wH=�O���"�!�K�I�N��j<5Ё�/2�H%��IbA��KH,W\/np���K)���pT�*�gfD2���=�2y�5�@^)���E��q��$|��L���Ͳ�r��#Ϛpe9Bx��T8���y0��_��g�$��C;�훷4�^O�믪���R��N4��H9*!�]�}�L�E�=���B��']Q�Sњ�\4�^�e��s��Z�T#o���x���
QğW4��P��M�f�Ƿ�@�1���x�mp�F���^� ���;��c1��W:��d}V=%�Ac9$��Ӿq�q�O�}B�qsuٸ�kr�&���-��H�U�4L�Be���c�0��!��Ip/Y�$).\c1��.�%�B�X)\�d��Jr�&�n�3%ִM�[Ŕ���(�jM���������ґ��°q�#+3/g�c�<,a`n�-p�jhkTf�V�b,+B���mm4@��XX2�+��y��m�Eef�BmnL���ݥ�m��kTt�R��0�}ݾK�\ݵ��?9<�� ��d�A-�;�x�D	W��@g_�8�A ��&�=H>� �$Bz���� ���c��Y�ѥ�F���z�c���<�H���fg�cZ=>�f�@y��I�C�;����e{hI$�;L�ă��dO��,�5�s �xy�<P[��)<U��L���{�Y�H̩I�Ȍ2#��*2+ȧ�ƫ��\���-)������Bx��R.��<�&� �c�K�#�\V映����ۭT^Ta�d����M�.��T�":H�sɈ�*�Ѥ�=J\�q�
�J�℞^c�y��>0\# �����$��B��>TH��tAw�l� �W�2	�<�m�;e��o{$I�FH"2�:ОO	��6cS�uH&Ym{8�;�Z�`�nz��}=�.R/G��`��<^ԩ�.C���
6��mK���)@ʅel[�d��5yNI"(�n�E{
1 � �b��q�i�!��b$�k���Z�eMk���9�u�4jQX9Gq�D�O�5(��@,e��nD�$���'1�5W<;u�� ���+�5�����LH֛�%�^ �x�Ms�a^�ȸ./�	&mG��3�W�CA`P`i�"�t�Y$��=+�-�y堗hW��#k���E��m���!��D�i������8'�弶*b�ݓ���s5�]nRƅ�b�f�o΄��ʂ�WK�+�1ep�B۬L��H��Q<���PnL{�p�r���}�G}2 �3��fč(�I�铷J�|'*�n��w/&�2�Ɂ1�7a 䨄
EwL� ���Ή��=0X�3�}̙`a�'z�db��.C�N/E�C�&�6�?9O'�ww���VL�H%�fz)�Ɓ�w�x��l�J�
^#�n9����A�,�ݘMk�mI�C'w�B������~-�Ѽ���f���0�=^���-.[��&LX�b�9��~%{z$A���|I�A��A"��2s7st�^X�I���	�$����e�OTF�8�f"}++}]�]�A����@��iu�.�(��=/[%��ó2"(ǲ�R��I>!�#�=2����=�T�1M��O=���܍�ae��pW�g��NI.�ڦ�ɡpk�5��]D�h-���:mϿ�~|�����7v�ze��e�ԒA4�y��J:/-�7���������s|�
i�UL��K�R���O�$:�l፭�bX�w����"u�� �o_��ʷ묓A��fBA�Q	�X��,H4n�Z  d���"o�����Y$�s��ج���@/˧�^A'���J�g��u*a֛���H/���S��H+�Gt�}��c��z�[��oۛ���i�,���nj[��W��I��<|_���P��IÑ�}�t֜����ӫܟ|R�wEלtΛS)���,X�b ��b�j��<B��!�=Qs�����c9�8�z#Ė静bX��>� �J�t�Rq{lk��0|nS�@tjm\��+��dñ1a���M�KYb��ileuTJ��筷K�"T('��l� �X���p�P�oL�͂1Md�U�|�z�dJb��_9K4M�
H��ǽ��2H2�Ԇ]��덙)��#J�kPDXvGL�+XGR����I6m��ё^t�$���t��V�$�6$IUu���]�����)�,~����݂��O�SD�4� y��e�ƿHE�"��2I��[��bG��Aw��$���{r�Q������R��ə�=.^��f�|:�c:q���z�g�.\j�1���	���[���մ�_EH9�5�&��ʷ	��ž�T��x�������:w�L�Q���p�g�Ǹ�b�/���d�O2�/)_gGu�IDJ4Bt���y�k,X1bo��H���+��:�jAf)�l�M�W,M6*J�1`;:\`��M��-�LK�n�D�ջ4e���"i�4��Bk��i�Ք�8��c��U�c���ikն�a���6�j���Q�� �^�cڷ�m�ni@Z]b�]�6�����e�B,vJ�v�X��X �[`V��!4�� _1�|0�W͍�K���	���#��=R�s4Is)P������C�JП�/}�I�vp=S��Ɖ7�fBe�5ˬQ�_zjZX~�&�bU�q�
E�@7��fI��C.�Q~��4k$O�;_GMl=� ����-��*h[�7wբ�!�����hK�x��L�	7��IWU��螘���O�Ǚ�/��� ,b�.W2$����HB����#�=�ˈ���[���x!�"@�V+b$0$Į���GozD�����+Ȗ�|����Mu�	9��+����
�(~��T��ə�M�\�HN�w���w{�$�3z2qp� ��}|b�}#������6��t��k3"\�W9f�5��N5j5o�����s
��|��>߀b6��H�0ϽuBM3����(���� &�ܪ$X�U��-��d>�D�	��/=�,Khc^�ʃS14����:���&�U%�Y8K��
Iy4��9o�;�{L�}���b���3������B��̀,X�bŉ6��p���z⚵��N�\����2G!�1��h�k�_��9*�ʰ��$r��<���u�$��^C �z2n��o\����$�� ��'�*}�~�3�����z|�On䴓�웘>�y�mՇ+�铃�F�Ѕ
����H$�΁4�/ղ)9
����Bc'/�I$w��@=����4��*	O�QtRO��;�c�"����+]k�n�Ý^ui[�^��U����~���%w1[��1�s�� �G_t�K���� ��L�b��fIĢ}J��O ����x|��<��{2�_\T��H�̏H�@,N_t�%����t��=��D���"T!8NE�X���$�5{^�I�##��ϑ���e�&��Qd�O������{l��}?�n�J_�H���d�7���LW�z���Qclbbb�&@���ď�}"I=}������ss��-�{o��>�6H���H${s���#���؅%d�b�yIl�K4��<b*���X�$�t�a��ˣ�)5�Cם4ƘE;���$��]"Lr�%�:d�w=I�4L�@ٺ!i���V]\+4heH7v/0��Q�U/��<���P��_��p.ɵ�w����}��/S��vz�r�5��'�=#tBA�K�:��D�q��ק�^�A�ڨ,q��d[�6i��igs@3�睤H&j��P�·�HB״S�* (G'��d�S.Uq �_Uz�\����֞Iwl� �ޮ�#�=n��(�r*�N����@M��,z��I%���%�v�@��]xf�k��0���W�����g���������mǒ�>K}
Y�y��m�I�52��\J��ݛ���r��$�e��^mN�b�ŋ,X�"����k�Վ���38�ˢ=2I=��z���9L�S�M��%�e\�7��$�iM\*����bNS���P�>���f���R*u��K�:�0!�D�ڂ-�B!� P�s�%:���YS$�o�e��NozD��^����ؙN���b�tĉl���JB�
E�]�$�ꗸ���~	��n7�I�ˇb$Cn��52�z=�J��[��]��v�Kc���_�� �������El��J��I99��IbFoT�(�\�
x����i���:�^��LF̳I���OFeט�	Ͻ'���J|o �F{�}7�l�b�a<��T�H��{bCS-�Z����&vjd뺁$�	_tH�V��g��/a�Lx�T�6��闚��H��8�����_}D��zf��y��{�u�W�����>ګ�o�������j�v���u��Og<0n��ׅ�����⯱��9n7����X�i���uZ���v��ʐ��w��˸��2QN���$�^(l���w`]��#pZlZ����ŉ����pO�_nL��E��X�{�}��Ӈ��ys4vlYӛ�AOǻH�/P�s<�A<��o�c�D�q�{;���r�����c���g�x�d�I����}y�/;3���{^U�}�7�5�����t��A����|f���݅vG����?P�Ѿ��Ǿ<=�w���pZ�}`7�綃���og�F�T�,�<9k��X�4V)n��_�c�4�ns�ږ�;;���~�~{��������3��fOYh�:�g��yPvl��pG��kPܽ�7&���n���밪�;�z�61�dҰ���Khe����0���<��<�׊�süڏ7��x�P�h��3O��I��՚}�}[���ZOg\QQƥʋ.��e�s����tx��VA��s����^��%�������|Й{�����kk��۞7���Q�Ǯ��u��=ܺ��ſz���u������%��H�}op6#w��m�T��\7r�3 ���mw!��/�l'�נ"�s!#
/\}ӧn�W�^�x;	An�߃=�=��LG����:r^*"���:$>Pvӗ=�O���=�1�P�����s&-^�?�����
�
���@�{��������,I�B)@���j	�&�7�f�D�u�"W�NX�������DQ�| �b7�ax,0���Vn��4�Df��'���������z�6��ǎH��mfM$��d܈�c��*�QȢ*9TG*�Y*�U�`DAD$"m��><i�q��x�z�x����t4C��Nx��W*���HT��[�()%x�����ǏZ}}q�z��Ƶ#�}�XUFd�	��H���(�#��E�˗.'�La��\v��ׯ^��}q�z���]�Y��Y�J��˞	��YT3��TU�����*��U=q�>�x����8�ׯ��K�<Z��9epKUN��9E9E3M&���%�!<���S�5ӮB@Rr��z���4:�h���n����*h���6�W
��pw̪����F��2k��a�!"�C��T�NP	*��Òv�dz9ޟȢR��P;F\*��Ib�[�E�i	�������"��|y��p(s�S뮖t J���(Ix���0�[�[�X�G`�v���ִ ��n-��fd �XG)n��U.1��-#�M�:�;n�6����YhFk����[X�m�X�[b������z�n�
3n-�#������R��MK��L6b3bWL�V�e�k45�a�Rز�\۩@Ms]f[�s�t���G͉��hH2�AE��fn#�,�!j�Y��tv�մf#��[�c3�f�J�qs+�I�nR��2��䁁���:�nk�T�S7��v�lE3L$�KM��l��c�Bm�����؉�7���+���u�cT�R�"�v�*]�4�n�hgd�YCK���g�k�SM�3���B�ܴ��i��6j:�k��z�n!�c���ZT��7-�e�Qv�p;��v�lE��u�YZ�H�ܴ(�135P֛lM,ܱ%�r[,ͥi�ge5�#3nAQb���J!�5�C\�F�۲��mb�`5�k�f�a�2�jˬ�`�%��X�L1���,k��#�2�&chi��0�قm,\�h�JI��h
��3����H�q�{S#�E�*a���0�mŢݣV������E��n�43�����1v��%�Y�5�t�t*]��Yeve�8��mQs��[f� fJG6gK��v%�B�[4�6�nC%en��S���:\J�hG��CZYlB�q�F;�q�B�B�4[u]f�yM�KaycR��l\E2氷� �c
���F6�������u�3x��ؾ6�.��m°�Q�:��P���ۜR��V�F9�2�yɴ�6+
l+v6��w`�\G:��4.�+�N�A+-�6��e`�gfm�t�.r&�c!� h�������]�L0&�SaF�#�M4ê;Zk@�V�m�!Y�����#4��׿��8�M�yo�CU��]�d�l
i��-��eo#.1X9�ݨ] ��������\�
������p�Rl�RXK�h�:�#uu[�1M)���b��3M����끉e�הg���5�p9;Q�q2L�Ek�W�ĺ�	�%�4#�׌��cX7Y�MƉâA6vu�XiJ�v�3BSn� ��JZN�+u��X�).��G(��c������*58�F ��_8x:&DLD��T~�.ٸ�$v��%���/E�E�ZZپ��Gp�S�����=ޒ�N8�Xv']�,���ޡ �d���@,Kw�����X����B�u���`��^�ZM�i���z'�(]�E1�ty�a��F �g�<2��ys �4ɑ랙$GF�P��.��V�s�{�kg�g#��� ��?�`sb��o�^�	�@�[2m�O
O�)�� >?g��ٷ�	�z����7�1���I,j}�0�s����͓��~82vU��I�ĒIeiK������5fW��B^܍������C���:&�S	����D�H$��H2e����J�Y��0sx�^o�ӳ�b��dNO�W�ծ2���"�ՂC��Oq����}*�!MoC��b�V����+Y:��9}��h�칣�@�j����Z�s���%�O�Z��,X�bŋ~���;8D�����$���� �}}��J�rD��u�D��&��$��LEWWT�#�?KIbX�>�����| ��y2	$���M�X��!9�
���	�ů6����:9�%=�$'��� SwdQ��WG�x� J�ý[2	�#$"�=QQ�"H�!��#}9�z��ut�`X��H��os���fvJ��Bg:�B��o�X�:�D�V�m����6��q���)�Dt����aՇ\����WY.����s,GwD��\/�������Y$�2�ބފ�n�]èI���h����4�3=x{��v��\P$�H��L޳�;>49#q7}�q�1��eN�r��&DDE
���)��׉e�&ʢ��LF�׆�?ѥ��$ę���CW�N��:I�#���S�\s��'S8��\������XwW��2�SCИ���x�'%s,X�b��i��o���,n#fX���,H
�$
�,�r���ή���lv(^)�b�zD�	՗n�$�wL?�Joq����S`��P���;�����t}R
<�tY��/d���z�p��5�A�3L����D�jcku՘��ݤ���p.T8!�C�A���ͭ9�S�u�*P���XeJ���3�<�@���O��2��O@��!�5��d���Uq���W?���3E��aĻ���F�G����uRsa�<w��=P[]"@9F��RQ5�誛��]�SK]q�$�*f��D6�l�l!,�_L����z�?y��X%���sݑLj�����Z^g���(	>�G��@L���Bl�u1LL��S���>]�ď;�$�{�4ԁ������}/*���ghd�Ȍ��1��Sǌe6�vх�h��LYB�-��P񷰮#�N�1M>�ԏ
��㵒}�76(��C�� ,X�LxU��hc%�H"�Um_�A�w��\P�{qUU�<�7#L��&�%�����I5���f��D�>��@�Rn=@��M�+"e
��!�(��2Ț���Ў�ާ��ϊD:1	�}�שD�vlW$-���w=�j�d��g:��C�q��Q�?d�}�P��L	���H�k�7T���_L�k��$�kz��Z7�f�p�ëe���+��u_]��C����Q�%���H��o�n�;���42���$]�"M��"������[1�U<�-�ꍄ��	�K֒�T�6�wta�����o-�,��zd���n��$����c:ٸ,h�=ʩ9�Z������2I$��N�E��s�z�ER�b���+`��{�Ӝ :�q���\T�4�VN?t�|�1�=�&v��w�c~�vm�?����<�l�<��QD�O���Hq�q�z�B�q��XD�ͥ�b;k��[�GhuI�)�6��%V�;�I��
Ɓ{@�X\̦C�֤�R[Jl�b�kj-4��Cj0�	e�k@�v������a�05�c1-�\٢v�E4I
�\�Q	��1+]CR���+,rvf�*��85��V6��0���$%�RT:�BR�g ��)?>�I���Zu5�5���]J�кV�q4�2m����^��}��$�.TQ�;Q�&e�f>ВH$wt_�Q��vϦ�lw\�����$}���s`��(P���'Q�����/�B���H=��!2n�_�P��0|��>�]cp�gz�< �a�� ���t�z�R�v�<���I�G�Z��_�� ü�Ye\݌U�|�tD�nmpC�k��� ����Kr>ގ��������FZ����5
��dc�2r\ü��}�D�sݑ#�)ʎP}�1��@W��2�,��An�́i�vl/n��ɒ�	($�=����7Fc"�G%�8[ze(T9I�leusD:���v�·x��!<O1�w�Hd���!A m�H��Y�������h�%�"����0�:x��[���Z��c󤦸G����TG�ׄ�NG��?s�V8/3�CyÌ�	p��2�Z��W����4l\����=]`��%:Isy�>)��0K�Z}�=�$�{~��Bj�X!�zw��&i���{T%�çQAo<�%��3�Q =&�mN'eD�k�D ���,�$noL�"Z}�1�(�]��uo]��j5�Yy��9�C�j�H5��+m��G
��
���G��ӞD�O�>;�A�x
Ȼw�� �]W-8�]���N��Q�fIb[��c,h�o���=_~���4�R�av.yW��%���,!,�-���@��Ld��*��z��=�}w-��}�9P�(;%�܉�A��y����ް��w=�f�$�wt�m�Ô��S�A��>+��$�=m��"9�'��dX�\��^d��?�^cl�M��L�<Q�uw�InV̂Ǜ��_b����{����,����o�/	����+�y�q5p����7�c <Ysַ��&f�W]��s�ZB�~��1�My�G�X���$	>z�ZO�G�AQ�t�*�~竮�����s�L�s�ı$�e�̒Hv�鳕��:�S�����v���5"ɦ���A0��ǝ� �.�<J��E�v{�Z�$��t���e����=�pbW��A,z��wr�PѠ�eT��&��vWD�G m�������<��쿞��V�P�z�e��F��ZH$���fN_[鸊����e�$�t4�`E)k�C����MASo�ʬ��'��N� z�����aD�r(��V-eRL���95��6I��ۉ��|>�z���M-��x	)aո0�	BbZ�b�!e{7A#x�o�z-Cxt����5}q c�^��[�	F����xu˨dnv[$�����w�,�;'��ai<i̷?��<ݖ\�[3���a�3$H�tY�R }謾5w����)x!��葺_Vk��I��1ݽ��tv���`���.�����r����>y��7#Vz,d��ɧ���CY� �*�3�9p(���H����kE�Zխ��~����H���ДB&�E#��V_Ѭ|�Q�$z�GP��&s���x6KLozfY�G{��{L�(Z���8%�$r��CU���Q��B[�E%5V��Pi�M��uЀs�Bֈw)�~Qi�� ��Ad����=��&�u[�����ԉ�!�7f�)�.����" �PE�ߺd� �ò��>��ܦ���fA{��(�U	���s˯�$
��Ĩxgr`�w1;�2e���(��=���G��_[*�e�#�ˋ-׽���j�<%/	:x����3�	����bJ�z�%���?l	 �%uݛ���}�T�s9虿���;�1���m��Jsd�gNV����c<i۶�͵� �F��*{�	|���:}*���!8�Q�f�K�F�G�&܆|t=�L���[}��v*i�͋'��	��f,+���w��%:38"��i.��CE�)��R���F��s&,x�q�;HoIO\�4��[�
�ib�cB�
; ��6��e��h\��A��ՎF��R@��Uk�Xj���p�X��$�& ���e"Z���Ts-��1U.I���T�t ���*�@j�4���� ^쩚7f�v�e(�H ��6�ZЗ��Y�N	��t3��e��������\E�5f�K�5�;CiX�\;�Vʲ����)���J�cNԢ �0�(�ǅ�����$t7�*_ҥ�D�gD�I�o�e1fK�p��Yf�稓8�1��nd��HX çO��Lt�4�{�\JY�[{Or�2	n��5;������1�>�2�Ͳ����"!���t�,I��v���B��+��L��_D�d�Ot��h�rk�'&���]OmT�˳�'�6$)=1�%���^.��X�%6x:�X�\�uO��'O��� L�G����y��"%/ m��{�ÚL]�ws���V;�TE��A"$:�y�jUaHkB&d�˂�2����&4f��k�(\D8��k��<9���3}�X���	�tY�m�z��ݼ�A��d�ښ�V6�j��Pt�c0�s�E����Ǽ:�ʷ��,��on� ���'�v��$�HEe��P�|�v��No/=�	#�����_���_�L���{���3��G�����ŋ,[�U�Q���I�c�i��ȝe޷�_Lf�C�A����$?�!\	ܼA�� �F̖$/��	�J�6r&�{��KfOL�7�Ӛ����5�ƵC���T�X�s'�}q����ǣn[(�H���$�+���n��ܮ��NϪd��"y�9�%N�l���͊�Abz���׃̣����ײ)� E�oU�h��ތ^B�� �$�T�p�0EB;��7m��5t���611$:03��+�J��g���Ii@���`J� �k�2}��0������#	��|3~��|��>C)4�{s��l�
�������bY��B]�"{m��,Nm��$ʾ���<�3�32D`�����t�bG�ru�Bk�葌��a��̞���K�QAZ���4�馢A�̈���U�3ĿqE�E�{Y!AǩҶ��t�w��6z�߮e�Z+|���"�'}���F=6��u����L�Z��=vK.�*W������[+pya�ȇ�x�.���T��Y^j�;Z��ĺ��F����ܷΉ�����]�R�/I}�.{<�L�{ؙ�<��I�4>Q�ط�)�};�dAb��2{�L��N��T��;��Dx�˯�{T^�r��9�s�4އ�Cho�{x�}{�M���!;E�c����0�|�>��
�֡fb��xe���v���� �Oe�+�+�
�,Ls��gr'{/tm�>M���ly��8����?9ᅚM|���z'�h���8@��Q���MK�������1����ɾ���0N��V���Fi�gx��1�7�_n�,�m��s�̃JN�}�C�ȘN�;I�ɏwG+��=ƫ-�g?J�o����e�����Iː�s����9kHEו�z�I�S�.��.��u9�L���}w��x������u���έ�R��\�z�{�|<�{���b���� X�O�l׺ea-y�1�T���#�4we�V���jw!�����k�2%�';<6�JA��#�a9���}�ٸ�{�wWZ.�Wt�'&@Ԭ!��IIi@��OX"!ȒUT�q5�y[��y�Ҝ�a�J��e��EȪ�������z�����O]޼�׿a���|sYqz��)��%9�ԙ_v�1�VAT"m*�)B��ΒO��}�w�8���O�8�^�k�j��S�H�rY7$��EB�ʠ��+Me)���&K��tj��}}}q��]>��=z����H��*T��V���WSe	TV��q"�8�IF��T�B��
��]}v�>�z���qǯ^��"H3T�*2K��eܩ&Y�;�=.�]�j-jFF�T
*���\q�׏\}}m��z���j��#R�UQR���.
�s��"����
"L�Zd�Y&,!9k1;P���HIQ��G˅�'�9u�v�B��hG�WSb�-�dTʫ���ʹj�-e�tW�N�e��]4@�j�R�3�̄�		$�Q4���S�\@��+��.\J�bMu�G3�MZ+�>�E:��YA������(HOq���9��]#*#�E�H�D4/�O8�	Aj��O]1�cy]��MT��]�ƂvC{*�i$���D'r���O�ns��|<�� =�|2H6��2D�Mt�Ff�U�{�̎�O�{o�<�18A܇u������2A`k��NѬ3��H�K�#1��$,��,kg��+�>xߺ{ t~Sѽ1-����f��JG[ ��κW�Dr�J���ԛa�������͉pg����d�;�&�&ۙ�ꈘe=����nΝ��ұ�Gr:D�Z=Y���˧/5V>zZJe����.��I�9�4ȐG�zd�$��L�}6#s-@���1=�Ȅ���"$�UM�I �OM�@��&r�λ4�iD��̑�H�o�dN`����-6q����_zx�L7�Wn��D����OH�{�쥳�����/��<G��9�z��.�r'}��^8~��p$[�rþP��C�g�c�J0��׭q�2�ةx-���H�Y�����LX�bňۑ˙�'����Z"p� �ߘ����	>�{���s�Ǐ<H�zo&M2dAǞv���2x�5x���a [��2� a4�*��܊�%����-]^�F��U�!���~�/ߙM����q �[7"H�H��d���{Q�'����"�W I��{/���Aq	C���ze�B�#��NS _L�$�I���![w�Ȑo	��	�*I��ю���2�������.�{�]׻3x��C�
�:D��d	)�ԵȄ���"${���­NU���-�ĕ��!�� H���SA;�>�՛Pv���J!N�(n�ղR^t	�2��7�X��ؖ��lWnF$�gL�z<��<p����t��j4|�{�;L5N�_Qg���o~�����Ο����>'&'�z��z�Ʀ�W&C��Q�|PA�Å)`u�xg���xx�����߽x�8�>����.���a)��uf��ɘ�#u���<�����F�����X����ܭ�Ļ�٠�jF�MI\ͨ;�T��t�R.�=�˝v�0�El�)���%���4��&�0�0飣Wu�Q)+Ě���NԷFj2�e[�2�q���GB�n�!����E�Di7`�����,Z�ti�vK�a��X��A��kRؑ�֩m��!�ㇴPx{���!'	<S���� �����LP�ΐZ&�t�S�xW�v�*��4��fY$���u�������$��3>�b(g��z��X�%�wdĶnt�#�k����o*˹"[k}�]�xb���v�>J ��Ȣ	�s��Ǭ�y��3��dInt;���i;�S.�f�We�+�}P�]�H��e���`�1D���M,�k����|r�Sh�>k��4���;�90�C�DH�g]��@��]3���S�_��ReQd	���L�A�GL�E*~͔���)qrX���krڹ��.���Tј@����@�_��|�i
9w��35BP�:w1��!��I��I�.�u��l�r�"0J7��o�b��G;6D�F�qt����/x�p��E��N)�'�+�ą�n���w]������8B1g�zG|琶����R���������\4n�oO�,�Nu?'�a?��,X�c��5��w!�rXI�L���[�Q�T�k��x�ᚠ;*�>�O=2I!2�U�u�4E��1�6|�,s}X���b��o�������g�%לFV"Dբy���$+, [2L�L�$��H�G�����5�oG
�W���4�Ed]�e;�S0�u����N5"7��	
�p��z;%���O5#�YMB��ދ3���mM��Qܿ- ;����r�\�I�i`�(h����k�K�4���"���Z�N��"1���=2�{]�@�{#�א�x�[��@��H�H=u�$WHHtz�R��A�q��_҉�u�Z��OD� ��\��1]�f]����q���A1�.��.A�����5�a���̒u孛פ�P���4�P������=��1<�!��_��ib1�k�<T��;<�n��{�.�,C�U����]�FM¾���K��bbŋ~h;�����A#p��f����8<)��Ap��� ����yF&����$	��<D��{�qW=����ɳ� n��$����� ��E�|��,v� {\G��-A[Q��vL;��h�9��L���n���H�-��!��(�u,��.�b��8ŭr�[�G e�h_��Djts�@SB�����ԁ'ۯr�d׾����1Ndh���y����D��H���m�����Q!�u��Y�qI��b� H4��L�$�}���uJ�-9w2B�ʸ�x�'I��z=��9� �ݔ��b�_�Z<�)�&H�)nz,=�L���6]9�	�����ͥ]A�9��9�U[;9>h��lSc)m��P�j���J����؂}�{$�6.���˾�M���A���{R�]]0�����ҏ^������`Sz��6���_��D%��N7���jbŋ,CcD��	j���t!�y?�D�,{�r%F���vm��{� �j�eAۮ��Fc�Qϯ>����7B�a���Kmq��M�����΍�cWBZV=���>K0�h�_���9�72%�1��&�T�*�:_�N�
��S��i�1O1L��[�Be͵Jm��;�im�#3v$�H5���	�7#+]Ε2��޼�VH���3�N��"${ú�d��������X���y8�/2�Ӕ(S.t�="@!xr�C��@�qL_W_��m.�s�$>�A��bIbh��^s�/'��=��CΎ���>eqt�C�
/S�)β��Qb|�쬇^�"{�� �$�Ȳ)�z0��B}=��ǥ��ç���ULo1��2��i;{��8��4	��\����:�0�l�O�����e@;�1������gO�:�`R�	}��g8E5����Ǽ����8���֑���ikd����d
��T�u)���δ�c1���(�陉F���e�����٣J�]5U����*	RW	6X^)Wh�YS���aMj5�W��B�x$�5�k	J]��ƺf]��5r�h<.&h�SV�Z`I��&��б"�M������j[#�vcD��CM�&&��U+PƹeQ�2��eH.14���7)u�%�+u"�J���R�N5j{���K=��s�y?�SKLAȹ�J�7���c���SQ���$s���-��l!.!ʊ��Or0��R����D� �MĒ���Y�S�]�A�K���|ޭ�E�@�<�3�g��i�|2I9�Y�	�fT]{,�OH�b�-���3;�~�}�|���ZM���wA�\��ަt5���b��4H$wnM>Θ����&"�%P��w0�0�(k����:%�mc���E��Z�2ı�sْI�Ιb��ޮ(��TV��)*��!�&k�f�bB��i��&�2%��nn՛����ᓑL(P����� ��{2	���(���?x�#�.���5}e2M\��b9��T�:d�W{�������
��%�L��xz�r��k�6��R$���뾝{�r�M^�/��؇���P���i�c������y�Y�����0d��͕>�+�m�����I����E��{�AvK;2%�>^�\;|�.�=��D�4ٹ�D��c�i�0�b���*�K�{LfկJ��M�1�y�
���x[Y[ކ{�m���8��:�<d9>~�Bu��{�p'	8���F�~��~n3�d	m�ْX�ީ�eDğ�٘	�wX�-�Vi�j��� �ݰb��m1K4/\�4ڸ��a�� ���v5��șA+��B�L�{e��DIċowL�3�Br\�MTj6fD鎺� �y��"�� v^L�$��w��K���a���U|\�bA��_��,K]~�%2��͓{�3n��#�0��A!g���A��{�2NEzO�i�Q�Y����^��(�$i�{vl�����.0�4�bŋ-{�Dq=��S$Mw{�MDko
�HAp��r�� ǩ��}	G��>mD�hd��e��cLN�F3!+��oN"��A"�QE-��r9:l@y�)� �]	�������G�sWL�N_x��ɉa�팴ٻ�@P2�vlA0z~�֋��/�m�0A��ch\��e��b:ؚ�Rˆ]����p�h&L���mh�����<���u��%�2�$���,om���{�dI����ww0�JH�1���D����_�7ղ���w�B�"��Gk���/f��IV��F`�{��pKG�h:rPT=P+��$o��(�d�T����bk,^V�%�;=I���a����& ����GJS�Mt��X�K��i"Y"}��̂A#o�{SI萹H)�=�k���2��z�j�����77'�2r�� ��Ov�Ţ�h7�bYG�;r.���s� �ZX�b��bǉc�ن�/�'�Ђ��D����e���b|�&��w��y�a$����e.�����ʖ�翞���Y��R�jf��(��M�\r���D1.�1(E�,&�<�__����1���	:w=0I%�o�������Mⵀح�1nz��K[~�3Uϐ^.�"*���$g��=y~T������P%��n$|�o?L��L��`U��"�;2i�4��t�IB���7��tI&���8��٭⬴�	c��;��,_;h:r��<��1֢�ޓ�P8���N�~�m�3�wZ*I
�r<(���H%��3
�B� :�����2	����^�uI���e�1����E{:l�L|��zD�j^��z��"��ş�4�tq��;uG���u}�y����҉�O��v��0X���A{�ެ�{������L��;pgM��%	�����0
[��1`�@��/�wM�8��k`{6�ϽL��w=}��_:��C�#��� �ۯ�o���@�yqQ�A@��f>;� ���%c��_��^�~�q^��NK�����wK�|��3ݗ�险!�V����������^_w�a�0{�;�q��}��-�-�7S�;�uyOwI���.n�r� K��`�<:w��֒l���*�����Y���qW����Ё�$ugd�9�|&�ժ�4׮��#�r۳�@c������W!p��M�'�j2��::����'Mŏ����Qi�r��>�%��j�t�!������o���< ���`������aP�k{��>�V�j;����]�Fﰿ �3�w��&�ړ�6p����Q�����[������{��~�/z��яJ[��|�����������W��r�vȏAd�O]��wh�t.q��{����Oe�O�}�C��pYyY�O�j�=�mF�����'׸�L�+_���9��篃�q�*9�mLo��b�^���:�v���[���{��|�X�O����c_gR�[Ц��W�b�s[ݍ�������Qoؾp� �ՙχ0b~���7�
1�0`g	�c+C`��ܪ�����&����\�'��l�c�����.��ä����<qv�O�2<p9�%���j	݁�8��~���+�m��θ�F��#�(�Ё�$H��p��(��D�1s�[�$�e|�XNAm7z�OP�׭v��v-"���8;���t�w�a9�49�Y�U�NRd_it�r,���Y���������돯����Ǐt��Ӥ˅RBL�H���Z�\NS��z�SI"���������\}}m��<x�䚪�F�J�TK*O�>v��E��J�P��4���5B���ׯ��=q����x���u<�8jG"��˟<�T&g*.I0ڗ*e'i2�C�&v�&棨Tv�����������<y�owfZuD�$$jՊ��H)$��AO�ݧN� �
��.FIJ��M��B��*%oΜt�Q%P��Ad�L�Ǯ��>�
�����g	;(�M4�Jp�i�+�\��g""
�U����ab%�p�:f����(��Y	�B"�TS./W�O��"�Dp�o�VȪȤ,���s�<��s�)	*��/q�/Z��E�>�*|a������QȫX�Ak�UEQvQy�0�ݹsZ�G
�Q'!�t�&��>m�u��ֹ���KWr9�3Bܫ3�X�����F�p�LElչ����Mp$tSg7��9,�!k4chGb\��-���Gj�F��	��9eS+�@��&��#�dA����	�L��m�����mpP�WTTvf�����l��׉��� �̈.�%�i�2���X��a+�n�.���h�k&�d�ۮ5%��u��MeQ�2�h�6�b�WcB�c]6іh�*��r�LKr�8����cF��«fQ��)[0m*���f��K��U�E"�J�i�f���qi.L��l�г4�{T;0)�v�ɛJ%n/.��0��&]aV���[��3u�T�hG@#f����G:���bV��U��e�6�єbL1��P5��j�g�kt(��
�v�K����h�ºn�m�0TAuk.s�e�В� �#�Qݝ� nؖ�]\�M�
�%qDsD��;.�^��Ŕ�45)X[Qu��B��w���B��5lɮ,;B��M�!e���]3��i�L�P4%K.��x�n�S)�.�Q\,&���RWL��841�`F�b����3��.kW�Y1���-��]3��iE����TL[e���j���b Y�(��Z���L
�j�n����n�A�b��]���:�ٖR�]�0c�,�c0�1��2nBR��,%��n�6�P�֔�����[�飵 �i�b�MG� �)f�Kx��遍*h5ΰbðhkf��We����:�e��Ԥc���b�Q��Ya[�@#.��.�7Y])@����K�Y�e�B+��ͫ�ƥ)�]�K�]en�gde��,)uҚ,t��#f��T6Yj0m�-��ԎP��dH�b\��d��B�GfR勝��r�s��m�"xyO�X1) �u�Mm����U��l٭O^1��4nN>O5w*KkEoV�ݭdr�ɡ��o&ma��1���5-ͳ%�02\���vt��۬A��
�F1Z7l`�?��y_jf�g]-kS[	e�m0h�����l#Hl����M2�vriDrJ�����u�+$,]#p���i��D��*X��n��a�E��,����+`�@�Hj1�.��ћ� ˦�$������X%�Y�تC�����4�����BL��H�H�ؐm�&�=2K���sUJꘒX�v��&�����`CӼ��+�$I9��Opo
�;k�[B�]I$;�� ]�����A>����T�lI9Fq���E��D
��3��	�Ωi,I�}�̏QǞ��r����
��g$�wzD�����t�IB��}`���̌��S~���Cv�,g#�IbA"�jD�I�����7Vf
M=9Tĳ�]NB���8��- y�}�3���bM�a�Ou�1,I����޸�����ۜ�E΃���I �9� '#&p����
9��5�0ʦѴEj;:�cYs�׹����mq����ڮd� ���KL�J� ��$&W��YJ"��� �&�tܺr�I�$�[�.q�]�&��I����y8(��Yħ��~ag��X,���#��uvg|�|mʁ1Pö�C3*�SҀ��Wr��]�o5�(2[�7�W��1�a�5��Hz�H�����h���y�H�̷�/�mT������	(���fU�$�칂1G-*>zzN�ǻ-�,b��d�,q�vc�u����.��곮�k�Я�1ލ9��L2=K���H-۝;�Cّ5�d��2D�ֹ�+|�B%x�vm�Ec�'3r$�}��E{�1���f� Kks���$��ɖ75�]�{�J	wjw%�C����,M�c����-���j-�����ׇ�G?|�����#a6�a끷�� �l��� c&����+��iR�x�׋�4�qǷ�H�����9����aM�"vd;�[�W��Yy��H��[�$��Bb�>ǳ_�{]xN`��B�\@u@����ّ %��|7�M\.>�����!>M�/x�;v�Ww�WWI>�����)�1�N{O��]�����{#���)l~�I�wN%�=�����6��	.��1�c<t̽]zBW�C����vd�)�*֫.��F�Kٞ�WgD�J]�_�Ts�1a�'� y���H�A�����t����98�<�H��'ׄ�0�U�u-'2zD�=�)���r��Տ �wݰ�Q�]#�S#=�.{���$���Z���y�*�nT�m2B\�l�Շ6���qq��R%;:�D��*>ww&P�;�2�2^�ؒS$}�q �u>���V��q�y��B#�^e���z��t�	x��L�P͝/�+��e`$�Yy� �$X�祧�F��~��9�T��^��%�LNC�C���>�h��H.�_Fǚ�i^��4��a ��ɐV�A�"�m�`�N�Q"��y׻�}���&��vL�:"O��S�s �d���]��D�̟;o�ҩ56n�6R<b����n��v>�O���	��#�i�&�z	:<X��k}��z�����g���c�W�=��J������0"A�,�睙��]Y��HËSA��ǦH$j뗌˝�r�#͘��Y����Ok���wT"K�܉�$�⟟-fʸ6s7]e	�k�d�hإ�h�]EZbRݢh ������0�wt�d�hg��I=�d��2����1
L{F	�ڞ�̒֐+&�M3�m�Bw&P�=�j:� 	���{�,��d�|��2@�s�H5�N��c�Ѿ�%��K�H��H��U1譐��7��̓�t"͝�읒K�[��a2���A0�\�s���o
dL���l��׿�.]q�1�͊�}05�0���<uWT�@,_��#8Nx��. :��=O���2$^��{t���	���7v,� �gHx����J"_ϐ��ڛ��x���V��F�8�zz=o�*ɾ����d}�fr�����<��X�ԼhZ�t {
���� `808[`��d���[���8�8�ό	���فjn+�sD�nP��`ڒ�0�3���8�16M��3J::�n�򴷍k�YyF�u�F:���y���KqԪ�A�]+�V䖏6���R]�W�C1�W<WEh6�+�E�Ri��5֕˕��u��VR�5����Yf�Zj��R斸\V[�faMD�͕t��`�J����=���ؒ�mt"6���1Z�A���I������HÎR�c=����M���
��ÐK{g�Ma�w�����oL�KvdY�%��������w� UI��۵ޒK�tYX�3��A Ǻ�ZWL�@�M~�F4�͎��N@*ċM��_%�,o;bi�]��xߝN����� �g�2@�݌2��$���3l�ӝ�.�"!"�B�s���$)��HU�v�<<�D�H�Ζ�[<��&�x'��Ȗ�
��D(��`���(ށ O�����z�rrz׌�w�[��'�a-}�"I5��%��O�k;9H)$P#�����hf�Y� "�[k1m]G-"�ƻdդ �z��$ �'��2���"EvdH$���-Tb��9��k��2f�̂G��������SL���� �V�����E����r�4M�<�1�f�>YZ	��O���o��3�z��_y��
W~o/'УcDP��Ttx�GKUˎmbbbŋ�=r,	'6�dd���tb��z���]dGA��#"<�o]�M2ˮ�$�q�z��½4H���c\�2G3��}������G?���������=�X�y禄�"������c��ƌ��&���h�����B".�5��Q]-$C9�ɜ�˧����H5s���� X1����4.����L�&����&-��dΪ�0��,y���^��!�<7�"!�!GwEv��bA-��dH$��>@�3�n�'>S~��� �ue6�VYF�q(�Bz�q	�V=���lgn�P$5[f��ĀH�\Y�#3�a��89>l�%Y �xb��! aũV���zL�6��B`X�]�}������?㨾n��;��\@�^5b/b�d��[>�����_ߊ�vO��~��zQΞ���u?P�u�J Ko1b�ŋ�G��wy��+1���T������MA�������"H$�kْ쥝�wgQ��ݧ�ڵ��1��y����	����M�8�錦D���v�q���{I�̉ �͋2I9��MAC��zZ��A�E#�l�5L
`m��,,t��j�u�F�ôviF�3Uم(A�H��ь�_��7��!q.�\=�c�ȇH\���igl�M�$^=�����!�Gd�2C������6br�� ��Yk�CYaE�����A4A�k����{��0��QTc)�P�A.̉ky�\{��j_#�l[��Y"7�Z{s��$<;�~�ui(����Q��'�^��#��҉�e���P'}O�(���Y�F��>�2S�`�t~/ǡ4l�16�v����m��[�Y�Kf�3v�g�ϱ�|4��ӝ�!{�MW�Lc�0�7��(~{�>[�Q&!���i�".g�@"M�|��O�7��%�	�� �<=�I�=u���u��ڽ~��<��"����i��[Mm��6��Ƌ�Z�dDb$)ê�P��'�Ϳ.��_��u����H��Ċd�s�L�e/׵�&P=�3,�{�,M7mV�F
�
w����d���w�����z�E2	�ٲ�L�}] N1@˺��wp��)(n��4	e�\lÇ��!AGt�R!� ��̑�H�:2����&"��$�$wgH�$�}q��H߮���DaX�.���[p^��B��j$�I��� ��x�t�`��ъcX����	�Hpnh+={i�I��ejui��濌]��GTL� ��NL�̓-������]�d�G�	Ė:���'Ǟ���F�}�r�� ȿϘ�=޾V��qEҮ(mU�JmDC�$\��r����ׯ�=�M��9~w�8�8��G���*�-t�m�,�ߺ���c+���	Sl�h���d�un�+.veikD!p�뙴�9�V�d5{lv ���50�^e�\8��Si��א�#��H�4�0
K6��L�ab�Jhm`-��/V*B[�b�ِ!1�v��d�\�t�M#w!f�jA��!�陶ʚ���d���7+D���Z�#WL�Y�R覬ٴsB�s0K6u�J-��X�ri*�BRmMP%G�i�P0�@���\���e��In�{P�zf:��V���$I�GKM���&��4_���ƺ1���{��J|�[*�$�Am_��C$1 ��Ȧ���t(�k���|� gV�tD(0�'z�'�ؤ�u������*���b��mme��i	]��,J�:xÇ��!r:Eߑ��˩a$��b_t��Kv�cF�>�N�tϲNY�w�j��̄;}�ɪu[S�57=,㷢[/�d�on\��B�d��1�m�P"R���8�mam���j4�!-�ټBj1����㠊�k�2=��Lr�fL���8����R%�bz�<d��4{�(P!����Nb�qu+1F�S�׳w'^��\�)�+��_��x��K{h����#=2��*dÇ|���d�2��g����o�Qs>��,X�X�cP��I�-ݱ� � ��ޙ ������n��]{f��[��&�u"�z!�!Joft�9ܤ���D�������̏2@��Θi�ugXH���'zcRy�&/m��n	>�xca2� -��H=��<�����,��x"EG�@&���.*�B�yt��2�m?[�	1����<b�<�C	��2K>ݾ�ꖺ������=�u�����̵�0�6�0�\%�m�u�h-�*FV�0���o��=�s2�w?s=O
9Yq$s��M^�wX���f�#/.d�A;|���bK�/`���Jz�v�.��K�e� H켙 �j��.�1��c��ҹ�O�!
�>��ˈP�"����H#�[2A7ԯq�i�)�`�¯mM֣��+}����q�7������P�p��Zto��<��zt]�Ê�=W�sF/�ҏl����E�u�>����fVӛ�M~��C{Z�΢ 4p7Qߞ!����t��$��:��n��<=�ݹ�
'�g��
�u���3�n�%n�b {p3���i�~�9�f�K���S�8��M����Чi�.{\�~C= �F������@�����g�q�gL�7��˃��*�����������Lxi�0Ҧ���,�y�r� �k8�j�z^��/�l��\����ǣ�ٹ_��m���
�qN���>�{�X�xq������7�_M_�X��ӽ�t��hÒ?�e�٬N���'���^s���Q׮D��ߐ��qL���jR���ո�+�ٹ4vUU^;��^ ]��ď��ܯ��c=�/�s�ʣ^���׳}���{�Çzx'����'#}��sr?M���zi��\N��S��V����z-�ܘ�|�o@/��N���7zI�W>]�W�N������h��g�I�&pW:�#B���'Gz�����gc��U�J�D^�s�b���A����ڽj9h[9+���H�Vy������x{����2L�o�[ I�MY���G����`\�-�ydv��?m�@���b�9F���V����,A?���n���l�� �sݻ�T��l	;�x�Rw�٬�^�諓�!�>���zr���v�A��'=�Xe��UE�B�TUG�QeE�%J!%QOv��=z�����~o����u�d�j\*���D�Q˔E˗J��{���P���o��}}}z�����o�<x�M�Q�J%UH���Es��/("�2��9�p��r9��I�����D�*��o{�|߻�}z�����<x��EFI!"HFI	�D���	0��kB�����";".zʑ�T��ׯ�=}x�����o�<x�Ҩ"��QWLR�ȭJ���(��Y��S*����*\}�W#�`QA��É�r
�6GKJZ��#�	2"�B.BBE˅9��ܖB����S�}|�h��er	+
��*RB��"�g*�AT*�Qh&r�$wGTXjEFt�*����Z�	Y¨�1���AJjHAL͕�Qr�HJzl�P8��*#�fYE��+A���* �DJ�*@��P6� ��q�p�z| a�����N��TYX�w7�8wP����ϧْ�n2��Q,^��I$�VL�o8������:3ݷ�Č��ޞ�	���P��?��K��yc��*�z����z�i"s�����?CK��x}��3�=��ˋ�l��U��cL�s����Q5��Z��[y������WUl�3��-�+*�̑����3̑4��2 �{�fhN�e�̚b����!@ ���È�C�0!���<Lg�"6��|�A$��L�E��os�:�K�����a��&(szÌP��a��#gՂI|�Ux��6'^��K7ur�la��tc��:t9q
 �UOz-�'�*.oH�WL�!��ۣd[jd}s�Lr�B..E��i��Z�?xm�G�1���ԋo,~=�u�{���F���|+}���M���Y�8v��9c`<���z=��mbŋ,X�����UtH�}���A1�/x�����K%��cY^�ϘA*�2$����2,H�oL���ܘ�|zm>5���/�]ٱ��l-�H)�ilb�[15�٤v��'sw�D<8�t�ݽ��dɶI��8�|�gsϽ4���g"�"�n!v��i�4a�2SU��eC�xA�@��uL�2��û�:�ۄ�^y�1`F�t�Iq��a���*gt�To^W�Ik��<�R��� �#^�	+��8����|���yC:6:��q��!ŨPB��T�'c=�v��8r�9���i%~|�Aa,���Ry�"z�{IZUq����;_���D��a`m4�=��L2���3Xoʦ����vC|q�L��d�H���[������jk��=Nx��T�����٭c����N>Y���Ǌ;��&�X�٢���iْ��&,��;����"a�N���X����I��O�S_^3��c=�P!�=y3~��C�8��ׯ=_Q�$�4\,r�	cP�7lWW.�Y���i��s��[]�R���,��)KW�XItl!����� �t�<�A��ِ����������5Xř�ԋ)ps��au��X0eIP�)��ь�.F��͌�fh�m��[�l�c�g�c0h�t{8�܌\��Qf�)78(%�Sm/�|�;�g�..�L�k�s\Y�H��Y��f��s`GC���Y��2��������a�O��O��Y�H ��wU{�X͏VX���꘾dd�#k2��1�w����������b���H=;�)�'n=I竬Cf���9�C�8w$;W��dK}=�%����f�]�)��C�k�촞�ə�I����!�@�����N�D������NA ��A� %us,I����~;���9��(�2C�N��";*����ƫޜFe��f�p�!W�� �L���@�KWt'��{ަ��mw��������P0c�Ҳ�ų-t�tڵ�jK��L����}�>~��E��w�|�=l�$�o+�X�e�� �k��uϖ�5�O*� �A����^�HnN�/��'t!]��݌��,K<���m'=#
W�����_�;���2k�:����疳鳌���ŗU< ��]�h\<ߔ��l��V�%k���+��3+ H;��	 )y�6%��W]F�g�ÄK��I;ȼ/u��f��g8�NwH��w�(@z���������>�<(O�@��1N<�L�%�e̊��x�&Q�^7d�W�M����tXF.�z�Ywڙ-zI=��0D8�`��`�S�I��D�y6y]���A���fI���� w��,e�{qa��L箊E!� �g�`�P�^�������X�Ӊ�4])\:|����`��V|�}c��HIۯ ���.�'��o���t���5-k�\y�'�'�T��d�,]�I�R/ˮ��,��r�L$�_tH".c.��z�m�Z-L��襥��1	�^�^Za�cY�52�6�V,0��K��>g����{=sNG�����S���y`$��q��ފn|d�Ջ߻��˧�Jf���!�p���>	�G7��bŋP�;�H�m�����UYp�RN�G{��sY @�^�E�2	{� wOtt͋ɹ'�9�7:�fv���<:q�,ڦ�@=\��V:��đ�~8�X�t�$�����&�~���08p@��Z ��M4iڬ2��]c5 �&�f�B%Z[6�0�������Ϧ��[ ���r�@D�+���$g{��J�xuE��Kr!�e�w�'w�[��!I9Qf=��oa�R��w3���(k 0��W�,FW�������
oU�4%	������L�+�bD2M���H��5H�E!`;ofL3�p{��K�D�)�#
ȅ�yp^�ێ����=69�� H$_VL�d���@���Ɏ�v�'x�f,�xELϺ��U��{:�ד�w{�f�����߹���qzB`V��&��N�'�G� ��pŋ,X#��OU2%cgz�8$��Iz�WOD�d���5���nW�P%�<���Đ>�}3Q#;�	�9��(B�F��	WA�KHܤŰeq����ۄ�2��2Z �uB��(s���	�>w�A ��ɒH$ot7�V���ή=œd�͚d��{$MvU�!�a�Pf��S� ����<ǫ�Y!�'���˔�H ��.m��^�&��Vx=�"�'x!pjL5Ϟ�$�y�m��s.T�>��[̓g[��BbKv����e����aB�Rx�v:���3ޏp�r>mi�	ijˁ%�[:������O��H3�s3�|��K�:"��]����,n/y�g�[\�y뙶HRvv������y���f���yq��&�WB#=��&s�G��|�/��rb_����^ﺛ
�vt�f�*�O���6��-Kr��:J���<iG�"t�譧�<��(i�SA�պ+f|��8�8�z��ތL��u�U�$s�&k�$t���T�� &����\W���f�չt3��ְh%an�MA�ms�<�
ܡ���1��f5b[�[ahv��ܔ��L���LL�͹[j��[��e[�KW7.���5��	�Gc^Ъ����<����[j�G�:���Ye�\�۫cj��q,-�P�a��\�Įe�KE���r`�T,�a��B���ɖ{�\DD$���*祤�$-{S�m��]��Q���,��dȐA�\D5�iC^'�w0*�e�Q#S�<����۩	>n/�% w��$�����k�}�=�^x!�a�Pj���r�]D'�&$��0h��w��c��TJ�e}�$k�+p���!��4��y�A����Jaq�$����R����p{"��_zv� ��N��VL���@/��'�n�qC���)�"sٱ � wk�gN��پ�	(Xb�M���X���SZ@!�U��Kv�I��"K(L<D"����8O��C�!l��[�7�v$�dg{�q�zb���P�mf����I'wve���c�@��Iz�u�I���8b8v��A�A��a��t�n�T���k��!�}�+�ǏofW�l��(hO��^[4^�/v�M@�3�r��z�1���+'�C<�w�3k�H�����eb�� $ �鴇�e��A����0�ޓ�Ʊ5_e]��Ø�dn�H$�kk���n�����P�>��Νy>�uT$
��9�!L� dz�A��w@��u9�*gǰWdd�9�vwqܗx!pnh!++$�K�q��˄j�lW��1 W{�C|�l�	9����c����A	� HE8���9(��L�)6V�X��<�Jҳ]�������`<9wO��n@�'^ؒA���t��]��������_�r$���Z�>���u����/9��.��<��p�켙$��p ���q���ܐ�vO'oN�;�(�H���y�j�wb,༰�s»�ҝUt��L�9���/��t�`�{w�>����+�)UծB��{9m@�`�O�� � hb���1!2Lz�s:���-�0 �S�x�O�`ck]�w�^�++`����]Y$Ez�@E����q�`v��鹓/����-d ��P�Ì�m;�X�,��^ăx�e�P(b��ξd��@$X�`�5��%���8��*�Z�.ؓ�nS<��!4��Pa*��ص!k-r)!��icf�MF����z�^�h|��Nw�I���� ���M+^r��*^�{c���z��!�6}o�fʰ�'P�:xv����bAȚ���r�|��cG�A�A�wD���U��z�}ã�d������BO��뮀�bgdI=�Iq���=���b�l�FZ� D�zD�l��q��0�<�f�(8���ɐ��2	c���4|���Q����/�ѳ��,�gv�l�C��#�eY�?*���&]�hꈒ\�Y� ���skL�Q�{y���T���y�ƒ�L���H�l'=t��I�ox;�L�H������o[ʘ�2|ɑ^���mt��|?|��u��p[d
R����F2�ۚ.��xr�e�\V&��
#m���ǒm����>�0xJBq�T�	��D����C�U^����$ZQ  ������!BrjM���<�&����x��ǜx$��dI ��A�}*�����55/�wP�wx�o�� �K��i	�ԕ.z�)�~�i�dݾ��O�6z���	<v��7�[�s�i1�>{����A�w�KOed����:���y��kZ���|���X����Bhx��<��r+���� �5�3ޝ��w�pK�T�$�ן6l�ϔ������	�UQZ�B����_����4(������ER�q��[� �
�+A�����FA���+����"�������b0b������� A�b��b 
��B"�`B
�
�����`��� F"A��FA��� @b��F�b��(a29r�˜���s��1��#��6r�L�s�˜s��\�.A2&G1�����b�dF*������\�@3�)���ˑɀr���c9s�&v�e3�8 g����\����d��� �FA�0����`����\	���d0�Ld2�v��pd�r�2r�q���������! `�(@b A�b$D$b$@`�*@2`C8��!�0A���p���!��!��	������(y������@`*���
)���`��( �� �hHQRA��@`0b�@��"	@�U����U�h@��+�+�+���+�+���"�WT�H+�+�+���+���(�EXXXAZրt"�������������
�"���H4����"�������d"�
�"�a*���A�+��������+"��*�� �P(�"�dd����b��b��!�� BF(�
�BF(������o�(�}�ނ�H�� �"Iǡ^�����?����}�����$��������8G����A�I�M�������?r��+���?���?� DE�R"��������G�@�������G��(!EW��~�����I���8���;`W����Q'��F�� ���(���"�H"��+"�"�X"�b��`*� �X"��+��+��+��� � ��+"
�`��b
� �`�A"$P�X!!��!�D�A`�T"� �a0�3�"`p�@�1FD��` $A��d0�0�a��&�1BH�"$ $��H#�S� ���Ü���UEA�YD �QX��QXEU�EdQYVdXDU�VAU�dAYV0EcV,VY�� �0EbD�EoG��?��~�d�QE@FE�@	@g�>��_��~xH?w�l�9�~��DEWA��?O������y�E�O��6y���|a�}K?��QE���?_��_�2���dEW�?����������w��:� ��+�@)���P������a�?����}�"Y��<(�,��EV�?C�O�~�~�ӟ���+���?2�w��>���?0��~A�����������EWǧ�C���C��R"�+���6N!��?E�o��G���m�������B%�lQE�y8���?�X� h6���!~�܀""�#��� DE��/�ϭ�����d���d�Meb��hLyf�A@��̟\�~|0=P    �h 2  
�@   �ښ���h5@  ��Ҁ�Z4   ��5� [��EoU(	"* �UI$^�HT�UA�Plʄ�����U�(RR�T�!"����jV�U"��+�                             =       �   � �  �P�>*�́��8�.wUWJ�gF�+p \.���m[��&�\�v
�s��Z�\ ܶ����K6˙�R��T*��  ���]Zsw��b� v�[��=����t�b��� {y�� {7 = ��=� �`:{Xްy��`��I*R�TT)�  � >�        �f���se� ���z� ��`�0�y�� s� t���a���� ]�nm�^���ζ�$��(�_  ����aub�n�]P��땦�ۛkVڹ��5���x׶7w<�ֶ�#��r��M]{�r�c���R�׶�G����YCRQ/|  >         >�}�ֺjs-�.XP��v�H}���]� twv��suڲک֮ձis�u�^ǝ��{:� <�bS�V��WeH$�R�_  �={�Z�l��ڲ �ޕ�ɴ���4֔�j�U��j������YN�R\���&�)S&J�k)J��  �       �T{��&��9��5���
�Z�7V�ۀuvԧ6]���]�7V��m�w6���.)r��(.�V�Ӯl\���`�@*	UF�  ����e]���h�V� �r���WU�2��h�u�m��i�RUvW 9Tt��ib�m֧m[��TWu��H*
UPT��   ��        ��ٜ�8UM���+��t��w[cp 3W}�7�:jֺΒm����m��W6�[�é�v����
�RU*�V�  ��/��$�n�J��P=��Oz�֚͜��T����w ����5rݭ�����V�9�v� ���)H  )��J� 4hb'�R�IH  �~�M)P  ��JT�(   bL�%2������������ M��k��yƋ|x���Đ��%�Y�d���%� @$$I!!K��BB��I	LH		�\?���Q�
+F��e�_�f��YU��H��Ӹ<�J?n����̣{w`��Z�Z��͹�=6D#@�Y���2A��O^E���(LE�`�Z��V�5�,*�V��۫�Ӥ�5ky��ͩz(m���aܼ@d��Nڋ�D։��oiV�99s��$�Yqs|�'��s�����cdJ���kp�pm�mX|w��mgމ�4�w	^��*�ަ��!��Y��r��I�
Ϋ�Uz�!��M=ɗ�ͫ��6n�Tl��텘 i�"4�,CJl�I���ژ��Y���dE�QK�ΥeG��[*K-�آ"#u���ZԦͤ�}��ڽx�4��:��qZ�A�N()�Bܺ6��M{QL�|	��sRg-��.�c���ʁq]ݥZ�:�82�^�1쭉=6��zk���TI`d��V�(��W�)b�w��ړ%d�YvpT�ř,�l٧G��	5*ZxM�R`vV�%wwR"��Z���ūT�����`ge��l�YR�=5�A��!��0��N���ǁb �w�.���S7��B�I�w�n�J�5�&��l�L�Z��C�b����b��ɤ�˭�n�#(��7^�+�*9b ����-�tw4�dmA2
1j�=�wy��ɻW�/1Jv*PW�P�kM��%��ks A �"*�R9�%�ӑ"�/D媆u#��V�`���#\.�n�N�5��yH�!��4t���7 ���&�2�1�߶B��Z�[L���i��I�k�-5�E"U��^l�K�.�j��5��)4���Y2�)2V�6J*6	�z�q�B�ٛvkt��̭`��)ɚ��i�yY������k2�̦"�N=��T$�"��X�z�J9�EQ��Z7th�+5���Y� V���^�r@Ϊy��ڽʩe�`�tN�q�(j����\�5Ϟ�P������vQA,��7N���z�����2^P��:m�� ZH�����Xpŕfi�{)�.�]���Q����}X��ֻܦ[d1u��+Ub)�@W���,���6�Lf�j��[�(��{�ln?�!DS:V�J�˛�܏Xͨ"��ݱ���h� a�{�MZt_�q��T��u��ޮ�\�S��턲5w�\�[�p-��X*&.TY���z�/��R�
��h���f|*,��-^�h!��&m,n��Lu�IǛ�7��������;y/+hnn±Z�2(��'0��ZǕ��`�v��-䵳J�͚j��mek�(a�Ōݴ!�V^%u�Q�0c��hw)hVX�Cm:_^�+eE(�X�Tj^֝�gUAuq�9
�M"r`8�;�\yZC*��CZ)C-��Q*��@EX;��7��ZfI�.R"��� h��r�X��V(�$&�a�m̵����"&� �%]@���wE��n���f��YF��k-��,�a�B���ʬ.��p��m�f�1��F#�+&]�-�Mۼ�c9Or�]��Do�����$9�#/�yyw�}�&�ͳt6�8^��eǨ:��ua<��k`����Ӕ�P�ٚG�E[J�h�ͽͬxjLVqP����G`Wy� �рV>��D��T1v ����-���el��*
��bnF����c&��BV��⳦�k�MCi'wc��"��vig�R�lh.-�ņ�|��퓈d�I[j�2نZ
�V┤�f�Gbڲ�j�M�v�,�y@p�h^e$&�q<�%�2�!Wy����ݐ-[���̼��:ځ���T�aˆU��cVX�
Ζ
�r\\�Y�ÑY�e�hz��f�n'Fj(�Їf(D��+.�7���F����]�1ʻס*��]��0����ef˼[5le3z��x^G���7%+�l4!����	 ޷��#tkhDֽZ�
���+ yGa
�+&��u��iJ�bAU��w\�7Ϲ�޳�t�f��h��)�VnU��j�S��O���\�.�7�q�i�7V���/�zSS�F��Xݼùi]01m��w����İ^X�K)��A1v��WS�'-��h��j�`�l˪&�@��eC�L��7�&Ǭ��47鴎��Y��Mz6�Z�Soh�I�3fʱ��h�
����2���Y��e�Up!��aܕhl�.ȶ%<�um�u�B�!;ٕ��q�Cwe±y�6�<x1V�MᗅGQM[�a��ׯ�v��i7J���ّ�nɵu3c��F-y��彤	ʍ�2�T6�&��I�W�Nfi�)�z��/B��t���N�F�N4�4++a��wMi)N�\����C�n�D�0K���*� ��F��Lܕ���kig�͖ws�#�'V�T�wK�ݳF�Yx��$�&ʙ>y�(C�)���p��欚M�_<���,�D�}k4���Ųކ*e��$���9V���^Z�'mfX8o�O>�ڴvd#&]�4q,v�4u+�R�L4Y��Kh�@e���{5*tjnY�6�:�yG#� S �仐�H:ݫ�M���M^
�
�d�x&�R�4lflx7媝k�y��sZ�ZU��/]� �ljn]���hہ�����׸&3�ǺF�B�����4n3�:۫����2�*Sf��9�TlA��wFn6efLy�9� ��*�Z���Ekn�h�YW�%u����)�bWR�LK�;a�J��F�H�ֳ%�X�h���*�o˸�"Q&h�7�\5�h���3 *��:>��^�i�2��\m�7E@�P�%�X�os-`Y���� f��`���Wu�Z��� ������e�:���;k��1��n!�� �+T��W�dz5��5x���nǼ�U�̳2��{�VYV��X�^�X�׀���
0Ոl�;�33=w�V�p	ۏC���Ǩ�3�ƍ[6XHs�6;)b;sUi��=��<p�`=
Lqg6;n솩�ڻ�0�,��m$��+k���H��	�ţ6��8꫇2r��ݵ���YO5ˠ�b��((4�Ak�n�m��@��5f��{[@�=��]��<Q6����4�)��4h��"IU�%%	W��+��N_�1pWq��u�kMU7�v��@�ш��$���V#΅u��\��QՓ��-#WiT"� ���l�U�1�v�X�mZ���Z��h�jLYtKF;Cl۵� ���u�{Cm<�E�eD]e�����2ز�ELX��h)����±�\���E��8�0{�=��\��48P:/^�@�q�G}�n뀥6]����d�j5b�ͦ�X�{�2��]k�Z��
ʻ&���(�Н��5-GO7��Mna$ء>87o>���E	��e|��p��'6j�ܚw|���m��e�z�<|��6��a3HK��ղ���t��(QB%�sj3-�h<�nb����.��C��Dû��-�J�bic���]Zkmd;D��o���*�Nj
�T{�b���f����[J�i��JѸ��ۡ��(��f3�L�ǯ�Xפm�B̏!b�c,$��<D���7T��u�x.�A�D:b�㸝M��nĩT�0ʒ�[(�K.�M �����j�T1-�Gp�B��n�Mٕ���Tp�Ic�h�D�W���m�֡6"RaJ=klg�0V�y�enԠ�\�ѹG4�4\�")y�fV�o][�qw��N�pZs���״B]�,��e$UL�N�mZ��5�x���y4�/N���[�8V[�
O$/I�7cʔ+k/4^}�v����ڌ��j�l���nÖ�;am���$!b���v�§i�N�z�l�@EA�.ˎ��v�ֵ�m�9���69���ѧp�A&$��V�^H�w)��#�@�����۠&�4Y�3)��m
f� �E䂢��en	�F����`VlN	5��I���Ŏ:�*���;�/ %�	�.n�m�+ގ[I���㘳�[�3 Ϧ�v�U�P��̰4F�c�VK�jQ��(ѭ;qܡ2:υ�qC��m�m�:D9w���i�b+� ���/i��9hT��k[\ŧr
ԥ��[lri*�㧗��ֲ���n���	J�h�n+��T�&zJt�ĔÙN�cow5�0�6S#[�C���](�@q��Z����BO���6�U���	�۩,D�.c��nh�*S[{M��Aո��m�4�K���f�#���X��L��D�uy�.�� �Jڐ#.��3F��B��9Y�C*�],����I�y��u���˰u���i՘�Dl"��)nȭ��j07k7��]ǫ)E�[�i-X��Z�]��HkS�{�;*�=VE<h��PNQ�[����\Z.��Cj��2�`��ss>�K��GV;�M��>�*��l��*t��(��H-l#+I��+`�ԩ��s�P�Ԡ��vx�v���aޢ�kff�������u�@Ð���)Re����V9;u�3+1D�NK�ʹ�.Ec0Ղ��t���dN��ų�:�&�E��b�`�iKt]`�/�^��B)
��t�T茹V
�̼�f����rūv��.n62Ɂ��n̑OrĕY�kM$ƪY���B[��2Z�ܓ��!�h��ȟ|ݘ+�9�L7m��f��F�P�s��8�,J�I]^�ecZ�XS"���L��c��aĘ�n�o��:���e�rj�$ɒ�ư�ٗZ�Yo0IF�$PiS��Z��ȩJݗ2<T a��(�X�v�+��b�����p`黵WZaz��w��Pʙ��e3��W�`��7B "̽��xԋbiN����`���X͙Yuw�73+n�7k+@+Zc�Z+,�ۄT^6т]-��ả�
AF�tp��k��]���愃S,�9��I{N�(��Q�%��4S<��K���ٳ/s�q"k6%�[v�GIH&�^�80�ФXRk��
6��oc�U���L����K��ye8�b�s^6a�%TN�c�ܭP�	;�e�׹y`�FԻ�⥦�6�Nu�-��O<R̦/"��)�ƴ�&����z�bY-M{s.�m�%F�1�\�28�sv-ʲ<���zrDfbE �t9M�����FMgk]�Jf�[M �FVօ�e �����+�D��M�oD�֌��rm�'v12�T�,n1�c�V�J�о��i��̔���Q��W��\�BL��	U�[5w�̶�����'8�@�f^�^��s@	�è�ؕԂl�D9WS"��ch[�i�g����ٛR��M��i�FZ��*�?E��[B�\*�����Z 5�@��yY���a͛�����X%U�	����j�L��b�]�i�F!�jե�^+��s3���R)
��Lh�+p-�c��O6���n�B$�C@�(�����5�.VT�4+]۬+u`on��X�H�f�9�>M��ʰ�eH�jxc��yw�:�5,Ɣ&���řf5f�ṋgrB�4����Q�g	[c+r�Z�![К9�(b�m��z1ݡbh�R��P��~ȥe"����1�t0]
�)]���1Y{��ub�����`#a\5�/�T�SY��&m�	Y0n�*l�A�y��^�ekB��/H�ua�*C�LF���k��f�h))SN]
��RK�Q/�C��%깗ͩX���71<r��R�C �1P�n�[��9�� h���y���*�ח���d�Ӹ����C�r��*y�^�O)��x��y#Ъfsmo��܅XZ�����+T��}Yaf��a^��]�����M�A���:�oy�߲ƴ����m��K�ˣ���>�u�Ig[w����fn�w �(bTl���7X�sl@36m劻4�7�nc�FXb�͚�6j(���/-������kH�(k������,;�ʔ�9�2%
J��P[ՔY�Mʘ���x�P��c(p�z7գ,��}�����|���E��P��$nK�T3S6��D[ՙc2�[�6���*��F��L݅t�3H�w�����^:��#,�jU�Y��-[�Ղ�w��̷N��v���$���G"��*L[&MSue��Ӆ�Hs��+�z�4L�Rj�F�y���ڎ��f��J�Z�]��!�]�R�DV�$3��y{aZ[n��6��>/�WMY�`�j�TiM�ͨ�YkV�ld�mL���ɷy2h�^Fj��V �V�2zwr�V]��Zl#�5<���Tn��֎���8�v��5m�>�u� ^8c�ZL�@��lq-9�)0�8���ҽ�h�U�4%ޥ�������N�vFhP�l�A���q�:kf`����*E{�LQ6i���hSu$җ[m�[�ۼ������b�*-���6��� b%c�4*�(��V��R��e-�#[p�gC��[3�Iұ5��s6���̤/2��ۻ�B��Ŭ�X���iiVV��&7no�SJ�3N�f�%Ʀ�2NN��g㔥nU�	�1H�p�ɸw`�Xͫ���n�J�<����=2���5w�*^j�4�l+�h;��[Z%R������B�o9�l��&Bn4�/7r���kij�U�G`��J�0@^E�����cɖ�&�0i9xm\r�^\t���w��a�)-NY��N�T���V
a')LpU����Z��z�$��Ű�[�D��јL�V>Y���&��D�TMf3y�»w;�.�bċ�g(K.��v�fQ�w�>{W���Y����-^많儎P	;���x1��Yi�i�n��S{��NaE����n��u����WQ����ZT��>|<n��*��ꎮ�㫯ػ�..+��;���*������.�*.�⻢��;��*��:������:��ˮ�.�+������� �؄F��Q�@��l \]w�wvUwXuU�]� �I6��&ā&�&�6�:���+:��:�:���ʨ�;�������*�;�뻬�:���뎮�6!!� H�Bmm]�VTw]Gu]�Wqu�]�\]Uq�WYtw]�uu]tU�u��WUG]q]�u�tUwGwq�G]�e�u�wVwuV]��]�u�WVw]��GWuUe�U�E���hH� $� Di!�����@�HH� �$��߻�������s��	�"���)�qP�pAU6����5 ��Y�l�;�������	�on@x�hˊ�N�\�z��
�N�4޸\J�3�v͛�yddÖ�ɤ�(1������]N�k�nk��I٢�A�C�H�R�Y����w-IN��,\�����3Y���@K��m�؝ܶ-SY�gV*B>�}��b|����bK�mL{����u�ۻ||BOE���WK���gS�rӗ��l9�{xMґ[]�x��|�Og�^�Z��EQ�;�ަ�����n��\�vL������V�OrJ��)�3�>b�t�<��邳��g�S��3d띆t�؋�̙�sA7XZ�����M�L���*�H�m�팝����oX�ߒ�)u���9��dwRm��i�c��2��6�EP�w(��,��,܄X���>e��D�ːn����7R�q�X�.Ҷ'�������_W8�I�[4�zc��+S�3V��E��b�Vf��F��g-cUŷz��(��w��)N��j=6Ej�8��5b839�5!���������P�{����u�-�5:՘1�V�}�U�K��+6�]jStj����6����!�o,?UQ��X��+n���( {i��zﯮ�rT��3�vB��ٔ����#D��AJÙܱj��	�xRn���_):e��2e��Yt�#̕R�뭗���x�]9����o#���۝1Њ���5}8��튩	�Bփ�R�9ܰ�|7o�/R]	X]������۵b����5���v{����89�������3{����i����I�V��凬h1v���� 95cyRsu��.RH,�����T��*�t�uh<"<o.ZSEɵ�n�l-Ll\啜�3w3r�7x�Vݩ���R���L��J�,; �M��9Ah=B���v����﹩;`�i��_-�}��&�A��ފf\�&�fW)�#����X�C��זr饁���\%�ݰp�z�P��pn]���Ju��l�k7^u�u�]�
䫺��52��]ΐ�I������m�\}��Ąj�Y7Nl�kM ��[Lem�C���h,���ٌU�h�u{�A٠孟X�FKIj�`O�)������u�]�9d�2E��%c�W;�6�nm�1݈ɢj�l�J�ӣLÎ��c	�d�)�&��nJ<�����L�3�r��o�Ď��{˅Y�繂������Jd�_9ԋ���f�.�v���9cIۘ��o����6N��!SxWf�X��;��%��:���m���[�Z�V��[m�Z��`�>ىf^�u�U��̛ݼ���fP�f}��N<$v�����%xS�e�9�p-�5���f�1eqYw�6�H6�s2��˒��i�C9�ĕ���T�f��l�
�b�n���R1[.$���d��!��a��W7eq<����O3�'lVJ�p��YoP����Õ۪�9[�7���*MX��h9(tu&�B���zc��ʖbO�TVEq�}]1>��׊�;sCw9m�`˩)n��ǙR;s	��q�,&~[u�^�R���`�Y�R�W�'�25о�w�2d��}�wM̅ݓiP�
�"�Dbխ3G��oN �E8{7l׸�w�]��\�uܑ0�Tn��+�͡���hb-�ۏ��	���/%�a^���J;��N
����,��f��L��
�45��noqn����F����/*r�3�(�������u�ꑻ�z��VE;Ǌ�1r�er��K�g�&��N9NƬ�_Kf��V,.�v8���A�7��lڳrc��+�cz���󮷝�:z�a��%�c�І1w�n�-��۽�GdP����N*�:�X�)�ۚw2��*����IH����3v�#(�R�a[��5�o6��qn�\;VT܂8	�W�uc7�@�2��
p�ct���<�x���u��d͚�%v�m�lիs��7�P��IqY�۷F}�6B%,3\�Em�Zނ�LC{ʻ��.D��u�˗1���P�&����w�U!�����"���u������ɪЩu�KÛ�[�Y��^�͔�>��V����ıE)؝�����su�l���r�:�o3��¨=Q�@��yk�s%�����50ͣ��>E��m.c%�S�kv�b��|+���X�Z�fm&�����c�V�I]֚��c�䗎˺��LJ�l�4�`�c坫��2����*vvN��z��#���^f��Q���h���e��	�x�AQ{��e���=؝u�"�n���҆�̊�:�g��w��t���^�Q5N�J�M�`������j*O����FmC�h�͸'�--H�7�1�v	���!5�k����)�2�e+�eԑk����hc�ږ����v�2�-|�E;Ϙ���&R�XꈔO�4T���9�ync�Ά2/\��w"OL'.J�	��әʰhu�0�{/���5�a��N:.Άj�6�VC���(T�<�֛+UǘJ��+K͑v�ީ �;��.:����6[}e�l������Ԉ��q\c,
њ-��굆��ص7�P�\���)ի�8�ݼ�wk���u0�=UnչFL�޾��b��1a�8\�}�JӪ��ܯm�[LhL���)ǋ��g5&%�t`P����#�c�އ41�.�R���K��-hQ�;n�j��y�E�j
��	�&��iXu�@w�n@��L��b�ۗ��ZS-������U��sD9�f�����\��eC�����&�n��j,)Z�}����H�5*S�Z��7E��������P�/]��,q#9��Y$�UBAb�f[�Tq�3�2��}�b��N$��]:�x0�t_6���}Ю:��ÝN�i\zc�#�P2jYL۳K[�w�|�[�oZR-�8�<u�T�V�]��b]&�q�5��K�v�	�c$��5�k�)79��ͤ{zʚyE}�V�Q���G>�%ws���3Ե\�A^���E^�P�9���tK�v�q���%�^Vd������c8�,�h=���[��88Wi�w`GV)��MU˪��F�N�EiN{xn�QF�ˣ6�`kou��L�ur���b�kz�N�']���	!�\������u���4���®�������"�<��ޞ�ɝ)y�sx �]=V/P�`�v-�fZ�fG�t���k�}���2����6x0���с�(�\^�3���#��*�l�	�����Y�p�W�7r֮!K�)%Ch�����ӯ�}V	#d�S[��B��oMȗ׽z�M�3i����'0
��.垖%مv���c2�
ɰ7�L''f��I�u*ѡ,�Ǚ��J<NV�1��ޖ����x^��"��X�����_M�S�}*����GuU�o�aڮ���[u�9���T
N*u)���O�lY�e��ғXY�@�wN���a[C�-��]`Wu�Y��+���
1�l^f�(-֛�/���@j���\����`�-ٳI(�pj���7ƴ�1����ٕ��a6D��7׸n� �u�WZ�҈æv��x���M�X��|�ݫ���Km��"�2s�;6h5��mo9*a4	E�(̱�.C]s*����oQ\���K�j8��V���Mi;,pˬ|��57+��i��k�Q��GMwͫh��9-v6F�)���t�r���Iy�/����e��{b�Q�}���Ƅf�f�t��m�P�y���8���@�k��!`�� ��^�92c����e�7���D�m�t�b�����Gp�1�Պ(ج\m!\��\wSz�=�Nޘ������}7�<x��rFic�:����7�;��e&0��(��=�yڸ�eC�)0	����).3���]u�%���a�s�$cM.e��	��jӁ,bw\�u�f4s#:��ՁKWQU���͎��ڮ�n/���٣uvc�F�%��|���ќ�e���ϴ�kk�q^e�Ԣ��*f��/!x��1h���~��:1�]�U�>i+ۢG ���^n]�Hj�۔2��R���{�jA{��͖�ݚ���1h]��NWU�z࿪��.��wҦ�*A_NMIm,��k�e�t�_m0��B����%�)ov�k���X�Ɏ�l��[�3R��N[�F�3`�u�����L�7%I*��]b���^�ƫ��l�'���^aYBnH)���B�:b}ݝ�7�s.�r�Գ�|̣��x�6F t�9b��SNV2u��U�s	��m���n�7���x�'����9fbة��|ӊ;8C��_+��ʽw}A��፣�ŵ�JQo'���b��K���{s��3d��Ur��Z�/wR��QLvYm+T�2�%WQ�5�2��n�6�s(�ʴ�V:���G
��+,�p}���]vŴh��;U�T:�]4ee�BS}#o>)�A+-LR��֫1�f�C���	K)�gL�qVvJ�'���5�wJDx,��}�%��w�8��"�y���5'�}W[jP�{{I���,�k�������3qJ�H�a�-G�7OS���>P�l�_`�V��AӦu^���ꜮSL���4Y�,ǭ\��:��M�ܛ�"*����p��8�w)�Ⲯc��̵��{$.琢Ǵq���T����ά�A�n�_eM�\�J�
&u�O���Ԓ���Is���q�֫�fEP�#R����oq*��W[X/�L�%K��%$Mՙ�M�{3U��hf�����r�S���t��fq�S|�I��mgu�$�u�-�R�vO/R��F�n����ƭn��u�B!���[}Z�� mjЎ��j]�q����5T�Q��4tg]��9��B���7���c!��"�����!*��a�уm���fu,�1�/o_:+X3���犮�����v,���Z`��o���]�!{��2�Jb�5��������\�wn��6�5]A��G�7�Ggo*Hhڝu��aK�O�i[*���=�,RP�u8=5�y���:��W�j]�+�Wo�$o.�q����6���U,lC�R�gT:���
�Z&�ܬ�܍��3Zz+�1/U6n�Śؔ\��s.3 V^1Ckb��L��T㷐$R�/����ς�֩��Z�|X�c��r�63�E�h���;r������)
�v�n�������0�e�5�:��U%��Y�b%MD��Ø�ثչ�p��F��K�u,:�E�ɝ�̢�T�9�cI�}��Q1ccJ�Mš����l��U1�,������j�%N�i��t��Ê�JF�^�Z�+�Pu���'�ٶ�غ۫�1[V#<�����whdg��/�l��^֭vr}wh<���n"PZl�f)�ZL���t��y2X�=L�*L���;|B�M���X�P��J�0�@�yx�Au����p�dVj���oE	9�3ϰ����U��˔e�@���:S�.�f!��lN����C��WU���鏔ɯK#�{Y2�C��h�ɹ�N�6�U|����U��R�P�.�}�:�%X9��z�%WmY��r��q�±H!1�w�Va.�k䤫	EeC�+m;�<�9��~$���5��ޗ�u�zp�
�v�\��5�b� ����]��1ě˜Ŵ�Z�����ݗ��J��Vt�f��j��{-ɲ�������w]�.#������Y6�&ǜ[ύ$���#���%���J�ͤ�������OE��ywSVi�U�k�4]��
�<��b�v�r9�M3;[�pv�9b�h���K��\'��e`��9��j�]ܛ�7u���l6�y.�'�u�j9��G 8�ַhs�RH�Q��9UߑZ��WZ�W+0m��sj�`�U'o ;sI�H3�-يM%i�D)y��RS��*���}�{Dhέ/ ���(h�|B1�R�/���͋}�[�}�R��<��Us�͋q�D^4�^)0��gv�h�!/i��6�VG�Ni�V�¶ȗ{U2��Pn����T��3�D6��Ab�R���!�U��1�eK
l��h�wn趤��*ŔV��- W^ �viTAٱ�Ӗ3�z>X�{�+4����gӷ��alʙ�Ϣ���]rwL�m�o�5�ot�5KWI���da��\�6s!�S���i5�YYR֭f���+v���F���.�Z�Wb�<«�N�D�]G���)�cz�Pݘ�x�4�H��϶�T���7v��gϮ�s5K�_�ҙ��\E�HT��+;��YW��9��c�%j�'2�mt��a��.�m�hVKr���n|v)����ڽޤi�E��+��߶��T�m�wU��_e���y�F����(վaUt�'z�n�Bd��Q�����q��AN��Q�^��3X-��Ҵ���X�Μ���q,K/�S��r�X�{���B�0���ð<���3W��̱��˓e��-I�}TD�|���W=[�����A��,w|fb�4��J�fHIḰ1�����ᮭr��oiͮ쭔����4�F,b6q밂UT��[S�s^�fhOQ�!�V0í�d<Rin�3�V���\.
ʳ�U*�rt�{���z9��x�퉠t�و(�9ڀF#�9�1�&�gn��Y5-�#s����^�EX�P����|	�}����_2��Wכ̼�ł��)�(>�-���Ѫ��%�2���rwv+�{��] )qtjF'��v0&��wX�o��˷�nh���Zֱr��3���$�k�zF#p�����e�x:X��N�^�9�)EGH��b�5�3WC �o��fV<��jq�^>)�}��)��gv��dݙ�1�v�M�>�;4���º�N:<�fn̟a�뗭����6d��g�I	ZIeJ��W;2\��\��N��Ylv��\�]f{��npv\�å�v��v�A����#tk�	�[4t!<��Z�E��g܆�[�r��uSv)�WSBm��A��c[r�"w.-�'h�M�Vnz�S��+"ެ�(^Ki��`Z��c�K��Sݳd�t/F�v�uzn���<�kv��[v;�iܻ<{=$c�R�˲J!��=������*]�t����籘��M��v�/��p��'[o]���p޹ŊwGav��8���)b��u�	�\m��.׸r���;\�49kr�6��8�6;��xq�ݛ*;�q΂1ض���v<Z���Ջ�;���k���s��@ۨ�88�=Es�BK���F�>۫<w;	V�ոӘ�nE:9x���m��'uXd݇*ۚ�;YWX��<srI���x}��V{v��Ke��@	oO��#�:�B.�.1'�:4�#��V'aC�<�}h�w=�����7ZM�n��-�N7dE���[��/�Anހ��O۳�mm�;]g�3���-����{3f�Gaw��*gm<��;�Nxyʡ�^�+��-���ێ�.,��.�tn:�d�=�n2^+���xgI��^{9�i������lp��i�������M�{l��(��t�����t��m�lj9�}{<���L[GT=�m�8�k��:��y�n��=�FL�\�st4�=������)�ݥ�!��G�lٟhms�}����ۧc"�q�8�m��a��]��ӝQ��v��i�����]�\;�zƓ��:͔��I|]lm���*ļ�읷b�n�k�M���Vw>�����b�Jx��o��ޮm�vw9��D1���O'�yN�.1;�5�M���	(\.ʼ��i���j�!���'u����u]�-�9$����ܾ�����;��M���gt���% s��Mnz������M�om���<s]�<=��О4�{vL�K��E�yw�M�ڭvɝ'v��M�a;w��G�v�����l`�=�4v���n�aݳ��'�sv�4�[�۵�Ǧ��N�O�oGnf�x����9�f��'���l��gKlpV�n�%ky݃�<y�l�'����B7��J��DC�"3V����l�#!�"-g<�k��]�vێ���&#urg�9���%ݸѶM��.ڏa���"�� �a�Q������6�;�춀ɹ�y��{n�,�G��s<3��x϶E�2�Ğ٠�!u��n�ۡ�d�t��3�!���#f)k�Tb�O�n�Oe�b�ۇ���;kmWio#�9<�m۝��x�z�ӡ��,�]1������.{v�ogs��ۆ��F��3�y��/�3���݇p��]��t�)�y��8ttHc��l�sv��>Ю�dMb9�σ�U��͹W�L���$2��q�˅xzݮ�On�t�����v�A���<�O�;c'Q^+�#n�ي.�&����wom�ۜny�U<sё�wA&屵6Ŕu�6:7`���s�����X;�݊���W�糲��n��!�n���ö�p����	�z�7e�;�Y�	�f�����;�nɷ�wE�CJ�8ݧm�xK����Dn�7n}���ʮ$�x7;�ݣ{�o�Ě���r,j�l��;:�㹊E��|�g���gs�l\�zT�tp6u�����t�q��5�u́./l�����՞p�Ć����꼝Ʊ�����pV����qb�m��)Ґ:��b�>-�v;Q�{r�a��hz5s7{l�]�tn�'�B��*����k���8�0Vuq�v���tr[n� k��B5��g[�7�y�S��^y����������n�{%�����&�K���.;i^d�3a�ɻ��xB9����[l넭mV�;j�۫n.Bv�s�nW9��Ѻ5�kq����jF �nu>��l�ܛtqѻA���j+D�ö����<v{��,��:�kZ��]��.��c���:����G�v�;Q����ν&�۝�n�"n4-ҷ:ٸL�WY�>����^z����C��ݧ۵V�v��ϥ�j�ϨВv�kQ��e6[n읺��.�כ\뙦�/Ru�8��N� v���rM��xy:�j�޹�.��B[�ԛGc��S������x��ݎ+.�ֆ͚���Y��gt��N��4�8���3��c��ݗlb�g�Ǳ�m�3]��m�c�8�͹h�:��G'�k��r����SI���:��:��*<��B0Wl�l:ێ�����z�Pr����ց�=���!�أj㤍�����F��v����A��+gs���ݎ{�7��\�ayxe�퉹]u�`�WMt�"5twl:9%�Zu���!�qظ�:ѳ������^܅����\nrX��P�v�ct燫t{y�K���5�5��㍕����xneq��嫋6�̓��d���۰b]��ͻFB�[��;nk�N(���˽Kml�\۲����S�펋nt��dN�cNz,<U�4���Oq��u����;\�Fzj�v�M�[�亀;�3·:E^��7nꚎ3�w<���nu�[�k���^-5��+n{��`;v�d<M��t�5�u�ϟB�cn������6�m�;k��]�Dl;n�n���m��}�:��n�ѱ���x6܆kη����OZخ�]�K��nN��,X�>;h�n�ɰ����ٵc�;����6��+n�s�Mcɯ5���\�Y���f0�퉙�k�Q�^�+�܄�6�d����d��еN1�t��o;�n��#�;�5�W�O<�8}�g� H;Yz���e	ӭ���]�tܘ�s-�[���NM����Y��>6at	\Y�����m\/k3�/8���n{eb���#�=�G>��n��`�L�G+��u���l��)e��ݓ���v�aK�L�5&GM՜X���uo:%�x�.쐲�<j���һ��vcN��<a�ʜ.��q�qֻ@
ru��`L���6�%0�ۮ�k^��>V��ù�9ٮ6�k�{���<A��o �<�(��q��Qs�G�l����g���N��n9�û�3�c����\�lRۓ�c���@�u��&%��v���王=t�ۄ99�s��,����\k^�-�tqڵȂ�������#������9˝�,6^�=�s.���uLn�^��겻l�ʡ����e逸�͏n8�66�pH�lga��î�����c4�^ɧ�����m��Z(*x汝֝�VG�ں,�< �ع��˝���؝�M��V�v���DrqC�WHɸ')[��ۇ�*�ؒ��;:��[��qXuna�-�c(0��r\�!+r{����^��E��kk������[d�1=.6��>Gl��k9A]�Un�e�V�N�5��]���ǫ�����<�룼/���S��݉�M���֜l����^;h�^��m�a�7fw ���Ҡ�;��:�]gm��=q���^�v��Ycr�7n3�Spc�]N�˛�{m;c�,땠x���=�,��.�(l�5���X�9��N=�s�Ǉ�Bݸ�1��.�y�K-
�;uXGb^�s�;�#t;qN�;���nܖm��m�j���1�{ظ,%k��Y��C�
:��[�aŞֺݮ#�c��Y�e��*ާ�%����\��b�u
�Y���=X=��m���o]�B��s�z�<�D��p"��ԝ��;:��ۧ���և�j��P�>��<9�g���:ֺ�屜oc���Q�42��Rӷ�L����^�=��V�n����r��Hε���6���kn�l��F�J�d�}��ro �]�v�^��#e<�e�&�.��,�PHR}Q���F ���e�R�CI�p��i��v�\s��/m�n�%��q�9��ͨ3��6��-�!v9a��%��,��`x4��E��7E蜝O�p��pxw�r8w6��h�٤� v7E��%��۩�Kوf�:�yK۱� r�i��n���;U�%�Eq�Z�Ӷ�n�`�>n*ŭ;�� {s��n{<a�u�h�����E��⍗�6��˺������yع�l�Ξ��:;x1J��[��ڸgt)I���֖ϭ�׳v�n�u��q��[�-�v<�볹�l��Fz^[��ZK���v�0a�ܞ�q�G�<����/)�xv�(+��9ڸcqa7t�LXB-.ݮqu��i�n͚��<.�0b�;M�&�5����GE��W�\����a�B&}ۭ�k^�t�sv��(%ô�Kg����vn�;��k����=�����v�w'��Wt:ď;C�V���8ŋN\��]��LY��j] B���e��VǍ̡҈��lm��C����:y��ְ�^:�x;b<�^�.�웋�	K,/�aqz<�Qw�.ѥ8�Oh,u\&v���,9عyt�J��k�l�磳f-�0tJ�q�V����e�K=�7fwYtm�P�y(�������U�����s�8�n��0��90G�n̺Fx�\6��XzTw�p)n7�7<�9���h�Ƌ�bp{;]�ްgUp��Vݻ��{r�����[����ۉx�-ع�B�8�x;PsR�.G�H��s�o/.�ۧ
>�ι�d��nNs��r�t]�,e�e�k�v�����c�Ѯ4��g8��n&��۷kC����ҷ*�a�m��Ƙ������Tj� ������$�n�U�Ǳ��{c�^u��
��Txճ7���'��ɽA͇��u����]q<6�=��^	������&z�x{��\�cZ�<�:1u\�%Ê��m�l�k�����/:16wU���λZM�W]r��a��չ�6���\��\�Z���^ﳎy�gduE�	f�)�[D�q�my嵌��n�8�9$n����B/l��C��[T%=��D9�P�I#�MQGvvq&]gI���2ͺ�I�(���tB��)8�q'f�Pq�v�pf;g�۹8��)Η���N;K@�9m�������0I"w:��H�e���J�($:C���" C����p�m�:$��D
=�'!�\Np^݊;�٪�+-��+.N9.�9䒲�䀖`�(��ܔuvv)H ��pG6Ȕ胡C����$���{YI�\�9�rqv���$�"��'�A�'Oj��q8����$�8)e�p�7B��N��K̃��	*8��������g�e��պ��m�"�g;�I���nz͝�gu��0�br^�����k����F8.���]#��nx���;Xu/=��ۋ�E��x:�b���u���p��$h�]vn]��73%��ޓx&^�;p���1Uh���*��,@9J!4�{]E`{��7C��k�p�7WX�����x��vX��N\m�Ź���3�;\H�}��^ܽyr�yxlk�Ex�;���7�v�m�,��綡��ی)m��F�� ����k�:�ʰ��=a�}��xg�����4q��.t���0���ux�ݸ�X��.�`p������L�±��xu�!Cb�;�={[۸1�Dk-���I��V���#R��j���K���Ütn֣��QΫ�e��ݬ�Ѷ��{d78�1��-8��.b�^�GF3Ʋ�ێ97:�M<uvd��;���q����d�<n�ɝ���9S��aiA6�i�a��%]��ݖx�1/�|�@�$UEcW��A�ֵ�Қ��:�6^�p�)m����q��k�X(w$�N�����k8Rv;%찬��^f#k������6��q��*�SՋ�GG��f�v3����[7l*,5r��׍m�x���׳��3�l��[�s�D<���ݻ�;�n��ƥ�{[`.�3B�Ppx�8�8�Y���ק(�h�4T��m�0DnO��W�u�V�P� ��鱷<ǢSv����8����۳�nOX�/'@��;dT]�R����8�\���\�c�Mչa�k�^N��Z��e��.CM�������v6qY�:O\���8�m��N��>׍�l���n.�巣����ۢ��N���"��І�/@�����x���[�F��k�%Y��V=�)��9Q�@��:۶ۖ�px��tnzp�ͽ��������r|2��,<��@(Tm\`��e���z8�����:چ�s�o{���L9燏"9]���<��� ��ݞ83�we7a������ � EmO���	<*s�pyrg)�<�xx���=���4�zmA���^�< �0����×�ƶx<���X�l��K�g�v�8E�=�����˾4[�����ý��¯&y*����y\dy����pe7�<nG�g!�+���	�#!"�y��t?Z���g��s]ց;<߉��������`˳.T_�����L�&o�`� ��T(���T~T��7:Ō��Л�F(P����O�(Ws�T�e_�Wכy����^ʺ ��t�6:�ϗ� <9γ��7��G���O���n�Io�~�uU��/ �����o=m���F!�LX���~�y��A?=��������&���囚��S�߳k�WrN�7\�W���O~��:�7ޏ���޺���C���@SO����p`�5X-DV⫎���a�N�l�����#c&�2Gki㗺�����j��߾벶T�,+������MP����)������Nm睻�z6(
��T������F�g-�'���n���򋩸P��������2�ֹH��>bXEh�gw�]N�ey<vY%�Ȧc��ۤ�q���^K�LƹcW-�k.5� �]؀�����髲7�0�n�q�$�!��+�n��˧�A��7�$�D���[3�$���	#o|�~;�>K�@�C3Ϸ=/&ӗ��� �#������^�� ��L�hu�
 �~x0��wU_Z&��V��||��t���L��.��1�A��* �9� �g��dԵ�^��p95u��98�o�w�*+���E�Fї�s���yX+�tl�����Ϸ?;�~/�lXB�]9�D���I����>$'��B��{��v�-Hs7>�I����	���v��h��g�߱�G�p���ix��{���kd��=^~ѧF�Ԃ��������hb�J�JW[�/��#��f����k�xj���Y���hݬ��
6�����g��],�p��Y�2��3uR�o���~J���I4�7~��{; �,�5gVs:8tś�y~$�ly�H����A�B:��P���פ��x�k���w�=[r{\�6�}��n� V߼��u�L�.OU�`��tH߼Xb���Z�{��i �;�3m	o��}[�b��GT~������?{d�GK�z��g_����W�s�6�"����<�N]���gq�,������;'C����P�Q��e����3K�Ӝ��?�|���T���
�oQ����GTst=@���UQ\eu�&��ִ��+n��^ʥ?{_{I �M�߉���0�O�j?N��}�{i7�����@��W)���I �����k�x]��s�����sى��_ii��i��b嘤߽���=%��^v�$�g�ׄ���{SѴk<�PiQn�|wI���y��CM����*E�K�Շ*j���]�c��y{�*Xi��1�T�q��*�,�^&�M�ap�� �W�y����T(u��7�m��~	[�Ѥ�#�cč��f|�.^Iyy7������F(�Ԯ많	�,5�����M�G[Z(�q n�B61�K<���A�H�C}�z�I��%9�	;��ia�R���p�罿o�z�ϰ��eX� ]e��r��'C�����������c��O�ܖ07s�t{6�x4o}M�z��}�M��Ջ�j�7kt×���A��M�H3����՚��$Y�L���5�f|�����N::�v)M"���s�h�e�b�𱝪��ۜ�P }��M�m�R�^ G����+R5M��W\��H!yɛ�ϱ���k&�{����'�l���Ɋ̻7+����{/Z!@�'Vm^�B��K3����c�+���Egy��7B���v��^s����tW��X���&�YK4.�` &�'٬x�i���b���J��㙴��t��73�����y�X9��R�맵Fn�uv:n�֩엕�2OZ4�5�tݞ�9]u�� �1�ѓ�-l.�qv��#��{I��N:�n����l�<iꐦ�ܪp�����@�m�C��7P>�t1�i#sx���qon�t���v$��ۢ+���>Cn:zg/��s�󉣮�;�U�p%׳rEgq9�1S��.��ܗx���*�Y!"�Q4#�u��Ҷ�~n˳�h�<��&���$����N#��W8Oxs�E̯�\��o���("j�F�����h��Gj�m�w��Y$~��@!Oy�A��&EM����wg}gWo��V7�aV�;�ޖ|����&�N��y�Υ���^w(
ϼ�G��3z�[ל��Qi������n-2-��ɯۤ�H]�v�$��tE��!ލ�+��x+�^��F��t*����{3�Ƚ��}�w�|������n�I �s�3K6�q��U�E��r�UnZ���k�v<���U�mÞ( ���Z��Ǳt]$r>��3�y�9� $�z𚺱}��eIA+o{ݺ	'�$��H8�
-Y!�������Key`�g��ѵ��ޔ�O�P�n���4��_V�z59��p�����;ٖT���x�2����x"��X&z�ތ�������F4����gj���uut`�`t���F�#9�� ܲ���R]*]�<2�a ��t�	0��!��R�X��;
���w��{oI�lg~n�dZ�Ψ�������~�����k{���}٬�g��i���*	f/3��U���v���-�����{S�>3&f��:�JWkBܑY<b�Wn�9D�]��7j`ۄ��r���c]�޺-�̤d9�iڄ���.��U@�S�/}�� A��X �~�ty���r��`���� >9z�:��&�Q�l����Ep���#۰($~^���ϭ ����U�P�u�ǁ��(�D�,.��G��/���F�H7%�R�{�T&[�n00FL�˦9�Ra�yOt�8���9y��s���/9�f����ɚ�I��[���9���޴+��4[��� OĀa}�M���E��2�(�VF�������0�LZK.�m` b���w�w��5CXt��5?5T+�X!��Y�D匳����������OF}E:��
�{����!��Ѥ�OM����n�����w���3��m�s8<e���n\�<��g�{Zv6Ķ��~���J��$-���淪���{t�IOM�6�)��M���RƓ��f�m�Y��7<�Zi�F��\������ �������lP����@�'���I��gOU�w>�z-T
��EU+;����i#���	OH�]Yv��� �3|�I2zno��n�Z�JH�Wg��s"��X=�{ $ײ=�	&?MѤ3;���������HӞ�{�O��2�Y����wub�.�ը�z����	����P8����3
�ŭ'l��Wl�(�>$$>�Kףtx�}D�4	�#w}��I��/��A:�d�r���MLP��6� 
��նd���w�9>�~�v���c�h���ds����Ŏ9r�ct���f�C�>�񫪻4
�7j������'���A��h9����䡧)����������gIV9fg��kz�����a�v``�~��A Ó�,L]J���ٻ�ſ�c�
��MN���m5���,�_X�z6����� �H�~�a����2p`�
�nk��,�\3�o�fC�"�o> ^>i�B�.���^יI���{:���s�٘���G�&�n������ �rg=E���C/B̺�����>�w�P
/j�f�}B��[ 3yF�z�8rE�s�C����7��Q�h��X�U�r����_P��X��ɽ��9�F�&>)���"e{�w�.�7d)m�6�$wt�>��#W��]�g[����n���qc��8���7��#��x����G�n��^��1��4r�!��;���c&&6�1.�i��ǵ���0�ۇ�A�E�9�sY܈&�.�h�079l��&qb561vMV%��;��y(����;sct�n�7s*�x0p�lݖ3ku�#MIg�=��Mε�]<��^�8����Q$��rlv�n���Z@�UdQV�ķ����0m��?T�����r� ������n��e�۠�OŜ�� E�<j����ڱ�����Hԡ�Y�=.g� �~��@J/kt>^�Z���"G>�mp�ѝR��$�b�6�I��s��`���{�37��VVw�I ���,6֮�����um��P�Ҟ�7�����םTr�N��X	 ���h���ns�G�{ ���V
����oI$�����l| ��i��T6Y�a~u$��{tL��wN�!��7Ue&�����q�M���z��櫍���OU����u�H�����_��8׈�/��k�μ�X �%�]1�;ލ?�o�ê
���U��$����^�X�VhP������A?mz_�Cr�]E�sW�n8��ۋ~���XH��q�O�Q�l�rn��or,�Z����5]S�tWɷ��:��F�[�߆�`}�  %;]:�{Ѷ �هd�ݚ1��+��Y*u�Uv�9���X�O���K>o���s ������?Fd��������O�Ë�TmXV(��Z<U���>��� P�F��UC�?_�)ɿw�Q7�7�b�=(��(ԥ8Gۿ�$3}Ox.�2�%���74K��� �D3}����.�ݦ��7Z=�t#�Z�[c���Z�h�v�gс����N�IE�vX����n�?��T������I�;pi �7Ն�f	�r�^�ޞ���VCD5H���uW�P����M�@�7y�>` =�6��7�/�Rz���)�۞�E ��UU ��n���}�	$;,���4�n8��o�PRF�倸�V�GEG�m�ͬ�oJ�T�a�yR��ր�x�j.j�+�5���5���b:��X���{������.'��v��B�p�8MlN��f��i����+#�[{�e�����R���+�9�l�SX�v���[�@-�M�"nú���ü·2<Wo3"9]�.,2lJj���':����c�����ʷ���z�{����3�ݸ�f�7,�v��éO/7q�����ұΕ�v�`�0w5�q
�8�}��Zy�����nЙn�>l��t����v(�Ub�ɹZ�"�;"a�)9O/oձ�đ�I�h�:�vŢ��)������l�o�-]�#2W;���D7�lv>���;k���R�a.f"-�Z�h�C45w%䱡�.UԷ&,���:���]�����÷{U���$T+�;5�n�%��[6�+��;���7%��h���Z=��[�AX�)�ܮx9�utN;�fmY�u�Y[b���&�"	��*�,�;��qL�<�unmZ�ꁉF�%�(U��Wƭd��;��4ҖT��ޅ��h�[ќ��(�7w��7i�.]`�8&������K��ޞIe7��_[ϯ��4:�;�YF�g٪�є+���R���f*�!����m`�_D��Ө���d�oU�ξ,�8�MW�uy���gQ��|o-��j�Hi�m֑�q]�{as ����v�O jGS�N���epc.���=;r�A)Y�.^�Sk9�=Y�������"J�n&.s\�z^�z!?2�$�DLE�P�����NVZ �H�8��9�7i9:I"�J]�X�"�Z��8�&�$����Q���譵CZ�8󳎎:��N/.�r(���8p�N@rPRPG�ʹ��(�Ր�M��m���N��I��'bmZ�Tݸ �"N::9	�)�r����p�'Q9���G�tDz���YJ���y�^ڄJmnC��8���۴�Q�+
&��"Sl�$p9ƶ��'@R�p�N�'R'pQ�Yg$':��w�Qqrw%�p��&���(K˷#;�:H�+kD\QskNR9Hf盋�.6��=�М��N	"ΫN#��+�N(裻�#�;2�ﯷ��~b{��igɴ����V�����	�E]���Ww��9I�/#��I ��VI�3��"�̳κ�H���A#�msd�T�9-�����}ZM��{}���y3����{������k>	zkb`�����.�����WlE�ER��ї���;k��vn��6�*5jd,j��]���4h�R��Jkb�| �5�� >K�[�xg�OL��z�t��ù���Q����ct#��T�u����^���C�� ���@V��1N2^7���w^q��1�IcQ���m��gy�cjgl�jv�n�;z�(A�k�%��q/q�쀈�v���7�y����u��dՃ�>/M>�she�u{Ҹ�)����mP�&�q&eX�c5��ʜu"�C��kh�s(Q��Gi�x�V7�$Z��x���M��3w��gj��<�I��rk[݋�J��"�էy���� ����v��罹2W"+��̬ �sy��O��`:��|,\�.�!p��5��:�O'gm���c�b�n^ۖ�)��<ާn0��G�D����2P�U��y���T�	l�>�;��צOtM��,��F�Ws�k�Q����f�6�v�>�M�t�W��0����@ *���L
�b��M�r��j�"�H�=P2����<pi#�y0h$|h���ÿ�iw_o��'�s;���ɺE����IZ��8E�=�V�u�q}>$��٠�%�I$�SۥN�9�h �]�th���I k�w�����$G�L���:7p�@}��07qyӠ(W_y/��b3h>�MI�ַr��*���q��W�l�e{I<�����,�H�c44q;���S�Z�C��&�C�v����*���A����%���^Q�-E(4Ӱ#N!��#���zMi�K,m��Ϝg�&OS�-�v���ɘ#��K��*�j�v
m�m�l�^L�������1"A���˸wn�=�z��\�<#&i������6�uOg=ͻ.�,�&��qj7@O*�A���:�^���n���;>�C��m�kI3v��ۨL�q��n�:����v]��O��i��5���ձt�-�=k�ֶD+���d�^rd���E>�$
��j:�����	�B���3s����A$�eO^�}ݗ.l;ՙ��R��{qy�>�gB��k�[fbk�sZi�W�]�<=$w=��#��n�I�� ��'��9�9�ږO6����gM~�ϰ�I�jME���30!�ɺ���!PՊ�(K+�6wOo�W��/��2�@���piW��$�s��o|�ke�v�Rf���4�E� �j�]"�z�r�=nW��AXv��,��7��W_r_~�ةө;&���{��*f�xɂb����L�X������c��W�"�!p���\9���{���A�S����s���,0˘��o?�1`�{�F1c҃Q�Q����
`]��M�=���齽���6����8<h ���k�~;��Y�z˾sz��I�қ����r���r��O�uyf�L�Vr���P�	��UJ̴��I�Eg5OD��9������s;E�PDb�A��Z
e�bE��>�[X(�6����}��.�_����a�!���p~-UX[i��?������H��lQ�b�#E���"�X��C`I�Bw5�}~�~��!�8�6��v�Z�!�"E{��R1�A�����&�q����F���-�=�z�=���4�Q���Qm+a��%��h�!�bh�Pg�w�1�{�1��ܽy�������>�RV�`M�hn��޴���24s=��[A�1�z�^A�=;�se�/�8�7S�Yh)�0#ڌ��cX�Q��Q�{�~���S�O����tj�����������Egu���ű�:x��c�v)�0�D�P��&*�#�����6�Y��6����-�#L#E�;�"�X5���]��``24=�繹|������ƃn7�wԂ�r����ݤcƂ8l:t�^���޶�A��}�[>`F�ҍ{Y'�>�su���W�5�M���GZV�Q�b���vьCb���F1`0�(�k�c��g����w{^�.�>~��M�=�Fnj=�j���dh��e'�q����E�F!��F��~���K(�����u����*7�
W��P���� b�Z�F<߆���� �vw�=86��$ף�:�x��_[�پɟkU�e��O�y�3�25{�R1�Q�Ҍ"a��~����U����ѳz���)�6�w�O\��;W��T�>�� #���ƔMF!�!��r�`c#A��kޤ����_���w��O}�$��o��x4��n�6�����ޭe�z��Q����J5J7�����l+��v�q�^Ov��E�ѳ\��э�4F(Ͼ��ŉ�bJ5�{ԕ��>�s�t�{^��Y�?��߾��#c��\�a��.8�jͧ�����M�X/l�u�8��ݮțjadu�^i/�#G�~�'�q��@9��Qx��h#���z�S,`Fg>��j�W3�q�3�W9HƱ4�PiFa����bb���I�����浽R#��{��F)����W���4�;�}G�cJQ��w�[�q������A�!�Ms�f�>�3�[��[��#�C~T:p����޶�A��1g�;F3���7�_v�iS��1F��߾��v����<�Ѣ1��s���0�Cb�z�m�w�Jg��܆���X���Y�����j���}��ӌD�{9�^A"�~��i�c1��{�=Hƾ������z���o��u�1�y���-���K[�۷�֠(v�Ӹ5YyW�d�[�B�g����5�����O�h�7�� �����W;��1�1F�|'w6ލ�����-��߳.��-�#a/y��0k\����g�����.�##����21��7�����$DE���[{$?I����i�d��#�q��dCQ��E�Z�ݠ��z�ē��.�=��q��9��o[z�q����#<�,���c��ҌCo��R
alQ�Ch���zэ������}�:�8�=��1���(5��ԕ����/Z�v9$�۳��˿�H�!��g�fk����/�ˢ�A������i���{�=H�����}�o���@7vfG�����A�R�����ZܴF!��{��F(�F��~��Ɣj0"d`f�m�?����{ۻ��F�8�A��}� ��!���sԋx��<gG�I	��m��ٌY��ь׵�_a7��4�4����QcJ؆�Q�^��֌h�4F�����{�����g7�p4�6�5�{Ԃ�~�����5�M�֬lF��_(0x�A�"��Qx��Ӝpwu[���u��'��h#����
e�d��/s��kQ�l"a�{��b�G��2��lq�-��&^��t�]���h��u�L^�3��}KNe
|��vj�cfWX̎�[9XC}l&��;���r��r���Q�!%[eM�jHko{������q�ʽ����m�=���[���	�O�no!�c�tt��s��3�+Qo.�񮹪zpv��'�,��P{�[F��cYJ�[ �z�Ed{q�֧�5⽲X�h:�m���K�\�u��8c;��^7�܎�qn|	��j�lNZ9��y֓q�/c���v��:h�A<(��F�Q�5�4(GX�hj������#��㓦��|�|�S��P�d�;���y�T<�\q��ǒ��Pnև�?������������m��P�bF��wԋi`�`A���������������{��m���w�r�X\�$E���#&�9�O����[�OoV�2�/{>��L�Q�s��ϴ\1.7����i[�F(���h�!���{����iA����O���-�u�m�k�H6���+ZNlnOn�bFU}�SƂ!�!�9��[��&�?r�3[����_=�g�����{HƱ���^����Ɩ��#�1? �SvILDh��:���+��R}���]�6�l#�7Y|��!� �������6���z�{�L��|V�G����D>�D�#���R1�A���rM��-3,�gh�b`F�ҍF�~��h��0���{�����S�:����э��3�{�F1cҍF�����A�׻��z�ۛ���n��ܻ*��M�"��'avG]��x:�+/of"h��6�{|�xu�(@VOɴ���Ѽ�2�4q�����QyH���7;����l̭�����j�>���F5�(�Q�w�ܣ`�!⯚���pқ7�;F4bh����,h�!�o��==t�5p��ӕV��j��x�wá&P��|6s�雙�K���껭�;��q���)��*�����x��J��۫|5�{�,^�j��Bh�{;H����`FF�����6�>���A�!�N3xv�=����s;H��A7��o{��ksN�6X���ܣ�5ҍA�%w�[J�D�A�4k����[���}�uh�h�M����0�(5Q��+�������ޓ'v7�i�ٌ9W��oV�h�o;��m���W�E� ��A>����l�d`F�/��Ԍk�{�;�=���|�%ָ(�>�o�c�Dֶz9=�����orѦ�M�����)�#F��s�1�iepn�>;Gs��!�=�s�[��q�m�=�Aj��/��ԋxЇ�������~���
VV;/�m%,�7���V�q�lpv-���E�}TzK�~��zoOp���,���c5Q�4�}ϻE���b�"b����Z1�m��ϫ>޻�)�L����c#�Q5�}�J�l^r��7�ӏOzՍ�m�2�8<h#�GyQ�]�z�_{���A�n4�s=�AL�dC5W��cX(�6}�׭^l�׍���<����|��	ǚ��Sf��hƌh����1[��y^�"؆��FJ��k{�Ӿ�$1�ZC�nfch�ב3L1o�04�4N�ǽ��!�#M�G�hә��Y��������T��3t;n�W��Wɛq��w��o���X��6��z�S؇q�~���Cy�tW#{��ǳ[֋@��s(�9��]zs���!��n�]�ƕ��b���ԋbF&���粌b���ֻ����ilj4�j7��)+e�!��#�&Nm=On�``��˿�A�Ƃ1H>�e�<[��s�#���M_�h)�0# ��D��~���biF�J0=��QlCh�r�TB���hhN�A-M��k�G���A�!��v{؛�ƶ1���8�k���4��ݒ��ƚ<��{�-�&��{��Q��iF����r�``��Q��>�}�޷u��ۍ�~�ALCb��sԌx4�{c��e �cU��c0`F!�����8׻ľoY�R
a�(�1F�^�޴c�1�1Fw��Q�X�4�Q��eWf��}��s�3��}�X�BY�ڋ���2j�����y��"�b$�z��QlC��Cu����'��K��)�L�6�/|��6��F���cLQ�������h�f��hƌ#~��k���}��u��wf���6/!�h�W�FXҍF!�'o���6�h �}�z�ww�^����o��kf[[��f��;Z�����c��U9�n�ܥ�A��^·tc�8��O�qJn�e(u�ukVmr�>�� ��lC��>����x4���t�=�zc٩����.�?e�L�iF!����AL5�\���O�Y𩇘�D���-уDh�Db����Q�X�4��iD�o��RV�ly�^�J~�Ϸ�?�@}?���\vZ�Dwj1=cv�S�v.i�X�Q�,�Ea-U�����>}��	�_���;w��-�lC`{��QlC���޴b_/������ �T�}�}HưiF!�������6�,�c$�m��k{��4|4GS=�h�(0�_�����Ϲ��;���>kQ5��;��,�&F��C}��R�!�Mk/Y����{]G3�e#��ATc�klڴ�b�3;F1�M(�7�_v�m��F�F�}*�������4q4F!�DϽ���6�F�����J�L^wQ?�>�G	,��IcC�]�9�����������b! ϯ�^("B�CqwU�Z��dC5|�z��v�;������%mhiFa��ޣ`�'��&���Flַ-э�V] ���Pa/+�Q�X��ϟ���|!:��ld`B���Y�Ch0b�W{H6�;�$��sԌx� o�<��������nqͳ���o�/�%ي]�����g*�,2�&����`�S_opAN�b���j��)&`m�R�E�DW*�.Cv����t�M�.�D[�]J�Ax�5�A���+,؊к�3��ۍ:*��M�Y�J���/#}wZb@z3�ɮ͝lGV0��H��͒mi���)��Z���f���M]��,��G�]��X�c�P�6V�s{���*;G]A�0��vL��XW��i�*��R+��}/�ɏ*�\�xRgIaU���\�$�N��V�]v��N��'��p����bv/*���i�|��ɗZb��j]��X1*ΩV�A|��8n�qUb�]!����pGi�}�"��+��@����wk�VUJm�@����s(B�S��U�`8�X����ygk,���c#�z;��X8�Z%��:�,��+�M�.�%���8��&^���9�
{tm"�g��yB��in3�g)2هP��͛B�_A�݅�ӈ�BސN��Y�fPT���@Xq��P�����ԕ���p��C���3�.�s�3q�'x�k70���4�a$�:�y�]+�_0S�X�Ntλ��,��#s(�#��v�G3,�>�fXz�c�^�q�H$x�7O�觐KI�X�"�Y�h�)N=!��j��ͭ�k����=
��������P�hM���ն*�W=������v��oe�5��.Nyp_-u/@0�S��t��rዻ;.�Q��vKި��T�Gla��vT��V\�Ԡ�R�f2&m�B���i'���%8�:�mv�I\��N�H�䎂+�K�����Dw)'{d8:�98'"8=�m�8���(�8��rH�J9���8�9m�8s�Ϛ��RQ�TVn|dQ7c�Ӹ�:$������N#��:r�:�#� ��8�'�8�>,� �Z��E�pq��w�!^gpQ�_6��㭷��Dq��!�w_��D\I��G'yݡ�f�NM�
��@�J��)J�/��"�(�$J93m����e�BT]_6m�rw9��Gq�I�ڭ
::N;ktG	9"T�qs�HE'8E�D$�PE9$���Fۊ$�6n��8�{g�ǳ�vL:�wh�*�
�]F��WXֺ�p��h{cX��;i�.����g��R�m�E��*�v�.���.��i��F-K�g��8��n0�[]q�y�ltL�w�q�x:ݛ��&}��Ć#ȸ�f���Sۀ�m�]�s�J�`oj���7��^N�%�7v9���wg2ӫ���uYʜ�exY�q�F�֛:N�ZݜoN�l�ӄ�{3'��	��l�r��L#�]�����}���HJ�m��FB&_m�s�	ǵ�|�VT� D�b���>{Y��ˣAT��n��r��<<ѭ���v�|lA�.�۲k����n6�3[�vh��rd��h)j�[�]Vm!s�Y^��;��y�u��F��;���Z��BS.�c�����{pms�m�½�F�X��!�9�1���n����q�3d6፜��\�C�[rg�����>�n^lL�6|�Z�յ�[b�q;�������8�n�v�p��2#�v�K�d����Z��^�yGq�8�xL�d�������8�H2l7:�!���Ű5�MXzxW\۔{cB��֮��I��s<GI�#��w��p����Ln��b<(�n��<�$ش���<^3$R據��9�0V1b�[v���*�1�وN܇u������[�U//o/h�8'L�v��������DOnq����\c^^�c��U<����b]�nu���)aS��c/�%]Dj��읬�2Get��cnx|Z��� �L1a�p�n̽+��b�mxy�n��X�n�t��bE�@X˺zgF��.{2C�4�� (�:<�ĻO���A�h8��3v��y7N����GQ٭�h[m��N���n�2�h�����r�՝P��n�ǞS�Z�;�����,"O=��*3ϵ��w'��L�3������o'�s���f8b�d�A��dw)Բz��y5�U������+�e��U4Z���ww��GZ����Ӑ�sϳ��������z�yP�v|]]��F���.۰&��.kmԎ���=G&<�-��z3>�\�<��B.	��n�H&۷+��������*�\��G�p]�3�t����G`��i�8��B��xظ�����8W]F��G&�ѩ���ۓ\n�	t�* ��Z�;���Y7�^f	�{��[κ���q�X:julX�=�V�:�O�/lS��q�{v+l�H���L�:g���������ǳSz? l�U߾�1���F�j&�|��Qi�LCa�D�W=hƌM����N��[�f��>b�3=��ła�҉�����V2��!%�����٭�1�����z��N1��{��{܊��wu�-�}�#��G��ݴe�d`F�/��R1�Q�Ҍ;���9�05����!�Ig#'v�zַ�H�����)�0�Ch���Q��b205����F���.��/u^����A�쯽H,�!�"B"�^���Cx�;��z֤��j�c0b�/>��|9̝�>7Ck�(�Wn�iS���%����0h�h�Q����1��>�Co�oZ�n�x-���҃Q�k7��ƴ�Fs�ҊЌ$�bm%�57��P`�1@9�s(��'Y��?��}���Ƃ8�W�h6�L�6�e���#ƔjJ0=�s(���.��ǜM���<zO���*G<9��ї�ӧ/mˮ9��vg�j�c`�=�����f���FoO[בmh��Yt��#E�>�5�C`FF��e����v��|�n���޾�A�������r������1�owR����3M��ދ@����-�&h���>���wW�z��?���'J��Hv4Vm0������X������J�)�|M��h+h�)G]e\+�X��=�dQ+��ɡԋ��ի��c��u�s��B�Q�=R��1F!�K�~�1�4A�1A��{�F1��Q���G�)��}������ U~@�@�V7��nY�L�����1�̢���4�׿?O���c�eUWPm��m��ԋkJ5�`w�̢؆ыZñ����ַ�h�E���ޠ�.K�o׻��>#lQ�b��4]��kQ5������1��#A�N7�g��8Wo�>����W�=�D�G7�}HǃA�s�kZ�����A��/r��1���F�b~�;E������߹�]�O��Ch��W�э�#Db�>��(�,҃Q�Q��=IZe�^�����d���{���Vc�]�c�,���N]�9�n:�P휀�n�˰$?__[�!+iT�߆��#F���E�8�6=��/ ��;����[3�(�s���}����
j>�w�F5�(��`s�̢؆ў�y4N����=M�1�#~ʺh�(�F,/=��o���F}��ƔMF!�>�ٔ[#؆�}��\�'wο}��������&|!����S�!]�{57��6[}߲�f0#ڃJ7�g�����Q��C ��}�����<��x`���y���G�g��{��{�faOX��^�@Tv�e��V���W+��(���J	F4���M+D�p�^�����?4F(�~�e�6�5Pj>��m+lW ����h�*� #�{�� �^�Δ+$?q�� �{�^D���_i���`F�/~�Ԍi�n��}�{�=,��!���]%m"Y�o�m��i�E1Ws�
ii^��-1��λ�޻쮮�>��{�cF�8�A���v���AD_��R1��G�/��l�ܦr�y�5&ۚ�k�1�=&[�����1������ެ���v��~�}��֤oskk�1�L^���1�0#Q����we����b��W>�cF�;ɟ�}X��q����F1baQ�҉����Ҵ2���+��7�7�M���-24n��A�8�w^��f�쿻E�$�#�s�gi��d��\��mcJ5�a����/Z�پ�a�(�9y3S^Ѹޣ7���F4bh��W���b�/�ߨƱ�Q�F�����|>`q21����g���r�"/�ϩ�/VNh�7��{5�������(�:�>����k���s��i�lCbD���hƌ#DCDb�=��Q�Z�ݓQ�S�����vr0Y}cuՂ^Ӧ��_���Rz����ظ��y�"�̹yPf�A�,L��[9Swg1�s��|�<֎Jx� �SK��iF�u�� ���du����7�E��?W��lCb�>������S��kEg;]}o�p��e��!����_�ݤcX4�PQ�a�v�a�Q��Ԭ�r��˃\{ޞ�Q�rn��3�����#��W<\�2�Z�b���o���c��f���yh�Dn��R
b��!�h��v�Ɣj0##w޼���x�}�m��y����pD�E��#4�A�tֵ&�{[V��W���c10#PiF�]��n�WE���lCh����F4cDh���z�bKQ��r���޽y�������u�i,�E+@��KC`Zdh����4�"�yE����GW�>����ִ���
g������ԋkJ5J0�=�^Q�Ch���f�oF޵��E��kuA{+�5�]���#L[��|�~�XҍF!�!߻yf1��8�s�R^����j�Cb��}�F<CA��4S���=���R�L]�}�c1��(�6���Ҷ��w�����0b���rэ4F����s�^Q�X�F��(�o�?g�h#Hn_U���VZ��:8�����ھ�R;���כu�հ�\5�7���fr���A�����ە��rNl�f��k�M�(u<�������|�NyF9$+C@QZ��84�]dIv�e6Xw*tt�=�#S׳�����ު;n�Iz�s3�]���m�ϧ�c���\��nw6�-�D������fx �`�������Y�&��j�5�y��*��S��[y���L��q����v�׵�{'<ݣƦզ�R�����X��s��]��[i���g����v��V��"���C����&�;�+sG��*�ݪ��Q��A&1h��A֌�hg��l`�?bG;_e��Ab"�}��/!G��}�AL�fo����O�W��� ڡ����F5�J5Q�a�޼�ch����1Λlֵ��F�,h��;�A�+C�ݾ�Q|�^��~h�~�R-�ld`O}��1�m8�7ٟz�YPC��2��8����#�᠎h>��=kRnG��h1��u���bXҍD4�����T�6!�w����޿fjU�}G�1�4A�1Fw���0�(5Q��3�RJ��f�/��-�+�i,M�������;��/��b����[�A�h#��{փl�����~�v�m^�|���ꏷľb�����Km-���Fw�"����Z�>[k�ߦ�T�l\F(�4_��Q�XҚ�s�w^�^�s����	{������mN>��i�ࠉ"/���1��G�����>�β����덎7ŢkQ�tgn��m�nɑ�%;������2�EE�v�;�����[m������<Y�s�c1���Q�g�E��0�Q�LQ�_���cF����<�}lV�e�(�,aPj1�_ޤ�2�[���Y׶����������?�E���B�����zJ]��s��(�J���x�ܗ2�lx��o��i3S�h���SA����TTVi��շZ��^��$�H_xe��_�IF!��j�z�m�l�`F�/�3��kQ���a��ﵝ���]z��u�h����nx�f���Z4�m��z��)�lQ�h��v�lCbY[�z9�eON��-��F�4q�_ݤPC�D�"���#qh=O�z֤܏kj�c11^_����]�ռ|���piF�J=J�R��(�Q���hƈ�Db����Q�O|�s��޵���'��-�F���3Ԗ5��~轎�l
�)q6�Ƈ�}�"�q�� �w�^A���=lc.�F!��v�h6�`FFj2���R1�m`ҌW}�-�m�{&��'��˙�m��]�+%�-*�,=;��Ŏ�v6ݸ�m'd����!8ݭ����w�@�ֵ7�|���%U�Zh�(�F(�F����kQ���#��}E�1�����;9Z���͠��w�AeAAD_{�Ԍx&�8{sVɭ���o{�h,b���Q��b_s9��j�E�+~�yH6��1F�}��Z1�#DM��w�Q�CicQ����ѯo�et�i�s뤺2��|�9-{Q�&�ݘ��dh��Pbx�A�"H+�r����4���c�w[�����"�ܨɴ���ѥ%�<˺}e���J�t�߁7���z���~Fƞ�j5�b>�F^J(���� �k���l���Cj2���R1�m`Ҍ ��w�(�1F����Hۓ�jk[ܴi�n�y���3w9�/#a2��h��b&F���,�!��h ���=H5޺��~�|V��D�G�w�#4�a�y�kz����A��+���c0`F�ҍF�~���cJ�a<e�k\�sӢ��%���F4bh�h�Q3��r�b��1�����%i���<ϱn��Vs�2�����p��͙�����cx��%���<7��m�emXE�&�Pk|�q��[��w�m%�F����<h �$��yE�$h#�u�z�m�����z���5=߫�c]g�_z��cJ5�a�{�c(�(�8��d�{�5�=�1�D~�WAm�F*��&����gC�f}�"�]j0"d`OW{�1���h#���� ����J2zv�Z�q}��}��y�[5����o[�h-1w��(�!��o���A�b�Ch�2����7��"؆���W}�-���(�����%`�`Mo��rZM=�1�����y��0��O��Yџ��;�?��$~�����$PDph#�j���-0# 0#Pe���#�����YS=��J��T�{|&V�pl�(1�ope�m�"�[���m:`�d��^h9Uas�W�r�2�j��Q�q�$;�HH_���~�;��(���GrumMk{��4[Dw3��h�(�F(#E�;�15�/q��aX�{�{+������6���/��PC�D��w��b����z�ַ{�~ޖ��2��)acn�Kq\�p�]��(F�Ʊ��b7n`�:�����ߟ��\�y�����c��ҍF�}���i�LCa�DW�w��hƈ��N���F����^Q�X#JF�����%c)��'�ͽoz�f���c`X�?�����>zx˻sٻ�X�{���!G�G��v�m�����e�����`ҌCa��q˜��}����(�G8ru�O{f���E�`��U�[E1F�m����McJQ��k��1޾պ�����F!��w=H.��"Ey��HǍs�󚷧��=���Z�����c7�d&g�٘}7�jƔj4�����T�6!�K��ьCb��E�f��~q߸iRj2O�v�@�d�&��N�"t|'�ژ�r���F��{ C��P )7[�*��y{[���B��q9P��k��������J�U�o����*W\�����^ז0�v�����4:mvfy)�%�V<uM�����p�4j����|=Ϭ�|q��t��%%�@�A�'%����;�k
��)Ƚx���.�	i�h�������r��<�V�����6j��S���C��l6m8��i��)F�h�:��gn���8v���r�n�����<��mh��mw���R;vMa��N�y뮶�B뭭M�q\�ܱ�L�5�n�׊���� YL;a���9���·F;��;i��r�7��byx��F��	n�ɪ��Ș$.s��o�$W�m��$s� ����C�^��=�<��w*7><e��I��=߉��mD`�6	���ߗ���W�GZF��
Z�۵�=��>��=o�林��?��^{�����̲s�HZ^�L
����ʟ�m�>�����߉��7�4�{��A���Z5����f���P*,�n�$�������?�ن��h,�$z17�k~�~��)c꥟iv{��M����K>cBZ}�T�m�n��{�"t	?Ol���˔�B�Y�IZ͊D�K�mݭ��Wp�qb����X:�[��mwU۵ӧ��H �F�� �vpO�詉�0(
�=��4J̺����G�n�ԫD���$UGe�LH{�Ř���Κ�{
��Z�L*��3����mfu�Y
L�����Hi/yu��ذI����C:ށU��]wDs�&��e'����I$��[Ͼ�m���s*�I$!���
zg���ٯ'����k�����6H�d��g=ߵ �#Ϧa:o��:����M�$�h׽#l�I5ޝ��f��y,��I]Y�^�7��S�a��7.m .sX� '�o���/�ѷ���O���&�rZ�̚V8{qO�~�Uq��ֶ�;���+���@7�y��$�*zy6A%��7>fv{��s�9��7�cQZ@v�9뜼�]�v��3۵;Y�ڮ��
�N�2�3\,_ϣ�~o��	��_�����~߳0A �wI'��b�{�u�j�u���d$��No�M,���"͌?�����$D�W����AZcrn1�|@���:$�Ϥ�Q$��z�⣎����,&.���$UGe�� ����/�'{ӷ��IP�W���2�m[��wE
�c��� ڴWefU��Գl��M0+�&Y�'vۼ�u��5�+qÏ	ӷ���(�����+\�-ℽ9b�koG<�SF�1%CجC�\��;�kP��Y�|I���
�5��1�+:V�?���"6񉘾�޽�b�����%��.��V�t��J�}Ժ��n1V�c4���_�KGݩ�Y[+F�}��,�0�GI�+�ޛ:�"@��;Yx�
�4���$<؜����i�8��5�*�9:��e��7j/�R���ХM�=pja6%��tV�YX��m�t3
�p,��QJ�q�_�9����-��iu=��U�g��k33��F����L��Q��r�A�˵*Tŉɡ�쉆iv����6G^��vD��r���oRƩ�����].�8��]Qt7V&�xh�I�ś۵��ɎqwǗnKb�	���ѫV}�-��-�Q�Ց���f<O�l`�R�-fL�.r6Y��v�n�i�8ދ9 �#	��b�(q�G{�xL���3�xņ���:x�[��f$�u�n�5+o�,�R�	��!�c���Zϯ-͝q���b^�gn@i��qZ�TG.�-c�t/N	y���5�ٖ���Mwj<ZKo%K���.�j�ǫq;��n-a�W�Z�f���G1���6��[��v&�%�|���oq���4�UU�ώ�_j�AQb���XC���e��_�������߇ۿ
'����\�e��\t')N\��$�q�E���RBm���/ӊ+2�BD:(�:�*R���vU��� љ�Nu�%�q�v�I�n���m�ĝ����I�� \)AG'q��N����緽��觵�6��9."�� ��qr��%�qq��d�
r����۳�H��,N������è��Z���9:I
 ��쳉�,��	ӎ�N2�8;�K̢&�eYeÅ�rPpAq){[��(s��;����;���e����
N,�q:�JD����#|ϲ��$$�>~�.�8���﹙�$3괜����`�"�B�{����f�+G����D�^��`O���Q'��������cY��CI/��Ǹw����:�q���E��w������������)�k��O�Mi�{d|I�^]�]�I<��:M�d����xj�;f�Rv\��6�U�rm�ӟM'���m�b�d�7�>�L�D�[*���kx���^���I$��蓢oП�,[2�9��2 /��|O��N]���X@Áks�l�}�ޞ��y��h��}�(�k=����)�se/%�w�@ ϵ��xo������y�X	!$����w�n�d$��w$�HB��3O>�]�����1 Y�t~�z��ۗ�Ť����$�I|mǹ��$���w��D]��3�i�'A-E#�̬�:�*��'���8������Ùf�rD�2����9��f���r�����5a����|�k��y�~��⇿VVT���	�|�&���{έ�}<;ԥ�n�K�B�{��	$#����od~K���OvR��V�s��ܶ�x��vxp/7/6�Ks�ą)\N:��rYj�"���8����I8=ښ'�MQ'���i�=ٚ�a4�d^��~$`�j"iX�ݶʠ�U����Mf�a�{8��p���L��M~$���� ?����4O��3�Q�L/���m���E�&� ��:<�h�$;��hNd�%��^5}�vƑ)Y�퓩/�/�w�J�w+�M�}���o|������/(ɯ�$�{^2I%�{�	�i;�U/�Mo(�uW�2��62�e�l�;ܰD��s��<w��7�;�w� ���t$�P�=�IѾ~�ܓ{�,^k}K���8U�����K�P��Y��ѝ�u��%|2371�Ff�u t�Յփ�uu3s�fWp�/�����UN����A�� v��w�ùwm�ĖH�d0�2��!`�t��!g]�1�hd퍷Gk@�Gl�0kϙSqY:�����*S�������P���Ȝ�Be@�V�baXXY
 0����/g���-�3r[h�8��L>3���m�ܮ�0u�;)v=�����+���XS�uv.���9����¶1��Fn��'<��b�E^�q!��rt��Iaƚ���F{D�ö6Sy����sM�)�I�ۃ�������53�k��X����f��$�|�;�%�՝d��])����C��f,�G�w�ϴf�_!�-�r7n�tq�z1*�6K�״���x�d�I��Zvy�$�/��l *甯����߰)��F�pr։T�;��h@Q/��؄��ey���7��XÅ���g�n�$�7�ӻ�K�O��Z ^�sli��ivz}�IA�tѢ@4���J$�j�r�a�d���*oHW��b�-W��f}�����F�� �5��:e���0��0���� �������?�8�7�w6v���"�����F�u��mIi�����ܝ]���3W]�u�0!To\^�i�AJ�-�>��:$�K��r�$��M�����<���RZߞ���S�R�f�DV�C��wR�&'�˝'G��Ԇ��MN7Wb�!4Ե�ޗ77���l�7e�{�!N��[��[|�4q�9BH'yW������v}���IQ&���� �_��l�L������r�Fw��Ņ��6W�ֹ����o�M�H8*,��猓D���t���k��֞*�W6����Z%���q���f&A��H$���u$@����Id�V�\���ywI	ד��AU`ܦ�
�ٚx�������j��ɽ��7��l�BM+s� 0�\�g��������rBvI%�T��Hf�۰�r�:8[m���3qv�v�m�
�Y��IS�⒵F�>�?M}ܗ�=s�@ԾH�?m�S��]�#�&�����@|.k���Sjk��J�-�!;��G�'�w^�<^��{��{P��p׷�� ��=����Z��f�ON�8��Vw�$u�(����sU���'�w:h�I�ihY'{i�I�4iVJ������EF[�z��KbtX%l���U���/[K��Di�Y���=���uEb̢�A�/���|>ۘ�ߪ� ���ȂI���E�9﬎�l+�����k�n�M�/� ��ruH��$����2I&���B\�s��<���-r.mJ�%��Mb'�H��Ā��͌�v@�^��&�b�H��e�NyǺM/"�E�D���S�6���`�m�0�9�)��w>q��y`���"��j�'���T�V�i��W�f]H��L}�ں�H�%��}������� �{��� ���M*���_�N�`ŗp�߻�ɶ1�4I��?<�/�����2J��}a{;�@�-�߈G*��y01��Ś�=��К$��o!F�{M��=E �{7q_o���C(�	�*�٪*53��`m���k��v�
���F�$���l��TH�^�U�WD�|1Q�k+.�d� Lm���{�ݑ^ˡK��A�s��������Y�;t5��ڽ�^��W�� ���F�C_J��>޾��#����>�*@��=�Y��E�y�"�~�����׷�T��y3MeQ63��&��{d��O��m�@������w������#��פ�w`�YK1xx�n�=��=���ݝ�jy���W���9*����޷����w���$���hoT�Զ��h�k���Kg�����L]����F�a"�� D6�u�<��Jh�$�O}�Q$��׽����yw����=�
��/�h��u��Ft��� 
^�̟��K!/_7��w��O�K���w$�_,~���iv��न��Ɉ3g}���=���I�?Q3�����J�`�*b~܅;�=i�$Ϟ�;��Z�IeU6(Z"���<c$�J���fk�>�`O־$ֽݒQ ��<�~��o���,;ˇ���e�����M��^���#Z�r���b7wOt����������+.&Uv�\b�'*]��5�12����}��}�tM/����{n[��D6��c]
�"�z\jv80D���w=�����)�݈;�Q���S�=�r�:8ƌƯ:.x(�
J���n���<qr"�l�x�8oh��l�׬LaY��f�e��.� p;^]�{n�rR����mMB�x`�vr�Q��4b���Y#��n�a���猽9��ewnvݬ��U�7k��"�c\˞:��*��{;>�m��k��E�-�Cх�s$X�w���󤎔�,C��.{|�	�&�Cz,�D��ny��=槮�<7�<�j��� ���ѴNW���ʳd��tO�����c���3"��&��=�z��$�:��u':״��y7�"H\�c,Z�$�֝L���D�$����$r�'�W<w%;�w����I%�ӷ~�I@)���)X�B%?��'.�������+�w�{��s��cXĚ$���Y$�O����k�77�mk����W�Z�[oѩ*)�!�%��:d�Ě%�v��-����`V�n�&��G��D�ϯ̀�??{��w�oa7�ߐ��s�T�vX�En�h��[�g��9�K��2�	�"7[M�UT�����	���N=;�״  �rw>�c��I(�-��"���^�Q�ǭ�	">N� ,�,t���Ybb.{��=��s��h5b������ys\�ո�����k\�zՈ��� ��i����%����N/1�Y�[�2N%}����Mޞ=��\��䐒�W��-� ;���F�ş���� Oi�)�y�I����{܏>��oԪr�2�0;�y�N��{7�$�H��)�w����x��{�������@}<��Ū�2��o1�GQ�btߝ�!���:I'4�7��@{ϛj���w׾��'ˏ�#:o��&ބ0ϵ��x��N�H��Xʍ� ���r+晴I~[�!'�I�6�x^��M׮����ky�M�@]�9õ�g&�2jr<��jBrP�Qlv2 H^��O��*,��F�����D f���6۞=�N��AmO6���kg���@}��w{oj��v�)
Ah�ӞX��i$s֕�a4G������ 3��om� ��ٙ����Lq��{w�{������x.��������s{[ ^�e�����ub37�ݣ�<��-�K=�m���o:G�|��B�vF���5�f����� ϐ��FW�����-��r��oG.xI���ޛ쐾_}��7&�;w{��[�*�������z�^��=�I/&��$��7`:��x-���w��z|A}��f��oo��T�1B�fC��a$�t.�k�̾�"�����}D����h�G4�o ��ͣ�Yǳ�O��ݯ|m�~���r&�O��KY�f�u��6��.�Q��j�T�B�J!>utC}؀�*��&�� /�沍�ֻ�.���������llh��7]��4�Jާ>{�f�s�ʕ���G�o��$I!i��ߒIry4A�T������I%r��W�ˌ��Q�����̯�w� #����[q^�/<ny$��Y~�ш��#��'�.i�ʲ�e�ˣ�D&q�l�g~�>u�i���j��8k�ˈ_���ie���D��m�늈-ec0?zgkX�ѝ��蕏k�֤�&z��j�}��';���=�%�9��̮Q|��W�����vT�ٚ�c��Ff|����h����ska�a˶G�^2I$�~��j�4����~��=��ok��i����(�Z����qv��,�9���.L�]d�����0�����������?|�f}������� g���H��]}cΚ,�ɭ� &��Aڴ!�|i�dU�{���v�m-qh�L�����U�� ��� $���J$���Ǟ�ޡ{m`���%Z�SߙS�V�`gN{S ޽���	p��^�,�C���'�%"�n�m�g���{Ǯ���)cW0�㙛�Vq��"�� $���OQ$���I>$�|��3l�_�҈uM�Ѻ���=�+#�QB�x淞�ll	Ӹ���/%�,��t4I���h��徐	�~7�ͼ7_1G�2���y�=�ʼ啕�Y��'e��w~�X�x�f˕�9��'*kh;4l�4d�)
������7Uۻ�v�p�[*e�V*��gRu�qE���Z'mqC�p��q��EO~�=���lb-�QC�f*ǫ+���o~ ��jv�}�G��G��X�v^CSt��L�on�+fZ�X������k�*�eh''_�4�2�ne�1Ţ�ڧ�D#�p�;��N�UY�W���=�;�wn�Q�S	c��L�&������Ɏl�h�������t�Qܭ3��!�8�^'/O��8{�5��}e�qtZV�y�1���w7u�X�]z&ܺ��v�\�jݽ����`��vs���5Z;=��.��H�-��V#����Y��P��K�bW�pǬU���t�&���뷐J� J�:���_l!��Zo���.�l�uX�_n��C��̩%]�'N�Vt�]-�W{Y*�Nǂ�֑|�!{h�6%�a�&]��W�DKysV��v��R[�w��`\�p��)�9݅�'G}�;��e���Dn	�{6�s&���@�M*�ܽ�=4�:��#�a�������O��X����W�h��H�F[[@`t;a9 ��KL���:N�'E��7������3wb�6��w$�p��M[�_bx�J���{��e���T�*�]�x�\�84S�;o_+,�!�ŝYF޸��R̽�_n��r�ԸV͈`�(���[�3aj&+Y�NUƇv-�k��S�n#f\�}w�Ԯv�v6=�1�����i�iA�o��0n�llmE<�Q�Ǟy6Ƕ{Z�J'$��t�9":����P��'t���t������P��$N�;4����iܜw�p�w$/2E)H�$R)����m��Z�G�el�'��j����rA,�I���hf�MjD�'aP��N�p�"�� O;�m�q!N�'q
�ձ�@���u��(�L#���㓘�w8\Vu��;nґ{u�u�ĒY�iH�N�K�����'9s�'�<�vw��������8ڋFC�]v{Y��;sf�]�D�[nܱ�\�<g�y}Q�g�{v�tl�l����۷mыv����f�#�Ŝ��W����ټgv㷵�!M�q�:5����+�f��V⎴�&�K��㨢�7�n�����۟m�qf;����F�r���^�ۍ�C{<���`�n7AǴm���j�m�4u�a���:��g���n��e�p�sI�V!N�[{og�u�"󇗝�M��v���1��%�͹�t˹d8��Н�Ke��79��.�u.�jx称t#�������m����3��ɝ \�ܯ�%6���Sͧ��5G[)L��c�м+�qm��v� 1.�3���j�y�l|�#�9�����6�{ud��g�n�2��C�w�θ3��ٝ����p
�X�'G��C���f�u<�v=7\tnz�ޏ� ӎ�{9�O�:�+ϗ8��G�2��Ͳ7�G��tܼ���9w=�.9=46�sC�	"8L�;n\�y�\U3���L��ư\t��p�A�n6�w�����X��.�=l��ٞ�h�N:���>�8�=q�;���۷�-�m8�%q=�lf��L)�+����ϗu�n�m���$۶�MU�vZݯǩ9Y���&w.y��b��0V��e�]���S��us�d��T�=�:㭟vp���Vț�:��\6����1Oh��N���b�4���Iײ�8�@��m�W�/c�a�]����+� �)#�H�v�;��=�,�ݎ�Mzpk����=ن�e���΁�Wf���ݹݣ��6:=�brK�]�x�Ʈ�*/l�qk�;�.�ۇ�A��s�y��)K��!���a��/]��yJ�h��9j��;��-���n�gZ����t��p6�uc�8��{������[C�B�LgGq�:�v^�7EOB%�J�B�uk�u� ��� �w|���;������ũ�G��ٓ��N&�L�bF��7���yz�>�kr����s�ŀ�o�.�ֺ݉�q�u�t�2۞���R�#��5��'g���=�[i!��]������Q�v��	�<zN\:ݎܯN��a�'�k�fq��ӕם�5�ǡOf�[s�oc���1�:v�6qܮ�좮�çvA�D�zv�y�m�񌮸�2�뭷b(�[��; q�2�0������;]6�����Ռ��,�\4,j��m�sѢ����ӣ���~w�gl�Һ��p�g�@g5����|��F�����-��G`?�|��}�iRU,��,��M�\��L����8�x��s+`f��o{�G)��� �M��Ƽ�Gi��"��q$��Y���^�*�$�[�i�&�z�*J�ޓ=/$��Iog�w$J�~�ѩ�,T��uVNք�ҽ
����W:�#�;�f�� |��5���n��o/��*��*� �����ukn���v5s�o��σ��.,=7��~�����{��$�
�����H.����$ߧ�9޷�aUd�O�M�Ӑ^+9�
m��>���ᎹS*��	�
�G\׷�ו��h����sy� 8���m�	OG�u%]��*��\�B*�=�� G������VrX���d�1�ytI]Lw�w��˕wWc��K��T���8{b��N�Ẫ�lo�z����S�:jC���M%�Yc��a�{�{��aq�	���p�k����⾪���}��� �~�eπ����`j�9��Nz�����x��d�[*qK%���$�;��t�$��V:V�ݩo��ܒI/�����AOl�В������ȫǟ��͓^��M��'K��:A$�3N���-�9�sy�ݚ��;8� ����Z��c��C,�S���{d���9�ꐮ�4�|qǌ�TI��{��~$�-�"A��y��VoY�U捔b+�r"�a�ݍ�Vk]��O	t�t��Y�h_]�ܘ��>�U��(:�j�<���Z w\��  �-�%�^;]`xQ�E��D�.� �XToxH�8���	�'S�"��~k��	;���$�O�zHI�X�s(i�Υj-g<.�^]	��@z���ŀ�7��{�[�'�K��c�YǦ�O�ɻ�)��ϥ�S�\�)kKk>��r;@���<�,)�<�����
ϵOn^��/�S�{��b��7�x����9kI G�g�6����w{ny��L���)K�zi����,pŠ�ǝT����'��ޒ|H�׳�29��&�]1��O۔�2*�$������^���B�70׈���<��Igc�$��qo��I$U��t��x�Ԝ�j����]������I�z�v�1K��ĭ뮋��&�M�.s��蚵;EV�f��6mo���&�4=���k��n��9��}Fs{��>�wٍ�o��������E}�f� ��%<��V�v������h�[��d�e��Op�]�]]p������V1;�oj	5ܚl�$�8���~r���~;�hs}�f�@ ���fi�y՜���BF<o�2�g�'�^���zH ���Ģ@47�4�?On���
���K��̩�Y��+w3�K({* ���V�,ݵ2��;ٞ��ԴҼ�X!7}%h0��sB��S�;�!V,|�,��ޟ�S���}��a$U׮k��;*�:�ɉ���� ���ww���gd^R޾VI�I(�D�5�Q�A(��mu9)�Z��[5t�Wd���N]���u��e��R�l��g��y���Q�N��;�ڀ�}zy#��s{�`���D�$�M}۾L:'|K�^���)��3� ���g�J���bj���n�}��� j�3�ٓ��I��C|�L�D�=��n��D�{/�^��~_������B������3O��0 s�I}����Oo9� !{����s�1�o���P#�H�:8߽{�S��y�:�$�Q�'L�$���i�%���V�6��"���58�ߥ�$�:A�3����` =�ͅ�N���>Ͱ�hD�>��6H4K����u�z�<G_������@+R�n�U#���r"ƙ��,����6�99I���FJ�.��M�)kܫ��w/pUC����{=�Ũ�/3��w���7t�0�O���b�tp.+Gu�;��듬�=�M�R�6L)�B���9ۍ�`�U݋�dڹ׌:u��D�ľ�m�p�X굍�i8�g�� clg�R>�5g�l�n�N;(kj{/\��Y{�����WWjy��ӈ�v����E�g���z�a%z��{u�lu� N�E�[n����B���l�b��c�B(�k8Wr�C����ӹ�g���e�7����>����^0>�G�v�������i�N_���w��� ��o���_��ܢsH-��OD[^���6���)$7/u$qiŪ��j������ ����+�k�ÈI;���$�o6�}��jj��n�^*�:�-Y03��ϲy�s�������M�ܗݙs� FssٟA�3�流~5%`������X�bF�&�g�އs�xI��6��$�%��I	4H��kvB"�=Z��CO�V�=G<d�iY5F�>�iu^���k�t���w?"��H����o������]��Cd{�Ĺ`�e_7@��/+�5v-P�ou����[�]'+�M�H�r� q�]�m��<��]��)%#v6>~����  g��f�$$Ov�57�R���r��T�^ 3��w���98�p�T�I��k�m2I��y�7�2��)����So�(�����t�|*�1iޫ������D�Xl�����]��\�L�Y�Ķ!�10����}�S����O��%���������y�� S׸I3����[ť�4Ū��j��7���� \��7�H$�	{�H�3�Su{3$����>5ލ��r�k(���퓝��p�4͗��9� ˮ�6��{�I�I�I���[�#�7�s��O�7}���Ȅ��H�*��^��i� �K��$g���R��L�$���$^�ff@��=��O.���sE��EN�Ѓj�FQ8�>�{;����[f磕n���@uU�����V�$�UŞ.��n}	$
�m �$��dzZ9~�sy�� }����םY�`䔍�����*M�<�&I�����D��M�$ꓫۿR(%S���m���`�]M�*-�3�k��i� 9��g� >Hxk����`�8�n���C���<�R$���'3��ָ�k�#ʛfd�I�6�nYRm�\��b+a�e�˃E��R�l�/z�?| [�~H���=Ѩ���N�۴��FU�C,$�Q�B�|{)�t��2�z�����dIޙ̺�Oė'�F��c\Y��ў�7�){��ϱqj�S��.��%����$��o��:�u[���\�~'�d�M���Y�Ks�&�	��=s8*��*1�9U��D:��[����<�k]pY�ꐠ�n9���\�E.�������`�WuhS#of{Q$��7i �$7|�w%�=�	ui����u�]�n�Ih����r��WM��=$ �/m�D�{}�.��jA$��^�I:7|�q=�]���SPR�����:����)���>J_Wo�H$�Kw�or%�ice=��r��7e�vA��M�zID���e��ةZ�S��s<�����j+v� �ɘ� g;��`^��L9o<��7��ɫ�\�'3�y|[�T��L=ԕ����wv�WU�<��JG�����M�k/�\Z�{^�k�V�]{��K~~	!.�Yw�>�w&��[�h��c,��l��O���M!��������>D�s�̲I-�s`O�5F�ɷ�>|׃���
'e��~*����F��������� 2�u���i�n^ۻw�~w�;��
��3|�Ő@ ��=�[	/�@�f�;���C�;��lyo�[r{3�0�������+d��(��Mm��S,Z9s w���t��%�{�BI'�]����I���]�1�7���Mw��>��F�aG�3��~�*	5�� �5D��v��z���u�_��I-����H�^i�ɪu�ٖB�WA]Gu/vWc\�p�;��K`�TN�qϡ4I��5shI�ӯϳ���X�α� w������8��ݪ�;r`���3  ��=�'/u�ev�	!Y��cxI�n�\rH����wf�3J��M�w�|���{�a����o�wN�[�(�@�gsF3 ܺ4�,feU1�t��'n��.���{%�p�nj�c�����e��W},��W���q����n�`٭`Gmd7kg�ll.���;k�k�ۛ����]���9N��.�G��:mn���؞W��|�l<>(��vN�GVK����p׭:p��s�h�4;�7E�^e���͕�y-���g�\��^՛m�<u*���=��:��F�;��XИ��ӈ����i�ݺrvQl�q��n����]�96���NƦ���v��=�&���n�'a�ϰW�jٵv*4��8�҂{|⟘+���=y�oil 5��, w}���^C�SW&�^�~��ܑ( �n��%RL�H��%�_�;$�]N[;h�@�_y��I�m:$ϯȀɼ�Ue1ӏ^�;��wq��Ye�/���30=��̇�$�6ik|�i����` j���� >;��fC>7��F��#*�]!|�2��K�I5'�uL�I5��̲M~o��=�S|��X�����!w[�g�Uȷ�`�,���z��%���$����"���a&�O>i�I4}�~n�����D��.��/�1�%��w23�����c�u��nɝ9�7���EP�J�s��G$N���O!k�h:$�N�"�I~��!:7���O��T�����l�D������MkA��@��61�g����������u���}e����8�"�W+�T��ūs�;�㾠��/2J�c���y���ʑl�yuvk��ډ��w�Ane�/G7/7����tQy� ���"�$�_��$��	S��ȱ�G��S�g�W�J'b��;��YA�߻�� �I��f�3�Y>$�Os�7dK����`��.�^^���G����Sx���$���g�@~���ğ�'�y����/8����g�3 }�N{�(�eg,}t�����$�N��7�u��'��~4Gy���R�,�K��nQ&��:�{����2��l���E�Y��F=��\�������f��5bVJ�Rq1�-$+M�gW�,l�ȩ-x;�M��| g3���I>+��������<�?��L��� 3��s���E��H;SV��bB����o���:��ݞ��|�,߷��`~$W�@2W1~J�~w�t�>�x��d��V
����3���` /wy�ԂH��@����9�Ϲ��h���+��{�Ώ%��I�&���h����h�1k����.�.�0S룘#pgZg-�c
Λ82��/ ��0-��wM���^>�`s�U�a�lUsU5�ü�[	�j��R��Rg��3\M�����3����y;�/*�
�����(2��H0%ZHX��YY�%����6��_h�!h��/ga��ٶi�O}h��[&�|��G��w�3VYϬ])3,f_X�]ud���Z�Z�����v����z��e�өƨ>���S���ۆna�����+�d��WjY�q�ɯ[�O��k�QZyK���3��uws�<���]��FV��#�H3�\&8�l��aG{��7qfV�^�k.���-�RqP��u'J��50i^�U�0�ou�s�Z���Ui#��f�u�����A���]*|���|U%��%����9�����q�-��ME4�\,���W�o�S������y���V0J�ʒ'JlJ8�t���@�x-����1%�x�X�<�Zn�U��lgq+<�r�[cv���'U]��PsSZ�6Ӛa9;:���}��$��u�ևU�u��}U��dodě{{��w0:�^�l
�Y747.��=�t�sy�g�M��Jآ��y`�=Q�;����n��БvL��ZB�-�[�l&�ԯr���v�!�x�ma	 �)�;^ΏOi�����ءͩ�$���\�H�엝��&�7�C+/�<�T(����[�͡���& �rtg\�8莎N�#.��m�7��rq�����S��JYi�\qp) Ry�NrDyn(q!�$�:�#�㎜���-׎^v�6��Җj�M�s�!ggk;2��;�..�'�v��đr��ݜ���;�	#l�^v��w'	FZgv��8$��$�ns�q�tX�3�%����gf�a �e�Z۳�(K��յr$�*8�"����$�{6��;�"e�ͭ$�gVu&ۧ:�':��Õ��γ#���%�8N(J��'�ڴ�+��m�D����4�84�?���\��{���"��z6�/��đ�c�,��������R䝇�$���9P�$�hwF�$�O=�5�b�M�dN���I_]k�u��v�b�������;;�$7��,X�7(�K�!&�ލ:�@�:��+�-��V_h<Ҹz�ɱf�����]n��%����4le��n��]\���8d���>ޞT(��t~���{ϻ�	=;s@d�~$���/�n�gn����{>~Od� ���i�ؽV�9"�,����}�S��tֱ�����Զ ^�i?�$��nߛ����������rf��l�qV�vܸ.�9�l�I�^Ѵ�&���}��o���[��� ��f,�>��-+�$�E4�o-�g����.�T;�tW���Ēk1rA�I��?v�s  ߧt���^�TxJ��pk�C���|�$�]�f�r�j�����rE�\�xh{Y��mz��W<���.�pVo{X��|+I"��MG�^i�_��F�0��ݟ�`	o|�bvc��FF��\�M��=�|�Մ�/�zHI9~,@���4i� !Q	�V��V��ؚ�yv��t�q�ݲ1S�TMF�����H����e������$�R'7l��K��9��U��e�
|)�o3 >=ӝ�T>Ͻy�(�V#�>�n�7ތO�/zlkH���I:�O� �t�ք�K��s��H%1����ދ�����.ŇlN9`���X���պ$�O�o9	$�3��y��3�@oĠk��h�����	� ��J�Y"�f,^�o���X �J'�t�$�I�s��	/��v�W�#;;t$!��}�fhҼ2O�R�u�f�#��;���	���fzY�x���w���Bs~���I!�gn�e�O=з+}Y�u��9�V�\ʚօd��QϪ&�x��K	E�3x���e�*�U��`�kV9WU`�0�/��������,"o�7l��7��ݓ�!�j�� <M�c��{eܾ�9)�v+8$�[���Wd��vOn�Ez�6;����ۡ��Y��>0�7A��ۛ��>�KW�����^zr�z�<"��m��mv7k;��c�۲uvO<Y�v�wc���o�����G;=��$O7N9T��6v�K1�������16Q4h�jc+�����ܺ\v��n�B�׷�ѻl�[rcf3͚.-��E"�������P�� ���atܓ3������'��.�H��|�����+�g��~�IBw���U�zAN����u�=��<k����rxg��D�z{y�D�$ѫ��@2pKW�o}�p}�ߴ��Ej�X��ֻ��� )�oX�  w^,��ѐ9��rU~%��nh�j�Ѻd�
��bc�
�H���~p�L޸�s�>��$�/�d�$�<��˛�J��� $��=$����4tY�b�>���:kh���D���Mi�Wk]���D�[�$��$X��"Ď=� a��nV6ܺ�ԥ*ł�+T�v@H�Q��<۷K�Iڏ3�I9;ݻQŻV����}"�@ZZu��y���� ��ޫ��7��r�sJ&N暣z5��g@HG��f�֚��:9
��,v��h���uƭ����4㔮,�!YU�8��nI��Sc�u̾��X爩+!b�u���=z̴jZ
�I,�/�O�˦���B~$�~��7��D���g�Dq�x�C��Ac����>���G%���c׹��/�~�%�{1>��t��Uݾ$�D~�f-���U�ϧ��i�c�,��w�������^���  |vs�/�|�ؼ��K�_��`q�;^-㋜�Lr�X�X���1,�b��l
/!�gpZ4���(w��I�I��ͲW��HM���x���#�U�I��Żk{u���;a���Wa�I<���`z��Z�����"HG��.��<��e�O��l�hD�^��!<��q߶��ėyæ�Ɉ���}3q!���B�ժ$��ã=��}�P��d�KQ �j����I$���I>$�O|�as��7�W��}��tr�b~�f��M��6 ��=r����S�n��VI��V���~�N��F�f���"��K�	x5Z�y���He�\ĭ*d�$��Ӗ��x�93ذ ������g��o{	��\�ꌖ\�N�����j��ET�i�a�O��s�2M�;�ω ѱ�o/t�I:ӭ�Ҹ7�=�Ĵg�;�}u�c�ZϨ���!4I���8����_ ����:$�I{;�	4lw�t����Ľ�Dm�����"9�P; T^�b3]�[$I&y����*�ٶx����~����z�c�.~���m�{=������NP�nP��K��������|��'$#��l����޹�v�M����rSF�$�N�r�?~6;Ϳ��Rܽ-��wĆ}y�4+J�]�:��N�I(�fA��|�����c�EݜI$�;�B@5F�y�H����g���U��hKL~uK�d}�fsH���� ��Vw��@?<�Tlj(f^�
��:����``��5�=���䮷q^]���A�S����j����l9�d뻺S���c�
]�w���Ӽ`>���e��#�̯D�t�Tզ�m�yɤC�]n)�J(���n�"�IB��givMP�nW���isOB�n�<�	�q�n��X�:d�T�t
��UZ����|�R{�������*2nYԉ_D��d���*ȧ�y�g;�o{@ G��W|����r�I0���&%9�#L�p�1���-����f\��:��fhg�R�׵�2n�o�� I�sdn8F+�v\�l�f|- �	isZ	$�P�J~��W7<�+ਹ��$�;�f���
4.ɵf�a໽'Uޫ�����UXI$�MXĀk�Ӟ2I-�|�܃���0Ձ]�s�=�34+�t���A%qC}�tѢOķ7�C��<�r�Q&��:$�h���� �~o��%�S8�>ۖ��|������k#\�Υڔo�,��Gq��`�:��r��p�y��s6�������[y�k�ۃ�u������u�%����@���8��۱)��Ŏ�s��bzI���t�vn;ݶTZz�8��ϫ6S��:ܶ:�m�<�FgleӸ;��J�q����1@9w���wp�G�E�l�u��\kqx��؎C����8���X���m�7��zy�`V����{(���>gN=��<�<61�n֮�r� �����o9��fWUB����53�\X6I�a�Hd�vʩ
;�[m�nK��yDܛ�\�P�
U_�ߺ�7�T9KU�ӯ��D���$�$�����H�ޚ�(J�I��zn�)%��7F%�u��+�2����9�>��$�Db�:峣۫�$�L;<����I	?]�5/wm���g:�9��ؐ�ݠQ��ȳy��3@	g=���NZ��d�<���� 8���hb��������v]]�3�x��`��s���zX 
�ѶI4Io�� �c�ه�ͰQ����ɥP&.�],��:2ot����M��N��w���w�#a"i?D� 7�̀ #�k��LȺ��Y"`�Q�m��� �d7>۴�@ݕ��\�K-,#��}�=��gPI\P��No�6I4Ks|�$�Y����9��.ڐ[4��t�4Inw��I��y�� r��KU�1�9����9��^�qK�J���p����Qv�`]�`���������aEF���6�+Co�b��d��Ѣ1L���.���|���I����Q$���uH�N�^����9��K~���&�� ����w�$�&����&�4N�x�J�뷁j�k 3\�6 ~�ey|�_%�4r��6O��4O�^�][�H�c�����p ����˾w��;�g���f����	?k9#hR1߫�:1����'�M?6��z���hZ�׻����E��V�$���5U9}��9e�<��t��>jV��W{v2�mˡv^�(��+l��t��:�٩��LV8�����3���i^��o��~�f��@�.�"��eR�|Ǯ�1�{��	D�N�ϨiWߪnqBJ��}��� fk8��+�{��D�U*n֤�ALu�D�S�Y'Y[�*f6_W�r����h���#<g3(��N�� �<�|D�2�0_��s1[B�gW=�z�"e��)^yS�V(��Q]��̸���l����W�/'����~�=:FI%QM���_�{=�Pύ��Q'U��ް�������U8����'����[�_`� 3�緺��]�=�u���3y���w����E��1u��� g����k}*t�kث]Q'��v�$��|��A���s���w�9�}7�OmM�m���~�3v@�m����J䎷"9�+��7�G���0�}~~~X�>/��y|�a�f* |�Oh��9�̓���Ok�3��F��w�C��v(�2�^Y�ã=�р3m�x�fh9��Q�\�^�{w�BOĞ^]�1Dz�z�q׾°W����BR�h��OfC�>�9����o����
9~���:�tI=��� �_�}$$�fu�B�}�e��[�5͹K��Ii
�Q$�]qD�$�{}$ =�=BlN?,��ձf�g�߄$��	%_�Լ����e��R��V��	�"���w�G���4~�n�1G����b��N��Q'��(P�O�%B�o}q?���4i�ښ���^ɀ${������{�y��͇_��o��\'��Gm�nSn荵�n[�v�2V7<΃�ޝ�I4p}u��VI"׃�7��$���� ޻�-���5Mw��ou�~��M����ޒ|\ܰ(��f<Q�׭�?�����m�K^��=�� _M�} �\kn��f�g�>�1i������
���~�t�B��g�'��I�R�8����[�� =�w{�6#��y�@���mêY�7VYd�;�蟇����d����u>�B~$�r���4{L�9�*��qj���>�C�=�ܒ���}]���G��n��$q��{u�u�[K�-�.@-�;��� 	��%F w��u�����.�:�rfK�u�����V�t�����E>ӗs.�7e��%�.�!������〆�՛��uf�SK�[���bv�{��J�t�N�ުuwU�l�I4X;�ܪu]d��K��8]�:��3�� ���mX��:fX�R����-��F���n�(��ҴWr���o]�Nh��׀���s�+��v�^�
��5}	ܙ�)��ԯ/��`���or�ڵ�<�ƛ\��)��p
j�˻$�"�7/%��tU��D�Z�tR��IR�<� �G������4�#�!����p˓!��>��N^jyE�#�kD�4PJ��i��[C/c�#&]N�M*&��//;�d=ټZ�&:�N}Yb�\k'f�&�cM�<(*�|^	R�7X����]]�n!غ>.`ȭ
�q�L�܊e�c*�v��'��^ɡU�
�TbA�t��g}u��ݏM*��r�n�2����8�9�Xkpda�����K��=��#r.��R�g�u2�W�v�}���_%����h�k��Ȏ��m,O��z&���֪����o]�`�A�ضV�k�Ol�w���R�#�Z�[�]�JɊ��KWR�����=6"�^�,��y�Xɐ�Ɏr����5n�h8��;�K��Г��W���yy[yQ��X^��2k�>�.鿬@s�����I���ȭI{(�fl}�9}:�&�]==\BH.Y�r��&Xc�[�k�
�qn(
�'^�9 �dj�j��~���
6�r��zZ�:	Z��DT�˗� ��$���r9��l��nv��7}�{ݢ�(�(��B.H�2�;:��f�ԑz6�Z�v�vQ,����fK8���l�G'r�[Z�����SZ4�;�Μ8��A^gy�t�셝n���� 	��d�䑝��vֻ��Üt^U�ga�sX�X��0�h8�����vY8rvVL��G(�ӽ����#���EgeY@��t���fr�Ds�YE��6��y^D[X�Ȏ�҃��#�M�׆ۊӅ���#�D�خ)���p�n���r�ěZѳ�����<���������zq�n�ݺq�j��I�ݝ���ې;���G���U�r��p�^S�Y,v��6�*�h�l]q�kۭ���Ysշ'W2�
ϒ�\�,r\y���/�{g�v�C�x��y�� S�O���4%�0uͷr�N�
{����=��\���r0X6�{l��qr���;j�B%��75a#v2�k�vC��۸�b�-�;u���<���q��imd���m�-��u9S��ݺ��Ӎَ�[��� ^.��%�r����d�b^ۡ\Õ	�.ݵ۝W�m�jN�D��n�l�v;��6`�ɱb�}qM��v<ɜ�%ƪrGN��޺l:�ض���X��iY�i��6!0m�w2�~?;�n���ǳ]v�,��θ<'���9�<�7�<$���	q��];v�=cK����v�׷;h�"S;u��������p��v���#vq�x��\bZ�݇p���8���s]�ܮz{y�6.zǓAp�qtY�K�ɇ�t��Ͱ9x{�����gѵۖ��Ѧ�3�Z���ѣC�r�G=Eȝ͝����ƻN�zƩ`�]�.�&��G�uc�:t�no=s����&ގ;�Ր�v��^w�J���ݰ�7&m��z[��v[t�pZ]���k�{V�̱s�����n�M�p��^�i��q��k��������zn�5m��J� 83:wm��\��B��X涞:�b�ʦ�x鸪n����v�h(�FS��n�����S�R]��WQ���O�k��k�����t�M����ƻX����� i׶т�t�ܰ'C{<c��m�K�:M>�&�Ơܐp�Cs�٧e�(:jM/�9ӌ�J�+3ћ�&�ڛ��<Gk=j�u�s:ۧ�&�v�ٍձ��ݩ���v�6�����4q�\��W m�[^p&��v��܁�Y��<B�c�n�U8�[�'�]�#X��r]��'m����pqCs��n\c�뫌���"t�Mۮ����\���h��n�SACuN
wN�@5cqKD�6m��Ku�ns��_]G�����.p�;���u��nՁ��"냛��i5����훣�M;\��7n�����or;O��:;vz�����(��u(q�L���Z$B�$�d��X��z4Z�15��XsM��=�����ݛx��n1��֥9ϔ�h��S���3���Ǉ�ks��2������q��x�n��u�Atf�sDȚ���W8�-�I��@�]k!�l�l���W���[���K��G\�����ͺ�i���.���� /���D�$�U�s��;��.�z/d{����[�-�9,@�rzσ���%�`�=��_�͎�Mx�G��>��k>�y�l�_}	��s^���M���'��]�.|i��Z��g�[}�������6w���x���f}C���HaQe�,x�������3��vMN{�W{�f� ��w&$�I��ޒ⋺y�װ5D��6=��Q�87)	H���x��	o���͑I7�K���(���]�$}��E ��s��Jl�Sno/�i��_gھ���.`��+i�ڎ���/[qln�jw`���>�|X��1>}�qA	�����瑞7��?h����?~%�o����U;
�������27XA�M���/��=b�"�$��'��_��u"T���@̓g]C�=e�Y�X6�u>��v����t=�t��Âc��z��sr�]����k2#f�]%�VI`'��=өX�$�S��� )����I'���.���R�pߵ�
�վB��B��FGO	'�^�y�@$��;�m�޼Y����MN��7� \��I�>�v�Y ��>���ϵ�>����\���g:xI �Nv�ITI��&�}��ssܠ�}w��F�w��P�-7��TYe�#~�{���� �=�F��&���}�h�Y����v�����I$_��h���׵�{@�	���j�.N+Y��MѮIw����]'v��m��F�z@??�87F��(l�g�w2�y�sٴ� �=�F����yj����og��F�\s��J����@ϯ�v��a$��$�;b>i���9�����n�I%�<��Е�o$ǌ�Sޢ�߻|"TPu6�as;���7��f�$�J�x/5�3�������3�%��1}Q]97.e]�oa��srP�Cv���y��4;���d�*�1wȓԛ�;ֶ���-u��I%�oM� >���ZyվB��B�6�#&F=^�S�d�W��ʄ� !IǷ�$��w�n�*��������w ���� 9w�Krg��w�ϴ ����Ux5��?A|O���$�@*>���h��g��{x��m%n[o.]�-��%�;n�ch�zM�O�����W%�s��v���+�-���~
;-�u���{�� �*3�4bI$��{h�������co7��"t�3�k�8uG%�C��Oh��=�`N{'n�3k` N�s& �Gy���1�ٚ�=!���޻��S�x����j����G��%@$O�TѴ�A+~�u]x���{_��	O�e�;��`�����D�Xr������8{^髝��4O�aВ$�_�h	/�_oy��J�)�����
/r}�y��ֻ����-�����Z���iWf�6�m(y���Fv����_p8�6Wd� �S�i��}�Ҧ�ۻ����9��kn�����&�d��D�%﷜����]�M�p ssٟA���=������;�kvyF��B/)�]`�|u�(�a��핫��6J;9jc��n��j��||�������G�����7��bY �w��k�����Z�0>��DM�T�vh�F���6.��$�$�2�֎D��P߽��%�I(���BK��7��	 ��ڮ�EK���{��
�A@p�K"�뼞�� o7�yʄ�$��1�~�G�M��Nc$�"n�t7� ��緽���NO���-A����k��Kgh�M�����-�;��IF{�y^Z̨'���Wr�d��N�H�*e�'��u����@ ��޳�6?�55cz�s��ޒ|H�c��G3��ʹײۋf���t*�P��qT�]�[�H/l��6=kVɈ20;y��í�˾7��):���V�b$�-8t��\MÉ���X7�x1�˶�kW2���(Z[GV��GL���������[�=��n7�[�k��cl�=Ԛ�Cr�n&�Xu��f˳��v��8r�R��r�1�u��׋���j	���9�Z��7�X���������� ��ʀ�wK�݅�sgZ�p�m�޵㎰=c���a���m��L���^Ӻ��F�j�^˳��wϟ=ne��D�7['z�H�]���n7������Ü�}
�,
���̙�!$�o9P�I&����J���3��^�޹ ��{{���9$������[�&�C�α��ڗ�$�T���	$�
��n�E%j�nwOM�W���֓X�~U-�c{����>��:D� �����q��$���I G�o3�֙ s��%�CF|6��7��"�~'�{�}	��Nz,tI$����#	ت2�Z'ğ���7����'�ӎ�S�F�{��h���wE
����9�ed�I*� �po�h�H�o�٥�l�Sx�5�<����Y�D|ts�v�<�äCu�M6��<�Uv�J�j���.���H��2���{�ڨMh��4I �<���~H	Q�;��q���BM0w�h��"h�31���3Yټ�d>�y�=<���i��Zk�%�d%����Y�ŔxfXm���>�M#w��.�{@-l�P�k��Mb���廨�,!�����{(bԵ��$�'�ѦI�$���ݖV�s]��˿s�A��$��'~��(�����IMu��_$K�{ύ���6$n(o�˵q�"�|�n�I�3S r�ffS��{zҾ��Q�z,�@�<���&��9�H[�oi�Ύ�yj��B��sO��P�q�H������I&-�9�T�z����pp��k�ԒK�6W�iP����wx����;�#a�Qj�H��B��r�/�6ݍZ�]�W1�>���bj���r���w��,P�ڞښ����ggs �w�w3i*�3cGe9�ZC<�w�E$�^�T��/
�vj�0�]�Oޓ�O��|Cǆ��/d��\ɩ�I�_��$c��HI��e�z�����S%_��/�k���3kۛр3��o��|�)ypo4IgFϲ�_�~�.Pt��G��l�N���j=Yx9J!t�R�BT��ՠ�h@��y� ���Ij��V���7G|W^4|I=�|݌o=��{܏��lQ;�,�g�糙܎��ɠ��sز �	s=��r�$�Y���������Q'���Y?{�����n��iй�;O�<��)���{�"���/�πk��I(�D�Y�ք�n��`����k��{v���w<l����\M�2iǬ�2�ά���hҔ���F�D��O��8ߦ�'�_�{���^�]���L���뙐g�%�w����_��C�'b���������}�|\��WA#�_Ě�zn��$�h�o��d=g�G�/t�y2��.��RY6d��7b����W��o{�}�k>�� �����3ׄ[��50A$2ON�I|�B��ڗ�^K�R�[aJ܆`kۛ�k�=�m{W|�^�{�	�7#�В	%ӫ�n���Y�{��*�;�|&Z��#%U�R�&<�|X8i���k��i,���e��ӽ��z��zz�z�^˗����EH�!>'�%m�wpInp�$DQ;�,�g�糙� �������3�z-���Ě]'I>$�&���3M��}��g�[d��D�3����;Dln1,�u�|(p��
ZN��֫MGmM?g[��B*v�Vߑ�w���$I�y��I �E��'z�ԗ���W^?wpI�B��3B�)I
�t�j&j~�%�4�������l H���` o������v��[c}"J��b�uE}j��+=1�D���h�A$n^P,��v}�s��+��1`π7�~̡�7C���ڡύ�7�J]�#�N� U��w̟�4I��v�$��sr`�V/;@��M^}�X��EIe�R��ox��4J�w6=�9��̀m�;�y� ���J&uu\�Wc��`���_��G�}ԕ#�e�U��z��<��1kw�n[c��T2/f5l��K�85���z�u�}�!A^�"Ϡ�*�����g��k����O�):�-���ط�o=���vY�q�n���4�3��[/7]$饂z�01���#�%�m�x]���Q����r+�\瞻<��*e܇ݴp�k��fxlԀ�n���ѧ>;k8Bm�`V�cR���T����:�.����z{Z^	��`��&�����<l���Fu��`�-�&�Nys����77<[v1��#�{��D�P�Ɨ�ݍ���lh~��?3�DE�Ie����f` w���)�I%��N�	kb�L��HK���IK��7XMtL��F�����������$rԲ��պعu2I?w�y���IS��!$��e��f��;�3��"���
GaӞ̠�绛[�A,\�,��<��$�7L�u� i�{���ݚ���Xt���{���V���[��$�r�@�I��'q<H!s�U��7���ۀ��3���9�}!R����=�`r_$�H_��#K���z�+CM%��=�	$����� �<�@Ú��˗�k[�p[~D[�v�J���C�!�����NUZ���,�m�m�42�Zo��w�*B�(��א{�S7��{�Ka�&�#;���^����u�=Ǝ�t�w��c{^��8H8�w�,�b=����
�] ��,oK�)�Ό2Mk�ҴԷ�Xκ��%b6Ɍ�v7��/e���&�#�sP�j���F�,Vm)Ԝ�j-�h��n ��$5�N�	$�B������j�q�s-T��vE4S�6oS{-��k��dl{�k0 @����^�ǽU�w�>ų�wpI|��<�q/��X�UH�5GQ9��jo:���0�-ｽȔ����'@Hƻ�s��pE]��E�6G��=��h�.�m��h�bEy��}H�O�����Ý^�+p�<�T�}=�ܢ@;ڝ"	$���a�Ɗ�����t�T�V�rϜg�U���wF�y�k&9	����QH��$?a߻�~�;]�ۋ5��|9�Jϣ��)%w��$�ZG���.j�,�wI(�D��N���s�rB�(���H=���+~ޗ��]U�*U��l�$�i��I�g����n��}y�]������q�8�w�yx�:��I N/ΞI=UO���Q>^��:*W`7��H���ջ%cĥ�)�7��\�W}��50:�o5��.��kS�k��R¢>�X���\:sA��6���N�a�!�U�/���%��ʣDT2�\�s�|�h�?k���lp�up�e����+x4u·��`�݇���4+�oe�F�k�]�Rm��u��vp��;uܖJ�:�.7n��)��U�E%.��:��LS��N��Ϊ�u�nB�V�\݆R�0X�y<51��MR="�1f]��;==-�Tvr����j�gb���X�&���_��K��:L�:��|�Y���Va@�I�dQ!]�a�b�x�Pz0��\��!5�Z���ɼ!�=�yK]�Ki;C�X��X7�P�/a㝊��e$j>���;��a��̲�bĻ�a\C.�KS�ݼ�����Q�Pc�(����X�C�tO��X�y�Q���Λ��1���&�G��%7&��N5d���񎾙��]�7���z�C������nPmi�<v��Lm�w�TjP'�ͽy�e����Se��+ջˋi��ա%W̇��Ժ�l*�q�n�k�G]¡4��#&���[��S������	K�f#����`���U4��uZ��-Tp�9���F��v��Yz���'��
�h��՟(a�#6�}��j��[��H%\
�]��aܗ�c������WE�$��8�+���_��>c��t���t��Ҿ]�np�5\\*Y�G$�v��b�6} ��X�"�r�'������| 9$i���EŞ^GxYAmnˤ�Ћ3���$\e�u�28�Gf�yyG{l���)h�vZu�]���^�{�z���cmu�Ʋy�{#���`Y;k(�i�f���J����3���HV��;ʲ�A��h��k+9���vGem��:��gy�'^�u�ee���mcj�*γ[w���;N��<豱m��ٲמ����Ӱ�++;6{�yy�F"wl�۶��F��{Ǜa�k[kU��7�Y^t�&�m��t�n�:)/mf��RH����l�e4̳�^�r]��̂v�Zy��ԃl�-�v�ݵ���ͩ�l���z"�כۙ�6��ړ�3���kYd�q��n24FF���]��)$���Z���{X�w5���LB��jǟ鳹>B��X�K�<�DƳsm �*u�v�I~�t�57�0�������� wf����ze^�A���޻��x�D���!�C #�a���I���vA$��������9��7�7���x��$ź�[:ۮNۣ���#v��g�Rݤة�#E������T۵�����|���N�Y�s����o�b��ק0o�2{2Z^���hu�3�Oތ}Skp߼3�]iZR��h�k�"�$�i{}�(�?zc}���9��������EQ���7`'ϻ���~$�Y�Vѿc-�����b��w���ڛ��A�D��WW�By�{�~�jx0B>4�����D��I�L{�Q ���<G�G���qbO"���j�t�Ru�C���F�z�Ul{�*�C�;C�p/kR�ÕP�nٕM�ܻ߷�Xuz6� _rw1@���C�N!U\�c�{��w��@ ׻7��9v{�J�ͅ|I���e�$�}�nPH�{�ۿR�e�*-�N[Y�(Z�~�u�78+=�H*ӽ�c`B�L�������m)�D9������uz�#�G������ ]��{�	$�ޮſ%�P;l�l>��k7;�x��������*m���D�ߋ��`�ޢ��]�2�k���,������� $g�7������fz�k[������(:��}��ql ���( ^�u������;� %������	 g�o1PV/rq�$�[^�[�WK�}�Ur�����I%�5ϡ4I�K����5ߚ9u�׽�����@K��{o���R}��n�<��~��	$����6�i�<�/Vs�!���$�Gd���I.{^��[�E��cH�BtR����Y�o�����r��u���R�WH��Y�>��7���5���[k�-�f��8���ž��i��׹�COY�rH�r�s�חc��۴��{/X�B�<^���Sn�^���ݐ)�f�]��Y����3SvL�5΁��i�y3�/:�����.];]��X��vs�Wg�s=�o�ձ��t8��qd7ZN��rd�Xd���7X8�{m�G���\\���s��i�Qz�;K��۶��3�r�=e�����Ͱ�lv�j��Ӗ^ɪ�I#���;��;d�>ֳ�㍕K�EE�_V5c���^o��1q
�嫯�#׽����=ٽd e�oڴ%ٮ�o;�u��y��� �g=7�擮G�dD���w��K OG�ǅy���j���$�%�" j�.�	<_���gx��ڵ>$����u7
|���� �N���	s>���rw�c|K��[�Wn�H���ي���rtE*�i��o�$����^�n|̙���A�d��$���w]�\LU�z$�]�Ov�Bz�wg^VP˶���v'�{�	bQzs{̒���]����d�bPg�/g���h����yun}�����+N1�s��!�w�����l�����-�j�x�����R}��n���vs3� >k���I5��t�d��k)$��Z�N%}� >9�Of@���f��8�UrՍ�g�t` 2�L�D�y~��0��ne`2���q.\�\FKz�är����ÝM�6;.�>�7I�9/rfNM��ve����b�]T���CS��P�Nm.�^�I$��9� y�wH��/e)��z��Mo�=����]��ǆ �9=�!�7w��7� 6B���w�j�>�mo� �
g�n�H���I��$��y,�"����d�����ޮ~o���A��s>Y�@_{����=��r9=�-�\����ٙ��j����yXH���9�}	�MQ/}q;'�l>�h�T.���{9�D�u{�$$�$�z���a�Nץ�龇DGl��E.�+��:�RZ{��(��7f6�=��� �:7������!Yj��9�377� o^�3u�$��3�qNkQ�vn��tf���,�{;��hj�8��W�-��<kx���IQ}w���ջ��I��o�t$�"�O�A�\d�X�fߛ�j5@��B��j��s��}��o�ޫω
�;P>¶�z�u����%�V()�#Ү��l\'�F���Pz���W���;�"�8*��]!q���gc��f��Ҽ)fflG��$��>�%��ލ�uPC/��n��2�~�]�]b�eL���4M�{̀ I�N��I%�״T�^g@WRLCh��������v�]�o ����$�J�t��ǾOBUݵMz,^�O���%Q$�F��ȃ�$���Yz��j��s��Q��muA�"�:5��Ƀ�\�k��Wh�d�֣A*B����}��$P~����} A��M�n�ГY-ƻ�E�Og���A$;tbKQf�Td�e��l������c���&r���{{�$�D��� 萵׳i�K��P_�;׳�u秂H{)f�#R��mǟ#���Š���Y�A�~�V��e���h/�<���﹘���k��́�i٦O��9j����B0�W?_���5D�ED�I[��]Q ��D��	��9���<�t\�ʣ0��}9W�N5e
d����&qu]�]!Sk�_U1�K�w��X�MYV79~U�H�����Z�V��ܬ�Wj�o~�р���ml��*M��̈́�-׷�$9Ҧ"I�5���z�o͑�>����#�uEAԪ�!;jhP��0VH�hR����!�����FvzWG߻�z�T,���{�o��@��vw2�ĒMr�l��kS�b�i�<���#[��b���m�r�<ϏG:H@�B5�yw�·�\J|��M���_Ā{_�@'����{ѢS�9�Rd��l�g��7�9��sk`�ʏw`ڞ���6#y��Ϡ���Q>�\�&��^P/1���_w���,>��rY�Ys���{ X�s�%��Np���շ�C�Q��Z��ǯ����@|���>�����f<�$�����	/�Q������&��x]`��9W��D�����/5d�x�,y*n��8}���ʍjX��oub�ݹcz��,ݼ�wK�r�ر�����2a]z�����F����۬��wn�gs�\�0�&G�k��M���:�7��윖;^�6������nl����/�ʆ�o.����s�;�8qyj9q�O7t����5�cv�[��۶��+���{&G8��8�cs�9\�۱��:��pr{���<�ft�yvA7=�ѶzD��n'��cMm4k�:�v���Թ��9������Φn��ƅ=r�v�]]v燹7��X�z9]�❌�wW��p#�@�T��؋�w:�"I~��D�@j��z��7/�v��5N/s�����ϧ;�UB��)[�5��̠N+노{��Y s��s6 p���Z(%�{\M#s�ױ�d�EiơUs瘌�o�ǰ�w��6j=�RB
�ډ���q<@)��tZ_fQ�p�$�nS05���z��p�����_l s'�����)/��2��|�s��{�rn�H�A��a���� ۷�Nį,7�9��߹�̀�=��1 o����|�|�����$M�c���*S�8�� ��=���=��T� �Zݲ9�4�� ~���m�n���0�u�� s��jԲf^�%�^��ؑ&j�7�i|���'c�Z����h��K\��4��+
�ʮ���U��d%�p�5���Ӫ�"F�x�m�7�m��J|�h�*�PG9H��Ԓ�<�+���VE7-0�6�>lx�k�s�I���u��H������=^G�Ɇ{����ﲊ�l���Z=��Fσ���%�� {��eu�{��{@ý��x�s�ِ1z����eUߞg������}�T|a�v	A*jnQВ	!�2�4I��wIw�����nIs�TI���fSX���l,����X���bI}�O�M�C�z�my$*Wn�:�Nm�Y ��t��h�>�y�N��U݋U8�'X!�;D!�\QF��A��nv���;`�ݍ���E)7��N�(�/�Kx����G� L�:v {��BUU,�7��y*����s�<KU=:�HE��o��g�@���k��,��BIm"~$۹�Y'�L����Q ?g����;��n�&����"(]�v5h	l���$��&�"PK$�=�/A���tv��@ن��""���.�kd��u�mP(D���S3���0�ޒ͉Hk� u���p��0F�fz�?O��̀�3��h��{2V�#�JV��{�w^�Z~ֻ)�.zS�;7�Z��Ԓ~������{=0��b��������)-��7Q���!X�Dn��w�h'��M������m���۠o��0(f�E��;�3m���s�/EJ�lQ0u�4N�H���]�W����&8�㎼�^@�[����_g�N��ҵhx���~�	���#���m�r�)�iUz��x�O<��K�=��>u֑�6s�8sh�{�RR����8}�%�_y�ߏ�~�tA�'�(r�g�Փ=��w�qeЪ
�+�����'<�`�Akº�	(���q�)zo�$��	<�,�_���F�]�S�^�6�t��G��L
)K�UP���^�v%���s��2����4Yma�l�'��:����b��{~�������+�[[c�n�G��nWd��2�"[�spϽH:�x��+�.�GN�޾��B��������A~��oUg�fk�P�AU��� |���P���а҇m�x-[�����KJ��R�h�,N(+l�H�=�;n��q<統t�~������.D�S��U�\��/@|�� �*v�6/�g���S:���I�w16׳�4�o��rYd��8p�����p}]%n�zr� 7�ؤ'�ܝ 26~Q�F��������,�������u���=���������}[����߷At1q]Ъ�Tj����Z�%�%�9��z�L�=���I�q�w%����!Ԭ�D�Gg���Z7B�n��=�h ��y�%�����@�I���v��C�U$G*�iO�5[�Z9P"ר�WcvL0�h��Ӻ�xi�Q��
|��"�h�.�;�����ְ��t�7b���w9�ϔ��E:�<�_Jj�YS�r]&Ej��Ub�2y]p��#��� x��p�k��S��휻�H���v��Ŋ�9/��X�4��;�O7&E;q2���R��P3������j�0l)�P_+��q����*Ih�-F����VXߤ��x҂)��f����&C��7"�U��S��Nh��u�5';B��&d��q�{��u��"/X6��]�V���lu�@*}��c�v�e�1��b���C�:��,�ۈw^S	��:�u�EV������I�X��1�<��ν�һw�E(���uԅ���+2���,R�r+[{6�L�`x62�n�$5{���U��dAu���>�y7jm{�q��2=���;yYwE�7s�W�X�T�$�}�m��E�ԡ�*sd.�H�b���Ř��$�J��b��طڬw;*	/��U�w��X�n��kfB�)�A�Y�Q��O)ptN�qf���w��u�*�Z�q�qr�}ͬ�.�B0�����]fȰ�a��`gP�����M��Q;�Pwnm�P2r�57NLU�q�5�������ّ_(���BC|�mu�5t[Ҕ����^f��.U�������b����}-]>ɌI|�_NԬ�znۏ���d�Md5�U�W[o���O*��ɏ2�gw]+��������e��i�լ��T.��p3um5���vH��5�*��8�� � �m��>�~e�m�-��Z-�6n�9ȭ�֎��8;�l�!�Nٲ۱�-��t��{͡��^Y���=�<ó m������98��C�4{׏J��V{ְ���w����؇^�t5�3���s�,gN۰V���7-�o^����mv��Ķ�9�ցM��Z�Q-���8�H%��$m�e��N��Ͷ֎�nr�؂l�n76���ۖ�i6�$D���0��[�۴�vd�j�ְ"��tY����[b^{�۬�n���H�ՌÅ�[kd���8�0�r�m���vl6���H���%�[4�Q�[�c��ٮ۱m�"�l�m��&��9�)��m�)���[s�I��m8m�r�gl�vk#L�����@N�B���؅H����n�/[uv�Զwp�`Ո�Ո�de^�pۘ�x����#��g:���L��6���)�6y�uα�ڄϭ�ݸ��h��C,�=�N�n���Aغ��Z��ٹ��m���
�������uf�m��Ӄ��G��m�4���t7d78ݮ+f�Sk@{
��9K�;���gn�J��U�<�D����;�<�cm���5����N��Vd�WGH\v����C�[���q�L�Z�]vϽ�vNq�8�'P����m��\���˰�/iʜ�re�P���W]v3�TI��N�V�Gk�A�g�δvQ7]������nت��J���5���R�83���t�y3�l��]&s	�a֙�:wWv۶�7)�q���N9���W�#���v��wW���8�<ǫ\w!v�p�x���v�oj�5�x�vzl�v�ld��s۷ݭ���gc�d�5;��7<r�[�'n-�y�\�\A���,XǠ�\�^��^����܄��݈�0x�<�^t<�֬'���ɬ��	2׵�ø���ݗ\:G��;^A:{w�;-�9kuˎ�K�A焥��/i�V{&�wx��V��N9�^����[�+U��nm��';-a�>ّ�<s�v����G"�`J��r�-&ix��n�Oc,6�Nn�����3�[s� Q���"���1q���������r7b>�����n��g�{n����K�7�ni5��!�X�`�"�Nmʡmn��l<���,��]Zv%s�=�0K�;g�8�ţ]�Ý,�m��\�d�2��:4��c������96\�=+��[b�ҝGx���![q<���v�J�X<\۝�R`�`��9���6;:1p�x�7n0M���b���i�@K�b��N�6m\�0Ց��n��c��7�탂}�y��������w�l<8�.�N'��]Wc��ۃ�:w�pk	)�	�rp@�g�x(����W+4�U��ޣ<�.-�]��'���"�c�`����F�줞�mhVS��Q�,[Na�l�g�)�F m�C/'��ח`�s�Pۋ����ź�<��Y3�C��6�s�s��/.�N�3��m��iy�ཛzO��͠��{G8����^6ˮԇ`qv��b;v�G;=pcmgYRH����<�؞�۴���֎l]���:�m�u����B덞�#�v4z�t>���wON�������߾����L5Y>7圳�O�H�h$Gi��)6��u��K�S滿sس���q�T��՘E6����lm��{����@^���ĀO��tj[�og�����%�ϫ����4���ϋ�wf�O��4H3�j>�~����z,�G��7~o����;��ڞ^8�Y�˘��g�K��]�܃�
��͊ ��]0�����u��צ�T��t��
�]]Фj���z4���s����1����ot�O��F�_�j]:]@�{�lP�X�h�{n�Rk��$'��
��xغ�/H�+Ym�F�v��<V����[Z��5���ڟi�v��{��+Ͷ*v��Ծ�:� ���E��
�)hOKQh'7��NT�(8�tM�Q�r��T���p��'-Ĵ;�_�
.�J��CgC����k�M�Ah�L��\M��Е��4�H>o�4�Ag}�Ri�j�Ox{g"�>�j�6/�ל�t>�z�`�la�:���޻Y��OyǺ	 ���k/����$��yU�����n�Q��� �����z7����_W������LxԘ.ȱ��8�"�@	;ܼ�[/|�>�3q���A�~��y��n�a���ѥ,�텅�Ң�,��ݕyq\���g/\`�X��tn��%㚺�w���/l5���o@f[	#}�����Ǎv]�u�����V<���%h���՘�^sۤ��_E�{�ӝSl�(Ľ=���x�V	���ۤ��/q�mz���@�ȩ��B�4��gw�~$��F�@+������y	k��� Y��K]�X��3��<;�n���K��R*�t���P�.嬭�e�Cv�����r"������knhY���.���I��@�w6{t��d�Q��#4{w��=�:����m2NyY ��H�I�'�{����F�đ�����uV.��#.�r���Ӣ�]yt�1Z�|(���3��'�q�*����ƅ�����D+��{^2�s�Cv�e����k`����\E�@�<��Q��W�vg��I��{��@��{�w���k=�xH]��#���,�+ﰐ5T9o�=��6�G�����w)��H���8�I8��S�^��i�yWڞ��+�+�f|�~��`'�ǚA/W��Nk�`T�z�@&d��$<��'D"�+$UQһG>"�"��r�΀�[� ����l
w����Ygˉ�5�&G��L�M��]Nlw�8��ٙ��d��s�%_�~�)���n�M/>}���5��6��WO��zm��Mo��~'e��5	TA��B����l {V}�=�]sY��Z�O�W����y���Oe�+&���jL_��|��tW0�s�Ta"D
����B8&WmmR������IT�F2����[�'�ژ��+��w*[<�(<�]�$O?v�$Yhh=t��{��������7:������7~ H��4D�W�k�st��U��lP�}�TUؤ�����[�o�}�>-S���5Z�}�	$z9۠�~�ʿ��15��`���_BE'���μw���T� ���~$l���i���k��J0HWz�ϛ����[RF�G����6����g�̭o��׉ku@B��,O�f��MC<���w�dկ>��ѬWРq�b����"�;���"
H�E�8oz[[/6��E9��6��+,U�M��&���U=Y����l�ϯ�n��]��R�t�/c��{�lt7l/mzٲ�7z�M�,����n�i���Nֹ�6ю�*����L��{g��'�7���؇b�ca��8�zлz�p��.�A�]u۬����a��٤��j�aǟi��c�;*���^�s����k�BcGX�k�|���3ñ��F]��nJSV�q���Bs�C�b��p�j��:�4sX�������z����㮋��H�j�fokq��a��Nh�^)R��#{w��?Dyb�ē����:2Ǣ�����G�H!�NT>�IT�(�����׵�&�}�mU<�>��1�$�9�Y ����o��c�Br�q���:�|��6�`5~r���� ��uN����y<���Xѩ��o�cm�9[60l/���
;W	j� vߏs����p~k�ʫhW7�ء^��~QL����}0���f��ōU��Y�;������q��~�z�����I��I��t����~Y��z���ϙ-BuV�m��q�E�9�tӚ��;g[�* �j}S�G����H���E�`����H�&�ᶦJ�;�<۞v	#=����(����F��۽��@6=�_�߄�7�[�3m8�})��F=����p�Ff�FH4J��!�t��7�����V�v�
�Q{�a������9R�3������I��&�$���w�_
�vG���I*�D�E�i?[�ō���w�X���~0�eBA/�^��yɺ��i<6��Z]bM_g�~�p�9�ir6��r&(Oos`P��m���O)1Y����M��5�&�ߵ��=���m{��EX9.g������'���$��,�������k�=��\�T7�u�b�nϟ'gnm=u��J�z(0�q�V}-��	�f�==SV��՘2����O��ǚ�VL'_b���U�uQv��;���o�t��<VE�E̰�W�̧�r�׳*5o;T$��=߈$ze�`�rvzn^�Н�Ⱥ�)*@ݛ$g�6c ���AOa�y�g=�\�'�wQݺ5uax�t�e��;����x�bܽ�������E�s^)Ȑ�f���'2�g7Y�?d}w��'��;F�H#�,V�T}�%ASpe�i��[\=���o�>=�>���� T��)�O6.�ǐDޓ�7A#�|��*�}�7�Eͫ�(6�ͩ�c��S W�&�(
�+�?o���J�g�������Ԩ��v�x����n#�t�ʛ���g���s�OMҹ�M<���	�����%3��,M���X��߻��=e�>��{������h)��"��f�����o���9:�wҞ�A��U�v�{tgv*Bt{�k^�śN�hL�i�c�ɯkwd�G�O�ݠ���e�U7�G���k���O�#n��42����懷!B��}�7 �Uɟ` �l�`|{z<7����ܐ��Q�l`��A��7mN�0
p�:i;K�m<���Y��Fl��o�׎���{,52�t��7��ÝY���jw�*6IPT�(�CoѶOo4ŋ�h6�ΐr��Y�o4�G����/�څ|Q�b˓v���[�rk�8$�=����kn��:C�0���>+2�����}e#��[�ꭷ��{)���N�j<���	t){s(�ڱ7=���95`��k��w����<���ë/�
 ��t�}�o6��5�s���s�I���= �ڕ��^c���t����I;$��f&e�u��O��N{��y��'D"� p�D�j�~�M�|kc���\�` 'o�`P+��4���U~ms���y�d�* �R�'^nk`��>�.��o9M�Y^�@dǻ����wI�'���n��9{{�V=���~y���o!��<n��`�n
]�U7rݤ�Lp�Z�����n�I���,]���,2��98����{���F��g�����%V�]�9�A���nw Hu��H�z��8;��ׄbv����x*�,<����=����s�I1���nַ\��]�^wd�8��z�n�����J�+�����]�X�G^�\9��˷X�/n�t��z���on�+��]�y1����x�'u�=N`�Y�9���b!ݞ�[�n"�����s�qV��m�ns����Oq���{e5�8tr+�k����7{pWv9�Duy�����_��[��U>2��F�OǛ�� �=��e��b!�r����$�<����edU�UѳGt�g_�@>��pȲs�� ����$D�]������c�%쪗�u25v�&�
r��}Z��� +|� �ǘ�K��<�� 6��H�]�)�D��I�x��T�6���C@/4��*�j���5�j^^[�5�{�۳��Ԥ�H]��/�b�/7�@�>�Gi��(o������'�łN����弮{qd�r�%�Ct�2���ؚ�3��oq�3����f�K,M�=�|�D4�}J�gso������;�t��V�>mR���(P����ҙ؜���E^�&{y��g�^}v&��Ei>��V[�<���P�%�)���E�
KVœ�g}#;.f��<&<�X]>��J�]g��huf��s�Sq{� k9� 5�kb��YF��₶��ʴ�����X�a���L����N�!�DhH}���$�xͱ@�7'��&f�PH�Yig/.��v�0XwFPG�� P��`|w���g�3�,g����}n��$��s�Θ�>��?��NRǍ;.e���С�8��(
�w6�xr�o�׬׭�X-%P��VJW\l�mk�f^)��ル�v���	�KQ�7߸��|�h�JWv|F{�}��&��${�n����1��+�5K�Q�y��!��2��W��?I�Ю�{���ʦ���-lP�w6�Pե���y�N��u�^���;�r:��~�����o��w���@ԝ^�r���R�X!��l�=��C�n;7{kS�yu3h![��j#��o.�q}�ou�9�#��&I}�ղ�r�u�����5?9yu�#9��ʤuuD=CXg�D0t�s��b���2RP�+�/m2�Jx����·V%�]#�rr#^I��M�ug-�_��6��ڤ��3A����n-ʵ]��!ٛi@ቫ��V���1�NP4��^q4U��ԼR)Y���gG}xէ���T�Q��w��5Mk�s�^��۬�|��8δOr|(X8�Wm>����9ԙSn�2�����gJ�r�N�}��:7��/�$��Hc�s���ϣ�u���]ԯe�h]Nk��q�y���66�+��v0s����F��C]f��9tYj�K�PzWi����9�*����S�7��˪C��PpJ�[�2S\�A�;U�L۽S\�3n��5&��i�Ҏhse��w��.��rit�^>.�9t��O68��]ݔ7�A%�..�/�cNͿ�k���|�
C�-��*i#r:��cZ[���mU�2h���\�N�p�-Zå��Cn�w�v�Z�J��v�v��]�x	��Sfh�\U��q��yiT��foW&y���T��l1tj�S��̉�j�U|c}\��&�V�^���.�wn��4m��
{1F�ZC75tac��Н�;v��h�f���3�obA��EL�ΙB�w%5�^�]�#̱$M[�-t�n�z�]oHe9ɣb:q���E��v ��j�l�.š�e��w�:ͬ�c�;V�m���l�8�lbLc��H^��'cm��m���٨�嚽�=�M���bvj9&aD��iy�=� �B&V��iq�`vV�Զ�"۬8���W��n��nӐٴ�Hgh��@��-�Qt�m���2,Ӷ��rr���Gm�̻H���:I�,��M������mi8m�(vs��m�$�OlDtC�
�8kIN��"N*s�
��7m�٥�q8)m�6�n@���8\���qG��Ʋ�:Clw�pG�n$�8�)H۬9.�L���HlݑӔ���4Q�%���@�������D8E�%��)/<8H��:n�Sl���m���g[9_.��;߾���ip3�B��]y�{W{�����&�{;t�@��w@$����;��T��`�E{Ϳ����$P������]��
�Oz$������٠bn6 o�ͰA ��كz���~���42�hث7}tl,��6箸���+V3'C�i�{v.��7j�P3A�IOQV��
��#�h�O��������銅���wt_�-�B��M���
 �Q����~�a#Q���C=�khf���i��O{�w@$��>�C�ީ��5	W�: �ת�RD�(f�7��F�A�s�3d,P�g���G���H0�v?�����n���Y�T��+{�[V���n>�$�>�}�j��<���3�����6h��ܴ�Sh�_NwR�׊#x��i��9�zƶ�V�j���\�fWml�!TM��ڎ�7��f�ݓ<O�V���6M]��EX&���J�N��K�|��wK����	�5�ݾ�}��~�������mG�r�[CO�z�n�P/t]��ۖ���������]{�d�n�z, J?kt�$ff�U�����4i?�N�d_ �����pؼ�׹��� ً"ٓ�t��eV_�h ��P�Nv��~#r	9��*���x��D�������J�\毧�f�8�o��4V�
��D�|���@*�3�w�XHc���Me�.�>P�#
�n�(�\�[ �G�I[�p���$���{|X8��,Q��d7{A�=�����}^���� cs���l
��m����ډ1;s������G|#wGZ�{"W|"̟ܠgN+�����m��t����!7a}��`r'b���&��E��خ-�2�ƝT��>tMQM�rf{U(ʾ^�R`�K��ۆ�n^�B1�ݑsɣ^��۲��H��3��nص�x�z��Ám��y��X��)\Ⱦ7[�'>N�U2�Fܷ;k�U�)ϩS���Gvq>&Al���_���dBQ��tMu�3�uփ��v�m��V�\�m��1�C��r���b������X�6{\VuU�KjN9�Z7���.�z��y������Z�;��P��|q�������*���u�ϵ�E:��m[ll���ښ��_��m�L!��Č�st_eR$!V-#j��z�;$�|�:�J�|����� g�M	����Iy���Yο@��|�u�O;da�8[��:`=��0(:���W�坙: 
Q��~���t�J�J�HJ�����nnxYOA&�o��8�t	���Ƚ���yk/*���AT�{��X�i7���$�� Ù�Wۥ�5Z��ލ����F�~"=����Y�\�wD�;��KT��,@��#a,ny�ɲ<Hk���w��rѫ	>�oߟS�uX�Q�
�&fz:t>�kN��*�����g��l)A�קn�OďI7F�`����nȳ�x�]�U���7�tv���y5=�o1AW�wƇ���9<=uy���v�c9}P�͕���p���`�$+B�`b��XG���y�sZ�������	'��M���{�	�,=��>�fm��~�jA�)��)-�_z���M��k}�f�"�,�oI��2rn���Oƻ_�!��Q'���������\�{fߦz�U�<��@k�*����=���7n�ߵ��=�����-|k^~�'�7�����nŲ[���@�f����{�u�r�9��AWUv�wZ�<y�Kt�n���N#<�K�<���<m���/z���A](nM����6f� �5�W�u||p[�v��7B�
��|����tE��Y�+^��gI*W��-���CX^&� -�UB����
O��M%���e3������`]B���@PoϝS U�
�Ls������;��mmwnʕM��2<�kM�Mc�ud�C�Ӥ׵vq����e�I�u�ϤtC�F���h���rx`$��}�t��E�Y"��^]/����~
��)� B�g� o��A �ޛ�t����=���A��}��ec�5y@�9i�Sϛ '��uC�k��;<;�RE���_:`{���َg{���r�kv�K~��~�V���]�K�Wuaq��Nu"� ��c�ڣ�������^^`�������|�{�t+�d�wn�<Nυ�#wc�$h�슪�"գe��sѠ��	��(-��O��~$�=�H>���A��no��G&����DݚB�RUv0��n���O�����演F��R5w�7�@z�͊w�Ͱ<��l��?fa��oخ3��nng�͞L
���ؠ8s����b����>p�|�)tWu�C�r�KY|��}X�uҡjị���s�����'�ņ�^�y�Iw�	�G�EW,ШU�ތey	x<���{3�׭�(���YmZ\��3 �x��})��:�Wb�;�y�I#���~'��g׾B�5cN���PH�׃`�|�s�����N&#ZX9�̛���N��F/�Bx���U��+��^��?�z�
 q��C]�S\���Ҽm�������O�>� Z+�������Y�^(!�ؠ+�'�[� ���( O�M�X������J�JѲ���w=�I>3f$*�x3iT�p�pGz=�$�f��y�D��J�**��2n{��>cԽ��r��@PCϭ|((��Gg)vm_�&�������5��^�� ��ӯgn�wn�z'�S)5��t�����b���٪h��d��x6�¨��*�ͻ:^�׭��U��N�-��8X��I��
��'4�^�˧Tr�ce�'/�ٶ᭳E�;���UW���t��)E�;f6;+��ӷX��I�<뵒q��Lݹ���ɹ��_V���*�]���5��7�`���.1�vӞ�����4uѩ���:C��n+�n�:�[s�����t��;!m̜�q��tc��u��ly{�=�ܞn���Q��n6��Gd�3�9B�v�mv�ω͋t���r�d1�����x�g��K�U�8��g�/Z�v7m� :���Ǝ��5���k�H�e�hT���w�Q2?Q��Nn����}�	��G�b�㶟׻��m5�s��Sm����SW[��w��_��GY�ŵO��O�c��Vy���8�+�m���<�x�̤O��P̼��VOy  �s]1@||�z��mc�H$���`�O^����*�!*DZ �v�f��XK(����(
�r`|=�sN�s���T����s�R�2��j��ӛ��o���7�j���V�b�zVI����m���ig�����߷V�L�	V��lP��ݻh�n��/;v�vD�l�1����x�j%}e>��{z�O�W��4�o�����F=�XW/G��e�	��{۠-�(����lZ����gͤ�u͗l��ߔ�c���=:��M�.�]$�h:��8ѷ^����3��?�i��h̠;h>�`g��-��'�VZS���X�;{��^"N�a�f�z4�F�	��=�9ffc�� �יW��u�vOo�H$���A�}¼�u�Oa���d�nOn�}�MѠ�Р�8�"�]�_OU��Q,����'h�	$y�n�?L��^����& >ݞ���l���dU-��k��G��S{*r�f��ٱӪ{�� }���a��7�RHdE`f�Ud!@Րj�]�"kvp��rݷ��3��/E��ud:n���������mR*�Wc�Ww`ߋrn�~2o��5�'�5��s`��^�sn����v�j����?;���v��NZ�k/��� ����L3}C~�+L^��s�[\� �d�
�Ť�}��7�~UX ����<��m�{�q��@�{�Sf�0��2�%�!)�j�TL;�N]ϐ���j���Tݼ*�&�����U}�޼�'jG�J 
�w���M�����j��3Ge�T�1��l�U���(n�YH[�'@P�U�Z���*7�g+%��/����������6��Ѕ�N�קy�W�i�s[���F-��} �w?/����|�J�=w&o��}6���*���ɘƹ;t�c��4\��C��o��F�l� ��-�7ӻ��7u^e��5����؍�[�qr?^��n������{��5HQ�*�O���cNmukk�%��R��
�*���#~���+�{���+UGw��(��/���⊀m����D�� �I��ݬ���~T��kَ�X��vj�̺_{=�֭OU�9@��<~HP6�:t{��箔2��<{�Np-��/އ�W�{���p�3��a��v�\t6���1V��D�Q%;;q۾S�0� �������R�C�'l��{��=ʺe��ﵧ|�O��*c����;Ա���w5���·*�S����{��~����ӛ֦��=�C�֙%q��+�s��d�-kv�{m�WoGn�jQGD��ߟ]�v�߼M��f
�<�� ssS�C�{��N���x��'��xT�e }Η��:�$D�C3۝�v ���^�~�����t �l
�>�ys�Cxx�Y��5�{la�?<V��DՃJ�X��٠���˕0>um��¹=��.o��u�{]��7�+�'KUG�S�z]s4il[�v��V�Iپ���G��n�AI��7ڼ��\ٜU`S�[`{1V��tl��^�>l
�S��/;��'_9��k�T6�9\���_��HH@��t���%����%�����%BB��$ I�B��BB��$ I���%�)!!K���HH@��)!!K�!!J$��	, I_�$$ I����%�BB��$ I����%��$�	,$ I��d�MdT���~�Ad����v@�����#��         P

  @ (      � (��  (�HP    �(��![5s��IJU
��PR� "R��R	 �( T�@���$� ��*�����b+3!�};����'�g�'��7�'g�t��(w�[jE������5^۳B���U�i�Yrb��iS�;������y=6���"C���UP*��=��:rv:˛3j����/��م5��t��S�$��e��Au���T
�V  =��]����|����� ��BB������ �*N�
&�fjU�i���(�x�P(�$
(q�9�GN�j�ݘ.�]�V�%�2��zݘ�nyE��ɶ< �&���>��Ȭ�M�ww�3�Ol���)s�A�D�Я^����Nǻp)*��=}�
TR�R���+l!�m=`KѢ��*3�;7�mN�z3��J�� 8�@�  �@Pr���g��h�7��kz��(Ǒyj�m�$|  ��U@)% (�*��.XT��ͽs�H�ԛ7�U�n��z�&�A����'1���A� י��jU���/{�rݱ^�t�����إ׽P�
ֽ`�β����_      ��@RT�L#	� �	� O�Ĕ�T�L d`  bi����H�%S�C hh CM�ت�0�H ��	� C 2a��ЙU*�` 	�� @��I����	�(��z���h�F�O����/�Y��Ϥ����&�y�����Ӽ�\��I<��j��  @��IdA@$'� H�d�q���  nH:�g�����:������0���I� �;wd�  z��0�d��H @�!���-�Y�dA?��~����߲@  w�$��qp3���X���}���Ӕ���~_��oP�K�޻�չ�����_���n���񁙼�pf#!��Oeشh90�]L=�gq�� %C�����h]Ȼ�j=�\��mq��41�T��H6��FP�dC4ҡ��,����vGJr.����n��3k��V�M6���^^����>�.���u��+s)z�����y��2��}���L�Q��M�n��w�B�-)��M泰=���&��D|�̎����dmn���n,Mo%�oӱ20&�����{r��4�Fm\a1���N$ǽR{���pXN"B/��	��1ۛ�R�6��b���ݏE��2xv�{�N�ی�[�lː;����8n�����z��W-8pdz�Ύ+pװ��(���dCm:r$\� xl|�OM��a�f����ծ���'�N�P�F�$D`�ӑQ����-[F��cՓUA��t.1&�J��[  &M!���.҆�D�&Y������[���V�g�aWvn\NW<8����m������j����˕ul�8Vٻ������.t�����I�]JI��b
��a�c]p�cU�n��9B�nN�1�p��:�x��{._%�y��+;2ފ ��9�ob4b�3��']�C�&u�C̘�#�fw,�E��bx�ӛ�� ]9D��7��K��� � r	���gq�LKxYrB�"�˄ ��g��޳pr׸�97���s{b#���/;���5S75�����G�!�ϛo�~}!6���DQ,�k�*����=���;.\-��/�M�<|�m�>�+ם��-m��9�d�7&��"z�t-�d߄+/�;�g��-����܇qbl�D��E�ڹij��ŵh�7��sk������9{sY�.��$�8��<*b�U��VQo/�B��8n��{u�={,��2J4��`��]#���^՜�ވ�U�c�I�ze5��,]s-]B��.,n�y��
�#�zs�/��+�\J�8OErN�{$��8L�����+7+R�81�X�&�ݛ�P�mS4�ڑ�9
&��ޝf����]�Ɩ���\f��fo^���As�"��ۇ2\� �v�λ��J#�,ӡ�ќkF�!e7�#w�b�3^�74��[Gf��3���x�U�c��a+U�PX��LMM�{��:lp�����t�-ά��2�Q4�����8Ɯ�>�7�)�2�&k���Qtb��I��X&��7u�Sj�d��ƵLx��K"����z�_��,����� h8A�m��h6n�BXN�@�:��n��*j���`޳�v7����\��݌���M��܈҆>c~0R���Oq�K7��Di�[��4�Ƕ����ӎ�{>\Mݜ��:�"('A�N,�=p �tzJHGy�N�5�tHtc�y���t"�͕�xw|d�.�#/yۉp�[�kvŪ>��>q��B{��4��5��/@�8�=����p\{acC
,�y+�{t6j�cy�׍5'aq�㨇nV'R�p���{�J֪�Q���J�扩���F�a��e�Kp�#'�q%Xl���F<*5��9�h�Bh���x{g��$l9�"�p���y;���]��z%e;oJ�E�Q]�b�ٸ>��d2�ӍW��i��ٻt��7ٱ��Ͳ8ݽ5T됥�),����u$lp|����4�>��)n�UJ���}!3��ն*��E
	�3�h|
�{��S�����d�]�Z����J�>Z�)�BfD�gM{��	��N����2&\cn֔��#��̮"h�>:��7���s�i1ճ5%�SdȗZ����U�[ڱMY:�O�#/
o�kД6�u���� ���^ �^�E�!�hL)�>�1��9��a�-�#M�.NVֱ�]�-�BV�0;I��D+;�n�{`���C�<3��7��|9�j}5��n=�х���x�w�s�Nz�3��ðe��Z�ޣ���M!�7E��5vs.��K���
?u�}ؖ��I�,8����b�0%�v�6��"+�,��Ƥ4T
驍j��:�s��ٍ'�8f��1��r��q� ;dm�ZsF�T��;�d3�E��G,�E3�!9δ�m<�;�7��"���sNU"�5���p��9� )=tR;�)�$�����it��7Nȷc7Z`X�� ���}�3\6��1�9on�ơ%�"�hNBq'rr}�oA�^��Vmһ	X�i������i[�m�Nr� �	�l2�Q�N�NL#����Β���{���8u�����@vv��]�&�����N.a���x4<G�� B|��m�4�D��<��]})�STo�n��(]��D��{�GF�/�1n%gX��y�y������h� %�{C}�b�Qٖ���ճ� ]�h�Jsw�R�]�N�f:ۺY4X�^|�Q�Q���R�ǎ�*�7.����(�9�N�ܝ�ov���f�e:M[.ڱa�wq��h�]FӸ��[�����>��j�kLB0���4b{��" R�Q�����6��5���r�
�;m�I�
���QAU�O>�8:qu��9����z�%�-gp���Q�Z͊��q��#��캻�T��_`�_!XKoM����Qr#�^6o�6oJu�SX�=�(����-��/�&�{&�xmx�J�\�ޢ	�D���O
"�2�$ntu\/�Cfpj3wu���z\�[�����[�n�P��`�͌���c�G9
rh�:.�n^�r雗	]�r׿�R����;{#٤FoG�����.�sͻ1P>��� m��"�ȸ���C�S|����;s{8v �O�P55��ΐ�0�ݢ��L��������8	�+��K�<ќs���,
-��t9s�t�*6��zܝ�<�2g]k~9�.��2��RB��1lh�xz��Q�%�Ecl����*�ۮ��+ު�)��`��N�����9�&������N�uq^g,�T=n��=���=@WF��'[��siwC�N��	ó��8��/J�qSk��nE�sE�ul؎���Γ��w�J.\�"��� D\c�;I�z��s켛�3��7:���~�5ݻ�iIt#z=K��U���r�FW2��@b��JA�	vn�\��5s�-�Sǁ����ˉ�;��8/v�{���Z�'A�sZ�r=����d�R)�m����}��0MC�)v��L�ɹҗDo�o=��~I#�ᗇ`�]{�*��Q#p7s��.������RF�xh�O-F��s}�����E��S�7W���a}�|����vL�~�M����m�Zh�ܧJ;8�v��ېl[Z0�}{u�Uxt�,UE�`��R�3lzHK�n���>��C]'�C��	��<������C2v�{�dѝ����-͓�͓�a��ʲ:�@��h&m�jTh˛wm��W|�X�X0�{ ��g����ں���s��`��(�s�����`� �v���������q�j��w`�������`�ֽ���q�F���&��JN.��3n��:�2���rpe�zf�iŅ��D�EI�-*2c����9�-��щv<�������/��C� W� �(ɑa7/y�k{8�����7Dn!�̬w��iZ���FjE�WOWVs�t�sfT`�C�A���f[w��$n��Ź��J��'p����q
SK���T���T��;9話�Q�I�]ݍH��@v���3�]S9��.vA�ƃ����M��g���y�f=����Ü�3�;f�8v�mg�YC��Y�� 9�9j�м���#��`3��7V0LP5��ܳ]B�q|�yIX�C65�Zf��1^>K���pQ��pF#�A�p��|���-Dj�� �whX5X��xpP�@��OȢk�~��%9�Fd�����><Q9�^��_��ofϰ��$ D P YE!��$�H,�"�"�$,���I?{
��� A@P�$*H,�I��E BT! � VB
Aa�, T��@ $�+! )	�I	%H�� ,  ���E 
�,�$$%d$Y	!"�!d$� � HV`IYR` (I�@Y$
�HV Aa , �d��g�����>>K��}_Q�Ϗ�??�	  @�N7�kp!>��B}�=��2��!� ?A��w7�>�快_7���g;9��7��*ks|7@g���. �<�dXh�ă*)�l�jDj�ͣ�A[=Ń2�m����{�⻅҇,}��<��������R�Qt���=/��ն��
P������[^��;<,.J9��<{���|w�9�A�|v��^�L����<�߷��_9��[�"�]5�,'�W~�h��9��yuj�?Y��!'v�#>g�F��b�@���[m�}����t$�p��,,b7��>�E�ǰӫ	Km���_y�.�I�\����n�D.<6�/,��ݚL<X���;�=��bv��`~0 Ż~�۹������CFS[s����j'�{&5�����g��>m9;ȫ�9,pD}��hr�<��r�X�y��wn�[�͝M��%�4�<1n�4���s��E�=�+5��c�L�%]�j������� �l8<��o��|3;�!
���ʈ-o���>3��w5��� Q��\,�K�:��~��Wܹ�x�%�O�΢��x�׫r����[�"���f�ݼ������ЖC@�K��+�Aӌ��VoQ~������>�6-WnNg������|L��p{�?AY_�^���<�e,�Fଝж�t/�
��b��ۍ��+���刍賏8�k����(�<�>x�M�г��zƞY��f�X0���v&���y�V0G��ܑ�λ�eXM���k��y ��K>�|�CtT/�d���^�����o�W3]����{َ`�'���v�|��.�z� ���t��7t{�t_m�gc�ݝ��u�Z��nnnk {d��]{���ځv��H��z��E�+b0U����}�j�N�Ƚ#���ÌPϼ��F6z��&�x�8��7Ƿ�~:�S�����<3��K���ٱ�Cs�N�"��p�-ta��K&tڹ�K^@�L0�[#�odGi�G:%�R޴�~�ӛ���{��W7�4"X���Xu��j����6���ZN"��l����B�^8����6&$���u9��;5��N'����ֵd׉=V�A���]�3!f�j�p�N��+3�{�
^�����AB��Ni����3�Kh��_o9������o��c�T�>>9�ju�����4��s�K�{ؽe��Y�����eA��fM�Fi�a��.��jr�u���u�o��'��S�����	-Ė<�6)�d�h� �&�(֓�	�A����������®y��ӸԒ�Q5��nI�q�ɵ���co��X1#�����~�sÏ�}=�{���C���z �xԞ�k�d�+Sdv��1:۳5�"��uF�_r��<6��d��ҙS�ah�~�M�j\ƌ�0�\�����䠛�z�V������&���L�#����g��U��y5t^k����E�f&���
�[I^>���ձ{'>�(G���U��Ztf��Y���p�f���8V+d��^��#��3�+U�zY�o�W��g0�rP.�8�mm`0���r+ca��ڐln�׿n[�^@_�~ɏr9���)țbl���<�����y����7�������E쾞���-XCgg�wEkA�˖Lj��<�Fx�VVF�����c%�,��,f�qk�=m�7{v���Jp�C]����`��и����uk �0ۋ[Z!>Շt�m^3K�ki$�a@�m���ʭ���oek�Iȿr�|���W�|������+��׋.�;��ܕ�7�BxJ�|���#93�Y2���9�����v���S�]<V����2�v?����gz����lX�'vi��A�cb.�2!M���eӘr+Nd��u�$�#3N�x�=~K����Ǟ+�L�T�Xg�9G�2Vo��k���v ,Fʝ��07���{�c�0 �M� ���#��@�e�W}fy��vC��潬�YT�uX��!ʑ�dkm�o%�(�6ל�MT�MN�c����&�xw����ۏ��Pw���w@I}�hxzՑK�o�P>�����,����qŗ+��a�f�P�B>;7�w����Ok=[�1��4p_-���;���Jw�g>�����^쏰n���;�蛋���=��/z�����N�x��� c�b�-)v��Ğ�r^�g;�d�]��_|͞�~�	�����{ժl	ӆf�3���|�e��Su�>�Z�2X|9�8�p�e� Y)�&��Sd�,ʽ����y[��"5�;g���8���{�秎�g��Rˍ�黮��f������i6V1�:k�\��MTeg�w,罺k�gC(�.�x�{�Ɇx����y^ua�o��(�b��@͌��8���n���[�+��p�d���G$!�{�hK�����^G����AE|���Ϥ)��g����`�3�:��[�^8OD��ķ(ʵ4/I�H�� E��A:�iE��sܴ���Nyw}C���.��J���s�%�7��,L{vuWO�8�~�&��h������~&�S�}s������Т����u�*���y�L��z_=���(�_����Y�˜c}�yx/��1:7/��[)��w�Νy�����]��:w��%��a1�q�6�cw�<��s|2N�;�f���]��fNdg��<s�7��,���֝��{�,���~8�}`HyM�����v�<#l�^����H����A����l�1*Kf��E�UY�}�׉�ܺM�̮p��vr!�z���顭�9FR�z���:�]=�9��޷9�sz+���^��;�O�懭C\�	��<���_e:uvS5<��fܸ6��[�e>96-�����Ӽ4d#0�t�8�;��G�;���ay?nǵ�,^p2�$3-��AȟI��ӽ��8��l�{��^=��Z7"�4����\�Z�NHШ8}��������'����8os䢞�֖V��� �d��Am�i���Ӻ@��>�%�榢@iuͭ��I�;�z�����o���X8y��q�~�h��<MmS��-�I�l����g��Mf�Y�L�}Vv5�1Ct��L*H���kq*�[�޻��^���.��L6v�4�ͫ���８�<�wX���/��	�r�����z}��D�i��# il}�ק�0���ێ�@b:q��V�K��Y��h�kܾ����*�63���'b)����;;z"����+1�U�
��c\�/]
;��i��=����0��9�@�^x���Y0zݎ���W���8�>��o{;���v{�p]t�}�̤pr��Q�ٶ����
��n��FŒa5Μ>)Q�{7<�x��`pK���lxͮ�#��W�W���Mo�K��J��Y��Pr"�����>�rCl4��@��x�X�i���j�/m����:���R&���M#�H{�v1�;��g_Mhd�rx��wY�i����Zz�ڟ���e/���_-������{Z �;�`���}y�=,4��U�{��y�ځ�����3���-z3��d�s۾Q_W�Y����ڵ�ۺy˾;�K���o�K� л5�I��ł+9��asb�h:v����.��wQ���J�z��X:��n��ۧ`��]
1��9F`��(S�Jc5����a��"kF��%ݳw<}�㼧	�R��m4��E�)�SC�^��wqhˇ�:\�k��U�N������wI�%�S0��*��(_�'�)�ʜ�v��3�U��)��V/-�Nj�f �ws��<~��<��cgӞ�@��(���w�j��:,��$k����'�vh��y��|^"2�FI-��������{X�.x���;B���H�j���r�xF�=�`�f�&)9����	�@.t�uo�lP̏�g��Q�ild��MZ��Q���Ř�Z�
��ta*ZLN1��uh�Jq�x͓uCf�ô�3sU�;ސ�O���9��k�:��C<��Ev��sqka��a�"8�@�M3�}���uu�y��[�1�n��O�  E�W�@�� ,
0}~!��ᄣ9��i5k�<9b:�5VSV�ðٓ����y�<D����]p�1��Ɗo8-���s��`�00/%�ж45	w� ����x�����^�f����b�5�1�˫v��g��LZR�������݅*]-�oKܼ��W���o ���U'-��v�쉇�ڷ!m�k����˴�CK�h��;��z%B�苝��w\ҕ�gC�y.$���[v�O=y�zb�v`�]T�ē;��׎#k��d%�¤oXW���
�g�.S�`���n9���S{]������<�Ť�F���<���d�4��e��q���9�u���M��ɰ�s�.Q�OE��Ψ���3��ek��c,�i7�i�I+űŖx�0|s��v�acg���v�R����K�w&�d�@�����ɹ�N���k۷H�9녙r�F�øL0�����V�W@����q��.�P����:v�%Jm]/[3����.��;P=��ǘ��m{�NA�3�6�q��1���%�Hu�M˨ƀ���n�1�D��'9�����΃�䵱k���w74��Hp-C�
��p�{�F�]>��yFv�C�їHA�Q�a4�0��-�Y���8�����1ɢ�*�Κ��	D�)&���iyf(	X��搭�&��`D�y^-�OE��$�)�\���6U����a�87u3`	nM)����&S\F�eL�,2�[��d�,,K'�@�Y'Uu���<v�-��*0�8���B�T%�f�C�I�]&3J���`�e{]�w�_�l3�[�Z7PY��k�u��^`��p�($�#K^[ks��i솺��s���8�>//D��1�'=c����T#�{u�/5��m��Y^D��U���[�.���@Be�CtX�*q�7��^[
��0�v��B�ؘ��;]��)�wc��f�#�cy�r��mE��ź�n%�[K�!�6jK(
l��/"p�"k)r[�]�������H�i�]&x�[�`�bZp����,���!�$GjF�e5m�6�B���X�ob�}�ׁ�X�.Av�aݶl�V��n�8Hzxy�Α��m�ɮ��1��X�P㡌0
��$��/Jx}�ٞ�I������q�����p��qŎ�G��]�x��=.Nl�S��r��;�a��8�-֍OI�IT�ⓞXLv�c�L��	s����'�	�Ġ��<3nώ�׫��ţ�n�����A��eȌЋ��2!�V;#]2m[`St8�Y�mD��4ac�3��"3]c�#����3�1`�r�M�m3��K	��a��U� ��T�Sr�V�P�"Wv�=d�3�onz�r�x�S�H���9��h�̥m��/Ol��=R����݋����bgJ�6��m1-�V�hk�����)����Z���em%͔le)pq��Ȩ�r�4���Z;Mn��W��0�\����9�ٸ��q�
h��)��,34@���n�snxY��r��Z8-Tu�SA��/���-��2]��i�H|�u��X����'���3�`�Y�����Z�`Ȑ���L3k�0��ff#e��xvK����r��ק�Dы깋n��.�R��j�vWs���'렳��n٢rݸwgp��{>v=�na�����L�ճ���1lqӓ(�9�1�1f�.9G�cYmWfޞ#.��2B��'��g�>2�E
��'$���d$%��k�a:8�Yk���-�qu,ۘ��ĥ�V�.nu�f/ "r��n��E�H�W0�fB����i�CXpKG��cKgs�v��)��Qq�ntیS��ۆ��#5��H�!.5ѷMqJ<hV؁Kfu-K����{;�lbv�t�`1��ζNE�9�ge���A;�313�uϥ�5��nx��\�ݞ6+�zCn|y��$sέ��5㭁���Re����֡[MJ���y��=�ع��<&��*Դ��Pb]�2�f�q���+c�.Q��ю�u��v�0޸N�+r`�מ�v8k� `ڀ5O>n�Z�\��F,�YY�'��O;p��v�3!�Sz��۲S�MM��5ڬ����Vn��kh}���r���\�6�t�ѹ�6ۧ�K&�Kn�H�u���)��4��#��B���ɸx(Sv˵����un��nPK��1�ug�Þ���]c���Oe��l�c�h;LG#s�Fp\��d��ݵ1��`N�'��ن���\8�hzZ��i��r�6a�����lнh���<�jYV:�]�p�i�������MJ��3P��X����ņ�Y�$����;P;-�ʽ{v�q��bW;�']�NN�u��wlW���o'6&t�%�hc&��|J��;����������9������6��m��nB�J��LZ��D��
(��6���,�u⤎*ƈ"C�ҩ��G���n��a�`��싶&=���7��0ȊR��Z[��/�5���q�t��4��g3.V^c][V��l�Y/\�つX��[��Fh2R�]ؠ[��ݫ\t�Wb������������V�������\�Uu���ڮW��p���l`c/Ω7Gn�G�0��Ѳ �Ò���l�eS`��+�Zuŵ�T#�n�m�f͒�
�T���`M���p�Gs��{X�=��]�ks�H�@�Yv��k��dͱ �n�p�l��q�&��r����F���V�니*2�v\0���Lrp��b�������6^��@�@�Vj�e�*Yyf,�-��-�ڨh\����G�p��iD��F�#�V�mܽ���Gp�lԋr\�_��Y�wOR1,PP�,'L
�
�X�R��!D�H�QA�� #��ԣYt��b2YX�2��t��+��ųVVI���&6�� VB��
�i2Ң�)m��)P�V,�
&!��iaQd+��Bc1�b��1DPr�R Q�,�)���ԋ�m!�����b�`��XE$t�d[l����B������+!R
,�(,U၎ �J��"�� �`Ͱ�1*b�`��U$cQ�B��-P��o�k���˘h�)J[:�s�->|@>Mv���D��qX�j��&$%DΕ;OM��m�u�k�8�T#�p�鋥�K�+γ�u֝ͶPw!��>7��ro]��\�`3�V��Ŋ����#��qke���b�k�#Y�jE,��w�d��-�����69�V���uɍy��kY���Nt�͸|F������@��#>��n-�4���EOK����A��P�ӱk���qp�B�;��+�x�\]a`�XP�^�ShE3,Ѧ�&��n&���.���Y���a-Q��v��	^f�Ճ�ꈎ �M���ϙ�]�.�p����>:�:Ώ<֏&���ŉ����5��w��<�v�	ms����Z�R�ݑ㣋��BR��QIv`�fҭWQX���&+,�R��J��aT�6lܚP�6hc��k���b-�8�u��s�T�ŞxwN�Ov���h�=����)�x���:�ۮ2ay���Et��Ó[6	ӆ�UJ�U�	O��6xx7Q�P6�5뉡:;>W"�pg#.��u�˦!Hr�4�0NIɑv��2���G�&v�1�����P2������s�/c;�Þ�y79�ʜ����s����w#���y;r��0�r�Gs�����*=�y^�痱� M�{(�/����~x��;!|K�Ҋ�6�z  ��Ƣ/��f����;�!PQ�u��&6o�"�v�d{�A��FQ}�>gΔ��ȑQ ����OĒM:U�v3�\!�l&�Y�2��܉��ˋJ�5�����"��"g�B����_7^�[ӹ���Aխ�#;dy���/}N��[���u`9�c���pg���We�/�{=�6�~��(C�� ݭk�,�М�E�"ɦΈ�3D?'�?��	�E���n�w�\`����ӚU�b.�=�MB�\��5=�sc3� �[[�)�I��uQ`�n�D�C��z�!n���S���d�@Z����|���$��#%�j�����I��l�qT�ꉐzy�`�	4�޶��a]�V��6����gW���e����x�fMh�A#-e�.Ź\U����&�_{��d�5��w@�ns#6z�����I���/�Â�u�D��z�fcV	"�Ҙ�� ^�yd��z�#��b�ֶ�wB�E�wL	�q��Z"�Uc1�g*r��3�x����(��r"7����=U|}9���B1�"!Q0�T�wzl���.$��D���Ƕ��VJ�K�l�	#��@��^YV*¯r��י��;�������}V]�k*c)����:eṹ.�2�|�}q�̤ӑ{K���/����q�{�y�	p��(F�
ozU�]mNL����`�B ��򑝑���F��8)'TET Is��tC��ޗr�� Og?a�(�a�����2r�|}5�D�6^�A�o�нq�ꛘ��������'��=�(�Q��>)�)����*���|DO8�w͠B���oma$V���ݖ��Wj�r�q�����۴=�U�=/3Sp���$�G�#�>=Լ�3����S���3�i��rOe'.׺��j����<R ��ϻ���NrA�\F���i�ަ �rdr�����[ry!�؄w��4�62��e�k}t����b����|i�]�<�>��m�����o�bӦ3�;Fe��Z ��`��(�y���M�/^�f��pa5�K��>�B���&��*oF�vU6�A��ڶ�읣��Mq-�`���u:^�[#[r([r���A�ˠn<�*��K���t�,h�mD\�c��̠:�`5���O7��\t����gn.���Ocb�)�Y�m=vn�9�qMft�.�jLF�a
�::e3\�5~�߶��V����`@;�%��h�e��e:��͂@��7���j&H��ㅷN�f�
��� ��A#���n��Xɗ.�������΀}kz�OV0�'c�WE�%CM�u5+�lLK^}Qٺ�v֨�����9
IГ&�.y�t����H|�l�=�������7�jm^wkR�9ӓ������᧠����H�K�ڙ���ڋ��hآaoDB�a�UO6F2{�v$���L�Ǹ�_f��ug�]�oD]��{�4�*�1Md����^B����u��i�5BF"Hu "o���R:�A �歰ŉĶ���؝O���d@�����7�>��/�%CM�J�A\��{�U�=Q�^����+{ٙl�)���6|���1ne�ѱ�0��?>�{\2�w�]/��n�E�Ub!�"�\�x53������[�sD�������H݅�;�8���� �m�+����ZWW=�r\�c��A�ȥ�'M���~�`���i��w�d���j�=u�� ��D��*���G��&��"9R��lI݊u<�؃ϛ��l8M�������&�ǯ_u�"ܦ���-��b��Y�U�*���g5��<m���l��dl�p�nl��T4��lUj~ F�J1N&�nSV�Ŵl8&e݊�$�D��E��=��nā�E��}���rfA$5C�4�z&s��׬��v(�[��D5U�}��j���jS��=��\lJ�S����VR_��t3��2�?;/�~�A�����{,�7�L�F0�&>�F�r�V�O��s`q(w\�s�߾���5.p4nOî���(6Z/6�r�s����{������1È��5�g[��e ZVj ��L9o���}>����L@*�Hg?GRr!�7�ʨk7
I�U�1r�S�T������ā��gڵ3����S�ב���J������ә�4�FLZ"��^��l|{�(�L�&H#�����r�e��S��J���W�_jq+���՛pA��G�����y��z��觼��C���::�:��<p4%���13��/�N�����y��I��bj��u`▧{t�����c���+����n�6e�V����lX���S�a:��r�7k�ܙ����&���Ξ*
D��v�,>M�\Z�Q�1�T�5�G�M=^J�"�D���:�H���#�Aͤώg1<\{K��%��e�Z�Kn��&"�ٕ\b��,ۭ4�O�Ҏ�Y�0E�L9n�m��*�Xtx������`�����n�읇$�EPn���]�	�>���w`D�V:O $PF��h��H�*U���&4Yu���^�^~9���B�T$ԓ��0�򝱼�<G/V���}~�y"vq�w�� wd� �Ğ"bI�����'o%I�JEG��Q�V� �S4ۏ[g��Q��T�Yڵy�zӔ�V�aE�j
-����I7؃$��!��H�;:��٨8M����LA��O���b�ր{)�nĆa*;�0�Ꚇ_(�$��i�����}�rX#��~�h�p$�׈����!���=\� ��D_j��/~����y;�)�δl\Z�Xl۱��7F�9U��>Oy硊�`ͦ�D�ݬ6+ܵ����y-�aTqUU��1��p�ٸ>$�B$��a�n}���B��\�'0��ח�_<�4������'�05�0�=�����~���Aj{�i��S*�-S,��gF����7hgr0
pz,��|��8R�j,i���kY׽m�	��C"����c>��--1�/85q�ܟ�}VM�k������H˗J�h��o����q����nx����W�)S5���'�f>�C�z�8���$n�Z��;��x�B���;}F�8������ Ck���U���Eg����a���6��EZ3L�յ��ߪC1�j��V)"�SQV
&������(�p��xHc�W����}����m{X�7�=�0�7(��Nb�����v��\��GN�!�&{��7x�l6f=(�3��｢�z�ol�+�4u�V���󹬍�k/W���gv/=�۝yv��@��M���,�E�Ȯ��LBJ��x�Gطϴs>��S"F�ݩ��k���o��&�L��A�4������ P<J1A�,$|��bm	b(���ċĈ�T�0��0��J�Y+ V��U��:��"�0"��X��D�͵�����3v�DR
�X(�@�
H�
H� ,*C2�R
*��e��2�I������� ��}2?~���ɓN�",4�u@�Yr�͂J^����#{�?�P^�?@^����h)�o~�0���v��>��Φ	#7[3}��n�tB�����$tw
��S����YZ\6�ӡ�3/>���%�wkhC$F�)����/}ԉ!�C�lA�|Par@���lwr���8��C�ھi��bbmgMoG���/�}����L�(Q��y��⛷>=�|@�o�v1+�c�NW�;a:g���.��=�+���z����X��k������i�C����"_��.�:���n���o�Dr��̱����p{[<Q�]��͹ȷ	�sfƮ�%UK�'ƫ�>�'��/j�ʹ5����cw��h���B��W���c^�6�w� ]���}�w�H�~�bL�?2��^ޭM�S5 �6��iҁZ��8�:�W��U{j[���I̬��W̡:\�H#�"Iޤ�GX���z�!\���
C������Ԫ��c�s{�7{�eIؾ���L��z�!�:��kW6����R����@�1	n!���"Lu�z��u*r��pd����agj��m��3��s����[��%�����#(��AI�X�L�����{k�9�	l��*�M�	Zhi���4a��X+j�jM��ۮ���퉮���Gjb�r*."72VHM&۾����m�"����INf�B�ڟh��[B]Ġ[d��(��ocb����{5��A�.�i�=����ێ�)'^��'�X$ǯ����%���jߺ�$5C���n{���usd��ٚ#�9
���e�	l�U�;q�q�t}�_�\� Fw+�GcGU!�C�&	���N�H�h�Zdۍn*���;��l���I� ��l�g���)��E�6!V

�m�Tn �b 8Jn��.M��ڊ[�1�KV�-��n�H�np�֝�͔��[���� �J}br�����'w�`����z5D#��T�C�f���v�`f�29g)*^[�`�gqy��a���4�'TDЇk-,ɛD�Z��H��>;��y,��,�W�HK�`!wL����}I���^gv��Ă��@�I/*�[�h�W��;1k��wϞ�Itq�5�23m?Ä́�-R��ħ*� ��l��$Pa%�t����@{��7bPV�7Z�b�lm��^ް&��g��-�WNwap���w����N]�;���<�b��i�/�V��̺���{U� ���2AߡxJ�y�.%�]���gEaV�ki�B=蔁ݘ�:�ܠW����4rp�'^sH��Sr���.�y��
����ݟf�:��w�B�k�����f�6��.uͬ_�s��f�8����;��n�ݳQ4�����i%Pa�К�.UubƳ�u�J�ġ��7��}=���Kɩ��B���gGz�z�EtJ����T����-�Lw �t��%^��w�q��1���}�"'Cy��5{�ΎE����(�EUY�}�Im�d�d�{3��=�x��"a_���p���+�_�B7~16	5Ј#j�dn���S94*���	�"!@,����pҖ���WUr�w��y�v��xGS �X��g�f�2U\+F���\5
a�D�6�kj�ء��At�#wX~s�K:����})�"U	�lA��b�L˭+-eBfn�{e��M�fb�������T���`!U�`�N�T�7B��S���ۆ�f�1Uǽo�U_�g�WkM	�W�"*�kw��ޙ������,�ӱ1U�5zr���w��fWFؿ�x{��?o��cB�k1N�v�3;,p;�Ȥv����}\�fsQss��-��7c�ǝ̝��5p/�����k]k. ���]O=3<�w=r��[�!�E�Лsp��N�e�՞�)v���K���4��*���:��SL�CF)sV/��~�㝚�n���A��� ���s15)�R�3܎f���$��!�P:�bK ������v�>cOb̈
��B�}֯=;\�3=)�;�{\8��1*�^��v��
���\}+����P�mrbd�!h)(���U:�.����lAމ@���ц�Cy����[O�pK���c����`�WB\�������Z�O�~��$��_5�M���iZ��Nt���mlW�OQp�B{|����������m�}"�N���J�S��7�d�ܻ͝�����7?~d�+�@���$��-SѪҡXI'>N0�:�"�m����$����n�G��)����:��}���Lw{�_P<�-鉄���Bk�� ��m��T�N�yn�ě�C����aA�v��O$s9�i��]�i���6�IG�c�ݤ����8{_��	����4,&�74v ��W�#cH}��������;	�Y�7��u+ ��a�atNs5��=�4R�F���eK��\;�.��nxO-+�oH��p(��{�x =�ۏoZ�	#�l�̈́��:�w0�Q��S�k_�͉�9����s�(��F?C�`�܂1q��a�+��{�\J��~Ή��Q�4�B�Ke����4v�f�Ek�������߾��� ��õ��H�{�bY����j|%"�IG����P��a$�F_07c�3jg\ŴxZ�-�n��O�Uq(�%[�r�>�� �v���wa5э�l���Χ�W6Fo6|}�x��j�k�Ƚ�S���j*����뙓�u��,�k�g�0e�l��]�I�ØkT����=�{���'�o[��a%��Nh�<��� �&g�d��^ �s���]�֚{Ϸ��%�lT"�e��a��tn�ʮw��m���j��u��.�J��=�ixu�M+��g�*J!�P���&qd�u�u*��CI7��;y��A��پU!K�ff(]�;�y�����&,`'�j �rd��B�m�uGw��^$I'f�>����_Z�;�Q��͹lr�{@_7��ۜU����o6 n�p��.(��,�O�y<�������^[�����n��v��I41Y%�eL���v����>d��v,����.#�����;��b�釼|����]���M^�ӭӝ�_5�ygZ�9]}O9p����j���<�rt���Dh�dߖ��	?N]s��t���۝2_�F�y?�`�b�;d��h`,Rp�>�	͝�j�5%П`�5Y%����laOe!0����X�9�l�Ǌ���*�n�\
�wU�кyί�;Z��4���H憹;sx[{5�$��b�c���>��B�|�L�މ����G!Я?N�T��=��!�#�ش �M�&hy��٭�$�Q�b
�S�*f[�z(����[&Z��/����"�8ϐ��KU&TZՒYE${�O���Jn]
j���T����C��s`c��}��s+9sN98���a������}9�ۜ�������E�s��6w����D�ʐY#핀��3�UV��X_�������+
����*,��D"ʀ�����Z��X�XEH�*)"�$ĕ�14��F�R�d�L`T��X�nd̡�P�Bi!��Bi���P4�XV�&�PXUHT�J�����VEXT3,�$�����m��b�g8w�}��I�X��	�NZ�A�!q��#S"t��Vu��I�PΒ ��('v���-��K#�e�5��2м�� n�pB�+�2�%��sejE��Vd9��g�8,t���˝�I�oe���㛚nl^v�rp�t��T��ST�;���2�+� &�ÃT��拱���ש��{y�s��v[a�5�u�5Rl�8�ݕtGV�J�m�6s��O!f[I4xM�:��.p�pu�]\������v\�R*Ba6���d�����i|뜖\d�`cdŅݠ��GK's�%%�ҹP�b����#��g{C��a�OkS�e�s��磒wO|�[Zb� ��%c�q��i���$��Ԛ���B�3E��#��ĵ��(�S��X(H�[����9�.��c]���v�c��6��A���21�m�җL�#X���<��wn��p�]m�&���9�d�}`D悷N������Wj�,3uP'4q4gY�Ë���2����>�'��3
۳�y����YL�ЖD.L�UUUU�f���l���;,�۶�MԌst�n`-7X:HL�D����fP�Zi�]֭�ۋ�c��� ��y���ɼ�7,v�q��lB�=�ǂ�˛[r���&<��{�&P5�̱�\���,ff��74g�#<ۥw�6��r<v�o~d�=��H��LT˩�4v�c2t�ϧP����멘9`��ƭ�҆���r��������l�؏[$6��2	��s��c�k��M��T�5H�����W��@wt��׸�a�R��>q�iyt�u_��i�Z
W�^�4+����l�b�IEݪ J�$��g6	��m�+U�I��#4H��p���ZIIQ�[6gz�T��;X`o@a�f�� �ώ�+�78����[�kp�	����"ӽӼ�M�U.$��^`�Fr�;��~���>"��՚�-	5��P������9�䧼o�>��5�mX_+%>�~��A\=wi�"f��1;1
��d�}�x�{�vb�'�ڀ��(�5CF�Yf#����N6#�1�}�ƌ�$��l�5��(�q55���"�`�{��|F�yvs�&!�I���"6J(�� �R~��̬��&�$�sd�x=y���&�K*Z�3��5�t̻jʰ����מ�g�V�S}��+��P{�ٛ�ձ��}�����T�u!�<�v�9�=|�A��-�~{�]ERR�7���6��( K�L�A��ssg"qC*ӝt�&������i>��G��T���56����͋��_����S�I܏-�l7B?�����D��q�@�v���j���^���(@S�MTTT˞a�s���kڢHݤ}u��<���k�����:9r0�i+�E���]�����ɶ��O�n��@=�mV�?�wB�W�mvhZ-�nh�b���3ќ�fJ$;�'s�`Ҋ艎�<D���#��>��7M�iwЈ���v�w�����U'�S�W�|�/Zh[�k�y�L�>�fX�����D9��z�-(�"�V�WV:5<w�]��o���M_�?�� x.�|E�t���>TI~AEgr��+g���g��z��0C|e&�jLf�3F� �ŮFlާs����[�U�`���lI������:uAV��iEIG���P*���T_���� ^��U={9֧���p����$UB#�"a!hbZ�NI7|�Ч�9�@��v8v����B+�P�k�WH{0�?[�%h-�>n� �3�%B��f�d�7�}]�s��l�LJ�s��U��f��2�
y��ۄ۾s�8sv�<��G3����HI-wKͭ3z��2�,�����͑�Y]̄]M�&����v` -8ې�U��ŭ�$8��;�3m��J`���k�v"�+l�t��[��ŗ**L�-u�������\���]=O��G;q˰`��-������Ÿ�X�skϽ�7�	�_�kZa��JokZ�w�ɫzr�; w��蘄��W6A��enS|-�R�n��O}4gg���S1BQ>#9"ޤ&!B��(��D��7vhZ-�n�����Yʅ�K$m �[�?y�L�P$�Bl@܆����g�\�����B#bE��]*>��Jq�t��Ӻ�P�
)C,���,qj\6�J*��]��6��|�H�],|{�S�1to�uǐ������GS!8C�Mmr4�}�mZ�}Sx7R��!�s����a�t���\����x|�?e���^�ߍ�
��h��`w��옄�}Um�Fu�͉��ܜq�3����͟�)EID�;�����ܰ�e4ދ�����n���-�n��bg�I;7Wk�o&}Y�?���=�����p�%��2��օX�U�h�.j�묜�iAi��Dְ�N� cr�߻���]�l�}Ρ�whUP�[P̂�^�폠�����(�d'ISɒ�H]�^lM
����X��0p�4*E���}���v��)�̩ �^�l��mi܉��m���r��*��|F���D�%UU�S�퉶|A9�7��VG�s�>��I���$�H�^�Ou 7.K��$��Gg7��T�㐽���B�'C����-6b��K�Ư���'�[p�|w1�H�A��)P�����;���|�%>�VA�u�0�~��� ���+�a\����u�r��UUt���}b�� #�$��a�Tu'	�T�=f�j������d K�b�뽕56�g-�{��`=�c�v����
s�Mu�8 ��TK��{�� P���'|�	�b����H���n���'wXy�fz�Ӷ����X4�K��6g.vK6�`�)���<;��.��!;�� �R��l�c�ꁮ�	&{�/Eи-�nFWc%%�8r`�	u����~���[�Zk�jG
N{m�Uv4�{�ނ.� ����Gw7{[��Պ�w��{�,ޔ��u�*��{�i���}٪k5�,:aS^�6��R�rɱ�FԵ;2����H���|�>R������]�}�!���U�V�}|�~[k��UjT.���҈�ٻ�ETj������>����9�2�R}��YT�-�NV�)\/0��S
1&�fsU46�d���э�iݛ��c�i�*@^9�)8b������.Ô�(�.�2��D���񁦉-��L,�:�N��U8��Mu=s�0nN�k��wK��;JTx%���h��b��k�g��з3���'<���q������6�IR/~j�L*N��z�o=q�>x {�xi��T��S�;�4�����y.fpbA`��N�
Cz�����4�^c��R�y��AH,�_}�bAH(q���<py�0�a�9:����n0�0���I�*A`��C
��s�ߜ�f�� �-�>y�l7H4�+b�2�|�c#�҄܀$����BH�莽y�����S�{�"M�RT���9�1��%B��{�m���9Ï5η�SL���Q�;��&�����z]k5��-`��C��-�=�I���� ��<�@m ��d1��T*J��w�m��V{�����jK�s�M�^1�Vk4l�X�c�._�O����g�@��7_pI�d�+����2VT
% ���`��u�n*���"M��m![�y��C�s}��qH���da A�z�Ӓ>�j�P�1K���&���5�3CU��\�M뵱��M]�o6R�~�`U��>���η�:�>$ �t����m ��
��纆0�
��T�;���n2�N�z���<�4��m�Ǌ�]��X=���� �)h{�H.�����9���ǽ���+*_{�bACI*����m�a���:�l�>|,#�P�������x��Q���Xhf�
A@�q΍�ڐS�}����q�$��߹{`T��Ns�Y�5� �p��z�i�
�YFJ�s�I�9�}t{�������;aXu}�VT�B�u�8i�l�x<	��zH� �狺gk���3�5�e��97gWkR(i������i���>0|.) �#��H[@�a���R
l��4�bN<{�@m��
�FJ�P8�4�l+����W���aS|{�i&Ь����<߸����a�1���Q*<{��jAH[O|� ����=a����]~Px�(*T������$t�R
w�Xm&Р���+A:��;�D�����͟��A3X��{z�]$D�^	��nz?���ϖ܇��Yrp��$���R3��n&�m��~�<o��x���M��[F=�6E�[�cT�+j�n4N�Uh�l�7#m�J@��=��g��ߴv\i�����<3i~���ָ��jg����7����>�c4�o�ٗr{,�������y�HO `��w��`yx�Ӟ�d���ۗJ[�3˶��?{�H�t��ƩŁ���"��ı��n�z��pcd�}�l⽈503Kt��p�h�ztTEOnԯ�%��������l�"^B2�M���K6���F.���ލ��yRܽ����p��=f�z���>����F���G0�Zz�|�׳м�
���q1/*����T��*x�j:vܭ���5�ƈ���Nވ��l���& ��!`"��F���/y��}8+ݷ`��8Rٍ��Pi���E�:��C��0fF��q�������Y�~/I�[Y�"�k&2EI+1
�!r�K��	�V��\m�!�2u�a^���*"�Փ2�J��kB�& ,m�Trԭcs��)���`bD���X�.3#1A�Y�C��f��A��R8ܱai`(-j(���R(�̵`VJ��Zҋ�+ TE�+&ڈ��
�i�Hu�o��aRT*?i �m�����/p ?���s.�`s���Ͻ;��Hsi~���)
сZ0*u׸�
l@���y����uθ�M!�%@���L6+vq��sZu�Æ�=��I�l�9��c%���H(��4m �6ԅ��y���
Ah�y�B���h�׉֋�tE���c��ە�6�"�"Ӯ���� $�.�G�#��8��I��+/�
�Rs���Ä�O}��m� ���p�hgO�W2�Bπ��◄���޾[y����H) ��|�@m ��+�
��
����w޺�8�9H,:��߮�e�R
o}�IȅH,<��c%eH(�_��~�O>$ڐ��}y�ot�i
�s܅t0*^͞W�V�� �9�8��6���=�z����YY*{טlI�*J�XY�{�VT�
�n��>�d���&�i�_F|^�5tnwT�ފ����X�yS��x�=w�;�׷_ I=���2�VT�|�@�����2�c������ �||s���*��
�uߺi��R��<�2 ��%@��0��|"F�
�����
҄Ae@0��h4v�
]�5���5v���<���kN��8a�
�{���J!Ro9
�P4%@�}��i��7�7�AL�x�t�h�Y�B�`T{��=.��k`m8I�a��͌��pj���8���=á&б%H,/ΡXhaR
^y��6��YY<����:�=�.۔�X�k`�c�.�%��������HV�*AM񝷏5� p� T�e��!R
T��$�����]q�*o�p7s���8R
Aa��ى �Y�}ѶƤ��y��^���� �!��!]
����{�r�8��'���h ��T�ް�M��]=w�R/�
Ö%�,M��H,�ed�*{߸�2��-Y�J���!L�{J�Ru��s���us@��Z-v��G���0��,[�_���	DED"e����g��wi�'e�;L�s�b��YvN�1t�/��p����j8X�� �.���NSY��뙛\`cn+����ΧY�м.��Ɉ�<;��G6��!��K5.+�SN-q�|k����ƚ�񦀶׌,��.浘�kޏk��s/���Xw{�Ӊ- �{�8kt�l`V�
�����M��^���:�޲ ��J������.�89�u�]k�r�S�z����VL��K�\NXwy�VM��T�=��H,�HRӯ=�6n�m!^�����xo���=q��5}�׽e�9�p�<��4� VVJ��8��Hm%H,5�~����ޡXm�IP���d�+%ed���~�$$:�
�\4�Y�TJ �P�t�R
:�yHT��R�{ހ�AM�VQ=�r�w����� �o|a��+�֝���]q �{����
Aa��3=�^qy�x��㹴J�N��F�jAH[N9� �A�!Z���B�4w��7���Nk꘿E�n��r[��m��κ�e��hω��T5�H��U�G�>��R
qߘlI�*J�Xw|�T���7;������@X�>�x��$x��0�M�R�n�9�e�Ă���@�<" xxP�΍�]5�?����a���f�Y�������on�5��.�Oy\
5+�T7׼�6}��4� �<�[��)
�H)y��@m �n'�f�*AC8�s��t�9s0�C
��Ӄ�GZ�ָ�)8��I;��ea�6ɦT
����Y޹�wƺ8H)!�N:� �A�!Xy�:��/X�Nk[i�O}��!מ�s�sv��{��uŒL����]�ssI��ʞ��H��_L�N��\�n�.�
B������l���`��,�� ��� d؁R(�{a�i��D�
������W�����=)�Y��j�P��D�]�ř]�X����5s.����=�I ���H(�P/���l�`oӾz��Hsi�`7H6��=��FN��=�"5 
"��_�I�'�:�ۜ'yԝ�{�I��+����*J�IS�|�i �=s�s�|wsZz�<����<�c��.e�Ăÿht� �-�{�8ke!Z��`T�}m����}Ӱj�Me&�܉8�;%m�
T��*h2p^ƍ�_:�잌�.�I�����+��B�4��y��m�aMxps��iָ�,9T��0)�y{�r�Y:ea��!Y5P*T8�06H)i�~`[��"���|J��<	;-JsZ��w�8i:@� �����m���s�~tN�x°�gZ�a�%B��;��6ɶT��S���4��7Ϗ�z'����6�遛Qj�����ZB��s����F��|' Ë�G��7ǘkt�H)/]��6�S�����]rL�'Y�B�C%B��Q=���v���W2�)=��m%B�y���뉌=����H)��z6��5�Z�S�}�7�AH.��}l<猅v��x<V�9�K�_�1xI@�@�@����AH,=�]��|�{�x��C
�RT�a�M��J�׾�@H�6T%�} 33��I�AHwh�5�B����;�H	�A/��G�N����+��(s��5��J�lNmN$�Y��]ݖ�q4��7F����g?�����H�s�8m��VkÃ�F�N��9a�aS�~06!��
�YXsy�VO�����4���^�i���,�����Rb�
�S�q���瘟�iV�HJ�3�ne�GdPa�	�a>��jP�M� �>#�f!) ��$+/�
�Rvv�=֯�㐩;޷��&�Y+*q�xM��<��᫬��.� �7�7������^R�
�R��ր�m�+('��B�4�����+�8w���
ß\���̺�����P�Ad��<��+&�T����=�a��m �9jB��u���)
û�B�����q]:́�r$�0�u�{��Y�J�2T��p�I��+�w�VT�B����O8w���߽LH,��ֽ�4��q��[�x1��Xu}�Ӊih��H/��q�n	7�h��*T
���B�C%H(T��$�I���ww�ѿr��l��ׅ�S�]�Td·n�r���;�U���m�r��2�!׭q�xz���a�ۗu��!=p�b�E���R�T�p�ԕ%����60V��Q#��kfl�-�n^2�s�v7���Ц��6�ȑ�K�"$�K�kc���{$��EDMՙd9�\�.A�K���+cM�u��i�V���-���N羅S?�OO��I���6��T+%ea��!R
A@�{�I�q��	΁�G�#� �0 �HV��{����/|{޳3ZsZ��{�8i:@��νԛN��8I��°�=��*AI�*J���d�+%Y.;��5�3����qh�/Fg���\�9Û��H[H[@�a���h��`T�����x�@v�R6�gY
�2T*J���p�@O��8��(Jx<	�@]=#҅H,=��+&�T����Ƥ����p5�Ϝ�� ������H)�ᾲ�́�u����I�����ł@Q����o��m��-��;�F��r.~�a([pp�rg�.����<�[����0$��0���تY۾����B3t�|$U�CfP9\ؚ�8�����V[�7[�ˬ��w1�4��ɋ����{��7�� �/� �+~lA��C�w�U&I�-�M�m�u��(���*����mG��@+�� ;��v�4%��N��ё;1�����'Ē*��Aæ�㹳���Ȇ�
I1%�?0|x�P��Rp�]m�|s�����HuG����n]>�4ڲ�D6�F�RTeu�a���������L����.��/!�T��4>7=<j"f"ѧL��Nk}^��$U��P"�e�quJkr|]	��-�5h�k`��P =\k������Ve��6�U����¸V3���J�ۜ�Y�d��H���wO���X~������[!���-�Vt`����Av2��UZ)hm'Th�A�U�d�&#vp0����fv�z֕�Ϥ=+�%.F��\
��`��i@i��k+y.E$��uI����?de��@��lv(�t`95"m��!I\v�7ӈt`�{�{����D�.	���3F* ;�X�z&+e�q���gӽ�?2��CdM������zl�cL[��QP��8�kh(.8j��SDӂ���T�#-d>��6��
�"Mzez�+k�� ��?�@�ݍ�l�n{�lO�j�r��ϕN�3���!�Xڄ��@"�WmT��GM1�,j4�o�1B\I�4����`�N�6z'���P�#��Xt4��~}Selo���� ��`���ڷbd�3��."Q*k������0O&�g;�WB�����i�L�	��8쁧�ν�� gt�/1�q�L��Tk�f2��CdM-��Ae�\/{e'���cJ}�1���9K�mIYݷ���XX�n��u+����F\�{�c��"l��A��v8�}�	>�}�����Tm�U�8v�g=�������F ܘ��m�hQ�c�]zn��ݻ�ga����@ �'�A.v�3�qD;��Nw&{����1���<���8��!���0xS=]j\��Nŗ׎�-��t�^{��{�o�<��j���z�s$�\�aͽN-�:4<��Y;�^J3G<�h�-��Ī��t�l��:�u�oq���TT��ui��7�`�J\��#�z]��]�n�>�O8=�'��=0/���+�R���2�E�Q3z��۷�j��A�
���o݀��_���RA�n��U�Rg�a��a)����o.�rW�W5[�n���>�u���t����\;]������ۃ����^����9U�M���Ӭ�y���D������G���d�f$�h!T�$��E�ĕ!��Aet��N��XDL����YV�)\�m�I�E��	CaRV6�A�2)��]*J�ƸŴ�M��C+UՖ �r�i�B�kQl��X3*�EJ��mkb�]\b��
�%��[%/r���[Yl�mm��-a�m*�x�a�Ә\4�L�:8n˙ 0{x{�5�6��,ؑ�B�yfs�[.{3��ܦm�\3�,BJ<q��ؗ̷�x��k��˭��\�ܠ3�z��.�9���"�Fѽ��Q�-x���fCC�c��K�-��:�h!6Y�GJ
�ۛ@���A����Wf�[u��U�B�����pg�m��Ǌ7�i�Y�볁��Y���z�V����E��Ů�ܸC2��m�lg�ݳ��d��s���읎q�������=l�v��Ɂ���s��eu�u\u&當����=^��s9+�*������ ��	�4�l�d��Ecu�s�ۮ���"x���`�c��k�4x�F��ƕ��m��Ѻ�1�3-LD��������;�mj� ��8]r�w�u��q�q������q���Ϟ�.
+� *��[�qֳ�m�e�)H�,s9qq���&���h�X�T,Ԯ"B�1+��5p�r�r��s�
�G-�q�T�1�ȱ��=0������cWf8���]����r���ڨ�;�lwYԚ�(5�e��O���5�{G��p6�ܓ�1���[ųm��-��EvҲn����Q�A�!M��s��Twa�w�;qo0x�y�� nz+0Z�sf�U�/Л[b�up��CnkQvz3�(n���EDU�2�uX\b�xo�s���u�q��뱙��c��28�����_��&�6���v�$��^{Qgd���f+��P���u@Ѣ�Y\eY��U���FG����*c�4��V7ܿ���p��eWOb[������iBPT��r{9�	=Q�7q�;(�i��K ��^=�!w\��}�{�Z�ɰ@�ȐA��C�W�'\���u��.�n��Z32��n�湦�j����|=�K����ERD�39�L�eD3��������p�0���\I����~�\�¢d�4���s�Qw�W��o=���cGҬz3���?��2	�k` H߹�O�V��{���:��	`m'TET�L1*�sJ�}5[�����i6��W_a������
��#�wkorA�P�L�G}�&�%K�VI'��{��6|�	/u0}{�9����@�z$�K5"��Yt-�6�r�P�a�<6
Qˎ�'���7ڼL�-���1��}��A��E�مTz��V���]I�	�����'Cf�ތe4a��H�X	������~��}�\�M�c�`�7y���e�;`��D5f�;R^ERЫTݚ���=�c��A��sg��0���P���u�I����N[O�7�27a�M��d˱���,g�چ�r��#y,ܽ��f*��$�g��H����a+ȃ!(�L��h��f�f��}����(+:jߙ���>$��~]����\�$�r}��AJ#���3/ogUwGpٴ�$��lwB#4;]s�T+8�1CdM.�� B�������}�����DU�����ۙ��H���x��h@]Ā%�ם��:3���U'���7�,�O���0�jY}����y��U�����R��{�~��,�ȥ����g$��L����m
�ģ��[$34=�Q
'G '(�K65��p1fWf�ǯ>����m1��R`�: �rg�NOyu��L9T���@���J����6	�9��`�މB�t�x���[=u�\�W�Gݰ��z�*7�Y�c :�P#������6Dݕ���-`��H-�������Zt)踋�CPۯn?�]�32���@z�o�s�F�Õ�.��مRfE�@���k�j�aLc�����0q����������o\�����D�#�+�Yn� ���D���k��؂�6���� 8��C�m�乚��V�c��`�7-��A䎌��Vɑ��s�3Q�T��`v��"X����fI/=]�K���v�t��2Z�S��1�"��Z���}��evz�'_ �:����.*l_\��bd���\×/��lFE>Wk=� �y��o�F!���Fz������l�2�03�VEU��ŷ��7�l�
M�b([��OMx���`]��oE��j��Z��s&.�Cf���	H#��we�� 3q���^ݏy]��eІ�v%��b�734*�uƌY�Y/3";�Co���n6oD���e)��=Z�ۘ�V�i:�D���K�}L�(��:C�(E�٦�-�ˌ�e���ܸȜq8#Fب��"s��+�I ��`w�(�%�����_Rc�Pqm4�1&r���DU�ڒ]��S�=\߈=��V��	U^�����YEU_���`���%�'P��u��RarA.ِ땞m��D�&O�=���!ej�3��& _�z�q~b�|�9�F픒��;M��c�Alï��0�>��"�X�P=؃�>;��2#0b}ԅ��t��a%'�P'wX~4�1.7u:ɍE`���M �$��d�o�d��IXs�$�Y�����/Z˻r�l�/Uэ3nq��~�jk�	�D����X���8j��eJ�^Hz �d�͟vｑ��Ȕ�Ъp��S8�`�ssY\u����U�|�M���!��׋M��r���D#�0k��W�����1K��J{�X v���$�s�)�M�|�LP���֦\ڧS�1G�+[@/n�Џxa�C�(��І���`�g�X�^�����L�/���Ѩ��sDM
�I]�a��H$�j��݇B3�9w��&z��;����*��� L���p��a�ܹ�Q? �ՠ��>��e�3� �G�%�素:�H�i��KV]�4���0Ԕi��҇)*��Q��Bl��F���U����ϳax��W Ȯ3y�M�	;��ArAwF!f����g���,ti?λ����)������׭4"˕>̎V��靤��4<B���!�۟w[�T�{/���$�>�Ԫ�.�=͕X:
�'T
,RUt��w)����`
�ā�Ӹ/���u �ֿ��捃_�qy�&��2Fg�")��=��݋�;�������Y���O�D���3���0R�4Ɠ!��0�fK
�]xW��c(�q�AG<�.�v���Ѷ#�O���o������h�b�\�5���Nx��k��ɋ:D��g���:bj����C(TJ��3<���N�gq����ֶT��r���/����e��&�`�8|�w6nZ<��c~:8�\��v�eDݫ�l[W��T�؀��f�h^�u����}:��L.H"����� 5�[{=[������=���P�.�����uZL���6���C/&Ю�R݉AQQ˘5-�[��@.�m���e��<����$nr�z�\pj8����ks��;/	]H��^��+D4��I\�`�o9�2�����cJ96S/���R��61ӖV����PꏖmdݔHq�5��B=w�b{�>�H������A�b����©�BTְ�ܙU��2��F����gsL�%C��>�[t\�v��^gwW
�v�֑K�L�4g�?ETE�ڪ
eI$n�`��ۋ�8��y��(X�&I1�`e��aܖ08�����~�05-��cM ;2ZoB��ϻ�Dx�cn�t�Nh���N��v!�b�I7ܙ>#�>0�j����U�vҴ�-�$��d�;�2}��MT�����YHJ�ߡ]{�`�����3��W��Ͷ��ƫ/�����X!o�VD;=�{�.��8���N0;�L���z��nw�/�\�Ȯ����p �h�ɘ�h�xyx�5������5�����X}Jk�uGu�83|���wI�U��댞�e<��Գ������S�O=��#\�6.�C.��m˃p���Q'��n��3ܥ{����g�ի�����V���	m���RyTP�X@!{�F�ؙ�����&庇�6�svl����%K��+�k��ҧ�@س۝�zE8�.yo���m-{po�,��9���v����z;���r��]�vX�G�F角�r����)�;6�:�ced�׭��9p�C5��9��ܸ����wz�.LSs�h�Iy�n���Ei;�2]��qE��ξ/J�A�D]�����(�N��H��A�
��ZΩH,T�k/��l�̻��lNr��k�D���2��ʥ��AA�b,)���D0ee�ᬻq6��R�T��2��j���4�#l1�k�eb�2��o(&�SqX�A��m���ncF�����f�ZPwKm�j��*V�SV�Ә���"X���ue�`����q�.�b��k�(��Q��g��E�����@�`��TZA*�5�j����8��`�;�Og8�r�I�H#����I}���ɿ
��`������~ �sg)דV\R�;�=d����L�Xa#P�u�cW�NC�C��H�Ng6v�����+��	P���p���uݏ툸�c��SФ7��FE�u��K�dbNt5��D���s���d��@D��l�>mCE���7�ظ� �����6 �m�fgT�혽��Z��11��ZS ⴛ�f$9��:��噚�d��2��{�ă��67"*�H%55�2'~aҬ�+B�L��7�- �nk1�nԄ��3"�@�ո��5�ٲ��B���pGA�`����$v�fҙ*��g�s�L"A���Q�$�tr��Ո��L�{[�L�ɨ,@ۀ�u�24�x����������tZV� 7u�$�V���r����a�# ���w-	;��c -Zټ|چ�e����#�Fu�-�CU�$_S�9�0;a;$�c�-�D��n2���xTT�G�ħ�.���
���l}�v~��>���L�τC~p�h�A�<�=��Wt�����v���*�ó+v�u�_h:Q�[�5�1�~���(jC�����,p8k÷�lF'�!�;�M�q9:-��u��F���+T���Y��ڍ`<-�"�5+i��ܶ#(�fn�̏���_��~���$�jd����g:�k��5�g���RtJ-SS���B�y��H��f�#/3؂ߢ.rId;���l@�w �-m�wTn��Jz�]q&o���5�rh$�6�$�Ow7X��8G#�+VFA�bs�:AΦ���������{}~������(X����^q�a���ffWf��yﮮW�X!{�D.�l=N��(��j�r������1T[A*s�YW���8��>qʹE�]�yW��CB̍y������bMM@6�y�U���^TN*�����t{w�@�n�����+�DI:��u�{��՗�}���J+$�|r�Ff�r�+E3h�k!nu�N�$���m��v�f���-Z�$lٰ�Zm�ζϺ����`0�#U���F�|[�މ��w-Im�).9�r�7�2`ͥ���ם���5s�7W�:�LFw6s���0C�R
��{P�����Vϋ�K;�DT�.�o�n��n�u-�1�d��QE��:�~3�ߪj��(��	.�f�]ۛ��8��8�z%q��<1{��zpď�T;�ʏ�$����o7�Qɤ`ǻ����:xu?2�%�����ّp�;=��"��5�9́T�J�CʐL=o��������)�@����f�s����t����.�Ĵ�}}�������-�ޭ��
��Av�<�8BС�^SH	��CX|g5�A����ȇ��\����Á��ߦϷ�Jֽ�"�Zh�ؓt..�r�j�e�L@�t�ؔ!f�Ԯ��;.'*'�+�֗ cx^v(�z��R��/�q[�D���#�B��4�6���a{��5[F�4�h ݉@�{e�vw^��B?	cjq���~��z��M��;	i����z��+�����P�w*A�l�t��;�����
��ap�m��B��D�Qo�����{927ڄ�Ꞡ�+��(iה�L�$��o>���B�R��n��p�l� ��dR�`D\�w$A>'�<��v���P��0��N�QM����}�j��Yn���W��@�����u�fGr���w"�?9���J�\ezb���0�y���ð�y��*#�o�n�@�=�(�8k�NkX<X����&�uu��o[��Nq��3��v�&q����,��̫�Ƹ�	�n<���:�x�u.��g�X��ѧn[���\�ZZ���{F������G�sݑb�1ϓ����.��v��\!��G���f��Ԙ$s92�v.�Ġ�i����Y��l-�H̊�`nm�C�z�`��;�0�{��`�r4�\t	}L0Gw6Fۍ	hPӪ!�
S��3bT}~r�n�Ż���ˀ[V�+���QU͡!oL���U�)���}}�{���Q�Fb�
4q��72�ma2�j������Ϊ��I'���\�*J�qXS�i_���!��P��Q��lmu�fz�]F+螉��B�h+�efěT4˫����>��Z�vNXl�����|=�1�I9x�>#��Mʚ[�IԃW$Ҵ��9�r�ERD��'��LoS�A�����&dd�j[yݎ<1�3s��s��}����P'F)�g[{��#�\�f��~P{ƨ�w���̰�&�[9��7֜�pш�Tz`��p�$�0�qg�)�US����}��^R���H>��3c6b�z���n�E�0ɛ��i�o�LT?s�������U�ʪ�2kwq��"�Y}�� ��X�G;����]gz�7�f����՚����w����Zq����߼9WzM}3�l9$ҸP�:;B�|E�@g5I���]�r��Fć�Q��!�m�����i�v��D�H�-wl�Љ�V�x{���s)y���g��y�8I��u�ࡧ�C�DL�`�����;��Cp��{�gN�p�lk���ͺg`5`"D�&I'{��R��=Q$�����*�5��mr`�Q�>��A�͠gt�t�����
���K#;��������9�6=�;�{޽S�4�wk��p�?d��{�����|O�5�M}Pi}
�Tz�Uuy?]v� ��bt#��f�n���P*)���1�!&��;j�\ۋ�qW��7��e~���
�%�7�P�����8FgK]�	hPӪ:�C�T)�^�w5ݏF� ��ݱW��8-�$���y���W�jk�A �[`������Ț��q�J�y
���ӓ�� Ф���\�\�;���P��A�,���]W���w, �B��T��͙��t�=7r�F����ҵf�����{�v����yo.������$�=!=������ �s���;�u3{���n��P`ə<w^�����y�������o}�=��w�+ګ �.fE[����h;P�.�h�W�Wcd#{C.���sG����z�ׇ��:%��Z��*b�'[4�����v_6�+��Os�y��f�w�p��=��G�8�ܐپ��{�i��������xmg^�ʶVi۹�K��5�`��Nd�ĚA]���|R`գ�<�Y0%�=zy��y24�y��2B�	%��5n;*FNf�%y�C��J@�7���{�;i��V�f�aD����uwPLwJ�|15�di��S�{ao�ν�Ʀ�
�A=yD�8�M���TLd9l�PvL!S���}�1_cӈ����Q?3����!�np&��v���>�r	]:���P��1�\�^;Jk�O[�f���t�Yh�2飨#l̙e��īJ�Z*��Eb��WM�J���� ���%�Q��*�n\�ڻ̚MEq�bYEK*�tɑ�����v� �K@�	��˭5�ӎ!b��SY�(�-\�B�ۇ&�S�nL�܏���1��Z�܋** �mA�[J���)��-*��Q��5������iYDV��`ֳ#�G�Q�V5F�U)m��z4�m�C�[�%�������Gm�c�"X��vn�Ŗ�VyD;M��fl�@���*ɠLV��<uF��ܼ�f�Ф0��'V�u�n,�k�)�`Q��ۖ'64����%VS՜�6�2�Dgl��us�L=�ŝ�)�^�J\B9|طm<r]vvE��,a�;]���
zy7���4��ѓLq6�,��3��#v!�W;��<�gsϔ���{a�N��ڶ��Ŕ�L�Q(V��՚a���7 r"EY3 صl�t\���X�Q�2nm2b�K��j	���Մt���k]��Ë��.��8�aw��U�r�a(G�VcMU�b��2���#�5t�7�R�\���g`�Sq`X���X�f���F���e��Ѭ�17��-�X�1Tm-�hۥ���ӄƕ��F�"f0\�\i�]Ӷx�D�hL,dь������x�M���l�u��,7:���;|��Y&���qe�V�f�4n"E���u�%�ڗ�[���;�;[�j8��cr�O�o=J�l�Z˫�맥UUU��kk��<>�]�s]�H]56�i���aX����Fĉx3M[7
m-�RY����
@#���lWm2W<A૳�f��7h�[�\<��"�v��ݎ!2n=�K����c������>�-��>Fv��6�8k��ڇN��0�{)FN����[Fyz�m�s۩�)UT�N�h�N��F��C�<8��=Fm0V7\��6+W]��=��]Z�#v��IP�����t���]q?��!�m��ƙ]�Y�r�� �sd��q�P���=��SN�N�Jl�#�6��=��� gG�څf��p�X��a^��XwB$�Z�nmGXǗ���{�E�	0}H�0����#�{&W��"*�MD� ����o��*�9��	H��Da����C8�&�8�u�L��~O�#�$p�'��r��{����V�Q�X��0�(jߏm�y9�OQ�&y�%������B	N&�x�.���$�ٓl�6����<o���w ��� �J<4��M�ζϪ��D���V#�,gJ`�����S:�r�����v�>se� ���������׎vxٜ�ÇcT���?�鍌o�T#�p ���qċw�ח��g�a�5�}η��SMl�DFU��-774df��Ϊ���4W���Y�/�Q��>B>3y�^aH�Ii«K�^}�*���6�I�λ��� �]�3�ûF�6|�);�w��T��2!�߲'=�ȹ�_����u�[��u����������?"Y���6��G`�����Z7vZ UJf��z�D��$���hKAM9��L�`��M��wW���LH����Tb+v��T]r<[��9A�m�;;N�i��!15����l������<�#����Ǫ��m?��$5j������֙A[�?�4k��%7e�3<���0�y�BÅ�޹Ly��y'EC��$��O.�L�1�;[�ݕ8�7\�&T|:��{�b��u��{���z���Z����&r���2*��R�Ѯ�m\��9�\g�Y��<=��ϳM��ц��KH&��������F)g6��zp�{.����s�xA4.Qܲ�L�Z��V7ݻ$΢\��2�*�� 7���$�/�T����]Ӯ8«�b|���P]�07u�����Z�D:.&(@p�O ;�X$LI�o1�{�[n�ul�������`.Ζ#�I鉀]��Me��ûGv6��*�^G@SqjC_7�|Iʷ��$tq@�<T��h\���L�Av�0�	�[�+���;��	;m�<�z�� {`� �QDg�-��cOŽm��ܧ��cFǖ����ҭ������-+B�v#r������ke�OW<]��i�<�uH]��2,c5���1'�ۉ�ZWUU2�q;˻[����1�1j��\�R���tᅔ�t|�F�~~3Z�$���.7���d�O���r1���E�����b�8|^k`��_�r�]	�i�h�_��������r�UO?i��{a�ED�)�\��j�����$�{�V�0��o�ZQJ�$R0�P|��O���9��p�� ��@�t����tE�BV��f��u:�[4�:8h�Y�)�%��}�����ۯ��4��ٚ�:}�`�[�(�t/CF}Ա "�mB�Գ)�pＲ=Ҽ`���j��;+��	��u敄B|A�0��5�x�ߟ�?9�0�LL�6�0�n��`�h̡�<�$��R�v�A�d�����ꚁ���]}�Sy�|Y;`��Ξ�Y��J�-R1U�8�����v���uucLP���㹪sGk�咊J1��nm/�%�bn9��Ö8����d�ƜJm�Gǽ���n��B�(�H'�<�+(PJхGu��|��WXV@/{e�g��|V��ث��9"��4Sov��	��љ�'�\�=�\aP{�{�=W��.l�E�=pc{K�{�ۇ�ts�:Tz�]P���_3��;\��o����:�N^O��6X��kh4��T��{����8-�fq�i�!Y��VH���"�%4i�ǆM�
�(�Q�	���ne3�x�ղ�N�kR᱾V�]�N'��W;������wz�n��^�Ϸ�����[ �8��u�������h�F�V��[�!]	J,�Q��f:��u9�t�t�΁#��4Ss��|���|�\nll��� ���d�w�缀�8���+���(P�b��IÇxx{��W��б��U�W7�;���m�U��ճ�u�]���u��s\�,�9�2��ɢݴr������l(��C�wUeV�E	�ܑcA��p�_ 7lD�r=�x��.�Ӄ��X�3 �0���5����rO������~�� D��T29�dx^���5Y=�YP-h�*܋�A�-�TN�395��مsd�z�c��  �~�8ҏ����F���*S�Ҟl��Q����߅)��Ԟ˶!+�F᩷�8G�^�����nm�M�󋴇9A�9�k0h�;X��m�bNK�r���s����V[J�當���l��]��\J��v�b��#T����I��G��� zܘ�]Ψ��R�X�:��K��F볕_���7�����C�j:m��Y��m�ń�-�bgP�-��}չ^ջ<����ęI]^ΥU�vN�z�n/&`fmw�1��^���dU`�an��F�Q9����=��nV��*�U�fS�|�>��gZ�C]���c����;L�e��6�_;�;�զϿ2������f������H��v+¬,D�O���gc\dnK�wj*栧�
���3�M���Jv�u�(⺻5y����xx�|>�C>�}s��8��	���aˑ3�>�FꇵH^�^�h���I�zp��K�P6R��c�zV��SwR��15�2��צ�5����؝�;�V���������֌9��l��"�����b5�n�ɏU�Fo�P�:��xUw҄���B���Pf!jN��\�1�U��i�8�@p��]u���.T�lʉ_ǜ�N���R����^�H�T/�[�<�	ѷI�����>��xq��@ɨt�t��{�}��~b�)N��c-�ˀ�#������-�-K�\�ԩ�ٗ��y��	/S��sq_r�8h����CozLԃX:9�)�޽�bklq�\���<���9�h�)�q��3}Աd*{��|�J,.�P\�)[.�^�c��HU��B���xZ��7��\꜕|ϻԋ�����v�bEo��{���Em_-�����������jPV��[I����7vj9���r����"y�w��ǤIV��N���-��Ι���� y�����7y�}|܉z(�E��<&���>}���}�Y�Զ�^�^�~��b��G6I�V����;��Сg^�dŗ;�N@�?f��ѷ|��om�ޣ5^��y�~Y0dQu���DQ{f�p���pƸaE-m��X�s[6)l-�mRԺ�1���c2Y�j�bT*�QJі�V�)Db)R��f�M4,m��%�E�j��Gr��X��5���hV�`)]f@[Z��ږ���[Z�1̕�J҅��,fH�����lJ�ڂ�Z�TեL�l`VQ,`cPL����v�&�i���wp�JZ�ժ
[F�­e��ڪ��2
[s.e1��mq*[TF�Ŷ�ml������4[��*�q��R��*���b6��QH�f`��ʭ�+ѥ%�a�GHZ�V�U��b��IY*)�ͺ�	���{ψs�}�������[.C�b�Y�k �^f|�w;���s��6��H�uO4��w�u	�ۨ[��a",�(pL���-�X��6�+k���v��`���P|����=�: z�!�>�3��y��039�[;����P�ݝ�u
/�.[�� 2���=���L4�gw�VF^�gr5���-ԍG\�����y$���A
��K�I5n1|4)�C�!�M����dN�Ѐ�?�� .�6T^��'�����m�m&k#��X�2�p,��6�eoA�8P뽹K��3(��3��ts��
�GE�5�vW�mxf�Y���3N�"Q!�s��e^C����^�T5ن�$�n�e��kC�z`���^cV��L4�)=B�?lj���_,<�j�~�_ϩݍ�U=��9gO=�ˣ�;׹�#���ڭ#$� �P-��τh;J9��-(���l�2p�6�egn�t/Mm��6\-��6�!ۻ
f�0�cB^���贙��^S=�����sr�t>41�r��E����Z��&+')��ၼkn'Y����Ri�2�Ͱ�3��p�7�g&m��4���+:�ܑ�X�|4}�!6[��s��
�iVF\��d{n.�.��8R�;�>fW�m�7k�Sf��X'J��3n=��Y��c��f �����'^�ȟS��^��QJ�uG�x�-��y�`>�!�w �Ο��)y�����Á�17����֤�pV�	�Uks�������pޯ����ӧ=�K�!�M��i����1w��0�G�T�>�
uj�>٣�p��Y=Lٚ���ɫ�����Oݚ�u�fU�w*�K�s�]���Sd՝>����-
��{���� ݤ=�-Z�ȩ��Ԫ�u�I�y����-��u�;�
�C2�L������@!��i�s�rq�l�d�t�g��}�qm$���A� 7`e)\d�{k�F;�iƇ��Q{�bw��#�Æ����x��&˙�^�Mh���BLT���Ķ4&>s�~�)�m��vz���{3�@ƚ�r>�����wјIty{������{ۜ&���u��2��A�q�:�ݑ�����l
��2R�'��z�X�v�Y�]QqztfIp�17Cw�Вq�>O��P׵�/Ln�5�VG�,T��I9��'��{� ��ىW��]:��v#Bӟ.�y�@R��4w�gې/uu�v�	����e�xj�R�f�R�ꩰj�m]����I-����ܳGQ�{�|o�ʌ<��_z�+h��͇�uۂ��i�Y����|��/I�뿞\�R�͉�B�P׎%�-#�lÆ�p�<��ޅ�k��B���ۮZd 󕬔�\Q8�Bӽ�5�oo�呋�-��	��s�Kϩ{ׂi�	��n��� �A4�k��`-7�m��2m^��H9�z��/^�o��s=HЗPw!;�װ"�"���]��R� >����_�߿[z��j6v����i��ة�G��(��{�ߺ�|/���s�H�K��-H\���Y
p��w5�t���0�h�.�.��!�Rl�&�1	�2������f�ϞK�l�p	�;��]e�i�2 ї����+#1kD]GdUZ9rX;G��Xy��x��2p�D����Z��Wk��(�/^��:��g����M�07l=��f�P�!lz/X1�%fz�c��o�=*�(YO>^ـ-�U�3rk���A4�Nwkk�QUҪ�\����iaȍ���NG8	���/��^ʀ2����o�����O�1�Bm̵Ք1�X�m����a��%R�MR}���R'c�__tz���daLή��E�Ol��u�n��i�uy���S�+#�R�����f�bx�DE���z ��*y晡�e�!P�C�j��Q�������J*�Z)���x�z�P�쓡DE���FPM$���^{Or��alG�qW�x�Ed��M��㳺ɛ<y^oR0�܊̃���q���C��܋SN���B��D$��V�MI�,wr�Dj�f n�T���&�����i��������W�������FM����:l�R� $e]�mT�ح��5����N*�C8�DB�V�C�ŭ�u�rl�	�]^��3�D�GJ�EdQ�X�O�¹�1�~Z3��䇢}��x�����{Qu۰uRNd�|� �N!�o�GhM$��YK�2iG��H��䘗��] ����2���i�pm��;�LD��;�я��(��b�ȍ�6;��>{ ��ܨf�-�%��3���H�Hu����
N�;iI��|�ū=�ڳ�K��T�N�#h��l)���B8�C�lLiNb��ʻ��ٙDB����=��-inZ�J ���}*b9��ʼ�}�3LB,u�#�l,]n�j�-r�gu���k�]o���S�����gJ�Tye��%���I'#v���1Q�2t�;���/M�Q&��b�.[�
�u���T�(���>����#t�U�BQ{ǻ����(�  ']�p|�C�OfB��@ȟ��ظ�V�~�E�J =��4�Q_j܍��GEl!<�ˈ5Ee�
���6�#�o����e��n�F��v�cr��	nnv���NI7��x�g�z���^)�;��wpɷC};�{VE[��ֻ����P�57�%5�<f��SX��Rt+���p�zp���yn���=��r��sM�^��f�;_�zpΩ��}�V��t��~�C���3�k:����ޏ'�o-OdWL�����Nx�������ɷ�1U�K�3�k�η�%�l�Q:��4�� ��؛^>3��r=�_OJ>���{G2E�0�Ec]�7�Y���`��ՙ�g@ڊ�J�͕����e^��78�{���2��}矱{W�X|H/��+k(d݋��DM�{�C��֘ka�2���ǲP���診Ǜ��#���3��X	�!�[�L��v0A��d!پ���� ����S.d�����|<��G��_�/<N�Χ͛��}����p�f%SG12TD�X�"���*

��
�2�)AamE�T�j�K�R`5*(V]4DV0(��UV��
5�R�e��:k�\�"#liT�QV���,�V�Rն�Z�Q�Z�F��)��*(��1����4��"�2��ar��"�l��J�v�ĬX1++X,���e��Y���e�m����f8¸(�fS�H�pH�Tf"�-�EE��q�1Y�X��t��@��Rګ��b(�1q�@�,�J�i�4�Eӌ��eV(��LLk1�L�*�YQkl�b3L�ed+��ԊEZыNcBN`/@!�s��?o�q+�6��CA�cf�	q��u��1���K���'n�8�V�� ��/Xd�����l�!l�̝\��O2\��b�N� �vc���7U	cn��h��sM��r�Dq�%�m��
}���eČ��Km JݡJ�ښ)('o9���rs�ѻ#�\:�ǆ"��L�Q�\a�2�	�}.8��c=��N���d�m���+
.�&aݱ���ED�k��4=K+YՎ��9��v�Q.�9M�qá�O�M5��^�1�k)�����p-��݌��"��c�^��%��m�E�	w#=���7r��5kd#�jh�� �7����-�q��SO�����[�nܛ,d5�E�	T��	@ƛV[M�аً,˭�M�]csBb���u[��|�u���S����`Kt���[��+g�٢1�5�	��%�GcW�ٰX�6��x��OR�.yN9,����3y,wet�-x�q�8Z��m����<�Z�\=g�B1�m�;��in#�t�ɵ��JXy����3�8��UUUSEظ�Y�zڱ�b��׵p��z�`���	n��9��t7myL��É�uӐ-��������b����tԘ�٥(r嶲�4� ҝ�u�q�xv!�r�vۓ&��=���O]��i�r7<�%�{7`Ě$�c�<�
f�����N�B�s�[Q	+Њ�U��6ٷCE�s�|���b�X���F�ݶ�&�Emb�����YOu0�$��+�v��f����󈨘�L�Q�O���󼮈�[ҙ�FY�������K���^F�Je|�Q������2�?5���o���i��^���^�(H:l�����v�_܅-��p ��$n��{b���@��ӷ�/�H��ǃ�>���-���
��<$t�rۗ.=�o�@ȟ���8��B��f�=�@Ti&)��mAS����Uhή�PK�q[w�8 ����E���P��ټ�r��8K2UL6��oqd���H��Y�/6���G��F�0�j$ kVQ�9�qs�i���$	v.�iBN���׶�èA դ	f��\/L_�C(�4M��U�9���������O	�����}q/C�̂��l��Y��JMY�vm�}����&�|TW@'Y,#we���λ�q���+t���!y�B�]R����%dA�� ���0LE�^G>�#�h���۬lI���K�WC��^�J��U��q��X���"�!J�r-����s��-v�w��Q��Ygܫ|�|,�l�%T���'���U��3I�I|�A��J��	A����^�2baݛ�� �ç�]��MSb���z8�uqB|�O������@���D��Q��u��p�������9n�W
��4��L�&'f�o[�Y�S-:��.aV�W�\\͟�؍�>�ˆn�v��J���B8�J.1���
#�[�Q1�$�*�5kk;���𻱴 ��J��͝D�?z~��~;�TkKb7}�����{e�N�z�k[�8z4������J4�J�"�/y0t�|�D��[)�l��c�~�ׂ�N!��Tp㗐��Kk�������p����d�(�P!��×o�~n�<�o[@TY(�_#�T�n��O�o��[�
�>�����<�\nڅ2ӻH��@��"��_u{Dq���B�AF��8�$��G&"�����U/0o:eE�^Ӥ%HFi��}�j*&�(�DMR`�w5vԯ�p��9�T��D
��s���}��_W=l�o<D�sq6������ｑK�����jRl�>Ji�C�a�C�L]�V闵�L�;����c�cnxq��H�pf�m��6Y�6�X-ˁ��XC@�Ŧn�<)rL�υ�!�i�n�<�[@�:)�)�=�W>ź����k�;�g7���e/]d�c�KL��{��_}J4�I�>/�y�/9�V���!�A�b��dDû=�-ɫ��g��@Wt���{�?똜ý�h�x`��I����.�� �)����8����7�������-���2z ���ӨAۓ���*�#���7j ��B�yL���@���D
�߈&����8�����C��[�%���fa �	cZ���9c���[!<��w�� ��`�>��B���h ����ɶ1�oE8k�y���d�a]**��{j�tm�JR3�ǹՅ;�~�G�%en��N�K��x���tJ{`O.�uUl��DU�b:Ԇ4� �s��2�]�	��������&���{���²+ �shn$n�쉈�;��3G,e�*��`�����>�h��$���q�t�׫�߀��Sl�qnw<i,�h���X�|���ͻ���	�s�e���g�) ��LUq �V���RR�B�7�s/l2}=W��q�=Uk��e��6�9��gL��h@��_�]��6�G^�:�$�ޘkO�S�>zb�l��o��7
'0�te�(;�);���H ]�Ӝ1Z���u^�X]*��=z�����m�E\B�*�pF��ޕd�U͘���9O�t/NO0����Xr��N,% �Rt��dn��L����m:��x0Ӈ<ER@��d����^��v�.̨�#���N�J�S��A�ڵ��vK����"�u�L=󜋌#�!<��N������\v�:/��m ���&��q1B��׈r�6���tE�hܞ�訷<����]��R�OM�5&�՘ٝ�q�cUY��wt�f��{���5Z�D6��vJb����Z؛��hA���-�z;$�3��N%o�p]��;��L��S �Rp��#0�Є4��a�*�ށ��)m*�l�A���#Ba���]Ě����\͂n��)+f>��ݔa�!ϔ��� ]Ҕ�]q1p�m�-̟���!6��w�&;�sR��ބFo'Ԡ�����'��2UI�p�ّ`�{�D3i��H;�>����_.���6nᦔs��P�q�5ˊò_9�Pfn���"���0"u��!#q0|��A�+��͡0,�:XֳJ�n�[�1v�����鹘T�-�ZX�ݲ1�,9f�.�S�����f���40 V^m��k��sӍm�bku\�b͞����m	L�5ǎ�ʶS���|�r�-�U�[�.99����vQ:�h<ʆފ�_ERD�����{�>�Z.��$}��#��сi�ަ� �f��=r�1����`��ݕ:��p�֊�e��}C�ޭ�u;��}#��<j�s�QO�����R�[@,��{*!x>:��9
���um��(dL �l"6�F����qfGTC`�&�2�Ca,Uے
�n�m��K�&���R�Rgװ�T�ڔ
�D�m�U��m���{��Ge��-W���RP�xO��[:��C��!��_AwC]	h�x�2�q�ѭ���$��M�_j��g��Z$�it`=�#�!��6�"�۾��1
����sy�Ʊ����vu�]�4��)�wcM�R���M�"땓��ĭT?5���rU�PT�$<���޶	�/�j�>��y�5:l����	ciN4�6�M���5�ϰ��cﯟW�;���sb
�i��p���&)q(���U�=�s2�{���
L�
"��#Z1��]�+ŚQ���v#a��b�}�әS��6tL�9�`�z`���P����KOG��j�FG�۹�D�Գ�=�ְץ��Nq\߰��ya�N���D��4�K���d�i����vY�bEБ��g��;�(jNh���̈́{J;��;D�c�����6����Jk8�����w �x�a:��l��jƚ�9���[�E�߽���H����{ -�]=�=�%�EZ��ɒ��{;g^,v�<�TV��kގFM��7r�V?:��ԏ:��R����of����oo9�w�8#����Aʢ�]�V�����>:�i�y���">*��ۯ�t:xxo��.��	6�����w(�dl�{i��1������uΨh�JЦ��Dc�y��n�7rW�3�G{f�h�ΜH��)�:����l�|&s~�(�r39���}�;�L��m�i�ޅ��׸�������K�\ᯧ���v�g��T{��q���"��I͢3hE"�ڡ*噁a�f6��Y��LCchE*TX
E�UwaX�UL�E� �"bX��Z����鐨M�RiQP�,$Sl
�YY1��Cmf�1�`�J,E""���XB�X��BQ�E�*��,R)���"�Q`(,Qt�Z��A`�Ю2�m������,���,��ek�i1L��FڨV�X�V�RE�H(,R�P���2 �)1��P�5AJ�i��B��w��0���2�GD�M��T�c�ę�^}QB��XYV݊6��k�u6C�vYr����"w!VֱnԂA�g�sX�R�^��h{)~iK��j:[vA��˱6ɣ[�sz��/��MY�!����� �sOs�h��i{��lxG�8�j
��Kɸ��:��@�8�{ɓ�B�7us�*QeG�G�y3��;d��?�
P-�7�Fk!��n���1t��"L �����o��]���l�$���QQ�2!�)�^�r�	�)�����N,�U��c��E�ˤ!�x�����s�q!z�������ק�
�}U�B,e`��n.�I�fjͳ�k����5�)	=�U�t�$n�eR�rTz�?�4"�TW�>mU�_Z�GG�=8��v�]��I�݅LO�"��T�cb�Ƙ}	��1�a���#�۳�0�R6L}�n$�_u�����@s�R�p-�`�N�0�fP�P��T����ws3�HR	=��
�[B6���|c5wM�Z��rj�l6��v��^�oD>6����^���T͛*_�e�!��l��N �cp�6Pvv���E��\'o5	�ɘ�׍�y�Fݭ�`�8xH��e�ض��;�M�"h��g��.��8F"�ri�;hA6ݬ�F�r�l�tT%6`�Mn`�I�.VYs�.�nw-��l��GK�1nW|�}�����K�$�LOt/yO2c_ۣ�y^F�f�R��|�Kw�ay�Wsh�[���)F �]z�Ebi\i��1QÙ��*~����Bܔ�;Bzf�FS�|�"��Ov Ξ(��Y�C�w��#6X{<���e@Ӈ�yi���n��W0ɸ�����:�|������BgM�:7M��hT��gs\����sۮ����Z`�4�{wSv��2��ߏ�(�����{͂$��mN@U-���"M�ڕ�8��h4���]�'�ܚ7���k��0㷳�~>�&�!a��{�s|�c��&]�e� =�b>+V��w?3㷥=��*�LCT�]�_�(��-H> �~{%�#;�ݐJ��(����`�>���m�ᮻ�ٯLo��@
��1wse������7����M����Zc�`�N�i����~y7��I�z�Dٜ�:��Vz��`��͂D
��(mݛ�-;I�qG��l ��Lr�^m�렣��ZM�W0*�������q>�kj&�ķu1�K]�O��������w�O��}>~R�#y./n-�<H$g[�7گT\hh�ND��bD�d�ѹ���iڟX:mh����k
�o�:b��^��Հ�<�@-�o�4������������D�6ڃ�F2��WE�Gk^���i��3��`�`�i'lfO��6 �~g�tѠ�ED�ǐ��fOe�4�'>f���E�~�U1=8�2�9���w�n4�,�@=s_Ѳ�75�r4�8"8b%���s��L�QĈ���̟9��wXV�lE��щ��d�1}�n��|�ʏ8pN��?��{d��eݖY =�f����- }����{e�����D�vy-���-.��1Z�CC:Se'�}����TC�3�3�� �t��d�u�UM�*,��5��U�%�}���H:}L@iĀw��Dg|��2�ݸ�9&� :�~eӿy���!�N,�a�e�M��z�hie����h�՝��W�LZ�D9o^� "��u-�����E[�� 7u��;}�)ȅ{<ؙ��j'�эC݋SGi��K���Y�� �{�r�-+)�7�j�{[�%���4��Gpɥ1�]��sz�"ʫ ��c�ikeY����B{]�n:sӹfoI��5&XmP�K�e��m�3�d!==��pf\��ݴѶ�l]�2ݐn���m$k1������7����:�<�:cl����9�6�u�����&O����`��B�Jܺ�Qv�"�`�<
�bA���OwV|M* �/���_ɠ�ܵ��u,��T�$�9s��m����޺�� ]�؃;�L쫚R�$�w�v�X������cOnvDm35�0#L���&�W�u��*M�5@�Zh>/|��Ms��ʾ�F}F�a�6��g�V��8�����9�K��1]�@�8��Ts��Sd�]����C	'Th�$J���s���"#��j��_T#^%�ո0��d�ސ�Rg�_es(��&�2�x@_ca�(	��:��A�FQ*!���O��7/�f�˕�oW�9���dB��]�0�R�Iݤ�#r �j�უUͲ.����T[)x�GO v'-�GKu�U&� //��w݇36���*����8J�#��N���݆KM���G-���6��%n�y�����4q%yDz(�-�]\�T�ȅUo�?�(�wuEgE�ʶ�g$�P4h�Rgۙ1�ٶъ��"O?hf>ZX�hU�܋��b������T�x�Q�FX1�EOO�4��eY툅��\����:��O��e[`-��{�vz�*q$W�V�%OZ:�>ř41���dA��A��f�:���>V(,6��-a����M2MTvS]_}>���c^yߺv�d�a,��ؿE@^;��*����&��Ͷu��yOn"Fw&A�����݋��UsA��!��eY�W&A̝�����#�Xf�ƍE����ut��{�<��6X��i�F�GMFf��3S�{�u�)�U^^B��-�������w��n�⟱��H���n&��\Iˈ��J�bLζO�������9#=-�I����������B�i6Y�Nm-%!s�R�6mV���==�O)����I���lJyB��]|�ۭϕ͍����ǯ��A$��a���^$�b�Ó���&E�1	:��h2&����:v:���m�B��*9yL9o��m�����6�4tJ�y������D�t����XI9�*�$:�eԘ�ݩ��B�fk_���9~�_/��B�ҕ��AT�-$ ���� �~��� �Շ����0�h(f�ί�Xi��X}F��D���;JLa��63Fo�6�@+ @������a>$NR���(|Fk�_��7��|�����@  ~�"��P��~��~Ǐ�~��!��0<C���2q&͇�B>��:4C����y�x��AJN�W�9�����l9�3Aτ  @�؇���?G�'w�BD���� ��� ��XHAad������_����?�	����?��?�����C�?�?)�����H���� @�?���_����$D@�r��$�Ͼ~�А�`Jq��7 �C��lĐ��B��gD7������/���p?W �Jb�"O��a  ��V�<�7�\6��p"`h I k`		�{$���R|�(l>
r������3D>g>^��揃�� �'U��d�?0�C�7�	����A��1���gd�}a�l>��ߤ������g��?����'�ǟ�8�J|�2���,���`~r#��!��?������S���>t�y�P�!��_��}��>��'�M������ ω'�8����Ó�?@  }P>�����A����::�A�'��@����
2�|��   ��� ��O�'`���'�ش��`�Q(|h����p�!�6����d!  }x�,I�0~�H������,6Y6N@I��l~}�i<�Ì�I@@���By�"C$�q,��bKHw9{4u0�����  <���O������C� �3���H��~?T�D�����?�>>g��'�}���>�|�`H~_�>�>R?�~�C�}�?G��O?&�Ą���C_��|C�k�?�X@  }��>{�ϛ� ���ZR����!�� '��q�A�a�!� @;�z����Q��a�!�?o>�:�s fA?�� �`L~���7��x�~�τ8O�C���ڿ��d9'g������C��  3���}o�o��}>�p>W��c��������	��>�C�?w���@(l��>��B$  @��FI�̟���v����s��g�w���B �O��$��'�|���N{�I:�� ~�͜H|��B���H~^�'�9���]��BA��4