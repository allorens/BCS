BZh91AY&SY��CP�4߀@q���'� ����bB�|     7����%�+5��  kMRT-jh2j��5UFB�X��R�՚��$���CUl����$UJѶZ���w1k*ZZ�J@�M4U5���d��ML�R�Y�%��l4%���Vb�ZR�+Y�6Қ�E���cR�KjP����{���L�6�hЩ5Vf�fڤ&�ŕmmTƔm�Q*i��kZU�����T���[Y��M��ͬ"�T����Mk����eR��Ѵj�<  �}H�͜r��Wv�E�.�6�v���5�
�����\	ڂ�:k�Z$;�c�s�WN��6�v���ZĞ�@��b3ceb�Ym���   gw� n;�hУ;�p 5��t �nPP�
\��:��B`  7snv-�hp���㺀��)Ɇ٪f�jщ��4^    �o h((�.� 4�G��� ������h��;�B���wP((��'Z�7���u��s]��� 9�t.�hQ��Yme���jl���h���  �@�ڭ��*��<���5@�sJ����w��R������K����y޽(����@zh*޳{�:=��(B��bl��%��V�2T�h�  ɼ�` ^�ݶ ��]�(Pf�t�()�S��T�Rk�� �Pw*��@W�����*Tp���l4�$*�t�"R���ix  �����%�`wg hU*��`(F�`R����@�g7)J�sF����:kBT��,�J��HkC-���(�Yj�^  3+�h4Ѧʽ��I�n �-�9Ҁ �N�l ]����9�A�:�T``Cwj�� ���fI����j�T��� �@v��  &�n ��P ˫�g\ ('8���+� t69� �g���h��ձ�U��R�j�m  n�=T47.] 쩵��4N��u�\P ;��h ]� �;��� ;�8: Ӛs���F�kV�ZkX��f��FE\  vxV��� Q���5U���5� Wv�� �m� :9ݗ �u9��g8 :�    � @50T�R �  @���)*���&�4bi��F�hO��IR�`      ��$�J��  F  L $��M�S�j��D�4 CA�@h��5$�4j`�=�FF��d��g�
vu��Y�6ܘ�1��m��W�SY��b��f%1x�e/B�E�,��� �]� �����
�x ��G����?�H������T��( ��j��~��PW�������P�+�����>߻���?&P��s~�D���3�3
|aɑ;e�C�D�;`N�ll�� �{e�G��{a<0���l�
��=����{d����=��l�� ��=��l��;e�S��{d�`^�G�Q�������/l�� �½��/S��{`^�G�U�{dOll0l	�"v�'l��
v�����;dN0�l!�v����l!� v����l/�N�C2l��
v����l��(v���l/��D�!�"vʝ�'l	�v��l!�(v��0�l��v����l��"v��'l)�(v�2�l�(vȝ��l��eȝ�'l��*v�̇l��(��=�l��"��/�;a� ;e^���{`^�P银 ;`� ;eG��=2l�����(�l�/l��l L l
�� �(���"�#� �v� �|e ��"�l��l�l�'l*'l �l(�l(�l�'�P�T�T�
)�*�()�"��
���(�"�@�Q�^�P,��S�(���ʊyeC�BaP{`{dE;e;a {e;a;`@{eE{aQ�a	�;dN��D�;aN�S���� ��<e���;eN��"��=��l��
vȞXG�D�0���l��
v����l�� v�C�`;`N����x���v����`(�v�v�b.�$T��%�'[{8q����M�4-)�E[WC��qգ������ݸ*���v�E����^�3��g�V�XN-��gT�,n�U�n� lm:V��%�61�ہY�.Q��h���6c���U�PjG��ӧnQY�����8K�C��"��F�3��q�gk���:��w�\����ا�zdW��.���]\�(���ՠ�����٫�N^���^�O�&9�[�1�\���3��q<g@�9��V�B�={w[����Ï[��s�;w�����Pe7m٧�j����}ۃꃗ�%b�*h�P3�;s��LCE�b�B�h�63������lڌ������X���o0PL�X$�3rG����w9�Gz��[
�Bl�tt�`J�`7�i={~첛{oM�+�Wu�DFK�����H��UmYۢ��<�vi���=Ŭv���Ǳ�[����,�Yo��^�χF���L�[�D�n�JɍZoZSes�$t������M�����.(��1���-��ZwU���V����gA#��R�]�fK�&r�fèayPT�z/Y�lD����7"Ѫ�h�C��Oc���VNks������W伏�ٱ��Zn� �G�$r�{�p���3�ZT��c���U^�S�c�m�u��;:�m�Eخ�c��
sDX%*�j]:)�\�;7J;�>�,Dq�cQb���.�͍��2�(������$��TǙ�nu,���Sɦƅ��ہǆ��w	j)�ĜR:��جu�O`d�m�w�,�J������0�t�n���LS^��+���g5q�޶�ݝ�;��M��+��j��Wv��y"��w���8����5J��]�H'r��7h�r�^6~,M@�֔+1�r��tuf$�v���V[�1��a��V��`;�4��iaI}x��@>/+�`�|�mXV.�6�+p��J�f54�w�sB�^�V<��,e
�ulI_ӆ��V6�fG���	f?��{�tm��kwS�Gv�n�]�����T�1fEu�r�z��*��y� �����0�b-H������lL��}�����7\ױ�7����\��|�mX�L��A���w9�8���ϥ���2�ۃ/0d�Y�xfl����rܛ���Wp���j�A-T&�*R=�S�m2���h����'v�;�n��H��7��mӋLZ��r�5�cڦ�����]G��Ӥj���l��u�W��6�+����*���N;�9sM�6��s]���z���r<������(ò	zQ��u`r��8���H����H G�νTR�:���m�i�{	Dw/u�{�di��/3V�����S��<���>�f�v�.V^�,��nֵ�{c7���}�ꡳ�m��{"+s�δ3�ۉoS�rZ{��Y�I�4�J�{t�yM"�G��=��뻌����+�B�����mS,��^��6����҅��[��
�z��ݸbY,�(ű7W'U��-�v�"���{�YE&�I�����������ю#�eY��{)�]�j�[f�dk *�A��3*��8Q ʴ�k�����C�BA�9�6^���E&�.��U����pnъ�J�����W��������e�yv���a�M@�`��E-�c��(R�H��GdYv�`ӣVT���b@�����6h1���%����F�k\K7��M��U��7_A�dy4�pִ�U�#姻G:� �Sŝ�2�*�[]a����2K̭K-����h���V軂���ٺc�ޔ����MЪ�q�k�֛��L��Q��Na�u,ޘ��#X�Yc0Z�en̛��ػ���w8�2�p��M���k��opF��W��ۛv�r��b�A�S(�6n��v�U��5�7&�+���%n�.~�üe�X}�� r�u+�T��%owU�lV��t�'>�-;�G�[�77U*N�>M���T
y5.Τ"v����f���8�j��kC�5H�HP��d�p�:;��V� ��P{�	�v�rL�*Q��$f��1��\�i9,��j���Ό�{N�A�G./c)��:M&V�D�m�E��V��R�|�B�Hj猕Fo=c6+.�������+�3(.q�\�C�p�X�
`u�SW��ΣVp�3d,	�%��{4V�DM��h��+�K��ѕ�0+n;�7y0��I��2ׯJ��*F�u�����$����ޜꩣ0,�c2*:��5�U��v2����7�ݰ�2X"t�����~���:��&o� ��Oh�q �۫�)+u>Hem�o�qcN�u�G��ؤ�)Z@�
h�{;��\V<K�t� ���)���3�b�����s]��8.<`u2�㝽@1K���m�>O]9)x�޻U!�u:�5�u�:h�L�Ӹ����k�T�g3.d���Ŕh�;�։����3��CGuoO�i�ȣt�j���p�u�O��;�3r�e
�<�����_;״�ʣu����:`������d���ݍ���V��קq<���Ğ�+ܽ���6��l�3]��V�ŝ+��;�f�7�;y����L��B4����+UnK��*�����gd"5�зl"�x
���"v�#�!�0%a�7�0AgqEcu��w0�����n�+#HkXwwp�M:�m=�eژn��,��{�pЄ-��gۆ��"V�j��.ӛgk�m]Wf�#�˶��I���:��<;$��D!ګh��UL��87T܎�종� ���F�����U_�`� j��x>Swr��9[��fҭ!��A[T�,����VYe�H�w,��.�=�s�k�7b���1qdB�Ȗ�����V0\{D=�d�)v�tȐ�4H�C��"��:(�p8��KW5��#$�q�/9�D�y3�q4,V`�]�Z�=m�C��hq�Ä�z�p�Y�Tx;����G�2�o$�.�q�t�*�A�'N�ǏJ6h����u�!����Aͮ�Ϋ}�&�D�!��B�#W'�3��z[�[.$jվ4����Y@��僃ȳV���)XWݍַ�{���ZFpi������G�$79��H��o\�� n�qM��z4L1��z�����Qs�A2�
����hH��ȍw�\�,-�ܵ�������ܷd2k3�մs���th�O#�C�n��]<R��㫰f�N#��=���{�t������O����酫t&l	3�VV��#S�,�?#g-�M�	aoX(�-l
�=H]5&;��Q;�6#�(F8eT�f�U$��G��l2���<d�YVa���H4%c÷�n���1��� l��,�o��9s�4�皩����p�TD�Y:u2"����Y���{v�8�LD���6��)2�5�au�Yԣ��Q��6���{Q����g;R�i�\y��ADS&���U�D/�n������M7�=��c��ߚ�5e�8ҷ)^^�ה���sL�o4�8�}"��t�����u�#�e_]o2~�7�YȎ�I���,�6���!V^�w���o�6�e���G�N�\V�Hc'�������L��.3����/�&n���p�ڛ96H�Hq�$��M���Dͤ��[W�1��E�9'T�I�D谾 �'(�����>��חH��7h�1�]t5+{�>�Wt���sg��]U���9�j�d�m}Ƚ[�JTMJK���7����ݕ�]1v�F�<Y�J'��.<�����2��;�;��"�CJV�ozd�lD:4��S�5�v��MI/hhAv4,jT���dT��ɩ��եM-SQ�%�S�x;f�̘40K�x��p\£�@�;tuf�Ҷ f<+U�LiU������w�Ɋf�Ui�(YijA���Z���ن,�{��m�u	�{�LS��R�W)z��]�ٵOtRL��嶉�W�u��q��TkY��ϧ\vF��՛t�]��-�3F���ui$�5o�w^���Ƕ��E}�rER�0S`�r�l͡�BwT�kf[�a,�%��t�j��vV�#t�VA:�=yi��Z�E�b���
]N�p��z�uЂh�\Pl5�왗���paZ��Z�r���Uf�SU�j�Gu�i�w?��|��J���h�얿��*߶PHa�v��Z�[��^�K?�2�*��k������:�]l�tm�e`؋�{���{`#}%��ڬ�u��x��E�e�32�̓EX��±D`h��h]j(a:i��&L̇K�J�2j�H�92�4�2%�R�W�0-��e�MbK���e��%�B��g(��m#��L���D���5����v�lX&��4)�:�R�	
f��3{�s7Y��ʟ��L�;�$�m[N�81�OY�5V�> ���5�'\�c���O��y��f����,�}y�I'5՝��2���Ұf`��(/Vgv��Z�M��.��֔���~[��ET]�U�Zx�U>v��q�Z��7eA%�2��,��3�Hwb��ݹ��.���#�F�����u�MBܒ���˭��
8XȪ�FF1T(�3o �d���^��K��G�ە�N�^�%��)�s���ti�In_��`h�����Y����Z5l[.oK�LI���Ψ嚴W�9bJvG�|��N��Y�{�d���àņn�̦w�r�.�+���@�sĈ���f���̀a�4��0�ѺM]��aمḏ#Lj�k���xX�g,4;d�1�u\�c�}�U�أ�~2c�v���J;/ ����A�m����Rb�Ep��S����;� �;O��* ju��I4��Kmޣ�pdK:\y�{:�G�F�f��{�V6�4����6ٚ���8�сh�)��$���_J�K�d���K
e-�dv ���%�xw/��e2���|��[������݋7�MQ1�t���e���s��n�GH�`D�Sޛ9��n�,�l�A���{RK[� ��
�� gnN�=`�����Ƽ�j�a�Z�l����^����U��Df��E톉�n<H$M,$���C)V�ܘa{�����Ȩ8,�D��ָ9i�eĹ���c�U��f���Zg˥�P��o:�;�K�Y8r�&��U�ʶj�QdwW��򯆛k[Ǜ���qt�eo:�%������B���Z·xsR��y;�eǔ�&��5�\��qQ�����J���+�Ou۲��`���yt�u٫���պ yI���Z��i��.���Im�5x4����*���QVܽ���o������iA�uw#
?U]l.]u�����R��A������`�6��T�Ud4���"�K���.�o.HX���eTdu�c^��c�;@�R:�Zp`����f�r��>��~({�*߾ځ�79�^r[gk�����֩caxpP�p�|�N�%Vu��(�o�D�Υ�L
�1��2�+v�R��v�f���d���Ƨ�2�4�(�Ev���3�/4���g{�ض$���P��r��j�3.���j�x0�-�@���Ka��c��R܋&*��X�yedޞ�ы��j xy��-�C����["$��t�Ѭ^�Ցm��Y�[s�rH�)]�0⺟I�ivjՍ�x`�Z&��&R��W�q���!�XR:��ڣ���S��S ^��.�\Ur絸�.�H�;4^<*LU��J����H5��r<$�\�8f��������:t��5@�s8�4�6\��DPե��۲��F[;a�J��X�uo.3�-l���)��k���m��[�6�%Rb�O��LX4�Cz��c4�0�CN�&��+/�wH�ռ����x�v-��V��@��-�
��O��8��sZO4��u�����`�rq��v��~��Y��)�x��ugvj9+x��q4���N��s.�:B�e;�#�l"����퉵lDZ6�e�$���[ͤ�'�H��rS7޽g;�6����o=�����&̶���&^�xY�;)�I��6ͺ�0�38��Ҩ�wUõ��*��a�ٵ��x�ȸ� ��;RgK��=���q�5���ųvv�9'wl��Bsd-��]ͦM�󸝱��k��
N�-[�ٯp�-2����,�)�wr�
ίd<q.Q1u�Hh��{��}kZa�,��^��m��u��/I�Y��;6�N��Qa]ݎ��nT�1A�P-%�x^��w3L"$y[.1;Ezx�2��˽;r�)�Հ�;p�^�}wTz:�K�O��lsI�t�	M���[c�5`��s�s��oO,�������Ż�N�kfKF �R��Ab)�k(;�4c8���C����F-;J�fZ������s#�Ӵ��wSa�l+�ee)�ⶈ6�E��wj�dL%`�t8�����1�(v������^.�MJJӋ�kY˱JLiqz^C�w<0�-ϑl�J,�O�K�N������=�I��å��5ϴ�}㬻=$�0ygQdSV9v&�\�YN�m��iFޑ"�L�Jb�J�%`�Y�ZiP9K�P/F��Z���(J�����PO��2F���&a�v����%��mH�D��6�G��],J�;:��2�Vt�,��50�IZE#���H'|C �&�Š�"G��7��]�D��ú�`L�������3ݾv�~R�64��ePƩ�����z�y�C��Ϟ��N���>��h���4�w��T#��e!*�.\�V����J�W!1b�2:7�*ܑ���ѵ�{�ܮ_s�b=V�2�L�{���<�"x��n���:�CC$�Y�};]s��@�C]��gs/��$��w��#�E�.dm���T4#��^]�.DZډcM�G�.9�Ҕ�]D��ɜ"v���a�5��˩&�p�I�����X;��2¬�97�u#F�%w���"�VHKΣF�S5�f���8l��^�ؗLH4Y�%n(���5��4���A�/Ki���8�K�Z�)Oz^;�مS�K������/�њu�K7��nh�{&��ѧ*�rW�40��k�m�����瞛^�]��~��?m�{��2��x�q���3�(�F�=�T��e��g��tb̡J*`@�q[hI�*�����xF;�NsP����ȋ���r!N,���� m˴g\7@ʫ��s`Ar����L ���a�/.AcL���R�tޤ��y,�P����hI��2�^��w&�k��kW�)��/o;�7�{�)B�K���1q�������udܣ�(^�/&���[I�j����\~�Y�3�QУ7O�iQ�qɰ̝��~�U���=7��d����z�6VcZ/8aj�C�f��	wN�λ[�9M������k���λ��K�D-,�ӈ������Y������}�����-���E��Ps��r/_ �X����F9;Fp��!��>(��G��1>�|�|��!���7�'��A�LLqy�Y׍�Z>������b��)zf��~�s�M�j98]���%�_����{y���.Nх�\��T���lⲜ��rh������	�j�+	��OD���+X^q(J��ہ?1���W���+��{;��A�v���|����<�R�{���O<3��)�e�^�p�r�a����S�o�r�wJr�����ŜM�h�|�+���kR��Io;j�Tv��H�t�_a����/�`�m���7\�j͡�
Wf�uK��m�n>���I'�5�w��v����q�\��*�N�)ƌU����:��7%b���V�#TN���� 4nf-jo=�DY|.^1��zF�v����x�n�	`���Al�޵��܆�KXp�N�)7F�L�O[���3����x���]�em�s�39�
�r��#���R�U��hC��)�g��`�k�4����!���Yܞu�0�Yk�kM+�2@���[��]m�#�J@��
��r)\� Y;n����<R鵏a�ά���s��	{��<Cx��s�3���e䖩�X�0���/�'|r���`J��[�]cW�8����FϜ��v����]P�b_
�Ģ+B�+����{qզ,���*kNV��g�^���/z�Dt
��L�	b�P��a��.�h���"��z�[�֧�J3�{w7�y ���=���ڥ\������MPvy��Pk�R0l�f���Tz��3����*Jӈ��d�HM�9�;�2�^����8�)�:�"nUĘ剋|O��rA+j��,'̶�l%(�GBX5�7�)e�;�����om�E.�����Z&=�kySZ��� �Ҕ��Z0���t��;2:�H�\jm�����+NM���;�Wp8r�T��[ȓ�Ε��j��C=1�g}��I��r\�m:�EK2��`K�9�SgiA�����P.�d|��s�.s�PL螴y�Mq�v�g��{W	rnU)f�wF�g����)��}�#ݺ�"9E����(���i�쒕����OgL�0-�,{�I��}�{�牽{���䤙���۫��;�qL��9ml����Y�*pjBT�]�^B�TMsѳ����6��&��ŖU�M��-�m`M��^��|7��������j�G��;�ȷy[�`�Cp<d��$p3%��>�o�N3sd�-��*�[{��3̥Ӿ�&�h#�͝�{}q�G˯¡�%^ݚ�/�H4[<#���׏װ���4�x�xL)�'ZnU���):ܷ�tz�]�+B��
�(�P�ޚ�V�2sVi�+��Z��D5����e�z�F��yJqTn�{����y��!�/z\2y���N���r�ߖ�Uy��M@a5�J�f#���g��.��;�+���<�R�IO(��rX�r�H!ӅXV���x:�Ӽ��j�쫱��8�YXJt0t��vܡß;-�g>�=mo\�pŮVE���cY%asz�m��^�Hظp �����.�6n���^]�JS�t�tnF���Eش��-m������y9�M���}2��¹��]n#����W�e�V`����0��w_��;�[Ö���H�%_?\����T������ݯ�S�i;�s}Z���s���z��˽q�ٸ8��)�flR����/���qj�"�u��b�J����9�OF�z�Km�����=o���xJ:u������=7�.�j���s���{_n���b��"��˩�}�iJ��ǲ+��-\�yew9e�S=�h��b�$}���^f�{ɬ�P�`vU�ks�:�z�ZLd6��*�ob����m�n'~��������;��9��ɱqf��1Ǻ��b�ڼ\��r��X�ȗ��Cv#�� [�_y&k���|^��z{%�x�	�M=�wy�}yn
۪p�.�go6�hշ=���])S�_LxB�m̚����9L
���� �����z��
u�ڬwN��Ӊ�]G�r"N�h���g!A�^i�Éh�]kQ�&^�����%|ze�1��4z�s~��=j�C|/;E��3W����y��6+�h���\R�mЮ�`�kp����{�\kGR����]%�ˁ���Ǽ�S򷼏��_`��߹�||'r�^����T��y��P�ņ�#k	5�VS��YtC�p�g��;.�͑�9��S�أ�0��G{Tv�	g/�|����
]Y�������K�P(S.��wEp�c���֙�w�j�d[(��=y��U�H �8�~�wm������_f�yL��1X���s�C�].WX�'|)>��gI��w�ޫݽ�=7b[O34��t9��3�ғ���zE�bp���c�10�a9�gXyҔ��7�6�=������B����Ʃ���{:��q��M�9H�xo�] ��`��N�xv{ټ�lInXU�d^I���=o��x�⬓س�l>9����ĳ6��9�].�mM��z�g����ŇoF�.�J(V�ee�7V�c��������kK��]��[��d
��J�Xm&��� t-�Y+�g��p,��q���Rm森�9�w��uq�뾫AC��9VY�S'3��A7,6�s��&iy�����uǗ!6�Ui����,�[|@Y��)^�e��L�ɽ�8WN.�6�U��r�b��圛���_��߶~�P�~�%�P5Z6���]JP���r�p1�ڼ;e�����sg\c�\�Okg�5��Z�xU<G�Ȳ��f�fُ1_"9�Ls�U�v��|�8kd7�wx�*����X
F�X%�i��d��mٓ��H�p���iݚ����F��
2�n���O^)ž�A��׵#�	APɐI)�7O-G}Q���]5��Ic	�\�u�M��"�a��!�J���e�o�����G=�<suK^�f/uLp77���0s�! �8B˹R��������_=~��x�`����M��Cv�g���!��62v'�IhY��xQ&e`�m��l�J�a��SK�kF_"���t]�bl���D�e �R�Wu-��dq:#p]�D2X�,AS@r��l-��Z(����b[;�;}fo���}�TV���AF�^�L��Q��\�Ht-�ʦ��mq��H�+}��.dب�{���ۮ���1c\�-b#-���YP�٫h�RG��o�5�%Z�z��.WmF\�qbÊ�[����7��;��%P3n�K�7�sm��=��i��zw����+�������jAt�����~���5�w�T�p��5��<pm�-uMڕǝ���w��5�:��T�֤ �9Y;��hk(��c���[x�)���z�:��$_^P;�� ��V�SJ=��W$*6	�[�0���[�3j)�L��Y��u��ffP��"��f+�v��X�Q�ATz��;�rA��難9����_#&�ud�F�ұX����jtv��9�,ɘ(���|"��2��6������)�{r�����[:u��Sܤ{ɟm�. �|Ƹ°;�p���@VۨޡCF�{eڈ\3e<."��z�����aS�J�ϻ��d�������}� q�3ə��! 0�ɝF�s��(la�t�J�6����K*5J�4�×m��s��ì9N�B�	�Rx��Ҽ��殲]���Ө"Q-�-)��*�]���{��3Ua[q��p*�h4n�g=n苕�6���L+�:$��zmbR�mM���7{#�;��짺�X4wO���f��[��";����v�=�9�K�A!���6���r�H�^>�9��]�{�b:��]��)�����e��/n:>�]�6ȋ��{;��m9nI�w���˲l���q�R>@���9T�쮺#GB"�X�V���[���뇚�:�!�,N7��������ՎP-[b�f3��}�\�s�1,��9�?XQ���w�+��-�";�l����{-��ak�Ƚ�����zŉ�k�a;˸a4�`y}v�gD�%��=ɛI�;�Z�YY �Q��[���鵵s}���y	����4��I���/mTY�*)�v+�;����L�%����,=M��N���T���e��of��4�����g}{�E*���F�O:Pμ5
��Q�[�AH
����t��*�0EJ�v\c����"���.���w!
���S�U���n�,h���>��d
�tk���E��EuA�r�m��	n��9}g72T��0��y �[�d�DI�OQ�=0���uf��)u�7���v�v-0��q	M�z.Xɵ9m.�aG�t�8w;FE�x4}�۱�0}7����!*q��vV:��oI�ssB�|��������\B��G�j����}}�Z����gT��qR�Y���V}�ة��t�K��_�t��Y�=�!h����w*Ie�^���l�SImu<є�u{�%�{m�r��B���P�^��ƲWP��}ʳz�r�}��N�]��3�]!�+�hOU�}fEt�"�m.��Ķ(-C9�;��ty^V�rPQ%.G��ˏ\��3�o��5y8�^T����`�j��l�s˯���=���=��l"�y�gb���ӟ@�u̢�vK�=Gl)�M���)���.�VN�7eq R�G;���[`��a
�.���߆x��`q���S�}+-�+]�ϡ9u�������̜���;��~ŝ�s��;���Sx�w۟q��:󱂦cMw��9�%L�<K9�U�Xg^1��s٠��'pY��DP�U��d�f�[�\�u�����ݚ��i�w��h��4x����v�9	�G�V3+��6�
�A[��v6���<2�ٚ��iP��*�\���D�,�:�Wj�ި��iG�H!���itD��}�
�es�v��mT��o��=���Q���q��ׂ����~;F���y[kB�QWy!����M�y��׉����K�`����g��3'�KRwq�7�gc�l\: SM;u�3D8@ժ	�9'8���� )t8����*�+*�b`V7>�l�9���{���|,��b�\#�pdgb���w������u^��H�L��2�T�٥Eٮ׸l{)������t���
�m[�,�4�,�����uT׼�͙���S�n�*��D��&}�A�T�̫}5WW��]x攷�N�w.c`ʰ��Kr�Х��Vvj6(&C>�X�m.]�H��f�b֏]���7!�Z馳hm[=��\�����8R��S���:^�,c�'0X3���x_g3����*�>C{�{�4�E�>��=�On��[�"F�``=����`ٰhܥ,�+�Z(K�>�h�F�=[�i�v�,���^����]ݔ�מ�[�j3]P�(�g4C*�V�
LPV�z-9tr��gʾI9YlsP��]hIö�=�%9OY���n�vUlm��h�S�٬묌#��,�R�`�G��)�/^�"��L��V�����,R�;����kju��4(^�H�ZC[����mG�&;�|���q�Y�;�㐻ne3�oP���';Ȳۧj��$՗�)ܖ�m�Y���t�Q'�q�]��qj|���x;fi�������mxM;w)̷`�b˙�1uF�U�I��5�oj�E&n�&!]>����ÝJB��>缙7��r=�^�������$w(uǸ�
R� ��n�ЕD�R�|�>���B�C���7BW�udqf��i�b�7�R�wu��c� ]���3��s�sݼ�����I>s}���B3�=kD�Mv�Vʫ�oDǎ���i���?p�e�bڶyy���x��I"n&���N�>x��������U�F1�0��ܮ�������\
��1�oXG�� �?�Q��� �4�u����_r{�y�����)��.�ā�|�O�B��<H�}O#��<ϘE�����y�z޸'����ԣ���=�I�<�������󃄔�ruz��u����u��QE��q���� ����ϯ ���G�"�o���q�Ji-ǭ[�1-m�[E]��z(�z������x澂��<�X3�#oL�<��Q�9]�V��	.�����QZ��G�j$v�Y撷lۙ�pQӰ'��5y�6��G��8�Y���\�yH&���ul�íQ
��U8*,.밯����Wז��-u�Z�`����ye<b�	!�f2ߕ��E ��W�i�: ^4�q��[�oT����+�N�c;{�b�Q�Թ�n#�� {9闗���@r'(�he�.v'�G��S	s�r��L�;c�,1��o���Y0���`��E]Xwkڼ8�V�(�NphͭM9�1v���˞2�$���F�.3nE�o�"��}��St�o/������3b/+�'N�<4�:�*�Vw�yκ⨓e�ڲ�6_�ⶠlX�����{`~�,�C�>�v�;�_t��u���;��N�|>��w/��0��M�^2��L���Z(�/�7s����a�ʇUu�<��.m�h\�e�^��gv�:X,��c=f�7Ԕ�$�/\6s�=�}������s��uP��J+i�����]f`�4���AZlǗv��T���a�\������m�y�����ETdm�%9���s+�����Kw��Qt��o��F!�,�bҔZ���y��:�n��̈���T��\�}�q�4�����y��>�՟LsF��Y'E�/�$�D�x�Q��廧8a�8/x���5.{db�Z��W��jF�����ЍN��g�7�o�Q�PP����L��>����b<�~2�p矸�� �ו}b���L�=y��ڒ��z;f�>cǟ��ʆy�5��Ç�nKb�譝�L�&��@�p�3��ӖԬ<����Cz+�سië^,����%�t�p18%p9]gsK�N<}@��|"����ѧ��B"���i�q�D�,"����^��X��f[�(�`oc��	��[���a�y�-�|�^�2нZ6V�Q`ڰ~��\މL�!�.��4ܖ�z��Q����rx������r���`�Q�͚���">�ݽ8��n���p�H�a�٧�M嘬ݾZ�M�50� �(��	btt�BT$�4w7h���d�]��6�;��浼 �Ee�/&[}0��3fR�8���s�[����O	����}�s��O��퇣�>���w�N��e�ŷ��C��ț.ΐ���l�p�VJ���n�c���ࡻr�����Pɜ�]�A�_GD~}��F��M�����=�����^S�ږ���*O�\{B-��j�1ӟy��MepY�g}�g/K�Z�y�{V������S6�j���l�הkź��T�{jyo�[3ym�,�o���9����w�A���ì�b�$��uWva����2���5�[�Hi/U.��n��̖�N�^��9t:��3� iѴ���A�z�G�j���r_ۧ�a�Y����U�4��6knq�ޯ��[1�oY�7����O�Q<����l@�%�0༝��s�0�:��{����b]æE-�M�-sӔZ���w&k6 &zG!��/w*�սG���#W{*�i]����Z��7�B��N�wZ��`{y�OЕ:���^�p��g(5�2�b�e�ߓwX�^�ʁe�T�6��&���ʼkHe��R�j~A�\,�c���e���R�QZpS��W*�B�ww�0V�����F@���R��e܈o���vǬ�:p׭e�'���l���T�U^�\��އ�S�6(�V.#m�&�� Nu�R}���)Fٹu8,��{�b��0��
w���uX�u=��=�S�����nN{O�w^��N�E�մ{v��W�z����{ým�$�e�=�
�� �z������ ���=Z����VfȲ�^�M�{dݑqJ2�'�4tZ��0�q�Szz���xt;e�srV7T]EW5[��Cһ1/ܬ�^��\Vt�$oM��kx�ono�5�*ꤙ�li{�]tca�nD��;}�;���O�A�����:�:td�̕��u����^%�'x�K�w-)GAא�r�ca�H�+i�ݷ�%��)���)��Lsr��VxC�=7�Y�S�;�����|���r��|�Yv��x&uf��c�:��1v�m]���'jM4uE>Y[}�ۆe���{z��[��~��䦍�/���������Ը��f� ���o5��Q���W�o��[�nm:h^m���3r��q9�V6s.!p�65��(-+k��}3�n�֮S�h������WG������*��e����e⤕�R����x����Sf��&#MM��@�d�qƉ�۽���7�܆�l�w��_>"�')],+�Z�.\�c$E��D��a��ٙ]�k#�շ�dKẅ�����-Ū��2���`��n��u�;Yu���_`�i���.��ư��x��\�҃�wL��[���>j����Lt�a|�ǝ|���!xWa�uw��&�4
u�6�F���]n}0�I���gyg}��B��X�s���V�1w0��4諭+: Ǎ�U�;���k
���������7V��q˾�|n�U]�\ܱ��L����;pzw)���ERT �t��5��?/M\���v��jʼt��U��p�c����/9�8��r)����������$,o��JE]�����+�҂�[m��d՗[qV�ִff��_�����b��.|����g��6�Vh]Ѵ䝖>0f�ۛ\/3E��V���JW��L��p�����s/*���_�.�g{�LQ.��U����=��8��Ž�'V�o.��۳A¡Y�U�v��û�^Q2�禬��vH6�!Fb�P'^�P��aF����.ڱ.N2
��i̸DYK�?��}ɛ��7z++ ��4b7�-z��z��5`��y�s�q�`{���}��:��a�ʻ�ʎi�D�"�!���c~��u؛���6�ȫv£
��y�����80�v�m�힝�my�������.�٨;��n�nHz�x������{�/xOgO���M�<ڝ5HϜK��"8��^�\���N59��0��zۇsy�l�wDE��+�O8�(�����ze*l�.�<��Rܧ�̗��|xm�X�o}|�l{�a��X��k�ئM����3�����10��rB�k��1n���p��rz�>e�����7ǛJ����!z�c=7�yV��|�v��u�w5�6�()�볚(�;�m�~'N�R�~ފl���$n�>��I�'����o�R���3�'e�E�'E#�0Mew�D���Fog�$��kB�k���!ad}��\���7�J��KB�m��m�|�/�sqy�Ю�F����ya��*������C�'����6j���Y���Y/�U.���2��=Rފ�����V�w>嚒J+*=�D _���w���6��*^�p�^|x*8G�&��I ���Q�!q��+h�P{���u�L���I��Y�7���V�Jz�^�})m�]V+���k�:N���JT�B���!�j�RZ�~�K��}Gq0���f���靴�N�@����3y������^Lm7��O	�O�ky�d��w�jՆ!�����d�[hP�.'c��xjt�o��g�zr���uŞ>�3d��=�,'m���))��HT�ݷ�����ڞ�>��\kG	�ۤ�^�����I	Ew��M�{} �cB�O����%�Zw{��H�ޥ՘�3Rt>ƍ�t���Ph'��U90�&u=��t�G�=-��{�=��2[�G����`��m�v�'�#�j�n�G��c;˖Wm(FR�̤]���^�<d�T-J����7��oI"��9Ҭ�ndna+X앖	��Er-���OQ�xR�1�9��~�<���s�.���|_nZoS������9�.�+o��F-�SVX�U�d�2֓R���F]��3C;@���;�D��bw�P�&����԰�#7f�43�e�Uݞ�ޗ����~���h���n�Ǎ�V`��K3�q��x�~�.oH���́O��<��Z�kS_fLQJ��#7��ՙ����k���\R�#���ȰT�~.D�x�������6����qŎt�O"�OI`͈sq��ښ�n=�gwݫI&W-oɻ޲΂_)�ׯ��.�(˽������{M3i�v�k��@�C�X�����J�e�`^Bo��0kXk�X�p2]O]K�,��z�5���3�cy'�q�^D�*��uO�
�D���]A�h�Sx]�U����B3�����4�p�F�p�n3k�9Ͼhc�-u���+ke7���RP�Ũ���9f �Q�̥�F�J������k����X���<�n��f�A�o�u�;հ�����=�[��:[V�J�ۈպ���w=�s}ޜ���z�����y���g��@�g�\�����w_���vN�L�� /=�o�.�Ё���n���oB�8Ut�	��X�5�������� �L<���>�/��q�R�Q��q6U�:ëb皁���[�}���9�u;�ͽ0�U�Oh�.��������m�=�pp,I�$$�zM�ik�<�]�u�*���5�t��5Ã��;r�Pp�������s�~u}.�F�v�t�Ҳu�R�[Xyq��z�g��3��h����&�3[\�;�E�Vc����4-'+`G������_�z�0�Y���%��r�zP:'�&����h�Ǭ�t���X������Ȼ2�Pȯ ������]8���
��-�z�>:����2&��M���u�V�ު�i(��P��ЖwS7�?;�w�N�ʍk�k|��u���\>�%L�wC~;������N���R�y�U�偝�Qd��V����y,��}�e(������q�N��r�z�^n��b+F�����:p�,��Kwa4]��P�,�$;x7	ʰ�ʳT�`��)���u���׏�N�n�6��`mir��rR�;�Od�%�@�ۆ�bC�J��ՓH�o2�١O �2Y��P��7�̋D띻Ap=j�Bf.�ѵ-�7W�����o�����Ec��HW
##���HT��\w��N^{�)�w�J��y��a���=�a^G�|��>�%=*��vM�h��bͯ�/mS7!��|d��rH�	�8����P5�gF�ĕq�8ld�[�ȅ���J5�}]��4�-�N{jLf6gQ/vL�s���xX֭�>��9�O"��V�S�����Ӭ,�l����w�w��<,�c��B���sz�H���R��%�E*m�+��Սv�`�&�E�M_<�loX�j�:$�ԣ�y�S��qq%r.�I�swz�� ��꾮���A��'�sw3��f6e�e�5���r�vx�o����p$�����!��!^)e���~���,�'bZ����񫷽�a�&��'��3n�4�ň��I�Mi	��8�	�]]��:��#�wE쾢�޳���BA'��ɒP}�Uҗ|,I\m��S�9� ��I���եxb�A�ql]�yY���̩oyה� ���������:Jܥ�{b�ܩj]�j���A�8�R�.�~��@����#.�R!���K���U��$��Z�{��8< �5���f�u4`�����y�(`[ſNQ3�Q��vŁ�"�wD!2��P�[�	cǴ���6;W*��=��,n�Ȥ빚��7������MgI##�I�9{V�s����_��`y|���o�������LP�Yp�2��Ƭ�B�Q����/W����f������d~���~��@��ڋ 6ȅp罎n߽H�FZ��l˷|-颣ޜ��2��(�ϻu6հ��+��
Q��PAS���e��
L���gogI6��Z��h�W�8��ݠpGʡW�;/��7|xPZ�� ݻ����>=b⢔)b��M��r������i�8in�N.
i=[�ȹ�iԧV���j��ֲ�����'&��*���pS���:����5�4.c������j��q�Q��{�{���y�>7��Ih1E�-Kʱ����d�
��sSz�\_u���4�6.^T@���gm���#A�P�%\���}ݶ�'6���E�SR�Ȯ�dV�q��\yh�:��2�=i ���������)�J�k$�Sm�N刵���;�C׊���m������\k��%�-�P(1Yx�Q�;t���݈�6���Q�;eY�K3�f�{�d�aV�5B��;�� 1�5�:9K��Zg���kk1zK[���M�G\i��U�̣�1?ufKa%X;�� �ٹ��=a�7ڞ�:G��3ٷ�և\u���p�T���T͇/fڮ�2\σ�"*]���@v�,KSwm��k�����%!���3��Fhw5�@�̇�-˥w)K{�R5okTP
s0�pSt{�34��e��+�a��.՘		�/��K����Rܬw���ј�{�J'hI?3��2��M}��U��Ysk��V�	D���]곫�a�S�N��V����[�⓻���9h{E�f�oVk�T齤,b�9#u�6�N���hт]�$�,)qz���l�J�u2�k�!�ͳI����d$)�{��EŖ���y�crx���y�{��郞Kn>���v���N37�����,�7S%��q��I��S1l��bٹ���pp�����v^��a=l�X�P�"��V��&�f�"��&���)n}�($ $��J�,x��<=��H�anXN�-�޷-�T�R�O��}�w��}>?O���߯��a��C!E����BRq@%%�B2��H�"$lA!GIF���
(�Whm��%2�R"ʑ%a$���(�b!���5I�?FK�D<������N��Y�%�efɿ�.���.�qܴ�k݅��>y�h�&zv%����o�nk��]U< �jJm#�9�|&��#돽:�L�q+�ݗ���,t�[����$���7olډ�f�]�J��3��̈��#���.�>�}��Jc�D���_� q��ާ�W�zDf,.c7E��\�J�}7e��|=ta����!ڥ���ӧ;����S��sY�
��f��g=1ʪ>���v�2�ԏ�3t������xJ쑼��p<��H��v�1+����i����2t�?I�4�ث����*ء9�i�˹��6���D�V#�;�<�Z�t�^z꡿,��p��B��ntD�����y�@78Jr7�Ш��pK�ri��_e摎��a+͵�dx��n5�.Q�N~�^H)vs�tkx&�oG=�}b1S(�4˸C_
!�*�T���2\{��J��*�n��"Ѯ"�κ��.�[�ɳgnO�D�@�{[9i=]�ͦ Nզon/z3o�D���M:��ͮ���	����VU�~��`�3����F'�b�<� S������#�'������F^Z�u�7*My�"�Ǹ�pħd~��u�l\�f^H��U�G5w=��ׂGSfm����J%���~�-o�?f�C=�Mڲ�{��5#ݘ�rm�*l4H�P��e�h�i�
p4$�1Z��D\A��1
aOŸL����cD�i�e�� Xq$B&�
@��B�H"UB�M�e�L��1A��D�p7��#f$T!��0��
F��E��6�l&�q�qE?�(�Y�Q��mcU?W��\S�����S���:�ڶ�q˝X�zj�b(���)�F�9Ziv,�6�j�4:)�����QK5�N �Z� ���RrtM��jh���AC�LZh4�4��ZJ���5�!���Y�������X����堂J(

��Zh&(���lccPQ$�U�UPEQ%RDW1�XbJ5���(fbt:�(�Zt�f	�c�u�UE3� �Er٨��j��๰IPTMSD�6"�9�DӬ�s:�X(�����͊f����Q���֚.X�6�S��QARRQTm���M��T[���AN79�cIA�Q0LTܱLL�TETLQ1MKE2W/
{����HF�d�N"2
R��;=�-��gw�8!\��a�3�{�.�����=2ȼBל���Ϸ�X_!�Njd�IlI�)'6q^ސp�IFT�$H2^����� u@��b"#$1�n�K�=6���%8�*q���y����<����.�ș��˚��8^TF���>��t��/h����>�m �{I3G��ڜ����lN�4km�{�(j���Dj��v(��`���Fm{^8�'�2��&�f62	�����=t;&Ȼ��g�I`���ϡ���{�>��^��sڝ�7���E��'Of�5+���<���j�Y�|�:�`�o,�y4���X���{��s٫gt���DE�������E�Lc�"����陯s�����3yH_��\(�{��>�a^�l�k��=��Up���pyM�����ĭZYȎOE잇7���u�p�}z�ѹ=���P��;:]�hޚ���-�t��gPz��xɳ�s@��Q^5�R3�k���ɽ�����c�|�-�A�q�y{F��O�w���|~�߷.�<��ly�����|Ʀ����¤�}������Y�~���oQ��gK�����^>�k�`ŃL�'���`s�]�Y"eY{Lu���Uy�Er��]�3Y����z��g<���~�X�3�f���T7Du�u|K4��F�ZF��f�iOwu{&��ʷR�*� ��U��T�z7�r����+���W�ޤ�x��a����o�t_횳��7�Z���T�A��#��U��N{Օ%J4�QV�C�������t�v�4g�/{r:��b�3�w�H&n�ot�ޯ	��ig����~K��r�F��u(���}��}>��ꉋ���l�FWa}F̓���]�^��1O*�y� }�^yj�>�;�7|�pֈ���k7�3�&K�ν���)���o���K�Hs�gｶ�Ϯ}T�xz�*��{8��;�㶤��*�:z�⍝c���q��<�����L� �]��/�Q��٥R��kG��:L�tM�?v�M3�	�T�{>k�25������^��k�>�������A�۞]����}z{����&�N�}h�u���\���9�4�.k��ܫ�`ȭ� p&Yskb#��M�9S��.N�1�����c�	��~�G�2|�6�~�A�e��nK�0s�D���9�(�'~���:AP��ߪ��ߖ�v�*]�1���n��`O�S�����
=R��Ffg��p�Dp���O�G�Ͻ��]N��﹨g�����aFo��b�F�f��rd�3����ޛC�G�~y��ߢؽ
ކD���9t^Z������ٿ��C�y�7XC��٤tGs�Ov��0fKE0g1B_	�$�n?����t2�d�{����0��Ծjo�{�ޛvH�N%���ϟ��P�~��yo���/*>����w=w�к���گ�Sչ��X��|ڿE�O[-����u�&Ն,|��;��g�I�Vd�o�����g9�<O�M���ѮRd�����f*��o����7{��\ܡ�~�@eN��:�?��ڨcrVUOo������ƃ�U��=�|�N�8�3�:�[�~���H�7~�T��/���]��FK�kTa�^.��e9o�ן�_-���ycjq��x���vH����~~�?�6H��&�l�Vl.啎���ރ'w?^wh�����s�J��Р�5��/��;�(�e�u�Ǉ�x�<Ғ�W���ؔM�BxX���G�=!�H$���Ùe�4�|������M�\[��9��73�9;z%��k�&�}q�촄�z���3��&�w6��{M~��L�����ߺו������Of�o�d<9��=-��Gm\����{/z��zMz?�%���(8��m�V�������鿹�F��>�n6�dk�hx&�&(��!���8[&9�j+W.�{�xyY9"�FSh�����'y��x쪒���ڻ�s��(�ƕQ>�z
�^�� �ᵮoo�n}<k �D��ѱ�zz�c���7Ֆ�d��$T�y)�<��ɿE��������{�^�6�ǻ��x`�e������������-���]ާ:v9n��3��J{Tܥ�3��*}ut���̒�Yi�Fe�>[q-n6��� ���%��ӴOuW��{��N�m��"FlͰ��՝����vy�T�|Mm��vN���{�FOtl�nw��|���폾�
��i��S�1�v/,D��Jr�˥n�.��w�h�x,��E�2~b�\�}6��u�'n�|7��o{���X���ZF�ʋ��9�Y���nZD<te`��	-���!�{%�J��d��2��!t�o�4�Ҽ��"��.��h����!ȃc+�]V�gD�0bÆFF@kќ`��r�������8�/��22����0�ݾ�Ow�����ʍ�q������m�H��BiQ������U��~�l�)�Ί;���H+bM�(��>���S���*�g�蘪�0<+�W����u�f)�]xuXR�4.ݧ����I6D��tu�����No��䧈;1����]튷��G7&�����+�����s����|t���Z�վ����$V��1[��� �����ENW���#3�>ݍ*�+����=]��i�ϳ�r+ ����΍ ����׽=�n���ڲ��>���I�o^Q��^e9�V� T�$d������4���޽v�l��������Rm��٤1��I����j�2c�bv�u3T���	�b��U޽�<��ǥ���I�d��l9������m��"�ǟG�_�a����n�mpO���0�V��ɾ�� u���=Z����n�t�D]�1�i�y����c-����*Z���¥z������{��1��7�<���Lr82��Wxf��I{��=���?m�A�k-��Fx+ݦK���H�M`귷��x;�z, �L�nL��O=�E�;��l�=��ϼ�y�t�n�������+�r�u�G��Hr/��d�3|ߏ��j�.�B��e�P޻W�~���9����������F�`܃�w�t�Z����\�3'!��k�F�"�=�a�Y�ޏ8�Zv2��C���<�a��C�61X*��dOWe	���=A�=��8� �
�_�RT�{z�3�)sHw5ޙrd~���ʒ��Q��<��Z�@���=�bX��k�S��=�RdRޘ�߹p?7%g�T�T�i�WGKߑ����^O��]�ь� ����f�{�,����)t��o���z��kV�)��:�v���3�s|Hj[��6	k�뉍�z�$Y�7fI�a���8ՕPj���z�����w�)��r�93ߖ��{J%9^�=^����XV�;@�9�#�����e��:&��aʻ8�`��b�/9�0�T�?vG���Yw�l{��s�k;z���#k�˩����
e��O�]C��Юqa	:ꃟ`QIH�Ö��w	��1u8��ڱ��e���+��
��F�ǵ�� �x�&��_�_�Z��9G��fe����)X;�mG��׳�˾�g�It�;n���'��6gE�̠6�Ǧ���1��A"��o�N\�6_3C��89������	��Ǹ�y��C]9��0�R��]곛�W�^���ܛ���+��~j���7����OS>�%*N�@u��Y���������������4Aď��F�<���gy�s|���7�8	��`�������Z\}Y��l�k�S4;^٩��;U��z$���P"e�Yi7�|�Ժׅ�|���I��ۯ9���&o�����"w�ǿE����c�ïxF�M�3=3+��[t�Ծ���9��_�S�i��÷�W�n�/7wq�{�Ϫ��\{]�ʶ_֩ܯL4Zp���Vٹ\�l|�>�gp��=��x�L��rʩϣ���M�LZ�>��t,ݟmAy�T�6���i�m~�S�,���-1k(Ϯbťk�*�ܻ]l����Ȓfa���g�;�=����66�-�+7r�,�i����Aqؽڐ;�����M�X�(T�۔_&	/�h�BCI��&�0a]!�Y{�qd4��:H�>�mR�=��<�59����m�-{�¦�1�������ا@W�Y�}�3�#lwl��ܕ���>ڒ5Ei�u.S���1�Vz�/g���2-8���W��9Shf<���55�DC
�{�4c{t�e�<k=M��� �K�a_�u���+��@]wQtr���o(�
f��J������ި�^�^}�mʪqw
xz����ℽ:�t����S�e����c���5�E̡�Nf��,�A�������K�R#�@m�l�k�w���i�k�{�ι'�,�)nܽ��G�Ϣ��~rDx?M�^�{vI69��l�{��:�:��ל׷�!�~�1��xx\�vb��d\���ڎ3��{�6 �c)�.�M�����ȱӷ�w���7����<�p��:CugZ���e��mˍ�]�S=����{�V,{��d�mc�*	h�[��!��z��ڮ�y��X����uw�49�x���s����;��J��q��cd٢���5�˳|����1����Ҷ05zN�]v�/)fwU�P���O6s��:jWQ9�g2��z������zu~�jcȌ�tE��p���^ރJ�rl�(V�[�����|uȄ��I镾o�~��޿%��m����PQ z��9�|�*���>�a��{gs�у�^����=�Ǵ��ջ��3��S5�;&��di�|�l��2g$vH��6Ga=E�r�����r�}�i��N��lwZ�Wk��k�i|�>V�[h>���n���ZM+�Ƕ���������y留�X��ߊ7�_B�K���M�+/�18[
�_�=�|�e{ާ�}o��8X��+����_�$�����N�{���w�M��('�]��{=X�(�o���yb���Լ
����1��^u]I=����gk�&�+�..sI��z�s��{݆�t���*��X�����N��j�:;"�O38��Mz26[x�OO�������4��7��7��e��듫���B�1��L%r'<��:<�3e��+zH\�����53N� �YS���{O��VD.L��W��a�gV�}��.�����_l����9&r���I�Fqo�T���U�hҺ.4y�.���M-1�㾪�xL���r �|#l��o����0;��~�z~�>c��ߏ������~�U�<
�E�p1��o��7n[�}�r{wпm�'(������zz��}@ݪ�f �k��٫���s�Xݟ%d���'x|��r��W�C�c��0�o1s�_��;=�X�*�)��^��Ͼ��c�zO8�����ac�PU�sw:�9���x{�����2(�OC*���ﵿs�i�̫���f�]�X�	��;�X������g����fA�+,gg�oH��s����o_�a���9{F��'&'Vl�u��bVV?6�}-#��
��j)�pʷR�*�4
�_���ٽ�[ƛ���s�
��N�<p��~n~��+�h7@>���9�����x�����~?Ooooooo��������|�|����^����O��?D5�����m9���4�i�,T���:�H�O�P*�a�k7f�z�|6mGgz���,y�ȴt��n$�;�jZ���ġ|�hR�*���bS���:��v6١��>̱����.���oMשza��p���FN������b��dԻ7f[�)��X�4K4#Ӊ�}��v�"��Jw�kU�y�f5��SR�@.&j����`�+u0�;���w�b9thͶy��[���/+Gnn>(�*���A���(M�+��o`���"�������8S�9�<�=���z�'����3���҄�;��܅c=�z�N|�,�H�d9����G@�U�t^���:��&���9&HKWfq`����QK�:���z�/����!Yk2o)\lC�[�.:�����<��B:r�]�D��{g�U�Y��Leܻ��D�ї�C��h�n���u�伨v���l��|��1�^��:6�mp��2Ցg]�e<�_I/��q~����:�{נ���kJ=q^
n�i�щ�G&��኶9s���@�ٗ\9V�k
����D����Ų�ǣ�W��=]�7����S;�	e@u�2r}��+y0r�Ϋ�Tz��#�95S{
�v㵺N���l���ո�l���L�Y����'k8��;SG*��+8q��[l\=�/�:���s�-�[[��u`X�ҶUn���}v0��*;#�;��¨bn~�Z�<0剈	uT�,�I�����߄�X�g��CQv]�/����ſY��3�^���PZʎ������O�$W���t��R�5���QfTYz��k/2��VPs.r��%��v�GV�X/�iQ�n�k��F��L�A՚�w��}eur^��<=�X|3؈}�����ߨG^c�?\�p�]��6�=���o�ma�0ov�\�Nl/_�!)����/�j�xp��U��4�j�@�Ӭ:ٸ��a{
*�ؾR�FP3��������I�$�㐽wb����4m���'��[��=�
w��~#�6e�������E`�Me�J�V%�8쭢	�"�LVp4�殶!�U��.W+�r�U��P͢�1�GQr���#������ж�[D�ܦ\{�P�����W,�6`�MLE�rl|Ft��&����L@�>l�1-�ӹS�f]�9;giE��(K��^��!�M�L�z�e;��Wn�����oMf���uk�)F�(��,�E�WeR�k0 ���{�2ȵ��J�kDlFimp
��p����5{=u�?{�lT
�ݛ悢�n��	�.4�� {���{�R������0����E������d���_�ګ]D�޻OGM6�PT�K�n��d��Ma��B�L���h��=�hiF�dG���L�YV���]]�UDPEQ!�lDr0m�cDEQP�Ak1EQr�=['\�M��"j$���Y�����Q��DT�TDUVي��Q1DEEUT5DUW1��(����PUD�6�ј�
j�����*�&&�j��Q&
�6�J��A���������MT�-\�yLE�%MW6�&*�(�
�bh�M:"*�"�
h����� �QUͣX�Vኦ*�����a4��h:âb�s9p�tj��cN�\.s��]�N������Z��3�p4p�g�A�6l�N����O"���(�(.c[m����s��f�Q5F��ئ:�]�QMSV���N��r(����4s\卧�s,��W6� �m3��mrpG&�G�j��ѹ�sA������U`��v8�Y�W)���"��j�Fu�*6�E5T��N,�LUQE�E1�͈���1u<�X���8�UP�6
����,j�,r�ͤ�9b	��Ƶb��W1������#���}��~��b�̄?�ϡ���)�fOXt���;��r�`�=��cy@�i��V-�Xs�4
��t�h�.��i��WNGW�x�Ω�D���Q���!��mcxCH�C��M;O����b*�dK;yR9����F�������A�1����T^=��5�p�4o��������%���׳i���+��~6﵍��������� )�C��!:m22�ؚ�O>�@٩*f�eT�q�`&��;�--|��W���&�{+�%G'�=[�������O
���	\�W�o)��W/�{*��<^]=�S������s R�)=�ޝ3����>O��+�?�k�L}���~!�l |�ӵe���vD6�*XM��y��ac'P�p��$���eaQ��~��|njgO����	J�.͍�	W4?wgSɉ�YP
�_[Cy�ˎ��@�Oi��"S��"��e0�nO3c�:��|�Ő��J�c>#���[R8�s<�f�;�A�Gd�#�L8��F�|1�<P����\Ø���j�ɲ��[&]�n4J�{e��<�)����Bm���n���TCt�.����2�K��<��bUX���e;��R�i���t�GPa�H`��}Ü>�2�Ϋ�n�v�� B/��y���8n�CӬ�̹�gS�6��9.��Vẁ����e`�8��dpy���\�*�������|���]�Lk�b�(Mx��e�=d��Nj�Wd$E{B޽ɧ;U%9�d	�;���*��Y%_,���$kw���v��&[.�p�=Dcl�/��'ćA�/^C�k����4b��Ϙ�tf������j�0E^��ۣ'�w>��~�ԥ\��8Y�1�d8-!�[�4ux��������t��R���j{]�BՃ�è�k-{�=>�2�.�ׄT>ɴE�.�]	b���ڛ��c�����[!���mg����~㴓�~Nf�W�"��s�z��[�|��ş�F,��y���3��k;E���X����k%�!���@���@�f ��0]��G0���T݉|W��B�m�ё.���hq�"&
u}R���>��ݛ��<.�@�w�d�×��ٙ)��+n���v�x�e�s�<*9	[��7�شb5Q���+�z�)���'Ml��}��ʍõYa栕�^H�3�Ųѐ-�<���������wlǖ Fs�w	�/�o��ͷ<Ә��e�0�}c��sj������[�Vb?����?e	��3o<PW��+��s���㴌3�Z����^~�c����(�*�
j
�r���8�p[Z�������8]lT�nt���v�:Q�kƭ�價���.���������:�;�խ��v�f4��Eg��	o��y�N�g9X�'̛˱�������{y/h���������X�����`v��w&����΅+�"��P<��;���gWno�m-�=�|<��˙7b0;��r]�Od�殈L�و���J��RS�Sy��r�M�{����0��)`����&�ӭ萄kO���rH�����鮘i�u*L�8LS��{F�q��ԀZٴ��l����]����/A�-��̂�>�!9�sཱྀާV�C�Az8�f�kJ�sLUR��5/wM�.��i[�#h��~g�l����U���_�K�<�߼��)m7ɜ���ERz�
�r�I��M��'��RX��7�<;�@܇Ǘ��d��F�9�\9l��gE�nt9��I��V:����q�+ITXZ��RUְ��u�nkp��0
g[�����,�]�w����-���cO�(LhOO�6�mx�{��4��&�@k���M��=Bu�է;۠2
�[��;s}��G����6'9� 3-�Û�u*��ֽ��f�CˋO0�j)����=u�7\b����A�g��>a�B��{k�L�����t'��Qo�{i�5�
縜G�X]�R�u{���hv}C������L|<Ěy?�F�XE�0����=�^��SLt>�&��8��gH�Y��
e��YSA�!4r�U����E1��e_�5��s����Ň@�_˚`�w���'�O�U��x�6��^�f�k�"�t�)�W�ti��Q�E�m�[�w-��̷<�s��c�0����j�C�,ù���������e�|tE��W�*���f|��_���a��������7Φ���۱�#2 ����J�� y�\e�j1p�)������ջ��,�D3�΋����k���T�5�HZ�]DYB�Rq��Ӎ��(OZ�tv�ëe-o߹�E1��p�k����g�2�/��UR���Bk�R*��B��5��83���r̙�>���=[�S[;Z-�!�&B{+�4��<���Ž���ˎB��7.Hά5�l�v�}@�-�Z�B�F�c�m�'�o��[Rt��z`�Gc@!�4���Ě����~��5L����(�d�ctS*H�aO�|�ݽQ	��_Z��1	��k�=Ʃ��]vNV�틤�n��T;(Á��]0�U(����W��Cqs.@>~���� �j�zC;p�ܺ�n����̀�����YR%/��s��Q�]/Vb��ZPX��0����\8	����]��9%K͐��G�:b΃���vh���`X�ɟ5h%Q��PK��t;��y
�:���Ǫ�H���Y 7�Ch-	ξ0���\1n)n��G�e���ʞ���uUuo��ؐv��H��~@tŔ�G�5�y�?q��B�/g&�K��p=*uk�%ru_u Y��SN���zCA�k\G@^X�s.�p�<�?
T���qF�R?����lKj��7�fV���\�7�{g�`c�f!=;�������'yQ���_�������!۝4��f�z�3l��p�b1�N�����l�����Τ[�xT�eO�\��mrY�{�,7��K�j�`<h�^\DN�ޘ��Z<�MWO{��ڞ^� 3rQ~���!� ��DlZ��GܚT>��:�^{�B�^ϯM�V����p�s��f/_�&��ޭ`���q�s;����?7��p�����8�Yw��J�u�KH�S�^��%��Qx�p�5�p�4m���7�e�-B�3���=3��'9�jK���o�ņ�`�y�cǔ�r��ʆ�u% 3gx�ɽ�kf7i�m��9����sV�ȧ-��_}�V�ht�vx��a�w��p�6���Ko'kr����[�w:�\P:ڼ�5_)������=�v��OV�Ę�|�Lp6<C��;�n�v�m�i�ab��x�((9E��a��$���d�ʿ=��c�W++�?R������Cg����LE���!Of�O9�+��컫�=�([<�/��ء���x�{ä����u�h�SOU��,J��k���g�7	]�/��o3.˧�c`_.u�f[�u�ls��$��wC�a��#s�;y�c��Ʊs.��z`���iO�d�z)�|��Ʃƒ4���㙭�7�h����4r�ш{��62�%,Ƅ�{!�,�'��f�r���St�U���0����;W�;����1L�~�>�����C�	��1��}�<�^��0�7K�����
0{�\=�8�ڂ���+���;^B�f�A�at!�������,=p����Mݪu���:��^/Mh|����(��2l��t��4�Ļ�l`� /��?s�쟍xOP�tިivnt��}�x����oF�ԇMx�6gI�_��6�j��T�el[�0���������>�î��-<3Go5�0,�t�ơ���B��D�Y��9;� ��$��t	�A:�Y�s� �U=Q�s:�������!����9�a^$@:��3�@�r�v��w�L�;ٳ3m.̿0��&S�a�E����&9���wHn~pЊ�3E�92�X������8�ef��Zq�U;�`6�_�R��l'�A���?�__Tö<�Ϗ�w�������:.�����.� �8|�m%���Q<��r�$�Q^u-���f�7<ٌ����=��^�AK}�qM��#�jV>��.s�vu����7[*�i�!Xuj�^��,:���:
t1%�3ic�X���+.��-�3������ j=
���=X�����y��r\T3!Q�ʪ���>�D����7��Z~���x	�ь'��-�{W>�+��m.5�T\�1�66�?v� %�&
+�aMI\���}��� [:~iw�,ޑ��p9�[F3�쵣1y*eg�]O�	as�M�E[P='ְvOi�1���z1���/M�c��
x��U"�����mَ)
^D󌇍�w�nW̛tizaX�8�'X��DJ��ˮ-�Qh�/i�J�m�Y~xsL���	�oA�,�^�I�w%ۄ�J`9��2O��Ju~IP���mq󞨹�ص������d�	�m
�Ӎ萄��K�;�*�6_D7�J�&�{o��!�3-[�r�ɔ��Ɓo\�����F�AƐ!�O���|�%�y�E��Vyz<�BLos�T��Θ�����"�<^2�x�;5������bu�$����D�,�r��tuҸ{[]B���L(�.yj5��܂;P�S���7!���[���<@��	���Ϸ�ȷ!5�z��b������:�ɏ&,��e7�}l���}njp�_��[J!��v�猺��*���Qy6�<o�+���;G�����<v�rf�G����N��v�ء�~����G4.*����N��u��T#)�II�	we��N�^)�O��ݵ�Mכ!�ʺ*>�7��ly3/�L�֎��Mk��}�����On�X4�\���4��`�&�p�����^�4-Z�Z�'�\���K��6
Po����V`V���ͳיakSPw��lDy��69�6'66��ol����u*��ָ55�m-ن����W�����~g�z3g�=�g��`�@=I�}?���	���&D~�}}О?�d��v?t����ᑖ�~>�3��p.CwU�2�'D[qL���˺�h|/���tj��jc�\C��������L� ��!滤��� ��˴��-�UC��~t~��^o���;9G�_��C�}��L��Tw��g��-��Y!
�#^k|�M��.7����m���-u���A�c:�	�zä��4^F�ε�zv�������� ʭe
II��v�lӳ��m������_������߉���<�\���d�f�~"Se�7�T�ðλ� ���J�uo��|��k�~�H5�ni흀�^�Ӊ!�0�^!�݊y����p�������/v�T��I<J~����jT.�g1�_q�=[�Hqm>�� �@Lx�
�y�.����]P��SM)����oȭ½0�`{F	�cK��1���/c�N��U�{�O��W��wr����S�H�yLS�����]����h���%5���`�R
|�����}�>!=�W-PN�R�K���Y�����j[��r��+��BQɳp��T?�{��/�Tb����13L�� �<�K��tS*�F�xP~���xa��+��_�т��o�=��psQܮe�<6�춁�ep'�(�a~�R���L���q~��!�;�
���*�@p*/2�gSs���!��@�!0S �vt�(qU�qWK՘���9b|�L?03jV���v>��'���n��A���¸C��!�����y}��lR��v
ĺ��Q��_۷W���f! +r�-�wK��oy�݁�)��r�Xu�ã�k��vi�\��V�V �L�%3�� I�X�m�qץ�a���/~W�ܳmt[�!�?��0�����&��ݎ����J�!��6�v��sy�	Rei������&g���z���;ᚴD"�m����ǩ�ګ!9-��^����~uCvC6��K���zHz��;D�zG�;>4:�G�s����^z�6*_o۳{H���1��"�"T�}��r�����8���?������i/��{�U����n�]���w*a�\K<{���2;[$�g���5�s�����h�}%�*� �^oJ��8CS�;]f=���V�[�� ���OhY���od���x�g�8�Ѳ��������9m��6}��eY���Y��h��P�~���he=�udފ-AIb؇��JMn�_a�:��vؑq����{/G
���d|�E�,�l���k����\9���{�|�xy�9��Z���u�?���Z] �ڡLX|a�������/8�>X��5IS6��.��������|Ż�\�7/% cj�Gh>lZ}ǫxU�)�08��Ȼ��8g�V7�O����(�3�j�u�"Se�eMV��{�q��ǫz���������Ϻ��b�Ȕ⩦3b�\�?t�v�Tb�j~����I�$f�Z��d�~��|j�Ξi����V�A��VfU��%�q�!J%;6T�a���p�vI������1�_�H�4�������<�׌�\2�Jx�/����(��P�m"�m���d��@�	�4���1���ꖔ�a-!�"�#��I�6[����K!�����������k��v�|��8�s�!��m��F@<�U�۟�7HΛ��k�҃)��,"ї�Ԍ�L'ǘ]vG��>z`xr��_y�����i����ò���c����_BIĒ�%��qxw��6O�?s�2~/����V5]ɥc�57u֡��[R)���հ��d�6�a\���l�����l��������//w�������x�������o�������}[e�J>P��梗�����q���e�l�l�:J�9�ou�y-w���{gz\�Xq���&[[l�kݮ���|�#K(�����nh'�t���)}(�t������]MY��ȵwvƧj�t�_�>kp��KN�B�s�o���*x�_U�6�k��7!ݛ:��y��-�4U+0��-đ�1ͮ���%w�=(R��s�tһL�}���}�i�k#l#:��s�^��z.-� �|LsTA�u��·r�sR�p��(��n��Y���(7n5ZG%5lbk�z_j�u������X�=�|��U�z�ԍ"��!�����k���U��W��9R�ک�w�XG:���HN�9�t�ٹodU�����R�*{WKS�RJ��f�"6�Wu,�D4��IV��;�p�da�G���X�|P�p�+:��ܲ�'nP6Xh�	��M>���G��Jh֏��=�$-+|�"�n�)�_s�1wm�p5ԂM�,�3f�ܓMk��Dv��FH�$�A�f�h��un�wX!�DY{��dR_)(��:W:.;��W��+��ȬCr�:Xѡт��*0g���r�����>,��瞏v;*�{pP���H��f�������d�����w������~�%.�f��f׋�^e�7�$j�c����f�H)��_)[MJ��9���QZ|���}
���;�jd<��_�o8uoe�]ٓ�-�znf%zx�iz|^R��k�L)��׾��a������z3ߍ����S�o��v����>���F����>���Խ}oW�hw(�\��}=ך>�E,���>̓��Ž\�}co�U��UAh��Cד�s�W�g;��"���e],]H+�6 	�l�,Rŏ����8�
�ɖ5��K��*�3��Q�����:��zʦ�Mb��(޵Z��W�v�_#�!)��\� �!��Yi\ p;�f��U�T�ON���k���鳙�Gcۦyz�zm��qg��gG��W��8w�
(�R�����v{�^j1ir����T^=r���dV/
�/�9�ˑ��sL7w�9�ﻔl0�ȷR���˟��,ւ��9w|sm����I�'n[��6���v�taՓ�����1�7\^m8�iWa[�:�̛��==.�=�|_2��\�=�bg����S�5u�ny�e����;�$��1G�,P
���ڠ5mib�߶�y��yi������R�{�^쭻IDǨ��Z*&�p��#SS�P!-��aڵ}��m,��"��][B|����.�S�.HU1�	�ŉ�ھb)�џfSRmn�4�1�p�n^]3e]lL��j}Sh���N�Q�78[����7D��Y>8��)�C�2�H�G��J2u��3���y�:`�`�
�eEn۷/����M��{��C�a���G�I d�F�Qm����<�A[W[4��#�f)�N�u""�*���+��b��IQnc����*)��rh��ih*c�"����\�UA5U�C��E�Q�4�V6���Sx�8�X�
��6Ʃ�8p����QΌQ[l��)��+gDS�����n��PM3u�WX4�\�MI��Xt��6����I֌cTTѮsQ4�li��F�KMP�s���e���TW�����
�1bqTĵQ�ѵ���Y*��f�v����\Ί
��ƍh�D�Er�Q�TV�ETG-T�����Q�9ǁSQQ�EQDEL�E4D�����X�J4��)��:
��tV�UTr5m���F.[m5[:��bNh����h��)�����(����s�	�)�(:�h��(�

)��ib
�#�$���i�Y����h(���U7 �A��r�P��REBUrtUU-QTUD%T�4�EQMRQEU5UM�Q0�T�����מr�����I2�1�	d���f'���xo��}����~���KVI�z��5]eS�x��f쏦l��/	t�˗w��E~��]̻ED�L�8܄&�1�'G � �E�۝n=\:�ni������L<<<��x �:�'.L�ۨ���ܜ�w���� wo�}�N�ۛϽ�E���u�e�OG�{Ƣ��������Ç��g�D�^U�V��L�:mgd֟%ؾwi��;I86s4�� ��`�cL��V���ׇF�d-�;���3�@	��',���ﶤk%}��A�4"�L�vow���u�k0U�ֽ���e��x���:��y����,���![� q����������ж!��l�<B�Pzۆ�rfRƂvvQq�֔� �I�i�ִ�9����{��->f�,�q���%�p56�dj����Ќ��#��zN��2a ����,�����f�2�Ο9���1����O�JI;^K˨������=��=s�
����9�^��A>�zO|��	uc=�|j*.���8h�b��W�5 ̴���3*+\�5N�j���^~�c߸�'V1�Ia,����dO��-�2iۮ���p���RƲ���?j�M||�܈���|��D&I��N���9����8����V�.P�9��Oٶ�'��lt�z�#� ��C-�v��7:@��0����;����Xӧ��/�C&��7����w;9�{�f���M��
�;N���x�؜��h�.���m���h�;bq4 H�˒+<1�
��EʇZ��#��eǠ�ܶV6�[�����|u��Ŷ\�CF�(���� 1#J!J�4�RyJk3Ǥ���������n�I�Ɓ�l�|����a!�B~�1� r[p�3Jfq�m�h��%�o*���)=X� [&�d�n[�#kǧ�l�����=�-z��g����7�&�\Ȇ�u.��T)��x�yk5	<�RX�;P�3��n;ہE��?DZ�F{xtl�-�kmw�xל��Bj�Y�u��*�
���`ں�݇֍��]�^���]�]���C�B\0g��LZ`(Lc�s�;MW���c�}�/�G�BOl��1�N���]�Y޷�\ªD[ �w�pÃ���~A���0��Գ-��,9�J���W[�d�w�oy���2���\��N�����0��X+�z�����!�����2#���t���1f�(T�ڞ�wS4�&�
W����%,˝(���:�ː4�*�,p�OqWo�75ì�[9��5�ry���f/"�y�� ����F]��D[*�xc^���U��W%!�[M��% �̃��oM��cĥC�?gzw�%��F����p�z<��C�^�,�,���~��Mx��,\Eі;���U�K�{n������wa:����x/n��(JT#�}w�P=^��/Q��'tK�j�f�F��q�q(>�*=��//;�,�L�{$�p��Ĉ�ggk�xx����]�|�������r�<�s�"����Q� iQ��ߎ�~�|������Q㑞�����b����q�~�~9����򥭵(�2� N��Z�������1�\����d�-���z�*��3�鱯�`$C��ig(ن��"_��1��H�q�^�/+1��m>="y��N���1Au���4Q����BpX����pm��\k�%��nKN�P�̻�2���ė6L��M^�U�9�^��	��$8���΋,�vC�m,ؙӛ����k@���=�%:��,�ɖ�7����#I��p�Q	�k�r3b4@}�UpM�];;#�7(�`����7OcH��&{"��9T��s�.z����ަ-8_)�rZ�dmM�y��ǉ2^�nt=4X0��"���bݢpУgiC����^����͉Ak��-(M^�v1ym]�̣ud=2����0W��'�6����ؒ�A�����`�F^�C
��m�/SW��T�`�_�+��T>�8�*A����|&����~�٦�bd�2�qmQ�Z��֫�Cd�|;-KOJ粠��uO͠��6�@�t� ���(�����~7��(�pK�*���K�-tw�gjıY����X�˸]����N����p�|��j!n�|�N�^b�y�C�V^���G��_�����s���5�������ɰ}
�^�M,��b=�h9e�$c*�v�Z��˱X� �*.y�*hTP���Q� �l�Uܥdm�k���f�X��1����|d5sؓ3�磹,ƌa���g��W[8��虭Dmb�`��C�~/bv��`3n�J/�Ǥ��D��b� �`uv1u����kIY���,��p}a��\H�Si�^�� �df�0��rC�$@"x�v�)����R���*V˿š���*"���D�ǈ��=2��՟�U���;�i��B^�O�sn%�j�:g�Mr�jy��R*u�<��_�r�����S!�?�R��������fL>��������<��T��͉A�,�`��Gh=f�'�1���N��-�Xt]��9.�Bb����*t����$�I��(Jl�2jF$��`�Fc��^@��t�Sk��Nu�a�nߩ�����߃c�<�; ���a�j~�����:F%��i5����s�:~����=�s���֜\�j���xN͙0�� ��y��xN��1�^�ƀH�kj�HJ0��U��0�fA�^~��=>�_�(f�t��sޘ�˲���0�L��b)9U�c�o�`g)E=8��/>5�W��r/IC���w�t��s�M�^�����.��dF��^`]��GdOS�#D�ߦ��N�(��rf��ҹػ�5%�T�m�;�}�ma�sy`��Q�T��ݰh��q�=��HΡ��{+�����
�a,�b@hۨ3.�V=��U}����F�(b
@��T�@�
DiA��=��lI���}ڣ�ir�KbEY�����L�__#ϳ�lA�@9�Z��ܜk�Ƿ�ϲ�|z��0B+�R�2�y�̷K�ŧ偔�^���:��(��a��#�~kÐ�����m���k��tj��mMy>��Y� kR��E�}jF�����_�I�wm|go
A{����9/7�k��T��f�osk���Rkµ��H�F�Q�I����6�j����Ů�'`�AS;��K�Y훗գT�,���0���ϵ�hZ�(�ë��Ӭ��>���ͣ�3��.��!7�ݨ��nw1�v�*3�~g�!2i����.��{MW�:��N6���0$88�b»3�����#skk嵨;�<3ƈ�v�
H0���d����pȉ��c*ߋa�{����Qx����:g�|���{C�..��~�"L|e��8��}}S��������F7j�k}��SV��fu��%S4a�]���A���h-i��~�����RX<������{�n%U6w+��X�Φ�}F���X`��ˠɒ�!��Fq��gP�Ο�]Ϙ{����^確�K�X^����m�ȱ;���E��fU�8�ge�&H�Eپ��H����o��qh��]�B��<��2�;� /I�z��,�	���������z�E������K�Vf�c�w6�|�q��-!z�-;r�[r��J��hPF�iJ7��=� � ��U��8�9�!���1���U�Ec.r�w��	��	c^7����[�e4�j[moU�^;�Ƕ�k�~�oØ%1rÜ�P�r0o�Jj���OЃ,{b���
W+8�[4S-��Z���g��,`�9��Cj.U�*����Md|�3��G���Ǎ�m2N�O1���6Wq���uF!�hY�TS�����S畃��� �Ƙt���2ۅ�r�7����(F����T2��T��O1W�����q�r�z�[����g�9	�w��){�,Q���.�qN��	e^�5#����1L����8�>�Pmt�T���g���Tg4�V��C��3�yЇ�Ƚ	y�=&D��;I�Q�\��,ܤ�iIc^Gj&wvf��k�h�S3j*���橴����if��@M��ӑ\����f�7�닰J���G1���W�x�%�ܲj����϶��F�_@��:~��1�BcBzG6�i�j��V���_��2w��}r�y�'��k�R��J��\�7�S���3?���p؜��2��m��~O��I��4B�d�qP:w+)���7�
�~�ڍ�i�Z�x�)��4�{:�&�-6t4Ez(?j��Y��m>��/`�\�InT���ZgO�a�V_�
:<Q�9\�v�]���fn��g:{��As���|(V��\��N�ȹ�}aqS��S�*5����ˣx{��D�*1
#J�� �o�0���7���j�5�ʶ�y,bq�*�k�Է5��轆r`C�p04Ba�6ߊ`���ҕk髩ў�mN�O���)[>�,	x.�L�z�3.g�;>�(�,TI�1'����EN�J�Wo>�#�j���K�w��C�,�����_�z�e�oD[*oj0���-�9{�����!@��O���o=�՚y�����=@�C���B����EQM<W^l�����r^?dv�P�E1��[$?|�;�^WU��9R��5o�πV���M��ev�~�WKf���jֆ��p��zq���۬���x��pL&�C��c���NԷ7R���U:��9�������
ObWe1���z����v@�6�C�L�����b�Y�Ό͖R5��2�RZ��)���N���L������i����@E����~�ӗ����<�08����v�t	:,�]'U�~pޛe~IV���qOw0�:�f��]�/J������m��.z�7O�D��#�(�a|�Qu��L��oT\_
�E�K��_�P�r�����:.�iU;^3�x�dc,�V�R��`���v�0��RyZ���:
�3.���ʀ�S;��^׉$���bU�w�w�(ۚ�kɷ�*v~�zK���'�v��z����!�oe��ʊ��'n�+]��_8|�Վ{���]z����2���*4
ЫH��"�
H�B(4 '}z���}�o�^z���׾�$�k�*/��N��	�_�����u��(qG�����]y�WS%n�a��0��-��X��C�A8� v�}��=�d�����Bt	���M�-@;B�N2�ؙ��n uI����U��&
s7�t;�c�m���8qA�,:<A���!g-�^+%��Q�㰥/�-����Z�����A/r��q�&�Y��-��� ��}�iLf,Y��W�}��5��9zn�f��Ͳ�Rci���ϧ^�&g��ܖcF,3�.�$��ψ�j���gc��1^��gv���6�����=������!� ��D[�UOk�֫�tqg��4!Q.�XR��DJ�/cj3],&�ͬa=�HrC�s� 㺃[u���[8������B��"*�D��ZZP�,�l�_xL��zgݿ�	��~�y\���ev����
���of�׹��u�LX|a����ӯ�6��*~�O"�i>x�U�U�~�7�t	*�����ʂ���MI���i�cռ*���h��E��<x[�\!Z�r:�"�sM�K�D5��K</�X�\�~�2���{���/�s:<��m���R?y�M����]Y.���G�b�x���de�۔�w]��m"ؐ�	G���Q�@\�b��a���y/{��g"�=�7����o�s��ڊ�iE)�P
Q
A�i(@
Fy��e~w�����_�Gٗ�;
�uQ;���>�c�E w�}�?��e��1�H�"SgA�h�'��m��f=���|��uPşz��
�8�-y� D���[ �1W3s��o��$�K#(�k�����s}WS�S�]��!���eZ��$�1��9�|G��`�ܹ���D�V�E1����PS��XWm������j��uT���������]�=1����vo2�0wQ���wo��L�=l��:9��}���E���b�ן#ϲE�2��D&����#rk��_OWr2gZT,m�R���,��%��R	u��w ��	=�{�'���qq�vsg�o��'�O�x���{��߷Us]��^j���2��������t�Ļ�{@�ga�Юےzt��]�eWg=�m�yu����
.L��:d�5�����2m��ύL3e�[�6�\�:Nt��[5Ū�L�KA�;�7���ϴ;MW��qg�X�OO���W28�Cr'h[�@��A�^����Բ3����X�����d�^�4���Nf�?�y�������]Lz���S�*� ��U�Q�V{��Jc�u��蠾�)O��@G�zHn�=�*q`�S����:�%�q"���Q�`|�^:���4�5���b�t.Ra��u���mp
V��x�;��k�Z�c����ѷw?��[n������{��!)"TJT��ZT �0�����E���e����W5x�^5���C�*�,`���ؽ��?";�7;8�
3:�x�ٻ�Oöuމ�e��44�0]ă�,���"�{dK��h��	:�����V%�L�.���~@��fY�h�zIv�T� ���2֛�W)i��
I���`_���4�.sk�99~w_�a��;7�퍌W��Y�5x%r�PH�3�l�* [:~
�J��z�ٮ���\�G���`���1��@Gg"��.��t�Z�,i.��;����1[��c��%헮���^�>��͈��*by�F��MB2;s���x�'V.�F5?|�E �9�D͖��BU[
j]��]Qp������?Bn���`��|x����h9Jq�d1���8m��)�%"�U��:q��ȶ�C��|k�H8�F���ϻX�֛ቿ*F0�*�v��o}0�Wԙax	�����W�~D�&F���<93�z�f���G��d.e��)����s="��i�c���q�d]g�Ǉ4�o<����;�?>�#������y{=�/w����{|}��o����������z����G�Q;����u�;�v�E��s93\jM��-O���v/&�wq�棗L�zլ[��/���ѹ��H��#�A��N��oU��p΃��ѳ�rJ�ǯkK�A�o�,���Õ�u=$�er�k��W��鹽P�MہT�0�=��n�otv}��[A�]':���!Y�9����F,�J�>:X���f��wհ;�cn�50�1��
c��ՙ{ܹt�Oh�6��4y�+��U���TOr��܈gr%F8��Uqڱo���lã}ھ�K@�U����_+`)��s�#��7o�6\��rW)e���ν�
'��w�΃����i**�7�-��+�6�Ǯ'ފf����nwt�,��=�F6 vvV+o�L�{(��/��V�:�\<�[��(�#���N�R��õ1���mA�;`9hd��V�].wW�(v�t}b� ��7L�G+3SqC���qӁv�`[ �K�^�����G��T��I�����$ �%u����F�"T`�0�#V�.zJ{珍�� H�kS�$cA��,WX �x 5׹X�o����z]_�*@�6�r�xS�鉑�\�o(kf7�M���Dm�K�n�#v7.ヨ��\ Q�qL>Rބ���}90pN����k$�k��x }��]h6����8KJ�d_Mi3ǭ����c�Z�b�~�j(�s�)a'����A\�з.nU%PBdՃ{�n,ן��	�W�٫���u������ڣ�O��vC{/�����X�]p�J;Ƕh�b���nm��f�J�������t9��X��K��m����%�="� �/�/!��o�{_�N�U)&LbA�,�j���Tn�͐5E7��5�9��CU�!ݜ�F�i���R;N��ak:m���@.j��&��6Wpfg7�^�Wv�0�|�n�ׂi789�t�/�J�������I���`�g��k8�?�/:ߛ�7/<x��P�>��t��n��U��Ĳ�:������NCsMh�Bˋ~.rxB��8Z�a��96�Xnh� �>��p����<f�b��-gt�0��l�й��e2ND뗪[�x��y[2�{so�pcJm�c�>�4�ƨ�v���o���0
��)�cc��Y�n<��i�h^��cPT4,��X7�V&� �u��+/Ou�OR�Rj���uɒL�vT��f]S���q��c��s�]J�����,�/��j����e�n+��=�d�4�͡G78�Y�ȡ��0M�U	b�M�ciPK#���\�A�0A����t�gl���򥒩f�M}ko�ջ8J�$����u�r�+kW���tg
Đ8]fdN�&p�N�L���;i���&C�E'Q�����E���s���{��U�����b���3�S�`�j]u`�q[�ڦ��u���)9�\ ��N�����UFڊ)�J
�)j""�$(��*���i�j� ��* ��)�j�(j��%�h)%��"&�*(J
B�(��"JJi��f�i����"
Jbb����)��f��&X�����y�����("j���h�4SAHDm�H��f�i��B�"��""��X���*m�4lb"��h*��"j��������h��X�����"d��H�����h-:(i
�JJ�b��J�����(Bf�i������"��*�����i�(��*������� (��!�J

��h
(I*����j���bZ�&��
�������(����J
��$�����&���y:J=�Ǟ�ߋ�}tu���΁�N��n]��t߁��W4�f�U��=P[H/xءF�:w"<:���m2,{��7�Ͼ����]\���ܪiU�ZEb�B ��@�����(s�����^9���4(���x����nRy����`�X���ĭ�+����n��8|c,7O�n/�δ�o�$닰J���̦��܎�m./Ϛ�p��a��=�}`�� ��,[�D	�tm��^7>hW���{S餝���̓d�L-��~*��|���4��a.�sp_�~����=�,�n�F�����#Fn����/�̋e�PV���=��h��֠z����ȗx�`>�Lы.�;aQ]��7�>�-��&]�9�n�E�a�&��c�@��T1��׃�[9y�חr�N�hc	�[��۱���6Ev�j|��.a�gu��~
W��=��F]���V�4��*Z��s6�՚���l�y��W�0<���ħx��m�Hxn� �W �6��>�Yk�����k��T�ً�T:)�0Ao��8�sE�
�Ʈ�9R��5)_��t6�;�OE�ڧ+sTW,Ȭ�[eQ��쌸�P�E1�8������� ��f̈*(�L.bb���Xܷ��+c� �::�B����U%:eu��A�^�냝���Ǥ���j��W��0��x0�ɓ ך/��*˹����^4qɣ9Kͨb�K�wNRn���;�L��Q���ɱ����E��Q����"�q|l5�7hE�����ya��i"U	�i�	%A�o���ϯ�����}r�߂�%6_���P��R{���`��4��KS;Z-�'C���k��;i��.�sO�d�j~"S �Jt�	��U}���}Ǆ�-����'�bsp�������k�Иsϻ�k��2���wΓ�^Z��,^��n1*�S���vo������'��N͗�.xb�ݍ"Wd��F��]0��x����5�;�v�~����2˻o�ϵ�-$�����IBt�p?�W�n�vNʇ�⮗��,��x��SV�Z���ʋ�$���]&��q.ka�3���F���l�/�z��Y�V�s�]��ձ�fsr�/_R�-Gs�U#��,�� �;��7 8�!G@G?��vV{L'�Y?k��W�ǫ�V5^��S���\�⠗���o���N�;!t�+�0��3�}�1k6suyt!۝6C�n>nt�/�*�<u>X&} k�&g����i�ؓۘ\*ew�շ��D3$2�u�p�����m�_�?���H�t��0�,a��u��Iʗl��v�.�j��\2�9f�ˠid����/�4����M|���S�?97.O߯e�����r���ӹA�^���%�����;�-��f���.�ɋW=
9��K�n�K�2d�5%��7mg��
�@���
��R�H�(
ȉ2��OϞ}u׿�9�>�����1o��;�:a��Se�����[�4�ͬa��Ԯ�q�h^����N�,!������k�ë�8W��f�|1��՟�]b�ou��9<f��U���)����K+�\��z��S���9Iw ^ͧ�xkזx��Q#��R����b*��ʉ[���.���P%*f� �ʀY8�5y#��gױ���N�כy�:�ʄ�Rd���Z��bZ 3��u�&��4ߧb�#�	M�aLm��%t�A��7��I����Þ���zX�5iJ���`l�as;��ղ|SͯЂq^��=���+�i5��SC��Y��r�jܾ����[�:zkw�H�*$�r��c�+>"�i��vN��?��.n'B���"KY�t��3m��,V�k+��6��p� �&�}	�>��.�vA�l����6Mi��5�`*Vc뼗�t�5ኹ�1/E��ϚE����!�m����8�i����7;o�u��5S�7��I�M��8ŧ�]o<A���"4c�}j W�yR_j>��f������9=/x��v�s��P�F&��AB����
<ȳďE�kw5����K��iQi�H��1˦�
a��N�<
x+�����_�[����n��^�@�9C�6�Jͼ�+���4谂o�L��9��҃�	@"B�R���V�� ( �i(�=�z3���As"9��Kj}���:��h��l��BԍeA(�t��;LK�k�9���~eP�y/n���Þ���ޣ��Ҏ�<��	bA�Y�|�2��Z`�Ҩ��l��e���^�>R��v���� ��S �0,#��򶎯��#�w�i�jL8��,}'��`���7��Nn:��m����b��A��j ��5�9U�>���"�C֚�AŞ���2M��hw3ٳ�ϙ"D���@yp�����43�)��^������jFkI��E^�l�VS6gH�������SIڡ�Z��w�U���)��"O��,�e<z���{e�;�������~��>����k�Iv�T� ��˵��'�sͼ�.�:n5S�3�Һ6n��ݣ�BRXC�[�髟*݉Ơ,�A�jd��A�#8�C6q�^d}l��Ye�[`�ߐ��yiw^�`d�������#��X�A	��� �ӈb�-�9�$�] �*��vb�tc1�P��.3��\؉.2�1<�:�Y3�}~�c��x�����%��*�G°s,�Z4z�'Pٓ6���}�#е�qUq�nQ���.��n��1G� Ә�|Os��Kڪ`oq�ΝC�x��|���&s<?��I���Z�׽��l$�'k8K���͔;c��>��o�B�H��)D
U�Xb�{��������u�e��>����Y�F�QaMK�q�����\c<	[�f�	;#r]�\�C�ҍ�C���3��/�*�(�˝;�u�$�Z�TS����;���8<���Q�OvS^����Ngo��v�����n���F�"���Rz+�pf˳e=ˇ������ۦ�GF,��C��P��z`h/=�%�{��4�T��c��"� c�B�x6�ҹ1����>�*���9�R�ڛ뚥ל?7	=�r��^S�ul�¨��-^�޹I�Ғ�����XҬ��|+���~d|&�,o��A����� ����u`���cߌI�`�E�,a|̚3^*����[hOh���R�֑�NV�z���!i⇗�rzG6Ф�j퍡]���b�����Gj�q��J�I�zc*9�����t����<5��π^%}��J�Fk�6�g����	��T�?Mk�v��R����0���dȗx��e�-� �Qp�ݜ��'�.`����r]���;����Q`K�v�8�����̻Ls�[9~�u��2j��{ɹYp����g-��a9�	Ln�Ěnr�q"��o��e�ݡ�6Gn�-��{�Wc��Q���[5P���m�>��M琟�����`�(0���,��ם5�z���VN��5s ��l��3Sh�ŮCu���m��^|t}ȏ��Z(�i��xx3���3x{��u߭$�*��":
��@�,"�˘}����߂�;��G�`+�ɗm�5���\)g�ޗ�����!t�n�3�y�W�b|���ߦ��x��7c1�>h����¶�/F��a��-�#�<�!�{�ך���^:=5������a}�w+�-��(�\��I��x��������;)Β�j�P���p��l:�*׶)��9g`���fX�DVVn:8���$Աj�%6_�HL�ZT+�������M�CZfR���y�ڢ��Xsb2Z���˨3zy���`������f(G1��N��I`��B�b�;\�;}~Y���8��k����.�pZ=θ>C���hH� W��u��K$�s�.�H�a��fw]>.݊���ۘ�\ �s���B�l�D&���(��<�L7ܪQuvY��U�z����z��xf�C"�\���ׇM(fƑ!7C�ݝ����P⭃cv�S��n��Gg7S����ش��T4�L?5y8������G�M�1�5����.��=�l8�(7��K.K�9��z��Q�}/zwg>{.G�j)_�z����G����b[ꡊi�V����kT۳��y]33!�E�����?���������4˾�:{F��ۓ�;�;�h��2iC��I�wydo�_Ap�/�+����}���قR�ih%JQ� �f�P�x���׿~z��}}^>Lz��L-�:���dˑj;�<��>l/al_��B!B�ҋ��A�FǊD]����Ӽ���=!&i�X���Ԫ��J��+[������;�A}C� �Χ��7NC��-[Lzv �p��vd�d�6����WRca<u>?�^�z�3<��{%����S\d"r�^���P�~�	\9���(�����?.��;d�1�Ǥ��p@;�U���Yٱhs������Ų��� K��h|.'�*l����t�94�ΰ�>R��e�v8�j��ٌՄ:!D��;O��k����]X�_���?��ʇS�{6�F6���j��á���"Y�3E�L�������O��o:����O52	飘��$�5~{�ܦ8��F 2ߐ��Iz��WVq���{2>Y8�5$v��l�z�=[®�N�G
�j�fk���w�]���s�%�!��D\ztW�V0*�b�>�Jl�2j]]	]8Fc��%Q�r2Q͞xui��]~w��@���" V�#cs7:	Ɓ�%�r��%��ǧXZ����3b�6�4��݋<i�Y�"���;�wr�ݐ�ڞ7�fi�u�h����'3��P��΋0��3�cBG�٤�L�m�V�w\� wCus)�]2Q�8�F��j�Kj�>j���e��<�r���NU��}帣��ew�KvlƏzuC<����C�J�i���i���VdtR���5�ݽ��^���=���]�*a0R;A�y����sMF9��U[S�����T�n�k�f�d�qS_r���2l��Н������'H���p�ւ�6t�W.���"��I�WU�9�����`��a�@o4yȄ�m:��;6�̧oeF�.���{vKR{T�I�M��^��!<�^��Ժi����-�ڲ�ZZ�d'rvq�z�����dĶ��VM7_�Ms]����Z�����A�� *g�md���{�}��u*���+� E��2/p쟕OW�s��E1�&����I�XZd���+�6-�H5�`�=NK�{�?M�6�'�ZD���)��ݛ]�:�����hZN��ø�e�e��Mz���=ק݋ʢ���A���lC�.���ǋ��S0���K�rz5����tϰ��>�J۹QpQu4�&+��~���$�L�,`�������=��FTv�cuS�N��BZ����-�B(���z�;��hU�r���`�?����C�~��?ؗ~K{O_��"8���Q�)����J|FW�W��u�����hMwQו��&��������z��y'zh�Z5�z0�^�,�ZMk�Jg
�Dvsr�V���V���n��y)��v�A9������֏��_d~�H��DB�>�f�8����w`ڡ�&7lmN6۬�Fe�f��t��@��A�F]���>y���P۵T-��ڌ�+�R�
ȼf�O�#�����Z՝	�0�&�%r�P	�s���X������7U�)nW�� '�{��2Dc�����¢nA79�^]���`=k����K�#���m�5�r��z
;%�e�J�|��a�(!�`ߦ��<k�=5�&v��<f93W����kw�0��'V%B�ʢ��'����\c<�-���$�S�D�5�k��&׽�#����)�7:d���rOH��QN.����V_���c�YvC3��s�̠��\�Hp���ݗ�7:a���e�/1V�"��q�n�zw�x`�=oUWggp�b4X|e�~��G<��ʻCH�%=_�E��Aj�瑪P�ʮn*��|[�{�tV��UN�������8Z�!�n�/%���4(�;I�>�^��W8�y\4RFz��VP�'cb������ȃ���D���OB�qz�\��H��1'\^yǴE	���(�N�12�D�k�i|�b0;
�޺���`�9���+Va�ZˈZ`�+�~ ����ϷN����L.\�sM�����1�y�U�Dg�oWO/^�=���ʒpWun�_c�e���'\"�PL��(�����-λ[��M��xx�z�,��~Ě�0��-���<���\��
OO�-=��_����%Ăݸ�!�A�����}��71+\+�W=����*9���:�9�;�8"�?į��_�^[�Va��>�6��"�zQ���Y���,9��T�������F����<����`hT�K����a̚��gv7d�A����+ubr]��¿wK7I�1%ډ�c�@��i �b`�m�=ս�S��B���F8��#9ݡ>0��s��t��d<�t�C�Pi���C���y��T�<2�{�ӷPzb��&�k�k�2�.2}��Ƕ���3 ��ذ]�wJ,M7b���[�7��,���5曌�F�Gm}@s����C����fU�uO�jg��͸�#��`>��^S�ML�^��A�z�P���p�7�H���:��hBll�1��V38�d��%�Jn���%0����D���!2�iP����
��U�`�e�ק{�F�U��[�)[C� ��^!�sk���x���RX&�EP�����!�������}�^�G����{��>�w�������~���_�<uw��f�u��9(; ��õf��t$��숩�[�7'�f�/0KT3�m���Bu]�p�i�2��E�D�P�]6�FI\���囄���í��{n2������N��ಟny�m��[٢KbGpe|y.�rǮn8��8Zr#yF���6�@�`��/6�K��_eذ^.�:�gj�j�TA��A
kY�2�ʾ���38
Um���s�]��,���kb�=���o�J�Y�V�{��Tpι6d�5��'{�O��3��\|r�9-��M��Vw*�1N�'^ь2�K���ǉ���G�إ&�^Ԥd�*�e�����g cj1�N{��L�Mt�-;`w
$^��
�B�h�;\�]�K�p��\���KE�M8�E�N���U@Y�̧B��w����t���YO�,7��'�V#ٛ����4�I�l�����-Y�w6�Fl,`uO�I[�q#yݰ�&Q�'�H#X��[L��T�m��Q]��X��<ۄ��z��TYTL�����8Í㦩�egX<�M��-o
x+7�Bh}F�҆M����#�>���]T��4���3���۶3rS�(��+���ʒK��|���_*ԡ��v�Lʵlj鑭0ޥ��Q�r毁f���gQ1���g	�Ę�
�j��[�s��� Q�����M�u��_��lw�M�A���.��+��]��r��8�zx\C@��0FF�e�{ٿ��~J�<�d���g��ɻ��{�T:����r�����1�˸/y��M���9�4Lt�A�R��*1���^��h�G������V�x*��s�����-��N�6���~�&���ֺ1"+��=��}y44+�r��˽e�:��el�ˏ���@;O{�*�����NkklA�P�%�vރ(��;8�I����7���ExeS�>v���6ޫ����}Pw�E:�{�����F_�]��}ld�Yg;j�(h���$��H��B�f%gh�%i�y�,�-T�(�ɐ�ݵ�+6KS��Z�����-Ν�ؖqR�0ň;���LC���)~��>+]r-o��q�{ֶ�9ϵf��7���ܵ�m�㴺����lCۺ���5��9�ءG/+�<�Ӯ�Zc^���1�H6lQ��݊��u�ۛ��@!��;�K�V��>t�ec԰͑�r٥(����~{,��g��3p"��/��9d-\2���|Fq%�)��S}(������j&»D�f
9��U�\a.lO!�޹q�T�ϖN]��{e���v��xo���3x4�ٮU�>Xuu0!Et�6��@2�6��ϵa�	��s���% 뭮�����䴱w��d
�9q�d�o]�3��{:���A|$��.`I�s���Kgb��Aj �3/ubNns5ذjr������7������|���������"��(��Zj"�ђj���"���J���B����*"hi�`�������(`��X������)$����������� �"������(a;�E5CSQ@TETEHQAALAMR���RDPSEDDP���U,��RU4�KEADT�QR�4U%CT!MU4%!D�DU1MQL�QT�Q2�PRROvB��Z�**
b�>l��0QAT�HD��M4D�EAQR��Д4!�Q@TE���T40�AJEE4E��U%5S3DQ5HDJU�ID^KR�)CQ,q���^M���n��2~��
I��~[���U�Ȯ��ЎQ���A]��d��ٔM�)d��<�}�.M�tK�n��xC��1�խ�e�$��r$�\F$*2�N���%
L6PI��Q����u\��7WW4O�/�"|{�ߨ�6��C��F4DN+׍�/��:�xcO:��O���>�5��):��,���v�I���^ȿ3�hb�e>�2N�.�*�>Wq���.;C�N���r��x�0!uɇ�Ȣ��;E�����j�FZ}ҷ\���sfQ�NZ���k�ji��#�&�`&��4(�T^�k�(6v5��6��P���L����X	AcK���PN%�;`>�a�2mj�p�n7�dA<�ϙ���k����T�/6���ܺ��F^���u6��z��ť������G00��������&vݷ6�����sBri��	�-l�J�aA��S��.�����m��`��0$�a�/:�v�w)sUx~
aP_b���q�;��:Y�ߕ&7����`����զ��򸪊����o2�1^����f�; �>���Ѿ�w��.���ݐͽ�����/�S��O{����"r����I(�!�""+Y6+�b]�1aCC�q1)�6^����g��Ŧa��Ӆ�s�+2��،�l!��t= �˶�-�;P�^�Aiidv�IϘz����]^�U~�wP3�)�I���o��۾�҈]����`SJq`�r�jp���>��'���,���y�Ɍ��Z�WY��y3�H�L+�D������A�[�,u��;y)o�RE���n݊E���:wz�nn���yQqDw��y�Y����[~Hi���ϊ��k�0���O}�&����h�}%��U�C�~H-��U�Zf~�
�������Ʒ�G`�o���_�(�W��v��}��3m��ʂ��	�#��l�|i���ԉ{�=+�A��%���t88֋KϢ���%V0J��W���׼eM@Z3I�J��[-W��z�tFT��v�����Bޭ�[� `f�~��հ��\���A8�1,����Mpӷ�Gˣ�/J�Mw��Ưs�:zkw�H1>l�]��L&
{A;$��6O#�SH�?tda�}�@�J�w��R1��Mf��ic����d�_|�܏��t�������Z�m�ó(`�zT8�z�$�b)9X�"�U�9�^�#ϳ�aA���oc��r;�	�=��B-��HܔԞ��0�rt�q�O��%���i������n7�y2�j&���G>�37����GLK~��n�ګ����ͨ��J;����3��e��/Cu�v�~6{5C�}�ga�+�y�o��	����Ԋc^2k����\����2|s�<n{c��3�xd�+��S����c�U,j�Au���'�f][��������d�����@m����-0���#i�u���������������H�����9_ֹ�rH'ovw�xX�'�ǝc��n����w0K�򥄛/X��K-�?��2�a��.7}�qR�e�ݛs��!���  ���Γ�����V�S���R��	�Mk�-�� O�����?yu�����+B������j>�N�_[]�ҳb����\d�y9�a^$@:K�1m��$��Ƈ����k�~oΩ�KRZ�_]�S�Lc����|w&$�i2�ZG.��z/��x;꣭Ov(ȫr�U5�ں�u�c����l[<:/��8�ns�}2�3Gt�TS�ܫơ�_Z��ؖ!K8Ӽ�1�s�6���r�\�w�p0&�HN0l|dkт�gջ����P�qB� Ũ���.������ݶܾY]����-���r���C�Z�`ғ�[���.��,�����Mp�D�TO.����\ps�[h��g���YQp歂P���ÞC|���o�'��+���,Ӟf�á�yW;C��O8�/b5�JĪ,)�.�Ơ��d:̍g�L�Y���5����Iz�wcUn���Wn��!;�[��~��=��Ju~HеbU��:q�c�BΕ�7�z�D{���e1�Qz�bBt�x�µ򐠋�����s`�b�l+�������B�]�уNu���6r��V����t�[w��c���[��q5n������n���
w��\�jWVpi�˪h QۖK��9屾�F�(t�n]�i�醑�J�"���Rz�\h�6^��ק*�rg�<���%p `B1�t�z`��s��,���4������6Ⱥ��7&:���MS�����G�܎1����;F���u��!�z��Q�:�
6v�
�����cz�[���泝m�_����Lkq�`�I�K�b��Xv�=�ι}c�t,�n�F���X�q�#�l��D_���<>��'��v���, ����mnk&*e���21�B㻥�V�mH"M��1+\rn����=4X z��V���~'~�Ϫx��WJ��8�����a~�eK6��������V�k��z�hj[���^��g7t2�L�C����U9Qo{��DS�C`<z�&��d;��f��ۖ	�.��1��f]�/1���qW6�4C�����8�~\Z_��H4<���(l���wBGȲ�C�A!�	׹]��Uڍr��pd
�v��-����U��>B,�����5�t�~�\'�_�|?����Е��?�/�8���������7��[��.��CpL啨��ϱ���V
���f�m�U��o�θ�R��Ɛ������QCi���_LE�\��{�u�C{���*$Iy7�jR o,����!b�T�)�Ř�Jŗ|�Slر��[�.,]�R�Z���¥�"#'e4�uST"a߯������@��r5曌����_P�E1�������#���pV�O3c���Az�:.3����C��P�R��*B׿�U��Jң�z-�\�1��g�!	���s���LݷDm��m�P�-�E��wX��njJl��BeV�
O�Ei�sn�z��������SO�T�l��2����	�H���أ�_����x���RX&����ʸ@�qE�Z��vw���~׆�)ZO�|{�]��)hpco��ݓ�D��&��`֮�l�����{k����
Wq�W�Ky������>�v�l�^����8L�!z�����5U����{��2���L2 ����l$D3��'���F><��v�������͆��B�<��Ê���^�ŧ洠��.��@'����L6�&�B�d����q�P��ָ�r���jNл%Q��Q�H]�C�c�T�cq��IWy�K�,����; )a��8t�<l
���%��%8�Q�Z�9A/r��9���:�!�6��2O��X?U��Δ �\����gB������0�#Oc?�`, ��}�p�/=O��Ҟ��!����1�w�\�ʋ�-�0�J&��e@���ў���a�h�|+���]�P��K	�ݐ�nQoZ'[���y�̾�ϙ~�+�0x"y�ra�q�:)�*�OB���=�p/���x�����\�ke��̨��"ᚇ��(�Cν���d�CvC6�B/�[��i��'\��kNN�>`�]$ n�*+���-C��&щw������ę��6�5���K0��2�����4�O0�Cz	HpF�4�4cF?��P�^ؖt�r�,�닺M�͙2�<�[3z��[W:5�}��CZ�uS4P����*�!_��䂗����Zfj�}41Ǡ��[W���m��-,�0Y��_��j})�nL�W��L�|z�iY�6���z͜Oq4�mS)d.֝׎�1/�%�hqms���4���;ӱ^��%6_A�Z;4��6��ޤ�9�mZ5]���[��j�?+8������\}�~AA�hB1������'d�>�ˑ��9�S�R͊��n�Pٮ�3LnQ��b#�����[��J�.͔&=� �^k�
"�:[��z;�V:Q�s�xN��H�4F�[\vO5ȸuC�� �5��Rͯ�Ϥ�������7�8������&!��^;�/W)K8�{1�%�l�x#��c�>[�P8u�j�vc�L��uXqu;�CǰA��v�����3T��]nd�%b�qţ�Uh�;YL��z���$�z�g����٫,�:
ebH�V�~�jN��sA�p��R���2L8��F�|"��:��\Ú��/@>G�d4[�g��- �ɛ!_db�C��Xyl��ڀܞj/`S �&�~/I��	z�GW���[>��*w���}�0�a/̡��y�ud�u���e�P5�?��� 6��(nO=��X��ƫwo6/TK�=|Qxk@B�S�G˽S�W/�z��k�McY�I�����0pZ#b�T��=վ�*��~`}U	�T�;� �ฆ~/0������>�u](�l�myGoN7i��^9������9\�_�?�u�Md4.+�||Q�~Se��ƾ�8��3$κjzC�h:;)8%9�a^��׉��_�9j�{���?3�w2f��ݧ��/)k+��5K(��s�X��A���pЊ&h�P&Y�O��w���9��'�Wu���{�w�D��`�à88��
5��ι�����A�gٷ��$��v%M�\��T�LSp���q]Ҏy7�Z�ռ����N�L�HV���Ʋ�5s��ݭlN�q�!-�a�Uo���R�� ПKN,M�G:nt�;=8m�Zc��8�Z3��qĿ�ݾ�e�����c��X'.݋8�-v3ö�(^�X��#&����}�g�e�t�ab��������I�s/!�w�ܭ'W ��|�[V�u)O7Uf�\o��X���o^y�f���ʥ�~��k��![c�UA��`���I����L*&��鶢�ܡHK&�L�]�;�/��j�Ϭy��V�KK���;�ʋ�5p��(>�\d<s�Z�B=9N�[)����KY��;s���y乳�$�TXS.��Ψ�tޡ}��r���k2�W[:W�n/�zc���l������nK��[���+�R��Ruc�j�QN.�t�	�d[BF��Pη��|�]ս��m���i�H8�C�ܻpmΈl��&X^b���kbr�vW�`���]���fk�F�4��?|ZdA����<1��˚��g���3�0S��\�T�m�6�Gr'"�������7^B�f�ӿ3�ˇ�����0�7sЗ���dI��º���g�.�f�gwT]��@���_���#�'��D�Ʊ@�������9�/�(�}j:Z4fҹ���z�m/tI�c��½k��M��`Z���������84��z�!i�}ؼ�Wﾥ��x�gwA����#YV�jZ�'�\�PK�\�#�H=Bu��;�tx0�8��*mt�r�l[��3ܕt[���{�f�/�˵K�͠�WV��9rMbj��|}����Y�h���Y
��:���m���T6��:���"�;w���;�E�[��:��t2Vr��iJ�6�Da�F�q�Hu�6,·sMkI3���H���Q��t�T�����{2�}w��P�ύ���7��U�P%9��v�h����0��=���X4��k���D��Xxh���Ta?��M�2#��;�=�+�P&$�P&Y���̉ѕ=�Wsb�m�N�~�ϫX������y��g�����s��{���^E�a�*
)��+�b��~����Q���%CIF]����e^�xc^����5R����O���Ƕ���j����n �g[�i���W�BҸo#^in��b���g�0Aa`��mv6.�2�M�����i�&_����j7�ʖ��`,~;2�YB��*:�V��%�Mz�k��{��o��S�E�l�ř;p𝚇����>04�?g���;R��:��|d&T-*�Į�g�u �uo��*��c�6����D�.��s/k�		��{�S���xN��`ZV�.�r���:o��u��7�C_q�=[�Hqm 'H>P�'����; 5��I��VW_<_H8�)6�K�n^Sd��Pٯ�2�n��&�B��*��<����B.�����>��SχN�X�"�*�rb��O�A
K�����J�Ͻ��yĮ��L'�{�y.��]���{+�{����9M�T��w	nO7�p̜��j7�h��c��wH{ ��O;���<����\��V��ӎ�=8��q�rM���ݳ�1�zXb�ګ�xy^<��t}p�j�N�%0����P[�H�����.��<�AYc�l�0>���+ݻfW�YS
�WM��k^����*�qWK��E�,���.��^N%�������LW=.g6�]�Q�9��~G�мy㚻��8�vA_{�W���Z���R���1ip�(�%LUH~���+�뫸\���as�
<�����m==E���U��Z�⠗�{Wۖ���*^�$u�ܪ�[Oՙ7�����`0dA���.����m�s��\��3�|zLג��q<&yo�=��3ƾ����} ��a=�|Tjj�zo��7�vޏ���T42F��(~G,�l��e9I���A!my�L[X�c>����.u��ӌ}WMO��~��m������6��7s�A"�&����N�T?PȖx���ޙ���_��8�~�Z���7�~i�}��zZui�i�+��X�B�K�y���z��xj#Ix���{�ԃQ�c��)���&||�Q1�/�rg�%L�vd|�q�j	���7����{�>�/w����{���o���������~���vxP�z]��]�2^��uc����һ0�w��Yz��"30����� �wj�o(K�MV�K	��(2M�O��	��xa�Z5G�h��z�̫ȱ%Y�VA|���ŗ�W~�c��^���yLk��L��XTj�K���ɪ���t�g�x&���ynzan4�ޞQ���m�̶Oo�W�(����3���Ȯp
�j�܊j�g���6~���@�b3|��7��"�IT��(����}��+��.p����X3u�/�.�=���"����	���D�֨Y3�	Z�_s���{��]�ƭ�[���ܲ��_���/�=k~L��N�%�:b\5Z|����eRu�BY�^��B��>|pf�m;��(y'�R�2.�4��o��َGze�s7�0-�ǃ�0W� |�)�u4-V�q�*`�#�w����^O���w�3��,Y1��ށ�e��.�7V��il٢cŅ��^�{ �� jUiGF�8����������F��կ=������7�{�D���9�]`硤,��wNܶٛ�_��9�r/G��R�)�Z�q�c��vP6�x���E�#���11�knx�u{.��{N�e&��pV��Q6����#�4�k�_s6����^Pu)����rqv*Y�}�oK��^�#��=O�+�;+�T�����Kz��J�8�{c�y��r=Ȯ�+4ƶ�	����Է&m2�LdНv1�l#ztL���՞��ex��[��D���Iwv.�K�N�2��Ql������u�{G���M��ε�R�}W��)�W}f%vnǘ�77��ۚt;��􌹑�<o�iW;c{;r�vqw��o��9���"
n����.ўq�Ƥ�v���?l�d�=��:���Vtu�mԨ�6^���Z�k��鑒Q��&1��}v�{7���^�&�<�\O�V9�z��_m����GxP�N]˃���Ҡ���G���Y�t7v��N՝t�n[<侾����4;��1%C����n�"��0^��We&EN��\\��TYm1�WMn	�C/�{��6noS���%z:\�,�V��y�B���cP����w��e�4��,cщ��/����W����-��7��K�'&�t�V�ֻ�!����S:+��C�fB*�u6[���{}�r�}������&uIK$�w���q��5$'o��[o�a�Yȯ3�q�C:�Yg��g��\�P5'*�A��w��� �u��X��^W���;]�xӻ]��B@��E���G'��Xw�֯d#m�ř��h�S�,�H�\C_CCD�8)[���%�\��ca�M>����7HM5��<�|�r���Z�9RF�rT͘
��z�j�>�Xv�G3�����z��Q^��VD{1�w��QN$��ua��#}^q�EW��M�ܝŸi8�t '�KE%CQW6�J()(R����� �����(���*��((("�&&�b***���)�(()�Z��!� JZ
Z*����
	�
�
(�(Zb
hJ����F�����	�bih�)*$��(����%�$
h�H��*�����
a���j*i�h((*$)��"
J� �������H��R�U@RR�%TMR15IMT�-MQ4P�PM4�R5UT��DMQQQ%D4$M4�-U%RT@O�H$?�~��#ϻ¦+�3y��J4_,��v���1�k�3%���-en����m��#�e��^gV���� �t]����$��v;��xA�CP?��)�=�-�X~O1q��S��;��"Se�3�2��v��B��?a��b[.��[8��{i���ǣ!�0<0����[ ��U��Pa�����m�Ƈ�����7ð�F�Ȗ[�	(��(�7a��ڴ�++�?R���|��8��}RM���f�Z��Ԧ�c���i����(�;�t���rt܂F�[^�i��X���c�C5��=�ew�Rә�ty��6�Lpc;���I�;��O��Rr�7H�^�\Ø����}UZp`q���9؜���C�1;�zM�&86�G4��S"�6��8ŧ�����;9��$���G(�v�����Y�
��{`|�[a����&��ݪ����/6�k(}����[dU
���2�9�jĆ��8�`k���~=��?.�t��ZjE1�5�|x0k�!�̼�q����6��p��Jvޯ���T�eى�k�q�����*����@r�Q�MK��f���:הJ`��e�OG�x�b�A��۱�6�~Bb��Ͻ7+�
ӯ֢C�����nt�{�Ի��=��/15��� ���;֫nn�Y�;�W�u�f^y��W��3��1D���D.�0�hy�-�1�;r��E��W.���OH?xkXa:�F�u�=�*�n��;FS/[3n��2B�m��vv��9�l�����N;U� �$���|ha`Ih(��oQ���� s�<{]]N4!P��n�,��!k; 8TkO�ac�ڑ�Wt���hEQ5e��L�kO.�|tE�1�HƇ�y�ǒukc�[[n�;��<�Ai�Lbuc�q�������f���%��T�`n2�M1��O�2�n�NȽ��֊x[]�`0&B���ɫ�W^�kbt���[�`�i��j����t�r�Ő+'CR^�U~͘~�1� /��'c�f��I��{��W���J|�i��L?v��'ֳ��z�KK����c�d�C���
�"K�Xvs��y��cgQ~�g�ݑ��MB2z�C,{��X�hR�*�
j�q�^���g97А��jQt�w;�7�
�]Lg�;Hܗn��M�A�$�b%:H�y�)U�b:q�q�����}��M���)yN��H1�0�$H�a2�&�ۃN�L4��T�p���$�]N��1s0�%�a�;׈Z�z����w @CS�gb���0%�a�m�)�|��T�B�(<���=��v��]���� I.Ͳ3E��^ގ�iV^�Ho�����	���'�޸�(I�P˙�*Ϻ�J�ཎ�^O0w�eEle�>��;�͈­����EؗKlMҡ�i�=oP֌2���L�x�bnG0n��>���S�+i)���^�sx��Y�7�j/�8M��瑵��\�"#�����|-{�9���yO�&�B�}�N�]�ڹPCM��u*ah�)�T$�srGj&wvm�{|p��,7L@M���ORq�.�>$��[~M/k�WBՎ�Z������̤�u�$�}j����3��*����0�wT�g����Z�@0�����dR�J�i�W=��s��A�4�+	p���oP_fe's�k)sV[/!fqAF��|�U�,�{d��8��I�k^��Ӥ�72��cv���<�.wt��^b]{�:�w�����~�9.�:�;����QaC�sȼ�����J�<�����/oY=i�ӯ2� �n��l��k˼ `L�y��a�K }B���%s���K�Ud��pѬl���B��� ��˴�l����5�̀���e��3'�$���j��W�qgו���p�
�Ō�1�9��xj��Y!
�k�o�鳣���Ί��B�<7y}�%ew�TɃ*���,�;�����*Zڽ��-{;2�r%jTu��ޜap�c�=�l�F&�lBn��:}�l]��^��~�^#��{�bw&�i�2%�`�
+/s7�m�f��DL<I���JEDD�oI��H?(�E��Dd�
�Ymh�~�#�2�8�	#�S��!l�(1�;�724��`{#��1yT��s�+k,V;�k�+B��\�G;O�N2W�ږ橶�"�U�	���Rx]r(�aS��c0gW����w_Z�uoV���{ght[O��/�&B{+�4�ا�����x����m�ua����Z��S��؍�ǭ}ǂ��|w�Hqm �A�	����^bP�������/!�W�h�d]ctS*H�aA��!A]��ZX�̜K�>�/��^R\�MYH�kGf2+z�<��N�_*�]ye෮��Z��mxp�Ђ�lnU#o���#��Ci/�6���c�&��ΫeP�vT8�t�1i��(5�6I���'��Wm�<1���@�S��B*��N��0-�:v��*��Q��e6�α�3�5 �5KfS�ۻ��p���N@q#�`��:�ꝚmQ�Z�p
Ucz����~3\��T�i�^t��\�.�+��W��2Da����_22vdnt['*Sv���$lM�Mql�:�tz1׸��P=��h���Ln�����u𽍨d�$���F��Y���������ݔ�z�3��y}���&�[�r	�R��e$v�[}9۸�u���	ц�]9��|����#������`��j;r���`͌�Xy`Ck�׷,��9���k�]��U?˦f��M���A��3�~]��3O��Iue��^��1^�tE�j��g�]�|��������9��9J�z;-��G;Z�t:�9��M23kCw9!�8ot��o�؊��"Y��B���u��uΰE��C�D=����gui��L�W�X]+Ô�p��I�dXNi!��Oeg6���r�ʔ)�|a�����X� �����q�8��3i�A�Y8�4�����Q�Vb��4nV{��>�!+O�|+f��b�O����&ap<������X�,��V��D�S�wd����zべ��Fo������^��Uj���-bO���2.�	�`�#3j�d�_.��,�{��Y��\ �K"��DJ4�����9쯔�J���?�O�9���!<�y��XRƽ�7Xcc����4�$�<��]'�)Յ�)��&���͎�P�=��P}j�޽�S�Z���������a�ИA��K�]�a��F�|��`�)V*��	�/7����"����^�y�<�VY��C�	������I��a��j}b��M �oq�M�ͼC����PJx��[��ܣo�|�\v�F�Q���{�"�s�iQ�iN���Ǽq�m�B4�v�����0I����)�xRr��0(w%;�v�@���s��#u7�ىQ/��v��sx�<`���x����ž��Igm�"]L�+��ٵ��.����V�9J"��������N�ׁ��.�8{�N�vB/=�uʚe��`�[ޗ�k���g��k�J9?6;��K�@��v���{쟛ƽ="�՚�LP��ly�a��@yŻ�D�8�I���)�Z�>�W�럘�T'+]�N�d�q��ĉb�!ڝ'a�!����*��٪�6�S��ȣ���^5���z}]~5\�_�?�C�u�l/8x��E߻�d4]=�|N�"��C�qzP���d?p:�l�Nf�qg4��j/���?����N"(PuwA=��(6x�:��,Tc<9��)߶�ʶ"f��6���pK�w�sZA&�T�!Ѽ��y��@@���Cif�EE'W�8�n{�?����I�O=>�M�f�6�Y:��jۃ"�]�[�Yz�xU�N���!�<���5s����/�fp�y�L�+��d8D��Ed��3���8ʆ@�t���B���'���S�'a-s����Ӓ�|�$�cP�'ְvi�1�����v>S�����\g(�>os��қ�*����WP��)�́��䴳��V���9w��-��c�·4R���Թ��n�l]Њ"��+j��ʶ�<�b����d�V��y��3�����nʉi��]�Λ�m��?Z݃	%g��v�Pç����l�k��M���.U�@ؐk �h{����>;:ɨFB��2ǿq):�1�J���jꋇ[E��gU�l�h���]�z��p~?��Bm�r9��d���&I˼'It�(J��]�C�������(�sf�]�ԋ�L��h�?���~k� k��6�<�6s���ȳ��m�4;̣p]�C�T�Э=�·n��(���0����0�'�q����C���V���*��j�,�.�N樚oR�z]�l��c�o<�~�D�T�e��T��=ʿ�˪c���kD��g�?=�U�<�P8ޕ�@Y�I�ҒƂ;P�Sû6�=�����p�a;��iO�&e
XKs�[iԘ�uc��Z�u��%Qa@Z��S~WZ�|^�����>��[+2_g�R�(�pޝ�Wy���>��X����д�D�q���{*	{k��a �	֌��ZPi�Zf��&�;��;���4����s��w��j�ԨO�Z�]�3*Ä��V!��(ܲn�n-b�2'�ܬ���"O���a?��4���"):����.y�;�����.U�C��뼑<4�F���K]�&1�s���(+!�G�Sd��m�[��Ӝ.�){N��
4Z�u���~,����JSR��t,.���b��ώïm�=������6Q��)��8ͬ㯵�E�p���u��d<�0p��.�S��_�涎�������mע�]�lh�l����bhY偩��(l���n��	׊�`���E��u3����D:NmC��hzk��6�Ɔ�f�\D�{0"1�;�햝�\��S�l6b�u5^��lkf9Aᷲ.U�CB,k�o��t�ê�E3�5#Ѳ��*)���X ���D]�s�TcR�9R��T��aUk(RJN8~ӌ'�-�WJΰg튶��o^[���ygZ!66~k�9�qN2V'j[����g	�ҡI���-}}�tnNY�˒-x���ۅ�VQ;?ycC����AB1O5?!)��`Kk�Q���p[s�'z+�kp�q>O��8��)*��l�=}Ǆ�.="C�d�� ������JF�wv��ݼ[��;S�D�a�;��ĵ'C�YrF�
�|ᮢ����e���p���ս.�f�k��x��gN�Ty@j^�i�2�<�EL9L"�y�)�-���\���ׇM;)���W]R��۷'\rf�^���Lc vl�(qTqWK՘��֔+���&�(�~ڑǵ��k9�� �apBtP��x�����_5�8����]��8���Hd�;�Ǽ���{)^���ٛIS����>HjU)1�j~F��4u��s�C)�[e,mU�m�aVE-�o� Ѝew�C}Fv�8]vb���dE�=$˼K8k�O}��=�:b�!���Iј���D��еΦ���~�Ȇ���E�ڸ�!FZ�R�9���}���/j�(�ϧ�2�V0G�k��gN�(=��7;�=�$�.�2�\sO�ܳm�`�>������"��h���������@�e�I��Պ��gZ-����儧ӮLG6����@G��$����_�?��SV����\Ց����{�C29�{����^��y� tE�j��y�޼����j��m�vei���7<^����	��Fmci�Hz�H�z���K����o�F�ڻ��
}E}��a���Ljϼ���+��`��L�W�X�WA
�).���\���dx�K��ؾ���r��3��S���M"22jMO��r"����l�C�`��NV�VRw�y�հ�^�A�g=�g�e+���!+�Ô+���*�|�ʱ�Q�>��H�
Ҫ��Ņڶ��������ǟ��є��[�{lw��`�as	�������6g��>ᓭ�����䱞*�}�Vl������X���i:�ݛ��O(Lan�,,D�1�ĨL���lFeoZ��*��\��wt�;��zͺ[6��n}˭����G�aC%a��8u�J�u�3��Y� �ʜ�9�I��8
R�*+��޾��]�\�v��#���A8�o�I�$��V%M�̙�}j�=�򂕤Ǩ0A>�����u~ys���yٺ�r�iOd�z)�r�	��S	Mmx'�msG�b��*ZF��7��m��;��[�c(JY�0C���I�;��O�"���7H�X��srb�Cՙ�a,������nWnb�u����������M��sۛ���+T�H�M��q�O�n��1���_�:���otu������.�`y��y�[!�zg�9	�c��]-��;~�7�o�KTpZ�]���O<�zBn��Tw=y>;���/��(���:r��z��B�}�x(���MӀ�����ތ�5�c�ڗ��NZ֙6�j��j��+b�ٶ}���|D�^�
��Q2?`]W�ܳ�n����7=Ӡj]Wi�i<&Y�:�WX��A~����!۵�4��+O��ELy�C�[!��چ/�;M�;I86��8����i~�H��������J[�����v�,'?��
ˑ�� ����;#Y+��@;�B(4]�,Ż�>oG�������y{���w�����}�#����zET���wM�(�6R��Gii���0DlVjz��be2K�.Y�-V֭�A����^d��:����ޝp1�:S�w=�Ơ�ｆ5��C�}��J*xg��ε���=��.�I���zQ�����ۯԤ�����e:ʄ�Նr�gd�D-�0��^�}��Z��j�V�j�`��u�`@�d�3��p2w7�>/\s;�6u%1H��䧡r35��X�gK}�7٢��f'x�'�5���ևw�T���F��/e"\�[u�twB϶��
�ǈX��;*��[w�6��B�֖����3B���t��  ޥZ�������9�]�
?m�l�;��)���w�+r�UV�a�pŵY�� ��ܱ.���+Ey�Ҹ��c�H^�aV���\������lo��0�Ȉ�-L���D��8JVp�r�D�h�]�h!y����c���7��S�Y��j�S���2�`�;��1?�����mvlZ3��0�}|��(I��tY�$l*9Ίɘ�W,����XM��NN�Z����)��;��L��2MB$c����x�%ct��vh��Ƕ�O���Op4*���ibP�f�@x�k;(Vۛ�B-��n^��E�KL���m΃M���n��Z|�Ū:Ԫ��툙�+(����Y�ܮ���F��Z��K}�{;�݃H\|��ۓ8�3��}���$Mf�Z�~��W`0�Pg=�	�n�Gy�;ǣI�깝��!A�v*�^�<"��7��Q���~��aK �{����������[�UG���'���o��ľ��*�ɢ��9�b�,*{؈t�N^�8v��\j�Y�Y�B�BB䣭�s���,�9|��-��f�Arjt�\�]*����9o��E�̪���:�د���7Yԁ20}v�I�r
��(�;x��9wGQ3a���Y��XW�{hm�\�uC�w3�I��M(r��YsvM�hU�*��U��-G�`OM��\j�l��Kef=)mt�vP�����bY�f��*0�|bXǌ�Lӑ��tP���q�Zݺ�$�wZG��j�w��Jhח5��=�������P�@UARv���5��S���]��x�f�������o�S�"׮�n�4ĿQrK��\"�Z��]�\��s]e��= =-C�]&.L���r�=�sNC�.�pBz���^'}wg��K�����Շ���;�d��������t�����c���KbCY(Y�k�/�zjW������x�dMS.^j��X��u�[�\:�r,Ƅ����7\	.�_����y�M�܍Q��<��:�[��79*Π���u�)���R7kȗ]V�W{��8�ʯ�N�����ir:�o"�����R/�^��wZ3rφ����EdS{l�jd|�C�d�G�N�fW=������7�:�p�(0̦8��ĐA I��i(�����bP��� i(���&FHJ&F$������`h)("R�*"��(�*��)h(�Z��������)*�I���B"��hH�
�Ib��f�� hbB�����"��
�
)�������������(
JJ*�"	�h
�J*��hH�J�b��Z%)&�*&�
hh����j��J~K�*�%�)h
��	�***"�R� �����*������)���V�*d)��(&*$h(
H���g��Ʊ^>u�u�us��[]ޮ
��+��0�b��ä�j�5�sF�v��KaT�Nڝ���-U�^���oʹ2�5��8A�v,��0��!�4���3�d�e ӆ�(Aʺ�s?�����z�C��Sn+[��66�e�C�h!��*�-?PH�M �ڀё���:�:�m�wOy���4�){;]����δv�f�.�b�/茵���y��);���c��|�{�d^�}]-]��S�8�uؙ�m(n��u�̒�A�1�����T2�����W�%C��)-��{8yN덼�ȸ�����D܂lNEcr�p;'���]X�@�c�y���sB�3>��r9�ͷu���c!5�!H�2��봍S�Y��~b�,{b���hR�*�
j�q��\�驆
��}x~�SK�T���e�Y�0>��r#�vO�\�$����E9�<ƞgt]Q�u�g��渵8�w"�t�z����2�}�̠�o*�����r�Hy^�~m'l����1��)�E�o�f˳e<0��B1��O���~�%���8��H�r�+Fd��g�qJYi�)�Ʃ�E��8���
�t�D�\��
�>�9��f�t�9�[ZՏ�5i��Wkk�R��x�yk5	<�RX��5<8�4�`�������_O,�{��#��ޭ��
n2�ϩ�s\��gDy���b���̤FT��F�x��0�
!N|�_z����@Ĳ��um]t���P!��Y���є�*�{��%
ݭ;�R����+��yE`�b����+��۵����;�Aˀ����| {��1x}��;�c��N�7�WB̀bN�y�<J�a^��̦º���[9���"H�l-�^�Z��ˍ��!�"����Bmj&U&Am����Q+\u�?J�T������=QQ���j3WM�R��Yz���#k��tHB<���4�}Oյ,�-�Û��@��z�3�WP{h#$������J���Ǡaz/a���@p04Bax����쓫�L��iq�^������_����s�{Rj��N�Q2�uɈvâ-�tg/#^]1��~���~j|����i��>u�D�2c"�5{T�Țfy^hwH$=%�a�q�l��m��̀���W	evz�<]n[��ӮK�"�s^���Ƕ�؁����xj���p�r5�\m�j鋇Uo�jz���,�k�[��c:�	�Xt�=�Lx�z*1��NT��*B׳��*��)_���d�M��rf*���?��������1P�W�)��cH�0�}#��F2\'j[���"k��W����/��!<1{=����!�]��zWe�Ӻ��V��)흡���K�	�����#�O0��㪧i��h��*���lY+]*�s� .v�)�W�qo:��*T�<�,�޼��9���zυW��S��3���bȽ�po	&6��>��r��S��M������e,�襊v.N��&�.[�����*�k �Z7|A�_�<-���ޘ/c)ď�kG��%?_���5%P���x�5����!��yO� �s ��ث`�wf��|����m��O��I��d�`n�eA#I�?E�w0��=� f�M}����U4�]t���8�_��ihvQ��vEL/ܪQu��L�oT7Q�NZ��k��V.�[��ݗ��р�.��Bn��[��У~;JQ�=/�Y�O�iAcK���)MW����Ŋ9Yv�?=n`C����?��Y�}n�	٢��M�-GNл%Q��Z��S���dġ|�p��@�0��>T�`n0��zGB9��_j�(��-l�J�`z����j���U�N��T��u�
{��q�>7rʹ�E���t�
9��3��������U��H�F�&T8Qyћ����t!*L����ɟN�fy��f4_�a���8!��Y���8�?scߔk޿K�9͈̀��Y��� �x���D[���@�~�_2�.F�S'�Yػz3�-`�?cy���M����r����6��4��$= <M;H�[�o��Q�\���`��|i�E�^t�����c�r�S/�N�=���T�p�ͳ����;rH���t���c��u���v*R��*��K�v|3܎��g@��X�^XU�6��=��+x+����rͺ]f�m`��j�g��o�yxev�X�Z?��R�y��[�������?41�߇���=�Fk��z���f�����]%S�"�LK�J7�Ef{��������MR�:YT���l������y�rg)�jJ���{��dNJ~��Q\�1@���<��C6q=���O��)&0 �Z�B05������L/���Dq��P�h7���:��D��&Pd�-)���]8��z��x/B�� �d�Kؾ�i&��f��Ɍ��~�"�:9�|S͡�N8�2O�H�2�e5;�s�:y�=����v�z�(쳝��������&��iOd�~w��?x�Juk�SH�kk����Bt��Z�f�r�aͺ�zJ<�3]y�(fݘ���;��T>����$�b)9X�R�B�_��By��yc&�~Ƚz�dy�CE����!�l?ܸ���!��Bn����6Y̹֩���
�Q}('���ˎz(u��a ��=�>O��F�혖\�ՓM�Y�`r1u2��C�9��;)KZ&Jy��}A�K�J;����q"Ƽ(���:r��y~����]����=�����o���+*o
�Nk�u��$P�zJ��$��49t�z��+�K�N��ݸ������}zd��0FU�a=�f�O#g%i�1�]���`�+yH��Lr��t��(�y���G��GpV=P��m@����}��<>~2S=�$�s������:��ڑL�)��=)8Y����\����v�,a��>H_�^漿z�{���&�C�t�����i�j�JaşYc���>3:�϶���u�3OA�쳉룍oew4�����Ƒ��׆�1s�Mxu���i�i�qhIy�y�������O�x�\���i�KD�!��0(�����	����'s��]�TP3ОNx�+jǹL�1��梀��,�>���*��E{iw�_ʸ�Ϩ���27��=�I�Zo�������ͮLҸ��jHA����`�Zz�<�����ϐ�a{�d\���sJ봞�#�wm��r���ƾo9!��AZ��II>��e^�Ξy���q��6B��N�Pۇ����)Ї�zaQ7#���V5�I���	ͨƒ��tq�Ɋ�U,�e���9N��[����d4a�;>�Z�b�n�ϟ��X�8�eV�
S��+��>���L^��[q�}p�B�.i���A�k�L$�#rG	���Ι�b%:oo�흊^�	��zBOܸs�(U�*;�m�q�u�I�Ts�$z���}��֘s���u3ڨ�e�����
��Y�;�y�ug]Y{Ͼ�UԨ�uxy���l3a���=Oz��0�tR��[�\��c[,��W��n��f�sG�}5ez=f�L�=��|@X�L�}m�=G�����B�!ZE	���g�L?�6����2ڇ����ΐ���f��t�9[��:��kZ/1V�"��\hW��r���"~�a�����������Y��B�5�^ϴ�x�?Vo�=q��|��/}����}�rА:�
�� ��Ň܋��vE!6�B�\���G1��w$���:��Y�I�r�oL0,���ې��V-�<�VnI�:6B��$�'a�J�WBK��.�TXU��e6�}l�K�kc�N��7bNK^)5����P���8���|��6��2)��=+��T���7le�k��y���s�Bq������<���g��&�nO0LqѭklŨf���4��!e:bN��R�����V
�����-�(&��<h����o�=���V���#�w<��zI�½�$�P&Y��1�Ƈ@�r��.�1G�Ax.�v"/G���៸/�?6�ߺ\��`�C��sv��<{�$�-���OՐ����R�7U4�,��a��/6��f��꾨kE��:�g^:��\����m�le�����e�{�Ny�h;�b�M�S&i�4��-��9��эX���(�\��k�*UǗ%fò�nU�����x�q�gf�>3�G%5�}��ޣ<���޶
.=OE��^�kO� ������B���\m�f��&�r����M2�4��{)6��
нHx�B ��y8�;�KcW�)^��A�Z�	v��K����:Yma��ӇG'M�T9��L����v]�ڧ���nXH�>iMd,�α�es��<�^�uq�ǤO:��B�Fcз�xjkgk�-�8��pH����di�c�\�UBp-c���p�gǠ�'��B*�j��L��M��#2���Tr�j/�Yq;K����lDe�gE�I�?_Hk�S��[��������F�r��q��=��M?o����I�b�y˼ً��rf�;%�7&�p�,���΅�8����uXH��P�F�4�M[Vk1Z5���R����(@~��lO�;V߮�(ğ6�*�:�G8Q��s�s�\�/]�����Ϊҏ���Uo���J���������{&�䚻�W�8�{��՞�:�_,������S���<o덢|�g���i�I�����T�M��b��۷���q��0�3��9
O������N�5[4����;p{�o>+ŔL��I�ݽ�p5���s�� ���<��R.���WP(�j)S�tȯ]e��� G8#���"�݋�}v�Sg��m��7r�P�yP/vԟ��fzuCV���R��Ki�9틥�eV�my�,�q6���&���̒��ʎ�L�g���w����a��y�e�1G���W�r�f���bw�H1���8S�����e�L�	}���E?H�g!��WC�K��N�������'_�֢؈nr&X׽)��V���{^]o�Y��� �᪑��f����<o��f�������F+%�\��J�GsmH�e����q�a����h��3�k��oŲ�x�B���P\)GO�۔��d�ә�AU��O�/qC6_sv#&��Z����KQ���P�)RF@N�0��5[��˧:ff3
�U�7�]1ۑR#�N�p�غ}���x&�J�^H��7�囹D�ь��j�m%��x�ވ�)L|"���gqU�c�E�Z�\��h>v(��Kn�t�ݭs�>YiW_ u�W��]Ơ�n��v�Z�홋� ~���)Qk�ח�{��1dN�KM;�xh��s}���ms�pʊ}�T�b��e���w����M4�]�OU��_z��L�_�~�~)�f�<wJJ�:�yu�_�6�W�a}�4i:���fbT	� 6c�g��e��kn�m;C�B7��/C�GQ���{�=+�ir��c�5�}�*{���������Y�޼�9R*�g����̟f��gbGZJh%ܻ .�-��'˭6ξ�֡��zU5��چ�c�M�J�����tɕ��f�ňLXf�	�W6�5�L�K�d	AooS�ᕦ�u������z3��2�־{�h5w�k�-�ހ�}^og��ìF��[>�;'��U,wvG)�UT��q���JiMݞ���+��ʺ�>u�n�ע�%}Î_��}�9��c�i�Å����1H�tQ���2�@����Е�������=�Q}�v�^$�4�$D{O4{�ڡ�ngCz��B��g���{^9�JwuzLS(W�*r왲��u/�e�}���lm�Wh��@�Oor�M�-e�}c'�`D,���D�Dm�W8RݷCZ�hM�ղ�0�D��Lw@b�U��hh�(�1@��}5�ivi'��YE�I�����������;�9�&�����W0K�z�����OKf�J�~��x@���W=��7s�=?2�gǒ��T���|z�:ٽ�����~����7����F�ohW^#��O��]AN��q
���=.O�H��i|�~����U�w�.����.@����6�Ϡ>��
֙�Y&D��^�F��3���������#�t��M����vd	�!u,��ps��˧�����8�GDׯ���:I_���@m���Ngَ# K��7�M���횜�;L$��J��^:��q�Ԥ-��==,1z���U�j�5�j!�*�m���
�y?S���c�݉Ux��F�����R3��2�$0˽ʛ�uKͶ���t�W�d�M��w.T���u䛡���GnAᛢTX�Ȇ�b��.�Fv��4�(X�VH�z|��w�����{���w����{���￳��o��������kkg��-���f���ي�V��C�͵��K|4\YiR5}`�u��J���]f{w��[ ����vz��4a�U��V
��!����ŉH��	��-u�{��ȯk��>˥�����3���hB�gGؒoct>�.�iF	+�6���������}�M�:j�M6�����č�ckE��.���P���Y�n��U�A�O�޼t�چ��B�&��Ol}��i����ϫ�8-}�j���g�7��ܾ�Axl��ކ�C���Ls,	>���Z���F�(Ơ���̮P6ö��u�{U�����<��h>,�:p�ְ8��꥚=�U���,l_M����#��nޤ<;��ڴ���}����^=�&St�+��v��ʓ�.�=J�=�o�R�f[�Y�k	#	M\���u�s]��D=ps�y����,�hj�cjxV,���
����I�cQ�"�����(Z���0zP�^a��4H�:*�$�7�!�f���.�z\�Qޘ�qM���d���b����!��k�d>���L�y���[#D�w}ݫR<w�`Uh�FO�K����,�}�YG�~c6��cб�>�z�F��:LQ�"R�b��=�����S0�>�,�r�J�U���j�n�^.�wW�����ѧ���V����o���H����*ec[�ITT:eě�� ڳ�,���5?���͙��Gڂ�oj޴x�̹[�*��7����.wU�A��'-\q�SP�[���@��jǲMf��y��������wJWΜX=�K��,�{׸��k��M�;sw�ou D����;�l"�!q��M_LCm�Vm��B��r����v+�&�R3|;X�zkH^���W"zw�қ��ұ�{=���"���O�X��;ܟ���K�_8��"�X� {�*�EK2�=Y����q���X��MCe���'�r�Q�^�����L!�숑��3N1C4�z�;#Go.]�rӹwP ̚�9�r�C�������z�����e�]/,�����w�\�_��`�}8���'p��۬T�Ƌpի���R���=��hg�uz{�x��A/!s��О��s܍��FTwGaP֡��6�\����5R�j��s�E�oZ�]��ߛ��qS����կ�����r�T��ģ�e��y���R�g4�ԃ{�PR�l�	!4�ÃQ�ΝG�s�jM�t���c�_vK��4G��9M}�`3i>xCj��8�<o��5h����H���jQ��sz�ǃ���r/:G���&�W��B��,mS�|�q�nL<�U�7��GM�coȖ��o{C	=�ܫ��s|T�ݯ��^=�~}�z�45p�}�E����CNC��Q�w��!`��vDO\)�-gj�'R��\��c�����_.Ȥ��)�%�9V~?>ᤠ�
R��$�
�JJJ���J ���
iК�	�.`ґ#A��4�
��ѭ�D�R[�]UZi4�H�7.M4֊]5A�H�AL4&-%1#@Һ��1��J(b��8���t�+b�P4��)����h�(�4%V�.�q!�kA@R��i4-)Dl�Rh�.چ"������4��颎G#�Q.���h1@h��!�5l:"le-�mH���!��5mV˶]TTh<9������:X7��������R	e%����3s���.�"WX���1�u�r�U�����%�IeK���7S����3�����t^�C��;�#��F�H�fP.�}˻�rDѺj�=i[v�i��xq2Gtl�,4�0�������-���;����k��9���5�����(eIS�}�l��ʆ�-�ڇlz�z�o1�:��<U�ɼ�}â��=��$o�pTk���׈�,�],�c%�O]���Ȏ�����(^!D`��=##e�W]{�1���W�F�L枮(lu����Q����/�y������$
j�8"c���Ċ�:��B��<]9�u�r��[n������������e����?G	ŉP���HɊ�ɋ�~ޘ�p�����><��JUB����7�p��Y7!��ʜ������Kvm�RR�2ЧH�;�Iz$�������U�f�w�z
�L�߷�K�O��K�����R���*O���?_O�����x<���D]�Z2/�ϡ���H�̆���k�c9w��2�+��/����b�n�U�ΐ�NQ�G�P���8mC�g�w�}N�̝�;C�c�ݦ�2ǝ�W��Ӷ��A7c����GG���@��X��{vY�v�p��s-U��r�Iʐ�2<�#^�[+e�n�%~�Ԋ��R��e�j�f��ۗ��]v�Dɳ� ��8��o��q<x��ޓ�����2�1¨��Ά���;���2S��a�t �cp��U��ڶ��U��83FEndVjj��=�_��\e��t7���y��}�L�<[L�/���z�u�Fm���R��.��y�97��L��O��b8�>L*muP���kqԺ�i1[��n�ܧb��=C 6�6Jj���R}xU}y]����lE͙#�wl�#�����;�{Es?_7)2�F�:M��]�i��n�wd#�,׶q*���χvx�`�+���C�ͮ��]���4�b2�)ȧ��C:�B�<�����7�׻��5�ٶ�OE��ܓ��xc:�E^��g�e)�FK=�`fB�T���w�B�찺x�ɣ*�65�}lLnk�~����XJC�̰�т���=�0�ޤ�D�����/��-��D��k]>��Q���Zά|]��3���ytl@�\��}�!��R����V���4�jr3n�,�*�O\��������3�xվ�˸f��bp2*����^��_��&�H�^R�]2�i�p�[;�>�x�D^L�~�X�h��g���Ҏ'ii�ɹ�4%�ND�\UT��A�qS��(�a�L��� ځU�R�����3�>�pV݅V�\��xBD��5+��:��n;O��49��%Q�=>��SY��l\�]R�9�5��T�P�Hg����ڧs=��	&�h}�w�웍���e������3��WQ6s���m�\!O����܂��tUF4K��y��U9�EMy*M�I�V=��>�n����-�#z�����R�݄�[ާ�>ٹ��gì�W$���r�| ����!�9���'�}�{c�=מڶS>�)w1��]*�9G��{��4��\�i��@��;u���/f�k�*��=��iQ����� ������R	��}�'�T��%�uʚ��vi��@[�{\b�bZs6��]n�Xz�׸OfZ�!)�'z~�����xԆ�C��ư�o]�C����0,}�tl�����3(��qU�q,!l�[�t���v��b���E������!��=le��^e���\�0@��F�]��È��*P�3:�n��좻��nl������dڿơ��`f�
�z0�Vp�v�)��R{/��l��oF	Ô����¢����`�����b-�'3~����ަ����ȉĉ(���nYK��nd�.[.�8;UX�k��oWs�K�'6������Hwa�'���}C6ԍ�t�ˣ���1<E�ɭ�͢��,�T'�=����y,������[��ҡe�s����N��{�p�K��F�tňP�@�h�����t8��=o���=���Y����2zi�M3�Р��Hm𽵩�hNz�|���/)V�g:�)��>ZܧYّ"�$��(Ox���A�=o�j����D#l��� �ݭ�'��*|Wm�.o12���4�jB0�ҕ�h�v5�}��s��Od��fL��d>멾��=`f��T���YC�u�h'�m�z=�;gi�!ޣv�f� ��J�<���,\'�-M-�-��uc[�͚2=�+�*�7لZ�冪����1ʚ6�a咹�Ml�t�B���m}�ț�EҘ}�z���x�QV%J�5.[ϲ��a����GLt�]���a�+��.����v%<qtMJ��k23��L���mïs��O��e��}���>9�]˕-��!�iM��i���ܮ�)a��}�6k�1�����Y��(V��Y��� �aލ�橋�7�ұ+��dl�7o��oPq�.��.��٠�Q��ۛʑI_�����>&6}�rK`�`E��!�lM5k�SX�lvɷ��Y�#o�W��$���]#M��9�?9Qo4u>R�'j�\G]�6ČR�Ҟ�}���=>���\rVU~� �O�ズ����rf�U�Dn���m긶�O���^P�3�w�®��7va!��ʈɦ��ncW��g�?m�@�;���(w ����Q1ӗ���m�t�=u!��d	���y�蝼/��U�y��d����:j��䰋j[��k^�qp��)��r��e6�F��W]�B4 g|��f�a��$J��q3x�J����ǣ����4כ���{=]���:�ٲ���H�Gz8L��.�ʏ6g=��7���#�l�I��^Z��s l��)�# ?G	ŉ6�ٳ3�#��tV����9�\kz<���w�u�ۺ�sb�� mdY�f���5��m0�
-!;����#A�k��U��۹>�R*�]3��Hٍ�Z(����d��l����ϒY��yt��M��e4�?�J.���<n���X8"��[S�[.�����J(l�4�\����}�0���Ƿ���ɯ�  ��H����	ΓG�6�&�����l����6�/���Ă\d./����m�0����|��j�l�C���X��k��R�ӿ���1&�	ݟ] ��g���z��	(���Z_u��{��][sO��lU��ux�j)S��E�R}��o���*�V-������e�7:�9[͆��a�1�X�t���{e78��2,bl�{$�4��I�K�7SZ;7T�47����1n��ܛ+"YZ�)q��P���\�|u������c^�B�:PT��p���7X��Y����^�{��^ǝ՘zи�`��?D{��sݐ�͟_/���*S:�Ғ���ݞ�;�l"?`.El���3�^)�$ƺ�+Ѹ[g���3$���_�E�()�B�J�NJ��UA��<AP0#
�l�T7F�����CV�M;Zz��&�΂��cOn�+^]o��t+��~䕙ͭ�����;�����:�p�w��J�"Ţ����������᪑Zbk�+�R�ە�c�O[��p��$�H%!ց�c֕�u�:��]2��z�:~$��5M��Dі�kz[�㽔^���v.2O��Ҏ�v�̑sNjJy�*�Fξ��<���B̍#�v��P*��R�~�����ʿf��蚁�h�y=k��Ə�[��g9ӑR!>܏?	�]8�+��}ޭXF�Z�%YY�}g�(���%y���͍/ ��H@~
2�T�s���鹻�拝9תj�n�9�M�x�� �21�n�!��.|G��ꆶ�~Lg������?y��������e�]Gsޤ�މu1�����v��]�N�#xgն��q�{m�ձe�*!���U�/��_%}d��И������3emrC�uD6n��>����{�(�s�+$�ކ��rB�eÉN�����/��o�]}������y�H9���T��޴�y�
�V�����5tF�ɡ�fz�{�/\��%ܻv2�㔠W�������#�j���.K�Nȍ�=
g��� �R)n��iA������Qћ���]�����H�q�FGOd�T`�����`�����H�X�u�m�����2�پd7b86B��;'�/R�z�����:{�E�ŷdq�:|v��1�q���*���Ժ/x��G�n�^���t�;�����OtoG	t>&�^�^�����P���=B�KWDJ]s#6�'��<ut��]�.JSҊ���Ǟ�3D�m��5�8!�k�m6ã���g�&��ٙ���;)R���a����0Za�����R���u��.��S�"n8��\��aE%��vn�cC���g�'!�S~��n�~<�^�b��Q<i�`vjf��T�MX��Iu���-��֖ޗ�-,�xrɺ�7$��;��F��	J8���޸�<��˼�xI�ܻ��peH�p�}��-���߱iȁ��I�Xf�#�\�w\�c��=�Oڛ<��Y�]��^1t��k6��5gc���n������7�Wf�'�� �g@�("�А�m��؛0����Ƌ����xI"���-N���-�B��M�u�/S��.靨{��_F�q7�u�Ig��O��!�vZ���c�e���|�){�h;ۓ�L���m�t�ð�\�j��jw��}�zx����[��={g�'M=��*�<�.�=�3�;�8�(�Z�b�-�;��c�Q|(�;ݷo%���'�����~���+A�':�;�'���5C]>jW���$�flX�.�tİ�a$f���gj��J�������N�_YM����+�{�\��~���{���a�����L���z���Z��5Ѵ(��JNu"���1��#��l1�G�~�z����8�ٕ����䒢EX��[w�r���z���� *��?aFh��{�͝���1��a�@�j3�6�N1�����nԧ]�����,'��[8�SP�v��6��s�<�Ӗ�?�ѕn�]��~-z>��7�W�3E,a���7�m�9��5 3��G��H�k�d$�rA1�WHm���[����yɞe�Y3�W�xM���/3�6{���"G�G_Z���6_T��ro0Q��^�jg�f4��5=�n�f+g�=�
���ko�(y^�'����:�!{y��O��B�J=绒�����-��f���q�y���G�ڵ)u��4�F�:A��[�}Ʌ�M���
N�9���:7�9l=���JS��;wQ.n��/���8L=W*^���d���pˡ<��� ��� �L#D�U��۹L��!��٧i�C4����[�L@л���b#o��JJ��o*���)s)�۝�uڷ73�3"m��\R�-��u���^7g��ʑI��6F��ů6=š��k���� Gu�z�t��B��[�̽�N'�{������~�7�������{���o���<}~�W��<wp{���̼�=�����ܗ�d|�d�.F��a "��n�X�䔄�|X��Q�p^��㿮���=�x���g��_ٵ�ꋉ|r�F���ه��j�G'���=3��ȧg���ymu�X�ݡl9na�bƕ졢�%��B�}���X'��a�>.us�����'�;�l�{c�����+#�HF+:p��l�l�q��:p�|�q7�_6W�j;d��[� =��6�9Qb���>XW�Δ��p�a�O�H���h���D�_w��^��tN�"�v�v�h��
�L�IQ�1b4B&{�C3˕�ѣ��3�}ŏǣ�F��"蛊?��:��ֿ{��DyJ%�q[Zi_p�R��Xyid$�Mel�9�;��/c�F�tR�:���V��嵒e1δ�
���W0�wy�������v�5�	�eX����Y�'O�U��X�"����
h�
:�� %�l��h}�z�-��#��6�\�h�z��;��wZ�35s��^�b����ɣ�a�h좶��'�Bjtm\$n:ٗ�A��pFV�9���*V�y0$�z����-�ɖv*.���ys{����s6����b��I۴�c��D����L=�x/�@�LR@t^�r��w��h��W��l�k��3$�[8�n����79������Q�g|a��!`"�˝�Cׁ��S����~��w;y��˒t��A�f!�� nvY��(*�^C�߇�7�X�#�/:k�.��θT� v�,�q�s:~�0`}�ƭ,��I��2�k[	��o��f�ʳpf	��R�rݗ7w���^����2�!�=+G��]�y�QC9`���T�xMhggҬ�ƹk���M�7���nb|����l�^�kCo��{^�j[��m5d��c������sۆV������bw��+�I0�8Rx�"�a��8����A����[���{�}�#���+.$��A˛�����[qА.�]H��ʴ��ɚ1�Z�Y��l땷���U@�f<}�����4O5�LuE��Î��U��2���Ң�;�F��D(�ǘ�v";n���j�ۈ�%r�;o�
����޿g\��
�X��{>��/N)�Ḕs��K�NoWb3$�����
��HjD�쪳X��dñ	�.�R���p��+�Y��U�Y�ͣ6îrhP)M���\)��.�]��������n�G�ф�ʇ�ۯ���a�^�y4������[d���żX-k��6�c�#���٨ޡe
���X�hk�G�L�n>���&�>�{��i쪃
������E������Q.S��a��}���Ԃ&�_P�5RSk��4Ŧ��r.S[�&\<R{�Wc���T��w2��;Y���1ʮ�9HC�;��),��}ܺ��o�G�E�sI��4�<�!Y'$�w�J�WwU����`���:SLD@Fڧ��F�AAFوu��61�a��$�*�&�i
6çT�Z4��18�)�j����`��6�D��֒�4���
hiM��4q.��ɤ�@l�iu���CSM�T�AE�i�Jb6΍m������T:t:"j�J�A�)l;e* "i��k�!DK�֑�f�:le5kiҚs4h3!��4�J֨l�&��MF-#Ak#M:
@�:J].�W[j	T���G�~�2N�\I$�܅P	A$S�Hfzh@2g6�>�g��Ec�͆1��WY�+.�oE�ӽ�L���, ȝ�P�1
�:�wV��ٺr��QI��iC�!��(��$��i�%.%fG?Qq�L���ٕ�ȝn�i���v�@as���i+���=��WC��5�~�ܚ��JO���*���=�x�P�;TJ1*�����6�A��(o@#zMdr����^���n�C.x>��3��֨�\Q3��d\�)>�����И�e�k�h];0U0�K�#r}�ԫ�V���}��&8�ona�cw9��u���p�k	L����!(}�#$,��m�_�=p�����"���~]�ש���#sЮ^q�����³[8�Ѱ;#�a�ps�G[��Y;�/o� ��y��JFϦ��!�hB��J�o(�)�̦t#���i�ڳ��v�w�Q�Z�ȵd��FK8: �e��t�<f��c��: ˭xQ����P���iPH�H͵"�l��p��՚�!ݯ�w��vs�\3W��̈VUE�������t��ڠz�|g������Wuj%�lJZ�vl�Q�6纺�x|K�1�"}�U �v"Z���+E���QN�R�?����֢JU�[h�Ӥ�B�~��[ͫ(�0�t�l�~Щ���]�/��C��{WA�`�Y��xk�i����Æ�ؼ�d��Ze峌!Wu�<��s�â��!\�;�Z��l����e*	KW`z���u}==�$u��X*���UB*F�p����0ٵ^�فo��]�N���]�FiUu��)��uө����[�,?�ڝS���D��x-�:P����\�z˞#`�]^&̶cǶ�B��^��ҟ\���r�%�q~���c���_�48��a>ǖk�d,�st0���o٢�־@U�C��u�*��Y�l�ɱzg�lMrJ(��.�,Ó桒`��]ëk�U�y�"��ת<�W��WA���ʣ�H��b���\�桓F���L�2FT�<F+Cy�G��F�@+���`j,���>C�/5Tݬ"{�W/)�;C$m��0�๻����:���u��\��YBr���g������"�����l�u�3�z�x���껽�&8�C<�km�w��f�`v�{Y1�aX]|W�cVu�3p�8�[�f��Nة��oP��_JL٠�R� =���m�s9��i�E���7������b��Un
¨�xӋ����tUb���L�W������0����n2�c�!p�R��ŭC�]�
/�?��q�Ih��G���!� c�~S������Gt��Wp�^m�5yd@č+<D�<��_mP�+�L��v�Ut�_w������w��*�2���Ǜ�ve+�)p��ͩ�C��=�ν�cW�*��t���T����=@FE�J�݄���#_ZN8��y��	j�yr�i�늉s# �Ön�V� W�Y���w�{�_unj��'(��IK�>��hA�TfH駚j�\��E����d�#7g�}�3a�=�F��T�R�P|��N��IƁtY�D���.l�_�e����(�$Jn�O:��/tyC	�~���uI�)�Uӝ2��#��ڕ]���rU2��mIo>�hu5� �����;����o	pK'�A��:�3�;����4i.��ۛ�5gr1�k�z6p��pU_�r9~qVGi�Վ��9���J	��E�l��C
-�Fu�,�q�ZZ��Nћ�]�+��2c��`r�s��fr]ʤ8������f�'���+��]ʯ��X��`��L�)U�4�7f�ܭ9-f��g��/qԘ`�q������ѲU� �x��inNf�h7m��}�橍HQ�U� ��a����o��ڢ�o!��K�i����O�5�e������Psڼ������a�n�Ă+� H�T������ȵ��>��5��J��E7E���_��w	�����:����ʽ�n���{F(
�F13���d�4L�H7��v
�xvު�4Dwfr�~��P���{F�g@�eF��x�����#&��p��#�9V�!.�J�������M�$���L��0�*�5���{���q�����l�� }���n:z�{P�O&�{jk��F�?�w7�k�6"c��(�v��A�n`�=����PSJ�]M���Ĺ��p�=rZ�ڹ�̃ss��Ld�-�*�u�*2;ӮB�䑴�P�� �2�͹���O���"^�
�t!��q�P4��X�+�%~�T��]�͡x;��?Rx�Ο��o�VIFӟ����^�.��lJ�63��^B�a$�U��:8������]g�����&�ENI���Y��X>Cv�E�o��]bj�i�[��`��-���[ň������+������0����a���;�nAN�F�<�B*�>��F��֙Ra���U��C���7�+)�!(�b m�ބ���ا��Y2cn�[L��u�������ۿ�6|>9��%mO�����;�R�6ԂQ��.�[�Zzo4�����Nkm��A�d�5l�t����j�J�gb%� �v��.Fw�MV�2��O����<º,�?��me��K�퇭����箶�٤�v��%�x`��KI�������m�6�{���N�N�#'��̩��4y.����O�"-������lV����5��x�O@�z| �T�*L��>��;D��
7xE3��U����g0T�58Y�-�sd,�v��G���M�'��A��b$���}z�� �O�{�<�h��#�0#�^��%�����;4�ӻTE��LΡ�X���?9޿0��q>�el[L�^9�5�<|�W���O+Hn������}�`�x��-K������Z��~����ˎG����!4ۭ{���7"��MdB
��w<3�:��\q��[9j8C�Saм=կ:*�ݷ��I��:'��W"��E��E9��q�Ю�?$��,���=�6�{����qSZ�cw�*��E�Ք�lS��랟<N��ꌇ�1��������_��(D��Ǽ�HH� �J�H�O�Z��2��z}�Ǫx�Z�4t�U�a�l�{��
ѯE�J�WҎ�v�V=v����ߺ�∩�3A�P(B��F�R��CjWH�T�9�ӑͭ�˳��F�ˬ�fN�w��O�=o �NEH�������覽X�mW�z��##ӝ�!��*�$UW���]X�� :B�7%�-�3:��<љ{�-�,���$̸ͥ��&G]B��^mׁ��!|�o`ӁE�,�����4���|�G<���h����|��*{���N������rx�}��h�� ��=����g�kbErJ+�wH]��ovb�L�r�=sbt�7w|ʾ�ESF�gw6�Ej�Y2�5��,:�\mS�N���D�C%�Vs�1��6�T,S��Qu���v��|3=�sw�����lk��UW�g�g6*�o.ЪK�ra囤��ޕ�u�Ņ�ԮY�N��1>yt�x�vm�i�2w/m����C��8���<ú<�q��ߨ�D��<�H
[�2]���}���oz9�R�r[�����3a�pQ���#pңt[�f���#�u�k�m���;�U;��N�m�o�p]؎�[��lݪ}jg"�Cv���ē@�ʡŎ���l�<�G3�N�Ks��![�:;��\
��C��˸t��z8w:Ih:(���a!�[3�k}���g�v;X)Dm��	O�*��#��W�������U=�1pS�.�;�w��5�{GO�x?�Wy9r�f;D���A�%hGOo̚���޾k���`����V�GK?���yꧫ�6y����,���(�t�{NS��\�i�J�m=p*%��� ��0��բ�\ls�R�����f�=�1 ���zM:����x�� z�u���0�s�)���j4�G3�ͅ���^IVl�z�1�����V�g'��j-l&�c�/�H��2�$(�۾�gG����#%a6�0n�v���a>ȵ�z�vo�����D� �B����������s�-=���� p&óc0ɻ��W�G�o�������S�ܷR;1����Y��n{ʲN.�J6�a6B�C�m��ѻ	�I+n�>+���;;���0o3P��L�����*�|c%�F�̪��J�i���R<�ns�{0��Ov��s�c�BYn�"<���`�J�G�bK�5qw��{ۼ��e����$�I�u*8�l�0����ޡ%W��/]�+�r2�֣��;*(�� �]�
��{���<�8��p�\0+�m��|+���h��"{��ʩ{{�P0�F�[C�u%=�hl����ݛ�d�?>Z�h�:}�\a������xH�~��|9��h���Պ����bwV���SQmN���z�g�Ty�Z�#�������&H�A�_�8j�gz2g+tC�^`�4�̘g'��0��M�6;�E��p�{}�Z���D޷��%���#�͚����XyA�u�jO7�݄S������z��߲!K�| oK�{v#���Z�v@���c�&&�u�=aG>
���V��a�ع��LK1l����I��؈I��Θn�PoTo&�2�@=F�� k�]@kPJ�Iޥ+Vl7tK<�fa"���ȅ兎	�5���_�1Y�=%#f���s�'�eWb\)�܋��;@�F���4D�O&�/mOE>�P��	C���
l歮a�/�Y;��:q�5�▝AV�%�ה�%{״~w�?_!o$����z������!�X��wX���A_$z��B\���TӔ3.�&��]�dc�ev�{��d{܇�5a;Kr
t�4N��x*B֍�����{ui����>�cL��Fd%��r,m���t����b�V�i�ɋ�أbvg��l��um�O�����pE?�Њڞ
=�ˬ��k���7��M�MUM���EXn��wGu��q� ���ץ��dn:��2CX��T:ɻ�tg)�_�ޓ>��L�kly�t�,�`��˦�Z;[�?F�M%��;�D�x�A;�������{��������Z�3��������$�sS��tC�bўN�O����bk#�Mcޠ�c$�[l_X�u:�!4�/��,�{
��Fl�t��a��F�?<��&U	������_��5,�`������A�{�Xf�`��#ʧ%ʽ�Ӱ#>aC���Ξ�\�D��]@�j(*C����U���w�W�����/��+Ճ$���5)#r}�hל��φ�N�զh�z�yu�_6:��n�`����6Ctjg9���2HY>�-�؏]�i����k/gy>b��v���h������3���Q
�xl�I����6L�7����p���3u:�$�;b{�].������𮳳M�O�A�s��)��<jz�tg�j�^�y��@�BG"�+)Hا22[��7.��:������}�B�=B&�V�d�JBEr�K@H�H͵���0�c����'^:r2�
��Ǟ�%�Z/o�+�[��J;����`9X,s �4F�ު��H�d���U�mȃ�5j���@m@��V����f�设�9�y���2��X*���T�R7�?O�����?O������~?o����{g�_��r���Ҭ��(ex�Q�{�����(��N��,Ӛ�,�R`�RE���b�ˋ�ux��/�.�'V0��ϱ�*�w��Eܠ�0�y)g��Ù���keF�5���� fȶh�`�ڛn8�9L�'{@�,�˛�6�ci[�0%�͚I��t^����kӢ�7�sn0�*i{@��7����v`���V�=.�+���{����6�2Y�=|fvs��M9��5��.���4�O=6�n�쫫�}�e��mv;���r\��rb�YEd;V.V��#KAK\:�xboo6��u=ܲ��*�;^��^L��x�(�gvz��f�i��QXF][Ws:�M�ˣ�]�o��?g���x!}=��97����x-޾���%8��u�� I*Go[���/�j�����l�g/#�r��"}3�;lU��n�˶�xt0��2,ufʌ.o��u)�I�F��A<^W�)�#c[��+��מ��.���fzy݃��ɰ�l�'6���xwr`�%��f�]Zt#na�6;o#�`���Q�̫����Y2��ٓe��y;PK�3[�8�ܬ�r]�ʖ�vb���pd��vU�p �:[�]�x�!���+!��S���ifr��gJ��+��"�����B'aQb�{SVZ4WV���öM�9.��2_Nsic���nѰC�m�c������Yr^p.��ֿwy�ͬQ� �e�O��gg:X��^�ߗyE�x�y\��}����)0�7{)����yQw�F�R)�\�RiWz�d�X��m�:�т�#�e�t�J4��3ԯ� ��^l��2�����sRق` �sCO+'���;>��כ���S\��W}�=� �����UhuVh-�T���w��k��N�HO�Ѷ]A��;��{g��~�둞���p�$����I���`��r�@!�o�P������!F+��ܬоӷo�bf��dQb��5v�|�"�����^<���!��ۏ �پ���X��{�~�k$7|�S��*)��sOX�ܷA��M��u�9ð��mhE���'�Y��t.c;.�L�uB��3��o�j�D���&�J5r�ѽ��:7]v��߈�kg��v	�z{�F	z��Re**YqB}�)�N�8�Զ���F��l,�v ����k�ݮ���������S��Fw��z�yv���Ćm���}�i|Wb���]�ª�����%��.���׼��R�ܥm]q�h�l����Vؼ\j�ݶw�t�����^;ԟ*��Is���M����}l����5OI74i�G�����EOM�1c�
��`}���^���;n������$n��A��j9���鹚Eb�K7/Y��q{R��{}�z$���lO �N���PhKͤ�*}��G)���篜��狅 �/��-C�M��K��N�tٳ�(��N��-�Q�4sX���)U�%(hM;`ևIHLm�4>g�ļ���ٱ�:4i�8��)Ӣ�k����L[s�	C���bm�
�V-[b�Ŷ���j��Z֢��(�5N����k�G9��yj�����kl�j6j�h�٤6�"$�Q���@h�+Q%8�#m�b�A��lZڭj ��4T�ѵ��X��62�͌�m�:(�"hvˢ#Q0C�"ؠ����[b'Tbi4�cTV�E5�h��)�UN�/9�<��U�Vڒ���cӇ��K�����{��-��:flc���{��1
C�X�^ݕ�M�h�����z�B�k�x�m�睚��m��rv�x$���ESuuK�K�"�ΐu})b�m����'{��v�I��%>�/�-�\i�O]��#1�m�P�m)�rl�v���|�=��;m͍��d��i>�b��,�levJO|ԣ��������ћz������X��j؃������5�(����럡��?�Pn�`�ϑ�ߛ�!>���8��.�9�1���I�FUx�]ϙ/�ӭ��nS�9��dI���&�&Cs��a��`�#x����T��^5���И�n�ν���x�-������>{V���J�./ޡ�`��O*2"��Զ��hL�_�O�[Ŏ����׍u���ҕ�s��p\��`Z{��؜�Z�LZү�t���øq�K@:(�G��qK˿��	�o�һ�pDH}�B����ث&�M�;��y��Ə��Y_\u����zlnz\Pt�%+�!�a 3��]'':�칶㻺�g��]�L����܄��j?v�^j+�Z9���n��{b�v^ج��}6�w3���.�D�I����<�܂g���]���ys(�ڳ-���]el6�[c��#�!�c�
6�h�M�]�:�93[�̝��!�4�(�/;[�t����T硨��=T�D�ꌋ�iT�kN���/7*v�t�m��<GM*��i���\K���qb;�n���2�n��n��?9p��FC�$f�I�:��ftKԿ���R9�eF�ܥu;��ti���o�jH�/	$W<j�-V�˅��g��0������狢�s�H\�Bm�X}݄���$�B+z"��6nh]6�٬�՛�r�b1�6U�u>��C���lm�Tax�\�����z��i�Ɩ��v/WV[�zzXc��X�p�Y��ؕ?R��>�uOe=��G�w}��OI�y��н,'��v!�oTl��&���7}y���-���k׋͹=Ǖ]�+ʷMǷS���o��ս�5t'���x�r�G-;�Vv�˶�k��;7D:���&��9��U���%���˳����A��{ڿ9�����c�n��w�ܺm����ه��4l���P��#A�/Ҵ�Tr��	�]�����Y0�7�.��_y�]�����}�s��nL���"8(M���DF,��U*B�V��=ԭW-������x�Fںf�i=y9{�˧`&C�\y�Qp:�e�*R4��4����Ѳi��n��5w�3�"������5��P��#�� m�5�L�H6Z�M�l"�XEn���c��ܻ�;j���d�
��x����w�彬�U�/�mDf���BK_����_6>�_}{*�n��=�\���������v��;�z��g�v��Y�S��S�P�����x�{�'|�au2�����u�&:}��ܖ@�J��.��yjE�^�^��di�K�X����^�A����ы
�Ȍ���J���W�u�v��p�o���?1z��r���3�v��μGd-���Dj�'�t���L"O%u�94�;:�?m�t�������1�&��Z"3!(�b#�d�BJ����{SS/�%����R3�9�Yh����k�Z!FM"�j�<�&���cܶk���3y�c�)A�tVP=Tkel�U�����&P�`EV����R�Z=�
c�:h�6�ŗ��/8'�t�t��%ڔ�kl'���ѝ5��
�<'@1J9�R��Tf2�v�*T�r������},���Z��?�����l���ƻ�MP�Q�=ʚ,q�n�r0�*�T�B����b��A�e�Q����ܼ3R�7���=-�*�'6�3��Q�a"eq~����m�����+���Ǥu�i�{��4��iڢQ�W�$����b5���(<2�y�n�I
�b
�
��i���@tʟtu��<�QD��y��zt�s�i^�]�<�^o�?���b9��1����I��k4b�q�S�d�ɡ�7��;dOp��}СG�c�6��g9�E���W�p�k	���O1�P�??v��6���@�S ��#�6Gh���Ϯ��a�YcҞ,wh諛�9��6�O#�@9?q#A ���(����-�0��zA�f��X�t��jyp���t��\�W���Gݾ��M�hhO��VR��r{|�(q��U.ZXG�V5�UN����K��i�f�wC�vk�S�'*�]~Q�W�.s�4��V
�H:{!2A�u'N0P�����B[E#�#�gl-��nu�1���sn�����	���g;6)5��cN�ˬ2LY/;��,����>`��Ps��Cq��HMr|M%~���]�oL��d+����cW�2�vY�+�U�ܺ�v.2|���8��&�l�;�m��͗�}�-R����9�(2
�P��x@հ��lz#D�F��_^b��CY(�FUB铷r��Um~�]9誖:9٩�Kl�"�89��\����Ti"�����֜�c�d�ɾ��j��i]�빳��c�L�]>���(��\kͲdq�����|�)�j�#6v�'wq��E����v�^�x�%MƗ+O�5�C�=�q{�s��ne�B��[�� t7�fWP���b��Z��U�J3a�|�
�Flb3��'���.�˯��3u�G�����{}�x�n䬾z:"��s�{�6��A� ����3g�o@pQ~vwƪ=>c�m_N��r�0�^\<X�X�2a�Fv٫JI��Rp�ׅ���y>���ݭݼ�G�!�5�Xh���V�EN��ۛv�,�k`皥����}���w9G���.TIar��b���i��AF^���\�E�râ�MWG
�vKW}ǖ��?Q}-�	�����c|���D�H�Wb[3���!װdr�>]�h�x�ʮ,vI���g�A�t7{b.��=[��S��YZ�'�Y���#�3���f�w�r��^��ðY�K@:(��y6kV2�׵6�u����ݲ�'"��dlU��{זDOq"J>։c/���;�z� �ocv�r�U�n�CX1Q��F�M]P����:${o�Tٳ��#;w�z� 	��ʺ3��t5�oHK��z�l���U�
b����ϧ%���9M���PT�	v1꺉s9�/,��Y]6'�봷L��[�j��rQ����+�H��B��{2GM<	����sy�rg32ݸ��.D��mn6����x$T��M��/��ډ���{s�S���5�7D?[��Wd�(CP� �6@��c�}�Q�t��7J�o�pC�7C�v�T*�N�rmwr��c�Y<���|��/�$QSHa����9��0k�GXn{=�xdC��(%Q���sӄ>��[��m�
 �EC��h�"��UL������!�7n 2u�^�#���t %fe=��-��g��{F�Agǒ�;yb�g��J.����f��=#|_k$5ө�q�d����2��磲JX�O�ף��'�]���;���1�#^\_�:zCpK�
�~�GY��ڮ����g��ug7g
t��$R�����B�����p�6@}[�Cg6�p2��:b�	~뭸��27U{��Z�P�wMϷ��f0r7D�jg�k9W�:ͼ>�oi�ZiP
�՚�V���hl���7����{k��kV�Ux��B���u��.�ԍ'��c'�5\�Y./w1�s��:�.�dh�:	�B�}Q����\I��������G4wX��|�8u\.:#E�xThd�#%BWxC�~�{��,g�VO�r�c���܈�[��y~�k@�,��ZXfT��p5���s�M=�M%ݑ�Hyǧܨ���M7�������3ǥ��fa5&�~<��"Ӯֹ�#�z%y]��2ݝ=��/��,~�H��Zi�cȽ���1؜��@4Ap�G,Rf�{A��!!k�wR:����v=�V���;�؟��d~7�eCq�6V5F��\xN��8=�k�yM�{d�aɞ3�I�!r�nSW7�k�T��]�Ve�@MF�\\�4��uJ�[Mז�\ӕ[V�Sv9�-u7]�r�K5[7�Q;�?
ň�dFq
�y�P���T.�{rªF�J�N����SN���뀲n]���\:<��0�i�y"�Mz��p��]"�iS�66��dU�������%��X��qZ���}sƥ+�ލ���#�a��x���t�Ey��[���<B��m������'�c�{�����t��7_���)�@��<tS��E��X��=�y�v\�qJ8�M��z���>\_�#1��w�0�I�f�ɞ�ϴ�gC���	����Y$��JY�$YݐmvL���SfE�V��x���ŋ��p���z�k�T�u�<�Q�ަ#������E0�^���-�؛>X��#�!�mφ���v��4�9Z�>�rϊϊ+��~O�w�"��	k���WX����V���}p�{ϻV�{,?}�F��~�.+��������ߜ�qy�Og�Ə�g�H����a�jg�u*��ZrEQ�Bj�b�%�'������z��3�Y[*>���	��o���Ov�NI,�-qY���g���!�7�Ǝg!�ryn�ɺ'�o8��nw�}��5}�D��{�^wF�h����� |;�"2��Bq;��{�b��������ۣwݖ�Gq"|H1᧚`�Mt�c."c�墈7=ٚw_�!ğp�d�諓ݷtC߷x��V��D/�����xy{���G����Ib?�2�bN�Hעz{q�5$&� �I�B��[VN�j�����.X��2.��5W�ߝ�(B�j.2B�e��,�5�y�NQ�1]cw��㶨�eĹ�PdE;(�Q����W=z�ᧉ�6��ܐ�C
�#)RFUB�;UcU���q �r*up|��l���YpM��J�؅�zG��49��%Sx�H���q�u#x��Sdn����.��֮��4�� 9)�����IX�\i�O\z� �o���ُ�����j"Y}w�k_l��)olM����Mr����Wdp�5oT�7����{4X��nh���ŗF�w`~��!wfy{]�5|�N$�=q�n����۴}'��j[�az���C&;�+:ά4�ex��]���WQd�	X�/��9Y�|ԅ�\y�[ F{�@��#m<m���*\�j1N�4�_y��k1��y"�V�w�[�ޟl�R6��stKu������F�����4a}�����G{���k��l0]�ȍ>�_,U^T'h�[¬��rGfF���&�Q�1F�����1�F�8(�S����%����ݣ]u���Ou��2v�l����@���QS/Y9��8u{��wd��vN#���*�I~ög�A�;������uv��4ץבσ���P�p�9|[E�Ѧ{���UL��6�.3)V��y�:e�]�ČL*C�1煳튴ot��R{�߆�z�.�q��뺷y \���G�m��R40!F�ݣB&��fd��������Z��x���N�u��I͕�Ԝ4� ��4��N�>������^����=�
�
�� D_�?���P��E~\#��<ϓ��2�ʳ"�0�0,��̋0��+0,ʳ ̣2,ȳ(�2��3�2�³̣2,��2�ȳ�0,ȳ(� L0,��*̋0,��
�+2�0�̋0,ʳ"�2,��̃!"�+00,�3"̋2��3"�J�3̋2���*�02���2,��̋2��3"� L�0,���̫2�³̋��PL L�0,���̫2,�3 �0,ʀ�Ԩ��A@�U^�"0(2�0�0�0�:�2�2
2�0�2�00�2�20 0�ЀUXe aUa� !� !� !� !�U�UVK� !� !�U�V @UXeUa� !�U��aર�q� *�2��� "���"� ʳ̋0,ʳ(̋2,�3�'��̫0,��"̫0,��*ç̋2���� L0�ʳ
����Ǜ�h"
4

�L
"����������26t~N{[��M����?����pC2���=}�Y���
 *������� �����H�����a�@��?�_������pPW��~�����8����	�?c�C��{�����C�_�?C�DX�D�
P(�@B�%A�%�%�!� FUVEV � ! @UYXUY  �!UaX �U��  @R  ��U�UfQ@�$�@���?�����(�"�"-@+B�~a����>��(;�ߠ:��z��aPW���_�}��sПä����ǃ���<{�E ~�C����c��ޞ�W� U��~?��"QUz���=� �*�?��&��|}p0`����N��z4���:E o���������
��{O����#N@���<Hq�0��@��I |�'�?/�"�
�px���I�W��1�`��˃�?��^��=�	=~o����Q0z}�2����A��OK���;_�ET��gǓ�
�+��������?�2�?�b��L�����	�� � ���fO� ĉ}�>�F��5�k!la*,�EHU��ajմ5i�ձ���U��l[jT�MjJ�jх���2F�!T�@)U"
P[2D��6�-a>�Ͷڡ�Me!5��f�l��Ŋ�*ҵ���L5����ֲ��T�Jkl��c3-ڶ�J։�kJ�)+m��[af�s\l͵���e���(i`�*Z�+�34�3kle�ٳm�RSi��[mmQ�m��dZe��6��[Qa��+Q2֦��cTFUm
լ�m���5iYKk�  �[kv)ʍ�giH�kN��]���ev�:�]�+�-Ҷ�ku�][�ւ�]�\wn�Jո;@��R˥ʪH���Mqv�k�)��4�m���՚��a�؀�    Z����+M+B������>���"����-cwx^<���d�}ؑlP�����С��K}���I�.�hͳ�f�J��fw,�p�ږ��R�[�S���B�q�5��wl�n�ڱ�ʖ��kL�e�5�   g��=�M;��ڔ(*Vu�;v�ֵ�w6�]j�;���Wm�S�MݗSJN�]�Ε&��l�g��m:��q����kmmۥ�Rh�v�36i������հ�%5�   <+҄�3�ݽP�e�2�Gf�h�]\�ĥ��n���kCw)]����ѷv �E
��q���`��ݵ��nE!�C ��h�Z���j�[K�  'x޳�h�1�
*��9B�Z:�m�{��\9�Y�k��	ɝ5GG]v����u��֨��շj�+76�JKegs:�*m���_   ު���k�r��V�NuP�ʌI�ӣ�{��b�'npئ�\P�i5ӊu�=�{�r�
]�m�Z�L��٪��i�-mfV�mU��  {v�4ս�p���n��ή֭8jY��v�s`u�g������uT�
�O;����RB�O7�JT*J��a����lٌ��ԙM����|  1��U��BQ$>���@�ֽ�vҝ��^��+٪��4QAΦ�%GCUoy\ץRBS�����C���UE
��k1��훷���c���  n�|�*����=u{�N
I{����v�Q$��g�AU*�����!J��ʢ����w�z��0���3��$���u$H�U��t�B�m\p�$b���i�m��6Ū��  ����UQR��׽(�TQ{�R��X;���K֕R����PT�ν��%�/q��P��Q�*��+����T�Qjz��R�� �~@e)T& CA����@4@��BR�� ��!��I  ��ڪ�a  OT�I�U$  1??��������I��&��Q�3pM֏T����Q��+��r��8�功�_}��U}_}��o���v�j������kk��m�km�u�ڵ����ڵ�Z�[mm{����|����+c�*��I�c�A�r���933t�e�D���+L���ܐ�Ʈ��>��Cxt*N�0��_aV���tt��u!��û0�֡C*l�@9R9��� |I{��u���M��q�$ѫ��Q�j��*�Ut*��&��9JU�kE���e���+(���p�؋��C2��cX���B��j�mq���X�+�[�Y4��2nLzN2��f]\�3P�����`,�h&[��P%g_̋CpmY)�ұt���b'Lz��Ⱦˢq�(�/%�-��Q6%���ղ���TX�xp�ũZ<�kw��&��>���qZ�JŸ*K�Uf!`��+�F�RN������;�/o j��x�M���Ach�F��pU�9t���)]LQ�H�� f�J�ҫ�JPJ�q��S�6�Սἅh�M�w�!��Ws~�I2 na l��Cn��ħ�e �)ciP �˚a�+�7NF	�`U���י��hZ)��e�I�*�Do,���	�Y�b[���"h�`��i���n4�Q�ǈi��N�f!�sC��I����`�#�)�1J�a�o�N�4F��z D�f��C+�/1��lֱt s3`,�Ljl-������$
��� D4�A�sK�7��z7%C��̗I��[��6lVM!`f�-
�`ۣ��`Ւ6��J$n�m�2�
J�����]L`�R-Y6xf�h�a/�>%1+1S���A��հ]��ږ�X���j�bd������V��XQ���4\*=J�L�X�a�2���(�rY�b�j�r7w��&w.������68[�On��Ԗ0���+ ɵgq����9f�JV�,{��ʸ�T`��FZ5ɹJ�"2��`�,cݚBm�`F*��Ar�9,����x���r�U,]�Z�
�nf���y�PM������-�e�2���4�@�m�#&e"�J��]A�ѧE��(�\/7,A��i�/A���"���	ӶA�;��r�4���%�[Q4[����6��5�n=�4��w� e�E4��Kn��.���$)1Թb���[�Ӳ,��x�I� RD�TyCl����Nd˘����Y-f���d�	0�Yr�LVE`�sn��4	V��:b��a�pYL#(T7�d0]�<�E�c�ۥ�&�B�]���i���8��V��g>W���u�)Պ��r+օ��p)z�j�a�{�2mE��R1N��5�&Y�x�<;�U]�]�c�q�6%F�o셬�n��g�Y6sZ��*T�G$���r�Ïm�У�V`��6J�g`�6Ў�S�@ᱷ�RKhd�B�b���0;V�f�ܬ�bVf�{�M`�����+,�V��D�!pdW�[�xr�e���d' � #V��XHLw��`E�"�R{��oqV`���엣f�/<����dM�I�/XI��4JeL-�vMi��tصaa�/���i�-�Z��6ҩNY%�gr:�Ď�jc*���o6:h��aF  ��|�;.,�x	�1�33�ƓJ�>#M۵Gxg;;\�*E��ē����]�SPx(�$�w4��^�cLn��ѭ8����AA�6>ˏ �@b[����J�2.��e��N�5�%�Fs(�v�h�ܬb�X��(��^�J��CiO%�Pu���ƲH�/#��֠�,��̭`;.0T$��)J�%l)�n����C$`u���-)�,)��*���H���T�2�C�{Ov��7Y�)6��7���A�F*���2e�1дnP(	e�yS`�B�fb�&=���F�e�Bn[��jSo*̴.-����ݹe��{B��2��T����7���n����i�d%3A��F�0b�X�&B%��� �0
�)�7��ז�Ė^����D��Ե��qmIJQ���riW���8�n�[�tXN��/Xb�`���=ڕz��6���˕s.$sc�3j��d�)���(��|r��,�Z��l^+8��O�h^j0���&&+V)��8ay����ո��5TԴ\��5
���s-�%]�9p&5jb���`�ec���݌�!NG�m�A���^��MU�6�$��E���1}�om��I5��e�
�D���l`*�6ŵ��i�9	
��v�;�$�ٺ�����D1d�i�U��^]�=��Pxj�.{λo�#%n�v`�%̒�G�hմ��sJ�=�-vjM.L�Yuן5V��%rV@�I����e�F���t2�M�S��I�v����ێT�;tD�b��C��ddU�C��a̬���U>�i��X�m�̽��3��H1�%��̘]�b�ft.�´TB5��X�5
:�:S�[��н��1j��m�7j3 ,�!R��E�J �vp��B��ưu��p
��Ʈ��������S���)zkn͓�!��6�"mڽ�V����T��쳦�6���d����K��`�e�\;pe.�\�W�vR�k�,��f���HtZ�+�L��!hi\�� ���N[sc��35Id�h�4�U�n0[<*/�c8w0c�M�c8K8�F�\V&�ƌVw9�`��zr��Ŗ���Dl�,#?U��)h<K6U��/��p�d��D�0���d:�ج��4f����CѪ;Ʋ5�☍[sR������c"NS���s��,)Y(1e���Qq��m�ܹAC-�<UȖ��ОF�4���C7�Ɗ���K���2V !��-��X�cqn��؇U�����e<Ba�t�K�Y�b/�؜X��R+&B�=��\t�E�M�<��A=�[�������j��(��[��H,��!dE4�vN
6!.�KP��.]�u�j�d����l�*iV6<nbm�A,b�2���,��)����f�����hdB�+̀��t��y,!_1h/��CG����p2���� ��˵�V�9X%xM--Kh]���]�ANB4 d��^��M���Q������0�}k�n)[y4`@0�hɘP���o��/N�Ue��蚭�n�л�$�/��W�n���g��K ՈQ��9��C�OM�x������Kh][̷Z����
����x�E�5`�����#�2�(Ц���Jd��yWlծѬ7�ۖ Nm�N�
��£�u��I#���5.�f*�:�EC^ �r�AS+�a�&ݑ�,��ˌJ�[���)��Z��<Tp�-M�Ӈ�)���%����5+!���
�i� ��C�����iC0��#8n�ʤ�jn�
����)7�&����⺄F����L�ӳN�zY{�xvBd��n�b�E��kl�݋F\3E�n�0Q=�O$p�[�T��z������1zM�<V��9j����BT��X��Yo+e] ��W�)&���{Oi�,�K��-J� *�Cx4�X�%�+�'M�F9F���U�Y�H�6�K3U�J�c�O2�( ��6짐.���6��&�<6�`f6`W �R��bZ�͞��r�55��5��l�
xw�LC&��Z�n��&��,�4���eei���8�NfYX���Bm�041/��&,�������wR){�kE�jm��%��L��XP:S����d���Wa��Tȷ�J�V�z�Ԝ$]��l[�b#*�Lw#9l[�ձ�IG6�%Zw�t˽���.�UҤ����`��X2��N���:(9�
�t����U�"��n��Tҡ���D.��g]�E[����n8۩�X��/2���1��E'�j��-��6a�m0��Q������U��ޚJKȅ��xmi�+�V���m�f�!ݻ�76�rO���"�rI��$�un���Y �ʲӨV�+*��*�Ijfm��2��P�+58[�-��~j��Kj6(j�A4m�n�n�a���w�d�
Xe\��&�"�rAb��m��.�*�(2:���m�Na�[��*(�ًZbMu�(Ɍ�t�9Dw!��a�tn��l�f���;˺7��Kr���U2�@1��[�F���,�s �+)iy�2T��`;f\�CA8�ay���10�,��@F�Rr���Ż �|��kԦH��Yz����@���U��uu���C
��4râ�����Vf�j���N�����h ��������;��uU�iK�1��)�� �I�2�z �1N�i�u2P��XpVGn���G[�q�+0��^��S��T$�[�r�u6H^k� i�.J�qY��༢����	��Cqj�Csrt�>��6^���Rk��16c��;��9��g-YHGa+� yKtEVqwa��ws���
�q-���.�te-B�5�-�k>	h�p��7,<hF��)�����֤��1����m"��!@%����N�J�-������.Ea�VƖ0��eA%��f�I�h^���F:�0��xMͦ&=�m`5 z��ooU%^��&ͣO
��ͬ���4:�ι`����qF*���Fjy���t�A��,isY���N��[ږ-i��j˒���C6�M��h��-&�
�H�VS0�!���kp֊���4n�uuo0�~sh�Z�	�R��#�Xc5��k̋R�F*�n=2�摹�|U8
�n���SW)m�$�w�k2��e'�w�� %�jM:�,�n����&��_Z��ڤ"�uVυҷ�qd��6ڛiaB�,��*����,GDB�:N�m[b�!vR�L��y�мd�]ŲL�5M�2䦝^;&ڄk.��c�B�cv��q*k�p�6o[O^*5guk�YH,�5�{@�K������ֺM��cQ0���Y�U�A*��k2�E6�����vW9b��Lr�_ķ�����(�T�e?�5R���i5����M�����9x+*ďA��{�:R;HX����y��U�K�#zsc�-
2�M`;ˢ��ū�*�AG�X)�R=����k�^e������
�"�5s�. R�Y��j���5�\VnV`$-� �l [xZE�(��ֆ�X^^�5/;��\ql��*"/r���dj\����3n�*�3>�������p^��J髻uj{y���[�3�6d�Me�S��k /qhX*��:�d+�?S*�H��k>fL��S7M%�T�p����nب�Pn��/^�V�k�A�8Ӭ����	F�゚� �9YWke��R�_mb��-�X��Q��=A#7Crm�׃M��LM�xZ���4QW[�ņdՖ�*a����x�	n%EU�fJyf����r�0a�.+%�Q��i׸��'R��C��h�$��7I�q�X}*:�D�Mhn)�,�c �`̅k�Lg5�R�aeM�+52�:�/O̒�(�H	�b���3��q���nt�k�B�n��4�X�hhW��B�����&�h0�c�(��Cw0�Y�)��CBe�;���V,��v^�6A�[�7$O5d�E@�iMyQ'��i��nhݘi�G6�]�Z?��0X1Kܳk2���6^;�RH��4 `����$#�$�-��ЂMڕp=I�d�DL֠�ö�Zێ��f�d�0�ސaN�nKۃ�7
���AܒZ�����"BF7ق#W�Ԛ�
�#���R��l&�+T+v��Pj����Z�7���.��)@v�iR+c��/*����{�ȴ<c\�&�"�1#J�n=*Li�ʹ�J�t�I���&��2����Zog�qKP7���g4G��̆*���w����%,�nbb�&�*.�ծm�� 
F$7���^;��n��M��j��+��rY�	�n�T���⮴m���Ѧk�^܏jJP5M�a��6�V�hIm����sv���ĵ	���R���g�g�P�h���^iw�<���Zu������	�B�Ďd�3>9���ll;교ւ��ƭv�����VtҗZ2�vuQWZ�x O�Q�cǺSְϴ/�c�3qU�b'�b�ʅ�B�C����4Z��c�4�I��L�]ZF��]�%e�ֶkr� �#.Lx�%�ɲ�f�):ʷ�/ka�Z�*�U��%�M��3&��wx] ����Wڨ<��8]��� b��b��1j�k-�*�׍-�mV�XA��FK"J�'8�:)��̗��l��� f�>�nf\�ua;r��͵��.�`nI*�En�$�+M�c��Y�JF�/��V;L��?aR`�p�q1��ӣY4UBV�j�-W(�[1}*`��Yoe�]�N)����d̪Ǫ���lVV���4/�Z�]�+�4�]���GZ6�&��r*�eլ�[�B�d��mҺ���ӀeZ����&Pb�NL�R]66F���a�L;U(��V"�5�0���+.��T!�ۻ�:����+F���m\��cG@řma�%S�!CB�\�ǘ��{kmV�����;���"�Z�	h���4�󎂪�ߛ}�ə�#�i9p#�h*5�KY{�	�gL�,�űI�
�Y� �G�j.�6�9����;�q��G�^Jԕ��o]�G^^&��4�U��h��ʽVnXu�C�r2����)Y�.����:�V�MN�1I��ˉI2�x�jeC�Tt�X�6��(6���jR� ��I����Q�r�tR��
��U��\#hށ&V��'� ��6���3B�4�b�ef���)7(�r�	��lwN��G�iǲ���܅�7�M��gh�Z�@�PE8������GӋ��R�{1PU��;�Y�iM���^�wwC{�*��#C�Ap��w&�{ n��ȩ�W&�	��}&9����VLn�_�OD,9����@1���9�$&���RM3����;���Vq5]�;����л&� ���'���dWV�S`M�����Z8K�s2_+�����J1����Y��E�U��x�5,��G,��$]�%������i�a��v7�r癠l�I�������(g�=���;�}p���dŚZx`;ћ���/%���@���jU�Ch[�r�r1v��]�|ֻ������9nM�W/v=鋸k�Wh��������Y�q5��-��ՕY��S��)�)tٌ(K�]���v$�$�l�bI�Xk��C�ݥwR��r�>g�K:i�9m�k��	���m�Ϋ�ذ�*�C�R�
�U�;)����#��
Kᔨ�Ξ��d=B}�4�B�
�(�{q;F�$�xvq:;� Z��짥|��Z���:�݂�M3V�|�YI�rN�&9��8�ѭ.�W�y����b���3��l��X�������{'�Ob�mMՕ��u��pN�.RB|�t��w�!¯���.�(��zkލ�R��M���F^�w5�n㜴<�'Ap��KfR擤�x�Tq�Jbl(Op:�c�h���h
HȦl�Zޜ:�Vj�.r�:�EL}�q�\�
�+��x�yR�{���',hi��a lw]��*ر9�;��(�L�vmDqCm�f�Q�t��0�lӹ�x�U����J�15��@��7v�}�I�� �c���������-WL���uz/*c�4::̭����/wy��K&^�����������w4�/.�Y�`}:���!�B����xBY��)�����r�+�)�N�T�/�j�^��Dw�:Y*յz]Eԃ�TZ���e�<ͱ*��t�B%/�����-���{��O&�������ɵ�E�]�WV+��EY�����9X&e�{�i;Wsɶ�)`e�P�[X�eaҝg��$��i�%t{;��,|�gM��}��y��]���è�t��E�į'�Mj;��ٻq���)�*�ܶ:���5�P��YWL�[F�m	`ż�)��s)�r%�-�^ԅCo����B�i.�i�)5K����{�Z�͞D.����,��yd��Y�o�U����ˮd`bTqns��sٝ���A�B�,J;{7�݌�r�ۻe�J.mc, ����3b�hx+>�U�^��,(��4�'����ʮz4���)�]��F	y�T��&���"��KN�p¢hI��+K43+U��86$Ja�v��S����qR�(���qm�8�O�]�u����|��
w�Z�IU�&l0�{C�I0�AB�:�K͙�Q�s8�pC]vĬ5�i�_nщ�ޗG��ʋ9r3�)�u��W�b!YW�x#gWL���=y������9�􆞄t����	�w
�tٗ�#�}d�]ޠ��w7jM;Z��2'���߄��8��U�tS�o��J]�����
��Ss� \�l��ҊbEq����*����2/6�b���L��n��x��2<ހ�����2��j���α���5&����<tQb�rQ�� Kp�w��W� ��u}:���+jv�ks�)Z"��b,D��xܭ��ۓ	g;+��6�K�3F�1��M�U�<�ȉ=ۈ��h�d�I,��o�;�镼��ee%u�ǧ�>��j�ҝ���mVh��&�h�,ձW�}��in�a�b�=�\�&�t���jL�
�/xE�D�4ӽ��|��i&9i�m�XWS�;�Eh�m�Iml�&����	��V���&�ˉ��E�u��O��Z�X��琉�ɘo9�%�tu䙓a�`fE��da��Ex�#�3�lg9w8����o��3��+j�b����3�(��,Nl崖�|M[N�
�K�_m
3��ʱ.����&�wr��rU�!�QP�F�-BNbe�_\�9�LU$��M�C�WD��/%�pM�]��"N�@,���a��g5֛�/&�ךQ��a�\�*e�"���N���Jk��RhV��8�ĖKxtT�MjU�(��K�F���	���$�Vw�Ѧ�� .�J[�$�ƛ��q:�q�]@���x9*VFR-n�|��ݕ��sJ��roi
��j��mro���L��Zfd�B�®|�[�J���P�:���=�.���!�'8к�c��"�F�}��@�=���6�V��w��Ě�-��V���F�S��n���$��m��QY��6Y|������A�<��Gr�<]�p�Ώl��]�8��5��:�,vd�u�.ذ��/��A  f��(+�c*�:3X�ܗ�1�/)`.�H��Vg:�˫���!8"����X�bN��4k�ڃ jɨ�r��$�vK�z�'w�*�K����gl�ڊ��[��5�Rc��[��R[qՋ ���u�ۨe=ոV��"�J�h��mA�Jk4z��aO�S��69��m���VFL�7�Ȏ��E}#+m��Q9�묩a%����y�:��d�Y>F���O�x�#�QY��=\�VEb���k[�\��Ns��n�M�ݔC��� �ɼu�v�^���9���]`��ꃳ1�$�J�v#���Hy�J�:�9���h�cј�\SΕ ��9�ǒ��Z�%�5y�t� e���C�zLd�j{q�2X�y��n�&�f':�^<�"P��Gv����툹dU�������'M����mIyV��M*0��Je��Y�G�j=�ku����ԚVyXF�Y}N�'��2�Ջ\J��/|%��^�*g��������T�Ͻ����\�]<���w+@��>+r��꼾<��e6">�qzܣ�u.�����i�8�z���s��J�$�q�q\P��lJ�s7sַC-ڗG�ǀ�Î��|���:��w˫n��Zf���OCJvcs�J����6�\P�:�����r�����Bk.	#�U4�Y}��\�:�r���'���dݬ��� �÷O�*��]Ļ�E9n��ɇ	G*��,��;�wr�=����/���h�&w��+4,�R��=3��^�y��J�	�29�d����vT��Ţ\��������X;��l�7���C�ژeI��}S�S5����u�ɠ\�+�G<W/Nm��ԑ�3Jyu����Ȝ�rә������NÌ�
���4����3);۬�?=�/TBK&^W>��˂�>@EM,�y�<���<�&�"d��؝tVV����}�^>�-1k�7��I^H�'a�@�3V�8t�`z��֣������Lf���f'"�-����g����/�#�nH�)K�e�Y �!��A��Z�P��'9.�+y1�i��N�ƹn0�71��6��}�oB�/�ڡN֋O4�^*iAV@�f�Uy���R��'� �X��ޙU�]C�̺�d��ݔ"���앪���	�m�gE��Io0єb4�j#���[��)q��yO�6�D�c�ou	�:��S���yØ6�[0B��<�szi��׾������<�]�o1�6Cښ���_QX�Y�*��0n'�8K�ﯢ7�*#��d�5�к�V�8��з�-VP�|s'r��U���j���{L%*9���x�L��E��JD�ӥ�QvF�k9k�ou5������(�_b�[}�,�ccR�������; ��3��C��:�a	@o��t8����Y�_qłtbHtM���g��Ѓ8�e��T�ŴG˔E��Bv�Mp��v�2���_3ZzP�_=�Z�n��S�����C6�����"�Im���Ǘ8g�&R�jmL��f�3�dz	u�ie�3
��M.C��(��\�8�&����-�RK"��dQ�j�J����9�/-�i:��t�m���*X��u*k��R�[��>�K��;o0���TYG��b�����P�2JŎ�ƫ�C3�	@�U� �դfL�N.N���,
�L�9���k�(<\]d��Ԗ��BӭW>���]u��oj�D�m��Ƽ��)C��}K���eT�����yb)��A�����Z�2����L�p����b�-*c�k/mu횛PliٳJ�A�Nީl 3�[Ff�YǶc�C���A3\�J���l��x��tҟW(OFn+�%g��l�ں?
7$�X2��͞�Q�;���}�Y����ͧ�A� V3��»E�KAq�o��W�8%1;�ȕ�GU��l��O��c`�Z�Y�1�
S� �{�D�+MлN�=�68_Y>K��q<�Yyڭ]c\*�:�M	�fș`��F]C��_Z����h\���"���=�5K���=bT%� �A�.���j�Y��],�u�:,���Ѣ��L|�/�a֜bY��_v܁2��7p�YL0�\K}\���7_n�2ėz���aNk����ӥe�U�D�[�v{j�]�Ǩ��o�m\Y*?�T��a�XpN����~����a��+�Pn̚&+�����Z1��uڧ��]���w�⽲҄<���9ڍ����ͅEء�Y�ܘ�v�e
�z���P\ �;h������;�[������AХG+Cę�R�K_c g2��<�t�.�b�vr��Q���6o-ʔC����������)nRU/�J��
Nv�S��g'�(���]<hV^2�PϽ(h�2P�|��n�v�@d[�gNmd��5sE���"�x�"w�T��阻��(ayvS��fPD�T�����K�V0��mFr��z�Y[ƃ��i���Qo9���)�y�N��k��^<�K��#�/f:T�h{��g����j��)��*|,�4%��x�(��gk��	���^v(��Tu�e�G��"1�*�0WJ�h��Vw�F��E��2��Yw�cW�����j��'��Zڇ.��ħ��T3�l �ht���E�Y�"���K9���]+�����[++E!x�%W���f������V���c�������W�V���fq/�2��� o8���X6�d�%�׭bJf���.��Z�I[X3�"�;��ޖq�T��3���8n�c;�f�C�0Z6nn
ẛ�;N+n^�kD�!��_K���I5R{�-�3<��r�����nrv08ئaxB��ܖ�%�J����Gn�bc���)Ν!�Q�(��{w� �kh̎�^,�C �W�1��^5�]��j`N�Շ\��&w���fqÄ�]���c�rwhU�@ۘī�| B��w"��Ԡ�j�̧/zK��aP&` ���˩R,Z�扠�!v��k@�6�ii�9��u�Q;7j�S�:-蔬�}�Bk�2wIM�WVSނ
�حK.Ws>���.mI��W}(|�kv*U��i	�݇�_8p��Tt>[&���/b4�T���D�5M22�#��w]�G��zxrD˭|)��"�8��w-B���U�$�h��{�I�\8���Yz)�&�B�X��IUrܤ�U��d,��ν"�ٗ�ܰ+/��P,�1*gQ�����]/�� �F�ՎwX֮Y�W�RL���n�+� ��R(I��v����*�R��kL-����i!l���;��X��R��ڛƲ���h�#n�7��Ĥ8�ڜ঒ ����j�����b��L��42*�6ri/z���G]L��2���9�7����fcY�;�|Uq���Z7Y�U�ے�֒� M�w!c)�F��=YXy��Vΰ
��V�c��ý��7��4��ac�ؐ�e�����ܷ�7~S9��:���#1�j�v�޸X8C�A˼NoK��$z/��&�J��FM�Aݍ�L��9�q���k��3��4�˷G�a�+b,L�����;x���a�\j�IQ(6�l�(_f�+OggA��k�>�4є-�S�UƓ��,�&��٣RÎ��9���Eoj��f%y}t�ͬ�1�x.� �.�"�uh�a��^<�.���d\��vk$����N5�2��#�Inyq�u�v��Ñ�0���67����o����%,<��dE�7�d!��hƱ�r�()��ȵ`���+��Pެ\雯Ge��5�;/9S�����2��[#��<�,Oz��#��]�w�2�-P�)53�ņ4�؁�aj'r�޵�s��ah�4�p�R5�U���2���e����J�� n�r�i������f���P�@8��L�j��ub���%gc��,�W���]�ʽ�i����K��V�u�Z�h/�p����-ݶ��K�;j�(٥.t~X{�ֽ�K;&�${��Tҍk}�Ģ��!/n�!ԁ�ڏx��=r��κ 5|���L[g�*`�,�!v)[��m�5b�k �v��c�����W^���J]��dk+g$R0ݻ��2n}6�]����
vJ�o�}�� ��`7󑁣d/D�=ݝ���2�oS �%������:�WN�S��"³����0���\Kw�u5&t�8�E�s���BV9G1����j0�m�a��ҒG�gx�ĳ�-t���V��RS��j�	�6��\ì��={+q��d�l|�zk_֖6���a�<@]�B;{�0�p�Z�)�)�ʕ��,����Tw��l��s�[��)�u�d�c,�=�!�3�=T�o�l8#P�� ��mIM�|�D:#	�M�I��Ps,q�VR��Lj����"W��E�6J�9�r�3�7�vT�O�����W�}�}��������U�V��L�Q��Gj�v�+h�K����S����rp�bp5�ns�7[eg+Y"N�=C]\7���9.�$AL�udE�z�5A���]��Hݸ)�X��	����VWrd;v�)k���e��.��W���
0�c$ݸ��Ջ:[�1ح�5�Kͤ^�T\��� �z�"*�[3n§(v%���E�f�B+M
��z�λ�BK�g0;WP)��[�E�Ѻ�����[�Y[����)Ĥ:�"AP�ZzN^5 ���g������5b�Vg��{��A�+.m�OUє��A������d�d��o�h�81q���R\�շS���Rퟲ�&(;�ȓC�t�cX[��!(�-�#6�zp���lc�&�,�YG(˩z �+-�Y����c��r�ʈЫ�Z��הL�
SPk��j��u��d6�vB���ڶ+�m��M/2��1��%#;�e�$nv�c�z���\[9ھ78|�L��V����Y�;+Cf��p����
Z �V�
�N��J�J[�dT�r�m��T��õ�1�Y:S�ޙ*�s)���`�m`�S��������z`�=$Q��2
��We*��7��x��`��%��s�-y��DƝ��>��E��"e�1�y�p5�K�1)�n�&������ƚ9c��!�r��j������#i!�ѳ�[0�K���7�G�V�zTn�m��Q�o3�׶��th�v^�8믛��4p�ܦtq%�	�F�v�N��}�ڝ�e� l��BQ���.w;����)�f��"����b�V�C![��㭒��qX�u�X��VF��P"��m�jޠ�i�	YvrgV��糔 K�s���2v\F��"�Z{��1b����Z����C��^Y��4��g+�*��*���\��	�&,���Æ8.�=�Gv����fܩ�I����ֹ]*�T5Y���P�(��A��Vwq�L�*v�1\1m��pI �S�����]��}r�
٩Dt�ܶ��X��U@�y�3�KÝV���+��Y���Y �	�@���1�W��7�ɋ��n<�چY�,=	�o4���_>�k#���%AI��:��MM�{�Hk��\y΢�*VF����h����o1D���+lf\��X�̈j���u������=���Ku�d�H�Ⱦ�㻢Yo5�5ۼ�9���P=�]�X�U�5�ޭ�ӱ�T$�MD��h����Hn�Hj|ub�[���rZs�6��[52���x��5�;����o)���|)�d�H��Ӧ�뾮�^�c���1�;��3�a�yj�^�Kwb'^��B�>d��Z��|멜�\��w��\x"ynՅ��\�/��08#N��B�ڵ�o%!Jq�@�O�wG�W	5��k��!=GlLR�
|�q����T�ִX�D���A֢���]�-�ĳR��͈��`�2�ɧ�E�td�v��%'38Ӥ[��NN�Qq���7�;d\��5F�i�S+��m�xi�4��7�7�T��Av���7��i�[�Vo�]��P^d�|��}�!�E1�v��m�����6ܡ��gKU���zA�����qT�E���@��;�S�*�\��貗A��Y"������Վ���^l�i�8�VBy�.���sn����'	Xk-�&���q��S#J�j�B�
�WN��	���2�v�w�g�$R��޳�u������=g����S֭�s\�����p�wqogg!\�"��®��Щ�kn�K��Ԧ-���OHu�mX����ќ�O�N0����v��Ħ~Ӻ$��N��1[�����3�;����lU���n{�Nl����EY]!R���/�L�l-�S�c�띨�|�AHe�6�7X��L@�۵]�Il�����{[+5���r��2���wX��KʝCz��[n,O���O���*S6Mm��q��[����Ż$��A+}Vjs������KV6n\I淔`i�4E�=G~Dӵ�k96r��8���%�;��3��c����+���w��j�5G�Y��8*9����k9�,if���pH�
੤DCV0�o�a�����5,1���)*��Y�(��>|z����g��Yi��ҏE]�5�����O�n�;kW.�r���\ �)��"@ܛ+8]!�ia�k���R|\C$���'�>�-*���8�=Aֲ k|%�j���Φ�St"�'�Zj�
�54'nj��o(��ceuYۚ3jK)��.�F��P<�!�m� S�wȗ��m7A��(e���PX���+��;@�=F�ܖvwN3���ѩ���8HYOf�����"��5�[ɺ6�b9���;F�^�L
�&��7����=�ba�Vq�,5�Gv�R�3��_QL�Ϝ	\�u��>m@k1bw;�h��(-�9W�)�N�,�9lZ���0n��	�Wj+S5�m�X���~��Pt���0�gt3�R� ���D���C)Q��w�Rb=�)V9�.WSkx�0���BS��3��wT>Wv��ua��9-�2�@5��b:8ۡB��y����6e��h$(�V��[�@�sF�L����َ;Y�Wo^��:�b�b!SD��E�ip��wO��
T���l�7Q�˔k�n�Q�Ю��-�@�%ۛ��,�:,�Ya�IKWY���u����6�jt��7��4K=���ޥ�j�'���q`X����`�U�ۡ��T7Z���h�v5�rD=����f�Aڗ}"'#��R�W�M-�Q��RH�Qف�׫��>F�)�{ٵs����ݾ2쫉v)����D��4b��:�:٩��e������C�M���hZ�+���5��ї��yY`��M:�-ǲ�,�܌d��X��V�%�k�f�EJв��o[�,��.���9.���)A��c�;X�*G�
a��@������ƹm4����QV:Dt%8(�vnk��7�S{y�]�cb6�6*#L�c�c�ˣe÷%5]����n�;,����mH�q)Wo���./I�����T ��f"�$�r�7�Rו�sF�="o�+��,�w�kw;��VP�o����.e:o�՝����**�Oy$���!�؂��u^䗹|��"�^ݣ���E��wU�r��G��X�����rq���3����}�"O]]_͌�!�H0�f��e��Y�˕�G��V�e�ךҭ{K#"�Tc�i�r�3jW0kX�ku�	X+`;Y)��iI[�ee�vΒ&۾����7Bv^Q�F���'w�@Ԯ�q�/I
��{b�c�)�g��4ls��b���'�9#+!B�:���-��p��pдy��'��7��y9�Yx�w���Po%s�V��<a�R�_l,��d�):����ӱx:��;��z{�\����B���Z�yKd˅�M���Vk�e����s�����_Z[�����70����m6]t����xiNv��M����G ��kpj��*��J�iS�h۱قE��oM�N����:�>�듢��tF��N�e�����=��ɔ��KWi�P�hS,�9&Ջү�w]qv��[Y�K	� QQ���c�c�4�ν�����3�g8>
�Z�����a:1k�.n�2�DԩQ}h��ύǉݨl@Ф��H����7�n��&���.�v"�@�#kxg�]|����7(�X�kH]D#�-dڹ�NXK(��8(iVt1�-���]�;k���1]��ݖV��
l���wq�Q۹�227�U�vs�̚�+J�U(��Ƿ|4�E�ʻq��Uz�h�af\�3�u���^����M�z�B�=��.��D���V�Ò�;x�@:�]b�iO�"�l}ұl��Q�7��4"\�A��tR���c��5�$ӝٗ4�%�9פa��U3�2�#	6�+�cK�w������g�9�;��o�I!V�]K|��9t�`�ԗ�4uy6�C\�5A���i^U��I�L�;j¹��Y��w꿰
E4��>�9kp��T�ʲrΤ5����#b�]�@dn��N���`e�k�ʰ�x�]����!3]	wq-�o�����;����t��\�P�M�}�F�h�\[��=šuF�!X�Ci��}�;�xk���K��$�Iy�d`� h�n��0��#�Q�J�H#{�A��4� �y���v�uԠ��j��&6�˭���;�Qt�m%\ Ք]E�J���!�o\Y�7�o)ʼ[F�A�x۽��X��^G��T�(m.�.���}r���� �kEP�8�����l���ZK�y��p5�՞0�H��M�fwo<�����ʦH�UѼD�S�O,RU��w:�r:j0�����9[���+�7�v՛ڸ�[�y����v9�c�n7��f���c��\l��ˈT�F��.s�5O�g�چ��yf2O���]����(�Z��|e��b�Q�����aF���4J����o���]�.�k�Z�S���29����m;U/�����[�6^��>��o�����+8��a��km�ZfdY�l�N�\k@N��,�0c��>}Ì0���������²�F������{�r�2a���v�Aj�w�+R/)��yAU�催�y*î������/~���ʕ�;��[��u��P�t� ����5��[J�Xӏ�_��KBQňX���#� �J���Y�n�v�v���k�e�k@+$�(��t�,0��W�؁����2�ݮ�,�a��
��6)��:�ktة��_qt2���S���V��u]u�c����ڬ��-Н���w�Sl�7ӂP�|�osV��*�da�f�����8!�4����]��/����z�%9n�c��$u�[*�0��䣶3H���k���19]�!b=���\W|��oWCӽ-Y��A�T�8e�WC����Z���y�h�:-:m�F�L�5.0�j�w]����ח���o��fZ]��u'k������M.���wp3^L�N^p�]:D!n��^.���W=���;�u�Z��;E���	���5r�{��2����@*���G��Ҍpk{��ɯ�.��Uq�2�Q0�u�&ڻ�.�����`�he�|�9�^c5�͵Xt�Uwh����[�C�[��&/�m�68,��-��4
<Tź�wT�H�$��V��U���ɱ5��;�V��wƷ�2�_r��w֚�qJ����W�f�BJ3e+Ff�܀n[�f]�ɕ�l�>����%iG(�鬝�9��|�6�e@�TI�]v%bnWJ��J�;ں�����e.�8�S�d343֚�.�-�J��J*�Υ�`�� Yu�;s(�a�E���V�N�Cc��a[fT�k���+٫G&Ws[����0
.�%�um*�;vF)�v�����}E����P��p�4�ycmj�aeq���X�#6�EM����\Y�,�t��8"�E���@��5��O2�.���(��B�G�	5L�5�U��PWMe�e�b�`\GV��!��у�)m���`4�K�Ca�ض��iLmc��Qc�u��8wUa�����X�lv�_f��$m���Q�� E�\�d+ԁ�`�5:��
�����0V]ش=ǰ��ޘݬa�QZ��44�U������`0�γd���ȃ����TU�V� }8����̨ە+vN��b�#j�� %SM/K��mm�b�雟N�)�V���)k5��I;��1f��w��2���{�����1����\j_FHK7�GIu�<�iF�V��n���m$��h ���Ug�Q�7�-tr�ͭ0S���׻ʣ���F^�eQ޾��96t.����,��*[l���\w�81Yo�Eۋ5��(#��4���� j�p�w�-v���o�����GWe����E\X�	��e�ӡ�3cil֚\E[�Z*���'�#�!fp���WR��R�8�N��ި-Ё�P�PĊ��\�i����N���L]�p�W<��]��Q�Y�z=m�6�7,>����qi�����55+����	�Q�sSTC��:7����J�eb�BE���-�t�6J(p�ы��ەhs����լB��FD��x�V� =����`������ԝ��Nm��r}�Uu�rݬ�01/���r�r�pއ�'Ishq]3�����S�Ҙ,a*a�`�X�E3Iux�ԃ�0\8Zx��-)ۭ岃Vb#�EȬ�����՞��YC^++*d��WRF�|�D�
����6H��w��ãx;�R�4�Q��e�חw��}����N�tn� E���nK�sV�8�	j\�Z�Ug�:��i�2�ML��Y���(���w�������g��5k[q�v�u5u{$�|�8Ժ��*�#���`��%f�Z��&�MT�
�K�M�l�@�E��x�!6���ypzN�4J�>��j\R�r�<U̡P`+)�r�ؽ;�6˛�E�B�����c�
glt�nY��H:�f�-3[{9k�1�|A@��Ǧc6�5!��Y:0I=�k �K�9�E0�}݄��g;���|���)d�ht�B�W�g=�f�y�偧�j'���y������@km�$�W�gC��?K�d3 ��kiL�{���Ѳ-vQ���q�G�tM�mf�:J��udx!���I�c/(��T-u�&�1���=n����T�)�tº�Ԓm�hCm�S0��V��S�Ⱥ h�(RΛ�M�yXӄ 9��N�l�MNB�8��G�|�V�2���H����r� �u���u�yb	d��:`����S���%pQ�sx��)����}�W���z��ܐ/W%JU�bJ�)b,��u62�׽D��L�գ	8#ˡB��R�$����M6��ߊ-Z�7�ꊡԡ�-�v�jse䥳c�@�h��3�`t��ѹD�h@"�R�e\9���;o]k&���.��m��9��E �vRqI����)D:��B+UcV�t��H��rTw�t��]��kއ+�D�;�Թ����i��wQ��=+V�r,`�<W��n.�Cs�]".9P�5�`����V;09����O
v)5�IwV���X�YZ'.4&�Q�d�n���ʣ�%v�®;RU�Ei�-��t'Ġ充2�n@F���Kn!��U�q���(�Ծ=H�*����R���CF��`��{�#��������DћW�l��|潩9Û��x���67��7��:bc�2xE�p������aƎ;�r���ѽ�W=]=�Q���E�Wnn��8H
.������g�uܵB�_"4N��6�'0��ܖt;m�]��нx/QZg:mRݳ�����T��ݻ�����ݛ��]BQ7"��L/wf̻[�}�����sG�Rw4�f����(͓U�l^�XYW]����vP�=�%*�R���0.��q��-�������[Һ�HC�Od7OAqV]��WQ��d\��vd���s�ʌJ�=uʰ%r�4�ۙ�F��@�5� ~ ����u�]2�I�R�ۻ���n�nW+��g+��n\�˱r���.�W;��5�N�����tk���6 ��w]ݝ��Ers�л����&��n��iݱ�u�3].��ûk�\���.n����uڈ5�sv]�:�H�.%s��B��Nv���ut�wu�N&���.T��ҹԘ���qwc���D�s�5�H�;��������������˷"��q���ɻ�fr�\�!%ܜ1�:�Lwu�칸�n����v.�ۧuِQ.nDK);��\3��M˦G;.p����JHܸf�"a�gw�u΅q7wwuww:�r�wH���8E�fHg9;�1��܉'t�S�q�r.]wp�
C�D'8���:8i�wt	ˍ�t���}�!14�^�+9d�gt=ʼ�ǟ7�k�$��f�Wa��6�6�`ߜ4��8�D���֔.t���qb����zzw@��a��Xx��/㪗ǵ�+���2�
u����td;< �_w	v�F}���w���
<�ڱt=��.&:���+yn�����(��I7���۞k���;���D�&�e��˱q�l�B8i�C���j߆]8��� X�X�	o��Y<�ͬ��+w��0���N+Ggڝ�K+�PWX�@(�
��8nh���RT�ce�����=���΍?�/]��p��];�#"\�<����ޣ��:n�3�^i��\����H�UsXD���	�W���I���uM���ك����"���n��R��}JU���%��?X���
�Ƣ6� �q�U����OS�#��ݔ��w-�z3�u���_�[�}Sm���N�'��4kн5��9�H|��_^����vK]��D`TҸh��T��d��	��<	:��G]m.5�KTx�[��P�:5��\R�4dP���9Ie��?!�:�&�V�Ǡ �A(	<̎C�1H�T������h��^ss槰�׊�q���VV����V-�F�wS��@�k�"1�Q��+Mk����6����X�8&c��SA
�+r�wP��Xiӎ�����qʴ�Gl����5(�pS�i�02+2*2�o]E�.Vv���K�n����x`���v��r4�8��_9�!0���QE�u#���Ǿ��g��z}$��E��w`)�\���ڿ�����7]��=w�ĳ��}�r��òVo�n@������-&�/s���*����F��0rj�N]"bٌ�1�e��Ɯ��w��0�����
��~�ŝD%��͸�����xzpU{��Ȃ�.m.>���ז΋Ԑ4���
�3�o�N.&��O�v)i�5����=�����i��t�`ہ3��A���L���̈́��3Uq�0�YC��6��i�ya۰w�y+c���W��ey�{�T5�ݣ�~d��%���n���zg��j��u���Ӳw{'��&�@�K6Ru�����١��j�ddjt8����{����w�+�w��9�g����$�O�?)�0�Ʌ�,��@
�u\.u�뙋�43Jw�_Ok~�ԟ�Y{Fۮ8c�C�|�5�������s��uJ*�$�O�&�@u���
�B���(�Y#(�,�:��+�꾮��3����וw���c��{�7�yoQ�`�@�Ra�+�=�E>��F�q��@���]�����kfve��%�wl<�@9��8G.�>�7Q�m3R��n�iD�X܂�bɢR���2��>6�U�_�nz�滧�PL�Q�Tω�	�8V��O��j��n#f\ں+ں�1��}�m32l�e2��|�"��k��XjM��Ԓ`=D���������_���X��J�v���4�`��`2�[<����V��0�|�:��=~�������%����z�'n��D��%t��5ƕ�Y�~����Ϝ�Gi�p�g�#��z������M��"M��@�$?��>7��[�|(t�c��SF3��#\C��p�C���y'�{TmS�{�8'�@�5��a@	N���2��ák늸��8[���J6��N07+�;T�OH�\F�Dk�~	�rG��@i|<>'��7�Ը�߄��j!o
��<�h�{�>�q�%�L�����s�;X�s��$OCtZ� PC�`�C�0y���w"���gW_9��^m2��to��8C�q����HB31��m`�Ã�H�c$�ռΕN��P��+L\k��S�|_��vd�s�	�S�>�����i��U�yG}��=����b.:�R��� ��n��z��\1ܭg��-���N���
e�("z����.��¡�pE���&��e5Ywk:s�R�ٶM���{�:��n�����*�c%j́NY���5��b��9�'���`����1�l���ӈ|jފ�%�o��!��-l뿐����_�2�7,j#���z�hrv�T&#�����0��դ���R_�wO���҄>��cE�2�X�����N�2��s퍷6����S������bB(��x��{��b�j/ph��R�M<��*c2��t����l�pfFq-u}�o��u|��t+�"�:X8b��4?a�էu�� ���2����
]�.p�=�W�)�K��Zj��s|e
vk�GZ\1��{���������z�J�YBC���嚗����»�e���M�'�^l'z�h�t��n��Sh�5 ��iz������Gf�O�躙��Ӡ���Z]|������m���W\r��#��76����Rk�>�@W�6T~M)$~��2�}�џ>e��!n:F��=����5Ρm��L%��-<I�+�#��7�I���%��Og��T���w�(B�<�]�h�fx��;{�#T��&J���,r�
cGq���B�r�K+a�dQSx�l�]F��(̜W���)p`\5���7�ZT�vF�`t�E��T��hsv�������IM����t�od܈���I9�"�����/���;<�v�S�������
u�+��4+Ŵ�x ��O�
q%��_o0�:�gm�����H�C��;N7$GT<w#/�4��)@�U(�c��A�_��& zp��/�a7���6c���ò%;l�D{)��0E6�'-�3!QϕO��˷�_˫�ܝ�L~L���/�0�*��
Xv_���[2�\@#)���F��	~o<�5�>��"P3��M����ڭ���9���=��M*d��e���I[����R�e�W\�:�Y`S�[����C��P�G�V.��?j���Kj]5<��~���6ѩ��,�kY��3 X�i�0�gj�;?O<�D7�s���o�!ի#�}Reh�nom�Ќ���;'1�Z*z�޷�}����!�]ѻx;	��]u�C<%���^_T�T��{�ݼ���8ڹ�'�峝N��*a዆�V������b��F�Le|a�T���w����Y�&��<���>uSiQ�d1���1�G{����:�aF�T��S������w\-�L�`��Ŋ���T���fFRM�n���6s_f
�t�}hѥ�X}��eNˇ`��>��xͤ�R��V)�Adlo.�^��癲P�s��0�x3X����������.�f¶Q��hP��44�˙F�}�ӗ��ϑ��NXgd�t��>-�O�7/�ܕ.�D��}�S��tץ�͎�D)�f%��g�����*'Es����]ƨ}QR$_Jw`잤i�6�����)Ĵp�+/��C�'Iʃ*�����Q���U
�Z$F�tnΊַh��T�MT��/��Yc�l��T���h�l���'j"e!�T���+�B���Vo�	��Q:�6�������t��%�������p��M���l]T���x	���L;��� '�;o�ӡ2��ˀ���b��qۯ���x`�k]�v#��*�8���!
$�vr; ��\���l������n��jq|芅��hϥ�\3zX�n�����x�;�_o_ZJ�5ĞPfO�e�BF�Fr���*�۟u�����+C>r��
'�̣��1�
Ę#	q�ց<WF1����Dĭ�F�]�^N��zpu�ڞy#S.��\�+�&eN�0ҭGs8. h��7ȧ�w��ʏk��:͏uot4�ݙ�|&w�Ӆ���Wv��U_�Q������uPՒWګ��G�_U���aYY�����^�A���-��J�-l5���Z���P�:#<��6�5k����Z�G��	Ojx�xIZ;�yC]�jz�J:uu���lO�������0#�sh)�ebW׀�.�Ih���*Z�!�E�V�whʒݝL޹��S��ѹvi/%�Q�(쨫�~q)��y��-5���gܝ�1���O%���n����p��`���Fs	��N����֊�މ�aF;
��V��(;١��j�djr4�(}_�V(1��,��Qڲ����`R�(�Q;�ga�L= !��� F�bs��7\�L�P�m�/u��Π*�_1��_(�6�i�����P�/�+U����� 7��ȩ���w�{��U:R�pSϹ,��럎���I� �%����\k5^�;ڧ��F��k��W05��_7)���??�|�{EL~U�^D�O����BgBAf�������j:1�%m�?��	1_-u�.�,�e��岝:�x�i_T:(¸�wf�b)����+�K `��3�����=�(�폮Hf9���j���~�`��J���]�cX�=M
CGw�h	����O[�n����e4c5���VA�S�$3o��0���ܢ�v��_v�i@��i7�2���T-}qW�����A�J�W�������ȓzh{A�c�h��t$�+�NwZ8<�5���`d )��4�5�K���.��N��<�Ŏ)�̒���V:P��>���6��yΥ�+�R;�."oF�P�G�R��0�fv5�1϶m�0��11l�FG0nfL/9��7fڇT���d�� F2�h65t>�섮O��z�n��l6��A}KeqD؄�96��|6 �%q��R��`L��O��=�co���l�q���ts[7��2�9��7�s!�s8�x�h��"������G[}V�۪5ہ�K��"��z{L_���ާR�Ƥ�|�vd���F��
�,>���	�®�{�>�Xk�l�:�TWI:��ʠ����/�1|���/�N�E��s-�#M�Y��{Q�I��K�
�ީ��/���b�K�~��9��}��lh�����5T����f386�e1$��m�uE���n}��t�����;���1W:Q{�ne�|^O�O#�)�I���NuLɝ�L���7_.7���_W0E�`ٌ���Nu�Zn���B髞����z�Փ�Ù��������'~����^�BU��o�p�U�,�Vl��������ݷ\�fQ��\L�kh>�ٔ��5EBR�`�:l��\c7��A]���΢�Z!gn��w/�ѵR5���]��᷇��&Kpۡ�v�Y���k����!�mѬ���M�!�1r�]�&�JQm��vފ�{��8�z�uK����|B��8���Vkʉ��q��)�]&TI��s-�׻�n��ĩA�������UL���tcKկ���<�����*HE�ܶy��|o�X�'4�\-�ٛPч��T�0l���?��&C���q˱S>���Fz^G�3]�r���+�w@qdIO���i�����.y���k����oe�/�Og��ۘ���"���j����¤G�m����Ɔ�_v�,�� z'RP�1����P����I�[���9��|�*�X�7
f�9����r1�ⶹ E/�>D3�{+L�k���������0W�\2�������␲�0Cnbo~uLȥ2QC;睐������x�+[J&�����&J�Ρ��Xj��W>�Ϝ�e��+����s�N�&�m��8i�&�/}�r>��{�)��#�ȿ�����[]zu���}S�JY,�1QTWY����z���xl�n�����,;��+�tΘc+2�Q����Ϋ�U�'���6�B�fk$�,¾nX^#�bǈ�����!��o��jC�y�C:���r����u,B��gXX+��"�0x����ƨ@⾱�x��Q|�V�'�����k$�O��p�n��Y�����^���[��s�;P]5�&�v�]v���w�1]��S���[`C�]vf�H�c�1WK4,�-iY�@S"��	-gue�<7JOn��Om߈uq���ݼ��T+���g�j��y�]��\�ݏ���<L�ηaٍ��V����F�f�"��zQ1��TÍ�Mr��U<�k
xe�NQ��N�N^u +q���P�(���m�ꟹAJ��r���5��s�4z�4��.�EW���t�<7��/ /�s2:�w��6yuL
����Bb�ף���/�K�\�ʹ������\�?������[:��H�6â�Gk�Ϊ^�p�&guNWJ�V��M��]�$�h��\�#^�~B�X�7�=9;�����ᙛ)h�X\���pً���ȉ�����N��(	���Q�	i�B�浰�=
1I����'#R��!�,�9~Ci�\!d�*��x� ��eP��u���E��p�3aKG�UX�D;u��l��pֻH���F�y,}�ĺ��v4f
ȝ2Q���~�A�.ۯ��b8��E�jv���ڿ���Ʒ;���>�B1����Â����T)s$���z��N]�o:�]�\NPַ��ol��nbz�yj�yӛSh�Ú��Ɯ�2Jm�M�
���8�[9�����}"�,�핼��n�#'A\ �]������Nɋh(RӜ��_7[N��e��QV<Qأ�ֳ�Mc��U�'o-q�3 B]��N�۶^��Bk�5�$of�Hv�&rbϜ�L�e��
�!�]vU����7�®��r������D��h_-�)�aEIKː.�I3�v^!�Vk��ej��w6TM�[َ�<����r����d���f�iU�ڑ\��%ث�W+�K���4�H7�5yu�s���墡n>��ֵ���rw:���'��G�|�y�\}�צI��a�A��Nj�.بDf��/s����B��}�~�)���(޼%N'�蟆�{z�L2��2�kP`��X%�k�+q-�J�I��kZ���F�r�^���qW:ĭ�/fc��Zʼ��uk�	�f��NH��Lb~��Ս��I5�t/��nw�e�|T)oF�+l�-k�V�t����ݔ�s����Y�wь+�h��0!@������Vv����ө����R��H�X���6���ː�9]����a����]����}J�\�D�WH��L��ӭ=*2��r��9��'h�P[��=�p4��`���s+�)��1�YV���7s�Q#��L�utu�P�{��R�����WVV��Nl0�,����F԰+�M^���-�.w]0`��9c
9}4�]`����U��9p�T%��GD���重>��ᦁ�Ќ�����������z)�K�#���]B�<�mP�t�� �ސ]��겫8�n�n96wM�_w���|�6���\�3ru+���p�,���d�u��%�:jY{r�ǃ����V�v[T��]0��(�?�4m��dV,r�ݠ�Bz�s�z���D���b�ueIl��YQ��P��΂��,�5�Cu�.�,�q�h�+�Z�x�>�A;d�]��fT��q���+��!V�@@��U��R��m�'&����tt-Uk	�`30� �b]"����k505K7��w��b��7E�<�t��ţq�^�@��[���>De��y=�>�"�찒��Gx�	�Gv����z�Q�I�R�g�|y���͈�y:k��9=���
F.�m#}v87���%���|H�n�dP-�]�����\4�u�9B�GH�s w+�B�퉳�� M4�n*�ǃ̓[�=�48��l]��qק`i=뮢��t+$�po,�і�-��ʷ]�+u�@���T�h�9C(�5.�Q��="�vo�����i�;c�.+�%�W0<����)�6���L�7�S��m�8:��i���;��1]�X����#�ul��s�tZ�i�t��Lv��;�:����ml9|.�ݎ�
C��
�>�\�4�s���]s�F�'8�L��\� �t�r7w%&���ۍ�u�t)���M�ݔ��D�LW8�`�]۬��9�de˄r�P��);�H'u�۝�!˜��p��]��']wW9�u�ܛ����;�wK����S����w`�rqw7u��s.p
wb�F"%ː����.Fswu�FFΡ2d��;�k��ewwN�bB��%�9�s��9�;�J9��D&N��s1wvcI�c���"�g.&\wK�W;1]ۤ�nt�E�9��\�1HAI%΂	I��\1�7!�Ir�`�� sq݃7u��q!��Fnvl� �wL�.݋�.�������t��r����Q�s�I������wb�C�;��F����LҚ%�$�"�4.]�w@���n�tk�]�N��������qwt)��%�9p�4c#7wݺ;�pK3%ˍ��H����� Gu�w$�hB� U E�Iyh�����t&�K�9p�k �o��Pp"c(�}+�7%�^vG��@�3���(Ds�2:��GN�Zt� �cfQ�g7F��hޚ�^õ��^-�Er�����������^������ţ��ｷ�x�������}�~�E�c�s��|DDh�"��}�t}�t����//+��pJ�����x-����[��~��y��߾�{o��ݿ+�W��~-���i�[��7�^����>ux�y��o^u�o[��/ֽ��{^-������Ƽ_��o��h>����+�ܫ2O�o%J&e�Dh���������6�������ͻ��V���o��������Qo�r��|�����^7�7��<xѤ�ۖ�����^F����~�j�-����!fJwtI�|��/��5~k�G� ��+��k�����~���o��o�{Z�s��|�B�O���
���Q~����k����_|�����mx~v�/�_��i�m��/w��m�C���{7"buL�[w�7��+���>�ۖ��﷯������_�V�o���U߇펩��>b>�#�����@1�l'��|W�G������W��o���Ͻ���?��������_���}�����4�	�����{�hs�"6�ޯ���+�����~w^��6�_���������r������o��/~��(t a��v�H8G���>��}U��=�h���������������cQ}(�}��<t����3����z�P��n�ֹ�u���{^��/����}^5��W��W���������^->u��KW�o�y��s�w����v���ssn�߿�����O�y�ׯ񏘈��9��J�>�&v1ǹ� {^*�|xѾ������r�����~���潍F����~/j��~u�5���+��_�������o��7�_[�-�$��&� PR��#� (
=�$DCG�G�Dg6��,;6������6�[�r�޿|���m��[���^b��~�_���[�oj��K����7��m�~��^�{oM������<[�]����zo��7/�zZ7����{k�� ��6��1�Qڜ�;�f�{&Ө���W���o������77��}�o[x�m��o���Ͻo���>�������ϾW�Z��o�����͹���W������6����|W���^ּ�[�G�A���墼�#�}�<�R�(�X'�ɽ�t�����q>f�7��N���\$K�VnV���զ�Q��&�9t8�圤:c�{Xﯤ���0�}���{Yl�1� � ���1��-7��(LCv��k�l@"����ۢ�����i���$�����ST��b����������_���n��ϫ�������o}�������[{Z-������m��yھ�����տ��{W��|k���￞_U��W�s�l ��0x� D(��P |>�2�{?o�8Ծ�����������>�^G��~*���y׍�?V�m��ߛo�~�_�U�������o�����_�[����B}�+�����k�,kr5�<��J�!�}Q���$
�r���z�޷��o���^���W��s^��/��o�\����^�Ϳ��X�W T�Iq�Κz>���������|���@��t|�|��Y���ҟ��}�<0@���
��G�����wίm�{Z7��u~/Mx����EDW��޼�KO���z�{~��x����|�~?�����o���k������#F�Xۑ:tfzk��J�]�ݾ�ۚ�z�~/k�o������+�ͼ^~}��k��+���������\ޛ����zU����w[���nZ+�ϝ^���y�����3��"<#��=�Ү�w/3==l���zk��~���\�kE{��}[��_�o��כ����>����_}z��{o�n�Ͽ|���o�sr������-����1L}�ƾ�T�#V>�����C�i����#�ǖ<{׽��
�ޡ��b�G���1�Z�d����ӥ��龫�x��߿ޫ��F�+�����}oj����o�r����^U��������|��{U���^/���-��!�Pc������������弞
����KO���|^��*���&߭���_�����7����ͽ-�^-������s}[������ޗ�Gߝ|k��׏J�_>��TE��ߞy��?ݾ�%$�a�]�
iE;H�H���/���x�<���?��hߪ7u��ŧ�<�[z�7���������G���>b �}meF� ���#�}���#�c���D��0>���*�d��Kay�H�D��}�&>�"=���>ܴ}k��W��ۼ��~��7��^/�����|_�~w�/�~�Ţ�}[����x�����|�叫�������T��c��_\}����>����7t����y�T/ ֳ���a��P|�X�/z���n|�ٸܩ�ĸp��o{$}�l��xU��5�KY�ѩsY�|��vEJ��3N.��gm��׳\䌕�*@�[�Rr,fRf17+�����2�bY�M�'d	�8fÝ��S��j�3�H��@���DX�>�������}��*�����W��nW�����^���{����^+�׻��ε��������~�kF��������t ��T��"> d o��q�|j��3��M��*��U���
�\�o�_W5�y�}�x����������"s�G�",G�$��g��>���G�_�~/So������vߍ���� �}��)�	�>>���\ttbi-�s�=��� ����D��=74>c�kƼ}W��~��Cb+�����_E:��|Ǆ}#��D��������o�z�+��_�������+�_��,����>�ژ���#�H�R|\��3dו�Oo��h���z 1��0	��[�޻������ֹ��/���m���+�~��ޛ�n�����c}m¯}�`}̀��|QM *>p|����@�D}p2�_\�: P>f�z%���XUװ8���{G�#�$}"$}�~�~ur���{�v�*������=v�m��U�K��}�j7������k�|y������ߍ�W��}��F�͹����}^�����[ž���~������~����=����2�{�}B�몗_��u~+�x�^���W��������r�o�1i��^y����گ��������~�{�ڼZݷ������� ��ӟ�p.>���En�V��Y�=wǽ��"���"6�1�X���E��+��o���Qo�������_�k���ݯǦ�o��o{�����x���h6"/��^->v���7��}!�p�*0G������=��A�N���i�>��DP�� #��}��h���ޯ<��o�5��}����/��^?/��_ͽ��\�o����5��ux�����j��ޛ�wv�_���W7���#	�(|�|@��gH=I�{n��s�xK���aG�}�5#�c쁱�P_�V����~^�}��_��W��/����n5��?�߾�z�?������ߊ�.o�~_z�{��z^��^��n�>"G��  ��z����N��S�~|���ׯ>����6������F���祿���p��Qo���W���������7�����_U�x����������_�>�W���~��^֞�� XdT
�|�0OS�7ڍiu[b��v������!�ߡ��J{)�y�X�ǅ�-w1��Y�q[�,^J�u��2�[.�4���a��R�Xp�+��q�����@�i<@�lL�V^^�3��O�]�{�Bؔ��ՙ]4'#��/ɺ�&оTZ|򌆂t��T�%o﫯���������{W���_�żW*��u�����zom��{��o����s~��L� Y��	�~Q�쏨}����Z�����Ƕ�o�ƾ��k���#��Ǟ�B�.���_V�1�����b~�z_�i���W��^����˻z^����k�w^����x�{���n������m�ο�x7��uzU�r�����ܷ�q��ͽ/CPD,�jME�U����*&@p�C>�DJ��<�zo��ݷ���w-�w_������n�����<��U�y�s|_�y�}[�zZ7������k�_�����5�o�s��k�����i�<^��'W�/'�R�Rcc� �c������oM�[��|�nm�;�_~��o��Ϳ^}����5��m�ە������F�z��z[��x���x5��A@���M��1��LL�@Q���Y����[��g�Ӟ�����|�D�L} �4D����DE��1�|���~?�x��~�����5���o���^����v����_�~+������~���7�o�8����r�yߍ�-�]����5����٭��k��n����#�!
���>�E���#�$}>B$F�1^��_W�~_���_U��~y�ר��!|��=�u@����|EA�����I���|�zZ�w�����C��K(��Τn5��D�wFDK�G�����} lOO#�f�{�EۂهyR���&>(TU�a�,B�V�!�N���\d���8n�N���n�ۦ���^����K����W�bx�m�,�T>&��y�Ss�ٯZIY"����¥����J�����x��i�����h�u�#+�-%���^���VC�G+��n�5FhƥԚ������Cy�/	w���:5��iA2�ޛ�"МZ�=����NJ<� 5������:(�߈]�*�S�VLs��g����xhm-���C�vR�:����'��d�.��nS�ղTVz7)N��ʱ��;�\�(h�\F;��\�LnGӕ��&'�����l��N�5���qu*�5�S:cE��i(MF�o�D���?!�:��&�W �<z2દ{-�n��L��pJ0�3y��*�g!ۯ���x`���Gc��*�2X��W�k��ۻ|���Q=*��I�N��ZH���N�S�)k�j�LޟZs������&Z��M�G��`;���h�(�8�nq��U�'�֦�aɦ��j%EL��q��Ɇ"�%�8���jc��A�`�{F1 \=]��t�\V�p�+�o�G4*2��rk�m��`��s|�E���w����0��X�Y�9��uT�F�r�a#�o\�7�'���j��y�'�t<�j�q�$�vw#V�*��[)�(�������QR��p����ʈj�z�s��Q����mx��u{ܸm�8���S~��a=��ܕ%+������@y|-T�`�k�p:qV���f�.�����
��L2�K�]i�k<[X�z��G -d
h�R<�w'2�%�v����K�Pϻ�Y��W������Q�q:(w�l�<��M:ݾ*1Y+`Z���gs�mw����=ᢁ����S�녥��B�A��\��PƵ>98�]���bb�~��<o���p�lA��9��L=5�(`9q�h[����t1gST�����g'Q��U���s�j�TMn�O����/�+X���=9�G��J�vr]�8��;"�T�D�)��g�����y�Hx�/�,�u �ݦש|�U�9�
��W1��ˀ�e����_o�����3m�p�ٹ8.-I&27uG),�+W��'����=��m��L_[�&*��hr��0x[-�N���V��l��M�`,ԛm\�κ2 �P0W�J9�.��)������:C2�GY����,��s��m��S}Ef��<��&2��2�vc��s��n������3:C�YٌK�ց6fkx��)z�s*al������P$�ZM����*�����r!��\�=Aݙ���KW[���u�C�z`�ߝR�*s��|�n8��Y��C��M����O؍C��rt�d؆����6�ݿ��]Uā�,���Z8�.g��#��S|;}���Y���RW$���Е�:�I+�b�s�=+��<8.�V��f֛=�#t�e�M�e�b��O����5�q����!J8�mⳛ̣��`��o]�6_P_#�4��6�G�� Ƙ1���-K����C���]]����<R828�\�c9�:<��.�2^qz��_�H����ÿ%�6��=z�ST0��W,c��U�����.�q�Hv_��Iْ�����3���;s�����m�uya# ߘ`=��-��[�G�o���~YR�{�K_9�f�(���_*_�eI��b��VE��o� ej�1�U���?5�m�½2K���Ko�;�ON����L����3+E�����]WR"�0�r��̍م�VSDOv+.��m�8�-Of�8ں���F�m[��Ҿ�ume讹�.�e�*	Vlcxj���1��d��q{Ů�>o�G�J=31|��䩤�'b�b=&��tX��F���w$�g�
���%*+]gOz�,�%��%�e��5.���1	�S���\c7�9̣R�;�^d����5��x�PT��-�+J�L���"�9���_ �9B0M�Kr��g�-H2$��m�+��7�\�;f�����UL��?IQ˱P�`b����v��Cy��>�֣BΕ~�pe���������{Wf���k�ٳ��Ǯ6�A���6&)�s�9[>u�'���ϊ���tz��{ɺg��B�X;��ov�c�J�ҁ0��c�5��)�F-q���{�}M�!����J�^���������e���Z�|�86(�=�IUc���l�Er]SN��=�ݧ�&��?QN��jK1���Zm�T��U�h������.� �n�������)�8��ү�ucxⶮ*�e��Ɇ;d��j�[�4�ҙF��=����W=�Z�!~�̄�_��5w�
�2�gup��S��`7��Ȃ�0T6�'')5F�w�&Lɐ�'R�e}Q#���2��'�M��P��Rø/��Q��C�e������V����$'�O�Ӫ��\��PJ���#�ȷk��oR���y�Kv�J�m�]�*3����d���`sϨ��%:�"c�'j���yQQ+�t�l�B(��5��4TZ�ݣ%B�#���6�\��  �`ahd�P���z��~ZF}�����_n�|���D=�=�T�Z+s*:�'w�S����?eBYv4,��5 �8i=�&YL%������7�_���[q�]�h��{�����������Y��[��vx,���t����*� �!��62��q@�y.v}i�J�I	�˼)�s2�s���QY�r����/��pl*dI�$*��]t��B(���a�����y���Dk+]%گ=Ob�O�[me��Êw.YtW���D=�r@^Iug�����V�N\L
Q@���1��ÁI�?d	����:���C.���.q����[��[�ש�Dek7;�Q���8�\*�E@�_���)2�ar���R�>�9�e��J��+P�6�R���O�fD���硫�L�0�x	8��$�¯�ƾ�TN5���6��W��+qF���O"E��N��LG_Ϋ��ak�[���� `TF�*��[Pl=�����ԡ�4��َ�x�-wp�����a�:��)j�ܜ����'N�bWK�B7�f��r��z�ꍺ�F�0QA	�R��!�,�9���םP�|M��|���.Z�v�҅A�QW@��  ��`t�3�������ۯ���x`�k]�v#��*����n�~�"͜E�?r�Q�h��Q����-$Y��t)�]pё-��9�k$Ҥ�n����$��ӺK���P�����+�E�Ai4��ۊ8=�
��Sy5�;�����\�ʃ3Hqo�����&.������q"1� ���;$���^6X0��W|_j�d�<o�΍���
V�w/kyU|��j�9�!镕6Acg�X2����G=�&vj�ح�Z��ZVrd$\�Ne[ �}Wcw�����w��ڙ;�-?7�Lk�����*Esc}�I����"�z*gR2�}�W�U��Ԝ��''������|�FZUMCn���0�c S*L�J'�&q�����gc�=�Ǳ{���P�-�Ѭш���7�_�	�"�O2d�ͺ�3T5��o��h��NR�+=Z��PY.������a��_YQ�S�Ts۬F3�%YP'/�4m>qdV��T�ޞqE`�֋Gt� ߅�>�1�TxpTW*�ct��ȰÆ��B�v�N��٨��H��ξ_c�.�N��f0~� �hװ :�澻�)l�@��}�*jL�`�*sL�뙋�sC0L���Mo�<c�CܾTY����u&�k���}�BJ�]+�S�H����.�U�M��櫩�૩�pd8�k>��̄*H�}O-dC3��l�=u몑�W1ٗ\�%"�z����]CY��P^����~�O`�����ol�@1(��^������?,X-�^��l�N��˜�7	ٖ��%����Vϴ�z�:�=:��ʔn��Q��[��q�"��K�YSȍ(e����u5�M�\l���>!�AVf����[��=�j��w�;Ҵ��T���.�}�S���YZ)v���Ѹ-����j�>e��W�a�V4�詥����ndk����G��0�]�T��̗��C��s�}1�A�-�d�kt�bB`�3�zX(Mp^�yZz���ؽ�FH�}f'�Ӱ ��)���o�kYk�ɔy��h�7�y-�Q�.҉��J��X��Y4F�����n�ʓ(�v��
V&�IO:�L��:�tW9��;fm�F�TW[��m�F�fꝩR�CQ�o�<�9�^�9��/7E���n��H��������Gb��bcg[���o�c^��0uZW[O��b�-�	���o���M������Uҭ-��,P�d�P����2��g6\�h��PN��m�
��ṥ�b�����$ c{%C�h��vwYɸ��9�c�0��6R����V1i�uك+�ut"rgR�[�{c�S�ϔ�C2��[}����<%�=� �۱ �^k�7��kD�ң2��z�cP�eW<�Ǖ�Ӕ��K�سY2+4���� �k9�#2��Z�^��Ԇ�����ۺ>t�A�t���䛮� ���I�}/�Ѷ�]��j��ɨ̘�)�z.���ʅ��º־��r�֚qtU};K%	H�I���{)�4xReѱV�=+('��V�v�ȯ�T�X�����Z�R�V�Ue2q�[��ҾۥM�oC��ٕ
"-��[W�1�T���)��;&�B��W��ʰz��9ƠK� ojWS���q+*����M�x�-Mv�$�����7�1.;��>��*j�ԙ���T9y�,��i������$���L�d.�e��x��W�[:,}Ē�w�PJʷ�lܜ��XQ�&V�/�t�t�h.&�B��K�}�.C*^�T��kj���ER����ϰ�M����{�H	VA�kNu<�k2�Ш��"wMz!�'dvc9�=��[�r�>*�cR�erN	]j�;�ѫ���Y1VFr��߂ScZ)m�	�	��¬G%�m��JY�8��D-ƲP��AM�g�t� ����2�<ScXZ����^q�"��a���*�U�qSg��z�9��A�y��U����!�3(	y�v�ʥ:&�3�7h�8�R�P۾]�\�Q�Iv�æ}��sb��H2�n�;r�<���4����}��Vb�g��d�R�A�ڸU�آ�[Y������b�p��J�;N�d,���ˢyvo�}�;��_	mh4n$��}��VCaR
�ˬ���T��)��\vmD�W�������B
�&
(�[�����@]q��PS0���PZXwQ�Da�n�eJ��v�.�����N���;�Q���nCt�ެԞ���f`��Vtsfq�Tֲ��)]���I��|��޿<�~�m����ݤ�	�Wv���MӇw�((D��vM۫���,���fh�0̱+�\�at�K"��k��9ȗw�L���Hh��@�����n�d�4f�tӛ��!.��	��븡	(.����be;�1�JfI�L�IhҤ�a%,���;��e�D�2M"U��Q�
.�̜䍄#!L�K&IH �7.BY�Nr��nt�I�%l� �]��F1�`$�$�$��wCB��B�4b$�2��s�B���$��,#�CL�)D�&s�e���仸���ӵл���lú�`��I��5�t�Qc��22Y)J	+��eG5;����3%0Iˤ���`��7.A�;���(hܻ ;�h�]�6�r't�,��뻮pW7##	$�!��2U�]���U����J-*��ݣZ��L��R��o	��E�R"�0D����뛗*Ʀ���nQ�z����B�a:��\���S���ꪪ'a;=�U�C
��S����1P*�|I������R�zz��0�X�gWm^,��9[Tj���v�q��a�1�ᨅJ�\������`�ZM���/��kj爨Y�>����e!����(�Qþst��s�IOf�2��*k��}/j.H���vy���{3�*�oÞ�D��io
��:H��g6s�/k���؃�d��Un�;�&T
cOG_���]J�·�M D�
j/C�tE���c+�[�Cs!�s8�hN�D�lGtLt��;a�=X���|�_�Q���6�W���B��1�VNd&_��Iٓ6K��\�Y2�	�q22(�B�^`�>��5\?e_��G�T�&x�t����~�{^��Y��b�F%y�3�!��GL�r�&�����^T�[,��*��~k�0�8�W��=��nZ�&���Z�Kq�y��Y,[uLE���fVC��t�bFGUԈ��(����������)a��&�/;ݼh`�,<S��F�cI����U0sb?=��.��`����/D56:�[�k4��Z�Nj]ǳzѬP��o$�l��DǢ���f�]N.@��S��u���s�\$��`7������������j�qκ�7��n$9�������-����T\�����t9�C�()��:�N˥2�0tB��� �DDG�G�k�mԸ��S��O�ʭ6jy����ϮDJ�L�dE���}����RW����]�A%u�_�k����&�������e��+R���#R��\�z�9̡c.j�����X�6��Ӏ�
�R2�]���#eHEv�V�?�si�ӷ���K-e'0ȹB%-ϝ����iq߬�����\/攆�g�}�K����u4�>ŶfflG`ެ	�2��m��鹹����(��� >0�ک����&�4��ɝ.�Ӫ�x��Og��<9If6� ��ީu\���d��X�:�赧�v�(M4Qg8�_���V7�+j�e��9�c��ruC�r2��3�Z)�B�����WH"6 ��$�-��e��q���òS��g���D3"�CӼju��Ȝ��*&�Ϋ�^H������BFz&/�9׆����?es�a
��7n�'y;8�Q*&Gn>�Fi=u���\��u
�v���#�Ⱥ�k��l|=��:L_�g˧`S������U8���u5�ي��y`v5\��m�xob0e�F�x�%λ
���6�y��,�X:�%[�J�y"�At�"Q�m)�������˽G�s(<�����NzA�/1j��?�UU}��'���кq36G]3���2^3,yDF?w�J��u�(v��U��<{�c_�J�Y��oa�2�}��jyL'�R^ B�����X�Ë'�|��}Bb�?�]��G��8��9�v��#��lV�͍��F�!�����g19���̳T�x�~�1J�{Wt��|��~�E��֮�4J�=�ꦿ?�va����w{<�����̔�l󀖂"l��Ńf�D�Ad�
�(�Bx�r�Τ�W(�N�79�vd�s��8	H�}V7���1q���Ѡ.�\�C�Ӵ����\�c���n�U�Zn�f{����q/xl���0>�[o���t6<s�f��
���6�i��T�S뵮7��°=Uű��\S�M���u��1�7_Lv�H�(��d�+��x�����K�9�a��z��
�6�U��wTa��a�:��҆����93,gBNbi��,� I�Pc����Y�/�`�H�Bj5+|q�,���\v��ճzg{��ʬܾ�I�+��*��O']�����4�V!U�7`:�d��\�v�$6>6��za��+E�:F+v�I����u{���@�k�{'�@��ǽ�3l�&qal�0H������i����Y��׳x�L�b; �9"V�C>���磌��N^���V�e"�`���	@Gfr�G�UX�C�_M|[<0\5��0wl�(��ę���'F���H���G?�IF����Pd�-$T�jv���miYg�u]ѫ�n;�S���l����CG����+�E��IO8ͷ���uU�3ڀD������w�}@`�� �r�E�N�n�n�t�f_�A`������k֦����>�.VuNw�_:�����J�ɦ�p/<_�_�k U��*'���k��kmx�Ұ�X#�&}ia�?nS�Z:����}Zj���<ɓm��3T*����b�K��q�Ϣ]"�6c��rtE@�w�������r��`_Vs��oy�7��O��� E�_.�w��T�PO�/l�{
���|-WK
�s5�8�����١��9��쉅��Z
5��θ.t8���_�w�ūʜ7��ޟX�W4k��u�{:��Ow�,�q��RC':@��b�\�2��1�ȼ3���&״����/���q��<�'TweS�:��c�0+z�ԤGm�	LwWP�+�K�SiW7�>b�t�\2��o�71�����A�(�?F�l0i��'��*���ՏP�L�Y-���;�]xq6ߘ��G��8l��❝v��glʹ:���*	`��D},ygZ�⣺4{�3�Jϑ *��ȺQWq#�9�jw8*�{���KG�vka"����&W�V=�˨˭�f��!�����Y)������3o�Q��.Y��Q9ۖ*n�"�u<�GG�ȓ@p��������b���^�Ls��ۖ�7u� 4��/����|���Vw��W�GDj)�]� |+�J9�3�>T�{޶>V�jf3\U,�s��DQ����S��j��A�g�#��Y'�@_��*���Q�ح�*4�S�Wx����q*P�p�SF3�r0��9�B�P�\�h}��0�IJ���Ɋ��մ��ݷ�qR"���_p���*廎Ծ9��M�ق6�uHM)�����TN�L,aO�s�3��v��\�����̫���D-�_Trt��3�8^�۬���Bʅ5��u��J���Ykx�@Wq��E���w����?���6��b���%��rI)m��]�)�!�4 �m�)A0Ս�*a�h��ޕ�S�|_��:��c&�޺yZ;�����a���RL��eX���.Ǫ��ص<�f��]�d��'/��t˚*t�VJ���ۢ��zW��{�ʓ[���C�d�B��yRiTs��L��Z�N``\�P����Z��7�r�u3tt�O�Ld��R�d�������}�CSN���d�7�#W����^���T1}��Y�K��S����ل6gOS�����WOyE�3�ppӻ��s4ܰ	������9<�9Q�׉���n޵7�C�[d�󍫩x�;cE���b᪦"��̬�Q`�lČ���Q��,s8�v�ێ$h���NV���s(��Ζ���j��C�Z��U0q~{�-\��d穃���H{8��a�NY��N93�~5-�l�D�|��䩤�&DZ;�&���S��N��
�Bۛm���ޑ�e�D8��6l�`B_i-�3�՟l�h�b5)L�U�8���ME�����F�q��m�z�h�t�b�tW�𶗅=|����c��Bk�[qQ��T"����qU37�����Χ��f��.ʔo�0h�3{/�s�^��^IR�d�+���>Μ��8�z1�c�:������ƣ�$�3���ow�d=�mU�qs*�l�î]ĳb����vv��m���Z^���U_(OQ�v�T���]�i4�9�k�}���`�0�f�����J1C�1�p����"����z� ��}�V�l$bY�f����;0�K����;��ҟr��.r��Q��*Yҫv9�u4��0ϥ���KAt�w�kn���R����������7�-�r@
���:cDW�G2�X�8�����c�ۙ�;NBru<w#9^����v�S��L�J.�ޕ０"���.�Q)�F���Ƣ1up���N�x@W�:.����`I�s�+�W��x�?ua"|��L[�P��Rò����'"�����m�)u4�=�����/�Uϝ'
�v�	T��0ӤtyN�CN�	�;J������֣�V���GT�ҖKP̰9�`d'PDON���Zn ��`�|QâK��ڢf@9�.h�A��qqNa��چ#�A����`9�`ix�ՋË'�3�8��;gVb�X�xL��,Daē)^��������K�e�+��(�r�s���(�qVng\�,v|2~u7Le�R�-������P�^"�=X|�Mf�_���h�+j��*���0�QA��'��bM�u +q��6�GJ3yl�gLE�Y�Z�3�u�xXs�\��<�O�q�Uܖ+��{GZL��+�_���86��kL��6������:͓r���"TY!VT������6�X����T����X�Z���Z��Zr�a뾸�Ey{/H|E7G���Z�T��1Fn���7�'��\\'�]$�[�A�U�Z�^�.f[���C��\���ĵv*�U���+����I,r�7F�[fFE4��n�����t�y\.7���J\g�N�K���O��d�N;�qѭ�3��vB��՞�C��r����V�%���E��ۍ����^��{E�0/2{����0&�P8�TEM
�W�V��]�qt���<���6b�%�crr�q����uW�-�t;B�2L<>�'@�:���ׅԵG��<N�+|q�,�:>C7�\�D�ց����N�ĺ�f{�lR�<��N���NJxyx�v��6�4��Z¨_n��6fu.-�U�d��TC�B���(&�E |k��Ω�[�9h���uJ��E����zú33v,?�󿘭,cs�J�Q:\@�~�`#�@K>���?k�'�l���g��.������^��,o&��-�&/�b�&��Z��ufС�O~����S��NLMt��l�����ל��)�p�C�M��}�/�/�`
��E5j��j~����@��/�!�v)i�5���4�������UZ<ɒڐ5A�9�&����?��C�[37�b�0��،��Z9�;��;.B�d+^�S8�~�>��Ru��<W�S87=�ֳ�+����:�h�.�+�)ޞV�.�*����1A�'F��mq��.�T "r�F.��%6ɇ9�a��׹Ǵv�O������O�\9�@���,�1)��9.����7��G�ž�"�N79;�b�q��-_m(���$��qܶ�۪��l�C�+�4B�t��3^ÁӜ����\<�]�9�c���ZJF�u>��n�Y��Վ�X�yS���wn���
�a��-�JF�ެݛj��аq����C��g#�[�O|U��?mDѶ��������*]q���qvkm}�QT��L�G .tdk�=G�\�T�pU�c��/
}�9sO��K
ކb.�G2 �8���Pg��*�o�b:K���Yd��Je��[��W�� t�2V*\�������h��I�TO�0�����b�P������`��9����֡|k�:��z����eS
�1���:���\Q���q�ʘ9r�e+���ѝim7&����\!��u�uצ�?0�@��&?��!���F$&���3F:�6����W�Ĺc�YM��#[��p�*J��l�
��m���r29�� :��C��ڻ�N�&"ݺ��/xT.�����2�t�- ����=�6�e'=��i��Du�fJ�A����Y�Y��]憾a-�޷:����[
��o����{�rKFG�ˮۻȘHx�*��#��>���*T܃6�$�=~�:��-}qW���7O��t����:�%T�WLް�s�V�k%�.x ��|��փ��l����N�9�������`����R�>fc��jT�E�>��7E�6xAҴ���̸��W>�FṈ+Ô�|�%�.�=�G0��&z�q|H�44���S�C^�W�|f�{
��C��x���r�Y�XÇbfFɍ�Td�����h�dTl�2OOh��hp���h�a��:{k:�kj�"_��Q�E�q�p�i�Ȅ�s<ܰ	�s��w2Dl�z���� N��Z�������נځԸ��K�#��CDdܱ�U1��fVC��t�71B���EaD��zj��4�ٝ��R�wYI&0E��[������j�\n5]A��/���R����s�֠�@R�#��T��/�'w�p�MQ���^�+�d�Q�G�������[
q�b�|���t��j�|D�,��U� �/��Y�pz]xQ���R<-5��f�VB�D���3�CPd��2�|�V�g"(֎nU�J5�y���-g�A���+����&���W*Iw������t��l�c/EsneX�����lB�04����+��7[{�𤶗΄
��W#kV6j�hf�+2��hY �N�W�{�����e�B�������7�����.L@��!��\�a�5Ɲf�K��I��u�]JJK�v�j�ۊ�4�urFZ1an�;��`��J��z��g�.L���Ie3N���3��� ?f#_Z�J��Z�1+Tx>����W�����Jj�Cy�HhS�otG�|�5=��1jN��u��t~�Dxu��p?�@�M�X]��;u�݆�r���n^�¥��T�gmZ���=���p�2���Z���e��&�qT,U�T�) s��ǆκK�3�7�;6�����OJOn�[�y�%���&p���M�W&�0��;o���8�o]���]}ϟe�һ6�R��Ђֳ�B�H�^�@��p2�����R��Ur
n�lM򥛖8�]�JI7���<*�Y��m�]�q��[B��۶�� HO&���%o[Ra?
����&���Ɉ���[��׫ �����w���Ԭd�X[��ͪ\�P-c�.�S�w��{X�]���4��7|kW���V���u����,I��1�Q�fV��nT�����+��� ���*�0X�˨�JӰ*Q��k�ei�����Ħ��rՋ1��2�I���
���
��	������O;{�������|�`��m�`�t7ca�<���r��[V�#���=E���i�ݪk3Q�j���we��p􊜜N���0�3�ؐe��Zi�i�>�&&���[�2û�Z6��r\xZ��N���WJ�{��Mϻ��Zl>���a[�i���QAC]^�D��O1��g��% ��lP�����m��&�b�oy)`��j�vt1��N���ݏ�%b���j�t�$�e���\�a&pP��J�;�.��t\�S-,�J�Y��Su!׷�/���f�ȓ�xf*q.��b����HV/���v��qi�.ly��]�Ob�o�����W���I:��ԉ��{�$ﲎ+Jf�Aw)sy!�R]C9ʵ�/dy$s�k����hfZ��,�*�3KNs��`[0�K�����y���u�4���`�Xl�n���1�6��y���s%.�U#↵;��,��1���:p�i��l��z�t^e�t�⮁��|�G`�˘���������f���
Xlh=%2�u��s[q�QP�k�+�m��j�����ɕP��o.��E;�z�uIC)˔-�@m.Σ�{S��L���#�]Fr �R��.ּUܹ�n�t��Mu�]]��R���T=Q�u̔��cO]>�+:t�z�q�ț��ݸ&�4�2i����1�$#&���ؒ�8�F�7w
�]ܢ�$����L��H� �81"E;�"ܰ�h�	����)�I�)�bfPwvBH��ː�b1$P����� h#�c&��$�FP͑�cdP���bD��L� ������2%Bh����D�ic)&ED�K2H���N�A0���
Q&e*ha7v�4F��B3wk��$�6"�L�d
n�R2hh�#D��3sr1�e&14���Ћ�I�0���$ELDH&d��)wt�DdS`�2�Iw�]]����*�N�.��I+ˊ<T��ə�Ү�jP޼�9�LB�DJ�����ƧS���j��;�[4����n�Ͽ���諭3{��^V3��<�;�+��X��6��M�����!T�Q��"��Y���;ǉ�Gls��(Ce#��B�f��.ʔh@�~L�҆v✑˖S��	u�*��J�؎a���B�=��_<=7::���b  �o�ˋ�Pg��[����#j+����%����Z��!�,��c`v��lhm���ѕXE-��mF:�TM>��#��a�ѡ"�X�8�����c��a����Ν�]����F6ʴ/ܞ��@�U(�c�̄����6S(F@C8�b���)�g��U'ft
�&-%�]I�v{�=1�s{��
d�J��Cd��<�h_�ʡ��Xx��qҲ��өkQ�PfO�Ki�VY�Fq=ྫྷ��:N���J��)��:<�:�r��O��gV,�����W�YX}S�JY-�����%:�"c�'X(v��������Ͻ:��.��-Wi�َW�F���|���a`*����X������2%�;a���i�|7u��^�w�t�Ƴ�����\�˅����G4�n�
��:�]�{��ٌ6��������-V�NU*EW�wǛ�Q� ��\��_>jh��9�w'���6��6�0��R����o9C�����]�e������v(a�˭C5���}��7�,�^��9��G�8�J��}��u#������ۿ`�:>;F���Gǎ���H�A�;�8!����?-��V����_{��+�|�ʧ^.��[��$s�Tq�����B
;�~�øt}�xǀ%��p��Q��ʰ	ԹIݛ��~Ǿ�G=�j{z�5Oܠ�\w�*�R���Kڭ��9|��^:�	0���'M��F8	�ӾfFE$��p�=�
��Owɭ�;����}�m�����M.��̚�����F��\`{��l}c����Sj��¥כ������6��6�<�{z�Vƒl���]_T�|k�0�k��}��ӟ��u�/���4n�隽I���t����Pd׸�$�J ���Ƽ6Z���B��T��5%��1M�;��9��%�A��ŷ\h���GA��P���)�1Uc9�_J{�4G%N(���w�F��C���v���#J��׮aU��]���B�@��N=�k>���Uɛ>E��Oh��$ٺ�_C�J�n��w5�C��d�61V�Y9԰��X�����솣�kܹ|���{��3U_X�J�����P���u_-���v�Z%h�V�I@�S6�w=n�,uE�_�������}a�����4ȍY:0z%5_�ޖ7!��&޻��bY�Q��������V/ᨘt���:�f=)�h�1k�\��5hg�[�L[1aPۭ�;��0Y��\
�V����X����>D*�#���/q������
��J�ɨm���i�8Z1�	jc�s��������O����~@�����x�S�Y�����ޗ�{�/��(���c>�B�x���H����u^5`Xk���R���#�|����svUu
{K+�CF����5Z��|J�a�?"^s[����< �0��`�F��s��AOl`�r���,��5ӧ�l���C��NF���תy�wɒĬc�
������Ri��|
�:;K'����*7C��F{�뙋����:�~쫩}(��zޜ��;/e6�;q;XD,�_Tڬ�<L pj�K"�U�M�sU��|� f-��X��-
+2�Ċ%L�vc��R7sѽ�p�u)L�߭��,���W�eF`q0��\k��qO���W�)n;�-YcSk.]�t��#ģ��Gf��J�f?���
hU�i�v���M��s�XAm��6�x7R�sf�9.�h���f��1:OU�'�с��Û	t'\�ĥ]J�x�����������fܮ�{�����^�G��@pPN��_L\u�ak��it�ďN��n6�k 3]MB�f�E�)h��~���zT:(��� 뢸�p%5�d�AF�r��v�����$�	��_ؕ�����`#�ڸ|����P/��&:+��! UP��-O��e{&"E]�UN�Kn��@��4�>����mW*�l�M�Z!}C��<��nz�-�ޱ�(�to� !ik�
��K_\Uķq������%=�#i�!3=.�貪를ʙ�OS�b��@i}CG���cJ��|'��P�����#��pCg��K�xQ���v��Q�a�3�}�$OCtZ��� ��(��"�
N�r����GΈ�l��^yr�[�t���'�����!�Ɔ�E*����\���3M^��w�ɋ[��Q��|�\�3*B}(T��m;2m9��p�FC�^�������}f�R������u�w�֢sd���h��]���wr,&C���Ms�Tkʐk�OT@ɎѤk:�+���rxi{�)h�y{ك�.�&1��G�igpv��_���uum+�>�Fc�meQR��ӓ��42u���	�]Vo�K�LLv9�p�.��z�V��6�]�2��V�k����|H����kR��!��m,�=3�a@����ﾈ�i�=Ǎ�ć��.[�q���K��t1���%�S�N�2�E�����QWR#.�r�Cb]\s�����Y'_���l��u�e$o�1�0g�n�[��Ң5]A۽A5v��wݳ�u?`�x?}-Q��]��2�҉`a�	_a5G��%M&Y%�ҟGN�|.�ݚ��9@�!#O�|���Y��EY��N%�~�=���e�aݾ�`�Je;���)�733!���P9N�+q�����wQ�.҄����[���z��{ڣ^�У�6hv? �HE�r��w\�3|b�eJ7f ��?&r��	Nw��{�s�]9�GT��ԉ�ZC���B;~E�я���HY���M�s��_`a��N�qN�}��wڠٟ���cgL�)]TK.=��T�K1� ��=ꑲ{��u@uRݺ�Z���8�P$�n@椠&�b(hH��V7�+j�e��Ɇ;�P���ᛥC3�}�f]��Oy����^q6E)DC/2r�X��<+(p�]gG����q��v%�m���ᘀ��S�8�Ʋ�'�C�H���j�Z�u���k&%��
�-ԡ�h�ǣrX鼴ѡ$�n��9��5nJ��%.���!DG*�N�[��8��GڇAFd�f�ͅW>=�����!����K�=���]��9:��W�}��U&3�4&�3��=��p��M��˯7���<_5�:�"z&�^��-J�'���7}%���O>��?9j�0�S�/�*���ʓ�&c����
=+V��&�u��x=[�(E^�A�>VC�}S�4���,rX�S�B��02P���x_�g�&V�'+*+��ӑ[0�����Q��M A���4�8�*�%k�uz�z�qB���N��t�4}N�M��ǠRe+�p�>�Ow0T���S�=H���y�<l�C�����&:�p�6�3��ʉ�ou:��ĺ���<�e�\vרf�Ԥ+�l����j��EC�nN_b����R��{�I5�w��8a�rw�r����:ͽy�w��,��Nϯ�v����"�^��N>�9EGn�;�8߯�3r�b�7��ݸO;:��1���lQ���ԭrR�mY�p
����[N��=VR}�l��:箂��>�⽫<_�b�f*��E�(���1W��G������;xz�������ڮ�zՑk��٢F����T#3]5zq�R@5�+#N��#%�__�z�^�����I��5��Z����R�݄�#������<�\f��I������j�������[��3+��9(��y��_WѴ���j����{b���
���]a�p.j�v?����
*�_II�]_B�SZ�� ��S��b|7q�I�#4�mC�Z)-:{���P`w3����xq�N���//��u��Ag�W,�������r�

c�����+�K�5L�]Ѽ��@�J������ni\C7�q��O�Y�D.�%j��l�j*IT:5�3�O<��Wed��y�b�\r�4�|�͡M��vɱp��Y�Γ(d���Vڵ`508���t�K��6�6c.�̚�Us�en��C����8��L�Ѳ
U�뒷&�o���-���j�!�5SŒ+��B%,�� v�����ϵ��l���n2v����׾��o>螫E�s�΁��pӮ���j8:��F�7Z�E�˓�Ipz�4Xʝ	�ib<��V�g�9�\��U
�9�gE�Gu���%P���µ�-'|(��mb/�V�f]��K1u�s9�jL�w,hV���j�0��;�w�(šM�Jճ+6M�`�JG��CK��Ca<����P,ռİ�J^��ﾯ��g��vGWv3ɵ_nV;��}x�kY�uc�SF��C2�>�H��%��4�in;�u�'����/��Q���R�����Ś�w1�g�=�:�u{-m�[^��TY��������w�A�/�sNB��Y�]�57K5!��AN7���ׅ��=Q����K�Q��P�oopSC%dnD�ѭC�Eu9]�o:��dSG8��5��ؽ�Wc��5�k�=�}�VmI�އ�&�9Ox��v�����<��?	�Q��x�:����a_�m��t>e�ж���͵_
�ϏT�u$�2zs�~��!�nm�9�:t�jO-�k���}8�|�(��&��ʮ3�hwv��[��N
�7tT�>:�k��s6�q����qF.��d��ۧٽy��.�]�R���+Է�Tri\3z�t��F�����pا!*����};pӆ�85�%�����s�7Q�5-��3�ky���k�{����l.�����ϋ���d�:U�V��3N�2k}��AY����ܫ�����\ƹ𗼧YY�����ޕ�T!Ά��UUW��*�P��p_+�C�e���CA)������rt��Mn�T������F�t*g%���+�q�h�LB�&9��m\�M�ʶXU[�.n����*�Q��F��p�<�L��	��p�F�#����m_���4qo�B��)[�/D���Vr�|�N�m���Z���[�#s��̱���y�4��c̯���Ȏ����}x�2�흨o�3BZ+e˴�׽B�]O����*�"���o�V�O�+�E�ֱr5ҕE�����б/�b��L�GxfTAw�h�@���*/�=��N���b�,���ĥ������}�?�x�������J���O�'ջ�l�IL���SF5�q�)�عm����o��Tga�c���
m��<e������{��) ]O�]�4�W[W������Xkq�T��h��D�c[[���1Wf}�ٗ7�2'������Φ��6�{�j�!̉�:�[ғw�(,ي2���vr�.@�'J��u����}��%�6խ��6sB�l�YBdsr�&\W.�k��b�=K��6uD�'{�N�Y�?����������%�R�O��r:��q�.�������z�i��Zࡷ��z�8qR%ư:~;�����Ib�-��ߋOb�S ��U�ѸOR;�@��mQ!�|�(��LPԕ��O����q�	���V�&��&����J3�3�Q@+ﻤ�JZ(jk3ೱliq)ʳij4���_5p��X�m��r̢|�M�b�?<=�o�_�q7��*�����ޅ���|��b�sg!J7Qڀy�w�".��݋�ɔ�j�sF���jm-��n� �!��i0�̸օѪ��p^o��IS��z�Y�o�.`�̸�kj��յ��MQ��8F�q�T�,&�t��,G�%N�#���o���?g��������r{��p,��i��A�祐7����ߗ��-�������C�ʤ����-9��C����9��x�X��ku�dc/;Є�kQ��yf��g\6��x�[k��N��3^�+I	b�ePި��X�����{ԦJ1��hj-���m�]|W.j���R��ư�01~�h֮2��8�ҹ��t�j��١!;��7a�lW��$/�F�(��FTD�HƧ4_���䴈�EJ*�Y^��ݬp^�J{��C��\�wmL �պb�K�����N���B�Krs�)��]��Y]��gz$e��*��cw���X�\��Tp>��N�A8�w֎z��n®N�����7*'RvwY�,C�vyyB9[�dJ���6k2S�oF��$�V���z��ճD��l��ǂ�>�:���Fk,gR�������:�k���;��(n��Ot�W�P:��C�Φ��'x�=�C��GZ.^!y����#:EwMD
�O�*�+B��[é�����Dt�:�i�HqܹlnmOFج��D0ܙT"���*
�c�L5��JD��b�^��*C��̲O�ˬ4�[��0k�G����)��H�k�췭M�}e��6O.�;Tc�F7���L��Et�p���������C2��e�p��ު�=a���D��8r=�����x���2is{f-y�A�5)���{]*r�����nv<��6�]0�`6�n>��ެ[0�+���q�+�2i�umN�W%��r�cgG5��V�����K���P%^H)&E~g������ItѼ��`��ږ����n��έ׹�@�R�7v�-��Pf����2����L`;��)E[c���K�bZ�蛕m �H��f�]A(�`c2�_
�8R �4�	f�m����*�f&�y�nu���i�k�gu�7b�c+�nv��,|�1,L8e����x��v�V�͸����	�;:,�v�o�#�4�D�ȃ4�¹��w�{mӻ���bH���0F�B�m$�����<�̱�R�y��ښ�a���ؖ���(9y +p�To��3p4���wڌ!CRZ�88)N�MN�5��7N�}�QnYz���9Ǩ}|vt�$�3�>�<�s4���6�e���%��!N\�!,��tx�8u�wwv�_?�Ff�e=�b3d_���B�Лݫg7~pK�ЉC��y�*�ˢ�����&�9�^���vn1&Ŷi������/n�η{�gۀ\�"��#)�����B��.���ie�5y{C���|5�v���	���GV�$ie���o'>�e�&:�rU�>�LgΟr�)r�ų��M[�����MS�K"wGE�W�i(�����J@{\][W����6��uҽ�KxﻒB�=��jN���J��Q�����K����M��oײ7�l)�:�Ց��r1 r��Ww�W,e1�q�@�ڷ�K:H���=vR��p̨{bn?����꫹BD���X�A�BE��D(NEt�%0R�A!��2h&B�����	I��11�RHf�� �����4X��"!��I!!F�.n%�"L���, �!
D�܈F(wn�st]�ӛ�&�3����"%����77`�AW.D��S;�u1I�G7�I���AF�f&�N�)3���&i ��D���]\�QD���wP�nt���%wnE��EPl�	��D� H���Ir�D�B3$�}WUwu���I��a�v�p��j�'I�]h��-�C&ZȢ{|*, ]N=g�O��P��6�]m/�t�:ĭ���n��K���#��>��7�۳Rf{A�ym�ֲ5��y����j�S�œs���ؾ'����է��uc�yo��=땞1�Oi]��g4哢v,kv�^x�I���yw�g�t��nA�[�òOz�����.����,����&����ZW�����\w==��.�2���$�*m�î}���T��q��U�]�騫��=��5r�sG��(*�j�q[���o+\d�S�*����[N{^�A����͂��|�$���l���4�1�/jgނs��&ј�����y�n�B�LG|�`����JO��KX�����E:����y��/�K���m��)W�ﻧ��&+E�����{S��TMR����u-}���3z�"����?"#*��0�/�G�'��>�������V.9ɤ�|�͡M����"U��\��y���:��Aɡ��2W ��ߺ�ri���j�b��5y�5�zs�β��IW,���g\˨!r�N{��p��}��=�:��yX��I�C�u���̎�;��o[��:�*�r�樺�.�F�"3��0)��߾����Mvᡥ��i��.ȁ��^���]�q��>C).sM��*rn�u٥:/�~`�T���X���"9�g?-MgF���|v�F��h�,gK��`�n5�o#^1�tZ܈�OfT��P�]�0�1�-���ӥ��w.;�6�]��)ヴ�U}��k0-tf$��I���#n��E�[y�G��@Mz[Cw{����\5/��N5�r7��R�7_b���������|�}q�~�J�7ƨ�So��/Qo(�Y�󸝬F�.�e��qJ�5�2���.F�`��^���Py��D�\�6��m��lt6��Ǩ��d-�}l�	�a=�=�V���=R�0�:���t�PL�+��i��n���{Y]^眸��]��?U�/�-�#M�J��<��N��%�E̚���A�n�o���kg��WԀق��˔��%�[�=��߭(륱������u�'Sw��\���򖽎y��	q�O J݈��u��cT�_�GF� -e�Ms�!�e!��]���5c�+m]�~�3�V��0`�u3��Ff�
��\d�=H8p�%�s!�06#�r�WJ9XOt�	���}�u���Ç�B��C�=Q)Ѩ�M���5�B�m5{�����!�yu��J)O�[��L|;�<WE�{;��[X�g��:�q�R��$���B��Q	����P�P7�̀��k��u�6�r!�ѻ|.��/#*�ɭ6_��Y�����Nn�vw�=&�|+��e���y���Й;���_6�*�1��R���^y��J���铑D76���/�Vf	qo��6�6-����R�R;_Πs4;<wv�MN	�y����'�$^�v�je�7�-&&�Z�ȞCg�kEe�y����v�o�J�1w�z<��;��V-���%�p�6�o;�vB�o[�m�[wYy�D��1���z�'��ϻ��ە��j__؜2���{-�8=:�6gg-��hA��;6��T/���U6��J���ru���/Dv�L  ߐq�Z�zo�w#kr��f�G��4�3���}M���"���M�ҸE��ڨkW;Q
�LnEwf�Tab�\X�g���zfC�Q3��fL#��wt�*L��܋�2;���u,���}�p\����$�{qGG�}����i� _+�:�׺��QӀC�J�`�υ��D�D�a�����p���l����>�������1��P�lf�������u,�ŝٷ�᥊��/�=
��ؤ�b�7�*it��K}m�	�t��Y]�����0�O^��6��]\it�0���o���Qz�ٜ��ͿD�.N��^�p�0
��Kꏶ�J�j�Ɩ���o���i��F&{����7Ϟ�nV�Cg� ���	v�t]*[5�I��IIh�1w���h�/}�ӎ��s�1O�LAPBLW�RW�9K�{r���SR O^����V����n3���C�g�B�ﻃ��F��60ܦ��sy\�F�xR2��КLVw?�=�P�9P���	W�CJ����'KxoR�t�\K���ۯ��ʏ��W����㔫�Ϩl7�^X�Gh�n��e�ƺ����õ��˥pG|���0�u���?���r�h�}_1�xvQ�sՋ��h31��gF�;�N������p˸��I4��r�K��WrvZ�@�V��(�3Q�Mduw�Sr��1�Jp���U��V�����[��)q96����{�jm���o'_>A�}R�a�\k�����ƚ�yV6e��MK�C�s ��îb�Ü���[Z�����N��7�����d���<�5����{����Dj�1�á�t�[K+:�T+V�m�k:����?�s�i�9��w���:E���ۼ�Z6~�w�ڿ�?h�
���Ρ3�������ra���EC���kz[����zu7\Twl�o�����
��ȗ����+����;��}�Ү498)-��oS�ڲv;����	p�𨘾\�Ĥؿ�7�
�v�<�
��ʝb���t�JТ��:��s �,�}��-���7���B��gO@Sw���tj(�	�Mp8�Ѡ�U�7���BmT�4�C���9Y""܍�s�����"��.����V��?rB���)>�(��D͢��O\Z
��Rr���=b�]2�.!7*j�s������y׏H�˙��8��]��,�:v5ip# �v��,+	���6����\�^�����I�V�"��e*���c�h�N�r�3�*��:�d��#�Idu�����;R�5/l��O�Ė����F8[P�پ��}��'����u�9�^�Z*$�8N����-�\%�vk���W�Tڽ��n�YF"7mx�)�CչO�z����3೫寶ඓ�:��,�O.�P��#��7
�	QT9���?���D���X�1q���J�|��p�Orqj�C�?�ﲻ��a�3Q�P���|4��D����!��\��I99�Rg��ͯU0�N�
�3����P:�ܓ\�7���f�w�Q���.��j���%��n1�mk�'�C���O>���\"�ޣ}�0j�o%Yɓ��&�e>ok]b���18f�8;M�TF�7Q�t�]7��85�4�瘝��U�.%nTJz6�[��+�/��k!���yJh��Uf��ӑ�nӹ|
��ۘ�Soj K����r�;*^���W�7"R�1�n��ژ���!ݽθ$��3��a	���7xV�N��;����k1�ǗCx���t6��ҏ_a�y*>��3���@��1Y�7kJ�ݡX�
�'#[a>�;�:�9�Q4��Z��V�L�!���˙����D�Tٙ>�r�Z���ݧ�g�U�>���~�ڳuFe|z��_M�W�S�F���9��=�Uj����M��ݢus�zv˩���;,m�P3T�ꍥ\ip��<fb��VF��7��ff�Z�ܦڷ]��k��.��:�y��S㜼�:��]�K�-.�q��_<��\:^}��և����w�Յ/G-��]<v.��\�[p��)I����>e�[O:�_
 �w��:汻�L����f�X�����ٯ�O/汮������D{�L��#1F��z�.�;��Cg�����0�P7��9k��}�;�c�V�vE��Ʊ���p8���C�P
��0JZ#W;�:���q�.�I d��m���uy��^�Z�����öe���CA���Q�4�Y��*�Qv�?{��5���Y�~�*�5����#����v��V�)��*�?O_m=����	2���[r�����/z]�ts�Bv�Rᓵ5}�[l�
3��ܼ����F8��!��]��:�sc�D5D Xi̜�-��X�ދ�Fl
=�f@��v��j"�j����̏3�/77����ǆ��S�Wv�%E���W�V��.��t��Z����2�����M�>G"u����\N�Ԣo�i�ei��vPH��/�z���=��9�i�4ہ��]���HW-��6���(Q08�܁���y�<��}�kr��5/�18e8͇�r{����๗:j)��x���nS�J�8?n}Dt����;=l8Y�����}n��f~��CM�����(�w�es��*���=���*�􃽽���v���7�0�l(�^.�Mo\s�ɣ��fV��qY!*vڪ���⣻X��W��TaLT$�龘�U<f�d-���f�̽)�z�mE��\�Vs�+*$��p��+�b���o�s�[#$�Mիւ��VQ�L0{�s#�v�ʵj����z�1�k�5�pO.��=B�cf������>U%.���R٢��x��%�N��j��t'�r%ޜ��Sjzqc��JF�]x6y�t�oDٴ�����W��w��	x�cD[�7n�D|<yIv�]�=FJ�z���p+\� ��l(�M�㻕.m��{f��PK5]:�kqV땳��ZZ��*�O?���)f7� 8e��J�<㔥*�P���Q�&+�+��[ȳ�Ԍ�:|�s��������u<g+�r���S�wZYz�]Bu���|��~���o�ͮ�[7�C������=!,�Ό���!��ܝyJh�ed��s܀�������[/��qp�D���<%�fLiڽ�Ժ�g<F6��X�����u��ΛꖓC.5�K�z.*�[)�h��{�x[V�Xj��"'���J-�<�i�=V�:�Z�X}�љ��{cU�'ux�~�j�-��s��a�͸w�\�ه�wR�qnA��pӮ���<�;m�W<7Q�t�-��Sok������Y�����mm���U��'pT���kY�y^������UY�"��G�{>r�)��mը���<y�%����[�M�/_��1����&'@���{��\"g��cn���r�\��](����*�.�^*���;P;Ґ�,wr�{'H�HAO�\o�N�ۜ+=�t��ƱV<�Ҳ���jS�[i�rśSf39[�ZЯ��euQ����8���{s��}�9�܂��A|k��:lJ��\�%*+�nx�/�Y�v�C�¢~�\��M�-���S�����o�}D+��>8$t}h�K�?��%���alT-M�v�\e�ע�:�W����9��M����5�@��eAZ�RVD�ʠ����յU'5��Yx��i�ި:~�@hQQW����{�����j�����<9/�M�����c��9g|m*:b;��TR�ۚo5N�۷J�ʝ1ۚ�[X�>�-�ZX�dk�ꈶ�S��B��j��n޺�h��80��wE@�k2ΨZ�n ���z��ۆ��t��zOgu#:�F~��*�v����(,U�.9Q�W�o���
Y�fU����ē��'�P�E���R���Z�t�u�����8����9+�s+���&c�ȕH�CrN�X[��7�[��]��V!eu�-�'���r��R�#O.�u%��D����;K+[ea������L�k�;~������:���Zt����ά�W_uK(���o!9{Y�j�����I�;����7J��l�[��3��9���m)%J۩�,��`���[�՚y��xq�t�T�՛ж��9�L�[��Q'��/�W��鳯�:�Ƿw�75I�R�}�5���N��X]����m�+i��&!��C�WX�Y����V�*��K�� TS�ѽ�T���c�Q��.����\X*;����<�:�#��2mBՕ�b]���)o����]���{�ؤ�%��h�,b�O��6e[t:'S�dĬT%�\��9�Ө���$<��*�	9f����5����Pq�����#xs�t�p,v�2��CS�9��X	�`WV��,Ğ�x���;�`���:��Hj:Y���u����1	�B��R�;Y���N򦔚�xƅ�֞���뢙Y���}ث�Ӭ���,�k���}x�l�#���q�$ծ陬��*����5%l���eu̷H�Aby*�f %��ed��N����pkr�\��@ŲN��-�����E,��v���9X�Fb	TyQ�7w��(����E!�+��ݥ�˱�T���/��+t����j��)�.X�|�u����L�L!�_/bdn����P��L�2��,��>!x����N��mb$z�va|#Ř�wE���Ʀ#.�kaN�,�:��՘��U�IeLkz�TLSl�	�8r:S�G@�n�}0��ٷ�;ݹ�B��Bt�T���C%�{���Nf�R����zL�:>�L�E_3]Y�Ž�ZބK���F2�mN\�ܼ�]�w��2�B��� p��W������^�Ë�JcepeVe�n�wG����ӕV rT�.n��q*�t�}����=�}�}�xj꾾s~}4�Yg��>5��[�ǣtЀ�����m��I� F��-�eW>q�j����u���F�*lWc���$�4���ե���7��plN�:n�eВs@���v �YJ<;�����-�su
���X�	�m�a�Cef�n��24�];qW:�&�d_ S�8��0���컲Ty�5G��3�������T1�^nM���N��i��k*۵[�!uƦ`��R�i
�W��
sȕE�SO;�X��U��E���ve@@R��j�,ˏ���s�8���M���M�3���ofu�}��/�*a������2�E��+���i��,�iu��̍�n��9%ܲ��v��q�N�F��}�Nz��f�����o9��RǨ!7�����u����[���l�n���aB7Q��S����A�m�rD�z.�E�0?���fd,N���W캐W��P;&u %ɏrݞw��s�Р*�¨P��i0�##N]�W@R1�B�hP�PLDl �$f1D��1F&�$"�R�e0C"�RB�"�C`X�60�L�R�lc1*)BK��DC$�&&X�$�Hd�Q�E%b�0�&�	b"ɐ�$�I4J!M0s��1��D�#Q4��#�`D��Hؔ�FP��!�����eDH�P&4�@���X�#R �hbBR$@#i�2Dh�F̆A�1�M)��Bd�DB$�H����]��;��T>՚�qXO�K�.Բ����9�n��Q���d��]p*nԬ��n�����8��`�y��3j5�:�+�Q��>�io[j�}k�-����Tk"��y��U���h�[��\wB��"���_ҟ:�YѪ�\G']q��/�vp�/[��5u�^2Z���6��e}<�m�[���j_\bq�gϨ�F{�ڭ`��[QnL]F�|��WA�d�m��IX2�N[L"�����J�� �+�+ӫ
b����<vm���tz�Nj�:�%�����L�)�g+�h�2E�t�C0�~�[꞉�ss`���3���|uV.�u��..,��f]�]%4c\i�)���6պ��]���v�������m`����H��:Ԁ]O�]�k����x�z��}e�f7�j���&7r�g��7�tOX�c�+�9��ʩJ�F����k-�Z�x)��D�[eM�fc�8��g`��?i,WE�:{5��c]��p��L%<�L�y� F��=��&���;��-yS�ض/%9�iR��z!XG���sO�v�X�uLŵq�����l�ɥ����_VR;A��vj��O�>Y͠z�ٙ�սU6��p�ƻ���k0r��۸("�|�#T�OS�i�l�o��f!0b���p�І�8�PS�.��KE��Υ���}��O��`�~���co�;3k�5{����9Fa���)�Z(j��Y��f�57\r޳R�fD�|ճz�|�m�W�ٔB�)P�J}7*��޴��+���d�f��{���9���p�0�ȘT��#�9�;�ӕc9%��{4k�P�y���ޤ��������i0jq���vE� �	�n��&�S���Ϫ̛V�(FOa�����W�Ѩ�ᚆ�1���D�{��'�*��:�\�\���'��E���.�'������ڗβ38:��3���|��-	 \q��u�n�:��b� a��gy����s֥�f�)�7	�N��3����m�k#�����(�GxfT3�"�q�����]���'��=��4�r��)���u�kz��y�4s9܊�=�j�l\�5v���֎Ҵ���7�n3��0�vaY�J ���TFi�z"����dRR�sf����Au�lÈ��7�>�f���[�v���=���RJLJ��/*Ս�j����l��Y��;ٲp�(�K�v�1I�(����$x�ovK�o��w�ml�A�].'�� N��*:�
a$�P龵]�O�Y
�8��N��pg�>G�^��;˘������P��+�b������>���<ʭ�}����ہt���V����D��ڧ*���^����k҇�igA�#�2��((���3��މs���".�-�pl^�j�s_.�~2/k��ь�q��Ͼy�)JT(t�|�(���ԗMVQ�\�B����Td���}�z�h�o�ü�q{�<g*!�3�"��wIc ��J�u��/���.�6��Q���)�p��Y�{��g*�0�]"�wE؊�h=}���ͅ�0J|� &����;�O.w��(�hθ��p2�ғ�MQq���WF՗�k��[ɧ�:o�jL8;v2��N�r��ddN�9����U����"{���(������8X������&ב���������QӼ"εEm�y����i5
B���j��X�j<�`-I�P�;v���	b{ڬ��^9�G�&��C>,���5�)M������t�H�v��fK��X���Z#�]�:�3fj2(#͇雋�������1�n5�9Z�cz���ȗ�Q8���}J��+��\����6n��Vm��18f��9����vkX��[��f+�k��tnWEo���n?VD�$�9l�	�=^���i{m�rU7�j�N�T�Ǚ��q��S�x+d��.ʛ���^Fr��ϊ��.��'Y��8Mh<޷���[�ǝ{uu.B{eȾf�yQf*�=^��F��3D�طM��[�^����pָ�y�����-������.7dRs����P�ƙj�%�78�I���k��gu[���:��w;l�}H�<�9�X<����/#�ٛC
%��>\&f���	[z�\KO��P���ق��ȴ�a��ӞY�ӎ��(Guú=_Jtj#Rz�5�-��r�6�@����҃lߏ��)s:c�,��K�;���v���ž˄���q�V��r�u��mʷ��Z�;��(��Nj���[. ���;��ph׿]L���I�ލ�5�P]/B�۵�u;� ��ė�ϝ6�!��y���r�<��vv��:���9N��C�C��,s?)�%��������$�b�n�$�*t�h���邐�y]��Ǹ�p�����J3
�/�ň�m'������E�z�����~�7~F�1��I�K w�f�!��o	Q1=�\q����l�,�@)T@�J�5˶�y1��!��嗕x�](��.-�����̸�h�)B����*�`��Yo|�) �k�8�#��q϶�S�p��_Z�|ۍv��}��-�_E����V�17�[�G=�eD�뫌յ���u��3P���o*�ṷV��Nt\�Eu���t(`��VK�d�V8�%<{;���<��R�5�ܑ��Ƽ�j��<�V�b�z������E)���鷵%`ˌ��ӿ��z+3y�C��Y̋q��9S�Y���ꈘj��D9��o"�V{׮���5�7�h�M�������~?K�T�O�~1�í�Lg����T'?K�}{T-FymY*����ث{!�1�N˚�k��o���jR�ݙ�X�A�ۡ]��$Xpn�p��+bu3#��]5�����l��I�]�t���J�E}*t&s�ή�z�-lb(̀�����.��æ{�٪�.CjY����[��Rյ�q\�G�Tal$���V�]v��ʊ@l�y�	Yst`�
u��-�u=z�ڨU�]D-t�4�)�o.>m��t�Y���=�f+�;΄m�k�X݋�-�P~��������I7��Y=[O25���*����Z�M���P�<����K!]N���[X�9;�bI�/n���H.1��R�
7�z@�b�o5x����Tp*iW�5��~���I�/����u�T��c*�_!r��#{VT��0�Oɉm����޴R�2���i(f��pTCo*!�2�S)TyАHf�lQ]&��vmqr�7p6���ϡ���W��=}F�ǐ,>������Ŏ.z�=��k\@w'����ܚ��Z�u�M|�b�q��G!���Vb�$37��&}L2=U�<���c�/>Y=������j�:5���U`'m'b��j����0�1���*K-�)��ը���1C�w �nD�ћ&\17��W���WhW)�0��9��L�7�l�#0U��}��ؔ���@��k{4���<s+����b
�L��N ��S�*�8qC-,�k��jQչV,�~���E�n���{�(��qm#����cU�.*��n�~�(f'��׎��!��u�j����7���0aj�{==��p�su������'p\��i�Y��{׻������!�o�x̽a@�B���m6�W����g8��&F�}/Zy����2��F��p4����r�z��wS����v|���b�7�
�v�<���Q�[�&u����VQ�V
���g�J�{~�+���2���	Gt��sw>��h�z�l�f_��U6ʥ �g/��G�ʨĩ^��*2�r�s}=��#�T���ۃ{����!Az�Os���FTM[���5H嵥*�FK�Y6\}Qo�3dW�����P�*߬��^g����\m��{*B�9���:�>����[���:�x�S��+����s��ʭ�m��/�t�K;���zN8���E��a��\M �<b�r�˜���l�"�yJ�.���W�b�;�N��Nd��H�����(�L2�L��Ad���fj86Jy�}�&C��v�6l򌸀6m��Ժ�&��)MI�j��.����2l��+r�z���w9v�ҶoRyc[g*!�9V&�`�u��λp�h�C�(�#A���_N�{��֛��_2�;gۼ47�@�g�K>s��+���^{@���0���]�q��>BR�4�M��r� nq�cU�9
@��xd���{p\����pz�Qe�њ��h\�3;˔�m�_6�Z5���V��[+�ʑ�B=�3s�Ѧ��������9/N�'�<gi��vk5����V�(�܇y�%�]ڻ]�u�.%fT��o�����E��N5��t:�䩣O;_�k)��-�|
��nFd���%����c-��9�]i�m�@[|�|:I����7�_���mf��5���/�=J��@̝�Ԟs�L�w�N��S�0:\-��o:��õ�1�@ιs����Ɩ�8D�U 1 �;Ҵ����>��ʝ�n5�X�jfoVQ*�w�ʾ�#~[�8�U؂�a��G}�r�ud��IH	�^��ׯ!���������2ͺ��^n:ʹd�N�����ll3J�!}lW>jf��7B�s���3�y_'8�r1f�g9\33��OD~��j��m|�g����<��T��j�ZDh-�c�v;VI�-.�im�n�����O>�rϞ�r�����;����[1���{�F��l�ґ�[;�u^����!���W�+�c���㷸�zArﶕ?��������/d4�Rƻ>��n.��c�&v�u��(������\�Q����f�K_T���oJ�6/��ŧ"y��`<N�6v�r��yW,���\N���w��3o,��TT�\b�q���v��#f���yv��yL�(=��5�ێ�{/�heD'�[|�^�.2!1�lC*��9z�O,���j�*�H�%.%����&�'�k湃Pۍh^k�'�i�Z�,=w�C�L�{3��Ӟ�h��M�Uy�iuZ���8f�pv����t��=�e"���BnV�ܐ�ġ�7W2�ۙo��&JjJTѮ��
agZ��IX�);\�;�Ѐ=�=�>;�dP^^C�"A�;��3���f�|���u͏i��ݎS�b+��	�z2gu�KF�Hj
@f��F�k�Y�����:����%���W&��*����;ʲ)��>��'���Sf�6���s���Ͼ��	�6���|m�لl��o��{3!
$����[�q�%�k�3�-��9b�1ja�޹�o�B-U��罡d����y^qN�7���c#<c��?�G��?[:'e��O6�g>ͷ�c��W\uaLT$��oϦ����.+�^�F������s.:��8eD�U�ӅK],�a�I-:zW\=��������o�:�`t��GO�O&kf:R7������ˇ�oSM��F�"�XY��P.���3ju���B郍%����Of���[�d�0���~��|����*�&�إ��P7��Oӌ,��=%5gbs�|� ����~ے����9E ���=��py.32���#�,�Ö� M��_o{��
S�H����uoU���-����xb�1ݸ�Z3��]Y΋߳7ej�e�R�r��}�H�m��b����j�;!�3F���ܫn✎|�r[����zR�.����<_�����GUn޹�@������\~[C�[�6��ff��p-��,��8�S	�I�U1��ﲷ:��Q��-H��e����)Π��0xyedT�V\
���]r�8��*�@V�^|53�c9!w����j40�d1����dg�R��5$�ř����9����60�V��4FI��*�����ld
��{4�r�L����9,�Ѩ�6�	dZU���ێ�fO�^	b��Α�������IG�����<��d���V�Vu�Z�(x��� ;T����q�����NJ+9[���
z�ϖ���˴𜸣�<�"�N�l�m�«=�3\�#@�-
��w+b�W��f`�Y�\N/�q�Ԣ���Xh�{;ot���L��qa6Mӷ*�օ��Qnjú�3���hT%F
9Ϯ��ˡ �u�ɽ}��S<�><{��+=`�;t�-A�xl|�� �s���0�s�]0w4U�\,`d�E
[|;�2���O��>ܭ"��� n�.1�:g�(OX�*�Fuq�r���m7�m�ۈ+����@���C* �r��}z��ƷR��Z�ܺr	�YM-&PЬ�C�!��
�0WsPTD���zQD�J��;%FK�>=W9����V�]bQ�:��ݿ����{�V��Ϸ��p�����Pm��LY�x;����{����ծ&p[�8S �N�p��� ;��/X[�fL���4��5��LCV�jn)Z���Έ��D9�<6�c+Q.k�Q뵕��������]3Y�.�cWPo1
�vٻ�S�#O6P�,�uh���9,��b��h��4-Zi<82�J��dzT�0�K�C�|�)vS9JV��w׎X����0�������c�Y����)D�+�r���-���Wx�%R��MX�`1(�绑˺g"Zo�G�U��>*������f r��U�f��*w�a�Ȳ��f�U�3}K`ZB�sy:a�X珸u�����U�ӴWA*iG�+J���E�t;xWt����i*QhMExsS�%Ze��%|j[���V�B���-mঢ����K�����ps���v�� �zTaW\t^�6I_ɫG�P�k"k�D�7����a]ݔ�)G�{Q���؍�E��~d�]���Wv\ks�^��G���7B^�V��2[]��� �uekTr�-ޞ��-�V�Z��	]�$�]��e ��:ι٬�Gqwa'tr���£�ɱk���V��2�q���.����J�)��F���G�fPt�N�U��	�/��uL�2�m7��Ze�Pt�AVS�\�T9.hּ�J�F��X���dsoM	�N�ݞ{w$��h�+�@
��B(fB�HB LZa��L���F�S52Ƃ�D���D�A�cbJeݮ�4�b� %�	L�#$�P�%A�Je`�dRh�$��EI3I���2LM&`�BA
$��(�6�jB�4X��E���`�#F2S6)��0�"�0������(�"#bHؤ�	�E����2h(��HJ�����(I6#Ehجb�2�*e4̘���ɒ��,A"�矏~�<�~�x�hLf��ݽ�y�@(p�Y�AU���A�1������+�&uf:px�Eů����`dT�\efN)�oa7ټ���{�_ri1Z�<���H�nc�-�pD V��t�E���]�2f'{������Ϣ|��+g"U'4fۊ��z=/R�m����ٛɫܜ�}��P�T�4���k�Mn���,�2���:hT=�#�nـ�`��ﰿ-�|׌�=���^�l؇w���j��\olm7�_k�&9��kk�?wQ:��w-q�ݩWU��ԩ�33��}q�3O(�|�VЛ��|�b��|f�a��+s�lܷWv1�mT^�wK�i�Y��{׮Q��w0W����_�R�S�K���c��΂�:���;��6��	���ʳ�m�l2R��y{��Ey-O�ۏ	^}r�E�a$�N��U۵Ixd-�=�ĸlgz��ԟ	��C�V�O=[*N�ug�L�~s2^1��s -��Ӱ��CCw��5���L����Sn�Ә�,6x��蒤���U,}�޷����=�OZPy׹k�R����3xT��6K�9��~�W͌�.ms=�4�g�VD�Kͬ�+��x�(�]Xe�*��b��i�9JǽF����q�ZzS�4˗ཛ��f�c��`e�y���T��L��S���ȼ�r��*.��j&�N�\�ƶ�Ol��H��(�z�$�;7�|��NVmRޅ�����*ө�h>��-�ggI�{o�w*fŇ�c8q@��k:�	���}�x����[�j�nBq�P�eb�������)�ǻW)s�`-�5�����}�SJٽw��m�ç6�S走�U�oI<�jK�FL8�yl�ӫ���"֛��ڶ_�ui)�X�����׀�1��
��}O�k��yv��'O���W���I�}ШT�����ˍw�J��ɫ�����-��%;�$"��m*G]yaX�.G��t��z���ϗ�^|���Q��>��'����#��=Z渔�n���Y��N��S�v�ʨ׆׭��{�ʇ��wN��e�ۅƱp��۬�U�m�����E:��A�!�S	]�>��������~�p�QC����v�Ѐm��J���ܫ���gʯ��Ϲmb�H��՝m�g��Ĩs���%A��8�xPd��~`��:�Nwc]�`Ԁ`��BEǬk�*Z+gq�I��ݕ<�m��u�����N5��C�-�0�!���Pm0+��Uv܈{O�!���;뎦���tT�-�\��/ht�+���-Z�f���ܝ
����s�fʢ�V}�uVW8�z�Ξ��=�Ҕ0�~z��OMۮ�G�L:��D9�r5宵��0�B)�m��ۻ�εh���M�E6���y�gS�5��<8yJA�{�Jc@-���-t�Kuwp�|Zz+6F�7��ۊ�gsgS�e���ݤcͪ=Q=�j#y�������6����İ��7�t���T;���/�����O�;���r�CN�,k�\g��]��e��z�\t����;�:��	������m��9J>9Z �)�ɤ�پ�t���x� ao�W�3�3��o��׍ӫ8���-C)7Qgۯ�У�Ln��c��g/	�t���U!=�m^$����$��)}�Ӄ�Ǐ$E��I~�ݩul�[GD��/2�[�����iw�bF������9���#m�b���v�)�!T׉�m�"����N8t��u� d��s���Vf^lQ�2K�~���|��=рssv{5}<�r�f�Ġ<�9ټ��=�Ϝ�6�;e뿑ȘT�!�A󗝦���YK:�I��Z騛�ڽ絩�O��5���й�b���+ŀŉ�<�%x�Q�B��Q�gn�鶝\f��]V�9����[s��o�P��{iq���V�;ײױUɨ�E���y��U�O?�����.�[��BHMu�o)M�C&z����!l��;i���
NK�Q�yz���Y߾��jaTa[T��k�N����E�}�}�^ɹ}�g�N��xe����`�Z�f��ۑz���*�ۊm�X+�'����л=�2��>"S6��I6[{�B�͸W�{gu��an����k(���]q�%�F҅P�Ҹ�-������t���ˠ�+�F7���Ra�(\��7ԍtz�U�,����ҫ6=X�U�ߕ��b��K�ɡ�}@�����tOk�e	L�XXwVJ�u�d��*B���ut�2��7 �M��Z\Ο']������E��c+RԘQO�cZ[P,Ε}�h��l���yTI�ٓ�]]2�=�v�.��$o$]��d^���f�0�S�D{�N������������_�j(����~Ѻ2�3ҙ�x�vd�{oϤ�!&+�'EW@ћuj�n�e!�Uӛ,���>Ά�uC�q�P~�e�U������L�R�B��3�K{��i\C7�C���噄B��G`%؜o:�j�򉺵�0t�O>{����_6_p� ��r]�WT��*+1�-u/x��D�Su����M�ڽ���֋����i0�뉚yv4�=�A*&FD��8�O����+aՕ���B�����줹�������f��$�g��K�^?[���Z��;�/:��m�%��X����bԳ�=�zW}'�������iB;T���ԝӨi���a�
-��Nq+K���A'{�{:��qV���DS�4ٺ�E��x[�
#k�k��ޏv�;R�4�^S� ����'!��z�[��0�T��g=�pE���%Hmjbf䬴�
��g<�z�:mo�K] :h��)9	os)����3�!ru�0���=[98�Cw�dN�O�q�؝7���3�5�����w��6����s7_U8��u�a��u�ﳔLF[�eJ~���i]T�\d�P�8�'��ƯԹ	�۾^���TY���{_�u���2�a�{"��)\�8���A�1R�����B��[z'g���c�[*NCYH^���,N��
0���ܧV�5�Y����3ʨΑ�z��ub�]❭��z��Ŷff�����������7�B�Lrg�*�ePo�Tw�$�<�t�gw���D*u5�=|Ŏ�<�m*;�|K��jލ�s�!�IpT�=�ݦ���*����o��ƻ5�uC�r���*��v5oi�y�QDv��!�z*�Y
�c�	w8f��|�+����Q��ש	�+|߅��7� �D)������{5����b����M!��{�����Z6m��p8�m����taE1,��	��Ab�E�[(cF��A�W0�{3_��չ'2�.z=,��7��	�a��Vgu�qɛ.F*�q��y>�	[���b�	�ҮK	���g7]��8����u�o6�Գg�+����.�׉��C-J�S#�k�9��{�g�Y�(�ek�ɝI���X����e��O�_��f`����6�6cB�B�L� �Q�hDp�J�u��q��ݎ2��N����[˨��`��Dk�5�}�ji���(��J���G=��){{�J%3�s���x{�2vyx��Y	b$���{C��L�5:�`��k���p��#��uY*�X}/lg5מ����H^�N��w�����{ è�٤���'2�(wH��GW�r���oz�"$e�S��t��)}�>oyw�)��cu�1|k�)�Üv7� �n��ϣ�X��-xL��"6wf�/��������u"���n�K�H/�N��>%ٗ���B��U#��˓ǡ�>��q�:��׉N���R/��u��d��˙{�S���u���B����L�{beVz���V*n������q��J��(Mok���.\��^�ϯ�}A��W�|v��W�}����XK_�Oӟ�f����a�*��0fn�[@�6q�Ym_Z�*��n�q&pm�Fs5�����d�fmOE;;XK�O?�l�0.N:i��W ��Do#�}w�2%v��P��l���EeO�9Pm�����=�KE<,�PT�U܍ZB���9�,	�'ҙ��\j{��P�t�b��9�Ǩ���#���|��'��9ss�W���xC�#�I��$���"�줥z�'��_��E'βZ|u������uV+ܛ�9�#�������]=#�)2<`C�P[�&�=+��Q���jn�l�J�8��#�T�2�)��=�ԇ~�T���SNd��@�I-�c���G�V�>ՙB�n���ux�b��/_�F{�����Ʋrnr#Z�T�9"{Ɓ�l��"vv�K�Z�W��oZ�r��xK�ӱ�6h=�H�?K��Oĳa��'��h�d���/nGǞ{���(���>�6=*R4.���|�������H�����1;r��U�7�z�1,�D���b���^�%w��.s��o#z�놮�1����\c�L�������V=̕�k��4X��{jA��Z2a��'t¿�պn��>[	_��m5݈�� 8��kУ\�j+������o&��W*.�.'\y� �My��ph�`9ɴ�������U��b/��f����k��c4��*�[a�#䐥��N�,=�?1��뛃i���l/G%Ǻ����f�:QH\릥k-mmn� [7����F��+�T\(�D���Rl��B��͋Vsc�:��)��.���2���� #Cf���!`S��_J�Hd粏�[���U=&�}#;���H;Y�{=JѺ��p��xG��n�y��
Eh�kl���r��~����$�_���J�e������}C}~��p�,�h��=w�A�&s]f�7.'�ϸ/	�2�h��OF%����85�<˃K�Ϭ�Pͱ�~!�^���Ң��_K�a��	�k�d�ٖ2��>O��rN w��ϴ��vCN/��l�yߵ�;�}�K=[���梽!`5�=���,���~ �c>�����u��k,B�z�s�m�z�T��{�kh2,���~N�]~���99<������8�a�WM6^����QB�=աF�M��%S�]��-��gc�j���v���<��K~˃C��lZ>�7M�[:bZ�y�Fx�S�	��{��Vϴ�m>���e5<f��,�(!�R�C��i�6��.*{�S��JG�v!��m�K�wa��|p��M|t4�Qg��L�^
r��}�}^(�Ls�DO�|��P�t���#��A��y�\tsO�Y���'�����C�$��l��+'jhSy6j�QP�S�9Z��zz4�V�W3�;�|:�����u7���� ;�S[ L�E���i�mM��//�ҹ�aCk��}��ַ]˛��c�Ǚ���T�&���]���^T��p�0��O-��J�QVe��@�iK`�w,�P�ʚ�����X='�Lǝ��1Q/��o��k��Kq�w#���Wtg�V�_�q.� )j�4�TL���{���#��@~��s�,��������QQ/�p�>g+�v�i�n6��F�ۜ�lS�Ic�7�i��!�ӈ��-Lf��|�>�7��+�W��0��C��*M���~7ʍ����ܬ���3����E��Q;m�X�/fs����8��M�|���~ͯ\*�~�bzr2���'N�l�O�6)xE�bu��2����5�YJ=��^�~���&�w���^
�*_�&p9�YG#�<N_����~���O;`����VD?U���w�����hi����~W�?��'3`�{*�E��:D�ܴ��;^22���G��jn��o���@LZ7���#��B�mO�>%+�3=0��(�[���T!V�{<�w��u�_�JJ���>[-8~��=��ݱ�TπQ�*�y���zh�/��vyF�_.�uh�>���ir���Qe����~V%���Kc��%W�X$�G�,��|�驟��R
��n�q��^h߯��K&J�-t^;��38˦�D�t\-�!���N�ͣSSǭE����n��wܓg�4�ܛ9��87��5�f����8�5��fZ��yDU�}30����$��zI[��b�RF�9�!r��j�գjJU}W�-E��Wr�U��igG�2�z_��-S�����9B��qWmʔ�xv>麉U����T�hi�h�T.	!���ѫˈ��ڲa<C�R�^��vN9�й/ ��ɺ��W|��OU��!}�ݵiN�Z�QL8o���;���TO�3��x���`	��I>�r�x,]=K�x�8M0��얢���.������>]$��%.��n��$s���X���6���}w5P���ԨouѾ�2V����,���
�#un�Cy(��B�#"���:ni���`|�E}7���4�EK��@wFr�i���O�����J�o3��(�?��A��kUh5ٜ@��/=Ve�λ-�
ׂ�ևǩH꼡O�jX��˅�ڛZ�P&���{�B�v�Q�0p걯"�V��m����v;�i�Բ�)�ɧ���(�Y��P��
�P�ޭX��5&�fM��|	�a����=Jn�Q�+Ac���/t͟7��Nqt���|o�L<\�m��#�yYT�od���J��#�	ϵG};(��3!��mcUnF��0��ތ\wι���O���4�\��[PP�� �}g����V��
����-q`�3�G�9�S��b0�z��*s���4\�9������U)o-$� ��'{ڍ��1���=�b���\9�|�dߙ�=is�w����q��L�З�YK���5hrcs+��h2����;����u����E�01Ù�e'(#BKZ��f\�ԥ�S��2㱙L�Ǖ΃ȶ3T���UnX4�F�R���8q"�r�M��J���ue}�s�7;l����`1�1����e�Sp��N��k�Fs)#&�G���S��ڋ��Nwgh�t���f�Kw�k���sBR�Z�.\F���`�ܙ\���v�:���o.Is��f\�޾�jZ5�m����6�e��yj�����O-�Yٜ��� �Ԩ�Ť��YĆ��{~��Jb��M����anȣ3�i�
��o	�6l��Aѧ�j�ѕ:S������;[$�����. �q��.��z�kE-#{E�-�JN.���ӴŇ�<q�)���*�3�\}���[��'��T��:M��m4�6�iܲ�F40Gf��;�bms����KJ���O=A���gk���#ʵ]4-㾐�پ�n�N�K�z��:F���#�ݑ&Dﺬ�;w�>�#�9v�!��x����ښ��Z9/_�P7�
�io����4%�K�p;�V��WԻ75�ې:I��{S���[���B*C�u�0s��7�D�_~~�{�����~��6�!��L�Q�f0�EE���6-��1���`HD�33QR�����h2�
�虡�"Y2d��@bFK���d�F@��25	�
4�sD3D�`-&�!��2�h�R��I���#1���D"ƋBbd�bF3�X,��&,G8�!����D��h�����\M�u,d�p�&@I�v��A�����ڥ7�&���a�N<�wl���#�[��;c!yr�f!-3ݰ+
8�9�$.�����W���z�-��U�Qs*�G~���
�gǝ��W�߸�yI�|s}!��j�}�gw�6
7ۖے�����Ü����}Xe�5y���:��N}_&�ёa�:��}#J�o�'^H�l��7~�J��J'��9�9���"#^��ݨ��ϖg�΅p�և�}�lg�:�9(�y@���C��x$��}�\O�:��d�H�О&'�^��<Z>�F�ֲF��lL��B��u<��������d�q��m����z�Y>�[ �l��"e�z�Җ�\�^��8ss.�ñb�8��y��~U�+����e�F��9#�y>\N��R�l����$���S�H�^�oQ��U�b�.{�ѱ�=47��w�>�F���%m�'����.*��o��~w.�lN,j1�+���������hoVP��:�y�KF���-��e����Mț�	pbY���4�.b�������^��t�;cvz^�d8��^ر��5�9"��s�U;d:�Tf�k�w
^�dT9����|Ne|
s0��7/M��9�~ e���l;��K�b'�2��b(M�����]��_�R��;��\"'9t�g�[��񥯙� θ.���t��՞��w0��/h�x�i\����T�E%���4m*���{zD��L�4�������#�ɖu�����2_t���E
�xv}�Wi.^+{�0�w�X��4��}2�T].'2�(u��G+K#̝������$��O�-1S���/Y�7'�b��� ��п�N���(m���Fz�P�Z����t�/��yY�;�3ı�.Y5ܹ��)�l����3m�z$^�G"x�w�wqqwUT\����p٢�<�.�D�!��.]�k�����pi�^�ϓ�|U�IP.6����+��A�B��Y�>�I��x	�R>*��,ʖn��s��p�!�cs�'��۷>��������c��*���'�IJ�$�JJyz�'��������gy�A�ӱ��m0M��r=�n��q�'M���;%��D*�0�/�t�5���{!~2��D�s�2�7v:�����ޯG]�s��i�_:�&�̗4���������Ӝp�VX�������Nyi���f��Tm��|l�Kg>k' �m��SVʞH��ew�1\�*(�n{V<�Q3��O�bj}=㱸#ɲ�Ѕ��,6��f�X�v8�DOܫ����6��U*D1$��0%)&`c%�5��|�����_s��;���Ag*�u�"5-�����j��q�+:� �dI�5}[����.[��aSP�D\��ADa�-�1�mJ��4k&!13&]�k97���&�m���.�-i�Ty	�>C�����8o��S��V����>{2�>�E�����ҷ=U�.l�O_O��,3P`j�(���v@Ʌ��a��koFDV����c����'��!w2��ݍ|�2@�2��؅���TPג�ΦO�E��aߥ�a�>]��>���ƷپJ����8�5﨤�ǰ��L���]a�\-5�y5=W*.�q9 A��5�̑�7/Ŋ�S^�]t�e%/sl�dӫ'�Ƕ�x)u^�sΣZ��u���TnM��X:v�^��;FEyK9n�z^	��!~�T͚�"Q͙p+�^WϢL�NDS�2���r^�G\����#��e��ԧw��%x�~�ѕ�C��J���:S�l�^�~ۧ��s��{�g�����r�NF�^�_���K$ͨ�1�eK7e����g�S>F��e��U��}^=�c�W��q��_�䙨K\"$�[7�WHyd�0��Q��N���
�2�R7�u���
��ǝw�*��ܚ�{�<П3��{�Ǵ����F�d�8|��M6[��6��0�
���*����5Ʀ��03�ww�*������#�W5+�f|�����ww��c�f=��O�'��6~�=j���ݩ�������[���n;�8��T��ݦ�� oa���yƶ��}ɻd�vD�,��|��_V9^�5��xO�p�
K�nК\��Ⱦ[���j�p�p(����$0�j�FO^	>�3�m�7@�/ |=/�Ʀ/��O�&�u�M3�>m>��:Q��+9(<lޟ�L�V
�|�iwDR#eIvt@�~,n���7�R%���f�{�|[��n���إ+w�"Vz�y�x7���#�8}z���A	����/�����dm�������Y�ϟ�f�`�N_fC�Dz���1�F�ϕU���vMw�������C*�>�.W*c�N��������%�;�ˢ[�aǪX�71q>l���<���z�C�g�Q_K��9�l��C-{��J����]7��<����>�~�<�����MEk�P|Y>Ϡ�v����?�EB�b�����.\���>e��K�}��	�Uq_k��7{n�u��
���=O=bh�����מ���$���8��կE��Oi:wO3Y>���^����{޻�����;Y�g�Ώ�%�=���;2�rs�>
�l�w9G@�>'7�Ss���}.����z��:l����ug�Kr��Uɪ]�J�|J}vE���7 =)�7�r�.ԫz�fS
�T^���b����m�cMi�d�9p��.�
|X�u���̒.���Η.+��!=��.�6��Ep�:�D88ܹi��x�ogSj��u*�n����*�e�cN�)(�'�:���q�r�׋'2�C��ѓsZo�N���4���xȞ���aX�Zɼ�8_�A�]�[��n���O���+M>%+3�q^�F��tr.|�}Fjﴍ�d����X(ӱ��;"�����^~�CÔ�p��eHۋ�I�B��2��R��rT��s��l(Ā^�>�\�����Gd4��ǭ�t�O�����
%gХ�OnҘE⸪���3.F��7P�)v�=u+�}��Q5�����ȳ�o�;@<��*��vR���mW1����GР��<�R�f�Ke��s���ӟD�n���i�bΡ����0y����l�"�e~�|��ɆPO� �-��g�y��@s�[�Z2'�v�Cm��*3>��=q�{�]I�w�w�N����Ai�.B�(��"��u���hu�G�j}[��8�J�#r��j&��롖�K�YM6�b+�n��}2��=$��9z߱�s�5��z�V��i��k����r|۟Av�x��f�
wNL���e���SXB��6��8H�)���<*uE�b�it�5�!���i��r��d��bX�h�[#ċP�����T���]�ή�݈f�&^��%p�hr����DE��`��x�:��G$,��(��ɋ8۾��1�p�g[�]r�0���j�d�5�7�?{e�i��~s?i����|�e_/2Q�ۘ�w���.�=�(Z�k�$�Ki���XG8���
�V�[�������<�O�h��KF���e�l�賕&��x�.�C�,x�f��}?��,�ߥ<9ܴ�ѻ=����q>��Ȍ��֧�W��|��-��=��X�o�E�wr���x��9�ꛗ�����ODFϪ���T	˷9�S�V<���4���=a��f��}2�T_�w�� �T9ɝ9ؗz(�FX`r�VjВ�W^�%!: �c�.%JnNC��]9�n�X���Ʃ�=\��6�闅���>�of����RX3(���}J���r�y���}�arɮ�̽ϩ�l�H�����r){U��t�f=w�V�
�d�&��B^��I�
]0�v�1�\�4�K/��>�}A��o:]�D%����ǧR��2��}$�(	�"��R�x���z��s��pȏ!�c\���eװ-=wK�E�㦽���}��a���$���`�vRS��Q>�z�P��:�Q�y˰mP��Lj�n�W�a�jL�o��]��-��k�d�P�����8��:��j�Ҩ�Y]9��%o>= ��r���+S��=����j0��s˥�P5'\��L����Ș'e�W[|����h�+�
�҅�[�!xD�e<�I�"��I�;Q]&�ѓ�������*����˘}�,� {��C�/�t�4�3؅b���=�$�ٞY�=��Ho����\UĿ,C#ӕ�{}�C�����q�&��sH���E��#|��j���֓�R��q�;lC��4o�FP�:�,���g��lC5�;d���_����m��7���>������H�J��S�to/��܅F��&�Oĳa���q����}F\��ڗ�x�Q.���Ϥd���{ƅM��M^�{M�*}��H���F�,mdz<s.�3ݑ�'�0�D���F]M��tY�!; ��n3�Η��6z6�z��%�~܍�~
�������j���%C�qk��*+^J�:�>��h9�{D��5>]����[1��c���_vbü1S��͛���~6s�eu�����ɨ��QW���n<� s$v�m��SwO�ײ�u>����S;���|�}�]N/��/I�H��7�A���صs�r㥃�}}���{;�B�o�K8Z��<�_M��u��d����rex�e�3���r^�F���3�FdT"ktP�C2��V?'��M^ȅsFT�y��[�yy�p�7�t�n�����^��v3��D��>yu�U���1=��˻8/� A�Bc ��e�Z�ض��v0�Rl(�2&o+aU�v�}�b۬\��y!��6�'2�٣��J��
+��t{�t�(^	�
��tY�C�s�`+����/����{�G�CCƀf�.�1G]��*GՏ�r�)UMʝ4-tA�2��Tϑ�rk�ޫc�%����o��s+gt1�eE>���יY�����3|b�eJ7e��f�A�L\T�G��%z����޵{�=yޯe��i�VE���9od�m7]ND��W�H�J��Á0|�-�â�Kݙ�o�^s�z�B���{Bi>�i�9>sپ��=��mêa��V) yJchͦ�գ=��}C\Q�+��]��gMFx��?�{��Vϴ�M��x�FSS�s>�{|%l�癣m���}�u��1�Wp:_���TF�H,�_���ζ��zg�߾ۉ�u"��v��o�f�Ϣo�FE)�8��φ�y�<���E�Qz��歆&�G���-��d�\=��;y��Q�Ζ<�i=l���WHS��	:��A�NNNK]7���W>	;ެ�1t�f|B�30�},�ฌ~hdD���A�.'D�7�w"~]��Nm��;�n��WW7����I�oF�k�\�KtZ�P�7c�W��ro��3�-9X݄E<��+K�:�L�gwYb4�5�@`����<���ڍ;���i.b�k��4Q=�D����Dh�ʂ+��<x��U��#�zy�q�b���𩆙Q5+9.&�F�������p׺�1��ɫ�1St�4��S5�3��'� �t?�O~jvuF��o3'_ �����V������r�����x�5���,�ݗQ�֕`}x��W �����ŌzbY���WQ�#k����}=��7W3W����^|���{5�鲲�*r^��KG���´͖���>�����h�`}?�r�zz"r߬8��yۃ��ڑ{ޛ���Ⱦ��l�顛���1{yS�Nf���	�,\VMi�.�M06�.�e�JǮI�Z�ٺ��-2=���Ͻu��������ڞ4<J@ò�7�z�v�\hն�5v��.�>��f�C���dZ�M�l_���=v��ȉ��K��m��$�+�lv2���b�d�ł�z� �>w*��uP��/�E���7����il{D'�v���K�iw{q��b�y�N�e��;*e�|3�Yu,�C�V+��iQ�'���c�{瞡ڟ��ax5�Y5귚K��e��;�e�0��-�0gT�6�Ϣi7^����x�藻1�E��[�n����Y0}Y\ pV�m�0lx6��_Q{����`�����n�dF�*�s=mZ�ˍw`�����q�Ffr+;�"҆i2n���T��ѱ�n��Jۀ���q�.�S�̽�ؖt������uqE�����o
ɪ\/��o�ocr�V��t�m̲:�R<g��{�
�!�}$\��;�΅C�Z7��L�(�b.��wzI���?+u����M���M�t��(���({΂�ҥߜf�^��6����N�7�=�4�����K$h��WC-x��2�8�m��Pv�)��iz��ٳ�B/�1��T��2��b�yQ���v�]f��D����NM���̰{��ӓ4���?k�����+�����ۻ�SXX<��Ȝs�v������~wrq��d��@��j���q[����˃����p�i"��8�?Z:�)��Zt_կ���;��w�!?]x��bZ4a��z
�->q��|O)͛��e�Vh<O����9f��O�t���g����8ڦ���k�Gn���w���z9�{ʬJ�����l��n�⇘9�r���zrT�^6�!�M]�tR��!����r�x���z�MFi��'�YW*.���s(��a�o5Њږh��ѣxH��,�����,��#�T���;��қ��{m�:��'ђ ߚ�6n�C�B:q��
��W ��wVh>�s�-<�QrD���{��<ؽ{��0�HXˆ-ĉ�b�}��J7O�!�ٮ��
���q�%�-PQ(5%֭4��oN�F�ZZ��ݍ|�D�Xt��gnQT����Enp�W�a�c�ϥ�ΒN���B�&F������|����WG�b�0g4��B����ض��va蝞b�7%sG�'y���옷_r���X��Zh��M �ju���v�â�u���h��������q�L�Q��z,\v[J�L�yl5K�3�V��*i7��f��7O���oS*��o,���%F]���x�榪H��i$9
k���t��.f|���O�9g����R�;�����%�D+�(�m�D��0����t�u�d1�7e
|��ښ�5U�n����RU����
��R�+z��	�v�\[�}�5ZT�uWa�J���mQ �����u�Px~@����'\����J���ޓ�mI�lO�z�U��+6�.��)�Ù�>��u8
�����+ݖsm`/C.�+��P��ԥ�[�s7j��~4v�v�Fum����s���@�zha��\�} yw��E�/�kS�aU�4/WQ{���,�]����#�Q�V2��v�.uP��w�i�P�Q܃���I �V��wv�����SN�E��k��*�Je�a���|�i� ��!�8���[�r���>ܕ�l�Z�<)��B��^h�[�r7���29�ƙ�:a����xC��C�>`Ҭg���T2�K�gg7GB;���`h�U�IJ��0�RNܽO�R�m�kXF���â�
�+�W+��qp��^��x\�tҊ8��菸��6+C�&���`ZU�h�왐R8���Sol�A^�n��M`|�v�0K�Vu�riW�
���2v3l�%ݣ�oɗch@�s(+L�ޝ(Vu+)ڙi�p���F0T�9���jk��]o!�\Z��*,�x��FI}��_2���iR�t����������.R㻌�=/��� 2�U��E�FW,�S�@�BnΥp`][��t���9[w��w�R'�Z���1E��q�,�l7�d?R"&��}��*,qC���7
��G[��b({�Y�Gn\�˓�5/Ҩi�����F�ܖ:�ݲ9P}�k]5�Q�E�@�KD�y�
�7-��]ܻ��3]wx�Y�}ze�Lt��R3F"���C47���'{�7�[.J��`�vN��"��Y+#l������U�T��vsͬL͜�h:�;���2LE�Zc1��)⏙�՜�# ���uMgd�Ӊ�������c���`�T� ���j�]�;`�ڈj�TR��
o�Wΐ��q�.�+sS� �x��\��+��|m�t4����\Gb��Fk�=9E}���N�]|oc�	S�gY�w�?������@��q����"�	��&Q�%$�]F�j�
��M��`�)NqBM#4h�.��������!	y�
i\�&hιݹ�y�a+�t��1P�;�+��wu*^uםwut�s"�;�9�';F���+�ۻ�x����<1�]�.b�o�S4I	���;��F9�]�*9؛&�]����:7ew^u��)�ɤ�us�<njh���O;��˻���t.q(��g89��.���2r�q�w\wk�B뫻�w]%��w2JD]uۙ7(")9nn\˻����ݝ:7.��NuK�$|��(}�ӥZ%��s���:�T�s�����C�5�kN�r�s\i�����l�,��t��[ے��6�EV��46�����Z��Vj?�ˡu93�d���jLGP��]˙{���[�Pͷu軟s�EwN�݄���7듢�$�}2¨�3��O�����K����i��y%���i��	�f���g3j����ף3|"��[�5��;e3B��z���c"�R��Y�,�Suby��4dû�=���%Oc��4dg��Rx���ǻ �xø�\�iU`H)* 줧��|6,#S#�=���{�Jl�]q0}����o%��s}A���u�%��D a���u��d���s8X�^�W�Q3�k�#<h}��Bi7�C=9^G��z��o��ޙbv�sH�����^ʬ��EEW2=6�A�)_����5�葕�u�l4�Ke�W�9���w�#P���k���J�������6zH�n����4xv��r�y���m?̀��K�>�5�g���R���c~[�1�?X�����QJ<�u`�s�4/��K��*|n9��zߕܘi��w�����2�2}�z<�'�N�&|x�GnBvD���Y9<Vz�A�\���~���k	����>����[g��1W��B��s2_)+�|��Yy�q����˫M��Dۖ"��=�
WVR[{	�ie���f�n�`�����
�L�1����!�j�x�G+@�	���RptOEW�U+�"!3waR�l$�ǣ��*��U�8��<�"���~+9^}x����������E*�e��{/pɦ��?�Ӎ�r��[閎�H���^	�{�V.�H�,��p/����k�<�'����Y��~^Y�����<[=�]N$�}#;�zP9�g�w�S��9�?aŬ�V����bie����t&�p�>'�m.~}!�t��Y8%�����7ʔQu����i��i�PC�>�y3��8sf|2��u>���4�yN��Xx7O���}~R��-�7	�$zѿ;W���b���M�e��pe��g�3�n:�^q�Xx�+))��:�K2���MT�`#���79�g�W�"G��x�$��P�d������%ߝ�R�����/�d��k���ެ
=�}����}q�[�l�]E#�?x�'�
"�:1Y����u	yp��i�������	��S�m���� ��T��uL;�%J��ZfF�{f��'�� �@]\�:W����O�&�M׼l4��il�;����.���.�?���]�����=����U�LQ�;[1W�nV�QV�қ�;n/��=D�58龎�ck�޾������:��]�4�2uX��9��_G��k���#�4]�:�I� ���㴫'�<RF�����|:I�Cc�C�i�ޙ�G��>.H��끿�K�cX8��j�E��1�{I�`�&��G�S���q�E�%�:i��Q?rG���Q���4%9^:��_��dkʵ���Aڥ��x&%'�q�:O�~'��¬���8������;#�_�(|�nX��Yț���6�lzݸӞ�\��|�U1A�K%�)�k�42"y�(2=,��C��Q�:Vݝ~&�y>ך���3���i��cv��]��)F���O��8�.��QZ�T�d�E`-X!��'t�9�T��sn؜Oaag��Z��	�|Z:��7�m����v�k��7���u����\�uݯh���,�Zǖ�f,��p�n\e|'��N����{]A�)�1:�M�]�c�ޕ��Fo��з�������h���>�᳡�T��~'s�T�������`��ą�<��bw;��<���V�Ӿ�1x��Y�(e\�4<x��(u��z2mN3��y�ջ����ۤ��z@�rW����/�]{�d;�;�|�������gĥe�?�9o�5Dc�m�3I�&�ݿ�4ͩF���	`#�_�GGr�xHJ�sy��)2�' 0:�3³�g&��W/�r�,�x-/a��9m�Ve,�v_�,�h�h49���{���9̴��RI���z��rt���N����jCi�\�T��ʮ�9h�߰�dZ�M�m��<�T���
eHۋ�I�f7\ڥޖ���;�p٢�ŕ�1A��i1�ުcK����Yyc����=���׭��0�ћc�z)�5��J�L����S-φ|��Y����W���G���7����l�̸o��\ݔ�����[�9��6�B�Te�?+�c�e�����B��ֆ��%E�7O��5�M�X����}A㠱��v�#�|G� ��-��pzW��3�v��9����{��JK�*oO��{N7�i4��Zh:�D�3%�D@n�O��WQN���sb:���h���f߰�!z�?Z�����4�Ļ��Ķ�Do��?rM%p��]X�`���z��n��7��L�0���5>]�o�6_����94�HxO��ցN�ɖ)>�3W�����WȜ�R�5�8�jȜn_�o�i����o��(��1旲�d�`��Vz��s����#�2Y�="�6�Zt_կ����{p�������|�O�7���mI�_���]'6��G?!�Uu�,[C�M�2���v�h0α�e=�q��v��[�9W��׃���5�P�ʜ)�5Q���=P[�M��֞׽1��T�A{Y0�`,��c�ñ�p�n���I%<�ڛ��r��XL�vKT܂}^R}	O@��z��a�<<O!�X����OE}>��v�g��1��T���oQ�R퍏j��k���^�1�EGM%F��9�P�0�V���;��i���{ثΣ*��mע"F[�8<��g�y�Fi�{>��e\��\Ne P�>A��3���6�RU�*v�T���"V}��TGD�M��u�s�� �{mG$�������g�����qB��2xy��̕�y/ip���&#�.Y5�r�^�A���νC5���N�=�7����b%�1�V�EZ�:K��Kc�JO�P��ʻ\�u�.\y%����{$6}և��V:���I�^4���e_��(��H=FX �$�^=2���n�M����!�
~t�t���jMQ>C������=~��~0� \�iU}X
D�����j��EЪ�g-��{�/w�����ؘ���E��/������HN�.a��䲀��� ��eJ�T�Ϭ�w���3KȐ�Ҳ�ic����o��f����Ѥ�iF4��2\�&<qS}��/Q��۶��R���8���s�G�a��̭ɗ�J�
���(wN{l�т�P*��X��PMz���EYy���5u&�dҷ~sN��Z��r�6Z���P�s��`�;p�l�Uơ���|�>*���/Fʷ�Gyf��o\w%l��rU��> 7>��H��up7�Ƚ���_v�$e�u�l��l�l���BY[1�ٗN�S��˽���:�>S$���zH��ޤ*�SG�o�Kf��$e?S��~%�e���>���HT$��_�ցNm)zk�3����*��5�����;s������G�)=D1��E���k�20itQ6<x���mBvA�d�gӝ/MLK��kd��m[���.�x+���!�����J�4�����y*�L�H�C��wL)ן!]>v�o9�����y�g���G�]�s���_���0��j�i��hZ�����:r����{���\��{>�ZY��n}�_J]�ᱞ\��]N$��_�w�� �콄[ϏMT9���\����@R��^s����g�k��C�ʭ /�DdˁQ�����i����+�̥�ũ����$Vg�ho��,u?mc5��-]�;%���t��t�?r��tG�a�pS���r~���̜�{ ��=z_��\od:�b���M�d���|
��BR~46�c�'Q{0X�ʉ���w��n]O} �]�2����V`.[ˮ�|kz=w�jBh3fR1tE]�]z���*��4�N�9��!����Y%A�u��v��\-'���M� �]]^�גZ�3W-Cqxz�c٬��9����9JC�k��E]G��OA�yz2�r����C��nee�z��񯌪bc�"�c��ڮ�Q��<<���B�N����"�|'�;�{����[㓓�E�"�)^Ұq�7k�Ys���(ʆ<!�}�B|��^u�� ��	��S�a�/����#���J���=w'��y�C[36l��U����Dע���<����]ǯ:j3����M�{��J���m>��jL�Ad��?O�cl��_�'�>HiA��DO��p7������7�R�Sf;��M���u��Rd��F4��m�YA̲��<o�J�&y�LX�t����=�SQ��{�Y8���/�Q,[�8迚~��&��p�������GA#�-�'��.LS�1���C�bUW��(��.�|�L;�vG����b��K�S���"�9Ԩ:x��*;I���n��g#�뻙�Q�֠���>�aX}��h=5�{N/�M#W�b������QZ�T&(�8(%��&y����I�#�cG�	����~:��=���o�h�P�~ۨ����N2�kF~7�L֓�P�.�x��]{��%-x�>W�9�^�%*b|ٵ�\/���R�jRk�����w74��t��l�[^d�Sc�g Pq����5����ձ�=�տ^аu���&̺�N���v�E�x{P��J�#�(�+��ݙˇ>��p>����O���/�:�G���ۊ���W�ӎ�=q�0LE�6ǝ\q����<m��p��Γ��F·q9�_��S=v����%xd��o~�'
��1����}%�q���j3o�u�#&�t�,�ۃ0��.+&����j�S��&��gw�В�WW�1z�?R񐾦�~=u����/�((յ<hx���<:�
���6U?Y�ǳ;����G��S�(��j���2!v�[)��W��z��ueH�Zat� ��_�\�^D�>�8�.c����Y�|��X��ᷨ����'�ўN�h��lS���o�M(��l�g�'�&P��w2��d,��m۫|���G��ǵZ�B8t0����s��8�>k�-��q�`�(҂�,�
W���l�^uN2�D�
�?C�R���ϵ�RS��1��]�ŝ��Ae3�u|"��J	Q��-��g�y���:�u��{��{!�VR������q�ϴ��Bî\�?qG����酤Ԫ�jo.���8�fA��)蟶��G~�b��Z陙��)ߜV:~���3��6�چ� kd�ޘ�����bT����)��8���H�>��������Ŗ�p���n�HK�jo7��6��fW���k�ؗ�sT9��6)�ة�J�W])�)��-*����Q�^��`z�]Ƶ�4Z~vŴ�Ļedq-����S�4�:W�}ei����k��9>�������Q�|.ods<9�H���94s�-�q��g"=Y��5C3�o'r4��E<\K�%"���VR��9��~�d5U㌯&�7l�:��� �`V�fb@e�F~��&ףk�j�J�����v{N�܎���Fg%�ʗa�����)�}�'�xX���e��<<J�X����i�E'\Oz{0�w�Up�}^=��g.�-h���%w��<���s�c��/P�"���U�z3(�� B�#������+xF{�p�1�g'`�zz"=�_z�_˥��X��=~i�h�[�W[���np�Oڏ�Ϙy��繳�l����#+鹜4ey��g�&���T���C��]8��|����#.�g���702K���^B�(�J#��O�:��U���@b��
��d�R��hw�����{qYZ.�{ލ�.�Ȓ�_����,GC�I��\<�Py��mK���z�<���8�3���>{��_:&]��Q��J�6�y� �K`k�rԬ��z���#U��z�9P+r��J3�*Vd*�(n��7�l���3��V�/��!qa�U�#/`5�{]%Ԗ�/+a� ʶ��a����{�lkc�Z�Y�T�r�aq:+f^{/kmml�)�=E��������|j!�(����e�0�b�U/w3�fi�.$���j>R�m��p�N�1��ѱo��-�:�Hy⭑������*��&H��Ӌ�)��)V+͎�h�&��PZ���L�n5�K��j,���8_ΝC�%�*ג�޾Z�U~Շ��<!�kӄ���/2:Fx�õ���o������n}M<r�i��$��)�q����J�(��W���2 �5��&|끎-b�:�F�!Q�	��>&����g����}8l]��黭P�5FXm��Ih٩����"e����T���#˙���#+�?S���J��U~j��G����gx���Z9�H�Y�30�p:�T�����T������=R�Fk�ٱK�I���T����F�4�k����:��L�'dE��B�'��\���!n��w�?p֏ �9��Fږ7��w����w"��zf�~�=kבQC^J����C�E9�)��\��~x��W�1^�]�✮>[	_���}2�l�0���\-4ɨ��Qy�޸�c\�?��p�+R���k^ĺ�Y�j�����ĺ����p������<�;gD�V;��X�=�=f4XG�Ã.Õ"m֊(�����<�'HϐG�]��4��w�dJN��|C��(��<(̡���蕌b��Il�rr&��\��]Зܳq�l�1!�U�ѡ����l2��t���Ǹ5Ӛ�F�[��A���骼ӷ[_`ц�s��wX�jT�r��{jPr�5x�2���f��BsK�l�^+k����v8�.D���n��+�|=|,*|�lcv�xM0ki�5yw�\絛j'>lN)�v�@�)-��*��er�׵d�z�1���Yo{ �V-*|��4�J�JsYD�rV��WʮƑ(8�b=�&��GW>۹YS˨��C'e���Y��]��c!0^Ƒ��e��������7�7�;ݸUG�H��,u�u�w��03-%68j��l�*J��ƅ3bR͖L�27yⅹu���~%��Bpx��a�:���sk*�Wͱ���t޾�v)�	ni1Z�2��Ul�r����/]ʹc�������[��]���C1Z�竵%U�];*4O��ofC�}"�׍ܭ�W��	�n��6�/��Vp�§k�֓Q#Z{�7R���
c5^�K Z�"(�Ӝ9X��GO짽)OArl�6~�oD�^
��J�;˩�v���W�j���f�߇.��X��abm��L�@��,�ᵤ���r!3�Q�P�����G��]����Ɔ�X��\���u1���HN�f�N�8�J�6X��c��ӻ�X�&�ڗn]�v"���8���p`�E���ވ�Gd�Z*�vG�;Ց��,PWX;�z�k{�>q_,��}L��A�="'�sQTj석���!F˕�M�
���	d�MV{z�]N��kS�wy��պc�*p������	����L�����@���.Q�P_ʮ���G�vs�%���b�.��>��E��j���[Z�ݗ`%Ki��h�0r�P�����Bn؀b�YE��R������YW�$����+�MX�����Y�_�KV�/����[W�-��ث����SʹZ��č^��>P<_gmI�J��y8,�a��a�Nϲ�p�P���<3`"s�	9�\�p�*9]�i 
�Nb���t��8
�G�@��d�k��	������(�KU��%ͥy��LB�+��%c��y�A�(!��hX�����=n�d����B�u���z���Ȉ�cc�o���D����֣#'���d�,��جgA�R�P���W����i:��;5��'3����-�+��xb'�Bf������rc���	)�:΄_8�O�éǻ�)�hF*���5��=d4k�ws�0Vr�6����w%��j�}��l8��%y85\�&.6ln���tYU��+�B�"�¨|�{t���昉.�h���;����$�t���wt]wm�;�K�uܷ;�9\s�����ۜ�\�A�'s�f��7.R�*.N�s
Dww$�뮹�A\�����K�\�ɺ�\�d�l��uӥ�c��5˙sW9���������w;�Qss��wv�.\�']���]�K���sgw.��N�\���;s�B3��r�s�鋗wk�v���Qu�9t��;����v\�w\nQ�]�˗5˝71sS��v���(�;�.]�Fv��Ӯ���ۘwN��]u����Rwuq��]".��t�%.q�9�vn�(�wS�]�Ÿ��wwq�.mʎ�.��vwt�����s�\�.��.'9s�;�n�1*�$�E� Pnm�p�M^N}+��pu�s�`������J2�Uϻ��)�\�ޑ�,�!�Q���a$xSlT�A�;#�׿�� ͝ڎ���T��t�ڥ��ӯL�&�H�򿷪AЭC�F8i�y~�襀��}�9'/�<����?:��%x�*6e��^Wȗ4�|Ou3b@1R����}�� y�~��w�z��	�u߈���\Ud��G�l/+�ٖ��v����ݙ�<l�ϰ��@���{�g����:�b���MŖO���r �=��WMZ3n|�7:5-���c�|(�C*�<���!����=��������H�m��G�;%gXݤ���;���T�X�����T�3p�'@z�u�8�Y�g���C�9<�.J&��}~�^W���m\�Q/�4�C�/�t���>g�u�˗�'B}O�E���1��=*3v=�/zL��.�����	�9�4O��#Z�`O���1Ųֺ���;򸫟z�9��m�imv͝�]��/�#���/�MW�ә��"�}DL�\�:_��ΣkT�r>�Tb��#�����F�|�Ǉ���0�Y:۠��ʌ��҇uF�/)���/x�O���MqF�r��z��!���տ]پr7/�ۦX�< �EC��}�1������;�C����+ �JV���Ƕ��<yw],N�WSR�9B�H���P}ܣń0v��W)��W�v�S�Bd:�ަ0�����9����r�b�ķ�J2���t[O�Yd����)ۨ��rz��/\@������.z���ޭ���?IKY��ƹ�t��a� ߪ�)�K%�.#��C"9Ԩ><Nv5	�n�S�@߽X�,����+�;��8�����﷞Ӌ��Hоsʃt�4��Q�}�d��T�ộ�p𘖠ٲy���4q\:�0�=�������YP���9�����`p��$�d^3���
r�/���Y��F,�V�^}>��t�g�������r|�}=�˫�Pf}�����Dw��ߦ����f��8��q���:��rr(U�����P'+̈gݧ=vй�H�䝇�v���8���5����_e\Δ9�þ�X�d�4tz�@8��*W$(���u �i�X��M��z��+!�!�q�i�V��>%!�N�՘�������k�2h��/�E���7���"F��l����xy�z��u�sEu?0m�.fK����#}>$�CG>�*��F|��ˁ,�uP�q��6�^^:�w��:�F��
.n��^�دS�^��q�>��|pX����v�ک�}z�۝��w
�PNǄme��ƍ���h���h\�E%���2�^��b���Y���+'��JG�Kt�I�Nm3qM�-c9y|����]-늙��ݩR�(�4N�oY��Z�D��!���Pֆ���A�d���z��`L@�w2��d,��n!۫q�߸⻍��S'�4�&���z}�r�j�}�gv��( yQ�������c]Nx�����"���k���w}��a�u�9�FPx�,iq�K+���<[�!{w}U��}�ۧ���L�x��Y��^��	������q���I���Zh9r�G������ī�g�z�<�ʡM��[F�#���gW�޵����9�-���w���E;t��y+�^NfCw�1.�,pTg�|vH�����)h��~/Ɋ��m_�߽��lˈ�}�q�Ysu>ɵn�0�!�-�E:�(L �x�ǖK��v���,�)|o������O��5�t\TȹPl������J?�F����bF�`��=8ԭ:.+__��u>)��U�����{Et�K8y�u^"�6%�O��n��ixU�Y>G{d�r/�:mQQ2n��b��5]d�ˎ��U���{C�9�k]��P�CdTWUʳXx��(y�s��p��.nEJɐ�MJ����b[�nc����l���pw~��ކ(���z���j�bNhぎ���ϟ31V�(u�nd�nnVܣlf}��N� ������Y��;�p}+D�"vU��R$"ԢVƮ�n�9Ml2ӺVv�pV��nq�.r^z�"$e�S�].��mc>��V7�G{����K�H|X~�Mj�s4{!?�`2�g�x&�p�2�'�i�+�MY*Srq�F.����+�[3�<���U�a:���b.�x�FPIك�zĹ��\!�I�솙;ܹ�Ҷ�q���`_p�(P�Hqh߾v�7���|dX����f���	A�i~�W/�'7�Vv���+�I9�u~w�&�O��%�a�[;�:��Ui��v��&��>E���T�L�ق�L=~���u�K�\R��ޚ2�hO���ÆG��1��Oo�<�V��$���d�H+�7�<�_�_��S���_S�3�D�|\��纤'N��LR|�"�d�>�s|�z��t�Q,�e����Y)r�~�(p���4uy�̎��5��Bh&�~�\�mla>�զ.61,�E^u�Џ83��;>� 54\�1�p1ţ�B:Fx�o�FW��qd֖͉̍���fz��v1�
ē���FQ$�"JG�zH���B��T��Ћ�q�B�yb�~����Fb( ^�q��+dH�o�|t��l�+�6_v��M��4���2���dU���ر����X�Gt��un���,�aɅ����8q���<�u��֊cwM���9��;=����̷��<�sAb�*Fr �L�ӕ6�3�А^ |�5�W�m�g�L�/\����o��i�n����R��2�|1[�-�J�W������y���$jvQ3���š�_BvD��W����T����9Y:����)��y�����d'���iP�B���*+^J�#S'ޟ_�5U���q��ȜX���.�	���'���N6(nVS��=7�G��ڸ\o����O��e�U�j���*��(����?2C�7/��M��.f�+������*�'%N^�MeC�YS�����JѺ�9G��Z��s:k�+̟'�h�?P~�s�ن���]��ќ
O4�,O�x��>���:�j�ȵ�:v�e����'�toƝ)�K�"����]c�����z}]�ny���ec�q��ю�;*t�Yd�Y�2��,2�t��Cڪ////У|�^V}�Ty��Qׅ˃��E����S�~�Ui���#A�y�)`��N�Օ\�������|eV���F�뺉V�e�^�`^�>��{&;h7]M�kc�Fc�R�<V�P�"���n)w�,�-�أ�6�]Yk2�w�*��=J��c3ACR1rX4����u\�Ma�r����;�n�T������33��Q���r�̏i!�~�p��sԴe��]5tƺ���IlΙW�6��۬Bɳk��Т��>GĕFc�IJ���t�g�u��OhM'����_-���Gi�bP'�HH޳��EL�Ƣ��3���'�
@I�7^8�Z�V5w�qW>��{�}~�+����Iw�73�����\{}r7�Y�s �JETO���[��t�7a��Kw��A��}�7[3�'QL'�|E��k��kp��+��YQ#�<g҇p�b�>~S�Sn��sܻ��Q�����ø�򹌯?S��i��6K8��d`���
G��v�!�G2ֵ�zO��zw�MI��!��O�����W����Q��o�S��K�N#]�ƆDH�t��9�8�Y���ͨL&��Gq��"Wl�q>;V7hv���ßM#B��G*ӈ��=��LN ��{7O�B�4)��[� ��e__��a����Vy��)3�u5˪o�h��[^�{���OM��ZJQ���ꘜ���c��f���������7.2��{I�cus,{7��>�YWU��o��Q�R�5��xE���=��_�Vq��g�>;;q3���l�wS�tk�-���;��H��_ۨң,�w`��2n�۬5qq��ΐ�OK[�A�J�3���2�X*0sY&�^�ڶ;�8�������/��$|o�����W�j��S[nF��4��Mg
�ڗ{���o���:e9aT�"��!�ֻw�~�߶]�~���t�>�8����ߵ�x�ʹZo�Y;�û�꒼�޳c�ϟc�U�*}�hz)M#pk�,�L
��xȖ�^Ǯ��J��'��V�������5�9ݙ�^��eh�I�;�E�ezC�>��� �G�
�d\-���߫��=v���o���~�;��D�n$vf���rʐ�.x�ƢO��*��>Gc�\	f�;�ץ��a�,�EƼ���{��
۟}K�òr�+�T����2��UIn|;�Yu,���X��9��H*��7�����kO��>/�o�3��W��_`�JTe��χKe��)�Zj�#/����V�f����bO�v.}���Hү����S0��f�A*��Rϐ%�d�^��-K��[RG��_9��G��ףb�o���j��n��M|��OO�'~fK5�&������r�5ܯ%�.| 7�>&'�]]Fx��:�w�H�i����"}��:7�z�
�4u��^�t�*����L���䘃�Q��ˣt���ʡ��&*6�W�7�z�>�1��~.jm��b�༔�3Nk�%>\/-�5���T�����Q}8˿Vq�'��sҚ��ʉ+�+')���+4��@ˇ�{/(��V�4�C�WO('�vi�۾�Ζ���g�v�;�ض6(��A���q�L#�����,��"2K�J���+-0ïd6��� OnT���+�ցN�I��,� ��Tਗբ���^=g9K�q��q��� ���������'����Y(�nb5��3��i#��6�B���W��P����N����Ǚ��j��/}YCl>u^#9��版Z�ܜ^f��}"-�FNB���3�]�;מ���C�O������U����~�y�cZ�~���sqC]�N������ޞ��]�iU,����!w�u���3��9�tDH�~�K��7:�_��f�׳�>C�_{J���X�1>���}�	̠Pvd���Ν�5/Ĭ�L��#�T���;��Ҝ�E�w���*2��~~�\\�b�|�o�S�z���(m̼4g���G~��ljLGV,�q&���#1�[���e=����P|zĿPͰ�z���D�%A<}S>SND���y����J������E$�<����4�K/��>���yd�(u�Gbܐz��'�|�f,�Ab�9������~v=
�����,O9�U�����5�|�O����[0�G�%�K[�~�u�ٻ.e�ڔ�Q�� �XG+����ϩ��g�}v>����u�{6\I�t�>WV�p��$�b ��<�Q����˙w���7�M&Ј�Ly�Z��l���Ԡ��Z�؉�MV̓+|TH�f�X��c\���m�|?K��&$.֯Τ&���Ƅ��E��/��\�P'а�OH�[��K��A�U��Tp�Y�ǌ}h�-Γ|�_��g���I�_��W/�[[JQA��N�w[#*�ˑjg��SH�<��H����lt�}�F�p�
�O����~�8�p�J×�	Q2�H��=Y�u�ղ��{�>2�����s�D�*h��
_�zEދp�H�#�5��|.x$�����-��K6K.�ȉ��)zj ����:�{ƅxU"�1륝�n��x���o���s�H��+�1@>�E昍w�F	�S���'E��/[�=X����ʬ�"L���k���T��}��5Ua��U#��C�6�>zׯ"��ג�����ף2*�]���F��d�q�{�a�>��_	�z_��q�ە���L����]=����;�V����*�\�+�QOA�=
�e����7Ǝd��7/ƥ.�p�ys47+�ŀ�e�#o{"ڡ�9�!�u'����/b��Z7CWAÕ��0�G*KNKģ���t�m����/a�ߧ�G���ŰRB�Qp��g{����dp61�#�G6j���ޭC7/J3&e�siYT�A��,�*!�1����V�@8qj��	��|�aL.,S��Y}Q�We|!��t�R���V����\�ܒ�1��z<�-gs���γ�"i,������Y�O��͎�ח=+1f�%�WVũ�9���>�m���9^�x��j�yͣ��:o����sM�I�P\;:�:�ۆ�Z��I�|�P�w��G^.vC]��:é�?X*��ụ�sS�(?s[ fTη�X�X�"N{�3�.xeL�����Ie�XϽz3簟��Lv���Cӹ}��>T-�{��&�
���<j<x��� yL>��=~���r�D���<6"�o��g���{ޞR�@q�|�ǳ#=��`�*�H�k�,n|ql��ƣ�;� CG�9��wޔ��Qc�[;�9�����r7�Y��25�G�E�u�����;R��;���U���<)i�Q��R
��]�Xj��� Z�%�!^��TH�5
���uzt������m{�oR����r�w�s�iì~�^~�~���q�׍F��n�j�:��F�ǫO
~��ܽ�¤ǳ���D��;%Y�}�>VC��֕2^D3,�Q��[m�[o���խ���ڵ����mZ�v�ڵ����ڵ����ڵ���km���j����m�խ����j����m�km���ڵ����ڵ��m��m��mZ�~V�j���v�j�����j���v�j�����j�����j���-�խ���mZ��b��L��#���� � ���fO� đ=��@ @�   �P   (P  �    �(  @� � ($  �,�gv�V̭jSJZe*̓]nɛ3j
�Ͷ��յ���6V�E[2Q��i"@leUZ6�`֮��Fٚ��u�j����l�ՖɑCӹm���lKY�i��f�ɄҲ�c%�b��ԦY���m1Vm�S�Y��d��T-6���cl��5RmZ�Fm�TֵS[-��>;vY���.�vx  t��A������vOx�v��{�s���PuְM�����֛��V�(�w�={^��w����-�;��xz�t]�-�t��n�<c���P�AU
'�aim�m�kf7�   ���E�tv��;���#����kC� �=V(�  Q|����:::4�>��E@}z/}�;x�� �ou�� (�(� ��G�:4h ����*U��;6��P�Lko    �}ƍG`��]�@z�nӊ裪絵 �ӳ{��� �U[z=t��۴
H�w����j�{G����y@f��u�ʴ����mF���G�   ;>��6�Υ��ӣ��ڞ�x��L��{��l��0V�R��WPz]�U^��ozݩ�ծK�ӱ��n.�=�t��+[����f�6�ʉkR��j�m��  =𯮥���[��oIv������Ur����k��t�zע����:G�[=Η�Վ����#ݷ�Mu�w�u�;N�8�y��={M[���{��ޕ��m۷vݽ��k"m��.��Ҳ��o�  ���I�T�����hMkwWw���۫g-/U�靰��M�e6ԭ{���ηS.�x{��ݱT�u���^��������ݴg�޽F�]�{z�k6[�á�-dB�h�  j������t��I��me���֝Y����Κ��k�\�u^�z륷�]]��GYy��]we�R���εz����ޱ�]z��\��jm�n��o*��Wv�))�ST��  ��� d㩻���׻]��t���T�黼�^{s��]ku�w]�vݰ6u�3m[S۽��v;5Q����i{S���z��ҝ:wn���Sm�^���زm�e���l�6h�_  ۯ�v��JU+��]Ye����{���+n��v�ʮz��<�S�ٮ�e���A���=�^6�cv��v=溶]۽��{���{uz�ym^ڞƬ�\Խ;�uK��Cmi%���ՙ�ش�G�  w�>�wt��U�l4V��w��n�it�����F+�mMvyt^5��]T�հ]۱�����޴��v<xz�n������zސ�.��w�.�ݮ����0�R�  �)�)J�hh24 �~JR�  )�A�T��� � 5J*�(� �iJy0��T1�z!�??���Կ��IK��3�ޭ���QSfp��:�f?o9��}u�o����H@�w?�BH@�bB		���$��	!I��ID$ ߿�ǿ������?_��LR������*��x��)�*��/�x��{{��6���=�N�O{$Y�d�&�;ٻ�t�$�h�D}�6�Ő�@�莭țMg'І����٣CKTo<�I'�t;5�j���7�Y�9�����X��e�`[B��ŵ�k;y����0X6f�1��-A�k*t<L�`�v��`��g�7���e0��S}�`ٵ�+��9�f�Z��4��Sov��,�wi�ѹϘ�&.<��<�O�{Ն�s��Cx�랴Jci�Wb��݂s0��Ƶ��E���4�7t�srGi��[��M�����v�6vի&�us�j%3nNc���U��y�A^�V���7lH>��L;4�����MH�ğp����5œ��k���l�T��ذ�������\�7����Hz�%G�]������'S�����齳	�嫡�08�W�j���8�}jަQ�'Dx�Obv��l1S���uiX汧������]�d�-�S���r$�
�d�O��>I�m	W�cߤ��lu�j��x�N#n��=�/%�~��LYm6���I�b#Jl�j�3w�5d@:	X m�K����M�K���G�4�t�e9K�_i�˪ni囒֡ķ$�]��GT�m��>n�)�!��!�'
���űît�����G�CހI�S�w��2�4h�q���V��|��1q�֙�;��Ǘ��ޔ%�.O���;�j�%�3�C�$ɼ00���9�[ugi��[L�J��gm�5v6;%���1V{��q�n�����Օ�"�n�M��>	F��7bmɸ3��l�F��ۭn��N��1��F�Vw=V2�h((%�D=�(��['�w:b�X��Θ�@�H�1���4l/`�����w.梫��\l�y]��u�=��lnvC5�L���ܛ�Q���F1ϙA6p,b���=�0!��\�]�܆�ƒ/:�����M/�s/;�'���F����q'��q��,d�r�b�[� ʯ(�v�_����FwWxs�*���&�5m�شf�npt%��4<W-ѭnN�pi�A�� z�R�o$2�vi����0&ov#���U�MIood���qf�զ��OFu�W�>�s'�LT��o	 ���q��:�Dc�V���"�J�I%�rҎ�w�/rf��{�|r�s:R�1mٮ����O������t8ĝ�]|�n�Y�7`w��;k��st�oE��.�n���u8V��4��0@�#�e'��^�񻍭��]dc5;'JvcL������R����y�5r=�p�}�˺�
�l�H��p�w��`�te�`wE�d��J,]o+v���w4�,�'=����x�oao�7n
��l@�u>��Y<�Y#͵h LwV���ٽYJX5\�M��,��N�h�����R�R�.��;oo+�zvj��N;j��3���t���K(�}\�&�(��.ݜ���N :C�J&�����pZgbq62�ƍ��S�s��J��7~�uS��g!Y����N�B�q+Zyc�)��mq��n�N�2��wYv���0���Ctoj��n,�Q�n�.,��s����Я�;���R���ذ��#۱�O��s7��ٰ�k���x �.��nHй�8�rx��*�L�@�p�i.�wa:��8e������y��g+������8sd�iшf��إ�g�ǫ/8�
����#U.j����@B����u��B�����{�N]$d�f�� xS�p�ݽ��V!ږ��^���x�UNOtc���9U-��B91�,	{�p���Rf+�뤣z�}��s�����sV���Kg�o�Uu�%]�B���A��4]Q�CZ6���.r�� d2j;w� ��ݛ�[�|;w�G�Y�(kCɶ�KC7M���'���Y�W}�9yأ�I�ȵ��ȋo|�M�?�0��b�K�1Y���mia����gw=v}^soF.q�Ȏ��T�&��1�TlS'5�����8 \8I$wge](�&�>#vh��4���]���9�ђ���;&�c_��Swx�펍�sXks���q���7~��zX�4��C�][rv�\��3��ģ���57{Gv;:����j솓w�pbw稍Y�Tu2��Wz���f�4���laيf�鹺tAy�mݹZ8C�y��-�^{��s��p	�A�٦A�29����Hfl4��8l��	:(����y�..H*qRq׺{��~1�.q&�\,:9���xFp�r�xm�8	�;����-x�ك�#d2u|
�Z�bJ���qu[�o�4Ht���M��_E*��ޤ�����盒.�d��N�;Oμ�����
�XY��Ӧ3�E�!����L��p�4@�w�Ѹ�7��K3���`*�Nܵ���ڤu�	���=�A;4"��EC}�T�eN�:G`�a���}��1�܍����n���l�L_PX�^�Pz�^ ���v��z��RJ՗�@�;��J�F�t�,��o9�q�����rm�N��o)�3�xж�X9�w;���-�2�k�\z�D'��]О$^����aȫ6K�uy�V��Itwq�в���k�	��Q�+�V�	�n�<�{�Ylӆh��'КVD��d�7&�6���1<���J��%�G~�φ�M�۲
� Z4�>�N�inv���,'ۍ����{�e�S���k������x�1��j2�F#̼��˝!�h�Ňf#`���8���Ս��� ^�`=�L=�z�ﲵ�j0���q�jU%���ae��q���<��J�۸ 9K<�f��H�{~��l��<ZaBֵ�Ξ�5�нx:���	kƴ�,�E��dI.��u(Vn�fnwk�(f����4�n�%��p�Rǝx�3�]	��9�6#�^���^9�=�2A"��Yq�r\���
�\����j8�x��W�sv�ۼC��O˵vu���
[;F .5�#�����m0nA� %f�
�����E�sL�4n�F���B�	ú�AaR��&���161���An�ގ���1�Y�bɝpq/��C]P��_N����Yˏa��͘��G1M9��n#μ�Y�JX��,�x��L�Źƃ:w
���ܞ�t����\7�m01��Ǹ�n���� �����e���>�
~��"�I�߲���u�)C�ۅ��"�OE�`}`�3��Z���!�����\��Jy���ɽ�ܸ.18L�L�6�;�/h��1��b����Q]�'j�x[���S��qS�(����DU��X�W����!��Z"�&��+5����035c�_Jׁ��F.{�ohJ��=���5��'�0I�sOH����y�tM���!��Gϣ
e����V�W��!���rX�j�õ��@�+-���ٴWv<V�ac����Nӳ�ԻUM,�� �>Օ�7N	�-�ۊ��Њ��!v�8]�VL��2��9MS��ߖ�.)�b	̑��<�6Us��wS/^4i�3k�i���[ml�Z��@��9$~2ǗE��}17sIMu{�!�&���YF9�Q8����w,;J:��t��D{ĆN���ݽ��Y�\T�+�=Wd�t��@\{��I��|�ɥ����[��ŋrcx^��hp���)�E�P#J��Q���z=�1�'=��ǆmv,�w5s�弗5�ov��阳lܙ����Oh�Z*j��_BGv��wI�����VF�����Q�̌��&��u5�lfdX�G�r����`��]�����%Ӥ��H#_05�f#�ZQƮ��(V����y�$N�y��d��Zy�h/,�.{gL�z���BV��Y�u$�{՝��U{KYϱp�9Ю�u�������S�Z���u��omጐ���7���[�G]��E1=�N�W:7z)�a2ρ׺�҆8 ��]��t�����gL���L�OA�UNw������OQ;���0���30�^@��5����ns�<&��4�b ����Hu=�w��w��^�Vj�' 9϶d� r1ъ�Jon���\��VH�T�a���T�6�r�,$�)^J����(�d�6v�"Y�],Qe��������N�Bt-]Fr;r�-�ߦ�]�6�;"��i�Y) ���Þ�wΛ�+iEp
����n!�{5�ٺd�XOl�7������=�
�d��zs���v�vɑj�h8ZWx��tpl#�jTa��G�1HXn`�ť������I�+I��X,�Y�dRb��'i�ʶ���z���KŜe��I���p�0%�3Mk��r��=���5I�ik���t�a�@mӀ�m�;Q�ִ��&�=k��|��2�r_�"E�&��|�̻�N��y���T�Uܭ�Y3�8���z�pn$��.�踘���m�����_e6�>�t����ހ�%�;�n K�S;�QN�3�Y��0���L쁡z�}�Mo����!�|EV	=OOk����+t����=.4�S��D���l�N���7�ݭ�hh����U���~X�\�(�GB����N.�������z�Q��it#��{��t9�n������W�4���#cwj���h2�v2s�d	���ْ.t����g(S�v�.t����v[�rjm�/��p�EWZ���y�לt7��ݼuY�"��F�]�X\w��x� �v=��V�&��췔*�q�:�Q8u}�V��L�8��[�=�6sjg�и��{r��,a�#���c��Wp9�6p�;��m�Pf��z![ f�fJǚ)ބ'[Y���%���Y��9M�L�`�,��r���\�J�a�pィ�fۛŗ�p�Y��f(B*��ti�C��;Ƿ6���|�ٓ2G �4n�*�e��ո�$nMÇ��ܠ/���n��ތٜ��cB,����%��yڸ���gu�x�5n�1�z�Z��a�a΋��d�^�v۱�X�x�e�TB�ZQZ�8��E�ZTk7ٽΙ{.�ua�w�˚M[�a����Y11 �&_i%��j@Q�ȹ𠝏��[,�t�P�t�.r�ʳ����J������.�٭T]�;���2�%�[���)4$�m!j��&ό��ƕ˓�a�Q�{_RW�X>M}��Qz�H2�֜�t��fn��H��f��{z��%�v'tl���4Svoȼ�����M#6�ۭ�mt#l�7��]���6�ZN��Gφn�2��{fs��W'�I�w�G�x��$5��c׃�֩gó�t76���Vh`�n��ϖ������v�dᕜՇ�Wz�^�n�^ ���f��j�r�˭ձN�U�!b��=�eҏ�����V[o	��ۜ fob����������c �U˵JY9��4�X�:	tF�5��D!n�o!G^��;�B���Gf�i� ���Y-�0�xY�^l�݊oa�rG��m� ��l���D����]�vE��5r�7�W.j��1��{[8EO*�� =�g�>����h��P�K%3f̜)�P�J�qМ��ɫP�������"d�m�3b�Բk��
�{�d经.��]��5���ӽz3{f�����p}�F��h�>�!9�n�:�����82.n����I���V��xa�M�oWt�sf��<5*.�F�D�Q�Y�bޭL�Q;��p`ڡ��k\gj�(����L�xv3t����0�\��>���jܮ��a��=;���/U���|��7x	aַO=��u���M�βb�!���\&�їr�l�_q���Wh�����Úw���`yc��Lo��:�����aul�Z�5������b� t�:���ޛ��Χ�@�YR���+[m�����[�)�x��ϖPCUc%7�
�k�M[w�U�kq�s5�F��N�٫7�T�EoC��ïb��	ɺ�&^D������)����d�Dw�]�	��8��n�IL:�&,����f�!��qq�od�7��W�\Ni}�G��r�����k��k�w&�=b�mv��hx���kY��nwf�JI{ܫZ5#�E'; �5j�Fs*��͝e�	Qɐmc���:G��1s\�v�5b�`=�������vܩ�W��cHff�9�j��V���ŕ��߈:u`� ��:f�x��� T���VNa��~��p�s�^�Ǟ]�L�=��D��v��aW��+F�97{��f�+4�k����8̈��ú�O,Hs��C�a�nW��5[چ̫�cR��M�{���4��5$3tp�t�雂tO�y�/����syT�wp������Bq�viz��-��+�{���]����K3�r·5��nS�gx��p��qop*���ʟq��ݪ���#�T�)C�9�=:WL{qF�U�o�Swѫt�3��n1c��V����6�	�eLtU�3�f�N�^�\w��oPR�Wk�V)B�;J�H�ykvĩ�Vf���l�S ��}��$U���DF��6ԥ�a��͵PI��I�\>��Qi��6��q���h����]=����1�_;�#�[�֊O�:	[P_R���m䗫+�! �Se���D�gs�n�.���E�7y��c�[��A|�7�þ��P�,�p��a�o%al��>�GoLUh۝ΚPAY������5��'ǔWw3x:>�p�G�pٕ�i�t���]E4��+Rr��c�2�͊g.g�����W��3���l�a-9`X2�w)Q�����8b�
���g74шxUo=��&����u���Ïf�΃�Y����au�N1��=xM�縅�Tg��U�R���:�0[k����_'Z�=EΫ݂��\�;�x��S&V��}�l�c׎�y�V�sپ}��Nm|����n��[HnXì�n�A3R"�S6��,w<�]8������s�C|��Ҡ)ʔ/f�6��q�pO/co+/��	"lY��r��ݦ�}j�qJ=][w��rzuּ2 8���d"���t�+T��+���5A���c>]����{�W�@�(j�P��#��:�Ȅ0q���ʙ���d�"�b4��A7�G�{�qc�EtC��@u����[F�1�P�.����f.[��b!��^b�]݂�������k�C� �'�u�0�S���&� V�/l�5yz{�	5v�����M��*Ӓ��l�͋�pvJ�./as{smn<M�Bq��o����jmG�����"�,U�KN�$ޜ١�Ԗl23�a��Է�t�[ :��+4����U��o�l�E�:3N���8W�@{����0�q�o����bN���P�A9,Χ�ڙlJ�vq�ƪʰ���R�O%2�rF�L�{�-w��=���w�dg!o]��?k���`{�RR�N띌�x�0h�vL���Ȩ!������}P�j���pVbŚ��87*~��*L��V�jޡ�qXGh��	bmN��-�<߻�_�$KZk3<ľЁ"�lN	ҜV�0;N����k;m>B�0Vws\��!�ޫ�i�暎n�s�V�8;�J��r�x:L�I!{/i�ܼQ�5�K�s������Z�.���u!\&�����2u�Q��B�U96Sغ�)*�3t��)��*3dHjJ���t&��[Ǆ�+Y�f��|��W��Fk]q&���f��/���Ct��o�IȬo\t>���+ih�1jgS	�\�n�)��}`�H~0?&n�t�k���Vk�c�]�Xm�'�����#��M0o��"�S��Uu��ꢰ�|dR��L"�.��:iԕdt��y9��ë��^i��9����+gH�����\��f&l���D��3aٳ��z;�}0ڨz��7h��.tn�����׾�pq=��O����3y�-�I�x�*�m�$�@u���ݷ&L��#��w�����E<�E3U���!�z�^�FQ*�L�V��Z%�N�q���MҸ�Fwy�K�=tSy�}}D��bԎ�|5uv�i\�ݳ���o���ʓO0�s�S���yع^���X;������|�b�%�b��Lk�k��ur��u�����f� d�3ָ:F�+�2�y!���NShθ���b��ObYv���굽�V&�c��BB�g8�b~�N�k���j�}*����Z�t����%�����ź4�I?��x�F�:��Ed|��f���n�T�z�ܣ��[���Q��Xٻ�:{�����a����Xt\�S{;,�#c�Ʃ���M���
&vu����p8�&���(/�o6�l�8��9^ g8m��x�k��E�ߋ�g)K��oOd��宗��^��H��u#y��0g]oB��N�ח�����.>���y��� 1w�L��{N�W24�c���M7�5ٳx�kKcZ�X����u��ѡ�3}��]{-m�P��%;+n"p�i�jau�޳U���_J�܋y	�ӆ�ך����*=L?�w��U��eǍuY�eaJ�hWs����cq+��/��.��o�G���b9j�$���$�HѮ�h��@�\��#�@v�����mG]q<�Լ.@�������^Њ�����J۠j:��C�o�, �2��7�8Q\�X�{����:q�"���������:�q�4��y�Z��A��M�vzHe��Gsne��.�оG�aFfҚ�މ��	Gg(����㌲�[�Dd^،^�rw�O}��,��Q]촮�a�f�j�^*�e��X/Xw���.�)sDҒ�f'ٜ�Y,���]K S�r�&Ce4�����Ԅ�����������6P],��vL�v�,F����t�r	++]uJ{X��3��[ $��sỳ[���{svn��t����>��T��g (�<�!�o��NQZ�*J��ʂ)�J}�S�SG[����;P���o�Ր)��(����%]�c�dl�)�.ٹR���`���m��kT�0�Kٮ�5��}{����y������o_ʟ�-[�C*�r�w��\�r{4 �!o��w��f?$4r�c{ױ�\����/�ʢ<��M�!���ݚ}{�Y�$�,q�yV�"1h=������g#�S��c������gf�f�ɥvHA�;S�%X�:̇h�I��;X�NlSv�S�|�!�}�ԓ v�������Iܷ ά��,�dI�3ͮ�M`䢎r�Q�E��ko��]�]b�S)��s���hl�K� lK�[zm��y\�7O/7�����$�y56{����U�Xy�qp�Y[�G �)�/eY	�1!,��pd�/��1r�zh��koY|�e\�[�-��4�8J�t�zse�];�V*��QV��(���S+\mճ���C3�U��]]��-�|�"��R���0~�#Ʒ|-�n��Ŗ�s��&�����í�R�z��Z��Щ�B=R �W�h����=13�ӧ�)܆�<�2������\�ɪ�e�:Yk_T��c'hYS�E�U��MB�+/-�����%	.T�6��J�̅�ws�c�� �Ԡ���h��T{��Gxt�Rp�5��D��Eqὂ�\�yt�*����o<�_uOo�)ۗFZ���J�fĨ-�3h^�T�R�	�P�!5�c2 ��`��S�)v�ڧ��յ���o#���CO/p� \N,�'���'����ZK��w�a�0n��SwX���|w��x_(���F�s������g���zE7n<���9:��Y����&v��E��m�;y٢���O0��9c�C�D�����]Ĳ�kKSLO�t�����6t�..̤�t:��[s�x�J���	y$��ዲ�;v�J�7��J�?b�j�溂,kQ�x�՛�JT����㷅�$�2NW>2\��w$���̝���u}nf�}�r�F� ��S��
6��xCpw�3=4��ܦ��sఘܿw�'�N��}]�6����i��e���ՇR\�H���<�[��ؤ�ɇڷ�J���h��k��T]t�)w��B�l]Q��X=�Y{1��޷öN�ke?�,n�"�RYV:N��������S���E|!b�6�R��CY֨���%	���/S�Y��]���v���Oh*3/^�t#��'7{�����+-v�YB�Q�U�"	�t׽N�.vT�o���*�y��n��u�j�,�8u�D:��b�afά��[�k���q����Kj�O�V2.Cb2P�(�kj��P-W��}^�z�L˛����p��n>O�\'��w�	4!��Fb�n��%w��,\/#}�aG��@��&�Y�-��-�y֩̋�bTϰ�xݑZ�;yp�N�5�z��Խăzt@F�X)�a�/�\Q�P������N��;<��
�8]1����Z���bt�\ҵ���ޝ����\�9���.T�wG*��J������]l��WT�f���u��ٜ�~�*������`T���J c:��~��\г���X�u��erq��#�b��
Sѽ+��A�uuBM��/�	�v��8'Q�tĬ��/q�ұ��|�t��E���7;8�������%fN"�fu�ZV��%�|��c���	Lb�`��li���G3(ܭ�R/a\e��J�ƣSL^�՛x��^]�g�����ٜ���_�P�U�6��]�||D|U�h�����D�y��7<�Z�O<ߦN�2b���K9��f�C��;���9?iKU��j���0�vn�[�瀬��Y=v{����]����v1��xv�FJ��+��~��;dc+����d��{s���^�u���EQ�GT�{��ѩ�˫�*�g��l�`hI ���Bo��o��վ�)c�J�S �\M������P}�NO��]����1y�ѫm�p�co����#7�~����?yh������p�m�bG.�niW�ݍ��.ֺ�:�R���A��F`��b���yumյxXF��&�v����FI�B��`��M�+�c^���=�6�v����V;عO�[siA�mtV$��8��E�̢X	6��; m�ƟyL�"��k���hl�. �5|���e�=}�R�IIn��yn�5��t..�ҟK
e`���V�EY�Vҙ������w.T՝6�:(�sl+���6z:9���E��Rk�'$�9G�D6A�Ż�7��a��]+��o�]α�X���ij��ju��('��7;\ژw�0�:,oNDk�/s��G����b~�����I�V0m����f�D�ةҲ�a�X`K�U�NT�ъJ���]-���E���%,����פ��0��,�zQr�G;���b������J>MS����9�N��+&��-���y�����(�?�:�Y��E��c
˩y �w�xv���j�s�%���Qɖ�˕z�V�����mW+\R�#wݮ��&"dh1`{�(�m�S9C�����]�v��+g`u��*r�ט�}��ѭs����S] �O>-�S�cWG��n�͞�c�b��ؑ��&<Y�����hȟ	�-Ѩ1��������W�M�Mg}ZbNz��G��{�@��̲�?{uF��Y<΂8�oaG����0a!m*R\��k���w�:X��H�V�$�c�ڴ�"��ɳ.t���q�u�b��Y���|4��*��1��gi��Z+�vf�ն��hP:���x8���:o��_�;��a�@�ze����(�xz��p/n�[0��q����q�]=�e�ը8e�ݙQK��P 1HK�Ŭ�r�S�]��%k@�w'fI۴--�6L{�۰Q�>�d��S��29Ǉ�n�"���x��ھ�+�F7T�,臃���S�Z���
�v+0����������%��-���S���!�]��b�d�%��{2��N*���uc�5��,Bi���2���'�����{�znV�lgy�v+Yv��l��N���q�A��W��������q"�6�u��"���ZI��������Ÿ�2�4YY��!�*�>����dz�)���_ �0�zi\o"�W��#�H�	FV�2J�h_:�E4G(�{MNcSh��y&<�w ��o�X��T��+�셎s!�DkC��;��;�79�J�e�缮��N
e���������Z������؊��7�m����;.����;�i��M���������%8k>�l����u���6�b��m�]��\�:<1ǒ�Bh��f7�jc)�˞����AvP���6���Z�v9({7
��!]v�=�Du�0�ʼ��ʈ����9i��̕|g��Tә�C�qhb�6 q�<�/;�a�`�>��k+>���g�����s
v���V0�Qپ�_EDNE�m2)��t9�:�MG����n��9z����J\)�����ց�*��I���d'F�e��	oX������Mm|����6W�V�+��F��q�Y-7��P�Y���bMЧ)g�)���s��M7g�(��׊�ݼ!y�sͶ~�|u^9�j��$H9�͠�%�{znQR���N.��`��Kδ,�V��M,�/�6�rKP��b`��
ږ�Zne�sx�8���ՙxJ�{�ܹ|~�����l�F����s�i�\�ѵ��nvXvf#2���3[1wz�Aa���H}�#{K4�h�*P+�Ɏ�hP�n.����I�U�����Ԯ[br�mdȮ��;�J{�^=[Ŋ�/���vҫ������\�j�q�P��b�:���6p�+���l�r/�J�����oohQ�ؙ���z�Z�q8�tu��7=�����xjܻ劤P]P��(�>�b�C���c:����޴ּQ�ά�9oE�`�ɭL*��)7�u>��9 j�_w&��R��8a��V�e�űe .��^�\;H��)L��hv�};h�x+�`�m�2�*]�t�A��쭹�t�q�>�+o-�+��h�5�7���NぼkQ�h=�R�GnP��m:QB��Jj�4�%'wg[S1�(G֧��MR�quu\�-Zy-dcR�^[���6T]).�����c�V:�n�N�!�y[p�U8;A��m���wN����iM�\�.쨮�J�I�}����&�M�.��\_U����.�����/�/����m ��j���F�M��KE�ц.I�&��ƷϹ�BB!!�@�$�����/�~��܃��_�l.�u��k�u�11�&:�n�z���d�Q���p�ë�bv�(]�qlI�tz@��<�6q ݀�s��J�-�pT�A
����8��ΧO�v,ܠ7Es��[��\{/F�����)�7�Ƴ�x=ƽ�a�u"^"4UTN*T�7�/XN�Љ�[}�s��tK����"�%���ؼ�j���+ۓ�͙���ܽ�{�����r³��kK�g�O��^���0\�Q���LV{�(�W��qy����-�&8� �Q4���Z��f�jAt��W�D�����@��ɉ��rf�F��Þt���E�u���+*zR��Z�˻���.#�7<J������XfTa����zf�eЭͶ�r��$�����d+�6��������g7���������^���Gxep�H&3�n �E��g�����_@�so�*'��xGɍǅ�Bc�<t�pm��N�mu;䑌'۵�q"��Gu����Ů+1�ia5>�d��-L���`��Y�D=��R=���H�f�FZ\�0��i�R�s_&�hn��e��k�j�>�6��S�����zڽTRW�΂:O32v����5>K{�-b�Djg+iJ����XS��-�/5k)�닏����>�8�#1bnK�Ն�r�e�xN#9���m2/T���<`�w�Ss�s=&�rVM&�|͕B�Q��,K���&�m�?m�o�u�AP�p��fa(�Z�0�Ժ�6�� A{����/J�/�Sՠ���n���Bk���}EQSwzq�u$��{J�q�8[eSݡܓݒ�Xh�bGK��۹MR2�z�W'�`�]8��ѽϝH���]8��ܚ��OT���7�O�Ak�C^�d�k#��^�J����v��qo�f�Ks2�	�olD&���<���˓Y>s[Ii�o���S�7'H�����N��諦�kU�oa�������=
ᓮw��oh��/ ɂ��e�}�}�$�%MVBj� z��(T��K%����ժi��.	��V���H�!�d��.ݛ��h���t�_Z�}���_Y�'i�Y���o�k�Q��R�����QЍ���#�]ם������xbCw'����|�.�DYH6�:�ب�V��̂�ާ��M)*���,2���rm�\�eGE�8���S�*2�]��7
շ yvzq}yX�<�|�[{}HRK�(viS��+w+D��+6�����	�S܋A�hreZ�ͷ)\�Xz>���-��Af�˛3y�IYsE�k(f@�B���4��/J���f���Fe���\X�T�~��ʳ'C�
�k�	��;,WQ��t�"s����Wb�d�Lq��e��b�O U&��5j����n	�jv'W��J�"t4R�Һ�f�Ы$
��h|�l��9���)G�fH�Vy���4����{ƲJ�Z9�F����
�w��lQUW�{� .���f-��ם� ��w;�73���?>njb+�s��O4���I>J�ڜ��w/��H�f�p�RN�о��$cod�y���%�I�*��S������j��������Y�I�Vjw�����up�sj��X�	���e2�H�tT�N�:�ш;6�[Q7u��u7sw��[��� ^�=-S��X6��R�f魺��vJ@��W�Mje���q�홼�3cx��ۯ��ާ�k.&xY3'���)�[�����E��ӽs+�屃��}�-���m<��1�t3�S��#k/V��ɀ�Z��|�qK�yweٕ,a)�6,�o?pMt[�9�rdFkpt�W�N}>}��|`x<f�&��F*���F���Z����Й[D��۴_r!�w��8c��{�]� �_R��Ii�6�l�gIB4Z3']t
�fa���=1�j)��u���vü�N��i�k��fi"I]�R"�BwJ�����\w��9�������9�1$xd��'ě�;��t׍PWr�Y��˨b��:]�W���o�-�Y*D ��F:���7q��9͈n�n�Bw�3����Y���b���@Ou�S|���z��_hY�l򏄦1���|5�Jt��0e�%!�B(M*r�8�J's7)$6��q�3��aŞ�q��=��������~�Ơ]��P[�Yq�yr{����Aػ{�M�k��YS淡[f�F��7��a��_��̧�Xk��ev,t�
A�����r@�`t��9E���E/���(�ʺ���,db ��u�h���[�j^i��TK�-�*A�۱�t��]X:��.;�}��J��o��+��>�=*8o��D�������	d'��6b�Si֔�"�Y�t�Y����f�۳vi�|a��M]*�(��9���+���.�Ҏ�j�������v�U���k$�33YF|t���h]�8�`�5��d��,���zرJ��/j�ٜ׷��F̶������Rwnn�s������C+�K����/������Is��g�[g*q֒;E��J��Tjq�c�G��+q��'3�%�+u�M:�4�\*�!ڝ���ݻ����Y�Әm-\�oiJ�$}qN�E쩽�J����r�%q�Z8���WH����+7���;�z�
b��p鵵z����5j��U��o8�h�}v{K�v�e+VM��O�۱J//��{��b-�&��ͩ����4s�5K��3YsfÆSjҡ������������a�Ž2e0UB��	.o�:�ay;�s-퉼��/x�6��"jD�_X� B��&]2C"̳DIK!�ؾU���7���zO�Z=�8}���H�7���j��o5�<���M�2w3K#�rG�I��^L�n\��9,�'<_�M^�mj�4gŖ+]�Yos�`ܼqv���+J̭-�*X@�y��ajt���Z��8f�;6����u�f�\܂ ��7�63�R�NŽ%#��~u�E�5��G5�,�������0�{ y5�r(��rdS�.9�,�����v�^���qf��� ۅP�nom�Z��W{�m��8d�v�����]Xv_ͤ 7�Be��]	m�nDb�W�M�_o/�o����5�Ӽ�:L���ۅ��C��O��������u�Ğ20ry/p��L���qЌ^ń�����!�{�A��){iv/^�H��}�	y!]�Mk��`]\o6@���ձխ��P�k̕�E8�B17�$8��td���c+-�O��/��\$��1�o薁�m�����w+A��nSB6����ccM�].\�y4�<D���V�\��#�O���V'3p9�^��b���	.�%��� oV忶ź9�3q�qղ�TUNQ�:�7�p��4c83�9��Zۼ��b��d)z�}#���d�Sp-Gco '�ͣm�P��X{V�;p�h�����u_XJȚ�IQ��D]fn���9���}ې�r�ٹ��R�.�Pb�ɰ�G����>��ȹڔ
:g_K.�Z��/8L��Jg�1Goz�k�.)[�n"�IZ�������R�CJw]�'�d�n؜}O�Ú=aE'�,�S�u}��d̷ص�|�<0��N��[�0,�wy[������}H�\�k�N�l�;J˷(>gЕ��Q�����BW����נM=���G3yZY2�8�\l��gPVu�=PV'yR,��	���5�[tD� .�Ng1��>�3���P:�n;��y�n���o�S���ygh�]ێ�7�d=6FӽWx�"+��N�a��q��1}F^��M[���
'�>!�k����I<"�V�;�9��% �ܶ:6��䅞A]v�34"�N^4�onE6�����.,�%��?�� �X/5�\X�ɝĤ3U��'�n��ͱ;��]������B�n�c��֥vB%>岣�؟�'��C|"��E�M79�J`Cm��=��̇j��#���q�nwa����7��NTTe�\�bu�[���z>��~r2�ݠ��n�z�v������>�WJ��� M�����X�[wn���L7wKP!R�qa����1GE�����6ܲŝ���ޥ1�u�ژ�fV��xq��b�L��aʌ �ї���YTk;Q�K���*K�V]	����}��;���N���T-t��2��z��\��0e�����*ecF�fl��5��]��2���h4����J�����
�m�Z��C$X�*�~U�w�����U��3��Y3�FW�J�����o��5j�Wk��q��Ė1�YҺ}����a�R�����I�L_gfn2�S�w�ܚ�9�J��Q��=�J�(��x��X� g33}0ae�O{o�{e�v�W�˕aכ�e�p�(h�M G�QB����0�� *?;��<�X5���1Q�����:V^M:��9�@\`���j�*��f�*7�\�(>���X�S��� �.3q����ڣ���HO9��5�^�����z�{�c�˨�s%?��v�^VJ��w���V{K�';�qe�ݓM��&;�q�]{�R�Gx���ݖ�[#oL�^�vO�����['tS�|Ȣ<y� 6f�]c ��
A���)����=�f����ٹ�H�|d�%cl�G��1����7��D^�"��6�*�7m��:�$s;{�p@Mfە���!�6�o����� z�T��^��&�+ m7Q+�[x;Wu抓/y!�Lt�b����	�;~�(DT�\"v�����y#���Y��Y�>G��=,A�b*6�,0���&��������I�vk�] I��k����ȅ��A�gp<�ȧd_b(�#	R76̖C����i�fgw���\�ݽ�堉G0:�Ku3؝ca����G']Y�vެ��L��{����n<ծ�:�n�2���O����n���n_C	0���a%������[g9�e�ɓ(�T_!6��&yn�N,��ū-YݪX�X���Wpt�*@�AG{�\p��}"���������X�MB< ����sU�5ֲ�5N�� ��ܱ]>�OO4FP�$�M�Zc����[����S�~��Y�R\~-�־�����B�(��u�{�?���W�Y���qp׻)��
࢛���x��M꙳��5�En���yC�ݻ�7O����w,/I���Q71X���r�O����ۘ�un��NAl
c<.����9��ݪaN͵���W���%���4��p�d~�U���n�����l��S�m��e:��x@c��)��oE�:�����Pxa�T#���w9����6�L{y�;���β��siW��������>�N�ň�G$وK��Ĩ�j�w
������vB��<����sN�w�f���c6�e۹�9rS&
7;�W;��GSF�=��j�'�Y�4�����IwRZ�.=a��΁��32p���`� ovW3��q5-R�o�+�=@���<�^��U�X��f��些�/!�fNJ;��p�ڶMS5*��@3�D�	��Ѽ��N7��4)�U�F9�����ų�[����i�	�6��v5��}��:�O.\�u��X����՛2�m���1ۍ���vk��j	��E
O15�.a}&��V/V��9��-�S �����*)]�U�lV��U�lJ2�i����W|A��'y)i�\�}�&ž/������Z�Q������nbi��c�w�3�"��^�c��Ӧ���f��)�U���i��*��xג�cS8�f���ԧ.޺2�W�qvu��bx�U0��/��o�Y�_m�0�� <����A�*uvZ�?R�T�)B�{�ٗn�e� 8�n���<�Z'-�IT[�&gk���Ɋo���C�����F��Vy�[��J�X]����o6��7`^�W1��b��b�@<��y6zvzK����燒�=�BSp[���"r��*�ͷ���c�%�GT�KG1�ے�:���S�>N��-h�!�z@ą����[��E{޲c�h�8]+(������ aJ�M0z�xs����������ꠟn�Q���rT׊�%�A
T��n%��Oi}��1k[�_�,N�ϙ�m�v�ND7\ܙFm'3I���t�f�.1�/�y��|ƣ[,C����3�aӍ��ˣ�AfT	�����W���d�p�(3�I��5��$7�g�wn�j��Ǚ���R8��u���t����S����3lŗٺ9�M�5h1���Ǆe��t�+��J�B�5�n.1�ތ�0[�����K�	x�~���P��fm���FD�e��p0�﩮-�S��m����#�<Gw��Չ\���<E������$���kwE!}�u8�����dQ-�܁\�9J�s�pb�"�\��W:�J{9�#��n�c9:�e �8�u�2��t�iU|2��q��:	��*�ɋ�G�����-�0ҏ���.ӑ,q���`to.L����+��ƒ؉{�d
o*f�/��7ذF���k�P#����)��jZs��lM��i�y��(�֏����a�1�ͽ�s�[�7�5��snV܌CC��2�%3�vH�����]��<y�!��*��}n����l���vÐ0 ���~�����KXw\��;�]KG�4�397����,<*����`yO"1�7�E♳SlX�@�_<Ծ���F�����Yr�[ؐ[����Xj��^����9���2�*�v��Ž��P��x{�������:�`FV=��C�b.���P[{���i�� �)�q�9[�
Q�ƶK��Ŵ��6�³�<}n��>ކ�х�%Զ����2�K��Ɣ`�5$�-fCvgُ�fb�/���!���.@Il����ض��U�ݼN�0��$���ޝ*���ʻ$�t�C&�ŁD����ˏ��F��neI�ۙs:�������sD��Yp[�[y������Eؒ,����S���Uэ�z�ӹwp!~ZK
_��Z��XyH��wh�-F�#�ԭ�������:������7}iޖ�E���:���츳ֺFy7�_�^�FB!ww:!�Ē�t�T%�-�vtN�.�ubuu)�mG6�x�r�e��z6��9�5|�C�-S.±ML�z;�5�e`�Hr��wscZ��\d�N�/2>`:Wq���zMK�w�n֬\}y�ٛ�����7U�g6KI+��S���V�p�����>��u'oF�X1j�;%,��8�	�}�yӪJ��b��aYf��V FcK��u�@�R�;��:����UM7W9�l$�M���n��D0mt=6M�Nї�M�`�Z4�b�e�{.WQ�]�8�W�r��_D/��R�k��.��}�g�ދ��,��͙r��p@蚾��h�;�T�v�i\�
=���r�ީ9.���ӽw-���R'�\	4h�imF�Qh1�U�-���RѶ����TD�[B�DkE�-�,mK+,m�J�+h��elj�Z��Q��e��Z��֥�(�E�V#imm �*�F��)E�ʫ(�ثj4jP�֍lJ1���+UE
�FУ����+DIF�ƕ��Q����[J�Q+QR�Ҋ[BڭiiJ���h�(��+c
��ĵX�Kj1��J���ҥm-iU��*�ҵ��m��U�T�Z6ʋ�
kDR1mP��UYjڈ�J����-��B�m�m����U��
����5��JV��+b�[V�V�[Z*4j���EEڔJ�(���Z�b�ThՖ�DJ�clj�DE���֥��Fն[Pkk�V�ZZ�A�hV��EZ�-j�F6�iB�-�Z���ڪ*��U+D*�֭��mj��JRĴ��H�h
�������b�t�D�m{�qkvsV]�BT���nz&�!jTv&���q�u*�[�Y+�:����iɤ�]'�+�������ְ=2ӓ�L]KL?�Ү���@
�����dAs���'�������s���o�\m"9��.��098"�'C���D�Yд���|V�oM���I��vĿ�^�Lo�x<�s�K,('��1���0�_�� ��x)�Db����W���6���U�!�˷>�yG�_t�%m�lS�T%9^|H��vT����ؘ���
Qa�"�y��Q���a�]߯<v�[DW�\�&�s[��e�;��}�1��(G����q��]�pU���(/�~L�x<�d�?nN{�������{�N����a
cs���mc<M�ƍf��mZ�za�V�b����ݿ=���KӜG!�1!V�D�r�V�>����_qu#���(��!��1۴��	��{ϵE��\e+l���
��!9}lL�9�7c��j�=�-��?ϖ:��J����$y��批�<	i�x�5�f�N��.P���3��K���#�.�N^�V�NiXs�7Q�੄H�����w��
�69nrz��;���lH��e^�	���E�+Kn>oֲ�\�T��Ւ���9Z��I��(٢e����'8�2�-�{��
ü����ׄ4nZKv
�3���G%�T�6�h��O0ě��!�wBss'n,��sv�Fwzd�����������Z(l	�\�=��E�^I��8���z�����#RI�b|�f���jǘ��B���"�BBIBx�I+���ka�B��f���e���)e���͎3CwU����lH��<��`���Qb^;����j�W�s�s�OԴ�9����]MO4d�&s;."����,D�utu�&b�uc�+W����k��O�
B�	ܾ8��	��L��e
~���
�|�s���x�r���[k��2��qy��
�m�`ʝ,�Y��fp[A�a��|D�A�zm�1��{�W7���P+�
�<`7��W�t�\��3�F�r�U<�ƦP�sJ���E��շ26�Z�GT�z��Yv ʧ��z�1KY�{.с�z'Sx<wj���%��`V��I��6�8��,W�y��S~�e9`p��pc�3���Ō���7uf��޻]���Ʈ��5��S��!���N��!�j��7�j4�Tˎ�h�;��2�{3��c�S�YW�%Rgױ�&�Jc)ۿn�Z����7���`���{Iu�B}��Z_z���� ��Q�D��Ck��z	�X�Y�g������R�s*`�*w"U�9[s�tkS�:=�A�+T��Z�{���2M�:��'�����ݦ�9��%8p�S���ֳ|F�P�/�� ޻�
�s-�:����m�*�՜}��\ͽ��}$�oW7֎O�����h�5�d;����W�ap�я��3g]w����rX���=����:�>��F=ag���z]q�˦+�ۡ��t2������g|/��~ܱ��22Ֆ�$��*��hx�P�:��,�L�F��C�N�<Y�t����ZT9��޼�Y��x��2Q�~Ӕ=�ƪ
��0�j,˪KC��%������ WΝ/�W����J���x�^(�qz�Pr��j.��Q�CJ'	���R�� ��2��	�(}��^쵬�)]�HƇ�iʝ�%�8��ڞ�����9S�+��BӍ��K�Sgc���I<�rx���~v`�r���+v+#�V���Oc��=N̲G9�{�o%���O�R��v�oR�z3�=/��\gg����q=�'��G�����C�awg��v��݇���=�dP�#�^���tƲ��U.es�/8�w綵i<�ɠ� ��V3G	�z]�Mn�Y:ۼ32�o�OA���5�X���EK�`��XR뷘n���WB6���,�م����p۸ �p����A-��n��1��݂��VǢ;b��CՌ�b�M��kw���YƜ���೹9�}"��}�of�܃M�A,1OI,R�����1�Նr:�ެ��Ҧ>��ŅfU{k�u�L��f���=4�'"Jֈ�n��
M(0��Q���E�J;��6���ދg'�XgRR�7�0@�{·T�����0ƕL�d�ua������zj�����e!u�{�p/�C�r��A�j`���2�^`���S��xl��=y��Ǎ[��\�uy@\�"n�Eq�N+��rq�d�bMM��.���%�J��m뗸�vn���E����|;}��#���_vo�<ͻ�2���)j���=G�yeKM��;3;|��ޓ�5�6`���T8��p�	n��0��4�}׵LE�-��0l|���˛5m�i�,'��QL�]�?�5��8+�8Z���;�A�v6�����R����D��A�3غ.sC��/�G3�o¯�eRY��y���0T�{ٻ"���`�t:�H��ɓ�
�~�*S2o�9�o�Z�믕�Ư��$n��J��+-���XY��K{uP���XA��/�B����.��U��Q���VW�g�9S�p;b�v	)������H���V.)F�X���W��@�jj<�`l�d�k�.S螾7��LPE:|�D���DӬ����D���u3�C��1:�A*Ǫ�K>���7�n���y���,"]d�����F/�9���!�+~�.m�SC��i	�&7��t�غ}�v�'��?Z[�K��#��4�.�3��y0+���)P��k��򏗦\9;w��2���O�-w��O�{)�y1]��4���ʣO�X�d��v(ly��t���/zS�ד׷T����m���S�\��Q{Y��g1s�͹:䵣��;�����,��<�O=�%�g��Ͻ���`
�G�М�F_����#� ��x������w��NdyByչKiɾ�
�_d�˜��z�} �;ϋ��V�c�K�bP�{��u�e_�>+�����^:�9����bz�:��w�C3&=K�e%8Y��F��م����ȕ-�	M�WI��W{oe��l�����Ur�ϯ21�9�lk���J&J[rC��~���_K�q[�C1Z��'�΅d���N��ct�H~����{O�ݝ^��p�yq+�O�(�y�}�(�1����|tgL��5_5�:��=v(����9��@)���a�-�\u��ӛ)��dU>O]��1d��)��Η[�y��;0��5f�������W����5y��e=� �}M��ם8j�,���n�֣�	d|zM}��E�mj��$��s��j�k�-��N݊��Y6������A�7���N
:8�w+��IW�-��"���~��[����өrM��)tlw���wD�.��|$SD�U���Y}�sb��-��Ԩ���՛^��<��y�X^���f�']��5�)�{)@�.�_H�DOt�;�^�L���������s����U��8�;���;ީ�Y�<�hu56�%mM�8�sI1ކ��V)�L�vR���8�mL�ןLWo)�c+��u���X�q�̶�;�`�}����ʎs�/V|��%�^�4���)h�;ӝ���(��E��<ӭ�X������L= �5��)4���>�����I��9T�(=������2��}h�?v�s��j��i����>̚���g�^��K�I��g����6n_�$��]aۀQ6&e�g_GD��䖧�^��.��1k�;^���`(G�w~}��7��t�������v��-�a��^�R�*���X�w�����������ϵl�n��w�[s;lQ�:y��v�2���ӷV�=�+7�~jŽ��g�.�ԇ�����왎4�(�����o��(�J>N:s�+^ߥ��6T«wʞ��\dğZm����fod��X���({�q��1�ϔ޺�閰��,co�Y͑�����)<��_��[�'6X����9���i�̵wu:'���j^Mi��O���8��̈́%�څ�v�Ag9�օw��Va�*��ɻ����}�7n��gQz=n�u��hp1.�J��E��6�'i�J-_e��8�=��^�p,a}�=/΁���L����t�c`��z"�D{��t���4H�f]z�sݘ��U�Eՙ�J�]�Z�F{]���^�_=���p����4j/�qz8ж#��z머��<6�Ȭ�0E��=4Nl���n6�0Hb�=�b�e236����v����:*ܽ��E0l��f����m�GeIGR�v��^(���I��������a��=����"y\��9����WK#ӯ�f&�
�X씯���^�q�sv!���u���zP�C]��wɬ����h����N�h���ם����KWx��B�c)�C7�9������v+��
hS�؃�z�M��x��,ٲ��j���EO"ĩ��T����d��M�a�*/_�z�`M�z�n�ik�$�������P�z��&ɕ=N�?s/��{�+�n�S/�Dqb|Ī[s��N����>ί�)m_�V��R��5_��w4Kz�:[��8�f���wV�C����|$a�R�/P����!ؚg�����1]:�W^���w�߷=M����p'�l]n��Q�����	QWz�oU��]�=NEO *�_\��
YO�Sg�H��TW��qcv�6:̣���Gڪ.���hcq3\�,3�{ud����h��ʗM�O%�i] �efJ>�H^v۽�fN�4&N��U�rdZ��b;kX2�|c�t)�\>��[C%����T�CGR�f=��R���*؝w˶�[�)�����]S��sw�mY�%�k'�Y�|�������^t�Z����	��q��n����s�����3$b�ʕ�!؞�}w���TX'R�P?s��>
=qŮ�^ٱ�l\�cx�f!�3��i)ֽ��KD�TzֆŽr꟢�Aɽ�OϾ�-������h%5S7y=
�[>':BcV�tH���jy��l�3��ot�qZ�y.A�U,?Wxw�hU�6fŠ�k���z��^Q?ytx��o�w�d����X�Er������w���m�����w)QIŴ�b��D����2�b�x��� �M]Q�;3��G-��1�??��RzkϪz��s��}y2]̦�*�C��՞��ū�<j4�W~����12�h{s^�'�!���78(9y!�b���.��/h{7�r�N�	��β����ʄ5�T(ؠ�yc؝�KN9�P�v��.��w��)�dY�5\���C�ޗ�|y��B,9�jUl��`gK���Ci+�l��J�û5�+����L�Y��tv�E�vs(</)@u�weʘ�=ӞőF�	O�}FE�N��/n�%9���y�Ӕ��A���ut�ݻ�њ�>W��m��*Xo�����c�K�e% ���\�LԺ�f�!v[�P��U�u��U�Ù[^�j^:����Uwk��Gۼ|f��;���[�^��χvЋ[��5�ϔ��lՃ��%��L���*�X�����m�d�,������1s�^�}����X�{;x�3���tݽ���ܗ��2�����o��V}��+=��Χь�n��ӎ�$Ӎ��_�{��M�i��+�����jz�:[��r˗��Q�V�#ύ���ȧ ��9�o�yH�/�(-a�yT|�䢰zU��|�qG��>ʉ{r�5����t�֣jw��z�h�i{D����yc��W����L'E����CU�hxvP��ã��J�g,��
���n�|��Vzf�8�ʫ6.��z�f�p�6�#R�YD;�r�)���ĚVkjj�.f�S��wG����bk6��f�5(��J�_����o�aowoP��x�s{vH[]kta �B��w4$v9�D9�]����.�6w$��l}atv�VtikK\X6�+`
��ΙS,��/]%s��oDI[|3���,��+2�.��\i���)��j�>Qt��τ�f���$Pל�`�a��Տ�uw:�����!bΫ	t��������%	�v�R]�*}������+�;��+s��2Xe��(�Z\��)<]@��5!�G�fv7�Ǡ��km���p�:��p�5x�cќ��rs�w�#���}��ˀgr'����+�y������L�����Mڣts�`�W���j��PZQT'�vcO]JM��G[���Kt�/J���L`{���F�]� �Hqɬ:<Xy�{NAi�;��Ȃ�.���z��t�;:�'9mfH"fާJ��%�w8lr�����c�L8��2:M���}���چ"�&�
G�o3[�}(u�R�����k`�:o$=[n].��k*��G4���M�6qZY��n��hK�}��0�C}�f!�LO�7b��RC@E�oC&kYR��|+u�{�]�.�B[Y�˘�aLt�Z�o��q.����S^²&M>TW>�঒��Ck�P��+.�!�Rt��A��m`�<3k~g��{�����ה� ��Sb;ϲ���C������V�����	o��{��_F����;O3�Ɉ.��Zh7s�n��\���>�YXk{��N�U:J�9�es�d�C=��썆�Y�p�0����C�Hr�V�۲�vu&k>"T�o��h::�%v*�,��7돸�z�r��W���1�}�]bE3�xs�����I+��S��k˽\���nRx�u�Zҙ+�{r��V���H/�s�v;ZG&��@��D��{�	#s���[�Jx8�|�I[0���Ma&je��ń͔��qreˌ_b0�ȥ�t�2�;~�{�d
��>ɩ���+u�y*Z���$�{1"����g.�:���\I x�W<���'���j~�#������� ��t�s:N��H�q���6�����Mg(�r5Z�D=�]/g[7���]�u��s�ɷ�L�M�y]a����S2,�WoKj�U���{�t�̺��=Փ�@W��k���7T�қooDb�_Ugn��(p�s����BnlE2�V��f v5��؂Q]}7O�����#ν�lJ>bD�G٦k����S��'��y*��5��i��&��ZvF]�)A��+%�.�e����xb�'m��$T�}J5h��c�]>'��N{ϰ�59���M�Pҩ�Gm��P�X�fs��y����S��KjQUe��EhZ���DKim���Т��%kR�j-�[l�(���X���[+m���
UTbV��lmX�+U�#FR��V�T[jJ��#VְV�
��Z0XҔeEh%(�J�R��cm�V[eQ��JєZPmm�m��X�KQj�R��[AiF�mV�����B�
ZT
�"�µDTJж-F$X��Ѷ%A�X,+*��U�
��
ڔ�l���Aj҅AT*Z-AX�TR�++Ym���؉E"�%�X�2Ք���
(��ղ�Z�J5�UE�(T�m�ڶ��ն�PJ��e��Zж��j4��E�����[KU��ֈ�EQm�1B��
�Z�EE���6Q���"�eZ�iE
���im��6��VX�icK+Z�F�(�lDE[Q-���R��-�kb��V������֒�-�Z���b"(�le�Z4�Re�*R��j#A�im��F1�Km�)[�Tg�@;�=&3���g����x�����/x�&h����ʋ9�"
���W�����hgb�)w62��c�>k����k��qt�}"y�j��?�xs�wV�N�e7����v�O�ӟbn��w�6��yyT㻘$"��n����nh|�W�t����=�(�w�K���-��k��Iǋjd����.�{�}�����S��.{W*��*kM>�ݐ7�(�9��T籵+ҫՔ�&��ي���Ժ���3���\��T��^�4�P:T��R�l�C&��P��U7^ڷ'K3~x��XOw���Z�ԩ��V��I�U9s��4�9��c�N�k�t�mEv6zj�g������ڔ��}�rRܙ�IuĠ	����1��+���t�c�*e��J����yxe����5dھ�t�Mr����*{b��w^'ҝB-�n��S�n�����̠\ϋΚ�����l�^Y���{�iC�L^!��`��{�X��<)��/'��O�ŗ@P�!��q�RI�XG
��p�m�����޺����4e)�'��|������N��l��Wj�gS��f�ز����OR^þ�ԏb�.h���ro��˫�Xqt�B.��G��]/Ryy��˛�N1� ���\'o�o��]3�nl��Db[��x�ӛ��?=
3(����%E�x��d���v���>a�۲��
=��z�͉����� <�t�]��;�N�f��8]-
�r�L����1�\���W���|�g�#�f"[kRӱ.�;�N˯?@�բ=�|��8���̧�+�X�@X�=-j=�������k�EtJe���3�lA}���"˘7��?�Om��&�X�#��\ì���I�ם�/)�νZ��3ny�ZsG���:��M���}-ܾn��_;yk~4�oZ�[��r���:|�Zw�;��'z����d��e7�/�@?;꫉�:#�1W�W�T��q�����lϷ5�i�gk��+9���>Q3��9���:��2ּ�W��:�]�x����������kY�jݣ���5b>00�x�����n �����@N���yP����
�hY65������v�]��[�e"c�3Sg9(jR�yw7Is�7-c�f���nf�k3��&ꑹk/�p��O���t���P�t�,��+|�΋ƶwE��V����X�t�ut��U]u�w% T�Q�'9OJd���:�#N�/]������?<ܳ����IO\ǵ�jp�r��X���{xϳ�vc]	����_�뽷��X1�,ۿ��yoՙ��+u�|6�h�&��k�]}q3�U�V�����ݵNrW�0lEm��j�5B���`����X��Mj}n�rU>�)e�}=�L�S��u���0(�yՓΏF�/.�rk�9�V����=�<�(�)�m^��6%fK�a�3U޸!��6�/��c���Xp_Դ6.���R�y*p�w�w?9��G�N��O{���� Օ�tOK���Xغ��M��z�Μ���;���:�tf7��{:f?ߠ�*�K
�J߾�*�p���r�{�X=�@X�5���;S�޹�Kv����ъR�]X�� �|�r��r��7|���#S�%��x�d�8��Ūʙ�4���\9}
��y\§�W��K�˱���K�dݗX�K+�^��S<�I�:����12��ܥ���ٕ�䦯t)6L1�~��R����	μ��)�o	Hl�]>Rܺ�]/��Ӹ����belgZ֢y�eL�����ʩ�_��LxYq��]�����]=�Ԛ���ֹ��ϳk����c��ъ��Љ�ك���z3�&F߃�~3����Ki�'�_	�NK��s��w����!f�9Ov�{F;`�
���k�:=j��w1����C���3JR&�͋gT�k�fk�&����6������̝d9��I�N���0��M!��Ǚ%J�[���o��3������M$�	�=���'PX;�AC��%a�{�2~�p~d�a��bJ�w;ċ'�`~1C��.��?2u��Z�i�M$�M����Y��.3���3�k��2�d�s��	��<��*~;�2u��P�N���z�R|ɯ�ē̛͒�d��1	��O&LXy$��?kԻ�w����=�o8ƹ���|ì'���,�ağ� |�d����!�37�Aa>C=�2u*&���N��*��M�foX�O} 
k�!G���8<b�G��}�����ϱ�s_}�v��L��,6�q:̚���BsT�?2y�5d�2y��x$�C';���$����y��P�ױ�2ot�� |ɶO{Y��0x�s�-��>靸��V�%o�H�yt�]�TNQ]���C,	���������Lņ��0��ϋ٘���ev�m��!hPjC/�u�y*��{$՗��������me���vh�մ$+��"0���������;�E:�5ky��p�N/p��}������Ra���Ő�:ɔɋ:�>J��hy'����T?2u�!ϱ&��'���:��p�q<�d�f��d��k�D���O���P}�}!��V���O���Y?02��R~I�g'���ɜY��*~���I��\�<��ϩ*N��*rwx	Ԟa�k~ؠ��ӿ�ym���z������q��hq���&�w��'�4~�$�I���Vd>ed���Y��'S8�&��g����O����J���k7��~��o�ߝo�%IԙeO��
ɶ��x�y���'�q�'Y>�I>xɟgu��d�q%I���h|���)?[hy���S�hu;�>��s�ߵ�n=�w{λ����C	�I��~�y��X� u��P��bB�y��`㴞d��^� q�M2h�Bu�dϳ�VI��;�T�H~-�B�u�s��j��}��s�}w�����z��'�$�N��L2N;�2q�!���'Y=�r��I��xɦO̚����L��$�~d�l+	����'�c��>�s�{y�s��?x�	��<�d���@�O$�2`��I��[$�>�d�C]��N��?by�l';|��,6��i<�̟0˜��q��{��?�g;�~߾Ʒ�}�a8���Y'P��J����VN�d�b�ĝI�Q��&����RN�=��
��=�y�|� �}1�\x{n���8���q}	]g}iWvx�&�m����fY6Ś�p�m�'��Y'P�w8��a1�u�d�VJ��d��a��'ɳbjO2u�^�����|"�!�'7�R��u��]��J��9�e�&�S�I�� ����w�C�|ɹ�`��<�0�%J�b�aY8�8�u�l��J�� {�������؃�q���.��eX=����|�j5�G#�NYkX˫��8��HD��>�M�B��Yx�tܕ�XGOqR&�˷��)m�O����Hfe ��zf��y	�	�%ޯr^e6���ީ��K9#e;��>��+u���6%���gFԯy�)?��r��M!�Y�O�?�{Ǚ%JÝ��y����2��)�؂�Y>Ag=H)4����Iԙ�%ՒuɺE�ΐ4e���`�kYױ���ky�7�='�.Sܰ�&���&��4��>s6̲yNsd�+�Ad�~��'�u!��b|���JÞ��$��^�����cNe;�__�������dzc��"�N�<�1a�I��ɫ�u����̚I��`i��:���&��� �J��w�:����`4�P}�G��q~Q{g��ٞ�|��2��Ng��m��kWI6���,&��e����g�:�����k�,�I�gx��e��8�	2��l�py4}��U]����u���I4��o�p��%d<{��u�n�}���8ɞk�>`|��a���o�e��d�%O��y�XNi��N��}ϱ&���} F|_���v4��c�띧����� �?`�2�iC|��N��h=�d�']��ϱl'�}�IY4���'���P�,������ŝd�%L��
I?+�^�u;����l�Jf7����@U�1
���J���O!�w���5y�̝~a;��0��'�Y8�4��J���(m+'�fLY����ͺ9?3��"��/�5���q�z�	�(����qP�'�3ϰJ�̝J����C��=�$�K�d��M�{��i�N��q��;��J�l�7���9��&o���k}y�9�9�R�u'�zb���<���N��g���I�<��u��X��J�̞~CG��
��?g��݄�&Ow m�&�5ݸ�y�NWt)�_'3���iڼο��{�p9xǍ2
q�I�����'S!�a��N�C�3�I�<��y��Yw�:���=�!P���|퓬��w:�>����K�J��'!x�9l�Ͷ��1C�Qζ�u���=��{��֩��dn�YIfP+=i�s��Q\�g��f�7��M��^u�~c��z���6g)Z�{j��)Ձ��j������L��jV����v�&��m���ˌ��'x�*��p�%��}��P}����w�?�4�l2���?2u�VI���ؒ��0n�!Ru"�ĝd�}��8���48��'Y�P�'�$7;�@ǆGG��m���u�S]X����<e�i'�wxɦO�5;�I��&�e���	�e�=�"�:���T&��+'��~1@��q3��u�$�����q�����2�l������k����:�'�su�i��?2i�����2�h;�I��&�e׵��C,�k ��C���*I��ԕ��=��:<>�{�bn���O]�N�ٿw��������'�o���aϩ�'�6sx�d�|�����d����:��}Aa��Af���d��`�;�������N�ﱿ��g\���3�o����w�ؤ�'̜&g�	�&����'�<���/Y2�;߿I+*�w�<�;��̝AHw�
I��?������e�s�M��3���x��~I�k��'9dY:�X���i��C̝d6kX?2i��}�b�̚a�sI+*��O1d�O�;�̝AH8��r{�1�}������P�&ҡ��� ��������$��N�o,�:I���ì�Oə�d�!�kX>g�4é?n��~d�w���|�QCg�����)��*5AL��
ISӽ��N�Bs�i'Y>J�g=��~�g2O2g�ėV���	��L�a�I���j�Ru�֩�~g߇�}ԟ��|�8�oG\��j�ğ�Xu&�_~�	4��s��	�w�<����}f�m�ﬞ;��N2d9�m�y�3�O�ɶO&LP�~d�gt}��|En���y��H�~��vg����a=߰m2��M~� m$����N$��<�d�g;g�u��ϩ�N�|���� �l6�bJ����>@�����h~�6�?y����S��mk��#�R5��f��ϟ�Ec�!H�J�|�-����򥜲���V
VLm�&�D��X���c�b�f+���kϕ�`[ie\�M	{���c=��9[�8��t�R�K��֩��3�B�Eg]Θ�{3i;w�a�8z�ݻ���{�^�|�sy��߾�=���$�*~͇X�Lˀ�'�Y2� m�y*k��	�a����e����d��]��y���|g�I�I��?�#�����r�������xǽq�: ��d�!�C��ɶVq��>͇�RLo.��J��>�*N�u*g�b�<ø��2O0�{�̞��{�{{��Ow��=YM�vo�wc������~}K�����8�	Rm ��+'D>Ł��u���hD� ��w���+���*O2{���!Y<Ý�����_�~֌h�3�}�o�>�>�,��={�<��i5;�T��=�²M���ĕ���a�VN���i��fqp�q'S?�<��'�~�:����=�w8޷����[0��o�y�z�5w·:ɗ�{�ą@����O2~d��`�d�M�+	��&C��*I�~���+���Aa��C��L�$��]�W����s���_���Ά�	�{��2{�!�CL�d�9�`�'XL����Ri��&����&�e5�b��N撰�C��ؒ��6�B�y+'s���?��Z�;�:�߷�����T�d��0Y'y��kƲN�C�bd�솽�d�x�S��e��|��$�M�p��'�,�a�׵�0�Of��:������)�G��>��Q�^��di����UU�+�+�2��(I�N~�XN�m�����:����O!����I�5�`�2N�}����>@ﬞO̟ ����^�>dEB߉j��1����߀���x;@��$���J�$�ĕ'Y51I�M�y���a:�����4�̝a�R�O�t��:�T���4��'_���K��{DW��픥�|.=�D���u��d�p�m�!�`��<�'u�*V���"��X�Ru�l�?���<��C�>�i�M2u�Ӝ�g�4�L�O��o�Jw����q�_S�(���Z��U�����g�;��]6�ꊼ��6���W�M��Vs�J��>�f�I����;��\^��c���E��w
�jb�.�.ȯwV��������j�6���R�ǍF���9�&�_����n�qm�������$�	�2s�2��{�AC��%a���'̟���'Xd�%t�;�x�d��ء�I�I�Xe������߷}�k�{��k��|�'R|��� m2��9���o�<��*~;�2u��P�N����� ��'߾ē̟�$��'sbO̞M{�Ǯ5�����������o��M9g�he��O����M��O��@�2��Gy�O��7�Aa>C'w�̝J��ױ>IԛeCS���6ɝ�I<����#8EK�隻�Fo�y?��Ǽ�|���d�dņ�O���5C)<���`�2��(��$�d����&��9�O&Y'����N�Bgרd��O���WK�����i��V�C�T�4�d���O���M��g2�Şd�%g�4<��O��*�:�ɞ}�6�Y<�����O!�wɖI�wX^1w������3��kw�9��}������x�'�;�O�}�<�>o�%d����8ԟ�u�1B|��<�ŝa8¦P�$Ѽ�2y��RT�I�T�g�[!6�t��i���@�ǁ�1�{�x��<��{t�	�l����8�uɌ�J�l��h|���B�&:�b�d�Cɓ����Lu��?Zc�{>�~��g����2q+��	Ru'S=���?N��$�a��O0��N�}�8�|�3�ĝa8��q%I���h|���)?K`m2uk�T���k9����?����ַ���$��S��'�I�x��N�`o��|��On�ǹ�
���8�'�?$罈z�L���N���=�B�M�㿱%I��~�s��sf������w�{�k|��*��,=-��4�ԣ$�N'�L2N;�2q�!���'Y=���@�I�ݼd�'�M�X�Ri&^��u?2'�K�]�����{�ifQ�9��<d�i����̑�_���+5)6o�m>E�=�3��"����-;J2�֜gOp{��7ʱ�;�+wʬ�b����e�v�3�F��<}[X{>e���.�wr��u�\�1��	���[P�F�z��]�����mN�r�����xm\��t�o3���Ǆ����%AB|͡Y:��V�ԝI�g$�O&Xr�'Y��`8��l����&����؞d�	�wzɦeR��ܫ�%�f�;O�l�_!���c�����'�,���y����0n�%d�VJ�ĝI�Q��'ɲoX���u��ì+�O0ﻃ̓oP�5�F<��nG��2�����C��~���bO�;�O3�'�Y�g<��3�`I�;��R�������Y?LRu̜�L���d�~�؆ړ̝C�~�����w�Ƿ������= �I��a+8���0�$�`��ԟ jw؂��O�Y��Cl���~d�I��T�&ް��t��œ��d��s���3�����n��檳�������z����=<���$�2�&��2J�����a?&{�L��
C'}�(u��fs� ��'����u'3d��N�w�c�W�w�U�W纓&=|����c�U��!?;M0�����kO̚a�� m�d���<�*V�<��0�s��I��{�O�u�iXk��&�w�)�pS���rh�f��gg_����ǽ�ֽ��$��E�_�8�1a�I���̝d3�i<ɔ�a��L���/7I4��}�u�T�)�N%d1��y�^}��F}����u�i�iX{�� m�y�$�d��X��I�O&�XM?$�2b�XM�ɓVa���m2��I�w�8�Y<����I�<���ڹ����{��������4�d�Cǽ���J�k�4�̟?$�l�6��k�>`f}I�Y?2u2b�m�L�8�����͇�u���8��A@���k߽���c���y�No[��d�߻��:�{����Hk���N��k���O2u�O��6�|��ĕ�HIƲa�P�Ő���<�������}���ۍ���?��-ހ�=����%��kŜț<�&���ӣҗ�_V=�oM��Q�&�Q��^��W����;����F��
P�`��]��c�S�uf��ΣXRM���Z�YzB�nG6�'	����a�x[ W7T�oT���J�Ng���s/���f�/�L,H��T�����mWT=��wuoctU|o>�b�^�yO(ew�"l��="�]8��ξn�5q�8
q=�H�6:���l�F&��R���ʜ�M=�Mg���5�$��4*����y��%�:)Pþ�$q�:v�:u�Zs��q�0J�ۦ ��&���o�{=p��L�(��
}��vN4�v�p�'ʎ��\�k.׃�����T�=���������)֒,%�CL��K�@%,_DNڦ�Kҕ�X{�vGX�tEݍ�W3U���k�|��L�<�}BZ�'��ݓ5�+�.�FjI���n7!��fͮygt||�n���� ��`e�׎�n�C��]X=-\yW�NI���*�V�IYy�xv��¦�Y5�`�]�w�	p��8Zx��s�/dͽ���Ꮙ��l���d(���4�[
�mu�x�Ex�pح�/&9)�a[9ou�����q���L}������n˜�A:�T�ըd�4�w6����Y�i�k��T8�$̃�z��)��Y��6�d����mA⚠հ�nF~�h����|��mF�;�j/�22w�x�7���YB�MR<M?�J���g�AL�g<6�p�]����
Y�������K�nȆ�u���T��ۡ1T�W���EI�{H#��<{�ej4�$�4>���U�mj���˰mM�Oj��1��5g\�o\y��zN�H�2D�����yl�e�L�B��`�z&p(��{n.w+ou6����mŹAT4w���;|E�ˁLز`���ז�.~i�3��C��t��ڌ���Rao0p��F��7KwT�[�C���͂^qH��u�RE��HS��Eb�f8p$c%-���0��bǣ�`j�i������z�����hT�{�tVF/�T�W#�(v+/v��숲�֫�Wo͞#;��Ԙ�-$��=M�k�c1K�T�)0�����/�����!8���+���Xn�2��XN��PxW�ʒ���J�u�g�k�o�[+sp���7Ӱ�Ǌ�kw��
�a��m �9�Gq��T���]%����W��cN�K�����E.O�}>iՏ��fN�t�d�هk+z�2E�m��$�Q��-ЪN��0ɻ}�]{.G��Y��������3��7�+C�{����V;��\ڍ�8��7���t��[��'9���K]�l�W��C<�%�߭�=�6_]�^d���2'�y�Vh���V�r���ڏ���	Bk�wq0�$��;���W9b��<�Y+�����N��&����}�5������JTK,*VQ�ibԵQ
�4�Q�U�Z�"��aR�h�j���Uh�F��Elm��`�mm�l��+X�D�D�hQX�"QkUZ�XѤ�ij��emceP���YEJ*�E�Uj!R�mZZ�Ѡ�[J(�ыkR����m�m�-�-�)h)X�YE�Ue�6���X��کF�E��*2�ĭ�ږQj�D�Ĵ�V�ѵ�R����Q�єQ
VҶ��KD�������lm,D��QE��[X,mX�)V�%m�ڕDU�B�2�,�jQm�¶����F��*��cQlQ��V�T��5+`�J�T*
����RЩEJ���c%E�eQhV)DR���+h��-V����E*��Ym�V*T�*���h��-K�Դ)lU�����+lD*�Db,���,��b��(�Z5$X4���VV�TV�-ij6���T���+X�Z�H���kkJV-eKim�(ҨѴ�mbԢ*����A
����)[F���mX�U�iJ���%�t���S�h�zS���mX�o��B r^t
��r�vqξ�������n����\
=K�����������>�T�7{��@��j��A@�>�*N2y+;��<�w���5y�̝~a;��0��'�Y8�4��q%d��r�Ҳ~I����r�'��|�|��#i9��G�O��\2O��3��RLo8�q��X9�	Xu��Yߩ
��7�b{�I�/py���6��{�$�<I��u��z���
��r 9�����y����cã�<ZJ��N�3�P���Ɋa$�fO�<��'���u��X�%a�O:C��$+'����{v��o����3����G��ٯ��M\���~��ĝ�IY'���+�
y�I�
Chy��R��I�����$��Xy����4��O:C��$*9߾4y����%e��ߵ�^��}�}�������o*~��s"���u�	��I�/W����
�4q�I�խ�)��T�N'~U2L����=�b�3⚺4�w�*(�L�+�{�1w??I���^����S���d����N�?sl�#�mu��{��yt�Qrc�✥�K���]��9�\x'��G)ɲ�T�^�Vv����\T����9�`O�ˣ"������]�'#�]u9KiN��d��������vv���S먆��iʺ	�����M�k~w��J3XvB��gYR�PLh��S���WmSBO����`{���U��k��^�U���a7xD6c��J��.l����A7�����N[��x��*@�yIN{d���s������=��W�ߦ���G5Mتr팛ޱ�w�x{�"��HG�>̧԰�~3>X1�V��ͺܗ���ػ<���}�u�a޿6�jgûhO�kb��|2���l�X1�ͻ��]e����;a�ڢ%7���伪W�%�+_Fd�ݮr��.�GK����V*�n�d皚\ΉJ?SεGzJ;�'��29���s������;��{��mw"m�O)�j�Tk�GWKy���.���\qm����՗��Σ�w��ҍ��ǐ���=n�u���O\�~�x�g?m��k�g9��9�t��u��K�c�CDvW������卋��M��w���K���`ϔQg��臓�`P��8J����\���G:�s���s������)�=W9Od�Y�	��1��kxJT6{WboW@od>YۊN�Z��v���'��[��w�<�T��i���G!�x�AE �S�ĩÅ����vu�obc[siY	J�5Y����9Ӈ&j�9WH����[�e\`�Etv5��Aҽ������h�W*�mY�
�WI�r�
z.�Ronڒҕ�]�j�ܮ����X�b��+,���y@��]����(j���W�}���'�w�@0&1Iv �Ns��^,~���Rbڙ/�\��nm���s���j�R�F�z�k�������ۊ˶�����3b�5�CB]{���݈�T���Tvs_ũy��t�S֩^�<���N�mMUu�:������C7��I��hh�@�R�!�Y���M*�宙Қ\���}'��r��R������T�Qw��j�Ҷ?w���@츹e�׹��K}RS��1u�9�dV���6�mEu+n����_�ow���~^}~ٙ�&�m��kg9Y�>�_�5��7���ۖ�J����-M�V�>ΓH^�L�yo׾uj�Ү��t���o�b����7��}�rR�z�q��gQ�v^�\���Ju]�</�[<D�w��+Jlno��r������I�ؿW!��:��}�<;k��^�}7S��;��
xx���A��F����1��cSv6N^�e|�ؓ���
wz-����VkΘ�V��8�c;�nvӛz�{kn���GC��:�;}��nj�Eu_sW��yn�6ΎqY��]FR�pΨ4�T��9�O��UW�UY�!��x5$�I�����^���=0�������{�8�6Z�k{�	O�����M�3�Kj������|}G����n�6jI�5�*R�a�I�!=WOd��TA��;kp�@�6[0p�������t�ׂ���~��k��3�nĽV�g��yi�����L��{:f�O�Q�����?�[�=�����;)��Fn?T����ow��\�˾��w�޸�ܾn��U�[�=9�jj�o�LaE+.�:
��k�M,x��r�i�\��ލ�Y����t9t�3�ax��!wl�w�}��/E-tT�Z��ܝJ�b[�P�{��{jܝs=���,Q�=V��ٍ�ޮ��k/�{�}��z��8����9��#X�:Wmm=#u�V�l�>��ᔀ.j_5UW]�i��}O�RqӘ�j���Z9{�#X9���T�,R#�$��,8�nյw��c�l[X�=�&@�2�J�g>����C%m�͆0m�9>�-`-����eB��Xge���c�WN�ϼmk[���ۨpbۈR6.��F���'la��齩��{�  ��o���;F|:VHʊx&��<�U�唸vSaOP�	9-�=��'����H�G����޾Η�3�|sl>��e���_+���gb�N��U�r[}m3蒽\�d�ݵ+��������������_�`�Te��v�*O���K�*��-�^g��ӤZ�v����{��D(�;�.	#үyZ�Jv�8J�J�T�HS�,�r�x��9�����:���sY{~c���ěa���K�[.��Áhl*z'��e�C:����{;7M�{�Gej{�Q���!E�<�+W���&��=���¡b=���,n�|�w^;�=��QC��C}�:g˗>^�C�lO7 �Wՙ���^7a�'��9�*�5��㻩���(���Ti;E��O{5���{:SW����z��+��ԩ�u4�f@��l8����0����*���}[�+�o�{�ژL]���u��u�N7���Hܛ�6�[�-x�!��p�ɩ��2�����}{B^V��d��p2@�:��v�]�C����;�%��)�cغ�����-c:����>��8J}��^�ɏ
�룜M����I����x{� ]�|��_�ʯ?��~��l]��g@��S���ә���.��<BƜ41���7�������;{Pv���rs>2���r�
Ďoت�V,�&�v���/�����`\����퓾R��w@=I��O1�m��*���t�׷okD�~v-�� ���f-�K���ͯn�~ ����f�=�(6�(�m:���R������7,��zW��}%�=�]�~�1�@�f�בܝ��jt#�Ø�)[��>X1��iy.��Ԧ�߲crE��}�\{֖��Y��'+m�b�&��7�Ύ��[r+�7Jwz��ӽ&nȣ�{�k�:�g����r�\�n0�#���{�.=5f�o�@�Ӝ\��q�F/�����z�ut���E�x{��`�]���-�dT��K�ԥ^�
>�>��^�<v	�=��F�A�װ�-���Xr�Rq�����;m.�����P���=T)�������2E�e^ջ��/�*F^_5';f�5������I��Ź�y:�r�뎀��
�{o�
�<�t� ����9X�{�u���j���{ԗJo�PΘˁ|6Gb����<=*�fm��=��#��TCVT�2�c��Us	^2������'�^Ve�GSc�w������;6��{!�b���
1�w��ӫ�4�fε���|�{*!.r�S9f8�c�u�:O�ݘ� ^��\�v�]�$��4�zZ�{�3�n�Q�D����$�ʘ��2���p߷�ə;��R�=�QY��؃��vB�3���&-��K����Ƕ5?QW9�3ڗf�}A�>��j�؇��t��1����.:��{Lp��������7ٜ���w:�eG�/�a �{kϽ�v�G��"Ћz�y�}۱MӰ�-w(O��G9����:Nz�ѵ���;�3�NBq�[)5}��kU�J�I�r�_�SХc�i`�}S7ڍ�_�"���6�k��^��fvD�ͥ8_9C�W[�<�({X�smn�Sc -75y2�|�����g2TO�QQWv�HI��������ݬ�����:2���V���sAS����א���Y|uUn
�v��m�r�̷)�X���++45q\6�.!s.v@�����mfV^�vP�ܳ���5rOp�S�xxx{í��������X��f��s�fmǷ�n�ȫ���q����hޚ��{���ޒ疾j�SƮ�4�\��sS�md�xء��y��gz�'������K0H��mU��y�n�B�|��
����6x4�=��w����[M\�-^gܛ쭎>ۓG����f�����e�2�c���u�/U��E�096r�7�xk��1���S��f졺�N����qf\�J}���A>�#qEA���5]Khxr����N�n�A;ϓl:�K%��?+��ž�;j!..�R'�Ui��s���z�n[�����Ĭ�rw�������|��.��Ƣ�HT���Y���縝�ι��x'����������!��+��TNbyQ����q�a����w���bߩ侹k�򟝊� �)�4�����ͼ
sM �kX�	��_���dĿOc���Շ���a����/�ܠ�:Y�g���m���{X��.l��r"�6�Yn�T�Nư�F���=���>,�-�Q��7��V^���b�da��)=���J@�5;<�Z������N�W��A�s�o���_W�Ev�'M�Rd,���'�w���r_VUK�s)���y�=�qz��7���;1�_)�l��)����4ķ2<�q��ӓzg���w��CZ����TƓ�{(���{�yԻ������=���m'��WI�VI��S�u��+'GR��[UUu׻����)8����=�*�z���k�f#|$�ՍNa�ڼ�2��V���=s)�9W;'?������A�%yj`'�(Jm1t�����t����m����=�Y�&����X������G�;}S�<�糩�c&Mޏ��,�G���t^��1{:1��kv.��.$�ǣʮ��y��/18�*t���m��8�+ә���k�D�'oҋc�n��aJ�Z�>r�s((�s���ٵ���~��{v��{�c��O�O�;;�ew��|�6�ԤS�xa�Y��<��hu��6�	��M�7�NK.�Z�;��.��U���H ���Õ�`=��vH{]���`�x�x���=�9x�e<��^��Mk��	��8Z���b��F)Ա��b�j*�݈v�7y7@k2k�aV�v�m����J�s/��� S�i�9���9Ο�@E�wEy��O3
��žnN��������b]�}vdrf|�Eu,s#*68(��w�-[ j}v8eA-͡�=�5S[Қw�A���uۧ�L��G�u�'.�'!��m��_�6�~��/��n|νL�T�y�&^}1]���b�:�㩏�z�v�$��
N,A�ֺo��^O^��9}�K�ʙ.�e=��,!�&r�qOWj뚓�#���k���l�mu�.Na�	�=Wղ�o9��#�H��~�˔���M�Va����Ϫ�[��?T���|���()ą��7�R�*�z:��_L�����[��V��Ϊm{xKc�~z�9���>^ٶ�W-�䛫�)�w�k�Ù���娺�y3��ﻄ��[V�Z�X��u\�}OcT�߳j��A<�W�>��O���;�B
��_w�V���.�%j��S6��+�Iuu�9R�7d��r�/��2k���wʖr�PtZ�9�u�inBU��t�-�Iu�7�o9h�ї��ӓv5�CX�r�yʧh��rJBkvPg-0c��1���;�}��9�^�)��u�l���K������1��4>�5&����]y�~/9.�&�r2��t}x�O<�O���%��K98+�o���t��� 5�o;<�j�m�n��j,#����]�c+3ub���-�`Ĵ�e�{����1eF�mGͬk��SLǻM*�w�f���Kha��{��e���"�E�Qw(34�/v�Н��t�':pڒ17�l��U�y��\綯ý�sj�ߑK��ˋV_))�}�f02k�\X���r��3֢�Q�7�<<�Ń*9��vS����)&<�)>n:ӣM�4yNN@~��Y�=�c�B!c��}q^�B�G�U�Ԫا��tܫ����Љ��us�e����������쁈\^ݾ��q��^����
�n},�\���f-Y1�� =�Gv-Z�)ٶa�t�K�����zgk�s{xA�-�х�,��E����lY��m�08+�{��ɷRi�[R)��x,:��q�!l����3S�̯���9z�7ŵz)_^�_]J�EE��c-Վ��Y5(\�B��M�lpޙ�!��T��D�
��ϳ�i�{������j۩�p�S�s�LW9]]�}��)9^��F��-k oR���T�h'�Ċ4C$�L\�J��Ʒ۞^ǏŮ
�� [�R�H�Q�|z��9�l�g�;q>���<�}����y/y]��^M��f�P��y)������d]��pmO-�~y7���q��q�z��u��d#��*;��V�t��Ud�L�:�ʴV��%�;�{zE��.�{:
��U��N��(����r�hl�5$&P�_
���H%�����xcA�<^M8��!�����z%��q�[H�x�a�-�)e�ʶ��H���.���Z�Z��\��
Ü�ټ������T�z���Әx�-Y,�� {��bt|�N9.QG:�k	Œ�^����y�݋�:c�Q�DQ�H]��
I���/H�Y�?g�j/ߊ[�m_�E�.x*��ő�i����Ҏ
ɍ`��b:�N]��A���Ni�Kg;�p���P5|�ϐ;�՝�:�ȵz��qQ��s*t� �7��j�Z�o�����qvݷin����p,�U��`�c�0L�q�R^�R\<b��k�N{(gWs����s�8��*W������n�2ĭ��辶"�V]ۯM<ՅylX�3�o��ge��5[�]��)��[��.s9S���کl�����\C��)Hm|Z�*Ĳ_���r@9�[V��ޜ�yӭ�[��T�[E+kUm�Z%e�U��X,���FU+�,��Պ�V��P�������ڥl����֌��5D*֩Z��mkA+J��(�l�PZ6U+DF�6�R�TZ�����F����"%-e���+lXT����V�Z��()m�KcZ���H�+e[,R֭aj,FьJ���iTb��Kkce��ʖ�m�(��aD%U��R�1`�V[eP��J)Eh�(#hЭ6���m�Z!�Z6Օ�-X�[Y[[FUK
�QB�b�ml-��Z�"�j��U���[-��R�V��EYZ�lH�ՑUE� �X�[h�R�jX�6��V����mZ�+$��[B�UYU��YR-�-h�[*4��
V�R�h�*V���j���m��V��ѭ
*�U�
V[*%��Z���"(VThլD��Z6ւȕ��YB���"�klKJ%Q��(�R�TVX[Am�Y*PTkEDB���F,P+YYEm���kE�j#�V����k.����7QT��>�w�ER(�;�����n�T���"��*�V����ahyr���Q����Vqn��:����� =�ʼ�n���wL��B���]Oݒ�NV�����ݮr�Y�n�'݂1r������x�n�Ck'�x�Q/3��U���%:���^C�� ޝi���o����f�U��֭��-�⛾��fr����b����^��lO$<���F!�tzÁ\wFܑ��v�R}��śښ���c���8g[�Ǉ`�����ґ�K�{��vǡ<������=V�L��sC���
�XU�V��C|��X<i��v��m޽����s�MĎ������ԾV�\��~vh2T�zVg.�\^Mm�O��)-�^wK��S:��Q�dO=�T�2�y��귪[��ӓ_n�z2R���|[ViOv ޹���o���o�/����Op{�/r׋o�}1[먣~�8#���M[��V�t���h l]z�e��8�ڜ���#��.�oR񾱖�RΩ�a8�.�������eKv�Äϗ��Z���%�o{"4�ư�d�n_-�㌾we�F�E)&d��ݛ�ᥚ�G��
�T�P�\�Q-�R���R�t�����Ộ/8���d��#�]�8)���]1�Ѱ��h�Xˬ}�A�Bb���썷��t�'�s#�<�ܥ��}kс�be�0կM�C��͍�k�d�ֻi@I�r�9OU)[�~wK7wè�L����o_'Ka�W]s٘�m%�1)���(y�unk�)]�d�������N�0g,�����-��6�߯��c[/�����*�w�Z�@���nbz�p�5��˷4�Û2z�����Ox���hTUj�5n�д]�Z���;�#�$����;㙀�=.�����#�+Q�ǢLg��Ln�������r�)��+c��������GTqy���g#�xk������|�5�ԥ�At��.)��9g�͎����.OdƯ!�.�N߀�<���c��)�{��A��C9ײ:��3πR�Z��l������ե���j=n���o^��ЦЍw!��B0jB+�]K�S_��������*�U$��)q��H�bJ��Yk��_s�Ȯ��f?PpK�]���s��q;�������t�V����F�Q�kQ�GX�F]�3(&6��W
�Ueݎ;��<=�z�︷W���~oɭ�yߧ��6.�l��	닧��D�����,�{������/Wxu0�>�O�Z�F<c�Q-�p��iG�Cn�k��w�ۻ�N;�u5 �6B7�|�;{Z��T�{����+R��Ҹ��t�x��d������?S�G�bUЧ�|��y��zw;~*�A}�e�Ϩ9{�9/�����C��9ѱ��C�sX�)���o��_�y�R�
>��M1-̎�x����fPyG7�6�(��\M;<�d^/;/q��Υ�Wt9=�[���ԔT���s���5n����'��g�.�I�ff�Ժ�PO��YY��P��ص&G�>̩�I�{o��X1�^�����~�͘���IV�n�r���	N��f����Iu|��uNk�n��['���Z������a�-|��*l�g*GT$�J9�8|g漖���uV�^�s�Gۺ���V�c^y�$ь���/������{�moQ������
�;����5i[ne����ep'�	��q��%ebƑĥ7��͕8�ix-$��yGo&��s�@�z�Gqr�_}�}_<q�=ezs�#����?g�F/&�����;oty��}����=�Jx��ԖjkS'ԣ���WKzJ=�G�9��}���.^\��(v�ԣ�=ص"njOd�����]b:�ZO��.\ʠ�ܧ�����{�^pS}\����pKp[�=p�G��kCa���9��ewA����^�ٯ�g)RWN۳c�4Iey�<�+i.�����-�콱��=�z���|�𜥎dvPAׇId�~^Y޷�r_�1=��|���.��Z�^{���,��q��L��F��{��d�9��m�Iw�j�L�w]���x��N'~�۾���߅1�+����5���������^�B=kc�zkʞ�X���·NnGB[��8����j��ķ18E��]���1`��u���z�a%�A9�9��m	k)	�F��y:���󏯿|E�B�ѳ�v=�Kx�?��㓲S�`:Y �=����3_]E�8�N�ARÕ���2�a����q�����)s*��p�<�\��^LIc��ut��\�\뤒��%�,c�y��#���O���3f�����ǍȻ'b���5��ʞv����r�۽c�Fc��:��p�Ŵ���]���:��)�V(�}`E[^�Fm�K�w{`�k<n���oz�ڙ96}(�8�ܧ�ԭ�Eb�V\^y���f<~��=�s=z��쥽1o��s�.��{�5��+����j��^ͼf�o�K��.~9q�oU]��[�T[~t�vE�7�����ӱ�8-�ܱMl͵����-Q��E�	ë=.���[W�ޢ��y?T���o�t[���+����3"��~�\��u�/ý|g�E`���@���mǣ�=畹[������ٯ�9��>ڽz<&$<���b�G�8*`ׄE]白����x%rj��)NLU8g_�Ӻ6;���y�Q=������sn�]�+'t�.nT�-ΌD��<��԰���S;R�zǯ*��X���෻�(a��T?�ܭ���9������o{�Q���&�x���<�	[�@��IJ�ޅV���ǔV�H8�ڞ�<����G������]��T/]�#��-��z�#9F��ʔ�߷�\y��5о�S�ȸ���ꪯ���A&�I>w��\(�^l>�5}����z_+p.�,r�ٞg�o8���ܞ����T�ׂ��'�y��{�3�kQ:Ȟ{&I�w�x��-��^�ޑ��>EJx'��s�ѥ=�v ޹�+���׾+Ot]�CAVv͏/��n�J����}2����
//>�l�mt�K��d��n�\��w�>*ۦ^s��4�<�5���G����d��8q��R�k�=��*w}�Ks#ʡ=ΆS�t`���r�8�u�0��h�FÉε�#��M����n_�%���z'7��u��I��z���A�Ҝ�8]L�qb�N���*�.��k;�ɳ/��VU2�[�/E�%-��QU:��p�:HY\�r4�o�;_v����ӑ[h�u�B���hUה�B���X���C���_9�p���O��kQ%<}o���Yo�ߓ�#�-WS;o��LV������:FI�=7���ި�J��.��x^�ø�`�@�Z����H�]�m�,rcc4�c���]�/a�Z�tf�[V�n�+-�ײ��T���n�|����:g0v���XRE-��J��4����2IC�=��-�u�F�n��S�5��8�>;����_i�
��G� =㝗����{أ?S�0p֤�;޺�/��mN{aH\�RZ�Rr0�Hp1�Tf�s�4!'�����kc��Fi2�U�13��AB�׭��b\����D�6�P	d��f#�{��s�I&���dΕ����PZL,�w����7���;C��YwHS�X�z���T���Q	�|�|Y��1p��&U��ۀ}�$*w�6�F�Pr�/��]s9@��(�#�p��ݙ��40��x�PgW	"�K~lK��BFE�S��E�%�D��8nG��/,��a����َ���|e|�*�P��x�A����T�GV�0]G��z�k<+�x���y��˘�O_�ֶ�s�i�2K��z����"_���� �P'x��5:OB�uȳkv�jJz�{5�w���E����� o>���M����1jm��@ʥ<@��Z�y	��! �w�af���
��q#��%�̤��馾�zs�=0�lˁ�q.���p�Һ�d�1�7��y"�&�w���v����|P`�n[��d\P�M��9H��~��i�+Ðśt3�\��Ѹ�4=�Y��1�㬊w^aEn�b;Gq�Z�_?�WW�d�`�64���D�F��%ek��˱>�7�;��򏫹^V(Qu��,�Ьy�6d8����-�'6�Y��l�s�3�ab�ww�J��W�W�P��msg/���c�:�'Y0��	���%�,e���}�d���u=w(���2��t��s�-��;���|4�K?��4�N������g�~��xp��ZR�8�Z-b���fyQ��g �QWB� _y�-:�����]J��r/(�d]�� u��܂�F��I����eT����[����,�^� O��C���\�u��R]�<gz)0o��&�no;�jS�Hm��^�VB��gFS�l���]�����(p�t��ۏc�}{�)m�$�n��A	�`��	5p�U�u<n?]և�5���dW]�Z��g����U�Cũt����v��]a{�\�G�O��.z� ��8��N��w��i�FC�锶�p���*�#�γh{o·��8H���;�TW`�KGgbv��(������<[�q�Ià�N�'!�z�C9&��z$X��ps:>���L&/e)�;�u����֝����L�
��]=( �M$Rg����%@���j�j�ի��r�����W����~�g�vșO�	�9���/ �'x5���;��u3�	��~hW�+��9���������v��T�d�-����rط�O:.�vS͖�.��O6<�N��Yۓ��  ���o���*��ˮ�#�a�|�����琹��!��c�y?D��F�Ȭ��o�{$}���L���F������d���y����y�{?U�ds��gC���)��]k]�u/3zd�|��g�l>4.��B���5ޛ.��v�^_��|\2�X�9��y�=��N�|�яk�-�T$2w�?@�ށ-� �-�;
8]{۞�����]�@�'�w���kg�"���r|T�B΅�k�r�sBs���k����~G{c¬�6j��.�|{b'SԦ� 1THTj!�	ٔ{M剖��3�������w{U�35�j�[�ǦG�+2��D��<,8]�+ωS�h�"H�4��wЩ��_e�Av��Mu��<Cp�K"�6i��YDWk���0��v:d�f�����-Y����/�z�Lq3��m?
���=�`<1�s�^�fA-yٔ%U�h��9W[��c'>��e"�[��4�h�J'��|Վ�2��4���>8��������Z�b����}��s�d��YPZ���J�|NW~��K�ñ��.~ɮ��?nѳܟX*�o�[×i+���.�77�.�|W^�F���R��r[ ����E�2�s��¹�v���Y�X�cj�o��������	un�w^��2;:������}_}UA����fo�}���k�ӂ��;o$�a�e��1�,ؙ�eBq�*/2Ds]Wa�R�����x�9�g�M���.����}��FQ���R� �IZe"���^*�|�fr�);�ǭ�8r��F ���`짖���Y]��]l����<�m�mm��&	�:F.�}���/�U�F���E�0��yNC����"]v��`��ɦ�#���7I/��\܀�5��N{���'������8.��j]�&�����osє�4=\�D�	�Ķ���7S\X�j�| w����]�1����N�-�ҰՇ�>D
~wf�t�L�j��At9���.�K��^k���Gd}�س���{�.��y���V8K�z/���o�t*/��B�l�ue����SY�|%)�
�����S�Z�$�#S�n]&%��'��0_�2�쩶B�̔x�2�����Y�{^���s*�>yGLKf8z?r����j�b��at`��q��fPp�=�����ۑ�K����f�{]*?��'.�vI]���E�u�J��H�q���y��.��O5�a���zﻩ�B�o���0mg#yK.۽�Z��{7wq۴��cLr����r�Jt�y�iX^�J�W���-�J�n��/k�$c˕�X��h����C��b�b�l��_~I����$��ݭ{�W^d�i(!�5����t�Q�Ms%������78��vML�5D�*�cFԪ�t��iS���y�G<�aܹ��Oe�m<�
�3�*�n����\��s�kFp;���+�Rc��ʧ��7yކ�;+�N�zY}��pӎ��m�f��k3y�F,��T�'Tk+����n�����{�.��#8�&�Z�C��]�=Mwp.�M���u$�dV]4���=]@�t�Ӏׂ�^ٳ��b&�s[�&��ud��94������UL�qj�mK�Q���RY$6ѺݶXgi���e��gx�k�6�/c���sn����˼:O|��,|WtC_	M�4a����aS�����ַ>Έ�h�h���dr�C�B;�h�v�i�W��+��2�t\����/p��W��k��g�8��G72Aͮ���3}l�Ї(�u*1���Tvn�|J@�;0�����x�C7OxB(�@}qM/v���[\P�r��<����/x��XK�n��-o}�8ɶ�۲R���̴��,�A�o���Gb��>N���� �����Ĝ��u����.���f���͕{��FT��%>|B��Vd9ھZk�<�WR�Vcۏ=�E4<@գ63�C��(mЗ}mEo�͡s�m[����A�E~3��c^�[hR�ޘ�`�����g6��vZ|��|����t�a%�p������)�H7tw*Q�5�.�Q|F��V�:�ws�5ݡJ�9���H�lL��+vJ��ײG�>G�b|�׏vƄ����X��Ia��$Z��5��o�J�j�ۦJ���;�"n�u��L�ˣ{k8������Gq���$��ڽ���d!�j��4��S�T��g�*��/Ϻ�u����^�|r��r]'�ғ��.-��e�|�ţ$G]���(�v���9�4�N�u�ծ�+��<�,�&��Ż��/�J��wT�&���������'��n&�/ᷠ��.5[{f�[Y�*�����[�)��'Md�z���1�c쭽��ձ
{ R�J;���ʭ�Bs�ǹ�!$7��׌�K���p}�K��>Ë���kO#�3w������Y��{��{:�=�2�/B�t�ԥA�I�hF����-�Zw��rr ��]d;=��L����R����1��	���S0�.�fb���?�����B!�.�] ���&ݥS0��:��H�o���{�z�c]6�q]x�xĹ`M�d�ol������s�{�9��%�uv�i����J)�C��9�%q�Zf���KE�Nb���$�'0�$�E
�JT���J�b�cmF*Ū�YFB�� Զ6Ъ5YZ�؅KeR� �l+
ђī�"�1B����P����Qh���-�[,�cU�P-,*�VTDP�V)iER����J�mc5Um-�$RTPDVЬ����Qm��"�µl��(�PmeB��QPiUX�m�K[U�j�R�hZ��*�������*�ѫT���((R�YR�R�J"V��R�ګ��D��Z�T��j��*��DX�X(�U �ڂ�m,QDU�-"´Ab�,YIX)hҢ�FЪ��-���Ԡ��"(����Z�b"�����-�"UT�kVj
���Q��X-J,QFF )Y*%J��VJ���A(���Y��hԣIU�����DQXQ
����-���V����ׅ��៯�[ڋ�e�β����2e�V�����V\·uuH�8��'��3�2o��\����;��� �\魓#�O���c�>�^��nw�=J�;�̢M��+�Nf:�<q��ڻļn��c{B[����={�b}7�J�~�xAc-e�n�����`J{��a��G#�L�sF��X��W�׷��L����������o�� Wx��؜"Q���ZH��<ߖ�V����|��>ǖ��=��Rו嶬�Vyڿe!���ia�)LLL7{a�=�=���Q�N�V�B�~8l^�G{�]��~��l �6#�~;�W�k��vIJ�j��^]��LR��u�r0�����aѡB���pV������+����"�'�x�������s�p"r�]]=�C���aʧ8o�,�9���kV]���]o�c5�U,��pzgrqc��fm��׽���}On $N�و��Ze�]��l�I[�����$���{Mw���'�_�T�\%�?6$K�$uE�S���&g�M�wv2o�o�?yG�9q-�٨���MP��P2��xD�v�m������f�~����{{:�G^	B����š;}heq޽���7������,�-� �OU��֏rغ˚&ґ>��#���@x!b
��̙�l�{޽Ӱ^z&�qP�7���ӯmT��w8*��ќ�|��wT��\éYK!��_K9C0V��{�ֻ1�;Y���/�k����Xɞ����z�
$hR��� 7������}�+���jm��Ɯ�>��_�Y"��H���姆��碪��KD 1��ǞG�t\��� �㕐����>t3�5�u�	�\ӣ�K���v�r���ވ�H�srݧ:+�ӱ�,'I'�&P�7۰dZ��eQA�.�ɔ�{Ճ��`�Ҽ}5ME�Ogqy�ݛ�t��dO��'�"Yϗ�
M*�E���Ǎ���$�0@b2U�"F�6'����gm	����D7=�N�����-~Y,�
E������(=�J8�n���:k��} ������<����^��t��^��^��C]����-7�5����s}���:k��i�w�`��c��}�&���������>Z6�=��G`
qɯ�{�%'c�( �}/�yTX�[G��H�k�\\v5�ӵ��*�c>e
V�gjzܻ�z���sq�/��R�J%���1/P٫�b�H�k���x�=�ˍè�U�y�4z��[����勭�����c�O�^�{w��'ϖ�q�r[���Dt.Րwa�[�4d�̃�7�齇�#Π�gF�[2a	�j�㷊Ao�����b��k��q�lg*
���,�b��X�"H7��Д�ӟ^��_U}�ڣM��q�#�K��Z.��N����yh.�WX^�5׀݋��jGj��P��k{S��˻y�w����z�~U%����ܗI`�R�X3č���M�e�ƴ����Iy�3�s�R��'y��{�ɞq>2�&����쀊�e�ÅN�i~���$��cd�e4<�����$���� >��6;a>4#.d�ĐX p��`�/l�����K�jj�,2��L�|;Kv��+�o�W�<�[�s�<�m���K��z��#,�뵨����:a�A��8���K���9,��5�9�Uɿ;NMT6�Nn�I�ʵή�n�7:���"!n�ɐ��Ĉ�\�H��5�v�\g�\t8Vj�`�=̦�������[1wa�g��R4E�DD%��#���9�k�m�;�~e���J�mm�ˠ�iy��Z�p5݌���2����O�J�ꥲM-�ptb��m�-�zj�ɘؿ�9�]ؐi'�����������f�±}��G[K�H�uP�L�m��V�Fm�T�u�ټ�J��ۙ�lJ���<��kΰvKG�J����(p��}=i���O��������$4�g{��-�񴓔�^�k���ynΎ�#|$�f�U�P0Y�n\8y�cev�u��[}]�Je$�6��oWa��c�>��������]��7l͇�o�VbS(���A�NC�����#$�"�J��K�o2B{�{�������^�#��r�5�Ժ�s���t�d�8�[.,�{�+��������J,�z���uH���>�Y�,w۽���v%�
NW�%>�ɀ���]��V�(ϱMw�(z,�aR(�����U��\j9+Y��N�sXA�e+�s\{���:c�*��5���h�;�UM�ӣI_���<2����=�>aɳ���k��<�v^����9�2?S�YNt�Ք�\m��L\p�ͣrD��a:����s���b���:4*,�gˇ��)h�Σ~��'�X�2T����B�0��X�ƈC\oR.�M1�^>�yW��yM��eN� �g<�=�I�\6���춐C�m��rf���A�GH��ԕy�HV������5��;�E��w<pA��4rK\��}6%����«�.�R�"�K"V|�C�阑��+UμX8���'�o�k��7���e���l����N��dp���5����z�p�k�*���n��z	s��>�I�l�0�ܙ���Cͪ��qތs9�].��̸=����;U�.�mlͳ2�1qc�Z7���%�5�_WR�9�g+s����qW+ y������=���^�1���8-�s.���6h/��>��4X�<ɒu�\�s:�fv���^n�r��g�������ߦ��3~�3"D^#D{	�!gi.����᷎��ft���Z>%�O����u��K��0_�2�쩶{��z���2M8���r��9�}��8jR��vl�7�8�=tO5L�.�`�X~h8��aŏ���T���s�,���C�A8�֭���ס����'*�����s���-{h-+w�z�y��z=K���Ӱ+E���\��40����)`_��]FqK�>�}�9�o�����1?o��A<��3�U�hCO11F���6�]���o��s�%��l���k@�w �=����qj���d(H�7��u����+�m�߆-�5�'9K���kA���}�Wgދ�δ4^�LKK���o<�ܶ��\��jis.��S�v�g��C3��bey�ãh8_�߆_?� y��Pǰ�6�Kj�'�><��6�м���sYX��w�8�VA���U�F�X���i���U���1�y��yT���n �A̽�S�֊HccwO·i_
(1��$Ჴ����W�j�^k�2K��u��ŕ"�|� n���J��:�!ú�u#%E��x�\�79���zc�/�%�]�"�/eB"r���{��̅�\P:���jKC5e[�d�������>��x�8$�zߘ���DH��X�����-���7'���ߘu�l>5�*@�`�:�%�"�K����l���f���mQ�ĭ�X�����z�ۉ��񨧰�'�a��\ 	�tD��e�Kc�R�=3cs<�=U1Z�|�bf�v�g��֮���8=;ή)���arD@Q�8B�9��܉��;w5M��(��l�� �Z�q��տ?]p���ݭ���9�Sm�ʛ`As�F��Ӽ�ٴ�Rz�L %P�1ρ=3��!���:|�gCSdv�Blׇ4��R�`X�UV�.�z����m����0�~�~C3�j�8b�2�Oz�q��t�tT͉^�[1GZ����]"J��c�ד[HJ�aB�f�<X��d��te�8��q�'��K���]C� +(:�C�nGW���D��,��#�U*�B��#iy����
_V�A����ԥX�������'_�#i�Wft��'Y��E$Yvd�W>�N��>|�{C~?�Mk�i�����K�oO4��R���ƳmM��ν�c��J�������o��]��d�^�)��xP�˥]8s���w��s����֣�۲�I�z|�����<�F@�s�kQ>�R{nM���!�NEY̠��`�֨���4�y)4�]b>�}��.�K���[���K�r�K�շ�Pe-�Oz3ڹ��"�������#��Ih�O�vku=]fVS�Y�u�7��϶u��zOtnw���0�����ܽ��8r��q�	ta2)�����T�ޥ
w3+w��ar���˛V[I,����]v��Vo�D؞6��]U�����.���i��1���L�G=x���8X��V��!V�Y�>%a��sĉ.�S=�/�&κz�/	�r���qeM��'.��~���GM:8@�V���q3�(?|�s�.�t��k_xp�(��|<���y.�U�}k��MFr�x�r�	@�Vu����Щ��M�W	ẵwO�c(v�&�XE{�|����ʜ�*m��*ŗ0��ٹ7�����"�:E�P
�e�u̜v�YǢ��z�=�:��T�pپ��6.v[��Գ���n�{<*�u���hQ�^���f��N���\��3a�/�������\+�GH��\���[���{�i��=79!��o�}O1��)�;,Ea��M������~�{���ΣVvz�VM�`���vԱ�U߃����m�Y{ٶ��{�8�$ExkE�!.�Ĉ�z�"F��5�v�\gsoD��/B���:ZY�/O���L]K^�~�U���"���wM�s�����9�s�jV�n�Y�Ylu�3і\(�ˁ�tr:��΅��!/.���;E��}{�T����a���y��������@r����v*�������<�Q���:i��;w�l绖����L�S��<e	�3	��_ń*��֪=�嗻ln��}�,��Q���l^K�n��6;VQ�'|3��dv:qA���9c�.h��۫y	寚�8Jx�+[T|�Û�cw����ؔ2/h��z�j�<��o�����5�qY�F���X�x ���"�����dh�}��0gd{}�B=�z&<��mf��ȞUĮ�fr�����4n�o���N�p��<*����O�	����\��[aД-���y�����S��nO����(~¿��r��'�as@T��o�q��C{ܯ��7&��/�lm��W��y��׏����`"uֹ��8�[y�53;&��5w�g�'�&Or8�BX����쟑r �rd����ھ����l����޾tg\�����N��wwIMQ��5��|����ۓ�X]z���Tпs�pb?z#��u�q����A��VO{5�w���V�* w�0�ӒC�\IGJ(d	�a�[�����$É�g<�*|=Q&j/o)H�+�Ŝ���vfT�F#���6��:I��݃CH�^z�2)��j�dB�����=������T�
�$E��"S��<�6%]f��>������	Xߘ�x�yk��'�4^��c,���`�Tl�U���tyA-R����	��d,��owt�v��
�>~��W�]dmLdk�U�N���H��j s��U�����
p�j^-iA������0c�j�wQ陔�?Hxl0_�.ɶz�xC�ڙm��JH)���,^9�^U�4mr����dR���284�4s�4d�9�������<�C�2c�Ǿ�
�є��U-t�S����u�$χ4�)�eT��d�ؚ���\�����G����>�F�Ӑ��5���̶��>��Y�))`Oqc�ڮ���=�/�Q�mP:�ucq�勛����ޯ�s���ze��z؆uc��ny(���K|SbͧݖD��}���^$�G{����*M�L3\�g�w��V�LTI�ض��xn�p[�C�PZ�L�e䊝��|Y�n��[OZ����K{(�����^�C�R~�x�S��N$u#E֡xD�B��	Jl�nM���o&%Ϟ:Mrw������/_����|��G)j���!B���9�9��p�pP�{�b���7��%�޴?W��D���������9Q�Bߧ=�����)�p��Y��l�����<��^��w(g��C2�ؔ�tn,�{�N�"��9�LG��=��^oMǪ�ĺKY�J ��T�/-,ׇO���8�s�T@8b��MF����\����wHT��a��<f���t�����^ >�D�׻d(���]�b�p��S[o��sp��� }��j٦��7D�>	��y!7�߼H�Ig�v�S���������g��B���{Sԙ��C>����p��D� /+�"Oӭ�W�os����'!�����K�v�/�ǰ�/�v.W�F_��F�!��i�^�TѼ��8��y�0�����~�*v:'���5�/lR2���b�9��Ͷ2g��W���-��ꔳ7�nܧ�4���	����V9.\�A���oS0Ov���8�c����>d���Uv��>�R������q-��CL��Knj�r�rdǮݜj:z�C��3�lO���j�.݊7�=�����;1�vu�����Q`찄�i���݋)ɬ������1��T\ν�\�7ŵ	۶=�����|nA�n�Ph��8���n5�q���������J��R��KO��8l��HU����+�c�d��B�6
Y�!�ON�(X�/�,l���y����5�
��w�q��]nʋ��������.�R�\��++lu�U�K�إ�r≖GB���u�� �yD�b�}�A�>��1U�/ѣ,����v�(�����3E�Ww�V����� ���᧬��Y��Ǉ�i�
����8:��Н��)�jB�/���=�d#�X��mm�Vd�α�&�l�n����Wu�nEׯDbnJΓ�s;zw�,T�<�N�,pf��;z��3���֣�l3��֢Z�Z���ky{�oE�L�[���� �w��ZͰF%���v��2�gd
j�}aǶCp��l~�7�u1���Ht�L���(Р��Xp�kSG ��,�� :�:To�g��h�p�S�3��3"Ĉ�d=
ב�T$Q�˹)��H�?Y��.t!��&v�;g��(E�9Gwp����j�5x)c:r�\	j�A�J��{��uS�]�1�AV�HQ�ʆ_T��p�7K'��,�%��P!o�RU�qN�dҋ¤����|���&�8���ӡA)>^��a�88�#�9�F�%w�d)��+�����}�F��D��=2�E+��ϧf%3m����ݴZ�D����wYN�V	}HԖSH1zl���W��ˊ���bӜ���<ۋ5;�`˚4��gX����<�sd�%Q�
�4b�������s�&�/8Ǽ�����^�ԫ�\ p���s�Q{:la	[��.�K���J�d�5ڒ �Z��N�t����}�P��|������Z���8PB��T�x:��bS�M�Nȋi��kh>Ώ�ۭ������_�ɨ���i������s��&�f�>� �:+w�]Ԋ��B�]��7�\x���sGM7ʉ}�rc���U���MQz�Hײ]>��gK5E)���p�Q3�YE��/:k�c��11�S4��V�촧 �\�.c�I�`�9��#����.r�����ƛB���j�1���_b���M���{_,,�5�V���z~
�h�Vm��\�qgs��@��������j�r�r0e[���v�ui}�V�Nu'�JznE��f"C�W&h�]�"���a��i����nd] �E�ގW'Asu_��Qh�=ꏮ9�����2OK���Ӝ�� �}@6Ȱ��F�lX,Am*,P��#�QQ-�J�*E%`T��Ң�X�T��U""���(��U+Eb���E��)R��BQ��eB�V�Z%X���TA���Z(�"���b�(ZX2Ң%eb���Q���%�9��a�
ZV�[p�"a�`##��5F.U`b�*)PU[j��QTQV*+�UJʩZ�Q�1Ra*#Z�YmR(��%
*�����1PDT�h*�X+��1��F,X�1��UX��Z��ʁF*�A`&AE��*F"����
EX�+iF��F(#j���(-d���T�
)+QTIF�EQE"�2���*@R�Tf��}y��M���ƿ}��j:/n���n�|צ�y_���.ٝP�3,A���jҀͲ��6��C�hv̩�C�s�s�� ~�\]�6{`�5��P���d��4&�sN�e����k����eoviQ��XN$mB0���!/a>�R�݃ zՆs
And�}��Y���"��&y��RR�*�C��lo ���]"N�c��Ml)eE3�3����^ë�kz41>�&t����t1�[A�0�<���R�!�BY�OVns�k٣Tmquv����Rsܒ��}��RR�6��=uO��� Z�]�TY㆚U�rIҏ��c��֛y�"���>��͉�tz�����qY����=�V��A���U�݄=yy	�v�3]��.�9�+�T�������}���]l,A��Kd�l�a(��v���}�܈�M#(W�3�N�g<��&�q��b+�l!�����u�+�[�w�Jv�������;��u��b��ŦM�x�(�W�)}�
rS����N^�LR�lY�R1�9xm���W��EוIfD���q�ZZ=fP<��5y��~u�m�e-��Ϯ1��;�n���px5o�ZFv����`��UP7��
�:�\����)-��x��:.��pf�i��h3\0���Β���1`|u��9����&�H�4:�Z����-�Q���Vƌ�䷊51�y���Hh��N���)T��'y��-���� ��Vp*��+Q����ZK��w,��ʫ����n�A;j,"^K�uZ���fY!Ox�
`���]�{�Θ�TUJ��ڵwK�cibnńW����Ǟ�}�y�*i~ݽ#�d[��l�%;�s�_���F�+��4��d���XaE�ͳ�[~z/�m��N���N[-��d�ꃣ[k�����&R�|H�P��t���N�ڗps6�=��M�}�8�i8{L��0ՉfY�ש��#���{M�s�t �K��~��H{�ۭ�~䞀��f�}���P�Ӂ!�A�T�Bж$[t�n0E�ٯ�������D[솠ߑ������3��]'�f�
�=�z뗆��>��Bd؜���Y�=Ik"}�yV��*��L�S���e�급�~��]K�l�s��6��.�1$d�Qֶ����׮�D�v晰׻cR��+�S�=%h����V�!D��c�b�|}�oV�N>���v�����i��]�{=֚�}�rd!�di9-�K<7}�-ׂg<�|]f�ֱ���v�Nk���c
%�څ��=�{75���87T"��R�M�>&�k�t��t�(�RM���4#���ϖ�chh�H��o�t[5t�&�*�<�0�Pz�̬���r���C&k���e:�#�Nì��V�?MA��D1�W���6�mZ>��N��bW x�X>�t�9�^����s
k4Ӵlȳd�;Ue
�,W�o�����Oݽ5�x"����B}�b/9�2?S�X�~���xl�����5瀗˩Q�^/9�L[5>/���J���\<�8�A��o�|0�:�u�V6�>��Xe��	��N+!�-	�wa囤(�5��B��b��DN0w�+��i�#ML��zr��Ǉ�rMO�eAo!lH8��;�HvP2FL���"�xm�,��0�g;'*���ig_W\�A�e8.���=]t���W/�8z���٘2��=4��V�Ҽӑ )��hrs�>oJi<�FXb�Ȟh����g
�� S~�qD�a�,A�pn�M�WFZ�@dI��%���߼�9�h��~Pp��������x3�,(��c$l�nx�i��-o_lQ���\��g�=EDOZ�7���!k�\zքM�\߱E�����1$�7��>�݋ɮkv��][Y�B��Uͦŝ=
PV��x��Ɛt��F��)jf���R�ڔ���=�K�,=�汽�dc+}���}�;.t��.OO%��`ϧx#VӺ�L̥��C�~��2�\�l
�l�g��L]o�v �O<t��B�>����W!ؽj��$sT�����at`��2��+�k���Q3�QD���s\,��g;�P��'�u���nˊ���dsN���U��u����m�~|����8]L��*���K�V���c�vf�����X�)��{{ܹ���}'S��u(?��C��y.�ׄd��B���&�)��=��k�z�N��e3�V>�diCD�s ��� ��2��9�G)j���!B�sN2��շ�C����ڜ��W	�6ͳ]e��Vڽ���>}��a��;�����D{��q�����3-eq��r��:"��c-b�{�]������j������(��7�Z#��]c��f����T�©A�#���?��\�x+��P՗��Bu�mwtSfC�8�u�\+Γ�ۈ��t(w�	�\� վ!�W4Â���We�w���K\�9���샟Ǜ<�j��ޠ���F�n��ۧ�'�T,�W@��G��Y+Y�=���f4r�KW:}�ӡ�}b>�8�>\W�O��w�ی9`fg>�Z�;�kR2�u��9�ŉ΁�2.�q]�L[Z�Vn\�6�.��9����>3�zYA�amD.������(�%��N:�+c�J:�yNW_Pʟ!ݻ=яnɶ��Z}QY�>�{n&�Ƣ��Ȑ�>@�^'�T,��=���]o�>rnƖj���X�+�8þ��TW^����ײf�dr:�C�"9[�lr��x�W������B0���z�� �|���=�>��B��ݭ���9�m���=���mkS������曆� ����fr�H�7�a�|�gYsXGX���R9�+b%S4T��ߵlĻ
�2�A�8P�-h�$�	�@ش.�S��v�q� Y냱K6w��e*������hʦ�,�e9u�`�I=	���eE3�NS�V�[�ϛ�a�a��ݒm� s�t9�[B���u72��"��9~�9�'�������r��}�k[��C�����R�N�*� O �� 1�N�֍����53Z3B����>��a?+�[B�w�)���=~�.�:X����b�=�"_�믰0����[g̺i�:�x[ϔմ�{;D�^E~�S��]������f�����0re�#�gv���M��`���x�xޅiI��uŕ��/"��R�[)�l���#R���t�E!�H�{k�ε�3-v+�*[�i4������{�c�^��9��#o*�Bòxt�g��Fv9�]��U#m*���x�m���"�#"�1T��A,f��ta2)�:ӡo��J�;���^go��eZ\�����F3��;Jƭ�tV�i�~�l{��Z��0X^���P�9^Y;�	}9������y�����.q�G3Ч��U%�2�b�v�C�y���>��4�)�?f�Ƨ]����!s&��p$r{A�ro�>��h:^v��+�
�<��e��~P4�$��2U+Dϩ�ptVD{3��v�E����{I�.��3{S�!	E�� �-�E&n���<V񓃴�;b� �ȞW�}S=�}]���@����b|��N�C���S�t
_ƍ �&���c���^�AG�ˣ!Wc�/6}��,�^���(*�n��`�*4h/�#�]%���F
����9�t�Hٜ���e���U)���l�v�1A�th;t��"�"�^�~�]�w��@j1ٹ�z<��s�m�Ip�W�\ v4Y;�����ɿ�����=�~F�Y]�T�; �{˗��J�ϰ�r�,҅�*V��-HбY:L�Yhָ�g�wVj.��q��kn*��k��7�mL�M�n>z�Ɩ6i9��<���5�����h�,Fr�2�{B]���b4:N�>�I�IJ�]]��)��N�t�{'tGC~���j�52�{+��(�0<�=l���#y!^�+)m"S���O.�H����Ɇ�N	�dO�/j��9{ۮ�6�$63�ˡnW��5���Z�r����rm��G�������V`�WR蛻ul�ܶ��n�M{9�`*�7h���E������nЕ�8�x��b�5�����{s�n����(jy�׷�3�]��3�S�U��.x��k8�7�3q�9Y.2�";|}W*B�p�r���OE�t{�(�Z�dJ�h6B�P�s��td��*�u�pSY���9�&�ʯ*�Տ���"�ܢ���2�\e�>
��!9W���9�7j���Ez�K�X)��
���w�EG�����i�	��������.�
=b\���y�r���N�#�.�eNw�w�)v�ogӹ*JY�O[
W������KY����:�)W:��s�a�u�f#���� ��)Q���"�8�*m��~�ޠ��*O��Ԁ��B#��z�g\��yR�Ʋe�T��:�k��t��4#:�FCr�Uj)���o�`���n=B��R�H̑�5o/���z��� �d�당˖5^~�o�ֳϦh������������V���0��P�=�Ⱥ	�i.���|܀�5�>���a3ۙ~�$���fTJdô L�D.���=\���#����<�6&�E��ۨ� =떼���z��r��}/�5l@����ߦ�gp�ٺ�*{�f���'�0��m�Io��Sr+�x���jQV!����f>�+�9���!N?X�t�r)�s�k�B.B	qgU���76��I���l�^3�4`]Km����8��=�38-��0�ߡ����pv��^������?g>z��^ T���ʼ��h��.C��9�̢7:��ҭ^�Vg�u6�W���͋P������	B
�.�7�]=P1X�:��0�V�I"��A�L�R����[̱^��:T߃=NxU2�	����r C��ߗ�[vQ��͙�е]e\皩�&-�7d��*��9u�'����o��i�eL��u�e��xD�u��Y�G��^�w�)Â޹�kY�#h��_9��w uNe�iOr8�]L�Csu<^�wt��h\϶�k%4O�3�'��N���YCBU8^�~R0g��sClc;�V7u�0�P�n*�����J.}�5��9]8e7�.:�Qamb���yԸ��B�K!��X�����v/� t�V�]����WeC��D1��#w$�X���鋪�h�]�!��X��^���d:��u�v��Jz�o���Kcb�{zm�=�t�x��-T���,i�''���tn.9��G���G{|�c=m�N��h�Ӆ�����^I� S-�C�N�<Y��fgYY� ��ܶ��z����;B3=�uc�L?�j,ˤ�8I<=�?0�c�F��S�\�'d;��C���� �GOC���0�$g��:R�x�x��,A����H\��$��}kY66|��$4L*�w��X��/@ho�an��!�`dQ:O(�f�2ݬ򩷛׈��O9����&U�ك˜a�AX��-﹛	�y�6z���g��a���{�S��K�ܝ�B�P���h�j�Ֆ2���v{�}=t�]8�퉓�'u7EѿMy�s�ړ��>{`Ak�L�}B�j�z�7]�]1��1˙\��/8�����R%S>�
ﷺ���XX|��U��qQ^v� ��x�Ib��Ц;�A����?T���
Q��C-x�}�)wv,Șʻ�6���@��]kq�c�{wΙ��Ю���	h��#O����sK�3�$q��L�Q���R���֍�}Ywx*�羆h������ï�<WI�l:���e���z�j�h΄�(��m��f��7�9���gˮP��"��D�9�z]�<�V�D�t��R&l]9��������6=�5�����K@�	v�g�x
���0�m��D�7��<<���]/<�vF��!��V�U�����	�))d���~��Q`S�k��Td{pZ^�ƫZ��^kl��W>��eU���4ȟ]��s���d���v>�6���O8���JN�3���-�Q�3�,��u��]2|���>�~8�ݓ �V���ŕ�;�C�)�$���o�����5��eT]l%��8!#��p�Kp�y.�&}M8���b,N-����Ů�b�K5b�Y�Xg��en�L�_����g��놌�SK^�����A���YiE��������w *��`���!s�M|��jp�;Y�벽�a�HW���#(�-�ߺ�EѾ���`�����O��'>�pU�E�4?I�C��{��`K�ef�/Ɛ�������ï�.}��o.�,c,�|=��=\ _ָ�4=��[�)�q�U����$���b�(a�%�Ci��8����#��U�ѐk\�5���׶Kt�!$Au�����Ư�A�3;r�nC9۹��	���r^ꥬm�d��4,*�\���G�4:�� ѫ!�sSq���6�n�aӦ�M��m�1�-��x\�w�yX�[ɋ�pڻ���駈�M8-�"�$��,2w�nK�.a�,�kMn�$��,fU��;B�'���R\��M~�i~�X$�Ge�6�-g�?}����N��Wz���<R�2,ڙ��K�$�H�v����i
=���I��2]*Y��9X� ʲjs����VZ�G{�Jl, ���o{I�QO��cm_Rxƭ5�������^�y���6�V��;�o�{4f��3s�ؠ�l��ckfi�%�A?��ڞ�_f���тǶ��4�=�)\o ��I�=���ɸy�K���H��	.��G�Y%�K�0�n疎����Vv���\�n>|/�R��=(���F�:���o�6^$���G�s/u�z�y��%���y�JO,p�j=��46vj��
���r��듖���5�ү3(�":bT[0����K�(��s�厮��0Z���C�aZ/ �yݤ'��)M��qu�¸.0��n�N1*�݊�w�@�R{l������.�,=�i��6�-��+�}�`��5[��ժ�l�}���V���A�|�P�In �I���4�r�4��nv.D�q�@�۲{ۯ�n��#iZ�tBRaM���<Z3���������� 1�rQ�A䗳p��A�k��}�ј�����!���SO��@�Xm0�콝H�����q��\A����j�#�K�a��n�ؐFF�kٺ-����4�`��4��k;)mi2jݗ�f鑆>����z�v�+&��)'� ԩ�����ul]�Ǯպ��0�eڕtPY㴋c=�.�����F�����l��hrAx�[q]����Ϋ�-������}t2T����㶨��Mg�m$a���bʭ��evunյWǔ����2�Y�k���n����C]C\FE��C6'5��NW��뾤du�mL=YN�3E3���|�Y�q��Ü�4DU�L�M��պ��˕��)����s�i�4T�
��,�;�wH-o@k�_f�.aJ��v�%�ػX�/up������Ngv�U(�Ʈ��$r&��C^�]�,73��"���Ԧ�y�Y�,^������\%��C�6�jzL�[�gJ׻o%V�T�玖q�on\�1ҧ&l�T��L�NI֛/���d�$lz�ˑ��r7\�O�/�WX̢�\9;�I���������Zj[�5��B�87���nP����[�n� ��#�R�\�2�����١woX8���m���0���}����77b<<�Ah�n&@k�{\{WM�ż��g�Yh}4�7u�ҩL�ފ�e;���|�m�s"�P@�h���
"����|�E"�FEX�K@�DE�"��b��Eb�Ȗ��d�DQ�
��ł�dX�`V"(�QEJ����Q�V,�"��Eb��
�VJ,eh���b*p�L5"�V21Ubŀ�ʭh�b��(�(��
)�elqjD��F,QD��(��UA��	EQ �QDA��PS	D���U�� ��"�($YZ�1J�dYW	D���j�QEQ�*"��jŊ�U*�����TDqe���`��TQTE�iQF1TDUE��Lb�	��E�E�
�Q\%���R�G�*�r(Q�]{�����6)^D�Y��!�r�[�O;$�&jdd"�lҭ�>������!Y�6��y�8�[��9s���H��f�(�~���Ur�+x���X��E�AdO��{v�j%۔��w����zj�?>��ʙd!<��"� �4i�O>y��T�P�i	ޜ���Vg��j9�)vG���z��b�w��70(Th�_tGĺJCj��o���5���x�g.����/y�FT��ˇ٩���:4�:z��[��x�����|칎��.��}���Y@L��C���/�4%��`�z��w�+���Wc���쭙�&�[���L�J����F��k�糹�*���|�QZC0Aٵ�=�\�#Y�������z�ExG�z����G�>����W��xU��Q6�$6*x�m�'�wu��󢑭S]Dΰ8X"~�X�Z���n������a��uĈ�۷�̮��mPR�Uэ�t2���S �u]�pU�����l�>�x�;w� �Ϙ��Sm�O�ѯ�'��ę�z�O�*?U֪��	���x �_�]j�M��xӪQ`�1t�˺4���f��6��f� v+�*wCD4�i��#��`����t6�25N�1�kt:�T�r�7y���p��uk��0-֍�-����&{Z����+@ڎ��E��<�_f��T!�*3��36V��k�m�z$�9α�j��Q�#ME}�9�GU��?Տ8{������&$z�{�Ϧ��O���׾�4��IC���M諔X�o����%��\'/���s0n�wO�e��ڰ
{.5ŵ6�ʣ:�M�íU��v&1F��A��r�n�'B{ϋ��֊�ȎV�t�4���l�^�=�BTxy��^�Y�C`J�������%�t�a�zD���YX�"���4q�T���]�0�����B�=�ȰP��P������NQL}"��ly�S�:Lޞd��u�2�	�ȅ�<s�������9^�Ġ���+�2���q.e��N�~�s������<�s<��=:L�b@2Ddi,C���_e*+~�}ѫ]L$,�AǶəS�
�=���[�2���ڛ3ͪ�o]
eIRf4�)ٓ����;�B�����VUz�¿�m�`���5�ˮ{��~�xl0_/�}�.�6�"��M����
@
{�Z>��Su8�.B�;�9�̢.��d4ڰi�;�Zd���ܻT��t��Y���Ϯ� ��s��
���)�<�X㷔i�X��HmwR,���Ν�����F�Kճ�{��s��G�P+�IR��K�����s��l\�{���Փ�G(sn
�����5��	a���3��yʥ8:�e���i9�n��ғWQW����<.�EA\��#����گD��x�<���;�N����[��I�(W�y��9��VU9`p��pc�1*Ɔ,e�pw{|:��m�ˑ�j�[�Lt,u�3䥒o������s�����7U�w�pΥ�7��x�qof���m6�J�'�h��vb��@CU�`�]�9~z|��Z��na�Lei}=�E�D�������VnF�̆�zħV�Dfb�κ�0z�^i'.�v��<�:�[��+��3!Li7�p'#�T����g�W��e�������j�/�]��T���os�U9��dj��������}�u�LOd�R�i�վ,¯ K�o�����Md�/��fp�)��3=�.��uI���QfZZ6����)��
S�b���$�1�y���k�4>�fYzC�#����$g��:R�l�yzÕ7��}�ᴽw��%ܷX�d�v&+�	S
��%�8��ߧ�3�|Ŷw�.�Q�H7�X7b��}�C�o]�7gK�~�6�햨�k�n �ϱ*&���\�>�yyn�5`��r�X"���������^��!����
W���{V�ؕ��EV�r�ܮ�c9e5z������¡xԘ�w�2��-e+)wt3,�Z\S��gNbt�#�K��%�f���\��;�8���pV�Edz��3c^ǚ3g��ɮ���+Oo'Lx���qݚ��B�.�oO�vOG.Nε��;=��?�{�c��ؚU�ūy{㫯a\�[��9&��l.��O�� ՚�8n�P�yGY\f�.es��A�R��^��T|S�ȯ��;%�J��8��a8�P�/kG���@�g�:;ݰbw�97z%ܽ�R-~�v|X�2e˦���煝��r�#�6��։+���myp�d�%��sw_��'��gNvD�lN1OlwOc0@�K�C��-�6��|��,e�t��u��<�x-��T�/o�!ªUv�6,K/�JY驀z��� ]9^`�<w�B4�WC���^f��fc��W��9�ض�G���\�qۯ'�z�?�
l�P#"����$Gj<��cio8��9���eE`W�on�ţo�'8�{�lϫ��;vL�=]��y���H@sI�o�t�4MyC�Sj�9�����A�cc!�]���Kp�%фȦ�O^�19��L�u(7ҕ�/u��P�2l�k7�y�^J��Θ�9��"�.�^	��}���Ӳgt�E�z~Y�*[7����Y�]���W�Qm�ݨ[���>�;uT��"����G���AJ
��fEJ`pG˓��Z��[S�;�������d�M���;=χSFP��Z�Ĩ��堍��W�y��{�g<I�=��}h0yb�t�����29��u}#���!^g[�+:`��2>s�4���f�y���\!mB�LWd&ɠ�\	�'���w��{�ϦzM|�@�V�>�������
�b�<�[-�P�Ų�|W�2z�@�����`�ؼWzU�ƧlxR\��3�!�+���ĊL�{Ե[�NP�,Nذ�"u�GnN�T��Y\���˰��Mߜ��Y_�ǀ�~0��P��Ѥ�f�<��i��9�nj�V�Kmy�^�S��q�7꿫"y�v�o���wJ��X��A}]�$��M+7ĦAY�rN�s��S�ꓼ�]��켾8g�i�K���C��H���c�;}�mݚ��c��V���&=���A�]t�[`t8����.�	v�'��S�!�A�$��P�.9�U��<����^��i/��b^دMA�G5�ȉ��|��y� �ss{k���;�祘?E^�G�Q��Mn�v�{�[�Y٧�WU�+���=�S^#�bZ�ƛ�rxܙ���\r	��OvxHwX��ڢ��3x諾9𚒣s2�M9��s�z���27jU��B�ѳ�%yn%��W��iy��i'Λ;�萬�y�.��Fq�m�Ư�ڳa���fRS(��!�^�c��$�"�E�h{ή"u�e ϙi�=�,f����ٛ7冔���pf`�qb�q�eՒ�W���%�Cr��8_ݝpe�������*�<�[{}*x�V�E�ן����
׶ʡ*?p�jU��錝�Y�`���u�����@Uʻ�1��Z��[�u��Z�y������m�{|$#��"�.�n<��Ez�u�r��4����jk�STD�ԟ��FW�w�B����B�C�o	ʾ�&W���鬋�w���"�3W�:���o��S�m���B|mf��-T�GX���
N�"���`k8��_�����j�wvs̮��1�7;�U&6# �x�Iu�P��������K,�Ӥi*�XL�\&M��!P��\��lCի>��!�{�K#ABBIBu}~𥶫p���#�ow$%�{��kY\u�nkY,����T�aV�����<������Z�b���u~������ͧ˹�=��?ߣ�b?��j���k�˖��,�����g.���>���������c�(֖خ��}�m�TuA�^�]�]7kz%9jk�]5��L�u	��LC��˶��ӕ:����ܼ��|�16�Y���B��.��Wu4�?m���`c"��t��w��n*z�١ج^{N�����&b��o[k�*�3�&W��;[l�;�V�s�7:�A�~��͙�d�;9���{FȜ]79sځ/P� �p�2�㴂��r�qA��G=ZĻ�Ҩ?L<:����"�y��Z�k�k���{r�� �> �����p�Ϯ�k���^�G2���⦻Y����2�uD�(���2C��qC��t�c������l;�^w	A}6n��M.h3�ǔIp�^r�PP�v��$˸1CT@�
+�5B��������oo^�v����l�))��(ӆ��ĶG%�Y��F�3�f���fH�w�!ihVהÅ�Us�\g�rk�_�%��w ne�~S܎U�c6]��U�I��6��e̋`s�gt��3�9FxΑ�[6+6j�;7��1�xFmN~�ck��>��������a`v������"�b�t�j���|*G@[Q3�+�F2�NOC]�;�������PF�ž�\����r?S�~�/5LC,�Oǻ�d�۩�+횺L����/�_r�5淄"�Ц2J��y[8�n���ݜ��{�[u�;��U+KF���~��So�t���DƤ��R*r:������aW���[���t�����xk��\�sqp�E��S^	d�A(8��^��ӡ^��ϒ�]��������x�6K�pqR�����\*�Ra�:�E�%��I��}�AԺ��n�\��k���\= �-�
��Cz��#����$g��ĄaD�2/:��5y+"���o4ɭrO��h���(y�l���vh<F�=����w�?p]�~�gV~
�)}�jW�����끐�%�b'��;^��G����\��
�QY��ͅ���F��|..7{;\l�O�c���4>b� 0ѮR�Ֆ1۹�j{�}���wq�hy�R�OH}�7�}n�&��s~�lfM� ����@ �ѯS����Y\cS�;�p	�Υ�e�hmF��4i
��4��:���K�D?	꫸)��P$i5���	��{�T�5��1����fzd�z%�\s0��=5�a8��P֌u��z�(ͦJ���5}Z۪�ۼ�@O�t!���[JXg|��M�0@�{·9�+(?���U"�.�VVK�k��s�Mv�qʸS���#�[����Uv�Ρ�7r�i�1u��Rsy���x��ج1���<��t,�#JbnKH����{��������]	L�j���m��5	Oh�7ƺ-�i]:v�Z�m�hwX�<7�y	�=΋/��y�
$��.Ͼ^^��@����(6��0�%,�50]?Td�r��NZńZ˓�LOy��<��Ŷtӡ�e��r/+�4ȑw�+��R_�s�@���j�=�gY#�����u>�fw�UY�^���]2%�L�!����co����-@�Ԗ:d�ko�'��<:���'f������������	\o��c����0�_<.���^�qAR������^ў0���p$m��p�X�7�N�dO?*���{��6����R��S�r�c��1��h9s��4�|w5�q�EZ\/pG^�wC�=�L>�0����7�t�#�HNT낙��*�w���i���7�m,���F�*��O�B j=!1Йb6q�y����#�u�뭠�����%3�r���wE1k2�H^��a���N����t�[�N���Ѯ}�d����0�=N'�c~�i����A/�����U����Q�jv
�]]�P��yep��g����=�N.��H�p%�yܝP��b��bU�]t�V2Y���=Vb��&JwB��M�C��9�:1��n�ۻ��7u6n���,Vu�����V��=��l��K�{�IIQS%&������])��v7ڸZ�rvH��R��L��)�����G꿲'�fa���}2��L
U4D|K���<�>U3-Uv2��碶���#�!�k�]���Ȯ<�it\�1��tk�� uIi��.Yu�.�X�7���K�j�&.�]-�:�X��ޙp=�DlC��H�P綻5�sY}�b�c�I5�N��ܫ���F�h�~u�s� �`k�=l��ww���
���֯�_�u�
�u,^u.���]2���L�r�Cu�&�����[�y�P�%�-�beж�ω�R���D57�Cضڃ4�e�3/��D~p����ݪlBrsv�92�;T����\�����0�g\b�4lc�⬕|*�9�#��]�����뾆�f0��_a�6?p��z��Ld�l�2����FN'���7Qq8��80��y�zf�.k�W	�p�z_���G�F>������d����N�X�*���׊��4��z}'�,Ve+O��6�zá�7������.]��Դ�}��jj��Ϟn��|��ė]hum<6<]��-���2k��f��Ϡ�=X�/vnMQ���
�Ӂ�i��i�l.g���w"��YZ�bKH�1��
ť ��̽���R�&�ѣO��8�.��;�}�ӄ1��ƣ�N�0l�N�_�xٶB��.�|Ig&�%֦��<��o|x�A� [@m�-Q�iG9*%�Z��qF�z]|Ps5����'$�Z&�$��*z���������e��<�̌H�F��P��A�X�t�|8��<�!����&��἟v� ��~�Էtk=��	x�J�[:k+[�&j�t���:�XT���jՇ!�G��N��j��E� #�}��Sݨ�`�̙yl�z�a�;w��~���M�(�;��Z;�>Ì��hP��b�����U�=�X�&�;��gM���Bsm����I1���]
�4=y�Ż�3�+�vL1o6�_��n�yϺC
�X��&p�jdV����DV5Aj�.@^���r�vX�����K��J��۝|����?)=z�O���F��t���.��g`�7��D���M��s[�P�{&�/>��Wj�k�	�Y���#VU`ˠ�:+��SK�d����.�,Z��M������nE��쇶�.��hp�{�H��[�`��̧�-q1e���.@:ok�J� �c��4�U�v{w��Ol�������ZEUc�C~߷<�Ceg��/��UQ�ۦ�ڙ͠4͈�CB�&����ඵ���p\��G��ytEep����a"�|Ow�Պ�9��|��7 M� ����U���{b�,:k�.a�1;���z��=��M�K��kDǇo�E�I��0�����]q��f�n��Z
�h�|�Cz�U�إ���@��ɱj��&q�;��r�o�� u���ژr	�N�^�D+ 0��]�O��7ǫbCf�+�}��fL`��֫qK�R��t�cVj�~�֊�"�[�������ݝzb���ø�GSۗ���ke���ϳSGW\�KjJ2;aEAA[�Ը���2�\�"�4�'#%�m��#Eq�m�;tᢴS�>��n�.��8����Ԡ_U�G��:��n�G�~�1]�4!~�F����oH�V{8��mc�F�������},�p��Ȱ����qxq��>����Xq�&��N��x��qP|�L;��/�5�9�n�r��Z�r�:ƴ��:T�O2G	nWtj�:���r��}��>�i��W+y(x�AF���u$5�:sRC����sTB�=�5[BE:n+-ʚ��]y����]M�{CJ�	�[��9�+U)J@��)�4�4B+sT�v��V�k�.�d�+��5�0i�h�N�2��sH8vc��ǁ���j{)@���u�Cuw2R{c]��cJ���͓�&��:��*�]���..0���{�����]Tq���*YxT����z�[u�|�������A
��S���`�e����Im+UTAQkb,X6�IR���F�X�bDUcP��,�Tf���P�� ���ȡmX��*V*4T-�C��"(�((�֢���DF*#m&1b��FZ�b*��1Ub*"��DQb �D��µA`��QQ"+[V,cR�UU�Z"��"�hQ+TUX�1H���؊�Ԣ��EEF(�UX��F�*�TDR �� �RԲ"1F,E�*�*Ŋ�(�E�m�APDb�1
Ѭ�DTA��h��6�1��AQ`��KP�"((��
"�BҊ"�[B��P�kJ#E��KeA���*�P �h]����1�7O:w5�˔�LF�4-	l�o*y���EE�f�r����m�Y�i����l
�Mt��E�N�0��q��[��_a2���mf��*��T�F��?P��
vЃ˦�����	U��{u�s��)72�2:�M�c��]+dptt/ZZϭ\)Ҕ����ZIf���S��kcS���xB�F �58�n��b��[�q0#a��$���,�u#�NK��;S^Oz,j�y�`�5��;�7�F�Y߄	�ϢLUԱ���:W�t�:�Y
^IE&_n��b��fz��;�zk)�m��T01sS�3ɜ���� Tù&ѵ2<^H_6�d�N�Е�0������[l���
��x;U�B�~��UM��b;[c�2{˪ߔI'3ړ��FP��B���&��2�����L:Yf�9u�L���!��.tz�ȷ���wO	�e<�;>�`1t,\�@狅^}Wtѵ�\�j/p+�o���c+*æ�r@��W���;��)�2C��q�Łhϑ��*���pײ����)�.���7��2}�q)tIT砯_�f:Nx3ՎX.�]��LG��`Y�+<f�u��'f�ӵ��s�z^vf%���M�شʒ�\�oKY�������i��\��8+�YJ\�:�>�2�}�K��,�rK)��E�F�)X�ΦwS���u�\�$�4��a����.z��[ޣw�rv)x����jN�#R��9|/w{4N(u��$��)��	N{Y�oZ�22�\@)��j�j���r�����^@gUyt��}w��`}��s��w ���.5o6���[�+�Z���ɲ��v�ҙگ�^�H]a�m�2�W�Vի�2��	��#[�<���^D�8�Q��q���g�z!�}��_�L_�iq�.��`����.ιC jd�'�/o���՜��|s��ګ��FT��U�z�RY%��	�L!"2�8�͆�31�4��:��ew���dT��hF`�n��i�����Y���U�v9�P�Qj^Q4��'��.X���)��8��/Tσ����1u�י��Wt&�������\RM��%��h��.f:�L�L=��x�9�kX�����y#��+Q�A�u�|�N�ݘ6���	�N��-����疿
̯s!|�=��]�mtf�ڶ���u�z��)���#��� /�
�=��J�?��0_���9^Z�5ʾٗP�Y�ddJ���<pW�`��ՙ���=Q�'�Ao�JvV�[i�۲kRo����U�P���~��$����N�a�mX�Q�� p��>�����,M�ن�\�]w]-��2Ox�j\]\T6Y�3����ݹYNq����c�o�R���za�Sm��� �<�?�4(��k�ʔe*ի�^;Լ���p��z�E�.k��Ty�&�t⢼�/��]�a-(+��1:�y�,!Uߢ�+�9P���k���fzd�v!̋��I���C��K�I��^pǵ.}�L��谉��,Z):JZX�f�a��R�7L���:+(7<4�c}u+�9�᫣����Us�IBxfBkb����^J��Fi�tkۮH7�S �5����P��[��%ٮ�eDCE�:�ܛ#���B��.r�޺�w��n�O�p<[.c�ܷGT�r�	r� z_���[��qcn.r:��5^K��sL�yT:6���0SK-5���R_tN�ʯO	C}-��:�H���G����\p�0v�
]d���r)EK2'4��ݘ�m���G�JN�en�&��.�c�Ai�Z=�i�~f�R�sw��I;��&#>�Ew�)�.k�������\�_���6��{�!uM*�*����w���ϻA<��X�f��ꆗ�����QR��;�S���~+|�P����S��5���l�����f��N崝>�����\;ی5���>K�:U����5���.���e1�����\���u)�ѽ�u*b�3�2��'<|)
�s�=g���҂�\$s��	��)��NU�;�?a�]���{|G^^�dӼ��a��u�Rt�9tH���1߄���J�!~]������L�C��9�4���O�6���E0���oֈ������^���Q�H���7]�8H[�a-�
�&���zޔ�b�R�C�Oz��t�mX���:��B�E����4�8�U�����~~�׍��̜Y:���u�<�3v��J��0(F�]�0�i�PkWz6�sI6B�h!R�!t����w3njr+�y��c�Ӣ&)�th;v��~�)�x�dz���o��o��;ʻ�].��-�:�X��ޙp:���0K=@�x��X�eđ}��.�R�լ��J���](�y�~گ�A4�~}�ȂY��-Ic=�T6��[\����@�E^|F|X����
��ꊊþ���-��[4΁ܶqo���]Sֹpկ|��&%�͌ˠ����X�,!�,�uZ��m�Pf���h�J�E��Z�R޳X]E��fܫ3��0�y�7z�ϫ���zB�l�t��`8�=����e��2�rT7��^�ƨ��y��,��W]��GJp�)��3&]����7r���1Tj���jQ�Q�O�&`/d����{n6��NZ��lN���ncH��IԓIٓ�ea��R��+�WϦJP�c�R�������4llm��yE���[&ަ���U<���f!:�_a�#:)5*�s��9���'j.����#@岟_r3o��Z#���eH��ԱY�̎���!^��]�ܧ�5�l���>��wS���u�V�]��{��q�a}{+a�gM#�&|\(	�̍�S���9W����b��0�2�r[��^V#Mw��JȮ��4[��>GY�b�.�JkX���
Ui�����u-4-?;��b�3�g��_�<�����8aм=ik> �
�R�Թ)V��W�6ۦ5�w�_j<Q��DT�F��j k9L�6
G�YT
�!�WnBg,kw�����)o��2���qߢ�#W,�	��y��+*���K��d׭|�FE�s���i��I8B%x3��Q�\HH�L4��m��}MN�b�i�õBe@;qY�2��<��9ӵ�8
�S�48"xE�ˣ���nx�@<�"����oʠ����ӹ�e�A;� �o%b�%�L�T�]+�]l�ڡ��L1���(�<�$��E�pd1���+�yk��6k˔��t����7H�s���D���髭�A��A�MT�`{U������B��S�|�u x�32X}%�ǚ��e���]s9�w.���!΄ɐ���y�knN�Y��9u�f�;2;�xG���p��à~Xxm3�2�쩌`
?lG�t���m����{�UێLoucBrO���̢-�d4��K����1����:��:�Q�6��z1��3@�x�m�=���f�q1=S�3�IL�M��+�󙎃�3��r��u2�{�Z�ϰ�u��̏ur����@V�T,XW[���f��P�0bR�63��ds��$j��7�F�w����9�wݬ��뵐��;^�xD��*�1��~��N4X�t`d~ W	sJ/��yF������2��#��]<�\�:̈́o��
3�}�d�͚͊�[j�CV0yt���U�h��p1bH��o$f|�6���dVd)����E��m���7(W_�����ɻ�s��V�Էl7�K8:���͒�ۗ�Eװ,��b��~K�I!/��	t�ɏg,�|�4�|�z����F����mQR�����]1[u����yu�׀����2��=x>�!���Yj<ЁB�૚��ݖՃnT��^��B��!�*1Wd�ڻ&��Lʝ��Y'̈)�k���F9t�����'�z�̈́�tX����Pq�GKj56E��Jo~���-h�ׇn���t��R�p�IŢa�Wv����� ���*���6$^����uTb�υ�L)viq��۝��fM����0�N��~����<�v;�	S
��&8�����b�����{�s]�iԹѓ��� Be'��H����~~ӞZ�+2��Ȉ� �}#JO��ٓvfv�\U���d:���C�)�3�2Ֆ2���A��l�e@�㹓ekO|����*�Ov�͗4�Ͷ3*��]L2@�
b<�5u<z���^�>�7ϟILƗ.Q�Y�^�.�u�氎�hM�ӣ�a�8���'`��h�)�Ld�l����k��+�3�LE�Z5a��(tk4�C�C�9��b��zk��p/-�f�-���v����L�m4�e<F.�Ӏ�$�a��]�sj+u�&x�����s�Vи7�H$���˯�Bw>ih�)��n}�d�-Qzo��o{��ټ�0�RR�-K��dh�o4lx��q�/dU�@�� y��m�u�&��(�Ы�dH�����>?|kl\U5���:�ժ� �� z)]���f���!�Y�s�ҳ�O��J�'Ihʬ��w�ݝ#Mu�v�g-�|������];���I�wc[h�*>��S��I*put��J�}Ѿ��odT�-.�gV�V;����d��9ZdV�>ݒsq�!���sxF}Bi|N)`W�on�ʥ�o��{x�,d��˘��m��J&JoS�t���׻Ր���['6u��W�A���<3��>۶��"�뙴��,��8��9�.j�t6��T�ޥ
��̭��d䞃���ւߎ��ߎ��V�Ї=������.�Ԕ����]V;԰zB2�Z x����|��4�|Vǃ3�N�-8�gy�Y]*��.-f_�ρZ�u�<H�|�&��p$r{A�⌘d�k�n�m���~��!$�rg�Y첍_Ǉ���G�"�4����������Ũq�Xեg�B���=���	E��;MFrg�WR�.�J !OI���t��M�~���9�yo}$����a.oH�+Sϲe�:��!0XL�E(�l��9�j\��Ū*4��+�m�(u�����G꼉��ߦ�
˺��u���F���n����Q��$��%�D��S���9�n]������\3���ϙ�<ϙ	�7o���a���fnE�U��U<��q
;��1VBk`u-�N�]�ͮŔ'3Pd�[��:�ҝk5f8����6�UNr�����&��61a�{�c�o��55�y�G�&�e��b}�j<� ݊X�Ny^��x3�5��o�)��ٳqٚИ"C�'bju]g�nď����]��u�o��S,Fr��.R�
v�������mw��p���}@�C^ޒHC:�>\���sroM1�x<�Ws�&�W-�׼�V))�2��N.��4����x:��]*��~-���]>՛U�w+Qti�u͙Қ\�
�J�O�Cb�����)��Wy������5jŷ�Pf�%q�~/V �<��o/vw=Z'϶f���a�J]q9�9WF���C*qR��j��+D,x�<��|���Q���p�r�s�n����(mG�tԫ�ϟLd�l�2��tp��8�ٛYʔ����ʜ��r#k��r�7�t/�q�FU�𐍫W�g�]��}q�^�b�����D_�����f>Ի3���i�Ӥ�G�6`�)�x��	�B���;X�Jt|��z�mr�2�#�M�2Iu8�lw�VEp#�#���>�rH��i���ɇ,F\��W�\m��7x�<�1�i�A�u^w�9���������J�м=%���\+~9���u�Yw?^ӤΖ��Gd˃<�d�tmz�]|��<M�+�`��Ԉ��.9eY�,�Y�g�Ci���'
�=�e�u�N~cB���V���s�D��ʅ��efK
a�i�Om!���Z�ɩ��\��o62�(�{3��W��k5���zK�Y�N� �b0<���jʙ�!�{���,�p�����������h�I:'�i
�J�X��iU�7���t@�̪�]AO�*ۑz�p!���6�vwd���xό�V�A�����wt��9�7�@���hͩ���:��ڣ�����q�^��q0Y�Bz�a�#	�3��	t�A��c��ڼ+yc��\��`�]]~��4�ئ_������1�{n���!Й&7���gnY.Oi����Rգ.Y�;]��r�iۥ���h?L<6/�ʙpvT�����xH�wM��(�3����m�:��\��s���m�tD��d4����<�Qc|�q�R�:�Q�6��ƅ��iNm�crgdi;��~�����{ԬC�K�J����s1��s������̻�e�g]55�}
��m�:n?X< ����w{4>���`�JY&�ʺ7�N���sM3�0�EݛΦ��2��s8-'O�S�9ό��߮��͹���]x�`��s 3��V�`�Ԥ�Z7�S�]>B�7/%��f��(=8��]����|�\4�����L��w��V�2[	ڷ���6�Es�U5�s5��
��� ��ͤy�lv��,��l�iCD/���=s�gJr�z͇��;޸JSػ��t��;6lT��)�N�r��J�PT����d�&�st%˨�@7��5����2�ǔ8���J�+���o�=X�]�ɼ�����}w���.)��s�[O�Fvt�f���E�Y�*�X<��a�]�k@,��NN����y*o6�I��s��o�8ȹ�h��{aλ�*Lc+� ݦ���sغMiufj��U	���*Ĭw|� 9���{z�G �׭]�~A1�̽pL;BGQ�;���\hk$�[n�3[Yt����a�+K�tGL.���;��4j��`=b�T��U��q4�f�b\���f'�۶�Bn�����S���2g�{M��ݼ�U-r�rqsr�%sC}Z)�|!�Ӑ���;�e�[�-]4�dU��ojջ���x���٭FFH������R���
o��T w���V�&q5������.c���s��
�28X�}��kX=.��d�yi6јtz�2�e���}��ˍ&��,c�Ƒ�Wˉ�(&�ګʤE=@I��af�p��[P��m>lZu�I�3rʺRJ=¦|�p�y�Q57gS�l�On���U̓�'�i=չ&IXN�<Yv,Z�&S�n��8|Z�,A�3���v����e&^ՏK��Μ��K��Q+����0sܻ�d�I���2��i����g�;���~�i=�}��8�4g.!�&��X�`(�
%6�g�I�3����DSC]�7O+*j`�Մ�V���:鞑�0Ӊ�C$�h��i_nh5p��lp��b��.���l���Z")�J|��O�Ջ�t7�0^���-g�s���3I��&�/�
]��7%�֧��Gi�:�8;*�Z���x�=Pڊ���m
Wӌ��G��DZ,�7�B��o����®����G?Z�W`޷�pt���'I��nB��CyM�$��֑�E���w��~%�h�v�����fN�$KW���q�b.��)�J��ݘ\�.�w*r�!��&�-�|u�CohI���Nl,̫��pL������<e�-�Bhs���`�O�W9��_a�;S�]h˞ű�=�F���w&-^u(�R������M�۷rS"C�ϕ���Wo����*=��Es��y�A�PU��F:��~�(ƀ��=�tq��ňЯ�����_]^��;�v�I�u��B���Q]J�w#�t��tU����x��s�'JICZ9��[���p
`Q���0T7QeZ�(�5�Lb��e,��5�#
��ݮF��Z�6[P�D����+�X���UX��P�e��TE���YX�1������k(�m��iETU�����""*�6ؖ�F6�T�YF�5-�ZҥUU��mR�F�m��m�����Z�(�-m)U�j�Uh�(�U�֊�j������X��l**��KJ��-(�X��QDm�("T���[IA*Q��X�-�[jT��"�(�DUb�F�ʲڌEU*�+R����Q
�QUHĈ�m�VU�
�b�m�m�DJ�Qm,��X�mV"[aR�B��ijŭ��V�D�AeQ+щKVҨ�V�h�ZQ�R�V���� �F+F�lKem�Q�ZXq+�ѧh�I�9+]uH3je�GF�L;�f�5������pmT���7�k�ƕ��ѕܳ1��Q�rL�s�׭�7�L�~�܈r�:��z�\�:ͣxj������`Z-��5Oi�[����,鱭���x\�^B����7���H�	����uw�7t��K��P||1�������+��[��ˬ��&S��tmPp�9[%�]�c�����c��ps��r��/6�q�B%J4�T�>����o�K|v�f{Yt�m���k2�����LY�/��L0�<>IA2�X�X= ��6S�n���)�=<�1u��;˥�}e�D�����J��8�q�\��H�ߛ�~�" jaS�D��qk�!;l�8�֝���Wg��1�<��J%вzh�����疿
�B�wsfFR���k�|�M����挆�����q�B�P�R��z_ʕt[�`̤�<Ay9���HQ�O��r��)��ps��*�Ov�͗4���c2m��X@t$P����٦�)��{6s�J*xe-��ei��2��5�u�	�\ӣ�a�8���'���C�g��y,�vC�
�k������,Q@�����"U�e
]��t�tk�M�j:�u�J���Ra�`�=�1��S�je�:�;�{�=H҆����.��ۚ�Ʒ�y�*Gj@ݪ��i�V��U�swj���;%[%��	�U�S������~�d�t�N��$H�	xTEЯ_np�*�1�P�ޙ2��wZ1�;YT��D�Й�2͢�߮Hw&̫C�$�|������c���;�,3�>���X����%����������ϻ���)����q�[�_��&��'ōK2�����3�aϩ)d]�Y�w�ڣ9���z�*�@rR���Zu��gK���|���~�~4�5��a����������O����o��]>�τ���ߘUY�\�+���WL'�~���kۻ^i��}�)�>Y����>��V�NQ�ϥ�r�u��z!����7�������3vF�U%%����b4N-��{�$k'�Ȭ<�>���#���Y� �fR�Ш��'¼#<Z��О:���]�������-�+�^S���$C�cF����}I�ĳF��3Z��G��F��s�f�^څ̘��	�^' ���8;�&v�䔩�����S��5��>��i�q��N�'!������:�b6q�[֌Дf�G1�d�I���kj]*n�Kq��rX��N�sǜ�Nea͔�`��;�|�i�af_j���<}s�n��L{k��V����ۖ�g�r��gcފr��ݤ�`vR��'RӶ�6ʙ� ���:�r���V�39C2��\�{u�K[�Lf�SwY.�A�_Z��1d��.�B����tJ���D5u�n#���;�{|Uaˮ&�f�'o�a]dO+�&{��\a��u{�t��'���iU{�����6�B5��5�s'R�C��u+by�v��
�əK=ayJww��͑o�|������$���F
��eM�!�_�ˌ�`9�Ȯ<�it\�06��=����Gy��嶌{^�<�C�(���QxGuM�wj�'Z<g���2�q�+
]~����	Z�g��[�����+�8� �uI$!�I��l7m�wj�5NBZK�"��W�|z,�ΖG�����V3�@�+ψ�0A�PH�A�ж��ӓ^�l���W���:�OU&����zeG�+1)�M����.�|�y�9JX<af�WxM�y��ޢ����M�x����/wVl<ߖJz��U�UѺ}2P�{�o_�y1��{ݵ�ܝ��E��!�v��ِN�}�P��®��u��錜�g��M����s���k�-��\ܧҶc�;�Ow�4X	d(��WW˺�=�m��-��:Xn�;g:Y{.]@o������Y	�g���wX0�2]u.��m�t�ƫ��͔�5c�d6��D{�)N2�������^�b��v�"eԇJ�V��̾��7�Zs!{x�M����Vi��{/)E��Yn/K�_��x�|�z������k=������S>�}i�_%��y�+
o�/����,o	��'zS~�y9N��i�z����O��|k+c�׻"���4[��f��"A�4ϐ�"���*�+e�S	�6=j�hy�s�pb�
��Z2�s�����b���~�Z��t���\-{��Q'��۬��]L�W'"�9;�و���L��=Z�f0�U{E���2m��z�a���,�=@���X}��һl+!�g���K: L�D.���ps�sO�����x.�$p��Dz�<'��0y�q�.�u0�Ŏ{W��^�okw2;C%,V��帝��V�bY`
�R���L�u���Ԃ�{k�zK���)���jm��:��qמ��>^���w��xr��!:&Q�;^Atn�d�27��tK33f���$͔jSr��fg��a��|D�A�Sl.��(��`�Y�/9mXոT��]��M҆�o���ۥyŇE�ןA�;Z3�(o�ъ�}�L���n�]���tG�{O��]�����^��2k.��v�t��l��z�+C�͖	A���@�3�mLǨA�!�S,J����Wl�+_4���!��{1&���=��Y�f�ʽO�Q�*���1Ϳ�:$j�p�{0TX�4d������������ד��s�!]��3���ġ����+�%2�6砯_�f:Nx3ՎX-Y�Y-���3X��=qV��y�:����4�d��� g1 �C�9��E���<S[�,��G�-̃ju�>ڧ`r8��K3U���爧���2uj(��c���}���@2�� ���{ ߵ��[{!�#GYЍ�	�ؚ2��5�d"?��y;h#^�ؕ�ow�uKw�c�4e>����]�j?pYJ��dP̅1��j�r0�nE�<�c�yg�`��o�-����v�b5��ʾ�#����Z_ղ\�r�hʚ=��Xr��r޳n��v��KRfٹ�0��F�`�JIf�7^s2��o����.���}����k	��'�p{�ȳ	и�K�����/ b"@r�x�bE��r��Y�̺<�,��4���>�L��6O�,؄$�3C�[&(=��x�7�6z��p��^�>> {���'�Kuu�y[�ĭ���J���'������y�7���ݐi�lu%{a'�C].�zKɹ�7�p��4�}G���B[[�`�D��F�ueK�G��	Eռ�4M�ˆ�X{�l����f�q[ݓ9q,45��:�6AP2:O���EluJ�=�vX�E���a+��U�\ww�����b�T��qV��2��H���!w���bڅ��*��h鼯ٽ<�Nm�bS�s���\�z�
q<�'��m�ʛ`Au0x� w��T^7[}k�I��F�2��tƲ��U.es�/0��	�\ӣ�a�8���'���>���SR^Y�n`D{��Q9����P�;ݰbZ��eP�L��B]֍�z��%���q+�mz3䔉��e����}]���Ri@���>���ϒ�I�`��G����H��׏�.�����#�z�g�,5Fi0���tǫ3ٻ�9�<ju��N�ݎ ��Z���BT�\ eS��Rmɲ:���]	r/*��!*t6�pM�jj��������:o��c�f�}�b�^b�	Ԗi��@����	��:-���]�w����ٕ���[}u�Ӕps�l���;�8<��/�����۟����:�_Nٳ�����>��9��@P]b�W?gN���]�<��$��<Nv<0$��z������f�t�C7gW�ɔ\�A�r;t�ʌS��շ�`֡P��'L�Y$k/����R-�ӥI��W �[���n���*r{����E�o_��ûw'6_�N{��h�^����C�y���.M�Gp$F�n�p?Mٚ�A�;ͫH(tV�V�7����à��������x>Z����u.�
���D��j
�.�w���盨�\���_H��,�`6��e����[P��!9�K�,�7b���{d^�L�X�m�97�c�Yƃ��kʤ�P1\�"�|��p�L?�X���w��%)��kXD��u����hz3�<B���P�P�����4r��D�]�SV)a�r�}�2�C��;~���/"y^3ܷ���>�d!<W8�.��{9�S����C�"|,Ѥ�^4�\��~~�2���G꼉��ڛ�+/*fR�W���IM�M�gg.z:Q�Qd�N���$uC�y컃�ڗ�����T�[/����D���kKM`�V>���pз,�NR��4�;{]v07��=2�S�����~7Kx��o�0m�!BY�2�'C����$��I�.[Rq��7�<;�+����,y\�B�
��@)�š��M��iN���{�D�&a����LJZ��T��Uf�X���w���k��`�O��";�k--o^ݺ��A7l�i�4b��:�VrI�����\-�%p)��/�+��)p�W.q�y�ԅ8�n	�����bo���!�f�O[ g�W��:���-��t��I��K>-����j]�l�7J]�6o�Ve%2��}�%�B����r��:͏/�Ft��ч�"�|��T֓���/�5����s��h��r0��bA��鈠͈�~��q����V�����7�b�l�^��*���;e���̂ub��(mG�u�U��>����n�����;�T�_5��
+�GﶭG?C��:�]e��.Sǣ�!r���V���wW"�t{�U�-�k+d��ﱬ�N�V�&Y1���e2�ۂ���<��<�puMOs\��=�v^����v;�Ʋ�;�z�z~�#E��z�ϼz�]�E9��c���f;�)`��2�!	��^w�h�u�'+����J����+%�}ɶ��fo=<��f��a2�t�]��E�gY&b0g��L���jɘ���_VEufn��Ozs�$��{�`�;����JP6}�=�k��^Qfi�ӓt<:��́ԁ1���6U�+%��w�s�2��Ƈ�TGR��b�7)��Y��ag�U��W_ 򜚍GLZ�/]-@3��I3Vv\滟�
���_-���z.�v^7�4��TB��)�N��*K2*C;�������*�dTE����t�Vԫǳ�,q5 �Q0��z�
��Ζb"S�xOBmU�ĺ���WQc�տx�@l]���(n��MWs�
ٓ1�jCv}C�2�@�y#A�D�z�ĵ�ə:�o�Ms�j*n�Z��&�]��8����y�d��*(�P����:4`��y���h_&��e)l�u
�L��C�{�dr�љ��釆��2��`1V �R�x��w^���G�H��GrU�8m��ڋ���]��=��ڡ.{�
c4c���2[�����������NU�<�F��W�u7�ĦQ%�y˵AB߳�k�x�s��|��>�7� ��G�Y��vh�X˥.����:�IK$�����pfg�ǘ��l]��쏲������7����=	�����|�R���J����
��Dlj;�y.�Kw�,\mh9�U��c�T<�|��ō�w�Q�H`�c�]����f����%=�Yʶ��+�����ჟG�fŔ��KA�>{a������x�7v�w�C\���7@��*'��]G�s������@�9Op�D�r����,��sv.y�/.U?v�~�����f�4�X���Y�c2YD�wnuֺ��tnȱ}�G����cWhl��62���C]��)\��(��(�U溝�㡋�L�D�'��ȹ��2���*
x=�CQ��V_[)��:6�����.
��FT���㜫�z�d��.�18g���>���]�T�©A�b0ß;��y���z]���7�ޓo�%�r��[<�l�\+}I��=t���K�������]������"�G���@g�x+��wl�O�#����*ÿ|�Fq��t�#
�-�T�R>A��.��w!#*���-<&��W{��-2G�)�`�������90z�"��Y2�Q+��f؛�e�0�
=psw�����K��-pVd�B�s��L���U�$nF�
T8T���|G�>��Ɩm��^�qҧ�r�
��0��'���̰�l��7��d��<����J^�g��%*Mm�d(���� e�Hto��m9�\��{S��{6nA��>dK+�z�}�7{��s���F4Y2p5�љn-��e9�)�u�hpK�ݳsn��kk��X0�J��M{^��g�:Ɏ�~Ml>K�3˽sj+u�$}U�:�d�:�磼���o���x�"T�YqsY�f?C�$�����m�]��D�K��"�X�H�	yظ+A��c�I��m�ݛ�I��ͺ=�ǳ��-m�{�$��/*v]�gDm�I	�A���Je*X.��������5e�.��<U麒&�~�ykHt�r�Wt,��G�My���svZM�m����~]��
���K�Suջ;OE�5���9�E��j�Xzw�\��v���
���6�KϹ7F]�w��<U+�ø��kl��i�A,�	��a���A:�pg`�����@:>ϻq���s�Ιs0i*���[R�l�j#�F!��*Pu�n�&��U�M��;X�E�Fvu�
���.A���+^��Kͣ2�vl�H|����ۧ��z���� �Ǝ#��!��������W5XNE���O��/vbR�;l���]Q
�zsc۹��o���MkrM���׺�Wl@F��0�p��f�i��V*�a���.�9GWu�(>�1��l�"�B�>;c�i�ŏ9�-�q�j
;ٵx.�7v��;�c���[h����§���ځ
G�d:��#XË/R�8�9���/[��ݽ;��sk�/�>b�ͭ�jj�m��Ѩ+
�f�6J6i�U|Z0W��i���#��w���!�٭��P�PbU�7�{�
�S�o�L� .�k�㕳$�A����OF��䖖�&=���Z3e0[2{S�v��P��d�Kn�iW�+�Cz�f�5�e���yh\5X��2T/4J@G�����OJ�bCp/{U�F�u�ju�3��˷aQ�Ĥ�l����K(OSma�uG��w]��>�[C����B5K&���br�*�z�Z2K������k#��j���Jŭͼ��N�ǣfL�Y��D�.e�b#[C���Ig[��C��:����&��:���+���ے���A��k��,Δ�����w��[Ow6Û�UՑaq��U�i�,���� ���d8��n�E��G{B��Wb����J%����C���6 y���\�c��$m>��NM��:�����q��!;��=���{g$���g)(�f�J;�"�Ztz��*X'
�6+/j�3��YN��F�#����i>�ɳ�y���
��q�
��nV��qn�-N�)U&�W��"8��
��3�u�6k��q�vZy��C�d�3�u���Ջ�}����b�:�L��Q̜kII6�r��e��*Ñm�el�Ԏ��gx�X��K��;A)�b�5Y��X��Ѱ�#=K��܉)��(z������j�U��_^s�/(!���+A��E̦V빊����Eh��fl/�=]����=xA;t>�4-��k�&��
P��M�}�L�]�u�Y��3�ѳoN\�bs;d�y#I�{bt	������B�P� j��Z*+R�*1Pb-h��[UaZ[ik+�J���V�V�AAkm+QZʫFV�jX��DUD�Զ�KJ6��E�-��6�#J�m���-�U���j5+YYD��-)h�l�E��X�F�ZЭ�[Z�YJ2Ҵ�b��m+-���(��am�kK"�X2҅�E�����R��)F��ִ�l�i[j5��-��ڠ�iR�Ԫ�JR�+m+ZVKZ��T����m�)Q���Z���TR��%���KUm-��ڭ�U)[-*�[Z�m"ĵ,����kmIFѩZѱ���h�ѨV�lmmҋ��[RƍV�j4�UQlR�j�kZ�U�X�UADeTR��ڃm�J�F�Uj	D�Z��FU�,��m(�"���֖ڔ��F�jV�KK(�mD���ؕ�������ִ����T,DI�
oM�.�l�0D�W׏���\w��Hw���rE�"VPAn�#Ak�:\��r���OpQu�8:ŗ*��)whIPɺ0/�	�(H@���O!��n��c$���^\3q��f{7|�h��C�:��z�]4����R2�ް��Ѐ�z� :����e-�����b�u���eLu�`�n+]�<7����S������A�s�@����&���{��)h���j�1o�=M7�l����6�'F9�m֑w�#�Y�<;Ӓ-������v�3����wyJ�y���މH{�>��G�h%�j���f�q>�ڦ!a�r��Ψ]�g�d) ���C�C̷�n��I�A��kcEh���������hW�/x����j���L̔��xu�6kǔ�����/����ߋ>���nK���<"��.d�u��V��]6�5��:��`�&r�*ߢʔ̛���,t�YF���1�%�k��u~�k��
.w��^쵯�C��(Q7O����E�L��*/�qh���!\�!<=(#��/y����=ؒm
�&e��yJ�2s��X��Qa^D�Z�œ�A<���~�pg�����A�|�疝�]V��뻒�l۲��}��C�t���"O�*3f�#PH�{n�@ru�OG��c��Y\����5�n�[,��U���m���-�6Z��o� �}�G��a����a�Y�Z��-�ؕ1�1�s^orz���.�B�F�aOU��7�g�5�)�Uɷi���ut`���r�)�S��V�W�ABa$���@�쭉C�狭̸�6��'���Z�=�'��e�[�Ӽd�<5aٖw�J����	t����v�<�	�>�S�^tƄ�۱�g�[GL�e����'C���D�C:�*.w�~K��u�����I&٬/���vD�3�� u9^|F ��{ v�������mI}GAٻ�L�&��y騻Vl=Tߐ�ʤ�Q7����ˡ9^|N|���Fǃ%��R�U���}�,��j2�W��㛞b�vf���4җ\NW9WF���Bi>7��ތ���ۢ�^g.��k��0`��{���㕸�$]�S����X��@��$\�ͳ
���Zɼ�}���&E�e�Ύ}�6��P|�#�ue�*��B���!*HE����=]���}�c�c<�`�ߚ��"��[�=Mf�Z���%2c -�Y�H\���E����3m����Ռ-��]�|�]fm^�Q�|����b���f�K�������LgF>�u�5�w�v�ڑܬ�_'4b�벋�J9nҘ�l��w�����5YX�Y�����^3|�3�.V�JH���_-R�qr�[#�ն��g%�񦛗)���Xt'�"�>�1���Gt��lv�VS�q�<�L\O�!K5�rH=�̢�i����%�Vg�P���K���j�<e��g��y;Яmr�Bh�O�1P�ͿxL^�$N�<��(�4�y�M�>���At�F��k���6�2�BJ׹�}����A��ш���<'��K���B��\܀�WҢ��5����V�+D}9�}����
��TaV�����"S���F?�6%�n����"�CeA������I�ז�%7�4c�&s@�_��9�##Ib/�WGPAt9sĳ��z�N�Ne
�Y|�:�z���o/K����6l�C6��ß�O�W!Й2�:f2�R˝y�|�O%�R����0c�e��z��33��e�
/�ʩ�eM��`
��S�ܾ
�-�+])���,�U��tѵ�\��z��S�@��T��3�ls
c �Pu�}K7z)�2���k緢�z��95�z1�Xz0E�*���0�P�t	3�i�\�xAer��Q�z�8�Kgk�|\���F7c�V���'8�M"�T	F�Y���5��������s�<Q�����߲��%7K�w�ب䡭��Eí�;�fn��r��च���ި��ͧ�:ל�����QP�"�O�{���9P�u�C"ǻ6
�Q��G���^�,{��:���`�b�])p_ۻ١�C���IK$��:W��}�����6�++�z��i�s�a~ʙq@u�e׆���$�t�=��4�0$�O�:6�z_����T�rw��`R�� ޻�
r���kU���:T;�������{�F���t����y��=����jy��uc��~8E�O����=�h=|�����������^���m��nH�sr�̦o.��|�]�WC)�}lL�w0�����~��Ѡ��}�G�!;��3G�Ĵ���J&�F��R�v#�_8W�̃h�o�u��Frؑ�S�x��~㭦�z�*
���c՜3n��n�%��T��]ax�H����{�U���=��<�e��[����3J��*��}�k���_�͉F�$
��7o���u-�Jaװ�$t�qk�ORg}Q$r`�+>���t ^>Ufؕ��9�xb�dY�sU�4׬��\��pV�VG�����y��F��#>� !���b�8�������⦕l0�r�W��`7�j�:��A]���[u>[��@�C��lӋݿ%3)�\�Ga��].�[7>홯7�s�P[�\�&s/љb-��P���]���tJ�[q#R��M���v�@�+{U˷��:�6��kƯ����ۘY�U���}[��s��u�ϧ���q=�6\ӛU6�̛`A�7�����͇f&�����x	Nx�<)��^��v�tƲ��R�W;�sXGX��ٯsN�S��b�b����rrr�|����-`�	�������uB��v��=�j�9�QA�W�L�Rwy��S>���޸�2�H�,�'���I$�E�����1l��!��]�m��������\���R$��8 ��.yYA��]Kn�Z$��G�]R�ᛍ�6��{k�_ky���T<���o����� \�( }�FU{�5;|��ӯ^k��nE�yc�(�]��묇د�����ܠE��<#(M/�ϔ�+�{u��q�������8�x�~�2q�l_U�2$]�P�N-����f��`�Ƚ���\	G���۲�$����(�FC�Fċ�p��W�q��4�}׵LE�-���5�\���B �E�b*���s��G�I��k l��A:<+���R���zͨ�W`��l���fC~�5P�����;z�� �Y9O���r�"F�j�{>�tӼ+m����h+1�Jo'��A�-�R�j#�Bړ4�K���ى����C����C�;�d#��Z�-)�0D�7L���B_��"#����|�@�2/DгY6�T�кS)n\������~��;M�s��R�=4���/��f�elq���e����Dd�L�9v߽3]�I;)x�v��ǣ'*u���b97�cB�4�8�U'H���)ٝ1d�9���*s���_�����r���{���N�ȏ%��-*���L�
{�!2.��k�k1�n�:ri��$Tf���,�o8;K�� uY��ʙ�[�py�_^�U�Owgj�os�!�Nǀ�L#h)��N��|Y:���(�WYͳ@������]�[��*�eL8�y��DByL��C�H��VĎ�r�ίfx(l��;��]��\C�� ��;���Zlu�DLS���v��!lDB](�#�����@K\��{w;mn�'�vo^yp=��0K=Q^t�	�A��HC:�+�Ú��S��oW��g8���k;Ƽ:��6Ҟ"30����U9^|F|`��{ v��M��^����r�>N�q�x�yWj��j͇��!Y�L�_\� �����'Z��c+��VeZZ�ͭ�Z�����R���72�jbky48:uW;8�������(1�`��.9y���쳰`����������(�Xʡmf�K~0u��v�7)%ɖt�X��
�����Ε�7$Rdi9F=���K�9��{&��q.Wٛ��Q��gRrQN,@0�1�:�P����K�Eݺ�pw-�7ZN�^�L��u�5:��&�_LD1�ՁG��cǮg(/�W�t�����p�V�Qb-��STr�53��#sz�^S��#�Nð�0`��:��:�A��]e����@�'N���N9n�Ě����YN]�ܪ}q�Ym��9Mf�Z���%3��3��,�lZ��<��f�]�q'�eh>B�9}lL��fڎ����5��"��l����6NZ�S���#|�kI��S�+�2�0���/Ӌ?V	�NW�mU���|�)O}�/�^�'���!du�N�E�!0�ή�Oa0ªv��F��i����7<��-�=�!�ԙ�@lȡ�C<�éJ���A�"�xo�Qd����).����T��b:5^{:��1�:]DJ`�&�߮6%��a��J����ۓ�ގ�G�4�w�A��<�#�eP�ٸ@��vhz��e+�3E�
�ud�yy�qM���73���n���]|G��83�MV^W�H��j����c������������^��O��͇C�	�j@�G�źi��9�T�sas��E\2[w�5y�M�Iof��sk��ηA�.ʷ�����s�n�׮s�[�.ps���߽}�S�k#�*���U�W�s�D�c�� ��L�	� ����<j4�s�W�\'�N�Y����1.�$��d˃�m�Ŀ����%o{�ǖ�1��i��������#ː����ds(���L�.����k��#��}uT�O�E�	����\,�S�D�k�W�j����?3���K���b}2�\3��U6�H�}mv-�#������e�	�;��+�X�Rອ������'"<�vP:q��{q�egɪ�NGR��Y���C����.�#��\��4!��T��Y��[Y[�t�-��zZ�������#J%��`�� U�S���f�od:�\�:ͣxj��툞�|�2n%c�K�=P�9,/ǵ+�+m^���cF|�<#+g]w���b՞6xnL�G������i�<��5Kda�R6�g�V���S���]����ܸEg�FD,M%ulf��Λv0z����&:��e������R�]aT���F���&y�x�a`*�+��9E[b�m�T���j&�VhL���7v��G,d�M�n���s�*߱�����t+/�5�(����$t覥n�r1wPNQ�)�	��%G��ۺɺ��֩�0�=���'��u�H�>~�f����O&�]������S.��Ux3���]%��i.�����D��Ϫxl�����~�B䗟�g�P�=K(O9���:�o��ҡ�����Bj+��~lK�]�-��g���ܘ����i��"]c�X���L���X5����D�OC5Z1����B��x󹥋�+�2U�Y�˜v{�
ؼB�����y��=N�����4)����|�fiw������* ;(Ѯ閬��N��0��箐�q=�6\ӛ6���K���zske�.z���%5� �
a�5�p�jLk+Lr�W=�/��=u�~��7�L̎���N���֗��뢢�:�q>uƲx�K�j3�l�֬3�*�	�c~���Z��8�eNq�"�ܢM��9M{��p�k�ю�Y� K�!E�����7$�i'a��ęL�τ�t1�YBx�1�Sm`��a�yE��!>��w}���`�6��Fx<9�%,�԰=�?Td(��t��S)m�4����-�&T���_-���|L(�ՈK�<�U�����ё.dy��B���@��f�nS������Ș&�D]�w�C���c��c��7�&�]j�V����B�)�
<������J����5))e��[��e����)P*^\��od��"nQ|sز��vo�ev��C�}��5��ܠE��<#����,
{|_��^�f�4��w��6�I�m�Nq�`ɟu�5n�e1��X]m��Á�:-��O�3�>�u��%���_�l �@�����[��fX�g 1�d�g�rҢu�cqO7j�G<x�d1�M������ւ�8+Å�t�Y0�;q������ b��`X�/(��*jSt@��pC�H��^ds=�k��(��6�b��R��v�n+~����2I6���{��G{r�b�!s&�p��\j�ű�l{�ϡ�_��5Q��`�}%F���=�z5���3�c�]�]e�o����2z�@���\u���T��-涉��N��Ǜڞ��
�H��ܻ���2pv�'lXDY��ʩ�����8-���7�?*�Y]R��=�0�� )�W�;W1�d�3���.��] ��m�7��'�~}w�̘�i�ε�`��h����q��]�?|�����>��H@��	!I��B���IO�B����$����$��B����$��H@�����$��$�	'��$ I<BH@�XB�D	!I��IO�H@�xB��@�$����$�`IO�IO�1AY&SYp�/B _r߀rYc��=�ݐ?���at��ހ�`m�B���(J@a4��� 	��)@($ 9b hi��]�򧪣A3Uj�����m�[V�6Yl�l��}d��Rʶƪ�q��P�Ӷ�ywF�Y$�V�mT��m[YKe[2Y[!mm��Z�FR��j�kl��d���f�k�ɮ�獵mV�� �	���n�]84;�}�5��j�ٝ��u�W�^�)�n�[�,�Щ������V�X�|�����}�޸�׽�W���%m�z���[k7�nݮ�Sq��j�o;�:�\���ݺ��;�z^�)����sp�1Bem�YY�  m�W@P�{�(
 �w^�   z��  袀�{�  {�{����/oN]n�;үT����9�v���۞reUv����c,�ڵ| ����Znc���=ٖv���k:ҧMJ�\�{���vT�������͢UeE����3J��G���m��l͵-=� ���mY����Թ֧����]�;Wv��8;�����Z�]z�#Z��z����[��6ꣶI$�ݸ�Z�� �\�� �m6�U�]ۡ����u:`���h3;K�h-dvղ�4%�� w����6�]0Dݭ�t�R��9Jۡ˲�S���m�B�Q��Jѳ^  ]�]��n���:s��\��֮e(5�@6Xh�6u�����U^ښ���_ ��ـ햌 �t33��7p݇X��T��룖� L*��&��@��6շ�����5Ӹ�\λT���n�0n�t� ��΀,���'�     j`1R��2h� `� �� �{F��JI�40� h�M�)�1�U       )�M	RT�  �L��  i�0UT���(�L@ 4ɀ �I�Q�a1)��2d�&��2O���/�>?�����^�����1t�F#�G��.7�Y��! $���~� H���K!4I	>��H	�A����F�����G�#C��Vt�*I�  ���d�! $�K2�Bv� ��O���Î&��??�����  �:��_���!��Z��}��  @�_����E��S�BZ�i_�! �aٷZr��X�ꢊ'!s)U���n���z����sn���H�J"��-՚���D��QGaZ�a���V�F@P��#�7tJ�%!��!���zͪ��V�De�%��u�·������$�L(���kw� ��ח��Ӭ�K�J�c��aStv�O��Ҋn�lOq* ^��B��n�
�e�-�1�a�yV�#\JRvV�[z�+�Eb	�zB)��T@YǀU١�oS����E����jK+)��ҳLRR�Nݏ�ل�4JʈkјB�ݵ�fdu��M!�r�Z��j���TXW��ǳT�/��n9̽ $3~�1���1Ѣq�qe�A�.e�փuy�h:Jȣ�+A���h�kT;�4)��[ɦ�0��Z+n;!�<ɢ���젇ݰX�өMvVrnd��Ӿ|CA���P��QnGz�{W�@JB���Z�ѯ6���Xow[��k�`���9E�1%Xں�5k�X�^��Z�KսDH���R�j��>o+�M�k��/�Mr��O����eotu�`�9N�u5E�$4�:���]�����K��Y�{��X���<�-�U�3���5*�u�U!����#@V���U}y��[�(U�S��˻�PQ�G5e��S�b��r��ͭf�L�]����V.���ݘ&��>Y�˥[J1�o/U��y�[4�x��/��
����#;#v醵�VÃk0�TI��qe���X�J9�����,֋I�SJ�����I8j��Ll��F��3�^;[�.�y�E%�b�`%J�:vRۙG9��mcW|jQ&��cj��&���v�V�o�|/�hܴrK�髒�	kfv�i^��)q���*���N�@+��X^b��ޓ�k"��6	�ݵ�
{@��Ŗ-�آ�h���(WV�M���ˤ�K�����b�6�*hi���V�E��Enn�D���1i�.0e�j�4��Ae���J�Y'_V��l�;��t.�{��YKX�E�f��	K;� wi6�0i��D̑���D�f֚wR�VLs>Z�����*�F�j�+y$��˕a��V�v�}�Q·l�;op��]�L�/#��R[&nh�P��L��B+v��8B���˫Vk4��<1��si���qռ�i!b��W*���bzͽ�/
�H��;6YMfZd�ۼ>�
�',�v���HJ��zu2g��W}��Ŝ�f]7�D+cV��.�֭Y�6��(�sk7$f��n�
�*ag2�\>?en�m|��-YG^��F��R�ǮSw�>�1�kC5{M��������Yu�%��փ*�ˢ(֍y��v��,!JVi7B`�>3@;�$JX��ax�n��0Qw���f��^��v�V�N�7uv$�DL�ѐ����aLh;��nm�VZ�5��vN�)�S��+��R�
��]]�r���|��q�c��T+�5���s)���v�i�7O/n�#t�Mjz���7�M�)c]��uWa`�����x�`b:1P�c0<WD���V��%ZXM�ͥ��r-��6���&�[pP�z/X�N�*b�M��2��]a]E�괳�լ�U��mG�{��Jօ�D۫��d ��[�tJ�E�q�;���Y�.�}r��d4���H�l�r�Xf����)Q4��]]nV��v��K@�ze尨V�83t^��ȋMɌ+3��n�����g�0��'�m�T����ʣ�ih�jѿ�9b� ��P���K{b����W�N���XE�5ͺݼ��KI:-P���\�1R.�ښ8��n7l�T]i�D�5ؗ���r����mP���C.5�`1le t\�͈�k���F��Uh`����4�Dh`��N�)�P�"�n���`��M���Q	B��3�wI�{D��@c��$WJ���/A˼Ie�gm!��������v`|M�A�$�ZMLra�b݇6H`���Gۿn�oʖ+m�o*�X�)C{�.��(4Co]��nQP"jj��텓5iy-�n�B$�l�Fd�Ԫ�n��Uvz���l]֝'IUl/r����$�ѳV��+YL��e]�}8�f-H�Qfл��j��-�h5�I��V�=�p�h#�]�ռZ�gDh�U�Sj�2��ڊ����yhl\�ͬ����c��ʈ7��8����5���D�h���ŀTz6���JJ.XԄvq��O��vq�J�cvj��r�f��(Vo赬�j���r<z~n�"40ފ��5n�f�8�C���Hw&+ڊ�R��mnUm����(���]�R�ۧx�J"x�#q]��W�;��bN�b˕�fi�P�gp��'��lU�"���[�m)�kU)g�n�˧y&�iѵ,A��bI�f�Ӻ,�ӻ�1I��Rv�z���,��*kV���ݣ�R%�X����CI!S�zu����(�5t�vһ{E6,����]]��T����x��Nd(,ĚI��j�RpT��N�Yn���&/��ED���a�U��� ��N��>FC[ET�PBԄ�m��6���[R��L�����5�ڄ��Z���,Ư'bJ�c	_����6.Jeja��ͰUK8B��9��1u�)toE�o��V���W��!;�7lm`��f8n����r�ٌ;܉dԫA��Y��+�WW����S��Fκon�fTvU��۷��^Չah"U�I���Z��a���l�|����� �۰*��{�����Ҙ�&��ʗN��Z��,8�d�]�o$�8�Ӌ^7{�lP6�9��!���P5�l�j��t�Q.��2����j�q�L@�2��j�ڙ��=t�K1���FEr����gA�M�� T�H�Ph$꣣%K"2l��5sEn(h�50����;Y�sXU��c%����P�
{7]Ը0�V`������U�m�
Q,ޯ�i�E:!]�f�]�8/T�4-x4�*��:K�zĵF�ډ�;7+0������}E�}��m��v���7KlDj佻�+�c�ѵ�$�0�y��j�����`�*b��[����cUՐ4��6⿖<M�Ȭ��Y"�)37AK��ܶn��02^���[�^R�U�iCvc5nL��-V)<��h6v�m$�^ �"�2�^ƭf,KYJݷ�(K�s9Ipe�;C�+VHn��j�^�Q�J��k����<ܩZ��J��X��͸NY(��f��CV^�2���[�Wq��;oWl&�[t��yb;W_҅�P��u��N6 ��9L�jLQ4�C���Ǜ2[��3��nР�h�SN]'u����u�܈�:�MT����]��O�2���LPJn�a��1����u�k�� �`ҡwr^[��W:1� �F�,�j��ZU�k;wD��h]u6�V(Jǖ�[�ie"7i����^<X��%*��7ՙ{�6�y[�k9q���f�:��j�h�j�&�����*r
�Cf�,!ɔZN�;x�v2�rz��.N��/9&)՞�[�%���|tm�e��t��h�,�Kob�,,���ӦE�T9�l�a�c�(��*�x�
��@�*Á����%��w����`J�Tt�
�; �d���̭�V�T2%��fF�M�Ѹ���j0Q���NKIՒ�BI��/��pV����f�cwJ���R���ۺǁ]+e�5�]�P򵒬�u�1K�%�,ZeeK�I|wR��$�^�TơT>�S5e1� �O,mj��(oה�X�3��3��W/1����T;���u-|@ϭ����I�|Q���q�Yb�e�2�u�I-Jj�����2L��V(��Bm1����mӊ�Th�,�H�]C�� h��iI��5��Zv�W�����t�ǹ�-Z$��1�/�'�����d�=��L�j�)Ee2��n�"�l�҉իʆ^�%�r�RN\�`��+�M�:Y���=V;��]G�1�.����N�%���)��S���uK��.����R��v�c�[m��)�nh�N�D&���2��mdV�Ye��ؗj�j:��ɖ�{�oi��I6��i>�\5��X�]����-f�����mrEhi4Uga7��˳Ǵ�0�Q�#j�卒���X��3~�����7x�C�.� ��wh
`4e���˔�ɂ*�TL�5t�˵Z��	1��c����7Xq��&�#NMz��uyh@�0��NC{�=R���&���6�!�b�q>���1�9���oו9'�z���>��/���pu��?��.)�� �b�9x�A��i�H��� -�������Ճ/�_^#�>�3���ʘ���ȟ[���Ǿ�7+s>&�:�!�m\�c�)�ftSy����#dn�ֽ.�Bk�O�����W�ҝg�aas�f'�X�,����ɹA�����7�A\��ׯ�^jQ��J:����M��c�f�,�ü��CIF�/�de��v�Ɣ�4��9"�q����ub
�P
`�މ��4�F�sՠ������1P��Y�h�,���4�1u�'SU}�/��M�:V3�K6�wQmkte�٭n�b��U>����.�(�n�|�aA��)�
��I��k��䮊FE�U����q�*Ȁ��͆�.m��6�6�:m]�uŽ�͟py�& N�� h-ap�]�	��J²���,�u.6�r��|���[�!��R�b�� ��\�,;"ʫꗆe���g�i�z6�A"�SX/�j�̍��.4��踝��L�"�\,VN�{�̶!$��c$�
s^^�jIB�f�ȳ4<X��n���t�of����S3)�@newC{B|mM�L@��׏.��+0#���L��%]`
Q�Ǩ%sH�ORWQ�sa�5WYc(�C~螑2�,�T4�E�N%A��(��%9�� ��	�1�8Ý-��$ːP|��Q�&�]��[g��i���1�D]�Ȼc��_����KO�穼̋�f>T/�����.�B����oL)��Ѧ��񓚻���+虱V��үv���*��\�$��|K��椈��k��4g4r
�ut�u��ou��C�M:�1r�p'd��^��A��Iܥ�%ZJ�j��Gg9��E���[ktpĝ�<ۿ��[|.���tDh"E�@<��.�b�8��+u>] �/�>7���`��U�r�r���e���@���Q��|7G|V��9�uG��s��^h5-rׂ�_5��c�������.a�'Z�5W���5�O���)��6���P�L�EV]>�1	���ܓy�*���!A+���g�B�-�Px Շ��+5�)s���l���/#+S��*����7D�y-�%q�58l������)�����7�q�*�qͭ1Y����q��̙���W�:�{d��k$��*@�����P�oM�a�1[�0������m�۬�EQ��e�1ɫ<U�kNo|��IX�h`��٭�?�U�f�co/S[�e-/kROav w��2K�1Ȱi}�A�b,����F��ε�bɕ��L��5E]M!n��/8��#���\?.������n��/�o)��c4*��u�k�D�aSƣpe`b�b�_V��u��+�C��a�twwo��-���5+v�t�RBuv@��܃�J�^nx�ٵZ	���RC�q:覃]a5R^��7�v�H8�4vCC�`�;L��6yhQ�]��C�^R
�f:��n'Iv*�;)��	u�i��}�[�N"c�KF��Z�A�{y���X�[�"��e���5��oh�S��Q_uI[4�u���Luh���,ö��� B��\��8���uY����_�6�.
PLvU���QgS�����F(r�lu���v�zɕ���J�����y&ݼ�"ޓ��K`W�V8��<��I�S�B�ܰz'�J��|q5�h0�$�;�P�D]m�&vP+B��]�U����j.��Q�Mk&��G�`�4I�(�M��8K�Cn�Ȕ��ck�v�sǘ��aVP�R� jgs��=o�.+�"��JO�������H���kn8w)�ѡ0
�~�C���;Jh[�z�] ��y���5����!���f�
q��X^�}���B��e\j��̫�zB��h=	�{a��ZL2�[�5�.L����ִ�k�̻���O�gAA>�>6��8)5��$�M=�4���m��}��<���Cx���Jb��롚�ncÃJ��t&4��&��of�Q������j��,�Σ���Tl��y�yfi�8m޻�,�hG�p�9��Bj�e�ĆY�t5�ԋt��/i�1:کB�3&h���r�H�a�n���7BE�s���nGb����ɣE8�*TKf�m�.�r�)Td����C�v�PiZ4n�VHF����;cF<�W���;h���`"��c�j%V����R�*#_aL���\�}��i��1�)�2&s7&
���	{ɶ��ՃKZ>����ٍS�su_Fk� ��oD���a͉s$��b\�u�լY�.�uJ�T��}Ț�v�YWSp�ʈ伻�oi�	�}���k] N�� �o0�d������#unp-��rʀ�Q.ޅ�%�K���42��:�8Qz���6m�LV��oB���̏5/�Tb��{�|CWf/\�N�-�N�R�"gZ���i�ts�h�qB-�HH�Z�2��Z�,�k^���L������4��� n��)n���t|s.�,�-����* �x1�o&T��1�N���z0Xe^��c��3�h=�mk-�NJ�e�F^�=�B�Jz��C��Ld��Y�Ծ�ڗ$*�uy�k��f_7d�O�(�Y}�{Cw#���W��;�F[���b�c��|��ٱ����4:�P�4���K-�2�a�+���:�m����Y�H��g-D�
�E4&b�P�`?��ޘ�&j��}4�K��L+���T�\�Ʒ(��ftˁ=�
u���� nr%�|.8�bLͬ�븾�O�D��z��J�#4e�S�.��:���/�-T�Kd
"򌂥[�S����M�NÎ��|u�BT-��^:��F�OfZ��8S�쬵ѲYG�S�P�CE��jX�̹E��	z�-w$�Jsm��CR*��u�Wsy��V��-j�b���3�u�/�n	�*T�L�Ä7ƚ�׳/zV�"�z�]�x�v�KEr��g���Oq��V_uӬ<m����&��#�����:��/n�؛��NrWmp��(Q����>J�¯}yr��_=��&2͖ �]�t´Ʋ�!x3�+K�C(Q��-���<�W`�oLn!�Ctwl�j��Y�q�(�൛���ʝ �ڢ�F�t)��1Ɋ�\���ۥ�	�Y@}|F�H���D��F��ZR��3o�ɦ�5ǉ��gO���D��t>'�����Ec�=P����� K;�Ⱥ)��IXו�K|�$�9���!#{%SJ;����c+	��V,4�:�!x�&-�3h��R�{�΄y��/v�;DU��U�L�ɜ7�F�sf�޵i�2^i��Q�K@j�:�`h�!�c9����Wz[��t�M�	�Wq��2�ƺ�]N9��K@Ա�V��8�022P(�mK�.��dĮ�B_<ujX���B��Vs��[n�ݥn�WN+�M^2��V1������M��7�`��N$�oo�i�x3��h�ne<�ە�pF
wSﱖ��}"Fu���W�,��!���V�����q�U�JP��h���TF�Dsɀ�M<���Ǡ4��
��������В�;}G6�	���.��\#���*k��Z���n+v�%�EZ�y�K�ڨ��Ձ��l��+	)u������c|�V�1��z�tM�����mQ�E�nU��j��yt�r-#�9���v۷72i�;�����V);�����X�e��(V�����uW�-3tIĢk5^z�}��wǨ��[ԏ%�0٥#�3�^PCb<�B���`˭���Q��ll#j�e'��[>�m7��L��5�ʉ'�u��KM=�;���UAb����=��/���2���❩V;�S��\�h.�ƻ/6ʹ*�
[�S�#Η��^�Fs:.T�`ж� �Y{:I�����������J9]�D�����hd�eS�Y2�{�8���ιX_ͧ�%���^��r&��Wԫ�5&�S�˜��\�_'�w+�*��9rM�d���$�:H��\��pq�\�QE�.&$%��Z��ӥ(�ͥJ�i�
�3Μ�0��)��0b�
�F�rG8��JK��V��IY2�Ⱜ���{�r����ZIN��Y��%g�$Z�����YȘ�3��a�Ԩ�P��P$�;�cK��fM�7���\�P�CM��F���Ը㩝QT�P#���"��,��%i�r��9���v��؂�:"1�-�L�yAg��|(Wq�i��쩒�Z�gi�!/"�n�u�J�`�i[��9p��ADѷKz]=�ڴ;`U2������룷���㏎�I ��g\B� o�p$�'g�H �Ώ����=�ɻ������¶�\p�|Z5)��S}7����j뭤�6�Z2�xG��Ԫ# ���i�4K�s�m=<G{B+�}��a���t�y��nRB�H+��񗏝�b��4>�gw��$�V��&�m�vh�ǫ6P�޽��t�ʪ�{X�� ��5<���m�Y�ʹ�7*�S#*��=�%�<oqY�o��,��S���j[o(4s��3m��J��W�.G{��n�1�>OW=f���\�t3sn���4B󶳤�Z����NQp�m(��������D����`�u�i/�>DBR��W}��ɘ�������4S���j��.�,����د6\�OG
��"Ɏ)4���V��p�)����1��޾ɻ��RTGvЮ��3'uFFw>p�̲.����,��>�ڵ�"a�;�v54uO�3�Z+)�nq8l�~����z�h8��V��v;y�4R���JJ�w�A$�\o(<���a]��*s8�ɥ�!�u��Nw2��w� ��͋TBz�U[SU=�OX��F'R�]�@�z^`�ٔ�|���:9��7,d�dZ5`T�	0Ă�4_ouw@V�f�)u�.����^0
��*ԱMz��.�x���g���;8[�����ݾ�Sj�6[T�j�S���2���A�\�(�q���m���D���9�gj��7g�q�!�&��*�t׶4�yZ�Sx�ȴ��\˘��7%m��xWBưP�0���n��5�cǣ��%��'!˪�z��,��P]5LX�8��ʌ�#)�a�c*�hn���ۿJd��Mut��8`7k�ʙv�f��Һeb`n��n��^�)��[[��2�]�k
�dw�+�4X@}�c�/���הV7���"��4���E���ob�@�{�oR5 �6��`�x��pQ���Z��MB4�Umdc�Y�'>�J�P�9ܙ��5�]�ܽ�.��f�2T��aɖ�`�[�n��r>R��4�IR�lf��p�]�f��B�98v_ MK#fu!�B(��nY�x;�ϰ����h�Ǎl�(1�x��g��U��;�jݝ�jK��iR��ҵ��2��!T�mu�)�i��4g<��NCC�ׇj��o11�}�SF;B��:�}��ŗu|�/e.�s�2e,��[�e��xc_*�oC�ŐN �+����|����i068t�y *���פ���wgF�q��o��[��'#�8�e�N�����M�z������EG�͌wtp�m�S���q�s�cT���C�%xT�V�5�n��u�`�Ó �򺘮56�J�C[3���`Y*�OѦˡ��4�e�k M֖�'�A�Wa`��9|fjC�j�Gp�(P�7�:]�M�����ϑ}�-nh��N��Ŧ\6^|��I;��k�N!�7j�N���h��qyV��U���C��'��r��ٯ�^�d�h���pD�_C�/���Pd땋�_N���׎�)n�]F�e���Q	:wab*n��0=�����Ī�M�b�Pm��&�������mR�ݭ�2��T���qf��<tޤ��Y��䁈�
W}V ��,���]��������B��`�vܝb�&���oT\��i�Y>�.z��s\��*�Z�y��ݱ�MhjU��� T��͎��4_-%\��������<S�S��J��m�ڙ�Ɩ���u)LC� ����J���6�]u<�s-�Яn�V��՚�-�(�]�qi$R�R��%=��a+���gvNE� �;�2�)La�W	�e-�E x�w]�,n�D������Vhٍ��%�%��Y�\�j�J���q������y�AHojpX����
���n��v���m.e�v�z��Kj����9Vl�Y|��f�C��K6��p�R1�b�N��Jggk���g��A#P�n�vj�Q�Y�5n���وr��6r�3������0�0f��''D�:��:�Ec�Ը��Bt���Er��=�{�A
�ev�=:õ�V���
I����3�����5�1�����{���K*2t�]�Y��^���oņC��6,WԷ�dAQ����\zHo���x jg:�V�;�M�a���x��W+�WL�娷���2.[��d�5H�圇2>G����%莨a��y1tR�ð��W�{��{&����u�L^��-Uq�owd�v�Kb���;��eF��iE�$���F�k�N�4;rRe��!��2���>7{��Zޡ0��u{����Ж��T��)�]n]�)2m���U���F�Q��TK+���M��(H���������F����)ྸ�%"x�1��n醙{�������ҹ���L�lܔt��a)�e*����j��CJ�k�w�<X��]]��p���2Ai�V�i�i픅�PN��]{sk[Bȅ�VFfd�x�eq|��2J7�s���L7Uõ��%��O�/�<{5Z�ϓGa������c�w7]�����V���Y#i�n�F02���^ҡlŴd|���KH��ÿ[�L��N�U�V�c��-���ss��l�WOj�(�V������7�l$�e;�rT� P#|��uPi�7��AV�9��"�Ը��S(���t����M�WH&z�X��
��0�B�lM�&bߺ��(浲��͊���-��vέm2�"{}�n��÷yrs�#
Pe�G�ݔh�,5D/)M�JP���&������>$+��eu�M�Crf��!Шns<���-�|��D^Ó V����83��T\,R
�Qb�H�}��f�P{w$��i�ަ�<�ރ��������έ����8���v��{�UE�9J����,�%:[��ݲ�,�-+a���ʟ��/D�bF�N��kHP�Ό�3�C���/����`�6�����o*p�s�i12�'j�P��K1��ףuvX�P��k/7��7hȖ� }�N�[���;ox���}�M�w*��k
�\j�����Hm���ұ��D^#}I[8e����K!c�)�Ŝ��/�����h>�k	�+��޾:vڣnm�f�j����VE��{��Dni38;p��j��Ѓe�S�=i��3o2��`�Y�T��Z�Xա��x�^�I	��ʖ��6���8�3D]u�m��'n�@4�WKZ���e��,���f&�F�����W�(���a�w�mpo���MNQI��t¸Me�+E�,�j�-�t⿱���.
)�@������u�ցׁs��R�K���w�.�y����ie�G&�H��o�W��%\����l��͢z�v�p^�],�r��S4`�i���C6jH<ة%ق��<��e1 ��eˬ�;E�B,��}/��Ҽ����L�D!����T�rv+Q��w�k8��gw`��Z�KSJ�i��V�䎩;N��f<�Sf�����t;�5�8�6`�==W��kb�h�(�{��:6�:.�G>$�I���ҝ;mmm�w�=54M�*��s�vd���8E�^d"�ש	O.�F�6�T_)�h���ͧ�6/��WG�dn�lf����u5�/�G\���h&�V,��`̣ ��p')��ԁ��vK���(�&�=�Kj��஘�Z�m6�1�o�@�r�5y�b�6��qN����	�� �t]h�O��}����Z�9;q��di\��Ʒ\�� ͂�[߸]�|ѷ������.���jEu�,)��]5e�C�
=I��c5$7M*��������Fv�Xm l.�p���FR�O�\�
\�R-�Ġ��tgY�����"��󩼦����ds7p<����Z��t���m%��'Lgmq8��@t�������Mc}�>�+��Z�ŌQي�T��t���nҍ�PìT{k�-ΛG3�
2h�i�~�)��W'�z����ښ$ܰ�� �C*��¤G ��li<�)�K� � ?�hǻ��A� �Z���ϲ���ˣ���0h���X� �w���z�9�˳��%�e��,t��vsX RzQ�:`K-������n�D'6I���K���f��-a����%�R�7J	#�f�=�j�}q.��+�T��f�Rf�̨��m�8�Vqt����6��LT�`��
p�:v���d�����2J|�*-���/��Za7���r����-�E(���o닊U�^��.E����lv�L����LKeh� �{x��t��kSI�-��Geb�mk��z:�'M��<����@ $���~�{�eP������?�"�g)M�D���kD���cWf#r2�.��
fJf���%r��w���:��\I��[__h�`�eY��g���rH2�p�z���.IXr�m	5�M��ru�`��Ç���XJ�3�:���1�+#�(q�+z6A=mCEt�z�2���`�'(���YD'��`E2���+����l���+��nJ�(D^��a=�,��:e�D��tFH�^�Qe�etGA�f�9Z2�q3���(�E�!zz!��̙}�V��bdU4ѣ:noV �v�ĸ��=D�5�r���ۥ�췢�(��l��nT��G�"�!�w���3ufaY���w1u�o�a� WJ�l�(��Pr��L6�����.C�4��26ۛ{ŧH0�i[�m)�0꽮�rTrbrIA��T�s��=Ïq]�>��VQ�@�3��]3��d�q1�[��e�J��UEs��b�j--ї��8��\&��ۤ��jT\�3M�t�m�t�R�,Ym��Z�-.����\i��Z��c�MZ�q�%2!�W�kh��S��5CI�҈�ir�m����E��eˊZ\�F�C,���)n�䢢�E�L��k
3i�WfZ��-���㕨"�C���lm4�^5�u�ԹLl�k�Uҩ�*T�Ƣ��*�����Pb�j���mU��r�Au�.k�����Q���Z�b�-+�D+eac��.R�1\�ª��U2��]k&E�,�,M0jŬ�R�*TJشe��i�hѤ���mkXj�5�e�M\\��-��
�DX���@#�����{�ե=�7rE%m���)ێ�z)���J1�>vh�<��ڢ�FG�e�R��A�ዙ�Ҫ����.�|��7X댫1��j��5y�x�g�&
�=5��E#����FOw�؛�)���A�rC���P��u)�v[t6{�B8�zJ{IQUt��34����r�VE�7�<�{��u]>E�N��Մ��K��ݞ`؅�/{Fz"2֗{WzQv.*���Z���s�#P�K.bz��񬫷�V\?9��t&�fRj���)U�>���7��b/��v��k/��0���qr@���F����&�[��B�����.��kJ���ѣ2��ÙCb�QUdو'v*d���m�S*��/�4���G�$ȥ\�c9�����U��PWC�^H�2LY�E��;�k��#W
ZYF*��3�)�^�}˦,k͵�)R��'k���x%9��F�K����P�զ�Wt�S��a,��Q�F���{���u��ִw9;C����fy,�YU���<>��P��Fjp��/�;*��s��Z�������X𧼢+7@3���#�� @	�:7w�j�w�mP����f�R�ܑ�pt�=6���4�Kr�T)�M�Pz�[����c���wx�n�d�u!O�	�\P����Ù�:n���rE�_gf�PDoQg�3.X;� [�X��[O�����\�=vʇ���<�^�.r�}�l�҃�}���ѧ�H+")�^A>rGT{��C!�ex5D�]ڽ1�s�x֢�1�r���g�:F�Azg��1��/)�N=�Y��U�c�;3����]�@�i-?9�a,����[��A��<s"0c��{Ń�;y+���gGI�r�ӻ���o�1C5g�$Y��d<=c�Ε��I��tOnrq��/һ�ւ�P�+�⧛�,h��ğg�}����CU$V������	"t>���Mi-�]b�!W�[�w�_���%�����L)����#��GN���'7`^7wv��mXw�,�劽���
�R�@�˔j��Oo�GO���w6:�92mu�D��"<�:�H�8\��7��`;7X��Q��?b�%��RC=��x`�q���ty�51N�	�D#=<QR{~9'��wBw�������m�g*m�M`�#G��n͕[��ǘڋ�U]x�{���H�ώ��F��2����X��oX�	�b@�60P2z�&GV8=s��K����к���}��th�Fhn%����O0���ƶWV86L�,5W�DP��t6���`��k��,���9HV�S`�MѺHD�U��dC'�ofV&��ǻ�8�Ш�]f2f�]�x�7=/$��2eҺ�y¶�f[�����c�z��h4�cz�sæ�Y���N��n�d��t�*�53��]s�(z���,�rg��]�i4�:�v89v��9��IdTj�qEj�F�Ӫz�9F����S2�-����I�)�D��-Yb��b��Ӳ�Hc�S=>�L�Z�^L��N���HaΩ���W���Q�Æ�Zj�P5������y^����hT� �ؠY�cf��O���]!D������[��sh��@ו�t+���94��d�]z�>�v�Q)%��1�U�!>�G�12�N�q(Yc���I�	HK�M��}�$�)�V���d�w��" d_�%C�
Z��A���p� �Y�>�ύr�;PC[�i��x�'�r�N�$�o��71���Qo�`8�����PO<�Q]���d�$3�����Փ[4:�D�<��s����<�Ty��b�����AV��X��|1�]�Ҝt���W��N���&����U�J[ve+��U�l�OM)n�+D-��Uf��,��{�C��^�Y]o,R��wHt��(+������eG��^��N(@Pf}p�FN�^m8���'����V�mΆ9P��*o�T�Ǵ@QP"���W��.,�P#S���N���Q갰��E�����dʏP��&�`�s�٭�7!�����P*���1��hT�kF<A��\�*�έ�+:�H�V��@˞2�ݠu{l��t��^�:W��Jˈהj�cFj�r���aU�K�U\��� p��[ӷ;�v*g���/�: ��0T|�xW���
���u�<T����unr�7nȳ�tb���K�3�u�q���JL˾qjn�$���@�!C�y7ȸ�AR��Tf�E���. s�{�.w]^�(7�ۤc�0��d��A�U�jn����t��f)8��}v��m��q��2���^�y�XC	�nI�$��HP����/vw�`�����_E���x:ãa��+��v˖5�$�w�<H����l�r�#�at�k� ��{�=⽓{�W  ��_,�\)�P)��7Mذ���
v�^i��ߡ��������Pܼ6�^D�0m�P�Jߺ�eZ�wP��]B����VUŹnR�y^o"�;��2�΍G�_�E/�B�{�M��{�7+uY�C|�H`v�V��n0�H�)�)Q��Sv��]���oy�|�]8D���[C`���>��EȾl=�{tg{;��^�Y�`�|�_S>n��C����f�nܘݑ=O���!���1("wO]5����TƇ�cp��M��4��z+��;V=T�i��/P�W��*�Xk��Dj�k*ی%�s�b�E.��c�Z�V�K��I����Ewl�Y�r�w6[�8��5�:L�1f��<����GR��YX��#��V���˙���3�	������n�ĨP1T��錮^lI���@�>�Q��h�oK�YK�+¢KhI�5�����[\���Ð�z-�C��2�e侸g^2��w>ć9~�~�u���d^*�95B{�Z���9�<4a?v��*��ʈ�<5��錿D)�\�(���.�	�!�)�`r`�A�2�,�¸�4�p�Nn���u�,8�dPp��- q1�Ý{V��F(�z�s�WA��.������Qce
�1��qJbo=O�Ou�t�RV�.�9aR�nJX�X�P��P�2�7��pv�M�V3V#���y���Jv����uA4}�Ƴ��v���ze���h&'*p"ֺ���,�)M4ٻ�޽�����T*�Ey:"+%�^� M:nv
@�l�Ҕ؅�����Z�j��0� O��t�BYC"ۯ�l�`��OcPs�����SB���
��TV�c5��0�aoNv�\K�Q�lq��	�.�f&�:��a�+��O9��/R\Z�#��`թ�
��C�u�zZ)���S�����f����{N��f�Z,;���U�8��Uȼ������
�*�U(}��g�;q��ǆ���xh9�zǶc�gu�cG��Bj�U���V~�k�N���5����'̤v9	�bA�T:1�r3�@�ʷ?@]#��������3Ϻ�B>s����O�.+� ���`�5��h.ᶦł{�4`n��v	g�hb9�I��n�Y��.�ĵ)(��`��]8l�뼥w)*�}=ͭ+��v-jL���C'��+�0��9�'�üַכ��L4X�j������}t��
��{�X(vb�$���E���v_�F�ǎV��Μ
R��Va~�pW���oy1��3�j��N���;��p$�@gP�:��I�jC�K
.� R��1�̈�Yn<��ra�x��K�]M��g5�:Mlx�"1�bb�e��Mȱ����J�5�d�ނ�y�����_%)`�F�%�YB�;Q{.&���Oy0� ��]4^/a�D�>�(���{m}��|�ݛ�s4�{����c�z���\V��Ѣ���K:��X���
�A�i���j��B����g���/��Z-��;@y�=����r�����u�Y]�I�\b�G�99k� �ЎJ>c�d?��}֗�&���KH�5��r��73�|��Tټ�'^���omd=(f̧t_͙�Q�Z���{�Ћ�f�����c�4S6�-U�:��(�*�u��
�g3n:�Gڊr�tʙ��U�.��M�F�M%����������M0f�K8�Qj�^�ʍS̩�YW��nnVoFz�T���i��L%G�+��+-(6�Ǌ��6r�74�Vi�WIi�amgkĳ)�b��s����-M�o�+[51\�9���n΃�P�n�j���ʖ�+H����U�>���HfĶ��W���U�dTM�QH��ss��h�i�8E�� �u�ҢQ���.�Y|O� ���7juV�:v��څ^*����p�����t�[&رq�Sb;�t�&��������F\��-ԝ@�Y�&ʲ�p�NE�t�vԹc������:�XW@��C�V�V�C^:F��4v\SX7{r#���T�T`�y�R�r�I�~�ެ���VSهͷ�����㬯g��h�!&T�=30�y!t��%�����H[*�K�J��{f'E8��7jziV	0��q_r����q蓥�U�1��Ї�2�r��ˤ0�g�"ج���j�Ӛ�n
��d류m����,��v:w��A�CX����1鰦n��/5�qB+n}6�k�:��2I7y�m���i�8�`��v���[7�7��Wv�yÅwg��|��x%4�sUmc�(���2[��Y*�m��Yx��/&�'��������b�ö��{���k�!�Z�*x��^��+�i�+S�ck%Ũ2�S�"�:6���]%LW�K >�P��[�-5n���VV�o,W��t��3n1��*�㮛��+����OR��]���F���Œ�N\�wI 0o}3��H��>�pf5ֈ�͠k�L��Ø/*5G��C4��[n�V�9��33Z54XT�Қ֫�譥W0��J)���DZ�Z���X��kU���C��Q�Keb�8����ĭ+n�Z4�A �))�E�"ZIB�$�nIX�F�%Q�P���*�(��[m*%Z�L[r��S�S.DѪe)m"�[(�ie�3Q��Nj��F�r�DFi�%
��YXZ6(�+*���V����+�V
ڔk�&"��FVi��cY��S�L�,QJ���P��R�2�8��I��Ud���Z�Mep[mh�+B�ţ@��{��/�����c���oe�y��(-*�Z�̞�?�j�<�������/�����������[F2:܀����.�X�K3rUs;ũ�$�{��D���	�G;���}�~�0�?��O>�m@Ⱥ��:����w}L���볬0��ۭӽo:y|�3��[�Ez�ל(�F��K$l#>�6��" 7w�ze��I�W�WB�ҕf�Kp}�m����A�0�o�_��eցB�}�.�G]ND�Р�C�q� �ص&Lܛ�Kð�#a��D��QY��%@�P89��07�یj0.?g���]�_t�\~�U���O�4o�]�.�F�1-�x_��u[�j\-E'�h������Fcޞ���z�B�R�:,h�fK�{`���=�.:E>U+�_dпK���i���ԌǈgY��E�KFRү��ʙ������OzQa"��+�'
�, ��3z�C1�A���^oQ.wws��XZi�Cꘀ�Ax�С ���JT�����=�l����DX�~i��U��eZ�C4���_�^Eh^Ğ��u�����@[�j����c/(��u�>f��&/f�X�w���<�ss�ɖ�Z��(�ZJ�� ��<�8�[�zSj�����T �pB��c�
ˀ|�h�r�j�O8Sk��>|�`�����E]V�>��/q"��ϔڒݷ{K	S��͓�h	�冮�lGF�k8 9G�^[	��	=]o��!�e^߮4f����m����ĘHN�:3���!�>
�k�uW��Ms���xօi�|�0c�R�Slvt�l��dkT$)��'��yyTGa��pº�d[��q�.'(�=��T��qzs-�ʜ�1���7�r��H.�,7*�|���{�z|�봓�v�8��G9��jއU�[';ͦ�-\VxJAB�s��$�=5��~���8@1
{�U�=p�K��:N��oDGf$�ʌr���a����4{U�8�� �t�LL���}�ܥ3�P���ʊ~!��8w+���}���zY!�����av��a�8~ξI�*>�޺ڰ�*3�����jշ=!@=)HUQ
�f���2���9�"ECګ���F�w�C�"�8��d�Krgz�?!�E�U���Ƭ2km���<�0�/7|�;�v^ibB���	���WH��s�J�x>��A��8���f�o��7�W��g[�N'�P�Ĭ�aB"qv�T	��z���E�s^p��%+gǧ��
wX�����me�e�5�xs0�z��R�-��ᮼj��FN���3��l�ֳ3jo���>�ʙEw��ޤ�xz��=�mLM�}j8�n],6�5�QkG	I��L9p8�p�G��l}�o�U*��?X�,��ǆ�b�U�u�h�%mlS�����@��O��ئM��Sq��^9c2"�"�s�ys��G8���<��=���{�˺wɕn_ݔ���w(mI�WO�c�"}�����TMo���3X�'eI�Op�w��ɺ�t�P�4�X]��HX������o#G��x��p�}�U��t�( ��:�)z�\��T���|�=a�$f)��;�!�,ZZ�Y�Y�W���LW +��ΒU�S���<O.��
-p0��R�V�%��a�ɧjz<�T�2/$��Z�����@*��ƥؑs"#���??G��/��5o��??z��rF���@B�L��$�*@�ElM�g�p[��E�˅E�]h|���={[�!_JR�������1��]$��]Y������&�U������M͍�(���m�e1C�PB ���U�k������
��Y��s�zҁ��JMCKń&-�N�����t��#�7���Z=��
ەu�R��R�בN}qC����޺�_aҊ/4�j-Z��4�^C
U��.�MN^E1�9��RaQe���}� O�mt:Qh���5F��PVa��<�d}�r���## ,c�DP��ȕ�����t[���<�gT�������0:�\����RN�0�Xi/���8k�k ���ϕ��#*F�9W#aG��$mHE�Y3{m�i����B~a�z��V�jM�7V��XhɎY�V��X��~
`UoL���^p�`�0˰�ub�[�q��zF�YC�9+O�6aODh���_�ö�Lu���Mu]�٢��f�y���-s����H�����vt�C�I���6,�����G0dw3�vr2�	�Z伢�*F���S���8e(
��D�q=e�=�������� V��4:����S>�ʡ4[�NLl�,���#��K��G�@�4��PP �C}p��x�dc���Q���V���ƪ�nÅK^�T�y>���w>���:c�V�!�����}�B��\έO^l��]JC8�Dd;�]�n@"O���T���="κ[�N��u������c,�$X���<)���.�3��Kna�3V�Fʏ*�k�'�����V��To��}�LtJǨ�1n\z�~�e�0$p44D��R*�{��5� ���eL\c^t�`���O��:+@U9G�n����;(�4��ߛ-�ז�>|�Ĕ�:������׳��Q���zܮyc�)$�W,���� �o��>���n��r�-�������UqI*�0�R��/認���*<lFkF��2���N�27��d�b`��m���<���05���Fx��bxs6�ȭ�� ��`P`�u����aF ��c��{�#���ԐX�=t-�R����A��g�htXv�]I�Q����񴕄zTS����4,`X!�<�@n� �DI�p�|TmF��'.v�S�>\YÀ�@�j�H8��p_�[��J�{]#�B�-Ɉr>0�n��!��\��󑟀��h�����>5@zV*5P�hSW��}��:�iTĎ�w�.f�l��Z�&�7=��+e@tM�_8wƏV)�q�� vX�I1���}��!�h��FW�c�;M�$s+��3�p����D;fv�/uR,����Y����1����L�� R"�kkX���l`,r��nմ�Z�+nCo&>������o��Z~P�P�*�p���E0��Z�5��v{:/��&GEFi��Pb����y�X%�5��^T�9䑊CΥ����w>�)W�Q5]�
(p#��}A�����+t���U�@�2k�΄�f��_`�xkEh���{��J[�z��|��#��s�=�9sB��>�8,Qجxp��Pkw6�&�TR��V4���~�P:���+����l�0���n�_�ث<k����
�%���n��hj�Q?K�'u_i$����j�Q:����.\(Q��Hgf'���Rn��`���pA~�p���l� (��>�H�0�>��\kU�e�
�EP�<<88j��9p���K�Q�Y���w����N`��="�,3�˚D%��#����G��n�5�'�/m�]����.+aT�r��"7lcwM�]&�s���W.�<�P]cb?��{i�����93=�4+� #62TZ�~���B-9�v�{,�o(�r<B�]1r��Š_���Q$���]-E���z�ّHs[n<:/�B��w�bb�e��M�#V�Cla��Ȱ��J�8����P�f0�q%��S�0�f�#�Ϧ����/�����::�M��S5���!��g�ޤ�+�Y������f�����b�pѢ��&J�k=Pu�0�=���x��.3M1�vk�T5���U��+F���﹮�ζ���S����.Fl� O�yM��WW�s���_4�Tц6z;'ў����0�b
ϙ�?w�AY��y2H��=e$�t�X�� 掱Cg�$J��+ʶ��r�1�d���a<�Tt0kOs�I<���En��u��{Ӻ��z��ߝcT��d�Mr����y8&J�Ϯ&9�é����sK���qos5e,�y:�6��w)W| ��i�{'��3�!R�Da�0�%b�0N&M�C;-Xuv��\���<�8P/}#c���χp����,�U�KO��B>�l�zT��>g�_��a�
�<0hx֎���u�:̝���C�P`.7at�*'p�wv��F�?@B]8�����ͅ�Cc�ʲ�p�)��<���ۛ��J�����n
�E�p��5Õ���r(L��j���B�j}�A��l3���4HQ*N
��P5�[�e\ǝK�#�Z�D�D�@!k�j�W��5����K�~�Wb��;W�˗�N�e���!󾻿}y�rV�܊����2z�qq�nۑ���+��W�~?o�Nc(�@�'�R!J�.�����rN7g] x���#5(6�u�r��v��֯���c�]�[� �,�-�������swi�v|����,��A�I+
��VT;!��&n^@��p&s���r��ipnv_[I�R�f��sw�0��ݕj��72Ա5�uYp�|�c�EǕ2�5JV�%�`W:�d��F�����t�P����Z-AHv���[3G��]GsN�ST���<�ʻc![��
s(���+�X�����j�\�� ���f`��	�w�1�X{��h�ۑp���ʷl�ui����#A�m���ꓑ�=,'fuq�Fq�xӱO.�vp��84�Gk��.�L)���5�
ѭa[���pi@���J��Ǯ�p�[9��`���e��Tu��[�o�9��`}k�8.��
X�Ïa�2�IÌ#s���=�-lE-�=g8v�n׷�,�������,˱�-+mr�Rm�8$9�_MC�G"�e��gV,��)'r:7w1P�WiЮ�#�N���#�3V@x�]��蓷w���:��P�(Y�����h���Λ�1{�[�#p��[�䙴h"�Cg^ù�D���Mcv��q��1_G���S%D��ƭb��Սh����ҷ�H��c�c��	��-�-sg�R�5�Jy��NAN���>�y>�v�Y���p���Tٳ@Y{R�;&A����(�l�O�,��(�N�@�sv��5x����k!�g�|,9���lk`W��W6��m����?��PW�9��B/IǐV���6We���!ɕX�����11�nWJ̧��[p�(�uϷ�5�.���ǃ�IVwCS2���s2Kb7��@:�J�t

����
P�]9j �>�����V���@�%F+kkiFإm*ÚP�,��,�V�x�aDI��+ZZX�,*���kF�T�b��TD]4�Ҭ�J�QҶZFTF��LJŶ��������b�J�Z�(�(�i���j���iJ��1f\�J1�X�J��e��j"��f�i�k
c0�+,DԥQ���Kl�(#2�kTJЪ�am�Qil�E��j\n
�0\+�X�Z�(� VT2�6��m̲cX�
��Re����4�E���[�Y+��R���7
(U�:AֳV���������Y�z~/��*M��pд��ATU���=�lr6Ҫ�	+��u�E)^���xx1�[�C����I�8,��m<���)��\ ��X_F���h�@wHc������]�=m@�ʰ`���_72˛��T794��� ���h�30$z��
fٙ~�,�Y��~�\�F)q�vL3" �ԾU��o5����Ɉ�5�&$N:�7g��ô9�� �Û�&�S�q;��Ad�ى��������qݓ�%q�ή�η���x�}w潎QH(�Y6ʐx�Ձ�*�2T��Y�`p����v¤��b���IY�1�2T����錏0�3[�b����� T{cӬ�!�a�6²m��v�Ϛ�T�ő`z�a|�+�=��AH.�)��
,�J��*NM�ă咥��~��9�{���}���]�a�g�1E�aSl:��$m�P+�T��`Vx������J�AHk:ֈ=��n�G��#� y8�oYy>�t���Ȥ�K�T���V
A�hx�a��R<V��E �wE&$<Im�d��:�I!�̞2T��y�7׼���߯{���bp�|�q�4æ��x�Ι+�cuE ���l���<T+��+��4���hc�V����.ܮ�yz�:��s���[���e�R����曺76��Fmnv�����z��z�v2	�%؞��I���H4�nT�Bͣ.N�h�3{�YSEi&cr�j�g�����^5����l=a��ŝ0�AC��1�2VN�TP�%t��)�d�=ót0�a�,7�Ag�8��U �8C�Û&uHV����ٚ���7�� �o�c4�i�
/`c'l�k�LH6ɬ�f����wm
�=�b)XV6λ��Adά�h�V��\���	\��G��~�� "�����a��i
�0��AgY1�$�Ĝ�"�X8�i��H9uœi����wI���+㝽�>���]k���}�~!�*AM�@���=�T���+<d�
uiP*Ag|�18@��ca���i���Y+ǶM�Ag�VLd�z`z�o��#N	ϳQR<&<D{�9�H)���x� (���La�
��*A�C�l*ANy���%a�l�P�%xI�Ă�5�{��,+5�����{�{��q�Ag��� *�J�X��u`g�CS��<N
E�����w%eN�*A�X�f��Ɍ�=B�^�9���X�.e��}�������h�Xo��
ÖpsM$����1E�xɉ&��)TO)�0�)�s`c<I�!��)����s�|�9��7ߜn.0X,r��c9���H,���b�&�6bIRZA�Ͳbu�;a���]�c;d�;����,*`;>�M`?[��u��_o��,;a\a��M$r�[����QH.���OPR=R���H,}���1E8恌;aXk�H:��8�Y��T����˜�~��~�:�1%g�����C����Ă�Þ��!Xt¼j�ީ��k$����*A`j�*Aꐮ��&�
����22o��x������/qѭѿ����{�9(5�>o�P�9�]�e� ,DA�Y<�#�Il[k�N1��ޤR�*Yޠ�ĺĩ�r��hZg/a9lG�Hmb��W������^���� �b|qt�Rt�1fӶ�Rm
��v�$�u�*H,��&yE��d4�]�kt�<d��v$s�~'��8��}�YH<�zqCL8a��=jAgi;q�������ۦ �@�1��P�[���S;��Ă�l1���2�H>Y�L������zѼ�;��w$Hp����� �O�N�xΐ�t�x��!�H0����Vs�������kZ�޹�y6��!��a�,*ktH:�}�����LCi+=d�u�1�W��,�Ag��u��;gF餆� ��J�U�_.�zoo|q���zN�
M��ăՁ�Vv��R�VV�!��&$Mn�H);�$�Y�x��
��+5�6�I�2��@�~��-��\{���Hw�
��0�Aq�����J��S�����Rt1&0�7���C*L�9�M�R
m�n0X(p���ot��o�o�{�u�=�����%H,ݲ(z��ÛH;�k�pö �gl��2T�I�PĂ�2jsu�!Xc
�퓄�Af�f��
v�ߚ���l����c&�lĂ��kۤ�i
�՛T4�Xk�f����*AaXs;�R��ö�6�Cĕ�0Ѫi ��zc���5=�y?�����ﳫ��t<&!��T4�����8d�]��P퇎$�qݚa�;L`vԂ�a���TH,:E� �uֽ�|o���{ߞs��[�,��=NXl�H):B��7�i ��d4� TR��W��i �'Y4�Y*Mn�>�+G�ZA�v��4�2����X�=4��F���ͻy�+2���wc���SA�	xS�`��u�6f歮4�6��efc��.s^Giuγܸc���d%gFdp��u�<����&��x��=�[&�1Qq'�QH|���X)��g�0�oPĂ��)��RT5�aRVh:�bA��Y�a�
����2W=ַ�u�������������bAJ����
�hrwt�N
h��&�Y7�Pĕ �s���A��
�S�
����l����>�L��yߝ����6p�R���<a�XVrwd�=IY�9CP�bcX ��E��y�*�L4���q�gl�u�b�R
zɷT5�n�4��u�����&2{Ř�Y����(��٤�æ�%b��v�H)*�y�b�*,*m��(bA�&��a�
�[^8�����|����Ι*�Cz`VNYR��^�
�L=�t�R<M�Ӥ��E���1��X,4y�Aꁉ���1 ��e�3�IP]�>����<y��ǧIRWL
�x�\�4ö&�����������Ă��H�HV�ُ��&$r�_Y;�(�"�G�������������>�3z�T���Ι��aQH,6k���
�r��ö����=IY�였��I�wCO,
����8��:X�0z������0<:��%gl��UT���y�<jA��j��3��j�4�R���R7�&�R8d�Y+z�=�@��'�/�5���߅ǫgި B.���N�*AH;��=���Vmk��J�E�C��ć6��/��a���h��S�Iˉ=J��3�xߞ�C�-`������aߖH,��IPR
���i �yE�t¡Ǵ��Y�5��=�H)�8g:��=��b���Q�q�!��W*9\���u÷R�.����	�eK�E�O��\�fR��(�6�⮥�kl:��w7,�{Հ�_	�1�����Y�]��=��HT>'Ua�L�&2q͘��_=�q�a �wa�i �`��=T*IR=f!�P*)��TXbAI�,=a�<C��x߼q�>�����Ԃ��*���E�0+',���� t�
¤=�ߔed�0��UH,�ٌ��9�V3I��wdĂ�'^9û������ǱNP4���T��,Ւ�g^�l4�Rt_p+5����4¦�+��(�i1�aY;:���GwH
/�
�p�^�ǻ�}s���6Il7�搬8N��R<̝$�Ğ%E��ɌZË`�P5�4�{�Ă�-���IY��b)S]P�A`=r�/z�^�Ϟ��=�4Ɍ4¼0*Aew=���V8�I!�f��d*j{g,4���cMXc:d���N}�B�R�fI�T�͜�4��B��ޯ�]��s�<��]w��l����iE ��l4�P�%�Xc<�P�AB���x�PS�RW
���OsܓL���9޴Agl�:�{����x��ݓ�T��s�`m��搬=g�����YO5��p����(c'���R�J���$8��ydĜ�"�L*m�8����[��:�{��Z����/���F)q�Xvu� 8����_+J]H�� �s��>V|У�o�S����j�x�I�f�b�6�"1H6��s�*���+�0&T�{w�L�;�!}�TD}�y2�:'�_�0}�����@X���d�M���r܉ud���^M7�.�O3�D2�
��Ɍ�ͅ�R�%�t�y`�U�/{f��"V~x���y&�f6_D�W	��p����]+��^�M��m�J`d;��a�s����"�
��kK�#�1V^��Ǩj~�x
!T�**����v�� w�H1{=K�v"=͏n\�r>�GŏY���2ҿ8q�`��z+�Ff4]kԉWudFM5BԘ��EP�	Jrc��B</�d�|:�������*�8~��R�fԸ�9�t:�����խ�-�������t'D�J�E\�>�tۦ�`/gk��̜$�% dg��ǅ`��1�ƾ��w�G��d��{�e�|7�'�)�G���I`S}��O~���ɵ~唵ePB���hظdt�#�O����C�|w��;BV['��Ҿ�WN�4���.����&�0�`�'f�鸥�cώN���m��qE:f3Gq�%�v�p��y��v_��	���}_UxM;-&�f�w����y�S��BCT.�Z�y&g��Eq��O�� �P�P��ܼ�P{�D��h�Y1x���7}���S�V�~TN���$`r\��OEd�3��Krv��<ʸ0���dQv����]6�<Eْ+B�]�z��+�n=�+��}:(��6��#pUN�{'����x�d<��sP�B��x}�|��n�����X
�O�{�~"��^!R�ѯc��)�� (0a����U,]Ż�\Ñ8:�4�ՃÇa�~��g��.�n�*y�%��Iu�t &��&aJ��P��Ƒ/a����ł��{��Ղ��	��Q$<�.[8��
����g�Y���+�v�L����wK����ӖP8�	�RZ��/�k��#�����}��>�wE).�(�+u�cƦ��J���O�x�%[�J1�dIT~ xz�E�r�����+��*���&�����=�J_7O5��Hmk����X�Д���OW�D�x�|\p����Z;����C�I�z��ab�a�Y����xi��"�&Dt��s.�^17j�yU�b����\Vx�U�E0��{Gκ��I.��XG�Xa��P�A�]��gJ�b�S��e��^O{�V�Y�.P+�M�(8T���h'�Q�|k[�g\��o��k�z����e�-�^���V�<!����-T�W��/|C����Noi�=`���D}T��x
�F0��t��M�w��Ð⽓�B�/+}
�°U�*�`����R�e�j�ddPr:�tnH���r2�9W#!t��aCS��c,�P��cF�U�H��j�&���G�.�w�B�� ^QIf�)<��3�I��:^���Q��ŵ6ըI��9o���2��W��xT�M~u�*d%7S��
%�G\�.}�Ր�S{���v��R#`�¾�³Ԗ�ѥ\~~>��]�l;أ�^���裖~�%��mXb&�4��t�cP
�9��n��$h��4��O�D�\1����B�%N��Ǭ�W5}��lJ������s��V%[��*��t*A�i~��<��e�0��#Wr�['�l�g�d��gMF��$�j�j��T�@IW�J�q0� pو^�19O�t��%d} =��j��xU���%��5[Cl��j�-cE/@���#��nV�۽"-_�w�z�i�|��n��-��X<u��/��i�sL)���if�F��:��VR~�9��B�C����^�P���w�Vʗ��#ii��b�2�P$�P%���z[��b99�cd�����(΁�y��q[�,�軕��z0��  z2�6�. ���� ��W�
 0;��CDљESW�x{5�[������~�eXp��ڼ�F)q��a�W���S�0���X4)�ة"��F�%Ol�}�^7�%�F��&�����ԋ�Q�,9q,O���$C�iת6�2�Bqx��s����@}=!9��G)��c�:��3��fN�����+����aAFよժ�B��]%��������B��͸$tmeS�*2�(�t�[��$�
3xa�q�3��s*�u;��1�kì�3:\���h,4+޷W2��m��;�Ȏ���4���WA)X��9O�v�xY<�Ȉjr&���=>��:DH�͹qj@�}!~l���'{�6R��W�qN$$�K0]EU������� �i��`��7	 pV�7�K@�&9��*�k�7��h�������Lt�+�#M��l&��D-4�z�vF`�+�iT���[�Omc`���ܷW���*��7GŖ�į)�"�E�G|v���ӯ���c�"�)y��1f���H�[�j��ͮ�Z�����t
w�I�6�\�F#WW1c�W0�v���̓�d,_l����t�J�CáYE�1��7`B����ì�R$V�3��H�14+�v6�u͓�{�̜�F��1}{��.*]�l},�]�8�!�
NX��ƺ��O0�NJ76%��
;T�g}7�'V]%��u�uaJ�M3f�0#�s�d���!`
Wk��t]��^}Cj�i�����j��	usA���d�b̫��ll����$��]f���]Z1l�ݲ�� ���P�C nnX�z�|���  ��-^S6���/�Vf]kN*�R47�+Sl�y�77�t%�=A���X��#ܩ]��]d���JP��}Ɛ��&7�����)�i���u�u�;N��ǔHp���;�>�k�����ʱe�3�$7��|�l��������o}7��7�2��|A���W�����	:̦��=O:
�f���tYR����`�/��@һ�@�e����B��:��iă�]w4�$�h�S����w��.7G��v��upF
x:�/%�S��ܕ\ĽФn�l+��`9f��*�)]H���R�[��Bo/���('G��o(�6��k=��"�?jH��j�m��[��1M`҄��r%��T3rv��˂�aT�6٦�ν���;WXI����	�*qj8��Ԛ��k��<�ގ�Vc����#�#fs�]�YN���L<�VN5y{��2���=�)X"�'�q�G�3�eYV�*[Ec#����n#l���qP�ic1���2�]&9�.S�f\1�ӥA����1�2�V8Z�r�)dKDVkj�-�e��F�bTr�e@r���ܕXV�5J�8�ƥ+QX����&
��G�U��+��JffI+.Y�8�Jֲ���pfT�35�ѭa�"k)��T֍f������6�l�c��Vi�HWVP��`Z�*T-�s�c4�&U1!�bi�
�s&\Q��,1���	J�����)�޵I'Pa���5��c�tt�k����n���Bd��+�=��N��m�� �3�Ρ#D���6,L�M�^� Nzݷ<cF�m��{N8r �-�'L -aI�&幂��E)Z���S�^Y.+&��@�i����J�U���jÞ���c�H���u�w�q��T������@���@���糷za4����C��p�^��}^V�Q�R9	�<�c!-ǭ�ճ(G��
3�]�9��qW#��}^����{�9�j�g��#�,:Uj!��81Pk�����~�kN�M�W���׭�_q�E@�b��v60R��T��UL4Q�֋C�c�>S���m��]
d����W׹3=v�j�G����r�[�t���c�Tj�D�;����%�艠�F��$�g��5�v�_b"�=�HY3 �#�����`��𕕉�F��r��]n4�aK�7%7�L=]"b���''�M�J�`����K]�6�j>�nk`\d8���90���X�JE�Qy/2g��]����ߤK��+��ᶠ��,S�G�8e��ss끒9u��U��@�#��6EzfҟR�c� #9
)U&��F$�{�EzXC���k�"�#�LZG��S����OL�E�r"+���b�#���z+��!�ƸN�cҘݛy�y�(�zC��1#�n+C��PP��U)`�J���7{΀d��3Kup~��*�Vi�øi����Os��#�P�T�_x��v�f���[.W��؎����=t ��4�ۿ�)HJC�"@Q�����
MB�/��y>�?1x!B�hǈ3Bq�*|��3[B�Q���)�L2 .7� �"���۾�u�g�5��=ΥY4o��jJMs���u�wj8����V�q56�[կ�5���A��Gyw�W�W�m"[r~>4��f�:oez*b`��]m8���olN�{�`����&�sC�a� V�G�X���8aƉ0X�m��o�k��`��pu��X��Jv{J2�W����1��j��i�&��X�5ʞ�>�k�ƭ���H�+C�9��7����Q
����^��Z%��gݍj��6WI���ǩaç�,,���bYJ���
"�ԡ�-���SB�ҩ�_�%������>�I���ibE�W�#{��A�`�pI�@��7Mر�,EG�O��
د)�d�,�.N�LUz@��#�kȞ�<�_1�
�]!�;P���JO�l�婻�9�C��ǫ&��r�TC �U�F���0^e1V����*���W�5]�u�>Zo{8an*�[�z��H�r Y�&뇸G�k} '��C4l��U3'�Y�d�%�.�vMZfT�������]��y�R�J�+�B�{�?���V�j���Z����r���,������l�nR��*.=Wj�r2��U,���>U!��iA��C�MQ�@�u��D��5���m�����@�B�%[`O���蜑=�QBg��b!��m"��1{AE�5���{1#�aX�.�M���i�+J��1n��B�"�\u�y�:2)'�2������!����PL�W�.;�Q�_k�I�i�/��I�70��r�btp�LfH�
kS��3��2���2��o���/Z�!c�q��5�~�+���]��9w���2^�Q��P�Ce���	��a��Z_z\���f��i
��PN�u/4���Zݬ[[��2�t�*����^97�	n i�H�����e���+bkLC����,3��fs�7�������v�Mעdd*4>=���q]>��np@BA�$p����N�%J%������K��C����Q���;
UyÎ�A,giuO�U"��HR� A�P�n�\{"�BR��.��n3�y�}ިIÅHC
�\X�"�38�ũ�G�s�8�S%)A��^O��T�X~t�}���=y��*�$��u�� ��P�jn{���wC��|h�D$d����-�x��)<$S�sT<V] �b��6G�n�7,��#�!.{2�y�V�en���c�n(4l\	2+�DW;���\N�M�}G��BD���=5l�v�G����TԊr
����JO$��fi���<$��c⇯��׷>:��sȉcA�4�^WFJ/8/-+,�����^�k���-�T�ѴB�8��/�P�C��ow1;+1�V��qgwTQ{L��6�U<����=�ì����k�,6-���J���x}�k����.���n�m]�(��ãC�P7�"G
�غt:ꀕ!w)VY�k���]�N����۟yWat8,��qG��l���I��:ZE@S&<�(~9r�O�N9��^���>��;
$���g�x����I��¸]��+#�uq�"�/H�qZ���l�azGD#��U�~r�E�dl\y'�Tp�gMbm���}�dv 0�/�٤G�Z������}���c�mz\� �cz�Ԏ����Pg�C��f\'�9��^ȃ)���@Q>�
k�}�����9����R�a�劾��X�^Z�	�i����/��{���x<�ҼX���E^�O%���4k畔\�xc���Tb�9ɰv�Nᎌ.P\�u�a������uev�������2W������M<q�
�|��T�˃��[��٪����͔TN{}�(/�W^�n�*ϥ�a��J�(�S�w	�5x���B�TC��TGP���	q����P���<�������rnnҧ�U�
���
��tfV �#�*וJO+m�緓xӡ]L������?;4F~�N�pm(�/�A閯4�up�CT6����R6�X��^�p�VV�U-�o&�mC#���(OE@�7�֠P#t>��E�ktd�
C���kG
ۧ���,��5)/��P2�6�Nˌ�r,G�@�(D@.z�ղ-�)��r��s���SV�9�wJ(@�./�t-:+��-��IP�����{�|��;n�����xyD������x�<�����f=��k3��Y�EcBvn6r�n�&�r���d�&��޳(�ǝjӳ�(��cDqn䘿>�{���4�;��ʀ]P[Վ|�\x�� 
�M�+�k[6�g{�p/|"��$��P;�F���hR� z}��(dPJ��;�;�k�2]z�v8C�옄�ßs�r%�l�2;�3���'	eU��$0a��\+GξV�|}��@���
�~	��E����^`�G�4�e/�<(j��qJE�&���#�����Q'���=�}�B����*5�C�Ϯ�7 �ݹ�͖�mn�>��qA���j/�4�� ��f#����Ķؼ�ߦ�tv�u^_�bگ1[Hc¯�����U�us����io�ա^����l5[��秂h�e��㼿x��JJM��*��e�>f���E�x֋�0/��\��<�T��}�Pߦ�ՠv��^K�Gk����,7�_�o�q7>�of�����Z��q2a�3��!b��V��͠��&� �B�Y�s<�)^�K~��އek-�f�@��b& �T�A^��T=�h	ίȻ��	��ֻ�W!�j�G��j���H�)����1��.zM�>����-u�����e�Ќ1�q�0,�Y��b�<4m�<렬vTov�@��Y~�*z+�8��̌SJz��BGL�P൨Ӈqzm�S��9�F���QPl{n۟ d6�dU�)6�Xb�������Û�yFNz�aJ�8qUJ/\�̤�4C�W	�qN� x�K�yaw��0{q�w�����x�l�*�Q´��w�U����^@�nt/l�
0�jJ�=�GNP��sW�b�B�8�Ӣ]��y�So�\����X̶g:BÀ��H*_ʫG]m��@���*�m�i-/qm.���{�[8���"��b�Ȧ�sE����C([��i�s{o��X�ye����o��9�4�	o+j2��Z�H���ݞ��W�������i�7~^:���P�T5[��8��&�Vh�z(���α�+�&�բǧ�wH:A���hظdgtd��,m�"#�5�G�©���T��3�-ڭؾV���n#cj̋���>��u�H�xF}�z��Au���~��Zd�r��P0�Fl�N�3f�!ƈ5S*�~��ݑP�'��l?t>
�-u
��hi�����*�IU^��
�㨷P������Fo'β�h:�K
��E�g;Tֱ�r����ʷtd�yڡ����s�����1ת5I:�V���Sٻ�[�^�7=鐔O@�r:���PtaX��t�7�x�kZ��g�=ˍ���!��):��r㦈�����q�1@��;g*XZ"|4�B��݅W`O���ɵ��!���$�VN4j��?�j�%Hܭ\u�4�E���ѻ�P�U ��P��,��c�Dt�{]�7�¾4 k��q1����;x��+Z���F����N�fn�n�һԢ.;9������T�c�޵(���g&m��1'{(T�/�a�U�p*�ٰ�zl�4����l+�l���eh!S�f��`a0��I&R�:�'c[�Z�P����G{�X���h�]T�"qt��T�/e\ε��F'K�j��'k#zc�aB\w���
k�f�] O6�J�I@X8���]�0���t�i.p��FrѨ;Jp�(^�C�j3:� 7�ȺZ�����%"�uA�QE�[��^�4\���i�fT�h-�ɵom�����S���{����[��q�,�A��dAM(�;��8ew�����k4Ve�g5%��if͓����bᲴS7�RA��ޟaA<�1�Cc3��_ҖU��&T�(�^�ڶ�U�XI��ٶL!��>вlf��M>�B+��Vd+.�ɏ�-º�&!�P3�[�#=���]v&'��/��r���hU×�1�7���2�}IP�[�3k\u�ViY�f�l�kp����YnY���ƅ�U�;/V�lD6Q����Y7Uƍe�:�Gsz���H9ՕA)�7�fX���]\6�ٌ݈Ŧ��Σ/\����go�����X�>����4�$[�]M�},A��*����c��,k�GB�Pt���wfң�w��^�Fy�$�mbo&����ٚ&�򷫠�8Z���#�*���t5�2�"��sy�x)x�A���F$�Q����"aE�h�10��tɮh���Qb�l�TV[Qbhlf��Tċ+b"�A("���2�Ea�����US)EY��3�-�QDkD�#h��)"µU1�Um��-̨���M��jc"�.���喴TDTE@X�V)l�E�b!m
�DV�1��Bҋ��X(�[V(�
�AUX�eB�J�`�T�Z�lV:�*"e���*�s

c(��Rk.(֠��E��AE�1Z�*Um�"��(���eH�DDAV�T��X[Q�[B����X",V5
�,��(�YQR�k�D��Z+�VJp,=#/0c7a�J�e��0�-{-��[*i������ {�׍sm��~
7��.�2'�,BTH���}��ǲo��@����8\��h5h",��D��/���)ۜ�F��e݈b��=lײ �|lH��W�Tx>�fd�ݩ��� 
z���Xx�P�hs�	B�1guP�l�����k���lR���f}p�F[v��q�jHD�0�y���o:��܃I��#��#����W��qc$p�t�0�VN>Λ���kB�>V&L�)h�D�|�|k�4�Ц��Q�Ξ��#o��]���y�̠if��qf'*�[��l�H.F��P��v/�v��W\t%��C�e�=��l�ÁP�ClH�E/Ѱ7���P�t�߃�.�$l��j�k�x��=�.�ڢ3��a��{� �g5+�n8�=&���[�:�!�nVd�Uelw^@�Or�=3��d��J�3v�t��_�j^��޴���ߞ�/f`p��f���P�b��HO��=��*F��od(
e�:�B"�A�w�c'�C+���`���z��(����Rp�!$QV�9�,$7�����%@�+W��B�H�m<0m��-[�n��J]@"f/\Dꏚ��6.B��e�]8��Ss�4ъ�v�	�k���niJ{�hW�}�b����[�~���
���F�y�b���Մa����0/%F�;sy1	K����Ojī��G�5 >��|���>�Ԩ�ZvҮp��OM����@x- ��s�򓽽Q���Eᤫ)}�	dwk�H�g�bIS��9��VWW� ��V/��B�C�5u�¯�H����؏��;�r����uf��6'[1h�i离�1���xl.�V˚����L�q��db�6���Q����t���g��� Hk=�}��oYƩ�ŝ�s�9��qu��j/�8U�0/E,���=����ИͿm�8��lx��Cj��S]";r_��E��S����Hk��s��썍�.�Cs�L��ҿY�Sy����3̾��lm"T�	���NMlX�q�>Z�Ń=^]�]�O��k*&d=�����@��}�CCAr�	Lq�W�e�Z0�כ�����0`��\+�@�")HUn�ڳkʷSLgl���_*����(r9B�Y����k��
�g��\\���Ʈz�?a�~82	t�"1F�붝�.������oWBժ�꽵#b���ؿT��9�>���\f����ޭ������<D0��p�:��3_a��H;��|�^I�W�b��lk��Lf<��e-X&�L��J0CI�[W�l���n��	X�;"�'D�%����OVW'����e+7���
��o.O�K>�ޅ��4�2B`G�EyDl��1�f̗��g*`�������%�4��2`��ѣez���VA��0�X|Z��/ �_��ٴ��lՊ�N_X�e
ы�a.�>��=^+;�'j�.���5�{�1 l!�)"zp襄�w�ݭ������LG��n�Y*��:�*}fQ��2Jܪ�+��˒�0��dWm�y��#��b`���E4lb�]��;ɼ�7"�h9
���ÊYw�݌�#2B��(��Д�ķ���s2Z�[� � �C����.��(o����}x�~B�Ϳw�Q�����hcE���N�Z�x�����`�;� ��}s=�2���~v}��K�Xxhzj/�t ��Y_X1WGv./D<��~�)ڀ�؃>���mi��:H|8�V��
o9C����sVK�m-0r�C+�؇w'ڲ� !�cE�m�]��~�i����<���1�2��Ջٮ��Jї�N�3bWO����7uѧ�#��b�}3���U@ӏU�1`~�{V��$>�߫�~�dy�����B�t�����"*dbk�\�B��;�J6�C�N��dd���<�������ե� ���4�R��u����b����}w=�4���ִM:F,�c��Lx�1C:0�^:�έ��h�H�^8^녈w!���AZB��V�Kr��f�y��o88��h-G����r١�,G��߶��O��Cm����0�p�J�V/F��O
H]�)�]����H+Sz����^�C��K�pB�x��u�T��5x`B���EW�0�}����G�����&��J����>�ɇ��5���	����JO5�����!Ӵ���R]�f����m\B���0�&��k�&��6;S ��}\B��QC,�����$��q&��lbYU/ׇ���2�`�{+!@1&L	��s9�J�j}jP܇���w�)8 ,��W������+AF�խF��[�@��u�RG�v�VH0��[�s�lߧ�^[�}��U�lR*�E
^��2��:�b����	�E`H�V6�FI�q�Myκ���VP��)V��;�W,89&��B=�D_#�Y�����q	�����\$`3�d�C�/�2:L	��{��NP�
9���؍�d_�����PTMw�G�T��]��@r�>M���ȨP�u�Նn�Q�cA�!S��U.��S;���eV	>Q&D��\��}8��ꛜ2b���n�[���n�0_��8��^C%@�ND��*��jX����n��2	ɱIc��jQ<��D,��[��
���Lys�5^{]vw�To�1�䊞�K��JN�<��WtW+<����J��h���r�ݵ
p-����U;�[w>�שX^?y���M���h�]�;��
]R/����x�\��nF̨�X(I�Rr�8�
=Y4g�r�bf���sٹ�tS�g�xi*�_W� �w�}�x�Uf�9��󧻙'uB���� 0xU��
r"
�)Q�C�B�
�ج��fƟ�ϖ,U*����x���|X�0g�0�������'riK�Q׆��*n�Q⺀�ںzW����r{�,�;�cGޯQP���yJ��n�~�m
���t����N�_��z�R��!���f�zӋ����i���=�sG�q��!�<� z��^hh.Td�'�r�g+9[���ٹ�ٴ�?N�P*�:5�3�)V}�^�@:��
��	�����q��,�io{fiY�9X�6�%��\%�6����[��؊���5l�=Rjy�rF]c���n��X�{ݤo.�B��tO\���G����3��Q��l,�v�JZ,Qfy}��Rm�٩]b��gqR�;�V�8=G�I_��n��zT��JƲӠs�co6QZ셽gJX�Ѡ��d"CŋjmIeḽ��Q�{�0D`���V��E,��w��}��^��{��U��S�ֆF_c�-�!{�I��z�M.�¦@!��i�^�yD��+��)��$�%���Ѝ�v��7���bkn둦��/��T�A�ko�{z+�y�LV�b�L)y�������G�C>��B���ۺn:ә��Uoz0b8�4i��5E��kV��]#Y1���-hR�N`��Ht$_2��+j^NƦ��A�km�&@����#R��u���2�/\�f�Һʫnȼ����e;I`�`fHF�ӡj'B4��M�)�ұ�sH��6�{ݽ���ݾ���q!ٍ�`+f��}�s].�bkT��o2�����q�˧����ނ�,��ѭY�F����]Em=�[cB�2�k�,�����&v1��֔����w��x���(�aE�o����\��ǜ޸$J����.#t{k$U�Hz$��ĩQc���)lh$u���u�Z������S}0�a��:�Dr�=nAHc��iޱ��#���@T�`�����]6�W/i5=t��5d�6�5B:�n��TI.IsA
�;N>��5
�+�z�	�':�x�`�+�x	gq����$ck�sa�Ϙ!��Yy٧�Uhj�LNN���M���177�db�ͬ�`=٧3�ΥBj�*bc>��S"�9{�l��W�X�:��k�S�dć�m2��YS1��gu����Z��x��OVv���/��w�3F��,��6,a��F�,ԗ�m+�V�+=���)�<z�_�ڳ�]�i^���I�Ӣ�R��A���U�ɥ�7|��1��"���WB������-e��8i]�4��<T���d���GX�В%�}��h{��Cދ�?_]w�a��ss��,6���:#�'!�:�`�V�[p�ep��Ղ����b���ֺع�B�m���a�܂P�m���n�������2�r���EM+�4��{�E@FW��vB9�{�Z�h '��%[6��kG��]��0�����B>z�Q���ƨb��Zn��h-W��4X���Gl.S��˩YĎTZ8���_]hU��mL=*�v1-��'�vf�^�ί���&�����]�z�h�5���ݓDčm
؉8삧w�7-쓤�t�|�n��'C�Ձ̧:�Zx�]�p��Q4�(�v-M��cHw|u*�K�]�ǻj�W#A9Rh����2`v��h���Y�l	ۦn��֓�&v��ð1u%I�(W(��4���sqӣa��2�ir���ڣ�	�4���MT��i=�U�0e�voJ�Ϻ��W�r;��h h�r��^�ͩ���B�B-yk�����@Hr�o3�D�7Bޱ��!Wu��G��gFR�ۈ\�Q�r��K޵���d��opZ;N�u�]�䝂쩱��Sp�ަZ�'�m�=�2Pn�{#mSI,ùL���d���^�TR�*��9N�;��ť���\ �ۑM��]���f�]k\J����N��&A���@�V�ٽ����ܘ�/���,�饦�(�wׄ���T�wJ�i}�2	���v�[��0�[S�"u��nl\f�xi<�* ����<���y��Y��8J�I�ҕJ�n	�!|���s�{3����b�c(���r 8�w�޽ ����^h���=޴�!
S��Y����Wm鱔�+4���c]�	���N��O�m=2��i�aRQ������.^RŨaO�� �V@ʽ�ɬG���J�KM�ݡHoR��&t(�1����>#�?@� KJ ��Rµ �ڱ�mVZ�����ԫ�H�hUU��Pm�҂�Tc��V�
[(�EVҨ�%cjԨ=Ҩ��"R�5*�X��VUDPR(��DF�PUTX�U`��b�J�щmm�R��T���,�Z��+��*��mlZ	l
"�,�UkDE����Ң��-(�QQUQX���ڶ֔+-iV���c[mE��[jV�X���DTm
�Z�h
֍h-lX֢���k�� ��k�+椬�]>t�8��y�W��[�Sn��QZ5�������;�Lv���/�m֢n6xt�!0�{�ǪgS�t���
�E�a�(�2	�}ɪ��]�%m���p�Ƚ�0�u$:�Xtݡ ��+���B���[��c���߉���k��u-�Ln�r6su�)V�&w�B��Պ�ʡa$��#j���{44�F��@�7+�NQ��*�&գ���:4;&v0o�QV�ޮ���P#�y�w����<ϕ]|�E7ש�{�������i�%c}��ί59S�P=
~�5��<�ǣ^N��+:�X��#���Fq�S�S}L��"�m-��l���{QAW�@u���^�1���dZ�6��qwiŌaҹգ$��0��ێs�T���� Rm��డ;��S��{^ޢ_�j`�C�D���ݏU�T �,�g
!�/<[0�٣S*��}]�Qr�Qz���z�i�������Mn�rs�׎Wf��v�c}ö��	 ��a���X�t���^��7�Fq��������F�b�1NJMr[�ޫR*{��W��GqR��z�vY�;2N>/~R�jR�b��p��M��'��Z1*�'j����^pI��F[5Bx�eT�G�Ysv��&�f:�SHH"0w�Q���R���1�W�`����{\��墙�vrͻ=��r<�ӊ���}ܕ^G���~����ei�sr�A6���1$�v���3��BEW;��\*�������Ys���E��v"��O`���`�)¦���@����Þ�&��ÞLelч��H�+���7�v�w'ShsM]�m��{(_@����a��K�Y�ߙu9,��&"�����6מ��-_�܍7~}�3}��E�k�Yy�shR�Ӽٕ��B8EM� �=3��N�n�Շl����7���FP����2w��c~#}5��qkno2�z����޽M���	��ty��=W԰�z�]��EX��ی�����L�%K�l�Į_�"���B3+����w�\�X�o؁��v�JF������8`�f������;=m��g݇c{���(�Jo�{��ε��,����uF�R9;	\(��������e�w]~?�>��u�G
��ڡ�l��7}��iX�ark�?��<��<W����Hғ�p�v��Sֺ�r�'A���(S����'[U:,�R��6Pއ�7�.;"&^��-��\�(M�C��ۿ�^5�|ξ�S̓� ��V'5E�\��|A�qQtViO`?V��&4F&��Ri㨪*v�j�)���'���b}�Z�<)H�Y�j�R��g��1#(���rL`���hN+)�Iv2^r��B���\�t:�ؼ<J1C$�lD[���&�(����%��xM���bq�jF���)���5VH�շ�~��J3����ޚ��܎�BF�R�d���4�^��,	��L9�}_d�<%^}[}����l�ej՝��7�w���3��̌Ž���^;���3�H�h����b��HܩA�Oi�liv�
�շ�S��~��d�H.�8!�$�n�D_k�8�u-����m��M���������k)��W0L�'�xfMM�������RM
���L�N��F�R��0J+n�9���`1��uN�*�C"�щ���l�t{��U����7�Hm]b�2��K�*��yJ�
k��h�� �Bq��^��_���z��T=�t�0��zV�=�Җ���D7`7b�<e��#�W�f�r	�x<>W��n�u��<�[E�y�4�9Z�J[θ�0����+���J��/E����P�:���&VC�&w��:{���>I�^��~�$����Q#MP�Z�����o��߈z�<Ia��r��M�]����}��Ǔ�C̸Ǿ���-�"x��m=��=����凥�|�K�*o���gC�X�=���ZS�;j�Q��&蜮����g��-�9��!��������87R�i�9YS�nx/f��P��.��g8�T��R��is|���*�:��Wʆq�=���e��O�'��sϤ���[��'2��	y�Q��}��2�bb����7�]����4���R����썡�u�^�u;$J
���-�;�<G�!�ܹX�$Wa�(����˚�v����%J��+��Y�7y�|��8�IU&Eq�N�cT�#J�ͻ-A�=�lK��l@'�D.�fB.�d����fe�țlRPWo�H�:xl�2���i�{�����R��,gF�^�3��[��XoY.��/6��`�xT��V�e��}�X���U�sJ�������P�˓~G��4�\7�A�;���#��:�����=����Ľ'��_Sڄ�9�:}ܪ%�>A{QjR��ݑ�B�mF�&�̭����3��P����[��U�V�4"D�bnmo_�k���d�N;4�F]�<��^9�q����*�x�z�ٷ)��ХΨ+�јL��ц�:'��%����T����Y�,_ʦw~W����[m�}S�
K�����p�WD��nh5	3����k�hsˋ}q��O���hZNZ���Zz�uW���}��C'��Y�J0����)��Y	�D�Am�|p[?�nS_}]1��)M�r8kQ!��Z�q��ޮ�0X!�{��*�����ƑZ��3Rui��wa�%P+�xv�[�]��HH'A�L'W�ī�mPW�,�R��6�bX~�z�m���]�k��&��C��y���egOt+�ֆ�����-������T3|P���*j ��7o\��xSɕ#R�'�h�5�<9>�k˯�b�}]94�NO�tJ'2�2������msT��J�y�5�
o��R���A�o���z�RnE��r�.h��D�<Un�Y��s^��׸KS���(rܦ,-�u~K� �wqM�Ha�R�����9���K,j5攰��<y7��%��^͔K�\�-{�����B�GW_/z%
G�8�����]�ɳ:�/5|p�En�yCgD�Nި����t�ۺ�77|Z�ݖR��}�Hܱ!��&�E=e�*Z�jrz���+�8����D��!�"Y"�g����7)#����΍�HT�[�y^�������Cr����o���E�"m��V$�;�u������w>|��:\s�+�D��u���1���v3J0^��۾q].nOt<����u�{f�A�s������6˩ �
�wX�S���%�w��۩�B7�҃��=k��+DD���\����N6ڪ�j�'s�Y��}��;���Ѥ1���P�>�a�N�x��-��Z�o���`��(���9Gu���O�g��'�Fƅ��p����6�TfM���nE���U_Q�)>@��y-Q�h�!NF�}�`t^��9����B@�CliSG���T6�th�2�ȉ��p�N��퓏�t�Nb�vyp�.]�2����(jv$Ò�$[�����,�7�_7�{�ab��1J��s�u[�~jôu�@u���:�!a�6���gQҹa�v��(D�Y�X<3.��7���Х��#e�]�]!�+�v-m
G��<9�Ő����^rT�-���i��J��wDv�YZ��2�]��^qZu�\5�� s�����;1�(�U�6><q���j�Y���c�~]��U�����ʵȆ�G
�65F�؝l�-X�A4/�4s5��D��z��B1jrCQ�f�$�t%��>'�}���k{)���2S�j��V�<C*޴��b�0�Q���oP������j�X{�-R�I��u>�V���[�-B�m��Z*Y��#�K��#Υȱ�9��b��蛉e�l_^�:��Q�n�2eJ���D,���{1�W|�ֺ;��lj�llcsqor>�(D+Q},l |��^�t�1'����e�p��j<_D�U�9��rP�v9���9�����,��LݷM���9����(eu4F���ˤn��%c2 ���{*5{����bv�sk���qP���.���.x�K<��W�z.����>�Qp+HދNW}��m2�p��A����v���/d�6NI�n���]���K�*<��c�ZI�� ���1��M��Gl�WsfW'٩��sZa�v��ld����ì<�2�0,u��7@k����#��F��#����+��ťmL��ྮ�m �5�Th��u��{�"0�딭����%�6�<ގIo(V�H�Z|����mF�u�_=��'�����bp0�&y��e�S�vp�2Z���ε;CYa6�f=�.Z�\��K5��8�j����W�s8m��n�J�����ӗ��H#Ԧ��ɞ�c
��	�]�yǿ9"��ƶգm�3��kR��1��eh1c���b���[m*"(��j��KkR�%k*
�E�,�*"*�V(��*U�k*�-�ĬPD�5TE-)ib���*�[B�B�[j�aEj�(%eJ�#Z�"�\�`�

���(�"(e+Z���UUQA��Z� �"%kưDL�5*�*��(�Q�%R"�IX�\1*��b�(�A`�3(�+eQ_����JdA����䶣C��X�Ғn��+0��Tst]v)Y]cp�.)W~�V����]�����l�ZT*���(L�l�ϖ��]�,;z�_j�S���.���f�چק'=����]l�K�/��A����f��ww7��R�:���f��R�v���"��l���2K���]R]I��N�	Xӈ�YI�:�'9.�Vsv�g�>��f�!��O�p�����˻�5�o�H#p���R�r�h�w��u��v1S|"΋��N�Y�!o79���'yZ�l�h�N��ݞ`؅8T�z���w�&�[c�����f�Ocn�!&��)n�S3�P�����*"SW�Y�`��
�=�M�ݶ���AG�<�Ƥ4�Jfh���Z�4ɐ��nD��C�"�������d�a�q�VI^���xE�-�7�>�g��15��Z��~%L�<d7ݳ�y=�Z,|�u¢G�BaT�ܲ���������c�4��a��e�@ם���+�Ϡ�~L�6�P����fU(ѡ���t��}���4V���V���Ǭ��T�ge�K��z�x9����Q�>�'a`푫���QY��4��y� Hܡ'c����#��}KA��ʷ�QsO����##B�A
���T�q�Y�ӏw�k�9<ty�/��h\���ɣnoX�E��n$��H��g}�;2��*��������r�c�x�><�r
y�zن*|NJ���6�y�o�/"���7⌸���p�#BN�\����o�lb�ݺ�z|�حI�}_P���n�|&f/t�yD�Sֹ�He_[��sv�j�;�C��A�p�qJ���8���֑e���!0
țh�6lڋi@x�fel	��w������Q5�-��,�tY�=���F��T�T�B3|fZu��x�#a�
�t�z���Wfu_��&����!��IJ��9;7�٥��dbm�u u�U��$��Nu*�-��#y`�o�θ��X}B�9��e	�]l�}�V���k�Q�M�<���v�������֦=�!�k]����z?��w$���Ú!���;r��,�ɝ���IGҬ䳣m���L�2,�n\��J��gx�Uk�+���{��,,Q$��m�Y����2�n*~�����ӫ��*Kt8��NF4y��Z�+����]GO��龑ݧ�n�n��������1�9��[��}�g�i���ޮPG��G��z"q�������zDg�z�88�Z�]���m��O��������4'Z���k��h�zZ�e��a��p[� �u�ۖ�;8��s���b��\Y��4B�oҺ�y;�|�NcK���*�,hߴ>�p64:gGK�N��r�i��b+(>6���)���j����{�V�ĥ�*�1�S5)�t��Z็a�jM�轙���� z��8�ۚM1���|�2�c�u��+JS-��n��9��ӚNk���L�3N��u����o��<�r��]6���ޕ/%�ƌ��q�n��g$��!��2���<g9�z��!��a��+&�����c<Oe�Ⱥ,� ҳ+@�1r��Ʒ\OnV���I�N���X�.'��Xu�E����3���e}Z;�qEW{�g��s�'��n�/(O	�PMd��Y�C��Y�u���N�6x��a���H|���~��K%�Cg�?A����d����4�̂�	��M�w�����>�@!�e�RSv��y	{%Kg.����о���G�f����e�WFI^��o�C�3����0Қ���
�:{�ws��[��C:�K�]�K}�����/���"=�����o�ŭܮ;�}ANM���W�a��!9ѽ[���Jh�����m���[<�"ڰ"Mw$�N�[()�Bn�S�۱����$�/N��杍�|����V��ִ׭����A��$f�f�LH�:��"݅ ��t^�}C�3�8ݰj�X�@מ	�d��{m�S�j�NJ��3x�ѥB�O�#y������$��X�y��s��_7���f��]��G3.�c⻡����tо4.d$�	Შv�h4"ԧ��薳ʌ������sq*�>T.dLZ�NV���n�⤬���t���Ʊ测&��mR̹���}E�G~⑕�s��[�zF1*0�Qyܜ�p��*����TC<��[�Y�*]�rO�w=�K���e� hSl;���d:�Ü�W��������}O�B��-x��#�k[�V��̃Z�N�x��@�^��!��~�
�D?BTT1m��ֹ���yv�RT�Sy��c���>��Oe�l����Rw��m3k�u&���CZ�;jH���y�/ևT �{@��5�&�pM��|��yV�~����gk����Ɩ������y�p�j�N�k���<"����:�^�aW bYX(Q�+���V9�l^�
�׃3�&ғ-vKӤ�nW3]���4�s��n��&�5؞����削9&�>��ӏ��D]���ݡtmJ�gVF�/;��ڜیt]!w�4���F�Δ�������^�CS�-��Es�MQo�iNq19-��5��}V���o,��=�D�FK�<�=ޫ2��j�ܧ��2�CT$������:�[�Ok����2�r���-��tI�ׅ�>/�{"�0�ڇ{�}�g)��}PI݃�&˱���X����H�[C�╫sL	2��.��^��t@�����iOP��\Z��y\��hp�!���T3G��_��ZB^}���_,V o���m�qJ�0�>��1u�c{��@ڙ��d7�T}�'�9���asdW>v2-w#�"�j�&��%aW��h. �c܅5%��'���F�T�t��G&���Ԡ��*�rW����b��ўR��WQ8N��1J$VZ�/��>�����!�وܑ���|[�o�N�U���֩VK}�Z�y+���^p75�o5��1y��mh�ʴ��ᔆ�{Z����3]b�ƿ,ˌ4�[�4���g	<�o�<�� �W��x&@sǮ��;Op�&p��[�
�ߍ*���	4')�ֵ�^�����r�k���V�*��y�:��]�Jħ8&������V5��I�C�]K�k������}����>�ʜ+LFI&ԏN��p`�+�`ut���"jn��̮�WwM7�S`{D��)��8�b^��:f���l�G�);oޯ��(:g��l�5�������)��ʲ:�9J���5�	/)��^�dI^����:ү|��<�����N�k{�s�gf��TEG.U���V6��Ox��w[t��s9�Zu��g<{�n�c��[��9�(u}[yܕ��"�q&Ԣ�3b��9�e����E;�l8�r��6Jr�Ch�0kLN�欺�%��%�>���U�S��hcn�!m\dSy,���W��ݏ�kfms=�E���/ZSZN�fu=���_S�����֧��3�Q���S�E:;>�"�ң�h�kj�cq&�̲p]AkU`�t��9'.���K�¬�m��}f�To�۽�����0�׷w��E[M���|�B��Ø�<��M����78�IwWj���x�ޭ����Mn�O�QgFIITU��	Zd�a�K�Aa��ɹ]�e�5{��,X��f��^���7l�y�Y	��a�=D���zF��v��7���N��f�Gxb�Ubr��ٳ�!��&<��[�,�r�@��Y���퍬�.���.�v�w��h��\�����"����_[�
ܹ9v,�fw�˵n�$mQ�7����]V�*�-��mp�x���m��A{Ԗڸ��h��n����V�z��x��f���s9G���}gAZ8YR��T�^��=ڎ��H\u��GpYVee����=W��n�n�K7l5�0��[�Z�b��[�۫��M�PX�8���n�(���3���5AȝZ��v���Ns��Ǫ�i����ӿ��
�(\�C��z�((��Rwi}ݍ�p�{�%��)�gNB�IE��h���L�<���<��A�uċCV�3Y/NL���k�Gr�Dj״�jI���En_ݭJ�����A���x;^�s�V���8�}؉y)�3B�;-�����;��c}D�Sm�����R&��x0��(��Z�=J4\j��`7;N^��˥و�rFY}�b@un��k67���wcC/�-��D�e�����J0ƻi�.^wHؗ�"/-�1��c�f�f�6�Ц�Ws&�Ӗ�*���Z���t:IL>k��u��Z� ��n��U1=1��x7pW/�H���ir��bqY��P�՗��Sle����Bh��b�*ᲧACI/�+�8�(,y��'���n�gSt%~�e
 @kA�LJ�EEm�,QY�qDUX�Il��R�����"�ʸ�a�6�qj,F�h*e�*�E`�3q��#1�J����P�����mF1�TD��ԣ�f�q*�"��lUb�Q
�-�L�����R�UBۗ2��q�e�DAQ�UB���*1kS,̱EKlb��X��V�,+cULJ�%��E�,�\1+%aF �5-�XV�J���b�T�DVڭ�,EX��.%E�5RбQ���UUU�+KE��VeTc���j�ʣl�F�EE]0�ի1����|���@  5��go�d=k�Ǒ^1�$�\$"Q��V�h�}�My�[��;�GzP�rI;�i�{Z<i��3^���).�u�E����(�N���o*�o��t3�j�-7��z�}|����Gg����R'���Ro{����WS�Nbd���J��3�����;=�w���R���Yys�(�i��E�g|�{"t)FЗ,�uR�p��5\��H�����Hw��J����������i�vR����I���ul��ߘ��w�*W��8�-k��k]D�]�`g�vB���\)��Fm،��ts���$�g(?_��4��y�|x������_�+T�V�RϘ}>�k^�ٚ�׈��|�j�D:�nH�|�.����Þ��;���T�Wh9C��d)��su�����}op�=��WPN",�H��fH���^{�T
��I�¤u!Υ�𬵢#��+�'��G(f��ݕxb��sSN»Y�<��7wV��"FR�*x�YM�//y]�\}CV�/d����_w��-L;��B0��A5�����g�&-%�X6�*4^�1�胳���B/�M㼫|�8O�������k��PGp��Q�3�Y��[�W_vu+�rU��I^NoCΨa��'�����q��{%Ɋ[��>[V9�<�+�C��B:�S2��[�X�Oi�V�d��`R�"��b�Z�-.��[�JL]o[r��I���2-GeS�Yƞ�{N9��s��)r��P,>Q7���I��I��V5u�;��ݾn{R8$����/$�'��#w��[s��.a�;C��	�p!�f3Ae�m��D�_*b�Ж�9�0m-���o��lA)����f���[�����V��Wl�T����Pv�^�tr�2:=�uA�gve�qǵ�j�.��U�$ۙ�ޠ�Dj����I��F��%�p�Fi�̴�;���PM�:���e){FulFڟ`�9�R�Ǽ������,n�H��|��C[�1�z���\sx>�.��S�h!����(ĺ�qG-4�����c�b�qU�j"ރ���יL6��p�y}N�;i2�	Ϻ�yt��,3
Vz�/`�]��սI�N3���%���A�j�Vz�J��Er��	���qx������#��9�aYa(�9����x9��:�MŲ�:����H���+�sY�܃�Ô��NB�V"j���ݨ���M�Tf�F�ɧ����-�$�E����L3:6���=��kf`Ї�p����M�q�9Ս�P	�ހC�67.A��K[T�L���^Ƿb��\�C�nx
�[��+�?uwM�h��J�>������f�-�"s��g:5�w;\��A�$n�Y���&�����!�s}����Dm�_wygjHHYw$�K�w�yDW�[t	^�|��fyY���pO�f@1�9�ؔ�]5\6?xu`m�)5;S��
/`K�N5J����s���U�8z���tH��j���M.졇�m���2�u�2k}�Ȝ��;�qӳ����4�'���ҭ��7v�9�YH�	����%:�8�.�ӗT&����v�yu3[�u��&�=�W�*T��=Op���H�s1�}go�;�ȩ�*���7��a��̩��"�����K��ljù� ��
�Ǟv�U���-����38o��s��U��%�hh���<eX�
slh�#���F�U:k�4��f�
�KP�W��#�x�t]�m'�pmt����
�.%��2��՗0���;*N�F�99��
�%�M'����yM���D���/B�u��z��C��(�<��?N�EV�7��>+�E~;�)3�탻30�<���ֻa�z�,��.��܌�����Y����y'3�r���ԥ�#\*r��K�A��a1�UW��Ϣ�=����1F��(ܧ�"�v��y�U�1Wl��G�'�9�::�D�<�-��UÉ�MZ�W�t�8Ɠ�l�e7d��'sy��a�y��wW�m��')m�J��0�����w�e��ѧ0$/�����Gh�8�Hp��O��9ν�(��;��vҡ�G8s�������rVۻfrd�H�Q���,���^:]�j��w����1@r�6��YjQ��`�u�J�'�͍z�T�iNe���6f+f��6ši�pi]�>���bqׯ�"D��K�x�އӣ����N��l���T�9�;���[[z�XΟgQ�_%vz.5�x�U\V�|]�b��R(��Az�y�j5U=��6�jp��.&�aoR�s�.��RzW'����g���LԗS;�^�lewoKk�*��n��\�O���YO�P^[W�n�U	n�$p��^ly���&+kV���Є$`͉jT����~
�>���3P�p
�
=5�;P�߼�:Q��g5���;]o�]<1NltL�c5����D��NB�벸>�o&1�`W*�EaԾ��m7+#�P�{0ql��K��D�&�j���o�!$o-ѓ��k���Ví�����̴f�fe��k�Sv(A�m�$f�C��@҄�=7�3Ԗ��H>/����H(�I��a�R�n��o#jm"Z��%�ud�=0�+����ڨ�fֳϻ��^1]7;C�ǽ��M�X�_-��Y��{ǮT���9��)�B�FOnC��T��e>N�1�����/c������Q�7h��q�隣��ꌝ��l��b'��B�H���J5��^�,��Z$I�a��j�զX:�������j*���p+�!�M�1��oL�&H�Xl�e��\m�̊�A���H�4��:Kłz��gF:���}퐘.L��t٭�-��W�*�e&om��dw�'����y�V$ŷ!+	�ŷ~�:�XnR��K�V��|�x��l�%X���ъ������K47�!�z�>&ٶ�6�Dd��r�
���h�4��Ʀ���ױ�Y(E;��KӪ�X�ԅ�f�o�Q暋�`�i�E�X+4f�^J{(���[���D �M�`�]��ל�����[��m\ �2\۲苴w��ݞ;�h]G�I��1S(�O�.�;�kW�ӻJ��A���l�����v~�mC~S�������
�m�+�g]��������yH�앐O�s��'��c�	�5 S��/� ����w��Yt�w�mF
��[�s>	��[����P�adE�\���l�{�#r���N�M߹��aw�좵y��G,�c�u�s}p�R�l�8g�p��٥_e��}��K�L�y�I�]��e ��U�D�D�Q�)��G����LMr�{��;BSsg�Z���_��oc.��8:G"2Q��p�q�i\����筋O،���#��B�dd`�Ӎ%����
G9��1E�V� ��`�M�'��{d�w'�rv�/r�8��|z�#�r���[��I�4
�{z%�-}�ܲ/q=;@��Nѵ%=��(�$�@�'s��m'���:�`N���A����s8IZv+�o�� ��T�Q����0�y�Cɷ]5��s�:ۺ�Q1P�uz�%��*��W�k�v����	4�) �m̤@u;"Wڛ#�S�E-�����P4&9M�ڝ[�h��ZU���"$s�L�AiN݌c&m3�h�4� �C)��08�=�<��aEjRV�g���X�sZC+�(�8�]��M8/2��<�
YN`o�C2I���
T�q�����f��U�"J%a�[�q�q M�'6�e))�̛��h��r
s�;��)��a��5BC	�֍�B��O�f.��1e&F�7;.(�h�r���.Bq�}.!|B�A�)�O�뇪0ElZ���2�įS�^nX�"j� )�K�g�S�is�3)�;5���b���O:[��%4�����V�s�̈́AȜ@hH"���Ǔk��ډm�[&Bz�iJ0�Jk����e��ZJ��u���+ ��&���D$��d9��,��%6�(�nJ�n=��m�G�c��n-/7�������ׁu�6w�����H�m�n&BBd�w�{�+I��TҜ̠��T6 N�j��v���s�(�}h����FWs]��[+X�[O�>���JK`g2��Ͱٛ�:&���R�Q�\�0Xw���P��*b�k^h<��2.ۭԻn� ��� �Ko�n����[*e��a����}�4e:�����5��p.R�-�]�J�����7�{
D�.�3+9�b±.	%>�g�*S4N�p%�&%�;o�t{�\���*H!sT�Jc1�d����+MgCm�ˎgUҺ
���C�>�V�40EE�m��j�4�X���UfZ���0��U\�A��YmPEQ��������*�V�d�M\J*���uJ(Ƀ++��U�qƌ1(�DVR�2ʗ�&&YL�r�Ƣ��V�B���2�֮��j�!�ʹ�pY����AL��ʕ.%1�U-���KM3SMƈ�E5��d��ڭ����jKVƕ��:q4�[e�[\Lʵ1�([kr��A�T�m���l�`���&�V�����r�P�[l2኶�[mZSHS�t�[���%�� �ɹ�#]��rp�y�ff�$M�}�G��������9%��Ee_����w�	�8L� �P�z��X-�b*�;R�F="�G�����i�+�i�S�WH������s�r��O�y�5�f)�]Sj�%Nװ�)��4' �Q��z�E$):�H�)X���	:���=�)�ŵ��tVюƉ58��[0��f���5����۴��i" �s������4�Js�rc�<��+>1m)57JV�.'�{�p�r#Th�>��:�Vq��q���gELc��Xѥ�W��RY�EXŀ�<5Q�]w@�:�xN��בo���Ϣ!����ݼx_p=���YCp^�3��Y��;���xp0JͣAeR��/1�9t��W=�2�&3kc�Xt�T�N���;�)���bw�U��P�"[�&"����R:��m{�W�5]�0<E�j�\d��xUν��9$p��S�)�*��ڱK�ɤ���b��:�[�W�HB�W&xD�-��{P��vh�Vx�e=��4�hs��ݶ���� �w�_(�ħ��z�fS�36�ưĊ3�O}��(�X�9@�]���<N�m#ʥ��g��盵�'ܧi��gFoXd��V��)�\R�T���*�=�`�����K��xoWo�����?��5Eې�}�g��I_Z���èwq�7:l2�1�:���ֺ��z�mb�s�d�f��:n�]N��� �drm?z���(&Y�0j��I�v�JK��{��{���M�aN��^�gdlș��JV$�M��[�O������^�$���Y��֘��1ώ>Q��"2dܼK��[x��B��jP�M�{i3���V�Bu�i��ίu*�E��:�6�"	5��ʻ�����tg��4��ҟj]a���t]���U��9#|���-�*V�����+v�"^��WD��w�H28D�6��5�1�M��k_� Ї>�7�F���,����գxOIa*�s�NS�l2$sj(�ݪVUJ ��BQ˼���aX4U�*�՘���]=8�s�](�#��͎B8��&F�޷Z�++{���]��-̷8QG#��ꎲ�������-�ۗ~�o*=^|�ޘ}�m��N�&��>+;���)���u�a�/VQ�v�����˖Q1���ݛ̮�a�`�Qk-��2�)�Uל�"UN�z�* ��B����S����=�"o���+a�׉ S�����*�]v�~so�]�F��y{����MɡۯM��p�#r���(�{�}o���b|�e�2�aOd^�͗����,�.�9!��������i���Aʴ˺ܤ�oP+|K��P�dy^���G�3��0�t ��#��M+��ΏD c���D�V�Yò�v�Eŀ{��N���bN�β�9��gypiZ t�FC7/��B����7�B���뚂��,�';JS�g͓'b*7Fх�*w)�)LO^1̊���jB�eE���=Pל��ٕT�A1�/�0j�� ��lQ�o5�nn�6hd!��F���׵؟'y<��Qb��k�>�q�&u��ۮ3�ImV!������n�_�Α<#�L���^i5��O#PY/�Gf#/���o9J-������]~yd��3֜:�}B��Q"��>�s�zLֈ��k���:���Qrby��>E�}�u���*c�3�[�m/\{�U���ė9��-\�%,T��xGV�2��٩=��<3]q~Gs����c;�l�ց��hެ,'d[���j�g����4�ɬ��슜��k;�ݵ����>ŲHɤ��s=�[F�]c:s���x�)һ۲������`�f}O�_\�(@6ɸx{n��Ώ֝9��{�&��d��r���>�X��2&�����6Vm��2{�,���F�]�R:����>��
1$Q.���FH�G��L�<:"(T�5Ħ�u'��h�#*���>�!�����im`alJ�'�M�m���"���$Q�;�P�����_�5�[��m����4�N�w�w�g�]�Ǐ3�/���f�V褮�P��<�+i�u��(k쾲�(��OIٳE�od7�uiF̆Ø�vqE;:�j�3`p���լ�rb�����~�١W����4~�c�F��y#�oqo� �ߺ(	&%����RF�I��0+�i���bj㬛��׭��U@�7=��V͙;{���`1�E��7�o�=��ʶ�\OML���n&^��f&�hK%ȭ5s!�؟Q�g/3��3}#���K)N�F�q�[S�C�5Qj�%>�Gc�˴mr��P,�+�:���s�1��^��47����U��ý�X�Ɋ���̻���H�L��F�ts�i\�Ue��{9���4�=#U�4�o��z;P5k�2�m#��v*X�|�f�cy`ĮBoN��9�'`������JjI��%`�ڬ���9%���1�@NI���Ѩ����zy�{�Ь�索bS�ip�{ةq0K�MqM(��3�N(r���]3J��o��hj�V(��^eM�{�!b�ޝ*�������ֳ�WȦ�ɓ��m	�k;��fy�0S�2�D��bk(<�I�-�#����فq����U(*��)����9�d��e���;5��./6��3��	U龳Ka4��k+ݓ�=�X�4��hQ�y��t=�m���f�-����Ё���w���h�s��F�N��%b=�Ā�NY�b�\�n����{��\D#Y�G[i�+��k�f]2��d�ғP{D9�pC�lN�V31�r�P�+~������ͱ�8�{��.�푪}���#r��}?9]���9�i�vQΗ�ڙ�z�fϝ�b���"�W�5�����V�IU��m�y��7���= V˕ҋY��w�y������-9$��4$�EB�l)��'���8�o+M)�݃�pC(j�t��i��H����[�Ď1<#�[�U��f���f��)s�X�j���H�1E�&tC�|$^�d�
�kcTM]��hR8F�<Z�\+�������aN���[�V1Α�rcD��������W鸉�yu�8Oe���Sቧ�6�А����&<0�ϖ��"s٬V�Әî�'ņ�ª`�5�U�#����p�*1'Qm�Rȉ�ha�� �#����7�9u,��˺穂��FOF�V�]k�mI�|��t�E͔1���g��h�=�lAk*�$������Xi�6�a�����Oi�'��Ӛ�ίq^d���=-D�eݙ�ŧ�Z,k�
�����Ȣ�+<�0�<{�xYO��}G�F34�����r�f�'S�*r_��Gn��7B"D6Mt�iٯq[�Iw�g�'�τ�L;_p��%��/�D���*��i�g6�Ox~�O�\����dmv$-W�v����ɂ��R�VJżnUORv��|GRut�����:��a���.�'!`���髄�wQ���d��>�j�2�8r�������y�7��"~� �̧���Eb�F��2���R�y���*󘖍#�5n�}�bO��iff�ռC��+,-����U�l�cI5��.�&�s]�H�WpV�ʴ����]��WK�2�����V��{K
8��Q�$	�)��7M�U��R8�.����WV_s�e%�����Գ>�9�/��&0o6�˖�����U�)l)4q��\x�kF�3y8T��j!yt��MtU�j�Dk��9�,Sٛ���d��i���ij������V�^(`�j����dm���Mu�V^n�u��8�<����5N �n��j�Ú�,Jr:x�9�9�:�8nnZ�@�{F�	(�<������+��3^m
*B,�d�����Ү_+�cq �2�9髅'�v֓[����8���HY���Edߖ�]���;����Սr7�G9[�
�b#��́}v��Oow���we�g�ޖt魕sc{k	iK�{���o��k�fR��L(���jJ܉��{��gV*�J�q�q�B\�Y��\��<�;%�nVh�����o'u�Q�}y�o�=�KN)��w���B4o!ƎD"�s�� }���{�.���1Oi=���k�e����\��a�𤆾�"�B�7�4�����k���Z�a���oAS��9��ymg6�;B[|�5�@6^a����̫�"� Ӵ{�5�������Q�mحU�M^�f��G:���]���U��]嫃�.N�6Vd\W�@QBu�W4�drJ�ͫ�j����R�H�\ޒJ��V�'���^2�7�V���_�s���e�bf\��T-[Z���1�X�V�x��(���QVa[�1�UV"�5��FƕZ��p-b��2��[Ae�a\��GT��!KbQ��33I�S@��p�6�*F%�@@�V�(���b6�fV[D��m��Kp]f�ikkUL��*�r��[��jҭm�LF�(னMe���e"Ii��`��)$!�˖�X����Ɖm4�Z��(��E.arܡ\X�FW���I�id"�a�`$��(��QMe1SJ�-��--S�0b(�a��ft�-��.Z�m�%m*�1�Ƶ[���29a[jbZ%�j$�Ԧ]5�T��j�㌮Eff�T�M!��(��Km��˭iV��F�X6�=��u��W�|ᶲr#9�Sh�FWv6cݍu�eᦍ�-7�	�msr��I�����-��k�%�L���;�E�yZ�n�d��J�h��I=�T�f.<��a�	D�0�p�e�GC�!M�����+\�=R�:	��r~E;j	�Ŭ���\�Z����r�V������v���#)��*h��W��2��	6�^�7s)�Mk�9�xO���b��Ɠt)#��xܨ|;=�F��7L��e����̥�5���c�@���(�������� `����z�t����z�u��̆_et�4�R�x�k�㺃��*TX*ӓO�Ej1P�5��n����#.������H��IX�n��)t���ݹ�Y���h�Ǘ�<c̍�%o�,drYI��*�\p{�*�hg����G���<�;x� ܴ)��:�^�<F� �s��~3�V��"�ϟe��3:7b.җS�]�)�&���R�GZu�^��]����).Ҟv�=P���asj�T��"A���.)'��z��Cp�����h��A化E�cP4��z �T�;�'7����X
\`Ѕ�,oN��J����x�%�;N�Noh*yR󬮔�=,|����|y=���nډ���n9�"��ǫt$K�S���b] \]׶9W�k[�a��.��s��M�X���u�C�*�fX���8���gr��	�h�z�ެ�6zW0��l��@��B��|渰d�7������v<�����q�
2q�"�
C�RLC�ؙc��^w�U��Fb�$�u��ͲI"�V�?u*2�N�R�����:HB}�{���X����kz�6)q{��WwP�x{z�a�˓�ӳ�Ǡ�w�cZ�IĒ�SGh������2�
E.��R�8�[P�cB�%}����&�P$gY07z//w���;��DW��=[a����%y��{��&�%�W�� }I�����,�4o^�cgx�?Qe����ے#�pw2,D���wqE����������oέ��hOj��=�y�&,��X�51��&ǲ��9ތ>5���_&:^B�	�Z�z؜�-��qx~jJ[�L����{�*ZᲘ�3�^�S�vk��۹�É��C��۳��!#9Rɓ��V��OҧLVRm��C���C�˷��ՙ-·z�U6�ʭǤGwv��$���=Q��DU��b9�Wuv�� ˤ�홽J����p]D0�ب�n�~��)�Tg���݇�r�KEy�A�R��+�ޅ:{�ngy�^���Sh��^���]��Q����D��e�-�ʡ۔{-H�ٞ�S1��/�I�e=��Z:���vO?r����|3%�eFK���A�'6mk5�e&C����`�ns9X�M���g�ݒ�����52��S;��8�mwS�����{�o�M�x��28�w�3�[��;>3t������6���Gk�415�����:��آ�wYf��b�y�f�R�'�����3U�ZW	���F��4���mߐ�X��nuesD�Pn:�u~vՌN�ծ���+�Ûi��C"N�(�%@��I=�2���z�D��������l7K]�T�2�ݝp�΁��h��MuE�h�u�Is�+1����t9-Q�j�գ��h����$&�I�稵��p�[�}k�,��m�3ݪ�	��ͼ&Sپ
ޙdo���ůF�O�u��z�	�c'7�c�{�EdY'!QeuT�Ndg��F���N��$�7�X'c�	j�����Z���f8��{_�Bc�O��&���A�,�W�U��ձ�V�k�)ͥ]+��m"��Q��������N6�o^��ķ��z�����z�Ü�s9rj�Y2i>iI�c\�$�����r��pژ�5V�#9keS��~hq��}��s��Z���)��[bY[�<�(�`=�G��/	֞����J;oR��O�F�Gt+���EQx���w�]�-��b�":Λ�-�1=x��,�� @2��l9{�t�(P|�>����j���Z\6��������f���i]y�;��c�r�)�Ey��	��i&75lI�y�\�̳r�!��Y�d���pU��9�O9B��W�_+�FF����6��������0B��6�/sv���%�>3��s���EBG%�)��3��w��V�?��[5������h��@�"�Y���$�'���5���0u�9N�]��v�}�S��..S�<�7zplM���Ya,W�+�$lm�օ;|��oQ�0�0�2�L=,�k�:]����Z�lT�*��7<�N��3��Oj[{I�j^�Wt�e�T�l.s�8��*Ɨ.Dp�vȣ�T3������=��3v�	g��6�U�g�0؂u�F;M
*W�c+�g�M�������Ȗ�n7;���B��XZ�<3C��խ�2�3��+ǊФ�"�f��C A	�{��r��#�q���N����믟��:����z�4M�{w{I͏��釤<d|��;S!�����=�̝^ܟ^�Yjz�[rGu#�n%����^沩?V�FH�h◌�t��1<)�i�W�j��V9�5���d9��9����u�"r�KXy��k��&�*F���m�xT��[�9{�=��t��z4v�m[�V��XJ�e�wm2b��>���Юٔn�ڍJ�����=�l<�[\����P�6��;�6^od\�c����MJ��EWI�2�g֦������o2,O��RSn���s�e�(#Fv�`F�t@���h|��������v����3$rB���7��\���[�p��
�Kv:k���K��u�ۃX�n^�*�GE�U��[���a��1*�_Tby|��mLe�p�ܗh��e�:�$\�j��>��NC/�8@́r+E'ulv>���:a�I�>���U|.��E�*a4�g*[t�Ѩ���t^Mgsj�1yP�
R�P�kةX�&{_#N����ҹ�/hL�����Z��m���Ɏ�'֞cbݡ9 ��r����\6j��{�������`�d@lߩ*#*�Q�;�d����w�"TJݧ��3��Щ\�-��m���-�Q���2����os)y.�������ƜV�|5�\��j^S�b��������|��3��J4h����&xD�6�v+�7�y���r�;j�l.�C���3��'�%�=U�i�|đW%�4����Y��L���Ywl[OU�64�=���/�{�w-���.�.��ż4�T�̱�^�����K%,=(0���u.��ɷ�*�y�'�¥<�7���Ó]��b�{$�vQ��zW��ٱ�D��e��c(�k%�iĖÌ�e�5�W�;!X�k��v�pܩ{�d�S]ǹ��su�����˜VϿ���x���T��h"�$�I��  �1���d @����y  �?�/!���~:�����k�;�mI�s�  G�9B�� ~���;ݒh4K��>t?�@ $��`�7vO_��^q�q����>�ν�?�Øq�ӡ�ꀆ��$��{;�s��s�א�A#��ߧ�:5ׁ @��=���Ϗ���!C�h �?�2x $���XE���o�����C����O�&	�^�?��������}�>��@ $����X�������� `�����N?���Iďr����}`[�g2!���'��o�"��h��8��?��@ $�>0���W����u�Ā H��d!�:U��S����s?�:��������$ @������~�|��|�|O�$�~?B,�2|~�>[�����'�}��}������I��'��� @��;��>S��?����������l�
�~߳����}S����h}��7����9�~������}�  |������ȡ��a����x?�	�y��H@	�� 	�?|����~���B��������~������� ~㟛$ s9>X�1��(|���>g�I $2qd��@>��NC�5����+R��^d9��'<��0al?wF�5݇�����  H��~���T� H�q�H�!��>p>������^���?���a��4>�0��w�7����g��`}[�����a�B��C?���;���̀ HQ���y��	�T?D� H\���q��ч��23ϟg����'��6��8�r�G�s�"L~��~����hy���?G����:�3��q�q  �}M}p�}D��_<;OéS��>D?��C�����>��Ԓ�� �� @@�h�~���a��P�#�|�_����������a>q�!��_�I�q��NĜu�}�\�E$�PO�(��y��rE8P�;��-