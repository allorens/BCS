BZh91AY&SY�T�r�_�Pyg����߰����  `�        ��  tUV� t     
       �T(B�g�`o�7S >���UX0|%��������]��.a��6�9�N2���܏��u��}�r��|y��u�����7�o��eA�ܕ+�}h퉙b�k�>ƅS�� U[�q�C-�A6���W��λﾕ<��YO��l���N�<ś�����G�;޽ǽ�.�:�wm��ݺ���k�t^=ov�z�{��{�A�m  �@� �49�ٻ7b��o�y�Sl�^㋼en;'qG��ܑ��an���^���Z�z�^l���m�����窢�HX�*�/im��������^���O�_{��M������ zu�K֦:�.�lٹ��Z�z���m�f�75mx� Ac��z�5i����ή����ɏ[��Ǹƽ�^p
��F���ٷ�.�u�6Ξ�0=�n���6����T$�E*(            �O�4?R�TF��1=F� M �1���DIJ�44ɣCM� @%6�@�T�"i��b��� #�I��2�P� �ɦ�b2M`�M ��&�	��jhjmM12��=OT���1�M'�zz�� �3�U0�&�@h� 	�F u]���-{�-j�\�Z�e
$L�}���4�� ���PA���u � ���� A��
������}���ng���$���J��1j�m�RIA*II��$UPa����8@1jH���w	��W���~ş�M�ɸtԲs�I�:Y�'~��o��v�rΧ��8�D�������N'<C�^���Y�*�MB�M'4��=ĝ=e{���'�O'�#�ǹd�5���6�V�'��N}�Bw�%���tI�J:$��a/������	�c��w��E�"n�N|�N�VJ���n�o�iod̓�$;�'~���K5Ϭ��2s������l�4��F�hIG(C� �6�CIF�KJ.��Q^�bz�=z'�a�Q�S���ɲ�p���-%'MpM	�}H�A���9�u�����o�"Q�H�C�����&���&����%��)�NtO&��NK;�(N���쏤Mx�� ���K4i�>K�=��Ӄ�	~I�;(�͒��$:"w�"'^��>vO��9����"x�I��vO��B&ɮ�ĴD�xI:M�ZI�ZQ���H��
�%p�"6YC�O����H��'�i/�<p��'t��;hI�<'��vO��%�+I+�)I�E}Z�6���(~���$N�xJ��n��Ҏ|����<�P���	�"'~�eǄ�����=�;��M��A:��I�f��'S������B膓z�"u������p�A(�?{D��|!h���<�<(�{'�%��N"��	���>�	_P�#��N2��\�9�ӽ��tQ��rj����o�7�����<�ZzJ�'g*tޢ;��O3E3�x�p�#q/C��G�:Zx�������Y�w��b5�J6x�]O�S�n��m9ө��>����h�6W`�E}��s����yU��^؝l���s��(��ǕQ˅��C���{8o�합�]��0��{�L}Q��N�Ӆr#�TG�����$��R�">�J�# �;��gx��I�y/�O�rNhw���<͚5��CȈ�8&� ��k�K��Q�]��45DMy�D>Du��� �j'��SAUDFOv�#֥�Y�p֢%������L��%��t�!c�uQo*P��DNm�dA��5�%�#��8T�UDG��G��x��KO�hNg
�"u�K/S�&�:�D���6�(NF��?j".�P���ߪ"'�,����j�o�M�#�TN��R�<�".�'��B<�DM�e�4Ϡ�j"h{��4�"z��� �	���v�'�Բ|���O�cȍ�q�N�e�Mo�tGܨ�by�N����o�lԉiB&�4k���jQe�%TM�:�ODzM�7���	�����${���W�֪t��Q��Q67��#���D����::���z�5�C���7U6�J'�>��z���2T���!Ĥ�)�h��}_$�?n|��� �#��l��7'��}ꍥ"!�Ε��݈�<J9�zN��N�9&�#�j|�}ߺ|��Z�U��Ӑ��^#W�s�9�s����'Nl���NE�l��b�+>��_/�f}�Y�d�-8/��"�f�r��=�G���'�<nN����ؚ��;��yQyR���^��+��؆��z9�k>�����w�y�5��fz���Ⱥ��y�=�W�o\�S�*%m7iI�;iOO16'}·��jX��I���}��9����y�꘷�C�����x��ӏI	}}O������NIrk���=��~�֪v��3�>e���]3W�9�6>�'��r1��[6��>�W�l���>a���=>����}����t.����w#/����}�j/Y���ul4��ӯ���|��)���u��}[*����>}��|yoMc H��f+,��h�u$8u��C�|����l~�S���eV��)�N;��ǒ����ӧhDi��C�pG۪D�6{��~�u8�RtK<�8'��e�q�>��6%�"'��4w�YC��DN;���r�hu��DM��8��V�>�E?D�n�"y�+�J��Cȉ��DѽJn"P�"p�8P���;I�U�6�7q�%��e�D�"#�t~D�Dn"S�D�jR'����ץ|�ڕ��%7+bqܤEܮ\����D�Y\4X��唝7�W���D��"h})4y�%��+���"i�"_u)�ex��ҾM���4;��DDy8P��Bb%e�Y��G�ĿD�l��e���BT6;��O��%m�C�*x�U]d���h��{6<�7�|�g�qN2h�d:'���'NH�\(��Y��g^��Ύ�-_U}��=�'��{4�|#r�)�Y��Iì�W:'G�w��=9D�q9���,��ӒX�ؖ�m�W�m�MI<'���u)=Sl�"j�5:p�����a<�'�TO2%οDn��O�����!�d5��Ono܋�O�_M�j��'�	6W�5uMr���5ꦙ_Q�w�$!�CP~n�x��[_xz��+r����C�C�ETUl�j��B�ӥ��� �r��'�����ᾇB�P����ݏ��\��R5.jSȔu���W�7X7A>}O��E�M>_B��>���g�k�p���q�U5G]��	�?STW����mC��>����"��;ΪN��}�{-1��?���	�>�����9a1]۬Ua7)a$�*�W��S��go�g�|�!ۓ*�� 2�0c�t�̃/���=ٽ]Y�&3���W��t���۽b|��t��'���iog�(�o=��z�œ�(��x�� u��ԝ}ɻ9��O�=�ǻ�<�;4�3�G���پɅ-׾�h���Lє��g�guv�وV��f���y��}]4���y��N���nbӧs�"^^�Y�����g~�ϲw�5D�X���d̙�靃� JA����wv�%N��{���<������^�A�w��U{0`כBv�we��΄Z��gN�kDUYCl=�oc���]��e(yAoM�T�<p�Wz�e�� �O��ש�w���3g���������eU˽�>��.�>� kؼU���۰�B{��'�q�']4�z<ɬ�qfN�>�v���>�X�������M��i�^�>�;��ӓ㣞���۾k���=��`Q�ڽ��y59��;��`˄��Y}ܰ���N2��~񁱍��M~�Ft�]�v�t�O.\�!��7����f=1��nߤ:w��~�=��W������d��)��G������ ��!�����vj��;��{�~�����g�zt"�a��2ogۙ����N�z�;sK��`}���l43���$�NL!. ȝ�Iaa,���5k��@�P8ڒ�S~������sm���(�X�Y^#s�0��r��0~�z��3�{�7rn���U.�w��t]CƇ�n���7��<y|�`��Λ37��0���G�(��:M ��{�gvd�9vi�A^��`3G���TYg0#I������w���揽���]�-P��%�{ǧfE�`?�;�왕6��K�fߞ[ɯgA}�"��ch����}U��jՙ��:,yr<S;��f�����5[���H��I.�|��).,�l��J\�d�eBe��v{lO%���<{/��5E��޸�b��{p���9�m�E�ܢ�EON�׾n]']��-|��2\�1^����>�L�����ֺ�l�������{�FnNf�1w]zk�졙)J,���ah��L��M��+>1o	"�˕a�xḦ����]��~�{e"��O���kz>��K5���{>n�no���wٸ�Ͳ��3�Y~�.9�KY��~�WC��㎷8���]�ut�!<��.��4B}��&��1��^)�x�g�]3�.���z>ʪ���EN�Wq�'�w��=V/w���^����&̡���2�_e�����߮f��rM�/�17�CkO��w�13+O�߯{L?��=��˸g%K'N�wgwgs�}�ݳ�ޟO��~_��o�,ݜ˪/�(���R=o��oO�q���=�'r՘�:3����_�}�q:�$�����~~�ݧ�L�s~�X��LD�d�M��7=����FY�U���u�ɩk3ݹ��o�/��`�&��y�w%��$�Dhn�ېu���{$�qݙ������ڽ�;6kϟ���5߶��o��.���䜛�N��)�Ձ~ɝ�ےg������o��L]�$�$�~�������>�l�t~��(b�3:5,�%�=����w���o�Ϋ�o~gG͓{�3$Wg~Ҫ�1wrng��L�����~�ũ����L���j+��y�.{��n{�ʨq�;s Y�����@g)�Ӄi�����gۘ>�ܳ'*�Ff����O��Z�ɞ��F����k<�}'�!��h��(ưY���,��c��<;ro�7��wS�ٓ�9�ou��[�D��w~Ǻ�ڏ����J2�V0�~�`�sﻘ� Ou<˻3��&��vP����rcY����t~���JN����r��'��N�H��s�!�T�9ww�O^���m��K�{ow�srv���nI�3pywM��-��y}����d�U�?Og;��Gd��y�2�����M��
�������'� t��<��
A�g^M��<L�$ٿ����p�&�C�݌��3������֙e�d����g�G��u�CaXڭ��=�џ���҅�0;s>��v&�)����5<i��m� 7Z���rbF������v>g��Cw.�4���%ye���,ɳP���w�~����Oϻ�r=;���Ʌc>�>:t��q���%���׶ɴ�##�-�X���l �y��͛4�d�c�6g��e��L�lg�,���.E}��e����A�3���!�Tڅ(�ul+Á�d2�2;�m����7p 	�d��rn��ܚ}t)��td���N���u�\���UL-�$��=�%{	�J<O7G��iӶ�����n~�{���{�X/{���-��������6�}�{sF;'{������p�1�k�y�S�7i2�s��6�w�fvo�5�Od��?a;�7�ɒ;�����]��l�f��ooN��T-�k�Ξ���<�~�/���
j�l�[mʞ����gٳ��s~칝���fx7��5?��F?l��?L_	��g}�B�(����?dT^�97r{rl��6��p;ud��e�d�N��k]3Zu�q�����l�g{&v'��3Ɯf�k77nt��6n�6L�9�O�w��Ϸ=�q�,�}3�7�$nGf�jߘf�$��V�������ϟ��>ɋÝ�5�����Q�svI�cύ0�܊޼�K��Z��v�N�<�L�֚��������M����c��dsM�v,n����-ӿ�<kv�$'�)�0K�rgn���Ucy'�~�g��cY��Oޝ0?�,߻p���{3=�]�f(F;7f��2����п�/��Y��|�1��Mć�䘡ɵ�o��In í?�J�O��o��Ȱ�XXYmec�oa)e�LCM�/��M�#Ve���Ԋ�k-��k�*�+V�����uv�Uٺ�mDݨ�;u�cc��@M�ӱ�I-v�˷f�nkZ���l�jK@������>{�22Y*8�+t��0O���Jݶ�
ՒE$#
좭��)"g)'Ti�$dc�㲻*9G��)jeR��PЫMڜ�r����찖ح��aJIU�DR6ݖ�C���j��q�,�V~����)�7Hn���FT�kf���ai���$��s�ňLqd�%�j��G�#l��p�[mB+�_���/�a��J=�K�,z�I$�U�]m��j�h�3�@�Wlj�#LUBZ�T:�'-m�+�X�$�#M�/��E���ihF� �Ab�6J�	9$�~0�٨"�&<�R�O����0TjlR��Y����*���������[Kܫv[�J2���H�l�VeݻeҪ1 ܻK���8�C�L��+v����噏��@�܊9��K#좘��!1 +{*�G���Q�&��u1�"TKƫc�m�m[JQd�N����9�lTj+H���cO�Z	>Bdt�Xף���4����e�I��+�[ee,D�,��e�[̂�p��&,yV���̧8e_J��T��:�6���X
G�R�i$�6�6~��fI8T����땣�5�TF�X�U�PY�RW,��8ډVYҘ��k�U,����?\��yI���ڶ�.�� ��DͶ���vR��U�hcD��j����ڊơ�%��؝Vj��@�F�����Y�=k%*�X��OGV6�w14
i`��-�gEKS�X��r#ϛ7��m�]��)-cJ�~s���u��'T�6��jRa3!0PU8ȝpuݼ��W�v��㎕�F�x�mX�!����`"%o"�h�T�V�v[��-n�/VpUfKIc@E"pQ�����jo��(ȥj��T���]dNw���F����0�PW=4д��k��h�{�dq�������~oq�??_7d�uDj%Ej�
 ��߱�_����S��UW��UW�J��]*��t����]*�]����U�iUm��Ҫ�WJ��iU^���WJ�U^"��V���J��ZUU|�UW�UU|�V*���W�K�}	�>����,#B�H��&,C��U�	j�	eC��G�CZU�Ҫ�UUUUU_1U^+�Ux��U�UW��UmWj�j�U[Uڴ���*��iUmWjҪ���T�������U|�����������}DU�*Ȝ�$-�,�"	  F
�J���d
��'������>�ꗊ�b����Uz�*�رU|�UUU_1UUQUU�Uz����������Ҵ��R�U�WJ�U^"�T�U|�*��]*�t��V�U괫�s\�B[jR^bI�����B�*21vZ�������;UmUګj��[Uv�ڮ�W�U|�Jگ��Uz�������UWȪ�եWj��UUX���v�uT�Uګj�j�UW��U^+�Ux��]���>'�Q_|HI�����P[�%��l�Z+Q�H�P�YL�!?X�[h&,LT��b �/DL�7��Z��横B!	�����w���oSS��x�g�?AӇ�?Aå?d�-��tD��tO��:pK �"lDDO	�"AB'��BtDD�bm�b4&� ���<'JD�"lDN	�<"%�,K�؛4&��	�2| ��>A,Je�bQ�Q����8A�DO	 ���'�DN��͉� � �$4&�	���E���"K��2o�j�V��+"*$+���c}��pI8�B:�R�+q2��R��ƒn���Awu7Ym�[K�m�b�U�s�p��
�X�(����.�9l-ԪI�ܲ�i(i\�T���m���K%;i��t�i���c���v�P9\���:�hn���5�:0(�䕑�Ԓ8X��p�W�-���[*;,M4+�����ۤ�TW���[����1�G+��+U�UȜ+�r&�f���Sn�&��:ݱ���-N�e2�.�Y��j�RZ��Y����a��G�k"*���P�v��'-�UBQ�B�c�Q��
�B�N:�����b����H���,�;j�-n�D0B�[J
�娼�#UE\%��ta�n���ͅ�B�in�֩%i�]���	�"	�J��I� ��Y)j#9Djke���d�`�
�Q"Wj�v�݂R���͊�z�Ӆ-�a�̈́�I.��z�Z�o{%l����v��{�U[���Ͼ��0�����V���s����3333U[������������wwv������ŝ8t�Ӈ0�xN����8h���nf�R�M:��,X (�����mF��V,8"�∴���#�V�V��cFd+�_.	\����Z�⪭9̹T/� Q��SCE"ڝt�'8��T�
(b�uuB������f�
�4c
J�2�Bʆ��S�L���J8�g*�&�_�X�_�i+v�*��zI1.N�����������q>��#%�[�췄�����I��e����ӭ-_,��g�Y��v`��(�%ߡ��u�Yq֟8ۍ8ٶ��_��g6���?"bA��p�t���IM4Ԧ�sf�ZL�j%�#��sL�#e��!�D�Q^�iÇ�!J|nB��N�Ed>VV�eqZ��s>,��ʤ����Cf��E�}�d���s�c;�.���`�d���c�4�l�ۛ���Ӎ�mZeg�9UU,�R��,���P�;�XE0e�5Uӳ3&%�!�N/�QjxϢ��2@�DUHXk\�,�8e;����>�17�Q1���0O��;2]��N�S���V�tYW��>�Vv�̒n5=�O=L���m��M�ۍ�Ӎ�^B����� |��OF�l�-D��
�ڎ�b����$�r>��Dd�,�&d|V�4���iZJa�}�j�������.X`���fanZ���X���n�WL��y��;&z>�Ӈ����2�IsӼ�8zs7�3ĔiP[�4�*�T�=X�6p����[m��mƜl�j�/�[��b�)-)h�m�&,ذ9��q8��$a#����Mk*C�0�5�|Պ��$wbhDEh�<UF�⥲�����64��$!���#�hEr�$�� W����%��R1��w&�H4���-�;I���}��p�&\q�I4J|'�)�9�O�ĩ(�3ҳʦ��-�Dgň˵�*�9�٣�E7�ɒ��,��s'h��zC|cwZ�f�5��#$Q�3z:�YbLGw�cOV8�����[e��q�q�6ڴ���YŸ@S�%�3�U��D�ga�fL���
b��T.#�je��a��Y�ꊺ����3,쐢����(%m]��"f���̳zVR���1t�їAσ�0�C�ʆ%�g��YUY��3�76r6s˖�4�E�5T��c��gFf{e��4�-��n6�N6m�i�ʥ�U9��4�M96d��A�0d9
4t���ɖh>N��3���$k���h��B�L��]>mn3G$f嚇1��E.`�EA��ʮ+ivfY���G&%�>2c�FF�ɖ�m㎲�n��n4��yy�TO�o�tes� N�[�	M<9,NB������z[���$�me��w(j:ҍ�ZpT��GM�L��.�s�����fbd0&q���l�gN$ޞU1��Za�S���g1�jWVg��ft���m��e�m��iǒ��V��T�C=��홠<��N�������걎��j��)M#��1V�"q:� ��Ivً�l��jѲ�6�C��5Y�۠Uki�^�UՂ(�  �)��G+�N��rNRUZU�`��#ph����,�ѝ�)��G'Lh
����ҸUfg'!�n�SW�L�%�Y�m�dy7O��:3�z�mK[���K��7�)��gդ8�k����(Ͳܛ��
�ˁ��18r�8�3���D�jA����x��[m��mƜl���gE/����ʖ�YakJ�  !N.�Z����c���H�`(�t7�T��!a�Wػ�ɸ�@��5�>�6^�H�1�tf�4~7B�9�t}�Ço]�2�����FY�P���u���W�����"!�'��fwIJ�V�ɂ�V�tlL����M	�e�>~U�|Ë��
����n��:�^�ë���^:�1���WC�����>+����z=2VƇ��tK:WG��]���kJ:t�	ћ^������(�`L&RD³�V�a0L5�X��Ҏ�����GG����~;O
:t�9K��^��:f��J���Fգ�M�uiN��(L�#:(�(����Q�:!���gM:%�ΔtQ2%�(��?)�e�Һ=�;k���~:V˧�]�+�i���=giz}K��Ҏ���Ҵ3#kғ�`���d�b3�S���z��	�(z'LRΘ*`�Z��S�M��s�>�����O�w)x�)Dx��>��[�����>�.z`��<j�q�Μ��Gl��U^(�:���r�����c���H�s|���O�TUw��neW�}�S331�QU����}��3/331�1]�{����fL��w�����{�|��9�Ğ2��Yu�]u�xN��������	�UT���(4D�7���t��(dbp��p�Ș���� �!��,��k"�������_LH�Y4'Pâv0����]�[/�1��^8H�46ֵq�m�5p�L<���L�(��C�.�}���:�Q�c �R\dD�PJ�U���jU;�A��' ���H)�UU�0́BA���D(s�R�z�׭�m�4�M�ۇ\q[~i���^��UU1��~ ^�R���r|2zm����MDF�ѓ�2x̨M�g���))���ej�\��B�3�&f��<�����wK��q�� ����R�/i�����%���Q�c%�.�"%=<Q��4$�G�UQ���mbT���`����&��#1�pI/�U_��0��c+E�&"P	�!���nX�+�T�,v��G��ڬC�n$�d�b}.8��Ͳ뎶�n��$<h�F�kU�2�e5�*�!#���i �Y$���>NX�I]b���l��j�XmWU׮@��T&:#�tXL�EE|6�iQ��(�ݹI�Nۼ�o!��!]�*oC=UUQ�╶�r�li���^�%Z9�>�M�Gx�e�4bnlR��%!L_�1|\�Hg�U�/TH!%��dF	�:X�wUe��Xƣ1�U�*z����	�z�c4�(�"�.CB��dCQ�q5J��ac �@9���v�v��b��e@�'���n��b(�y��^E������FA�<M�ۥf�0�L�9��$�Y[S��Q��W6X�u�*�C_k����fΈ�<'���D�f�9!n	wUUTpĤ�b�"7)�6%��j8u� T8!Xj�BT#�L�U ���ɔ,f)��a�M)�"ڬ ��I���6�v!��X�:�<qX�*�d갲3SKߑ�o�=,��T�?�.e�1��1�7y�u��S�S2``z0:0�x�I�(�,����� �ʨT<����DC�0��	��PC���n���6]b䂤̕9��b��l�u�.���:'��	G�6s��o&�h�W+I�I"�B�7o�n'�UUQ	�4�F�=���*��'�YE�JEу�.f�) .�=Q�щy	9�~���@p� �ʙQ����RԌ)ߙ[s�Km�,,k#-�=98㋔ɟbl`z��8!�� �(��v(���3ՠ�aP�V����6�(f*Ib��y2@�;S���֫ʜ
iF��/S�M׉���N�ڍL�K,NgoT����4P���Q#أR��_����8�u���qƜlp�Ҏ,��a�"�1b5L*��(QM
����
�((�0ZQ�z�UUUUQA.!�M�gnL¡�XwlZ�H~HH0���z!'�h��T��90p��_Y�]�Cw#wIv������l�Z��xf�a�b��j]X9�h�[ݠ�٥��RF�~���de)��ұ���<�(�`X_V������А02MA��ad��b�V���[��[�0�[F��bR�H0��*I�K�)�R��d�򾦳0[DoNCv|T��22ۄ��0�L,=u덶�n:�:'�ǌ(��f�s��ޯ�j���{�Kyb�(��F7\D�� �ܴƌ?(,3#Nf���f�V��32Wpv���$���"D���Gg^fe���S��ίm��m4��wm�v�J��++�3�Z��W��5�!�$�R�B,�XF21�v�*������3^�#�q�2�L�M�P�P������Q�၈���fml>�A �IBB���#�Oe},�R��L'�.�N�=p08$��j�6	̙���2�|��6�~׆�q#��ћy3�L�g��fi�����!�̉9�h����ˌ���[q��qƜl�n��O��Vk��4���_*���xn	�����*B���EYs�'bF%Jc5រ�,`ñcQ���(��M��H� �#O&袨�ɢ��\��a"3ѐ��H�������q]��)���Z��3.`��[1	��"y
��&�+֩��Bi��f�;�dnTf��@`X���Q.m���+g�+/�4�2㯛q������xvi�d�Gs�UU>�'``�
�d��F�sCc%ˆ����П���r-N�C����!�z��rA���`��4�ho��DS4�B֖Y��v�d�QoAy8řs;��@ٓ0j)�,��2��u��5���&)�FVf_�)�������'�����r�%���0D>�I��kTv*�I� �%�\��m�n��n:ێ8Ӎ�m�h���x@\v���u�,�Pr`� ��2CdY��6jRAg�x���2a�<�0�����`�H£qI�,2�~y0ӽ���b�/��?H��J��[jl-�cm�h��q�膡P�j�����bR����T7,}$��b|%C[,�0`#
��VI�d�`}��G	pҘ����O�&Ze)p�>a�H�������.$�4�:"2hd�(���LM0,������|^���K��~Y��]�n�ˬx�u�\ba`�$�0��a
x�[0�=�K:_G����G�[�F���>R�|:	�<|WD���GG��Ҩӂ��V�G���/K��u�:�e��W���ilz+Ǌ��x|>�׏��O�iz?A���Z��t�GL���X��:YSe�mz"�(L�"tDN�4=Vh�V=�:&GC::^���:�^���x�sm��0_G�i��zWG����6WA��z[��X�,uz�u�U����m�umhL���JG�/JWE7MR��W�SC4%D�S�
�s��r>n���:�Wq66G'��^iV�[r�$!�h�ܘ�:0�3(2"aNX��S�-��+hȣVQHտ�K�^�U�)Z_���l��Þ�W�*�oy�^tc�r�iE���Lu�Q�N�-r�U.�7�')Rڐ�kv�҂3.1��J��w30XWu�*fWct���Kp�l�X��"Dd�8�Z�Y1�u�R��s���1F��J�5��^grJ�N[J��,6Uqbb�'�c�Aئlx(�䱛\(ԏ?�`W�:!X�%��F�#1G)y�v�H�Ƞ͛5���ʭN�3�6#���dk��G۳W�L���r'�9k�v�M�����A��;Y�����̮Px�ފ��B���7,$��0��R9�.�ZØ���[�,	sr��vCv,�4��6���&��2Fn�Q&�ͥ���Űn��c�G-��tm����WS��+���ˍ�L�,�5_.ZK�	�`�6�i��>�r!���� '�*�,i����Sr�^��]s�#v�Y�]������r�[�ư�
<�8T&r�m�2�#c��^o�qt໳X��s;2���C��=��������̽�{�~�ə����+33����������z�s3�{�g~�̬��ǫs�wy�#�e��Yu�]u�q�6ھ<;4�t�����GMڛlڱGdY�;�"��6j�lݵetf�f�Kl�݊�b�;��9P1�m��c�M9AV�vUU޶�lm	\8-�)����Un�7fư��o6EL��C?�g��s!��gZ���2�7�9Y�K��B�t`ld��ɽ��j�,�,i`�IY�Gc�d�Wb����}9��}0!�2����eS��{wMT.ML�y(�,�M��$P�.jy���h�17Ê4щ7M0�e�,�Lra搎!�~���ո��yBE�vw��r�@,��:�Q6�D62#/J4},�9�6���6㭸�8ٷ�;>;4��{뇾�����;&f��ɡ��by&�T#<T��3�ME�ґƘ�ǅ�aMXbS�6�X|�Y2����e����Ew.x�Ht �D>02q��!@��.0��e���J,e�a0Q����Y���v�&J�c%`DĤ����2$��2q�b2P ���p�S�C1cm�^�螟<~m�o�i�m�i�Ͷ�:��lO�1N��b�6�]*����a�3vu��\�)f���.hՄѹF�6(��)1��Uj��̤Ԁd]�m�KL0U`�B	2�i׮��ۭkX�fm�-���91�cu�9�V��]�¯*�Z�>�'@3�ɡ�D�҈A���&%Ȏ䦌*�����6Xp�h8���U��z�\y4��~��q����}�ǝ��)R�T[��������Ɇߞ:�/�q���qƜl�jӧf��$'}����2�L70��n�˃"����7
�7��	),d8�,�j٢سn�sR3��NL�e�a�{�<>�F\p�94T: j�@�=�޷Ʈ��%�F��_�n,���y0���zM��9�L�
'�{�T��~杖����\8f!���f���7;*��9v�s��Cl/��L\ȉF�$���nv���V��aY�����[z���
�ѳ�����|�1�1x��z�o�>uƝ�L:'�ǈtæ��}r���n�j
Q��%oU���q�C��ě8T��,t5StM˻ni�,`�AY,x8�j��1�e@M�bto%�LFd��nP����Ï8�e$��ce�B#M�,Jl5��c�Hº[tm����i6Ef�_/���@w���aG^��ͷf�+��rs�����!�*��rhC�EH7�Ų���CtT#3=�6d�*xə��aRR�#j;k�����:��釩#-�����3��
��~�y�m��٠�&%��a�1?*8����ժ\*T7����jM"	ȕ
5f�R�=:6n�-T�IZ;
G\����s݅�0�Ùs��D9>���Uzm
��R��d���fc���O�q�\|�8Ӎ�mZu��Gi����c�1��	*+#�K�2��UR���~�����2���N�b{(�N���g���M10�#�lOT���:! ,���%��nmb���s�4p�߾��m)il�<l�=z�6�#Dm�ga6�0L�����7	��	��.z=�ns����1�����l��((�2��Q�aq8Da	Y�4-T�fo�{��6|��O�4���:�8ٶզ]x�C������?xS�{�>�~�U�ñ�T� �.T���雝с�����LLB���g%C���\731����YH��e/sJ�퐻%��届�;�a���7�2b(�0�c[�����������g
�(����`�(�F:�,��YP��pePP�pT�4fw���rfh@c�dY�^/c��=z�̾u��|㮺Ӎ�mZeׇ�31�����1�c
�3?L>ێ�:�ٝw��0�r����GM7jפּ����x��ށ±��꡾+����'�f���T9
��.�y�E:�FlB䌘�@Z���B�1K��d��%�.���
n�Av!S(H�
 �C���͟|((y��I�c	'�Q7 `�}&*c�c����ɉ�;u��4㏜t��gN	�E�>�i�)�MeU�WY�2�
�l���&5YJ�9���R�1�#�h���cU n�+(�xۮZ�]���̥` �*�V+]%)Ri�+$��yڪ��/RK���t&�V�E��XI�x̒��9��Gc���0O��.�J�ɰaf���pԭ�TK�]F�7(ܐ��b�ш\:*��f���Ň�&��C��O�
P��.p��.SCߗ����V�wTT���s0r[U�չ Q�1��!~|��g<�Z���C��xi���6pɣ��4x�î�뮴�f�V�~r_.-a�'�y	���&]���e�4,��L�򪪐<���曝���8<�զ���ˆ�f}�,D�����bžS������=��Ra���s,�n`�{�ɰ�gI��u7�30�<��R�d&�X�����V�R��!�seĠ�f�(��}�J��;�@�t�1.��`7	�Ϧg!�Qcɷ��=W��,Η���Z|�k��x�n�������]]�RCDL(L+�RO�6aP�L:U�+��Etz=���c)�F��c�:8:Q��6WG��GG��p��x�/�C2x�C��R���lzY��=�����?+cbt:WG��������=����S�Ժ>#'GçC�Y>���|M'���Y]Z*WE^���tQ�	�O4��<3ñЇ�C�2Y�D���)��~�\�WN�Һ;:WG�Ӷ��=��Ο��e��Wn��o��:���I���+�G���خ��<�{2&P�N��:`��ƳÿQI<�E��uj.�y�w�W|�8�$�����@Yׂ�*�����CoS���@���gv�Y����ɞ�=�׎v3��Cݭɻ���{\��w�~��̬}�ǫ9ww�������z�+����fb�Ux�+y˻���t��V�����rx�׬�˭:�:�:ٶգ��6|�����蛉��G)����`��e�ψJ6��9ȧ&�`p�.f��~��~�G�ꥃu��!F�#Lp�-q���qy�q�7jg�-[�����q��s�?)�sm����0��Y�G�9��Y}q�,L���~=���8��:tD�0釃ǈtᣛ+z/mUUUUP�F�:�+3㪍���١�A�}���if�est��M-��Wc��9F Ð�=<�>�25Į��a>k�]��;>9�P�8���ì;	���}cK��v�s<�Ç�<p�_~�V��Ø8�L�K�CJ�'�
1ʇН<a��N8ˌ�㯜u�Zu�m�L��ީ�I�Ҽj=I�(��W1�K���l1amoJ�G�Ԏɓ#��9EE�dq,9b��u�Z򪻚.�ma���:+�(dH�b��c�̔L�$�q�DʞI��NDnҵ�a/%��j�H<���5n6nww�fS��f�{�*���pX�F�eU�;�o�8�Q�Ʊ/5Up�b�l,�j\��s�R@����`�,��ƕ\7�Q�{,0h8J)>;�0�L�!1r�0�W�#q>N�{3��ǩ�f!�9�Rǽ��"�t�H*�NET�kv��t�flmn8u��~�J�i���X�.d��*���z~z��-�|��]m�]u�\8�ΊΦ^s�UU L���!Cyk�¼>rsG�B����`�2��d����v7�m0e���^LəBQ�����d��6{��u�YB�8:;i�i�#�
�h�a�	��>QL�FSqE|#���Ⱦ8hB�	�����H0��9sCO>q��u�[q�]m�8������d��@W
�@f
��% ���raI�ߕUT�8"{��= ��o�R��OY��
������35�20��p�:d=��������&[,�b�-P�GL�:�{pH|��s>Fl�?fYWlbr<}��U�ժ���GbUW	��]�G�U}~W��|re����/����_6�n�ێ��n�q�m��"5*L��1�c�WB��������J6l�g�$�ADsb�B}Z�?倇"������J�F���B�L,ѣ)߾sUW�(Fn*w�wY���O�B�B���5�L��Q�j�(J����2l�J]��va���?3�½j���f��9+�;�I��i�ԓ��X�M�=���T��q�n���a�]e�[hL?a�0A8h���_GZ��R)/,���I��Lw#B�5r�k��ݢ��
�B�6��.�Mm�r�,�v�ej���+E]v�2Ie��4��@cai%A�����(��Ͷ�o�nժ�F�b��NW[E��Fn����f�uV����4f��ᢍ£
(GF��r\��P��`J�����\�'9<Y��I�Z[���`��\3,�Ϝ�Uj�K����ÊƥgK����}x��֟��8�&လ�X�x�>g��9(�=�n�ꇸ*-ۛ&͖Iü�f4��Ba>����~Q��HM���GO8aӎ�ۮ��n�q�m��$c�%�Y�A�z�����S���7����y�	�`�>���o����b�/��N�p�S�âv^"����&�.D�m�,��z�i�6"'bQ�ӳ`J��v�繬YX�L�Ac��6�/�.���,Cg��`�5+��C%ʆ���Aa[H��0�a����hbz��ǯ�?:xL0��"C��YP���w~UUq �a3s�p��<U�2%�A;,��h�9���hN��Xvb<�����3�p��i����p�:M!��ǖ���bMwu�%�,��i����M������[0'�ʟK1�Hz��*�����!̸vy�/�Y����-RQ��U8d�/Y^̙���a�Θ*|�0����G����?��_�.:�i����]u��6ڴ���V������K"�D8��:�(밚�jl1��ߕU\D��V�^�Y4l���ß ̙?7��fv!)��!$?F��*H����#X.Z'�U:�����D�$�|�ˇO/O+��*�p�"^��H%	�$�7�Z���g8ddN�N�96����1/��r&DF{�j�j�Bjd�4P�IG؆e�E�0����!��(�͏���V�a��>bi�WW��7�p����W��luv���X��u���JI�l�&	�%a0�XL0��BtQ�,��8:Q���N�U֘��x�Wg���u�[��^�D��z`�C�zt���GC������=�����'J��lz=:V�����^�����S�)tt�GF����:h����`�O)��(A�ҩ|P�b��D�<��6t�	֘�].�궽Y��z�Z�_1��L�WE>+����|W����t�?/CC�zv��YҺ=Ӵ�:WD��=+�8WwMV�����=��ة�M���b��Q�^Oͷ�*j�~������uSC]7ws"ݫM��n�.e��+{���-�i��1ʝ����+n�cY���+aJ<%�H<lY�&#(.�[� �6��[���UD�\˙�����A\�Ɗ���̱�'G3�/��.^Y�Z�^߽>�w|��~���-y_T�]��\���d��I6���ج[�O�7��ެ]�\�l>3j�V�%CqK:jT�&�˒!g������ոG����svWz;p��j�^H�Y_j�!�<���k�bi�A�cJ����{ٻ�W��;�N˞=�M��b�}����b�o�؇���:��.+*�DWO��k"�.,�5��V\㌟z����>o�y�Oo��w}��n���OYtt��n�9�
,^35�޾�#��[����{��z��x&e�j��{rw>6�����ߦgu}��ם��o�Կkv�Ok��`����'}�{��0۾��~f�wz��N��o{�R��w=���ѓ��f�1I���&��-��i�W�o|ﻤ����nJ?>[��71O�;{��*���������s�~vt6bʧ&�*[����M���>qT��3�@GZ�M2��"M�HKFYV�,�(�Kb�W�E'r<�m�[��]�o��n^m�����.�t�Z7�+�4K��rXF��.��(9+�Pvƭ��Z:�F�ʚ���(�˂��B94�L���dr��^��E�|Q���% 6�������$��AIy,-��(�tR���FI)��3�ʫ��t�qⴭ�.�331Ҫ�ZV�w����UmZV�.�333������]�h᳅�8a�0L<<vp�w�<���]�v6l�"0��rJm�-ۭf]-��&�K��aFܦ��[H�Z㬬v�[�V4��Sh��Kx�ȐA*kaY7uDR�컶�U����ͻM����eۢ����fv����Cz��2��m�l�h�Z6�*��:����$R%�\-f8f;J,N�0h�(M�l�3�pXY�*�̔|/�Vyy���{13���=Ue�.S>SP�2X�2�<0Tab{�w-�鞹�7*1��D�]P�Təsf ��3=e����6�����ǎ���i�q�]u�Ͷ�=~9���qdU�UUć�LK�S�*"0��-U���Wf �0�陃й��-���XX����~V#
�!�v,y;774�*�/�Kf�Ul���H�����!ŸQJ�g����3xC��p�9���2Q�)E�%HI�EMfm�=}�L>x㭴ۮ�뮺�����g
s���-��]�����3�ĥUWa��ȕ;,��2dK��n`�[�5B2p��6PɃv.�z���E��Q��ǕW���͝z��N8�F�Zi]�n��N�mpx���0"'��K��L�CF��3/C&!����FDr��!Sp�)��dT�TV vY]\N=&�gǏ�L�L0L<x<x�K4%^h��G�U\H��<�1d�H=a��	_C)�rjP"s=;��AGm��Q"䛮�~�2�	�{;�S$��P�49�`�,��
'�!�f�bc�L ��S�h׍q.T�U�ab}�5C��;*	������"H`���?â~&`�<<C�d��ZՒ��f�*����0�\j�Y%���#x㛏.�$�Pdr���f���'j;VɈ֘�MR$��2J,rT	���:�Äj���6dڧ1��1���UW��ǲIZ�B&���Q[\�G)�l�ʚlm�[�����I���%C㣐��DJ.Qf�>򆏕Q6pFO�ڦ�!�5;�B�	��B���zl��4U�fDF��YG�/G
/Z�MST�Wwc�sy�'��+�z%	��)٧Y׹â^�)X�X��]��U� 6ڰT I�j�F�j��^?G�o�ʮ��c��Փn<i�ζ�N:뎺덶m�i�蟫 fI���UW���:4D�,>��T��IP�T�T,�,Dgh2a`�&���s���V!�p�
�R`��/ަ���wWr�C�r�7
�,��ڿ�M8�I,�,+$�٣H�U-J|��:p�%�L���z��Ѻ�UaP�=4P��.xa��eU��X��q�_�m��4��\u�OO���;���UUq!0D�t�&:1T���6%���1%	��\:�QE<sFL���˸}(��g�d��$���$VbB~f1�Z��ƷN4�Ӷ~eXa��x��R�M	E0�#�DȘ1�2]��Gf!�&����<�o��z���޵'#Q�����,��"t�<x<x�Nu7r�oj��$'>��Ә{�0�4!p���$=�ז$r�V7Z�(m���͘9H|p���8���Ӭ�Ě2Y�ϕ0`D�7L,�E��_nJ0b56*��i��DD��G֯٘:3e�^��lO��n~���ñ)����}�/#����θ�N>u�]q�ג��V����lxXH&JXÅ��i5ja
�+I�;�R�#x�#�ر�[�MM�"��V+L.T"5�
%��tMstx�9��R��6K���],:D��_�U\Hp�7�khu�j8�r�N>R@䱻[#�ۉN�|Çg�ϳ�;!�J3mF�sm���'�o+L0�un���2&(��W��J��2"#*}�`��P5&s��B����؝3��8;��g;P������%;���R�%j������
&���:�m��.��Q��6��~=��nU��:묾q�:㮸�m���.��i���EG5Ђ2߮Cv2�P��olH�8�lcX��in��*������G ���rIJp�c��0���C����h��"Q��'���"j��Vr�:j"f&�̳q�����v��m��%5͌Ҍ�M����"5L�74r���'R��Æ�,Љ��x�0tĳRu%N�h��UU�M5�����L�靏:'D�gY(D��tO	��x���4"&�D�DN�D�P�,DN��x�8&͉f���D�BxK �"P��"tD���:X�%��6%�BQ.O��<!����,L<a��!�f!�0�0��'���D�(N�O�ㅉf�AA:A4%"l��ó|ּBUTh�����1�{���_����~�Sz}��ߏ���}~����~��z�����]�9�O=$�|ry}%^S�WIj^����˭�oj�/U����v�2�O}7��ʘ��GK��������������3�L�I�3���ݝ�7n}gG��f��]�'�wd�f,�euZ{�s�>��OG�?��6����k�G�߾��,�<L�v�@Ǘ1N��ܡ�{���]-�r�333���������fff�3U���]�fff6��]-���gM�,�Θx�&'�vtK�ڪ��!�4�Ek�*}?>ȉL(�Fx����Zw8t�'䚅1����Hx}���m�ۦ�n��(�#�ĊJض�ώ��s4�&�%˃:�)kg'U.�9C�D�9E��W)n�3P���8`K�,�1=/�T�!�=.C1,٣G�����a�a�t����9��t�ܫ��w⪫�s�)���)�~�8'���\�.dFw���Յ������:��N	],)�s�g�#F��[�Ʀ�V"��O|�ri]ɡ=�[����(�A@LM�u~i*�/��*�ȉ�xJ��|c**(�D��aa����0���w�c75==
4#4��}��i�%q�Oδۯ�u�]q�\uyyyɮ�R��c��R�)[��v�D�Y�U���z�6�Db��ƥ���ڰ���q�N��J�Z̆7$q'�^EH������V�v'yT%N4(�l�p���%P������)ƣ��IlIr��ʪ�$5�z��+T�KH�׹����Ӝ9���`�]�f{��"&<��0"_ڹ�����٣"p�֩hVUxܬ�
 ���2vn�#�5H�4r2!D<�l�YbT��r�EXP�j`�6���	������|�6�]s�0�nw*���s�2}�������e��v��15��6q�.:�:댶�j�2�w����#��⪫�3��\<��~ӄ>���X�>a�"x�a��w���{5��&�0ffh�8�faY�)M������ӡ���B��r�ڍ�+N�K9N@�8D�x�F̉�8�aG�뱕\<X�����Y��'hQ�F�IN2��.�e�ϝq�\e���4|Z� (��L�\1X���̵ےGXٙ���UV���s|�4����!5:Y��	(������'��ٸpЕ>,3���$DMvtk-˫��)`�ؔ]UV��.����&��T��SBr}��ѨS<yu	�`L}y��]U����3>�3ș���1i�{Oʇ�$��s���}�m��;��<`��٨���y6���>e�_>|뎺ztxxxC�;:>���a�^*���c;���f�u��;��.�Z�I�8��%|���]� ���`�]���jRP��Ss=��|63MƦ��!u%7�L�f���d�Y(N�>�0[6��fDa�n��N�'D>@D~�H�$<�7�mTx��^?8��ϙ|㮸�������	���'�ůk�b��i��Ijj�(X�*�A�j9]�(:r���1$kI���(㶊�Z�1;c���Z7F@���2V�r:��~m��ća��i�	���%�Qqmp�Nw���	ʞO
��&B̔g4U5Fe�MR	���.���*���|^�\f�ꦒ���31;�k��)����-x�u	P�Ԙ��%�0�&d��U&��>4�jLԲ{�<;�I����9�6��b<x����W�sQ�ǌ8��Ͳ㎺㮸�-����.[���U\c��d�3p�ɬxC\�[<MO�2�^�Ǒ��e���h����4L�	��V:*����,���>�˞1�KвE�c�V0�Pm��\�^Ĩ�C�PR�,-��	�������+��|������6�
m��jy=�x̹���b���G'��æ�|p��G��>:t�ᣇ�F�F��V�ݥ�ٹd&�Ҫ��u����3��e�fm��s�#�g�%};z��^x/��Ȃp�\2{�~��+ӧ7���*�\,�
�!TH�#�R��RD����t���{�H�we�\��Ȟ$OL�K5,(�5\�ʢ�\>�77�������<r{���^G�_=q�:�n�뎺�o[m[a�Z嶥�U�1���/�,��$c-��Io���	1<!��9$3�$<Oޓ�!�}�'��Ξk`ŗ�m�e���2���,+r��t�4��z�e��Ù�!g&�/�OC��D(�/:��gpl�`��QJ��S����vf/vR47aJ����_�����ag��Ի7>6`���m��-�m����q����.2�BtO�A<'���"'���� ��DN��4 �M	bX��8'��b%��6&�	�"%���� �"P��"'����ı,M��L��X���>A�%A(K8P��L,��0�<y�_�q�]m�[u�u�q��4'����8X�l�AA!D �d����UZ7�Gf"4,x؀N�U�fF��E�eV���v1�
�cQ�2<�q1�&�,�%ݎ��#)w�eL)s,)9�x���N����Ѻ]��]��ݥ�H�����UFpBbZ��EN�N4�+h�k�����i��-�m�r�)v��>uF�!Um��B�S)H�(���Idu���m�܎�����������X�dV�ݚ5��MZ���H�m�0ٳt�߱<�<8,�����Y#����h�1�$��rۖZi��*�Q	�=�oj�xC�z��Ҝ_��q��rѳm��[�e��K5��Wr��ij#+V�dTKU�V�ٲMH���%��披�4���;�(H1��K�6��4Q�T:��G�-�6�;A��7%"m��ʜX��`Ь�*E%j�B�����h���\��+l��º�Il�J,�����mIe��9�O�r���U�wy�����mWj�ۻ�����̵]��n���3331�Uv����k��8p��`�&�^X�����V�z��~��%[��B쬒��(��b�V�h�n���K`�t���e��(���$n�GX�*d����j:�BƘ&���I�EE"M���:�UU�.���R+
���RX�ԣ�N�ل^x'�gga��5����`�o�2zzY�eKd���*àX`�u,�֎�3���'�fe��T�
�긆�̘��2dw�y��y���=��}v�6�fݷn��[4���S��nf��ì�)6p`����4䫫[:x���>q�\m�m�l4�N�Ŵ[r����p��;ϽÇgY��^͜��-jh�}�9Oٛ��=�y3��X��'��1�^��Na�hS���n��Y ���ܬ�"&���'Ӭ�3�\�&��ڸ1>�.>G��֥�U\m�\|�l�~	�a�x�ǈx��{$/|�����Q����𺴝��������u
���i�ݭ��黝3Ӂfe��0��k�:������ئ[c�W�[�ҭ̵pMud��R�����d����wW�b�!�gN��Κ��V\]�N�pe�͛����?,���y>e��]|��\|�n�덴����vzY�qg4��UU�ɕ�$���=0��5��ч��+>�md����-o�]���-�kl[�1���}�ΰ��;��ͰXpٳpJ�t���2d����g�w$���!���'�o��,���C3�!F!F������7:�Fa�\jf��0�g##Sqv�e��q�uƟ�m[a��p���O�`\c���CoX=������2op
Glq���������s8���mS �r*D���"�QU�m�U�r�i�Q���']��[\�����_6�W�^[�Ml�R�K �B�=�Ag ��+�)i�P� ��b�~�]nݖ:�g�w�ˀ�g1u��K�K`��L��9��)��\�A����J:p�I�r�@��i�,(��iVv��M��v	t]o�}���|�Γ&����c���[��ߚ|ˬ��N8ێ��JxxC�;9�c��0'9Ҫ��L?d�M�g2W#~���}>�O�6�K��8{5XqeP��Ѩ`�`&g��)�(a�����UT8v�}�rh����@����蟘ս��v���
��ӡg2d}<L�J8��y;��K-&�* ���S))�%�f���[�Ç�0O	�������vS��?������' H~�^O�p���e��'�=�˜0��p)��)��	�WҒM�R�؇�&��S��D��c������730",颡Tqg~�L������F�Ǳ���L�c�V�UU�C���-Ql�Qg�:㬺�N�ێ��OͶ���ө�9ΕU\y��8���zL���鋔YgafgЩ�W@'�5�豑�4���D�J�,9��e;�=Ί�@?w���g�ڳ"*n�$=���s�i��B	�K4d>�����|%*�!����!��=8{ޣwv_TrNB�Hx���>u��Ze�m:�n>t�짇�<��w�a��v�N�)���GZo��v)}��wk[��̮�Do^ZH'��l����1;�ԭ����)X�I��c�CD���ޒ�q�)���r�MNn�򪫂r�\KT�K'H�0f��;"T�</���:;�2\��
3�}CEPв�����EϐOCu���J�d��3s�3��gs"xރPB���樦���zt,0y7�jB�����N:�h����4"U%�z!��Y�Dެ�n��f�q�N�ۍ8�n>>=;)���<���棚��l�l*Cm�%we]��U\��|Lr=j-��>���9\�rt�`�=qK��FT��r
3%�$�B�L����w,��D�� �)5EEk��0q�ږq��Xl(2��$Wp��x{���'��4V�n2:bw�`���a��|�a���?<uǮ4pÂtN��tD��x���<tN�P�D؈���J4 �M�<A<'���&�؛4&� ��""'DOd�b��K�D����ı,M��BhK4x��R|�(�|��BY���p�,�Cǌ0т"tD�0�a��0Æx�Ŝ,K6P� � ���	�5���9u�桽d߭�ݾo�'��^�UY����W�>�s۳��nE�����.������M��]��0�?;�rO@�����:Uv����fffc�t���fffffq]*����fVffffwU[���̳��8p�0O	�	�G��GMVꪩWy��C�|�<���喥i�����\MɊ�yb��vz��j���3|�����ֲI������S��ԧ��{��[���R�f\��>G��?G�c]�g�`�8x�.���g�,؜�e|��Z��Ԝ�n�{~i�:��\|ӎ6��\i��նm���h���c�UT>�!F&�9�d0`L�AN���NL������z�\�iY%�S�V��>Q���E32]C&C��<{<�~��<�F���W#S�͜o����*���a�����v�9\f`�F�s�o��签i�Ϛu��|�?6ڶ�Nc~'eU��8�Eg-M�v[�B�a�p�T
+]b�
�[Z�"��"lm�]�GmcB��f���l%��t��Z���N)P%**��(�`'H�{�m��:�V^�v���n�ΰ��|�C哐�����ڵ�w�g���39=�8vbp(,מ�}R��ocUTу2�.3]��w1��d�r#�E͇�|}����Fh�x�ɣ��fC'����b{0�i��]�m1�⛗[���Q���e�t>�z��ok�u:�׮��/�4���u�Ӳ��Nχ�_���]e��ꪫ�M��K�CE3M��%1�<|�e�LwM�p�@��+���1�#�5 ʽ��ޞ�������,7Pnm,�vٳԶCdV+XG����$<��<ݟ>[>���33>]�rd.C;�
�ii��j�70ی4��Yu��q�u�e<<!����ꐙ$��Y��n��aIk��J������!�Á {��73,�ڡ�j�\��w�g�NK�J��+��J\[�&�,MJ��	�I�a�������r8�=���?G_0z�쟁g�L���~�.P���`1��6��o�|��q��u�~m�<��gp�?#��U\<?}�Ϫ�U�K;6T8	���2��_b�R,��d֓un��Z�0�}�fI���l�0�;��j��14x�11��S����f5�l]FO���;1�+)��)�7��j1;�ӆM�,N<t�<&'M<C�5�g̯��36D$��ݒkQĶ�B�*�E��hV�����ݢ�4�7s��3�GJn�,��8lt���#��GtV�!]�UJԎ�$��C-�Z���m���r=��v�&�Z�^T�՘�VҚx�&`ϧ�6}�unkEL��ƙ�G��72g����k�y��������2z�e���)�>�C���O��Ӑ�A����0�%nB�m$���}��a�$)�dX迶�)��ǰ�~{?x�׏i�[i�q�\i���x'gi#ǥUWľ�9�0;`!�t����,0:�>�/ت�Z3?���^�:��d�N�N������Է����(�8��!
X�&���9
���q>�x������e�p��nOc/��o�Դ���ʵY���q�]m��6㎸�k��^Mu{�<�d''\�2��6�n��>��TSP�a��	8�T��OESc��&jY��~��^��M6 (�����+@�A)���h3$7��+�Qum�n�*&{MV麱!���l�d1��UF���ԛdJ���>e���2��O�m�|Ҷڶ�K���X���&6RC-��������g�v0��g�v��Ð6�%�LN�R�^��a/
8[*��٣�Kn�SM�;ì/�L���x^�T�O����8�A�³㮲6ˈ߳�m��=3:|�[�8p;<|-�ȣ-i�a��	�t��u���o7��e�,���	�:'��tD��tO��<tN�(D�B&�DDD�B"AB&��<'���8&���f��4""tD�H'DK4"pD����ı,M��BhJ,M	RO�B�>Ђ�Bp���:lL,�Fx��0ق"u"t�H"&�D�&a�	af�AA��;�z��4j1G}��a$rdY����2��'�n����ޮ�G���nEm�KxKܔU�]j}��OL����o����v��,S�	%�M�����z<��Z�na˘Wy+�[^��vU��v7oY$�N�;�y��]V�x>8��<�1j<={=�aSk{wc���>䓹WZ�	�8�b�ӯ���s3�B��vH�ojx�nV��{2ֽo�ݣݍ?:��/�	s�nޱu}��o��e��bܧmU����� \��E�ن����;����}V����܍9��7w"�r�3_�n��I�Kf �~v�gm���J�/���o�N�Ǫ%����<�,2���`��-�Ȼ�64����_-�����)Uv�r~�#���d��U+�4�-P����]ZJZm��Ս��5�ه��V�C��Qe%�l�3�I�lp,Vg�"�W["�ҏ#��#������WO�V,B1T�m��ǉ���7����D�$Ah� ���tw�F�f����j2���k�3_h�W��$�߮�/W���iUn���3(������J�wwv�ffffgV�V����������U[���2Μ:t�Î�Ӯ6㍺Ҷڶ�O��g�g��?f̊�2�E,d����.��78R�A��I��+�N7Ij�;���"R"!WDܗ�2mWK#T��A7lm�f�ڪ�-���\%I��@rX���ﯪ�����n�Ѭ�m��n�u��6M����ԧfg�p�����P�oW�{� h���0�~�$"�gxs����s����i��r�*hp��d¡����d{��Ei�|d���8h�v_��>�b�Z��kJ륌,�+7�ΰ�	�fxs��׮��L=e��e�u��q�ZV�V�պ�T��Kb��j�aP���0��gCKj��f3�j��\jL����|�y9V�41� �a��Tnx�\�d��o?|��v�n���lv.i! vc{�MN�C���̍[M�s��UI4zL{��QM�$90w��>�4�֞��-�Ӯ6㍺ҸpN������6r�SdY,5�,���o��n��F����<=˄À�9�XVYH[gͭ���Yl���`5�S��/s��}�1��F�yxy��^{-b�
<�>��iI�r���A�J�99=�S/[~i��\q�m�:lN�mPu
�4�ʪ�g��p��HC�(S�\9�)�����%C!�n�3 ��R2D�\
V-�4j	�x��S3=�f(5$>�����ȱ�k°�qcF�1t��bmᙿǯf�T_C�:���C���>6u񬢛��[q�O�m֝q�m֕�ձ���'��.�狮���NV1K����فѵ�ɶ��fG�u�5��;Y�Q�
6�E���fݶ2n�h5�
ݮ��H:�Ket�̷�Y�awv�BZؠ���v�녜�*,a�s� R�8Z�Z���%䤲9�Q�Ș�%(�(Y��F�῞�SLQ���r�)���'b��WTs3.b^STU&Ã1j)٠�*�f�ɀ���4�~��#�;v���a"�ōF�~/y�t��ɻQ�g򪒫�N������e�8ӎ6㍺Ҷڶ���]�&�x�M���(>�S�IT��9;'M*w���$�J�<�ǣ��q����|뒞L80��!vϽ�Qmݷf�5b�)�[vlJ��N��诡�N`P�La���~<D�~�m�Z�ŏ�||���l��.���q�����0�����vf�Sa�1�A�.L��>�f������|�T�U�5	&��ֵX���pc
Ë2��3�$x���mռ�Y�S�B�������>\L���z���4�gM���񅱣NUU8fIӢh��8xâ'�Ot��	�e���PiU@lɝ�:x*p��Ns��~���^�O�0�bz��K��^^��8l�Y&�Hy����?A�
�C�*t��|��XѸt��bn`��jX��๠��.~�N��&��zqA�罆>E���*���1��m�ϝz�.8ӎ6��y~]B���TG����
�;nffa�r7d���&@�;mvs[�lv�F�d���w�����l�Ƴ%�3�0c�e�dTtv�p�\����[$��փ�k�ƛW��� T5>�4�J�u6B���Y�wu��u�$?S��Gg��8C[�}2geCJ�d��4Ԫd��f���6h�1w�����fd�&N
�ɸhɠ�Ź��Ex�/,���NJ�lLQ��pfx�˓p,�C�17��YW�d���:Q��D��x���!���s���ْ\q�Y�)xKHC	pV±��o���;8j�pnK;���������� �,�0��5vh�bJ���C3�#]�jUbQ�f}0��a����9�
Z���[tm���e��F
xvvݾ>y55 ����Sǆ^U�ɚ����N?;56e���>m�[t��tN�㬝<'���"'���Κ4P��<'H ��6"'	��tN	bl�Q�Bh���:"tЂ$b$�'�D��ı,Љ��ДB�I$�6	�	dԖ7'D��6l�?�!�0�,�<'
D�"l\q�m�u��4˯^0�ӧA(��}Zod�u�sW�ק��-��n�u��w���e��\ݎ��m�����n��.��y���wf�eTg�)����W{>�vU/�w�[ъd߶[/�Z~X��m����2�u�O���:�:ȴ��u�|m[r��p���_�Wl����V�J'��G_������*����������5�մ��_w���q��7�V5�^�����{���{�ʳ��ܻ׷��|5�,W�M>ǒ�w��͝~�O����~�GZ:7;��O��}�x�m��{�7�{��X�;ݾ���}帽\�Q}�{����w�O���������[���
�V���]��{}}�n���n�J׽�}cWʿ{��vN���>�k{;��c�5��_���5�rW{����{Ϙ��wwnfffff>b���ݹ�33333�U[���������V���p���:t�0[q��i[m[i���m�,�Kk�lO���4��tx���8���ݚu�w�M� ��k���wf��32�v�'y��|/�4[n�ik%Ҳ�E5�M�d-jYF6���

$�h�ϻIU�adЗ10��̗3G�XbXvnT��tHfw�kL�yWm����e�u��q�]8'�=�.t�������-T2O3�����Ӈ���OǗWMݦ۪Sr؛-d�B�kn�3Os��g��oѹ��ʫ3�F�4l(�Ӆ0lѹ>8�c�ٙ� ��10|�~�j�惔x>բ����@��$ü9���]GO���aX������|�-6Ӯ6㍲�^^B��/U��H�Z��%�u�n�T��E�#v�ʔ��M�6�cN�:�"v��h�]o(<*h���Q��4�&YB��S�Ƥ��J�Q�)lLT,�E]�� �]p�n� 8��*���#Km��,�#0c9�)�.`+"ƌ��58�43�Yq��^�~�Q�u�Of�L�o?,�:|l;<bl���6�Z�c
��aa�s�x'�҉���>V<RG����U+��c��,v�F.���+v���:4����y�}rڼ_�+M�댾q�\m�4t8pN,���e	��L�UZ[-�a�j�J(�+��`�6QY�D�}�!"��S9
,��P��/)���w�r'M�_�Z�����:d񑘆B�Ջ�՘��%�[bi���"B6R	�J�DV`�r���p;��\5��,1eTF�F�8}�Ě�����M*��M�ˮ�델�l�m�^]Q@�!���Pc�F&���o���E��G��L�'�J�(�DT���2`��L���Zj�%��5��FHΰ��:�!�ϯ�Jz[vg~�ދ�hF�a_U4ОH\�h�D6Q�x2>J2u$�,�Po�0М:x�t�<"x����8l��ζ�)�����"��f/<UY�Qߺ�%%F��a���[���
V��|eS"!a�UQ��*�����7-����/K|�wUu>���OMO�=�\�����̤P�_R�F͌4U��B��B��'���EϏNMC$�S>T�ﺵ�ѯ��t���9������m��=e�ʹ���i���V�~mp���a��:�G�YSB�5�2Ie���a�f8V�r��,�F퍃�˒?[.����k�ԏ%q5H�+��8�n� ����-N@j�3#cƜʜ-��N���˕��یj46'�hvD�SD��q�*h�G�쓘_��0���®rP��M�0w�	U�f?4Ya�|�.�+bjQ�Ɇ&�SK��̸&��4ߍ�=��~Q�8�B���9��D���E��S��P�T<8v���4���ϙq��q�q񶕦_���U��OCD���%p�����]+EZ�U4gfͥ§�60��&����Jj�8��=��0������i5ģ�,i)���-"B�}508��'�&���`��e�Rj{<앦|ӌ�q��6�G����gE8a����R���j#�y���,�.��%�4�N�G�<l����`�J�$�%�'���8O:;��kOnۣ$���I.�LT�HE���˧Fh�
P{|����MN�3b\�:S����荗�4vY���ʓgHa��&��,�_-�8��Ye�u��N�O�ò�'���dk	��Q�A�mS��F����]�A��.�Z��՞Ga�rq�5��i�_�p���H��$�B-��+$��FMLBvfb<.O�M�8�t�277+ҵp�7�p�!�rL�(��3��K�c��`���LUk�-k���wB�sL�3#��>������ʪ����H��s����=����}�ŉ�Q�T�!�e>{^�L/�f�@E�l�؋bJo��Rʲ�1�$bq*"! ��0H�#�#DD`��b�F �#YK,R�X��YK��*�,��YJ���*XA�1
�$��`��K)b��Ub�ʖ)QF	#`�`�F$�RʥX���RX����T�*�b�R�,���K)b�URX����UU�K)b�URœ1)b�������K��UU��0H�!����`�R�*�ʪ��V*�b�Qb����*�eUYQUeUQUK*��UE�JX���X��*)KU`�#`�Q���Db"д��"1" �D�*�b������V*)V*�b����*�,R�,��T�EU��YUVU*�UE���UV*�b�V*,U�UeU,����Q�"2""#""0D��0FD�"%��U����J�c0U����UU�������UU���UV*�d��YT�*�b�V*�eE*ʢ$D��Ȉ#�"#""0D�"2"$d��J�����T�%R0D� ����Ȉ�b""A��1F$b�U����Ub��aV]��"#�F�0H"0D��Č��� �Ȉ��DDD$��"1J�UURʪ�UTURYUV*��*�T�Qe*�UTX���J����DH0DF" �H�`���R��U�Ub�(aVUUU�R�R�TUYT��Db"0DB1""���U���)J������b"1D�"1 �F"�D��b"1"#D`�dF��D"#�DF" �D`��`�VUU�UbS
LQd�*IE�(���EH�ĔR(�E0��%�ED��Qd���,J*IE!B�(�(�~	�E�$QbEB���QC@�`�H X�E	E�T%DQd��B��E���P�(�%J,���(��X(�QQ(�B�D�ȔX�*IE�(�QR(��E$��E�!EB��,Y�
E(�QRQd�T(�QB��E�B�E
,P��(�X�X(�J
*J(QH���T(�P��B�QbQH��IEE�X�Y�
,U,�0��JR�U,RU,��e,�1A�"��" �b�K�R�,R��Ih�E�e%��K))JYJ�R�J���)b�K�J���K)JK�,)R�)T�J�JX��,�R�J�R�*���J�JR�)T�R�T�R�,�)b���R�)T�X��Y)T�R��R�e,�1PĔ�YJ�)e*�JU)Ib���R�)T�J��R��*�K%(�)JX�)e%JX�R�R�)JX�R�,R�U,��Y)d�R�J��Y)b�JU,��X�)b���JR�)K�,R��IJX�)T�K)d�R�K%%R�J���K%*�JU,��JR�K%*�JU,�����D`� Ȃ ���e,RU��d��e*R�U%�U,�<�`�JR�*�)T�(�E��R�YJ��U,�)T��Ie*�R�,R��JR�*��*�R�e*�R�T�R�e*�)T�YJ������E�R�)T�K�X�)b���*�X�))K�YJR�U,�(X�R�K)iT��i*�Qb��QiT�����YIT����R�)JX�R�,R��JR�*���YITYJ���,�R�-*�R�����E�R�R�eJX�P�JQe*�R���L,ŉeK)TYJ��*�QT��),�i,��Ie�YIb�b��J����(�D�Ib��*��YE�K�(U,RX�b�b����G�ǘ�1U,RX�X��E��J�b��K�R�),RX�X����%�K�)RYIe"�-,����S��K)RYB�<�<�`RYIb�(U,Qe%�E��YE��Qb��b�(���TU,Rʖ)e%��R�,�*KJ�UV*X���R�X�e%��)b��K��D�I�?ɢ�3ٯ�ɗV��0P���ӌ�1 A1P�DAI! �wB�$��U���i���g�5��\�u��r�Zk�W���r��l��q�:���g�{}�{�,��{���+����4�Qs\`�'�����7����z�x
��^��P�`?�܇�DO�@�|�@~cH����'����|�>i���J�e�A?���t�?�'od��QTO�O��G��	 d���<R'Oy��@��!f'D�~�|JJOjg�oi�k��G|��x�2�o�䗆R�`�7͎��"��(�o�d@l
^
�f�4��1� =Qv�h�!"��"	"��|˾
��3�ZA*���籀���S/����=O���)T�AiT�AiU$�e5�� �J���  ��r1�}lD��̸?x�����Pm�W ��u2��}?��Za��HT��@gR���~3��G�8��<��}��/�!���G�}����0�n.>a"}����_k��xn�Q��z�Ȩ��{a��â��}]�q��f���~�z����*��{r�^��c�`ye������-�rM~�$���!�4��&NK]rB�Y�p��Y� i�წl��9CLª�I)(��%=�D��rs��m@�g���x&��O��T� x|z��(Θ^�**���!>Dx''� <�{����nc�>8,�l)��N�T�>d��r��.�>�{R
t(�#�>q���M��qQT���J�Z��޾EEP���4�����i����Xq8.�/�93�Yyf�i �%H��˘ܸ,P\[��>V���� �����;!�M�X�a1�n� n6�n��QT	�'!�;�])*��:� �����4<�0|�{��Dܦ�$�B��p��,���x&8oNPB(�	��OE��,r\�)��r���f�'�J��w��LbfRu��z�$�;��C�*�,�)�������]��BBES`