BZh91AY&SY0l�۵ߔrqg����� ����  b�  {�                                     >  7�`        �              �             �                                    �         JIW��5J�DTY��DťUt 9�R�̊)�BEbj�*��R��j��1���   �  R��5*��+�3�P��� �)R�N�u<l�T���+��I�3�R��2�4�'8 �;cs�9.m�]�73]QV � ��           ��sc� q\�8�
�` ����^���\`��s�r�6P�r� pFlsj��f`  ��PA�ӈh^X�B�� �LNᆃ�C��݌��Š�q� hR��sF��C��.�ɠ�pP   �      �����gjR�cU�j���\��T�g ����0*stĸ���.gUAv� ����� � P���  ���G*� `� ;���`U�h` 02h dA����uC�PP���<   �         $r �07`9�V�@�p ;�us:���@UfX  �T@�   �^   @�C�  ��9 �1 �d 50 0� @e]9 r,�                OcѠr�w0# � :#��w0�9 21 � �ꁹ�����  �   ;����  N�ɠsb��8����@0 ;��4f@��@���)@�   jz�*� L��& i�Ʉb)�M5)*�d`F !�`0��&L�2OBz�&��&j<�M����T�
J�0�  `&�  �{�5�U(` �     &R�P)T �&�@ 7��o��@y%0�1�*2��S9Ӗ5� TEh`�kX*y�^s��D[� �����0R���[A��|�~��|�����s�4�vgt(
"�5P��T�� �"����h%�?�.���AWD<��ZiO󇠷g�e{��zX *w�A�`)� 2`�����%  w��@�b�v
7b#v�b�]��؈`%؊F�*݂��b#v �*݀�v*�(�`�]�,`؈b"]�-؂݈-؂݂v بb�]�1��� �b ]��v �`�v*؈b�v
�b�b��`�]��v� !f*` f
����*�b����]�(؈(]�
%�*�\*�2���*��4hǧ����L���/��&n���s�wL扄�Gdт^�=)ǐ�N������^�=���:ׇ�L��{/��mBƜ���P6��Q�fn��I4��|��b����p��z��W̍w������Q�{�B�j�o<KeƊox⧱���}J<�C��Ə��nF�����K�R��r8:��^��f�Bb\�c�����{ݩ_��f�MA1��Ӕ�SEЮmߴ�<�F��@ao���!�F,C��v���@�PC�pvD1�Yj@a���-�	����k�*��d>܋{��/&�y$�I�`W�[�@.սqIG�9�BE�=H������}{WCΛ�%��Q�j���}	o\�R�oӀ�o���ie<�t��^_��xӄS٫�{�	���8��"�q0<�yJ�1�]rԔ4�;�㻭.Z-�7a3p,�f͓�� �Dwf�]�Sݺ��f����:����v�7�磸u��n>��5^�8wt�q�bI�����5��� h�*,��Á�2R���e�n�8{;��xȤ��8��ܺ��ޡH��5�o�t��m����$�Ź�+��	��p\xz�|�'7$\m�b{�uSUק�r��j�d;��P= �����u�P�[�pc�N���@�$N
!�u�qڻN���[�43�s�)9!7m�r����OgD9���ʦ����o4��f��Փst0b���#Ę"l��s�W�xC9���Ӈ	�!�R�t6�l$j��n�5�?�\bcX��R�(e%��d�u�1h/7��C��� �ƃ��+�z�qN�3w���^����Nyq���L#��'$T#v�ynJ��{\9�֭�S����sX�����|�w4�՛۽���l׷�9��[�jFc��*6�ӲUӱ2�C��Y�"���n�����gr���j����jZ��e�pŖ4Ǻqo�����#��;	3gN�KJ��Z�ͼ��(�b�ڸ�g����:T=�a=���@2��N�j׈��V�K���u���m�q8��)��C Nc�K�+�e.;u�:�ٹӠjb}4n�4Jı�k��L\�pS���y.��m�>�a#37&Coq���Y��(��φ$��2�O[�t�ˍ�,Xi�����	f9�@r!��`�!���u��ة���EZ]�T
�WF��:��Czd�WeOy���;8^�P-���,���Ggd��N�{�(�2��twEf�d��q9���������y)Eb�qŋdܪf���}�X���^fk��$zw�{5�<��]@�s��V��i���U/���{nm��a3s��^;�{�F_Y� �=���x�sT�/X2Y�!��Q��v��ڎ��m7��%Dn�04� �oe� �����|��B�]�I�[��;�a��Gv�3� ����ey�X�jPDN��I\�3N��c&%�
��=�%њ7���u �N�4L���̘��&��-��-
ot���gn�f�(86؜ 7�v��`��צ�}���9�Y���7/l#��s�o#�.�+����2�]F;ز����GM�
�ͬ鯡湉.�,�w=7�s�2���4�\�"��9%�t� X�t홥A��h/Jy6T՜���Y7 1�@����f�[>�&����&����+�,�ۅ�޺,���Ӝ�qE�+$`3�����4��FB�
oۣ��ͱ����tYǴMetFk:�.�S21���q�ݷ���;�{�t7W9;t��/����'��{��K�]S�u�oQ�Uiρ/���2(l]x��m��b�{�Μ7���b/|�:G�F+N������W�4y�z��a镋�줩F�`��\��w�W=0����窱#w&��W
��MW�sC3��f����/R+�����Q��E�Pۿo�i�x/H{7��v��:H77��l�i7��0��~��o�DY��(¦tes��R�9����3�y�e���]sk���qk�ůyM�5�d�W5����ĹϷ9�Wm"OE����xGa�wv��^�Z�h�D"�ę&��Y76ܹ�'^�r��L�G&
�k92��r�!<�9ϷZڭ��{u^G��6ˍ`�<�N{E�c&�V�s��n�}�O�,_��]�p�r�
�xiq]���J�ѧ����������y���7.<�� !1�_nD>�1إȜ�d���d8�[Kc�I�����r��o#u=Ӗ�xlZyH���)��'&&2���D����b���qs�.Væ�<��8����j�;�L�1tO�� \�۵n����wJ=;b۽hWU��ase|��R�Y�����
2���ށ�6�n=٧�GJ�� �in����b;��c��m��A���_>�մ���#�CP�8��Tn�Ԩb��\z7�Y�(��cN��
���{qZ�kԔ.J�`���-�!�lX�#b��賺��&�D{n����|��aO�8��H_^U�\���;�i��	 ̪k�Y���2Ӑ��J�ռ��J��	�2�p51��g�V��Q�yn��p?�!�r0��\��`��Vk"9(D�ջ�,�z�MR�1�P��k�F"իI�{�2��p��˿\oq(�X���+C��@��X�I��)q�n����;���8.�9x',�]�϶�!���)����e6MY9�4�}݂
�,���	�i3��7H�:8��"�^��7�۱Ud@�X6��������.7p=�C��Ӝ�U��;f�����8��/oiC����yU8�.;�t����c]�K�J�5���v�sޢ��N�����%wP�ba8,�ނ��S"Oc:�r�2c��#M��)u���o;58of�b�c�{�����TW�-:ֻ.<�LJ��� �O�3qtSn<��flNڬС���{�ݗD_qZ��e�k7�;5}܃U�k�)�ަ=�X��-�ћ麡���x��ڻr���=T��n�����̽��Á�b`����vv]]a{�x��}�$Nm#���sM�J�D���ZGP�6�|�t��xIN��I�{��W�H���v'x�bʙ)i�{��,��ҧ�-��9^Ź�ۧ��w�p4N��x;4n8@d&q�<�,��q�x�� �0�F�d���W
�Eˇe��Cy�ݺ�N�zp�Z�w'��bVr>��3l�&�vv4�����>�t���ǥ�"��ov��yB�*D2mo!u�y��&����ۚ�;6Eݡ�u������n�:��gW��y��a����q��iz��5~\�]�F�����.�سt��]�"����Rf��l���ap�E�m��뼪Y
�+y�h j�����B���kyC�uv�����ƻ�f+N�z���z��ߙ�͑�|1��ޗ�d�ՃM�������7�Ŭ��a����w!����]\ݼtQ/v1w4��}Q{(��{����>+|�ܱP�:�Le�s�So2[SL!�wݸ_�z�7 X۵m�l�wCv���@�۠ύ�a2p��BbPs8P�,��VP�!�^�#�;����WB8!SH�h���b9�cV�x�m�-@�a��/)]�iÏ�y�wo��\���\�ٕ sU�޼G`�Y�sK���aU��,�K��P�H�TQ�Qi��÷;��Tv��� |�U�.sɧgf��%��౻2�ώ��ӽ�m�Kp�-yN̡p����Y�v��T�=� ��0샕[E	/E����Q1���2�&낝�ǰ�\[�7.pߖ�Ow{�
��Κ{y��{U#���|�Q�}F�p��d'��BO�3;��4F�]Աw>y9����y�c/�m�6Z&��8p�f���qv��z� .&)�v(ɓz����^)�ʩ�Y3f��@ޜ�p����B�33�k�89�ssB*��U���A9�K9qcE�X̻����Y��:�b
1j�fv��p=��ʻ����(N䨥yA	9S��0	�����:�\B-9XPP�mӐok7,&T�F9�{�pv���'�څ�^��07/�::�,Ӗ�|E�;[F�D%�ۆ���XGnl�kzkJ��kՐbm��O-ZbC�L�(#9&nl-�A��wXq�&�E�j�rtݵĮ=�ɼV߀Vf�5�����v65XTyVMz@�	N(f7�+�2�z���s����(��G��0�f��N=3^�΁z`���Vv壚I�݄[Sw��ۣ �u�����A�p�pc<L�����a��ޤP��^�Dx�Z�=�4,��+Oz�|�졮C��q�Og.�nj�p�Ws�棦�/^�"�a�|���8�&�9���ᄡ�G0&�;{�k۸2��]�]�J8�8\t� ��܌N�����*F���>ӹt9�w{TS
Ã�Q��Yt=��:�S�L�Řz~yn�i��8\���܅���`s�;�9�wTfwM���G.އ7w����W�o$]v�79�nN���}y���&�r��/XOP�γ:�ӸF���1D�tY�!P5�5z�ן@3l��]�
W��?#����5� ҋ I���;�˽H��w^���'q�h�.o���Phw]n]=�%0�m�lѓx.ɐ'��!/t�.��Ѱ]8O`�d�a��Y���P�_Zη���tx��ރ7b��!�]Ŭaܙt*2���^�G�6�bŏ*~o���܏C�u7�� 7/i�[p�HQ�3�*���w"�̞Bܻ�ꏶ�Mۮ|ɷ��՝��1�9H��f�1����M�oA��z�p�Y�t�3�9U÷j'�Fs���'m�ޜwv,��\J-�C-ɮ\�p����1��xaĶ�R\��9�1<�N��"�l��#��7w���a[�\�Xzgu��WWk,=��|Qڧ,!�#���\�N�@����^�9�� �zv*�����*{�����o���l3�e�/
��7�>f�v�+Ex���q	�7nU_Y�gDL�;7Zg]Y���BZ�7	�O^�'�L=r ��-{���ٯx��;�Y~(#.J^2��+�!���݈�f�MZ#lm�7\N��m��U-�0V#NZ{ly]�b����y��d�D�[�[ˏ�{�:b��&�h&���q.ۂM:��� a�έZzt��� ÛQ���{z�Nc�X��}�Svc�nDgr};^I����ƥ��-o锭�N�G�:z�������5f�5s��`���ns��z�����i�|y�س�]n�'{�wi���^�n��]y�Yn�
��w�b�02Q,+��0���`X�ow�E�dmR����N�!�m����t\1Is�hR��č���7�|��{�L�k�zނ�<gL��U�ezŷ�������Cw�7&�Q�x��qg�Q�4�w9�I��e����t��������g�Sy��vv1&�G{@�G>Ҟ� ���,e��� �vӝ��!�4p/,r�)�^��Pш}���ó�p��+v8rl�b�$�um�Z#�n�1B9��Fwd)�^����^����4�h�8J7�^�:o+�y���^3��돏b;pmBG�kSyhDַ79�%Z梾�LeU������N^�G�k|��:�2h��BWLrQ��z{��&�%��u�;Y!T��v�gj�?k\;u��`���	�ˍL�.�+.�Ty�X�����s���Jû��4k��Z���Ox�QһcsɌdk�oiǌT0q�}M��׬�3�L!�K֧<:5�Ovl�a��}�
g��n*�^�m�l�')��ӳ����LQcW&��FwX��fp9�X�X)�B���Z�
���6�VK"LMת����դ��:����t0�nM�S�=ئ�<nUC�tvvɹ%LK�"���B�d���{�W��p�;�<�3�}���ZCmFlG7�B4=���v����ŋ5#.N<�i�3G��BЍk;Uќ����9��ͼ;fm}p(--��"�ۥr:6u��G8V�EZӮm�JUoE�p�z2��֑���+�B/X&[�ۇ�W� �-�]k�M�ݼi��Zú�q�tZ�>���u�A��}S�s�'s�nѽ�d���[Sׇ�Q����3.c��1�Y;"c�mm�����k�5�8db��լ�E�̌������Q��cT�'s��m��l�6q��͈1�Ou07�ڙ��h�� hݻw��mʝZyo��ܒ௖�5��V��ͼ�0;�{l-ΰ���\n�5�N���p�	Y�B'=���ae�D�	���߁��&�E�r��y�f�Z0�K���뽢Iګ�Pû�b�4iJ�hHrWF
&�V�.K�Ns��$n����t�>�.{��%4
�xb�}�歎)�z�۹�t�	S���LsM�4�:x-+h�Gk�L���[s�m�L�Gf��������ǧ�[;�n�Br�9���d%v�od�,��`t�G9��invt!�9�D��A>B���* ��q���}(J/p�I��qwa���g�c���rv/>��0o�^XGˋ+t"45bG@�ݟl\#�:�3��3=Nw�%��_y�j�y����2�צ�&�*��=�{�9��7����Ц�6t�\7x��0��ܞ��-�¼���o�2"���H�h�H����M��`64��v�	 �'&0�e�aM�	6�cE�.1�6 P��"�m�aM���v�`\`�)��P�&�!�(�]�C`��C
c(`�`��	4�q�v�����v�����&��M�N6.6L0l. ]�6\.�i6$)�l�0N�ӗc��)��ce`P�q��M��	�m���)�]�
��ce6�
 ���Sl�H(c� Sv��!�q���cl�L���l�N6'6]���?��w{�����g����+�����_��3J���Zo�V�TD��r�v��\p�w�1��%JZ���" ���#���א"�L9�=7��Y ���'J+�ǣq�|�S_1�;9q��J[
�����\��l3�
��9�u�yh֚�@��Ԋ���m�6M�sb����wv{�Q!�ٸ"�`�{3]���_���B=ZUH�{����m�� ��l�Ḷo�ص�EE���C�;��[��CA�-.���2Y��Ӷt���X��1��]���'�c�I�l�;<E�����n���·`���*G�8��O�媮i=��Ds�uE�"��8s����Y��Ƌ���th#��<���ɄG�^��$��<�%����;�$�꛶�v�+"^����|)�ݭ��\5]�e��a��1����ޗ���+�"m��%Q���yg8Ry�'�Y��;�^z"Y����b��N�:ּ��x=Ļ�������%���Ց6B?��~�V���8��[�]q�pؠ��sU���
Y���n��U���D�~�"q��^�!�w��N�����-¼<o�ۗ�����X1{Yj��3e�k��3���ri�n���_9^��aD";��B�!{��d �������F���w�w\؄�>�yoN��\tQ�ҫ���qD��;���������nˤ�烕c>�%���.^�ʗ_�5ry4$�|r�2]lTt}a����� .�I�rpMC���g{�@.��:P;�_��%��'Q�#������b^�		^��w�S����C���þ�g�zA�6��Vzy��t�wt�o�z��Fɾ��>�Oo�'�jp��}��m[�=ɓ,��C�T���=;���é����c���O���=���I�T(�0?M�� 잜8�v��R?x����=h?[/r��&vL�@{϶C�,�Og�z��(�׽�v�	�joöL#)Ly�Mg�W�*�w���~�}�?d?1��zc�+�����6eΗ{���y������a|�f���h����`ܓ���	�L���{�=09������H��"O�
;�����L��׻�����I��k[k�fﻮE��f聪}����qv�,�
:R���c�,a�P�ε{<<��\�2�D�6p֗����n��q׺Z��x���4,�Nr�~�Iפ9j��wa���{٫�l�uH*��\y0��K�?f�����[�_q����*��+��gmcӻ��n�ͯ���t��/\���)��߰([�/{���lj��zN���I�&8�({<<�;��h���lݸ���{�h5����<�v�So���+�K������Jw���sy�~��*2c���B�痴�}�X�y��-��u�m�����ٸ"p}�]��1�6�O�7����r=.oGڱ��V�|���8�$	��D�.l��ц/)����v䦄}����l롮~�h����I��[�;7�9<BMy�����P���\�/��p�a:�Zy�����jN�������g|.i�ዟ5n{ݹg޻9O@2(��Ify�'�0���c��d��K�hMۚ_g�U�}���l��j��s�>�����=����S�x�,���n{f?O>�0|s��r����z��.j�����y����] ��l�=s��]�k���l�/\%9|�F�ysȼi�H�:{j�w�۾��[�{�KC�o����9o�N4�n��H��.u���'xr�t�Y����FÊw���vx1T�������ū~�b�Q�c��>��Wy;Џ�x�űf������s�tǽ�-�QC���C#��X�)1�:'/�|�s�����,wN�QEn�gTȜ�2�均Ϸ<�3S^�r�^��P!��=�4��/3�#K����a�����Ǿ� ��W[��{7��q��}�'!��Q�w,�k�xƴ�|�8�	o~������T.Tz��ʓ;�+Q'��Xq|� L>޺T�[C�n<x�i��=�|�r��-��l׺�Y�g�>�ȷ�9��糽)6�׸j8��8���!��FhK�|�H�=޸J]�J��z�l��z�8�(s��8]�Ui���(�w����W���Y��=:|��/5��O�d
#G{�M���o�>V�;g�����oxz=�xv���K�%�zju��J�1Q����\ֺs9E˸h<��s��Kn�r�̓7GD�:���$yz�Yy4>��������:��c�4�J��/{�?}f_mg����&U�� ��dmՇ��j^�����l|�D	�Op�s�@�vQ0� *���>��~x=o��i��W����{�,���P���yOL����
�=T�]��z�{�W�=�!�ѳ��qwG�����ݴ֮z���8�ou8@�;����8��<��oU3x������S�o�����}�L�ۮ۱�ெ��x��(�盚ύx�j&t�h~��vT���;�g�/��R��L���t���K�Ӻ^G����y�P�c_���z�x����{�h�t��N��5�7��t{}���7��yz/M��M��M<g{o��)܂9�sï��a����l�&OK�}�S�@=l��3ۻ��淦��}��"ΒH���^|�$g^w��^�sH�{�<U��C�O-�C{N��Ѐ�՘7:��/��������~Z=�5dP��� uK#�T��{�c,����{Y��<���!�����R.�塎�v�F�ހg����fn�A׵LrX�o{�6���B�B>�njcG��4��e8.�ѧ�ā��%���/L���+�����2���p�tsE�-���+<&u��������7�[P��u���G�w���)wK�Ӟ.��1��0�����Ǆp���$�N�s}ʼիފ���j��K_ia��h	��}���y7��ANZ{�?w��1M�x,��{E�&���X���� Ҭ�o�>7�or�b��&`� ����3z��No���������� ~�;%�W�c��Gڀ�h��`ݽ����xz��1�w�ĞH�@
�y\�Ϛ�B���r.>�J��<p{�{(�B����f��g+YR.�5�������ٓ�Y7�V-l�9�\�{%�K({�W�L����s�!S훜�bA'�y�u�77�,�㱪�����e���h$��T�T�u[�{$��Ѡ�Ȓ�"��ۼ���;�f�{���|��>vR��ť��5���x3,n]ͭ�+/Yʊ����A:-�B2w>���*]�g��wxh]�Q��"'o�t/v���{s�F���}��֬�v��yFg)$�s��J�&�݌�����Zq,�}H5���z'O�zG9�a���bG��x���泝�IF�r�]�r��#�{Ĝ���pc��9��\۾ꢇ�=�yl�����;-}y�jX��_zו ���Q�}�x��W�u���n����������@{�=����c>�+3_�;{zo��Gv�gUǧ���Ӯn��7|#U"�����<q�����Ӫ����(ᛔu���!o��ҥ���K�f-Fؔ���d�V4/x����=tn�أ�]!�q����O����Lg�d��p�.���z�Cm#�����FCՖ���Q�%l���$���Ӫ�!�E�ɳ ���Am��ԣV�޾��"���N��l�Οg�\���͎���ȲY��=�^�j2�g���J=��za�{{����^��rK��.C#�2whjb��Ru��n��z>�nxm[�<CA�=�o/!:i�xݞ;�w����=���wϓ��U:�������qP�{�{w���w������I����j�����������ۉ�Ws��tY:y�d�����|�M�M̴>�n�����gS��&�Zss�W��v�l�2�z�H-\爽��K�Ȅ�c��\�8{n�^��N���;
�Q�g�D�׹��e�o���x2*#�mx�Z��`՜���׵��~����@,�cW�p�)n�k�}��y�A��s��fϻq�>2�PreV���a&_	�XޢFV��$�x����!�9(ֽ\���A}!��ږ�.v+��%�/H�:��snlgtKĜF�Ьs�>���q���^3��I�vs�^�����J��{#�����M���ʌoV�F�3�yW�/:s}��ǰ�{��NS�u�[�/v������C ��'<^�~��qZ'�>{�wN��Sn�q��b^?o;r�,����y�sپ~y5{ ���#c��0�^�wZs�_o��x���f����B�|!c�_X|������Ԋ�-��*S-���L[������<!_�����ܸrw��KfBw�!^�Vr:����n����{���^ŝ^{ҵ������ۂ{< Ÿ�\Zn۹��F[�������y�MB{�'����Ԃ7l�L��]Y=�F �����A�I9v�j=ܖz.�y�'YV�6́V�dР�K"�Jk»x���o��|3ݹ�n�q���5L�n��\���=���0��NR����o�	�G��^�8�Kǎ�e��j>
���<�3\��Q��h�<"��s-֞�_���O��r�M�K�''�r����c��hOw��^X�_�<i����G!=�W����;��ʿ}�1\o8(8G�4��<`�[���:w�>��x�z���3�S�ٶ�>�&z�����pn�9Q�̙d�N���<|�=�P����=|�{�[��G�9�(t����u��ǟ��OI-�r�x��rU����ˮ>�gg���Ba�s~H��Gp�пc+;���w�l�i�nRZ�yh�LG{G��qΘJ]l�zѥ��	�XJa��݅	�Ƿ�_b6��»#�ދ�{����=�(����f��w�s�>\|�]����!�U���6��qй5YOw�vhL�w�'m�����׍��x�5r�zyl�n�KZ���ׇ��t���S�3�,'���!ۓ9W^���(�N����}*����->\*�돾G&Ө�p�o4��<��>��|7=��^��<�Vk�+��o����#>~>MY8v/V�ξڵ�����r�-<3Ɓ� з�V��p�{���nt<��_�x�^�|m��6���Y�72�3V��.y��XVwhY���p<����!}�z��;Z�?�3������[�Moiܺ����b���E�.�SeM�x��6/��1�z�Nvz8gQ�x��TS�=dk��k��|<�ɨ�к���>N��&k�r����oܶ����Y�y���9�{��O�t��2M��9m�h�(�<��A�q-��������a]w���@`\Fy�o��xsA�4秡���<��7u��t;���'L���]��A��臒~ڞ����^���.z��8�劼�f���Q��['��&n��lY�n�6�ve��ޓ��GI��G=�M���>~y�h��{zKT�wS��՜:yD�0�#�#Yx{|��[�]��E�O���8��w�K���zsS���vα�1{G����c����΁��H����Q��w&�㇃��Hm	a6캩��s�`��{�{w���]��7�0��A�{r3{݃.y��6Ff�ݸNnz=������}!�����hS<�Gs�ӭ���4���(�|9���O���kpw�Z1=����o�v���Ww���m�*���gu�y�X$�gZc����������;F����h���aJ�XIsw��9{c�������]�y��r׫pn�����x�7���A�;ss|��:�ߕ��]�@uyA�N`ٹw��]>���<(O�q�u2z/z�"��!�hq,s�u���=s��/�^�Ϫ~l�K��=Lh����1�ӢI���w���g�<����w���Z�.c��K�38�(�q�xI�ҕ�0��"��xg�Zl��_���r�����a��ñ�}�,�޳�=�|�y����sM�s�>E�ط�5�Q㪠�����s͏`�%���X�&-�+������^������l�e�{�j��<W�i��v�b�qA�o���������=W���\\���ݹ�ﭘO`sͿvl�m��}�e'���L
��㔛ۍ�g��Xrg���Wsݻ�h�=�𧦛��ih�=���qo%�${��}�����5P��6w��w՞�X�}��b��'"mO7r�/i�0���7ۗ�z�}���Ƿ��{��eމ�)Y�a�ͬ�ю�ǫ�a2墾�%���z�?��f���M�w�`��rƛ��f&�x�^�N��L���+�V0�X�H�=�s������۝��J��.�׻;{�G��>:����^����\���7��RWz�͔����=�yf�h;�����vwN��4!Ö7o:gѽ�K��/8iʧ��X���.l�O��窱�=�&b�>�����i��m� ��4@}��q.��;2�x�������(��ET���7闅�jw�ڶj'��5ǝ�/��A'�M_nAw�
H{�Z@<����0��}�ބ���x*D��7�ӓ���=�%�N�w��5/\s�:�wtẵ}-GI�х*g
��`���z;�%踖��q>�����lS�̤���p��=3W�S�q��<��aY�ьn7v��J��*~�6Ӯ�u�=��k�X����G�y����grL��Ӧ��f
��緎.���^��Q%�>�n�#���+��Mg�KYԷ��<{�U���Ǣ�{)����k��\W��w�Wr��WGI��%����P��^~S����1�{1j��.��9��7v��f����،�ݲ:p	&�>�6�{IBn�3wb��W=�+G���aI/\�y٭�s �ww����\�u��7�(���Ĩr���㧹\'���=������g��YQ{ʫ�f�}���m����C���m�>Ȯ�Y�0b!y����X�eJ]���ઈ���=�/o�WoC�����}���ȥ��|7}^��|�|��������p7�rF��㲷\=A�TrS��G)]+춋���#&�]��k��b��"�5en�z�ǷJ�&�=�v�m�W�l0T=�ά7Q��	�*����7\aݳ��0���8��y�O\��U�%պգkW5�v��[���<��]�[v���zѼ]�Ƅ��:�N)-E���#��Eۃ�C���닳�Ol���9y�^�s�n�� 8�2Y뇞��z����[ϫ��n�ΰlMm{a�]�۲>N�	gE��9�r��	z�V��2+ay�y�y��{�]ix�˻k[q�L�m�
b]q��7Tp��m;�7S�v�]��j4���`�uc���!g��R+��:�9�j����E�w<j���1�v9�{mi�`���|�o`������w��mv�­��.{��fv�{]ʛ��iqVM����	���8����mۇ�s�p��/`8�\s��s����"���9�dv��y��Ǉv�.�8�.'�fŦ×�t�l���'�-��˞�Y���On���yxoY�FN$����^�\� �e4'`m�u�rn٤'ou�7���(Ȟ�;pu�T��m�4����n�J��ų��[��n��x9]��Ll���h�\v�t{DW[��۠v:v�G���v�g]�q�i�@+�rh��[���M���ع���;�2<`���xe�y�[���	�6�w�c��G�:�]R㶫u�r:6�N���ni;M؜v��ݺ�gg���:�� ��vضM�/V.ƹ���c��;��`��N�#=e`�C�e�u����JM �I\4Gj�wm�=��=�2�Z�^3�υ8����Gg����(=�v0�.9w^��t(F�ܯg7D��mv5�7<΍�D���p.�r�7GX�;`���d7^���*��n�ŹŎ(s��ˎgGtp�Q�8r�v8��!����v$akO"��g����Xm�ۛb�����m���ݱ<�t��Mы���v���8N�'6;u��$�����vcsm�c��M�nn�Z�Mۂ���vKF,�z�7����9ur@����Q���'�c�"{m��>x�!�2����̩EPb'��T壱�㓶��>�����8�:xɗ�	�ڹ+��ƚ�m4�-����k=�G�va�wk���z�=��^0�����Q�N1���ۊx����x��p݀�z���w�����ݼ�\�vyLgOl��+�v˟#�Y8�4�&��vx��&.sg\eᛶU������%�<�����l�,�{jʾ"�eۊ��_7J�<W�\��mÑ�c��68�Gv�=;�3�q=k�Dv��v9� r�Ӷ{���M����{v޶�<�;]X�������-��JN����Oi5�Q�Q��[γ����y����D	79���n���,u��q���A����G�����n <���Gk��źsu�6�ؘ�t��v�ӡ��kn��j6!��]�ݻ>�={����X%��v鞷�w=���pr׷�r�e`r�8^��%3�c[u�\s/O��9�{q�n�k��Ѻ굦y��1OGN�bB�9��ː�yKQ>,v�μ��c�9�v�٨̦��Ɯ�v��ێ�Bsr*vz��K�q�v2{'G��D��7:Bν��Pv�F�w1^�6Ϯ�ܖr�s��Tn����{1e�M��{��ݸl�����Cf���u�u�[�u���Y68˷m� Sdf|�k(�I�ֶ�l��'�q\�͝���2)�c��e:n�Hz���:�\i�s�iݻ.{u�w9֞�p��7�a�֗�v�3�S��#�;rj���;��޳���u�qnw����7F{LU:�ͳ�9-E7�����i�����{v�y�WL�VK����0��Z��/t�z�i�����\]rt����5�9��8�v:Jz���=7h�p�C�pP�u6��5b���g7X�ڰq�O�=v�ĳWd���S�\�v��Z�;]BA>���8�#9�Zw[����n8�n��ѽ%�����J����E���]b�E��`Q�.�g���ɀ�a��j����W��8�>�<f��rql�.��һpm����7b��ly���`�3Ԣ����Հ�gml�
M�E;Wm����dCn�����f;s�&�Ǜ��n]�>��<Q�uJm�kU���l�q����ϭ��v���<q��,�)�kϮN��Ӯ�;�c��x��s<��JB�#�v���`}�3�v�lՈݛۧ�e���\�[=����Z^׎��u�[��X#���;�mŭj8��[�]��f���؜;�񗇰��`�Їmh�A��֜��n���u`�w9Hn�j6��F�u�;]uS�6�]�n��tr/l�l=�;�Q7/��:޹ɞtK�[���sgk��\O+���B:�D��Oٓ��vu��az�n[��m8�Oos��n�܎����z��'Vpn:�97vy�.y�b;)v�Ssc�{��ӳ[^��S�z^�K����7Q�<��<�Fù��;{8�,u:�Q�M½���V��i�ՉZ��k:]��:���-����,\���t97n�1��ˍ�-=+���]mӋ��wn��u,�u��t�[�5�j�:��Z�wl���O;bʛ�h��}7�]�U힖ݹ�dp��+���G;X4�O�y{m,u�;�C�N:z��;���Y�V�BWnr�r����r��uI�����ݮz�5�x�d�H�jn�n��'z�%V��.o%.t�8!�g���ls��M]��ӰqӉ5mq���%���fAɳ�d�j��͐����m�v7��C��g������v�!t��YD0��N<s��X��xeY��|<��|k�����}�N<,���m2�&�l��湊n�s�-gO��s���WT�[v��6�rk���Z����mZ�tM�kz�������55K3�Y���qL!�77F�yӵ�ۮ�-��� svm��z�����T`�z��<]n�����\{lu`�+�S�/"m�s��سƞ���r:���..���Ն���l�{9�ld�7�7�ę;@��K����r.�ݹ�ݷn�ns��ɨ���Uz�]\v-�ڄ���^83%�{n��F�3��O�㑸�s�y�Fl��aË�i-��v�F��q�j����I�m.z:�Ɲ���z�h�1c�C�]���v�l�8]�'���[�b�f�]��<�n�֥qv�q��3�]k3��9�8�Lg�{���B��㡛�	z0�^��q�h���[�lf͝�v��u�h�/1�@�Jn�ݖ7P��;�)�&R(룳�tt�m��(=%��V���y麷��f��>��]k6�ut��:c��vKg��;�s5屜tO])�e�6�M^�n̠�s��P��Z�m��B��\����<۳�y��������3��/S��s۝]�;'m�:;L]<G1�(��8�%�v8��l����t��=��Իc��7�l�F��]�A�ҽ�S��6uюT��0�[:��ܰ�n�4���jr�;�dOA[m��!��^3�@���������K�p��wSc;\�L��Jۣ��mw<D���N��M�g�c��6C����u��9m������f��;�x9�ۅ���=�F:ϻa�:r7n�������*k\�of�l�֣��3mp��؉��rXk�ι���Uɓ��s<��ȹv/n}/l�۳�v���d+ �=p.ϝUz��Xn`8x�s=ί8v�x�Ď7]��2��n0vݞ����M�h�t�fSu��[u�ob:ݓ<�BAۃ�K��xyzN&��;���0���u"i���U�Vqư��[����az�n�$�pE��)Z���R���[�.�ۚ��ꥹa�v�y�Ħ۲�U��v���9�컜Uʁ�'���T`:{N���:�D��,f�16�GN�&92��	q9���i��$E�i[�nm������k����ql۬���b���nY����e�6��v�us�g��b�pu�rی��gI"(B��mҋ������p�a.m6��t=nu���Nv�Z;]�,.H�<�]8��ݜ�:���6/9y׻%�Uu�o�,uv��M�N��n���pa{�ƻ�K�mG;#ݺ�q�n=ץ����ɔ��X�X�N5��ڮ�v���űg��`on9jۓأvKI'G9K8M�X�S��۬��|ݱA����&�k�v�#���10F3�&��.�rj��8�.h���� q��"��m�i���8m�v�N��e���hqsk/A���zx69�s�P�]tp�u����W)Ɠy���z�h7*���]�5b���ݨ�<�<.�Inۚ��N���G�����=ָ䨺w'hv����·;SLn�|fp�����6��A�ݜݞ���x^1v�����q�My1�ӎg�c��:郰�]�܉��[a�O�0�Itgs����a�|;����n�sF�K�v�]v�.���vCa�9�suأ8�v�6�4rO��:�$]M��p��N�E�W�nɦv��p���g�Ӳq��t��8�۷&N}{cv�uٱ[[rJlS��=������u���r��^\�\aөr�i>O�,T�B��欔=<X�OUu:�WY�ג���gQ��Q���L��.�Q���#�;"3��n"{i5�FW�{��v��׊w��9Y��m���x�8�[�vaܯ�tN�����M��i���u��c��y�V���Q��S�<�GYz�x�<M�`�����͘�6����:H���Q�-�j���e����wn���=w��l?Q9UG&DE\J�~�c��G�U�5�\�fTG(�* ��C�/Y`s�W��I�!E�4L�2=�F�E�s�qAdE��J�­�x�\�
*(��	4�J����&DTG"������I".�H��DpԨ��䆨��¹"|�@��Ĕu��C�*"��Q)�Z�r(��Q��L�g.DQDgI�M�i�H**�,���Qe*"���L̈�A�eP���9�dpN%E]��;�a%TU���s���D\��:Q��Z����j&q
�3"C��9Vj�U�DqD(((.U��ʢ��3�(Ix��Ap� ��'�.��9f�r�*Ԩ�/2'$��VE˨�VM"�"#��9F�$fY�H���)^�Bf�(ʹ|��~���~~|ϸW�m;��[51���x��M����t��z��mZ��`�x��g�-�8�k3ۋ��k熗8nkR���a�'c8�>@}�ݸ�:�4�:���s{����5������7ύ˝��=���l��s�6��9��j�%Y����̮�-з�"������G&N�
��= x�FϮY���S<Tl-�c�&K���sc\�l�Y��J����C��vݵ`�v;��nCEc��[mX������n��>�[�����]uO"�,,��X��:K��Uϓ��;��g��nom��[z����-'<n�率v��Bv��kX���y��֋�z��E�;q�*V[om��.�� wϝ�G�8g]�f�}85�`^�<kr]�t����w���v�ʍ�M�t��vu�e��z9�ۛ��D�;ֆÔ��d7k�q��=��#^㫲�0z;=��O �P�n:K�ݗ�[�Ɨ$m[^8��[�!@�zz�|�����q��j�Fwk��H[�tk��xWlkc��N�٭�U�ظ�;`w*wK���vS�Z>ξs�Ka���V{f..$�^��8���u�1<�g�v�gmνr9��C�l��$�z����F�0�ck��#u�|�h�u���n	�9�������H1m�L�hk�E����	YM��;f����[S۞@�5cSOo���s�d;n��dpv�u:�mA�x�&Jb�e���#:Sf^�7`�Vw2|����v^M�źms�Y��<�9&�Z�n�=��m�۩��<��[���q��3���:�m�[�p�D�:��6&yW�1�<���C�����21�l�(t�ں7Y!��^[�n�..Z5n�k]	�6k\�`��6�1�&��*��y8}�vۖ�,���s��V��7c�2�2�u)�]����,1Sm,e�f�RL/A�E���+�N��Xp����^m��<�]�I5��7$�wvbl�"Q�MW*�!ɷcy��ܘv�<���^���c�����tt�*<="Ŧx�I:��\]
U7U��Lv��q��Cm�.���^p>>6NN�m��Qn�NwK�{�GWET��s��<:::�q�y�8As��AA�q7�����Y^]�@���p��Ã����[������V! �O�^\	�\;�t�kM���2���w���ɍ�C°�2`���CV�ݪ�L�t�"`Q$�F���$����I�9:�(�H#���L�d;ô@v��lNP�	�/��,	,%C���Z��~"��܉ć��2q�0�"��6b��)�6��r&�$I� ��Q�I ���6\A�ݓXH�6]=э�xZi����h5��F`�g�cM��V6�>�U2	�=��$����b��LK3�S�y�����A��v���G<=��2���Ӵ0������ҁ!��m���؂��Ö��VNϤ�׏�H�[x�
����p�┩�-UD������/�@27�o��7�������cV�e#�Bq��ǌ�QQH>fZ�fo�v2�j,viDdάhd%w/)YHf2l�V')����3��k�h��e�z��I|�	���$�v�ϧ��>l�������h�޿�ce� Z0t��bO���&qHmgE�b����+�:����R��#3xv�����;+1b�4�@�ʰ��b1�S� ���Akjh�h�ܑ����'ӹd�k6a�D �HdEH�H$�R%�>M������bL��a�["I�`Z��,M3)��ª(��_ � x D�2�;/v��[�z�w<)�F��uu�+q�������$��I�t�|3�AX�=$n�H�u2wglf�'������?t��3��6
D��8��
�P}��vˌ}aXcKV,�$��ځ&����e�C�g�`�i)��Ah��|��$�A�ʑ$��4kº���|=y."2��A�[����O4��'^G��A���6��x����{��?��%;�[�3���
����ݽ �m+�H#wjfj� �R"�h�v�R�~?�р|��ۀa"�j$�A =li˚zʼ� �{�	��2���;�gh 쬉�^��C;��ݪ�Qj��	7�S��YdV~��eڲ?�- "0�����cM�w����S�tn�.�Žv��}�|̙�O�������뫛�lۅ3���ʟI �[g��alƙ��t����?~�n�n���e����n�}�#�g"���&����U(��r�|O���x�*9��F�:H����)^4�cr`��7FW�������j��*vha$f]@�K��2 �tr�`��dj����;�����u���R$��	�ڟA�!�وL#�i>�Ø��T%$^�ɃB��WL�^}�=���s��n���ܨ��������,j�
��ǧ8?_Ә�\ߴ}���LL�,E�ѐt��Cw2�Ivǂʑ�V4���$��̂I���$v��O��ұ���f~�����{��V�N�'N�8u�jc��e�z,X��
n�}��w�}{��Ur�H>��������ځ s9Z��k�S���fn ��h�炊�X��x���2$MVK	������H%�nD��v��I>9L�ŏ�B�f��u��њ�u6�d��3�`��>K��YH���/w�W�I��	�v�F��b~�$�[e<8���~�{�+���k�>`ח�$�N�ԉ��A#z��~̠fy����T.�_Če45��{�S!Bu��6�8̚�iܺ� ǘ�QLN^�HM�]��0++�Re���l^�f� �eL������n�S�@O�gY�#"	������_��w��ߤ��/���4ZGG
�眊�eM��=xQݱg�;���uyড়NV/>g��ȀRTagv�-"l.��/g����u���={�ۜFڶE˞��ٸ��]��P���	��
Z:6q�����d���keS���*�^x��fGhX����Q�9�j�v�ɴ�oC��v0�s�n8ȉ܊wR��uۂ�Nnz���!v�%b�u�o����=;���蛮�����"��[=��B5m]��т=����߼ù���ô��,��Ky��yP'ĒN2���w;�ȐI;[R$dn�Sm�D"�Ÿ�^���������لA9{P$x�O�n��@)�ȋثM<�r�����T�6��~���� ��S$6���ܦgg���	�ʑ$| ���{��~m��	�L��8�i�۬�m��JC�� ��S$Y�jh�JSmJ�'k#$H%�Z�`��l�'&��h�0+=��'[$njz�;9��'�U��Y�$+L���>{�����D i��$;<�;��`��0D��fݻw2l[r�8��__��b�xb!��]@�O�3�'���	�j�{9��KU�	�S� ��R$��6^�@X�,� �?<߄���)��o뎤��)ۍA�S��&�zp4&v��v�w�SY��^���%��N&�;��H��iSUp���Fk�4�YG��iŭL+�K�\ �M_)�@$:ޟH8����3d�Ϯ{ �Ge��m<XPE�߇�s7����јT�VɆ�H$�Z� �|�vD�O�dc�v0 C�%��2&��dI�'6.D�A/ur$@'v�Cք6��<�@��{u���,��4�1���@;YP$�)��z�,lLÒ37fA �Us���u"A�
T��������0��+�)�ٝmq�Ou��p��O`��l�Sn�vܷY�����_���d�P������ ��ȟ	�9��H\e�����}��{�����,2�$c)��~��$����P��C������_odH�읹F9u�ٶ#Kf�3X$[ô�ᜡS;H$��@�H!��ɽ4����0�3e��9m�f�il<4.zYZ���M[0G��н;:���;x��K��v��gi�ӵ^ٟ���+�1 �[3�����9v��㲫L��][L-�t[�\��>1��c�ȟI����5ʆ���z&]��S��CǍ<I������k��a�n�d��X�I�͑ �	��ٷ�����v�7~l'�Sڻ.)����n��Uύ	չ�sٻl�n�-�F��W������&b�!�6�\��[H$�ݙ�^�E����O��D[ʹ�	Ur'Ā��gm�������˛���|��`�SA���H:	ݙ��>�A椋Ͻ����y����Xm$c)���zD�	�ətу*��f'Ăm]ȒA ݙHEhB�×-�����0"��h��� ���A �j�f@>�݊�zJt�	3݇u`�4Ļ��86�0b���㥒7�������?{N����S��E	9m�9���%;]U���p޵2lM8di>X�D���s�-��x���ŋw�@����g�z�V]�k�C�)	$��̂H Tn�l2��Z�?X�n"c��#�q���L�<{V�	xnCl.��y#u��dњVݞ~������������L�>�ə ��Q�FDb�X�N�y�׵eȐ	"��D��8�ƙ�>��J�_��zm���MnLI ��ؐH̭̓Z�Pd�L�Dě	0q9>�M� `��{t|�n]��ʌ���f�2�"�Y��ϧ 9����3'�n���G	ؘ����'E9�����cTI �QWH'ڶ�:��)=��`v'dI �	��|�,��h�v�1�?K�WdJ�m>���{��A9��IV����-�}׈�x��X�<:dV9��4D�i�~�>�k�~ڍ�W�ý�Ot�N��rC��L��2x����Q��复CW 4��e��`�@[m�e+�9���7^s��pQy�l��ܽxws��u�1��fV����n]���Q��|ח����qiu��v���#іw*v��8�r����9��c��q���<�aٸ�v���j�T��61�7��a��x�� ݎ�gM�s�r�n��G;�(�r� Lm֞5�p�)�*��-\�!���ܶF���Tpvnr�̯����7N�s��g�6�I�F�h�Ke;�츽���a@'��]=�h��o��I'ض�O��X>��8ђ�U^G���Z@��)B�Cǅ2ql���h��m�e]�A���I#V܉!��.�LEl?���������Gx�8�x�ob"܏O�6g6K�D*��jm��N����(&�LOx~��M^w]�a2xl�pG��*��IwUj���~�|��it��K8`���y�@���ۣ7�U˱%'�i$�Yr$	w���4���Hg��b/��&�42�r&����LmȘgm�C�t� v�k��=�?Ͽ����h.�;CCA�q�K�~o6Td	 �Ừd8��J�z��a@ڭ�&p�k"�8w%�8m��>;���5�`;���o�!D���}=�����΢N�/�	3�5�	�ʣ�&�-��V�щ%�;��/��7�(J�Ny1�<��Y���rf�-�5�V\	$��S��45s�M��7��~}�M��
�ɱD�A�� I ���Y��6q�I��\��$��ꉘ�&�� �2>�hm�NЋ����L��	 �Iz�|I>���W��a�٥��ZC<ջ>f��C9x������2A �[��ѳ��zH{ʑ �	9w'� �E�Ɛ�C����3����@�B�\)vs��y-÷��m�.M���mi.2�j������GcH�v�܉ �{�"I �k����E�N�=��Ϫ�$O�'Ʒf$M���o]�v�v���O���l��kڊ��00���댍"N�X��y�G��
$\�c�D;<��U�'�dk�A����{=��������n���N���sэ�	����N��F6��t�T����xK1�r�966��-�{s�����s���۲ͺ���rg�R����{�x4A/Q�R�}J��xo�����'�{۹Ǫ�.��k#<���pW���)�����>���Pԑ��4�rї���x��N�O=�� �����Q�M}���^=�9��z���B�ܘ���X�u7���]����D���J֍�垌�]��q�n.������`_;ϻ��t���2����a��|��|8o����<.�Ϸ=����qx��NQ�e��}��1��$<��������{c��}q8ϗ�.��d�#���!Cz�ȡ�����+@�6h�sj[��|�k�1�Nz�:�������}||���s�P���7;�q�]�����x���+���t�|��m�5_v|#���x��/t�ç�2m"���?3���>;MO�M��Tؐ�oS����u����-8.��b����n9�yv�{���A�{DN�}�zp.���㚷}98������\c�s��}�ELj�wuC�O0\��;�7���hEO n��L�پ/�7������\;/\�ߡ�/��zx��j����77�k=�ó7�S�x�n�گr�O*�,t�h gw�r�cD����"3�M}����3�y�]��o�������+@��!��W����>�p���>����5A;OB�|���4�H�͘��]/�sH���L����>�0�K#��dAT*�s�%�IgL���T"�J�¦kU�%˔G��PUW*s�I�6��'�'L:AH��#0.��4B��!*eI�C;���
�%���UD���eEEs��Z]���i��HB9Dp������#�N�����(�KΦ�*�7���u
L�:@�TX�˕��#�Q�h�\ �fZ%TE��C�&E9�"P�E�j%'J
/%�QN��Bap��=�w�(���-b\$�	�����TZ�q�:��B��r����U �$�NG�۳DrTa��Yt�8Qy�-D��/;^u0���R
"�T��S�]hfEeQTr�E�+������TMɥ�Uʪ��\#�� U��wACI��NKV;�G�d�^y��Y���s��|q���߇ͅ1������������.?>y��Ӱ�j�p�8���(� ��RO���k6;���� 9� by�So�;z�;N������&�q8'�7��}�I��b�]`0�;�ݼ�@���b��{>O�y��F����ϓ����>�c��b��Q�~��~|O�	�������7"�|ޛQ���@��;��:������N��	<��I>�y����k��f>�=���`��mē�J����Eϳ��.-�Z���oJO���5�~w��s��7M�o���۽�yğ_���=v�'k!8�������;�I�S�_ߟ>)�FL~_^��_�����aK��8?Om��\|�����	 �y��zQܾ,������}d��$� c�  (P/uo~�#�w�}goP��iſ>}����o\N�'�@�[�d�y��� ��u��������e��	>�gw�����U��g>�����G��V�c������}<��G��>��������Y��t�_?�=�e]�!�B#�]�I�Dy��{hkc!���w%�!�M�q'�Ϯ�C����~w�~;������7ӧ$�)����ϟǬ�.��a�Ώ��<|�ˡh��%M������xĶbO����uq����^/]��r��'Ȅ3!L�׍$T̶��3�"(��U�5,� ���7�	����������pI>��k��"��Ǿ��>���ϯ�=w��@��>��t|���wYOh�����}��dw�_���g!�����o��Ǒ3��t�d�Z%�!H����v۞3��p��1u�P>�ۓ�.����On1v���~��9{�|�������ǜw��>cѝ��L��������LN�K����\��1�n��"�����u�  �oR�P�����&������a@��/����C�`�#ȏX>G��D|��&Ͻ�s�.1�@c�Ϫg�������pI&?~����c�ɈgaO�����^M�[�x1�ÓF�\��ӻ�<H������N��f����Ͽ����	�P����?{����'iĚq�_?�<�<�������o�k8�~���|v�Bv����oT������;��1��üDxP,|-WL�^��0�8e��}���fa���q%�ŲbHpI���}X=OG�t&}R<H�OJ��������� I]Y�"<������P�w�%������z�O?���=�=v�	�Bq�������t����G����������N������S�bgb�����`��aa0b� E��G���#���uq�n�L�[ӻy
)љz��\͜��3Vّ+b&�����zg��n.G�)�U�a����f�7����*}ѧX+�y�>���_yWu(��Q:�h�S�D��m�f�6�j�.���r��8�g��kr�#��v�z⇊�ݸn��;q�[�������:������4��{]�GRf��\����#�v�V����Ƶ�<ZڼnM�4L��(f Yݍ�)�t�q�·K(r��/f:��y[����N�ӣ;��gc�q��=��wnϭ���a��^oR'1��5�f�I���Sh�`�"!��'l��m[�[ub� wQ�>�<�� �<<:��ͧ�f�K�/>H��~y��~.�@� HN�}߿V��|��||�{�<�>G�)��/eӊY�gޓ���$�Ȁ�������M�$��sb0���1Bb<c���2<O�7�*�+���Z�����L��&'aK��>���	�Fw)$��1���x�`�9tw�rO��<���dck9l^<(zɾ�~�_>��q봄�N<���������`C H$x6�{g�CĺY�c��Ŋ>��ϫ��av<�����aO{�����p��y�{�H^ ��$���+�CM\[*��A!;I��}�Ǩ.��\Bi�����Cď/���������$�׻�噷���>�>�8!$������=LGϿ�wb�O��>�'��tφ�������۳$��Ǚ�Mt��8��NpIc�����	�@�'�ߟ��2����(I�~��{�q�M8����}��9z�},<L���*�bĢUF��붼�1�� A#yj��xdg������������7�w�ܽ��o8�����G����y������8$�I1?~��$x"�xt��ꮒ�Q%c?6��� �?~�?,���	�ǟ��>O\Y���g	c��<�
"�@�)'Ȁ����u�B;�:(�U4g��`T��(U�x/�W��7����^�����q�0x�I�>����w׍��^^�0
BHҷ^��c�	�R�����������밸�N<������op�M8c�0>��RO���������y��o{��R�D�y�C��"��
3��������El)��_��>/�bM�}�H�~����n]f2���m���;��y�����(z;HY�BM����ߋ�ri�y��7�����Q�zo��NG[u0F�-%�͡:ꈝ��h ����ϯ�7�v�$�)������T�Cŏ�	��a��M�/����M��rbd=�������$w����������@�������D	�P�����o$
���r^N����P#�|/�����)�q;�;�����Õ�1�C��M� B#� m��jsGO��sב�;����,a-[�&�񋞸��:Q�m�:Y>~~w����������w�g~�|��Fv*رF>~������>�'���~���|^���7�~�l�� a� FN�#Ā�}� 1���	��}�O��5�;43<Y�xzz�8��������av�{�����C���ߟ��ԓ�����c�ɉ��	���O�	��1�Rc%�j���L��E3ŭƒ�1/�y�E���~.� N�Bv������p}�@oy��	 f�aGN;J��=xN'�o��/���o�ͭ�%xǆ����s݊E�H�Y�I��/�!e��o?o���|�w�g�g����.�����]�B@���$Gsu7��B#���lD�y�C��!1>�s>�g���	�3�	���a�����ϋ�i�Ȥ��ߟ���`">�������G�.-�.�������&��������
b���0"����(�1i��>�'�`|3�|��S�H�Q}�>�ϧ�&/~����1�Ɉgb(������l,��w矿���U�n����\%�E	����AMN|��w��n�G ��E+�%ͻv�1q�)�����s��<�����?�>��}������'�￾os��NӈM8�����Mɽ>G�z��"1�FN���/]���`}5��.��'apBI������z��~�3�h�x���
�c�i�'�x���3{®%��-�N�N`��S$�X�N	/���φ=Os�t�:�����=}� 1������M3=/C�/Y$��N-������<�ů'�=7���$�����z��'!��������z�0!��y�C��=p�N{Gs]ޒ=�L3�Q�����w���bd.����o��pI�?[�ş'��o������S]�׷���e�{2հ�"}�v� �n�Q���e�W��/�/�{1�O=�V<��ٔ<�i��xE�]
pT�J�6L6d8,Y=�/M���e��ʨ/�J�63,y���fG����sH&:]2�U|"�&����;�m0A~��i��\�Yw9�}������ �{��3����^L�����k).z�,@�o�s�t��^.!�]K�C����v�Pvx�Js�v�M*��+�^��SJ��5�Po^[� )�e� �u��%�Z9΁2�;�����3x��)%�Q���DQ#�����	�� ��s߹no�B�����!�u��qVs8�@퍙��A3_�p����<;Ë�a9��	�����$�br���޾���1e��>�R��ܻh"!�v�L�²AQ4�QI�
�v򳾃N=���+�|��� �|�I��7y����YS��+1��%������H�(U7�"o[M� oy���>���|}8��/ۮ�=�i��F�5��n��q�-L�WJ���D�y�F�Bd�`��yWb^�F�ֈ���Z�U)��}7��(�@{��t�ɚs�j����1�ۘp����Á��u��9�GjYn��9��wg�t�ݝv1��*��YT�4��ݶ5��ۧ��b5 e��'�z��]xnx� � 3ɰ��K��`1,n9.�̝ƻW����v1=�����{7�{�ϷRh&Z�Σ�=7&���2��5���l8R�v�^۟9@6�NJ�m������������e����dI���;I�:z�Fb�9#�yWh�`�@su��0ݛ��v�Kg�G]�὞��UAS�G���sL�=�Zi�b[���$�/33"c�p�6��-B�w)��t�H�GQ
iMT)��׶�02VK���n�~V  H}������i�DE�����k���p2ӟD��*�Uv������79���,�������{�⫝̸{Z�~�� ���i���2�4|h�����v.�
��_��$y�n/&`���ղ$�VC�'���=#UC�E_6�a�Z�� �SJLM'M ��m�>���mQ�E���4�f�m�(
��M�F{�i�@��fܰ�<��U?��������z�eF��	x��>�B���0�c.�U�:pZ���l�:+n�_�_��?7~��R�S}��v�� ���[P��n��U���G.��o�]l�x�i2"�皸��)yW�(*b�����P K��P�����J��X�5BVɪ|��&գl��=�bq��^�-��ìA�`|3����G�q����9�#s�)�O�R��1�-�����+���74a 5�b	3c��N�11t��u�������Q�#��4���q����z��j�Cε�r\]�Ҋ�W��! w��W�yT��t��r�"E*U@*���|Gk���V������|�	�{{�@�s��}���LLFϸ��t��d�~"��M&_����)��&jJ������"/ۖ�L�G+�������� .q�M� ���_7Zi2�U��������j�PpU�C��v��/���'H����/iv��n��[S[��x��TI4��w;n N���|�i�u�=���w�qv���u�� N�k ����D�JS�y��<'H/& 5�m���.�T�( ��Zȇ��֮!��s{��H�}�M����7~��҈�AS�Z9�W�|����6��2 ��8n��>�/Ci�C�\Ƶ��j*�[�O�$K���G5�|���"u���0��`�o��Ē&��l<�y*�}�;����\F�'�ZƀA���&<0�DAx�*�3u�����w��g��G6��R^�Zq ��kW-g;��Z�f|zC��l`/�K��H�O�B�l�wZ��{y����kZ�e1ٴOy�c/31e�u��$��ͼ���'�c��,�)Α��+;;n��gccX��� ,����4�;\{\�N�&B`^�#*��}5%J��{�����e�� �[�Zm�=�l����s��� {���Z�eG�QQUQ$ҧm`g�9�r&yVO���Vs*� �@|��i�;��4�s�-�Wk\M�m�Rm������D�JT��|D�m4� ׶� �Ok�f�c� ���L�5�M&�C�p���	��\���e�#{ �f�m @|1���V�\G��.���v&�5H�*,��Ғ5
j�B�*H-��u�=�����o��f�X�Zi�^��v�u�w��s�l���ڤ�Q�q�&wu./-�A�h�c��O���s�	7L��ӌX���<UX�o�� �{�[��dy��m�{��<�Աt����Cd O�m�A��������?�6@ �x�x^��L�\���`�>]��b�c���h�nɹ%;S��~�n�P�/Os������/����v�0�_�.O��9�P�o�6A������~��&�1�k;��e�ra'	��_x��;.�Z��` v���}�W�EEV�0^�fۮ�`L܁�'<`���i:h+g�K �ʶ�""��׫j��ZpK��'�!�p�q\�ř�3jဇx�����U7�|N��J�^�q��� M��,����"!��u�J2���L����� �_K���h�0���G����M�bU�H�C{E�f���{M���6���� y�i��G�Y?�����y!�w���2�On�3��NAb�����^|��UE���c6w�no)ң�w�X�kcro{>;��ݳӽYR��	ڨ%�{����������%��xA��Ϊ��<X~�"���=�X�=ʗ<6��{nD��^��O.���䇏���f��������'e�Y�O�]�W�r�B���f�|���6��eARp��������%SDu��l�]��z51X���h�:Α�x;^��/�wgM2��\�/�{����DM�Ooh~[)�$���p�䨶�[��4/^x}6j3׊G�~��g�Or.[!����w��������n'=�=黓�Y_w�^s]���'g��n���b񛽕:i�?_3��x��!t+ywp�;Z��e�(:_�`	Y���h\�ow��4�l���:�Q��{qT��,�e���śK�ɓVFa�Ӟ z�\=�;{ܻ��P��ؒhg��}���yX��0�����U��5s6���c�^��s��b�q�=�w5�`���~m,Q3#1�P��)��4��f�2߮y����(��Xｄt��}��+�Ǘ�c��Ix�P�s��ڙ��W��7'2r�b�6���j�!
��r�>�0��C�w����{nv�O4�ħ֯c�|���6�ŏ�U�z4�������Lˣ� 3{�Ys�r����
�v{o�+��y�i�ݒB"��}�ak"�)�}�쓧�;t�k�I�=Y�J����z6��%����q����Ԟ���8���Ǐ҈���BI%��(�/VQ�y�w<��d��C��2��d&uX�E
e$�����H�H��"��N�)I�#֑f�J*�NM�*�D]��;/ ���?B"*:Nr�;��HfTr�p��>!�L+$��f�w\� ��5��5F�.�\��\�V��.�u�#��=*p����xG�5bWF���wB�*(��y$Py�&z�8J	��Q^�U��|o-+�<$鑭a�;U*ҹ9�L���9�(E�ΐfU�I�r��U�<���'�x!�@��N����$��n��.;���Br�\8���*l�P):U�U�G+��5[�teHp�)AE3w��\P��wU
rn�t�-8�J�s��U�r;�x���Y])&S�����v>hﯯ�5v��M���Iqn�gq��g�<�Ȝ�i�us+\�P\�n�0qs�u�g��&�z��&�6�^3�nl���[�G�H��혳�9��q��]r�ݻazj�h���b��k����X��;@o|v<f�q)�&�i�`S���{k�Nɥ%нf�96���el뚱��m����.M�\6�=C�6�\�mL�z��ݻ���{Y�Of6gn�Ѭ:<�6����A7ol�h�l�_!�d{g���WYi�;>�Q1�0W=��c��i�p�6��c�����[�k�.Yi�wtޝci�ϥ1[�κg�ɺwmfM\�;Z獩���s=���������s����/���yɵ���1��+�bS�b��9��%�^-�zN�Ÿ.���Yj�c�x�Z��NM��%l��yF�����s�{m\��f�N+.0���K\p����NN:뭺�%����s]�ڄ6ʡ��m���3vuǹ�s��GۅԷl��j����<�>۫��n�ѡ(ܧj7aՎɼ�I�q��66����9�ٗ���ؕ�ŷD��^�͛��җ֔�ݣpa5�<ְ�ph���l]���;���竳q��W�s61��6N8�z�ϫ���xg���f���v6�X��p��sƍ����`��gu�V����fw\�;���ܺ��6eWq*pz#n" �CV���NHZ{[���鵻V�mi�ga8�ke���o3�4��89��X����m�V-mAQ5c��:��:ǎ��-&Ѽ����[�T�мq�]�Թ�f�b�uѮ�wn�!:k�]h;q�q\nNVIL�������ۨ999�ko[
�C]�C�۝��[ta�j���ӆnT��ݻr�X���[�ĂZ��I�a�ٕ�qa�ݻ\�WY�G�%��ط��\�:�d:��'<z˭�.���O�5�W.�ivzz:��u�lR�p�m�C\�Ļ��qm����8�BWj�=^:���{��wϗ[:"􃹆��uk�ڔ"�ue�5�ۢ�i}���n�8��sv���m6�,�-[V�#̜<�[��71�b�s�x�<-�����(ge�\:��o-�s��T�Z=tێ�'���s�Ѹy��EYлY�dڡ+��s�iݎSw5��/!��O+��7��y90��t�A�ت.7ony�+cj�ێX��ϟ)2��m�֭�=�Z �� x��M�d�Dm��f����+���mgk����w���MD�B�����z������%��u��sS�^�ط��'��?� ���p�Ԝ�R)��DT"�Ƒ�{Zi�{�����r���` r����C�� ��WFО�־��S�@���b����q"�ݦ�@ {�i���K[�ɨ�ܩ龦v!��[�p��_��0~`{��i�e�%�/T�Y�~�j�g���"!��w�8���:�d��� _���Wt�H^�6;���J����m�ng�ݞk�q�͋�ytk1���@���M&%���i����q�B���ed��'\���O�l��u��>�Պ�z��<��7<[[��ٺ�f�xf,`G��ʉ'�1*�d/& �{ߥ���t��1���^��4�=i���5s�)U5P���|�z�#�|�ޓJ����6���nL�Do��@j�x��<(�^9F�=
T�~�&�t�}��s�ҟn�t�c<���.�#���{�]r�~�����[@ ��OK��M�gc�^�ˉ�T��F}�OmD�f!R(EKGy��i 7%�l����3{k.���π����L� n�Ѱ~�(���*�%s�Ew}Oݎ�F�j�T�� A��� �K���az�5��,Q�b�W��3oZ0�����������l1ϺԱ�S;f~�FW�:WY���s��u�Zm �U�� ��r�>������~j�m��;�mJ9����[�o%��^��݁���5lfg�����_~r������m6D��Ʒ��>ٙK\��=�{�>�_:�飻�i�BG�$s*�i2^�TDzaE*�b�2�kj�2�8۟n�lOҔ����Èd�S��"!�G�,��L��q�}~�༙�<V%����U\�{���, =F忨^��5^8�}�"�ْ����B��v���k!��A����B��l�|0��	�;����s.�.��~��/^�3Ǌ�?{���%�}�f%�_D��"ީ��������E2�*�aA\�|{��aj Q�.}�=` �{�K�=�-%o�������PF����Ơ+�ȻJV�2RO�$�w�+�u� �~�*���qF.r#7��6�H����> {�j♾�~���eڅ���s�}Hd�Z�G\m�@s��s<mk�l�n����:9rs����~w紓V����<�:[� �=�� y�i��r=���o�������j�L�K�bD��5���� }�/���1���b���*w\� �{�i� �}��G:��v��q0R�Asߢ�_L:����� >��M0@{��1���}S� }�>� 	7�4������#M�nۘM�ht���o��O�7��� ���` f��%�����y��-��4ٔ*U8!��aH���e���u��\�OcV�,p\\�X�\*����-	�����fRt��rm�V�#u��  >3�����N�3z�K�!���Њk��	+������gD�����s]}MH���i��>ӈ$ۖ7WLM��OY��.�9����^�s΀���\�O=��u���*�=���{�����	�E}TT�@�t���0�G>9��q�BP-��M�͎�{τ��Y������|�����}0U��v������Q}��a�:�{�[��PT�C���� 7oZi�gy�̍�EO2b"��f~���U6�ʻY�` oom�b��ؼLz7cd���{,� |��l�n޴�/T0� �U�ų(��ss�S��}�yi�H ݽ�l"T湟{\P���[��@$n���SI��b(�*��W9�ז�P�z��j���΢��e^DO1egvհr��d�3n_�'˜�حGrMQ_f{��]<%��A�����S��e�b>��{�p�����o�ո�2�%���V4�4�^�X}��͍L���A�� ��`��>xx���x̏r-��n*ĆF%�ۡԌ �=�������zZ[=s�J�uͰۗk�+�э�9є����i��Zx:X�h9��'S�g�����]�����n�ͬ�/p�Wg�s���}9�d-��'S��������v8�{7m(�ƶ�t"nj96�x�=vq��r�zx���7\����6�ؠ��u�ߵ���q���p%��A��ݻ�v�a$h��\%bN;wk�5�x��?w����-�"k#��9�i� r�چ|�s\��ר�8f�#����i�@9��W7߻�����m0wv��$���ou��omy&"��֛A)�V�%i"��E���MSt��L܉�=D�QJj�l/{�V�DN{j��>�=|dx���������O��>s�Q �R�f�1�Z��v�R�/*b�Wý�DfCw)�]ͷ�/w����z��}̘��9���a/Af�͞%���n(37�!	�=�*9�D7M�ӛ��!�;؂Mk*�+-����;�0�wga(s��ʨ��[k�Y��xze[��p�w�~=��[�C�x�">����ҁD�3�tJ�D ^�mwb;�/[}�ˮ�(��l�	�z�5�w�_c\B"fa
�Bx�B��}�+�3c��ǳ�rǔ?S�59Z�v�nJ}�=ӷ<��a#W=����4���7ד�-�������=�Q�3xg��:���񝿱�G��@Ms��߾_|�������6�0��4�d����s���^�5{��qi0������s�Go�N!���2��q9={�^]���o��@ ��4�q�O�&fj)C�������/ټɄ{�|ڸ� �{�8�3oZ߹粰92<�4ն�� �}���

R�T� ʻ]��� ���J�d���j�}>^�� ����l�zy�[��;ēT��\C3�.�Eb�9����,g]����N���=��D�'��8�����L� ��
cu��8��/��M0�"3om[��ssgs�8�JX<�yn"�r�O�L�w�F�D)UUB��9�o^ڶ��g��d����.��" �1����z�LJ
^�'�Bו�6�Q�Y����8b�剀HxEy��]�(
b[��=��Q-�c�'w7�̩eQJCӘ��v�.��z���'����~�juf�Y��̑x�.��}�sC��h!>Lj����M;�S���&"3��İi����0��Zl�o��D�4��|���i��3}x)wX3A�=��|/<�iA>ͷ���Uu;j��ã 6^RP�N�s�.� 4C)L�}r%0|��mdO�q��z�j{��aՈ$����(�2LX�6�N��=C�^���Ұa��RG�������ut��+�܎�{
�T�T��f�}P��*UM�wkY�{mC �ٶ��7��M���	y�4�d n<i��w���|A%!L6���6�A���I�2��j�#>@s_�o� S��q�>x�E�k��E����U�N�Xг� DD0��q5�1��O��o� Nq�{ذ�ە����K7\,dX>oJ(1o=�?K���HxEy����jw ;�Y|�"6��JXN�m� "��"}�q��Z`����6-���;�A������M���{��{˽ͽ���|�q�:��9��po-��I5yۣs�1?�� ���*/�I���vES1�Ҫ W�����`�_�e�̝^\��y��v�\�=��H	�v�4�֚LW�e����y�9n`5MG@q\���	��i�ێt�r\�xά�Ħ�����/"2��.����D7O3[-��;�V� �u����y���W���g������ۆ|f�2�"i
UM���	1#M�.�M�L�����4��'{��D^�m6DE̳�z�8����N&� Z�ψ�)J�m"s;M��ʑ��i� $��ź>�:o���<ܷy�i�U8#W��P""<U���m5�Ϗכ,ľj�$�����ӈhn�J��˪�Z�A��W�}~ܷ������R
TE(�T��kM�6�XƟ7����r{>Nsm��bX4��ɉ'g���1-��P�������Eܣw�A��];<�Q��{�=���'i,G�Ӻ�oo?=�u�)Ku}5�y
_�����q���Bɓ����zii��G����2�y�S����(�nM;c��n�X��Y�ϵ���:Z�\��G6+������gQ�趜��Mc���fě�����Ԗ�-<]G<�n�[������q�J'��u��jm������k���t�u��:��fgvo[r�q�Ld����Z��u����t3�L��5��p�bOE�&M�>�Bݩ��k ��/X�q�u�{&�wiN���Q/&��]�l=��s9���6�vw�E*
��d��c�* \���� ^{-4ȁ�^��h�Di�������z�0"��y��%�#*$��35J�T;h7ܮ�� <V��x�^Fs��W�> ﵦ�}$JF=��� ^T{�ޯB⧷� �21D)�4�*�����i 9{Z��	�U]A�S���� ���d {{����2M*a����9���=�)��Ns15Yr�f��;<R�r^#�Q�K�N���]�l�ݫA3z!3�T�UT)�r!���CDO��l#W��YWxw�f{Zm ���M�$�nۆ�#9ҹ9�;\�u�TC�%Q���q]�ݯ=Nw��ۯv�^;=2���1�7$�Mw|� 0,  ��⭑$���s-�` O�m�U3��9�=�{�����=}�W�z��*����+�����i�@��r��#�L�~�㍨��~\�v>���'p�싸_>�]����N�{��A���?h^j��~�$K$7隫+��7�M�� ���?�󖱑�y�8���W ����zyܾɚ�.�V�HI�������D�J�M����l�N{j�)|���)r~ffc�7=�I$���.�"�h�B�QHR�o�'[k�n/s����hH�붸r"C/r�"��!�������su�!�r��	�.f&��1q���� >�m6o#fe�}�r����֛�j{�b�!給��Aoe�K�SU* ��U"��=;Gg�OT��'Z�`�=rmz_#ջnSX����;��*R���f��f�P�������J�3��0��l��뮐��3{�����Ip��a!� ������O�o7������{z�&| ,��9 �{m6DD�a�!p��w��]L۰[�C9�4z�U4[u$=I+�dIA���?�����zT^Ͷ�;Y��C&��pdֳ���k7ߺ�y���K���,��vv�T�{Nu���SD�ǹ@=Rg��Y��m�X������W�>>���@"e�gX����s}�r���#6==^{xu�2�4xཾ/Q7.z.���y�7�y�x4�u���=fB�Q._f���w�ґ��,����w�D7�r7��5槝��ޕ�}�z��f��p�޳������g��A�%�gȆ:�_g����1{��IQx��O��x���7qY�����$9�Q���<�Ox���s���\]7����y�}�J�i�n��˷a��+C�=�vaW޼n���O��y��u���2�F_�N[}<gC����4��s����۴����<(�z���Ǻ����_clpe�\g�n{�x�n�@�u�h�q+�qm+=&�2����cޯջ\����KS=6�w�}�C>x��k�6ʌ�<�p�r���nG�۾�4�l���&�,��<\�4�{����z\�ήc>~�cG9���B{�\���f]M�z�A���n�m�w��_���.پÞ�k��������D����Y����{}��|/esw��kO=Q� N����X,T�G�]�2s<���j��r�>z8^tƳ����/�mԻp7�ؕ�w�s�*�Z��8�+���
����{$�o���� ��s���:��sO7������z�ā�#�q�@�V���3����	��0�Y��zwg�\9��D]���=�[I=d�G�$7H����f���y�T����������3ǀ�O�޹aei�N�S�Nq��w:��N{����#r�q*C0�wJ�/'qj��"���M�s�Pr��öN��y�^�lٞ)�'���I5�+���GCs�u��]tD^I*���uu����]tq$�\��uK�8A|�<�a}�dx�����z:�W5/Ju۞Mr1<��c��꒢F�'�"�D��B�<�ԏ'!tn{��@���<��Y]U��r�dn���^l��'D�n��Iw$-En�����)���ЏZ��&�r!���m�w;��n0Ԓ�u�5��J�4�֞��mɓ϶�E{��C�q�;�C��J�'q�w�E��q��J*s�e1�=Ii蜸E�p�T�%�ADDA�fZ"`���ʁ Jȭ���c`6���{��_h��, �ߚ0��bD�B4;a��nv;��.ϻ�  �7-����ӈe�ڙ���Q�Y=�De��'&vXb�C���:<ϩ �����ۇ�����j;�&"�l��Z���ƛ""6�o�ُ�rg��b+��n���հݎ��vv�]q�Pg��Kly���e�v�\d���]d.�������;������j� ���  _m��/Fg*�Ma�t�9�r� ~�4�UC2:)�UQ5B��8���o�`{�o�L�h���	C��h ���e|J�z��]Y-9�o�2�{�3��@f�")D*���i� �e�h�+���7�]���� }�6A�F������=A1����Ȟ����$����ō ���Zl ��i��{��w��i�]�n��L�-u�����P����z �� �#��Y��`]O���a�������Q�[��G[k
A�U[�����˙��ϐA6#�8gĠ��"h�a��m��G�Gsa�J��[����}}i� ;~ƚL��S��g2�F�m��ehJ��tl��N3j3�;Fܾ��ݛ�ԝ[x֮���7nf������D�"&��T��;wkS
�fC��mCD�9�Z@��>�ڟs��+o�?� ���',��TL�jd&-�e��>@{k#��S*;W�>��L�ƛ =Fm� <�j�'�k�u�X�}U����QD�
���r�m�H��tC��x���g8�yz��#��i�@�6�V��Ҥ�C�e��C*y?Q}WpD��a��y�-�" [Y^dC���։e�ro݀�x��%3�;��D�I_Q+��^��[�H"�-6s��V�ЍԪ'w��H;��[ �k+X��!ﵦ���Y�h���f6�:Ri��T�3$=�E���5�N�5���'[�{r���C<���)�o�_}��V�Ƽ'o�=����L9g�9��������,��Hn8Rp�s����cۯf��vM�u�P����ƕ�n6�.Mm��d��{=[��u��|M��axn+nN݈�^���͵(�j�-�$'��E����d���Z��v��n=M��qO+ݸ.�ۊ��Gl=v,���Wy�-k�i�L�/\pj�ѭcn^��Jx.l�g6�۸�w{OJ��#Kd�|��!��#j�c� ��4�';�H�'k���nl���uڊ2F˲�[0�RL��)̍1�A5"j_����m �+ӖԀ�֛u��c=�t�x�L��v������)�DM!J�i�m����"�	��9�wj��;[9c@ <���
7����W=S���+��P�eDȢjbf.;.v�) >�m6s9Y+������՚� S��1�~��O���?�UC6:}(���W9���۸�#�-u_`�� H�s��	{��h ��Ϣ�^\�E���,&����a$::�����N����a�߲���Q�f]D��dCH�|��N`[�?�3\������o���7-g���a���hN��qYǝ<K��\'���������3�9�K�*��G��@ >�e��� }���a���M������s��W�֬�j;Y��3�ROb�l�<��]�F�k�俍�$�a
/�^�_NK��w�}�J=`.�#�L����R��uN�[��S�<g�����ڷ�H��f���p���6r^��K��MO�����/����� "��i� ���6@�d��x[�}z��c�u�:B��D����	��2 ^m����Q2,�zV^È��wр �cM2 ��$�,[�2���Qm]#�5����˘��gD:����@/_m]��e\R��t\�ڿ{B9��U�x�QET*���e�`DW�*�sڋOJ���eo-_> /���0{v�4���$=�P����w I5�u���<��v��v�gML�p�g][��8��[���G��qn�E �"��ko޵iF��/2چA^ͷ>�w��l�&�K\���X6�bəe\�r�zU׼��"���o������ o�j���p�3��d�����ߘ%��FeG�MB�MK��o��pπAY�h�ߦR�K�^�̂;Yq�����yh��j]ٱ/���n��{��.sK�+�Ǿ�7��i�8N��ܽ�x�-j���
�TԦ����7�{����O|�~� �5����n]v2ALg�T�*���o[^ݚ�y��@��w�s����� |�e\4$ "��k��Q���,����L���mD�T1l��S �m�����˺�|�}���Y�̪�� ���o�i��*:�;�#�!�PI�.�C��;dT|:z�텀����y<<W"�v����P��?7���<ET*�����| O�*�  �r	3<���f����m�z�t��3��h`��հ���G��/��s�Bp�#�㻑�#��]��v� 
w=n ���O�@��zlrN���3S��8�1�aHW�4����6 D_w-6�gSxGb,��f�f�3 ��(�@&/�D��Ҥ��A,�A`��5�c�W��跛V�Q�A��j�� ��ƛ@|{����m����p�dT�`�Q��<�,L�~����8�����&��!E-1�f=][����&<㇞���Ie�b�P��y��ɞ�6�>������{¸��]ܢ��Lq�f��C�qB����� ��Z����8o/����n�$��cO�A��{����7f�̟�g��]zĪ/�+��kix���M�맯&7AS˜W�������� ]���W�|��M�kݧ�vV��$���](�I7�F��Lj�8xj&�U\�>�f���y��zA�>s�q� ���i��<�l��{܁T����9k��T���D}4Ƒ�wZ�h ��5L@*(禪zvs}��HH���WѲ�f��,���ML9h�TryD�gVN�t=�OkZ�/0�2m���f��g9$���0�Ay3xm��}���é'�*�b�Ή'k��30���|�h�R%0|�FK͛�`W�m��#��������{����ڽ�5�3�Y�l~�^�8{�����c�
�G}�1}�
�\\��ɍ�qU���+�B&�=L�C�%�~����$@��nյ�9�=�<���N�r�;�]��V敫=nw&�����"W\)`�9�i#"�9���N�]][rٵp�)�P<x{[��*,-f��=�g�C�pz����h��q�y��ð㇆�/!�����C]Y
z�"�Au���ol�GJ�G��<3�`:ۣ�r���G�-����:�/kl��7%�����z�Il��G����z��ƭ��.,�b��n-w<<֠���޹�E����H}9�UI$T���M�i� ��f�����i��ezƋ{{�9/}-&	Uj�V�12E0�k�O��3RÌV�⵰���٩�9�� �ݖ�A^ͫ�����s�]���n<�UF���)SET*�s�³�� W�*�����}�(�Ы���� :^d��>}�na�wԪ��c�jl��4w��vL�\��ff���N 	�ڸ` y�؃���Q�DDI{��y؄I�M)��\���8����#J	��j��Iȁ�K��3�&f�����`! /}{�y�G2��L������Z��c�uFW��b�W ��ȷ��V8�q�zh�I��x{��	1������%[ ��U��H��nA��'ӗ�Gx�5��� 
}��M��1�S1%\�']�i��u��]��r9�;ܥ���w��2b�o���Z߹��Y�$��w쬠J���(�M�t�0��i.�mn� ��`�S'!���8�3OM��\\�rY�W(���}��~���~���	ݟ�0����2���5���-��˝a���Al��RD�s��N7 �;�lq���L��3c�oD癘>�y����`��N�f�*�j�U�p8V麟�>�Ȕ��=�]�  W��M&� d����鈍S]�+g����X�V�����R�PW�@}4Ǝ�1���x�9��ۘ��π�u�0	�֛ @:�[&�f>O�ߧ�����יW�ݮN;�Y��k�0/E��뷒7��(Q2[�D"CR�S!T��G�O ��M�2u��;���?lݚ���ķ#�g�5_I*��<��Yk�3K�a�; �d],��~�p ��M���%&Ȉ�x_�}����
�:zALo�T�I\��>'[i� |7x��y{�g�j�A��26<��otzc���k4���>Z_�?n\���l��e�Hҭ�ٞf��ew	٨�0��bt�e{iy���x�b _�ߚi����0�U�W1ໆ�f.� ����s���J�$����$�9��� ^��O* ~�DMs�@#�z�aUx�SQ5B��83����Y��՗��;���Z��#�}�i�{'l��]b���t���q�oa&ǣ-rN���g�c9{u���+�\Wm��Z(�532�����ȪPW�(>�Ԉ��Z�Ј��ɶ�}3%�'lu�[�ݾr)��Fe�[�90 �oe��<��"Y�����U��ę�ѣC�����\`� ��9-���c����r��v������sc�g�5_I*�l0�<� �����+��Ǘ]{���| '}ɸ�흱���L��3⊒N\��'[k�}�ً�r��6|�h������\��D0>/{�_�K1�����Y*�b�踹QR*G2&�E�,XD�:ۇ�����U�mb}m�r��vx�p���b�'Gw��\[���n+�x{�1$�k�S���O��!���C�b�R�O�bJ�Y���c���#+3�d������c��֟��W��ӰS*c&�D�UH5X��Ȧ��o-O �+��fλ'mۧ��ň+��:i��*�j�U���u��4휲{ݵl=���u��W>h���[ ���&%�E�Ã`�-��5�sWs����(4��,�<��S _r�� �E�u��io!i��=7����Oױ�Ԫ�d*�9�y�� �e�� ������}����&�9�|���|("��i��ّۉ3�Q5_P�����n	{��|���W�����S�jA ��V�~�N���d�L�9�W�O.��	�;0H�ꒂy73�"q����O���˽�L��;��@_��6A�	8�_����O���y�±O���|l{ʧ.�%��1��`��K��G}�k&m�n�s��N͞>���m�WuL�^��2��M=��.h�7��(M��,\����Kwg{�5�%�"�e�j����6�y���1���7������ w;�)�;��e?5T��m֘�u�`S���)��t��.����TV��+�fú�+Y�v����ɷ�zr��Z�SY�����b�O�_V5��=�xd��~~��jdէ�R�>���7ۜQ�=۝��ާ�+ʿ�F��<��xL���s��J���s�Z;�Dý9\ -J,1*�ݾ!z�?L�Ϗ\���G	Y�!���iȱ�ԕ��)���I-��
��պ{+н�"�/Ӄ+�}Iw����d�ܾMX��b{�{�מ�x�wm�J{��������Lo�1���� <�L��M�VA����u+8Á�����̴�^b�x�?9����ٞ�3���W�c�8c�: �^4�J����	Z儴'ǿ;�x^��J���cg2Β󓺮��s�w�SA����ҧ
w$����փFp��p�9c)[&8o��W�窒�(3=a����^X���w��>=�`Ӹ�����;��|VM��<�#n����}�\�g�Ux��	2�6����s����n]����㞷�px�����Z��{�gf�6/z\��[V C�/�ñA�l�Ĭ]%U�X�]��3�:OYs�O}�lb�Љ���8��v��A�������M�Ha�{�jY
ɚ��_o}yBBs{��3���U�%��z*U:%&^�$]ʝX�+��w\�ʮ�s��t�y�Ъ��Oq���#�\����y\��֫H*�:,��bM��s�<�2�z���T���f��%�8L�!��XD�)��y�/Gu����D�)dL�W�4�D�*���=��$�1"̩���Nc�q�H�T���ۑ�{r�X��PQy��Tg�N�b�F���s&�b�Bz*�z�-[)�j��(�QU�f���D����ejw)v�*��6O�y˷�Mn�:͚`�T��;��*�NY(��rs�;��"��a	&DP���Ix�Zj\�w"�7^H��>=�'vi�YQ���H���<"������:r�)?1���/���-��ƱWc��w��-�//0�b���6l�pO���V�H��7v�NvQ��{n{2�)p���b��v�v�;Js�A�gx]<q����wk��q�mq#zJڧ���=rl��A	ŷ�nC�ʧ]�H8�x�n�m���s���W6�LO�\�tg��<n��۹K��y�wY;�|���;0�����{����۱ѝ�	t���6�9ŷ`^�Ṻ�̜7>�Ș��Ǩ��k�Q�����.��:xn�Ō�[��;Ōnz1�y�m���Ek���\��V���<�O[<�LA���͔��k��˷��O��{]�M�Eɇv�q���K�j�\�hl\짓n�G<��60vȼwI�K�G=��1b��Ufote�l��>Y��1ԯn�i�����m�x�t�LlN�7=��t̼�D[�8�u��v+�V�!L�����<��g1�:]`�7[�y]گ=\[���u8��]���&�7k��u�Q��6������dB؏3���9��ƥ�p�i��s���=�=u�����77[�}sܖ{n��
�u��κ���L�e�2����@=����fJ&r#��6^y�e���Gv�Y=��s��ؒ���م��ѓʘskq׍q.�'f���jn����;c�X��sͷa����E�(?Y��v�h�>y���/ lۻm<���G�{7�;ct��G[�yݎ�kS�=�9:tn�����m���r��n��R���+�n���y�Ϙݶ6��nֆ��s�GQ��3�'%��n;u��[G=��T&���E�<u�Ah�񓶋���k�x�����O.p��@crq�SF��4޵XڷZ炭�n���4�;�r�Vy�r���b|N�s'Fz� 6rǊ�a���</Goq��(�8\A4z0�pv�9���:-��l��i��Rx{7q۵�s�� ��%��n�D6�y�Gn��;4f���s�:N����y�ۑ��q΍wA'<.�N�q���hO8���$J�O6��|¿-�Cz����瓕�H}��c�t
2��q�A��mM�)��N�p�u���w]u���n�q�66����inq�phnz��=.��ֺM�[vdロ�
78�n�ۇ�.5���Z��ۗ:�y9&S��u	չ����G=���.�۟tu�t�22��j�V�_nT��wZ�Fx�Nj�1�[��z₹�l��]�WQ��@7GF;l���m�쳲D�n������DY9xٽ���C�|�#��K������?!��� �����e���OFû�y�LW��]���r�|~*���vD)���4Us�@�oZ� �k�`�{��<�< _;��!'�	��2�ܮ8�����߉+���`i�����=�6D	�-�l��g38z���L��� }�4�dD	��0��9����H�\���(������r�~�+~��;ݴ�rd�-��>�ejh�����:��5���w6�ɻ���0o�gva?����$�����|������.z�"��m��SѦ@�����a5���;u馻�K��~���Yܡ������z�O���ݪDy�x֯`]�q6f�29قE��l�*l��|�M��|��K/�;csy���|��En�Wy�\C@#�OF�]j�V��&j*�bfD�'[�@{��rWNŷ������x��O�a��$ ��3s�����v�����ߩI��ߌX��T���q���J$J�w�n�>���yZ����m<a��k��ؾ���vMh���k��`����DP@�����_�rڒ AH�v=s��O�m{�8�H�O�" O�ZȆ�oqp��Cy�y�2kY�:�}Ůi���K֓� ��c��/=�5���y@"�64�'�� &}Q����P���L�l�R��A�պ��^�A��o�^��� ��A��L���.�	p��;�����b���6���2ݷ]sێ�S�H�����C��;��RTDMW�3m�9ιq�N[�A 給®b�<W{���y�s�총�"d'��1��g�	���+]妩��A����Np��yT�t�� _;Z�@|^�Z2lU�2�T��4�`�`gx0!���'��@ ����L��zqs����+��?R4�M�����)�AmY� �W��2,�`=����` >}�{:v��C"�Y��<���|J��=V(JD��x}�O���7ѩ���3��4޷!��������V�W5�L?V[Z�w^���<�"�֛H >��(����*5T83RQɉ^;H8戊UB�}4Ǝ�cM&  �Ǖy�ȝ�}��-�fa1i�%��AĒwWBMW��3d�i�I>��؀]�v!�X�u4�'q�ηd������ϩMs���@�s�� �}�E�j/#�%��{��B �{M��ő�;���-��l�n���̵p�����"&�Ꙋ���:հ=%I�ӻj��~�|�_� _3l h5��"#�X��z�6{��M��I0��B���-��i��Go5�"b7�Om�6��\��:� ���W�^m\5U�"�O"f�R�	m��p�v�8��v
��@A�}�� >���
��\G��V`r�7.�5�Ax�a.�D��n��gU-��d�=�����[|��0�s�;kG>�L�6�B�t2��8��K*a������<=���v �@�{�3�Aw0b�:���~��a>�W��Y~���	3NM� ���3�QL΁�Nb�J���[~,5x�ۮ�a��{:�ۮ	q��7wl�k�QDDJ+��)XMU
Q���ǘ�L>e�?��"+ٵp�ik�v�Eq�"�8g��$/,��f��*��p��_�e S�?����H<{�^����\]��  >E���@^ݷb����y
�bS��uWm�L�x�&DDMW�3;����m� ���V�����i�4�.��Ws����LU�I$�f�ǐK�!0�+�j �/�'xځ��]���E���մ��^ݷ ���^��ؓOP��}�e���P���;�$�B�T�;̦�H"/��O�o�Z��c$�s�� g���
�ݷ������>���p[W�J[+�����+�g�DU�B���i-/�c���Ci���U[�A����|V"��کԜB#�{���5�m��1tRuD���,���kr{YH�ĘYM��#Ƣ�촺���/��B�/�X�Vc-��e����q�Ѻ68�_��þ3Ymq3�c��k;�g��ktk���Z�fǹ�e��H�V(!��ޱ�;ۨr�k.Oe�2r軶��=D`-�}�P�Ԛ�tS�':�s���<k����mۃuŕֱ�08��m����b�p�	�xs��m6�˭�V�`�y;�p6�F�ۃ�?>���?|~�J�_����=�� >
�e[|ﵦ�w��R㖮�Ƭ�u�D�OF�J)��٢����
Q��:�Zi�z�{����,���̃�� �_V��က���6@����g��~���q���@N)�D�&��#��S�h��M�@�������G��/�^��XH>=�v{�:��cL��M��yA��s����a����g�}�h >���M�YY�j�6��@*y�p���	b߮-@]M��M& ��k�^�p÷��#>�g5�����I�VNiqɨ��j�<G��+�U�QH�*sյ���\�{W�Xy������Jv
ys����m�y<��T��sQ=��iI$��M�[Y�h8�<�=݀;��K�� {�i�.o�~�*���U�q��yT�3?WSu.���{v���[tC@�C&tw7����t=�G�;ՇZ��8�a@����44ݸ�Fd�ة��}p1��	��ń1T ��mI��0��I|�7���Q+��i�> �����n�N��Vקmr"Wf�*�R���g_���
ܬhq{͚�{��nTv�̟ �E�u��n^����5L�$�L*�3%�#�Ƿ&T�J�{s�|��M{�(.�Y���tE��QoWd�Oe��^�X��jMQmu�X��e�]Ż���1��M]�A��ѥŃ3���3mB��
,���o�1��4C9g��X���xӎ-g1Ȼ�uǖ�T�îUۄ�{,��o����LR��PS}�s��� ���1 �z�n���ӻ��MTo}���l� V��6
�b.z���J�%�,��i�c��%dG#j���k��+����`}��o�$fl�_�����R����
d���W9����3��^��l%���c�+���WK��z.�6�A��4VF7g�N4y�}��g�_��7q(�TY�*�Q<���6DMFD,q���dT�任�[����Ֆ>'�]��6@z�~v��6�R��T)G�L��m� ��g-Nd�ܠ>W��"$��]�0������a�G7j,~�FJ�U�vwg��0�.��TVu)$�=�#lց�v[��駂��1��b���=}�� !��e>?n9�����s��]%��'o7F���6�g�����o&,����i���?��ꍆ�4oߟ���]c߲�d@�kM�6R�s�y̛"m�O]��d�oq�CN�q�(q�D�f�y��� ���ڻuw~�˝�_� v�����y���bNn�m��Dus]]�i���3ĠDz�*j)U����m0{�{2�>`�H2���k:Vs;����Y{�qy�i�R����d����S|VV�<��1f9��ǲ��%H��z��?w�6�$n;�H��,�ݫ���3}������r�j�Gs��Lo[0�o��z���*n8/Wb�ޮ��M�}z��O=}m0�^�v^��������}����?G䀏g:����MJ6���J>�cG^�i� ���<�~U{� �z۶�@��W����F㽇�9Vx�Q��q0 a�E,�^q��E���z�\s��`t��z���Ǝ�?{�~��j�
����q�!�e�dA����`�<�N��?^O'�����q >�� ��n�����ߩPܲ,�by�t}��з]�� '��M��|nL�Jf��b�;�n5<�����P/4е)��o�m;]L#޺֐� �qY����j�����͚�1,V�"�Gv�a���
=Q5��m�'����*߾���ȁ �۽�����k0�s�;��Ʈ}*��b�*�U\|��E�-�������UY�Wy�e�4� ͻȸ���|�3>��*����?qQ]�p~#?~k��3��CP�Ww�G�;��~����'�ɌTOi30�m��-�=�� �db�k��a�Tô��a���>!�7o����f�{V�ŷM�n�F�b�N�Gt6��vB��<Mf2��]�v�\pm��Y�3�.�]�z��mJ�/����vQSt�<6�\ޭ�k��8�p�mtl��Dm��pz�m�+��f�^����$���x{#�A<���Dn��<v}��gu�c��q�I��uB�@�e�PQ �y�9��v�={�x��ŷ!����&����/5�7l&�;Z��\�;={�fOF�+�ƣu��*؏Ͽ�������?#���� =�X�� 
3;�Pfḵ��ŸfPk��$�Pkɜ+�<�$'�"�AS�B~�~dG�5��)��y���ڸ �n�C@(~�v�	9r[�F8;�[�3|uUER �16�݄���~$�G~_�>�rXH�w�Neǧ��{�^���w�� C�k���!��tM��*��ӵب�MZ�zJ�� cu�3�>�v�/w�����Y���D@��_"��DB�TEME*���<���`��̎Tw�n^��\@}���o���.� |^�4�5aa�S��l��(@6Y٥�^y���f�F��A�ڞ���i�$��W-��S$�TUP��5�ֿ�2��Q ����H�mn�4�����ѢA"v���5�����6�i"@y��Y��8(�vU�t$h��z��^�H1�m��^���>^�:��n
֟ދ��2|�jgw��_()]u�xgP������GV��|��~9���ĀHٚ�������ix��`��3����4:��S��c�m"�ӗsu.Z��L-�H �v���èj�PJ����n6�-��42�1�g�or���f$�|�A;f8���X�h3ڱ�2;BV�3��4C��n��.�1��O2���ح�۴dx�ā�u�	>ݘ�%Ӷ+'6~�Ǜ��շT�7j�ñ�ώ{sY��M{ts�z�gO��n�(?����o���Kn曭H	+6�D��מi%�;'87�1]�D�˔�o�;�x�kO4��]�����^vo��i @ �m�y �U�Z{�dm<B�w��O�$Pp��"��F��/"	#�vF� \o��|�����5�u*w�t|J�jy�o/���o��_w+[�x���n
����p=��x�����y_w��nqRU�|%���=��E�}�z���G����B}��P�G]��o<9�� ]0�n�_�=;��z<@ٜ:r�������g�8�����`u��!���=]���ul}|c��`{�b9�<�݇���2�f?xq#f��4�{)a����B�:g��Ӕ�ID��VۜV��]�f�5��
��`~PaB�;^u��/_fq���z#"�O{���	��޾[�K�7����ޙ<r�a�ui��o��ӌ��(��9�=�Ivy{����}8=@>{K������3wپb��e1�.FA��5���5���i����=���|�z�Kv��$$�{�	5w�R������{���﷣>��I;W�ޚ=�7��XH�;ؽ�����l�j�o���T�l��g�w���
��5ճ����%{�� gv�ud���\�����l{���6�B|h�E��a��u����ǥ��C��ڻ��]��[0��<p�2�L�dU�^5���'9�#��Mo�����E{/����)�|\�q�	���]�ި�@ص�wQ4�B��c;��.�Ya�t1^�{ܞ������~�l٩���Ϛ�Z����M��R���c�g|��D�VN,�/*��P��-���u�tn�߽�����>\_�⯖ܮ�؂�dȱ{/�Y;��ݲ����3�yFo��=�"쩝;8��׈���g]���W�}N��KQV�G�DJbf\"Nib����s�s�2�VfEX�m���J*�h�2Ӗ�8X�^�G��g��V�Q�{����0�qD�5�$EgN��RJZ,�\�%�nզg4!3)�=B�8��DeB')�i�)"(���IiE$EBd󻰲B�j�Z�X�$�HF-�����,ºI��,#�L�9���,+��$YI��,9�(̥�ʵ�2"J�,�+9bE��/=���)�Q��.�r*AreQ.�Q�\��W����g��U���Q�'0�3*2�T� ��ՐHI�i]�q�*r�:T����%���(ZiRU�9���a$k�uDԫQ�����[�J���RZ��3&�����@�(�N�J����H�$�RNY���N�F)��+�qZ�.uws��↗��������������߿}$�����;;�s��+��W�Az3]����rqbD�Ft�H$�!grX���K�q{�#��9��h�Ax�%"6-@�cs:P+���u@��ԑ�ȐA�ܑd2j����)����ݫ�1�Q=�[�[����*�V�n(3�|7n&����\���BĦ�
����MD.��$O�+�#�m��sM�]�%�l�H$GT�������lWuB`�e�cV�f�� �W=O�ӷ�TO���l�j7&�a����Xw`�</OFł|b�B$�4v�uP�j���vr�[�"����� 7���Q��"�7�[�tH��|�ԉ Lv�O��3ݷ>�6{�es;2�-�Y�ba�j���/'J��7��~�$U���'sVU�G���w�F#�B��e�5T�n��*��x��N��H�3 �,&wr��>0�Һߩ I���X:��J�Գ\z��@$�#�1 A{����ǸQ��i�|_��x��y�[n�k<:�{M4=���Nxڥt�s��~��}�]���o���w�$�y�� �N��7��c�>�@<�bI�'ѵ��2��a�h�P-�8�-R�P8�hsj� �#�� O��� �s=��T�	
�oulEx���A؜&Cü@5M�\� ���A9�WZ�"%�tH$���HH3������Xw`�!��H�y���t6C8��J�||&��/|O�l�K�,쬂�~�� �|;�&�0�x���g� ���ʂe�܁��Y3iMv��;��$	�����������E���O��t+�/�Cx�xd��qS�$Л,�*�bR�||RjE�Ko��aM�w�Ů���/�x6�+?n;����v�׿����ȓ�nM<V"u�˹k`GnW6���*V�u�I۱�\l��<57c�m�냬Q��^�t��$�]��l[87a�m���`��m�k9�u��<�t�P�6��qn.{x�n�,o�ۋ����E��g��β�u��ڶ���qϷ�����lw'0A�WV�T��/0!v����x3������듕�������z�7\twjZ2�HpV�êksQ<�K �K��=v�n9�8MԼq�v�u�~��2C8���h��m��ĀB�Ԁ@�t�󷥍�cy��u$� �w��;�n̄<�Z!�C�ܽ����9o�<���!�v�//kl��$�U�`�tꩺSQڼHR:�� ��C��g$�;=0A ��n�ƈ� �AU�I	�y�H���N!����ʥ�3o9�=�H9jy �f<�I$����x�Y�7[��&:�OՑa݃���""W�֞i ��ΔgE��T듚	�Z�R$����$[�qh�s�;nK���UݧP8������@�ET��D�M�s��m��W ��jۍ*�kƭ���o~�~��<~75y�{ƖmH@�� �H���-��tn��3\z�HM��4�}9�E�g��4:C=�˒�!��Y�nE��0?=}������9{7B��2W����V޸p�{"p����.Ec�-%n��,�2�2l\������щ���xx{�V����$���O�����_!i�;���ū F�,�!��Axv(s�̀�}��$��J�^�bD���k�u�c+yq{h!��<�nS��]�	�P������0�����G������crZ�G�P�3�U��.ԇ4�!�	I�z� �5�h-�x֭l9e6I�C�a "��D�m��U#��E��@J#�PQ$LR
� F�pc���u��u&׶���rى��c/���������r���"�6��>"/7ex�"~�;�6ٙ�7�Ż�����(�45�����6�i	M�c��1:�f���^vJ ����@�frn�Ku��`�U��;�b	�ZqW)H3۶��-fobGC%�*W,�m�I���\f�ql��b�"�j���l���
/
~���}��$/{]k�+�g���㍚����� �嗢Ę�ݕ�A �}�(n���4R��h�>���s����_�W(|	۶� �מl������	-�t�$���F��!��<�-�mI���;ON���s�|Xї!����j��j�ݎTi�&�B� �Q(�%ѹ��M�Z������Qՙ����)\�~��9�����Opk��x�igZD�Ns�0���]� ��O}�3�p�)oZDy���(;�x"�H�K�q&�.�Qq{W(�I�ix�[6g�'�y�9wc�6�O�z*�A Di���DDA-脼�� �>:_e� ��!ŘkNGF�U-D��inZNt����o;�bLZU�u#��[��憞�@/^La�A�����SE��,W)���Z)E�|f�oY�J�3q]���6��n�A��AoK����Fŗ����ǂi�P�aq�Vܿ���-n�s~Q��K�&�i �}����l���j�I=�d	r��<ו��??���[�i����񍮕3s�a�t�qѮ�4<+s�{a.�+[7o��}~���z[�!�D<�-Jy"I��	"r���+e=ŶSQ������]1�OUH`��"C�er^$��͇T�W}�}cnc��g+y"8wwq�����N��1<�env~� �߿n@3���49�3N�$�gLi�9[ҁ1L\5���%�����e8o��s9gˊ��n%��'�woeI;�ߴLf�2����FTq�5�d�v'A��U��%�|I�ʹ�ۜ�n�FW�d����A#{myT�����D�4ַ,{3�yd݂i�����}"�~Y�k��Ć�&�U�A��Rص�l���j� ������g,ǡ6;��3��n_9[�xq���c��}�n��Ӟ�'3r�C�����Bx֦8�s�Շ;L�q�D�������܃��8�ݍv��;#Q�[�
�F�g��{'R�Z�氝�u�;\��a�7/G=�=�Y���9� 5�v���oXl��m��OS�^�6�>�ѱlX��Ug������R����v9�컜�&���Y�9�O��p<Rc��֬��)ղ̝�t`6��Fn��`Ӫû �uU�����u6vX������0�6����u,|DWf�$>i�ٔy��-5dk�׷&8����r�`e�%���C������X`�o[t͖8_^A���@�om���i��s��i�^��7�,K��-R����>/]���������zc�n�	�9/K�m���=�f!��P��	���^uԠH$��yiI�l�ή,K�{�Հ}���'�c��!S��`��[�!x�K�dr��٘�c�Ur�$���K�Nt��.��DB�o9�Z�u[�Fy�Ƕ����fۛl�suAN-�v�^.4vhn�1��\&,���������K�Nl�4�le����W��ۤ�$���}=���c��&Dl�/���*w��f�ݝ�h��,\p������720�W�3"[���r�*u�E\2�[*�,צY8"����+�����/�Y9���,!�&	)��T�Q��d���$�>��D��g�?4�a�6��ʎ�Ɏ@��6��>qb!����$n4�>!�;�a�i����A�z�@����$uQ�\`1�Ahb�F��<��,.y��P7�)
�$���$N����T�]�.��y�k�� �0�����I3ۻ!og)��S�|�M$����ȟg�zQ-S����43����,��&�W:4�rc�׻ka;��z�y�����b�q�<C�-�㫶����A3��/��F�n6N�s�x��GD�2H�M�cCx�C��9�l��.ɧ8ۻ�� ��ȒA"z�� �pn�ۓ��s}�m�Јgw!ؤ}�2I3w�!H�̯���:�FUL��z��å�7z�ܞ�߹��}�}�5��n�=7^E��*�f�:�J~��ڍ�;�:3m=�� �T����Aۍ�$�ޔ	wÛ;�8�1�r�m���j��h�F�t�>$����O�/ܶ6N�8���09&+2�ѐ\`/ �Ahb�i��1\�,���+cj�^����O�"v���A��?+�\,+��(؎�R%T�*���vy���6b��Ύ�vU�4vm���czK�����qf�C�1?z�g	 �7���>��׌��j�'ē=��x�މ�b�q�;��/芠qZ�&:-�fV����Mt��g*� I&w��Goٓ�M�Ӱ�;O	�DkSx��fhz���HW�쭤A>0��9�n��#�I"j�R�3�Iy��ؽ�wq"�D?Zd]li�k��ޝ�H�ܤ#6z �<���\Q�귛x2k0���d|�\�89�sMƷ��z쒽y����@���~#\"���ws̄Nx�cX�iK�/��3�+��z8�`̐�X�C�-�m"�'��I����u�D�fr�3�Ԑ �l�H,ϋ���R���Ji@U�Q1(�J����K��ח���W�m=]�=��7Z������=�ٶ�,Ở�ԁ$�5�I �OD��l4��\��r��P���^D	�L�x1����G���b�l��	���L�I$�=�H/1�yĘ��L/!���Uؼ���~�f'�!��&��r|mgRD��� �z\�[A����	3ݕ!���>$d�u�a������m,sר��Q�܈�m�F�jAO���y �Nu�x-�&Z� �_T�v�u�I3*�UI���ͩ���Qh�[x��D�i��E��H�E�N<�A�����W�����0CSWd���Dbz�?��25�����N3�;�-����x�ѫ�T'�:{�t^鰤���� M�̴Ԯd�����U)I����ػ�k��E�'�o{�V��;Qw�pD�_��)ZZ�F����9�j`P8���	�],���
����(+U�[����|N^��q�W3X�޾�j���ooyl����!������iP��- f��`�H����5�]G���v^z���a�\�O��|;�m�I�,7�S�Y��Z}�<��E7;=3I�.&�g=��=�����gy�1T�騌ꊬR����˩.1�ٍ͈�gR�����l�wrQw��{��\���h�=�Z��r��v+��Al�/Mc���C��;�
fB�|���⧨-����
���2��ņ(aq
0�Ƅ�{����뽏N������4["'��cޫ{�_1�`��s�U��c���v箸�����Hhf�'=�Gy]�������QMr@{�}%}r����V=��x��y�u�T���J����+��
��%d�q�T�R�mY���E$.���>��C�L�{4g����]󂝣&k�(^M���ww���ur��b���q��<'g`h�~ۦd�ug�jC��7�����v�>��oY�+Z|�<���1b��I�O[�������ɏ�k;ŵì�^�oJ�Crz�������~����[�(��Lnxd8�X�S5���db��v�S����Vg���	�x��|:c���\��ޡeeHr9����r0K	P/�s�	��$�J��KIT�hm:QL)"�T��	z)h�p��Lȍ Ó��)V��2[���r ��2D�QfQA�YʲRȢ�J�APV��v�UZ��O2U��B�]�.EO#��+@��Å�ea%(�y�#��RN�ʹEЩM2��&��P���;�h�=\�Ad�<2�%���9�%F(���Qg.$�;�X�eHs�T���E&ʢ'E��B�Y3�w/H���I\��䜫���W
$�в�L]v^t��"t�5�NEG	̉P��&z�������Ң��(��
�@�P�8Dr�+����Vl�$�T���rp�aV�V�QdT]2*D�9%�8��"�(��;r�(���V�J�V����I��4�VD�u�;WΑ9�,3g""�d_�%h�%�kIK�Y��e�bEм���?���!l�fع����q�l�O=���ck4yۅ ���Gf�n���|��`�
7�0�Q��Si�����z��;jg	:�=�u'O3�U|���sO�8��wl���ݘ��g�v������Y�Y�f��竗v�6���rK��ֶ�;![ջ���.ѯ�ϟ6�i�]�@�Q��A, ��^3��k�nݠ��X�����!�&�dݮ�Վ�d�x�b�y��t>h�[��)��g�i��9u��q��\�Ͱ�+�>M�V{��-V��k�gN�^u�x�8�^���C*`xr<����-W���Lh޹f�v��tsk�z��;��v��mq����a�`.KO��Xڪ��c�cv(Vx:����Q�7.�)U��cv�5����[sa�n�&���ݞ3r&^��i�Z��f���[.�=zGL]hP�Ѣ�f8q�nג1�n����qДu��^�%��魅YLj�v�ă�4�f�	�򞺄s��d�-��<Qӳ�`�f6BNۄ86,����ͱ�<s��zۑ6�[����͎@�P����VJ9���r����Jt ǴS���s�3�[����Sv�\J����'�Vz�ns5��.5�E��=u��=��Jg��v����k+�`���)]�W��q��>���cfΎ����.�&xm�y�;��t���c��q�GC ��J�A�m��Dc��l�<m�f3�'�<���=��8�c�t�n�[f�˼���l��t��7n���a]�{5=�Nm��bz�Y��i;�%���� �+u���<�{\ݔ��U=vf9��in��J��3������������1�v�YkFh�c.�z�;!�,rd�����X}�Y�!r��D�p��V��S5�dXZö��Q����129���Xy�� v���;Gv��7��,�6Ce6�[�+�ѨN^L��f�D㰱���M�<j+:�۩/Fh\�-l7��n�i���ո֮�n�d��v:ݱʹ,�B�z�kSv�]]۶��g���1u�crO�,�0d&М�� �v����۶���A٣M���6�`�r:�7�7F�.�ݫ\��c�r��u\�Ϭ�s��0�9�������=d�������S���n���<�����koO�Sۣe	����˶8���O^��pm�vl�8��p��p����:�|����wO^�9����ٶ�8v������r�Q��x�������v�l��}�~o޷�|����h���k��'OL@$	ξH�WA�.������&ۧA�BAq���Ag(Թ"Iث��'�G^�INN8�9�҉������ܻ D<@�C��H����@"k�e�1%��&��j�$G�^I �u��Hx�b�m�˘��脍���jz&SVg��s���쐁&{�����u���-;�>&�d�������v��H"{6�I?*�gԁ��o$��H�L�m��[��<�����5LsC�1仼D9x��P�ą��=�;������Ӳ>'k�Δ��Ͻ��D;;��Ǹ��S��� �g{m wc��pbv`����	�@��ԁ��< �4�\�4��S�"��������i�T�s~78Wo{M�o�ЕY�v{mX^�[���7���'~����HQ�m��X�i�<�UQ|�w�!�&�UC�"�xA� �;��N�����vA�=�oheE��9X�\pv�1\;'~��$���H�V�J��x��o�$�˾JY� �ԑ�D���6C�自�S�o{���-���,'�y�� ��=N�w&�i|k�ZD��1t��ዘ��芯]Լ�$gN̠�U^�jSSC�W� O�ve��1�{/j�t��/K�Egfn�*��$�olt�k]�ve��f}]���vIN:�;�;ZWP�Y4��������}II�ʹ$��Q ��3Fp�:������RD�H񋼵�s��gB��D�b�!�nd�>�V[iDuj�vY��:	$���K����Q$�	B��W:�	q�=��b��i^-�:�>#s��$��-�}��Wג�{>�~W�lG��.$;���Q{�l{���������=M��V9	�j�.����1�#rT10�Iڎ�I2�$ H9��A�A��������Px���ݚxm=P�TѺ���\���N�(�H$%��#��9�8�ه/�� ɼ�މ'I�p4c臡�t� O��ݔN���.�JV=�̍�%A4���}+;�%��ob�l��hn����=l�+`��sɏ!����B�x�D��7Ge���=�ܱ���g�w0�D@w�F�K��u8�Y������0ѓ�Z�oɛ��N5�y'$��A����������g���ā�k��A�;����^����q��}��2�3*�Q@�.znDL��J�>����}N�ו�$Sn'�I�y/�ˑ������0a�W�uNt�S;�I��Ab�s�}9�� I����'��89eW�1U�vOT���|[�ԯ}ï��u��8S��[�l�Yk0���H���7��|;4"y��IK̨�����{���CG�
UE���׭�}
��igeM㋹&��_��Wܐ$��iVuj�<��m�&˹x��" 7/<n��w�uѮ:Ԙ�w,e��s˘�#�o�?�[}��v��˗����_�;���$�L}�iΤé�q���3�q �˾H��5��D@w�D�k����B!����3���H���  /������M�s��a�9����$�D�ȃ�f��/�)/K�m &��;��Z��ͤ�7y�����S�����hwx.!�yg�sBR;:d����"�tO��{�Q 	{���i�BDj{|Ŏn�/9�xDL��0�+Ŷ�ב�����ϣ/�WD���'���gR@י��sxX�-3�r�wɮp�tO�.����ܪ��˵a��{��*ߦ��Щ�����tƫ�t&���5��M��kE-(�x�7,ο�D=8o|3Rc0X��
2���C�����;�N*7I��8N�9:��W�;�;�v9�W]X����Z�Ƌ���vln��=OF�ٶ7�u�V6·\g����Ol�Wg�\R�Q���]�ݶ��gJ�ձE��lۋ˴Yܚv�n��s�c<�c�8MX�9��B�3/&��[���Ku��cn���N�u��<bs�Dr܏��k8�W����u�g��i�Ѻ�r��:�'=6뇧n�۩E��2]��FD*��O�\�_߾Q\������#9�A����g4�b*u	1�ԑ�&�Ag�#��������n+���I>&+�� �מi$ܚ�f�OB���Qu��^0��D<�k:�G���4��%7,�܆P�V���s ��R7��d��� �"�"2�So:̮s�][��H1��yH��'�V�M�1�d�>�$�u%�".��*c-$�ƃ2���F ,������
�n�ŰW\���I�O&@$�[|�xu�b���<�:x')B���k:�l롍�A���6�؞��1��W1�}��}}���q��0a�xڝH�@9��,A m_$q�U�U��]�x�w1�A�LA�耥TPIoz�۝������](΃;c��]	yU��X�8��ڞ��e�G�����ʡ���:��ۗ�ˬ�Чw��c�e��_H�ߍ�����7{��G���� <O�꿒�y�^D�k�#w�M{<ވ')�7Ab\<Dz��� ���D���Ӑh�h�/GGs�a~@1�Wg$H����Y��0s�6�j+{Y5ϣ�.z�T�#+g�x�wm[=H��Q�m���YH�W�{h��H��
� |�6�]j2���b{��I�SA<�1�H+�iyu��������#��$S4(�HA����m�Oe��l+��è9.��g3�e���}})�ӧw���o�D�H<�6Q��ڔ��X}�lZ�A �j�$Nv�� I��0a�A��D�G����*&g�I�"�n��|I[�I����h�D*b(��H�]�D43;J�K�$
��A��m��~��&����EW�h�a�+�?w�3��DnDh���L.�E3��2Z�}V�;��׎�z��Pd�;��r#�����6�1�H+{j��Q�GUJ��S-����+��$�r�D�	Y}IA>9�W�/��x�ڻO����Y��0s����@"H##�D���� N�W����K��	��"|r7�Ah�ӛ�g�ے��ǿ��c����#>8�۝無{�`�@+<��/[�oS�gf�4-�7�����7r��H�H+siI�� ��ۃ���@���w_$I �ͩC3���1��a�2DEr�%��	r�M��U\�������F�AvPۏlvZdLe�B��ı�
bDɇiE���$�63�	$��vq�EuS�xj�$�w�!㑽�G*`d�%�Cgt���'�)c������ݵR�$����A>ŷ��8�4����.�ֻ�%V"n T�a)���h�U~�{�ޑ�v"�jҤ�ǡ/귘���з��y��qܧ)͉��/l�i�L'�jOw����J$�@��}`^'� ,M<J}���� `��exWDt��=i;� ����� _��-����+��p����C�IpS����;]����⽸�$��
ۅ￾�x%�340�a��.�AA�$|N-�K��cNs�,��{�_.��#z$��{��pa��]���Aw�QS��9���'�� �qu��H+�f�9�=_�Zm� �{��1�[I�&$���Q �uft�I �7�������6{�&��$qm��%���^Dɇi@�T��0�Ğ��բ��`ڪd�@J�$A]�W3����!MLH'�&I�]�D1�wK%.H�B��JKVQ̍�v��G��d	�!-�H��R@8Y���(�.K�TM�sm甩Hk5�!��eJn��������4��)�������h��/������ʵ��"�w��ň뿮ۢټn�%�	Rv�Ms�f}]��=z�����yыX�r]�
����R�3�p�h����>L�����ɷV��-�ѹz������$vq���=/E�\�nN�_l;x��BpsU����.�N;ۧ�7W=@@'gs��c0uĦ�Q���
�<c<Q��੎x�ѷ�Ι�ܗ����:�	�wn�ml>���#�����3�6�;]���9˺�i�#rpnć)�G�g/�_�Ƀ�bi�_�E<�����$�=�R���J`lc��f�� ��� ���H��q�f���:^�u/"	cs�c�")`�͑$9���$���Ay���q��n�Vt��|�1	�۸0��.���HI�ͩ@<�'j�g�4���A{���#0�!ݢ!ɀ�R�":��{�E4i��"z�%x�	�Ԑ�3x������ous)�������@�/+��%���O"D˼�n���IfOL��8�.�GT��}�}�w��W�K�O�l�Ihܦ��}Co����|�θ���	�zV�&�p��F�݇�iz�sU���-K��}~��o͒�4/��ĵ }5�H"$���'V�m<��.�ԉ$��H��
������;�j��$��]��4"��|$��G�s�s���m���2��	u�囂$���z?��=Ź%��ˏ������0Nô�{w��8� 9��l������[�xH�ݩD�Nl�y��ep�{����������T���q�A��K6����As6�r9L���g
��P$�4�u�	'nz$�ìBr��I��d���(B���e���skĚȮH�|ޞ��;��#u5r�����;��z��wh���`<�jD�L��J;y���&*�h���w' I"{o�񦠌��f��j �0�pa�C�%�����c�����Wl�델m�6d���_|q����2�<UOH��$��o�屜��;^CP��׹� |I���'�1�p�h����\�&�����F���}w;	�:��"L�˶ml�1^���,�Z����w� �����H<�vQ>$�����^�o���������f�!���;�^m�u`f[��yn/i��~�Wy"fnQ7%BC����8�k/��k���M\C'fsZu�>#�וb��pN���&{Z<z�;�;�o�6Zx�9�Ʒ|'f�2�񽽼k�;�P�Ǟ�w{qw��u_|JnW��������ң�BŃ��q
C���!���hw����#��Ɍ/y��Z���<Op�?2R����{������&'��4�QI6@�����7=2Kv)��C,��z�ҝ�������~�v�U�,�z׽�[�߽}K�]RƄ�\����r��-���8zxh ���qxS�ȵ�*��OI}�ot;�چnqŃ*��,EΥ��9d�>�s�}<;�k@Vi�s�׽�w��9�߆9��ċv�K�پz��9]Զrʁ�{p��5 w�h&{�_�~���~k���x�_h�E�����]/������1kJzv�_n�۸p٨n^��>Ý�V�,=���.÷�>��@̆;�яR���}�q}��'n����{�ܫs��źx�u�c��A��ɳ=�!v�{�j���ߔ��Jg�����r�r��y�1d�I���˞��y��9�_%1+Y��b����9!�}�v��Wg�/f菷�����)�g:]�9���}�a�U(��V�o&�*�����ߌˏL��:�o�ӥ����|<nn��{ٰ�7�s��r��\f�=�+`g���;�b��]Ke#�(x�%K5�~���[���|�1�3�"''Y}�%�FS�d3X;��I�~��L������ɾ�Cc���:���w�I�RE�	6A��y@���R��G(�+2
�u��
ud^�a�Q̑~Gp�2"(�SN�LB#X&�t>r��U�,B�J�,+*LV�r(�J��JP]�Ut(*������g�fSBV�T�eʴ��
i�IK�Pz���֓��Z���ᚔSB-y���K4وVJ!U$Df��ʐ�\N�2yЎr�,���9P��#Q�&*�0����f�X�"�gybEQW��'�G:U�&����T�,��H�.A2�QW#����Qb�S(�YFWSXg��]dQ�Q��%4�:HDE�s���$lŅG*:r՜�d�Eb��Y�g"!Z����B5
yNN��Y����.I��C�Q�uL@�#��UDDE���(3D�W*�W��jEʧ'9xt�@��΅���QW����16EȈ�L;$x�1�f<��_*C�/��I-���뷀Z4;p�/k��5�j�xa���#�zȐE*��I����3gvY��._}��:'Ĉ�b�\0�A��d�eu ��ͤRh�}�r؉ �%#�w$I �v�Z�u��n텇�ͦ{#�\����p=�0]cd��r@�qfNw\���j�0�r���}�o���.�6��='��mnl�	 ��Ix�ݻ�Q�x��H$W�(#7S���O"D˼��Sh"muul�卅hI$�9gbD�1������*����tH$

��6ļ��]��"I+���$���-����:���'Q��W|� ���H��l�C@0�@��y,:�r�6�Y�����x�I����$�m��rq��fI�w7TȻ�d��*�F����_=�y�C��u �+�x`�Bmؽ
R��PM�f�O��#c>��Q���-a؈<<�s�R�H8~�w�e��ۛ�b;�u 	 �f{��GM��Q�~8x�!��q����T �˲ݷg����-��k+�g�8�O=������x.�h0��!���ƃ ��,�ݕ��$Gf��<�<y���
�,�p���S�>�ޥ���l������/=jD�#�����1K�ΟE^T�zq�vp�ݱ���w�����r!<�3.�(��0Ë�"8*z����wi7�y�A�~�>$[l�ω�Ldb^��@�Y�{y�W&r�^a��{�2I>��ǒI�m�,���xjƊYx�L���2�GbEk�.��<3�x�Tt����oe���6<m�1�V��'��:�	'v���7E�bѫbf7SG���{t�����WB��,�7�|�������vp�]�.�3h���Č:q�O���0Y��޹HJ�/9S���ûc�=;���Ʒ��n�٭g�֎6�{p��&�#Ϲy��lo�mgr�ff/:��^t7'Z<�������r�OD.��f޻ 7�Ko���"��y�{Zy��!��&�qƜ=xM���՚�{3��Gnţ퍜��{М���^���s��q� �j;kq�\]�m�m�q\�g8�=�s�0��FM��lF`{�^���x�28b��x�ǲ��Ń�Ǆu�ɟk�3�˺g!���������|���79��$;;"�۾H�������A|�ԁ �ͳ�>&3X�S�0v�Av�UuF�S4&0������k�yv����-æ��M�V��A�˴C�v."��ܙA'3/�@'����A�g�?`���9��w�Vn�&�OL˼�[�s����C��*��ٛןH˻ļX�]�m�\���T�}�yr���E��Ji@���ۧ��IU�h#S��#ڻ��t8�l$.��"Iwm�Dd���nZE�w��8ڶn; ̝�w����Έ�m��ud�X'a�w��1f�L�"���5������>��{(�A+��H�@��B߬D;c���ZA�/��^�C���79Լ�+d��z�4��,�G��,u�cV8�j� h���;|v��M���{C��+��6�ЗL5al�;�gr��	�b"a�ǟ��fq�'�{a�$n���V�Z�#�1s�I���Dճ5�x��G��%=�H"J��H��n�b�/��m7�u�b@��:�"�ք�����_��&����:���h������n�@�9�9�+��2m�3A>���';e���"%�I�w��-�Z�$3�1���2�Z��/�4�$,��3�����iw��X���]�3P1pm�g����/O��(��ɳ���hۀ:���ٞ<P��]��9���q���� ���ܤI��<��y�^�9�u�z"6���$H$ۘ�@\��]�4Ax��A�� �u��dP$�׸��c��A ��QՍ5W@�땼��������$A ���|H(i�a�њ�ّR�1�qX���MF:�5��%��-���g�tae�M\��͐��-AD����+�<
F+�'�_n�.��r`�xd%b�xz�p�Ρ�;� �5ے�&;z$/Ӻ͹�3�G��U{V�#(�܉��>8��	&*�$���1hA'�b���A~��#8ք����$Er��l�J�y�/S:)�SX,b��I��$�Or@�e��w�����|ƻHk�q�^��1�A�X�s�G=�b3�K��u-�F,��~�~�M�N��;|���-�:�@���>�	�+'� f��t��*�;���jHK��	�%��g,����x��4�D����ȓ�K��I$����v9� �hf�T�鰞�k<8fx�W�u�H9��!x�]ŵ��3���5�\�S���]Y��/�Q���6�`~�hR=�|Fe�� �Z�D�.�xnk-�Vl�ϒ�N�-�����z`��۩�Nàg�#�{�w���n8�o�~�țvl�����.��=γ��Wp%N�6d��ݚ=E�S���yf�\���;fs����$�B�\�>'Ǘv%;�Y�b�Ő�9��`0"gx���t��wǧ�E�Ѳ��ls��T�tX���X�� �h�#�z���b�@�H'ڻ��̲Z[m���͓)l	�#z�$kH"�����;���2�6i�zA�A7`�6D��I�ŉO���Ax��q�م?D�:'Q~rAg�Awf��mV�H'��f �$�n�uעY�T�����I .� A��݉<	�6����h�wY�S�-��Wi ��ԯ�6srQ�s�Zw8Ý:��N��	��ۈ�L�A"��r:������_�3lTL����X����m�R^ ���H	ۜ�ok�Q>�+�t���\V�⿑x}
fh����N�Y�0]�T��|/��U,�TlK��c;U�g�u:*�2f�X18�­��]�{���Yq���$2��ֺ8-�^��Ϲۍ�5��wW�y9�ֶȓ�GH�Ml=vstt�]fZN���u�țu�u����S=n|]������T�b��x��j������C�auÓ�#m��=m卸ϵ���6����鋣��N��{V�q�l��y�N9�-�#�cs�&�=�`�,Fu���Rq{n�F�u�@Ui�,���u�ڮt���;�;�Z���_h�-ˮ�3;z���x���������1z���ߛ[H"6sq A ;nsɾ�gڦ�h�olԩ��$���A^Ѓ4�@gq	G�Ȃ�a1�2��nt�7�ā�;9��dU����i"
y��y:��
���.�N��$7�0	�8ju�v��o1��-�H=7��>.{9��*Nñ�%��S:�8m�(�q�r��'���R��C�o<�b�9T����Ԑ��!��x�"�oO��|s�l�*ц:���n���95z�����	_.Hܾ�M,�΋�K�.u~8gĆ6e<7���/e����N�=���h�Y�D��������n�n�?p1�Ԃ>$=�"3��$�Y��DCvSV	�K:�A�C�n��ӍX���A�Kػi I��Ec��^��
�ֵ�$E���ʗ	��l��ǘ�XR��ww��`�r�`/8��K��OeVRzd�j˼�ݽ���������!�~��/����eּ�/�d��z
 ���! h��� �]"�h�d������H.v���](�gY���u"%�P<�:�y���8��WL	�^.H�OWv6��r�uů��o�J�x�bD%��\��>'ƫ�N��B���s��Mُ �Vjԉ��we��?Ma��Hޓ��\���d��T+���ţ�6�]���ݝ��%7g�K\06x�A�@x��r�$A ��{�eI$uwbG��er��k�y'Ċ���c�9.Hw��<�ٛ;T��`��L�Ax�$e�Ĉ'k�^��nwr;]�>eS�"(��f1�G��(��8I'�7 �Q��hghfm��=$�Ie�54J�����nOh���:���j��S%O>�wN��y�!�<�⸐�;J��Dv{"�,��\C[۔�����"�/#�݉�m�@- �Ec��������I���`�˳�]�(�@v�瀞�Zom�"/���)���R��uj��<���z{o�:�}x��;�w*0=[�����G�Ah]e5�1�B�#���;���Qҋ,0jw+ؼ��Y^���U�mV����������v=�RZ��Vn$I ���� �Di˾��7F�@�GV�$|�$6���%���.�9��)Ȃ�Iz�8	�*�1 AϜ�Knأ�"�.z���$L�5C���Axt��_m �'��g�r	2����'��7(��	����	>~|����b���z4�.�P�L_s|�@,��GĞ�k��� �VB�v!�"ْyć���Q]
n�ҧpD`�Y� Ż_h(<���x����Ҽ��N/y���z/�@eE�9���ݔsdQ�W�	D�A�m�A- �;��B��,8 ���E�#I�[�bd��N��V֤IznƟ|�W%�s]����6�8��AxLXX_�+2W0�gqi�:����u�p�wkۆ�&����_߿�Zq?�!�]�����=�t��$���x��f�<��UF3��@�7��$��;6�Aw�$���:�$I|��wd��witΒO��0ψ>W˒ �{���쨫�|� �Ē�	���}��$ful��3,'f�[��f�^��� ��ky�����0�"��o��ٽ��#W�'2_�1�B���$�˻(P��f&ʜNoD��Lކ/��9a��,�H�G,�AcNnTH�c���I���H�A�݈(G�����z*s�dVv�"����({;�"��<�.���,b�"~܋���!�wF͸'!D�;�m����7�rs��]lY��9��X,
�o�'��,�}V{u%i/�J�P��&��ɣA�*�7��(�O)��{h��ȩ���A��خY�&`��d6ݲ�e�}�K�!��T�ٻtѳ���ݷ�}w�1���K�<<����}ڛ��y��o;&��=�TN��}$ש[�3�z����3\��^�{�{ ���{}:4�S}�0��8s<�Ǘ��x�����c�g�l�L�q�� ~�2ף13�1�پܓV�C/y��^�<kߎ�0u<�ƻ�}G��M�
c�ݹ�m��1���l�|�޹��{E�*=��_)zo�{�ˏt��B��)��-�Nt@�N�۞	�[�����⻫������\��Ż�wش���};z����Y���s�yޅz"ǧ/#�U	�wA�0����%�pPX]�g�Ӫ����ݽ�=/x��8�~��Sw��-g�[�l��$�w�����j�������p\_5��
Q/�ŏ�>�a�͏w�׸R��y%��h���h�2��Sc�t��GL��vO��:�����s��g�P{+�`��e��3N���!���Z�/[9@>`���Ӿ�v�{���P�ξ�^�N���f{�/7�²���=q�u�.�ONڻ׽�|�Vxnh7�=�<n��]�0(�Kk�pt�UD��z�G���ި��s�����ެ��I��ϴxiYNVqʜ�,��Z3n���̈́5�,�V<#�?%��DPЈ��L"8\��P �eE�*E(�)j�G#�Jr���-N\�+���8hh�!ʹĒ�*�s��(�V�L�r��AYI'-U4呠\�DΔBM�uf�Q·B���H��FR�(��M�L��	ӄAEL�����B+3�@�p�?�r.N��2��T�2�镛xܒ��s �r��9]�"�aeR!E�HUX��W�f\�\"�����WQ�+��r��Q�h���� �"�����hERAM#KL.vEL���ʋ��\����ʳ��8�����|�E�T��3Cͦ�Y�'y�9�edAW.\�Q	�Qʈ�Ȉ��@��ԨU���EI� �r���r��9E������h*��*��MJ25�\�*�#3�\���d��#���[z�F�[����m��gM{<�����h�B�}�]�������7Y�:z�e�rrY�v,�(4�"{ ��[,��d��Onta��'�t����{S��p��toWe���b{-kq�>:�8��݁�m����n�u�aLu����g��y�������95�׮�X���]`��36r�k9�n�w�ۍa���7N&Zx�Y<�{U�u��s��3۔�=t�,�.q�m�q�����<A=�`���]&uٮ7<2s��<��wh�Y�}Ռ�M�`'q�����D�\���:ծ���M�vE}VZ�7�\��W�D+q����a��n�rd�۰l=�N_7]#����#��ݸ5�鰯kc�r��s�6��M�/I�#N6��a��k������}1v7G"u����������r��ݙ{q�4����\N���l'q�k��cp�rGkbD���q�c�n�b`w^��t�v����%�ʺ�n(��Q��x�v/Z1�^Il���F�W={EF�i9�^y�GH��]j���ȴ�q��d�
�ރ���m^�X�#��V�]���b}�A��p]��G.7s�YF{uΕ��v�8$�&�[�{NX��1ҽ;\��ݯB\p�ݚ��X9�x���m��w*����7lJ.ݼ�od�쨄���v�vaܞ���qq�m��l���۞)����bļq�h�d9�u	C�:�!��s�6�uc<"+r�e�m�����po)�����؆�6Dd�dI��B�tg��qε���͗�l='&Ě{;��a7Ty��Ӷ�*��urb�X��;������`�5G<���;p3�̯;��G�u���-mս%�A�����3���,\.;N��-�({z�Mu��mg�N,��G����v�G/:��/!�Ql�������I���kwj�p��r�0	��y�Oj7��ۃuWf�c�����+�:�-հ䬷>��{4�N8���h����$1��Nh�g�v{����e�3�
�ey�i��+�>3n���&��kA*�9�}C�T�F'#����8�S,Y��y;9���N�tW\$H�WX=f���Y&N���j�3�#�6)�y�qoc�����	>���������A�ˎ�u�ɇ���n79�x<n�$�[������]���6����h�v��V�B�-�wZ�{ c��e0xt��G%۝�+��lݹ�s�������m;����x��̆ og6Q> �Wv �ѻ�����#rsR&o�Y���:�2�+Ǟ�W����!��m��$��l�A>:��/<�b��r�5Ӝo�������x�L;��9+P^$]ؼ�$ϪFt���-�d�HU=�	:��^$��M�10����]k�V����Z�w$�oT��|H՝�A!�c�,�OɁ#qZH��k�,�?�0���J�%�_L��B�����"o��q'�Wn$	���bC���Ű,�kL��eM���l�����s�k�ěF�;F���cp��q�.&D�M"�q�w|B���UP�(�\�7���H�O���3�V]�LJۜkz�H�	��9��� �p���!#]o2>c/�z;M��&X\�{*�p�4��OW��a���_˝��f��V��n����z��*a�$��'�34�[&��5[,����p�A"�s>��Ikz=DD��*n�1ܼf�(ujn�<�n!Orv�#�0���g�Y&��@�_���$t���"�w)Lj�}�obN
ؓ:�ץ7�&)�ZA�0����wL�h#�&�y��	׆&p�r��A�͙=��!s�ł\�%�H$�vĂ|HY=�X7V�x�l���w�K�Yru�y���Ž��؋��6���tjNP�3�h,b/o�a�?��}�mfԠ	!�v} �N�^�3TA�s٩O���	�i*��s�D!�:�$h3�9��p��Ý�r�$�MF�H$���^ڈ�a����B�"/)��ó���w2$�7':Q�f�=��33���]���V"e��1�dC��Q�!6�s��{q4iE���9m��&��_jŏe���O��ma�[���Ml�I$�.���f�fgx���y�i��S|�o�9K���$��S�>$��������uG��#5�7�35O�N�w�a;���`�vܝݐ7��2'�&$rv�"@$���I�3��/\!�Z����j�a݋�� s��nu�u�Wkq�G�����5���𿝁����}�.��}kwe	 /�m e�1�M�=�^R�$��o7�ָ���a�]����bM�X!.ݔI ���	n��4�H�WV�(��m`&!�ȇ"2Bo������H���(�ڞ��֔i$�Uz���ݵ+ٔ�B��a��B^!u�;w�u�)�� �J:W��9�IIΞ�q�����઴��z��A�P�j��fOϭj�����>ɉ�6�[��ۛߚc���y��O�Su����������"��,*;�'�{8� Ov�fw�Yʘ/2�(�T�D�7'��37��q� eF�@�D�u$	��&���6*oQ/'cΞ8�Ookv4�a�g��Mێ��y�=pb^.0�(p���ot;<;�����=%�/f��A>$�OD������<*�by"	��n���4A,"#j:d�����e���UM�^-=�I�Nl�O��4��O�fns�3?�� ��H�;>� �J���כ�� �v��@���$��qX0���!ȃ�W�U)��L{�-�h�� ��r$�g�y�t�z���FVՠ�mЁ�\;vw�ɂ�R'�u�(O����3�=l����W=$�[����[�֤�и�wdI�1�a�#�R������|������>c�f��U�����[}ڷ�ۻ%CI:<�k�� ���%i݋{��ñ�C�.Ν�c\�-nM���=�Z�jk��흗���+��`Z��Ԝa�؞���I=H����3���\<)u�;9T��+)�r���\����P�gn��7K�dܤ������h��x�4\��݋�7��آ]���z:��Ճ��_v��ɝ��֨�9�r�ְw:�gm���p�����w��v���-�8u�+��{Q�m�b�wRv�%n�IW�����3����c7��t�:]�3����Y���]��eN�$�;'���2���K�Im��^�t�O��M�g�q;����%�@5�򐨦]x�GĒ��I ���@�Z󺫄^NG���M�EUU@*��ڍ���v�	�v������C���A'c:��J��5��Y��Hxq����4���	nvD�A��ļI �w]8��;R�H�D�4���b"��Y�i/��ptm�%*�	�<�؍6��t?�TTH D�g%�	}�~��6�j�_-�C%� xg��3a��3�H��[�h��
�P5Ny%|z�bb��}q��\;vw��ّ'�E�l�A1��!�N�+m�es�����I�}�x��ډg0�S�]�Q�gc�ݣ*���w�źu��w���s��^�mWPמ6�>��3�\4]'�a��P�K_��X��Ե]�Os[}(4�,�@6��7��%.�	 ¾�D�z;�y�k�4rJ�����}4]�ecM���S���>��
���Ж\��}�;{��	'їڂ$��^�<M�KD��f	֮ᒄ�MdgW�\�d�@'�"��"C��4�*��%�rn��g����hr�0�/}���$�7l�Y��@�/�jf���o��P �j/�y�_��+,k�1jȞx��������TTLIAطm�9��.��%�p�f�n��m�S����#��������.C��`� d^WA$����A��j��9W��3�#wR��z{-}����(.��ó���t�2���[_�&�j���$�}S�k�h�-$�;�̭�݋��%�}� ��L��&�K�2o�>�t�ω0��$>�sռ����w�r�oi�C:�%뇙#o�s�xn�?��:~������7K��t�(��`� �G_tHe�z�7Z�ܧ����bܹ�Ύ2Iٲ]�C�3�f�؞�͐�F�S�ۉ	z��>$�[�Z:�#�N���x�^D<N��KD��X�%��˚A ��l�Nf�F0�b�������$��1��.v� ^��V�~��C���#���%�Cg1�=rn5n�x��y�{n3��"��;[����������?��̒�Cw����\E��!Wl:-ޤ��HC��4�_�W��Ap���e�R3�Р{;eߍ>4"��I�>||ƒ�_%�Im�OK��gSUn*�A��ػvw��m�r'f�A�*�v\�*뾝�|HWd�E�_$
��KA�.�2��\�<�7�m��u��7�E�HbA9z� �z��/��gf���Σ,���U�d5CMū5�\n�c[�L�l'7��5iUYJ�����T�]�>^S���z�'|Tp�Kۻ��s�<��yyw�u��M�V�n��<�p$Ft# ��zp�x0!�ܳ$)\�>$�wR<�Zx���`�6v0ω�,����Ig>`�쮛	�/�(c��wO=#��l�\�nd��ѷ-�N٤�7m�۶ӛ���������lV�������:d�oWl�I���A�࢈�k���7��2O�X� �qՅ�9K�q"���HT�^W6��so_����+Ԉ ��AAU�UGj-�Q|_11��fҽ9�h H=Y��!y��4j�O�NoM��Ex�~f�[�x�:��}yc\�D9.���$W<�4�g}�#_.�x�	9]�(|����M�X�T�4OV۽5���|g"a�1we!�&��S��H/��!�45�q��u0��������"2��	/o��J�I�{��В�,��q!�Sx��Ĩ카��pm����1�y}�wҴ����6��c�����jw��+��@���w�ܮ��]��]aw5����0H��˹YuH�la����ӌ�C\���u��T��a.��V#[;<�'d���ɳt�\�C�۞��3Zg��:wWl���#�Gk�["�n�g�qlf{8�v���۷�C�7n�5���!e�����n���r�#{v�o^��5�k����)��'n;{w��k=vv�m�.K������'��71��ti�=1�ul���Aȃxz)�i�v�b@���J{�̌D�R��$��]߯�ƫ6�$���a�;�1�#q37#�	7��d'��aM�����������h�����ex�H9}Q����A ��~��;m ��x.i%��k��遅�#� �a�S���&i��4��k2�	����)�����d���3�����804���$����m ��uʧ5�}����o��z�ht4�a��B�"�s�N�WJ�x963�\KE�wə$���i:�� tz7�qNީ���ܨ<ETЂ"��(Q
e۠.��yMc�ggu]��;hv�`��b��{.����4	 ���$��ml��
Y\��壷�\T	'��ݴ���c�xjU3DJ�[zӊ���Z���^��lݝ*#���3�t����e���Fw�sC+N5T�
�+f����܉�I���,�m�D���>�ec��I$���$����H�H��/�آ�<d���:�3����"��7T�$�ul��M6)�����će��I[\���P���0�"��6��wI��^o1��ד�ĂG\W$I'{���F��ѽz7���U����n���Y��2S���'ăٷ>�n�^o)�u
5�gV�	V��c��'��76��M�+p� ���3�-�G��d�8��p���g�1��rwhEsn�ۉW����]�w�t�قO��-��A��s%�`�%���I ��\���LJ�&\ڒ����>7�-Z|��M̒�6�%�3�H�Ų�'ă�� O��{���;�[�q�"x��������2C%-H	��D�|u��o����-�fh�,X��4���~�M�I79��^�V��ͱ�I���<����p����(��5��7Lk~��l���Y�ydJ��"�����L���8�n���w�f-G���-�=�;=�����g�
�~�2x9f���׺�7�ḳgx�<[��vs(��:�{G��v�t{�=eng{r��P��F�u)��b9X��ʵ(4�`Dd:(3�^^���3vh�{:�������;�A�W{��	5ryh���iW�8�w�f�P^��������cڄz�p��o�Kho�7���OvwY=�0M�6og�9�ɭu�e���7������'���^Z�h{4N8�\���gw�ě��!/YX���f�N>Щ��8<��$xn=����1��|i<��[�N����{����otAx��i�};���rNX�|3ݽo/}LK�%J�����w�C�Ϳo1��a�?e��g���c3�sV�=�8�-�̲����q���G;����˞��]^�4aI�2��^S}�X�w�I���������O�ƕ�{waў�zx��`����<5�A�wi���wr�C0�7DY}z[�F/���ٽ�}9q[��>۫�=�#�{R����0�ݾk^������$T��l�L��>��|�u��s��=ǧ��/;M��5w����K�km��ςc�{�쳸d�+Z�˖�x��eغ���RϤ<��K!:U���,���ӻ�[�C�H��YId���͞�ӯb7.e�y����xEW�{�UD/��� "t8L�����ap�����0���UL���Qa�hh��B�N�H�*�EZ
-1h�&.�W��W�!9P_�(L�U�R��D˜��:�VBQ!�U3�9!E*\�P��hgJ�g9IҒH���#�XqH�!�x�0����r$����yE2��9QZ���K�Ы�E�+��,J�ZȠ�(9t���:y9ed�T_ ����&3��g2��GD��(.r��꜈�"����Y� D��g9\��(��iI�:�E\Q	$�.�Dr֙��r�眯[C�#�Es�s�9Ur(�*s.�$�^vㄇ�y�nO�G"�"�/ERp��A�dL���i�S$�)+�Dp��<l>$+�\�9ϔi���UQ��
MHs���(�������<w8s�|.K�L�p�"�s��yNl�8r���\��8Y�������rj�|� �{`�!�D@-	=���E�ࡶbz� ��t�	/�ٽs ��W?��|�%b\�v����C�a!�Nt邏�毦.x�z�y�
�8A"��A|n��H'��|�����R�j�+��BL�CX`�a�,�MS��������o�=r��{�6�)������v�l�<��K��Gf��'Ļu��(_
�;���b�O,H�wz�M]q.�1�.H�v(.�`�Y|���5ц�rh�wr�|H�u� �n�y��1Vr0���y�0e�;2I�sۮ$軋���=�t �e���n�q#d�e�c��,�J�Tϭ�j�@/4�@$��$��\��n=��S`��+2<�a& �R�zl�낍[�ts�.�;��z>'p^���K�҉���y픉��M�{��$��R�.�3����`�ur�$[�;�
�x��C<��Z,{j`����!�*+1��bC\\ω��<��v�r�ƣQv��t�ﾃ�c�/��~�"�j����ٞ㍧��^N�ZiU��,�t��������!��Y�@�	.j�@��IZ� nv�l����I���b`��
Bs���bf�q6gOM�$C�_<�I]\�%��7-���2�U�X.���.H�.a#EGH�	=�]!a(�j�y�b�<Av]�>#ioJ$*�F��'��P�v�y�ӊ���0|H7k�W�>;�wv0)c2��QB�"�����������@D���D�k��L�w��R��� �3>[��o'<O�{�e�ҋ�/�LGXf�"V������<Hl/��cd�E,�g���RY���}v̈́m݇l��z�a�}�uWj�_Ɨ��#w�
A�X��+M�:5lg�[�&��\&��+֮�W��ͪ^�l�ƍb�ة9���{yL2V��K�Jv��=���n�"�N�3�1st<K�0�*=ʘ�i׷=�v�)�AmӞ��6���m���nݎ���A8)�s�ݹ�I�Y���N.���;�wcvu�ўj�d����0&�on����욮��60>�q��0=�-�[�)�.�9l�l��n�`�ެ�bum�wg�㮔+�mv���??����DD����7�0I�7�rP$�O��2���矧Fh�5�ē��&w��wp�ȇ�SWuB{�e�e�c�r ���WҼ	#��e�X�m'�؉\�ot�|�`C�ř�;�IOf�H$w�`0���Xs)��쐼H;��v�Aش9ba˘��4��30�T��	�=���'6�$|K[�6E�@��'z;c��mj^$��A��.��;Cȑ�f�$��Ο;ܜ#�ʼH������ �����&�w5R��	�#w�<q� ��S��N��:=��x�6p;�Ӏ���T�Uw������D����J2�d�Z۹�������ދ{�#6��@�g6��)�Ȃ	�UT�������>��R�7��,zw7�ԥf��Kf��`�I�>�Yּ�7���}�W�=�t�4={��#�瞙��L�Y����A����F��X�
�$��q�#��9Ւ'�<�=��I ��֙߬�d��7��rsNL�)L©T7�<������ZQ$��=:`4��O�]d�>-�6��%�_@��DA�����M1>�v��`�uϬ��>*yO��A>k~�	')o$��� D�s�	9u�>����f�!�9sT�E� �{t���t76��X>T�g�Ǯi�3 Z�t��u�u0^ �����nө�����N��":+�v�������N9n�E
���	�s6cʦ��&��V�c��ڒ	��d8$�urOZ�WAЙaF�쾙����I���^��3�t��@�o�';4gc�$�[���H��֟�+�=��rA�c*}�J�� MQx�.�	杗$�ά��o/�(A�y�Zh ��.��Qk"e��Cb$�+�z=�����g�J=�Wq/f��+���	Ǥz_?��9�Vi�L5Y�Rh�J�Ɛ*Wq$���Iy��D+��c�L�*d
���쮣U�0�^� ��&�	$��H�A�6��.f�����i/4.DY����H|{+g�I�t��V	���A���]>�a^�!��'Eow��݅ulTip��n�(;Anh��� ��R�Ԩxv��&/�����pF�1������\��سeA$�z�d��H1}��f>&�I>�Y��hB�)�D�[s!��Zّ�
�1��\�|MZ�Ax��]�Hs{Fu��f���̆�m���٠3�b%��x�MutI �^ӿ�O�j��S`�^+ļI ��S=� ����I�����|�Ⱦ��z��w]6<H�3.�dI 5��u�vۮG���}9\����D{Ո,:k�v� �cFA`���/��Uk(fX�i����yՒݛ�[�ǯd�BHVp��q�^����� ���e%��N1P�<��Q
���L͋�G�%='s��緒$�y[I�[�0���m���ͻ�C������I���p�sWN��Ưn�a�I��m�g�r�b�������筭����O�7+fI��i��|�Oݲ�Q[a�m�A �VϦ�视���Mɤ��m3�O|��:	$��Y2Ao���AV�5[8�+��v6!ዲ���J<�bE�������4ٯ�ޓu�^"��g��k� ���ݠ3�b*��ы����݌�h��I�4�#��.�94�����,z�g���<CC��a�CO��]�,e7<a!�6d	�}>�]��=��u�e�&�ڠ�I�Z&9�ʬ�m��ݱj�ܼ+���+ dq x.��rm�����_P�JW�V}����m��?"���I�.Sݧ��e�ٹ���E4 ���q���ogh�ݐ��y*�ͦ�`�vۋ�Ykb�=�u�yƹ�v��nd�x����W��Ƽ���ye�.��5�Wc��������a��.��/A��l�ss�Ŷzx�wi6,%���ead���n�7�y�u6�����cnq�<��oK�v�ڭ��C.� ���ZS��n9MԬ���	�m��F�G��=��=[o���X���o-�J�����{fv��EL��Q�$��$���IKy OhM���w��Ϗ�.8�/:6�q�-�3��'&HS]ƺ�%7'�'Ā�ѥ&]w$	�f�F�D������gZ#K�I �ŝ(I�SZ/0�W--���$���"I�u.��(.9��Dq�xi���v���*ȫ�5�D���'Ă@$g-�'�{��Jgx�Ά�^ϧ�[y����Ad�b�"A ��Ȗ�M��	�-�
����{��vͬ�?�������a���������Z[������j�:ճvɶ��<���7������
C���c�>'ƹvJ�$�}��2�FW��]3��O�k+��I$��L�c�C;9�vv� z�L�GV�w�:}C�b���[їy,��X@Yڙ���VL9@$x�`�|O����7D�V�
�vF��ӹb��٭k&�fjX��S!��_5�v>�QĪY���'�Nف����ˇZp5t��ü:^�Τ���KMP��|�*V���2Q>$�u�������4�iK�Hh�[;	���=�}(�I�s �^߹�"3�����G^�H $_`A����D�gkg�|I}k�]*��̪@$y��<�;2d	��y��`y�����;��ֳ�	h04�W]�v[����n��u���wEr��\���������~�Y�rwF�jDr�`O������N�뮿X�C�H囩7w�2��ŢC��Z9�ک�.Ɠ�3_�u�dQױ �Z�8��-�Tu�Sڝ�B������×q!��ꞑ$�φ|D�ԭ�ϟ���`�@��9)۞����
	�4W���{°07�|$krf�3�^����\�����7�Ӕ��|ޫ"�����u6�c3G+o�A-z�d���g&����Υ��wMK,�C�L�%���}D���TfkUA|���� Ī�I�b��v0�C��H��DI�YҀ3�P&X�쩟Z�8�$���#�:�$bw�x�b��"!�bb���<A��Q�TX'�P6Չ�O`஡��_]�|p<C���!�O b��I��,�r�s��E>�m=<ڽ�[zfA-X�d�%��vw�0!�,����/O�����t��_jI>��q�	��Ž(���{�+eh|�#q�L�7Ėh����!"�/�I�]��>'�p�;����U�,� I$���/m�Dg��q���Sa���x�r���|N��Af<��ޚ�����|9g�2Y��̵>����ˋW!X����v������v��Q}<9��/k�꫊�^�7i��dN;?	)KِK�<�b4y��g�Ht�R��ض{i����=Y�FDy��+��>��e�d�۪y���w����n�j8�>n���Onx��i�ۓ<7���rv�t�ŶnΑq�����:������]KM�͔��s=��J���
�$�U9�/H�҃�;D��D�c��O���>���C%V!9�¹�X�H�ɼK�u��e�>p24V��)�0����#��I��O��ڧ��X�8�$fM�@���2f{b����T��PVN��^�Uɻҏ,j�J$}y�2O�!�#�h����︫$n����w=Dg�@xt�]�$�>H�3An�=1�He	%�a�=:,`HV�,��jO���8�ݐ/Z���"
"���$PW���YR�� l�M��o��������zy;��`�����#1EcV1cV1kGc���EcV0EcW
6��ѥV�AX�s�l��
�&6�M���e�X��AX�E�X�Q��V=�յE�%�����c;lv��C���h�E�Q�PX�E�X��X��TX�E�X��E�X�E�TX�E�PX�E�X��X�E�F0c0A#� �V���8���O���K�H1�`&��
���`h���c�ѫ?V�0�6{��'����ﵟv�?
{��`�3���������i��5����{?�N���f/�w�
"��ǿ�'ə�?�� EvxH�(�Ā�?o�!��$��O<]����x?��ؙ�({T^���<��qoq�@�)��'���W�V���.-CR��[-��6uChsJ��Ȁ�
�JGP>����Ã
 0"��Uh�@B#@B!@B ���P¡��ò����>b� ���"� Ƞ3��6��,h: }����1_�h�1�,�������;�b@Q�t
u/i���t�� r��I4v�kC�
m.;��K���M,4;�;29&�DW�b�㩄��6����5�$a�؛ ��+�@Q���(��3���2���+�P5#(V��b�DQ�@h��8�Idۈ9BeB�� �B�>Y��F��5�8� d@*���+mc���yp�-��@Q��V
nk@9�?Yǎ5���O8qy�j��i���t�vI���������Xi_�O�(��:��I$���rPEhXt���@o���|��0n����p�h��bt�`�4f\!!�n�ϯC�\�I�V���=\r3PEb!M�i�4�ƈꃰ1,@m;$�T-�,�xS�ק�.����0>��zZv.O�w��d� A�6,u\��[����P�}d�a�����
�2��s4D�� ���9�>��7  � 
 	   6�  (    P�B�P   ((   � � P 7  wf���R��J�����)RER�f$��UD�m�J�U����T%*�ٴ�@J�	UR��4��P�l=�                                              Q���ALAݚ.g@�W�� :'r�>��� 2 ��o =t&{k�a��M2�Ceh�  ��@7�s`� ��֠\���U�5��ũ�2QJR0 3J�U���hPCT��J�`�T��-J�Ey�H�!`   x         ��B�c�w
P��
�͔*�2P���W��*�Rz� 8�e�w�*�J�a�OYT������J�� 	��2�ܪ�/-Ux4��H�p   8ݼ�Av9:}}� x}��u�#K����Ѷ��(yp ��u��=::�G I*� �K|   x         ��}�}�49�}��t ɢ�` `��;j���0���A�t� ����qf��ΏaF��յ��  =оc�K���i$�f� 9ȩ}���`�;��.Z}�a��j��8 �(f72���S�ܕ咔�r���9�D"�U}�
 U@P       ��eh���o�Rk|��n���
�W3v�]� c��s�=o���v�}��zTU��+��� oi�5��Ź����*%|  A���-�����t�x �L��y����n�������/�U�ͥҶ�{x y�Ur3�TW��MK��y��1�WdzB��UIEo� �B         7_o���6��Kf^lN66ܚ��[siE�x� =�/s;� sh�{���`�֜�(Ty� �
����J�07���(*B[��   ������<](Wy� Ǯ�����n5Oa�p���j�����{m�� �U=�w/p:y<��E<�<N�t����RT� 4��M1IR�  '���T��� '�U(�JJ``j��&U*   i"jz)J���`O�_�����|���UW�W�ۭn��6�X��O��$ I=�9����$܄ ��$ I7��B��`ID@�=��?j���?��z��͵�2V��u����Md7tӏ���[ ��ճ��b��r��O%w�M٫�oh�����	^1��fm���(;P���J��n�:�%���rTRU<����N�]뷠����8ev�<z[�LU���tp:
뻈��Y�(���UzE�_�7�K�«؉��xV:�ua���gr�p$6� Ɂ�¶�Vnm۔J�s��&F�{5��`��ө#^Pʥn���cn�p��Ct���n��:����I�������!�	�agh���>A��Z��9��F�������`d��(�O\�na�P����*Lb�z���m\yE�X��U
�P�n��:�׃*u����Ⱥ,k��p<)ō���`�І�R��̲�\"�B�츻c6٦R�6��Z�ǵ���[_A��:�Z�E�)a����wx���;�k��@��G�>�����x��A\:$��n��VҶj���Kxu%��Ez�s�l�յ��;C��ɇ�5�|�U����2�V��5`Xh�o��Ջt.J5r=��Y�,/t�jZ�r�0v��θ�k��V ��(��ݍ���Πk����PlNH{�}݅w�f�$ 'H�ugp:*����f��6i����Yn�T�&�1%��ԁ�)� �G
:[ݑ��(Wx��Bm�wVEǨĸ�}�%�����(c=���ۆu��n�t!� \m��8z̴�%:�Ki����K�^�H�s���V���)v���K'?�a��0���p��^l�D���ؕ��S��f��FX�Gq��h�o�<��-_�Ė51�cV���-U'����p�7���B[9p���-=�G�S�6>�Z��ݘ�ۼj�A:��l�w�t)��#{����b:�y
DON�`�\:f��{g�;�Gti=6F\�a��e�T\����ʱj<XQ�!�7�}����n��c���J��;&���\S m7�^#`Z��n��h˛�7!�p;����8!���,�I�b��E�I-ڶx���	t:�*έ.�F���rt�6�Ъ�-e1��2���[�˿H�&��l�mP���m�~�ao?ϗ=Z�����61�-�6��AC`��⎬v'�yb�7�t�ܢQ�V�o$�ʴ��WB��>=�^��H�ݻ�f2��æd�Z+�f���93��c�]�;4v�;�&��Y��oi�444#�ۋ����­*�Py���I�d���EY&���ٴ<�?o��ܣ��qQ)�����F�=v�ڂ|U�Y �JBkg�l`�+C�S�5��@qG�f��kٕ,���ޙ���䕤/ef�a
�73@u ��d�[��@'@��sф����j�����PY{��W;1�F�2c΃4�����Bݕ]�u��]ٺ�unU��3j�v=�#:�ئ���C�)�0�.Zv�ʵt|ї�~.�Q�4�7(I�v�nNI���� Ī�x�%0���&��"�r4�b���S��/�l���w]Ĩ���ޮ��&�/�9X;�=�,'H��f]��-��)�{^»ݵ�Q� O��l�ck����LV]�ܴ]�.wW
K.wq�R�K��S��n��+	�z�:k���R���H���� }��D�L�wE�:�Ǳ��J��QL��PXf�������\|�Yqv�_�=ь�yB��!�Eiq�4`|�%/����R���Z��	��ǝ���P�?Fť�8�ff�ņ'��o��㼷�7v����i�;�'˜��b�#c�c	�B4��awf��2$H0�jCzI�)��P/[[�x�N��B1�~�B�t��Z�UƱ��٥	n��ξ�M��F%��Y��[�HH+*ӹ/q�V�]'[F�3���p��ȵ
�tkS{ss��RA���!�9�UYlg.Q˷�ߛ�$''t�i!��|.[UN���x�ۻV��c1�AG8���h�Nw�}��b���1���2�ď뮽��{�ob'��j;�Ս��DnP�z-/{qJ�5�����%C<"�BhY��y	��C뀂0 �`؁v���,��4{���VR���s�+��b�,d6s�M�';7�n��+L#4��ϮZ�� ة�-�z�s�G/y��z�}'M�ٜ���ݭS IwMlܫ��ۜ���s^�àg��`�(4��)N�4X{s�>�/���Ő���B;0����3y.VqX��%�'nHL�s�ݖ�Ûm4+.����L9�U�@��:e-j�����75����R�<�erM�\��]������׹wwD�ʚX]4���v�o��m��B�g$�zΈ�a�?���y�+��-�.Ҟi}��8���Y�-P�;F��rb��KԔT���j���{/w�nͽ�z��o�;��l�!�9� ,��7;R���{�m���z��4��#�T�n��ݺ��7�ó���ZG�c�.��wL7�txr�[��mt�}����Dw,�U+J�)M�%<[qs�N��8K4ܤgl�G[��oQoY�i�N�aC�#m
���s�k��DRn�ӁQ����署8z�c
��6��Ob�b����hM��2l�
�<��/`��75��Z-�ТY�kAE�k�3���7�u{Z�U߬���7f����v��K� �{�1�����{#s9n���L��� �d�Z��7�7(��Y�"�B���#|��&��\�unō�s����tN Qf�tg<� /�!��uޮ�祋����X|pP�[��n�����ܷ7_`�F=#��ŕ��w��� 'o�c��<´S5�*ױ]W-�m�d��%��S���U���W�[���K^W��[���P@g=���q/ˍ7uQ�mY���\�(���2 �C�{���0���9[_<��+�ـ�D�y!�"�̣�l�f>��o@�p�]��g������^��{/w7�8$mʆi.�)ڻmGMn��C��a<Kt����p��"�����8��7N�a{8����i�XKm�C�ش1$�F]��Y��n�%l�]k\r�8,O�݄�ƀ�	 ��k�:�E�8H��Θ��A�(2�0Sza3�dNK�gF�Ci�麷��&�G�O9�h�r�#��0I��g=K;�5���X�C	ug]+0���$i�Wh�]�!"7�#����LC������~�7@z��������p�6�1.�q�Ƹa�Eژ��\�nay#�4,o���Iv�F���3���v2~� �ۅ�(7q�79a]qAj�fL�c8�rӸFlT�s��x�R��Ҝq�{�c٥�x/Ǧ�4맥��owvwE�p�cK�8�9�a'n�� K+3B���8Ñmfn�F^(f�M���O U%[Kma=�C��2��Ա�Ő����/}4Q�������E��8z���T�۲p��s	rA��Z����I ����<�@V�Q!���˛!h,��U` nۼI$ �;I5���V��x�ƍ���=�z��@�]���7�oc1��{rF�gy����'v�_��c���
;S��q3�s�ݚ�Duv�W.��[�S#[wH��y���TRp�!�����_sPC�A�׬j,,�)�C���7p6�`��W�鴞�2X��Λ&[��ɵ��SJG����Rf����=�vB\��"�Fx2z��h;/^��ȫ$��M�͖i|&w7�)o� �2@x��-t��Fn���M�W��W��ò�Z�3�p�c�N/�-�b���!�ӕy9���U�u�[!�����g��7�
������g����˕^���8���d�5�{q�9�s�s���.uI��W��[ɭ��P���o�3Tε)I��`da�8^s;���Uz�z���:kt����[o�b���ͣ8�}���'�p:����=��7�^-�u@��<!�����{���؝�q,u5]��]�K�YⳫ'�\־Ok9��Y� y��9K����5���ǡ�;�� �Z�wJ=���i�rvnvl��>��
W�gnF��.�G�oo8��2.�7󛹨���u^���ַM�qq7�s0pͶ����ٴeOiT�A	RT�`Hpw,��!Q&t�A_�"�,��^�:���s�u9$ܮ-��n�K%�ݗ9�]�G��j����v���L�XHX�o]�Y�8��׃^�ݎF;z����gh��j�6�7T�5�UT���9v���Vj��7���f�ʟL�#��{P��7p�'HF��9�aQ�&B�h�.!��x��c�׼�Ѡ�'4�]ua��M��z��g"2=�;�'H�^\����g-q&?Csc3}zs��Kp��$���=���*�۔('T�r�������;�X��5��y:#�@�eQ��QJ����+R3^�m4l|q�of��"lZ�b�� -��B�*��v�[�.�mF��tm�㽿�K��n��Ԓ ��9q�� e�q�@od3S��J��횻.��h��0���_@W:$�s��+ɵN��$8X���|`ڡ��-4�(���|�[�tn�OI����p2Y� ��&�Ӧ��%��Ū�K�e���Z˺U�{�Z��1����r�����e�n�5����+6���oco)��W6.�I�-��<�sX]{��;�Y�;�ȝ�-�Is��W��ôӦ��ocO�oC���g\a�ݶ7ۗ��L59����W�(D����]��bHT:oP[��A�j�CHss� xܺ�ro*C�)���)l��v���@v��ܺ;:�Y����n<��Jr���r�ɤ���C*�u�KS-�V&'���YyϷ��e�s��p��J{�ݜOt%m��6��p�<��t�.����'=r�A��,ڭ.~1.鳻q7t]{����-j�9��q��mz���3)E�˂�guѳ�A=�|sgu�H��~���#�:���6��'鋬#�`�_	�ܢ[�0��w�q,96I�5c������}w���I�o�ۻ�C+�	b���mʳ����\6��:f�ʾ�)B�Os`��i�rGf����k�zm� ��s�%�HR4Uӥ�ܸ�!4M\��CY:��:c|P�rם��n�(��bg�ho@2��=�\�w���Θ��N��`��� Ÿ�ͥ�m��X�P��ƭ��Y���XX�����{iZ��A�� G����%�w�t�ۃ	W�7K����ql���T����3���5$_��o��U�l���7�%�z }ъ�"����\'U���D��Zj�v�
�X��Zwq�;�Z˖��W��z����jׯV1�]WKa'�rWu�y3��:v�˛��W�F������]׃KM�swc6��_��U:��Wɽ���s��d|��Cū^��ͭ�N�6�{B:�����0�q��N)��rUwUo�n�����nw�j�#un�	7���S�A�y��\k���D�M�v4x#̮@e<z�۶�N����]��75)���l�3�ކ>0�cpf+����OMT`�op!��Kl��F����9�Å[����g �w�O�<8���ׯlł��Z�l%�9�钱��~�&�P��ŶD�,a�����]�*��&Ch�HE0���k��Ot��yL�j����`����Ҏ��(�d���yLz�2�q���� ����!�p��xi�'*M� �c�J�m���oG�S�Wggn6U��d��n���P�&F%�C$F�a\X`��{�M�x�wv����r�b�)���Y�;���j/�v�I��ºë��%��L��1ER��ЁB�t3q�Rf[^��;�����̘uP\�:WKFs#M�y�ƚ�	;�����Y�Z~:����KyL��;��K���l�0�oa1<�?9��f\����c˸ل��/,}�5�4\{uo⺩�n�r>i>�I�8&6�:@9�Zћ8e��\޽�H�X��0���A���������p�Ӥ*���ۡs:��ǐ�:�6���ӧ�:U��SH���chm"��v�Z�~�&�3q�O�q�F>���x���u� �\F✯"�ݘ�O4w��5�43��e����Èˉ<(3�-[�wao�h�,�c��&;�ſ����R@_���7� �p�k�u_��Dh�'r9��;P��n6$�����G���V5N �^��PdkK����6���J��:u��(�է;�OF�Z���j��%l�����W�^fl�C�CtU���\牐��yqX�q��/pӣ��wy��W��Ԃ	�Q�N=s�mh�����;�F7���"H�0��l�ծ�wj�q�Cc΍b��'�u|�c}k��w��1ǣ%���Ͷ()+J�sF�cǼ�]B �3yhO�s�2V�<�*���/s�rK�9C��7,����6ő7V�G���I���.�4�m�����կ@Z:'$]�7�A��4�ob�d͝�H�sXCy�T�ˀ�/Y�U$��:�ӹ��4"ykT�Cy�;Wskp�r`��9aH&���ؚ��WöT��F<vr��	qxѶn(�bbn�����q����d E����I�$���� � B��I$$E�����$P�E�BJ�BV$P� � �d!TXAHUa ,��Y ����"�$ RBAB � T��H� T�RI!	Y$�HI@P(H,�T$
�B,$ � ��"���a	+  ,�@��@ 	+$����!"��
�@$%` �*IY$��P���P�� � , ��XH`H
 H�A@��d YI
��H�` E�%B) *�RR�$ RBEE����! ��� �$�������S���ۙ��;^��Z�R������<k�E��'��#��m#ߡǻg,�NE&"[�������ñ�Tc�7r=���P�g2\�� ���Y�x\�"�_Y���E r����a�fH�>�N�f�[^�\ �bzn�B�qg]�	���f]�IF�2�G�@�� ��
�FM�}���_#I��Ʋ�ڎ��Y2"�\W^=F+�<6~7)�zD�jB�[{�y��*���b@y�֮�Z{+NkƺT�5�+�����Ń_��i��$���ZƂkb�����s!�c��>���.���y�Տa{�*vrp�| t&��y���c���h� ��%&��&,�:�&5�U�gNY��6��4H*P��8iVovQ�xt��U��3BsL�9��V&X�Et��DG���wfPұ+|l��1��e�s�K�=��e�~�yOT�Y��1�]Qw7�r�0���W헶6*�	���l�1�	]��S[�m�\[.��l�w����E+,�qQ�E�EY�G4���]�6�^�*�EH���������.Cd=� �n;4��Iޞ�t���)�{I`�4ެ�R�j�-�������Y���G��<�z�@W�i��g�٬�ov��+��J����e�'������_�����-�����~T��]UN/�.�5��q�.xL:�o�Gqȧ��I��o6{��s~�q����&��-zi�8[�ծYos���0��O;���1`�9K�r��&�*�5�b�q�e�+B��#}+7�����S�����u�IՐU�}�5	��5��g���3��{;{�EK�
�X����YNky%jC���w�Z�-Vef�d�5�y�Ǟ�p�$������p	7vwp�1�������ۋ7J���:y����=���'+{4���:��m�\^��*�5.���4�ܾ��i�����#���`��8 ]�#sF��gB�'�F�-6�sM��b�FF�Yȧ	���8{���8+/w*���w��f�NI��U�`���iV�ںk�gv��F���v�w��R�)��xp��㢸c�	���[I`g�ٲ+��[�>���K�����H-\��-)hwx9�Ʃ
���]#���A���켗�X��ȩH�st�={<�v�p��0�5���Z�ڬ��2��²nT��}+�綶��l�d
#��ի{V��xw	ƀ�_d%��&�_�&�B�qw��Z��ZbL�dm�p�<�e'�ز�yd��0���j���s�w}�����G�͜&�艩6�6+�i��T��5
ʄd}�7���K'c�
p��T� Eg%@,��X7��HQ����r�1TU�Њz���u������u��xsS"/"���\�~|�ueٶ.<�z�4��Y홡I��}�4G�-�wn�r?M37�p�O�Ϣ<?�K�/�\�Q����R�A�G�ci�q��rX�q��_ѹ���N����'�{lB�x���"$}�Lz�Ax��ܛ&��-"�j�%�	2���+�L��u���s�ɱܞ�ݻ�;[�2�y��JҺ��X�r���p����Էv{�x�%��J�22h���wrA&޼9�ǩh�Pi���ު�0;�%��7[1��K������nj���;�y�����n�gf妟`�駱�I����y��Gw��oF�^D���y��w0����炋�`-,���q��7�N���f��{�}�����-tSR��}+I��/�^Se�yN�LY�˫&]�<�{7#R#�En�e��fΗ�����ܯ3��w2�.x��gqT+�2�d�ݣQ��o1�,"x:�m��,9&�1O��7���0g�@ծ$���z�zN;މvز�&x�S��\O4��a�*<z��n3Ol�pX{�4�]$��
\�]��m6�9`���X����|����T>�5����3Ը�R��a
�o�|w��ѣ��~A?U�ɢ9F���q[����� ��,��V�aw��>yEA~�I\M\w\���=���I��n�I/|��ٯ�n1#z�i��v[.����2T��v�k8kٔc��4��t+pa���4RN�oyqУ'��Y��[�݀d;�xRתn0����LXv1[���
=x9�:�9��f���\gf�r�vC�΁5T��nLx�n���0�<J<�8[\�h�a���[�_�̋�ir�g0%S*'�W(��w-�s9F���t��Ηi���q^�~֜b��%䠤n�[���f0�&��1���6u��q�M�y:�o�lULk�alЁ�<��`=���{{
�r�,��R�]΁���BV�>��r	ר�t7��%ͺ��2�S��x���u0�Ҳ�:zr�Wl���a�s�-�G��
,�9�V<i����� ��'�R��|==��Kin�-�pp�
̨Cn�k�P��i��V��
�����f۸z���YŽ3��
�Z�,z�)g�<���7-����r�������gײ�����$<!喂�:�����ּ�y�ɻ��y��W�.�N~��V�\�;��u~@�I~tJX׊���ٷ�	�^��>���+[��sa�g՝��i{�yu��=�t��Z��#7w��Cj�3���
D�H����w���L#0���@��:P+.�ܵ
e9ꏳ�Wz�������(աa�3���$]= i)u���1=��N\��06�r�;�/����)K��*��V�y��Uv�]�.���.����ז��`��}n��t�42)j��
.���^Q�V����Ž�t�r�Xx�Yc<K)j��e�zv���z��6ؔ�*M�����S�^�v�f���3=v���w��i�n ��ܥD�9�=��%��	0��0�8���m���SFB���;yV9��9�G!�e�l��R�On*ˡ.��U�����Ճ;hܑAWVm�f�G�B-���7�/#���{~��gڸv�ly�0�Eϝ��J�+m.Q��-��q�{�{���� �Ή���95P�j�s5-^��������\�:����z=Q�����ڈȖ��c�ݕz(���wS�r�
�2W,��2��ĖUsv������B�{um@&����M8�ѽuk��:p�p������W�^^��)��U�te�H�g�\�J\zl�'6��&Y�I�[�ذ�U(���nؗ?G�kW��z�'�=���\o}$��r������7r2%�Ї��Ʈ���-L�2��#��}���:Z�|�wrI�\��bA��y��l�W�K}ӭH#6��uԂ�ֽ.�ӶZ1��<�>�(�Lu�yy��ˍ��1샫���c'LQeqb��.��&Lw�l�2 �:!����.c�w
��\�
��]]r�	"��f���ՏI�~�U�2k)�r&T����)z�pO�gfc��q�՝�)IV�{}��[ӟ �{�(=}o�]�C�w�e�@�B�)e�;���7���5�*�ĜQiuƀP�{��16�&۰U�V7{U�rgK�eS��T��oHx�����i9����:v�M����Q�yQ�����:a���~��Z'�{Ť��y7=���4Lvw�;�'v*��2�q\2���O��Ԗ({n�ꈑ)Sy����ݗw,8��u݀�o'�xf�E]�ٱT��i\.�P���� 4Q���ӫa�cV�Pu���ꝗ��ֹ��.	VX
��y�Od�m@��@�f-�<�J�us�4ͨ������ �^MjMCyeS'�Go49����������c��V�ޙ0��ny#�X?Y��Lr�	ߖ���y��:��C\�n�I���ŸNO]������,�_uճU�t��
�,�Kve[�WB�F*U���r,��*�7G+���(�Fu��~�Z/;�i�9D�'��3v�J�O��9�<N9���"v>���[*c�cg&��0���:��{O��+b~��uU���|��p�̥ʍ]�/�f�.�����R;��pe�\�������y7Y�R���$�T�5L��DP���4�G�"����^�-L�Jx�\L�oMn"Ax)�;����:`�C70)�jB՜H��θ:�%k|.Ru�"�y�,��W�2�=v c8��9-����d=�{�pP�u}��T��EŐ^�����]T`~	w40lsa
�C�{{���mJ`�����!\�k)]��Fn^T<�C�ķ��L%�<�qd�w?Y�	��{�ٚ���7�~ǝQ9��NL옳Q8��vV��i�4op�i��;p&�j^�,��V���ƍ���G�f֞;�S{u�gELO�w�$;�*�߲�J�mx�bnr{��{:rg2��ô�y�j����q��CÕf���2nN-�$�ަ�8���ɺ9�W�:�p����˵�n��{x��4F�>�m�q���O��Kz(;lo�!�k�vw�Fc��~7 �P�@�ḎH�ҳ&TD
K�9ed.rxt-�'����Lu&L���xV����P��c*:�Ej��}��r�i�|]n>�vLT�:0�ɂ��ڙٺ��jl@�V��PlÉ�8��jf�כ�[���
5����}�dS{��H�^W�wY�vt���z+:��;�����~.>�"�W%]�N��2p<�SpT��l˕F�T��99M�-�������C@��0ŏ�������j��%!�2�kH:�r��zI��o7�L���?v��,�^�'؊�m��u�J���kOn5��m�&�z�(_-~��[#z�$�0��Ƿ@䙎;��\�:�,[��|0YVI�-̗7_�Ŕn��u�������t2��p2�OJ='��ѭ�W
�|x"�G,�b��6�煦��3�m�ݪR�E�8����Omj[lj)�LG=���1�u������µu�̠�m��5Ȫ��9�N�QS�̷V�82��~B����[-��u��f��e�tv<1�}4R�
1���A��}}�4�\����wQ7�;*^tի;���[Lw�����u�Jd��潦-,��Nn%�Oyl�+c�Rޞ�ik�l�����c��H����g����z<�7��Z�#��FPU��f��8V�9�3���w�6=��Tv�2f����c� u��-��i'"�vQ��2t�s���/)�z#�����G��W.͐�����)h��8�廮A�i��y��C*�G��;lǨak.n�J�V��Ml˸�=�c�th�,S���(�|I�Ғ��7��Ϻ�3Kc)|M/�h�=:�{�3��x������˧<��<�3~�D$Tǃ+xP`����vjL	����I�A�'�1�Z8(�B�9C%�{V�`��9�ޔ�.T��[C]Z1B/�-9����Nu�f�k���� �<F���v�2�ӛ)y<��<�:��m����eQ~��7)��ڥ��]4�]�����z���-+�sZ9���f��?\g��jݽ��f<���Ԧ9!WƓ4��;,l��+H��v��y�q�cL�����e�e�:�x+WML���9/=)b��8tUh���!Ͻ���W�]�oI� �/���+�S7����j�h��B�˔$�ǥQ��LsMr���Uu�b~�aM"��D9(�sͫ=x��Sm�:v3Pó x����ٯ���6���wW����j>o&X�>� �_r��}<����+�熥�|��[������j��N�Q"G`�U1��*����+'@���f�u�}�~+�v��v��|�P�R�	�*]�}���Õ��P��t�P�/\�Ǖ�/W�=S���B�+�	v�W��`X�"���o��ߏP���ڻ�֙+�#���/l�L��U�&���z�b\��
�ܕ3�t���-�]W>�����әν��=���V�)�7fy$���s���ig�,�\z�U�m�umL�wφ�eH���9�l�:<�U�&�������oIzGC�իg�_�
�P��kTag��/���Y�]�Y��m�N�
��\v��d��kZ.F#W6��3$D�q
�l���ǣ��I���HĞÕ��p��g�kQ=��^��ֲ����K��E��or^;�=�ç���X���I1�bch<�C�0�
=�,ݛ띧�{݊��MWܚ/jHt�6�5{�+Qۚyv*7��7lѿ��mn�1+�}���@k���sj�UΦ���!�y'��w�%>�$N��<��7�r����-� �O6EJo�S���,��&p�#�} \�6�Շ���|8Ug���F�{�F�a�_=������{0斒�F�������t�h���A�ՃP�e�W����(�����)��9k�o�<2V����*�e��D�@�+Fᩊ�خl����	Vww��Il�����t��]]�]s.����}}����k�v��6e�鬑�I���]�Y0�fA���R	�w�M�{k���zo����4V���G��@"
V\�J�F�v��4.TA���$R���{׳prwvK��#f��Ӂܻ��2�����.����LS��'c��"y��+
q�U��F� �)i���^��}�V���9x�
Ӄ�ϼ�	֔�D�z��D�w��U��_���1���׺�����7
�����(�B�tsɣ��`�Lk�&3t��Mk�]�b�ŝ���jĹ:3!o"}hɆ]��P�l��a��-Ե�0�i�[�!٢�1/���BbR
�
�g�_��	!I�$���z[�C�i�F�(���l[���V9�&����h�x��z�=�,�;
��<F#�67���� &S� ��7)�/3��@��[�ݙq����w��l��8N8�!�\�;]x;��9<۶d׌b�6�^����W���%��v�1�`�m/,r�fn3��q��lm=Fuݹa{=�9s�����r�Jk)כu�n9{s5`G�f�]�H�ۑ^1ϪN�n�8xn��K�Ό�;u�s�y��/�v�d��f��'���u��xN�@���/7=����<#�\v�y�qƞ�V��uj��o>s��dƣ�u�.8oV3�uf�jj^����6:ې^�7+�5ۆԝ!�&��=�#��i��m���[c� z��8Jw��ؘ���S�Y�8l�3��[��N�i�	���7\�O=��z��.��9۫=���<�]��kv�7����qQ��k5�ls�o'Z2����ZwLq��<7Zs�uu��9���kQ���Nܘ�]q�#&�6�J�j�9�I��ۋ�%���2���1�����������㌽�m�oe�퓹�u���n�=���ћ�f���ʛ����[q';<�^ɶ�]J��M���5�u�%m��w]z���gz�9��c��v�j���dn5�X�m<�\nbL��v95˘|k%s�;�}�[���'�4g���v�f[�t��5��C�A�Z{�}��-�tk�n=�L^v��E��z�s��oJax���U�L8nd�n�P�s���S����I3s�[[�U�۝�I4�w�bt����f�{�&;;��c����
^�׋�m�o
w�0w���<�F9	۩�̪q��q7^�܆%��ƃkiD���eG]�1�Cɼv�g.�&盷c��x�kz֤ή���v�n6�Ƈ�E���a��ۓ��������smYD-��狵3�u5�c���nF2�t�ۓV�>�Qv�f��m8狭�����q�N�MoIV=r��(�N��d�;�7I�z��x��o;�����/1m`mgv��ZN���̹�ج��kٺz]�=�8�-�GE���m��3��:�I�x-x:�N��>���;[�q��2�[^�z�u�9�<���r��v-WBij�7a�����ѡ`�������ٞ\�\t��{Z�۵����Z���vܝA���&-���VuF��vu��v��n���<�M�m�j5pI����ف��gk�
]vw�mR>�W�x�61�g�P��ps뮮͵^zW�Փr�������u�:i���q����v�N�sbWvw.�>Ş\�Ŵ�s�{qH���vgnz8zښ��<�kyD4rh����홳�@�L�V�9�4[v����볎���q��Q��fNCn��=���.;g���/����ۆ�^[gc���5�j�GfzƮ�=&��v���nSsƌ�n��-
$������:�Gs�n8�u�kj�Y�m��8Z�J-��u�t�۷hm�9�=p�k����u����ъ�/Okf�����4�����p�oFMp1�˥�8�,#0�2�� �K��u�K�[t�\ڮ:���F��\���M>�C��lk��kj^�#���I�v�=TSvq8�&ݝ��km�d(H�\,eN�]�%�;���]��9(+Wk�mzsm���em�۝�g�^�]�h=�����I�ȓ�e�Gn��ۍ����=��V���`�6�|���5�D9��:#8ޯey8�x�k�kq�}d��O��v
0���X�c�;UӸ8k���t/��0�s�^���ܯ!ݎ�k��{Z���E�#�xm�j���qvtb���Ls��i��{r>�l ����v�vi�F�7�W^ۺ������7[ƀW�5�����F��s�[�';�S���On�6�;�t�`���i���{/PN��k�&����۫���ǜ�v��<��.���Փ����;+��)2�e';��AW9g%\�]����;�5���9�^��9�X$��N9�I�E���[�����Ɍ8�FaR��k�����(k]��=t�r7`g�k�3֍��v�Rl۲<��6���c�X�z�+�	8<���3X2UGK�7���\t�>tv�v'>xŭ��������f���7\V<��]���;�q���`�2�'.�ہ�M:�Ժ��`�׋��^�ծ��j㬺���	F/olv�n��l�i�wkg֠��lF��c�u��x��n�3�=��1�e�=��ۢ:W����n2P8n�eyR���ח�8�z=qŔ.�fMk\�n����O&�+�p�/����6�u��ne,�l�V��5����t�����M�JL�ψ��	U<5�ۮ��!�[�qQ�\v���f������u��vb���N�ܽ�ٝҞ��4;��m�ۇ�͓���:ۍp��Y�qgWc�5k�7*u;eh@�<`�,�2�������������r���ۮ%�%�@�f�=�k^��۷`K۫zM�áՃ���c��Cu�/k9��S` ��Ak��]�v��r`z
��Ӎ�kb����i�*4��k�F㭚!{v� �wf�q�*u�[�u#X�^]pF�u�����ׇov.�d�^]c�-��vݯ$�=�ܤ;���c%Acof��v�a�:���-/��X�D2]�mͶ���Cb���C���+����+��`���j�k�i�wgHvg�g���<Q�n�m�/i��)ɹ�^�O%��[����Ʉ��0�ٺ�:���pJp��ۡ����z��S��l�/ݫ�n6�\��`��9�������r�]N������[��v�=ԝSN���Zg�������#�v5r�9S��ݱ;=�ݽ�j�s��b:zcrh���ۗ�n��Fw�=��l�:����b׎��n�7R�Vͅ�cۮ�Mٶiin�f�.��#v�xwd��&�¦�뇦��VB�zr�^�s���nܴ���=�<��g����۸�[�qj�����VӹɁ��j�����vl�c���Ok*�6(��m�|4RG,5����8�Hd2����FQ.z�O:�v����l�H��1qt��Y{q�v���i�.���;�>^��ݴ�>yT�^����;D��ۘ��s�t�6�q�=���j�8ގ9�R��m�۸1�.=��롐&�� T�>۫�f���lu�mN���fgY������&wf��Ơx���ڤݎ�2�Y��t���	�m��7�x��y��|�;8�C���N�Nɸ��ٸ�n��s������<'WS��v�N�D�̫Ӹ����i�q�}���=�����n*ޤq�-�i�;%�m뷱��bN;hN��=��v���b�c] �v�i^ۛ�M^Cf��$���^�nv�sm�"[t@�7'XfJK��#n������`�c��뛔g�i��>�����iH;m��q��i��g;�m')3�m��7lnW�����;c/G6Y�ϻq�v��.d��y=i�k��ds1���m��KY9����Hs��v�\���l���v��i�q\,�gttl���6ծ�y��p�S�\�:�ʕ�Мu=���v�oo:;�s�����kns�s�On��e��q�}�=�:�ֲ��buٵí��=[�8��ٸ�մ\���q\#Žw��c�c�<��]���V�n=^�����l��Y+hr�\V��klX���{'[$����8�g�4s����X,f7r��Ө�sc7>ۧ����@���mj�Aa��m㱧84q�\.���kGs`���۶-n[��ݫ��;u��l�#;RK˶��J���j:���Վ�ӕl���ݸڳ��]Pݷqs�Įv���\���:z����/h6��#�N!�I�fw*L^�C��(�N����h�ؗ���+����>ɁW�v6`ӭ�ko'7]�(��[�C�zո#�m\:�]�n�f�ݞ�8�N�Y��ց�9��wl��4O���f-�;.:��ro6����Խ�r��wH��[��d�p�����q���FL�h�i��{O�p3V�=��gCks�3Ɏr��8�M�67�Hs���={m�Gh ގۍ6�*���3,�<�s^۷m�L\�k:���n��]�e���0g�hUM�|���{���q<��kb�5Ǹ�v���{c�Q�P���v�Na3���s����չ4;Fq�\���h�ri�V�����C6�Q��5[����N��wu!봞�{$�{&��Aڶd+rE/���b9�;�	�KUn �g��zx9�d�������vϝ���-�ٸ�]��ݒܔ.�潱�h4��1P\��,15p(pD0{\�rG1���&9-FL��񵧶��t�Gm��x�n�w@�Wc㇄붬;\,�̓��s>�]1]Vn�\�βқ>W�[v�k����מ���k�b}ƺ��ӗ��)���e���q������d��6�w�3ϋv��l���-۹�7n�TZ�cv2���x�\8;X8v�]�8����lWag��+ӝˊ�޲<��&��sl�<kS��P]7�mӖy�]�ZM<�c1�z����ƭ���O&�V�V. Nzb�;[���v���\���nw'��h�+Ͳ▭�j����崪ꇗpAw;�ZⱸJ�t\n�m��؏v)�񭷮�e�h֠5�����Y��k�m�OZ�n��ێ�ך�qBD*9ˇ��:�y붫=�p98����ƺͷU�V�Tڀ7[��U�+�kΎ��n�g���{]W5�j��u��tK��y��Wq����Ű��mE�z�㜐�۔�C�n7Pm�6�[�n�����l���%��]�a� �m�ٺ�V�t !u����3�����x��:� g�i��M5�c%ֵV�i�Кѭ9ɋ��U�h�!h�iF"-[[F҈�X�QQmVʬj[T���+eDm�G�jG#V-���9D��V�Z�\¢�� �Kj�Ee�ZKh�Z5�V��\���mb�ҫDV�"U)e�����V�Q�-EQ�J�-+E*9j*eKKK�DEZ��0���[l�Z�T+ƉB��+B�b�J6,kV�JZ�[j%m��k)e�R���QR�JU*5h���s-jY[P����jZV�-U�k�-k(��h�5�YFԵ��F�KVX�5�\�`1��f*����ڶ��,���[R��cZ��V�KKhĶ���m)E`-KR��R�ƕƬ��mkB�6�D[J-�,���4m����V��m��m�օ�R��mZl��ֵ��J���T��ڈ�T,J�bUq�2Թ�-YV�[ZR�Fֱ(�5KJ�KD�q���-��m�[�-��Ԣ)J�eD��jږ�����2���$�����i��KuC].��g��4�Ù�84�i��T��2#L�p�4-0�
��:!D�s���o��y��w�/k�#��>�Ľu�^�v�V�ݡ�&��{W[���C�.C��\ZF��c�^݌�A��������r�4ćk�p��Ƈ�v]�n�Ƚ�'m��'�ݶ@��j#���S��#�Q�!	�r�q��95��mw\��"sv��/N�����9=��|R&������ZcU*�,
�d���y���q+�؏m<%���|��l|ۨsn���/Z�v��ũy��a��E����V٭���n��݆�{��]A�mý[���lݻ3���1��k�2]s'��)r������{3
��vϏY�6��nk������2��yv�ř��Y戝�{<Vظݹ�k{n.�.��Ŏ]eⶔ=�t�ݗ)�Og��<�W:O<�u��j�D�kl$Ǘt۞.wC���;K�f���귤��4�7F��{Kz�46��q��[��Nm�	<��3��W]f������{K�:�^�E���&;o�Hk��u��[�)tq'b��,�V'�j�в�v��q��`�ۋ�x^���Q���%yt��<�9z#�|G=a7��7��ܽ<�Ay���h�糠��W7B�۶ݷF�&v�˻h����x�h�n�qvA^���eM+ɣrV99d=��4u�O�"���/+��fm�`y�Ht�o9�;�	�c\C���l�mu^��z��Ş��<�f�ˈc�z�������J{uM��0`tv;q������`k���.ůI �B�p�Ŝ7+��E�][ni:�I�L7����%(���Glv��]ݢ �n�xj��������;�6�m/]f���F6ѱ�����oGb:l�� ���u"+��o-�I���6�)km�9���]�/<�p��FLubEx5 z���3�IZۈm١}���/���<p�<s˽�;eGvx���@l�{m�;/�q��r�� (�N�3��N�{!�v�d]���'.��v��s��L��vW��q�'8��1�����֕[j\r�3+��E+�'eP�p��۷�9�q���-��L����K�mr����J���l!�3����Îw<�����ۗ/a�xp��ɲ�M�o<�����5�=�	����5� P���B��Ɂ,8�ܚ�Gu[�m�O^wPf�	rRQ�&�d��O�,���o/�X ���l�|p�ezA3�.6��aC���S���;=L�"I�1[Q�m����$�e�2���*��I/;���Iõ�$����
DH!A2$P;�wv��	����t���	���"�$��|�������l��ݦ��Q�&!)�T�<r�� ����!��$U	��o7�|H:gr� ��ھoǰ��fns��ф���:<Z�d�{�QZ�W��j4h �����<�C��D)$G;���|p�ey �t����81S����	���=�$��IS�aHoź�~b���c+�S��6&
���O�-�bs��K_��&OImSf ��JcE,}�.4qo�w)��S��z�����a�z��ł�g�iK�`�B��n��~$��j���s�@7ZK�Q�Q��׍ݡ$��l��Ƅ�s�QL�Qљw`�A�9�>#����>��;L�"I�1Y]λ(ҧTnQ���A6k�zO� ��l@'׷����5��n (U�`���wX�H�$H�ݷm�F��S&�6�T
5d�*� W�����$_^�~h�mY: $7g�o���.�8��P�uۮ�1�z�n�1s<ܵ�pVv�������Ij�}��ݗ�� �� �H�������r��uV�z���:���6t�$A*eH��|�>$���<r�$�!�^6A���� ��P���<ji�>غIR`LaHbjs�ξ�`�Em�1�o뤭\g�[i̹�7�Mb�����z��w[[�LoQ�^�Ӵ�flN+��b67�!�����F����dn85�#�I;uz� ���lm�HF蔕�!l0���h���gK��fۙXH���d��3�������FL�S�;�L�"I�1[[=m�A �ʝ���qY����l����w��?��%x���M�Y3�	>��8|iR��c��ۛ`qj9ՠ�� �]�O/]��5ҷm������IPL��dB2$q�ۺd����� �F)܊��d��獓�כ��7
8j�(j)S����~W����P׽�`�F^w6I'�T�Cs�=Q;&{]E�"�%I��=��?0ܯIj҂�ۙs���	'o7���p��	 8�IB`J�-�u>sN�=ٕ�,[��~$�3��	ͫ簎U�y���sm6r�E�I\�v�ֳ�\��bZ�ĥ���F��vI���*�[Vq��}}�u�[�1�c�أWU8�Vލ�ޝ�m��01!���~) O��UgmI&��V�ü�d���w*A'6�����DZ���2v߮��ԃ�r�qZ�ݸ\����95����x	j���c^y�b��~~��'Psmiz�cm�|t�e	$��W͂93W�OJo��|O���5n8(&`�2!(��m�k}�I��Q��~ ��{"� f��dI/o{NC3s��k�:��F�����K[^�0oO� `��_ �5��9�� ��s�����:b	D&B��o���Kk$A��t$�Ğ����{��ݼ�`�8sn��.9��IR`LaHb�s�a���fͮ������w_��r(�w]�`�H����K:\�,�����Ѯ�f�:e
YY�}��Ǝ�Vڽ��[��-�}���k����9�ز���3䑃b��,�Y���I��ul}�,^���V:w��ڨx�K�o7m��,���۟g��7;�t��T�7g�8�)��)�[��99��<Gk��q��mۮݠ9╥�v��Q�r�:�WkL��Վ��=��D��攋<=���t=8s���Eoa�غ�J��L�tv�{{��f�k�]�c�8q:펍���ҍ�kc��L)vh�l;���l�ԋ��o+�#��xx��V+����յO�9�Ǧ��ߟϽ���H��_����jH$��$�ަ�;*y��e�9��O���~۾�Rd�L��MGu��I��V�e�Vv��F�	d�{����
]x�X�[@2v!��y LD#"E��l2H;{�LA%ި���Nga��{OĒ.�y�O��*��eDCg��d󌢭7n
s���H����$aיʈ�����CA8��~$@�V�(��H@����|H��ȹ�Q\���l�}��͒Iï*MtE׺`]�: (&����M�����Njj7]ۃ�s^�{����;�v}�i��	%L�����[��`�����ב^oT�k�
筲A>�����ۮ������!l1.*�~
�xDY��Trk长�E{%f�U��3= � #<�k�ۏ4���+�=I~'�۬���ۤ�ǖ����EΩR�nM�wƉ왦���y�� �p�ʐA��*{b�옺�o�"$�J$�&���l�|x��2r�݌sS�&�Y�\I9y�߁�ב@��hB��T��H���qs|'(�v]U
&[�H$�rא(��\����w�H&&v�c��(�DJ�3���E3�wK仹qA�H
���A>8u�O��wͨ��M��&J/颕�������P�Tj�}�m��z5l$�:fJ�c��[��]�����?]�Q!8=��0Iï"�$�;��-B�5$:[u|�$�l���Z$�0�
2)��9���z�`��w�;k�p���既I���s#D��������aMG�hI�]x�� �tH��x7��>$g2 [�=�i��eZ�=�c����;ӷX�)�de��Z񚇧	�un�g�[���U̶T�[Ob�_La��w�A �א(쮾l�]=Ȉ�d��(LD���۠�1D�xĺ�;]z�$���2/O���^�	&�c���
AR
�"���m�6�z�n��m�x$B�آ|NW^7����ɌD:�Qƕl4V��,}(A�~D��ݔR[]�4�nSKok]�o]����~�߳B�GF��w�����/Y�0 �ose���Ր5�R��w���6F�#) f$"El���5��r�Н�&�� �@����A��o0�kk����jH��	%L&FC`/:�$��u2I5Gu�d�ʮ<�8�]e�`�H��� ��ѐ�%2`�Nԝ*�&n� Ի��$�f�?<H8z�������F-Hɘ!���I���{gF����ڛb$\XÚ�0	��ꑛ�����<��^-�Mc�*��%'ٙC2�5�,��C�
뵿�t�""A��L�1[�t��I><r�ܩ��4,�Tj6��$���͟a�ʝ��MS�-���.QQA�cX�p�]r ���b���@ŵ�:��[������t2!H*AR$w��v��ަ$���"�5�g3�AjKv�$���a��7
8D����*�[y$��5q0�t�O�/t2	�gsd�A�ו� �Pw�os̚S��FOw����P �HD�:��I�÷�$�NM�31�Jr������2|p��I9��I����D�l�:��;t�og#&ω/��?G��#^E A�w�N7Z#4���Sn�����,T�����3W[�w��5Y
���[�t df�Aӷ�+Č�|��Q��R�R�v�/�N���M.\����O2�f:J�tT؞'��)���'��x�.��=�8R���F8�r���n�������O���7����[m�[�c�|�m��cv˖h�$�Lm��/i��G[}L�Y����ǖ���D���!ۇ�5�ڵ����[ ����2��|u��Q��R�xy�����Jܾ����mXB�ˣ:�v)��wI�n��b۲�sv�OGl��z|cs�l���8�i�����sF1�9��=����65]1��j�1�N��N�v٫��f��#��=rq��RG=>��[xv��Dܓ�^�q������n�a	�������Aӗ�$�	�w͞������D{!նI =yBH57�U)) �J�ok�p��Ȭ�k�6u��Nw�o���Ȣ�w͒i^j[�?�NSN����t�:������sd�P��q����6'3	$���H�w͓:t�@�3�"�ξov�*�ʉ'	]פ�N�	&�7�/v�ԕ9�ޗ��-����	&T$��0u������r�<ǘN�y�A"��6H&�k.�6gL�Yo:͓qه�gG�g��l�q�4��ڈ��87�w&N6n�������4i����$N�l��{���=O]�3��U �r��`1��
A��L�12�O��W����y���<l}��l�f�ı��W;G	�x	�����}�wT���_@7����AV�>m���)}�ݚhfŪP����O�����$��l�v�N<�e���IU�p�""BR�vm<� ��ަ	'Ʋ��C��r����$����>$��l��Q�$�GAI��uN���{��g9#`���� ����i��zd�zr����Y VE
�s���z��W	+��	�c�U�kd������N˩����߾_�p�Ӯ�i�j|�ړ��
m�V���=�Mb�\4�h��s��Er�4��._s� ��������ՑEF�S1���&�T��wX�$���lբ�1!JdL�Q4��$�׽Š^��[V������$��� P!7z;,s��V�����������|/^C ��;���>�ޗZ�Xx��{��}m}b�wf{�.�������=jÚ͉-l�W6��
gz�i�zR���˧��H�:�y�'��_7b]ӇN��S`:fEi궂{�R��]�����Vɗ��ɹ̝���1�K�k�衩�o{e�
K�:�k�}�sj�x���tt�:�ba"A��v_ozVy
�=�C�_�չ�Ɵ�=׋姞�T'`�	��2A��Ѻ7"wSw{<H�͏���3���g�>���w�����v^���Vz|������Ƈ�������}<���HN,5F���5�.FrPǊ��t�|E�S��={1�2�Rp�'MLӄͶ�j�Fe:�F���[�P�o�d��p�3As��a�X���Y��g������6K�y���!tQ�M�Ǫ&mY#㶻���������鷊\�\W��u�<��/Mí���NV1�K�MbM���m�������0�y_v>�xQob�Տu�\�ǾWU����8e�K��/����}!�0ɿAfz~��L�U����B��/��0����P<�;6��������&�ʟu�m��΍��Ysq��ѓ%���	�*�p;d8�K��]×��x�g3�%*���LX2�Q�X��	IC�OeKt�N��`5���y�V������k<�����������Tyw(|�,�y�N����h�K.ܬP�n�ӏ�Y��ܕ4B(�-�J|k���.�!{*�%��r�	r�����۝9v젔��W2��ZXQj�X�-kP���LZ��Kke�h�enZ9if\��ĕV�����0�"
���ѩmZ6�K��ԵJZ�JQm*֣�Ģ�(�[\�m¶�*Z6�rՈԹ�V�ZVYR��Զ��b�Db+KQjZ�1��U�e�0��R�mX�s3
VƵ��KZ�iQ��jUT���m�6��J�mDF�Z�J�R�J[D�DJ��%Tbm[V6���m-+m�-�eX��W2�J���A�"�T���Q������-h���1h�B�R�KjV�TR�+E�kKe�-�kh�KkA�aR��V��-�#l
������-�6�Ҍ[-m)V�(�Q��V(Um����6X��UV��JV�cim�m�)JҔ�j�ԥ)m�V�"[EF�J*�TQihж��եm����J�Z5�Zح��j����U�R��VҬZ4�Z(�DKV�ƶ��|I9���$�p�dP1Y&f!D�S"B���2�����]��l���>$}�k"����U�ݪ��Q�@�����v�5n��6>�C^���Fb�s��#�n� �=Y���������:fJ�ɢ��)A T�<(�a���z�-6S��Zv�q�����rx�?�����*��S�9�z�'�a���H'�]|�.�:��=�T��J��{ѹ\O�8r�):�$ϒ2P���Y�,s�x6T��UH'ֺ�=Y[��#����Z�w�l�lF�P���D��
$I��|F�f?2Df��7�(��1۳\A6q�H$���l����0TH2�fCu�����d��<���E�nS$w�̅�����_\v>���{���������e�2ʼm�@���<[6M�8�p��rA+��v.�ޥg��;�����fbջ��´��~���|��SFC�Z<Ƅ��(	����ǉ&�6���"2bD������Cqͱ�؎�pNȷ<�a�ױ�W\�vv�9ꮮ��h;����Kt�٨�[�$�^�����A���� ���lBٍ��=H{�|l��	�f�2}�2g��0�O��7i�d�R{I.R�we�Ԓ@'κ�	y��$�^roe��r��VW�2HHD�BBo���a�r�����Q��)B���A7]|߈���
�X(HF%D�RN h��8��P�?r��I>������������[UUd�x�D�1
`Toc��D����xy��˦I>����>$<�^�r�9%(�2�8���^���5���P��"�<]���Vq��#��]�* }���%���>b&����H:E�x�B�*`�`J$>A��<;*�V��˪ۑ�LX�lv�]v�1�oY����n�OGtg����Lt�v.}�7B�f�"�s���s̸q�T�z�uR5��G<�l�WWn�n�:�y-���q�x6��s˻P1���jKTW"��	x'�ݼP=�Ìr�gp\�ӻcn4�c�Cu�����[#I=m�����K�溓�{gɃ�L�9��c���ټ�wI����:��,���%���F��5��߿��I�0�IQH��;��	����`� b�Egq����#�6b�t��d�E�w0�9�Q�%J��"T�x��	 �4��;wʵ���2H$]��g�y�/ݦ���o�/�}���T��#����O��㇞T�fʻ�6�n�o\�ea$��w�����W�:�2�	�(HT�.2�c��L���!���L�N.y�H9Oz�@�*kW��_��o� Q+*�eX
�t�X}���ȇ�X&��7�H� W�#)�6����֭[ �6�>��AD{r�vz�v�]���C�d%�:���1ή������Ș*%*T�/��	N<�>#)�Sz+V�������d�<�
�p�aH��
�4�v0�6����:��!�:ݝT���Wt��rx�IV W��T���▯Rs�Xk���h"��e�F�i3_8+��G����ؿ*���_xI<��P�H�|߉�� ��(Ǚ�t�^����6��b��P��(I ���d�Dr�}]y9��y}��Oy�[|��0��Q"Q��D�n��֮2l��HOfԟA!�^7�Iy��=u��X胴If3jH]\vf`������p���\��=�0U�Ȗ��Q$��^6O��oP�"Lӕ����/�]O�H����v��Ȫ7U���7����뙌[�8�<�mv�Ӄs����}��א� V�	���J�� _|؂LuD�:2��SYa���2���n�f�
$*(�"�m��?��]geM.vE��I�$���l�n�z��7ؠ�v�{4�4�KV�CwIX��μgă���� 䩋���]��r.(��<�ӗ�q��(*����{䢴L��;��	#��(7uDƊ�v�{o�����Np�}���,���sj�|�W%Yx.G���p>'�/Xf����#\�(�QGw7���K^Ͼ}�>���Ay��$A�ՙW�2�1wA*��£���(�B�W���|p�e	鶮���9W�w*��|z�$����W�5	��%ZXh�"�.Т��n��v�d��j��݀����wU���rr��������fBR2P���s��#/{��I b�ȣ�磏2�(���7դ��͂D��P�!j�7@۠��R���|g�N�m^�� �M�o0�	8gr��{`������濗��bT�%B!iow[d�̡$O���Z����d���u?	8gr*U��D�J�%D%"���������t��})���G�"
;��l� �+c������x! G�~y�x3�Z!���#�:V�oN.��QҺ�q>�}��Jި*޽�g6mo+�M�����Ҍ���e��'4�d��E7A�r�Õ�`޿�{�}�y����_]f\��]]\�c�!Ă�^��a�I@���|7_�g�}﾿��뼼�H(�w�}��"V��]����t��Xw�>�����WΝ����_�����{��A�3iݙ)�몬N�m�=���֦��=]�/:�������}�q9����S����l�p@���Rۿ{��M�RT��ϻ�8�X}����y����I�w�y��������߽ܞ%��]10�(��FBb��'�����6|�Dx}\j��PG�G˖> n�m$JB�0+Osw�O�@��w�>���pd�k^�^���>�>ȾU���#��!]'��3�32J��!�����?6��T�
�߼�vr3���Ĩ��y��G�ߺ˟o��D�
��~�������A��k��>1�ΙAAR�J*b��g�sg���}}t}��{�:�ђ��W��l�i
���߽���^>�"3;��dz^i��X(��E�?2yR��;�<����_ؚ�ӗM̷G��<�=������F�$ �����!��8���=����V����@�x(�YS����g*A@��}�g�p�+}��;�����S����e������X{�Aú����q�Ii��5���ȉ�z�TMSU�ef�w�r�Ȧ��,���=�d�:�X6��ڵ�����6k<��x�p�n��ôa��(��ͻ-e=b�^ݝ��i���0ö���U�9e��g�}�����'j��z��nQ5Gk�[��y8�5��)��¼�����Ȱ��x�h�l7��
݊1ǖl���w��N����ǟ<1�xN�ͱ�'�h�;���$&?���������*ty�xM�r�n��8�|����(2N�k����k�V�=]\�<޶2�u��~˟����a�u�C��
����x0�J�H,;��ݜq��� �o|ő�O�\�]�����]y��y�AH4,?o��p��nu��nj�U�k/��$�~��g�� }�}�C�����
��{��=B���%Bĕ����wq�H),����Iȅd�+'�{���}��;4�w߷'��
f�v���Uk���/�8��5�}�<`pjB�~��l�!iOG�-�s7�<z,8��~�E� D"eO����8�Y��P��w߶qD���gN�p��Y���6�����@E�`�l���T��H�>�{��8�YP,J�w����%`V�(������_����7L>|)
��>�̯6��b��(̒�#�N$����'+(�R��{��ޢwʆ^|eG��s��@�<��ge׃a�°�
����߶q'+%O����_mx	 wG��dE�+}�W�:�<���{</Fקr8��DD\'��뫨\�f�9�B�7�v������ݷ�;��n0>����{��<�-)
G�+���$0@���tZ����~��~�<gFJ�2T*�߾��8��β�bT�(B���g���G����QDG�|����0��b�s�:��2�0��L�z\�1Ӛ�ݼֹ�.m����;6��4�Э�����vf���ih��Y���%���r���@?�L;���x��*A@���l��X�
������)����b�f��0�²����`�Ti��q�]�a���$�~��g��� ����<6�T,IX_�>���Ƽ��?C�?
��%��l�ND+%Y++����Oh5ϯu�a �(�)� !����䮪7Z�XHR�=��{��R��h��?f��4�R���ۇ��Oe��y������<g�����8�V�?�ᩎ�Ct7�m���|��݇�6��T�������8ɭ;���k�����*=߿}��%`XԂ���$)K����x
��~��~�}�����o�a�7+�6t1�pf�ƚr�t]�]�sם(�-k<ף����￟�p�N�j��8�$����$��FJ�w���hQ%H,)�~��!�aXo�w�ٝ�>�=@�u���'P��� �]��������:��s-ѳhD�=�ە�π����r�����z� +��
B�`W����'�*eO���^}`�ȏ@�����־�����V�y�3�8�Z�)��א�0�׼���IP�,B����vpg� D}��܆�{=R&�乙�2>)e���I��6�̭��I���"#<�����.�^U[�1�(�T��Gӗ���y���s�����J��H/n���y�A�������Ï��w�2�10 '�	�ϨY�}_��5����@�Ag+���l�2m
$�T�����wq�aF���팏^e�NV���Y��|���׼�E'��&fIDD̢�G�>u���H[@���g��m�����mgVW+��"�F}��I D�������r2T��C���g���ޛ���M�H�L�2��&T������ЃE�u���D�{$�yK���L��ݯ���}w}�ˬ���a�a_.����IP�(�a���vq�d�*J�O߽�� q+z�<��=��$Wz�p=� �HZo���8�`V����u���X�.y�Ĝ��~��� VVJ͟�Y��2I�{.ۡgޢ#ȏ|V}�C� ����{��8�Y82�o��k{���گ����H�I��T%��6��%a�~���AHR�=��~���x"<	@�w`�=�Wՙ�GeG�xH)�@��>߾�p�8�YA����w�,�`�#�o">
fR� L~|,�#�oh
��C~t*7|�%�?y�?l�g
J�N��߼8��%H,
5�w�w�4��~����ؽ��3�����n\npԿ]гu����ή�~oHv�Fsw��ɹ�`a0�7�x�Wf��6���Ŝ�70��x =��<�K����8�^f>��ZtWF�Xa|��}������ VX�YA�������6}��ww�:��V�;�C�9VaRT��}�gr!Y(2���ݯy�� S�\�c>=����!2��F�Z��Ti��Q�-nU���l��ӣع�/[s���w�lL��
&e$�@x�|�}@Y��!e�~���l�!m!Rf���$�s~�rz�i�J�hO���}�Ì�%e�����g�������N��47C|������~|(�"#�}���?tD%�3@��9�:�JʁD�}��~���+X�G�k�?Ry?c9���<#��p��_f�y���\MfWE˞@�q'5�߶q8�YY++%}��<6�IR^{�w�s^����8��¤���{��$N��~���5�폑%L��(��1D �G÷>�e���s3�
C�@�~�͞r���+X�����ȁR(��߻�q������k}ߗ4~���%B�}����!�%|:o">
fTD@3&k���Oʻ(���AID+������d��.w�~��P)������
5�F���wI�B�����8�T�����ߺϝ��хo{S7Fw{
�7_��[>�T��g�'��ԹSe�L�o�S���.	�}�<�؛�u��%���4%�R���=�ޜ�/�=|��[O �bM ��F�̫��X]I큜�h���1� ���3C�o�J7c�ؐrɏ|������\�7R����H��� vr�������mM5�uޅu�C8���t��>�q�$[�� ��v��Q��/,��jd��|���0���_̱9J���32�6A/.=�]���l�{:��j>�%v���[�'�ŜeY�#�6k���/O�Xd����t��M
��[�2��fL��a��9�Xy^�Oj��	��}zG������:�e��2]b�ݤ8Ӌ��2�������&���}]��j��&� ��~�'/��k�LwPW�Ug��Z7ק�w�z�Ib.qz��6��\�y�e׼ހ��.��]n�d��;��[xz[�ݙ����v���n���n(Ũ������(����g;���Ǯ�fTt�9o���V+�X�ޚ�o:/eB��3Q�w.-g���N�^������VA���7 t�}�K�� "�w�ݔ�}�w���%8n�����t�=m�j�qʜ�`�Ը�clKb�������
���օ�:��D�����	`��q�5׺��(k��Lt�������|�ẁx�tk���跳}�Ǻ������L����ZUm�
QDFԵ��5l����ؔJ#b
����Pm�V�UFڌ[c(��YkTb��Z2����E�PF���U-�Z�T*�m�h1E�kTh�YDDYcX���imv�TjV+l�cj��V��m*5�kmR�b
"U-A�J�R��\r��Ջ[)VT��Ѷ*�-Q�*����m"�+iQdU�J�D�km�h��эhX�R�m���
��eʲ4m�A-[+mP��"�
�V��A�5�⢔U�kE��Z�(�R��-ZQ�9��2,�֩iQUR�Z*�V֋
�UDAjF�U1����Т*�X,(�kE*6�Dm�j�h�F�*�Z���APm��b��QX�[V�m�V�ղ�Y��ѭVҶZ[V�P�ƭ���B��eZ-�P��F�T++Uerـ�ԭZ"�m���Z�+k`�2���������eZZ�Zղ��b��V�R�j�l��+Q���
���Em*�m���FѶ(�8۶��v%/W<�\�B�Y��t�lnm�c\��:{������mɲ��ە�s�\�l���pw��G���=��ۖ;��q`x��m�<�7&��wŝ�zw��(s�a�N�]�^��͙�8%^��9�9q-��`�1�=�����"Vg�ͼ��p�(���,bq����٫���n�G��{r�ݬ\�n(c�����X<mM�Y;m^�ѻ	�p]��T��q�'�Hvmr�ݕ;t:Ξ��9�rv��v��Ԙϥ����Ʉ���B�5vm�Y�c�L[�ӝO[���@�[�쬢�����MZ�,��Ǟ_�lma�"���^�ŮV2T�v��;;���j^u3onn���s�9A�s���0v�^{>ݣ3�����]m�\n�vQ���6���8�u풢��5�7nx�a���_eƔۚ�eVQ���z�t#���w�N��ݭ��oՇk�>nS����也k��h�c��yy�����"\����m��u�ˎ��Tx�A�۰*�����f��ѪL��l�t8^,��{'gm�:�@p<�z�\+e��1�˧���\W��N�&�AL�܆:P޼�YLΑ�M��%��f'��4�.+�9U�lٻ��a�:6�6q�kNn��n���Y��v�>��b���m�B��l+^.��}n���9s��i�un]u�B�)����7.�Ր5�k��j�.��:^<�<�b7V��6����o,lק�n^�#��Ej�s��%t��rl+����]G5�7��u���z�����ڮɲ��l���^��ؠ���v�e.��y��9���{m�r��� ���C��]�Ze9�kvz1n����{KGGl�k���¸؁h$�ཹ��N�v���x��u��A�ګ=���z(�Iѻm���/\t�<zwf�u��vz�(�0]��y���R>�.�u#�\ezÞZ�Z�����b�����j�:j��GM.��g-� ��>�U���w���{��f��`']��6�V@v�,lj��f��� �� 5�Δ�ܰ�>�]�P%^�k�{r:�l�ކ+v�4�7X8�Z:�b8�<�$([�Y�8<��n�3m�d��[	�ݻ/�uVi�],ź�{>�d�n�oS<#�Z��-�۸[�y0��4�6�9�s��y����y�^9��6��Ú��.G���/��&M2��nKq�˥Èv�2۱�ۍ��Ӂ�A���	=��t�4S���?߽���k�t�/�@��<O� VR2T������
Aa�������+�y�5_>u�异�I�~��gr!R%e}�s���3|﹭a��nkN���Aa�����g�/G�E��_P���ns��)
�[��;��I<@��wϾ��Ă��g�{���˾珽���|��8�Xzk:}��A����Cl<W����$�
��X{�ﻸx���@�@/�����-����b�u?�:��Z��_y���n�iHZXwϾ��ǌ
�G�~�2���7E˞@�q'5�߶q=��^w�_�u����2W����M�A%B�J���}�|�>�G����,�nG/���N�hɶT��|����o�v��ї-̷Fͤ����{$�@������<�Zg�����|<8��"�3�~'�@�P+����3�%e��x37�Y��>��\�ս���O��t]��� ����=g�v0��\N�&��i�ٶ�%����_�Y��9�~��w���|����
K�;���gq�����߾���7�y�0�������7���������8�>�k�3))&b`@O�#��P���2Va�9��g�sF��y�K�i����2�'���Ð{;(�6�W��ٹ�0]�3�	�@�Ykm�wz�#F���ٙ��F��ƛ�ЭS5u�#n&��!!$���{�v�B�*%a�����0�0�+
������gpB�Q��>���ӝ��;:���r~M�]o����5��iվ@�Vk���$xZ@�����IQ�����>~g?@�t@�P+*{���p�9+(2T(�{�~��8���קJ�4��T��|k~tp޲6�����H)>B������H(J�O{�~��"V�`V��ﻸ~�;��?o;�����R�wϾ��q������ٔ��.�.n�}�����H���围��D����s�a�V��}��q�V*J���l�Ad�+%e_�wrx�@љ��Ͼ�s~�?��;�$�q׬<=��E�m9�v:�N�N%�=r]΀@̑> �̎�ϒH̉P�BR>@Vw���px��R�=�����B��)
�i�?}� i ���o�߻���^��a���w
AC�w���H,=��3�NkZ5���5�x�_m��8
#Ȁ��㯾�#k.s8O�s�}���2VT
%@���� r%O|(�϶���@!��[��mT�F�xL:���<	Рeq��T�10 _ )�}�y��$q�������vxɴ,IP�+^���~�=���wZ��j˷��9��r������9��)$�V_eq���7���V��M{��X�ź�t\á�.q��H�� 	�׿C��°�*J���l�NT��FW�ﻩ<O,�����a��2��LY X!7�P��k��lJ�˝���ԅ�s�}��)i
�hw���� T��'w���8������n��Hpd~�9�rx�3��.\�vCq&�wz�lH,��߶x$>St~������@�@�,�|��{���) ��ﻸq� ��ԫ��?X�a�zfPPe��u��l n�/"���C�%�:�u��Wk��~�}S��Y�C�>��9�y��� T��+���P6��J�V����0�
�9�|�}����8�bg��8��
�O���;���2 (s�RFdLB1Hb��'ó��A�<	C�Z=�0u����JB�B��_�w�����+(���wp�8�YA���K�Ż�����y>��$�ę�""D�0�a_s����*%+�wg#8�YP,J����oZ�����}kӨJ��`V�~����yH)��w���8�^\5�۬�n�\�ž@P�#�}�P��qϔ>g���#�"<矹��O
IX^���Aa�@������ꯍ,��Q�5T�U$�
{�7��P���J�}�����,�A�\��7k�g%W���%��N4-�38n'욼'R73���� �2z��c+˿��<h��������kWV�q ��y��ǉ �~�}A��j{��Nm��<��i�׀���@�=�~���82VVJ�n�}B��<��E���P>��P�0"=+��3�+#K�]�1��YƭN��q�q\=�M�A��`��ǥzh5����a�¾_��a��i%�V߽���'T
D �w�b��'�}��w�|$f��
~����i �H[a����8�]���s)���.�.n��I�~���$pd���u|���s������g̛H(T������$T��l�'����ӗ���W���_z˧k���Q /C���3(�!� B>gn��(5!e�{�}�g�)
�Z0+���RT���/��I@�� G�Ow���8�����D;�����q">t�D|$SDD�~G�<���@һo�5�� "<��yBϬ�R
��� pJ��Xk���+�eÇ{6<	׃�~��g�"�K�sY��.�Y�|��{�=�g����GVvPgޢ�����l�]��G�����~��0�(¤�}�}�gr!Y++%_��=� eѶ�����.j`��)P��\93YW$��cS�o�՜p��ӎ&�F��+f*�o�*1���B�CYoRo�f�g���v;K��o ����7t�L��ݕR37�� ?���~���ؠ���C^�N��n�ȶ|F�n�s�iѽ��v��
��H��iK;�m]D��\O�N��wO[�:��M�;�κ��;�.��d��.P��]V��G���>+�wn{I�l���HGF��ll�Nn�ݦ�.���q%�M��۳PI
pn`lݵq�n헵�)`��<lٻ�vV�u^�nI�-n<��.��e��A;o�x�;�-V`�bJ�s���zȐ��+~����e�q��C�w�����Xy���a���H(��߶y�B�B��[�?s� i �s����k���Y��nH,�%@��}�g�q%aK�N���k3Cqo��W����H)-��;u�����~��YĂ�bT��{��8%`V�(����wɺA�����_����[�ۇ�#��>�FA"b�
��,��P�,�R
A}��ݞ2m
$�T������y��O�s���=V0�*}�����8!Y(2�VW���w'�m�s�R�&e(��1D �Gþ���W}�G�An��-��(��+�Pv��i
����?s�@�AO+('�k�>���"��;�A���;��pIXY�o�gƜ�ֳ1.hא�0���l<m%B���{����8�����_�����D��ﹳ�%`V�(����������W�^o��#��E���z���A�	z5��3ٰ�ֹ��DA��j�^���c-��{]dv274�%H�2J��>������`�YY+,d�o�{��d�IP�y3��_����Gú'�̓�k,�x�'�g��sgr!R
A~����i �s>��Q�fbb��G��}��g� 
#���6Fs䈏��b�f�U)����������n��ҧ�v��j�@�s��ff%T@r�DwS�ʓx�)Gcfwn:�|�Y��0ć���x{���;�����␩�
�_��p4� T��?o�������T<��s�Z�ZYT�f�6��G�> ����	b$��Cl<a_/w�����T*Aa���г�>�>D �B ����ҫL����:%`V�+^����y�A���xgW�^G�6{���R(~Ȳ=|��`���ӊU� >>�}�eJ�w϶x2m
��D��}߽~G�#�����G��>��$�8d�ʐ\�w����@��׿7Xf�kV�7G�������`Q����������������#���@�AO������Ì�%edD��P��<����wt�S۹χc���n�nN�������-���ٺwl;���7\�u�	�i�~��_޶j�p����0�o{�a���T�!Xw���8�2Q��@������%`}���>��.}�h�~`z�/<��i �HV����x�W4������in�)�N��Y }�|�g0��:�z��B��T����~��q� ��~��~�Ĝ�T���y�g�k��֗�=�*����(����1 �"L�B,����݇0(ԅ��}��<���AP>��g85�ӍO�}f�M�I�nצ�:�ɍ:���qZ�ə�=qh��ism!��*ǅՈ꺨���R�3�P��{��G׿����R�
ʟ����g*AB�?{���!Ȓ�{ǥk4e���g��Z���j���h���=$G�B�������8�P(���߶x�O��|O:��wfQv�xZX~����8�[<<��ێb�X�s3�N$��s��'++%ed�����gޢWS�̊�>���=�y�ꇉ�T�=�����8�d����8�ux	 :��}�����Te%��q�rv-q�Nr=r��uK[�%v6��y(��;R�}�TęS2�R>G�>���5!m����<�R��k��y��<�����9�3�3���>�Du�T8�2VVJ��w�~�ĂÆ}��|iu�kY�sF��pa_o{�a������U���_t���$�ov�>�� 2�T��~�� q+Ƥ������A��;���w�r��}�~z0+K�w.��F�kZ[�<}�{��'
��YFJ������AH,<���?{����q��°�*J���߶q �q�������w'��@�Z��Z��HQ31�d`�|��@O��oW|��[����jB�����<�HZ�H-�<���4� T�ʟ����8ˮ�dW���X��X
�D� a���)r����Yٞ]l��q�qj�e����"=Cx�sn���Uf�2Xwcw9�4����@�'�2T(��߿l��+
�?��]��fao����l<a��B������vpg>��.�& j%@��}�|8�X�^�?wp<7H6R�����8�W���~��~|��ҫ*���[�0����c��)s����:Q�zy�k��߿�AD�N�+�������l�>+,d�������<d�%B��)����!Ă��������<>�=�IS����8��VJ2�VW��k�`� Nw�d���B���O�}���g�"��ۜ�(� ��Pv�[HV�
��<���4� T�e�����Ì�%ed�o'��|��x��g�:���>��=4��kZ1��^C�8¾����i'�B��
��w�vpg(ʐPg/m����~������+��F�����xn�l�-����q �a߲�Ktj浥���bOw��l�w����=���S�ϼ��|gY++%~�����<IP�+���<a�����gg}B���h���~��4/�d�VJ2����p4��߾�kW)sY�������9�}�q��!B��>���!�Į��]�bL�hww�wI<+(�����q ��}�@�w���>0������8��ҷ7�YW_�3�2��4����oi�jl�Ω������e	\�=qtܳ@4�r�rۮ�W`�k�9�ww?@��j?���Z�l�)�;W��%���۾c�n.q���m��:ֶȩ�Y^#ZR[U�vvz�D]vXú����uΛW�����K��.]۸Ab콻q��n�I�Ӹ�<��C�0<�<�ln�3�f��9� �W=m�0vkv��iW6�k<vs7/��s��ҝ"��lnG���sQ9Ӹ�]�:
���E���ے�덆ts��]�����0����v��݆vk��:D�!q�qu>�x۳v�����[��֌�-����
�u�퇃��T�B���w82�T����1dd#�8v�O�?W����>�O���&���w����ǌ
��ϻ��f5��C��@�pI����N VVJ�s;�zw|�Y�����}��M�D�
�������0�¤�O��߶q'"��VG�w��]}�og_�����M�Y�5�m�h��Ӭr����J�߻��H[@����r���@�rm��_f��ջ��c~Q��'���H,9�����r2T���~����q%a�q��\ֵ��ѭ����[�@+��~^D�_}��@Dy!Xk�}��Fq���%@�����	X5�F���{����=���̭󼾾�zR�}����H/%��.��F�5�-��	=��g�e+(2U��{��O���ϻO����IX_���y0�¤�=����8�H,�e^����/��s��o����(��曨�񮬅�5Ιo*�-!�۷<��;�
iM.�h���Z��2�k5�_��%a�o�
A@��}�ϊB�B�`V���� m �n��������Y��{�y�q�d���
!�>��H,��	H�B�?
>��s�^�� "=׃m:Ks�2�%����l8U�e�F��ɶ���9᭛G^�8�`�����p!����&�fi�-yzq�-˚'h����������,�o�}͟��%T
��s��� pJ��X��=��y� �B�7}��{��[���s����F��Ң"JV��3p<N$����8�++%eDO�v�DG�������b+�a]s�:�хaXT{�߶x����������^�!��ns���& ��O��ve ��"����#����@���ݞr���*Ai~�����@������3��s=Wrx�P臻����Aam�|is5�h�sF�u�_��v0�%B�������g9��ٻ¾J�Ĩ�����9�+Xj�ϻ�yH4�-���3��g�#�}QѵX�%�
���J嶅�:�v[�m	��*b�8��s��r�j#vܚ�����HR&"bA]�	=o/hYe++%^����d�T(���y���`�#�;�9�'![��{�<��y��9�������=�������3"b"S@B>o~�p0+Y����Mߵ9�3�<�X/� ��� >ڿ�~;y�з]�k�'d�J@�T@*}+v��W������Z�f(�Y��*�''j�왛��6z�4���Dx�Gn$r[��H�� ;��S=�ݞ��LW�n�+q�����:�ɸ��>]�%k8���tv�l�(�	/�c��m�F.Et��t�ul�����Y=�]�Y5	�T���쥔�jvp‴�-�(�/2��.�DU���—��
&AYV;��Z42��H%�\�yc��];�u�ݶ���G)�Q`�4-��foW�X�m�Br�"5n��N�R�:p{+2�:�$%�}�hf�t��ܲ�����]�z�q/Ғ��ǀ�-�72v�11H����=���S�Gj7PS�C��]�@�s�s���4-\8ˮrŶ��b3����7��+�j �s
��U���<n&qЕ�l��.t�\ْ����HM%�gvk6�x(M��fF�3�ս���5<y�i\�A-���Vq�'a|��,�{��	��5kPU�˫��������dmH�r�������M�-M�48m^���h���|�=[2�"��N������[�]u�{�p���Y(N4��;�V`�v�k�샸
]YS���}�*L�G��P�+���3y|�`/�="Mg�bt�g���~�����'�B��&η'�*��/;]��#�
����o�4���ѝ=�֮�4$�&2�k"�2xfJ�]�]��{���ʙ���{��J�"�E��`���՘;8M��M���gMH�m ;�UՃ6���P���.Twr����b���w��|�ՠeKVҪ~�ee�,�D�X�Km�kj[��kD�KZ�%e[J�aim��b5!KjFVնҶ�Z�R��YR��Q�e�ZZ,R��UJ��V
��)Z�Um�4�b���V��m��(�Q�+m[\���2��H��D��iH�U@R���X�6��j-�,���j�э��RT�V[Kj���b�+R��V�-��-�m(���R��(�E��,�Y-Z%�l�%����mZ�$������*�jF�,��b��U�4-��`Ċ�*T*�����-��im��[X[c*��" �j��B���������-�JPmQ����EF0[h�UiV�)X�T�j�+V�Ke�Ҩ���FҪ�+V!P�,�jTb�ƴF"
��bҭ�"�(�%J��KC��QXbV,�,-�؉Z�V �dX�J�Im�D�**�q1`ʊ*�ۍ�fZ(T����F�UET�11E��-�E�Ym��2�O� Ṯ��I �e
Gm_���[�TDz�(����w!^co�ҹ�@�n�@�yW��>$^_s�G�7Z�5� ����w��ú�Z4�\/޷�¤���fCB�bV5�G�o�xʽl���<bN@�W2aI��P�GNϯ\����M��Mٹ�#K�ۇFm���--oj�
o��p�
fbD'x�ד��}�d	�������Fv�q�A����B�'��e@ͅ"B�1
3�XO�y�sf-W�u͂3j��$���l*��M���]k�I�i��-��Y���I���d�|v�5�<�Z]S��w����v����p��*� ��Tf�0�0&\t��I������l��w�n[7�B��K�T��
��,n��{�όu���MEp�;�]YG�9��+�$�Y�2����Z��ͧ�4Ⱥ�W���;vÉ��� 
�®�[�>Vv�L�0���m�	#��gw�>�h��x� �okp�mI�S�mF{���
R���rt��F��}v���nd`7[f�u�rG^�)�z��ĉ
`��"xݹ��;��LA��[������o�v�kOI��Ғ՚��>�ō\��}��M�+n��o����$7[R	k�n��O�r��ͰH16�
D�LH(WO=l@8n����StwzE��)�� ���l�I�u�&o�L�^B�Doź��/_oOE4��ăѵ�� �آI۞�.�E����p�]6�&���)��d�Jh�����A���%{b���:��'�7���I�u�>���h�c��>�u�7�6N��NS��n����fI�^1ʗ	�����ݹ��C�כ��3�;��U��1�wk���\�ɱ����$ K�G~�e�ĺ�T�9��r�l�x1��A�v�r�0<�{t�bؽ]�sayӶ���e�,k���ϝٴm���id�g�p�w[v^N9�]������5�ت���n8��q��yr�b݀@��6K�ۚ6 �P���\�t�㎭���(`4t�J=�^���.�l�����e6�ӽ�^P:�n�Z�m��s�ы'E<H����7]�NL��Ftݕ�r9�ݸ+�q����~w����*�$B�y��I>#n�h�H۞�UE���\�]�`�>ڲI�u�DԬ鈑"`�
`Ț=�x�$T�w�[���W�A��l�;s�L��|m�����UU}cR�V���]��S{_��$�{�\�e�R�ts���~ �����A>s��$��R$)&D![����D��*�\r���6f�Q�>9ӹL�ov���f^�B���2�LVU��13)yI�)@��u��$�wm0d�r����k6pOt�S'���kx+q��9w"��ȴ��74�+p��Q+=f�z-<�2�u�q����L������o����ߪS�*ɂ��"�v�@;���';�hv��sd-�>��@���s��¢#Љ�"E?7�l0s���bn�J�*��쬥��g���y#��}֩�ӎjR������4�8o��o�
��H�qCn�	�`�GIá�ݓ�q~+���F�oޣ�>��)�N}�m2M��3�Qw�g7��߻9H�+
µ��\��A���~$�Yr2��۴呂'Ļ���$�Π�z�w�bdȂ�d�{o�9�o��p���Io3h0H"��վ�U�2f�1���u�����
D�"`�Ȅ+���A>e���}�	w����Ι �Φ$]���+�����-���~�������m���KL�v�!I�g�:�6�8��_���߹��D�!ź�a�H7۝A�M��׍\`�$�{tC*�귭��Nu�6 ��	L�D	a�+'f�PS�o8VU�tof0 �|��$�g`��Wm�;nlv�waQ�D̓
!�>���'�����:t���}�a:�5k;�O>�2�:���
#F>m��;��G�ٲ��Rݡ��-�p�9\%檸��eY&���X����xggv��m��0A��hQ5N6&&%J&B��f�v^r��ɞ�&��$���`�	�׉� v�c� ւy�c`��0��j:�aR�Y����y����v�1�O����H��P$��l�V�Ψ�:1
HVl
�H��R�خg�s�;q�����[t԰����M�����R닧4�B�5��A��hI'���c
�c�ү�w=2s�?�0P��"�g���B*D6[��ω��iN�e\�N�(wg��"4�T�����X9��7c�UՄE��B}}� m���;ƥ�z���$�.�x��=�0(Wf �
d�Q���XJ�$�ɪ�	'6{�y�����%ВY�&����qn{�R�M�p�=�g{�D�l�˯]�I|0�}?�)S�B�Lkz�2nԉ�b ��1c^�A�)�t��Cϓ���z]��5�ZuWF�4f�?}���#s>�g;��]«�L�M���I{;�� y�͜USS0+&�A~)�w��ӎ�G�)rw/�׭�`l�uw.�\j��`�肥�_�W�DJ�Q2k�8�$���l�H���6�yѕ�td㪐@9��O�D�2&���P�޶� �����'�Gd�ef6A��߉���Vt�i�|��|�z�|땓ufe�dCSہ�H7��L�
����V�$�̦>'י��'#�M��Uuao��'ev�>�2tǜ�����$�F�o6	�/rs܅_^�Fe<l�݅D@&�&C`>��� �y�<b�/jg��2fw6O������K�[�-F�M������L���⤚d"�^����=�h�󽽏a���_�(���l���xX�� '��dL�Ԝ�MDV����_~��=��JG��6��[�I���F��[�Kv�X����q\{�;9�L�	��|����ϓ��vӤ�ՄM�f��NM���D[��v6�;�;q�����G�y���$��g=�i��;X*¡�}��t��e�I�ρ�Û����]�V�,v��Q�>LWL�T�C��G��v�۸��Ny^6�#���m��lkW�n�+ٸq�aܗiyRq���=qq�����sUucg1l������^ԅ�?�����*]5��wo�u���w3�� �}ko"�3��o��.v��N�w0�K��(D��%���(I&�_O
9]�*����0I�fo6>6v�p�v����p�޸�o��;�(ȑL�B����$y	 �g!eL���sF��H�����ï*H�ĥ2Dʔ H��:�5�f��A���`	$jǑD���8�B�[;�(��|���P���@�"�'cnH'�z�* f]H�}D��A�yR	���qK��W!��ozTf)%J�&f�&GB��u��z64�M`@�B���(�U=<���q�����)*���)g�Y}�0 ����6�;s�;�`���q�A �ו$�9�&�)MUL��{�i��l�r	����p���N��
�#*���U��1{���}�vK�Fh߅7�єHso�Ogs��fo`)�bï��O���:Ţ\����x
�-�ē�F.y	�>�63��jUU	�t���T��3%D�D(�-�5�^�e��`�`�;H����	��*A���~$�ؐ�HJB��n��!�U�����+rA"�$A!��l@$]�s����%�)'R����Гq\v%)�&T�D6k-�? 7{�Lq0�2�ǷcI�wz�$w�͕�gRk&�B%�����q��n���u��.��<�9��9�ݔI�os�(S�"}�E�P�F��l�w���.1IOP�(��	�]�PbF�a�(Ɉm��?]�i>9}6Nc�$�c��&�;��9̾]Ip�\7�e|�ZI]*7Jեu�]p���d�n�*�F�������0��f���ð�ev�٬��GROg ��e�CX�;�����5�{���2D*�wX+� =�x]�l|��0M�w͒*^h��bBD(�,q����ynEP3�H=�� �ۛ̀A�:v�Dv���i8+�����	HS"��u��H8v�#E�d�J�9=ף�v�6$��s`�4��"�����ߗ��hΙ��f�� �'N:����w`��/V�eݺ��Ew=m�n������bu�ND���>l�o�z� ��Or(��Q�X	{7��A��q*bg�'Ќ�4cv���21�1W��I���`	:^�	��2[N�dWn�C�p	@�2d�l>�� �y�$����[��;��kc���� ���E�D�4�ZV��g.��ʃ��6-�(�c�A$�}�D�gso�>7O��5�$���>��i�m͚i��yp|?T�y8"�*r��#7�\��B��-u���k7<uA2f�\� Գ�6��}��< C�ٟs
+�1蘐�
fM�U�O�]_��>��,�>+�v�� ��	��_6{�"�f�j�9�c����z�����y��]atr����Oݸk���s�$D�Q���dHJB��<ym�����~٫:F��gP��m�	8k���O�SeD� H���N�������ϺF��̭�ƻ"�'��o��%�s���vʈ�2�}0"}H������a�L���<��gs�V�G I�=�'�9��̍y�� �&R�a����*�⾮��*H$���0H$_ws�m)騉��IF&�I�ظ��$@3"T�M�ُ�w{���R��9�Ö�Ex�v���'׽�٠Ga�t���hO��n^]Էw
T��d��47��IӸ�ǹ��wO0l�p���`�(%N�^���m�ه=�/C��p��k��u>�3SH��$F�^�8G_mĪL���sb�D/4�~)�ڎB}��OZ�0q����!]xs�`��׍7B{Ni���E�ԋ_J�]a�j�"�2��J�ܻ�9ע�tit=5�@]wrw��{:	��l*-=|Ĕ�A�S��{u;ן���dE�!ܙd�}�f��/������J���,轷�&wc�/�q�f���ڼ�Y�ס��ɻ����Z�8�Jou�å-{������r�-˻�ռC��slQ����9�!Xf��=�R�Z�1��t�5X{m҆�ŕ�=|�/�zǚ�+JOu!{9�c��ӎ�_�%�������۰�P�SC>�Do9�0��GMd8�;&��I���rrؽ��^ؙ{��� !�[��t�;�x,&���Te�qȐj�t�e�v��1*�Ȯ�L	/��;�LJ�2�_3D�\���B%t�$��5�V��ݺSQy��8B����W�����U aW,C7</R�h����Ύo����慸..|�w��?g�+��Ҩ���	�& � 7N���3�#F��xGZ�dč�ln�㌍Ŧ�Y���іQ��a� L�ځ��t����w(�x��Xչ#�4+��osȍ�t+	���(�5�]e��b�cض��H���L���ݧ��)8��xF=_i� a��=����c���=Ssc�v*Tm�	�#
�R��Uv� ��Y�QQYU[l�U-�K*[bZ�cYUm����1Kem�F�C1�YiT[lF�DTbƠҖ��\B��e�lY���Z�V�U
�Z��Ke����Ң�R��(1��JYKm�+++-(�V��Z�J�UE��Ԣ��8�(""��h�H���L�Ŗ�R�l�B�h�YZ#2ڰ�,�R�mT[j�ʩE����Z�),�`�Yj2�-,�E�R��F�[-mP�*­P�+Q�AjUl�R���h"ܸ1ƈ��J!Ym-e�ڢ*�P�Q���G-��*�Ցdh�Җ��U-�-khʕ��V�s)�k[Z��U�iQ�1���Q� ��ZE�
��P�eE#���4J�+KKKUl�0��cT�B�*Q�"VV�ڂʔKU�)E����յb�ѕmj��2�QH9Ic��ZƖ�=�}��t���TK<=]�=8:�S�aS��ݬ5�aQ�n�a��j�GJ�;��7l#��nx7R����n�۪_�1ά���;[��Z��)����u��ڻwl�1�8-�{��Q�n����!���ŵ��#m��+��֗.[k��LsmK�4�P���i�v�;�pK۷��u�U�v��C&Y���]Z�m�M��Y�U,�[m�T���g�v;c��.�۪��z:���\�Cǹ��=����������}u.��J''K��qv������tu�K����jx��dә5��H���G v���Ƿ�@Q�Om�!ϋvy�:�Z݂2X�ݽ��yV��#��w7OH���r�o��S��
H�5it������N����6��3`F�n����t7�:��l��>=G�:�펜k��\�|����l�<�Yɱ�W�����@��o
P�mݜ{1zݺʝp�Gb��;<y��+���u�8f�<��	ګa��'��cr�T��)���ϵ�����v��;�r\�ڱ�|�o��`�[����{]�����s��+�B�����[n��uƜ瞌)Y���6�]�"]�75���S�8��X�k����m�Ä��q�4�1�vȐ��q�����m��۶6z�k%���re��·K��/]�����6�Nq�m��J��筘�q������h���k6��{9��F:�:e����n@�;F��z��s���Z��n�T�t�NԄ1��tr&�y:���qn̕�$V�'gr��=�M� 6�vu�z�kq�rv�6�;vc���zE�')`���r�zpF6H�g�mv
�b{v��92@[��j/XnX�)Y�w-s�k�X��z�׮����]�ٮ}���]H�ŷ��x��y�}z|V�\]n�퐹��1��ݶ�|��q�.��z�8�-�����]ۆe�K�q�����nD���:6y��2��/���=sx֛R-љ`Liš0CiqZ����{�����|���J�g�S.�V����bn��fn�[���>�tt��7Y\�V�q�{[s�n���E�2wͶ����`֌۳b��]����m�;t^9����V���w�n��� �v�������]�;lq�nl��1��yt��=l۳%���0Hۭ4�"�6b9Ƃv���)��Wn�܂�9�<�`v�lz�qtA��p�[a�<�s`�׮ND�FA]�7=�Ng��nf#���K������c�3%"̝�l��	>$�]��}}�͜+"%x���U ��]u������D![���|z�h����b����l�M�w6	vd�D
U�Z�+�D���B2$M?��L���d��`������>u���}���Ĳ��߭!~T��8�d]d� /{-�H���`�A���tD�F]f6H��r�R�e)m��l�|G^9�g�����d���l�Ggw0�$e�sͰ��iv�EJ&h�%B�'��t�jx��v[�Š�S�tm�F�θ��l�d�}�����(�I����޼l���� �H9}s^;SL�!��k��� ���l5�eyL�H�)�:��	���%f�U��}���ү�7�B���cgMhuu��[*���U$�V�.�	P�2��Y��y����؅�{����oo�������.��P �=�b��Q.���(IwI� �2!
��`�e�РNP�G�"a]Yd����lI{;���]KI�J�,M���_@��u��V(ܾ��H$���H����q�/��w���-��&Lϔ��"h��u� �s�1�f��U۝�W ���$�.�������0��ʅҴ��=�y�'cU� �!ۍqv(��#v�Re�l��P��QV���	A���IO�y�� �F��I�>{=���l�[|+�?D�k`�o�P��鐢$@0&eLM��l��xfnl��1]y�+j�Iw�^'ć��!l���P&�����-X�>S2R!D�l���	Ⱦ� �r4`ܨ��v��*
�(�`�u���Fn�	{;��$m���^uɧof�X�:���uֽ�S�����"��#	>������Q?s��6/��߷�-[�d@3̈B��Ϛ����F���$����H'��~'3��,��1!�Ag��T標2�TAFD�lԽ����D�jA)0�Κ$�23��s;y�lL^��ɷ�F�DD�#&D��*��9���1�E������Qa��չ�v������2��0LO][B��;��g���fv�`�-����EG]
q���D�{����31��|�&�O�@7C��$�FGf6O�3��`�76�2.�a]�,'Vn�"�\�[�g����IqWR��
��rz:l�C��l���͓֎��3)$�L��tx�v����vn���c����l�I}��M���p�;���2���a���0�ν�,^q�¾4�3��J�MOi�s<�Lgj�VGd@����Fj�)��d!G:�D���A�	| � /l7�� �EwI� �2!
_u�I ��ʥ�S����f�D�*��A��� �E�e
<����dcI��QJ!`��vw�lw�X3sV�a�B�|�v�;��������ꈑ*�2$Np�޿2	7۽L�H$��M١7p#hP}ς�l�H����)�$R	`+V�.��~}��_��jD�*��]�������+��M_;��G;�*F ș��u��� H#�2�1��J���z��9���̳�݇��P'W�ÉiZ��J�&�K�b)7d����H$�ۙ"�]|�!q�Kn`�	r�7�}Ո�ɔR12�mm�r�����&���d��_6	$���7=}L��q���*b���2wʜ���
��h�r�ἆO�i>w�̣&�LL�^��+�r�m���mB$U#�3�������Ё���c�k�
n�{"/\n����Iֱ����!�c^���wE��4Ar�֍�;n.\��ca�m�fx��l��p`��v:�5{`C���'�y:X4]�t;����n��ٗ�A�qZ^�/k=p�s��^���u6��;��.J�]N$���xޞ֞G�Gn\[��y�WW-�9�nx㎸�Miy�l�#Ίm�z8��Gngr�)�O&�+��<��ֵ˘۞��Ml�]9�5+�dI(�R/q�&"�!����$����	����6y]WSt,�6�*�D���2��A�"D�j^s���5�Q�����|>'��d����~'��p�:�9M�4�9��S ��������ds����n�&r��O;6� �E������`�$k��J
�S-���hJ[����d�s$�[7B��ް�M��>�Ǐ���`��}TA��Ȕ�%	L� �m���w;z���b�Q�ѡ �k��zn��$�v�0QjhA{t�b�(�EF���~D���]$�`�x{F�ls����w)��6�6�e�'�O�������2d$aL�|���|ɻ���o�Z�ڃ���r3č��a��F�^�"�![]��$f6�����]e�.yg�nMߦ�z��b
�:��/[z˓o���l�{��
�.�fn�a��j�Y���Dւ��q<g�m��п <<۪��$�ӗ�d��߫���z�0/�w�Ju ��V�Z烓�`2	7��L�FuR����\N�E�����}��2�Ԗ�Ҵi34EOm�b�h�NO[~d#7���$��}��Qw�2;7�o���[L"���PP$J���+m�`�I�+ԧ�i��6���h�ݦ�'����d}�H@�������$��4D�
 �B���7��콯5ZsΓ�j�r�Wg�{RϿ߯���E	�S��x�$�v�	�#d�4+��g��[l����1%�D�)B��o�v��(�#���Z��au���� �Gn�6A��+�9�Z�Scl�^|�h$G.�|��U�F�}W�\�V�ū�"��W�.}�*^w�Z�%�����L�pn�&I��:���g&��,v�8o>�/�7�ur۹.�N��CL�.b������{�ߛ�1�W��Ol��J�T�3�f�����|�8}�#3wi�H$�ܑ^$\�ck�5pð]h�Js�߉�mjKV,:�N���yd}k���y���n�I�cd/���O�{�����~�_�m�J�$��h�AH+��%:�=�qy;a�f�M�󊗧��m������������ެ����'K̯I�@����h�8��.�w���$�e�W��4�a�PXqQ\-�׏���S��Hut4�e�E7;��#E�ë�"��5�߳���:�o���ro��	Q��Q΄E]���w�$E���O�w��J�v6J�	&!Ck��p���3~`� (���'�=��$^v���,���A�bĝS&]�QZ
��qw\����-��F�)�7�Φ��)�( ��uy�m�o���� FN�Nj�S��*���ผ�|<=�?��i��9�1*S�i�R�����S���UF�9@j�&��=���7��هYScGtRhOm�R�!z�Ѯx8��hv�ڽ������u�ރ���8�rm�k����ffdHQ1
��ES�F��?3�A>����&C��}��s<G;��x����w�B�Q�"R����c~�����plF@k�d[� ��ܦ	��{�$�9�Wȋ�bS嚾٩n�KA�RҾ�_��>'�w{��I����Οtn]$_os`�� ę)B��o�n;�s��GV5�K|��|H$^�s`�u�Ud�T��b�#u�a��#��H�`B�]���HevU�B�˝����m�	'���$��R$�Q�K�6TUc�sBbQ�f���{�aص�=va�`�-$�������WN�Q��P`�Sn���wԯ!2p��Hp�m�����G�33?.�����HsC*P��v����v���$f|�r��O��Xb1�l���;N��uӑ�����{��:.=Q�u��!8z����gO���⑺���/ls�PaG�������!�2]]�j�m. ��yR�u��M#���C��/u�Xٷ���Cnw�;c4����d�gz��c\u�"�������e�6�:a�:�KQ˂(z�c����\\�,[ٛ�μ����F�*ޙ �$����fbT��Rؘ���2���`���d�1��9M�=�����oĀs.�L�Ȑ�b3�ٰA��O�Եj�f_V�	'�3��� ��ܪ�O�X����$P�!%)�lN�7᳗��$T�b�n�b's��I���d�A[�8�N��Դ��ZW`�OE��w�ɪ��P$X���A�ܚ���,���ŷ��	���l�� �2TB��l��t(r����y-�N.���l����	��f�n1S�1u�k���w�z����K�51j�L��n�jy��n�]�5�)�s �~����zy;�r�H z�`�{��d<�T�wB��C��dC@!z�a]�Z�V�+z�OI�>��]��w��7��f�&z�]��xh3��=�@�;����=F^�Dv9�4��u& �o�m��{�%W�h�	$�=WΚD�/�{vM�&��	��TP����_2s�Hu$�,:�w@]�g_�̀��x�>9Orwc�v��f>m� ���f$S{��"D�30��T�t�m��ήɉ�&�ݴؐ�����7���z��7^�V����{9��|Wd�%L�Q!R����r�Z^Iy.��H�e��j�r��v�@n�����ަë}�������v���I��rq��� ��i��˧"�gT/Nn[t���_>���}�ź^��@��4� {���� ��h7ïO�T�X��d o��f�:gh!P�`B����崉3�WWe)�Snj����d��39�݄�IyooK$�$kcw&w�g�]�3�OjիQ�J��MW=yi �9��L�H��٩��6IV�0�f��b�M����2(w,�or���v%�.�Z�u��͸EŲ��G�P��wvbw�@w�N�S
^��-h1�e>���V�����"�L}Ûn�U���
O����M�x934~sv���y�!mx��g�y��;��ϰ�5��T�XZ%\����Eht���t�P���
�i�n�Hծ�����eB:2�V3eS�%��ɩwJ뽧�	l-Jx�Ϝ2��s��A���|�՚m3}�R�<��˼��yu��U�]�	y��3n*�R�u��gJ{Ҡ3q�y]�_�G�^x�v��j˥�=WǬB�V"��/�.��t��@]�����e�ӫ�շ���W�J��Ξ7����F$YG�8:���²%2-�����8x#�ĜP�-C�Ƴ89X�z ���P�} �WwY���vP���Zإ�v�c�e#[=9o�!J�a��]AMNO�0+X��Z�˹�T�ԯl�E����ȊS��UÃw�ى�
�z���b��i�KL�C��C�:������3Q��o�����u#NU]�=,��ҫF��-�����Iq;�3��@�����BQ�J�l��dd��Ѩ.�I�0��ﳞ�Feܛ)�A���ʑniVu�]�Jg]�k���s�s9F^é����U�I�R�rY*��K���"P��b'39@ع��:�T����;�y�Z;�M�����;D�bk��cN��V0΄��5�H�o��f+�Ǜ�����^X��I�d�>�]���G#!@5r$�)�+���:�jTF�i[j
�E�(��X�q2Ҩ�T
5Dmk[k-�UZ�Yh
�e��DQQETPAdQ�QJ����ڒ�A�m��e�J(�m��[aR�kAbԨ��j�k��Z����e���P��b0�cV�Ң�,m�� �D�[J�2�*�R�5��-mH�EQR+h�T�(,�**9�������r�LJ
�Uh*6�PX�B�����e��lDc+DTj��ij�KD�-�QTV����(ֈ�J���R��-A��T�J�Rت��ۙY��X(�R�VD`��E-�-V"�mR�Z��m���E�UR���h�JZ�+F-f$�QL��2���j��V�`����j�%VX�r�E\����TU��hQ+2�j̠
�/��������73 #7��`z�����&�8�����9�5fw��A~��ŀ�A��W ��z��m��O��gfb�{��%R�*�[/��� �y�5M�Z�T��W�ݙ�|�=��l �	ȧ��fB�w4����$
CZ��X��G7D;me�ckj4�z�n�Ŏc&�*����IS%THEMN3w��� woU��� ��2�]�We�Q���F{��H ��o�#�rAP�e*M7����G8D���75/^ZH�o[��YY�� ���̻"�u,P�r��@��Dl$D�&C,.�rߒA"FM��$J�+c:���� ��m +9���Ev�U5T�)AJi�]_k�[�{�� ���4K�D��ʧ�Y=�v�׋�Vj7��C7Рǋ���Ѝf���i\���V�V��u�^o5z�����Z�
E`��s����鯼���f�O¢f"L��	�ăyͲW���uݫ�K���t����Ia��D�$���ۻH�>)Bބ`@��{0�v;SǍ���`�bءӼ�[o@ж����W���&(�)TU/�.��� �l�?6�A%����M�u�>��L��<���D@-��lxgD�2UDHT�)�������4�K�R����2�M�%��Ly$���ɰ��t�7v�\�b���$$�@Q*Ka!���z���` ��2"���7�ǧ68���i� ��kx���'�H$D���sP(�E�]��ϖGy$�j�%�gmݤ�H,��m�)��rd��m��	+6J���J
SNb��]�I [�˙8f�r�,�a'��v� ������zܞ�uE�z�����6���|�"b��0�K�Ы�w8p�E��4��2��e�wYs{�z���=�7OE;���Bkc8�{�l>	�v�m��q�4��À��n�!ݍ]��v5���qc:�;J#�7(.�u�;rr-� �-�l�.���Xnr���;�g��q��x�u��U�S�nLms�k�؞���ֻl&�.#ӻ<=yi�Vܻ6z9Q�Q���)�U����7K��]<*��,�n��n.��6��c�g�cu�H�.�-���bڽ f{.��:�s�+�C�S���v�u5�u��&�÷f[��ߟ?;��g���� M�6����ט  ����_o����>�H����@޼�fg��C�0P������©���"J�6�N��#�_y�%{j�n�$�9�H�@>���q������d_�!S�HJ*ٻ}�� H;�=n@ /#}f���h�볮#����ȌH����.	�|BeD#d����Yj<�z/�k���@ ��\��DB��W�}9��ǒ@evm��%�(؄D�&E�P�"PHd�0�E���=��|�F����D0��o�j����o5��ve����NB�&���GE�uph��t<a�m���7F����q�/��������)Mz{��ss>�@|�mP$���L$���"wm��컰�H�-�����J��DʕN��kl�d�W�7�*�r��=
kТ��`��d��"S��?��V.�R�L�<�(��嘘7ju�| n�㌀EX�Mm�Sɛ�'���^���I^����$Hl�:%�1v��i�y՛����H)S!_QU2�޿*"k�m�$��'zd�)�[�=� ��� >���^� R�J@�QN7s��}��Ί����dD�a�@�@G�������˼S�{���=if��U"x^���Pb�4�C��l�r�uصR��ʧ[��ͅ�ۄ�Oj0$J���6��ݭ��=�la�wҍ�>�����r+�y�F��]���h�y�ӳ��O!`���p+�ٲ�I@2�G�/Wz��{s1c5�U��<f7D !mo�a���%T�R
 *b�\�������i^�Y@ ���I~��ۻ�Iy+z�NoJ��K����J^;Z1&J
%D�Uہ�~�y���9z.�|q�*�)twW6,ܑ�`�]WyC:����:�40�|/�%|MXڸ�Wb)�Q��2�f[�*�*hNq�F+˰��E��M^7O#�I/!���^Wvݓbp��BBBS�S1����s���zl	 �,���@ =~���> ���]WFO�:�V	�v��]q�R$H��I2��λf�'�wS�&��a��N4o&<[�t�Iy$2�����+��;��v�*-q!S�{� E�B�r;l���u�؛s�[;�pc��kvR� q>:6���� UD�*���@���q=~�x��>ّ��Z�;v�T���C3�Ic��o1��O�(���2�;�w1���e̊�z������� {�<�;��ə"j�?v
�8=+�j%jGv
J`�L*��w�D�����/$N�,9�W�DO����� ���3�>G��͈K�+F$�H��@�.XH7۝�מs�]ޜ���^`����aaȽX����0�6!ۊ�����y"����zBg����y>�S���H�kr�E��J�3ɤ�����t{��㬑��U��F�<"�<i~��JǇ�K��:��Iy雌��A���3-�]<�hk�i��Y���՚��;y�����y� �,��8��Y��bܒW��RJ�0�J0R10o׮�Y:�+�Ot�G=�qʜ��2��/Ͽ���1uh�&�+!���� ;�=o�" #+|탼6R�_�����vt�j@�8�eAP&`6�k���r�b�ޕ�S���� �l�� �V���$Ƿm��#�ra�M��$�N�*(��"e�z��R |+�Q�g^�]�_z�D��5@�o��� ��ͦVuQ5S$�
�qU�����@뜶��	G����o�ke2�J���ݳͩ}�U D�̩T� Un�d�%��]�H�y�)c���om�n��� $)�y�@�>�dC��?���M��5$�4>��^�Z�A�U�g�C�@�gs�t✅���zkke��t(�鈼;:�w��H���<����:�v�m�yjnۜ�i�4[�<��ԃ���]�f�o���/a��h��]kɈ�*�
^;.�(���q�q���Ƽ�ڹ� p�n��ױ�!�X/W[ת:�[�u��؇9�o]C�-�&9KGNy��Y������:sͳ�	�^�L]�;"ֻtZ1�l���^����5ǲn�v�s�6�ۉ3��)	����Y�D�/g���\�XW*ɨm/CP{4���ݵ)���=7�h�7����9�/UT��E�ζ� @�}�؀���fA�i���i[�+�9�]����������T#0bA��%�wm�$���[�\l������eo��� -�ۙ� �k|��5�Qr��R�圐*�`����.�y� <�^}�� a��]�������Ͳ";_kx�*+��%QRDˆtk�SZ;���@�$V<~m$J�}��������k˝fV�{+�{���m���UUQ$�
��46�s>��"=�uu�s[3�n=D�s�@}�}��@��mYf\{���-B6~vN{7�=�;z�V��Ԝżu�\����]��!%H3��x(�F�''��o���'z�]��Iy%�����NV����K�!��ph���]�w䗅麌(!�L�R�qϝCA)�����"v̴8�]ɾ���ؤ���3{�������V���i����O�/{>��mFY�>�#,�ڛ�7��)�r��55���(v�m݄�H���ZVi���ݘ�9s�<S�wHZ5`D�x~�zI��$�κ�����=޷�;�׀����� >6;9�`�b9g$
��&��6�n{��_a����1 �=�D�vs�� e�{1�"s�r-�S���ѳQ*����"e�GE�J��z۾�O+y��-�o}������PB�Q)�-HfN��&"$ɓ	���)t/]�z
�v�ؘkl/�Z����ms����h�!S���b� A���t�% n�]ns�n���b.�{n��^H���~��1��F�%�"��lA�/�0^&^gk����7��9a"H�����'�bv�[�^���ǀ}���R����J�ˋ�nȁܿ4��v�htD��뾵��܎�{:��l��4�j�bo��(Df;��<���H0����knd�n�mE	Z]]_�:_u?R)$�����vd��)L�J�G{�2^����l�x�@$�[V �~�`���k�2�e?on�Iu�)!0N�*�3!�����M�v���G�������;�����m2�w����7(��Ў��\�@J=3��ᵍ��cxhuY�	�O>{`��j�.�N۩*;;9D� ��JR���V^[b�	33�n �:����<W�ꙫ�b����Ր ����W��S3E)
�i��l$�"��Vh��o��G���I���ݒO$@�ǲ��I r��D� ���
�?�?f�� uv�d�T�����ot��a(�RM��B����A%���dؽ9P1 #���|�%��/)���� .��l����fݒIӯ�s������z��̝�f����l���#�:ί��"S�B����b�H��GbGX�7.�;�S�#���[|����O�Aq���ym&���$T�LS!J�;��1aF�[�Οu�j�R`���2Ny[�!$����<�-�ӹ?>|��rv�6��K���<�y��_g����-e�1�Ԇ�%�����w��rW7}�Y���q e{���79���IS����'�[؏7kK;�wa(3~:��	h%������ �:��&dǸ�	�ӹ�w䗒@-;|����"	]^��&W��D�M)���"��s��s��d@�ڨUؽ��/��o@}~��@|���j�(��b�(PA5":i~�l��d4�8�@hz�Nm��ПĀs���M  �������ᐵ�j��vfg��6�E*!_�´�����M_nePb	��$�飛J*�U�ѝm�I#�s��E$�{��������/,�ۻ��!���w�|�75���o���!��=�%���t�Ə��ʮO7i�MҨw�����A<�I�q�nL'I�nT��b�MO,�>�^o[�]7�Kw:���\�� �Vfʱf���c1Wi��E�xx���j2��7�ü"�[�Ξ���Q��G�/��[�9(��<^;��TC�����QT����Xg�k{�u+]Ӻ��c]3o���lE���r�gD��/i}�E�k�5;�Sp=s�#�)m;�w7Gzz����?)O{9��/�x(ug�Ȣ�i����ڛܡs=vO+Α�r�~��9���#7��,�$V�Jm�<�:=N3M�*�Q��[�wV���s(��$�|��47��z���ܚ�m�Ρ�����^G\�;V*�� ۺ��D��ϳ9�2j
u�wR�z,y���]B�+��@�.�u<{��}_ٺ�W�d·��%Y�+��x�v�]W7�xn�ѡ�"�cL�귪����׮�[A� ��޿k����a�!�$=�yEe��M"�p�!�x������U��Ӏ�ϼ��*MA����ANo��dNVn+��r���n��l��ܙۈ����vv-7'1�k7|!�Ӯu4��%e!3Ѕ���4����W-^��f�|*wo<*��.��H��隄fA�qa��lu��V۱d�Nٌԏ)C*@ X�;�]
V���0Zz�F�v
O72�)=�}r�.���'M�$j��3��e��AH�@$��ރ	���F�2�+eT��QQs��9S�3���ݱ�{hTb�DpnV����
��ܹr���d�V((�S�[V�%Q���E%�"b�.qYs-�
���PX���«H��*�4n�UJ
�����Q1���s�Þ�9��v3�+�V�
�b��EeZ*�3)UT�,ki-,AYR���U���1JV�eDQD-1����ڨ�\j媢�F�U�dȊ�((֪���ac1,q��J�TQ2���6����*�e��f%DfXU�f��Z#�LQDL��\�R��E�0�%A�mdF�J�m����T��UJ��|=��c�o9�)��Vdq���e��.\�-f	c�re��mݻd��C��Z�`��8�9j(���-��g�z��Jb�c�޹Z2ٲ/�N�^�n<)K�v�K��]�x�r���hd8�̀q�;Y�ka��Sms=q�	�Q8n��	��r��Nk���	��}q��96��a����-������c:�TK�\�LTt�Mipʋ�R�f'������s˰Yq������϶���zs�&]v�5=������ۣ�nka0�[�R�����yH͸��/<۩9e;'eoB��m�Ƭb]uu��Hv�-�}�n�q�,T������{lo>�M�nH��<Ӎ[\ص7�7m�c<��G"�Ş�n��N1�xݚ�nu�� �'Bo�(�u�;^z��wX��;��\��$�H�Z+����scsp�e��܆�D"YYc;�Nz�<��|t��=xBvݮ-*��B�c�X8���7�Ӷ�<,9�ޮ����f��ɞ�qό�9�\�W�=����ͼYˍ��3�d���۝��[���"nd9�M���鞓��O������3�!=Q]�`�`ޑl��A�۶���a��qt��v�����VCU���5lv���5��y���Ҝ��.ލ��M)��(v�Um����lZ��33Ln�0���Vڡ{7qƲ�4�m�%�mA��va��+��a����%u���.��A�'���1�ζG>]�&>	��]�P�)�)3�6�v7Bܑr��ݻ��]=��k���w1�(����;�2t1�f�a,n�:���fzr!��kQ��D\ƌ��6%Lh���;l-�1wa�t��g-ciݲ����;gf�\���n>o��w?8Iv'�ۋ�\��:�;v�M�[S�s�A-�ٞf�Z�G���<�n���v��λ+��<�6��3��Fv�<��[�V�u˸0�8��n��9��.s�n\):7-��s�i8���.:�fݴc�T��/c���K�Os\�q<l�ݱם��`�����[{[95i^�6�ɸ�F� �g��F^]�^8�s�P:�y���m5��;n��]���˹�����L�Շ�'rcg��Փ�4U���z�vM1�]�Й�5Iێl��v:-�Ѹ��3A:�^�\[Y��+�hD@Nz�s��4�ö],�]b�"9�g���v��%f�i$���t�<v��9��s��>t�ÊN'9;Ve����.-r7ލX�Zw�N�[��^7l��,�g�,���u�1gL\��U9-d{6�Z�^y�u�`�����v,���Q�"�+���w������Ң`��0�K�o<�I'��WR%���;��������]h�}��H�0�s`RAH<;�d�
C`$:�k���K>�$+�~�~'ޕ�@8I�_�xH����	7!��}��{�=��{P)�����p���C@ ^�y��]�)�*�w�sۺ� |lu���	#/���]��R'V�@�����=���պQp�vZ &1��0#�x餂K۷�v���I�ѝ�x�.��G�v	D�n)"�&hP���5� ��=��d�M߫�bܙ7Pu����{<�!��{�3��w�Q{p������ML�(JP�g� ,x��e;�sRO;M���hѥL���˭����_jeH�L��|�z��$n^?6�'v�&\vg�k�i���H�$��ܼtXR�:d���IS!J���繋 7;�=+Lϳ�ذ���`�b�x*��V��DZ��UwV"�>Z���o&�;�0p)���w�d�z��	�"ID^��.2���o�������z:r+�U�I ���zd(�
C`��lH�=��` ��]ǥU�K�j+_d�i$/��Ey%�y�d�S�IBI�e(�;������v��+u w�[`��f`#ѻ�o�2#;j%�m�- �����)��R���RX�I��&B&�{�|Z�כ������n� ,��f`�=��%y<���H�QH�0 ĉS1�ζ���w �nd�{ucr�{[�K�/6�~�~�y4vؒ�
r���6 �=�� ��r�[����vpǂt�h�$�m���	'��	9�DD�d��(�u`��D�q���뇻�=��lH�[�����w�V@�}:�ͮ���~L
{;2(��QS%LSgw=�X  ��%��H�^qȪ��7�eU�P3	�k=�y�[���Q>V�m�ۨN�X�l~��wF�,WC��}�p{"K����m��>@)�g��fi$��w��JA�ļW�B��d2GV�vB��ol:QP8> ��kŀ i��XH��w���I`%]]��K�W%	A&��(����%�"p���j��^�][B�$����l,=��"�Ia������s�������:lB�#)��M۝cv='Y�ƭ���ֵ=����Ŷ�7[��f��K)#Gž���@8Vީ$�����/a�5F��qT:�w3 ${M��NG�I}��
]476���������n��  {gy�@$���� ���~��y�������FR��'鯪��m�t|�G������^9L�͋������Ӷ�T@���vE?N̊*iT�SMwv��Xc7](�ֳ�%䢖u1(���:i �����vmպ��N���U�$��~�%}	�nW�9B�g��gG��D��9�n�u8��_��mA��f?i���Eӂ�@#�n��K���+�%H�	q��$3���`tT׫'kIl��q� �o�	+��'�8�<<4�T��O���gp��6�؄�VM�v��+�ܳ�qnׯJi�ԤE�T�-}�
j"TQ&�|c7A�����b�3��3 ~���͸��r�lJ($x��0)/�ܑ"IIbR,2�}��%�}%=�=�<��w�� >�7<�� ggkq5�
|�^�#��K{���D�(R�q��Q���׉`| c���{���^��$:;<ݐ 3s�3 _?FZ�;�y_����a��J�.RCsāq^�Iؾ���o> �i�ɠ�t�:/�*{�@.3�ߩ�P���12MU�wv�f �w[T{��gz�㻻>��� �}�� ���`��rMv�;�e�ֱ�m��T��da>RqS�_��Oqj������5l�m�A82��/kl ׮ײ�ۍw��}?7ζ?1mu��E�V��]���Ӄ��s-5�K<M��'���F�	�S�^� <u� �no�qq6��Ӆ� l�����n:\p�ruu�K��z���Y�\iM�*j�Ds�0�ݪ��:����v�k�f�ͫ	9��s�F��&�텥v��38vE:�8�� �Ŷ�����.�z�c�;�<[\��^n(x�ġ	ی����pt���-�]�w=mw\�m���|7]�jy��|u~{��ߩ�愤H��KN<a�(�k�D�$�͎�,)�fh[S���e�{[��|�[πۛ���SQ��GE�_��u��쎽����y�> 3��f �F�7`J�'K׼>H��AT���Q��Ա�*����Wۙ� z7��'��z44v�$��Y]�݄��8w���dcĊA
�D9i2�c�5^\����  ���ϰ	����#!�>F�ke��ò���=������*3Ј��H����lR^Ix%��?:��]��*4=� ��{2# ��osj� ,��t���-����q��7V�%i0�������t$t��c��c�3]q˜��"�)i*�n����bէQEO��}�$"������ �3�4�y�]W������os�d�9zE�55Icd�OG���D���8O\��s������ZCg$�o���7M��d`Q
�^�Lk ��B[���!�,�/��Z5ّe���v���J��	$�/��� ���Ր �;�=�ي뚊���K�Q\�%� ʄ����9$��w�:%y"�����iQ���"R�́H�$l��I�]�"fJ32��WH��ܞ5n,��Oٗ"���A��~�J�Zn򤖒��v݆!L��]i3q�7}LRFE�H�$���ǳ��6���¬鍙�g��Pl�<�@&	+|@"��I	���}�}�������(���{X��+�Y_7UÍR��ttؖ�nl<6k���;o����=�y���/�&=����c3�; ,�����"�qf��ǆ�Eso� � lfs|B�|t�Z�j��\����&BP|Ε�o(�sU&�H$�]��^��ۻ�I-ݲgk]��Q�p�@�蒢dHl%��ߝM�v��D�czv��@����egt�.�FFe�WF��r��t8���0ٸ�@��U^t�wZ��Ni��؆U����#Ԩ3ʽ��z��s �9u�,��4tfsv@�K+�s3��zI0E"Q*,.-�2hS����j�2\[u-  ��nf��{�3ֶhpl����{XH���V�n����K4����_I	$�G����(�,yJ��++��C��n#G�{�پ�;�3�{��l�9�q�sZK�\(�EҺ�'Lp:�u�9^wmp]�����F�u�ӽ��&e�?��8y�; Aם�0�x��L#�]ފ}��4y�����ޒa*��TyH
k�U6�1��� ��+/p�b��J���e��h���բL3U~�A���tt�R^U��15D�DU6u�nb�|�u �ݜ�(TB�<��h �=��� Aa���·�Je(�)��^R����|�>{�0���:h"t>Ƅ��or��g^���ʅ�3Oið��f�Gg��"�Us.�Gc��q�EV:��j!>e��$�Z�PC0*K��A������T�"�(�G�wՔ�Iy,/��]����ݎvI��/o1 �>6;�� H����Y��$�[��}��ÿ�,M���fzx�j��h�ݪ�.���W�OWI׎v�|�}��Zc�6qI��;}���Gv�CA/�}�O�:B�S�"��N�]�H$p�mI~E�E)�1 9`$��&�*g�ʞrs:k��A"P���"O�Oԉ+/��8��g�6�	�8]$�O�D�7�z��"R\^c�A"_�.��d�v�lzo| ��6�������"���������"�����Ag��p]d�J�ԒIc��rK%v���=�
 ʌ��݁ԍ�TD��j����r�#�9����}�|��� �C�[V@��}ّw'':�kgϫ3�A�p�W$cǐ��+���m82!���i��k�p��"ߓY ��8>6����� 0'�h[������^���]�y�n�q=��� �c��I��&u����a:�!gwk<狻c�V( 9����!�XM�:��pݕ0��8N1�<v��9�v��Ku�k�v�xnW�w���cv^�K���Й�TMۜ��=t�i��VȽm�S�����N�k�{:�Z�A6�{mu\� iz��p��r��v-v��-�6�KQu����|�@�� K�<���s��tpg=c���A��cKО����S���+�4e�~����YƸyJ�gଷ�K�H%��T�Һ���s�]ģ}����u%�3[�W�^V^�~�%���$@Өh+K����O�l�t;;5�۾�@ �{�Q,����6;��}��6;=�VE-z�
�
f�T�t�u������ ���Y=�;��p,/��
D�7{�dߧP�r
(D�dL�j���fTv�ڪq��n� U�ۙ� F���r/+�Z�ĺ� �t}�7�t��:Qڨ�	�*���ۘ� :;�o�;{iV�b;,���x� Vf�f@��sb��j8l���27g�� ��I�&��w<�����-�θ�탬�.�[�i�dg�0aM��$�L)�4�q�:I$��9�~Ix$�ns�Bq0�2.�(Ƀ���Y�gnf;/�TLJf
$p��ؤ��##K~Շ���2���B��5Kyҳ�WY�1��,�<bu�٬�5'mKTdC�8<vJ��i��$f����T�qXsN��K� ���7a$�a���H�#�f��&&��k�ωKo�"�8�Q�V����! 
=~�������?|���A�|� 1 f�s1 =�uH��T(S�䙮ݛ���;{5X�ĉ���� ��h �}�5ZsF�e9U�^�%�m�Nu�p]��,KX#�:�I$��S�����w�_�i�N�ý���$�}��I�x1(q�Ĳ���?��9s�.��]���ݪxz��=;����E�tvݹ������f5,�k��<�ݴ�I$J����ɛ:��u���I���A���>��Ȧ��T���]?�ݱh�!NOU�������w�4 �>�Y [;�@}3~G9�'��a�ad$��Ά�ڲ C�4�� Ͼ������v1��S[�D�Yc^��j74Uν}�p�=�֙j��%�ĢV?+mQ� t�Qz" ՙ�uY���۹�kM��IV�*�]�i�a=+'A[����/qZ�=;<0,�6y��y�W�9��X�;(��uвy��{GL�BZt�d�[�u0U�_1�kR\Zˊ��nAV�Sz�f�5�}MM���K�opY��֓2����\�.�9b�:���Gl�����n���=��}QCp��7U�����Y�ۭ¸��$�i{�
c��
7�h�n�Jkm�Z��l�ud.���17��vL1�<��]K�u��]�h�VzFl;Ӵ����+�Q��V�j�W�y�ecQ�񘤯��܇2�:��RZ j�7]�s�v�G�U�R!�-�D���Ƿ�s������*Y��o�Z���J���	������E� ���bQ���] �4��Ɲ*0flx�p�6�λ�eQJjT�nJZ�{}�� ���-^��2ܧ�zH���m�����b5�qkH��Sl��k�%��oP2�� M��4#�kIW;	ñ>(<W������;9�lܺ��#ee�Ckb�qR{�f����H5�Թ�n\O ���iy�-�cX2I���+�H��9��5�#�5�F������s�q���Մe�wz�*�i��`�%��*��	7��S�r�nVQ!v3{<�9Z�`����_`o��/cKr��oG��E%�KE�}}�w/d��� W��y÷����xӾrR�-s�T��4J�eS
ҍ�cS���+F,U\)b1�Ҡ�����2�QqKk-��ŭ¢��T-�Ɔ3.�X��h������-
٘\*Q�T[h*)���-�U�c���)T1�DT`��Q�eW-����0Z"������8+33J�`�)�V�*�e(�*b�lT\Ŗ�bYiTU�TjU�ģSTr�V-��mī��V�KJ�Y��[���Lr�2�Ek)iE2��1��)U-���alA��)J�Q�%"([Aq�mS(�F�Т��3�Z,AEEj-QXeZ9j �"�Z9h�r�F,����)�U�J��UVbJ�˖dAr�,�\q��q�7wU�w+��l<c.1����F+���T����8���R��TP���֪P��%�cUETr���3+1U�3,Y��[h�)Qr��b�����{m�޾�[�a'0��[����$�8��ѫU�g_�;6LL�i��	$���t���ΘD~�f\L�gM72$��ͺJB��"��L(0�F{p:H����p�����g��3<�!����n� �m��3n��V��7|��-��~���ʦֶ���C�ە˹:���ݘ6Wgl�v��[��ڻ_�����߮1�֥UO���mX l?y�b 6�����X랃]��9n�Ԋ�H��68��}�V�Z5������zɐ��|�e��۬��u t?z�!���ۙ����Jl�Y�����K*PI"�*�RmF箟��v��O��n�9wY�{v{�/$x��b�&{;[�l�TL2L�����ߟi�7:�^�DP8�Ɲ�|����x{��<��D�l��ۭhMb��hZ������.�ҷ�����@�SVI��{
/n��i���x<�5�*T��6�=���a$�;�|J[=���X�V�+GnM��|H'��߁�{Ku=(�>�ϝ0 �������e�3������T}��xj��
�*εIѭ��I�&���nZ�*�����u������3RLJ����4�� ���v�Ia�ʖ�����b{XXn��XIGom��$�� ��H�"f[A޷%�C%�e����Ʃ��	�3�3 >=�n�w��`�7��9�M}%�R��U�n��.��������[� j��Q;N����bz7�mX}�Y*PQ"�*�Rl67�[j��+�� �cŁ�D-7���ȼ�7y�=H<�$ݽ��/�1P�
���DM��w��I%����D@Tr��4p�u�{�����/$��rI,f���F�.̐k8L�݋U7���C�؍�|$v��K�).�ε�us�by�>�5Y��F�˰�C�\�w
�4��t.�&��V;7�NY�D��v�r�]�x��|�lF�7m�z:j]�K��U�������c���jp���Y�q��|��1�N�����X�D�rm����{z�ri�9x퍠M��Y��ݪ�\P�ڗ��h�`p���y��Wnn�m�\T8��]��ݚ�g�]����a���@���bؗ�n�z��2���g�۰�'�c���������C���P5�y�
��c�g���X��Y�V������$�G�-�  ��DG�.w����{s�[�߀=�ڰ����TR"S��8���H�T�x�s�cgK�/n�[�� ��ͥd1:6�Q���S�_G�J�� SJ��U7�:v7A��:�$�)��rݣ�ɣv���p�~?N�'���Y�bՠ�ҰjГh���z��3o���e<@�g[T |����nfٙ;�X�u��K
���r��X
:sBA��>1�A"b�uص�w����7[�7�Y��я[V@�	Nwnf ��U�>��s;�TG�����n�kB�m2.T�rK�{:�v��ђ;�q�N��~��ts��f����!�n��я�NĀs{s0=2��A�х�{g�dSm� @L��y���uj�5$4j���w�~�0���:������)�s�I��Z[��o�陠�Q6����DFV���k�y�P�z��=e�����oSĶ���#�+�u�N�ڄF�� ��릀s�s""3�n���ǃ�$.�؎�d�@�X��e��>���A;���;�\��hz1�� @}9���[�*=05bL�F5�T����ı~�:$���vD��{\	٨��BɀHϾ�wU����QҰ�&���d��\{�����z+hۊI�1�H�';w3 @|lokv�jz����ֻ<߸y�J��NS�c�a����-������6R����gc5����W/�����u؄�V����n{ͳ�>	��n0 4��QYq�D\sS,fjo�B3�n��*Δ�1�PS#��o�Ȍ���P���w~@|���� �F����._z��n}j�d��iի:�ӫK���� z7�ڰ@ ؍�OH�匬�k���5򆍥l�?�S�bK����=�T���l��k'6I���˛��]�;
ۈ�N6pG�ۀ��V_�w���s����=�u��� ��3 �I9�;����H#s7[��A�ݷL ��9������OF�+��/�.�{vM�� ����$L�ju�H��;���+�����a�=��s3 ��ݮ� Z�`w������G߮��w�P<��U��-<�� 6%7b�A���<�(��fy�/���߱U"*b�1U����f` twm�a� s��K����o��)�o���R㽮Kep�T���!�;n�#�^�*�˭�{��v��	!���,%�c}2㜩�ט�kx%9���R�(��*Ǝ�zڰ�"�sl��˳��0!d$}� �o��	;�mY^slҝ��M*	��&�p�7�����ݓ�4��m+� �y�� �3�3��q�Ӆ��b�鵤Fj�u4��Y�5<����g��Ȼ��+'?'���Y�˝��z��q\�9�u�G�+����o��čnS�$=:a��Q�D��L,��� 	��y��^�e��|�S�r� �<��""s7��X9{
���t��m\�")t]K�^��v���v��%��&e(�e	�Nq�AI�"D̾
0�mP �k���+3���3������3����)�Ccc�/Tf�LL���TA�g6���A*=4&���Yt��w���,}���� {��j�oԸ�"f�ŀ����*)6�<�b��ןa|ܝ���m�V��o'����:� �3� }���j%��g�/�b��u>]9��ѯ�v  ��=�� #ѽ�9q[�$�Iq���(��"&$RAH�gz�I��=�����h��a��H릀@*���Ā@%�{[�!@�&{�.}W";8I�١�1z����q�f�۽-˅��t`⤵%0�~�鴲:�U\��/���i�+���'�a��" EAII�R!(��������e�n&��3Ԛݯ-�;z;����ŧ�������u�&��]��ڷ.�W9۱t^G�F9ΆJvĆ⭭�8pq������]��v=q��;uuv�������\v6*��+��M�tS׭�\E����uOUq��`7]n{vM!�[l��&�{su[���xzݥ6�.�Ƽ[��A�u�MƱ>�2ny;6�!�����:��Z�qPc�r]+��u��.��݋���~�~�؉�UQ+�����Wf�ŀ�	 �ok���:�ߝ\�	��n�'��HI�/f�	 ���j`�|���I�����G�x��s	*O�  CF��"J�F5��A7=�)/Tv���Q3%Sg����@|�mX| ^�"�+���h�U�ݙ�@�F��a�M`r�A2�"�����N{�my�ڧ�� f=����ۦ��H-/��Tv���}�H:pǒB���`W����P��*jf�gE�a���������.�$"]�ݤIݴ�(l>��&b�*0��ĊT�AB&>��a�� �7I��]�k݊:�.Hy��7/;W�޽sۮ��o����R�QSJ��29}ٙ���m0�����4�s}�j�i\�P����� �{[`�z%�B��Q5�4&k�����&�p��Z\�0�ʽ�wvP��jz�w��;��d9�F�+��q{v���φD�k;Yޡz�=-
�30�&��f�')E�k�h ����l>��""{��Q{龉��lG��D$TO�b[B;����Dt?y� @��y>�G^mϫ/|�@F�m6�(-/��b�5d��A)�LD*��k�ô�\؝,������ h�Κ@ g{�:zfTyB����L>]5���MA5_D�I������D��s�-(y&`�.clM�H>�]��cs�����f`y�Gi:G����������᮴ݏh�lJ�Շ�0�=I���t[إ��1Ų�>�oϲ[�6�%�?|,��l> =�; @_{ݙ���Mq`���r�[��"�:y�0) "�BR��R,2�feV.�|j�
��l;�$���e�_�@Wfu݄�Q{��h*�!�!�R�Q$�_�q�[� �����^��9�����T\��\��*�cj�[�7�yc��"{�N�#6`�T�Ԫq#��ئ�.e�/"g��>����[Ź�ä�����$��ʒZJ�3���/<9B1(�I(�H��B�u�� �*"��݀{��� {{�m?y�]�9�E$���\�7:rba T�%U7����8�ww���˯�k��@+2��@ �ٙ� !{{Ͱ�gY�;�Q"�Pؘ�$L��`A���@����ƞMnLiG\��#rt俟��M��i����I)lC��s� �{�, oc��!�7�.����RK�ݝw~HG.s
H"$�3
i4:�v�pf�3��p:%�f�]�	$���	�f��3s�V_G���g��PX�H#� �|ظI�r��wI'桹w��Y�����j退W��fb$f��i]y$��T	&�g�Vg<Ϊ�:< S~ǘ���l
�G��‟;�o+�x,��D�$�w:�i�����j8�I��-�:-j�����}�ٱ�t i�<\_��ڛP�x��u���'*o�3��>	� ����6�=��`�	G��AyD�5&�m�Iy"3{i��$���~���Ѣ{/��:6�
�*d��:ۖ��gܝ7b��4�mڶ�U��+q�]�n!^o��J!AU%S�v�{1` .��0@ >^;<釕Ǖ�����z[�vf ]ݮ�GDr�TUW�I"�./q�^J;�H�;�"[|��I�.�۶ #���Ր|�u�͸;���]�DH*fT��C���� =�i؀
r�[���q�����  ��[d�=�n�VgT�E*������,(�ν���p��$��hF�P@
w�w�a��O����u>�T�hvp��տ�ɽ�|�i;�"�E��L���)*��wj��x0�k���+�M�7�Ey)��l���G&a�����{n�Ѫ<�A�+[V�`ˏ,�x�����|PX�.#�Z]���\��{mܓ�{':j��Wz������b��;��P�޻2͢��3J��5s���ٹ����c_���F�g}��Y��w�N��l���N��lX�3f���Ҧ0�O*B�.�˓ɏ�[�t%���*�JW��㕛΂s��ְJ&��>@-�9�F��Vi�g��eA��NN8�_w�+'�⇡���EE��ݓ��z��q�Z�L�:vff��H�/7��U�@(T]U꧕��w��!B[�^v]�9Ӝ�em�(���\=|����Ɇ	�<&v��P���'��<�Ҍ�����ɏE~��n�X���骒�L!0�2�swb:,�����,�X��B�[��'g N胤Z��1�ؼ��E��p���%����߄7��h+ѥ�)�:k�|/�L���}�[�ٳDɓ��9 ���5՞���D��ۂyCx0���i��5�����W݇�)�'y��{�C��p�vyy���9���[��-m��3%D4��79hƯF����$�Z����\��d�q�Lw5�).HY]Sz����/�_r������L,{:�!�G���rC����uaOd�mk�3�S-��b��(bWގ$.�R����N�3���{�<]D���!�Dd��H~�{�9yE�6/WV;O_t7�,@g�]~�<�;�f�T�B� ��w��	۸b�<�yW��*&N�搻�A	KT�5Ҡ�f�C)�w�\2��I��I>HS2�Q�m�����TĲ�Ka�2,Ve�*ҕ�ʲcb�J��(��X(� ����Un\�e����q+Q�G��LkQ.d2�+��iF���.QE�%��3
5�r��1��W��4�B���0�-�0ȗ.!�	E*���X�\kQjW�[���r�b��̥2�V�kmV(�")Z(�ұ�2�҈�%�+G�Z9KY�k3LJ�E-VִC���
���S(��幙�Z5j���mj��U��6�˙TU����b"W2��eb�T���S�E\�Q�J�Ql��b6��5�P���+Q��mF!YVV�)ie��LT� ��K-�EG3"����"<�}�c��m�ve��"�[F�YZ�U��X�������b�aB��`�Zb
�4�1-̣Z[�������	��{v6���7����r�*,QDB�QJ�
(�5[Vѩj�T.fW(�l��c%�j�KF�EZիZ�h-�U0sۆe�ch���<~x-�of�Kix	�vn�s������u��������m�;��:nSs��Ȼh[)zm�W)9��x��s�vA�ێ{�4o=N9v�Z�0��Pŷq=��`3��l����C�#��V����=���\���<nI�������Vs��ĝ���������yy��ns\j-��vݻF��W�t�zcgC<mm���m�r㞳�&݇n����`�sc�u��WY5c�v��r�OIm۹^rFӵ��꫔{vn,���'m�o�%�s��a;d�Şv�W�ő�ǀ���y�3�k��+��z3�h�h�9��d��<�{=�X�.^�6������.t�[��svP���A�ZڽWs;Qt<� ��ۃsq�[=�`z7��]����d�*xɌ;�#;z��!+0$V@�e�+gq�i筽6:Bz��v��h;z6�.�@����c�p8�<ݸ{dZ�D��Z���p�pu<��c��9;<v���9k���/�C�xz���	{g����v!8�m�M��9�ѳu�*�c.��q���8h�s�ݱ �М�鎜θ��w[�WV��%�;m��ºb�ױ�<i2S�˜j�mp�SѢ��g� y�ƕ���x�
/c��#��gmv8���.���<���5�v�o.�s���]�<2���u`nI���PN�*6��:���A֔kv��n�XQ�sP����B*^K�2��A���Gl��\N�b�㗣�';��х��B��m�Һ�;>֢�f�t��\&L�Mcv�����u�/Y��twe��m%;�����fL�k�F�m�{6v�ն.;mqB�U�0�3f4� l�v��d�V�;cOg=�ͺqێ�V<L��;�h�v�G:[��Ҥ���S	�v�̕�c�n{k��=���:=gvw;I���bݰqȶ�y2uۥ�y���/�rm!�����-��\ݵn���F�\q�ֻ����ZF�Ǣ$�u�:
Ӳ'j�En���9c��06��˘uq][&��mv;�]�؄��!�;QN�m�nb��n8������#ϚN�Vl�X79�͵�E��=P����)q4i�;&�C�s՝J���\r����g:���s����s��n���wF͎*{.�we���a����=qu��;B���][n��Ë�&�κ]�d V��jvFˮ�8�˹x�n�w[��=�Q�d����`�Ǒ컮떍vX�n;7F�rޱ�A�ݯ�w��~��(�H���A��%�N�̩i�7��w�N�ZY�u�����T��>��	'�>��/FO�R�*$T�oy�g@K"&khTt]�� �gy����rB@_;��O���8��gq`ԊK�Q�� ̝���M�}3 J�L�muN�:��=�n� ]���*�e���B�RKx3��^����ؒ�_a'0��`��v�c{�W�z��"�q6�q�4��q�b���IZpɮ�� ѽ�v{��x�;�c�� �[rI/su��@-;�ߩH"c6꿿�����~�9}���
VuC�f$�]mUX�a�KU�sڕ�ku����z������ �E�H��q��; A��m0 7����&�8kN[lR$�v�0�ӓ
)J�]%o=��s<�n��g����o�tf�{�Y�1r�Pڄ.�Ƕ�q�|��ov?����eT�vw���]Ƅ�2�G{#��JR�mM׮/��; {�[@lwy�D��g:;m��0R^��8�)�A�-�-�E�"x��I$��Wk��9���ՠ$����lwy���8��`ԊK�:Vp�ﯺx�^�B��JoQi�k��K
;w��:;&_'��I��ߒ@�.�"P0d�T���`�F>i;c����:����S��� {��!���|ݬ�YB̘�d�!(% ��0W��m&C�G5�PTs���֫���8�v6���Ͽ~�E)��TLёȚ�m0 ��m�%f�T�w,�r�WS']S)�K	/!��豌9�0Q�R$�._�g/����DugUs�#��鄉K�l
EfJ�չ��y�f �:�2f ���&�B���L:1��GS�����jwn��Q'jp �Ϲ=��۾��޳/w�2��l���E��vx�[�F;�y�����׿wb��vuu�z��]:�I �v�a� z1�v���B��jaDʪl��}5���i�H WO��G�]0 Ks��sR�,=yך4 �ߛ`�r��X5"�����e|p�,�s�A���M�($�2�]?$�K�M�rK �sl'�Y=YY=i��ns(���s�W]{gф�����x�'lF���m�����u�i�D��w�N���TL��##��F>n���6��hz�!e��Ew���GM��Iz���"șQ�~Q��p��j��{~V |���"v�~Jz'jd���0:����Ü	�"L"��_7D��_u0��>=�w��^�s�{�� ��ͫ s��@�=S�	�k�$�e�s}��Sҷ�GR������۝Ͱ 6;������yn�IHjŵf��ygE	�l�]��x�Pj��ݛ���,2�77	�b3~����m��p8�y����Y�m�������Lb�k���i'�}9��2��ۂ�=q@]�xwNQ�;;[` >6;������o��٫lh��EH��L�E"H�F"k���g��\$�9���I�7%�v����?���e�}D��#���t ��a����b�Z"I�Rl�5C���xu���%Ks�����g�J*&b��:��a�K������7�� ��m� H��~�IH=�z�eGb����()��ME}3QRMP����| z;�ڰ�����q��=s�3u�� #c�VcN��B���UC��u�U���#z�';v��I.=�RKI+��������$��d�*�p��k詊��޻���?7W��E웋L��޻h�ۍ�G�|��~Y����g`������Web�?7@'b�!��-:TY@����a���sC�4$�Φ�+r(e�m���MJ�K��/��F�XH6,\�V3��[>7���Td1���gBǎ;F�p�9���e���$FV��u���F��.*�\ps�ƨ1����C/Lr�<7fi9u��wq��onl��t]�@�n��>z�$�q�b�Z}��b!�nn���"�Ru۷�n�DN(�|�-���k1%C��l�d�"�Gn�9Ⱥ����6�|�d\�<N�6w��w���	�'iƔJ�8-\��̓���=aM�y���B�sڞ�P���<�LL�b͝�uD��ӛ�P�@{%�]��&���z��3���w��T�f��U�&���ܒj�s�]��fW4�D��D�$��|�Kܟt�^�9��"x�⚩ED�LR�?�����|�N� <��=.!��z ��d |{�K�7�1&}&b"e2c'�t`1������z�.က]���|ݞ���e;Ȏ��'BK�uo:/s�HB<eH��&�>�)"z��������ʫ0��۶����DC]�����.d��{;=����ԑ҆�R%&�]L�J�b�76���R�it
�z��l�����p.	��*b�	��` �/����m�A8Ś�G��[<\,�]�@�F�|ؔ�9<qB�0L�b�=5Ձ������>?m��k��s��Zcv�T��:�V(����/��^G>��}�hq��Uݣ34VXU���4,�ɪ+מ�[v�ݢ��[L> ��|�����;b�oS1FU?2;�� ��**	�Vð��� ��i�� ����wLS��ˈ��_[� gkl�6qMT��`&)K!s���������#ْ�A���t ��� ������ůVY�}9��ݖ�������SS%Qp������m3��V�^d>=��@óΘ���B��m2�����&�x��&�~y�5m����;ӗ�M�Y�c�:(�}��v���4)f	����HB<bLJ�r{�3׍;77����F�7m��K�w�vq6;X䖕�uQ,=3��%R����-�W:$�M�=��@�۫�D���ߒI�]L4PK��[L�&���m�'1UEԴ#R�M�?s��� �z��� �,&�\e�տ|x�;4c�mە�[�eeÝ��=�qӽ�[�M�[c,M�5n?��^�U{��Uv�F!=6�[Y��59h�D�ԯ6��~�\�3y����7e��\L��L(2LD�O�Ƚ��8+���"3��` ���G�_+܊�j�"��*�r�j�"*UL�0u�6A%���,���պN��l���[l��F>o�!z��W��Z����-���v�k�ծ���7g���<�9ͮ��}"0ngD̉�@��S*� ���-"Fo:a�RXm�KK�SP6���E����@�Ͷӯ"��蚉�P�q���}u9
�[%��{|[�ߘ$�}��q z1�jȈ�8����{�=���@J	��
T؟sm0 :1�� *���w�����[X�H��t�)#��S�����B��2�Uu;A9�xq�b�$����$}�=t�����϶�)j�SU�N&�yĨ��p����*i��W�m ��;��m�u�:gEn���'.�.�Ӂ
ؚ��{V#�!
����/�*jb�L�l6�rK�YٵGGJ�ћ�z�O�^;�ΚH�yOԉ(wf��T�����Qs��Z���t8��.�\���GUp�Y�m�Rt�$�Bb��0��$7WTx A���v �����~��]������Ή%�f�6)*
obfD�"`�*��������,�7�����>t����� <�=��=6�=�z/1�m�����9z�� �w�m���ά�;8ޚ[��~��c�v@�[ۭ�^��\�%���'�ܸdb�4v�#���b���m��c�1ު�uu���� ����!9#2& ���2���ߚ^H�ܶ��W����r�b5Q�Ο�$��L$���tڟ ����ޝ̺G*2;t��جTwnS�j9���9�(ֺۡ.��;���y�/tFʓ�L����$m���
������.��Yޣ�s>���9�p���R��J�|��elWNݸi�j�\�n�y��n����vCF^��b�7m��tn�1��e=M�Y(��� ٯ7m��v}���]��vbUs��b�m�UF9��v�h��+���y�Η�����m��m��ܻA {;G5!����q>�n84z�κ�uOn:�vnHӶn�\�qX��6M��e�y���tu�/l���W	�v9�P���=��2q���@.��06��������k
%%A������I����I�;ݎ�H�P�5+U�){;j�H�-bbfB�R`@�d�u�G<��rFR�~]}�?; ��owfDb��� A5ﶫ<�����|����f��}3TEH��W_vg�  [��i2 A�^��.ׯ�u�{{�0�gca�l�A�Dx���R�x��}������ ����[��i�Q�w,{�I7��ݥ{�%`%DR�b{ʹ��A�=n�y=fV�q��J~�{�� ���m2"f'͉S�"ջb%�6�H��3$�'Yu����4v�q��-v&���u�0\��;x����S��"����{31}��!{2�� ���;^�������;����	���@-�\L�3 �2ĆOR���'}0�P���h�{�ݮ��m ������qw�}�5U��26 ]�sm��E�~M���}��L�|f^<�Bc�`�t�T�������HQ����z�, G������t@�_C����Ȯ��H�kU5T���(UN��`��tGVt�t���٧�O�I&�}��RG->��(L_)��
I�L���|��Y�}��ޒPI;{m� �/�X�n�fOd��tw�� �C[��F6�#���S��u������a޲̟N��S��7L$I�Oj	%�����+�|�o�������;�
�.\n��A/`�o#�u���u<�ܼ6:6ڴn�e�����ݯ߿��������{��`���N� n��x
���i�f��
�]]���=�@�}�M
�T���T�:��b�@Mޢ+6���cw� ��_���@.���π�3v�\����|v�TA1J*i7�k=� ��x�K�K<�@�ؚ��zLKi��ʐENT~Wa�/�1��dL��u�B�el�.��P�;��H7��� �j�;�4��2p�O�q�6��z�,8ME�o��͡aB�G,�k*�N̼F�T��#�Wqc�c{���#����ZĻ�YV9ߐw��1(r]=��d�^�l"��:�}�Z�R�۽���ݙv��(@�	����w} 듃��dnYdC�U�NǱq��^��W�=@����w�rK�8S&Q��u� Nx�Wu>��omMx�-p�pK�1�뫔�P�"��eZ\�M���r�ǖ��R�S���L��*KEy9�/����n'z�.��U�gI��1 �d�ϲ�����j�os�M$f�w3�X�H9��]îP�'��.W/W�������p`Ŏ�?=|��y��,Sq͏fsW>:3��t�C<����Þ�wS�&ٖI��L�����#�C=�l��Q�~���U�Rbb�,�xO�B�s�1�غ)�����(_X�.�U����o�ٍxZ9,��7��}/�ڽ�+��G���7<��&K�[C��X�-��AqP�M.���]۩��
yx�[��e(���7����L=oLo�v�n�{=F��J����f�f�����u/����U�z�Dn�W/�9=���{M���<t��
�j{f>�P������$D~�쭽�bt�v���px�]@�JXI�����睼����7�e��d�OR���lL����20/��)(�ꫨQJ[�hk_��e�*�iU�b�j�*�(�������R�Xަ&Qm�&ƶ�*�T��,Gff({�����s�0 �ȗ-p��q."�`�q���e��n"�6��T�L1b���KR�F��Q���V+kkE������4�-��-ܷ)YF�j�����������(���ҥmJ�h�h�s
LF�n8`���mkl����%��e�F���.fbQ�m���.SaR�U�Ʋ�Kb%\��J2��W
,�-
؍�iJ�ehؕR�ƪ���Z
e��-�E�q2�A�VFV�Q��kDPB��(ڥR���U�����V�m(��إ���h�JE1̫��ª(��b���KTX�#[m���lJ5Q-[Z6����-ZV�Z��X��L�-�"��)E�R�U��D����--Ym�f�[KUkm̹iZ�eUEPU�R���F�U�J��l��+QkcU�����҂��RƵ+k(�K1¸�-j��[hօ�eʔ[m)J �jQA����e��U�Y[V�AE""-��|��n�T@������9���ԖKp�ĸ���f��g�|��,"��ٙ� ���2eF����^�T�߀H�/[TZ���T��&�,���z�PHm�S�Lڔ慠Z3#�!�K�go]ߒ%!���<��GHD�\ h�H�7�KBP�����f�V-��acs��#u�]�!y�Ǯ������]���`�2��- �w��` �����
�q���lf�zy�D����Oz�"PJ���T���� �U�s�U�������{�{3  ��[��hW���7ϡ�T��?��sM
�T���Tٵ�30	F��Հ6}��[�����b1v�7��:;�m+n�U)&)D�&�s7ٲ�[�SE�|{�" w��` c�릀@|{�N鋊�Y5�W��ojv�45��&KRܺ镕��
���0 ��ι��ta���-���}33@FL�S��)��ֽ�eG���L$��x-ԳN��$��|:WP��9�[
KU�ν��{�3�7����F��ͫ A�:ڢ�n2�
�����[��n�p�T�D��C�\]������{�����B���,;��{�̿nf �{�P��d�9�`�+�ھ���^\w1�J��2�B3J.��9����3Y|����ַݽ��}�M �G��s���Q�r8��Vo�zy�L�L�dKa3��C��kt ኲ���Y����� �67|�!�>=�sj�T��A1U"��T���6'��jwd.<�κ��,��r�#ۻ�ޙ��]{���,+�\L��D�2D�������<�W��s��{ i�� �y�	7����'ݸ�淑��c�O�y�M���ډj��w	*Y�n#��!{CU�'Z�L�D��,���D�z����z�l����Á�w����~X9s�+�^��y+r����"i'�9�8(V�]�6M��\/NÃ���{Zw�1�m[o<-��W�n��rd����t���wl������펋��1q\]�����zń�gY�Z�k��ϔ�v�f47�<'M,�y�b��n,�|K&�{�tQ�k�v��+����F��E��"Ga^1���r�nûv�@����7X�&Wk�l<�����Oi���q�}�}��j��B�*��qO��X �sN��H=ۼ�GG����f��w��d #��n��U=�&�!D�TAƻ��X��co޲�c�X�ϐ��O�"��I�{w{3> (�g�j�Ҍ�-��fr�#Ќ�S�	<����$��y� [���y�=�ّ�]]� �>nB�Yۼݤ_B0�($�L&{�Ñ�'���to�H$�!��@gn�f@tv��ɳ#��p�'M�td5#���n$�~;��I |=�Δ���O�̽��o�w.u���o]�π����j�Ê�-����Y��S���u� �L��G�m��;sq� c���vλb4/O�"&{9o��3b$W�%�fT0����0>�8���?OT�7u�T������v�6M�Q�b&`�I!�\j��a'�zvV�%���apf
}�J��r�u-5ڈ;QA༹�z�;�d� �}G��QgڃA؃W�48*�;¡��]��`��ue��Q�($�������\{|�V@u�)�]�gfm�S�"h�B����1��c�@�{�Ղ "U]^���q Y������:���7B�������K�}}^_�؟�"^v<X�:`|�3��z��6o�hyZ�ē=�9� ��ɥJ��q�۰� �3Zt�<����A5ݭ� ����3��D�߯�? �3�|� �Txب�pe��� $����m�&�Fns�v��M?��ZâR���:��b 67޷`@{'9�A�s���fvWa�z����y�3p���4���L�m3|����}.�����n���@q���3�� �D>��W�>��� "iϵn��wsS�:V��I�ϛG	8M�%%z�5CР>y����v�^�S�㣴�^n�&�[�vtU	�x�S�#��Q޻�~��?/��]=n�{����9�,�H�I��n�$��r��=8L�H1AI� ��������N�0��[�a� }�9�X��ٚgTx�5T;ۨz�1J(��0�q������>�߲�ʚʼ��8�7L�636ڰ��fo6OF�F��U%8�T(2�%nR��<�C��z�l��Cj��;�e��vjB8�""H&D�	��n��H�635�b 7��o�#{h��"�9��I8~V���C�!����n)l.�뻴��Fd�w���`���H�x��KH���n��'ſWJ��K��F�po����2@X�B+Ս���^>$�o��s� vON۷�\�����r�^�ՠ љ�Q���0��r{�ZRѻ���Y�����q�u����@ ���̈πGG:���>{����:y�&�����-X' ��xn9�z`�ڝ����W-����3��M��/1v�&���*B0l�$ܫ��)P��&�DJ%&Z{��� A���Ջ�!DC���Ofo7`$���v9$�д��b��x�=�����x�ݵ��sSQ��uص�s����3����d�2T�	L�&z�g���� ��΢/�0���p��,���I~���I+�HE�$DB�Ȗ�3�ߩ$��"�xudڪ����1@���:�h�6�{����yYFa�
�U"�U[�����A�{�h �o����LN�>����l��/�mv ̉D̅!�ƶ��b���$����̈́K�t� ����m�[�qHOI	9������� ja��u�$�����4��Zu�i�ىvgcv0#�}���{ͪ/Ϫ�,�xf ��m̗����R�W����՗�|�[�N��	�Yvo�����-F�ud�b��Y�5��![�0��)�:�J-�� .vxF;{C�U��l]���p�Y�p�Տ-��r�Gk����J��1u.X:�z�����#ew#���vl��q�����Cuwd�,{@��;����@K�x�R�.��Bs�����q��Cn������:�2oBn���9�m���s�0����y���ƺ�ml�;����2��{cT���;���Mz��T5��ju�Ohk��v.��������[[;k��������ݹc`��39�b��ؾ�iX >�d�r��^٠��lLF������[��+���d�&0���O�r����ȑ7�����Ǹ �^� �7D;<�H�3a��1��p)�
�̓J"�7�⻛V `���  �}�m�E̿= �E �>sꋵ�d���0&[�ʎӺ�8�dϼ�A���� �/��� y��q���&��t$���9,+���2"�U"f�a��4��}��t�e4�v�Z�ۨ��`�ڢ �ޒ>$�(�������Q�sF�p�w�e����u���q��ζ��Rz�8�?�ߪ���2�IN9##��Շ�`��B�>y�٘
�algj+sһg����VA��s���V��b	��
f��p�n>���BI��}6TL�s�Cݨ�Op�=��}]� �{+�r�����(�ѳE���{���t���]�����)wE<%DWN��vkc��@r}�OG��K��2Iwg	$��v�f$�NK�u����*�+��HT��@H�4��'�� >��y��3���v�w���y ��[R@����fg�"��Lb)&f�������ee���B:�@̜9 ������uW����S�Ȉ׷��J?CPC�"4-�K�K﬐�����OU�F-&C6&����� }�ّ:/�ݍ���Vym"���+���sd�����W�Ξ9{\���.�c�����U2��E(���ID��!����A���0 q}�O��V�6�q;���7��\6�W���ݤ���F��P�H�!K'�M�RA.�ɓ�g5ۈ��1]�"�~��f ��}���Ǟ�5yY�G��(�$iZ �DXf��٘޷a�D|��Po:YSVg�$N֠��FocVn-t�{�(��v��m`�1�dU4Iq�-EW[�M�>.�ws�Υ�g6w�wȺ�׋��(��wh�A�]�鸺GD�
D���L�}M�Ffq1]�	3�{LH'�ExN:�s�Kn��G]�*�;�� ��j�(��[)� ���[��`N]"5	]�7�I�@�q��f!�^򗃎W���`�Z�v���0��͌m�.��d�+o\�y���{DrS2B'��f��$L@�`�@��7m�A �ʒI8�y��GEuOI�z���=l��A㕔�kY2��0�Q�ζ9��l<��ˇ�����V	 �]Y>����[�w9bj;�w���F��0%R��9�^$n���A��1Zf���ZIrr�q��`ѥ`�(���|�B#���xaE�'Ǎ�$�N��� .�����&ˠu�2�h_(�a�����E�\����y���y�����A�(�	p�{�z�
b�ggGn�I��$*"
R�_??e��?��݃%(�خM�	�������<�{ �Ãe ���iW�q�ԩ��۶G��=rY���g��m�6�7u�8�bA�w�Ƅ���D���hI$�{�A&�{����<�n�ܚ˽�mW{�������&���o ��ҍ����3ے'��c`�E��6	 ���mB�j��$V�d�R$O�FE՛m�v�$z	հ�;w���_��o7�nh��J&�*i�x�cV:6���@���'.v��'ow�$4�dg>���N�A5/5�$FO�LD��7m�~$���(	�[�&v��%LHU@:�=�����$��B���	!I��	!I@�$����$�hB���IO�H@����$��B���$�	'�@�$��$ I(B����$�XB���IO��$ I?���$�xB�� IN$ I?�b��L��,�N�zW� � ���{ϻ �����>#�  P@  
( (*�  

 
U	@ U� �� �	P P
RJU HIEI@U@  P  *J( P( (
H(P)Tn�ЂR�PH�$�EU
�R� T��H
���Q�)PH*�PB�*"�RRJ�$��  gB�P�I)�(���w*P�jUSwt*�\����7R�VlUrҪTrР�6
��R�:T۪E%ݹ^� �/� `��R�fUU��x���@3`�T�5R%ݎ%Eݺ�QM�Dn�wuQ��$+��UG�{�uA P�@Qx��Q*�
�D)ET�
){ҔL�%T�ەJ�f,ڠ	��%�E*ݺ�f*��r�J�۪�����;�U���^�ux0  ��   �� >�Ɨ0  q�$�8  =�7����� � �0Ҁ�x�<  ���e��9� �� �`�  �
 To�  xPQ%P��R�"�  m��} � �Xͅ
���w�(�*�-���J����W`��q �"�p۩(�c!T��(�  �y5B�}n��p����6AI�af�UT��R�0ꃝ7w$
ݝ"#��
���(�|  ��QT�*��RA�P�&B�ɤ�2�]�ʒ��\�s2�����QN��2ª��(s�XTQ� ��  -S�ê��4A]�T��T̈́�(Tb1E[���3���m�����ꈍJ	U ���᪑*@�$��
 �����6�n��ɔJ�j���(�:��[�;�:+wtT���"�EWuU,�
�݃�E ��  ��h#���7�R��E2jU�ઋwtR�6)%YҪ��QY0�S�rU�9E	�����@   ��4RUM@      ����IA�`F h�� ��Rf�J��A���4�@ OĩT����ʀ &@h &R�T h@    $$h ���CBjzM5='��#1&ړ���O��s���Qx��HH��Z�/�ַu�|y3-�H$,	Q�C� B�O�1D��$�!>� I
�F?͟�2/l`��m�Ͽ��7��y������8��`v���|�<��llg����0m��M�À�
��@a�	![���'q_�5��|�����I	T
�uR�
�T|�5��h䂥�j���$r�&�7������ժ.������Z�3//J�����R�aX��1�l[�S5��d�3F땷�Ud��$Zu�1�f��1�`U-Z$0�PQ������1�,���Z�)t�nM�Xi(�\�u���k�����wB�5Z(Ă7%ٺ@�b��H���cw��t�
(R�� ke���fR�[*�D;QVaPT���n��^݆E���Գz�B��t��	���c77�
Zv䙂ѧf��f�U��ő�;�T�X�kg[7�=��{6�2M<���0�`N\834&�:n�Ʈ�2�&,��Y�x"7(\20Z���<bM�j��j$�D6nn���*�]A-.���E]�m<���Zzn�Ǘh���8�����Zk#����fe)�UJ��ݻ�9X�3e%�/u6��v6PE�o�7QU����,��31`��Q�/sD&ӽ1�a��;�ʱ>�x��k��y��z&�4�֜��7�{Q��p�j0Bys-�w�sQD&-k{�hH��b���[&�wv��_�
բ���Wl��U��ޙa0p���^�Co1��ލ�� �F���ɶ[�9��ʺ ��t�n+|�ض��|�x9&p�e�N1�*�-��Z�k7M�3X:�k�of�+Ȭ�pa6*�z�0� ����c�%���u7.��M�iޓ�#p����OE��L�����R�z庸��H9�%�s�r]fL�h�u�v���n����;b��c�%n��t�걢��K��BPX�ۼ���1�����#��Ki�r"d7e<XG�	���If�ث��f�U�$3Y\�`(�?n�!��ۅ݊X��Ne ��t� ���^�)ҹ�K�Ko[٤<)�.�Z��t��zٽ�zE�b
��t�ʚ�7$���Lk�Wx��ܠo֞�-�Q��]�,5��%�w3H2�N�B����[i�o�l��n�
��1&�x�T�M��
�NX��M'����1��嗹Q�.����7�֔�/�ٚ����+�@-������xJl6"��(S��	zئ-��1l�н��'�;)�u�$���2�5�U��@Q�6ql@Ve�h��9��cFZ�v��e����@͎6�p�Q�� �[�F�r���+��M�C�J��6�+���Y>��o�Ғ.�7݀�vi,m�Y�o�)Y�f[AV�!B��#Ȫ<��d�@LG(��j;-֛yl�.���nf����C�W�Y�d e:sf����qe��X�Lj�ˈZĽ�Jm�6�mͫ۬S��d�v86X�b�#3�owBV)��F�Y�#�=-�{2� �S��Ͳ�cr[)'�Ù�e�w��P�a�fYV�|,�i���^T5J[�n�Ͷ��M��'G��,&c+�G+��y�sk,�nX�@��9��f������՝aʒw)",��#	�P���,�9��J�S2����Gt.7�Q�4,CVF0�[������8�MسLW�By4@��b�X%8Ιb��Z^��>4l����W������i�p���8A�]��Vw4�hR��")��R,Ϛ.�tQ���w�k&�F��U�y��Fh5[B�6���"��@���w[&EE���? �Jˢ��1�@;u*Ҽ-ѫ�b��X����#p��L*�ʚ����WY��
t/&퉥�"�	X�n�����鳮A([V���`�-f�q퇭\�x!�t���3Х�{Ww�C�EJ�g0l��&�@�NSl�>"�79�!'W/+���,k'�P�Ku�nZkf�X�.,L�k�/Cf�T��#!�w��ɣ���;b��[f6)\�u�&���j��,�%����z2���]KV���晨�4�&Vl�wwЭ/��:�������J�����sU-�
�m�U�m��&p&���.���s.,
%�ڶ��M�塱���t^���bf^���-jՌG.,�����Ɂ���U�:R�e��I��Η�X��4��;���'S#���#�rՓj��ƯoX�Y� p�Oqh5�$�P�h۳@�
n�5�aP�̕Y��b*�CV��R�Y�T5KD�2�-��i�g ��Uo]������d#u�+i�!�U��� `�+`5X+�h�W����"o2sR�l�TyKlAV��;ڀ���r�<�vPx� yH�IЫ�+)�1�/e��
a��r���ٴ>U0� ��a	N(<J	�7��Smh�ݽ8ᙠ�c)2b��a!p51���R3�I���O�1ͺ^��D��t�3KyH�
��ӻ��4�9��(H��f�=�KcrͿ��]�`�2Z�n]�K2򶓶�N��o%��Byxv�!wZ��7�]�v�ٷ���L4�絵�����
g@bFݚqok a6��nЬ�kq@��\�mX��x~ݸ�X��%<!̻	��C<�1��9-�SIRk.�9�5���],�R4�K0�m�mU�F��
ffc7bY��V,�<������P��h��U��֒-��.9��*��ov]���'v�e4u�d��xU�xUfDd��In�A�1�d���v�����u�6�59��e�Go�>x� �ȵ�����;�
��+��Q��lf�J�������L������3^��n���q8"�kI^�Q��{[�1(p�Z���-�,�J�%؀r]��6^B��q(R��c`��j˄F+^m$U���Ͳ�Z� �A
�:M7��w�U�nVh��ݥDֹ�&V��B���ٰ�RK���opV^ٹ���9��Jɭ*�q��W-`/\��5�B٦��q���61�y��ŋ3^�ː�-�\�9^��-�hNa�wa�X/��$���
VȘxټjT��`�8,����q��}e�Z��p�JYYHcR�F�[����j�Y�u�+�<ѹ`�,^ ��C��cS�P��F&�2���Ru{�,]Eee�	JCm�&��
8 ϔ��P|k+0�j��ØE�H�E̻x�����Y�Yc2Z-ҕ���Ӭ[p,���;64Í�t�gV�.�V��m^�E+�Wa��Z�� ^F�e9�����.���[Yw�ˆÀ^nL�0�#h���ͭ�I�7��ށ5QP�,m+�ϵ���ͽ�m�V]�d�V��]
ɛ�Z��x���IKNK�T«ws-��-���sM�EH�XU>yGv�	��VQ��D�	p �V��1�A�0��ݗ�k�,��9{�y��2�3�w(�G�h��b�m=�k-��2�	pE�4^0�j�����'5��N^fĵ�r
�ln��++/K��Ǐ2��y��`�q\����tJȨ�4F}�ԑ	�D�j�KN��RM�7+S,,IX�o�҂Y�2^=У.�Gu��r�j��(�u�q��oDsnȭA���[��;�@��̍ U�qhل}�4m��Y�C���͍cѶ���^Sٙw�F(�&�!8r��Ȍ
Xyrrf�$�3�W43f�#[��Nh��i	�1;����J�>�Q�^�c�m7���1E�v�mIbeF5�Ҕg.�0�+��E�7	Zf(����0[K�Jw��YN���4$2Z��	x,���@N��MĊ�v�V�+�ì� �2{wJ:h�ZN+�2�@ꊥh�bA�6��鼗��ͬU-�&�.�d\	�E���dR�]Y�1zkw-Zafǵ�WM%-�g%Vc��*�E.b�tRv�T�U�ӷ�taۻ
�le����*s���k��wZ۫n�mL0��U��qMʽ�v��{[v�Dd�Se����P������B�K��%��s볭�R��Š�ҽ��`��`�&��[���h�n�TV�ۊ�m�"h%�^U���&��Xoƪ�-Ҋ���Z���g ͐�~�I:2�sf���Wś�#���<6hT�ʫIS��ҰH����)�:m������rm�MN��,&c�Ȫ8u�������n���r��+E]i�ԌM!q�r:E�F$�w�Y�W*n�
KAeK�Y,�z�ɍ*�Y˃2Ѭ�*�*m���[�&2Ճ�@UK�1�YB��-���n��2��(Sܗ��S�p%��A}�l��^2mK01aÄ����V�"w�݆����F�٭�.���ŒҫՎ-#>�]Cs4�r\��Z�4Y���b��aNnD*�dE�(N:p2&҂�Qݙ@�w�����qй��!Wd^"JA��V
�5�^�n��R�HӔ��r�a�E��Չ�q�E���jGJ��׌ʲv� ;-C���zc.����ņ&�TNB��kq��b�$��N䊤
VH�� �H�ra˰F�W�ɁU�
{D��`�ljKY�y�Z.��6Qi�7v��j;�nUXOi,����F�J��y/ff�d|l͖ڥB���M#�\(��M%���H0�Z��[�����n��5�x�l����3j;��U)�}�VR��X9YI���2l�@7�0�srn��;����x�7p�p�����VK��63���JP�j���d��S�bmVAl�n���	��Ʉ�[ˬxn��¢R[7Tl�/Y����@H�d�a7[,ƈ�:^cq��3X�L� H
��V5e���Z4�t��*ځ��{P��Xa�U"�m�Wc@`2��ѹN�q��n�Ó�-�i�s/qd��m�0V��⍻�eH���|޶��dUq���l换�[���ePpb�;���
�2�������~�|[ke�@�b�{f�`ou�܏k�� Y�&�.)�e�w�j-���[�a{K��x/kaS���ww�\Gt���k����Yu7T�!W�h�t�ҧ1�,$�\�h��7k ��������7 rnK������A3�f�쥀�'j*1�wYRaa�[*�Ԟ#S>.8�R�wod��E��'��QF��ܧ�X���K^f�ؤ��cJk�Vhf ����ҥJ�h������#)'6ⷑ�9"2n�.��Ij�d�.S̖��i
ӵ�R�
��Ѽ�-Bv��@��kv&@Q��J˖9���tX���q�VIM�S9$�4�:��4Hp�fC0�%�`�R�u.dyeA6�$�q,H��E@F�ؑ�*�]โ�́�̛��!3i�Vʹi��Sm㶫ob���ШK����v���l59{Y�3���sr�8mY:�O(E�)R�6�d�]E�c)Q�^*i�	@N�=�Ճ,��W��m�[cfdR�����D����K�A�ј������V,�R�M����3���a%�ea6P�ʫ�h��.�L:�����ĭ�"z�`+6�92p�&�nMmcfX�i#@$�v2"�
���"A!D�.E�L!�(�PA�I�y1,��b��-ә�n�t��F�2�K�J��6�����yA�u�-�n%�K��E@�4�>k1\�MDw�P�T��ै���P5/	��f\�oR.-��W����6�^]�׷,a�f�m�`Yhݷ�f��l��m-p�j�e較5�L��͔�c�V^T��f�ڹ�.��H+`�H�#ul��W�CiSBV�K0��T�4�{&��N�`�� �.#!�b����S�l&���U���}�vSv���흐���CFY�d̳Y$'�����z����/5���O����a)�x 2F�Y�-�GZ���Z�GZ+oٰ���`J��r!�K�x�e�oEm�2s��h�x�FD�kV��a�uj�VFBu��5V���z^���6�۠w6��(V�.ڦZ��{��o�e����Kf���l�fC�h��N��"�Sr��oF��.Ṷ�.jIMn�+��6���0lU�v�BD�c��Pt�}w��(R�
 �X�l�j:�k,�.�q�A��K.�qU�T��C�sZ7,�Z�V�1[r��j1Z�v`ݜ8�,�U(��,*9�Fj�jF�\�v«FKȝ n�Jx�c1R�ԅ:.]�d[B�-69�NRڱ��ֻL�i�I ����>ߎ� �4�����@��3�03T�0aK�a�>�J�yҊ	�H���~�,��,������߁�P�e�P `?e؜�@Ć�m;`˶�P��`˶)�e�Cm���ci�6'
��M�� ����2�bC8660)�0N�a@��.��.��H�v� ��
&��c���� �.�8m9M��cHm��m��c
M��m�	6 \Slbq������v��@0���6�����66]���]�v����C4���N�8�2�S0`�6�˶ �Ɛ�i�.6P��6�X	�B�"1$���~���>�F3��1�����$���/��Vn���[B$����R��H���9k��@H_����CG��� _�W������E��k�݉�u�0dc���JY�u��!��*j�-��cA�"0"�X��52c4D\��Cf�L����z�������(*��n�wE%�ۇzNc�z�i)���h̬�uv�_0Ħ�*���֫�cB���.N�!���wp�:S[�mn@��mT=�ln�}����q��3)�=ܶ3�����ۇ���q��v�gWK�Jv�����R��in������]�wR�8˹t�'v�֨c�{�X���c�OZ����=.d�;����=�j4Q$�Ь��yhdR��;���q�T���k0<�Y�6�k8pL��#!�g&����x�����`u���`Ե˻sgL.>�wz���a9�������9�{C�Ȳ��K�Z�:U�uL|��=��Q�����/
�v<d;7�xO 9iB�6�]wt�Cl��־[��Dq�WVmKzF`�te���)yL��a�.Cb �!��`}����A�)�_+7Yu�s4%���,���E�p,,��wv�>���ے�m��+���]=Rɧ)�I��V�c٬��ֺ��XF'5p2�r�2��Hg.k�֎�u3����R�76��d�k]W�XAZ��jH���9���;cu�o*S)N͘��x��3���o�pi�4`8����m����W��N3�3y�*�u����G�_u�$�,P��{���%#ã��K�{�(2��>݋c� l�%���R�b;���իEh�bvͶ�(�4.q�b	U,V9�0�od��u*�-T��v�>�\t����NخW�&��b���w���5n6�����;��<��NǷ�V�/9b��7j����p��V��u�2�`��\ܰ��Ow[��)f+�M`�[Q� ��e�[j1���l&��U��i��W3Zx#�CVw	׻�P#���-(-���E�^�X���;U�a���l�l��;�q/
�A�&�#v��J��V�
`m;Ю��}%���U`�9�w�J皊(�˼�6���l76k��Pgbt�[�cV��U-��w+�FeZЬ.�5�Pɨ����Y{Mr���=0`4�� ���ss�5�Yr@ٚȹ�0�LKQ���"�%�f�k{���CEa��^��um�U�Q�C�r�&�������u�:���	��<m�?u�.�R�G�D�vr�Y���G�������s��؎鱕�G��yEe�?t�;yI��&�N�H���ua�V^_p���\,�Vnp̾�Y�;�Ͱ��)��DLO^n��e氼�hC[$�ivW!*ov����L�Q��}�6Zorgb��%�kI����wV+��m^g.�f��6�MWKF��3���
K:ŋ��5�k'3a�ε�tO���^�����/�������^�|�ʹ$渼�y�-��ؐ�)�k2s����.��j��b�N��Z:�G��2��\%"/���ݼ���sp�y�\�g>�!�x��E�����#���J]�L��w�o�ۛb����)𺎛�-�9F�3�ᕅ�3���1��,1�0��ee�.��s-8�k��qy�N��6'O���;b���)k�Щ��ݣ�_h��e\ze��ǵ�8�(hüȂ�Ŏ��UdfcK6���2�&vKʃa�\<XՇs ��E(���6e��z7�t��ɢZ�`
繛�5�sj�p�����U�5�e] �i�+�:�k���J��YǼ�������]�+ga�hJ*�i��M�6��d��嬷��p;[(17������4�>��{2�g&b���q��-Lbbwe�`�M�4,�jŌ��]�Ppud��=۪��ٝ[&k��Z��f.�j���J`".����%.�nZ���`�v3�!�&��Gd��n%�/��C���tچ��,2���U�/7��j���v��������(���%�'rp�Bӌ�؁a
��ƙ�=�Z����:.�ef���OFT�{��I��"���)��,ra����β\��������������@-��Ҡ��-z��0n�WG1�t.�yxL��]�ol ��i��w��ۼ}f�*�5Zb��:��wV��7�������*��ޫ��o���=�O�3��`aɛ4M�M+ƈga�͈x;2�V�����A �,8z(fa�v)fNA�	sWW��7�gm�s��8fbt��g+�΍��#��T3�v����Dȹ��)�x�W���c*�mN��I�G@~���7�wueAy>:����V�.;3��J�xzm�Jv�j�x��j(��k2J�{�]��b��X���NA������0mvty(�m�,������}r�nv���4��;n -�Lp��Ȓ�]���[:�(�]���\�wٗ�[�Q+�ۂ�]�o�ἴ�������e��طO�j-�y��[3��;�Oh���,R!��委�n�9��u�6t=��ۖ�r���������D������I���sp�7pu���b�����]Q:�z��;���(�	�wgJ;�SOvݳmK�KbY}���ms�u�ou�^A�S�p��I���|ﵡDa�2�/�:���ܗ���������9�ʁ�MA0�P�#&\�9(�j��.�9�xo���n�m��2���t]��dfkҾʆS�K�V��i7yZ��kv�uq�a(�/s��>��6���|��쾭�%r��y��q�S�b�3:5�_D.Լ�����u��)��u���Ǟ���z'\���`��|�k�KO^��� 1�9L6��>�vj��+����.�w�l���ǆ_�C�S��7�X]i��1�.�7����|�ݶc�3R!�z��{ �.Q������d�#�[n����4��W���tH�V��vz��2l嫦��uWbA�JnD8�����㻺�<�^'/r��I�;-qetȴ���6�Vm��on�?e2G�,�ŵ�&w�m�}�z��W/��@�t�Qޭv��ހ��"ķ�{Np8ڍ�j_������*���`���f��@i�)���oy����ΐ��tbYg&�ʘ2�+f�`�hՄmE}v�Ԯ�7�ݻ�n;Xi"��2���nΝ}���'z�����S��n�d<q�E�7�-Μ����1��і�S0�|uU��R3u̲v��'ܮ�X��/��&.J��b����7����P[�ņ�q���7��U*[�)R�fn��P��Z��N��ʃ��Lo90�ڱxy���R�sz��m�=��X^�jt^��u:n�8��"虦���O^`�2��ZT\�r�T�ʺ��b2�J��n.1�\v�ZC�-�+*�R�}������;cR��S�I�eFo02(�RS��v�2&j��2\�X1�Keb��)�8̴�kΪ��������T����o��y�;��אWo.�7�*ѐ��^��ᒮ5����+�i]n��yP������D͹���Ϋ��m�Sf��V�C)��k8]7+iʼ%�i�D��nNrL��ML�����:3x^=��*���1e�����AY�d�ųk���Yt����ƪU�^�8/�nhq�<]�����
dn-���X�㸜����m�Nl��=�wfͷ�g#����j_p��$hV��ލ�n:t�
<�M�kV;|�`la���+�k1]�G384�n@I�;��j:��s-WZ��D���0��3ET�XK$sZF�4�̮���"���΁��]E_\�of"wGS�	'591�IX�]��3�1-��clov!�C�ջ�B���/7I��Z���^M��+JN��e�fĔx\nQ���i�uA&Ή`lV��U�z���fZ�n&�8�l�JrA��62�)st@Gs�D^*25Č����g���.ʩn�K����zGf�������)2�«��0����rge+$\6�hF��/*}s�O��0�l�ݜ8�`�y��s�ha���X�O$��9���gW*/1M�٤pGF]���C7"ޜ�ŵ��Q���Z �S[{q�f"����ᢶ�4�[x���3+�պ��-5hvK�Zv�koFQ&��邰u;ŒM��;u�Z(�ƛ�G$U�'u����w`0⚹n��`���Y���]��(wm������Q�d8��MBf_^��C0�o�n-gw/EM�Мz�1�2b�q'P����s1����24Bo]�T��c�x%N��sr�f�/{R��% �����a���9�Fն�Z�#�]�m=��r�w�FM���7I�iZ�`�Vh�$�w���厍��^�aJ��uf�[�O^ţ�#�IE7l,���M[�Jg1}����B
������]6��%^��� �:��v�.�Ô��7g4"�Q|���7V�|F�M�r�']�<i�	�A��:���u�䭈$[��Q���d�ɱ��z=Ba�(ň��rt�E1���r���Pi֣[�Wc�䦩�2OQ3R}+_db�l7����`v ���Cq�I��<������I�4�/]��C�����?an�V�=F�p�[p�b�*$��t�~�u_jQ�t�i/�͒e�cTZqbr�Smc��ĭf�	��.6��i�&�A�{�7��p���G׎������1�Ý˶�>��bx�p���
�+;�{�뾱;���x�U�y�HᢸUѸi�sU��Au��s.mu:�0n�{�N�r���d��vtA�s]�,��V��
�Տ��Mf^�mT�h�m���"2���3O	6��
��� .����<�c
'uv�6Iu�+jLݍ\݂n��8�&���W&i,��:���4k�y%�ܠ��}:�Li�X�].��R剚���+1�ߜk���u^C��j�̱���+�Y��:���<�U�2��u�7��S\�ԛ�\.^��|-btr�U�)u�ԡ4��ݸ�a���ƜڝR\�[��W8��7z��Bt�Q��nJ��
K��a/���"TT�ܣ�'m9�G�?ܽ�|(�
կ�w}ͬ��	��4���}�]�u�7��Y�mܘ��Zkw*��rb6-�U!Y7�֬��8؀|����Dl;8U�
�ʚ��X���`�����İa�1�]};�׶Udv1��cV:�m�0[/�.6s�=�O�p�t�U��4���$��v��¯	U��Kܚ�V�b��8�͙HP�+�oT�դ��r�j�Up�>'���6s�d�ܽ�Ĭd�+[�?K���E���z��"jU�rb��u�g�Cz�pX�\�ڬ�ogh�F�a��R�o;Vh��R�76��wK7hOe��䤘�{���(��*�FCa�<C& c�,�;�˸�������XQ�ۭU���Ө�V#Atu}W�YW�V+*`в�yXjy�W�T�S��qTMmw,7��;�-Uo��v>įr]��!��PZ��	C;W���w���eI�𽮤ދI��u�J]�YICt��4��s�_]�1+a�lKԄNΧPH���%^���wzE{�L�N����+�������[�,m1A��R�8�7�h˄�G]n辉Ʈ�b�Tp��H9���|�X���K�+%��!<ڴ89C��[��X(LdBc�75X���o6R�[E��Y��c8����^<�Մ�ܳmᝈngT$}�b*�#��aB�ַ:��$�t�ά�r&7,�q�7g_ܷ*t�������S���:+6\^�z'��!�N���/�Ɖ1':�E�� +��0��͚%f��غ�F�m�夥��e���-+m,��Nb�����^m.���bKj:��w�w�^B!,��V')q�lqwf��6��-#���p����T�i֮�#���z��p�qβ�)��z�ݷ���t^�Ҝ�ݒ9�u��+*e����{':9�JM!��=}wVizk� ��r����l�/�5��+#r}�r�u�S[u
.uYX6,N�����UkG\$��[r���Z��;gY�.t����L�wmU����=i�����/�db��/7E��&&u�\(d8�r��3rr�c�����{N�d�Ō�6ꚽ���9OB�cSwZ{�/7�/�I#c �g8_����_0.�8}_���;��>O!ݥ�/����UUUUUUUUUUUUUU UUUUUUUUUUUUUUUUUUUUUUUUUUUUUU UUUUUUUUUUUUUUUUUUUUUUUUUUUUUU UUUUUUUUUUUUUUeF$ۣ@���k��2^v�ct���\Z�����b�--��e�� B:�R�i�ZEk�7&�[��bmv�10��-�.�dl3�#bɁ�B�XBg7l����W&�4񻗧	�x����"�yA�X��I+�\��K�r��l5Wwn�CY{g�	7���$�ju��xM��g��J�B������Y�w:�Y-��s�Z�BX�J���Ansۃf�v.ݖ^75�A"�m�RW#�A��H�(��%e��H����WJ\n��
Nj.wD�͎�v��DƬ�l�SR\����M*�/2͜4�#y��u�ꮩ�raW��5����%ٚ`��q4v%,ڶ�I�O8z�r`����v�e%��gF���H����/]vҊ��p�g���V�-�Q��w�2���q��zn Ll�dtpF-A�r������ҽ�ώ2;`����xN�؀�ØWWQ�c�`�r��Uc\^��ؔjF%&���d�y��I�ۭ�9�:N�uĶ�8Ǘ�G
7WGk�޹�l��!e��W�K��ь��Ńqnh�Buq�s��9�6�c[��8�2���Lq���r��0��A�(���3D�].na5�鮛\�����\1�XhN8�з+���qڻI��mH:�Ě�'Ub�6�������H3`��:����*nWXY�������uNx8�b6�����r�<m�v�3J�L�<!�ݘ
�p)��bN�n8�IV�F&0E4�K�Z�2����̓Z�ꘖ8u1����A�ܣ�����S�|;���k�f�
�3�̱�.��0�A��BF�\�WX4�&e�bT$���K���/���:h��l��(�1PV��#�E��J&�vv�pP�v�l)S��o!���X2:�����Uj�헙�i��IF0Sד��:/nŌ�-�gM���� 㗗SջoY�뵪[e�1b
˝]�����n^*�tjŉ���n�5��d0-�bSKcҗzv{]���Z8�َ�7��9�A�gtb'\x�x7h�!��p�pl�Ƶs�dH%�dX��6���5ѧ��۵�T<�Wm�������i	�5���Ǝ����6����Wkٕ�K̎�۪[���`8�.O!u�k���z��%�(�(m�s�K�PMo�^�dˎ��ź����i�]�O=����Y�U����\Bm5��zw.Sk�$��un-���b\K�Iqx"U��&�B�b� �f3evcm��	��J�S0�����n�7�MvwI����Uū�\�M[��eE������r#�a0];�m��}.o<�\��\:�b䅰��2���v�c\�9,.In�.Q�v�N1��Ӆ̼-�������bư]��`i��a��dՎ��%���+nxxA��n�C�C�힬�Nm$�l�"b�:�7Xؤh�-'dw@��6]�v61�8���d�v�s�.����^���Ӂ�ⶃkV�"rf�^z8v���;e�v�
v��p�����6),x	�`Ԛ�\��&I\=i�����0f��餱�L�!N�:�R�5%!m�=v�i��Ĕ�uW��.�Ŋ�6��s�F#��#֖��(u���k��v�أ�<��f��&�J�I��T�s�ڀ�(Jf�mu�m�F��v�ֶh��c;���r���eC�� �n�����JD	�e7�T��xStlp��#�L��vx;sv�,��Cb��R$!-%�5ь�m���uc,�@ᮖ:�J�qq��osڇrBu��-�۬G-��v�i��Ř��'��ZGe��l��<(ۀ�����=������9�������;��7��0�z9�ݗ<���Qp4�dJ��JV��h�XM��\��e��Ս�;*[ �Ir�^�u��n9�5����]C���/m�:㳎X�͖
��]��G�E��a�U�¬q�띒��i������Zp��U�'G%	<��N�˻pm����ܶK�$�dj�3*�����X��&��3�m����v��F�.5;\4�/Uq�Qlns�	��%��ͷp:���Id-=��|c<�j�tFSiXs�M�.[�����íן[�����ˇ;l̯F��ڽ�[�M˖����Z�kRg
���:VC2ݘ���C�9�.���OdR{�m�y�Jr�L���;o0]�rb�`�,{Cq�[��z��92z=!V�nG�ܱ�P�2i�s0�eJv�Z�wh��)���^��p���C#�1:;�ү�6�YK�J���� ���j��hMH�Ѷ�\��둩mfl
N��m� Z�\�C��J�v�3� ��j�;<7cx�b��0޳9�1{ �٤���f�YQi��<<�ћ�us�nϡ�ƞLG�܈��oR]����SGER�U�[��kŉ �Av袸���;lV�J�M;r�\��6!ݝ��ۉ�9�L�8�R�Q�5�"��c�V4�l],�f5%�$��̺������E���1"8�͵y�.���m�iz�����Z�dĥ����x �
ҖZ�%u��e���]����ܱ��lf��"�V\�%.��z C��ئ�����&�aI�)b1�˭��P�4aG	tu&�U�v���,[�e���TN��˝+]Ό���WDX�m���f�㋛e�Sբ�I3��B9T���F̓�jJ1sb��q.���kr��^%�(V H,m�2�y�0��$���l�F�]H=����$�v`��%����4�K��H�m��6��i�2V�3�H+����i�Si�
�˨��-��+�@ȅ�m5&��T�R�'
�V3�>���s�p0ah��=�ɰq��)ؕ������h���C�%v��v=h7�vW
��	e2�pg��s��]U�ى]F�h�c�٘XR1a�Ѷ��e���4ҹքn�Bd�yMZڼ�'i�I�#�.�5�f����ۙlS[����ɷ%��kZ��Cs����#+ǞՐ��og���اGg�����U��b�lJ�K�m�yx汷b�!��g���ib�ѳZ��n�[*Ld���r깳lq���l��6�ܽB �\E����3D�L=:�9��y�\q�^�Kn���n�K�]�����E���a��M6�GTu&Aˌџ�7[[#��JY�u�T#�\�f��&�e�.5�5�Qɠ�3���M5.z�7�B]vb�[��9�E�4l�3e��[ �k3����m���#%�.D�-�0��}vr[�;j��l�������l��<튶wO=�Gm�9���Nn@�6�7���9i%�f;ZSItqeYM3��oW]C��a��k&�z]��v뇷DpEN9�30�e:�=�YbY�1)���\�J��lش+W��vvS9�T��2�l�d��*z}��;���������p�[<��M�C\]��bJUl-U�	�`8�����6�q�:Ƅ[E�,ڍ�����6�Kn�R9��+�]]�a��h@P���6����&k/d�Y��p�u�c՞W�+sωu�)Y�t�q�}z��vFn��KK���,h�R��]�x�������v�a��\�D������)�6@��6�q����l�;o6<����̳��pG�W�����9��[{lK�3bw	o�rڬ�z̒,3��6�h�R0�Բ���1m,�Mc��ʦ���E����5�ց��9h��A��YXl�LfY�u�3٬aV%Gq�2i=���n*b3�F���������^��nVĤ*�K��Qq��tu�/7Z7,O�s���8�#h�ܽ�oXwu��ltL�h�R�V;8ٸ�M�),6�2霑Һ�fZ�h��k�����m�GGb,3�����/. ��m�0�����gk�ɮ+۝����03�M\��E�2ȠY�ۑ��D�=.�ZKny���F3-��5ȕ5�s�i�q)�+���d-aݟ;�c��=��+Xp@C0�;!�w.�.6�2+t�ɸ؀�Zن�	��r�14��,[)W-�ЪݶЈ�m���ێ�%�㶧a�K��ڍB$KS],`�$���\Fٕ��.�Pe�vP��e4��:Ļad�zg8y,.�J9';<�E��ykK���!���n%Q�����Ja"�!�Yl[-��û��܋�8��;t����c7Rh�6\�j�6�af^��#��^c͸�3���E�-�+�(�mk+� �� ��������������1�cK�����-�����؎p��X!'L����!aw3��C��Ap��
���J����d�*�!��UƐ�:��w�_1?wiDON��J�;*�\���EU=��q�r����aA*������5�w�RK��F�PmvUA�y���\���4��r��"�f9ܝ��/9��-N�s����ȗ�N:�E��z���/]�(�#ԛ�$��U�?HzApr��*�"��;�)���@S)Ը\������I\O�z�2eTd$k\�*�I��E�Nk)=FU��B|aL�Le �PW)�#�<��eUPSdM�˄vW&Y$�C֚�q3���ʋ�H�Ӕ2���J��(L�(���ޙ�G�hky�]"�ȥ�D���H6����d���k��1�b�UUUUU UUUUU UU��0Y��X�g�rn�=m�ɱ�#��{㏸^����KP(�÷3Mtق�';XL�l�k1��y6zZ�T���f��k�]��6&̨�92����f6�Xˈx�ΓՒC���l�\1U��h��Ѻ���/j��Љ烁ꍹƥOp�ڨ�m)�kb�ՙ�p����ͱr�Y�sd�bmu`\`#�qtq3�����s�m)L���Y�%��4qh��:{p�+���'Z����eA����e��n�xn�;��h�p�Y=cd똤ewZ�]�C�Y8,mq,cfц�`F�s�e�SO�W\څuݧΦ����*��$zSF^9T�]ۣ�v.ŻX��kp�1�)3A���T�&���Ou��:��X�F���(c�4p�X��!HiI�4��9{��r�O��hy�]��j�Drz6y��m!ŤV\��]�$tl]f��g55416�HS.
�
Yy��C����a�utt���Ě`�0�RT�*bvC���r���!�Z%�ΐ����sq�6��wȲ}өܘ��=��&�uر��]��d8���n���;[W`"FX�6�����dk��t�EK�ؤ�zM�wf�i-
ZM�#�H��`f.s!Ō�=������tbzNx8i;�Lhn�ݹ��<qv�����zqHCC�F���$�ƀ��(C+���a8���`����B>:\&�;n�V�^�{�n��h�Y;n��)N�E�r�Og�q]l��.ڽM`�f��G�n�:�qҎ޲�&�8vt���Dݓ=]&�����&\�ƹϷX<
�6]��Y���H�t\��5��etZ2��K�PU}�ӻ�z�  ln�,��Z@"��#�1=O5�J�u���/)L"�^z��#��ye��)��מ&=MuQz�H8���P�=>|P�Ms�q㫂zB�s<^��.��(��M����q<\�M
��*$�E0�#tp�u�5�3W/\
�4�<=�-���}u�����JXB`,ؘ.��<��׿��4�$��_���/�mm#۔&�I �	_DHK�7ù�^F�T�]M���gг4o��-$���~H�7{<��J걶��0�{�9D�I9<�$/a6(�<���A	u �%Ʉ"$�`zr}D�@٩�� tX+=��2�@�$Oo9�Z(���J�t@�3/�ϋ~��"/v�sM ���pTQ9{3I$�]��9�ƍl)�$u֘�^߉� � ��)p�7�=ۮB�=����W��q�����Rd�I �9��N
���0fbIv�"tܲ��E�����Zڝn��2庨������,Bm%�vJp�h�:y:dTI����;/a�xNWs �1z� 'g$�My�ڣj�@�d>��!5D�;l�W�(�����q��R�t��E��K^:��ֱc5{�4eK�:J�q<K����$ڼ	o:�7�>k�[ݔ& �:��V�I�&i$���TI/���B6�m�P��*�Ǿ�i$d���d�)+�ʱh�m��==8�D�{�4�	%��tm	ځ�`�� ��#ݛ"��z�[�m|I����d��5�v�BHK_9�~���Z�K:D֜	$���$�a���bT�>�3<�I$q� ���=3!�4�Jw&h$��Z�.��K�9��\q�0n���2%IR�A�e�m�İ�[�j@�fd��0!G�9�e2+��<<1-�A]�]~$9��$�D�� BG�ژ1������ ��ܓ�M}�)qJ�P�&�PBD^���m�`{�\��Ow.�%�Z��a,�oDc��oL�S�~�Wj��D���܌BM;ݪ��Hȫz�Aq�Q;JagfI�q�KC5�S��h�N�N،�l���	%-Xbt�U��h��ۮ{fh��f"&��P�gDd���A_<�&�F�����'��*��}b�H�D�tT�Y/�e%����I%��9�	 I{u'��=���X����+Ԭ�� դw�n�$�'��*�Ȕ�t�ZKsn��D���7h��\��������Yn���a��nFWgGW�:�us��y0A�v��EQH],�>F�R)]�_�{�-$�H��4M���4:��\ﰹ���{2J� �j����H] n�
�R�!�O�I4��{޻��3��&�4H��N|I��D�&I&�I���s�y':^�K��Z���IA(�d�I�&�$�;�!M��sǡ$�9�怕D��sؓ�K|�mUڥ@�Q2s�~���ŎeS�	 =���V�D��$$�}����<��]*ў�Y.��*H>��{�{a�x82l-�����d7�^m��(q27�S�4��za̤���@ ɋ�	���"���b�H�HމI�&g��W_�b�a�3��G#�!$�N{R�$�=�Z�gGwupܸ����$�)H��**e��\��tĎhZC2ʕ��nV
0'�>���Ų"H5��٫I$Knj�	 ���vLhܕ�o�W�0 =��Y�49����(�$�Cz�R�ޏ,�N$��Rd�I�{d��@�c��\�BwnrB�t�VR�	rA���n��I�T��2t��d��H��I�����%d�^V��D�JH��$}�eF����ͦɢI'w�$��D�';ڮc˧O�D/�{�tIo���]�T
!�nI	$�H�v��ev��@�� 3ݲBI���P�����ˬ�8Ć8.V��9�j�YIm���KS�@]�oQ۽�+���aL�&�du"�QM�6�ݶ�I*�d�5�J���Ԩ�9Ȝq�nn�c"��8���P�^�.!
�k٠8qOlAH޲9��`+���{�=���+F���Evo��C}�熮�G��l�vF��jm�3l���-��ұ��#����B�"Vw.w 
����[un͇8�X3"ŭB��ۡ�r����tʛ ˰es�2�pM-�y�e���m�K�$MItqEelhmgM�ʌ7�~�����X�I#߉��3�؟I!f󛴘y7�T�V���U�f�I#��ؔi.��m$*�
Q#��N�R��e���W�V�) ^I^�&�I.�sv�+:=T���
�s$��,( 9����(��BM3}�� f���J�ɩ�H$�Y���$��o9��?g�rB���+���$M��m�"u�9�`-��|ߜ��I5G{�HI)x%��!��Q]cDe�97�b�o�4��D�K ��8I4H?&�~ͣ����v��I�����I,������w���fu�)X�Wv����6+�Vd{8�!6�!v��;��4n@�(����Պ�\�)W-חD�Ov�դ�'/�I|�[����&�����$ �ojbS��b�(QI#%5�6M�d��\d����k/��1�v��f��Ā��.�v��_ws�����I���ޓ�3ﲦk�њ����<oВMOwj��$�''L�K�9e<Us��u	�{D�A�H�f�ZI"]��A$�vf,��}��N��k�$��Y}3I!j�@�����-��Sw��޵� ��O�I �^��	 ���T�l'y9D��'��)	���$.��
��JX�XɪH�����������Q��
'���	;9'�$���s�i�e��,�3}�寣X+j*�w$=��p��su�v�[�1�@�PV��~ܯ"��D�� x��$%�MxR%$�����J�d����=Ы��*��5D�rL��J���Z��nI	�$rNv�nvj��tS	 �	u��	$���v���1-R����	���߁W�I#'č}4"PJ�X��H$�BPg-Ύ���N��� �?P�S�L<	&�j�0g��b	��VƎ�1��ī+wu,�!뽘�	$�K��I�=��me�o��u$*�
�U���&�A�Iy"r�j�$����%�-���w���y�����<Y�h�����(��$ '�g�-�Î��'��$�7���G���!Λx�{���������̥n�3lU����1;9�VRg4�],��J��
��J_���:dWsuv�Ir�qW�"8�c�RI鹝�$o�\��̤<��H������[��Sԟ����@?Nݒh�}}�4J%�qcHӝ�����R�U@�d>��* ��d�	 _�N�QUE�3a$K���Z)$�wd]��"X��U�RH�TH��b��pyD��q��p��ܢOĒs<�2���F�����Zb(�:���Jv�l�x{J�F{�N�y�|����y����DuL�+�p��]n^������PBgT�&"H6N����$�%㚦a�[�̗+��xI�ٹ$$}{�rI5�9�I�w���T�ά�Wj�K�n�q=��b�ެ�w�>�x���atsk����g~�� D.�LO���|-�i�RI�$ɝhb�%RI� �H��mϪX��*�*
�)r��?�4I�\<ff��;`S��7�BI$�����$�g�d�t{�ﭶ%=��=}�w�R��H������ȡ�I o�:d�h�����fGMr��H��7\]���K9���O���	Z��L�}ے�� �Kl$����&�Iy"_9�I���y
��[mֽ$��"�]EzG��I"�7� �L�k��>�}�Xs�I�n.�%y,�3I/$��eش��^׎�7���<�]�\wyT: �S�R�?^S������me�;�An�-���gAԶ�0L����^��-���_5~}UWTY�s�<XFb\oKC�<y��w%�^��m�ng#{d:E�^<�l��F*Eŕ��) B�rYe���.��}X�Wa��{qm�4=k�9�A�\�eR<�m�-���q.�ٓ�|�K����8��;s���8N������6U�f%F��s�����������-��p�휲��Y��L�\�E�jV`(��G�M�M������G��1A�-W�bl��&�$J��v��y��Zs�hwֶ)˕P�j�D���B��#hZ�XSΝ����&�.��6�@$uk���Anv]�(%v˙�yY-!��R�.�]�,_,�H��! �-҈��2;�-$-k���Gs���^/���&��pJ&fzBb�D�g��G�M4��$�=��� 9}�s����,�r������E*)QD�>��bQ$�;�Cg�tm�H�El�I>�d`J$���ܪ�^s�D����ظ��Rfౌ�f�ll�Hڷ�#*m]�˫`4�����G�*��3���+�D��li,��i:A�	�t�⛵�=1I$��c�BM%뺺#�RhP��3�l�8�}Mf�]m����5�.�a���E�[OTY�;�|û�!�]|���{��fn@B��Գ�%88̱����z�%����%ydw8�h����f��0�\�@�\%L��\_�W;�H�I��sh$Mi��;�e��0M�[ے}4I9}��9�*TڣJ�'s�*W�/�8an"^Jf��Z^I�F�$�It71��=����eB%��HĬ��Z��&�J����@ =��}G����l�Z��	4Hݿi`BR�n`���}�_�&&"I�$)0T�+��hxd�v���nN��cc��G1�~y�߹Z�d)Ky>yw�D�%�9�Z	 ����0��>}R�5Q���P��$���>�;ub��MI[�O�D�Dɪ̟n�f��$ߒMεv�(���4Y���<�=Ǚ�%��6�!v�;���]���HH�7�S̒J������<>�����?��X���Y��M���j�.��\zә*EI_�ݙ36�̻UZ4e�}i���zՄN�]��¯��s3D3��c��TV4KPt'b�גgQ< �q�ĭ�2��'ۄ_	o�Dt�
�#k2h����+�\��O��1����$�4`3A{ۃ^�S���ck���ԧ5�\�+�=��5n���Ǜ�oOVM�hd�����
5y7Q1X���j$�;ak[y��BS��N�Ǔ�
���z���`�vhfv�>�S��vK��^m��!�LȽn���Lw��\�P��Z��w��çԁ�[���3[b�oX�*�8����VLh.ӛ�2\,��N�̽vy�3on����ɏ<!�Ͱ�v0 �a�bL�i��Ff�@�6Ϋzn���ae���\�)AC5+pS
���^�ŉ�!c���*<2�U֎ٽ�5�ĕ�z��$��Sk(f�w�+���5���՗��K�=�B�t�T�2��{}��#����;�{׽H��`�e^P�W�;/BǕ���� �j`�P7�^@Q ��)�/��H��-a2N��j��B�д���XT�C>��8��x�u�t�e��4��W��.����r��rÑ�+(�#�����dwY�3Or�Ҙw�#}�R��ne�:�s�J�����1��YR�;w�$@���P�p�� �?' ����J�W(��t�˧`QE}��dE��O$��I��yDȜ� ��QUGu`S�O*H(���#R�p�g(��$Dt�(NSs�};��72����=3���G�g��.�Ą��.�7'&�u��\���p��epN��&�.S(�Wiĩ"��:	Y���I��_DU77G ��M$���U��Eʠ�#��t"�Q3@ҙMU��˅�r]MBP������1%B���9�%�VU�F��M�q5V�۹��5yp��EzQ+˻B�E�C��'�r'�5|���R��*�I4壻B)�BDأR*��=�ݝ淝�H/�O�Z($����4-J� ���Q>��W;��G]΢I��XD�Z�(~�&?�բ�r�^Y�h�Z��a������ ��LD�F�_MJA$��*š�#Ѷ/�H8��.��'��$}��>�yf;��`��@ٴ��n�	�Hѝ�/-lrX�\�ѕ:�&�-�T��<�љ��*f,����v&�Iy#˜���	/nv]�J,Ow+�Q�_��+�ߢŢ�^^��l�U�H�j�TQ0~�a4H05��*���o�my"PY�	���c`BkyS�nWy8v-���H�hZJ�'OD�D��c�P�M��Fj�ro1.��|�jI$G�b�I�쫴����<�#v�ω�^{ K%��B	j�`�	����$�K6y��Mt�SG���l�F��%�:Q���]���#�M�/�8l聓]�S��*�X�6�#{�]���yz�~P�W�@~R��H�&&"}q~U_�߭$�n?;����<F��3@I,��(�bt�$����,��/�~�ɼ��7+�F^2̶�luH��-�&"Rf�J*����ȟDHBTL����+sR��^K��Q�$JΞj�)Ӥ:��y�<��Z�X��=ݒBk&|���6�$�	�2_�>�h����
f8���쟨�D��:&�I�<���B���.k텓�^g�߱�W�#�A+F�Z����c J'��آo�,����V��H/���D�r�~۟C%�U�A hZJ�����\���1�x%�=��J	.����I�~�E�F����\R���G�l�A|��i2�$�D����Б%�sBj�_l�ut� %7�j�뻒@��wuw �威��P���^�ݧxVa�ꕵ��=���r��0ˬ�%�c��ulj�[0�c�#��ñ*`Is�^_����?���:I���������jeJ^L$KuЖ;�v��f�m��͊���e��l�4R7�t
��Nލ�gv�l�yܸ�+������+�8��������s&�V.�Tn�����mhl1,����g����n\j�s2�e����E\��Q�Ý�������t]2��mƘ.Sj�4%�lN����;�,t�t71Bf������)�ΰ�b�I��G���~�/�������i�M>w6�%,�r�)�\*E�)g7$`BM�{m�X�� *�Q��(�n��D����������א��Z��Q6��Y��RD���q3-xժ�^����czg���]�A+��$����C$�M����&�N�I$�����s�QtI��{t�wj�L�}ۓCs��^B�&�E9)@O_j�D�Gg���xP���pLq&����&�E�e�H��(�>���$	���p�cړ�O_�\�h�}}��$���{d�T�M�x�҉*��D&éj�������Е�i�Ick���X*�|�����I�$䷣6�גA"�sR�I#���(��*j�U#i��U8��d�Q�x :�%v��~�*�w�����y����t�ol�`�\�J
L�v��.����:�m�l�=Љ��P��c��)���x9��H5ꣵ��N-u��#.��-$��	f��I�]�;�Z)(W��7TVGl�ک�G�H +W�D��S$��>��� e�5�bc���	Ok��$�Ks�ݤ2����� ���(�/��/E���$���RI$�몴�IygO51�\���?�ֹ�hj�ժ�v�$�Kz5�_�tƔ�ԒW�3I$�׮��%�<�W�:=ծ
���������WcM����#)�u�8!.*�-�b�����PT���6��t�����#�d� L��P�@?g/i�A��eъ�D��2MQ$���B<h��!�(8Oz�\$����2�) �'L�@�n�	%%�<�~K�o�
�nfs�&��^�I]����t�	$��~���H�V�rE�N�^���	k��H�)Ղ#9��g�^�Vz��Py��e���2qk��W�0c� �v����*r���}w�?y$�Y��Ţ�K��ՋHb�Ҫ��j�
��(�&�ss���.�?I}�؄��5�]�J�@=�2��wd*0��D���HMcϕ�$.��	U�݁�^H��5KF��oQ��	!�n��D���b�Ey$�vL�IvOsq�����,Q(#t�ڻR�Sv�����q� I���9��yF��߿~��FWo_f�ߞ�� {��. �sؓ�����u��|���A$�r��P�q;uеF��� 7� �v�~�� ����F�I��Ȼ	$�Y�2M ���ǔw��\�%R�� �,J���\�6*�$��dגId�u�eI��':�"E����I=�?�5
$�ԒWk�p�N�s����}􄟉Gg[ N�$$��w��M;,!0k�J!!WXk�6���V�"��pN�R�t�=;H^�S.���nh�$(s�L@C�R$Zױb�j��"	
$f&.�#v�I4�5�7�v��ey$:qd�h��H ��d�bV�r���2�	X��[�������қ��Mj��ݗ\�X�#*(�����@����,͖�$�7؛%$���ߒn�U��Jqܨ�	�Āt�
F�j�"D�}���TM3˹"����UZ"�I$[�3A$T{ےB '�r�����q�K����B���	�$�TL�㐀h��L'���"oj�^I%��4��H-��!%�+��6:��B��D�םQc���I"w�kԐIy%��˻I�\��|e{�%�H�&I��
�$���\/�� �Nm�%�����}�ʖ&�M�tI$���F ��/a����ᛦtF'��F恺#W,&��:�Le�^1���a<\ݼ�͓�v�-��Sa��Wf�z��g�7ى$�IV)b�lÈPH2͑��g`z[w]p�޺6�+z����w���#=�^�����آ 6�p�;����pm�]6�i��z��F���\3hDf��A(L�yڸf��w$\ke�ѷ%e6�q��x�`-.f9�˴�J�g��.���M<��r:�ka�Q��cFŨ����酕��9��-��K�X���6̺�0R�DZ�#�5e"f*G����� +W�_�D���؟JY�خ���]��;d�V�ط1A$�O{#|��R�T	6� �2��+iTi�V��NnR�K�>yUi ��Ξ�v�%���)�5�b7���J~�v��Z�j�!���	�_ap�H�L*[�K��D����!�M���2[��]ThZJ����\W'᪗�r�4JS͈H�˰�I����E��כ�_dtI/2IP���t�R7hP��}�Ο\$�F���c���a�weyL�~)yk��v��I,�s.I�3ɥJ��*��b�٭�t��/@�	�p|��Uˤ�d���A�߉�_�$U���_��	��N��Ua"N.sYV��g��o@U����O�vP���r6hQ��Bю%���Zo�*�O��B��#�,E���9�	�rjޞ`_�.��̻�{q[�n4�25بn��I��3�x{��9O�WZI���"ɰ�	g�f��	c���&9�Z[Y遲&"A$ڸ!0Α@ }�I�w�ע���wd|�	��eϪj�$� ��˴n�V�R$H}��|�b�N�I�~�J I=�2M;ۭ�z��>����L��r�?H�X���д��H�D�$�&{uϡ�VsP:��I�y�i/$���0M��n��q��(<���}�Ҳ���ebݙR��r�r�	m�z���6m��$!x� �&"$����ι��%��$�K���vz��z��tX��5G�uXH5�+�R_D�7h����9Y9";��j��d��]�	�$w9�a-���׍������-���D�'ݺ�П�$�����i�P�-x� xǎGn���'�wn�V�����d��KS��R���I�o�eߜ����5�e�_�x�{��F^nF�O�8�0 �~ǵL�Z@m[�g��{�Ȫ<�� ��l��$�v�(�H���`���n@&��rN�4��I(�V�$>��!4I'��b�ڙ���2��}d�I�L�H$[�Wh�$�Gs��:Of����Y� *�EZ�3���k�=����ҙ�0��%�*>�����&[�?9#�s&��B8�j�$�K�;�I�[v�	o�3I�滣aL�u@(F��� ID��t��Ҩ�_�1a�kY �q�w~H����a+��n�K
�2M$��+-R_4�~�D��lP 9TY�z.'sfh$��7�شRH,��U	�����Ѣ�����D��*����Iպ�a"S��i/$�G9��^�y����^t��{��ǣS�'�?�9a�u�E�V�z�>����Vƃn��mvY:���w���}V+�>�9Ap�UUr+�AL}|}��vFįL�]yR�T	6�	�0��( %��ԧ�}�Щ��i�ݤ�-v��Ey%��`��q �5����nT}2�I�>�Y�Mr��k����0�a4�[vb8�n[�����B�J�T����rJ� 8��($����d���.F?)�������D�;�P�q�GY hZJ�|��A.h��v5�n�ZA"W�8���4r���uD��q��5�1�R8�#��D�n�K�f�i��$�Jj�V�ˋz�׋ ǯݷ*9~�l�'����QI|Ԣߺv��/Z�?�����H�ڬ ����ګ{dr�zD�.�z؟x�r�4h�(!h�(�g+�=ۭ��g�պ��v�$ɹ�	 �[�>��(|I���0��5HF�gM=Ux�9{�:rv�:嵽���ɓP��f��x�]���.'�EI;��؀+��qJ���u�y󫄜�V�޵�뵂�Ӎ����חg�S�:�s����FnK�闝63ss3G^��l������}��ec���Y�6�)��e'����B�߬=:t�C1�ܚBQx��	+lZ�ԓg��y��������1x��C`��rM&sQD��9,&Iy�b�M���h<�6���͌6��\��,�ѝn�fR�=���u�.���(n�Z7^6"��6�4g�90�;�(B�SE��o"'d��ռ� ��ZN��Fmtݑ+�v精�36���f<�b	;C_G5�ǜ�o���s.R����{m�?�ܮ�n�4�m�V�ܠ;2&n�Ub���f�MRMN�ܓ��� �  	U�v����4��뻗�z��B�{v�P�J���p];�}7W<�YH4��6$��E�ͣ�PyΫ�`J�kC�	=Yj�sl���=g�`5W�\�w�#y�[����/�*N�M���ͻX �]��Nuۢ����T��ɋ�`&�J��芬��	��'A.�(�jӹ�c싚F�73M`Z͙.hR���+�uy�Cok�ջ���������;O{T�+���+͇����!�FU��n�~B�o���'V�ʢH��6uH���S�<��%D^H�>�q��N��Nns)m=GT(��t�[Nj���S9t��瓆0�1#F��Bwqq�P�3K�C�ڝ:���11eI�TN�An����ΜI�t�a�� ' r�(G4�7sq��-�B*���IrK���s����"���A�e^�QQU�ޝ��U0��s1�\�#���U��)!�P�G!�eEIGP9��B|H�E���o��\DY�w:Y!��.I)D�r,&Y�q3M��$ʧ'3��x�#K��N$��N����s�9�I�GrM��H/&�sE_:t����⪪����������������\� F�X�*�7�fY,�s�m�����ɺ3��>�G�s
��7n.-&\�l�����ej%�6�Ѭl#/n���ݜt��+�jw�&xN:�v��p��ə�^%��읹Kv7�4ID�B�� b-�n�9�<��2�[2�HL�\mЖ��pM�督�m�vS6���xi�����L2�:Yx;l���]�#í �p���5�)�l�*Ae���X�Q�f�v��nLX�8��v����19d�{Jd����va6�\]�v�ޕ�7���8圮�E�L�EŔ�uF�1!�p�!�z�K3-��È^*�ivc
�R
�[��t��K����ik6#��!��������]�Y�٤ݖ���YH����WB�ۮ"�#˃��m�W���魞(�wk&��3�%�JRT1f̑"وM�˵t�b��h��4u\�5���<���L��^�t�������k�����9���uaY���.�����#�B%K�1'��ۛ]16qVڈ$p1+R�P��
�i��Z�k�0��F��7.�wi�ն��[����&�SvZm��ɇ�j<`b[���4cG�7k�ٽ)�ԔX�,���&W\���ی�-�Weӳ�-�,Ƃ«i�0s�K�5�u-vk���.G��b:���	���u��7��M53s���-�vI�|�)R��a4;�8�כ�67�ˌ�n�Ճ3Z���&���F���y�G-���xe��.Wa��&�ƷK���s��R�'6^6�M�mfWd�1�K������!TCa��YB��Zɸs�l����6�s�6a7�ƤM[u��0�Ԯ,ˬ1�Z���]�mfs���c�4X��1�F
����;��>�UV��´�Z�/d\�8���hz�{���9��s��zIy5����fNL�>�:S�;�]sn�9Ժ���Dm_���}��{cg[�)��*�ڄĬkWj�<�9�o!���]8��G#�z�u]b,�܋\b<qc��簩�8��׏8EAk����ٓl�5����5�Jh��[+Ll=[q�kk�����b���v8�3%l2*�W�9cV�`H
�n�H/�����HڠI�p:��t�+@$�GW9�+�%K��UiIu�-M��x�y��|z�j�D�o����H$��̒N����)�{:n=��Iƹ�i$g;�h��lh3���h��Ǿ֗^�%F�� h$���t�'� f{\� ��k���	�s�-�s^	 �9��ȓ�Cd�Dτ�D�����{��]�$���4I$�=�$��H��ێ2��fX #m^aG�ub���B�	{��I4N�v�;$pP��n���؛���#��Q6Idw8�Z9q�#r�u�M���2-F�؊=���,.#Bi��K]�tJqRJ����Ͼ!����J�����5:D�H��*Hw�U���|�y��m"N����	�!ɟ]�*F�M�bQ0�$P���u'�.���"��B���*��=%]z�䫙��Z���Mm{���Ρ� ���N&����ųT,N��{���SɃ�D��ݒM���qb�I7tDuŃ����~oz+V	I$� H}��- �KS�~I${%D50M${9Ԅ$����	�z����FO���8��P�m��I$����^Iy$�� ��>�wW���d��{d��Ha��whP����)�I���u4w���iu�����%�ɢl$�G9�R3��T��pH!1�Mz!J��
#�����z�'v+�HH1l��u[���{��5��s�S���Iۖ*גA#���%v|���t�$�'��R�8g�]�4R)Z��0�M�:{��8¼���H$�Acܛ��I��`�J�у}�z��'^|��� �j��D��vZ	/$Z�4%��^��QP�oݶ���KP#�UܥX�̱�qg���]�׽�c���y]�k�������������=��s�I?��@�_�V����`��I�}{�	v.�v[H����ZI���0M�[�� 9�xD;:�����"��6M�-�>;D�I���2��t}�C�9H�s��$�Kz\�	$��n��NYn�9���p�&�*J�5b�/�"��&�F:X�*�j7F�e��kZϳ��%��P/��k���Y$���B%���%��;=�	��L 2���Y0#뺰.�nЦ���B~'����}�Mp-�p�I$�刀�4{ۑ�(�Z�=/�d_�Ő���vh�T��j�;�d�I'��Wiy"wg���wW;�$�^M�J��$�{rJ��ϕ�(Z �j� zG�t@���*�$�/�"$���r�$�y�N[�͘ݩ�Ŝ;6��bû5�;��}{w���9�%E.��wCg����Os�Ԯx�.��s8�B�=��}�}��K��Mؿ"Oz$���I @���� �߲8Ǣ�p���]�IY�r�$^Wۗb�^H��ɿZ�޷����]~z�]���B�X��5WF��دW:%��H"���TRB�g��B�M�=�w����ʱi$�AgvM�X�_��]a�͛E�����!-!^7@���$�G_lդ���1�𸎔I'����I#��)P�D˾��:d�Wyy��a&���n���,ݡQB�tbh�����|���+��n2� m~>�����s��Bp�r�`�_/����a>����H��T Gobr��D�9~�l�iI��0�g��Bk|���b��pJ�D��I$i��H�8nd�3�I�� �7��*I}���wV�c��<�q��ƛ�����$.�졜�8�XoK	�d	����`�n����{y&���Z1��w6i�<kp| ����UU�&4��i)��Vc2�koQ���KfNkE.m��v�yۮ���e�<J<`���]���j��9�A�����`KcVvQ@	f��WIV��f�.v��J`v�x�n<s�����X��U&y�:Ӯ��X6Ư&�{o���mlfs��:�ӝ��6�y���r����+�2� �ܢ\��I�V��P+����K��Hu�ktp�omaY��H�M�e"@�vd��@����\�	s��Y6�V�Au<���J	k�R�*6Mu��A$�O��I/-��S����$�Ϝݤ�K#���H�Kوl���W`ZBfH�(�0�$�d���k�!�m�RA$��f��$��x�'�?I��Rh�3ړ&|"0!�QEI��GVn�y$��̿
�PIy-�3I �]��Q��j�$<���7���A|�)\`�c&�'����".%�?$�u\݄��H$�̺$�;=���{�.�w��i$P�6�L���=�)�\���ʝ�yY�l*܌��O>�硫��Wd�|=D����h�7ڛ$�Og:�K�{6«�g�ؔ���&�Iy,�����@�J͠ ���cI�*~�������c���J.G�'��(h�]�v�p={��ӿ��N�)�o�m
�aa���g�FS'��!��[A?�{���7�Y)"w���I~����$�a]��3'�l*0�a!XF�I(���I&g�ʄD�=�޺%�N����O�$Ns���;���B�H���,ݡB 9�������� �ɲI ׷�HI�$���S��� �I'�$�0�[wV.�j����:O�$�7ۖ*��k�!�O��$�m���E$����m�a�{.��x�"%l�-��崕�eԌ� ���]#�5e"f*G��<<4�A|�)\~���&ɪ$���� ����P�#���@�Ķ� L�r�>W�IR�m\�a�K`G���gV�9L�H:$�D���	 a�����J��s���[�4&һ�D ��_db$N��bl�8�q�`���w�2��
�6�,���Q��������H��7�TTk�ӗ����*�Z%�z4<5r�TLW�����̘a%���t�����P��`1ąI|RH�N�E�z:N��x
�L$��ܫ�%��~$�0�U�_L�����⸒o�d���x�7~�E�$��3�nIwS�csc.�D�۷wi/$Z�ȻE�Y�(%�h���-�dH��*$�(Ȍes�bⳈ�о��o���f�T֭��U9������
"H��W[����-v�U��H,�s�J�U�ffeQ^��'/ݗ*�z����TBF9TK3��D�hZ�<{�ti����LZ%y&��*��I��b�4L#��U�{'{y���~@��+%+c��a��J�$�4�S�OĀ�-,j��	$����h�$qs���V��H�H�� 	�l�(f��3�|��I��b��H�s��s
�E%ض2����9Vgtx�_\��.w'�'���j�/\�n���_QI���ͭ��u�qKkf�<�iY�"f�{��L����mϡQ�KA
����p���O�I%�>uv�WPQ��8պ��]��	$����^[����|*ʖ��#6z�9;0;k��u�x��
���ak�%�Q�e6P���5BQ%� �y-W�a"KM�H�I&��� 9u���/*e�o\� ����1^IFO(0bE��UwIP��)L�v��
˓�?I'/ڭ��H-����T�=x;"�7֐�6ύ]�_*!#�V ω�v�	�PIe=������p	$���9�$=��*y��R %J�JؔL>�^���ox�E���JI �cuD�GvF��m�)���0�e�V�-��6��(�g�����I-O����JN$����y$Kɽw~�W�8��(�v��a��8�7V����x����u��Qdd<~�Z��g�^��\2��u1u��BaLnթPx{��VJ������]b��m���K	YlB���6�t����nv��7+�jF:� �0��Υ��f�	��gjNx�QR�6��;m�qf�49n�2�6�*����KnR앤x��F�G���<M�f�-+^d��)�:�2t�c;��k�����O\:�@k/���z�P�����;@[�qM��g��7H񶋌ú��8�c���4���.:�#)$�{�W�T��$�O5�I��۵`Z%%��"�%��`�z����Z�5�tH��rM!\l����(@8�wR�vֵ�1dV! {w[|I9~�]��Ii����;�1�%h��A�v�D�=�H}�4I�u\~s�5͊��	 ��Y���)$�7�/ְ�<x��TBE����7=����7	/%n�Q�$N'�i$���0��Εv��gF&��_R %J�J���$�$i���jo����š�2�7���I���`BI���d��Y�W<3�n�,�ǵF�L\��g��V/8aJ�L���Q�#�����ʓ"Q%�u���	$�>˛^Iy$�9�P		��\���wwh��Y~�\��������$����>��h��s�,��ua��OϹ��:r��N� ��[
���%�1>�+ҳ�7�ӘU�������� �0e���x'J9H渲m� ����>.E$RN�=���(�/��$�2����Szc�����#�}`*�B��O�$�4��&�4O�&�*�s�x�O���eʄ$a���!.�՛�*X^|�����받���?���R�� q�V� ��n�fM���<�Q�(�K��-���ȒO��;\�i瞳��+��i �Z�ʤ�Ao7w�T�6�~.��M�d���3 �k(3Q�T��h�\ĻJ�]���E�(���;'��5D���4!$�Ky�ݥ)Z�P�k<Ο=��I�-E�IO}-V
���]Ѵ������[�O�AE���a��5M(�h��9�-SJ5��TҪ�}��M+j4�Q����q�9W\����ụ[J3Yն_�u�	���KMF��b�e�O*j��ST�%L׹�[JڏC5L��j�8�M�}�˘�n���|%:�Iv=ְ�gt���4A�`9��)[:�@�Fs�íꊲn�R���A>Ug�'�,hoTR�f����5��չmn	����v+�ޝ����8M�κԑ|@]zVI�Q�i$H/������^��g-��&1�]:�{$9̆�f���]����]���-�]�+6��O*�Pöe[�o�[�iV�Yb6b���"��!l���є�2V��{���C�;��A��U�n4�����}v��*�f���v�fRg]7-J���**�T�s���.,W�l���<�t.�y�r��9�zT[��N��U��a����9�q(��J����~T6�)�ʏ0q��e
riݏki /9S��Sؚ<�岖衏3CӘ �{x�'��u�#�1L}ʬ\�#p;sf0m��=��:��{"�+����n`$<z�ų#�fJ�%s���:�`7Y����^�[Nm�-���i��c%�ys���8w�ذ��cN����nv\���ZD��n�>����e��|2v�/E��;_���f�K	(�v@0ok�32Vf��m�w�k��{}{q�Y���"�$[��oo�R!�3���I�G��D�N�ʘ�wU��me`w�q�����)��R�]��Q���n�o02�c��h�h�ѫ8*)?fvǟ^}�o�����,��V�s-���l�a�oA߸��<���H������#��'n*ei��rN�|d9ӅY)�z9U8p�Ǟ=y���CB��Yy'�$�4�'\����nYe��8�	�bh�I9�����x�9
�(�NNE�$4�4R�L��!e���/DUS��!S0�����t�Ca����tԬ�\<�Zr���ՔB�
.��R��QJ����;N�f+��
��;M��ܯK1S�T))5JC:U�L����vPk�^�����NT�R��y�p�*���eFp�ֻ���YEi�Һ'�^aB�q×=x�*q2-��2�"]=�N�(�<���숥ZUBDAyT��������(���x��!�T/?Q�RN\��+�3$�M!:jQ̂�[-/����i�LI**�]\�"3��`>�~��{�5�|��j���5I��g�2�4�Q��STҌ����m�����Y�S����,�i�N��v���'])�泜�3zk-*�����rf�XiSQ�2�T�5�w:ii�ҍF�j3~ǯ(������}�[j=&*j�0�o>ɖ��4ST��3=eT�~*Ua��5�i4S/��4֓5MP��5L��d�XkL��Q�]�*��մm��4Uc9ՙj��t�1S���U{^ƚZ54�Q�&S7��YE=�J���z�<�~��מ�|��YE��olE	�Sh���ݬ&��tu�wGa�Pȯ�Ϛ_���j�����{4K�o&Y��MQQ*j��S=�wҶ��b���4ST��>բ��44STר�N�;���\k���f�e�amST���&��潍4i�j�)o;:��V*bI�U�j4�Q��kY�i�EEM+�{��i�WM�h��=�:Qa�N�M*j4�5{�-�l��L�M*j�C}ϵ�SZ�J�����|����{	��2�2�)�ef��S�3�����3CE3�ױ��0�TҍF�5L�1�d�XkL)�j�)��4jd�9�r�OY��^o�Z��j1i�TҪ���ƚV�iMEM*t�f��k(���iS+:���%`�u�b饦�D��y2�^��\ii�U���T���ŽZj�1ST�M�3�ǵ�SV��4�Q�^�y�-X��?r^�<���(ѝΜ��[�g'�-�H�U=�l)�uV�:��MX�Cv���"�����^��c+u��z�%L���Y�D�!yF���>T�s^ƚ4�5M]�%:�L0�#Zb��gƱ�܆��4����AQA�OghU��>�έ���QX	�����2���:ii�4���MR�o����j�Q���MS�a^�y�-S,h������eN�:=I�JAPDD�;Lm4f%�R��M^$<k��G�>~�/�`l�������w�5�j���0���g=��&��ZaCT�4S)�h��9�-SJ5����}�g���4�=�������MFs�j�Q��jݕQ�`�����N�+Z�re��Ҧ�J5����Ǳ;�%�^}�[���Hb���4ST�[�}�E5�i����j4Owɖ���,j������Fsu3��{^�6Ѵ�5Ms;:��V*bI�U�j4�Q��kY�5��TTҍF��c�2�4�Q���T�kS��?b�Ҷm:iSQ����g��)�-D��ҍF���2�4�Q�f�٣���5��g�}ŵ9\��q�c���a���Q�����{�4��ZaCT�4�Q��߳�2�1[���������1m/s��j6eSJ5Q�e2�>�QOL�J�Z���:u�	��.�Zf�M�cY2�4�Q��Q*f��Ŵ���\�ghη����ҍFqs��֙��MST����9�ڦ5MS
j���go�Ŵ��������3�))-��>�Q���ZXtGT��y��/S�s���>Է�7%�-�lq\,^�R��>��3��̵�	�����I����Ҫ����u4]Mn�����nyC��e����%���%��1X�m�^�e���\��c��o�.�Gb�9� �-�8|��Ξ�c�\Y���|wŨ�T4���^J�5f0�
��T���*������ܒ���G��';g�m�G0�XJ���v@�c]V�k�hM� V�i�	�ëq�Ĺ����'��G=���R�X�Lں闋�������?���0͟�׿,��S;�{�i�EEM***h�+�2�4��SJ�2�T�_��4��'M*ge�}����s�+ks=�QMij%MG@�MS��9�ڦ[E5L�T�ߝT��u*��F��4�L��x�Zi�j�ST��z�~ҍi��/�4��J5)2���^�9�ڦ�j4�Q�eC��cM+j4��*iS�2���tFL���S�4ҦQ��oު��G�K�J١�F�]�mSJ5aQ*j�%L�︷�-5N�*j�I���s\��9��<��u�����j5��5C;�s�L-5MS
���5L����Jڍ�w�^)�Tē�4�b�t�3^�����.��޵�k�(�if���n��7T�iF�J2��|ΚZf�4��:iSQ��=����q��{޽��|��ڎ�*j�w�mS-���f��d��09���f�)�޽�4��֓
j�P�5L�1�d�XkL+U�C��}������)��4V��d����5LT�iPT9}�4�֢��j4�����������>�sgw}��	��L̥%L�b�%���T��\�%f*���2�������
���c��Z��^�M(ת%MQQ*f��ŽZj�Q��M�3~ǵ�SVҍF�W,���h#T�z���0���iF�J3׾b�4�5M��Y�Su��T�,�i�N��wX�rxkO�G���G�9��P�@��̫y}��>5=��RB�l�c��6�[=��r�%ދK�X!=��8/^=�dhq��9#U9�/��$�
|.�wux3�E��:e4��e4��|_�3�����L�M*j���O�Y���>�>G�o��5��ۑ�SJ5sf���qԪ�2�k��L�sx�Za����0���g=�`�ZkL)5MSE2��3z����o^��Íq�l���w8A���md5W{�:xX#�%��X�w��4�����Sؒ�g�<�1��s�Cb;��9o�;D�7�=���T�iA���Ze�'q��b�
�LI1��LCh��X��")@�w����#�|k��#���1�� [,`FA��;�^m[J1�L>l�>�>��w�#2�a����*���]V�m�vs�/!rM�cmŕ.+�7?�y�~���`�"4y4Fw:��[F�j4w~�5m(F��̖�6���s�w������X�da�v��v�FK�H�څ`�r��L���`�!�m(�1^��5����{��+ah�Dh׻xFZ-4F(0�Q�߹��V�bK����o�{������X�pΒ��$�S�48���0�������2�6!�MgV~
ah����doR�VܳqeĶ~�4c^�tf�Q��1�=]Oo!�3����<*+����u�{2�� ߊns�Ú�홮o�B@��{���`F�z�yE5m(�1Fa�`�!�k�'��r�J�3(��4F_��;�m���1�X��4�j4V*����1�#��0e�m��I{\��뚭�\��ot�!��a�c^�)�A�q����2�LW}�e��6�4�=�w�[�=�g9��v*bGz�;h��h�Q�b�5����j4�Q����
�[��������ב���+�@`X�e��T۵�kD����5��	aV�V"~�y�}J��6S�}���^�Z�yሒ�@=�sX���A;�s [ٿ33�݁���{�E1��`o���Zh�7�ˏ
�<h��#=�wcb�����71ù�ya����M���������2[Ahq���!���0���f��|�y��ǳ�S��y��!X)9XŁ�i��ְ[-��J1��9����A�4D�;3�6c��p��)��Db��9�s���҉�ҍFw��c-���)�a�0�#Ac���2�v�z5�#��$�k;���A�s�,�d`F��{�QMg;t�P�;�K�s}�7X��,�K�$&G �ǔ��U���r��U�S�ۖ�lɘQF,�Q;�ӫbs'f�{��|%�	�0�5��bE��0d�>1���Xe�Mh��_pX�ұ��ϊ�X�[���}��z�x�����7�^Kh-Ƃ8�Is��\�
�:~���g�"M��.-�c�0v�`-�:Wg�Z�[G�5c9�h[��k6�6j�F�P�y����Om�V��<1f���`F�Q�Ҍ�������Dh��wڴa�ƈ���~��5���)�7�����҃Q��=�s�[���aL���ʱ��aG����؍t���ʛ���`��Ƃ84��}́l�����C5]���1�dy2� �lU�h�G�>\�c�¬7������_�����m����4����#�z�;��s|'��,Ch-�"){��\�F�N�YF���vN�X)9XŁ�i1s��f�|9�[s@m�mA��o�-��F(���9]��bح�﹂�^�süޯ�ì׷��4��iF�+>�l�p����b`��h���(�jA@7�sl�#�9�ʿl���#�A�ϲ��bQ���YF��a��^�0[E�|/��R�$ �����Ϗ�[�ىm��J�P�h
|�2�U��ez״=��=%8
��`���z��;��坩.0���f0x��u�xx t˙����Yd�4�q�Y����-ns����!Hݷ]��{vn�\�݌Dnrq�����v�n9��^WF�nКU��\�h�ۋ4Q8+[&�t�t6tX2���R�tJ"kZŬ�p�,�6�,��.�[��c.Z��i�0�ԥ�3&9�y���E�16@�:��,�(���IGKX�-JY���Bj:8�lܶ V]s��5�o'��T�Xg�-�l�s���أ�6�OsYFV5��{��lCh�_���W�3:�X�H_��e�("8õ�k(ö�2j�6�;L�LV��[o��l���(�{Ü��xm*g����b��4F��5^��h���6(����-�cQ�m.q�}�>�w�U�[���2����r�)��Xvi�Ӎ���1���9�,Cv4�l��߯�vY�0##4no��0մ��D���0[E���3|}��۬7����#=}��y���y:k���!��F�O{�,k-(�����2[An1�l��� �\�<᷇��Dq�kz�Q�!���MT}��Rr��L���`�!�m(�iFk�� �����k�h�Dh��9�a�lV#���-�m+j1���#�@L��;?]��~'�ĦT`Mu�K�]u�Q�
���H]��BX�7��e�?�;��Hc�3�h<�Ge��yb H"H��`͐Db�d����l�f�o����&f��ej�Q�LQ�a�s�-��Dh�s!�:ĩ*�̢؆��<�b����vs�X���
ٕ��\���f�:M������EM�][��؞'7y��R���S�[tƤP��e��3c��� x��	^��OYiF�20&�=̖�[�C�Cg�9�j��"=�w^���a�-ׄ�>��$����B��@
"Ȯ����ҌCg���b��4D�3��\�����a��Db�#g��`���Q��(�g}��V�l ���Ѱ�Dʑ*%X��0���t��n̷�x�l��� .�dQ�A���wy�lȘ�S��Q��u��gՍ���F֯���{~��۬7���ƈ�_w����iA��ɿk%��������;��d`B���!��l�9��pC�F�N�YF�����r�;,wd�C{"m��V�d�4��2���LcM	�f�D�I�_{�OҊ���cL��Y�j(�iFk��LV�6��&��գ4F.^����&���)��s82�6��F!����+l����:�1��dbG&}̇�$�r��i�]��o�Y�`�؆�6w|�������W}��XҌC`��9���ӡ5�`�G�����8��<bT�XfQlCf}�`8�ؠ0�(55}�B�}Dx D" ׿l?�i2
���x�I�ckvkl�9�[�&jY�nMa�$L�(�ם]Z�"x��'���Y`���.�a(졝��<πB��_Z��!�C}��X�pDh��Ʋ�;h#"�\m��,PɊð2�b��p[*�[��ke��6�4�=�^b��4F��5\�h���F(3��0[K��s14�x!��[J��҃Q�|�
�lw=کقcr�,�A��E��yyb$���0f�"=gW�,�OH)�A=�� [-���׽��XҌCa��|/���Mk��eT(��"I�>�X;\q����Ma��e�2�mW�F��Z�����n0�t`�^Db5�� e��#�97�d��ҍFd`E���-��Ɓ뽹�d~���)�:�pC�Dq0�s��0�6Yy�]vJ&'1�Xf����e����s�y�g��_�L�pXu1F��;7�eh�������i[Q��Ҿw���c�uņcz�і���,l�����#�;3�d8��6"H��`͐Dq��Cd�����\y� �8���5r��eb�û�0[�,�ssϓ�*��i�M���=�ָk�ѭ�X��4�Q��wܖ�X����k|�Kh,q��1�ﹼ��~�>^�1��v�f�&/�헅��ǚ�`T��0B�k9�3�]t}&�^�ɹ���'b�£=��~����'���A��}�Q�cA�3o���G	���e�W~�e��Q�l��w�2·y�W	��:��cDh���Z0�m�#f��`����JF�j3���+e�=f�S��m�*������GL.Ukrh=�4���PKs���:��	�Lb��<i�m��yb$�! �9�7F!��ﹼ�l�����t�J�kl�c��0Ս(�Q�L9�s��7�06�����Ѷ��_w��alQ�i]\��֩�ҍ�޲�4���������!��	{��pCb���y�a�k��0���w���(�0��1`i�b�X-�0#Q4�PiFk�� �b�#G|����'q�ާ5�a�l]a�5����cQ��;�o�[g��`u�Y�����C��1��t�t�C`s~���A�2o��@�[20#Pf���Q��^��nsIm�l ���p[E�F�{9�o��*��i�lǳ��F!�ro��me�R�7=]�ѭmm�lﵒ�q��1C����� �����^l �����O�7U�;��Q�A����܁�ā��멊�^b�PL�w��IڷwZ�2b����us�&�I[��L�
�M���>8���E�D�'�\�6n���*DX�|Sj�){�seZ
����Ω6ʣB��Y�w�wR��.�=�lm̃�Vl"�-B����m�����U��[�y�g����h�a4e��0-ܲ+ӂ�[��Xv�@�a��v���@��na=�7q[
/�f��{u9w������K���]X�<���op2�'�q��{�j�19c��N�/f�]5�i�v{��gk	j�P�Ȇ���d9t*�eS��}�x�k���b�Ba��
��ob]K��2�oaG:���SW^"�˩,,λ!��t+�#+,U��l�,gp'u�*]Xz��X�B�Wm+Uݗ�锓 ��1jur���o+5���x�]n��h���{f��&/]�^	g������o�$;�o<�1K�'
�M� he�.�Y��Wӝ\5>�2���Y׺K���(�����u�����6��"3��\9��i�ZiҖK�Ve�����$�3$��h���7o�y) �S��#l�A���N�Y�Lf
�]���{ճ�$XK�Tk9ǖ��7���+I���`9y؍���l��r]�-��j h c�P�/�&j���:��o5Ӻ6|�i��dcjIf�QO��Vj�M����kRX�TNQi�H��:�t��"�C����M+3��u2��WK�$�2�\���U�b�(J',�H�-4���*�O)܋�l�5�iX�S1�DΜE��e�iL���F��r�U��9�W����ٻ��&Q2���Ի ����Q�̓��ɗ*�G,�D	$�йJ��Z�FB�qV�ADq}<�	0�er಺�|x�ʠ�KL*�$F�q0�ӠU撊[ǶQz�9���(��L�Bզd�rv葙VC�:b�Oz�HBåE48P����慩F�J�q��L��Wf��Dr�dfBE�f�����hm<�΢w�q�$�H膽���ץ��4�i���ڪ������������������jM*K[��6��I�֣1bݲŻ7f�Ơ�وL�Ԯ3��+,��2ۜf.s5�؉qT�U�X��e�K��6�l�ϟw��}�v��̲��Ze�6�d�I����� �{G8��Ӹ�mB=���йf׶��<]��� ���t{�P`�^�z����)n�7#tVw]n#f�@:��h�5V]�Xb������h�jS!�]�vxSg�y�-�p�np^�ٹzL�cO���s������mc�fJ�鬰���.ph�oV�箃c��4�Im�Ñ��c���ݍ�8Dskj8ܪ�!v��7X]�/Y5n����Ms��y��ӛgK��U��zZҞ�����$�����ۮ�W<�B�@k1�M�GnC�v��9�[ek�v9�ᮜ:��E���Rq���n�i��c]3[�	�����XMWf5��*T�PI���#˓��{z�d�ǥ���^q�6/b�1t����=c��,�Tbsj��kk� �1쑷;ύ�,��<u��;�k��Ԗ� !���4�6��d��苴7�t<�\�l�8�헍7a9�����:����ؕ\�N����v{O�z'W<�gu��/�!X�lźf�L�<r3X�pu��x��)q=so�y�u�ә�˷	
�ӹ��R,��GYn7�v��`�0oc��;�v�xL����.��3�a�3�Z�(�vk��9��Ӧ���-�������Bbf6��[P�P�l�3E�����ôFS�5GlG8u֎!��D����\$�(K��W��j�e�lKY�L0
]n��#��w[*�[4�;T�xqJ��Y�a�Wp[u.ٚ��5�[D��l��C;aq\��U��QUUW�;�wts�Ҫ��n��VM�5�9�l�ڥ%��۞L9�����8b�i���mݒ�+׷A�\
nu�=u��<�ㅸ%���&.����v�t�v22�u&W����N�R����ѕ둚�Z��CXmʲ�)j�[^�b�](9[.��iq�F�����)�j�궺%p�)��ۖZ,�\L����e��V�".��L�Y��k�v_�}�ko�o魺do�$�g�J+�s��b���x,Ch��4CU�jц�#�Z��N��Wk1u��;�؆ұ�҃Q��w�[-�5�mT��1�X���i�m���X� �wװ���	�{{G�1��{��l����L�w��0մ��n�|�?C@�h�͞��09%0U�1�ϵ�2�6!�r{w��e��C`j�c[�/�x�+}:�X�A�ﷀ.�� ��a�ﵔa�A��>�M��u�b��41{���ܽ��bQ�^�X[h��4M׹�F��c�{~�iz����4kQ�m-Fc�� ���x����̑��q����Q�"�	 ������{7���������ޯ [�c5v��ejƔa����0[E��w�7�Wi����W�t�G�(��.M:٣0A,w!���y�9��1���=�LbT��3��G�#3�� ��V�h�ߵ��YiF����̖�X�Aw�����n��HW��w8A�����Q�mkS1��;���1Xy,����m��(��^�]�}�i����⎵f�j�,�iw3L�?o[�ڇر*v%�>�C]'5mջ�)Ǥ�����o4��O�:�>��/2�{�𘭄�D#D_��F��c���s���(5^�fo�7�ٵl߷�C-�V�F*�*����J�t�DD$	 ���b��G�3����V1�J��NG+}�c20#Q3u�k(�V�Q�LQ�{��h��ы7ܷ0䎌1�F�h���xj�Wq3����-��Ch�޻���JF!� k��Kh,q��1C�����&p�͈z�#Gf5��Ce���Jo'X�,3L]ϵ�؆մ�Q��sX-��b��㚼N�^̫��6��ֻh�E�F(�1F{��iZj4�Q��;�k e��e͘����v�A�����c�Y18�ֲ�v�5�5�E�c�]��!P�Xg��6�N�2O,D$��9�7G�6O{���6w|5~���V��8�SwܣCa�(�׹�h���5yrݓ����-h���_0�[�O�g��h��u���JFd`C��2[�b �;�k Z�!��V��a��޲�=4�r�{��x$o�`e��w��!�cJ5J3���[��<��'æ�j����Mf��MOR��kz
���+�ɨ�ٮR��u��7�Qޡ��F��7�1'�ۜ��S�UsF�d����sY��0�����07ώ`�J�Q��J5�����,�}��*�V1)��4�hh̿o!ӎ�{��3z�{�b= � ���h#�f�����0#Q��{YF����6<s~��Za�(�Ƴx2�6�͚��0䎌1h������[L#�9=�d����w�2���i��5��%����!�~���� ��W}��Ƃ3�כ��_5����z���e+��j���=b�G�=�R���5Xe�"A���	�&Q��� q���E���ҍA��sx,b��4F��5]��h��19��{�g˕3u��Q�����j4�Q���y�
�l	�~���`u�Y�����C���I�|>㱴r:��Sr(�lƂ2o��@�[2�����a�iFb�5�׏g���Ʊ��Ch�0�rLbb���-���3=�`-��F��F����+j0 �@<f=�ܟ�ɨ�����Q��<Is��pC�Dq����Q�cA�)Y_I��lD_����"ȝ�����X�֓J5�eg\�lV�Q�����Q����F(�o�d�{Vy���ʛ�b��S��!�6��.�[������G-�����T�rDJr/34���y��N�v��W� k�/��b5��
�[{>�O�cu��LChĿk!�划��|w����#�֞��t��q�h#!�oy؆�6���sYF��أ���0[E�F�c��y��u��OS��vb�G� �fd�գ�I@�j
�t�W'mg1����7F�#���X0�(�4�Q����Q���FL�������	O���ǎi��܅gׄ��ǻ-�����I����J��VWˮ�^t�$�]��A;��Q]�]��1ݕ�����J�+4���n��|��>$�@��R�o���$bθ	�й�B�L��)�]L��Ք�s5��'�EH�n��Gs��ʊ��w��B'�c�$r�Iel�!&fwd���Yu;�N��������YG�~�=J��fi2���\Vr�]釥k��C��"T�}!Ӄs>������r%Q��D��$��!�ѱ2�n�? =�v��ffffD�D�.��~�v�����[���y�\������z�s�%6���UZ��V\C5:m�<�z4�Źu�I�<�w;xA�v���n5��.�x���u1�C̭��W��pt�{[�`n�0Q��u�Y��V[�h�Xʭe�]���,#j���p{o�v+��_g<v�q4�ap�)��]���!��h���$��#o/R�9,�v�b'�?����32�);�FM<�$��P$�<�1؅�L%�m���L'Y�� ]*T���تkY'����4(3ڝ@P���Cp��^�GD~W��v������mT�O���Q$s|��z��+*i����$�wr�Q�,�3L�2A�==���OV��3r�ē�[���e�DcBأ٪�� (״�Y�B��[ �����&��*�t�(߉v�U�|-w\P5;';Y�
�.��Rd�3Z.瘩^\'=prm�����t��i���%��d��D��ڢ|I�� �H��q@�۩�����ǓB�pX;j��F�%%=�n��]��v�<���[O�@m�.��'F\�գ{,�"Ft��	�W������귫���! ��<�m���L�\���|I���2p&��>�����ID�4�e
��u�>$�Rp˔ߺ&ɋ�>�NT�N>e���8�A�����4�d��j� ��f�/�iW�$��t��g�|bk5�$��U;L�*�
�B����M13ژy2/eB{�$OeUF�:B�s�Q���k�����}�e�b,W!�]E-�q�_��$Z�ҚM��U�E*����Q��
V�ݡO���9��xA��$vs�SB"kH}���B�q�.����@�A6���p�K��E�Mk� [��(��u�*�=����ϯr��WhQ�I9Buf/v���A&5�٭�9Ut�id\��]�Ao4�S,u�gU����n�� ��ٺ2����}�c�d�:�fv��0���V���_��xOd�ē�R���B$8�T���"D����(̜rI9��P$��ν^=��P�B��4�6@�]���y�� 
�]?/8$!T�PM�[T	'��
$�uY�����u�[��-.pJ5��(f]AF:����ۇ�keJ�2�,c��϶y+Y���_=o�����h�I=�ꈇp �Ml;��TO�#�]��̩��QE?�!kۺ��G�U@%��Q��4�+�3��t:�� Z�I�����
Lצ�j����I�m�UsL����jr�*��V-
�T��Ax�M���{�� P*b  ��N���fl�%�ò����]2��Vt���\�����8�'��ŝ�qM��=�ظo��G:)Q�}���;Ip�_}�𿉍�T	�O0�&�h�_�(�Ax���F�ra�0LgmP �y���Ԩga>�ڨ,���`���n����1�a7W\�e�^��Й�]�ϟ|�y��p+����x;5�B�����zo-c�s�E���=��|)Uڰ�����k>�u�@�Lz:纺kĒM�uD�oc�W���y�+����2	C�S10�$��kv� �'J�q�nU�u����"���B��d�6m|YAZ�!Ƕ�sɕ\�]xZ�6 �>�_B�{��g'��q�R���D�T�Vt��]�J@�s��u0�Y��=w� ���uB��=}���U��T�4E�eD���X��ru��cg6�X�]4��]�i� 
{Ԇf�&�봱�d��*�fR�z���Ѱ1�ބ������\�I$�X$&H`&�[�I����]��׬��Y�K�gh�Z"4�j[H�j��5���z-*�ɫ(̷.]e���4����}�'y�t�q�wO��v�A�=��9�㫲C���]&�%�����WF:r��[�׫Yk{p��nGvp=pS=��(�y�ŷ�s]B��vOl�:���!LalF��莺:pq����f�s�\j\�.�a��E�ߟ'߿�����D�s�?�%�ۨ/y�=�ܙ���q��m�
C�D��t�R�DL;���9I��F��Y���I'�m�D��u@�����
������`(�=K�s9Ƞ	9W�B�b�j��F�u�@�_s�@\�%bfeDIf��dd���,�E�.�A �=n�������h�G��*�CT�/�O���Mn���8��/;��@%�uD���
�Y�Bɽ������n��6k���nأH�<�3��7�Sg�.-k�㷈��`đ"f�5w�I;��x���ۡg+���>�~���;[�����#"D��=[�AM�
�Q�p�96o�W���X��(q}a ��Ǘγ*(7^�'��1��p�b9FqV�ܥlꕊ�e=s�;19gn����6Sj� ��4 ���РA�{���o�(�p7H���I��'�[\rDs��ۗY/���su@�����"��"L�E�纃��MBxte������{i�b��`���T�*����"�
��v��P�m�����0���ϝP ��ޛ"j&�9�e?~��}�p��,imm�m�[,�R�ڸ��ִ�Wv�%�� �]�_( ��~�L
��LN���"_�[� �{[QNgIUhUڤ�_��G�"�6g/X>�����kē�ޛ"��(N�ew>��f���a$�;הC�A�I|)R�a�s�b���6�K��WJ'אtͳ��7e���Q�Y��r�)ݖ�fi�A���b�-�-��fsN�sn�K-sÄ�%��sD�ȕ����Tvag��;������*�R��"=�y y����QPqV:�����X���y��%ꇍ��,��;�6��X7�y��r4.�ͼ��܊�,Еx&�������ҵӊzȅ�xu�7��pi�s*th���-|8*E�&k��$ݫ�rQ;�'Q;'v�s�oNK��q,އufnQo7Yx����Z�RoX�psƜ���eM�ba��S�cT4:���	����oY]˕91l�2���m���5ok�嵢̇��.TM�6p��LJ���(`���,�uh��F2e>}���l}Ov�ls3N�RM�����\�qr�6E�T�{^6n^u4�'��e6�ʈ�㸪h�kF��c4� ��+�z:�����z�m�)]�P\V�d��Y��J�!8G���w���YsV����WἺݳ��(��]ܩ�	-�>��<�*�V'2��X	�J��ݺr�ewTT8;�qD��U�4u�j���mX[�Ff�f��ձqYw�
��uy�p�Om�ۆH�7��^�{�$��8��#C����ɻ�/ҢC�f�
ܙ�s�"���7\6��;��z:�+޾GZ$��"ddN�Q#q�'�kv��("�8D\#�$I0��皈r����WJ ��D���ү��t�VI$$&'(��(�*���Rꕕ�IEAUH���)���"��UD֕i�¬�Z�DYYe�f���T�U�Q�\�j�	9qyGC�P�W��0�#��]T�4+2Mb&Y�a(&TU���CR�fi%g��J����bF���aJ&u�!�˚��8d$�Z*\�H(k2BT�	eDI�s�Z�u@��1
O�
�̐�7</I*��E$�eZՕ�YT�>�ʝ^7.X�"�2�����U�����%�^�Wd).�8R�R3���Us�յD0�)���$��߯�g��g#�|V�^9y@/��Oܚ�<�*��_\�ϟ³�X@Wg�������e�({���.����
'Ɓ�f������ᮗl�$ݕ^'��ta�Gg9���f��t^�	}��M�CK,���d&�K4��,&�uά[����ffeLI�5/�Q�q�$�;9��:���h&��@Z�I��v�Q(��S~�����g�ܵ��Lo�0�'��s�G.'u����]X�'���*�RR�x|v�B�8ic�}5���O>�"�g9!ƉB0��p��(]^�ӛL��^^9���w;.��G��EMա� Ǝ�]dLm������.p���p)���ò�͆\ᳬ������cTl��u��wZ��JA��>���ܼ����Z}v�s��n�����f�-'U�9���� Gf��O� �vUf3���'������c�n��J�]c�盈r�Ӷ\�b�R�f����>���Z��_��]A	�\�$����U��]̒�S� ��l�x��I�F�JW���8v��:��]G��P'ĝ��3�Z�{G1�3B���Պ%���@�yTA y������ouˠ ��LTr���*�
�T��{//�]*�I��h�H��	���W3��1wR�;�3C!�B0�h�^P�CΌ�.�te�oP�OV�P$kʠI�8h�T:�D���I��q�V_f�տ��6o{5\iv�����|���õ���a��ks��k#�W���d��4mʇwW��r�i$�J�]uθ���- 9��[%���ڑ�%�x�I���v��:�v0۞)�/�;�:��!�����*�Y��.z�^���,�i�k���:ȍf�RC��[W[�p�kTw�nCR�f�9;i��.�Osy�����86�����c��e�з8;Q�Y3��܃��7&�v����>~�vڳY66�=e��W��eR�u���2�L�e����F����쿵��>����U� �vW�������Īfy�gt�(��E%H�m|��d0�ffz#K��A#�r�B��B��^u�W���K\�"��b����TI9���c&��"�k���q��P:���B�
견Q(��7�r���.���&��P$���� �79ו�e�yS��K˛�Q�=eU�hL؍Wy� ���ؑԭ�=Z	�n� ;��(
��������#p�YW�7a�Ɣ�]+ך�`�z����M�i2\:��#|%DB�dI��ʢHqvP�I���률z�s�����4����/��R{�7@|(�>��^גX��� �!�[RŜU��m	K6'r(��Y��)��dk���Ǻ2EZ���N
���b�A��{��\�AΏ�Q$��uD_�vpH9���Fl
DD�H��=KZ��d�A<����T*o�x����(�����xu�R(+*@�y�q��U;��涨A �}���	��Ed"�f��,�_EڠH�K�>L
��	����
�Mt��+��D��O�>�'��@V����d�v#,w���I�w���)�����	��f���<
�a�٨��%����,��ׁ6�b$L胗|$�{[��$���C2����k{\�v!V�Q��&���""`�Gl�z�5aڞ�P��_@�va։ ��4	�'���{�|�:ow{o�U�`aT���JM��S=��n������nS��`�3;74��jjHK����T�sc���V�����my�L6v-�S�ŋ�����ߣ�I?n���ϲ�EGl
DD�H����=������4	� ��5����$��6�s��j�oA�9*F��E=�5�lC�&�5��P	�U@�N��	�EQdK0uIn�����EF�*	Q+��d�L�L�В�Ye;nsf�5k�?=���vx�j�=�	��Q��[�Y��o.��H�%Ͱ ���N��#�l��B�RR=��$�g/��:�K3��$���TA�ݐ(:LL�r�z?)@6<���"�X*�����F���R��]y`�m���|a���с�RT�i)=�9 =M�3c(�ﺅI�� P'�:��/v!]�S�r��o����n�l�ɶ)������!ks��i�M��2)�;|C�%�ZO:�'���U���������QQ��""e"�|F����~O�b��0��&�r[��=�t�fy��o��C<,�P�B�Wv�ٺ]h;fSn�6�M߶��>T��p��2ٶ3),3���ۍV(D�DW�5<�
<�I�Α�DK���N��@�O�+�ڥ�3|T�!O|�P�}��q߱` W�t���F���pnz:ni�!L&"i'�����
�(9�q'��@��P;<�I�W�j�XV-R�N������F�$����:��y����2�J�p�m�>��%B��II�K����u]-�d��]v�Z��qD�|�6��H;����!�+	֧����$�����mpǂ=�L�v�`�W&V��U�KV���#�f�XU>y}W�"d�tq�e֘t�O�2��O���آI$�AAQ�@�47jbku���LU%�6\�%Vꦺ&r\�\��.�i*:�\��Yh�Y��+3L<��*+���`�f�X[i��r^72m=���put����g��'),���(���n������0�xм�2%��-7�8�Z̄B[��)�GX�B.4���Y�Q��M2��
�`�.���Z5�e�#��ڍ�s4n��[R��L��$�#w�
D�TO��M>�$�I�Α@H�n�1��98�~zr&0�5�/�#mjՒ)�ϝS �����"Nvԟosf�'��{��a۞�+�z�P��0�T�C~*}&L��ڠI'�]
 ���f4�ۍ"���n�����x�բՀ��I8�f-[�X?_��,
��8� P��ㇻ#c�@���q|�\�MQٌ
(�
$I�����Aӝ�鞔���1QN�ĀGk�	ý�@�c�f4�[���ߍ�6yP�ؔؙъ%M�A��,������$�KӽB�Ȫ7�ݥ;�^�B�L�UGvE�o.�H�[Y|�I�';�J#cA
D�TO��=�$�vH}�;�a�,�����	l+yZ�O����܀����������3����;�П^��U#[Oq�}�s�$�Gn�P�1w�H%���*��I��
ؓ(D�D]�juȠp��|H4+�棵��b� H$o$Q#vE-R� �*}&LЪ}Q]5�.걺�3R	5ݔ(�kEx�{3�L�Ȩ��޹��F10J
�	�ٍ
��N�����0
��u��dP �gP���>��{x�I�mý��^d�x7i�j��X��3Z��*[tB%�ԓ�uƅ�Q$�9�s^!�܊���;P����Ȣmk��DV�0�bB���)�MmB��0�����{���ٝ4H=�k @Yf/%v�Q�5"RJ'�3ؐM�t�$_)m\�]^^�U�Y�]��v��뙗!y\o+1��1����"�����V�����.j�{���y���<�쥜�ɾ�� ���H�3�n'��\I�"`�]�]N�++S�=>$�t�I�T	�{�]4���d��O�uհ4�Z ���A6�����T����C�x��P���	�������]�F[��t ��n�� ,6��6��h�����Űu�f�+lK�Ͼk>}�I\���;�R	��>�F�����ܾv7ڹ�>��6cU���)mRy�t��Υ����A���I��
�{���9����b���ȉDD��MK$��(:���[f��b�,��:��s����2x)	(�#g��w'�Z�,�]4A=��@�s��s�tw<2������d�2��t�%Z�l@�V�����KrE��Оn������vxN>��&}v�B�X}e�xYYB��Ԡ�L!z���
�;�E��b�hW7TI'��
wE�s)�5/`��z��F� ڠUq=�^762�0g���^|!ub'��6͍��~����9��Wh ���@P���СYމЬ\33;�\
W���m��3ۭ��P��}j�"�EH*�����Ď�>�^A�	��^�޹��Ռ�T;z�����V�)R��΅
��lP�[..赜�Ē{yРI;�EEI;��+wiM�k����Tr)�^�N� (L�L
����?�x٭�o��)_�[ĕH�R�1Z���ᙞO��Z�[%��wB� �w"�"�:�Jx�3��C72�\�a���i=��d,ǂl�͌�[t'��&D ��6,����2M�m��:u1H�ŝ��\�rNK7FsZIeJH����n�fQ����c��(�s��
/+���-a{�K�_R�*Hl���)ge	�}6�R��]1X���ӆ
�n��S�`�o+g]A��}�2�R�+��y����Ns%`GV���Z$��tQU�Y�c��F�%���ۍ�����|��W�-��{ �8vV��t����v+���]JXʬ2�UEڠ__G��	� �Ѭ����S�'+�kܩt��K�(N굕:�YE�bDd]>�����A`SB���:;�^~������%�Ǽ9�x��uKn��.�W9c뻁fRՕ�4;��h`V����?��t�]F��KCr�ł��J�Ō��Xc�J��+"�E�,əW�5��s3Gu�ھق�nص)����|x�NUt�>ƺ��:p��f�ԱaXң�3����N��������pmmgM�u5����f�LlD�p��4��0�9�����C)$�m��c��n��t��p�[Y�������_Q���/G�w^�R�:��|議{�	r���ۗ�����V�x�m�;Yt�e,jv8��]^����Q����+�Y/fC�z��.��=:'�xOf>�����()d�(���y	��G�|Q�,�T�L�X��#M�&&WAadY�ZQaR�YPY�#TR/��q乪H��W�%��h��A��*�J����VՅ�I5sR3-,YV$-E�9ԥ*���h����jV�`�Y^xw+iV\̱�ʌ���AUI�$1DD�͓IT*�"���r��s:D�Ue�fʩ���k�;�Օ�(%�A�-BHI�	~(r�"����)
|q��Т*"�\�Qs�E�\ �9(�O�z��(�@�ҹ%�1�Q��B�����0�I$���6\(�6A(��ּ�|y⪪������������������#��[
ʄיte�FA�,b��{�#�jW��h3٘��]����e�2�H��VV�fLC�?m�փew;����<Qi��msm���V6:�..P�#l� �gaHm��:�*U�љX�f��6��u��	�*�M�V5]�Yu�ckSJ���Xu�,���j�h�����Y�֒�`��0�"	�n+�<5�x�"�5u�:�t�����(�M �m���b�z�pm5a��b����۝!��pW[��3�s�B�[c�W�ڶl��.�V<�61���5�kr�V
�J!Jf2.����v�y����1����������vR6��\]-�
Y\luW�'���xe�A�C�y�8��ݱ��(<�yn�K�[v�f<�j&�[6��Wz�e�L�hՆ��M,2�FmRQ��mp��j�V�YG��=�Ԉ����I��Ԏ��_[�ξۋ,|�Z;����)��+�����M�m�K-N�H�z�
���q���'#f���v��e��0nݵg��C�.I��S����\�Xl=c{�����c�L�����8l�sۜ�O<��Z�C���nj^�3�qF��]q/�rF��������'kqv*<��e�X��6�mV͒�ù؎{qRiA֕�mV�䲙��]rʗkF����0�sq�O�;v�!�뚈�l3�{e��0O$�%�h��������=v]������[�< �����ÜUFFf�7;X�a7*�Gt�r�W:�j��-�lR�ۙUyO��ܾژ��Z�(���@�L�UٔƝ�����d�iٺ���]��l�L�06�j5�9�X9�:ݓWd��`�	�y�jcWL�ګH�bd��UUU���*��N�2������&��H������'1��"�mA��)3�����zw��ts^i��68�p3s�=j�JKtv�kd�%��܌��نj�.��7�Fz��2���bɢ�um�7�W\�i�jVl��qPA��m�Ex;9κ�Dt�KP��+L�0Djhjh��a)�3��:�X"(��h��٩.��K�2�4�%�,-j���0���Ω��������/�b�X?g�=~t���=�LG��Sfz\{T	>��P$Z��D$i4�̀�6����{�G�\�ۊ�H�Ϊ#�{5C��U��F���D�2�fbn�̠$��s@�H3�[�'Ş�@�^�U]Y���$�3��k6]���`��H ��H���@�f.n������h�@�3�Q3v���/��i4�	w\
���	�n���upr�\-B��i�y�ܶK��闃7Q[Hh��n�v��F�ƶ_��EH�IL��:g���Ffl�$;�� �u(��38�Y�(��6��䮆�+j��Jϝ0r}j�t�� �����=6�ﷹ;�]tqw��φ�E�E���ǎ�H&�,W!��ӳ��B�5c/^��z3k�3���~Ϧ�#�8�ۗ9yP�"�\x�8L2����Gf��	��$ؼ��y�fktC���(Ev���&իRP�نs�2���C��>�$��TFz_�c��N�t�h�n���� ������	:s��ƹ�)I��}2����z�8{�(��&dD�nc7�٪MRf����l�+��i���(��a�Pe�����*B�B����YTH^s� �F-�*�`;�6_Ux��uDD��d�VIK��= -���FBōxl_K �:ۯPŽ�@��z0�d�N� �	�"`�]�jwhQ��; )��f >�s
�3��~�{Kz5%����9Ok]Ij�5 �Yڟ��\j�	�m��n���qs"�K���Aϵ�	���	��!&��)%�NOs�z�^�P���� ��r�M�u	s�Hݙ��>5u���Є�&իOE���B����_k���x~���*�]:{<�Co���Pr�r议���0�kJ�^c`l:`��d�3a��;�ߩh"
_xv�� p�� �&�U�*�����4�U���F,y	������Jo�Z ������}x�c�C�9� ��&)��S�ԑ�y>dDr����|h��u$y�"�#*��8�»s� ���z�3������L�^�1����j�xv�#�A �c��>$�v([���yrj�Tf!BG5��3�_T��ۂ�I`�,�33	3�����S;��.�T
.T�C���}�Iټ��#W�!L̑&��@�	��7$_f�M���=BO<�t ��U�ٿ73��"�x���.���W����u����`vbL�`j'���DI��bbw��yB�$��@�G{q�>�1�Զ��r`��l��R"�TU����ءs���{̭����Iٴ(��(x!j�E#f6D�M�E}wi?y5�*��On'�>3��Q2�&�uQ ����A'Vȅ*�����0�b'��$�oMf�O��iٞ���Y� +97O-�U")!g�魏�}���훾����;��=�(z�Nw\�еO�w^�̚[k� ��/:a$��	� R�����*i�&�Mrü.��EL�N����Fo�������UU]�Y�]���%Z��OYl]q���eMu�Ɯ7'`�s����n��bp�a6��h�Q���!��Kd��b{��=���a8qj](	B��cM���y��9p�֌�b�-���k��X����]�L؛jsi�h�-8<S�og&M�넻Fl6�9��ێֶa�+4kH���L�pL��V�cW(�%�uhf�t�<-s�܊v�9$��?olx�8L*g���V��	� �vM���K���Q�o����m�1�(}��]�@ڵjAW=����wJ��T���I$��r�Iͮ��&9�28�畵��Ԉ�
��k���w��I9�S�����I%��@�w\׉����.���Ҟ��ʘ�μ nU	/:��73�� n`�[�h$t��}*<�DL(�3���r�E�t�'���r��ځ�4��|��vg���_/��Q�ni�\Tŵu��4*S�}OV:_@�bj��AQ(�3"%�+���$��|k�ТI��@�}ٝB,�Y��u��={��s
���Һ%�v���Θ�q�t�� �c� �eCE� �7�ksv�@q�W���K��j���k���B���&�x�׻��UծQ�l��&'拓H��4$���Q �Zr�L���t]�
��IH*�����Q'��(����ödcy4I>��ıԈ�k�Cݐ��~�����xEK�G���3q�Ggd��ˈ�A��V ��k���Y����n�"��.4�I�?n�����(���tݖ�{�}ك|�U�JV�B�s���]81`�T�+�c
bYRWJ,�OϿ%�q�&B����]4	7��D�;;&��a^<ɩa��i�@}^�k����	Q_D�^�5\�R0J��nƿQ �H��D�w;+�	�܁���g	�N���`�����>���T�z�(�!��r�$�~����P�{7�虼��6n�O��2;ʾ���	������N�9T1u��2��ª&� $���	?g�5�V��"�S3v��y,v�W�Hؗ5�H�@��^���_ރD��ŗEg��X/ DZ�k�뺠H�y^��զ
u�|	��@�=�����h�Rw��;\�������\sv�N�1��=4��3B��a��"ثr���L�bQFL�{S���r��A{�4�hs�l8���W� ��t(�OC*aD)�oK�dd]��Fwaug\�|I8��H�����:;#a=[s�ۅ��`��ib2"DP�٪ݪ>'�fvP�H"2;ut�A����I{�4l�G�%�&P��=*�vk/9���w9�*��$�y4H$]�U��3�$k;���2ͼ��Z�J�]�iL�Aot�ws �9�*&hѡu��k��Փ�DS++-�E	]����Ք�����ýd�
��IH*����C���n26�Uق|+{*� �דD�}w�@�[���O���Bfd�& q01��"�48�k�v%�J�e�f���r�^}���]F��O�빣盔(w�T�i����ʭ�T�T�C��:�>ih���Y������21ᖽS����5� 7=?��;Θ��� )�����Z@�%���W�k�c�L�`Q'Xszt���X�t���h�����jT�XF�җ�J�陝��ǜ Ϊ�$��U�I;��ƙ���hD>���%��QAK�ֿ6 �ڗiEI�l�jf�y�M O�wΫ��ۻ�7��jٹ^)�K���kG��@N�U�n���nf,E�Δ�:��O�2G�;��rov�9W_��D�UWpJ�i4�١G��ZL��Z��{Rq�A�n�B={z�]������@A�88�����I�1E�\���T���Gn��/�GnyLe厙���]Ͷ�-�L��:�2�VX�ml��6��­�U8��]F:&�C�N��v@��4���RkQ��C�VR�i��]�s[���E�ĭ��ѻY`f:ǆ���٠E�T���m�rG��7ߤ�b�S3~N��Q�#o���I��c�!��b�-���]�$9���aB��}�8�s����^{����&	� �7>ۀ��-�Jy�f&&Y53f��&ͥ'.���	���P�tNR��t��}����oz��N�sJ�ԕ>>��5�)wT9�I;Yrs�`�K޹y��R�y�U�P�e�2&P�Bz���� ��t(�yYHw�B�Gsr(^���1`��R��Q8pkQ��Qlmc�י�
!v�xм��������)%�I�&|�r��Gf��A�a�#�a/���X��Y@���OY�v.¤U����c�q�{�m�CnN~�N�Ż���w���Z^h��>��D #�lKq%S��9�޽�'��y��?Gf9������ȣ$\ϼ[�:LY@k�7�R���|�=�s����r�@�٬\b�A �t�3��$T�06D�I(Q3vU���f����`��Ϊ�� ͉��{<�u�/X�3Mv��5GLT��;L�$#��
$����t�\1�O��7�u@��o]�x�E�uW��.-X���b �A\$JB(�E�=�d{CU���]�x�0y�2Q�?<�f�Ⲑv��4��I#9�Q$�}�T	�a���یG[�@��s]�{ �)�*���@��H+y�����Β	7�sD���ûƵ�j��/n��6��v"�fj�"72�H=��"�ヺ�!n���_[ʺ���v�!��8*!gC&���gV�<��ם�$�r��u�/]*�>�{�Yh�%L��u]�7���2[��B^�J
���D0�9o�̃��pc@s�u�m�z1Iq��F.ݝ*C.@1݌7�<�-ʹ��3��@mg\o��ק���}t�*�{6m9�At(I�ÂЛF��v,����x�%ʩg��fD$A��rƌN��i�ډ��Z�S�kw�]Zfc�Y��\o��z���)$�H��@p��2Z��W��hN���!הXշ�w�|-��Z��ݜ+
< g=�y͝;���;�����=�FK3��Z�'J��_ћ�2ȇ�U�N�߻��:Na����ɏ\��T/U��v{��}��>O�� ]p��Y[�Wy֡�n�n���Vj��H�z��0'�!���+r�#���a�� ^�A�`#
W	�X'wkDAY�]�0mnCQ�WKp��h��3�xf������Ӽ�$*u�v��%��ht�ka��kAŉ����1�gnTлN6�rN͢�ѻ��S_;k���ST`��V�D�/�khgY�՛�rwp����xE[�t�U(n�ᦙ�q�&�ˑ�ć�U:}�s����	�Z�ʹMu��+��pދ�B\��â=�Ú��8�`ɋ�ܘ�"�$I �T�J#R�
��QEI��:�H�S$����R(E����֨QF�Uy�at�9!2�J�"�G�y�PAGe�EYbY���7AUg��
9w2T|D��U}q��YV�bR
���Re����*AJ�Wn�:����w
�%��r��n����VY��ȗ[�����r%陜��+�O�<����)�(/8\�.�avU�AVI�s3[/�9TETWrTJ��-������� �*�X�Ȃ%h�$)!ȇ'!�	7�ȝE
y�K.TfF�Tf�g*�6�V�"�><��3š�B �'/a���Q$˴�ꊚ��s�*L��\��EQ��B�r���L���|D(Q	�?���~$�v�� 
������t�"��>��҅�� �"�ТO���s�/iu�ݯw�R�kh
ix]r�Q$ٴ��qӠ�����ʠg�� ��u@�yB����.�����B�A�32`"^t�����um �lKIQ���9j>��-�y�""H=�{jH$�f�Os�+4G�^�u�A9��@�pd.s2���=v��^�a��Cg��{.4K�u@�I�y^�0�`�q�qy�����#i4����� ���������5w%dWLw��6h'��VM�&bAT�I'Dy�ѻ�W��ު�
��L1w\�`@�g�O�t�k$�򝜋Ұ�szz?	��duw;2eś[2PU �����lė�;�WA|(h�孁���!J��B����b���?GJ�+�����8�o�Q �{�(�}-���U�vx�E+�E!v�T��3.�GQMa�[3(-�j��`6�[��υ�1�.gx>��$o;*���ȯ���Cr��Y�U�I=�(Q��ݔB�h:��{Zs�/)]�{���&��.����κp26�P�21F�DJ1���Q� <�(���1�V�= ���E=���	��g�����:ך;�� ��`P���;3�w�Z����/2�^�V��s��eR%ZS��{�S������7�Z˱� ��b �<�y-�ck��m�^ʹ@�����٬tމXs�ţ���9J��r!\��n�R25{%�]p��޿$�I$��h�j�>A4p h
^J���EıI\�i�a�Q�К�Ļ`;Qs�.�]zm�J��ƬV�y�]ss%j�K�i,9��`��m���1PI�5U.��X��5��� ��fT�@IB��]������:�l�1p
=�+հΝ����/�ڣ�;�q��y�c��I��rt;�O$8�a�k�+�ʵ�ں�CFh&��4�Dὂ��m�I�I��b�Ͽ�o����Q��U~�}��TA ��,T,�#��eŎ�¨w���`yR�tݥ%W��z�*�.[��A�����T	<_v�ڸz�أ
)�AA���<�P#��:ED�h�:3ϪtC�ɢA#�:�z���P2"Q��٪�f��x{��R�S�m�B�ٚ����6��':�lY'_t� =����f�*�K�� �q�]=!z���&(N�6 ;=��@e�/f��,���(�E�ـ�m���X�34X��6�ѹ�0�&Sa����S
D�13�D��	�� nu����OF��A������`l�w�R�H�|��"��mza��ݫ/Lv�N1k��+�G:�2�ѝ��-���!_)VԼ%y�%XK/w�c��v_O�U�|e@��UB)�;s߄���>Ϫ�>�>�E2^;�ݎ��t.�ܞ5=PK�"`5�7,M�ez�����f*ďe�#�6h�{/��P	H��*D�#Ls�̒WT����>;���=�l���:��6�e�^7� �.�p'��
=��x�"�v�p̠>���������ݑ�*��R�XS�=l*�%#*�e&�L�
��+�ζ�WV�g1\G���`����3��Gv:�A8���~5�����,�O�>����p�&�YT�V��s) 	W;�ٗȕYI.��q�ТZ�ȯ\ي�p���9x��*���_:�& �˦�Jqs���d�M+����
>��u��I��+363�Z�G,�OP��J�5R��LH��S�l_N�Zh]:��P���쿁 ��l��]�E�P*Uw@��RUr�0t��2�c%=�|	�ۑ@���Wļso�f�O��ˡD���DL�@3�(㗝"�(\� �p	�W�k�@�O�����w���{���?%;VK��p]�0ܬv?��[i�zD,(ư0��+������GZ������D�<�+ĀN^�P �����g �I�.���W!��0f|�K�"������_O��q��r���I��b��w�f���+�V߬݋*�% ��[�
3ɀ :���N�.�(=� ��N���B��Bʵ��:��N����闔$�	��TO���ν�D�Lq��ԙ���&b���skX]o._c=n�8��_��g�jw}e���;�V��%N��y/��G��������OtWodr���F�wO*'�" 6m'9{�
����hv��UW�|_9�I �s�Pb��F����ɋ��6���с�\���y���"�GFx�$�H�V�(&:R22��$r�I ��t;X|{2-e�W��Ѹ�oE�R ]��O����U���פ�.��A���	�3��m��ڎ��ȸ��3�.��{[�Q������`�-�s��}�U�|I��7�W^ٺ�D*%+pA�����W̐bof�$���(���� �ݠ-��L��B������7�t�+��@Rz��\��>̞�D[�@�NwdС��������^>x)��67�id{�1)��Z����Wx��@ޛ�f�Q���̽5=)��z�u]���ԒIm��bN�W���\\����+����ݼۊ�xvj��"۶�]כ���lj��ld��E���3"+6��=F���s��=��$ܵ�Fʶ3@ojB]��,X��Fy��g;s zS[���wl8'��駖���2b��..�\f�x�SCk����e�k��w[�[���n�&W&B��zΤ-�P�w<��cj��B�;3x�v� ��������Q3wVUI�ܪ�gvH�Emk:�/vt�k�"At�B�J����b���r�z�wbc���]z�s�'�WEBxC�]�rXQЁS$��P��!���h0:��>�$��s�&��p!�&g�^�\Ӽ�l�s	�ѰC7ؘ t�;�O��͠>ى���]���B�LO��juA1 ��$e�O����5�I�:�<�sl���쾨�&fA�]%H]e�2���
�n���K.�6�f˲�|���b������s~��*�on?�>�lx�°L�ν@��y"�Qt�D��ѳiI^]��|˻�+*%����<�q8��ٕmb}tc܍�X�e.;�P�x)˒ݳcH�z|m"���dDM����!o�3�?|{�&�$��>��$��6�v+�5��@W"8BS2�N�H�:h�H75���o�a �{^Mz���@��LG�D����Sbw�������6����>�z�J�q���d��@�Ԡ�!��"f}�g<H$�r�'�wq�}1>�ɜ }��� �=���i*F������~Ƴ��N�8��v a�9�<���}��u )�S1|�ܚ$�s��>$�κ��=��BQpk�0�:�A�z�0"	��$r:t]�nhާ����T}Θ�g�t뼋�e�����ݪ&���JO���СT&z:td8�4<�/)z�+<%����SF�v�1T��^n�JA���#��X5+C��ȱo�Ί9���i;^��8�uj�p/eo���
�����`]�뫾VHWiPcǩ�����{D�{�&�A'3n� O�>�1�C�d�㕃�%2IQ�5΅,�dJy�ə��$/:���5>Ȯ?+���o������;���Q)���duXY�,/m��fZ��T�Tj?<��l��>��u���}�FC�W[-T�>گ �S�DXh���)销���ɫ��t9޻���#[��4�Ȣ|Q{Rp˙������V�)!N�t��'�<�I'�ި��9�S�Ǆ��H�� D��v$J(���ܨ����u�|bj��˷"�$mgV8�Bh���TQ
vLU����넆���T�5͒}ܚ�r��JVե+W�i���D�[W@��r�zxR�����Pc�LP�c�3*Q���G�����h�+[�����U	odQ>$ugU�|����:H���(�B1R'ҐJSt �cZ�д�<C�<�0�HB]�`��0J�gx��D�9���VuP.30���w���"�彑^7ʠB$1LO�NWUf�X�}db�ɔ��	��"�;Y�D�����4Tϱ���c�4h_]]�)]��́G�\�!�s��;C
�p�:ݯ�����<��z|���HS��N�yY�6{�^�B��
�z����5�	>K� LCD�H��Q3Y�.�L
=y�N��?�.�@Qg���({=���|���VS"M	~9�y�&gs��7�"Q��J��dj�v����H`��G�nb�y��5bM�)p�'�6�S�Ȳ��-��N)CWm?U]c�9Ka�ō/-3��9����m��$�QT,��;��fY����LoW�	tԝ���o�v�#�� �,ei�}���}!� �zNwDUm5mZ�k��@���S�(��F�CebZ2mG��k�oF�K0=ܵV�1�xN�����n�[7m�:֝j["�ub�j��	pM�m��*�a��[*m�r�PZ��6>��r�&���pj7gw-�F���;b�=��aW��bѫ�O��W����Ա���/*���{7�o�&�4�����/7U��9R��̻.�d5� Ъ�[��#ytz�\}����3O]gU��Pޱt{v��!� �e����H5�iu�&�H����Nk�]�viޖ5md,Y�Wz^��5'j���*ZU鬰�z���cv��%�
̵r�oem�̬��3Gom��h�`��|��j�.Ar��s����$�Wr��}��8�8|u����R��R�!|7�_\���D��k��ssjVc�3o%��W;��&>qӈ���S���w9p�{�̀�]�MnmG�F�PD�ܽ�Жe+�Z4��ْ���c't�{�>\u���y-L�n�1@�b
(i)	ݱ,V�,E���;�r���/��[8�m8[��|v9�S��Ύ�̳B59�RɅ7'!�����Z���B�G����'9EU�W�i*Z���	P�NXrQE��>3�;�E绸meQ�9Qfs6rt����*�����P�!T��+�2�P0�L�DO����vUQ��:aDQ!S-H2,*罠�#���j�5H�4/U�8��#�\�3£�tK�.�$�G�8G�T�(��")��P��I�U�t@�8PY�p��r}^t˟�8��9ˡ�r�Qd�J���e�[�E9�E]���r��ds�^�\��{��
�*Q*Ӫ��eTQA*�ӈ�ǀ�m7R�e�v�o�}�UUUUUUUUUUUUUUUUU[Z�B�%�.�{kɝS�(�,u�s��fفҜ'h�bx�v2�^1���V���#6MD%s��4 �xH��S#s��ϗ��������@�t^���d�(xb�v�ʶ�;�Nz����0�pŪym��q��34�{�J�a�T�6��dr7h�˴#�]6 �-n��^ы�T1��C��x�%'\&���Jwf��:�Ó��]S�{<���h�ź��K�wT�2輶�Vt�
x���dݥ�l��$*�a[�]�-�R$�0�Wi����!ԧ;{K�DvJk�7l7��=����v�c�3�:x�c�#�m�pN6�vk�/)�l����f#�n�����H�3t��2��W��փ�t����pn�+QWFMF�S)5�F�-���Yu�u�c[3�s�%ʕm����:�G@a�n��^��)��۬g'��zb�K�Nv/
`���S��<���8�;]�1�fJ��m\�m"�ia����F=��[s����V�	���7Fn=#؍�c�Ყ9�ael��i�H�h6:�m��0Ąmf6 g�j[4u��y��n�x���W�a�j��:W�����/>�oFǷ�K�x�%��vvM�v���[ۻD#
d�u�������[�Ş�͆.ܭ�7�e#e�3k��V�V{L�u'%��`�5���M�����L45n\��G�饵�2�Q���.����;B�6���#��ؔ�q��.�4ɐqu����NZmq�sv[�j�lƨ�uGZ�+U����v
�퐸D�ˌ�&�T�	�JA���i��Y�IB)� Ŗ�����k)�]p%%�v�:^�������.���C-�Aqs��J6�am�B2������)������@�A����f�6���)R�-�8*�e���ڴ`K�U�\[�P�2g�52[�͍25���4")e�mX���G�n��c�z録�;d�A&Ie1�M.�e��[�"ې�v�]z6�^�e���\~Y>�L]g��B�b�+��'En;;���^�8���α��.Tɴ1Uɜ��3���$�q�����A���j�5-�5�5�r�}���ʑEXWiP�C�{�ʀ�9S� �g������)�łA d���U��Vڰ��O���Od��f�9F[R�=;�D�F�]P �fV)�w�Tk3]�8k�d�#A���T�mQ�k��	;��F�_)�mm�sb���N��DU�ڢ��
~̬f�=��r`#��݂H�ܙ�]�`$v�UE�8PHVRB��)$���7��b��{}��9�O���X ���h��mW�����).���Ǎ��q����%S<�hB7��v��ER;�H#`6�{���� L�wd��ɯ���a��v��A{ݳ��j�EXWiPt+�������}�u^EK�X��f!E��]��h��,�����c�{L;7U	�y�3+z�,G![v��sO�;�¾۟� ���݂A�ɠt�ڸ����S��7*��f!H*=v�vز�<�D�g̕ϔQ��.W]c'ď{�łO��ɢE�!b��AG�xL��npX�HV^ӱd�A��W�3�w+���֝ .{rUA\�p�uv-U�v����L
�f�!�����F��l���؟�P���g^�K�ޱj]

�
����hV3A5�[�ʧ�Lcp<.�p�k.��?�Q��R!L�û� �F�ez��'���t:��F�����( :n'B��$��I��<l�ƌ�av|�<ʔ ��ؘ;3ɀ.6��ur�>}:T�A*��H�V�T �/��3?*P>,Ao�"#�L����`�*�!G0+�CYE���`'�Z��3�2�[��< ��RI47\	6�r�"��� ��ɠO�ٟMx��T��"AQ�;}�V�[�U/t�W�<�	u�7Ax}�Ts�&�� ���AG�C��}�uط��/0�'�7�h�}��t����b6�QM�EA ZC����j�!��u�4c����l4������HUi]��<��|�ݚ�`Wv�dݍ�k�Бr
�����*�����F�س�<�de�Y��gh�x�$���ذLg�wv�{�:�b��2Q@6��Qh ��l�
�I�������uD�^�wd��eB�32�9��qx"F�@;w�@�H'��]�$�nE���V�Q���G�b��r���N����7Oˠ�^MQ뱐/Z�j�P���k3����������=û��'��[Ҩ��"AQ��~�����ѡydI�#B��S}���!�d��y=�{���SQ��.������������-5���f�m&s�}���٥�fPQ��x���v,��K���ϭ迦6���u@�|_�s�,�7�L�"U���,��뻔�vK�@P��v,�^vM C��b�G9��O��Tt�
�U�H�=�� 
��6> f�@�o�}0+�tNos�`��h�ai�2��j߹E�}�p��rH �q?��#�:��gٹ�f� P9r�_�@q*�@%iPb�{]1�fy1s�z{=x:C�}vH$��MA#�:��8��J|)>^��KeG� �Z��˱YX��TS-t��mX/��P��<��G�!'cB���R�$�I#c�tpp��!6�ݧ�W@�8ϷlaSvy�)�`�M�ٱ�3�%U{�R�-O�7�^��nR�^P5�Dꮴ�{J�6Fb"gZ����H��f���,��)-#�t�=����nM��e�[�D!��fILi	���l����6F�*�`��7R2�ЛA��MbѲkV���vXq�g2�gNv��XX1��uq,V�(Z�]s���oX��,j�!p��	k�����D�DH*}A�k�d�<�G�ٝT_Cz��������w��nvMz��t>�I7�io� z���ŭ=� 	 �vM	�Ρ@Vg�)d#S�<�\��5uv-U�v�O�N�1�vj`�LfC�zƿX/MA�ΐ�F�1"$DD�+��c�����A>':�H|�噱q]a��.h�a32d�.ͫr��:�f�[g��X0fPs@u�M|H/_;���uS��I���}ޢ�1�����XC2��Q8�ؗ��ū��4fPm��z��>���mPm��x���OP���A�/�;[Y�>��5=s@�N�t�"�m�F�����������m�:k�������F�a�H�.shf�=WoC,[{i<�y]�
#,:kS���#�2f�:��nVW�*;>�A��dP$����`�%T�lJ|z��A����<�����yD=��Nv� �{��m�٭U6�tFfuP����7ڄ�"f"M���̫9)?kn�Q$����	/�H���ػ[V��Y��5��Uj��J�>�$ ��ww$c�q�uD�|o7]�>$�y4!�x��%*UBV�" DD� �>�)��n3��:��b6d�yF����&�si
&/��(Q��� �����V,*u�R�7hP#�yݐb�a�$��I4Gu:�c��.ȑw�;o2��6:��	��w~$�ד��7Y/�b+�`y*�؃1O����ز���D�px�LTM��W۝��	��s�NS���؉;�n_[���-��v]3H�ٺ�V8u�5/�[W�$���$��&�7Ѕ�LJ<�3�E�x�^�A����A��h�{3�<�3o�O��]pu9�Uv-XJ�>'c`��T����3q$�o��ĂA�y"��Ρs\�����<e��]T��T�yZ68�tq���T��J�H���p�BʫTU����Id�k�$���4���/�G�컰&{S�[W��	b�=��������7Ҡ��;u0>�d��9ĿU��o�}����Wh���WݳD�y}4$��s��Z����ل��7q: ����.�݅wv�Z���b��}WC��Ă&3f�	 �7{TI%����a	�ܣ2`+�C�p7ϲ��xŋ��_I��f�j�]-ۡ�o/k�꾻���iNj��T&a���|]=�$}�!��	�@ǔC�IϷ]^n���	2zE�׵^$��%?X�^O=��X	�t��s��lc��iJ��c�ٸ�e5���=���Fb�T}�73+�H�"�I!��b�� bѫP���t'MU�ؿ+%�V�|=��@h`���ۡl<��Q� �^Ȣ|^�rP=�}����'�4��� �w*�NHd���زH$dl�[��D��sD��& lFLʉG������oVH� _N_1=��(
 n{�(wdV�y;��>m:��v����|:Ot�(
�[�����qzp+]�#��ۮły�4_��I���;q��(�n��.e��}�;�z�x�;�2��:fWw�^��Rzu�mT�e^��
�fe��+z��������?F�I$���
� r�t���mE"T���l`pv3�!�eœ�Z���s��,P瀲ڔ�{+���Q7k=��=g�zM���9t]o�s��r�j�E�4O��y�����]�\�������pҖ�2�����ض+�r[4�EQ�d�[�n���%n.˱F��1�g���n.M���mׄ���4�u-0#�9meVV���7R�����a7<����η0\����a,��)�?<��H9ۮ�;&��[���=�d�U�3=�si��TlZ���2P�ٍ��i�v�y"��� �|��%�d�'������Ȍ�\���d�)R�k���7;&�'/��,ފ����o]��/;�>im�� ����d�=u��ۼ�$��e�`�|{;&�'�:�F7��d�� ��ʂ��a�*�*	D1^]�����L�&;���&� O7$�
�>���{�:�xO>�}�$�^D�\!ϥx��d�Չ0
`6�K5����0[6D0�=�%�.��^��{TI�y�^�͚�E�=Ȯ��_�#�gbt'��V Ѝ��*/��7�ʢ8*E�Ko��}I��u������*�3����ے��W[:JC��)�n�<��]w�GO�[*��_93�� ��;W��g�� ��������mI���X�a+��Ƚ̡^��4An�X�����q�v{U:�����/�!�V�S}v��ﻔ� �ɺ�	���4I%�s��z��f�a���D�ݢ��$0I��رY��:苋�	ٵD�y����{qR��R��LyI�3sp��eGO8�:�ԥ�u��
9�<�1�0YZ��=�(�/3f�'��������r�wD��~$�wf�x�J�Z��"`�Pٮ���0gU�����A�Κ�$^w;�1�凕=y���B ��TLQ�$�}��o�:3�>t�v��x�i��v�H����PI�F��O^�[�z����%���i����-]���/��:�+2������Z�5���h�j��kx��kM�V�G�)=���.���)�8	�Пg<}�f\�v2ef^h�t��suH�[��A-��0Կ���!����+�L˻w]��}�K>yl�l���չZ+��yN^�wqh�� ����ᡎd��'�mn��F��&��B^�Sh)�k6��yq�Z��a��,'�,�,�un��u� �Bj]oYr�,�9Z�v�G�2���DG��V�_R���5'3^DX�+.`��[C+*����i���HF�9d�byրX�/sg<�E�鮼᜻�ӻ�GL������k;3�b���k���+��C�j���x���84���B�,w�9;�	t�VE��~�b���:��n���;/#&��^�؂�ej��zD(n��L�! ��os�8�\��Y|�vgU�ƃ��:+BʍdU��D�т�b�.*�T�Ь�k��ٗ�}��L*+��#1��{�ؙ���n�u�6�k�Z�>r�=Ψ��JZ
讹�9����r�̦ �b:������G��A�ΐ�8�
B���Rl�Y��4-�t�Į���l߱>ɳ���;�Nۄ��m����]�D��+�S�/X�,�m�J��h�"�M�6�����tsS3hub:�L��*�c���WC�	�TU�	"�w����z�ÂW��Y�sY�I��͕L�d�t�~��nI�BJ���4V$��8L��uG*��$QE�I�̨�$�zH�s��wH*)��M'VS�ז��Vp""H
5�U�g(�ʰ��%�訒���f�(�̒wJ*�����C�DN��r���VKs+w���� �����P�Wts�C�'(��<����+�=C�ˑ^��D"̇$���3ZDQ(.|�X����PQ̗R'2��#6�"�W.��vU�*��\����p#Ք�q�p��*��qs�DG*u�8p�z��S:��K���l��H>'������I��Тw�틶kʅ]�V�ʡS�=�$��IP���$��uݐK�rvn.�Us�y�~�l
��!R��V�S�{��P���B�R�=�*,��ڢI �|��$�{S��P��Ύ���W@�R�aq���ŉ]v�c��B�h-�j�G\U�[翛�X��""V��u@�7;�H��k������/|�l {����xU]�V��!�9�a��[4 ���s;&�Is�Fq�fg<O��@�)�AL���v��|x���zOM���]�$��vM⍈$�J&A�*��#f�U�'�k�Ւ	/7&�I#���y��k0A^Ǖ����nw;˹m�J�<�qv�|��^�S$�����sCAPV3(���Ko��Ǐ&E/�`?��*��Yl����
�C�L�kT(�Oٮh�:���!�wS�$�{9�w���˾��`�æP�0g�W�1�-8�#,f�˴]�[R[4�6e˴Q3��i~�3$�|&������ؠ ��릢k��ך0�{v#1��ML�'�HR���Wc�n�Wx���̺~�	��� 7ۭ� �4g*NQ>}�P�yj��+V>��k�'�S� 
�}�y�Q>XŒ�9�|{��W�PIL�$LO��;7�\궻t�ڈ�H"�h�/��$��s�h�.�Q�;6kĶ`߮��m*�k�7@ 3}����^�<� =��P��l �{$|�rEbψ�7h���n���۷ٙ&�O��b��9� �7TT����'1`��c��X�>�=�*2���1m�͑-�_�w�J���Im�Eĸ�ۑ�'	'j�aq�ݦN�*d�h�n���V�`Wv)a�f�ƺcJ�
��%X�b�7��ͬSF���n\XI�3�f2[wa��c ��e���5�-��K8���7X���v�&艜�E���ڑF�Ԃ��(���8��e�D���6n��[��&6�v�\�9��J�j���d�mnn�jK�2����0!DJ�c$XV�����j���
��銠(��4||�y݂����$����%��t��_�R�d�|7��@#�C'd�(D� �|�:�O�y���,M�ӳ~�3+Nj��K�*TQ5wh��5�(o�� ���0�W7
��x�'<I"���/;�Y�c"B�DL�ɠC��ݘ�ܝ�-N�;�I�]�#3��`ʠ=��O7`��$j��W[�u@I����;��2!߉��H9ۮ���sD�	�L\#`)��zD16�p���
�(X��c5���1���b8����Ŀ\�d(��&s�Q ����H$�r$˜�{�M�LQ!��Q���w���P��H�����LP2��������]pQn���XzU\@�����kys���p
��(��Xo���ۼT����	�ٻ�M�3^&Ș��2���YnG�$��~wd�3>s@��jr��6O�@G��T��+T��I�<�Q� ͞���X����I'��ذI���T�Y`r�EWv�����~x�H���I��J���7�1Bw�����rI���(U��O�����j��)+H:}�鏀�f{o�@�ux.���:T�
�3�: 	ލ���Hve#(���4�Sa��b�[��g�-=����3��i���A&:L�3�6�|	#1���}��t+a���Y���J 3;S�����JJ��]%�o�N�q~<���}���ݞ��	�ۆy�I���:����i.��؝  ��3�p�x�5��I��FS�* ,9:3L�M���M�}ҟN]���:���#�>�@�ܦ�ϷVD��f6���o�1:��ns���}sD�q
�TU �j�;=:�3@���}G��P�	6��$����Z�Wս��H��r(EN��"D*J�ܩd����%s�,"��5{�@�^�ר�w:#Fg{�sw��$UݑC��Q*�.�{1u�w8�%LڧC�K*WJ�o�<����Ww��Ϣ�7�sD�@��v9|�M�lׁ�ѱ�С|-]���pr��U ;7�v#�Of1@�M㺢	��w`�"�9MX9p��/��D�)�
<�L��1���N��zDl��d�$�=wB��β��%D�t�($�S��6��K.�Ox��\����݂A'���B.b�������n:`�.f9����i(2N�A�>u{oX)ܡ2硷��S��^���]������UU�5**��R�L��� W��o�S�yt��@D_e�A&�y݂H7���f�?=���[�=�PRf��%u�
��h���i@^֥��]/��
No_�T�PFͣ=^��� 
�:�	'�3�����Mݳ0���7�T	nw;�b�"$���U��ׅ7�b"��V��� �}ټ�ϳ9�c��AO�^����s��]iF�Z_I�}�,�C��'�*�+�\sb��$�y���Ng9�o��D�)�
<�g��/;R� �ӥ@C��0 �g����|�k��:y�Ҫz��H�M��3V�̚$��#4�&&#c�D@��r���%�s@�M�:�bN7	�b��_|A۞w==�w��CJ��J��/���z��\�t��q;�s�%�沭�M��d��
q�������bI%U��m�XRَ�GZ���%��f���,�I��sѱsFө%m[p�$�MvxP͡Va*	����f��aձr+��u�ɣ��.�;��]�ku֗5���#ɇ��L�En�^��n�v[�l�i�ֻ;�uk����x�˫��N���oa�.DaMV�P��g)�z=>�E0V�TsÒ2��1���-����,j�u#��27,g�;�bA�TLO������S�{�T�>��JZ�T�y�)�Ͷ+{|U��X�d�llW�V����f綠��_vM|p���8�e�b�
<,�I$��`��� �bb����iW���,�5�xY���@��ɯ=Q� 5*��U��}�N��~j	4r���I!�eQ$c�֖V���<W��RH�\�)Q���b�(���1z>&���Ӻ B�ȯ�ɯc��.w�F\�`�������*sP�j%�ubP�kR6�a���+)3����2	P$ʃ3}�&�*O�;�&��F=}v{P�r�\�P$�ɢ}�t���Yժtzc�P�r����s3J����N���4{lgT;�KpI2�>R�oh�k�{�����:���勧�,0�c�D���pE��(Q��+�?��,�H�aETT;��&_�ٵ@bђ��7@
���� �x'z�/'\
��ʠH$���ASe%�"ffUx�u������!���d�:�g3�7v�����nP��]Xڢ��T!>�ѷ�d�����I��¼��Vs������P1��ާ�t�l<o��@�A��t*�"|��un��P�{'8�kj�!�ن\��߾��a/�����*���f�@(3��a���w�o�	7���/.�qP	P$�@����H=T،'�ԁ���$R��L[��@����hZ�dV���2@)��:Tpz����%�� b]8k3%������T�&�����إ��{�fYtxջ��V)�����̽L�B��F�o��I�����i$�>���L��v��+%�d�N	� 4O����@$�y &�{���}�9��� r�z؟j�B�$���?&�$���L��ߌ^���I���J$�9�	$�W��Ŭl\�*E�+��;�]��zv�m�B��USKi]a`�l�0�~^h �B"H9�j��%$K�2h$�J��U�����A�]��(����I��:$�:�Ы�����~|��MϮ�_6���@4N�tI�I�팛K�ɧ�M���ô���iP	P$+�J\$N��� n{\�I&���x�C9��I��$�rL�I3��!;����j��6��Q6g��YS;��~>���D�9�K�$��Ui�{�3����Am��U�W-9�4q���e��s�;�f��[��$��9�N�0��s�Y]c3�7Ѓ����I�&�Y}J�T������;����˃3"�6�A+�2I4��Ţ�D�훵���́��d�� �"��իF�u�ق�d�����Gh�[�V�i0"#�ϾM����Fx����$��9��B����N��w��OE�a+����@&ۻ���� D��A�N��կ%��'��L����-��I$���wa"RO�f��׋��_g^��s4<���$	S0�\�����$n�c���+��^u�S��>i:$�Ng�J�A��N�ڤ8��� � ��'p�;у�+���M$K�ڱh�^M󛴐I%��9�͍�3�i�8��I�'�R�J�P�RJH��8$�M��Y�ﰿ�3TO�^srI$�ޫ�$�K�V�����~�/��?2&L��Q��Q��ccs��$���.	$��"_�11�_�`)ETYJ�> ��@����Y��q��Y�I�/F	i�I,��l��� p� "8'����d4�w��`��Ũ�Q �d"S�������HH_���Ơ�������߃��$4��Pj�/�A��+!���!��E��(���Z��7�

�F� �9����� y(=�eΖ]H B���q��~��O�!4���@ �����H߀�evqm��c�������~����4�$[!�.���^?�p��K����I�����I		���d�������44�/��P}�Q����,�QC�������C�FR?�U4�?��Oت�Me�g����/�C��?��K�Ze�La��~ �I!!5��eE�ŞT�-S�X���𲐃?��686�ö��� �E���R��?������">�I|� ����:$�HH_ -
�&����~i}��-}�����~��!D�0���q�k�>b3�/������������?�����0�������Q  �h�uR�?�G�Z��?����>��0(��0��T.��i���O�������~ �Q�FA��W�h?�|��_�/�����h��	$���|��Ƅ�����P�5�C�,�kk+aCL�� �������� @�MR���I	�����!�d�օ�87}�����$���6d $|��?�+>T��B��>���m]*�$����&�B�id��Z����B��b���]�LWQƔ����B�.�RJ�@��T� .-��[T��cx��I	�!����~G�^IjE�$��?�?/��I&E�|	rh���~��w� ��.�����}�(?g��/��'�G�c
��~���?�?�B�ޏ�F?���c�O�0RI!!}�澺����P���D��?g��x�C��I$���9_�=�?��/�������/#��_bB��#��_i䍚�[I0�3��p���O�����b��� ??߁q|0����tk�_��M��7Hи�}L��~K�BI$$'�}��V,~�����A�3�_��83�� Ϙuw��}�#�5�k��lȌ$���"�G������� $���LK����$q�Gܟ�_��b��~?T�$/�_q���C���������j$�u_��~ڬ�#��4#��D���|$/}V����H�
aP�