BZh91AY&SYr�,0�_�`qc���"� ����b     �  @ )@  PP ��      �        @      �@�x   =        �  *�  
  �         � ( P �BUJ�)  �J��)RH�T�*�RJ%IIETTEJR�
"$BH�%R%T�%R���T��� ����UTRB$�- g����cP�ͪ�UU�J+9(�b�;��U7s�En�"G(F衖� ���  �� C�r z��� �:%�!� n�r� �@ k 9L �� n�r��� =p�  (M� ��T���B��J�-4%G�l>@�����=�� �u*�` ����v��c�� ��� �W��0}>    �  .� �� ��ϊP���|��S�¼�wB��z��ϐh��|��pӓ�a���^CG��P�4(  � ��T"I!�
R
��p�vr 8����u ��n�(�ފ%. OZ{�)����<�P�z�Q�P݇���z��   ��^���M{�:��T8 M�@z���v 9=� �x�J�B��c��)�7Js��3`W��   �  x �P�UIJ U"+�҅2o�h!��� ]@�98z��{9
zê ��'��z�l�%R� ���SO{���i@P �  ���XuG֜@\x{��vD�C�Ò�wp��T܅%p�.LJS���6P{    ��  �
 �QU%�J� �;����DSv:NZP&DW���sb���'v�]�
WQ��Twa� �  �  w�d ��IR���!�������J*8ॳ�Pݸ@]�t�b;t+�� 
�   ���*R @    6LE%J@      =���� �    M��	TP 4   h OT���Sj� 4     �=&���4&�������24ѠڏjF�}�_�}+���� *�)������]:��[o��UQ_~H������� 
�[����������'�~����~vlS�$UE`�I�` ���b�"+���g��lP��P�X���C�"~� T�q�����������b')�
q�0��0��8�1C�P�8�1�`%1C��8�0C��8�1��`'!�"q��`'��q��3��8�0�툜b')�
q�b���*q��!� q��0c���S8�0C� �8�0�1�1�@�8�1�@�8�ClDSlSlQSrEM� ]��D6� x�C$ �`<����
i� �B
#� ��(���$"*����A��A� �rB �� ��)�"t�8�Px�x�Dx�x�@{b<`
<b�<b�� ��A�A�A��A�Q�Q���G��� G�TG��G�l8�9!D� )�*��)� )� �$"��b��` �!�DC��4�1��8�1�� �#�q�`����"q�`�	�)��8�N0C��;b'!�q�f�	�q�b�o���To<�a�_=緩�~w<��������*AxѼ�K��ɡ��b(������աۛ����nAX�L"�Ҫŧ
�6Id����i����z�9�<���
ܲ�8��N�u���m:���݆@4J��R����Yv�%��4��ݓ���u��V \7��e]k`��]֊���Y0e$ڙ���"���Y{r�w�b Q����U�,��0J�,��9�2���RWJ�Y�ΉB�H��"�{���L,7*��=i#$��hl2�5i�kI��d���DS�5h��E<��;� �e�7(Z��'�tm�7>zӕz�1�-����3f��6*D�Z4�m��Oo�#�@�A�ض��5�e1Vf�46˸E(��F�(�$�� �⢦S9�<���O$�5+t^L��h�r��W-��Tʌ�r�X�Q�P�i�����v˦mՀƙ���,Zr�Co]�36���Ӱne*���dT��:Ap����Ba�[W���e�wX�ǂ�P�Am�z��h�͐"�K{���6{Z����Ŭn)d�m����D���U)�mf��ՃM�M����Q\۱W����!6�ݕ� &jHښ5��Q$�(l�R�F��7TW�6����h����b�
dܱ���r]��(^�P�&N(��nd�v�V"�#��@�7VY�f'oV,�m*Jǖm;��5��#VQݣܳI�Q�h^�rDa�5x�S2֦�C��<�&#A��Z�e��{mReнN��m�#��1i�ۺ���wf�뻦0i�+wb"9��_��L�g!9�3B��@a�v�YK\�9����xz�ݡ�M�tU��3s޲ǷNY�I��e�D��7��Z���n���
e��ʼ��L�f�m��Ж��y���F��1��VАP�������E� ���V����P�ԬZ5�h�V��j�2���r��acA��h��dn���x9�[�q�󺵴�WH(��-غW��ld�h��ef�+a��'/�
�xT]�Mw<�`�j*V�H*���]Gb�Ų�&/�e���	J]=��j�Abi�ou�f�ܺ��8Ǧe��-4��0(^)=5�+H5�=ͺ� ��h�fT�t�wee*56��Բjv�]���Uވu);+�
Zb��ݒ��<����ed�ڣX)`g%��n,h�6&�)*ӯjT)CHXgcDc�sv�7f�N�Ճ��w�,f��	�L4�s��n�^��ۢ��
����7R]f�&�#��X��Qc2��U�@�,��YFL��,w���KWZU�`LA8�	
=
�2,�8Q̭̳Ie���1�qY�n��9@d��Eaź3"��f��{k�0��h��t�����*�z��n�"@��;�J7!@�F����U9a�m]�I�WB���F�꣑�`f=�Zˢ3V�]Ay���Ĩ�(���a�;$�4۸�H"T�4ҢJRJ�j��h]�X$��⬹$�y
��Y[��h9o��b�d���ZY;�rQtM�N(�Aj�JP�ݫ��f;���u,��VvV�e��w���7c�F$�;{���Ρ�t���=ìd�MV�3-��N�8�1��L1Y������-�r���n٩%��C%`�7�^�ȍ�dr&�Ѹ-ܩ�ijɓe�k+sL�dT�iܹcoh7�V��nI�
����Z�����"����A�6=i^MF�A�w�u�TӓF��B)�y�M0n������nJY�S7d��ug6���1*
<���d��6�݀r�+P��Ip*�Z�r���ܡj{7f�,QԲ�X��m�T	����|�Ku�e=�ʗN�`�O5=�X�ڵ��O,I���ڻk(ㆬ�tŅ������%e�2�&m˱���Z�rD����ek���Mi����*��%�<�+4k��b���l;�Z�YIkv\a�F{Zm@��[��[y�4>�!+
бu,���BA��
�H\�M����t��)h���n��oM�r�pL�%��l[�hx�te�I������A�-��[�z!!IV�N����,z��e���R�x3q[b����3s/s4PMHfQeS�0��%
̃CR�L�\D*�)#�+0���@Z�[���%={�]�eh�{�����{�`ue��v��i�H�m��/q�Q���#nLJ�+��y/6c�:�bV�{��dƫ=5t6��h�ɰ�����S2�K�`h\�h\�B�F����&�͔��[@e�d��Ѻ��v�*b�:oƛ�/,K���R�fU�Jt5�݂fMt̡��7vA��bű�`�h�.&�+�k	j���s.��J!N-�p+Ly��f�Q��^�[���UB5E��Ic��Ņp��:�L��=,�B�%D�E*��0.ɝ�5L���*D��l��1�ە�r�$M�3�2�9���VX���-Jt�U�N��,�=yE�l5cl4���i�Y�h3�fa��q��m�FTмv�VըV3�F��X�X���3X{j]�U���K��kv�R��1�&��zq�9�/u�2�2�v�ʺMߖ�6�D�~�d��t�z�a6���oFK5`M�N�Y�q�ٯiY�3p�wݺ�6pV=��(���2`�x]!.ϳ1�6���|�X�İ� �I���D�aJbY�E(Wu�5�L�X�%��6�(V�oj�^L:M^f��3A4-L�Ϙ5�e-§ ��#��A��*�Kc��˭N<�l�t��췇e[Ȳ�VR PĶ�%��Z�2-d���,��n�C%n�D+��j#0�fV�e!m�B���՜��4C� *���[z�-��9`��5�4<V/1R�yI\l�)�xYL� ӣe
���ܱۼ��pRXӪ�^���x���J��Hࡾ����Q.�Vq�"�ˉ��(��{q��&�����Y�ǎ7[��Iv'Tܽ)ea������.7/�oB�u� �)C�BEd-w@P��с��m�.	.��8���f������3rALް�]j�9����XpV`�ց����P�9*��/�w�"/3�"���I�r����(��-���m	��Fji�WR���X���4��p�0�� W��[:72�<�&�YX
Z����.�GW��6�lhє1�%mkak��b�kCP��/j *�oo<������V�
f�w��n���Z��E���tj*򎥄�� O.AF@ ����]\�h5�2<�if��^T��y3�����G0K��uu�pMѕ	)���`ڞGs�5/-E�f+��v��t����˹J@̺�U�I�-�V�f���ux�i,��ڷ.�S�U���=���`��	�[N��6ʭX]F�Z�7�YT{Y�g�j��NR�,�Ū�b�VfI��3(�ݢw0�[�m�+S�v�*��ɲ���D�3wS�ʈ;²�z�n�ˉ�YuL�ǔ{��`��yz ˡ���s�5ֺ�
��k�)aJ���!m�ݢ5�/n{*߱g u�',^^�kѻm����fml���Pk؃P5x+md &YOn��^&��&�j�y�J���][���[`!vŽܕ�J9�s[{�F%B�\�[��-�4q�6�߉��ʬ8f+���ƨj%�ܕ�1���$5/0;f�i���zQ!�knL���U��2�&i�z�k@Suq��^�P�yz���2�Qzr��4-RҺܨDע� z34�l������d���ޖݍ����3o�%��a��bY��.��*���1���I� �&�x����Pa@��׳%֦\�p\��5�9H�i��N��4JU��T;
�X��p:IT0���6�0ᕰ��������fP�9�i��4z�J3!є��XY��*�T�%�@�� ɋ�T�P��V�k1y�j�;��S[*��X�j��^:܇J�)�{sC��٠���)��]^�pL@K�X�ޜ���5�c�Y�`'Q�-�;�.��sh;�O��R[��V��̧�]Vr�/ �{�<M��+�Ve8��YC6��t�Q46��in�-����PƳ#���{���֣�z��MwL�i",љ*���N875&�d�3��b���nU�ܕ��d�8�bZplDQL�4��bnY�6X�8��E��csHĥ��2�f-�Q��0���J#י��kY��na���ŉ�@i>-pԘ�����&�5o4�W�j��[��ջYZ723Ce��ô�)S[���� �l�n�Z�����.(Vi�c��6ƹR6H#D:f]�$�%�+6*{���=�:�l�[w�mm-�2�<�RH�ov��7{�5B�*z��l[��uU�˚v=���	[���n��#��;KHnb��(6�X���ܩJ�K�p�؊��ऩ�{�X��HP�(�sp��V4�Û�;��0���WpK;�@�2�#5a�f�����W-ի��
1��g��[���4$I˭�GFI�ټxD�6I��r�Fl���� nV;�%�Lc��fa�7`q(��ȆVLCtͥt3i]LލݛX�q6��J\ B�M�M?Z�R����k�bD�١���N�^Aк[������a̳K�F���Q�z��/kA5��C�R��oh�S�m��M�DʅfM����E��Ek�WtX����P|���G^[��Z�t���G(�Zve�Hc�77s*�ɖ���R��*e)
�h�r�W.K����Pf�&Nѫ{)�� U��7��4wS��-��fb��.�[˷��C,\�=ʰ���[��$�(���cF�fRQ����(�����V�P16�c/e	����V����l:Cle��� ��V��r�S�����ۛ~Q��&��ݳ��nxղ(��s-k�V/ak�ZR@F۳F��]be�}�Mi���bˏB�k�dc�=�6��jlKsL��rm���i���4|�o/rab�ڇ.�5bٚ��9x��mZ J�Ժ�*�h�Ȳ:�WW�xsv����m%�kh�2���1�����JHe�la��CL��e��p�Oe�nb��	yjn1sE�we����r+۬$�2݆�i^��6�5N=[���	�m�@5��)��ܣjŲ�h�,y�t��1��TF�۸�4!�iH�(en�M=R��Uv��]9�2��u���5��J���{��Ԯ�fVP��L���W�����S,��ջX^f�F�z՟-j��G�д��MfE�0Fҭ��ڶ��n�V�6��d��C
A��(��lnPV�u!��/Pb��O7P��+�#mԬ-�p�/+e��A���&�7/D�3V�W�T�/r�e �;wz�r��[��5��3#�q1��gsPf�V��N���Kȝ�:h�0���pM/*B����⻲�����\�a�m��aKЮ�.Ν�r�Pav���˽����v�+�wC;e=wj�cf�ݡ�V�L�4f��NƤ�3 ͷQ���!R<t����]�ҹ&�! �!&�V@.H�Mu��ܫ�#���KR��Qe�L	4�Z	����h:,��_�5YG�)&h�0SD�Щ!	L�UՔY)��o+�60�/��
���2��8���*�)7s=w��gL����j-�uf�7��m�7R�큳l���HM�����܈j����P<w��Jܭ�b'
������$�[���.�0��8���2\��f�F�cK��H�w�S@��(;"������p�L�鱐*�R��iL;lfBp��U�69/̴\�K�R�� ��Z�*�4�e��4�&=x���qÛa5 UM�6���"�e[Fa�+L�̱�#4�Ԭ�Խ�p��I�Ĳ5��A�ۑ��j��*��P8¥�67���PA���NQl�lVY�U{o]ܡ��Y�{y�~��ZW��E��Ȗ�!uyY=�"�jmF�Z���{�{i೔�Y^�(]�r��H�+�+7/34�a�Tj�2�ɣ���.�`�l�cje�A�&9��leSOBx�x'�f,{Y�\{V���;a#a��f7����v.�`1μY�%E-���iؼǒ9�0�����p�X���+e��h;�F]`��1��&�
��m6wE�yc-�ڽ(��K��zN`^^��5q$F/u��v�u��]J��暵��Z�ٛf�^��ƚt0Ƿ����7^�Q)mJ�hNX�#��SJZ�"�*�����0KXu��=9�� ��-�$[3C���X������-a��F]���+����d�wP�QK�aٵ���{[�3��`�S��YR �5t���-IJ���[��"��Y�\0 �7B�H���ӊ�����#a.��i���,�f��B��U��"��Fnf
Çr�"�X�[Q�`ӷz�r��f���F�.�r������JL��b��=��]�
��ȢNZOE��W�L�f�yI���!
ۦI���y@�a�s-���Ҧ�SҶʌ�����Y)���[��O%ё!������$�LFe��W4�٘�'r�X��ŵ��F�Che;�v��2�G/[��
4��Ǫ���ܘ��ֺZ��z6�V;OBl��m�&f�љ��D����Q��7U��:����%m�L�m�T�t؎���*b�6��X�~謷!�ƀt`-ST@p  @�Ww�����2� ��ҤQ ���X�a��!��U�u�J����,�<�ɀV��`@������"������ ��3l�A�kP��@*��Џf�¬7�R�ac �#phK�j��ō�6�@�3��0	�z��v�'MNx�ur�3F�Wj���O�T䘺=G �=� �tz�싫u%�`�`@@.��a��ш ��r�l��,ɮ?� ~=�YY�}���:�;��4.W4(!�@��Tdd"�cZ�[j�k��Z�Qj؍�ŭ���-m�Z���b�h�QkE��UZ5�����Z���h�Ѫ���UXՊ���ڋUbѭ�X��mb�F���Ѷ�ڶ6ն,V�5��[h�ck[��"$���������cj���E�5[F�mTjض��kb��kl[[X�E�TmQUQmTm��cj�6�*�+j��X�h�[Eb��*�-���l[m���V6��������-kTZ֊ƍ��5�ص�U�mh���+F�[F�}JK�뉄O�nd\��r��������^Q�nn�Ws#P�@�#S�����}7Ã��Zp}]g��v"LLw�w���V�<CՓ}[���\M��w�*�ߔ9�w�I��e���t@|��9E��?�UQ~Ϩ�忮���b���O��EE��������|��+�o�֡_O��&�}QW��ZJ�ؕ�V��Q	oB�]o�u�9�yX�����)�<���x�g�L� �3;8��ͱ�D�gC5r8DݛS�E[�g`��a��I��M>��qo9|�G���=�u[N�Ͷ��טCʺ�nU������;M�j79��.��o*H�*�}ٝ��tc�����c:���غ�co+w�������i�m��������g���۰yկaUx!�aLTޜ΢��l�n�fS�=�y#T0��r��`l�36f�c޹����FE�kf�Y!�UY��r����RV�K����ń3Y=���ᴯ��#r_g1K�m+=u�����]����1�.�t5yv4+]�\�̰.�Z�w��yY4es�������a��CBOۻ� J���qݩ�g��TU������ �`��4�εCkp/D7�Cmc;İ��
Z���0��$��]nY��u�J[Z��;�f�غ��fc�3z�4���dx�ee�`���J+6�e�#3+���ǐ��cb����}��ևu���ګ<haV�5o��7t�� �e��9�:r��`eGԗu���+����v��(�^]��b�f�x)I>(Y�2;�oXD7k�`�2ʵG�z�L5�fw�r=�%�g�����g�hTMŜXx�qe[�f
OD�5è�[[-u�u�))y��%��z��N���i�ܷ���{�ưV��A���V"kn�kMJ]/e������r����%.F���-zyKL��[�ב�fɖ�;�N��ﮭ�� ;z��[r�=KC32ԗ�:�o�ޑ���]�ۗ[[�_GImH�ixw&�0֛W]9<�e۲�� "����B�=R�j��`b�c��.�Y�@Ӧ��/+��2��
��Qt5���/�ҧS��fxkz��ͦ��T˳�]���L��lbCփ����
G�m6�\}7��PӴf�O��))t䦙�ʳ��G���i�7�j��eu�Fe�+��y5�3H��F�;9��Cx]t�rà<��{f�N�V5�K�R���@��}��A*Uգ�D�L��5N��`w$�i'�^27�������9M�b�`���6U��9��w����&֛����Ƒ�٫x\:�V�ذ5Y���Zxmح�ެ�{*m5,椲�ǗE^G��H��m�kպ`OU�Ê5���ɚ��r���: ��}n�Ar�iS����B�����^׼�H@��5sʛOܮ��{�i��*�oa�/V��<Ƿ��ʗ_b`���ׄ+���ʧ;����QD���;{SR��hMR�u35�kzi�ᷖ��w�6�]��+L�V�q��J�oz��xŜ��7+!��K��Q���&��� ��o��ތ9iW
<���7��{cB#39P놞�2G[z�X�$Ggm���*;9�fYy�5b{K\��_R���7eҼ�4�83O[��)=��:�'����٠Pй�Q�W���Jt8��������-�l��&c�<[.���0gtح���uoU�(�7y%G�*
Jl�W{�Yw�h��Ǧ�Ȥk(�a�p�EI���Ҏ���p#�a�ّ�tf)�,�	����b�� �0]�#x��ڬV�݁eZ�ԑ[��d���(�f��kS�Sh9�h ��ow��nn��Qiw��H�v.)q`���.��n��G�%Gsc�wъՁ������Çgd�C)qk4�꣹G�����.>5ծd�B��;�:V��q=F�]Y�z̞�BWbqk^�5��r�2��/�J��Y֯��Xr�v�X������v:)�/6�oV�k��q����6���=��1����u�.}9!jg[���pqZ}�_P��HV���^E/̷ ����;|v^�$����n��@
�8�gg\��=x7�n����V�b��a��Zm������[WV���l��k̻=�u����q��x�v�L�F��]�qr}�n�D�X��T��J+��4GgR��B}�ګoe���8"�m��Yj�%�֫��ys���y̼����G��a�D�,���ۖgn��YR]��Z�vsmU�#&ǛJ��4�s��`�X�`�L[��,�a>M5-��+�R�98��Ł��(��r���<���&vu�uCo7·j�r��)�b�=��e�*�}ښ�OO�T�Yz���B�f]�[��K�i����j�����rM��lه2��7��:td�u�$3jB����l��m%�9��u�ˠו�MoZ��a��C����f>{g(:��j\��ϟ.����2u,��L�jܡeU�'�������#.i��ԟoV��[!��;�@��iқ���m��v!�cUpi=����Cwv*�-��2^N�,-x�]9�.�ͣ�ǩe��c���U��ҐE��}���2�� n#㕗XΫ�neGq<Ts�P�;.�C�&��g�՝Â����V��f��{��9���p��>���l�e:r
%�����^r�Rǝ.h��[�ܦ-��va�vtm��M��w\��[םU�䡋 ��}ؘ���]j�obV�]�/��%)�i�a�OV��t���Ff"q�ݝY�Z��D��R`��Tjͫ�MrUAx��5_ww��)��nn�.<�.��&�֗m�d��W�NvjRI��18)[-�%?	�� ^�Y��9�۸�).��ɫ��Z��Y����Jzc�:5�[��!,�Q�z���D�)+����� {u�FI�j��\���E�m6����������f����L���M�dnqS��`�k�+m���Շ+��7�|u<ݭ�e�[*��q�u2�g���}Բ������ф�[tY�pI]��q�/)��^Y���`\�٭�x�\"�ܝ��m���gf�v����Шiږk�]3��
�ݼ{[tI'9|��e���=g����^p�2֑�䥽m��|6��pe����; �pƆ�k9�9f�u�x�q��	u�\�WP� %fe	X���S��l��!�gtH��V�zn��X�f:�W{�wf=��㨻$R�-����Wy@�x�E3����R׀��!MJ�ΓV�v�i�wͻ��M�``u�fc���}��t���Yu��vV�fQۻ	�r��[�=Tq��S��{��e&i���2i���{Wc3�-a�'���;3E�X�n`�<��[<'Y�[��X@��2w>�E2y�[D7Vef ����%�B�V����5�Z<gU5WF�����÷|�	AY�*�4��;^w:��$�Y����8���ι�\<�F���˰�hwe�F�����+�4��h͗�XQ�������;j�L��S\��V*�l���Д�]í�=R��Sh���,�����X�g*T�RWq�+��H�Fɡ�n.�%�r=5x�K�(�=������1�nY��Ψ�<<�.�C/ �V+�e1�Ê�]�<o;�)�>����K͙����в{.�Ds�Óo+D��`���0�&��ێ���f �ɚf&��"*�Rl�R2��h;����Q�p���d#-N仪Ϭ�.��+o��܆-+2f1�l`W�-�]fm�i�DK�-�n2���**��W[\:��W`��Z���7ua�N����9��=[���ϴe��=ڨ�퀺�d�("�}Ie�9����_���JsV��/1֘q�	��.��a��{�E�����[F^^�	���脁�+�Q��y�S��m���ն 5�P#�x10�J��6�3���A	+(����n��+��f3J�F�)t[k�ܾ�olNw65Up��m\Vw�a��;ۭ��;���ڎ��Ӽc�2�9X��̱]d���M�D��Ri��Lr�w�<��X�77<��P�V=���k7���8�Z ���(����6`�M�HQ��1��Zw{�ݭ��8+w��Ehs:�єqW�-�L�
����͢/���G6g=J
�ﲇ.�ҷ:tc)���Ci�	]`�P��R�F��;qJ�0���hE4�W��\��� W>�%w>�s*�����0����r�;0�6�M.��a�6�V�{�־�����m��h4wVޘ�ŋ+xg��w�f+��.��k)aj%�9IM����<��\�E��N
�00iF�F�dK"�FT�֖�Z8�����Y�u������T�f�hf>H�|�Z���K��!wQk��qF٘��<��'Xfvbα|v��5�f�;�]�7��Wf�"Cj���/�)Z���'��Xܸ�	H��no�6h��z9V�FW�PLd��U!t܇"6W�N2�÷g+0���2&ʱ���Z����l���c�-�Fhצ�݇Z]��9u��./��4���H�ٽ�3s�{ t	0L�G	�ç��g��f*E���t��������P�.��Ng7get�CD�O�Z7qŮ��\���`�s��������.���2��n�#p
�_����3���,V0���=;������(X-j��%�X�wC�N����϶���ݔn�q�8Ӑoh��\yӶ�a)0�.>`!�4v�vF�v��W4�V�{�B�V�v��ܭ���eF�G�4SwVB�Ż0�b����s-(.�p�G|枸��`����[8T���7��;t��wX�ނRnQ�SۆX���oR��X9;K��jԘki��CВ14X��ʑt;���ے {�^��5�� �.�H*j�磆���fT!�xj�%z���&e\��ǽ�6e��kȨ�ܔR���}�Ý�s��
o4��jr|�'J��Z!M�j�s}��Awt��y�9:��][��*[J�_���]/��Y��16��ç&h���u��ΏBm��*A���:���(Kt3z�g6���2{2^vsde:kkupN�m)�e՞��9�~T.��r�)�h�%�[��fTP��� AkI�>�{oCeC.�&���IYD�3P�H���@��NI�$n��/n�T�Bd��/��� �[��Ơ9�L���nr��NE�\��j�n���[���[�xNj��[��f�]�stx3�t�vh#��uq�DRJ�az�ɷ���A��J;Z��m��3K� R^�3pթ��0�l�$`=����f�ki�puf�S���S���ھ:k��C�o��2�	��<VG8�ӻRgJ��쀥�W`1��t�4��W��ڶ�0��̨��ru!D�J�>��5�5V�gAҚ���{�+*��r�ј՞�w0,�m���\qӡx�6�n`��VXǷ��N./6��6��̣�;Q��w7C�y�,2�MT<�l�&����Y�Cse��9����Y���=9��שj]��b��fwh��GC�+A�ܹn3}:P~�[FY.�:�.�������U1�o �r��v̿u�WT3z�<�v��-܄��"6:�jխ'�4�ѳXs��+����>�8wf��`M����;u`��Lq�{YŰ�nY�]���π%�v�+t�e�|�2�V�
ջ�[L�4��r7ս�r(�nҼ���%Hn-�^�ɛ�s�ՇE��y�QdNa��^�r���ݥM�g�)�.�q��B�b��M�oD;���Y̝X���z��YWxmӒ��Q�D6,���m�`���/�sF�� ѝ&��9���έ廛��k�:j�f�l��U�xܺt����y���%33Q8�N(���7�7;%m�u`�3���eq���l���;c�L�1G�e�NK��0T����b�XMn�FU���z�s��}gS�]�k��F.�a9���-�ٹҷY������p�AJ��x�F5ZDHj�D�l;��wCV���8�EGo���1]���"p�ܱc�d��v��N��2�{�N=]�wV`�٘�]�ӗឰr�b�pYk��u����Ÿ"��oWf+��IŌ@/��,E�Ix�R�GS"�ۗX3�����hts���I;���!�r��V��X�K�}A{²�Y���3M�����Y1jXT@�� ä�A��x���CZ�:�������\�o�<�T�{�v���d�s_|�vgm�*�f���8q�f"e�h�����EJ��혆���^ä��OÚ^`I���Uvl�bV��z-M�#��׋մZ�J��(��=�f���g5�鍾8.�k�d��WC;y@�b�_Ibԕ�����8gN9w�[�s��gflɸ3Q�`�z���s�v���~��n\��ˌ��}�7t;��X����X<�PD0�%Z=��\Y�eI���,�2#���P:�����'v*����W<�}Kh�J�W�a>���7}x{��[�9���'3�2�/h���>\1��s6�Cj�se��h{P�tCݼIow(��\��(t�f����wn����uH�v�Ad��|t1`o�����:m���y��Ǚ��/c�5���]�' �΄��X���W�m��{GsP�4Q>M���e�r��ݏ�©T#f�O
F�6���-٭ٱ��k�<lr�{0��.l]�r=��.�{s��#E��b�7(Y|�lQ�i!S��r��d��]�؄:໗]8zu[��1�r�f�\�]9Aw�M$@$s��;0-�ݧ����󃺯L�ZS�^��,|&m�!C�@a��mn�� 3z=�玍�c2�wg3���_d�r��,+�}�Crl#�o��i�[2�D�9c��/�g5�G��d5;tv.ژv���P��������W����=%�s�ڥ�.[zQ�v��uy��^Q}J(��^�%�v���ft���������x�T���ط�й�������]�I�U��b��ѭ·^q5�|��:q�=�Z���}������~_���������� ��?7�~��~���8�8������wԙ��*Z�{-M
K���f0�ښ���yၴ�@�BF�Qv!Wf��y�䣚ml�4���Z\]�&ԃ�*X3��o�q�wk�.0�΍M��D��s�kS��a���ʹÆ�Kb�[\����YU�v̱[�96�
��T��q0lÊ�E����"+���t&����a|��"BĦ�6u�2��LYw��v�b�W���K�f�\bX�A���ٴ�/������㩭\Sb;�B�bXiT�ً�Yfes�-�&��\%�H,���^�\Q%��u٦�rьh�e��a�*f�jJ&�9�ֳ&P���a�7KԻ �)Z�u��]a4T�!H׀��ݙc�s.P�]*�
Ѩh5%�B��d��T�hF���m���,Kk.�.��Ά���{c�E3,
�j+��
*Kt6��Z͛��a��K��k��n��r�s��5�KE^m��5V�lh)[E�[<��o��нY�.��百j�Z�͜�[1kqF�M�TqVV(��1�$%[Yb�c[���!�QԚQ�h��5�*e�璒�,X���6]]�֨�ib F�t�c[+�d�"�Mb]����\��@��#e�Av	��-%��6���e�3x�%�K
v����f��T�k����2��9��bPhMS,&Z��V��2E2�c�i�+�f���2!����ׄj��i�fل��Ʒ�l���x!P���[�a��ْT���k��f�.�v�F0���F[�b�-K�4vҀ@H����/=��������#� B�vk+�J� ���($�#٤e.���ٮ�Kz�K�
%����,3mM"��ɘ�G162��c�ns��JEo ���(sv�L�s�-�S�`���c1��6&�L�AmB�fV�몬�r�m��6�4�Kh0�)(1�Dh�GF;Z�Ym�gB�lt�M�Xi�3�[4%�k�(���GXM\���	J��Eb:��ia^0X�R��J��5m�e���an"K�tYE5��m�%�n�`51 F��D��P�6��J��j�@j���ʴ[i4 3-��З�9Z6N��؀흥���.�a��6Q��i.��vҴ��^X��(p�b�#c !.(�K�K� 0�g�n&��2�9����J��v��]v�AJ̃H�Ү�e¢�[]�%,�oP\�V턶*�ՍH���ܺb(¶���M(ې��P��E�6�Me�f��+�9tKZ���c]LCJ�F�J�R��]3I �,��E&����3�m�X5��\U�7=[,J\�̹r����LUe+�9��n%b��I�����Tls�Su$R-0#q	c
�U� ��pm�6˝`*k`V��KL^�t����s��]`����c-�eq�N3�j����դ�ZeJfgj�if�դ-c.]��R�l�\���թ 1� �\�F�c5���]n�R��`�ɂ�р�0N�9�d,��P������ѩ��q���*�r�`���)��`��Yx���ȯfU�v��4fj�΁�L�֝t�akI��% ��#VŲ�n�Pn���aD.la1���e�l��Lc��&�kFSP�K.��-�l�:��FPl�p�˹�K��F��	4%�u,ne���l�Ό�@%�������ՌUL�#��m��X%r�X쀚\�@�B�Ggq��b ixe���u�Y�I�����n�	Kٱ7l소t.c
#\H����R���,(�\VX��,.,k��-B��Q��%%,Y�$e쀃�uc{Ftҡ	c���+�bU��OC��V&,ˋ��@��)1+i<!��(�`\KX�yv+Q��㊲�عvx��Qη�8khRԽT�ԍ�u�V�L�N	�X<-s���-����]
�B��p�W�(��%�܌%։B7�U��1���\�3��a曮l�Q[��l1�hʭoR�0��@�[z�[5���,u�tѕ�֨��cM�\˦�멥�f��m�KHKv���.�fȺir�KJm05.y0�е5Y��vis	\LKp8ܡÑƍ�l"�AY��a�5m��8��ݶZ͊����Ҩ�ۢF�ͻ]��&�8��5�uuؙ�ȹ���͛(�eL˞�H;m3Ї��s����ی�%Y��3W��3cTc��hl�d��4T\�E��R����
�j4Ά���M������K�t��E��<h���Z�Y�½j9�EŌ�]H�UjZ��R��X�j�Xm&�\�bSWB=�f��
m2�\:3ŞP�y �uw^�e�Fqm�����S@�̒��MB�Y�Kim+6#��*5W�]b��{ɶ([�˝�A�#�+D��Dz��]H�n�@z謚av�I��0�������F�[�vP��P-1fUq�����-�X;R1�x��	@�aq���t`ؔ�k�h2k�[rX��]R�M������B6�Q�+W@���NRd����eю�ĳV��P��]u$c���kڹ��&�a�Hb���1��K�4�4��[�a�u�q��G�(�J�]���Ԛ���SY�X+j]J�rkV3J��޷J����ɉiũ��h�j�F$��
�պ�s`�n� �����b�[�c(]
涮Z�K1	ct��cZ�5�˲P��KHn�uD6�W�8eL�L��\[iR��#�W�(��鶬y6�j`���v�\R�&e,�V�5�a�jJ�g`"(ƒ�P�e�9�e��sYf��]�k�(gb �`��W�����n�b��PњڮF�d��f��,uv��u��Ք��õq(�k�̶e5�Ҕ��u�"!A���fֶ��i� ��2*KE�eqM.���$�M��7T@�vE*[J���(ؠF�&%�K\�	��X˳��1G�lb�:�-��d�@�6�	f�s�YZ��]v���f��mY#K�۳X��Mi�L��u6L�<�U�!K�8�U`�.Z&��Sy�ճ�,6�`L큚��j��5��Vd�3L��b�H�AR�1-��2�m����c�Ͳ�VZ�#��L����j��ųD\�H�`j�L6l]E�*�s�e5Q.�����JWlͪ9kV���e�En��n����Qـ�&�n�y�6l��Y\M���Ę��馶�=FU�0�hv���n��5%4�.��,*�a��T��aj�&QK���THŇ��&�eJ8�ctG�qXABSKF��h��[J�Lcn��&w�G���BV��5eh�ڦ��l������"F���u�"���.F��Ʊ��bm(��d�v[��a�J��F�3X�3TphJ8{j�Ee�+�u]U��+�̰1ԇ:���&�%s���lY��h(�Ie��9V8&)�Ԥ&�;,+�m���P��� ],��Z��X�R%�KFi��.�&k����������)�-֠�l����).&ej2nмV�v�1��c��MSM�JV�]��-�Ss�4�aC8	��Y��l��9h6��(9��f��d�	r�1�5������$%6FL0��2�^܄1���0��3mδ{F���]�`�\m"d�Y�WCWL�p(�b��k����k���YW8�Y�9㮌&+.�N8�n���3]\��2;F9 �CP�!�Xfن�i��a�CF6�h��#�b�']Bh����tX��R6�U�"�8�%��h])�p͵f6ۚ��\j��bkP#�
H���*���	�43-d�KB��C�vZ��)�B�[ŻP��q��2�ʦm�V��z��d�b�^��JYʡi�TZ\8�ڎ�âa	JV4�)��:�k�@+pjM�Q4���ZL�Iw3b�f�L�2���9���j6�Ѝ��kx��icY��9�]R.�-�ZJ�>e��[�8�4"�)��ģ������/g���-*�ZȔ"j]R9Mb;2,6�MP�ֹ�����]� ��qu&��#WV�YG�ah�&ΫWn�4�f5(��(�X�(2Īݦ�\P�[6�2��1e��LlZa��	�̴ji�D���5���L�גka��%lʻj��
f]����\�qn�l!.�yk4�d��M�]Z�ф[&�"J�W���X�ͅ�����)]��Fm�:��Y�,6��	U+b.���P�kK)��YL0�SQ��]�Fecٴ��`	KX8�Mx�.�Q6	��f�ZhF&��V�#��j���UD�f�..���J�!nw<��CX�l���%N�&����ڱ���13j���%��th���ɥ�cF2���6ƚaЎ��&��p\ԳH�(jV憛)l�K��q��;G`�(B��%�
d�f�%tYH:k�2:�)�j�z�ѭ��I��i���Jʃ�N�\LEƴ���e��J2ؤ�%1�Z�]u#i��b�Ѩ��D��]�M��
�$o��Y�4�Al��f2ᆁ�G��g��m�17X�-����n����-��֑�1��	�}i<.�[^X�vr�f��*�TװĚ�v� f��llE� ;L/Vhn5�K�rÁ*iR/l�2m�V4Ҵ����n���uŚ:��M%�.�Uv�$ �j�����Fgb����H�s�mu�.,t ��Dl�iCM4Lp��%J4�c�ɥt�q)�ʃ]y��MWL�sn�	v����54���#e!u5H#-�k�5�,�&�Y��|e]��qq�GK+c�u�b[B4�v6e�L������2�V�5�ɩl&�WD�y�<��lV�l0.A�6l�cv\Z��.JZAX�l�!H��isY�m�٭�����
�seVܚ�ƎsXU��U���e�L�Վ��j�UU+�
��daX
�����9CUT[n�,�as4�֪L��̥�d�=]el��@ŮC6^� [ָ�X�l#����Ņ���ST.��K�&�T�t��֎�����B�&C*4�V�Te�g:N �	�1a0V6)&b�)ch1_;�R�����&4�QX��rɋm&�>�sQ�4*LTc%3DT�QF0��Rb�)�EA��F�IEb���ym��cF�h�(Lm��+4mQ�E`0+�(�1c\�Zƍb�cX�mTc`KE��l	lb��j5����6�I�E`5E����mk$�chѰ�$d�5�,�i"��A���y]6�����p�5h-�X ��A�$ �֯%�j�W.��	C�*+b6]�.W$�^ne;2�ipf�],�f�6Z˙�V��G`�Q2mT�D�e��-4׋�ٚ���"S�v#(�%#�ֲ�j�:��%l`]A�61ti��5BkMM�U;k���ْS�K��E����L�P"Ūfһu�فHlPY��G�3bї�SR�����ٚ���%�0������%�l�h�j��3i���)Ʀ��	���X�Ac6~]|�<6�71��l���GZ�-�J�&�J�H]��*��`�M���%�q��sI���P���%k@f�ך�n�\��k/�v�#�]�`�� V�@	��G����6#)�.f��������Xkl��Ў���Bg�5a�.���IlR�&���T�e�
��ٛ�ؚ�ؑchgP7��4�\��ZmX�B�c�.J6���R��^�Â�:kPV�7��R�&H][�I�m�h�;E��)�5�S4Y67r�WJMf�Yk�������G�ì�	LIfc��]��U֛D���v��1d�nU\FbB*��RJ��LZ�F�4���	kuSmZ�sr�ST4-�+��2���뵴,2]3u�@6��˧��M/,]�cqt���H�¹��b��ԋl��Q6�m±0\���u�Pl$)�L��7KPYr��\�%��뭎b�%Ɗh��G5��JSG��	v�m(ڌ����Ts�`U�ʁ,�2�{"��XV �&u��+��LlM�,��e���ڵ%)[v��[�Q�XT������q����D�`f����)I[�1�`q�`v�	6�R��U�Ԙ`��ܕ�8&���\0����̔s�I�WK,%���Yx��YM�¶���a�k-�(A��[�RJ��B�p�R���i�W#X��K�MT̴Yn�"�Z�2͠@͛MR��j���4��Ѷ��.is������j�i��À�모T�F[]PԀ�ǇI�#WT�U*�$�I(�`S���o-��J��e%��ڕ6V��XK`��V���2�b2��Q:��QF�9�VR�
�V��m������Fڰ(�l�j1�(F0,� F�b2���^�P�J�!F�ai�� Jij�oZ�J�X#E���e�'���XXhSY��@.�f�4��:�j#�-�s�&���`�eF��*���$>>��y�-�v1Y��gW7Vr��Y�%�4��G�$qvȤ�o���h�F��xV�f���uu�a��{e�k]�Øz�}����$,�&mwj�Ff)F�������ڑ���ｨz��d�*��>��~ɟoU}��zk�O��wǸ�_>���nf#��3�L�PU��}���-qww������'۴��ƻ:��l�/�����J���喇ޑϺ��Y�f���#�a�]��t:�n�E3b����V�Me�U�L4��4�^K��w���Եf띈���ͫ���8�l�\^�_�jA��ԋׇx����d�$��֙����^�.�ɱj�?M�\�v`��p�svJ��"�6��<=ڴ�����R*ޱ8Dw-W��$�������ע�PK�$Wݧ��%">��R��OfHWA�!�{�^�6S69��Տ霜\�����g6.��.��^�u���D\mS+o]ܚW��"1D�$�3T�HɫkgNQMuwϓ�ޒ)VzA����v���S���f�n��&4Q��˺���z�m�QA����h;��9T.��� S!�D�Jf���.�J�*:��,�K�j|��1�ׯ��o]�aO!^�lT-�cC$�Y0B٭!Nof��w_�wp.��#������40R���z�r��7Dk䨨�K34)`3m� �On<@��2����}���LCB�}�]Mc�V�itѦ_C�%�[ d�w�x��qEi�S��huwK¯�ὝC'[+_QJ��(�S�����S�mؘF]��m"�פ��k��w���׵�~��j�T��*3m�:���X�]��T��͝��Z�X��}�{��ϫV���ҺWp�I�'�2��	.���{Y�#%C��Y��%��wH������NF��dVY���@&��B�W#c[�gh$�ť�u�J�JR:A��_��g{�Owo��J+5�a��U�Ī�f t(:4N�>/w*2H� u��<5���O�I�
�[��P���ǖ[�Z�v�v`����r��t��I�TjJnm�W�ukP;�*"��ff���ek������ǯ�f�A�9
��p�z���Kk_Jim�%��/Un޻�=���|���lǬ�wb"J�Bʃn�TƲ�)G�����;b3�w�7�Ҿ�5q��L%�%f`l^Lk�7��)��o�I�} ���J`�����P��t�߷Wg��o�_!^��T�f�����}v�O�_D	�yo7҅v�*`mv��V��˱q]M��f�˻"�_g���U 񐮊�4h[R�&�bv)�,��-07)��z���%o�u+�0f*={�?�zn��/��Y��g|6���o]ʶVde�}\�k���W����� ���,����Ȣ� F�j��-���m����v��T�����)�U���5���$��E;���4)��̽�N;SJ�:�-��P%=$5RT����]�K��:���%;��$��)fR��k����v�Y�uH�1;���r�Ʌ��&/xB�Awf}��Z�ȴ�)�DCI|KJ@�5դ��;��"��Ύ���%�UM�j�]�oj��b�����(U�E�M�r�M��[xfy.���ge���b,��P�v`i�U�j��w�p�8U6Ps�Sk��&o*��f����[b�X�cu��6�9�d�z��:lefz�	J�l��pR���B��g�(�E5�k�G0���ejh�h�D�E`љ,3J�niD.�\�W@٭5��1ȹ;h�������R�VU|��C�O�Bk���vr%��! 2L亴\ia3���,{P}���V`d���+�>�Iu����;��p��C�`W��ԅ��0����v�~`m�
#s&��<ޙ
5lm�fh�����'+7ލ`k���
׊��.w��q*�<���H*HjG�g�þ����er�v���/�禾�A$5 ���1�{j6 ݷ��.L½�;�x�x�~�χ�}�*a����R
�T����ފ���'>k{﫷��u�8��_!��R
�g��?���tC���HQ&�;jKs���[41+[5"�r���uf�ͺ��2�-�:�$���R�Q��hͶfR��lZ6v��x�����ݽ�wb�ݙG���N�?a��W\�b&��3/#7:v®5t�tOA�G��γ��[� �k�wXyד̱د����� ��c�2�{�v)���;�>pVA��u$��T�2I�$�u�,���I:p��e�ŀ�ʚ�9+F�*ۊ�ARC�e6H��+wMH��}�M��(7��K�W�g+%��g�+ ��޻`.����n�cf�	��à\0�%��rν��d��o��=�ͯ$��5��K7���}��5!�J�@��b���Slt� �`�bd݌�-��Vf��ܞ߽޾_~��{�<J�sp��&]RÐ��!���k���5�I�AY�c��}ڎ:n�d>��9�;��lgԠ���g������+�V_ۜj��Ԡ�h�I��IU�r��#\r%����g�A�N�o�d4�7�.l�-}�n�h�t�������K Ydl*n���&nX�9)�LYvVRB��%owwK���T?x�>5[�ER
�{sg׮#]���u�[x]ہ:���Q��
��_f��9���r���墜>^IJM���ً�I�-ƵJ`�ks3���F�V\F���m��o]ަ�;1B"�>�׭�v>K��
(0e�B��kF�	�/],66�� U�
5�X�`��Ԃ�AF����K�pM�_pa���s���υ'T�g��#e4�1^3r�
V��Vj:�&RÏz�zs ]��1(zXP�D�T#��>H$�J쿣���?l��o:�˷3�W���<�H*����w�+v�$��Mo��zj#׌��Vm�P�kƦ���o8�5�+6����c�;�yN��%EA]��ѾV�9V�iq��6��n��rA�,������nڬ��8o@�� ���M��/�wg�wo�]�Zx���tP��6v��W,­n��Ͻ�V�>�T��=��Ͽ{OF����-e�B�f���:�bss0����#�	�4+*�Qʠn���*p�!��Nﻬ��3�=�Tɡ�8�Q���`RT����/����ͧ��G�Y�ض��egBƖ���
X�-z��� �6Қ�"퀻k��Q�Lf2�i4jX�𣏕­v�����*���OI���֬�<��)͒O�o�Z8&��v-��l���p�z�Q��2
�E�R
2�>ͼ��d68. ��qUuQ�	�6)�@�oe�����!�r"(d�;��S�Up��X)g>	�r���:bs�8.gX�]ܻ�&�h�у�?�qV����6�_DI�w�AfjZ�}dՅ[�߷߽��v}���[�BW�X�ئ(�W�k 5�R&e�Ճ@�3��1�M"��M˛�+	�i,B\Ē��q�7-,	u�F
e�����%�֖P�/2��"W�5�4�6m��!�� �Q%WKK����P�WM^:�5�6
Ave6e��A���ƾ`HZ�hFP*�SM+nL��S1�ۉ���$C��t�UWEx��J
ʯ�O����"|�eH�8�j�Z�WP���x٦���Cb*%9d�tHYVZ�E|^ɞ�7�e���xy3�(�yN�'{uM��,���^�zI%��Jg��k�Nu��up�]ov-ꤷ�'��Z�>�����}[�us��xR�E�}H<�ٿQz�[)Ox��V�l��,IP�WpU<d�q���7���zH[�/����y��o_n}�K�]��0�W���A��I$���np�]��=�,�k��u��NK��>�I��f��yIw'<>��<��+̸���-c��z��tլp����PpJ]�D��H�����i��d� ��]!{�-j��Sa3[��4=��-��
�
�>���{u?��M��[����\����k�]$d'��Ȯg�i[334��0�N�ںH�h)���T����$T�v�X�dR���s�`�]��I�X����.r�p엃3�(�2X�]�n'v��x�p16�'I8I]�ª��c��U��v�o&��rr_{T>|*A�!����A$��ӍT��z���O���O���'�_!O
$�o~t~�#+��=���zAU$2
������PS��~�}u�H�;�v}�B����*����y�����_~����v�tM�X۵d�h4�e׬��L&�l^&`P�}}���>����@�-�֔ݚw�9U���k-��̮�w�]�h��ܒ*�o-})Ӝi�	L�ʤ���j���M�-��zIZ���̂���VG���}��ԝ�{v��O;v�۷n8��x���y�ֺs��W���~���cm�{V�C��{nf/8��y&�"lǱ���5v�k�cU�(��q&+���YVr�'������W,��:�7YwE��	�//*u\TZ@+�u���N����v��tv�Vѣ����홡ɝ6��Z��h,Jt�.<I�W�gS�]�Y���qWeJ e�fȹ<��wq��l��9�nh�6����W��7Q۬=u���"�ҳ$~��7K�M�u�B��=Z0S7���˶o
�Ʉ���Fм�왡�;��e�c��뒈\��f����Pd�N p�^ڿ��p鈭+�m�]�-魻�9\nκʤMy�w+8���w�:s�_LuhT`�n�.^
⩖m%|�E�m
� �:{�l)cE4��L�:�o[�T<�u3��ꬻ�\��j�۾���Φ�������4��t]e�_+!�tR���NS-z�:�LәN��8��,]��.�wWXjP��OI�����r�6���u-\��N���P^�z܆�m�7��먬V�����ز)����l�B��nR�ӄՊM�l�љ��]�]	՜m>��9V�mV��pZ#Q]-M�ּͭ��\s]���+(\�1lҸ�B�Xf����W�Q�]ыyR2�)�P�q��K�d���ϗ)��b3g�[Y{�{Qt�X��5t����&JMm�V�4��J��)�-����ܕiUC�g�f��D|��]Y�u`'����ح�yǀ��*p'���� {�r���`�dT=c���QsBR�`�@��k���ʠ��z����1�Rn�{"0G�G����F1B����md3"*$�ة1�j
660i ���I����IE��&�A�r����J#EF�&��E��F5���E�(I4k2�.n�,bѪM��FB���1h�(���H�(+��5sl��\�����7���*(��h�,Tr�v�[�h�\�D�v���7*�scGN�u4L��]݈��E�w3��n��"ƻ��>u��.�չ�C��@�wv�{$�������&�.���L)|6wv&��A�JX%+r�!�+��wW���#b�ۥ�7-Μ�p'��$sP��ַ�Ye���幾<=:���cC1`���?���	-�њ%�ĥ�4{c�����#o A	3��p�$�@�a��T�ONv����S����
L%���:y�aWU��ۏ��x͌=��rs���g>�Oy&^0Y0r�fd����7��)va�Z������jn��>�8����pT#Ĥ�
�3!�q���e؀�8"�`�����%�BZ�*����lH6䈚����0�l̿o��'}�� ��7�i>I<+��O�j%,9�}��h�{�}�T��A��kz�p�$�@!&p|櫷�A���oxI�='���:����Rz��N�Fx�nޏk��9�I�-0�dF��}|>�k�u�?�>I@��:O�F�=����<�Y�jn�J|=�Q��9��p�BQ%&@I��Y����F�㷺^H>8��� �RO^vd.�ܼJXs����;L� 3Y�>#)������*)�-Mr�bx�GZ�飤&h���dh�L�JPo��ԯ,,�9w�ma(CW��O� �\�;�m�-s짜�j'��S�"��A	(�HI�r
N���L#�����s
O����
n%,��HI���g�Id̫!&e��\���Vy�^�$�Pټ�QW��sE��&G7��U��]Mi�h�s�����z�9Z��&�=dU��cqw�V@�J��z|c�s^�@>s�>�L�8 ��x>�Z��g�fg��Y�J���w���Kw�;��SJ��7���j{c�i`fNN��E�9$��	(��x+��r��C�~�z�������*�ηn �+�0k�Rg��I��'��L�Z덷�0��;����/z/y�qt�8r{��]?%�7�����.���o;�&*w�8	�b=���M �
I��9�,���pZz�Dw`�)y�jYp���Ks��fz�?�3�JD�)��'�^�f���q�ղ�A����M��wD^j��nݭks9��?������|�ۙP'��<Qq�x7P��$N�pk�+t[E�Ұ?{��W^z�G��n>��7kK�"���UL�bb�X�b�Mjk�r��`ia��P��Cî����Ae��m�9�r���Q-)Zl�],��4#�u�1�ԯ9L�E!o^p1`uִ�0�E��!�a6b;U
�'SPѨj�QVX�p��(Z�"�Cf<�E�Wgh���������	qar��m,�F������Z-e�\��%��m���Z���\b�Q��h�x�P�l\b�L��a�@�����z���0������0rQ$�>Fg(�~&2%Ngn�|"��'�Eqhlm���s7�@ ����0pR`�>������m�F�{1�$]FV��/WM|��ztGS95�I?��0k�A1g���x9�g �i���Ra^�4��)����*r���Vb����RÝ����j ��9�IDxC��i%�Q�5�'�����"dfr��1Ä�D���-��
�q�w̻����O�E��pA=���|N��� ����{��Յ��K��Ӻ���U����4|�k�!%���V*�ڝ$��W�be>�XHR���9�bE6Ԃ�s�s��r���K5��g}�a��^x�&ϒOy�k+y�)�a�`�-[Y�2i]*m� �+�T�GK��p��� �Q��)��Rc���Ȩ�0�U�z���9D6�lW�)�x���;&�)֝E����}��
�Uy�V�ù���ˤew�ʕ���l!�F{������G���l,�����eD���v�A^�}m���I��Ӗ��t�!@���"M�wZ�`
uQE��?�ZŇvLpq�;5���(]U��gN84\���J#Ȣo�1��R������q8��'�m���}փ�NV<���d�1ea�,���pn�|�zš���R��w�4\��I@�@(�� �'I?�-em{��9��F坒b�C�����)k� �z��)3�$��熗7/����0>��@g0DZ������R�p�\��
��tZ­qqUҥ�O'����,�n�&�Iç��9��B��w�w\x~!2�Z�1z7�1���R`���)'���WQ��M=Ac�����|-�c��幝C�:gV�����8�8�BL�&,�`�p���ycQ'IDx��xW��h����6��cQ`LR{����/���n�6���G��l_��۝���L�s��b绲�كjl�\��A�����ڦ��<z�qlvY�"�4��N�	ּM�)3�A)'��o� ��8k�o� -j�8���9y��Ԯ�87�u���g� 	�;�r�'c�^�0/;n �w�9I�@)'����I����R�����,�K�Ū�gP�N�BY���aǥ�qz��z�V�]ry,d9$0d\��+t�i6�{�R�ft-3B��sI�0-�c"2��A�'BI�)7���Q�/�ܶ��Y�;q���Z�y�jb��ȇ�gRO�&r	I���r��c;\C4�^�x��� �p�'���y��Ů�;���.E�!$�骭��2�_�sq�[I��Bd|��A)'�>��ئ�u��IR���H�.�BY���vy���!n@�p�r
N_�&Q��9!8��q0�N`�M?��{�!2!�r�S��K܎��;���okd�&�r�%s:p5�ƠMj��*��vpY��}���]
2���/��p��1�a����c9�>w�o�(.^���.�P�I���>��χ�;M�=�<�v�8>%EjUB]	�K��1G�ջZ�#��@&y���ÂQI��.���6D��
���+Fljƶ��Y��e��H�vH蘌�Z��!���j�r�����o ���)3��JI��7-,�%�D+�n���SE�_0��4���z�<Roy�NJ��R`��f36�SoI�F$@��e(�N;řg)���q#D<���n��>:����R`2�C��Cs�m�������y��rS��
[����cu���':,z��Z0���G�;L�����I�I�fg2�Mr�WQ.���ێM$�x�ܴ�dt���1�������s��V�c�'��tW�Zo"� �QpA�N���m��R�8������}��=��1p�"afv;q�x�[i
M�)'�=t�:$�׶�s�x�b���4�������l�+�ɷ)ǋ���J7����~�"5:��9���6��A\MʢU�=�xt��~S��_�́�(xi���˫e�ŔWf֕�vv�a�H��\6�%ڈ�q��ST��3�0����Wl��v�B\B�R9���6��ؓ6�9���e�q�����ƅ*[v06�Ze�Mі-2���1��.˭`�ڔ1�u��;��Q1���尛k��ic�-kԨ��f��6@�����I74l�B�kR�]4���*�����?x��*�[cf7W'%��3��7k(�]�a�2������& 4�OW��å��9�I8�QE�)8�zI�8���\0�����+H7;�Yu)4A����Ra�A���1�������XW�Sy�k�ӗy�:MèW�7�w�S �PL�Nn��N��������#�����-1�P#�T��N�R���k5D�󼦮��\7�9���>k x ����H>���w�g��=8Ӕ�3����>հ#�n�!'o��h=7/L�a�3�#i��=�QcW�`�g�z�!!�ٍ^2Ro9���`�ϒ`'��#��tH��U�����m=)�9ި����Fb�Zg �'��]�U����كǌ;��\3��0KY��a�@�]��&k�е�,f�%�a������g���{�`�$�zI����=��0��eUfv;q��'��sm:���>V���gRO�;�R`��y��itӌL �-��Hc�=���Y(��0�k���F_j�o[:T�6�>��cpO=�k�8���]��;�����ګX�<�T��YYY�E�ǀ����Ea����8O���O�m4W=�u�@'M �k�i?�`���qQ~C��3��^?�7��䚁�$�d����ئ*�T�i��!�$�y�=L��E��8����\7m���WA� ��G2���dC�]�{��a�U5�����]�y�����Ầ�1[8 ����#ɔ0 ��Ȥ�AE#g��6hs������<_c�9;t�\q������OV�rQ��(�3�3�뇬����Ϩ%��U!�Y��]Q�F6�,���:�7mIZ�D륁���M���bS��O���W����j�k�)(���LsxK��j<Z�eʷaD�ӆ�!'���#Ȣ�
��䤓�o���B���	��K�����
��f�7�N]�,�R`1eld�4C[a�<�_ä9��8IG�F�#=�<}�-��gX���j;�U�msW���W�m�}WR�A`���� r��V��_�4����Cm�K�C7V!pՑ/J.�,�J�&�3�����w��F?pqS���6>���:h����ITx�ȇ�I��e1-\����O�"�gI�z�/XoIV��,f�1��=L7:r'lH2t� �pBI�x��BN$�S)�	�j��f����yg�B����op9v�A�����$�v\(m�#��̰o;�။��V]��]4ȡ��nul�V��\K��0A��Za0w����������O�Eu�s|θG�|��8�3��9�K�V�<S#�H ��<|9��5Z�Vf������}x�={�il�*�\��&9� �8 ��� 4�U�3s�8�b�����t����IDx�2>1�0EʮJ�ϻϹYs�e�B�
f�;��r���Hr�9��E;xVX�Аu|�<Frq<p�$���O�\Eu�s|κ=���^>�Uqײ\]��r��'�=1�zvK0�O��{��\��k?��xmv����^i�S&`����b�Ys�63ΠY�fV!��62�x  ��l>g�����ϒOȇ)0�.{��b*Wx�j��no$�N�2�Xo8I��{���
��"�o��bm�0��AeTy˔�b
@p�L�5tY�\iHR �.�6ͬ��5����Chy�2r��A���%^���t�:{��p]L�gc�	{��Az⻝��2!�s��A)'�Cy2��8�7�O:��/UV,���|���O�\Ew]�|��3�	�`����$�{��w����8+�� ��C/��W�7�۱�������N8&~��EL����*{+�+W��	f��`��i��|��!% G��j�5L��0@�ۇ!^���*��-�S�	���v���y6P�a3�`V��A�O$�r� �(��hl���=�G �Íx���."��ܾcw��z;L�f�pBJ4�{�a#ۧ�on�<v��۷nݻ}w��<�Iŏ���*�Aw���M'�&r�����_\V8l���ٖa|{�$VJK8�Z�0�>�9]=Y�Y��<�j�n��cV>^�G�Z�)��\��hX:Al#�s`��_�%������c�"��H�PEm�*�Otܦ2aڜ6�j�s��w4H{�o#/�Z�s5�]C����'!T>���A�?EִAL��]��_J7D��jJLB��f��[�+�b��@�{{7��<j��7n������<y��I����oF��b�b9�v�Tݘ�gB��-",s�0�w+@7��5y��壮�ω�2Z�Ŭ�L�����u�̢�{.�h�yZ����,�k{��<�*��^��غ�ll��kg,����m�Sљ��·&f�Wyܬ٫���po	��MW�4u�7���hP�̚�w9�#V�I/d�l�L�3&�F�.\��\n��}w�q�XE��oe ��B��8h�ż����wL�ko�����mZ��;�C�{\xnA7�����4�,�A-k�yF�cgU5�)h��͓�k*{{������>����cqo<F:L�Dnɺ�W�׌%����Hm��(���NA�1捔����Vl�T�\�3�M�Q�r���E�yO:����9���Yc��f3ɓ�lMF+�k�A�&�[P�fK�S��wҥ�۩�k\�Ё�k�m���V�C(]p5"�e�m+kr�kӖ'S���P rhө����܇+_]���Լ�`�,Q��q�L���IU�-���@���v�!�7�(�D1r4�����Ad��l�Z껙;�nE���JjA���7�ך�����\�5r�M��W�|m|Q�ѱ�v�|�W�F�.Uʹgw6�A\܂�e��l%$�ە���y�j5��ص&lXڊ64VM4X�t�E����\�s׻���k�����l!b+Ϗ5&�����v�w\�{���E�7��Dky;�E�%���Ts�s\SE�w����͸h+�{�:V���5�k�T�U���ڋo9a�%���#r��2X�F4{��.s\�墈�����Ũ�#EW.o�u�cQ$'P� �V�KQ�A4�]Q�ܻ�9�6�3s��=]�Bcj���V:ؠ�M1t��3Y��mu��m�Hb���-:�8�JGV�V�������|-���2Y�Cm��[� G2��D��W@�	�K��9�`��"�\P�u�β�[u
$�� ��L��[˅���[��pc;dU%a]\�86҈[�˥��K�.�^w[�X<��N�#]�fs1P��:³bWl�#Q��kb5j⨚:P�k���b�;K<��_���l�5�%��2L��u�uuXf�yZ�[��iQ\gB7�k.�+ �R0oWiSif�4lc1����n���^���B�eqv���YtZ�p�Y�IK4 %ڋ��¶�L6gR5��LT` ��,!)f.�L魰��D�8�t��V��BMx��Bb��Z�T�p�,"Gm�UlJ!t*/�d��gK�]2��l`�8�#�)���D)*��Ό�J�݂�]͍Hj�j]1�b7f�Y�i�y��iEv��m-4(a�GdB�nIFSB&��5�b�\j���3�T����:gW.��T����Z��Q�m���v�m�6 ����@.cJV�!6TƖ�7qs������4�ͳh��u�!Q`�slA�L��Y`9:�6�قk�)�u�s��HʳM��4�t�V,0Tv)e��é��/�d�,�B��դ�/��wVS`a�q��mE�f"�����ٸwy���e��c�6��#�]cɳv��l��1�aa�1�7e���Ѵ�B�2� �m]�l�i��2��g/Q�%v��K��ȩ)�,f�n��Ť`�3^�Ij�CB���6h͛1�B���R� ��P��q�,�V��+H�L7m�^�m(`����(�!<��w���+t%������$Y����E���jғ9�J�!��Û�M���p@�����H;.�H��8�%����X[U*ݤ�p�1��Mrd2��va�)�s�&�GZM�UvQ��Z���빅MhYD��w�j��)�"��=���
����,SQ�@MkH�6J6�T^]ɚԌ�κ�j-���M�Vӛz�0JC&X�ok��Kt4+؃��H�k�/Z��ە���ޕ��FĊ��+�6i�\���%�E��n7!`d��q��нm�K��%X�S����MH8]���q,7�.�44A��u����s lȣ[��y.�66ʎ`A�z�=�nS2��aHK�]1ߵ��a��cv���qjҍ2�"6�.��]���F��l�~� �����I�	I<^vY��ԩ]��-��Y;�����P���d7�Rp����f0ɱnD
Lk"��W��i����%]��e�J{�Y����[o �/�3*��ve��I���|R`� ��&A	8��c�x��cK��V����Fcw�� ��9�J���8	4�\�;/�ʥ]���u���p>)'�}�*�:O]J��7�(�Ǔ*x����`�E���ITQE�)8���R�*���B��ў4t���[�*_�2�U���L����&p|�~�M�\"XñzM�햳�D\�K���g�Tl%٦z]F0���ct��v�3y١�3����cr�/�\QE8I��:�M�^��ώ%��+��.6}^�p���l!�Ro8)'�C��7�*[N���k٤��V啱 �6u������Fol�Û�K�D������RKwAV�a�c�o�Z"��(B�MK�x  �����3��Aϵ���{�	멥8eg5�	����N ����������.��t�pAIÐ��#Ȣ's7R��m�Cy����T��J��V.N�A3��xϓ9�M>>I<N<´ƒb�{n4���
N���n�h���?y�x@'M�Wi�eF��v�.�ǎ7���O�'���]d��N]��`޵�<��4�Щ�A��ט6�� ���AI�lh���v�7x5����� ��g�3p�9v�qvB qE��D���iu�D(h�1���'Ͽ���G!s$�G�o'Uۜ*_��z��n!U�>޼!�`)�} �?��3�	I?�j��Z`��ݶ����>vށ)�O�����c����� ?�>�p�$��@��yL����Q�7ƹ�@;��AL��i ��z��uԶɹ5�v�;�B/&0�iU>��KZÐS��
�]�L0�ݶ�0Z�<M��6�Y�@�ʳ�j�����vm�6>�m�z���3Y��c'T��cJς7�y0r�!&rI����@�;���LeJ>�p�V�������-:z��]n��;o �y�0A�����	:�/Ds(�����e{]��בҐ�E8q�3����;��!�?y�zd1��f��>�%&��L�������H{�Xqv�ZCE��5�h�e�\j��B3A����gWLG?M�&�����
3c�\�d���)���rE��@�x�pBLJ�Ȣ��J���6یFտ��+�ܸKI�=|N.�n>���|���)5
����B3t7�:xq��
�BI��4A	8�ۭ��{[>�~��ǈM�-�ϯ�2}�f�rQ���dC��8"�)�aݚv�˯F�>���Ow7�B͎|hY�9�,�0 ��r���A�ju�3����R���w�ύ�ʍչ���4�����2f��ύ��v�$��������
uү%�j�_����[��PC�*�{�h��E�����E:ND��Ψɗ������߷��w�)�u�q��x"��&�&O;���R�[6+�����5%��VUEn��Ҏ�J;�Ձ���\\�݈08Q�	�`����G�(��)8t�mds�t=?Y���;�F mc������DK�㷦<Bj!�I�|RO �w���wg=��x��h �w����l7a��YY�����LF� ��=�]܅8ͭ|��-���O�`J<S":p��O�h�܎+a�A�5y�0��n���pRg ��v��(�!6ʷzE�ʬ�`"' AӅ��8�7K�^c��넬~���^��oCd<�99R˙�����Dx�j!�L��x �Q
M��Oo�9�4��V�n�[�;ff*�o�����jP Q�I���^an�u��Р��7D<�=��j���u�2Ch��X��3p�&\�ϫ���+N��"�t��3b�	jki�Ob�1�������t�����y���e5�=���W��m�Z��eѦ2�%ڴ5%rl�i(b�ȁH�Ԯ��k���iMv)Q�c��Ze�]R@0:d��2��md��b�k55P49�g&����֚�ք�˱�2T�K u4/$����6*4-#ԛ9�MA\�1�f\d0��f����MfV�V�-9�)n���֢hX�man�̺y�Jp??>|���&Ѓ�R�X�$J^�]3�3�(q)�h����ZMX���K�������G٠�$�<|����'����L��N�E_[sޖ����X�F�!�{Y�A$�B(�)0r1�=��Ȁ���Ȣ��j�<lCt�
����ў,t�pFk��UI�'�]�mf����Si=�"<�I�$��t�	����bh�Ɯ̅���[ ��@�QE�)8rP GE^z�q%ԝ.B�n�x�ȎY:{*7��m��6e�����1�'������`�wq��pR`��I��%�u�w4V��"v��#�������hށ�:l�#5���̈�L�6�~�2\N\�``�`a��z�.�M�a�mX��\�u�K��8f3)s���o�ޞ#�4� ��I�3wx�n�vcV,���Ree���1��(vz�����9	(����"�}�o�:����i�t�`w+�NΔ��ť܆U�x�e����e]��<&
<�-�j����=]��&7v�0�H�y	�|""��>w���y\����3ߏz���8R�Έnwu�x�`6�)1��8Ӥ��fP�ESwXҁ(����8.m�^1���N��W��6�_xG��p�X��IDyC�1�r�W�&*PZ��SY��O� �������\�������pg�"Y"ϒ�[l������	(�|BL�!&BJ���X�Q=���P��y�F�6tCp ��^�񃂓8 ����-����a�Eߡ$�☼wp�ۄ�+p�a(��*��R���k�3���&v�9^,�M@����UL�eۄM_+l=�}�t��sP-��6}<�gk��RgRO\H�s�f�0���~7��d�o�{��������z�9jP#�$�o4�d��`y����0Jg ���!$�$�<|���v�D�;bޔ9�{���,Y�)�BLɥ�vd6�ʚs�kކx��Ϛ�-�j�)]���d�TA��X����]k`��ٚ���vMj���w�fp�|�����;|�u�g͉�,�m'����.��yleN��4v���BL��[�F"&��1���:����*�KK�̉s��W�
��lƂ	�ǂ�c ��#kc�j��t,�xs�͚�m�-F��>���F��<I����D�6w��[�dap�Ę��g#C��(������
Y����ÍI��̤�8I���>��@$^����_@r��R`�k(v�4�~pj(fe�xn"y�"�z{��hh7��gi< |�� ����vqP��,��F�J��gu<DO%9�;�X㈜g� �8rU���A�x�������o�ާ�AI��x�o8)'<��*�mx�	�G_3�6�ˌ*�����{� �+Q�Q�|IÂN"\U,��C�7��p�_tG�dCځ�ݽ��MT�̟s�{��<x>�r7�sk�w�Dx�w�X���F��)�=���T)�O(�׮�ܽ���V���9�6v�tS�[uĢb/]HO
�*��?U�w���\ N{����$��BI� QGj�>�J�6Nha�\)9��C�r�98w�yހ|d�r��G��".�*�`r����v`���f�
�`!���Pюi�b�f[���vF0SY���>��p3X��m�9Iy���x�[Y�Zy��cἮw�)Ȳ8Lc�f��ǰ��$��	()0c,X��;f�͸$�J �O���G;��I�&�Vfs;q�x �9I�#i#�ٯ2�����D�ʞ��g �����(� ���Ӑ�w6�TvA��jrp�����׎��)?��{�9�Ec�<m<�S�8q�����89��Y�++��{��`4E�-{�M����s?����䕈�S ��� ���|���DS�1���p"�E��
c�MP���v�|���5?��� ���|t���c@�ށ�<��8�R�.т��Iyk�&�@�u��_f_}�}SM0 ��,�5�9��Ntڷw�]�ٱve�"h�eB��EC�) ��~���p�iR]�w1�@!akh�2��Ɩm(2�UmY^�jՊ�լ�(`�l��$u�䥺�-KR��&�W�K(4el
+�9.��b,U���Y�+����zbxCr�ٷLD).W��ݬ���������4�3p�$j˫]u�Y�+1�9����L�,n�\%���-�0�7��4�3X`�G\�ֶ�45�X��{����|��[�Em�F��4vYQ1ʵٍ�if���7"���3~ �`����
L�$�Қ���]���<��;�,`�jl���i�n�<Rpi�x#�i�13��ۭ �s5�lgV�K��Y�+'��{��`� ���N�т��]��p7C���������x�'��q��fg�w��OE�\kc42�5���m�|5?���A$��`�@"7z�#*�lna �e�+�'���~�<�*����m��g?��y�.�K�mB�������lƀA3�3��A����]SǶ/���]��
����'-��6ӈ)0ra5Ո���UV�3!�`8vf�ŝ��me�P`��j��8E�3�4z�ߓן�~��$����	(�y&�ڋY���y�������~k�c����O� �3�$�	0	0�����0������54c�ܗ��q��da�����j־�\ֽ����Zh\m�"�Zs)��(��Lj޷h���t�}Y�bJ�x �z�E��^�٫Z5����5Q[�G���N>��}�	Mk7/�Q�˻��޸�	�`^8pE�38���Ь���s9�s�9I��9����{xC«o��T�"�q0����@9l�R`�$��	'�ͻZ�_�f[A�p���c�ُ�{��GZ����in �����8��D���+����N,x$���L�J���N˗VAx�9#��cs^��n˻�þ�N8�0o�G�I��hm��ﯟ���kY|)M-��R�Q��ݕŔư�(1xy�э��/m�a����߲����B_?���9��ǟn]Tv�q{������Ucd���ӜM��3��� �E�AI�IP�"�����Tc�!�F�{[qk�,}~��Lf���yoq[o���D8)6K���t�a�Ǐ%޲�����S&��ѽ��ۦ�zq�Ǌ��<��������a0�h5On]9�.c�*�!ѳ9�eX1��C]��@����F7+ڑ�zgu�V�v�����W碍]Y�w�d}}�`�fd�|i�طs ���Kvw�ʻ�c/]������)R�7����M�^`w��ge�s����7�WC����̖���fP��Բ�Tx��+B6���Y��0�˦ �/�A��]��K���p�������Ƹ2&gD��#ae6�m]^�ۏz-���F��ky���|1TZ�;Y/vU�O3j�C����jr�E�>�r�'m�������u!�Z��O+��{W}���6�8=?2Cɲ7kr�;}��%7Y�f� X$T��r=��mT�B�GJ�u-�Z��r�;��*����՛P��L{���k���-�K��b9����2����v�SI�vۧ2�A����-����ڴZ�}VAU��c����p9r�x�l��toV��{�{�l����6����qs���n�iU���gZYʪ[���1��|�iq�i��J�W���	�gJ�ԹoIΙh�ۥ|�M��ɢ3r�C�S��� Y��&e�/4�1��؜"]B��ؽ�d���y[k%�U��BxZ�H5;tr���{�V�q�ok�ج�4�݅q
՜A�[N�N�ױ[�&A�"�,����D�{lX�hy&�˧l��n���H��ۢi|�3Wp$R�E��Z�(;EF���c�ۗV^��ƶ��7/pc�W�,k���률�m�!wj�i�$�4��D���UL��yw�~�'d��� ԑ�@��IW�u-����(5��X�QSݵ̓[ʹ��r,Z�Z�Q�b����{�;޶��i6���1�[��[��r��CX�ow[�sh-���{�F����u�1Qb��$�����ɹ������7+��5wvƉ7�rƍ%<�tƂ�͹�Z+���bMF��ѻ����DF�j�X�lcQf�X�V"�EV*9��#k�U͢�"����k����\ܭ%^sT�[�^nmr�5�ID]���QQTj�Rm�Dd�DdD����'^�p�}W�wy8{��'��/��(�&�mj��m<[�F�!��8 �����\�\׎2����r�?��+i<�Ө
���pBJ�j"���4���^���y�'�٪���yn���x ��`�&pA)'���C����?����96�u1)���S�����n0��]m�"��g���z�<BL�$��ܡ|W�i��Q��T���q�O"[ټ�����&pA)'�C����N`����l� �X���{i�C_=���>�@`v�?�1j}"|BMT��Pa��F�؀AGO�f8�G�dF:�!`�����&q�U�Ś���;��x �"�9�$����>�y�f�2t�U��l��#1È[�η��]I��*�@&�W��etJjQ�;Wv`7FiY��T�H�̽0��	BS�`͹����6�2�}+$��v)G{f�|���h��p�N��U�w}�����$FARAYdEd�BD_.�����;�G{��m'�
dC��^��l��S��������Tb���5۱�F[g:}�������Ģ�$��(�#*����>���c�F]���0�U���f�Y�b��J[2g!Ƣ ��C��r[ �:_��J�x�ȇ�ט�[�[�������P�y�3dm�~���A�C���|�"�0 ����k�!���0W�/�;^�ӽ��3jy;�����������!��ă�_w|}-$8;,�$�A	��M$���,455�x�QG��1��Q�����`AT�� W(
(� ���d��ɏg���&M9�,|��7�z<S"Z��nΙnr���gT7��r�#�m�Y���#�JdA���0��c ��ym��=QHW�<MP���7=X�{��='�^?��BI�	���sy�ſM�2���bI�4ûԬ�N(c<X��4��P�^U���Re�nֳ6�Ɩ�`��N�_z!۽��}����.ekT�> ObB H��"�SZ5J6�;��I��_��u!��͓�4�\K�X�<��@�)�Mi���f:��h�kl+�rA�v փ*�8�4W.�yd�v�IM6iͷ2��YQ��ٚ.�\�[�6e�2�j`e��E�$�r��չ�R�R^�;%b�e���gk�1�ma����R�cC7M[Yvؚ)�da�n˵����3vTB�ҷ+(�6勫 3���³[�^���_��B4�e�7,�Ƅ�p��ZT�M�v������%ߟ~��8|��[�i ����<����	�c�}o\PX�&Xp �*�@9���8!%�L�u�5>o[:�����]y���-��!�3�[�e�F�&ۼ���+^X�`�����
J<�
�\�]�֧fj1�s��N�4L\�ca�Tg@&q��x��	'�$����m�ܐb�����6Y8A��)2�Y'�/�P���.ݑOy��5�J��q����o¹],s �jp�!%�I����9�kE�d5/������r�	ř�-��2���o?�c8#<͙����uʧ�i���10K��1�XU�����K�V�\�a��wXLFgA	t��L�����p5�{�#�P ���(.��։���l=���e�(j�9�[aK�#1Dx�'����!{������5��P�gV�i,�O 鵍KVNV�}:�y]_����w��q�4Ո�,zݳAp��l*uF̠�.ˡ���ʝ�L쬭�w}�gz�? |1$I	)����UՋљ�$���^�7�~'ǟ�דߏsƎ|����6[�>*X��I�Fw*1T�����?�
� �@)0r
Naw��]*s�r�5]
1��3�3�h3���[l̦�eYON���^_uw��&1��D�q�����Ad��������I��5(Q�����nfU�N�\�nfW^wU��TO�`CL�8��r�ׅ��1�l�x|T�j�9�`��
�0��{.(:z?=���� �@��v�"�ĴE�4�5;[W��V��IZ��Mx_�l�״\!�XfP�*��������k
r�g]7 F�g�:�Ȃ.��
L�nټE�H �ݰr����5^��z4l���e����1ʱ������E�"Lk��y�p��l��\3)��VG2��yʣ^R=�)�m��c4DRU�MfH+��uASp�6ά�J��HN����?}����Gc�_jgK:��.��z���X�*Q�TEE�B2BI�FD���0�g���O���e�>R��l�E�"��4(Vl�X(���Wi�u8x�:R���k*�`v��L�!ے�;��&��=���3�	�g ��pA7l��������ݎ��4���32�44Lr�|=�q�u��Eˇ"�������}g㟟L_��L�$� ��Ne��4q�"�t �Х�#mt�-��qp�X�ݣK�����C��r+[��8 �v�b3Cr�߯���1�F�x���ӧb
qS��yu��mcN��Iﴷےˆe�@��\7�~�Q�;�4�n�>��W�77��,�Y�V�%S?�;n�d⑒"�����n"���o�9l�탑v��,��D��DɊ3؄3�f[��Ew�`�r�p.��f�sv�:_�:#�)�?4Ə�4�M�>�e5��ny\]�Et��|��[��Q+�_�����L�1�SU^�{Ob����k���}4u�)u�YXQ��*�{�Q��.���L��NTY�PS0{���f$������$�4hɣ)��,[��Y�:�����3�$ɒ�tљ��k<�_v�~���!��K�M���Y��m��U��|������JoAI��צ���{?�l}f\mjR���!^�#4ٰB��i�B\��eF �!�ٜ6�5�*X9��f̐n�k�5���=���|��q��#��%��)Ñ���-���Q��9B��ޣ[B�⭢ �7��j��c�N��i����9�K ���f��j���a�yeþ�ɒ�L�,�e6YSS��w��3�=(U�6 ^�VNg]�$��dI�g���8"͸a#m�j7���`�3�8|�n�ku�&yV>�� ��:\���ǹ�L�������d}v����A�C��j���J�]F㩟/���1׮�-u�>0W0>*�9l[2d�G2�c*��d�u��=��S��ތ^�V�������C;�ʗX4���&3��
�Vv�;�����M�?�bl��̆͢��B��8�=�E��}�B(�I�
C)��M����}��5���nI�ѹ����QB�9�c�:�6-Zhf���3sI�.X:�6]ķ�,uW����@p��tc2��ƴ��gcp�G9�lZ���&���n�ґ����*@mա���s������!��%����t��e�\\��KH�I^,���D�[ "����P%\�GJ�=����҃��Pn%��ݽo^���z�;�^O~��Yc���Jg��p^1����+�:m�ە��$0S4��������O|��k�w/��k!�b�7s��/k+2����j�	��%�9{t���0m`����탍�
�R�2��u��p�+�<�u�rr��L��ca���pA��>]�q�.˲��\ay f�8^m�CH ����Iݶj��G�5Ю���p�"���do�w���p�Ñv�"�ÀEۇYND�A��;������n�8�]�79����Vu�p �Rg"b��b�s��gݍ�>I�^�WW�h�ߥ��2Nio�/��4J�{���bf�y�������$�I�]t݅��|��y��$����S�Y��͵ˑVⵘ�[���8.K�F��~8��	�g ��G��}v�&-�j��
c�GxK],�2�Q\�*7D�I��nʣD&��fn�a3,�3:�2��=v_:�����-�Ԩ���-w)2&4�v�P�X..l �9c�]�4����u���,��ϛ�2إ4rڕ���Q��_o�3 �LL&�O����}�����z���;�),�2�e�[p��޽oO��<�w��GA�����8#q���`�]�pn�8 �v⦻�N?g:��ԭ=�R���FV6��y����A�p�]���>6�7@v��:����K���W���l��̬@�Mkp���8d7)`�"�9e����C���q����6\�p�"�]6B���B�BF��@ƒѷ���o���N^e��p ���#���}rޓvձ7���w�SC��hS`� �� A���leʲ� �7#@v�Ak�h@�m���\8Q�0�0pAn6\v����՜�=uX�{�L*�*FcqYz3X��#�; E��͟]��|n��[��uoQ��$g�3W���W�r���Ok2$p�<��İp��C'�ΝP��y�����(�2�2��-�k)�mf�]",��L�2\&x��.��ׄfT��ga��sz,�����$m�A{w��7�ܸ��rup،v��0��k��~�H>}l��;]L�-��M�	eM��뀓w{ ��pE���-��hO.a����[ ��ý�ugv��꣫y���"mҝ�+�����Yal|݆eu�ʶ�9�me+\lK�C*�L�����Ț�k28d7`��p>�"���`��v�3�E>��|�z:�g!ÃDG�X��7a+��m �X5M�h�:
�-
����������0r2���ݿ�vf�]N����/f��r����a�z��SzM[9l�>�`�#���5Μ� ��p��6R��UX�{�\����oz�"q��_������81L� ���A�?��g ��M7��8�w����v��h��̎�>�`��9�`�]�r.���A�V�"{=ɘN�o4x�o�]y}�+�P{̵��m� �M����ę�=���MU5'f��3㙟ź�R0&E˕wj�n�ɭ�-�U䤲��C�Y,�w4��d�vz��V�/&"F�[�� �N�{��y��g]���탐}v��n���}/m�1ü|�\7i�*�:������;,�8r.���v���}J��k�l�c�������i��P���8BP[Zѭ6�f��l�e鰳�����'���m���pAf�h�ݬ@��l𷕊8l72�[��іLݮ�BM~>7.7lk��,���І�޻oH�ً�M�,���m�A���O�xܚH�B{☥��P� �r�zְ�ۇ7lEۋw������NԶ�5dUTe���=s�vX9����?�{w*����j�we�ʍ���|m�]�լ�D��m�U�8i�ot�vv�m��� ގ�EX��E�6l�7��kp.�3�ͷ�Ƣv���֠�A2�Y=v�A8���Hpn��)1I۷N�v���n�|v�۷o��rs��MH2�e�t�q�>=�2����s�sE+�V�ݹ��/Kw�	ffĻ#|�∥�nPlT�B�+l���$�&$����)��!/1\��Y�x���{3��Z5����5�F�_�3�jw7�གqb_i�N�(��U�\����b��up,؅n0z�e����w�2���̬��P�G �o;q$s\|^ͳ5߭�^e�jH8X̃J��񰹛��2����/Y̚�vtl�X�Ƨ2�;u����Z����ݕ����_L5�ax�M��e��
'�1p�}�7y#qgi˷p�
�m��$ZyJ4-T���C�q�5�WeU����Ҽ�$n]���ݥNd���_���9e-����9Y��3��`�I]2�Gth�wMN�IC.in*�sr�� @�s ky^#���5u�7iyEpF򞁸���Nm�S���ɶ���wyj�5t#t̶Ʊ�ۦ/@���ٖ^D���5P�%C�][n�{"N�hF�X�i�T�v���"���\�u$ ��7�΃��&�6;7;9uD5^q^v�9ѳ��/�ۺ�&���'5+^9�٦�bΥ�`�Α=��Z�R`�lXzn�{�2�ފn�]������f�3AqZ_!|r�D�]=�Q�}�+� A4�
-k�P�I(�o����{ �,�KFٔ��^*��]��բ�hk[�Ƕ3-��� {�&��Q�r�N�������c�N��WŶ��-n�vӫ���gr�e�L�O&d�s8�n�>�u��?|�*���
N���쥶���bE�I�Ř9�@�G�$�Plm�7-�ݘ�����;b-F1���X؃QF�eF���6Ɋ�ch��Esh�Z6
� U��;�3mҮmwb�6
,�
�k������j
幬h)�cb��5&,�����j��wua�,jwk�S"�ur+ssb1U9��k�TVf--\�Ur�Y�uo5ylk���I(���W(�ks�wII�ӿ;?_,�&���\�e�\ymb�l��jr�4�J���Be�l��rXS.�UɱWgW/U`-v%�:�P���e�cΥ��!@6��hh'�lkl.t��"�DA�1�J�dm����#u��5����ی�Ҭ`��ՅL͕.�J�m�& �٘�2���i�Ě���x��lԬsk��V� �Me��U�j\�"̳mFf�#�R��\�f�W��1v�39���Q�y"�؍AKj�VZ�ge��]�Ռ	�2�����2e�D����G��;/vbn+�ڂ��m�u�\�lbhF��Ya�kCTf\�mU�L�C����Dj��me	���FnwjE6�ڳ+f������Z�.&��GT]{i�-bڤ�qU��0ˊ�5&q11c��,[S�+�[ �赋��,�G췷ƍ�[klMBҲl6^�26�F�H˓JZ1���ծ�4Ԧ��ڏXP���UY��YP�W%X��1�6��vuMlx8\��͒�c���J�g�a6��P7��	k� �M���.��7���.�X�<�Y�	1���n�����k�M
�0r�Y�R[�����R9���MǷfXA�5�h2�`��m%�X�=b��J�.&@��7iUr8��`���-�]B�U��e.�Jg��S�ca���cB��KB�:��ݐ�g4���4S4��;��ٍt���9"�����Z�M��&A떋�n$���j�)t�sIH �s�Z�X��	�MY3)�� j�@�L��TK����ͺ�hm��([V�s7b�J���Y��m��koд�(�C�&�GdfL�ȻYe%��i��͍�5��-�+�SJ�$�Rmv^�q��*���K�B�aT�F3h��Ƭ�����5� ,��;cY�r��	���X،�f�cj�kE6��t"5m	es���v�f+�����]E�"�p�L�[h4�6�WBӛ�LZ���Φ�e +��
�͇2ܪe�-��i
��͚a[)��CVRXm�Oa	���O_G�<�J����rJB�YIl��1���ZQT3qkB����)[^�,9���Fٳ^*��rF:�(�	�1Wh�de��h�.��ѢqB�M��ec�[]eG�-6�!��e+c@���*��Q�l�2� �B�+��4�l���g�����u&�bh�-���h�P&6L1�6�Fi�u��.�Y��+ N�e�p��R�%�I�tM��R�M��Z�	LSVT(��b�4��.0֠�Ÿ�0��t��*X��>{��w�KuU?YX��#!��B��&�G A�c��o��� ����M�}��a��woy���A�gz�S�~����-G{g�@�`����ȻfٓX/��h�a�f�����.��v�.���sA7[٭A��O��:�&pA|= ��J���>�B��୺��3�Eۇ��q�[�Z����4��F�9R��<7(@"qÁ����g �v�ݰ&�F�/��--A��g��IL��w#N��w�y����F�v��ۆxfi��ϕ!��u:�3������i`c���kCC��j�u��,FP��i��I�rg\��o���`�fb�֠�ɓ�Y����Wpj�Z�0s��� >�H(܂����߶�ޚ�'M���i�0 s"l�]EV?9��Z�µ9|b�f��eic;���)���6�)ř9��Q�l��N�adL�b�i���}�)7�bp�����O�2��V7y���F���kދ�/�g#�=��C��ѭ��p)�������t$�t�Sλ��ʩ�l�e�F�͗"����q!��s�~�Q�A�p�����k!-̼�j<�>$��ۼA-�.�ˠ�cj�ko��p>;l�]����v޻`r$ɫ�hуb�?�����٘z�(�x� �r+8]��.����������</���Ⲱ�ipVb���6�6�L�ƚis�u���~�eγ��q>0�9�)�]�RRa�v��>T�M�U&|f�c]��0��-��s� �����|ٌ �~��*f���0����-�Y��y2|I�9l�����v�0��z.�T$+���z��'������z턂�q~>8��j[a�B͸`a��OQ�x�����zs=T�o�6�՛��駲�'I�{uz�p5x�_�,[;ɟ
�C���q�C]v��(]�Al�D=m&�3������ؙ̲��3*��7~�y�y��}����'u�A�gIV)0��epYS|57{X1�`�cN��#6���(Q�`*��I8 ��� ݸp�!�r��L֨�L��@�&O��5[q�g �����]�ܗ}�x��[�s`8��� 	�Y�e�6T��l0�l��m4���@ �n&�b�D=;�!��Cܲ�e�fY�ɘ{B�x����7�Xu[v�`�X�c�~Yd<�̬��52����d5�YJK��73�R�ѺEL�jg���CG^��eE�Ӝ��aG�86d�ǖ;x� ���n�w;�.<An�]���[Y�[yֺ�Ѵrd�i�K{�XG����&-���H�6t@�w�t3��`�Z`+|A�ۇ����2��������F�9��&��v눡���b�M����-�*s�ٓs�U�u��aA�ve����C�^��Y*�5��%�;i��֭��}կ�P�B8�^���z83~f�ߟ�3�'�Ql̫�fe[	3(?��i��쟻m�+����9L�]�p��Wr<L_{s���<��Fc�l�]��Q}������G�����Kc0�m�t3K�kns,�rL<�X�/+�c�Mlf���o�y���,�=��n�&��_e���%���mgU�íp���]�״F��Ss2�#��	�`�"8�M|�%РD[9�Ë���\�O}I�w���g��OX�fYLLn�t�<f�M ��z� ݷ	��n��r	>�P�j��2l���g���{E��G����XBovXJff���Ns���+Z ^�pF�� ݰq���th�����m����r*���|l�9��k|oA�;��{�� IÑvہF[�ޛ�B`6f�!�8�S���n��l3�e�P�F�"����v�<'��{�Ǉ���]Q5:|v�b`��/���碡���;���Rw�)v�#z�,+fQar�r:X8{�#b��������7�oy8[��/@ͯP�Y�PX.M�]6����`\��B��c{jv4t��Uu��!�����asIm�[J�+^E4`�kX���5lҀ'������5�kPf�1*�c�@�0HlYN��,a6�Aa�[���G��,�2m5�@m�l�!�W�Z8�7Z�ҹ,���(Q�\Җ!�l�S�mAĤ��0�m1vϪ߉�D�rcE����]F���v�P��Sd����2g����������ߗC��ټn���S�Y���P���K�6�QFn���E�� �;8!c8 �v�]Ϝ��4u��f���':$�����n�E9q���`�M����]��v��r`WH�;Z0L��mÂ��l6\�������<&�z*.j����o�Q��r�
�7�5橽.�[$�m��6���si�A�g�쫌fj�޼x���`L�Eu�,�[1�`ӧK�A��BT���.)8r.�1��F碙σ�r�i����y�V�'m�G�xɻg� ������ӱbL���˵ۊ��V�t��̨kE0�ض��LCfAr�Ŝ3�y�\�1��6dv��!m�]T�]_M��O��sŮ�Fټ�}������d;�|�4�A)3��>��_?qN�DU�J/mzƊZ`��e�Dv��=3s*��\]�u�Vhrν��Ju��49��q�3=�h��/aU�^a�Sn� �r��za�G�p �g+j�������h�Äq�`N6Y����F=��x���p�d'��l3(���+!�i�ΰژ��]��Rl5��m�v�Ⱥc�ѹ�\���갠&��Iѫp�� ��ËZ��s]U�U��q�j^�c%�<�27�������̈pn�� �pE�!�n٘gsn-u�~�\2���Y
���"�8G�Ƨ@�e����p�ø���ii�����YI��ר�l �L�l\5���l��4��r�~6F{�ye:+,3#�l�w�^sgo6e��S,i�۶��S�ogC,�l%��9���l�Y�7l��,eNt���A� ��W*ռʨ�U�,q�k��� ָw2�F�Σ��}����G���ed,��p�̪c�&�]@Y9,�}r�<v�CeÛ�6%KjAyc�I�'6E�Խ���W&ʁ!����˫ m_��^��A��}VZ��w~a��|t�'3�8Gx��qWW��4j��7R
7R4��a�����-7���^f֭ٗ/�әԛ� ����o�SM'>t�A �3�f�>p�ln�9�g�Ѻdh���N,ɾZu]�����;�|p�p�`෍���!��k��UmPѴ��+�),���b��!qΠ�Xf�\F̔ƭ0M���֮WW��=�V�=�V!����]���%�[cE�I��Q�8fx+1]�#���p���� ���.���>]׭��&v��DK��C��kz�sg��Nc�gR`2���[q�=�{���^ja�#��\0 �`� ��Û6\�.��	tOz�Q;�X����垵��I��Hw�-�e��+!`ݳ���]�m��O�[�&�UD���O
W*�<0�y�����Ǥ�=\}>���{�$�k��9(`�,	M�_��w�N���[ǷkQ���t�cyN��a��b�g	]L���V��}S>�u2Y�gE�d�p̢�fr~���A�����vU�vw=L��̈������x��C��M�o\��ٛ6�+F�F��`D�Үa�t�-�ZܩY�����Y�J�Â�`A���>�Y�$�����OV&j��8�5���I��Mc+��NK�9�,���̬��]B32���u�<n� �Ak?�֪xl��JҾta\��ȼ`�ٳ1n{� ��;35eï-�ɹp��Y�l��\�h,���}��"a�"3:���7�m�G�sv��3[��v�DC�.��鬘a �p�ްv��W=��TX���X����9,]
�Йo	�l��1��>>���@n��5R6g;����>1mz��eե|,�I��zX8 �8p���n/���m���~����I��z3!Ӟބ���S�л���a��롇�����[�Qˮ`OD^�Ml�pB�9O����~��e�Ұ�^���mMt(Cq�p��&e��i�tM�\mPH��3G\0��bHhV�W2����V!�RlA3���-���N��V1�5��Ђ;�e5�
 �ݙ�1�Ya b`����v�Z��(%e��˃cntճv���3b��-sD�<��5!�k���Wvًj]sb������pvr[�^���}����T��d(�n� �C���ˋe�Yl��J=���/Z�+R\�k�������awe�2�v�^g_.���fFgV��i��w�s)�߶�]�̧&t�I�E��WP�����������p��_u��5|gw�s�p�pEkw�m�r��\'Ǝ�����=��	���zM�f�1�(1rqT��/�,�U��W0'����͟8�p�]��p����w�ǦY�Lx��E��>���ݷݜ�����fukw�'m�'��s���r��*�Fw��23(/2˙2w�s;�݃��8�ŭ��\�5W�)�y�?��rk�"퇜[Y�sT<_l���y�"۱�	���&��1��)&2��%��B���/Ӎ��Y��pn��A��NoK�6��t"�s�S;�r����#�)Ú(� ݸr��6\���Ջ�n،5��<��:k�Ȝ���uq��dD�B�̸|y=���m��bW:�'-��h݉Yl����ѡ7TLU�$ʍg�Ʋ.�S����)�Fe�n �M����ݱ�<��^��fw�V�ӏ���<E�z͟Hn:{�.�!o,�H�SFy�o~��nu.�3�ܙ	ә~}��̄�MRL�`��C��pA)7[��t��]f��"��qU=��$nMx\��9e�2�!2d�fQl37�DoǬ������9'2�5ٸ�&������	�g �M�9�g �ݱh���a}{�����'���"݋	�Q�Q�{8J�M`SG�y&�gM��骎
0��S�/����|18Qn�?�EwL�8d�y��X�-19aq�� ���w��p}v�'�6b�����!���X�T�A��)vb{.4#|�L���8�U�C��e:���MΘk2ˆ��fVC�1�ێ��^<w���{���o�߽������l�$̣c�}w�PX�T�Q�>�y7i*��Vp��;\wB��27�MK��xV]�펕�a;V���c�;e�Rk�Ź��d��C��_�w��>R�xV�ʃp�lhwn����a�-�;Y}x:�8�g�R��ۈ�ʝXW:�jW=�#xX� 4mXͥ�V�:
ve�5��.��3(df��
,l��:����4�:j�n����:gV]'|fv�X�8�:A,k�j�"�=�q߮#�M<N�� L��\x{(�{�jݧ{�j�5K�PE���E�]X�	��s�1ش�wu8��޼u.��c�WWW%O!�4k��C�]!�ڲ�N:t֥[�Ma�|i������݈띹Eh�T���ef⹤T�9�q`}F��8}����3���Ӹ2�E�\�9u ���N�-�<o2hu�Kp(9"PZ∾ҥ^!nee�I�M��v�N�[;�v[j��6Fu���b��Tfw�I2wǔ7S���Xy�|�)=՗�6�fY�[56ɇɍ�h�� �v�w�d�u�<�g��	�	��J�E1ca�f/��}��ԋ�)?�v]�=c�Э�m�*�}��٢���IYPi@br�+;��[0k�y׉�f�{��-j��+KU���׵�kӣ:�Ӓ��L�x����ZwN�J;V�7�k�u}�/���� tq!u4ӡ��E�m� �yS�2V�k�ry�xu2�'k��t�ދͫ�b�h����C�ʠ �B뀼����_�:+�\T&���u��k���Ù���i6��5F�6�Q�+r��nj�5\�lQ�˜�m�Qmʋc\�Q\��TmERksZ.c��j�#���r*��[e5cN�F��ͮ[�q�F��k���ܶ-wus���ʢ��Z,�Z�u̓��5sr-�ʹguQ�r��ԅwu�Λ\�+t�5����}��a�c(����m�ri���gI��YV�&]o�߲��o'�ha;���v���Ū�E�Qk2[�냅�>؄�n��X]���C�v�A7l��-���X�Yg
�r�w�kq��C.ŉHЍ�	�`� �8prd�̳+��V�:뫩dyrB�Q�-�a��瑰��6ct�`��H��k5�cN"��߯}�J."�Ñv�k!ﻵvts�LqFgN��Yݘ���/��A�C��r7l�Y�`M���t�n1���;�c�������yk������Z���e�Y����A�%и�/���,+�Q�8ޱ!�o��"�ȟ��>56��ěxI��0c��m^�5F�[Paff%#���h�9�B9�.d�a	�e�̲���V���}f��4j���%�������!�0�Q�C�[�A���C��Gl9��T���b)��1�90�a]�:}��Z�\š��������X,�y-�%�;ΔA�AQѹ:*��V�K9ճ�,���7l������ ٳ�>B�b��<�wl��7ZL=;�kt{2u,��e�3.�ed=ky�]5�j.H$ ��Ėf,a��zˎs�*4B��9xk�3�T�HQ�SZM��z�D��6�ݳ�7l���#�xK��̹0�0�W��:t��ɮ���s��l|�(p|QE�"�*���!�u���l!�v�f?.�0b�Νow�[?���?��>͉���9E��i�q>`N;s�.c)���d�d!�eg{�����Y+��,SBx]`60^7y�8&̗�[��4}u!>�%ѹ��,?��"�f�e��sI��n��WV!��K.�̹0�y�e���p��C\Tؒ��qI��y�P"�9$�$ ��yY�f�
�󈾽�����p�Q�ӭ��w��oP)7�����
���2�SR����%v���us�2�Øg;��˝,�N��f@ն��E'�r��Zw<�z����8���gZ�{40����~>Y�?gޱ��Ou��Tx
[,bKz�����("mE;p�M���Ms,900����R�rnv���5��K�3�j"6�I�\�q��u�;�8��F�Z��͵����{;8�+�������4(l�-�\fi]�&bM��R;X�Ɍ$fE�$m��	��
��f˄#����J�15�%s�M��"d��ЋSev�XW ������_>�?Wf�.a[hl��ȁG��X��٢�-M-�����M(�A���߽>_5��T}v�1��y�E�ZN&�:aMU�oR8xEۇ����ݳ�M�z"�M	9�[wL���H ��q����vT�����0�y� �r-0pl��\Q�7��հ��2p�_=Dx��<|�!���N��d&��&����~�����0�Q�ӭ� ��p4�C�n��n��mǘmo���u��; �p�J.7n�2�����<N[w�0�l�pE��Ƈܺ���78�m�9�gn��"���Hά3BT��uݤݤ�z]��-�s{%��}iÃfː}v�|�~�����M<�?M�鐢����P. r*�:���i��P�ՆĦ��q�?�c��V���m�6E�K:�O2�#FgV��p�\(!�b��	k!������9m��v����5ٓ�v��L$I�OM���ņ�'ixY2�nn]H�Ղ0\�+'3>Y�&[%�otwV�S\geٵsp��v>���ɲ�e�uѕ&5�x�rۼ�2g��D^���#8��r��AI��6}v�&�'mڝdw>t��2���a�no����6�9�e�l܇��ǜޭvf�.}e�[/�6C�K:�u2�"��s�[�ku��q,ȕub�"K8>�w4ђ�k��h!��&N�=�ټ��禩@ܵ�§TҞ�ɹ�c��n�pI��l#�,��lr��U�99�4_Yߞ~���zdg<����tm�������%�t6�,�V6�ʎ�ls_'�^ϒ�/��d{{����ݳ�����y�5k�O7�����A��4G#,�����7o��"�Â�k6`��)�v7a�]�B��l!�-�]��%��c��N�	�g ����۶?iL-
�[q��;8 ��`A��=�ό l�pAn/�ʍ�E���GvF�}n޾��I�{�n����Z�ۓ@P�3M��U mJ�{3���>f������}e a��!܄�f�bܙt�e0BL���d��ȈISÍg�냂l�r+X9o���!��glf��;L��c��oQ��́ݳ��_&��]��xi�`A�`�T�l�Ή{�����Ȼw�]��w�@�BQ�5����vSmo�5�uo+Y�n*�hc�gN�	�g�?���v�A ն���BM�����{�X[�_��]	L��]պ�X0���)��vJZ�`V6�6��|�=���Vb�����pE��ɬ�ȍ�,]{ИC^����0���dN�����v����\���[p��Op�9��|e3�M[ ��Y��j�f4���8 �pA��Ȼh��9%(E4A�2�9�8��v�Ȼp�&�y^k΍�坸l�]P��Νow�S8 �Z�Ǎ�9ݳ�]����-X���\�x��Es9lf��K�Gr�.�=�\E�9 �7�9��N^���")��"�PJ}/"�I���e�ٵ���8s�T1S��N����,����y��Lf彨�$e��/��� �e�*�ꮍw�9�gv�	$�nۗ.��mJ{b�Y�o�Ǻj�Y�ծ��ׯ3���;��G{��w�d#�eY�������{�:�O%^x�	if#NĀ.�Mrv����v��)Q,M4�;��r��߫/Y���
��`.�Hĳ�gp��22.�n��RK���h ���ŲƀB�3&p�8 ݰpE�uk^��.�L��d���l�4���.=�\����rs�v�
��Fc<�췤�
���`�=T�T��3v��pΤϚ3ʯ3��m�pA�`	����rۇ"�Ë�����N���~"���w���ن%�w��FL��t�u��m�!��޵R�a�x'�v^(㳐A����	�`��]�pE[6���y�"I�0G8p7�ksfz�K���y��A�v���v�||�[�y�ؓQ�	W-&MN���W��<��yehM��V0�"�v����-�]����6�9}�ne9Z��Y����9��}\.���̘�`�+����-�LA�;kq���b����@�]��r�j��5��Q�\`���s*�����٥�V��k��`�U`j�4�]��ڇ=��Ya,����ݦadNؚh)3��fP��CE
̅�0=�4$�g�8�Ƙ�Y�L�(����qFm�U'��۳�spp�f�eu�s��)��5���څ�-���m.#�����翿E|��ya�n.в�M1���,<]�͍��H��M�5��%�ӗ��Vߏ|gϻX8��ݷ_N��$)��O'}[�q�Jf ��zXH��{VB�Y�,�3)�u+�y��עb;��h"1���0q6�jƽ�eT��|�8� ƻ�A;l�����y��A�g����`�����Q�n.9�b��({��WL��.{7(��a���~�i�m�2����W�����N�L�v���==��\�f'�ޭ���j��r�k[VO���v\3,�̦�2�!���n�GC2���p1o+M��ʩ����8�A;l�v�9�gv�ËS>a���'����s�2�0R\��x�\63Cm�i�Ъ��!+n��HX8������޾~�u%����}`�!&pE�ՓX��\�Xnw�îp�k��Ɇ��N���1n�v���v�A�7l�?������	�O�6��Jz S?��̍Im�^o�闹͐9��o��O0�9�C����]��`�d�ܳ����,T ,������μAY����;y��� �5n������fd��V�vX8 ��Ȼe���	�o=-|��A]�d=���=��̲���.�t!Sx\D�l�To^���a
dc�gN7 A;l�Z޻oH7l���;�����o0n��o?��8K����6�k��\\��t���e��;X�;	��d̫!	�VD�̧2�5�:��NƇ^�j=K�#�����ȁ�����`�N.�����k�lfS�E���ҫ.�K(޷J�h�f	��3SJ�J%�s)�	�7�pH�i�0#�Ñ��M�
�ͳy��!L�w����![#n�r+i��Kz��?��ۇ�Cu�)nt]uz� ���p�D�f��f�f�Ry�"���EZ׸��ݗ=T�}@�w��@�ʸ�Qd̦əQ�מ����z��w�Y"��kN�O:��q�I��k�b�"���b�9W�;�s���&+3����ڭ�s���5��$�nWmm�<Nc����P�FB-wYk"{o�rި-�~h�3*�L�,�ek�6V��;�@���A�����v��Z�En�0�R1�3��ַ��a�e�cו�9��m����9��Qd!nf�̛v�̦fsA�����V�hݦl�#�������g ��Ñv��87l:�Ij1�����Y��ap�uݰ
j��q�aT��(#.V���ٙI�o�=߳��� |�c��r	�k܌��~L�uֲ o��b�fk[��O����Â3������E�?���5<q�e�[E Fc��A�`�����7��B����8�e7x������3N�k�U�ܰ������8"����e�یg�?;��bЕk��4i��Kpf+�9n�&탃v���ġ��ܳ��'q������׻Y�������� �����a�g��:��Y$?h#2��xh�de��-�<2]����e������N�78�ڻ�t*�t[#�ە��ܹ�̭���hѠ�X4����$W��������	l� ݸr.��E	;�k�?�L2��������:q�A�g ����zM��K�Hv�m�ǘ<y;��v%������gMD�Zma�RQZ��R��̴1�H���_�����*��h�8��CFo�� ����G;A�p�;{�472/9o��U�sv����`C���M�&�c�w��v��k��7ֲ`p�p�=,�3
�|��s�g�p�"q�F�pAnv��M�Ui���	�>���j�Z����:q�m��r뫹T��||��"��h��l��=v��s.�w���x�;!�e3:�����6C̶��<�2�����\��_�����`|�W����'�@����L�g8 ��q�c�v�E�	�=�8����۷n�|v���ǣ�yF����W�`��z�Y�1�HXt!i�q :W-�ff��|���&vg_t=��Щ%T�V�m���~�̯�П&>���
�&fE>�/�c� ����[z_h޽���[�Ggr�R��_K핛��Y�:��kDhե�;&��F�^wL7K�{v	��y�r�4�OcY3J/G��mm�/1Z
gV�2�7nl��93��4<��i�By��,
セI��e��)�3��_h�+�L�|r�Tk+��[�)�m)�VQ\l����4S��:�v�P��LεwƋ&��Ãt��p�����֞�Ⱥ��)XǮ�p��s[\�����w[Ά<��:�W)��v�;�[����N׋u���E��!㎋�qҮ7��f����Ѵ��#v����w�WL�Aׇ/z��N�f�_ucA�|W6�Y��U�{��"��x���s,�8%q��w3�\�����,�W�{wl�ŖN)��C��-M�1B���8���r6�%yS;����]>��6���U���YW��!հ�� �Ҿ�W�ǣ�8ڼ�	�YoԻ(�輘�Lu�U"�F�p̘�;�iz��j�/k�{3���Q�mϺy�Gc<7��SG1KYhۭ�ӻrG�U_x���r��K/���s�%�Z�hF�e^�F�b9Ӵ�4��p�ܕ��t�{�,�EBw���u;r�X/�g-��3��
�.`�ygj�E��dޡn�JXlW.F�؊b�(11)eh�e��b��^�U�_z�F���-�j�ۛh�XţQb�`Ơ��lg8���S�c�Mˆ�� �\�cF�ŋb�͝�\���[���+��[���ӗt�Ȇ�(�wR��h��h�hф�1�WM�F��ȍ+ţw�ƻ����v�IQq�gu�4FM��4[ͺ9�Y5�ģ�����b�#C31�=�fX�&"���s���H�@Y;�X�&��h�)&#	,Q�-���b���-��"�D�\�Q�$��s�`���dƇw,LN�&�3ߋ{���k��mA�3�Ff�bA�Pu�jS[p�����=RSWv��!��]�M��t0���Ʒ��b��a,%� [ɦ���ìP8�&R.̳���[q�KLvqz��J1i��͘ĺKE���$+1Z�� ���n+�k-*�ڤ����eD�T�0\,�ķ[��O���S�k�˭$L�T�(l���0��v�Zpf�6��a�kаB�mIZ�%pٜ�5����f�aELA��+R��q�ِRY�hq��r�$,�L����T�-�ţK�#`ʍ���]G0�M`̮Ղ�i��RLa��`YoP�P(%ۓ��c*9����XG��g�V�\��4�C�]�L�VEBB�6-���pL,�tm�كz�`��YH�F&����śT���j'R:�!r]CJr�XM,؆�f�Z�����No����v���K�A���I�I�ca.�(ͣ�KV�m�1G�8&�%J�u��4;E!���L��g7�2=��9�鮉2�@�et37�,攌�Ab.K4��%V9q5
3gWaQR:l������&rJ�F��\�٭&7t��&�+HgV�]�ƹ�Z�fn�&ui�s�X+��Qťݍ�"�F�&���֥�D�;J�ee�DfC3��ٰ�* 'i.7���)<|�0,�j�ik�1t���KF�XBm��X�í�(M6��I�ݭ��ل4tUvZ�Z&1�1��)�c�k{ j6a�l�鍡�eV�kV:��6R�5�@��ML��3Tp����ee�Au�e���[X�6�ڣ�)�f��i����ZqD�BmZ0�%l.�f���Gm�1FY��ƚ�!0f����u��,e�P��-Xl�.٦�����2��l��gY�{+�N��5꫐��Q�LU]��t�敛��SZ���,�m�klclZlB#�-��\�FX�-�ڱ���  �2l�l,�Ȁ3E�����\mk]��p���C���	n)q)�P��^K��ϓ��g�/�䙵�gX��K2!�+��x�)�&t��I�֡�m�1We�(1�	n�ѭU����M�J������%��u�Dz�ia��j�s�s�1�����0;4�#��۹�hfW9��B�9�╹P��4acl�Cs��jU֗A���62s�	R��Y�Xu���+��,M��jR�
'$��wm[�Zh�%����eW�W�O����?;�	�KZ��N���Ǔ,Բ�AaRa9�ցU&�SV2^��{���E��ָr.�?�7l*�g��W3�p�����sKUl�|wҟ��I������fe\s(��E���K�����y^�P"������fX�ϹE����!�"m�����yav��I�D��׹�ו�#7��@��\̫1��en�3 �ݥ���[���������Y���������E�8 ���.�8�%�f�lk!k�FӁXޓv�����G��
�+:q��np����%�ra~+Y�!9ʸ�Qd̢�f]���{9W�/��	ë�b�:�-��������Es"���2����Z�3v&������,%����c�[4,D�9�[4е�y݆�29�G�c7l�|n��([y���뵗#����85B���xg��wF���ᜫ!�M33��ʲ3�p���`�d3���N�=�����.���V�?wVa����b���we�C޺o`��3�)G\�K���.�Bi�z��)�U�n��8�O������mne^��a+����A;n�e�sv��#�4g<�r˴w��p�����d#�e�3*��N_�9Rw��b�=mX���������,�]�����y�"��v�+�M$w�9�gvժ2�Y�;vU��c}����rY�֣"�6�"u��n�]�pE�y��p�]�g���y��;��*�t�#Y1�Ӎ��pA-��v�&�O���G�~����~���;�0��
]�3p�tۘ�1�K�y��Kn�g��K-�X��f�f˒H�qZ��}�M�����r6�4�p��"'9�?��`��]����O�9:�|a0mIL���ʻX��Ba�e�p39m�Fi7�W�_,�Ǝf��VB9�Y˴�v�<}ZsuvN0An����8�Ӧ�_(�/���?�3�oU���{(��ۉ&�f�u�s*�C�EP��h�q�C6M�&������'����5.EhQ�Ի8��N����t��޽G��Ɍϧ���9m붒	�`.����l���A9p�|>/��!&�2��Y�(�77�$(���i3����:�+�h"���ǹ��m�5l���3��r����w�wb߿�๩71�g$d�pAX��E�?��]���_WW�d~��~�O�D-͹2k,]fH�`Jjnh�\�b�b��)�u����z�O?}� ��pA��]����C��݋/Q�fG.c3��d&�]���/u��Y���A��Y�o]�z��#��Tvi5/��%�A��k���?e=�sNs�d�s���ϼ�_$���~�g"|W0��)��v�x���E.�x]B
��˅/97y��C��	�`���6}v�Anb�Qo}�r�0ɐA.���md?���˽�ݕ��8���:���>L6sLY2,Dm�¼���bi��zIُm'gpL����lf���	�l,�\R��r�щ���yT!fT��Rhͦ�i�kw��̧&uD&e�fYlɓ{���{8I�ա�[��0Uз;E���S�\�l� ��] ]����FFB+'6#�un� ��I��pŋ@�-����fL	H1� �XY�&MM�ㅔ�)T���~z�{��������Iݳ��T�zzf2��30�s�����;u��ax��Ӈ8t��I����pA�g�7���3��B�sq�՗z/��Os�Ս���FϮ��XU�9�4-%@�Ɲ�f�0 �`]�6|�n5���
Th�a�!���i·]���nY���^S�u��˴���-��v{��.�H-�~"<k�� ݳ��U.ޞ������<� �������7�dB��qw$���6l� ��~`nȳn��;�̈y���Y|z�5N.�op9l����{"<n��ƭ���ݛ[��l{�-J^���7/c5�e�"�n�Cjmݰ9�E2���}(��t��T� �c�	�K&D����T��Q�4U�u��)c�L�|Υ"���y�ߎe��H/�Ulz��kSkY��2�*g6iq�+�]խ�)4f�!�hm�VYpՍL��ے�X[0S�LJɌ#ni�L�j��u���Q��ne��a�^�H�m�l�(53�s1�	q��wia�lNl��R���sc.���-�#qU�����l�.5B�)e�%mDK�JK���8�'iV���TRZh��Cm�>;}�}>o^�#��u��D��(M�%f�Q$�.���Ҥ��x��c�T�����`N� �?�ِA�p���C�Aʖ�<k\�XV6E�Gf��5nv��m��� ��x5��A9��9�o9\�V��oO<�Sե���y�%����ٲ�*!��&���-���gK��I��A��0	�cO��R�U|z�4�-�n�<0��A�޳r'7}�����C��oi�> ݸ
[=���Q���Ƶ�n�f�9϶^�&_gi��ʹh�D���?�\���܀�H<n@�#\~�K���0�"s�OD�S�Kh|nrX8 ����	 ݸ���R�Yǀ��#�	ô]�`4�%����q]�x�j"Ѯ��)f[�p&�jL� u�73tXB=�e�̰�f[g�����x{��P�9}z�EIr���ڻɝ5��"S��ސn����<G�`����c�U�S���@����}r�)�X�=��H �拶�a>,*�U���U^<R	K�ȶ�h�XSK�oz��w\8�۰̆Q���Ƶ�n3l�\�Ȼ�ݹh�n���p}��n�y�7l��nۛ9��	�۴g�1'݈�����?Q����n���F�FCU"4/h[���B6�������L/ <��I��{��oab��r��z���r2�n�>��J�h-���?��`.�I��v��:������٣�8p�����4{�z�\&a�Ű+�?�7n�]��/ߗ凯����^|�|JC"좲�)1"�YF"�L�hТ���L��`��[��r����,�~�0|7��붫Ȝ��\�4�d�����<9 ���x���H9nǓ.�9n��6}y-�}�Ъ�0��F�#��N�w��83������[� �3�}}���!TF�Χ���l��{�z� �oP�q#���A;oV?�P��[h|6�;����Y�Tם1�����}Z�Kc����e���]� ���d4�V�3<b%�7�� ��l�Gw�s�c}�6��`�]�l'gΓHPPq�)�ڝ�c�p>�`�5�M�8�����xR�5n�_���9,��W�vwDp��A�Â.���r.�9grrъ�pY��ll���{��1�4����ԙ���7l�;؉���c�s�ܖy)���hh$0ت�fUb�R�!�.lx륶�MMY��Vk�Kn���=��y���/�8"��]�qN�j����ox�w�w�v�.�P~om0��?�7m����pE�s�VOuc�k�� �TFjs��s�V��}z���Z��Bh'rOONn\��.����v��n�&킋�|���T�f��A�'F��S8���Ʊ��m�vޟ�q�o$��1�7	ؚ���` ���/ g!&
�N���+{�s|W8����k������ڵw�U�jO�=��hmf]�9��~��Y�b�vpf���nCbY�n�=�-��)F��F���N���hn�c�4�t3�S��<<O;���z퀻`*�X�l=OU)�飼��l����m�s=wY��O=J$�.�ud	�%��e�^U=�����~_;��g�!.�Ф2n.����Fk[��N�#YU3[�a���ϑ���^{�4]����u�e�h��c<�g^�&�����Å�A]^�>���> ����Q�ݮ5�g�.A���Ol�kxg7�7�L�|�����:杍]�zl>�i� ��3�RtD���ulN[n�v�6�hlʊ˪�:���Bs�-�m�zrd�{�-�B��Cy?���`�7n����!º���e��fu�p �r��p��{��	��7�gV@��[�,�cGIU��1�Wx�&��&�|W#�VC�Qp̦əGLk�\�}9��)��/�Ɔ�yX��ݑ�"��ۼ��N;+�`�oN�X�	�0z�f���wm��SK2���������7�{�m���{���z�O�LB� sq\��ZB�ݒh�:d�3ZjfnUU��@x�l�YD�V�(h��tî���3D���@�r�P�Sc����7��l���3Vk�4vk"�efv#Si�qq�*K���[��Rkm8�4���l0َ+��5�"��J��a]r���,cf�j�nƵ�Mj�K�å�K�%f��m%At�)�u�kvGCmO=u�?����S	�]���:�n�
:LMv4Pz�mB���9���z��|��!�__vG�[�n���t����cތ`�M�h�j�(�pX�v|:�<`�M��ˇU�r}v�D�qb�J|���GS�� �p�VGm�!�3�[����m����0y�R)��/l���#۬ ��]��.�;��h)��m�Aު��$�� �w�ppA���v���8 ��Q_�^�)oG��{u�G�7��?�&x�-���q����ce��5��<���3�m��z��n࿘]��X��U�(��3M�>0B7f�;���o �^���N�p�0p�8 �ݵ?$);c_*b��n��h0�KCiK(����N�h䴎�M��j�/[4�J8O!~v�����u��Ð�8 �$����o	Ȧ�\;���+�Zq=�Ήt93�G[�'�vəE�ʴ�2�e=3D4Ǻ�W����5�#PXj;jv-�n�"N���wU�?w���ъ���=%we�O�T�1�8���s;W���=�DS%�n4ǒ8������
��o~_�~����D��q�`�G'�ݬ��a|j�hH��p��ĕ��#1�!)��֮-��S��0C�Pכ:�A5��_�]\�ߤ�P>��i�ߝ�Yy݌$����1(�"��_V윊i5�HM���+��`��z��W��&^��i�Nym�2��I�V�eds+�s�;᫾^y3�,�3�L�����'�����r�9�e�l9�,�
&��z���	�tR���D�En��q0�q�Jڱ*Ö��uUs\z�$ɹp�9E�ؙ̲Y��+t7؍�F�2s6�b�s>�Um�|�B�E��̫!�,�2�Y4K �IE�$��ݕY'�����loQG�A��E�-NDЭ9�T]Z�n��뫩���܁=�������nݻv��۷ׁ[�5z���<��Z�~�&�Z�]�9ZB��=�_g	S��\RDn�5��N-��h���}C�ri8���9׊i��Ֆpf陈n��IԢ옷D�j��{�5Z$�S[�E7j��Aو�	W�F�">��704�bpraQP��7DgL��%�4��uL቙������Yb��q-qҶ��s�Ghź*�:�A��S��ļ�'〉sY;���Ȩ�eo#w��g4�ig�����$�z̠6\��f�eq�,v�t��XjZ��.�et�}$E^-ҫӷ����X������J���M�#R�/
�9,'27�1|�K#���j;R׍�Ő�R^����v�R�O��n��@��D��ד=Iw�h�CBX�L���1L�(�L���b>[Z^=}�>o���>ǥ5u<�����ʧc�}�n�E�8��}�GR���"��Qu����H�ْ&�����E�I�aմ8;�����73y]^z�԰\���N�X�33v�
���z�:�1�`�]^es�{
��wG5��1,δ��Ǩ�ԍ@���m���#ݢkq�)�]ͣA
��农aֻ�V��h�yz*�b���,rz'C�u�@E)yŕ��]c�lV�TC�Xw�S4#�X�禁���Uf6���w2,o&��V¥v*u��_��g�\h��6�7�Ӯ���p\�l�|��ppqȩ�Gz���䶳�E<�E���\�ҷ�`{:��
Q���J��<�*T�vW*�v�j������\t^��!��/�o����Y�����e������d5��G��Ţ������K;�ݳ6L��+��A4�Nq�$�79cPT�D`c.���4�N���s�	)m�ѓ����`�4��Hrᑀ�1	��HJB.t�\2�8a�R&�˒AGN��FC(�f�\AE�\�T1 �S(L�n��	���u���("D���J�p��$�)`e��� �#0�2(�#h1DFB2ȂPL�ɠL�k����D�A���v�d�I�L�䐓H�&a����Dh��Ȓh1)� AGwBLGf�.�ȆQ���B$(������$�-����aY+�_��2VQ88^�����"�Ãv��>n����"�9���ǌ5��n�>*����0�tkp ��gSv��V��מ�='��̮�d�h�3(�fQlɒ��~�<^�!bӇ�*ٸz=|�~�g�E�^�r.�?����܌x���)(f�slyI�$ �\��Yc��P��(�b�y.�_^�:[f�=e�O�=/�b �v��y����+'2��d:��hp��M��	�p�r�}�p��QE���ڻ��@�og2!�]&�U�x�3�a�ѭ��
����n��Z+�sG���̯>�e��s,�fU��ی����
b�"�IV�C�\�e��la�;�7�����3(�fS��絹�jr��T�[�K�A�gkR/�C�7J�̦=��rI�`�w��7����x!�rSͨ���M StȘ���{e�=/�3�#z^��=�����W���l@�Ȝ7��&�e2�U�T�H2Evy���½���<���l3:�̦��y�����9O4�Vz|u0����<$���k�[�%[W��4��9����x}��o~����^4hZ3WR]�D�[u��b\���-����zК1H̓���y}^~���(�p�6l�턏:嚫.��]cw�(:i�:Cm��&���zKAeÑ\��md87m�휊ȃ�A�v��gY� �v�6{tDsu,����� ���gdgkW.X4(p�w8p|l��Ǯ�@\�[Y%�N�V��s�
L�K�2�`����*�H�3Yn�� �v��n�:D�jh�}y��+Y��p�8p���p�|�ګ.�c�/�������"���C&P��р���u��WL#3*���e^����/��uy��c�:l�`ؑ�fPnt����}��fSfe�ƽ���k�Q�I޵}d<�n���5�:�n�/'L-��$'�5ph/i+��uu���l��'l��/fgJ�WdW�U^�����O����v�2�1C4� �k�<�Jͭvf�٠:[�(��ګu�SC�\�����5\�\a:�B����L�C0-��#���3��!!.�M�ss[k\f�`M��-�`eq��6.6,rZe�ճ<@�aT�\M
b�ɜ�!G��0-�-u�[��!c[*q	�lh���獫qn�c�؈VYR饬����7Ϗ�W���f#��b��	�Q��!�v�-˭vCk)U�R���>���Є���'߻1=���7l6�4�-\�"C��5�m�Z�T9>A�>y�B�_������j�����;T��4p��S���s�?�5k�����!�7y�E^0�.�����c��w'�U���*�C+!l̫H ݵ��1�v��F���Veᓞ�';��G�l��d!�a��e�;�4����A���v���I��us���Rq��|n�Ȩ�ۍjR��`i� ]�pA7l�{�mj����Ѷ����׾˫��C,n���+g"������a��Xǔ���r��(�evI�JBj�l��a6�E�dT%�l��Qi��I&�h��������Q���@h=�,�x�+)fXn���\쮔�
���BL� ݸr��vޟ+�'{!��e��R��a�n�΂'뺚�7�x��ʩw{�QK8v���;�����]���vBi{#�!��Yv���-N��3�2lT3��z7�,w���կ�����"�u���n� �0�aS:/%u��	������3�,�̰̮�G2�<��R;ƕpS��ndf�x��p���F��CG�W �ruk�_J�R`�fg'�����lN���獠��e��\6���/����秀Sc���]ہvؓ
�L���J�θѹ�Ѭ��&��X�m�v)N��c3����9"&d5�M����L<U�-�6h��X��	Zy?=U�޾o]��ןc:^�l����x���8���C�ej�ce��ݸ�$��Q��=k�����jz���-bA�xm6�]�nSHkm�`�m0{�]�@�����q��ڿ�~Db>;Ӥ�vU엒�j̢7=�����8|E�{7�)px��F��ڠk�Z5E朹`��t�c��݈rn��{���f)\`�������4��H�$=�6�����c�ԃ�~��r�n`gc�n�-�*����q��N�z���cw���jA �IT�m��E�����gS�TR�@�.�oo]���q��~��i�����@���������\ܰ�C�6Ƙ����,��2��0�BŃy��>/�RU	#���{'�(2B�^Nh��P�4�U��q�­�wo�,�1����n��cft��Z�耷���>w�R^5��!L�u�ڝ��z���wQ�͑=��k��a{�Ee+�^w���޻�����m�f��A~n����F��ێ<�{Գ7�����	�xD�
���6I����1?�V{�w���u�t�k�t��Pi�ɶ�}�8������]kUY�ШҴA�4)f��a�H��$�:�J>V칕���ߺH������cnɮ/�s���U��@��`�z3�~�������w�vO� ����\��`A���V���Z��u�s��1�� @SXX��bm31/m�צ��j�m�i��Lv�)�x��\B���)�jd��»a�H*HkNM[��-����˷[k2{'�g:����T����A��N��ʫ�~���V�T��K����G�dն�������s%����unc]�ݸ]�����4���[;c��O���l%��Pa�[93�,���l������f"���q�w���o]�ۧdB�=�nޫ73�z�oМ�4
��.�]�_�����lLdq�Q� �ɒ!Uz}3��IQ{BJ�����ߕ����p��}K{�R8BKa�t����R�� =v�8y�& ��Zg��3N�5�S�.)40BX#-��m�� �1�L�"%����l�ݚ��� 25�4�­��U�9���8�LB� ����L3B.��xo��M��ڵ��[�7�kX��r�����	�K���i�k�d���1k��֠���D�.��ڮ��Gv+��X���52S(�i2�<Xk]!�͟S����S�!�k5�c�Z�b[DT�u[G*V �+�����������Bl�����f����!����}1J1���cf5ݽ�\�F�F���m���`�4�l�7�g&o2��]��_0{�qm�f��Xay���� �I+��ݿ���S^���}�k�������&/�_�T�b���ܶ��l*�C���l7;i�\K��܆pWr�^+e�/��E�T�{�9�LC�L��K�|C�}gX��Oc��k�|s�.�;e��k�]�w^O<�ڦ��s\ϒ�l̴�j��͋1`;LV�l`�\��bl�Q�ు��o�)|��v��gu�����N�r�����bo���,Y��5r���M�?H�u��sc:��cz���)�|x?��q�n��5�ð�R�7�\�k�w]ڵ��"O�Pa�y-T^]T�	����@^7��M��q�����²�����R9��UW�
�H<�� 8���R�Q�]�w��8l��w"����!���uvz�:�v�f�e�M�n���,�T�1�Ժ�u���1
��E ��s�*�]`,";Mq,�F3���TJq���]�h��Az0D��.b��r�څMce�3���V��i���u�6�)��ܯ�l:���v�^��aN�6՜b���4ۑ4��v��ݎW��{���ڇ9EVsׯ����-c,Y3����~����c�Ws>�>�LURO?>�M����k����1�ʵ/��۾�:wG8�\iЕh���z ��1
q��˜��S]���F�F���a�.�G���P)��	A�	h�p��8<'�m�wovMeyME�it���w�s������mi�bv�Y�
E}���Zx�T�5�����UIH*���5	�Cp�q���̬�-c,Y���W ]����\�_�/�R0M�n�v��6c-��[�ف�ʍ%�����!�׍wov�_p�6&��h|vQл�-�F;���Bk���w�t�ש�3Rni��f6{1�5Ecc��p����{s�R�ܘ]ٚ��.��
uqṮ.�]���?�٨�;d,Y4�p���f�M7m����]��[˖��Eí��G����7nf�Gh|vQй�8�G��RQ�a��W�_�Z��)����U����#�����c 6r�5�����]�)p�IE��o�o�b��jP�6E_��������4~�2
�I��3>���t��j��Z�O�;f'V6ۜ��5ݿ����6�^�@��`�`;[�Y��m���ۥc�����͂d��Ձ1p�i�׸����$RC�۫~��{�WC����GE�I����\�Z�]�������R��`�.u>m��F��k�v��e��S�I�?�)�j���5_p��T��$��;ze��jE�jJ��uc`=��S�=wov�m���Yv�������ԡwtҌn�Jś��-.�l���ۗw"퇮���Z�șB�t���L'/��;e\��8]G:��[w��z��z��=�q�q�n<}cu��9��������yW�xn�d�I��Nf�n�I��M]IsRݫ��z�Ȧ�P�b�Ӳ���ݡ�h7s���8͢�.B�$4��z��x�Æ([�)������z���;�r��w[#_[���\3vv�2��
�RM���(V]p�V�˫W�SE9�;hn�n�3���P����ɛ�s����`��H� #��B�#Gu-$�%�RwTƁ����un�Ё[Vy�ʼ�˵��2�-��D���	�]�5�������_NǓ�j�y�Vgu��,�dݮ��Hd�p�ޡ��z�멊��@hc�Wvn=�
4�n8��m�AǶ��c�	].���,����������u_h퉱�[r"5b�dN��~eIf�m+�m3rW�������t�ۚ�Z.�FvmZ�cR��[�܄��+QC0���:�P�E�/ΎolX�!Z�������{F��֥���������a��<��R���R��Y(�f��9WO���(l� hW�+on�l�}�5�+����w�V����X���M���b�����r*T7��>5�e�E�2��\�0a��P�ERX!���7"-PnwJr�=Y�n�+���wgl�w����K g~{�9W��]�N|�sƶ���z0A�y�XSw�U�,̾�H[-�jC�����N�[8��FR���ک@ʫ�Hw]s5fJ-�=�CEy�sU��6{lA��t���N�1�[��8{�u7W�<f��n��d�>
�9eqhKCp��	I�v�������@%&�>�HB HCA�R}\cC&FRlCHd�I2��(ډ}���%e�3&dX( ̓2�$�L�H�$���͒#�A���,��R�ؒ(�M�,��9� 4��&�$$FbK��J23E2�jA1#4�$�DD*��&�L�4RFL̒I&�" B�)	2M���@�Ja]ܗus3*dW.������ ��!���)!Y2�d�EI��  �E�$FD�(�,f�ɌIhH�)�A��M @�P�$!��o�6/���׍��CK+\�30��qt��c3s��e��Ɇ;f̪¤Dy�,-�ڸ��i{Glvv��KB=M�Y����Ѳ�mKa���bD̤����f�ʠX��u!�`�b��Rme�n��Z�+Uom�5/��5��9�,,�o;A��6�k �t���ʳ`�%�z���*\K)���P����lL�J2ޯ;9����ĠY�c���sl6�Z�s!�ցYX\�bEu�X�L�j�+-�;��YZ�k�,i{%c�.4�`m���tL���͑���3V�*�C[����[nMj��m{]�� �YG�u�W,1�ؒ�)�b�\�6�,e� 6���K.Q�I���1*����5.+5ם�U�cp��-,�]Eh7&"�l�Ca����h�F���6��`$�iq&鶬��ˡh���0*�hj9���x�)2ꮼ-�MzƱ��w��B!3^��д��k��ReД۴�ME�X�Y��UVhҼ��,���W;+e�����-����]�ζa�H���8��WC0�����õ�6�D�֑�ڂcelu�*4h�SƀWl�74TX�"�ۮ�m��
s&�t����0:��d``
å&8�E(��0���\�� ���5h�1ɷ]6z��d���1�Dh�l�(`�J]�	��☖�&�1��FX�4�mD�����v�R�zČ

�]vٗe��P���LU����jj������Vm*����K�Lq��b���`b��u[c�Mr8ԍ�gDю��p�bgB�����7.�V�e)H�.GM\\�%	�1�ii�a�U�K�vױB�F
C;-n	kk�Ǐ����S95%�Z���.�a��5��-�$+�[]��5���A�2��4u�%��I��탎Ui�66��+5c 
܂8 Nc�GfL��B,�f�]c*e̷cX,1�9L�Mn�mvb�]l#M�(.a"V�v�����_���Ϸϳ�)
ZX�.�M/m�.�4&͘�Z�4l&g#e�Y��K(��k��eaHP,��֪��B����u��ø�1H�GT�v�1Z������q)�̺�J�b�\1Q�,G��]��M@��m�\�e�,��JJ�0���%&J�bWg���8j�%�Xؔ���3�83v�-��*�/A��A��2�e�]eee�� e�/����\p�T�ב8�͛B�-4,T3��5�ăF�Y���w4\������Ƿfe&e=�z;������V6�}���o-V�S�ܷ���z�߯�a��}����v�O%+{��h�PZVfh�n�qwO�����22[/���]ہwqЦz�m̙پ�$f#h�&A�S����~��j��A�!�z���V#)O�ښ�Wm>�3\j��{o�]Rl��~���`s���(әxɬ�2��Y����6��dc�ݍ��u��ҳ3@�a$Gs��k�b��f��]����a��OX�n��aEBUu�[՚.��*��\���R���X�M��`�y�Wo]�&o�=\w��"E��ݿxO0���>]������1>�vW3��L'�N��V_�9!�X�۫��F�7vU����̏��P��w�뿱_غ�u��/��m|��U��m̛�2m>k����e��@��~�f{՘��W-ɪ�q�y�8�U5g���.{������N���fnۛ܊u�ұf�S{����zͺt�ιJ�G�7��}I���kW=���G5���h�6���SR�i����n�]�ݜ��b�f�m<y&�����2����\�/��n�����h��o�ό��#� հ�m�ki��f��\ۂ�֘���X"�7��ߟ=i���mws�����x1!t�qj9�t�gѬ~_:�
�H}2�=�dW1��竲�V7�l��w=�i�:S��O�w���w��y����qv���v���aR6�(=6Ądǚ삂���M;�:^6N�
�)�I�/�W���GnZ�l�}�e��NՂ�󦠬�b�/x�9;��F5�z����N/Օj҉����3�-X޻��3xB��]B���Vޘs���L�ۖ,[둜>�RCR
����O��	@/���j��%Q��s�g��e7=�k]���#H��}*솘��� �C��m[!L7p�5s��"��a�+l�!Hi���o_�o���?�v���#;�M7:�99�¢�l������d�]����-'�ߙ�'������n��{g,]JŜ&޷��3�x��1g��g��h��UI$_��((�v���⮳9=���%.<�������wO0�y��.���
��<�Ȥv�y���-�����n����I���H;�.�!��,��o-�в�e6�;F�����4�K7��]�L�V��9�9:qmL�i�&�mJ�Xٍƒ���0��^kQ���;��O���I�ʒf����?-
}��]�!^�˛iX�|������w��fnfɺ�F�	j,� 8����1-v��h�.ƴP�g-X�uh�Hi�t)�����a�������z�cks��y�i�Λ��abк~?�z�A]I��
��v��j����oKT
��s�V��=[�6����0ŵ;�����1c�v�mRO�Td��n{� )��pl]O�+{{���������չ�H(�B`�p�Vt�X�~ڥ�SM��x�pUcˇ������#V��a�$�'+��s:��0�ָi��D]Z����������^����ܹ&YU��Z���<�1,[(� ��%,��4�q(5ɫ�!�u�ͣc.CՑ���7#�;tm<"s���|^	�«+nS:8�]Y8�3�Ա�ͺڀ�*��@Ų��g�����T�P����0��6��2TI�[��Z�R��6��Y��1b+���x���8v��8���qt�����$B��]���./�4lA��c���M����
��tiT���i]����-Q�B��ۊB&ŻeRWl4�V�%�*�¤ۚh՗.R��.��|��[W3��	���0Ɓ1%�B�q��Y+n��.���p�J��>���������RQ��,��VMT,Y��C�Ӻ�{aʟ1�v����������}ىF.:�ԟ���]�X�FuJΙ5��xtc����͊�##����e�V�*H} ��\��gB��~�N�_��.ȻJ��y��v�]��`�4��Wɵk�n��wn%neo?2��1�P�sXeBȦqݷV�]��]�mwh�1X_�fx���NN̮�q�������w�~�OO�_^}�XR9M	Ae�6%k,�L��t�K�SD	cqn-��N]`�&򅚻'j�у���Gl�#�sn���]Y��ݪ�v�D�z�l�z��}�=��Ղ!K�ɹSTc2��tW[&q�fټ5y�ΗU�r�K/�+�F������!V�}��'*bq����8ło-�}��y�Y[�9�lWS��C�)���qwϥ��tDtĹ��GwO���]�܁~ �9~w�=�qB7�<�,�x�]�F�Y����\�]�v�lF朚�������o
j�:ݷ-vֵ��,3of%̆���	�~)%�I�.���u�*ݢp'#^��s��Ӽ'�^zU�;�)����v2���?CE��a�jE����*�n3�6�]e���Е��Z� ��xn��{�����IT�*�j�H���]�f�Y��SJ�*]޳jc��z��z��o�$����k�9B$���d��4u�Z�#���,+�oD��������Ll9�1O�$�T�|�[t&��<_C��u����YH�y�2CS��ulT��|2/sb�H��bu��[EF���a�r�����Z�,�3W	M��	,fM��^!8��CҬ�]�W!�ߡ�W��&^8��c�8�� 3n'��+�҅���̈́nq�xtc��~�ޙ��q3*g<�޻��<Eݿ�ë�g޲��t�1��Iܸm�k��Gm��[��p.�L��-!陼5��%�n�74u(-�j�T���4��͗+DPulf��xl�1�ȋ��U������U���<�{�>齽5��:,����>^�IH?e��E3~�N0w�c�	�핰��3z{�Ἲ}v���61y��s;�Uw��H*L�'Mb���L���SMz�v��S]ۋ��ݱhv�1PĲ.�����w�M
�-f�>�,)WNm6uuC�B�@@��gJ%�cj��jj�qؽ�놘�*̱�J㎑g�o۽w��z���J�Q�Dg*G�r�s�wr�v�W�/��o�ERK`.�,зj�P�Uˣu�Q=�ҶB��i��_0�awv�U�zHg�b �H�&EMD�VD��,qD�vH8��5#������/G�\de����'x\t���dv_E����,
���-ڢ�E�T�Hk�?^g3�lK>���KkxG=��4*̵���mݝ��)�;}��J��l.���m���o�9k�#[j�.����/�퀻�p�5�6n�+��`(~����]��'4=��ZY:�{%��ˮio���N��z��]����6�Lvk���q�KGG5�x�̵����׻`.�xy����CB�,��������4,&o*��5=[�����%��M�1��́�1�h���	U�aYxlwL�c1��X�s�J�U�J47.�W��m�6�*R��ie*�%�dU, �����@U�uR�e���d9��l9�5٢�a��@#�	�F�n����Є]-LLYj�cN�1�Ս��%�c ake)Q��kq��)��j8$CD�CH@���b�&�q�K`e�7g��ݫ*�fpf��SGY�v:��q���KV^Δ���54�X��R����́�/�~��[fT>��hO&mSU.��I�����\tЫm�sls���kD�%Z�K���׿���/�v�b�f����k�i8�X�+�y� �_:�$�]��	|m���dD���� ����\ǖ��Y:�{${��%�P���J~�����x�I&U){D��]R�{w���Z�f�.�-f�(a��I$_~g�����V1]!�����7i�ڹ��v��x���§f��:ŵ�V��x]��wwm�R�����ha1:1�;�N�˓һ%��0��hxx��￼�>)�汤-mR���A�*�< ��#J�,_ji�Aʬ�v���u%X7LUFQ�J�bb3�
*%��1�ݫ�@�k�qv����歃:� ��M�y]"3�hn<Z����(R���a
|�@�{�=n9�p�`�)&�K�͙Ʒ:\�=T�xjRsI�l��X���y^�>�/�O�?{�#���5�S5��0�[���I���m�')�H�Y��ݡ��|�P�b�Ҹd��o]ۿ��z��8�D�� �|��6&�I7��߿T�x�e��g-�2�Y����J��}�f5z͸�o]�݉m��XlSֵ�0i��ı����UVc��;%ǯ�޻o�c8?��],���,�5&ݳ�ns�X͔�ŰR̊!��f[uڇ��<��w�Y������Ĩ��;q��q���=7�K�O;��;^S�qv�l'�l���z�Լ5[���op=�h�bĳ|�������S"z}�Pee9�c���M�zq���8�/�{����Y���"
���ju�+Oeʛ������"�M���s$!%��3}�����q\_=�ф��ף75���]o'��z�l����-uc�	�iL�Mm�ٽ�3i�s(�N���|s��f�E��3#��Vl��T'7o,�n>W���9n]fm��}�j�7B���,�op�eF�K��ٔc��AYF����W���r�e9��Ԫ��!�q贉�8�L���o�(���kxO�)��'ػ%���s,W_�%���ü�����^Ř�zI�1^�r}ҷ/�������Q���^�w!-V�D_;����k�T�����v����!r_WMR���n�
�ܾ|/&"�Nvr��(6ڼ���\���*Ǎ,�~�!6EC�K�ȱu��nsQu_ucL]����Ŝn��W����X�1���#6�>��<�ؾ��ňU��T�Z�2�:�oR@RX�At�Y�u�]|{:7��軾������Z�y�Ls�����M�+���zo�V�Z5,�� c,��\��>�0�j㼪a	me��Ͱ2��(�4���k�����c_c���. ����#�^mb]y�K%#��/1>����g�.7�`�]q�wt�a0^��k�<�+ ��tVb� �����E�۝��p}Vi�rR��A��T�8�I���O�K=W���`�mY�u�%��zv-���l�}��c���͑Q�k���&A|k^n�����fՉ�f��3��h���� ����ʮfh�a)H��(Ȕ��)���dȒ};�b`��k S�\���	�͈��FF��O��"lhQ��Ԥ���@ɒLj,b�j
`��H��a;���������ɢ�1&�l"5!d$��0D��d��Rh�b�X
�E�mJ4Ad�DPL�B�(�"" �j*6��)Ơ�#F�ج�J��4Y�T`ɰwq��jQY$h����F��V1	�Fɱ_z��HPhQ I�I�m��z�7ʫ��5�y���������҆��y���n��z�|����t�n�kY�'����mő,���������붻��A����ek��g#�h=�h�bĳT7m��x]�<�y��W�<��	�jY�,Ş ��&�:*h�*ARl�Wj0���x��2�cA��'�=��y��e�ݿ���[o���gUk�fC��c!ai{�]��T��qv�]�P�n����e��ަy�l�8�9j3����awoT��k�'l��[ m����=wp:��]n��-���:��7s����Rë\]���]ێ;]�ۍmr�4;�򮾟������s=�=��>:�;i��|}x�*�i������F����XF��}O�W�ݵ�6�o_eg�o'`jO^X�w2�H��<��dZ�����y��|ʻ�C6��]h�aݮ.���ݿ����vLX6q'���?!}����s��������V�Dڕ�Ҭ�"��p�x.u1F�D�B+Y�k��H��+����j��H�F�k�"1x�e��v�\���ms��b�a9���(��ـ,�z����m���J�7�=�䁖�q{��z�O�u��+���$9~�q��Y�c8�f?�7�N.��9O^(z����'-Ve��,;.�|.�]��g4c�C�SP�w0v�%r�x7\�Ά�U���,)'����/	�6�+���� .�]�{��+1��nt�=N���:Ⱦ����p�ϟ��p!����^������#��H63ww6tX�û�a&��ԧwU�wR��;Տ����V1N���gm�7��R��[�btx��f���IB��u`�7��V��KvH�s�+4 4]q1��kQ�h��KV,��KJJ;X����,h挤�u	K���u�i�q�-Eɥr�:oi�k�^G���T$`��ܠ�"ҭ�::�7+	k���I�d�����؆K`FG�0\��P&t�3�m�i�l���a��9���DJh��ʲ��](푍+����ء�6[���6a4ċ���~�|M���M�茲���Lk3��e�.th�[�ٷM�fX�����b�	�a���P�u�υ�,�ϲ:6kf[���7�7��A���S0�R{��o�wn*�2ٝf��ѣ1��������r�:ƱVfo��ov���aսt�<�w0l.��v��:�4�o�o'�\�R��]�ծ+�Y.��Gd�C�L��]��۷�.ڙ�_?H�٬Yya���S_��sV��[2�1�|�����I�I�v�u�ub�66X9c#S��Qk8WD��1�U��7���퇮�(Sdj{��LĜ��r�QJ��+�KWe��Q&e�����Bf�f3l�"�A�9=��m��z����Q|��<Z���k��!��Ǟ R֘_�7n.ǽ ��������Ft��g���E����Rɏ,Sz̒J��m��>�$�r-֝�E�Z4�۩��L��8b%�]�� ��
�'յۍ��-;z��ѳX�e����Wd{�N���[r�=0�i��H�$8�L��?#߿t���7��b��v����w�jARI}{${��sC
6�-kWk����y�1j{H�SS���s�M�M�|�����a�𻷻�[Z.`4�5�q�[��5���z���v����v�:����h��ڲ�hWk�uP�:��^�k�Z4��ծ�Fwc��||}S�/�]�o��)v��ҭv����������^��g�A$>��!�[���Vϳ�n��j���b-v������s�ýMrr�:���$���x$��l.ϯ��[�*v�z���X+�̼���Q�_	��]�{���֙��ܵ��#e"�E�ʄ�+O(ͨ�}g5G/mM�0^<�/2�P�!�2Mgq�&�����X���� �k�]�e�C�sK��Z����v�	�.���e���W���}��a[z�2b�n������
�zAR
�!-�]���ԇ�-Gr��rn#�5�e�w^�t�����fj���kz��\�""gfr��lX�l.#ciS+GMH
�Fѣ�v��ajWF����Λù8�`.��O�7�2U�eab:k�s�(=B�ߤ�P�2O��_�E�T�E�a"�걤��L�IƵ%��:��3��3|2[ݶ�y�;u/�D�,Rq�wwwv�"%�l��j}W��~Y�5�j�r���v����kvt0T�u��o]�i�׎捕x����7`�w�֊�"B���?~�)V���З�C�=�껕����]�&1�_&��5S��.{���R�����u'VkV�^����8N�
w �������zA�v��wcy���O�d�cp�2�`�+���K�wwu�OյS���p�H�/j8�R�i��]mT�u���C��$"mxb����Otcxm�ݸ�n���{\�~Y�5�7�#��E�ͱ���u}��$>�W� ,��բ3�o�۽)�)0�y��舽�̌1�]���k����ۺ��͗����쪃��RI��"���������&�I�}�c�f�d�m�����v�PLeé�^�m�u�w;����5]�\N6?>�w�S��v2Xu[ݵ�RC&���;m��3A��:x��C�:k��a�ws�w~�'��m����V%��峉��F^�9F
�K�����N^%\�,��2k���R�֮�B��M���|�h�5d��� ]�}�ߞz����@0��a	�F��h䖺����1���9f����cj����Ьh铔��-��hM��t �[zbe�K���Pf��iXŀ�]"0�sq3mT���7nŋE��=���.�M�B�3B\���bY���D��n°��։[��S]J�3V7;�:jڬ��s/��6XM�9���JĻAL�� n�MeI��cs�fP��׼I��'>��m�>�X���,�-��x&H�a[���,��n���`i���k#���=^�"�7n'�n�p0gl��y#���n��ܖ����.��E�1Ps��Eg��#��5�3��n.a��{�5�j�\��(��Y�����5�T�HjA�,|KIk���7e��6e�t�{��kz���
�?�;�X��4#U�)誒�&�ͼa��&1^b�)l�3��`����hI����(	0�L*����������A��\vf.a��{8u�j�oc�Z�mwo�@gއʱ.C�g�f$��"-�\� �LZ�����f�scֱB�JP�kL���u���]�mV���t�f[�U7�f���Ҳʬ�Ր�j� �^�&����x����vғ>�z��Y�1�A�	71֐�<2�� 3{�X�H�L����]ۛ.��mh�"�tl�\�*��]�����ku��0��c,Z0Z�{~��%�c9q6�j�^���]��]�+{�����}��e�o3����F�kd�w���X]�����FH��*~��bG�S�o]���w�u<�k���\�}ק�gB�W<Fu��k=ۇ�o?��ړ�R�����o?46Sc�ŋ3�~H+�.���]���@� ��ʬm�8�[i��[�b�Xɰ��� ��"�+�{�����]ہvԱVng1昨Ӛr^�ahX*��ڮ��#n��zn��m���whHel�o^���e���D��9�é��&�m���{;����	 ��س?Yi:K�P~{�ԬQ�#-�M��.�m�ƛ�bॊ�8�S�Q��]�4 �D�9W>J�w��.�8��;{s7�v��퀻lIhC�P2��m��?��/YVvv��h�Ӄr\*��s��Ԅ ����'�)zARC'�����Z�K��NԪ�3��}���.��v�w�>�|��o�}���y2\�/2m�9H7@uZ:�l$�!b����ż�e���߇���޵��][�z՝���-	b���n d��˜e��.��G��}�]R�B�n\��]}Y��Z:�j���ُ�>>�p�i�O�8�@u-��oW�ۋ��B�j�in���ͪL[=��oӒ���!�O�޻�wp;l��s)z��L�.�Ľ����w�Ǧ��nk/��h-��E��0�����Lz�N��P���\��^=Ý�,�Q�>�� ����>�S2���)����n��<�,^w>��\3�Õ�ȫav���Dd���p��^�^�k4tT8է)Oxvcַ��]�����@�z��u����m�z�&.ڛR7�6R�jf�¡���W�; �`��!��=���=�����턻�X���{qO���UWE���>��`���A�Oor��|kn�֚��}����3{f/*ř����]�1"_0�4�#���|ݶ�ܛ�ww"��*s�2��3;5�:A���S�ݘ��q�wov�)���	
oW��3X$�.�ק�u]nAÏ�_g�4��ӉX��x�U� �p�������xҦ�囎�
�^.�U�Y�Y������T��UU��Q��?��JIT_��E����]t��E��Q�Q��3[2�f�e��Ve�ͬ�l�l�Y��6�-fke�ٖ�-fkfZ̵�����[3[,��k3k2�f��l�l�Y�Y���Y�ٖ�-fkfZ̵�k3m2�Ym���[2�e��Y�ٖ�5fZ�5S-fmfkfj��̵��f�����Lf�f�f�e��n�2��Y�i�i�ieY�i��6�6�6�*��L��VY����k3m3m3lF*F*F =�}�� �*,b�����T�-1DX�QcE�E1AX�WtҢ��*�*��"��b�` `��
�F�EQi���(��,b��"�(�",`���"��P�����(�",b��� i��L0DX�cE�]6�,b������
,b(��"�(�
,b����,b(���̭��l�Y��-f[f(�7����Q�Ef��Y�ٖ�su�e��Y�Y��-fUL��k2�����`u�(�~ࠊ�������
���
��?��~� Ϗ��N��~��u���_�=�����Q�%u���}�|g���UE���y�B��[`*�+�����"柲/�����������}��}q���@+���L��C�	�_�x}r�>�(
�@Qd "0@�E�DXEbDX�Q)E�X�E��DX�E�1DX)E�E�AcQ�H*�#�>�����O���"�Ȣ) �H  ���+����� �9�|�@����������A����>_����t��>�?����?�����'���5�M� W�UE~G�̃����"���o  
�� ����A��q��#a���:O���}t��*�+>�?����O�*�+���g��}��_3�͇��B'�~����UTW������@��������PH�EΌ,�(6����ϧ��lS{��t������#0�Ͻ-�������}~�W䨠���L
��(������y���?�Rr��d�Md"��<�!f�A@��̟\�6|0                                      _  .�   
               P                  ���JPP ��!*(J�� PQ
AT���UQA*AB�%E) P�����B$*�R�� �D�P�H��@QT�
M��C��U�t��w :�D`u#�� dh�r �6@Ǩ�{�[� ]�:    /��h(�  �cO�� (��D�p = �4<@h()���� ���PW��s��w��J޽ ��{ �[��ݎ����h���  7���JH��)UP�
UU)J���)]���^� 裑�G�s`.���(W��r����R�-R��]�p ��IU�H����r2    > �:�}�xP6��t(	�IU^�Ҕ�[��(W��U+ݺ��V{W@Qxxp m�R�{׹T���E�
    =��P*���$�R�(*J@;� ww ��{����:���x�J�:݀�@���=P4��:�R%n�2 �    � ��` I�:R:�����@堠d� ܩ@�
7w
(�N�@�� �  <  �A*�
T�$"�*�7s�(ݎ�2���wD�V m`NZ ��ҝۢ�J��VZ 7g@   
��  ��gР����U0 �v���w` ��� Hr n�C�� r��@    =J���U$ D	< ����n`��Ί"��Ѷ�����0wS��d�I%�%w W��H(w���   /|  .��D����a��Es�
��������n��G���Tr�WE۩��
���%�����5O�I�*��h�A�~�%)P  �ʩI�L����R���`4�OT�ji�@  3PI���JI�5  O��W���G���I?������
;����M�[�I����I3Vy�$ �y$���$ �~�O��I@!$$?\�������W�֫�[年*%�n�c�-�'OR�Y�!�M�Yݲ�y��<�ɘZ�fīҲ�^�CN����	4�J�1��]�`ٶ6�n���4�%�d�jku�ExTӫ%�"j����em	Yck��EF�k�+b
�=������E��i�̱�j�nk�a\w��3��T����N���G*!�Pa�u��5S�*n+�P�^:بA܍�{�2𭽴�UHV}Gr�Ŋ�{�Pݫ�o���m\��i�-��-÷�y�*S-��ͭԬD`�x�]Te/��s#(��ݻ�ZpjU軋!.JѰͦQY�v�3ov���o
���"1m�����+-�Sr�Л�4]K;��܄mК��`5�C��vA	̧�t�PM��,���fӪʧ2b@�ܼ9z�e)��I��-X�٬�fJJ���+l�
<R��Y�KƉ�.�bɗy�w`턓u����fU�h,k.��Zf�b]���f8��u�n��zt��Z��@�p�i���(m��v!c v%G{�S+c5w�ܫCf,�5D�n[ٷo#6�Æ�Wr���ż�ʫ���pn�V�ɛ���L��ջ%�CqGkXz�U��Mfƥ��D]*j�j�֔a�T�Fɏ5�Y�c5���^��ىcf���w�)Ry��(��`��Y1�ӫ̧Y����Δb��nm��b�t�7p-��J̭�s`˗�`��n�3�s�4�ـV��gU�����{��¨�h�(̚�2��j���W�0��{{kb��]���Q�x��vɛ�%�'j�#6��yv�!�#wuu-S�;���m]݇W1-fn��#P�p�pe]��8�C�%]FE�����nh*ݳ�4��F]S�����L5kt�7Q]h�����6��f�o0�;a�Y�k���N�)���o��363[T���0�W�6A���%@�35�HP�]26ܫ�%f]XL)L%S�Z��ڬLX���[4���'.;зqVY�Wj�M��%��B�'`�!<Dūh] v"�-�*�){q-S3,�d���Lm���[�V�L�e�����͘�]S���Wa�)W��Zf���e�<wH��D�ʤnM��O7M���4-쬨�%���e\כ�Cx�i�ۻ�z+,�B�Pj�+7��n�-�Y-+5k�%H��L"�ղ��{���Jg1Bj򨽭WfY�.n[�6-�n�n�%����j�n-{�wbH�8�mY���Z)2r�V�	&�Z������N�
�*����Yf��r�e�[��*�J�2�Ɨ�nRW�����4r�^Z���H�LAoB��1�z�Y�l�ܹ��j�^#r���01)f����v��ؠLh�L:��R�ۙl�8�U7j�:j��^�XJ�P�RÚ�.L�܉�j[�U{�i��*:�+�«���V�;l]�N��{P�`�)	a�/h���ۣU�f
�w�^#lMcJ;��&�q�%lA�ߩ6��P���-��z(Lr�pr�~�`tsi�iٺI��]����7omZ�
�\���,ӱ�aF�흆���-3X���C*�VH/&��̫��/ zU�v��T����TZ��&[;�]�+j+̡E�X���T�;���ׁ�� ⍌�y�C*[�3.]����CJ�#R�uRv�X��kb��쳘h�н��	���3MM��:cؚ�����H�f���p����!�V����n�.�'.C,�2��Xշ���vt�Ҥ��,"kr਴G2��ӂ�$+ۍ[��h��l�UQ�ʬ�n��kM�R���˗���"�B��V�f���.C�X�!5��j���
D��v��!0�J��ʸl��d�Y冥��f`ݯ�]]���́��+�WWy�e�4�����A��)��^�e��ĉ`�R��
v+H�:v�PWb7J����bh�J۵vj�'��5�����$<�bw�-)���I��.�Ve`yt��ӌ��ś�U���o��6&r�e��O/oh�ū��ZV�Щ�ƨ��w��1P��l����R�W�H�ˠ�߶e�	r��a�w���d��0�ˏE`�*��whY�I�j��K*��ѻ	�c�M[۵����Kf���]m���s�ܣ�PPU��*�ݑch)�qɇV�h�C2�3HÛ0����I\�������-��m��t���ѹ���[v�*|e�
�,��F5�d�7dY��5;ܘ���7���m��%�xb9xSŸ^F���YXnM	��-�uy*�ٴ���-aѻX#(e��+]b0��9WH`Al�v�ܢ��ZuCQ4��J]m�v��T,`�H'�Ӳn�wZB���u�ma%lݘ.b/��R-��Y[�Mѫ���{[%R���jǸNʧz��ܭӧ;L�VU��B���ӺT��I�t�TZ�z�MQ"�B�-�Xu 9[Bsl��Zv���҈f�]��Br��X�qҺY#�?!+4l�wR��/0�a�6YK+(�=�A[b	x���3r��;�<�mZ����j-i���E�V�
�q��W�R�Ӳ��,f�Åd�˷����aW++)�P�
�Z�Q��
Ѩ*��V��v��C�Õ��zU ��Eml��l�,M��F�u����nf�h�v.��b��1�WI�X�ꙅ\�
�E�TJ������vR�QLg��	��lf:g�Z�WD��	�Q�� �mٳ[	J��]f�[�!xK�W���$����H�i'L�+	�$*�u����s���a.�Qg4TC+o\�ɽ�Y�a�i�����iQ�:�+M��̶7���zp�yY4��(�n�͈��`a.D��Z�p�x^��3n�m�p>4�u��bKZ�z*��>C6���Ǖ��2�����3Oe�4e�e�-���F`�W����I��M��n��X�.��d�/�ׯ�1�J�@��L���b�,:U�mg�mHX[��5I��i"�
;�(���A��;��j����a%U#x��T�v��<#j^��%`�tN���ڊ��˼�q��yf���S���陆m�s-h����bݣ[�i0M�cW����ۺ��j�Z�{Ҷl�;V��-�#M�L��]"��R�9��`Ӛ�'Y���g+7�V������tol⦈d\pZu\��m��{b�õ�Ys20'Z3f�-�v�%��7�Qw��`��5�F�.I�2�]���ѡ�F���-�4��S+����1j2T�]i��3n�0��͐��ɚ�*U<���h_I7^���&�bY#5������R�1]���g�f5�m�/����saYt��4&�m��u��E����/r5wZ^�5����L��.�Y';�ZD7�g��'u��0���v�b�nfQ�FN���tTVWո*K��<�H�p[�F�I7�F[{X�9�L��(���W/hcyzfIj��̈́���69��+҆%Kf���}6�#�YE�0���̱3j�F������T�)�URy�u���'��ג�N];-�Dv�Rn�{#��7cLG+�d,nb��e����7hʒ�L؃�R�ދ�A,��b�U	����B]*�QplȮŜYn��(���Ug��8F���dEj;��kie�zC�v�%4P�"��kkE�Nv�&��^AE�TɻH�fݑ���t�i�.^b�V�U6~�ŉh<��~9��ܰ��m�J`��c�A�%�.ĭ$<�ѧs&.Fi�,��Wz�Ƭ�[u��,Exv�WՐ�T�(����Y�1�ڦu:�[�f��Q��V=:eP�a��2+�q��;2��1m�V���
���V�Kv�/m�ɕ�*j׀�����H�C�y%}���V6(��m�U/%j�b��7[G�u�R�Q�ƪfX6�,2��EV�����n#{��h֞��/j��h4H"����J�;��[j`�+Eԭq�M�E1B��cxMc�)��JJuV�ʳ���c�6�6ѹvAڧiYŧ,ͼs6�ʻa-�M�JM�
���l�5��x*�@�Sp�.:�t\W��f��,^ԅ��r�T�r�ha̻U{H�c&�n�i���Ӆ1+(�����J�U���X��U��Օ.���B���N��9Zqa��7M�7Vse��Ď(�ݻ���{�S��1�c(^Į�	�b��.l�w�\�q}(� ڗZQv3�v��Ge��n;q�ދ�m�v]�
��l��l�ݱWe�����[�NQW�H�ۧʆ�+�k.����:Ż�Kq7%�Iy�h̸�M�bV���
;-�ub4��z�-z���m�Xlʨ�+iڙ��W���v-Yn�yW�,��.�`��Ǫ0��mZ�k$�:�Vi�t���U1D7�Um�2��m���Β0�"��T���V'��KC �Q�f7��86$�\�F�f�U4��i��F�w_�=2��z��������a��T;UQE��V���uuBӲ�b���R���e�W�j�2}��i^��IcBaʗ�W�W&:ȯ˷��z��jiJ�M����ä+]�%<���,�5�Y��MgQ�u-i�q@�k�яҐ�э�2#YY.'��8w6ѳu�]:���9�Q�iclܫ�����3`_=��zs5�9�r,KY�N4.�����E��#�)b��֊������٩y.�]�,�	��L�i�o �B���N�%��P(U�K02�k���W�\�\IVS;N��#E���JW���׊���L�:k]�Ǝ^Ԡ��:�YV�<�N�O�]�˭�����Z�UYu��ȁ��4(Ʃ���sX6���hSʤo(eV�cԨ-Z����v�c-mk�jm��7v�jC[�N)���.e��ɓ�3m�o3.&�{5^c��®]Ŏ��v��tƬڊ*�����S��b{Q0���[Tr�f��a��yU��m�3pY��jmKLXnJ�.��W�m�z*�7��m�7J�0���!�Zv�e�$�TV�T�w!��f�wF�ұ{h<���6]ҋ6����P`�S��t��M������Fd�10�I(J�;�A�*�m�,�:�5E��vEҹ	����,�Ҭ�-��9 k,"�ܑ`�ӑ]�� E(�0P!�	�+F'@���Zʳ���bƱŅ���'�����w/I���j���X˂i��9xb�1ne����h%��V�ɏ
#r�.VD`ڥj��n�Q8�e��i�e�ʹ%�n�+U�D�|���ӗ��j���slS	�tݪe��JȾ�jOR؃�ا�q�{0:7u�)f٧X^K%�o�Ya&��{�Mt&XGD��X KFH.�h��S�1�Є�qL�N�ں��Sw35:\�UG8�;��,��q�p�5�5��f.�è��b��[.f�E]��K���*�]��ȕ�F�t���sd��B����VFզ��#i����]9���T�љ4�]�Е-"�S ���ϱ=���׵ oB�
�^�4ɑ�z卥{�Ɨt�,�ܵY�mc���$�Gb7K��{[�G9^G,e)�u^\7P"�7��]�����/�0Ǵ�����ޭ)��L�6(&!���N�kn��.��n���jejZ�n����L�I�]��]	Z�bCU�$����L������]�r�J����5��m�M���M�1 �T6�(\Y�P9�T.�r��Wy���*��A7D4�f��d��m�Xde���Y�U�ղ�f���i�8�Y��y�<�i]ᰖ;ų,4���tt(�ehn����n�E�'ZИv��śY�w�aH�feI�VnK��bR�7u�7C.�'��;���oE��z�ǻ�CU/
���5�F-��h�ʑJ,􁛐+�+�3�w�v)ǒ�Y�$�+M:��A��tҽi�nX��W�D&К�5�n�S��[�w�ۻfV����۔l��*���MتfůL���]�:�{�I|0b��5�م:�r�Κʎ�ͽ� ���ѵ��0�����Ya{N�`W���ݰ���R�k-^�
����kE�zɼk��`��;Ò+��X��+,oB4�dTܡ�lї1UY��GD����jVӏ"�c.H�#���\��G2�~��]�HԪ�n+�ȘKr��i�Y^�[���/qd��h�^��jĵk��w�.�]���p���F�t�Y�:�,c�a�U�f���Um�NTqM^:Ů�*�`�"�ޔuf�{��kaɦ:ڹ0&f]�ځ�Y�/
e�U�֩-��g���f���ڱ��n��WX3nZ��E=���//571,v��ѷ�6�X�gk\ͽ�'�"PHdG
�v´2���1/C.^]�th�w3s/��,EI���[��Q��	��{���й�qC�S�"�Fϩht�n\2k��sn5���^,�"؅,�i��M��7v�H��uv�Xv��jm��*�r΅�����U�t�ޝY�^�u"��ޘ��N�sVln�L5a����h�}=֯6GK5�
{��*�UQ��B����X�q�xƝ�v�K�{���FKn��I�^,l���ةZ*E��DԔOFYc3W�`�z��Ī��3mb^x��e�y�%�zrƦ�����5�<n�ڻ�OQ�3C� /\����Ǹ��&I��k
�w��Y
u1�b�2e1*�R{o`���%ۭt�F-��k�e͖RW�w{Y/t�3�ie���U�3wi�^dM����U�hY�B�ͅ�75�6��"���MS4R��0�ڕ&8�\�$�|Y��|��x���fř���乗KX�ܪ�D[�ƅ8��B�J�̻�ZwRI��w�CR�=w_3��QٗC(fҲ�
w�;y-�%&2j*T	[4�;�2���H]}c�i�D*�ʨ�j�e ��[��CglB��抦�
r���0�H��`��!��[���ܪ�쫴�w(��6���-Ӎ%�Y{�0��mK?:y4�i]�+q���Upi���nwY`���Cv�:UU�:f��
�5mf:����u�d�/P���SpI��;�;�!ł���*���@:�a �,��QEj���Uklj�ŭcmcZ���mQ��
�Q���m-kk�m��cZƴkQlm�6�5m�j�m�Ƭm�-�bت������U��V�XѭlZ�m���Ս�X�V���m�m�6�bն6֋m���ѫm���Q�k��Z�[[��մZ�m��m�U�Z��F�j-Z�mj��Z�j6�Z-�ŵ�����E���Em�Z�ՋQkZ+V-�lkU5��ƶ�mU��h�գm�j�5Z-Z�E�Y5��Ċ��	!!�$ �W��Z�k�O���.8s����1�sN��pA��I)����M��pn[���6�'v�|~��x�xh\�hU�Yf��S
�]�;��vSKo�^�a�*\�F���U�֞��m+R]
��x���4TS�!\(��mC ]]^�˗z�ڳ�n�2��w�j�n���5�g��j�t�۽9҅���U�!�-ś8v:w���VY�U\�f J���jaǆ��!���8�;�Z��Ӫ���j�ۚ����cw:N*�Ϫ���0Uj�����Li��]Աe<+����-m:��ܗ'N^�zqg$�������1�v��K$�#��2����擖k��q^���\���`ØEi춄�v3��&�w��m�psr���W��{��33S�N�ʔ�l5�A� ��7�~��O�\ĩ�+�n�p�vB�]��p=���[�C�u򧔆�X]hL�q3|���u�`̪ڍ�W���9X�*/�������o.�ܩ\QWt��9x�VbX/��.�xUL����j��W.�-�8B��ïH�yO+)�K)��G���QSյ���n�WN�����ZchR���t.p}��%^>P򚬓*��I�tkw�ժ��[B�]�[�k|y*�\��f����׹|�e�4n,6�Z�J��7����W�MW��8�{��$���B�1`�T_nt1�/�gUG����+�P��#v�a|򆶭��T�s���lgo_Vu���օ1�ͧ����gf��vb&��_R���b�nfN4�m4���X�)�.�����T7`�;r�����3i��6&X�v����0�Q,W��>�ӓ*��ц߬����=�WSI%����T�Nbw��_fU�.0�j��F����}��;���T{j�Mwpk:�	W��z��im���Z�+��C�����R#�/��~�(�.�s�yZo.Z�Ҝ�un;(H�1J��W��������b �w�gE��9�vyi��L�к��L�̃u��f�u�]��CZ1ꔯ�t�78�V��TMD6 j�����p��b���/�N�a�v�mn���T�c���X����<U��+x[;݊�s1B�o�]J_"l�����f�c#2�3.��uMè����%�ug���b0��+�W�&��S�1P�s$��%�Y\E]�]���3� ]80�wV\|.�}�K��h^S��z]CQ:�"u�=����]�[3b�nR�԰:#�˴�
�:����Z}����-.9��^�y�r���=���O�l���l�
�/l����X��٪���rм��]�w��N�lp��!��^V���4��M�҃�fUS�ۃ3wE�j���f��N�ً5F��8��n�W\ݭ�֤�V������g��r����]��Ś%ɝ�/�n��	um�if�D�N۰�BB�ɛ�T�j�}3]��&1}Ӗ��f!ʮ�v5G呃Pm>i��mnV��Zj�mQ,r��p�ʵ�Y�ci��IfiH�s�&�f�V�|6�ռ�W�L��P���)=�����|wj�٪���ko����t�ɶ�7pS�d貣��M/i3%R��AmK��ʑ��;�dgFe<�_��X��.��N�������{�wUnn񚲐�h��B�_f$�iiB�����mi4��YCgMś�.�+���R�gf.?e�YTyՊ����4�EW2Rc���W].u8��Kh-�j޵��B��0e�p�-ROu2�&tL�������ݻ=6�>g�+�y�7� �MyjK�Xweb���l.�Kkk)kt�SL&��<��X��BvlZGs��b���c��+����Yv�/��G5ݐrPk5J�m�9�tU��=�Zc���h"a\j+������8�冹[�lO*���:2�:�$/(�}J�T-�Tzn�}YƮcb�����k��^ns��On���$8��΄e�}��Zͭ���6o�W	�H��B�fDUJ9Ck)f8���&��3x�Y�EZ�+*�t�uV���)RH�ׯYoy@��!�Eo;���������)�œS�nu��ڄ"���i���lF�Q�Ν�.�k���u�7)Qi��gf���Cr����>p��S���f[ګ��,�C�uᕊ�}o�3+���v����s�WEӕeTg�r�F�fE_׻�ѐ��\*�����n�O�T���&�SQ&6����ኖ�j	�����kr�*;8�s%h�N�(@��W�d)6B/6Ӡ{�v.����lڙ��:X0�;��n���]-�iOkO:��`��2���7j4K;�T�r}7x�wq��n�u���v�z�̈́\X�+�ٙT�)L\�.嫼�{�F����@�ԭڣHn����Tw-����W�J�6½#j��h�wR����.��ҎW,��&�S��m-U&a��t��m^j��O/Zo�f��٣�J&O���U̱�Yҁ�u]U�2B�Vm̮����p����5F1)�*���ή�ւ��
�؝U-��f�YM�5*��\�;��:���T�uԹ��a=Ͷ���Ǐd�VCo���l�2�V�f���5M<��<�ޘ��÷�r^P��w�m廨�m�vf`{��u�+TE����ZA��zx��=��JeV�_�h+4��g\��vv���N�ǔ~�KI�J�;�8�*��>2]�Z�N�m"#���k�\��;˸��j��v�S��o:"�.�w;��hb�7[��]x��54�ɳ�s^X�l_^mR5���[W:�/��qo�wγ���Y5+��6_V��^�5R����>k��,��R.J�6�)I��5>��]�
ŋ�{�z+U�u9�ŕq=�j�|�v��k{4����9U�ժ���oC�U9L�G��ԡ�@��Bx����o5�o[���:�2"�1,gT�1U�w�Y�ViV�5.��.=�,�����.�3wx�5�fnWs͜ޅ�dy�.�͛zc㶙:H�c7k{qX�U�Ù��Y���kkze6璥�&�{[u���b�����ŋZ���5�qi��C0[�Q��K�i��6�\ut�k�M�o&/�ԨoFдx5�h�}�-�i��FhM�T/�{خ�#��T�;ںT�ַ�SQ5Յf����s.nv�t�4K��+7�o����Ϊ�e�"�&�^q�3������-ޱ�l��6�oC*{��_mo�Z�+�I`;i��>䪉��B(�f�[=�Wu)��"�)-雧����QU�������X7L-vR�g^k��AN��65Be�u�f�e�yye�i�t��:7��[X�Z�Xc�������1c��S�Jд�]�X���\�ӡa���`���р��l%��n����m�Һ��츭����8�8��|�^3�c�,퀥�o��y���S/.��qvU�ML�y��;kf�r�u�t����cn�b�cnAg�d��ͪ�����^���WS
���C���FY��A<쯒"b�ʂ�;d�x��,Vk�u�2���:��V:��+/%|��+�_1u�&�-�39���\��񉅤�SE:�c��5w�s�ũ�a�ʭ�5enU�ۚh��w�8�x��0�����^bQ8�6��6�e�0���ȼvm�z�KI`�z2b7%����U,8�����Җ}�Q�)�x=dU%Y+�+MQ;ۈ������k;G�Nj��/��-����t*����\ D��=z�."���ՓQם���`�z~9���3x��d���t���ʫ�P;{4R}��.T��vM�4c�ު�*��mr�]
·P��M]�1��D^ݖL�4�mf^dZ�\�My5�j���
�YVuL�AT�6�^��y}T����/UT낻(���w�-��60���������2��\Gc�8��*������ğ�΅��x�]f杆��]�(Wb7nѲV;E�T�0�V�D{�Ӕ	},>��M.t�&n�9�����S�j�2b�X�E�q-���#�BD�\7q������31�[G���zWwMe䭙|�u���!�t�s˱H�S0M�A���]]��s�$�m��&�`�l3��f�a���9B��:<�/��mSJ�,�ARz�Γ`b��te�<�.\��M>�i��.,4/dGݺ�0MO]\B�[�����X�ۛ�IJ�m�L�زT�n�4�:_of��4�،�+Wq�ӗu��s3��v*P��H�^Rٙ\�jko]��3n�8��+WLᄮ)��V/���*pӀ���L��P�+��u}Z��E�p�Ρ���p�Zy��w5�X�X�Ys�o9 �1ӳ��-ԟJW]�[U����C�y+3�l�U[�����ɍ,�¶gU�ͅf2���7���yuN�������f*i��U�w�z��s�g��d�]jMJ�[#�؂�q���c��q������e���`ʷ���2��Pj�K+!��<�Yb��U/:�}#S�s]��uWmT�C2ʽ�s����7�u�T.���*��a}mvo\�Yt�N��+*��+sDV9Z��!Ü���wlpp���ՅU�=��):�� ��}Z�{��y���q���B��@�wV�ϸgf,���.���.D�P�NU��g{bܴ��*�͛���ӗ9���u����v%�8��v��N�We�p�7Հ��[B����V�Ց\R�졁�բ��2�pnZ�����>��+%_X��0��P��/�e�b�}�v �K�S�]m�����[������zΎ�Tv�ە�(����v�"ѓ�V�V�V�֊����U�GQ�Sf�"�nKo	���}�rѧr��;����u���:��]��`�׏eb�x�	�fg$�
Z2U	���%�NU����u#��jͬ� e!}�r�nb'v���W���驟)��`�Ɵ	�_�vu��1뽪=}�
uV1+ۍf�	*sl��v�or�]x�*��<�ޤ�r�܁��Վ|�R����-�j�V����г(XD���ݻ��:H�m-C��'LJ����s�j�1q!��8n��P��db����-=h+s�PΣSx��i�x�,���=7.�����!�*cύ�ڤB۽�����c��/V�lsv;h��i?�9J�̍(��\�������i�ܡ{g몾�8���Ed��r�O3�;�.��17��ƩJ`�5�z�6��M��۪��mou<�jXܫ�$Z��vV�P���-c=��nl���j=U0���}�.�"9�aU���ـ�����A�ZIr�a۹]nV���?b<�J���R��ֆM_Uf:�LW-�����3jqqe���J�7���U���6�����ʹe�}��y����#X��[��I���Bw`��t�}�Q���5S���@���}��١ѻ}����)s��y�r�y17i�^��i�Z0�.p�x��C���Y�!��XE��բ�%�z��w�����?f�5WƕG�gP;�������흾NK[����l�9�z��=���P���8�QQpb��KefU�p��0f]ޡ��κ�s�S���۱۝�Xû�lN9}��Qs��ٸF�^$�W��k�Sզ5�O��'.�c���=+b.�;�i޾L�;�&,�N��t��6����א�Ц8��5-&��]�;���r'�4M1���`�w�q���B�OL�y�u�]*���&�r��#LR=��I�5���Ԅf�5l��]u�f�mm�ٖ�j�c5��� ܊��e[�7
z/Y�@tB�ʰ�W}���=g cqwz��+���E��ˡ��t��/�^)]n�
��r�1�����<�WZ�]*ܬ[/Ov��[
���ܫ�+�8�w.���;�o�Io�x�gZ�wl��L&B�p�uT��w�MT�%�<ouPcc2�Az/w���}��zLyO{_U�N�寃X��oQU����UYY���oԝ�n��,t.���J��Y1P��w]����2��8����U{ˉ�*�S,Y2��v_r�{;����?H�s�_4j<W<;�[��V�j��	C�K7��W��E�>�77�ryM]�M6�m_Kw,�X�]H���Z�����ݚv��c�	
T,mQ\u��T��WWW[Dp����YB�w�OT�t�b�����*mr}��{o]��(e,������Y�Dz�*�e��6��ʧ�fml>Yj���1`�dwk Z+Z�y��b�Nу{ֳ�>�a���ڒ���=}
���Q疺�mn�j�����ڃ�XpUV�;��;P�r��n�2M�9��l3'uA;��Qyxld�7n�(�n
�q-���:++8��ܟ�N��Rj�7v��7d��uM�,��ωs>e�ހ�apƕ�K�N,�������uFZ{�q�cqP��nj�UF[���A�2x�f�ޟ:�Z
ㇾ��1��T6V���U`�ظ�o]4v��m�4�W�l^@U�ͻ�%V�æ��Q���(�A�;;:�f�T2��.,�����������݊�H�]2;i�5�����|��R���$6���Cyb��gO�lb�->��n���u��=�ݜ_W��Z��k��	7������T�v�B^f�Wje#�{Vg��*ПSJ�oZC�1��c&��`y)�YC��੔�*W>s�޴�j�U��1���]�7N�.)(3nXN�܈Qu�r�Vf��Ў��Ve�9�����(Q���y�<hɄ�K�l��}g���ܗ��V���%����W���=+u���刪�z�'����/;]�i��er��5o*}x7�=���[���Z�E�YI��wgE�(+��z��u2�w�ݵ_T�J����i���Ǝ���+��5V��n�wsn^�T0h�t��62��0S�X�ө��N�5v�ޒn�����)��|�];��1�cr��n����d��k�6k�W+;7�9�*�T�oE�	z]i�v�S��3�BKpL�߅J(��WuU����7�{�kۚ��u�����s�<Sj"�S�k
�����<�ݻ���y��I, ��F��N���Fkv��������؋�ev��;\�L�;��1����sl��N:�:��v��٩5�x�ָ��� �1�3����֨�l�u%)�Z�;Jk�Kf�x����m`�R+TU�jciL�]K�K�c+q� �s�Kq�m&���=�X[��Eg����� AN�iA2iv�X+Y*L)W0�})�;i2�=s\׈{;^��pn[&�x�6����ٱ�1`�h^YF�1Mk2�f9�Ý�Sa.rY��� ���㎺b�Ж�����x����s�I�V.�p��<!�o��|N�����㇮m	�v2�]���WTmX���bd� +�*v��$��|�8۳�z�\���m������B$��n���T�t�x��ݔ�pm��m� ������Tt���gpk���n�[	jS$O�5�#� �֪�Or�$�g�,)�F���r����u����^z�N�ql�덥����@�[�����:ԕB+��=i�޺��{v8Ř�qŮ���	�b�����Zc��	q��MRSP���a6��uL7WNz4�콸��h:�L�[��NLp���n�71V,l6AZ�JL��φNK
����h�nv7���5+��]ZN{�x��3�Z^m�ꌔ"���&�i�w�فx�O=lkc�ƩLɥyCF�kAU�!�([UL��\�����e�� ���.�Q�	�͑�cPkv�*suv�Fn�a�&�����yԞM�M�Uɸ�Ĭ�d5�Q���$�m��c�1ѓU�KÃ'aqB^���Ki��JrAi��t�)�f۵Ñ1[�46��csn�ֺ���+��]\���3��9��{{&��jὣ���aָM�ƬN���ֻq�F9�:��CsUJK�0�CƌЕ�)s��^��Ld��SMY�(Is�(���2v6_`�/��fX��`!����r�÷ǧ�j��>�������e�ȕ[v8�l��r���wYMIz��,[q�$qim��h��b���.�vt��z�G]�����Q��!�����b�c�Wn٪:6ֺ��^^��������&�fE�YC���Ż]Yy3�u��v�ς�6��ù7G��+1H��"���ՠv��e�ȱ�[�U�ɜ��c9���Hd:�[ۗ-��� j1zs�z��t<�s#�fU K��n��ٱ���Ԥѹ���`X��i�prt��Z�[���p�B��TW[P%Y��bX1v9'mX�;��Y�6#���&^��h�[�Qt�3Ms��-�K�֎c5��ll�h�8�'n��֜���Y��\�=�S���B[�gt�[i����Mlm<v�.��v�c�'�O`���i�y9�d��p��v����v��+z��;h.��ϔ|~N�0N�=a�ʽ�����[�h���1ćFٛvضR[�%��xB��{�n���]��U�,�S������T���u������vCv;:Y�P��n/<���7\mt"�%^y�˲��}ݐ���K�X�Z�!�:�iH���6�n��#v��!�n�gټC�d���{^.2�n�#�x�v!_0��M�0gE�U�hz7Q��YwP��{W�8��P�<��b�ūL緬-q��cqˌ*u�y�݊y�����y�y]��'��+rK�h�0�f���[�bǄm�`ԣ*0�m��횃,���8�wT�rZѽ�p4c,��4��bz��*�`��nخ��sѮ��ڮ�K�fpt�^۲緈cf�&��|���Qlp)�kաm�tg�ӂ�s�}sv��iV���z�y�-�"m�X�ym����r�.��e���M�6������P�6Ӏ9��
"r��/e��6�ᮨ�6��aFY�5��4m4-%��i�eR�`(�=��^_Y�\��F�R�N�3]5���EBR�/"%`�w+36��hd�;Z�b�v�5�^����5<>.xs���۫�9N}�J͎�U��1k�sNsl��������I؅����7�m�k]]v�x������#���1+� �Y��uf6�Z.9�p�è�Y�-� ������Ǡ�h!{=�jȥi���pu����U�
#�K��q�N�h��xݹ����J�vgQ�@��M��v�CѰKE���c]C�*��7���8����<�g��q<�W<S���:962v�E���k)�5�P/#����d�0u)Lݵ���b�%�kQ%"�(�31�l%����.	�8nԃk@��0������5�K�s�B�S�V�����f!1(m#-��ܞ��,b�'�m؎��n��9��W��=�nJf\���L�E�%!�JĖVl�V-܍e�L![��.6�7,.95�݀5�SFk51��)�K���y�m|:����_�r�Ff/gm!��hwl��Zw$��::5AKɛ�:�Ӟ�Gk�K�[�����Ȏ�v.�Gmd�3q�C$.�J\;�y�{iy�ބF�Q�ù�fl��L�F������{$�mon��j��0��.�Vv�iw��JD���~vw�/ej����ݣ�)U�pp'/&�b��s�e�R8��"jD���MK�v&��Ծ;p�u�칛�r��[[���kc�KWvt������hѮЪ�Qі�pl�jD8�`�#�3���ju�'oY��R� ��>,gn���m��q�RB`	���5��L6�m�B#
�[-��"g�������%�ҭ:���q"4�w�����^ƍ�9�v9籆�t�\�{<[5�`e��4q&btCp����LPk��z��yc��l��S̳��5	G�g4�BYb���<��y+4�Z,�\95�	h�XwU�]���n�{c!h��DɪaCY��Mt!4���:얺z�\L�"����v+�;t�NX�5�Ak\#N�@8�4M��n��9K�����iv�t��+�B�æ��	�n&W��L�K�c����UF;Jlq�9��/8n�ŧ�0Z�.�֕�.�Œ��gC	ӗ\Iɂ�M�����q'\�^:9�oY�z�S]qM��m]�H��2�cRm���RX��]Vamh�]��vۢn��մ^6�<]�qd 69*ޑ�Q�[�ˮ
���\�Fawn�8r\�#��\F]a4h@`Vպn������gFvb�<q
�cĨN'��L�;]Gf��p<3��yナ�6ا��c�77�׆�]��;S��"�ԻQ�VQV����A��9��pe�MsŐK%չ�sձ<ݻ�o,�n��E�2�b�<ǚxvtu�,.��˅!��B����Ź���px���i��.ͪME�.Ӯ��k���uee����8P�Y'�v&z��#x�ֵLw
����y�������,-ᎎW�IK�4R4��M�س�=�N��pع2n�h�kاgm��K�=����A&���<�J���0�Bӝt �^T3�����n��ۛ!lv�p]�t�Wn�j�ťP
�-.���Ԗ�0t�t�LV�fe10g��ּqx��\�k �j���"(h�y�+�g�W=Fs��q��c.��Y�V�V�zEH.9��x��8�z�&<o:��NM��U�%M��l��n̽�ؕ�W$���j�1��`e�p����v�5qtQ�/W���`����n�iF�vOc<X�w�OO�D��˛���SǱK����;��R@�v�mucu6;[]u�<�1�:[���݋C�܃�@m�n:�:��p��#��[�FP]����H��:��-�����eQ�4v�C�o���#�f1� �鉌�E�ű,��(YuMIKk-$K��>ʢ<�;�u��Pu0& ��Ӷ�r'��,p��h��ݺj��{c	&Pn�v��!	�t*�f��R��vI��(MǷ<�F�F`�������A��a��n�4��毗����R�1�	��i%qѳn�@��̔���]�`�{�6�,u���m@ŇXDx}�upL��bջkW<�q����r�o��y ��e˳�:z{�KJ1�qO3��3e�!e+�<*�%Yь�ˍdC����3�˨KE��@)�iHp��ء����4#=��m�ѣ��ъ�1.:���{-ɻp�$�����	Zvh���cv��p�4����l<v��,=<R�Aƹ��u�\�T�u���A�e�CQ�VŦ@H�	Kv��m��W6ؔd�9ϴk��4�d6J��-ɺg�ݞ�Z@�jp�h�5r�f�t�����h� 8��L�J)�m�۴�1F�45�X��ye�ͬ
�U�e��Z�`ٛo�|���xф���?�]�O	p���
6mJu��� ���-#Ĥ�^�]=����6�^��8%�������z�퓰�wC�|ˎ)��Ġ�v{����ncG�1ض�.9^x�R>̴v!�s�Hj�T�nr�e���uB�9CDM`\;
v�"��
�+s�Z��ɐ�#Y�ڮg�tǝ�'E��{�b���)Oj��x��s�ƺp���c��/�C���p�-hu�2�1���[�p:�㖸��4���pźS_7m-�a��=�2֒��KP��x�81,�N���u��<���[%im �\s/`]�	l�٠KX�l���g=Z����h�Pv '�Ma��I]�6��lxY,fݰ���A�qg�4u�˥2W�'�a����۱��X�C��F=�X{uE��K�2OQ�Ζ�Ŋ��L	MIY�Xh�k��',�1�&m�U���p��`kg�*��r�;��o�N�r7M�9��"P^栮��1	v��a�m��.�.���V陁�7nN�%�6^6�V��竌��y�$r���cy۳��z&!��:�s�8�gLru��q��xzu\�V�9�{OZ��nк���dz�r�!�ښ[�d�")ms��i{Ǌ��b�j�b����*1���h1-���"��5d�65F��RE�h�
5!E��m�*65QE��جmQh��*��h�h�K�6Ƅ���bh��[��m$!�Ѷ"��mɴi6����X�d��j-�V5QkF����Q��b�ډ6*(ѭAhړk1I��m�AXBŤ"�`ȉ"  y��U*�,F���s�x���˔�\)���`��Z@��r�Ўhb��,���_;Ȑ��f�W�����Q��m�$�����k�y/��ɘ�G��o�c�ݹ��ݷtkdz�X��ݮ*t�vzN�l	��][,&&��Y\ �,�]�	�U0X����� �����u���[�k\��ױ�k/I`��W�ۧv' CM�@Z<�Ч[,Uږ�)���w8a��̶��u3�����C��T6��M�pL�X���H���z��A�E�nXH�xy���L��k]�q��Wm�H�lkn��y�ļa�T8��e�����E:�d�ͼ2q
�D%3�M�GG����[��ݳ�kB\e]f-d��'��LF%�u�fx�,tXgiAB��q�.5��ct��14s�d�3L	\�-������S0��˳�⦁����=Xx=�m��V��ًF�xi�=��6�� �"����RT����MR�1l��Z�]\�僦���15v�uw	\*U�l&|fqӪ��t�[n1H�
�ె,�Ҕա��W]X������F���щf��[b�Q��j���^ǆ1N�O �a��r3A�lk.45dq��ɘ�G0E8W�[witŶ�MԇN�դB���ls���4�:Yq)�`{Ys�=q��8���z�9	�E�F�[%�AݻT:"	���ݍ}]�t|�F�PaŶ�r�������!�G)���&o������n�8o���T�۷1Ij*�p��>�S[��b����4%��e�::�G�1���������>\�j$�p��U�[c��.��ݮf6���t�<.�pC��vڎ��Wب��mX��������{q'P�v���]tJ�30�h϶��zP����=��)n8�V5�N�Lc�5�f��4��6�[�;�cm۰��f<��\��l�kI$��
[+T�H��mj�jrr�jж,�`��[P����`2���
T�F�,�ŀ�6�eR�J�A��S��IԲڱ�����I�xe�e%�Uyka%N�l���(�k*�AC�r���P�'q���VZ�Q�-,�Z�`T���h�@%K������[���6�l��=�v��)�,�]��1�rn�[���fZڵ����.'%����e�-��w�8*�36ƚ��R���i�D1W���_�Ae�c{�𳥌�/�%�*>�Y}ޯ_J��յC����!�!�=�Q��Tr�*�Ah7���v��y�Q�ef�w����:��λv��|QH���Y@��@�L
.
�d� �p�F�|��Dy<}K���v4ׅ�/��mg`�u�fy���!_o���?YD�E�(u����e�}���e���{V9�]P������� �\~n���o�o3�󞲅7_eBm5b]	������v�Dq�i0�Z:�eCh�`���_ķ��e���2�w�|��nmg�Q{}3�f�;����֐���0��#�� �YeH�t��n�sx�"#y�axU���&�Kdvp�ן`���%\�ksB�ߕ��o*��p�{{t(PZ7XM-���Gݵ�C���o�Ӈ�ճ�]�5�(=H��!�\���X��oi�P�h"�/��Ў�k]	u�5�[8��)��q�\��ȷ_7C>!�@�ݭ�ݞ�}=\���A|F� ~���MQ��b���ʧr��5��*�v��}�7;�?�n� ��A�[��n�_�o7�N�MU�P_Sx�;�kz��U� �W��� Ct��Л�=hVò���U�VK�D�c�ae(�Q�sЋ�9�z$���s�=�U��Up ���h"�#�t6{<�M�띉��ꆺ����t=�f/�3�|AmCt� ���k��:��B�?�UE�m���:��w.�4������ [�{�l���5��3�@k��eC,�t�-�]p���>�Iz�gK�>ͻW�(�}OY&�����y�Uu}����MS�[��o:���v��GM��Êռ���j��C6�t�G3�3��z:h�|g��"�B�-��n����4��?M�� ٲ������:�t�p4�/��~^��5�:�i�pzP_j���6�e���Ԥ���.���/w+�E�~��y��k�>?)_���e�am�x�����ڨb@ڤ��v��#w>j5�>�m��e���7mx����M8ٺ*�q��PC�4�-��ОJ�a�3�;���t4ׅsT�v]��Y���{�=�W�Z�K�	e�~C�v�ՙ|�h>p8}z��f흟:�n���@��C<B-�AYy�-T���c�h G!u��6�!����Gv��2VA�MO���睻^ �>(�[���QiF��*��A�ۄ?]��j���y=3A]7p<c~	����9�f�6�GƔ#T5Rj&�+SU�+L��o~��B�)����ԥ1-����c���њ����l��G5|d�nua�<G*���-���f�]��q�ƪ��lA��}[A�c�;y��s�=��]q���B��!���������B)�����$�g�dٺn�\�����긙�.W��۽ߟ���e�u�mG�p%��ҹ�v�]:���~���{^3�� Ȃ��H��e�m �-�DgWx^���޳UDw�:@|�C����ǝ��a=�t0�>�D: �!�	�Jf�~�؂7ԁ�K(��h/�t� �Yg�y~�'�F����z������� Ag�_�@m��;��ǵy��?=A��|��G'��<�<}�_x|P"�5�>t<� ��ȳ���� At��ׯ���<�Bp\��;v�Ǒ��V4�{�5�@��"D�+���]$3�U����Y\��@�^����}YLK��)�M$[Y��k����i�WN�Z7�[���q3^��1������|��/��ݟs��Z��kKvA˞0lL2�in�4`ҍ+Y�g�j/`{[��n�h�E�V4*Hjk)���.��9���ݺ���uɢ5aKq�.J3Y�RG7.�-�K��L�[�Ɲ�򂻛{!�5Ґ�흥�,qt����C3,Ƣ1�+k{�;`)�oh�<.�)�!��cE�s�p�[G<�8nr-qs�G[n���z�g�{�=vZ��ˬŋ�&"MB���b�ui�B��d#�L�/�����A��[��e�$��2{��9��a��#������>*��� [�� ���Z	n���y���V���!��ޡ*�x���n�O3��n׈ |W��A�VMCc���AӇ��΂ �2n��3����^�zU����V�}�qqM�
1�\"� C-
����H���I=�>'۳�t���/a�͔7Cܜ�Ѫr���_�]h_7��B����
 �2��e���D7@2�ݬ1�_dh/�R���]��d����x�>(dA� �5��Q�����b�$BT*�¨V�g֭�n�j��6���q�v�ps6�/GjZ����}6���n��@v���������&�"6=YH��:��N���tn�E�P#������곕�<<�������Rm�T�c.{Y�|����{(����ot�v�41�A�X��$z�v���m;Y���թ*���G���+���fcӪs.�A�!u~-�_θ�u�\�;�"��������A�U���9�_U�WG�읜���fdۛs�4�v�~g�� �-�,��8@���6�_v�~�d#/�!�{}�&FS��sWv��^������Ԛ	�z4���:����u��|����-��2�\��A��]'���ǹ��C��P	���m�������M)�j��G�R�J��E�qMg�7.tΦ���%���'=AҎ���M~�T����A� ~!�<Vnxg�3�)��i����n�^����z���#%/�?� � ~-�DV�`�t�>fu A�7[4��.�>O*Do�^�>��n�r{���e|%}+PGv�G]Aւ�_Kt��1a>�O�ګd��V9����C���m��6pz�ӗϬ�:ˬiЊ7������&=Fk��vb�1���\7����w]�{�����Aq|�n��u�#����K]�7�Jψ7�)�m�w��/=r�:�O�ւ	���^ss�]]tE3�� ��7A|t��� �C�nW��fCv�������I]2�t�U�>�/�/��|~!�M�6��@��v.���4�k����U6�������#������Xc��q̢�>��w�����s:��o8w��y�Kt�|g�);7���yP������n�n��-��@�~6qrCn����z���{d���o*7�װ�7p�-�/ѕ2�� D�w�/�n�E�_ChP��������ϯi�%web�2����D� ���k���M��T.M�����ޤ��
��q�^���C� A���{lnVw�Uq"����y�.^�B�!�U]b�eU��i�/qHUp��x-]wGx�^�'�n�������mLr�U�/^��`��D|{�|_W��Ct�%�_͠��tj�f�χ��X��y�׍^+yQ���}�n� ��`Xu�/�>n��V���1�q��<�z�4sF�H3�vP��\V%wD%"L��i�L�k��� ݠ��kV�!�vU(�U{����u�o|�V AƂ�:���[A����O��.lY/`@ΤA1�\<'���^����,��	2/�n��o�ۛ='z����Ar�?o�[A�k��Z	�tO��n����=ӓ���� �_�"�"�/� �AH���[�0��܏�=��W>o��-����A�����D�u藰����HAn��Ch [�[=��G��@��A1��r��1���ǥ�H�@�H��hWt]��O�]��gZ��uY�be,�v�j��[(*��m���ʭ�v�m$��W��uP����mg:w���~u�`�^[U����bL��Q�v��[���� � ����:8��Ob��;�&��.��x}z�m���#�n�H"6�w�&��q��u;��`r9�3x��6fIbA�0[���to�u@4a@ce#h�m	�l�@���l՛)bh�B+�YD��s�����@*0���AV�-u���q���n����sq��{dQ7\\����p�[]��Q����_��'���1Li���]4.Yvv�	�͹�m��3��^����W�������X����{��A��գ�������F��S�oܬ��@+��.R�Ch-��&&:]��_��R��Sy���lY�0�M�Do�簁6�]�z�{��Z�M�G]�"�(�����\v���I�����OQ��s-�ȼ��P� ��[A�/������n�l�0^T#�A=�@�Chyj���y���9>O�W� �PDzWI��X��A=(��|��� �f�ۜ��]��{X��a�����A{�����ЈPW�r�����3d�H���f .�Q��^�XL�s��ĕ��;q�і��U7U�����#�[��n����oI�|����ȼ�%�:T�w��^I@/j��"h Ct���Ds8!j��U�1s��M.�ز3M]�ï���N�J���J7��۲�TaӨ��
#7�u_ev���ET^Q�N��KN�UQ�c+�������x�F���o��v�t��d��� �quڷ4�y�����#b@�d��6�G]/�Z	�R�W̿O)��}��wc*�ޤ3��h"� C�Nm���2u�?t_y�|A �Axx{������^
"g~_<�<��!�f5}��� o�@��Kt�-��䚼�4�"e��MU���Z�;9O.4��A�S{��;��NΗ^aTYm]׬�����{�q,�7R�k���ѱk�&*�z��Vn��k�e �����!��o����<��ycxP'��]�;LC�#�*����Ae�e��^m���=�:YX�V�[-ؿV`�%j���u*��rŪ�R ��_�U�u�j�ea�~�Õ�:�
���*�̷%��
�S��I
��R"��6�Qk�Um�#u�:��)o^�)P�Av�0�l@���`��m3۷�2u>p��$��	�Gw��[+)�cdY4�6����TL�3\�U��7�OX�#�jf�檤�6���no��nfr��*�_k,�$M��kMɏ�v���CuClon�	`�3n�ٷ�^_e�oJ-$���z�hN�k_[�tmb�R�|���ɖ�F%U�w��.d�Sy�wؖ-e�/��՗X��ҳj�����˭�bꓒ�����ʽ]Խ�������0�2+�$��������.�#��ۣX��h��Ó�K��L�j����wY$��īY��)YI���m���T��i��c��:�or���l��:�)�Y�j7r^��q����n��WdUx���j��wR�ʳ�u�����`��G[r]��Vme��u�\ڣ����� �5��V�E[:��u�L5N����pҰ��d��+uu��˥�������)}*�U�f���ƴ����}����LӪ��<�`�b�s{O2��L�����P�}�7�o�I��-JR��W��9vɝ�V���q�e�#ũ[�ﳧ%L�X�Τ��uUc&�7uK���-���{u�<��YݎvR'H�j",�H�C�\y9W{b���|�m�1u�BR�ʷk$��B��y�U}T�f�s������C�C��ʧ�:B��u�{��:}|^�[���a{���q��p�&�:򋐠��h�p��r���>�H~�%#��[�4Z-��U+E�Ս���Ƥ�ѭ�hڍ�X�lEڊ4F�QE����j��0Q��0jō��Pk&���,jM����Z66����-E$j5Rh�b�XFX���6�h��ƌV�0Q��b6"�UcZ5�ƋQ��3DZJƍ�H��`��&�E��,*���~k��0��kyǜ�g��@�Qi�$��}p) ��.H,43(��B�%2��������2�Pt�Rg>ߟ7���o~��΁�Qi(�$+w�
i�}ʅ�C%$d	#�O�k���W�h�A���=�� ���
H)>)�~�[&�I2�c��=��s��� ����p) ��C�T4�]
@̢�Q�*2S�wCI) ��2ᤂ�L)2�H�ϻ�x���{\����%r_ HCzs����O=���I!ATr�H:�B�Y|�
H)�
a�P�j2RA@̢�׽�t�Xk;n���_�v/8��������Z��OB�dm��e���Iwj�'�M�ֵ}�Ru��I'��0��ɨ�H(o�i �4�Ar��h.�)���P�A{{�o�kZ�ǿq��Y�`u�E��$W��T�쿊��{�d����RRAaS̸i ���I�B�%�+. h�I�e�$���E�B�
��]hr��"�p) �D
aܨ[4�I
�w�i �����}y��}O<��z�$ڻ��RR���R
��4�R
Ar��{�ϋϹ���AH5P�ꆒ������H�YL����RII��$Re�@�$��e��k+���2���5��o�y�No�y�|RAa~P}$�@w(���R��j$�@��f�) �HfQ���@�vaI%��<><���o04��*�R
���H,$컁�T@H��̏���'�{�n�T�f�7[��->��YL���p��~�4^j�HG�fxQ�3�zh�/��iHN���d�ɖ�݋�+���TŅ�:�dTT���x�,�uM�;;�RGD�Ŧ���UV�#�L>aH}E���Y(e;��Z����
B�Te�uD) �f\$�@��c$4n���|7c�����;"<���� �#���0�g.����� �� _ϝ���+w��Yz/F�)l4#�s6��x3����U9��I�3�e�:�kz��Z�E�������В�
7ۆ�
@̢�i
H'���G�" �7xk{�>�.�{���A�t�R�o��^�<x�������}�H)�r�l�2RAB�3(�Aa��$2�Q��
J�Sʅ�i��P9^}�S�u�u�a�����Awځ�j�)��=����'nw˭ʅ¹��.��4�Qi ��d�>���JH,(�\4�Xi� fQi=�C��ｬ
H,�2�{P- ����
B�P}E�Q
H-e��AM Sʅ�Q��
̣I�x�j��E�sݾqn���3`����WP- ��B�>I��4�R
As*��
A���P�At0)2�M�Y��x��y"�ځhu%$�.H,40���B�Y)��T@��^��9߫�{���|�>) ��(>t�R
r�H:(�$�8n���o�׎v��:�S)�wP�i��
!̣I��
H.e�$��2�l�e$
̳I�����Ttx��<�������'��||=^�]�*������s(��@���d�>���JH,3�H)2�I�B�
As*�y��[�WxUl��מ�ѧ�6����.*�%-;کW�]�[��:K+�����z��;�0�8�Oej�Zv��o��ŵ�A�^���pC\Q!H�����ͱФ5::��[�g� ;s�ak7i��!��`ɠ�@;6�6�7nkY�i\� @�%A�j�!�X�\�֑���i�mx�g����Hp�g��	y3'im�����c$��[K�YD�+#��ՖDW�uے{Nr��5�P��Vu�ڒ�ָ�.���>9�^��5�Ӆ���ŮG�zPƆM����}�{�o��ϋ3h^:��j+n�:�s4���Pp����4i�k�q �ި?@� �*�>����$|����@��f�%$*!�F�s{���=�;�>���7���A}���RAI�3~y�m��T-���H(�- �4�A{۸*�)��eCI����- �hd�2�����XwwϚ��t�܆$R���i
H)���P5��w�;ߟ���o{�y�I��A�� �*���R
Au�֠)4 Sʅ�u�����y�x�P;�- ���^e�haI%!L9څ�j���A�f�CI̻��� ��/#�$|	���5�H/T���_�+��W\�Vs��@�Qi ��Jy��$��rᤂ�Q� fQi4RAd���]�P5���2�C���u���s��`W(���!I��5�
AMD
a�T-����P3(��û߽���_;�O��^n��݇�
H))
aߪ�R
f�]��j����|=H) �v��Q �C�i ���E��
H)̻���%$�$aH�ZF�3�o���� ��Mj_ H�[�z���N��{D�&j��� �*���uD) ��H)�
a�P�i��
�d	#�O±�Tn�hG"+��Q�bDK,{N�ݐ ]����%`Ե ŧ��ݧ�q��R���
H))
a�jɡ��P(�l�A`i���]��Q 1��Ii�/u�K�Ck)�����- �h���;����}�{�����XVrᤂ�PaH��HRAd���]�P5��:H)2�H:��W~N��5=�u~yw��Rg�FHϐ}m��\�71V�0����9X��7�'�w�����z�$�j��uc���a4��+n��h�Hw=��S��fT-�) �s�ZAa����˽�z���|o�y��$ۻ�RAIB��ɦRA@�v�$�H.e�{���w��u�
Aa��- ��
@�Zh) ��%;��JH,+2ᤂ�C
@̢�j!I�� �%���j1�wLQ1�v�a�wu��Ғ5A󤂐��;�ZA���ќ֠)4 Sʅ�C%$)�4�XhaI̻���;�r���a��- ��E�����p5TAH4T3*O�3[֫�!��-�����H�G|�YC%9�� ���k��7��������H,:;��HRAd�S�]�P5���
B��̢���$2��SH�2�l}�]�}��R
�(�@���{��[��#���|<G��I�RAH,>��l�I���@�As.�h� �*�$��j[��LL�4�Y	Y�ݚ=sv�E�Up�3�	��jm,�%	x �-�s~�����E�b$P�O���R
Aa���I �fQi �2��0w|3{�c��;�#�O�� w�I!�w�i8/]��E��B�^f�H)�@��B٠d���fQ���PaI̻F�RP�0̨[&�RA@K�W��w�߽��N$��As۸*�)��͏���&EwZ�Tpo��ϻ�5�E��$S%9��	) ���- ��
@̢�]���s_{���t�<H,�2�ww@�RAa���R���
AH.�5�
AM Sʅ�@�I
C2�$����]���o70F���g|�����`��V�5��	Ns����˨prWi���6��/�sq��*�y�Cث�oUM�9	��]������K���� ��{\�g�~su�~y�o�$ۻ����
a��d��H(�H,4�\˸�D�EC2������E��) ��f����;~�����A%${ۆ�
@̢�i
H,�Ne�G����;��|�7���>) �֨>t�RTr�H) �{o����W��^u�@R
z�L3�f�) �s(���Q�$2��Rj!L3*ɡ��P*fY����i ��p>��θ�F�+�s~ߜ ��B��Ϸ������_�<�y�Ϡu2�H)�FJs�p4D��XVvᤂ�C
@̢�hB�%2�˸
�3}�#OP��EBQ�f$ J�2Ssm���f�N7+t���a��K�6��3�FΖ����t�R
{E�Q
H-�Z��ЁL3*�FJH(P�eG������+�/r/�߽t���>�H0����>{]u��=����0����RA@���$�I�]�Ԫ ��fT4�]F fQi�@���d�2���JH,*��s�O+^n$R���hB�%|~���� ����Z=����D�&��I �w(���D) �gu�
AM�2�l�w�{���O�k��Ă��h���L) ����
H)(B�sꅤ����f�M$2��Q �P̨i �}��KN+�������x��� ̢�
Ag̔�n�) �垹�~2P@���Umb�u�u*��� 毐-� ��]��Y����ݩ�cՃ*�A/a|E���su;r���k**�Qu��E��-��M��c&ߍ]�&x�U��;�NdҜtl�c6��#�K.˾�*]�^ӵs�k�]5=�O����1��3Ծ?<�-�ȷ@ ��V���ص%�r`{��֦)����� >���_7B���gU��h���'P��5w]��n�h�k)�aڣWJ6]��GfX�Q���� �B ��������5u�l��x�wQ�z7T���l�z��Z��'��q���.�E��챎�E�fm�Y*Elb��J@�()������ˎ�Ǹ�eW�?� C���<��}�՘�V^�z ��R?k��?6�n��-�6)�ZEԣ^�ד�����|��_y�@��|�t��@��k�V��}9�z�W@vׁ����'y�{UÉ�x�wQ����F����{p�/�� s���[�� ��E�D�^<6VR�[�a���܂�Ӷ�{пz����Ń*���ޤC���~n��6,����K�na�^���!WT��F�wc����U�5m/pV���Z��K�ݝ�}B=��v�5pѡ�6+P3m�B�>]Y��Ӥ���!��񮍳k�W�3�[��znU�TL���Ы���@�ʼ�f;Xg
�V1/ �W`�ܯ%����뺻��H�5sڸ��{H	ֺ�o��ne�śi�:�3b�,%� �rOۃ�;q�1�+��*Pm�X3�cf�[�֋�!u�h�l7$�]4@��\�n���ǱvKQ��i�B�X�Xk]��ц8���Щc�����/��kK������v�G�TSWnv��4��
Ԡ�5��;��������n��,�6�K���sǷk!/(3���{Tt�wʰFovZm�\-�O\��%a�5��G�/��"�{qV*1�8T�N�4��@����]�+:�V.��wp?�QDo/�'҂L�[�!�5�Y].���/3:{d�������}�@@|�2�|[A [�8;��ȴt�?H�>� A�W��ԧw���=����@2����T���z ��(�@�� e���� IA{�+t�wr��p�n� ��2 �t�̳۽z��e��eo�n�"J_@)HFJ�J��Wvz-ښ����F��.��m�4��SM
m�zN}�����[A}7t⏇��.����Y�W���y�ި�A G���"�#�,��P�u��-�+9=��U�����X�������f���s~�ב��H<��*�/�bו��gC\^#چ�s��-�59myY-����!$�v|�ʴ],��Ӱ���/4���Y��;p �\B-רym�^�\3�@�y
�_&���|���L�`��|�jiڜ;����]�^ ��g�D�"�"-�D6��^s},���A|�G]/� 6�M�w7ç����`��|A=�@�8c�<Mu磨<�R?� [�~n� ��n�O}���c~.�!yn����nI��^|�"����HChϭ��{���ϑ��+j�á���d퇎��y���l��e���D��%��O����H�;�@� ~?6����o��s˗�C��H��9ll��Lcg� ;��]"��[���j�;�ƻ5'�}f� AY7L��==`�ܗ���i�� A������C��?/�P_�~�� !�n� ��E�ٻ؃U��hj�S�[+v���)^ѕ+�2�>Rî�kc<Xڔ(]F�;u��f�f{����>�w��/m��/!�h1�[�[?��|>��t��<f�ȥ��W�t�-��!�DKTl/v�n��0A�"6�v��=���MwO�p]�^��G��ͼ������@�[�m �w���.gӒ
�t���od���R&#�/a@��"�?���_���Uu"	&��Ҫ4R�F���%[�j�{K���J�\݆J�fՔ�.o���e�|�}E�@��n�μ������m�d%�7fYU����o(i���"͠�� �� Cwfy*�S���U�?��C�v��-��wV��Oލ�A|?	�әk������u��|P"D��A|At�@�_ ��]yʥl�Q��~��}�
��.�Y�<{ԁ�!��|�|�g����^:��{y+��:=�"�#�,�3׋�;����˼�!-���L�^3M�Ԝ�u�SU�^��8�ږQ��Y�J�h�n����{�s�zV���
v��S�E����Vk�{~o��}o��o7�5y�$�	�-݄!�l�n�@�A���g>���[~���+c~�b篛�2���� �@�H�n�����͵y�篾{u�6���cS���\���/`l�nq)����g��&1/�Q�K��6[�������#�|�zɵ� ����Z�7��E��_�h/���W�����,��V�y[#�����vޤA0�X��n7�o_�M�a	j� ��B��ZrH��<	az��9�yP?z�M�x+�BG�𺹗~�+s�/{_N�ve}�ϊ �E�DYg��*�7YU��a���li����Cj�R�m���U�`I�����nM-�>g�Ff���,��r��E۶�;ݖukv�����wit��U��S���1�(�n���7�({Os
���z��k4�IwZs�Hq�����w*�U��&٨unUF��\�+��\�.��o�ښ������y,�A�����{�3�{&Se�y���{��Z�5�ǖ&f��e˝��# ܗ���le�
��Yx)+��<�U$Csv���j]�ȔәbsvMǳMI͐� �r�*={�;���	Lg4��)<f&�e��y{mҤ2ř�wv$��lt��CU�%�)�b�e��7;c�DN�
0�k���%$�wL��]�3��*�J
�h#ݏ�]��@t�B�Rc��V4�m��+lgv�Q����q,��v����k�*;�U��]j�mX��Y,)\(7�׸�����q9���[�]y�ה�M�ofܫoe\;�.	ٴ�Y{V����0�ڔĮ�+Pc����gm!z&��kmwWVL�L8��?�Y2	��]lŶnk��)�1껾�����]�M�{V�eޤ��;O9'Y.���t��y-�(5]���77)\�Ԧ=�v3�kT�}׵��ڏ4�U�(���8�\��z��̺B<���J�|9Xs])*Tx͇*�wi�i�5b�wWێ���[�zV�
N��vݻі{~��A�|x;�α:�YK���2���X9����v5�������R���ļ~Q�|�D�os�!���.�x.���N�1f�M�]��/�7
�9x�h�EZ�Z�3�R��UW�XnME����>���&Y� Ů���{�a�׆5�j�|i�\���wmҕ�Z��Lm��s�d���:��\u�z.��|�yt�(�
E`�#hf�#fj-��¢�FŤ�h�3*�h�	Q�F�$ڂ��A�AX,Q[�űQj-b�-���(�1�ƨ�b�m�j(4Q�!�(�KE�d�E�Vѵ��ō�����c�����Q�*���ܲ���sa��0�A�Ο��B�;qq�x�uqv�귭c��Y�M��p�f#1k/+7�1�	m
��R��ĺ�΂�t���at9�7k砌�k�-�.�墅��"3u�
�U�SfR��k��X�$����N�N�ҕ�[���j ���:��T!���B!i�ǯ�s�p���W6m���Cѫ��#�G]s��$.�Q#�mN�]0���	Y�º`[)��c3�����h:�����w������q�v��EsXqё�8���[�Ik��|�4e�m,[r!�)r�3 ]C@�b�˖ i4Vj]7Z�T/5��D%ٺ٠�� ��{%�z��ts	ٯX�2�g�-�p�o%g�Ɖ5��^�nN{u�ά(\H�kav�t0B:��nC�%e5�-�#t�4�(]Ԍ+��BXؗ�1����63��%pS'9&����4t����[�q�c3im]�.�,)G.#�H��aq1.C9DS�m{\�xf��^��X�ꔋ	�h�[u�h\[q`����Ԧƶ��bޤ�i=n��N�!{��p듪�X-!J9�J�xGx��痌�\�q0s���^�́B��T��!���gI�v��ەu�C���
8�%�I�[j��j�`�6ݻc����E:�e������:�ZC�O\��[�Z�z<]��wh��Mە@�0mC��n
`�E��i���3J0���oyr����U���>;����q�+ g�����Z��Y��ܲ��`��%��#��aBN6K��ѷ�D���_X,�;a[7�y��oYf-�O3�u�Jv]�ݞ:G�meġn<8��8���+����GD�쫚���6lc&��ͺͰ"a=�`]1۝Ѱ�P�����1�;	ړ���(����h����WN�Y��O]9��6h��<Z��+Tt�C��M�{
`6��8̱�Ę�m�F8Ib�%1�p(K�;�v�V�vs,j�o�I'Na���n�chR����>�Sbu1����,֭������r��[��ɕѮ]�����<	���tp���u�0���������)n�F�q[Kv��u�0���e�ء��ڪ���g���{��(�c�n�rv��t�%j�̭�2gY�J8��I���e󭥼x�{h}�,��FV04m&�n�5�	���8b#AC�u�~���<?�\d����${)OE�)�n��kv��,⨺�iiݴ��"��Bh",��]���Z�4��V��Oލ"j#޷;�`��Th�{ }ԏ̳�t0�A*��Oy�&���G���:�#O�W{��t,ר� �h/��z�n��V}�Z� �R?i�!�-� �����%US��	��#SF�k� ~>��>_ [�A��n��y�Uݞ)��Q��ۨ ̀�hy��Z�XU^v��]�^��g�/�q[�y^UWw�&R���HǺ�7_7C> ����ڨ�Ϥ�4P�Z痦����A�j�L	�� ��R#z�n��мw"�p!||ڞ�Ű�ðKi�
��#zk������M�Kț^�ZkL�n��/;E���c�բ;��*-��U�j1�VymK���ڧ]@e	�(Հ���%��"kz{}�2^����U��c���
�2�Uf�۪Y��x����}7���y��j���27>��}\�嫁#y�}H�=>��P^e�<������5����WfP�x����\������Ot�����}�P6�@�H�CV[��9{ոYyf��=`�j������W�sA�����H�V\~�y.YB|A�/��#��'r"�l�MTZv(�����W��h�b]���>�n �"������a����۝�Wz鴥��CA<��[OtL�<�����	�P@�A|[������{�u/h�[���(���L�Pкh���o;�.���g#a���(XWA+F��_.�1���6�6������b/Hʯ/2�D����o��Fr�:@�~mn�n�`�����7c���}B�5�����h�Eo�?z� �����<�齫�����r�6�!��`n6��K;~�^��w1W�M{:u��岧�í]�:$���A��qUM`w]Y�(���//3�8���9��՞.U߀w�#�m�Cm׳��}���&={��J�?L�}�_�'�� ��q|�a��6�Bj�r�cYΩ�j�Yea���_vl)߽��vH+t�5�wa|E�*�<����wv0�Q�k�6?��A�f���t�U�p��V�S�������"��n� �����{X7���QCBJ�_6�0� l��Qd�U.����f%kH��6Q���/z�|��e"����h,����N4�k��ٕ�%Q�zFLO_�@� �����_�[����&ݺ�1�>�k!|E�|갧��zw�)TDi�� A|����s���ϟ�W�F�HAޠ� 6��@��
�tL�=���A�v�,o]}�� O�A\_#�����3�j5���ǽ\�A|C�G�v��[��Z��٧%�cAt�7+2���R���n���6\�t����ڪU�gq���{Gc��W�޼LϽm�v�.��}h!}��nA+kK�lvu��� ���~�\E����칽�Y��_����m�/e�M���9�ݝH<��7���mE�@G�]��:��6))����ؒ��G�TMثca).��8f4p�c��*�0���JXc�����I�����~�e^�;�N��\Y�Nc�B�B#��N
�wtUA���Մ@2�
��-瞥r��>?hm���<�<�\�:�˯�Dtn��	���Q�e�	r���2-����v�YʛKyb�[��؇9��ʯ|A���_ �n����"� D����z����A�؂e A�VX�Ln�٨��Nc�Z'v �su�w�O��z�2<�\G�a�ב���mCt4iׂ�|��A?{=V���k�3�˺���"h"�"	n���ʊXA[�%V�S��Ə���dն�dw��W������P{VO3��=u�Nva���O�Nŗxt-�:�q?7��:^W�=7���O���| �����6Γ3E�6�JYl�P3����N.�r�^���x\=���Q��hᝮ�X��ع[kkGn�����.�0W��4eK���[��Su�9{�o�9ه�A�G����x�-��^k4Љ��hC\h�)T�3�WK(�۫��:;G��εt���Y���s^����\���{Q�v��z�e,�_\�6���.�߽ߐ�7�U�SeP�2�ƺ��=�ͼDtJ�e��:к��5WCς�w��v�t��Y����|��C�õ�2��������~�x�#]#�mn�_���<��~ow����R�������_j�����������Щ��l�6V|Ct!�|��ާ��U����̿����v�S;���{�؂-�����wَ/VLvةA~�_ w�|Am�bw�yw:�ۆ��LF�A݄~��jZ��b�t�5@wP��"-����*�ɕy�<�`����'n���P�}Ё;��|�t�6�ޡ�V��ҵQ44_���	�p�ð���q�2�C���=y�T�Z���0A9Ԉ�@7Y����������n��+��Ϋ��s32���ECH?\A��-��ϋt�{3�V3󒟩Qhk�� �*d�W5u�f��۪)���S�n�����ۍ���gI��!}��3�o�����9�ɿ� }��|u������1����Guݸ�����MW��Ծ ����)�J�r�T�|5?�g/���:�!��Kt/���Y�������C��{P'v ������a����F�,�%` ��9H���ګ|�·ݮ��+�|A/`��X�Ki��������@���@ ����f���(��0vP�5l9OF��Q~�QP&#�;�����7H�h_�e���̷����J�Q��m�t[�Z��Gl^�rq�U�q�y�v�%;?]:�?9@.h [������q��>��*��+(V���g���}t,����"h"�A-�ճź�g,�$M�;Ay�Q[z�V��2ߣ���{A�-�brD+%A�Dԁe���-�Ё"��$��䜒�m�_c-E�/i5�r���{2��&A��h�G/����D��+Wb���Rڎ�
v�U��K݅�������}�e�����n�?Y����D�@�����t�#*�Ul�GjBƂ2R���ӽ8e[>����Y��\���q��7sR �v�û�t�ȷ_7C��Lʥ�[��h/���ov��-���A�(�+E�@�,���������Qi'�[m�x�y��>�gG��ue��!��n��f-9.�U�
��@�nP�B��H[A[�,[���H~�QP$ƈ<'�| \-�|�e�|Gͯ�� �����;y%�(�BnyOX���F��\I�@����[�tX$6u�<j�"&R �)��n������k¬\�Zr�n�"ۧ�[�51���/`
���,�[���%�Y��l�?f/�n �v�nѯgjC�E@�� �z�Gsp��+��a��[��oC\T���t�"�T�3#�K�mQji=0�9H�-~�5.�����u�y����!!���`�7�����Ct-נu苬�QP��p�Ũi�1�:4nD
fH�j� Y��[���1�h�)��Q)WR�WN�:r����S���#�[��-���Rj�/���^�� ��/���n���j>7h)ɍ�כ��Ɇ�z>�U*_�]�#6��Ẃޯ�e�m �-�@�TV�p����!�۞tk�OW���pems���qC.}��b�wRO���R �a��m[�?Y˩���}��U$qQf���`�U��Ȭ��҂ ʄ"�/�-�dbY/���w'���ab�)|~ 6����|�}s��ݕ�+��F+Q��^�%Ϟ�	m ~�6�E���Y�kp{�=��j�ۜwV�9_xz� ������z��u��)0G����kN���S�Y�;WW�牠\K�M{S+�(���b!�P|� �\D�K�Ɉu���m?Γ����,�����s�tR�f{u)؁/�Ͷ.ݒ%ڷ/�w4Oe�W��nʗ�O�=a�J�u�կIWHj�,)�E�ِ��ػ;Fg����n��0]�D�kHz"6�]61�!^�V�Mͬ��r�7L�a;F��l�����/\'��n�Sm��q�U��3�Jl3*���R�H�����C0��@�a�PlU�����mw��ݸ�R깧;����^��녹&ț�wm�k�lً��(s���v�-Z7qMa����^���Dn� �[��tPo���a���#�Pz������;[�������v���_� A�@������x֏|F�/��n ��^���7���ɧ=h�A�/��N�w�yr����- OuA��-� �hk�V)g�t�vz�`n	ۜv�V�9^{Ԉr�7@ A� F���iδqJ���\{����jp?�Óe5$G�/����/��5uT����e|��� �[��h"�4�9o��O`���$�E�>��~s��˫�+��P@��t�&�{�e	�oR2%bH_ �e��6ć6�"��sm.�5Ynۍ�l�Og�YxF��/���_&�_<�\Ͻޭ�����2��;����rmB�F�����Kt�o��Uh��Ŀ+m�m�e�u1X���r��j�v�g7���Ȣ�4���u����Y}TL�-<��4�.�w3re��| �g�p/!A쀷���5ɍF˕$/j�^@@�3ȷN�;�R(��ͯ���� �������^��V��U�ƪPE�����zw>���++��PD�|�g��� Ck�U
����U�����H��#�]�ޝ�s��Pʠ'P
߽0g�s4��;�_V|~��-��t�6�-�5�{Z�ȿB�n]�ߌ�1����V�Õ$/o�^@D��E�@��sהfה�,���pV6y*}H5u���s+nkU��n����jop�f�핚Tl���j���;@��|~#Ze�{�'��N��]R��CG.����
���B��}X%���n�>�W�gi{=��c�b�pb�n��.ǅO�z#A�� � �q��o�$y���5�J�ޠ� 6�n��[���i���g�ҹ]��4~�����[YoNNyg���Xg!k.�Pv��R^n�V���	;B�*8��U��v�d}��X��W�.�nU�8ڎ��Ƙur���R���]��Y�,�U���ĂJ�8�a�Vs��+Hm�����=רiٷKs��ί+!Ǒ>�λ�:&z�V)WE�:[۴n�VS�nSv�c�d4�+�vCD�e��V�k�
W9�߻�n�H�ݏ��P�ǎ���Op�D?m�i�v�;��<T�A����`�wZ�D6M�q�`�g��p��Oj��!�����SK�z�)^��m�<���;R����a�kޙ���S`,�Kh���(��2��D��Y�gF;��1�z�i�D��.nY}Ʀ�\�����p��奸���R�n.{�MΥ\P9d��$�T�7ث���6K�#��m��&�
���ȶV�;}֪8ΕY%����\��sF��c/��q�<<*����ήg2m�ƭeپ.��x���t�mʛ����;�CW��3\�u���o�����G��y+2���i3b�5L���D�%
�Z]�����[4�n�2�r�Ō�iִ]Y�jq)���r��w~{���wD��+/Oʍf���}�E^�aۙ�r� �G�T�q,�"�M�NuK-MB*]J��f�5!̻Qog��LpҦL�H��:�������U�����콛R���C�CA��r�e���K^�w7�[玫�k�����zZQ$�ͱJ�ka�����)�vf��,�}���{�^�lF�(e��Qmʷ6�l�̔b��cX�5d���h�N�\�k,cb*"�F1[�nX�h��4IX�T�ܮ�"�(ڍ�������(�b����r�s���[�[EsRE	UQcTH�3|��[u��wH�ݑ�C��J���  ��7H��#I��V A� F�G��m���wo6�w���^G��݀���p^R��	�A �P_�|�[@7O�NԤ"hW�n�b"�<ݨ�c§�=�{�� ��?�@Rզ�?x^��G��BҢv�:zz�=V��	��V�Sj F��3��4ƍ&�ʮ#���ye��\e��Y��.ju�	̢=00CQ��u���gN�� ���� Amn���_���C�^�ґ��CT�����9N�Ļ�W�?{�4-�$)�쬚�؆�{�҂ ��E�@��Th:b}�a���s`���4�������h [�אǌ�^$X[��EA|D�� �B{dV;oW���]v���%El�_��)!�ۻ�:�#�uf*��S�}UT��j��G�.�*���jKws�(9_
�?m��q��=}g��v����%q��[[����}ʱye������K7��_��&j?�'ձSn��浍�%8�x�}��� [� �B[�'c�������`Fhch����`n^���{U4�h3b��`Ͱ�a���'�w�4�|�t�!���V��w��[o(dF�/�CJ�jR��WQ�D:�ݏ|~�A [�� A��v�}9.���q���l�;1���Au�#/�\��Du��o(+���`�wh/�n� �"���hV�;X�����v�5n�����f4/`/�ˀ��#�tа�K�(Y�|\�Ct�`֟x��y���+�{Ԉ.��I�b��n��7�܂-���A��t:�����C�AI�q�e���n��F_�%� �q|�t� ��9u����#������yf��uSQc�!���K�c��������������U��F]?$��Y�{[}%mo�i�b-l���91=���8	�C*5Də�Zi�o3T�4/ep���X�x��^���<�\�n��X�/L��	L[6�[`�شVjC9��l��U7bs�F�O���{;�y����x�|Smhy�P�V�B RXL츊Ji�ݴ���͖piGbX�-�lqH��m�O���<kd��5��J��.Bie����0�r�@쎗�.,��cGNȗMYv��o~�}��1��Y�諬�l�UZ<	<Қ�a��lԱd�i����{��Duʱ�l�7��c7�,�^y�so���W8�x�� ��i�x�mꠁcA|d� �A��FE��@���~��O� A�_Um�KN�n�͸N��v��ǽH� �/E��8���izW�� ��-� ���lMc�P���S�Ōl���#Ө{\@7X!�u��n�a!�fV�@IX~?6����ޛ}�����\�1��Z��/��:�����n� ��_곽~�A�� ���;~�t��IGs(��� D���=�y��ﯾ������:�D�[��p��<�=Zm�I��m6�V���G����Yw� D�n��C��S�͸=�Eu�#'P����d=�� Am|�� A�]��7����Z�����ׯGN���Jg���#B�u=�6�̵�����XW�Y�+]�{��Տ���wU��n+�( ��.ӝ,\�D{���f�2�������l�?{5���M�1���A$��n���wh�>z�k@ A�@&���}%�и��a_;2��nmmT{�� ���$A$�~2Kd�F�'�g���+/R�eA� �H���gWK*��EK�B�gP@����t��з����% ~�+ �$A|D������/���3lo��wӚӼn&٘߁�����%}�Ji����9���]D���s���v�.�#^��<;6[�%�Oc<�g�N.K�@��X'�AH�D�'��R���ʝ[Y���;T�R��}����`��j����D,�HL���q��E\z9���(/���/�3�F���������s1P���Ug��p`{P@�������Jr�RK�B{��^L:��n�)��{Z�h�v$�CwV��K��*��Sc�W��;�Ŕ6A2z�{|U�^��j^ݽm]����f���/�����(��c��no~�Tp �^�f�s!|A��A$�`��key�ת�=��sZ�Fd+&��ljy���ϐ����;���-z�`�[{H�zK�� �A����7�X�:E7��Tׇu�S��[�CS0G�v~{~�_ s1_�"�����{��t�}B��(�Rf����$Y��c���]�����"�xx��U�j�~��"JG�$�b�h�o]�ksx�����L�y��&���@_gzŗ�@�d�$�,d��夕|��{��JH?<A
ɡ��'^mM��ϐ� �z��A�Ù����3ej�jC�z�G�D�}%h �:<eW����qL�Ru���~�AD�BH��(/��*��3��U{'��5����I,]�����{���Μ(�A�(��~0D�0��Z�yG[6o�})V�}��FS���q�����m"��e��c�7���G�K[����9�aR���u�}��Vo�P� ��$�/�( 2�"�W�y��� 
�[C4�����tg�Q��������$����,e�+g�߳t��"���<q&�뫓Ʋ6�ť���H�e�7�5;��MW�Sp{�X'��s*��8y犥�]I�v���8�]���7&��k�Q�#�.X��^�2�Lʱd���WP�*�M�'�{h����V���~�eݸQ��`"ٮD���,>�qg��C���E����~�ឌ�L[�o�<н4{��43��k�;��w ����H��)�C˺���G�CH=�ř)���3��)��Of��FVz��P@���ƨ��/�f����)~2E��@�)eW�]k����7r��t��f���]ۅo�v�"Ā(4��W���-e���˧�-�K�
ʹn]�X7{:�ԙ�(�=��r��z���XI.r�6��v&��nw3]L�z�g��N:�8}������78Ѹ]u,���R)غ��/���:Q�h�,&[��k�9�Ie"�[R�q�^��3��C:�R����伳�7M6���Dv���{bݞz��@�E�S��xpe; Q[����b�-�M�xx{1X���>�7:s��9�-�R0s��m�@�c��!��n܎���]z��3������`�.�	��ظr\��}~��?)���#.X:���%�#��#��Y�a�=�=��V���!Wll��9���	"������<�Cx^ v��~E�o�ݢ��j�j���R��@�X�% A2PD[/*���,�7m݈sk�d����5=���h�Deb>�\_#$I��{j1����z�@���D�"J@�D��v�þ���Ӄ3��s�s�7ԫ���@)�fJ�(/��]��S���ު���By|�~�d"X�N��H������A�����ϼ�}@�c�ܠ��d���A$B̕�=[N��(mSm,\�������/Eb��������_/��}r!��й~}������Q��_{-l5�쥫��Rs玤��}=I�<� BD$PBz$���	�5$����"`���G���;��U���gO^�8�;@l��:�|�"IX?( Ecc��ҳ����l��\�B'�:\���浵��W��͢����V6�m�7*}s��n�{�ނN�Շ���5��z�5�T��X&/����U�D�3���c�"��*����ީ��jDl�y���H*~����2R����PD4)L�%��b�2�Cm�����k}-0�@5[ �p��_ �X"J�+�Ov<�C	�D�1��)��Ku�4޾�~�����J n� ��{"ε�o�7qb/r����Ўe��,s2�;Y��5�{�п{'K|�w��3���׈&w���IH��ǍJu��o��[{��+5&��0h����9
3���u�`�۔�6c���|�����>��_��8p�4M{l~w���T��V�#M�����Bn�����A�D0��+"�U�^�����e��6w��8�iF�~ӥ�r'��	�~�}0�<�(�݂{�T!|�I�6�&�&�\߼$�A��k�{�ڷk7'eR���4e��w��M3ƴ�.[��7_vZt��*H���^9��Q{<]x�Ncn�Q׳.;k�8�tEz�;�;�ȝAU��JG���]ĺf�p����Z&x%[za<�W��LEl�̀�%8�V�a����@�bH���� D0������f�?z����͹�9���9�j먽z�F�4j9�h�0����;W�iƑ�RU�iB���L�2��-��&�I���3k�=�̬�7	+�����C��#$V"D�kQ�:/l��Х����<��_�Ȼ�\�O�;��+���ř)L0����Ԓ�U��0q�Y�
}��'���`qS�Hh;�����ul��"�|�+@? $�)MF�l�T��Ƌ���բ^yf;s1��t�@�z����0�_�C���w��gP��B���%�u��{]�c
"~��w��E�*<�sn�(��^ݩ�v�8��8"[ښp|���n�����Rf=[��<����9�6�ejَE;�U7��_����k��QK)̻ڟ���9b̔� �% A�X�d��5ƫ|������.텫kf�$�Uʷ������2EdC����gy4��U�)�"gz�cI��ή�n�{͎p�������D��՝����F�����%��X��VƈwY8��c~ �o��[9'
�`�R �a_$�,%C�f>��xF1�޵d"�:�N�~�}���Y3�����n��yݱ3i��_$B̕�0�M���Qew�#%�[γԶ�-C�z���x�d�� ��"^d�߽~��*�xC� ���i�y����wk�ϝ׈ ���D�^��$wn�43iK<~�m�d��2��w���V�ߐ_J���N��K���F��T�[@C2�.K�t�H�K�[UuI�����.�IW������RN��{�lT"�P�n�j�[����e5���Y�;CB�kq𽠜�Z�1���p�~�c�v1�w�8�i�f�8����>�־�k��,t.q]��#E���v�6�Gq������Y���˫�̷9�$S�:��.�ꦆ�Z_X��g6���-�wv���m��g�)�*k�U%�n�l��c�&��1�ic��U.���6�X�;)�*�Et
R�XRB�ql�8�v��7S3+���Q��(��:URi�e��e�;��oϯ;(��^�-
�`}�[µ�u�+�K���EU}$��ze����6����Ҿ�0��-Y[v+V�N�&�qO�&^���bO�o�j�֌�Βi����S}}Qt֙�O55���ݭ��.�u�Y0�����ڸr�j����ve�m�b�e����R�]į���R�����ۥ�5JFʽ�4�өoL�rݴ�ũq�h��r�j�s��X��kf��eI�(��u}��̕geNuj�M���Ir���fM�p�vw_��L��&7��w�6b��H:�&��*�=��w>����}N�ڧ��yƫG2��=�Sh-߮�}�P켣����o����dN�"i��`�׏�%��>i+�2�;i��3��i�޾l�Ź|q�șͮlY��{R��yu֎����������!#�//��;��Ft�顚���T�0:��6��p��gEF4�k��͛v��qwL�W�Św-�����J�:0�h�c��<n����_���[���@SQ��V�+F�Q�MQ�[��-�s�͋%�F�V+ElZ�V��X��-r�Y5��ɨ�E���k&��嫖�F1F5EnW5r���F�%W-�nb��ʤ�5͊��U��s����+��TE�UsE����st�w5½~�,W5�tv����HcS��G0��y;�j9�����*c �n�u8�P����;u��٣�ɐ��-�'9�n���K��<����Q�-ל˽6��0�A���0cj�P&�A`:�e��$<�\�؞�;���:�n;�d]�9+���<�sŘ�R�*Z SZ8���;T��gq��pi�6:Gt���8�8�F݁8��B:1��'Gf�$�Ν(��zcNoLv��o-�Q��5�n���]��pu�ܑ��SU�V�\ll�1�Iݸ�F�HKd�Z�V<���ѓh��`��vzJI�L��b�5c@��m0G\K	2��*o�@r��t̓w\�չ�[^]�t/<P��u���uո�6���iN�bá�B����{&���ͥe許̠f�Z�: ѷ�J��CYV�����*Żd���q�t;�ɣ����K��f�%[#�)�;s�j�/<۫����wE��<Y�Z���v#�d�Li`�
E�z�=�; ��N5����]�qK�8�=�90�9�0n�{<��q��=���7a���p%�̶���*��k�%�F��p3v�K`3,�^�c��u��A]a4�6yl.Ddt���JJ��K��a�	u.%���2G�X�F۰�Y���k1^9:��!�\��Mftv�v�C�0�L�Mx�!���ݭL�rZi�w<m^�zձH�Ð]�n݇�c�'v�#��l��:�m.Ĝ��1���۪��f�^�����MJh4��Mn1iZK�fd�E)qq��\vh�y��1D��Kv#����K-�z��� -���ϥ�ׁ�gq���t���`�q5�=�s��׭ʊٝE�X�g�Lnʤs�h�	�#��[��� nBݽ�+�ʇ
��`��+x֘ؗL��UIb��-b%�k'>@���n֜�"�����Ş�@��Bn-�Qr%�{��	��h���X�&t56��j#�=s.8r�����@Ǵ=���t۝Qjgcr��8�:��vN���Gj�$�V�Pݻu�p<��썖ypX:��n\wS�!�l�9�B����Cg�A۰WO)�B�LC[�]
T#-���4���������$4��A�Ɂ�H�2d@���u���6�j��K���)^����jNS�؏1S$�E��Fb2��UbR�N`�u�5��[MAXHw��C�g\�}w�آv��x�	M�'���������)�e-���':���.N�*��Y�@�}b̕�0��VOO{�c}g�:����S�|w0���]e���VP__P&H���a�/>yCv[�Y�
�����Q�L���t�Ѡ��?!�����5������A�AeC�h"J+w�HW+�uX|��~^�ӷ0�/�	��drU�Kd�CȽ9�п�(���X�����
��w���s���[��� G<��tJۼ�#~9��{�DC����D3<�m%=�?���Y�o�F����gvM��	��@��X2R �%U�k%ǔ��-=��.���	�4cƱ[�������C�����\�n���V��Wly�=���_I�H���w�>�Zjۘ~��֫;�WJ/|�`n��?O �2K�J�I_K<��gf�Γ}v�F����f����c	�ꬱ@�u�޾����]Y�i�K*��!I�UPK���,���d̷\���̻����B��% ��o\hx��Fd!�מ��U�c%���D��;������Y�f�ɾ�cz�����A��~q~�|�Ib���r�di���FnoGy���gvM����"�b���DIK�$��96��z؀�P�	��Gފ�!�ۂ�|�gg��nL?k�w��*�UT�㻧�2}^ή�y_/�N�`�H$�A�X�%HC^��lv��C�j�#���㻞n�Aɑ���A�P_����d@���p����O�
 ���iA�[�.�El�\�ka���i��L"D!��)
��V/��� F����Kf������7{%}��=���Q���=�b��D?I7�`�+�Ӆ��^��VGJp^n�T��v��s��s��=A�o�����gz� ��A�IIZA0ý�|8W��j��{n�ێ�N�p����rk3|��X�OUoʂ]mec����)�����4��K$�T�]+o�a���.ݐn���(�t6��	�P@~u�#$_X�D1P�	�y��1D� {�"��K����ϘZ-��:��	ӥ]G���sEw^��ܫ��lL�֦e�eˆH�d�}Lth '��ۜo��7ni��������%/��D���������w�<ͯ6��D3��`�Rܘ�q��۸��A%=����/Ͽt���2^́�j^��U�a�AN�T��!�]xW�ѠL�K�3/H��.&eZ.f^�wN=H��@�|Cp��!'�k�Mâ�[���u��� A��'2 o�LwB�]�O���&;���*��+I@��[lvl<�I��~G��(�7����(_9ۚ��&8�33S2���.�磮<|��3z4�q����={��լ�(N�T���gH+��V����R�H[l�診�O�&pΌUej��ປ^to�.'5y��fg��G/�nX�D��j>���J��GL�fLDx�jȝAB��+ �"�d�8��W�ک�{P�[��|3׼�G��+����J�a�=��YU[�ߓ�����h�cRV����	�[syL����u���	��5�&W�饾}$�~��� (-�{�{s�ҍ,sH�����7ܻz�/�� 3�W�D/�%"0�V��O�ؿ};N�;��E���qW[#o}`�� �/��(b��W��)h��2�;��$y�^�̲�2�bfe��}y�1Jx]k��m�_H�;%{�;��?fE	̀��2=짻��q���@!��@��dAf�kܹgޔj��#�o��2�U�*G�#����B�2R �a��Kd�Ӻ��ιU)�t�-����~�k619�3w�ǽA]q"�J�^�u�u��%�Ky��iQ�����;�3t\b.f�ҳ#�����Tݬ���;�Y�}:R�Gu�T�>�;��a~��?~���}��]������D���z��Ʉv�[�H��&�p�ܹUО�ŝm��<-v��f�N��y�a��B	B�4m�6�&U
J��ؗ �n��';��:n����u�����4�Yr��t]�۹���C��x4
�fx��w=y�q ��@&u��<Y���Mh$5���-A�,Τ��8�]7t{X�\0a ��:T�مjh�������va�͈�ё��{��b���t��l��+�a.3������{{}����|D�Ō�Ufs�W���9�d���sx��T�K��w����g�|AJ$��%�#��{�|������c�ϐY���'��o�1�9o����1��<���j�H;��&�A�X�����@�&��ff�Q׳6��hqi��X%� � �_`m ͂;�{!����a���A�>@w�K2�Vv��<6^�6e�:����#�b;{h{Kb��|g�"$�X2PD"�$C͛Ue�f��c}�4�6����|M��#x�|���J��Ib�?'�n$5$��z�Y�V*�QDZu��I��b���[]�Yj%n�A�4l��|�-����o�_�JJ��s�y�=����#7}cT�Ն��A�~� =�/�DW���F+���I.��>f��Xd�W��ʺ5o;������~�z��]d�ù�b��}v�Q=�wreP��7��y�g]̇��u��+��"m �o�a�{w�z̒���u�'�� ���O�;�U?'y���y�Ǻ����$_\�:^^��kV����/4A�<�{C]}���`��A$�~�!`�HL}�z=�����L���W���n͹���7{a�D<�UZ$�#%tP���ߟz���V~��R���_�"%{}�V؞�3־ė�{�q������{��u� ����������tVvo��!Gj�;���ɫ�j1MA�lˣ��`��4H+X=���?t_#$V��������َ�������ԕ�xP�x���"'�������(�4�o�|�URΩ���@��f޷�~�z�=��#w}`��:��.���7*K_u�`�0��r/�H�C�I,N86����˗R.d��P��A�S�OU4Xʂ��L�u��N���	�\�ྷ�h�×�}�8�=�|7VU�O�����y&)�z�{�0�_GN�)	�D��&�׃2�t�yC~ �a��/�D���^���/&:Y��y}r��Cg��!����~��d�&JI,X2Tg�㚯��}`P6֧^�ٵ^�����CKp �_ d��Plv��w�\����c}E�n�^{$�5a9l�������B�S!�{)HSL���}�m� ��"3!�fH�������U͇&�����S�ˬ�#slX=)L�K��WC8��V���>7���"�ͫ��<J�x�J���g��;�_%o��Ϳ��C�Ո���fhәV�s(�Q�]Q�P�n�3{���.�B3w��u�.X�e�̲���dM�p����=Q�÷���r��I,_�:���_w��k����^ ��"3���_fx]��72)[!�7���m>�t��勴sݻ��=v��45B���w��"B/b�<�uur�ғyu�o"{X(Q|D��y�㒀��aK�~2P@~�_/�f-�{�3�u�A�nV��1�x<]�����yY������XG�l�꬧�3UФ�q	P�We|r�=���#�2���Mf�]4v@�bS��y���?P~7� �u�JG�(/y�<�w���깯�uf��U5�¤�0���@ܯ�$��I_ d��]�����lɢ��R??r�=^�{fO*��G��J���ӬX2Wv���f��u �/�P��+��X �"	gU�Ϩ���9����f���ד�WA���?Ch ̤~ I/�+Ane�")� ���Y}@C�<�̞��n�Ϋ��wP��!���V}���_1� ��!@�d��2 !��;��@^���m=ؼ綺Mi�}��A,�DӬXJG�a��+�W�u��-���4ȓ����{�t��V'G.�v��u.�U�uӾ���~"��"n}x	x�t3WR�7*����_&�*`Gh�S5l�M�5ڭ�v����MI)�*(�c�-�V���c�.�a�ۓ�[�5x�e*�Ąqo.^�`�ۇ<�Y�v؞S��m�Tx�Y1LK�>��*��tu�m˻n���5�x(�����Z[����,�j�4�kBPK�(J�R@�!��e0՚�Mp��%�R�`�G[=�	��RA�nnP�#��_bb��r��&��/;�J�n�W���*BKƓGm�(g�����>}�|p:�~�-[��W�i��n)�CK��E�Xڱ[�P��@�8~C$�`�HA�G_�r�m)��s���ʟAg�������ҳ�:�����{�/�?	�	"�;y,?����D#ґ��`�$@IX I*��I�^�~k^{��ڽo��W�I �O+��)�>�-��P�o�ʙ)���^)�������t*�/z	�UY��Q�}%}$_I��{6��Z.�z�eɾ������n��$��"���S�����\n���ŁPę�"3�ƈ8�����x݃p���P�n�Y9z��å	"E���qo����z޿z�=~3�+'۞_w��$�~V�k7�fi��Y�q��sy�c�
T�>4�C3jr�ܑ�#�LW�հ�ܸ����k*��k:$(��$ȫ�hC�v����^�3���ɴ��U�roj~���N�!��ݻ��d�5��������"���x��U�{�7������_�r��vlΞ���/��	*H�=�m�k(��C�'��$C0����������^�}�����[t��X����W�zI�IBH���{����7�+�^�L��uVٛ����}���)"������0.J���h�l�5�M)��5�#��T���,g���xAF�<rl��J��0毆�_I@I{Z��?R~}{t��๷yo���tNr�J�H��t[�0i��-^����<��x}<���{�Tf��~����BG�Ǌғa���x�j���9$��y���W�c��3{���Dw\q��m�窔�7r�fmd!ۥ�:n��r'�t%:EմZ�J�֢OY��q񺣼�����dI����h����Fq,L/.���D��:����ޣ��hz��[��1�|��]�z��&��Z.�UJ�}utw0U�n�����n�d4Nw�4d�*��u[�v�u���U
�zVY���w{�Ӧ^H�{]qP�#�Y*��h\*�Ἣ���:���(<U����-<��"���eޅ�dV.橌�[L�F^vo9P-�Y`74�`��j_H�����E��A��o�&e�a˓��n�5�[�CEP��si�`��]Y��]��sx뾼peB�;�:�`恷:^�륲ힲ�έ|p��RF�Gx���hN������tZz�޽��3�'.(uIg�eE؇b��V	R��y�*��'�̣�g�;�$�T���.�	��L�`����w�+v��0�^ W/e��D-of�ʱ���t��_-��6r�F�f�>����#�h.n�k�2��LL�Td��@�HD6I�4�S��؛.�ɐ�I��"s�A�ݫ�q�U\�)�F�N�n��������k{Ayܞ�K4X�n��t)�X��wD�;��Db�%���tz�-�pq�q��q.�[��j�y%�WZ��{�ː�۽	]n��RظB���w��5U�h%Ul㪸М���ׂs��Z��b��P��7V�;I�lҴ�Xl�wr����G��u�p�i�M]Qo�]�SfI��T3���1r����e���a<'F�������ܝ!]��>�@��w5d6�Q�XӷFܹ��\劺s[�*�عr,cE��j)4QI��ni���͢6���n\-(�����F��w\Yݭ��W3s�h2lb��M���%�HQ]�`�W.�Z,�����ĤP�L�"d����K��B���4nni�S��*
�p��h6��R[�BF�X�S6�En�@�1d�;E������X��4�� ɴ�B`A�"����#PF����������r�mn�����:��}$_I��ǫm;�Q�wP̀31o�ۭͨ��w8Co}�uh��ʮ��V��~_}�r`E��$��Z�Uv1�����n��fm��e=55��/܆�)+�&#N�v����=��]���k��Ûٚ:R�;���"���:ݷ+^T��ti���ܸ	��辒)*��kr�=�������W;i�ʱ��k�z)"���ALv�/)�]��o�f����|�;x��}�@�$t=~�$���l����}=�%	"�H�:-��}WV=rsY�ݻ���!���}~��>_IBH��/�x�����yߧ���J�=济�~�r˶�y���Π� ��q�Ç�[ʸ<j�`pVq��a�d;oMd�d�5��J/6�M�}��ǩ�Ţ*/{g��޷�U*�D�K��W6�xL����	+金H��OE��u���w{���ﵹ.q|^o��Pn �_I�N�.�*IQj�*�]Z__Ȟ��9!ە����S��lZ�Z���֏���~}{����w�!��3�_�5����Z�~ٮ/tzd����A���I4IAN�ʹ[��hm[��o�"wmU��wq�D��;�o�<����Fu�A��}��I_I6���^��v���:����C���H��"�[�np�~�a�l�������}�ڞR/w��c����������E�V����$_I@I$����2���`�N�v�yw?u�ݬ�m���/�Pr $�l��fT�_�g
�䳳v�!�;�rv���d4�e��]&���]:���<��[����o���U�\���˻��wݰ�%���v1"T��Y"��Q���:]���ۃ�nk���B��e�/�h�p�b�WJ��Є�YT��;$�lhx������78�d��"�·���ճ3��,Cg��i��v��-���S�9x�c7���ѺAY���m�®xS�<g��a)�xe�Ya+y�J��s�30f��
��fX�5�&�,)4I��ee�ҳ3M1vl���S��-;�n�f�k+a�,F,05*�Z���т�91pb[!�AV0�{5}��%I�s��w�^�:�{�xW�����w��y}%ICG}	i*���z���9�/|�YX�����!#{��K��q7������& 31f��w��qR���)r�ۭ~������>���I�H���|��*�uv��˻��$\3��{��y�>�|�qH�s��p=� ���RP�r��U���JK0s���ۙ�$�X���!��BJL�U�Z�D�d�@�hp@�7����5�\٪�YW��3G�nĄc�v�W��n��r�8�U�+wֺ�ܵe��m�u�>�t�ɲ���?wv$RP�H�9�[`�P�.�'��b�9Mך�(&D"=�8,>�h�u𺇳0�Uqᙓi���SX�Vn�r�"���F���Jr����ڧvкS�oE�k����e쏶�	{������n�-oR�����_���LI^�F6)U�q���c�{��}&�X���s� E$[I{1�:��*�p��%e�f߫�{=][���֧xvnn�wI_a�9�MӜ�/��%	"I�O+�ׇ����i�o{�ټ�G�S����P�~����g{FX8���hOw:n�[�f�e�-.��u�[�݉`]��Е�MP!�ѠEի;W=�zT�}$C���'_�������آ��Ǣ����'�v $�MJ�h�.���7���7c��:��;=J*�����P��_w���2u�{�<�I�����Ռa����L�1m�^����]G�\֣"�v�;��x&$�����B��E�F�pr��J�e�J#Ҽ%B?m-��Ϳ�u�Y�~�����5�ζgsS����W��~����o����Q��3c�����O0��Wg�7�\bky�܁Ʒ��c����R��A���%|$�I	���ws6��	����<�˫kusx��o��"�I�������/_PcǑ4!e��]��D�6e9��#���,]�*jj�n",���Bǘ���o���E����]<�?:x�g=���fk�ʭ�/6*q]�P�/��|��zM��m'�"�3d�~���q��q��9'�w�S�wZ�^�wU�!�z��I�I�wt��c:�r��+��3]�k7���>������$RP�|k��K[W��Z`L��I��y�<�i�����߾������&�HW����r������VvP=B<���rw)#[��a�,n�\�I=ʯ����?XV���b�7;[�̞l�Km����+3����L���$�$��%$�ڙ�V���V������ϱ�7sý������fn�����A5į���]�ؼ۳�y�-=�����S3��sa{Hd���}2���$BJW�u^����;ke�ߒ���]����z�D$�	(I�'6���VG�돫uww9��5�7u���[�>�8��,�ۦ!W��Ȥ���I�;k���((]�E;p�gq׳����kꜾ���	"��(�߲���o�C��	(yƶ�w�K�۽�~�˾Ӱ��gC����t��)"�K���#f�b��os�zvOs��#���uG� ���v����J`��gr+�.��͔2;��;���A����#ڥЭ0���o��%c9XM��e�Q��m�]c6�&�����/���ΪuH�m�gꫢ��nZ#[cm������*h3h�^i��u��X	5��a-Y 	t»��	畂)�Rl���7�<�+����1wK���)��Bi]3�u�%k��E�p�Ons�y)Q���,����1�a��.��C��A!J�99��%D�,q�a㚻u�XV�]Zg�u���ۮ�;�<���P�b�չy�s�������D��[u�)�@̽���0c�R���=m\䧌�WF������31}���=����]T�������^O�yN��h���GP��n��|�%��|=�5f����}��>��$�df���5A:�|��I�	#|��wf��ݽs'��wipu���V���}%}$Uu�'�~�z���7�t5��fb�5N#'w#qһ���h���N�t�N1���~PE���g�|�mz���Ɂ����{N��׸�<��ޔ$�I=�'��]-P�B��h����9�쥎ך�Ǭݔ�13][ˣc�kn�J�龞�yHkk���3���[Mֺi�x�l1C�m�?���� $��@I̚q߷w��VS~4��6�*V��	;����7t�^S+�UQ����Qm;x�_8y�i�_^:���W"쬽*�G;}3֑p���q�g/ES_
z�W������u9t��xw�}���^v�c�:]���r��I�7�:�4`w��7����^���zPE$�<=U�%O!����_���������mf1���Ə������3ܪƤZ��k�$�$�I$���f��g�Լ�>W�G��B�՞�@l������U�i�'+,U�4M�APʅ
�z�0�B��[��[x����,H͒kl�CiR��.W���H���=US2>����߰ȷ���}W��^Py|$�g�Es/S��Z�r/�������G��l��:Pn)$�G�����v����%	"�I���ԝ�R�U�e��*�S�'QT��4�r�r՜�R�Ѭ������z��neM��^g�s����ۺ�#P�î�Pζg9)<��O�v3���g!%I�D���^�S�{=��^�����y�R[��BUWJ�t;�:o�RcC^v��*H��&���=;6������}����p̓�׀�@7�D�U5L�3(�9�=v7j��Gh��zCUf$K��Э!`��@�f�g|$ht�$_I���u����/�7��
���\c>�g{7��S��I4I_�9��^��ۀ{b���N���V7en;�ß�ú��F��T��4/k�/��}%	#�W�t��Y.������vp���׺P���� �L���:�����c�(N��*�����I�1n&��kևڏ��j��5��G���Wt��gr��c�S�/�u\��}��u��V�.�F���>�YQ��*��{0����"a��#���vԢ�ݐ�9�z�N_I�W�I�V罛�ݿ{A8;�{6u�^���߇����L�I+�o-�;v�"��V�"�3�Is��n��#ui��a�Mإ�j3=TЊ�s���>�"�7�IC�"�V��w�����R�9m{�*�M��P�_?y%}$@I��E1[[��빓��OX�^^rv�t��g|>�r��HN������/{�؀����M�K9�\�S�Y�ޗ�Ux�U�}�����I�!"�y/��'�bNCޯ��MY�N�߶_s�Z�-���J�J	<�*{;5�$@I�P�{*�Ks{^|�B�d�^�{=�]+3��}���}&	' 0�<z��U��5�4�zv>,!���U�ާΏ^�W��3���Zݶ��|�5!Y�P�K�Ud�8N���[z�Un[±c��D跫`#���`�]��]:��Ý�kL��X6뤘B�C�h�P�z�VWp3V�gJ�Q��7]ك�'V2<7�]v'��;{}I�Z�s�,��x���g�g�����*k�H���D�[��r.���g{7m�S�ge��7p[weo�l����|:U�&�~F�z\`A�LC)��׏�m��JyYl����!ZNnk,��gU,+k���:�7W%m�Y�v�o>гvR����kO:�/j��}�����lw]E0�8�k;89Ԩ��8O��wF��ҁ`3���U��yئEZ�꿝��e��Ṗ��=�OJfӗf�0�N3�B��om�7�$�,	�v�3�6�Wي��R�*��mR`�M��]���%egZ�j���w�س��oC�\��U&�M�[a�b���Sή[k��oU�컶����aG���w_�87sn�����xc[%����;)���r�ʊ���Yx.��������j���m�X��N`��Q�5qCw:������T�� �':\���[yr�A�&�|��a[��}��9����PZ2�r��K}�ΩZz�qda��TP����3{����;���V���=WGM�K�G����!�+;���N34�ܻ�pg?�ɇ9#��V�Ӿ�(��*��39�b̺
�ϩ��9⤅����0�6]b2�D#��^a�>$�� �H�I%z�lc&�j$��P�1P������Ll��PX�A�J$,7wXIQX���c]��1&CI����#!�)�bLP�b"�(�H��1�IL�We�2l��(���t0�4�BP�F��ɓ$�3L����$&��#e�(�e&BQ%�aFY����%1I����# � b�2��ɄH����S	d)3��IR	�g7c���DDi�I7cMCc1�A&��Ѐ��LJ�9��Ffx����8�g��=$��n�Zx�n8ݭZ�s���̴If�c�)-����1�����)Y�逭��We�2:1�ذY���n����b�Ѭ��]I�Tm�8���/�y��5v�>�pv��n�qv[�=�+���q�>.2��,V⎴%].��a.���&�W W/8�9Yi�a1K7M�m�'�ڤ�"��X+�a
���n�s
.Q�nͮ�S�u�H�Ǳh�d���T�!ݳ-q5��n.,sq�׈U�E�s�&�B�-k���,�ۺ�1LPD�%�
�j�Kh����mzձ��	�v�v�=u{�`c��W���N��)��c�],$28���׍��:1��E�8��c��e+�n�����y�6�^oCmf��nb��y�nr�=�8�����"�e6%�B��i���xz3�N�{Nh[����[R��Έ�!2�rL,m�i�[#����ѻ�f�0RSFy�ѓ�T�^_���]��E}����Ch�*;r3���wg��x�F*.Kg��v�`���B����k!*J16S
ۛn�+�l��:`�ճ �nzݪ�1��&��q-��ٳ�wk���/Ĥ R[ae��.%��v�Y[�-�s�;���W�`�ţuϮ�������''s�X���{6fn�����z5Pdҽ�eؼ:��;�7fN;g����N����W�e���6��*ĺ�����-���V�p�[s�#1��&��[���r�Z��H��M֞7P�6,���ϴ�X㙋�^-����B���)+���,&��f����wiB�Mc	�X�֌Iu�H�B�([wk6*�[\v��G�ѫkɡ([!����6�d�{�B���<]m��_lW-�����sa7=�Lt1hUdc��)[M�@�`�D��<���n+�s��40�Jb���.fAum�hLZd�#�7&Q��뢰IѶ��dRz(��{v�g%�N��t�[9���U�h�{\�r:��"�ӵj�=���o[9��u�Ia��3�1�:VD�ox�-�,��7��Y���Mc���ƃh%��,ʚjmKbk�i���	����`�m"��C=@��Kl`���n�+��,u�F��1[kd�Z�P��]�Lfm��1ֽ�!� c��8�u���M�.��6N�mp�.g�>�Y�_��a6��&��D(F]*�æ[f����Őŗt*�WE+*�V�W_狀I�J��ޜ�c��댉�΀vaxi&����q$�I>���{m��oҾ��՝�����I�V��k��̒K�[�M�f��ew�o>�	*H��Y�sS������[zu������;7�Z���fb�H��~��u}����h��^ƞ�M����g��߇O/��v7��տK<7���%|$�I�=S+ޗ�C�ebC<�};�ٲ�/��յ�·��$_IW���������6r:2�s�[{Bݭ�\Q��\�y #y[�2�(+�3��xC7��Oc��C3..kK}�V��������b|�jl}:���/��J\򟽁�x��qݻ��3j��)���US%Ud�{yQ�[�:�U��gF���[��5�}T��:m�!z�&+F��i�܈�*��{�}�/cV�V�j7�%ϩo�5 �̩�תӉ~WW'wb�_?rI2Ia{�d��V��q�l��,um{�΃rI�IRE�+�5ވ������_�Ks��%�ח8?{��^���J,���H����I����d��_{˲*�3_R������<��D$�����u�>���W����St�v�Imi6����� �k8��J&Ŝb��BJDŞ�{�쎠���Ք�F��Y��uG��9|7�	*H��+j�tt�x[�N��w�O��7��%�9��g~���՘���)ɥ^=��-�_I@I�E�{a��MU�]�4��Bk9�Y��赦��>R���5����c�sPݫ!�UG/;���r���r���]��O6��>uʻL�+�5��Y���@wPE��I��JrNV�5t�$�+���Wo:�ac�+�tr��܅*'fMBI&}$_I_I����m�K�+��5/�<������I_I6��;\�d�u߽���z7�k[f��P�^���mŽ��s���[+�d l�Bū�������I'���zg�x�L��,��`� s!��w����}$RP�"m�?JU�Um[o��;}�y{y�>���t��_I"�f�߷��w�=��!%	"H����KwW��s����2�����/���$�IƦ��������u���_fG�}e]׃d���,��:y�q<�e{ĚŵrS�w�+4�D�͐��}_#5��/����]\Y@�·%v���4uѥUL��N��l��^�.e��yui@jm�}y8l��H��C	a�0+��.�==����L�1����+��E���奉��������u�Mj��mf�͎�u�x4��sm��O]�*�J��}u����zI3�#��ao��]��{]�|O����G�|�P���}$_IC��_
�z�����۪J�˽���R���~��uI	�^�y�tz����/��)(I;ٻW��puS�پ���qd�wWVW�W���I_I.ySLV�gi1.�'P���'썗~�m\�76�ߞ�������<��u�^o��!$BJE��*:Y�z�.��|_���u*R��8��<���$C�&�55���ʊd8�LB�]V������3ê�*:S#w���2f��f=�ط������̭[�R��,R�����+�`@�K����2�C����]4���u\x�Iv��@14ٴ���%ݦ��p���tX���h�s-bV��C��ė7[�2z���9݊i��lͮ�=C��a=*e�#��&�:��*�VYH�e�ҹ6,k�fS]m��%��L�6�/5J���۶y����XL�m�Gh�*]bp]k<G[�]d@!�q
�ϯ_h�>�!Sk�v��4��nzJ'�m�!P�����aR	|n�X�����ro�IRL3������,{�6]b��/.��U�mR��/�M���*I$fT�u/U!�.���:m{�qܝ׼�g����&�P�~���W�PE$RFOwb��}���{)��~�R�����wy|;�	"�I�"ך�pc���.��H�W�<��{K�}��X�;�zv������ju	"IW�Nǲ�s��%U�c<�Ѿ-��x��;�9p�{܃褡$՞w���j�����}�����mj33q6�l=N����
]����G`I�ʨ���߼$�����Ǿ|W�^���~�:�;y�%�f�����+����I���-=fe�,]��^D���W/:n@�ۼ���g8J�^<��Pq�՜�y���t�gu.��v+0vj�ෘP����v��_c򬮽�yP۷���>��{�{��y�n��^�q	%a��j�8��d_���"I0�=�u���czd�Ւw^r����/�I0	"D=c��ո���@K�רfB�z�+!�l<��`Jk~y�3��
�y�B�E���C2��/���%kɾ#Q6��L��^�{�ٝ��$�^��n!$C���ޭ���a�	ƍ<��I-{e��띺):�;Kp��;f�z��RJл�_�K�y�}߫�"� ��c��O�U�����o�+O�o�e���������96J
��6��y��C�yf�{f���WL�F���Cޡ$��j�������� $�'�����+�T�%W#W�x�9��y�t6����+�'r'X����WTޡ�Uiy���S��-���n�vݱ.v�NK���7^s�{ٝos��j^�ܒo�P�#@�m��������es���>�3Y�d�}��A�w�}��͞Z��H��$����v\�E˨c\W�Rܣ�^�x��ܙ�����	"I#�>����5_"�+�l�B��Z�k�{e��͙��{	�N�GC��Smu��v�:t��!ک����s�छK�W�j��%�{�	</\k_!%I�E���<����!����h����"����t_䞱9����{b�׽_I�	�����v�fd瞩ݬ�f�����z�� $�}%}�U�VS�㠩{��}$C�W�o��[۪	rm^����"��[q�~��'�-@p�=Q�V=ݪ�p��j�ʕ��{cu�o�������`W y�N��T�������	�"�c΅6&D؈�`' ��oq|.P�!$_I@I.q�q���aߺ.��}���u�&3��!�t@IBI�z����>�����ka���J�ejC ��Ԇح�<�j����j��$�*��V)
s�n�|����B���r�u�Xn�ϵ�g�ȌڗGu�C��z!$�$���|$�l}%�tҽ�.x�7�e�m�^�u䑍+ӽ,�������@I_I�HF�[Q��]�}��mF��.�m�~V=�=hx�́��$�@����^�5�{�� $��^��l:�׎��xϷ��W� �M��kr|>�E%$RE&Z�e�|wV�8מ���۲�x�߀��� $`c~�Yۺ��UP��[�+�bH���Vs�o�f\����ˬ���*�S�(�C���yu�jN3w�.��z�W�6�o$s:��~t��X�
�������������Ⱥ�z,j,��;��ۡ�kϷPdy���h/Z���6�	�<�=���1�h${��n�v��*v�'`�:�rvu�Uٲʥ��Ȟ���X�L�k]
*�(r�c2�o#!îu6�G�੝�v��u��\r��cQ�]�u��"���m�4��]��E�����^[v׃�5k�}ul�39��~�/��ͬ!��7�uk���ys`�[��Հ�6�7�i����=�����"x�RHk��;��1�{�r*��=O�}��ɢJb�%��'+��zé;�����~��=���k�xdi��ֽ��8�D$�#ƍ�]�U�����o=ه&n��ú�n)"I&p�=�I4o�����ܾ�L�T��{׍�v����w�@_.���og�O5���/��$��'�]��ƫRU�=ET�^�|�S��]��|����" I-�/v]��^�v����yE8�J����j�Y�f��d�83;(Ly�dٴ.�Z��i+��g �!%}$C�V���ɭ�����TN�44�V���jd���I$�"���z}�|cAfÂ���\�Ő�U���Q�Ε�3��WY+U>�6GF�����3^��!�=��j��z-�:��u�T����쩓}����q½�z�z���wM�fࣳO�C�]���}$_	6�°z�6�(UCO�I���8�{�v���}����	"���yW�WLݏN_{�$�گvJo׾{��.n�����+"�m�������t��	*I�A�aVs*��}��8�ޘ�wd�{�� ;�������o�>~�5����YD�W@�۠/9�ʃY�7s���6�Uu`*VR�UVz)���܄�	+����U�W�wm�/=,"q�=�9~����f!�3�p����s��OD;}k:��ח�V��^��n)&����??s��J�/��}�b�Yf#�İ��?���V�3�y�*V\�6�2.�c�k����8+��r�U���r��~�d�{Zl��.�It�����VF5w�M��T�*[YX��X�t��P<�&��ESO�v;�]u�e�k���T컨�wzH�U�_c�ˆ��bu�li��UY�
��Y��*��#�,�0�x��;#3*>��������1*W�O�8�0_��,�K6�f��7\��K��5���z.:���o/-��>Ѹ�.1s���j��賢��!KE����t4��R�K���^�֫�*�b��Sov�W����܃;zuf^`O>uCL�'U:��z)����N��h��*�����`��F%�t�lK���'ò��9��a$��Y�={X���;�N��m��[	�{pu�U}�Q2-��n^�:��=�Nfc�Ts�"鍝�w7q�7U�a̺`�-J�"��,#����o8��,��6�"�7گ�g(;�U��v�\�F��}F�Ut�3R�@R���B�q�vmtڤj�n�T�1��uQ˚��*b��P1��#�5��Vl�&������|�%�C�����(�Je�"�pf��;+Eu�t����k}7�[�9��*�JY)�gV7K)h��7Y6ifu��gk-uAu�D��轙�KuV�0wN��Y��gr�n�]�,d	���9|��ڶ���xd��^-��)��\��x法�i�gv�W��aݬ�ے�K�_�Z̺o�B�sAS�fX�S��fvX��k����]��>\��[y�^{�6_<�
��"1(��Q�4@��� ��B%�1d�c)4S&P�&&E�$�1��`i" 	  ��&!� fD��!J��b�H�Q0X��(E��S2B4FD����ъ0FCIh,cB&6$ 1���,���0�H���!�0��"4&���AH) ����L	�� �TRl#���a-$�6L#�A����RF`Q��� �PE&*f�"4IA��ĔR�L,�$CF�4��L�Re�%3Q�LlQ�1b#b�\=��oU�g�ߜ癫�=�����	(}$BH1�|{����{�}�3��*OV%��7ܵ��މ�
���X��A��I@I�/��/�T��Zu
�kԭ��'���Sy��'Sq	"S<��}��S�aZ*����4R4�i�u�PݬwO\k�4ôn m\�,ƦtNw���M���߫�$�o�ߢp����%��ٵAx,����[ʹ�&	"��v|��<eb���H7����T--cLՕ��ޯ��ev��e%�UiBUVw��f;��Ȥ�$�է^��.��%3}�{�i��m/	��n $�I@I�%�<�GD���P~�$S4�K�w��얦	� sD�6+D���jT)�&r�J5"����x�>g�f�|<�>��y��Cϋu�>��b���.��ܙ���@~��A�Z�t�7�gP�D$��%|$��#���6�Ӥ�o��4�3�ҷ��_}:��IBr��^�l�*?Ul=q�yα2]i7e�ɺv�qn�#[i8!�v�(*$I��C5�{ᙉ�NM?SOQ�t�[ҽ�=��}C���{�"�J�)"�i��:�G���M�|���/�d�0�	�/��$�x��3��ϳ�_{�I�/��:;oc��;[y};�[�8��=3���[�9�	�$��"WޱB���N�,��x���I�&]���y��\�׾����OJљ�Ϻ4=(I�H��������w3u'_�__h��N^����ڃ<'��Ӣ���mҘ<�*Gۗ*��蝄ՠ��Y�#7�W)�MӃt�x5'��ΡWW��S9o�h�a9�o�)�E�
.߸��n�¥[�l:��YT��Ԑ�۔�UJ�/r����O��KF'k�GgM6�i��d�'�pܸ�㥇��.e�� 62�Q�퇐��D�� F�eo�a�3@B���W�r$�L:�k��6v,4�Sh^ea3���hZ���s�D��0u�S�X����J:T�g0�[z��6�qt�j�6x%���#�����.�Ͳ�m3�bi7�s�/߷G�V��>C\	ț�8·<��q�s;a#s:���;�]�R'���	"�N���O�7��i[��L�칩׀<��/��	(}$V����<9L>;Rn����.��q�F�z�1����KQ�^�}|��܋�辒��	#WKi�������w/K�}|��}=��褯��I��tvD={���st_>�$��p�pT��:X�9�t��z�v��C3=�O)(I�I+��Ϫ�����V����MG�5ﻫ���}&'��f�xUW�c�f�(�dqC���M162�`�&*��)��K"��s@t�"H��m����w۝r�z�<c��^@zj���H���(��mڊd>mp�E�q5-Ϊ�7F�u�$�}Ǯ�������$X8�*�� ��[5��	`6���T�)X��^l@(�A�V�h��^^{��C�s}�@wW�K�E��1^�7n$RI0I��{h�~����]ҽ�S���f�>�9�$BJ� �Ow�����t�~��������ڑ�b��^�d�˯9������E�Qh�J$o����` �r$���?�mȐCn��'B}�g�Ԃ�ov������WEZ�A8�};�/�mI��������y��u/�L]���9!0�4��.�#�#��R�LzN��eD�%(�S�ބ9M?^l��}A�"{9�����J�N%O�%�C�l�UwT�������~-��k�-�$S��):��*�>�R?�R+,Uo��{%\�q�<������D��Ǯ�/Bu2.9cY�'�6�d�CnD�r'���P(�>;�G�����*�S���j�u�UY��y��QVd�wK�z�a�3)���"sq.�T�L�Yh��i�f�T�{�i���J}]k� �m�A� [jA�ԂHNޖ��<:(o�!�G͹[�6�w7������N%OF%�O۰�g"�?T�Ȭ����m� �ڒm[j��u�g�V�U1U����&��-�x)���!$=hIn>_6�P�z7#U��޽O�{�~J&�����H�/ot���kcq;�f��n�Ā�$(1t=�	ڄ!�Ȓs?7u�m�n��-®�����~���5�z�/����#�m	#+o>�.�.�1��� �Α;�!Z��\�צ1S���� �ClU_�4ڹ������ �h"�@6�&j�me�shy�w��=s��:&y^��uȐ[���n��~��j�u1���G��I��O���ۺ�}p�N�����y�Hy]���i+����˺���B3+�dJ��(b��}��iwc%�r���g�uZ�v�N];ܶ^�-:sx��ԃ#:��ܺ�ެ2�z�����Á�jH �k��m	���p~��؊��"~�<�s��zTԙ�O�Z�^��ZCng��hu�e��<��U���:m�d�#f�V�g7��wHWg=�%�@&�fL�2dD"'����K�+W��rڐA-�#��ݾ�o�g���<&yn��9~� ��hH<� Am��,��44O46�u�$z�}#y:���	�W�޸f����A��� C�-�ٿs�V8d׳��Z�@@��Cm|�}A�"ht����ݙ^K���;���S��A;��Zm��@��k�ݪ��q�=Id�T���܂9ڧ�~m�e��}~����n'B�@����+�T3F;�J&�tH;p��Cn~���AmȒ}|�m�
�����{_F>��u[�iq�\�9O������	}ʗ�+�*״h)e��P+��̌ii��ː2�9-����8s:���-�]��?��Җ.)ި�]ޓ��T<{�9O�Z��[��0�ek}�վ�� n���t�ۢ��	O ��:�n�r�:�^-�[
[)[�����ʐ,Յ..xZ�d��d����&�7c@�tL��z�5��6Ѱ�����G;u֩㍼&u����W	ۻLJ	oB������|�w�"��yhk<�,�=wYӳ)�$���L��Vn<��ͣ�/P�]f�)Y��!��Ň���>p� ��BE�������,c��.-��h��S<h�s��4����Rb��gBID(�?�������v���͹�U�s�>�x�U�"�"���ӛ��(�y�$�ޙ���-� KmI>�����Xh�������$w�OՖ.�m�x�p^8�08�B~ ����Tp�t��c��P#�̂l A��"~!�����������4�\֙Wv��.7k���H ��m�[jA��� yq{�Llg_�߈:�D����ݑ��i���`�Ȭ�����wF��l��K�=���4-� �m� ��͵��LWosM`zw�|�lUV��t�L��q:&yn�$�vD�p��܍ݵ�bI�������<k5�{<�TT��!ZT��1���bѤ3�,{
"D��&"�z>�}"A��O�6���l�Ɉ����?-���D��`WF\yI�m���Rm	m����[*�s�3�S*�8>��&rl�}]/xjT8�]��וS陴v����&Y�>캳��ѳf�ٜ��2�=�38a��~}��q�܎ᒝo���{�eΈ��'��_E��$6�����w�o� x��H��@ ���ԟ�i�ӻ�٤j�����jtL���$��-� ��H!�2�;����{Cf܉#��~n]�n{d�Uo+�~[qk�ռ�evr�΋I�΍}�H ��K��A��"Kp�݀�;�h�y��_�v�xtU`��s�ԡ�v��odO�6�~-�W���z+O�����/�v������' �OO;��t��8�ү[/
1%H�fO��<��wq}?kA|[jO͵"����v�Ffz�5<&y�px���Y�O�ˏ�U��f�fYb�B#���#�裵>cH�k��]v���DҫܮL�q�]� ��_N���I3Z��'z��=JAi}��H �܉��&܎�7�p�f (���߁�W���4�f��т��>h�Ps}q��uT�>�#u��XC��^�a���f�õlM�՛���X�HC͑$6�����-�$N��_�����5?Am�˚�u���f],s:&y�|АEX>�$n�������H���?���Cnz�#~������Ƃ���ov�}*�k�f�����ܧ�7`/�m �Ok���D/�D�	̈涸�vll[��rZ6��%�,t.u���!��N�����rA��dH8�|A��&��{�;�¥�<-R!�����Dq�	!������ԂŶ�q�*̞W$UXp)��_Oǳ�;�C��;�eg�_�B���B@!� �r�
�2�1��Y�"A=Ё6�O�6�~n�i�y:�g̾~�zU�t�5�7K� �}�~ ��[jO͵�t�oZ��{v /뫑 ��B{�ھO���`禧�/t�^�"0ch���E�����!ru����ӵ]�v��RP�
�]T���v�T�]����_Ld����N.x�Nd���
��p"�ȟ�4Ŷ�����@��%�G����f*ݣN��7���d�N����	�vD�[��mȁ�����8�q)�͝��a��ڸ��woG�獩C�+�F�]�]�)���ù���^�!����_g_���'ҫs��5�7K���G�v����;  wZ��%��������ב��/x��@���'�W���)�p��H?��#1Ȓz�U�4,q�O}`L���b�	|Ԑ~mmH ��I������{F����WYw�Y����}�/�wvD�[�AmȐCnd{��<�nw'|��^��p���H#���m�o�}*��9f����A�������o=�e�Ϗ������t �П�m�%�kϣ�ncS^)�o�N�W��ގ��H?���� 6�~!��}U�rW�Z"iI�Yb�nDW���L�Q�֘{S�}2M7]U���b�r��e��1�ݧ��w��&��*����TS�-���z�jkk8�:ҭ��ٕlTeS�c:��<ɓ���;R�(-�6d�w���;n[[Oc�pf�D��|�V��Bf$�n���@����L�jq��9�k�c9;���������y�uN�tP�F��X3�����ݕ,CX��8f�ȷ�K�z��"���٘!ʚ�����F�6z���X#�Cj��Ϡ͆�J�]�f��5���3!��fWVK�wb�N�[v,���2�g|���zlk�:ﻒ��4p�j̉��h��ݛn�Hێ���X�Ͳ���DA�J�|rgac�baə��:�۽��:�˼:�f��m��޳�\���.�*e�����~=l�N�n��tVm�jm����]��B艖�?�ڭaGNj'B�N9�N�M��ɑ����N\{5t�]㼍^?Qe��*��Zrd�ϵ��յי�6�j��S��������'[u��4��w`S5gkJ\�(uۥ�Ɖc�2���H֐�Р�K�)���j'�ٮu3����m>��~���GYܭ����=u��ݗUt���=�6[���]�4��g��u�.��;�!ݼ��3������9�:s{9%m�����@spV}Wc���n��!.���WS/V�]{U�6�ȟd�'&�Ꙇ�Ҏ,�q�B�7h=��p]L볻�����/;wt�Kw.��Sn�W�9�R�ȢB0�̣D��"0L�����R�D�Id
��e#B"�%��T�E�c%cQ"b�`1�I�T��$���bJCY��M��Lf%L(�!&	�!Rd�#2�Г-2��DE�ěD͐� ����h�3I�i$J"bB����H�h�BPb�ĈX�F(H4TJl��B5��5&CI�lZ-3d�a$�h(�Di&6���Ib����!3X0Q�	����lEE�)(���,1�`Q�$��Q�����b�H�EEF��ьcy���O#r&e��/f��ri\v�b��]pq�������j�k�n�����kh�é[f#qH�W]��ViE�E6��;l^r���7=9��S���N��nn'n5�\	r�sll�ƍ���ٴfa�5�a����R�ڇK��Q���YDa)z��0v%�k��Rn-nq\j��� ��m\��Э�A���GX&L��&֗r�z�nԆeƑj��Jh�Q�ݢ�
�`»���.�-���J�����4�V�MWzJ��D�:,�l���h]�B��e�Z.��m�&ݳe�0�!�`5f��^e�rc�����ې5;!&T��0՘Ucd0b#
²�pm#�	62��2��I*E�L�b��es��j�Yn�a�-1���%��,�PD4�kIJ�;J��f%Bk6tr������.th\Y��N�Ng�CU۳�z�[Щ��Gkm��l�.���^4t�6���e.&�6c�y�]�Nd9��7\b|0s�Go#2�>@v�;h���x�� ��Ƒᶹ똹���[���y���%���E��u4[�/V{�A�n49,2:٪�1�,3\a�#��g
}�Am��;oQ��ñ�=':�%*�3f����[�n:̓�����`�Pa4-�sk�Ѕ�vw���n�eWEԩK:9����󭇏�����9��I{<�t�n�g�M�6M��k�nrFXp�MaA�/m���_j�j�z�7%���v�	ve��As�be��0�v��R�/=t�pb��f�.�v�q�㞑2)�ь�M�P��!���I�D5�jX��aB�EĨcGgN�㮠wWnp�(;�7��n�x݋��9�x˦z�cO/Z�2���u;�۳,gu�q�]�Gn۠l[�x�nW�ڽs\���[Z2.凵�9OL���<>H�9�(t+����6/bF�[�מ������B����8�!�sg����e��B�q�1��M�t�N�(�bԛf��y����F7,��t�Y�4�8�rٵpYp�l�t��R"Tį2E+�XQ��	eȋ\���X�<�Mm��|'V�"quԡlӹxp����T)�sc�uBZ.�ŭ�3�M�=��ɔ*\U��x�T���O��6��j��ٮwH�q��]�fҹ��0��Chf D�v��Yma0�nw����l��GS���8�������k�i<M��D�;"�� +�;��ڢ	m���y��d��~�p���뼈�A�{i̑'/�-�CnD��/�n�W<���F���熂7�?��6��>��|��W���g/����[2�/O�3��/�AsB~!���[�A�"��⹔�r6���&;7/z8FWH%�"�r$���?�͵@�$m�l���_@Gw��KmH�v�5�o��s��5��П��5�-;�,Q͏�ۛ"A����!�"A����g���	 ���6{����uǫ�)}��j��!����[k�3|�yv�r|�>��>q��X�`���.���e�5h0f���!H2D(J��m��9V����p� ��O��mV��Dm�U��]#�{���ˆF���Cm}-��k����s��1�1��K��^�P�Se�
ʜo+U��&�Dܬ�����[Zi�wf�����ř��e�Z(ͼ��7��P��7	��]���)��S�����G`�cu>��_v�$�5�-�0�<�d��í���7�~����@6����,dҸ�>�(��жۨ������Z�W͵G�ڒ�v&U�{A�~�A�A���6(���.=NOl���1S��=� �����l���y"~;��ڣ�mI�m�{��<c��cLkR�q��z���GW	�hO��dOŸD�r;��
�Q{���!�&{P�]c��퍘4�Q�7q���ƣ�-�-,��/�}?d����zY}���<k��?lż�G�^�F8�m�.)�`ը�U�4�ڒ��z�KmI����O���&�[n��g��l"1�;�����&_A����A{+�"@!�epɍ3��>[A͵$q�Am[jH%������E������^d@����j��x����f��zo�,.1A��(Ң��t�'�;���t��5�^��WD�'���x���5��f�@�{Z�wdH-� �r$�܉�o'��yw��!�H�/v~��mw�F��V���]qK�'�T�<'1�0�w�h5Ԥ�sZ��6��[r$�f���>���F�ȝ�_�Q��6������O�a A��Cm}!�=U���r�ެ���Z�.��Xf�t���=���d�m���n��=A�8����������?����jڒ-�#��_���c[�\*�*�P:�u�_!����I΅��"@!�"A-���Z��(s**}04�]��Fj��Y���o9X⫍��ݚ�PE����xY��x��*�_chH �nD�� A���\�T�ُ*�0Z�QӢ�S��������"Hm��6���y�"�+go�ET}���?6����y���61�3K�ͯ�� ��%�����;��+hZ*�֖M.�[W���D�`Oi�e]��cm���R��t֣�0��&�]U�C�\�qLs��[����/u>o=���O 31-�܉���̸�q�=����z�"}[�V8��_p7ܤC��ԃ�my��&�:�	$�O��&����j�G\a�e����j��9	��ֽnd�3�	��$��g���܍�n�Et��a����!M���;F��#�dH#9���-�'�ڑ�א�.C?{�Q��H'�T�w[�s���[�f�
�@��	 ���$�WVTi�L��J��r'��@�ېk��w��븙�h����+���/zeۚ�5K� �{9}/P_ڐA�ڒ@![��I=���!�-���}_6�H��A�	oFR��簈�6v�ˋ
"z�1�s���_7 �s1H � �̅B��4�3�np +Q�zd��~Μw<*��/��Ȑd Fd	���%/�VR���SNі���D�#Ki跂��ܥ[�]J�%{�a���oi��x}u���3֨3DFf�U)^���8|&���S��5p�ٹu2��)��:�����e��%�J,ڸɧ5��I��Z��"��we;YQ��k�5�Ç�&��c��/U)���k�%��é+�/;@32͈p��h�9������)�Ҍ�b���82�6S��"�l��^64y5v�x�gc%�6rmj����0�v��	t���4ٕ�q.��|��P���`1�ҵt��Xk5��Z�:��Ʈ�v�ŹFOs�H?8D� FfL�Fb�v{e��|oB�o��5E��Ry�+eYٵ�>�D�T�W�s2�&e�#�E��^2*�Wo���s�p7P�-���czt$��2|tC��qq��W�}�Y�}>Ԃ=���辷_+�d�]�*���<���Y��^�����ȓ�@�A|Ff!Y���ٓ¶b>�@�E>_H�A}�r��>�es�.5Dc���D�|eb�������8�U�~=ܬ"%A�Ib�����fӇ�j�h�A�gE��;'{�2|xC�z����DI.�2 �d�e�}������\b�͘/Q�v�;��3c(Y�ۛGd���2L�q��y�!�s!��b����~ks��bvϫ��������Y5�}E��w�4�b32�34h\ʰ���W�xP��&�V%�dzL�x*��E�v��e�������&V�wm�c�Uh�l�˳�;c��<C�Spp�S2u�T6F��`͓�v�-U���}"~#Zun��M��;Ηz#�=\���s#��#Ƴ�Twey�
5mI��Ǻ �d�21�f͕ǌX3#�\����d��j�	�v^���ɟ��_fG���9���ߩH ��A�@�1H�ݽ�5{��Yn=\=p8��@5�n�[&�G�:����T"r2K��J@�$A D��[5m��}@[A��OI[cFL��Q�Dp ���$r%|��n��4p�_�Ŀ�B~���9�h��s�]�w��u�'z�鰭��.�f"feh7?@`�7\�2 � �h3�[��������t�����#cHw <u?f@_�D��A�U*.s�ܴ_�: �mH�{}�w¯�U��>n ��"Nd\l{�""{�b3@�}��=��̲�ff�D̳��w߫��-��O36�|l��f�]�U����F*�H��G�=Tᏺ��Ѵ0�I�x:���DP����;.��Fߺs�C\H���O�Q�%ܹ�eW��{���#%"2EdH�0w�>s��&:�q�5["@;���=h�̥�8኎���A���"9���>��7q����@�H�d�Ȓ�2V��=Z0r��^���__F�^���E� A݀�f�s!s�������ah�^D�G���|�Z�a����,V���!��z����c�A=p����?�C��9b�\��x��a�y�:�8r�Z�� �{�	��$f%�dx����gy�cD���g �����\��8�H'v���fa磦B�1��r�@�w9O���d}�f*��fGr]7�;�o�.��d�\)r��@�ք�s!s@�̙%����?v �"��O�f ��z�XI��W7��Q���;�`zx:�9U]�$��R�)O����I�����MO��]�uR�
�l˗e�q�ڃ��=H��L�9R������B�RD����">2S��1�:��1�����B��8�	����#3&~#1	�A����{��Ӂ)Z����3\/f�<�
M������3ƽb�r��'���.��|�9���b�׼�:��]I��.�R��]����O& w�`=����$�% A�d^�����"~{i�T�+`W~�w�����A���מ~��.�f�I����d A�w���Ϥ�r(�\g�[n~�����})�H��G2�(�Ab����b����A|�\"9���ޞ;�D��fIu N��"��u��Y�8;��/�#܂I�d�A�D�y��ϲ۞_��+��.PU]��G��"��+��Tw���RAPG2������T�<��'�"R�ۥ�T���Z�׃3��T8�Ww��س7e|BM��o�S�I]��+^�3��
T�~^�=]i�ݏIj�F�hFk�h�7f���8�s�E��p���Lhۡy!�uń)E5P��c]�n�	��Pnx׵�$�z�bJ������b�&.�$�R:F�����*���<�CR�ݓH3 j�N�L�Wnݞ8�����F��9�������Σ�g�����e�m�S�@��PsIm-M��.l�qT�����h������Yg�%��Ÿj�-��r:Wz�l���A�0�`[ ԹŮ��ڡ���}b��� �"�7O��d���g���1��sdºذA�:���_fG��b��fb��s�����+�P|���[�P�c3$��J>nF�"Ā8���ى�;�N*8rH
�B��� A� FfL�s�*s���y�@�KX=y�
*ӧ;> ���H{��	�� ������w�/c}�/���?^EFb��1w�Q���q��\'��_�Oi?Q}�P"}����d�~�/��FJo��ڇ�<���eWwT%i�x��K��[B�̄I�bBs�{Y��q��}ij�KRƪ��ʱ�����Ք#m���EF�p�١|ʸ��)7���-���{ǝ�k]����J5~;{�~[�>� ���3�Fbs ";�h�w�����SדD$��Ÿ�L�9�z�V�Ġ�+����\����Q��}�6�̙��ve�����N)�H�-�Nw�k�#��_s_&�tG
���p.����"32��b�'�x�� ��j ����A�#��_T/g�z�v�eu�7*��:�K��|A�q�ّD��I,X���92�yӎ]��J_�����"~?f ���c�[9+�#��ۜ��=����/U��ѿp�'^��)}�s2~̇���C��fb�v�1��Ep.�	��"�FfL�Fb�S��}_c���;m���1�l6��<'N�i�XM<{�xPT�2�H��(�S�ƃ�y��/�d"3�n����o�9ye��T=:x�˺��n;����"$�X9����A����բ���􁸇]���� �\�ƶ&8�w9};�/�d9>"�/����q�8~��� �">E��t��g���V��P�������SA��6���%z1�].��󹽯�9�V�a�*��Kw.�yY��Wj��ّu�R�BU_G�lUZ�+�&�R����f���Ȏ�W[�	˗��[Ǩ�t�7�l)���*΢����`����n�os$�v�۲��l������Q��3ԖX����T��QkP��1Y�{Nt�]�l��ЩG�wY*��j#t�εp]��Rgt�+:�UtQ��1E+�0�ڛ�颴�7-��]W]�C76�,�U^��w��M�&g�:{D�fֱ�"Y��gky�A-�����mA�Κb$�5�Af���̭ojl�һ/f��s^%Wu��M�9����k�2��Ȇ���4����v�,�����U��d�z���v�*\�tv��fl���nA����;�|e�_�	�2��sپ���La���'fw.or
���:�+�Fn�˹P����tX��]ٕO)��m
L��I�
[Usu�o��ou���/�7��{�3��Y՛�����{W��7��p{s����nΝq��vh�WSJ{]/jbq���9G��O.��DY\q���Q��9s0Ҹ�/�TV̪�:b�:�n�O,^�S���yL�MD�\"f�V�\�G[�i�ܽ�ά���ި�2��Uǭ�mcbz�UɎ�ݲev���k�2�N���}c�*}B�Y����m{χ?ziā��𗚭e*�n���M�kwEX�n̊�~~�Vٹ1#l71�M�.�~�/r�¹\������X��,�E2���2�Alb�(�d�Ab�X�,V0X��`�
5�0���b	
Ʃ4��E�ɋ3�&�X��FƠ�Ѡ��j(��c`��#��X�FjJ�E��F�TEX�T����ţ��4���5�X�Qc3F-��0l�E����+FȚ��Ѩ��l[�����-�h�b�4Z"�F��A���Ѩ��(�Rh1�Ih��i6�ڍAdړTaT"���)�����UV�}�ȯ𕿯���� D���"�H�����O�^��ˁ�����;ٻ��|8?^M�Ȯ|?����z�|n<�~��K���2 33�M�=b����;��ocnq��q�1�����̄�b��9q��ʛ�W�%#�	D�0D�����ư�j5T�[y^�%oXh��5��	�m�=���/�d@F�'2>Y� �ͧω�{��S�"��Uu�z*黏��܂!� O���d{�9��/��5���n�ݽ�λ���1^<��7� ~/`/� f�s"�t��"��#7f~�و Dq}r!!N�>W]�u�x�����(�q9n;�;�	��$��d{��f)f$&o���K�\#�@� ��"~7��d�f�������te.�A���8�.Yh��۳3Y��~�?%��/"�c�ͩ������i?o���[.O�T���ڀ��h*�Y�GTl
�<��~!��b�?tA)L�YW� ���9�M,�ǹ[��D�+�q�| ��3dĪA�AD���c������ީ�'ݶ�J)�Ԙ�+ez��j&DB#�"�Ms2���V�+IzK��k/���W�l33�Ff �m�1۷�.W�_G|D�A�ګ�;��_�E�� �\��4 L�K��z:��w{�C��ﳟ��̉�r�	�����fd�<����,��r��w��Fb��|d��{W��X�Vk�~ܝ�ܭ3���b=�"w��̯`��\35�~w��ط�Ssz�>b|�Ss?���}��=���m?\>>����������I�߆�g��/���fYb9�Z&fh�9���vsWw�/=�1������ ��<�H&��#3&~?f!Q�9į�w��^��ū1퟿6&������-�wT��
���ӓscm;�%�����]Ю�\���Ky�!Pq�V9�m]���K;��}]u��uuv�!�����z�Etsn��:IL�� ��,n��C�c�H�k��|�a��ގ۫��R$��)�=��^�=�!�S��(����:�Vم�<���[0��m��0���R��5R��f��1Z�n%EN6g�K�A]Ž��f��%�c*�Sgm�D�IW�՗ {Z�Кk؎��]��Z�4}���\*�%��u6v�k�퀘y�b�C���iPw]2��%Қ���8Aε$nGّ� �R�7��ݙ�f�^;S�o������6�K�A=��=Z?H�"Iw���̼�ݏM]S�R��u3��
���S�Fr���p��p��_Oۨ#���*ߟ;;�ݬe�ǥAKd��D1`�]/��P���T����9<��]p	ۄ?^���ɟ��1d/�|��0��+ւ=о ��R7q�NӾ=g�ک�u��GD�ڼ!g�Wop�w�A�!`�H�"$��]�j��TBw�?D73�9�s���7M�;��^�����H�����V/�~T	�HѦM�yh�Մ��Ga�&X�.��h\#bB���K]��W�1�(�7�ʸ��e��7�:L%Թ���s��v�3��FG�u��H���%"2Edz�}]Bg:��p�WەY�Lo��.�,�w��Y6%�w��k���Rm�=�*���Я6���5�|&�6|��Rl �p=P�?��n�oN�nGY�mT�����@~��O�2x}�\�?J�/�}Z����T��"I���zE��4�-5�=j{1��L�'���c߹z3�[�A��30���ì��u0��_=� � ��;�|�Dr�<%����A ��!�Vt���ަ �џ�[���?/�����+"J�O/v����=��oU
������^��6�O�@�w`/��П�d"وP�����׏���+R8��)��2�aV(K��4\�4mĹj��ι�k4^wo���u��d������~̀�ՎK_o7>�t���3;�*�O����8�[�sA ^B?fb�3_f@D9�/���Q@���gb����7�)���t�u����ͻ7�qk7Q���B��K�;<��(/����H��DRM{��3�	���	[lb˥wlv�F���9N���*^t����(t�.C�h��!a����8:�r�&��j������k��7�5A
�wY>�m��W�k�����D�"@9�� ��]��=����~�}�Z9��?f!^�7s;�<�];Y���o��'���Z��x�w��D��3���"�J<^C;;�
��������߸y>�]t��"ר"32D�~|g�^�	��g�g�ͬ����&�V�Ob�8'��E˦f�km�1��S�w���e����#ud ~�Ž��gw����;�>�\�Gx�Z���J�@�A���O��/� f ���	̏���{!�J��c@#ΤO��U����Mϯ�y=����g ���{�i�́x���AK�������ʳ�?>h�;m���~&�O�8��N�|�P_��'㘂9���
����� �/����	��/r�N�o7>�˼3<2� N��ͼ����ǎ=�-�T��������������_��.�y�9��S��cczw��X�����I�mY\r�S:V��vy�>kyi|��>|ʝ�33SS2�D �B��.���H+�W��ߓ�>�����A���q��9���b��^bӦ7�"��lUʙ.PB1	X��F{N���spڛ�,�Ʊ��a^]��M�.w��ˀ��D��d/�̀���r���4�k�Et�y��p�F��>��P4�y"~̀�d ~���>��SKG�n�G�/��֤v�s��FU�<2� N�"�Ȑs#�S{s�%`��#�g���� x��_Nb��$�����:b2�;S�~���ʣ��[�A�h rR���Y/�z-��T,����ZA�(�̧�o��m�����.�������u��y}%` �$V��̉[=�Vne���概�p�{��܂��C���<���D3��ӌʱ��v���f�U��%����ӵt�N�B�uU{�+;gT�۽F���bTTF�ę�6�gU-��3`�f��w��Π�TM h���H�E�Bq���wL��6^u��qN��\��y�Ė7[z��}Dr����M��0BYH�G)f�X�skf8�U��rJ�bS�t�;'��8�����]����y;���&�l"#a�+b�v��-ḕ�;�l�fM!��C���є�x�3RЂYj�V�רK]u��rp�;��i4	�5uJg �)�m�k���B�����6LM2�[������T�b�fɡ�0.� �k�Lo�g�z?βޠ32���O��B���s^j�禣���+}�倃�Z�~��$f/��|F��X�Lu��\}��L78Ɖ�ȃ�&�e.;p� ���yOc�J���I���ӑ����ِ()|A2E��O�x~p]؟��b�f�O���݀7s!~�A��"k7c��ڃ�YU�}��D^��?���턳^�>��V�zj8���H*�ݾ�!��|y�?9��"D�J}$�fJ���cٞ}ŉ�"PB:����4w\AǓ|WH �� �z�fd��� �f���UQ��L�"%&$B���m���g^=K�r�P�0�[��0E��(��_�}����@�B ���~�����w��ʼ��+��x{fV_\7@g��������	&�`���Ñ�^L[Wzr�Bu��H�|j�٧�q9��o+-}״[�/�d���YY�0ul�Vs��N]�TGm�ʖ��)!!mزi{�.������E���/�S�Ks7���5n�f��'o��A�ّE�vnnV]>���/�R�@D��,�_/�B����N������_��F[��r�H'r"�"�&~̀�d"9��������;����~��/G�[��b]^`����� �ak�*u��2	̏�by�;���iyTo)����	S��W��[�٨�~�� �5�dx���xO.���Qз��0�%��.�q�����q8k�%JP�BͶ
���FD��� >�e��2(�3.�(��u�����s�F׻2%L�w��܂?K�� �2PE���O��j{�ĝ�@���/�W��3b^^`S�+�'�A����(�����2m�{�@�D���~��ْ��Vg�!�)�n�d�{?f��o��*�	Εa����Wۚ
8�ql�/c;�QB�����8kMeY�b�3{S�V�ܔ5r<bܬ���tۉ�z�[5A;|����+�H��$Hn����iҡ���'v>́����Ũ��no��/����a�'u���/����?I�s@�Eǽ�1��;�9ڧ�`�����n����p�D��@�3�������>J]������4thq��y��p��5P�Ǩq��=��]�8y/?���:㏝F���'�3�Pީ��s���e�[>�{̌��t���>���� ݠ�?�K�	�+!��%A��HZ���,x�_m�Ep�ȍ���-��9�8���^����]2+z�ܞ߲<�5�w* � �̄��}]ϓ��2v����	�y�Wd:�"�'21���{\n��
��`+� CΑ?�+�:�w�sS�>�w>���v�I|���܇fb&�o��Y��*���V�劔͚�6U�Wr�{�	Z�N�����b��N�*�)l�e%F��\;�� Wr�Fb@��FfH�s!�u{�6=:��(��N�/��_3��g����X���.�X���|����v{r�s��M�ꤔ1(�p��X�ke�1�"R��O� ��)��̄�b���~Ӟ��^����<�{9��a�م�z����ݿ��AD�E�d����y5[�>��x�[������U����k/���q���A���A�� צ���OFv.�A��${�y�D�2~̊ ���	}���_�>���90��ÚV�U|2+��sa|7� FfO���A�u�I���$���x����#v�I�y��g�������.�ҧ'ד�Ws,���քs*�2�30���s�D�E��=��kW��7>��C��A����ʛ�hE���B	'��6�Ŷ�Z�~�kU��m�V���kU��έ�����Z�m��֫[o�mj���6֫[gﶵZ�|��N�$�$ �{$�o���kmﶵZ�|�֫[o�U���V���׾��km�m�V��$ ���
�2�Ȥ�֐���������>��������                      4( �|P�@
���UPP �v�ƅ� ����B���
p�GZ� W�|��� �@}�� Y���P�᮴ �^�b�>��Zwx᯦� �υ�����:�]ŀ(S� |�UR@x��Сqb�
w=�뎳��z�����x�y�uv�>�v��x+�7l�{�`�a��� (`k�f��/�;�x<�w�M�s:��޻��u>�G ���Ƶ&��r5��zm�� i֌
})直��Z(>���z֎�� O�M�cA�@ Ӑ������      <@j��        �~JT��H` ��4��O�*�'�R��a рd4�0A�~�P��140��&�C	OH�j�H` F   0 B� �M���D�Q�� ��LmI�}^���}{}:�ϠPN2��`��"�{���DE_���&A3���щeUQTh������}?�l?��?��	�TLu�PO$L����)P��&��վ1޳�,����|���ʨ('?z��`��2���0���Aw����� �����6�`0a!�?��|yɝ��׻�}�ǐ�*h�Ľ�.��Cub�ړ9F�3������W��=9���"�f�Џ�l�O�^�B�D�2(�����h�ܰ�������,��
cͰ.�%����1��-j��Xt����b�{8����a�:��p�e�{]�gN݅�y�k#8Zu\OåRP�<\���=���;;��t�9�LC3[��ןNn�S,<�LwkӼ;6#6��}�(�}\
sU�@����g���ŹD��V���M�޽��Djж��g�Z��n�_A�>x��ڻ�;�r�Aкk9�,[��+n��4�L�\�]h�	Mٔ��Z��f�k��6�w「8��Ca����8W�xv��:Q�*i�p�o,�a�u�Ds�d�.��GՀVuD���Y(|�ʩk�E/s:� 4�Rs/m��Y�&,���I���d�G���QW'��;)|�J^�����1J������:p��҉8$\�/)u������G���@e�B�������y��ȼ����+�ΰ�ͳNh`J���;d��R��P{n�I��6S����ޝOQz��E3������w$��m��⦈ȁϺ���/�4SԮ�o&F����f�^�&;�f��s
�b,v�S���"�LX�hO� .�F�d���t����N@'�����3g����s�O�w��5g<J5���Qj�z�és����0B���e�yi��V�B�9��y�w5F�n���3V�`���jy�ycfG����W.h�|r�Bv,�s9�j�r-j��r�L�;fv	�"L8�R�*��������`���2X�-+��
M8�Qb�%4%�$�͘�0`�k�a���s{�0�;�cTHN>��q\"
G �ķ';;ù8ʻ������sCׯ!d|���;��x�����7����0Ζ��k�6��-ݽ��n�f�Grn,Z��+��aob8��w(m��>
]�`z��X�c�yD 6Y�y�kxp7{��oL#/X����ˏ口��Z9�3�P�['��
赙���;�Ё�[�'6h�b�H�N�@��F�׳��a����Ǿ�s�0tv��j�X��ǝ�xa�5���#"������9dO��.������,��wr��p��EQМ�ͣȓ�q	��]�/7�Ę�_7�Vt�׏砽�8��@ŧl�H-�h����_w,5��0��w�,�Ox�!�ż�ޙ-Ū��$m��V�[ӓ\�$��O.=���:c��ѯ�K�Tf�R�V�� ������zUNj�&'�OUn�чul�;I=#�/��wX9�@U�x𻹯M�q�
��ʞ���s�,J�[�~�
^sX�pcs�Q <i⹮/Ov�1e��ieۋo>�,W�E��+f��S����_s�-�F:��xm[UE����O^O/E֫W�.weŽ��[�Y��v�����Q<�b�B�$v��za�]�ea��4@f��B��4�v�c�Y;���w���FS%+d�~ŋy����q-�[˳5֣k6
��nm  �Y���{�Z��g,5gkt�Gp��ިnȫ�*%�����w��d�ǘS!�3�-Y��z�f� ��� Ivy�Ș'���KZ�D�ĻFu�V�.q:������5`9,�3M�>PNѹ2,�_t�&���Q��ѣ�a�2d�I1s����3fC��`�[��QV	���xV�{9]ޅm�	y-�-��iˉ�W�Z�&'n2��Ws�XQi{uҋ�(�O�3pgNE�7I�z Y'rPOM�s��qŴ�rYi3���ѷLR���*�����O�y1�5���Y�$!�����`�@u�o��:Qy9��Y���o;�N�=��^p-�d1:���,mj��ŧF��������%y��sA2��kՔ�V�h��#N6���YI��9�G0�לp\�Ȫj5Y�J;Cy�G6�yM���¤ΌU�FLr�uZ���)�;�a���Ds'E�.�)��ݩe�7:�����w��vs��K�c�;t>�0]��/�	ug}��y��{Q�ؙ|�a��Y[`��jvhSO$��N�M֕�\��nM��xM�[f�9�sX�*ո����z0���b�1,�.]����yb�^�{d����v��c 3������L�;u2��^[�L8@�s:�CX��9i�I�yr3D�跎�@E^��쪬��ߑ��'�m�5vq�D���5��
�;�l��%!�G�r����?n0�3k�}y�.�������t@G�{|>>1��;4v|t���
%   �@ ҈� �-"҈��4)@(�ЈR��*+H%*% СB"��P�B�R��- P��%"�(�@�SB�P
�"(?���>^>��ݜ�����{E�� 
(&=$o�{�Qݿy�O:�V'�H���I�������{w�<�����(��m�����x>Oq5�.O/C�=�a�}�39H��H5��*���p��������w�r����ُ8��"���l��SÍ�^�S���5���6����p#4��VUf���9ܹ���V�uM��.��f�R�#g�����8|7C�/�G]`��^��r�9ؗNgQ�ܶ����e��M�]Bu��k�<uz=�;�\�g�s�{+ȃ�xI�}����Ξ���q�'/���r���m��^C�8a�Np����<7wu���������&jo�z7�Y���B���� �ٽ���B�#�
3ޠ�ۀ9�_,xU*n����r,��f���>�&U<S�".���=��eqW@�_x{�|�]K���8|m���V2��\U�M��ӗܲwk��*vO_�}�x����L�%b��g�J����}=�Lw�h��N��Ǭ�<�=缵v]{��,���1^Xy�$�@����^�t�k��j���M�M<�ƍ@�>�mXte�_�z濷y�q���Obz���$�=��æ;g����^��&U�l�ݺL�����슥�������]����]}��u�{���GK���Qjn�n�o�i�=����8x���n8;�#�$��p2|�sU���";'9��Ϸ
��.��e����vዴ�Ϭ�d�1�!����;�G�{�c��(�`�˭S6�Y
Ûˋ8,�sD��%�H���)����v��Ճ7ô��착n	*~�u4O����p���$�@_rYa�D $<y^M�/��ي�=o�����t~����4y㼅�=��<3F����Z�"Hc/����_����{�������H~kӻ�����]�D�,��������~1�L}1��hE���|�j�Giu���Өus�d:�.G<Eng��8�~�-Gg`�N����S����O���Ƿ~��VE�{��콴�m��p��Lۛ�1L�3��w�ԏ����Kv�)�(0������7�����=�!��Y8�B����ۆȤ��\��޴!#׎���ڳ��B�z!�z��{��>�4�w��j�Km���e�~+ݱj�a`9�N��q)~�R34�����{�ӣ�l�/I��[q��4��'�c4h��LIݎmd�;@�\��s�:h��y��|d�G�6����y�	�����A�]și�{8�{x�:O�H�3	�s������{���!x7~Z=��͍��[��iY�,���沇�u
��q��=��v��k�xʳ��ó�E��c���Ft7�V b{��8&j�G|)n�*���o�8�''�G�NVf���o���N�p���ֹb�Fѻ��U�y���Ʒ�e�~��P����O�/۱�0F��.��Ӫ��J�o���x��Z�r��򓚹������A��~8�񝛫�_��8Zⷯ�xb��Ir���t�s�(wv����*ȏx�j�f4�2�o�F���#��_����"yg{�l~��r}�|v�<�?v��b�}uvbgF\S��&�U�~�N���+���O��������/4��fiX��b'c���܊��Q���+5��z�������~�7�dI">&M]��Ŝ�,mq�,dc�p{���<�j�w��n}�����|���h]�����ɖ��o\��ڻ���С���/j����f`^���N2nJ&��:sN��x<��̾���ܻ�0���t_ë�۵�0L��Z�}Ь�P��$���wo�.:��Ϸf���a����v{��٫}�����~���^2�V�&^�H�#��֍}{s���0n(B�N	� !�~o�'��4�E��^+y���1��pT�ǐ���,Z7����7bU��Co�瓉��,۽��=�<t�ׂY�f�I�/��5��B^�۸b��<�ϲ`eၡ�/���L��"�t$�~��õ\z�� ���'ӗ��S痭��i~������X���?����d�u}��Y�>y��5m8<�¦j��M b�p�fr,�^�FY��@�Ub)�/�}}>�������v��7�a_D�-ٞ���0�����޻��ft�L	�@f	�@,�F���K���,�s�|\0g��<Iy�e�&G��1'��m���,�8AϦy�=*��6#㘷J~��63\��wXYV�&�_{sY�:����+�}}��u��\�n2>y��Ig��E1���Ι;@���qo����6��\i�:��շ��T�k��ʃ���	,GYI�s��	x��y��b�m��қq��������n�K�W�i�Ë���5��Mo 's�<����n[�cX]�X��Yh�m1�$�0K
���N{g�8����׳�^�G��WW[���:�<�R�����v���c��;���Nd��z)�э�i���nn�(k����]��s�\$ݍ&Ő�$��4�\���p��m���yٗ��l�;No㵼�غ����'�N�+�<�G0���[�Z�La�n�=�cH�<�^�Q��/J�q!9^ub���Zݳ!�]%���"N�u���7g6.��ۅ��[��ug^WR-�jz�pC�n#%������J�4��%�-�67]�=�c�Mc�W�ź�\�</�J�ډw)�+J���b�i�]GZ��\���v����`4�<60b��b�\�Pf8ɇ��c=�4s�#ݱ-��j�GTq[�2�.`�UӃ�v��;]u�ֈ77/�׏z�7Y�[;G=���y�'^zS6 ���ݏ�6�-rH��)��&۵0�f�I�n�C��lG�*Գc1i��e�+�ܳ�p&��8�'k������WFvC/=m�:��i�� ��k<�r�]�7p��B4�lc��sȘқ�ر5�.�aK��+�c]B��>%����Ԅsb�Uǋ���ڴ�l�e����1�u;wGc��jM�Zc�;�����4j��{�qv���m�8%i88����R��Ѩ#�r궻n�E��; 1D�e���B�خ�Fс�3���m	���h�[ u%t���Q	�4��f#8�����xۀ���S�����8L�эi2P)6������33	cm�.��9��8;�3;�����uM�U����}���n����t�gI�蕞��v�-C��mڊ��M]����87Ou���%��]x2�v�+P�֜"����$�"��2���\D� �,e,W[D2k�l"�p�Nd�cݶl/��p���6�nz{z�)�@�MLvH���C�nV���o��t��ih�Gu���^�u�O*k�Nc��B$�N5��j�af�@��Y��I�Wj�f��P����y�·kVB5b�9���΍Q�d:V�7(�-��YJ�ܺ_\�]Gy��V8E��`�;���3�!u��N��u4k-������S�|�Yv�������A	���Xk�%Ĉ�Gnx�9�.uƏ;�f�yJq�%v�iƓ�EZ�N��Y����t�O���bD�N���.5�q��Ɨn\���>ێv����Ƹn��<�Q\Ӷ�Q��ׄ盶�^WV�ġ�kH��N�k���1�pv�趱Ԙ۲#N��N�N݈���i���z<*Y��tpBg3F6hYb��mC8%��'�����B����=yu���q��Ix��C��y�<ܒ�J���ډ��Ưf'��:�m9�<�t��s�g��z�nT.[�ԝt^^�Y�k��ղƻ%�B�fMY���~�o����*,Ϊ�]z�u������������������������������b�ny�v��UUUUUUUUUUF��᪪������j��U���]fZ���������������טu�8�7tNf�sT8�69��l�,����u�[�ŵ�:`�T�`Z�����n3|�|����Gw~g�!3$��Z�A�jJB�����NѵEV&�F:����u.*�̆7¦ iv���6�Ir`�@�2`�$x��x8��+I�����H�v�m���!GQ��a"CiN8��WZ(�U꠬ԟ�s_t���]ܻ�v�o��t �c�[`xź�8��
lUF�O�)Z�(:n{=J�v�s<i���Y"��R<򫅨5�}�(�]r����EKXSUϱ�[=�'�4��]gŃ�y��.�n+�u�3\�]�x����N��޺�z��.���L̴����+k�45���]�y���2�������f͎��lzݏf+�՟i�C�ў9��V�����&H �����[��:8�Dp���n���2grџ=�R��!t=����[c^|1��x��%�N�L��2c%�̝�*��ݸz�j����ن����U����n��*���q'x� Ԉ��	K
RU4 E^*�U�B5A�%-�T@�J�%F4D�4"*��m�>�F1\��zy22Nk��N���~�	��g�o�,^$�U�bi,ɧ�Ӷ8BAHS�e$U���U;��l�AfDګeM;���Pj�!	nm��B�ͽ��Ͼ����>�l�F��pf(�lY�[��9���$P�+���t�K�D�U�0
	�s����8�xu�T$���̷ϧb�$����v��|���j\�%ByAm��������R7ݷi���k�ɸ�0O M�j(8��~{�1�.p�䷽�P���vcmv��*L$V*��E=u�W9(����*���3�o7��6:�
�rV�d��5�kr��ZH%� d�^6�9��ӡP��q�&�<I(�R�!T��ȪY���"����B�$��ƕf���������mG�S����hh�	��V�N��µ���{�����Q�`�W1�_)[˚XPA/)�'6��.�)��GXo�ѸB͈)�em��s�Cc��w��P�d1(��f+ǛǰG(�A��BH���׭o��Fn��1B�W}��ܾ�C1��jw������A�aH˝��k/�k����Sv�̳[�o�}g�-����ᑙDm4l
�WP��YK��\q.Y{��d�7�92����^�n�L^ˎ�\��]�fv�m��������1d��L D(JRǣ�=uoZذl�0���U�/�9�e�RDҘ��s���!t�ڸY�W��z�@W��BQå����s�!�<�d7s���٬��K���nGo;�Iy����M�p���q�r��m�c:;j�v��3����OwJ�����UI:6���z�Il�SB�V��o��0UJI!�C.���;�B�%��ݐ�xW+��j�����)�7]�5�&���),���h֭���}�ɼ�LXA)o(�mc�� 3��le��H]I����su:�ę}w��.]O�:���iB	����{Ǵ}�(�L�$M61,E��L'���&���G;(n���q"�UQ�յ�ۧ۪�E-�[W��Y��H�{Te�[�W��z�z�:�&��0�Î�l�zYH�U؊	R� ���76�HoO�&d�b������IR�׬j����^I6�T="o*�Z�!�D�!	$r�<�2�u�e�Wq��k1(�M��z8�E#.�;veV���=�¯f�ذ������ObZM��cH��]lLd����t����k�=�pM�# ��Ci���n���ٍ��=�7s�}V>���^�⫊!���UVh����B� ����ڻ'N�����ͧc1	Y[F�鷖���&dD��pMfwj�䒬�xsB��;���<��a%7��u}�����%���{{듿�ʘ&ی`���b��ގ��oZ��Λ�+p�d�l&ΜL�""�H����w��k7V]�i�Ss2MB�7���x#�J��V�T�+n���Κ��I4�	uK2����0�>u�;�r�a¡3�L��yH�Z�;����H��(�ŝy�vNr�5Q�$���C��G�?}=��_��FH�|�sik����r�Ơ9���i>���x'm���M���
3`��ۛX#�v��ȕ�8�nx��a��}�z�Ӧ��̀�����!��z�)>������^V��L����B�þ�9n�av��x�!��Z�s�XO��o{R�/�������{�˴ѐ0�9n�^���9N�/���$�!�'���V�\3�=Q���dԠ��L
q�z�KYѰ�3%WYP�l��5
�*�k���N/���'|���e(��t@fQ���z��q�3)�!��I�\�8��jP����m#�(fW�Ԇ���0�&*6��14�U(o�Q�'hLAE	AA�qTBv&���:玻ϭ�3��Z�~��V�g������&�TH�	ڧ]��������=��u�_���6�fu�b��3�q/!�O;�������G�
�.����3��oc��N�z,$WР(���{�]������FZ�ok�o�UW�X)���l�=Q���=wٛ�q���N��ѿ��ē?o�ɷ������Nl��O_���v�D�0��\+�:��R���^[�,ZF�&j�v�������URIl���W���ߛ�!��!-<�c�.�6�d� �������.�Ҽ�ܚ��;p �� �
3�N�|�ߡ7�%<s�*[���\Mgt��N/\$j(��f���5��۵k�b��1�5ہ�<��~���OČՇ�U窪��E�~~�]�Y;�9�>P�*Q�9T����j��������ݯ[O/���])�T(��f����N��HL��ҋ�����ʇ(�� �/~to����lg">ϡ�3( V5�D.%\'�^�����>y��	!�8��)��g쐾Y�GdT%�1*�`�Q<D������w|�}����_N��핂I��Y�DG�T���]��<��=舩B�,ݭϟ��בwQ �!	T�K��b#�����i�#"I@̄<T#)n�!�}oZ����y�35{.��v!��x5b�$dF,�#~xUfM9���딷2��������������>�*�e�~]���Q	';�V�v�M���ET��D��)eu�-�dv��������%X�D�"�EUZ�M�$�"B�<������<�oA܀f@3 y jA�w�{�2&Ё̀j@��sל��!y �g]������ly���9��Z[#���8�pm�`�5dME}�"=D{��@9�$2�iR�k��1�������Āw%h�@�c@o�jϮO��\�d��f631a�Yr^g >J4�@���μ�h<�5�m���̋�5�2.�}�,�m#��o u޼뾻�w"RH;�&H`�<�����i(�F���B�4Ʊ���m�߯:@�A�� �5"�H�5 ��e�2� f �v��<�� 8�ĉ���7@1 �`�EԀj5���͐u k���λ�B�=H�Ș�Ԇ	P�^k�3ͷwo����&8�h��a���ċ}̲��8��v�����Ͼ%TP^q�|a�f9�q�˻�����Й�I�2l��Qc ����td�:趫����ג�<�!�]v溷]UUU�����w���B9���8֍f�LY�s���"�8�Hd���9@�A߽��;� �D̏�u �$+� ㍻<��i�<�u��uמt���o#�"^`:��[���Ps���&�R.`ԁ�����ߟ< �H��܀j3 �|ߌqͰ��D��̋�5 `�[s�y��P�����>n f@6�8�5��"jD��8�&2���z�~|�ΐ5 ��`:�Hd��s�c3��\-2U�y{�-���q�v�\��6�:�A܉��i�Z���:�A�D�	�S��E��iς�� ]^ޝE�����l�W:����0���#܋�:�7��w�~r���q H���mc(���hH��"bR�u r`�]k�=uǞx��;$^$pH��H�25���m�H��R�םu� ����T�͌y���f�s��U
[�o�K�C���I�Y-�"�$I���j�Z>[[_g6����o�$��D�O<�z/�@�"D��	氁�*K���	i�b��W>fB�(�̉��Gߣވ�y��޺���PS.��S�?��U��At($P������g��Y�'�|�l ʹ"eڷ�����b>\��뮲&�l�!!��2��zw5�\`nUK�	-nݺ}�޴��(��N���R�#7�/�醪�g{�w��7�m��� J�*�Ǟ�g9�k��~����&�����)A�F`�(�)L��	'�V���Vgu���Ҷ��J����0p�M�۹ȑ�	*�"l��[��P<�
�>��|��R �Q�:�-���E}�O5[ ��O���� ��	3��)�9*ܫL���;���iOg<�xP�<U����_TN���oE͚�y8}���o@ޝ�
<���^g��@{}��xm�����M]���z�zU�W:���,���{u�� ;�l6q�Zpz�7x���)�y��;�Xy��V���d�u
��Y��t���ӑ7�9��r���N�2]�����B�-����ܗ�q�=�H�[:{�1�\|�����Rk�N��ٶ����?ԏu�G��@��m��4�&�zɀ(.=d����c�T��N`���W�^J#��J)l�#r!�0�LU�UUAE�& �1؆�����������iJ�(hh�ZB�hy��K,B�K�(�����)B��i����y�1	A@�!ABP;�CHU-RPā�DEϣ����c:1�͜�&+p>bc���v�U����y�{��<vTr���ӑw�]b�m1�q��"��%a��Y��.���!W$\·<K=	��i��鮮;kՎn�r��ϓ"����Vz�3nlY�ְZiy�F{t�v�k!s��ڤ+�n���ʪ9�H�m#�;���,��6O�]���inE�]���ͬ�����.�W���w�����u;���:��x̀ܧ��H�q����8��V궺��p͍���s��g�WK��)�(��6Z١-(�)m,ci|�1'<uݰ�8��n��mVf�o[���jf���z�UUUUE�5UUUUST�Ui ,����W^q�?�ĜN$�-�庰��#�I�Ӹ��d���T�rc5�$�S�yS��]��[lxnJT��/]X7-Ջ��KsUUVd�������W��2fD(L!B�J�c?���=����Êz�*�Ejd�ڝ��5��樊	Rj���r+�+����<��g�̻Տpb�y����x�F�	���ƻQ�t�Tu4W*s�S��z�k]n���Q�9�Ϲ�da[TsVƵu���}sc����ڮv��J��������v��i�@0$D���Y[��w�e��U��s�=���{܆�F��cө�w�˱�S�m��JCҀ&RG��L"
�o�*�׺�����*�z^e���zN��q�P���1x���]TI�3Gxޓ��c&��r�ݎ�s��z#�G�����5��I)f����׻�P��7nf�	I$�Lۭ�W���u-�H��H��H�)(�[[O�1\�( ��▻w��ґ	��X�I��k��A�1o2'�Ns�)�c��
�۾��/L<�W�as3�Ȉ\��P6�@כ��g9�z�K���\��:�8�;���|sl�f��Z2�[����|y{I�t����*�Bq��YYO_0�5����NSGfkr<Is�,��^>]���ۚ������{�?[(B��;}�� �	�}$pW��������jz6Q���%@��ވ��z!c��d�*Z�KagOg��W��\DIv�dI�a�.Ԙ�Y5�C�y�`��M끮����W3UU\4}�~��a�F�K]\�f�Wn�!�}���g.0�Q*���NJ7�|��ʺy�n܄����9��3dUT�{���!������.����<�y"E�Q�{�#t6�ղ��k�W��k�+sF�I%ܳ!���.�=g*X<�˛j)����@[��ހ"#�����ǿ-\��隊%�vu�g+�y
�b��������c7h�J�·;5�~�����m<�͕�U\+),ZPB�e��#�H�Ґ��{��sW������!�X�3.��v}�}s7��G�v}��fN�h���Tj�ވ�z�'�	d��%W׽��w���BR��u��K�EF�;f$�F @��bc爂�;ÑSf���m�Hؙ18��y���RVi)*�kR��b\0�V�j�Bͬǽ\�o'����##�A��9
	dԮ6pGP��{ކ=�=�XO�Q�ur��w�����],�|�h�q����V�J�N��+k~�z��<�`�S��V�U���u���O�G	�v������f))����u��ȸ�a"����y��r\#7g��] ��*��f	U�)ֲ���UKT}�r���y!�ZL�j�1��3��t ��J�Զ5ѹ
���r�������1n3s�l��:�����7}��?���HA��%2�P���n"�}oZۛ��)%�o��t��s��n2��O�9�m���b�����s�|ErR!��/�V��{��N)��ƫ q꩓!и��tr�yq�g{�>��z��B3#�/L�O�<��x��,Y�����炊�W�
�5��۞�Ϝ]Q���8�[\�g�����CIL����Z���������������):�o��=��w��������6��� 	*fƓӷ���w��i$!.�lE����=���P���ʵ~��Y��1;^���*އ_m 	�L��d��`�,g��槛\F-{��.��=�}�ikĕ�_"=�7��Y�f�A�Ɍ-��#����;������B��.���K�s�*Y������t��p�͜z���G����_��#zTg3������m��ӕ��ՙN���+���T��%r����ꋯ��+Jsp��U�GF�f��4�/h2�����*���;�������;O���`����b��FM�fiRK�s0݌ɪ)7�am�b?�3�DzG�'P��"����J
J+��8B��&�����B>��E�5B"�������7%*�"S�W.�-�4�`���)h�%sR�k�����-�!��M��#R�C솷���0j3��m��y�H��~�㾵���JjUQ^S}��7rq��H���d��������n�N�Ƴf.�U�֨JH� �Uvk�j������'�W���}��.jW'V(zQAU�-F�ygy"�� J���\�`1Nˉ���s�{����x�
�ݘ���w0���2�J��(
s�~g8sg�L�ݎ6�~�뮻��F�{z�ɋKQ��ٴ�%������׮�Ha�BB�D����U>���#73.)lTɹǭ�r��GT�I�W;����ޗH�	x�����ϴ}��j}��/%����x\�1vd���~'qCM!TU0��R%@�-*����B�
��P�(Ь�޻ǅ�}��ͮ��L1E�u�{G?�<Q�\]�UpI�8�zLd-��p8�/OkM�s�5�]��ͮ�=����GO{���&h�f6�4[q*�і��^sq�k��C1u+7S=���.\J�B(.}*���}=!��Twe�#wu�7�f�i�U;���}��^��kU�o�>���K@`i�DL%)fƈ�Pk���}b����!,y�A�3q��؁k-���N.��P�*UTU���{w)����"�ͭ�`ڄ�;Y:����5���^b�	�W��ӏ7���.F����J��(L&@�%#1)%3c���v�p��U�R*8�2��˽��n��&�W�a"�S�YLh��y��h�5\�)���G�j�q�K��v�Q��׎������a#��7���O}G�'�'h��M�i��E�DA%L��]Y׭��[�O�*�UZ��WB��5��P�I�z��v��Xa"��&���6��d���٣8~�,>���4G�x����'(����s�۴t���9�vDHFB�����[\�1��o<�z�﷓�v|ňA"�iU]l��p���R$륅o^�we�Ѫ�T�#rk{\�J(B,�-u�����?E�h�z�g�����4/�NȪ��p"/ޯ#̿��~�xW�vZ�T�Ca�0���7\p��.��<y�g\k�^aٮ�n�9'[\f�y�9(�F���m�WO��{�Ѕ���W^4�(��%Y[�]i��P�I�-�Pj�w'o���Q�1:q`X�I*���W0�H�Q#Іe_=��VCj�$�*���"��u�֜g$����JB�T�	�dL�	JG6�
�k[�6�&��C3��r}�[lR�ƠU�
�H�ڎ	��"g��O�߫�q�Wܐ�A�wK
��.��V�Z�����|�>���&FMWٻ�{�+v��;p�J�+�B�/=y;_~��>=��>$z�H�oKӣGc�o��@�2bD$��ѵ�3}�G�dN����2EV��~�z�g{����L�0�_nw���z)M�Y;��������z������q�tæU��NV7����|n��1B[<�ً������u��S����nM^c�-�!��켵�6�=����b+!���WM�~�"�~mpxN����z�舎L��V�D9t��o}����;?0���,�X%��#��:��w1�j��3h$�^Ws���q-J�f������)2q�9y}��Ugg�<h��o��f��3��s1s�edU�	1^��-�S��E�8:	�vq�X��"Ϸ����ֲ<>4\%2}�Q���q�=.��1C鼷���Ö҅\��p���[�⏱L�P��Q��^�c�wcq�׸-Y� �.k�=.C睜�y%i���<�=xi��n�|�:���wQ Fx�)�ɦ��m��_f�ټ/�c�s>�ա�1go���INO��,'
��Ms�_u
	�?s|��iNf����:�E����y��<��˷����х���8e�������..>�0&�������!�k2Q�E�׮�	�u*��JՓ����C���*޵���6�
7��3R��JJ��솮^�-۵c�
�"dwk�u��{�7ɷ��Lj^Yo�`��&����ų	������ӵ v��:9����b��D�mnԍ�7	�ۆ�:u�ݛ�7��
��$�E�-��J�d���ۮ6�qոb�n��N�@�VŨQk4-b@��Lm��wE/c���7E���p��[S��8m@ipM`&��:�8�;��n�qm�ZԆ�mɹ�)䄔�YZ0�P�h��4�P,��F1���.T ����b�޵q���m�<E��&5�QN�����|��<e�������Ӟ�%n8�q�H���\�2]u��r�8n�%�$�bA�aԯ7Z�'j(�5�N��v뤻UUUUU�F�����j���6�cS��h�A��7w��|]�/P Ų6V�X�"�!���Y1��K�Y��Y��-�w�8��x�2<m�7n�ڈ:�9�Fy骪�3w����}G@��l�)I1( ���A�5��þDm��V7��8�D̡"��f�w�-�2+��V�i�:NI@�(-��l��"���m��&�J�SH�LQ��T�D�s���T
t��f&$C&�n|��m}�b��b������_��P*V�m��$��x�wc<s��.��|�ApQ8A��5z��bk�ݸ�)Zxp�$L$�)J[b�A����ӥ�Ş2iUl�}����5I��s5.�KGE��ڵ���3a�u�*?Gj���RȂ h�Wwݟ2��@�MLc5�e��O�n|�$�+�%�[\�->�JR�����]��N�}�yĒcD�j�����y��kp����"	ݡ3D�w5}�k؅���Ԑrp{�u�AdOF]

�G���Inc�l��U�۶�Ȱ6Lm2���ٽ��qH�}W�f3:�M�)�"�TzAN7�<��9�d��
"���o��X�$�3��l]�-o��*���y8n*����xA] v���<�-����e��7lڱ��	���fE$�\a8�h��:�mh��3X�c��=sB[[v�e�:Ni��=5U��;��O��5�٬�M���~K�os�Z܃���=�{�������AsO�v�=C� ����} �޼��k[�J!|K�NfWcm�Þ����9�kv���rq�mr�R�/x��̩#Ǣ�����\H�<eȲhΜ�Qzs�N�3S��_G�����׿|zA �A�������`�I]5u�gfӼ�Mi&6j�f���,==^{�G�%m���i�l���M�ۯy��,ABu�Ս����:n�Т�dK4�=m��YJ�T"딥Pn���Ƒ`��!r���~��zO��'�wo>�>�O�;[�-���&@�z���QAlZ6$�n._'�t ����l��
L��#QT���m3wۣ3	5=��뭚pA�R$��{̼��:Ae��L��\,k2lV�9;Y�5�?{��Dϧ�Oݏ�=������@��e�+Ƌ�κ<���{���'D��!�by�>��ٮ�WИ�ͭ��~A��H�p�e�i�xȘ �qA�
��;Y�C�3PVS�����i���r��m[,����,�����:~��c4v�:��7"񵶽v���Y���y�Z�0��{uU��s�n�n���GL�/=5UU����}}}}Cp�K=���
E�}�<`D}y����&���%	��4#�S��bl���Q�"0�a�{��b �c�! @�e���1�s��c��.��i�ڶ�A�F�s}p6�_s����WS����'^'~�����u`c;Mf	*f������bw��H1"�c��fj�ï������"x�+&{l��h��訡��!���?�!�0��5m[E�p��o۟{[�o����+�A�jд�eƢ�p�n��~���f}��1-�j�����g����t[^���=<>O���X�L�i�Gc��k�[GSicD��~��/�o��F1,{�z�uO�B6mng:C�D1 w�z�H��!�<#��H���F�>���������;�۲���yz�=�r�1Z�W���7�"�[ذ���Y��	���r6��:܇r��wk9��Л�n��۾�S:�TWe��򐧵_���\!�m�/l�'�ޛ����Ld]��a���_q90�e��_j;ru�U��]3��Ty�;�Ov�@������юb/aG�G ��n?D�8��`������kE��d.�m���<pZ���r>yN��Ǿ��e�#4k��yN�ð�y}G�2umF��謣���j09�	�=x��ΗՑ��/0����Ȝ̼K[�!ƭ-���W"�,9��s#˷0l���eTH��hP�9yu2�ADU�5R�i�3r�=z3.
H�h,T�K���|�����^`?+rbR�eX�i�m��m-�J�"⭱�����q�7�=�׭�iՂ=K��mk\�I���"55�o�Zu�A;kuzǐ� y!CY�}Qf9����o�}*ڴ������=�.���l����dfe�����ڴ�}��~����m�O"5i� ��7Zt�3�k}��5�:ս�t�-�im��y�{�����O$m�	r��!h�|Q���o��(8j���S3|.u��{y��}߲�M}���4~6�PK�snvs��-���:�np���،�Np~o��(��	b��\���6�Zk���j�����m�W*Dv��`��u=���A�b"�׬z���m��9y�۾����k�]B5l0 S��(E�y���s�=�)(j��%ZF�y�i5�����z��E�#ЄPYu�ls���*���Dخ���Y����]U�h�n41Yc2���@����t��9Qa�+�=����\��/�VZL�+V^zj�m�����}H�j����.�BR�h�|#� =���1,�=bZA���;�f�ޚE�L�o�ｫk���Nk!ı�ڴ�9�����]k�W�m������:���i� 繕��w*����㬥9��o��-� ��m���޹�/�Z助�R%2�����j��>Q�Sj��X���<���#���H�d�}Ry_h誁��6�Y���-{��5=�}pm�1�3m�3��pg�̜Y��s�z��]�͘����]�yw�F����ް����,�Z�Vաi�U�7����q:�-�.��9��ɶQ��.6�iA۾%�y�	x���w�e�|ԿO����ƭ-�D!KQ"G����|ף��7T�ǣ��j�CYϺ���d��39�3�7W�|�r=�0�# ��Ӛ�"G�G�
�f1g�s����`�l������s�z����!n1R�6�j���=��j:�x�z1�Uұ\�&J��8���ȫylkH��U��S{���N�9'ɂ-i�i-�e�_h��Mg����{-�+�u��+{���i�H�<�mz0y��<����d�P��5���H��2:h�4i�{N����{��`c�r��3�o��[�#��sb3x�e�u�>k�:�Wp��m��w�хԸ6��be��f^�k��ؖ�Ͻ�}���K��^B�n��%�q�3��}��z�E��os�85\j�Q���{Z���G��C�C��H�`Bnq��j8{G�9�uX�t��#o^��m~���x[\N�!�G76"
�������8��fL�qb
�]*��D�up(�0!S���/�];���r^1;a�w!]Ʈ&�ـ*�%؞݋��\v���Bc]�fv�m�����*4�u�ma�����%�^��a�_{\���k�Շ�1.Am	�]����o5���tq��@����� 6�[Q��2}�s��i׭U���=�{��Z�u�O����}���)�~��-�Qj��j�%��w�}Ͻ(�_zUK��}��}���SMqq]�Ձw.^}�q���,�}�}�#w߯_5[j!���7�u�^������sm{��e򏽫��V�ﾙ�#e�j$D�����+�l�U{�}�ϼQ���UE�!� ս��G�F�-}q��M�[j��N�Ͻ�c^��~![��^����+)��)�"R%2��`B�!�!l�>��p���p�ʶ�OrV:Af����-�'P[N��{G;�X��4Z}�]U��s���s�Z��e�]4*A�Ǻ��^7;s�<�ֵ>A�b͂�k�o��cR�3��y�J8՟i��նǐ��\ŏ[����h�#�y������Sk��6ŤGq���ܝҖu��gy�s��c^�}��McU�e��5���������{Љ�[���[���r��[/vw����N�H�mZVL���$`��V>s#��7����6���H�X��y�=]��`r�<�o�o�=b � �=���1ta�^}2�D�#E��7߳��ۄ���\%�0.*�[�S�F؈ׯ�߽��Y�u�'Ȣ�R�E�����j�i��s~�%y ����V��X�E�����3����!��;]LEXH�e����-��R߻��6�%X��"���u����c�y^e�Μ��vv����v�ퟋ#���J�S��=@7a$=���zz��<����=�w}�r���хi��9�g?����85��Fy?���M�}�<�!�^�~]H꓁k����g@��gnwWMO��q!@&75wvf��fFg�L8��6�w��o�hrd��ޅ�M���a�'�}wq�o��<�bT�����S��l_���us���\=�ޗ7s��T��_�9�o��wI�;��wC�_,�l�>F��9V�g��nq�b�Tv\�82\����dH�"ݖ���'%��_n�Pgж���m"cG.
u�*��r(ҍu���R
� B�PJACO���P��qb�&���2q8����J�EEy˼�ZT]�-*���q'!w]21K�K���q�klU�J�޷P&彄�]cc�VY4f���sC)*P�7=L��4Tؐ9��×�� s�#ø:8ܧ<���%Cvvyz4,K#��fau�&��� ��VkR܉K	���؃6�w$�R@+ը���f<[��n*qp���w2ݶ�!q{��T8��[�q��ocm��86������gG[�mZ�1vW��;�y�9��kj�E��,;K]�n��<�M�{Z��_����my��m#f�!1��s,�؍�#hW�l�B;U���5����\�D�5ƍa�r�Q�[7X9�.�UUUU�5UUUU5MUQ�����Cz�M��������T�����Ϟ��SJq�4�ۍpD��K���cȝQ�k��9C�%|s��������>٬Ey骪��o������r;����e�̽��-�M_����ҏ�����������a6m�"ׯ��xZu�Tms,S\jж��~=��>�������EJ��&�H.1�9��}�z5�'=��z"-m�j�[n��9���}�;x�h�"\>��޺�{�E2�Z�����d����Q;���}�^5�����U�H�dnK'Q�w�g++.�s�s�\�t�Y���:��#����<�q=�����	Mʶ��<[�s�s�5��5ۄAcmD-�Hk�����x��j�c>�b �B=�(�ޛ�"rs�]kǥU�c�z����rɆ-�̷%ݒ8b���~h�8ն���_s����$�>5h[V����E��N������E<�����1֒�jڱ�D�lv�U��?oB_ND?gz|T���TtPw���~�����<�k��o��1_^{��]%qwg�4�rjؖ���s��NRHC����jG�D|��ۜq.���aE��Q����	���y;�q���E(����4|����u�`�N_��p�[j�k���ڴ�Zl���{wn�u�#�y @�!�"G�A�d��m�b ��y�7j��Z��:R�Mɕȷ��2a��>���8�"�8sTq�Ɠ������ߗb)�6a������Sj��͢�k/3a�18�Zg���߿��ʑ�DKH6�<��mop�w]���Y�\jz_�陶���UmF�Dwʓ{������}��#E�hZk>��cMT�k��5�z�ɻ��cV!mZ�o�k�#7*�PǰA���ewi�o�O(��w&��������x��O�4�+��-�Q�i���ڹ���p�W��q�tz#���!�o0ͬ[CG\u��v�랪#�����C�����[��
��c�a	vi,���F�"�s9Ͻ�i�N��櫍D�E���Y���'��y�}���B6��%�)���F�g��{�w��ѷ���j�ݜ��c��^o�}�I׈8H�#�!�";/���Lwnuo5#����E;oW�O���dHإ�xx�Z�e���Ԉ�lKM{\�����X��� �������O����D�@m������Xa̒�����#�������F�pk)����MI��9����|�)歫B�7;�fڭ�n�:��C=M騱 zǐ�y�̓��;7"�h�� �!�����Q�%�R���;��Ր�4���s��c��=���[h����m݋�����ϵ߽g�xאu�X�6�!� Fb�|Wt���]��f!x�[�n��嫎��#_|�{"�� � C�D!��w��{�;y�����p�������|����ih�m��V�3yϽ�:5�#�F�I����l��Y0��K�ʱ.���׷���J�-���p�^y�>B5�%����s>�8��뙿��ƾE�:}���࢛�+"�mZ{�s\3�w�ﲏ5�'�b{�{�d�z�A�}�w��Az���8�(j��D�����TI�]����x5�Ng0bs���Z�?�y<մ7|���X1�,Sc3j��o�K-�6w��{��`n�4>5��V�j�s�ޫmZ4�����ki֋T��lKB5i�o7�}�w����c^}��B1���B*��szǳ;o����>CЄ!�Ì}���8�0��1�JC�}�C�}���Ȏ����.{P����=N�=�31�0�v�)�hZ;f<�d���1{vp�4"獹�]��pF�D�/m\]��m���nˢ.j��n{���0�k�,��=��j�,�\����~O�	汫B�� "�V��o^｣Ȼk�w<!t�V�--#mK��~����j��Nw'sn��#B\&�ϵϾ�c�")�9��cE��m�o9>M�3��k�Ep� !v�#qZ�&&�#f\���$ �[ �6���=�R��y� @�=d-:�r��8E^�A3Q��P[ݳ�MvyŎ��::�u�yێ��Z��;�فKjдFڴ�g9w�{�����#E�j�KH�Dg3��xk���g7�ު57��lKC�v���r{�Ͻ��^8���0����ˡc����cy�����؍�k����{A��~�^���5R�90�Zj�f����N�H�o�}�og�-�.z1�N���(��nR���ѺYY�>D3q�&&:ʈJ����$t�V���劖c����1�ތ��3
p�u������|�bCC�����I�;��16�=�����y�V�wpɹ�3��/a������G}�n�{�<�o��͢Fę�Z78{9�m7̀�a��r�i@��'r����xQ�A{ޅ�I������!lw.N��x�~�wv�}P�ebk��{���u��z��8:���w������C�?$:ft�#$��8i� ��w���yL�o$��l[ؚ58��*��E+� ԕ[b-W�)KM��8+X\�3o�%6�0DDhD�rV�(��
�fL�ł^%�o	����8F�j��q0q	�{k2RP��8�n��j}DG��3�3�mF"'S�����s�{GȺk��{U[Km�)i~����
.�[��]��#E���4j�|��Q#b�L���B��wx룊�������ٍsk��J�V��6�=͙��&ӻ�3����k�>�}���բ�ʶ�סy����IרF��B�l2="�<�m[��s#�ZP�Y�E��H¨T��e��q_{޸ٌ=�! ��:jv�\!�����D�=���6�;�?]�s���F��R�@�a�=�{�"��,���#Fڶ�4�3*�>��޻�^5_'�uS��R�"��=y�J�Ӯ�r:jzUB�[cY���Aď""�����tz�7�_ٽ�jڨ�KL�^���� c�yQA�w���HL�%~��j�f�{���e�t9S�z��>�f��X����ȵ�6����-C��t�Q��1��pMG]7)4�+���V�+�K\�UU�g���}}t���,��D\�>�J�#Vէ��{�L���DZnU�hve�5cSYϽ���[g%�adB5m[US����/���w٧�P}*�,KM�LH�Xզ�����`y�P�Ym	���A-�]���\�o�}�]�Ԉ�[R����ݹ�:fe�q� �%�u;8ᱛ���>�٧��w`��D�6�=����C����Ae�彪�\Nr��jO�>�FD�8a�t����H�p"㶅 j�֚�j�#y3z���}+�-�p�g��ͰM�����׻�f���>'���QKH�Ul�>����L潞��ۉ����6c����f�J���-�#	ylt�"<�m]"���߸m��N:�VH�b)��\[��]��O���g���>Aܒ�oBCwr���x�O_uQ����?y�e��՛��/� �|��<1noM���׬D A�*jfJ��ۖ��+ʑ�nN����-M�����K���|�@2�i��A�Hj���X�#Ȓ�.���ϻ���&���(��y�[�G���aL�3z��C��m�T,��җ��_{�?Nl�������px�*c�y�֢H�+,ШAr��Vs����qȚ.�"*EJꋓ7��y�y3�vu�aO���c�(�}����yX��$�%+�v��� ��ɍ��9��`;_�zK�s��V����N峿�;���M-v6��7MR��9�PY�7�*j-�n}�ջ��]�hۍ�謧E��C���^�:�����Q����﫪I퇤�\��L	S;�������F	�bex!י��t3Vs�ه�J�1ٯs_&	S0�0ܽݝ�ؙ�$A{0<9����sO��q�<�R�10T�Q&T���%3`a����&�Z�Q$�J����"b��6��^޵�vB
퉚�ݒc�y:�=?6�pҷO�D�j2gE������I�)� ��=�ߗnȞ��"I��ݪ�i����P1|d� HR>F`�T��+;37�o ���}"%Vk{̸tf�z���nX椬��1FU�f�Y���X>������.0���|�=�0DW���]�1��D�"�$��T�-�6�3{�U���b�3m������)g�z�ǰ�"F�MEnռ�i�'R0��&�Ց~�-���!����z;r���B����}�zg�؟�S��!T�� �&��GS&���^�_kϾi�;|�x�P͒�8�ZA�;�7�{����E��t�.�T��� �ɑ���um�Y�y��2H���nz��mg�Ǒ$�X�B����������Oz�]ܹ?T���v����
�K`��n�;�޻�'o�=�[�U�,�]7=��ޛ���I�V�����C<�ۦd�{��aǭk\󸎞�E�g�L��Ԝ���W�d	c���;�(C��g��:�:x�' q �n�vּeݲ��:�uz�J1��p����a��,� ˞6��=�q�}�yd&�>�����WP�iߴ�壻�:3�,-0�pu������Lc�K�b���Z�f����:�J���3�R|��97y5��&{�\fh#Z����7��Ͳq��O��n��s���Q�H����v]i�j����G��5��3-�hs��M%Nj]������7j��TKj5h�҄M�]��h����S2P�m�)ěC�hmX�(�N,ΰ��x��<I��N��O�~�7l
����6�U6�M�I�w/M�QWl(p6��ؤ���:� XS����;�����MAWKyf�@��\Rk6�P�mq�ٱ����d|qr�#��4�q3h�˛�;e�j]�l`^��*]�E�m�/�[�k�3Br\[�]�p���㧝W��'���p=캬[�n:�0�npv�g��L��jK4�[z{Y�\[�㇬vػ�����Q�8]����i�H`�͖0���:0���+�����x'�%��c>��c���.�;�eօ�9��X��]�s�;s�.���"��jz�mzA��͵�^z�⪪���i�UUUUUUUTM�P5���v֭�����>�V���2�
��Y&�� c��]y
m!��-ic�ӷv͊�C�U�g�;&��\n��
�j����ߟ��@�\���B�����,K������Q�v�B��=��y�$��!9K�Y���u�9=}�H�mD>Cr��z4΁:vaU��0�Y���is�}N�w��>{˘���` AV��60ץ�R'�oX�̩@���R�z#_�o/�k�0d(
�E�<�3׍�L�7�|�{3�ٷʻ:$D�$�MV�{Ym�m�d�޹�sq�\j�.\Gb5v�� ��}��-"5ĲIK��m�h�5;��ZU)�Q�ݡ�?%:ҵ��nȮ�������{���Ϲ?���j�'1��m�R�K0���i�l�
�y�ۤ��O9�6h�M�V���1�GM���\˞��Q�Lp�M�����y�z��xmb�5o�f�ĝ�>�<F�=��#;�ޱGb� ���q��䙩�͎�Z��*�[�{�tO�s+s�o����!��S��*'Ҕ Q�j��$e��H��7�}��}���H�`�8�EWU�si�lτ� _6�l��A��_f��B1���xŮܽ�j���Ju���x��@��d����I(��((������%BL�RD�)���.;s�%�^���ogE����p.�g�n��nlp�Ոuyn��)�Gd��i�2�m��j��{���+Hn$���
	
2��Бw��y�E���,&)�Y7{ܷ�#�l�&Ϭ$ap1uv6�2K�7wr�^_=n�D�R��aYH�:t��1��U�k|�,G"��yӷ���>TN
k��� ��%)ofk���Td�*΅"�Nq���hA�hbYw+e�5�DG�.tp��k��h��vd8�������[|�%�Fu�$]+������ڈy���:"�x�o7�8��N�u@��M�T3,�Vc�o:/U�o���^�U��,$�[��Y�(>��|�tC
��wnU#�%М�-�Ut��3�6Ѭ��uj�{3�z9�}�s�>H���P��]�M�=
�r��`BJV�(�
�sj�5t��$�2�R$��2a�p_�,�z�0=")3!u�'�j�ytP�y!�.D�{qc�mS-("��>W���r�����>�G�y�jNÛ�g���;;��
��W��H���Sf���=�RTW\Ӯ��sv҂�h��z�uuٽ����CtA��W�q�9q-M���ѩL�sy�w��1.f[�Z(m]vw5޷�or��(D%{��{s_K��G��x�>!(�WR���S�Hlû�vq75�u\�]�*+L-�������(�F��<*���k�S玄Wo]��kŮ�Y��
�r��qg�.ɘ:� ��n���ٻ�����M��$�K�-&����=��]�����Cڨ���E?���W���X��ŭ�Eِ�YG��ǭ�KKБ#�AE�/{˳ ����(b�k_Y6o���մ<�����n{uR�Y.	�	�H����ZӘ�U�� �"���;*�(R%���˜��j�̕��~�_C�u{�S��W�H��g�:<'s^>��4���:=�0�������`��$�$oǖI��77���!GMO�_&G�J�(�����a)K/p���_>r8���H��DR�חo��SU1 L�AU��{Ok��,�+L ��jN6=�xd�=��r�탽��Y�\�������oipd����FG����=�����s��䗪I�{���y̒���Ք�������]磴�{}��ħ5�cTu>G�؆�;wB%�.�����x��=�������_b����d{h��np%'�ϙ!�F�+���=
�P��xW���9m��W%�
��ӊwGo�����}�s�;/F$����]��5��20��vϻ{|���m��,(�)f�u�y�b~�y��h)����(8�6���"GhCBfM���C��)M�D߼�s�14�8�ؠ4�ih�D*�9%�.AM�Q��cT\����q��V\Z�LJRlKŝ��
Z*�
F��pfx}�s�|��[w��9���C2��{���N|.�A��o1�m��}w�}v��T3,Ȍ�.��f����]�(�(%}T�:�7��Xamć�9�JH��^W����I�*��Z��֫t�4��3D�&k�Tc���SJK�������t�4}�ۺ����� �ǅs���3cs�,�w��q�IU#��z�klr[đ!�<ɠs#�Kyκ00�]*FTH�!f�m���|��A*ؘ�v_n�.���E��B�k����*��h9�}@�&TLW]�v�˗dq��JV�s�Vy�{q *�7D �B�b�m<ݝltl^,��)�=禪��f��~���k�Yu%��Nnw�>NF��s[�De�!T��.�X�cn��S�-��s1!(aev�o/��Id�&n�u��H��*Ss�O7�N)���uXS��R|�� ��B 1 A �F�ЂY9z���fW�R�uz��T���4�%�0ި�z�%�}q����7�tF�+�$�G�Q�����e�������ܶ�f�TR!�g�Jf�����].�⪏g�H!1D��� (��5�ҭݫ|ӊ���P"�I��Q1X�5�����B��N+�}b.gk4TN�0�#&�Tv�}�w.�0x�ʏ���}�[��HfLT��1�ke�%s�	]�oe^o�E;�}�窖!�6��7E�{��{����"��胈�@�뚻���l�U���$���sצ�4P��T	�V�w�~����o{����w	m���o��߇r�
vE����gK�[�z����0�m�9JT�BR�!�S �S;pE"����#��Z𓽻�>��j���0nE�	)�p��0��;��H�9�q6aoOwo
���ZV!�W:vu��������|�(��%�Ҟ.7`���u3�
p��}��/��~G!b�mRz}/�<��g��[����w.�ݧ\Gd��y퇠�cP���s�<��G4�g������~���ɜ��
�F��"��^��O'5�e=���i$lh�U<����D��$�NI��Ӳ�$V�yAnη���J��C&(!B��oX������M��"^6��1<J#�S3�κ�LLKI"���#�l��V���Wݘ�#���v�Ǽͳ�YFQC��<�˗�+x ������������f1�M�?��������C�c�O��(E	H�� �T���+';���\�`h�����d�����Q�]����rϽH{����J����b�r���}U��Z����K�*J�oX�p|Ča�*���;o�������!�q�ill�Mk+m]���U�������³���6G]�9˻3Eo-��n�AO�`�e�uZ�*�
*M��8�[VD,�r܉�Qx&��o+В!)�|m��6>KD�ַ�u��	{~�S�ƗUٮ�4�����0 ����[]���H���j�E����mv5LTuڋ��Z��Ecw�W4!9N��k1S��ȼQ��v`Σ�u�<��:߬g?���A��?�*>��UIO�AA3`���PPO�����
	�k	�2D��`�d0ɾ\�F��j��=Ə�C��#�:�:�v@0m� 1J��s�:3�':wݍ�&��H{,q	�l	��L�=���/v6M��0��>aPPOĆ�� z��ǝ������>!��<��0De�v6�D~�`Ό&��?��0`8�2�ѓ���������0�!�i�q����A?�'���3�}��?�,/ H"('���
���B%&'�>��Z����}���p~�?M���!���S�?�������>�ت
	�U?<\��"�6S!�~D�EM���Q�� ���׼;�K�?y�c0�?�&1���X6��O���$��z��vC�n��5���c
���������g6�߷[��~G�үAmT!��&p�`�C��3��B|�������j���˸;�T�>&��!�o��5�q��d�bo��p�;�?|��M�{�6 �P�����?���S��������3�PM����fP��槱�����|��\������#�S�'���_����C�ka�.���|����=�>����!����y�
��{���`��?o�0A����NC`�2D 0x}|��q�5� �	d?R�('���	�� ~�`O��5����B���rl�=��?17=���	�n�1$�\����GٮA0��av �>'���k���WhI�qb����{�	�w����a����4r�+����pPN܇�>��?�O�O�T�_�����
��~�p������=�B1���=�� ����}�������������O�?!�)�S_���9Mw���O����|/�_�L`���~�')~�PPL/�o��˓���C���������p���Oa>�Î��p9 �r��~x4LA�s}��� 6�`�������S�����~?��)��vom}��(&~��O�M�_$����{c��bNH��������O�Lz0q�&�i�o�A?�_�����?��@��~o������|A>K��h��A�7O����lۆ�ی��C��;���'�#����z�����]��BC>�4