BZh91AY&SY�Ɏw�߀`qc����� ����bI��           ��m����h5ckY��ֳ2�Y5X�`ɶh5@��M6�[U��j��H&�k[[J��Zͪ���(Yk*�Ң�F�Rֶ�f�����f�ն�Qji[b��&M��l�	�IH�T��V�P�!�-�M��E!�f�����6��I���ed1��ճ
@�@��J��[R�炪M���m�����xR�^SX��b�]�WD��Z!ZҶ��"�j�F��ZՔZ��5�֭�ٔ��06��[�%j�fhWc);&�h@�  -k�y���Y��{/m����-��^�5��D5N�i��]�+^��5Wz��{qۻM^��[i��wj�����n�]%�V�וw�;験Rڢ�c)#FmV���P4  �
P
�,w�ER;�x-�$�����jQQU�W��m�b���}�*�E^��$R�j�s��
G�ER�{n�H��km��o�|D�R����UZh��d�l+UZ�j�X��@  �M��R�ھ۾��>PT����b��Wl�J�w�f���ks�pSM��9�>�J��R��W��}�j��}��J}Z�m[>���=���/'�|�}o�w���g^���Ֆ�X���R��P  w9�ѶյN��
U��^�Ko��G���Я�4Я}z}�t�[o��|�ꔦ����|���T}�}����!Jz}�������}=�Qv�[kN�;����lͳA�đ6�1���� ;/�T���}����}އ�E����}�}���x��>�hP���|}��@:���>�Ҩ(>�s瞠m��U�ݯ{Ҁ�=��@��8�(�J�s���+Z[d`�Z����o�  �>�ւ�����)Egz��}S�C����V�JR�>���z ����F���={u� ��.;ۼ(���㸧T�B��y"�4���mh����5I�֐��ك�  ��נw����=��ѭ*��u��{ҝz� z��.� R���[h�{��w���:/t��zm���q�
�����S�23m,4��Vl�  ��{ ��x�4�}�@�^��������zC���q��������z���=;�m��B���6���QkE(��6��J ˾:CF�^y@hj�{n� �u��݀=�f{���;��t+�������x�z�<��zձ����(��X��UH¢�e����� ���:�:u1�
��k^ �ֽw�=� :�(N�]P�֌� =ox�� �Ύ���`E�     ) 	
R�*T�      ��a%*U      )���H    4  �~%**�@ɀ �4j��4����=S�S�44h�6��A	I�B�Ɉ�L&�@ ������%��"?(y��ʣ,O�*�sun�j|����y��@W�<������?�E U����� U�Y���������'�������O�� X?۪����?�	?C�'�Q~�����zFal.fa3+�\���.ds��2f0���ds���2���̎e��S2��̦ds)1�\��29�̎ds#�I��L��S29�̎as#�̄�f0��̎es
fG0�`s�L��G29�̦ds�3!09���L��09�̦f`3���S09�̎e3��2���`s�L��S2���`�L�f29�3��fS0�as fG29�̤����9�f09��as�&09��.es#�\��W0�as#�C0&dʙ�&��W0��̎es#���2�.es�2��3#�\��W2��̎ds�\�� ̮as���C0L�ds#�\��29��d�\��G2���as����G0��3#�\�f	��ds�\��29��̎`s#�\��29��3e�\��29��.ds#�\��\��29�̎as#�&G0���`s#���29��Las�\��̮`s	���fW29��.as)���0̮e3#�L��G0��̎a�s���09�̮`s1���G29��.`s#��f�L��09��as�L���2��3(f0��a�3#��� �.`s#�2L&d��̎ds�L��fC0���.`s���G29���as�\�f29��`���G29��ds#���L�09��as�\��2����ds fT̎`s)��f309��e3)���0���f`s��fS09��.e3����2��̎`s)�L��a̦`s˙L�f2��̎d���G2���`s#�0�Bds#�\��0��3+����G0��̎`s f0����.es f ̎`��P�0e�3+�29�̦fas#�\��@�.es�2as�\�L�̮as+�0`��@�2��̎es�\��29�#29�̎ds���g29��̎ds#�\��0as#�\��̎es�&0��̮as+�29��L�2d���!��́�C2�e\��"�dE̪9�2
�D2���,� f\��Qs(.a̪9�W0��\ȣ��3".`̀�� ̠e���W2��T\ʬ¦e̨��W2��@\�+�Qs*�e3
!�s&f`3��� �.ds)���10es(f09�̎ds�I���G2���.ds���G0�`��3*f̮as�I���W29��.as+��� ̮`s3+�\��0���.as fa3#�\��0����?؀�����j-R�����!��6}e	)�@�,����u\���¢SU�� dbv�,��)miR��V��a�Żr`M�+wf�iЬ����H-�ON��`nރ���An,@ӺS!��&h�`��[��l�P�ܥ[��,�"��	����-V�ٔ�!��d��0ٷV�KZ*�@H�B�Yd���&�l�b�.��Va���+d�V)�������t��e�8��0ʕ�[0��R���e�Ҝ�J�b�
'@�X0
jdTm5�+D��(F���2VP���m��fD@e�f�P8!̬q=�{kM�҅��զ�� �ݭx�V�)�+�%c13+��3uh��L��=�r��MHPyN��Oʻ�VAM�/n��d�V�5:76N��a١e�MUj�f9�����l�,�Nͥ׆���ч1����6�V�\(b�&�p��5���M����:ZƦ��l��VM���*yrY[���y%��9�tcNI-꥗�޽�*\ؤy%�{+/rh��L˚��	,*U����b���B^m,i������+t^��v�X�{�vaw�OE�נKS�n�;T^�B�!*Tw�r̭�.�c(��Z�����\�b�oXߒ�Ȓ�,cKc�JQ�R\��楕mf�a����]�ZYP�t��1Ǝ_��2�mأ��"kj�L����i�yz角L�jS�����Z���Vlb����L��k;AU����Z��:�e�x� e��i$}�	���[e-L�d��ʫA�7#���酫�&;�ɠRvVV0�U�L��^
�:��ݺ
���r�ס��V��7��[@�4��3U%!�L9u.�D^#�-�jM
)�t1 "G3T����FD 6J�s(U֋�N�te!D�����S2���L+D� [f	]��Ģq�!nx$+��L���Uq�am� ��f%u�O���r0�21�d8�&ѭ9gF�v�K[��uml�l0ո-<�X�	�YP\�AȤ��ԙJ�uj���F��[�EZ�~PҼ1`{nT�ɳn;��
�GB?��@ѭ`<b��l4��/V
�f�n�e	��5�/-���)��TiD/V�VҧR^�5]����f\��ӊ�8c�C#��f��B4��	daZ�̪7KT�k%,��b�8 �_H��Dr�)@�j�܏v�[fh�s.�BjZf%Z���S�=�e}й��.W�3E��� {m<8�1y�+K�ŵnÊ����[ �2�E�t��m��P�ڽ%�v�A�NQj�!w.k�n��7m┒I�&6�B���0F�T��M���1�thܷ-�����T��	W�i2Y6íU��E�[dI�7������ P���H�k��Xʘ��t���R-�$��\0����A%���1<�����M��&�
��<{�]7+Yچ��hf�Yj@m��U��L�߲a�eѱX�|�HҦ2!�4f�y�����x�dP6�2��`�]*iv�h:ܡ�L��݂ ҁ��u[�-��j�E��JF�kv*��o!�rբ�h|����b�>��u���ED��H�z���ٽ���^Pa�e�&�h���K�
��Y�	X�L�:��ԆS�p$v\>�n��;�D�ʍ�ڀCuF��R	h�R�WǤ���6�a�6p�F[��M&V'���u$�ʙNQ�v��XpC��,�"��YSt|�:�Asa'kn`iT��a0�L���Zr�(-̊���E��\�!\���K8�k2VS�*�*��
+p+Z�@	���F`o�]fZ'�鮜X����@�;��fّ��1�i��7��2���(�g�[���7M��A�eI*�6�z(�״)nY���n5��jʊ�n%V�p�mTMM$�3U@��FV
�W�[E��&��z
�TV���#.\H&��e��a�.�PҌ[e��5z�I�#�.i�y`�W�*� i�+`yB��]��lV;�:�&�	�L8@/&]a��D�Y"�P�0YV����b�Z�R���7�E^�jʇ�{o�f��������q�f�-kx)h����nMk6T�%]f�`�X�wsHY�c�`ἑ �m�ܛm� �,�I�p s2�Gx.�b�������+fЫ�=�(�yV�+fY�f?�n]�t2o�)�b�ըmfM2K'$B��A��i���YW�JRڗz�E�ۊ��a�ߥ�9̛N	�˩J
fm���d�1���}�[�CY�*1�a5�Ͱ��Q���v��v�������7l� kHH4���X���rU�TT��,E��P����ټ���t�y�U��ɚˤ+���]�g7iJ�7�9�7)���PJS����LK�a���+>e#�pڎ�x���1���ZfUEtkC�ec,c�.�J�J-��⬴�`��.d�����o��oP8�P��Bn$�2��/\LG�T�$��������;dP7�wMm�ppcT!wx�y��jB�gۘ��\j�*$]s�ƱUȰ�eb���3.\1,�v�) 9cb�1������i���)#W R0Vl�]ZӚ�j:��3L�%
�[K\8"�LPp1�/,Y�Vb{�j�'���aMR�'i�mɮ-�,ڒ���Z�sޭ�̷+5T�(�gsI�AH��VE��c������5�8`M:<��WP	�i��ٺA���Vģ���t�j�+*��(�����ɍ��Z�2��k��B���C6C�����{�i<�"n#XP��U�;�!�܊�ly���[ԴP�Q�jB�x7vZyY
R�ʨtkyZb�bK� z��(�X�M,��N�ȴ�i�H�G��2Fԫr��d�sYݔk~��%m�jL�v����1Y��X�A�k��m@N�R�R�)D'¯2�ؼ$�oq�g.�h`t�$��Vk����se�
ɡ���kS؍�,9��#$�x�m�on������΂�ݣ���j�
` �a�FidB�
&��zsW2Z�ksV�$��am�R�D�N0�,�l���)�
�g
ʘ�1��"�0P������y6����kk2X�A�klR�)�[-��&�w.� 5�x)9�HKR�-��J��4�nIl�R;�e�M��dܐb�m�bLV��W���mJ����Ƞ�ջ��2	�ź�D(�+"ϜX�b�y�gs�m-x�Xn�T��cdt��5��Y2i�w�^<�IV�6�V���c��J9i��kX��6,3����ڷ[&��V��6D�(\ȳ�ur�˭+K!J3���C�cc{M�K;,�_a���	���lX��R�.1l��7Yd��ׂ]�Or�=�JeB^Ǩ�ZNL�Ќ�D(ܘ雚D#D6�WI�u����̊��i��&-c'�/���;2�sF�M��Ah�ױ�13je��pԄR6�+v$C*V�R�`���e7 ͱ(����ku�~�&,Ukuk�$Q8�a,��)Pr�mh���<(�
9�J;Re����5G#�Z�A�W�@*�7�.0�̎�tY�IJٶ��Bj�:�""2�t��q���J*Ȁ�Ku*��xvl�hP��r���ͬ7l9rn֓�a���Ζ)4�j��u(r�e�zڀ��/a�Ԗ�U�j������o\;z#	(Tڏ4�2��v�bI�'�|��!�WX3`1f�RO�.�ںT���ޛ��Aj�^FLW�m��J�☳H��n�ʹb�l�־ˠ�r
���6�7�iK��rg���P^�����Pm�Z�� ���rR44�g*���{̠%9cMX�V)���K7E�#P[�m�ڳ���f�̅ȕ�4rī�զ�Y� ���][�FMB��{��ڼ'&�R�ƪeӭ�F�
M������"sr�Z�-U$��
(�C�WX%d�/j%���j��W�B"��c��O.c�Ӗ+6��"���
�]]�.�l�vtʊ�A2M՘��'Su!�f�a:Re�
�dUa�l�y��%V��Rʺ%X�p�К����̆aݍ]m��hÆ�&���N��QɌ$qP�e��g�^�q#2�B]#�#�
�!� ���d슮��%�i��a���~���E�]�yѓ4����f;$-�jW��Ȟܚ�կ.̵��)K5nT�Ҏ8][m-4����KKh�Z�C{H��4]L���x����`]�d���cf�ӄ�9Zړ[�����]�&TM��` |��R�b�R$í��wb�F��Ѭ4��t�Z�:���Dj����<�h��ui�-�*'a��)7馕k��IBv�b��gr�T��4%�4V^��bȕ),M�N;4U�L�ws5�I����^��ȫ/%n����ԁ�L)�j�5S���e\�&V
�u���#\�;�l*J�N6j3n���,�+.-�䫼�	[OdW���A�K*n�F�
coJ-!�.R�����ʺ�!'DV�5Ϯ����
��5�5x�"��95mdD�PX��u��VQG-���Do�{qt�tb՗.K��K������f�zj���Ǥ��M�RXV��1ּ���m�)]����:Q�n�,͘d��zX����@Rl0F�+v=�U���oPå���M��T+ne� ژȻd���L�y�7Sb����x,��8�*&葢L;�
5i����Q��	��˨�ސ��`�bM��֋@Iv��6������Nń�Rh^�J��u4�AwS��fTP�3@ǩ��N)�nPVPV]CP}Y�R*��*�3ɟL�xA��Ht�nU��u�{O r�^��L�z��Qb�� �h�]\��3@�
̉�Ғ�Y�l�SՏF�Da�@K
�r0h"�Kx1g�jV����6fi[1Sz�y[Fm��ǉ�ա�y�b�¹�Ԣ!�w%��r�
�K H=w�h��3d;��]��8IӪ���	(�,p�Y*8� �ld=˽�]�Xa6�yR^�_1��A��YX�V�
�5*�� �L晰��Y�r�:� ��.��6B�Չ���Gu�2����n���IS��re䩉8vAN��xq8��*�\�����V�yQ4�7U�l8#U*B�a�6�X���l�	�)�+w[��L`�w6�j �Grml.Ҽ�L�4iF9��R���<oHE�V��6���01����d%)�xj;�Wr&+r}+0*��Q ��*%�����Gt����܆܀�V�v�=4����Y �Q��X�۳V-�oS�	w�Q�)m�kYL�U%�A�*j٨�0asK��
&�5�rF�h6�ݫd�R�݀m�p�@i^L�)é�)�,Q�&��a�e�i��L�&�K��%�Sm�p�"�ڰ����z�`���qVK��� JI�ZKNA�)mX���a�M��ő�ԝ�%���1.�H�b�g�w&�h�H�-�L *�u��]X9�	N��Y{Y�������2��&�^�o�LR�Bn�e�a�5�v92Ь;b`�W!�/wb�`�2�
bV͗��f�jH��FZ�k÷��],�ZV��i��5�\��d7VnF�t�]����Dk�)B�V�FnU���]G��ܭO��y�Sm����:�i�-^n���"zi��m6N�p�td�5�$��IU��\�����{`(-����
�6m��m�ht��k*Q�T�Ʉ�"�V`mk��q^�m�#/5*�75Fż9>E�T\��1��.�@�V��Vpe�K ��t(^�B1*z�0(E�+0c�HDVY��p��&����6�k�rL������X��Xs\�n���2�U�G7�K�m^�{N�d�4@sl�+b`T����^��{N�=�Ǉ
���\���v���qt�\� 
�+%��:�(�Cn�B��^�3n�1 �R�F�\�˨U�k�t�[�H�p�H^�e���ndLK����,钺�DF�e32���]]����7.m�)���4ڑ�����4��p=AP�O+'wY.���5 ���)6����e3���U��x���K�k)���,F����|�����wv"@�
������Q��d%�%M�6���H������-�Vf�����̼盪�j�b�4�r�5���f3X��r5,��]��s�����h��z�y��-Lk4fA��8SU��C�S!�ҝ\I;H�e:t�j���i�mk%W�|�5��㜛΋]�N�.�#6��m�Ff<��GcB53�Y��G+f}9�@�̼s*�n�
��+<��cC"Nfc�[x'���&����qq;���7 z��Z痂1�S%%Dr�C�|��� L�Mz����XT��������<�ϯ�
sz0H����C,�����|����b#k�
��,2����(��H�c�u�c����+-*z쨀ݍ*�9��<������=�z6J�<Hb�J����q	ʥЀi�+��V��S5�vz��"w��;�}�ݘ��ٍ�A_�%J�3:+�:=�;:����D��v�(VU��.��l������p�Y w����b6�]��e�G����p�#�g0�\PyO7��	�TF��C3��>m���}J�o��{+�"���WWg%+�����	ROb��X2�Xl���M��X�πc�@X�T]]�w��*-S%��F������Ą��u�4ju� LM�͝J�v6��6^���]��VLj�Y���ݴ@���D�Թo�����3�F�r�)�-��N�X�Ѫz�EP��q<4�ʶ*慅�b� �$*b�%C��0���O�^��������;C����?>�?O�~��`���J�ɛ����n���Ѯ#�т9/.%V�OHX	д.��Y�����(�w�eD�ըjW\ޖ�=K;vpɂ�L�*Ҧ�9�r0.&��]B���Fӡ��U�k�����o��8��t�V� 4/��,�4�裵�"����c7-n]�ă\�l�
�Ox0*8.�a�}��왗:-)�`��C�{��#+�u��ٽ�boU�2v��V��,s���v&���0���Oq����,�!���(��d���\�d��bJ�6�J��9����:V����U�ZʸG ��0���V��}�	8���,��uk3@�4;��սz-���.\����)ua�`�;��H�A�+8FY����&��ޅ6�6�9gLz�*���yh<\�e֗A���e�zVT壷�n�!��j KoٜM�d�V�C(kw��f�h�֒#��gɽ�x�;#!�_V#�w"(b턺�B��M!�~�}Y[M+�f9,R����w n�ܬ�}�fP�g:�Q�:�-�Ja�J�pi�����2^j�!��r����}Ƒ�����dM����Ȉ�%� d�̟X��Gl5*�HM#�;����ع���b&ެ�z��w|�G���ݕ��"��,e(-:�A��x��+QmG��Y�n�]wn�y�e`�K��3qT�P(\�*[�q]�|u�d`*��C0`���H�Մ]�y4�'�q)v�kl$����b��{�\�������P�����"]W�C�:8��nvm�����:U�	�]AL���M&�t�C���mmv�7��Ғ�6OJ�/sz�]QY���g�P��!|W+AnY���Ek������֧�m�m��\�{M��=��j}���ȳ.��;��'�e���\��7(����]��]��tV�k�7( �ԝ��wXF�ꖵ�ʃ�W���F��w\[��gr�Q�E��EmC37���h��c�H��{�U�O�jd>4+����0I��w��PgVD���a9@m�*��T�7�ڡ�x>�Tܧ#1Qq񉠞���Nl���k-Tʱ��!Ic�t�θ�dw��?�D�k�j�Gjf�#��s.�X�0U��4i���}�����oc�!ā$�-Z�u��3gX�}!��Ǹ��b���cȌ�%�zɵ>p�ǎj]{�:�d�;�a��s{�%G�/�uT̺�le�<�ȁ![`���҆1#�l�4��n�u������}{7�m\ך6@wl��g�c"�GA�NuB9�f��\
��x�>�tzl�`|U��E���n�rM	M_gp�=K	޵\��;P�C�T7Q�m�؊�����]��^߀��=�ի���V�k;�ɾ��2��w�$���HĻ&��@C}ƍ��Q�I
�����MFZ9kwx�roM��O0\��h�g-X�rV%j���������F����q��$n�V�U��^�Y�����a҆bŨ`Aх6tM|WR�<b}�Ƕ���"����c��e�g�BGN��y�q�JV�}W��X�Y"q�T��rR<%`�${gU��U�6�C�Cw.�~�2��.ޢ^�4���]�Q�:���ܤ�6�(�u|OP��qĝM��K�aRĶ�A�k�jd�% �pZ���j�g��p�v0�+���r]Kj�Qrw���
��S��v=K��c��2�18^(�1L�r:P|gk�Ƕ�.ީ�6]Noy�� !);m�>�ObB=* e�H�=u{����
��*�!�2���_M"�ŕ��F3�]c[6��<���ܫ���eE]0X�T�p�,�d�B�22�R1O`[���5���6H�W�^<���]᳅��N�56�mC�-�Ϟ�@ܑ�M�����Ar��}:X����+|� ��K20��MV�MS�v���x�Sq"6�l��W�J��5v&�%u�N��d�BdH�Jߺ0� ��F�7��s�C�b��k@Q���+��s] qe%[w��k�L8�B�3u���G�%a����Γm����LXX²�Ơ]{��ѡ�8!����i�,w/�!a��&(��R�@rqs�tYֳ�E���:���*Sw���b���])�u:U����e- ����s�5|@vJ�gS=M'+̝wP�B�ش�A��4td̜�	�~��ʜ�l]��%_!���m��Ԝm�{�4s�[�����ҷI���u���3 ��e�fT��-��z�K�OkNVa��$�,t���*�lx�o:�]�2�2-�+�Pm��;�1C����ҥ�9c�.��a���6��Ɖ�����uW!��yIe�m��e�ܴ�'ϲM6�<�gqo"�X8#�θ�O��w�	7��睔����&d�������],�O%
��\k��i�E<��l�P����'�gE�u�Oz�VF�[�sf�m��V3������Z��>�f5��8�{\$3=sΒ�X	���~��c��M�DP��4F�FU��b�UX�_Ϥ=p�ԾƳEC��\Evq����T����Ԧҹj�L</�B�Ÿ����)Ջ��Ù����(��'�:�I�%°�}/���\]�1��� qڼv,:B�D��Ǖ�3hI��ǀQ��9%���^pBnY2�vw`p0��v��8���N��Ԗ��}�XwJf��QM7��ǟs�ܻ]��VjX�J��4ƣ������D����1D��wv>X�8a�Ȭ�,��
�S!%�<}�T]�3`�Ͷ�
��Y��r��$�u���
�q*&�Ț����f:G%ǵ�ך�+���wZ���S�DaT(������z*wZ���T뚆��R�����]��>��-�x�gI��ҽf�7�Y�1�h�9�G
�D��e�'G@û��|G^9P����CLtMei���{��43R�;vhu#[�@!H����]t�bI�,^LX����j<71��Mx%�]�4	��%��2�j�uh�y[E͊���|�QH��ʝc�5N{\0T)�ռ6��BA���3�b�lw���ܣ[f�l4Ka����yŀiT��Ǳ�*ww4�!.�/�;1n�y���ͻ��9��$���w��,��j�8�$�{��U�lKٺ��I�(�;���&�tN���Q��3�l_T�F�	�;��\�i�nn�/�-\�5�K�R$=p3��/��5�z�2t������h$�T6s�g;ەc��Jڣ��5�v����/V�W�7Y���P�^����uV�u��R�s��;pY��=�+8�У� �z�w%�(�d��e�U����,T��!�n��%\����7롣�W)�{��i<�����/`|O���� �M�0�����+���Y��W�7O�$�WukL� x�l�]��wu!2�xs��x�j�,�,o&�o��r8�$PδWe����JO2h��-48.�dG��U+�ή�!LV㫫J�B8�f�J�\"�
�f�5xk��'\x�ck1q�K����щ������/_�WՒ��:u��4���:��ҵg�*R!M����\41j箂u�s���'w��g�,.fؠq';IuމF�gv�����wP���^E�!�����*��[��`��\v��jq�S������휟Z��)a�^t�Ҹ��:��]� ���+����f���p6�08�<:6(�8V��;8Lr�J��Ab��}�r��+JN�2����:H��Ĥ�'aη�\�d%Z�j<�a��Cp��m�Ov)p��[��E���j��4��8S.΍r�7$�|Y��+~����6��-�	|d����/�����T�>��ژ��{J}�[���V�.)��Ĭ�e�V��\֭�*r�ľ2=1[;|枏��N5C(�N���q�-�w���fN��я��.�e� b�]���*��C�Z�f� ��S�|����Ne�Y���w6�T�#�EZ�.���Yʾ��KJ�p>�������#C��i�I�[ېZƸV�ϳqX�4�ʘ��Ϥ�OU�3:�u�!wG�r�zj)dLk��;\���-e5��i[�cT
�H�3/�#�:���h�αۙ�*T9:ִ��/n�]鵏x��t�Rs��T9=�gY}k���
�j�j���y��ėu���| �*���xw[�	Ȕ>!.��oN�g8�+��)ʻ[WB@���B^V�^d��1M�c0�K����2PI������L36�ѻ;�֟���K2�bܩx�RC��Һ��3�?3K�h=�nE�4��79�<�e$.d�9��f�}|ܬ��#Υ��o_�X���Yͭ��`��@���"�4+w2�Xu��I���׃J�����A���\�N6���J�}yC�����Y6��,�x`� �g�]x9�
�Wd�p�F�
5{{�osP�)�aA���z^�cY��Hj�&�S|	��_��n����Vo�7MXI��g:��vz����3z�ir���wЇiԵ;r�gZ�6� �l.{��^b���b����<�gP�J	Z%ÍN[�	9U���S��lV5X���n�I��H.�u�y;6�ؐ0��S�f:ǳ�;�?.�Sy��6�
����߻�|����+�E_�K�v5(�:����(<헝�sk.���l�
/9������ޫܞb��T(��"ec�I7��=�+S�$�<�yuӫs�]*
�m`���	M[Yb_[/:o)o��\4��ӝM�8�4�ۛ�m�����k�H,]���S�@n	���,��p�u"=%l�I/�F��
�`j��\�Ng"�J���n�4[Hb��ُ�;X��Fp�.U�m�\U���8Oe.�PL��7���2� �vF.�ee]ЦM�j�G)�[7�jh�5wb�6�ϔ',崱S��4o�V�u�-��*0�'����SV��뛊�}	��qI؝
��E��];�����:�b+Y�s8�wm�1�p��.68}{�qC-�K��!�Rm���@JN���B(O�o�Q��W��cY]WQos��+�\:��o��Rϐ ��S^*}C*�*��Ū���^��3!�Umwt�����}n�)"dpp��|`}+.:=tS����H�n�l�%�N(%�O��"�N�X%c����O�5���Yz�/�[��"M�(hs�9�����
�|��PS+`��9���O:���뫖�N�:�&��H��ˡ�ͣЂ�u`�z I�šX���MN�gI%:μ�X�S�2/�%H�� ��z����t�>Іͣ����U�*."��=;➍�L�}Q�M����B��s��/��S{B�f�9 $�kz�R[����"�@ܳ��%r��w}}�1H)I�yH���y׍tQuF��tx�X�&S�xQ�ϩuЄ��c�]%�����ʞ�D�G�� �ةdd]p����gVk_(h�G����n�|�d� f�u�B]���w�<�ۻSNԸe����[T��*��0k�"��T�F<	�Z���}�S17u{��z�����i��q�z����;w ���&�"&�λ���P�m(B��u�в��vn3#�QFv��/�����G�ć�e.h��� �V$��>׍�!�z�/	qwz�3t{X�<H}];b�br*A�s]t�=x]'� �>B�v���
9���e�����Gk�]�˭jw�7KZ�۴@}\�!q�8��gP�V4���B�SbC�\�Q�� ��c*d�����������A٢�#�}�,��0����a��N~Y�\ǵz��ynt�&,DX�'&:U�LAw{�P55���"�C���J'�\����:�gWS�-��c�]�uj�ݣw�>N��H+L1S�֒�tA������s�o��Զu=��7�N"��	-�¯o�}ۜ�T�*�n�b�qm� (]�2wVfour���$���'wwwwwJt�$��������)'���u��Ή�8����'pk�*G.!IH1������Զ��U�b9�u���M�1�S�s�v:�֝Die��ꆵ��+[iI��
,m
wW N����|�D��2H���y�p�n}B�n�,�C/eޅ���C���׮�<l�M7�xph]$�"i)"Ш���j��A��@�Y����P�v�2�# ��0S�H���7Q�i�4+UO]�ץ=pPu��%0�M�tf�CT��s��D%��t>�!!�R�W,F��t�th*9�y1�D� d�_5�m�E$#���n�A�:�:���Xi��E�M�ID�X�7`a�?)fS�.;�R\7u ��*X�N��Z�bB�S�B�RdP��5��O�*t,�&�DN��-
0j�Qt�`���i�EIJ�Ѐ�R��KZ���	
�"�0�2�
�C����iݰü0J��B�"�
��D��/�$ ,6.�N�E�M  3�H����V�-Q���O��	I�E.��Z&:4id0�T�t�th/.� ��)����3 ��4�Al�N�"�>!���.�T�D��n�R�B� �T`� �O��Ѣ���e�(P����<j��T1�@��J��B-�qD��&�I3�Q�ʌ�M7�O&sT*��(Ы!���!�M�F 1U�V��HQqM�x0��2�O�e��P�17uYS�a��`$ ��}���o TAC���E���װO����DG���?���y����wڔC���|̕��Rɱkht�+ó	�:����Jj���gUCt��1�19i�pt���C#wv,��]d�'�ap��TfL����ϔ�,�Ҭ�F�!�Q�M^��%�4����}����k#B�j�fbz�2ُ年Slj�+D���l�[�+���K�xFM�"�͢s>o�H�:�eYQv�$L�y�Ln��׸l��X��s�a��iF������ɘ��M�Khޜر(�p�,�t���p����6xˎ�;	��ŋJ��̤C��8�v�݀�肮���bַպ�kr�ϫ�zAW@V�i�[�z�R���+7�E=�VsS�b�雼�_n�1h��&4��]�=͐�<&h�4��sz/���Uer�f���S�����&�E�Mk�әO����d�ƭ¨�S�FL��ݔs���V�^[�c
���BP�8�{�]}WW������}[l�s�6�vL��:�l_P�����fQv�s�O{�Z.�2ˑ�k2Q �*��;s�,�A#5\�.��iC��bk[�(�.֮���T\;�@��i���l��8~c�I�@r�/#�T�/��,8�X�h��>X;E*��u ͛2�
h}�T�@�;����2�.\�3�Ն��	�BlЪ�C{��٫����0.�K����#���|3�ǯǬ���z��ׯףׯ^�z�����z��ׯ^�~=z�^�z��GN�.t�ӧN�4t�ҋ�:t��M�:t�ӥ��:t�ӧNN�:t�ӧN�N�:t�ӦΝ(�ӧN�2t�Ӧ�:t郧N�:d�ӥ:t�ӧM�:t��N�:t鳠�ӧN�:u�?^�ׯ^�z�}�z��ׯ^�z�zt��N�:t�ӧN�2t�ӥΝ:u���ׯ^�z��ׯ_o^�ׯ^�z��à�ӧN�:t�ӥ:t�ӧN�?^�ׯ^�z���z�^=z���ǯ^�z�z���x�=z��ׯ^=z��׭:t��N�:t�ӧN�:t�ӧM:t��N�:t鳧N�t�ӥͽ�:T�X�G����| nh��_R4�i3V\�(�B�W+w\�E2�l�	�m�l֍b]e,#w�ۦ)f���u�n�f���jZ`> �̥��7��6l�����=w��WC;01�g;�n���ݒ�ь}ԛ���ar"�+����O1�Y"�έ�t����l�D�\5�Z+�$\%����J���b�]Bh�e�԰9e_^�ɋ��d�3,T����+���\�.���K�����Uh �EX!uw4��}�1�wJ�(�ݓm� �Y��"��w6��B��]����Z5�"V
�m�9�t�T�f�E{N`h�e�f�V���52!y�&�x�ʽ���x��.}���Z�@�v��뫋�٬җBv(�ͤ5��ݤ�#-����Ma�UU�������z�$�U[�v;�*_p��_e5K/,�R\=�rwQV�#��!����%w+���HI�9���#ĭ������n�e��L����-R���_`^j��P�$Ւ�w��h��34D�!P9�ZkZ���%q��R ��WV�}������L'�2�Ӈ0� ���^�T�-��o���PB��5�ˌ�p5g�β�m�Z����Jr���k���j���5�>���PϘ��nt�Q2�lcMJ��6%�+��-f:���ֹ��ΐpV5�4���R�h�\6�>0d�GN�:t铧N�0t�ӧL:t��'N�(�ӧN�:l�ӥ=z��ׯǯY�ׯ^�z���z��ׯ^�z�z�^�z����ׯ_�z��ׯ��^�z��ׯ�^�z����=z��ǯ^�~�o^�z��ׯ׬��ׯ]:t�ӥ:t�ӧM:t�ӧN�0z��ׯ��^��ׯ^�z�z���z��ׯ_�G�^�z��ׯ׬��ׯ^�:t���N�:t��N�:t��Ν:t�ӧN�:t�Ӧ�:t铧N�:`�ӧN�:t�GN�:t��gAӧN�:t鳧J:t���˗6t�GN�:t�ӧ�׬��ׯ^�z�����z��ׯ^�t�ӧN�:t鳧J:t�ӧN�p⮷j��BZ�_n�;����Eٚ����H;j�`L+M����R��uUS8,d�h�ӯy��+��Wp�ۈ�v�i��ص�뻫pG������g�����`Ǵ]
5��D���Q�Qf_>��k��}�g�}F�"u�Ƴ4V:��Q�׊�Z���:�2��X�wۑm�
���c��}�v���b��1gR�5�P �E��"k���0]�8ML�P�n��*44[}���6��Ԥ�+��bGE��Q_b�N`��P����k��7fu���o�78+;s��t��M*���u޼L;\k�>��}�7O�K�
Em���/��@�.�}Q��I�@u�ʱc�V����Uu�GF�Ls���C�r�g�i���vZ�2j��4Պ޿��J������s
G�<6��c��2��Q|"�o`{��49Ն>�������0Hl֊u*�,���$�
��+���baס�[��#�FZA�D7�<u�[��]�Pѡ[�=��,�9.��R�:ep�S��\Y�[���G A7>�_Uwu�q��ۯ��SB�k��}ul�kd�u�*#�Ns+�+8hT[(��PWZ�ÒM9���e3�)��wZqH����YT-�����ɶ!إ�=��.�-�Z��V�
;=vա��]ek�	-��Uۇ���e�_e:9&���C#I��M���L�2U�JF�@ۛS%B|�Wt�,=�ʫ[sdY8+^p���3&}/��{�j,r�1J��/hȈ�Yop�+%��[�Of��ٱc���-�ww�V�3a��]uܻdW�&������]|kS�gV�� �K��5e`8h-y6�ǎ*x�w+D�u���pD�@�[7��)}��WFv�y� �BR�S��z02�:40]�Gz��1��@�e3Z�yV����4�i巹�v��Z�qH@��e��=+�'�E\7Z�8v�Ֆn��e�#�`P��hvn�t�^Ws�z:�(��Y��D,c2]��{J��ψ�QC���pU�5ۊ̬=�D��h,��M��-VjBU�G�vER��[9u�K�S2��^q��ˉA�(�sU�D�NC��y�=f�3�t��U��qG�r��븋���T�I-<}���z��p�ћ�X�º������ߌ�;�]�S����z$������i�6��6�j�_Q�ܘ��{�t��P�F*�7ǘX�U��+��]l���s&�K���L�;�a���r�����ac�N��Fn�;
n �<1��-�4�Ʒ�Wu�.�w���h�����Ƒ|:���}�(����$MK���L���n���৵z]���5�r�]��\*�\Ҕ�������~�貉a�U��ZU�'$t÷�p� Xqe!%e�-��k�r���Ts �\E}���N>���P��Lt[�z���v�nKU����U���>9y���+v:�u�}�f��]>���x%X��`�q���{���*:�w�h���z'��Q�2�j��hQ�nZ���g����wK�j��
�A^�<�ѪL��duP|V�#�%�	F�3G��[�v�쮖�yD��4(��Zr��J!vn jm���������4:��\���gr���i:�G�tZ�2���,����&n�t�$ �qN83F6�,�����;"����
�Y���ư��������`&�b� �P���lPP��ѧ5:���e�����~$�]6�
{N�F����`� ��3y�	��J
<��72�kz�\������4m�rҌj�B,eD��,��b�5�w'l��er���G�W��2��2�0AS#:$bW>(@;���&�c����� �@��	��ҩ6>
���"��{W^�h̺Xݱ�e#35�!�6��l�]�8[�U�R|lcr�r�m��z:N�puX��C�)N�k����]Z�R���ufN=P����ܦYQ�x��4�^�Uwat�oSB��u=W�Xw�M}L�X`�1`_9Z�+���3(��ShC���w �'��d��*8-Ժ��
30�����'@&�+��\�*�9tkp���i�`�*�"���U�d�D�ι9whx{����;Ij���vѭʥ��a�l�wJ޼|�"�rj��p=�����k,IW�+7�,��	d�/I[h��Au�\�i%�eB���%�hҥ��ӡ��e$o�����$OD��Yl��K�ˮ��������e/��b���-0���I!Ng(7�T|�oM�e���	9(�ѡ��r�KO��Y'mG0Z��wvִs��(�UN� ��t��w3B��u�T�*Ȝ�f-&��t�gV��]р���ō��Υ�{u�dO���'	ڳCޫ��F���*ھ����C9PVu���K��N�Z�0v]:<�"�TM��7�M��wwۅ�����Lv�^��M�H�}axE3��i^�V�	Z�<�q� _ U�ý�h�tنwWܠ
=@R�4�m7Ư^zk/g�iI]C�N���]�Ij�4�+F�X+i�� �E�W{�,]֍w�s��Ь������ƅf�O4^�N��:i���]�˂4�`e�M�b�.�w���]�FWEړzam��9-��&�J�|FVV�r-
����n�:x��$ծ=�@�Cw3���%��L��ۛQ	x���G4����c1wC]oW-sٵַpʧ�W)�	O:���u��i6�e�I��Kig�ʍ@��j�sV>1��$jfp�1(l]��lzC�CZ%��CP�R��=�S疅;���{5�Ŏ��4���0x�fE��o4�PP*�c(d9{R��t5�e�E�LC�:q{8k�2z&�n���c�5X��T�G�+%�{β�.��$�J�X�]&/�f:+j;��;���J�}�J��݂U�e3\FdZ���H�#w�	2�\��+!F��Z�Ol��4����F��b;�)�S�z��WVW	�fSj�]��?^(��M�G�Μ�[�2ΐ��f�8��]�z�qt���C�}�8�+ͭ��U��+|+O	j>HI���K��®bb��{J^;�����"vu��eYP��U�S��O �,�*�>Us]�2�gd�����&�����R�N��4��n��D�b�S}.��Gg'�$�yQ�����b
��j	-9tE4vT�j,���YG�e[�n��=?B�J QԻ���D�>*�=Dq��b׶�e
�B�D:���lQP�mc�ۺ�u�k�����݄\�7hۧN�TD��ԯ�3E�V�����9(�댝��7s�r�蚟L����l�(��T��زs4゜u�רH�ʺ3Nk��釫7l$���Kޥ&N��i�-�Έc[��enZS7]P�)��(}g�X�:bc�;��ʪL�kU�Bw7��IX63�.o�{z�]'G�)fK%��^��k�U�}��B���x�V^P���M���P�G��#��h�WIӡx�V�;��?��+�2�1B�����w/����ó�8�ͱ(剄�-G(������[V�]�ʊ����:���u�n�}��M�s>�*�D�f޻d�m+ok�=��T����Պ�8c���J�[ �2�xms1�U��"\�����P��ٕi�B������c%<��>Χ�e�OoE�%Ԡ9n�Ҋ�0���yҚ��ʵ�pS��7"���@���a���!��s�/0l�떚N�2y�g�퓎�y\��H����aV�-�ۡ�g�fP���F9f���ae<<Q �d4X�0�:`ŷ��UU�1�W[�q�YY@ߐf����"�G+r�#3"3�x�W�V�l5Q�gw8�4�*�,�vЬ�"��yP��@Q	��ZS2'�-ڢ(�5����[�e����M)�p�ڏ�̳����Θ��6��Y�[��}2����ԊҒ4桻�ʴ�2� ��m_,��i"}�ٌ�W�`��i2'��W�hc!T��"'s�z<��Coz�"!C.��f��x`_QV]|wE�����84�����Շ����y]��|0�=*���xm�ч"��gM�޹ yϦ�p�*��汧\�(ٶٽ���3p=�Lwe_eM
��!�h�p)_N;�5՛6��X����A9�d��!�h���v�f=���(-�K)�6 �!���ݫ������x��b��k�د0v�
�X���Ul<T��'b�pU�C{�.��fl�,Wb�eQ.*.�n��B��Z뭂��^%��'d��J9N�排����N�,�Oz�,��%rӫqJZ71�"�'XV�oG��ݨ�c�{Z��m�<�zxG����M��n��a���s͌��:7؞����a ����9S#��w��e�m�2�i:��p�T(Z��:�3i�vD+��L�=}���������s#]WO�T}�Z��4��h�16�fN$2;`�3�a�}��ޣY˅�kl|єsCB�kL��P��[m�3s��K|�}��1+�����8�M;G3�m2���FtKk�t�!�Fݠ��98��6�8_)���o:>���ݣ{SF0`�jT�MM1�_f��e�7:愉����+V�$:v��C	��f���V%r:��qY��ϕ�,�� F�d�n�R=����&|�`-�3oP����aʱ8�5ь=o�rT]�-��(w����4�.eguX,q�"3L ����\��R�;wԄ��wU�|\����ف;���vk���;����TV1t(/�� �e��V)>�}(�����@v��o�_6z�;���2;x�3�Mb�Q���Ǧ��J[�~��ܡ�xvҍAboY�G��i)��A)�g�>-w�+�٘o��X���#Q�	Gj���4 Q���uu*�7jN�i��<�ķ�Du�B%I��-s�����Ĥ�� �u&�A�v�|L�O�]d��E.�UώT��+A�OǤ9R�fI�����n\}>���s8�(� 5�m*�lP��}�V-³�����mp�gpB�ws�[����Q�ݺݘQ�X��zeؾ��D]hU�TdH�� +��,��P���Ś�<�CWc���]�b����׮|5�rĚ b߿��  $����������П�@�>��X}��$_�?��6�1Si��f��BB�.R�[M$�	��aҥ�}"�iP� �
��Ca���Wl�]O�p�����3>��|��q[#����X�d���7�������h�P�*	T�0�/��H��]\���nC�Cм�wR�n��7�gw$��t�2M�kns�V�q�Y��(tk32�pJ��͓��ݤ�bg�75k���ۿƄ>��0V��;0��Sę����fQȨ��7O�9Պ��b�;�|��+���r���������Ɔnco���٘�:�u�~ѻ�����O�c���k1�#}���3���&��&&Px�Q��Q���eM�Awi�F�K�c�E�Lpŏ��i ��j�ᙃ�u�\��5%�CY���DGP���Y���`:���՞ל�1�oT����:��Ҭ��
��+b��5\�{6^��?u�D�^��>�A�y@T��prz�X�%lu���V����.v�䌉�\QO*nn���@>q`�KR�wKM���tW��x�*p�������
���L�j.�h��;����9������o�d�T��Km��^�=UfӴ��g(�-6y7w����nsƠ��]*۝�;Jif"[ټP�T�`>$� !���LP�1@�d2��!�i�o�@���
��)�"�t�|Iq 膤�!��,
N�IQb�,*F��5[n�)��#L��|��uS`� TڧI�$L�bY�q��Fɡ��.|��T�@�����=Gc�16�Y�lձ�F*��s�׌珧���������ׯ^�z�����z���������Ȋb���4TQ�h�Dѣ|P�88�d��������������ׯ^�z�����z����������/{|ڢb��1s��%�ۓ54\٢֢!��7�M��c�ֳ����p��"�cUT0MQ��y�m�8��Xڶ���;�6+lQ��*���:ūj1j�Xv�s�k�8r��p�AEE��D�٫{�ƎV,b)��{�
��5["�rb�j��9s��j#��
Ѧ�'�l�Fh��5l�X���N�cL�Z���gͨ�l�O"���51Z�\��b=m�h��I&ڿ9�s���h�q�1��+�	���&ۜ�ɫ~!��}��F�%H���X���wF��{O�#�1���E���.5�mʼ<���&��[Zo����A�A(*�(��5�m��k<lr>?�Ϥ<��������X�N��A��������]�:]�%�j��]�.�r�N��{_�l�~>E-;��W�]=�]T��;2zU y\��x���Y[S}���{�͢�������ۉ��z�d�zM�{�����9'V�=�~{����ROG}�=e��4�{ϫ�� �v����.�{F�z�H����J�Vs�{ھ�O��/����O9�5�%��;�zsԤ��u쏲7�x�>�g%��q�=�w��z�6x�n'��j�%����^GOgP�v��u�7{� �4#Kǟg%��9��r]�3�a�h��&z\��c�Lz�y滽<o���C}*���;.}��	��⦋��{�y�_��W���|�����u�'t���Ʀ�W���ۘ3�э�Wۛ��/J;��:K<�,\�L���5�z����DQ��r��+fjwoYwPq¥��Nq�s7�Z�Q��=��){�a���9wK��N�l�?tbu���K
�P o�T�J��[vGPy�k��<���Q�7C	�R,����\4�/w�iγ}�ѫ�������!pw6�N�a��o����&c��C���8�F��+�ys�^42�s}8�1�}����M�����w����\�K�̀������z+���հ(W�bu��\LDG��<�Cx���	���wk����pϳ˕�.B=�����|�S�Ϯ��kv�R�	�S�VUw�_<��6�`k���{��G6����4��Uu���n��V�uzs���.�=�J[�&޷ւ/ޞ2WQ�=��^�h]�=Rِ:o�~#�Ǫz�}�ק��v�ոȁwf{��ՙ�*QKE��E�~�i�U��w-�07��F=?Vu�1�F��U��l�G�s�4�~��Y�6j���z�(�����:���ٺ�|��,v���zc���vzC�;�}.�>&dp��scLg�����q��,ʄ�|��oӞӺ�/�w?/O?k�|��A;d`9ˮx��c/�U��n�6nU����S� p����!w����Z�Wά���\��B��V<<@�[�6e�8q��;�o���0�t�.��Q�����q��gg)%��i��à{�&�&��p�go(��J�D
�_��û]{ݯ"�7L�Y��n;���:�I�����x'���$ӎ9}G:�4��z��`K���6��kei�z���ۛ���k9����%�������1�W7��(.��UH�����O*��7m�Ғݭ�-��{=}��M�<�5�m*�b��}���I�sZr���+��*��;�2`�0�	 	s��W�WU���t�i��Xbr�,L0{o۸�u�!�Ic	��P�=<�N��jQ��v⥼~<��"�����<=n��~��'���td����y������S���7����|.����9����s����~�e�؉�(�H�Nj�z�Y�XH���_�3��uM�3���1�-�wV~^ͣ�>_�J�J�Gu���S:����]�r��>��5�Ʋ�"mL���Ɓ�ͥ����-���i/�VQ��A�Y8�x��Ig5�1��eC����ձ"Ə:pa��6�S�-�l��b��f���^����T�)
/ԬT�`�ϲAok:bv���r1����]:�x�$Y��8��R�kYb�u˓���ioT��oS�ިC���UiO;���^��I�m�L�0}/c�Hz�&7�z��+ W��}��/�C�/J��x�Sxm�e�,�����ͤ=�2c|xw�x}�+�A�i�����-]SQ�b���d�ۭ��;W�4��ѷ�O��iF����s��{:8� t91���$�N>�l��N��o\��3""�q4U-ұ�"se�̺�`yޚ��V�sڷ��g�=!�?\�6���Ns݄�Q�e GUy���/g����h�9ʌ-'/��w�_�g��~���}�[��J Ec�CP���{6b�چ��./1�/��&w�zN�x����z���]y?�M�/�J�����[5��WzGgx�����pv����Kv*���!�^�g����ɗBV��57�������{P5�N"}��v��w�����+����o�=��v�qg���kv�\�_uN[՝���oD�cmG�-���b�� 7��>=ڭg�'��8V� K^����;}[kJl'r�����'��V�2�v�G�_\����>��Y������Mn��C}��1|-��ͤ� ]: <�/4�CK*q2�������#K2)��O/��7�"��zP�5V���K�Wǻ;n$WK�1t��z�m��v|)��ʡ���,��O�(��V��������1���̕��k�ꬴJ�WT({�R^|'{*U�9�-q���q��w����τy����1�������v���[�ǎ������٭�י��d틫x&�w���+�8m��hq�D��K+��o��q�3���P}ʨ��k�F,��/�OSd̲���������������Z�Q�cy�T�L���s8����]���y�i>���B��&/�Jl��zc)��lm�}��}pr�����C�{��Ve/�]x��a�����9�b�z������/q�R���>��y�y�,M^�z��>Lb�_���wO��������WVC z�Vפ���a��\חq�_�CT:�����X׮��_r��;��hJX��t��<�<8�7t���U�r0��_݃��D|�Ǎ9���4�6�T�{N��V��81HR�R��da�9�ծ%��uA�����ѭ��6_P�w8c��0t������q��4_�c�:h%�\q9��ݳx����D��]e�'�"��Dh4�:�]����P����mt��x˭>)'/Hiد�;j�c7�,�Qޞ�s$C�3O%ܝ�9�\T�z��{���r�Y��s�b4Ȉ�{��Y7�]�Ï�$��x�����2������PB�ˮ��=���{'�yR�6����x	���K�ڨ\^H��8m ��J+��\�^�껤��J�]�y�E!Ej�O��j��ܽRI�����x]f��c�3�}�޻-;�`'�u}���r8#ƌ��C��;��Z��/z�ES-�������1���A��5�>5u�v���S��]�w4���*���y�����:|������r)K�T��~�z�}SmC}J�~�Y)�~����X�������V�t%�[����b���Pї�󜾭OTٚgP�tI�������,�����AMB�'dm�pu/�#v4�o8��L��@�R�|D4�,;�ُ���F�}�_��F7��s]�k�Uv�j��A�x������zo�����D��J��Q_r��GΠz�(qɑf��h;���W���#ͳR	Ȍ��>l<�I�;���l�Q/��پ�'kp���7u@qǏK�	�:X��>�j���vb���/W��g��9��?{�r�gŹ�y�ï���j�9g�3�9��xjɲ����3��7de���,�Cf�8�}�m{�7ܝ-�>���~�z�����Dp�cF�w4�ν�ӝ�ǈ��/],O���=[���\iΟn7�[eó��=����b�'�������ыe�;��:k���H��=��[<m��^3X�1���G|o��Z����G��ֽ7���F\d���ɍ�p6�\٧7A4�`�Hw�P����������x����}����9]�֮(�̩�w;�UH_��<�o�!4�.��5�+),oHok�gv����F�{�iS�M���=�zon*qgP][ �3�b�A\T]0x�1ݙH�E�%�<h*�[�a"N ��_6Yk���*o,�wv�KA=�/�t�M��[�,v�k@l�c���^e�=� �5�z�o�+��-�N/���~8{~�hJ�o�vv_��4M=��y���f��Y�@h�y��J���|���`�����+�V��~^�Z}��q)�d
�~��� j��fW����ʺJ����Sg��G���<�G��(vЁ�NgF� �3��3t�WG�9(�[�ބ���u�Z#��V�UU��3��+��S�x5S��dM��o��`�K!!�4y_ϾD6+�����j:�bS������µ��uN2��!�L�Tz��X���fNߏ�r����m���Ɓی﫶!~��b1��kx-P��;��� f����{�9{S郶�7K�Q��]�������f$�� �{��)Ѕ{n_�p���ݜN=Սt��y���gqF�m�H�PN\k� �`Y�@n���dc�S�p�u�6>wYFm��Z�~m:~�6}��6�}�������odA��Cһ�T�I;Jg��Of�.�0u����{s�3E�Õ���T�x,`f�!݌�J� _�k
��-r�u���S^��T�bW��vHY�X`#[@��~4���C~��f��fwo���� Ԝ6���.w4q�n/o�!�VK�G�3~ۺU���p#P�P{g��|4��Gz{������m�rr�c�P�9[0,�hfBߘ���I��[�ƨ����;�Ӻz�u�wh� �V?��3\\lw�e=�{=��Ы�Z��#�Oj�'Ƅҽ�\���u[�υC�-����δ����c�6�-�Ì��Tǌ��5�J���NC<�l��o�s�|�r.�;�΋0��l���o\P������tq;��`5F�����Ϸ�����oWH��(63_X{��a�D_̦�ӵ���Q4���T��}ޱ^~�A;gR����5W���CUP6��|�O�X�t.I��J]]��}Y��K�b�����E�h�k�6���3<��[�Vo��oi/Q��������t�-�ø�r��������i�S��x;���v�l�5c�C�4�;��kzd�<�������B�_oǺmoqʴ^�����c�sJ�C�R�@Wʙ{dg�GZ��yu�Ԥ�7�5ڝ�dYX�:�6�f�s�7!hn���x�RV�*�L[ʬ̚k�Ju�n������;;��}�pնk�k�V�O��~��׫��{ɞl��=������/o���͑9��}U{��f�U��秽���K�W��u6��!�ӵ-�{�������;W�����7jؘN�y�3���'�S��u��>}��/��On߉��Y��q=S@8�?��b�Dv�E\n�i02���%���m�o��2�O{ʪ��^�ڙ�{�i��斝 A� OmV�}��c�q��~��$ɝ^v��\���r��Y�*�i�*��9�|�<��z��^�kɦ2{;J��a�w�y�^���F���7�������E�{ٛ=��(���tߕ��՝g�M�׺�w�qh��Z�}y}�y��jm�\�3����m����ձ{/}����k>�}yx�}��c�q����=��=���7��m�W_�!6}��#E���;Nz]�Η�^3�.�	�ÙaQv�5+6�uZ�_r�nE��2I��JJ�]�'C�uI�V��[2�ɋ��ǗV�*msv�\m���;_��yl��b�.�^V��
��)���W��@�QA]����Vb4���6wl�/H�I(��ެ�2��oV������բ��B�'��z�x�$f��)w�,
���O�6�ʴ�h.V���/�v5�i8���K�1FB� �k����g���f�V�U�)�$Uܔis{�%\n��> _Jw+{�[Dk�̖4�u�;][�$�>��"������[3���5v�L�psF��LU��6~<^�j��m��T�YLwe�R���\�ٓ@��t_ut�V˸�Gi=��6���PR���lPpQӊ���Y��3��_
�}�%*!�{��s:�)	Ks�ږEAgU+�=�Vfp��G�!C(r�Dt��GR3����l��&I�>W̢�8[/�Ζ�Df���p1�pU��|j����L�V�b	��ڃ���]�uv�*H��k+B�杼7����ټTyM��g:�}��X1C%�;��A.ԛ�;ɛ3V�5�x')��o&8���Ĳ�M|��.��Z�����0��r���L�ٴ�hܤX
�b
�I�nh�s��'��d7W,Qu��R�T�>�H����V��mu��Q뫚Nv����(��,�	��2��{:�2ĄJ�d1T�&���o��y�K���ҿ}A�w��Nq��/Mt�� �W�{�X&vv�]��</�9@�5�`ɒ+�����*q��)���s%�VA�R�t l��%�����h�WKi���l����Vhށ���Y(V��r ������I��<j��\��b�/SWD5�f̃�ǆ7�hVo������'s����v\�],V�ǩ�k�х<*�u
�6�Yw\+x�4"���𡽜�E9��Y;8��}�;؞R��E�_t/l@�Y�,9e�iwm[R+�I�� ����Iώ����#\uX���Y���� $��p�f��؟kה������S��d��Fv� �V^��\��GV�^�Y�[�ԩ@�p��>�ͻ�+QpC��4�����OĭTC��ll��gB�rgX7�;`��nZ�jZe��R��N�ڮp;1���jE���l��E�S�´��˴w!�� +&��t\z�R�b����5õybζ�슷��s���ܛ+�R����Jߤ�0�Wx�ϜX0�� �acOc9�@M;�5 ���Y�k��@t�.���q%���>0��[��Yt�[����r��u;�MKo�����g��sZ�9�Wp��i�&Z���F�D�*��7$���h(�{���9�%ǆ���9s̏yD��P��Ȗ�nO8k��ر�b�����P��m�U������l�����||||t�ӧN�N�:\�sǯ�?23�-�F�1��bSm�˜mm��& ���9�¹4f<�r�S Xƫc_0h��-���mˏ.X�r���y�5Z������>�N8||l��:�:t��Ǐ_���[lc@žm�E�oP��:կ��F��ef(�A;!�n'�qE�ض����\گ6�ҰV6ћm����s�8q�F�m�ܢ��bj�Q�
�l<$���b�5D#H�7T�)�ԙJ�_^��<�X��b�Q���q�5Eh9�r��T��9�o1��8�r�y��W����c<�bno<1�TA˗���Tp���(�ǅȽ`4^����<�1���W�1Ey��s�yZ ש�s��ތj|��p�9�3�$���9ǕQ���tTT�F���"*�ibj���+p�����=�pw��
���c�
=�'�b�s5r�MG�蹍5zǣ�=A�9h�DTEAM�yp�9�DRy.��G�"�[4<���q�1C��J�b �#W1�m%Dԗ������"<�(�"������+^���h������'9������*�:�yZor���\��/��m�w@p)N��W��˛�}�L�ʼ���a�;Z��+b�����.d�QGH[W6�M�8]�\��3�J��ږ'�z|'L��b,46�?7��M<3f&�
��kl̵]}Dy�ò���.Q��:s*0�r2�׏Ɖ1��T�p^���#v5*�����]V93C����b�s��h���a��h�7Y���h�A�2�
�e\e����kT�1aG��Ꞃ=:Z�WQ�=vm����@@��K*[����QL6t�nNbx��Oγj��������2�y�@�]�ơ�_+�� �;�z��C�"��&�^L��u�t�:9�5LM,���C�z� �sU�d݊�[J���9Ƀ�F ���3q=�a�;��x��čm�,5�������	�=�O׊E6�S��#3�O7���ö�a@<zD��W,B�U�6SwD�] !��?l)�@pj�l"��P�x�Z��&��{jl�36�Y9.�o4��c�i����C͏�L���JoH�b�O��/�3V%2ٮ9?�1yO��P�s�i�1��<:2bh��b��(y�fABVP��1~`������ni�ɦ��ռ�f�b� Uk��Ѷ�����-j�w!0�/�5v0ܝ���j�ed'p����DǄR��bR�5�w���O�ŷYlu;��Wb�Xl2�IzJ�!qҺVnn��Y�}ŞM�}�t��E	�]�d,	�Ϩ��gRɸZY�0F���R�me3(�g��3���e����٧��x�c�vK�D,w�`��5.��S�Hfnt��8�5Es�o/V��N��5�u��mZ��r4���s����`�s��(���kѸ���[t*��0�÷�z�.q��3��,�J'���������h�4z�R0p&����1x����η��b3���N�!��Y	q}�@c�}P�`+׻%8�'Ɔ2�p�t�\W4��{&!��8ml������y��^%��zZJW̪�	�{�l���X7w�HD�M��»����q��3e�g��w=��&+r/uo�|p�(���v}M�&�{/<03r�mأ٦-���q|Zl�S�Q �Vw��P�^8���NN��h�(K:S�`+�����o+�:Y�R�����c�Ƌ���Ռۋ��9�j�{f��/p��T����)�1�5�x.�^��z=ʩB�\���{2F!m�����Nj�0*�YQ��}9pn��r)��I-�CvZ���r�H���߁�*��s��hq��Ƿҭ�c<,�Ƕ����mo%P&�N0���H�0��_��[���$�H��F��7��8/S�ASQ���ms�$�|�ö��׮�N(e4'r�ڢ#��3OZ��B�_"T�tk�[�xo5E�BZ�y"t'���}��#e�)Α6R5� \ʜjp���y�)�M����z�%h}� ��}u�ύ\$X��S�H0�P��`�@���f���X޾���������|!�b
|�T�K�� mD����c�@Y�O�0��%9�-"��t=wY���Yz6b/j2�6ьi��=�i�ħ,�D�
� ����"|*�)��ȯ��������u�=:�y6��c��s��F�k�+y퀂�_����^vi��
)��Q@��'��$�^z�(�W����E�.sȪ�s^m֣9s��@`	[9�̏kȕ�۪mI��~��i{�DY��e�o�mG��.�`L�n/�j9��5�7Le�*���"�-(5	r˯�	�(��Հj�Q��"����$��aa#%��20��m�\���١N��` U��g���P���ƚ�����9g��3wP�ڍ�}y�庈�=��;��F��ftOb�n#���ؕ����i9��K�C&���{q%C,g���Y1���Խ����{��(3.qc�Ԕ��㩃g�>fp��(l~pɫlTK&�
1�>G'��b�����[�z����V�GK�EJ��ƿ*<]"4�!I��ccЗd�l��UT�����v�X�[��{�7��x������,�B�/��ݎd���8͠>��D�&�c�%�������W�E���K�7A]MV�|�����m�U��Kq���.C�.��v�Z	Ow	�PF�+�1��p�k��p��RPc*��}�
ZZ�o׫�޷G�|*L.!!�9}Y�k ]�O��� E��t�W����`DLaq�}�5�mtY하���Ӏ�vN0Ȇ�������=|\5R0i;6О�LGE;���l��z��y��%4�僵 &a5�/*���B�C�x��-�eC���e6�Q�LM�U�(M�;YY�RVU�N7M,�^��i�5S�eG����e�&�V/Em��u�<HJ�nVm���G�Cw�R�4 �54.覒�C#1���9>怡M5n)b��_i�0+�tY�]{����,��N0;�<dN\\��Rf���
��BT������f�vH�N��o.��������W�0a��aR�W��D&�&e����3bK+����Э�S�Ag�̋t9���\��ʩ����F��P�6C�t�H�Ͼ�GM'L1L&w�U� Z�m�L� �C�vŴ���XY�94��5�v��0V��e e#,x;���B^�s@��s�Έ�[�\�'ְ�su�k�Bp�<\X�M�'��ϯw�����sϒ�#�Y�6+��R�a�F�Q*�;'�[�dn�d9��#����f� !�f�����[����#�-^�WF����>�wۣg+5�ޛj�kAY�y��q����1�b�^�6���T�y"I.-���^���Z��q1�&x̷�����Ī�e�F��m�����E��g�w�<����ַ�l�θ4%����~i�3��!����m��ǣ����5��2�bv��Cկ�a�z;L1j�p��'��@\���F�i�63�D�E���=�4�vwr|��ߚ���z=f���	�i��1���d�%�5�`Ky���Z���]�3>�Ph�m�:����B�ZCڝo&����u����z0�
��QQ�C˅g�g���wmhuީ�{r��Ɩd���K\8o%М�cC�$D
kiȎ.zG{�x��?�%X��%�|Z'�r���߼��Z{�W�-�5@v���K��c3d��|�.18�zNxQ�c���C�^�:�z������_]�W�ք����	ڣ��N��޻��Tݺ�ל����Vt�׳:�n�ݴG���Ù�â�i�����D�]B
�?U��w�?t˺��5�Ɯ�B��b?��:�t�#�����S���%4۝��7�\��+��4?���[*w5�FV~=:���j�������3'�tr41e��4����[(��D��[���k�Tz"����+�����FK��c�I�T���/A��ck�:��M<Y�b�;2�+ 9�k;��5��ڹ�� �ĳM��`��mLTy8��^��>}���N�N0�v*���Y�*�9�jǙ>��V9�B��#76܅έn�4ɤ��*ovsm�NB�6K2�l�@���\����y�Š`&��&Gs9�w8�˟5E'8�KbQv�����Y��}�E�jK��Ե*�m��N��m��-M��	�����cXH��+�U-t���b�{^�W���o��g���΍أ�;nun3x��p�5HR9���H�3�>vO�24��f�Oӭ�9�1I�r����4��cJ��N�s�P�{�V�=�q~�t����l��g����2Ж���c��Ig��=���m���ۯ+j����a�Pul)����`�_�ɸ��y����y.j�{1u������ˋd���q��d��E9�BƉk����Ma�s��5"�@ov���S��l�,e��uNY�hțg�g[�?-샬n�ѭ�JQ��A��mK�z���OF�쾓������M�2��EEz/>�F����OHƣ�"6�j���4�c�};ya�4�ܭ�\���3[��x�ؓB���-�N{�/�fk��>]�w,	�a�xv���f_i�[�f���ݟ���v�|R53g"�G��+�)��?{�cEB4{*�u������F(�.��ٻx��u����G�I�iV�a�#Hi4�v'��m7��u3�9�O�9}�2���;��1g�%`�
B�Jk�dE`մQ�.t�l�Y��o3_�%D#��/��e��Ѩ:�uL����]��:ed��iӛ�ܖ�
P�C�"�EH�(� �T)"Qb�W�����?p���ʳ�yT�.�zԏò44����-�89��M3��l/Ţ��[�yv���̞CZ�*���>������
g)W��qs7����4���O�u���>�:!�^̇� �}=l۵�Vi����-���[\���N6��Q���Q����=��(�^s�K�S�j�t�����͸��n��\)�݇��[%�k;���<,� JX8F�c��EL�%t+/ګ[�dí�
]��}1sW}Y��&�<J{l�%<�,�Y�<��ip1?4������9�q6�	��SC�nnl��{��c�<4�j�w������t��Wʶ+���y9f�S�6����gɵ�!��'����%�[Rs{s�q+��׫��=�'%��`i�4ļ�kp5��T�P��]^�4Y��8�+�S(|��il��j=u9��[�u2���8Ͳ.WG�WT�o�U�&�T�asv'mڡ������6tL�+��;'v���i�먹���;�1���2� ;tw@H���L(tƏ��9R������c���$جz���[0��;S���#ʞ�ư�c�(E�B�~.	�:�A���d�� 0>̊lj'}1���H�Bj�5Q�J�J%�%��?kQw�2�����P��5��e��!�[Ȟ=<`M���ݷ�.�X�Պ��R �����w����r�LtO�.���.�����>��k��V�::KF�e��U}���l�*����wD)��~K��r���q���V��3|��������q�*ѱ�S�Āof�C�w<y�Ғ�p[��<�������y?4D�.͉�>���gM��vQ��L�k�~�X.j����ZL�����x���ʦ�u��!��h��]�M����>Q���&� �����8|k꓌.<��Y�&�fT��f1e�]yZ�����
�\W ӯ~4}"M��v���� 6']�D>=�;7+a1��|�)Xs��;/<Ye-������g)O��C�MD��-�=C=�;T
�k׫�j�W:{���S�>�1�*F���Ү^�ZT���~V�2!1�"F	M���6О�a�Ⓨ~މzO�E�UWuv��t�Sҝ�S�xH䘏5=E����.C3ۖ0��-�eC���5M��;�F. ܍xW�J�N�C�S�)�e�2&�'���[��L�R���%�Gt͖a�#ށ���*Y�0�U������\��Lxq�-i��u�*f0YSS@[��mB��4�}����
i�L�#�Ev���=;���r�%�m�Nc{l�7l]�[Q"ݙsϒ����f����\�nv�b��<��|�;J�^�<wm�/{��+ĊK�ϴ��I�R�ɣyq�A[� �r�%����w1��:��k����kndM˫R��Y0�$��T��ݥ���g0H���mB	\	�6]$�ork1k�`���{/�}��r��r��$��6�;�3��:�~f���>�e��S*�|Fc��bSN0)�^G��\O�ƚ�s}|:X1ǉ˼�+�H�a����|�={Q�	*8��酥�I��)�����k[e�8�};� �:f0��Ym��Oo�0�Sp˃x?�)�b���x�ڄ��7ʊ�Er���9�,d{�ر����r1Ȓ�NN��7,�z!ò;�y��&#_g�U�k�;)Q���@��z,B�mQtZ'n��O;�^ɥy�ݻL����*�"�q�|mi�0D����8�}��W?�V�����H?ڸ��z�NAs]�Ou���T(�U���0.N8f������&�&:('6�<逯K�sb�c�+�[��"34�(���y�"�Z2[lFNןN�;Q0�qk�#��cl�h�a�A�t�(v9�5�#n�ѷ��k���|��H7H�X����^�o���g7��A�F ��lmxT��y$�V�=�ױ��X�4��S�Tbz��R1H��lx[c`�<��eCW����y'A
����ٔ���=��ދ�>�**�����e�����Q���P�0�dm[�,I,Q�`����5Ŗ�m�s��r��:��)Kr�j�^�<x
�u��Z���ƪ�mxeC���+qҵi� UX�o�>|�(dAԮ�1��3r���X,�{�6wd�zJ��lMUc��,s���n���;������G�?�ǂ�<x �^��}�Y�<�!�k�"��-`�,k);T��������4���a�����0�0f���/sw3�jJ�=L}�ʜ.)�sP�q�9Q�h��vmR.H�z�-�FB/SQ�oH��ۦZկ&;Y��Qx)�Pd�xc�M	��ͫy;U���yZS�R�yNC���R���^��K������dp8�qw#,}=o~��Ŧ�K&W䲩�Jq��]�vK�މ�o����gMe���]2��Tk>��[���[��Ηl�z����F{Q�N�c�[e�{�eV��ba��̱�)�:���m�,�>`(�[ �`h���4�R~os	�U"�bQ�	��*5�-y9]2��m���z����ء������H�9�0R���KHC'���h{A���5���D��	:�����M��qO=c�ޑ������C��U��o֖L6N�&�-��T�[doub�C�����9�c���\ߙ��$��N����0Ƃ�$����t�qͱ�4Rf���՗�G��K��KH�]��~�L�-�7\���9��s�7���c�4Y�V�$7���~��Ԟ�WWv��mkMY��A�U( ���SY�+w�V�V|��]��j��S���ϰ������Y���[L-�r3�^�i�EL'z��;-ɯ�ne�5��7�Ӳ�pn�F�[�MB�9�Xu>�����e��z1��amB��-�Y�[�cf���ξ��%�%�㨰��	U��<�� �s���a��RJ�owyq�tI��V8�a�QPWW��;0V i�ub��ed+Ř�(�����)�I��^a�4:����:O��҇g/\�G�i:y&���N�*3� ��tZ��3Ya��C���w�k�ܬ���ze+�!��&gf&�r��B�r^I����y9`/�`�`\f��1ؐի
�; ]B�E�j�!8�� P�wT�;O<��+��D7>Mݗ-�ݚ:��#��Y���Ug�Dڐ�;x���L����J�[=})�M�斂�Z�^����Ő�&��)�(t�x��ˉXnS����g.�n�89�s�����[S�ʱ�һYIu��5Q�n-qۮ���[O��;_u.ӇbZ�z���m�f%m�����k���|���W�v�����< �1T����P;`K��Ke��'c��;����V��gv���;%��ò��`�H�ۅ��m����D� �����|�9$���u�p}�5�GZ�8�mv'OH�Q�@ѣ�p%��Z�{3�,�P��=d=���fC�h�t>ư�y��N��-��扥�R�T�#xX���ELZ���iФa�E�3��c{�/�۾t�k�'�����K	)-�r�˰��j�A�28M��7c��E�J�l�]lnq��&��i�(n��p���z�q>|���G`v��3ڄ�(+�9�(
ѥə0��N쮽cD�j�don*K Gjޢ&ުu�K��w���K��P:��bOjN�Z���E�r%����fZ��Ҳ���zj�,r���uΔ����*=u|1��,enY�;�Ĺ����*c�˖ɣ���N���]�\�J������|�MuC�/X�:�kMF ��y�(Kwϱc4>�M_knX�Y���j�YPe��R�S箘w\`ܼ�L�R��db��������v�H(.;Κ�W	i= �g�̾̂�*�g<��]�eweAǟ��l��-U��Q��
B�qΙ����X��Eve)�'a�.�P�� �)W-�
H�o����:��;�6����ts/�-���a�A89�3�z*�)g���ik������j�a=�rՙr���/�1�j7A˩�da��ݖ5l���:�t�5�wQ�҂�'(;���3�[kK���k�c�au�Y�zm�;!��`sr��Y2rxe�]-E7B�,q��GZGn��S]*sJ���Gb�MN�����v6����7G4z���I��uDA���*e�Ӗ̈́�|"�
E*?;P&a��D�./^�tgڡ@��l2H��`#A�D:4Z���HDF¤R�@WD�Mᠭ��4B���p&u�܉�qA�+t������K1��=#��S�LQ�M1��߿/�(����գA^������s�>������^�ׯ_�������?�����Ǐ����).j���H���*�\ړ����np�scl�'�`�Æ�:t�ӧN�:t�������x��������j}Q�MQnq���q\�͈���km{.sE,AG�8���KW�h孳�Ms`��V�^���)��`�%6�y�3k���g��"9rA�PPQ���AW,�U��N�yk��(�8s�0TG� �� �Zjf���*�����<��UQh4r䜚B���W<��"-�O��W������Zq��v�ئ���t)���f4�ձ��Mh�V�l��6K`�ׯ7�夈���s^sy�*j�gc&!�gb���To2�^r��i�3��a�C�g�5QUD4�%4��J�9*Z��9�5�ђ�`��UT#s:��4SITUSA����4^[�������Q�>y�/Ԙt�Fp����i��Y�sїb�	}{��G��OMk_�8��;���R���k�QN��n@�
��@U1�A2FT(8�P�sC�����x�S�~{����z�c�	3.���aG��`�+���20�b.v��z��oy��{!Z1�6-�ۊ�ޱ�э/����71�dqT/3�9.�g�I��"B�wf�K��<OPƭ:�#h�m��^�l���Y���r�:���r`�g���;2q�ғ`�(%�9��0K�ׇ4��(�B����j�ژ���]��n��Xrfl�h�`8��3g2�B�	���>/`Pt�M;5�R�0}m7�oB��P�u؎�g!��� s>㢠`i�Q�b�E�'�t����U�@~V�S�����X�㨝�;.��=����Mi�gBfo�ٳ�]3�X:<ڢa�^^��b�@s@�z�>�7�)ǳ_��1߿|s<�4���	�q��� ��lpm���E��(�q��>98�����|�iȄf{�vs��xف)z1Ř[
�p C�սc��2��P�2�)���S3��~QЪ�~��6�^��BO|}(�����,�`�xi�����sv`z<[[��_��ra/�x�a�~��Zq��g��s��W��)��R���ԃ���:��Gt
���G�i�����xJ�ʈ��w߈l~k*i�
ܙI$2�.�+��"��F���.�eZTۮl�⢷�աu��9F5ժ�cJ�s�]>��&�*t�}��;��a��v2�����q�4�*%,�+�pF��{�\Q5���}ƞ��wa����.|�>-������><L�<BB`	�ۗڻ�8�j߄{�����V (����
�+HK@T�Y��Z�!�I�{ piVi!3��z��r�pl=Y�z5���z�I����᮸�1L����>��]���y;%�R��40�^�u\��1v���w?!�h��:g�Pz�)��RX/��D��Ԩ���c�!���"��6��I�snٔ���j���g��p[K�y/"ѿPb��,4�T0H�d[�X%�m�V�a�c��滖Vw���B�����Η ��6�6�i�8��|���_}�5�����;�։�g�3�Q� y3gB{-�kgϴ����(n���Z.��Cf�{��4�zM�哄�AȀ�{/�gcy�8ߤe�#|��i5��mxN-���ŝ��@w���,�M2ǁ3l�0���s�x�n+�y	�p9�F�m�S�1�Ba�pͅ��d�Tla}�óծV��9D�lpݐ���$�f-��C�f��/�&y���	�-F.ZG��;+@y ��t���w�`0	��ڧ{!,�|�&8�T�=ӈ�򺺄�A���KBfޜj:��m�>� {��3�;}�m}�a1+vA�{���7|�YAe���.}�&�l���P��U�o,�ʠq9\�-�&�ʬe�&O{�	�P�C�Pؤ�{�%]os�@��9:��a�k$'
=�˒�2遛A���]*^�0�]��O�..4$�=Y��eu� ��)z;�|�ؿ`��xϏ <g�D����N_p-	Z�Rz)�WE��]�q""��o�ή�Tρ�����S��嚇C�KV�����q/�RK?�o��"6O�c]�g��f�O֠���.�~i'���W�NǞ��ۗ\�J��NG�,)B�}�����˧n��)b?*����*⦱�~�S��P�v+"[�xf:�)۪wg���}p�Rf����b�� �5�~OpU)q�"�ߜ(W�.N����u�q�츥�2[�GDW~*��=�m��Vg�Y�;;��+�\\��&op��!�8�G�\%�5��r���z�%���]&��W�l�`+�^&���okZ�\�6��;}Y��7��0���Z�1���}l�n��݀���|�I��3�-<z��Q^�����j�C ��x�e[n��)y�9�g7x��\�x�3�~`6���)���ޣB+Ī��̵�%y;S]ֺ�O8�P~��H��ɧ�Rw��b#ε�B.�ٴ*e�}jD��^�=�GR�Ż}ڇ�z-�����{�X�{~�;L����8�С�D�/!��2vn�x��q�n��I�-t�m��o*>��&�s�m[Y!"�|J�ĩ�}�s�%N�݇��瘒�H���a$^�=�������`���'�X��QΧӺ�:�ac�ͬ�+Auw�w=�8�t3 ���s�^}�x��o���E��(�.X�r U��sDz�8������ ��"�n�~��	�E��X��y��5�Y����.1�-�מmJ%�n:!�Nv�Y6�N�����'��Э�:�=��x<qQ�N,�A�Y�`_��n�B�)�r~��*婏�!囟�kivp����y�	��:��&0�c�%Cdl���66@��z�f���H�����|����/i�;Yn��S���@v�7%�K�TP�fÙ>�q���[7<[�y��q~�@���_��(R��P�> 8j���$�pV�h�~hxzm�;��vO[k�)�[��\��Cٽ�ޗa����;������׳����S�¦-��b�D���C�D-��Kz��>�g�ۨ{Rc�2�.v��1m�̞	��;PՔ�'�\DH��e��ʟ
��ZNK�MaʎZ���[b�	<�u�4���r( ŨY�d�h��n��6�����FU�=L�[ۇ��e��!�b� ��K�s��#Z�a�
'�R3��W�9�}n~�����y󠲏�����I����-�ړz����y婥��@���̽����;�D�Z�T&�*K��k�f�ȶ�����r��.m���<��\U7H��MѰ��{s�}�*wr�P���s,qC��v�D���z,�c�������g:Ä��>�Q�3�42YGI	;t�;n��3�}S��c:B���;��'9�y��e�N�PWȪ h�$�N/�ﾯ����K�(�b���*�lz���]�rֻ;�42�\W�|>y��;� =��HS4�Y�γ�|A���ŀ��&%R�I���6ʆʶ�ۺY���0��Nb���49�ԣ�l���˻�N0�����-�mkgd�l��ӡ:Ei��GY����Q��=S�� ��}H� �6V���0g�q�!��4��>`xE�c&/ذ�{ZL�u7!�il�dJy8�H��1���r�1k	,��ǭ�Z�����,v����*+�Y�*�h>��8<�b�R�˩P����@���<�+ݓ�A͙aod��Pׅ�b2;V�כuww�����f���f�0E75.4�Ɣ���>/vR�@�dSI��gn-��9��=:�W<���0U,?���hp|��-A߉kd8d޶̸�3��b_NP�>j��ԑs�*�LOVb�~����P�T�'ƃ�Pr�2�f|N��L�V��tvk�#翞T�������ÿX]�e (x�q��x��3S��S䦀�,-3�'�h��t�傝d$M���~���N���x��v�1�̼;�B,s��b��#Y�*N�Pi&o}0�jG��Hׄ��P<���*����3R�^=��Sv���~w��B�t�mJ�@�@^ON�;5��w55X������cQ����9�ZNv�Y�R(��\�S#�0)��;ê+��7:����{Gu���=�ѫ�(���?����3ǂ"/��������.	z���5��]�v�c� C�(A����mr�wp$��qhڵ���8��)�߱~�H���`1?}�q�sb�h.�WS�m�R��r��O��<�� ��MЬ�v��K�ȓS8��-��������C��mC���P��B�kCU?�E!���A�@MMGr[{V�PloOF��Vw����9\r�ב��F�3���M�!=1q���{�\H�@g��Y1�i�y8ef����n�V��[�خ|�^�+�9d�[㸦���g �j�F
mSыdŰ��ï�f�P�0�ĸf����{�/<��o�����Q�E���B�AJ��{��=_��Z[ނſ,�o\R��F�� 7��`�k9��i��\��p�a��w�@-���Jm�S��
��?40<͇}w�CM-�ͫ�%�!�a��qͼ�o)�ё|��,4�U�-#%��9�asF����V���N�<���˝$�B�����dþ ��[r�X��]�Z�@/�k;�	���邧l�����[���kS��} kcK�k3^�N0��f�P��3����OK��Zۭ�[�,����c�S�sR���˂�C��:�a�@�V��t�sy�w�(����R0��w���i�wYwwwW������j1��)s���������4;���� �gF����ϑyvpw]Euը\��HN��5��i�ߞ�U?ng�<g�_~�	��u����a�������-�HL�8�p��ja�c�L�~�}�aq$nʪ�Μ��)���^Z�����	�j��y�^����q�0�}���f�~��� ]��t���z8p��s��6��v��"B��k�^;�5�Tp�ʰ߮xx��(>>7\�H�.�7��#ۨzX{D\Rg����"�����-ـz�����X��$#
�'�����/�ff�����iwEI��KL���21�3&�O�0����&%=1����PBg�ɰ���owYyX�q5��KE�����p�� ;t��xk�@e�)��N�kD(m���E9���R[g%^�օ�2�7"mQ�ƀ��u�*ff4��-覡%�T;q�m��
��έ���#�ޖAGM5b�f�5z�K-���U�
����<�T���������K�BO>�I�G��^�0;��f0]@�<&�d�v�*���5�m��V0�9N'2�X�h����xb��2M�[�e5��L|��O��<��H��n@�s�$-x��+�z�7rSM����9�ُ�Z��D���;�M��D�.f�ڕ�)��n�#�.�]�Ԧ%�h:�[S@w0���'�@ *��7W�&U�:��4{��w�*=)�m-'���O.�gw�.�����hSk8��k������Ͻ��\�����?��><P�<P@�k��Qݴ��^�}'�66Pg� �S�	�\�}�qJ����8�1I��*���!ٸ�D�gov�Q�yj^�>��h��r����&���q����dE*��r3��nc3��1��*�wc��m�=�<Cͽ
�!�e18�7^J�`���y�t}Y������%�o�Ci�qDtp까�7+29��=�q�,�0��&�Q@���P�h�ƙ���������/�Y�M�[�<])�%^��7K�K�&EJ5l�倭��u��QG��1�{�q%��82l�p�}Oͫ�B������ߴ��f�<3��S��m
�yU�md��9��^c��cT��+z��!���dڞ�0M��r�-6���#X�Z��N���zF�&F�l��8����=�]��%�1n���r!��p�����!��U0��u�>Y��?k��ɱ��}��ͭ[Ѱ��CӮ9�C�o2 ��qC����@M�0�1�|j�t���F�~�>y�C� �3�La�N��w0C���:<;���;�f"�������-��_7��&�Sg?�
C�|��C�����d�ٓ�x=�	�!�5�����@�Y�����y���.���𻷔��e�]�ÈO �LA���ҽĠ&fY��q�Z��Χ�k	�K��@����)���/��;2�Ι8va�S/������(��|���*1�y��߰T�����T���@L	$bH���^M{�!�(X�I�!�<�}����p�#�C:X�W)Lڧޓ�Gw��v"}�1�'���n��5O��ư*V��ȃ�(��]	���+�p!(�z�d!�r��ЖU6�?�Y/��p��՝�]�xj����l8/S�T�Tӭ�a	�a�2ظ����t�^��}XUn����c!v��nӄ�!_���Q���d�q�/-M��R-��О�`��*ziZׄхjez�9��v���r-�`g���m�5iɸS�s8d'���0����-��<�f3��ԟ:�p��eu]ݝ�s^-k1ps��6��G��J롖'�
ǜW&�a2���;�ײX<䛋a�Eg#Vk1җ����vFl��M���r�c���hૃ>�ԮШik~��� ��S���"eE�����v�����to=xv\�M~H�d�9�,;Ke�c��!�j�g�2��F�f�_lճ0�{`X2��<00��su�U���m������=l�ľ�]�]��-�TS5�ӧoO6'��kr�1���7��r�������h�R'�8��=^ۡ���n�[1!��vCt���Ef���wJ�v}���}����X���=瀟^��@����&����`u�����t�g5vm_�����u�����4�}{\�J�J��3�-Gt��S��ys�f�O"]8�]�74ȟ|&嶺=<^q�>���~�_��|x���<x��`$\�Vg�29�o8=�9*q���"��~LY�@3c�[�4+�.��)�3���e�rr���w��Tv����x����fK	1Bc
�f�/��:�އ�;�2.��Oy�7,�4m.������@f��S�\ށ��^�001U �`_�qd���+D3Ζ�_x�������u�h	`���j~�"�.�%W"/�y@��)A�T�e!������T�!y�p��">S�~~,���P�6���T�SHKH��l9D>��f�,��tw)�Z��sm��Z�LI"���r�q�q�J�pw6᳠L��}�5�]C�?~0]VP�j��=���o��X�%��?n{�[�	�%�T_Qo.ޜa-7�ueػ���55@e��jv������d45S��{؊���p��^�����Ú�_/�x�(���8��M�m��E����ɽ�� <���GCK+�|��>��;_|���.��-��=���&�
�jffT7�2�X���J�!�y�ڧt6�n�{�e�M���a�4U��Mtpߓ��e�R�l���>�3�1b5>xY=*���N�bm�e���u$��R����]�u�f�1��B�x����ċ����|k�����agV��N��Aǳ������J�
f�GR9a���>��I �^�SK�T��������:�Lȴ��b�.wqڻ�h�l���]b �A}Y�T��ihJ�ja�ue��
QC��x�/���Q���+'u��Y$մc�sc����$�j����s��,_�Rur�![�qMa ������{��\;���k_|�(���@N�_V�[�PI�|0��y�.�sx�G5��T*���Y>����s�-ࢪ+��{څh�z��̇��X(u�%�����;I�l`%Q�ݖ�f�B۲����G���:OX+5�n�r�,�X�L�t��^ �I��h�Ii��n  iX���Z;�Z��0�J�.�{�|�Ѽ��X��i�;eMr��T�&Ƀ����;F6ۤ4�tn��T���륿m8��6�"xˣ�[>���8^v��<�Ɔб��;\p�[�L��!���<� �)vi\��:
vg�㺲������%H��Г�[���6�1���Y��� n��n�H�ަ۹cR���蟤�x������6)�|Ef�=jK|�c��y�X.��}ݞ΢���fQ]B� X-�Ϲ�W����O)^�Ȥ�q�b6���pC���i�}���uC�E]p8�̢2��fQA,˦)�E"���o�T��Bƾ{�V������k�|��t����&�PiЮ��b�]�/�HfE��jf�\8(n�;�r�Ǜb�]��ܳ+�w
�5��.M#2]!��m}�+�s�v��7�5C_Z4J6��i��Sd}�I��H3+�V���7�r�
�G�۵�m��{5H6�8Bw�̾�Y{`�ȫ
^���8C�}���z䅼إ��D��)�W��EᎢ�v�:�}�82�Y:.]J=k)�q;\r�v9pA��kkz��ٝpcq��FӔ�$۳��xQ�֠��\��|�bˤ��9#�K�p�Y'^ �Vg,�m!�ZV<I���[�����Q�ν�C�O;�vD�\z��Iٜ���-�]Գ������j���].f�hGs�gJ�@'toH�.��i/5��2���M���y1yu)X٘�i[<"��;B���O$�֬�Apъ@)"6U����I�t����{q�vxt֫&���劝��L��pڥ�.�<Y�nc�zn1�Gȫvf� ��<Й|�u���BSk�y�h{����<7�H�a[O��f��W������1.X+��ѣ
�#-ŝu{��Y���YԠ6T��s�aH����]ڳ��Bv��6����3l��Jܲ	�0���"�1k�;'/Q�3�EEFڂ��jM�.sj�p�T�EQ�(���Ǐ������>޽z�^�z��������?���?���į-)IT��0G*4��4R'lj�i/�C����X9Z�)(>��O�����N�:QӧN�:t�ӥ��:|d���O���QD_3���L�!5^��d
��9����b|���1�)�y�
����ƋmM��J�����ms[>c�0RS�|ۄcgM�hb
�C�(����f(i9���jy� �(��(&�b�X���F��J�jj�* ��mI���y�9."���J&��9�L[j"
��Ӥ�t��9j����i�Yhhҙ��<����AUMQG6��XM�4[+�q�1Un��cy9������&`�=[����EDׯ8q�U�PD�^l�j���P�[d�uS4cU�A54Ѡ�%P�AM	TrS� 
�^�߽Ӻ�~�/}ک���SA�X�0��L\4���
�"��[���vu�v�(�G���;�V�w>u�^DT�f�T���_@~X�� �\�r��	6:w*�[Z��:����� �2�d>{p�a�c�ۚ��k�n�iR�/azaЖ����"��F�k�w
"XD�ۘ���zǔ�iH�vg���<¼�O7#���-���S���]ٍ1jXp�zo4��d�R!��k�.L�u�DD���Z2y�����ɻaO[{XTb��Q����.RqE�-����v���r��G'��S������[��y�<sGE�� 7�oH��"�мuQϲ{.�}^V<'��(o3���򢶡6�����&vbo5K��e��-����O���wAk�g��<�E��r��utl/0�3���)�1Uq6-d�{�z�!7+a���W��Մ��}K�w*�~��+��D�y�^䮹�9�x�PgN����"=�-C��6*�w ��U�E2�*�i���8���n��j�H�Srb�U闵L{�F=�}Zi����׳�q���ǡ�y|�	��N���C�����߮~Oڭ6֝�W��j�T���6�A7N����S��J�?	L���AU�wC������yssKJ�c�Ȭ�ӛzg��G��g\1h(u��"/�/�rR��τ��5�CU\�v���}�
��O	79��7����Ժ�Z>�A��'�PT���Os"?ʩro��xa����{���{��{��*��?�Ҭ�<
b bH8�}�z;q��
���#��.���C$�	���	SP	SSK�6�P��4�E��Wd#Jv�޳�!W��)�h�馡إ��<�,�2�	V7�z�Dپ�wP) �ڡ0!U,�l��v��	+��W��3#S�q���I�z�ۋ�3�F����"�-O�����f|�\�P6�sl0�̘F|�IaT��3�oO�	�9qu����@��+�eQ����MݞJ����Os3�Q[x�#w�w���T�k�=D_��ngƊ��E��j�`,���CT�๎/3�0��~�ќv�w�d	�\��{���ӊN��%@v���ɻ��N9�O+ZLy�TI۠NƱ���8���xVw[��
"P�>,������ڭ�!�{�6�yj@9|qp.�y�]ٷ�\��!7�s�tU��Z�GU�c!�%#}OV�m�v@�)S~J9�2�eV�f��l�M�P�ݤ�_���ǧ.Է���/7���Y4���W��߭5��ڨ�;Q5���-�&݃��u98�Nd�{r�<��L8C�|��ի�ˁ\�aų�}�t7`�O^Ȍ��C�x�vKZ>�ۻY/���o��c�|�޶�7[�Q�J�\�1E(��S�;;uu�[[7�s�	DV�"4"��Wg�SLYVJ��i&�Ƀ2�9�*�S�����+u�)k.N�Y��t܉���8aw9\�k�
h��ԣ����S����nB�A0�aP4��z��y�9�U?����	��<B��`&.�m������ԙ�FO3�_N̛0��y��@g�Ĉ�� Xw���AJꝿ�gxi����;��w�8'5Y7E��,40�� ;agf�-�!2�5�%�83*dH�/��x�9�a]�W�r 		���	��o�wܱ�^,��J�ȯ��t��*����j�+�M���z�g��y` R�@���e��U�����u���e{�8�8���C!��s��s/nr�m�W�3QL2k ��o)c����/�O����9NDE[տzLbM7o[��ꮾ�J��^r�[�)K4g��{�щd�~'*�R�R���p�����V�goKQ�x`��Y�mrj��r9�m�e'�+Ň��T-Ec�u��)�U1=��&5xsZޜǦ�Ѹ�ϋQ�zi�p|�������S�w?�ܬ7"��֚���[L���Mk�1�O����c'kH�s��Q�3����A����&�|R�V��� Z<+���z������ ���fӁ݁ui�r�ؔɝ�lCP�g�f�c��<9�S jb�W����K�m�33�=��6k^�yO��N����E&���N��+X+'-���%yβ��n�f�o�W.��X�b��c�������tf@�eg!�u�i�ɴ3�[��d3�I���hc�]�j�כ�
���\�b '���F�s4>��.��ɤ=%�!�z�Lv�Xo9na�����ے1�Ĭ��vՕX��Z'���k��<��M3�t�>��|�<O��E��]^�e�d�䌚t�̏,g��0����5'23�/Y]���9o
\�ˢ���/=d��(]`�@1�5��p"�d��|�����3V�vb�1���l#��٠
�C����{����T�x�>xuߘ^�~���镻U��e��a����ӭi��&p�5�p�y&����/�q��|ng5{6�5��#��Yy֪�^|&�\�ވ,,tP��6��@eT����_�q3�����{;��������e��ɶ}j}�������`Xi\��b-�=ywU����uT���q�s��<����*-�����^l!�fqO���>�f��ٰ������--�x�zK;x��/6t/Cͼ�@d�������[B�ȳ.юX��-����jD�wXe�d\K雌(���M�g�<�2Q��!����K�]8�@m9�L/�b�E�9��n�Wˊ�u��r�������q�!���̺��m+ʝuƦ����GU�D؝��:�hJWrF�M�35�%o^Iw|Ȥ0U@�cdN��Ǣ�|��]���))�:��Is���䷴�S	�u���R����F�ZCS�q�w0%q��}��-�PO��(�ǎx�)��c�Z�t�-�nv[����kxKa��z�u�
T���0�`L�p=��9�&C�����6��2��@s����_\��=�weȻ~�vj�7l���XHۉgn.;��ځ^��x���\�9���n0X�#zГ�ų��k�㼬/���~{��`Vޅ����<��B�Kδu���v��kI�p��P��A�Y��4
��z1�蘦\��)�O���$�d�e3�ܤd3�& kAU�'��XhC1ӹh���3���|�t�E�!�i��z`��5)������,h��wL����~���;�6��}��z�ᱪM���%�Z2,��{=�Qm��g��'.����E��@0�Ŷ�s�BMLÕ�ȇv8�%��\�s�ށ}�������fƌ��{�[n0�At%s&w�׼���F��ƨƓ�b���Z(����T�����~��`?�<̶�^��kN��UKya�C�{)��d؎v/M�0l=��w��9�<��|�:��5eU�]����F@{dj�4��0ӏ��wAkoQ1���P#�	����ó�🾮P��53㜨x�؉�j̗���1?�;��������jnR	��mJ�e*w�o=��>���Ny���y���}��X�ġ�p��Z��~'`�O��}��#����}FR�g����015s�L������튨e�K^f�=3�$�����K1 1s�<B�J
P�P�����߾�^���z�Lt"�%ؾ0�X{o�^S����ǁ����Õ�fz�$'�N��nљ��V�T89A���Ď���!4@��r���ah3w &��+h�7���f�`-�֝�V+@��C��3l|�m�ƪVt�e��g�JG���8�خ���A�u�o2/��YW���-ge�=���}4_�r���B��Sꃦ�^��2�%�5coj&�\�Z�z��@�Y�۶���q��B�!2�%�O�{ա��Uo�uI�ڲPp�hQu��0�=�r�u����P���)6��C��6:q�5K�f%>�S��*ײ�/v�� o�ﶯ�+H��c�y�� 1��ב�P@����%�Xg��S)�	U2�#Smz�V0���3Yʦom)ۧ�3�����!��󮧕�C(��mf��v<,%��B:$�aa*����d��Є�-���;3���jL�� �cz��XU)|L(��^�0��e!��n�P0��bx��;��i����3�����A�W7�����K����_��v��+>�	ۖ6�b�M�=y�S£��7o����1�b�V^�z�fs���7���WW���{��}y]���V��N�4�p�f�;�S�!����Յ�G�Ѣ9� �j�2 s�ٹ�Z�١ڎHA�|�]8j�|0*��G"�����q�X�����MVo�%����~����9�˕�9p����������+J(��׽��z˥ךf;�<y�j���U���M�Ny�ϭ�@�������]����gZ�З�`��'UȌzO�3m��T�j�	e��Ke�N�c�
:Ҟi[�δ�,�b�����1�`hgޖ�r�v�K{e��QQz�Н6	y`5�ѝ4�1Bl��օG+��"�5�C�\�$,uZ�ջ�Bf�6�!-��_��{�R��^�l/C���OO��k�s��Mz��@�ԫ��2��=ګzZא�R�倡��$�L�1k	u����f,oEotᕿ�|j���ǝ��q^�%����ڠ���W.��^��b��L�ha]�i����œ;�F�Te�<�f���؃s���������^R��8-x8�G0��$k�?�uBX�ɯƓߔ4��L�a�Q,k�<�sM[՛�r����s]��Y2$PC*�,��hƤO��ڥ�N�)w}c{�3�Y�����A|�h�B~��*?~�+�R-1.0��,�ۓ��s���N׆�S��򋈈�c����������]@׺�z�,:��\>���H�~�jbY5�K�0<6��3�N�H;�ho(E��;�Q����;�oN���_���c؍<�s���v*JIެi��SE7������f���L�Ȱ�Ḣ��]�5
�C{��bQhd���A����;
ۡܒ�+���{9���z���n�V�2��$�8x��BO9� 1"��=z����������B��9��`w���|$;���P���Ic�/��_�-�@�'���%X�����ѳ�/���m������a��]T@�1Gύr�D��h��*����S�f��><+��P���� L)~0/�VMt�i����C��3�0w�������0��g �iʆ�g��\��[ʙ�*|��ږ�k�L_��yE�y*���\��c�(�7\N�m%����3˶��F��l��K�-�2nj/#Xt�Lk0b�
no�q��ɼ��[d`Q�k?�;�w��UE&��Pj�O�&lq���[���	�{P%����=w)�`�)̏fƫ0�[�f�f������~���;k å��������6kԼ�E干�M6g�Aa�`g׎kD��͐�glsL�Z���Q��ᡙ�e�d��-A�y0~��P�W�t�i���>�ekN��]���������qKR��s�F�n���\�[<�͇���A�H���'�v��&�f�\ݵ����EH)�,{�wA��vy��=y��!�e���2$�ӝ�U���������Q-���EPܑ��j������/���J�32�.v8~Ӧ����y���w�剧��"�m��;i�W�+��ѥuq4���$���8���y�q7wQ]�˫jugf�i_ UnN:zՂ��-�|�������g�� �J)J�R�_???_��ן~w������o��5��z���t[ex��	���i*�~@ݡk����٣D��zh�����.�Gf�p��lD<=7j�az����O����ى��i�/qX�_�d�_����K��x~yJ(s�(�O^��qmWp6�;c�~�n.��|�k����ó�g��7��"����u�$T0�c��JW�q��D�`��x�N4/Dy �R����շ��RL�Y3��4dDtC m��M�9]-YUk&~Ƒ}�������_/�q����z�y���, ��<�l����ş�b�9�=�Oׅm�Ot�pZʆ������k2�K] ��*���Y<{��� r�T�y��lt�N��M�;�y���J�G+���|o;S	|U������S^�_D!�Q�a��3^�4P�6<�c�O�<��I�d\��4y��#�6a���B �M^��\1EL�]B��%�k;`c{��d�v��L7�o9jV�ku-�`k�ܼ=ݝX/���N"%��Q�جTxOͮ��j�)��1���W�b���a�E=�KFn�vt��t�ڽ���'"�+�[o�8�=���M�9]�u�k�^̭�O%���k_]�^��T�������Y�T���_<f�bt��؉M�3�����je�%�fWD�Xd�sˆR٬�ݫ�T�]�O�'���1��(��`�{��xU"{Q�M�x���܌�J��k� 63w���5=���c�S���v�o��,�����E?��61=���XJK	Z�:��ڼ^�	C���f����jc�mgj}k0t����I�Nxhm��7��+�|zp6�/��K�h�����(o�G{�L>����_fS���nͷȲ��	����\���,㋿�{�7�k�|�_z*@��usm��f���ܺ�f�t!ڝ�lC3��i����
�`W@��Z��o?w@�l���4)�ݚG�Y�|�Yt\3���t�pm�oF��7LzU!1n��U�a�Wh�g�tUf�����b�1���ǽ�΍��g�iF)�����׀���j}a��Ț���j�N�m���-��-�i�sjg��̋�;E�`ޥW�o��E׽p��M���������fy�3z(ʛ��Y Z��R	O�bZ'���ebM�y��[H�b��j�.S&Y�����v2���?�W��(q-Sp0����잚��{�ʽ��X��a^+�շ�<��Lv�ѕW|��P���Z�����|o[}A�b҉k� �N���v�4ڗǮ��S���<��U^̔s��sN��R�2��c��M|L-��w#g�xk+X�g0ʒ�8;Ӿ�{�Sv^)zNl���
�����*����5���k7ŧ;���`��:-M���m��+Z5�"f���W�B]��{lf��*
ވ�o�L���#T�( .�>V:����S�%%���Ɓ�oe�����ª|�	eE�b���W�5[�hgc�6'��۽˭K��ej�|9�0�ܱF��_g(d�,�xC�՘@�s�a����j�I��_M��{{���Y��L��l�v��X���R�9Av��(�.Y�����A,�7C6Ķ��溕ܓl���"���5��@���A��Z|�պ�Z:̇XLJ�u�2Z���$cg���kV�AA�_X0�OS��7���Z�nfUE/���Y���4�12�֚�q��"��Kn�wp�i*��S����=åv
�V.%�w_R�A��g�a�ӺmK4���:p�Q�������+*.}Ը7���e�F[��C���J'���$����S�gZPVԔ���}F��0ry���9**W���{���{�^)C��G�Ut2"#-�(�P��Ak�.�[M@@���ls{�ϴ�7�7B��j��l!�O&�V��n��銿�Mă�M�*������(�++ >)�/ba�+���J� :)%Ɛ���̑���hT�X��h6�N��,1�խ�3� q3C	�ϵZT��Pb�dyЉ�s�CQs}�۬Yl!�:��2��T�m�
+�ں�lw�3J�\���-�{��+j+mr<�3�r[uô8ը"3)�W]5K�윮%(_d5׋v��3��7@�Xk���Uō:��+�1>�t�����b����9�6v���i��S`p���sGɺ���u�ȕt�*�ۮ�,F�Z: &Dգ���� jj��oi�@V,�o]7�(�![��MҮNl�%�ġkU����R�[&��0��F���q�Vk���nb�qf9/��.ȧ�$��8x�dڀ�6ι����Z�.�ż$ͨ[!�*y�u/ϩ뇆M�k��\=��֦���}-\,:���`/2�������qxފ����S:5챋�q�'L��y������Rn�!|�����l�4�'	�a�E��.��C���z�8�l�]��M����R=���S�d��_i��Kz�:BR\�o�ĕovgmYȗS�s�g]h;�N���}k_F4���,P;��k���sh�Oq���k���u��,�n�T�a˺�t(�&k�uo�:M������8�w+��j�E�ZJ 
?��G��P�(фl�BN�2!B�k��B��ņ� *A) bT�&4�Ȍ�(�*�L
���)�H�%J�Bͼ��d��1E�)��.�b���<<��4LSEP�Mv1P��h���^mE�%P%;��Q5G�9����}�t铧N�.t�ӧN�:t�ӧL0||�ɪfh��h	��)��TR4|�W�5�m�E�4A�EW��Ǐ�����~�>0t�ӥΝ:t��GN�(���L�߿�X�!������r�UDESUT��ljf
B����DW �G�Z�D�G6Z(nX��I���i)h(�
���,L�Q���a���Dy��I��͂�H�b<�PLT�4^cCTFƖ��*�#MPp$14�.p�T1U'3���[�EQ5�Z�&*
*(�����i���<��.�� �J�hB������4QK3L@�z <�)h�����f��`������%4r3D��AQ>X)��K�o#EA^l�%�^X
"+C�2 �"��"�&�QD���T�Er�/}�ˑ����w��=s�5��*fhtb1��e�2��gkqJ; ���Re|�z'1qhRmr�h�r��V���gwf+�ԡ�H%��7�Ó�.��o6��RO���O9�$@���|v�,�rG;�YTi��c~�$�,;�[;w=_��꿶��r�z!2:�eν�����������Z͜ᐥ�c2`P��9�&�Í7#(D������Pg�L�m�=�JO�`�¹�5O2K�E���y���;�
�V�V@�m���6B�A�;K"��0T�͕n9��`/k.X� ��6H��r�f�q;�9�f�nr��J��|k&9���K���rC�B2+d3�����F5����7�6&ꮊ����̱Z���Ә�����zuب6��S���uVy�'�lP.�b��G�s��[��I��P�DG27S,��CX���C���n[�|ڱ�=B�Ӳ�MSC�6�{�ܱ�t�����D!a�ّ>�^���-YL!�O�B7���Bl��փ^9^v�cY�Sچ�N��glf���lg! ��c)���I��ͅ@�<�������i��n�y����ά�pb���̞�vu͡����L��c���&�
?��61�R6��؞5׊�vgU�Ő1��D����7��J�!N�"3Ӑ�}� �1x 4��*{i��h��|aW3*��D�W�T���y�c*��"˧�͜`�X��s���>�Y���P|���JZ�]���_����~�S2��A3���Dj=�L/���f>�b|y�YQU⩳'^60q\;���*��l��T��=����'����0����,���S�*�
�Fk8M��@�#�;�\��� y�7���<�,|�s����L�ck	�n�� 4�7T�Ƚ0�*����L��vmK�aijh�ANDL.�=��s���0u�j9��i-��l�LN!��Q>�O3j��������NӚ�^���Ώ�^�㨻@8?,��ʛ1S��F��GTh��Э�ِ��f%�e�9��Ų߮�l�7���������爡�B(��p��Hw�qT�&�Ydk��`�
q�ѩ+5k���*(�^�E*�|la�*��u4{=f��"}nC)��^D�J4��`�['�;�������X 1t�p_�ְw?7�B�\����mk;��<�v=R��Tya{.��N��\��g�t����3E���5��#^S�m$�`-c��ˑm#�g&�0u�-�<��L��\�{-~�c?�>>_��/��H�oTחA��y�P���e�<Y�{*]�;k'C��>0��a�
g�~��I�Qz�g���q�EfL�Mi%�RT;���=od!D+��c=�s�i�]�WD�ӝd����,��gÞ�0 �+���{������*������1���
5�n�ݐeM#cA�����5jG>��^�C��ќ��=�u���"�ֺ��D�v36-�e��6��D4Hn>(�b��ha���w��������~����?ÿ�yo��ք ��e�A=j�Q�w�#�9�w�%����<d{k.�_���~s�"�·.�]g�A�{hf�܈�f�p����B���&����U���&�8N��,��-=C�@�38�����y6Z��6K)��
g�s�P�X��Ý�	��ß[>�`�;K���i�}���LP���f�A�|����U�����˻��@J �+<y���������-Wo���G��-=�Z���F��jΖT��'�~���=��~x)��q{M��`�Xכ�cn}� �e�e�ōp�SU�{�k��d5M��_�B�1
�J��{��5b�U�R�`wM�~��v��|�:�l��q[��8��ʘ�L&��`Wz"�L);/M,����ЦZ���>�S�Y���c־y:�j�V^���1d�>�M�C*j�$� � �P}xi��}n��E)���[׮���@ډֶ����׬� la��]��S���,,wF��l�{oLn.Z_)��XlHd����8��v�Ժ:�f]\��\qA�Ukb:�vcΙ.�`�iUqu��:rykS����u�pr��}���=z�h��^�V��ܐ��M3/8����ut�f��zd�G9ا��{?������<'�J������� .0���2�jD�gc�>�:f�ɫXGH�=2S�Q�6��6����W&\�]u�M��ڨU|;����D�Q�.��dۏ1fs^p������>L�*�=K�9�BS�I� �y�G=N��m��}�) AE��V����ku/#C��������`�^�t��߷�0����=��{���g]�#S���{��%����K��;C��)֖���1\�p��Hǒ��"��=4vf��9�7�pM.����𴌺f�3�=6�6;�
fН��6�b�a�	��Y���7�'�c/J�F�V���l�zJ;�',7��1�S6l�kh�c^h�L��w;�cӠ.�p���)��oN"��,ӑ`�i�Mi%�����e�7Qb�N����ӵ*���]���2z�,DZ��w��<6�y�
q@�Jl��}y�r53ܪf͊�̸��lC�ҏ�3]�t��9��s��쒍�� M�A����m
6��ʞ=��4p�����#�E����}�G�A��D��=�I���g�8�r�i�;U$�P=�~����h኱��D�v���0�֎P����)��3״8(�NBʂ���0Ф�ݐ��6�Jt{;�G�
Yy)��p�"�D� P�T(��k��U8N������"��Y�I��];�C���g@��n�t��d��q�U8,��R�-���v��FnŭG�J�܁N�LR5s�<����O\���𦤒��y�W����������[�,aSlG������"[h6Aa0�l
��Yȁ]�/`�Rl+��R����>W�R͏��/<�T9w;���#]��.uX�n{��{��{����u9^���x`Ze�wO���ަ2*,�z��q\�<����i��`X^�:;۰��z�ՇF��V3?.���ɍ���Y�e��c���]P�=G4k=�Y/�/-�]�>H���&B蚁��{ŁN:5�f���Ʃ���̭�e
k���ù<z�QjC^���!�C7y�q��k`���K%���*L�Lt>����1k˭�j����[ӊy���R6�٧q�Y.+[i�iM�T��O�|D��1�z{��S]���]��(:g��3���b��$���+_��4h=��G�LB}kLq�mj�[w.�pz�fZ�L`��ͫ��n�9�l�WL����V�è,y���TcsP+RX���M�&0C�w;�n:�t#�%b�?��FƵ~��~��G��������|m�{/���G��إ.�yu
	#���P�ή"e�D��-�j�['6Xޭ������C�[M�����DǺ����e�8&Ui?xT��AN��o�1�2��ὧ���6[�nX]����9�	=��0t���<Y���7K��+�^ ��)�=���?�x�9�@EUS)5���W����h��@������xh�L�j)��4��/uT�����J�r�P���%w�+�������!�"��C�(`Dղ}2X�O^�����I��dCN?'��c$��.�R���}�^�ZrDeU���'c����P!�υDs��O��Y�1��1�ݪa��v��b ��Ľ�;��g��^J�!OR#=(��~e��An�	Ն�i���9�f��'f]"�/��f	�q!5��Se�z �v�C�N<����6�Zj9I>�d+#�DLc���-9��jD�Tˌ3l<��=�NH�}a=����_���3�� ��@��*��G����5�
�M��	O�L2x&;��?�[_3xK�Ʃ�]��%�!�."'�qp�Bݙ�M��\
k��8�e�X��� �-;T;vZ�Z��K	�6��NM�nm\r��GhUS��^~`ڣ}���'�&G8�C%�36^�l�w��3Z[�P����n���O�nE6�oXT�C^;�������y�âJ�Z�@�n�֤�=�Geiᣯ�Wӳ.p��,�^�����a0=�V۫��@0�:J�9��GWo�� Eg2�kvl���λH�\*o|Ҵ��o��+v+�l��4[�n�po;:�kl6��[y[1b� �Å� b�� ; C0z�s;���{o�9��i���c�P��)���cw,�ǡ�sS��k��R���^��(��<C'ڸL�}!�
},��ސȟNDGz�wh+l���6�H�}�N��D0z��S���Y����<�=HB.476m��d�u��>�D�T�r�B]3��<���3�Ʀ�v�j�(qn���5=���x<�.��d��ӈkѼ�;.Q�^��o�3�X�Rk2s�3+,hǼ�|r���-� �
k�l+�=Iz�J�]�sce<T#|Q���\)M�sfX\x��p������G���imp�aTs{
��� vKU�l����]�z]FDzyO'd��s?o��;���"��Ţ�|H��m0W��ٷ!�W?)��%
F�y��
�Iw� �,:��8�¼b��~fmݠ�%�WSl�
Ǿ��7�r�ms���CH�^���f�vkNtdy��hn/��a1S���:�"��u�A[��K�y����V�s󤼰U���ߍ��H�Q��N(�b��r��iښ����p�g� E
m�ђnPre��	]p}� |�	�k�l�N�����&��*�Uﵛ;+�ެ�,zzG^��Im�*���i��U�}ڲ�X���W5�T$LM3D92�8�(����R�lT��Z�e^uۥ����ٍ�]�uL;
�[9[=M��2Q(��v bE�7/��ʜ�k��v���?�TT0o<���1�Q�X!1N��~[]�τ�V��o�'"��B�W��ը��׃T��������ɞ�����>&ƥ�w�{o�J���{����V�Rl��/�b����2��0X�&�Vj����Ɉy�m�{k���Ϙ�_ZEi�3�Ӓ�OV˛k����q��Y�Ly�a�O׋+�h9�.�mC�vսh��t���X�l.o#PZD:.%9f�Jq���c�oD$���ˍ��8�l��Y�'`���1-����LΊ]0��䄴f�K:�޽����`3@�R����0}n��GbId]>R�'7NuV/J���p���O��P�xV���{�ZyE\�B�?0j��,��V.����s����]sn�>���R�y�@��dK�l�0o=y/%�8�n���γo�>��C[K��3�;�9����N�������!ϛ�̣Xÿ8�����V�6�F�Fr�|B���F�����t�Ln���n�R���0��Bd0�I.�l�)��6G�:�U�QQ�4	F�sf^A8���{xM�Il�]�ϻ0uJP	�S\X���M�U�췟`6]�:��3l�����QǊC�չb����غ�����������c�̶[o77c+��&Y����Ҽ�������
��D�[(�L.�	��������9�^@�)[ϑ_n4{���b��)31f�0�K�R��1x��yc1�[ӄ�d�FE�� ��6��1�`rj�w[{�[;o/�`�D<h�C�(L$�}q,�K:ͪ��;�3ͳ���Y��HOb�;O�vt�v�9p8�wXΔ�p���^e3�aa��-N4�;�k������gi��ԷX=x> +�n�������N�ג�����i�S��I�K'����ݼ/uBc%�+ww����&d-Eֿ\Bc�@��Q�`�ql��]�����E@���[��]#��{7fgA�8۸�VAgi��\DՓp����$töm�l�O�6N�3mŖ�T��������/�fj�TPc,��p�M�2"jD��i��3.ׁ�"v�%���x.w�f��^P�m�0��@�9��d�%�{�,^��$���̤��:c�oPb�v�gK���o�-�i�@��� �K&��}f��3E-�k�	�L��&м�Yv�Krun�l֝c΁ymF��)��[<�"�a�v]�64T��+&��ԫ�<Vd��p6)�Vs��*í���@�=wO�9:`��AVuAJ��N���܈���X�7��r)y)#H�0R��|~�Y׽'M\1iU��hq���]}���3�^�ʘ]��@{-��!li�0�Z�2#n!t�"ml+u||l��r� K�3i�^v��{1?���w�X½�s�}���ZVQ؋k�/^Bڠ��M���M��LH�ОM�6��g=r�t-�[!�T�8��<^��}d��ǈR��*�o@�<EE����v9ל�{�&�C�+��m��M��z�2#A*�=��e���5��q8��^=��e�kUOry������b(�z�
�[6�,W@����֡hvs��}m�tA�2�cy��V�W{�՛�YМm�΁�̠�!���
Jxh�T&�yji���F�M��օT,o1陭�*'3;Wf�I��"�,��[��P�aؕ0������-����5�<�:4+n؄Qؖ}fSɞ����;J�)"pW1^��_A�+��>[фxJ��0��U,��Dg�����D����Ħ�����}�e��)�l1�b8�%���36^�ɧt�Q"z|P��D_��8�O��Ϸ.�j2���X�f�9��9Cl3��7C��:��z���Ж�<�3t�rGEN����am̓-�&zǆ�<�<=�9pcT
Lʷ�#9��oCIB�G��D�m짙TXd*B��u<���E�{
����d�zQ��u��gjO�6;�2�j��k�|V�jt	�ל]�����<��pZ)�E2#�A��H�U�s ���#��ڌJ�3�fJ����+��e��'���{��v�"�t�����r��~Xw��� ^�q���f�o4h�ع�0i�w�}���f�������XR,d��*G Vd�+GW[�c.���a�S���v�����	Φy�k.֌R��Dk�+t�l�v�d����U�R�!n���:���_.���R\�v�j��-Є�������J��:��h��b����D>��;;�7�ǵ�AՇ։b���u��s�A�Jl�u˞�ߟe��5�mqՌbT@�����V�j��$P>��h�w��1a�� �[J��3>rA���j����|G-���$����cn�u=�W	)]6��N�3���b�Wy痌�y�%Q��v��@[+3������;�H�O���7g�ՙ�p�dWr����u��e�9�'`�&I�^�{���Ž�|�Oh\�**�"�A�
�h�]�D��l�p����{vV��|l��'��']�J��EL�%���T#��ٓbá�*`m�wJvB__Y�-w:�MN�B�ŀ�DȝaP���{�L�H�z���D��[�Η�� �G!RF/��0�����V����f�t�J��Z�4��H�1P���T0W�RL��3�`�N��Z2`|%���f�@���|�ǍǓ���lɥiU�0�c{�*KC��5���v�̝6�Tp��k�zZʃ`�~t��xk&��Ȩu�Ei��wo$��Zs.�N�m<B���rY�Ejٜ{'�a�\��՗ki桯k��6�l�s���'��zl��#y�E+f[+V37;�ŀ��M"�Ĥ�xw<����+�9��!d�v�������J�2���+�L�����H��[@Bk0k����9l	b���F�Ra���,Y�`�Vɻ�]+��Hل:gj�d́ʺ��4�S�y���ݣ�%�i	`	��	#|5��n��κ7]�|��h��Ew�z���f㊹H~C��wيc�	.�W;�2':�8H�]>�V�z2�r�]�޸�,�Ui��μ$p�e	CM��%��v�Ș f��p���L4@�`�"U��a��襢��x�������R�X��H��ka�����l��,eqnVlI���:���Q�n��� z/Fc���g=����,,u��ͅr�l�ao-���y�Te�3�1jp�����w�{�� Ю�����[��=΀wl&���k�V����뇲����T�wb�����B������CTT�UST��LPP�x�s����������ׯ^=z��ׯ��^���������~����jZ�(��F&�$���(�:NlAO6b((��*��?\���~������|z��ׯ�^�z����ׯ�>?�������}�LIT�KE%PUUCKT�S5|�U�E0L�&"�bh��0�H�i� ���$�����IK-!0�EE�T,LA1IC��kCͨ�J(�)��%���()9[�D�AE-,EQCII\@�'"�墋��QEEU\��4�R�4$K�3DUAU$J��REI��dĦ�XH�LKBsh��(�hH���d�ѡ� �$�4�PU�Z�4�QDM�I��g%PQI��p ��U!M!T�QDlm��P��QD�s�k��a	Έ�3"���rJڰX�y�־}ʼ�3b�b�+���͹ԙ��4�D�(�!�Z��cc�����3fAN#R���<�Ĺ�2�i�sB��O)L��7�|��x,�:��_eO.k�cr� �^��Z�V�6���i��I�4}ў��)�u'g�2���޽�ά����݆i��*#|��hWy���X�W�ɓb��n��jO������b��
����,6����-E�b�O��R)�}�9��s�&y���"Ʒ�-L��Zy�zN�]q���vc;4�t&�u�_A��}����Ef�U�5���ki�\O�T���gQfS=ʘ r���,\�Af�fC4e#Z��㑂Ҟ�R5�?��bVm�F3��;�Z��]Me4[�+֡�[i;sA��M�zF�\���������~J.��i�ݪ�MY�r8����V�A[hm�˵D.ol��:��|��#�y�wX�vS�;MC.n���V�[\���y����㭞Z��d��XF3y�B���/-�U%��0y�Q��,����ht-#%�P�k��X;nM��4�T�`Mk�3I��7/7���G�r�{��6O�
���{��zOr�`��f�%s��+hd��{ω���u8y�������P@<���� ��]q6
���ݍM����ڒ�Öyv�GY�o�Aw@�r�7�88�r1E$ͭ}��gEuܵa��z�8�4P ���Y�":=����\C�O��^}7`�d�j9�#k�h}�a{�W^"��\>�r��.��ݡ�k:l:�p���y�C�uB��⑭���
�o@��@̖b�&9��h�9�`�q3�z⭁d��wd�1�8lOn�8�\�77�3Kl�;�TYz���kr%<q�L��v���=��zXΗ�7'ί�<�8
�yY��e�8���A��6����e�Ț����/l�tG�uC�mQ0�>{2$FBOR�n)���ޛ��$'v��ѫ;w6���2�~j���������ߔT8�0��=��*EP��q�l�z�el�� nث��=��ד����E�a�1�n�e�aM��!��T�m3�_0�������&r%�¹G�<4�=�&�k����
�\������\���J�\f�v=,9����Uv��l�(ea����C�q>I�&i��bٱ�7��I�)O�7�V/]��E�U��Ț���Î���M+HK5'-#8�5t˲����|}����g1����csD��~_��7��WI�lDZ�8�0��U"�~}��wnX�1�K�uf�F��h�.���Jr�fҮ�ZFL_]��3�B3n�lL��<���vv��C8�XN���r+�j��E��|7/-y�s��~���z��p�%F�,5E����o�0	ҷ���hC�/l,u�u7�LЗ�0���i6�B�ޥ$r��y@uQ1�G�&a������ה��	��_���k����ւ�����;2-��x�+hK�l�G��R)��ufv'HÏ���%��
/��x�U�0[�g�H[}nf�������*��}��Т,���^��?<��zR��5y�A4*�����61=���ZRXL���f���Of5���1�+�a��2�R��S��D)d���T�$�F=m��<іMh���jɊ������Q�p٨<ht�<�@	���}W4Ŧc6?'�Z�9u�4�31;�w)]b�u��ߚ�o<�,�m䙱7s�j�q�������<��]y�5�9�vF�ξΫC��܎����I�-F.ZAxg�4"=��ȉ���)�)�c�
��܎��w7/<������\CKM>p���1�#<�iS�AN��9��	�9t�F��z��.�<�O�=ɨC�-� �������4�i��~^���AH�E��a0�Ʉ�y��ZB2��uu��+�\�Պ����ۇ�N돼�ՙ.㦆P���3sܰ;�E]N͢��]��MS퉢�$d�m���H(r�Kn.�I)ի���\�0���}�.jL��E�s���x̦���<(�>1r�C�+�u��M�m�455�t�}.-��"��Y^�C���	�r�^k�l`���H��-�	�D��u^�-\�M���Vt[Ht!�q��6�R��ƨb�^^u�@�n�ټZ#oߜ;?7����g0~�}�~/n��������k���XT�q�����g3��Md�n�
��t�6��u��N0�����(^C��w4�ǚ�	��q�7aI�4+���s�ֳou��Ja����$�a~�[�MД�m-�m&1�L<��tdxg���o{do�*�F�%�ϛȿ0V�\^��<��<�ߧ���ڞ=ϥA��WJC��Pc-�Kv9����d>T�{ٻ�`��&A.:c!��)�d��xc4���|M�Ur{��\�����o,w�zk�V��$"�=��2^Z[��� �?3�;��M!���5��j;HR�'��Q�v���������8�\��y��G��g�C7c�/ϾRaF�i0��� {4�/������)���gEZ��z�5��|����T�`�ؐ��l�W��+�~N��r�����~��Ӻ+ᨯh�-a���@\��� +�o챞*��Ybub��,����r�P�V��01|1
����-{�Cݴ';�+F<�U�ri�7��(fVu�Ve`��pǨ�S��'|�gj8�[6�+��p�1��O�� ?��7��f7{�HQ�X��:�/��'���v�8��>[фv�J�#
$�0c�&_3��� �%/w��f�N�w�hXui�O��(1�5���9=T�&"�C	톞�f��z�dR��hA���ho�7��z}c��׀Z{��o�W�.`��U���9Q2�:�p�D[y'f1��;@��ȩ�{i�s��N�,���[�2�1��n;��j� z�3��rve�G; �Uԉ؁�ͼ��i�/o�-��󔘗3&Y��t��Or%�&�.�hK�3zL^��٥������K�.�\��-�]W�:�J�ͤF��.�P�-�s.խ���]sہ�^�te-~O�ҹ��+hUZ����q�tf��6��\Tմn������cZ;9��Al:��׆�<��)?X�"�h��{�T�8�y˃�^{ٔ+%k�K�֦0�Eϝ�yaV����K�[�b�{@,oV0֮Y9/��^��>��\�^�F#����J}�
X��G ��C6%���A/I�o�P�oz�:Wv~�	����0�f�=�I���ۚ��mk<P�  Ӄ{	�3�T:h=Ѣ�+j��}�ݽ{�� ��H��hl��q@4f���5��C���ܴ������nu]�(�K)!�Q���tb���&��6��p�(�A�a�sb'i�`φ>\�m��톌a��R��dS��]��7�D�T�rI�-�����ӧnyx�B���z=r1��wV�z��'�R!si��I�3�9�F�:�dF��n����ń%);2��oT���X��[wX^��cE6W�1�;`i�L(�z�]Rڟ�8\j�ܦ�����AQ"��\�x���׎h�ze��F��͋p��2k��dܪ���ݲr�K�&1�ң.t�����8�'hcWgH��U������ʺ͒��D�ʹ����-y�-�H��5��yLt,�5�{��ϻ��8�y�s��a`Y�V85k��VF��.9�q�.�2S��㐳
C֧��N�M�"�L�Mx�|��k�bT�y�]����,2�s�C�-�z�lT<��~q �6�¶�Wa���w�τR�*t��;]�N-k{� Ts1z!� �}���tϊUz���r�U�-�d(off�j��r).�h�}d���ق��� gE���]Am�wu�-���)�G.��09(k���
�L��Fn����f+�-۹�
�u)(���%�zf���3qFr}e���w�H���_�Qމ���t�@U���0	���C�*k:��f���:�[��T�|-�UZ�[%N���xy:��ZT��Y�fV>p���P�YE�*�E�&�� Oɺ��(E�!CP�ȋ�t�nl��
��ة����PO��P�]_?����W��T�	mLC������g[a�kN���S:���KH� �/�;Y�Ke�c�g�~�YM��*s^̨wT�8[�nf�Ƨ0�x.�e��y����E�',�ju���>��O�
�.;�F��\^%��_�t�e
"�ju�]Ĵ��R���[i�_l/�3G�A�����;�uv��oMd��C�Sio?`J}^������̘��.����c`mu�骋Y��#.���yu�Ƽν����¼��[��Ԧ���E��Z��Q�"2�ŀ�z^tWgC���jVf���=(Ce:,�-)_��iN�2y���~�*�N#V����<ާ{��
9����w~�ї9]�GT�qG6a=���XJK	�ֹּ��6�Z6H���;_�7wnA��#��,��8��	���򸇮R!Cj��6���ag��@�3�슚���]�y��
��M���6� ~2|�M�� �-k�<75�׶k[���!V.D�A�8�U��#��[]{�-���!K=�_N{�
.m��V;/.B�a����Mz������
�',F�5ŭ/$v1Ch����s���u��M@.CsR�iR�L��N���o+�������m7�g$z[�3)5a_G���΀�ۦ���eEG�j���\���m��F�P 4&��3aw>w�U"Dlaz�d��l?{CE6�wT�t���E���L���㙳��b�����@��`EJ�.8A��i|�/����d���Lǘ=S�p)o+lK��/*m�O���'�Tƽxl��} ѽw1/�s�Gun�nd�;Vt&��E�r�[�v�Q���#'L۸y�{ۑu��lc�����V�.p������2�1ie	=a ��ű��a�fҚj��ʉ���t�b���-8�+��X��F�&�ذϼ�H9U�]����~t�7��[��Cp��Wv�B�[ݮ��G��" eE�
���ב̱w���H�Bf�P��n�Mma�R�DsX���X����ݬҲ��B�	sze6�j���)��YX����1�3D+�w*�n�[�O7;�Xܤ�]hn;��e���S	�x%V�V�W�*�}j8���=�w6���"�йw6T�� �!6W�^;�f���I����Q������b~n�T�}kT��!��\��C�֍�R"�,��3�ú���Ո�����ᚂ��wNnkS�E�����<4eY�n�62�܅{�J�oX��Ĥ\wM��Õ����Awʻ���{`4�bM���K�Ws�
^�����m���*��UP� �(�Q@�@�������EW�h�LA}<����-�Ҟog#"	S���a˘��{��P�̚r�2��b���>;��2Yθ5.��LG6m��2֯�C7k�(�9s���!Lm/��Ke�nѪ�kЃ�q��Cr`5��EK	�!G��Ϲ~�p�_�u+�U@P�3�fo0`޼Vw���E�x�g��7>"{�����n�q0i5�(PW[:,1��6s���!�팧U��y�r��Y�3x.�P�sH����t�0��s�l��G}0ε��Nm;'XEܽ�~�x�%��&�Ň��Վ`)	=c�)dl����6#��K���͗�a���b��K�r��/+��Z���w�66A2�}n�sE����Yk^�^׀ZF��c9?�����
nevcn������yw֟D'��p������y>�w�|�#Tg�u,�bvsG+Yf��m���-����<�c�*9�Zf�E0y�b�S+[ʍ���P5��(ϸ�Pb[���v�Z�����T�7�y;VuBa�����R�).���~P&Ew5��l� CФB���%If`~�m�\�ɝ�M�:��䡴GW�W1��'Z�P-�KY�H��o��s.A/�[�n�푶:
�e'S�7%��nM;#����=�Be�9b1���4gs;�7� �F����%�Z�o
Q?�#ów�ٕނ>�����F�MVbY6Z+n۰-�mM��Vנ:1A�+ϔ�%y���5<ݔ�y������W8�8n(�⍵N�y����7�ڬ�5��*���&�w���sc�z��;��~�oC�r-�r`Shi/l;/�bj���	���+dR�`}���2 �.���N�T��veS����{Q�eL���^v�)���3��keN������Ǔ�I���>Z�oN��r��r;aA���%�ih�*=K����xd���k� �6Q&�=;U�ѫ�1�s�e�̺�[4vð�wlaM���x\�%�`�^Ȓ�L^�h��jl�(s׏([!h�O>��,��2X�1�X�M����>��g�k�nc8F#u��Bxu�F�iЧMh���<�;#Z���g�NC����u���?{����X�Y���P�2�
��\b��b��H��)�^qg��^9�#h�kH��A}����X�e��W���ln��ƥ��)*C�@�ԶM9�_C�H	�;��^���P�"V�up�+��(�u�Xx����\�j�T��ޚ�L%��T�l']P�C�_9�yɲ��[�y����B���;n�[;�p�bH�}+��`�u�`��7 ��_ii�|�L�'n�k�meZ}�\�m뚸&^p�&��f��ٗm�,>�:��8�Ï.���b��yi4i�xȏc8�@�q�-�+�;�S��?�L��2�XvN�e�������y�,5�ɂ�]c��Ӓ�ạ�.�!��ܻc��bB�R:k:�u8�v*n8�7�k,��ޖ�}˥�z*� �,ۂ�WT�X�D��}��7S[�u:�<�t�z�o-!YNlR%��PXn���םo�^�{Z
�yИ�N��eu]�I��e��Y�fH5ΰN5���5���2�M;IroP�R)I�wj��(��B��lD;.����\=JB8���5��������>��K�`��]ѽ!��N�Rx�n���``�Q3�5Y���M��f�:������u�w�u�:�8��UҮ].M�ә��{�u�}v���!�e7,���;=)���{uj_S4T��*
�{�SBKm��uv��(=�BXK�	�0�!y���<%�KV>�x��\r�jۭr��Z���w�����K�a�B3��Z�Z����uQ�2�7�/:v�pJ�Fp�9����۪�.�b�b�>٦�����}.X�)�*� �WX6f�i��E��k��&T�t�k��GP�h
�! "�Q0QK-�@�R��U�"
�����ZS4	�4��@>���^�"`����c�σ�;e�����n6���w�4�(n6F.HM�3uBҮ�H�2�Q��:*]�c�^w}ܳ��j��'8*Z�äm+ɢ��q�=���īH�-"{��-�e��j��2nuf'[r�ymk��|❝/>箑��1ok�zc�a���]�n,�K�T�[PUu��1����ү{�>�ձ08U�5&�;)�.&�kV��{�����Ĳ��x_ʦ����� ��6�;8�����e��5Ŏn������3�.�<w}�������g:��U���F�q��c.��G�\n���ѯio| �,�2b���[[I)�ܹ���;�{�Z�{YJ��1uW�(�+��??aly�N���;l��GqZxv���n�!Qs�M��[Ӗ �o���8�<W���W��讝{+w����҃t&o�uı\�nL3�ՠ��:�d��h8Ѭ�X��f���B�Uݸ�~�����-i:�MX�Y%M[6�^�I�\9��|5򗢵��2n�ISSp�V㰺Q^�],��°�{	l1q%c0(�)m_s�W0<�Q�ר�@��t�ݺ�=�) �Cڅ�30�ٶ��HrC6�t��Qn�]�
����3���FZn� CT�E67Z��*��5mA!>�hJ�:�V�TS�R Bp�s�I���_aH��D�a��6�dǢ��� SdQT�a��Rj�u��h�5\��p�����������R��4�44S�~9�����GN�:t�Ӧ�:t铧N�.t����>?�χ�P�"
�b�h���2�y�#�ı͵�
8\��'8||\�ӧN�2t�ӯ�^�z��������?��AT����D3ACTD�Q4��ICAb\A$M�0ELJD%���T1P�P�BTIK_-D�q%L�MMDL�5ET�UHRD�T���Fى-�QIUA@PE��$�"���b��`*��h�����98���*"9�	�X )*�I*������"%�i��h�*R���xLUAC��M^����sT��AEy(h���y'��lW->l-M$E��AHQ2Qlꂚ�	�
�\�QIG6Z))4���|�CW���9��m����[�8����'S������̇��f��ٔ��q�퉨^eN�+_H�kwQ͜w��9E���9Ż�u��MW+��8\��眱�<�g�9�����?"��Z���]�)�@���Z5�)Ma�xG_#��_N��?;@X�V����{4շo�b��K��;�����Al"��<�꧁�����D��0�l��R{����cl��z�*�=���Ǟ��3$�^{��P���@�O~Z����/~T�ߺ���K�3��j��uh+�[=K�$�&r���ܩ�������.��M��rg�j�����>}S0$ғO|�q�w��5^U{9l?[k��V�f�y^�4��8���UP��};�W_���x�n��O*��t��˲:"�m�y�3-vӮ���>�+j��X��n�K[n#jo����{w{�u(q���cU6ݹ��>��a�<ޖ��C%�31f��4�0�A����9��J��mA���`)�H}f6��K�^���޲�}Y�d�hGWB��eb��	7�*�L��6���.�<1׬j���I�۱M��^���p�fM���Mݬ�;k~�OXb�/�<Ή�!r���\p�� ҽ�b���
D�((���7�N�Q�f_!](�v��q�PO��o\�ظ��7�r�I'>�EЮ&I���Փ�y1n�?�(QD�o�}��sdCO�>�s�
����J�~H��<��
���4����׊a�����B���H��R;��zf}���x�I�Yi_������Z���u�������p�a�o
�imU��q�O=�hٜzK:�`����UkQ�v@�VO�����Cb3m�����ɫK�U���ԇ#s�y�|e��y�t�q��
�.��	]�O>�=�6b[� s��u^5n����)f�R�p���E��|y��m��0�Ƀ*c/��f|���H-�-�d��=����W�itvӲ/95_4;�bi�S7y��ݷ| ��R �H��U�G�0��[���2̯�\Й|��b�7Gr�˲J[2^0(��L���Ut��O���Rf�z�7-����Γ}8�/i��#i��{oX�繩��UƳ�	�td��$ilx�[��7Ϯؤ���f��[;�ofr�W��Vv�p�4��A��42U�mXv#I�t�����ӵ��֌r�	��)�f��Ͱ�:C�SgZ�֋yӅon����4"�,��kƍ�kk�R ���(�z��{�7�9�������4��w�ƺl�Wa��癯߉��	Lxx��vwHK;��Ĕ���B��5K +2/Na�>�ͣ%�x�\��U��Ң�k�qKc8�x�%Kz�W�/sg���l��/�������Q�*����k��>%��z��Z������uusmU�{h���q8gי�gE~�Ԓ�_�����j�E�\��k,�*���MU�]��7U3S$qXj���!��8�0ӻ]�������r�ڄ{�cUu�����u���=�ӧ
�onn�e����\&`����Ug�Z�H?a�x��rډ��O-�sKN���Q�>m�+i[�;dz�b��ݗY���@r�)ɹ�s��"[ʜhv����e�d��|;��?w�.c�6s���[�ez�̀����m�[�g&�:</����z�Y�Ӱ�[N��Ty�Rs2�
h�C�|q\_W]�C���啾{��,Kj	Y�Not�lKiu[;�|n�wi��%�w����k�RH�2����r�˦��{�B��8�/��kI�������!z�=qQ#�p�QE��z��ޕAڭ�� b�h�)�*��l �ky�7M=��]]!��q�_��G����f�T|?X/�:�ܜg�6�4p����-i9���ݚ)�6�>�	6͆�G[2}j�ј���^'H��R��]=c���|ܝ:ܴ��N�}ff(��V�y@r��A��ߒ���v��6�w?wF5�����\E�e��"�V7�u�\X��J/���9�4��>hoT�'KT��_e(�rX�ϤS ���� s�N�;V��nq�����oQV��Un��]��.���>�\��n��G^��݃����3'o�>�����:���i�V/lю�ݽMp[����4Z[!��x���3_x�̨ޙ���>����ӦT�^Tu��^8������+y��i��v�SPlۻ=�ٯ;�z[�]o���(�ǀ&������� �q�&�c4�<�3J�cэqS.���d�V�P���R��wČ��ɸ�N$�NL��½�UEDם
`:]-�/�R%TQ� 	����L�1jV���`F ԋ�T�ؙ�;Ql�R(tBe�ɜb��'f��Y�v��n|GQ�{B����ץM�@�G�R��0*��
 "�?S,V�z7ݕ{x)�@�����?W���#�+y���9w�5_�F�l�'�&D���V�FY�@o\���맗�{�>��̌:��]	,�͙��	0cVH��o��p�l�@��Z��<{�5���n2�>�P¯���o7�`����.�4������Uw�������C�I��G�*ٮFF-o��"����l���ˣtub�>��3г��8�e���
4��财��%
R��*��M���>s��g���)���}L��ez$Lax�W���A���t_wvu�ŗ�������,�ĕB-S�M��5���CZ�聛v�=�[h�􊽨�5�7}|�x�@��?;���gݖ�b�$'�����y��;��`�R��O�b��*�5�.�1�Vl���uѳ
5�h�Hk��~����zLSi�g3�ܶw@PzW{��n$̼�ΦGn�׊WI����A�͇��b�Q�%cv���ɡm.:b����%X�"�|��uvMe�˕�&�t�lցe\u[�%\Х.Sw�r���$��&8��wsԘ�5>�5b�T�m��c���u���S��O�l̸�P��q�%�(�{���ȅS;�Sz��f7t{|�{yo�\�D�6/c��ӗ����	�{�x�9��w�#�Ҋ6�	�d=Uz��Sz,�!{�� ׆�w�Њ����{���d��@cc�z�݁$��h�Tu�t�C������;�ϰj����C����c�T�z��Y^[^��q>k��r��CDe���+_s8�l9��	#Y)�<dK��%+s������5�e]l��W�5�t�1*D:�~]S��ϯW�����cme��r��kZ�q۽����ĝ�$n��=���[���Q1}�W�<�Q���k�[�#�u:���n�zvOc)�cB��(0l,7"df�,���Pl���%���őϽNr�o+�\�&{�;�����Cn���W�&������rF�oئ�z$=^6��ݢ�X�'����tV����>�]��y+N2vM˳�2-�qe2��X�'�\��{	(V<o��y���m)s����~���#��5�[�w�zG���En������J_`�����ض��J"�e�<�\��Ӗ�6�ջ�v&.\y��}u̷��)������׆��wm|�Ƽ���c9Ri*�{!����8+�WK^��ոD5��CF9��Dٺ���3����w��#.':e�r��]�o,��Lǥ��%�A�e�J3���fc{��r�iH3��3��g���l��������?{��/��s��fKr�,�����i�ã��(�%��FE�^Ns��ބ��dF0�o gO��emm�U�פX}�/O<���>�����.\���g�4����}Җ�iE�Mگ���x���"���^\�~�z������@EYp��$x�l�4Le�ڣ�.ΎwlL��7g��`UC��&���� ��Ըi��L-$��|��жO��I���'spvG<q��֣��_����1l9�J+�n�Tk��wd�ݜپ���!���-ޏC���ޑ��c`R��%1����^nMO�ܶ3b�\N���Y3h�*%3.nu
������2��lW<>٦/]���^�F��H��S&�'��uh�qX�&��Ab%�{g�����[f�w#��@�ҁ�*������C,�U6��W�w�����?��U���ױ;y�������̚��7c��Aw��QN�\x��ڵMU�m��^���z�ԛ5	�Y�O�^a{!�v�_1F���R�,�e�����u�}���-��o��tZb�v5�6��u4S��~qCi>V�v���O���}v���!Ƭ�b�Պ+�v6é鷁���w0��Hſm�d�џAIP�}�n����:�?�p�io�$��[���#E�ǌ�������\�=v�Z�D!'Z�Ȕ��ή�M`�<IV��:���Q�R��#e�e�l��-�v!�[���ki�$��PI_��p���n�~U`�����uXw�8m�5��Y�)�>���_�����C�o:����4VLڷx�ڽ˶_��q���5�w��t�}�����U#p��ff��1X���G2�?LJ�?g�*鸧Q$	X�G���FlW0"�
}C;h��^��=�ou�uZ���=��}�����,|��Z]t�W�x��o�;U9�+$T����S�k�(�+1
"�&�5rF^��!/r�S�ϻ�N�`|�AY�rC7����z��0Wj�j,���nJ\��^�/���h�&���D�>I�K�A�4�w�<̏��Q�x�vu�#=��7��$�
��5�8{�Ͽ�]��mW�x�'�,���zv�$EțȮ����[^�Ϳ�ϫ�ނ&�/ߖ�e�3ɣ��U��U���g�[S='f+A7S�m����^�ݢ���Z���}j:@�Q��L} \+Lys[����z�i��x���6�jIu���pQ��<�d\5�s�9v�;2ƪ��wS\�9�*n�o����=��W�	t�[򀱫'Ǆ�g���U�D�X�ǯj�d�o]�1�f-�+�/v�7�D�jú%;md���3����fpr�C������>��J�wi�;@��q��8�z�g3ҭx^ʧ7l��d/�;�kz �e\�~mW�����HP^�����ۣ"9�<�ͻ��,��J��C��p�r��L;�a�"M��]ԙU�軋���W�l�̒�z�c�8��]mʝs㷗����Vk��HuD(���N�ɦ��:�0r�?8pS1����>�r�+�7)�7�� �j�z���^��ou��
s�����j��U�̴��d��ؼj�<� m+�RZ�*��'��e<s\�]ϻ�((n��a�g^>�8�����Fvv�)e�ܾW���SH�78��;�$�ܩ��/x�<1SRn�8G����k|���}���RP`��=;�Vs����P�.��4�� �|�o��mxC����mTE{��lP,p/<Nxr6ެ��.�$�u�lf��;�F���[:�7�0���P�Pֹ� �E@���x�=\�һ�;�u=CJ�t�l��{7sa��k7���n�1��-�*�>y��=,.d�p���5<��s;&�4V����o$V{gbUw*��Vƣ���9kwcT���S�8�v]�v!�Bɋ����A�3=�Jhû 6�'�����ԍ�6�}\ɶg�yzlɗ4�u;������;F�����g%>�D�a^���mh�γ$=Y�,����:�CsÜu��2R1볧�jKw�v�	#�h=C>��w��<{-�)��#�(��9J������,<5q�X9��7���	׀�RY(͛@�QH�=U{Bib�y��Z��74-��,��H�n��
��V��8U��fa��
�c���ۏ�$l�{��n|��4�ƍo}����:4CvU�Q\T�j�;x.	�L��>}%��C(��p?���" �<t|�>�Ȣ��}&�f��i'�b�n�-��Z�K��>W�,��t��F�:�txND��;�8i`Q�.��־�|>��Ɔ�m�b���얅v�ޡ��%cr�U�+{%�{��o.���,c���ò�p״x.�#v.���8��O�l�]��Sh��$�,�p�I�ac����o�-aljH=Q�pu�̔����8�\v�ʽ�.,g'W
!��׵����!Gi�!�l�w3_GW��̮�����Ywq�.M�>=1���*�e�owe[h��3��Ko`�l�:
X�=$����Y�����^���/ᙫf���������믆�v��6�]/��U�-�gZH]��q�]���a����`y�)�)WB:ʺ���Z��Xb�/z�*@̐+*o�^Zۑ\r�>@�L�5³3j*�^�(h]G
�B�J;��Y0\�c=�M��S��ƙ�w�Śnf�x��f��:��x�t���qh�Izi@�.���X)��]�S�Z���U������w�L�'�K�o�D�ds��Ί[MR�(0rs"�۱Y���c���"?o҇Vf<B);f�Q�0���y��iV�U�P=�3�>�$m��`���ĮUj�����͝d;�Z��xVr�y�+�'�q���E��Cҥ���қ�|�\Ǩ��gvWM2M9!Q֪/�������ݢ������4qj��g9w���T<�u�8tr����]�>J�Nk�Y�����Y� O��׎[����ͭ�k���B����%UYv�Ai��T��vݭ����aC�w��8I��3�����u[�ط��-��q���r��Wxs-S$��<��ȥNn]�Ԉ�P��Q��n��el[���\�z��d��4���"�]�ޙQ���'[h�͉8oN0Ar�f�h�N��^��Db�Y���!��KV�V���B�"���>ۭ��Z��$r��r�.�V�Ő|����#�V�N��n8����Z�a�6�7΅돺KM��F�5��Y���Y�M�\#��fN���X��e�8��M�{��mjMU����:`����t�R����(v�p�^]�m�}�3�� %v����V�]���*�F�v(�Br�ڢf�h��E�9�����	�7SJa�X;p��0sɒ�)5W�HQ�]U�_X�z�fB�,��wov9����c��Dy���}����{�z�QKM�M%���$�*�*�csX����/'Ӝ�|}=z�?���^�z����ׯ_�z���������?�I}�������)����j���P}�%1yh���5^�9����~�_����^�z����ׯ�^�z���������=���u�$��������4�4�P�uDLG�uEr��M$�E>@j����DEAS͊��Qq[Rx��D�QTE�i�Z�)�����:�4�Pi��sf���gDi�AW,�m�J�h�P�UTU�1ʩ��("(��<ˊ�ibZZih�tR#Qݨ�bѪ��[DPUSD'1�(���"JB����6��HW,���H�!�5E%>lD]ZDy�Vä��*(����D�>W��,7�:Q��y\v�����R�hij#]�#O�\���.ދ��3�svEӎ��N�k�
�|�
(��rn��U1�k�w�q�i�:/ό�y�ӆg�C
���O]�e�A�tb��M����%�z�`wh�b^㯛�~L5+��tɤ2ʹ!��{��W�`�= 1�]�Iolz��L��[�Ȼ�ꌨb[W����ݽ�����})r�i�߹�t��^^�C ��f�3ꇸU��n�f��p��ɳ�!b�����M��5��+|�
��h��d��eD��oN�;���,`3���)&��1���E�=��{J�_gBmf;<��ܮʢ(�S4^���m6�dz*g�'��Q��n��ҋ�ӻ;�d��W�\���7�q���/��ߢl�|od7)�=���(2;�)��
zg�ݞT��X���S��mm�U���f���C�����eVe����G�h���#�7��ZT���ݚ �̚��{! �s2�^?X�xQ��Ck��jb.|���P�A�5J��Ľ�jW9�z�����x��w�}�^w�\�[8�b��ۛ�|��o��)�|`�A�^%���^��0Tl�W��N��N�ѕ)�dǜ <3�.���'���r�Y��x�Eعr���m[n��X�ڌ���X+"��v����1䔬$�!J�!����C������4"����߮yw�9�+�<�6���xt*N��B�[��t��q��̻n=k�M����@��3�Pߌ��E�[?[!�)��{uW����,t�?�gI��D>��2ّ��D-��Ƶla��EWU�tWcEp��֌$���J�nF&���5�����9��2g�W|�Tɀ�7�6�2:����-P;����?;U��sQ�+��/Ū�I��f�]W^��F�T�Wޔ2]6Byv�삦c�#+���h���nfԄ{�Xd,a�#/͔r��z����Q3M���r�i�v4�H��.3Pw�b�WV1�j������Zt���ȣ~\��Ӽ��v l,�A�� �x�Ufy��p]i�;�g����ؽ�ק��;ۄ��\<:�7�'&4�i�f�ÿ����>�[A� uI}��o��ӣ0�W�)͡1٢#��tq�#Ho�	��o�no	E̜�r��um�۫S�˃��,4y|��c17���t����T��ݦ���+��'!�_)�A�5T(Qa��D���5���ߏ�<x�� ׿�9�y$�2˫�p`�S�^�Vdgw^2r| �f�.��1G�;�!��d��i
�\iY�}�����':�eZ�#a�
I��G�ꁫw����C23&&/��͗��s��U�� ��C�Jj�=fVP��r�Kj�گ[���v�ɛ̬��rf�M��f���&W(���d&���@YU�ҷ@�r�&����1�kd���Zq4ۑ����[-}T�Ίװ2�"��	cf+h�ͅ1�w^�U�<N�׮���z;Ǻ����!nι۟e�r��9w�m�m�����K)�,�rաj'��[%� �4��㱪����uOu�;��Q��l���T��J6Ű\V���{i�v��w�~yߺ�[��7� =އM?~JN�E�HKo�šjƬ���.�uJ��:sw9��A:��	S4'�S��/��{�tc�\��@�-vR�>B	�pՂ�b��#uk�Ѳ� 罽|bxV�L��]�;}]�ƠK޹�(�pEC5�:9b�e�c��걡\_`�뤭y�q�{j��Ů\؝J�Am)vƋ����k����fCF�7�kJc�e��s��=%�<���*���}��.\�� .����:�˾=����ň�F�Jm;��a=�nH}����^�dmWk�E��qph�S/7Pc~�m«��g���xuUn8ன���y����:�����>gc�/2�`O���ap�����bt���1�䀵}��-�3ή;j��g=���7���<�Wy������U�H�kp"e���#>� �X��m0+S:�܈i�-��ʲ���-��!��?v<R�k�e�'��¢άf��%�Մf^�
}�ٺW}{�xR��v�n���t=�"zlUg��^牍��9Փ(s��������]�zs�\���Y���v��:��u;cm��b�y=׽՝U��x�mx���hê�\*���?D�Z�"�"*5�땻U�͝�׀�������[J��]�=�����mʇ��[��O�5�dcm�}`�X�+ifMȟ{smj����������6]!�:�+���	Z^��Y���.H�}Ј�.HX�չy����n`䥝�%��W1�2�Q����d.�y󉯭�@�ۦ���xC��|t��\�E�k��*����k����@��h��l���G�n�%v��p�y,ᪿ76�2�����wOtF�R���h���g���xߘ��[��r��)M)��aޣ��SU��_\�{�6��y[����¤�Wi��-I�gi�^&����}[˧�nE���Ғ5�,@n�v��tv�7��K����海��¾�P���흁P!�h%�{��-j�3`>{{<��Aפ���3!�k�@�S���';���<y$t��"w\o�9�ʹ%贆�t96;BxYu9Em9۰��t�̐��}�n�D�d�dݯ�`w�5�(SN�w���U�E7{xk�͵]�go3�,b��6�ss�i�v���^�@Xj��{%�!m�.��c6*�_����:�!a59
l_]��^�rdo�T��o�{�7i��/V�&a��5�A*}f����i{��'``�W׃����ӂ����SO�:�\�s�,u�َ\��h"���uf�e��NF�c��QwNaJ�[�nu� ٲv�;L��NW�Eٖ�{W8�i;�N�2�թ��e=�4h�c%�(�gc銨�%7�=��v��Z}/����zF@��%�[�։vSe�I��l��bJ}��׵cG�S�l�wʚ�d��V%p���X=�����H(�O�����?��ѕ�Mߖ�fV��]�
�������v�MnA��W�m�'�o^��|:yu��iP�^��s�'��v2�Zc3�p���Q���������{�h��Vn��IJ�IV�:g������ս�-���d�YB�AP��
��ѩt���5�$��w��`�7ُ{;q��Kyv�����3,�-�::m�4���ul�-a�r�7��5�m֓��;A�2@⳨g��ǖ]G|���L����veWc<w<�/f���jN	���m78�`n�e�N޺z{�l˕����ƞ<�
;�y��0���o���b��G޳����K��De�cC�A���Ø;��j�kF�Aη���&�Omu�p�2���&J�x�����P����_>j����h!*'��R]�s�[��%0����/�Vc]w��^R���T�4';X��*/�vp��7��L�.�r�of;�:�(��wI��`�@��2.�C^st���ng�p���-d�Z��u��r��r2��GN4V���Z쭝�-����D�݅�w)�&D�׵�?�~N_{�r����3 ��ϊ�wNmqGƽ�a��˺��p��������nܥ{�76�Novu���%��oz���sS����cͅ�B�x�RZVJ�vëFEl=�`'��8��	�Ѫ����Lڥ��wu%�
���2��s4D�Wu�����r�[��0���$�ϱ["��}-e�8�Omq�Noi�!�fC쫩݋�T*��6a]�R��+%�g��N���ڳ�{��n=;�&6���	��B��g�|���a,�q�jN�W��dm�_�k�������8���@Uٴu̫��ׁx˫��~;ٸ������]�r��w�A��c��}����x�W��[ۣ�dH9�-n���M?R��z�o^~�)�o�jtF��8��66�K{l�mn!:�ޞ6��\�<��^�0��]r�C�$�]㭰���^U���iK;�=.'�ic��:,��謗Hp�O��	� jS]�a�NSFF�69�{h�l�@��>����x޾nHn\M������wF$-�B�g��ļ����^͈���b`:P�w�P�`���oJ�m<��� ��]?��7����9Xۨ6�s�zك��d�����%j�)d`+j� �zw�L�q�<Q�Y�Y��:�)�½=��+�]H7�q��pB����oj��-JA�0����W�C�a�d���:#مX�ܪ����U���Z��Ҷ4ߜ�-�Y����;w�Z�F��8yVz��k�3Y����;��w��:h�3ӈׁ�2^��ׅ�q��F_a��U=��ٓh�_<�P�Z��W���h�[�c\�vá��r��v���r�U[ߵ9�|���s�*w�}X�|�c>�,@P���uf�S���ֈ˷�npM��Ł�X�S��`�ز�Kߵ H�1���jj�s3f��ah�?:�4����˹	V���CD��SU���ws�<��.�f>x�'+*�ꙴF5�4� `���0�fG����v ¹E�[V0ws�f�����sS+�W˂�Q!����p.�v�ӽ|����ڻ��N��_�E[^/7=�S�!��zS۵[uדW^|@T����)��!=��2�c�jw�+,vɦ�|���o�+;�����WnU����% G;�ג�+^j���Μ�h�>v[֯$wT,㩼e�}��W��@{����-L���9�#�x��t���8�6��*z��3!��\N�K��U�_v��bH��+=�����`&�2�m�=��/EQM~G`6� wd��tJ7�d�FE�Q�)�/zr�7�O��Ж�~��M�y�rR��Ҳ���+��nc2.���Ȥ�շ��!q��1p!΀���R7GK{}@u-S�騙��_'.�T��Z�Z��3���y�>tC�;�j{`Z2�z^�+�����f��w���g���m�Nb-��o�k`��h��F��NGM[���S|L�v���-\��y>7/��6h`������J������7YN���|�"ukv��i�S(�=V�{�4fG���i��z'6�^գ��R�n�u��0��g�s�h_`���Z�	���#@G}3��{&XK�4�v�{LvM���*=p �l�Z멕8d{ۯ)�'e}/8��������Osv�ɑr���,���ܓφ4�x�� ii/.Z�6=�+	7��k-2ۛp6�i�b=��m���3r��Z�ͽIN<��2�d�LVu�_o3��K% �V(рfz��ચ`�&M�T��vק,k�/SO�񝼂\w��.��ͭ�F?�����qU��$�����Xs;ESD,y�}����"^V앮�`�35�*f��]�5���i��@d&���$�%�gS%kZf�fa��ݷ��mzRq�G[ܖV�f@�N�X�f��`��{�KV��w�s'n>˵V�y �;=�]T�p2+��Kd��qڂfky�v���M� �Ǆ��7s�@�R�F�< F!a�~;��<���R7�&�\�[S����M�{��1�;��K6tԇG'נ�c��x���y-*���V���՗���jm��I�'m�y\�R�p�:�:�n��gv��ب�u��T'��	�i
��X�HB�좏M���˯������tƍ"�o.*w�Hg�ro����9` �xeÕ��2�̌�9�,�����@.�^�=u.�Hj��[�ܐݍB�<:�;c:����*gb�v��r��<���@�-��|EN���L�V��WZ�#��/NuLB�5:��{����7o��J�"��1��V���ۗ�7��O�eċ�쩊�ή���-����ʦ�.�*nrCMΊ�z��&��K*Yޗ�d���`�	���x�IW��l����7��3��$�:��F
��u�ud��oL��,v���rm[�:
�f�5h���V��=�]v3|�o!i����,D
$[���`63��fg'/�ޙx�$���
d�{M�Z,�t)}ʌ��~ݙ���YW&umG�+dFH��GSic��\"7Fr�oh��m�2�7J��siә�6�wIܻe�\�Tj̕t�u��id�~$g(���1kU�*��q�j�[
�r��u��^m����À�EL4Z/R���p��z[����U� ���;��.�7���ہ�:i��I+jvZov�:a���W7+K�	._k���bV��u�di��f�6\��Ƽw��x�5���a���qP=L�^��Xs���[m�t(�Ы�1ZW_��l���1�б]՚�2u���]�]H5D��Y�2��R�c��"�n�L���`�J-���L��RPPI,"��袈T6����9�V�yC��*�V��̝f�{�	Du_̜U�r3�Z�T��i�4%>��STcts#y�!�UFl] �`0���Kq���W�
0k艭�
!�E]r�=˔�:�Ty�WN�]ͻ5:�W���bޕՔL]��е��5��큒�_1��J8u�v�у�)+2�,Ι�����S5�D����ty�Y�ܻLC�9��}i����=��h,;�_VT\��d��h�y�m�tR����C$�Z�Q�3��֩)duزCA鰻��Z�x�wBץ��RX/���vi��7-��C��K��5����ܻ�X$�����4ޜ
s�Kqc|fSg-�ujbv����ʋb�ݠ��FƩ�i�M�ֲ��	�վX�:�au�X��繛Ps�ݏJ#���]�`�ܫ]��,�~)s�pU�(2�U�YNwr[�ls�������:K����OH7�:ݾ/�����.�IV-�a䊟tb�jI������L��h�ϥ�G�5�U�ێ�@�H7V̳��С�����|;����k&�c�X��{��9��"w6��I���Sb�;l�G�#�L����v���(7�FۑM�����d5�8ݗ��&�YƢ�"�t�p�Ϣ�AtN\zS)M���y��E��{"W�Ev�}К�wOxq�=���ɏ"���6.�ݛ���PT���h�)�n�
$P?2~�X�@li�@t�J��>�QZ��ʔR��F �H@�LI�H����t("�㫧VMY4� qy����=n^_q��=�嘞�'��Mz�ڊ)�(��Ѥ���f��/0o3��><x��8x�����N�:t��GN�.t�ӧL>>>>=��Op芆 ">Ζ��-� �"��j���QE�8p�����N�:t��GN�x��ׯ_����l��Fa��lE�:6܍,ID@Ly��A��h�%�4�/-Z��T�y��͈�
"9s�ZJ����@RZX��c����<�"1��'U�sj(�Z�_W�[̇6c��AT���y�����ۜy��r܏a��O��6((9���l�Š�&��܍sgQ4[8�Z|�h8U��[Z�lf�mmC�1:Ko->��}�����-k%��*[��@b��T�#����:��w�i���opv~�{��^����D1t��a�Z;���"	��t���A!A�(2�e{�2P(��*��q�wmM=&�x��m�� _��Ng���K9�|=Z.<e��
�O^2-�
��^b{�ة˶��x�)ya���)e���c�x������z|]����w�l��d�7�P|>�}T-����{{}خ��Xt���׉��H��)M�8w;�^��H��U��n�{�x�z�ԓ���5��Z%l���;���o4�Wu��3�v��(|̐��ӻW<���J�+7�;?tQ	骳�Ľ�<��:}���.ͬ��y�X���U/ј�A̡Ѧ�:|6+�z�p�_K��&m�~�"�\��+V��J�Ӎ1�D@y�Fkxw�W�UϹ���3��Ǖk����b7���ǜS�rS������ ������+�T��`�f�ƝO�bg��+��&�6���1�/E�"&�E+2�8��W�E��l�w�4�!~���٘m��U����U��'>����U,��\�k��V�bl[g\5������=�H��6Ԇf�����tPف�B����S�p�0�Aݜ7��צ�q��˯�MF��@C#��S�-�٘H2\l��b�ֽ��]�ji�
�o�����ة�~�ꆻ@��r�>��Nتe�9��x�YF��ǎk�2�ً��ۆ1��57�K���DTf�sǮv ��"ze�o3{g/�5N$s(
r�����f�+�a�)O@����c
��鳻Gw�ou��:hY��Q��9fD�ږ�V����2j����ؼ�z=z�$E�fx2D������<�cҺ�Oe��cǟ}�!���j `�U��ili�/D���
+������+��qK��˹��+�o�Z+a6U�o�
�˺�+� 1�b9�:����op���W��ܞ�x��k~�%gi������~�k�߹Ғ�,�EY���ͯB�)�9�N�t��E��wY�X�Ǹ	 �^H�`�2��`\����M�9�&g��8�����2nzNv�i��#	Y�:��6"�o�n���-M�qg� �:*��`���ʹ��Fm�G5n�ȍؿ�"�ñwf(�Ω�����u��T���@}����Z��%gc3-eqX�M�2:y�&V�C�i'8�g��h�)���d�|��<��)e��J��6�w9s�y1ܖ_?�Ub]]��[+R�,;�5s���e�L��xm/ݦg�N�8�~�g�p�.�8���#�������8�`kG��WV�o5���y�ʪy�¥����^�s2�op.�IlȰ��ZB&�Tgf}��7>���f�R쳵�6K'���3�2�M>���T���.�v�k%�R��n��T>3�?g��u��ϛ2�L�ŻJ7^���i2� *���t�m�������M��
��{,���6�ջ��m�P��|�zC�Ԣ�ۦ,bx��0���PD�ʠV��Y���8��̫6�op^��u��wȘ�U,�c.^ ���p�z���Ֆ	K��J��ܪ}�^�i73zat]��Zo�;��'��O��f}q#_��Y�A.P�v��ݎ<�-uӻ����,�b1�:`�<%����KFrS�]�D���`��T�2��9�GKվ�w�ǒE��P�;��*'L��(V��r�}���:�P�yV�)V�䵾�<�0la,L���:@�	c�C&�=�N��(���8��©���Ǌ��M���A�R��c�P�:LY)���/w�̧V�5�����{���c���o�ёrڥ�Ljެ�I�EzF�%�2#��4��{9G-!�qW��V�F��ɣ�h:�!/v�n?_����z ~��,XNwzv�#2���Ub�͗�3 �o��3���0�l��l���g�+�M�z������+��0����Q<� �Lwdo���L���ius�LY�j݋�ʹvtD�5�@W�.@�sp��v��y� 3���s��2�����58��������3�k=>Q�Xn1�N���B��yޥ���F��k�X
�-aH6�ws�實E0������4���M����"�X��Li������?~���z���*�Y]Ȇ�js�/��
3 �}�\zP�who3�l��da�3�}���f�iԌ�g�������۲�ݨ+�l�c�A��T	��V4L�M1�.��{��n��θ����.�������n����*���QnvĞ�`¡�0�j���T/yJ�:��PF��ꬍT�F�M$��*�)�V֌�ECP��_vS�eCjq7JNޫm��pQ�gZ�6N�S�d�m�cBƯK���qa�D�j�qD~�����5&*�|~��|[%�is^�⇝�a�@�b���v?NI��`�1�4�GV]�`�?e x��Ysj��A醌j٭ڥش�#���+��G�J�-��3��Ko�)K��{}K=��3�b�S�t�ս�߻ͼa�q��-������l#�$w{#rUu�Y�Q\P��g�����k�3��lp��y���d֨��&t����k�&�tV�פ7I�iwH)gW��z�q�c��O�u��xD���Wjkz�$�qM�/<W*����n+8�^m�� �m����ε��7�FL�Q�0��b��	Lcۜ�w�IV[����oY:�dHyt�T���ݜ��
���o_��l�@|ɜJ�n2�'$ �H�Ut*xU�{<�)��p]Рd�А`��9�t�X�jn���
�p�r[9]��n��H���r�*���2�d:��?���c="0\,8.ͬ랶���|j%�uQ�g�r�/�{&bV採�W8�#�����t�H��Y���W�e��'ˀ�V��C-ɞ]�LE��m��!i���N�J̬�b�u�(�j&��x�g��b�������^ވ��.�n�P�l�����j�0���	�M�9M����.1س��Dr*���S���չ�!���}Ms�t���F|=9���a��L����Խ�h_��9�u���7��ؕ�5��#xo��X�Ba-�-76+����u{����4��'^.7�.Ԭ�y���r��L��Z��F�3�����1n�|e��=;a��U�鎶)��8�+)����Ł���{�x�Nv}���6�ϧ�=k�cg��3Rd
́{|�����P�_���{��W���T#X�S�:_*�fQV�L�C5w�*=\l�4�͗fV�s��٭Iol���	-�k$Q��Ἔn�	ݡm����1ԈXÌk����8�^<����عc+v�K`J�ʎ�Z��wv��ĲDLW^?f[��s�ݯ��ׅ�r�\��+��+zۊ\ݹ���ˢ���l�v�M�0����խ�t��vpz��{��^�A�$�"��72���.��uøΖ:il��DbZ=��&XN�=�d��jb˫��������3*%S�=)g��ry�_tY]��L��{:���QANts�ɏ��������o7�:���	t3o_S0+F�o9�ˍ�J[�w��2�%�H�a9^�Wt���۴w�5} �v���;��#�kR�q[\4ų�eb���Yϫ�yf0�#5dfk�c����h�v#Y?���q����1q���N#����?m��>���֟`��<��ݢ����r۹��Zy�t����������u���5#�sŌ�?N�1�y-�қ�}��7Y�P���@J�6,œo$�pMpG�#lU:O�vY���cm3⥝zF������O��)��w\�<E��O���V-9���@᧶9��I�:Y�М
F=]uw�q��d�L,!�W	���W�O��"�Q�j��c12��C-�]5�̷�����-	��)�zܘ�K���[�>��Su�\j�����4��-��M�,9B%����y�gF��r�]��m+��zye�B
|u�»��Ou�U��2�Mk5��Kή��Y�wO�Qu�^,���J=-,�I�Tˮ�''R=r�H�ͧ�"�;�ЩͭP���B9w��R�Wl���x����{/�ځ|�����K�سd��ͺ�e��j�dş{͇V��Dw��P�Gn|5�5Ҽ%.7�}[B�g*��T�SO��ݞ�w��,�	�.!ky	�����.N��q\Z;S���za<�����US�O={/w�\jhĚ����%�����@��=�+ʁ�g���{+oq�v�;gl���%�b�<����D0ս�-��>���Q5G�rLԛ��o]�:���	:���A]ק�H��������N�Y�8�RFgW������Y�F-g�3��&�߻�^��-�����T���t�{�"�I��{���6h���Z�'՝�{~ڵF|Z@�*Rq�p5���,]�8:�n}Ɵ��{v����2���mp�Jm�A���`�8��X�^���+s� �hx;��m�B�iܬ���4{�R7��wuZ�tPr��;.��=�5���b��1�J���8�d���9W�u3U��а�_@�p(Qڸ���rQ*����.�X�Vɭ�,4�n���κD�!m�Qڼ�S�͛ӃH��YY��J���H쮭<�I��|����]�wTu 8O	&wd��\p�,X��^�w��ϛ!:��-W�_���Lx�k-�lK��b,��k���lXx-*z��u-���q�zEp� q��8۠'��Y#EP3.��?��|�������w�*%��h��Ω'��V<�A���L�R�!�����ʖ�Y�ۖu�]ٮ5��-�	L�����9��<�JA��t�b��7������6Fl��Y��;�L��K}���.�q%Ցٚe�ٝ�0nW�V�J�|P76�&rf��8���s槦Ul�YJa�{k�,�T�X�W���z�q���F��P=��x�	�]��4�� �t�۝��ѓ
�xD>�+�	�˞�����S�<���݊5"��|�-gG\��÷9��4.��c84��d��46Z*���~̓d�>��_{�� ��z�Y����8/k�m���9^�"���%��8u�����U���������^$!�0��w0�����^V��c�V��RZ���Ӗ��3����]��Pa�#S��O_�ڔc�n�`�b�K�[�!��C��]ܕ:=��^o+:5���O��{Ӻ�#+�x@�$��t��˸�K��Ŏdl��o�Z&�s�{β�Dz]f��P��q�����ζ�Ɏ�ݬ���&~�n���L�Q��l�ʎ�(]�s��Û�fz�ެ���#9�[�����6�ܨ��Y�{	�s�vYn�-C>O��4�����2$קR�@l-�Jf��1�Zm�Ζ�v��L��zm�C�l2�;�!՚�vf�����s�e.�A�w��W��9�(w*��:텞��׀����y�gtd��KJı1��|��m(�k�z�5g�]^���|U�Y��ҩ�6el���cp�����1
�_t�����@�� �z�xw[���+n'rrZn��K�l��*M\� <���z_����8��.c��{��̎��@����Ym0
mR�pйU�z��S��D��c[�9K�$]V��\��Og��h��u��(�o�9�Yu�uwMo\��0T��Kr��ܪ�҂&؊��L��ܺ����V	��[WtE#�CSgU��X�h�Ϊ�V�K���R|F��x8���oܧ1EH���` I�ɫ�Z:��.���?�; ؍��(f�v�f7��j���*#�Z����
"��b����3F���Q��%�m޽���D�[��r%�P�l�E�s��c��g�P��B9B�#)�ҋ̩��x�4﯈C���!�8o\�e�}��t�-��9v+[�\�(Uv�*c*R�|25���"��
�<��A��b�m+�u�9t�"o[�w�m��ɯ!�SqI�qz��giU�1RV���)�[|qkjG��A/xf���t�mi/�D,|1��fpԟb9g�Y9[���]"3:��G)���᫑b#�`#��wY���rT0c�Y9Y�]�9����X.��t��Ǡ���«S�E���X�W�;�%{��fo0d�.j�"�5k��u2�^���;��_ΉUu�Vs�о�M�v�h�׹&�R��]�R=�t�JG���H{�KP�gS����k��`�dL۾V)��
I��h�d�ğm��ȸ��dԉ�˩�&/���s�6lu��ݮ���*�Ͷ2r�͹�M���{3Mi�I���g:Y��D$R�?�u�;uv���;&��(�%7� j鴘����a�����"�V�&V+�l'y�����:�1�p���D�eȻ�0l2�8(]�kZ��e6A=3�z����L�ܮ `n�u��]M_�VB���XY�wsLF��򽬠�>���|���O'��6!�,��!�&X�Kyz�Ӭ�"�K{+9��q1X4$�ު�_su��N�'BdZ��������,���/���u�_LGy' �t��"�������Vf
䭕	�gJ���I�z.�\ᩫq�+o2�4V�3{4�a���e����Τ/A��R�9vmX"�0"|wNԾ�5�;�(�d!uL�5L�	���}�F��k�U��s>
��2�:��:�����d�%�r���dk�=W���<%���8��N��W:0u�"Ds�d����R��7F�� "�$"�Iݣ�y]s�0�.�N�]��w\S�7�}�ף�8E�����wN��s�]����+4�]�}{�gu˂�+7�.,t�W�|h�E���	y\�J2��y�cx-��`�⁈��֨]�Cuᆑ�*���Lv.8[]R��w�⫔����:��d�u�*ͩ�Km�Yڞ���u�ԝ0f�z��o33O�U��k�mDF���%�#X�k:�̔Q�ڣ$[o��>2l�ç�:t�ӧN�:t��O^�|||||z�}�,ڣ��nb��+N�э�:����l�np�Ǐ�������?�G�^�z���Ν(�ӧN�0`����������h��1�F�ѥ�@�c:0Z���\�mcgj�[cb��.`-�Z��5�kX)w3�l^Z+ͩ�i+[[F�,m�4��͹��yp�j"6�h�4kk��킵E.���U�$�� �v���8m���s�p�LZ4�hڇ���95;ۑ����4cbڴ��I�������IE4�Q�gZ���&��,F�O6G�5�(Ę�b�X�"�9<�E)TMP��P�H�R�ט�.֜����8�uee��fvЛ���-R��΢�2bԫ1��u��w����]f��e*���=��X,YTzv'-�k=��`u*��t��±⭖σ�W>r��&Wbߋ��;�5�i��P4�H焰����%z�����X�&M��S����;��F[��+eՐ~M�z����vb��#a�V퀖�����ͫ¦~1K$��Y�]@����35O�Ws@��#ao)#����� ^���T��/�c��`��@�Z��g$4��2�;Ŷ@�ؤ�@�ޞ��$�UK�9�qOd��t�{�UO�e�BƬ�2�GՓ�)���ި�y���l!p{��w6�C�~�{�D�j��f��v��=���s�i���۶�G;�n�ͰC�<��U��� �3�����0ih��n��ll��{{���0��D�[�r٘5zƛ��q�l1��$h��Q1�o�Ɦ�'N���Ҟ< ��P�dYs��������>�uZ�dp�p}�lc!�s�m�J��3]p&�d+���\D�0��x7�ŏ'V���B�[� 5.���>(�ѹ�42��Ua�Ư�,@9�X��z��3�"��O�X���t�s��a�^�������o7������b;�� 9�@lOp�2��;X1��E���vo.��T蝣��8>�#r�gSjg�<D����;0��&�mKsט�O�?�����ck�7�@����f��4f|������]x��T��b���E�v����C)z�[������j{_T@m������Tff8��[�d�r�s�齁Q4x�}�X��+hY�J�m����B�M&�9�%�����h��̔&dL7�YKC��5�dk�V���^*����>?;��
�*���u����0�{��]48�Y!��"�qhq�]C�3�yX9+�E�|�}ޣd���MߩVvU��{)��g�]�Ի��h��I�̿Si�$E�'8��0���!�w(��#޾�09��M1Gl6���I�:��8=��5����Y����A�:�%s-�;+ �4�BQk��-L�zbb�BqOvmۆb�?L������*i��pƺm�:�v�,�Ƚ���b���u�lc����5��Ƃ��ZU�}�:�U��o����.���w+h��{������H����7�����[�_T�TNp����Z�A�}�\}6˂�J@�I!a�@��2"��_�?��o���i���hau$������=ن�Kɵ�x^�|!��@C�ъKa=�	�j�wF�G5�b*��\ȶ�����{/ei�w�ͽ�&�n}���<��cÕ��Mɀ�Ţpw�{"S.�������ʱ�d=�l[�9O�lȀ�͋�X2k�79ؙ�A�e�vae����u�������K��%�B�:%�¨`�m���f5_\��3	��	 �Tcb>�ɐ�}<�7Ժ�c�U��|!ƞ��NE-�×}��v���L�x�N��p0�7t����//��j���6p��T�;�����A8Bx�*&ϫo��d�!�k�gaY��ў�fm�gZ��R�����d�٭;�}�+��0�ml
�j'���?��ݏ�5z�a���.�Cm�f���esE3�R.4�aow:Y�d���̀��N�!Z�F���9�.��[��";{Z���E�����lI�!�NՈ��:6��ճ �U�J��u8.�j�B��P�,՞�_%�����8���B���f>Lk�U3���\2�ֲ�}n[�J.�2�m�CS��|�u�9�^^�y}�մ�oIW�5�)�ԇ�p�[�i�n��xG�w1���w��HQb�����`WH���Qc�Ե�C���Քv���ś�f�]Z�Zѫ�[V�C�Iv�,��^���el��%���F�Nw6MK���Nb{T�r.W.�,&��d�Y�y�čjM=FY=��;gy�D�!�LAޯLlz�J�����*�w,eu��,5��66���{���s'Q��^e��w��靍��Z��x��z3m�Z&����nl�W[�hha�j�KMw� ?d�~i�$sk.@�t� �ţq����	���Q�'k�_d�+�>|�k#��>�7�l2��OI��!�#)��G�C����}�x��ku��$�1G�F�t0d8����{�t|���ۘ�#����l3V��[i�4]mӞp�g/����lδ�Z�9�1nC�5�vcO��UU�{&�8>>�ثۧ~K��v`�9��9��,�����T�جt�tNla�6�R̘�̼Π9˶˓�0o,��LY��Ts3��g���:~�eh��k�Z�s��mپ��y�3&�{F�|<��u:y�50�Z�A�����n�uAJI���ލ�Y����_P#22;yT��^.fuI�O$S��d4�.yˮӳ{�5Qw�M۲��%�)����eO��	>�^�]�8��ͦ;S6l������j��J�ڲiK��122�q�$;��_��.AQ��nn��ܶ.�O^�c^۳��a��#Iݳ^��0��W{v�x��6Č2Z�ݟ	��S1F�o_4�gʽ��6��	,��b��̮�w����s����{�m[�:#jRr;f�G�W����ȃ3R�]Y���4��wP�����1B�ϔC�`���3r�ӎZ+�f�hf�m�ry���κ��#3��j#Fv�0���&�ή���4���f�y��W�=V��љOy�{���HZ׳����v}o2GO>�}��_���
}�{|A�G)�R�Kvx�}��n���!�C�?��]��F����O��׋�I��.���:Y�S��t�_��p�V��L)Ώ՛p7��f�n[������:�`���37���������k�8%#��n����z��o<n����������3�{�I�jh�8oXM���+a��lI�2�w��k�E��ҏf%q��N���~�4�΂�Mo5t��ˡ�OY���/b��7����84ir8�inY ��i�Zz8��(�e�>Z;]��}�o[��P��Խ#�b�<"�b`wv��ة���e�F��vƞ�=O��k���W;gB�Z�8��:hMdt�ɖ��t�([N;���:;ni�9"�{��c�\�l]獆�iH����<�ZVS���!ts��Vp:z�E�ѥ?�֪fde���v����u{��O���bɊ殷�?���۱�L���^'�F{�o�ы�:Y	�=��+5b�{��
�r��}�)��M�]��u9�(�Y��V1f�ۺ���m��9��7�6Т���"4�"f�n�t���q�T��	��:���L�#��o�uXD�w	�hȕ����j�-H&�������SX�of��gs&����w9!X�
�5�&�{�J�E���5�a����]�U�HNV��k.�+�r\�W�)���Ӊ�UNT��
�,��y����Gn�����衑.c�N�M� ���-�@
�l5_����|����{3ҳ(�ME�/⥏��,����^�-��6�)�9~��CF��ov�����(q΢ov�H����|[t?�n�n�����w�{Nkͣ�s�YAn��8��<>�Kt2�>q<��p��mHr���L��5g�䓗gy�s�ꤻ�,���a��f~YΑ���薽k[��9bjPw�u)@�&�q�H7���ue�N
֩����<�n_<���9ۧ8h�ZS	�b 숅/}؊�']c
8Ԏ����a�Z�w;6�F�����y�0�sˍ��r`T'���g��fq���1��朩�h��y�������;@]�T0e^�2�<��f�᭮����NL�X�0`��A��]ۃ��w��x?d2/�׫�kɋ4fD��5$4w`���R)�v�s���B�9Rh���錄�4�u4�+j��,:��֥$RwB�w�i�T]����f��4j�W���>C��(�����ƃ��To�Q6�]4��_RI2}ʎ����/Q{��1RV1��]�"����Kή�F�S;a�[Kp�t��#��w��	����k�Or��,u��}�꼬�<cn�E���s�.x?���W�Gu��m9-gS�K��g�wM)�<3�ZZg�v��fj��Bx�*��9Z����t���ו���b��쵩�=o>E�.W�QP�a���ww��WV�#��Tx��Wc���e*�w+7⭘v�j����~7!V����v�M9�w*�Y�!���b�>&�ɜ�n��"oT�`�^)�,�зbW����lk[껉��Ò^:�E8J�*���;��=C�X�T��5��Ե�Ա�[�����CK
�EZMJ�5�ޠ�Աb�Q��<�)���k)��q7goo3�X��1�~�;�|��Twy\��q�G��l�0&#"��K�5n��^�tτ?)���;�1��ю�4m�A.�Y�J7����gݻN'/Z'��#!�u"x;�H��I�&%*����L��0���M?8��yvԱ�T0m��S���=� mtOb?�e<
֭]���U��Y�����S�(�Bjc�!�.��1fP�8�{mg[;}�Vv�K�鵈�`���+2T��o�,����]�+T�iW����y�nq��=�|�����������!��ϒð��oj��Ȉ�����K�W���/�/Sku�6B�7A�p���|���]y��i�Ψ?m�����G�>���N�<�x�Ň��l,2w暤��|��ή��h�0����.��^5�N��X�w��\����.���]��n:����vf�m3�8�k�D�++˳��o�{m��c���s��ɗ�f������N�Z>���\!�����ӑ����N9?W�)R{��彯iy���/��@���J���1[�m|�ċ�$��iv���hŹ��
:�K'W\`�N��˥��x������e��Z�]i�^����O�Ԁ��ȍ���Y�@�{�3����IG�C�I�Xޝs,х��S[~K�=^蔮��.7윓+7�d������A?� .���y�2�a�RSJ�s<ݱ�JEs��a#IG��k ���O7�X��<̙�@F�>���ux�oms�)��rږ訸h3o�Wg]���k�Z�O>�-�	)�j��A�D�Ɍ�w�ٖ�}����4`��4��h�,o#�dE,܎��o-Բ2�E��<�F%��v���~�ը68��D�nzۂZ��ϙ�{��eq�>�4k��������y>jV�'' ��e>{6Ӯ�7 lW)`~r�Q���{�#{�#qq�=o�5f�X�a6��̣@u}�j�������ٳ��:��Y̬��>.Փ��6�SUt�w�����ج�9ݻ���Vm�k�i�+p_�U�����֎w<���B9mխ[� X��8��@��ĸ��n�v��f�ӱ�=��Y���w��4��a���P(��p����/j�1s���bw��]{S��S�{n�A�W��; �m2`�����{pѯT�=N�,΅�}���J�n����{Ƅl��al2����Ϧ%������ 3 H  I+�AA�Q�����yQ�TEM�nS�����0$!(��0,2�2�2�0� C
�� C"�*�
�(�2�2�!*� �2�0�2 C
� ʰ���C ʰʰʰ�0�0�B0�� Cʰ°��2�0�!*� �2�0��C*�*�*���C"�*�
� �0,0�0@2 C�����2�!
� �0,2�0� C(°�� C�*�*� �2�2�0�ס���7�!�aXeX`@�U�� !�a�VV@�U�U�U��T!�a	GՆU�@!�eXeXeXdXaV�a�aXeVVVV@�  �U�U�@!�a�a�a�a�B!�a�` �U� !�a�a�B@!�a�eXaV ��! � !�a�a�dXaXeX` ��``heUY�CC@Ȁ��0
��!
���C
�@ª�0���n� q���@ dQE�FB BP�!�6G�ʂ�ʂ2(�42(�1*!�"�C C(�C2��42��p"�2!(0��(0,� 2�2U��``U��`aX ��V��,�*��*���*��� � �U��U� !�a�xˆU�@?�{��`��{���B��Ҫ(�2�K�0��/�_����}��c�3,?��?��?`9�����ɤ~d$���\}����>�� � ���G��~� _�}I U���� �2����8��#��}�@�   ���������r���W�H�?3����F@~_����f��H$�J��"2�� �� $ʊ�� �(A"
ʊ"(A�K*(C(@B � ��*@�$��� ��d@	E� $  �Pa 	Q�  @ �H@A @D� !X@A! V �a @H 	V%ZD8xE�����8b��D�
 �DK�=��?����f߳� : ���  $�?4���G�_���0� ?�K	�������  $��!���o?�>� �� U�*�C��PW��@AE���<�0� �����	���/��Oǁ��A�='��|4�>��x [���O��h?/� �  O��ixt ������o�}�}�X��$�����0�;�	 U��?�?��d@W����x|���/�ڈ}���?D�o��`�f �_�$ _I�g������ ��8�~���rw��
/�G��׀
������?�� ���1AY&SY�ݘu�)Y�`P��3'� bE��{�ZĒ�hT[5
�Z�m4���j�EU���TF�T(lIHQHV�B��	*�cR��[55F��*U��)$�͚�jV�����!J6�fJZf�mkZ�K[(ڛ	��Y(f)[���4�����SZ��ԭM�f���m���1��(��X[iw7lEh�m#Y�)�M��T�jA�d�V�ي4͙�Z��-�C(lҚ��Vh��U*U����յ�ɍd�Cm��f�
���m�-���jkF���`խp  ����2Ui$�ڕvիfrV�fZ��kwt�٫V���.�օ[vmv�ccn�����Y�N�u6�,��qn���j�%��N�v�[E��ikfV�mv��V��<   ;�z(P�Cж4��E
(Q{,���СB�
=-��s���aV�uv��f��9�mWjim�uZ�c)�)9��mۻZ��;i�qQ��J�:ۺJt�nq��h�5V�1��F�Z֤�   r��i`iM�w;Y�-�fstuJ֩��Wn�-��k�s3������`lijm����n��keV����%J��ٜnUuXS[Du�*h#UͫT3U��k�Z�-�  wz���uW1B�Wiv�M�Z��]6�����\��UT�n�iU
���:����ݭ-�n���J��J�\땬��Xe+,��6�m�Xl�    ޻=5[�n��ҭk���n5Tj��u���rs���5u�㊉��V�U6������V�U6��H�ETPn�D"ҭ�M������  g���j*��ʑ��0�s
B�k�qNƪl�Z�
�Z���ݮꐢk:���U�SQ)7V:"�R��I�T�4�kZf�lԶ̖���  7
 +jW�  -�p  9�\: ]�Z�  3+ : .��P�k� (f��E �ipv�mp٭�J�hڶͫjѤ���  �  ��  �� �pv  us�  ܺ���XP nm� �Y;� ���5�@��6��V�A��4ٶ�^  ��  ޗ7�@c�: (i��:  ��: f�p �ݭ�  eۀ a`-�4��7  ��R3mfI�ֶ1��f�i-�  �� :�YР r�  �n�� �]� k5�r�)���: ���  m�� ۋ�  D�%*I�  E=�	)*D� �T�ؙT�# #S�A)I@ hc&&�M10LL��UP� ��_~���������ߟ��N�1i�|�#diao�8Wi��և�-X��W�W��}_}�����f�1���  c��co��6��c�   m��������_��C�������6~�;N,(@��@��;�dDon�X@����2�S��4n%��p	n%L�j;_Lc-�Ab,	<A^�.��ȭͲ-�7p�i��+X+#f����wS���7Xt.��Cݒ*��H1���q�� �0�ي�R��BV�x�$�d�,F��w�hK�uk�6$0$E+*�ˋ��Z夠j �+/3oKD�� ��2۸66HqJ����(����N^�蕻z��1�C�e
6!��t�G,p��ձ�u0��)ڰt��і2�L��Akp��N���E�#�kl��ܸ��EEj���U�R�z���b�%Bs�o[�0G���朻�5.̽j�9�l���1��kvT�uo\ƅ֘�N�'N�X��
�Gw(�خ�coV���.�Q��ec* ��$ݖ�����к�ױ��,+&���Z��2QIC�弑�G�n'3ft.СR�*ޒ�g�Z�c%)E]���^b3��ut�\j!
J�pD	F@)��,Hܒ�sp �,YE�۬�[V�Cv2
�-�N�ܒV���S�S����0�~{�L��n��P��xv���f�A]�˹ER	}��������Úc�m�VJ4�:�(S6�ԔMh͹y�DU����(�* Չ1HM5�Vm�:Zu,�L�R���-� �X���f(�ҵ��i����iV��v�V**Y�`V)�Pzko^��-V"�o5k����JƦAfKT�I��	����Xn���2f�cݓ��5�	>N"'�U���RpH���e�66��[C ��T4��o�Bٛ�z�Y��Gh���M�J�p3E��7���"�f,�*aa��IB�Ky�8��JS���Ay�em��c�ͶQ�n�%	h�vb���ǿ
�,Se&U�Wn�n](�[tܹW���s+n8mU�t�����p3�7�4h��t5K��?������G���6(�V�F"N�l��Z̼x��+��X��D�Gi:���XnI�aP4t^�������
Q=�2�)���a[&����SV�T���3]]X"`u�Z�E	�md�l���ږNR
:ט�X0%������ݑVT1,���ܤ�47N0�ǻ�E��X��1`svk ;�����[�6�[ܬ�n<J1���{F�vǡ���\�-<VcR�������k����- $��ź 80g�*�a
�Ե�$�@b�!�!�IAV�ˣI
E�7�],��&V|Nj@�F%SpZ���Pf��CM��j�E����[/Az��vt�ǸP��c�F�kA�pm��j�ȴ]�x�u���݉�Эd˔�ɉ�܆�paߵ�Jf�����Ԁ���.=D*���k
Nꠊ�w5^�Uح!,lW��G1m�'wݯ6?�8�O9��[�||Q�6��-=Vm��S�Ya�F� hC�u ()��lh�bR���pX����^�-�e�kNZZ�W�t9�{��ℙ�kix���H7���-`Yd����U�+XE`�Rnn�1�J�-9�ʃ6�֡��6���c�5p%�vy(t��ss	��ǔ���]�F�̦�eM!Ϧ���˫1]��ݰ�Zw��"�%����ƍ�Wf�� a��*�/�ފs-�n՛�a�j`��;�RB���
�]�v�wo�V��n#��'۷)�6� ���[��JX���BSaݜ`�j�80a�{X���M����El���SUɵ� kǖEi��O����*�/o�w]��w�t�� ��6� M�R�=�0�+r��km��x�ϲ,��R=����r�=��yZ`1"+4����X6�^e1���m��Vg�d���Ќ��@4�ӭ���`T��f���2�Z3�jcZ��եW�Ihڔ����-f��wVd,Zɘ��K*��R�*nі)8��"�>�����Z&ŷn��P*Ke%2�y�j�7n���@LD,3W0)�0L� E�d�K4I�%�ݻ��V�0/7h�I���o\��Y�Q�����S�$���;xq�j��b�� �DRj]���yod���%�e�2�G�M*$�F��n�" Ɠ5�n�+F�Uzc(�������&�S�9nk�,�]���@/  �`Ф� W;���l���-�.���H��%��F�<.�br�w�+����!ljW�j �uFM��V/Ey-
�"CQ@�m5J5�4�gw4l�vZV�6_ڊҁ�Q�f�ڙb�NáW�@�M�2�ϲ��2:���ܛ���x���?4�2�E2�6�M�)�7�ӡb9b�;p�z�H,�V�Xdn
���t�gU��nM�v! H�Õj���c�[�*|��U���C ͂��NM�9kEC#J�a��5,O�`[Wy,EOq�Q!N��~�u)iHJ-Ʀ55;�yx�T��r���u�H�@WO\��j�Ь�Rf+I˰Z2LM�˴�/��!�zY�R��ԥ�7,D7/uC�!����U��Cu� 3a�
����T��m��"{8I����V�W��CQb�i���ŕ/s$i���k�tI�[��6��)Ҽ-�{!sJGFU��H��UXv�Ȯ����lY�^&c;v4��R��*���Z�[I�]"n�^n�=�5[�
w�c�M'bl�w3�իmԵ@V�[��e%(��d��.II��/Y�F+<6ot�(���)�+L��̲���X�7 ���;J@D3{E��]���f�%r"�Z�Ғ����ᩔ���N6F�-ˋ ���Cnʶs#&�|FG[6�u��մ�����ae 5�+U�ɮ�n:W���s�L�L��"NK�vP��ܽ��.��R�L�%k��7M��K��"�ܑ��lv<VF��˭�Bf����k�������.�U�]�vFJ��0� ���d�vvf���	��}�.�U��K��z@�"�A^S�r��h.��,[Z��̣yR������QFb���Թ0hP��ҩ^�5�]0�
tqۧ�r�S��Tj�P�,���Ő��vB6VBk���.&���ɹ_A@{J1�Ǳ${�Gkt�f
;)��T�bMr��n!l%�Qyb��/U8�Ֆ5��G��v�L�%@��X����*мć���-ܱ�B8iհ#RMe�����H��"5X�tŭ�@�u�TQP7C��Bf�:)��h_D�w��ܰ���V�kwYP!*�%�:g>q���g%�q�*�y'ț�fӭ��G�+B̦hbL�1@���ʛ6#r�j��*�l���	��
X���e�'(f�TH�Փ\�Y�-��fa9E�&j��&E���ڷt��6~�0�ed�4ԥ6�^��wZ���U��[1��m޶N�i�J�-��j�V�fΤ��4$
h���UnY����i*�3*�C�`
���$��ԋ6r:���х�֭<��F�Ӛ����Z	�
����#h�D�[���G+-�I#X���0����JҶ��V^�QQ.���߅^nB�d���D֋p���AI����i^�wK�p�e衴�ˢ$�+R��H;��J��Q�Lf��_�+͘���Z���v��+*b�d�����l��Z��bH%�.�m��O�ź��p�9&ښro��K1��3�{�`,][�V�y�hrݷJ� �V+f�+(IRT�YQ�1Lf�sJ˖�?-��x�Տ�Aa�PI�,�k͊G	&�Q5��y�EZ;�n)��n�B��ܰ�έ	Rm�^�4��;h1���������Yj-g0k�1�vR%Uթx� �fFif�˩2`-���Kʎ�#�g̪�;��N�CR�N��znY�2�D6,�Ɩ:.���u�$�kSVv3Ux��A�$���Ei��@bvM@wu�m��f`��53.9z� �
��A�!(�^�>ֱ�L�;x���kcQQ ���X4���3Su�@�]WBC��q��/j�G$�I���C�h{f��ZW@�&iY�$W0�wv�z�c���F�#
	��� ��.�j�ՂB���BJ%	gu�2I%mǷs%���ت�x(/�L-��*��wu������A�vR�n��-�$��Ӵ��N�,4$��[+M��`�35h����q�1�U70����@���;[{.���T���93E����8�5x�f�ij�e�+2Q��I�LON3R»�AˬJ��R��n#&��hV�mnX��-�`�0�$ڭJ���ƨ2���K]j�3h<@���h A���%�2F����w�w�J�
Dڱ��,K#�F3O3V#�Z���Zf=�sIHЬ�bC�İ6����9�۰(�r�V&���r�ɛ�"�+
%զ��t�M�S*�?�/<�{�5yǭ�}�O���"�L�ɔ�n,�YGC���v�-7n�A\r�9(B�����J�r���uz��U�5Y�Z��b ��ν̅�� ��^2��WI�[[�iz�5%�7t�mn�A Y9�u����8 .�%j���f�o+�4�#T�.�p��������w*�T2VQSYK4C��$C�Q
�-���p�Ij��/X�����{W6R�$d�%0��f�ilrS�$84^U�c�F�˽n�
��
N��y�	����Z�Q��<������e%���離����HH �ފ2��۟jׯM:�i�!J�ӡ�r��M[�X�Jv�=Fd��(K�����X���7�$.��&[�Yx�$��v�w�����,�yX��n��MR<B46�����0�7�S��Ja�+3+T�ͤ���\���ƴ�KT�̗\ғ�m�0�Y��Aچˆ����R�2��{��ir�r������-�Y`�-.���1LkI�9yV�4�4.������S^�wJęA��n�u��Jn�(M�:E�[F��"�V��۟�%��L�^��`@(�7r 6��Ą�xP�F�`l+x�}��R�C^�AE�����"l��(7M]��M��h0uqWсoG<���u(^#n��\+��5���;1�6q7�iq�V�Ƌd�8<jR'��{�-pA:xǅ5���_�4/�v��5%��4�$��*R�k���2��f�h��1�±�]���`�Z��DHZb��Tє��bݭJ�0e�&��-�2�[�$˷A��t��ZT���T)�LqY]�t���z���XZFB~qTn�G�Utw
�5{��5��ְ��SjޜOKb"��ޡq*3hlU�)��T1kfB݂4�m�iv�]� s\�7E�-�FݷW�Ӱ�1����*��h�)�^�6�B%��ܸN`A�oj9-���]�ڬi��&"A��G�3&T�R���ux�E���J!�"�@ҙ�҅�-�A#�쥛��)f�eL+@��.�קOh����Blr�`������e,�@Y���kn��K�ZP6ȭ��YHC�3a�"��%���Z��z�b��1�L�m��6��ZX�j�H<{�yv�`Xq�"�o&hZ 7i��JSS,fZtS:�r�m�U��1Lyz�f��"6u����ޡvl[++��EK�� f���B��.̠�b�Q�M��p�vh&*�$�!���;�yT-4$V�(
�V!����fb����g]`�8��%��̞�Ҹja2X��0���l�8��jjU�2Zb\�/�J�5�Vu�6C��8�=�V$�'���GDZֺK��g��]�C4�\�×u�^�����Y�4԰`t�ͱscr^�p��Y��f7xD�մ��[v��6{�f��1��SCa�<����*Ҭ�ݽ��Ԋ(�]��n�>��n^3��E����f���D�^l�]�y�4�
��za�uTKYH����Di��ڽ,��%F��I��M���V��,V*/F�D� ���)��aJ����Q���(驘��إ{���K$!
�V�x[r� ���V�9�˽ᅄY��4�r�W���-e�M`��N����U�ߡ%SwE��j�3��*�"�
.vλ�T�!M�[L\*�i;�.�	�y����Z۽t-CN��bn�Ȥ���$n��0A�@,<�\.,��I�^��!/J5M��o,T�R�\��.V��ټ�&�V<ǧ��Q�9��G\@���r7guR��͢�xE ���]~)M}�I��t�7�6�O��ìe�:4�ڥ�
�Ut�(=T��d՚�*JJ�+sP�����,e���[�h8	�ج��+UM�J�md�Ʃ4dkt+�"45��Rd%gq��1���aO)��7-V7 ˛Q^���i��ZƹL�q��7U��DFya�+%aJ��ۙi=���Z�R�5�0+Y��)�^kX{r�Ͷ��n�Sx05F��Z�	��Y���`ъC6���n�Nõ�)��8S(�(<����1�J�tB	���T�@���2�n܂݌��u��d�t���dʁM�v��V u�MYP�ܨkmm���p�ww�I5i2�=��=��75�=YkfEx�n��U�v����F0oi��"��C�w�f"���գ��B�
cr���S��PJ��& �\ik[�t�`@=Hu!�i϶��c�����h�����P��DE{�m�-7j�ԫF^,ni�A7�"��me�x�u^?����ҕyX�kGq��Hz��ؙ���.��bd��Q�ܸ)ոF(=�j#�w{Xڂ�&��x���N �jŗgR��[���RF�ӡ����ֆ�a����wM���/I���zu�b��&t�k�g��pN�z�7�|j�*�on�ب��#8*�X�s+�sJ�E������%� ���r�������;۷��ꂮ���_.w/�{��y`�g��d|���様���}n{�h���6�4۔�*�.�
���V,lO�	j4��?s�c�|Y�m�]:S���\"\�8�Yܲ��
�vǒ�U-�x���4�whn��3ٳT^T�|՞����F5�v��|v�w�I��F�:L�颫��^kE�S,��>��'�|�ˮ��^�:[�m4n�w%�vȴ�;�nMlk���m���e�t86���Bv
e��1p�1i����t0u+�Y�nkl.o3�S:���mG5X5 �T|�j��@�7i+j-o�����h��h�.8`�u��IC�ŚSumr��F�	w���v�\�S��£�ڄ2���H����%��S��-�
ە�S���_�x&��ZI������m[]I3�[���ƾ�N�K�=b�tʊ���Pe���Р(9���g$�ح�����Z�ʬ�����y�밇�b>�q�i�Z�����5��hM���5���S�=(������|U��Z�<1�þ2�Ѵ�Zc0�8Ng��uv]��&"�Ґ1���XoM�Y�i�3�����r�v9��g��j]{pQaxW
�q˽�yջ32v�\a��H{^i��xe(�!�w��Әy�`ھ�y%sc$ۥyn�ٙ���Na�YapM�s��k���uɛy�/D
����F�;������`���i�aFS��xڲt�Py����
;۞��I��+�n7�Ū���њb��l`�^��m�	��O�j+�X^vldՀv�X�����L�|�9�W�.?<Q����b'�n�|�r������[ٛ�-�^CD�[�3tp��DԁN��*�tFM�1�;�wCV��uZ���4,����]�7��]��,��K�6k�D���\�X6�]�D:噎���i� ٙK�r:�} a��/����sٙ|���1�7���;F�[8b�*䄻�ݨ>�A�XY�9v,Zi�k ��/�-�V*��h�y{�*�.�˴���ބ�D�N$ҭ����-�����I�i�1�8Hc��lP�`z�6���+�U��u6NR���1:�"�՝:�H�v�go��A4�Ӡ4�0�)�wj��|������v��Ρ3o��hV��s[�,����E���T�S.�U�l����t#�+� �)m�Cw����w���|5ׯ�خr�/*և,'��
������#����;Z�#+-*[�X��Z�0;�JK�hu�������¹����\���[7R7EF��1P���P��b�U�-�F��Uu-=q[�͝�EW���5u־
��vR�a�^O�9Z8s��ݠ��6���o�V�#�iogp�!��}�:�{���f6�f�!�,��#d�"��t=B��y���Y8O�{搋>�3����������d���a�6]F%���Zo�<��&u����7&e78�|{*^������w�V��xd��ͮ^��U!g�Z&�
���XRޔ�c���}=��eѵD�� �u觰)�A������1�Gh��<�j�/�
6��ҏ���^�"(����O���4"���ݾ��lB�n�;�)�z"w�RʎP�B�5�E˧�sn�o�7��;���&L����`'�msv�}���JAoi�(�ҙ��l��zO��tH�
�F�w� _)�-�y�&{s�):=æ{�ই��&��J��3�Ƭ^ܭ5O}��A]K����J4R��ǆedË�H,���ps��5�e��إe1=sPC���|�y�&^w��b��s�͇�{([�l���e2Ȓ�k_N�y�m��R[�۽�"�\0�qB%�M����#�j�7i�];p��
t,u���C�Р�.av�"�㘡Bb�']:�d�o5�ej������B�@�4�(��p��u��&���V�m��tbڴp�Iދ���zFN�,ᴎ�ٗ�h�z镠�I 2*�I>ە�[]�c�&��6��rh�y{)�J3^������͢��b
8��+��J�q�7¶dz�e�"8��@�(����=B�=����}At�n����̾0\fl�5�':���sq$��h]Nj[YL�Î,�Rw�c��n�֤���s�ކ3���>h�2�ϖ���[�x4��+�}��k'o����d�]���]2��7�s�Ż׼e
��6��[5������KN���E�<�[��i��,<��P�9�f]�V: ,�YyY�k�ܮ�"��<(�Rk3c�{%u��J!�]˺�(��i`+N��	�,�Y�;2�xt'�]�����
=�[_#mӮG���l���xݠ�yR�XDA���]�i-Q���돦�q^�ކba��+7�T'k��l�4ɇ6f��A(�i��A�9���"ˏ;�5�8Y��\Шr��)���g
���u�o�����{KC�V4^�WL.�,�φ�̄���r�lMkj��빻�u���$fU�4Jڼ���7č	g%S5�],3��;AYx�����&��;��M溊m�G�P�XF�omj����&^����s=w�O��:Ѷ�ۗ�VlS��6&|T�a{��}�W16�ו$n���{	�q<�KJo������v�769kN]��;Y9���bL�$���S��a�5�ƊOe�iz�䴍����ʀ�^j����t�i�o��.@����}�G.���X{�3h=F&&U�V���$���u/��T�].0LٯJ�3���g,�[�V��*v��c�Bu��>0��xQƽ+�f�I�x�<��r�r	7�I�v�hAy���ΔpTp;p��\�pL^��%����sop�!L�Q�lY��S[�9�8�$��힢5�$a>�5uLAV��r{F�5��Ұ��� ;���v��9kU� Xy���ż��M��n¼�Eh,��~�p<<ftZ N�5��Nk�ڄ�Z��A�T�f�X�GH�'Wb��s��4\�nf:-.�Q'x�Xx1F5��,���ǣ6�v��@��Q�Ь}��X.f�(AX��|`�>�m���1�JL}��0՞�B��6�����y��9�ū�D�N�\%�*���+�l�r[TYNm<�l��GrЧc]t[��,:}�
/:�1���9K(ބ1�@�RS�Wq��l�]�{a�E��m�үp�[wl����Բ}�	�kj*U�
\�VGK�f����+���Z�y{�3�����/�:��lF�k�q�*��nt�)���a������G<��љ�ތ�%�>��ߎ�"�����8�6n�ԙ����z�I:ҁ�8b>�7q��W��&w8$�x��i��5c3�N0ڡ��D�4�����L4K��{������07�Ľa��W�u��ޫ}�ǵ.BR%I=\n4��޺�c4�*h@��s�c���7�,�W��J�u`� ��\S��(q+w�@q��[�ֻ0��9eb0't�/	"��H�{�ᝌUӬ��q�&�@q�3K����5�K����)�uص��f�1�@�i`ӻ�q}ʜ�<����΃/��@�4*V&a4os�k-C�3�s��i���r�}e1S������/W��1�/_75G�l��L�+����p0�]Y�?�U��cK��8汅d+�sw�op��=j��w����[z��
�j������r�X�.!NW�I�\W;���L$x�©��/�}޷�����\겯*q�!�`ٸ��Z�6��������A��}���]�|���`��i�DnS�c�8$�V�����9����V�>m)���Q��}=����3�d�>Y�D�s~JWK{��Zd��|������I7���f�wI_���Π��<-���6��q��a�v��m����²�p��`�ޠ�0fOv��dPZV{X��
�0܇z�j\�ӈL�΅	\.�� od�W�jz8�g[|F���ч��YJR��o���m�� 5��o��q��f�ض.�EX���L������To#���֏�E��Y�ژ�����`�%r�34�Kp��""�/���ȴ����v�f Px^;s�L�gp4��P�Z�ʷբ\�ܦ�^�scN��}���Ŷ���vȾ�>4��8��	�Is�gp��y�|�+�	�8�k�+��S��ը^z݁�emX���z����d�B^n]�`��{3Ev��5�O��|5�O�����C?{�f7c�K(��2t�J��f��u��QＺՖ�]�5$g2{;�M1�xA�fe�!ȶ>��*;��-��v)����c�<����e�t=B�UI�q�:�)�+^S�u�P�U�.���$fI����+�f������a�}8"�N/I��+FLK/]�����G��`y_�z[l�ӵ��OGW��o_Ґ����{�
'@N�q��FP�ȫ��v�d��ܭ"n���u*�x�}�j�2E�6�^92���3�(F��كE�65.�&fli5���W�zy{CɹCۯH7J [�]z9&�#n���1m��(��Ok����q]�1��.�bH�r�pS(�*Zv��^�+���.<cw���$3�3�e����ˑ�{X��;}��?)�Uy��Rhc�2K�f^w��H.�aY����h��,��C�E	xn�)�-8��quy���\;~��(���m���E�]*�����$Y�W�a����*�� 8��PT4,��V�R���v���g� ܣ�N�{�]���R,f}T�ݗ'��f�7�rl�w���>}��j�����M�/*t 1�v���zﰫ��d^����p�P����V&���_..�L�-'A���4��-��{ס�m���I�a���''RhG�۱7���xWM(����tZ����|����G�'��-�-��^�fOr}�-<�\�Y8�}���є��v
i<�o�]�5�Z�A� �ʲ��b�<�b���Ye�	g�X��\v�ѣ�D����-�]aS�zr�17�:��q���0p|�^i"�J��N(Sa�h%�U��g���2,�u(4v��ɵc�X&B�h��2����N��n��>�o��z�b(����!����:�}ʉ'�ݱ�dF�U�i�����<:xw��(#>Ӱ������.=W�Q����]:�i��)�us��P����B��o/;([��J���,���_!��+����b��V�]�wB�u��wӉ�fwLlJu8�/�<wb�s��w�䕔VʃBڔ�KI�'Vu���9�{Ņ"堣��u=���P9�ݮ�c	HSo�a��1����(h��;��,�r�Ж�4�#�w�fJ<���I���<���+�D�}FP�+���*(e�5*�j��ok-���/rYMoZ�R&��/�&�2ļ��ףc�F�*�]�Uk��R��=�T�ȵ�i���+���cx2�9�,0m�t����d6�������o�g_����x<i�x�\�J�GSWR�� 3p����]�h�����h5e8���P�9����}�Ҫ�X�$<j��eA�W.�Vm�ϋ���<��h�v���n�eh!Aca�8���Ӳ����\љ4ֽ�A+v�c�s{J ��6P$#��A�W%��������ן��"�v� j�e>����]�6z@��N�f�
	nb[�����{�Y�r��Ő�F�0b��3Q�N:�w�)�͜�mk�a�Yq��v�2��3B���i��D�?��b���tm�B����fL��}�b1}�r!{�ʗ܌{�!�[w'�X��P�]Op���|r�B#�u��$e{fH���Ǟw
�ڻp�x3�h9�m��s�7�A��;a����LY�ˮ}�9�T[�'Vwik��޳Y}�{_� �pR	]w�I-���U*����{w[���S����#!B�V��IS۝lP�F����c�߶�뙐��3�*�c�J_:+ᢨw���P�=3:�3K��c$��B_� @x���J�N,ˮ�9YB�[����� 5���!�w���P�R���ќh8v�uׅ�j�PI�I�N����r|f��Z�1n���4��h����oYM�i��V�Ѧ��پ�����v�_KK��2��Qy�8�&�۫b�<�O�]x�k�͏U�g8��.�zoi��w^T�ݬ*�p,�����A��<ͩL�1�.�z�#�kmlH�)���E��o0oj��R3����H0���X�X�/>���:[���>�bu)�VJ�WJ+~�3�Y�W`�Mp���^�ne��n�x5��^ۺX�s|'��_+��Z�����k�=r��E"��v�u�YS�����&&�5��H#�Ӈr�uz�T�����x�QaK���(��6�nէ�f���W&��ـU�6�hٴ�q��mf���0�, �����0��Qֈ��j�B����S.�wܐ������}<2���9]�e�=*�K�Rǋg��A8}��Ʀ$�$�w�8��i��I�N�:����������U��ǯ��Pj���5��.:��]4޽�^��ғR+;Ne�_e��v�Ryz�I��b��w���������
���y�x�}7����ݪm��e⑍`�Ձ&���y�ӫ^����.��[�]�/��i��咻%Z��>�V�~
���8wA�צt�����C)�Iq}2���5�sD�W9]>������  �?��1�󿯜����^q��J���e�^Q��e�>�3��V��L�y���1I�n�r��ӆ�cT��O����i���Ŕ ������F/�i�}��$���}[ y�J��6XW�r�h�K�p�CH�t	5w��s6Q�6n�V��Z���1;�<Z�H���g>��`ܝ������*Km����[b:�:R�X��cu���;��X���Ę7xw�����
�E�uΚ��'J�a�W�L�MXB����t�b�j�'Z��дo��{7]c�)h��`i���J=[���;3kb�ɠ/uf��.H:_mR:_�K�zW�G����ɣ�M���]�T�oCeM4���:pA6��#��V�45k�c��Y7��|yb��[��uBxq���S��^��f�w}Y�`5���B�R6���<�8��*kLs��l�4oM�]��o_iofSF�Cf9Əx9�/)K�vt�ў^!y���HVq�)XkX�ܮ��m
Cr�T�ر$�E`[3%��f�����̓rrO@�ү/o-CK_y��oY��Q1�p�F�lA⎽)�MNu�����VN��5#���Vs#+�V@��'cW8�CKՈ�]�d:9�"����%]K���@,�Б�w=�7x���L�����1�u�H&<9g����kF���P����(�䛕�1���YP���I��MX�l�P]՛p������(��䕋]|Q]��@�@�O6�绛�+�&���݁��܏3�M�{g���̇E	���d�F��|�wt|����Q�̽۷�����#a��/t�x�)���[�QT=��#��k���%��
�ӻ�W����vx,��g�lj���,7����5vU�7�,�h����n����A�
k�v�yW%Y{��D�]��c:��wPBԹi����# $A���b��ZR��U�k�4�L=�*Ewi��=|�>kn�9�S�����Ns�L��0���=��K�lܡ\o^M�����j��N��Βd5}�B͎����\��2D;ar׬��Wu꾍�8���Ƶ��Mp��W�	oPiP}�Ӵ�&�Kԕ�n��g ��4吖>l.��ZK������-�xj��6�D�����DV��T��3�H��X��1e�����=��^ɳ�N՚������y�r�0H�KW��/�/2a삵�.��&�o�n�X���b���	�Q�Y��SI����,Yf�tOd�U&��ě#��y��LS �)\����7�'3M�y�1��1n���6�7.�Y&f+�t�j|�1NZMüo�D�Ą�s',d�̎�D��T���ST�]�h�8���GFh�L�}�v/�$ﻫhn%�uڡÅ�TDN�ۺ�]���c�`�`.��3��pѽ��&��AY�*��֢��ߤs��Xl�l��Q۸�$��qfە�s����)IgV��������A��p �o{�*���Y��osP�`�ک˧Ռ��|u)~�6���'��zi�V�!?���E�S�K�o�@�n�Z$`�K�K��C���� 7�c'aG.;G��v;�Vfٮ-�;H�M�cR�3�&wT8E��>�&ظ�+^���ڛ}�	���x8{�H�z��:�۩{��W��>RlsH�;��l�P�,�<w����r�u�qV��.����U�U�Y�'�/vS�Щ��d�t�b��۶��n֭���&,�+�1* (^�ԱpKv]?&|��qhv{ك��e'��N��m[l���S�/續�i]v웻f����C!�_v^�k)f9W��]t�߯�Lut�"��n���&��� 7ӗ���Vu���(�
����@���j�Ez{�a8z��3����#�a�禼u(f�1������K�����3y1����8'�ծ����U�`����Uն(nk��ώy <R����튃��g��T7�.�ˇ)��< 8h�d;���N�x���}+�b��͗�{2y�hl]���[XDX!� �d�{��E���t�#�תP1��)�7�����!5�H-�Ew�e�e��=*��@EXuܼ,���)���!�h��S[�"�|2g�1���>�{�H�i͉�f�/����N��s*�W����$�b�B`�<����'7O�9�1x)���W�t۵)91-����K��׍4�Öུ6������pmi��A)V���CH��gx��rel=���S�}ikY�wy3e-u�j� ]�{2�����k���ˉ�$v���:����v��`ɢ�pw(^1�.�,m�����5�sW�8�Ѿ�Ƈ��`���E�aK�.EÙ�.>�\%Y�+�����볯^�ԡ�0�$)��tdͧ\�&�?-y�|������I��O%�ۣ�e�y�RG�x)=�\�8�9��B%:���>�!��4l� x/ںͩ��֠�]G]7/)Ȱݱ��`m���n��4d2uͅ�Lf��e�b�B�Ӏ:"n�Ǹy�v"V�w�>nU�<�m�]l�4矘��*`5:�B�1����t�b8��f���������J�޹�����2\]��h��sSJ�Aո�w|��HVz-sڷh�L���^��
�s��뇻����*��h��M���"�9ș� �,\�&=��Ez�j�S;'�T�B������x
@p�Tֻ��X��m^�D����9�"GH���`�{���r�]Ӧ�w�V�4�<j�W���@�ˌ��i؋V�h^v��T�e�̻�^t-_CF��z���*��:��YY9�����6J6���4rI�!�h+L�{s�����w��f@�-��ŐD�!��z�m�z�.���C�N҇0��f���<�+xv톣D�3�����=�Z�� ����Ҽ�ӊ���o���]���Y�٧�'*GQ�A����w�.f,\�C�)w;� ���5��_[�콑���.�7,��b>d��S��X��Ef�8���n.�v[���@�i��2����75�e�l�%�ƬӹU3;�F�M�	c'`VC�ψ��p��Hiܸ�n���:��p�K��;ץ�B�f[�$b�q�3�6Wo�Mt(R��;���Ƒ
X�9>G�qh�W4�=�.���ë	����	��XZut�(v�GSa���԰��P���|1�EDq�w�"l�h�)J�̃��{���%[<�B�9]0��&�HP�E1�L�{k���O�A���t��`��.���|���X]�y� �4�w�f��R�vn���:��wFC�kZ�L֪5�P%���n�~�Ge�5��+�D![��秧Y�0iI;�֭��k���Yف.�@�G�R�{D��R��E��u�sL���"B��s:�Yƹ�o�h*�r[�C�F4DW��֯2hU˺�Ś��vH%�ڇx�G��}�fp�w� �T��59tͷ�yM��)�u���ǼVm��ȳO9A���1�Y�v�GL�V���0����Y��P�Lyi3�Z���n���ؓ�cUL.�*׏ۈ�t2�$��;�Y��!��KGs�9�x�,�#�֩Ǜkb��ә٪���"iMe�]��̘���w2V�]��޸�L�l\�'qq��OiXq�[z��N�\(rL��M�H�����E%�*g|���FK��9�3��'D�s[�;�u%�<�t���7h�V-��'+�5ǹ��[��)��Ѷ�b���|6�>=W������#b�Xw�͌_�!	�z/�ԋ����2����^�ݽ��ڛf��Lz�D�-R,�k���k4�T�`z�������83����}��'�{����f�n�(��<�M�\#�e�Ej wV���΂������g�BŸXX�%X>%���x�X���ib�L���	[[vi�l�X��9��d�m9(B�r�p�p��W�tM����έ�ܸ����7�u�g7$����ͫE��{;>'(M�z�hn��[�B׶���%�<����g)�2����9�=�<7�o�W&�.��Ο�~2b�"�A�VQ����7�e��^E��D5��Q�z�٤��2�3��i$"�3���>���16M�{�&�J|����9���=<Q<ūw�U��锹��:]u��U�sQƮ�h�Ӕ�r�51.�+ǁM��|�v�xG������O�d���8Yy,�4I�[(�݅Vw&��(^�L����NJ5�63p���xs��ǚ�A��#^y��4��,ʎ��2�EaӅ��R�*Q��a>��)6<'��.�Q��Ʀ�rXVx�#��c5�����:3ݽ�D;�0�c;�`}6�7����ү���H�g���YBŪh�a,��]��&�����o8�c,��ʺ�ڢiк:�Rb�f�tt�;��N'�O��P�#����tž�,��ŖC';��鞆�i�w�8K��^��H<r�L��:b�#��n�e�V�w)�J]��%�LDEOxd�3�ƺ�R���tٖ�|�[� ���ڕ��:��Ir�':U�S,����z8�NՇ���3H�|�����m�&ׇ������kS0�J�`�������o�0^�Q��&h��Ɋ��m�ڵ,�Z�/<7Ѓ5�O�2w�M�t˔H��K�iP�u�n��(fj��r^]hL\�n{�}^��v�ߏ�eAN;����m�I�ys-�w�n�F����(̱�_ �W�XEjVS�ά��Jf�9�;N.�&�N�+��� ��x@�spF��ܽ1i;dn1�G��b �^t^�+W5��j����b����Q�C�Bh=SA5��8�|  ˺y��r���.�i�~����c��s�?<��ఄ���29i���υa��͇*��d�4,e&�ink�E��E�BY�dH��n��ە�ud�lQ;0y�f����{�޾�ܫ��i��[���ej�6��|��L�\/Gq�q��L��a�X��fr4�{z�y�hX���>@֞4Vݭ���T���v8�/d�7s0�Q�����밫J�h#T�I��D�f5��m��`�'p�[�W}�LW�]ό���I��p���{
�[l�t�6�f�`uI��OA��b�{
z�
�[�ěyW�HJv��sx��OPYZ�у9�P6�=K%_^�}p����k��g��H,��Z[t������ӥ�.�Xi-$��j�:ӛ�Ư"W���íc��ti�ʬT�R�w�2]�`���\��jP���+lRvZ�t��QY���gܶ��p�+/���Z�ne�� G��2��#��=r94� �Yy2��:���E��`�����k��#��p�p[�'[X���P�T�g<�2��x:�ֺ3@R��B�s���=#�c�[A�z>y����3\����e��n��8��ekFda�01ή�-]�4�<|\ Ăxե�4˱on��*��-L�����=FV�v�T.Oo;��9�����1�©�m�7�N�˰&��AM2�B�1}W�6雴��>x���".���3ì�*K=z�\ �׶��$ఒ)��(�-�"�i��v-����nH�$
����:�f������͞�q]Bܬ��C��؅㱚r	��~�sy�FA=��mb{���뱪m��Md	�+ �0�����Gkr��j#���@�T ޵��ҍ.� omL7F��M��^h�͡ϳN桉m��&�tQb���kX�[d*9�أ�9}R�	�@ڥr�%!:��y^^�K�,@[�-�o�L�r�"+H��c�$��C�����z�V�g�2*��ݜ�	��v/8r��u�����]���׬"Y.wv�K�%�W�@g�bL�f��,�*��������'e�� �^�T�]R�)Pgp�ۖ�
gJ	C2��݇�]�OHn�b�:��R�c��Z�\u��E���N�>yw`��!�\8�*6[� J���M���񱷁0�=W]EنԵ.�3H���Wϸ�\\�Jt��26�rw}I��};��B��ʓ��jd��u�] Lr�վF�9�RIq�C���.��?DV\n#d�͡M|���w/7�{d��qxo�\��%�O���.Z����ni�C�F��Wu�4g/Zt/4��IboYO�u�mq�o:��y���l%jWv�ފ�\Ȱ̻�6��=�T.�c<C�|�%=e���f�L�;2g�` �++z�d��/�R���Wi��c�kT�lH�72�7Z�\3����b�k�p�-V&�\6�:��aT��9'��X��z���F��N�w{��sS�!ռ���=:y>���t�uifq����	�h�V-��X��ԕ&X��`7Xn�`�8�Z����v'ڌ匘_7���ź��	눈�L.>���Y���oE��|�*�I�����z��s{������བ�m��e�K�*��냞�N؜�6�I��E�!ځFqˁWq��g�7S.V��R���K�s���D:�D��WUÉ��$|��A�;�����3KU���ykm[7�S��G�wv�5�-YG��,��v<hb�	��H�2Xڽh�'8<��q�/�I��T�M���o)������uo0����}9��;�6��a�pʳJ��b���B���.}��P�h�ɗ�k�8��ss�z�Fe2J�`��Srz�ܐ�۾����FV�ؐ^AR����uIg�T�O,�����ej�R� m��g c� y�p�=�c��m�n�56=-9܀��ܰ��z*���3
�t�<�����M^�������}��>�����[`�e1�zn��M�Ώ>��o4�u0������+���]�Yk�frű�����@5��f�wiv�NT1K�����8G_v(�Mf-C\}'N�TD��h�[3wwN���J[�
��;zc��U���=x��b!�5/&,�$��}�mm��k��B�Ɍ��j2�r����d����i��%�������~�پɶ{�������-iHnަ� ���9�)���A�J2sѷ���}��q̍{�@g�C�z1j��P��^�WB�cM�ۥ}IE�p��&=j'Փ���v���9����8$�`�@9��֑���K$0ffm1ci]��LU����R���MjV�`9�R�V9>5D}�<�KX�T�_@M�rHo͕����ֱ��u]�G-\FH�l]�,Η�t
�A��g�|�{Kh/�,�΂7��������@����02��R�oX��P<�������n�h��n�&c��̥FK����)n�C��c�<jƨ�Η�Cr�6�l➂B��+�ʝ�.�\�t��!��Ov�-�1.��S�{�ę�7w9�+I�8�[��D^ƻ݁�ְ�ks���ɃTb	nl�Q�M#Em;����r�-�۴v����=�^Ws����V���*���~���������>��T�}�����jD�*jeQ�I#.qP����Kf)V�\.P*"���+ �)�hD՛J�e%fj�EeJDӖQ�JZ	%C��Z(hl����E��:���q#�r���3H�DRfk+%4:��CD�4�(�-��,-
"��:Vt�J5(��QZHU(T�%Q�5fG!P��.,�M6ed�[�<�t"����F��P�TU*P����i�h�anp����eIrL�D�Z�+*(��0ԍ,�m38J�b�513�W*AH�I1#@�eR�;�
�l�Hp�ȫ���J$V��������䚆$feaQI�,(�+��Ó"ʄ,+�L�+�$H�8�@P� "� 
���h�w{[�r(&T�Ӽ�g�8P�T̙�
�_=�N�5|iE��gf-&]����<�^ۙ�m��.���������Sb�JĀ�2[��՚�w(*�Jg^��Y/j��\3�^�ė�t!���9�/�i��ր%U����.�#�y�	l}v��wc6Te3��T7	��y�/ܖ����`w^X)��@U���exU�B�8���S��
^�1���!e��,^G~�s*�+�@�~�r���^<(��i��mQ���WӡK�e_e��W���˗^���f�'�-����7T�ˎ)^�a>��ƥW���@���o��s�1�����Ʃ���v�.�vX��k����Yi���ُSޕ���9xٵh*��S�����U�l��/�_S0V���C�/ث®�s�7���uޚ+h4�v;�!]���]CsK�݈�*���q�jC�ľB����0V�	u����J�U	�MU����2��E	��6�c�	����}3Һ}i��׳�*�ze��V8`U�B\铳�}c�1>�.��t���0����e{��k�dJ ���#18{���{EQZ�*E{L. )��櫫�@6�}�~�2ߪ���Z�z�ug�V1��/f����Ⱥ<'�S����M��|����J�8q  �Ρ��׮J�K`�{�	��>������#	'[��dS;,^@/��S��{x"�ۓ���#�}�k�7E�1��J�b&��DE��
6��a̔on��c��sǉ�7wگ*�MW��k�����S�M���p�^�C;�2T���ż�݋�l�̣��/gv�g��>l�����[hX>P_,6���c��R���*$c _^|�����қ��I�B򖛓��E1��ª�'�(#�~��rb��}��ƼfY ײN�����-7t�d�e��~���9�Cǆ�����,|k&/�w�aP���������P\|����eKc�����w��$���4;� v��²��C��[�B�_%�;l���c.F3�ч���ʠ�Tyh�1t=^���G�x[J�aJ�Cbr�u�o�,n)=��Ϩ䷃�~ߢd�#ʷ���n/��#���fj	p�}�ϊ�4j/G������pO��8�h�|��>$>�@bQ�a�VpK���ov��w'�>�TЏ5��"�^�*����T=�c�Ƥ�W��H7	>��"��j�u��;����t-�D��=x��5�M� ���"=K��K̬%9/s��
��������qqC��(Sp�i�"}��>=̲-`��#��A�NXu�.e���(M�ݾ�\/X��1�"5춆���6v�̽�0�|��v���pR��=<��FIڏXC�m,�ڬ��qkđ��R���[�[-y�Vj���V�4k�oa�9����9�c�k	�F_�G�ǖU�M0VX�����,b<#�'g�����i�ֻn��[�\���������ߌ��x?���׼����܀�u�=���w��`�i�
�J9qU�\%H����W�W�qB��v�;����B"�u�}��L�Th��Y]a��Us3����^�27�^��	�a�-*��\7׏��| �d�p�h��쾱1��\�z���������l��sU]��ҁ]�S�x��h9�u�9V�\���G����F߷�=�N�sv��X��D�ڼBw!��=P	�邆��$ܟiiXwV�g�t��ڦ�=;���f��GQ��C��q���9)�(i���\7�!��厓�s�v�o��ޗ�[��"��b�J���⮔��
�Õ��*�@Azܤ�����8�M��@��jv.a�'������yUt�to���m.�8)�f��w�����b�c�M�|"t����\�\
{.��}ւਞ7�����Dr.+R:]�D������2��ս�^�a������yݙ��
nC\�/f���&B	t8s��r���OU��7�W�*��f]�g^�~O��}��wˆe�\-�k¼�}�/�r�b�ػ�B|՚�e1�S"Z�X�,��Mq7C��q��(�[�~O��ug�y:����X\V
a�oy����v�x/f`��hhk��	8pk�ywu�`�!���7�Y])=�t���ew��w��e��%gk�O{#���.�����5�E	�\���٢9Պ��2�qN���"��D���>KN[9|���fó&���5�"�w>Ԥ�Q�J�X�e� k�@�n�[�r�xW/��þ�ٮ�0mۣ�� ��{T>(�4l'yc2ͺ�U�~����QU���b��.���u�t����<��=J���v�e։蟏	W��uz��b#ו{88��5�{��j���m[PCB����l�f��:n1ĳ�5V+bU�]g����ϯ�
�U��^g:�`ġ��LS���g���^lb/s͸��"�`�Gy�vK��8�|�8��0�KTB}B��g����"��j�s쳙%��-�{�
^�}r�v�Xf��'�v�f�UO]R��o)WB��Wv�La�Ǔ
Fʎo����x򡅫=Y��L��t��H��wٖ��F�$m{��N�����Euu�	ł@{��(��g��{{�l��Jڜ[���C���C�S��t)��f��)p(�����V�c�9r�=Y22<(���j-ٙO�T�'�`D�6�����H'b
���nW���Ǐ :�B�.3 �y��h��)N�)b�/q_$2#�{u��$2.cp|v���;*f}�R�`x��YC����[}l=������]�и+�g�:��{�p�A/�����~2i�J���6q���>��Y�6nY'�=���Dyed�E[�EmP��@t��u7"'j�U����:���B�!��ӜV�V����^�l!ь��u�`5o���k��PU³��wZ|^ז��{}@��q�'==t=]�����>����}�r}����Wl�9���}�
a 9��]�~y�3f�t�/Tކx������O�����q?
�-Է�:��SW����Ǝ<^�>��8.�S
�׶��_
S�Z��o���d�CE��i�g��̀����u��0Q���b��ҏ����n#.S�6���O��7L�T!�^B�]/��m����G��� .�v�����P?|��C�s��a����<��w�<�����\�e���X��w�<k�I	��7�W�J�Ǎ�>������9�8�i+K��Q�,�; ��Tn��=�6�7@_p����q%���)��w��[£�M�4y}���|h��2�wG����p`ͭN3R�"�6�]���+��KY��_w%���ۄi��ǻp �=�ސ�����e _�xW3��o+�ֳ�`�(��^�o�v+�v�1/�W����%bέ�����
�:�q�<'��k^�����E'�s��{�^��oɇ^��}�����dp���o����J����a�}z��ޞ]P�8!�0�	�`�Z�ׯ!D5��h#���>e% �^�Jt�����vwc��PHצ���4�g�|�{� �n���3F��CkĚU�w��C]α�B��F/>k%�^�Wz)����õ�;l��/C4�����ш=��['����Wa�f��.�N���|���؅0
��Sh`k��6+G�պ�u`����n��pᛕ��4cĀ�ޞ싺���[ă��~R��Ɵ�f�{�� ��T��^V�����x�E��u.	����g�N>�R���P�a�O-p�������!v���.	�61"�ظ�k��&`*�>C!�ሴ�,�}^��訁�@��y����#�7w\�t��K*��;��r���-�P��H��(��B[��Eo<�B����X�	����2�'a=��X�Ft�|��,)4:M�sS�z,7tW��'�GV�����۸'�'�׮�j���ق��9�>F^;�O������d�Q��4��Wh���]ܕӞp�%�pq����Ig�jĵ2���O*�%����t=�c�b�<L��hޞ�9�����ϰ�z\=���6���o����]jd�Cʝoy��yU�Nj�3J�*pͥ���q��ݜc��Y�mG��p�g֫�]g,:U��S�z؀C�.�6��SNdFZ�NY�L)t���}﫧�P3�=�@��߷�j�:�=�V> *���_om�d��%���'-=R���oX��_%�{�e���4���M�+u���<S��U~�����LC��mEZFr���w��Z����^}iB��h����x��xHU���x�9쒱����i�SylV�E�_�^�f�	��Lo���Vz��8Պ�>Q@v̢æ|��מ�R^�l�꥕��Nb`�̐t�?��C�h�#1Z�"�t5��=kv�[Bڧ�15F�jR9--��A��ip�i�d��p�^t��^'��~�J��=q-l�\e�޼��vz�M�}H�5��|��+����Aw ���{�Kߟ����mK��rS)�b=.ͼ��f�.e�GiF��9��v��0��b�A;]���˷�!��V�Ҿ��Ǵ[�w*�v�+�P�F��v���V�����w�E�`�G�s7��]��#B��ge;͞�X�ͦs7汅S#�rP�E��uDpD�a�yѹ��h/}ݾ�g�Y���8t�.���\���Q�4]㾿��q䖔����ɜ��զ�&���N�~Aݑ�°������x�#HP��58����x9&��Ӧ�=@�����eB0-�b���֮�ɹ� ����7���_=Qq||�`��{���e+�0�5�+���C��ᯕNV�y]x�r��47�}��dw��G'	����fw�ve9z���P�_=�H?��xf]������O�W/1�TDxy��ʏu���R{vU]��Cj��;z7+�Z��7��Y�^OX\f�
��ܙ��0�!Z^]k��m�y����e w��p�[��7�&���'���1J�C5��I�'6ke�N��9�%�br��n���V�nE
�.xb�^�u�ꑯ�֠�6�t�1����fwm�0D,�f�Y;L��#w�H͋*�LVkaT
W��w-�d\�t��t���{��AK�E�ٕx�j���U8�����/e[�&'��`�"��.�ul߂��*��GL�Z����<uG�=�}��xiӄ\��Ev�Xc>��C���)���j���,�����x|72_�k`�y�8���jm����<xU���jC,��{+��x�N��+1fu	�mՅ#���~Ub(���S�}1��Y��	���h[�Ĳ�ԗ���N%1L*��6�]�7�#ƽ�v�����]���x:��z�;���r�LuR�~ĥ���SJ����OZR�X�wg��ϔ��G�f�E�ۯm7�U 㲓��<�H�.�B}B����싢fĪ�m�ͥI�k��*���>�{c���+@�H@5�TϷ����:��/��#ss�.��ц)���l��p$���I�٣Y�9�L?-`v_͡g�rӾ��/ޞ��Oɫq[����wL���j��]=��Uّs'E���4�;*g�P�U�O����b6xO*������S�!�-öl�W��V�k���W*�����򿽨�q����������0�I��JA����s���ԍ�C]3��}�;����v� _h+Z´/��i�ކ'=���z�J��}�F��{���3�*T�^a�k��\)}�É��Hѷ�o����B�-���f=|j 7+޸람~�����;�<�~�}��G���w�k:����h����^��Y�ve�)웹���v�̾寴�u�6F�ˢ��ʯNlo�F�R�����k�c5�+	���ه7"�JU�-�e���s�)��H��՜g��k��>o�M�ѕ#7��j-�4����*�v�A�N�����D:omY��t�eήs�
�ݳf��i���?�2U�~'n���V
C�����oNR�~�U"���;pD/6F����ό��/a��)�`F"�k:� K볾Е0�5��+,f(��JlŦKN͘����ɨ���g,:�|����0��^�l\h��p4�����돻� i�B�[V냇p�AaYw��\����w�y�]��ڻ��A6��{�����������d��cߍ�WRTd�g.�j[%;�G��ݧӒԃ�)oU��=s@���]�i�ׇ�y>�&�0���v�ţ���~ڢ)xo�u\�5�q���[�*j�Y���[Õ��D
k�]yO��(/���k��^��[ۈ�/3B��Pv��ZW��?�5t�dH�kh�{>˄�
J
F5(mr�]��y���5ڷ��'����=�ڎ���r*��<~��Y��R�u���A��}\��Up��a��l��N���
�c\̢�L!$�7m�a\)wݶ��U�T�o�<\+_���l�W`�@�*��}_+W�U��I�������d��&��&���>��9�.�n�65�0�{�:�o�pC��ƾ^�N�.�[�2���y���U����
|S�F��Z�Ʋ���t%�2gP�����uyI�:���f����±_@
oC�{W7�J�ޭV���:re�5C���0�Yu�=�u�j0%\���'V���� 7+W� ���V���Wy�Ի���W�]\U���m�rwS+��(cМ����k�a��р���t��!������볮����Hڏ�j�ðf[s}/��36�+��՜�i��S��z��[���8�.��vQx<�f���#��i[�Z��8>��=s�3q�ɚ�WfT��ȯ=k>�!{$�w�_�����?=��@�4�p���i���e#���R�)�L7�M9�zr�g�jf5��� )��M���i�Y����WCx�@V_���+K/qe%���l�ms �)�ݖ�����}�0e��F��.��R:)�A���m���6h�+	u0��w��;=���5mWsф؃��7X̼/:�\;�G�a��,�;+]O���~��|vhZ��}�Ԟval�b�j��5�7z+��=�5��xE�Q�4a�͚#�E����k�Ԗx�=�D3\�^�r�Ո��h���HE�K��\�K�p��
�2MOs�,�2\gq�����8ǌ�ĭ�����D�%��o���݋���]�*_	�ѷ\��wDг,�8%Z�\��e�+���[�\�!wt��M%o~A���p7F�`��R���7
Y<J]���v5Ǎz����n�2Z���3*���v�� ��Q�i-6���z7��"c��]:�bҟ���V��l�<�o��-��:�a%w��݋��w����=u]��kt��
�kR�ւ��n���0Q���sXirt�]� ���K��"�}6f�25��|5ٮ�M��t�P*�4��6+:�$���p駵z��3'��̣A]�F���jL�c��A)"��Z�S�V�NV�!Ϡ�{k&f����^,0���4��m�Y[2m�7M3����<�$��n*b�(h(k,��TxF�4SR�aᕥ_�2���ܝ���zq"a���+�x$s9�o*OB�!��o�I�V���&M����k2=;����Z�^av*8�<����v��g��š��X<q�it5|�?5�
ي�뺱��t*B��cgs_w�&���ְ�}��û����ú�C��H���~���ή�Ü�TO�}��U�#^H7����Gm��e����f_#o�?:�Y.��c`{�N�����ɨ����<<=~���+	��3$\��$�=�0�3�	��8��es����R�S�� �N����"��ͧ�hZ�k�v�;.$�𫌕C�W{lW!�ڍ��/|<}�D�$��-�*+J�0��t�i���fU�Di"�����ˉ�2�MQP�x�xʹ4��J���MD"�*�J�a-��e�#���JYK�q9
���d�.dG �U]0��Zp��t�NH�j-D�"r��aede��UT$"�ʢ�q�pIR���E(��P��QVeV�ADQ�2(I�GLdE��l"�-B���Us�&UY!�Е��T
���Bq�*����Ԣ�B�9�V�#��I�J*f��"ԲM�e�G
B�H9d�Va�,�:IfRePvl��W�
��A�TsP��.J�Y�	�Jѕ2Q*���ȹeȢ�ʍ�Ts�����U+R���r�7(AW����,15dD��"$�"��a�dp��vR���)E�J
��`hW.fh�dp�#��1�33�QT'(YU��GD�R��Rg �� ��1�a\��M$�O�PAD��$�r���^΢��"��ga�5�B^�˯(Tk�w7�L�;�yΕLV&�;4�[Sp`yƇ�%s�gG+ۿ�~������o�~�i�;L*�kdM�㸛��\����?'���p}g��C��7�~>����OP�������;>]��&�<I<�����<v�5q���M6�8�lݶ��[���ً�~N*oo��o�N��v�׮�Ӵ��}�z��L.�>��1�I�x�hU���<O��ӂx��>!�t��'y�8���C�_��v�U7?�ɛj4�tc�amU[V�Uv�M��?��0�����������:���7�$����n�$���W�|��@v��N;�s��>u`����nА�8��s�v�
%��v�W��W��:=�C��ٸ�]ϳqf�_G����&�<N3�w��<w��9�N'i�\w�~N�x����;뿰������9��v�:w���>�n�>���=뛥wI�ts�HI���v��|��}zݙ��;;��"�Z��x���9���;�ӷ�x�;}x���7�t���'�ۈx�~���n��0���yÿm�>�I��{�]`D޿���ۏ���?k߽hN�{�N�ݡ�����: ��J��{i�R�t�z�I�8�!�a~!�>;�w�������4�N���ѽI��i�X�oP����p����&�st�}{L.��n$�׊���=�;W�3�?���.�1A�FKEt�Ʋ��_ޟ�8'��u�����ߓ�}:��!㸇��u�©����>��8�_�q����ߠ�:M�	8�aՔq닯�q�M��U����x�T�Q�^Z�ӢEc�[:������bC�8�~�z}�÷v� ��+���wJ�]���i��n?|��hq���ߓ�_�v�]�o��lz���®��S��P�}B|q�J��V邪�(��#�)��^��[�߯�8�9������]��u.�[�������������ޡ<O�n||�|M��'�����;���徧I�o���Gq	�v��~��Hx�~������a~�������)���>�K���oߙ�a������矕������~�,��~�����	'n�s����'��~��>&C�Ğ�|�!�a{C�=��8���v��9�;C���~v����N����I�i7�N�#�O��uϏ��>q�4'��:����%n;��/TQl��o�f^��t��~�Iw�bˬ>5}��/7��{�*��v��l�1a��!��'aQ�M�����;�۸���h����/�����Bn�Lz2M�ޓa��9�SfJ��,){����6Y�m��΢Im���|�pq�{�:��פ���;t�o�ߝ������x� w���z�OɽN>�9�X'~C��C������0�|����O�8���z�}q ���oC����xn�]}ӻ3wR��^����O��c��|��m��Gv8������ǈ~w�?@q�}���G��&�<����ߝ���|�ǎ?��9��޷okC����9����K���;y����l�I�BC�9�/�o��:N��i;N��\ߟSqē���N�N;�t�I�B����ߐ}M������Ӽ�c�t�;<M���g�j0�n箃2�I�����v`����\���ć����u�t�]����ۧ��n�;�t�D�ω�u)����s��<C�	$;>X�����ym���v�\8�G�~C����������{1��K����U}�1wS�������4�O�<��$��׾�����	��|ۮ��!�T�?�H�çx�$�Ǌ��L/�u��<N&q�wN�ǩ����<���|��屳�7cq�v�;�]�_���܆�s�~{����=C�߿����ω����'I��'�{�ݠx��O�u�1�qM�w��:q8�<�q��������~;���;H)����=���|�i�"�n���c�O�3p������������:C��������x����7���py���&�BO�@q����}�}��> q'n�>����4��vfN��}�K�'o���3q&�럿����
�+�DAX)��٪B�=���.�����r���?���w¶Sx�������w��w���o�GI��u��ۯm���!���@wgv�z��o3�;3��<�}c�ӯ�.�������N����;w�#�w��z���w��)�aq�;�n�F�L=w���wI�v}��t����~E�<I�~9��7�O[�8~v��3C�@�oK�?����z1��r�X)����3�?������˻y����,o����'����������q��{N��C�u�8�L)ӏ]�>'Hq���|q ���;?Gh$��0�jp���3'`��L�E�Gc[�u�� ��,66gK;��)ɜ����v��i��g���gæ��A	
��Y�\�_�8y���h�̒�`�|��y�Wv���Ir͏�����b����;!�űqξE^:��}�؜�RJ|�3�����ٙp�������������u�G�4��=N7v:v���t��o�q��I�B����w.��	\~x�7�?'��0������ާI�n���}I����/#K#G���g"�O7��_�.O~�������z�w��7?�sމ�t������:M�	�?kϽbN���M��S��3�8�{��=I<v����9�M��ݟ ���\ٓ��F���bژ#���3K����:p{�q�;_��zN���C����]�0����yç�?'�qK��������'��ލ�t�U�=��;N���=��r���5�{p	�o�e��u�gǩ{�87����"�o:I��yN7�x��W�C�x������Ѹ���u��}~�aT��\|OS��ϛ�H}C�������|L.�����8�����v��E�b�*�*�'Q�������>!�{��m�#H.��?:��$��t|����=I�}��+���8�O�,~?A�&������>>8'N���q���븮���[���G���N���`�=�i#s�n��H8�<����n���aO��}M<M�~N8����]����㸘|��������$���t�}}M�7�z�;N��!�~��t���'��?��=}�����?��ƛ�*�@	i�1Sy����"��;���<I?��o|�j�S}B{��޶�v�pH}<��ݳ�~GN�-;�k�n?����aW';���L/�|�d?��8���8np�/�vh����WdS���۬}��9���|L*�����'�>������ߐ���Đ��}���?$��矺'j�S{��ӧk���:�hx�t����>��}v�N��j�@}@_|3�<����rO?��������:L#8$>���O{���O���'�<wHx������T޺C�?����Ă��ϟ=�o�$�������?��çNҽ �n��s�S������]��y�S���u|���?��i�H|N'����:M���R���+��x���_���÷�RA�ܜ����O����}�Rx%]B9���/z��g���V��$+��oOo�8�#u�k�d:�y{��<}��Q�|ug�+p~�+�O��ż{Q{z��,��2��qÂ5|��O�E�U����+}�0�m�=�:t�]}d���4S�ڥ��Aw��G���"�zpO-�K��Pa��W�Ҋ��ӧ5\��,�s2��g�"�a�Ղ�����@� �2Q��y���)9�2^�ʙ��,�� y��V�eoG�]Z���۶i�8=���՘z�l�]x�=핲�1\������˦����P�r�- =�}�>Ֆ0OwO_�NRy�jf�1��(��^P�n����������u�+�J��k���+�s�����i�~�"�0N��O=:�A�i��T�<A�y��'ր�����q?
�/u�r���KA�/�w�7��������gA���j-��׊�# �*�N�Y�eו:}���ɘ0W�,(����
u�X
v��=u�AUo�����
������~�0��3x�%f��{@]f+E�V����<%
˫��E������}��{]*���a�sz�w�ts�u]�U'�}��KU�W��捞�����]T��`����U�W��˷����tW�����|5���k]�Uμ=��or0e��|�<1ռ�8j�P��~�jOYz&�X��0��F p,���`�4�ҍl����m]�3�(�v�m��"<���HT�yh}��yH4��O�Z��ʲ�ì6b�&�"�(�Z.�7�>�I�^4]��Jp7��C���B�C^�} Λ�xz�c5�`�w{���|���S�zϒ8}{�FP	�>R�Y	�������݄p�x��0�3����p�̆�qzh2��g���Z�6����u⥂���d�޶wݺ<����k �/����<,��Z�g�|�u�!� �O��^ɽ;n�[��++�v�׭*�x��s��6���Ӿ<�
_S��|w�}+�/h¦�)h{�M'*�FK;�i��m{a�z�čQ�e���Ϡ� U��WM{]S���`E��,]W��:I�ð��.'��40O�����ׅ4��V�)�(/�y�;�½��X\���bd�������u�o-���	QSn6��z���d\���Ǐ4k����ğ-N��òǺ�;�{�E�����c��2Kш�hY.��HuP��@�	>c�.��]��nv.���|��֔��9z��zc^&UD2$yCޡ�`*��������_vۧ嶻��66a>mW���\�V9�ሱ�ǃ��o�L�jT���5�]Oj�g���y�{�
�"�g_>i�zf�6��g��f��eA�lw��n�2y�t�D�ȗ���z��=�Ca.�ڌӸ�=5.=��sj�`;��^��Žf,���Z
Ffn5lP��Y�h5��]�j>,�JzEuʸ;���&����({hK�G{������O'ϻ�|��&�u��2��q�Q�p�5�������]~����B���+�W�����ba���$+������3�7�6���⁵T�x<�u�2N�q�B��hÈ�݋��路#2��4z� ����#��y"6ɳ�e[�Z$�;g`�ؓXR.7a6k"p{�L����t�ޓ�޽���pV��p��
�/ 07�<��+8n���f��U��2���>�b����W�f�	�ȥ��׳�Y�kI˒�)�=Ѿ�����p��(�;�o�Y�<3�U��=}�n��7�3�	|<��V�����D5r��[�'h���b2��kH�c�En�I0'�g�	iWO��>��Q����ͿT�qx9�^	���0�+�xo&�p�&U��a��UvJ_Jw1{��N���/����C�У'O9�F��mt2�>�2����ut��L
���Ex�CK@�@$3��Z�e���OS�6M��&�M���&�'�J�E���g���:��8][�:UY@w7��5�yx+#����S���tnJ��9X��#��w�%݋�od�u�(�(Q���n���*w3Vz�bO��q�S����Sr���[��M�O_0XZ���v6��'��,�a>|q�0*���L�#����U��ُ�l�o��_`�%�Ώ���Uf�I���vzCs;k�^�Z&�e������^��*��䮩H.uR�i��L7���j�H#F�o���U>U��㰳2źLfv�5����A���4n��׾�Y(ת�����9�K�ȡ5'!���|��2vO��k�l$����\��s��jg���w~5�~��^.�^�t�Ҏ�-a?c�_�xW���ǍP֝fd���ٻݬb�<)����g�� ]{���R���tTz�%�3^J��a9�ؐr�I�������z�ĳR�����	�غQ�(u��R���$W��X�?7�εr�-N֗�fg`NDD�`۲���N �z��)��=%\Ŋ[ �T�
�7��"�Oc�����7�����ָ�;7�/�~��/�IT��_��>}��o'^i�T's���[��6!�U���ֈ�ث�U��U�S��؈������a����ǎ{G&jƏzv���#>���p��ZV9�`�7>J�ˡ��q+�~@W:ć���K
�nU�@V�k�U�5ˣ��Y�:3��%�}��Ɗ񎇲��;����Х���:ɳ�B�!	��{�m�����_�Fg֢��>�r7�.����v�!l��+<����V���{�D� ���:�k��>9��1O�&��N��RuZ�_U}�3Ҽ�=<�������_rߝ�A��鷽��q�T��j�y�J$o�������Ob'v&b�H{E�e��G��
�3%ۧ��s���2+]{�'�v��8����b�j��G�=��s�h�z���N��תX�铂���
�P���=l^�|v��p�C���y����R��3��wL�?--�C��B|u�eQ!�ɶ
{v��H�(�h��wp��޼`���m��Z;��v��JI�K|v���^UZᮦ?��*��zb�t���5�ʣ4�N*�Z`�xV�����t�K�eb����f�8=	��~���5���*�c;�W��<��{w�{,TX9�>����Z���~씳.����^VV�� +֗!��j�m��EV�6��i���dJ�(Q�P�^����@?���ܯ'��J��~T���,�KY�zzl�
��F�hז��͛���$@]n z?-N����ߨ�]J���t�~篳�Z���E�S���%=��?���N��L�{����D���l�N׆�����w�;�}�J��<����7�`�o��GT�/9eI�9�cޛ"Y�<��!�T��U�.D�ڞ�b�ǷcY/�5��BB`�OR'�:�rڗ9�#�v��ɘ�y*�7zhl1���ǆ-\�38�'�n��T[ƚ+����y�����3y�(�ꛍH�;;Ǝ��"��l�j�N+���v1�z�d>U�\��;�?N���kK���x/}=����ۙƮ��3�V�+u��C�< �����E���GC���{�W��n���˻DNs��uߪ�6���G��ް�{�-��L7�,@������ֺ�e��,)!~3�'.�V�2�wa�{=�������|�����<�hL5��������ό¢Z\�wV�Y֜�b��	�[:"�9{�T��>^����J���kL���S�JŃ�=�wi�y1�S���qyZ��i�\�c�DK�r\'(W�����©�!��x�OEJ���iz��3KZ�Q%��:j���\Ck��>2�t�X�J����T[�F�1^i42kм�l��S�3�Z���MW =[���
~68eQ����1���C_���|��l�s3V��ش���2���0�3��(�����m����f�z��Beo��TE\g�id��Ei����l��-'��Ob"�|�}��+�
i՚��H{d�c��ۣ�ﯡ�j�o*pw�<��L
J����p�P���Ϳ>=�*�۳�O�}������ǎro�P��%oYN�O��NX^� d��=[����[{Pbы,ُzNY�N�]n��F��h�aBY�<|$�Y<u>�o��>�ͰlY��M	�S�xm��e~�d��3�6�*q��OFG�P�#+����R�%��L��j�l2��$�'%�6�/8Df`�["�1��~����]�es,�� ���W�����{{� ��;!#�4m�������aW:�����X%��gV�Q(6"��|�Jl��pnգ��k)V�U���/E�<z�<+H�K�ƚu�z������Zl|W�����]���n{�Xw���5�9���p�����0�e�����of������!�>'ey!^�/���'�:r|��Y��9j�8Y�x������-8��� @��w%^��5�$=� ,?pGx�6V�_e>�@��{�N��wtZk|���*����8���>*���S+|r��r�m�e��y���y���te�����E�2����C'��4�C(�ۂY+����^L�����p:s���B�ǔPϛ����c��_i{O]jA�Y��C֌-�f�{�N���e����ND�Ѿ�����/r�C6���xg
t��|6�}�5����!H��t�ѻσO���2�{�e��7�_&�[NC{��ݍ�U�2�\T(��[�ֵ�)��fe*�ͧ����G�-+Ž�r
�e�!9ݦ���g$�զ�d���H��/fJY���z;�":w�3���K�S�4'�C���0�+ch)<x�u���;:nd̜�t�$���
�ُ�%lQI%�asi���Z��{����V�q��ǘǝz5�`=t6���4�P���`3����*e1 �ڞ��J��^W�S{���/ٗ2����ت�$B�k\U��Wy�Z��4�q��H("�2�VT����'����ml"�7���6\�Z�{9Z��S���e�h�a$<�V��>'��۾E���ؽ{�ޥc8Џ7�����;5�s]����wF��C��ޏ�7���z?v]�^4˷e'�>��=�i�n�ϳ�%�X.�ὔA-��.c"��p['��g��4��ՊO�J�S�q���a��8g{&�6�m& ��a�ɽ���_	�B���� ����hG[X��Ѓ�HP��^&�X%�ˋo������.n��ꜻtjp9��H��M.mZ�3څ6l�A�m��4�(hs&AfmoRJ�]b�:�l�c�g&�`>��#�]�7G�����"35��Gs��G}��	zG�o9Kx�]��Uׂ3̟fW+������=)����̺X���8b!>j#��u���Xfe݀�A[��#[5���J�$Ef�,���;Hݴ����ݎ@�q�v2��0\Ki�˒f�ѕ.��l$��ͥ�:d��)�ߔYs�c�t%���G�����ٓ��K�"��#�Sʺ��KEm�d�B�r��Zyi�.XH��8=t���z��KE֠��Ҝ9�.�1zp�̫�@P�9���=�\7��}$-��k-������km܀ھ��'���X@�t�y �Y�F�����i�7܆fPE専�3��1�pE�.����	Q����o�5h����W�ؤ�f}r�Z�R��1�Ws�o!�x�r)�.H<w�[ȷʉ��Q��n�vP��ΰ}}��aV���z�i���8É�f�����OU������a`�����x�=�p�A���99�8Z�+!) .�EZ�4c^����+r#�:Z���ݸ���{�=���YΩ3"�m�<y�ދ�yb�G��0u�S�8vj��tgu'ͭ�(v�`����$L�c�h�'���;F�0)���;�Y��e�c��ɍΉ�X��q���'}��79�:{Njk�5cB���c�v`�)�.��7�V�eLC7 �%N��u��L�#�(�0�8O$�OOK�Uðr��$[���+/I�5���h8�>��(T{�a���p�!��9�c��g��t��Ka�(Q�� C���$QfI���W9�#2�5(�Ib(*�2+�C�(�UEY�Z֙\�e4"
��.W
UV��S�D�B�ȈԩD.p�9j���(�G"���+
J��SRR�r�"�������y\�!UQYA�'"
���,���R9r(�e�(��Ws�y�DQTu9�Q��s���f�(�JՕ�#�1�r(��܂r(�AR&�Ure��(+<N
+�TD*\��,�G ��]ǈ���S"�* ��r�"$�qylY�QmUB��Tu��ET�����")ZU]²��a�L�ʎQ)�Yۜ��(�D˞$��Tʢ��W#q�*�p���#��'(�!ʯ9�ȋ�!�*�]�s\N"���\EN+� ��SYEEȨ�*Qp���Qr5*(�
eEBeDȓ")�*��U2(*�*�*��D\���T ��4(P�W6�F����cV�3�q�Ī�ks�-S�8�)���{�N~\}�8���b5��[7OvV�[��ծm��|>����r��OC����tg �΅uʮxv�6Y��ɮU᾿�����/0�ͅ��q�����{}�KG_���r� N��y�y�����P?.���{6�F�z*m��2�i�����tw��-K*�g:�*��ܿ�����yۯ�ǧ�;����5@�%��s��d���$Ću1�1_�Y[���2����@v(PKU�l�]��e�T�]�
�����uRl��X�R-3LC���~vO�U��s!��h���ؽ�������)����ǘ5\/Z�}j%�_�VW^����t��ׄym���zn4=�*��׏.�����sM���5N�T�D�{N��:c�J�c�U�����^��jW��x��?^E�^�~��C�Z�r����ޟR�����si�+���?+F�
�ʍ�yX�mɵ�<C�j����iy�P�
e�P�
5���<h�X�v��L�gX��}�S��;w�j����E}j��[\/6d!L����<�L�V�nE
_<1{����+��C�Ž����Z�01�p�����v��9���Np,gǢS�s���E���{7Q���т���^�D�x]��Pڦ���zwL�����ư�Y�W��sr�J5��v�0z�KLV�:�o�f��a[�����0�^ۙW(���� |�{|v�)��͹��q��� N`ͻ*�ʵ���w^�r�߶w��7�I��m�g�6p)ğ�R�}k~Ų�S~�ó/��)����T�^�*�x_{� �	h��D��d���qa��þ`��{p�'g�����cC�/g�C7��0D��^I�,)�-=|�{�Z�.�=|�v��]c�Ln��*����E�^��r5�?���J.h�:sH���N؂�ʖ�p���<����.tǃ����4� ��������f4(�(�}н��g�1��
�@��ZT���6kR�.�����w�"ޣVݕ��a	Y��j;Jջ�fK4zE��v+�nX��65���
J��f����-�n������v���6��=�^`f_���>��5�g����Jҭ ���ώ��$��mӘ���7�yge�����;[��&]� [5�<"vW���sh�������������Ӎ�u:ls�Op9��.o�sPf�
k�l��s��7!��c� v��@������!�����5�z3�ӌK^�r'��R�aZ=;{G�y��N����_�ҲK��������]C��lU������\��[$����x���$��Q��eO�$��$����y{|8p���ζ!找I��H\��z���IM�o�Ͼ�����Tq\N�D�F�|���&1��Qn�}H��r���[V��WN¤�]����Hk+���ݽʠ]����|��Q�\���޸람~��z׾�a�o�f_=Oҭ��p���5�z%H*�j��l?�y��mv0+~����L��r
�^0��-Bnѝ=���)'�����*�)X���ΰ���g�7��倮����,����r/�6`���а6*��^��xS�<����Ҽ7�*�8cE�m�H���Fj�T&e�/�L�\Xj� (��+u��C�<'�³||(�fu��^2�;G��=��<T��ٜ�X�j���\�^��b{�=��L7���/~!]M>�Ej��=ʄ�ȯW��ܧ�ӯ �`
�Ok�����<��W�/���V,�C��w���R��6�֜��&k�O�Ƴ��@c�>���[������__�dCW�VS�.VW�fwD��� ��WKK���S`�y�uA P�>���8��V�8ro��tg �c�O�a\�\˷Y�:�y���[��5�b�׀X�^��×Z
;\�G�]ez@���^5�]RP�*dįS����|��O��8Q	���m�y~�?�~�)����i���nfᢣ�w����w<��1�y�~���f�j��YvQ��6w�z�|es���	��T^���̩~:��Ƭw����� ����ݮP������C�wҫh���y�<���Sv���N����������[WY~�N�-���T�Ҥ?z���چw��T��߆�5��D��β ==�w>&Y��:+�V�ަ�{3ݝ��V*d���E�a��]Xo>S��{�7]@q����Te	^/P��zGI�i֙%�ݚF]�'��s%��H#��@4S���u�D?��x��l�R�/s;�����e�
�Y�%���0Xĳj�����.@�&�w�A]�R5�d������}.�-ۺ;�
�i�Q�S��T8m�������aі&U(d�+���-2�"I��#"}���*4��̝9$V�!�"/E��~4��[���$ܮx&���vy�Q���s+����K��������W���F	�m�]�5p�������ܝ�V��]:I"E�lp����̟><<N?y�^�@�~Ў�+͝8qWC=k⸿'�gB��lw:�̬���+\V�ld���TC�FNwq�E��sѹwy[��M6�L�Q��ae�M�>q�&;;Y���p[����Y^������&yc��n��4*��V��.�;���[��zMw�7u9�I�C����O��7��f���d�����0��{.�w7^g����1�+��`�֎~H��{C0����<��ͮe�=�?,�xX�^LuZ�S����>.��^ע�����p�[5�g2z{��YC�o��H�蝞��yT����N���p�]=l�Ⱥddbn��%b���X��ս�mĸ��U���+P��k�LpTE�`-��;d����	� �	F�S�:��ّ	�[��fR=�r�:���58�I��Mpʨ���w���YIt'�
��p��o��f�%�R�iu�^� 3ʯ+�a��UvE��Wv��:;���e���;e�;�d`�k�����]>δJ���7/�8h�2��k� r�%�q��i^5��Oo(ŝ�&�����xU��;S��Tc߶��$_��v�+̱	Ǹ0]�CC�/���8�gwvBg���M!H�{MJ_P�k��|�z%���mujҖ�R��ie���;���	�`�2�R�ؔ&�|�����U
������\��UM��A���	\3�4]��\.\��:İA\)��`]�f��6��"\v��c�Qmլ$�y&qŸ��x͗��٨2���d�<A�c�n��7���e�i��{{����aa飖)���'�5Wx��Yx�M���x�uG�����������;���1�!�f��	7�;�-��v����(M'��|�3.��~0P��C�Z����g��e1Hd�������B�ޟR���%-cڶ�+��5��V�bp�S+�-&L���碋E%�bǐ:.��S�������x����/Ƒ>xT�Ṑ���~�zOq���]��J�g�+�6�4�Z�f$(���,��5E����ft�8�d�eZ*N/����@�v���^W�t"1٩�eS+f��;�jRl��Q;
bꑳB$���3�a�MXz@�n���kº
�_����j������e��&q���f�С ��`�ג,4�P�)�`;^�1D��~T��vV4=�o��o��6��$��+�I����wa�b��[~Z�6�׾`�^j�V�]��x?�W�4��y;��j˺k�-��zq�	�W�ʿ\ᶽ'֌�c�ר.L!�N���"�q�f�,���P�'t�m���pMD�-�̳a
�y((6���oK��t���>�͆���Mrf���wX�H�5�u.���m�@���n�s�:!�Bb��^�v���	C���̦c.�Q-9�Ʋ�)�|��5�y��n#����%�~�Ƭ��zm�9���6�2ؽg�;�Xx��=�2��$u-��x�C�Ms�>��U�U|�u��r�j�9�n�.9���Q^�rƛ�4����2s����O�Z���@s3|Ո^�w˺�\,����A(�֑yph��Y�۩EQ!�ȹ���=E���v��Iu�|�Q�X+e���T���\�����[�o�ʼ$�\6b�����{��6��r�zI�ԃnw=���	���
��ٝ�B�rb*k��PCX��z�U�|_�����^��h��e;R��k�V;�kWl�QȇF(���W�u՚ip�4"7j���tKy|M`��Z)Vx/]�����X ���<�y���jݡ�A5�=�S:�k���|;�g�>�sL׃~c���@۾e���0=����C�ίB�Y~�������K$�fM�w�s]ӳlx[�o�q{
uk��N�|�M�)����&c&�ɺ�(����Cm�kx�#�4ͯ�j��ǅ:~�c6��ܛ�^�E��\�}=[��j�@��}=�oMO5�W��B%U�Իj�puP�	B²ꯗ����|=J�6���.Z1�;j7[�Z���L�f9��q��V��r*�{).�J-��PM>&� �����1�G�,/���5�9�^JZ�=^Y��'Y��{�Ck���JVk�I���/X�p��8Vּw+����d�Jn��*������ۭ�FO�� >����Ij���[·y�w-;�(g|�f���Ǻ��;^h�ȱ���j�-׼��E 2��Gvg�����,z��*g��_���M�C~��u�a��%bΥJXő���Wh��m�/��|�"lk>�N=ώ�@Z�/T�l�^@�<���hI>T�i[n���nIn�iX�z�TΕ�V��5��>�(wJxN�W���є���6��
dV(�3u����kG�q���W;|(�J �i�^��ɭ���1��l:wTY�H�dm�i�{Aa����1��U�O�Ͼ��ԠMW վ<�p�g��$|�Y���㸍���}ƺ��h3д��'��k��$k(�β�f��Ǥ��2VPk�(�o���U��9���Ä�",1��]��(�`�!�ٴ�(��Ø�l��p�r��Ih/��T��^}����m{��{���������7\j����՞�i9��)׮><��E3�`��6%�l�X�K��A@�B�w�H�lV�wV���MP�V\��o0�Gu��l6�������o2_N�j�vU6��{#
���B{��[��kI�0z;�_k�N+f������h^��[��2��L뷙z�^��仱��ɲ2g	�{��3y�c�+ۣ�OQEDǀ�s���R��6�ί����ް�wt��[��}^u�]�f�cQ����`����2U*A&�Z2&��A��"�,x:��~��K�ɢF�c'5=�#�`c�>C�3��48��1���K�g������B��,�0��tY���{���^U��PxLJx��|No��^�+���k��x��	��eM�BU�n����u�����h��熠�Y�8�?  H'�&e��(.02��s���Qx!�Z�N&1nb�nԄС=�d��\Ȧ��hK`,�צ]���{]2�{mR�2�[yJ@�llΐ��86�۱t�d#���cG�D�����ʦrjpy\���<�l���9	ЕP��k��:��j��Y>Y�1��S�#T�ۍ�i�m
����=*��O��'���{�q�7u^��<�1ӭѻ-u�+n	��(���<�`O���*�C��<�{-3[��jӰZ��t*�ș�bU{5��]z/��M͢8�?y��sU]��҆�F���Q�R������2z%���r�V�e�|�Cwz�%{��&E�1��EcY	0Q��a�07%���Z�A�Oi&nP������r���+����ةq㑤���,QXϯ��7��q�V�U��¦�fi�6�k/��ח�u�(uN|���{���5Mn���9]�jP������]*�s��/i˯o@4Of:�G�F
�x���J�Wc&լ;P@�ǁ���Ԡ�CnO�ĩ$_����^X�o>�F���׻[Y�-�s$�ZFd�$�B�q�4�/��i�B�o���Z%�v���J��b�m�"w)��ҹ�~�/��z~ܸC����e5�8;���Ƽ ��-�R�p�ǃ��)��b��\�5ff�C'4����O\��?2�=ٿyT� 4�-:��c@P!�T ���`�T�)�4Ө�����,�0[e+g�4�CY��M9��
�.Ιr��i���<���M\6è�O:S,r)&sM��b�anKC�hs7N��+آ�%�f�j�Z�E�q~���2f�Nϒ�%.u倥u�e`eE
i�uQ�����,��%���Z�.Z�8�,=�)S6��؋�^�ld�D�7�ym��~����[�u�[]��\t��@�]K���gT��nZ���m�y��Ǔ��m���+���Glʻ["k �f��9��&��N���\�ck&��5��eZ�@��ivF)��h��fVճ��V�n��N�_7u�o'h����A�٤[m����o����1d�4�s����ۈA˾7��?=�w�<�%|Xڄ,0蝝z�h�*3����w�qR�7W`�ҁ�8^�C��ʄ�F�Z5���bP{��[blR`%�vr�Fb��:J���VMM�ԓm�.��#�PMxx��j�D�B��kct��=c��$<V���T��^m��	�[7�����8����j6��{�<O5{	�rV���;�hdT0�r�hb�7�]%n>�ر)�����u�(��2�)����Swl�����g���v]�}*휭�<[G�$�A��l'��#��Q�kT]�P��E;Z�+�VU�ۈP��@*��r��oDD����5}�����{]�K�/�A��C����﵋ڔ��^L�~�N1�s�E���{6L��5�@�]ΰ�:Yv"��b�dh�Rx˯N;G�{��{�p29�ܕ��cD+\�N6�,�[nd*t�L�V��S������e��U��,�ØY5��uI�o[w7A1�znӇ�cv��tl�퇄:	�|��'�'�W���n쪞�X��c,�W{sEӸ]�z����F�ӽуr󱭸��ͣx�jI�����a��.�6۷�2��) c"�v��ċ����>�HI�c�C4��*�XE��B8��bu9w}���م�h,177u��J�>����]���`3���e�Z*Բ[N�c�S�!L
]��	k���rK0r��'��:E��w��u���%.��C�.4�n�˝�. [��Y���	��?'�Ϋ����
K�;�s��^
�q��Xn&��*���3�ᴆrޭ~�;��z��XA�W�㻎�̣l����:��4ԣ��P���g:���0�(�;�y�gVu���/zXS)���e�=�b�2�l��5���-�Ė�W�k|r�cP=L|ݎ���K2���B�:v��v:J%W�U]2o[!�B�Ak�d�r\!i�Ow*:}
i鴰l�ʙ�� (m�L��^��0p��V&��.���h�;�ݕ	<4'�>�Sӓ绬r�n1���7{^t�SU@V��
�<V��Qy%8��t.�����O7�6�X��n�N��+�by.��8��c'T]lgmj.��z�t��s���ѕ5��O�J�],�����7ٶ\e�у�1���.h��Gpf^��8pԆ�gf�@�@�}{܇*���r�N�Ռ_.�'C���]�h����ػ�oVUpL8Q�u�w�Hg�9�N��6�w�ױ��$rww?���31�'�QE%Bf��Qʕ
9p�V�D�����t?��C�Tr��$� �W"����I$TD��TEAPr�hQer4���\�f�r�QW�"( �EA��#SP�
���"�T�PfUQEQ��Tp����*�G,�V��Qq$ �����Q"(�gB��*
*�<��2���r��\���EI���I$r(9��Pa�AUI�s�**�\ ���9Ur�D�W����Tr�\.r$�.QW�]S��L
2B��A�ɑ8Ar��
��r����� (�V�jE�ʣ�s��d��g*8�xˑNR�\����M(�*����(�˕Eˑ�FB�2�QW#$$�dr��
u��AAL*,����vU��"(�QDL��"��+�\\(;gٙ�������dN���L\�p��NL�87}�/6n0xN�Ĭ��<�����z�[�l��֩3����:Z#�����in�7{��o���p�ַĕ�V߅�8��o��w��g=� ٓj�[�Dޛ����ZL�	G��3O�NF�?��\9����N��6�)z�st��Lu`7'R��Q�Uog�3��u��v��/n&��:��V����@����Yx�[~���5����b�^^�^Ys��g��6eE0f�-'L��*�і|;u㎵�{���:�w�,��r�Ŗn#�a3!�p<�ZwQ�;�*ԣ(�Q�Hg�SM�p�l�W��u�nfJ����r�����7=5_O�{]��q�~8ZZsMM��j ����,�4�%A�B�Ma���)����S�}lY��k-j&���Q���$��s��k)�5:44y&F݊��E+�z�:���Q/󛤗�u��:7tΫ�'$�i
j=u���J�?*��2�N�^�+�Nz/�p���n�Rߖr˧î���Ms��^�Ni���s�6���%�؝)�9� h8ݛl'ss��pW۠Y��`�y|����z֍"o�V���uٖJ����1�5�%h�����l���vܯ}�(1w�*�i�.b�(I�����y�M�Y�H�5Fs(�˧�i��^9�k�s��
d\�af�d\��*�5E��/uߗU���/�=�h��|�.V2�z�_��9�ź�{��������5|n��>�ה)q^N����Ԍ�;)ƨ�5g�1����l�J\�$��xr߻��1[>��|�h�^�>P�J�x� fOz�ޜbSu��Rx����D��V����2��m�c;�O�F�@'���nz���ԥ.��E�-�K"ثͯ%�%���<�$��@X�-E��h\�[�G�#m{a�6��T�TǬ�O��V�*�����h�� �@�J�x";�&��{�j���_�H]�zq�bS��s-Af��{�L����ma�;T�͜�F��0$F4S�hf��h��4��|�h�o���q^ů���^��r���bt�>�9L�)���a�{������<3�YZ	�t�B����nbb�V\����n}��IyS���o�u`������ɖ��a�=�M��^�4�=���M��|�Y�yiȻ{f��L��{73�c���é.�1�}�n�87&i'��gjƺ��dJ��8+�a�ۣ�����oz.2̡��X*wy�o�kqc�/o�����^���\�=�ɢY����N�{((�<�vo_�q/LK��~�\�j���A�A���ɐ��tn;`�����T�յM�@�6���U�9�LbU�r��}���OХ� p��oݜ/NW��}�!S��6+9��D�_~~����xˇY�+i�c
�������O�L��J��7�����w�w�*e�&/M�����]ۑ�}�Ԟ���	��~��f��(��1r�Q6s��t�㍷�%�E�Ւ,��ҙm01j���*��ku^^ܔ_�˾���/%�W��U��+N8��ٕ-{Z�{�J-1��^�p�\/;=i4-Yew'��A��6�Ļ�]ST>�ؽE��^Hm{����fT3����jH�w�����[A3�^<
�Լ��3�6x�������[�E���r>9�]l���'=(��x�wɮ���~[�\�ul-���� *o@~�{�asҽʃ�[�F�s��e�κ�9���9���:�3Թw��:��܂q���#�|4Y���B��|�~������aKGqKt�a��fXRU�e2���h5B�е,��kZ[����jb��c�ݏ�7,�C�"����y�\��bWye��:���_�Yg4W���e����lj�;t�J8�f���*��LQ"��}��|�������Ey���iu�r펳�hN���З�c��-�/L��x?C��5����K���k�[=YU�j�v��^���)a�e�l�V^�V*_�CI�����Vo�=M��<h�(�5����^v|Z��b�e	�癯�Y�R��yqkԔ����.���5��|�)��;�yY��(5�i�y^:ٳ��s@��pdf�i��S�8���n���`���SgN�Yq&������*��Ni&1!S΄�dN���v3��NّwJr\�Y��>��Ó�3�C-s�!2�f1m��[C1�P�5��>I��;Dx�4]y�ǺY˫�1�1N��7�*}��
&t��v3���5�Kb'��0��8�Pb>��Q�gO^���V�/�j-����u����<L�:�M�|V�
Oc�O��J�JN�lŬq�{5n虨#p6�IR��eW��(F5R�w��i�.#7\<��[X��33{��^�&3�Ӑ��Yb=j�O�އ5z�g�e26�1:�]�DyR�~��ĺVΊ/��z���ӕ���){J�r��zfr��z��)8����F��u�������]1���vK5]�j����!�hK��#�Q<��9�V���u�.���&�Vׅ¨.:|�h�K��u]�'��<j�dA��+w4��2�*�W���f[��R&Ҟ�*����]x;﷩�7��MÆ��V�u���dRXgگs�Գm��y�gd؍g_�����d�ܢ��KQmX歎�t֊8��T�6+��+:57Z�9o�"�߲7�ck���CM:վ�Y�Z�n�n�1���}�o�����(��AOR����\�a��V�v�w����[�s�F��j��������l���6�W����v.KcN�1VvU�	�n[cJA�6���$]�#*3k��@��Y^��r]泽H�Bs��rj��YVn�oJ���c�.I�2N�-�<�j�^����nƦ��ؒ�L*5	8Ff;�.��WZׇ�b�)��#��B�'�+�/�7���</z��������wZ���[{�ͥ�r�a,�{~���P��BW1zD�&�x����p+.���P�^�8+����X�Y�>D�!�@�FZ�a�h������3�=�7�F�&�w/��s\�2}��gۘg�1*d/i��4�̃��"��L�~b�zf�u�}�~��Ԋ��h��sP׉Ա;"|u!,6�%LNN9��=��Ĝ^��ez����i_��!�K���0_={;���JHZ� ����9��K�DmI�Lu���8�)v�1��X���So�?:�9y���e\��(��F�mn3�f@�sN���K([��%�]����\.�,�k5h�,�e�^8Ni��eu;ť:ikE�Y(��Bmk��#e��꧳�G�u��:��}P�;<�r��Ny��(V��ls�Ԧs���i״E�љ*���K�b���.�հhz��l���݌�֧\3V�2�1�s}�b�N�-[޹4�5���#� ��I�x%�WPܬ�EV��aM���3+���ˀN��ڶw�
񴦿C���2��m
��[]��s�*l9�^:twu3�;�\�Ϥ<�[��!���k��������5.8�	_^Y2Y�؟{�l����O�4��k/8w���o3Kb��+�k�w�]���p�QjZ��-�0+>�I�+�*GV*��{73F���o���+�6�-t�i�=����fZ��^�L�%By�=�I�����a����]��M�1w�Y�X�e�Q"��3ZV�s���M�k4�Xۣd�)�F��f;��Tf&���Ǿ^��r
���\0���[�c�'o�ma nL#�M�ӘX��e�p��^}�MXbe�,��B�-lmѽ�Q��ͤvi���f�k;�d�ݦ%Se�T���gM6E;akzf�FZD�h���@�v��MZs�ī�^>׽�|�t�fz��s���;6]�)]=f��R���\����=�|��t��v�i�ꕶT��[�h>�b����@E�7�+'Տn-���s[�w%Ud�d�J�qU�;/6- �ml���ZT��s=�J]��R�we���qϞS�V�"[����xcW�v�0����_.9r�`�v?��S�X��8t�T3�<]d�?���<Ovq��TG3Y�i�Wkf�����C�2�L��أ+E�:u��R ;��1�=������o7�SϷ�ح)'�j]N�0�S%@Ţ��*���)0��y`�e{=|۱"�)��U����b�j^��u;�~�A�?h�2��%�^��+;���4��]�7��>�)SA3i�{�jF�4<�v�7u6X[S�e�R�|��\[�\t�Gصu/k�YTgV�o���/}��\��95-]$�MfyD����zc�9Go�B���8��b��ؚT��SV�Z�չ�����[��(�z	��_q�%px�;&hY��OZ^E�=��Kd��$vɩ^#r|�J�kER�Y�N�QO�'��"����w�\ñw�Vv)�R�,�ްr��:Y�e��ߕ-�3Fi���2M�.�Tz�ڔZ{۬՛4Ϫ�Ь�[Ӻ,�zc$��E���TQ^0�1ЌR��ʬY����)f ��f�P���(ƳY�i�2J%k�J�c^�<�8���n���v)^�,ܵ�M�N+���be3�'n�.%�-��J��ol���&>��e8��;�n��T��O�<�~ҚO7e��,����+:�I�2���Wټtt���[J��6H�w�l�bS3Ax�ʦT��ϴ��z�r��>������N��Iq�s�^}���������К��+��#�vt�����0W6}3�I8����}]پ7�L��^�*sf����萔��z��n�ѵ�ـ�h�Q���E��K�*v�cH4xk�e�Y���fl��U5m�[�N�lU��Q��x��&ZYE�Z�!Ch�G,��Xf��$��՘�W7d�,����V�=����y�)����M!���zy��=��՜}�9��8S�����SV�Y�U�Uy[e3� ���A`ѡ՚�J͌�Ǫ��U���{E/iX�w��ɾ�GHױ�4z�����(���/_d��O��k]�>ܰ�'ϥ�WR�ᗎc�TW��S�v����=S���3��ޖ���u�gLu�q�8�Oo��c-VLe�����Mb--4N�Y�f�j��Ńe�ۜB���V�F�v�Ϭ,,�v����wݮK���xQ�y�͌؄�V2�ãmAg)�x�c�f�2^Yz�a�}�օ���N\n��Vd��3 �p�J.��N��1���+����Eh�}[3�x�h�Jp���m*�Ϋ�۲�]�7Х�����}C���w��}�W�B���$���sVM�٭m3�ܝJ��:9��Ys�ŃNK��D e�)/i��a�SLꢘzp��4�V�|*��t[�A���oP��l��,���3�?^M�/-Cz�H^��U?gX�}Ioy��}B��{��s��O��������+L�Y��������cZΌʘO���N\J�tȌM�j�����ҏy�p�9]wJBW3XU	�}:��)�u�y�j��$s����r�L�O_��-r��%I�T�6�Pl'5�Y[h׊��='���_r&�H�����oc�!x�^K�*xcPcʚQ.�� լ߷%Ei�N��n�4����F����8�_���oI	���
.db}&������4xidr�J�f�u�,ڶ;&_eT��}�-��,4�q�Nt}G_i�y	de�i��L$��ٟ5,�m������B��~��Me���p9ӓ�0�2��۳Z�r�׮�spk�h�k�y��:�xɾ1o(=���BS��v{�dǑ���b�G	V�:���k�V\Lcm���������t�і1jB>�E�J=�h8b�<�z`��+3�GJG��r�ɏ���N)@e���i�/��]۲ӄPu'�P�B^�C���7p�wŽ�|^�0�Sz#w\��u퐫"I�fei������n�g��t��,��b����}L�k�F�c�����������B�顙ۻF��N��f����sNBJ����0�Lo�{�[B��m��t�@�F�ws�0��YX BZ�:�JR���7�\�>���0w��sD��hќ�O��5g+͵��y�X��'7É�A��T,�Y���YN�-o3���}�Eb���h�V��"��8j��&���b�2���� �π�9��n��4�9Օۗ/�I�q1�Qz7�j�Y���3M���L�ݑn�e<�X�n"ݞ���/Z�w�K�����<�[�k*'���ѥ�+����a�����F�.�ɻ��3�V(+��>�Xce��U�a����>:o`��$�L�Q;N�C7U<�(f�NR��i4�n���D�'Ky����v/C�Ŭt.�+k9m�hJ#-D�I�,TIkuft�����<pnB��yha�;�Xйs����v۳�������ﹸw"�:��:��ň��8��%�FT<���q<�*�]]tp���VYؕ�<�	k�S.�t�s���fN�)������j[@	�zA�����$up
��2R�k�A�ܟ*�Ŗ�<�Z$�����W�4UZ��.��!#;��"�)�8��{7zXg%3Ԫ�h˹�8.���L�aə�zĊqs��=q�#�׫枨��&Je�[P$��ގ�O�G
ˢ2֜��t�Z;��!�cy��U�h��*�z�T4#���l�J��$r�	(n��<C�`���L��*�3�J��� S�mYYSlf%9�<n���PI��&��4fr�����a������ �e�#�͕��Zy��n^�:�OL7�h9�<�;ؘD^���t�(�{����y��j��6 Ⱦ/�eз�V�"v���+BZq�����h����,`p��͜|�W7�O���Z�}���9B���=����,qh��;���I��ߵ��S��P]�	�1ަ��Gp"o=w�=k���T��s(�~�
�ͯn��X����S��_�u�q[NVR$�N�{�{4�x�ûn�	T�/�9On�Jƽ<$]�M P���)�Ԥ��"�@��So3m7PQ��턽G(�L�+5lźzv!���|Wdݚ�uc��S�$fV���۠:�^�����r���]�u�"� t��1�A����u��v;�x�8�ňs���Z%`aiO2��F�����N���J4���P*2��y�ۂZ�00ܟ��w��@��U�TU˝���2��*!:W(*��+iQ4�(�5+$*���Ը���*���RԎUQ��I.b�\�������UQÙ�8�UDQp�Qt�#�UQG*쨣���U��r�s��*a"vE�#��&A��Tr��"PiPjAE�(���щQU
҈�����QDJ�]�g�(����9�r9�0�"Ι,�L"���9QZ!Q*��U$���
��IĨ��p�:UUL�J**���.EUÄUf"�Ar�h\���A�8Us�R�"(�(��CD�E�*��R(���Tr�\��.W(�����E��ED�r�EAE�*s������W"�*�" 9Tr$�K!"�ӤAUFeUQUUQDEŗ+�«�9M����6E�G8Ge�U*�P�ȎQE�r" �.Tr �"�#� ��(9ÕRt*��9ʅJ�G(���>��:j�yqrVe�-���-�K3.�ʉ���b�}�5���5�@��f�\T�t�<wH�W��b�!�?	��K9����f���]��v_~ba�U���y^�p�{=�?2�i�g���:�!�� �y*�<_e������V�V��~�2?��ؾ}�=�o+ϝAZN�	��iHƾ���d��?u��y�{�O��\����МS�Y��)�/+v3֚ԌMs����i�u��!~��>�GOo'<3GyE|�LJ��г~�j}e��r�RyjEn[ښv�O+i����|�����Q��F��v%{��<�:���>ޕ����ԩO�Q"�#�sMN���RYrQ��U��̱�Ɋ$W��z3Z%iƲ�(��p���Z�NYܕyE��V�,��|bt���u�W��W'�����D�Yy�zN�!�ulS5���fY�`����˼eM�:�
��2˞��-���ӎ�1��Q,���r����]2����;���/R�J�mN�l�`�k��,�-]�b��T�gk�n��vd�	�"��4O<pZ^<��)I��^�����E^�����z�M�k���1㲞���)g�Ϣ}�S����{���̓sk#�Z�"���i�3���P�/�s�F/����|=�a-�U��TO ئ�j�h�l�9۩W�_;�ݞ�x�CuuJ�;d���Of��ɰ�X��46�F}a��/Pq]3���sQ�8����ʧ���I5f�!H��S}�y��VЕџ���J��lnД��eU's�1�u:��b�)P��C=6��^B۟	9,�vfh�k�Fb>��3��$����ئZ�m)������#@lK([��)��j�1�8�I�M]��^OJ�_���U��սc�oxk��:����vU	�2K]�+�1��{��O|r�m����X����Zv�b�V"��d=��2)��D����'@�<���w]����ąQ�2���Ԡ�CuE�5M�_�S�74M�J�i��x��O�lª����B����;��ܭ��H{˃�r�$�ZI+b�U��+��Ctݹ4�.�e/Z���5Cb��]��;3hW��	c	�~�9a�i����$�|f+�9\��D$��s�������9�օ���#J*hV������:B�A܃� :�/+�܉�b{�t�n�˦��.��.�Yr�$:Mf��o0��G	�'y�w������;i�(Ќ��6��ԪijYl�i1&�U�l`a�Ee+dU���&9l�J�4��F�5ٹ���Ua�>|*�j1x�p���s*���7ۛ|&��D�+
9m:��fW��j���;����ɯFkϟ�f�}����_�����g,1p�-ʖk0�S�� ��ҌU��N.��woq����������s�]��A���R�Ma����r���V�9�Tֵ��j(��\�O3�.v��26���L���*ε*x56�df�i�/M���bB5������2��PW��x�c&�E��K�R��P����ܥ���=k��A4����$æ��,��S�����%�,;�U�3�=N�����q�j����P���H�~͈e|������v�-ڝ��?��s�1>��x!�9�ʽF��m{�ZR�.Vzft�L�T�{�E����b���x'�*���1m�.y_Y��f^|r|�Kh��x�2ߧ��׷�~~�mG+C�- ��V��z�'0*·�2�[�pm�JxjJ�t���p�Y�ܸ�'Pbsr�d�$b�T��u��2ۺ����{�'O37��V�LT��=��b�[}�M�G,��WK�.}g�E�x���G�T[4��}��]O�O5��w�[�v��츭v����X�h�~	��!�m�c��}�u��G�<�E�����N��m׺�g�sr�t�;�ְ�*O{�����R�o�ym���^�l�3�;�j��7��c��r1i�Q�'vn���h���Y���g�ώ�v��>Uy>�GlkA��NZ}����Z��/��q}8�����ň�o����нۀΡ6��ge�3UV��a��~�E�5�4Ҭ��O@�+���ڟ>��O_G��Wf�L�@�Yc)��h�4�.Zr����=Μz�P}����Tk��=�^M��Z>eD�F�i��L5c��U5jl�2XZ�'t�&S��Z�i�2an���c�4�"J��25�c�mD��N��p��x���=�*����HMoR�agH�;�"n�o<���I%*hS4ء����=��;���0K(�qQ����+:�괜"���>��.so�	�q,뾛w �K�x4P���ܢ:f���&�p�(^�]�f]�UU_-��/>v�7�Qsj��ݱ[vw#Hf��d��J�V��&�{�=%;��}��b��yج�F<�b���Cbu'$�1�͡�Q�n�� }���yP��9�6��#Y̭�������߲�!�K����/�_�zv|Z.B׻r[�I|���)T�rXI٫�>��͸�4���qׯ7a�ץ�����^|�U��uk{@���[�|�ri;ʼ�x���ua���hf�Jpæ�I�ҋ�*���'>��6�,F��%��5�E
^��X�Jƶ;%��U��_6��J��,vq�&���'jT��ּ��\=\�Μ^�髨���,���ڝ�Y�]�1ۘo<t%���1�z$=;��	��gj���C~_V����xq�؄�Pr�[�4�s�ȧ��ڞ\���M䯸��O=Ϊ�=����[*��)h�;��qO:r@O�@����d��(̫���Q|�X�ߎ�fV!�Z���J�\��}@̭���6�)P�����!�:�g��v��<��Tw���T�O�A�'�cDN�#B�s��Dif�Q���� >*l��a"⹟U2���XFe*��e�X�*)�f���+
ܴ�.�i:��(��^l�):�U��[��O�N��9:��۵\:��tf��Y��v��ޫo��}�5�=YZ�=���.ڹ�w�ϟ��:��w���mQ��[mV������Qj�@���A-yj:���M㒤�w��+԰^��~�e��2z����w�Ϭ13a��@�mW���U���F%:�j6�T����Gnמ�ٳ��x5Qde�6���qӭ��r}w��ɤ���=�^�doݳf������+�9��3U�>e+΋�ͳ�33��^v�Q1���&{�P�����ml�Υ��J�}[x$ܰɩ�N���5"v��j�#�j�O�Ƿ$��Tͥ0��cM��ck"d����ke���=�̌>����G���ϩw��[�C��xc�y_�#P��a���p<p��l"ys����ۊ��rdh�e>l�z�á�r�g��+����փrR�(eݸFl(�\w�}�[���dz�=��v��/��ߡFf��y��<y������E�\�N��8��gQ�,Q�����
9d\�"*p���36'��F�����E�T�a����O�Y���k+�a��J��L�Yi��K���i��� 윿VfZ}�/��]��n��q^���n��aj����"gq��ԫ,J���ŗ�~�=�]��B^�wU�o¹-*^k2c�'oZa��o,֕�F�GMP���p�}�U��p�y%N:��Wh��#`ݶ���7����s���:�բ�)XDej����4��LS�31;��o�,0z��y�"v�<_ۓ�ΔqIP�*�T娌�[Yd�r�������u���2�ϨnM�e���u�m���EKL餑5T�Q'[d�a�O���9C���g{����t��G��o�a�;{�� J�̹PL�
�m���|E>�z~�=	��$���H�"���Q�	�T�[c���6R�f���Xl9M�"���J٣��yTu��j-$E�.�6HVM�@�X�+�\�����9�(��cm�+��)�`$�8�xZ�'�1�b�Wf�c���y�{�̢5�ǰ]��X�8eGk�IS�BN���7�����S��͋�ReE�c�pH� un��ػ��UJGts\�I7f��vm�Rc$�i��%���UO�A�"Ƞt�L4,�5�u�N�������sΧG��!2�cڕ1�}������JZr.�Q1��SY�h�W^�sҬE�Q���eΧ�2L�K���i;xsQ��Otф����=����c{>��)�n�J7�3�Gi]�i�����>Kj�T�i�~�<����~�җ��[K�X$�ֈ��ZŤ�hvUs��L�쫁�)Z�*.+]���<;���!.�..�y���$��R��6o�OR�O��^Am{��+�K����"q)X�7w��=�Y��/Q�{K{�R�<�����|�W��>W�kF�Js�&f 1�K�)V��T��ѷ��-B���i���WV�9j�0nT�zc�ra�����}�q�ɉ�e)F�{���A������U+Q:<Ȥ�!١H��`�u���,vn�ugm�%��7�{O��	���"�c-7�r�R]ph	�{M��7�b]�[Y��-���s
/'�SXyX�N��M��M8�T��R�.��ۖ�Nu:+�q�]�$8ٻ.�e� $d�K���}�G��[�{"_�g�vN;L���X�E0�։Ze�@�X�l��S&8lKl�E�����vy��WE�^K%�$�}�r�����4
�Kk�7[I�\fM��U�7f�i6�M2���X�	JTϴ�Ն&lk 14�x��W3�櫉}�-������9�l(�gU�i���4)#P0���fJ)���%�����܆�TVW�g8v��ݱ[vtZ>��;��u�y5��^���
s�y.�T�4adf�b�h�.��U�3����Ǻ�-�^e��u�e���原���/\[jֶS*F19L��]:�i�m^9�	�x�z�:�v�9�b/2�S-sL���U�:��{rQ}n]�¼��\�'���'8���+���zN�[�.禸}ġnSY��y�ѶT�J�*Y$�윻M�E���6t֋�2Qq5����D�=Z�Ɠ�t����vlF��5�ܗ�.r�ֶB�D��ia���14��E�L_}�keEY�~�h*	������Nܺԭo��)�j ����8�tcĭq#,��D�S����}}Ď�n	m)��*�7_���,�D�7�r�u7�0_C٤N}����ฺ?tVw��;E���~��c_P�S�>�|�W��JӾC���p���W=�1�E@���j/g�Kfl��lMu��L���"�N�|uQt\�����i�Rk�TA�{��kؕ��rʣ����]S����br�'�=��M��]�2*�I'�u��|��N{�����Q���WՆ�����ܕ�=�|	�4d���vɩ��L�URE�*[,bv�u����:FE6ְ�sM8ae���'2�zIɠt�a��U+u�Y$�nt���ڛ��+��U�m�5^|E-�F�h8�'I�;�*̳�ݣ��+��)��Qŝ�맋�^���>��>�+�� ��h�4�J���n�t��r��bR�1r�sR����ZƉ7�����k�ކ�k��k|����T6d�T��OI=o�pR�����ϸ�c"��Xm9QN ��LͩT����t̐����;\��uCU7s;��j���"_-�7�X>�Ζ�mvWiZ��1������2�mdnSY�qV�,��ڵ\^f��TR���u�pW(�h��s�WT|eX�kE��a��� K��G�*=��Z�z`v'�9��N����Ҽkn�L�DRZ��L�-u��j׹�10/ڸ��9�zn��Yʗ��KLk>| �֊�T5��#��&��6Z���j1�w"%h�������ܧk~U�Wn����H��77D��t��Z2�e��b3��b
վ���U��^��Y;h��ժw��;x1����-y�(Pc$k��Z)�Yw�w	w�Jm9��l�����x"��M����L\ʙL[u��F���ŅMSƋ2�\"�[1t66���4�0�]���y�����`�+v��yU�*��wy��/+�0�yF���`�f,t�_QX39��sR�	i0Ҳ��E��D>�l�ռ�����4�N�q�w,����Q��6����lDu����]��S[����ѱ��ƾ�d[�5}�r��kOaf��& +x��wD��۹�EV79>��ٕ��n��8@�g,����;)�n��~�Xmӂ�q����Luv�Z�0AɩN�*�.F`5��9A�]�6,�#v�C۶�;�mxo�f�#���ku���.��E�K���bP��p�N-�XXˎcW���f;r�ᖇR�����]'Վ��f���Gn0^[7������!	�'�}Ӳ&�U�㢮N:�nWBR�������E�R9�2�����v���c�u�����A
�ܓz\B#_p6�up�L�D�dNz��0:H^B����y�O�m�$����r��� 5$�).�TN�38�hp�7k���|�@���g�{�O�IY}�f��$KO���2.olz�0d���2(��5�f��*�w�ty�ڴ��4N�ͪ��k�д[�����c�'�iud!`דv��ʎ���q|��=��C�+�����]Þ��z�Eyxn�uۚt.ۮ\PێMݳ��څ������ܒ��5�}w������ܞ�fѐ�Dh�L%\��U`̽n�r��e�W,���]�hj�y���V�U�� }�y��f�u�z�.SAy���D�[����N�;�%��l�!�݈E�8u;�^��vZ�[&Mfnβ�_6�t��Z{��*����Cr���M!�E�3_��/�p�����C^�p�yy�^w͡���;�iz����M @�����v-y����ÀL��)\E�\3!�k[�z;dH�2���y.�9Q�r� �Η��mASk��O^���]Z�`�!�0qS0�N@6�}�a�*�#�[,��I��ԯ�����:x���@�(��\(��OY+kעx�i������ö�U���WN�`�y�N�� �*VB��`�F����3ڏSa�vӏ��n������h QE
| �Ar���.PTPD.Qx��QL��*+$
��DU��T\(#�ZQ��d�(��"�\"+��C"�h!AEQU&\�*	S�\";)P���n2��.W(��R[XTd�R���G*�"��G*���B�����Ur��.TD� ���r����ȮW(��*""���
�� ���Z�W"�.PATr�<�.\�r)�.Ȯ��G9UAG �s�UrV��U�(�\�(� �3��q%	ЭB�UT
��ds�:.QUȹ��DG)�����̊%#��@�p��"���#Q�Q^6p"(�%*
�J��TQTEQTTQR�+�Z��)�fft9q.�B�YTU��W#�+! �P*�������xȪ�(�+R4
��r<eG<NlLȈ�>�t~��9���ә��D��.����udΰk�A��`��]�6���]
Ή ���u:K�e��V��Hf^m�}��Lj�z�2�4R��[約���)[�7OG�^�/��`��9��f�>Mv���n�]��gU��uA�b-��1�K|�����j�;y��Sw`����&s~�~SLc��i�eL�ϔ�����>`-��%V2�Z�4f�Y�L*�̍�.Ҽ��;��n�T���޷�ܜV��������[y�7���m�3mJ̳U�͕�}���e+��0�*Iݫ��54u��/��2i]ܲ.�h>�Aq�8��)u/VO[W^C�pe7IJ��D�ۀ�a-��V�3�j�.6��YP��r�.�ټ$7��g�S�yٯ�R�LE�_�6wzfx�U�(�?!9��J��c�;��bM�׫V�~j�Ct���:��b(��J�18h�ʳ��Qo�@z�cS}���OQ����~��Y�T�h�>k5n)94�2B*a�ލ�
E��A�@M����3�D�,ђ�-��]]���Ș��Yöu�G�	�u���I�ޔ(n����ԍ�Q��2����'��-L��:�5�� ݢy���c��k��n��yc�:p}�%NU�;s$���f��g�1�Nٱ����/egV���	�N��&5�TSh%�V���~�Ky�yկX� �.�'^E�9n�^,��K>�;Ma���S@�`KCN�v.���5��j%}�b����z\��g=�:�}�~B��
��Vs�J�(���@a�mii�QI��
N-�!^9�I�K5	���Pdf�������hN�r�I7t��lVnb�1�k�_������@�/*����-��mn���n���K~��5���l����S���Jd��M���d�!��ۧU��k}���a WWB�7��J�7�e.^��}1�^���K-���Y����ոZ������*anW����3V�5�qTD�!�Y���PgwQ�EyI���)�S�����6x�������R�@�)�
�Fo,����S�{�(���S��ؽE��o��=.��`\y��Ѻ���&Z�P';5�ڡ����h���3����:�"��Z���B�Q؟�]k�cu�������`���!�ypb�mH05ɯ��Va��+�}�F"yܫ�}��y!�S�ܦǱ_�D��Gs���P�&wn�1�(l�x���t�b3Q ��vAÐ~�{�5�q��(������kƽ�,vKO�uZj�'6�-��y��}��b�^�c��ގ�~��V"Bj�{�.��Lyo��f�>x��6��a��[�:��#����xn��j��Mǜ�������ꝲg3S�:}=�!nP�=Wv��%.U��;[4.r�7��c	}���t��G��1U��2l���~	�����t~�zoa����N��:��4)�5��in�>m+��\��gu$ɹ)�I��[��,��P�9+*�}cr�&#��`�4v��4�K/I9�kwҭ"�+_w+̱�������'w%�W�ޞ܏|������I���S�UMga�0�[�J����T�6n�г~^���8|�>�*s5�}gӝ��3��d�%L���s���AH�i��kI��]mB���Ϭ6�p�sE_y#|q��)R�~2���J�ps�k��m��� I�E�ӽ�MKW`���fY"��&�gM�'�L#�#��%�J'�;T��%�V���X-S�R�9E�bt��wzZ󏻠�t�$��;6��&.�3�U�c�Kous�C?}�8c�й籩e�����+`f�4�c�^QK.�F�ֳk	�
c�,��XK�1!U�S�3�2�f�K1�RT�r�I�j�&(Y$��99<�gF���ئ_�w���b�m��jYB܍�6Ϛa�<0G5m�I��k7���Î#�X6��W�0��HTuo�ȃ��ʝ]��*u���� ����j���[K�ƾ��lޭ�O/Q~땽��,��=y�*Y�y3���_�������m���+h.;G�>�����ؚ�nZA�U�� <��x��9���O�����k�[gؕÜ���kΑm+NsBZ��N�/q+��:�N�Vғگys??!6�+�=�\X��~�.jU)���օ5���Z8���T�qzSlZ���Vѳ�D���l�ȩ3��M���(ݵQe6�Z�ՆN�t���$��ӌϴt%4MU�c��M^� ��w/J���ɲ�Rw��D�Y{�%	�[����S��ݛƝ���wl�H�[���d�s;��1�g)F��]��Z�wvW?��nfV�,�������l;���u�lǖ�6\�Aj���z1-g��d����v�R��)�A-��W���,�0�[r�h�!���{ox�Ԕ����R!���8�����fS�PiM��r���خw4�\�-q*P�*��͆������C�w��Ν�ѳ�[���co2jC5�&FP����Bd|M�`+��#gּ����7��ڜ߻z�AL桘�21��Qm���x�(i�џ����>6n���5M��'�:e�;qhݱ�Kn�5㐙Q��1*�t�̩̌Nŝ� �Z�(�:m␚ݢ��`��:��L�P_�z���s����گ,�#���ݦP��������ߊ\W����U.�T����_S���h+�>�2��98�������"b�v����̬Z��k�6��N：;�+w4�m�Ek,%�|�.�R��]���\V�Q�4���ḻ�^i�l�d��IP��j+�f7 \0S�PF���zv�Mw5%��՜�����{k����k<DnbmSD��C�z���˱����C� y���t�㕳�Z���}���-ҬR ���3�e����a]Na�C�T1]u��%%_}T7C�mZ�޵��W�KZ[T��*̲�Q,�����8	P�qK<9�~�@���@�I'nr�ڽk2��ai�VF��«o119�}ƶ6(�:r򥹻�w6H}#�}Qw�O���u�[�c�]^�G--��M�w`���8�{�����Wa�*)�b2�CL�:���l*��j;8m��p�0����2�}Ca��R�˘�4Sh%��V�j�i�E�0�LaA�,�oړޒ�g��Os��?���*-��%���$�ߔO�}Y�	��ŅF��Dϙc�m3,{�RLW�$�Xbf�a��o��T�x�N@e;�F�"���ʳ�9�Lb��Y�j�a��O�����e�j�N��*�(K�hշN��ʏf�fdO����T���vӬ�h��U��5�b
m3��ɧ.'�Ve3���蜂]2�����c+`[�֧�	�j\�\�\ Kq_�@��+ ��}��?d���w���~��b� [����2_!����>���+�8�p�^wb�݌iyd]J3�n$=~���>��eԻ&�Gt�G�� ���(oQ�����������5n�z�g��ށSiɷ���O�͚�-xO7�I��RI^��Y�nڝ��]�����!����v��(�V���&P�F���nk�
�4�̌�`�nz3C|�<���\�8xuݮNa�#zKͦS5'a��L�,�Z�g4�?su��)�gd��j�l� �
�[�98p�$��c*��Ro�\�~���p��`�;��v��/�N�L����M��*��0� ����R�^�}[3����~��X�Ab�};ܵU�PDw���F^�R�*	��%K#�Y����C4�JKL��M�nّ�~������\�|i�����(������o�r���+FD�Y�'�\ד��eOa��ȧ���<y���H����`ӈ�3�V�	��
>ŬU6N2��p���%C��i�j�c���ހ�`ї���\��r���ł�ᓬ�v���d�I�J�h��'�\��9�<��wR��]��u���	�,�P6�9��B��yE�Π����D�:�N���r<��D�	�ΪH����~�t��~��^��({�唡5C�o1毻�:1��F�)v��j��p�ê��-������ݓ�/U���y���V�c��}���FE�rk��mj�;��"�)N߱nO�% m(/0�;�b�ec����Ji��R1U{d����O3�W/n��f�����+��S|}�=}�#D�<�{�����|��H�{#}�����.�gF���y�׾~��(i�!�,�ڬ[���u�r����b�.���V/Uޓ��{
��,�Lb�e��5��T%t~�M���d"�ǫM�Zv.-3�CZ��N4�E06�|D��2a�z;Λ�^i^�h*H7��s�?��y�ۈk���{�Jg���Ͳ�}��[jbdK�n��{e��,��'pT��M]�j��͋E�	KE�j�Op�A�Ҳh3��딴��Pu�5k���}��R԰�\\���8Xy�d��կMl�����Z�5'b�)=O����c2y	l�G�W���n���=V�F-��h�@G.�Ҙ�c:i(<L�gL�v��+en����`kt�3B_����@ٷ�V��T�3G��ߕNk�ʭ��� ��t}��yr��)���nۦ���ӣ��Vms�OP����o��o���
^����j�UI�/����0��[gؕ��\mz�GP�/���-�N^�BmrڋCIӊ�^K%g+جl�J��bW�pv�X67�+����<��U>�j��h-T̀�gĪ�"�Z�����*��c��/1�0r�va^e�t'�S)���Un��V&[s^���3g�ʴ��h���땼z>�06�u�������['�"�\�t���;Z���W{� ^����^{�dm�N��,�e�晁-��U����6����ma��ܭ'�,}.{N�}V�f�&�PF�aXbg�a��zG�[T�v���.�g]�^��H�R��©ˇާ�������j��7//c��*%)�r�J$��i�.���)f0v�6HS(�2���#�NnC+7VP;t����)��z,�^�f��}2�$�����49W���_33s�#��H\�;1��Y�U|�]V8�;p�O��j�l�����j��_y�c}%-������g{����q���]zc���)����U�xl���Z�:�Z�*=�n��{�dP�Q���Z	���:et�H�x۬p�ưy�a���Ŵ�����U^��c.5#9�¬�«j�3Kzͨ�ģ�ʘ>ړ�B�1/>ᇽ{�s�2�U��2=�]������&��]�7}�¼�
\|�3sۆ�{�[�����2�}�j�,ԳR�-W>���-,P]��Ni3�������e�2U<��ݑF�Y��E��&�@���h���I�j�mS�YFz��g�����5�Z��̍�e2����^KI@5$ ��������d^9�B�){X�/���p���9���'-e�)W����`�����A��l��fh-5��Ԯ�z.���qF��y��wq8��L�g�7:q���W��F#O�(U��E��y�wu���9�+�[��D�P���3��'���GW=�B���}8�r���v�)Ңsl�)�ަc��-Bl���12�=]�9��S�|�J� �u
��N��m�t\�lq7�<}�|��TU�5{�g43c����x�;�uBy���	�c����;�����*�/P�4��`/������Zv�=wF�Ls�c�C4M󆯏3���v�7U˵k�������,��H�,�N�^�2��=o�A�f_
=��"��������N�vF��{�0s��f�qZYv��K�����BC�d�Yv\�/D��3]!VͣL����O)I��Kņs:�<�rp�;�/]}�k����As���`��4�^�;׺���n`��s�= k~�תQb=K\�����`'������� d�X�F�8��y��a�c�2R-ñ�:6�9�x�����}�};�����윆�a�|�G%�c��\�!���M�YaB���ܲ`���q�gΘ��(��[���/�;�������K+\��j5��[�G<���i��0���W�����/UXf�q�&��Ea��4�,<{�=f�!������ے��8#W�����w�&s4�q'Lh|�o#x-�}�.E��o���ȅb�B�-%K	Jw$����K�e�X��!�p��hZ-�H׎3=��yЮ��7 ?Xy{T#�.6����sc��[Y�Vws�������_�\�%p{)��5�W[5.���y�h�7����u䱸:)��dy��0�!F<"q����R�HW�1^�XpcJ��i*{�	�\����(Y���t9e1ql�R�sN�:U���oj�U�q�余�<�NH��a�Sta���1������j�XʠO���ե��o���&����q��zEqо�79^`"�n��Ebt����7	G���]�-7N<yc�s��ŏG�M��g���1^�q���L�ܢa�3�8B�}͓-�i��]�C�X.�S���)� ��G�#5ǏE�}` p+�hT1f����/�.��qP��Q�$/o����m��+C59m�欬�u��ч�1����bh���Kk�X�;2�^��e����0�<�,�F�ۋ����r!څ�s��\U͋sf�zy��[Eo�K+�j;�Y��Y�;X���]�`VἭ>F�c�[H^q<ul[u�;�_)�����٥;.�|��x���	 9��8���:���I�)��V]�>�I>������+z��;k��4��i^9��G}��5+�����>�47�HWa�]�d,*Z[m��,�hf�M�n��ͨr��w���S8r��5�ێu�-���E�ƛ-�����L���w�4�o{4"V�4rޞ���!w�k��!uт���n��:��;F�;��^г��B�\�4zֻ�6�r:����2��Jt.���a�	f���W�b���|�Յ�ଚ$��w ���oJ�g. �k:��֌�^�v/?f{�%+P�Nk7�hf�Ps��,�ݰ�kn]'`��z!���Ll������q\���WKY]{j瞌�h�<E�=��7�u<��v�e��?�����"��+hEÜ�*�EG9DU-V�"��$��!��AA��˲�(�#�ETA�(Ԍ���8�����*�N!���"��2��eL�5;��Fl��"���%t
"5�̹̐\�ȻJ��L(�U×�)˜�*��TU�9\�W+�(�J��W ����ʣ�!M��eDE\��E�p���*!!g(�hp�$�T�J
�L��J�
8Q�#�\��0��˳��9W9Ȫ���Z�0�(�$�dr�9�\#�Tp����^B��2���9E�1$���S(�"*
�]:�M0��Rq ���(A\�9ª=���E<eQ\�
.ȋǉ�t�TTW
��)D���\礏�&� (  C�*^��]���Y�9�y��gMr��:_p��F\t;}��]rz� Q]:q��(5p|	�>�5n4�T;��O�>#L��%I.�Tv&(6I�e1eQo����m-G"�*�Ϻj�ka�0Ɍ[^+5�5��-J�A�/ff쫇m��Mv�N�d˶���t����Df0O�vu�鑣V�xds�M�\�Zo��i5����X�K/=?gO�.�Sly���C��X�:���[9"��.���O�<s��(AM�}M���n�K�bnk[*����y�D㻪��us�.��2�ߦ&�>[fHu-]9p,"�B�9	�ü�F��Iͭ�v_�;J�B���;���L�˼��O@S"9�h���k��Uq�"%�ط	1L��_zb�i���"ޞ�������j��#GtE�k3��B�����鏸m��ϭ��Y�\���;����lVEP׋����w�]m�m�s������<�uM���]�pI>�δa�V��G���#Ge2s�K(b���)�NM �z�����7�;X���۟�� w3m$�����s�����{�v�A�ݯ!�^׍/�/�v�5��d��@'yO�?�?p����Q4��b�K��!p��{�{>ɘ�M]�EWђ�슻��J=�lB�WYZ�����r�/3M�eN�vp b���F��wq Z���Wfa	��WH���Ǵ{�n@�~�u���o��$�*nN1}�M�_sN���mCe�f���ѥ0��j�ܭ���������6�^�1�>�L��1��̲�/�5�g(SlB|�.�{�Zy�X�m�
�1-�c�v�5p��i>����l�ʕ��x��7��KK���8V.�u�g~���K���1��6��и"2�8�Sf�%od;�	I�u��M6Y�a6�N�l�F�';,<�F?5�.�)����#�Z/���*
��g70�+�ҨF�s_\��ș����}�.9�o�f��C� PR[%9���~z�ʓ�qx$m����=-�)ʎ�HSp�Ĵ�eG5�~�Ȃ��m3o0zM�tGQ�K#,Օ�'\	u�8-;�U%��U���M��f8<?]�V=���n�o�!�-�i��l#1�.we�E�Pǟ�m�vǃ4zŅ���7�yFIp�˫]�_T��s*C�)~	�0<3ZnC�����uջ�s
ۏO�*Z�ឈ�[���T
d�]Ք]�3w]D�l;�2��7\���!�?*����b2j)�}�GN�!͙Fێ{�/-��	��+���B��Y
�y=s���5�����;�%��}L6��1�a`���@rU)P�r�*
�
����^�e����VK�H�æ7�Ktʢ�YbƹB�e��#cͮ��/`����x#�����s���\���tG`݉v^�W=��ͧ���)�;g�k��[:1�O�S�{k�O��t8�N�w��l�,�b�{زn	Fm�H��6�e�׮s*����ލq���c����d ��xV�4�f�MnZ�&8��ܷ�~I�h�S ���eb�a����X��N�FT��j��Oq�7�nk��Iq���r��ſw)h�`XOJ�)�\q��	�:*�ۣc�Ed&z�m�kH�λۦ�摛᳞]M�r�-:��+]+���}ӓ�B{Ƹ���a�\V'�ט5�蝆��s�OK>����tf���Vی{(�x,���l4T�2c�;t��S$үh��w��1���,B-��>�p���S�nu�L��6.���aOL�1ڮk��m]��n��1|6/�6�1�;����M:r��ׯ���m�t�웃�L	ؽҢ/g37�[��k�m�;��qlw[Q-��Ҕ�Ϩ��!��%�yʒB�%���Y��9�l��3N��X��2Y�WW=�s+l�E7D'~ع�,Е3�T-���/V5�W#|�^�E����{���:aè4�pF&+�*��7N�1׺�����\Cj"���\ҷvo�)�>�טݘ�.W���'e����J�gM�#��ݨS����@��g�)p9��ˇ�wq�Zr����xs�FF���i-��Y�kd���A�݅8�r�݌z�S��zB��5��)�,%O�,B�����f��}R/�ջ-��v����#4/�B���!Hw�ø!B_?;y�b��L��=�]{m�̬�E� ط�аe��ޝ~�3���FOtE���um�Ms�q=!�&sVK��r��E�ꑜ�7M�y8CI3�1|�xOrrjzc�(!�������J�5s�S���d�p9���Y�J#-���U�`eM};p,5�Ϗ,e�<��s��l?-xV��5V�;�|�{���w�d�L4�3�vلS�
k̖U����@��\[[S~��5�o��ğ��̂��ψWt�?[:�)��.��C�ѐ���q�\d�h����ϵWW�zվ\B|w�WQ��d�s����E3v�SM7vP�Dp����SFJ{Lx������Df�q���t���'��
͇��;䵝X�[���κ������Cr���S�Zĉ�<U��U��t��~��k~Y�u�Y���;�l��W�i;�������}��E�7�-��/�;��1`��s���SLk�������;0b�1�9�N!}����;�`�o�='a���_?!�.m	�zd�l���!�U'w�M�P�D�0{�ko�K�H6�s��|�z��F�CS�{�䗏8\!fvn��ݞ9��6��*<������-�"g��f���jc0�c,ԧ�\F!Mq�_�a��2=]�7������[9Usr��i�3��޻��Oh�5�ƙ"�źQ~h��xiަUb
q	����Y@>�
��'������K�n��/L��'����t�ʥ���ȷxf���j8���L1�3g�Mrs#��i�l�$Z��Y���k�^i�� Y���.�\�=��B�V{�*6oxh�@朎�~��D�ds���uL�RA���(_l]J�7Tt��",ȝ�\���&s:#,��X�oY�3s胠ؿ���#��ƺ[3��dh1���)�t]48�]1M��.���^w�/N��R,�g.s�t�����z����vie<��|�"bX�WcM�m�F:�r탛��B��;��N�l�u�1�*Ǟ9���U[��h��޽3�d�j��M;���K�w]�K���Zbi���2C���́`�f�f��F0�m�k&���/�:�u��t�B�x��~"��?[:�w�xwQ<�@��x�y8�J�<���Uf����{�d*��z�{4h��F �r���[jb���Z�Z%L&^�m�%����y�2�)��a��YJ��Y��9Rr�B>z��-�w�t�伽Vc� �����|�Ɵ��)�ش���K��b����C��nu�����w�������q�U2�3#��s@����~�뜱A`��c��s
g��z�oP�͌�ӽ�f+�����y�M����N��Ss�6�ζ}�C`��%�Yu��mՂKV���.�Һ���߫@_4d���Z�5�N
�(w��N��j�w�=s���p)��� �̎�پu��p�'�̱�N<�����e����K*���
����0��z���U&�ꈵ��p�$�U���r[�c��_^�{K�+ٌ���oWL�c����*���U�g(GV�=�r�h7�sH���G�R8-��l�,y*׽�\��w�J&�873n��,�,�zu�n�b��.����f�5�L6iF8}k�(swB����El��r����e*]ֻAܣ������إ�������<��8�\BC�E:lE�e��t[wt��=��vaډ.y���5�٨�7Mn��}���=�BA�h��ٲS��gV�=�r���7kv�|�c��b*��@9Jڶs��+��#�4Kv8t�["5�m�����a��p�}Q�	�����l�P�~_�U�L=W{�{pVeجty%��S�����W�F��U'�xl]f��Ow�3:�5���2q���
���j���+w,t#�G���'��i�h�k������}���k]2�R�ɖlqq&�k��m�Bf���������bK��M��q\z���WWT=yt�S+�~Q^ȇr�!����[ �̿3�.�7-ͯ�}�3a毮�NY���]�`RQ�7uc��k���s*C׹K�OM��xm��x��;��햴�75����($9�6p�L�F!p��r]�we;����]�~���C*�l��N�Y�^�Ӑ��z�pC�gFp�p��H�Y�{nخ���A?K2.���=!H��L���n淸���}�l�k���p_`Kb�q�)�|b@O-�_���WK��f=���s��E��y�f����w��xL��"��_���������3i��6zy�MPA�{8�c$�z���a���~��v�yj�/���ŵ�/HbZ�g:{�]�9� �Cs,�;W+74���%ӈ=����̨zn�y��p4f��{�M	��%����ee��`�a�)�����}��Qތ�|�v�w��
mw[r6Y�"���
n1�4�{�~�z���`���o{";a��9Q���y�)(oj��݊�o{*���$@R8@�m5C�w�PiF�2�{�N��*t�R�����a3�Z���L���b����od��{
��"9��{�R�$^ɏn���=W��nk�oO����g��;�L�z����ε��^d�4h�̤9ea�Ӡ��CZ�
��'�4{��x��@�N�H��������#���qB��t�����9��tѦ��tvM�X||���g�Wy�5����h(���yC��(�Nz�eXO^a������m;��%��Rܞ��
9]ou%��66�w4�
e���D��ĥ.�F7�ȉ��d)�V�Ɇ׮��ưFv��45!��q������Q�8�ʉ���"�R�mP�wd��l��U][7ѹ�y�e���*��#P]��Ҧ�O@X��!a�!��!�v��q�fk�R�&�����BBkvYR���}����y�t���Z8�I�sr��Q�v��p��y�� JE�_��{�m���S;J���1�曻)��ރqz�0�S�%�uq���#OL�~�cBᶦ��X��-�QϺ�=f��1�+�:_��%���������ߍ����j�i�Y��ю#i����e�Z�};[��^��ǖc/	��e�o�M��5�9�z�7�șw&�t��*󕉂&��y�؊~�W�,��'�S6��En%ݰ� ��7&��3!7W5���s9*�E�-gU�� ��1D5e<���X�q�t�zh�ö�����a	m�9I�:��[n%FM�H��K�w�y.��Auhg��6��N�2����S]s/~J��Ze��*v]����.+��r��[�I�6������5C���0kwL��T�/�^]2��Ou}8�af����P`(s^=��IR�w�}؍t�F��_������AۙM5߲3�����n2�u���6���[*��sdOMp^pb}�;��V�4g����˪�E�t�K_mF�QޤF����{}�'Me0,a�/X��=5�gY�zUkC�J�� 9���ſ��t�Qꇧ��i��-ļ��'=�Q���1�!l�1���n�-f�=��P��lç��=]�b����#��NѨ%A���W<撫������ʊS�E�%���z�SX��\Bs�5[r���˺cv^�j��$���i�3�9�oT����\��!��.��6E��JT�L�%�������Æ�v�|"�K*g�$�e�8�E{�����A[`�t��Z��q5�*1�`a��Zv���Aw�Ta��{!9���E���cokH�zҥ�y��H�Yo&�ߞn��^c�ㄓ��T(0�Y��;��l���Vκ�3���!Bl�w��f�~���!4��Y��5.�<?�l��**�����HQ�y�9w��E�T[*�4�M�|V?[%�8�L���TU��#ѣD�o����ވy)�B��z�}|T���� �b��NhZ�l�WC�zz�ܘ�a���`�0.u�W4��I۳�*�7׍p��+!�]lE �+g�X��g��&7G=2�j�n�mG8�pSk�3)6E�;Y��w�'���0~��q��A�~�^V��ҶrE`\7mᕋ����SM��^�jwgU�;��TN��w�j'��[*�s�`O�1���N��G����b�j�v�4��Dq��Oϧ�ct+H~��4�Ӕ+�J�w�5Dc�=C����
i�'�H���|kwiC�X��v�E�vy=�Y�x��F{~�5Tʛ��j��#E{�g��ȡ��:
������wꪧm����� ԏ�E�#�-��cc��z�C�F��S�7���T�[=�����i�.�c";�b�-m�oN����d<���K~�o��	x��@g�Z�����W;�wh��N^M�ܳP�Dg�v����5��+�į����[��7�k�~�A�~˷�Sr�[�1wg��Q�yڤ��1;��]Y�ηuk�b��9��%�\2�d�!>KY�eW�8q45�:�Ş�	ܘ�����g�� �Q�]�8.:���3�=� �^[.�M�pm��;�~�÷���g]_��.M �i�w5$c�(I���v�Wcj�˖�t�G$斖��C]$�q+j��>Y/z��`�̎��#-U@	��G)����P/xa�5k/-�ɽ��V%ٜq��H�q�u���/8�q;d=�]�W������������t�\�8�[��ɄJ�ն�Dr�ꚵ:����;�0[�.�+��;� ��FFf�S��G5z6��볷�M�ʊ2S��7�Ǿ=��y;�gvW\CY!m��-�KIC��U��)�j�Σ�(f��{u����O�1���7i�6�B��;�޽�����Lh�y��k�&y�O���rd��T$���=�VI��m�$�[�*��u�G8�6Ei�j7ޏ��%UX5��v/M�	s=�(�I��n����M�b�T*�N^fi�yhg�o׳}�*4�0�*$�ƹ�Ý�gl�1k�׾3�c�Z2]
Rk�}�5�Ytk�1Pj8�Ӷ� ������D\BL��i0�px�7t���ũ)�5���/���p6����ɞXѦ���p>����R�z��G
7�Pc����q�,�gKg��=��Rw�h�b��r��
��WReݑ4xm�$���A�h��R���]���fc[K��_b��aא�9C3Ǉ���gTwjR�|~JfwF+L�Ņ�+ǕXMfTF�I.����� �P�рl=W\��^��+-�m���gCeX��;4��^n�6NS̔u'q��o�l�ua�hz37i�pV���͝��[��������{C��͜���3.���uMg�HC����3��EΠ�C-hl���&w���E��ڞ,���S���Mڮ�\J�w�Y��JB{F�7��6���2T��qQ�i�y͋c�]X�D��}��A��/��gDp�S�:ٔ�Zf1;@l��U���_?�k��0ۓX!�b�6��ޯ��Lf|��c�.bA��0�:ݺZE�01*_��[ۇ1���'���@� K�b����n�a��r����u�\u{z��NgwD+_�xl%|�M<[ڹ�*��ԟMW���p�lWjKH�
�hv�K�È9�я2[ҽ��јw`��&�f���|��G���F����=��hf,����<l�@���od�fd�X��j0ӣ�ҩ�'N�6��ʘGNg:���z$d<<�r�L��tV7�n9��E��>�}5���\�W��U��f���ͽRкS�˕�L�a�j�G�H��Ȳ)n��0XTt���.̓zv�������}�f=4_����p9�Эw͚25�c��ǚv+c6'*k��=wJ���u�]l:AN���ysuA��26�q��ɼ����|5m����/��$���;�+��h��3��Ţ��Φ��V�곚�O$�E&<���뿿;?|���S���ADDr ���UT�rˁ�E*�#�Zr�U}��E�AqӡE	�Tz�*
qӸ��s��<x�*�EEE�(�EgJ�r��x˸�8���:����L�9JU��<IUA��4��/MՉN��Z��az�ĦSNU¥B���<K��zz�.А��9L��FV�r�A���*�G3
��.J���Dȃ�����W\����1*e8ʠ���Mq�9���*ȋ�g5�N&�(��B�"JUns�u���!ʎE8�&h�E��fTD[O-�,�NT��9N�E.EU\���ԓ��j�Zۄ�wk;T5������%�=+/�7z"��K����0{����2h��4�<�O�Cpn�
:��9bb�dNi����D��\B*-�C�|3�-��pDewK�^Y��Q���d�Έ�:��k{'u�R/�,��w��N���5���Hv��M�h�^Z�'E�tv�S]M�kr]��f�܈�ժ�N����˛J�J���L���! �>����Ng�����)O]��y�:��ɮ��Q<���ެ��.��d]�Bn#Yҹ�{y��lX���dg�;�9��~S�y�ȍ�{����49�-��_mז��P����L����VD8t�l#2e�p�Y\:"�k�]3�&�6n��C�F�5�\�꯮�����U?�o����i�G8ְ����$���3�����,ڞ�-�B�Fp��%��\�⺞��]�tkR
gcw�sh��ue-��=���!�����őϚ�=ɗ�S�&xT1���a4g�d����/Fm�)��S��R��R*GT�!�-�y6�Z�`N(�9)�LH	��SQ]6&BE��
I��{_�3&r��u��k;�N�pR��6٣e�j�02�����b��_��~�ߌ-��֨em��JEdy&ￇ3R6��Y�g��� 5��|6���3;-��J��4c�i����Ä�&r����D9����b�t^+{�ے6�f?^2O�*�������.�v�����:�!w��5;Ԋ����|w��j]�`~g[����(���Th�w��hu\S�p0WD�%���E�&pS`\6����ʞ���k��g6�C��^ѧzn1�:9�빇,�q�\����d'�k��+��棪��t���q+�c���h,�-{��4T���٠��M5��)�,��^ۧ'�n�D͍��`F��'[Gl�θ�`b��a�=����z�%��-�2�w�����vN�UT�g���и��"���P竈�*�8��:Gϳ�-���y��"૽n�O}Wu����o�����-i�)LY
")���]
k�Nz�U��6W^9h{bn<�]i�O�4�m��ϵK��l*c}��QJ!;����x���Z�
o%�wq��Р��Vz�p�&s_y�t����mǖ{�70��`�J+��lC������y��s�
ڻ�F�	��]�,H�׆�]$�Q�5�s�<���� �qoX�t�6CBC[!�5K�մ¾�Nt=�4l�n5�����eL�k�p�[�B���,�eHw�;���=�N?ǃ5b9�]`��\�73]�n@�e�8˵�u8��Y�Wؓ|E>�.XU���	m��w��s�,�jv�k�S��-�\�؃�h,��Mۭ�F�������G�^ɜ6U��At��fd|��U�pcm�SaïW�x�I$�7e��A~�i�%F��c����bY�zK��)5Ȏ���g9��y|������曺�韈�n���l�8CJ3�+s��<'�1 '�zi���3}��M�m��y�p�ـE��?U3����z�<F�EK,���� `X:v9��3�t_5t�`��6�x�EL��]�iL:�M�9N�j ���s������%�z�{@�k���J��WS��Xt��F��׃�c��̎M�yƊn�~�gW"�{��"�C�	�>�<v'�hg��t^�$�$�[c�';����k����Npw��<E�v�4�%wHtCO	���3< ݇���kU�w���Fָ/8)���];�L���3ߗNh���i�y���K�U�-c<��7<0��+�>w��v�A��Os����q�w��f_��e;�IF���V=cT�p�������z���O��uM췄�{� m�e���Jzk��,r���I9u��Y��&�m*��/��V8��Cq��ה�Ƕ]�K�o-���b�(�4K[��K,f���W�����׸����ǈf��9H�x�H>';���^�/��֪{2Z�
�]J}��o��M�5���'Һzp�|��1v��Y�1b MfepX�؈q��Й��4�
�F�aF���}3F�!�����Ϡ˛�Y$=�'l�|�v��3���k���?=)�I�ggK����lS4�wKv����y�ܓPViȞg�+E�~ѭ��ʙ�I"���t_��h�鮮{�70����g`u�{�{��{٥ͷ1����{�S��BNBs5����H2n�.�cZ��2�Wn���[fs�������S�t4w�D�h��ض`����3[:�Do�v�
O��]sA�W���.��L�3��=�v���E1� ��Sd4[@5���9n�����qld�UY��Py�j;ʬ��̣$�V˺˿^]5����g�2��tC�`T�ҶrE`\7wy�ҷ������Zu�9��O����~���w5��N�Y��C��~/�N�-�$:�r��2���gu�ĝ;�v�ޱ|���$��t��(��~"�
g�T;�r��Q7橞s��G2���"kQ���Od���j-���f����>j7v��L��j�h�+��8�n�E	�w���̨s�%�-�M�$����.!�F�>����W󂽊>q�)ܙ�n|�j��gބ6-8�W;�.���F�����w����P��d��b�*��;�ȏ5��T��)R]�nu�8rF�n�P��x�"���(��m�4�ܫ���We���-%G�򴸡+�B�,��*�X�|�ϥ���숽�{��`����b���ƍ���XIz����p��/�1��'x��Q���;Brב8+;�l'|��A�S��~²p�GU�q7�s,�w�gI�m�M��u���X�-�`X�~�ebnrYS_NЦ�������cG
s���:^fw�RS|6{�I���� ���FtE�����-f��o\:J@-'�km�f�j'b���{�G��^oJ��k�����U�~� �L�]�щ�N�:.�g���k�4���֓k�1Se3\Gj�Rxk�:φ{��B�����)�٦�fG*-�C[$�
�s���w�9�z]�nf��1�=B}���_�U�;���2n���������� ֤� c��'U;ZfsL��R����OF˺W3r�	yj0x)�NMt���.T�v���Um�ٙ�i�,_#!�X�u�;��E�C�gY�Y����#��Y=���ǉ����GL�#_�����\+f�w�{P��SMĿ(� �E4�x'�x��s�3j��"�9��1�+�h[�ݾS��-�2u��wV�����eH~P�����ci�R�\�OQ��ps���v�J���ĪzR�Kf��R���%��1~Ocq���w>�k�cn�R�L��
��X�I4h�{R:V�;:Vz"������yfh�Sލ�.uۗ�Engd�2���&\���{m�*��Aٕ�u�A�9$D��8��I����J�g�`�:��<7K%�H-��7N˺�r�~멙�d�t��V�ޒ^�i:M�z��6��̐�5<�:3�ۅbL�2�g�CS��b�c?Li-�=�t�/9�&���R��Q'��2rX���Fߢ��S\�W�[c���O��b@O>�/��8w��}6�-��28�M>�|�w�4�H��#n6[��,2���[z5�Kd�w��[�m�+g��r!n������g��n���m���t�2ʌ�V*�mx�{�-�������R�5{2N�b�ёͳ����6�g��=gJp�u���v<�׻�hr"��SFB{��n���,z�@��D�۞i�=B�|QM����K�QS|6q�Siܰ�Nu�hԲC�K�gt�%��;�7&z�o4�>X�����ʊ�2��g�m��7�=��䩶[h��]q�w��!`�
̧'f��xj�����5�#�W��>�p���<�����~�ʄ �ʵ���]���k;s6�v���b�Q~��x���B�O��eXOq�ݘ�^n�oSeS݋���k�FpY��a[��c�)���*+��i^x�Ճ�+�1�{W;�5���̻��%��3`U�(g�z��EǍ���Xg[Y};��C�3F� ��'V�o_�O���|�x�鱮9n��{�:#K��AE� }%��=��;��7Lm�c�xDj�|,�K��t*m��t�TS2�N�D53�4�.��`�R���.�R�9/[c����UjYw��)c�>���,������aC�R�%�~�t���^-2��Q��أ{����~��ג�En�-S�H�.�AB۵�k�T:莐�`�t�U5�.ؼ�0��H�f��록1s�S�]��8/ᵻ,�#]��hSwC�T��A��Uo{櫐�׍�{!��ةm*7�=��82����N�R��P��2{�*������L%v0�;x�=.��s-���I��M���tݶ�8C4�9"�v��8Og"`'�OX:�e�v����G+x��ll�dSp.�,��L�'����O�a��]�[};}�`�ZC�.k��v���^�v<?\�[�3#�����)�����%�<�*�g��~��y��3TK�L�#z�n�#���@��nBX�O=f���ޙ��-��g^+�ȡ>������6��R�.:�n���1]}jq�z�'#!�5�'z3�ܐ����MۙM5ݔ0��.[�=ͳ�ܴ�2u��E� ����Mk˒l8�XhVvh�R�M� ��f=R�a��}2;
t��#���4�̩�}���M�7W�{:&�y�����G]峞[����o�n�6���D�+p�Ɏ�o��u+n.�$��S���^^���ޕyA��O�5�u(m�Gzw���m筟�ν،��O8)�C�EF�w�:��Z�����OR!��c�u v˝$�S.dv��_[��n�	�OX��=z�3� �kva�)�i;�!�+=�y��ԧi�e�m�!�[�@��;�f�n�>�R��#�\G9Q����UqlL͡��sH�xu�J��R�Cd'�˪�>7[�sX���_�S�]�z�T�6��]��z��dVhq#�����z�j������r���'sQf�t�ʯ(��"�9=L6P��W\⁸;o��yd��w�=L���b���ʽ�I�����1���ֈ7P�:�;��Xm4�L]�)�;���huGK����f�)�}PP�'s9螒C-}�#�`>7��c_u{�!�Ƣ��!���vg�o��`����֩`�зIo���g�]b�ϛ�5�M�U��+�dr����;&��P��9W����!,i�zy�`�eL����-�Fe�'���@���ۉ���H��=5��c%86��Z���lY\�S=z�1]��)��4���[����]z+t��|�KmW�(�^;�ty��yj�~���j�vgM�~�ͺB3>̂����.��[�ӯo��w��cV2���b��vc=֢\A1>����]���4��w�־��M(��i�>��G����a��S���YoM�<���ĶqyOL�%
fQ���~Q8��ݔ�=�qR�C�9�N�e�#��Ea3�n�kNENv�r8=�E���p)͡`�/��z�
+�߈��3�����Y�T�=V���)�V;n�0>�:�nWC͎��|��~�5������I��U�j�C_�4�2��%�H�S?`�7tN�dg���w>P���G�"}��ቮ�����32�pә��6�iMFjq�\����>F�jn.�+�M,��'-y�����)ߛ7L(�����H�";��=�����e`��6��}�q雖<�n�0�4�+�9,��dXk��R��;EnS@VrXf����_/����᳞�sL{(�����/L�$!����b�B|��ƹ�RxDwS�Մ�y\��b
k	��O��z�p\.�l�Lg�^�{�0�~[.�a�5�dr��ܮ�0�����v�^�lE;�Wm2�k�*�#�E�1/ن����h�WGh�6i��N����S��l�P��������]�
d����v���E��������|�zH�{e��tC)vs�4�75��4�4��֨������+S0f=Ա��JH�h�rb��I�Wx�r��=��j������2U��e-��ݥ��w��
]�1̻��/qU��F���Ws��/R�I}��QXvf{ӯMk-�=<j�C��Ni�t������������&����H;�<�o�	����_��,jr�5e\�s9ۦ3w����ѹ��p���=��QM��!Ҍ ��٘{yoA�6-�G��X�j@��;�љ�b���S?RG��2�$�]�\.�����P�L��2�(~��@�b�P쫕ޢ�k���r����m�$���t]�<2BX��%�@>�\&�w]����!������-���H��Ek`�'���y��V���e�Hf�
Ķ��t�[T��t%��uӻ��3��s�sQ�/�y�H���.��7\�~̐�>�8!�أ8m�Osf��Q�ʆ������p�����ޜ�7�4��g����y܍��*�;A��0+�qF8��J~" N�[KZY5���or��c�nHˍ�nQ/�he3��w���c�ۍ�����'�SoF��,�q��1��K��f� ���J��Dr;��/�7��)�	2�-�FK+��,�/@��%;����8��b�K�ў�rz/��oJpEgfT?u�[�,��m�d=��3f��J�]g3�У5g��;�7#�3��U�q���#e�B](���������c��OCΆ+s25Q��ö5��v[䔥y(Pze}��
����g��N����y�,�=�ʄY�4�����C1��[}��g6fS��s[����#J'>}��i�(��om�xD���T��+�{}P2��b��Co8�!�
fIyo�`�i|=Ա�bZ���7�\�MZ&�8�=�|�
b��ƶ$��:�<U|tjA5׉d{�w{#��w�ۆ�+�(OGw8�:��/�-�]��E9���W�� ��c ���ܧ�d��3w\іz����w'��'s]�=�-{i@�Lp�3��З\�x�u�vҭ��H[��9����[���۫Y���!I�Mk�H���,Ԕ�QE���$�i($:4ְ����9�WPx��1,5�;W"k�NkbS�c��f�u��J|�ҋA�n�[ou'SN�`n�\�+)�a�����}�1V�/�Za�+;����{�Z]%�&�=i� �Mw�F݅C��l�a���\��þ�m�z]^������z��\��4a�"�V�h��z�m�F3č�7�F�*��M�Ƭ�]�� 6��ٔ���\V"��%u��c1Z����5 ��YX\$a�i]>sh+��<פ%��&�6��;��ٸ� �n����l��ݑ���X�-trn�#��[�u�J�j딅�\�q5�P��"�L�������V��s�u�t���U� e�z8q�݉cl�'b6�YnPl��c���-nm���$�h��Uc���A�e�T|z��?oZ�� ��B&�Ȕ�8�칩m��x�zo��{����ݱ��t�Z�]H5G'3|����SNc=
�h�94�%�E7¯��|iɕ������+�	�J����8D}�GWf�����-`�����U����{�ᡅא�w1�m\:�"�V��R�#��J�ǁ�,17C��vjH�_mcݭ����Q�53u�,�خ	�6R�2R��1Es#̢R3v�ݦ�p��c����u���=�n7Lz�^aV_l�Ю��pZ�DO�1c�RR�W�Њ���S)��:qc��QB����-�4�]��'Mk�b�i9�6XU��Z�О��u���Oj����o,LXm�֮ ��.~�����+��g���k��{}pm���|C�y��ǸW]|,�6��Onҡ/;��q3�7`6yJ��4"����ܓ�0�m��y�yKoM�LZA��$m�m�z�|l�m�W[Io^w[͆��0�n<��in�źؑ�-��i��׶��$�'N�� ��{Ǵ�m��}���R�ZP�h������d\lH�֛�uV��_��cL�x�J9s&\��<��8qHe�m�.ʴH+9Dk��*�WTL����T�9Ȭ����&�f� �r=P�
�t��\T������]����<��@�� �ÎD'AE��W ʓ��Zp�y˖!UERt��Q� q�+J�QZ�����C*a�bQ�79D(""�rp��S+�D�Мg(C	�"�*�H��/&�:e唒j�<�79B���✊iY*&�Z�:axXV��Bv��T�LH�bt�ZShL�4RL�N��㜚��y�y�$���hf�T�Br�(.�q¼�2)Qt��!�H �;��Je'B���S��8�r�:��'�����Pl�$,�Ks=��
	˧�Ey��z��;��l6����[vưLg��vuk_}[eц�y\��un̊��}ӹdW���d�2�\QX>p�{G3��|���l���Q��c��Atw;nB�3ת�^�5��uɜpnd�X�=q�Պ�����[<Ғ���j�������2����u$a��&so1ܨA`��rq���w�To��\F!W�+f؇J��{������j/,�K�����sV���y��9�֩����Z��􂈌wٍ!�k��W��?�{�����g�S�b��&:$S��~��7t�������/��!;��4K[<���<��x���p커L8*v�6��h�$S-x�;lݴ�zy���L����s�r�4қ�ڌ�y��4��=��y�$%m�ȉjݖT���k�P��xǟWR�z]3���p��;.*z�jm��z�޸h<6�!�DV3��߲	��eL��hW���*�~�Қf%v���֧`;�l��A���l΁iQ�1�tΞ���_��giCOn�%��g��m~��ݙ��#�Lc���l����Z�:��X�T�����n�^o��$����)Z[8zpJ%\��n��2�N��D��G״�ƅ�&e*���("��STb�hoc���j�P�8�����˖��0N]�bZ�8�>�Vأ˾�	��5���&�O\C��^/���	�32��(��
/�x�c�3	�YDվW�D$r�x굦�I(���SZ/��=O�2;���w���L����e���ʯ�`b3 �p��-��D����Ղg�q��s���1].�m��|�l���[���&��y�؊~��s��+�`�ٙ�:s���5VB��;@��K.ƪy��A�G8��n�U���B���u&�y�;5��dU�R�O ף��G���hҚ�Ա��l	�b�}��ܙ�����s)���R�6M�}633�Vi��; =�s�E���֞�V��}�C?)Z|��*����3̸�+xF2��E8&h͕������T�Xr�Cr����0,a���-q8��qC�*ه����z3^۪�v߅��;Y���g��	ʋu,��]od�Yf<�/�3 72݂Z�Jzk�� 6��e�yUq79|��<��L9}�EW`��S�nu�9�5E�B������1nT[D���g[VI��c��5�i\%�fg�~�:+���z�YS>ʮ����m�l󗦂g���@ߛ�]�M[-�蔠=������Gs��n:E���g��T[�:/��>�$[-�����Mup�_�i��FJ�bsa4=�r�Oc/�v:@�t�ގ�%eؖ´:y���.c�;fE/��u�o���xne�m����|6;���?z>}~���ݘ��B�L؁���%Z���
����hA�-��<Y;2Û1�[�8�v��t�mvtTe�[N<����v�KmVf��:0_{;�
P��m����5Bp''՛Z��JA��F֑�Zs��mO|�D���ɭ¦x#��̕����	V�{��K��t��#�ؿ��ds���u�E�Z�Unپ"�-�;�tS�[$(�gC��f��`�TSn��l̀�Ҷ{����sF%�e�-h�x���ݼ��z9��'�b`-�S?uc����wX�>�t�z!ߴSxk� ���0��_q:v�)��3���ı�yd�i�~6�q��we;ʺ�z�~j�-T+q;�܍�M��Na�����$9�j3�'��+�	2����
WK�h�Q	���vS������*�4��Q��3ި�r�ҋ�/�m��S�^Ra����%{9!�ۋ�F��.��Є��f߅K�
�;���Ϸ"����zc�6>|�\f��y�X��9)�	���ݎ����c2�v�a�1G9��z�1~]�� ���dςu�kȭ���y������R[��"��:K^�d�Eߙ�&�w�G+��h7�k^���q���wE�����e��X���`���h[6�V��`"D��z��r��i���:���VLH�M��͉�-S���:���d�|��g˻i�z�3�z3�*Y6	0X�8 K�淺�sڽ2N�c�y�t35���q�c�ه�	����&�I��_b�����IS|:s���A���{M'��xO��%���-�t���|������{��w꽒�U��T�9C@Oy�z��t.s��4S�Z���0A���31
!_�y��y�&ߜu�ͻ�V�n������8�[h�2�4�p����\b�Cl�~�;��Ճ+�g�P�kȚw�.;���w�Li-Q�'����[{T۪f}�F?KwSr�u3�gɸ����ͅ��كXJ�\�na�obiT)����W�w�����NE�D&|2�O���c
��{~��\���% te��o��c�J� ���L����cw�C���B���7�ed����bf�tsה��-�l�
۶��ϫ�T=.��el�!�EdC�[#�d�n�"���a�F��Mp~g�w�.�2���Q��td�˫]ߖT�ʹ�!����MxM"^��kv��ZNg>
~��AѱP�Ln�p�f`��xn�[2��t���j���L.�S�ۣ�'y�]��~�.�F_M�>�d��8!�ggOXe唱3¡�IJq���d�2Ln=C�S 8�ՙ=�ΐ��?M�kZ���Y���e�{N�[���2�mL|�]�Vn�����k�ol���z�a�(�/[�m�h�Y�⡸�����0���F=�3�9�U�o����e��_�&u�>f��aX�0��C\�^-U���1�G!4�
��Ci':q�;&m�ʍ�Ӹ~{0�|��K�ꎐdkT��,���s��}�8�D��]|�wћ7���w�oX�إ����Q�hd���qw���q2���Tד��7���N(ycW5m����;͓������28=6)�6��_$W�cͽqx.�d���e`u�C^�ܕ+n������O�����p�3�v��^V��8:���zf]�8�ܲF��Y�϶�uV�Q�Go�� ��w��)��3�;�Eh�|�^�w�j*o��.��9Y�������u�^m^o�����Zn���z�o���ҭ,��Vy��z���Q@��s0���ٌ��uٽ3�C�3i��D��	e98��ͻ�F�OW�U�q
�b(�;{g*����{څ���nu�L��6[.ʎm�Ze
e1h(��w�i�!�Z�
9��jy�=sb�S8L���;g��s�^�����������z&S̎S��Q�5�+�kg�}�^s�2b)fl���'"y߽J�7��D��%�9RHZ�af�������l� �å|�18�v0ƀ�����Nݾ����=J�ez��͑o\�`�9�gV���0�#/y�VQ�#����kI�������tv����$z���7F��kj����sڪɝ\�
�-�+��A��^u�PWn�G�q�#�̃�RuWۙsۚ�9��ދ|�C���n���h�@��5Gh��dD�첤k�!��(c70��]}p�unHɮSr�mљ�sSܬ�t��@���;�SLC�"�ӛ��\&�e�����^�kdLS��O5S꼬�g��ԇڈR�`���h.��f��Q�1�à��p�巧_�䋽����Ӥ�9�ܺv����*a�q3!���M�t�r,Ɣg$b��)qV���&�q��"H�:�(@	�܌�e/�/У�������%��/=,��s�a������q�<#�t�%�f���ǖ2�Y�̎t;���T�ÅC��70D�G9ή��lQWr��K��D��L�̎O-\6u����\$�O>���b�q���q����Px5�ƀ��SD���E��Qm�~\�u��2�Y�~����t����y���7c!�ޛ��Bَ�����{(�v�y�bЇ��h�X���Ǿ�VkV~�`�MC�E6���*��e�*ǲ��<G'÷ns{&��~��Lw4�vThnV�7��6�)�Z�p'����M��w5�ޏ��?W��0/�X|'�<�#�~�P6ٗ�,��6��M&��7�I��8d�w;E�J��=�<��0湌ߕI�XB}rW\�=�������UӍ����w �	W�9��|+�ẓ�q�睯6�q)p�ZVJȏ�� ѻ�����U*F1����s�h�=���[A�7��C��ԝ�Z�!\D�1�|�Q}��!�f<�:�!���R���8;�6�SeEu���Z:�1�^�:}�G��^r�Cz��J����̻�+Z!�-Ҍ��g9�sk�s[�z��uX�"�!9�m��j����x#�}n��O^f�hv��w�+9|�G��y�v-�[�4�S<�����tSzs��2�`p�أ�]1[�UT��&w�j5mj�1���!����u�f��y�(rl�	���:�%Ԑc�U��u�/S���-��3N��]F	j��el�s�߲��]m�f� �6-����#��~}2����WA����S9H骄_FBП���}��_]0yn�QLy�r���L�+c�u�-TMFS�6Gd^4e�jlJ�<'�e�=2��B�FO86�ծ꯮�<���g�AiDS7D;�cDCZ�\���qWǉ�~n�RS�)�r���s��֣4��(�w��c%�̮�w�W]R�[�[��s�5�b�I'3�gzbi���$?M���t�аKxe>��(Q].�E�� �u֦�'����W[1���q�����A��;/W��}���e�l�C���*��5�y#����7G =�ۃvA�usV�&I���)�r�����4]ݼԯ��ȯgK1���/iݝ�2�P���hzs����`�D�eh�%��x�zU��S��'X|?65TʳMP�e�@b#�̈�mA��lTf�tw�fu晸ȡ,�}��L}�m�g��o\f��ǜ��#rS��{oyMp"�&an�;d�E�g�j�WlKĮ�����n
�FW�%�׮{Bz���|��[�9]u�#c�7��+�λ�D��{'��WpX�v���nֽ�[����1�nnl���t�t�'ny���P�0f�*�S��������5��E���Ar�$!��ߡ���9����Nڗ��ޑ��}Tʚ�1Ez�3�+b� z�oB�ە-|
�Uϛ]����Uu��xevj����6��E�85�w��e�T5\G�m��p�n�\�mCÿkTM�M�T(���:��d٦�na=��(S)R�"��i����\BC�E:k�7�Y�z@��<�Mgi���R#�v����P� �B�,�]ʶ���h�����
\�Rve���k��In�4�����.�I��^	lݲ'��ۤ�[�FDk:؀�����bǾe~_en��]BP�]՝3H�OM*�W㳒���#ǖ�4�H�O�T���}h��N]]�4����� �^	'�|�K���]E
���Q`o+]R��=�j��%кlW��n���ݍ� G����8��ݬ�bǴpAP�:�h쳥r�o7A�$O*0�]�d���	�̧��� �]������Տ}%�X��1w_5�J5B��%�|�u��"<3'P���.���F�p>n��po�����Hw�>�"�1�����O�{�!��_B|ٹ(n�p�fX���e�('<:�	�d��e���n�������p��"W =�(���G�aA�{�U�Z�����8F}��dT��\j�n6Dv��^��~1m������OT�"�c���EK,�����9��q
��<V��VSt������盢@��_~����"|z%�'�g|��{�9��v�e�PӸ�v��ۮ�4�-W9Z1�\k���O=6���b�i��_$W,y���h��FS�L+�2%����/<��z�K*���X;��6�wz2�����m�Ԝ}�0��^q�3j��`���x^b���u��f~J���`u��=��]М	���e�t�!T�hU�����{��Q��xQ�;y���Tp�e� n�����=m�c�O�ZY�T�!�SJ~�dz��L	櫗|ƾ��Z�r姵7t�GE��ӿ��"Y3]֩ޭ�돐66���G���r�m��-펋�啬��Ś���'��C{֍�(�\%5����R/f���-n<H�G�����7]�ַC��|l�8�_T�X�ΔYv("~�E5�:��vjo5\���|ԣ4T�m�Q�,�!jrq���y�9k��*�8�
���"!<�fv�a�&c��s$��Q�e��{E�M�ݕ�v���b�Qm3n�4�s�Z�+q'��"��C����m����Տm���m�O>Қ��큰������)D'u��b�wAcƲ���u���7�l����k#���dD�_m2�*R�<���]��OJ|sp}�<Y�y��Z,���7i�㙮!;����CܴwS<�-��>��eL���lˠP��xǎ7x����f��쥦��C�6d�^��
l��C`�hS�]�Np]�B�5�,���}O1��=��w{�/���ٟi����HuQ
C��h����P*7�;�6/Y�{�:�������k��/;�!��d����g5ݔ�U��z�Ј��n܋�Q��	�����뢒�c����=ϻ&���P����b�F��t�;���-
x�qR�+���|i����1}�Nt��͆v��;���^�a�+�t��
e��E˼�0D�3b締�^���ᾢ�*�����vn�ə�vhQK��`����-X9�5�J֛<)�Y��匌����)�JWtm�*���.��H0���Lv|mR���F��	��r�NS���I��&c�r�Vf<�X�KY7�O������®�E�Z�6�w#�p��6�[6�6�Ǩ\�ذU�@��^�׀L\��,�_��`��er�����C�řH��D���N܄&�!r^K��<����z���ֳ,-�^�B���f0plX��ZԠqeF>��L�d��KaVti�]���"ueO��������6޸v�(0.o�c��w�n�V��[��Kl��G1k��OR�W�d�ceC�¬#.��Q���a"$��<G$���O|�®_EOoמmз�����Y����C��u��&6�0߲�yB�ozu�La3W|��Y�k��j��6��
�����M��G��h�e��z8%� 5�m�3S�725(����`�}sQ���U��p\����ō�Q��v�F��ʻXx�WL%kkz�Ksc��ݴW5N�v&q�Ôz�X���Eq'��F7.�ǯ,v��]�������������|_r�G�A��ֶ��M�mf�Y�ye��i�j:��ipBb���A��	;��`��W@�y�1�T5� E�_ZF��Ǧ	t����gݶ��r�V�,.W�v���.�LV��7~ƫ����cr^�<]��p��b֭�"0V����� ��tE�3G_A�8>��)��M�ǲ���߳����֙�Np�b��suw�Sp/�[�xjS�̣��(;y��Lx�_Lpp�q{�r�)T�ٚ�@k�^�Q1�$���)Ĵ7&�ЀL���+��c���h���|����E���|�S��qۓnJ���j`��i�}l�3oy��+:%��;<��}��u-�\MXa=���~��Tt�O�vr�di�Nfw�m r3��������@NJ�O���jwn���!=|Ӿ�^�XGl(t|�)r�)�q���W�D.-:9;�t�]5��ҡ�+�vMΜ�M$�ea)�L�g�8/;�Gmwq!M���4��X��e���Ư�#̊�ʉr%�3���\��ٔ�(�g����X�m�[�Nr��Ae
%���+�۹�\׳�od����j&<��#>�ɰ;�ˣ���H�JOD���>O �O.Z��̐�ݣ�=�
6�f��a��;G��"q��b�_3[���1�n�f ��n�Z��{���]��7���kP&�MRH�\~ut^G��.�i<=�G�	��/W,+͜�n������_xJ6���(����ر��;A�cjL�]�m&�<g�a�y�s���n�;drIm�ǝ�Yy�72�Gp:��k[%������+M��"��m�8���vaQ�����u4�H��y��X���xqe��l��
�S��VOm������-��>�t� ���j��g��9��#�s�ծX��S��9�;W9'r���
I�TES��n��R(����ǎ�#�.�H��J�0�Es��y���r��㸂.8ê�T]%Nr��J9�����PUDi�4U3-J��J<���i).��&���β9��eF��$�]�DIl�!:W�T�Ĥ��F�D�����8*&T\��s��,Ȍ�Q$2��R��(I*.,��a)��$��0�P���	���QE�D���J"e�:�e	'NV�i�"��D��I�lТ��uI
��V�R���T���*���maI5N�V���(�� ��!��gc#��+�/.�Gɩ�V�F��W2E��v@�L��a� ��W��`K��1�vs��T���՘/��%�����7����|���Kuz�N����D��F�y�̄=��ܺ�^rtrC\�}/G�r�]a3���v^B:�,s��[�j������"�Bw��]m�����!������pú�Oj���6kL�!����g��Td��k��lsŋA��;��LD��ݢz�M�;|��R����8E6��[�pC[+x����1	�=q8��g�A��"/)�zg���1�㷼�S�هܫ�.�-G�q���}�.�/���PCS,ǔ�@� �L�`��q͖���k.�^D$��/`,�N{`:|[��9�����﫪K�q��2^v
h���q�X��`l��{}/u����L��,�mW,��O`�����\��Ѥ�,��B,�ܾ87,,sͻ.�D�u�r-�<ҕ3��lC����}�I�8+�5\_.x���9=T;�j���A��8wHOA�r�f�~�(r�95���������<�E��I��m�5{��s-s%�l�ԩ�uGHOa�!d4[s0�>�<�`��6�_�����TN�I����3%�p�w7��N��7L�g/�.�pt+�"��k��Ϯ0s��:��Ɲ�<�L9hj�����Y/���TI����m֠}+-U�\*��e�������vta�ox�=�{B}ٵ�3/5��ӗqgH�|����TPO��B�n�ʙ���3ʴ%�zzy�a��)�&�{^��� V{fȍ=���n�P��l�I���Jvie<��uk���>W=�^�.�&7�{Z��f���:��w����'�$S`Hn�3�+Ǟ9�ؔ7�g�ߖ3�w3��`SG`ՐK��߶�]|��f�����-����̸��� c�#Y�,e���)���~"�yD���J1���7������R�P�D��My8��y�r���O�ƪ�
�fdҼBeQ8k����u���H�^<j���.�{����m���6�?>�\f��ǜ��"�`H��y��o!W��g6c�ߛ6����g���]�/�0Cc7x�� ����WL�=�<һ�ť�cK�81��]�HK��r�Sl�x�5�޼��W;�����c��v	ǯrǝ�m���ߣ:bf*��i|�ds
���
�wίl���3ުw�¦�l�q��]k����%� 	�;��c��*��nOq�6:A|�5L��#:-����'��*�6t.s�t٢-�a+���K�a�u�3S�_��������0G��=wQ�֎�F���c����e�B3�A<�C^!�_9����W�N�ݣv�x�Vz�x��X���l�13,g(��Zי kk�����7��r���X�N���fiu	�F<�����}�m=��G�2�q���]�~�(�t��ͻ�V�2�
��;zh�2�������h�e��Vf���]��Ez	��na{e�P�*]��Lۼ4Ɛ�Q�'����K�,����ю�=�I�����c�c�~������Mu71��5�4���R� =[D$����M�9{�����@㢧�멬U��~�R��4N��f��5���톡-����D&u���=	�c�lꯦF^f��Ooкrù!Ql�FZ�t'�=$�]�\.��=*a�.��dӜ�0�؜��{&&��q$��|�渇s���-�C�"�^p�$�+�k�Sr�pi����֜�{ɾ�l���[y�'L���w[���yk���m��<��/.��V7�7%�(v.�q6p�u�/L6�n����B�p�{Ǯ����2�ފ�|�fH~�pC�b���p��D�mL�t,���'%�G2�H\5���L�g�fu�N�ʣ�)�;�d�&]�����6e�����vIG�i���q�o� {l2Ꚋ�q�Lz%��gyf��3t���-��?9�v���00 �\U�^R�#�r��멹FS�f�;�B�I1P�m�4�P?zHdV���6�z�僔�&]�w�f�Pv'��U�85���5c�<}'��ë�]��ۜf���YA�N�!ڎ�[u�a�Զ���!n��\2�72s睛��N��k����Ѯ##��c����A�5W o��/�)�x���BF�����#� ����F��h�eb�vX���
��66�ɕ.䞜���)���P��{y�:�J�x�Ek��_�rB~3!�z2�\�1���Q���`�{>�.�%M�R�N�UM�;�w)���K�5��)�6�~K&�����Ϟ�M�c����ig�R�C�����>Dh{�a�����+[u��g3����ƥ���6�oeA呀$-�NN873n�7�z��c90v[��i�j�+���*�4�c�G��r�(�-s��pcM�%���hB���|�B*6�cw�\g-�Nx�w�
 ���V��Տ��af�}�5Eӹ���[�_�'V!�<�L�eV8k�2wn���D���I�w�PPS~�dD��%�9RHH��:�u�廫��5\�Ax�r��9a|Όn(�Q	߶!�մ%L�ꅣ��Y5�,�OQ"�@ �Z-�1:y��K�T��4������~f̭�rb:B>��
��0������B�5�,�`Gk�ph��^��<��s�h�����c(��N;�4HV;9ǭQ�-܎p1�̃/�Ct�bkVp��I6H-�t�l��]��ܴ�^5s8��ovAʵ���݅�}Ց�efuR��8o$�	_P�-X�����Ρ����A������p)@й���U̩�ɣ�����m�l���t��S���U/}Oy|X�2�+ɇ�f���d*;�:��u��2������l��S��N�h�|�3*1�[9�n�H�nƾ�sܘ�9��-�t��Q��O�L�,z�)������J=�V�m�&s<ٜ�+k3�1����ǚ4�L@�;��^�X7.��B���J:r�N�t]�"r�tP�k��[~N�U�K*����u�F��,j���̄��yƊOoo��]�2�}9-+h�"g{y��P�$���pW�!=�E�����	�	����7p��nڷGN�ɹ��۾D;��9��d���X�� ����d�P�Z�pV(|�h�Y�U��s��[s�5�pw�L���C>��Nh���i��v�V�o��9�p�V�?��
c#��zu���(���͙�v�ƽ�wz§�A�8滲���1ee�=tE��hV�~V�?�;�:.^�����f>�.U3lç�dz��)�7:�X�Q|{j��/�u�/�װ���F4��Z�[�D����)��A*@�B|^T5���3��1�vM��IR��kKҞC���8�w%@��bކ�!�.�3;�񗖺���S<qܨ��=�m�@L�V��lI��y�A�o:rc�,�%�'rs�A����m�2���u^���u�	���Տ�P�+q�m�'</ĩh��]��z����W<
EKƆ�jV�j�5�qd�y�=�WL�	󠪟�e�7���L����o8N��܋ �/d2��;\0]�f���Mus���)tG�9�a�aJw�_��k��&�g�-�ѱ�kR2:]fE}��~��!�u��i
9���E��m4�>�D��������Og���|�a�'������$(���-]T��ǥE1�a��h.�5>�<6LL��v�H�$��ݺ���l�i����,�7CI��Bّ��p��u�W*`���L����V_mh�c�E�zNs��5D;���V�={p̶xeb}���,��!j#����ws�Gwr��aL?i�z,���+��ٙ��r��m�!ԳWN@���s��/��-�VK�whۈ��N� ���B��VGAM��oQU�n�K_��{	E����6���t��h;��=2KF�v��-�\y�h��~eP����L|�ߣg���[!_��Q������Գ���*Ռa=�~�y���V��y�Y�wH�W?JV]���wo�c�6B	`/MW��Pf�V;'y ��x}V�C�[eO?zO(���	HW}�� �=���1ݲe����4ى���껹��f!NV&����/�sv����8�]g�<���Y���1u����<�w�*�.Y\���-]�'�S]�ς���--}T5�X��k�)�(� �LOes��Js]�V�����7,y�A��j��6Q8Ng
��*.2�v�6(w�[-ϒת��ՅVp3�8�[yQv���F�h��x�[������ ��\�<��|1�[u�Q+���P�3R�2��z������u\���Ѻ���hs{6�k�iɂ+ݐ�*S6����w���eMq4���P�`�ѩ^L14�#9>��W��3�=��K�7��Lx� {a�*a:ۙ�x��}Q�'�V��T1�zH{�Ӷy<��e[�g��2����Q�L2�a�l�M*�{�˺؆�N��2Q��˽�3��ӊh;��6O9��v�Q���^8��v�|����4�!ɉ���'hE87W�#oo��t��t�=�;�����F|n�	�JBۆ�.�o�]F���m���O����~�m��K�1��,˹犴e�*x�� ����d�N�p�td냃�y*;)��4v].\[&�[�Oj;Iݢ����u�,ٵB�|�,����n\���ԙ"�T'��ĊN�ѷ˿J�}�-�J���bߟ��[��g���6;H�y�}�h����)�|�Rwo圹@��w+w�϶��YT9me�\5���q�'\!�[���?	X�p����?�p���ކ�tm�����a����{0sdE�C�]Rə]OHz�)wDoEO>o�$<H���c�l���\���"���C,ٴ����P�74�t��S����pz:}��#-�*Yez�0.�X2�SU���b�:w��l���H��i��k[��W��_"��3�.w�b��8���	���e��k#-��F�ª�k�:+Tk���K'���zl3!�S�m7t���7+y�}&�d��\�|
[5]N�j���Q �挖V*�7M\͋u�#Xl�w���ǅ�}l=\���|�WQ���Խ#��^(�~Gv���>��2H����W9Lj�e��w������˾iz]��YG�j��\fg4��|�߻���oe�[;*4r��7�-��'���
�q�؃������hk�YU��G\��g��'���j�����ԍǲP	hȷ�[b�x'ݫPk�]V4�H���͑�^�:�-��o~�S�nu�L��6[.ʇm��2E� ƹ�;2�e�Em��pt�� ���~l�{�ܮ�B��T�Ս]��"]r�4(,����"$Z�q2�u-1���>h9z9c�]u��<��)���u9�������������j�Oa�2�y3�J����z����u�Nql@kr��w�A�����	�j�Ǿ&y��y�4).��r��e%��wFHM��y8�GnѾz������=��>���_�;�,���$Z׎s�ݴ��1�C�e�B�Ƣ�s�"Ɏ�����S`����@���L���u�"ka��]D�L︄f���n�oQB����'^�WSSv�@U鸗t��	����f��N����0���H���'.n��7͛
q��h��}
���<���!��G!Y����7���do4竵'�pm��*��\�>ϱ.�#eCR�<.�w5���2�Dm7L��Sj]ڐ"V�LL�-E��4�9"��h�gQ��O$��̣��Ŵ(�y�gs��,���&����v��T3����*��Z��	k���S�p�{�8.�9�)�\':�m+�g�g�V��U��'!Ȟْ�lE?`�k̖T�y<���,�KmT���28knU�PTn�k:hH�ۊ�Ū����fq���H�/ ���8*2�t[���د`\�|feݤJ�q59墅fe�~WOn����g�����@��Vt}zU��,��b8;qaF����C�1�ֆ�޵�<��!���oم=p�gpQC�̈�Nz��`�1e� j�Y�d��9���գ�5N��$E]��ƾIy���,�H7d�����c�J'��R�E�d0�n�B�{� 7t��h�j�WN9��y���с;�B�=���{ϕ�5�+�3�]�˧4Wnu4׳���Y�[�`���̗�������v��}����'{(5hX;�a�l��U�'w����E�N>�B���CY�)�L��jf���;p���{�-�&��=z�1
��U15.�m����~��/�[%�z��8���8�ƛ�]\�d��.�'=��/=
:]�:�Ոז�煶�e,���_t�,5�ع
-t�ڢQ��{~��ML��!��.�D�u�r-�L���i���)�;��[n./�]��ª�h��������0[p���s߆���}�
�R�٦a�}�R�栿�rYF�O\�6_&�xf��3��u���� ��̗��b[��2����	�!��f%��m�n��xo�W�k%~���OE�C��B�!�''ѓK�|n�(t[�|��`��Ң�o�9������4Kt�թ�=�����i�i�=''l;�.��G�3O�b�.S�Jq�iU0��o���F�1���c�����1��lc��c�����co���6���1���1�cm��c�����1���c�6��6� c����}1�co��1�m��1�cm�1�cm���1����1�m���1���c���d�Me#�M��f A@��̟\� �zP�EEP�"�����TP���Q	H�B"�QI*�
�T�PH � %QE"��QH�U*�j����+�T�P%*R�R]�R��I���i*�E �R���
�������)IP%�RU(��k(� �㯼=$�
(�T�UJ�!D�dJ�B����B�����m�*�J��(�UR�QR��JD� "��0��_m)>�=5
�(��  �^Mj4]˶�*:����kMNΆ��kj��b������S-���]h�j�j���)M����]v���J�JIEQT R��Sx  8ݲ^���Zփ��U���QIQE�.QD�(��(�+�B�F�QE�7QE�(�����Q$�(��u�QEH��t�4h�F�(�ꢵ����T$��   9ɡ\a�Z�YD�T6ʔR�ҵ�N�q�����N�ڹ��tQ��A+m�j�S���WE��6����n�DT@�(Q@��   ���ԫ�U���ån뫺Ժnv�d����ri-s;v�\��n��.���u����j���kM����9n7:�w;cv�8ƍVG.��\.ۺ�n����*�E�(
�%U�   �U�Q6f۷U�5�'m���U+�ٛ��c.��;�C�ݻ��ۘ7F���v��43���v�k�]�V�kL.k�n��ҵ�rvK��n�*�qR����U��w�   �w��iu��[���j���qE�Pݫ��6;����wu�Z��%[R�54wk��I,j��g]۫B�k��7K�j�.�uÙik�]�7v�R�R ��H�;�  =r��*��]������[�E�i�v�]��7S��Gn��Kvn�0�ڭ�j��r��j�\��n�Z�U��WZ���s��uҶق\�ӫmU��R�2�$�JQDG�  �m�ۤ��ꥵjj˺�n8�u�v��Zݕ��v������w-ֆ���掭�۝+��Z�N���ۙv��[n��S���T�w�l�K�51	)%R
K���T���  C�zj�Sv;����][�:���-D��j� �]�2��T�MswkUw:�]sSv�����[aR��gwu�jv��ٖ��;�n�S��D��R���BD�x  ;����k�l�3-t\����m:��θ-�u���Lq�ʷr�7m�+�5ݕ�;a�S�P�\�v6��[vZ�v�W��e�i��� ��*QT0�x�%%J� �U?��BT3H  "��	J��@E?"f*��L@4�a&�@ʢQ��پ|.�\�qo�U�1�'�,��7���ŷ�^��޼��uם~ �$��	!H����	!I�$ I?XB�!������~����_�ӧSZ֎�z��	ER��D�q�S1Mˉ���r��kk(�aZe�;�Vj�{*�)Y�/60�cU��ڻ%��3��m�5�i��M,7z]$S����/E�ZeE�תc�U�³(����0��`x���J��b�Tv,�b����fՑ�RW�јJ�����ec2�B(f/d�P*CF�������i��C��O$��cҢu_�\�[�'/v�%� `bg�Qf�^�fA)͠,X�IV/٤Y��P�iz��%�wv6��H�v�u�{GL%)t�-�U�p����m�0i�x�Lqh���*Ma���*G1H���,�H%�%����n�	.�ˠw%�Q�TX�d�ʬ�3!ZI&��ի���j�Wgj�f��Z�Z�Ca,�B3[m�7l��]��fKUz
��q���V@T�m�61mf������EY+k�v�G�(ܓd�M-�V�Auu4-{.��@�Smn�f�ŷ[I���S���Q,�[@�)������A�-��b��;�(u�b���8��oh� ��Ouw��Ո(�٢� j�EauM���t����O46��r�է�Zgu�Ed�(�L�V�']��5�֒�摦�AP�GӉҏdݵ�u �Ѩ�I�Y���V��7v+�R��V$N�MfU��IX6�SF��m;�쪚,��tj)Bb�k6X`�B�W��!�jj���E���i<��h&r�ѯ`
�L�L�^���"�Fw����`]"��if��Ă�՗��
��`U� ~ڽ),H<�����EjKl��D)̰�*;�h��Z�n��*�ߞf%V2��GY�242�Cn��JB�Ť٥n�{c	�<6�9�n��ۃ
^P�4S{w��9.��hM����Ю��������w���1<2�U��YOf���z�O��gk1Pv���裻��x�u���pԀ�j�w��j֍N�=3T�t��ϓ̍�,�p�V�@M�*�[�!D�Ǔ2Vr�F��(kE���w.��	b	�!b��S�s*̈,����n[a���Ѕi�m5��If�
���H+L�Y�,��d���僷L�T�ݹ�K�e�����Xݘ�nS�`�>���T���`'�,���BeE�B赭�q,�Ӛ&���VӃ���F�����H�)�b5|cт��nˇ4\Pf@MJ��T��nS�j:��Ȫo)�l�p1kj/�H�p��5n^�7�)�t.ES	��-��YEݿ��5Kr��u�a[�}�{i9�1ff�K�Hf�ْ�7%�@�b����Z��6�u2�k�i�����ɦ���M�N�K`��6U��ֲ�rDe
�6e<�Lm�[����~C-¥ێ�C���AV�(�z��+oF�ݽ��R��^����.5܅`�ƂM��n�nٰ��`�$e0�<�{t�$�i����m���a��Cj7L��vɢ(ِ�M�,zB�a�k�F	�l
y��5Y/C?Ln���I<(֯�MYa�ZΤ�EhV�i4�����#��w��AJZ�n�.���ͣpcO,J�Vr�͐�5ch|���Z_]�.m֣u�Jf�MKU���rVar�Ce��wB#C�i"F�Y��Ќ�Cr�2��a�*uz��4��ꢨJ�^G���o�nf!$úM�2��n��9�v��"�.�8&`d�!��� ��U� �Q9��$hDL.��յn�E���X��մqGa����2��\�H���ݰ�.�ů4�N�f�{&����C(ʍ1��&��v�l���4vf�[1Ů�̳���t��v��7� �Ɉf�h�b����[�A�WP�Q�V��LB6ƪ������K[B���/��/��d�(ɛYM�mGg1�[�F�ח��=f�f�nJq[��d�������7l���*ݣG`�Y��/u�y�(^hjt`�.#�u������n�<I��S*��wkr����1P�Q��/+A�6�.��ΜH2��n����ԚZM��S�Kkj}f�&3@��h;���ɴ��٤.��{�1��&�S)��ҥF��U��4�w`��mf��b�+�B�heA�0�9�9P;�E� �L�&�w'�n�z�.�J��9��B���)6�V:l��;�ԡ�_�-��ě$Y�^���ӭٙF賍A�FZ�{L
�ZD���j�WpŤ��3G.���YWFv��CߎǁeJE�+!02��Kkj�,ɭI��a�˷�^@�a�,:4o(��X���\ M�+A�ڼR�ʭr�U1��(e�%)Gi��� Йq=[�p"��kr�c[�bX(ދz�)�7�	,�{`@�C#0�l�K��i�wڥ���L4]<��t��z�K͠��.��ra�q��5�b��V�Ѣ�ڍ*o~u��,Z�g$�b�M����q։�m�p�g�z�!���IH�u��%���If�9#XfG�R�It�(:�2�mԕq�[V+d[��٭"7�ᒷ"X*�=h���P�~v��Z���ЀܱF���e�`��2ӫl˳���uC�@X�MӫAe�6�x�Œ,bͩ�8YlrVK��Z5%�����d戵����O!�c�(l�u+ڒ� Mn��
�j#�1Z6�^�+B�Q\�jĕAG��[�o�7V	w��j���W��fv+���	q��j�t@�����,�&��6�cx��]duj�p���d��A��-^�'Jq*����I)�y�řKP�3U$yM#yx/n�Y�f�ͤںx~I���抆ڋB��7i�@0Z�Z���tѺ5��aT��_�eS�-i,���0+����e`c�p����/P]�)�a�I�9A�IAP�b:�}!X������pw6�9Fؔ�&�[Y���ڳ�hF-�
8Рd�Ssa�B�m�Ď�J�qNb�F29�.�5�8�%3j K�
��,.�Pl�-˫'e�R�e3��c/E\�BԠ�C*47{)R���f�����[�WJ<h���1��E�˭�B"hP���vAse��{�Xw��-�Ɨ�!�F��nS/�&���l	1b�+[mJ�u��-����!�h�Wh�lѻH"M���nee��a�mٚ�!%xw#T�7b%��V�$�B��Y�+[�ělXs�Ĳ�)�QZ���q��+ז1��v�d��X䬷��1�d7&� Q���Ԟv-�6U�6�7�G`�D��*J�2��
f�vi�-Z5����ѓn�®�fI�b7�5�MHg�i����Y%���쏍am"J�t�h7�B	�6������8@:36ѬݗHn��¨V����Q%�%�{�����vᢷ&[�� imX�;k"��<q!��{O�u��7.�ֈ��ҕ�̫�pJ%�z��� P���n��F �LZ18��e;S(��e÷�h(*!�On�;�Y���N�UN�^Q̈Lu�꥖��i��fB���ɘb��%J�)��x���YYh���)�A�ů
�h���/�z�@���p�SF�63s*�%N?���bYxo�Q�!�85w3^*ݱMh9����5&�e��5 (#��M�kio�B�Bq+��R� �fbM�uԵ�AX��ۨ7rS�%Ǡӫo,�=6^Fd��m���QX���4[�Y���I*��2I���M��G֋u`^���j��+��R0�	[���-ʼo�o��mFd��6 ���k+%˫Zw�P����TZ�9r�� T5�t`���%e��/B-��e��$�3�\3�[�k�,�+i�efI��u�����^:�Ԓ	l�)��*Q�R�����A�*<�o&�${D�׆�Џ L�//
0�:��6��P�֐���f��<����^�p�^��p�G+.K���"nCk)�5jbU�a�S0I56Ԓ�*VR���ۋU4ـ���m��ahǁL�R�n1	ve�n;���+7uOX/�,�i�X"A��Ы�-Ay&Q�[N���V�F���G�����-_`h�{�lݗE��k-�+Xxu,�{N�0
�2��E��+]=�t��Λ��	�c5�Q�����7�4�S�r��t����I��:lj�{�7QS5@'�Y�K.�;I�)Z`��V�F*��) J�`9�˴�I�����
�F�9[�&VX'5�:zL85RQ�(U��@&k+�8ԫ4�K"�l)��c!r�u'�B
nl�>D
_��G�N��h����)��ea.��t%m+���BZ�<n\��:%����jmǒ%N̫(KNc����̀�j�F�2X��:�����rdsqS"����{Y-c4*#vjd���r�LVޓ�Z��:�36�MA����R8bJm�y,˹����RJ�}#�%�NP�u�DH\R��wCxO��@��q�Q8ki��`���,Lr��C����r�-
m-Ov�sC+-��&q	���	`��˂�dc�Wt���M�˕�Xst�yj�:�j��5f���	�)^�/��2]�T`֔7)f�=��"o�m.�WHT��m^�pe�ݭ��f��u�u�p�9v���0'�e$�`��"{o:�/Z�^�YjU˦��.EN���Xλj
��v(���V�lv�R���
V�64�1F���r�� �cv��L4l�m��h֡���b�L�"<qc�z��pu�Y��&Ղ����{����,f�J���	�̦u���ņ�=Qc$Ӥ(�βK�	M0��CoV�0Xx*�F���� �j����7���I��Q��ą줫KX�ڗ����`�L��	�h�Tn�H�4;�����jp�ci qE0����e&ɵL^�M�ck#�H��3h���D�i'&�v�F��rA(ө��Xőt�j�xД�����X�ݑN̔f�!����:�="+�z�T� x(�l�7�U��O� �,��ZC�sr� ۀR|��F�O�R�FRw�2�e� %��mV��FA54��m������ܨ�us	Ya,���CTX�R�u-���e��'ong�I�~�B2�'��B3<Ui��_9�lZ��*ģd��n���c�MJx��nn=7����Ofj����*/,j�:H��Y%ܔ����"�xpX�U95lW *n[��6]挵Y��j�xRJ�z��hd�B�+iռ&�Y���.��Z7%�����B{ES]f /r5 %�b��R�ۺSoN�V�V�X��� -�nZ��*Wn�J�]i�}�!�@�3W�����K֐ͬ�(;4V|o��s��v]��J�=fU���ҋ%')5�`�D�SM@G�(�J�ê��Cm���Z2n�s(��]e�4ŭ#iX��zn��d�Zp���KpD)8EdY3tB���V�����,�D�V)jn��w��W���� �� ��jyv!�+��,�4�[�F�ky����x�dJXr���p
��wH�G{�&��i[���)V-꽻T�Լ_HiM����֢�WV7F�h�ˎ�^^f'�V�1�Xlc$��I�0�A$�\���n;b�o��te��z$��\��P�%���4�㡩EfRvK{z�^[�4�t�ݣ�P�a�?h�.���Nh�ژ��i�eH�ŗ�+P��Ϟ�%����n
`R��Hjuf���ElǠ3�D�I7.��t"��#k^�gNy-QM����yE�	{6�E�r���^�	w(�l�uj�W��Zl�@�2�j�%9k�W�h�5]<���
��1���[f��ULP0���4����e&P�sJ�{tPH���6��3(%�9a
2f��vh?9y, ���>^QT.,,@��L��+y{Sq�2��T)E"���;���OZ�n^M��l^�x]�[[���p��ejW��U���ɂ:p	Z/I��&�v��+X�n�MkRc*T��Un˱���Z�4I���l���6���ofY��E�Ih�.l�r�V�v��2>�D���A�Ar����Y�Z��ƍ^��ӡ��uW�p�7|����L���8����w��+n�vjoͷ�Rt�j����g9�)$�u���-��Aq��́7�Y	b�
���Sq�6c��RQܺ{dE��ֈ0&&���A�m�5��+å���n�	kh*�v~1������=yt��X.�;��!�2h4%HY�m�N�f��蛻",!8�<��i�"�#��E�#6⻷�*�l�`����Sm=H�!�o*���2V�u@ҊX2�fmc"�=G�jR#l�i�ا���%
wJ��2���di����*˱�g&��D^e��MV���3�-��o�q�TM����!+u�%b�1r�(����Z��Ƃs q�"G��նi-O6���"ur�e/�{��X�b����8�D�j��SnL9{-\t�Q�i!���1J�Tif�$���V(���:���E!PPR�˛�e�zp��#a n�F���Y���X.�%7�*��ax_d�m^�˟2Ƥ���ڵ!���.�;x-�"ݝm< &]&N�`���j�/�ؚÖ�^ӄ�;�W��h�r@�rRƘM��Tme^��J�P��f,ct����4�.�u&ހ�c�f.��dVLVʹ��&�q��f�C/(�p�@���Yي��T�A.v�ut>ͭg؆-i�[Z��C�	�qaAY��&r�ӭ[?������^�j���޷��77)�\��A�*�Ӆ+�)�Ղ���;�e#�p7O{2��b��z^c�'�Ŕ�I�
9�t����m2<���D=�0-��JDn�R� s!V����`(Î�$r�
�[�7�u;+��ڎȧ��DҾ�ɬ����e;Z�w�p�W�B�*��7:�����vH�^Cecy��{�dh�UWut�׫F�th�NQ� ���(te�\}�o�L�q�Mnݫ+	��n��u�k�����*-�oe�e7F���*ۃws���k_G\�;��L�\��Ë��ۡA�Ҍ�|J�y��(�N}�muSW�q�w�����J��j�6Qf�сg���/=P�4��zq�-{������쭍8�@ģ���Uλ�E��rA�sù�ӓR���3W��j᮵�%�ᤩ��G!��.�[��`m��2g,%4`�Q�Y<r�Q�tt�j�8؜��7R�n򬁽�]��ael"�0�N���)�{Fs	b��[+�Hkuet�u�lɺ��v��D�ں���K4�oCrT����I!�3$�O5�R�5��V�֌J���}��w�8`Y)�Q�������%K ��4�=Y�/���U���7	�FT C�hH3o͇����g+Tw9��Xp46MӀ�7t*%�kN\��b�3/I=�6l��dt�������-�E�W����8��Tn�M���Wk�7|�ډ������v����ޏigj4�Mˆ�PYfq}J��ͬE#�6v��e�v^ū��m&z��҅�1�5���&�l�*���`U�;Y�:�.�LC���5�A��oc��%nN2���ZO�=���}r�	��g��mY���6�@j��nU��|�_U���
{�p�[��D�&m+�4�����ɗ��^rF��VWn�E`�U(L�Ӿ��FAv�*�/�<������Ą:�����:��5�A:�hZ����6�5��M�4a��Y�dH�Ʃ��8�˼(ƻǶQؕ��D�Dn��\��:����.]�$�1`qY6z�3;�w7�t�\2��S��*�o`���\Ma%�1�s�R�u�����!��gN����I����_˵�iTL�Ê��K�:�u���;Z������g,&�[��;�[�$�X�yh],�3,�

���UӺ?��"���ʙ
�ߚ7�B{l�,�z횴;an�	c������7�e�
EwL��o�	��v��uw�&r�AZP��}K�V��סl�+��w�ִ[7E�q�Ğ��]�t��j:��<j�N�}r��"�u1EY��p-�Ivf��`��km�Y�����\�����r��G�)Qnd��c��T[�ףS̡���%5�^J��z�=�>��V���}�Ѽ�@U�2�'���DT4K\��s�.�w�N�d�u��e����n����qV>kY�e�׎��a��H��'ׄ�B�����t��}o] �k@٠.���}ge΂̀�V�JW�nR�u�X����6��"B�ыe����y�.<�+MI���X(-�%vl����;&0�>G#����3D�̡>X�f7�ԍ��caui;�E֡"a�ͱ$49f��p��U��-70?<-����-�Mp����J鍊g;p�,X�y
�Ҩ�*����zc�]wY�U�Z.�d��!���u\�/�vghR�V[9� �s^�cy�\ʆ�2�������Eј���;��;�� �Mf,�3˫�m�TÔ�>�ǆJU��j�Y�6j�>�Wc;�����l<3m��+�4-���L�y��
�.u��-���G9�6K�s��v�$���ڀ�{7��i���iK0+�Gk��8�+o,�u`� :M�VrtU3	۟m�0�EP�.���,�Ԍ��Ker0�����2<�^��2�S�2Dd���$#��%���H�]ZF��ӎ�}n�H�w����0�b�Զ�>�jqM������)�7���w`�R+��*������K��:kR{ו�����[��x+8m�qkW������h�1˥�#�]*��=X�C�9X�t˼��S�X1�C�.�Am�2�)w`�d���SW:ϕ٩Z������j$�\G>�ϴ�F�=yo.S��=�˱���N��Z���]�����T�;`<����<KS�nˎ��i����;��i�N����;f�&��X��oLgQ��ِ��ќ�x���Y3H��V,޻p��:Yw%3P�`�K���b6�ENlct�Z�nd��X�wE��g�Y�j��N�;r\��s�Ѧs��t�ї��l��f�X'!ӫ��V����8�4/*�˼똩&r��5�qn�k�pe��<��6��L�z�4�QW;��	a}�v9�.ڄ)����yԭKG[xo�㖁&�P�^�H��N�T�L�A��a|�.��r�h�++U���52��t7�.�]�㧝A8��S�$�rծp͇:+�{/tP<[i1��v�vk����i��$.�%F͖>�aP5�����p���w�	o2v".̹m�}ܦI�s#�+ |dV�|�>�����/oLQ3�8e���Vn�JC�.o�97��O��8⧡�[ �2:۰�����ک,�if`��%VH)n�ԶR��*�U�@��|e�Ummg	��\�N�˥�\�K�r��ǎ����;kڢ���;^�n�]6O�wA�-���|/yl�p�u%�Y�]����mEtw�A���gw#�W��\�v0��34�w
�N�Ѽ�(q닲�쀷��!�sEZ��9�xf�����V�U>��M�x��B�N阠�FW:7��T��Ԟ�(�dQ�'K�`[[j+8S����vͤ�G��aC
��VA�e$��롭��PDyɶ���_z��O#8��fas�û�.�|HU�6�9�V5�^>���U�R�W]*��w�qN$�.�n��erݗ[�d�&�'��0���EO{���Ӧ�WWX��̒���g̉$�:j��|j��ς��ϲ��^)�)n�`�2��y��}gZ;��F��z��;^i�%{�Ȩ�>5��	��D����Θ.����w�=}���-m!7287:��]܀�ݷs^�d�9��bhu��,�]5�dM][�>�C�b�dl���F�v�K0��E�_v��]��dW�U��i��)+][��m����)t[�Nu����fZoi���Jˆ�u5dY�����r���f^����)�[�d�.�%̫�/4��t��/5`�	�@�z���ŴI�Dx��+b�Tߎw^���>�Wll�nu �' ���D�6�,�{ 4�b��� �R��=mf}Ҟ"��]N������{��5�]K�9���[�M�5wM�gbU���И�B�*��j^t|Nv(�#�ɖ�����V��%� *����ݍ��w[�pӠ^��V�oPC�;(�q��ܕ�2�n�-�h.U}�bg"�Չe1H�2�;�1��X{���,,٭r�.����4 ��ˤl��ܵ��Ӧ�����t�<v#�k��2�!W*k�h�ϒ���M�^J���	L ��|�y�ˇ�8��f��²�
J�[�o�F]����]YЇδ�Y�Xl�MR��_u�V���L�7��&��ou�F�l*�V�Y��h_������X�c����[dF��'R���Cqb��]Ջ&�.Q��ʔ�agm�����<�6��s9� i����i�g�1Ljq�{[XE��،{��X�ԗ�.�Mp�h���EgP]��<s��r��q���Usrm�����2�;a��.����<KWa�r �ȚG W�t�d�L��X��^m��[�K&��}>�Zj���v���]��t�®��zAQ��6�j��V���Rm��4kF��^�e�s��jO�����$�ם�L�ևBa�qY�!��)vV�"�H��F�;˯9R� 3�7�wh��]m*3f!�»'��Y�����Ԑr�T�%gWg(��溯6�����:Q�KE>E��9�ՇCj���V�m])m��lWv=u���X���RS1���ĵ��H|���������"�$��;,�b�'��ה�ݽR��PS}B�FX���z�6�h��m9��sl���I��o�Ӆ�G��<����cVR��uv�M_Xv�> M��'��U���^�w��	���ڀ�y
�D�B�eY&��7�YVﴀX_EذMO7%1��!���>��_c�r*U�y��k��l�l��i�Y��` F�\��[Y#%;��79r���m*�ĭ��}��;�r�a�����@�����t���pP�N�v��ٕ���������������S�Zu�(r�S��րB��.Vd��:5feLNA �G����7rfun�A��ky�kSf�����nZb�[7`(�S5}hӻj�}ف�X��u�
�=K�4b[.�Ge��]]�3QmC�׊@˸WBV��ś8�.��X ��[��`4�h�����y)����4�� �c=v�H3!��L�pr�G���9.˾T�kq����r='�Fɰ`�z'��Ξ����.�ҫ�g�o��`��,���]i��J\+u�oh*�^^��5.r�ž�T����S�Wk�w'�������i�Be�[��٦��ܺ��a�|0E[��e��]�������_\�O����+�/f�X���t�b�;���;�1�ö��f�,��OD)���V��d� �u��K��uV�W'%K�}���"���s������^
���%���'�ogV�/��)n���n���2�bۚ��0�H�2�uo9jDv�v��ӽx4�E	�L�4���!t%K_.�:_V�HQ�g5�5en]�s����+J�2�|#ywx�Sq_vg���JQ�ev�U�:ohÏ��3sjF3jM:��5 w�\�L�Ve�n��6�/�b"墻l����o�o ���^�ܢ:r���srd�!\N�&Q����O��{����N�<AM��)���u�&cM�� ��jg��̨6��j"�iv�׉(i��T�y��4&����P�6�?>Vy�f\�%.n��J��-�6�ڃ`|6��5�<�:�M�}��4j
�:�B�2��	J��׺��Nv� �����!{�"*��N���}V"4���aG��-�gdZ�2���P�������<����%nӄ{.�w`-ͮJ��+��n��S�i�J<�L�-�*�/^c]jk�X�sS�"�d��WV������C۸l��>�s}�κ� �/omWsN��w���L��a���"�ˊn+��ɼ];4�<��鶪u9������Tti����%͚�v.�чmv�S�
��C��9r�/�Ve��#KR���wV5��3m*�i��<��n�e�4o/!
�A^=��3Cٸ�<�2���{k�L�{����C$��u�"�5��b˙C%�!�vݧH��^���N��f�;���@���siK��`�cʏyY�b�c��Q�dw\�c�q`��N_^�-��P�1�(Y�Fҹ���C��n�i���Jmշ��F��ڹQ�L��٣�P�۸��)����q����ɀ�50�#GЪҥxs��H�|��p��ʚٕ8��l�'�mw��vE�ͳL���`g�%}��w,�r�l�_	,l$D���^�c���a9�������	��|����,Xyg4��k�
��	�Ma�ԭ�7�M��PB�z�{�����:r�fJ]�u���Ev�`�*�6@Ç�qҙ��HA;%N]X�C�y#}ٔ�f
Ca�e�؎^��uoG}ϧ^�_ujI��I�k���:�;��|@��mwl�r���9����[QHT�L��XqYU�Բ�SG	�����Ee+�3)��\ӻ}�)��a	�=��y�1ۚp��M��V$ק�φ�(̘E��e�R�����8�����*6����z��S�:�|_�z)�r+,�H`��޼.=@�*FM�&	��bt���%C��ڍN��QaEq_j��_n��8P�t���iN��)�#�0z��o	㻰���K����a�[Y/p�}��G:���l��R������<ýT�kk���Ɉ
��Ά+�Ɏ��T��5�^�ِˊ�㏆���Cfe��Nw�o+K��bzTH�}��5��/��u�Z�1�o��D9,�EE��}S#ʖp�]���Ua��Z��5t۵�l[̚�g�;�N%׆Y�ǝ�=���Dckj��J��V���U�����{�鷢+ɳ����"h;�J�i�٪S�/v���2붎��u�1�2�b%k�G'Nk�yY:Y�Wk���+5�e��;=Ӛz�,� $�l��
�m��|)d�o����K��@`t=1�6��ܦ��l�ڝ�Χ��I��Y`�Cr�k%�ɛ8:L�u��3ݗ�q��V�sU��)^)yY�IکZ^f��*���yV�St�v��/Qu�<%�.������dݛك:1X׈u _K���h)ۅ��+��atO�8T�kr}еV��b�"�{���S�sŧ�N���}E`��������5mQ����;�vn��V�>��b�Nг.��)���e��*ӶQY���vu�賢p�A��͛���xs�kLPwK�@��H���Y3��b�]
��^B��r�0u��#
n,���Z�l)핪��6�,T��r5��̓a"�+B���U���{�m�m�͖�o�-��6[o��+Sܵ!��a�%�봱g_�������$���Ϲã�����j��JG��*D/*�!oE�����1��۝��������ڤ9�фR��]
�ygM�y)Ĕ��4����E7�����Z�iτ
,s�Y�S/& A�����6�꥜;R��_A��"�2V�W����(@/'}���۰BV�:�C@����a�̗��G�:��-#��ԥԆ��XV�ܬ))V9e��stץ�}��P^:_����8�ݷ������/ef{7PZ��m��7��-�[��� �k`4��Ms������;�_.?�&�.��]+�� �YCn*X#�Sm���Heh�f��ˬ'jWH�]�;:�B�r6u���.D����R��7"Ͱ�ƴ�]��x�J�n���Df�#kB
��°	@��W]V"�J��0A�j��m2:m⪋�(�L��"��W{��q^e�ǁ�Y����*鷹�5�ST�SΫK���������Θ۳���Y��ңM���Z���h 4���c���w�49Z��c�N��6az�K�{�H:0MZ�9��y>8W�b$C@��Y��\�Gk8Khfj(��#_�L=��{�m�2�P5�+��t����ˍ����-hF���]�(�f��U�S2��Nv�Y��wo���ю$"2T�=Y�mb![t{�Z��Xbg��I���K:�S(a*аy(3+;6��]���'w�$ �b��y�u:�3 ���wYu�`��be�E���쓞�2����6�f�s�i�ڳm��1����
L4Jc8I��8�]�j\�x�wܯ�����4����Yx��юl�=Y�+r���]r3�[R�o-�:��ݺ�8�gq���w�A�fQٚ)��f�l�ȅѹ����m\�4{*�P}���)���؝XewecW�]7)�\�U�]�]������:�&*�ۊ}MAY�w6�4.)y7U����l�7ƛW��k0�2���d��N����2`�+$���[��r�"���gqV˖]G��W�%�]���)�YŗRų��]�E��⪗6�>��:�$Z�]ؾy`>݋{��W�@?>VWu�v�_a��w6s�?f�36k��aN���T-
_:��Z�$y��(TX
�y.S���tehw̃�7D���p��_mҳ�����R��M�+X�*W�H�'M��F�u�L��wur�qZwYq�����ܖ�Cwx��}H)}�WAR�nrrj��KWnwwuI\t\8Q�y��%t���Ib�{R-����"c��s��㣑�4�H���b��OfIm�[��a���Fڛrj��-�#�0EYaό��:;���%#��)����3B6o�o(Vm&�p6�٧���4DK{泗ni9;T�iq��lʋ���;��C7&g]bX���8�X���մ��[&��j��ҥw� L�1
�#V���vdA�L��=�v0`����i��N��>w|�<����һ\��)7^e�9V�[������tG)�X����VE�sH�ʊ�1�5Q���I���л����eb�nVQnB@��cZ�|��zy���(ڽ�]�Ŝ��*���],Er�Yi1a|_�3SB�����JM�Ε�3�d�N��w���v%t����M[Z_Y�y��R���:n�W
2������Y��B�f`��4���l����!Pui�X��F�{ƕ�>�;�"<� -~dPw/�@f"L�̺pm�/c�L�2f������5ޅ�EIY.GD�*P���"����:�J�������!���4+P�)����.ݒ���r$��$|��/v�Qa���\�_U��N�g%d��h&��Nly�;��{�&I/geX�@�7�� C�^��L�\����r�vfSu�E�7tKXkUrz����zr�Q�1I��eb���=�O��Μ7��E|hC8d�ĸr�|2E���^��7�ܥ��9��@Sk�M��=���ZUf�:5������FA{@nz��0ERQF��1&���Zڛ��m;�8�q&q\@i�V</h�-��
闵�@�;*�$�܀E�v�)Yߎ��T5���b}�V'������?�x�<�Yq,�G�uh_CN�{����xA�Y�l6%�2��a��%�8���J�n>B�S=\2��,d�q�n�՚T�ά-���4���q�o����]�aq�)Wf>�{������$�u�=���_-��lC�;._*�|*�^�q��I/K`�.�u�]��&��z����;��S���zky�z0�Agnp��^�8k��>vRZ��c�`�#8cݦ�:�+Q��i�H�ɖ�.��c�T+R� ì�=�Vd��zj�m��TJ�$A����+��et�k���6]�J��9�gY8�!�hܱ}/��+�K�O3��q�J��1q�c�k�����殠���a��__5����y�RɝԣN��j��n����h	�&�(�%Nۜ��ɱc{ְ.�
�칓"������RzV�e�h����1@�
�K,.y/	��9��n���jpe�(S"XH[V+K���h|��J¾[���{;T�,5x�'5�+��=Cx�A�7��ݹ�w�lRVa�N21Z�K�;�un�/��k��7�c1��D;��^�
�4�M뵌��@��F��Bp��Q֝w���������>��]�ʮ��WE�VeȀ�/������c:��_J��8�T�B��D��U%�:�-Kŋ�p	\�gQ�LZ���9-�)�&�@3^^^/ �>ě4^6�b�sj�!�HΥw�|rÃe�EJX";X���S�y%i�W�le�`Ѫo�=֦��PJ��t�lճ�����Vh��ʁ��Gy5�BCZ�0��+W����[+m�2���ʅ�R�h-] ��"�%bϬ�͹��Oz�E6�;R�m���G�W���b�o=�2�RA�9?��(�����i̻aB�d	O�wy��S�@��[u���A����B�O�`���li�- �i�������Xy�����B7�ѻ�C�d�`7|{��ԫ:!�4F!�!��J�*P=���ej���L�)Y.��HYhF�e�{Ҷq��J[G�ٸ���w�PPف��۝�8����MѺ҉Q��`inS��Z�7��	 �+��^��ޢ��礓7*�q� ��n΀F澤���+m��ص�N驪��<W ǂ�#3U:�Xu���%�\�{X{�gff�N��O���~g�`Y(��_lc�Z�״>�PR�J�Pr9�&`[��ln>5f��/���V1�t[��Y�F���'p����Aw�hud��z��0S�v�3"W>��g��U˽6I���V6V�|�f���M�Ӥ�&ĉ)a$\�������Aͫ��|� :<��`P�JQ��Б�o(�n�a�ƴ�87��ej*�2q��l�����]�4qW&1r�9��5�o)��v7h���p����Я����+EŶ�2�{����TQP	�\��-[7+�����K9�[�%eU��0]���f��j������c�2m]:�ƨ��j�5`̽��}S,n�xl{׆����Ƅ���::�%X��[�c��}Lѡmi������m.+l��`8���d�u�3^��p���kS8($����+C5�i*ПB5�"����/-:�*[K5L	/k1�%oH�c�Ŝ�������2�����>.�#]�`��|Fn��(oحH)���Gk �]��҆l�W��c�c=\�r�Ă��6D��K�N��_r��d�3���,�ʊЭ@�7���̔�=A�z� �v�z3-��3�yR��V�g\2�ޢ�h����,��fL: %��5+x��s�ZIT·ϖ�t�i�/��U�h��HT�v��LL���,��^��ƫKT�l���	����Ap #o���Q�Mv���y`��k���3����n���Ջ�#��s��=7XkoZ�	��b�5�\3}�jb\��q�mh�#i�Lm�]���e�2�ө�z�\��(�D-s���u�KO��r��p��6V�l��jJ��1�ı�qߺV7��E�/:���)��΀���r8� �e]"���Nb��ŬW3}u��,����W�nS���$F�d�Ꭰ�j��L�����̗2�6�j��*�4&��g5��	�%'ěZ�q��7F��D�P��Jʸ�Ye�wr��K�N�z��Wk�L��t>���6� �z��a��X*�ʹۅ�l9R� #ڶq�t��P$T.�+�/��J��ߥ�a�j�\X"V�r��*7���v��kE_n	ݷ+�ZN��]R��x:��pq@h�e@ ��J��<����hi��n���NWc�3O��64J_(�^N��y�6+����C2C�,��xn��a9��*͚;��x'NY1�\}���*�Z���,˺6_X�)�;�����jG�sJy�!x����ճfN�le���˵���{�m�ڸ6��Z�,V6�+�Iݣ��S��^��,�a��dD�Sڼ�T�\#+c��"�,[H�����[��	K�+��O4���G6.��jfwMM���V�	�C���͇��Y�\G�(��@VY8���B���z+��<B3���$4�g<Y�[���*�D�s�껫ǌ�t�g*<x;�)��Χn��=�-�;e(٤��O�<]oA�ei�yk⾊���JVsFX�.v5q!�΃�����DܹNK�J8��s��E#zM��������f�V$��o%�i�Kn��j�ڨKclu�f��)�˝�'aj����m�ڭ��R�";ٕ��k����{��gK������@��*5*J�:�[C��I-�#���I�H�XN��"�%���!x����&���66�x��;����J��*��j���_�/H�I/���KᕙS��'�+wd��t:�o��nǻl��O�R7�Wm�J3t;[X
f&��.�Z=�ڭe�I��*9׽���r��3���p�G}�l��܅�3Pm`:�z�I��(��ηf�mܛ�J����}9]H�̹�8#�i��[s�.���t6�b�-_]��y}��ש8�o:�A;�A;4B�,;4��>�{�*im.'x��c�]��?���B��r0��f_U�m�j7َgd�-�e7.b7(�QA��zp��oK���k.�6��㝲�,�X)*�L���U���j��L�zM�,I���V���Wؐ:B��:2^�Ks$ui�w�`���k��ޚ�x5��X��2�X��\�o5�嶵4f�Sp�ڙ*��ޭx61�8^���9l{��#�V�f��q	��& ̽����ɤ/�(l���\E�h�W�[�4uV��6ܮ�tI����%^�,�ƒ��H�G��nͥt^�yڀ���	�l���SH�VJ��}�ZE�QA�;->�b�p.���y�i�a�u�7b�YM�mg^�T�D���sW��f�Qߊ#�iWT�5e�6n�{��t�%i��B�i)��a�@圭���zglpB�vP�����)�
���9����E�ps�;��7|0�(���SM�\r��KnP�����fc7����^��i`�\)s�3u=�j��3�-�Q��kF�&�\�I�2��!Y͋�t%�$�<X��ev�z�n�������nWݮrU�����J���+n��ܾ� �.�����3.�uyrCa�4rG�f�6+�{�6'�p��M-��s�q)Pte#X��9 Zu����FwR\oFF�$g�%,
dBwQ�m�c5cc��}�UN�m��á����X4f�Cz+��w��V�L�V�ҧc=Z�-1�k�c��K_�H{^T�p�]iު���a���C�"{ՠ��$9%6�p{��+'.�f����:5v����KFX��!֋9�g���ӹԏG`�Z���f�hsl�F����*���j��%Dp=�!s[��P�r�<�Wq�����jr���+4���p]K�*<tm/U#t��՞f���
�Yg)Mǔ0n��_�ʐ���WT��X��o��c��t�d�M�#cǃ�XD�1}���Z�η!����Q�3���ý�N��=���9��<v�^�Y�差+μ�{��J����C�v���Xa]��ʨ�.�׽ø#�T�%K�X+n��Q��C����Nh�!�K���7u��r�6�n�R�玈S�eggX���B�ҁ��J�è�m��\'ʺ��l�x�x��������l���Sx:J��g'(�+���L$�,��6�sYԸ��U�Aj�Lr���+$�9}��:,|�{�{�ԌT� �d�K�U�ʁ\�Z��I�����7��jp����7�F8R��hevT�8*%3�*�v�ih�\�6]�f"�ɺ��c��V��/%�-I�>�FS�{csp;�]�HM��!�;)^t�1j���i쩬�l�Ku�B�q�-X�ZYX���]f�h��৛Y�oLWMV�	�R���)�&�R1�T��K,%Nx��|'����?
Q:�xd�!t�5�
�L�÷���n��
M��b�!YB扇U��)����Y��|��-�h�|@ٺO<��g�)Z�t�|��3��M����.P�4a}�+F��d��l����1lQm�f�W����O�w
C�ީb�:D�ݙX�mѼ��A͙*�)���;�t���b�F�5i�i���� ��<��ν�}-�mA�����Q�)6%M��'*���[���L�p'\n6�>�%n���9c�q�⭺�Y̝5ިBn&�$�(c�є�f��}`�J��J+:�X07շf��{]}� �TU�]��އ�K����l�t�����C5�;u��*!TN��O����ϻL�yY�t.�XY��3�y��t۩�K���U%�챩��("h��= ,�o��n�V�`���P�BsP�=RCt5c����(|j<�w�I�3�S\�lU�J�M5ީWw�=��B���k�k֨EbB�fغۆ��4>4'������H�Q,ܪ�"��`q�{XaW���E@��塆��M��K�/PR���Bvǥ^e��t���`g
�8k4�����;8�-��@cj�t�����ɶ'rb�ZLT)��(�Bг[�}n�'�_h�h��ʔ4��i�hP��s�x�כNF�{�K*\})��p�Y�C{�8��K���qP�Xm��pv6��\�駨��T]�Tܝ�@�!Uql�%��)g2Z��Ϯ���8��%�Fq˒��W�Qf��b��Η��;�C\��i�iz��Ñ	&л��e5j�h�q�7��>|FA}ʑ9��%�کC���M�4_ϚN�,u��!
�]*]1�:�p��룄ǽ���Ô�|uB)]�4�&�VC�����3hx�n��mwe��͸ӕ��Y�T ��Yץ�����rwR�C����&��]��}P�x�u�'gmGt��ԗn�괖�P�!&A>�[Q�LT����.�c�q����Q�Y.P�u��S��j�(Q�KicD�j-��PET)��%��iQ&e"�YV�T�`���b�QV�֨�4���b��J�U0��A�]f`�Q(�+J&d���������ڴ��m�.86�e�S*a�k�#���2�QDbն�T��j�%��F�JkY�P�Uĸ�us�j�Jʩ�˖S(�aciVブV��fe��r⹫�-���T���㙚*����naF�e�iauLc[R�,f�2�6����R��Q�N%�X\\j�)�U�5h�+�r��-��L1F����T�M7��(��D��-U�?C�U�HV�:��̫4�D�<�.3]��GS�V�6ep�X�#'S���Z�	�֚ê!	�j�C�R+�΋��\'G6+��AU�T;�R�B^�Ӌݖ��+}�{�f]9og'�NT.c/�z��j�"�w7MT
�>�� Zf��Q�t���ʷ{��1�w�x�-V�v�w�bV��M77.�L��İv���0. �<�LQb��e�ʣ�Eq�B��xp�݂��)4���T�ﵟn��ķt�z��o�b8�}+�;K{�L���Ŭ��������V��b�pu�P/��e��v�������z?j�V]��E��ӱb_�	Q������.�	�`F�T���(�AN��
]cx���;%���v:�I�h�Ny�0�/��̽�#�����:�K�>�=�f�՛ca����������4������:���G:��/�����d�=I]1=5�yrċƅ��*�C��{לm�2/i�{�=�z�vYε�H�Vu�f�|���)�.�"��
I��1^XDͯ��_{(>���QAp謮���I�[G��r�2����Y���#����O�N�\cْ�^��r��t���e(z����ʧ}�vQ�&��|�d0t˛ܱ-@s}ݺ65���TʅV.����~�T�Ԩ��	͋x�W_>�_�=�Z�9ѣ��ܕ]���e9�ʱ=4���V$d�jX�ɡ:�L��^�I}�6�5���Xe.�I4˧�J�n}.f׾%nJF�	��Z�Gޫ�8Z�_�N�GEؽ���r�+�헜�>��pҕ��2�t[S|��+��Qj�ڷ�l/BՓ�οAϭ�b���><wؼ�%k.orM���i�M�<LL���\��s8)�GXP�œ��f�[���Ɗ�M�yӼ��9f����hc�?l,g	��w��0^Xn(<ϟ�#�-�V�3��}hi�[����"��������c{�������<o�^��h�f�|��f}O2Ɨޞ9"V��t�giH{/VT��ȩ��ع��v�5�F��b�y�3>�%��X�4��8fn�u��ny;�z���R�pv�*3�[XIf���=]�ы|tT���|�S��nmյ	�{K��CX}FV���׉o�X-��Y@n�U��$�&��V_H�nv�Ûܵ�#+�@��o���v���(V��4�K�����A���Λ:����X'���T�R��)�'6���<����iVە����8���{r򮝌f]+050��;9$:C�h�	�:�;0 kP?>K1jN��朶'L	�N����\v1����	����})|a�gwg{ܛaR�������Υ�>�
Qp~�>��jp��v���HT���(�Ԝ�B�ц�m��&��B*�ᖙ�s���a�5���IW��Q�p�W6Κ���>��={��i?{\]J_xR���ٱ)y��.2�b����w�Nysz~�!U=�,�Ҳb���:�	�Fi���\䡗���o�.S�o���2e�ށW�R��Em��0��;&Y���~�:|+x�h�T��ÞNé��ĔH��'�Ef��rwɱ"N厢�[Tb�6�^u.�Nz�j~�h��<Z��{�]~��ڕ�=��	�}��o��ܣ�QW�	�#�,��g}���_Z�rݾx��ńҬٖ�$:voi1B��]�٣{uLh;N���0r���A���+���*����B���ڳ��˛�Bs鴦�by܉��)#sqM���sX�j�p��sq.��s���X��|�:ڂ?%����Ǹ�l//̻u�%OR�]����ۃxwem^ֿZu�`S�A6q��4ȩ[���s�nd�yqՊ������k�B�I��r�@�Hϡ�N®�8%=2�EN�^�L�SB���'Vv���O7V�����jS2!	[�8\�k��R�6��Pb�j��Q�W:$V)��U�r&7�TS�A�ps4�>��3�K"���ѓK/ؽh[��m�	N+iEԷ�O���K�3�����r=�70��z&[��y<�Q��Gz���Ã![Y��K��<5ɣ�5ɚ��=�ߢ ��1��U�5��!G}�G���xȷQ��D�L�vk6)�)�m�O�'��=\A�[�v�@oR��hn�]��=.C^��h��	���yOOC�Ś�m��
�J*2��lv]o�d^�/{�$�dfƐ��Q��j;x��	�h�f�-
X.4��z��ΆG �-�9YN�J-k�gR�ZOu��^E$�9`�U�V%�8v�NՅ���Jו��W�鯸�Y�k圳��ך�6��9%bݓA�;i�o����i.<��=�ה�&EF���t�i��Y|�F����޽�I��z��7v��aE�
�:�M϶]p�#�E1�I��Hȴ��M:r���W�^-��u���,�w���eN�t�)\ͯ�Y-�]Sכ�f��Cܱ���9���{�&����Zt]GNeN�U�������hKLu�qBYʘR��viv(�ʹ�6��m�P/,�:a
��|�C�R´���m<=����'+���e7P4��ւ$Ƥ�&D�gm>KM��/�/*����b]�Z�:�%Y2���H��:nB����U�����Ԯ��Jʯ�¸��s�m�:ۢ�������r}K6٩U��.�Qw{��Yj򵜃q��/��{����	U.ܝ�u��5fa	txV#�V�f�g���zx�W#��;��dV���\f��>��hz�7;��hR�.��j
�N_SP��/�.�`AC�^�R��"��C;u����V���8.��E��P}�iR9.�T��f^�+��d�OgC�U\���i��+J����e�n�p�HMm�oq��nw�$�O�-��V�:Ԣ��ǈ�Y�{��V>uX���>�ne#�CUx�+nr�:�t3e���s6��M�����VbCC5��7�2�Uk���l��+�fU;��y�͖(��S�;UM�r{���ڳi]�U�ɷ��ʨ�B��\�78��� ��su���{B�K=^EJ~�?{�-E�-Yn�{�:��93Hm40��ԍIĈ�ä�\��KQK�/�E�'�5�t���1J�������!�I��H�����;�eb������^�t6��;�]��3$v�Ƞ�-��;(9u��E1��U����Q��M)G_e��N�^s��q����P�ң��iR/��@�s�hZ���{Vr�Z`Y\���zf���u���4=�}d~N��3g�2�9�u�y�G���|&�g��0���;�5|=�p���ˏ@����Ն���λ8E�I�&��C�2��	x��m�$p���{ǩ�L�ঃK��չ�2w]�N�	��e�{y�G:�|D�zJk���gm�����	u�dv�<�2��tՎ��� � ��:��C�����o[
뙩���|γ����ΜRŽ�sA��\+��ˑ�K�^�3��ʚF�e��&=k��.V*����߰<��.�|i��0��'#�y�q�YΔ;f�y����"�le�VPkq�Cm�Τ�[#v*X��I���Y��%�-�S�)�
S3J���@]q�����SB�NTU8�����Bڢ�;ઃ�y�9�I���0!��
�?�6�VB��]�6E��Vt�g'u��`�!2cژU❚h�3 B���'C�#g�f�J2���b6�É�s�-�ܔ;K�b�'��VN�q�ǫ�2T�^ɾ��ͩ�L���񜓢��u�M����.P�2��#��a�$4ץ���ۻ�Wy�8K�/V�7/Ahf��;�뷔&�
Ƅ��2��fs��_���v��mz�)�*p��̈́�2�i�NL����oK�NE�fz�⤞�u9�*��"�[���>U�;2W��W���*祧��N��o6��S�� �f�o,�� ݴ�Nħ��3O5���	�����Wo�jB͆���FV{{k��u�gɾ�;<��׉�v]���u)���.]}�%��MF
�ʥzs��+|�Uӏo�mg��MS+k�%�Ҵ�F���z��]&��g!*ox�*Ҷ�i�'a�v��J'��uWEϬ"竲$2�z�H���dU�/��y����ET�&/���D�*OE:�.�,�o��t�4��Ž�^�"����X��3z0>��Ǟ̓�F��x�qT+���"��!��6VU yMm55�Zc�@f�N��ӆN-v��w�����)��M�1��9镚l���n�}~B/��B������[�����:�	��lC�hik�N�P*��d ��~乜9��'�8��6^1�+j^�9۵�XN�ϥ3�v�� ђﳻt;W���qɗ�>�R.K�E�'y��;�Х-wt�-�ś�XT�y���+_�P��f�y�����1�\����V
r���q&�(���u���@z����\�ݸ�t�Ц���k�����a��������jtn�J6Ŀ71��\�����}+�D^�>ṥ%&����s������mI��dǄ�	�p���&Cw�a󗼸���Ìh:����b˂�{��U�O���O!G���w�n�d�
<{C���8r�c�OF�VXv�ۊ��zZ�����3y+g�Gڬ/=�O�K]���C폆��N��:{�1�+���#9fsg%�sk.�o.]��<2�����>�W�ޞ��8Y�6ޙ�j��tfj|@`���ܴ�]D�����[�=��ek��z1�G��Hx�L�^ɬ�i��8���*��Mо~����:pTv��E&z�F);wɺR��5�elG�\��v����M�9O*v+��=��dZ=�Vt�)x�Pt�ܲW���ឝǗ�r�n'=i~���!�H=�U�WOnJ�y�yg�����M�y:��9������oz�Su	���)n�]#�+F{� O�"S�z����s>;\�z��[��ͤ�n��g�򹡌:�R}�8�,�B�����'W*ܮm!v`����#u�F]�C6�0�k{��)���3���x#$>���/����u;"�׵+��j����V�Sq�����k��]O��������fK�nŽ,�y�Έ{%��%rO�&:�܄߫1���g^�3z�٘�&�׸��q�>4��G݂$mm��M���d�k|�5�WYNs��m��8�OGM�J�J[ݺ�j�5���.��u�(mմn��Pw��3	������c��dɘ���Ĵn�̇,T�Zm�zy��g�[Iz�w0�_WB׽Y;��&�J�$ �jaW�vi�pd�����l��;�ҎM�H�׸<��׾��o2��@�u5��uR��	Y�t)J^��ˤ�z�K���i��{��.�Ks�_�Ǜ~kv�jc\��<�����(��^��ۤ�Èw w�J���@M>nP1�q�I���y�S���ӎ�/�m������ts~�� ����:_{\͈�VoCKV����&v�)����~����[>⟽ZU{`@��Lw�{��-m�a����ia�T$܂�V�k��m�����=��F���ۨko��w4�X�Y�6��\y<����߼�/%�sh"��$,��9V�;ݣ,*_r՘�ϰ�ZE�w}F�hb;M�ry�A�)�R��U��|'���$o2�,<B��J޻� P���BPt�q�/��Z���;���ʴ����jF�v;2����%BZV�p�]�X��:�=L�%0H;:.��u��c	���(U����ª礪�����Rqh�V�	�9�G�E�z�_l�d��;!6e��T�61���5@���&�n�:�gW&k7����q���Й"1)X�X��3b���w���zAU�W�c0�R��.}-���_i�5$�3��V�4y����Ĩᤅ!W�xu�ҥ��T�� �$淕�B�c��WDE���)��&f�ڲu�׸� -�y�*������u����vU��[�ʋ((M�F�%�f��\�'/]^h���r�'4f�/��U �YŚyd�e	#��!--b����B-zBr[�˹ۛ��TDǽ���}R�(�<ZH�ھ���R�s+8D뻚E\�ђ6��Zl
�Źњ)9r����L���wW%H;Kl%�(�c� F�yњN`|i�!��ta��4�{f��,d��S&�����!o{jj�K.�v��2G�Fu\��0��I�W9�y�q�o�"�d ֒l��;7k9S���EQ����7�|r�;��'zAz%sF�rՋ7��a*�fJe�4m�E�(�G��h�I���
FՊ�nȻ��Ō@e�$�DɕwI�]չu0PF� �� ˬol�$K�>YIr��vY�*10� ��ѥ,K�N1�19n��h�	��ԸH6�aB(-�n�Y���/b��g�HD]/�1��uu);�%#F6Dd!�1t�՗�a�I�����n���\���aY���������3j�Q�b�:�b� T�+���*���U�5�y��&r��b��Z?����;��pT%ڂ�n�+0eF	ߦ+��@�b�H��Z/k�7�@&l���z]�7K��m��t3
Z	 ,hY�t[n�(e�W�n9xqZ	o0�n�#;4#���bA�K�%��:��w��s����j�JV��_�]����,\FÊ�m�|:�n����kjT<if(��F^�
�;���p(͢��V}f�o\�o��v嬩�;B���e�	wa4T�}n��SH5r�M��v�(/i�ف��7v@��c��ъ��3��Z����k�mr���[�N���W�*"��i!�����UYr�]ڢY�Q̆k��9[��a���Pǅ�k�r��(�9
y�¶8�\�Q:+-_4Z.�!/�fh[٪ry�}���Ԍ]t�����_�mݵO�KR�m��w{l� Q�@��m�6�T���V�0RۍlJԬ��1���,PJ�DEJ�m-�IJ�r�-+J[�LeZ҉h�������-r��UF�Z�S)���\a�q��ƱƢ����)p��ƭi\�A¹nU��\Ƣ����n&*+is3%��R��-�LŪcXb��ڍ-*����T��m)JV�mDKF�c��Ե
�Z�[TT����R�[mkj�hQ�EڋX�-��-leE*�j�e��km�+U(S-�h�ڕ(�iT�ij���ˎQ-B����)YJ����)VT��X�QX"[VT�*+�5��c
J�jƶ�jR�K[+�L�F�R��EZ�DH�Z²��5�ѣ(�����,Qk���몼�U�ݠ����n��d}Y�1i)�TЀ�5v5{�x��wg�8��50H��Q�Yƭ�z�u����/�o��u�&2�̈́u�e���A���Z�%�/���qhN�<,6;��=kޕ��?{��6z��~�s{ⵙl$�?��L�i����+����oږOV�2ZsФ���%�{��>�M����o��=-ćI��#t�|�*�>e�_:P�.�u<�{�fq�4`��q���{e���z4W�u�/k�`�q��N�w�5���Ad�9���]��mbKt��%V���hi�9}�+���[Mߧ�J�8�F]k�璋������8�f��l�|�2}&�F�l^J�`�8��u�1�[�a��s������΍�礦�5X/��@�)��!)�����J���[��j,m��*�������զc�TS�M<�^�ɔ!��X�i�-�ښ���7r��s�
�Kz-2e0��f���m��	�)9W�z_�ϽܵFb����S8�(	��K�˄;��v1	;3�]X\ٷ�<�,9��G��x��^�:�0�k�FŲ01�u���Di�n��;y��sUm5$�v]�n�{��Nv�96�];M`{+h�ٛWwԢ���������:�lH+k}I�|�� �k���k"�H�lW_�4vwY>�~��E{R��ݝ�e��Ev���j��|���G�:�T۝����a�#��J�?&~������EA�Y��k$Q�Ir����ScN��y8��7�L�
��|���y�5%�!_{��iN�x�X�=9�[/��C3��Z�T�߹����~��92�K�����mu���%FM�����`��Č�%�NC��vH�egV�kO��x�z*�{�'�h����ɧ<W��Pī�l���+z5y-����w����Ҹp�h#��л��EG��xOS�vf�L�\���n��c'D�U4ڨ\Y�2_�42��x�9��2R;l�U7��\O,ɥ�r�N���1�ɖ�l���}hi�R�B�ٗ�Oeq��uˡL�c>de��?%Yj?+��@$OvҬ�Y�Y���2`���W}W�]$r��m���'����;l�e(�QS�:��w���p�ʖ��ros��rW1��(�WAg��\b�[	b��I�w���0�qк��I���Js�\�!WK�e��Ł��>�<;�kw@����*Q�0��ә.�����n,�nH�t�,0c�1�������):䬤N� ����,�U���/U�8�J�Yaʡ|e�vcy�я+-����iuy)�.z�q�P:'���ʔ�Em��\�z!H�����]Jz��W�Bg8E�Y`4n�Z����W��������c��M���r��ڥ!�����7A'���ɾh��7-�~����EMî�뒎���x��Ym��S�ڪV;�Kv��9�e9W�0����v��~���s	��Dc�+{��^6(f�h*�^�i��Y^yۺ,���¼�(JT�k�k�:L�����4ƚhrex��KGN�ɥL���ۦ3���}`���szx�bu��~gh���C�<`h�x)'�5��N[$��l��Hm�ĝ<O��}��������u'N��맺�%�J͊4j�Ǻ5�뉪n���O]��$�ܺO
���Gmq{iK��!�}��3w��^]�}fJy�����WpvE���5��k���	��k��o��׼�Z����$ ���q�y�A[��j�v�\�n~�|��">>��'s|փhm�2r��CS�`��I�u=�'�!��Xq���"¤>I�'�\֤� tf�5$������Ut�R3��Ơ�-;5����>������Lvξ�CiϹ���N$�s0Y�&3i߹����h��,�	�:9�O�Bh�2m'�<E�y@��zb���F`��^|������Α'�٫'�:x����6��|�w`,��S�z��4���6��1�:�Z���'[�VI�9�,��������w� �Ϸ��*�}�g���̀ x��$/�N0�M�Y=C�z���d���3��t;aXL:��2v� vu���:d�Y�P�IPߞy��r�͇���~*;.��	� }�|'�t@���h2yl�M�;I�����`h�܇I�!������Yf�OXq�r�>>���g��� 
�֝�+����ma}�,�]y��{���O���N$�4g���d�a�݊OZ�k.�=a��&$�'h}��m�����Cl:<�;x��:5x�<aSz����t�c�낗v�[���|=D|�
>�O����N$�&"΍oq��f�ud�a���Xv��s��$������C�c5:�m���0+=d�I�[�믲���]����N�g� �4��F����A93܇�q:�xq��,�o�vɖ��o$8�Xj�XN2t_�,:OM��:gl�����΍���X��u�V�-Eb��ح�����!�:ö2v�$����]}I�L��!�d�N��z2yhM���2���
�Y9��'9~�a���2�Փ�S�X���v�7�=�9�XN�k�0�!�'���q'��'��I�^�ԑI�ϼ�s�$�:7��z�C�����4�\� VU�_i�߿(Эջ�e#w�?J�.���Lr�!$���{���ٹ�J��Fv7XI��X���y�CԂ8 �y����.ů�A*�g�"(����k�=8+��������N��[��X��1���@Dw�;�|�8�B��qZ���0NҠE9nrՎ�EܗonjYW�}�� zO��_	g�@�9��vɯ;��I����q�Bu��06�'^y�x��8���&O��o��z����||4��r�¶-�}q�}|���u�^�x��'�����B�����+�������t�5Bx��4u�$�0�w��j�5��q�h�x�ԛ|��xzϽ���/���AЛ��������Op���x���~���=f�vs�'��CΧ>�Rv�9��|��:C�VC�4���$�'��l�G�7�<Ͻ�G�|幻�g7������oa�{�Ǵ�8��>�^�G�|eg��N�����'i�!�s�jC�=f�w�y�=a>N���!��d>C�O�����y:�$�&s��k^SN��ًj��������q�����iQGt��m�i��}����z���'vo2!�=d;�3�'��s�m�z�e�'��!̳�4��,7��}��b��]��|���Y����>�H'�Ȁѝ{�>�I����;Hh��I����y!ć�{־fМd�Z!�<d�6�i'�V�s$�3Y������*����f�^��Q$}�G���E�@��M}�$�����3g�>@�8��yCl��>N��Y'|��0;a�O����Y1�|�s~s��%��1V���)e���D>_H$�{�{�'Ȳ>̜I�'���-h2k���M�:�a:~I6���$��i����;g�������c�c�ͱY0��f����/�H� Q |/U{�vɌ��8�d����$��&��È$�;-h0�:�d&��{����w5d�������a�����*�s3u���I�}� a�2N����'��}o!ĝ2b,�[��T4s�(��I����I5ֳh���N�Y6��'OR�!6��o�u��c�7��Ɵ�f�en�Z��V��X|�Խة�����od:�����s���ۧY�� ɭ��o�w�L<G�:DW�V���͌1<���[��"������mWB���b?<��Ը�«NnQ d�.�8��a���E!<���#�d>�0�zȜ�}�P���8�Mo��:d�R��C�<d�YѾ���Pѻ�M��7�}�����\�| �#ٔ�	��=��{�u�}׼��N�c8r��!�{�Y�N�|�s�gM{x�=B�F}��Y&ޮ�d�\�C�<d�a��8�P�f�:��d���ѻ�//]�������%t�n�0H�:G��xL�>F�֬8�|�3P��	�CGt�t��vyH(c'[�a+%L���8�$��t��d5��T�cP������3���Hbau��+	����M>�8�e����N�Xm$���\ԝ�l�L+'Ğ�d�&�6�G�$Rq3�> �I�cｽ����Z�����2n�y�@�n�{��Y+'��v���yx�P�J�����&�'�w�N!�'�S�dڠtyd�_�~����e����1D3����G��]�������܆���C�y�[!���C�������*�߸(J��O�N�q=5d=a�'}��I�ʟy�H��A�ܸy*��pui����^��םw����RN�vɻNO�'�M��7Մ���ĝ�!>߸z���i�;�2OYCǣ�`�+7���� Y�T� Q��	u��v�b�sZ������Or��RNN�=d�:<���jto�	��y���	�}Ci:|Bs�~ԇ�z�&ά�2N�}�}�>G�[���6�36���nZ���;d�3����&���d�����E����ɶM�]����<v��������0�a�)��g�G�}^��Q�'8�'���o�(��]�,�z��z2�x���`q�L�+̤>I�'\��|��[�9l��2M�n�����t�Oa�d��gC�|���0��>������?g.�"�{n��Z	�
�u+a�� ��{L5���$9�x���J��&�;��ص�j����}�}���6�j�<z��5���p���@o�8��|F�l̛y�Iw��ZĹ��n
�E�f�lub��}� ���]���KG{g���I�{�Bm�0��>�B�2M�yE��P�fM����IX!�γ��� u�'��m�$�N��;a��G�F��?qs?gvu_� �xq���Bm&퓌;I�q���OP�<�|�qe�OQB{l�OY;�M���u�ē��'�&�ü�����]�|�f�g�2 ���|6<ϼO�#'��	�o<x��@�9̓l:d�m�МIXw�(�M�p��R|�x��'v��h@��OW��|��]�O�?<Z�j�w6>�>�=�I���>�'�ힰ5�m�ĝ����y�Iכ���4���M��&+5�`N!Y5<�
,&�w�,��	��O��v��0�|��Z�*���>�{�=��#�O�H�a>`y:���&��v�Rt�uM����u3y��I�sL����[�q'���u5�	�����;�|��j�����������^�����]x$����m�����H|�k�`Wēhk�aĚg��I�0�rg���\xI�	�:x����Gs��s�|�W�B��&Z<� T2g�:�M����Xv�a9l�W�OXm��Lf��m!��8ɦm']�
bC���0�%L����Z�u��.��^s��k[����I���C�;E!׿d��e���� T5���q���L}a6����2tY�C�{}�>g��쁤
>��������R�w��=u�~w�4�;�J���"�t��7��-����+'l�l5�o@T�C[�%a8ɫ�
��&Ӽ��4�_�'��i��g_,��jv�~G���w�$�4�x�!��"��(��'��	�f}�:�M3��!�Om�����<tð���T��;J�c�����	�����^���Z����U�����>�NGv�N�i�uې��Bh��7V�xs�;�c�Hޖ��} �J�̑gq>�]��;�m�7��`�:~�vG�ܦ�P�X�t՟�E��}�Tn\[���F\[	��W��-��a����[ܻ�Av,٘/�\]^r����ʽ�������xa|��O��C;�I�8�x�RqO�tRm���}a;@�h��{I4�q�I�!π�=����=�>�9Ӹڨ�_��5�qw�
���>�g�}�>��x�<�ܜa>I�;�I�RN���@��P6ɻN��Bv������~#�G�>R#�x���▿�5����>r�{+>G�#�>j�{�� ����d�$:�!�'�t��d<a�MoI�Ms$�,'�yd�'-��OO���8�@;�xq����������Q�}��:��z�xß{�����C׌�hw�'�;�a�	�:>�'L�!�5���<E�yH|��N�E$�'��䜷��66=�}��*v�Ⱥ���Õ���_go�Q�G��>� y��>����C����'���9��	��5E2OS���x�t}�8��O`Ɂ����z�����sc�u��7鈭���ՙ?3{�~Q�i���'d��N�3Ö�q0�0��!6����<d�q;=�	�
�سl'���d�'�ͤ�N�a�{�s���o��g&8��%����� ��� �=�q |'܇O�&ӳVORt���$6��;�� ,��S�|��4���d�C�LC�a�d'�*<�EY&��:��*�k"6˶��Kb��s�O�D���@<d��w%�|��&�_kP�H_l4�a6���䝳�S,�!�;g��}��<aXN�{��L�G\�6�L��������Y4���G�����QI>C�h�{i&sY�Y>�N�'$�o�I���O���'�0:2Ͱ���]��d�|�>�����~��������>�>� ��������:5���G9��$��{Ȥ��'Yv��N�<5I��:z���d4u�g���tyHv�2t���a ~x���-:g�]��2t��F¿��
(T���}x�;����������-N�g�)�B���כ�d�&��_w����K޷�븭��[��];�ĕ�7%sZ�r��R�bS����ﷻ5C�6 m^0*9����p�Z/{G��כϓɬ���&�T���C��	�wy�L�"��n��;I��F��8�Xh����>a�8`�����+�'�T�H|�>�����oIe�X��v���,����ˮ����=I��c'P��I=aSY�C��6�]�q��X�@�-sy!�J�Y�XN2?X��4�y�>�}�ތ�]�['�J���B�vɌ�0�!�����q'�+h��I�L��!�d�N��8�ݡ:9�jb��htn���~s���>�F������_}�e������9��v�:5a���_a:C�N��v��8�$��'��I�_�N�m0>�!ά�L�{ÌZ�u9��"��.;
��1n��r����@�
Ú�8�&04y�
3�'̰�3�O;����w�������M2mN�(��N"��	�G��ǽ�>���,�hS���9��S���_y�!�_����=`z��Hw9�jd�<z���M��'l靆�OL�`q$퇙dڲL�'6A>��" g�� :�3T�Z\1����ּ�o^|��!;d���P�'�>��������X��4Ü�x�T;��ڊN�c\��>d�!٫!�d׭�'�����̂G��ո����F��n�u9�? π����� q���Y!�����ē�;�2a�z�vs��C�=f�vo����������R��i��x�sV̚Ioo��w拚���?e.���vf���{�G�������l�$�0�Ĝd�6���Hm��to޵=x��Oa�3�C��gOd�}`�����,Y>gik�o=�>�^��{���b�b��G���A>G�#�D״XOP9��}l���'v�!�`m&�'ǜ��8�sY�6��'s鐈�>��Q�* {ȁ�/\��<�7��ooR�'��C.�PN~3f�~o"�txc��[O;��\RU�:X�ǖi}Z���8�{�|�ʔsҡ�V�1oi����$[������E�T7�1Z����9�*ފQқ9�}j�@���KE�%$.�l^��z�_җ�ݧ��;.��i'���� z�M�O�|��,;2��:�d��O�I���gFy�|ô���6�l�:�xAd8��y�]|���|^���2���t�%X�������.�M0�&3���m
�;�
,�hs�Y8�!��i=d��>��񁮾֡6��g0�?$�N�d��I�������".�ʞ֍]U���w��ڳ{�����q'hi��rO����Bq���(��6�_Qd��M�Xq�5'a��m�N����o�z��|@������oӗ�juүs���<`p3��I;g���L�$�{�I٤���N�1u��Rd�u�(��I�[�d��MN��@��>3�3�U;������~fc���B��?B|���2Vx��O,�!�=d�;��$�
���I�s!�N�!���I�&"ε�!ĕ&�yY&�u��O���֭ʬ��nX3Z�|��֮��T�'&��`v�3S�y��d6���M0��`,8ɤ��$�
�=��"�4�nÌ����7��O2�X�#�� ����"�,J����"��#���'!�@��$�Y�=aSĚՇ����l���t�`t��vyH(c'F�J�Sw��Y&Ӣ���dG�#s���Y�
�,�յW��^��P6��;�x�Xjg�h�'����'ܰ=C�x��Ն�J�rɦm��k�;a�'Ğ���A�>������<���\V��n���|8Oך��Yw?q9@���G^E��r�e�.��.��ǐ�V-���f��2��ǏKWw9��ܭ��ӻ6|��ϥu����y��ݻ��K.�e2��V	Օg��kCo�6�lɱ2K
��)�������c@���e+��3�vm�q �(O2M��۱����GT���Q��J+3h%L���g"SlZP&jA~6&����M�mU���T�9٢ģ����5ݩK�;{�*�U΢Wxr���1'r��]Ǳ�`���VLY�1MϦ�H��߲U ���rc�\VZ��QK�J ���9#��Y�k�_	�&�5�R��[�0���Ω�3-��P�l��(�ڀm���q�{�Xv�]fak�Qw��1ӥ��w��*1w]�%wDv�r��n�1�O���HNt=H�>�t�{Q�w{WrX��K��l����[���]�W�����[Պ�|&�#�`��5��'�d�������)�w ]Ӥ����v��ٗ\z��eU�RͻQČbab�	̼�g�p�s��WR�F����^,���� ♇8�/N��u�.�{gP�חMRgG*�]r�l��`��@!�ۣ�B���$��A��;��:���J�UH'D�v�S���g����]bMa�q���7���7T�b1:ۼ�uk��g�Cɏ�D�͙-o��t��何݃��W���:,K�N����СSIF��&r���Ǧvwm��Kr%��N�
�x֫d\[#L룍�#�K=�1q=	Z�ۓ(����
u��}	����cujY4�캽�7��_,m��UwY�y4!Y��y���e�R��݉;d�z'tǋ�O�lCn�-���t]*ԷM.�6��8�۰�fXhUKxtZr�e
#��͵,n�0f�,X��2����?`�*�@c�x?]�`��*謖d8h�V(C'R�H� �jZ�([ |���Ae�	���f�n�+-��T�h�ƦY��0�7+l��:Ie,0� �b̔�g2�E+4սH^��Ax�F����,E(�U=�1����n]A���tR�?*�K�	�,݂��1��$>R�%GX��n,�l�����vfPa�l��F����ϒ�GR?]jR���F�B��[�^���:��˫Ǖ.Ѵ	K���1��o�#�w��ߧ�U�uk͵����ĵ��FZM����so&�-4�7�ff�Y,qu!`�ѥ�Mhɴ,�t�;���q����i��Kb�RR:����z���p#���ÚQ�u$UOt�q�ri]�Z�庴v��E��h�[�[t���KW7�w���DR,:� �a��(����W�[��	N�
7���ɔ����{�J�8�L������c<�bce�Z��4�v�.`+�c���o�O74V<�&í<�q ��b�xʤF���:\6/
C�T�1c�+D{��T(�����'��J�t��o������:�]�����r��}�4����\]5#���"K^}��x�;��F+iW�3
�Q���
�
E-����ij��Z�b�*	ZZ�U�,V�D[lDV6��J�+FX���6��)�Ⲉ���Z����V,bK*����Qkb�,kq��"#�mH�ڍKb�R�m�$jڈ���D��r��j�#U�U,h�����[lDkA�,�E�-�
���5*-(��%�j%�b�"�T� �DQX"����j
�c`���QUDTB�
�$Db�m��U����*
��ڭ+e`�T`��-*�����5��((VV\�EJ�J��cTQX�����V
(��QaTUE��,)�dQ��
�����*QU�U�TQ���JVB��*�1�X���D��\q�X%��T
[R�k+(�
�iEDb-�X�%����"(,���ւc((�ԋE�cJ��Z#�-��������5�fG���-u�铛��QzU��9OJ9��MM��pŔ۠N�W,+0�7�ƨ��V��b=��{� FkkSb���p�������S�ث�kͰ��ec�oAW�����E�gut��Ke�(rR��z�}��<����^�����Kr�a�B>�|�����Џ��>�� w۴%1�Tt��i?)g#��s��F�<Z���f&��K�9���#�A�:�=6��_u�	�ν�w��mtmNi��K�wӋ}~��g&TLҭE���
����b�eh��"�����[��խ�޶�r��x�u�9Þ���
v�+���h̷A�r�	M�b�͵�H��[7�]��>������c��~X-����h,5X6��Ūu���Qջ	�߹c�1�ɵm����;�nWA��θ3��S����Fc��둪p�<�v־�N�j�g�r�ȉ��A�;����+o�ԫѥT�u"�
gdc�1��U�W��~��K3���ͩ#�*X�_%[��s=�P�{:����<�-&��s2��C��;�MHn���z���N�T��<�{��v��������Ik��[�\����5i񥖣)�l	��X뛝�;�cfٚ`�N�Ԇ_/�_}�UW׈Lu��Q�nb��%���rfMb�Uz�4���pXnr�Vf���,oP`>7�pX]x�Wy	�V�.��Z)���ju�_^+ޠ�S����<E�@'�*�af�o^>O���sl�4�;׷P��cG��<2Y�a�1U���}����/���w��.�H������B���=O;UM,y�fT�+�=s�w�v�O�j�-�_�L�X�%�.P7����I׹���q�ݸY�g���[%��$�wYu^�P�lf��]u���poF���9�Z��K�	���f�wC����x�c�����>�6}I���&�m��KR[ٖ�����NC��c��l.mŏH{ vԂo��Yt�Rjv�����m�~¦lV0!aT3��%N�0���vnB��-��G�n��YV�Ѩ�t�����w��r&�b�4�����zv��t��ǳ���@�w�ms�v��u�*�61�
�;&�y�U����׫��;4���m�o>�i4���N�眉�=D-�9T<�������S��1����ptOv
5/������$�y^�U��Cɨ��&&UͭkWQT��Y��@��[���)�k��p�o��YO:K5~[Boa����N����s�~�;��u�g�噻M�'&W�=�g�hJW�����s�<\�,�����?WM��4�N�}ٹZ��F�ls�)�Tm�4!t]{y�~�-vE�.�f�٠;��b(���O4���A��*S2!	U��r}+�ۼ.�j�_l7���d����#��=L�x�I8�41K'��½p񫙷�����Ӗ���m��/tV�s����Q��bp�a���2P�}�E"
��n�3X���Ç\�crX�+}�m'�+`�y����aY,^i2:�ϸ^#.��X[�y(P�lUT=M�J��ynd%;}Ŧ�z�+ӛ3~h���	ۨ��o.�^44�e�&�f�â��L�]���_Q!�)��U�Dڣ�����2Z'r�YIm9W7d��%����7$UH�������u��td�N�FW������ol�#���:�Ձ�y�wz��V���AYy#T�2P0�
��f����x��IZg�;oh�����bp�\�{�+.��KH�[�������*%'^�]oT3��g�{ٜo;��t���j��ջ6 W�ؒ�� 3˺��Tq�^��\�f�ڰ��yN7i�]��Ht:ړ�G�9>�����M{<�J���.ե.��i�����묻p�ա���ٜ����5��\�]*B/V��U����g[��g_���F^Mp��;�Ä�*%b��n�gk�{
맍x/&Ƌ�K�{�"���}�3:�Ȥ�V�M�cA��́Kj�f}���Ӟr��|�N��J:���Ps���6rZ;��rS��Jnv��)ߝy0&VF�h1Ӽ��^dQ��֕��L}����nĽ22y���	�y��%UL`9�GҸ{��.�b�FϨ�k �R��K�צ}¢�����ی�ج.rV�6���2���z)�+;��z^�Z��wLN�x0+F�Wp Let��)����k�wIJ����u>�{5��2�X�Z9���i�E�T���腭��y§��uZ;�G���Ys���wi�@�^�5l�\r��x��ړ����?�7GgX<6���k�^O=�N�Sҳ��Ro���9��{X��"�@��_1��\ư���o�*ᔸ�����Je�P�Z�Nr�^h��>& jˠP�wySk(\��ٱu,Ԫzʕk����)��1n;M,zk�'���vZ���>Z�z��{��g6��!�3��C�j�)��#�\Q�G��<�:~����WC���6�̙������db�|1�&�<3�+*�ר=���׻(Ti����G�]�*W�u�~{�L_S�luH��v�|�N=n�	�C���<��7�w��oO��\}�MO�C�&y"�+d�Z��Y֕���wm��l��E��+�h��`�A�T����Q]u��|Z*[�N��>��vkV)��ާcr��8y�ƙÝ#��.�`����kd�ѥ�c��6s7WV�V�*�i1��Ū��Y�Y�����;!�́�=?M\Wx���]R��o�FbX��G��h�4��8��:��M�)FZ���A#��qn�c�;+#�T*��^�	P�S]aY�&N�i�ّ��'F���{����O3��ۛ�B�螦�j�! R�sjڸY��[�A	<��|��LN}���?w	�������ac;��V�����U�JA���Ns���4G��
�����:�ݵA����d�R�J���g�0�_WVU��i��7������\pB��g@�qP��1�6$-oپ�e���s���߫��n.�SB��7�WEb�VZTŦ�W���qj���>R�̭�x��ߌ�}����n�w�j�W�#dg��[��|+�ۍ�LTc�X�
=��I�h�Q��PU��{A�\�M�V�cq�_ez���b�[b���l���� !������n&��{W��3��5�o��
;��'�{'����/'GVg>
��.��Z�z��꒯<�"22��(M�c5#ʭ�:ʀ�ol��}�4�k�H[gB7�V��p�ݖk����>-�����WeL�5�Fi*$!K2�/�t�A�ue���)���+�������:�re�Ҳ�,���'κ��M����b)ڷ�'�ݩ4��C	�'G�����R�Ey�ʎ^����������.������5�I��I$�M��|��'&i�)�ؙ�p���}���iڽnF�Ν������7��#�@�61;���G�ꕛ�Q���G��"�[��n1>Gv�m��c����z]p��<�n+\���V�i�g �g�kY=]ҦD�T;�z�𒓂�s,��V��mf�^h��Gnמ���U���:ĳ�Pr=o{&�u�i��[x8�C�{�*��yŁ[�7�8Q[�ة���X}Ҷb=�y�^�\�r�yI={�嫏���Y�����J�u%��G)ɴ���3�n]n0nk�i����T����5:ɰ):�R��ĻCN�R�2�+(5z�v����k����m�I�OF��6(����z�A�i�qȧgd�����՝�UC����;�
F�3�¯�4jL�B���,�a�h�͎�&M���c��.���lu#���]:mv��5ϏXe��M�tsV������^f�B��8�gy���{�ҟ8��S��S�i�y[q�����:Ŏ����6,D�ݝ��f���̜����]�sje��r_:���Y%�0��a�U�ݙ�v��x��9��^���s{� ���_{����k^��nb��g*�-���㗺!	�9	�%;4���Wu�we.M�wݘn�I�8�G^P�r)Ү�on��@�u1hZ�*u�]���&�s7v�c4��o՘h^>�Uϲ�W�G�^um�W�f�!8.a*)�x��{�_W=�Ο��g�+Rab�=�=r�q�2(S�^T8��\6�ٕCw|��������zj��h}�G7�!�tN�����{"X�=���^�}�F��l��I��ՙ4�כ�Ħ{*�q�nǁ���c�@�L�Kýqw[��y�k�{'���I�y�����<^-�'X=Ԃ��v�O`Tr!ꊇK���g�[���<��V6���=����w����y���R��Pq�!qY���{Y���ݸ-KZ��nNL�~�;˗c�v:8����	��y]*��i���0�پA-�������Э� �C�J�EŤsy��bD^!�SS�B����ٵ�y��ʷC����$�h����
����u�����머�57+�z��oX��e]G���N?���C�ޤ�y�K�F}�K�<�������䆗4�s�g'�����g#u����	�=�^�	VxxN>��&S�)��u֡�����W[���Q�^U�5��6�K�y���	<4�xE�Qa�y?l�`����T9Z\q���Y����s>��s
�S�n���7iz��q�K�m��!Us��~�9"yĊ�7N��ɒj��D�c3T$�,r�����_�F|G8	py��[������^�]l����)��"Zxk�h��ĵe�C5���WI��Z`1�y��1ӊ�Խ��Ym��}�g=-]��D�-��L���W�g��,���Ql�ϒ?c�ޠ�z�F��>*}\�:{�<�}����Qw�1��NrdV��r���3Y�@�?OC�Ŋ�.�CG�����u֊�[:p4Gl�y�x[��ݧmn���3z!n��l���R��♜�*;]��7w�]��KJ��8�Ь(՛�E��)Ső�����珐/��]�eh�u���ݧՏ�&�7g��.������K�2���=�٭��o��s|�CӨ��M(�ݡ�����ky��,M�zmߞ\}��vխ���Ǚ*���!ey�V�(wRw.����{�΢h�e1��}���KNz���ͳ�2��t��kh/md�7�S�	�¯d[�M��F/��m�:�X�=h=�;��<:b�s��1=
+vp]6�-�|�s�������W���6�GK��V���k]�F �*����q���]0����+!��qi�߼%��A�V,�|�<r�U5A]>Ka�G��I�z���v��mb~�]�h��3�'Oz�F�����*o��W�>"B�g�	����0��|�z.s�,]��׏<���gq\���;�4 ���C�j����]6*˱���<�d�<���'<'-��疄�d����Xu8�a��R�b��f��t��������lz*���uH��e��v� ��]yJ�|͡ >z��`̬4́&�W�q�=O�Sv��H��1��}������:�00w�[�x5�մ�hZn՞'�Q��:�uЕ1VR�M�P�W����z��w����o��5w]lάm셛�͋� �f����jn��v2��YMk�8=�m�"V%��B�'C�M]Yػ����%�2�yz�
Ǵ�F�PEQ������x3m�Ղ�W^�lƦ��GH�sJ�8Y���� �Fl4��|�;�ӍIwP�	�i`"�s��Ŷg�)�8�U��$��b�ߖ�s�a4��Vmw�|�uZG~��=���`h��yYxҘ��`�
����`�9i�Z��b9����uZcuj�t�Z,�]팩�h;П���S; -f�#�%�,T�!W�2��+�Ul����J��NR��oִ�x�C��&sC w^�rFd
�d&a!o�b�:W%݇����tnQ�E�z+��S����O��zg)�	�A�g�t�cs�ol��6���)û��&��o!kV�a^��m���j;�j�*��*�=�It����u�cY�F��y۶L��V<M�V@L�0 1P�O�x���,&>��n�r����G0
�W8�IYM]��b�]�vf�����l��p��>%h���̚������������\�$�Y�7�y���.�ǌ�	��w2`Ո�B�fmZ��>ݰ���^�`��8����WY}��z0]*.q��z��'tEKH��p �υ�S+4�S++)٤�{����Ej�O^��Hb镟e,P�(��9D����
ad`���u���Y��f*)80:�eʼ�X�*��Qt��IR4���l^QI6��Q+˧F͡�j[��+a�e($m=+EᇷYu{!�e�f�h�ȃ9�q�Ô��ư�6*�t�Ѧ�!��w>Y���DIMf�"\��������15���h���3!��o��$����n���f�2�c��lv��V�ȫV��~őFY6k��ѻ۫i�l�aTcOE]C�%���[��0^���+��A�,N^2����>c+�*��0YxY)B����% U�Y���m����]��K��$����Ab�GoS{"V��@�<g�0Y�*�3�B�� v�l�u�:q^�s~�n��z�^KGwq�����C�8�/��Y��"��X�H�ǐE�e5�;][���촓�,�(P��EuY=r<������Ɔ��Z\/]ܥs��z[r�f�Yb����Vٌ����
:�d�e"��*Q�q���5T&]K*�c ��GG�[u�	�8X��I�����P�w}y�F79L|�qE[}�U5�q��-S����"��2���lX�ł�"�����S��QD��%eE���kZ��m������!EaZ1�E�,TX5�*Q���"���Q[s%b��b���q*���+ERT�,Aj҈�ʂ$X"%�U�+��e��������U��`��e��Z�ER��.*1bE��"��,���(PIP�� �"����3X�J��QUDE�ZTF)m�F
1�"5mR*E��J�ѵEEQ[jE��"�UdcV�"�J��6[P����ҪE��*�PFZ9a�ȱb����db���R�EP33E� �VҨZ[Z�amQB�J�U&2�������am��kZ�Qe���R��R�F(��)DJ�m��+"*�FQF(�D�ebł�#��*�5,�"�aFLkU�Q���DaQE����b[c-��b�-��+X�X*����Pb*z�3�}��ϟ~�̹����]A�qQ�#V�n�W��u��\��ޘ�X\�y0�,��-���#
;ӛ4Q��-�_�����M]�ӽ[��DF�+
�|{���#��k;Օx��@�;��ϣE���J�֊pz����w�zQK�~+�}����n$��8YbԒ�̑6������H�y�K�<��E3�q�rEn^z���#I͖{�Fۑy[��E�������˨�%�^�G�����ie�(�7!��허z���~(������@�8�C6QQ�9��TR��������Fߩ�N�g�t|�o�p��W�8<�;1'�ֈ:�j�{�%�E䩶�u��εu���e�xO<B��۝7G7�G4�Ǟ��#�-噂6�1r�Ĳ�e��	��d
W�P�*gDL��`ߝ�j��2�:�'�7Q��!�ݺң�������������C��0<��m��i�}�|J��5�VuN��Na���A\�t<N���F}9��5���#DN)Y��D��ֶ(������P�S$�ƺ�%�K������y/�B�W��7D�S[�)j�>�^����s��o����s�ى�Gyh�w.%������;�8�0�BE\��m��؝1tQ��kD�.��8�[q]��o}fU�iݥ�J�%;k�;Öes��=�)���2��R�;Ƕ�����}Lr��Ȳ�OD������_8�M��3��)�;��7�z�7���%�R��tSp�B/i��{�{��n��T\μܾ菹m3�.�2,9f'Q�BI���]�����G���0�[��a�L�M(ˮ��=iՙ)�0X��u|O���4��ZW{�f�Sn�6�r��gJ���.\����Ce�X6Խ��ܘ4,�(�n��.�o<Ww�G�bw�;݄R��i�����ݒe��Pb�b��\��S��7.2�������٥>�X�2��u����xg���)�`�����(u=@KWR��� +�h3f�s�rם��N@��V{�])\���F�Y�?*�7(Z�����%��Q�;�Tg:Ŗ=��yi���%oP'�d[�#^hmqy�ȭ�Co*�#6e�D	el��t�p��,5�~��jt�F0tvA���d7]k��t_W���T�ۂzz^q/�p�x�+k� �@o�Kf���[��`s�|��0�s���}�@�{f�$t�����jſc��@�l�MdiHŅr�S�����{6�P���hv�3n�m>�J�0�:{L�ׁ7-��ƩN��X7ž����݈e.����"�ۊ�/];��ۖF�(w\%��T��гc�i�[0t�$������Ti| ��c�K��X�W]N�e�S�5�V�z\%���������-�<�A5�l���|r�e(;Kz�y�[�}j̬�U��]:��k��	�#�]OR��.'���8�ƹf��Z�.�M%��VrE��/��J���9�d�� N�*5���]+��|l��y��u%���=Zzܾ���{�m��^���U.b7�q��]p
d��_�� �cr���V�<�}m��_sad�˚V�����C�$[t.b��\Ob�f{_��eZ&�(x��:\���J+yr{��W	�Y�`����Ϭ��}H����ؓjD��ADPo҉ʧ��wj�D��v�oevT�����)��(W�
�8U��m���銞v͇��RȀC�mfeEk���-V�Ee��̼�R�N�f��xK����)��}f�E(3�Θ��`�뽣3�c6�s�|�^
vI�M�2�Pw��o�,�-8�>U�1�V\T���c�pof`��rE�k۲��t4e�I�F/E�^u�J�[#�|v��֖������U���@x����V������1VJ�A �b��Zѵs�y���X�P�t�'a圪n5�^��<��:�r�N��LN�Zg�2�4�;Bl��=K�W*텹vɧل	]��O5_�Xj]u�7I];R���Tw7�t�13@�f�����O�&�.{;4�a��*���8��N8ȊÕa5�`׍���Q�~nŏ���!G��SW�ekJ+|���A�-߾ײ=X^+�P�UAη<�9]��Mt0Fo��H���k��5�^��a>[���ho��{����wb��rqU'���ζF�})ȩr>���s��]�o��Z
v`�E��Y�gG��:�ү��ơ��cr��b���f)�~���Ӻ¯����A�]�6�TP(��N��e��`����E>
9��dx�,����E�S���y�����/�`������G�e
�ut�Pp]Ž��4+/ZE�DY�I�AT�y̎؛ԭu%�=�BP4�GFL��ƄL>e`�'VΈP2vߴM���X��l�����-�#�s��
fR�
3��q.�M��
ޫ]�E�p,��f�+�Cl�xX�ty4r8ϳ䫄>�@��vXjL$d����N�^f�l؃*G�]w��Oh=\�a6|�IC������=q��K���cu{��1�i��yFܑs
�ڄ�li�(m��hY�JR�@>{nq�}P�5�D!b�#�0ct��P�ٷ�:�E�v��QCK��ְ�w7��s���]:k�xc�����[��N�\k�Ҵ�Caw�P�̾#0�;s ́]��QB�� U�.�Wv�T�">�"1|�Ӑ�i�Ǥ�ǖ	��f0��W�W��]y�%kع4��W9��خu�D�F7�D��):`;������Ꮕ9���
$lVz����n����@��2��Y�h�͡���g1��s��0{i-&�\5O�����8�S���,�~b�>�9��ݵ��NxPV'z��1�Qf�Xi��D&,�w�6PO��S�[H����w���ܦlnM8y�L� jb��T��׹(�^�����^Iv$`�~���7&�({�9K���_K58��_�WU������mQA*z`G.���Vh⫫S\���;����mh��`o\�<+�H��In(f��J.,*��DXgeWV�����N�Dd�=�R�g��E�o���� !U{3e�l�.�^����\�O�[T�S���^���̻Q��M��v�b����!Vp�t��^T�bGL���!D(En,�$����Э�����~�+S8p]\�'��9o��ذ�U��|A��~=|ht�شL�<�ư��h
ӚYp1���B]�C�W��^5�q���0։�d��.՞��˝�^��ޕAg;͵O��Gt��]J�Cn;=��2�����$kkp*���Z��˰��:3�v�;�;�q��,T�{&��ᒰ�6\�N���ѵۑA�3Stv���}��{���w6�so'M�!(��Q#�F6��p�.�ޭd��S�GAPt%;>�b�cw��a�t��l�n�L�ƭU#b\��cdYF�J�y�tK�N�z�6ȁ�"��{�qۧ�'���>]-��}U`�=t���K�r��傅��a�(}�wH�+��$����Ek�ë�]7W�s}�,u	�Q���V/HT��>�u�cBء}T��M�fV� �^9�3s0���I�h�&r"�:g*)�� ��?c�
41	$2�Y��C9w���C�V��&�Z�"{�=T�_��~t���i�t����T��<��#��u,%�Έ�N�eݎ�qg����z%��m1�W������~�Cb#�����ڗ�"�S0k�+2�u���:�8u��)Ai�t]�娱c��!�@/[堽}�r�ר\vG��V��IK4Zi���n�Q>�*F%VQ�zRZ/����.��$�@t��0T��=���:��6��6�=��π7����VI�����+����u�5l�#�2,J�����I�7D�x-fBŞ�0�@<��ꊟ��a|�*���k��҅T3��H-�Ko�s�Yk���b��ϵ�P�t�uv����+/g��.>�"�t�	Ţ��x{����Z��>7� �k�X�{W��>Y"��}Pa,�2Z:Zf�+ێ���+�@
L����M_Yy�R��i\Q����3��S.(=R]�#�T͸� �1�w�n��D�z(P͐���p������:ޭ�Muq�BF�\�s!��TH�)]:�žNw������Ń+e��o��{�Zx6�t�zc>�9�we��Nnԇ|OxO>��Zi���s�	�&�؞5j\B��ˈ�3�YJ��S��Ke,��(�Ҿ�i�k{�����̭�ԍ��L*��~>��0�al��Ug.X]�#eI�;{�"��z�6Y�������g�*���C�7�
sC�J��GF�xW�����#X�j[�Z�ul=�G^vO�[޼Q�]!si�`�L ϴ�
�e 6�c�i��B���z��v�����؍EY��prS ��W����>,:�'���f	�y�sMv��U�.����eF�l�0��S�s(ۄi��1+�B>^�T��'39{3Ү��C'I�|��7�z�S�If�O�c�Ӯj��ډF8�͘�˩mY�@b!�yP�n�}0�
=���iz�b��[�q���ƹh)*J:�ju9ؙ���ӫ(�O��l��T\o"��������u�s8s�+si�+6�����X���K��{��n���./�����XK�����,\�B�Ң�����R�O
QF����R�s}Ϛ��u�F��:ժ����0n;:W�f>����ʺ>x`6W����K�j��i1���nMh+�T�p���&����҆�1W��5μ�?
_LT��;o����g{�^��W���V)B ����^�9Nz����6����q:טo�Gcd��Ot���e��̪�P��{X�4N2!�n����!Ő�C'K�<+2���Vgs���3qy�`�͞Qʳ��N�T*I⨯���}ح>��i�:~k;4�*�qk��,��g��`,��Xt�c�6T�hf�,lYd���U������6�!8PfT>��i�|gU^M�7�i�F��Bv-����V�W��Bw�`�fAW���]���-��g[�:�+{��;�6J;b5����LDu�:�b~~��g.$w������X����Z{���U�i�i_|�+
e[�L�g��E��"���2���T�^�zY���,:p��Ӗ�v_q+&mwu'la��Mmd����s#j��tӺ�H�vѯ/�=���F���v+�7\��t?���%7��˻�C�_i,(�c��
Z��8:���v���O	;�R���yX��-���{��Z7=�������5��U��(�߆�tEަu�Ys�H��67���p�:���tΊ=y��b����%��{�Y��h��EhK4:W��k!�}:���m̲!߶(lE{8u3f���V�T�ʮ;���U#bb�b�����TJZ��,8
�u�޳Y~���'̓�c�)��Q���xr���:n��L����Y��,��垶0Y8a�и�<���.ۚΊw��ȋP?Ht-Q���L&���+��>��	��r�>�/��[�B�u.]�/���Ň�V����Q�m9�"�*F(9BF��;5P�X�DU�,���Wjw3�g%U���L㡑Q��3���N0�P�l�	Tp��kÄ��'Hϙ����77���g�.��pfҼ�դY��.�<�]>��`7�[1�b��`ϥa�pR��%>D�3��l�҄�>�)�@o�n
-[8�}x�^�LU�R��d��
%!3�ٺ��{���-�D��G���'���Q�����4Pز����d���u���d�e���W`]���\�0qa�1����I��1D扱-B��M��D��\��,�F���[*b��	l�H�&����,�^�[�׫yK"�����>뵸�މs���ͭ苭|���Ȭ�-؆qQ]�S���6⎁����
3���ꯨ���MI��^W��y�_��2K�l+p��#���ʴ�o^C��lCL��ρ�4�Ĥ'�TݿM�=�j��Q����{�l��fˆ�e�>�.�IO?[�0.�kiJ�*(�:\Z���)㍇ʴW��vw����I���ӶtZ��V*�vk[�iOt��_��y��6Vcu'�5�>96g�o0x��R��'P�/M�������Wt�m׫w��hOpH�)�<(�8��R����LR����p����>�ͯ*S]<�+_82�.'�ᔼ���V7Pp���6XQ��#�Os�k�ӜZ����2���HTו��%��:y�0a�e�0S�oJK���4��od-=���'��8n�t��s��N�
�s�Izy]�Q�`�Vt����Nb�k_{��_�q牺�y�߭*�"�Yf+�H(ϭ	$2ʳ�_��S�W!��%;�S	��k�~�����TK�����`��̋�:f&^u|M�U ��xa�y�#�����d*M��8Q�]��Y�h���RZ��♽�����r+���A:��(z�*���6��颺�s̏�r؝�j՛R��&YTՎ��r��^Y2��5|k�x��:�A,;�};����4�<]i09������Ӎ���썥[��b�o5�O-���Y[Z՜Рg�]Ytu�sZd
��q[{�jy���FL�f�#k5�����&Y�Ӡ��!cu'�ƚ!էp�)�`�Y�C(ǢE��TR�CP�f_�j$:��[Y�Sm�E��/�w}z�(_m�q'׋
}{v��]���Pܠ�*�f"�6:��U���N �1�7��������,��!0]��S�{�1�:VՅܻ&��k�«������J��9R�Z� o�ہ[ �I��R��7��b}��2���y�쐚5�f�:=dv�o9�Nٜ�7�5E�+W2ڭ�v�9w(�Ҧ��μv�����l� !R��k���$��g{s�n���K��ӵ�+�5�G/�>�eW$�2�^�R�.���ڙ�՛7\�%ޚ�n����򋝋X����ڌl*�v^�10�)�����+��k�`|Т0��W��3y�K'��]��x ��R�-��I�����c��rr�;!N��X}��[af�y��N������GVJ��9�F�A�m��G��bik�>�t�r����ҝ��%Q�F�_o\��ZqejE\�IY���
1@��q�e��]c�o�8�������[��7��������p-��;_���/@� b�W5M�Vrok1Cv�_�"������qq�h��`�gpL�<��
��t���K/'T=7lq��˧�{@�ٽ���d���>c�+����ch�,⳰t4%v��;��\��Kf���q�/���a*�HNǨ��i�xK��� �4���#|ﶆ"�5��v_D:�p��靖�y抱�>��	H޵JFA�ݵr;��Γ`V����8Q��Fc�c�Rv)��8�K*������q o"KT��o2	Iv�(���F�?`��|�H��uk�:�W���\oM��Y����l���L�T��ݸ�g�	�k:��4$�帴#�u�R0h�i�g%ˠ�ڵ�g�vf���g�O�����ĩl7�q�R��N���c� �m-++{�$qX;�x���x3]#�d� �u�7i�l��r��f�v��J�9ڳ`��+sr�������pA:B�����16^=5�#��h����.we���``P�ӥw¯m� �YX�soh{M���^Z�4u�D���B��3Qg��\�p�wg�F�/6��:(��r�̭�CF �U�/���n��ڬi�ko�I��xҩ�[x!�ZM���۔��U��k�����?��5�*��=�˭w~�&�^a�7o�ּ*��>��ն�H�'�]�;��ZP�'1.J�� A&�Z�-�Յ�DQV(D@UV("Q�J���E�"0b"(�,`�U*J�",kX��@Fe�\`"T�EQX!Z1b***�V4�R������1`�X�EX���P�m��X��("(�Z�cPZ��R��1�"
( ��т��-h�J�\h1�l�*��[R������b-#Y
"���Q���(�Tm�X������YVʬP�b+�UX�%m�h6Q�J�mJ�HƤ�Eb�-�Q�"V���-
ȱE�"(VU�-j�E��"���B�[J�����+
�UTal�Q#(�E�Q�F֢����AU����QQkE�Uı1EH�[�UUV*Զ«QH���X�"�(������"��R�B��(�k)Eb1U-�E*QU��b�UA`�-*�Ŋ"����b"*�@T-(���("1-�J��*"�*,�TZ�m������Ȣ�E�TA�.%QU��QV�m�X�A��"-B�U���V(U���R�DdPH'���Lʌ��
xr�=�&H)q�Ht�B�-WZ�pXgc�y�=r|���=���U㭕i'1�:G��meİ�/��  ��\�kg+W]:k�G�K�Ãۊ�d��XK]��7���H�J���;t�w�VL�n�n�3n�֨.��ޤ�Ir�j��i��L8�a�LXv\�㪢Rg�lz6N7˭�<Ksx�`�N�U]����Yϟ/�x��p�O�(u:���q�F9wu����]^����I[@��"
�v	^��z�.����[��2�Y����]�K�Wc8��е��p�y$���(�p��4`Q��O�����b_��X>k�6��O�S����qG�n�������7�q�6�ތ�8Q������,���N"o8�Ogkէ�(�<��ٱ��S*�[���6��zl���:}�9ͮ�w)�C�a��9s:d��4-�6&��!�)-�4�z�{������>�ſ{{: ����p�*ϴ��xl9*�4X�P�j���0B{e׃�� �mچ=q�͇����M��n8���:�T6��4��0��dP�'��Q�������x+B��t��T*�����6��Ȼ�`n�񑵲 H���7��K~�ur����*1��ے�^�-Y��&k�t�����o�^+�H�wV��o#RV�]5).����gnuD���z���KlcOa#Fi�Bi\��L:��ћ��  	��%��G]�o�����N�� �-�a�T��p�u-�|�
F@�v�H����̇ǣ|�;5����s�w$���/k=.b��)�k�4X<���KYN��2��%෋�;�3�_�+�>�a�*�����!��xH��T�
�K"P�`��>��a�:���s{&eM0C�E04�_��������x��<i���H�9�cQ{��L��8gx7ӬD��0�o˅�'>����ߖ	B�_�B�����>��|U�� ��P��]�knN!WN� ���LE!2�tC7�Q�~�u�oe��9����������k7Kb�L�y,�83��嘡(M8El��Ԥ9��g�e[J���i�u�qk!��%R���A�Ġ�3I�F/E�ui��E�R���2tFT�Bڔ'���y�S}֔cy�l����CGH.$tk&���9��at> Qwn���ԽޤR�J+>�v,g���eYkG��תe�Q�����|�Z�WRD�򏦪��ݎ.�YI��)����tdv�^w��.�+�}��?Gu�`AaMR���C��q�ZhonQ�N$�i�$^��]�㸁������ӓ��3z{��ý�����гC���9ڱ;�����c:h�O`��g�̆yy;���꯫~���E^����ן'���;v).�R�c���`�,�#���SC8�V�̜�y�\�nS9{�:258�"߶��E6~��91��v��	�`��ƴ��>^�3��s�	2غ�u�],���O	"���`�@���P#pS�ڨ���fM��Z��{���g���H����i_i;J+E�ePuE��h����(lk���|���"�zꆑ�`s�u8��(��:�^u��q��������Bĺ.��s��'�4�r����S�4�ԻC��l
A�i�jk!������әdC�lP؄o3�\7�bެ��1.��t��6�S��)4r:ϰׇYٜ���{`t�;��&@�=�Ɂ7�E�c&\Eb�C����;��M�*Y��������5F'���� ���(JZ�{�"��*
�����h4W^�ᒄ�<���.�%7o:[��W}�+#]*���8�[�8��L��*F)Ȓ�:`;��ɒ���#3ssz�x�=���wk=X3�l�6/18�a�J2/y���7y����-<gݼ�P���f#�Cb�^搭m8����gF��}��ӂ|$�}�2q���ᑭ�5X(r.�D�i��%	8F8�=Y]1�M�ͩ�MZm2*(2��k��?UU}�/���8�{�F#����I^R2�p�S6x�`E�����3�x�<�d��i�WW�#���J"K3�����^��5�0$'""7������ᘩE�.��^�=Mj�5EF���q��T�x^�#~�L��I2�V)$HLH��ᅱ�������^�_�^;'�'�%�B����x}t���&q�+����LuLV<<,)%������������7/t��ݏ����r�$�X���xU�~�-�{6h�X��#�r�U�h�t��r�¸5�U��S
�>���|���wpk�	xϽ�U���UC�~���{�Z�;�c�{�WD��zˋ���H�_)�;�v�b�U�5�7tJ�b���"��8�a�|�YW�xna�8���i�E+�(�W;��-F��˪;n��'hZ~ݓ]���t��|��fzպ�ղ�Q��BqZ��Qv��Y��ʱc*!-�4��U@�U�r�nWee��`]���Op����K�S��/.'�ت�ኺ`~���$��\]g��G4gdI�5|���uq`���)gv���u>)˅��[�73*٩�'qnu����܊ӥZ�
vskj)V��ح�����oӸ;Z�bͩ��[
R��&��3��6^rx�bc�>��
ۘ���-���mo=4��cY*ܣ�^'�_�v��Yo;��0��b{bz3��E��r�W^ٔ�AȕZmL�B\ڇ�2��>t�A��~�q�v����O,�-���-EL;�+�W�*s�O;Z�%��`� �iR՜��m��{8�Vf�//�M�d��~��Oy��bD�
6�C,�F�ݩ��7j`b��O$�=���^�WY���3���mK����nٕ;�Q��_��#�>�+�N��,���<[�tQ<޺!�����T�++�:�N���'A�v�Y��3Ґ�z��R{�-������2����"��娺�c��S���88��rܯTg9��8��J��;��z��.�W�k��	��S��,�ϗ����.���u��{�Ӯ�Q&�7W�xMT�=(�)�1qA���bS�h�����K�Ͻu��JN�պ+!p�[�(�:����4X��K�x��3�C��������X��Nx��7�:
�	���}P
wA1L዁eϻi\QZ�688Ӧ͵$]{)ch�t�B�j�~��Z������]b�9�p��ږm��qt����2�"c���yλ{M�A�����V�O[ӷ�}	]�]%K�y�ֆ̱V0�\�[5�U�e\N�v%����t�C�:��f1��1��fd�x7��c�X\��������{5���q!���F��R:pK&�C������[����,�w� ���������{��3}��I�`��{N����F��<jܰk6Y&���#
��]���`�rN*�3�pmcp�9�7�9¤�1S���U��8���Z�s�=t|<L�Lt�ɻ<t%��{J֜��v��}@�xT��{�\��t�0=��[ƽjTB78d�ͽk�~3ysqu���q�0J�lO}1yq�W�B�F(C�S'��J����]k��e�����u����x<�lN���V5�>�[׎7��;�/M�vX��BP�D%�u��G]��󒰫1u�gd �z��5����kf���VxH�n��X�=q=�E38���8��w�G�R�X\tY��0�:�1��z5�r,|7<���Sޒ��{a����i�wne҉՛a�X^�f؞����,6מ>5��Ьt�ׯ����VD�Yb哋����r�[���'��`WK"�*Y�B$,�hWD3c-V<?j�/z�,�x;�{
b��uX/|ڪ�w8�7�������÷m�&�c��fq�J�mc�w�GXPY�B��i�!r����[a�����Z�4m3�j�|^ZS�m�ӓ����8zcZ�#��Ʃ�v��G�͏�ϡ34��#�!�A�*<ǫ��߀����k�a�d�t��`�5�3�$]l�,�4�$ԩf)�b��&�GD��o�y
�K�CV;�:&���1S[> ��l�(1�Qs4���.��E��*�8=��9��y�G�����6�M�[����+�G怯Y���5P�[����XL��bߵ�C٤�f��qC<g{�1����T�o�[�c�YL鼧Lح˶x�O�G^�ua�y�:{W��Y�J�4nv{q��Wgm��hIC/��x<�n���hoU���g$�E�K*��.6IX*]�O������<��e;dl���+Ҏ^��u�
�U?y��Pw������s�nlfU��ם5�G����J���ڋ�k��L
���f��ee
��г[�`�@�U��罜�r�tU��RݔNr�6l�1=38WR����$s~Q���}�~�b�`����<��=�:���ƽ�dut�+إo�"��l2ktܪ������B��o8?)Ƕ����ӓa'@U���*��`��Kq����,?+��WS*ZfLd4� m�rY����&�5ԭ� .�sNۻ�s�x_���T����zׇv�yf�q1h����:S�'���,d�f����8ءD����p,�A�<���(.Wǋ�x���v]t҆Z���RaSz�P2�ȷ�> rPTZ��՗�}���{˛�K/0(���쁬�t�[|.3�1��B��2�@�����Qq����{�u��V(�ō�q�~�ՌW��9���R��Qfz�I�#�թ/n7E^_c�n37UmE����'W�T���21��Z����،�:n˖Q�l��b���$�uiﬖX��t�<"����e����ft�P�g��!P�E*z��w��[�Dʭ���H~W8�B"���`l'������l�N0Y����5JH�V,VQB�Kq��6�kE�&ɞ���ϰ�U,y�`��"b3����:�m�8f$�LS�͖����I�v,�D�`��)1\+Y��,�v��p�J��E�+��eY���(T�6���]�ݜx9/���l�^�D/�X>�Ҽ=i},�8�nyߋPܝ,��t��"�1>&��ݑVJ��U�S���!��@!��#6����t�ե�)�ٌmţ@��:\)��u;���0鴶�"���mY$/efˆ�g픢�=-Tȧ� �MÞK������G�P��U�tss�Z��'Kf�|���J��9�w|�k�b�s[O�Jם�4J;:���*:$�{�v��E�|�N40��nf�z�����TYnj�����8dJ)����������,9�u�5����Ά���  �����o�u�����E͖�2���Eڑ�8��a�̊��tpb>�)�]7 4�s����[ۛǪx�_
h��)��6^bu,S�@��5��}c�[^�a8r+����A�mҭ޷c���`�IC%#2/�"��s:o�ۻ�ڣi�{�<�ĭ�����R�啉��82�%��\��vb�4_g��s�<N��ʷE&�n�q�V��W��Y.��}2�Pϕ�G�tw�c7.mC�YR劽�GD�>�A��q<ۜ�g!�Z��}��a����G�J@�>ʋ��F���O�/Ȣ=���:M�܈g�W���S�xO��3zY.�*g*0[ufE�e����(ױ	$fV.M;�j�j��������0|O��Ch���C�R��'�R�xI��yQ�B�3bt�hS/z���h����z �Y>�r� ���.=9+�O&��Iv�
~3���j�w3˟�\�Yz���<xk��:��薂)|�j5������f�9���*휪b���Т́��>x�*�wm�{L�0:����-=�FuwJ�Þ�rmJHb��u��u�=�d�e�5��wL+f�:��]�q*]��Eۢ`r�l
���W��NXI���і�}1�u��%�I���Ǡ�"[٘//H����iy��=���uO�'B6��T�@�>%R�o�m�ږ��/���`�����u�l�e�I������v%x��l����E4f��50b|֛ʓ],����NF2��'3'i�9V̕��ќ}𰇩�Z����,_�|0�Q��Q���2:�B)�9D��	�yU9���s[[��\�yC>�����Lf�}Xj�\͎�+þ80A=ȃ%����$s�J�Բ�A������:o)�3d k#Jf»��[��~{��!�(�����]���j%���c��u8�Ӂ޷��:�����L> *�e���b#O,�&�!"Z�<��qao�����C^߂���8��`�jf�\��<qWc��xOL��8d�����]"�*�e�	F��fT�=#XT(ad9�\S���yV�.�=�x���[�̔%,��u�0g��=O��d�{P��,��,@��C-��������G���>�YԬ뻮;|JT���gVvO�[޼P�Ιo�)�!C���Q�u�lTn+X� K�U�BV0���@oAΑ�t�8�e��D8(�c>�m��6��j�>F��N�$`�/K�LX�lr�p�ۋ�0�j��3�c�S\���5��v��w��ǲ�i?q�e@	�����Mٖ�	U���-�+��`;�&�kw9<�F^��;3a�*�MM��n��i|+.u�g[�tӴ��n¾������3��ңI���)�
����Y���uIB���*=�J�ŷ�Pܰ�5+u6Q��ط#4cN�(���$��87�<� �9F�y��0���{�Ŝ��O1G���:�o@���񨌣'1����u��\�����T-����4����ϝ�@�{���÷Yk�j�B6d�×�vu���݇���91���h��t9��i	��[W�JD�;��&� :����I|�4l.xq�j��Ñ�:[踚3+�]�9��g1mĨ�4��4��IGM���1�ٗ�з�����Wh���n�.��|�<��������g-�4����Qy�Bt쬽��ƹ\�lwVP]�ҩ���4~&ugoQ�79<�z���#��Yi@�O��`��X�es�0%�J��/8���E����C�����Ù�%so7䥌�Ɩ1�85�WC�v�0�Q����mѣ��;#�� �6�|��'�a�8J{���-���L-�㧣̫r�| �3��F��-�7�� �:�����C �j}b?�]��Fm��>�
�a�zH��yeVt�q���3C3�y�}�Cw�K �p�����.�5�W�)f�Z�c�tބ&���Yup�,o+&h�*�;m��#�a�ڹÝ�b�@RD<�_e�}g �V��w3��oɳ��[�z��crN㗔�&M��Pv��Lϗ4w'{�.$z�\r���F� b��J��8Z�,	�5�p�WA���{�~鞽�g�+O�N(�]fV��oR�@^����y��R�F���l,��
�4��9c������Y��B���RF��e�n����RV2V�iT�8����Zm�T���:Y�/u�p;d��S�7/E�ҝO	��V-��4T&��6�ɩ}E���`��Ff:_nr���/;>��ekب�VX6��V���7��x�V� Fׇ��,u��
���{X��@�d��ƍm��NwS|V.����=��t�և�w{����G`��_p���m�\F��.!�[J��(/�I��V����\S6�c$�5�w|x�W���{��g0֮�N��9�,\�:w�9oK��u w9RλX]�@]��K�}i@뼸5��P|qX�9�1�cAf�����5ɾ�R���i���AV
wN�w��˺(fe�f�k3B�|V��RŮUǋyۻ���$:�f��i�H��1�#_E�s/�Z��pҭk�5����I�܂4g���֖��?a��*�ӎ�Cդ��V>}s��p��W��:>bpk�� i���ح�G����0yݔ�C��1�WXW�M_S�wGj��[�[Z�m��u�o{��ATQ}�-,b�EQV
 ��F�����U�%��X�������"E�kDPVҠ�ED�R*
�jUj[e����_r�q����E�US2�(�KeQQX�"1D`����E��*���`��RҲ���4�Rڨ�QAcZ��$U�[j+YQEҪ�
Ԩ*�elTX(���m*�[-�Q�Q��X��-T�b�3+fR�F!YQEV0V""��*�EҪ��KB�mV5�AZ�X�V(�QDPEA�1AUDH���#PD��(�2ұ-)Z��H��ZJ+�+R*��e+Z"[DA�*�m,V*#V*"�VA��b�AF*���F1`�b,U*�*�m��[h�#@��-�ED�X��!iH�������`"�2�D��EX�S)E���P�X�"���AUD��T-(�-��iR%��0AU ���QR��[��z�y���i�w���j!B�P���yޮ�L=�F9,s���3]��i���+������&�{��S7��	������mzI�&L���ּ @F��k��^�+��b�A���Mȩ��;q,���.��2��61�׷����s�l���`Q=��2��=��2��F8
_E���6����B��"��eW������|�_�i1yhVq�`��{��k�r[�'�-2]���ڏ}|.�x)E�^h5���~�+�Դ�Rk<W�
�c����ų��DE����V�#��T?p�j���1>��
�
�pp�a�۫ʔ�κd���� ��˨l&�OE�$믕�3FX�L�WB�
�Z�1#Ћ9;،Y8f+΃ ��0i���\���I��7���v��՟nŌ��[�Tx�e��f�!�G�t!�Ҳ������wpV��s�B*9V�z�-�����>��ᐯ�nΐ�W[�)��N���;���I�GfQKU��fY�ޔ2���x|�v��Zo�R��f�,lYd�� ��^� ��A�EC�ϩ>��A�o�;dOyƑA�2�x���Dg���~R���\�[9�}$\��K�@ѱ{˾�V�����K�k�Jr�
��v�e��6�]����U�x�ټ���^��#�����]�W�.�,���N�W7�z#�L[Ҷ���\��	�I�1���ۢI��+3�ǟZ�R�cUp�5g���.�A�auf����7��Іw��������JK�8�����)xBhY�rcŚ�9�gh�YGޜ��.#T3o��E۪�4�4��>u�S���:��M�hͽI����� }ϚF�FYb��Ut�PpY��d�,[r8������8�q����5�U^���P�nkP��Պ�e��X��8�2��V!ښ�E_Nj<�����DU�s]�iqiwc�GҴ�2s],c�2��f[x\3�1�, �3���|�Q��-<Fu���4�7�O&���y<ڌ���3�"m�B�%��%�e��3W��S*�w/.]xS��1e�Y�d3C��X-�7",8ҿ|��sE��<�FOor�2�#�r�����{-	��=\kx�U��Z�8���2%�f:�0^��+$>���wb����A��~��o`�3��DV�p�ê�o�8�1B��B���X��N,��\�-��������%��k�Q�xe^9�u�#J�ʉ<�]>�9�@Pot�FF+�z���+�t���<6��o)ť+4�x5�i����*�6f�����KJ�qL�y{3�MW�"��\S��(��E�U�4jwa�������E�Νv�Z�3�:���5���+:��]\P;G;L� �\e���ĸ�wj�d�ݑ#Ά��P�������Փ$�j�s���t�UT
Oy�4½���b�
��ch!]��t�"fG��>�fP�@��*"on���Z�����yv������NΛ'"EК���+������<���Lu1����G!گZk���m6�%ϻj���0���y�_�W��8���K-P��T@�0]sx�t�,��Y�gA�ˎ�].�qV�X��<�r⭪F6�Փ^��˅<j�G5tR���M��{[�&F�3���0xf�*,+�.ԅ
��h�};����'�r���K�o�ü�،��o�zP�`�ږ�p#�8� ��
,
�(׺��,��0P�os��+=�:v�z*���9�*!6�ʚ86e4-��Bܒ:�JF0�g�xh�:���eӌ��:�=��ko�L�ӎ����P�ؾ��ʴ�`��p���y�*����ʻݣ����'���� &E�O}���v��j
��PT��Cj���ci&��^�B��Ϗ�� �'�n+^��i[�<el^|pm	Y��m�s�)�K�P�e���x�g�6�j�>ܠ��mAXYK����)�A�H�eֶ��M4+m.\�T��;�Wմ>@�'u������<s">���(��w*Bwe���w����*C)��&w�x;uy�;�ξ���]S7U�*�yFq˗���s�����7�������( *J��t:�zm����b\�H�{��X�x,�<����� �i���nw�
��z=PG��'�3&��� ���K	G���k��uG˃�hX���\�y��T��f�����q�O������X�U,)f12̀P>f��n՚��נ��{]`\%����r��y��U���0��6�*E�O��>'S~�R�}%������>0�IC��|q^z�P��H4,>�Ib�Q.���,�)�u&+���Ψr�����ĩ���6�^YU��^�6̇���X�d���`�_�*�{Q�2�����w�o7/��A%җ;9���2���I��f�c�,_wR���k�ؿ8GM�5]dd����|�nfj�k ��U�1WZ���V�:+-�퀁��3�v1���5��OenѸC>o�u��O�Ӡ���`��{i�|�h�+eN���/P�> Ac��\&�F]{��x��v,��q��&�n�䑎��s������Ըme�R��������8'�t�H���!������[Ƿu��U�}$�-�^�x$��v{p��m�;����+��%�{O�v�m��7�X�r�Z�K*��@]2)����%�}��OE�hi�����NU��g����ƞ\*/�����nz��GFN^'�1�Rvx�c�~��	��s=2�������%(〷�6-�C�*0�pF�A��7ǧt�{E߾���:���5�6q�-]h��*چ��Q0,��.n�x4}^B6��?sO+hJ�j�7H�D���U}2}S �(y2�:���޼��Bӣ�� �$Tv�dQ�����P����=S�ӪĽ�	�mй�v��>����5�-޶ot[J��d��Q7B�����X2���0K+�k�,v���T��|Mjޗ6�n]���	4+��H�J�D7�gF1=@]:�;Nt߁�.���=�r�S�9j�u���Y�*0Ô��Q�߽JYJ�b�.�)��u��7�9�г0'	/�b�E�=�k,A~׵kbY���l���g�͒dJ�S¨;.M�%2��s=�����GD��F��+��]�+�r)F�:�
9	�DXh��t<Oi��]b���}���g�8J�B��%ܼ	�����MW%q��ؑ�8VZ�*N��(M�l0����DӮ���E��ϴO�Y�ӳ%v�c`� ��3��pJ����]{4���陓�2���i�]�B׽r�]|h����Ӷq�p��*T]߾��Ow�(�S,]��V�}�3�޷�����T��;p��{X�4S��g)� �C��ype�X����囯^BZ^zg�6�YH鱔����D1�"�J�q;vwY8-�����E�����t���5����Ј��L�^?^���9����o%�0n��C5`�*ۊ8IY�������{��4���Nx��+
��*�Ɋnx�\�PY�����%�L��|�M����X��{EetYڐr�k��L
���f��ee� ��_pWK؞�t���Eʕu�f��ݮə��Z�z�}̟���+<�I�|kz�<k�݋kW�̙�Q�^��֠qٻf2,pȑ\$q�ف��b�C���E�땳�dv��4Oa�ǚ�����Iv^�/.�B*D uK�td�;W2Gкd��n�g����{�Ii�8W��"�;��"�۪dGg���|:�r!���φ����:5��pImz�'��r��K����³��`�kO{��ltˈ�~��؅p4�Gb0z욾�[��z7��&h|�r+�CXW��]|`�.跺eM\�-5��i�y\Ŋ�V"�|��Tnmˠ�s��Q��������lv#qj��<6^��,�V_KLHFGkP��]�# ���]���<Ƌ��
[��ۼ��:u�2��q���v���
���1���lG��m:fP�� ���\�؅�z���UPV}'�0|�����k ���â�C�]o�߼�u<�EF\F�@sJ�t��"�"w���7k�^Y�鍄o`f�ߔ�u*�Ŗ��~�i�~�H�9C{�[�.��j:����"��>�yK�"=?�DۤE���{`�8�ddw[qGN�3����*�/>��Ȍ}�$I�����B���,'Q�ژ�d�~;XB5u��|�e?n�	�o-Y�1H�g;{s%�ᘡ<Y����D"6��T��(^�#{�NA0�t�jl;�ܣTS�ԶJO=�,
�g:ʼ��:��_�����|і{R�Ybq����;%����ٖ�Ds[;Yt��gJ�Is�ڢ&�����ʝ�j`ć�nMNl�kq�j>f���ߤk�N��!n��m<�E�{�ˋ
��]N�=��M�7ָ�<�E�+�y{k<�(�����r3����#~�N�����x�q��t�k�m�!�NdV[f��B�<��g>��i�&/����ك��+����C�z�:����#\(����}\��}�
Ҷ�v^��[�����'��5?b�߹�c����"��������v��4\�s���(������x��5���� �Y�C.�mQ.w-E]YC U�d����g���L����.�x�l����8|����]X�>puZ\0:3��O+a���Q��{�Oz��GKS�z��J�d"t��]�}N��ɔtպ�n�Xoj�.�h������u�=ucD��^3��Q��OCi+�Y,�)�or��J%��(11v^��Z���f��P{V���fL�/h��������<i��8T��g��N}�맕/�B�6��p^��J��1e�>�D������	xf��)j�>��ze//�M�d�r���sFC�Y�X�+[n��ݥ�G]��L�`�'��5�6d���յ�HYw�ד^�aEc�]��rn%ˇ��
�V��	�q.��D\�\-��r��+#1ͪt:"2�cD�v�=+�
����l����$J�`�,�P7��eW"�2��(d#l��*B*��I9��M��'�%�7
�لBC�\���7&)�Q@!2�B+a��i���9Y�1t�^������1�o����X�X�t���0U,�)�7&)����Zh;*Mt�:v^h>��ƬVL@G�ےu��8M�o�s�Ɨ���u��F�#=�>D@x8�3�?f��(uL����@;�f,�[G� �}�(^�<U���W�;�T����FY�8��u͎�o6���.�N=3�4��v�mN�~��^Q��7/6#.~���P�L7t�b���Y<|;��F.�/*vrs6�d'v�uff�-r4�P�̓%�
x�9�g�ѕA�Y�H6�,��qF���G����EN/�Lnv胃��A��R!W���m`s���[�:uo( o�T8���8V�Ccj�8���j"ޫi��{�5��+��>��wy��q,d�Z���׋���2��$��}^���y��~�4�g��3�g:�k�������:̆�z�s�h�C�&O{n��غ�<)����ҙ=)_NWr��7-�<�@��l��#���,)AP���`0.�w�'9<�͸@1�t��o\��7�Qv�7�m�a�ͰD��0ˏ���(�i��6++�v
Uf����4T�ٙ�)��>�psߕ���xʩs���]ƥ�7i�R�^J0�t�Y���K�$�B8O��	z��fƩgVs�F_Q�v�&�ڒ�K��J̬W<m�9�t��͕h��\(i�+|U����'�m�E|+�y_��'�3~�;�����]wD�����C~8釞�Yܷ5�:�ϻ9r��e�־D�*�;��8��u7�����Z���+j
�eܤ^ggΞ�˩�Sw+�r��h�ۮ���9-)k��}ڹ!{}��.T�x/�l�Pn}q�G�έ��x{��Ry���U����~�Q"�*
"�ߥ;+>��h^���Lmv��E�}�ͮ*U����(����|U�l�p�`��� ԩf*P�
���<1�����6t�l+��T�/|5�42خ��f��Θ�=L~*Y�m�'	4���(M������޻�E=b%��{K�n�{���_}t���Y�=R��Ġ�3I�F/E��݋��^􃌉˯Ub��Vq���vY�Mp�����n�&g�j��=M
�V���:��_��ޚ�l�f{��U�bzAC ���f��v��^�0=W��
�x��EsHz`�Թ9�����7[O"|���Q#q��.��^ �	x;[�V��l�����cӷ���k�ˮ�V7Sޜ��{�<(�n�cB~*�m��Dgi��Z�������0��5U��K�`[,��w�P�j�[Ү4��]�8N�ۖ���V�\�t���z���K��QbaTW�6��x�Q7��x��vW
��Q�!�LH�W�������]���r���=�E�w69���)�����d���f�.�ùW�#�,o��Q��;h۶W�v��}Z��ƺ��Y]-|�*�
���{���!��]d�������UJ��M���{N�(�#�q��6��`��CQ�}	��Qͮ�4��g >#(;�
nc��Q�J�[.�͂fN�<��s��x�?�k+���Nl��</>�;ثw;����'s�BV$C�gH��N�f��e%r}7���76�6أ 1��[�ĒV�
λ��2�02chk�Cv]�=��uJ��GE�_
�"�5�E�7Ҕ�D�v;Ffr�k����9#.���Y�4A������
ed����1�f"�b�0Wjq1��ŭ�[��[��=�f�� ƛ�|��|qD�|�ȃ���%_[���o�^q����wC8D+B]U��ِ2���ǽԲ�}r����
��X)]��={�L�9�.y�}B�sU�{h�5�;udZ����WG�T�0g�ВPmӣH����e��Fm�Y����Ob����T���\r�-�if�7ʭi�.e�=�ږ�#̺�t�{QU���[������ P@��4�׺�{i���e�B�]��h��b�'XQ7�d�+%��E&<�S-l&�m��M�u�x4� �7��΀oxv_�uS;X����V(���T��j�wO�us�.�[�)�N�
��*!tՋ����[��|���У�Ԩ0��+oF�Y�C��p!e�Ŏ�
x��UM�f5 T�#dd�ZWK�Ö�s)r��rf�c�](�uu��[�M� '2��.
	۲^eZ
��W�Р��7�#��2TR��!A`6�Qw�B��Kx�584>��T]Ig��A���oΝ�� �G)��ϕ�Rշ�2P.һ>x���f
X�۬�AYgj^�*wApeo��3{��4[�wYI�n7P�e"*�k���ΕJx]_�(]�1`�3��͆\���R�W,Q��X�<z����
�H����U�E�]CV��ͬ���Ǐ��ܷV�x���[v�]�.�����t�_'��G3.���d�O�x��|\���1��.�t�b@1�,@j��ν֠��1#,�[�OwE�v��K���Wk/XJ��h#e�k��u[��h.J�;�mN5wԤ�u,�7Z�0Jcb�j㫘ԕw���+�pWԢ��H���`���:{��t��e�n�ݿ�W���:-زF�Σ�Ճ1�ף��7���P����5�N�V�d��Q`�@:�C-��	"�nu�
�&���#0�Σ�]�z�Y[a���E�sw+>�ɭu4��Fwd�#Zbe��]�wuty��Az;E�'t�۱5��z��=M7:e:�
c����G�r����ܼK�@ ���A�(**
(
	��S,��Җ,EmPTA����U���VX("!Z"��(��"�*�Q�(��P���b�����*���h�QTīl�V*�����b�jQeb�Q�����VX�m�PE�bUPEEX����Q-������� ��DYm�XT)Z"4nZ���-�Q���Z��ZT���Z���mX*(�+E[d�[KAb,-��j�����P�QeB���,F�R��
9h*�"��ZUTDJ��1b��DUIAcLeb�)EUb,jQ%�F�(���e-�������������%�+Q��1�Զ�������,j�ʪ*.4PTb�Ѣ)���Q"(�"����)m�33*Ѩ��*Ŕ�6���YDm3%�UUU����Ie��"1QUX�Z�����:*䆹"��s���4�*��{9��.�r]vAJPz��ti`���Se�n�LIZ�.LiW����!�O�EU�=��Mk{Om���	��B�pȱ�Ǹ��Z�`�7���ﱿ.�a��V
��"p���2�E��"���L��J�E�B6��E�U�ٜ��.���q���~�xN��N��/��¡,�H�ɔv�d�0��Z ;R)g_����S�����;K�g��/]t��w�[]�2�%�.}�+��T�}�K�:�����0J�4X���33�����;Q2_�ع&�l=�j-y��0U�N"��6�h4��;�C�7�4��J�	X�m6�wsb8�3�
ؖÂ.^����߯�s���*>!���!еGL��֛���ǹ��3�M�}G��_Zf	���O�s(ۋnh�6):�"�*F+Z�;�B���z<M���"���:י^M�*˳���vY�Dϱ�Ȩ�n�n�Q�G��.��_m�֏TpZ�<<)�Դ�S\5SJ�z_�F����1��nV��]��z���k]J>��C��\<_.��'�i1]d6(o_��YkG��'�}�S��I~�[���>�ޕ�y����s�
�X>㴯_�},���b���Ѱr*�,���-��}՟m
{�0���V�.Z��������|��h�)��ޮ�����zx�g9x����s��Q+z�[@m�z�MCK�r���у:��N�[�Ҏ�(�ˉ8mie��-l�a*z`Xm����g���e����a��oO(�MlYZ�~�:�f�nqʰ��A��hھ����%��'�����E��{=�K��w]�Ῑ�`�ϣlc���*5]�}��M ��٨`�P�6g���lZ�s��בp���:Uj/N��p�7�7)������#OGgj�����_��(�B��R>/���^ٱ�vr4�!7�~t�Έ�p��Z�`Rʭ��.Щ�����͋φN]�9m�1'g=��o��������m��b��%���n���;�2�~���(��~�4�<��9��E�����=�d�5L�eb��h�3n'�	��@�Wk������/�R6'��<(�1J���D��>��DSsSx�1z�҃k��2�_[m�m�o��y�w`��^���T��9�3����i:���*�&x][�I���P�ަ�}rX@�B�	t@�q��|.V�ើ��r��M�\�5
i��ٕ�i�&V��N;  Y!}^�w�k{����'�t��c�G�TG�4�Ğҭ��]�Q:�h�,�ϱu����ג�2tH[���Cu���F�v;��\{7"㗢�rN�:�	�f�j��\�L�#b%*��t�v�4�ٵ�͛��+R%|�D}|b������G��� ���K	T|苀�E���E�+cq��T�-��YGx�]��Uf-�B"B#h���y:�3��)�WPx}�ނ(�hυ�y��rp�� ���D�OK���O��p▁�r��"�j ԘjB�������<sb��ږ\�Fj�H��O��G����*�+%u(w 9`���ǂW�\s�l,E[-v\�xܹچ���r�G�V����1�x�z�P��s���8���,-�F��˽z�2$�^jᗶ�-w��i��^��v��n�\��Wf��ļ���Ưw�o����F��㓪ȵ+و�9����-��:�U���.5sU�&�s��*�+�c�*��z�xk�槒� ��
w�����	h��0��KC����ڽ���i�ս|��/ٳǙ��E�U��C*�o��+��/j
��;�È�E�CO�|�wN�Rf��|�^g{���2���]qVm���q�[�ڛʡ�J�����TsB*څ.��KKng/��"��"�YTnX��P8i��a��-.��RZ깹�t��'�ĩp�ߡ�p�x��Y����|WF�a��qW	�6py�e��Dc��ӓ�|���:g:�/�:ڽ)�/j�	��ۃ����a1���99ׅ�\Ń���\l(Qױ�8�j�l�Kb�����:��`�d�v��mn޵tle�α"t��8!��yK���3�WK����>��g:�C����/���
b�E�gL ����z �OYF�:o�eu�G^��Cޮ��8���$��r��D��4.bVel�~<�˃�Ϩi.���3��X0�c(v'��%\D������yǭK
1��cwbM�r�$J��5�O�������XW���j㚀˺��W��%��v�d�Z/���`�r\pK}���I� ה8��*���(�I�k2�s��+%f-���aӜ3{,�@;��C5PΘ��`�*Y�m�8I�*]����-!�xuf7=��#*:�Ja�ZZq/�x�+j��UY��E�A�w(1���X���<��{��=�������\�+l��tv����-��?���`W���3��ڿf��5ީ�弦���sA�;�l ����:�`�9�;|0Z����O�p-mz�A˨�We�7��y���.�l�I�v�n:}�*'��.������O�ٛyȣo�M�K�^����ܢ�0���qK�.�f�pⶥ��OG8:A,x^��7	md뷽Ս<���hb1\�J®:y""��k%A����޾��0�����&���o������<%��bٕ��u��1��~�����8Z������g(��X�w9P�x!^<Y'���U����� }<{*p8�E����UشTf�ث�W��$s{�rfK�����[[A�/3W���Ib��,�l�ӋT���M�K�v�J��>�.��N]VNP��npʕtЧL7��D_��a��Α�y�|`țzPNq|����=;�j�_��xxZ9�HB�Ѥ)�k��+]��fSE�)��|w��/����%�:�Ev�����T�ם	�h�L��2�؈#��\h+��ʷ(̭	)�R�fm�5kgr���\�B7�Q��؍�p�f�	@җH�`2ΛS(�b͜�5�)ݽ%M��ׁ�g�zQ�&��tNױsͨd9���C)�����.��cTh�B�٘��ny-P��U��4�^il6'˗��=���'eʞ�nD2��ܕZH�kZ�֢����Q�L$q��xM'�a��,�U���Q�lRu�GE���:�s5��Ϯ.��M����{	9�{���@U�r��������bnKz9z��ZF���1'D�n5�6k�gu�����ő��5ѣ�� JtzX%c�����a���[��<`v�G�9�����,9�FŸm�d�E�5e���N�_7v�H^x�m����8�>%|)��O
��ߝ^c��[���}����Ҝ���bv��Cۊ�-��/��3�W�A��-&��3ײ�f�V�=�f,��8�o!uH[m���;�b"�4%6f,�)E�3K�?v�±�t�"�e� �;ֻ�>|ۗ�u����"�l�LH���ޛ&|�ȺA�
��,���=���A;�{���^������}]��W�p�ŀ��!mQ��0�̩}a�����[����5SZӴ+s'2h�1�H=}#,L�3f��%�����y�V��0���]:"�\������@�Ep�~�)��t�G�0U�:�����se��R9����Č}����N�x�K�|��U8K�~�Ag���0�ksԫC�P����]/ge�F:>��y_o�dj�i/�(�����J��i���Õ4tX�G����g�wS	zȸsx����=�$U�C�ø�
(�u���R���C���
��n�n��?}On�$U��{+�{��y�agB�R���#�ěy��h�H�Ѻ柼��o�=�ƶ���K�(��[��ݍ!�٭���;h��#��䵐-@�M����u��I�	S\�C.��Y]�H�'BE:�`h7�l�����k�X���I�
�[��8����^�ـL1�V�;��!0R�*�����a�;)j�w���B�����*Q�1B��(��ֶ(�l�}+J�{��6j�D����w/�8�>�ު��K=�l�auS[�>��x����vL�V�<�7^o �0���4<���/�����2%�1^RAF� T��g�/YsUp_M�8[>�QyRڍ�1K��r����s5>�׽�qɣ#�:f&!�Н��R �z9P^u�/k��]�=C�����)�b����L��U`�j^ċ�3C,�B/a�Uq�+Ҧ��jք���8:�*��%���4�[w���w�:�]q�Av�"�j�_�.�ұ��e׏��|��]�m�mg�߳C��e�qz"J��]
�$X&���n^a�F�����v�s��#������;x��V������z��IR;i�QE��!�N�;��v��X��
�+�|�����^�b�{ZzB�hePdVmR�1��bⲮ5^�f�hv�O�9�����<�j�hүhOn^�t�h֚n�#�b��Ϋ�]&�wQ���B�0l%q��O�2�RY�.�����y��y
���ܴ�s��9�Ȕ+�9f�U�u��E:I�DD�Qq�N�{*i��l���.J&���%�꓃���������B�{f#�eT���-����:yy��n����@������n(U(�ޭ�]��i���^|*�<�h�+eN��q�p��y��Y����?/i�C�t4�p����Kh��eꑻS�oz����1�qJs&����Ԣ��S�������cE��n	��_�v�w��{���v��n�Ts���O���޶�
7�*6�Ⱦ�}nTB7�q��l�Zu�b�ߖ��N�����,���;n�
F�w=Nhu�+�p#�s�$��F��zv�9���H��y#>2�\�����p�]��OgQ�zl���٫�lHu++�l���bZy*�Q��V:���$Zr2���kY��񃪶U�p\(i�)����Q�r�]�dn����&x{�;�V!�6c�X�ؓj�MċRC~�s�r��|�����x�If�e��:�gզp��y�f\i�y�,�6#|)K"�J�b�	��F��DTY�B���6����:��N�8�}���D{t�a��6��>�lW�O��x�7&N�\v��W|�s%ц��}�ھ�ku��5�r�}��Ҥ�����§\�>J���t�:��?V�`����]���t�-������lz�c8g��.
_t|j�#A��@�K8��&ge�>����o�
�p.x")v^zVm!��&*�t��|�����N�*|l}�t��%!�a*l3-w.�2g!zz��dx��v�[x�<1?���@�\�f�6���0Dt�ǫ�\��9�z�}L�QA�+%���n}���b�u�k��s�%[���nxh�}lj1���s[;T��~���)_k�+��I��ضe{B"�i~?^��p��v��RSl�ǵ�������م�N�C+k�Y&z8��j��%oyeiё�^<(���"nW{�'k7��.�;9���ܹC7��O�\��������X���LH�K��c-.�V5��7�Yc#�����1��7)���Q�,�wH��gd�MwX4��I�evn��"�ܝ��X�Uy��z+_��4��4
fV*Q�Q�+{M�f��I}�6�a��������q�o�S�!b]A�hm��]�@�.��&�Zt{V6��gT��[6�َ\�9��z�v�3!;qX�+��Wj��=����<s�WO��zxS��W$s릕��)���o��A�T`3��ĵb�ј&x�͚D.���J�A��lN���OV_�5���:�y¶M��<g{�x��ӛ��#9di�s��B����s,�zdlF����H�
�<Th�t����N�#7Щ�$Ϲoe��U��oƠZz�Q;���C!�X�X�!P�p<�pfOm�FU���i;* ��_��t�-�������|/���9N ���31.�qq�u��L\h��G�Y8yh�>���S\�{�Hlz��>�����=��\�6�������$:��:`<����ꅑv�"��~ �<�4n5{9��=,��M̸�_�U`!�f4*f&U�YQ{Ii6�������~*�R��3�tS�V����[��1����~)�{�XE���B]a�C�����t�,�@��<kt��(����{��e������3U�r� W9WV�����;:l��5�0���|����]�T��v�4�.�ӆ��8͉,o�p���Sα!Q�?`5+ݏ1��r ��r �U*����WW�}�d��4���t0�n7�6h�orQq~
��]N��:f��S˾����ϻPSwT�6D��e�*��i���� ��ҭ��˂q�
�v�|6��i>5�a���7�Y�"�����Z��D�[e��\t��*�wi�n��`���zNvf^łxH�s}c�rT�k6-�[c���]-v��\�x:�
�,�_��3s�ͫ"�	�t'5�]*QQvtT��r��ܒ���LÅ]����:oV�-��C6�9C �i
а-z�����K�Xs���N���eA�:j�Q�,���f�7h�&$ȝnޗ�vч]��$Z� ^g P&��
�22+�B�,����hC���D�t6i*Q��.���wN�f򺦰~v�s4	$�cx������w�n@A��E�9Y\��ZB��X���
b�JY��`�衒_�����>�+�*����֊+MM�!pa����v�I
[4OuN�/\�$����j�r�`����Wqyc���-W&t��V,�uw����k�fԫ�F��'���r�v��{a�kV���u���w+U�$]��9�	ԑHճ�eg�:T�.��+!�/��^��bG�1�لt}qa��גX�.�#K�Λ�뵠��tq���P�I]IR�wh����#8�wX��J*�A�e�g��������v�W�cޏO2�92j5{yB˭V;/;���s�bي���{N�I�Z���L�iꡮ��v�WV�����El�Z|�V˗"�����s���S���vJ+��1�T
yj��S�e�|S�^��#�n�kgt�2:���l ��k�[w�4�m��d�b_����C&��&@p�1ـ�RF��vb"�tM�4�DҴ���
�m=���+P'�e�����/�*�t��%��4��[�n�L���Y��.-K]Xf��-�-�PX�H��)YG)T`Ѥ�Q`�Z>wD�1�Y±�H�Wv��CQ�:uh�r�Uta�NU����a��Ѻ�S��[��ΰa��6%�Ě.�e,UfU��-�����D�%���DM{v������NF&밈;�1il����Q�m���0g|8�x>�$r�t�^R�hA�ڭz	���H���l`�,��Cd`�H���e���Μ��{�<�bpǑ��p,ͽ��N��J�n��a�/�]�D�<��o�HX�]$�v��:���e��7\�;�m���R�}(���˃�A��p�XC�zk�\�T���y
���2ȳ��Q��]O36�s�W�5M��V8��e�6����4��Ć�5+�3����P��Y�Ŭ*(t�쾃H. ����H���Ԯ�VJ%�.�&�5ٚ�d#w1F0ftv�ZZ�R����x��hY��*I�
Kg*糢Hf�ʹ[�Ywy7��ŧwso�1���{�ֵ<kx*(������^=c��nbHN���6�L�<2R�3�o\h��ܾWWwq�DY+**�ՎZ ��ĭq�_.cuh"��Z������DdV* ��:q��ETQ4���AQFڢ���*,bT��]%V���*��lEX�X���6��5j�QEƦ��*UEX���:c��-�������Kn��A`QTAQ5j��TETTb֕(�Q�%��U+b"�ֲ�h�UTX(VֱY��T�q�,���U��V��Lj��2�EEe��U��ƵEDF7�mbV����c�*�kH��[.2���*2)�.�*�1�,EQ�,�j)���"�lU�X����ĕL�TEQ�2Ҋ��r��(0�Eb�Ab �Ԡ��QQGIE� ���"������PX�Z�#��9h��"�1TKB�QWV���*�D]R�*�l,c�	�n֜��y��C�7{!��9�����Kw�t�ϱF2��iiMj�p���v�6n���d�ʾ�'M
��+����f�$������w�8&gp�V����/PuW��]%����j�P��Ž�Ѯչ�h��Y�r����^3^�k���^5��YHeW��K6�\}tUj�K����=��<�D����	�Z�u���������	�Ja����%��7�I�rGש+`V����!=/�&<׬�N��:!!�t3dK����΋���-���ԎĠRX�|�Y�f�c�X�/�0	�"��Ci+�Y,���rɥ�v2��K;[�ʼШs+NP�����%��)���Z �kϬ�rͽ��D50�h7s9E��ծm+�T�V`��0������R����}+�|�O��1y}2oK&<��K{2<��蕍g�������!C�ڂC(�%�c�#`um#u6P����E���{1������_g��s3p��p*���.�/ τ�8K\���\/Q�����	����R�}�����ܩĩd+�X7��H�,��,7�>Ba���O��Z>�)����=�^H�{O��R��	}����37`��GI�n�^� e6��WT \��o_�@����O&Z���4����9iN_ыo�f	*s	i�a���xө��
�c����XWdn�n	x���:��1@��йr�7�۹y�p=gA��>�xx*S�>È��G�)�C�a�0�8��S<��[�b3ӥdXs�������
�6Y��%
$��^*Y$Ph��ˠ�Yv�ڇ�k��2$^^j��X�y�R��U����3��o�o��4��`�]Ƅ�{���7�}w�Յ�~�!�Z=�e���'��xS��>�~>���m�:/9����p�:F~��qGuNlpq�M��S���H��X�̿������*ߩ�6+�G=��kGv1�r���N#P-C�w�5<� ����?JаW��@;7�3�'�D�p�Lf%\���V^K���D_��E�U�d2�f�z�wT�ۤ����x_�i��L�Nr�o�Ex�|�M��q�=�b��.�T+��Ӷn�:�l��	v_o�Q7]�m��:�o��e��EaՏP�F��n�R��S�D#�-�8f����:�E���1:eL�����g�<=�� ]O0*5��V���əK���3�v5T�pں.��Ko�g.� ^e�E�]�x�3g�5Sf������`�r>9��n�e�H�t�e�P_2v�Wt��4�3�qX���������^6�z���C���ؕ;U3������k͝����H"Z��܊��Θ$�6&1��%
����9Y�ZO7c���;ܷn��?o'x�VS�2�#�tAf�`�dt��M��r�#�4��
�XO3��i�^5���e3OgOY�Yd��i���]>�6QDч���lVЪo���س�q��7��A0��-�m��w�c�C�n���)�"��=KIn�/�j�����ǝ�0���<
Q��V:Q�Y�g�<�.����f�E�RȀhK�`N�M��Y&�w4��a���(L�Y���j�E��Jإ0C4Y�'����g�SM�c��zÓ��4�f�`��d�Y��C�]���M��O�S'�!G��P�}�D����1�tÝ�;վO݂��_O�4+�:�z���x:��9)�����e��Y�^K%k���j��s�3��Z՜}Zh3J�Aä�b��X}p`�,�k����g�6�)88�༔i��8_��Uj��2��T�9NW,��eu�̯hD[���
�~���Y��/Y;y�lBc��(������62���f�,^�I�tYuڪ���{��4���"3��,L��6o��W�«�<p�<�=C�G[[�is~Y^9�e�HW��� �eҶ�Ux�4�ۗ�	6�6���;�msG^��1G�s�ɧ��	�W�'��sbbS,_}Ӻ`�z�ِ�WYpt3�֨N[���r��#���_.��+:�W����gLCl���%���!��"u�2�ϩdqS�Uz��T."�e˾7��ܥ�m��khM4��d�%YXp:�.PC��l�����f��v�Q�S�k��Ry��%��j�~��<pQҥ�tR���h}�_�ω�F�y�We�RzWc�׼ĽL@S���݉�jV��<�ᜑR�拙#���{��a��ڷ��ՙ(��-^�&+\��eT���(�U�+��J��BP4��;���8�4��[��{^���]��%��Sh�(�>uF�:�ު'k��=�8��ٗC�t�
qwN�gV�F�.�ȋ�<nʖh_M��g�4ܩy�B�f�7w������)���C������$:�H��0.{]��,/��p�d40��Ǔ��ʳ�0������(��W�F`w�3�7�Ȓ�(�wS���協F�;L���h�BT�G�k8�O�rЗ,�2֥\:��q�bU3*�B6�Y���V�n�ᨹ����7��s��q�����d�:��'�fSO�qg'%�HR�6�{33�oxq����F�Wd�k1ͻ�Ü`U��m�'�`�1W]4r��a1T��n�}��cY�Zp^�+�"%N��x�B��j;϶�L|^G��/����e���ץż�&�^e��o�2,��̫')J�y�~wB{�����$���tv���[��F[�O/U}����ɇ�s�6%��	�2s�u~o'���s�őt9^z�Ʈ٬�c<�_��9�'�zQJ.#�p�6���4P����-I-t�.�Y�>�plnu�����WA:Ot��-B��"�x��'�\i�x���t7��y�g�d�������d�E���{������.�Ӊ��? D��޼���Y޺���43e
�{üb��㓨�3�ޚ
��o���d�^�x��֥��xϸ��gÁxP�5Bء��q3�9�{��=��u:���0-0���BjgP���ɟv{�87��>\���`�"���3��֚�z��J�`R϶�>���w��b�qL�Ӂ�d2.C���+�#�]����m+7y�Oo�%�h��D�]��-��]u��U�ǦuK]��m%y|��9���<��Ѕw�k]^Е�i��r�g�cf,�<+5�Ҷ���k�,9^�8s9�v��������H,l�Bŷr�h��ڞsr]��Z]��-5�q�����u:r�۾�N �/�s����{8l_��A5Z�3�4�_c��)ں�L��]��F���x�5{����o51/��5Ga��RQ�.�+����4q�{�G��>���='�Q�
*�$�K�zѤlt[�eE�o�ϯN^)�y=z��כ�}�l�uiՙ�cq���&��&���c>��y�L�A5�T�� k��/�pe����N�d��FwI���aR��>��|]O	�K�n�+��;�b�|��ɨ\c�;��n9����=,����Qw�S0hJH�l4]ɩͅ�0+��x���l���R�<&���V ��-�)��\��S����(�w��K�J��Z|�3��u�8"�<sb�9�O�j�X6Y�7L�B��.zC�W,����XN�n��[�O�����7��w�T��g&;6n����:.���,J�`:Y����q���F���Y=�@�W��Uw\!ub��nZ�/��L�D�ʤݨs� �-�*��"7��O�Ƽ�g���>�xp�sȃЃ{�ٖ�矆[4=[�l53�kB���p��d��4�l+����&_	����� �]h��g��V��00y� �'m��غ��ӯY��F8i���̆IXM>c�/a�}�jt�)@�:^dn��4k��d��f���$wAG*rb��UKs��:�����|���W��L��.t�K�����Br=�gFHbSiM���0�C��6\�pt9A�V�K8+�[y�h��J57ԁ��I��#�(�S\�s�Y/:F�JY�;/F҂&�[��ʾ�ÿ#��7��aͥ��<�OO�x8��t�)T�\�m��ĥD��Mx��T,5�=�G���)X�W�*��슶'�Z����X��hз(����}=ɇ��x�'Խ�j�,�`��:���U��Nht)�s��%��[�Y���g���󥂘����x�|��x����� �@�x*��cp�4�������w{{s�:�|�敄�N�MΪV�d���sJv�^Sl���ȶ'b(˄r=S������v2`�[~�g�~�3��Cbz}0���p(n�I�N]ċ�AD7�f^�9w�ܕ��mER���!��V����%^�X�k�r���O��hR�D��n���m�we�@��<�+�����ɬ�^0+S'*q�}�`�U���z��`]�RB��.X�Â�j�-u7^�P������JC��dhˑJ/�aǼ.9��C���N�o���nm�0�i�ui;��dWv������o����ݾ��j<���� R5\/I�}�K݂���g�蒨/6�[,!�nS�/���OK��:�ܩ���{��#լ�'�j�GO:��Q��ޮ�#3*����6�����<X.qa��r����cWA�j�Ϩ綦��{��AU�ɘ1�i@�-:ȍ'�:��`�xL�]����J;4��-���9x�k;��]:�s�+�a.���C�*�mP��9��at>2��g�6�X������&�5��Ʈ�KW5k�SZ=X^+�P�F�}��i��'�N��i#��aSfuzLz:��8}A���X��~Jks�m=���[�� =CZn�l���h-�u�ɬLɗ��[$B��K�B�^�
�S���r���%}����4U�샋C�����$�v��g[�������P+:�FLa� my��b�^�,�$:��7���嬙����&ts��޺ብ�6)������`�����G�g�� q�S0:�tb��5u��7�5w_IsS�Ɉfw��0T���ee�W��)]�Vt��!:%4�d4�N݇�r��\����bTw9�2>Gk�]L��bf&
34�i9��A�n�v���������s���4ׇ�^T��O�cGJka�5��vVs����5�+R�>�B����!3��;a�����ث!�Ӝƭ����!�+	�뼧 }|�=����{�A,ֱ�MP���Q��m������PӬ��sj�wR��ozdw%n;�<o4S7q�pw%��t��H�`O��WХ��t݀T�^��!^f+<�(?<�朒v��9k����-��n(�b�.�ʣ�#Ȇ-zC�r�G�0��<�H<�T�p�J�5xe�R�.�CȔ"�fgL9ƶ�T0V�=���>|�*B����^�����u��Ǯ��ʱ�Mu[^s���VD���DP�j�uX���+y&()�u^5O��m�%0�����ۼ�̝������[��3T����e:�l6g�	E�2%a�lG	���&�.na��ؚ��igyv���Y|%��ܴs����2�q$^�b�XR���6N}�)��ח�f�yjE�u��\ϯ Z�8-͸��4P�����L�+��3m�F�grk��f%�z��Wm����^/	�8)d�W
q9�E�\"⼩
���b��;e�14d�b�����p��}��/kΜ(��
������t*׳�r�E������p��vq o�6�d���]y�J+yW�æ�*���S��[8�ؗ^�T�X�H�]]��Ts̊N���z�|>\f�����V�4����[m.N��{*zh�K��z!��K��i�4�K�U��oK�@�}�y���[��iiZ3���Վ��ک�v�)�o	=�P�VP".oh]Ԃ��a�ˤO�_Vu]#��z�s0�1��,4}S���7��xgӫOa�Á�A�e����c��*!F����N�/��k��H��h��^9��-�+g��]9��Ey�t6L:��FI��~��i�=�t�}n����d�W]x1��1Uu���E���_v+�t�z��I9r�VZ����s�<��_G��M\�H�qj��l�K�,��������qn_���
��,�W��'�ƟK�P�e���4�R7=6��:�=6�c�y��~������[��sd�غF����+ ��@�s��cxTJ��V'!�U�byd�Gr,�5.F���4�M�I��T�8G��] ���԰��|+-�(�*j��^Ν��\�ag��^�3��7�N�DP�,�������,��,U2�kW5h�=�
���g6�hm�����k�F�p����mN,8�%1a�*E�A9�ra�C'<��)7w���ޢNRPx�)���^�|S�8�x?YE��*�^��Wρ��r�$�u���#M��+�z��w��� �F��ኤ���fw���R9��5-�M
��ab���*_w-���hsA�E���2�Q�x����5�mu0�	�;�Х�o��0p����)m�mM���s����S�����ɫM;Ҕ��-�r��Vt/Y� ��gv:��Ap1f���0�t]����46��i��˝ձ�5�E'-�����8(����~??��I�x�p�)�-Ǌ� �+���nߖ�
K�"��|�J��'|���>���,�W�uc���a=���e���ۺ*p9Y�W��g7!�h4.�j���B�]�l�+ee��l����B
pԬ��M��t��}���oeb�:���:+��4�iK�z�\ĩ�t:�wz����"Oj	Os��nX�6���.�������"m�N��$�H^�]&���A���՗.�q��⻐�۹�v�����!�(��<5���9}A�wۘ)G���R�b���Aݭ-#6�q��s2�=��֐zt$�m��������Q⿹�;݃�8A5�ڧbPKi$��i�L
D���<K��
�٠mkes��ÇE���C��,�ϕ�R�uȢse<W�nJ�|)qu*7��ۜ^,�$�t3�Z-J������'�k-�u�Vd�+�R�:�ԳV@��Η1�!G+��z�sY�T��޹y\�B��4'/��C`��Ib����L����jB�g��Zt���a�wGz�y/2(�]��ĚN��cv��n텁У�GBO*ݥu�F�O,�eVWeXv,`�K7�*˺u��x�XJ�V�A���KosKa#wm��1d]S�h+ںH:60�t��hᠭ�.��U0ٰ��ݟ+���|�O3*��a�4P,�_M+,�V�f���$2�Y���݉�7*&B7��CI��"i"�iyb�����(�
�f2�&۶Q�
�&��܁ Ӎ jk��1틥��'J8�Euxi��D������nT�s��vP�8�e��!(^2���G�'n��]f^��sPW\{z�f]	@�̢%�h�Mb5�y�2։�Z�h�ō�Z�s�stm�WAzz�����*�D�t�kH�U��<�X@����S�y���r��[)+
���Ἤ�Y�#�y-5|n1͵�M/V��Ч�{��`)��������l7�����;[b��SzP5Ѭ�ϻ���<��F��Y��ӆ��W��ƃن�ta�L5I'ܔ��/fC�+(��1�/nVʌ�<�|Ag�:uo���toX��+p��XAu��v��X�Ȧm�6�V���w��oF�7tF���̴4���r�Jh'�oS.���M���wm��h*�1e�ne�b�E昶UaP�#���TEUTci`�Y�TAY����*1T����("��"�j�`�2؋��H�:J
�*��M!M6,Em*��"�
"#���(�F��X�

��+�E���Y[FK��a�2��"��WƱGV�K5lu[AQ��T+EETU�����E��,�VڬPTATkb*�Fe�+2��.�b�,Q4�1��\�a�*q� �UI��2�Q�R�5p�1̍����e��Z�eՅ�J*[Fڋ`�[�eJ�ԵB��F"����Z5�)J�V��m�řj�LM!���\6�KiU-(T�ea��WY�LF�je���mUZڔ�v�Õ9���Q=y�c�:�o3��d������S���▄Z����J�of����g�!,�+��$�`Hs����wu�Kӷ��8f`�z���0U��K�� J�90�i�%�����rf�v�$�k�����>�{�l#�ёfh�ʂ0����Y�`V:`ePd\�uIȻ\P�4=}I2�NҩMl �Ys��Wl����D��8�,eS���F����D�u�%
v;�6]u�{�7��7�c� �w\p�͋Z���r0����;�El���wxb�}=ա��Gn�tɭ�,Z�f�$��ґ���;�*�݅�m66�kˬ�3�\Q�J�6ݩL|Y��2e�p{���Ҟ?+�4�>�My<|3+WWe�Z��ej0Z;�mB/���شU�B�f��#���u,�j�<%g���/ �/�`L���K�{�W�WR�Y��+��(�`���Tx@�:U�=s�4}�<�j�nf2<���{���t=�ce��7�����\~8�R���J�T�6"��vA�}ѳs�֮���~�Wcp
��7�Y՞�d��TE7=q=�)�45�Y�c�/t�(�L�uH�`9]R�}�+�E�ܲHQ��j�ܐؘ0�c+9���X�:Usu��J�z/Z���}���m�0bH�k�vbZ���n�6���R��\���[���AB��C�����Vu��^JΨ��r����.]�CЏ2�p�[��(&��`�͚�hz���C�[}���E���@k����~.��yy��C�j>����/���P\)�N�h�7���j�jU{���S�s�$��g��ٹ=��/��x��1�7��J�'�X�k�rL���o����j��=���iea�᤟{��ap��V�^�U��K��O�Ø�Dh�|r�σg��$쁁����?~̚Ҿ�U��p��dJ��G���RӉq�+��O
uViqir�繭e�}'Z�7�d��(A�3G��*������J'!�֏/Gs"�Dp�z�l,�vZ�S��ʃ�o^����@�")��o�8`ˋ!��H;��7V�C;��塆�#��V]�S;q,F�aWO���V*�w�^����#�Qu�F!��o��~�pX��Ƚʭ:s���f�l����d��.�5M
��y����yQ��׳��9綬��׫5h��JY�#�*#5-ޜ��>��Y�Rˋ����=V+�9�a=O�����p��j��^%>�,�8j��d�"(!�*���'՚�NmE2��/h��JXP�'��?$6��xE6��˫i Sh_a͊�����j��R�Vwߣf_�j�z�R������d��N�S����7�U��r��z�(L���'�I��5Zm�������-)¼�WtR�#�0Q�禰D#=HO�[�pr��V�j�od�#OD_C6ԆYaҦl27"m�hͻ��t%R��Jv\�ڭ��k����X�ݺ�>�,P��n\�<5	��l;��VddD�L̬Kd�J^Jq�jk7*�GP5:q��tլ�����x�^=�� ��M�;L��vr�8f�ȩ��*��y��V�C��\.�،�:hZ�h��3�pE��v�=f�e�(���:��h��ܗ��O\��5uO��c��Lk�I.�gT�/��A³���5������9��M,w�%>���yp9^T�y�:�N�XmJgE����R��׸���' ��C�d����8|g�2���n�C��BqfeK0�;7爣��q+62v��BmzO=Q��U��;��G�f�L��b�XN���1��u1F��ژͨK�m3[��_l@ی�g�0z�(Pr�<�I2�R�Dr������O��R�p�e�Y���Z�{`��F���En?-[��ѩAA^z����q�'N5s�+�m,�)��a�J�20;�KB���ԱQ�oB��/���k����i~=�ӎx��E��0�`S�NuJ�-eb��S5��o �bg��fyy:Y	�}7n�$T�`�r�D�p���<���/c,R�\�ڢ&�7��.yd��X㻜���Ƀ&^�^�"OyU{�4kœ�,ߦ=�T.�In+6h�67%�{N���ol}�RO7o�1J��[[�X�r�Y0d67�.$��GTˡC��}����gz8�
u�v�P�ܱw3�e;���4W�K��hʋ� Ps��/N��fyćXq��lüĔ�N_P�e��Y�c㢽�|Y�����tמ*�M�vr4�"���oU��
�؜���q���L����q���r���M�3�X�vͅ=]Ѱ�T�Z޻{�������:O��9]J���e5nQ�[���"�8�T>ו3�bega��B���P��[��1ovn�x��wp����wW�8��hu��^�T���H��h��+#v�i�Q��36tYO{|@�U֙�iöcF�9Y�:�~m
d���\��E�<|%����CGk���{Ӹ�7~����VEJ�ʌ���؆Y��Dk�D�f+ÙDs�=�~B��&����Q��Sss���{�#@m��ᇮ'�[�Ě��jB�T��6,��S�[�Z|��ދ�T��z�݌�:�˚��)��uE]n���p&�@V�)f%���>m ��W+\�T�WmVo8]�j�s��S�7SF�d���	s��a1�/�şX�6W���=�jt%��<qVdXr�L2K6�(��5����tҷ�5�����pʊ�l��p���o���P���Kؑ*Y��1�ɦ�|�+𭡡�f @�Ss�ڳ���q�^LPt�`�l��4XoS{ש��ͬР����$���Q�S��`is�:�O�<)E�.�I-��QR�sl�V��V�(h4�J$��3rb�Ԃ֚ARk����Ւ��[(e�=�C����K7��ܓ���%����,�D��ׅ�� ړ��u�Oy[�ٕ�(�K2�yS5r�˖�:q\�D8�|*1� Yr=�N��-uś6h��η/}��XT�w+Ս��Ie��<��t߲�P���	��cX-��k�j.���>�;w�X���[R9����0��W��2k�O[�	ͦIR1�\������٢u	&ZQ
��S�"�po�b�����#���`��h[�U�e�[�,�S�F�$e.��o��Z�ܸ�ܷ��;�Xͬ�{z��TF>�Îs�R�����} Y0�Eb���������
B���"�=�V�Syhgj��Zӂ�l�/�+��S�m<�c��2����Q�xBD�n�5��,��z��|v��9j��`o0ۆ!��8&�6g	S3dμ��2���i73����Om^��n+�6�r�.�o��Q��~����j����5�\����!(����*j�<%t�1����h������5}y�	L�2V�s�R����Q��0Y�T+�Ҩe
�*���-�Ҍ�%��̼�'M>�hW,�Έ���(�RʽtO��=����r3��=eT��]R���f�46�s�;��T0a��N�X*v���u9�+�AD�Ik�ֳ����i�wn�pA�P�6�V��aF�2�`®�;�]�6^�;g�'�[f�{E�yi��]-Bc~s�DJ�0��.������yh�����lt>���ly���qM�B�=U(,�S_18�_I8�60�B>D>��g�!T7ޥ��u�g~VL\CB��.���X�^�i$����6�c�:�4�J�b��4)��
#�'E)oi��f�)X�븢�M�"'���G���ភ�'���N�ߛqZf.C"!]Ad�ݖ��7Nl���:�^�M�S�����lܪ�ؒ�t��u1Rk�8Ȋ�Fl'^�A
�`�㭮�n����[���데�Z;�a7A�+0ܚa�]�v���6���Rf�y�2���t���^}9Y��h��0-�>�2��<����z��erˁ̱m`R^��p�r��t�-��|�%mpީ�5(��	���5�0��Κb,laW�kʽ����>�=:7X<�=%B����7c.*�z����	pvPޱY�����x�yڪçy��/TNg$��ܳ3���Z6ڿ��"�{i��~H�^�y&p��T:��o\ù�鬇�2y���l�y)_?���f����<��*`���OU7�!2��IC�E��*Y�C.�t�ŋ�왪�OU?b.ª�4ߛJ��s��
��t�@U���uo[��QhP�=�,F�����0:/i�oC6����*T̈́�lN'�\����z��-�Q�q;+]��b��$+C��1^z�C�g��BC�<��s>+��xnp;��=��H]���17*�V�۸8yݱ����[�QB���)���Y���ݬ�k�{��[ݖ!@�72K����yAח��t��	U��S�tK!��,�r�����vמ^M��q<�!�ȵ�WI��.���!N���أ5߬1�p@���*�O�7��Q�kV��&o�����&}�!������O6fzᝠP}�Ž+�H���n]��y#���m��N��3g]/`��G���8g�B�M[���V�Q/��4�G}���nŘ��0�m����k��A��c���{��8N)Z�]*������t�i�*Q��Q�ۼ��5c���h��r�9Ve���y$��m�Ҳͦoc�>�C"�M�8!�`6S�3*Y��F�p,�f�����o#<㜌,���r�3���/��S�05�&��b���ރ�'�zQf�L��8@i��Ԧ�]�Wb|v�A[�y�R�L^܌V����X�I���%��*�,�]��_�^;'�'�K������X=)/�.�N6�r=�����%(�z�MӅr�Or����"Xݥ����ٜQ�%�7&�'6Y�1�Τ({���chGE�����_��~�SZ
�f�����R�}��u�i׶��ެ�p�3��|)��F�ں�)�N�q��]������Hr��Ë
��!�/zl�n��Vy7h�b�p$9U�.����,��BZ�������8{�V	��Eyn�R�(P�M���&�;(h�����0Z~�Ϝ�����b�������R�����.�;S`��R�x�)��hyd���h�F���<��J�@�vA���fwg=�N�%�Q:�?S��$6w�8n����?����R�#�,ˈvU�ܒn4�r�K�Q��SɺɁ�ٻͮ]���j�b��h�R�`�u��Q��T\{4["��͗��7:��K�|{z ��xm!L�Oƌ��{A�be6�m҈X QFE�W5PQg�[��~xfߜ�+�J���`�L�[4� 鞈d20)��ٞ��s�Ӧ��T��\��e#8R����λ������ϢǦ�B3�_��WJ�s>�t��7�p�,	o�T�'�����r��my�&{��C�ry�v���p���R�7�5���`Z��{n�mfn4����(�.B4/mZ8*tߥϤr�p9*���N�ȱN���If �RB,��z�.�^]&O��.x�G&(t�3��d�s�k��3��X6�� �wF����&L��`�Q�S^QBƉ�q����u�Z[��6u��7�z��S�7����@��"���q�B���V��	�:kҧ�>�ȵ�iE�DIz<C	[��'����S�,���.�U�Bh]����JWRzi�9-J|��:_Ty�f��B=������%��RK��fM`�r1u�yQa��|Edu؄߮���^H�)Hs��������V)K�+4c��U�x�U�G��ɴ�6����0vҟ2�]Zo]����Ì�w�h�<�@]�b�<��p�-c����q2E�K�p������,��ژ��Գ���ܬt&S����r�E.���l�ENU0oƜ1B���I��4xx`��p��G��EN��6E�zX-wR�f\��0u�4�(��	��c�-����z1wW��PeM
jޢ#r�Ss7٘d�=S)�^?=-�9��/P�> 8l6�R�N�S�ge޻�7�����^�ޕ��T�K���#��m�a�ڴ3�K���]x<�w��g�˚�N�Y�=���R�o��Q��q�SL����N�:�%�B�R����OE���#�uY�ra\�=B�s�rX�}&�k��-/,:��p���]�F�r8 ���mç�"b�<�o;6��֧b�S�/\��tO�'�x�\��/�t� �AP�9w���v.3ɸm;��,���W�f=0�lvz�m͍R�vH�-:n:�z�����R�IZm'�zL���;#ϗC�0:!����2�v%	�n��k+d��ƛ �j��-w&֥۾`��ʄ�\[*����X��O���½-1�͏}Y����.�X�מ�XC����<�ӗ�+)eX�.k�t��5Z�M�����L���8��:ͨ�H�N��0�Z��j�:^�tu\�ڷM�(:�����F_�nByl{�����|��vv�m��Qc�I���}�a�a�	܏N��/�f��ވ��ei���5�>�V)N�=��pfvV��Er�nu�2�D.��Li������dU�X��n)ݔ7#����w�]�ϸ�8�M^Y�0Ζ��ھ�Pb]�"�j�զ��Y�I�Y.�	��Z���+���竱�"�5gz�[���C���mQ�f��vjO��>�6�8m�5�զ��:;t�_+UE��K�Gr�-]�CX^M�	1���;�X+�beV��1Txu����ϖ��@b[�;n����ߓKr�Ж�������qZ�rj������o����y��.�y�뜪��3�fgV@�!l�b���o{�p<��:MǠ��G�:y9T�5{�Z�L��	U݄Ie%N�B����=�j_Fnv��+��`����u'Y� ���q�WLhTj�Ҵ�ð&֩]o	���꠫�n��Or�T�%�|�D�s��}%�V��ɢ�bZYUϖ��N�c�B�l��Xq���YKp�g����ٯ�2�̭o%�<J��N틨��uh��ws�ݚ�u�^!�6� [�q��	ҵ6�Ӊ�u�[�|���a4 f*�� �Mm왙j��/&b F�U��	A����@B5}|u|�J��JOr�������U��t%H��:�;���X�vW��ɔ�Gn����w8��a�-�����A��V	Ԍ�-��e��a����W:�m�8IX��	��{;(,����:�-D�L�����W�+���?^Vq\-��5���r������u�2�4��n�ǲ0����].��NU�υ�aJ���v��v�z���X�꼮�'ӝ�+����=y8��]]��)dIA�]��`y@�52�Zؠ��@o]_u��u2��G'$	�fF.�����D�0���F�-�m뼫�R�@��ˊK\�VQy�p::1���i4�ͬ�.����繸�so�*���}2c�{�́N����C��F��j�O�d��{�,����ܫ7�V]_1`�ۇ�xɎ�	�T9�:'�Q3X�k�%G*_!���Iư.�\ȁ��-��Ep����Ȗ&��K����c.�%��YضEut��_WR��&�lq�V�7&E���-^c�TqTi�	�*"�k�R���:�ən���o�N .�%^���l����Z]q��;�Jb&0z]�]��U_\J��T5�3��)(ހ�8(��P6#<���켫kbﭞӋ��k�4��ṝp:\g�e�붜x���&�}�vR�ޛ۱+U��uK�TL#����;�%��z�%^�~53" �"�@$xlm�ZѩU�L�cUH��-�((��R�fZ1T�KZ
P����V�c
2UjQTE���ĵ���Z��TEe�*T�#M%m�����V�,�	���-�����
��+Z�m��J��֊�ꋪS.��`�Ŵ5k�UT�)
i�DƑ�K�ej$�-���kW2��E-f��1�m���AD
 ێ*�B�+�naimu��j[Tm��]a�V)��T+
4eT�U���#���#P����Dm��\sT�,m���Ң��-���c-�[u���P-�J֡F6��-ֳN&��[�ʊ�Բ���KZ��A��m�
%�jR��j�-��-V�hX��mթQT+��  4�.٘U�ټ!g�p�<�r�t���v͋m.�I�czL��wϺ�}�@i)>\ �̥ט.�"W�at���%ױrh�����U���� 
�К
�B�C7��6.����[^44�!s�WL�&9V�V`8i��O���`�g��&3*�W�X{]+vc�C������Ckä�L�f�7c���w��� Jj�0�F�	��Fp�P	؂$,�,ЎZ}qN��ĬQ)����kw1�@}�6d3�P��BRbp�N2"�FpȪ�y{���;�):y���n�MW�q�r,�n���T����1]>]�hV�<�N�)6�8�d�u�;��,�!Ph^E;�V43i�˦ll2õ��yğ_��O_(�A�ǜ7�ϳ:r�PҪ��ʜ4����pd-�T�.b��;�<xf�,ԧ׬	�h���^RY�2UЪr����_�%�~�<"�	f���`�.�P�4���7��[���"�8X�]~�E��/GUio�6��;�Nč�΋�6g��GB8������J36�4�1	�`m[����Gy�E�t��S#r&�V�ۺ.�&���3ifu�S�K��HndL{�eV�
Sh�p�
��v���ϡf��)Z�@j���"`Rt�E�%d![�6���|y��ǹ���ݲV�gG�o��F(䍍�@�)���;@�ڿ�~
��ʧ|��m����śd���VK����	��գeN`J}j#�/�vn�U��݈�8��"�5�^r�c����GTϋ{d]�%��v�V���p�EH����wlc�e�>X{�ՀK'q��6� ޮ�MĻ�ua���Lz��3k�:���r�Dj���{vW�_��h� ��I�a�kR('/"��#r"À�8�"�FD+k��ǖ	��{'�����k.,��}Kz��^��`R�.�U���Q�)��ND��z�0(]N�HC�Rd��J�Ug,=�q��dW��6� �Mǅ�>f�J�+	�~���o�!9��]j�<��CFʻ�v�q>��C`���"�t4)WN��P�H/E�WhW~��H爑%yy~�Zlb�P�#�1�LV܍˖��uA�"��51"p�q�I��#��nzjM������su�������%��'yN2�-;���_�h�P�հo��tVG��vX��"hgR�ڜɛL���9�땹�|�
7��b'���%jq���e�Q,�n�M��im�C�����Ghw
�.t��h�M����Yt�͜IVPcbW����ŏp��6����`]�0-��:>���\�F�ڔ�7�2�7���D��`�m[ϔO6��a��EU��o�8��s���n-����Uiv:]F�{C��r�:���[0]��z�(��c��V>ywfפ�%�Z�O��
��e޸!���HgMy�Van��V��m�՜��K�i�u��i�N�`|�F��U|(q�\0E��`#tW]�f�Zx���v��5*6IO�j�nz��s
/-݆pz�6��^Ld�.'���S��!#p���^U��C��O���4�C�ݪ�R�B H
B���[�n�Yтe4-�6�D."�5�U�O4�wY��F���>�+�ݻ��9C*�)ĕ�(�L�y]\�Į;@��zf1�ĉ{z��y��u�3�c§�v1Q.���iq��'�W�z��>������/��7�!2��ll]��Ǎ��.�o���C�X������?�pg*2۫30�1����	N�J(�D��6���:)
w�|z��)���p��� ��̋�ފ��OQ|��p� ���Y.�=tEϨ֋e�*O����g���%�^��7(K�c�������d<g��q&8�ޠA������ì��i񺲾8R(�J���B�i,W�W���߇r̬'N�y_��D�M���&�3����C��[;�̅Ks:I��uY�2Y����W;j^�j��9 �]us�gM ���GPvmz�0������=�Q�S��"E��:��Y5�EU�:-�����R,�/�K��JL؅Ja���\�+�nq�� ;Eѭs�nc���$�;!�d�A�7&(5 ������K8&;6n���(8i�%����*����`Ẍq�"K:IS�Lɡ�Y؋Y"̾�1�e���q�����o~n~:�#���)�����`٧l+�]E]q�pٷ� ���$���l �%b�z�w��ZC�WdAӕ���(W�d j�Bf�}����k�3xW"�>�:�sܰ��Տ��.�E��x�\K<�9��� <5�K~��7�^[�ܾ�r8;�Q�������T�x�����9��0�o��z'��Y��)��q1�\�+����C�V��z�_9i48{��n2�((�'A�1�-	�'iwt2������J��|�B|���w���E�u֋8�}Q���z�Q��Ҩ`3Ħ����qZ`F�tn�/�S��9�շ[�\��YW�������ۜ:����|#�T,>��5���zl�����4e�@����,m����)ݹ��nBS�{�ܸ�q�4e#��.<z�Fo7�h�r�I�zA�T����� �̖���>�p/s�>�n'��E�H�:`o�.��j����Rw&IV�6��dX d����(��[o�ʽ�o�
_z]a9%�U�����(uP���U�g�&1��{��>�V��h�V4���3��mb7�_��~4��uZ�}�M�	嫽z���,�4�2z���u}KĿ��тז	�
�c��Yɂ��4*�����(б���T�XU�� � �Bh+hWD3yj�b���[yѡ��P=�k�����A�fR��e��+��wЂ �An��ԛ��Tl�&�W��^�gw+���z��~�/
R�/P�y�Q���P�`63�a�dg�eAe䋌�7iM�����G�F�{�ر���{a���A��+��(�p���^����/F��V�a����3.�DA~ѓ�ؙ썺�GM�X�٣E�!��}�PT�e��eR��~�ԛdvg��Y�lʬЈ^��������n,oM,l�d���jv�����Gیzzn$�����z��\� �b����Zn�Q� ���Fi�U�5��|�5��8YE��&Ԋ���&�hU����:Vݹ%Ԩ��d�%3�QAfLᇪ#]��ad��ᘻN��{�
| ��Vk�76�Uf���+W:J>���b*V|�@�C��+�FF�m�j��X*3����#�d-~D���Jp�Q��i��U���'�b� [�X���Ď9|�T%�y�Ĥm�L�^���Z�EK�:�aiy{�5}@�~�Xz\F�2��.�W��J���wT�8u���39�������G6���]b���p�1R��R�5!\�R;�#�&�M�;\<	������u�yֲ_���l�|�ʿ��$+C��l5��՞=:���P�ЮԪ���w��n�$DcE���D T9�C8x\��O�1��[��g|�+�nf*�R���3�:�r�����TXP@f�Wh��}%c��N�1Ĉtw�d��J�F�yX�uX�+!�� ͤ�`�H܈�� c�m�����`��x N?,eIy�tŗ�h�,�X|/�So�ǧ˜��,[=₥ˁ񬺞>�)�?�q+7:C'����u��ߏS"��t��K��Q��2ZR�}C�l*o��
�F�V�@�3�&X��F7��K�|���ja�.�IkV�Zk=�s�o��m &o��k���:�����t��{��&�/*��z�+���գIR��KS�����1��lC��}P].�#.L�Rv��oTW���l�����R�b�L[�a�̎6=�Y�0z%�۪k���.���<o1i���o��O�����~ujj��l���m7�*�҂�V3-�Fd\2�ס����컬����-x�7�Ìh:t}oyY�&NW�u��6��ؗ��	��|]U�c�i���i�x�3z��жm�=^��"���MH���,���3Ep��Q��r�OM��x�;V���g�vR���.�N��,�jp�]N�=��M���"�5Pc)����Wqբd3r,׊�ޒd��F*x�r�;��x�q~Wx]�A�q���t�Ehn���0�Sbvo�|�$v$�OO\n
�5W(���E�5B�
�lus�,�Y�,��M��R�vV^�����BoR�g�82_��a�=KC��i���`�,~RW:�$�{�vMܝ���U6�2(��e��)lXt�Ό(�bQ�
!p�Q�0��ٷ���)��<���}+�1=�X���c�pJ�p5�]xJ�5n�}����S�����4^v����ۦ�b���ʗw^gRc=�M�F��l>�l�[E�����s�SR�0�� ����eq����'>mؾ5=z�X1ur�n]�۾e��Rj���Y+��j�Ԡ�9���8���Ʒ]b$�`�u�� ���o$�t��x�S�|4V�s�/��.�;ˌ@��}&��ʮ�W//��/�s��]�+�o&�����Cw�l�}��8�_�T�3�׹��}��ٹ�8���UR𺾸˅��z-�<��!-��׫���C}J�Y2	U��`ߊ`�)Wpa=�ok���&w�>�"�lʫ��C��ŔGx���l/t��̧C�+�T�R����*�h�[���T-�u+@A�w�C��^� E:��"ō
�x,����D,x{��E�Ŭ�k��Nч:ō����lD�|�K�m7�=E���ZO��|�<�~
�}~�=�ƹQs]�n3�ؒ�y:���,�)�7&(5,�zyٯ�7ַ"{Z��鴄�`7����F+��ʤ}�C�4Xt�ivJ1�4�!��W��G�" ��Z�Y�ܹ���R�gջ�Si4u��V�pň��vӸ�k]tE�p��У&�Y�K�R}�Ev^<�rS�s҆�ْ�LP���E�͎V5Şt�*y�N�	����tj)���Z����7��_�f#�f��`8}�4��kiro+1U����|mH4qY�(��X���F��/�{�i��Z:�W�:ɋ�"_K�0�t&m�n��9�V˲⹨o��������H�"�6WPPɜ�Ț}�Z��=������+J�퐃���G��k�+Savf縔!PlZ�(+��u��=8_����{���� ~ٺ:���)c�µ�-����5w��;Ƿ�isי=�eu,��8i�83�;$mc���Ev���#c��J��n���<��ɯb]�>�#�ɶ�	�� �R����.��4�j�Yֲ�A��-Pī�A�|����,���%�8C	�ڗ�:������j�`ûe���+<'�����v�-1XM�zr�%*-x���ZO�>�`��=�T���x5����[����foa�����mdخU�m��?9��+pߌ,�G�N.��x�Y�V[o�����:�X�P�Ӑ��)�
��`��߇�KY�|R�Y��,�Y�l�}�+Yږ1�~�ӀG6�x��^i���J�нt	��L�$�L���M�*����\��YRnkQ�qx�Cڷs�
78�kA;�EV����e��]{��]��&m�f�w&��K����I�+P�0���TBє5u�����VՅ�B\��\+�/�<�+)�l�J9��Mu�Ӫڝn>a�����i����NU��'���MS���ʺ>6����4������o!(�[j��-ވB}�ǆ�"Rx9"V��~��{3�١�=��h�'��B�i�*����:���jW|���Wq��]X�/vX���UT��`-���[�'��y��L�Ӆ�V�ON��_����|�WrCzy��W�� ��rE�=,���L��]On��)��֏o�^��,�I$��g|���	)��>헻��t�QE�]S~WbgsZ*yoN��6�[׻7��f��Ȍ�O�����==ȝ1i�g�Д���Չ���3|��n��]f	
��wo5�ވ#��4�ʇjo	W
�C=K�H�j�.�~�{�u��lů��R3��Ȳ��T��Z�k�4_�����IO���$��	!H�@$�	#H@�~�$�	'�H@��B���$ I?�	!I��IO�H@�~�$�	&�IKH@�v@�$��	!I���$���H@�~�$�	'�H@��	!I�	!I��PVI��pCn b��` �������v���T�UU���J��R� ��AZe	%T�$)E P�J�"USa���	R**	Dm��m��*�Z��R����(AR�jR�Z4�5*K`�*�UUR�QU��ԑQ"�ER�]jRIB���*-
�Z(T�PE�h� -6̅����*#֩Tl��5�* ��AT@T��5a���T��(T�JJJ�BP�T֔
EH�*ETU�'��m�T�h�mKG�  ��jR�ͭN�t�l�@�*����h�U�N�n�r՜�Vh@��flU�uq���k[[��v��4j�jGKgv�r�f[Tu��ӹ�U"�A"�tʕW�  w�䦃Z���Ҷ�]��v�msk��s��֔�3Zۚ�v���S�����\���wj�Ut�f��k���`u�j�n�nwV�]���s�C��)�����ѣcP�   ,�   
AΫ�P�
B�ݦp(�
 ��.��h  B���
 �@
8�]
(�CC�;�
)iw�V�%W-*�.�m�����n�ۮ��C�1֭�D%6eZ $)�  ݷ��t��r�Im�SZ��͛�N��[������,������ͩ����w5��)��tvZa]�l��se���Qݻ*�[����m�J#IT�H��  {OJ���&�1T��i���k���ծ��:�:��f�5���m�whgj��QC47ww]]�����㛐���wP���ACI��]�[�#Z� j
B�(U����  �=����:1��髝ܰN�n-:����A[gMۆ�l��)n�k�]��Z��w��m�u+�a��:
��۔��M&��Z�䈔D�P�@UR�Ux  z+�+t��5��
���j�k�΋V��lm�Jwk6��;A��*ʦ�:��:��un��Uj���]��Nۺ�����sJ
��%B�� 2�P	� �����\k�v!k����u�w���]�MWY;�gZ�A��0uCU5�:Mh��) U�JT!*�)   wsƬ�h��0WUvut:�5�:v*����[hs0u]SA��(Gt�Z$ ��n��
u��ŉ���i�P%D�(vҊ�$T<  ���;]�]�����+���t�+�A5R�tM��T��u8�Z��
v�S��V۹�N��C(��*w:��� 56�ʒ�L@��)�IJT   5O���ҩJ~��2&"��	J�P Ѡ&�CFM0i@�ʥ ��~�_��~��Z^?�����VUy�n՗Z~X��
�������Z����!$ I;w����"B��H@$$?�BH@�܄��$��$�	#	������[��1g�F����w��C,n^^A���bİ(�Ih��ىE*�0hOk^�����ƳCt&�,�E�¨-�r�����2�T��7-i���"T����Tv�QCBs��=:�7�3ik��{��]#r�AS��\QYhP�eжkM%R�O�QoE����ia�Ie��e*��T��ޡ�76��7r7(]�a�)mI������Vu���4�Un��5�t
Bse	*�-�V�ݝ���C6½v	,눗I����ī(&��n�b�eG.��66<��*Bʷ��s\c0�5ynj1\Up-�7i;a�~�Z���12�2j1*�5tH�Ec�̈բ��	R)0��I>�}�^u�@��)��������O :� uT���-nb�#hɲ^Gn�ef�"5��L1�P���m,��V�F�pR}�z��[�w ����Sl�-���i�2˼�˧7%(��V�
:Q��a�]L���b/`��V��E�����=*�-��e$YG3J�F��,ڶ#z��y�v�TV�F����^顶�	�L�fې\;�f���nh��N�20|Mͼ�ٽ�f�5L2@�\f�U��
ER�?��.ƌ���R� �'y�na��b�pfr�T�e�eřft��5]ky��K I���Bm�NcS�yB�k���Nȣg,�Y��
�Ii�J�\����ȳD`š���`�&
��h���+\�f�suS�%Ѵ�v^D�I�Vm+��̹�M��h���j�,f!�6Q�;���� �x+� _9��kLtaU�`�4����xȸ�4�������7��@WL����z�N�CY�ZF
r�K]̦�z���X*�`�X���Ն��)�T�X%Y8op�M�eMŹC\A�D�;u6
6��{�f��L��E� ��s0�c@�N�X�V�GYjw�`)�X�Z2Jq�j�����]9�kf�)�X飮� ��e�iw6�;�[$��lJu{�[IJ��KQ�d��Y�]���!��*u��G.��ЩJ��yh�����1	 hMn;�0Йr�^�ո P�$f]�A�a�P�L:�plA�l�c@��VQ-f���!��x��)ē��k�&-�tiʲ�p���"Y h����o0d6*��n�楸�i��jhuh�n�k@�ֳj�-
�Rq�,�F�[��m	nh�r�t:��J�� ����ˬ�R�m��YIԬ/-��z�c��xQ ��7>�X���p�!KL�с.�˹�6 �Ø(�B�l1=������M
���[Os:�y)�jT���yK~1�j�:m�W�����x6�5h�1��Vcȅ��=2����U��TJ�ɸ�IXs4+��V�T��[Zv�T"�)fe��At��X,���Z����y`6kf!�a!uw�)
��0��l[zP��g	�Ǧj��F�[N�[�m"Skn�;�6��l�T�齅�������4sMC���B���e��\�{c8���QGn�U��A�{n�W��f��-ڽ�� �-��h!�B�m�E�P`�Hl�jà�%|B�3t�	&Ź�u�;wC\��X���YYl^�6Tt��*ƌ����X��;.ΝeP�c~��x��܈´jT �c'.��2�i�pl&��V�IaXR��ӧl��0�������l�����h����Ycw��l873K�[,�ES��l�wS. RZ2��Y��\� �t�(	Ki[��-be�ɪ���mҳYZV�y��%��Z�RD�ݠ�(�w���ʈF�?Q��wh|�1X�$��ޖ]�.��|�C�,���{��f�kBFb�m]ml��#�J�N�v��{n��v��$�xK�B�)+lܔ��Os:1�@5&��x���I���gA�eݓ{%�R6L�Ea����V��95�p^	��"�YRi��S�!�e�<��!��ۢ�К�@���`Y���{�{9M�v~gK7dKv�U�d�"��Ƕv�A�Z����YYc���x�k��:5P�pbŴ�ɟ]X��XQ�&�u��"�Ď���-�DW,��� sb�M�V%La@D77)���fۢUK&����%@�
�^5t��.l; ���:HY��N����v�Õ�؅��n��b��KPɩP8^��껽�(�6�<���ޝ*;Fn�.���X�[P��[�ڰm]��F
FTL:։����;y$WEUk����޴��F[o�k����Z�3E��U�U�����5���"kE)
�9[�'s-`Ӏ�8�h�C�F�� ��t,�����W�q�+]-5���f
[��2�@�Г6�BiѣR(�^�[ m.�J�aEn�pI���-������$��w�8��J�\���T#r}u�lZ�٣�+�I�+�覜���A醬�r:��fFVݬ*�2���[	鬺�D%�X,�M��l�3$T5���0�܉847�n3c�A�%��zsu���q\u`b+@	�6#)��_f��y����x��������jG2��{�.#�����I�2�z�:&ɬ��(�b���m�ŕ}0���kp�t����\�!m���x��K��5(U��OnH蘉:�"wzcܲ��{I;l�,�E��(9��̄P���d�`נJ�
Кm}5����5�.�7����m[.D����5]�0f�+ȩkWHV�y1��ɉ��m[?���c�Qk��i2�P8MES��X����I��ځ �����4�)� b�n Br@Z�?+���ڹz�Vӑ[��2���� ;t7��cC��ṡd�-k�r� ���),��#BU���7^0�E"��eG���b�	,#FL�%�I4�d!��]XɌU�4d���e���I@k!�h#�ho
�B��Vj˧�mce��M�݈�Dr���x��[�`ɑ�n�AK������6;�eU�k��t�u�H�ej��VY��͊D��mZo�J�rТov����Rn����bo�"U����
�ɩk)��v�J)
�8�IYj=�0�o�˫��B��d��-/p����5Tq&me=F���V�Uϋٱ;�3m��f�5�	@�1j7��BU��������2f�t��V�Y���m���t�^f�m�@�����f`������a��Rag.�Am}�,jY�=���ה��Ħha��a�t�����5��ST�+p�]������%�V�J=ݺ�VP��nM�*�gItq1�*�;4�7��l��\3r��ՊDK�PÒ�����=1Y��KK�fT�v�\\W@ި�pj�4)��Y'@
֘�E�>��j���`�bH�˘�Yz,�)������#m�9��®��l���R�Ef$en��r�j��^�4\�5�*[p9�0[�r;GcT�Ͱ3r�m� ���4�H)ST~t��[w�#ö�V�ԛ�1ƾ��L6+nL��дާ�L��ZtkL��n�<���Q���AL^�����*�5+��%շL7��*=�f��x�F 7(`vj�R��^���U�o�M�5قM���!�@1�l�`$�������
tࣗ�6�S�m�A�C��
�M�����К�41�JeY91f��3 ��ہU^�J�X[w��y���dj�	�qZҚ�����C���x��F	��vI�SyoC�(*u��<x�A-+V�-���mP6�T�8ҽ��2�I�73-�)����H��C6�e�M�{X1�]m�@U� ���r�O nȆK�E�����}�V��Y�����E�V�:ڷ�t����>%ӻcFQl&)�9��f���B�cva�K.����]Ҕ�時����k;�Z�c��R3pí7Q[����c���̦�e��v�m�����r��f�n��U,u�E�f0l�.��`U�ڰ55y��覰$�1=��"4��bR"a�J��QB���в�=�R��i���饗{��"�dkrF����i��b�7[r)*VkU-�m�ғf];��!J���j��_M����m�5�N��3m��7d�ь=��,�Oo �Xp�a;���6��N��e����G�HE�ݿ|p�RK2Ish�ǉ�����S�V��Zb������Kt���N	7/,�G�M�Zow��)�o+[T�#���H�]6	��+ږ(Bs]f�J����Z&C����jj	ON�7�E������gu�u�l�����B��P
d���O{�Z�gv�r�-9����(jQ6j�^��tހ2�"J�u4����-�v��6���a��-��D�V���<�X��ͦ���V�"�����&f�De&@��O�d��`��YGh�W��*�������@��S��-�T���/T����l�/m��T��6S�ӡ��[v.�e<�f�Q�yA)�2D�V`�Ubuu�[meX��	�%ʊ,3G!�Yb[���;_![��b��pM&���o����,��ĥ��Z�ݩ���r�6��^Y����%8��Nfi�\�qm�,lݫ٨P��lm�B0ֆ�IfAZZ �cخ*٧r����bZ�/ŭ�f���5 ̼6�5����o"�^4�8��'SQjfܠĦp��taW.6r|É�n�wh���&"����I�e�+fb�ܡSp�V
���S6nF����d�(m���
P��XT��YGt"H�5�����V�4���]Rc�-'�3jm�%m�"+S�$�����ڈ-�i�0�������W-6�m��
6�z^�C	����jV��:�MKàǔ�2˔e&u���55"�Uj�ӂ`�R���Qۃ31��l�I�مԳ���w��ܥ��I*���(
�/Ze�Mi�Q��6�(�Z�$&�v�m�˒�9��3������`��L�e�/- eѠ��x�
ffJ��݂��M@]`U�^�j�6#[��@��Z��m5r=&)��C$���fj;6�[@�b<�:I�xX�R����ω�KT�$I���z��+0S
�?�eԬݢ^�옉	���q���K��x�fX�;ɂ�E�6�.`(CZ�����SM�ZH���f��,��a���b�ose)��j��غ�u��kɷȯ#U#�<�Į����a��b��6���0㹪��0'��c�g0��Ŷ�̬s���&%3��s!��㺺5-�v!����XkM��A��آ� j��߽L�ǵ�6�R�!Zv�э��+M�e-ԉՆLأ)�Wb���D��C�1��׹��f�J���KW�@��M<��8����κV�qa&�Ep1* �X]�ె|�J���Vc"��۷���S�9�E���#�wL=T��q���j1[0�k��ō�Z�܃��'--V��� R�V5n^L19CU�+Z7�٦�]-U&���iM�����H�!R��1b�LÅ W��E��Q0�R�`�e8.��eae�F��7U��De�� ���f�(d0�F֗�0d*����	@�g4���F��{h�lZ�X�A�<-ym`���WShɘʠ��mSEc����f��]k�)�ՇYK,���ֵ���-JR����r��6��-XK�8[���R��]D(\��3HG>-Y�^Pt�lY�m����PufU��	6�eĥF+M��4�E6��z��CA�l�5+N�M��e��
��a�R�v�,�f�	��XF�i쵂�T�QoѢ"l�a-�B��.�]`�)6T�VAGU������(�ӇnV��2�=U��Y�N�ڏ#Yj�]���hl�6����d���nm#�T܊��4N��ֲZ:��7�e��2m�V��u��Y�TU�L�j�
Ŋ�R�1Cf�U�a�P��w��*�9i�+H�`��gk@�5�^�`c�C{�ֳ�p*�aVܛM[���R�7P�Ŗ���OC-6�\{2�Ve�1���:F3����m��E;-Pt����p�G.�T�;�1V[	�R<V-��υ;���B�ץRt�J�-`��-��J��',�^C)���
p�+��_f3�h���!�kkH��%-�Ҩ��wal�����ϲX��m0��ՕP�wk����Vރ!�*�5��g1k��٢-+nI3�x��eQI&�!��v«��$�s��l��0�yFc�Lū5��	��T��rCe�Z0>�f��g&���njcs@b֜��%p�K��۔vkו���0�e���ü���V#�1V����ǕgZ���ZÒ��.kũ�U��wS��"լ��`�.�@,T�l�S[t]�e��*���;��b}(�)�H3Z��+0w���%�vӂE�	H	`�h7@hJŝt���Ԩ샎�	�z/i�st�lX���Y���z3�ƭ[D1y�bɊ�r��T�,h�Y'*�Qz��[@��1���*b7Gu�*�b4f�#[X>�6� �u�'t�Y�{��+E���K0ֱ��Pks#�<VZƠb`���z�ʗu��h`A;��)�ܧue+4ԉLsi�*�DF���1O^VƬ�\XM��X��Z�B�
Z6�@1@^6�C��pp����*;��Q��*j��,���f*4�<;.��r�$���Ʈ��d�s)�H�kU@I�sw2�iQA�����T�;�;�ݠͩ��%���%˾������$yX�j�k�ЫU3I�c�{�8Ѥ;+-�pv��=u>�Loh<ȣ:���{}�e��>�x��S��_m�
������9"��^Q]ݶMFd����j�>����C<��)��v���V��g��h��4�,;�]y����)u�$z4������UrcJ[}�ւ���2�[�Z�����u�nʴ���Q��,��k�����$fIK�ʱ�.������Jqӊ��c��w��N�t���ԗ6{!ܵR�t�Ҡ7�q}-���S���:�D�w�կ�D��5��!V-�u/�uq,%�vC^2�����jV�������ViA�E�r�C���v�u��=�L�۷�%�q��,Di�2�+U5�9�<MYC�м��J�W��ǲR�bU��(U���j�b��2�?eY�C-�R�)�bky�=O�wl�}��E�zR��Ut{v�4{��彐�-���V��65]4��6�������;;��#8VK���9j�flf���2r����,XA����*Ͷ{1�μ�mH�j��6��eeZe���KΈg�mhxy�
X��	yǎS32���p�G
s]2�6.�%y/����&��0�I�Ш�nh�)�U���
����L?:�\�{�3��_����/�*��%Xn��*;��4릝;��J��Z����$i�wo�X��i�ҲR�J)�Pϖ§��j����u���T���wm��7�3m@������>@�"��Ħfi+;j�f�d����D���73�Y}-)2 �۝O�j���)[h��4��{�W��΂�U�
�9�]��H�c{�`h�џp��Df��	+��6T��z��L؅:���|��v��Rک��q�Հ�w^*�6�W��)��S8�ŢmE%�SȲq������rP�t����y���Eӷ�ǁR� ��"�x��,��b�r;��]$�7��WrY�S�v�`�#�*��Dwo:�fB�]��=<fN P+���N��?�R�w�d�!�uΰ��}]Ը��ku�ƱI�I�^v�L�+�aV�ȟJ���fGi�4�;�x��Z�_���L@t|�1�Zw\.�� ̴�]C��#�ep< �Ⱦ��k�WpZ�����)m�M��s��7:-|V8>�ڎ�^=փP�y��RUclwmP�����ʬ=ڬg�U�om��,&�p�;:WbW�\]��)>���w&3�a_4�5%Ʉ�9=��+S�0oT��G���7b�_s�f�8�i\���g��,�Rj��2���f7��[����؞����>�#�=�vд�k�gjf��NN��ֺWX���%��,	�4Ǝ���b�ژ��;�u�K��Uij_f\���u�h�;�LC Ϋ
�ܾ��F����r���Bj��N�ȴ�{�o{X�[O��,���9[�����J� �`їdgP]��f�D3Y>�a���EE�`I�1�o/��&v��|��7[�0��Wԝ"{��H�]�?q{ۨ���2Vs4�� s��@��npqn9[I�ۘr�V��/0x5Ni�t{I�N宐��ʹ�>}��Ӻ�V��Np��4��6y��u7�e���e9�ZM졔�
JD�-aL�{e�f����e������<W�w*���QR	�;+��>r��ݙ�YwW��61�Ǳ���a^~�K�$Da���X��f��L@�:��f��a�%���ؓ��ѪkZ���{�UAY}�9Q4:�%]�ں��yJ�(����9�������U�d����wn�m����Rl=����}j݅���T0�u�-�K*P&���X��oV<��W{ݎ����M��S��Cp�Ttj��܂7C�̬u�&����kP�o��59N�wzf_���J�Ó�t�/�so/��K���v�� g�=WZ����*ؖM�+r�<��5FM\��sQ9�u5�*���	��}�.�m-<N�u]w���]%h��-�f�Dܗ��r"�k��6�u�g.�s�G�z���R���0s��9�)*��{z��;��U��\�h��U�.w��0�ݪ=eu>�\u�ݔ.X����sGxs�*ƫ�m�6�k��5���'J��Og1�v�;YWX��fb�~�F�TԹ5U��C��ne���;�5�.h�I;_oQ�Zw1SA����;z��΂+��Z�٬�[+���T5����nf�3�ƕ]L}�9��-��y�1"/�݇�p��㊓�Ud<��T���]qfJ�-*�[�BT[����v�.���4�pнjRX��5��w�
����Bkk/�AU���Y������k���!�Hr*��c��r�j�lfH�I�ո�N&:�ç����r�{��y����I��oK��ᷜ�z^u�Kd;Z�źʵ�oXŽ���B�&t��$���ψ| ޭZ�\��Si�}'^
�����)%�ց�	 �CC�Ϸdu��k��V��+U��}jj�"^l�in�
�����<^ȥ^�o	f��;�ZU%���Y�f�k�j�mp��Ҿ�M�Z!=ـW���k���t��s������ݼA&�-�EX2j@q|S��j:��v��5�3�3��W�R��4vyJ����-�mVE��xSƛ�Z������(*�Tr�U���X)�{y�w�n�VZ�lϺ���=BG��j��CڙYZ��;\.�<kB����BM����wF��0*�ڵZ����mܜ��ʊc�fD��ɲ{ɚ_��Z��h��4+4��+�3p���ř
p��T�a��jǳ��c3Φ���L�[9�=GFބ��E��C�n��}��᰽��>��T�V0��Ʈ��[ya3�t�,�P��E����Z��K�fs�����[��Ch����ū�eI��)�K�n&���k7y��jցp�A�Ŗo���8o03�8���[������=rJ��c5&M�t�2Ylm�p�-0�.����<;�%jCr��ݯ���c&���_����/s�+��u��r�3\�xO�n`�otjx�$X
L���� c�VB�Ռ�Jj�ƞ�7M�"T�/#�Z�7NWÃ��V%�N��`(�MR�M�5a̙��r�Q�q�к�f��Gz��,S�0õ�݌U�;�����ͣC�� �8�+hn��5�]+ j.�^��-�nw��c�;����\�V-��c��&I�s�5s��f��쒖��mC�b��2���Z��\��U̶��T�ך6dX�-t��a�D0�!���m��.���{z�B�a=^�%����<}��{M��`��!o�B��[2Ю5���}�ѫM�ĬPKW�9�k�d��r�'X��4!���՜�l�(������թ֎I�2G�L���Xʃ�� ����&̹YV'X��ޮ�+"v�Y4ktQ��f$�Z�\yc:����=��G"�9s�G��q<홱H�c����;�7 ��9���Hd�԰d��f��]*��O�9��N]F�-�۽�cĪ�Z�V>�;�����7�%��U(�S��4�4���0k�k8omb#(�U��B���qh��`�'vU��Q�Ze�������'�;]۵:#L�m�����פ@w�-4/H��1�f��a�EjҲ��k���h���c����D��]�sS�D������M��z(�;L��]�n�h
���*�nѻi���=�v�S����٠ �Z�K+mJ9u
Q�?*ZF]G{�V0y�e;��-Π5��3t�6@���&;b}�&����$ة��L��i���8�YꝈ%�<ة��<�*	��C3u[
W�s���g�i��U�j�<8�Yɥc��F-��9�YǴQ�{��[D���%��k��Z���v���ݓ����H��QlF��J�C�^˺yS_�:�Ņj���!�EբqV֖m+�V�.Զ��=�ޘwh<J���f����8�E/ct��]�-�2�JN+j��ޙ8�K/R�W��d�ۙ���ˤ�%���c�,��Mv��D�l�-���Xb�7��@�v�V��j���a�D�Ɍ���|��q	�9n�^ �[����h},�y�K�]˰�Z�fV}���S(a3:��S����O�6;�3oy`��Q*b��VWm�����U�	Y�=�S�eK����H�+�B����z���y����D��/7ɹ"�b3��=�Uyj
p��ԯ~ȅ�%&6]��9nh	6�1p�+��"U�7t��ֻ��y�BJ3���8������&��v������(���(Q����3|�x�Yצ�:�P�n�P|��!X�L��^տ��>��+Q{sEL��&K����{�鑍"n/.�f�r�c��,wrT��e�M��Nn�9���n�T�Hw�1��;*�D ��:c	Թe=z1Y��Q���Rlƈ��v���KY�5��'`��n��J�k����Z���!�����^�z+�*��/�'z������L�Vi�dwԅ�+��M��"���ԎAفg*��:�P���օ�}V,=�{�����4hfq�u��_weNe���x���l��TW�5�5�3����f>�'=���P�0���ےU��2��'��mHdF,�{_{պFn8�4!�K�~�O�U��%ZS�{�onѴB���8)�4�0<;�W�S�n��]y�.mAI����h.�LR�gs��j�y�aW��G�씀����K=:�X��볬�=�Z�2��@U�a���#��}b�֞��f	�w�Բ�Y�g(�g1�xz
�A�_z��]y�Z|�^�1�7G/,�	���Q��y��VʢS��G��Pq�x�r��E�\�6�Za㗖S+
�p�Sw��e�j���0f��)�]ˍVL
^N��Px��z]�cX�zX��>�]Ch���/-h�ac\Y��MϚ��6ذJ�;��Ԣ�ZSe���"��X��	��h�kD7`��huj�4s�T�n��jB���ߧ�O&�g$z=b�)᭡׶�]>�8�O5>�s�)���������;�W f;ҙ����W��֭*��y�o���O��T��9��n�㚶�ծe%]��z�g�wM��y�]ѣ�:��]��H�K=�c Y:w�;�ٙ
6�[�֖���J�����qdpV��5����ԎU����Sx
�Jq�)
ˏks9��32�U�ޥ�O��P�x&��������'vY�vE�M�eG\��Rc���PƲ���+5�.��l�E�;.�x��Wv�y�C�@P�|���2����1��_]cWw�P�	�����Ӌ/�,�yL)�r%8[v!}B�naP7�jq�#��q��w3Fw%٭��YÖ_.|�e�Jĩ�tH�9���J�h?hά��HF��%�Z�Ȭ��1����.�.�W��'o������p�`�$�����m^F���4���^2i��YE��6��`�7)e�7 v���f�A%2e������ה�Pĩ���8gWh��i�	���JU˰�Ӵv��f�kݝf�s�WfK�
��Ԩ���t5y�9�"���$�8+FNk��ɔYd^k��'3���n����f���1<4ˮ�-T�f��WA�(IV�{�h�����v8^�^���E�EW���샬b/�:q�L ;.+P#�Ν�.L��v������Y�dk���3�W	V�Y�B=�6: h'���׏0ķ�u]K3�Vz�="4�R̡�an��6����fA�5m��6�O'�8�4�w�A��q�f�(1b�����T[t�AYʒ���M� �NX�.5�� ����h�RTz���3
]�/�:nde�ɨ�r�6�:hwZ����c"�G���!vwfP䦨��٠�͚K��9�Z��v&:�=��k����@��#��m$���mL�Y�wb�v���d�Vꬭ7����zmL�仩����L�w	��;����]� ���Ն�� �!�D$��v1����a�pR��W,���t��bJ;�L^�a���OWoڹnV���v[��O\��Ȇ�s���ğQ�/j��b�V�5f�5�z���|�]�XI:�*�-$1~��6�'�����k�Ь�j�w�³�aR�س1��Lج��S�N�E4��)	������Skݬ${�i� b�n��q�q���Dqb��0v�U�5���gH��ڲ�t\��W]��W��+����g�u�횲�ʍ34չS`/%:���ZB�#\��[rD�2ػwN�)��ڬu�e\��iFk:~z��7^8T�b��ya���$�"�Z3��O-Y��c�E+��q�����ӭ�X�TV#R���Oj��u�ݠ����N��n�7B���	����Ȫl]���,�ϭ�ZA[�,kH���1;�jԘ|��3�tw�6'�n��ۉ(�2�#�w[It��j�+���՘��CZ�]j��%پ�ڎ:iV��@�����m�e����PXø�]Iv���i��j|hũhBQ�]�Vr͵�qʳ�;(�o/u���
��X������.�=W��^�q�ۇ(��y E;����h��*�H�s�љ�8����J���g.J���'�Oxz1L^�E�\�b��z�ha֟_�7¡{��#�"(6� ؍.4��Y�N�5b��t_Hz�U�b�d��ǡ9*����uψk�^�#�]�S�3�ъ����	:q��<���fh�xM�sB��}r6�^�J˔�VN*	:��@x����3�VUՂkm.QGib*�ZX���Ku-�8H@$$?�	!I�sc�|wGM��U��z�&�]��U��b������r+Fԅ�s,s�z/pv�O6��g��c��o'F��C�ъ�I=z�����I�I�QSG!Eu)��`t]�b�]�)�;��Yܗ���,�7B!rȹ��N�W�r	�	��k�
�wu�2x��k�C���-u(�Cb���Gq�ڗW�eCX�Z��)�uu�'xme�2ř����W�,�B�hp�XW1mY��dR�W
Ix�E�]`A����+V�^!�q��T8�[��jr��0p���,"��_n�+�fGI�v(��ak݃3�n�F��d5<�Yh�\�^��#J��;y@���X��� y�t�ڽk�d;�a;��{AŪ�H��%�N&��|�ܵl�|1-[GWUԳ
�2�R�w2X�b-�dy�in˾1ge��2�vϖ���6��7tz#/P�c�&rɴ>��N
���P����uCE�8'�(��wͭsv�^�9����i)d4�z�C��m�uY�F��C\N�;Ś6��]Ю|+�Aӝ��4^��(t�vtk{��v��#Vc�֫
s6�W\6]f	�ڧ�"�&���]���b�]R�M�H��v�`�F�Jj����9��<A��u<�a�êz��I:�*�������R�:�s#pV2��s�8#��K�ࡻ��ut��3�CW/�/M�t<DK-���dWO���@������L�)��e�WLD�T�ksn�e1�t����efV'��]:�X�hY��3Gwbn]�y-�	:�P�7�OE��E:�0U�;x�sO)ς�Y�/.�[�Xz�{�[N�4�n���E
�{�ۗQ �1�p`��8K}�CR�]���K4�-�@8�R]ve.�'3Š���X�6��Z7s��V�Y:�ܪ��HΊ��=jv�Qn�/QJ�#w��KNΈ��
�۠һe!X-v� �[E���؄����ޱ���}7��V���7�ۡ9z���@)�[f�׆���B!��s�̧+�ҸX�Ɠ�j,�pv���ͻq�3B��h�/v�B.�{N˫�kT�v��6�e����UZ��0�^L�Kr)O���Yt��Х��m�fS{b�B7w/B!;����%�]�\a�SNTm<�M�i&�Z�:}��yf�2ow5�Ԋ�Z�ܜ��%��'xͧ"�����Jc�����4;u+��儆�0Oi�*;^����u�r�G0�S*�\r�	Ԩ֮��LY-� %�m�4�
c��3���i��`J��;�lY����fU��R�l|(;c$���Ɨs�G,R�u�)5)��ch2f'WϮ�mQz�3��M8B�Q͋��U�P;�'Dt;M�Ȇ�n޼m.�֍bN�� �=Wʝ&7f&�c�6�׷����a
��^&9�t�=09Ҳ�L�!�m]���%�&���&^C�l�N��8E$t�|cd�9���- 9Vr��mU�*T-��3�yo�#�S��t̓����@�u{���?Cڦ��i헰촟c\��me
x�Q]��ԓx%Z[Y!�p�wkp]����:-7J�����v���7��u�[:����'��6���S1e�ٻ?,
�\��+y�yp\B�q���@Ǣ�����ູ��彩x��|0E
}Bi�w
��4��%�:�&�J˺5ǳn�-a"���+�����}`��-��\�Vm�5�DN��ձ�Z��`�m��e�����#¥é#{m7�n�v��*4�w`6ɕs0��0Vnf��5����էu���ڝ�v�rۙ9"����L�r�X娇�+s����qC��v��sT^,�Ӫ�X�zf,0��׎M�����Kz��7('�Y����NwD��sv��u�;���ŧu��x�}���m��>F�M\�+��My�g�J�vĝ}��ʮ�)n��gZ	�0�ם�3���*�6��yX�BߙZ����/�����]N;�İ�v�Dbg�j�"�2dOW+�}����B�j�w6��N���ǑEu�r�:KGN���n�U2�v�9�.xR������v����/��򫬒�R�������[,��]t*I:gd��iRv�Y�[u1�XL!��7FL�N�=�ʮ�4��_'Җ���Gd����h��3���xU�0)	%�yD�9C)����y�^�k'ɲ:�+���\�\K���1����s�K�������(�����֥ST��8��^�"����Xi�\+
A��Y�c�Y����ί�;�ͻ�E
�}��i����%�]W��ܬ����\,;Pw����z�AX�I�C}�S����<�a��{c�D���u��T�f��;4�F�sm����r�a��o�8<qǳI3pf�}hH-+�1�w��26�
Yg���$�\3h����i�H1��Q㥻@Q�اXw��{�d�@e�˒�Ń]H6vEV[U��
��{��0#�wvM#o{�%]Z����-���}&,��Sn�'�2�$�����:C��Ү���X6֭Z�8��#/��㻊��
�[pr͛�+�Q.�*Ya8�����yKYq_'��^�"��%�Q;�%NU�; ݮ!Э�յ1�!l:�ě��7�q����¬�(�ʉ�72�ӛ3����BozWN
�8x����ʘ�G:ى��Em�[�[�+�6����4��<W� ŉ�o���6w�G=�Kp�Z(Z,<D2$�Z��b?8��E�)s��f|�G[z��o�;yI�д�M�C�!-x�7�xdDOI��*ptt�����P��S_+�*.��)����K�xe]^��88��fYC����$k`�86Ҁw5|�ŗ�j-e�[��w��u�k��6��#�����L7�Z���� �E؟8�u����3����Z�����nW4�CZ��h4��`��b�=�t���f�=���Z7/�)��ޮ�3�u?���yA��X�hV�b��:��En�6��
�|g��*�k㹊��>��XtA�0jJz Y�����ĜJ����}�@�r��$.U�>��C�u>�.�sH��\�6�<$���44�����i����gz�u�43�˸7�KM\8�Yʾ=κ5��1p���Y2�p��&ޞxeEˈk�Vɼ�ͧ�]	ױ�Dw*��ι��[sr��i�<�P��ov��Y	M�3Iiz�|k$�fk����؅mM�a�;\�ءV�M�u�ʸt�C��Z�!Yt͡Yg֓̔Jƶ�ސc�g8MV�U����k�l.f�}��ߏcw��;���YͤFDحHó������q��2%[��zu��7��S��]^&L &g]S�WVs]ٽ���7y����������[��H��ti`����5����Է�ojwh�)'���q�b��К���aK�R�����Vt�]1e���m�c�9[J����OXTƝy�$z�c:[9Vj٫��roR�$�Ք�C'�wDlā�1SwUH�nS�X[�)�d���u��9m�) 8-��:{}�E�Z)�m��:��2�\Ɉ�	��h���� ��Ru�[F��8J�:��4����W>��z���w^��r	�ݷ��f�*�x�B�o^`�i����*_s�G�����P�0}�@'�ڭ���4r�S�M_R۟_^Vu�D�X��-7l.��[�.��)9����9`!۝87\\�W'Bw0&V�.����X�^���R�X,¨ྔ!Ń��7Y�%��~u%t͘!6%�+}�oN$�j=�R�`�r����t�D�8�!����".�B۸e�3&Tσ]?K��"�xWV%Մ� ��(U�Z�1h�֎vv�P\�-�
�Z�#������ѱ*�n��f<�N�f�p��v�#{	�oi���b*#3*Ꮸ�ʝi���ZKFW
C3�C���ǝR�#A9%�;ݢ���ݷՠ�r�]9)�L��Q���8�	�3J0TJtH�e�u������ĳ(*g�JZ�͹֫�z��GT5���E�:XW������hmjkhI�՞1����̦�Y�Y�h�@+U���ft�T�Cgs]���.L٧2��	и���(Ù���)�������p�p�e�[S���N��6v1��11(I%it�(&Q�[����Y�� �63�l�m�t�ʹmb�ץ�ܻ��t}x ;J`��S��;��� v;�pŔgS-�8�7�NsǸ��Y�ؗW])��l���[�C�Wm�'��a�]�!"T��.��w!Nm�sVhw׽M�:�����B��p��S��ց}�hZ
�������\V�������ԕ��5��]�W��l���=l���0��KU^YR����v�H��lt�6e�	\3t��smf�M�7���7i*L������`]�Ҭ!�;Ճ��f�D�����o��+��閕��軤�쇮�r�h[l.��
�x�:}��r�x��-v���"\���` �]3rۭۆ�T�[���z��E�S]��3�  � ��3w���"���uÓ���i�9w=xyT�燲qG�C�G����[�ϲ��LWvN���p�I>��.�ճ���#(��b�e���FES3Q����Ь��h��Rm�HÙٌZ�y�����f��ǉD�-�鹗Y�Q���B�vė������� �buuv� 5-}��$oz�w58� zu�z�o{q%ua<�����/��,�lZ�u�9Ъ}�"��b&�1��ٝ}��v�ԌדzM�uEӛT��[W����Z���ݰ��k-�[�~��鑹Oo5�V��t�i�}�sq�upweA���C�ڧ��5�/�e����zw]����Vv��,F�G�$z�u>���6nNĲ������H�8��Mk�b�HR*IZ���ζ��p��e!�ڽE�@f��z�Rx�j���Ʒ1v��7ӝ1�M���B��b\/��j���D��.�ȱ㲎S5|MH��Dؚ28��Z�{doa�ی@e���fV̽+�2�cP�T�*�Lݣ�*�\��qt��mu�4^��}܇<�Cʰ�Ś]&���`�"�Wm�2���6̛6�aU#�g:��7,Գ��V+��젥�Mh�.�/7n��F�i�	ch� 9�m=���B�,��w�];����[j�C�|����x�/wJӇ�}��ˁ>��K�Ձ���xz�|؃������4#V'F�t-ig�:p�\J�J;��v;?:x5Wn��xl� �4j1Wm>�ծˣ�uӫ\DY�Sn��F��\]��ua�1�9�y^l̎���~�=R�W����e+Ţ#b�E���9u�2���(����Y1��1�H��f<�s���j�O��x�65�e�拧Q�4+r�Eh�̫�į����c�u���3��u	ΈY[g59�z>)���\��G����>�L��6�f]2�QH�B��Ɉ�ugw26�XDm�]��:� /u���n����5,���Ǧ�+���^؝E�_Qm�#\r˲.vv�I����_*%�\|˾�:����3d�pc�5�W&G<�t!;�F��N�<RPν�v���TA��be���۱��{U���:=��]F����飰uDt�#��XW���&BZ�wOo���ղ������;VL����𭾻���S���8m|C��F�qS��2j��e�_r�V��)���79OQ�إm�-�N�z ���[ҕS� �0�'���%�C�-r'�'^b�ͮe+S0��\kk�k���[M��y̻�$8$zIL$�2��-%�;,��<'L���8i�����o��\s2;L��[�u�+�e�#���2m(�am��{�(�k�ǆ��;z���<���S��ܛ�e�
̲1�骺���j�L��ڳ�=����m��l�k�t�p/���ኟv�( ��%��/�U�LBV�$���ɱVSa �W-�{�:�ީ��;9٢�N�!<�\����SBėc�^�8M��6	��F��,Ly3��,��e�B�|p]]ǔ��J�Ά�<"}C�7���;<Pqe������JT�9��ʵ��ۃ`E�u�:Kb��yOusl�Ӂ\➽�dL֎K
p���.ΜXn|9aC0r�C�FdD.(wYm:"�\y��[���]�_	��w';�ŕD���Ur@��s{i�L|�F��Af��I%������PN�r�2��C�r�4f3{����[A�F���S;���/C2���l[���x.V�\�e9:�U�����5��Rà��X�zg1�/��b�X[���)���e��\������\�!��ᮜ�&��Ի�x�^�IP�h,�l����?�U��7��BѬp���$��v�j�tZ�a �u��w�o!z�j�Aw+�W�t�/otIs��2y��G���X'Z�ׄ�uPe���*-�r�V�P=��p�hV�/���x�3S)���%&��i/���lҸ�e1n�-'�ۋT�\��g-���dtgT)�T�^��W�]J]�`i�˺�����"�Ƕ�3j��mr3��ö�w	�S
5 �{D����KY�Zj������e�1<���jʵlfu[�I�:n���K騤ڬ�F�[��G�Yp:�j�i������S�quXck�U�#��qn_h�:p�f;�zn��[|Q4_aT{&־%Wf�����E�,
�N�{��B��������x���b�7�g0x�D�aT1�DnVP��(�yoc1GwMYK�N5b��9ztQ��x�
�v=�j]N��-�)u����:s|&�ثк6Ռ����xx{��%5���]49^Kro,������q�Oގ��.Yʶ�� 87]�s���ϯvI�����y�ʽJ��tBޔ���#��Qh�H��r�!��nYޮUn�).�����M�N��3�U�li��6���+YoOm�;O��|��q2�=��;")M\{:��7�j]a���٧+m�W:GL��ԍ����3kA=���U��d�P9e�����(���+D�P�3�f�)Bt��9����݈�E���̯����{�")�ݤv���dį�=C7�L�o�j	��
�����n���f����|ck3cR6+��ѫ��5�}�"��2|-�0��<��Z�7����t�˱�;��66�ES�cB���b$/*޺&f7Vؕ�xn��-t�����܀��b�g�C���U�,�6����'H��\Ij�q$�9�u=��q4��Y��w>/4�ЩX{�8�]�j2�$]�Y�gEת<x��Ŗ2�Ra���ڻ�4�z��V<|��X�'#5�cx&��o�>�{��X��^*C,��q�qo_C�&�O(嵻��w���i.v�����S*���5�Fc��S�(���vȫ��-���n�
u �ыJƮ�7�_��-�i�`rw[i��#�v�ߡJ��b�-y�q�VF�S(��8P�2/�͞[G����]�<����ԢM�]�*�s/U�V�V��9Zkz�΄g4��"��MNܖ�)GWA�0�S��=��2���f����~һ�>*�~���J�+
�e[V����k
$b�*�EF,+b�-����UTb����iQb+b��ZP������PDT�m-��Yl
�j����"�V,DQUT����Db�b�2DUm��Qc-,UiAJ6�P�F(�TDQ�Q(#Jث#Q+A�,�b�1aRVV��(��h���DUUEU+m�(���BҨ�aeK*��((���TDUE���V"*ԨZ�kQV�UAb(�`�X����
""
**��E�QT0Th�V�U*UQEU+h**��DkTDQ�EkX �Z1Q��EQH���[Db1��@��U%�*�aXX��EJ�E��TEZ�R�ʊȪT��-��#���V�kH�6ʢ�ڪ"
�"0PQ�Ѭ�#�kB�~��A�q�ڔ�C�ڥ��Z��xR٠՛,<W�;�Z�{��L0b<x�i!!Y����	Y�ޭ�S���Y�B��;�ҝ�B.�6f2-�����l�m�3v6��j�,wG,�j��ݨ>�}���lW��\W�f:�r:=7����=�Chq��A��EJ�4ֺCav�q���ה�<'�BX
��;QqxG#|C��U�Ь�D�r�Q8�2�b�K�&���[;p��0����N�n�4a�(Qҩ�w�������X��ߋ�:w%n�ľVNz�������ݜ�I���#�8������LOy0��?%;�Gy��;{�o%�nn��v�tҷ=>��K����R�¶d8���*.��(��yݫ݆���5-pͳ��4��/�eqdW�k����KJs�{����D�:���Mޘ;}�A=�>V�ӷ6��\{S�|����g�ta�;`���_M؛f�z���mE�W��7m�������UU�Ŧ��n4l]�(�wQ�����*����+3�8�࠽��(����Zvr�Y(B��R٫�D{�Xѣ�R�FN�,�=�n�y�u��hI��=Z����{�m���L|[����b�<�+�&��WyX�W��l�*��<�֋���!$E����.�ׄ;&>�[Y��v�J�����&����2�͢�x��i✦���RU�9���qbwu�Mp��u�@a��$o,�o�.2M�^2y�wݠ���w׉zy�(���<S� �����C.n0�����Wt+u�N�H�������:��9�;Рtsw��mzow��y2��>��z��88P�dVԴw<8�B���T��<���� ؁��F��䷃ܤ&Tl2�gХ�ʢ���g���yV����4��%if����ںR�|w[˛��5TL09K��eϺ&��}j�~��"����J�ܯ�לmwU�� �9e�킥��v�Þ�ƞN�-p�KE:�B�L킖�LМU�<�A]�IM�����w��41�Dt0�WC�.�^�Դ�w[M��( ��W�.=p��R="cA�C+��<+����/���4Zؔ)��t
������=J,g5g��mJ��Ɇ8A�v�˽�f�ov7WmK����Ð&��qw����=)NÛN����e��yDB��&']`]����VN�H.�酺AbE�dc�O�j9�3��y�:*6S��ٱ��a�b��ڴgb��ҍԦviS��9��]�����Y�;@I8�Ѯ�C�[pS��=���r�xƠՕ�h�)�i2L�w�)Mr�\'Dr�Շ{�V��}�֙�Â-�xa���������.���%��9�.�$5r�v!�˙�Q[���|^����V�
1d*Ɉȴ��
΍.pT��ݳp�h���l�vkt撌�����c�w8OX>v�����Z!�xˈ�A\�c/���쑡��kJ�A�*�tU{�qL�ث;�=�Y�_�r�eଯY����Vi�u��G��n��\��A��NrbVE��~��4]o)��Y�:��<����{a�����e�6t�������B")�]��;��63��{YsF�S��~�67�nҧ���BGf�:��B��)�'��N�ݯ�VZ"��B�Ly���;����+@];'�;u1)m��*�H�U��k��f��Kx �vU�xVM_r��bǟ��b�x7��_^X��ŎA�u�֯�Aq6;*�����=�KA�?r�V�^��`sm�׺j�q��(3q�y��
Uf����V�o���g�-#B��A���C��E�t%m�]� �y9�@l�:�����e�ԙ����*��q*+��!W�v<�����&�2�4��K0����y�>�o�2nK�K���ڢ�R��U��X�b�I��f�K&���p� �8��+��h���E\�<�SP�`kމ5���9��]i�j��B���lĻ�7u�Em`�3JM���O3k�>\2�s3���7�P��õ1[�2�D�M�7ܸ�5Ӑc\�E�ZU�t9�
��o�P�ڱԋ�j�*�F�UK��)�5e����L�b��@�J.�B⢮徜�r����Q~���Xn����C���ZǏ��,�hm{��]yN�PL�lpR�,|>�;�dd'�����MS�\r�=�;Ɣ]k��^�B��3��d9 ��\W?l�v�V@0d�ˡlВ�b��l�2�q[;���u�z��
�Wc��m�=Պ��E̎�k�3�o��
hj����FQ\�9�'p�+�{�%�����v��؃>3���L'�͟A�Ǖz'iEX�vt��6ԍr2�U��ą�t��p��WP������S��@����*{��h�xm�t����s�vjev&�s��aƸ�BC|OuNOk����2N�qvT����p�̴�qKj�Ȕ��l���o�ԃ2��!w\Q��(����ܪ`�.{u��á��b }q5��VO	BѦ���Ud�3*���V�aUN�2/P�9��(��/�YX���Kr�4�t9D�l0��[��Sy��q�q��MMd���g����F��g"Q��#�W{�Fa��a�c��Y�5�gWv���n��vc�
�M���֠��1�=0�R`ݧi:"e���uf.�vɫ��&�.k���[��.��'K�K����W�����o;	j:7A�m+�N���ӂ+M¿A�F��%���Me^j��t+Mv-����6H�2^l�5�U]�������WYX������ʳN���MP=o��lI�f��.�2�"�cʹ���r7K�" �lpF��nf��=���=Y��;�G2��%76��A7^�r�i��l�mQ���,�����5ˑʭ�^�!�qq������D(�zӥ�+��G�!��Qc�߷Y
!�>�Ʌ8S�X�G5�$���F�\G��,BW�B�%�G�l�|�:�Ӧ?s!�y��=��K\�)��36��7XHP:��B��c8(Օ$O��B��&�6Y��J��k�:�fR�l%=i6u�U��W��&=�T��¤�Ss�m;f�⌞�1���VN��nO���q��`,7I+qX+���Q��:$B�,�0���p*27
�:�9�⚕���]g��(٦�,�V+|zϷdh�=6)<qf�{|���^%�V���A�7��ẙ���L̦Fj��� z�gv���HU�
l ���e*����[v�����Ly�\�+�j{�'���{u��[�.X������̭�)㙝|.P��1n2bT�ӗdM<_Y��F%���XӦ{�R/�/N��v�-��ExKw�M����CY����F�jw������(�͋H�%����g8D���c}���I����^9�	+���Lδ9t�_.�m���]̏
\�w�i�ս��WX�8x����P��ް]>3��!�Ct$
W9�쒙�]WtE��n�Ym3F^f���$Ĥ�L'�2��5��d�B�K>(����κ�𹽵��:J˻��I�>[�x`!� 5�t=������(��3ҁX2!��%�l%	D:�0�V.�c��Ī:\pF��
ҠK2�ע�'y�`f����׽f&��n�tZz��:��{wy���c�G��Y��N"Z��՚�a�5�9z��g8�w��c�����u錞�|�+�n���bҸp����QK�ZXꋞ<*[�����.=j��������bxa����{�^]oe~�ba3�8p�}�?�l�Qt"?uOu�~�N��ec�����#ŋĭ���Ǆ����Wt:w_k��8J�Z)��\�,�{�����U-WA
��C��QV�g}ܦ�dS^W�{���t2:.�÷l*ں���1-Я���_<��0.�÷��b*`��Wq��=5��ǹ�/�{F_m�J =�uC��3�{�][�%��݅�����L &����~�Z�����j<x��5yܤ��kxHp�zkF�X7/�~�|{<�#(-'�cW���*��]�û�;�d؆��
�fc^��v1R�q8S)���=J.�����Wg\h�y1��� +Fm�ھR�V�ʁp��)`��v\U춤;������v|o:����|酊.��Ir�װg<��t���d�>Ŕ�����aѵ�2�V�ˊ�@�yւ��Vx��}��wKմɩ�{z�F
+O�Ǳ��D5έa}S��t0>8!ç4�%̼1m���cxYJp������?��������GJg})F���^��-���ty�2ڽER��4�9���c��(��i�k8Lő��;���̿�3\i���#��Or^�d��٩�2|1��A�"{��W�7�m�s�u/�\�B��>
Ə��W�ꇖx�tJ�Лw���RǙ��s�N�Vet	��x[�e�Ǜ�˚6��!�z��V\U��]�XJ�D��b�P8%Y�*^Vū��ϔN�����A�	=���:�/:��Y�4�U��E�aL���¨�u�8}҄��� O�v�qf�g�}���v[p�R��>�tpə�T<6��|У$X��x��l�%�}\	����Vҝb��TC,(����kT�f�w�� ��i[�iG�	�P�R-�Y���sV�C�+w*�4k�R6�C�+]e
C��;p��5�
�����0�~}�e�U*;-)��dt6�Z�k+g�#�|������F��e냨UvU2�H�j�4�i꜅ܗL���;m�Ǻү��K7��G/|
Ţ�$9h�&�
�a�bv�G �z͵�
м��[T�PeG<�V3��
*_Sd`u;&�������\�����]�R�}�k;!TeGG�
3ŉ.)�Jz��X��u�A�P����*��mN�72Ӟ#e^��f�w"v�TSxF3b�n�T���(�.*.�})�
-����lm{&��[|��J=�3���l����VZ˫� �G��s��ll'N�:Kw�nq�{]��f�z��w����ʌ��ب@�	ˉ`��v���T�Y��GSĎ,��n׮�"���uYN�N���
.ܸQ�2��7̾ف�0}�j.g���_��[~W�"�����'\N������U������"�!2�͈��wp`\8��'�a��������ڏz�P��Xc8.\�	W.	�݉��kըw��fy\N��(N.�S;�NfH��k�-�r]�.�<��a�5���=b��3��[}���'������*9�np�veoV񲣨f���%�c=�V*W���-$V�����i� H"F_����շ׊����(�UY.Y�!�b�b�l���v}���
�-�X���O�<��㈩�pT����._�F0;�{䕉f�v�{��u|/�
5�5�`"{�H�qMxd��n��y]*�e\J���RY�X6 N�Һ�X "�1���C�8�`'����H6������j�g7K+���m�C�l�ߚ�'��d�RX�,���6x��E9�e�\�����}cP��	ݬ;�,p�yX��zH<��{�v���-:��s���g���o}t=��k��8s��4w�}r��{[�̡u�,=��(�g�e_�F6�tg(���&��v�<9�#1ǡ�a#C�2�X�(��Eڧccp'w���[�x4e
�0x��x|�ެ2Ԯ=�WQ%K�P�;�EGD�nTS)��0�B�7*'2�G8���5r��Dt���������.�gڐ�|����\�+�5|��

�睿C{�}�jwn7#8����\P<'�B]"{��Ѹ�a�QB�q�qrr���JY���S���is&�r�dQ�]:�tw�7I'd!���ƍ�ʕ�;�:�|^����\u�\��:;�Ê�U}�����T��y#�˙���2ʑQ���mp�w|֗�K=�������iT9}�;'غ+c���1H���PW�=����mS�>��O=Q91bqםJ�}7�m֋�咡������CG��|� e{�d}�H�a�{~���r�p�O�jOeBц�C��++;�ꡊ�60��ǩu8�i_�=���;$B�Rak2������!fS��F�E=��L���(�,e��QiiN}�lG����_Ff�8\��Z�����f�z�y��T��?!����W��oS;`����r����V<��cKj�w(�'/�\�ɜ=a�#���UlB�L��j4���:�����Rqծ1�	U�b`?59
/Ǫ�J�j
FO�L�xl����8��4�nڱ=3BO.i�ws��yA�i���ޠ��/��13���i�1����^%J[���V���x���s����U�z�Z�j/����BߥX�l߲�B�u
��Sso|�źrt�"�ʜ���\�%0R8 K3�n���i�o�y�bz�뗕=������3e=��BEN����!C~���I����{g��c�i{E��6�����O��j�yc�=����yjW@�e��D/���v��_��_WJ��#&��qIs����_jXP¦v��t�[h%Ҹ�g>�a��0��t+�e���j��3ۏwoc�9��)���r���y�\'���}X���83�T�0b�x�L'��b���W�qL��[��T�ݘ��q^4�%ؼ�iu�Ҏ��%��w�mm3��5z��7V*^���K�>٣n�ۼ֯��
�J�P�A��wp=��������M�r��,�5�s���>p#+�նoen�"���6��ࡉ�k+vS���t���U��gn�c2�	\��p���uu��yAZ�����)T��s���xZ3�s�F�y[W�E�.í̴��/(����*݊�8ְ�p��V.9����iP����'P�u���{�x�0G
��ݵ������{Y�4��j�	��c���l�A�!ۉfXT�7g&��'k�IE�w^��-5+w��X��
-Vw�Sn]<���聬ķEn|N-��K�NѮ�N�'{2֚�3E]Lp!Zz����] R�sL�ĕ�e�$�LU����u�6��k*�JP��rw���Y��wZ�s0
:���O��x�wvhe�'u�ͮΫ�ǹJ�\v��yK���6((����WJ�[ aG���wת=�F��21�uj��u�� �qB�d�f���wk�]�rt��>���v��ү�%��=�ą����lfD*쾼��A�c�������w�+6�at�ρ�B>�:��l�!�9���ܸR�{�	��s�\�v�	��i�{}33棦; ���2�k�F�������jӧOKu����7]�	t�x-6�'�.��̉�Xu,��G3���膧u�6��emgN�s��8E;�+�V�Z"�A�Vܹ��Y��v��\�fT�
B�إ��,�|�{S;��P�]�1bJ�α+���QvWK����`8-cwfA���!��Ѱ����>z�������c�X.�
�S�5>uk�rC��`mM����h�xpZ(gU�U	�- a'f�T�L�K:��.&hӆQr���a�n��J��/3p����-'�f_,���g�T�m�
F+&vٍע1J԰���u�P���ʕi	]�" �S��Ȫ��N��8Vw@s��SE���pm��Ә��eW3"�/V�J�mÉ:�u�i�r�C�8po�^��;Iժ`-���-Wj4qZ����e%628u��AN�H�8H�Vv���yv�+��W5L�{���bH�壺ژ_����~˽r+GlUTX�V��T,b�D�"ֲ1J%�QF[R6�bAV#Z��KF�F*��X��b,FEʅb,bZE�YJ؈�JV*ƴU����
#,��U"1Z��b��[ �E)F�Ŋ,Pb�m�,AA�X��A�AQX�b0U�UQ`*"�����F�X"��Q2"*
[`�֑AQUX��X�b��(���DYZ���T-��XŊ��(����X�-h��PX�UEUUc؉UTDDX*����*�b�DQX�QX���V*��$b*"�Q�� �"�U*"���)R��b[b�b�b� �m����QH�U��"#E��*�F0dPF*T-+V*�U����*֤V �"�*�*Čb+AEPX��T[h""�Q֢�b���M}�\*��n��so6r���]8 ��\�w��Տ5��w��w�k���Xio���x���En�=Pj�A��N�aE!��^��?�sz*v^�l��Ŭ<j�!�YK��ƪ0��g�uac���/��M�u� �y��V�^m���vn�n�����f:
/��=Pq9o�NE)��f�u��8x.�:�|�u�Z�,��fp�e��!��i�4T�V�ծɞ�a�6�-z���{b��+Q���Ǵ�G*Up\jy-��k��d��u?��x��ym�yP̜�wN��t�"b�OB��רcT��S��D�(�GJ��D�f:9]�˾�q�}~}�u9�]�t
���'*QҢ�����,�l�0]]Z4�j;��f��bz`\��9�
	E@�㒢��[R3�E�W*�r��;�󍸦$ٛ�V���[�itQU6h��>��t� ��F�b����p:���f������jq�jR�pF���]Ό��;���~�*�W1���_{)���_��h�+�:��Tt�/m�L�/�.r)pn�c8(�|��y�z}e�ѝ��)��(��x�uUr��Ui��yr��oA+�GIz�+P[��`)��X�U��r��h�+Tx�m'�϶�_S���)0�YOo@޲��ZSc`���s�.2n��s�����;�u�t��ۘ�x�G�`�d�C]\R�$3U.�Q�j�}�7�"Y[e�9F��OT	�����[u��%��,|I�;_�r�fY�k�?���`��$��eֺ��4[�Q��OMi�A�gh!���)�3ULj�#��}�V���;K�s�I���P��Ď�U[N
��w6v/�t� -�C�m��Ǵ=����;̊*�*^�"�[o!�
c���f�/�X\`e#f��Э�={9��~Ni}�{��`���o����vJ|�a���+R��s���+8��1KQ��q����9>|;*�,l��}��Z��@뒱����J�K�2���~���E��/_f�fs���ޤ{��{U�~�)y{�ܫ�M���<w�4'�Ec��СaX�.�&;,��X�Fvm�u7r�"���@�:P:
<�3lߒtaE�/H�R#ywT��3N,r;��/twk�߀~J�5��D�M��:�t�:W.�7!�P���'-�H�lH��6�K�˒":�T��5Q���p
�tۥ���-��<%q�Z�{��kn��X\���,�#�^o4[�
�["e5��<�6d��&6	���������{{I�P�L��g�d��HfЏf�M�|9�}K�܇�o�b�+��S�@��O9#�ƞm>��޴��-T��5xu�]귢΀knSm�dN�$�p?ɩy@���e�ɧ��%U^z��*�O�:�����]yN����mG"s��=����uMw;���Gy��5	�Jb�.KmB��a�5�r�	ˊ����y�3�VE�2h��"�0�"�	�#5���������&t�,K��^���a��c�8~�s������qm��~�/��3�v^�R&ޱ��M�Ub��?X΍.DTeˈy6"V���0*�?OP�a׼���Jw2��ے����m���&6����ϰANy��m9�U@�������^��͓8�h�=����;��-�,W��4�X'��'U�a�\F0| ;����ޫ^�o�=:O`o]�*ڀ�(�u��*l�������f[��Pˮ�QuX�Mף'�l�	�8�MAL�~��l�+ޏR��d�)Y~�K���Ur���)�v�L��<.s�0�Z��"��:���r=K��\`w;��s�+i0-:���xx�S�^{w��-���ʷ��XV�_EB~f}8tC�C`ߢ�*׽��5锬`�'���.��d��=�Kp��֌���J �k'.����uf �1���C��v��^�lܧ�G�ߢ;�7��\�H���x�Q����Ԟe�y�z>��c^���A/R��v!���TD�X�I�=����6+z��yY*�ҝ��b�!G���v@S��Q������5+�5�f�"6�b?
9��a��?x�*"�ʝ��n�#h�dd���z��,��]�	Ü+�i�M���Ň��
/�&r��y��S��ژ�n�zL�v�ON��P�ʦ���Y�9������&��)����(��(�=�/��}�h��.ee}G�;@��N���P�u����3R�zezx@Ϻ�̕C�k���M�G#��ە�܌�N'#c����7��9��1����o���A3�)�ZjԲ���${}�o˛З���IdVuU�jC��d�'N���=J,C�p�������1��aA��e�՘Y��z�z�߫�k�"���-y|��&la�
���S��}~|��
*0B�eQ��k"�+s^�1�N����~���s�̥э`idW�k���*--?�u�=����>5B�固��:Qr������wŉ�Ư��3��`Z��i;ɝߏ��H�OH~}�>9�{˩M-�С��.Q����><���UUlB�M3�h>:F��]��}V9�$(y~�����6�e�I��ހ����T���5f^��JF�����.���oZX�'��C[Y���	^B=�;M���>���}i5�v�M?̠�S	[ba6�1Jv�krU�;�YY�[��[�1���bPX��k/-R8��M� �N�a�{����b6G�ƗUr^SPy������X}d"�t�����t~�876�N�0�m���C�$Įt&)�}��ϳ�gj�Lp�_%���_W˻�#z�)v�R�t��V5�6����:B>��$�*�5�@��ro�U�vߑ���!�Wdĉ9l)����<my�0�4-wI�!w����[=/_��Hw��І�Gw�����~�O�bs��z���D���ٮ9h�t�*ڑrs6�<���㚝�r|��p}�+�c��p�^O��/Y��B�������(�	��y�����g3�5�S�Ǎm�������ba�]�a�����M�/���~[��1po���3��,.Va��EQ�&�y�cJ�c��㴪;&Q�Q�g�T.v�c4;���BF��n���vec���u��dL-;��ױ�XR��X��<C�s�zY��<�T��>�k��NZ�~�����#��y�s�
u��@v�R����X[t���ܲ;#��l���_	��\뷚e1��!�ɂ�U���y���TX�{<"0��<���~����o�e�VV�d=ʠ��q�C+xK���]�Ѣwb*u86�u��G�y��{���I��v�rQB�$A��x[�9��R�,]���!Ь��X+�|�>=(��c�&KjE�:z2,W*�s����ᬞYQ��)����"+�'�T9�A�9��>�T��`6�e��z�L��FЛ}⇵�����T	��a)���XAW��<ej����L�k�Z©�zƔ�M-���͛{n�MQ̘�)���V���<π����8K/��C|�%n�b�f�TGv9�Ź����fR39H����`�gz��3�r��X��ds1|w�˩�.5ݧ!~Y�*��y����壶�B��BM_i���Pφ������U0�7E���-�#��GO��}�H��z�&��wZ�x5��t1׌��� e�`߹mG�Q��3���[����6��@��ϻ��]��!��Tmt3���{1X}h��_u�~��u"<g]�5mF�����EAm�~m�`�G^L���k	��C`L1�b�'%a�DT'c+b�^�Zk��s���н�	&�;w��}����Nݾ�޳���m+8t��TJ�`����5_V�`=�&6vR���^ vt&�����r�h��	7�w��u�E�w;ػH�*O�����iK�r�	�: p`M�`�|En#t�'S3&���
���&s.�������ޛ�5nC�K�{l=Z��6� ��`v�+��^����}X��;7���{��x�R��/�������\Z�����i_�sxsyWB��A�&f:&���n4
۾8�7�*�ΩM�@~���[tT�tyS6̀��Qb[vt�gcp��crTFv-��7�l;�Г����j�0� �S�Fz����it99ʃ���V��[��'KԞ�j�%�\[:��g��U>���Qw�;��r�N'.R����Sw��2+�d#�������I�5XF@��Eb9F�ʣP"5w��">��$��~������]��֗�˜m5N,;�b�$'.%�`�;�oV@�2h��zE35i�Zvj��z;"�c��o�֋Dh���ei�r�p���v=,wn2z�?C[u�1�\}G�-��S6����5DJ�����hN�~E#� �vlw*�p�K��%cup`W����s�bt�)L*�o���0�tgr�͊����I͎q7�s^�qB*h��)�7t��&�r=�h���pV��pO�Xu�����@P�^=ӫ�)QR�����÷ZhX��L-���V��Q��OLԥ���5���!V^�u��M��w��Y%��JDv:����s��ލql�Z_W
{��̠�MH��iu�"��n�����k�.���m����I����,�^���VŽn���A�d�ֻbV�~F��FpM�
4���w�����b���=���o*\�Y�s,��el�$�D�C��`��
a��nǞc��'ϐ�p[�L��}}����Ty��0b�-���Z�����,���q`%�~��<���;r?,�GQ�k��ں������<:�)ʣƾ���M�t_f���L�L?d�j�+����1�=%���m���m�],B��C�F#����b�U������o�輆�l�=������-��oOؤ3��dW�Ѐ�BT$��Zi��EBDV�S����m�edğ��k}Q�;���cЬ�K���ýW�>T���C�?r*;�0�����ϫ0��Ŝ�6e��"vm鬇�l�%�����U
k������a�Tz��EiU*�U���ap���3Q���X�>��@�"���vX�qQm	�dBV�Wd�j7^�B�X��M�]��vn��h��OGBEK���c�7W(G@B(�
��c9F���n��!�ZlsVè�K����AE��O��C��R������*��6�ǫ�z�X�+L���74*��m�*Sǲ�p����U���{Ev�,;�t*�� A�Bf�ڬ��h�,1nq�8��U�r4)�;�4C~N4�*�`�Y��7{�jY?�  z�r����[Y6s�1k���5;>�ݤ��a���q2�����:\h���J+ ��wm��{V��Y��ҫE?����g�(<wη��?�2�"c�oi<p�U���%��i��c
/rP����'��KƧG�1\�d�z,�c�Ï-��[����HQ5tN�Y�!�\�B��a���IMy>_)_/�B�؅��fu�|������`ݧگ2=�{�^�����qP�K��������4)�}^�3��kA��}P��*�zu�>R<Y<m; �?{�.b���$�]�t���Y�0bg�����мE"g�]ov�^�fn�<�8K6�����K�5�9��37��x���e~��w(o�� �]e�]	Uh����4�:���qqp�C,�
�p%��u�sw�F���K_=y/`;F���:�T����pJ�>��)�Y��p����˪�̿{�4���r=+��!�mY���vV��E�X8a����V�:��i!�c��6�1�el�̫�{�vt<�N���WK)}���C�{S�n��K���_j���v��S19�x�ݢ�,�KIGI��u�)�)�eos�3�͹e}II��2e�!����l�/19���.��C�V ��rk���5HFn��{������O��b_������q�f�+�P��s��J8�/����uE0@��L��λ�gj���\���r��y�cJ�d�O�i���T(�����h��Y�ɘ�r�gy���[<�U%>Tnڥ�q�zs�=�Q�*V��ϻR�NC����P������^�UF�_3�x��˺���Nڥ�����G�E��G�1-��Z-���v"�3Y�=dmOq�Y8v�E2����;J.��jFp�nV�;�7�I��Ȭ���OJ���Od.����(���|�C�dr-�2�9��f6<��uq�2�%G]gr�tGEC����������K��v|\�� X�f�Ĥ����ky�td�`A�y|�F3�f8��f�q�~�>1׷�Ie25�4`"�۪k�0Hu�����G۾�����Uf��e����r�&Y�Y0��-P0��O0���T0ɦW���g$��0�'cZͰ���7/q�VO�Ob��)4�N�[���-��1�X��sQ�#�ǅ��>�8��.R1��m��d��g#%g+�7|�E �d�)�Xu<̰4���Π��E���u�;�rf٤0����]��L&��RI}{�o4�`���~Į�[�[CWV;�l�N�T�I8�δU������%�u����A���U�Y1#F�䅢Ze�<)S��~�j�����Y�����Yx��9o$�(��p��뛔7�:7�4S��M�P��J�fm	S*���k��P=ٚ�K2#/%�ېkb
֒��}F1��4�[\3��5'��Ƀ���!�h�f�E.�%�r�/�Z��E�X���W�9�.t�
�\���O�Y,D�"w ����Mhu���X�@����,��H�o-K��e[;9���8��&�G�\�	�Z�[L�G��Y�c���+�RG��*P��7�𮳻%�1
YD�Ҳb����7���w
���QT&!F�iV)suƟwVJ��c���H��VEug-���%�/C��J8�[iDd:P禴ғ^�z�k)Ks�l������跷{�EM�A`���ӽۖ�6.R����=�w6+<U9��V;V���ڇo��0v�cKo���n��E;�2�8���*&�up
�p;)Uhf���~���E�W*���!ql��m:}�S�.}cwb�pV�Y�Ց�2�r,q��-gX�K4������B����A۳e�JV�p��#[��Z�p��*��f�傭}Ƚ캊��e�5���7��`�BJ:�7D�33An�;=�Sf�RD�h�y��U��(Yr���wGo7�:�Y|��SWљ�]�gg�^ac���{����4Ӆ�J���@!�\|�f_^m�[2U㜳5e�%��v*q|�	����ܚ�5]M��X�U��	YgM�5�j7b�W�ciQ�4�\�6/��9,N���Z���V.S53�4�݉V���Y��'A.И�vaBX�z�sn��=m�m��o�������+�i�'�{1������_��I�[�����L. 4�[{s]�����An��Y\�j�n��V��K�*��R�
��%,�H���˶�c��4L�H����R�{n�B�cL��� -�_^٬�3Q-�`��V.PLü�X�Ր�e���Q���\�F���r5�ű�N�:����վ�Ej�A>ʾ3���n��X��Ϭ�_�v��?:��u�	3�F��љZ�xo:ں5unO�:@+�H[�\q�U�^�	U���Zi��˶�������tS��M�r�{�6H��I��!ގ�,WL�vsv���#�y9׫�x�p�]�z�m��mu!J>�#�^X�����|�Ѻ=�Q"5{�	����tС��a���#��64٣���U�l��r�EZ��A�II^@���:�)���[z�Ec�`�ud�����q�g2�j��QR۽
��ʷgk����2sVU�F��řY6�E˵�0t����vS���t�1!N+�
쑸X��ܽ)s6�ƄUwp�-\��_�D�v�+~ Ĕ��Ѭ$i��	�O���i9���aԶ1��*|�M����u�8>�b��w�k�,X1EDb��������H�UTUE��b���"-@��%l`�*#Imb"��m�EUA*,TUF*��Qb"�X�"��T�Tb�Q��"*���Qb��*"�"� �+U��Tb�+�UDF(�(*h ʅV,b,F#YQ��UV(�TTQX�b�mU�*���E"�`�Eb(�(�b�QQb�Ċ�Q���X�mE+F21A�������ұAX1�����BҪ-�TTAX���V��T�����Ԉ�UV,QQE ���
(��Em� ��+b�Tb+�TX�+F*��b)1E�F�V����EQEEDcl
")"�cZ�X����R+C�b�-C���V(��
*���TQE��"�A(,E��"*�!TEH���TATQ"��[��AU��(�\e���q���طi��Λ��S;|��r��u0���Co ��ܔ��Z{:��������ٍm�nsC��$���}�����O����b&Dvn~ (�O�DT'�����<Ʉ���ZƐ����`a9�8�(q�\~����%f�~��ZAf?b�bԂ�79�I��<��'ݳ�R0����Y�}�w�~ν��0�L�����M�ˤ0��}�e�L3/V�X���\2��aE>�!�wvL!�S�e'��/�s��4��
�hu�i�
�2T��<̢��J̣��_��c^�s��q�s�qo��}$��'{��0+0�;�jO��Ă���Nfɖ��^�,�L8I����{&����a���~3C��u8�	7�a%gS�l��O�VM��w��|?c������>�>ӝ�>OP�!�L3�J3�~fY�'�w��������O�}�|�=`V=�3'�|��/��2W�t�;���8�^��}���)� ��ɦe���Ͻ�sO���}������}~��sy���m���&H,�η�(i�3�0��\��&����t��R
g����mE�ù�a����	??����>a��7ﵘu�C>q�9�bJϙ+4�{��k����uy�w�.�s>�L�Ag�<�E1jA^�<� �f��u�Af��<�a�TX5�a��������I�a��
��Y:g���ُ�L 1��0=��v�z`j��'�0g>w��V��Ci2��^!��e�XVO>jT
βh�q̨�'R�Y�e&����1�B�`VfwL������6��Y:�Y��&���$������5G�E�����\w�4�8��!���ĜM3��!���e
��N��ؚI�+&�e�2��%x�Xa1�%p�2Q�O�0��ϘcT���%I�6`�X~f�+4n�a��'��I��ߺ�����{����}�b�;o��|�_�/�_�*Ag�+�{�¦�H/����kvL�)>;g��7l�
l�1�������l�C�j��m'���2����ٙ=�@����T�E��Փ�9���o�l?<O̘a�o�u%}�&��a��ˎ�w$2�2V~��>��ϙ��pE
Ũ�0��S,�����i�v_��L8ʊL!Y�L0��8����������~㖯h�m���BJr <XT�@W9ov]^&���\ч�L��f��-ή�Տ��X��EnA��@̳c�w;�r�*S�1�}C�`�(�ʱ!ȍ�ͩh���g��c*̛��fiXK��͜���݋6v�N(�
������+�Rh1��8'�Q�O�W��ơ��:̳ݲa�g�R~B���l�\�*O!\����0�?���ҠVy�����*�R���u�I0�t�a�2��Xb-������u]�g�Eu�Ͻ�:* ���VM�P��9`a�I�h�=�H/�-0�:�0?m�@�Vy8�	���e�fF;�����a�be���a�k4�a���fn���t`]D�������� !u=3�C����Re7��i?2~p��^MPXa6��ܳg�&Y+��Ms�6�AfRh>a��)���1����7�q
�!�g�ﱉ�������־�w��.}Y�(Va�C	�}�2��~g��C,5��8�0��
}�b�Wi�L3p՜C(q%{�>��
¡�9z��!Y�J�M0�h�~��0�bԜ����qN����7
��Dǀ02&���ƒq4�H/�{ܜa�q�aQC��Y�L0����&R��&��i�
�ĩ�����rɆ�������,�N!Ryؾ~@���1�޾�?G{볜��'x,φ�1*fY�P�̨�'��Y�J�W��ٓ�oT�C~�6�_��M9I�P�6ɌP�
�\b�e'&���CI�1�Xu�`m�JΦ�z�����y���������� ������|�)6�a���2��%z����-g�/���d�
,�߽�9�4�R{��N2eæOӞ�M��¦3��g�3�J���yJ�Y�l�y��og9Ţ�V���U�f��B�L"�����ݰ�r�?5!�gΎY�eE�<��+>g��k$L>C	���~a���~�!���&=�0,6¸L�c��d���G�R#;��ɱ;]׿r����� $����_�
ΰ�a�aSv�^Lg4�b�6$�<κ�0'Y���i��:ʊ|�Y�L0��w=C	�M�׳6�?0�����+h魚����b:����ǌ{(��N�����<���i>B��o����|»�!�IP+5��&Xy�a�ө�~d�0�n��'SXݡ��O>L����f�=�"I:E����=K�_������mؽ�R�_ճ۸��g*1T�L����!\�ֿ8 ��lu�,�Wf�h� �OZ��z�00W���*�q��a)9�<9�N]��N�U�9
��۷�ND�[wo�Ov�k�W`�$\�=��F]��;��J��s4�~��b�E�hE<���0<"<�{������@�_�wiY���4{��@�V~N'�IH��O�a'P��3CL˶,:��}�e����9�dgY*A	�OfβVs�Nw;3�}��.�����]���'Y6㴞��i�O̞�~���>d���fOɴ���=�xé�Y5;�L�0.,;��g`y��o{5�H,40��+:κ;f��!�I�Ϳ\s�������W}gUFd��=�G�t8�� >I���_c ~@���Ǹ$���~�0���|vɦN03��'�Y�����
���#���e'_3l���*�����=?g�,��S8�Ƴ�2���m�|�R�?�Y�Y�F��,��Y�Y97�䂓�+=��I��B�}���0��7�2�ha�T
���y�L0«=�{���g�����]����x6��d�1��/�N&�p5�i�awd�y�q�L�����2�Y�4r�t�������~@�ï�l�q'ΐ<��M��fH(���p6*=��ۣs���K�r���9��~�9�8̸b�.���@�V|����%@yJ�̛ŝd��V
M�q��o�&Xm�O!���I�$�-��&�	5��?2i�&@�#�
<��3;>��~�e}�3�U��؁�RǾ֧YR6{��,�����ǐ�A�'SE�'�04�z� e8��ܶE����f����J�C�/o�a�
�1g�<딁�ti�������8��s���;߇�<�޹�{���>d���1�c)���{�g]��<���L0�}=��i ���k6�!���3�f�^��9�rɶVw�3E ���wn���6a�5�{��?7��|9��N$���C/�a��C4�\%d�~�v̲Va_[!Y�J��{���&S�r^�e��\Y>Opq�$i����{��H,�jc8�{�0ȷ�]�>g�qZ����J��C����. Xq��X�Ơu+7~����2�N�d�N&���&�_1I]}��0�5���ٓC2�Rk��e�a��<���M!S��>~��a�W
�=U�t8t�΢����6&��Z@�}]b����=�)�4����[�U3z4� ZkTE:9F��cp����z;���6��2�Ľ!�됥+sa� Z�D�h�=�!��+��@�����Y*��[]�jee�����z�0��+�\%�B(� {��>�>�:�}����� �����t�[6�_0�0�p�V�<�08���VΠ��)����b�gﻉ�4�\0��u��� _ZG�����"fbŇ_��ʷ���5�I�Xa����	����|�����8�ᛔ?0�R7���,�
��8��l�:�9L9H.�9�g�\$�>p���a���O>�\����iY�2��љ���1���?0۴0�}=w�8� �aY��`��2a����� (���/�e��L$��vg� ���0���0�HuqI�t0�̕��]�VB���4~��2�����3��{�~���s�������Ϸ�|ǉ�ayd�=�O9H,�&�k�ԟ��AO{�M�I�P�0��
�0�>��0?5�[�m?0��?b�)�y6�	3�2i���r��a���y�1��~޻�W^�Z޵��%C�TY�Oس�z}�L��<ɳ�ƞ�+���s��뤂��ɞ�2\Ҳh�2ϙ+��	�R���Ľ����`u���~���*����x�;ԥ����ݹ���\�^��1B���H.�y�Y�I��͹H)�ԛ�1�a]s���M��{�&_~�0��\�P�~r����tβVe�MZy��J�9����9�ﯜ�߹ߵ�ߺ~��=�.��fL��|é�z��a��5�u�E ��a�:�a��0����i<� �a]�s�>M2|�����jM�(��~��w��	:��4��W�P0����=��<�����}�������a��qC����gY+�r�EY6��dق�(WL�Lv�7@�0�Xk<�C�8Ñ;�'Z�CV̤ۄ��3��ę�b#��eH��l���v��|�m�g<�a4�
/��bM���i���y2a�����Ap�Xa��sg�J3��5�L"�2{u�)�B��3�~t��Xm�����>g���@��G�P��8A��e��Z��Q�g�>��J�S���"�^�.���ۆ�8��Y��&�g�T��0e�αM���y$���u�ެ	8��9CH
,<�W�u�	?!S��;�W�?>�.9WC%oH�D��ׂ(��T9<6����<�p5��Ei��K�*/���˳���tc�1*�d�$���K�?z?O��=^�]O��]�'m���Q�skgXl7��k˝]I<�����h�1-�LH��U�
��9�{�ܘq���xxxR���$ԝ� {b��	�?y��2�Xu��'�g̕�aSF{�h�ϙ*l=��8����'���ct�Y�L\�3(�^r�0�i��!����m�A\ ʬ�{��#�j"�~�������n�3�z�`V�m����(
(x���ݓ	?;�a'���2l�����8��'5��
�2V߱2��a+:��ｙ��f e6s8����0\�
>��<"=P߮qa�b�o��ʯ���]c��s�ֵ�s���E	YRe�O�a�偆�Uf����-I��:�g�� .��T%gS�0�;`��M2�f���z��a�����d�<�e�2�����)x{<Ë�}���{�u��:�hT��%��R��y�&��N��HpƳ��J�򕜌��d����R�L��ua��2��]���gPYY��!QH,����n�TH}T�9�tl�b_�^��g7�z�ha4Ϙa�� ӄ��=_��eE���/��&q�ֱ�?0���'Y�C�:����g+4��3�֐Y�L���C�ʐ\'0�g�\$�5��<����~����|�=8� �/�VeE ��0i���e!�;�L;I�a���d�>�e�d��t�!�wvL!�T�I�+��~�&�~aXr q��& =���c93ԍ|y�}J��뷝����ud�Ve:�	2�x��ﻓo�a�s�����<H,�~�d�l�j)5�`2ͤÄ>M&��H/�
��`+P��P���q�jj�EIY��c�k=��c�{���x����o~�O�VM��}=L$��?0�!��:�Fq�Y�u�=߷��J��T���d����Xw��2��|�����V|�\2]��!�q��G�m2�Ax���O��}���s��Ū�M�q����sP<0�}
J񒢐Y�����~a�d�˚O��u�����S���=d���ϳ<O̘I��wH|��偿}�ì*a��oH��q�����U3_.֣&�O��8��{�|��Ĉ,��x�
�bԂ�`T�:�᜛��뤂�3G=��2������|�<�q.�y�Cg}���`u��ϻ����L /x�߳ﱬ� ��c%��4|���7��oX��� 1]/N�!�v+,N�B����(��Kz/1']�Y\�'�a��p���PE�@tKj=�c4���*h$uB�o\\��
eZ�XB��m�8z��b��f��>9�kݧJ�y�Bz���)I("��r����R:���VL{��cQM唏i�wH\!�L���x{�X�N�%0�m{���Y��0���>C)?!_����!�aXm7q��@��&��C���'R�Y�e&����ŝJ��Xa��=�y<� ��6��Y:�Y��$Ǯ�&�/}�+�#u|*��+j��.��N�YX|�C��=�I��1�&�s��(+8�M߱4��VM�ﱗ�)+�:�	�L�f�TY��l2��Ϙ}ٳ��&��u��aǀ1�q��'��E��P��d)φǆ��'�\��{��̕�%�o�*Ag̕��*e��Ͻ�[��e�I��Β�eX|�@QH)�_�P�4Ρ�95I�L6���rM٤�0<8o�>��b����u��93��=� S�|���a���T?$�}dپ�'u�C�2��He�d����f>��ϙ���4��P3�`��L��.�����?_��L6<`Dn#w��7��T���dm0~g�2�a��<n� ���a5�`�����������&5��)?!Y��7��>B��˟~�a�
����C��a��p,8ʊ�u.���z�z`��&w�L�g��P�����?������O�P=�a��x�~j/�I�rf��$�M�aXu�`~���m����2�ҳ	��چRy
ɼs/�C�>��\j���������9�=-fTY��~̕E�&��C���%I�޻�I����
��M2{�,��d�+%0��3�T��$Է�y0�Al��y�Cg��+���[�A�r��9�/��-��� X�ج�+0ϐ�_�9L2a?3�q��L��ŕ?=d���s�Z�a]�Y0�3�a0��l?Xe�aP��N^��!Y�J�~��dW�k��nm�){�^7����]�����(e�Rx��p���?!�cI��a ����N0�8�l����,��~|�\be �I�l�Ɛ_0�J�3�C�+=�&e��B��}��� � V>C��%���?���0+���e9J�Y�w�`4��TU�_{Y�J�W=���oT�Cg�����&SNR{�0ͲcO��Ԃ�$ۄ��p�$Pٛ��8��Ƚ��xN�"B�$&n�PF���?O��U�+� ��@���r5������7{("UW�Q�]��Zu��䶊Sf�\����H�u�8���U^5xdܥ��j�SS�������|��s��jR��� (�a*5'�i'�V�M�/U�CL��i���̗G}��2Tw�bM��2T����'�f2l��rm��0ɝ\����|�_��v������9�>��w/1��{J�Y��3C/�L"�����Շ��e8['�5l룖a�@Qd��gX�Y�8�������k�}�O�q���?z�	������Xu�p�dƷ��sN��}԰�Cߖk'e��o���>� #�ҋ'��I��T>M��'~�+>a��,�
�����8ɔP����`��O3��+��g\0>k2�ɆeE?P0̰�a��q��$i8sa-�L����c�)��z���Ͻ�fO̬�6L3g��E&������4��*M'��e��>a]憐ۤ���ؓ,<ʪ�[�S,��Ra���|�Xa���2�����P��6u��߳k�+�W"~��ǽ�d���gH�m&����$��H/笘Vv�~=�] a+?'���&�P4�/s����u
�L��2�J��a�Z�0��dgY* ΤR�>��S]�v(fv���+>l�&P��O�v����0��N���;H,������ɴR?<g^0�aMc��~`\�q:��1���ݥ�ب,���³,P��y���%�J��?O�;A�_��?!��`�<����	��L0���,<¿��7�`�O��|�����	���(�����P�E3��=*�p�n��>U��Ƿ���K;�)��/��P�F��x�(�}�О����;]���b�&"�.:��r��3gN�p6���"k�h����U�N��">ޛ�þ��@��NRF��g�����0�d�ׇ��U�K�c!�;=��p��Վ�=gչ-�'&Ĉ�Ų�ty�>Y;p��N�Й�t��3��8P�V���R�r�R���A�Bu�؆d��M�2��=C%efp��_ëmr��I�n�r�ZL�Aϫ.���ʬl|kmcy�y������s����ŪK#��m;��W�@yr�i����(��¶�QY\#͘��=I^�-�_C�3���=�i�q/u,�8�F���R`�P,h�:)����,�2Jp}��"NHQ��p�s�a��v�5خ2@�~�Z�������s#o�����C�A�A�H�}^����em��⊭.a�>�`�s�v8:�;��;�]b��qD��:r2K�
n�y{R��r�����)�4w���me�G{�߬��8
0��
͖Ƿ��	�*^NC|��8��pFz_���ܱ4Xd`ޟ�d�rl��S���͊�VU]��\r��١���.&��a�����H�3xD��F'����9�:"��2��8���a����ެ��9c��%�]�W�KM�5Fґj]d{Cw���#ᢒ僆|}.}>)zOT[������&7�dm^J��y5�a��(zk�sAc��� ^�u���]�a�?hu�_
xս���};u���{ʇ�'�B��N�*#{G�iR�%�|w�Z��.�KK|�i�4@qr8+k!u-��,�9�� خ��!�P�:�!ᝊ�E�Sۡhgh�W�5
�L�����fg7 Ī�M���C:��V\���o �xA�o-�\�7��[�
�'o ��ȝ�b��r��7!i�~��� 9�����Ȓ�}愇@L��t)��>����x?ἵ���Oz}3U�沍k%�<1�\��EN�0k˘(0���z���dLR*��[t+���������Xb^�I�^��ε	Nd��6�>�����G�|o�c"�J�xR�-���!wb���u�����T}��[xV�+��~�;6�(�k�㎣�9d�y�d���h�1W������8۷<qt�חE:=�g����Ϛ��:�ŷ8 ;�:�
���(ٮ�ECڶeU��a����U]�2�ma�-��/Uz�lR;b�w��c9Fa���aX|� ��)�B���ε܋ݢb�ޮL���P�U��D����T�2���	��yr5���o��t.M������S��gx��Lg����s���+�3f�V��|еS��@F���+��o	���u�,��ɪ-9�5� ��5?���<m%��T2r߫�ׅ�*�h�`(�w�n����Ώ�~܀�T�#�>���a��C�#ck��8��qG�V��X���x*y�<�&WH�m�>~�~�bm��C�Bc2�J�jX�wjR�iТ�h����h���Gnf�+�]�ZĎZ��QЫ�v߲y�������o0u`�Ŏ�8�u�=�#��[��S]�����h)`���iV��i�������l:ډ޿� x:��HU��ڭ#�����'fذ�H��O�Z�P�"�+(}����=)���1�����J.�2���8� ��FFr}|/��c���q0n8v�xrYZ�|�(5O�R����<5B�3��~� �@~c`车�>��~5]���u;e�I���|r�|��oY����5C���`�$ih�����2�"��S*��\�dGӻ����ۮ� "�lZ8�[9ht0�J��-O�
jw ƹP�c�-�¸��{�hRO�Xe��y����&©�J��yh7=uI�U}���8=���]��ϖ��ٱzn�O�r�ţ�:+Q���9�.L �MY�m���ݼyDaf�.��܆	|}C�7���N�n�:M�*X휁��T Beİt�;Y�X�,�����g��������GS��� ���:+L��G�o�4{�n!��2<�r�{J{�Y�kw��lLܔX=��z:fԉ��;�a�Kt6��GD8vtr�pa2�|_��=��]���=��+=�D��:!s��>i����l��6��O�e�Q�U������lu�9��s���^�OcۧƢ5;RD;�e���\ZU	��v6����cұqK�Uq��^\T�;�SN�V^����e��4S���n��CWp�y���V.���M����wfbO���V�7}|r�l�J�W%�q�k|3r�kf��a��|��Q���
�d�O:�uoL���������*/�}�v��Uơ,,T�z��\j��`��9�S������#�+�j�[��t��دt�������t:"�Cw�Z?X���kd���
!�&��6x�0�@��Os�y�FwN����:�ժ�������_q�����n�WR��]���]O��t`E&��{�5��e�h��*ˮ'F����aU�v��gZe����7\���w4�Ky�� [�Ӌ���/OsV���9���֎�ZuB�-妄��F�h��T.�J=����%�y:
j) ��������j�����T~\tr�௵��ci=�a��E�dg
I�SM�b�;Gabј�m��Zn��Oj�[d���)�Ҡ�)�ɓ,�s��E���;u���0����޵�G^ڱ�ۢ��:���mz�Z�T���e2;��j�Y9"z0�ڼ�!�jtD��M�\���v���K2���W�%u�Pj���`���/�=L{X��'l؋��{rr��2�]�F@ �}�sqR�����MJD�n-Ao�R$*���41���]�ǲ)1m��ϔ���j�T:��6�вXB���Q������xЮSu[��SUJ`����ˏ�1Y"[O:�H_Z�.t�����P�4
ʹ�()L���T��t �#إ��n�oBћwv��d��`�l�1{Y9���!��о}�c����9�A�����g dQ��]P�N_�/6��DØ��q�OH�/	~�F���Aд]�F��g����P#�k#M�U�r�91�Yb'�P��Kw@%:vK\�%���b[B͋7��Lܘ�ЙKl��j��i��M�z)Kt���	7{��
�Xn��H��)�>��o^�u;�b;w$�w����t�J�Y}��;QbR��˒Sa:�A�E9|N�5Gj�Asf�\��5a�W��M���Υ�E-V	4�[�V.o%m=476���v�Z�je
�}D��bvZp�,19۫YV���������<Lq[�$��R�QɂPӪ]tɁU����}�R�p+�[�-�]���8��@�9g�����"�8�;���X���n��g3Rɵ�f2���nkPFm@�c�RT�P�f�X�5&B�b㲓zc�5r٨:��bc/��m��Q|z�j��Ш�c�ٯ6�)R��<2eػrM��0�[B[qj�>��}(�o4K���m� Ӣ�j����S��]�3tX;�q<�U��X��A`���X��Qb��F,dTp�Ȃ�(�"������A"�1TTX�b��X*�UUUb���b(�"��"�"�DQH�
�����*(�DDQH�Ȩ�X������� (Ċ��TE�k"""����*��"��F#E��"�����DX�����Tb�DA���X��*(�"�"1�ETQTb��A��B(��*�p�QX���EV"��0U"T�TAX��j��X�H�"��E���"DD���X+Ъ�Q�UTb��ED�*��
�,dX�Ub1b���,V
���*�X*,T(�$`�,Q�X�Ȣ��DAlQETR0b�!?��Df<Þ�7���ͼ��lp`�hT��pJ���o튻�-��`^^�פ'�� 9��a��bI��r�]D%�|����75��YJ�'�sw(-�U��
u�����G�|/�Fڛ�������Á�NY��2��G����]��t4:�:�9>��O�9<($���&���,;qaG�&���WlCH�e���'ڤ�v�����7=^��
��=C����1^�F��
a(ȸ9�K�Nc-d[S̠�s<����A��lc�j�Y�$����C}�������Ŏж�wy�43�2�������]�g�9�<;��}췈�^�`�C��u�!Du��P�WtOtSd'8����nr����:�#���6�G�;W��|v�A�g�M>��b:��T-'F%8�;��;`%Fȥh@h?Y����#GEՄd1��s��SZo-)����ϥ`˭��t��* �����_<GB~&�����ŧ���t���w�u
��U���ͬɈ��lޚ�z��y�j#,�Tc7u��56!_�uT8İ-�
wo����wk����5���}�C�������r1�M��6�����ObU�f�7��N^�.h�3yc��AO<�kH8s��&�E�=��M\���%����4t5�[���κ��8�d��]}�.�`ek��RG��ل�f�q��Rҥ���u#��2U�Q�y �Qֹ�{�M��^9�]�2�{�� z��X�%�ۙ��:����>��C��3�qz4u��ߴV�ct2R=�'2�.X�7�zbf,,h�F����^��B�Ð�ׯ�
{_=���ǲ�Pwa/#Ŝ�3�&�D�ﳵ���N�Ŭ���ޜ�\�hq��ݤ����]N'�#l^�5iF�o �y�X�ךj�!Bhs���Ƽ+(X�xGFY�s��K7RRO��K�[�L]~9�oh�NT\�����70!D2	��Q��_C�3��.��s�zejx��O1����h�݉���kb�9�ʇ��,4�4J�3>�^ژ,��NPP��(f�9i�!r�8�A�5֣��|�F�ˎ�Q�J�8������s�4)Z1���ks�v�SQ���Pf;�^*�Y��]v�у�~X�x�X���I��	��r2KX���Q�e75z}��)Q�xm�"h�zxo��j���߄T!}�!��u]��J'{�SS��K�����o⋩���,�y9>S��N�dhÐAy-����.���%<���t_M�Ѭ�[�M�r懓	%����X�d��}��1�Z���T��O� yv��B�c�p�q�R�2���z���8��Hqg&u2�m��������,.9��⎃�Y�K)�|:*w�xh�}s��܂r���(��:o�{�{ݜ��A,k㰨�>��V��dLo�ͣ��{jZ�!�zxZ�rө�	���Zq��_���{��9z��=ʟ/;{�v�p�E���Є�׏�R�;��A3�q�X����۩���i0�)
(q	��Lɹ,��b�W�	�J�?�{�5^�B��k�t�<�)��z������`ߔ�i\�z��ƕ�-Kӱ1�df$js��Gs�7yx���r��fz� �@��]
f�O�E�r7�6�Q~S�аquY�9��]Ʀu�솼p�"�v�t�}��`ZO�j�҃�\(%�����7b�b����[��.P#Цn��xM�+��><�����#�(�&��A
~=qp`eh�B�f�]��ln*����Td]9�r�yG{��`�ydE���s̃pr/��>�����އ[4�����k!�ȄZ;ǣ�ܹ踯Jt:,78 ;�*�@�`��T!)oC�M��������oJ��{ܾT0t7(^�Ql�3(��M�AO����XT_.1�O.��̚�J���Qu[c�^���gL��ˡn�^w����q������1P�i����(5���������c�Ż��$�v
��-[<��u�+��{�r�U�k9�nd5!�X�ɵr`Af�7�VW�8��[Yw]�����/k��^,V��-uu9�M��{kKq�0vHU���ݽ��+λ=\���Z�]�m�b�f��Eک��/�a2��|�WU%:w+X)j�ӌ2k��!�ѥ�˜t?R�Zϙ�ŉd9��ey�E�J{V��.�[[��b��a�����N3~.�Ѵ?g�
�]�5�v�0k^.<vug�����S�#�aĨ�L+�5Gg�B�)F^[���N�>��s�[��a��[���y�[�t��z��Γ�|�h0��yۂ\��b�:�"+�����Q�~��I$���T���T������z5��ɹ��돊�s��_{�;�{q�������W	;�e{l�뚮��"�)�=�bx���\y%>E�de!1L�Tpb��.քuEeE�	[��pH�@�E	�h�R�p0i�<�)�f{��n�"]��I[h�K`�˽y{_a�F���ϣ��=@ұ�'���*)��:��ڳu�����@�+#z�0�=*,;T��j��_	^:'����g3����qe�h[�A�lF_6���l�:B�n��ԇC��]�n;�.���^�vX���E�;�ti5�J[]@���·w������P51�n�vG�Ӡ�t*���xx{�g3v�Fv�ب�*>�ܧӁ9p�G@��1�W�۫s6�ц,r��h�F�gD#�\�b�Vt��.��S>�ң�ll'N�:J}*6;N@�0BeİkFNFP:�����:��'�����_����3G�hВ�b4�w�F�˕&�Oo���h��j���f2m�鏸g+de{W�u����0���ClA
Έp��)\�[�ʉ�h�`,�����p�0^��|�@E9��4q�K�,�oΌ�)�Uxn�_�>d��TQ�4`��<[s2[��9�H���'oȪ��$�N7I۱�ϖ�߻Y܄"=y���f>nѶ"�D�I����L7�9y^Nx��{��|�:c�q�C��<��`sN�Z�{��T�GhZO�S[�F��X���ױ��`N�F��uM��	� �
:ͩ��A��q���X(�/��@����3��7�5��5��뼬|����%W��"�K7�6�����o�M��éi��$Qs�#a�����?�����������13��wi_�3j�>��'̋R�"[f��������U�������r���
R��ݭ.���z�[�.��/-<���3�h��4K�ʙ����ܜD��R��i��]��N�57�N#�]˕]lle��殺�{��5�gu��Wd��E�J	]��}��_Uty��&�aOd�t�*E���F'���g��JU�U�Cc�h��x���ec�V��jw��x3�E�T�lm��<��<��<����H4���|�`>������{��CϭK�(�▍���V�Q���)X�6��n�ר#<Th���D�25	R��ij:j�F?��R���r��ƣ簨t}��V���r2P*z'y�qq8�SK�ڱ��\��B}Dr{v-\�j(Y�!ƫF�:�Ec譎��dy\ɸ��Φ}�ם7 �/]BN��9��YQ0�T.��QW���Zy�a�(��f##hN`m��,�a[MV�&��d������7O�Z�=m1=�p�/쮯]�hY�
����/.e;o_Tj�0��gr��[G��!\)0���p26ʍ�o
��p�T9lS��]��.��=>Pȼ�CpY��yd���K8kz{\`gz�sC ���5��w��Z������mT�R9�b�j�;=��r���K�/���a%pf}
�Ʋ&��z�U�$�T�;Y�����96�q�L�D4C�p�L��.�s�ҞR:�v�x� Eaä�[��Qm �<���4gK�9�����Z��n�f;�UVmjW��"5�����Ff�{7T��������tgrۡ*��@��{��/q��U�Yc��3<��#B�����<hH���yX���%���>�O/�u�>����
t���?������V�8�����fȸb+ÔI��	���O'{�����{�#g�������$��0miad�����}u9��E����+鋳���߻Û�s(��E���D!@9(������bY=e�X����Y��:�%��������*z�ݲӾ��p'Ov*�hN�H����F:�Wك�Y�/Y��N �wJ_�4&%L���J2��S̮3��"Ժ��uu�P� �F�&5�׮=(����o�Ӛ7[YE�sp��&(b����&v��p�,V�#$󍑸�c"�nzU���v `�u���vw�o�<k�"=������B{�o�������(�� �y�b�j2Z�q��g6��J�L��ж����ZE��	^�=#�q�?����3ƸNZ�u��5�ō?A^�f�E^�6�v���ɘ^��F*9C<�f0<���Tv�����P���h���yY)
�Z���	��Tyv&i
R��w�1�α�շ��`Uiu �r��	�*�>]���ǃ?*�^�?_�GG�����sW��W�3��n]�kx�'2��iVY��b�d���a3�u:��-�h5-R���z;x�[�5�p)9�7�w��������#�o!�i�w
�����~����ڕG���#�>��t-`�!OǡcF�Ζ��*;Y��k=֌Q�wUL8 �ϖÛ	ߔV����H���� Ѓ�xu�f:�%�h)�#+�����~�gb5K��t�9JB������ �� �ڔ�]����P����x{\�l�k�+`Xu�_*:��z�τ�穀<�|Gti�=�*K�V��s�9頋�GM���)c�D{��G�mU~]��
C�{�c�ɢMgsCB��LV�;E���,e�1S��x�0K����^pu������Hj���8��)�ϊd�r�Lld{�o�cՙ�!q�!��Ѿszi}���>�:�eV�CӃ#�2v,m�>n毇=���M�{ǈ� ���k��`�9��{�g�!��C���%YS!^���-��⚹S��ܾ~�v|�Y����*��=Cg<>,Iٶ,v�֟�����i�ƃ������9�xbH�峱P��e#~�x�*uqp�>��k��#I�*��9��� ^dwOo����T8ڢ�Ez�H'V_<V�1�t�7�J��v<�4v��2���=V@��^��N�p�r��t{���`���Yz���֥��Ӵ�Z��&B^P��sU��R��|�gUޜ�%��yy;��[�X4`����|�n����~���~�����K�t�A�.<�iᦸ��3WIO�Mu&m�Q��9��A�Jh�]�a��R��9ĝ5_��i
#���'#|��7�{4�@.�R=�q���v�$�{�^��5y���{���>|: �IX��|�<�>���^܀�bUh��x{){{6�T�]=�Nzy�L�eB�W/9Hq��[��s�*�"m�f��YS-��D�~���k�U�ˏE�zF>��p՗(�0�d
��uhI1�8�T�Ҥ:�@���mK�sp"1�_��#cѱ���n�:M����q\v��0A���zQSGy�Q/��'�u�k�%�]`ߣz��'��lԔp��;�u3<4�ǥ���=�5N��|O]���pqy��{_��qm�H�a��N�`�=�}�?W-�W�&^�ַ�X�Ja	���*(��%眸�0+��ʄ��.w������l����:�vQ=�'��t7(�u��we���x��a�,�=4vm̦C�X\���fu>��^�r��Wr�X7C�<��z��8x�yo��Ձ����]�����e,�>�8 �a��ܠ�v��//rj�Lb�r�-�(�+����J�������&��Vt�R`tOR<qeY�Z�o�%=��;t�ͧ�8�Sj�l������缍Zw[�/�l�ȭ��~�+�����'���玈f�gi�W�:��
���3�Fkl��R^�4��z��%�v9�b�(:�������@���6w�fR}���9^��)o�Z��sx�#WT	
{��l�?Q��.���Oz`�}C�}͏�V>}���2����{jvx,[;i�ת�V|�8��`Y"�7ƒ6yV�;~�+�Ce㧥��0�Tھ�y��e�gCnF���d�/�aZ��i�;�Xw�E�+BA��#��Ĉ�3X�Z�T��R;���i�°	\���ë�9��a��1^M��u�«�h��y��/�8�p�b�N�Ei�q0��F�Mϫ|�B�7*&�����:�H�5�B�P��v�X&6�Z�P�.�dF�uP�"�����W�f���C���u�7���*z'��q�v6�*g3�\$0�;1��+�z��	*�]�Ѩ���!ƥ�З�g���`�d�׀g�k�⻓�l`ٖ/��("�ʧo�c6(Օ(��z�V��a5n����D����U�L�Z�U�AW�`֪���sx܉ҥ]�;x(/��!��Sf�����V�+4ժ�<m��Ci���e��Y�;^��{��a�/�H�ڒѻX��\Y��L+v"H5@j�&�J��F��7۳6���P��랻/ZW
��%���@�j^���� �W�鼹S�Z����!�����d�f��b�����"r���F2�Azn�$.�N	����G]�C��6����4�)c�S	<������6��8^�lx/��3,�[�3�;��FsU<#�\��e�Q5f�,���2��3�"���#KI̗�"���� I�ܮ��r�bԀ��0�;���$�>{]2!����,��}v��=i�mJ�� �vV��N�z��ոޜ$4-�so�jq��>FLe��U�a��iy���a�z8���d5�`��劵;G �h=7G�k�2��	cM8E>��GpI`��Z��K�s�����c/p]9�c�[N�녕�bz��w��i=m霯���ִj3�nk�+e�Q~Qyԫ෺���V݀D�AԮoj��7��v�|�R��y�ꆷzo�m)9:Pp�N�v��6�LޅX���*RczA|d]溸�iq�rh^c�:�(�>��EE�����b���C7'ۆN�I�vA�W^�էqj�
��s|8'I�V^@t�T �6�1[DwY"�m^���.�^�q�əܨ�a��+�4������η\�7�t�2�v�fúN����E.�ޥw�6K@�gM�;�I�{3_.�G�5h��NL�o��h�HF�z^���-nG5\6*F��r���=w�ҷq:�BU����q��{v_!�`��}�;�����u�1n��.ݡ�x�N_�kiVS��s%f�3�bh"���E�N�j���euf��8a�adC}��;�@�'Xk�;�V�BaB[y���8�\�7,�nH�s�ckF�Rw�6g%&֦o�ĳKXw}�7{�"�4�j�B�6����C����SPB7���:���;��)������j}�7F� ۚ�7���P�{��t�HА�sD�����|a��ݟ��Њ=Rd��)�]�;9fi�K����-�%rz��x����k��6K��� tU>��덮��l�h��|�Τt�:�5pv<'3P)�m�`R��0m��H7���=U�����3V�س�� �霩��b($�TX�kW�1�rx�0S��Ć,�̺uA<b�&q��rJ�YrĘ37�а��nQ����� ��n�=��ZR�$�R\Olyl���D�(�\���ݤQ&jA��=o��n�,��O�NiJge�X[�R�W�f�>YX�_P<��:H���v�*�.��Y;k����~~1���S(���b1DPv����5�F"#S4�������UE�X�����"�"���TH�B�b �ekUQQX�Tb0UUE�QTUTTX��hX����Ub���APc,��b*�0b*�����0E��	�Va��Ȋ��#f-��UQUU`�jT���X�V`����AUX��\\&*��T�`�Q�b�`�(�QG+X �����Ա)���",F*�b(�EDQAR�Uk(�",X���6�Ecq�"#Zb�m�U0�eUU��"%�+Q��Ŋ�V�1J"+"4Q,F*"EQPJ�TER1A\[�TF"���G",X��U���
*
ZX��}_�\����ohY]���٭ࡷ�vM�o\冠�� �7s�)�H'B�N�뿃��-�&�S��i�T�}_UW�e�~���.��g_-��fx�!�&=��x�z�'����]�I��_����3�F�&%n�ぼX��D�������"YTaX�p+N�¢�F��&y�y��S��d��^>������4E��D��S)ۆy��8��d&s�FNF#f8����s�^jY(%
�%�����a��|���<k�H�*�,�*h�~f}
���D5�v�dν�=�Ɋ9<N�<
~g�����.���^�����Ta����8�]]�5jTm闃������R�NeT�"p���tU��)�+�U��a�V5�/�b9A02k1d��O+�/���e\]zr��}G��=�pp�K4�G���qX���� %��7�1s��ǡ��YV$CKr�����AnW���R"5ز�*���ig�(<%�����9U�8�;!���k`M�7R6��,@�ev;�ZuzE�|D��F'�3^��a�ŋ�ӁB�U���9x��[��tE��;B-r��ڨ���A�+������`dtJ'aF'DՈn���>�T��spwe�8�K.x �4�vȨv��z���3w	 XL4΅��ne^���Ҫ���e�H�7G�]0�� _]|˔��B�藀���
�cg:���ġO�z�[�����e��&!�7/pq��*�%�Mҭ��o�L�1~����ҧ��y�G���f������c����;}7
��Z��y���N�DM��s-�E�Ԝ��ҹOŘ�?p^�zl�R�G�/�SF���
��T�e���p]����7k�3��z��5��h�;h�[Tl�D�6��jum�����4��9yO��������͞�V>��o��h(�Ʈ>_AҾ4��Ңcq�8��R���TE���$�\�����ѤZ8��mu(�1�t�^*�%˓tȚ�����$S*k�gc�4��hp�d��Zj�N�1z��S�yN���v}j�����>�~��A*Lgc���x���!{����@�Y>RF��Ge3�y��44�AM�!���:���M)Fpe-����ln�\��GA���Q`��P��h�B����n}CJ�� �yʐ�(�0w=#Y�p����Goy�v}e�#��})JX�S��xʲ��P�8��5��o$��v�+F	M�l>үO�'Y�]���������犴V��~���B�[*ijzL70#��wb:�Y�.I+�M$�&ŲA��9�b�k$��1ßz�����Խ<2n����R��]��EO����mh���1�(<5pf�yCQG��`��k/0���|�rw��ٜ�Yb�.�z��9��{~.�Z$��y�HK��-h�(���S�f�\�`Wv���v�yZ0�9������Έ�
<�t�ѱ�oM""E;�y�M�c�Ku��0��$FI�y�w��ܷ1�W�Ҡ#�y)�^�Y(þ6>~�q3��5�c�i���1)�����#�.��䆹�z�g!���y}�:���y�!���m��$��d�ldUR�	7��b��O�9U�m`�jV��-S��s�+��ָ�j�(�ٳ����3֯�M�wﷳ����e��p�"[��9�c�K�2��H}�ā1�t^�u[��.�����5��~u{�d��Px�c��Ч�m��B=��&��%{=tM�6+��z�3㺟�8���ͳi˅%�zFx:���c����]!%iD�����jc�/���G;b����r�d�AaJ�"��(�l9�s�Cu��9Hq��[��s����Q�idk��(�}SZˣ�����O�.*(]�}8��q~G�tP�+�~n��r��xdlRn�{v����OaZ�s�5&�X&�N��gQ���N�tt��s�r��q�>~��%>xeK\Oھ2s9V4�vp�4[�y��ɭKOf.K�&��)�(��<�*�]֣�9�32*���.��s��<�f��t��eU'v���v%�$�EJHֈ�� 괺�b˩�?qؾ�{��q�Y��^�A��a�~�;�n��e���Rz��MÑ.��
X��C	����d`�����({_��1m�]2!�N��f��2��~�h�f��Rڮ�����W}e�"��EƗ��%`n�
��Ʊ�Y;�lz��>�4��Q�I����t���zM�x�E�89��pe��w#Y�H� �d�p��p��Dv)鑔J�׍ԩ���C��{Ϸ@���a�	���eT�N��"��jr��8ۉn�n���r{�Pz���P������w�>���^k1�d'��^���).�w��o������ɯ3v�B�y؟k���Q�_	��=X(�H�O�t��t�W�os��+T��h�X��
��
��L�FP��@vٝ����0�^�p%\`),�o!"3O ��XL�b��W�g�6�m�Ŋ+U�
��7�#h���8�{|HH�p��4�@�"Y���N�Ʒ9'&i�5}��j�N�Ϫ���BHym�#ϓ Z�3���v���F��]� ^>��e��s�w�A�֪��E\܊S�_�PxϞJS��3x���e�h�y빏H���T��ށv�P=��\�2��5�d�ĳ��=�O �D@��k����^ŋ�&FE�w}_������Es1������A���E�����F٠��]�9P���t#M��<�DNʗi�-[΋�զ�\X�ɩL߫���d��iҎ�����n>�8�����wK§
G�t�n�'����3xC3��H-�yM�_gĪҹ��F�8X�[�S5�{�h��O��1�]����;of'�A7�;��]A����iO�����B�P�ru��'����p7h�7]B9v~�}�ԓ0�)����UHf�7�i��у���/Uۡ%Ky��F��ic����O��������\`�D�j�Q�l�p+�v�gAC�����쾛:~W�2[�'�..nKd])蹺OCٱ�6��]
\�w���D'�]�{w8�Ԏ�,z���лD{��B{U�0߯j�H��݊�x��M)Uٽ�SWŵͬ޻3��Ę�"k�Ya��&��y>�>�&$[��pA�a)0�o���f��V>������<�<�Fl]}>� �>����[���a�c^�s�Lz����B↾K�yЭ��x�����~�q[����d�c��w��9A���^�=x�lmV�z�m��O���4��Z��+9!ԤGX�E ���}��5���WThb�6�C�[�O���NM�gqf&w;��ɽJ�y�t�.U�⧆��D�+�n���y��~�%a7�/�W�P��0q�����;��ж��/Q���Ҳ؝XnBm:޸�F�U��z���L�����r3��rΣ�:j>+�[<��fܾީ�Hẞ�P��1�en�����yBb��h���k���+S3���������?�+w�VR����9c��P6܋�N�=m�^��G�="�5YZk�ܙ�˨�u���3�o�j�.W�Q��Bglt��.޳s�e7̦�Wo��-�ij):��r@Ǿ��x|>аt���5(?��D��h5MK+�T��b�U��t���9��;��|����Qc&yhC���!p!T��)`��l�>�J��qF����+*�L'�":��[
|��-)��9(#H���B�}p��LW�DƸ��Y%L�y�b������)�Ttd�J���f��q'N��1�>�WJM�ta�G"j2v������ˤ�Ì��>�v�3�s�W��q<v�^�z�2�k�"8,�!���.�m����k������Ea:��Ey\�w3�SH�"��+�}�y�Y��/e��. 泀�b��;>n�R���x�,wh�S���3Aw��&m�{�p�:�j[�N��jZ �����%}O�,�F��T�o[�S;mPXT���q��W}�Ƥ�w���	g�z��<�,����͎��w��+��;ްG*,\=�����J��x{t⣧���]���2!�Z�󡃠f�z��N=k�r��O��ɜ(�;$�����VUd��paX����c.�`��w��-�H�{��>���c�V�Yň3�^����q7|���'�����������9I��+��,X�@���^�Vbf��5��9�lEl�^�.���Uǵ<fo)�����+�~���c�!�I��ԙ��NW*u'�U�Yȩ�P�y-ܲ����z��˚64p���v4t�$un�+t������~�Űϝ�ˬx'Jƅ�U���V�=[s�O�νa�z�;���� LS�z���ZI�Ʋ���]��;��XlQ	�]�d!Ip9��|��k{I�,l�j�<zΎ�֮�@�y�z��(������g��2@i���к��z;��
�b6��Ǜy��S���r���>���GD��-#B�㇠�v��[Ci*����dm�Z�\ǝ��J�pwv[��_�٣��Ů�f���;�25���dN<�t��u�q�h���s�r�<�v�?]�uX�V���Zf���u]M+o��՝����>�3��r��9�;v6���l�сI锏oqpڏ=��Z�]!��M�]~���O���Z�W��a��W���z�lo��0��G.�]V
e�����\㞪��c�Ã7-9:�(
�]���n���ޖ�;Ɛ��5����_��K�[�Yk:��"�w���r���i��m�Ըp����O���s9P�"�ha���_wF�u7�;�@k4U�d�)p��|vTz�9�o�66�w��m5N2e�r��v���a�UlT
["1����7����v(���T�H�c�����5�� ��'����^��CN����,�z��Sz�!�##�*�Q�p����̓^�6��	�`֛V�u{>�y���	��AP�߹H�4
e���%cwp`W���ؓ*+�@��kf8�j��I�o)�,t�^���n�69D�4�׺�c���ʫ�`DƢ;�NV�ߧ�=����;$�L{V.T˹�%�x���Y�ǹ�O+�u]Q��guI��q^���[VfD�u���9Cl�Ptq��b�C5�<^-�hޞgm��*��w���W&��Qҍ���9��$�b���]>�vU��}A[���2�w�!)]I�����ư�K�X�Q$��K���nuYx;�lLj��jg*���I
�����C�V����v�e�4��KE��+�m��%����.}�����a�_�#�-��~�g��.����V^5��䇆'�\9�Pm�iz�_n�n������2���V|�?�-:������G�2%9�5 �y��J�e=�9:w��n�ʼ�#i�B���[y܍�o�d]}�ͅ�+��x�cm&,S�j��t5=7~�z(4�P5@��#��U��E�\�%�J�ڧcc[�����7^���ľ+��Czr�57�����P6�`��TW�a568�5��z��ʅ�n+���j�7}��K쩥�͜�م�a�qq`MM�v+��X�
=iʎ�������g�8�|����"�Dcyy�(�&�������m����+�BX�WP�h�?!S��Ez�._/]���2�:�{�"��ڊ�x�a"�#�!J�q�c8"l���b�[���de�\/QG�ɝn^Dr�:�f;w�`3Ԣ�3�i�1�1�#��4#'p��K�W�g��L�r�]�1����r}/�R�~Ξ���t�ۧ���M�!�"YTa[2
�dnK~{Q;&vL��`�N/H�m^��dyi���oR�T�c*�ɖGt��Zل��8���}��A)�Y�ws�����ы �BɎVz�U!�w^Э�C�)�����&ज़�w8���6.K�V��j]�0��= ��	:�cf�qk*��ϖ܄����n8����Y��؃�}^ܖ��S�sb�����G�6��4�*�*�e���oZʽօ�1�X���>1�h���:!�;AC��T�<d8��E� �[�w3E/r����mQ�v��W��sDgN��8��3��G�*Zf��]���<hI^>��?yjft��[�ƍ���}cSz늕�^����e3N������4xgӰW���%�W]�!Fa��X��E�a���f41�,�{}�o�(��n�^���E��2���냵�a�B�!�w@�J�0���N�WoƬc�o�@��Znx�T�h��܎��S�����
㞁,ϕ��P��4�fo$T=9�5�������}�Ǭ��#��6��}z�p��q�(v��U'��0}=�s�8��>�m�����:b���WX�^?����E�����#{�ڙ�%��{�r4��M��>��2���=��:�A�+ƴ6:l�i�@���������s?f��[xgƌr�KW����6�i�4���5
��ۥV��|�R��]�i�β�N�:�[���h�.e����o�#C+.����J������Ïi����L4�$��@-KM�@��|�F+�d�k�tJ�'P�鴲��9��>n���p�-���Q=�3���a�gu
�[���[�{��5���������УtQ��<��Xyj��qFU�<c2�ݰ��WT�|������[���>瓯cC$ܧ m�;7��&"�5w��i`�6$�7�."=li(�@��/!Q�N�#Hg�w��u}��d�T>��V`��^S�QK����"f��aX^��a�:�7��8���ݛ��Ѥ]4/ڦ77��9�흧�6;���/��� v�9˧ntѠ�E���3{
��d`pd�����J�P8ȕy�	��l3�mq]w����ΗS��]�����;�w�d�F��������fg�>U�z�*�s"��.�,Q֩�����kw�x��|�n=��w�f��
`�"zG�!��2��p�D���pm�Ӽ�	]o���WFPc-�����7!F���:�#3�ᴪNe��q���e���\@�N��%_��:��+���`��� TkFα|uW$D5�oC�,��[��I�!�*V��#�[M�uK�+tD(��/��5m���u�S�{�v��Z���փ��X�v�2k6�7v�K�(�jp��P��L׋l꿕��p��q���A8��ʴ���[ƞὄ(M["��aMӊ�]Ӻ|�vLڕ�CТT� �Y'�-+W��bu>�<Tѵ۵��2'��(�'�R�m����I��򠷕RL���c��e�1�"�q��M�Fo�v��Y�@��Cs5�p������|��޲�����͘H�F�Q˒%�KM�P.�	�D�j��%�F�E���wJc�]�:�dzʩiI�v���5qw0f���{��#l�� ���j�|�<z��l�Q5̸�X�]�ݯ�!�/-	Ҟ�K|9�Z�+�}ۼt�UJ��x(�L����[�[��l�B2LF�iIV��C�XĘ�s��rl��-2ŧX���ns#��W��@:�m5�w��VÑ�����6="�욬�mS�D-n��=}��}��c��֥
�^��T�s��E����*jna�ۭ��n�Ħ�r�s���%�$6+��ٛ>�dt�8�v�C|���O�:�F�*ᖨ�%;@����<n������B���Ȯ�X��r����ŝ�@��G�jڵ���T��	�̈�\�W���t��ӞuE�ͼL�-�4�f��2� �Farn�a�gl㣼3&��
�|F�`ev����P��Ny��Wr�7�l��!�{z�0l��� �mދ��@k��|�@�K9����gQ�6�
�s�$b�9s�5��Wt"2}�V��Q����+8Q���L�Jʋ>��p�������n�uv�ެ��j�|�@dj����;Oc1O��2!�ݮ[ʤw0�Q����' ��m.��r�
�j��"��6"
���UEQA���#�a,A`�X���"+"����(��,*���EeeEQE�UV�E�a
Q�1XVQ`�0T1J,TdUŤU`�(�b��� ��b�QEH���,X�,V�� �EQ�-�$J�U���Z�,KQ�iUU��l����k+"�"��؈���, ����QZ��b�T��,UYR��2"+,���DDE�h"�b���V

1b(��*
F+��V#YZ��TQEb+�T-(��TX�R��TF��PQU"�Q��ic���
��"+YUATW���_ܫ�qU8':�V�wx��Cm�w�5�D-ա�7��x/B'�w2�Ě�,�7��ʡ{oc�x���sPJ�m�š�q��/Fɑe�����`�z���kU��%� � %�U�.2wW]�67od�߶z�E��l��Q��	U�0�Ù��\D��U
g�>���0��.'[��7���B��S�г��V=wǼ��#G	�,b���/��iǦ_f/!b�����x��o2�給d�����'*��V�7�4��+���ta��9���B�BI�[T�V�ʁpH[�B3��|n��tB�ņ��'���ױ��5��J��P*{��ǰk|��������,�<aF���T�<����,���釣N?B�2n��noV0�5��CڶlW���l��W��S��>����-޹�v�C�B�8|����8J����;�J7��J){�ꅊ�i �3گ��)�s�Ww���ƽB��/x(=�*�@!��|3���^�����{A������j}��4�f{)���~[��ˮ�@�|���r��H���B��γ����� ��euS��5w�,-�i�y\��Y@�<�G���4Z6Ht"�V��=��uӣ�&30[0�.^J�Kl-]�̫
�Pt�,�u�a��LB�=�b<&K�_S��dK탡��ܻ�'>�������l�O�V/�y�:B�v^�WsyZ��܅�����k���ۅՇ�y}�:�Ǟ�z�|�J����J�W5	B��{���3�%6L��T6 !;��Xo�EBv2�.��4����et�@�H9�v�5���쭒�+����z��<�n�GDJ�c��_c\�
����>~[��⹊n�	ݏ��jRZ|r{�8>[�#γN򞄬֠�H1�!���8F�@��)�Z���[�
ؼ��[T�P�H�9�m�˅-��0:���N����d�b]�z=̕���mB{!�e��r��ԥ@P'!���n�ң��&�"�l��89Y�:DB�<���mA]�T��!���ԉ��EÇ���c�08��E��`�&u��P�W��娍�|<��^S�m�=��d�r{�3��?�3��W�#���ܚ���S쇎F��(VN�*���=�6��t,`\����n��m�l��1]R�mRu�pQv�����s�`zU���Qs<ek�5�g���e��x�p��R�hOu��=�5�z�XN��L�k���yR.�Ӻ���6X���<���un��3����r�]�������0��y1��$t\�Z�c��f�dP7�E:W��R�`ƻ1��d�FF�D��l۵����O���a�u_v4v"��O��yF&�SK����=�phˊ�yX"V����,��ؓ*+�㙣�]��0�;r��C^�ZI�����<F3�9:�
N�1~2��J�%x󂞳�J�a�v��;wa�/:'g�$�����g������C�1��Cux�N�]�N��hͳ�amYspI�pdV��Z,JG(u���u�?�{J��X});rŇ��M/΄��{c��8�ն�n�f���V�Qq���l��2�2q���AΫ/�k����)[K���A���U)mYg��~Bt�������Ҭ�jc�Ӥ�"��{�*r��.7¬޼�	Լ}X���#r�B��^e_���l`��z/!�xe���p����6���+x�޻e�cs��	90��4ˁ|e�+|����A�~�* ���h�79�=鷧�ՊZ�N�髨��Ǣ��-	��6� �I�ð�_*�,{ϝh[8y}~�݂�:�珟͌��t̡Ξ�=>�J=7Δ_\�+�n>�8�
1��I��/�L��&�;�#��i���38�J[b��i���[�����>��0��ɧ6[az�R��v�+w�b:���SQ����s���Bx���U�Ý��ĥi��)ɶ������{�9n���Y��fm�t��FRt�;f>�zDQ!���7s��Z����(*�Z6���B�D%�
�u����a�QB�q��&r����7���A[#
��1tV�779��=*��ӿMxAGJ���xD������f�\oۭd�k=n�����(�Gm�u܎׉�� nz�~��*/�X�2C��ʴ���aDn�������P�M�t��t��}^�����;$B�,�0�3!�O6�"�5j��@�={u����=�%�%���8���G���
/	�<��"I�\����Ul���3̺�.y�~���D���K��q��5+�ʔ�d8U��b*%�)�����(���Q���\WÝ"3�*��!i�gX@a�N[E�9�:��.2t"��O'����$��a��Q`�U�Y�SPy�Фl�+�@��kB��߭�1��R�e��Ǚ�nz�Yh�sq�+�$ĭ�b��"��)�:^z&j:Ꭱ��T`�P�2:��np/Ep��_��5�r<!X�f��:xDr�-�Q~�@g���(y7�ԣ��wi�4�t�� {���j�(�����r��R��&vn����T��}
��5j����ӥ���+��e�v��t�Ɲ.�쇛c�:�����S�]����e���95�M�V��m�թ6��b��S�ΐޣ[`d��.����p����Hc�Ӑ�dW���"�d�
�@�d+����w�}M
9ذ�8L��t��Ɯ�ol�����A�ǑZ��߯P
2+jZ;�f�CDJ�[{�<;4�d����
eE	�w}�[!�7L��?����Q�=7�)�hg������bfo��:��f>Zc���	S[�x��>�1�j��\6�0|~��+v�{����
�t��\�-��;����kF�`K��j9�*�%����BS;`��B��E��^l�W�!K�[�㨱��zzß?c�ZS���h�:Ga���/��;����Y���ǱHu��ع�����*xY�)�NTa�4�x�6�ir��+-8���v�TD��������P��tA�զ˨��NCY�~|i|kSZ�3�1�#ۄh��I�Jۙ8P�H|P�t_xU��x��[�h���ԧ�e>B������.s���^**U�����c�獲!�v���w��V�}y�b]��~���tp�t�.s�1�w��xu�dd��d4o$ʹYY4��`��U�Y~��	�ylg0͸t��<�v�37YI�y�*�cP�.\x6p:�ȴ���t�a��g1�x���A�Yx3��|7n��r;u���ź��"\5��O�k�c5�qlأ0�n�a[upVD�0�5�I[����+y,�ɩp�s7�N�Jw:��i��*�O�Vy�X���I�o}�9��/LW�}���l�&'����r���X~���h��1�������ڮ�i��o�����R�/��x;ӊ���b@�!{%�h�s7y7SF�M{�J���;�hI�D�����.�O�Y�-���^<�cBì���jcη�0����e�����|���}���VlS�Y8ƪ�N�P���5LwJ�HM��j�uҦ���}���{�IV ��wv;6ll����6��:|Y����[��hC�o����K�&A�.C���op���v���ϔ���q0s�>�/�F�\tVbT�P}����P�=u����ˁ�M��Տw�}@��@�wM"��6�����N@A���q*�oY������zg��� I����F\P� ��Cj(D!_�!����FyNL)�Z�S��P}���U��/r`s��n+#�!;�K�Hz�>�Z:��f=%��	�� RDg)�O���<;�s��/Eɦ��V���;Pa���5gko���]
��`զ�]k���Z�Z�ʰ��Nq!֤&��ٯ�^[T��������U&Db�ڃꅑ7��k�U�q�Ņ�:7+*���^֖flu�5[�a���R���  �EZ8(Ֆ�]\	7:�����O^s���贍�%��	��Ja�k�qi��l�b�
�\}��b�s ���kh]�[��[��&G�J�"�jJ�ܙ��6�	q��hS]�`����cR�c���0qm�^/�E�����e��r=�o���"��/m3V+�;\<6)�S.+��`�Y�����q�'iE
zi�R�,����*X��GC�mN�F�M��S>�9�Q7�s@c4 ��͝hI��pE�);��R�ۏ����
Ia}�V{��u]���#0�$�`���^��G,}�I�{[��=�
��e�|�xx"{�U��l�����ԃ2�3���#�F/�����VC��lu{��Կy�,J++���W)*�]r��(9�g�{FT������E˻�/yX�������뷈��v�<֍�Z� .�+��IK+�W�fݵbvX�[X�ܾy�k���
�A]	�^��e��X��u��+��M��=�<�)ڨs��D�5`��7.`Z�'�:ᓣ�7�s���]�w�bR�o
�G�X�q`��}��*��FT�F�;����w�h�����CQ�4�g��Sz�p꿼���?=��/-6��3|�j|�C�+�kҹ�:W�^���\�D�����A�c��鯋�|e�E�
�����㬃��1�f܅���oV���&%��;wBzTz�N��r�B����F�MϫC���Ήz�P�2��E�̷��GL4^ͤs,_U rS^��(y�hC�Δ_\�+�5}!G��Lf]��7U�e���r5*6R=�6���hW���ʅu{)�qxG"�<���[ї�1׮��T�x���td�[�g��Ƣ�;<�dP:���A�d�4T G�΋<�rsE��.�������:w�a����ئɈ��1�Ҡ�;eQ0�;՗0�qn'���ԔNܱfѯK�Un�f��fRT◫���.;���J�(Y'j%@�_K��K�ұG|x��/�w�c+�����*�wx1Qii��|_�*���{-��)gd&����F� F���7r�E�j�]��ul��:�(!�pW|�pî�S�Nƽ�%�;��P���S�xS��{BQ�X.��;G�l���oZ��oS��L��f��m��Wb�X��45��欲��7���-v��:�{�Չ���p�{Zִ��lv�kb�zK��{�>�J��IU��V4��,��$�[�f	�$��I<6v4�<(�7Fe��ىq����#����5��{7����U���D����:Dg�'MܮE�j�s��>B"6�x�K��6��7^x��0�tc`r74UrXF`�"x�}���0}f+��Ǆ�~t�y#���U'��{�9�x��t���ޠ��B��
5~�
Tu��h[	agK47���z\�]��-��T���*�f���s9��E�����e��^��C�'9�����wQ{�^�-�m�Ա����d\>dmxd�
�%�o>�S�S���e�����0��D�G=s��x�o���_B�k�ʧ�q�;;Q��Z9���+�+]^@��&&��A��Un4$�nvj<ڼ���kE��!����mꃪ���|k���Gm]����P�*Ɖ+R���WEÒ����*ؘ����\��h+�QbkX����ɴ#)T�7�31rQX���ȷs�v�8�f�mF5���#%N��Bs=����N�)����8�g+T�:��p�/��&�r68�!E���Y�רc�ZS��\/A�Q��B�SW��gEC����!��B���x��h�R���[�*�ج��Ru֐�d#���Ӧ�Mu��p�~�:�]Se3FrܝKB�V��m����u�T��Vw�t���m_=�x��Tu��!�뒧y;����3��0�N��*P(Y�)�	ʀ��1�s���Zs������"����ژFׁ���kq�
z`�eB���"��6z�W���=�@���!�ŵ��*o� �2.�yDE<�!B� �Ȥf`���Dj9:q�y�r2���3}�V6t���ѱ��5{ ��H�5��{V�
1d*Ɉȴ��_8�0��ܧ�ŵG2bt���}Jc9S.+��x°ۀ�����{�N7����<,�O����{�wPZ��L����`�gz�)�br�/�{K#��㾬��eج�C�5]pŘO-�.�՝�(�f,��k��O����uT4}˳\�o�è�h�S�1µ�_&�-�2|�yߟU�sʼ�ט��|�D@E1k�5���g#�=���{i�7؁ˊN&}ܬ��`�;Y'�g�nׇ������2+���&�j讻p�{�rI��\O��v�{�6��j�ة��[>u��U�����;ҭ����U��;�ݵm�Ǌ?f�dv?��|���:�q��ժ�c��@INd�-�B�\�����I��mI��캻�D���.W\\���Rs��R�y�bu������<#2��k�rK��>���d��K��"���{�w-<7�@v	�q���I�����5�{ՂK�c6�1o�n�Z�1�y��8�6��TF��L�FT���
��\k��<�db�kK��d�pun29�O�W�է�rZ�C�wi��o+��j����7P�s��$������]m��s�v�.ck{�,�.4t5$X,so�{��vd���w�'V �q��Wf�G�"�g͇y��o����-�!�+*�Y�� 촸.�8�'�>ь�U�ӝ6l)*����d*qF7\����nM����I���޼aVڧ}OC˻ZX��+���ݨb���ܭݪw[z�Em�V�0-ǡu �Rݧ���[�3��V��ds�t:1�����,��T��z@�H��ǃN�0J:7%뾙)'ˠU}/��#:>�[W%ފ3w�[���	]�AmuB��du[j�\�ف.�/��O��wNxGǒ�\�in:�}��ԭ�Y�d֮�$��	ir�Օv�6E��$��ٺ�w&�Zl7y�����߮�	�E�v
��{�����v�e#�.u�=�i�2�+�-N֮@Ac�:�,	o����~VSP�%����a������+[B�gf(��+{\Wʣx�v��T�zq ��Շ���9��W9"�X�T�H��9�Ӹ;��9:���4�܉0���g:�4(6vفQr]��P���t��-5��w7����Ӡń�Ȧ�q;�=;;�Ve�s�S\�R�JД#s,X���]�Y�5K+V�Ne��������2�)��h�5�R�|@���c�z`em���kk��$�Z9\6��AT�x�lYP#�������Q��I6%�D�dg$
�ї���}+k�������k)�A�V��6��c�r���Ǒ�V�o9�!�'�Qx:K�1�h�d�̋V�v�P�&`{E���]��֤f�w}�c�+\��a_aʑ�7K�}��kn��ck���7w�/^�M=J�����)�k�	�-��P@��A9}2�t�y[3+p^���p�7�$%m��t�w[�E�x�P�r	�J07g&�tԔ(���=��yX�.^��5���]�㖏���%�y�'�i��~[�m�/u��F��<:��~����.�U��m��\�%�[�ic]L�4NP3ZX-�:�P�Z��[ǌ��c8R�B�!/�V#�JN�T��ܭ��m
��yt���>4��6���K�fխ-�ڎ��X��D�_Iͻo^���X��ETD�Q+EX����Q�X���j (�EAE��(��U`��E�%�X*��E�UDPTTQAE����QDEZ�T�Q��PE`�e�QQF���F�+Eb
��T��,���T�F1F�J��+Z�
��X)Z��ȌT[j1DkH��D�
�cFT����kB�E�V�
����DB�YFU�iF���،A�[J�ڠ��V�
�1����ȤYR�Q�DQ�UAJԴiKb�Ɣ��m�%j���T*6�-�D*F5������mB������V���Դ������J+"++%D[F�,QcVѴU�����,J� �iQQV6�A� |P����	�Xs�V���׽�+]m��rMKr��PX����I�W��u�a�9+}XQD��t��r��d��n2w��J�o�d������~���k�އ�W�k����V�ٙ;�n��w48�!��2y��]�ߵ�/������WV�{|��i���M��Px��S�S�4���C���/��T�ւ 19�V�^�NAG��UX�\(�K�L�u;&�*1ڵ�ʾ�b��o{{}���7�� y�c�BOEB�*�r��c�R�h�Ҭit:�t1���.j'S��7��q�M��})o�UƘ��AjdF)}��CvB����ˇFuLD��
]���BS�հ*����˛
]b�)f��v�[�F�`7:��yr�s^,8g+Y`��zao�=:��J���a�;���pX6:y�65�,A���{G�2NC2EJ��П��n����B0ǡC��]��;ݸ���?C��^1����qm򛒴{�����ˈ&�P4��#t"�����پR.�q&�&� �V\y+�[Y�Y��`�ɑV�5���=���W�Z�,ϴANw��>F|��,���W���'����JL7Is������)��X�d��pt���w��[��f|HeA3-������ͥo\��q�qk��ӭ�f��k�!cW<ȶ�@�)����>�(��ѕ�q����U��9�bm��i�GWP�6I��{W�Xԗj8{�r�I{uAN���J��j�z��ۋ
7�5�c �$�Y]�k<}]���S�Y��Ä玈�{��Z<��G��L>�rǇ��͜�H5n�M��Ob�I�R�
�?7�0b�-���w[5-�'��d�Ri����F��u�t	�U���R�g
u�����M{�C�X�c�wS�+dյYzY��WGk1p�`��j�q�x/(�{F���SW|a������u�}�];�{�N销��x/$��˔��߱1oxC۾��N�c�W���`��F5ƙp:
:H��*烣���qǓ�7��˙�[wy$�U�tF.+�Wga�����G����h�s��4{��|�{���̴��.U��ܒ����#XwCI��Ln�ר#<TmTM��*\���F��\U��I/��e+̞�]��CL|z��c�l��F�+��V,f�\CB}�"R'�Z5��wKzuy��{[�i�.������׫�뗋ы���1H���Q�P���V314Td��V|-
ޥBI��[ԯzI�Z��U����U�)���\>"E�eW�]�CSb�D�o��]�E�^�A�x����@�!W	x�lf��v�zŰP9��W�3�x9J�:;���t4<f!+F)�����vk\���s1l�2�8â���Ec�LjB�Ð����=J.��M�F�mɏP��kF�k[���r��ڝ��'j���N���}�,ல�W�����zjˎ�ͳ�t-����U����[��+~3��4��?qt<��MC7�ģ�P'r["Q��Rx�-�9̘YGzv�'m��Mv؏0���D�
vdZX�x��B��j�x����(8�O����D�Oe�a�
�Lzzh(���r� �­��*cY^��
,&��h>]"*�=��j:ꇩ�Lsn�G �����g���Ό8��qu6�Y����AO���eu�����S��|�d� ��~U�w����a_M�М��s3*�^�Q���Υ�k�Z���z����cG	f�a�,<Y�@k�Cժ^�&]}�i�ԉ1;�*���P�V�[	Øӏ��OY`z���e��B�p��Y�������(;8jɷ�r�)�pޭ����Q�|�ʇ#~�K_��Nx�Xx;5������˭Lv������7Ux��rv�h�Փ���_J�}6���U%XZu�R덟��*6��]x^��p�v��ّQ!$���4�HK&ws��Uη�������+s:u��N�#�^5bx^R&ݮ��g+"��K�p�����F��;���=�e���bG0�l{�uNdtT����B���TQ[��W�p��p#�>�㙫��Q�v+Q��Z���ba������Ct3��T̠G�Cmnl@�;w!G�w.7�Ԗ-����s�ǅy�{V�%�g�i�=
49��P�
��s(�^����%��=��D�Rc�Фhc�DڮF�d(G��..���aI�l96"x�b��toF�8^�7��ctj�@/��J�����5�3�ʀ���(�Ӓ|�M��+"2�b���㞯=W���Qψ�xk��i���Lj�c�0�ܪn�9�ż/";;o4�g49U�o�j2�`ՔDPY>B��2�E�"B�������en�!��\��::�;�`\�Y��P����:�?M�s^b�|P�9�tȆ��Ҷu{��.�k"��'�5	��1�Q�z���*[*�\P/k����*���W��_�������f�	���{����t�v�P�l���P�Niłz.�
}iϴ�i�,us��Ĵ��n�w�ܘ��w�������:��>��}�{S��5xg��貶�:����Yn⑫m`0ݣ�c�6�<�|x�.�IG�k���TVN���fT�o	���U�GHM�ډ�hX�S@���m�iaO;m��3qh�kOo>�;���}�����7���8,X�dS��>�bVE�r��rΎ���d�u���k9�L���/�jxa�
_m#�5[LѴsvv.�K�gd! ϲ[w��R�h%g	<9���>9#����M��at�!���<}�
���eص���F���)㿧�.{��rF��K�><$��u;�#�~[��a�T�u�L��X�����ņO����u��qYuU��~�>U��"��5|/�o5���A:�t��CK�'��QN0�/U�.�[,ryWQ� �F{ND�[ή=>V�����i�J�J�z�5�tR�SV!��e3��Hi����E!C`ж�r�oG���m���(MK�����v���Q9޹Y�Z���p߾^~|�9�%c�jc�.܊�U�,"���#��u�ajy��	��fǽ-�3��/������t�\����>5�x?�^��~"�1��Uu�w��BW�6g`8�I��4�l*ta�� O�h�Fbh��]\	'Q���Թ���.�;��;���rZ��"h�[5�׮7r�w�ve�}���zvqZpK�h{$��wu�U��kc��+"�ڽ���[G�I!�ܜV���>r��QÂ��RZW��;H�i��vl�ڐ^�[�Ѻ���k��t��[�W.ۍ�շ�����g[�U�7��;p�FB��[������w��P�ܸ,<��3�6J�+�a.#+a�BOFEx�h߸���*:K���v�'�b��4Tc=���;.%ol���������g��dC�V����A
��l�zqQ�S.(���?<R�ka��i��j�x�{��;YV>���^a�iҞ�b�/�����x��S��(��~Nk�x��U�<��c�p����㩓�R�JG8�I`�lVNBy��اbc6�{nB"|{o�7�x�x�p��8lq�W��ϐ�`�6X^���E��g����ꄷ]�>�u8��Q��z|5*�1K��,�X�wy��t����dJ��+6z�iJ/�b����܌�J+�E�o�=��/�UjV���7*]�b5��}*Ϸ�rZu��Ha����*�7�h�T���B�[f���W����c�2��B����ŷ#4�{# ɠm�� ��}�|�jv����Ե�b���Td4bw��*�3Ƹ�E�t23ϜX�e����7�v<F�Gv=:{9-]�ё|ħ�7����Ni�e��q��Wۣ�ZR�-�!��f�y���e��U�j�g+C�qgU�A���3�ˊ��8��u�2��5�����U�����G��]�V�M��ě��Ǯ��Vn6���W6���W�X1��`�xtX����9`0���a2��,���U������ޡK/;�ܸzF�����˶k�B:oOFMM��3��:<Zt��$A��~����J�S�����u�~���[q��E{T�Ue���|O����+�WL��5�]2���^v(fN���hq
5ZSjV�N�su�b��zT+�>��V��{��9�v�)[ꛓ�}�OI��B��p��s�t;�(�|N���P�1��>��=���Sy�ð-����p�i��|���/��&n2��IĦ�=�{�z!����맚d;p���i�U�/j�0�j��޶�Z��q;W����>�tUk��;V���ì&�;	yM�`8���km=���t-ǎ�{���T�)����}L�U'Y�	��~�N�d�ᝲ�m�-��>��_�Kx��֎�'-�'����-��ʼ���
��F�����Ň�������E*:"S["���F�����m����)��ڪ葯	���f�&��G
��*�U�V,�M�Ԟ��w���&��Ë̲��c�g�o�J�״����#Q�j�]3���΀np�6*��;=��F���:wCq��oOK���"�(�[�+)���ܝ۾�����Uڦs�G�T�Mo�u��;��y*K1����YƮ2�%�?t��puKq����gP-mf�$qy��~]K\7;D��;��P��2y���IÐ�����c�NwV�/��%is�o VhzWve[]��B�WTڼ3C�GH�94����u�ƫ�VV�[�qTy��wi�P���KR����l=�7A>�W��.�����I�Rį.�&g�j�v����%��j^e��5��7,z�F�4d=�]�!�Lf�ɜɧ�v9�mo.T�^M%`��:\k˯�z�p�pv����8��>C�d�/��*zk�'��Wu�6�N���Z��7
�e�f���ܯwY]rc��.���1)h<E9�Wg\���LOm+/�����-v�װ�U�Wv�5ʜH�K6�L�V*�N��}5����6Wh��P�� h_\�c8j�7�b�h���e�%A��W$م�m��ed�n�ϗ���gE���O�J�y�����r\qK�x�Ì�9���:���0����\�i����E嫚�r�gp����U�����3��g]J�J}�op;ǐY1�:���~�����|�Q���M�C��o*��Cw\����m�V�Ue�A~k��Gu,��L8�7{�J/Օ��0a�yI�ЉN�E:	ˡ�Ў��9pnk�3���/�s��~OⲣO��W����N�P�72��qcT�h�"6o��	�@���g�Rr9=;�Q�oٌٕ�R�\֡Md�]u=�fZVs�ր��q��_K���vg���e䫬�;���zw���B���H�Y��)�Y��xfi�.��U^���Z�Ǽ2n'X�J�#(u��Ԙf�f��3��q�����A����8�C�����ז��O}r���&X�y�����k��(؋�2��j��.-��C�ni�T�&�,�'�J��R׶���~B�`z�R��6��#֫ls�p���Sl4��`r�n����Ɖ�����U�*�!���4�k"��� ���L�N��V��;n$`����+.��teT�<w�u]�Y��܂ˮȥ-�l㼅Z��P<ժi���,GqY)��{�ۍ1�L��������\t��pT�y�ͯ���/�����W���DO^]`�������*㱝a�U�*��)���WܭPu�YX�Ks.q���^4��t��ޟs�j��5b�i�:"���e=R"��hX3�]��FI�_l��sW�jwq�[����_�&�s�.�WL�ado\�����Uإ�׽/y���ƴ�BԪur;kj�1!�,F��=��>��W�e��w:ݒ��naބ>�7v��ˆ�Sc_���S^�����'�����s�Aɯp������`���b���V�M�1�<Ӳ��_R��y��#�*�0�nח*�հ�s� �T=�[���ȥ�yG|�7����X6�T�c��'B�[�Uփ6M�3�,M�=�7��yyWe��I݉�c���K)�¼s����nW]"ҧtF�Ηak����ZzV\���Aoh������֙���.G��a�b�.u�ɝ�ٳ��eX���ov�f�<��\X���nP��̧GK�'P�����#�W�r��t���\FTv�	��ʷ�[P��7e�S�ͣT�mɣ.�:�ǑѽV�`��ḃ�����<����r�s���p�������-ә��O��slƢ���`�Z֍��Ì���6���ocrVX��G#���f
W���V��5�Ur�F��Ig���s)5�%�_G�T*��:/T%طl���0�N�Q�����u�D��^�(ܠ���}�vj�1��f�bɛn����i�VE��M;��ig;�x3e���c�2�Z, x�JSPY�VWov]f.�FVWZͳڮ�!�Q���9$��Jo&�D�g^�O�VR��#u��Ad#9ڭ����Y���PC&���l��.k:��k���������,[����O6����&�"p^�\3U�;��T��A-a;�S8MC��F�F"�a:���4�ݨ�gH��c"�F��Eu���M=��h 7��v�*�V���W�~�
�Ma���[4e����t�FQ�+$��a��	>N�U2Ɯ�Pn�xFfj�{QX*kC�|
�E���2�w4���$����a콴��.�]���B�Cݶ0;W݉u�X�U��ä�w��V�ڴb�0��7�{:�ɵj�%dM2�e��IX��!\H�[ǧ� ���'�u�g���=�B��O�g���Ɏo��ɺ�\��תgKR��Y�v��.Wwv�]-�]��!e�2��h}�=��{b��U|���(��&9Q$w�s��Vk���[�b�͋g�FZZ�����s�L��.�� �G��\�Kư�un�&��8�j2�0ɉ�[�t\O�t�M�x�,�Y�;Ww,�W�b���$z]Ô�'�4����U�Q}g@� Tt_v��sv۸/()M>�Up�gZ��x���غ�!n͎�+�ZA�gR���	2�B��L[y4�*V\�(�W��`�S���Ŏ�X�p��&�A��& ԙaX�ܞ�\�}�*�LS�Q�z o.�]g; ,p'\�Am�mi�*|U���=m�B7z_n���'�\̂�q��^8og$/������[Z�Yï郩gxfSY��P�������]��Z,�i����L�Ұ��'N̻;�yG�]�!y):g�����5J�w4%�C�*K)�v�_(��Ԅ�v��C��짔a�g/]�C�����;��)V������Z����l�T��z�S<h��+@���&�Ŵ��n�����_a���8P�N�����83�s.�+Q({e��뷡����]�%�V����(V2�z@�փ0�:ø>+z����m�RƦ�/�¸��	F����PW�EGi:ī�X\-�Y��6��;�q�͡y���}ws�ɥ�cRءYZȣj�PFIDX�k+-��E
(,m�++m�*ZֲE%`,���U��V,Z«P����Y%J��kKH�[@FAH�IRV%E�h���i�YX(��Imb ��+,PJ±Jb�E��Ɩ�m���+P
�m!Z֡UP��D�2���keJ�-m�B�����E�mTmR�����%mF�X����KK
��5�kjQ��*V+b6��6���U�P��Y-���J�h�Z�ED�B�J�["�eAb1V6�T+ ��J��U���J�¥Q+(��ZPF��)V�J�����c�����;湚I]E9^����;��f�ٹ�1J��d�P�Lѹef����ڈ7�[�ഉ�P�z�E�^�\.K��v�5š��+�n����O�v_���k���1�E2h���_G�]��2w�TW-{�3��v��>Y��y�ڞ���k�ޱ���.۸ي��x����T�56���=k(4�^ՙr�]|\e���u䵔�&�6x޴sk��Y@d�"����կl􎶮��c
iȩ..�\���M��a��@�i3^[��u�~3S�u�V�$[J�:S��H����_n���!\^{���}�޴}o�匢��^�73�2���r�33St��ƾ�k�6���8����ϖ��dwB:cz7�Y��nn®�ŝc[�|���{��R��_Sjz�䓱�-��l���c��®'_����L�N�J�r��� U�C�sqˆ>����ɪqۋ+�4����zdSf�����UcN�ud�ޒ����p�2��7e���Ȗ�#���X�h���� 75���w%BiHөb�j��*\����;f;�U�6�X������&w������{n�z􀷦�ֶ@j[�D5rp���S�/�
Nn��6;�giݭ�t��N�r�^���b��_pF*�M��Rh=p��Չ�����1�q�z2�:�dlA��R�R��JaI;mvXvߕC��<���X���z�oS�1,�)*9������݉r��4�&��^��Й�V&��\j�W9�n��Ku���2D�q`gvh�{��9�p�˱
c�y���=r����nڻ�qE֚��bj�-w e'46��Ib��S�g�m���	f!V��^}!��=Rv郝t�<��S�n|4�q��bV� �������_����n���ʇB������^�s�=�{�i��9OP��2�%����o6����y`��3�^�#hj���@^�XR��y�P�]�����ɐ��}���٪�h��]P�>+Ѭ{��É�Ac3�{'���:ؼ�[�uc��J�)y�]��Ӗ�{j��s>Α�0���L�@��z�݉5�)�<DYxp0�q���m�ƫM�Jd��F�k��k6;�y�F8U��f�z�;��l}Zl���7;�G
考rc��(%6�M}�n�ݫ�e�����B
]��kU��5%�lU����^�4ona�e���U˕yi��-=�+O.�Qg�Q']۪�:
и&v��%O�wD�5^O�G�{>o���=�}�U���Ru�����[�	�V�%uU����->	��)^I��sٚz+�|;�|��fW9q"�"�m\�5b���������X��z��F)�Wo���m4;o*����Ƿ��%Δ���xm@,������Z����x&�=FL�6w#�顽��@T,��#({MG
�;Pg�:
̵�"�9|��m-����ƾ�V9�p�A�[�Q.mJ�i&Y�ʍ,���"��k/��"S�QN�rØr��ۯ|�p
~�N��jQYQ�5ʬ3k���e	�t.�i���V'L��ʖ����0P<����M]�n�9��G�!X���F���r#9u�|3�&͗r��dc�ݺ���;�ғŁ��wG�N�i��w�z@#YQe��.�(xyv-*G��iaZ�F�OGnY�i��l	�y��X�Yb� ��*�1D�6�� ����-X�����S�1���=�t>�G%��3�5q�F`f6��dNt�h^�J���'
|�I��Ş��EysǳFy�:)�b؋T���{3�1��)�+��C��Ek�T��>����^��oz��5��qY����ӊ��|qۂc���*�g��wBe	&mU����=Ϸ����m}<�l������4���x2���F��(Z
}�y�
��6�ާ8�y��sj�(�[f�v/��nPIF���\��OK�iFi�h�(�n�O��&�0����wc���i�c:�*���H���ءI��}Xh�����o	fd^������}��ͻ�AJ��<�L�]X���œ�ll�q����u��j�W���wJ{��n3�T�n�ǁ�ʪj�rR�/g��������so���������Խ��;@V���If�'R�-W�k���3��6Z8���nme�k��ChX����e�l�S����֍��YV��c�He3N��9�Q�'W+{��u-x��a�ۊ(���+��5�u`$���^b_ Mz{yK~Es�kib��[W�au:�i*ڰ�Ro�5�*�û�fՑ7�t���T�u��ez[�z9�Q04I1j�m�����AH��TNtԽ�r+dX��sA��W���偹�5LHG7;�:$��3�{˘�C���c��u�O�s���ed�%A����}R��u�8�4��7�8�{
c��3�!�]ؚ��N�B�/g)��d�Q�t��FF�L`�ą�&�u��U�A��cn���������Ū$��z��>����e{i�:���|�k�O4�S�cQ��ܽi�X�=�*���1�G:�NSvJ�f��er��g*�r��9܍�%^�&#�+(�I�U���sh��9Hc\,��׃g���5�PJ�^��)�W��L�+z"ޓ4��f�3R�*�ċif:��d�мy�7��:��X��dn�7a5�j�Jq7������f��ꋶ#\�E�S��=�{��Ҫy��q'�;��_�{�X*T�y~c�d;�`N�Sc<�:�����h&ڶu��k�dMDl�rq�2�*�5�:KQ��HQ;�t\ʖ�!�4"o�`���a~5ܽ��6�ѕl�Z���݄
/��6����:ol�d��H�t���;��w.�H=o0"��\sp���ڂ�e�jnG
�رlF�us;��#ᜧ�KW�?n|����uͣM��rV�)�뢦�ܷD7�rD�[]�Gr�z�<��=q��WX�x�v �A�a`��g��vE�Uo�^'I�{�:R�BB��w=��ksڢ��ɩ����v)h4��7�^Ɲ^���'6ĝ2a�ʩ����γ�m����"���!�n!W�u�-��.�R��GUMe%�f�cԫ*Z��
��2�^��c�y
�Vn�A;T�{��]F�7�8�j�.�b\���h�Ͻ����y�J�h�,АMî�x1�u�c"/�ϳ���s�Ż�6�C[�f#�;�jJ��=��iۭ�~'���y\��-��:ں����{��*�U�ђ�q��.�sN1v����;����̫O=����޸;K�=����{Pz��,d��Z�R3����u�/�u�L���anc�i���[FWq��k�^�X:�Wm�i5�۴y�4�̽��S��뎷+V5C�niT19b>5�!�gLJ i>��ט��Ұx���͞��8܇y!�!���hCtT�m�̕W���B�q��De�{��%\T���RK6�^��G8̳���Z�W�ykXN�2�G��)�˥l)]�:T�n�ÓͿ77�Xi�
��]�76Y��`y ��l/��fN�\�K�)y����6�t�<ƛG�vN���cM��~�"#�X��U��T�I�����!Fͦ�z7�Ʈ��v�la��6�b^9AP��0_5C�򴧎��f;(�[q0x���n4�N�c��^SШG%BV�%'�u�ٞ�d��cs饾���Ӿ�=U������ԩr������f��U��k�[3�{K�e����)k4�O��mL	搯C����X�w���+z����f��}�!5C�l������{��&���s���2���k��5���^̖Pӿ�Ǭ��#�N�2e.�j+���rS�.]qmmȌ�t*4�>f��JIM������u��3u�睜(K|�q��{R�F9��Z-����З\�wZk+]�͖;;E�Y��}�.���F�V���Hp\���5۽4PŖoX�[�Mgz5^؆�T&؍}��s���Y��� j0I����q9	��1�O�n�a�ڟcu���NЗ)�������:6\ǜ�N0ɪ��6�ǫ��:���A���E�9-� ��P���m1��n���ssC��%K��;��>+=r����S�vY�3����}���a��1�h�m�	���L�Q��q1J�N5��YȜ��;�^O^8�va����U��.
ke��B�o&����=^�zhy�F���-�Zt�T�7y���78�4�{�e��o:+k�؊��]��پ}��[+���gVV��q�;�ǎlR��to��#����(���7}4#Zh}ճ�XT�8�T�Dٜ�oKV؊Yy�3�3=��z�Y�N��@��OK�-(�Mnȧy]���*�����e�!`��uo�� �Q�;ihP�]5t�*)g��ۺkFjyҥ�`��U�Ԓ֌#�*�S�wH�^qU��i�n�Қ��C�;8t�l�
��<��*��*��	g����^�	C���w+j� �dt6G:M��=�v�pt�%��[�{�6޳H�N�m�*���*٤��1��c69r*��a�Q�9=ڝ����ܯ���ќ�3�P�#x�z-]�r���
V7���눴ꆮU{��i'�}oc�@��p�I��S5e���+�&�PB�q�3Iؚ�#V�{��V�Vk�{�:�+���ꯓ�7�z�Q�!��	�� �������ˬ�Ω�ePUj��L5��N: �R(��':jV�$V͋3\�����xY��ۘ��\x�w�Tۭ�r�C�#���T���D��R�v�ue�<w��6�U�ή�"xO���Nr�}YO �;����X~9�+�\�쫿j��+�OR:�Eӝ�elwr1!sɠ�d�U�A���$\�GOS�c=駫^]q��zU�7�z��e>q����P�q���}�Mz�#ލ:x��k(g�8΃Vjt�:[%˱��mVЎ�4�<�Z�*Ɏ��w���9Jv�]��jm��[ӄt)��N�l�x�!��Z7�+z,�Qt�a�zU��L�d�
�ܖ�JN�C�P��ۄ�b�ל��\[Aq߱oyuDn�`�,81���L�Um�}c��*�M�W����7�{���s��^�|)�t���;��>�޾�d�x��|�;��������Ɲ��3R�(Z�I�v��Y�X�{�>ԍ���N[���������L`���/={������7+�W+�{�_V.�M}��U��}�^ti�^�P��ǜ;��J�K���eZY}ʺ���+�����=�a����w�5ї&81	uxB�t	���Nȶ���T/�;}μ��Q9���TN�l��@����YBN<(�h�ڃ��:��u��W����:`�\��\�5Ҙ�`5��Ż�p��}�ڲ�5YZ�� �sW���:*]��;s:���\��Cw�Xo�E� ��r+0�B3��G2�a1bvr'��{�C��E�Q�j�t�\u�:F9�kq��"f�.RS�=Ym��%�,�hD�&�Y췙k��k�ք�)+�x�-R�iZ���Un��kz�^и`t��@�)�`�/�@������L
�R�^צp9��Qr۽���+�7%����Y)�hQ\�ݫcn�o�5QWjة��lf�Nl�[3w�ӏ/���6}`uw9R�ǫmj�h.U �۠RH�N�Ճ38\��{��A��2�n�^R�/q�r�y��>ucRSIb�5j��2p
%Ԁ��������.�ps�y��&�����A˘m�eѬn%�%�&s�����T�u�%q�T�(b�}�٠:n\q�w�� �u����F����i�]�t�d�ӛ�'5��;���6�-&+WV����vΕ��}��XRe�Ő�`�h�:2��3)Z�z��L�`u�8&��(�\�9ǋWz4��H攽 ���>z+M�9De9�[b^R�i���O3�֨yH��EIV��U8�:�R͊�Lu\�*|r���;]�JWU�rF(�}+Z��b�}Kh�y����3��k���^���km�D�G�&y��P�	I֤埌Ǳ�ꀝv����t�׳*�:�oU�C�h���U%f��\���zS�6����*�N!��t6��$��V�=�ǥ�ҥ�̼O�Y��-!�ݧJS����[3'ěv,�X�SJ?$z�DP�������)��rk�!�
ᢰ��P���rU��mT�h�˻R�O�)��0����	�WW]N-\�؏�7�WM<��Ͱ]:��+�NV��z�J]��w�b�4��mL=S�� c���{3�<�����ח���<w�/<B�:S�� `Sln��Л�l�T��]��T��΋u�++Lr7[Y{����N%�0ظ����.�[�qJac�;����$��PU�Z�-��j���ݓ���&k���Į�JU�wU�©��3l"Bb��V�����LI�A�+*(~ǆ��umDk�r����d��t�3' �F^K���̠	ըm�`�(g "Vj����t���1�(���Ǳ���k�K-�V�Ɛ�41�����̫{�V�RٳiFa�B��I�7qnH���i}�vĘ8�g+8�U��6Kv�/�\U�볘��ݕ� 	�D�.�����!��fQ��C�n�4f]'�ݴm؉`q��pP�Q;�7)�U���ror��nT�`�<�v����:[ո֊�r��*����v��V6\WZ��C��>��$�I�("�����e"Q���Y�_�k�>��VN��kk3m+��N�IȌ�gB���r���\�1�J��(���t"�״���ny���dPj�֬)YYm��YZуj�����-��P��Am�"F�TX��PX���,��-��d-��-k"���������Ƞ")(±H�(T-�1�X#Jŉjª*��iJ��`��TDF"2ң �R�DXʕ��T�@YTB��`�U`�YTamR�QUb�Q�j(��(�)
�
�QP+"�E�����V[j�@ik-�
�*TT�ƫjT�D�J��ŕ��b"�
°kejB�Aee-�[AFAm�UX���[UUE
2�ł%h��*1�Q��TX-A��+�����E�eB���Qb�H�)R�T(�������V,��Y*��b��eaF[ZZ���Ъ�mѶҖ0U��%�U��[YjEQm�ֱT���Y+cV
��H	�x�ʏ�mMg4l�+`�+�0�{����i���[l�ڇ])]K�}H'%�xAM�9yǲI�va�s���l�n�CLu������}����2aU����w�r��-��8�js���˕�t�t�{�2ݙ��lD�@%�ys�y��)��TT��F(�=���B�w��L�ۉιu�JN.�y^�C�yt���3;�O�-��y�S<���1�(�������w�*��9Oz��w�85����zz�ub7ќ����ݩ��oj�P�\v�{ȥ���|{rSs�';[¹��b(��Y������uP�@�F;��C^��bfۭ�T�v���a��<�zR�u���=4�t<��]��O'�'����]9�u�,K�(^l�=�6ym��T���۹䷦�ލ�Z����Jv��,��l�ʪ"3B���4$��C�
mi�J%���{���W�6���v���@��I��H;AT����E��r�#Z�:D��G�0�Gx�L��􅯐�Ǆ]kz(X���A*{�Q�E{��V���P�~�5��sK�i��� ��M�v:F7Q�@lk�+x]�oq|�7r�:{�([As=����kolvk�ԫ]�̜Wܞ����7Q;����}7�
���؊wӥ��{Ѯ����b9U|-X����= �V�V�.��ū��8
�y�c�9�-��Q���3�7l����Zi���bdc��Ź}I��=؝�`S�4�^ָ��m`��#����U����FR�J#�����ջ/����7��oO��A���c�
��P5]���sK�����v���9g��x�5}�3�r���u�(1݉�T(B监�S1Yh���Y2��+��_������!.��&^A�y��SKc�:�'*{�YY}�?�>�Q�.�`�J�g*^��YoP�r�8��O}�(���C�j�q���אu�zj�X�jpʚ�i�r��԰wPξs	���q�j�]�ž���]ƽGՂM'�����޹`U�۔�y��W�<����5�vN�������s7��E��`��:�j��.��<�w}0-��4��}�<����IY�W<����'���M�M�R�27q�6#����u(��ЩV�w.1��|��,�^�~ۮ�i��Ӆ�r�V!ĳ3Evi��$��=�ьb��D������@3{}�x�y��:�z��V-��t�.��䇎�w����Kx�'�;��r_f:�����T+͂��!W�6{�l���J���me������P���vNO=�X;�����5�4�$[J�Su�j�.�nwO+Ӫ%r&m��v�-�
���k7/�Uz9�B�sZ��p�nn?{k&��.����tӰ�ۛ��mk��F���V˪�JBO��$�Ù}��>���9�d��v��ndS�^�z���+��E�7p�*����{Q����&��'b��ꪷʯu;�����N��:�\	���]��by��������oD�'u]"�U���՘��]�Խ������k*���{j�9����<��W�1�ܭ]�}�=<�׼C�p� �?&�-,\�0���T#{p<x�E¯��/ml��X0�Oc�r�d���b�Uh4���]z>�3[G��]��֚�oe`p��!�H�ͣ�c�0�~�̛��T��d��=��:�*t�:�6��u܎�!�6�p�vC��[.���eiT����8vEx2COm��YD�N��ǳ����6�b� �����%ܱ+Iz��]���WZ�m�3I��o�<+���˝����^I[5��@����C�
Ȩ+��T�k ?Usӽ��饎�$K�G7�v%��t7^Nq�fn]�5Td=sϐ�ws�'�����G4���J)v(�=�M�b�� �s頝d��Q��)^ou���u��9�Em�]�Ց�o#	�]�O�oY�lf��帽�D���&�gUw|PǛ��,�:����]Qo����m�2�ڵW���4���qz<�����3�^f3hwBr��s�]�Z���?k�9{�	ҷ��^����^>�x���5Qd��ֱ�h-�<Y7㗕R�L�h^N���t��hOZS�Moz����l�\���'fS]N�T]qűMF
i��W�5�b�9_n��x���ѵ��[�^��]	:
���6h7`�ID�[���Z=��Տ�+���#!ick/�VmG�پg��x�9�ua��v��*T�򣵞�4��pl{kc���N�O�˞�ۗIQ���go-4H�D�"�͹�۱�Ⱥ�fN�s����t��%U��M����rQ�Mt�~][����j�i+="۪�ʯ�S��y�E�����{���%9���j1�;�^e�w(�ʹL��Qڍ�kP��SGlbX�Ef�%�r�-�t���W��c�_2�"���0��u��2���*)�����jC�^_�rXK�o8<~Sv�M|{��Ĳx]w��m��P@��]!ίT��[^��u��,=�V�C����R)e7C�St�n�8�x!�V�"��k�Y�"S�%�˝k��{=����KG7Wy�q
x1g��LՖ&�e�f�)9��'�Їw.�N=��eD���������a:���r0|��g[]UԠ� �{7I�w�WN���YD?%��dז��ՇY�F�c��8���y~̤Jo���dDu㼼�(]ѧ�Ht�u*�y��m��ᗕ�f/:�l"̚4r�H�+e8�yFٚ���p����L,�s�����o�>�@e>���-;��zpE�����܌��/f��?dë^�Z��q�q��o1�S����Ԥ�]�/����k���Vѳ��۫�N��}mÏ�����*u�4�ƒۥ}�m\kΗ5�)��,�ko�J��|����:��,M����5-ڊ�ڲ�*�ҩ��ȳ�[<�ä��O7m%�r�cj�]s�R�y\��.r7[�U��`Ȱw��iE6���i�m��t��ރf�[�y�f{�kcgpy`=4 �x����z:�,)�V��;���J���7����l��gV��9J�Z&R��-�܀&��7��b[v���
���i;��>���<S,W -���Q[}K�`��{ݶ��e�b�Y��)��w��gg+����}�f���K:V��R�s4������ju���\����op;�dJmL�꽘��3%���+���Vg]�Q�h��[8|[����]{�Y)���ue캴1��ɷ@��G_D��މ������>D1v�Dt�Wr^��j�hS�>tA����yak�L���9�qA�<�Xr�P{]�����O��߸w{[k2.���\F�G���ݽ�1�[��� �:�����[qĶ�i��+ �rơր����T@fn�6���*gtM-��FU�5O̩��
�tƱ�p,����>�R���1Y�AY��{ܹ�m̴�N�P���d��5;)#A�n#ʤ��-뻦�m���˺������c;����{V�M�5�8�2�	U�m�CUw[N�y��[��Vd�im�,-�:_'q�sɧ��'�:���Z)ٰ�֊����-OU�%�C���ߋ�W�uE��C�}�Lx�{vdaSq�S�HGTV��0ҩ���f�l�Ò�^t�=�6R�r�e�rEEd�n�*j�lp����9Y������w�B��hH'Z��4�DY֨�$�0{��&�l�Lns��u�R��Y���_�*�B�=.3h�Y\�1�ied=\�R䑧=��6�nX�=�̺�|+y�w[�f/j�ǱHm@�ӬJ�r�*�wGr�z�>��n٥=t��{d<�6�@ڞ�>��^i�K�2�ugy,�_m�us�D���GDfG|�;��'c���8�qp�ݥ�6��Hd��lj�����.�gJt悪�ƘR�����"�doG0c���vN�خ��e!�Y���7��ΰC�)��r�ov������ ��s3G`[^�S�I�O��3[�{y�3;�Wn���Nc5ފ���M��l���j]M�j��\y���~����]�u5{�%s164���X��]����0��W�WW��
���:q�r��/F��O����]�y4�v:��g)�MY�i�k���Qp�D�Mz^�"uh��;�*sɷX�,V�o9�B���Ձ6��.�z����'��dU�V�r�Ĵ�ڗ:�un�
�}k�a��ވC=��s�3E�S��OHֱ��,j�uV��J��]޼zgi9�c:�LW�������⮦3��|_#j`ڍB�m�8�+.���@� F�p�`�fͪג�2�6����5�m��y�z����-���gm WT.�an�;��
�v�K��a�ȯ)K7^K̓��w\Fn�w^��+׍@��Ԥ����f$*;�\AW�V����Ո��g�/�&��PƁuJ�v�l�k���R�KR��o�U����}���Sh�i�,��gV�ō�3��������rwJc%DY�y\�$�A!z0n��Ntv�5���p��z��2��}�N4x�F��·��]�O�ұ�� ��Dycԏ�_'�k�e�1�F��$ZJ�S�J}]�^�}����ٷa��0���L�C�\ڙ|ƜɕL�>=�EwD��wZS��mw'/���ڂ�g�{�t�ܕ�vpT��,C�f�P�RQ"��u>V�WPzv���%�j�vzL�ｪ	�����L>�f����n��*��&�X�7�.�Y�ۖ��F��V�yˆ*7x:�y:|��6��O�"g^_fws9��lR�k��p��P$
I�[,��j���*����0���v*|�����_`Mon���t	\Շ�[���W�_W��؛U�w��^i1r��\�L?T�+�t���JQA;bJ;׳������[�O����A��n��i���]�#�����'8���n�,j�8XJ��M<A�@����%o;��N��
������ã��,��_V���t*6�O����Q���b�v	��Y-�9���B����]H�Ӳ��e�+��Շ�����|r�]�-�7���V�^��LL-�RJ�];S//���Yz�����*���s@μ��Yx��r���@�>���̅�1�S0����v�B9�k�\�������ϼX��w[�rM�;�yu"VdF��1��+ݯ&�[Xf���w���ק��9�g�����w��k���>
k��'�+����ypy����.I	؏��'m�~#"��o��eq_<��jgg"gy�M+y�i:O������[)k➌�roV���19{;�.�w�b����;�q=���I�-�N¾�hF��m��\�#N)�m��IBk�;ӝ�(���zs}������g����Y=.��|�/vg-K
EûWX��r�sֽ�Ϛ9�<y^KLñ`=�ƕH�����Uvv+�w�+�E�䴹о��I�;�1��n��
e��f�G�mECq���qx.rrH3��3 ��`�CN��qo�0%^M(d(�(�B0�5�F%v��c�.��3��.�N$W.B
S�4�K}&���buj`殉{g@Z���ױ�d^v	�艥i-�����jU
��+���A�쇃R�&Qo$����bnNeWm#X�a��,�Rack�v�R�"w���Iލ:�$1�W��vG�^w��7���Pz���nO�:�t�2��@C%��Ѳ��aܺjֳ	�	B����k�� �[�{�%*l���Ej��j��f�}�����O2����ҹ`��yo	�%��qu�p�N��rO/ *58�$hۺ��*�a���c���P�2.e�-��;��ۤ���sLg�u�v9/��gKnc*��d%&��c+_<:�����P��rF�|E�7l�Θ���,j?
X��):U�g�'b{hR�8�Mm� �Ki���܎���hg�Z�Nm���ӧ��p�\#�l�tu�ŠH��%�Ʋ�=C�-]���쁏����i�;��� J��-�X��`�*��ȱY�x��3��V�-�ũ`�VgmYܝ��V7.�����x
˾�Cx�LEF˔�=YN�ޗ�
�Ȯ�M��.��K�����mM��^f>����; y���`��{}G�]�)��8��Ҏ��ga�]�T�}ȭ��7>͠3�+���QE��b�p���l��*�5ժє�79JU��A����mA��᪑k^���TF�v���қ��=���Z�?(e�ͩ���\��q�!O�)|��0�\H�7���E��cp��ZV�Ƭ�L-;E��S�+���Lv/D�\�[�EJ�
++��U${sK���?$��Td�vFV5pE.*s�4��#����+��'i�q����}S�|���h�e�ۓ2 IE��c�R�$v�,ͷgw��'�.�K�8�,J�r5�
���'�V�f��M2���u����Sz��Z�U�ü}y8
ZP}*�'�]n��­S�sZ������� ݺ�)C�ֶ��$f�;���ZSRu'�\�VlWyۿA�.UX��zS�.�@E�7��YLֻ&n�>"ե�IwJ��\�����ͻN�1��5EPc�'�ۨ��P�㙆�A󩣷p��ge�t�=��o.�:M��t��=��)�f��J�r}���oV"3l���ƠZ�q���Ka=��c�����j����2ܱ���"��U^uup�@0h�����<���|;b\ܼj���G�{o���:Tj5L�h�)�壜��ja.�b���e��k%��u}�k5�<�������N#����f��U�:tETm��ԅ���Q�+l�,eeB���(�UR�Q`,UX
�#
������Jъ��"ƖQX�FE���,UU��X��"��EUX�Tm,H����),Qb��ej	l���j�����`�*��R�(1��(����+(#*J�ѩ[h0B���őV,Z�*�+[,c
ʊ"�,P���X�j�U@Am���#H�[J�d�+�Q�jkTkX�P��U#l��[k(�m�F���Z%e�J�B��*KZ���`0b"�PF,���k+
�J���,���H�E��B*�m����kA�hdUUEed�,c��(�FAA��U��ARШ�+*�`��,b�U�b�X ���cDej)+X�D��j�dX�9�����f�+��n�e<Y�3'	.ac�^~�%���'��f��R���i]�X�������3S��usC��[ӪH�=]�J�ȬF_�ķT-U{�ߩ�O�k�μ�)�5�b���U�>���W�es��s/����v���rL߄�H~R��'+���Y=���7�~�^��v�����ͩ؀9�{�l��5,vwBku�R��wt�iFs��W�_K�uNK�w"��6�*�����ok�N�0�{�O��or�ޅO��c��s���s�>��4����u���}ٰ�^pz��e����;]��Z����G=k�&���w�}�!=毪u#�/T\�
��Pʤ؞�bB�M��ӛ� �Tc+$f�"j���u*?���~̩���6�SC�Ϲ<�\�k�o�y��q^��׸Es݂d�e��`�T!����Ju{K"�E�&C����� >Y���fv��(f�9c7�ϼ523�qoV�2��JX����RtM\�A�Ss؊�������uôo7e���k��>�R��d��e���;1������'���z����a��QҐb�kH!ȵ�}�q-�v��ƀ�윖vX��ՙ��^��!n��P�(�:b�ƚ����*u��T��1�#��!�y���tmw�����W�23j���s�:���rj�e�b�Qe�ɼ���v��mݹX���j7,_M*�^3A
�q��nLrh�X��z����9��[J�ԹXF��<�O/�t%��O�	Bk;��c�1̈́�l�ҵ˪�wGr�z��g7L�9[�¦�v=�Oit�tq�nB&R�ʠ�c�N^�a�T���;���b��ݷX$$ᎎQ���W�n�WH:���u��W+��=nV�!�M�����ȧs��K��P���j�]�d�o�-̍ݓ3�P��K!���R#��#s��#\k��(W)E^�]��5��4�!R�wP���j��i;��e��]1�Q��hT4w�t\�����+�$ɞM�c(���s�@�Ou	��w�݆#��N��g�di*pc�h_J=����k�f*.�7NSHe���PU>�_S�2�٬�ٍ8�k2+k�Z�c�s�:��:2p1�|f���Ylۜ�9{���ƾ�Ā���B���[h	�P�6�ֹt"�׽Y��Ox�0�ǃ��liW]�%4s4�ukAd�Xl�[,�Ļ��Y�Êj���&�^e%�t��Of�2��g٧�>ipǉ�m1#���y;(wO;&�(���ٵ�FUS�G!�[��i���R.���ΡDv:�T!�\Rv&�Ud���ڙO�Č�3��=��
�s���*��:l���0�{�XWR��6�����u��My��c7|u��@�7�"pB����l�n��+B�i0�e�{�*}IKͰ���>&�U��{���|�?�nAnܢש��j�Oc=|����R�iZ-fpT�����;Ū�����AU��4#x]wD��T:�+)��RT��GE �v"b�R�tUv�'d������BTS���K�����]0�]Su��>JW�%��^y�C�TH�rR>�f��S�m�Z��Mܦ,�wS��B�Ŗ�i;��o^u�m��.��P3ih���UsZ�:i�<�R��
�b=B
NM&)���f7���V�U��H�𭌵Ҝ{\��6����m�3/�f�V�G/"�2Rd�G�˹J�Z�f�{�'|���Oa����N�noK�+�����7��5..�c�ڮ��~v��w|�!ZYqyK*L��ؽ�C�}"�l�$��,��=:�S���뮥�hJ}O�hy��p����#:�7&�k	��x��!W*��9�_�=Ά�|�.�{�����oq��gEz��c;��4j
���P��u��i:���}׌:B�*��;����w]���J��y��,�tU����Ҫ�ƧB��38E݌�}1���f�^f�1��N�����b+��8���W%G9x*��v��¦���-JF�;��^Jٳ8��`FN�c�A�qi�3$�KQY	���9��V��`a��AMt��Ob�N����4���{��B��r*�6
�lN���wBr�X��A^����J����
x7H�;��<{������*�z�ڳ�3�s��_:"M���}��w@��b�Σ�v�e�y��;e�O��#����r^�=��TWk2�j�kC
]�[�Lc.�8:{d-��5k��+2�*0Y(Д��ٹ�WB��w|�^�����q�M�Qɧ�5^��K�)�K�b`��N4��60��xCg���s͘���؍�P���'�{�AoF�z���hH;�}]�M���Tc;�W�{2UM�q�%�$Ͷ��4��H�_����l�C����Go�֛97Ǹ��Q;�N�T��F�_����ư9{�V+9P|))t+�L�m�h�u^����H4�qݡ��su�2�BW��'/�͛���:�%
�g��Y�|�^�v)�>T5�g^+��y�����BYݽ׌b�2�W�(�\�}��ڷލ�;�f��J�yU��<��Xff����@T�e�ƍ�����ڜ�eL��W(����Q]8�̶��NaI~��Q�`��Yp��h���	�R�ܹ�'�lxWe'J9�|�OuQMs�މ��1f��P��T�h<D��;k��o7��f�,{�/�\�bj�U�7� !Ϫ�����/xn��cZ�MJ�eq�s�Wv�$eU`R)�y���fe�ЧG�}Y�h����ԻyM	z7��9Ui$(��8$��N������C�mMާf�[�o/���Jp�-�+'즵��u7J��)�Ur*�Z&�E����B8_N7Y��*�TFV��U�W���26�3���F$�&��y�ڟ��6y֫|��L:���t'g�̫n���v_+���*\[�Pk��j)�p���&�_7]H��uW���l��؇^�f�t�U��a�N��}�/3������5�z���5�`��Ž[EL�$��}#�aӰ9Ӧa+y��wb5����M�,�W�dq��x�/�v�&�{սGe�2��;bԚ�Z�v�Y�%f�j2��k�W(B�)nw\n0���i��.��~�*�m��j��+�4ݍ+�4��ǋ()�œ]���t�S�X��à�5��T��[Uk�]=V�r��/���HMSiH��3��j���(3B�7'!k�n�i*�����*�������e�t8�9+j�pmF,�p87lW���f�3M�oU��;��#�ឤ�ˏ^/a�B�mb�+�}`��n������d.KJ��w���o�Ҧ�Fp}�w$�l��Z�6�n���ͩ.^v�Yea�,�����C���*��GVTZ�uf�&�0�s���c���`n��6��З8�cλ�l�X�A��'9/}K���S{��T�
��8����Ţ\�t+�.�S�(Mg�}���u����XW�ߔ��\��/mdP����)�oz��0Z&X9]�
}�[RXz!��6�*:�բܨԎ?Va�| :F�O|��}����N���Nqߡ͖�TwOf\BڨM�^�{/��V1җ1�-�y#��J{�N���ۼG^��z�M�߷��N���ލG&�|��f�Z�q�.�nv5�z�[��߇[{9��cx*C��9��3C��v �ס��0�
z/)-n-��z�y�0^n[�K��c��ʞ��A��a��M_����І3c]�Lc�wx������
��klt�mV�y�^�A����]p����&R�\1�	���y3�̻�"]1~{S]Cg��R�iZ-fr����н��OD�1=w�a/:W�]�GYV�^;�����;9.m�gH4uo,�X[�`ǜ�d���SUhu%R�f������ ���7!��E�n�V!�;υ�t������U�.���Q@�&�7��5D��vPsE�����?}^��:�`�	��'��j��\��7��H��'�;�'w�^dl�W�A�=+����A	`R��QAr�����J�&��԰|��c�|u���S�g��L�بv�)*��Z���y�L�&ݡ���{��V���I��}�mް������B��D�[EZ**{�.����~/��&�׺��-f�|�k��x����8'r ^e`�Ǹ�*���2/r�ۚ[YJ@:���{�^_�u��h����2ĵ�^�n�5�9W�vT��b�E���lF����-� b��%��/�;/���j�U�
��f�&rՙ���k�v�����
@�%u�������12ڜV#�ʱ�7J�u�Ǘ�Yx��]ų:R~��yl�r9�JT�cmA3ʶU�m�{:��:�U˚D�Nq��f�&q
�v2�	���g	n��ɧ#£6�o}{I7�gmC�Z��nc)72�L2,��3�WE&p���@�0﨤������.),؅ah�YW��ip{��ϭm��:���=ЫU�x�H��'¥꛸��y٥EE�l�#Gl�;-��Z�:�Y�n#@�:�G����h�!����ir��NЦ:뵺�IY���+�azr%pړf��_B�U�����#��_���VL�eฝT���I�t��p�ñSko�W��u����U7����_D5�f��k�f���w�ҧ���&�	:�|<<�ג��Y�'�z%��U�>�2@i����o��{Y��	��U����4�J�*7�DGD�v��7�AB�h{�qq��W��f�3j�k�,3|S.p�=#N�FWw5g|����cd}�A��Sʧ���.�א��Ɍ�Ԯr/�j��ү�]��=*1�S�ʤDet��<�k��Z��JH�yG{��]VϺE�QpE���
?.��^��^���	N�p�W���XaӵܡlO	 Z�7�ѫ)UT@���\�#ca:u��_�T���q�8�J�ws���]M�=[�И���x��E3|�?G�qw��M`딸h�W�0H͢�j��C1<mL�#e�a�,���T�#��g��`�˾�He�K�\��,�Ih=��F�5�Q:��E�����gvbƫ��L����<�術{c�E������b` ���꺊���E��j� �.�#|��6�6�tMi.�l4q��C����=�(�š��h5+�?�mq��$8+>�캏�)�5������ZV�A���:��e�M��ph�\W��U��)�������f{��b�t�!S��#y�g^)��a��hK>�t�9D�;	�z��͂f��g�ƙK��1ߝ	W��vf��S�D9�*ؘ��^�B�L,�5�E�����$�D��ʃ�
��۔�ess�=X�������� F��|�vy��b��>4&�:/��*^��7�9�8)���)��}w��G�?-<F*�J�<:���aN�>���tl�bz��f]~:_U{���y(��1�z�"�󰖡�t�V�J��F��:fA�w%}\F�6A�m<1�Im��Fr��l>��d�y�bz���O���J�"�� 4��'����g�k�v��n�s2,3L��f��D���q�:����@�:�Xu���jb'��ۢ�v�c&jc�ؤE�%��N�5��N��xK�R[6���-���B��`IO�IO�!$ I,	!I�IO�BH@��	!I�IO��$���$ I?؄��$��$�	'`IKH@�l!$ I?�	!I�IO�BH@�rB���$�Ԅ��$�	!I���e5�'�+�)I͘ ?�s2}p$������$ͅm�hTJ�kZԨЪʴP"��E(�-������	U$�6l�MfնTֶƆ�6Q�he��XM �0$�W6���k�钕)S`�Z�+�d�_F�j��s[0�I!�@P�Y�J��]���2�wQU��֑-�[1��R�c�V�)KvӲ��h.�USmBhj�h�R�Y1D�cKTV6e+cE/fI�5Z�ART�Y(��آ��e+]vرj��  ��KMP���#-��Wcl����S�\wV�Mf��N�o�=�bP:ڔ�a�K��j��ʅ�mP�lkkT��dU�[i �fj�����u"�@g�U�  �  ;�v��
��{��a��V�M��jբ�Ĭ�ѭWK�-�j��&���v�\���u��tlٷnwssJ�n����뺬�j��G=쒝�9
UP�R��5n��|   ���>��&�իnڶ5�d�.����B�YT��[c�h�Xf��J�6����v�m|���{Ox�
  P^��z
 � P�wz��C�    ��H�(�  ��  ��� h4Φ�@ P�hP����B�
 СC�A�(P�n���ض������hT�%`D��P�݇�{����oj���)I�    ��Z��eR�P��� 
� M� ����Al^ܠ钶���[Q�(Ơ MWT�jUIB�U*�(-Q�  4�UPm�h RԘ�Wݩr�Z �XJ���
H�M �V�jB���(Q�d�*���N��$�    }�W�RE�\S@50 �0Pփ`��IV��NQJ��B�٧��u����ㇽΊ֭����j[j��z��fJ�ɶU	R�٬m�|  3/���N��iVm���VT��:��WLt�eu����c���j挕)f�ít�RH�ܽ����՛���wvV� :�]-�m�k'�"�f��  � ���uvwd�v-%*�Ӥ0�hU����"���ws�K�6�]՝lm��g8Ul��M���#M%�cn�+F�;�EТɭ���U����RcWӖcHHj   �  s�%s*�j�7mV���#�w%AQ+�髺�];��l��d�*�%��4��ˠLݻ�����+J��m�t�iU�vmk���RR�@ �x`�)P  ��&)*�  )� ���d#@��UG�� �&�ةR�  �N��O����S+�R�J�i���g�؇jT��Mf�+�pN�2���N�bi����o{���c=���$ I7!����IO�$ I?���$d! ����e������|Vr�H��j��kW��B�v��t}���\e�r�`�a=.$�������?�����L_�@4��_X-�6�����#L�����&>�EX�K:��O1]�I�_5L�}��*u�t�I�g�o>ĒxA�f������5�2�g?����%4��$��-T���yM3��z�x�N�{	����>[8�O���;޻�,��]Ó$��d:^��d�����D+Z%�����e��NeeE��P쬶��{	|GB���}<ټ�N����FG�>�=�7P)����F{Z���u�ݱ�uںO<�|��rv=������'�����)l�F0�:���q��i��h5�9��Ώtb�ua�e-�Ge��f�sC���v��D�n�Lf2�sʢ�ΡP��T�����[�Ƽ΄1_�cN���}��I-MƮӞ�l�,z�iاe���0b�Mf��U{{���*��p�66�t������z�3oQ۶F�_f��þ���O����s�Q8a8r^H{��{���D�>�;�B�y�{�/y�4�l��%S�	������?N^g��Ϻ.;�<kJ,;����E�v��^�5��7�f�c(n;.�-�7������8[���VW����%�W�z�ܵ��C�aZ�j�;L)��t}<���8���uO>o9�a�G�$���˯�\�Z���6����I6d�*w<�!�>^~㽕wK5:��e�j��|4�����cB�����Q��܇.��پ�;�e���7KQ��X���%���U�;�˩�+F+�Y\ �$�ݧOp��CbPA%��.�l�o[냑�s%��E�x���i�Z�.l�sc���N�9VPKWX���}�p���b���I�w5�ޗ��`��Ϗ�j�<�k���5B��y˺u�o��DX6�i
������͗�׊ޱT+���^/�f���~}b�n,<�n�����-�kQ����W�ﹼ�I�
�懯�����y�E�E�3��g��P�K<�]���g��f4-V��5�Ѕ���t�%���	c�ۢ~�!����v�����T������;}n�#��.k���t������x�Ϸ)��*;�m5�q�U���VB��ov3Ƿ�H�8�m�3;�U�y O�i�����#�d���K���.IZ��iׄ��W�`9��&���O�{��4��}j����;��0o^xh���cv�(=�!��x`q�����e�L��<iX������ncw�������DOJ�N����{w�yu/��&T��x�W�C�8��
0�F��oC��<�]�gTS路�ٗB`�Q��V��P�]����Z���
έ��J�\�b�Iޤń�7��'W/W���J��E�{�Ϝ��N�֪��x�U���	�GU�1^}�C:^�{Ǳ�v���g_OmԱ�oj�ch/�V�6���qof����7��d�H��"���\c�֠��x*w�20�j�(��-��^�e>"�2����۸ar�>μL�hUd�s�4��}�h�x#��;
=��=�1��[��˛�:ב �U�����	�.��	�Ju����y�44����WN�sz��/45I�Y�v��q��rPJMN�T��6�b҇7�^y��&x����{ܪ��x+�}o����;^�t~"#�oww+N4�y�z�f
:�ҧ�esݽ�3���:����ߴ�t�"j�a�Ǭ(�̹��v��|�JwO9r��O�v1T��T}e��]�c��E���ng���pэ�����t\yCZ:�wՙ�`������e0��h��{��_u���.J�Kr�v���/Q86�e����@>�X�U͡��>�>�����#:*|��pq����l��t���W���Z{+d��$�����Y�5����8y� �����<L�e�tJ�����n�5���0	��1sQ��Em��i����,��胺��c��M�A=Ī�������k;�,<N�UϤK0ӗ�0�GI�u�3^Q�Eۑ��'NSw}���ܟ���%}����5Y��!I������ؙz��ǹ[Z�����`�ۓ񸘇,���Ά�&;�}����~ܼ�KSƨ��7�G����v��{�|쭸������X ���b+v6cyA�{��ޣ��$�
�{�;3�Ks<�*OL�'V����}�M�k�R���hӂ��DI&�S˽a�݋	�������X1=�y�Ӭ@�>�����5�M��ܰ7n�S6I�����o��W؞ԫ���OQ����)�4�ǋ�k|���u�5�����z�����ʻƋ�wo{'���!�unQhu�&��0�qAs"�Lx�9�����LZ9���w�+�83T�'�I���,f�~���v�$�BB�����ܑ��<�H��y��{���w0����\�w����o�q��\�T�z���z���O��RLK�fe�^<�<,Ɲq���y֤H�Ŝ9 �������-;��\Ǧ��o��Lo]R��9�����>��ם�����A>O�����ߙ���Ϗ��IN�����Z���gE��K>�5;��=獌9�����r����i��C���@��bQײ��Vm~^��Q&�~��<�?^=�U�S�<g��Hv�b�R^v�9��N�M����&Q�8uY8w^<�v/�4���l��n�gژ!jؙN�o[�������]�>���,'�^������0�o���)><�Vd��K�^�ܯz�h�^x����Ȟ!S����ܴ6�+���3��20�$�6��8���O�]^I�sH!�aX%fR�J�qw�:Ai��֞J�QE��Rw^o޿�)���FW�N\�_49<��.�k�	')GL�7�f���q��⬏ǍyO+M\�S�Ӥ�&4n给^��O�b�����Ќ2#ޡ�[��8!쇳��/g�k
������`�[�}N�������Sio�h��[�^/;J8dU�a�����¡�8Nrz+$�rw�s섳>�м���͌���\U't���Sj�V!A��j�օ�%ߕݽ&�7�Q��؎%4uBT���X��*]��39uP�ɝ{���Lt�R3ʱ��7�;lr���L��Oy�����A�m�{�z�;�	���'IS*�N[��\dy_`�����~>��W�������Lg>�4�ɾe���{���/���v�Y��ѽAa�Ա:̵�=��t�Υ�B��}�[^�.�`��h�9Q�
��$��Y�bw;驻ޯ����w�;6�ܰ�_gh���u=�^�)����ֺ����\��>e�է�wړf���Y��7aQ�H�����@���ɢf�#TZH7o(8��^�Ӆ��v�i|��Ž�H��՟a�64<vJD:Ǩ1�"�XЭ��6�|D�>!x��a��2#�^��25rXk۲muoׄ�쁜��¸<ʠΊ�����K�7Єؽ�ԥ0P�tA����7E��ZkZ;LZ7��e;o�m���˷hS�WFv(�v����>��v�c��<��̬��T�n���jB�o�^�ݲ����p��#{�?=Y4a5��U��#��2�՚�(nu�1e���o�Ԡ��	Ǽ9&N3���f�pC.��:��:{��n[�Y��gϫkS%�I�ޭY�4>x����A� �U��ˆPMC��Z�-�osq[�gr��������{��8ŇZ���C�{t����u������6�f��f�s�E�Y}������I�8(���^R����Շ��yWOi�gv����7h{��$�\�8;�,�lme��m����q�x�u��i��)���;�)�[���y�<�[� G�#�q>����=�7��׭��e��n���دܖ;�"��1&{.h��؟c�xw�2���/߽���̿c�v}ާ��9�;!D=<]����>�[m�f�o8�B��P²���b�Ǩ�A�Su�{y��9�����˺<�Z���_&����k���p�q����ge&u�)�E�` ԫV�.�])�ᘮ{��6"�z�ć��o�4&�ع|7���_��`jH���<��&�Y��i�ok��ˠ�Awp�q:uc���'�*����#0f<V_^��z&�0x�=�f|$�]w�-S��?{w�'��3m�Cu��Z1��ͻw���X ט�\���}�:�S�5>�C��{�{�C�m�,޷�<��1��^��t�Fj�ʝ8p=��x���Z����y���N�fm�5�%ɜ�k�B�D
�a��л�U����9}����0-�K���W<Eۄ�y���n�S����,�B�����{�7����W�s�J�Z�����{�'�}D7�uq��(��om�����ٿ����)P�*�޻-_��}n\�����έ�珮WR��eQ��zŖ�ދ�X��2+(�);�W'��k��b�`+u���u�1������jwX�=���/�5�Gt�NVs�q����䥣����|�S��c�A \AH�&mTJ�N()��b�\7��|��Rzx"緸r�.��j��{&4;8�����<⊫E��pe���ܤ��3�-�bE�8��<:�n�"��A�8��>�/��#���R��;�z�����D}��yT��Yf̴�%���!�u�]�)cv���ͤ(��� {Jf���?�wpeh���B�:����FbÂ��yGv/љ8œo��_.����N�.��<�;��t~���z+�J��k�̿���po�L�M�F��iR�m��0��֖Moh��U�����HEHւk��{=���:5	yw��h��l��E���x��}Q��¬Yf~�,����X�:B(HMV�Ƹ{��8�V���q���i�]{��N [`�C���7�����{��y��� �T�ܗs�t̂>�C�-�=���z�2	��~���
·��5g��˯C�w��ψ�"�r�(���(cq[D^��g>��_f�1�p�{��xw^<X����׻}�I��5�-��Si�E�1��Or���w�Z�ֆgG�Y�\`���FkMl�9��/P��xCt}AV�!��ǽ��{��p7"�� �{�d��CZ�M E�Z��%ʽ��:λ��߽�޼�bv��������N�n�p{�{`�w���]i�sIP�z���]i7x�2��N�ɑ�0S����vr�/��
\rxHG��>��f�����WZ��T��*�$�;	p|Zk�)��Js7w�����Ky�m��*L�o7����F�Э��ӵ� л�����ń�v�1=c��e�[�Ͳ�;׏��7O*ثm������k�h�6,m'Wy�*P��&>[���f�z�=�`%(�B�wt��#p�yJ�ǈG��)E��7>��	��X�jp���҈盝y��ue�h���ږt<q`�yOd$<�[Q3t1�}i�M������zwcK���D"ޛAýb�$����Q�ی�K5E{�ݝ����D�w�ً5��Zw��g������ׯ���{!SH�}����Nh�����ޥ3���\Tydza�t�=t�����&Sd}<;�BĈ�]��ȟ���gjvP���_"������NN���Y�Κ��	�v��<��x�7���w���5�y��]��gZCA��L��ٞs{�����:4��|9�ר_����J\=�1m�J�����a�k��rbA����1�x��x�z��fw�p\���(��ksp�
Ү����_h�|K��㻝���ɵ�^�i�WL�~���*�$�G�UcfMz\�ƴ�.��6.j$�}�΋�g���ɶ�.�Y�7V���P��C�\����f�V]{ůW�8�Ӥ��XAn���y���5.a-s��c؈�e�g[�F�7��
��9)���59k#�.5g�yZ`����7=�[��=����.�~���7�|��x�gZM%�?N�6�E�3����ߊ��<
�o�s]|��$-�����>�ho�fW;թn\<���m��%c��_�^wZ��n�;F��߷)l�E`&A��a��<�b�l�Q
��̺�_� ��t��Ҽ���N�.�˃�_~(�/oQ�:�[�����PPw�E����0��K���K���9#���a�Ӄ۽;2���X:�$�I�d�Sx����p:�������f�ϋ"S�{�\�Uڦ�<:�(-�ѧ��A-9�����	;w�1�{��s۸I�7tq�_E�]�N�:�����~烘4v�K\�p"�|�]��!��&�7�o_��{I�?�����[V:��N��>�r��*;���o�2���^Ī��6>Bw�~��=��(?%Υ�<���_KkF�cǘ4;wY(�r�k;k�$����Ů������t�5��A�9`Y��9�� �4�릴S�n��Os�n���Y�퇗n;z� �0��:^,�]Zp#�!c�r�[�{�����3B������`����-&T��dkw��ܷ:����Et�S�9�B;��e>�צ�������X���[dV�W ,�{Bض���Z��s��`ۼ���G9���_�C<�{���n7n��
�*.�E�׋��2���{����e�e�#����Y�	�}}�^�C�/5y��T,;7z�@�,�b���ø��6.1���ubfLѝ�ur�Pj.9�>z�(�O��6M�J�C��N�"�X�@���Һ��r�=��"AVs��&�_�%:�J�i��6x�aP���0e�ή��ͶS��6���vf�M���+9��VU�x��FBF�w)ٴ���ܜ�'�e��2��lTxyJ[2�5́�,��Ї�}���iJ2�=؝�B�j�%�*¹�cr̮��%�F-L�rxwn_�j�ʐJ�����˲�(�9h�7����Y��*�CHYxx��`�ș�0t�n�v�\`cNA�p4�ǋ&��rѢ�e��)�%�ڏ��Y�r`���奒x���m�7a�T�%8��?`�/|>?rr��J��[�����:U�<����['uV�H�\s�8���[��-��v$�����_|�_P�L�.�9Ae��J�t�ΌS�<�d�����%�_,ʹ�d��Շ3���eo-�q+N-���;���A˙W�2�����ohQ��<)}6����c�l���a_��b/{Dm��>K���or����;a@�'�%���x�[��z�R|N�<��9�x�7�*�a��:�b\�w%I��O
2�Xi;�i}Z����t��yRsr��ݧ1���d��Ln��L�
��iyxR�����	˹���y��drnn��bZ�e����¬X�V�N����S6s嘰�g�72Y=[��֣)&#�z�#d��I��=�I��lA�}vp
�lV��j���f�Vr�GE\�apx_s�u�v���t�N�kBs�����\��MWr�R�-?���h�\V�uK
���q��Ô�Ӵ&&. ���ѡ������Cp���Sx7P����*�8���wX��qq�׼ق�M�_�㎆cd�;��i<\�֖�aR *����[�$fZҮ���a����o!�<(5\��E��Wi�9���a4S傰8�sk��c��\V��˭����r�=W-�MI�f���kD���DS���*J���)�(f�f�e\��X�L�uv=H�9�Pр�>��V��2��{>2WurO	�z�p���K�P�qMB�VC��XmW9mE���@ʃ(ls75�w����� Q�{���`��j�{y_r���7+���V5�B:�|�g]28t�S>�@��Գ��xv>j�o"���o*m&Fg %7��%)�k�=��<v������,���)���F/�_d9k`Ga��b��G1,δ#��J��6r.�F�X�F�Q��_�0��[��Y�0��]�������}˝!�m3mE�iv��d"-<ͬvVVS*۸f_��Yy���νc[GI�ݔ�֦c�ޙ:��e��������k8���u*&�=ՙi`W3
TL%��5��w)�Gj�>	m�ۮ�%��b�e�%@�k���YG�r�)Ֆ�r�0WU�M�����|#�٪ܖ<����8�\���"���K�7n��1!N>�!s�v�3�=�I��(�O�Z�{�fS{�P��7�ZG�[��q�:�&����uȐ�s�Ñ��	ڂ�1��������P�8�~u�����/���O���̮
u3�v���,<o��êț+rޙB�x�S�+��G,�y��ژ^�5�k2�{��B����oN�^��Ss��q�����G�'%SO�k+'N�`���n:v:�ӖjG]�g$�v��p�F��� t��k]5ٴ�]���E4��Wm�z�Y��� `{�ӎ��1MF��D��n���&u[W�"9h0bop VZ��vv���z�8ڥ�Tz����V����(X�od�y�b��<�ԟp,�o��>k{�p�
��Br^����35�N�;�&���{,;����.e��k��}y2����d
�H�|ڬ�w*�1��2��q��m9JP.���Vk�{k�f+�6�VS�_i͊�ct��a���h]�Ct�V\�(Xހɏ'Q�f����fS�wZ��� �μi�z��R����:kLF s3fV�㹖���n�IJȱ짇���+h����5�F�%�O�����jօ*Ęis�ڐI��f�s�,df��b�#�*Z�t�3~�!�s:����f�x�e1�ܺ��{ep�.����%x� 4��P1ZVl8����<���:ᇾ|����t0�D������$���A���=��Ln��IKy�b;��̒T�LiQ��pSt��@�Klc77fR��b9d��T�qC$�D,��J�֐ZI��tk�k��Y����'�r���Ƿ�i܊�;����ӺoΠ8.��w�]8�}��4m�L����h�.�p��C�iY�>�B��Z���
�5U��D�\>(�m[��w�P.=L��5G�q��⅓�0����7�F����x�7:o0�.n;\�)��S�w����\��Q�q��"��:F��C�kY�ZW�E�k��TWMɼ�Yp��q�U�wd ����6�e���*�p=����)��`��|�(vl����z*^�`�z���y���F�v��Ix'Pj�k;yvˌھ�w:����j1�o KJ�%w�v�)z�\)������������/�՝�����o���6�V4�uQ�r�+�4��(��� 	��7Hu�#ʆj�Nf��Yp*��s/�̻ɴ^��Y��9�3�U���u9��Q@cV�N\���"�P;d�ۤPעi7c!���V'*稗 ��-ś���+�OBsYt�)"^��!���߬��7����&<
��T��Ӵ�VYT������@��ݭ�iP�9�W5i��`�J�A��])[r��F�<
�]�	�0�|��E����m�����5;J�^�WE 8� e�s{]��/��s���(�]���Ty���K+�:��*�h���^�U�	|�-th��$��s1�;T�wմ����tE�FF"2�5fs�����Y�C��/�ú��Wͺ0��iL��:�)����Z��!�v��[��kfF�����Rh�*�Mv�Ív�Y�側�Ճ���.�JWs"K�P�n�L��	���\��J5L^�j��V�EA��мN�m��[�e�����e�|����|n�l^\�:�����8���k��]����EЉ�]��e�E7kv�gJ�o4�3iq��.�O��wi(����7�Q �Ě�F�_ZI�L�qsk��̢i�i�`�7[�K��W�e�x�5TA(��n�WG7P|�4�6�l	�Z��y�k&��\�'b��u��G6�|.�����$
LL�Xu�`�]�^*׻���olcŖ�_v�=���7��+���k��2Y�*��$h�E�p�ʺi�V.�F�n�;/EIhx���ǥ�+d�������Ӥ¦�� ��Qsw��i���|7��P��7�ΎY��PUr���Z�iu�9[/��R�xC����ud�=vC��TOql��
�¬���:����:V88qR;�	�Tͺ��2̄���ԧT)\d�3T[����Bf��Eem�@�?��Ñ��y¿Z����|Ϯ����j��ԕ���-��>���O@�^Ĺ\}���`�]]ҥ�%��2�+:t�u-(V�Y��v��r�����|S�:��O{J7�1:�l�h	Wm�F�t!�U՜��,���b���{���4���S	��(G����d���f�m���F����5;0�5.O�"<:�]�ξi�4��}0�����y�_1�Y��)�][o�BY��j;�e�CT
�� �Tm��^7��o��Ϡ赲�o<.�F���g:���_h H(��}�]��X��0wW_�h��WY�A%z���,�+-N�[����ٝӊYgBZ s@:<*e�
����3
���Y҉��oH)t.J4�K��>��1 �t�5�(��|6	)���W�	jsE��؊X(�/��΅aw�M�|j�����!|�I�����l�g;�;�ئ�
�r�E��Fr��qb�|*�v& �A����w�b��A�esh����Q�˷�7�BS+����^a�U����՛H���+&��Z(�vI%�e���C ��we�2�x�ھ�����Kc�6:�f�Bo�wl-�����gQ�q�v�_WD�ܢ)�`6~��,gk�Rcy۶�3�!�뻌�;=��z��~��۶�i��g�d�{P�>��+]7�V��t:;�9��\*��.�<�O�4n>Z������ϰP����Jyf�~>q��S2��i�[��;�����z�~�Xl��Q���C��z�]c��R��6/U.���e�j�S��6Q�q�U�l�Oy��\UT��}�5�В��8�]�j�v��n�,��ٕ�Κ�0��S���[�%L�=�+�Y5��$�R{P�L�X/oj�;NF�X��O&;���Xzɺ�4:��l� dY�NC�j�N��]�#��ÛE�ܼ�>{�uv��84��U�K�ӥUz��m�[n��S�ʱ������E�:C��̄<w�f�nлIA6�Z�:��q��C$�s�YZ,�nU��b\dC����*A�`����ND����u�����]h�Pk�P�^�y=�48r�7�?9����4�Е	�b6���ՠ�i@t:�H�:y��y�zI|����8w��;�hM�����ݭ���J�u�B���IDbd�\��k��;�5V��gi8�6:C��X�] ���L�W��x�]Ù�\gl��N�Ob���P����O�E�.�fӻ����k�X�{�^Ą�+o�ӣA�=Q����S(Ӣ��։�X�ͥ�Lu����-B�0gS6s�o^��b��J���P[8e	R�_k��K�	��EhSJ;�b��E�@$s�Kc-�bA���Ck����v����AbI�#n��'�ޢ�p��{FBwE�XsCǕ�7���_T�5�GӾFf�tpUyх���`l�c�v�j�Y6S�K6��ޑ�� z.�8`�;v��U�P�Bge�݆�
82<���+mL��[�`s�)�*�-D�grҋ(.�͔R��{��ˮI�/�9V��pף����xqTu��f3����\�2���<-Z�ً9=Un"̤�A%��0�f۷/�ܣ�f�s���	�rį��u�/:^$���y�l�[�|.&�O;��4CW(#kV�xɓa1���^\��7��^����㚩Z����h�Ӥ���h���H�[�w:�y˯��H��&�s_d�2�vU�]��v�������v���5��Ö���Q�QnV�Q���Eq���ס���n�N�돮Wl4O'+�.��-�=�.�,D8�؈�m���A�w�k�sg8��]�w��tY�
���P�7��ƥG�0����1��*�_wdr�G���5�n��;�WX�(+is���5�;|*�Ѱh0����d�>�� b��mWR͜Mkp�B|�S��Z���_�C����P����{���f#�_7����xw�C��WۻY����쬲SV����M4ح���|�M�m�[����[�P�y�/�)���OV�����?n�p�y�:���>�G�7 xA��\շفŜHU������QZ�燻W��$$=���Y���J�ݳav%PX5��Q��O��S4��2}q��8�CO��MT�������..�t��৫�ʉ\��S���5X���3���O,Q�nvA���WF�mc�P�˼�]��XCC4���k�Μn��(U_"*5na�o1�k�b�������3�K���K���f�%<���2I���7�5&�|lm1�^��"�wr�t��0�� �hmU�#6� V��7oE�4��H>H&��n轃�4Y�Ɇ �x�}R�W����U�]�6{U�:�`k�"<�F���)Q���O���r�p��8�'j��w)�{t^<�L�5���o�v�i�4�����y�ofwXK��u#�K�42�1�GC��v��1.��]&s�V���A���7���YY�6Vw35R�d�o���̙]5աحo_W[]� ҧX��-�s+�g�M9�I]L�֩
"��TM�߅�z;��/"�'�CMC$`s�v�p�steC-.B��4޷z�̧��t�q�����h_�ٓ�V����ٸ৏0�W��7Գ���'���.!.���_Tnf鵥:��%/gm�����^5�n����=�{ytQ��@�c�4\��b(f<�Ea�N�#�՚�K�^� �h	z�Q�Q�G�΋I�Բ�R��p�қ��hv�A���BY��#� ;�U�E�p>T�����5�N��i�a�Ώe�������je�m��u��z��Xz���w�/7-m��	it|&��}������X'׾��x�;�A�z�g�Xt��B���;C0�{�rN`��q,���Y��mr��i��u�����o�����kv�P�ryC�#I[����[�$��r�Z8н� ���4{��{��L��>��H��1����"8�bw%�˼̜�q-��Nv[;Î�-$!�^�)]f������]��K{�g}�>�g�t3�Ш��]�!�3Q|-��]`1�U*Rg�/��A��-e�a�EӻKG=}��4�uқ���s�V�f�	SM�/S����.���x��m�fpzf=d��ī�.r���%��p2��߽���]��w�����[}��~�9U���B��;�A����,����=�&���m��i��3��� ��rv�d�!)*�(Y�&���o)���7�s�u����$! ���$�	&W��x�₿b�R��vby�Cges&����׼/^�oj^�m]�>h�E=��+��+�TӆV�x�ȭ]Y���nu[�a������;Poe'�� ��UL��c��F�"s5ԯ��qKz����<���p�ͫ";DT��Oyg�+U��[A�����GY��*��n�<]y���"�{�i������㱅	I��i��.�m3;�9��v�Л	}�< E2�_	�ʶ���O��F�DOAQC��}�h5���ՄP}{�n>{�����=8	�GA���:v���w���y��I��
��*�V��a��E�z^tp^s����Q:�ѓ%��Gu��e*Uĳ��D���	�$�r�f��Fo�姍��KYǦ5.�&U���P\����hk�܊#wWf�ڷz�K�>[�C��u��s�5*�Zz���:ߓkO�u���r�M�&L޾\�U�6]n[�#��0%�2ܾ�8LĒ]��{2�Lq���'��;�p|}>��A�32�`��4�����OhėS����^"�Ƚ���:��l�c ����3��t5�y{Z���M����`���Պ�I���X�|,goҞ�2�t&Gћ�u�[�� ʇEf⮋Y�5״XׄE۲�+��nSΝ��7�PDn��Ѯ`�2���6��'�Jߌ乌�L�;f<F�N��&X����uq}�-O|'a�����{��n��V�y��)^�in�D�)���F���LV;f�$���Bu���� �j�ٸ#��*�f�T8�7+����x���F�E��]���iN��}�i�Շn�j,�z����M���c ���yWd�}�\K:��V�c(��6kd�Ϭ�
Vk]�gG�f�ܢ5��L9�m�]\r�w+!�����lL�ִ.�=�GМ׃4�y�X�+�Y�D�U����[��^����-^�7���q绸�vd����O;�)�8����v.���WJ�BK�.m�ؓ+�'�ҳ�q� �1��{�osW\��9m֢⾫�B63T��ѳ-Ԍ�Q�Wy��a��J�i�ߐD����v��c$7�N쇒&��bw;�mG�C=WY:�1
��j��%g:�ln��)�#�%���s�[�v��7�7���V��]�kM|��D�22��3}:�y��
qn��g�뺾ut
�k��'u'	nZ��Tx�9�jq���>O���Z���\=���p�^�[�ض����<� ����b����Q�s��=C���`)�����$#|��= ��+�E�QZ/�_f�,�o{�ڶ}����G�2�^#k�;�4�}�v1Ok@���[��]\�wSY���%���t����W�]�d��낻n]s��%,��D���;���歗��Z8�G}���ã�#������=] ��M����^@a�����rk~��yP��.tj[�)ㄯ��?���+��SM��U+�\�<���)�hV�S��,$�-R�0s�����MZ2`gKl ���tC�<}��o�20OghZ��J]�RMkb�ݶ�_V�-�X�V�-�{V]�uc�������8֫5�Yq�5�v�b��y'
3�� �[k����ϳ�tp�H�6be�|���X�OPo�tȍ�@��>.�+����ħU[��L|UO�8��OA,H|����;���͘���x\N��k�x|���Mz�o�ct��Hl��I��M-��#��{k����o�c+-�&9R��L��LN}��1|�c���~D�ܶ|����� f/��joA�{Z����frxS���������eY��鲠�ף(sX�X��,�L*!-6�qAg:��'���t�����h��M��8G�ıɍ���[��;�|ޣ���'�1�p�/3���W"b}��=�p����#*�|Q�:�S:����;j���� 鍣she^���b.�^媏5n�|EK��|��q}N��V�F��j'�t�~�ݡ���L��z�f���.��ͼw�l�4ٱ���4<�¸���$�ee[W`�V8�08���f�Ӈ�f)+��~r�N�?��E�����m;uZ�`� 6�D�7V2�����T*u2��y�ϕLޢp/2`AM���sb6�=<�5xw�)���&n��w\z^Q�}���6�ʑ���5��}�$�J1h�*{�\zbOA�ғ+]k����X�Q0o_�؀6^9�gPB�Thp���YΥ�d��̚����e^2�R��+�b���-b�(m�;����ߴ�������v��p=����]bE�N��-�%J�C-2[|>��i�t۹Ac���vQ�9z�ٖxԢG7��kӵ�ǰ撸n�'SD]�nB�Bs�����p[4['�Tn�;�'qU��y���M�w.�WGr�9k)n����ش��F�NFy\��.�5,%mj#i�[��
U���Q��.�'<Xv<�=a��%��X�c�r��:��L��e[mP�q����2������js�(�6�������[Qk%������\O�\
s#8�A_�4�9��ow��X����Uc�ʺ��i��@>̉җ��O+l���U5�A�t��,m�B=�X�z�(�[��cPDt`�唲����G}��"�m�"M7��|V�V�	+���gr�^]jj�i�6͇��+y��e�~�ѕ%�CF�V�Z���m.��^V�Ր����%� ����r�Y�9�A+T��p�Ƕ[\�ŷWY�LBl�s*��p�o.����8L�'�[�v�ܷf�7ݢ�0nܢew4��=����J�ڕ7��yX�3�՘�(s��Z�x�/�ծ��2��^Β���y�1U��eL�oC��޽2{���n�AJ��tJ%���	�c{1���:��X�D3����V<(��R�����H肎��������&Z�q��lq=j\� ���7��ֻ$�&\noUшFl<�w^oDՍ.u��8ձ�&��d/0��xGCN�|�1l3��u�S�9eΜ�cA�[2�I8u:�ח]̌T�Z��[��O��s擗�����l�Ct[?.�hʹR�]��G�&��%�;�:�c)�6!]���Q|Y�u�@�7��̻X���&���e��6Ҕ��e��'H�X?i��G��+�}�Lu���̰��ı�60�k2��/B�6���9���w��]�8�s_V���&��S,:�{�m+�q¶+
u=��f�w�NEqϨn�w�:H{)r���q�{ե���3/��V�4qp�35�Dp����2vHS��Ɯ�5�@ҧـ�ui��0¦�ulb�Hr{�`��Y�	�8�;E!Vrw��hk��u_6�by���/m]�5���d={�&x������pE���^A]E}q�ǻ���RVR4o>�GAe�5Q,Qkq�w���;�S�D�ů+q	���4�.����f��YZ�[�x�"�D/��zI����1�AE�|��we�TB��f�JM��j8������D:_+w�5��ڛ¦_�U���h�ٱ����ل��z��������w�9V;�j��m�{�+mQ��r�K���W-)vX`�ȘѤ<���]��	�����u	]\v����R����8�2�]yN�Q��E���^t04`��ׇ!W�P�N������N�Wfl�ˠ�Kϖt�K��7o�*Y����<cWgQa�O�6�f���	�X��Z��k�k���&Q�ՒL݊�jp�y��.$�ƶ�1ϲKvu^ڣ�uJOA��勺��F�}zQz|�Nz#�i&oJ;�C,bh�o�+���
3ｾ�"G˪�]�uԐ�� Kf�is`�W��𭋹��H ���p�;�Dk��ք!�>$�]� BNY�����te��Uѹ��9��n����ܢ�f>�Ѩf�05�{��*wuTg8sY�n��Ntdu \V�&��ٵ�^m���)��sp���N)0�v\Õ�od���ջkm��� Y<GyXۭ�,���� �nb:��'MK��V�o5�pɨ_+�G]0�u�Sˀ^[�#��=�x��\\;!C�	[��:������Uֳ^)j���Y�0:�.�jjjq�[މ�h�k�u��k0�ْ�wW��>�Te=�Xx��>���+��ދI�f.(���u�Q��v���:'K��*YoP�To��6��7���E5�a��i�l�iw^(�k0�к�c�V�:Hn�'�h"���ht;��fj<O7��gN}�ݕ{[�v���	�Ы,
��Z�R�Zi�݅�jc��1ek���m�n�l;�(Q��HefX�R����v�d���R�
NSM˨E.����sUC-�CY���?"N��4V���[��j������79G�հ�f��*wh0�\�S3�d� ^��Ӫ�ց����1#x�(%�r`{+�}�%vr$	m���T&�1��#K�>�D���d��0GI��R�)C�+z�`>0ZL��4�}*�O�`� }hڶ��e��v�t48+�v]�G��������
�P��xRk�^�օ�e�t�cI�if�K����f�u�j��U���7��8C�F��΃�$�Rh�W�C����F͠�N.v�kl�;��;h�-ڽ���]����pS{��$�]��<��\�[]$�&%I�+�{�[G+���Y�J����/Ў)��E�b�_����E��㈭$���0�f�o)/a��&�&�uu�N�4�B�h�{(��t2��d����ʮ��6�U�`���Ldwn�v��֗���w�:h��ј:����D�\:fN��#�f.�����4].��x�����o�r�6�ޔ7:��ǀbf�R�]�8�v��(����V��V�i�t�!Î��Qu�*�#�.^��<�`�n��Rv����S��27�!$9�wǛ��n��Z��*�H2�J.{i���z_ܬ�v7ՙ��c4�3����p�fn�«�vo*++M:��'A�rY�1A��GV�S+0k�/�>�ه���t(�T�
��JcEgf������Z�8�R�Sd�e%s5�Jcg���@�6����A$q_�P�@@�S��k�|.�NBw|�:�\�Zq���Hꍔb�6vud�a�M�X�mfNv��h�ӎ>�Yѫ��q�x=N�u��KA/�Lɪ'�H���Ce�eJ���P�Av��1��O��:�^t76jf�vKmUu�F�p<����r��][��`׽x�o3o�`:T��C�Ү2�����K�ӫDXá�����i��3������* F�ڦ���S��:�:���%�`d��e���tZ���H��Dåno%-�u� ��W^3�;�T��{m�aA�
�|�"AӮ�h��F��s�.��Q��%��ƈ�l^�֌�Q뚯;��Z�����䢔v�*���W8�<�sr�<�!9�f�	�HU�y�{�]֤�Oe��&�as��y���R�񩫨ܤ�,�I�=�]8p�5t0=��Ҥ���û�	�!N���=J3w���|��]�h���.\!1ͽ����'\�C�G�K탴Z�z��N��B]��鯊���ݚB����h�b�����r�����f>�]��-�%�ܬ��LQإBu����u��W4M39���6I=y�
�#t8���si�H�,)��iY�Upr��YPi�
�;Z�a��\�	ؤ��%�fe�C5��&��9�[8�Z�����iua��wi�L�Z�vإ��E��2����O�b���e���y��Ux������aW[�r����w��-_q͜����B�k秱�}���c}��<F���n����C��\��gykH�96f�@��te�P�3�u�c1MMJ��]K��{��u��hi]�\��R�]]}݉�f�j82;�g�*��f'���]$�R)ھV�СzE�Ձ��u�8���G�3,U��ݙ��O�s���c�H�;�����v��D"WV�����m�(/��LZF��8�_uD�vnNN�I�RF�k�����鴨$�mҷ��n��6����!�U������Ɍʴ�b�=����x�sB������Kb��G�☻��_8���oV�0,��P��	!"��4��؇�9�=X�na��g9��g_I.5Ysh��W�k�ͺ�]I�a�ľ�O6�Zs�.9M�@?�� g7}��N����������q0�`P�%�ʙ<�3)�,����P��C���cHRI��<zݭ���-��S�GQ9��Qdö8�z�ڇ��џ�;�v���F������\U�mR̰�{���-��t�t錩��|�p4��w��O�)�ǥY2��t[��J�Yȼi���e���G<��g�� ��eon ��u�ڝ΀'�R^�7ؘ�˵�"w*j�F��ִ��|�-�t� ��avg�1k�GA����x��u>�PL]uڄ���+z��U�����4B|��I�J������q��v�%q����*������{� ���+��C��rha�	�H�܃e�xQd���A!]��?��|��AO�T����I�V�sԓ����m�)�a㊳�*�t��Vr�/�ǑGn��;;3PF�r�x��#���A��u�� �r���G��[�[Y�O�X����9s�o<�i�]Ȁ�b��l�U��xot��Fa���EoU�X�>�j�+�2�y��C[�Ur�9�$�y�UN�Փ��D����$6r���.g�q�&΅��ng���ﾯ����}T�hT��]d���|$�<t �N)}�^�jL��0za�J����v��j�-CY]AV��P,|��]�{����ٮ(`��q�w��oU�l܍4�5�ݔ9���Yӧwr�E����� �[{{v��iw�qT�:mE�*�m�?s�U�h� , :�V+s�eY�G+I�P�`4�p��ksWE`K��L�:}�Hd�Cg;_7)MU��(�j��y�Mא36lC�kn�n��YG0��s����5���[+�9���8���)�[3 ��HP�ׇt��i*
��-R�U��+�;��SXu�^�U��ev��Z�ӝV�'F+��ȓ"��*�����橈�c�8�0dmӮr��W��t��Ζ��(lNѴD��Im�`��ӂEu���[�������28�F�!�m�O�s/�i��u��ύ�$�������d�&������,4��C�2Y����8��c��P����E�k8�Z�?� ӓ�|3���fR+��I�Lg��l�
�2��fq�OS޺��KC�)R�č��F�/1;��}t�w7�+R/Xt�2,��s�'Th�X��v���7X�44�i|2ZU�1�iwH�e�����E*��t��|�k��-�+��LO�מ�j����vB4~�T_~�|W�ZxV���
�۰!�Çx�Y�5�/0�9�t���a�,�hP�ǳ9�L��Jje��s���kҖ�Uh^j�'gn��(L�C፷z�!;��*�[<��u#˻t"}��C��3���ff�G*�@T��Զ(2�V
��l�5i�2�����Knv���	p]����]�5�;2NL�Q�8�DE����)Z	mX�iJV�,DTU`�m[h���X�,����J�b1AU��D����%�ڶ�*��F��1ck(��-��AQ�cF�e���(�EF(��,X��A�[(����V5���AZ�QbZQ���"�����J�RҨ��"�TUJآ�h���A��#(��"�J��� *1��"�`�E
"�DT-�
�P�Ʋ�UU`����TEE���)�X�U��QH���#Z�(�I[
ت,�*�EPTTkkQX"�E�1DQ�ZX�#F(�1m�,Q`����Q��T�QjU	XPE�$Q#"�QQE`����V1eh��Zث�U��Tm
�Z�6��3����q���խ�J]��t���#��2Ժ׭�y�r&F4
D��]] �7���;�+6>
�`�� �M�w�[��� �0Vrwu���0Wf�ʂ��R��6+k�W��f����IeE*%���:v*U:s;L�p�ԷOm;��s�)����b8���S��3�ۥ�olA�s]:��h�ab�	��9�={e�d-�B;�.:�,4���u,�)�x ���腍G��$4S�/��8t���;��3zKQmZ�a����]��V[�⣓�c�g�)RO���"˪���JG�BnM��3օ-/����>�^H�j�l-;v�2Uʁ�ѐ�W�U%H�0���wr�][�R8v�z��Uϑ�L ��|\K�	XX�7^���*7p*
6���\T���n��k���N7��>�|��:P��FU4���	mP�
���3�|\^�s�v����R�֝�geC�:7�bP��r4%�DP8��LJ\T�'2�U����mVu��������+���`�O)֡k�Փĥ�%�"�+׎"�Ȗ�{ě�uߜ�b���w�T��aT\t�Tł�cC��<<|��߼�Ҝ�N�4iʣ�zR�D�о��,�oĞ�~����f���+�;ED#��jPu��J��^Tesdh�������ڍ52��b���ّ�(Ң���t����.Su57��Ahvv�=���Խ����]�dYE�V/��[�:b��;f
���������|�/��0<'�ޓ�E���´�O=S��w:Qc�����pT�lK4�i��+	���xv��g>TA�~[ә�6�ص�n�>�ҽ�Sc�ez�y<jꗟ�J^���0U� ����*��ײ�զZzN��"�~#�E���5�k �]���O%�c�,Pu�򨝬���(�쁌�p=��\e�q+T<��V���z:����V�a�sh�T���;�u6�����=�ᙳa�0�U��^�֮��R�瓐7^����
�vsJ�VC^Z������m���L`���2��}S�Y�]I��r��vT^��'���dAy}qMn�lkq%��8�y�,UΈ�L1���U�v��P���F�;�!�_*a���ؕOV��=�����=��Zp.w4OJK��t�UKnP��M�D8�#�%b��ef�캒+���c����y�Qઝ����1�����Z�	ŀ��>�j�A��յ�,Y+���[�x�u�p�K�W]�7�ɷ�u\\��9b��w3@4��CI�Y�Vx���͡f�LuS1M�)�O��q�[�t~4��38F�֮1N�ZA" 6�vY�����*���p�&��V��4I�{���Ù��1u�u�{�s�{'y;vB��&!#>Il\q)xѣ�_�)L��b���7�d^��J��+������Ϻ<&-�!����j�]��`������WY<�Mv��9�0�3	�=˸�6�!���=I��o,U���T�ث�Q5�����s�u��Q�G�3��ܤ'����B��Ďɮ6<yS�93ۈeI�-K2n�ɱ�I�������>3Ŏ���MF`�]U��YJ��*�묾<VTp�j^�ڎ�����Zq�S�ɍH�zI��I�]�@�-����ɢ��^�>x��C<ۡM�'m�f�̛Vs���k��ˤ�t]�g)NC�F[D3���L��|�;zI�&_�@ t�c�J�CS�8<�f5�3"c!�# ��"Ĕ��^q>>�u�����_�F�Y��tP����|/R�5~0b����}��奖<��N���Qɍ�wlJ���٭��H)�{��[�\jx��/J�}{�Ky�݉�Uʛ;��]*<NCnѯ=�z��J�����7��I)tXN�/������/�>������[Ζ�V�l�T����9�W-�{C��{Oe�uή�&Gc�^���6�U�U��S#h���-��6���H��A�%�����H��	i�	+j&7������Cg|k�.��m*���!��fW�5�E��5NM*�X��j�o���ϔ
�Z��x�>]�:ꊫ����}>Ga��ڠC��V9����x��� ���{k��]"n�ͅY�7ۘ��
Bn��Lh$��#�<*�7���QW�%��o��ާ�R ��[�����nÄ��p	Kl,�ڞ)�$�D#���+<9����f��ӝ��]�c�/�`;"|ܸ��H[ �M��ؾ�b=�D���w˺�����D3Y?.�5[����p�.�԰{��iC%%��o�zp�-�{~�Z4�Y��ɎVZ�Gf��yt����!ip69�pl��M6Υ��fS쐙�W���q��ŚKe�����GFW�	
�{Al�@�B�o7�=��oZ2q��
xiI?_s]:��Cxu�����oWS	��"��WaGL(�u[��-i;1��}�9Bf����8��?��:-�����w^4\�پ"�k�]��x�[[cpS\�<���
w���E�j*d2��}�i[�n����4j��,�m0�W�k|=���^:�:r_"kp&��j��8��i!�L�us��4�L��[���y[���X�V��D0��k����K]��.l$j��Z�a��ϔmT`H�!�!s�Np*��i����ب1b-�����oWA�M�j�In�]&�`�hu�jk����War�w"��l�#�E��>[r�'�(&�{�d��>ջ7�=Y��s=�0a���R��n����%=�/�
V��q�:g�U^-@�:!d�פ�5a��Ԏ����^,%�x+�棵u�u�� #��W,��f����&Ø��^��J����ԆX��Z
%��װ��S:&s�-2�yհ��y{*J�!�P��@wө�@�wSǆ)�xC�b�KǢ��އ4'�#:�^��nvx'�5���^�àvUt�R�[��+�p��(����^�<�1�LmrM��ν��v��Q�Gu���3�~�%3�*}�l�nJ��FiZvŪP�VZ�qѐ�j�{S(6v�gKy��T.�OK��!\�c,I*"+��F���
,,��]l��ꖫ���'
3�iU�v���q.���,q||�؅��@:;�PG��Tk�m�us���/' {�G�״�]�n��5ڌgB�4.���qp��Ak%��%�yR�2J���{h^��'D�#�{�_[�i�^����>^O}u�J1\xHzXR�W`�yn�x���(���nv�za�:�9�h�#�b�����R�t�C�w,������ �*fl�}F��I7��7��8p{�Cϗ	����}��o�����"��x1Z)gwV(��T��yg}Ro�d>b�gW��A�C�o��aK��/��<^A�����"�Zu#��,�z�c��G��3#�8�g��'w�0y䍧sBb8������osEGM�>�<�h�2�����o4S���N�Q`��f�S7I��V:�yy��و%�s�l���t�rV)gM�T����kT�<�l�4hru��:��p��J���ޫy~o��q_�=W�~��T+�)ȺR��d�	�f@훅M3���YzZ�7�fw<�ϲf ��[u��+տXkK�/�è�����b�5���x��W2z���.����<��fWz�fՇ��|G~��;�"ġ�Y䇬��/"���Ů�r��!�ʰL�����s[Z�,Ss2���`{_�Id,s��
P�tܼ"���Ӓ�0�ǵ�	�W�/W����Z�#3�/�:�# �r�E����r��{[]���A[d�t̳M�����E}��>�P
�{t7Q��-mE�f��\�]�\��-��s�29v�KE�_J��vy��/4��t@�|kǹ�9˺X����j�o`�2;���2T��A�i*E.6�(w:t��z�\=4�-r�ͧ{�f
RWJi��D{˔*9��\$��S�*_�gQ�b9.��:u�W�u&k.S=J���[jL	@J�;P�챽������Dht8A�y��@�5�
��/�ˌp�iZsM�z���<�q������8�g��(׽m4OO�:���Z��׻��,p���]Pg�=6����'�ɱ���q�����§݂�=�Q��0���D+��h�E���Ҽ�����rk����W�,^�@�<�#�py'7j��:� ���ω�:^�npJ	���������5+?���<תּ��Չ�Ǜ�t(Od᧖�U��/-��A
�~��)��w��ь�ьL���rv�'��{�k�ү�;��"^�@{��δX��y^#|�=\u�%�f��f����)Gą]+딄��x݌���8;��T���Y"��헴����U�s�ߌ�,w�ɡ�&�@}�B�C�$&�-\�eSղ�ݯa��ݰ3ֽ� �}[�^F�����88]?nM��K���mnr���o��μK�e�]�u���Z�)��۱�z����ff!\6��{����؜L�'�y�8�����+�C�8V.҅�e�Bv-6��L#ظ7�a���r��Wta���2�W݃�S틭�۸�\��n��ml�ٽ��6}I���ƽ�!�s�Ȱ9�Q���:��vlLX˜��[]�Q,̦�J�uIގL]L�K����,UN\�dj���eZ����U���)�ކ��Nv^5��X-�.�eM�a��\tߺ��c��=����>��}�`�P�u��4�����b�ˇ=������[I�H�^����}��/�oq�dW9zVNhɖ��������w@�����=	�:�߆�U��3Jl�8�n���u2�>wxћ�jMn��v�Ƿ�+�;b��3���}
�ﯱ��tUX�T<���k��9J{yZRr�<�p�QZ_9b�ͅY�2뽑
s��=��u��
�U���=�.��,�]=���`b�U�cE�R��l����s��Q�R��$��D+@��uq����i��ޕ	�vbO�p=nn'��=5	|z6=mˀ��r�W)�/0���ز���-P�
��rP�@늈�eو�*]H���(�4Н��>��ohPy�O��薘ɨ��պ�ܟׅb���B�':�[q>��I�䜛������xOB/�����c��9.���{*U�u*k3Px�r͵�F�۳2�j���f��X{v�k�5",a���B��T�j\��v�r�,����4������|NQW�k�1�R̰TQu�KyI�BM5�ȯs�cަ�N=k���}k�:�+�������w�S�[�;�v=���K��Jl�J�Z���� ��YqWz��k��kC�oM���s���.�-f���ch<����T��P�%�0��{+��N��Ⰾ���B�}�R�ԝ�X�7&��#4Q��X.[ ߜ���m��\'�SF!��|<�������n�}�]�x�x�N������S�]��Y�׷u$nm���Bf��J^d\DO;�F/�L�
t
5æ���9�~����*�V��oՊ������C"y:���F_�b)H�0`����T�!���P��E�U+Q6n�g�𩜬��:�!��J��W��V��k:�����z(Tv�QLL�bKݰ��!i��9	�w6�E,����K�hSx%k��.k�������Y�b'�lK��Q������Uꝭ��t6�s*ԇ�¢x@�i.�}�iM��y�xg��.��,R��b�ڐ��<����c�r�vR�f�S�3n�E��{�[U5q���O�k��APtߛ����ys��)�*,9��\Ƈ�}l+�q�@n���|��V����T�c�n�n7�5�K]H�sk���v8�@�p#����朑M���g������a���7�`-w��2a���h٘���qU��\U9:�{D\��*ɍ�0��4�p�=q��9��gj�,	��.(�g�L����)ϼlX�����]�E/-K �XҀ^�3�������ݝ#�n����.�җt���(���'�T��^��w����v	�z*#ܣ�|P����=�JԵ��\�K6!���dÄ�.��WT���W��T��<��E�n��˰uK��A��KT*^�!���F������H�#����hw3ݮ��^�i�0�jB�L��@%/�X����j���"�|�(�����Sn�=Dux��-zD�,�rgz��X>U��.���ў=*���DW7��(E��"!q�ێ�U��7c�_>����9�$@ڹ�r�o�%Fv˒��d��>L���m刪�b����Tl�{��/�J��TD7Ta� L��gX��s�X\Pң(t�*+��ѯru�
�Sp����1WV�M�Z��&�VDE=o�-=x��F<&�1M�79mF�<y��;q�Q �,G2��]�M�F!�6����oE�kf��d{�V\�b���qI0��-���qZ�����e,�+ff�J��`o���:�8��*�����^o�<t�g�U��9���gtCsF�s}w�wx+�B�Y�s���A��kw�m�O��ht�ȉC�Y�x�ۉ�^Ӻ�|+r,\�9}�vҷ�/qZۺZʶ0����e���y�oal�U:e,0�sx�@Tw]�{���}�Z�=�Hl��n�3����Y��X�U�z��s�7`ؽ����+@��y����\sU��qʐ�����ݢTspۀR&�'���,��]k�'׮g�t:M�}��'ҤJW�sj�I�k)l�"�{pmk�r���fAPo;�bw���nt�f�S"�L�$����ʺi����{[٦GW�$&H�����{��Q�vn�r�z����mG�R�/���;��s���.�LYS�B�sw�	�ݛ��/�l����A�;Fhc:8�
�7��Ѷ*��ك{#y}�������W�Z}�*Ɔ��8K����&(%b)C+t3y�������N�&F�����t��Zqi��O��-������Ӊh����V�2E��H�w ���+,f�Cl�"�ڙ9���-UjU��ű2��f`VT���M�������hi}�N�Y�0�� )p�Gv�
�W�ev��%�T�Wmf��*�K��\�ީ	��h��ᡧ�s������=Pݴ\\�	�Y�v1䦑�`����X��'4���Po��|~��a����p�8�tw$��Z���k<I�ݢ�s������*ͩ)E��_�ᚆ�p�%�WZ��X�$��Ob��m��!��)����/�OU:�"�/^-!hR��x�Mb�YԼ̏�JQ�J�	�β;������c��h�f���\�Ev�NT1�'	eY����KC��冉���2܇psB�v�땳�K�Y�_%�q/t�����;Ӡ#M�w!�<�JksJ��7u���wN�^|wiC[Lx��K;q|o���bXn��֗��uY�X�eQ)�La�J��RM�۪�X������#�1�#��������U6Bl��]ˁֺ �AY64�X���8��I�K�ȇ�d�tUT�
7@����F�MN"U+ߡ�K}��
7�]��\���ʢ�
�c��%ݢ��*��JEc,�D��է��=^ά��`�>�0��N�p�q�m��eOX"�Z5���\��ZTe��A(ݹ��f�^����'��"?"Ac"���"�F1V���J�1E#T��@QV1UU�DQ,���X�	���*�Z(��m,PX���"$F*�TUE�Eb* �"�eT�Q�1��"��X�kQj�1AQF*�
�UE,jTH��b(*�Ub�dTF��AX�"(��1TPYڢ�EUTF(1m*łĊ!,Q�TQFX��[A�*��
�E�(-��PUPX�֠�5��D`V�Eb����`�,TTR*���-`UbV�Q�k%h��h�0��cX��)ADIYX"��j���	Z�X��UF+�"6�QATDE�j"#b�kb2�`�(�j����)dDU��"DQ �Q�U`�V��R��µX[E�n2smP���ko��pc(�>�`>M�n���b��:�3e{E��W۹�m8`T�$�X�����M滜�X��G���hp^�N������ݣ���:��o�U��֗��@����TNn6,B�w^R�����FC�������*=|�-C�"uvr��(;�ז7흕9Q�.p�Y�#
@�44��N�Q���UI�����5=�q,5��9;}B�_`>!��vd�����ԾA�|�}	Z�^�ԬV\K!�K絰,kڞ2���
�\�:S+����م`�J��*�Y�*��G+��Y�.��/[��
�Gp�|]^p#�ӌGP|�{�|=�����}*�[f��U�ļ7���	Ɛ� ���X�7�_�͝�[�`�|�pW.���t���+�*�T{���f:�E��SB��
"�y�t凣n�&Ԩ\X���N�Ҁ��Yޭ�G�5�t�!�
*Ar��S�ذ��l�%鯌��(�Զu���Pgrl�<�#�.�A�4ݫ!e	�T�-�C[+���|Ūj�I�Ơn���*:����s/�XN�Т�Ɍ���
��Ӣ8jAZ��;;�^�*jA��2�����C�G����HSt���{��Kw���:���S&�}����Ğ��R�j}��L�+�9�y]�����3��r�
Kf�&��c�n+����R�b���욛�ф�A�n�V�.�0�7�2ܩ�Ti@zk8ʒ)�x��r߷Mݻ1o���L��.sݛ>w��NlG-%� /�frp�1T��֚��In�����)S��3$�%�n�[g��Hj�����f����ޅM�)pE�H@=��U|���+[<v������@��h��½�k��~�=���[���b�%/)���k��'� �W����|vPp���4]?[�мA��͙]|�]����0���U��hqG�ju�|��EC�`�>6gh88Һ�7;ͩ�)r�����]ciF�5�ˠ��J�CSu8ȨW��ʵd-���n*�1����ߗxf��o��v+�����u��f=@�S��IX]���(��i�Y�;U\�1��ܨ�f��w"]��zG���
Cي��Y�ʓҠ�@�:�~����b"��iMO��-]{c|���Qcl�+�
!�Պ�T+�f d(pk��m�[���uѻ���F����=Zߍ(��t,E��C��9�l�P�|>���]>$g�w��[��!���OS!mbl��6��f�Q1�1W�f�>�;:�ɰ�8�]6�� {kz����Ԇy����o1�.�<wm�Ne��%��9szaFAww�6;�x�.pt@���p�*���sJ��;��b�a�l�]��&V�ΦmAY��GK�n��wj��1{�j��ì>�!7J�f¬����
��S_�+;E�R��-~zb�	���
M_��rLذ �qV6n�N/�C�ҙp8�V��Q��� �Rz2���5�q�)�<��ĪIl"5�������b�p౜%q� �{��0)���mF�֫S���3U:C`O3`�b�3��"b��@���*�@Q�u�;o�U?%9ՙ��c��pưr�Ǟ��dX��H+�c�Y%c�O�7��ƈ�IV2�Mi�"Kgd�`�8q�|�f�R�f�6_d�̡�^�g9Ƶ�2�޲���h�o�`��VU�1�&x��L�c�E�D���Ū�tbλ_y�_o��-��){�_��sq��-a2��R����}r:b�l��gu�,�L�N���;.M�H��V��xl(*���wn�d%n��\ޚ���d��2`W��dO'P��3�Lm�ٵ,���.�*#�޷m*p~W%���%3�:�96^�!��v,6�R,9��g��E�=H����V׹�E�7wT��V��5D�"�#b�E���`�)^�Ug������=��r"�N/Qɫ��Ҧ�yJX�6�NT� 2���7��Z-#0u�ⲹ��s(Ps{\��mv.s�ad�J9�n��6ԝ&�"�$
ʻ���{�|���=���ʩf�������4]^>�^>r?b��u�=�7� =�� �/g��>,/����=H�K�t:S�ளs��#Y�9����b���p�/a!�;���e��{\�z����82�  ���	N��]Yk�z��^�k:O�{�Zɢ���Z>�˚������T�6����ys��)�*!��$|@��w�����n ������
|Ud�*��q\W)qJ���i�<`��$lAlm��ݭ8��bN���x��D)������̤o&|��myH�X�e�5����b���{Z/S��jU�]�틌��j��(���c.L� ?�������!OuX���[~���ͭĜ�]�D�^쎌r��q���Qb�����d@v��J��U���b�As���1�v-�@���/\�9r�R�>��f;#��m��j�eK؍	}Qr��.��S�K{�.�k��6��f�S�:(NlPvze)zJ��ز:�S��ֹ���L-?��`@���3���vi�Ӂ��b�n��	�� ����R�)�S%o6��z45^R޳�|�Ⳓ�-�1C��ys�E�u�9IV�����3yB�	\XS0ޭ�V	�عݒF4����[�m�iC�de=����Y��εI�A�#�J̿�^z/z�6*�����*X����)�6wb�h�!�o������L�a�{����}F�NP1>��nk�cD���d�IZ�Q���W5�\	><^�w5ޘ��qE%�˾ͣ����+͑���gC씅C�%A>[G(k5T3c�j�� ����Sͯs���_[�z���{Y�W�r�"SO��43���@����o�՘�����@Kr��"ڙ}~�[����D�Ly|�>���_K�b'��š��p�V<aپ�.�z�a�Ry��&4��3�W�B��T�Y����@�<�8��f�j.W�"�K���K74�͵���;{ g��=J�Q���8��B�3�w��cf#�ĵB�����>EwL�/�y��N�3��g����.}����R�瓐"�l�\găv�p���:��ެ>���{���¼:R����γc�%}ScY�{�R��e� �b�14�NFWF?��n;�*4F�Q 9�>�wL��\��Y�޺�hp�i̩�f�U�pS-mA��"ܫ<r������^j��3B�5m:[�G2�ς����<�}�c�R����%�.g��Δ�u�w
�gEw�jgm��U�;)"8M��������릩E��4�p^�h��K�5��2�GZ�J��>�����}�֏���q��\?dTꞭ��ޜ�����ʫ��6�%	^[�>鴵=o��!����T\&s9�ZJ�
#ng���<�ˀ�Zꊮ#:�ַ싧��o���=�W�Q�M3p����Wf㾍�!�vGeL
y��Sw�8�zmZz�V���U��	�q	DD��4Z�ԻN����8J�b"�z�]>�:\;���O�mwk�U�o6�k`Hq^:�;mp�;qA��^Y���`���y����ZUS�z�k]vg��EV��T'����"8:3���Q��8 ,�.���"nY21)N_uW���{^����*�)�����u��u��W�*œ��׶ժ	�E��S{|��5�ш��:)Y���qT��;�qO�u��s��N�oeE�xyN'��{ȍ�^g���$�-k.=aO�BQkk!Cm�x��7(Έ���@W�"�yW���b���eX�s�fzm��N��\�}2T�S.\�f���������+=�F]�&��d�Ԛ��uun8rL̹:�f�Ә�ݖ1:D��[�Y�Ħ�f&s��Jg���!�7�s�{�UwqK;fV��=ųR�g]uN�ɓ>v�>���:��� ��4�+WwF��8::N�����jM@n
��f�����ߎgv�:p.�f��'{2W��v+�M@����5+mx^q�rKd�32+�����Ę�>�����>7�/�̴qV�@�_�T�8ݚ��y����t�Ԧ]竊�f#S��/���8x��]8�/�����rԶ�.^{k�>5
�.rB�:΍(@Z��ޝ����h�saT�`?�˅Kw���傠^��:oض��.,9��&���ӽ�,e@��u����q�W��Fc_N�v\LO�Dخ��S}C5=��^��`�*�&hLwK�P��u�mFtwP�=�I�R/�0��ٸU�[��fʀ�IE\�n��$w��}˼�o���y'Q������_ri�'=�g�m�:��,7��ȱY���٬{���}��u�
}�7�3�sP7�ٹ�l�@�,@���K�}��4kn���fN͉�1����j�l\�����#0�N�j�KY�xBK7���{��C���ݯ�ŗLoD;oHG��*�{O7)R�n��!3�/o��Y��F@��e���
��6]�r��s:��1c&�ۗ��,�dl�n�[��WO�Z6l\�����@m8�TC�tէX�+�t^�T9���oP�����;�v:xQ��m�S���T�<�މ
5؇,W� �f&��}\B�2t&Ĺ��u��W�,Tν�����ǌ.��[*���"�}P��i�rA�2�3�Y�퐾�`��.3L��Sn�i��.��^���@]�Ӣ�h�����[ǹsq͊�?�V
]�������+ʠW��O�7�D����9��|Wc�B��/޶�#��Zp�l��S��<����O�b8��qQ}�iюh}���uS���9͡�b�82FP}��,.Pc3����>͞>J
�Cƥgy�򺝽i���|��6A��%9�,�f��iB����K���L��C���[^���p�V��䈥I�Hn�I	�^�j�X2�lv�F�	�8�cF�Ҋ'�ݰ�Q�xB���C
d*"�+�^�Ti+)���^��
��u�د�fU���6z=A����9�t���x���~�Y�3�q:k�.��hp��|���7��<������M�dbf����s�ί*MpU�i��È�/�%�`-/���1�a��:v86y�^nr�u<xS�Td�'�p3�\��k��4���D%;[��lh�+�V�q\W)qK��8���.1��Kv�]��q���4˒x؞N���FI)��'x�?g�������f��VLE�����_g�5(��ݶ�&F��|#��y#��j�iMoZ�aKSo_7�E��R�6u	Z�� )d�6 |=�{���������o���8�P9�%��B�J�XdTDW��Fr�B����U��N)�ԕ����䭀�	�;�Rm	ul���iE�G�5��D+g���U"0R��)�*9��qM�0������sx�y�z�T����TtHKU�^�!�!!�K1{���B�A��Kۘ��f�X���i��$$zg�K�Vx>�t�y7�(׹��4kO�m!w�G}����Tn��R���~ע���T3���^x��a��}&�������zv������,�-�!
�`��/M�����K%�J���y3R�i�����>�ɠd۔=^n��	�:��B��d�)���(1�| �V�O[w։�Ab/��x�,��	;wS�x�����[��aJ�[-M0R�F���rw
�gvw[/(�m����K�Q�Jd����A��y}�>C>ȩ��/��`Z�x]���7�1��������_U^��3���{(CS�g9i�T5󠴸K�2��Ru(��R#�����N�]�>�Y�
�Ou��*i�����T49*�9�?��m�M}`
jk��M*RH��q�$�լ��Ecۚ2�Q���Ժ�=�)��(0�/;��������)��Ӹ��0je�8'�q�����xyrm���[7�kf>�8�����6@�kJ��ԬDNo�9���Ƭ�:�����k�ʓ�>�ƍ�Gu�����a��
ǋ�e��2�Y�
CJP]������+���|��fcGf�tF�N+�N��U���X7�N
��R�\��	�<���E]a��es�s��6�z�w���1�U~p=�j�\����G:}*�;v�*�B|7��P��uԱ�lל)u{~����７c�d�r%V���v
4�RJ�J��.���b�k��5����i��cW$��Y���ʐ�X���3���|K�4�T�cS���7*"����{�ͭ����!}�1�����p�$���䧸�1��6����.�1U9ۤ��z�u�?��;s:6�I����
�eS��P�`X���X���;��aj}yvs��̥V:�8��5�J������n:�kt��S
<��L��-v�*�&v3'���*K�o�-�T��7O1�@H���q��E���a�{S�X��S9c�����-^���v�̱�f����,�%陚)�u�n,]atȖZ�.�.�\u����6'��y�!��8�w��P�=y¬n������F��^|�=W�{�Ft������ȱ��n��p[�S�npr�����u�Q��.7T�o˫���w	����x��ډ[u`�.���Z�Xj�*۲�=xfmv�7�+��pRy��@�MY��nH�����>ge�@��j�gJ�b#m�ԫmHM|^�Y��d[�+:vj����[L3��'��;r�u�� i\����\k�s|CK����gR	ihZ���`���cw8)���w�݋�fǕ8��/���9r���lV)m;�0j����f�R�mu���p&5fD�^{HW=Z4/��B�����t����J��W���N�UlS���-��kl�{�7.�i#�mC���=A�H7�W�l9�5bhc�w�M�e��x8;׺!�S"�/���ؘ�rDV�Sx��鬚���s��= Ծ��w �	U}\�[���#S!cFX���o�i暳a����x���5V��U2tE�-BZ��*��>Q}1}�7F�i4�"���kx﮳.���2��ծ
���z+���B&^7�oG.��*ݙx-*�ãբ�a����*B2D���oo FJ������R�f��m�B:���U�Ɗ*`�CU��{\��`z�zp�O������������P�wI/+-iT�~y2��:Ǔ2m��1��]��qɥ����X̎VM/�)����v����p��8��U��l��s�4��b��&э�wۗ��ˈ�iآJ�Wn;���t!s1�WG%�`<�$_c��軇Q�վtw.)�b�;%�{OV���.��f����P�{@Á�un�h�M��꺾�"����u�Bc��>N\�;݋H�+�J^ڷ�'���T[A;��4,u�\�!<6�&T�%��T&�H�:�9��_P���P�ǔwh�)��J���)ͫ�Kh���0�\�u�ϟY�	����PÙ�|r��!�v?n�g���^�;�59��C�x�.�|]�-��5�\|b�⛢6�kUݖ��8�y.��n��'1-Z�e���s��ˇ��,�i+�N<b� �yxt�x�=ʒ��e����TдU����j�M� k{4���Z�J��qڢ��{t͕<�긋j��܏N�WJ�NL��*�ed{9sV&�S|���#��K��TvoqT�[�1�\3�OXcEuf�`s��
!/�PE'��`~� }˙��o}S;�j�n.�'���|��Ć
F`$�.2�qe�7c���l�c�BNC.Υ�Kݑ�r�ur��X)L���P#��(��G���s��������Y������ɣL!F�-V UƓ�M�{z�{����=W�,3@��v8W6�LHtG��n5��Ԝ�k�a�z��op���Me�	S�f�^u��mE��B<�)�ܙ�j���tY�`�U�e��Ւ3I���<cE	тT�����%���KM�⮠Nt ���э6۞��4��Mέ��@`�A,-�_}����@��x�ym���aU`�*��*,U��AEZũ-��#""��XQZPYEX*�D��`�dE�ƴb���� �`*0QE �V�A`�֊$XČ�J�
¥UEP*B���D��H
�R�EX�*��EA�b0QD@D)
��(�a*�+YD��Q�*�
ʒ*�`�QDd���$PQTUPF	ڑH-�R�
""�TH�� �"iYP�"��US4*a�Ȣ
!+j�Eb����AJ�A�R*�F�*�����b�b�mKj��V*��E" �*����B,TTR#`TR6����b"E�YZ��DKJċ"��"��B
�E�ȱUbV���dX,QDDE�ŀ���Jت�¤E,X��Ȫ-h�,�*��#X�
*�`(��n'��p�v�mukݴ)T.��\ɢw���6�܃�fc��\���6=��খ��f���5��Y��C��'?{���*���5:���U{ H��e�}�����?
��)�����yA޳�& ��W�|+�ԫп0���o����^�@�Mn�I�P���dc����f��X��3��b�s�^��'��v�D��G:��mDD�:fx�m𳛼
y����9���T��x=��~k}g1v��.���*E{S�8�Z�Y�:D�m֬�g]�BsX�j �{Ȣ�yX+���|�5M|���<τ����4	U�j�~�
��;������=�#0�*���7�[T�b��`_��xq)����u������}� ~�5,��˰��o�`��pM6�u�J*�9ATf7R8+΋T��'4���鑲� "�@{yp��:�(�v��2��v�;��ű��}����}�����0w��=B���j؜8c��|3H����>z��uͪα����j�
��2n�j�%���֓?�����x0Gi���\u{R��d8�6��W��3b�X������V��,VbnS�{5�8.-���x��]�r�+�@�dg�4w���Ww�_\	͛[�QaU��E���G����N��9�	Q�AC�t��x0owf�r�� ��(�\o���} κR;��s����
���i���x{�ֺp���k2��a�?Q�06RΖ"I�1����w��הt��;g"�>yo��D�N����﫠;�9�R,-�)�+ǵ���Ё*������+U����w+Y��S�dj �"�!:�}&3�����/#N�:a���F�>�@(>:����j��H{��{xR�w�'�
xw��b�j�$�bU���ydw-�y�Xuj�����<��'t����[!צ���L�~r."�h_F׉}�x�sݯ��?v�3����q	���k~]�2�`�n[�c�s$�nn8@���+�b�BVU���B�[#R#�z�F���ɂ�R��|���t���S K#u:���E���ۙv�b��{�5�V�D'$���Aו@AO����M��w	�V�ɢ����tݕ
���VQ�h��+�9����Q��siE_�}� �� �"����NS Ƶ/N��vFgEbzV�_F��)8tJ}�g>~ڞ�q.���M�#����GT��W��l��v�1���:��M�s/���B��R{��8]�����т�3)U�>�Ć�7��T�ǥ��Mnz��[u��*���ɉ5�ýS�=|�����i���+�d'�/�]��d��D�;�Cm��.;���ghU]��������a�w#��{���VҜ\���њ�`�϶�>��"@e�����x_��S����L6 �����R��q
e����f�<����!q���b��a����P����C�:"�]���cñ
�x�D3�3���{��f����|q�BS��"F
�QWn�� DY�����\<�ig7�s3Q�w���T�n_a	�@�[�%E�'9W��Q��]�Jgc\{_ձ�T����M�ۨhN?X7F�c��`�<�®�)w���-]C�˺U�U0�<���P�[k�K���aR���ݬޘf�x.5uĢ̃U#����'\1��>w����>\LZek�b?����j��*
�[��'׮��=n*P�5�K1}7]Eؖ��9�ƃ98��t���;F�DBSQ,Aԥ�;�����O(4<t^�W�m�z:�4��r`�zK)��ՋR�9�O�ה�<'���q�beJ�zs�Έ�t�(O���M�<J����M�И�]��F��f��
���R�oD��,��N�P�/�Oh��f-����݀,�K+�h��m��2�IwM�&co!�0vô�M�5����[�kyW�7!g��)v
��f�z���b�4�7�_Y]N`̾k�a����t�6vCYf�i���D���^8�۾8U혮������{����[ŷ���&���BmX�J/*9����+:Q�JB����01�|+���k�y5��y��p�*hw���7����IG����l��)��Ȃ��e�t�W���L����}i�ćoN�&X�n
,t�F���?X��܏`s����4;�p���q[ u��Y�c���\�Ʒ���
A���L��"e�u�B�S�G �GB~�g�'����w{:�܅`0�n2�����rN�H�(D��B(��gMB���t����VqA-Xq=z����	g�e-B˪>�DU�ʋ�l�1��siDB��Nn��'H=��t%��e�d����jx�a�s�e})Jv��o�o�7�F�Ξ/w�Eϐ�LGs�|��z;�m��#��T��<�V�v�p����/ϋ�xB>)z�ӭ����n�yS�����ʗd�����g��x��o(\��CN׫8BG����Ȥ\�b����(��!M�b��������ϗ�ׄ���Wr��`�G�^]���N��qR�C��H��q]�о�=�p�L����f�F�	� ���Y�j�(�t�����y�V{��Ɖ�
����7�t�;��pb��9�W{I��A�Z2�*EQ8TѼ^\\l]wHl�����&:Ih��:�4��v-����{�v����1��/NDUK���rR����{�☀��m��9.C�uS�e�ˮ�Kzf��s6�t��Il3�JQ�gѡ�f����2!���~���Z�����J|Y�YMq�S�c���
��o`;j����wUF��Y2�{�sݚ:ޝqWÜU�"y9�-VȊ�1�È����qe���pfB��me��<���$l�"B���8pӪHh�����z0%kg�׋�9�_^��+�L̷��S�䎬9-�{낱]*�]c
�υ �7���� Ǫ����w��=&��ŷ��][�ܯ�۰��P��l}_Nq�>�1������p_u 8�M��Q�B�B����V�
�`������U�n�L� G�}2T�S.\�k58�qd���ý�0J#����+���H1��(��^tͼ�M@����k�{Sz�Lm��Ɋ�3�K���X��}���W\}�;�;g�g+�Hvb��n�m�<�|��g����!v=��̺b�Λ���m�'V~>:y���Y�]��[^�>�y]/�>/�6�EO3(�����l⫪J;DS����2�2�D�4�V+��y;	�Zq�ײ��8�+�L"�\\�^Ҥ�ZD�H��4��k��A�R`��9�R����"j�a��r0M%cu3�{����Dͧ�k�>�-�r�K�.���z��;��CI�>��.����< S��>��8�q�;�N�G�q��#x��)zV{�d~��	��Ñy�l�<(�Q[�;�Q�l�x@u홅��"�J�hJ�{`(ҵ�&6�ͩei�у�f��tL�ϋ�d����Red{�3�9��㯳����I�u�2������!�������%���*o;t�2���B�D&�"��R��!F�'.��՜<�)y2F��8�)�;�=��7���@�Krh���D�����5�vQ�-�X���:9�+�?)����ZN/.n\4������X��=�^1t F���5��=se���X�����sǲ4����-������7EG�9rB�0�����y�B �rv[�jTR����6�3d5r;�Un��N�Mx�d�S�\�+P�E�t��L��ϐO׻�1�e7�8���>� ��a��o�t�{y�ޙG2b�"�"|�˘�uN�WF�Bq�(����T�A׌�r�p���jZ@�;.�lt���S�2��9Fx�e���I��s�µB�ukh���BpXs`q�tw+���27PoجJ8��eX����!m��#$g/����Z�]֭ݾٜDD}G��:�A��sŚ����;�\bک��@�GM;�"r�"5 ��ՙr+%�Mild��)[�}�QI��\7M���W\`6��r+`����9�����
�P�̘nk���ld�S��5{BL8kA>̕맛@�C����F��`�����o^�w�����NO�\c�����m�v%o�7)y��>zs�[�Zt8ylO>�[�i�f��lT�d��3�	ATDH�6͆��tf����W<���3���}���X|\~�1�{z:�v�
��gg�_((���t��^<�|�b�^_�q���Q�:֡����V}ر	��b���|��?�E��f(y�=M��H�,���cԅr���,�8�sd�+����~�~<���~J��xc�+B��k��S���q�{x��q�Ag�=�eRa8�`s}�^��a��a6g�/�N�]�>s06�M��3��a�vM�L�/{`a��i�P^'�a���R):��=���u��gݯ��JβW�������6o��I8�|�f;��|�z��)L��R��`�&�d����0L�`6�����m ��6g�
i
��M��2�3�a���؟�Dv|�rG*��( �a@0��`M!R�!�~eH��y%'��u�(J��jg�ɷ�
��W�9��Lj��Y�b�X��nhǰgY*T�o9�$�+�I�sy�� 9!G���Fs�˫�(�X�V*���tU<�����N�y�1��9�G0��Ε\���>��zC��$�E.��v�,�KlSO�v־�;H�7���:���rJ�7h��Ճqm�Ni�vZh�[(�^1��1I� x �J\�g4h���($�+�T?%d��4��Y�>g�� ����Xy�C��0�g��2�C�P�{�`a���t���e�Y~��~a��0*NP�
½�L߻�c�+�gZ{��߹���PR(q��w���+%CA����HW,+<Ρ��<������,8��h|ϝ$u�l2�<�&4g����N�a�H/̛L'o]���*xMV�i�shW3�~�ժ�WA��Y�@��a���gRc�>�*H��M�ْ��Rg�:�t�fXl3�@�T���a����N!^��q2�PS�2W�`^\3���ޘP*n����ݙ�<��Jxk \(���s�~f����0�2�`W�>��I�Vy�C	�&J�L�Y��T�E�a�l�Nb\��+�n|Y2�Ԩ~N!�\0�G���#��U�Gm�ޣ����&�t���s)(|�p���oD�>d�X~?:H-@�u�<a��e ����2�Ԭ4c�J�~��o�3h(e*Aќy&٤?&��E���y�y���Lg�}��ܹ��s���sZ��}o�Μz@���a��e�&>J��a��0�v�!��}l8w8��P��\��;H,�%u�b~CɽR�7���f�;�&��j�Wl
�����
]i׷����I�I��a���a�'��9tf� �d�c�+��ֳ|��e�|�5?Ǳ?�L���?���4�(T�����'̛AH��4㔅fY�s�p �����{oAq�䞪���ߩWs�~~߶�Rm
�k>̟�o�
��J�
��ɶVy��ɇ/�i����`4��H/���P��}Ɲ0<�e�C�`�>J�4�0Rm
�]��������Ƿ8�7�󿹳�0��T<cx2��C�+��>��&�<���NI�׌$����>�r��b���_P0βT��P��i�+�4�L�����q� } �;���*�U^����;���o�i��yfS���a�@߻�~I�a��c����?!�g�t�`a�53�SO̘@��a��?0�J�_�ϡ�&R(y3��:z���~���0���1�|P�J��n��F%�zS�D�`��O|E��K��^~��bD^��tn��jBD��pʆZ5p�D�Y�mv����J���$��;���ʸSKEh��8"g+*�Y�������z�ή�ս�q�M�����v\���������w9�s"�DP�?�
��0ϙ�8�CG���4���,����2�	��IU'S�a>3���'����i �d�k� �aXns�2̳��0φL2V��
O�c�~�G���_�GL�?USHT<j�|�2a"���Y�L�%f]�w����ۇ�
��>>���R�`T����E�%z�����K�&�R���3���@���I��\|�tYsൎ�N�ShV;C.X��3���i)P<���p`�����q�̩��sA���X~;N2a�WGq��K������i��I�=��
E�N���	�9�/�����5��֒&r3�9L�8����N�v�Z��Xe�Þ��M��be��eC�\$ٙ��:͠���6~��Ğf�|��{��C���I���s�L�d�O��w�s���/��0��R��
��'%�4��V�~�3˨

E��u˦eCSVe�'�?8t���:�L�wa�e���.�C�Rq�pɿ���*J�<�&7�C.?&�������N7�}�k�v�}� (z���
����r�YY�0��1'R�VW�џs$�J�I��/SL�A`�N'S�%M:d������C�nX'�Y8�x��W��~�������5��ׁH�d��N}@�0�i���z�H.�6w�3�O!����f�.PS�Vh��J�Ƴ�ٜ���*L~0e���WL
��a�4)�S7�}��׿t����x8�8Ʉόܡ�K��	��u
ϙ1��wԙAH�C���{��Af�6~��o��<��Ak����O&Xh1�ˆzʆ�o�4��R�fu?0�
J�xs�����^wӟf��N���E@�G�.<�% �0�{4Y֤Xk�s���~tɄ�a��;��*N!XT3�cO����S]���L
ʛ��!��Lr���:`Vu�C��}�����b���Y�����v���x�ǀ12�jM�.x��C,��N&�L���L<C-C	�~1a�.XT����t�YSϒ~�1���VWE񉴘IP�s����&YU'��_�{[Ϧk�������(\�É ��3��{e�W?�ۧB���#c�a�&�:�U�>�DBL�s�x!H���[~�-v�m��9x}�o�n��������%�˪vؼYB���ȋ�GF���$�6Ҏ��r�<K
�;;�U{ݙK)W�xx{��͍M�����4�Lˆi'�8f�*䩟s����0+ڽC/�N&$��e"�d���a�a��4r���H/P�,1�L>f4o�օ��� c`11�2{\^�>W	n�l����z�{���q	Rz����f}�i �C�0��~��E�P��fv�̕���S(~I}x��)<�g�Lb����R,R_\$y��)��+�7{��~��]��cv��
�{�M.��Q��P:G��.?8AOO{��m@���3��L��
J��
Ԝf�?{�G��\�����R,��&й��L'�����a^9M�I:�aQ����]��}����PRp�0a�6~�4ɤ<�S��=���g��oVO̮�P�a����8f�ke�IU&o~��e �d��!���VC(.XT1�^n��4?�˝�����ǡ����2��� |���O}�<g�a%B�P]'�0��s�&Ry�pΡ�sؚg�J����k'�L�~`T�1���p��a����
E�ɩ{����d�����r{����}��������zN?�)�y�������a�E�:�&k�}O��4�R���:�z�`�Ƴ܆���M��~eH�>jn}��G�4�gY+���|���'����{���ou�������I�+8��kZ���)l�0O�p�Y��>z���X�'S/��u�>jJ���?��C^�Hu�AC/�8H/Ry�s�b|�!�������q���~�F�s�}���e�O{�y4�(T�ě1�i�Va^���d
�hV��*�PY�8�P�8z����C�q1�>dægS�P��e2|�Aa����{\��|����}�y�mϠ~g�*������6�_0��>M0��0�����ۖC.Wq�++:�g�d�@�VLb�=f�a%f\$P_v��i*E'Y��;��d���O\{�k.)��?��{<�>����i���w$P��C�{�)�n3��Y�/0g�&^�Rϛ�'�w�2�j
h�9������Y�m T��8��X(0���w�g��m�2�B��q���FLۣv�]x�k�ZZc��Tz����hQ��
xw��Č���k���W�aG����᭻�+�/+��G�)^����Jg:�9�#������V��A��F��6�1j�`Tzl P�u�=ds�Pb�9�x�'�<w9!5���ZWa�����#Ǉ��mx��׳��p^��U�ʾX��H�%-f�^ 'o.	
3����uz1�6R���Rd�3���יSq�Y�hG}�����5�^�����_,�;���ry� �zGV�����>g�ժ��+�K�������*��9��Cj�����Wni�Wï2�wP��U��MMM��v��RJWV����t���jۏx���M멲�������X:�EZd lZ(�Y5�kt����h��Y���������u���t�]f�s��tav*<��xL�b���(*Վ���;��fތ���ѽR�@f� V�fv� y�ķ-�+��oK��0��q�`M�a��͕�D�Vېl`°k��ڢmV*�*�˝���e�m���v�Yâ��Cw@�NL��$Ԫɍ��5��)�.�d�4�-8t��Nm9���s�g�U��TVSf#��x�ng��Z<�>���PKm6D��fS��n[����&�8�)�����c���P���4U����p�_C��p�vL�:W,M�DZ�C+�٩@��������e=��W7у&����u=�Q�K��gJ�׸k@n)�ص�l���f-��Ti�<h%�8�0�p���	(����)�f�K�m��;��gw"�D��=�T�q
���w#4��y��N^�Fe�opS�TRn��3���DH�b���Ư��!nl������5q���q
s�d���x�F)�l8�bX ���������k_=�+7e�>`�p�J#�i~��uL#s�n���.�{m(�����t?��C$���L���+vf�zQ�%��*~�u ���D0���1�@��F3�i�CYq.Lޯ�<��jD!�w=T-f`a�z"9p"����Ir���.Z�����0��f��EԜ�`�1]�$c��h"͜�Ksn����U�Ǟ�"]����܆�����G2:�KE��WKʊp�i�Wd�ǎ�K��B3Z�$�������NX��^��u5�:j2�h�����ji�\�n��ak�[tE����:���"V�&)ň��u����2E�(4\���<'�oj/ky�$5�N`��f�����[P蹨��䘷c������1%�XL�+"H2m�XE3
o)}ԭ�5�TG��y�b��D�83��ť�G��[�.�=GV/��n���^X��C�,)��$QC�UTD*��DU@X�E�������b�T�5�U���(���Eb(�
[P�QB�*��#*P`�UXԬ��[k"�ED++"*�IYF,�6�Ab[b��EX�K�*H�"*(��1A���
E*��kR*��cE��UEb��E���PU �bDV1PF"� ��,`�,b$X�YZ�Z�Qb2,�c ���AH���V

�������QUUQ"��XVV)���((���ł�1A���AEU@V(��Q��,EQ��PQX���(�UE���EUbȨ��AQ"¡*E������(,UX,`����AAV,b���cTE@DF
E"�ȱED���F,R,����}˽s�m�V�G�xB�W���J�b�V��D���c�xR�[L�-�c<���N��P�[��[F�vG��3o�{�y�����c��A���g�*�W����3/�T��8(u%'�L&��L��K��?��m&����pa����fR{7	���e*N�r�f9��6�]0�~�4�Z��q���W�닫��@�0`G���3)7��L��<���'�a �w�!�y�5{�y�O����o�����M{?�u_�I�*n3a^�*�{�a�Y9������c8����B�m��1��L{� P@���\0+1�ϐިu%t�ֆXq�?&��2�Yԕ\���T�A|͈~L���0�X�/Y<�Ap��V��YS���?�m)P��ߧ��{��������i&W��%H��N�j�Y"���l��9�L�%@�k�d�>�Ru
��þR.ӌ0֤u��PϬ�x�MG�� ��G�5��{s)��6���s\���0�j�B�+Y37�{G��e�C��'�+�+2\`2��5�s0��*E�y������4ɍ�������8ɔ�B��<*�ǀ0@��F��+�7�וz��x����A|'�L%a���5��L�`W�6s��i��p�eC	Xk�{3�<��6c8&��1�٘Ci�075�e��a�jE?�p�hT��7�^���r��7��<����Z��4����ݙv�	>B��0��5˄�a���}�i�d�|��{�&��y�~eC�u��c�}�*5'O���Ag�}"l�}X)
����ѹb���������������!��a���a�k�2��Y+3��i�L y*o�f_��L0���v��(.�:�AH��Ɍ�ٝd�?2Vs�
\Xk�ϰIP�5�|����ɳo}������ث�c#� z#�V����T�ο�I��i��)7�`��~|���S)���Z�~��m�C���e�_��8{9&ЩÿY�rʑa�߾�9��=�e�I]'X~��4�R��%юp�XI�+7?Y3�����C�\ j~��J���.�`.X�3�>N��Xj����y+�F�|}��T���'�=�Ll������ߚ�D�4�^�]�d��;�m尕إo��ñk�ˑH�찯����Kh��4��|�Q�\��R�t�t�ȡϱl1�49ef���.��j�][M�u�Ƈbp��X-�]��B���B�:SL\����ȼ�ȕٽǦ�`+�~ x �U��N�~��Z�&Ӊ�?��e��0ɭ�/e3�I��`~jO�T��:ɤ�a��bx�	:��t���-����	�'=M��H�,���t
�� �]w²�N�����v�o���g�f�fɶW^�3H,�*�0m�p�Y���+0É���e�&S0�&�� e�����ǵ�i���nc.&Y�i0�Կ��f3�0�n̡����o�WX}���;ǝ�����w��?��y"̰���y��l�ݲ~J�d����7�I��B��7�`��z��,���Z@_5 �����(t�pL�`6�����m ��7�c(j�,
�y�\:�����}�^����}ϟ��4�g�0���L�|��6}fi
�ro9�a��T�?FL!����gu�(J��k>��ް0��W�`���`V?�H���'1�Y�J�'^�{?�NM�[����M]�1}�t� ����y6�H-f��/̩�+&�˄��:����Ҥ����4��a�ݰ�Xq>eC��XjO�S���L�u+>1��i�$߽�����@��w^�{�ݿ�6��L}D}Eݰ�a���L��c�&�HW,7ha����<���0*8ʚ���:H,��eRy>L2}��3O�:�a��x� �d��G����˟����/{�n%[�àzk����RaS�pe���gRcf>�*H��MM���PR)3�؝tͲVe��0�ĩ�'��6u
��C���
���;d� ǀ5���������<��֨���~e�2_�L?&S�� ��"�~����At�����Hf�,
��Zγ�a>1�oD�m)_!�ł�(T��?!�()b\���>0�Ԩm3��w��o��>�\00��|�d�/�
���E�N�����4�̕*O?���w��v�ɤ�Ak��`8eC�Xk��T���B��M e*A��4�(m4��-�.���m�W~���W��>�H6W�l0�ĩ?&�w�n0�Į�:��Hf�;��4°�����PR(~a�.�����{�MꐮY���4ᇐ�l��y��l
�RB<:?>�U��
��	���I�X�Ӹ�"��X~�����؈����r��muw��'G4�e�[s>�W�G��[Ε����uMcMXF�x�y�[��1�Za��%�rf���]�	�w+�.����[L^�[و#z݋�G9ݪe��.����{w{k�a�ti�`yǜL�$���m0���a��?!�r�6)�'���a�
��Y��fY��0�S�y2�Y_fɣ����B�P^~���2m"��͹g�J̲i�Wz��K��գ��z7�.  ����ϳ��
��W���?&ߘ��L;d��~egY/��r��� �dR�e����A|���d4�:�@����f��1�>�L u+��~�D��F��_^Jxg���� 0=����0��T5�`��$���|ɴ%C���C�m���Ʒ��?2o���
E�M��3���u��L�CO]���,_0�u2�ם~�9�!���Fo�b��� c#� ��&��|��O���Ҡjo����f�a��Ґ��?!�fc�Β,5&��SO̘@����0�/���P�
¿[>IPR(y3pw���{�.5��ս����
*<�'��(|���ԅr���@Y�|��d�+�Af�O���~L$<^���UI��0��� ����a��wY�H.Y6k� �aXn�ba�|�&/�����mΩ�.>����>�boB]�C�m������e&P��)��u�)G�g]3���vk�&�?%N0��&0*O����O̙L<`T��a"ᒽk����|�ud���Av����{�OS�L�f�{t�r��!Xh��d�+8�'賓�@�WG��e��HVh9d��a��*nk��8��&�k����d���?&�*�8�Y�Lb�&VR�������I��� DDz {�O��a �l�5���v� ���/�'�,��\0+�T<���NP:��;C�����n�Ry�C��?w�6�_0�q�m�E�泿r�~�V�fn�]��]�᯽�Q��L|�G���
��&����B��+݆3˨

E��=�H,�5fP�Lz��������;�3/�Ax�\$�8�}��*��~L}�o����j����)�7����Ǿ���!�����y���? �aXk
³�Ra���VJ������M��T��^�Y0��v�8�Lr���ݲe�S�ެ>t���8�I�f�^�N��7�w�F��}$��@��:���V�5wԕ��(��]���!mnMK�]w�xRч�+�Χ���و��mEow�b��]N��ا�ssW�rY�(X�A�u*�{�����OHᘫ�����ՂN���c^�DQ �*[k!�v�h㳠��B��%�Y1^� ��d�z]����J��
������8�j��N[�K�7��B{��<=�\�J���5�߽���lz���
ΥO�o e�d����i�m �d����Ry�0�w�P):�f�~�+�γfs�B�T��L=B�Ra
�^!�;e����|i��w[���Ǣ<A�0��G��&:���$��`a6��V|Ɍ^3g}�i �C!��'��i�gu��I�NR]����釓i��W
��7_�i���v�N9�ms
�|�v�V�~�ǔ *�|$��'������O�E�d�5�,?!���L!��y��i��WnP�!��B�d�_[H)����z� �	���4��c�K	7�����CU&��8̝��a��,�U���~C�����Bk4�a�I�zā�u�	�L3s�k$�f0�&�����Xo�����HE��k���}�.�,�d��X�I�~p�$�_��m��*���,���`V��8�䮒l>�)��C���8�}g�S)�aqI���Ԉ��`{� ��[�*��EN�r�e�ۿ����7g��srԸ�{�8��Jܳo���u��%;��>U�}�V��Af��΂"ə�^o�>�쮴��e$4x#َ���m�S����k�b���� ��}b$��Yر�T���q��>�ƣc�^u&��[[�;�S~��h�0���޴����E�J#�y��l�����d�Y��|��+C}�V�Z��>ޛ��a���3c��b�~��\pC�d�8�����Qt����0`��֜m>�~ݨg�% ����Yod���)Y�;쬰x���������5ZH�ck��\�Z�l:� �=��}{��c)��b2zL~ �w�8�'*�#1\`����R;zQ#4�P�r�,v/��~|���gg����y���v\���ݑ
u=���ÉA����|TLZZ5�+�	Q"��T�bC.���qA�*�XY��]�x1R����^F�z���T
�]�Jk���HR�@�/zGE'+OFo	|{��.��(��'��\�;�#<niT��e'����V��٭�T�������A�;c�1��Q�	˒
=�N"7�;w�� /9� �����6f,)��!	³Z�ۺb.��ߗ��E�@�I�I�5z�c�i.�����̆�,�T��%�2^�r�Cb���U{z-ݻf�x�^U�z�5�Ž��sR��=��2vח��e�
qVi�C�CA���@S�맖�̖h����[s"+�� d\DH�N� (�ɝ�6�dRc��5k�蜎�T��NZ�S��&DYI�H�*�m�T��Bv�s�凈n��vC������n��I�Cڵ�}m�>_K����_���a^�9��p٩��g��o�h�\hVew.��Y�!�I�i��L�e.,�C1W�����;�7��հD�?ոyZ����_���,�\bR��Y��g��s�=�. Zj�)����C3�S4�1j�{���6zcT/;�":�Nd�%GJ���0$R.�uC&��&�|�k�f*�p�x��X�"��p�.�CP>�o���Nys�(T�t�����ji��CF��q��)�J�Օs��cf��_=u�^��q�\�ͤ^�YO�}�^�Ӎn�
>�����u�C:���O.g#Q�p���X׭��{�yQ���_.�k*�Bo�]�_.җ"��A�?<0�5i��ɜ5y77�ޜ�2>��:��@�J˫�:�����>O3�����A8֏.Z}��G���c��°��ނ��P�\�v�ٻ�b~��K�{c]���)pm$��ڂ�=�C��h_yK]���u7}��L��*O7r�P�S�v�n����:H���͍�Z���#�̻������<�R�|��3N�M�u<��y���(�gk�9�ܶ��{�~b��:��9;`�v,�k����8��Nc��m����o���rV�3#'�/�����b���;#Z�Rs�0�Y9�9��Qm�[�v<������u}]Y}�L��>�p�qL�M7˲�rF>���[�~�������~�5�x����S^����}s� �B;n��N���M�Mz���Rx�)ti�MS�ݎNçs�\����{��ϕ]������8�n�j�bmi_�#'�'�9ѡ��؋�H�� �+�zR�����\��Ow'L-�9f�oft��s#S	�S9\�	�^S��Z���[Eb�L��n��$�˙�un�'��J��LC���b�1�8ag[����ݼ�+Po"K�ܝ�YW9C9��@�B{�C�5S!�muì�p�+�%K�˯&#n�c�C�f2�w��2P��@�C<��[0��j������<I;���֚�,t��ܰ]�hj�nq]>��!�j3��]���(N�Ԅ�ݳR�>{�so�լ+l���)F�7<��Q��Lr������SU���{\s���P�e�YE��*љ�WZ��iv���EU��x�C��w���[���X�c{Pڴ5NG��Ƴ���^��R�O`.��u�`��Ḛ'5�x&u���>o���x���r\��{�v�;eD�;p�p��ʵf��<�,N8gk�?����f����}�z�Q�C}"�����$}�Χ�(�R��U��S�9ܹ�R.�s��/��=B�+�);�ҟd�v��r[]'�I:�R��kNo:qo8�;O8�A���#��R[t���kG]��I[�G3&��%[@/7fCt���e;		З�bb�˨]v�1�]�.�XaZZDm3ٵ����9�(r���U���@���Y�z�)GG^m�oNW�����NԞ���p>�����	�u�<��R�v˗]��e(�{x������to(O�:��`S�C�qeƨQG�d�Ά�gP��q��3nJ��ǎ�hY���do0���O��
ޝCWJ<�v�-�{�Ζ{���{�X���>�#�1��FľwnzL��Ė+Ȳ"�Ͱ7,]Y�s}W�xnF�����'����}s:��h�n�o�%�v�o6��w�����"#u;)[���8�mVu��"��s��%>��/�q���&�Z�x[f���݉,�À0:q:)ŋ�m���;�v6܊e;��O7��+�x�#wpt���
��8���$`������)5�j�g����+&Ԣ�9�\����	�c��f�V*��.�w3��W>]=1���J��b�]���@'��r��=�e�!n��9�sy�nk��J1YOԝVpŬ`�B�V3�<X�,[���;�
$��%�Ӕ뤩�v[ȋ�f�}��9գJڠ�8oűܹ���	gi��K�V�MX��\��ٞ�-�v��Vb�Lj�{�iS��}0M�y�����?R��� �%z8�1�V�zU6c������*ZT&�s�J�.fb2�����p�t�?ov���W�u��4Y�H*z.�P��|z֝qJ����M�ܼ7�N�7���v��N����!\�l:��󱹛T�Z��Jl���R�^��P�.q�=�hcOb�;�4��@K��G�2�+�Y�`�U��17�1����h�k��:��ށ	�u�.��K|���vI�^�b�WNɶ����,�ܴ�1ḓ�`YX�M�<��l��;�yJ���$W4(�8K�x,e�9z�>�3����l�ɮ�ue�Y�%�&5(3�0��(�]�e�W��������)Lέ�X��7��K�-���W��^�Δt����'".9�ʉ �7���\�z��uͦ�#+�Y
�u�umWjS�x1|��*Ft��s��9E1��S誵ݍ9#�e�u�3*��B�a]v]�,������pHLX�9ۑ]���J#��ؗ{4,rr��D�k+�L\�"�s�E�}>�pO8}��.�����-����غ�|ܫ��ښ܃"�:�}�Բ�7;\�Uk�=4�9�v�t�Xbg�K�K�,�`;ͪ���7���Ż���t��ܹ�9���gU�o�ͤf^$��H�QA�.^V����A�P�;s�ZQu;6E����v��)l��ܳ�û`�j5N��C]!�!��*25𾹫��׼�����_�36ۼ�Ʋ{/9Qk(C�z�>�j!�s�sկ%��*y�+pQ�ɵ�<���wy;;֑�EZV]\^9��[��uqQ�ܧ�#NC�9ҖM6�L]��3V��鳷�Z�s'�cv�F�FRB��+B��)����Oe�{�6���ƞȩ�Y,�ֲ����1Ѝ��yX��{����&�
�����T{���xa��Y��g�v��#�CHoXd��T�Hc�ኌ�wDi�X��mv�hZ�K����i��M��i�`6/�ڐ����O�6C��	ȧAP�پ��q�V)j�tb��L�ʋ+�m�<���:�Q��g"�G'a�j����ϳ5�#P1W"���ri9f�v�oU�7�Y�b��멂�e�@a2��UrT�@��)�s�+w4�*+��+utd���1鳌\4Ӯ;ʰV`ᩎ�L�˕u��'QGo�d).�
����r4Qi��a4�l�:�(Av�q[�j������;D�r8��k��
֕�h�J'�bB�_Xׯ�0nifV�GPEI4-�z��ݥ����%�ұ��܁6F�:�Yrƌ�Z��{oA���lrq�k�r�30�ɀٵf@j�̔�"�aV|�{�oXŗ�b�G�̽���7D��n]Z���c3x��Mg�6��~kpYܻx��9�҈8I�ϖ������%`wL�sGR�R㵟!"�0�O�O��t����}�5��u����'��} o�U��:��#{/3���kG$݁_kD�n��9m�r�E�ތֵ	wΠ��R��r*U�S�ۗQǼ�e�"o���J��@Yz/�؍=�Y
�=�1�zO��k�>����3$��0�H(�{�����`�3vv}�1{#��et0�.)V��%2k�3�l�Xg%K[�p
T�i9���컂I�jl���f%��է? ;G�(3����qA�	rou�"�Z�y4�m�{��2t�Z8�=4#®q����!s��ų��0wx5M�ҧV�����h�?x2Q��,�M�b�)n}�UxגS��@�s������P+�\���Y��b�&u;�n�d�!lj��Wa%�PE��2�?n��qxY����ּyp�^慜X���?Y�L�|�*���-�E�ir
�H4y�9L�n=���i����$J���L���~��Ǒ�a�^�^��v��o�\�Sb��r����Q�w^�f��.#�� Cs&Ø���k�vg�ѕ�Z��۔]�Ÿ���vq祼��PW��R�����6��I���V/9�hȟ����	�l3����v�T��|z��E۱<���M_c�jX��h����H �X�X�"#>j(�R*��"��F,TAb2
�aR)bŃ��*1`)bȠ��$Qb�@P�
�D�b�� ���QQQ������ �,�dDU��DTY"Ƞ�DPX��1P,UX�,"�+Q �H,,H1����F#"
��#j�R*ֈ*��1b"������"�EE��E��)TX�D
(* �EH�ŋ`"�@UUF
��ERaYUUH�ŊE��Q(*0X�(�	�A�URER# ��AE �X*0�V0PQU`��
�TADT���@b�(�(���E�U�Qb�lQUb1V(:��g�9�\o������9s�$#K.�m\���e9��"�N�
��"��~O�9��3B��+u�+;.J��Ɲ�x)�� W,�smW_��^mfl����zm��d�qқ�:�лY�V
�I�V���]�'��?Pm!EąS���]�S9;��ڈf,��}Ūm���+�jE�<�M�]����b�ع�M�e��KnD��3Ua'o�%g8�S^y���]��Ŧ����|wT[����-���ڪ�"�Z�n�>����c&�Z���B�Q`_�X܎V��G\{~�WtV�[;�\�J:�x$;y5�R�Wm��~��0�8���
�Y֜~Oua�he���G0��M����26�Oך�G:C[Y�SS@�[TT�V�w�gM{VOL)�g9�a�FUk%�rT�'�3i��ВmfP�G4ttV�;YbN^X��U`+��b}2�!�?�}^O��~p9*�ñ�w����Y��Z*+��3�q{��3��d��$C��� ��`�,��H��eA��|>D`O������Ij����M.Qynqʞb����=a��ˁ��:�珺E�"v�^WdͶ��1�\�k{�Ana�GZ#qe�%����P�{%�\s�nz�{��ԧ�ɼő�n�~�^�j����X��1��h�����*⫝̸��a�j-��<�Wzj"���s�{���,\�(�@a�]���j!:���Z��z��VOR���l�OU�t�{}��K���P�(�Y����)�V.���歽�����~�}AӜ�Υ�ߩ�3����(Z��֑�v�7���}V�M��\q&d�؉��~�S�E�4�J��̞�
��.J�� ]I�k��f��������E	|��N�Ҝ����������SJ֚�~9|���!����j�I�	K����r�l���aeTԫ�]ɢ��9QE����Ƿ��9��^���˯f4�K���QV�s;KMCѶ�T߹ʗ���Ѽ�[b�ʛ�˭-;�r����Qʆ�ks�������U%EpԦj�A�K��~��T��k0�L������΃~��^y��k��tm<�A�Q���X��l��zE悷�^�Ff��9��K���v��D�ua/6�A��.cVT�	���gn��B`��-�nqfҷ��nʎ x���v�tj��6iܫ�s�J7)�:�A7��U`.�#F�3�������9��<��6���8f�Θ�ϘI�.�����9���s��{�Kc��]Gt���!��
���;'��ɳa'z/��ok&�b�\��8qj�j�����*�:��%�ͫoB���Btlo0����nn2T����Z5�A��I�:��A�@_3�a��Yq90�-���b�O^Ne�1�piNo;�.��}��1�x%[�������rA�֧�7}�����z�+i�tsˡ� ��c�C�w'/UNj�ux��'u�h�L,�������pϱ��$k�Yҋ���i<7^寪{_m�`f�^�L�s'��oX#�T��OSdS�;]/�y�&:Ɩ�;���ҭ���<jnqX���J{q��5�W��ɉ��V��]�]����ܮ��Xz���+ �zl��b�GU/��*q:�\�LIGT�%ڍu���.����O_h�tю�֕��t	�%����[�Av��'�W���K��aZY��+H�_�ܽ�/�m���Nc����/�YdVƜyO�����֥�Fd���G{��uR�a}�cbT�����o;�_!�V��! �:(DΠB&�"9kڄ�6���VwL�����v��2Ct�ޛ����q���O�+G{�fPv�{������5դ���YZ�ȼ릀n\�9��[�I1k��{=���9x�2��tߪͷՍ��f��.�i��Ƃy�����ĎaVJ3�˕]��"5S��>�
�^�9�I$3�[�mxx��q;����M�AT��W��;4�U��y*��F�p9��R+����֠�DA�)���lbb����:a�F˷�odKܚ���S�%���.{�'&{o�saN�����U�9�>���v�<��\b��=y�Y�y'={���o�2��aO�Ksm�׹��w��O^o1,O7�}:���؊m\��⨼��Ku���E߆;�Ǥ��&�T�E)���g������j�fΣж���̭Z\�QF����*v��^L�n<^����@�v>ɾ3�W�i��Z|�����c/;I�Q������j��&cs�WAD�Hf�oX��Nm��t����e��r�M�r�h���Wֽ(y0e�=W��w^<:@{�D��YW9�[�@��A��fVa�����o.[c&V0\M�9\���B�j�s�d�І)��[Z�W��#u=|���Q����M�u�������g]�}T��Q�=ԬQ�)�E��%��'��f����S���wz���H¢�+.��R��OOdX=�pM`�T�k�q&+^Po�6N���&-|�˓��B�"�����ƻ)z�.Ѯ�����A��ޚ���h�� �.7�}���alt!���'�r��<�z�.�Vڠ�f�c���1Us����;��s�C�+ $.5/l�1I���>�;��V�*n���;�|M?��t}lf�b�+��@܈j���m�.����ğxMд�/1���6�t��wNQ.G{�P�0������nU��Ө]0�s����������oh�<4D��ϙ���X5֣-�,��;���s���:M�7�����7��6��TG����2�y��om<��u4���UȠԤP�'\Sv���\=۲�+�"k�0�tCt�&���]n�,�W�W��2�+��ct�v�߾���uC�=�G �4v�;ɘ�}�FB����ؖ�����*�m۞����������<��2�eb���ܭ�Bnd�*��l����%ۓ���L���0�~�v�[��W.e��[b姐L��{u�s1`���bpdbl�����\��H�#�ye�G
�}���tXR!�r�e\�!mV����Z�rW�3+Ն�(�{��x|3������k�ql\#X���w�����uu�-��*}���h���4k[3�<σ��8x/}�U��!�����)Υ���_G3~��(ZPc�jv�|���g�K1J%/<�,���>�}V����V��z@��;�i�*������[��8�{��7n	S+w}"Ĵ�YI��ĺ�=���Fw7g��f�t�@�Zqǈ2�-!X��Ҝ��%�$�u+/DphYL/�(�����X��9�X�Y���ZzN��@��1��}j*b27��L���'A�V&b��L�x���El�����+b/*W����qp2g�|��"~6�q�2���kГ��#F��g��-�Q�G�O��
���r��C\�q��V�["=]�Ƽ��1�oDu��n������a^����@�m��G7�¥�9�������d���v@n���U2��=Y»����=�X�`����Gu���7[�-��#x7�C��^
�HR�D�,k{|U�Cc,T-{8L�:�j���u�=B96l%)�m����b���9�����W�<�����;9�5.�k:ϯ��0��AU�#mH>Ե^E�7��lX��ϳ�������g���;Fx[��,p��޺Ix ��k���j{}�˷�!o9�b���$���ߤ���J���Ȫ��HoA�v�[���,:i�(S���j�Sڿ%��V	,��O �K�]o®s'{��O��t=�+�W�b}�1�z�`�C���C��Zt�=w�r���f�B��Nn��V�K��mv�䶜Η�͛\�c#8��|�[z٭:uŏ,�[K4cv�U�ſ_|�PT�����s��O�ލ��e\u�p%I"���1��'8]��o�����ݻ�j𚒡��=dG��"�$�wOL���"ns�R�c���C�2{���ޱ�w}I��O#�m8��/o�fP���V(�C�nK��r�y��Y#��F�<w9Ac��:�>�K���\ �z�lN쏨o��nYa�����!gdǏ�F�z�uʞ��}M� ��~=W�,K�27Ƣ��u����6�V��m��(&��_;�v�,�$x�^pҾYT��k�R#9�_�)q�z�-�U���J��������O�CF�t�
�K��a�$)K�]vק3���֪9��uJF�X=��>1����b�ǝ�Z��G(z8F:4O.��'"s}Q�+sݓ8B��j�j\q�v��0oR�v˗\#���H:����
�z�5;1e=x�ik��i�gw��i_���No�r(l�U���2
��O;hmޱ�H�hf85,mY��p��H�^�0p��F�
���+Q(���d����ˑ��36N|�n-��BH���4�z�f�r�$w+s����0��⥭�q�������c�n!�D�:\�g-��%�e[ثcs�v�ә��� �UZ�đ�[R*bi��z���u|�ȡ��F˷�{�ܔ�D�j��&��d酲�f���
x���|�s����Vy������eM�z��QI���LIw�R�^A�犯�6��i���S��.oW��f�����<5�R�V��7,
}��ӓ���N:��}��E<�(�����ln�an껐3l_t��˪�+�Z���Q�^e��3}ɧ����#�Y�����z�J���.Q�4&��N�-4b�g(�5��7��/b����Sΰ���Ԭ� ]�0�=7<�+{4s�'�*hu�꺼|u��.@�u@r���+�w�)��H��'=U��l���ne���;_�����3r����T-ve���7�㬧�geԭ�	���z��B��3l>��~����mvPm!EĢ�� �f�E��&�t�������o�{Q�ӼK��a�ۄ�����4�.�1r�
������e+w�&e��>��Zeǒ,�J˳[��l�!%��5_��Q:�n"^Z��̮���˺���L�2	���܁�oqV��'[���斡�žRw��T��؝X�dZs��{t���䓓{��|��NR�v]���#�]�y��x6�}]׺R��{F�Y�.8�{9����+c$n�m:w�����VY�論v�4���k����rhg���U.E{�P��lR��pU���
C�n���Sے��p�xs�FĆ�eȞ�[T˩J�mE�hk��P���b^�n�	W�C9�j��#�L��LK�1�Oh]Q;�}O{S������MP�����e^	V���O�2�q�����wemM���W�a����[��8;憖x�^*���bpg���<�Y�";v�/m�|Q�4�PΔU�mګ85���{�D��X*�	��NC�	^�*<���ӳ�����B���+�wƆ<7A<;����-D�ϣ��'���S
K����wa\VN��MǺ�=�Ռ%�v&Vn�c� �d���(tݣ��WTb��z���Q�ń*f'�J����s�'%ֹ>�2�]���|�bV�or��>@�w����b�s�j������S�<��#���*(��wP�ƻ��R�Q�vz�z{���ck}eG���lh����>����T;�2�Ǭ��^�r({m��T���C�̇����ɘ*��Il�@*汅m-�v7y�X^q���,.O�#�Hi����k�6��g������ƸK�<�M�L47����u�V �6��n��ѳ�"4�S �"���_s�HdB�����UpM�T͛]f�dA�X���+ik�ΰ�>�հ��nC��i�[y6�!y��;&f�8[�aq� �����y\+Nv�
�S��}mZ�0���"�N�k��o3E��R�*ݔ�w>s�vΫ��A������X�tӔ����Z�e� A|B��ݢ��iJ^����F����t��\�j�P�3���xX�˭O��M�����6���;�z�o�����k��1'WyE�C���U4h�VR���ݜ�ݛ�ެ���e��s)>*gd�D��n(��˽�V�!����GT�[jJ�p�2� ����:0Y�}�����;��j�+zq����d����O;�if���z����	�������(d��
�V�$`�mTa8^+ک�4�)�W��4��V�kN@�o��p�Yy�Ua�P�V���]�ɭhA�2�	�kfB��Ê-�.U�,5���\q�ZUC=d`��n��Howm:[���2��8UX(�� �$�덣Wc��m��X}Zt��Qy�o�_k��.A)���/��D��~Z7�&�j��Hݺ����=>bwV�]�)[yf������ej+�{)�{c�W�u]����؊+�X+Ma"�A\��K�U�΋]�{�y�X0�]��p����ӱ�8v�'Jo˪�Z{2�}s �x�͙�	�i�Ss�<�~|`��R*h<�on�� ��xTT��G3*��`�8��+�T�D
$��5��\��6�m���ڈ�"@�4�)¤���'Z*�k^�υ�U��ᄞ�Y6��A�+�ܑq��-sh�l^��+���ӛ�]�bCS}�R'�KA��仙�uff��-c*�z�i��+N�KS���2'��Jh}}�|oma����{�Y)��ew]�7b�{�ڰ,Kxatn�m�9np��@�`�VpO^���j]=�����v�ӂ 2�U�׳ig_. �Y��qۃc=ڵP
�yNg�|��K��J�N�!ޡ)����7I����S֠��&�����嫻��ͺQq�z��	����w{i��.�`C�ځ��˳�n;-`b�1�g$�!�~�xwƯu��+�>���0�y��oT=�n��u_e6�,��A�}ō�E{���w_wį�Y�ju]:; ˎq;������Y��F�ݼxbM����j�,Qξfj4�[Ӻ�U�4��PD���#O��-t6q���F�u%���m����}��pn�R9�u&!�l�� �O��b *�`��(� �Wm�"�E�DAdU�����U+U��(������QB1��"�",R*�E�U��XQ+(�B,%J�b�AAE�EF)UEF"�k"�EPQb�T�`��&-��eTp�	�*�"��� ĩb0�G�c��B�����(�
[A��0�A��	Eb��X,"�VfdŪ
�,����0�U�(X�,E"�V",U�((�,R*�"*��,
�AAA�ʑ��DX�P�
�+cU�1�aX�F)F*2"#�kPX,iJ��c���UEjJ�EKec��g��j�����	�	�W��]]!m>�T�E7�ި�|����d�̽�tGh�5J��pM�Cel9�D00�d��,`]�L*q(�u�c�vZVr۝��4e��	�(>'Ta_[S%_tr�8��Aջpuk���A���8t��5�:-H��9����U���I�痃��/
9�eL����C�5�]1�m�T4���ڥ�ջ�!,V���eq(Y��y	s�4q���P*�r����UO �w���.���Ʉ<ڐ��K����{�ab���*��a �ޢz�z_*��Oev�{�R5n��8".Bw�s�!��?O]�1�Wb(����{��-P�=�-s}��K�#�an)���#�G�ԉqC^������@Hv�{�������r��ѵŁ	m��3����O�=��n�0#��ԼP���c;�.{S�bc6��9[ҴcR!<�N����o$�M_3��(�}���
����l;��Yc���cy�_KLw����q�t罏W ���}�	�R�Ѫ9^�k��xs�hK���,u�
� w��J���A�% Y�7Kz^Pݘ����H4�Cp����mc��c�=`�з�tŘ�ȩ�l�}���s��˲rV���x5ϙBu����S���)�+w�p�/4�>{c1+DA���5}X�����o!���"F��g��w^�9�]��SSˢh��)YΩ=���@ǥ�afj�X�9��p\�I�\���.V5��T�%�ؚ��tޛ�������t�����O�5�i]s�BuV��u��ta����s"�y^�w����{��qys�媍�J�v����b�㹠��B�hM�+��[�u�=݂����U'M<�ki��.v��k2�;;B�u��*�1ֆ���\�ZV��N!�u���g)����x���$��*g��L��ƛ�o��t��v.�y���T8��iNJO0w<���c���1>����(�F�c}yt�Ѽ�.�xI��h��]D�G}�����׸fYE�g�Q��{,�L�朜�*v�W�db{��[۽�ͧY���i��u�F�^��|ѷ.F�.���}��	׎Y�VW�3��H"3�1�Gq�V!NL)^D�gw������J�Y ���(z��ތIIK���2���+5.)UA�*��D,��S��Nt�V�{Z���n�V�NA�"V��5h�v�x�b������f27����r��d5r �6ۣ�]�3��>쩻�~ђ��$��5Bd�{$Z�mg�s����淡��Ц����n]CJ+y=d��"��%B:��*�X!r=c�-��m��nxK�%��'c�������x2��S3��`x�ldv}7Ea�;=��=c��V^�����#\9\�jgkq���[�9��T���먫J�>r����WJ�ڻ�׻�����:ڄ<B7��pÙ�h�K���=נI��f��8>+>;�r�������9�`�݃�lHn�Sr��0�a�r�W9C�^�q����6��˼�mL.����Vߞ����_�2Pv��{��e	¹iƻid=N�(��^�6Q��Br�����*56�;Ҡ�v��:k:�yq����
=d�fNν�U��%�p�Z�u ��eu����kt�e��0�k���r�f��6�D���V�z6���3~�����'M��յUV%0p�B}�Ć�u��6��굅T:Xl�Zꈇ��ʼĎ�ɬw�q�66������V���=˓����ǽ�ΑI�)\�T�"&�H�8��/���1�}e󱶒=}w=�yM���P��\�3U��}v��\��Տ�߲�d�;�Y]�O�7妨6����r�մ^m����#z��{��C �����ܔ�:!��Ǯ��N��xk����'Z��[u��;sAd�3��LXTysyjr;ciOn���=���4�n�'О��wG�S���ub9I��8����L��o�<[���#2�oj��l�p��9jk�H���tDZyYTr��Q���]���tw0m�j�l��J�k�=��Ӱ�Ć�	[��ڭ�����R�nd0����۝��8���
Ƹ��2���Us�uZ���E��iB'vI��7���� bϦ3�������ho���Y�u��YT1omij9�1�o��F��x*�Ҏp3 ��	�\Ե�U�&P����Yctl ��Bh��wzn'�{�}t��,�&y0<y�1����q�����rk�P����^//.U��� �'
`�',eK�]��kLD��~�t�'~�&{��u�����Zpe<�|��pfT>��W�Nr[!�0�o�M����Κ���͘c����9{ۻ�{ۛ�jvR�qMc�5�������
T�z�7�A�%�_����yV�B��;�H�l�x��۳��'w�u[��5�xA/�*ּǐ��}�>��n���(�����T��Mjƕ�ܮ����-�TU��]��W�*MK�5o>�U�(v����J��V��w�~�[F yiV:�=��/��z��,�ݛ}%^������x�$~ޥ��z���CAW�t��Pp�w$����x���k{�З���4��׼��Vu:lu��P�%��ss2˂�`�����{���Czj�<�eh}��r;�Q��d�}42����@����G
d�,SF�p=�Y���D|�>�-5y�^�o&��DQ��e����K6I��÷�ws܈�J>	v���f��2��v��(���Tu�.�Y�j��jv�r,�-C%�U>B:�u����K}��s:�ݦ��{���{{�v�
����j�DT_Qz$F*5��r�U {������!b�k܋�������ʑA�j�dt�ȓc�ͧ��\�}����S�3W{���բn�6lKo+���B?k�,�o�J��l޿u ��>tg�ns����DA{s"�lC�b'���0��\��@�{;�sȤ�ԭe�KN�{oV^|ܩ�)��J5�N��eY������a��]'���߷����\aO�Kscx�Y��vS�*���t�����L��SJ��Su�OM��ϵ��(������5{�Px[��xW�ܯ)��5܉xR�o�c�ю4՜��9�B��wxs���n���������-|�s�&`�Z(���)��#��^V	�1��r����ȅ��,���(0v�Cn){�f��I롷D)�T�����ah!ln�B��]6����-Э]��6�����h1�����<�;j̐U��O�J������c">ߤoDYd�g��J����b!�g�N{|��	�UPg������/�E�\G�Kg�ǀ�p��Y�1gf�oϻÞˮ���!��>{���ӏ���M.������RڳܶV�N�w�r|
Z���Mɸ4@ۀ*�[��G8c8�NЩ/��.������o�r[�¢��{�f[�;���n[��51�"����:��m	Α�u��#�˞̌���F;Znvv1��k�*�ʁ}�1Q���Y	���m��T޻�gN�j�27�[v�T�9��#�z`���y��U�U�ߓW~^�=D�^pɺX�ͣ�Û��v'؛ؑ���ˌ�����d����U,49h�,h����="9���6$7bG;.(���0m.O~m�����������������3|Ň�/���]g
�'v�,Kr�5@,�$�r[C\	'SN"՜�W,�g���L���mq���q�V(Ȭ��KI8v�I�n��w��kv�^	z�����=KUSBw8L�N�g�:�+m�9��Tޗ0sVgu���_�CRFN@�Jݕ7�֒�Ʋ��0 �;�ח.�{����:�>�Πj��q�� .�m+ز��T�=4_L=�rr�g��+)8�#m�Ɗ�ƅp�� NJ�՗G��|�����Z�Y���J�
���(y/+�=n0�GޯGp����k*>]KS�t=3g�3�6b{�h�N��9�Sa��~�����MQAdT�#���y���;;ְ������ =�N�����ُ���w^n3����IPҧ��r��Z�����Κ���ՃϬ�����F�1���n��u�ҔN?W5<��_Aۡҳ��!��ҼYk;h��
�R
�uנĉ{�G����tښ�"`�H�v��p�;��v�ޜ��ăC��"�
�t{�	D�'6�1E%�B�]���9�Qn��v���	W�9P/���8;U�՘(�ۆ����w���+��]�(�W��9��C#����{B�Ĵ��������5���M����3a�n�"Cn��k�6k�5[`��%̣�_<@=�+�]�e)Q��[Fq��WL�5i�
�%ԧ�D秔 �s�˷�����
h\NkTs��G�k5�9�F�)`��;�+t���I��E6_Q�Wgl��U��g+�V6��+//^8Ν��
��+�ǁ.Te�]�̖c����u�ݸOy��~���ro����d:�別B���4s�ێ���Q��{���rq�9:���RF����=�mu��P�v���qp��oL��y`Syx�kݓ�sM�]s�T]���;0��dh�$V�F׫�>�n���>��8��\�k'w8�i�83���/�l�釴 �W�����sX��{�Ւ:yvss;�R�ٸ4�}�B'?R�d��\�>O�i�w��/G��������罖O.����a9�@'�B�>�W|a�8�٬ɝ�+�S5�����[n�r�vu@�҄�Ǐ ���8��7�q����tsF�a��wӵ���jdM��b��r9[5��{�$���K%J2��n�մp�[����{7�Dܪ������n��.E>Unm���rr�+=�eN���
�߈��F��xo;�obo�����p
|�!F�Zbp�p�{I�����-����$vш�uq�թ5�Ə,]�������7���}�MU���������%��vL��uvܴ�M�ZxU[F RQ�+=U�q��}�f�,I�V�X��Ḓ$��챳�ګO1���[�vzy�D6"��W��r��74��}�C���>=M-�/�C�������.��ٯ��
 ՐG[�V��gfؘ��@5�=����+v����^]N�+[|y��v�J�^�&���'#wU�soc�nAX�Ct��Nx�R3m��w��������9��0��\�[���z[���S��6qT�a�f�n�)�4�=��o��W_'
��9�'��l�]�����Ib�.B�[܄<��DP�oz�ߟ}y���Z��y�!s|H՗6X��y�M)a��á�r���	�w����L�:*���t����%��Uݓ������ ��w��Ջ�RY�pJ��T"
b�)��:��u�՘W�?��Oj���²�#�r����\&���0 ����*��CL.�K���ő�O;��F;��&����
ds6�?O�����_^�a�ے���1^u{̵}�!�:��w4,���c5���Qd����ц���[lX���،��S����������9�6]���ux�M��܇�cj�s�
[���+0ꃜ��f�i�,m��rUR�-}C��Uf��	�kr](�எ]�2'N���y)�zv�KF��\����0�YEd�f(y���F�]�i(��F�ؘ������i\)�]��6�*����*A�t�s)ӛ,���7��#6m�ˮy��\�"�n@����.V4���^�����Nm.�D.�ݮ�F+�K�/`��x��{1ʺ��y̗��i�KS�c��nsi�W[%��NJǋ �8T��|i�ϙ{W|����� �}h��ۥh��veݦ�qǛg�Eä��OQtޖ�R5Yv{�p���x8'X��Y������բ�T�r̼��Z�Oɶ:WJ�K��ӝ�0�{K��g4��u�
޺Ee����fe���C�k%�7:�p��ls�h���+�	X�g.��<2�XܵW�02���z��8��XW4Ĳ���3Z��y�r�c��4:��,�U�qQ'���Ý�,�9:��)V���VE"?��5��?I���\9�;A�>���a�G�2��9ދV�=baD�
�8ͅ4��t+�`�rßN�0��r�a/t�$�}486&�9�L���G��-	�S��]��V*��d��Y���X&�A�XHBW�P�I�����8vhn���[׬������ڪj�(�rѫ`���*j:7bG�G�G��n���5MB����*��E]��h��v�a9Ib�Ʀ�y6�s���f�6÷���A��$1��W�gϜ�iA&l�	ض���q����rψD�'uX�ʹt�G{��	�R��M#�[[�����B �淏s����Aq�z�h������K;]1���w=ϺY�a4Y�k����u+:��)ڋ�!2��н�vש�6x�\4�W%xdk�7ٞ���nSK�t��piش}�6�W��V�:�Y���$h�u�4᝶,�hXc?)�89ӎ�vLsn��2nѮᵎU��\��������~��?�TQ�U��c-�ň��Ո� ����V�QJ�XT*�A@Y"IX�AH��$��QH�Z�U�`�PVJ�E�PR�X(��Y�(��R,P-hIP� �(�DDR�XT����ȢȢ���������,QUH�(*�EJ�1H�T��	Z�X�QH��F(��TX��X��QH�"*E�(ʔ)R�mVV-����P�����(�VJőA`
,*����E`)����Qd
��+KA`���d�XڡZ�L/0��&��sl�6f�bzɲZ�����w��e��rXox����� "2�Tm����{���h�g@sM�ՑE7���+J�v�[��ė��/�tܙ�
�8��r��]�M��e����F�킦Όw�]3&�֜n���u�n}jQ}֠cphky���h�����D���,{2�t17xDo����<��Օ��uz�I���d��[�Q���&`�b�#876���ü��,S�>ǪQ�����z���P�*�n�:��7%��Ar��u#y�F!pL�i�Et�쁑<�7m��okp��ç��H'���ܢ6_�����{Jq'w�2���w|�;
t��@�t-�=�xGt�&��C,Êch���*�	\�m.���ٖUD��h�u���{*�[J�=]ٽљ����h<��G="�DWX��t�]u�y��]D<4�w-isG�x��k�o��r�J��*�1 F���N�=�t�Ƴ@�b7YO��.RZ�$��$7�=4���h�C�g����ˣ�n98_aj��ж��L��5�C(��3�1Z���aov[�t��8j�e��M�2���e.U z8�;n�=#��(�uc�N�rkP��Fl�#4A=�{���ØӣR��e,��~m�u����J�p��$�b�7��5žɝoL�7��	q���CrR�xrp�vw9��ċ�L>jl��[1~��,�ލwʻ�����L7(𐝉���ZE�R����>S�Cbi���ܢUeXv���8�k�+�^��sl\��=Ƿ9̾�g����<�1:6��'3/ҭ��pdz�ٕ�y[�y1\R�;5,�͉ڌ�c��� ���!����Y��I�y	4{��v�d��u�m�$Q�4�W�t���hnt1�6��u
s�C�ޞ̹w
g^���ӗ�7ۺ
~�sک�+o�)�̰X��I��sç���7�_�5P�1������hOsE/|!�-�f��T��NLOt0gLd���O�����r����+�X3s���lhM_]�mS�~��:<����Ti���ZY�W��6ZW�+��uPLR/,@��Կvu�==j_k���k��<k>���R��阣�+��H��gs��{�k��䀴�>c�3g����iZI�W�Yj�R.��j��h�M����VG:��Q{(�P��ޣ�Į��qk�Kd��^�o�,ȭ���7e&�.�H*��"A/�;���uMlI���.al��W����;s/Ú� �n�vCS���
;E�@�2�b�r�Oq�x�9�Xo.���wwj���nR�v��@J�g*�xh=`�u�x�%s��X���+#dft���V�K�29�\�5Ӕ�)p�"�D>\;%�սsx	S�6ÏE����9�ݘ��rq��N�Xw�����S���QXt⼺O+���eװ���T'�UNc�^���w�V��eH��>�:�q�N�+ر��s�Wֵ@�n�OW=�k+%i��;0k��H�n4_���#����EV���0�>�H�>ի,>��7}d�_�J�/�����������c*��Y���:�]�I�y���5<H��X�ݶvM�S��V��,�ԓǔwgW�ʇ�5p�v���s�9������RA�G1�D7���T�Mw&�)��p{PZXMէ���;�N��p,�|c:��0CU��29Ev�&m[U;bA8c��F�t��ϣ�ʣ:��W�66}���qV�/S�)�`�Ϡ�u�p��W�E��;4�[���[=�NK��x1c�@��>�n�w�8��Ѵ�����O�>c��t���X���&���ک�o����m��gvn��`�9�,�t�O��tN�L���A�+bZ��ULܪq׭����tgZ�{pc�f�t��n�:ޮ���ux��ʣK�"����+�7*�IUc�%��K��\��<�)��O
���8wvڎ�ц�dxڵ2�Y��GUV?#��e�+����V��u����~���a=ҷ���IA�~��T櫔�����wSw��d�I�u��Ռ���h�[������p�g�ê�MWe	��n�kZ��m,�I�ƒ�n��+��Tֺ�$oax&5Q�C]�1=�Zq� P�C��t�����]�H{��ˮ%�2�+���b�-�Mn��T�F�wܮn:3gSW�e0t9�7:�^.���u����N�wws�H���c�9��ә@@s�3}8/��xL/���k7�*�u��w�ˤ��xS�[g2��vZ.�j���?����=�o��Fl�S˵{E\����Ԛ�Ȃ�冓<ؖ�R�r(t��j^�ʙ�:E�����̰y��>���7��M��V��_V5L���N�X����t��(K�{9ŭN�l�9c-�ī�}����1c]A0tZͫ�uy��bE�P؛b�2j�Z�Őg��T8-K.ӝݘS;�4�؂��u]tn�8�奏Q��L��/�&np�O,N�=�v�����"�+��&�+Tn��Zxn��7(1�t���]S�)�"k�i4���\"����+�~�E��|<0�S�y������Pv/wreH���KQUO��r�ک�XnV!��Q�#�s��.�7~ ߶E��"b��a	�oM���E�	��Y�s8�9�I:*��{
}�h��7�a�wA�Fe�$u����8�oי ț���x?��}��t���9�M�ǁ)
n���-�xZ���N�9<�#����-ɸ�:�a�O�V��v7���֙P`�N>P�  %�e�����$6�:W��;0P�t��ՄG�[� gb��"�sz�գ3<z��wφґ�;�Y�7�K�_*
�����3��1";�P;�^&z+��׭.��z�]�u���<oqs�"6/h2k�ek����T�U	�"@��w�K[µn��ܲ�]��nNL7���O؆�~{�����C!-/��07���xk����`�&��������m�[���eO8h\jW;�RɍYƎnos[�ZhJ�~�"�)�׎OTrp�	��`�ܰ#���0G���:ym�� �\�y�(�:�7�-
	��݇�rIzko����ʄ��~
a��:��&��MN,sj�L)\O&
��k�[z�yu"�w�5��\2�m��L��jMym���m9s2�[�Őg�uR�&��w/&
�Ѧ�$�{_A����v$��ʹ��x��q�.��^������|��#�j�P�P]l�}R��N��Q�j��}�I�	@���� 9j�tǥ*�(a]����}[��H���O&�ҩ�V7�c�Vv�f�G��M9(o*v�n.詸��#��n�ɇ;T����$?��9��l�^o.��ۯ:l�ׁ
jWS	���o���=QQ�c���gJ׃]��yO�7+ŋ}P�-E���i�z�w��},K���{��K��5[)4����g���8x�S�w{�sV�J�"���ez6x��u+��sL(��K��9����T�Y�k[>O}Б���a���3
�!��z��URV%"����}3{�'�/������>s����Uh¢�Tu�zg��]|�=8C�bnA���Cj���^��)��zWi,����:(�θ�P�#�ż��e4�[��Y���b����;��;��nrS�lb����m��8%�u�LP쉈�l��er�����6�����=�T��l�գ�^ö�{�E��ǔ�V�����f��ڱ.�O�P�.�ĸW�F"'@1 2ɓع��͖w��O���N�39dS)$�7�]>[lR�L���.�n�Z��=�ч��Z�Aj�c2���Xw]t�M,�<�wWv�P`-��V�i!^�o+cfM��U�MԫD!j��v��.�"+ܦ��:t
^3y�j���w�l���T�
�2�H���Yۙ��������q���~�s���]{Y*U��9w=���ڲh�sλ� �ⶱÕ���b:&c���IU�N�6+�VȊn�s`����
j��!	��t�����+q�Z�ng�-88���hB��v���*�&}(ʭl��T<���a�mAl�
�]*�DwC�rlg}^�@JL�1!5Q���Ez����4E�렱��߻&���z�D��;�����wֲ�չ�}`�i�o�uη�ax���y�};�P����L��dí������ؑt�!t�(�g���;钤P�T�Ny�Q���5Ι�1/����pa�SCqq�T��{�:�+�5����*�-`�e5�*�xj������,��X<�3s�:�]3�yR��;�]�7\��T;1R8ݚ��y�Q�t���璏�O��lsiXGu:[.���SM��(����+�Kܷ�!j�N��Q/P�-#���m�)��Ek۴��t3^-���1fN�4%н�������k�a%�##�Q�D.Ƣ��ۺ�2.���ͧU6�7v��x�ZX��c��P���:���V_��
s��<9AÉA��s<���ز�mf��\��.u�w9��Ѐ�\��6%��X�}W�x�uF��.x��u��$.�}���������A=��S����j��\����#��ٸ�����7M���
���O5���C��؎� �9i�����3�K=,D��#_o��k����@��=����}e�p,�gt����%���L�N��[y�e��1niSԠ_���W��t�Bvǉ�gh[��q3-���2�'�K[��r=A�rEW�Z������E T��O.�c.Bv*�H@�̔D�-��N=�\�M�k�ء%G���]��1�߲��P�Yn+т0[��ZѶ��!6�d��#jn����A�9 *�zz!+�~dJ��ݮ�yϗ��=�b��]��y�ۗO`��w��f���^U��T�K�;���e�^ a���Up1NŪ����F�[�on����w�`�K�X�U�����B��OƗ�Ρ9�SQ�b!������t���P�)�.�˝���u5;���'&�%��y��\��*�>,ͱw=w�8��+��&��]�&;El\_�K虨���]�u@�46׉OD5�o�`�u��Y՟:�Ί�R]<�{�>/M($:(C�ܤ�����g.F��{~譞�����1��A���Mخ㻝v���A�Ir��`�W5DV<;¹-�茖�y	�Z��I\�a�TV����d�vZ��4����s�����X�)$ ���g?f}�S�r=�DR�_3�YΖ�-Z�?TZ
H���B��$�z#o���x�5
��"��!��69U8��k��m�Lq!w�gu����V���F�l{3M��v�<��>��EgY�~�~J
�p�/V�o�Pb��Ȱ���0@=��cn�;��t;D�hj*���aI�qZRR╺��i�:fл�F�Nβ���7�I�t��j�hyRb�=eE���l��W��8�3�6;R���[qYFq�]�R���ڭ��#/{�:���8�:�@^[�U�À�4]7��-	R��_Z�#�M푪���u\�.7Ǵҋ���D(��I@p��mWv=�����Fx�q�Ŵ (ҭ�c\�I���*,�_��8!�ůy�-s��.���Q��1�|-tmM�͵9�����P��3f���S�B�+9:]��i��{��+�<QS*����>;o�o�@.��@�����P�N':!���q:@��T<;��}��e�q<Sq�Y������2����(��pg��^���֝b����̛�`QR�TZ5~��G�c����(\��|�:��K�;��+ o
�{��<%�9�]Y��n� c]j�"���t�&�V#���fª	M�4�pG�`�ܮ�A��\�/jw_7R`U�KWlۮf�|��I���o�*�m7V�y�z��%$k��h87L*����s�R�i�*�
�7�'�]Z�m����2��Ec�x6M� ���g'}�`=�w�i��2Q�Ƭd����6�5٩��}e��gі��R��P�UY�jT�4��v��ڭ�12��6`�m��[���Y�b鴲��ݬ>�a�J���/:b���ӹ٫����K�	��b��%bp�N�
cޞ�C���Q�/D4��ڏruA��]�J�N/{.`��܌5�8|+�E��\mڥ�v0�14���5{�^��<U��LCC��MS���[���A0Dī/`K>��D9�����
VJȇ`���ȴ�f�rqH�x쥸�Iͽ�¼cm��,lմ����5ښV�G�8|����358i�%ި���
Y��S�3�ӕ`�v���_Psf�X+�u�Ӽ�Y�7�EڏF^g`ld��WIl��V,�y0�h�8����8î�+�� ���;�*Ww�� ܫB@Ǐ����i�:���u�U�u���¦p���[�M.��$�y�e���\j��.Εo���[o!/1�	ٲkZ�탉��U�M(f�t�6��Z�������ȫ8��5٘8�:�X�9[zo�����u�+�I{�bOyf&\2�kCb�-Hmΰƈ`<=	�
L��9�R�-UI�b���P�ѥGxkw4�H__R�ڨ3ʻĄCr��V�S@_|r����hv���d�s	`703�v��w#��N�r��62d9��N�z)����F��xh��:����%7s�:�[{��m^ۻ�t����8>oP��/T췁�i��Z��R;U��)fV�M��K;�;.L`�FY���9�F9L
<U�lU��v7�.LX�dna����=�z��T�{e����Ҷ\���|���������,K�ģ��\����4�N��4��y�\/�M�fcWV�7ǆ����2��ڱW��e�!�dov�t-K<w�
���$�D��zpX��8U��5T�V���A3}ԓma�N�>�V��MT�궕�36r�wwX�:��D��m�5�s-��ݻmb-벐i�9����QUɹGB!���=y��;��!|{���)uс�m+�̽��9���_IV��̭��DWי.���˔ �ٔ��n��x�i+R���<��x
ܾ�ѵ��{�#�b�(�Q�v_b�a�ۢ&1}T�Uk_v���χ_&���]��{��Z���\O����K=(A��,��{�\x�k:p�u�h\{��`�:���4ɛ�S��3[�!�V���/Ou5�n�3�8�4w79�pZ��'z�R�d-�J���{C3V���y�o�Q��ժ=n֌Ϋ��C^M�h ӓ z#�WwVe!b
�X�*YE-T)�A�T���ł��Z�X(�,X6�PX��ŋ`�eUb���+d+++RT%*TZ¢ň��V�eDU�#
ʄPR�DYjT�"2
��
� �����
��(
E(�PUR,�DX,
��+%-��J��YQ`�)e�R
*�E"�#l�ʬh��-E
��j
�R��)+�PhѶ���-��B���H�"�V�E�
�,b����E*%@Pm�ZJ[!Q���eeD�+h�P�am(�QjJ�#(��YD�H6��
���-�Z�E���+(��*��@Q��$�r��9YmVsm/�JU|z�u��W׊��5Z���U�\���i̓m��T��^�\��G��ي��P`�f6�"�S���l��ts��W3:����YK�����׸5KS�ώ)BE��ޕZ�%5�Z��gc�+)z;g��Fl��4T`�&�O=6Z�1���3�syj��7P��>�lVDG;.��UE��z���ȫ#)MaXL���0��3o:��0�����q�E
���h������Ӌ��{CZ\^~GV�������2�V��o]7��u��2���a�!X�M���d�N��\PY;��#��^�M�f�o�PV=O�݋Zq��v�@�5�Dt�`�nhgMB���tߧ����pꙌ.P�ݽ�;�{���� �D����Þ X����5WY�C�Wf�X�$�̭(�p�v�=V��y`��N_�uj�m��)�����ƅ+;���{_x�{d��7�9o�m��LM���{s�Be�Q�����$+���W�:��]�B�S�xo]cC����]_/qe=ы �KY#+UH���;nd�ޕ@*��-��~{���j��]l4��*X���K»a����Jʒ'�amQ�̦rǪJ�&���{Kucѹ֑�Gp�N��Ҏ��)u�Ь�;�9w+�c3�
JUwײU���S(y�EH�������\����n��z�	�^2Т�����>�ݱ�oQQ.�Ss
 ��j���)mxP�o�K��{L��u�(�ǆ�9Vz� o�	�y�q���om�\���Ѵz!���o�7��9�Oq�S���8hk}�h��u��ܘWk��3w��,qn�M��b��S� +Q�B��|n��b
n}���Ɍ���
�ъ�'b��߻7o��/�v
U���Z:cd ��8e���-v�=١k��`�a��E̙�� �8e)�N����m�Ц1��w"0�P$�3<'X�����	(	��tۛ��ׯ꣓���e8�.�1�� R�wQ�E�/mف�ڂٔ8W�ӗ�ޘ��2W���٢��>��Uo㢐Y���qV χ�$/�ʼ�nz6�ʬPpo۳D���ڜo�}��kA����gsK�y>�1#B��{��j�u��?D��U>�`_P|q�9�����'u
��ڼ9�s��
�Q����q�v:d���˜dLlP�p�2C���^�ng=��2DË�FN&{���M����vV�W&>��|'%��W�U�Jb����+*(.Ӗ�!I5���cj�WV�㬱z怖5��V�3����+��1�X!������a�����ћ�+�z����n�t�ܦ,�A���s�L���ݵZp�m(L47\�!�+/���0�Q�ی���o6�����x���=��fM@ǽ�Fa> U�;1RuN7f��1|@���뾬s.ĲK�\s">���1�}��/��m<�_E��[JE�s�ik�aB�����C
����ҳX�P�oBaր��p�ySˮ邰J�]�s�	/
2�:��&��s��Y��Y�>[���:�^K�c��q�{��=R&zG2���n7�0-��*�tp�����|�>a��%�mܿn쿻r��BJ���-ԭ�i3'.x��#��c&�mҼமSU��M]�~=�y�cA6�0���.q�*�?��M�7��z�ǎ��پx�|#��Ϫ\�!b�(Z�n
=Ǿ>^�Cutb�@ZxV|�U���\.�7�Of���{���Z�K��3tTy2YD�S~<�0�|�F�;تٮ�@��g���Ո!�--!"؝��^����Nncy���(sW���q�@�L��3�����<"���W��=;$dK	b�FL���,����o.b���ы3Zꇟ����9W	{�	F+���;2k��|K Cq�N���'�]��{���q��վ�s�n���	��j�QѯcֽҘ>�C=YV�J��y��\!��c7���|���j�;����2�¢]|go.��xkh� �ǷF�X��nøX�v�Hݴ=4�%C�n[TU�����-������GT��M��X�� �tC��"#l�1
[&1t�����Z�͡�b�?A�2��o`_����7�vX�q�ઌ	�BY!9�j�y�Q5P�_[���OFҨ!W�j���O��,�mu�
�0v�{Kg��"��z���U�Gt>����4�L,N��Q��Ȩѽ/BL1Z,�2W�4�������x�2`y#i����X�^N�x��E���ؕ[�GNJ^`u>>��v�ݐ�p����z�OMU)� �TDO���l7T�5��4-��
�1���Xbb��r�u��k��C�fNjͭK�]��xF#p9��P�P�׊��� o\������\s�����g-���'մ<�l>��@Y���0���+T��R8W�1Z�vS~g:���}��2`�J��W<MqQw3��>��^R1Rg#<#n,Q����q�g�t�q�o���d;����Q�J�#�O+bL����#c*T(�54������Y����o;2�sV
h�=�^v1s�ݥO���&�����?�Uս���)3^ۣx�s$䮶�����r�am�l7��m�:u5�LT�s��ƭ{f���fK<)�	�Nt��?����fݒzV2�F��t�2��@XhcU.V6����Y<����Y�8�Q���\a�4��H�*!o�u��8؋RK�h�k;���}�aZ� z��t�No-u�.�R�>�����'�b�KT�{4<��m4�ۗF�q�)���+�n0��9���ZnGN�s!�T��Yft��Z�a^�N�h���A7my���'#�qգY�2���T:���	��zT3Ӂ9���3�x-���>}���1Ȉ�a�ML=�@Xn���
���K�;ED#���y��/+;#v)`:�1R�k���!�s��h&`j�^ؘ����e���h}�2^z)E�/��3įxY`�~�ڈ���(s���TN�tZ�_����*]xb��9�������F:�ݦM"|�$p��@>}���}��Ff����g�k��me��h�{+7srP��U{
:.0��D�C�A�
s~�Ǒ��ʘ��l0%C&���B׺`��݋m��u5���c���Pf�9^�8xnz:�)z�AսO���\{�~�5lX�g:ԍ*��d�՞е������͇ι�q\5�X�}=W;g-�N�K�:��� �1(�^@; �@|s�6�jCw�Ȣy}Q�����8�g+��rR̓�V͊j�`!���m1[ً u+;w!�l
4�SXOhU(,é�*�%R��#(^k�2�O�c���U�,M�ldN<�����-u֬�B׽��Z����c&+}�w����;\����1'/Vބ��Z8��m�f������Y�
�?z� �]v_#n����ʀ�vT�bd���a��X���P��L�3�b9)061�D�&hevk�om#Vb���p�){��f�\���<�9��V��5����ǞE{��S�~�n���������آ~84�|p.���<yUvQ�5I좶.�m��+Ȝ{���6I-{�4cj�R&���N��]�P��F��0��҈�ލ�Ft��97U�w��<@a���9�la�IN[����=�b���:5>ף7dLHp���e��ʕBQ'0rK��%$��id٦qRn���E*l��Hw&8��rbw�n�O�7�S�j|�J�
U��GD� ��% �xGi��B��t����Dr��a���GeR�z��a�N�.�'��X���S�t�sG$�L
�Ybb�L����3T�OcR�d\֑�8�T����r��	\�㲇��9��-{W��9��ɴ��C�U5Eu���}c��Emb}�m_C��(C�Y=�)�[ŗ�4@��⋱VI�[[��2�y�̽%ȭ����z�kau�*�xR
�|��]rx t=P���*�4�=q��(8nf��{��^��չxg+P�]9Ƭl��bF�TPU�K5����>��>�`쬅at�����Ѽ']霫�,�=���I��m�c�2T�����Ș����{փ�97�u���Z[�z��
T��F��J����P<3���W�d:.�B�5��S���B|�+]rs�A��{g���Ō���K�݊���[u<ا���+�������u����O��h�j��C��$�"��^�ߵ���#�t�u�R��'$!ͽ�p슶�^g�<m9AUYBî�`=�\�d��/��-;��J��#$uJ=k�B�#vN��8aBo�Y8'[�s����x��M�����0�l���ݧ*D�	����T��mT�Z�(�%�BNA�	A�I`���n����.�R���7M����]A'*�Z���f�:2�����ۢ%��5��J[U�¤��(��9P���| Y˴�м���n��б�@͡aM��K���wM�Qw�u��桄^�����S�\�t]�N�p���w7B����=�/�r�e��8"<o���M8��V�t��pl4)ٗ��1�ܱa�}Wg�� \̱��Ϟ���F�'�w�r�vc�鼎R�1�\ܐ���<�'��� ��9��;��~ճh|�R�#��h�Ѐ����b��{T��鍚���*+#Q)�Bw��Q��n��P	˒A���ɎW�͈P�B����#�"�ؙt�_^d�;{5cjf��bv�
�&vXN�m �IJ'��|��O��7��z��ۍ�3E]��-&�V�i�[�BE�#�1�����<kǥ2�"�!�u0�fY=�1��s*�V��[���.{x�S13��m�M{A�φ�@S�막B.NB�Q��d��-�&ot�Cgm�j�{���/H�k����6�_�U�ZW�.6�Q���%���s\���L�ő�^��(�iBr;�7HQ4KA�riK9�*.U�a�����@6�vX>'��\��UکiO��>�Vu�Bz(� �ah��#��Ð�0��0@�^�Hv���v��b��x>LB~�%�a]�.ĭ�#�"��80|�^���=�=��;���jJI�EM�}t���8�qG9�yL���jV��sʘ����^�l��l�H�--��rή��:ȣx�e9A�O���E��V!O+��yw7xVj���$�#f����sl}*t�U�:m��=ԝ���\W���Am�d��n*;�W]S)AE�N�f�X!`Y��N���V��0N52Ԝ#��5�bRv�}�S:l���J�����YCc��G�U��o�ச����7be���r6��K{7�t���V,C�������Hh�P׻���:7��C����*�MQudfCg�n�e�N��,��H:]�RM'F�)�5%�kK����=��ޞ�b���ߗ���]��6��#0�d�.^R�cO3��g�Ҥ��q�BפȨ���s��L�P�gr�H��
�����}*2@uI�{(H����Ǻ�E��U1Ob�P�]�ݭhۿV��.����
Sm�ynY�f�Q`��F�V��Q~�r9}W��w4耢Ԧ�7w�=�����T���;��d=4��%br�Ob� Fan�e�]{�����O�\�G=���1_�VD��eH�;�bg	X�ž�1��Έ�C��DF�	��������é�1�"!q�_\���&���E�n�V^{3ʪj��Z�w�1K�d, ��$�l��6"�������4��tD���0*]�Q��Td�y�N��j���_N�~�6V�uYcӵ�Oˑt�6*'y�y����Ee�D�Sm9�7(�K)���Qoc;0�[�=q�`�Ns�Ot��^!��B3��废w\VF�	e�8�a-�V�;��X�M��˙VOM���X���:���f�۝�噢�fu��_{����������aN�������{r��L��=I�k�[���L����l�{,��t;iV�2�.���{�����2��8@��8��͡�xUB␷����(U*u=��q�X{��A�D�u�XQ��rz%�id�zV�YwI��㜯��X�O��w]�����F�91�5
k�/i4;K�e��o#�m4���':�'զ�T�vz�/�8�6�g��K��=�={d�|e���7�,9Oq0�z���0xX��>^Wf|y���c�i{Lw���>� �{ϲ�.ϓG=1ϼ��3�r�3�%���q�"(�Qp�p�^A�!X�!Bu�m�Q�Sk�7��-����խ�<���4ؔ�h���p��P�S��=>\��wH�uF�v��(I��Z�f�B�K}9�ۺ
ҡQ^������Ļ��OeJ6=�G�y�X&��f�Ģ#_�h	,i�� �.�B]<-�@�S�oئ =6�N	۰�y靼����n*�ȔR�V�Rݞ�!�9���:T���Z������R�.��1���t��yf��,��,V}[�����v,pfP7y�7SlpO~Y��(���oZz(-Ij��w�vt����4Iz
C�Xs&�)*Z��4jRTq���ι���.�q鷚��;����9��_
UX�ʪ1&y�s8���O�p�ڽ��xz]E�vS�A�����UpZ�ǝ}�al� 9�/3e�}�u��C��zAk�ž�)R��#���[yN�֦�p�p���zJ��`�2`��L8�'1��wY�'�������ݷPs��GCM�)�E��î���.k�,��p]%�7�C� b���z�S[�M�˛E7��D�)��v�쫐`�.�Z����j_`e:��"�>R��_���/�s�m&�0<t��@S/8i�'�ל(I�1����Ɋ����y�O��9������z�%:���_�����}ܡ����;k�����z����1n�ӺqR	Xa��x��b؁ûSV�P����!����%f�o�!XUiQZ7��Qڮv���0b����κLynV��t:xZ����2q}yn��yA׆����E���\���Tb��u�sD�triZA�q[���#k�9}F�i���FӠ��7+,/��2��ֱ}׸��]��Yݝ���[;|�ۇ�I�Z���/��)hҹ=�^��vo ����O7���e;�h��SM��e��%��F>��da?��۝�}Ƭ.6�n�r���M��������@�����e���\N����~B&�����g7x���N�>�3A")�-�C+w���7I����lh�'&�?��1D�?�@��\�:�G�hwp�:�&�$f����|t�|�����U���1Y�WY�e�*(b%�r��S�F�@��N�πx��T�c8>|d��i"!--����u��I��'�=_�B������ܸ�A���T"�k�-����\���E	wl�e�)!k�ੈj��;Pe�l����N�`�����A�'u�`�O�0�A�1�p`��
ҍ�o"*hK����g������Z�URLm���(�sag"��l�Fq<�8��G�\s������t�o9����V��q��?�N�M��)K�K�G�h;3��.%�)��l�h�ʾÝ���hK���(�����e�4S�r#���{�5"㭤�+K�+j��H�ב�����!I�:V,L����8d»$9q�-!��ݣʹ���b��2��'�����׸d��	Q"��|��y���g�C��	���0���S���<r	��a�3c4P�'�7V�ZS|��N�-��	�!��BU���(
H�idmZ�4eb��+-�@��iP�ؒ�
�KB�*��T�
Ŋ��dP�U���P��j!P�Vڥ����X��
X���
�V,*�*VYA��U�h��h��FTJ4+ZZ�����E�eJ�jҢ�*�D[[[Jֱ�J�U����T*���ڡUR�����Z��`���Vڪ�-J5-�!k`�+[B�P*4lPP��V�@F��kZȈ,�*��Z����-�-�+Ue�EE��m�Am5���KmKkU��R�Q����֊[m�(T�V�kR�TP�(��Q�F[J�-�P�aPZ�-DJ�J�T���UV�ҶQKh((�����I��5K�؛EX5n��UtbU�H*�ͱ\BZ�!�*Q�Ⱥ����M�f�<Nw@��[R�]3F��wǓR��U��Z�NCq���rSA��u�.>��f��T%���H�@�y���Uut+��m���
2F+7P�-�Xb�ܵ��2��{B��=}3� �B�&[�b��5`��e��_��ޗZ�N3�e�v4���.�X��|�	�=o�P0�hQΎ��'�oЮ�f��nt�&֑#e�"|�k��V��μ>|���<wG������[8����k�Ly#�.Z���%��f�������1~�u�)����,�H� �+�K<�/$L�fbث����W�M�]����϶D���
�.�a�:ҏ��_�Wᗽ����M�翛���m6�+d�-]��;AŁ3�xr��>ΧL���N��jEb�r�e6�5��9޻�۾��ޘ%�$Lo)R��4���^��;�Fe���k�ܘ�z�=@�ڙY����a���H�q�������}���2ϑ"���I�ݚ۞tê�@_�K���ӧul�CS�b({5��FxV5Y�^ܬR�R,���^Z��Q�/N�WTe�v("&�k��P�*��^�ioyp�d�u���܉W�S[S���1w�����+_x �٧�q":�u�yT��1D؜���O�H��]-��'� %ȊH�� �,�4i\��l�r)M���аQ=X��vp�[�/�i��6J�F�l���:)Q�/qg#������#�Pʡ{~J�V	�mi������X�R�O���ճIc�N3��(󒬍�=�B�B�88�*�qQ\_)c;	g=}#)>��!��x������U tE�$�%��i�C�������wX��t�\{��l֊ǜ�j^�h��X��{�֙^��4C;�`�Iv*��|\5�vQ��Vr�:}������}٩�[�Ffg�dO������H�,�)>^�L��.�	��W
q������p���b
��9��1�rj�6�󍴅����Y��~%��!	�q�v�F�v�Qڌ͐��Gu�n��NӁB;���)ᨿFۺq���d걹ngo'ϽF��O����gv����݊�R�جGFP$8�h3��txBdĲ:"wS��ю�/�r�o�����yq����au�Eč1Nˮ��L�	��Drad�Ls��
��+wo�P"]u�bÚf`�t�r�}�E�3>�X<�k��H��hx���^L�R�������ь�$���t�ku��Ç*��E��gRRɼu|7w�H���d�8ZA���H���{y��~}HV�(q��H-1�S	ݾ!^���ĕ(6X�1=Dl�ֺQSk&�K�������5��n3ltK,a�X���R��֢yԖ,�3��;.�B)H�A
���T���,�n��>s�T\<�>M<�s=K��l��A�X�b�E��a:��br*7���O�"�(V��*vՆ�\�.>�=�N;z�&ӑ��qc�q��U��ܚ�)3f��'p�Q
�����ڨv�%�*^'�i��7V��ꛬ�4Fvm#D(�<�Y�UN:5��xxo�9�Ln�8�e���Mނ�[s������ƻ��5��5M����P�P��@y��`�8Urg7w[޽9=3�hr�s&P�>�,��B|�u)�d>*�f���Rⷆ�x0i��lSv�o����yr'���������RKa�q��n��|����ԗ��ӽ�/��ܔ������C�+-@�GFB�K����!�+�+dTDW��F������߉��8�X�{u��rM6^1�2�U;?l�䲇Պ��H9�(+w�dO+���P绺%�|�����Q�Bn'��o���j����)V��i�t��i	j�ǅ	+b��pZz��]�,�yXv��L{GK1��osκC �ڻܼt�y�I�F�{��IKp�*���)��=i�z�r>F�޳B�íu�J��Rm�WI�.�o��W�����n\�pY�B�3**|�h{�h�<(�8B�I���_&��'g<]c���N���y�+�S}[����5� ue�*�1��:*����t��Q�{"y�L�nw6�S���{�.����w�H�[��wK[9���Z&Cґ|JI��<r&29dV�:額�y��R�Q�XY��ŧ�D��9[�2Քg��]��t��Q�'�C=%��rwr�̽1I��z�������Nz'HZ���>G��Y�*7��q��Q���tx���Q8/��;��z�!���Ƿ9Bp����a��Exblv��{")U�f+ �+n�ݧ���9�(�r�p��5[T��=�K/:"Ln����_R�{��\��-+\)��#L_H�{�uۗ����Z��3�p�k���d�^��At��z��ez�S�ʳP�v��&�AFn����pm� ��z��n2(ap���DĲ2V�᳾'ci���-��L�S{y��]$	����O��ޟ3�x꽦�(���b :s��5
7�%�e��S|��ڌ�z�9K''I�"�����t��2��
�D���^�9����m%��� �9�.�{��3�F�\K�n�󧷰8i�4!G@Zo��0ߏ>���C�|��W��ۧ�wi�O+�/�W=�]Du�c��F�+s�v*�݁��Pr7��X.����xn���w]�/��NeiQ�U���Z#ymD,q@��ܫ���{�	�C���k�s���xfz�6�Qså]�4�j]���ۃM�nz��Pi0v{�hx:�T��Ni���M64)����t�BU��������4t�9����ø�Y
�Wb,T�9���Ëڐ�e%�#&s,'a�YAŃ���e�~�$�yɠ�Uk@���%-�%a�/+w�y�6i�N�7Q�(���o]=O����R����©�:ι���.�pK]��R��f����lW>w�9i9auA�����< ��w��
�IҜ�&���
U����` Y�DO��CZ:o�9r�_mn�Þ�ǎ13���(�{��$;yb�\�f��|ϼ���BaB���HZ*R����[-��ՋVw����mK�{L�q�T��Jw;~. *u�DXTQW�sp�s;y鹄�#�ۛp�v��QP��d�T��(,77!C�b���ȼ 1�[�^F�m�/��U�)�f�*',����Փz���x��S�)o�N�uD�\d�_���W:��%�>?|v[;� ��+I�j5^z��}��b�a������L*�I��n�R�z�����]���Ԋؤ��
�W:n���t���h��Y-9��9S=Z����`F�����.!��G2΍�f��d&�EAqֽ�S��yWY��ϐB�}�@�^n__]����&r�#)�}��q�ΐ/r���jF�+imp{H꩹�~�'MoD�����UfJ��8�W]&��n��b��?2�yԓ�g+�|Ǹ�z��bU^���睍S��?��х����vb�������4G�W_i��[�t����J~�؆y���%CY�L
g�#���ϗ�hr�D]\�.���{�o���#����b�x@V	�6��u��Qk�L��0V	�e�}��>XR��y�=���z�F���엾�܏�!��S�Y�|� �(��⢽��9֬K(_Hěr�시P_h�N�nQ鹺�,tRՠ�;�bav��aqw{Y
�J�^�0��::�]�wY��j��̀�r���jQ�'.H!��`t��%�OB�}�/�k���b��.��y�{A��c�S�9�Yۻ*����?BWñ쑭�8�7*Eyd�a��
Q�`3Bz�R��331@�homV�Tqp��Y�j���l\��`˒)dL%1��.����/c�0�+�d����.�++b�a�J�S���>2��5�-`�ә��L6�Nm>���d۳��E:ݑ��pVa�%[S8�����^aRm��QX)���9S6��G�.�s�,2w30-̶�@�oB}I��jP)�9�tW<���%��v,J�зde�g0�r\	������׃�xj,�wA��#WhQ�"bz�kj�}u�;K�S�;�n+ ����B��d=����&A@�D6�LVޒ��lU[Wp�'ږj����'T<��J�����#��7�H҆ˮ�%�L�Dٸ�k@.�s�6��X4��!�t��f`��!H緰,K�̾X<���3�"�έ�X�hӛ}�Ew;��{��c<�}�,vKt*�A
��#�R�LW���g��T�V
^uގS\=F��ޏowi�Il0���H�U:B%�uQ�9�X��{�U��lO�6{�"���V]A�M�u��4+:�#~G4�Ce�OM2��g�3��װ�z�����{n��nC����Y��+~
�iզ��Qq��Χ`��ɸF=��`��"�ͳ\��(��n�ysCwx'�D:_���� ���YB��C�.��	���Ft�pk�@y�'	��Ѱ�ݷ�^(�g�_s�[��0�.x�js���`ysCi��z�$4S�k�zV$9�팾�^>׈�u��참Y�cd���97��]�\�+&a��Dr��$o1��W,B2���88���{�]�����s֘��K�Qd�.g\tR֤8�7w��Uxn�;��P�X�.�jܼ�.#Dh�=�VeL��-��;�x�saw-ȨCݑ�t�*ID�h�s5���]Ur9�}������N|�N��v�#��6;NݪP��VZ�u��o�MZ����\�/�V(��N�)����ss��v���{麭�Y�A�WJ���Wu��u�G���#T�^���)f�jq�=�:�k�.�|�f��w(#�FR�Wv�S�+������	^�E�^/���^
�����J3R���o�:� ����������t�K���:*wh+!頔�%g�X:m���Y��Mp�_S�3�.�ْ�>�0mܝ.�Z=�����V���Yd��օe=�Oswc��熛]��o_�S���A�;K�>G��D/������2�p���B�{�ts�(��5�ȢL�d�\��`*�����+;׸��fƄJ�=���^�������x��1�/�+a�aͿ}1��of;缮���p��-b�"(7��&��jl�U�.�b�v�)��R����БF;[��K(n��X��qxK�=�0}����������P�}<�e�m�U(�����3��$���(�ýJ��l��gf+=I�W3][�/�uVaf�|0�G���3{�)Y�P���/b�Vm:��4d�;Y�
�3�^vZ��[�Ā���'�+O�����t��b�Qʲ�g�B��q=S{�� ����ǂ��,:���:�]Q>�d:d(��h�l�'cNz�t�{�����3e��+iUv O����2x[YsGdV�J�U~/���:\�#^�$iN��~��٣}���W�1cݱ�R������R�^s.�p�=>��豪b6+O����7��M���C�WS�]�5����`z,��J��[��+k�c���'�����>v��x��� YR{@�msb���?Oj�*y��xTm��'�t(�T!ұ�>�I�<�<�+�^S��;��n�vfV���xls�pN��Y�����3d�/�v_Br%nl�9�k8ȸ�L�؉/���0���jTbR*7{�2�zC�[���M�ص�x/z��j��'o��
t��D+ Er�fqq0�J��rz��u��f;p�t=pqEo�;6�췒����n�D0�� �S쮺v�k�o	��t��9�m��Q�³��
>����7%P��sN��-�U�ͅ����\(�7X��/��^�K�ԍ���2�L��e�\�;�E�H�n�@8�E�\�ML�T�xE��7λ�a�:e]=�Q��Xй��EP9G)ѳ��c���lC�pz��@I.U�w+d�݅Bv �6��wM�@��w
{D���s�H��h3����h�[�.�f�9����S6���`�*�r9��z۠$'�9�so��7����BV*n�f胒���ē�ܭ7+��%i��!ezG
�[i�Gy�yZB��@*�O:/�}��)�q�B���5��کKy�sZ���X���R���r=G&�a��*r&'�΢Fr"bdB�~��6�q���X��x��~��'ئ����ϲ��g��'��<���z��lN�-�O.�Qs�ѵ^Ҟɀl��A�������n�R�&h��t�λn��na�gA�,&w�VbiJ�8=��3��T��{1א�v�p�p��Z�^�Y��c�xJ��BC��=�L|��Â^�����ƩU�`���Fa�ˁ�1TQ+5���������=k��c�Q�|�ݔ)t�x�]��C�X��,�������n�a�V���*�a]L��!�\�X޼͎��`"�ceq�,@\0�@�u^�*�T/l�`l^��ℱ�t&��s)kL��c�b{�>Z�{(��\({y]ic�/��H��*	���ސl���9*In^�e� �*����!�򂄦�[?��������E�Y���M��tXݞ]O���[o�ڇ�u�ם�-l�C�M�U����G�X�4j��e�$`6V��s/�ɕ�̡��&��@ ����y�Qc�6�f=p��n�QS2��f�$�}�l�"�Y◳��.�589*_�$T�"�r�j�>&1S��cV�ޕ���]�kibĐ�DW��ǲ�}&4xce�rn1q�6@ˬ�uueL6����D�M�l �=-�,�Owҧ7Z@�Ϻ��
��]X�e��1��f�9T���X^:���j��J�A?;���y���gY��H:�$׆���ݮ���&]a��E2�aQ '+kin��6��\/��Bn��v�7��\�P�0�0�����Z�PHr��j��q��u�}���(��f��ъ�t���2�/J5o��ң;�Y$�S��n�M�Ћ��aT��lgLȳG��\j
�5�3��upK�3;	u�0�����i���Y�p�z����� 1�6�BN�����t�x��0���ĭrGS�ƅi�����q��;�'��d�s�ͣ�y��::�If��p�.=�����3J�WSE �p
F���]�قV��v}��C�5g8u�$]&��&�p��^ɏyv�$�H�٭͡��tLU�pȡ�}��	Զj,Z��+c�J��O���:��G	�{�:]�>�4������0��TkШfw[���)�vz���������6"ʫ�8H��'�sv��wVM����#��=�W:�Ө"�����Xǅ������/�=Вhb��v���u������r�y	ܒ7�#��b~��;�hν�	N�p.���Ra���j�6�HӒ(.�uE1R�l#[a�������%g{X*e��X*��+��";�Zs�)�
� FYy�!"I��^�_����[�g���&o)��Lޥ".�i�8��s��WaQ�%Z׶������
}͑�fs�o=�wN�������L;.A�Am�4������f��簄��+$T6�'k���c�Oʷ�����=8Q4����������x��E�7���ػ
�a8�.��J/�p���R�Q\�l�'����8t$[!�!8:�
��9T\V8��[@]-
�Jk_qs;��_VxѪ<�tG���M}�N١+pَí§b���q�_=Ϲr�ޛb�M�3:
k뫊L�n��.eE��$�m3|��Đ	�H�e��,��R�-�����KR�R��me�b�T�Ҭ���(���ѵ��XR�KiKA�Tb!Z[QE,DZ�[Uj���DX�(*[Q�KE���R��1Ub��XT���2""d�Q`����)1��*�*�[IeJԩZ)Z�ƴ��h�h��l
%�b+"Ū��k`����������F�-i��
(T�*�-��[eEh���J���B�-(Ŭ���"*���V(�%�"� ����UQTQQQ`�0YVV
�Ԭ���@Um��DV[E�dkT�(ň�E��@EAdX����1`����K��QEQTEQ�ER,�mAF����"�U��D���",����̼�P����̧)�Ý�S�X���VTn�t��ٱ�8m�s��W�@=�S�Rw�i�l�k;^I8���e0P.���iq��5�S��]��vã%�ȥ�A� 1x]f�fB�:gk!ZT��S�����m�B���Qseu�7�;����08�3�t"Q�3"�H�����j���mi
ޔ�F�^�@�{%�p�޼�Do������sH������Jv�v���v��٭�$v�꬀�.9gWl��EpL��s�����͞llș�5,�{�1�;�D0\�����(��0�s��P�����vci�<5%G�Tj�U���j�7�sw�BN�i�L6h]m<��P��|0HP'����6ޙ�%��h� ���Ws��Bس:���.�C�m�"|P�����.61�.V.ӛG酊��R�ֽ/3e5�������A��sYA�� /�ѯ+[#����`��p��|�y�|3#�O%���uڳ�7:vg���0D���9<����"T�$s��l��>&̲�C�F{;7��;WS��
j{�U�T`' Z!��:��br*9��3��<��hW�{��ϖ�e7r�W�Y~�Q� ������/jѽ�6�%��M-�Ǹ��6!�ג����5V��e��9ϠL.v*F�lS^�Mǲ�Ӣ$��NQ#%͡9�J�i����/�T�=\tbJ�iCR�s�p8�,���\]v��p�zB%	/XY�vD[��5�x��Dq�\i6��]���gO/>.���L��B֞���R�����<b8B��0%el&��=��Ch!�DD��]�:.6([��X�"�p�i�[�V�ܘ-ʘ{�TE�}��N��Q�Y�|�
#��ޕ:T88�T��w�K�}Cq��2�}��VJ�\Zw;�Y��/���Ai�Uc�d>*���ڔ���v�y�\���9�얍A�~���QYs��}"�.�,���'����O���A�4��Ĝ��
p�s�w-��ʞ�V?	��t���C�ӷ�T�ܬ��P55RT��ގ�_*���V7hLN.���X�@]�`����uֆ�]�e�6��� �2ٕ��G3w^1�J�-���d.�cN�.���J��(O����5]�[b�.s�hS\X{&2)�ECrN��ҕk6wY��B���s�uo�*y)|nGN�s!�%/�X*N��pF�*����Q�u�=��Ｗ�<0ЗiRly����lOH�-K[�;^���%zG���E:�8��x�]�!;ffGZ���w>}��Ђ�FW��'��5lmfc��v�y�އ(�f|�P!��eK%(��紉w`P��^�`��8�턡t����L%naH��{�T��Blm�*�T�кOUΧk�iz^�5�ޞ�0�e*s���w
N4�gD�>���Lumc�n�5h���k��VL\���i��vj���]F��b��{�.����ctf�课.�>Ouj�o��c�#�x��Xw4&"�DB�E��;�O�d+9�.3�&�/��ZFlK��v��T�3aT�E��6V:�]����5Q{b`n�UT�ȁ����~���m\��E�k1Tc�r��r��ȉ�+1]��6��R�yzf�,+�x<�J��u��X9C����T����+Z���qxH�����6u[��'�uMb{�]�`��{���N����p�K4�c�'`P�������(!F�A
3S�g�u���\�������x�T���(e����� L���mL=�El���^.������͖���j::5T����\P	ͣ�n����k�a;=g�Y� h�b�WB%�;ljP�/b�X�[A�¢mHz���l�k����	g�犥bg&`(jX��x��t,�/˦!�S@ܝg��ҙ��J���ӄ�v)0T(�N]<"kL�Yie���v����5��4�*|O�*�g*a�͵W���VVq���(���ϱ=��]�W]>6���ν�Q3���ԣV�JT�*��3	ۣآ�ջ�;Bn Ij�%s�q�����Ev_w���TJ`���t�B,R���P���*�����L�C�U�W����c�ެ��7�V��+>��G'���A=^��]Oqv+(�Jpn�S�L��絺��b������%Z.�,K0g�z݆L�Ց1	=,���#!a1{��̯?x�{7�
��;F�D������4���'^�Qi�\����x~����;rT�Z����O\���Xŵ�,G�)�������	�N��;yb�]R��%��Ʌ	9A�;u�vk����8�4mf�׼�V��x`��8
;��ʙ/1q�� X�wk�e��cqkT|�Ԗ,4s�?Q͘A�F�υy�*�^����1�����,��DI��yU�=��n;Z4�������4_��ޙt~�«*{�(*d��n����9L^jX�>�D����b��mDP���0���L��՜��*0��l�	"D��Y{|a�E~铲+�uܹr".9��-z�4�x7��d�!�
�vh
+_��pg�x�#��F����u���Ig,H��;�gZr�`�Z�P�&���֜��G(8�	#o�7W4��A�h��7��t	.T��ő+r�_Q2�vt�f.��%4�Q��Z%��V�#���;,^tA]�8��ҧh�/������om^��4�---z,�9K5k|��<�j�v���DfKˁ���S����|���/�7���O:a��F+�ӈ�:y��dW)zVs�����v�Kŉ��ok+�&�gp幋��<ȋ������t�e��;H�0,�]Dwa�3ܥ@5=B��+��R�B�����Y3�ddez%�(x�1k9��4�ۋ={g�skm�@��N�+B֧��,����m��[�
2
�G�I�KG�{�V|�>������M�����X/�aH���stf�k�+�7�;����08�2���,Ug��M��a�̀	�aDA�r.$'/�F�K��v=���5*F�Mn�b�ڈ�G�&���rOVm�j�+�����˅8�{#v+]��/Z����z2MQQ�NJ"�y	N���J��얇d�wkB�bs�=Tq0C�L��2�N�Va
�i�����vck�)᨞�
7���V�Z�/�(4v=�O�Nu�pq�8��V�#�+�$(5�`NUq�ҙ"���Sv�+(՘���������޽KjPKc�[�Ué+'���]>=�9�g��i��G�gJ]�4n{�7z
Cp1qL�U�*/����۽��f/_>�Yi�K}�����c˼#9��x���9'Ҕ��-.j_ُ5Kct�L��oj�m��^��T^V�1�?}^��"QQ�u�f�9�u��)����j휮�*i��f^)d��E���T�k̍���@�\�o��R���/�6�zQ�N�P�}�c׾�fh����@DF�;ʡ9Rf3B�|H7�qpby�}7�3P�p�m��آ�l�n�*�:�J=���f�����f	�K�ʼO�y�����A*����_hٻ��z������݋m�D8j��PV�rTD��e���#z��]�i4�YފH�ӡ�Z�b�D�F�8<�>=kE{i���]C��u��}����E�Ƕ����]+峆b��.����̺<�����B;o 5���#��uX�zi`�������5:��,���a����x��N#�Q�����.P:v����i蹳��)�-�ͽ�A��򩋘Sػ9�`^��Cx�yx;�<k�T�Q��3�"x�˕�䘴���)0/9]V���i͙�v�yhR���F�Ӷ-R�`J�P,GFB�A4h�r�[����d��DLws�rH(�����̛���8��c��wMXy��*��B��G�Ύ
��v��e;��/f�=��3y�7jQ�����e�{��=;��ɇc:�`�YF5�S׽ر\���-u³�c �z[�R2�I��N��gG�՚7F�x`�g��	c�u��t��ʖ[�"���ݗG�؆ZJ��x�/{O���>1h;]��J�U���+�o�q����h���$c�ݬ�����mu�;o�����P���k��tn���V97�i�w�mE�^X�ط��~$EZ���a<�V�y7˳L���\,�} Ul�AQ�tB���HE*���dA�
Jv�= ���Nz'H_yP���Z=�!P�f@<�G�ɡv5���闍7�gOJ�.��2�h���f©���X���R,T`m��V�)ᙏK�Y͆�{��)
1�υm�����jd�{�Y������>ۦ�}�l*��4�c̆������T��`Ѥ�^��pQ5u��\�j6����['Z����o	�ֈ��Eg��Kp7�YN����fvM��o��7'`P�q�����@�C�2@�t��٥s���Y��V�N��K���+?^�W~˷g<����\^N��U-�>.����!0�ݕ�E���6�	��
"U\���M� һ	�w�RldOjC+�R��lF�2z$��G�j���5-F�ب$����Z��U�n�d_un���m)(�c� �6Ѩ;1�q˖^�"_:'.;�g&!�o8�n�lKB��-��}%ZI��e	�hxܴ��1Æy��}1��h���,��D4
�����B�mu�Z��t8�-��s�ک��ϲC�Q]��R���k`X׵<G7;����ϊ�cA�y�����hsc�E���n�2,��K7MV_��ם�,��a�{�"�:)j�����;��9
��2镖k�\ ���hpu����4�Zv��^+�#�t�
�'{���y��:Xz�I�z@W�q>���l
��o
<&5\���A,��a�l��+tu͛�c�۹�x�T�
���8��(���> t�k��;�J;uux��=;�4�x�I7� v�����J���t���	�b�`]
�iU��*�t��ݭX�Y=����u��e����B�d�Pׯ_�/��@���ȕ
���C�WM�=�Q��i_m�jv�*��=kv-�V�L`�D���	�X�S2��E�73��nZK����C�S�87,L���!eHpH���Òb�N� ��P������T����l'��J���î�Ȯ���[���
�ó/.�*&�c;ʹ�=�Y�|߉��;v%6o�u#�}DG�̦֡���FN&wf��,*6���ܥ�֓o���É+�{CS��vN�Q�al�v�:ĳ�7�t���	m��Ӄ������.z��LF`�]Y�^yJ�Z®to<�ņb�����˾���y˥�V��8��{ʹ�O����o�+��<ub�t8yk�Ҡ��3�q-��5W�vNe�1f��6�eƯ��~��*��z�#0ׂ��ݛ|�{o�~�&lD�;�3d��Vk��J���2���"��=iT����個��8'՞XR��UfJ����t �3*��I&fw��S���C���w��>��W�� {�Fa�/ )��SK�~}k۫:>�OCT���ɭ�� Oec�'����E�+��+9�[�z�茀�l���Z��+msv�V�F��{(F�E�Z��B��V���<2����*��7����fV5���ܮ�(me-2����^K���Ca�9d+�f�qg�oS�;�xz��ѝ�p�01堜��m�a�u���}��*�Ubմ�
T3���V�[�u�yo6e����`]��G(�1�q���a�G})m��7jx�r�R��~��Ȱ'w�eW���iq�,��f߹���((��9��Ҭn�{�4&���M�v���u�K�O`T���c����d]��o�}��c's��l�PWBW��l�gJ;�������.s/��bլ��Oq-l�to U���pWm�jIR��sJM�Ae�P�F�_�O�q�*.$b��Ѩ�Q��Kt�;�r�X�"ݜ��ӹ�z7�<���u�����>^��h��j�%Sv+h�t�Bu����ۙQ�N\�7w96�A94d��qMG<��U�H�/�#���Gp�tQ�����
���k�r�
��=~n�lh0ŞQb��2�PH���{����`�ІR������(���L�E���w֒����&F(hIw�����x'�^܆]^L؜ܺ�F��N��6�Iޘ�rq�Wɸ1P7*k�g�6qT��"�}�[#��Mt��0T�,�Ss�['o�x��{�{;�T�jn��yP����U5i��;/�\q3��Ni
�9MN5�y�x�_���3U��x{Kgë�H�A^���Pt~�V,S��}�r�_�o˗�{�1<ߠ���ʩf���;Ɗ��,O����#~�U��װ��
�vr��Q��W3��Bl��H�ȵ�֬|�\�V�\�|<�oÏ��q?s��	!I��B��	!I�XB���$����$�hB��0$�	'��$ I?�H@����$��	!I��$�	'`IKH@�l�$ I?���$�0$�	'���$��H@��B���$�	'�B���(+$�k=��DK�B
 ������I�*�)!* ET��%�JUU*UJ �"�UUR�B�U)J���	B�T���D�T@)�$	4%PTR�T�H�J��iQ
R�E4є�*�T�SX��R�Im�(�SYJHTA)D@єAS52�ri!)PP��H� ����RDJ�(����%U H�B����UJ�P�I*"GlH*
���P��ڄ����  ��f�m��kV��P���k@R֫V�F�[U �ګ��Z҃j0P��5AD  ��*��(��T�#K� �)Z4R�ZJ�5V�������2�T���l��(V�� �+5 �����U
D�l�QT5�p  ��Kj@d�j4 ���[
Y0 4X5�V���J� EPfʚ�3`5��ƴ�a�b�)J��R�*֠��  ; �j�`�I�@�k#�(���n(�E(�Ev쳀�ht4(P�C:�
(P�B�(�"�
9��B���(hs�b� P�P��D�J��
Hn  �)S�3*�L�Zl�h[jЕ*�Dhօ	,V
�)�J���*�F ��S[kj�V�؁b6������)UJA�T�HH���DV�  wkJ�[aL5���-���J6�Z�Z�m���L�((���R�M��2[�k*�j�a@i�(��-�4�P�Pd)T���DEm�   1�B�mYf4Ҍ�QX�`*�iXҪ��L��(ST*�ʡ�ZچV�����
�4��j )d��Mdh�IT�c*H���IT�   �%SZ���i�b�0!���BZB5T�@�33L(B���M2+j�T���Hc�5Kh-(i��c*����R(Z�
B�Pm��g  u�@L�YB�V���[5l	��Ҁ���H4he��SB�!I���P�mj���E�2RLh���m��T��D�*BUT���  1���6T� bղմХPV�+i���S5�(��STUh��JP�SdXDV�T�f��U���0hPQ��� ��*J��      S�0��MP     �"�S!3Hѩ�b	P0x���T�S�A*�       �&��` &	�  �H��URj  4    r��.jR���iz���-:e��+^���|c(��"1{�)|W,��y���PA\��`�Ax��� �"�PDAY�Af��g��������U	"a�K$� I?�� �:d5$�W��w��}$ �
�F
"Aϔ�3t�� ��w�O���t�V)����Z��e�1㴍�M�H�&��$˓1�����k@$�J��OL�!�FD�zE��x����4��a$�J�;Z�Y�R�+H�(U�F��a)I鵮�(b6~M����k-�I\�]I���+O�
�����OUC �1Zv	æ��hY��v��]��,�)�qà<`��,4�q1�N1���n�ej�){�zfК��l/H�9X�·X�R����֑��SukQ��o �(kb�!	իpǱ��D�&��g�
-b�-�q!*m�$ �v���b���f^*�u�%̬V2c&�L9Jc�RZ�4c�ݼԌ�����w+v�n�3j���!&��7 �nʹW�^ �*Z��n��Q��r��n�9F���@.�7���n�4�4�"kB9���0����(�%����˻�sV���!`��F��i��ZZ��x��������ĪM or�+wkqaJӣFՃ���&��جcR
6C���Tƶ7NJ�zثna"�i�6��ȶ��а�{Od�M�%�kA��G)��~՚IX�&��Wc/�+��֨iz��6��q�y�	�A��O��!�HHYvnã��%�#$�����
���ӧ���M�aYF�p<���E���.��ѕx���&f�(n%*�V�7
H�!Ԏ�v�w6���f�Vwg��J-��K��c7B�P����tĖu_�%�P�j&�l�x�O�%$�
�V:�nQvo�3E(��f m*:/j�ɒR�b�ݫ���zp��J��XB��B�C���u��P�+��+{Od���d�o:HH�t�����1�#�2ȨZ�ekW[nCj)���1
�+@��f�.V(�j�.��1S��(����� (�5�ƥ�j�^�ϳp�4�[G��l�1���� hxs4����YYr��j��%ڙ���C1Wn4�U��:)i+��jZ4rZ5�ͭ#��ZT�Q텭«+Yz�9���f%�F1�pAz�p���F��X�l���&�-b�CB��2^ݯ�L�5���X��ݖ�Ilټԉ�Z�Tm�ʆB6��8څ��-�0�4�VX'`�R�/$��iC3R��\5
�-�B,:`lfR�
��t�,�3a���;-9���3e��E��۔ò����U���Zur�M]L�*��H�L��B�[{�.� jU�ÖN��h����n��T�Y��#F]F��J�����{��:!��3@�>��Hͥ%KI	��{j!p��0��*$+��XB�Wm�Ճ1�,�1��t.��-,F�6�S�VN0�p5$a1�Y�
��B�Y��65X��A�D�����q�Vs-�cC	�޻5u��<��`�U(J��Y�@�ri�ySnފ�M�*�^P��U��6��7T����"ҋw�j�f��)lD�];��Z3C%�k�*�B�� �VJF��ˣF��.�:m��N��ƮF1��FP8 ���V�7�o(�U���[�m�l�xe#F���&�	�m͑�"@�:Xj�Zж��	a͙PP�ܗ����,�F��Z����-�y��e�6�LW5U�
X�:1��U�������M��ܲ���q�r��E/�Jx�9m�t��5�9��^�bw�h�eGCE��������1tX��X�� lU����]I{J�D�VC���5�h��k��u��ݠ��œ)�ZE�;r��,�+�r��!��*�=�p�iF����O���Q�Jpe�u�U�Ѵ71V91#��'J��&��Ũ2��jf����@K�cQ4wM;1KX �e�eAbQZ��!q��ܫ��"Ζm[�PDkla��&�ESZ��J�Z��S�e\��YF���Cv���t�ZT�n��&������]=2�(F�<j:�k,����Z�q�^�2L��d@ɀ鼐좋S���ք��MS��=;.�ƅ��ݕ�ݱ ˹8jJ�ܴʈ �۸�^�f���d��(�Q=�wPPa36�٤Z�L��0�g�^
�&ur��7�#'`���&�R5����iL{P�,!���4ٌ��) (;�ب�x�Wbfc*a�q��v^D-9N�wQ��K`NZ��f��4�fRq��K"򅈘���/yD�m9	�Y��V�۶���� O/Y.nG�&�բ�fSբ�c�]ӺW�si�Zu-t�V/sT#`.�1�mѸCk��U��=ܵf�H�嵡J4�[�����$�;U/
a��̃N,͖:6 U+B�f���y�h��JE�A6.�Wueim��[FVCWKp�e��)B���ʴ"�:�>��V
�8�+3N��� dsB��5�ZT��d�2b�Ŋ�=�'���-��x�cvpJ	��G�tO��ɱ�7TH�n�jXJ���r�q��[�������1[;f8�N��A%�j��S�l���v�;�᩷�z���)̩����P�n�$6�eX8��1����Ku�l�y���f
!bZ���3d.�6�F���]��W�hȰYn�niz(��5ĪJ��Zgھ��jXŘ�냶_�;+$����I*ϯ�͍�D��l!a�Z�㦶��+r��^��O�A���mf���ѧ��lf��vtG�8�G��5�X�f\Ugi��h�Q��L
���2��ĥyGM�Sq0v�`u{��i�TV�i��)9����,��"j ё�6ԡ�'L�:�Pà���oMc�g2��@���Y3$�J��P���M$K2+mR�.��]<�e�ע��e�U�
�/���U�2���Nݰ̓����U����V��k(C�a��&�ۘSx�٫�K�3ڲ*P7>aD��^�)�N��]��Hv��Jk��Ai��u�}z��֪�[� ��.-���@T�˓pe��qM9�t���*1�u�coK���Hq��a}��1	�hhɷS%ӕ6�4ݘ&�f��_Z��(��+@Hk]�w�	�3tJn�&e!Cf�E��E9v6��E��-�B����,��T�&Fv�*���zt�R���ݞ��}Ԋ��Va]�Y�#dJ�����ͬIj�hխ`[���'Mr�4S��ˈƯAT�R�~8��oJ�yYX�Z��sSWu�3t�Q7�8V���E�N+�i�iwY[N�5�$y����)�8CWr����h�)������يh.�(�;��i��ƶ`��i\�"[GS��n
�^���Rb6^�sa�*�ƃ�K�Z�t��%t���2��յ���sKw[�PN�9�s{$���T7	ݸ�V+(c�MYG�싆���^�Yv���:�R�m\Tp�n�!)4T�4�n
ä���Z��Xn�'����l�خ���u�&�;*�V�B��?���òQu�G��,��Yt`ͣ��sSxc?f^�W�;7Y�h�j�3@�JY.��nFuRه5�qäj��������:z�
�r�$9�,��L쳢�n�6P�Bkt��ov�yt�r����h5��`�@�M��]��u��m���	��ԯNe��k]�^2�[��!�x��R`��]\��+K���tV&pTnɨ��ë vƻ���[���ɹ�]
t��܁���ģ ��:!�ҤU-��×X��o6�����&�	���������W1�7q8�/6Fì���ܤ1�4�7@�];���>Mjᐻ%X�6d�Nf�{oA K������3M�d�*�%�k�ܳZ�w\ow,䢵�`;r��d���X.���+�`��ݭ�3)e`+!��R����
�gFctrՄ6'$"�l�Ub-J��6Y�r�Ĺ7x���O��DV6�טM�N�[��:r���{wb�!����:�;�c�ɔ�z����shLN��2͙"��iE�g-d:��(Zp"0U�MhDaGkq�c��,ǧy�Ca�w<��f��v��H���[Xt��u)J�ll�1vp�n[�p����.T�J�Z������z�[���n̼�
�q�N�5�1�Hƭ_�# �94b��3@= �\͚�w���,n�*;eZƝ�W�Q��Qf��A�.���E�G{���N��_Du�M�������Z6U�+jd���$#NVb��{��Y�]�c�+"Ӗ��ͺI�#kp)Zs	���@[��m�ݛ],��l�Kp�n擋h	��X�����n��l�.M�1eD�Y�iZ0��8������f�jM���h�d��
ݸ��%E�骕^���Ub��L�O��v�<p�-���s�iY5�d��؅:�2��֒�ޜ�����/�9n��2Z'�$��ʏ3v�1j�
�(o,�"1��X�h�2u��\�v�oV%i;J4�۱���B#h��;�]P�قŦ*�"�	D��2�S	�E'�]����7Ҩ�5N��X(���[0m���w���(0��YE�	e�+7k!5t��I�.�y��F1��y��/pn34۴Ԭ�m�!0�j�vv�ґW�6�1R����)^�j��,F�M�b�A�Oץ�q�x���PߝmY�B��	1C/5�K� �H-Ө�ـ�*��ʙ�,)��o)ÛWD��,�Ew����6cM�@�d��/U�ud�v�Z*��I����X�]nUl�	��@�kP�o[o^��42;���"�;���V�U�)��j���V�s6��m���h��"N�Mbolܣ��C��*�{&5M�T�lk�3�f��rM��rѻ1��2��ҙyAg��ٱ�������ne1����[b��&�U��3zΨr���2�Yw�����KC��0����96yokM�T�~/(oQ�4�%�b�,�F�YRi:�[@jR"�" K&cE���-_<�j�oƳLڗ�Ӛ^��U�۵vbMt�fA68��D1z�8,���D�B��ʠȵ��`5Kr)��cߍ�ڹ#��܅4rI���t��ZT]-F��l��P5��6
#jI/p�#ofM�zYX�yY�0�B�V�͎�j*�����P-�ȭͳH�Ƕ���PJ9�m���Z�a�b�?]hT�X`��v��N 3����CAl �F��K̀��XΓF��w��9����ܚ���A$�@�����Ry�z\�.���B�2��WCUho�N�nf�᧶��!2�(���Z�ZaYl�������)1���L��(]j�Gh)qh�ҳq�U�7t�(��#w�3��m� u�#В5��G�^��V�z���kob`��E�-8�j�����;���us7]:um�6�9[X4V�h��c0�k[�n�����LJM헵	�]��(�����F�ֳN��dJ�dI���	(=&�Q<R"�\�U�0�	���B�k�ఉ
���swiѩ�0"Ƙq�퉺�CC�ϥ�%��/%TR�N�mɤ��b2�Wvj�ʘ��ad+J�Q��n�D��� R�%nY�j�e���6Qe\-��/5f��43E�!Yp�%J��g73�h�;�/,�:����l��$�]�0Lx5��4����H�%Xy�{*K�%E����jLՀ0�fB�ױ]Ja�{�0ܩ�&�iiXU��L�{��+/M�͌���#$j�~Fd�V�z��$]X����B��[ ���7/k^=��K[��I��)��`9i�c[q8��&]��Mkd���"�av�"^�ޫ���gouA����ћi*E�u��P�,ͣO)��];9�Z�jB@F	���ZE�{��tL��4�e�zY��.��1��72;�#A���i�}61�w6�M�Q ��]e!��/-=�`�4�6���.��f�} �jGH�oUrM��L�AU���p�,���o^jUYvB���@��	y%�k`ݣ*&֥�
�wghku&�Hų^��۽JJ�[E��X�d"R,�&�(M ^��U��X¶�	k�Tܗ���*�`�hU�����eaw�C.���XF`�V�A"�yZہ:��� ٻ{rC��@�t�{b�����l��lcD�Z�d���m�[�Vv�/k�*�NL��Y"%T��f�-F�����G��G��R��mf���V�|��Z�FeYsM�eX���ڄy4
�f�2�*�5�5��@�:�ԋX2&­!���]��V�]`O,*��wY �+�ɷp�(f�D���]Qf���;�s7f�(c��x�S"��e#�*�C+Eй��1�b�3pݲ�`Qb�*��f����Um�P5�qQ�/7�B�֍P�,��T.;n�,Z�H�)�IF-m�]v�c�.�7���hhT	٧-/��l�*�Ee �驍Ve��.�՚�Ӕ�kZ�@U�&*ɍP��+�w>���M�Q�����F�%�Qe�Xݱ@�1ֲ�w��2^��cߥe��W����F�ʸ��DPJF��ƭ�5�q�up}h��<պ54�c>���&�)���9/KVD�۩a���ײ,�!L�����ǘ4���5�,ӣ�+�n�B/$P�R�ja×a��hl�Z�c0�AKǍ���QH^i�4��5��U�X���kh-��V��ӂ
��K�Z�`^6t�B�X�߳�RR�(nm��VZ�H\j��忐G1G�(��ĞZ�v�%�H*��)�ư��'F��n��$l��*M��{�e�&Me<E�6CV��]
G)ҳ�B��t2��pL�`-FA�cJ��A�h6�eK��Iٲ�-��IR�1y���6wV���9�+ŢA�I�d��4�$m���ٓzԇ��y�L�N�WL�\�!\��Ν��\�v�*�uk�S�[�Ȥq_/�s����-�JC��8�t�/�˼k3p�E�{H�=����u��3x,�����,���,<�<��珨=�\�2@Rtɭ�[|6���	�;��/0ViVOte键��V2��f<��s"q�/�8�}����N�\��$�#לJ|Ӳ/�+�M��� {�{7uB+a�����S ��T��9YżO��-�K|����j�c-k�qm�4�;�XMҡ)d�]��%V��"Ũ/:�t��Q(E]�|�D�J�H���M]�ˡ���oy�j!�,����J�d�u�5�/�b�����*����:���r�lC�J�<���rd��]ޯ�G�+�
��������;���K��n�f.bɩV�cܨ��eM�{�0�%�o�Q�7�}�3U�L�x���-�e��lP��ݙ������$6	�u����Ҥ\GΕ��o�묫�ޙ�hSj�ۼE<��ԧ�I�9w0�������4ֆe��Fp�h;��S�r]�}�\�Vj�b�u�Hw*p�g%Xޜȅ՜� o_wm��� ��S����*��@�,LB�n;�R��;�y��RK/��w�ICJO
:C�]�]b�V�v�}�j�$@�s��W�F}��$d
`�ߜ�g� ;M���;x�!���ns�#��lH����K8	֮�n��7��0��W2fd�hR�HT��k���)�faи�f����#=}#�[��#;�J�L�\�_d��x�-M���lطef��ɰhc��KxU���2:�G`5��H�iv�v��0T��P��t�H��&
��s��YRa�?6{�]u6��y&�Te���go�nՍw ��{�5������xT��u7�=T�QŽZ�J�-��*�˩G7���Җk�QB���h�)��޽��D>5t�d꩜����6�wVLOC&,�s��UW{Ӭ2!��z'Y��
-�<�K{P����u$̮rJ�Y:.\���G.��.�����޹��5�'W����0m��+��I<�0X�wL�����Y�ƕ�;]h]v[(*��l��{dS{[�����Zk�Mg6Bi
=g:���{�o�d��(���X�,q�V��"���f�` hu����|��ALu\�#u����St^U�ь]�7Mx��t嵎��Uqm�Y��O8n�5���kkm1[;�<$ή�����ם��k��������Iءu#���������ik�v(��EDeؕՓ��e�Gb�
t4��a��Όü�eD�iʱ�3�_)9��vom���8$�(rХ�k��g���Q��~�is��K�U�p��{O�����6,�2�%xB��ܪڎ�օ�]�P��T�����\(*�mn�D�­�&�������z���HA���}-���P�ɖ@��}���9�Wq���M�@��y@ܕ�Y������s*O�Ko^H�!J�a����Sgk��$l'S{l�e��3��ܓMlK�^��%>��&9Q��#��[2[ٙ\��:]���oh�e�fp8�U��1��	�K�p���A��G�[�	���4�n���fi�{X<��e�M�z[.b��h`rU��eP����4���o4�V��m���҄j���B�T7&_W�+��r�x��%`�/�0�1��'P�y֓��&;��i���}|�^��N l��
�@�'����=�N|��N�����oXx�!KC�Ý���]�T�Mg�Wʢ
�C���Q�@8̄�I�s����\z��ü��T�]�9cُ�n�{j�n�Z�Q���K2�4� 4sU�ij���jl���R����獛o,nn-Y"�R���+6���<���y�a�r��[��=/z�z��{���E".8_��q��Nd�Nq;a�:D.�eƞh�\*P2b�n�
F��3Y��j5:�L��S�_7�����{���x�Z�+v�xD�ӗ�":YϷ+UI]������ZvSX�a(&GM��))mC�:;��JA�F���d閧m�볔��g!�Vp�O��V�I��c�_v��v�ܹ�����avI:��b��J����m�|A�͑�1+�]��]fJl�����gl�b��lQ:�n��(Ax�97dS��V㕻Z��#��!�Ε{�W�{ZΧz��0�����h^�_^9�ݦ :���.���H���o����X��0�'k��4���]�}Y�,�s�2��s�jy�0����z�ŉ9���L�&�T��{$GP���)n���ޚ��,e�L�d~͢�g�n�u�9&�f���r�28�m���-�.�E��T�ᤆ eskx'yf��ΛY�e�T��W��݅rW[���iL�Jl��0��-;���9��e.��,Ӗ�6������b���h��ܵ}7�v�܋E����ϫ.s�A��|�c�ݵhuo:VWEF��tz��Rݹ;���P|4�%��k��v�)ccB*J�E����t��/xMO:�2m����]`��%��\�Q+�nEyҶF��:0�t�gr+�̭9��g����g��ݼ�)wi6�\X���Z�s�c�o5ZT�����	7��<ky:n�A��N�v��&d��l�]@s���q\�O��)9Ժs蹴:e��Ϭq���n�^Ю�}��Q,/XgX�I�GrSRK@���ι�{{	Uʎ�0j;���9�h�Q��iɰޚ$|�u<���9�E�ٷ���&�uY[ܞ�ɷ�ë��kp����sN�0��9�늝���`�zt�Ɲ��5���.y��͕:��V��m�8�o}\�z�g1��Z@�^���ĸiw����#m)���Mv9D�a�����lYo��s���5����������B�/��3�x�gK�p�d�+vt�6��݁�q�����4��&���G]+��6e����ս���͖S�x�_��1eȪͷ�Մ!�M�&�9u�/	��A�g��o+�`�����ɊsE�+s��j�w:ܠ�p��ݹ������u�'�!R������f��Q<o�#g5YϦu;�s�˞�nu�VY�P�*��"`������S����Բ6%݋�]5}z�s��;�*�[��W-��#g����0峘����o]�\���iv�Ҵe�������_4Z�b�s��:Ҳ僙��[W�`�C�$aړSTi�ʿ�@Rٲ�Of�����˜HU�:�n���������{��-��O{�4��W���Ȼ����߹��4a�=EQ��5}���o�B��ңs]<9�9,��W�U�]�(\�
8>�`Χm<�����Ev�4p���r<xE��,�����'��j:{��mtTt�
��Y�Y̨k6��uu��}܌K��aۡ'�0v�-[Z�vZ�O)��nm�,M_ ��~�Ó��x&bﻵel�p�oP7(�|O�`��V��Чu�����9:�V}9����<�d�}3u7��t��v�*/h|{a�钃�P�W}����7)�v���^�5�CZ��f��t�9���o��(��C�}������7j� ��9���Q᭾
h)����,�Cq�����S桬����$��:;�Fa](�l��0z���'Wf^+�/��Co�Wr���A8�P=+�)	���(����N6��z�Qa
0U�m�a-wƎ���Qdb�\]�@�"��m�΅܌�x(�5u��W�ՋU6�쉧�o0��ݧ�ُQ�n�(�Q&��m�xf���}��-�n��bO����V�ұ^�h�O�+�5�����_�sj=�^]�ݭ}�CD ����x�>�v�psX����6r���ae
"���j�f�и�j�S����U��o1�vG�Z�U�;����NT=��:�`��v=�w]M4Co��[��^et�A��'w�8�nNB�]n��n�v��J�]����}7��.ʻيݝ	{����9�w ����Dj嘶����R�C��e���XAe �a�!�{o[��{(Pp*I��#6���j=v��k�ԾZݎ��Zz9��&\�CiIXӂ��_m�����Zz�%�^d�A;X̔C��d�j ���*fQ����:˸U
;z�J�)o6��rVL�\k42&�]EKrX9
�W��d[�bP�&U�����ar�|)�tQ�T��]�-���$�*ܙ�������\��˳3�˱Y�N���t���|k�%*�`�s��/��/ �W���<�c��HT�M Н؞�6.+|؃D�Ow�f7�n>��� ��m^C���ŏ��F�v��.
6�����ݢ*�e'g���^���ɼ�ۼׯ'����z횦7���,C���k��Zڹ�����F�Ob�.ٽ���������fܼ�&�hsڸ{�ܻ���Lsh�|����u�����&��c�S<x���d�WJ�3x;r������n��n�L܂r���+��mY?�,���.1�)]��o�� gW&�sWZ�=֒���
��'��IhQ罭k��ì���N'�ӄYݦ5K�".g��zƻ�%� U�q����ְ�W�˷/�h�����N���[f���<oI[�d���r_Kӓ4p��]�ϗ:�k���vjD�LWD;Č�vˬϹeg5:���wf�[��n�OTӫ&w]R�.AJU�u^�(n��`P"�idf�Ӂ�n,٢���W\�_ ���R�\�ݬ]X���y��2=��y��WZn*�����Y��j"�ۺ�'��@�
���lp�ۨn���OEW�8�7��l�������WIP�^#��bv�2(�>�ﺥvU���"�VD�(�\κ�E��\d��k=�^e8sw_}�L��9f�μ�usA�\Ts1o-�q�Omݝ���a(�]nO6����oپvގK�m�f=x�9i��w(z�+WSg]�|�d�/�*m����=2֫Z���3z�ӳ���S��.溳�X�6]��1Q�XR�d��o�_�7���Ǘ
φoGrKg(���_Y�i9X��z�ڗ�֊%�`v`����1�͆���ɬ
$�/�/��Ա�1�-�]��Z���.*�'�\��x 2�Z�#��l�͘`�3�bJ]U�@���;��S�`�A���76��}ZxTLrl"�[��qxmN��%G*[6�S���o��Yϵ�'J�"�{vm������+�c=1�6ݍ�\h��]�tx��5z�о�)�[ �XG�S<���y���ΗZ�y0�*�����o��%l��d����ў�fty�n<ׄ9����)ܨ��v���ur��H�.���G�eEf��Zߺ��˗Ь�[Ƿ���/qߡ��Y�k#��	6�=�WZ��MR��w^qn:ه�5�+J�/�k.��[��9��o[X#��
�g&�qsR<�.gVov�y�����[u1�8���һ6I�����%ȦPd�lPC[�}�}%#zW�Ȏsϡۺ��o`���u��p�j���(U�F@E���Ⱥo6본n�J�1Ď��mǘ�������H
�'� ��,���[v�jW寲�љ9Ɩ��H�s�c�vs��yF��mp�,��kwYם���MT���7X�jr��(�;}3ؘQ�L�)a~E�\�+uu[z����T:�k1>՝��/ݾzi\�wj�IZ톴���O�u�.4�	ӧ(����X`�m�6�yZF󝭜U_m7:
�%�{ܒ�E��-uɰw�*����9�^b,_r3��d�^�Y�,�,��@����B���h�k�17Rn�C�J��8�Vk�u������j.ڝ�ʦ.Sg�$���=T�gDr�f�Iѹ�/���/�\&e�ۆTGy�]�f�f:��xs�sx:���ˮ�l�[�L2��u<��Ymq����Y��y��7lۭz+"�qZ�T��辨E:��Y=���z�m��1xZ���}������/r�@��'�JYۼ��JV�=)T��D�5�tz�Aɠ�5m�5���NR�<b(`�D�\i:.]3���pU�w��hx���%}ǲ2���a�͒�k7��f�8�ǉ�gox��w$ n�ۮ����S��G�YW��s��g|��-�+o�8u<<�w8�^�L넩����}�ؽg�=�)ɮ��U�O3�<��K幱fg*�a��(���.� -�]�̽��_f h�D
��}{�v� �mf��9�Ǆ�I93y�,��	��Ax<r�;���t�U�'���h���h˥z�..R0��r�{��G�Y.w]�4�E��q�O�WƇY�iڝMuwpq䬮f��t�s��n��ט(�Y�',����iވ��@�ʼ��� bA7f�#]�N#���Z�\g���"��7�����L�XWj3���zgv���	�sy�yh��}H`�R��x��E{Ɣ�T�+�or�I.IrJ��\�.Z�JS��S��r)Id�S{�V�{��C�q�Ý�z���g��\/�+Y���	�&�r���`���ɥɌ��f��i�T��0�)����* ON��Ԧ��eјy��&�<�9�@����wr�� �rv��$Z6�s�j�ct���a|���Gps��}��>�i5jh+8���u5��*��n�������\)���r2�����n�f���ݓe�P�kTT�#�j��΄.�X��Y!��ŋ�����[E�<�*��0U�Y���#:��q�:��r���c��]Ls��;Q%-g3�JU��:���/jW��yƥ���~(�+&���(+�i1����A��C������?�f���-抃�=ʤ���#��|%[C�n�8��86��:�$��6.�9��Պ�A���Vmq�Q�z]�-��}���eѥ4�o�J�&F�]�]}���ۙ'Wk��@+��e�nM1V�T����s�gT�ڶ�6�9�MF��p�>\K5j���fN�X[�����Bt؝M�MՈ�]ʭ��1��2%�}a�-�.��eL�U��\��U.䩰-���f��a![3��B����]lj���|�l�n�6#��<7rdϳ0�̎�)h]3���,x"[a\i�kpaŁ���.��
�ܘ
n��Ӯ�#=�t�+��پ���QF�A�W������o�W:�r[xZ���q�@9F,@�Q�꜃T�c��o�x�\D�x�^�Y����uܧBmj��յ�#гv��޵�o�x�t�u|5dB�4f������d�����F����r7�]���ג)�p��F\՚9���9K��2�'�P^�>Y}�.+�v2]E�%����Ep���uj�7��4�!s�T!/*.�ax�礂����8����uȵ�,1�9^�V�8�Wc�N�%�/�%C�׼xA�P�%e�I��(�=Y�Nȵ�.�`2����:�V�H'�m�#c��7`dSS��XՅ�*0��L0�.qޔ�\���h��:u�}�MWU�-���7y��V뒰��^}Ζ)J�8�a�FH����p�]\06�24Ucqs�	wRq��I�Ϭ ӻ���9v��چTi^��y�e��S2��
@3g,�pu�Ę�K��yݴ��ˣ���n���U�gq݈�ȡg�LhF^��;���n�+�x��Sq��-oR���]��+�Ǒ��ꗱ`lGs�LL�p,ٻNr��f�e�u�<��q:]���f�N�¨�򣚡���z��Պs�kO	ah�+��5a�OQra/�;�,�Ί��.���z�'�ut��u��~��#T��������t����A�v��m.�����E���h�djyf_>!��5,����V��ͥA��'Q��ˁ*�vY��+51��v6J�P��A���\ ���S��\p&�x�j¦i�7eo.��u+�[�[��Y��v(�0DZO4�� B���͡t�U �V�O�gPe6�Q�<�M�k�I�ttV��娈��u���tbua,���IVm�=�qν��;ۤ4Q@��#ҍ���Γ8𳁝���d ��э�r7�Gn�ʑ�����nқ�{�	�`Z�&�6�����k�R�ᴺųn��N�8�ʻ���70��,k����ҏf�E��	ZLEU���a�L"�1���x�Ju\�L�����$�2.�[�̅3b�/۽��Ò8>`'�SƶXX�Q�� �0�tyއ���Ȫ[��C�O_nFX��׷�>�]ð�q�Tp��`ðe�j7�MWK]�\��٭n=h����R���t�2�-`�s�μ�;�4E--��M�:n�_?�P8ky�n�ߑ_K�5t�����^�c��?��!	�=�y���gr'��G�q�%�WnM5�1����"���,��Ou�(L�ڒU��U��Ҋ��7v��w���ޢ��XU�\�ل�F�G�Ѻ��J�Wsi��+V`=ݶ�
�Ǿ=>r�X��;�t�E,��GxmƧk��K�Z�R�ͬzU�1�g�"|�^�3;B!.(TЗe:y��*�D,�G�<�c��b4�D] H��w%�aiQ�v��Qm6l�]�u��e��%�}�[Dq�)#BC(LC''�.C�J3�
ч
[� �m�v�|�@rνN���qB�nW#je�9Յ��G �2mز�b���٣��6�7�]]�es�pМ��!0uo��V�ݻ��b��]��eEk�5�a�6p�s*�8�
x+z꜍,�۩ٌ;#�\��V����s�=���ZOc鴨��޺��Q�/��=���[�V�oA7$�RU��=s���2��R�L��1�Q�L�.�v�3k�$�47p�)C��!���VFqu�J��gk�Ԇ-���f8���t��N׍}t�9���f�aixn��	6���񝖟�+�v���jO�Q��+"�!Qw�"���!5��^
�і���+&m��odB����pF_+�ec^��t�v�0V�Ū�����;)B���+*n���s�����s���f,\|d�󥡅�nl��湳;i��>��x�����Β$�F���Z]u�����u�A����� ������7�}*w���"Y�A7kHqD��H �>�-� ��E���U��H3VmX��+i%pH�V�p\�$����m݀�h�)�tM"_�b�y/�Rb��NW&6��ayM��)�L��)3�u?�T����oeYJ��S�r�G�)<e���tUe��n�ٺ�t�=�l�Y�b=��黳A�4q]R���M9]�{3���yu�FfU�K�[na 9�",�)��M��Vv��T{�Qr���h�S'j��pNۺ�7��F�q�O/o����N!{LZ�e�(� E(��4�G[�W]�\���wvT�ހ�Զ��������/s%��rWi�XɃ�r,\��ٙS��na��~W�inK۩��Zp�)��;�w�c�m�d���2��Z�i��\ӥ���F��p}F�1��$�S�h�ΧԦ^�*m�.�]*�!�2�s�@�&W.d�o"�b�qQ��hV8	���i-����|�fs�X�=����G�����͠�z����<
b�z�e��⭗�F�r�2�k�)SH��0º�i+6J��۝�YKP#ohk ��e�uP�\�}��R�����wU�re�_t �ufb�%n�!�O5I>�CL�O�'R�������������B)�t��-F.�$�\��Hd�|u�	�k��WnTf�C��Qk{Ugd�qv�c5w�&R��X��{������QX�P��O�%�9E�9P�C{�Kz�n]`��Q�݉@n�\z�23-d"�S�uu��Ҫ�,�v3A���Uǻefb���K�UF�2{���P@�{(�KL�guSd�,��+x����Kj�Wv�J�NZ�ZŴ*X�ٛ�j�$�#{�]k[r6dVQ����A�����&��u�Ʊ�U��V�t���h"wf
|@cgC��R(0��v�Z������[a�ь�i�����;-��D�rUfU�=�|{ ��^���7�;��aF.�V�/3�V��{�K����!��M-�m�o�f�BȰ[ၡo����qF}��E���۩l*l^L��F�fQn��Neɓ������������)���\V�3ֳ�-%p%u�Z�<�di�Ԑ�Z��
DsսPS��]�����Ѣg*w�7]�X��9�%�:dc^ʕ���t�s�RM���\�o�+r��@������v�{�Y8Ƀ����-�p�eԪ"��P��Q!���r�<�Q(qb��>}��e���9�xZz��ϚQ�Of�x�(ÈuF嚥yOn�X�o�+E���r�?f�	5v^9v�]�qR���TD�!��+��,��,Pwo������e8�mlcC�X����#y� �.٩����0�%Z�����L�Nd�l6�]nY�S�u�ge�A�n�Xr��m�6�s�ͣ֎	&�i�y1��v[�_<W��"��6{;v	��^��kN[KI��YX�5x�2���t(t�4	�g��<�v��ꦑSEj�=�P�)V��ps��;(
�\7�JѩʬYfdnWK�K�f&��m��ʙ�zWe�Q�;'M���F���rvf����)�!7)��V+�PĮX�}��b�ӥ�wVD�#[V�rx��{hѩ;� \D���X�V�9�o`���N���ۂ���ocۨ�{�c]�w3��4�zs9vd
:���9h�d�����D9�Ц�ofأ�_���|�s�">灛�$l�����.d،;Kl���쾋l"��Dt����g^d�)ǔS�������m���(\�k�� �P�G���h�e�+j+U��z%bۧEȄ�V5��OA ��"��A;t[���T�/]�H�u�g*?3�j��E�9�B�E��@��'�ƎnpXq��]W-MF�)Z����k�oq�[��+�o>�q���h�>�E���OF'[E;���r�5ms8�#�0S��/�3樋[Q�Y�bp��;���.}��
�%��
��:oayB�D�uL2eH�]�n�e������[�*K�q�r�j�R��:%r����̺�X�5:��M�+��FW
��ѷyck�p��ڰ݄���P�/�ʥ�T��*Yb�l�=�� ��f�eٔ���B����{�ͧ���ݚ�1݅H\��i��6����74��j���!Z�ÖD���Wx/����U��X�?,�2�j��jW,�p�����V��V�^fU�[˂o�a��K�uї�8�����z���u��m���)�@7J�ƐW�D���iF��:��]]j]_+�5�`��N�W�ć�oP�>i��d���ϐ�i�y�b=M�CW]{$��P^�8NT�.��|"�:ͭ�8�ǭ�8h�Wk���mp�G$ |��rT;����=i�2�+Ǭ��յzY]R�U�j�d�z��ֺ��2Zx,ڥ�C��fd�S���K��v��ޫBE�t�]w��#��]�>�����Z�����V2k7:�Φvu��<��֍+�o]������g;v��.�W^:H�O�Y�S�F|뮴��$[3��/�D"�L���Z=�2���7���b*p�t��Ɩ�S9.U��ǆս�\��kj��}U��̘iLT��J)�y����Vd������t-�N�`��RY��x�a�Ը3����nT��ͻP55��O�ͮ�H��6N{�]B%�tސ��ہe��4�r�w�t���K���#7�ɉ;e�ӻv�T�˨�p�b�\�&g�☫oBF���`�sŚo�N!�2�	<�m@�4���c@�O@=�,MՐ�ي�U�Y	ƾx�1\��1�ι�,�Bndu�&�PѦ��@�Gv���h���w;�)�W��\�.��rV����\��zj�'m�m��N
4_]����J��*5ԭ3v��.3�A=��;����V
��/]cڝw��Z�X�zl6DVK���"�+'i�iU���Q�s7Y9�d�G��@���^^+�Q��V
�+zZ�v�Y˫uҀf؝�5M�o��N�e�r�Q��E��OeΊ����~��5�����Y�"8>!���3��L4�ټ�cg�jϥ�uϏL6�7e����}N=ݨ�[
uѝO����*�t�墮H��𣦶����t���Tm��W[��ZF
r�����(0��]*�KK�<dݨ/�5�/������;��ui��,��:�	f���줧�eZ��8��p5n� �6�[���t��*m��n��k�m���$�١w\]�5�A3/VG��tyf����㝹q�X�R8���(W̓mޗK��E1 (�s|�3�v�������Ko3"�1���h�S�"��.�M���
�Q,��V�����KG+-5�@�;5��Z��]n냍Wf��)pV��'Yo3�__$��Z�Al�:t*����A��zc�&�p�5�t%J�jb�/T!�P�J��J�"|��<ƘivvQc���ܺ�{�v�U���&�Ec\0�����i��[)���4��,��4\��^-��)'
�N���''p�7V�C�)����!���T�nմ�)eDW
�]xX�oz���rz#i�a
�:�|���k�6,���1KzU5�\��Hc�@��fB��(�#GRK�T�������Rܩ�Ȏ_��������':�?vƷ���4o:1�����f�Ǻy�ګ'4�'��f$��["n��n�ҦvW�Wc8�eѭ&o���s���N�ZAs�4��3{2�՗�`��-�UB4�8��́��kx�rjk���}����.�z�u�LPu����# ΣK�օv��w3vTQ�����;6<yf�s�6���SK]�oye,[�wc�b̚΍�|���5�I���*4�^�
\��������|T�/��VX�$�#:��x7��x�z�W9�U�1���6�w*�@���I0�f��czf'�9xq\��9wP�=J�H5�:UEë�#�:�5n-�/2�##/���)MX�G3Cg�1>'�J�6nRT��P��ڟr�;n.�����*���B]m�5B��P��y��=J�8�4m-�T�Ѷ��+ƫ{2�.g�_m�}�Y䚫����s��P��r�Yb��U���XN�ٙ�(���Ս��`ɱ���r�q��n�@�K�����������]c.�Yf���Ɯ�U׿`�9@��Uï2��-�ϯ��
�N8U�i�v�Z)_ᛸ�:�`�
P$�5��H���v�#9�oC���Fʹ��vz均ZY�^��p/����\	E��ґ�,��Pg֕���q�Z�����9W��Ui��5Щ�L�w8V��vk�&��%,q��{5WWO�xEdF��)����+Ǎ�YHA���n����dJ]D�V��S�"��P����c�*+w_f1MӖv��+k)nc�Yn`�^Ô:=-��]8_(���U��N�!Z�YorP��2���F�V(ְVZ��B�'fB%p��c|���֊��t���n*{�JoK}4�b�aΤe��t�c�:��eq�&�qӈB��%=�����wAi���EgZV�,`���r�+	�@L�H`� ��}o�ۼtWdk�����A/���<hY�ZFgq��� t�7c�s�e:�iH.(���N�7���P��A*�=C�푼�����*�sb]�B:��
(�كo
 ����f%Ԟ�ۢ�òg�;cr��t����N����S��l��[���V_����<�k%���29�Q�f��P-���r�8�.*�����Z�t��Ut��v�5-��Q���;:�O��,�P�7����vj�֤��1i�.ӻ�ٽ����m��'�b��&�!3��y�g.�],ɵ���v��6�5��{8f�4\vg�Z��"�n<�zh�E7D�Y�@5��)�rvsz�MP�&�����m۳��;u��L����4;������9z�n�h9�umNXh�P��Z�+��Z�q��;Q2��Z����Ju���/��/v�Va���z�����$�lԞ[��$��
�Ďh�B����llH�&��E
YێR���L�|ҧtp�_'�\+NKa�ZZ�w�\�6�8m])5N�M/���riE��v�lDk�(=RJ��K&�r3�9eq�-���] rK]�(����\�'c�qE�U�$:5v�g�P�J�T���t�xYH�

Hh��Ȥr������=���pM�9����Z�˻����t�d��s�{��9�X3����m�_�\�g~v����Q`#��lgl�(�*���Q1��Dd��E�(�[m
�kd�X\Lb�*��ʹTb0::�+b��V
������X,PY@U5�&"�8�ɨ�I�\�EU�$���
�PP���h���U�K�fU���j��Ƞ;J��AV��r�cA`�c@mXz��c"�*� T1�����Ջ �REmb֌+q���X�v�Ķ����6�b��0��.ڂ�X,daEH��v�ژ���X1J�������ȰH��� )1�R(jU@X�1d�H��j-Gssd(�P��"�B
���=r��!�a��ը����=FZ���;�rheE��&%�O�g+V��M���F�{-IB���g��'���5��%'s���R�f������3ي���F�*����j�YV��)�4�E,�"�����i��:2//�h���@���N0k��K��y^dPo+V>�1�dDE]�FXT����c�I��aR6�b��.i@���쀎��Z�Dh���U�c�\&�	"��>����"��<��;KA�|�z$�V+C���x�v�'Tg�c�B���wJ�o\{i�R��[����d��0P	�8��ns|껥��*����s���1����ymJ�
�~,񔮙�^�d3�_H��[.E��ȱ�'��NQ�II���m'�NVGLD��y�^�NQ#O �^��j���e��J��{�1����j\>���1�.�u�RwpIʙĪq�Y�,b�E�F�9r�!ng����/j���D�(�x�}���n���^Ah� a�py/�Wi��]"ĩ�s�k�e�F����7��Rȫ�A�L7���7���x�T���ʬ�:�V�pO�X�0��캅��"���"�n�&r��"`V�"(�"�{�č�(��6�ĥg.����d��T�-��*T,�[*K[u�U��ar�(��Vtr�]�ԦR��x���[�3��s,�K�^ 9�ܜ\sR��?Qp�������`�U&�zez�G΢�$�]�D�t}nE��(8 �+�EM����CM�X�8��W�{��K �X�i��.�!�IU�NY�)߉L�^�@a-yhB���c�4�ǽ��&�n����L�VED�0��k��,��C%)g$ĸf�5�q�Hgg&�Z���9Ycc)�X��OO���4p�Ÿ��N��T�h$e�+��0�3/��8��o�[�S������6h{�R;6pT95t�q�r� N�"}��V�%׸/����-��9vgf�o6c ��ר�v���Cx����[����"����0}�. Le=p�:������\�!�Ç���0`�#0��Af��|���5�OqW �A�k=�އ�UL�մP��(P����ǥ\�s��eK8}�bd��#LӪù)�7�(�:���c�h=׮j�:O��,�UXo^R=��\;������0_@�w�v,�뢦{1WY�C=�=��z>f�(�����y�ˈ�oO�R�Sn7���q�~�^�I\��r�c�V7�z�Wiv($��3�*��,䣎�Zy����9��]r>��5����\��Oc*��#�&�-<8�aR��*�/Wbr���}��&�y����C,1��t��_�x��+ޢ���*Mi����enYݘƞ�1�Rs��3o��p����5�.R�q�kjo>1~�,����7��n��F*��E	�����ow]�����U'�Ct4�
B9B�hu̮0+�ڛ��L���D*���np�6��Uj�L-+6�Y~�'��3�{�W^̣� \����gd7�O>��nE>�ES�j>�[�g�HӋ$"�s�&�>5�d�H������+��pc�@����m��IDU����s(��}>�Vu2�M1�b�^��v"���؀\YbI���9�Ucr�cB�0@���G�����6.�@(F�2�ay34��`F��xfх��K�l��ȹ`+�;x2���r��!�,�����r3E��8}�嘾ڱ����r*�_��#pþ��f�o�3���1��̄h����Q������U�݋-��;;x�3�dH3q��5fy�Mp��V�|����@%}N����'�f�S"�pO��_0�����#eހ��׃;J�>A`�o��4�ܔk�sE�}2�5ff�8U���$ldu3��T{��Zjt��K+�Zun鴮wb9lf�L�ne���c���*=.	:�Z���JE���v�_�g�
�9���h�k�NJ�1t�j̀�q��ge]�l��^W8���k.���*��S�%��"�X]'oN[���z:��~nI�>�f��J�1eH��j �Yh_�¯�
�X��A~k�6윌n!����A�1a��1ꕊ�4:=g\(�W/!��dVB>1�b��-�u�u񝞤 ���N�<��Ne:�rU��D ]�t ozQ��V������]�MΘ�"36�G)g�d�6�(�Z`�i��OΫMߡ`��sh@���%��/y�|�V	�y��S];G��v����J�C�ǋ�=ぃT�vZ"�	å3�1�w^�9��b팭w1\��֥�
�;���ݛ��D%,9u������K��;[;�8u���Z,^V�o�-�~P�k�^� �W�h���w=0�@����^%q�����r���or��a������>��>��DgD��n��ϼ9�G:�S/�tbyC5H����Ʀx�Hf%G��C��<0(�_H;A������)�mO^�����u7��@�/���U�Q��l7+��GpٺP˰GfR���ܗzP�kr��LZ�AJ� �����1ۭY��!vi\��ٰ�bn�a�y�N��;ؼjy����#�/�\��sQ]�֗]<����}"��Ǘ�K�����ש+3N��@->*˨�Z�.Ս':Z�`��Sh0�9�>�=4{6�ſ��׌�6�;%�R�S��Ś�͞���@�JF|���t�=��T�.�-�T3L���DU~��_0n�A��w��K�@Kf|�ˮ�YE���4�n��+�5N^fE�8M��ɩքE�D��Ά�A��(�xxNה��sV9HOD�ړ �՜5r��閭υ�ּ�:��kb%&�4n��89�5P�/Iw2]��9�D�A���y@]s��B���X����+l�o3&�.N*�����W5���U�,wtD���,d��'ۍ
jF���~���B(�MF]i�a���q�߹���oN���G�h7]v=ٝB�	�3Y�`e��E���#���:1 �B�a�ݱ���׻7�xS�g�)OJ�4�"�b�ʻ�5^��\�\qk]�JyS�o�׻6)��	B���X
V�wݮ�ݱ��J|#�xô	���B6W^��Q�W�]C=Mn�{}�j����^^�~��Z�=ǺB��KMW�X�+��
����ݤ=�z_TW9Ȇ�K�¯V*���Wݜk'|n���wKVtWM�43~��%}�^���5;�j��%1yP-�Fo�6�o5#���kX�Z`�
;�5���')�Q�j.*��yu���t����7�
7����|�=��R���rՈM�[
���7���;:�����f��ܥ��2�v�kkZܬ�\t��t�:$��,�,Z��u�oН���L��>�;J]�����o�zC���"��+�-Miŕ��DLZ�'u;j�]��_�9�1r�@��&e�:v��e�T�^��-���/F�wb�W�9�-P�=�p�}�Ԟ��lʓ*��ޅo��U��s3r9���<���دh�'��3���e��-��)��kBxɑU��&��1�'h��ri��jo.��4Db=���L�P�u��"p���I�y�l{�J��R{����eg�WS��}B��e��o�v{���YJ��}��P�@��V�-��Β]�)VK����S�����&�q�9ݏ[���\��D��Y&	�ѭ�	޼�ju�ξ��6Hj���{�=�kT*���oi�.���z4Ӓ�멹F�����+r�源������Σ���
V�}ڍ7��a�1���ݱ*��-׻�	u�o!;��gyn�[ѵ:�St;��
�>y�:�>��h��y�m���>*	�Y�-l�U=�:1Y��f�Su�v���n��ݛ�=3��+���}�3ޒ�3�N��i�yr��X���f��W�[��V��̻��@�z8�Q.�����<Q�W�5�J��䭟Rfo�6�s���^�y�sV�y�5�I�7��<�����ة�9�:c�x�U�oiJ�|&���w��%��ٜǬ_Be&!�'Ǘ`�핔.�dW�|yJ���]Ө��ǖI�[�&�k��\���|��<'���YU�u�������YmcTr���l�[��Y���M񐴇+���P3}�=yV%�k��/E��:�r�J��[�9*s-LL�̾St����>��9�����mw�B�����ţae�'����ޛ�<<,��o�&��A��*�)�ú�9�����S�Q������v���{�h�-�}rv:�yjd�QԧB
\6��٫!.�ɹzc�<el�B]#�{Է�j�B�֠��:^��e�OlS�+�,�z!��2�#hm��Z�kj\�О8������2rg(f�[�ɕq��H�uf���,a�;�en��S��nq�.9RF@Re��YE��ɥ�B�H���D9�ҝZ�r��[��B2�/�	�2Ѹ89�1�7����M~'�Z!ަ���d�۝��������:ѻ�|Lr��g7C��� ��1�k�7"�T�lpܷ:��F0o��smǱMd�쌛:�=�1��1s�1�s�F��^�ߓ�õ��,v���]mI����Ϸe�W0Zl���v;@�B�3��yJ��ީ���Q&VC��ΎG;���[�.�<�����f¥WCpRf@�Hнw�/�z�aX�Y��|���7[֡�[ove��!(Yn]hp�E����v��C���g]DDT-�X�b%h5��n�]��7rb�&毜�Ն\�֟7xK�.�)�de\��oR2�rf^c��rW��7Cz�sGU��2�}�W�k(���$�ЩU=����n�d	�mm��g1lt���ݮr]W.�;ɾ�C.���VF���+/�K���V<��^���ÐR�+��Xr��ˬ�Z���Nⲡc�[6�-�%���O7�����C�6Bg���{�n������y�F1�;�E�|������3T�sw/�)3�2-��=�I�����ˉ�%��p���l,�K+i������?{>�7޹9��Z�[����Kۀ���u�a�"�le�Ok�-H�9ڼ��h+��.�)ؠ�}L��/��ҫ�,BW�-�
L�Ι�}2�3�}"��\8�1�
������|�"�a���H.y�[2�ˡ�k(�v��ɴ��!7��w#�Yû{��q�,K�h�Mĩ�t�;�:��yҮIC�[����נ����i3
;�j�j[i6h4n�Xh�"$�l�����щ���P��/ʍ�]7Yr�e��.G�3�����7b��W�C)+�x�h��u����$���}ݱ�7�cj��ұC79��b�S�<�P% ��*u�]�tN^>Z�['	���P��9+���i�ޤ�N����<L���M�O�����][�C��Ofm I�������R=9�=��r{2n��&-���m7o��T!{�
ju�䚺W��l�9}78Ӓ�q�5v7��-�@k����.6s^�r��&F���ظ��z�K����Y|ۛ�[�Z��׻7�xg�>��zr�*UB�h3�J�F	��/9�Y�_�z�sSʞ^���̞��^C��v\*�W��TPǁU������<����+淖�:��j���@�gq^� Ȯ�9w+��u�80=�~^Ps�q�iڱ�U�<�����O7�r�͎���c��ؓ�o�����t�۹��:���k3U[<
%�]�,<��wϵ����i\��#z���a���,Z�+i�ոn�]�g�:�!�����Φ�T
mzC�,:M-��U�V�^
L�8Z��UY)�����䩋Z��)�	�t3�ѐ<G�G��6 ���Iyg?Q��B�X{��j�w��e7w3WE�^�"U���{}�_�R�i��vľ3w��1c�������wO ���eپ��jʩ�;
�ض�5w��5HΫ��^�yʢ]�C����v�;Mt�|;u]�5�S���0s�b^ŊI��V�glίL�p����D7����y]vg
iEt0�ޕ�ې);�B�����Ȉێ
Y�˗�k����.&��i�`վӺ�F`�=w�w}\��M"�e26�e�;��`,�)��)�-���v���K��!Ȩ+N�5tt�)!�̭�a�s6.�hmlD���*��;��@�ʂ݀����s6*�߬m���e�R�3U�H�]s�l�2��*I
��f��u�}�WG���ۍr)��L�wc�ӨS��Z����l�GP��^G�Z޹W�9�X*&F����Q�s�9�7K���
[����]�ls���u�4�Z�ΫSDU���\�s�����A�/V~�t�N�܊�L�s\��-U�R5ƻ(ɽ��^a�*�ol-��D�ͼ��"1��bPneme�ë�@7�7u���]����3Z�Y⒊蹫�e�"��T�^9���V��zRj�ia�1� l��D���-)�h��+
u.����H�H��đ�]n[�H��܄�]ȍ�>�1����!������Kn�Sg�
���X���(�n�X��+�;��[�\��U{R�/R�A}�Ȩ8��uj=وî]�<�����i/��>x��yRx��)�Wj+����/����<�m�1�)7��P �.
@<��r��������q�Z�i�֣��3feQ��)�N��Xw C��czG�"����Z�\ȡ}6�iѨ[�{^���F��
S/�]�קw+��#��q��ڼ=W�T�Y��f���qn�=)!Ih�x��-�N��nYpQ�s)�!F�R�(o
#���|��c��#�in�c�U�B�L��ZTg����>qW
6�o_��Kˎ�#o����}�q�{5�6��a!	}���Glln�鷜��Wl�SJU}V̅$����;l��oQ�.�`��(�}2���l�wҘ}����˺���u��s�2�usm��Gg�w����U:�8:}��
�ԕ/~V����B���Ym<.Q
��m�.a�n��edD~�Y����l9���	tw,1�9ϝ�_8���!k���x���Е���uHB���$�Wt<)�.� ��ó��s���H�;eO��s��v��j�:?d����t��ح�����Mz�{�h�[c��Nu�t󒸚�l����,���5f��N��9�\�9�}G�v����]G�n�^�IqNU"]��P�VM)ޘ�G"/g=�A�PH �/�	���Z��p#A�G�s=:�m�ys{;%΁���G˺t@�9n��=��z�
�X�e�T�e�5�y~�>�l{�I bV((OVjV
#"�1��dPDR**c*([`�v�1���X��b1TP��;IX(C-�ʊ�
M�"ȲD˹q�1Y��+���I��bLk+(��A@X���*�@���@Y"�

$Qˌ&$�SPRL`��J�Q�H�-�3Xk����VB�BT�$̱a�IY%d��Y"��cY"[	P��`c0�
E���Y�R�16Ƞ��e`"VA`�&��*�TA�I�k5��
ʚ�2E�mK��k+�
$��+ Tr��*+cU�ˌm���w1�%EP�fYC���ܠ5aX����Oh?�D^��-5��0��K�Α��A��q⾫|�ϰ:�4��缚�ZeA�ͩv��k6ik{u.��{y&l�5я�GJ���g;}�\�z}����	l�Re>����]Wо��3��	��دh��({��bn'e��-�h���s���R�Z���>r�j���@蝣ϳb~ew��O����/P_�VK�?N��&-OC�U��f����Y�xfה��o7+��u'�~~��WY�I�f�8y��<1+�-]���"CC6�psv��T�K'dMi0z����Nzns#�
��t�kF�z9���kL�}6�l���X>�d����F6�=�Ox�Z,.�L^>��r��v���[���69�k��γq��̤��c�V]5J�[��(`�L�Q�U��ޫz�ft���5����n�D��/�ٻ��Z���F�9m6@�̋�Zw\�)士ww��OS�G{!�����a(U�ʴ_����96��3�Ηv������ߛ���P$����A��Y�A�w���*ĕm��Od�7z�^o]���ړ� �������N�ȮR�A����k�O�ڻ9?a�]����ٙK��`��qu�2�6��n�N7dQ{Jm�}A�_t��nqQ���}�e*�X�A�[�כ��b��-�z�P�����~�+��曆w�Jc��7r�v�_T����+J���0-#��6��
�I��=*.�f��5�p�ԧ�N��	�v����g��o�1^_r(\kМ_(��{1�E�b�涱\�څ�@�<�9�v]<�~YnjQ���I�zrtl�$xϪ_FZ��,Z�㊳1Ї�!��e�rT	8T3����ZC�{� 1-�&]{���o�n�dUڟ[:�`��÷W��˕#:�Q�;	��9[fT�t�Y^-�lJ�۵"�ۘɋ{#��VCjn���NH��0�#��i��e0`s�c�n(;yr�m����\�9�=;·�[q7Y�K�̙�{[1>	6k���ĪQc��u]@���[�n�[<��Me�,^PO��C)��.F�bB���{�6'3'*���TrE��V���HG����q!�/��)u���S.�����.�jЛ�J�7̼<��ëiڼJe+{+_`#YNNg[�ޱG�V۹�&��[�Q�׆�\��u�����#��47s��,<Pc^�S�[9ٰb��Z��"��u'9wun�.p�ˎ��p�7ض�Y��Ɔ�qW��,X�::�*S�7�§Zߺ������T�.�	1FOk���t����f��*Y�0��Oo6d����x��Qս��,�b�D��1�V��rV'�
op��)��<����P����JTݎ��m�ٱMAJ�Z,۱խ<�19
��j����dAa�~Ī��[��<��tSa���P�ܬ薕(�hU$su�v�^\�L�u�ĳ5o���;�><e����#[��v�F�j���J�-���P몯����S��=�󛅒�
M^]8�î��s�tȎ]��P�j}[Mߧ�hB���A"�	$���z�3;=���I�
��Bd9Xtȩ[`:{V-H�;�ڃ(-�̬j!�.�B+9!�$���@�l�0�gL��їT�+�q���Z'�u�
$��Wυ���C��*��[W��;K�u���~G�;�oP��c�y�=�(ޓ��sS��Ww������O�2m�&5�ɛ�y����?_wk�X_HK$�\ev�>���u�k/T�jڷ[�J�6����	I��L���f�y��N��N�lPI�ٕ&] xV�p�K8�q��k���eܙ��+(�����a�ҙm�>Mĩ�f�WH��/�b�G;��j�(lOH�c����Wd׮��Ky��؉&�����d�A����5T���wr�x��=yn��z��\���X�L��m�D�Wtt��ϋ��_��d�D�؆��&�:X��J7���b͝�tk�A��T(����yb�an����2���h�M9�r�����&So%
U��A�`���jg#�biM��m���י<�2}X�VժUh�w�s�]>42�޷yP1W/Z9��ܗ)w�[�a�ݙ|Gq�n�jM^IP�@{�b�{ؖl���PaO��"�#iW>\���:Ƶ�vB�1��X˴�,�X�<��L�{�B�s�!q�iڼJ�׫��ڸ��.r9�6�V`��m��,N�{u��w�W�e*��E�(����K:��bn3ԩ^Y@݂3��g��̠G2��蝥���4�ު|��C�mG�G��sm��i���gN;�;Xٽ�"�k���:����{H���J�k�(e��J�n�p\Vmfj�a�c��;`��=�E���=��Z��{~6�>�;�/�9����o�͍azGJâK}��P�j�]X��6�$�=��ʊ���'t;\�Φ�����2��9��x�0����ͷ�ج�,;+���jm璦!�����̺V0o��z��m�.{~��qm����ũ�*�μ�[�����;�l��L+�ڡh���n���7�o�v�Sȫ�7��0̌n'e����u��GT�K�r�;}�n|�zr:�	����4�n�˦�D@���[�6xU��yБP�Fnqa�pgX1�!��AA��[��{u("�b��S˻w���uN.��bRl�fdߟ����a6k:�.�M�(OGڇ'Ov��q�=�(���n���w�v�:5��Q��6O���^��b�����'�AQ�^J��ǉ��|�d��ի��L#}]Վ�,�mPv�H��Ԡ���[�峠�rvQ��z��+��Z2�MBV�Q�,�Ÿ6�[�u���<s����B�2R��7--�e>���m��¢ޥ'N�K��s?�ro�V%���^�R9Mֻ[aj�a��͎zm�ZŧQ��UF����D�ئ[V�����]!"�3Y�G)U���m��f��V$d=p�]�׼�WW��X��:�e{V��CpRfE�F�;�kJ�t\	Y7X�)g%�]�F�ީ�M�{�\;�*yu��k=�}7ӽ�k���;���2��l�mo.Q������e��[c!Z��1˸�����71����5ӱ����T�_y�W6��=#�y3�O>�6D��퓽6�F*��Z'�e��,���	�v��o�/�y�+Hr}ڇ�B�]��6_l���i#�~[��g:��h�j�]M�	��bp& n��o��sGh7��]�石h���jK�W���󔕃�v;��<Y�����v�	H�ReP�oh~Ց����᝕v�9d�����B�+�����}۽5�"	�i�*��3���v�D�q,�B��T����g��xG��7����h�=0�^����u�2����9Ҙᬜ���A� �L_hNfSv��t��&V���� �r�v�U�1.JJB�v���0c��y��e�eI�@��7=4�\���{�2��]=�w���[�fP>�BC♠��2�C#4o..��@o���^�ӇN��1M�Uvy7��~��JM�h���s��p�'���n׊!���� ZW��v~N��?�X�֌J���ʜ�f�������b�Qu$��C�3�=����\�7�
�*{����u9^ �n������G�3%��_D`�{���P�u]!"�3����K�P�ۭ��QУw�a'i�̞�������mXT��v6�9[.pͫ��9�s}�MEƖ��KG*n�Cζ����H��e�u���kv+imK�	�Ԛ�������c��-��C��/���rR�*�Gnξ��]�Zr�k�#;q_�=7��ܶ���'u��� %���z �I��)]l���<1QF�!O0���x0��Mn�)�i˦wQ��鮰{���2��ų8�
5ʭmsr�J��1�Y$�(
���w%/���wf��	��X7�c^Ӌa�Y ���;�� ���!<��5:;�a
�X�<��,��"_�
��}.��9�~ٷ�Y]崟j��˾�����t*����B��Y��<ei��{lJ����9S��E�뙭��SN���ғK�sc�쩥����	|d�r2*V�Xt���S\q0�rn�C��<�E�\�ވo����	l�ReW3�EK�ɕq,aI���ܵF]�r����נ�Ct�)'�a��L�&se:��2�֬2�].�-d�K&�v�^_=�1��b�qLך9Bn"y�"in<�E��l���Bv������B�O�.��ّ���JM�����:��Ozy�ط�ܱ���p����/҅����[�k�nanK��h�{҂�����o3&��cض"Z��i�eV�VS^��w�Ry�K���Z3����gk�c�an���7�_D`�{���!�ΟZ���`�(�̥^c��lЦګƗT��)O*��6s���P���{�>�i-�3#-�q1U9[����=ˤ�C��+�,Z�#�v�:-��Ņ�C��V���{-��0�uG\W^���5��%3,iy�v)F�κ�-,�
O^mvs	Iݺ�����&� +H��ܢ��ŝM�{�k�]�ixL[�}u��3���K���Ƕ:}I���w�r�lkz����SPvG_7=��M��9z58�QLGuh�)Yt;=I���W\Ԏ[��<��2�F�9ó��jMNo]ˮ��B�-�nVP�����iڿbUB�C]qu�̹{��f�9{����cX·�"�B�7����C��]M��O\��o�+��|ɼ��sY��|�lk�zGHXtH-�aeX�r�v�f��OB����.5۸n�ݮEgSr�`p��a�")nc���R"k6�'�K��ji�U�Y��Y�s�J��-dL�L�*NqU	��8*�¬�9�GNGd[�yBŹ�qW���4CxFX���ǕZ��6�#Y�Ww-���
�h�1B{VF�e��X�]�w�>��wՄ��К���*�B{t��\�C�1J��$+��Qx!D�5�
L�����!��?2�w2�Ǹ]���Ԙ�z��������1՗�u�Q��BL�а�_sѹ���d6%��.{˺W9�3rfd��\w
Eݕ�+B�p��WR���YԺ�N�ri�9y(�9p���fĻ�j���u��m[=b�׌FRU���Xh���yp�Р��o6�۩ͧ[��z���L��s���
����	6Z������q�k'7/�D\���R.j���DS
�͎[��oZ1�V��̩�֝}���s�5�V��<{�/j͒�X�R�_�N�9o(��E��v�wf�c�q�1J��)^�<�\��ط��ڰ�j��r�rf�R�U���;��7:/K	����[�.�BJ/>������/�4-;����y�r\^�w8=+:ޱ�9��U7	B��pk��.�9��O:�t�=r�$j�"��'T-9�-�aF�c:)2�e	 ��
�M�h/s���֮+*�yO<K(� S�m�zt��L�#ߢ�2��*�M��F3"�Oe�m�uS�P@0������-f��[A�P��pp�|�3T7@��$G��jv�K�nV�[L�����5{u)n[�,��JQ����Ǻ_3�Z��n�s�害-�"5�8�Zr�?�&p;���͹F�oN��\m.���`Z��u�k2[T��6��nЮ��;{�X�i %w&�5��f�Զ�Y�S���V��iT���VS圱�Ձ���{�6;���]{�`gC�5a�b�h�#�{�ӛs��*�F(ڶ��JI��Q1H�[=E�l1jcSsO|gm�赍�h:�l�f��}��P�ht��j�J���I����)L^2w*��x�{5^:�U�o:˲uW:��f:��B�<NGօ��Ul�R�ad�+�uڠ�\�ƚ&��!w�L�F"\��F��;=o���.l���j�mF�o
αܢ�S5 ��y��G��w׳������N�9\���<��ԓqb�W=�;�*>9�ZLc2e���@2���\R�KkVv�V�]9�wDv*����NƩ]�PHA%Me���d룴�6e�Wu��u�S�Y�y �s�����	�7k��.�7�@�f���ߣ�9=�*jH�E��+oM��+f��#���J��7K��4�wJ�(�Q���Th��37��M�V"���H,(���!�{�	6�I�A(V%�t��Lk.KY]�R�@���B�<�	E��R�Z	��+:�r]`��j���~>~�-�ӵ$}�,Px�[�mL+�8:W\�/����}+"��A�r��8}�����GVvsb���
�ɖ��R�P�e)���[/{9��a�yB�Ӧ:��8� �n��,�*�E�o4�+ֳ@�Z���[��t��uaǷ]M=���P`����������Iv�ϔوꬢ�dT.a�$��f��+�us�V����vY�j�C����xf q�����9�6�f᜹	�s��D�G{).���jy݈�W[�ҷV�T�%9���fP<J�
��cڽ���U�J�Wne!����*�ls�սeXt)�X&�&�[؎*�]
�]�fM"5�����ԻL�H����uU��1�!j����`T���+���]�/�["5tQg7��lE��j���c'�suލ� �hyq�Z��֖c�ْR��
�ז���E*�^seB�e�5j�E����῱R�l��h'��v��㹍�V(/Sˎ���F�晜o H�̰b�b�jr�c��{+_u�(�m�w�l�4)���'k����V�<n��n����w�q��w(�a�ݱ�P
7�Ə*r�ƣ��8t�ND�o7�syۉ��t�܏���a�Uٜi�M��v|�?L��A ���Zwxh��*!���OOwN��m�9���}s�Eww>��t�(��ȭK�㲞(��u�U�_��?��C�%�a�0��e�"ȡ�*c$P�$+p�T�1`((c�E��&!R,��Lu%efn`j@���T��2�&1L��E	�5�&e�2a���
bjUf7ZbT��J�-����U��f2�\�5����!�
æ�e��S�S�WXf�J�\�\[�b��k`��k�QDs^��Q�[e�t;���bL̸�������Z�\B�LBc&m*.��U�7,�	�v��F�MeME7h�ek5�"�XVV���"�X�b�f�YYm�婉�
�ms���\I3,+$���& T���dQd�U�Xbj��l�b�*q�J���2�F�P�j�a��mJ�Y��Ad�SX�@���j��s7n36�URk+�!���VDe72VV,1�*�u�Hc��"�J��5$��R� VLV�v�h"��M�
�\B�����t\�0���!.�-9ۗI�0"���^��k6��#sZpor��ϝ�:B��q��Sjs�����z{ǽJN]��>}|s��[����s��u�]{b�����׫��0>�J��z3��1!^V��.&���pϡ��{*ũ��W.��,��n}�U���TL�+�I�o��g\VX�eז5��:{Bũ�8�36�'z/A�F��l57	S�(6�	lʓ*�3{^6�ve\`�Sl�e.{p�YQs39}���.��ΣOqlSg ��yI�G�e�7��PudWp�8���kF�9U,z"-��g|��2�<��BV3��y0s��}ZI���,�m�[ͼ��ˤ�#u���	6k���>$�d��V�������C������W��̈́7�nu��kF%[ǕOVdD)�'��[�a9��;�8'��L���#}H�u'�{�*��{w�T��Ħ�G�������o���$g�h)��Jֺ��
Յ�u��5�۲Mzs�����+�lo�?�
f�1�ڔ� h��i+�<Q��gl��N�WP�����[&�AL�.+ܢ�
��v�1�q��	�Ip���Q���|v�8�v��0-3w��iC��
��E�T���E�Ժ$��{qv��Y|۞����ݫ^�߫����V�7%f此���ڤ���C���E�D�/z뚟r����m�͊j$J[�Z"�^NS��QyW�-va�_nK�4���j�*�-�弬(y׬gEûU7ؤE�ϥnl%1
#��{����]�P��E��~�W�T���F�����*�	�6>\�]V�/ˈR5�������ܪ�]BV�f|�%�>�.	����(����w�����*/�2�ވ|�o-{���pJ0N�'&��4�VGg.u�M��	|S!�Xtȩ[~t��Zճ��_]���M8뾖٫�����Y��^䩋��KfT�\Ι��y����.��s��SV��w�مν�a���I�-��u9� ��C�U��pg�[<�v��d�ڼ��t��q#e��qL�nW��9؝CK�h��\��q���bh��)or���x��K�v��u)3Y�ԯz�R� �4��t4�Wg8�үM�_����D�t'h���է�v��of�ė�Z�Ej/�#�_V���nQ��evc!�%9^.5�v�*f;,w��v�V���������gү��_o��=�F��Y�Oet��b���S��Iwr鵔_0yVYi���$L��׊����(^U�t2���U9}n&˵���=[�
ټI����Z���s��hT�q��e/n^O����[]cZ;K;n����:�"��s�kNDMc���[B�^Ⱦ׉�w�`�^4k5ϹM�;[kU�z�f¼2} ��{)d47;�®�N˷��P�_$k5�rR*yzާ�2E��7�]���P���r���c:yׅ����H贮���-�mFUBڌ��ת;�1��6�5���l%`<�C�z.�㞴�^%I�3�S��ȡ���GJ�5����yޱ�_����>J��ؘ{�G���|�c4�����1UZ�I�j��n��r�\'���:_z i�#�kFq�l*m�n�o?�EP�M�I~�`�7Է��D�AiwX�
��sx�nWC�s	�U�^�'����ݥ�)6�NSqU�m�\�v�l���j�\6������.�k�<��;��ZhoL�w8���ɮ�A''~����/��f`��;�^��lN�v�Ζ���A�^���NLe�3�NukN^�oe����M�w�mx�#��.Zȭ����nw'���� N��=�%��,�b�E3��as�6��A#,lU_6�"ʋ׳�֙��$�X�{�*�����������s�����3�oZ�J�0�9��J�$�:�y��d6̩�txN�-�n4�h]��M��Ш����J��j�2�$�j���Ѹ��h����U��W��(�j5���֔��F�:�(]�@ƶbRl�k3&���W~hf�h��Ug!�ё+;�/4�[�/+�O�6P��:��Z1![��2�CZI�3������.&�4�t�s�w+\!V���<��]��-V��#�~����urEa�律~�UR�+j��j�oP�BE�f��甩��T/cq�
8��9�/mb�,l��etO`�m-Q#��`(���u/��[�չ��Ar���m	��gF��L��a"�Wz�w��g_ ��_�U�5�b�6���F]#ʯ�ӌ�f*��(�w;�;]�c�O/Ut�;W�ܻ`}���sO*�,b��u|9v�z�f��$��c��jVU���̋�E�3-�=f:5�v�1y�,7�O..���/��H��e�9V��w<�J�ҽ\�ۨZ�S5��j��%UmϹo+��z�tW�-�2��yv�Z��b�	���'�e��P�N�.�`bYC5O���ǋ�:/6�r�V�ٶ����9�U��{w�+�r�F���lBw]�@��������UZ�m�Z���,4C�:r9��yBŪ�����[�O{r�e��MV�bFvR��t�@��2�;�T��r�.�8�fc�S�Wc�z2��"��fs��#,So`P�̅!s�	�i�T�YIǱm��NU���A�4f� �~L��5mbGqlPl����&�ٹ���lEa�4��1�-^^S{� Z��F�&;>U��7���7��k���:%՚}��!	#Y�����]jn+7`���#�e�}��M]v�XB���u�]�-N`=闘���j7i�Co��ZV�v�q�|a�]Ût	��y��J��8f}�F���И�K��A�/���S}��o.��{��]����V̢K�U�(�(�����]4�HI�Ѫ�al9�F��wu9��X�؉���r��yB���S�+��aQ��SC#���̱�Wf�ʖ'����?+��[�.�R���8�÷�^Y��5�ݼ:�-w�aJ��ޝ���n��xtk�g�uNֻ���b�Q+\���0�v���#�Z��J���ߛv�={�*�5l��5J��Kgp#sB6�"ch���*0홽h޺��r���:�m���PR�qω�7w*E�\���%u���uRV���N�}��}Ӝ����)x�j��S����`����^���z����վ����dbƖurv�h�/�ᵣ���r.g�Y�y}�Zd��;�$�i�9�Z�v%�\�QxF��({lJ���T����d�I�f4kّR7��}S��Fj�e盏2g�1n`7�jS�y�РWM����<d�A�	���+��|@����j0�G��"�R��"M����|6�'J�l�n���i�=�N�#'}�.�]��j�_�,�;�d�tVލ��9]b
�{�>��qo/����y���w�**�wН�s�Φ�/��2ä�ɽ����9d�qM�f����lVf��eu{mCͣ-��1r�@�l�ReP�t�<uy�ݞ����3���I�xg:�U�Ab��[��4��ɻ{<vѮ���#^� �L^�zLg7�4�ʢ���fq���'ø�b�i����ө��69��6�BV=�U����[������"�s���Ǒ�>*w:
���,6n��y�<�C6���(^W��ߑάQV��d�x��>^�7J���b|�����y�1�[!������ǒ��C3�צ4�h�Wu［Զ/��֎o�<v�v��ޙ����{�;ɬ�u�-O\�i��Vrߩ��d�+�����^~oWT���q�a<�W{�yZ��b�|Um[V�,v��/�;��|��T���]J��0{fb��UC^�)f��1�4��ׅ��]���N�9u��[��l�a�8w�|1�'���b�f��ЈǠj���R�\� ��ר�3�p޶�w�mfu5"+�.T��v�����e�r���fW\��t��F����uj��}�����5���U7��?
[�W�V�R�����3|��i]�<��e��0���gm5��vGW^��Ƶ�n�	B�'7G��Iɵ}|{ǽ��p�_sW)�/+e���]����3������t!�P��z�◷*Xw��G��h��8�<o+5H���W7�#/H�Xw�������S���a�����2�_M*u�}{b�ע����>��ї�=�ZVF=��.�bAɝ:X���~P��,�8�mY���1\{s:jk�lř��G���Q9����	�i��:{��/���z�����)ƛx:!���O�'�#^��;�v��>��*�E�7���C�����Gj���n�b3����S9[f|�!��׽
���Ok{�^+9�4�>I	�u�R�D�cܙ�4n�o����	I�MJ7`�^U~�c��B�n*�]�C���Ӻ��0J�7�`V�I�Dc���;2�Y#�ɱ1���*�k\�K0TpTSYv����b[a���5��zL�V�9M=19j�9�b�[{բ���͎�|���l�j�3=Wخ�qJý�/�{��������s���Υ�]O
ny�S1)6h�2l>&1\F���ڷq8���|�����sr8U�.���(W�ָ�h�+x�o�"���oU���L��*�o=��$D{�IU</�W�|�c\]J����9}�������m ����B�w��<�ͷ�u�eg�j��j��B�	��g5�¾S�Do15ڻ�~��~������_j��ve�bJ2��h�+(]��I��Y�A��Z�����F�n4�*a�>�\����St�H��e�*�nVO��(\@؝�����EeB�"ё|�^%Um�弬(�v���n����%Vi�Ù@�}�}l�{۩����į�j�y��U/N���3]��+�-��Eb��*ʡ�D;��o���k�n��Rg7�s�E����b�M���ˀ�ؐ;HR3�.�R�+ky�|z�����}N�F����S�9���Eh2�/�_\�k�B8W;�4h����G���5�ީH�m�=}�4jN=k����4�NN�� ��'��s�zq6:��X��^ś��	�5Bp�Ф/L�͝��Sl�(�q7"^��V^TL_L�.�ʮ��x =�����7��l�����z���2��K�{L��?c�9=������d�'3�T��ic2�����%�*L��#����t�:���o��kv���r5QX�φ'�a�űA��[eA�ǅg%�
{٘��L�3I%.�-fc�Y7O�~�h�|S:9SP�ܜ]��=7I��T�Ǝ���s�6�ԋ˦�nΰoS1>I��Sņj��ة�ڷ�ܿk&+���m89x��Էy!����<��v�[f�NCܳ;��+L=��c��ܴN�{�͗���Qά+�S��]8k�����g�St3��c���6ӯ�0[=�ANӬ���>U���4��S��e;&�wf�R����W�vn�D��(c=[[��ӌK#��������ݗ��I�䎋�|��T��<��d𦢀�Îu��h����_�g2*mC���b��R����V�GN���V�#�LΫߥ�K�]��=}��v.�֪낺 �ꌠ������V�!�a0����k(�e�����ö�sӶ��tζq��Z�-��nU����xvt�ق��ly��*ժ
*,�#��u%&��}Ms�n�P�k�u=�Z��:����RU,�s��g:c�2�u�����8	x�W$31oj�X��K�1Qw�h]:�ۮl<�{��0��u�<�	ۏr�\wE#8����rޠx.�+��4;����'�7����_Pu�Vc�L8�F+�.���87�V\���QCG(�)�=�[6Dg]kje�g(]kn�>�<Y�����Riz0Z �O�����Ż��c�rn��cP�,X���y�.�څ�6�i�Ӡ1m�ύ+�y/�doM�J�nJ��$����n]���M��q�� �����2�.��R��~�]~�d�O��)	ld�t�,��Sin���,u�֏��0���;�TMJ9��!2�M��K����;�nG.�pc`k�V{.iœlva+�VWC	n����.���/z�Ȣ����{k����m\���q4���z�^����6�ӝ�]Ū��*�`��v�m�j��\ ����bt���V��X�lɓ�*� T��˭���)�xvmoes��X��j���1���5���o|;��u���a����!�.b���f��t�s�K������QE��:��w��y�k��P~�V�l�v�EL�l����|u�G���h��;�j�k�J�5��s���Y!e���YJ���;!wku���&Cy]�.ݫ�Lӫ�{�Ƹ>��%�*����r��8�"���Ph�Δ�t,3�L&���*�@��f�.	p�\&j��=Rq�{	�%�Nիk�F^�AC��wYQ����ޕ��d5�Ҋ��I[��hFȒ����ې�f�����ҫKc�|*��Uٶn�S2�9�n�9T��sX"VJځ��՘t��S|_	�Ό;�5����Wh�q�|��:��������;���=�D_vQ�H�j������
�yW��"Dj2�����ԡ�UZv\;
ĬΔ |Y�e�Ú�>Ņn[i_v�9:Pbލ�LL�t7��\]|�����8O��4k���t��m�:j����&���R��܃��L�ir�[��:��T��OI�Z����͓y3sOy�2Y��=�tY1b���%�b�Yܵ�I��K���v�q���׽r sB��pCB+�Rw�	�;l�����;Kfs���X����S�u�n�Q�\��s^:扽DF;ޠ{na�a��I���˷*5�Z��G3j�J��h+:ĝC�N���D]mu'՝���L<�t�m��vom�9�+����wN<G(�`iv�Eݴ�=����]w�|����O�;UdX���+'mb�cr�X%��b��&��L�$5��&�%d�:����QAE��m51��(�ȱKl�-�����5��bCX���aP�P�2VXk�-aP�"�:���ē��˴3,UR*�4�ȵ�e���`��u��,�a��2�ԩ:jACQf�ƕ�
�� TnպɏI�&0�\�Rn����tʘ��`(�[b�Y��jTݲ����
�LzۉӉ��E��l��ȭ��J�E#h(J[Qꀰnb�Z�
�ՐĚ���m1�����j(��N�cu��+��JũQejk�=e��²��u�����m��Z�Y�X�+	�E�dĶ�eed5�L�F�j���k5̱E�e�$Y=Y
�MT1�u�4��å�0����=_ǝ}��u���وZ'�~�e�S3��݌٘<� H��K���WNտ>�r\��ҮCp�'��t��N��Rs�~�����\�[������h��e�Ը�v��kyo+P���q|��*��N��|nwT=CgŨC����z�z�.3k��%���������S��U�������������L�:a�l-�w*�:��.���3W#�O�:m�Y�7>���޹��F^�Ұ���YBũƚGU�l����i+���6�ۨyt5���o7P(K�)��a�b�4��@u�^o4�w!���jr��*�jmn��S�o T�eI��M�X�^7��nmy��v�߬�=#֎��/^�0č�ؤ��"�n붺tlL���i��~L�&s�ӷ4�n�]5�t��cq;,q���ۇs{H��Y�m�W+7e�r��D��u��tu=*�=�D�|Q�y7��cIZf���c�z��P,s����4n憰`s�{C�=�X�����＂gW%��%a*Y#ݾz��9��a����Q�ZN藼r�7�{#9��K�JT#��om��n�i�T�%�yY(�J��no]j\�;AR��'��9v[WV!��8��<�{��`�.S&T����2����E�9�j�;9��Ø�W�� xx1X���s�>�>�:����ww8�!������}��
�bs�V�qyDSR��1���_����㵻�-�ѯ�((z�MN/xf>U�\��Uߥ��Bo5��r��K*o�^�ў���ps�co�j��eV��;wy��V�#���w\�򧃦3geU�O��c{�m��ٺJ&���}Z/�VU��̋䍥Z�F���Z�����z�<����n��R��̩^]o����W�f-]ɍ�������`.u^�\�����觥*�P���t��/<��黦o+�;�ʅ�.�N���բ���+�azGJ����U�s�*��%���[��!���U�]{p��k�Vu7����h��1t�G*�������2"����@�jEi�CmY�s�S
+�/"c��>�4+Q-�{�f�
�1,�2�ZF���+c�*��@�P䣾������9�٫�Y�{�B�^�m[�\fl���q�+�C��y��w*�N��T��n.p�)�ݲ>��{�R����w�.��0bVzƺ�沗��Q�z�
ib�{��o_jK��+������c+s��gF�ϵ�U�\�^iv#��d�m�<��*c�yD�g�L����sERȫ�����n�&9�=��^�h�;�l!�R���8�1�7}��i��=�t��ז+ƙ���UR����lGre�Pq���:�n�hF+Y�[��/t�ۖ�o/��P�]�`���JM�fdߟy���I��Ddu�ԟf����!�{����P��o|3e
�[��O�/8�y�Vv�-���0=+�W(�����ϟK�<��&Ny	�:����p�74�r�=	R��A��v���R�k�{�y���1��-j���k�>U4�	�L� A�ѷW��k�f�����T�|��a�ݛ�D�%CV�R��v7y�$���㻑P�17N ���V��\�yt<��Sb���+��C O�!x��Z
�f*�U��v9�%	 ����v�3m�Kt�&��e=��@�n��{om.�W:�2|;u#�����()x�@k-{:���x��Tm�S#��>٢�r{�mǜyN(����>6v�l��R�9J�Wo�_��d���?�wtj٘뭨�W���\�{���&75M��ܟ�nt�k�%�J���-�j7��gE&[V�VQ�S�][��Ṉ���r�w=P���{�fj�x�ީ���v��`��*5:�[UU�K�S��]��6W��P��]{b��$ o�m�	}]/�fI��,�Ի��~���£ݶ'�zܩʞ;�I�N�z�_e5p2�x*m���_H�Z��xSu��2����ڕі��X��xS�yC_i��iBm���1,?���H���0Bx��r��q	���5���us �OY1��a8�SO�!v�>gG�d+�P�N�0?$��=����n��Nh
�ױ���K�
 O�����4�B�ԇ����*ɾ}��I�\�8�I�����E���a*��i��Bq��~�
�	�μ���ט~��ٺ��\��	�0���|v�sz�?2!�w��'�;���$8�~�d��,���w̓����k�8�y��xɖ������>�=J�o��u7��	�}��|���2��I�����*C�;g�;�d�d<OS��;H|�Ӻx��铈q�{Hz�Ro��d�&{�I�d��t����7���77Qk�qh�"yW���0@	ǽ޲=gS��d�HT�����ĝ��P�2�eHvô���	P����wgL�gY�Md�yHv���_9[|��k^boUݲ�1]<4�}"D�F�f5�)'�ó����i�1.Z��X�Hbf������[2�Z��v�*��rܺ�����������ܷ�R���XѺ2��9Ot��r�ahU�<	b���K�b�J �I��%l��'qT��۹�(-\������{����X�u�����t���s$��&:}�I�$;�0=`z��S��`J����0�1	��}AC�z���n�=C�������y���'��;6���Q?����y<I���a���?~̒t��y�|����2O�x�`w>���z�Nr�����1	�6w�
��~Hi�:��qφ�#�c"�?u_D�˺���]w�E�x����Y8��Rty@����̄����0��I=Nr�ĝ?0>�8��Y����CO�$�:�<4�#;��PQ���ljΊ�ߣ8}�*3�́�����q�ӴY'�l:�>�{���|ԝ��q'o�'�}����w�2N!�?0;�2q!�SYט��~㯴��6�J��� ��>�xI���H��C�:d�w��O�x�l��!�>d�i&���a��'��0>I��y�^N@�́�of/����d�����}�!����1a<N!����M�g�c'Ȱ:/��?2z�9��;C���l���S�O�a;��|,�����3�O��r>c:���o�^$�:W�{��>�>���9�=g�8�����O�Vo<���O]>�B�~E���	��<j���>@������2u��N��'�w�}ό��7q��gu$b�>�G���8dx|@�:��	�!�^a��I�����S�R��$���I�7�0+'��^P�䝵=̐����ޯ����򟢹���9��ω���>����?'����v�Y:��0�:��!�&���t��q'��'tɈ���'�6s!Qa8͟y�Y=�A����u��vn��Yڒ��πD�{�ʧ�����$�M�Y�<B|�y`q�'Y@;Oм�8�����5���~�d�I�&#��AN����YL�#���Rxئf���/7��6�;kjL���Q�RlT����y}c��=&��4�x/#b8j1t����_j�����䘡`��q�O�>���9�`oZ�%���>�E�7���s�}C)�=K&�-TH�d�:�K|rtQ�ʛ[Б����Gv���� � n�-KS�w_�"���>�܁�F𫬟��bx�}u�>`xé�;B~@ެ��!>z,P�'��$�.d�@4�ܩ8��Y�t��c��o�s�x{���?0��9��&�܅�Ă�����N�SR��$��������{N�����i�q���^��<f�!��9C�Ԇ�����/8�,���?��!d����ߪ�|�J���\a�
���VkW\N���N2����X�u�P��٨V9�����`��x�v��fN T��MT�֐����#�|d���s���g]o��;��� H�8s�,Ԃ��{�L>E�!��q�e&3�}���,Y��y��%eI���a�x�&2q���=�~@�}�&0��n'�o(jAa�x�f��u˦zӶ��>sw���!��
z�S�,;f�2q����%���}�Ԃ��y�'2�H)�}�q�'f0���yl��S�~�X�J��
�1���>�)��=a���#eȨ���X>����ye���}�3̡�N��!RV�z;�L��B�����}iX{���*|�׼��P�%N�2O�Ă�g��5�O&�~嘞�Wԝ�&�\!��w��}�OMn�`�w����������������VM~�k���v�;��!Y�m��ΐ���'���aQd�ˌ�����}uY;eC�Rw��C�|g�*0��X��y߾e�__}�7INw$��<	��T���jz�SyOɊ���<�욘��v�OY۞C��t���gI?3�ygi��e@����*�L{��?:ȱf��Md��'9�w�Ot}r�ܵV��K�0�(��}�#�RO�{����ܜI�=C����N�M�}���d�����$�����9O���|��a������}�Ne��|;��'�I>q��>��^����,�r�oU�����(���s �z�ߩ�=aY?2�ےq:O��!�9����9�:O�C�+��k5��HT��3X�yiS�7�|ʞ��wN��P����;o|w�����}�IWB�CN��V!�gFO����bQ��L6f��v�ò���81�u8��qUw,[Sx�䖋�+���x�+I� f���Y��-�K�|���(����F9�hqt��\��ss�Rk;D�<=ۊV��� < �������2�>}ꋉ?�9@ǉ;x�ÿ,1? W䝽�s�����������ϲ���8ʓ�{�Y������a�13�-�B�Ȥ�x~܇�L?0�	g>�آ�`�Ec+��O_�a���ä8e^�@�OS�i�N��`T;߰�����'��5 ��<gG�����S�d=N�!�a�9����0�ԝ'��1zH(.��aQf��^_A_�LƜ#"r�5�����F��T������=eC̰�}���dX�N��&�q����T���ɟY�?!�S�Ov�$�8��'a��R�y��t񒢜a�u̝2~}�D��?{���"h�Ӂ�{�td���%�9�`T^�|�]�{�bP��jq��=q��\��Ƴ�ꘂ���7�z����䪁ĩ�=a���|�d���MC�z�B���e�*��ۻ����q��>�y`ru�:d���&Z^���N2�3��`Wz�8���rt����H=���L{Mg��$��}C����!��u�0B��c�y`y�N2�z�����Ɋ�J��=|�V|>����1���1����'HT�)+��`kXTS��Y8����Y:q�>N��ΐĞe����y�t��:s��]XjAghc�u� ����V�b��u�}f�|{X��Fj��'���?[9����:u'G���� �u.aXqT���jN&��,�s��,�2��O�u��8�E>ˌ�J��T�?`(jt�Ɉvg2q�$���B>u�(N��>��k����z;�L�?Q䕇Ht��v�R
p���t񒢜g��k%eu�O>��PėO9�q��ί��s,ĝ>���OI�=}�;H[`c]��<LA`p�4�n����]��5\>ߙ���$a��'�k1ĩ�;C�_gl��Y=g짞�Ě�T:�Xv�:d��w���+O��*d�T��쓍�Pף�'9n w~¤����}���;�03e�v�}rǄ�$H����'i��^`Q�1��r����<e{7�E����vyN��C��N����t�O�a���ư�
�Oـ,�����2��2o˵���M�?���
�~��pBt|$�#����̔Ȟ�`��r��t�q��{�,�
��1���{5�<6-m�K���dlu;9��R��Ho��p��7{"�&Z�on׺��`m��g9����ŷ:wt/���|iM�tΪ� ���_2�b��=���҂c{{H~I�/���և��<s�<�d� ��O9����5'_�ä��*Cm��=aӬ��<ezH):��YX�Oq1�Ȳ��`*�y�A2�}?_�D[�2�Q�bA	���Y>�,�x�?y�$�<xɉ����t����3�s!��V�~�?51�;�§�t�d��O��$��+����m �����\H+���S�ޏ���^nߠ_,���g����qğ}u������j%A`z׾s$�t���{���ԩ�:O;�'l���ju>�s����J��s$��t�}�����L�2�C�;���u@9�7��X�|�o+�K������r�Yû�&�>�w�H/v�?}�i>@�_��v�;Hr��}�M񟙉;�2q�!�jo.�|�>���$>d>��]��'�l�u?�k&o������5>�5��:�pPO̩�>a��1��i��$�/̝�MC��v�g���Y��������>�N"I �} �F���*�pE�c������ϼ �G� |%HE!eIyC�?&0���-��T��uI�桌�Y���y��5'�*v��K'̩>ÇS�pC�|,g�!f�=���7g�����?y��I�1��}�@�N2���£������`u�O�q��H~�O2�{=܁��'�!ߔ��$>���gC��,����Xz¦�}$�Fv݋Z�2"�f��U��~�7�!Y=ed��2}��*I��:�5��]���Y?2�O~�!v��q��jc'��A}�d�N��Om�~�&$��u{N�
|�ۏ�:xE��EQ��Y&*0�͔�Т�� ��~f!ɶ:��u��Md�+����|�hc8�l��`ꓴ*j/a�20>kN��J���_��V��3�����!�M����P��"��y+�+��&k3>&����;B��?=�d��S'FP��
x�����$�8�A}d��E���	S�<La��2jC�ɉ��gHgT�����y��Y�%a���?y~'VdNlߙv�,[���J�<�L�� ��.F�N�&�w��kU��Ê)b�t5�۬l�Y-�O&��F���K�£�+�{�zp"R�["�	�r .�]����S7�+Y���f�֭f���aQoR��*������=��<���>�=�"��?��l������x��|����
�~@�;B��1������@����Lܓ��H(u���Y8��9����3)�� �1Ŀs�{��_=s�y�߽}�������L�!��>�.��TN�y��?%a���8ʁ�T�;a��2��<g{C�*!��M`V�Y/��Ɍ��y�'-*I�)��!�{� �$e�(�_�w����~?!�*xɶ��ϲ���'�&$��E���I��k�nR�L혏,�q!ݡ���٬�2�u�<u<C�1�C�����i:B�_��#�|�>����?X�}�K
W�A ,����:a�
��vs�%f��O2���ɨbJ�'��������������@�����C�H)�v��jN3�0?yqR�� ��o�j����iE"�����U!DW����Y�퓁��5e&05�u�,Y�Jι��O���y���1�&&�����T5%z9�^��cl����1��T
��Lt�܋��N��F+4}� �~��ė�'q�)1!��7ߺ��AN�;��:I�ć�N��$���Aa���z��V����*%��i��æMegSϰ+>��*?g����Z�w~�{�=�j�7�|>�� �!Y=ezJ���@��t<f�̜nRw-RT��}��AH/����:H)�z}�E�'oY;��':��������4����i�QǓV���r��+?2t���hW�!����'I�'H^��)1��Yúq�����������Ğ&�zʇw��~��T7��޹HT���>���Σ����<�>�|�S7�8�S��8u��T���o9�Ǵ�3�<�d����}���'i����f�?[����9�������"ş2^��>f��
����d�2|>�_~&{+=vY1�q'���g��]AUV��8}�k�z�q���5���1�w��QN T�3���:��9`vg��>IY?"�yΰHyhvζ�H)���O��~q���y��5��)ʝ~1@�\�U�|v��K��_��	�>�1�
�u�uiS0�c*��˧���Q7U����!	uo"pp��䣦z����T���j]���	��gdq��l��
k���q=f������L:-�ճw#���S����R��n�ʲ�$���x�1�\�X���Y� � �~����|e@������c'̥�x�v�Vp������hnR��yJœ�J�_r���������&��J��0�mE��O��Q�-�}��N^}ө>zMH)�}�5�N�&���'6�D<gG����RN�ݓ���eg|���|��c:On�!���Ӟ��b)+�^����5�y���O�>t�,q='��Y���Z~���W��x��*0�����%{g�:w��Cݤ�~C�{�LeO�*q�i�j���u��v����:� jV��sgI>I��r�*,�[/�i�=�}y�����
�Cܤ��p<zdX��Ϸ���<B�wW�Md�����i�C��a�<q?2~��Xx����I��*~�'��퓈��:�MC��t{�AjV��1�.�~ԗNM[Dx���>�^�� ������I��M묜����5*}u�>z@�+�d���ë8���c'�~�Y=fe$�_��M`~k:&nI��*N�M��TW>͜��͞p}���� ���Ͻ�*zɭ�}��%MOO��]�$OܳI��jC�0È��_SS���>�D5�wN���ui�q���^��:��Hc<�_��}ne��]���/}��>g����X����u>�+�8¢���	Y�<a]q:���v��T5:��{���q�w��+��HT��`��x�v��E8��0�W�,�<@��j�i�~���F�g�����Y|,�G��� 	J���Y�1'^}�L8�*CoG�|ʇ2��ϰ��E�1�=�L��&&��a�x�&2q��3�ACީ����\&��OP�����_op����󷺔�g�q�QB4l��B� T��^�?#�;��%哨g0Z�R�۲s,Ă���l�{I��;�̇���x�9���ƠD�>}�>��k1���`�����y>O�I�-f2z��C���*J���tɼ�*��1�'֕���5��T����f�H(x��w�'��Aa�v�'oY=���S��6EH����"��{>��J��\4';W��6��a�Gg^S�tF�L��w�*�#�@���r�qb����f�MwR�A�wY[�X6��2�Y�M�ֽ�������,��}�p�%bʬ��csr��(�b�-�WX�>����B�+�aT����y�1Rٕ�$݋©QPl4kdv�.�qn2iP��ٹ*�kk���f��M���_ K�d�وힲ+E�}�w��U��/��Q�	��X(�u�汖`Gj<�`T��4/��8�t�O+�R�� n3G��fٳ/���J�oV�T�:��L_Yj��z��Tbn�M�]ҹ�HYS���Z\��w58/��b���e^�;0�K�-\/���ͮR��}՚�k�@�2	�8T�`ܶv�u�9���6�ΗB���a+��Y�rk�뜮/͛�}ԫ+�6�
�.2�	|iU���|�f	Du"�+3�<7}e�黴�$���i���N�Ǖ��w�՛P�Es��y��b���+V�ȁJ�����z��+N�쭇Eu���ԛщ���Ÿ��	Jɯ����/��*L{�S�o
���0��)��_2���GD����&�r.RC�� ��A�0=D,�n��/2�K�yV�ͤs��J�޹�_jU��M*7Qvո�%�Hag�k���}���fɹ9�,�V�5y��J��,�w�x~,��Nx�U1����Z�h�K�n��U�Ֆk).�u��q�vzn�A�o:ܒbw��R�V���9��]�:���r�Y��&u��.coW�u����=�GU:��jT���>�҆).ΎW�Ǉ�e{�`�v/JVf��|u�897��Úf�)�+Ԩ�r�˝�x�X�*u�Y]v�4M�&�x��twt�<ѥc�Cu���=]\���GEh&���B����j��ɏA3ikv`X6fSp���P�o����ԥ�|�Q��6����6��:Y&���]��C��툟w���R3W�i<�x[rV������+.eti��>s���v�k����pmp]�h49��s[yܦb��0����	L��L��:\���p��ݥ�d������yҖ6�=�(�b�9���he�ײV�̾9��;X�A�_s�!��_Bkx�k{ �"�,����E��=�C�{[�A�+*%���s��S�/!��\��֕��r�mY�U:m�F�T*�a!���3E�f�MŒ%R�}�w[z9��._^wJ�J�j)N�:�&��u;���y�r�3�NmٷWw��v���;�:�57oK��':��k�q��(U;E�d�%�y�H�13���b������b�[z,��Ⱦ5�J5PG�^���!Y*nSJ�y�O�顦���}֢b��w��X��O`�6�}�k��Na��w�%"��]Z(���3��C�����[�:�����g��ӹ�eI.uwl|�ox���9N]ӏQ�N#;��ٗ���ń���1�����|%đ$�2G��.�&�m��F;T+�c�N�`)�Z&5&1�Z���1MaU5�2��E�Q`�RR��p
�-F�Qea�RJ�j��C\(�i�f�¨�.�k�	���)5�Y5�tç�]�r�mY+"��X�L�:�JʬB����nj��¤P��]���cGi:�f$ŵzV�V��k�N!FCEU�N���LMe�d*AꘓR�u��%���`�(�ZT�P5�E"�!kE����,��C�h�$�e����jX²�Wm���leJŷ1�,Dƙe*]ʻje�咢�6W30�m���Ķ�i�P���Z53%U%u+��c��*��kZ�Ul���bt�QU-�Y2�+��� �>�g���g�Y�#�"8��pg�m�8���ݼrF�ٗ�x��u_���Ҽ�tܘ���Y	q�Ǭ�O2uqQ�`��۰�gZ_��x K_m6n�2����Y������!v��+&����������a��$?[;<��5>E%I���]a�N��=ea�
�~�:@��T=�'{~` ���<�`OWT�w�j/�Ù��a��l~��Y�3v�9�S�
�γ�~LT�����2jb~a۩=gny>�HjIY�)�,Ԃ���<���Ȳ�tyO�d��e&=��?:ȱe��g?{���޻��|��}�ܓ<eI�sS��Ld�<>�:I�?e8�_���1��z�t���'I�&�}���d������+�'��;>� �>I}��;EԂ���Y9�bAϹӟ�Z�"���dk��T�4��h�q�1��Y>��C��PX5��a�?0��2�����ퟘc�9�u��v�tCu%�T4�HGk�EՂ�Ibj�w�
�9�F{!ڛ�E]���oB6�3�E��	�8f	(��:�v$wT�����Z*�~+R��Q�֘Q�-���m�k���6��ɬ��@�3���(Uu���p�)�5�ע�fa|>����\��Z\=fv�N��i��Eɩ����;���|�P\E	�D8}�=���f��gbv�`C�{�?/V�~6���6Vѳ�O1J�M	T�Rfh;Rx��k��2}uo��xc����,�����y���H�e��Kq|��`ۆt��,�*�sp�/�2��:���p}�d��]� 3$^�s�k���J����;��b��jWdx�C��9Y�+:��+\�����u��6�[���@��	^�T��zY������_W8��}�o`�ha˩���Y��"�F �S&wY��;+����lP�|��sҏ&�9�����}UU��!'����T*�?�����İE�L�ft�S�ȟ)�,ЎY{y�Gb&Gmkֲ�mv�lԣ����^T��d��B���
<��Pjc"b��`�J���:�#�m^�jCX<z�^A`���^�\\T]����:��<�6a��q%nE�=m�>�L-Y�]̽s'ÖEɢ�͊��� s�E���9�:��<6��
)��.�fL�'_���]��n����%�g��_��Oy�4��ȥS��N�]A�7���*�v�nܾ���O��a@gVJ6����Lw�x��<5�>�I�ġZ\�v=��s��ʙn\F��UH�9�4�n�5��a�Ō����40|y�u��9�"5��5[�C�ܓƁL����n@w\�#\��8�FtXm֙�t��p3���b�
٪��}�O�	�Le4OQϠ޹v�7�g6�t�s��u���͘�hX��M���q��'3��M��fP5��]0TΛ�eR708ϭOx��Yw������5��}���o�Z��&�^w~��p9~��(�5j%Z��!�z\%�	�&�z2�[�"�!����k"�_�%�8����ԃх3�w]$Y���S{�x�A��ƙ�7p�Ĺ���8-��ˈM�U��%��#-ϰj�4��+��|�U{���=�Z��vv���d>1�8=!ֺ�3�_�yh�p��.��)yAN�-P��")jX��ݺ��ֶ{�j���gS/)�6d��,0KK*4��-�1k�KM��U��NI���gT�`TqR�k�h��p�0[ufEӮx}�}aa1r�n���^���оy�7��F��S9!h�[��Ͱj��c�S2�$h�L�*��Fv�4zmWz6{WrAɔF��Zg*�����f��C#"l�t�bE��-�n0�lT���&��cr3��u�Y<�Z<n��g�����a˷��^[���
��VY'F��3zz��֣i�ޣfN`���TW+&�Ơ�J�A},����.����+��y�+��z�[L��};�m̊��Jyrh�sUx��� i̤ǼkZY��˶��b<���<
-�w	�\��M<�3A�v-�{aglA^�c�(xpb}èp5�Ky\^рM0���G�2�uB���Dq���-n֙��i�C_EHu�|t������Y]�w�(����M�rI�w}ulⴇ%0�N.D9��B1#f�4J+C��%�S��%�RC@�J�B���Ǹ�u�˼v�R\"�HXe55$�w����_W*{�Gw��U-	�gۤ��5*��3yg}��8c1��DaK|ꙻ򑇍�I�y)��4��5��X�
B�6�׶n����T<�z-$��#QD�hV/��73����Z��M\^V��edr�eK��̅���6��*��Փ�ì�%BjR�[%�
d+�0O�.#y�(�>U���ɑ�����bg&<<��k�<�	�J%yϙ�J��#���S���P�ZN�N�աC'p5���ޢ�� �����Q��w�1�,ޱ<b�{Pz��ę�u�cbٕ��m��XrY�.Kj�u7�5*C�ڜ�>���z�Yf�}K"��IF%�@<k�L��l��&#��.�sM�}���%]+����x�E��PdH���I��7ADF戛�qMٶ���5<94A��Fv"��{/�!�4��j�Ε{/c�	��9�SLEq��N��n�;hwwlq���s�*��	M��B�7��h_?#g�,'�|tm���8�I\��+ey���
�^#!�M�;&-ܳ4��"�v 3ӳ~�U麔E�Q^����a9j�"��@�Q�N�N�L�$�nn����q�+��쎅<���j��4��:����5��ѡ�n'���N�̹q�o��Z�O*.�[����L%�J�]��"�UˎM>˴F�ng^%M��;�
��u�=Dc��[��V�^�,�ż����J��㍌�1��{Rk�X42ϩ�8f('l�[r]��5n�E�rz�ﾢx�@�U�~��ټ�]}�8��e��ѤA��H��~Nt"�+��H�D�9Ɇv8mq����9���=�5���no�LB�{���k4TbP����j�%s�Ì8p��0T[{ֶ#6�+`�j$9N�x���p^�=�aɝ�������h��ɲ�\��e�|��$xK��
�J�*nnz��-�b#Ն�ʯp��B��sv2ͻX;AK\)б�}��e+E�����z3xfɳ�&KL_�7���һߧ��=�PO�\<�U=t�g�q�W�9M�ݥHR�����'�LV_y�(�������T�BI\���~U(��B:i9���%�nRM	�ȹ�T��1�9~R��x�c��t`m��wx/�sC��\� ����ev�����N`fXsClL�`VB�8QU��((ބmN�:�Y���3+f���;���[�3��-�\��J��k�|/(�GC��蔹l>�UKu�����=�sDU?e��Y��S8����3�}����%�#!�@r������Ҳ����t���ɻ��9a��T[�r��7�ڏ[4f|0��5����YCu�o�ݺwҖ.�L��eNʗ��'y�fq�a���ҩ�J���*���E���(Vj��{��]�sL]VؐO���<	(��G�w(��N+ҧ�����f�eAC��^�����M�gS�xGJ�5"�r�S�(,1�._F�X>6�\���k�a�5�Z���I<)��!�+�����.�:DA4�f+ə��)<`MT�t۹gl`�FF
�O5�<�D��C���d%�,�Gѩn,r3E�a�:E	r�PUQP��ڸ�v۵�Ʋ��ql��칝YT,�0c#"���Р`�D���`�lΙ�t
"&�l��nMVs)��W,��>ù�;PS�xW�� ��:!_�N��>%�������z�ٓ�fav��uQ|Lz4N�&t�K�o�Z������*�|�!gx:S���g0DT���V��Z�L�U��d]���A_oY�:x]yb��u(.U��蒇�,���#'D�D�}��g2�B[s�^YKa�n��EA�{'��C¥���:��P���/�s4Z��W!z����Ɏ���s6x�s�R8�>�׺]��=֭R��E>K��p���{aU�u�g]�þ�(��j��
9~��;�j�Ì-�/�8�x)KM,9��6�°+�L��ʶ�e��dP<���S�e"�	L�8)�/�˝�h�vr�Q[]t\Yw�pbj간�o��Օ��E{�	 �Ϧ�W�Օ[�V�\��¹���6n��Bc�^���UH���a�H��Zv����I�2�lk������X����f�u\Ez�I�E#@���X�땄hr�l�S#:,6�Lؼ|Vt�$���ۋ��d�O(���n���D�r��pR�����+�E\X�H��,�s[�vv������zV��@cX��f�.�FP5+�FTΛ�Hߦ�<m�����=�{)�1ǅ�6�z�ic^�F�2|g�="GhN��B�9V%�n%����Q5�@n.�j"�*N����#J3Y���t���g�Z`��c[��0t���msB��bb�0G
nrܣ��*T�k�h���z۫2.�#!�3 ,3�.(���WT�!-6��ɇg<�7~�X��9!\<���f���h�T���ȑ.Y�����x(��2�3[�u[YDqgV�.I��tg��;6O�׆��U
�[^��U�w�goc�C���>��^%V�ވv�Ǽtd���ᗖ�:� ������
x�r.�K�R������/������B%\:^9+wzq�n!�x��RQ�[��]�q�MS���6GN
���\��icW{�k:^��Ȯ�ɢ��M3Pf�jn�}X�b��.i����3�p3OZW���!kv!�ӧ?�UW��o�eBD���F�9&59>Jɯ1�<S�_K0{�é-\>�^8������v�;���m]-�0R�E��<L�v\�2
����S�l�Td^K���Z_CT*���&� ��$�hd^��N�."k�+��yXr�>�1��L��ck�p���\Ku��-/�^i��`S�NP�� Q��E�dk�~�J#�����[��[�0k'��b��9Ml����y��l}� '�A��D����iR9Mz�;V7<�+r`�,�)�	6�SެD�_v{�B������l99�o�t�?���O1X�:8#z�,tXk�x��<��ʎ�����k�C9�%�R�Z��sGE�U�y�xթq������֧��o!+�]^U餧�lqV�^��:�l9�3�uZ��>F�H�o��m�"r�v+R�6�[˿zg�iL�]�uS�壆7��b8�=�<YI�����%K8֊�3�C�n�O]Q���OJ�ĩ�s���^ͤj�Yf��Y�IF%�@<fA�vk�q+وnbA�k�V�L@�9�|:�C��"�unzk��y��{YW��[�)]_m y�
�@�6�l���0of�M2�Zͼ��..U/]�g+Y}5�2{�ԁ����}]:��O&���+8�2w]8�$KKf�i�]�{������rgO{�,�/�]8=kÑو���¹�������OX��n��w��6���}����}��N\�*��T\������23`���jܗ]����T�nkg6{Wh��G$?S�Jfd5�D˝2G
�Xl��"��B�6v!��W�R�w���_���Ɇט��2�����O�����[�f(Mxj���u#�M~^�]jcLb�s�wV{��Q��OL0W�2ϩ�8f+��3J��*MG�%��a�܁�(�ѳ[��)���e�Pfn2�uƑ1	#0d׺�.��|UVy�V��> p�s�D9��cRq=#&�&w#sԨf���˚B,dau�`�T��):q�,F���~���}�zslX�,yէn�r:\������6V��gF7�폓�v�>c��<�羞�"�U�c��ih:��݌�t����Pw�«#J2[�p:X�]=��(P��ݽ0y�u{f%7�g�jë�;Cu�4ʎ�ޡ���V��z"k]/7��I�Jұq�9�6b���b���$nI��e�e'ݡg_�o�U��h�Tf�
<r��b�\�q;xCX�.6R�����e��P\�ʏ7�̴D9����0�}��D��n<��c��}Sv�F|
�k�vgP���t�.���b_���0�X�OK��RTG���BR�j�q����q�NDg�W'.�Z"©Gt�k��j��Jb�`aܨ�^�t�/إ��!��7�Yэ��P�BU%�#%M�Fui8��Id��
%����D��2����N�!w��oB6�i����}c��Ҽn����f����\�8�)�X���k�蔹l>��]o��\([���ݬe�F35�Zks�vi��d="G&g�%�7�G�w(�+��r�9ip��7ޣ2�#�`0��μR�ihc�.\��nQ��H��/�5�8M��P�O��^�E��Ŵ�Ҋ�Ot1*_A�ed�)�"	�.~��u��!��ma�>�^�f�k&Jmv4o3G��Ɓgѩn,r3E�n�*\����c�FGpWhZ}�j�bX^����fr�cj�𻰍b2�����7B����m��1BYd]�;�y�]����T,�'�Q��ùN?r�إ.?a ΥDm_�N��>&}��ۨ���w�`2��dCY�j;bZ:sf�N.�!+��M�@#ٜ�7W�Z߮��>�˩yOpS�t�zC�.���aʔ��Y\ῶ��b��A����뙊�0�n�PH7MHf���J�sf����n��J��*X� ��w�
kI3��2���h�f��i;T�_hź���G��8�C����4L��G:�vi�	�Z�p�:�S�(�G�]T�ҭ�F�b��� )���+���˝�Et�����T�]k;�u�Ĺ7�s�8\��b���@�4�,-N���iG���p��k�dz3,gCKvFsp�\g���y���R�f�2���g��{�NYQ��]0غ+�U!غ&֧&T���� �G ���|��h�z̧��qL.�YN�'���Xr_-"�9.&9�ػ��s����]V������;��m��2�wh��.f֙҂��l�Ku`n�Q�o�:�*c�x �F��[����2�m�����`�v�^��i�m�tc{�x�B��_�9]v�y�vjr�J���o9����2&gm�={���\��A�t�]�q����p��ٕ,�<�\�M��u��z.�S�(L�u`�]a��X�?ku�*s��urT��nC
�8���IY)=c
&�S�{J���B�oVuf��l�<.��6nV;x,�\�)<w��T,mD 4;U]gZ�cY�Mh�6V��G_K�U���ָ�X����x��������컭j]6�>2��yVFBZ��]�ݔ��o�۾�Ѿ^�4��k	��8کg-2im��Æu��v��[�Re!��gB~Q�u���v^q�l�%eIeݰ�=���e��X��CN��;S�����2e�;z�����	����Z�Q@�,C���'�k����aal��/�9|U@��A=Xq#�w:�`g1c�3���U�=�	�ZݮPQ�N�v�fˣ������˖	��f��2r�5ҍ`�W�wn��Eӹ�r]�����Z���7��Y�	�wN��q�i��[B�Zk�U���72Σ,^���)����-��۬W��!��7��5������j��x���YJ���Q���G��CU]=Tz���r�Z��O"sG[q�4�h��6Vț��6:W��䝷��H�R+3�a�r�zQU��u��M�.����4p�����OUi�
��h#[V�W:��eR��#�jt��HYpiθ��}39��|:��V�}|>�%�(�w^j�.��V6�b��&3%4��N�;���U%-\�"�mWsжW{������[9��eSoL��mr�w�4g`w���n©�%�lfb�';�馪�FFZ��z��d�5���ۤ˃�Z�\:Wp.��;#�\�{��I���S����N7Iq&����y�;��j��w����5���,I+)�gO[G�'fJ��J5T�y�^y�����x���L�v�P�W\e'���Ƞ�*H+Ft�X�6�q�ӂ(6�T�X�K�d��X�J���6��,b�#5�UAIXTT�c[JuB��Db!�)Du)
��VV�Q�,UQH�#��X�dUQCF(���Y��B��fPX��֢�cX[LT"ł���X(#���R�E�Ĵ�m�!U���u%Lu̡D��$YiTX
*��U��ʊ1�k��q��Y�AUb��f0FEDUD�(�Pv�AP5�MtTv�%���2���2��LQ���U.�1���V���k+F)-Kn�Z����wrA",��iE�ZbZ�D�J�TDUzI��(c**miP��J�
4��SdfYiib-eX�B�2��KUj#j�c+VḚ�*�2X��T9a�����uj
�s�����-
��#`'e�r�Jw��O�o&Ld5Eݵ����n�^8��g1�4�1��%�l�W;��'��9M���.&?��L�5%��`�
U[��寚��h�)O`3Fwt��&�;�T�d�p�Oa�,s�d�"Oڈ;�Z<*��
ŉK�C�2鸱�4P��:���Qq�:&�;ލ����̎�qK)�<�uǲ+!
��R{���^E>~��;�����u�B�s_:1Y ���(�uXx������g��\�,R��6�ٻ�[��;cu�sn�8X u�11K����(r�F�9�4�n���֝��0/!�v�����(�1���H���t�L���H��|�#ʝ"��)u��k|�]y#Y5��]�d�g����������8d?h�|��T4;�c%q�B0�R��o,K9����%lb��&]� pGJ���Y��̪F���j8��f)��h���]��b�Q܄�kk�����c��N����.�-L��3��D�~j�.L1آӾJ�VD"��Y�c�p�Gk:�r�3����-\�%�L[O^bo}�a�yʤ���7���U�`IÁ۵��Ǳ>՚��D�A3��[WZ�4+ku[�.c8�Ç���|=�;���@�Kc�}sk���p�ө��o�!�ksf�#�[c!,�v��z������������D���uz�[�pT؅u�(��p�3��Y�b�#��W*籒f`��Gvuy��>�o�k�{��$-��{��Ͱj���e����U4I��7�D<�oOg��Æ���,؃°R���+m�r�և��-�͓�� >�F�X�/��f���M�;�!���1�D�5L��3dP>��Y>M�������~�#�o�k�p�wc����a'��f�9&k�Y5��+����NE�j����I��í��d��rn�Ѡ9	�<�JYqќȫj�ħ�$P(����dy���Յz�WS��<&ؚ)��̋qCX�49K��y^dW��Õ��O�uɓT`V]"r7�M�\��P����r>`\+����՚��ԕ�|L��X�k���v��z��a�{]�7vS5s�`����XˤjÚ<o����7��� �*G)�+�j(Xj�u:+!�&PL�p��|�{f��)�9��\m��h��ƽn@�}(�����6PL��ܽ�&��uzKU�ΜM��dM���2�/'̬C���a��VB����'C]}���z�G���|1�i+zV-"��a�Ӥ����C�}�m��g�0F�����gaUx��9�&)�}�u&E�Hdɫ���m�ih[�PN��M��������~�=�ض��p��֐�<R�p݁b��5)E��p$�S!\!�'�R�u�D`��9ke��*�#�C)f�F��⑇�Ǉ9�m�f@��P�2�p7�������]���q^h����]��c��8�P͑j^�<�z6YcX�1^{PGT28����S�X��e����Q >�Ĵl�O��<�T�r��y���ͤj�C,�}K"��(�Eb�}}�"��hǔ��˙��d�� In8�i�spNo�Y�:�za���T�]NC4�4�n>1�t�!TE��v����u���9�bxׅ�L�`�>���׆�2g-VY�çO<;'�����T~��_�%�9#�;�25A�RN�H�u�H��Xl�<f��B�w�6�it�D�r}Ԝ�$���`e.�t*�s�����y�����}D׆�R�����{�b��'=y��rY��p�!(����z�	d
h��NٚU�%�Rj8���̉���uys{��%�ۯ�v�ύ��n4A�BDN:`ɮ�\E���g�,��f�Vג`�R�R
��>L��Y�k����o^T�RkH�� ���7�fN��ʭ%w ���8$���p�{ޔ���ݓ}k{� ��)�c��ct'&;;M�"��I���:+6�U���V%��78e�,B7���L[�Tf����a�X��fe�l�����τ�����\Lxo��2�,X�. M���J���W.�v�RaofI�e�\��#������&w��I8v�Y�;�eP�40��5�N�;�m]����AJ�cT�9�7<vڿg��.�X����S����:3e�)qq����w���ai�6x��R�-���c���>K1�c��t��e²���u=t�v��{i׀g�^��g���ș��ˈޏh�!�6�[���:�v*�עRW'<gf��Ӛ*q�j�wt����)q�J��Y�P4�C��tcn��e�gD�\���m��q�U�d�
F��v������jld"��;dR��F��khź<��X�J�Ԑ뭰�ܿ5q��U��G�O�Qz=r�}x��u�K�8;Gu%��a����	�Y5��+Ľ"g�5��C<r4�>���4�Cn;�#m+N��5,߻��Unu2�S�7",7(�y��6!�=����`Ю^>�u��P�d-�mNR�&�oL ǈ2�]1{۔N��wV�U��mK��F�y�d�UG�u�٘]�Үʟ�i^nB-��������Q�X]��K�{��9�R�|�W_8Szfj�ܣ�U.�e,V���V�����<��T����BM� 3n(K�رY��e�D��L�f$-����5�$��o�k���ӄ��7����i�.��5�!�,�����bK��t�3TT.ͬ&��ktW^o&R��/Н*��]ײ.�3�̄k�47^�`�D�L�ft�k���w�UkR��v0��`�kтk ����]#�c+��闃d��$A���׊�i����m�ls�v���B}������9�5�$i�&t�K�sc��(ײ�8l�C��h��;s�&]l(&O	])�⏮�i���Y'df�93�a�(M���n9�*Il��s����d����f�z��4���m`�X����I�o3��~5yyjڲ��/K�{��/(��?9��q��C<�V�����8�.��nt�t��ꊇ�͞�w�«0�����U͡�����dj�S(����n�/\��٣r�L�s/���\_I�w'M�a:T�#@��t�����_�<�w��f���C/���^���s*wkgų���W<Xuۻ�Q�4'WԂ������6��|;,��B�"rûdK�ל���}ͻ��K:�9�{"6�f.�7od6Z(�8jy��c�F��ʝWQ�F$�ySki%���k�6!ԏE߾���-�*�1��&��k��&�R2kҔR���՞
9��2)ODP��V2QWJ��'�f�pk��ҷ�ה5Y�{2�.�B�(Һ49�p�̢�Z�v5N�\�&�)��b*�d�?H��+ٲ�z���ކW�����Q|kE���&���e=���p�Ս�fT%e�rl��)di�R�_�J2gS/)�6f�28��	x��L� �B�/�z#y���/�ʎ�>^�L'��\�@��p�0[ufD�F#އ�� ��!u��AX2�'��v�Ƹd6}:nGfJ�)�R"��!�j�j��Z�w��oq�S�b��*V
G�����#.ևW�S�6O�/)�+��GWdDu7^���!!!��b-�b(K!�J�T����(�FJM���o��^|3/]wQ��]5����̂x��A�7�e��1�^�/����^cPx�����E��Mj���t�{������N\>��Ɗ��%L��h�dU�Pa<�#
'6F���G�:�@�[<�cg �`���K�E�;�jL�O
z�� 3{i5���n���)}z) E�H�96�V�2�٘V��<h�dհ�Y�ُf�d�3V\��9�t�&��ܝ���Fk�;n�zktQ4�t/ܚ;�}s���pÛ#�,�̖�{
�z���� 1����^i����"���}�%Y�X�89K��y^d7sf�\�R0=��^�K�W�L��T��#66�)Q9W4�
8ZC #�dU�|N��+.�m^m�#��w�]�-8){���C���u|9�~KC�PV��3y)�����4��c̽u}�Е*;��#���>�UV`�'0p�3=q���7�'�z܁"�QQm���<:[p��ڔ+P����#\<R�w`X��#�_Y��LerU���wKF�h���d+�|��dt�6�̊�(ݎt�[R0�4ꁝ�"�%R�X�{�G.�Hj��0�W�ϔ�X۪r��c�l�P�^��hs��GoK65��������q;]����8rgH�K�u�a�3��ɯW�t����s�=|3i�f��Y�wes���M��c��	�����}S�k�{��X��þ*k�Y|<��k�z��s��D�S�<�j���`Pn���8 �>Xgb(M��C62T\��t���:�x�Wu
��1���mG�Iٝj���R���%�}S1P�g��mh��%zib��I�H��j���p�x�������Wޜ6���-ُV�_l:�-9�[ö��ĺ9ѳ�Mv���IR�b�Aώ�:ǧ*�]E[֯)��d�|M��GR���xx:q���LEdyt~	*�#=Mxb��>w�u�� 0�ߞ�*S|�|�N'v� ��A�o��h�VED�5*!��)�^��E{��d�,��r�R�5�����xLy�_t���
B?v]�O��l�!X̘���N�K���@|�w��sȇ���U4'��C�g�uz!��*��l֋N��P܋�8=���2ht"�)�>��v
�]�J9����[��`ň���z%r�7 �^ͱ�e�˚B,dau�`�5K��s����w��8�WlA]�,b�0g�	͋L�G`�D�u,����5aN�8�}���uR}f��*P�,�1�
�c��9��S�ƟN���Bё�h7w��4V�q��(�$e4���򎰵�SS9�|�if�UXo^R=gC�b��,�,�i��u��+��(�1c�'}{�.���5�,�����G)��6�[��� �ث�����AT�9�k�β��x�թ�8�z�(�\�D!�Y����~�.{����'^3�MMs/�R)��4��Oz�Ǣ�㍴�u��E���i����t����2�Do'XV���ܳ:٥S�!��vr둘L�ޭ+Q�u$��;�3{�����GBo��,�Zr��6�[���	�K\j�)�rn�PB���1Z;�a
�X���n�,}��\�G�G*��[�CI�!�]��2����������J7��t��=���ฬڑe��ͧp� u<�}u�p�F�:/G�U.[��8��`�ܚt�w���ґ���h3m�,��'��zD��&k���x�i�}��B#L���U�5a�w����ETL�s(����Y���u��E�(�>"�!a���R�6#<aƓ�r�cVM�:��v�b�0@�ù���(���P�o�L)f-34�=����s��wg�b"E�N�xqR����3J��^ �#^̐�x��hR�r1%��8|Ĺf.N3�jPs	�X�jVn��������_.g6�YrJ���\�.k��z�����KU�<�Q�䴏f掰�*�^�R"�?��'d{�l�k���������W�茢75��	{�Ȏ�g�P�``�Ң(71�1^NɃ%�j8H�JL��N�ތܔk.h����e���3'�}�u��y F��Sf>���>�1<�.M�͊rg�Eu4C3v��q��.;M/)�ěM��.|w7LĹ��3ǩ��Q:=x��$�y�[Jm�g�h��R�7�|�vR��J7XI�o�L�:���w�	�9=�W��Ew�����d��]݆*V�E��6������|�Bmp������6��n╧3�/������N�VE�����b��k��g\��Y/!�uǲ+#��,MULN,�z�+BM��o4UܱKz�9q��G��n�p��o�]&�z����Ɠkoa�{�&�>o��5a�i��,:�m2qF��UH�9�4��"�Ԫ���~}P��v��Ō��0L:�9��D
�OOp=g�G\�#<u�{V�=�������6�i.Q���R���՞Qۀ8�=@.�s�W�)���r��YR�B�h�Cn})oXH��5��6�t+��@Ў�ѣ<��y�H��%u�荻�	���e�!d#I�G�C6Q�ok��z��x�="�RuER8�DN� �fx�5ev�'�UC��R6%͐\qmC6�J5�,�sƌ��!i�^�*�@�&�o�A�2+���dZؾ���5tx\�fH���8Er����n��f��u��X2{���蹫HÄE`Yaa.������6����t>�\|��Po�5u���[OI���U�0Y��am&���ڛE�`����i]���1F����:�j�p���Js��Ev��6�AwƵ�j%p��(S@��ڜ]��o+��\�+�։L���ՠi��и�K�i�̭cl�m�覽b|֌B==�FlDr����HI�T�̺�*./vV�>��Kḥ�ͮ���?���.�u0��a_s��|�a`Y;������b�KH;��%�\�^hڴ�Q�9ūu�H����{Cu���u+�6�M�=�%"U؝gN����5H�����R��'�
Z��q(�9�|�L��لc)en^mB�:Z�T�X�_
=�]�k���K.����+��ۿ��c2������;�˕y�����w�8�7ؓ� o��Q�51NG�Ę\B�ۻ̀�-
�j�q���B�0h��y��	�:���g"K"Q�Iù��cs�w�d��Zoa�O�/�F���Ve�O%� ՑM�X9jhMVyw+�h��a�P��A�3P��t��Q
k��xM��Kb�[�h˄im�n�_%�S�ݷ Yy�U,���5ݜ/67�$�|.ʋ��,i�������a�y�m�yGL� 3fq��p��Y��S$�����%��Z˰*ݺ�B�B�nN����s]��Y���F�u������c:i�َs�br�K�����4Ӄ�iW'��Wk���P������r� B�i���ъ
#vqlom��\���	W�����Vt�\3�su�5۸���E��mrX&]�uKq��GS�@(d`�nɭ���켏X��-����%�R2.Z���(r͒�1����F�M��yw\�qc�	�>ad{3��vK��@L1��irIf���5Х���|z@�;VQ:��36:\4o���*Dmp�ή>�͏�Wjb05�;%��3`n�`��7sw�K5յ���� �9��2����� �rZ�	���Ӫ�s�u��v9�'bq�.1���Wi�f�,ʶ���-���S"�ۏ#U����v(�X.j+���{V���Z���5+x�k�٭l��WI9]5JV�*|溻)ʘ� �I ��㎴K6ͮܙ���Gi.���1�Lp�h�W��ξ��ܳ��J4�m�ʴ��2��'��]�2�9E����H9��͒�C�S��y��Xם���p:{f�CW����h��k�ub2�8��}��l^Q�ǎ�=��a���oت�s��9�c=�|����_7�&و�с�7\�+B� ���&��<	�GB�I�ՠwE_%
Қ�U� �����mL��U}&��
[�am�ENw`0
m��Աǀ��ݖs2s<g�n�,���;�iޮ��f�kx�A�v�VQ���Y�^ެ�[FJ�k��ݭ���'E�Y�\`��M#ml��"�)�0qz�ij��MN�����L΃��Ҙ]Þk]�6t���Dq8o�Z�aUV�ޮS6V�V	��� �b���YDe*��ŵ1	��lƸ$X�V5��0֢�Z�WY���(��Jҹj�1�Mn\����2ي��+iV���Re*��E���aa���%j
"��k�%�����X,���V�4����¢��j+�Mʳ)[j��DjTQ6�J�J�3ȍ�bܥb�����V���f5���Z�]skJ1E�e�"���"ֈ�Z�(Ȉ��5j(fb��wl1*��ԭ@�aLjAU��s*Ŵ� ��LE-V3�p�;h����XTUDA�"�c�T�TV*�Ҋ��*k�#*�-h8����1��[X��8�"��(��E`�E��TƢ�ĥ��B�PX1+Q��[`��(�b�TY�QEVm(��fҲ�	-*�[DQ"�(��[e�B���G)�Eԣ��mK��S-1Ab!��Z�+b��+*(�{���v�����TLJ+H�p�:��S�&Ɇnc<(��{�;v>��d����ـkv5uX�U2���]?��
v>���l�i�F����R�b�T3�
�I�=
�I��]���h�f��K�ƻ�R�&�pZ��1#ň�(.2��nF���q
L�7�fȠ��Y|,9Wo�(��A���Vf�pm�q��W W��Ug�
��w��-��_�ɯV��]r�f��a�X�ǌ��t��Y�(W���u-\9�ס�����@�J�q����A�O.H�Ov7�O�.��(�'�z��,Z7JL
���}�$�k��kg�8�O+���޷b���D2uk�ճ7w9�ȑۻA�k��Ë�	u�4�X�Qt��c����w����G����H�#Ù���!���&ۭ0hk�5�ER4}�3)
�j��
��)��)WBF�)|�61�p�E �hg`��J[���������Ò�NK�Z�Ы�p�jyR��93"}\�z�dr�dX�/T�p݁t�	�J-ld�t)������S�gv�[��s����\Eb�"*ԣ|�+c���8�%C,��P�y'����5zpCI�n�B2,Q�ۭ����#�9Ӟ��V��Q���(�A�Z^�;ILǻ��s����onL��,:���͔������u|���;��ƻ��Cuuv��1Q���%��m�P��Ƚ뮙��]ٌi��z����6K�|�=��&�G�j�u�.�"�)g�b�E�F���#����`k�!:1��Mf�Բ�s��~�#	
���u�p�v�̟=U-�W�_[��i���;����k�f6���[���1>j�KL�>��{��
�a�5��/��)}-?o�Y�q��T�!$;}v�m�`W���)���6#گa��4,\�W�t��v�(�N��#/�{��u\����������؉p�H�w�S3!�RN�T��$`�U��1�ڪ)���<�ת3/*�s�؎5��xЉ�Gq��JY�1��x\�=�3=�ۜL&7�Ǝ^n����j/S��O���X���e�u&�����@hř���1��5�Zj(���N$/Ðg>U��ٯQR9q�r�i�BV:`ɡЋ���]:u�hYo�����~���&$u��k��Y˧���px:��Q�Y��>�#WQ��S~���P�ǽ,%�	������A�D|H"{�^sN.@Xh�VY� (iPt�h-���3-]��^��M�Jq�S2\X+`����N���]��2`;�)l�Gh���Z_q:�J�Mn�C6Z����&��.W3��������o�C3n�{/�6&�L\�f�?�D�/��Pp/b/8���w�˻�v�{ѵTw�jha�{U��9�x�T�������pU�?zL�)�=(���L���g+.y�UY ��>��<hr�î�8UCY>̙|�LT>����u��]Ի[����%�!v4���_�`���`�t��/����!�6�p?o��S��{>>߮r�7\|�Yoq<y#�P~����k�O������57���b�r�R��;��:5[#�n7#l'{ɴjo{s"��f�(��T4�rۨ������M����t�B·Jfs��v�÷ّ��OPf����~N��6�(�U�׳(����7*z�"^llȝ�{s�y^�~N�6�C<�Y5�X� ="GRf�q�0�:�W
�a2+\y=�2��y��z�G+ ���W
!p�O�:Y}N�EFU{ˁu^�O���״�#�R8�(K�Ő*�q˜��_υ9Q�ƨ͊��,��K2��*��L�N���N���t�AI��ڑ��j坱�)���9�d�kŜ;@Է�I`�t���v;[��ݛsժg
�Fp�u���/[� 9���Gܲ��͜d]�|�{ Y"Dhg�x��D�Y��*��FX����kGa��oo�c��@��Г�[c�,X������P.�K�A�"���]v �����̀\]Fe�F���(�V�ؾ�6+�%�����Ϊ*6ƺ��'���w^Ⱥ��c2���SX�z����̥*��]���w���9V\gL�_$Ex:;Iٔ}�w|1�v>R��y�eT<��uj�Q�;����,AՂC�⋈j"�c�`ϋ�Ў4������Z�^����N�V���ܢ�[�#�	�cS4%)l�x�봝{QoY�W�^`���r�\�FF<|�S��"��WI��M/�g5Z~�<x��zϻ�z6˳��~�a���pqQ�ʅ̉l^�s1�K�@޹�R�^��@׮1���:�7�^YH��;�]���!q*���M4�5s�a�O>�l��JgMl<:�sh@�t���N��g�
bB+��&�\<��4�j��S�3�7rt��'��)Ȁ��xSWp2���W��������kR�Ҹii�Z8�΋m֑6)��/��y���e����3��b��d"w;%�4j�\k
Qw1O�oP\�^�� _L�T�!L	�]{w���i���'.�/.��v͐�&e*38b���nU��<qDn)O �zcN^�n�i�Ǳ���d�5cQ5��g��_y��꫅\	x�<��wύo=��Pj���elYco�lAw��mv��}K���\�'D_-�e䪬U��a�����M�|��eB�?	�ȵ��HEdVl�B���ކP|g�PzE��By�Bin����d��{��#��d��-�.��/()�Z+M���#J5�,��Hٛ�G��%�5�C�i���F��;j4��n���r_[�t8��5��Z�b�yxWa�}�$���|���7�;��̆:��̅�v"�N�f���g���C���蝊�2�*��fS͎S��\�SE�`^D��L�*��F�di*]pV��h�]���Z+}o_��{��>��i�E��G78x�bE��e�r4�C!�`Tj��:L��q�dL�f�@(��>Q����:�A�%�}S ����22%��hL��D�Ȁ���ͱ���,�^�.�4^��7�q�U���˄��\h�!0ds�"R�\E�g2)���UM�-�Zl(���>�wd7&{ XTd^X�-��%C"�V�8k���y>dT���в#�(�Ls��Ĳ ���ſM��{��B�-��S�r�P��B+ #:��Nx�l{�M�s�S]f{�N�N�Y3�uw�����C��jZ�י�5fT좹�����x�5�wS�쾱j�%\��ĵ�в���:�x��C옫Q�eDv:X�Mq�	o	�G��8FEI�f��8q[�g-}�3]t��
�-��e���\�0���>�ݭ"l7Z`־��X��jê�}���� ��ҺL�gS��TD���m��f�HV�޺�ͫ�0i9�����u�� �Yס�8�=0`j������Ȁ�*.p��G���tȰ5��8w`KR'})E���"����Q�r�1�]��S}�2���:hZ�^�>DU�F��!di�K�ボ�Q%�z�뵅��"��s'�[G�j^�|�XϤn�|�tEb�p��{���#����)��Z8�TM���c���I�T�C#�2:]v�l�=y�^%�H�*z���m'���{X�o5-����������X��H{PZd	��~��d�V8Mk����Á�N�e=��t�X��R8�+:��r(���(�pAfB�;Sj���͝.Q�@_.b6{��率5u�rM(Y	��6+���،�,�u�S3!��U:�$7n��'�[W�'�/{.gMB�qӝ�g�qؙdP�24�vL_��0���W�.�6�=�v�{qK��1����ӕ#���0�/^1[3�Ո@�B�,�mb�i�f�r���:��_L��}3�����n�*���;�Q�	j���	'܅����l���^��|�	0K�t�)�v���+��	l��.�@u+�Ir��':?�_U{7�V����"=;7]>��e#^8C(�DLf7Rk�X42���Ѥv��)��Co���[�1�����&���Ql��܄h�T�}=�H��'��|/�۾c��w��O��!o �ɆtG�6�Y��{6ǲ��C.P8h��@5צ\eax���@��ՓI�oO�_�B�D��J��`�.-��;��Ȯ�a�m+��Nd%���t��`�z@W/�9��S�ƟH��RmgC�ù
�۔�onr�,ec����0ku(͖}�K:9Ua��)�#J�ogٓ;�t�}͏^�s�iRT�<w��逘l���V�:����[A�Z8���i�oW	w>��j�ȩ��TU�Z��5��p�����+��!�t%��+�)K�/�(��,���qFzx����ja��y�!�׵������30�ID_J��ې�л���܀�NUC��#[
����86�s�җ�3c��N�f����c����:���G�ᒍDt5��{���������.��=� ]���vI1̗�������,��ݞ�0o��۾-�6�ٴ;�Cqc�|{[=N'��ףlJx���[1�����qe�c@d/w�д2S��ZD9r��ɔ�5û�vjk�ؚ����*sVwn��C5u�B:m��ޥ�qb_x6]v���"�.n;���mw���7��Mf�^%�;5��0�F�G�e�FI�Kw��3x��z�����\�g	E�r��gK/���ܣ����ٳ5	�e"Jǽ�^��v�D3l�
�U�f�((͊�AG,ا(�&�S1�����_Ǚ���Q���4��V�S��%վx;�^3�hR�_#4X2 �opZI�w�wmun��yyxH���a�'�����n�f22*q���{ʧ���g�_Xך/.��)�E�v�63�b��D�H��gi;0��p�S��9�[������ջͺ���ley��2;P�@�e�5q1��0d��G	k�L�)V��9m���(d�|/:�q�u��s���,߲0��$��lД��⏮�i���Y'<Y��b�G!<����)�E��V�#��i���^!���QK)�<n��Ed#��EH�+#9�y��b��%Q�$�3jtR�^��@и�ޔh'U���^YH�{y�ޑ��+�A5tW���S�+}1���Q����R�ٶ�'8����`�kN��w�}څ"�h��B�F��Mf�+q.�Ч�~�Va�»�l�!�����=s�n��ٲj�J�mr�P��'P��v*8����MD=}�
�ؾ��)$�ܼ�Ί�'\N�}N�9\�=(���N�N�^��ʩ��,�nm_7�WR�"�����֝��zf�w'M�q���U(���t�L���H�5f���fc�b��ҕ=ԩ�Ft[n���t��J%dk�Vx`�(��8�4&VB۪t�En�&++!LC �w�2QW��9oXX�{Ʊ#:e2�t)����]�+�e�;�l��νh���E�Ui��S��	��͔m���f�����P�fk/SW�n*֨S����)r"����s?~�"�O��1K9q��gS.\�Fn�h�w;�)�%�*��!�d�<�pt�ϰ�R��5]uO/�ja<lU��^@���r�����9�!z���)�1P��Xgb.T��k�g�E�g��PW������H���Ά����Vt�����`�,��)�1AUEG<+&��+�'F�ю˞��S�geh��fj��t(�[(��
�q��[r4�P�C�RfY��6E�q��}�5q�^�|5�޲w/7��]�}����n�Hr��Ym��zػVу�z�C�OL��ܻ�;��b��5�ռ��r�%�ܵ����F�>ǜ�*�D�<����,⵸j�g):�_Y��d}�wn��wg;�`�[�e֪DL�_e*��8���_��1[�J��#���ei͹e��&L�r ϲ%��hj`오�У"�7��9融6��{�jAń�>��:�x9j���������@����̊�{2w��Z���qhMR�u.��A��\�GI͑�c�:2//�E�� �pd[�b,�K�����n����c�C{;�Cו�*����=�ţ~U�����Q���Ќ!SG0�wF�_�H-.�x�R�F�a��6�ZE��kH��{&.�4׷`2芁Ѿ C��_R�+��7��l*�͞0�F�)M����]<����S��C�",_��ns|+|�k%�,n����o-��W�/2���(�ʥ��t�̀�BR�[���OUf]�4�f�Y��Pyb�n\ES�EZ�n��H�+c��(�;�}=����u˯w1'������(��pE�̳�#H�^uC�J�����Q/e�z�#V��^]���\�Bͬ�,s�Sڂ:��Ğ�=`�%�g�i��=U)r��g���ԡ�?9s���I�9�^�kF�ۻY/�bz�vB�s��ѹ����Z��õ�5j,'G��C!�a�8n�aT�Jp��7���社�D�R�ݰ�蠯��W`���-(��|k2����eb5!�w�b���1Hv�ۚ�D�\�9�ꡉ�����YL�x���zӕ����|��k�Nn�2^�mK&PM��k:�m·�N�Nt�j�aU���>�whֻ�!���s��Z�ot��4I�(S9�kz�:��u%��+[�[�i����G]�� �">�����m�� g(j켴�~�R
E�w�c���A;�ixG��|2�=��e��#�rmK���Rue:%}"n)g/E>�<`��w6w@֟1�_f�Y޹E5�Oc��b����z�BXD��1���wI"JTĸG[��Ab�tMlǗ�r;��zT'Г���$�*SԦ�Wsbi�\�l�=S�XXr��N�kwCWd+��z�W����)�cL�-B��R�c�˅�o�r9t���9݉�)G �;�n��J�w�|���h��bF��ݿ�uvM�D��}�MYC�e���N���������0�K��s/��\�w�#r�KO�(<0f��'i_(�b������\�VM�jc�`�U�+L����}9�t�a�q�[+M=[ם�|+�ݭ@q��ƻ@=d�%wV˫��'P�*�V�D9}-�k�p�d��!Eyu΢��D��b�K�X��ZQ j:��b��_I�󍣂(JQKc�[�])��mC�\Wu��84j�Ŝ����A`!1	�eM;}d�9���d#�S־X�h�s�eG��a��;*q���i�!(U��hMi%֐|y"n��Q�����;|��ؤ��er6����Y�e��ۭjwRT��ɷ���C"����	ʓP団�3��+:������t�N8I��.9�V��m�z�R��Z�o���YA����h�3srث|����[�Vۖhv���<��,��M��/+�]���} ����M�V��1uu����+(=|�<�8�e�w#�䱻AƂi�Y�xzXߢ��Gܱ3Qc�u,���e��(W4pT N��&��c�t���/��2�hǑ�����6K��[݆e�� �BĆ3QV��'����U��,��I|;g]	]"���w��wb0*�=m]s�F:D&�Q��fP���6�&���3�7� ��U,%Ѯ�w�@�)k�cG�Ʃ�����(wo[v�@m<���ëU^h��*6�sH"T��;?��[����9�.DE��u�KYIe3{�tg ��6��&��n�g]᫆�u���}6��d���}��q����v�W^��q/
�3�<��n�7�oo�=Ök��2>���D�t�\�R�}�LK���nɠ�u/���@�*1EEAb�����c�Y��*T1���
�&Ze
*�Z������b�K��]B���h���"��U�����E�h��d*����m��wp�4�W7RQ�nU��2k*e�UDKeT[j*�P�*4F3(T]���XPU��,Eb(�kmF�����T�\B�WmD�aEPmb�Q��\�
"*ETKu���QQ���ӂ��0��b��b��A�5EEc�TRV�QbP̢�*"��2������Tm��R:�Yl��1T�֬PX��A`���GhQb��ne�YiX�E�«K���Ȋ"�h;J��-b�F*���(���C���5���ҔUTE&��b0]`k�1���忿z����x^�ȝyN���MEY�M���;nh��Sݥў�8��o����*B�ޤrj��U,�ʞ��xx'��e���ҍ8�aE-����IF%�@<ii�$�r/b���8Q��I|�n�[]�����TU@��ba��+:��[�F7AD2Ag؈�>��f���)8*F������E�2�X�{bgٱB�\�[�坑~�O�]��zr	R�t�>�WvL�o\���qs��z��b
������	��;,����J��1~�,�*�^Q��G�q����Y��]���� q�9��r>X��]_���}B�� me����e$v�xՙ��ٚU�#���<ke��k�ӎ�(nE�}�H��V�(�su|�������8z!#�ƹ&$s��d����\b�oɚZG��Ϋ��Z|���i�S�\�G\ }��גv�/��8_D:3�/u+��iͧ���ďo��xv;J��F� "_�M��,��{��/_����p|��ihN�,M�PZ�}���1'���F������=Cse�W�4�@r��~ה�*���fL�.�I��[�5�-������eL�q�ʬ���+�U�f<�G��R�V��Nj��*��:�]V��wpޭ,�཮��:yKH��.�CVy�V�8c��˹��q)i9�v#Rك�I`᫾�l����8�+Gvn�XTnj�ّi���G�I�]����t��bNL�[��}0�v�ȣV�P��] k�ҋ���>��B5�Sn7���t��kz:�n��sy���j���|4<�9�*����4���e_/j�+���EݺEoj9�Z�ފ�ˮ<_��c�m�8��ΈJ��/�P�\�"u����W�(�I��C{�6d�r�B�(�?7l���F��u����'p�$�pt����̣��1��݈�I0��~�_u�*�t{xߝ��|��oh2�r���b�L�"GW�5�׌8�,VŅy���t~����T@�N(K��؄]�.�H��e����1�|EytR���U%̭��Aɜ��Z�8M���5�|�U���&�����uǃ�p�M��9٪�T����ɠ���:���:DkLW�2X�F��9�̐�p���l%���Q[���һ��
�9B�����2����fΈoϙۑ�eԒ�:��U�ٸ��bi�1U�,��cz��K��OqT���阆Y�33B8Md\7]�i�VU��S/�/s@Cnqֱ���{w�������B�%�AR�o����t�T���VS��Z&��x�ߓP7�6���v�rKL1p��4ʷ�b@��C|7��������F1h�K�ع��ȑ�����X��J�6��V���3�W������i��dҢ�rL�� �bF(���S�`ϋ��4�1���&�x.���s�sQ�ƶ�K9Q%6Fxs�`ΦhJS��H��j ��1��&��u�d�^c���b�9Մ#H�����N,����g\��Y/!���=�Jc*1�c��*���|��h|=ۦRw�p�tۛ�ר\����ޔS�����S��_̽���,J�;�;��������G��V�������l/�����������*z�^����QТp��#J_HE �֝��zf�Mܝ��c#³��X��OK���;�r&��ڢjn�L?(�#���8�Ft[n���N��BR�[\���$���;*�dܬ�'g������w* qu
�P�9��ް�(��,k3�m��Ǒ@��oz{Q��	�ڽl�Ve{[�]��U#Z)T�z�p�.�p�g���f�������B�}���?y�R��WM�W�_��We�r���7.l��<F��)g.4�5�L��z�$�j
�^��3ln�͊j�P�k�n0��C�Mz7�{/س=k���R�Hz���O�>Nn��ѭ�y���TL�����b}ks������w6|�齻�`���Xk��s�t2iQMeB�9U�WY+�l(�=]��|�x{�����V�֝3�"4���)dƘ%�Zc:g�B��WNY�P/b��8FZ�qGy��<a���x���=��mՙ)�1P��1�t�f7<���DU��睦KwZב�5����|et(�,)@މ(Yy(S�b����xV
Tמ�wRN����#Ac4�ƵF]�^���"�2#��,騖(wlG ܍1%��%Q�f�L�J�2]y��Տj��l��F� #}T�����|I2g�3��3��S1~j`����/z�����K\}��A�	��!Z�y��>�b�<1�{~ס�[�`�"�J�qNdM��e���iRg�o��c]A�YRFx�sd81����P�P5�n5���:SOk8��ճ9��*v"X�uy�M�a�}Pc�uɒ����͍�tN\J0�hC��^D^��������F���.#JƬVݫ��<<�����s���&��8���[;w��i�S5��p�����h
�X�S��}���4�8j�ÒC�a[��z�偊=8�݃eb����e���
\�ڣ��z���昜.����y�h�*�~6Y��T6�-��E=�Yg,�v� k�BRSD���yY����:PT�>��v%�;t�[�Xإ�`��um�O��G]mE*�WHgr�����ƽ��5[�����J5n@��Th���(��tȿk����k�0����Җ��ޖ,ƽ3G��͇�-T�W%]�to�9x�|��S���d9�k��&8R�KEZ~K{�k/jB��р{��7�pݣ~j�9������xX����Nb�m���
�u��-ׇ/wv~1�,ߵ�����$��u�cb�2kĹ���λ�f�YSk=X��r&�;��Qw�f�}K"��p{PZd	��x_�]+y�o�y��=3��=lA
��L2���"�����"�
�tEg��E	�^��ݷ�P��gk����d�(׭�үelu��6�s��b%�9"]x�5A��%']��dfU7ݞ�ApM�V��A�Px*|������ZK�U�s��
���� �oU�{ۏ�$V��'�#1J&�5b����H�1b�8;�Yw�4��`�s�+#{4�����!:�ՐFp�V���sȇ�A���m�B�"j�Ch�������NıZ9gy%B��9�f�Z��u{�mB�ڎ<�v;i�=*�9-�x�`�Uhn����6Yn��[�1�h��̼��y�	í���ҁ���}g5.�W�W,�4�
hi�IZ=ȭg���k�8'I�gPP�;n簠�r�yӆ/u-br��u�ɡ�\E4g�g\��&���ԙY��ٷ�e��[a��0ʶw�˜���atp>� JN�B�8p�� �|�!W����iޕ���R�X-�Oy�^QD�aԲ+vGC&˭sChǷ����<{*qƟH��Rh�]��6<�z�O{r�4Fzn���cx��Fl��Q�UXlk�G�F�p��k۳*x�:�A��c[[�S5s�a��j���j��詇=t�e��^�&}��U����9O�j��G�c�l�43����}�Wj���8Y�8!L#�f
�R��j�+�K�=�TMg#Q�;���=(a|�i�j]gFy�\�\�JS%Фa.B�hu���<p�e�l�y=�#UX"�XP���l���F��h3�E��N��70JGJ�LK�V;�Yŝꆸ��ќ��м�
0�7t�(u#��m�h[��s�&�X� ="GW�5��^����Yz��N\���X�؇�_�H�������n7=2��]��e�u��E�������h�?�^�XB�ιT9x�*�;cW�T��v��Y��B4$Iv���c����;�w�9����v�����t�,�����½�~�Ҝ`b��b�W��L���N4��3>����v�Aǩ�]���Y�n.�=MVX&��;v����ҥܞ\M>���%�5�8M��
�uOX�F�&��͋�Q�͈��bs��]ڹ�c�v� yy�9���v3�Ө�i�=�_�e#W �#Y��p�s�'�eYz�Sp�\?j3E�`8gO�K�aL���84ߟ3�R?�����*�3P�}W�&�R���{U��ok���]0l6gL�K,�
ff���E����N�z������tߒs�:��U�w�sd��B���
<Qq�Ș���<���#N�[�x)YFUB�sy�cA���||�MgG4xhV}=�Xϵ3Bk�Sf,}w2� �S����-<���(�:���
�/�+b.�ˍ��颅��,�G�ιQAe=��ۖ�f;ə7�J�S���s"�ώ-��c I��f�ߩ�U̠l�l"�uXr����k���|�9=<8��:'�Y��,իA)�C�1�F��!d"�-���s�O^³Y����R6�#M��#~]i��j��&�N���p�"���K������^�~LP�]N»'K�x�6h�KH�O�6�yؓm�\z��6=�&5�-��̮�N�̀P\b�R���3�fU��Il-�u`�:���b��7s���[MhK�����zd��ݐ���k8\�������q'��g����K�k#]rLE�D�ً�G��s���ݳ�dgE��ZDاHɩJ)lc�V{�c��+���g$�{N{ `O��t4t=*��U�|���M+�j}�H�3a��W-��뭸�����y��b: �.��S:lfU#q-Oy!�C6Q�-�q�eWT=�[�婎��7F\EC�BP�q�@�o��>,U�yh��x\���]���A���}�����¥N�2�28��	x��L
��i����t�ӖxT�1��9�x h�v�z�U�*u�����n�ȱN����@f|���P;��گ���b.l�C�џYj�f)��\�/X5M���h�oŗ�"\��U�,�"���fЋV1�]��0�}��UN:�Uk��(P���PJF��Q&e ���KI= ��5�{��-
��x�)h��fR5����&�x�I��S1mL��E'��Z/P5ko.j+�M��^ZMs�q⚂�Y�x�Y"�嫇���4mN���=�V��޻'~Q�i=�ًH+��1�[�N;��(�3��q����<�{��V��7�Jx�k<=x���3�=pQ��V��N�;ȧrZ��w���k�`��\NdY�`�t{5_}
��n��MR��&Sc
����C�+�5����éʳND0��Ȧ�jyrENl���-�\��
��4�Pvg�
Х�"�p�\r��]]����ey��͛��;W\�-��<`����D�sH@�i1p7q����&��j3��B�](�+\��ZD�n���k�4�v��^݀�[����;���m滙��"��"M�4cA\��ڱ���ͽu�Uf
qȺlP/��bIq�S�ш_'�X��J�>ʣ/�F�+KȰQFG+�E�k��Y�@Sf`��e^2��ޗ�K�Q{��\�:/ʨ,��tZ�C�Bԣv9�4V�E�����Jc]�U^��lc�Q�k��Ըnѿ5X��ϗ=%�},�1J"�ӗ[�@�Qɣcm��:Vi~�;ЎޖoX�1Oj���L���-<����ɕ�Kn�{۴	PrΞԑ��SjR�[��z�C,߃}K"��sڀx�� O�q�#L��m�et��X��c�H�f�E��f��w�s��uEgU7�r(���(�pAfB�8IC&�E.�z�΅H���-����w�1�g��XVT��hA4�/bM��5��
��_(��b��q��bꤍ�q��p-����`a�\�Ƕ2����n*J�K�S"���1Nk����d��h��CP��Y�e�Sy}Hgr��d����ٍ�����6*�zgJ�l���3��.��U��r�Ⱥw�t��LD��fTYt�jXn�w[�@i)�z��|�O�A�?#g�b�|�h�)��U����� ���m���;&9f)Q��r�����S�s���#�Ŋ����E�~�@�7��rv���ơB��9���^~��=ZB8;�>U��
��#�
�[��.ג�����c+�_�"{i�&�qџA��I��&<6x���Y����y��On悏�b�	�;�`�~w4�a����. JN�C6l�OQ*�D�ԯ���0���};�o�^��?00?�^��U�?�Aγ�ՈZ1�W/�9��S�ƟF�ٗn�x7rg�x��b�
�'^n�Y���mu�ϫ�Q�UXo^R=��*�<V��he�5��Y����9��a���v,�뢦O]:�q�����ef��U;+���fv�.�$t�<�������,�7b�ϣJ��g�h��Go0W�C�|�Dg��yk،�!�b{V��fG��ӥoӔ�Eg�SL�3���c�XYNݣ�`qR�\�)�f�S(X-u�{�ż�ML�b����ѱ�],�����XmN�<8i[�Sү60i	�>_
WR���{:J��{l��q�f�ٛv����̷8��R�F�7�ՠ��'�h�kk.nM֝<3�6�W<��]�Bг�Q�`�gs�(�m�)�1�,Z����]�*�<۝�뷔΢����b�[�:(N��V�3#��|��:{:��ʖ�|ջa�d�M`�d�Zә�Z]<&���]��T�9���d����(^�:}u��Uꇹ�v�'�x�L�J8kpqp��b�J,��s��	{������l��֬Ğ]�f��ZI�3�Zd�d�j�e;�o��;�/��2�E+���j\4d�O���[4��Z�\Ho#+0�w�p���^�9�U҉�o
ꌲ��C���f:�U��$h�t�����S�v܊�aG��Y[��ݞ����.N�rٓ9���d0ܵP��Y̼��`"����:��}Ϸl�*��(0�P��u��P�l�f�����)8Z����o)	�ׇZ��j*�J�����f���C�����ܫyW��4�{f+��u��5�wD�@��[�.&���~�`�w���[W[]»�s�a���j9���e@9��]�r�����A��νp��eRר�0��n���qbʵ1+47�,V�o� �E�S;=��~��i�vl8\�BVr�O�Ӽ�7n�J��m02���rm�v5�iu�+f�a�t�#�U��׊h���5��lK�:�xt�ݷ�h�ﴙڡN�%bͩ�z��֭���c^�p�gOE�e�f�:O��2WV��yL���	8Y��G�5��7cZ�>��bJIp+w"��T����N�jfp��n6q3^g%�~���x�ؔ���@q˝S��]�Y�!�8��rX�<�\��k����]��84>�;�)t�6�(>rP���avq\�t��)��
��D�`�!�jS�VW>�{��(F��%kٺ�v!���NWCJ$��u���NgY�l)���}S\�f8��i5n��0��72��&�ײ;ϋj�H��k&E��5iL�d�B2���$W֩��qi�6v#:��+����\{䎓VM��L,SQ��8e�b��;��;A���!���,�����!��o&V�b�Godg��n���
L{b�{���w�����P���"2�Z]��Q�wS:K�+�]�Z`�M>��%�`ۥ<_+���a=8��j}b7t��3N���������<��a���ͤ�N�ޤ��!����VY)�+�ͫZ����Z=�}cl�7�F���Q^�&
w7�s:{l��ٶq�(�|C���M�%U����T�6�%6���-�_wZ�]0��:�N�*��)tdț5
�AA���b+"�AX�X(��U��-��lX�<B�R���ƶ�S,�J�h�"�U��H�*UAUեAdDPF
��B��F#1�Y�Ŋ�,v�۸TQH�T̹J��%V�qT�r"��Ȣ�e`���5�m9eb��(�Ԣ�ܪ��`� �qDTD�F"����Y(0b���S-Q��ĩ
�Xk1�Q��M��(��Kh��U������UU(�������*)�j
b��*Ȳ�UV;@�+QT��-F1A`�UAQ\eb,2Ոł��`*�Q�X��
"�TX#
�D�� cEֳڗz9`��.�M����W�c��"�Zr��o�čN�b�./#�˒Ӯ�D+���1��\ 3Z/8��ӻ�-\>�{p��o���(Q�s{6�Vz�30�IDt)N�9�]�°�q2kq�guk3k2d�~p���U��l�Q�ڝ�αzx'pᛘ%=*��w������L�~��+n��gfĩ뇱�}�a{!�nyd�{X�/H��y�Ι�3+*R�W@�����ϫ�r�������ɔ^E�t�@��e�:�r#�gՕ��V��o�p�s4W�)������{N�P�`Y]��د	S��<-U=}p�mZ�ԍl�8p�](�&��f(&f�����O��i�+�xe�\2x]�����0�'M�lJ�֚Y�&/a�f�Ux�`��/�,��|͝ߟ3������")�G�P!696��d�Q2�Uz����m��0�20)�!��Y�ls$��^=cF����L�O���^]2�d��$A����\F�1�1^Nɂ@f�:�$�O>;O4+�X��c[�|w�=�,�sE��F<�3��ISf,�빟BEa�ʿe��P�U�J��4U��,Zק�'�������|�R9����9�]���u��{:�>�)N�������+�{z��'��w�����[�;�܂.e�k n�֔z�[I��ȦZ�����.#@iu#wժ�꽛}��8�۸b�xU�z��V"�(.����:�b�����.%+��\6��Em>��@�z�jK���l^���7�2��8i
����u�7��߷�b�ݹ��ދ��po9
u���m,�q��ئ�L?�0}l��y������������tC�*5m�_s�UQ�z!��\RUH�9�4�n�6�֝��L�n�鱱Ǝ��D598��ĉ�zk]��o*:E#��h�:�C��:E�23��u�M�N��	D��w�"��6x�u��A(��QUhO�DQ��䢮/����z��(��5�Ә��R�(��OQ�h�)�XVԔ�4\9}1U3��̪F�2��Y��F��q$�k��W4��зEdaa�,��P�N��
G���+#.e�"�� �
��\��Z��Y�T���K�Чi/�/)�6f�28�Zd��NX������Q�:�'��ݑ����ν���rwR�DwC�,���������}VdOҌ@e,3�t�f7�cU�Tu:ϼ��,���t<�)���i�"�&b�ؤ&��A͑R�y{տ!�%Q�t���e�b�,ך�M�z�Fwk�[�-sqmh�ji�O�#ӫ'F:oVw1.��qՏw7�&�4����p���'n�k�[����ɮ�a)'k�<d]�RU�>���d��B��5M��SE�~,�������*��1��S+�i�m�^��NqC��K,�%�6������o�<ċ�[m��R�q	���t>�{��$��Z�uF�RfϟG�&��5c2��ܦV{��29g!�e����x��Z�d��1�a`�{��Ɋ�K�?8k�0WH�:�Z�}�ס��$<Ƒ;OvN\����ޔ�եD_�3�~j�ħ�$QD��pc�FE����V:��&:H�Ba��r�W�"�	K��y^dPo+V�5uI��,b���J�h
Z�=Y�p�ij�§s�%G�7��X/R�|��|�W�1�m֘5�}&��U#B�O���>1bqʻ7��#�e�p^Jf/�iS�S@c�C4)
���^ٰ�0ى��;�q�ѕ�8q0��*�o<�6oقxз M�����/"�E�tȱ�^�D����"�#0��0�o����:M{�v��LeO���7(������VN\$�>�[�����J�o��MdBIZ�VMo�oq�v�jv�g����ܯvN�EH�{�ҭ��i6�`�@J��,������G�qز��w-����J.\�^i4��Q�,t�'���|;���#�V#���+���Wan�����oL�������Y�˲:��O0�{a��9�lC,��z��Z��7�������*?v[���Q�K�W/*4����B8oK65������C#�2:]v��(쫴�w�ij�}�7�;����5^�d�s�\�+6��y!�o����X��Hj�Ai�'Ÿ�zY���A�4�}�^Q�����K:&^��"�26��ۍ�Q�M�Q�b����=��Z�[��&x��F\��P�B��7�4��{bgٱB�^�،坑����<ETn�HJ�Ժnj�İѧY>���ЅJo��B�П���]�l�A���M7s�I.���!�gf��y�/����hS����������j�7R��2�{2b��.N�[��Y����IIn�AH� o�3�a:fuVܗ~*MG�vl�@g&��;��\:j�d���q|��j�yC�c8H�R����яA�rLO:ɆO�<����B���*+tOkM�)����M_��F/D0}�@�	;q�
L�ce�����=$S�U����
j���o�N��8�XM��.��������Mt���F�$4� �Cd+=H�D"^�kZ�p�㕜H�~S������}VxZ�Þ4�yb��z&��}�G���	am�vj��f#m�j���':j�.��IL��I�Q�N��B�Y�!@d�U�ha����yƝ�������Lĉ�nj�����]�Rk�̍�u�o��-Π��|�[6v�����c,V�~C����Im�|�e�:`��g9��یO(Y��#�e}���>�{y��ndtbjJ�����5){��7b�[�D��NX�xֈ�*�w,O�
R�W�iWE�ز:]�]��ȝ�~JY�B29H⍁��:1�[����Q�hp�w�`ʸ]�4��X������[���V1�g�C ;Sc!w���z��h3cX�=6w�&	@�]vbx:�����g>�/Lb~�fpf�����������ܵ3\([���,��b�H�3�0��ye��S\kA�8�i�}�re�	S��e�at����2�F�1H*������Fw]����\D��dF��_&����F�'��t5�0�\��ǅ���;��狱�0!�ϗ
 4�������q�WR:2l;�v����Q�
�L�畿p����Ş�u�� ��6��{���\r&[@ լ�[
'��pz��D��x��V5���M{/�n�g%}���D��=�3�x�t�#�tϕ�u�2��]nSu�pާ��I�"ŧI^qYח�Zg���屝R޴�*��:����y9[�Z��ݞW�tPE��gh�������:}R嘠TT+�FG�c�W�+Kv�� e������h�r�����D�N�@�`��.�63�b�D�L�ЎY��ͨ9��tfv����v>��eb+�tB�cb�(��LdL'D�k��x+E�%�]�Љ��OXrgM��3�=�(ײ�8l��3��ISf79�x;�M�`o�r��՜}w2ƹ�;��+�^`�6�R����҇U�<WG��HWZS�J���v��g9aJ����[��7\{"�Џ�=�c�F��NlK�/��P��z�'b�����>�~o���W��+�l��~YH�]��_y`[Z���C��=(�׺L.e��b-�o2���׫��Ŀ���es�i��l=u�j�a��I��8�Ң�S��u��Չ��n�a�rO3o�#��u���5�V�
dgE�ͺ�&��2m���]���ܜ��n`�9����WE�*���cG��W(��q��a`
%�Y��:�r:t����<R�<NuX�k�<X�'7����h����L�mg�ėv�J5Y�1�:����a5ZTI�0p+!	sog��ˏ
�R��M���6eM3�\"������W�nh��m�g`����V]�wq����uj�7[����B�e�P�`�hGJ�ўuL�fU#s��i�"�+ٲ��,>^���G�.~�@�Q��]I~�d�:�]�z�<�E���9Uv�����삘������bS�o{�j�u�L�r��dqL�,����Z-ULϑ��틦��31�S����ڬ�U8X���Z�l+�q��Y�b�#22���\�ٌ��o�e���gI]��'�Q��>�g(,��6�����h�l�ȑT阥U��$x�S���iNW�g
b��C�7l���2Y�Fx���ȇ[,�0ċ�q��XnF��
�b[�9jZ�"z����쌈n�S9(� �#lMS8j�̤k7)���&L�r ��C$�=�<u;�מ,g�\�U���0d�܈����\�����+�_K5�)�����Z��Q����X~���|�P�:�}ԋ��ќȫj�Ą����!����ȼ�4[�J{\�K\�;��oM��x[�����K���y�^�aZ���}^�=�бI�״�E�נ_E��6>מT>8��Ŵ��
@�Pt�Ң̽�g(�sN�{h-2:f#[�z��5_"թB�B�toWWE�%i|���̝�o6]�x5�,z�����]|�_Pd���{7eY�mX]���u��A��Ϩ�9��eh�5��#�_ѐ�k�z�DqZ�Y��J֘45�T�JZC(����;5:�S(�R0�5p�2�b�T�r��;V7<�+s~z��<0b�9T�T�3�#W7&	L43*�o�F͌�<j܁"�QQc+KȲ�29]2.���S�:��,���rt՞�uwV%BkҔZ��K�GE���ȱ�'�z�x�|��N�.Do��qԋ���{�GJ�,����8�%C,�%R�^��v��y���F�b�ۜ}�:�C�s�܄�GI��dU�\�z�oK:�q�j�Gdt��1�ٔy�5kv|�p�����C-���D��G��-�s졛H��Y���E8%� �eP����"�'�9e�h����*�,���0GVΉ�^X���v�h�"�
�Q��Ή&�fsXrh�Ǹœ�<��4ׅ�L�x����;+侼,C�hrUlF���d�\c�s��ov���N�N�2�r#j�q�,U*��<q�=>ń�?��F}�E$���V}�E����.�����.�`M�NG)àcB}��(t�'ϯJ˚1��sw��M�F�6�Qvu�RA����Gp1��Xo/�β�\2�.�Q��nPKnG�>������3��3$�����3�	X�B�>��ifZw�z3�A%�GRWiSp����d�,����/�i��|��^�J���ԏ�C(��+n>���le�����Ԛ�
FZ3�a:ft*ے1ĸy<@g&���]��7��!57
Qwr�4�c"}��2ht"�)�>�#\��&���ƥ�RQ��ywY���x��*�v|Q�z���T�P��ڥ�	Iӈ�8Ç��0zV �Ni}��pQ1��!=����oR�tк�E�!^ɲ�k�l�uKm��J�KԳ�y���w���!#V,}��-S�V����6����Pu{,��4�\��ͷ}�[�JU=x��*Tb6�#���2g|9Θ�C�hc�뜆٤����]C*�p�>�^W�)/�³Y}�ia)���}�:�v*ź�JJ��g�h�
��f
���9��o���,��"���Ã�U�4֊����+��)���4T�����qb��&C.EOa�ILn�2���ۙ@����E]��ބx)���bx߯�s��佘��c��q⻧��uoI�,���W�gw����{6]��oWM�K�&C�ƬIչ+�
.+,�D�ܥ������(XMN�﵁5��!�L��hۗ}�3]�"�6+ht��újSt���݃gu=P���wY�z���u���m<�}�%႙:.�G�.[��PͰ�����M.3���=�jn>AUm��,�HT5��k�90�9pc�t�m���z̪�_X���s:b�f+�X�����\nDX�r�>"}�Z����_F�g�8�V #>����Ƽ&���f�c���u�{�]Į�!�Q����� ������i��u(�T���<�R��Ǝ���\�qT]\=L��@1R��;@Է9��e�>�r�R���|�28،t�8����]'�Lt�L5v0�0܌��������~��1A�d(�!�;��"�왾7I��=C/!��Kc�������ʖ^��Lϱ
g�<<N{����0m*��&q��yo�3�#�K�V�)�b�ҫ||��p[x<�0s�`ΦhN/	T����OBe�O*��}w2�A��rkő�as�Մ#H�n^��
�VipFq��졘���^�۝��YKa�n��Ed#�Ǳbk�F��^p3nn���@��<�����)3�~``	�>ll���mr��;/6�D�j.���W��4��6�Hc���w��Cy��y�v��:�;���+�\E�֭���z̏5�7���W
t�ɽ�%֖";���]�e8B�8Ŭ��n�2#O>X�E�#���+~Yb�J�v����M��Z��*�t�y�F�#��qT��*��B"_Y}&�O�L��u�d2�&:M�G��[ZM��n���>�wt���eN�����d���Gu�����:��ɚR^ۭ��朏�
��¸��,\;��;ĭ�O.��{�\/9��t^PB����$֐�X��̊��*`p��j�Oz�YF��Kx�Mjnv��ۤ�R�L˵5RivP*����>WYG
� ��ܻ��n_TIdT�9.�%=)F�W��V��=����P��SFu9[�v	�v�B��ծϪ�4S�Me�o^(�r�����D�q���9�k�yX�Gc�R�V%�9`���:�^^�6��-2�bbwa�T�/���%��i��Ǧ��t.����GG�mԱľ�X�.����23��R�<^��{3Zr41$`ivl���m܀�Ii�N�+a�Ĭ띍�9�oe��ԯ{�;O`�� ��` ^r�x��R�A�"�ssT�"�*Ȕr����$V:�QR��JЬ����t''�������s��k#σ�:��8]�ً]4��Ór�M	����_c����-�N ܐmL�U�ê�әf+t{���lN�G
zT�ʎX�#���t��ۦ�Z�^�s�癇K�@/w�=\�Hh1*��sN�f\�3J�W����T��}{�6�fs�z��҈l�}5ة}r�z&s�)Xu\�"NT-�ႎ��-X��[�5�˖���tM;�{���]cAu>�ޮ��N�	'k�Q��*�[�7/u���M�+rJ��4ڡ����-fv<+Ir��/T�fQi�N<���E�ћ��B�]t<'%D��`N�U{5n$�1g=4���C5#A:�Z@���vUh�^���+o_R8*v�w�	�`X�ei�쎰릺t�Cw�[�땀͇���vt�8�Z�2��ܬ𐱪$����3u�.�U{�f^�Vp*�%_3d�9�z�\7��˱�]�x+v����ã��3m��&�U���I�M�we>��緈P'���\�E�4�ڰ�1$�a3�1�3}�:��#/֪�R�b�鳳�<����uՔ�2���r�����]��ʴT4�wI3�(S�Ai����n��P^�*��FFgR L��.�5#���V8�������b��	��5��J*��F�f�&�_$�a��ڬ�ۼ�0T��kR��]�'+���A7�#�7s�Ve:epGD���b��_pFnr��e�*`�0��U��[�N1�����Oz)���};���f�\�u�}��.�út�JjE�.���^�=��C��:n�Ѕ�>|J>fA$1�5ԣ+'��R嘨�@U��H��"��*
�j��F�+4q��� �EIZ�b��U6�B�V�m���12�X��Q�
*F�q"����������DU5��Tڍ�bc�Ev؉��*��2�]HSm�EPb�\�A���嘊�#�.R�7(:�j�T�DUT�1���l���fTJ�eK[D`��sp�nچbRcR���Փ��m��Y*,�a�Z���3j�Z�f2�CkI����h��E�Sr���#��J�5��J��&&m4H��]dp��hX*��"�"�lU�;Q���X*���c1�Tm��FTTUF,����ܦ55�AE���K"��rɬ*AU��FF�j��\�uGi��a�j���WDS]���h�G�����Jp�lLv��y�w��.�Wp$w���Ø��
q�˦�&8˥��uXo��唎8�.����q�����l�q�
�M�4�i1����w���(�C*"�F��ʩ��a�Az�N�Z�3I���ʍ�)Vj-�+3��N�fʘ���4R0&�R1�δr��{��g�΋�ZD�4jas�[l���yx�<���7��Ք8c�*�
�)�<]¿�UŌs��a�+og�=VJO7g�zV��@zČs6�z�@ף�th���c2�`qjxۀ���q��!�s1�Ό��L��Ӌ'H�3a��zD�Nc�!
G���+"��T�8�;|���e��ETT���,�Ɣg՝L��:F��28�i�Zɍ07��-1��}��c��+NT���ۍ���)��[�r�^�	S�k�t=P�`�Y�.Q��@ea���z�*�Ќ���ݳ�yjn0���`Y\�{`P�#6�j���$�x��$P�L�[�9�e߃Lc�>�uٸ*
b�[�`ĉ<Y���pSV���<�co=[[RlF[�-��Vn�1׹��֨v!�˹U��u�	ٚ�x1<�"�GB޶���}�Ãv��t�}%���$y6q�ޏ$�m��:1�d"�t�BI������M�)ѧqn_N��GY���]�f��/�~�w��.>��8����{���3:��JB���^�ɣ^�U�()�x謟&�Xr��uyoïP+�
^��������K�><{�,o�b�n`옠��'�r :=&�n��_K3���E��W����秢�^��WG���!)�\F��7e�s ���)��/? ��J�K������g��֥�.���;�7d>�8kc �'{������E7��+\�j�&����&�9vcu�Bb�u��Բ�H��b��sL@����!���w�t�8��ZBܜ"t7Z`�m�nJﭽ�6�\�D�ؙ,�W�:�7c�al�N^Jf,�+�H�ՍP9�6�[U�\�Sӫ�+�ݞ��B���XCW��U�� �U�i�Ua�ì��<��4���o��^f�z\������dnp8���j�ԥ�2\�:�W���9�ĺ�_p�����p׈R�wC�.M4�n��V��<�<9��~�Y)L��K���U���o������s��q"獭V���"��+����r�*�,��9�ABI�s�c�c05�+g�MZcv�L���uLHA�/�𵺡9QI��g���v�P�}t�Y��C��r2����:���$��L�I�1	�qqPVWk�9���\��R��je�Nᵛ9g��R��Q�e>S=Y����8{�]���o{J�JGݳ�rۜ;�%5�T�%O[��>�ͤh^He��U�'$�����w(�Z!VԵ��3��z�d6,�/�K�c����kf(�]�EgU7nEL��Ѐ��0a<�8��td�������w�EM��8k�.Q�1�d<�@L�6(C�qVz����)����[�ٽ�պ"z����L�^��%U7�
��>�PhO��썈fx�KS1���{�����b,���d"h%_�)�1J�׫����@gV&�|n�|3õ^���^N�O{���� ��1y�%��`�H� SFp����:�W����V�/�6�S�{J��Ѳ�!��f4q�aPfn2�u���!+0d��E�PhϠι&$s��g2VuX�[5N�SZ��6X�3���ٷ�e���#F^��R��Iۈ�aÄ̈��U�b��;z�8�{uB�R�2��uyc*5�[�:=�ek�p�zw���xIhݡ*x8�G���"�U^�>ϩ�^���)����FS�\ra�f�>�����P��NLz�q��.��P�n��P�N]��-��Ve�;�͖D��7�����CQ�r�+�pWTb�c������f��sFdڷMtc���]	گEM�S�z�^E% ����z��B�Pc�ގ���fsQ���[�K.23�P�E�J�N�������Ħ�`.��ՇU~Gb�oO]P�@���^^��!��%�K��RTB��JB:��cr�g\n�]��O�W'.< �W�|dQ��q`��{��ۅT��Q�|�D^)gtr���u�ۮqX.C%)��:h��[�w�q�<�r��(����s+�
 ;S~�E]��)F�#jv�7�N�Ntd�x�W��^�Z�p退%ys�����Q���*�-�׋�W��:���9�it�I�V�R��ݚHωoH�ԙ��8�cb�����t�m��K���4�h!OI���J���c�.cL�ܣ�+�lFy�i�n�����x���K�q;T{z�r���ж�,(F�7NQL)f1!����
R:2]C9cTZ�c#��B��s7��#��\#C2G,��5-����,��p�`UQP��͝��]����6}罜zٜ�����.�#X��k#"��h0X"{����阯:�]Ⱦ7�=��W'Öe M���=���ڊ�>z�ٍk�0*vf�۶.�b��犧+�7���F��q�:�K3t'��K��[e��n���X�c�fB=�y84�d�1M��%�m'�u �
H��-6#��r.�S�yq���X���꙽}�IL���F�c�G�<0�^��q�c�u�ו,�$�!"�lP���dEns����;kzb�a��`ϋ�h����0R�-SY�i��U�S����������l��,)ZP�U��g�S9��$rȹ4#6�,�6r�˦�����@��"Z}kލ�����=��&�S�mΝ���#�ŉ�ʣ`I�8�6<5�)�i���ʣ���}�Q�����ҍ��@Dm ���uwE`n��t�����\�9n�&o.�V�ơ����6�`#�5�2q25G)�ts�#KnB/ط�0/G�i��ê��=�i���:T�"�	å3E��b�<���<��<�΂1����o�S7��BZ�!���o�?86��qUh_>ZM x��y(���.Z���/3$����]��^ ���k3�ly��W�LGJ�ю��7�ʤn`q-Oq�q�!MZ<���a煮��K9�^��CW�ܳV������<b��C��B
��	�ĺ�ĸ/�U��ϧ��E�ݻ��$�뢄�k�-�5х�4��<�f��D�����g:����C0�VmԈc��ĸp��5Xw��0{r�{h�z���w^��M�V���*�K�8w'�Ϋ��O��b�2��7�A@�&n�q��v�e[xz7��$�v�W��;*�|+����X�(ϫ:�r�3����%�YQ�7+�/D���yc7���K��NQ�Tء*p��,����n�ȱN���М�2c:�q��Px2w~z������bl+�R�;��f�5M��SE�~,��rz�EmD@��[�Yq�����6di*]q�m�d:6��Y�|��W��>��E�^ܞ��5!�<wpC	H�BQ

�a�	�()�x謟&�Xr��w��t�%���A�}Wn&I������,wLņ�Ɋ	ϡFD�=&�l)3�Ȱ[�"�w(刈Qk.* >T�I���r���ޤF����<O���A��yr|�͑�rg��;Ko�M�r
��=����J7���Aٞ/=J�(q��y�A��9X���ɢ�������'f-�Р);^�{@Zsz�W��P���v5҈���'�92�t��ݸ��f�vL�����F�Κ�F�p�7����T���x��<G~t�W�����߻MNpCKq��qs[9�][i\�u�.�{^�%]�'�F݊���5PX��Y���3k1�)˰t�N�n��u�eΥ���<�F"ӼI�Y�%̖x��e��}��n��ye���T����W}��\"lC����'|î��>����5���3=q���9b8�f�m`�#NM�R����7��5p��z�HJ)N;�.��4%(����Q�~��Ϯ�hs����I����ܣV�Nn�j�#�C)f��R5�8�Q/c�8�K(�J��t�=�1ԍ.#�7������k���<�����W����Q/eq��ޖu������$�txOC(��	�Y�ʹ�\���Ѳ�?�<�Q��j���uxѡy!�m���Y��b��jc�l�u+����n ;� e��cb���8Q��gf^��"�24Vu�q�������ʚQ�ׂ�Ά�WA�Xg`�����^5�bS<.`X:b��}xo�$�܍Y�]�}�?�e*?�꿄`�,��;�3��Pj	؉�:d�J���~F�z7�ޜ5Q��gm�{��p��\a1C�25䩝��r�R�5��f(Mxj�*Nu�t䝉�l����Q�y�6C:k2b��:�C�X42��ќ3�f�m�v
�QǬK2c����/=^�`c#���NT:��"�� ��%K
K0�Tkn6�d�n!�kR�X��v�1f��)؇P�5��+j6.��� b�Rk����%vr�����w��V�,�f�0M�����¢ޥ'N��n�v�F�UݯS5�i�Z7"��P���"(c���B."�F}@�$��J\S�nbZrs�37�1��*E��q�)׳leYf��4�a���5K�A'n#o�p�dN���q��-W�l�~�0HWȂu+�+�,Ӷ���Ƽ)�*��9��N�[�x��gv�W.�~�j���m�����=���X�v2ͷ����Fl�p�������a�6x��V����iW�����8��a��c�v�T	:-��w9���vRe�M<�{�KvR��xq7��o�py�8��t��q�v��>I\���b�r�^���y6=���cY��%��;�J"��Y�R��;�Yэ������P����LY�_^y�!��r�%��G*�hu�����NU[�C�Q�߂��Η�2��ח�:��W��뭰�ܶ�:�J �U�׳(�N��8Ͻ��y+������7z�>Z�a�����r�M`|k���$k������|�U��Ů[g=���w�+�A�J�ZM�=��!Q]�6m�j�y�/c�=Kt�r�`/�̉���t�F������Z�"�:�����Xsx�3��i��i��6��6L����́WY�ted�
2��+:�>��e���r�Z�;[�'W\�e�YC䄥�[�̓���Vu2�M1r�S�+Ұ��W�K�،0�MX���9�6��J��^V��{�{���R6Ǡ3n(K�رY��,�9DA5*���H{�`P��ђ�U�����i�w(=<�0�V� �q���,�����Fh�m�:}�UQP�l�7������y�92�\qp�*��w^Ⱥ��fB5�ddTױ��x�`�����c/�����x���`m�vņU���"�:��'f��;�8�c��|�]2�	�BD�6(p����b��ǛI�Ƅ�f�s9Y0B���4��	w����7��;��	f�7�b=KB�f�R���Ul(&+2%�Rf/Ǉ�$�������<*� �U���Q�z�NS�edY�=X��_O q,�+�)��(���*"h,�����Ȭ��=.��g!�W�,@˼젳ʠ�����q{Fy���q����I�a�tF��Gb�����0}l�OlL>��ԋ���«5T��<:�͡�B.#��3�\Y[n�6�ӵ�
^w~��_�l�x�(���Վ)J�N��Y�$b��m����9,�����wr�%�J84(�����
w��<�m��)i$�u$���q���2k�.��;˃��3Z=A�-f�Z�\u��W6��:��w(2�sS����G;��f����c�a��	�qw$�S0/�#|�+�L�^ʨP{�-���ݢn��"n�#&�(����Y�D�v�r�)���Y���]����{p��IA�]��6�`�{X�}3͇B�L{�WF��g�Kw����%�{Zb�<�9=W�rM���P͔k�g��(�ͅ�x��#���!
G��l����rt`ԉ�w�5������T%e�ɲ(B�F�P���(��L�r��dq��.���L
T��%��t9$�`����h\�����wJY�P/b�N��p�CqM�:F&���}�6]���3�楇&�X	؊�u������8} W��%�
�#6�Sp9D�	�3�jP�7���ݧ�$?S�b��*�#}R��O�~K ��Vҵw�y����I!�sLV�_2��%!��b,7#LD2F*5L��0�q(٬�e#C7)� v0r��e�k���9pN���+O n���v�-�y|Wժɮ�!d��M+*�I�z���B{�$��
��@A_8������A��K�ˀ����.�Oe���ti	$ I�P�*�ĺ�����ɳ:�O�⬑z�1�Soa�d� ���jhڭI^���"��x�\-�1��=� ��ٿ�G�a
`DV�� ����7�Ѡ~�΀���{&��3��G@W��z�z�I�IC�<��%-󍡚y�e�g�qv���h��ԡ%PW@�_�ۗ��؉��z�@ I0�*0�5�x���� ���47>�'��O3�&�=9ɱ@��y#T?p���?AV���	pj��&;I���t��{c����B|���:�5UtM�%v�?VDڇ�	�ʻ��PA]@A_G�\*��L���!�}�@�$�4�`
D��?�p�� D�P�0;.�c6��!a|X��RB��X���h]�P��+��aچ�PV&>����`�#����W�oÐn��$F����z'�C�h��lI|>$�@A^g��]��ܩuG���J� ���T��{���;��d�FF�<zL�,��i�[�4�ÓS��������b�+�����Ky�rc�ʥ�*Aa�ӄ�^�y�	�Q1�h"+�)Z�����3}ق ��&��`+
�4<�:�� ~G��kW�����)��q̀i/�(,����s�����(���	���`Ld0 �  �4�&C 0L  ��H�D� h  @��O)��F�z� F�R!3BzT�3U�z�CLGꊧ��3\P���?D��J�h���(���U6����L@@1�05�3gc_o5�+ai�0]	��<��j�,T�!��Cx���2T��m-0����n3�o��g~R�FӘ�!�с�2$P��{�@�1t��,�k���'Q��T�h�3!��`1��n�Bt�J�錤�t�4���-��opH�V�m��!�(7���ҽ�$����QK7I�hV�Fo�I,�Y��(�`�a�H`AʌLCw>7e�~[ƃ���t�(H�r�BB�2ֆ�6tNnЁ�`H6�:��/偼��I�C����c�����ι��F��F��B˚@�S�]���L����g3�8Vm<KQ�1���CYl��6�/����~�NH������E�2��ī#�D���**(V����j�f"�`+o������$t~� �=8�1M���/C�Sԇ�N�	�qm��CB���N�`t��58\%�~;�t�,z�C��3��\�윃!!'�'z�יX�p1I��L4�������@���f��	CY(�o�K�
��N��W�Ln�E�J;YZ�!KC�"P�T�D7G̩yP��\��3�?&�.�;������;�jBb<��?r��<�#�0�����?C�,���q�f�v����l��٨���H�K�� |x!���q-' ����Ч)��٩%���>
n��ǆ��E�y .����Ff�����v�1�唆�o�2X+ul+�����.�p� �4Z�