BZh91AY&SY�Еiڽ_�`p���"� ����bK���        ��(*���A�R�%T�@E$�HPU"R�A�J%�A��JHUEJ	"�E)R{b�*�J��*�U��D%*J������EQJ�*%R��T�*	%UR�R��QH�( r�yʤ�R�<L�ID+"�T�d�(�Eb4�RQU%�Ԕ�*�:������JIJ�LP��BDD�*R
���� ��T�   
- �-����H�m�
 h�"ڕ@P�A��*4�ISl 5�(5�ɁaZ,�*����BP�(�   ��Р f�4  3L  :��@I�  �.�����  h;U`����  :]�P ��"J���"!RDIE�  i�� ]G8  t�( ��Pv�� A�s�@P��:tҀ�8� �7  t��  nT��J�%
��I   �@t3Kt  ¹� ��  :{<^y�P C��(pNp��9�  n.p҂�W[9� ꆨ�IR@
�TRUR�  i�  Ўs�� !��J��[�  7�t ;)�dP8@�.\� ���  �� 4 \R(�B*�R�B)p   ���@ �7G@ �\�t�ia�  �;�PU 9�p t�k�  ���� ;���5X�p ��B�IB�
���8   ��  ��  t;F Y,Q�A�X5@  cX
�`���p t�� tjD�)*��R����*\   ��N�  ��  ZL 
f�A0� il�T3  �sJ Q��JT"��@�G  
1p �2� !  �` ���Fр�` �C` h� 1`��& RT)	J�UP��   NP9� UwU��
��j, 5� Q� @5�Q�h�   �   �� �%R�@`� #Oh�JU5@ �@    �)���hL�O�M=C'�M��D�AIQT`    L	��&��A�   	4��P�R0    V���y,�1;�BCD����^p�ABJN<��':�~���! $�>���$�TSR ��Ԫ *�f�k��벧� U��LDDDz` �*��}B?Qk�~���S����U���u�,.,&,,.,3���������C���'c&�'c'c'bN�Nćc'c'c'c��N��N���ćbc�!�ɑē�	��v$;��ñ�!ؐ�@�Hv$;�bc%��Hv0;;����!���`v$�a��v0;�M�C���@�`v v v v2v$;{;;;;���N�bb��N���NćbC����������FN�c'c���d;;v02vP;;��"c����R����@�Hv07�����bn0�`v$;��N�!��"N���bc'"c���v v v2v0;9N�bbbc����� X��d�`v0;���bc�c'c'bc'c'c����%��bc'bc���ؐ�d:Fb��؄�I;��c���bc��؁���@�d�I،@�Hv$�@�@�d�@�@�@�@�e�ćc��!ؐ�`};�,gc�������`v2}��c����؁��$;�NćbC�$�Bv!;r2v$�C#!���Hv0;5��v2C���n0$�0}>�!�H���a }�; v0�;$ĒbBcC� ��Br$ v2;�!20�؀�!!�� v$v Hr �d�;H�$�$�&�!�C��!؄��HBv ;BC�����HHv! v2B�!�B#	��@�d�;;	����������dn$�;B���BC��Hv �HHv2ѐ� ���'cC�c	���Iv2B���I��$bI���ؐ!ؒ@�I v0v!$;;��,`@�av!v0�;;;HD	���c �Iؐ��HBv$!;v2@��$�b'c	$�Iv0��d$�d$;;v$��!Đ'c	$�@���v2; ��Đ;# v2@;�;H���� NĐ�c I����K;$;;v v2v2};;;2=��ćbC���d�d�d�@�@�I��$�IؐȐ�d�I�����d�`v2�#'bN�Nĝ���;���;;v$��d�I؁؁ؓ���'c'bbN��N�'c&D�ĝ��c����ñ�d�d�@�`v v$;����ćc#���N�b#�����D;��������N��7����؁����؁������؁���I��$�I�ñ����Iؓ�'c'c��;^b���<�?�=f�T��e2{�7�?���Z�nV'[W&V[Z��b�"���RP�J'x���a�b�A-ѷ������܄۠�-W� �ն��uj�ʷ��/a�)�Z%;"~c(a{���ZX�ĞZ(k��n]�Nm5�
۴%�����33Ҝ�W����m$)�"�E�{���Ɣ��T�%��^�g�K�.<MenLn��`��e�k(���������P��yC�F�4�d��[E*A��Ӏ�8�@��vh�4T�q %U���ra�"�!V�ɲ@�x�E���Mm�k<�����	����&�7[�w4:�<���Ì(�dދx��*�zv��Z��3�p�j�&Ӳ����$3E��t�)�gP4t9d8�f=�Z�q�Y������Y0Z��-�@�l�/j���S����-�1���� �+J��� �`R9���$kle�W���%�K&@��k_�֔|0uv%��X�j�,�I4�Vt=��n��m-fڅ�C���Xw/6ƆR *鴘��n&a9�830PpX�R�v�W��J6k\�d�7J��Ks6��k4�N<y���^�*B�S�y`�`Sc('t�Cla�Y��CJ��*��Q�@�
���+&;���բ��,������X����kh�k!�F\U�؜�+h��B�����&�;(���Jl*�͙E�tԭ�n��TFI���W��z�8�vFԸ,a�{[��lYL�Sh�X�K���^G[W���gtj$敂4�50�[�(ج��@���\�;�˖]�vl��-�m]�h�M	t����`�쑢,JF�4�Eܦ�MJ���:�2Q[AK-nV䲷X��b�5�em^Rw�vZOTN���4̐-	٣y���v�L�8�mc�kZ�xkJ�"�0�R���x�f��Ǻ0����5�����JU�骷�ٻ�X)(˳��ݘ��Y0����B��5Z�h��D�0�Z3r�e��^dd���0F���߄Gm"���.
�w+4�����2����O
�)N]�z�	(�kٙ@3��dauy/U%�R`
Y���M�@�kk����1�[z4 噒��^5��H�.�Q�f�t�@�����:j��N���,s�l[e��ݢjdvf�q漟,���F�V;�[���K��w,+q"���X�ì�:>{J9cI�%�3&�L������Ƒ�j����97 �)y��ͬɗR �UZʼ&LPx��M"�'��I0�AZwj�Ğ�$;Sw[(a�����mc�i*�rJJ,n�e%5:t!��.�`�蕇,�tXu �Gq��V��2eJ�yL1�ЀAJY]�/�F�ݭ$�=��B�w��H���B�H�̱��A�*R&nj�9V��ׂZS�h�";��L�*+�u�{L�Y������j�ՙ�h[nֻ�]�kb/sk�ܶ)n�Bo�cIX5��M��M6��hb���W3LF�Ն�[yu�-ɓ]�3j�b�P{S,�]���閮�:�Q�����r�և� f�'*���SF��n�Л1�ʽ�2�#Z����v�0��\�j��Z�3l�t-��nE���颮T�ײKڵ��\�1Њ��$䐴4Р�rhjY������ҡ������ԬY�`6�}��,��d2����@*Y�t�0�X���T��W�6\iD%���B�:6� V��jb���w2^�T��^Y��JWkh;��#�2XE��'�(#e!��-懰V��b]+;WC[XUnZ�2�T*�I��DG|�ٷ���;�bdJz��8��e��԰��]���A�ئ	��,�ٹb�mԲ+4iB[�QWH�WN�1�97F&�oe�!i]!��zrQPY��L��k-�*&i�Zvp-0S���nL��<�*�{!�/,�k(BK�"��T�Yiá;6�\�pȦ��6Ap<;Y���V6�1������%DkpG�XfY-��Ǔu�0�6�BAnv?;�͍.��3�c�c{��-]���.H"��TuJM	E��� �[���6j��',G���0���B���{�Bș��w7��#� `Sp	�5CXv�6�M��7Eԭ˷v���hA(c���kE^	�b��*�U�� X��ߥ�! ��/2%^2ꖋy �F]kaᥱ�Ӆ�MXi�C�]�[ͱ��J�ݍ���/�7���[Sde����l��mӆ򖳋v�br�W��i�r�ऩ�;�&���5\��a�
��J�h-WM�v�7���w�iJS�/j̙{�6��y�Ru��KH��3f,�3s(�6kF�-��,�6P[��7 6�sA-�y*6��/���~���tѠ�Y���+X��R,u�*\����6��������q�)J�;�"���sa��,_'�]�c����x�A�LJ�Nܸ��1�2�yM]�	\9z�ΪokbJ�q-����#SY����/oz�GR��\�׻�TL��Z��g$���`��� ��N ��N�2*�sw(\f@���W,cE���#.�"n�	��Ħ����;z�E��@�;ڑ�Q��AӋq@kiJ�� �0R�:�j��Z��:�m��+��^g4�vRX��w&a4��1VH���)���W�mT�Ay���2�A�X���k��b=
�*�S8���Jz�;7MRssu�jW%mfb��Y[Y �wJ��1RY%]J�U��NMw�^�4�,Ѡ�$B��%�.��36�G0���
��l��`�]h1o��ZٗM�I��J �qsS���\�J{���8��#��ʔ,pSC�D��� �V��ͻR��I�8�̘��Ď���(��]�(A��KR��NHå�Q��=�om"���*�Q��B�Em+�	�/bC(n��6�:�;D��u��B�1��$&^5�NB/�IOva��R��`0��Vd�n���.3��h���o^�3j酭!�S�x��)�yEe�6*��%w�՚m�j^'P�L�Ö�ǉ�B��ky$��&	��n���gv��j��6�a��Z���s��׆�ƴP��y�0���²��ֱ�^WF�jAo@Ÿ(3f��C)����1�-Y��oڀ'kC�EG�qޚ&��+�l ��̴���Z4^�J�݀]-�-n�ܢ�f(��F� Җ��q,e$&��Ǣ����6݋��E�j�cn�o6�tl`E���uɂ�$,��Usc���M'��n��[r�N���b��l.�yW{KQ)"X�j�4�v֢#�7k�si���Jm`��1.J���K���f�ٰ�4s.��C9���;�)��c+Z�pP�I�䙛tبK��$[
���[�8wNmFКvsk4���.Zxֹy�2+Rḭ[M�6դ@�w��[v���͙Y(��%��0����Sg� 
�~0brn�ͭN&hZ�*[�(إ�-/	���X�Y�IN�&�EU�xQ]�3d���!D�kaV�n���˥�&�+)<9EV�PӛDe��{j����m;J:��0�U+���"����0���9!���ݰ�H�9�-e�^h���(�X�e�M��.8UeM�h6�m&��I�����U���2=���������D�o�6ޭ۴mźۗBbj�@낆�wv�o-�F��'-&�:Fy�n�%�to+tʖ�ר
���CD���]=NT�8�&��7H
�Fr��i+���,u�1�C/r��ZA��R%��cӯT��!���`Ӥ�r�a���*]�Ȭ&����`cX%-.�����Iv��[j�WnS��ER@�:
�C�R]���a����E�����-�!g(��SqPu��I7�T�%�BL��i���Z�b�'.��t���Sblѵo��[�lX�
�[O0]�R��mۡG[\O]݇����Gup��v�����[J$�ͽB�;F��)FX���ne����!�@T5�^�%�Q����E�AS����^�,d
��y��g(*Ԁ݂�s�+�&�ɳ�)b�m3-�_
B�ږ.Yu����x%a�{R�-��	��B�]��z�/5�-n�C`�c`M�R%q����Ⱥ7ds\5;���T0������V�6�4%�.҇`�!��%eC��w���g�)����髻�`;CqX�-�An�����Ǣ����6�1B&S!,�N��Xig�&]�B�;6w-�5e֓�\`Y��Z�4�R�=�M�B�bIH;p��h8�XI7I[G%k�3��!X�	TX�\[V��K(�.!Y[�ܥN5�6���A��%�\[Vn����:(+���/4Ild[�"����l�f�mJ�f�3l�"ݩ��j��ٖ7e�m�(�{�5{X����VA4MOҊٴfm�[P,����C9�y�)& �Su���f��b�����gN9��J$��S��X�N�`G�)��$f5#�TmK����s+ZtVb���U���7�Z`t B��L�V��,, �	͓51A���-�x2�6dlzP��9���*�E -��E�29jU�s&�M�&�Cكm�Z�X�rBi���p)J��$�H�@��ŕo>�Z��A�zur��[N�Kv]՝T�Fn�7��E9���u��v��O���C�~j����Nn��ҘaX�KCjA��P�[.օ�=�e ��f�T�FYd��:�O.a�� �V���s�S�~,�zlB�@�ڙWe�fV��䐛7���$d֧E���;b�(��[���K
�qZ�^��E�fQ&�`ܭK+P�3RL:A�����yP(�a��M�;L?���b�E� j�+��E��]+0,ʶ))WF
��o �L�	�FX���Pci�Q@�����;6*i���Z�E�����WR�aV�c.�fW�jS1!1�=�1�n��Br���Q�-��r��T�a�5&1#�9{3T�>�Z�J���9�u��[5<+R�;��smȏl�k4IKZ3FU�u�qG��Y�"��,����#��˻�x��"��7I�@���L�[*�xo&�lL$x�`1������J�#L�Q55f�#��(%�b��d2�`�z4��NEN�K�Y����P�Kl�{)j����ʺ�.2��8�)Y-X�Zl`B������>��t$�S�E�GE��*����j@)���o
�Æ΄o2X��m�Y�'�boV̶L���Ͳ��k6 	�mރ2��bH�֛�CC�)�Kej9{����v�TXO)�{E۲V5g,e٧2����rL9+&ko;KN<,6H^�
G+e�%h�bfa.ˬ��n�'*yζ�\��R�C*Rc</@;���́2L sNԧf[DʵPԔ�*J�ݔ/sU��Sb��C��1�^�fF��A��snV"$��Z�wbr�8iɥ����F��.%.K��d)0�n��V��V���@��Tv޳�c�:q'Z�S3%d�Z0R�@�cXw���C���hnLKlީ�n�M5#6^d�yW�J��V��@Ų�'@lXv�&`�ZND�k,��o�V�!�njyl�Bn�"Umc<��tg!	���$Z1�b���*Pփ�rQk�W��f�WZV�+���
�D��$�im�e]�7��!����U�)�mi)�j�'�mfS$9�U�Q��nɢ�/)M�RD���;������� ���n=�V��Mؖ��k�NԺ�	;kMЂ޴#Ք��-WE:I�Enbyv����C�.c�����5���6��3�v�hV+�6��n76h�rF��,�Q��SƖ��3�i�X�*�Vk��V�����j��ʽ��%�%�ɱ��*[w/B�T�B�-:X�%��toK�����+�4�Uդ5�#����	b��̫�A"�6Z��x�pfZt��^��yw[��<���)�"�"BL,�[&J�-�J#�+:�Q���(X$��&ؚ�H��优����i�3hh�S%[Gv�� ����f��hX�^(X�Z@�q��s&P	"^��.*��voM�1X*��ɕ1�2�[JX��)�޹,JyQ'Z��ٮ�u�� �e�Fc�8��t:w�6�ۇn�ct���X�# nnIJ^0��L�ǖ;�iV7,ʔ/7�l��ly��&]6�`�Ս�-mX����KB�d�ݫ���n������z��h�#�`/E��Xw&j�K"�P� r�R�ذ��h���q<�>^��Oz�1㣦}/o�����D�h_\���4�̦]^�%����ѵ.R��^N��.�C�Ol��	%PI��`��s5��0�,��$�ʾ�����!��Y=`���Y��]qW�F�CBphp��1�m�Y�����6�Y 0�0�T5����{݌npDQ�ά}ȁ�)�Qu�m�4�/V�O�P��������+��uvCљ�+vʍ��-�ޓ{��`�膴,�%�e0P�Je������38�}*�T7ݰD a���;t����rP�E�o����i�FB0���8b&�D��.����ܱ7{�r��ѶK+X�e�2����n�m�h� ��� a�U͝c��_-՜	���rd ��W��97B���ud����E�pS���Zb�pdr� �;��4������w�fޱפ�L"���
�8�k.�6�����li���@���-&Ge��e���F�o�3d�Fƛ�ɜ4Qׄ�In��<'V��:�#C,nqE:]�mu��9Ч�}�H�\��<�h��.�[����5�8��P'o����H��� {�j�k;�cc
�qX F��e�*q�-�)�f>�`mXd�$d�(ӻd�ج�:M���"�(b�e�ydP�+:F����;fk�w1�8����Z�k$@�a�O���D-���J��ڹH=$��� �L���f����+�gp
d��-��9E�Ͱ��yu��p�>�Ԇt���9����]!,�95� jK�«��T��Y���V�.�ud9k�����4��g�' �w8[Ar� '��6��n�]v�Jv�ܗ���3��VN�%o���[�r�*�pkZOl��A�7���U�QC:��V@6:�o���:+N
_W�`]Ff**�k"NOT�D��\��y �EN�x3^����kH���T�_*�W!�+����γ3�e%:֌�q6kz�HV�Ӳ��,��tUv�O���8^bn�ג�n��*[S1�
@C,��/w��tYV} �7� 7;;{6�v#��+Df�]=�d8��E&����֗:��E-ViiYV'Kf�b{r��un,���ӂ����U6v����=��͝ף����u�]��+&�$.����WE�>�x��E��Q�7^܀w7�yE��"*+��:�x���WIgft|�9���+�#��8�T�>D���ܜ(��A�ueM�ܮn�mQ�=Oi'%�Q�#aʶz����j�SiŅh쏰���M#al�E�\��7:�uj�����4^ձ%k*[���ꕎ��`1�S#]�TN�B�xz��Y,U�y����rB�U[{:���%��u}��SQ�������}.�m��C�7C�2�#���J��"��4:���۩�ƜW5R�-��ڬ�y��2���9-k��ə��+1�`��J�3�V60��yl��٫u8��W]�uP.��ޫY���D�ӳ���:���u0��.��q��c��҈��f`|�k�}��O+E^��B�PF[K�s�2nr��LUǜ��-Y�}�y�Έ��t��'u��l�U�%jk�|�e��Q�����Mk��}C>_�E�{���wT��H\�qThT���XS���338�Q�ٲ������2,�π>c6ۥn轂��Q�孌����p����P2�Z��Y�&�|r}}/�Ck�s�jL�y-#�����mu2�����+���l�l���+�AS�ut-2����G�zi�H+W��z���<��t��x�V�1��Դd��i�ܿ	q�U겐`|���T9�\�c�Wu�6��_B�,��HͮӪ̔�e��������|�l�f|�������Y��۹�y9{���L�	����Q^.M*�^��e,�y.���!�4aئ�L֌Xt�r���B��}~�J,���n*��ˌ�p���gw��;�U�f��W]rܶgˁ��suj��C��+����/�"�ϛ��L�Q�^���b��ӹmrK���N���W���]�̤�=�!T&8��+�vqeĞ��k�W>�W�i��S�WЗ�2�h#����5��X&�$���u�巼��̤5���r���B�0�9I���f�$�B.�Tlڱ}8F�,f_i�WV�㐍T�̺�{Y��z�MkvR��z�h\r 3X/��o^bͫ�+

k��V���}R�U�	7�ĝ:� �U.=N��-�ˠ�wi��䚗Eݝ6�5�m*6�y�yh]��x�ށL]p��b���8���s�W^�-��N�[V����K�zޣ�����.K�v/���$�/���7�[:J�i5��gm�FU��V�=,M{̘C��k��~F�N�������w6�8�m��lf�k�Ǚ;�Ȭ��%���I���mN���Qɗ3:�[w��![�k4���R�*2v���N�ct,J��v�$1�ٰ�r�.���dԩl���5"�E*D�ˮ,�e�w%<�z+G�����[�x����Li_N&ޙ��\�����w#�nN�yC͇�ۨiZ ���N�uݣ�09#-:���;M4�n�ԏ9sӓ2�G��<���̆�]ޫ�tS;w�
~Y*506ݶ�JvR|�Y�ʛ�㽕/>��w5��:���ˌ�*7�t&��8����}S���Õͥ4u���-q�r&��"�A;�VBa�d,ޞ�:�R�<T/�m�k�KSء�t�j:��ܚ�A���}����n�P�J�eyxG�B�W^� �hrŇ��ۻyg�/a71�R��MnP�x���Т"�e.��c���Pjn�d�w!�it
�<�S;E�[*��e�L�<wY�)��IV
���|�L��5s�X�I`!NZ����+��6]���a��I�8Ϋ�`t�o+��q<o.��.�S�[��E�,�2)��Q��T�\�^_)U;OPz��M���m(r��������v2�OQ�������]�y��8�[�4*���o:��ݍl9)��|ծ�7�������<@�8�ܺ��Uz����Q��ֲr���]�YXSH�y̋����� �tZ�a%�u.��Q;f)::�Ό�u���pq�xz�6�������]�uh���9N����̻Q��Qiv�:�j��}Nֳa#x2��`}�������Fx�ӈ��@���̩}x@ڻp۹�5Y �1j[�wF�Uh��sdڗ[R�}v�u�fc�F�,s�`��p\�Y�s����w�� ���ձ�M��zeD�B'��N��y����ܮPTZ��ܷ.�Zu1��a�s�WW}�u�2���Λz�\�Sy:�ַϹ]�Gaܛ��S�V����՗�E��:�֊j���i	�7}�ҷo�әe��SVK�y EX�!4d���U�A&�K+��J��t]]�D�K���,�
��b�/v�����զ�V`P��$V�l��&��I��w.2�>@�; �K��Pq�6��/��f��1c�ȁ ��zR�e���J=��hr�zm<�G�o�!��4���e��L%*1I�ʀTlScǯ_n]��+� ������Ɲ"���S��!y����,�/���B�&��m��Sy�
���6)%ռPY���;��W��Gw+�T��`��8�/{:ڭ-�J�Ʒ1!`ٗR'¦)�e�]��X�ǻ���_7����X�	h�st�9�����.Noe)P 7q��Dj5D�i���@�7^����uN9�EmÓHUo��
��$)jyyo��Mt��)�g�ԏ�Û��v�֕���:�J)ug�����ʻIAR��9]vm���1�e�'����[;��,]��؝�ѭja��%v˳M��N���is���Y��U��ckUi6HE������0�o�z��"V���mٗRh��	�#�2c���U�)gM��C��.�����v������>�I����2��ej�Uw|��;�gq�v��L���Eʌ8���Q����)=��w$���It�G��.9�7Q��L���Vn�y�����q��wGK��-n,BK�3r�2�"���Vh�}�`�5���l�sHU���/���/04������\ح���o1����5�)U��9��r��T��M�@7�I�\��np�Z媞��wUγ����vo_+�=e���K��9]ل.�-�K* �!�C�v�]��F��]�C��掠���7�V��t������;D���.+�p�K,*k&���N�c�o	C2�qkD÷tt-��0�<�����aeh��ɫ�`��3�0��{���|hN޵�`�o3��qeة�8�m�M��#�N�d=��aW+�2���R�_f �,�Q.zV;}���o�х�:#Q;��P�8�o�즬�՘��ds��_4)�ÖTx�/���Ӈ]1�����s�͡A�����q�eNy�%�+E6(JJ�Sո\��-ea�X�C �Vʼ
�pPH�j�}�a*��6k��Ѝ�L���a����A�i�}�8=�s(�|*�.�d�֩�HS�,-1�j�*l�C�n�AOq�_�\h�#t�Ǩc�\���Kq�ko�[���V�X��&ؗ��JTj�e�j�WDUF-�ppՆY���
Te
�3_��K6���#��r�3d�¦n�o	���{�DQj�j�۔&��ܽh8^F��\*��ȷ��g�&u�h��ao/��\e� ��.�2FKp�)-}�n����J����N��-[�c�����#�s��1>��Y�V[�=*�߂� �����6.@k{��$�g^1ɦh:\Atj\q���XN�K-f��0%G-�A��Mm�o�=���czh��{�:渻�@�v���"�9e�Q3h��0tk�ۥJ ��n�[Zl��_֕�!�x��>�u�oMO1��U�h���yEna{z���:�W�I 7&�Kӽ�h���X�\����lN�sY.�F26�=d���JT�OY2�:8+FLd.�Y����u���z)��77H��it��e3]�)S�N)j�[a�Ƒ���経�΄Ꝓ��؂茜����)3�"��;k��YÁ[2�j��k;v����-hȊ��P�W�����G�ԹٗQ�����F�욻�1M}AO2&���f;O�uvOI�M����K��)�5��XGm]M.�oV쾙�L�.�>Fk�WRxwKK�%K��s������+��ݾ�)gQ������r�+���9��^�4��Q��\���t#x�ō9����J�
��0��r���7-�[�p�cn��o�/���4��%S�7NeY�!��WKPv�rsU��T}�]�Q�urގ���࠺��
��T�$W&Vou���71Y>����ke�Ɨ~�k�K�Ox-2ť�	�7T'�GQ�p��fڵ-�b�h��kb,Sz���~��8�2�[=��B ��Gs��� ���e��7�]å�;Z�&�B��C+!J�v`f������ŀy�i�w�u��r�R���4�l�9�r�&�T����5�hS��̔s�^&��Ŗ��kp�覵S���ﲙ���q�N�:��������\��u}��� ��ۣ�4b�E?P-2h���L�[ط���f��b�K�x�+�U�NˇUv^��a�M��ŊlCF"�M�b����8u(P,t�a���t�O�i燲 A�1W�Z�>����]xs`�0[_@&�ch�`�0ު�љF��XV�y=�o��C&�]�º�|�$����Co8�ҴG����b�Uj*P��Τ1�NtiAi-��p��R�@���g_vT1 %�꽗���h��L������
s���*����y �Mf��t�$�����[Z��;pIY:�� �퍙�D��,� �N�X��-����zJu��{@=�U0�� ��$��-���5�'���S�d��H;Ơ�	�o+�f�w��O 'oFGup���O[�SU,�r�9n��7ļ���
v����7�.���dΣ"a)G���#�����ɇ�����]gq
�rZG��}?Ga��nb��%�&���L8C�i�T�AZ��k��x���`۾d=TJ��]I1:�97ض����[��h`b�n�\�}�J�iJwX7���ۙO-@�7��8J[F��.���>�WF���Ұ[�X���z`�}�sz0�V3vrv�V�b�-����s���.��[��+���o[����=�B��Es��ڦX4Vz�Z�)ї�7Ba�Of��tN%�K%F�D��3פe��.褝FZM�:�I�`����W��ŵ��7��s��l�L�V������^�*�i��MV�M��v�V�ܞ�݌�;_3�:��N��3�ɺY�x6�� ��Z�\C��{��V����T�;��`=x�
j�ۅ�S��
�9gVچ��x�mp�Y�pv�j���	\[P�^�����ֳ�nu���b�r�1�Ճ�]��DX-s�;�Y��3���q4L�Z�5^
�'J7��%��g3[�5��;-�KV�=i���[lR���W�N�]��0P�G�l��U#�S��.亶�����ܴ�6pX�4Ro�٣G��78�GEK�ld���M�b򺹚�Ӷ����\yL�I�r��ò�c�.t�;��^��0�wd�!�}]����+����c���A���ܺ�f��;���.v�,�]ӝ|g\��9K�Y7�I�F�WP�ӧ0`��n��_�	]l�+�� %���O�"��͓��Zj�����Y�҃��3uu�ӖH�f�I[�]�ؚ��z/�ՠ�"gP���S��1�E>����M�'*tV9��5�5H�}���6�ݱƻ�U��#���o7:����˹Ԏ�wwwN����ݛ���goww\���FqI��1%: Q��Xj]��*	X�+�ɷ�>i�-�u��G/.�Y6	�IR�1���t�j�P*��ۤ2L�t)TAh�Q���H�J%^
�q�F�R�_EL�!�	�_Ej��,V���t�)Fth�r=�U�a: Yj��Ӣ@`H�I�,�iQZ��Ǖ�u��b����}~�x �6$tXE���T�Q����O&�
��t1�D��8�Z7�`�@���%V4�"�H��@"h�	�,�(��f��:���B{���p���u��j�tᚦ����89����Ц4��j�J�Q&���N��R
0� ƨ�E<��	�>��wDH�_r�%� a:Xk
{��T�s���T�%_
/�~f�1���?v`��P"�@� ���)�H��T
��O�̎����f���<������WV|X,"����V0�5�G
�T�#⊪*=Z��eTC,Ɲ:l)`G��lay�����\:��t��Ѧ�"�D*�%��5����U�wq�S6��]��qN�.��;9d�ح,�Đ��ɛV�鉷�ɋ��ոU����.��< �sT��-V�:�
��us�O%p��ZB������̺�aͰF���EDL�����=����zbw�<�ÛwS6�4r��5�Z�W��٦b���뭽��̕�;.��� {��x��G:\ x{+S$���#���]�]���W|+9Cu@�i��N!�f�ġ%����U��w�$N��!�[���l��p�zwU�E]�TT-��FV_Uᨸ�
ǐ�z������^��x{/�7���@�ҭwQ���r�Y��o[=�^Z̰��*�ki8�5;/�EL9�J�賂��6����X����kޘ7�7��|�P�C5z���o]=����f�uv뤶����͙�h�x�����Q��һ)B�\����niE.T��U�u��uw�4� � �ܕ��:�2;4�a��'ee5��P'�W[�Cu��Ƣ��.��]tn�ލl-�1��3K5!|O{-�����b�2K-n��JxkT��1�k�c�lIj��S؋�x��Fe]�\)i�}�Td��p�/�SΡ��L�.��z��3��_B����/��n��]7���}����������������������====7===,�ɒ�OOOOL�������������������������K��5���>��|]�R�+�o���[r �(bޣ�u]��ͮ>��p�&1t÷��J`�O^ح;׻���������ܬ�������- -�����P-O:l���8�s�d६����\)};Y��C%�k�N@F��ɥ�^־�c͛������R�l���,�벗Y{}ɚ��%�I�L=B�:b�0t�}�g�	�Y�yV"�GF���v�Y����kjɛx�D��o:_�^�n�����̜6fM7/�k37����h����w�ZV-x؝��b�����Y�DmK��#��]��-�x���R��Y,ab�3��$�Sn���m���S
CZU���ڝ���7�i�S��
.��6G1��w#��X.n���V�/�q��n�Co*[T�>vrmu^���u�$���*�)ؕpb�ڷ~~�҆�Ikt(P�-�۳2�1��j�j���XS%mf�-�ڸ���3�����mz,�F�`�Yt�)�j,���iZSlh�^�N�jNK6��<�;�GA��`9���B���d6E�ͽ�9Ey�=�e���cr�R.Dla5�]�[\����ju\��Q.f^)@�)������}��j��d����W�+���wwm�g�q�����Vt�ٛ#sΧS37!�l��mYÉF�t�
����rdɹٓ�����������������s����S����'����OOOOOOM�OOOMOOOOOOM�OOOMOOOOON��]�U��s��m��Y���dIK��<���1{&��ڴ=�M4�#1��J�l��E�1$�:31noT�+m�/���\Ƴe+�>�і��4����:t�Td��b`���:��T�c�V�.s&���s��Kwڻ�����ĕA}O� e-��]ݳdm6TmX�y]�m��M��7�<�#�N�v������u�*��J�衅�M�sw%Is�٫��N�u��yD�4u�L�dmZ�8JG�W)S%�n��Ro���Zg]pVl6��t��A�Wl(i�f� �9����j�¥��{�؄"̥H1�}2�n��^��+fp�@M�l76P���\1�sX�'.CA�LlW����W{�xÒ��&�=j�\�����+`�\����[ֳ+�t�Q�4��j���W[S�"��U�Uކ�H�x����V��8��G,a�u�$�D�7W��*�D�4�w��k"^U��_5��pr_N��+4_G�+R�\�����|�A��y���c�gguj����(Tmh+����s�o*�슳u7��%qI�T�i�V(1��g`���,�d����x
t^����{}<=��w���OOO���������������====2d��Գ������ӓ���'�������'�{����w��읖��<��U��k�݌[ڪ���g�X�Bi�����f�V �X��*����s0C�yEu�{l�gn�����$)	��:@�1p,�0�1��f���sO��YѤ�1��NR�Ԩv��!��n�� S�#�Mi3��_3��pՉ�._J�`u�T��%<S;Y;q�����r�������spK������lD����F-�\E�W*U�q�u������Y��F�^�.Z,�.�����bEf�*Mu�\�v���[	U�ge���X�ُ0�H�����4��	0��Y���2s3'��w�c|&*�-���joe��s.�˯����k2��nC�ARWk���n�9bv:�'y姝ē[:�I�s7��J���+�n��/(�n��NQ�8���⬭�-�T���K=�G0oN�R�ʝe�`h灉�3�q���=�^��+�0d���[>��0_r�����n;��cXy�xPn�p���k* ��3�p�&�s.��3�[\%X� ��k[ĥPм�۪�K�uos�:���1A}���S�LInL�Z�:�b�g����ݔ]b�Ǟ�I��/�����]e�b�y�\�v6_mb��ޏ��ۡ����p�ON�OOOOON�Fzzzzzzzrzzzd����ɓ'��========>���zzzzzzzz}==,�������XB���������$x4�
����7'e�k�n����=����������`+�`_�r�Ռ�!��c�uֹ�u4�n�"�9nc�6fr��ʴ��PȔ�i>0J�S���8{٨��/;9�ĎqG�Wm�F���b?5նv�C�8Ґ����Y����T3w9K#{��@���j�G�3z/jj�q8���#���)uӯQa��S���{%M:�w�w�._Z����t�Oxu�ءA�-V��;:%r���r-���'Ţ��G�[B�,�TY]�p��m/�V��|�R*���V�
�����G�FQ���I�Wy���+R�;���k���M&�fF���>}�&����(֠�3��17L����IG�aَ�PȻUҌoI�R��u.тJu�;�ޘR��K����7��]@���Q������@ع�V�x�;�9��<�h����1>l�ok;���^��4�V�U�}{]��X���_Hk���^����u�c9i�����x	S}��js�-��\[箝cQ�Ͳ<	:1��w���v)�㷪��D=
J�G��&Q�y�{M�Q=����=��4 @��֡�mʅu�υi���:����ڛ�<|V�'�r��������������w����O�����������g����L�2x�����������������������===;㥊��nawqa��hN�]��JZ%A�t�R�,�j&�)t3�V0�PO5���\�u��v�7�Z�װv�,�Y�����ؔv�u	��|�`����L�tu�ι!U�1ye�/}�]u������5ubD�7\�����ƫ�F��m�Zu힘w:�WlW.>"�{���J-$b�T��k7�ȴu�2��r�
��Cd�-!S�k�)����PS���,�L�·�#o2mV�����ghP��ǝg
��d$:��]��D�u�;�*�����4*���ʮB��8Q��=�v�_6�����(�[v���g��]&�aTLi��7��g���%a���IhݷuԒ湼�݋��4�C�q���5VY1�\�
�a.ñI�ṣf�7�k���.+4�ͅ
˨�1�D[[g'>U(���L�j�9u��-+����������p�q���gP��e�Sƥ1q�����u�����)&��fr�6�c5ǖ�*�Dn�"��]F�9C�{:�GE��}/u���\(v�hӃ�2�1.��s��s��]�ioo0�S�LWP�O�czu�����h�Y��\(�(�����ss1F���ReЖ1�E6��/��� 8�V�pbJb�b��Ҳ��/e.xwf�8��n�ie������D���p�'sorZ�u|+5�Gd���h��Av�՝z,��l�;������м|}��]�f[�nݻv�-��۷nݻv�ۓ����&L�<OOOOOOOOOOO��ӽ��w����W����ze�9�
�g�lV� ����ѻb��2p�z�:�{�m�mogc�����U��D0ܰ
o�Z�d*^�33.]K���iQ�k+Hk*S�.໱0�����w�Q�,Ƭ�Q��9���w:WVYydt�&����)�ز ,�[I[ˡGu���9�v�!s2ڛ���Z�tmy��/e_��1���U�3��ï.��9��X��v��4w�'GOh\o.�Ãr���!wֵH��@gA�]O���l��W���ٯ�Y҉��)<鱔/�l��m{\�H�'Z�΋�۩�&��I�w�<1�V���P�]�m�&{��[��N��\��t�Exzi�}��:��iq���B��d�p�z�m�V��k�nr�3�3i&0u����䓛�Xණ�����Q��ڿ�}O����{qhq8�5������+V,���t��R��o�MQ!���"#�V�׮�=����L^�}�ŉ���M9���F�p~�D��Y�pbX�)#�>���;�8O!�K0�KVmS⍗x�5`A�YZd�Dۏk�I�n#|�8��wv�{Χ���^u���N�Zʃr�v�Zgz���J��i���bVV�ۘ������3p텔�E��5����vY��D'6�X�'�H�Em{Ԍ�o������|Ov뮁�g�޺#�q���9>����zzzzzzz}==����������zzzzdɓ'��========;==���������w�����y��Di�}@ȹ:��͕�G,�_�����]��&X=��!n
0X�)R�S���v�z��|�^Q%nb�vQS���o ĲnIk���������P��:��٩�s���8�����=��`��1:f+z��-��9J�"���,��K$˛�fO{����[�S�ָYO+��`���s7�u' �]�EIW��>���Y��p�V �M�y�pVz����5�L9ynˮY���A^1*_���/s,2��HZ�9:��;�s{n��.(��{V٨��!^]5�o#�L�w��:ë�tG7E��V�5m�x^v��J���"gUޚQ)�E1���oT��5j���3�u���9��7F����򺯀����s+Wd�.�<�m�-�/���fDP�r���GOt����ʺƱ�0���#�u+b�5Z6`�J��Z3���Y��}�F��:.�T^�,H�艎����':-K�tp�%s:��/�Y�UR|a#*�B�}(Mڷ��{�ǈZ�%��"�-��a�ؕX�Klq��b��ݵG��jI�N�R�b��@z�i�vw�S���^��/��|%d�-x*�r�D�ҷ�P���-�;O�TX�(�u4V�h�c�20���q���Iw�8�Ĳ
ڪW��8UR��M�	�<Fn<�кYf�ղ-����E4k���]zv��t��>�ׅL��n�ytt�=-۹�~�97>������������������zzzzzzz}==��驓&OOOK=======>����zzzzzzz}===,���ۭ���M�lz��VL�zB_Ww5:�� ��38�7K����_k�|��{��}�sv�0���2ŋ�b��t2�Vӓw^�ݵA���5U�x��G'v{x�,��C�0$�:=�E���V�6:C�;�̗C����/�D^Bզ�-]^↕}�u5�������ju�*�5�ۇ��1֡��S�u�����G�s�CB��}Ogb�{�Rp���'��T��y��Y|ܽ8�u�]�j���|��J��p�=�/y\<C,[6y�>3��8�b��f�3���v�Ρ9�,!�Vk��i�����u�:ζkxq�V�"p���x˨�uϟ2���|�:)�<�q���G9�I�V�oB[GT��M���y�7�6�gt�YK��ƌԖ��L���A��S��c�hjT9�AH#��!�J��/������5��Wa��@Sα0��;̅2-h�}�A�2��f���86��r��t�m����1_�HV}�IǔY�3�FR}��1�v�BL5�fP�zA���Y�ׯiQhL�c-�Cj<0�%ˎ^Lܽ����TC�dWJ#���E6�(���zy��v;���\|���7�KeNb<��l�/Ir<�n㵯����T�g:�/�Z;�wJ+�<*���=��8�Oy��X^�"Y��4�˟}S9D�`Q �թ;�:O��nλy*
�N8������������d �� hAr���G}Uח�nT�|��وJ��0��m�r΁�|�fM�����䯟>���<Ni�2ej�C��Z�6>r�s�k:���I�%�VuO���U��j��ХL����ӧ�OW�D{ ˡ�i�v��)o<�G[�apRKn�y��]�:���=�j����t��.�����X󾛡��4�Jɓ��N](��&�e白���X�����|U�K,4sDS�y��9��o����,es�f77y �t�}A
�1v�b��9гԎ�L����ق��N��Y�5��k�^�kb�R�4l�۞KvW\]�ub�쾸z�X����̣E;�b��WR�m�������Q��V$��ph�fV.5C��{��>�-*��S{�e�T�Rq:4�)5�C-R����\�!�^F:��F^��gm@��{L]�Ƭ��S|^���Y�d�"�T�� ʧO��VX�v������X)0�!�2���)p�O�f�bgE��˺���l����-�*Ve�B75q�p�jJ������>[�y�.�3{z��
_2�W��Ơm݁0�*`U��3���lS�t����\����ب�+iPClf]9M1�Ԥ��1��6��u�t����D U�D��{ҖT	gvg��#���«d���>�і�����h������R�)I04	4Et�R�O�>��u�	:�=��]ۻ�o��K���W\�m�,m��9*el�u��f�A�]+.Y+�vg-&��Ei�T��l�2�(j�PU{/�J4sX��T8u�.��*�gS\�����kew[�S8⸄�m�4�#�����&��-B,�n�n�s�]������0-z�����¤`���,�Rٻ�^�����Ggc�/���oR�MX�٤v��K]ݒ3Qǝ�%����A�KV�0��x�4���Ȝ��x`���9�	���+uPm�a�U#v��o����n�|�blm�]�ڜ��ہa�;��A�*��hSۭ]-�D\Xp�)v�c�[�nE�a6MX3�MAc���vԬ��o��z9d�Ux�yY[H��Ҡ(]�ޝ3`�o.��-O�xa@#�x�+�oI� ���}X,շ�t��]��D�͍�.��-1kf�]�2;�x7�G�7�N�d��ۆ���/s4�)W�G�����* a���C��]eVʵە��0wN��X4_����mv�[��F��>��9e�%'}tUh�½"Ժ�$��&���yyGm>�l�l�ı�ڀ�h6��M�uˌ㵣.��f$�t�4�w���+(JMF	� 0�E�5�Ԅ6�L��6ɣF�LSi*i0����ai��\��E�K�Al�x�e�˦Z,RUA"�:4=4��ek�t��J��#��CX]��K��H9B��H"�jx���v�̙9=98��w���`�31���b�)'�w�Ϯ]\v�T(��b�������NNC�ڦ�~J�Z�J�UQ\��s����X��3TĬ
:�ʒ��̰���95;98Z�* Z�UV���]5)Y��U�mj��X*�k2����[=�`Y����N嵇R���݈��&�k���kZ�b�(�oZ�pw�m9l���ٛ�ꙁ�*c:�Y]��������a>aG��¼�auA�4�s��)[*�3(یm�i�ǎ&��F��]�i�M8�;99;>�C�`W��1��.�;w�8�D�5�e�Ӌ�Ki�A6�4f2�j�;�I�z�TՋ!UF%�HsF��r�F�[��ӋZ3����9�q��q) �eӹ������?S�-+mq �nf�pM&�G'�\
��ϸkn�ƥ��Ɛ~5���$m1R�_Ʈ[R�T�K��E�8ջrT��J�̳}��z�=2},�������dL\�7*KaC*�!�c4��b"�ʮ@bot֫�E�[,�h��3w}�>���뢀9ʄ���U�KF�֪nF���ke6ْ'�G����ri+Jߝ
&������9W�.�<���nӎ�Q�?�:�`Q�z��?�7F�
�3�aP���4��c5��`�S��� ֐y^��iWS�;�hUѠ
�TS���}T�X�z���h�h3�R�^hY�U�n�n��ݶfZ����ؙ�kݞ��qyZfhy���ᦊ�xm5ޞ���g����j�����j�j��y���(���Uk�^��<N��z��p��S��z]���>��m�L1�|�;��{�]�7��o��(�Ϡ�3���^����7���,���ޫ�V{����A�~�,>(�=溑][�J�W����cջ�l�W)��Ww�{}"��\��8����Fw��J���̧��"��W������~�a�������^o���=��>ѝ�y��/u�Vx��g��>�#G�Y�(ɕS��۽��sn�Ї쾌���w���w�Ө�5�sO=՛wb��_d��»�^�><��ה�k�gg�w��e{v�k���j�ެ�'^�Xz�˯w,��
n���U������,��W����oRG����}�I�T��w|4�v���־ͷtE^�D<C�Ao�!�	�{���'�����6���V�K[z�3YP�R�.|�I!�Oy��f��ä�&į�jN\s;�`��;���JW�Y�J��N��P��ݛ�"߇p��d� 5���#;O�a����,�.���
~�h�K�3�n����ht�{��="�F��r}��p���8k�aղ'�8�>��~��Ѱz�{u�?A�npd��ܟP׍ �1��;Zyu���fY#�N����Gλ؛}V3v�L����ֆ�u���X*���D�}���ᾝn<�ߪ&���]��
���#��z,��/���;���^��z��f���3~�����X��a��5��㽸�8p�zM��հ�����p
�8�ٞ�g��U���Z=� VV����p�v����.�u8����NZ�ӷ���?06�/�h�}�|�������_5o{�N���7�.��j����G�V?����Oýn�T)t/{�=�WuOB5t�Ǽ�{��ʽ;�y���A�k喳�d��L���YA�F?]n����=R�.횕Б�B�յ2k-�wn;��:��������Mv�����X���Yw'ne��M-˘dݜ���8 �+b�4r�L�J-�er����r�wk2�J���jop��t���ȷ�2�UeT	ݼ��@w�I�Uʝ��g�J���w^���u�W� ���r��C�ܗ��F���8�^��^߸uHG��KϚ��r7{zG6vHm��n�i�EX�����ӸoEWn�\�f�.4^����vn������E�6#���Qs��������Ez���W��Ny�ݙ-�c�������+ۯ��h�U���'���n�X�Ͳ�����a��E��l{+\Y1A�z�%��95m�n����ޛ������8R��[�J������k��Z�U^��#s��r{)w�.���}{õ��7�)�׿A��e���9۠n�q�A�=�O���x�w{U-�S�[ �q}���3�^��=¯׸��j|�{�چc��<b�*�j�S>�u�@h!��3M�sK6���������r=��Z��_;μ�t"�&���o�&`K6�w�'r=|��|�q
�� LV͞�
Ы�Q�t��>O��o�now �׃�q�Q([��\t�R*�m�}�]ou٬����x�=�ǌ~�|��^�"���c�����yD�u9�٘țKP�/�:����UZ�;�]Ki�
�tu�[ݧ{&���W���x�����K���O[r����3���r�^�^�s�ew�}dz��n�n�2��{}Ǽ���[�j���V�_��+����$egg�v�������]��%��H����=�x���C^�j*�{��esȌ�g�3�I^�N�|�����v�&�����{���VבO�}k��}5Oa�]ces$�d'�GW����Ǩ}K�T��7�9�;Gfz�s��y���^c��Z�A�#Y��d����x�O^(��L��՛�z��_|$0�+��y�.=�b�C���;:�K&Z�y^ G�gz�z�����~�<��w��;r����ت�C���g��oY���'7�o{|(��>U~���3����h��}�e����s�V���4��UR���=��ҽVS��O���$�?_����z^�r}�g_�v���*�f��r�m)%��{9��׽Q.��Z����,~=�1��ݷ���\ʻ�>_e�>��_V)Q���u�y��9AKZ5!`�Q(�v�����*eMy�/�qL��1XS?*��xg�P��r���h,�Z���ӕ�ث�	M^q'$$���KwٯW������3x���=�s�&7[�׆��|~�����r�uZ��s��u���יǠ�0_;� =����r�g����z�,d{��޿S�Y��7�_�����L�w��)ޒ��.�]GN��rw���}7ݓ�3D���|{ۦ��-�~��`]�~~v|1D�u���p"��l��.�z� v��D�Dg���g�s�w� ���RC��X�n��{	^���?v�ib�f���.mN�wa׍��5��o�u]��|6�徣�iڣ�}״����9]
��5^i�r������!�j\5. jC�M�o�xﺑ��$�/�{�]�ၽ'k�������0���;���\:����G�h���g=��ZN�nꀪ���C�er�U�;�v�N��_VqX3���UX����VuI���Hu�N��V�
C�2������Eݕ�on��zz��f c��86d��'C�*u��7�e:�_80�[H>��~ ��VnMZue�J5�r�9bu�� �:���j��-+Q�廉2�E�;]i�}��XK��ʾ1�����v�.�(��>�����je?.�������}*����yA��sf����g�z@]�XǗ�w^��V*sVx�����7��w�;����-m�x�y���N�|� 9c�������q�g�ݻQ{�~�ǯ�*Og���/T���+#+�Ժu�����@�������2n���}����n��/ú�ɿ^���+��l�|�|��\�˞�^~wF�5����2�bu�磺�j\}���ok�7`�3ׯ�;xzC��Zn�����J�T�����w��uԗ�/J����ޕ��N���I�_��΍]}�Vn��r�1����ֳ�OکrV[��\�:�?K�.���ٖ��Z^K�駳�o�E�γ�heg{�kK�4�.��z�{��4Y�w;"���.ȇG=O;�����]�8('�U�zN_|�j��ڝ�w9�@�ѝ�%�S�TQlMX����H�Roya����˼`e4Q���f��0,��I�t���H���:�1�qc�i��ttE����M0�wV��ƞ��ŵ'.N�nĠ�f���pt ���ݹ�L�}A�V.K]n�v��W����O��+oI��y���^���O��en.ʴ��0��y�ʦ&xx�=;F�w���񜵟y2�@f�2ɮ)P�w�z�&S��o���=D���go�s=���{��V�Y�{9��[,_F�i�:q{�Wm��ǞS�M�����ޚ��}�qW=]���ǿy�-S��ēw'�ꇢ��.�i�/}� �����۰:�?��o�ֳ]��w��ް<��^U���Tʢ=�J7�K�M�`4������[Q����cV�g�K}^�~?eAm�������'��G���Qɞ������6_p�h�������`Iy�XI��}~ߞ�r�ѓ%f�/��}�|`�V�����}ɏi�߁�������y��YVis�;/��v�~ꬩ�]\5���n�2����ٱ=���ך�
��������z��Mw��9���ڹ�ҡ��m�G�"�}�$"�X'g]F����NN2v�0�G
��/�����3��e4�jw���7�Յ�7e։r�%��υ�N��:��p�Gv�积In��k��`�X�56���7ӵ�ۊvtk����ݿ*�֮�� �u�s��3��ڡ���hNt��5F��&{�z����[�!��>��*\��d�1�gŲ絯{M��> ������נul� [4
T��}���7�6�����:�d�%PQ6)��0e�ܷ��G��˕+O^�G��f��/>�G�K��`ǆ��\vk��kݢ}��};[D�\�)��B���:��݋~~7uY�62m�_��U{צ��!��~X�6l?`�^�m�d"��*�x
����xi��F{�Y�[��L�Eia���|���Ϥ��U1����ܣ���A�'�
��4Y��L���9�jn��KhUe3�~��w'����xo��:�.�[�5�6�{�}�������p<i�֜�����'���U�������]G����U��z�-:���&;i�F���0ĝ��mg�5>��}5Z���&��eQ��yS��y��֘ECR-ߐц� �E��������Y���9��־���\W7���W��TW�tU.�H����)�5�p��zN�S�s� �m�؝W�v+�9�&J)gios�-ɀ�j��2�%(�Z�t(< �"ʦ
ڕ	�x���}Y�kzA����^����^�Sk�����~7n�W�j��\;�O�+�Ϗ5�>}����z����ʲ��h���v}9�]�e�?W�������b�y���zz��]V�w�A���^zq����۽�W�}:��fN���>���$�7��},���U����G�ܜ��-�{����c�\��0ʘ��l?[��9��o�O���7c�w�����5Sʿ)O�B��pr��}7�T���Rn̗+��m5'?�ަ��oh�{�t�~}�Af��[6���]���^m�,L$�Ogo"zx�_X��t�ނ{`�{�C=��кB���%]F��U���ߧ`j��W��iK��W
Ի����^l�b��_���\v��,�7v{cH���7F��"rs���pH��ޝ^�bN����w�݅��7e; \�̻�o:��,AP-�J��#W�W��c�u���
�������gc�����4n��=���Va�#w�"�)˛<s���xL8e9ט5Q�G����g��q#GPmM�A�T	wr⪕���ޜ.����j�~�����_K}��Ʀ/�ϫ��{}㏘ZqF��z�xdݏN���jL����	�������h^�)��%ßnm;]�I���x�u����/S�^�C���+�c����ס���n!˾χ�fo|�6{������5N�R�V��v�1�-o��M^�WmF牒����|�o���I����7�Ϝ��s��+�l/J��sޭ�|C��Y�{�٦w k�ݵ�'��1F���Z�� "�7~��+t!���:C��H�|����X�/ڸ��~�~�6y���=9@D�;Z�*�^��
��N׬`���l�Ft�Ɂ��;��n�<S~��ګe{a���n8�՗���\�˞[�j�=Qw�Z������ԇ�ޞf|z[������\5��5�V��� *.R��St���X�VR��J���L�h�bu8@5��J�.�=����urp`ݧ��چa�wX�5Z��ɕ6���:���Ϸj!��!'�vI�]w�mj�#r^õ�Qx�ׇ"���b�nJ�B�qK0�6�v6`�CU�w���MY�_I��������v;�V9����^�.��]�F�~=�Ws��Z�%n���6�� ��֭E8RZ6�U�0�k��I��/pjN;���O���o,���#D˸E����﯒>]����{H��1Yɸއe��课U�W�˘u'Rr�m��Y���<m�t�B_]@�V�ú"��P/7�]W�-���A���}�W�:��o����A�M�e�K�)��ۛU�pX Y�i�=ȑ��r�:��Ab$�"�*uK��:Kuv�70�A��w����L�O���q	��x��;��ik#W����m�K�ݩN]j�1l�ѳ���(Z��ރjV=�
�Q����"���N�]'r׹���H<�Ն�����;a��5�f���*���t��R@�����p�j��TpnL8^�v�*pCU�bN�z��<y���%��)1,[nf#�]�6L��a�on����j	mYUv��4�;|�nu��S��K��{�|hv,ʉ}YqQ!i˕v�m��3�W.�٫r��l`q�a>3�D�}�"-��-S�)=���kc���v	�����a��<c�'|�DmR���=Q�Y�N�k��w_p0E��R ��I������n�Vf�._yL��s�F��ŷ�������90=�\���@>�rX�CDQ{q���Umq&�7�pVCԬ`4/k���9��}��=oY��sF�q�]j��m<���㜃�x�v�1�DҷKuWGll��=�n��%̮�:��SB�4��\��]��u�7���2�������5��]�3K9��\J�8�b'-u�ٛ|���kM���3��u+AP=MM��o ���fQ��
�q/Frی�ru�\�\��83[�f��S�gm1�b=��u4=�9�͙�o�O)��lvxhK�ԡ�)���@�},�����n�R�u��\�;�t�[��b6{�����V�3�P��,ڼ6`
����'9D�k��fR�b"�W؞��8�T剾�+��͠�v�^t�DI�X�t+�μ���kcn��ׄ*�'n�V��}D]��S��;�8�r����E��z֝˝]�E�G�6#Z��&\�[�kuU�^>�tu]���0nb��s��n��ki��i6�_�[ϊ7+�(r�6�4L�ؓ�	�J��9�{f�u���n�,������G��fތQT��!R9�Nu��̖4Cc7y\��B�0��a��R�6JT�T3I��3:���WAchT��n%�f���ɓSӓ�����9s�i̺�&e�W�JZ[Z#l`[u�;�̷3myk�'i�;~0+�9��K�1YC'�s�s�7k�W�R����J�ӆ*�E+eNe��T+�2!�ְԬ���ݙ��Mϧ'-��<,~��\�LJ�P?�i�m���~8,�^ڋZ�:ʴ��p�`�E�\��s#2z~NNMr�PkJ��J�i-9�3�]R��uB啩iekuL�DKb�B������}999m�-����e�t\�k0�V#�Ċ��I�i#��%)�\J�q�aFV�{���Y�����Ȱ�k+o��,�Cr´��a�l[ǚ���V6��Z�Typ@ϩbbn���-Qt̖r};996���S_kX��kmsz�1-e�J#�f��9L�Z�%���k�L�
��֪�\M���NC�y^j�2�eֱfZ�.9��M�b�mˬ�����n��6�PT�Q���_�b+��2�ݽ�u�]32�2�)�]Z�o�SxPX"|�˥MN��z�߻��T>#�y�"��*piu>γٷ���C[cWP��͛��:�껧�[|rV�_�)�'��{��R�ۭov�7{��鞦ۓ~��p�m��q����d{[`Y	֥>|��$���3�~���o9c�X�m�Q7�\b1
33x���/|V� 9|������&ϖf� ��끚Xq�w��E���R�w/�V�]�nՊ]����a{��;6��c�P��f|CT�,f/p�Uڪ!V^��y�����;���l"tZ���=��c0���|�/� s 3g�Mo�&<���<7�hTQ���<zo��~�,�,�5�R����+�pm�B}�U�=��VUw���<�i'�&�1��/��DD�S��R�Gnދ%�����e7ɨ�t���͏� q�O�D���x�{[��6�>\�͇#�T��-�v��n&$�`�,��/�#��
����������yM��j$�}�1x�Kbݰ�x�T���\�8dΟTna;��-Gn8r�<�|����|���!�'�K9=&J�g±\Is���%k=T����_^������H��@�;{�M��M�Ɩ0+>�#H����� 	�%�����G�spȪ`��*"ҹ��n�=j`oޏ�C�>����G����>�b��(�뱿e� ?s�d���'n�}՚j�e��m�Ưq~1���$��Ђ�����ٙ@^{�$����2�+jwv��]M�O[$U�]z�mdl���6�y����to�(���4�+��I:j�]�pO��a�B����br��Sl�WI'S���=�]�
�c�̩�:䂇��=��,Z�|^ܗ����7�GO�38>��@3ys�k��nT��` U�tx7�X�l�׈QՔ������v(t�|��{-����]���
�F�0
)|�S_.�Uz~����!����{S��1d��In����Z�����5�U���t������6��H��Ԗ�^Dq�.�继d}_]4�>�0������@|P3j��k�aۯ�"��p۞��1����#���Nb����o��T�}ȝ��N��+e6���@�mm����)��m/�y���q���s��]������43nϓ�^���_��֟ho��n]���q|�n|q����:{[]�Ö-�|#~c ��w޹��P�{.�G43^�g��h��;��E<=Mbo��y*���\��:_tGd�q`�q'�k�b��	I�.ZEg���b�Hj�1qɥ��mĐ�IB�+)cq�לn
@'��CW��@�s�=~��B�g F�m��c������s.�eL���Z�eĩp2�s����S @�i��6P�r'+T��+v�x�쳌����;*�q-���Dܰ�	l�So��7.���W�D�����U���λ�V�b*��hO�Hj��)Q��AVܴj+8Ն���ڝ�E�sǜ��<O�Q��Q����1�%��QC���xX�<�1�Q�x>�.,3�n�����hv�0�����+ה�l�>-���-�dUc�4_Liouv<��hL����)���M�*�N����;;K�\�'!{7a�<����>��,R,,Sq'��g���i���5�J��s�O]ME�Or3S�Z�� ��GS�]>53a���=v��'o[ �[~�|MkdZ~ơ��S1�.��o<\\�Niye��w�<���7�z@��/�F��杇�si���xdV��Cp;�"�M�`*UV��8R8�?��)DG��8���t@[��4��(V�<��kǗf��>Q���6������ 5��+2�O_GC	�])�(r�⏕���3Ka��[�'�����y�z:�Vئ;B��i�!�e��vy��O�#:C�j�v����t�J}���a<|%a�� ee�͛�VDĺ����Ɔa`�69 ����<퉺e��{~�7�n�T2Ҏzy�'��S�o%�K�΍�jgm�G�Q������D=�����T�t| ���
<�쁺��%`a�x��Q�(C�:�C�l�ơ�1�`Nsc�ǔC0#�D�Ⱦi��"=A����N贓�jz�̆�|�������}����6��f���xo\�F����*]68�ͩVsEu�~z�F�%0��﫨���W=�4�`c������G�j�h��ْm�]�M]G3S����-m�ә8t/���<�����s��y�N��o1��$�Qi���)N��w��s�<P[	b�ywe��2��T�ZU̱�0U?���ߓa���Oq�
9Ec�(�i��T��ͻ糛M���Db���K�cYo��Kҷ�EU8bSq�n���`E���ٷo�������vᵄ&�r��g1�-~��G0Z�K9c��6)�F�GF$Y��zG��R&�c_F:i;1���\Ӌ�B������
#�g�:��f5 C%d;xl�HN9@����!�l(�=���<s/���y���WSo5/nt���ן��9�~B��?��� m^�w0!8�^�@�'��,r�f@xer��b1�ڂ��G���J>�ֶ(䫩�94�8���:w�3z�9���;�V�M��w�Z�����}�p
�p1Gs`���)���{�O3{�B:)���
1���wS���M' e��y�^9��O��|��E�ʆ�Ѽ���5�O�d%
�K�R��+7�sp��fpf�)��m��w@6��k�`6�ʺQ��osM��ܧ�c7s~����μ���
�ίnd陋�I:d�E�|�*�^j��{���y��eN]�
�6-��H�9�s+q�nE�7H����V�;�����,(8��³�b�؂o�Op��i���^ʱJ����������^�|E��Y݁S����G�[3�8��ç�ϤC���@LA�=j8Ѡ�B���[c�t���̰�k�g�M�c����t�=�-`�Ϳ�9��w5�����A}d\�ӡ�M������5j4c�c&��|�b�MЌ](�0�z,�� 1�� ���D8��5����:��oh����XT\�Ɍ�AA>�p�8��ө�9���D�@ב����rͦ��I��ܜpS��gF��dU<]5.�b�դu�?��`'�.��~�p����V����G.�byL�0d"�"�N�vryĭ˭U=9���8�@s��EȾO�����׃��+�6����Oq��+�6T�6CpB�5�����}�O����39��-I��$�s���z���*j��m΁�B�8�X1n�����5�S��h�/�;�N�:��,Z�7�O���2��o��<����f�*�|���:��>�:����DZzw}0|ƹ��5�(!d�$υ�96�՛�&�d�Y�E\����5��,5�����HI\��fW~����~4%�j�0:ķ]%ڈ�[�$��͠(�Ǩ�ū׈(�����ɝ9�݄��5�w���jQ���؀X=���,pp�!Ӄ}.%��Ec�̻�7�ڙ��nl3_'�65,]ӎ>�L��i1���y'C�@�g�k~�q�y�����k�,��?y�.|6�����Fs_�lg�m֏�aщ�k��sVE��~�Qg!�5�YTn�)��,�4�˹ݚ�#�bz4gϊ�}d(H�l�k	m������{����J~zn��Z7ߧ��&�n�A8��fem8X�xf��X����Y�Ŀ���R�i.+#K�i��㷜
�)��:��*ڦ���q��Mݕ�OL��h��K�Yְ�$:��U��ߣ��C� ��E�仵�c����]��{(�h*h<���>o'��g��`$��:������l:�!�n"bK�ܚZ"P���(`&����&�r���t:��n}�l�r�d�a>�u��'T��)NS��u�j>�&un"�ݓ�e����O�>i��p�I`��
^ aؖ ]����R9�y�h��,�]��&�V'��)�� d�lra��qik��Ӈy��e�vl��2�,���A�����0c����3��[zϻ3�֯=��g�`'y��dn�&gh�{���4���i~��8���mR�3�Y�?�ƭj��yM�6@�q��{8��:��d9����&`�J��i�hƀ���^��F������I���6���s����[�*�q1��P���ά3T�w�iN{הn%\���$��ٸX�5쭁��ۉ1ݳfu�;9�89��[�ɝ�}Sl+�]�*��@t�����u�("��E/1�B� ַZ5s[��%e
GS�����{���J�Us7��v_��w�鴹���1���<Q�����k���޻a���a�vb�>5�~t1�K�ia^�7�oa�w����U.Zئe3�j$�t5h��������ys��*���/|��
N�7��V�v�N���3��P���htS3�.���=[z�U"(`�ޛǅ���C�BW��)�Ԁ�M�|
N��[ y�y�2�r�𜡪l�+)��ꧢ�D����m4D�;����I�y���6�;B�4��9�2s�Z��a6��`��c�̙��<L�7fж��VuC�5�w=��<�ue��)��Og����L��R��9ɢ6�N�u�j��!�B��m���ꋆ�]��kp�E�v�@[n8K`Oi}�ǒ�K�E����pT�<��^kA\�|�%km�b�� fz:*�=��,�pU*g����w������Ky�K�ƨ�w��j��!	g����ᙴ��P��m��0���:�u'V�;klp'�Y�$�HȽڡ��P�PqC�V���4KEB����4g[�#�_��c�*�����]�Cf����M�-=�����#���7��7�+]�i��q�H�[�ռ�����"���AT��2榣^���%�k���+V�s�uI�8�z;ƴ���֦b���m�K1av�3�k��喛�{s��3s���M�=v���}��x3^#�B����-�,�'�k�@��;�q�D>�*��Y�+S�o��@t�)>��r�#F��4�����)���	(smC8�A0��y�a�%䦬�#۹�R��׷-Jop�K�wy|�t�p�?<j�J�7|�^K��΂|K<df�`��F:>���h��G�W�HR�ui�_5H��g/�:������j�Z�Of�����kLtœ�����Nq�;b�þ��g���8E,��̖�Q�;���0k�C�&��+��s���L���2�2�x,|���-�4�硫��C��W�������_�o���A����`P�G�D�&��ld�����m��u�21�n�<���_�;$ނ�pM=�=[Y��d@b�m���ө�9+��<ͻx5��)�ϭ���N���v�V�b�v7�o]���M�H
)��:w4lVh�^Ets��<&S�Z���Q_	������P����1��h�j�,F�4�9E<{�{EՌS%#b�ad-���'�h��ڳ:��&��z�|%z��D����)�T�DXt;���*���B��d�P�wƶL6�t�iK9U��s�F�wn��Ɖ���BT��-vC����)���Ymg���MR���+��V�D���_]��[�c��2�Yz�Z�Ƒ�Z���tM�n�ɌV1'�iN5��1��j�.����o�?�1b1�A��B���ᨽ�ӈq���~5�9�V߱L���9t�f��昢 ��aĊ�c�LM�Ψ.	��O���7�=����/k��c��gB֖׎�8��ڔ{�D��*����֓P�C�j���)<KD�Ko��ڸb�A��p��]�=� -`v:7��<�}(&��J:�-/%��̳�?���I�X�z���d��kkş�ߛL�� �l�x**��y�X�s��ܧS&n��q�jg��ǋ�m�p�\]��S%oe�b��`�݌:a�H������2<)G;k��%�4t��=�6P��C��=����������p5����
~Lz���as��m��f���%=oczک�Y�Rn����I�L��a��&}^~�!�8v<�4�_F˘�.�U��-��|-i�X��A9Cb:���z駹�_��G��6����8��NH�A���0`@�R�e��PB՘� '�i�ۣ1H����������tD�i�����򚝻��1�cO1�A��� ��r���O"؛�r��+�e��Oqqcp��L��r��/X�]�ɚ~	����Q%+Ըb�1��
A}�)�:V!��k��v.=%ďf���GC��	��=C �y�P ���̾Gf���Rk��NP��g5�\��ьM���kw�c�[|�"Y5�+0�}w�K(q����?� ĀČd�c ���=W��ڔP۬����
*_�a%�;�-��=�M9-�O~�ĳ��o���D���ү�]�v���[,B1�M�U/�#ZY�K8�cl �zu���ؠ�]{�}�� ?~�gc�5#r�m�,�.�r��*3��"q��b�b4ON���\�&���H|�%z��oAgFWV�SK��e����i����	炊�W2r���]a����)�Z���T�h�d%2̊Ǳ��xZwR§q�쀰�w�ϧ�)5��O)�c�7�g���y�N��.�8�~��&Q3[�ѯj��/�!��B�6kϽnm��Q��Bn�_�sg'����+'^��[�LQ{��ٴ%�S�E�.s�A���Ǡ?9M��S�/U������4�;m�;�l �dw�f�ͣ	��kV ;��>
���;+}� �0ii#��3�N{=o�v0��2)��z���ϹN/T���m�<��3u�����`�¿4fwuעM���;�ѿ�{��2����*s��E�xn�W����Ӳ����[w���&~��߹�׿TG�`x�	O�s��6��W`?��:)��gZ{���:��$;���6�(�4u��wΒ�Z��"��(�A��}��:�+6��X�ӡm���l�uǦ\�`��M�� ���i����w�V�l�}�iP�lm����r-����ёة�j��D������[�i8�|-֋�&[�ܕ;���O�����)�^��f����.�һ�+;���^�i$f����=g�G)��y���Z��Q-�M&-��v\[�\�gsx�R�+I�����;j���o�TTUe(-��v�צ�ަ�Ae�f�QP�|�>�.o0����fe�d��X�X��8�@��(C� �����j��Wq���M��eWƱk�R�$3������Yỻ��۫��\F�@ѡ��S��3�	�r`��I�ʟ�oxK�,��0��j�/h&�Y��Kg��oYti,�~��G�]���LK����IID��r6��Z�K���Fz,���H�m��ʊl�[tD���xWL��*q5y���i�f��T���e�S��Sy�m蕚���|����W��ݻ��g&w�NZDXq�8$��Z��Uܬ�)���,V�����R�Z��Cj�v_T,�r�`4*u=����
� ���t�¡Ħ->��I�n���J�]c��t��(��5Ժimk��{��L�Q5nJG%"ڤ)Ь��Eʖ3V}��M�	����N
7t,���tM���2�J/(4ZH�^�f�zX�T٨R��{��M�h�6�ߑ Nב��`,{n��\T�y#0˲{�0v��Gxm�|�-�@gvf@&ĕonIbH:��m�zbC$����H�h�|LYJ�uf=_WWn[҄u��p�/|�P�C-�ҝ�v����\�y�2*�)��t�3�T��`d�r��{����d-A���Zk�W*@u�]����Q��!0s��5{�F����8κY�0<�9�� ��uë��8w$�vWb;�m��9)ع�=��+h�z+����j��>��&�p.��;_,��|Q'ju5�gA���������z{^����(���������b=���EK��]��5����n��a8)Cf�*���3�Y�n�,�c��*�\�����o��yԷ�N��|Ųw��'�&j��Z��vXZ3jrȕ#�-bu��&q�m�;��h��(n�{������3u�����R��D���B|U������9.���B��,Ovr	���B��`��*^��*us
�.�9����B�r�Dp�J���"7_Y�9�7R�&�b���y�h�bm�B�uq�[�S#�'7x�X'+7��)�h������K+�q��m݇�oY{gzK*%����7z��t��ف�/�i-g�s�7��N3	R8��\9����ǶҺ�VB�	 ( а��y}|y���5ppT����恼�romm���,����A��
�(�@x/AH�hTL�V���R���'���Ƣr�f�0P�lEW<��˺b%�մz�:��P2ˍ��VM��.榧��'��J�+2��F,]0������C7nT[u�E1��c5����7��(̜���������#ml�j���J���1�T�j�W�Lb�ֱ|GN�Q�����NG��gr�q��P�f-��p�KMSZ>��D˂b��e\�U��a�]MOO��ӑ��>l��o�p�[/�U}Mej1�X*�U*�Y�*�n�ɹ����_�����Q���\��]6�p�۱ESH���~4w[�p�c����4U,IP��s.51��
���Y��~MO��8*w�bT�X�i��Y�b��Q��[D&V�����RϦ�������ڧ3٦f�f�p�Km�o�ȡ���Aw�ƍe��j��%u,����䪛�X��1����Y\���Qq�+Z��%q�)j���m
�cTQ\��U�Ƽ��j���6��O�|K'6��H }i��f��aTZs�&�7���;'$�O���@(;x%��5�3�+w������]6v��k:������ km��A�Nڹ�tkTO�C�2F0�H`F$�H��;���c��8���߽�|�a5��g���2�#K��W�~7�>_j0:��0��u��.�O�n�^b�Ȏ|ZN�y�0��n3:���k|�"C8=W�'�dd�M!���M*�x�H0vW7��n(�@sl��݋?��3�$tq���oWR�g:�gxs>Sc`V�h��+V�����a�������5�`m�o�9^�{�pQ[���q�6��b���O����Ɛ)�t�~�c@�J��U�]r�_��/�U��'�`�JՎ�����G3<�kMV�j|���նp`���'�{�I6�K���)�N���THv�hw�P�b/9���0��]��l���US�6��>~���By��QC��ضg=�� �LJ�,a�״�W�{�(.�<��K�$O"ڈ$�M5n��l�yM�\=v��$�ż	d0����Ee��{�� G42�v5���l��Od'��j3��\΍�	>֡i�6��/���O5�$nĴlv���}1V�o*�V�V�z#�3�,ϝ�Mļ�x>yp��-V��g�2}p�Iku��앆�,�Q��j��{'oH�V�?wq��n�nSc��:�ر�P=�vv�wݛ|�z%�ř�.)��Jvn^���z�:M�r�xn��gn�mQ�jpb��n�<�}���!كe�IWqvgh�m�s�����w�Г�2 �11$�`F0 Ā1���_~����P�4����˺�P�esP3����m��L58{�eۂman8=�:���-�k|
�T�JJ6w���ɖ&`�m�7�{!WU�p�tԵ�Yq�֍�~/��'qd�B������u[��"7��S'y�C��6ƝA:��𹇷�kW�md�s�*�%֌���χf#��m�V��EW�����ҝ"�t?���7F�]��؊,G'�ٝ�YkK¶,H�W�>�>�ͦb �G�_�ⳤL��o����_G���ʝ����OJ�����v-�M�!r3��H8�[H$��n�|M�CAV�}^���cj��_�<��/�eh���ťt���H�0���hL����;r��q���@}7�.$�e��v��<�5f�����SZ�L+9����LƘ�2�C�5�9�v8�s��Ⱦn�ō�8�*���7P����e�#�)�E��f
�$q�[y��|�x�uAfS�x-����=XfuUK'ꖑ i�E�֤0�#es
����^˶����E�&�X��<��;�Y6x@ޞͱ�����fNP�>�}@N��ڽ��^ȅ/� ���n�&��[�n��X��
��(�@�b�a�;X��
y�j�w31�]��;W"0y%02�����{�M���&ګ�Ȯ�� HF1!�DS�Rc�j�O>�?��U_ѐ����d�c	���=��]���Om�x�4�l"��=�&'=��2_ȷ^n�CPL���0#����fLy�n�mo$�J��s�^J�r6�M��� ��>{~��a�`J�=4����_{R�q�n��T����?}(V-���.�^]+�A����;֩���T(�i㈆V���n�m��%�:|�4�U�۔}��+���>A��?p@.ͫX;�R��K��*"��L6'�����g�RY��`�]���\i��"Q^Jd�n�kf��ʛ��_P�jq�<���bY��v-��-�qE[H�@���}���~dGra0�1o*��U�Sl�E��1�e�ܾ"ފW�e	6�aq�J���vE�F��6s�a�m����-	����t<_nA�;1j�OB�o��9�]-�z9�;@��
E��	M�y�7@����}=���ܦ}�����<�D����oco_<�lS���l�9�gOf�� ��s�/�C29���v�YN�&l���W^��'~��{�'V���$�uc�n;�`d�s`3��h��� ���Y]:�cF�ٿ	����V[(W
κ͔W7�_S{J�i��g"�"�갹�;[��%�*`��c�hY��wce�b�\�1X��ܼ��Ż�q̺ŋ_gGp��Ql�i�s��G�@f�@�m�ص�A+h,��;3�gGv�C���}�w��i�@F��$��!�����d�c$�$w�VoL�+A�?:ؓ7�Ҏ����4����|1�&�1c��ᷠ4�n��S]������s`�^�)�4�iM����jk��O��8`.��ڂ͇��=Ҏ7�qo0�F6��������[�!���s�4�d��KCe� Q�X���{��mW�O�����_�?�$J]9�S��c3��M�<蹁q�D0�O#p�c���ų��F���so�f٦� ��T�U�҄/b��c�>��hf�K�լ��rg��՗>�q�p�&�YsH����u�"�u1u�Q���b,:��]��x:�s�~L-T
��w~��V}���
��8�y-[����T��E���cϞބJnR�>j�Y,Dbzw~0�Z��k��ܠV���֑��]};��P��5�fy*��<f�ࣝ��NhUf}j-��
`u>_
��^3���J�6�9�{ \��1�Ɠ6-\>���m�Йcn'��K I��(�j��&�Sl����ͽk�Njf���/?���e�;�o����17km����JmУb�?K�j횋������ ��I�;k~�o>Ǎg� �7�g�5�8�;�q�][�OhB&V�YZ�A��M��xŃ��'��r4r}��k`2�f�ۛ�G�s��,s��Yfs4��,�x�wp��m�Zi1G�;��=��ݡun�$�Pcꪯ~�c$! �I0�1 F!{£��w��I�Ck�h�3�ꇾ�oT�,G#�����L_G1{�c|�N�w��-*XP{ˉ�H<�C�\�F�Z�#�2�P5��s��s��ε����Q9��(�s��j,�r'D�4������e`���z����K��Ph:����V8�-��p���9͕[9&����`U"S^` ߩ>�N�GM\� �ۣ����r��f;�Ax	��#p����7jZ�f?`�XBo��	��$|}�;�x��vF�M"�G��F�
�!)���Xb(n��>ի�ZbGhf�E���t�Z�iM�d�>�L7<���9��Z*��Vgl�ض��+��/�:�.�M�$�f4�qpU�Sz�n�07{$m�ed?UJ�8ѸwEN�V�[Y��M;	!.��%}-(�TB��|g����.[����!�jH�.L�KH]���q�fy& _���/�F��e��AԪ;<�:����ۅ��S_@wO�\BX�̼�郲�kD�G�ܲ����UK��, .tM�cau��E�^���=�f�_x�С����z�8d&�j]i(e��o��f������R5�#�W�Kyk�ݽj�e�Q�wW�U[cr��ܷOy ;4u�؛ΆG��M�|�l	z���˿�����������~��HD	���$�d c �$c �����\�cshK��<�9�a'�W;���)�u:;�9�O,�6��fsWbw3H�~�-9��N��DblnA���z8�CڷR�M�C�S�i�[�{}|қ4-��
ޱ�5݌[-�u�b�S�G�QG�m�>v��E���K�_~6���hF��u�Z�,]�ur��yB�t���/K{$^�t�0��\��c���_K�b�`�3��Ĩ�Ƶ�k�=̩N��Ww�bu`5�.l�q庮D� ��FV������0���{#�YLv�)N�&����5͖����W3�Z�|��
��eGE=�V��(�͆:eb����7�
&})9{��_}]NV�	�1$+5���5�"�Ew@h��I݇���]m��Rul0:}.q�����J�N�\�\).�N�w��FK����)�X
\�u0=,6�F������$q�+l>lu`�z^����L�G�1bE���a�L�:M�/��Y�y�evl�h�F��N�Z���7����{X.�QFy�9�����K�}��D>&�h*��q�Xs������nBccZkE�P�}-�<a����b�n����ϩ��=]�W{��2�01[o_cަ�tɫnyޢ�����oQ��4U��;}�|O���mv��<�W)�j�TѴv�C�+0�u�+^�%v�MA/~��<$﹮6㣽l�63.������d!�D�I 1� �I ��	2B@���{�����9�sߧ?�.����O��c�a���_�z�r�`u�'~���7��U�M{Pl	�3�9�b����r�H]��w�M�g��>�H���@o�"8�Q���߳W�-�f�D���7un����ۈ�A��
��:�+�^�o�W��Y1�G(�5Ƽ<v��� �9d;;��
�{����}Dx�G.��L,E�&�-����%����h�A���;���QD�}��g�@��]��z�(����p�'��m�m'"^�ޅ���U@b�O�v���9�n����\�i��5�J�����<����3��Lc�|E  6y5�l��SOF�B�����'l�b/pR���aq}�y�R&�
���u���j4N��N��q�!K;s���vWC9�hy^�m�%��p:լ�ݨj�>��*�j�ݲ�������5*4��F�`��fs�����^��ь8�[���B݈D�_�L�̱��r������Ì���rL׳�c�c��f=oj�T�p��M�z-�b~֖׎dEr�Gu�����E�jv9�ȳ+)�.o޴�����]�L�Ep|5N"v��f��{|�!Y���~~�2����n�����u=�������
���m��:ULh�Upի�d��\�8֤�_u�w�������;g�<]hyOP����x���}@��"�}i�x�@���{���x��I1��$��@b�@�>���~�(�)9�k"L|Qx���DG�C�U@F/v^�P���inyM�\�jte�ެs�\�u�IF�q~`��]x�ޟ~�՝Sϐ��e���_����
k{�xʆhfO������%��#�6���{gm'��w���cr�t�g���q�����Sa�>_]c��B���ӎt����N��.t�D<d/���l�g�<�tu�蜱MHJ�j*
0s��y���GFR)O���rcyq�cZ� e�pOL.m��/,�dpk�gu��/�|�f��n�M�ŝl~M]��==��f'�D��p_|�VF����5Ր�ٝ�`�q��^f/���-N��;%�'�޵�=I��ŗ��M�|����]��-[GEeu�鐶��G2��b+غ�\Ag����>��r{$�UG���\V���C��fQ�Z熺j��x��z�p�{��S����q%�I�磶<=T.=҇B|4��І<d]C$#]oVc�9#��1�:�z�~W--�&��FĊv�Ha%�3�v�c��z������/D�}=�L��b��*��+�ѝ�S����c/kl�vv�|j��kw��z��!��x\���0K�E�1��� K  ־��j�r�Y��� ��,-�5n#��X���_!O{Nٖ1%�[>�hV�ϊ�\�J��-�y����G5Zѹ��5s��'�I$��$2���1 M��<�����O��^����w������:&�=��D��j�b#ݏN���\��舷��V .o!S�вІ�g���yкp�SO���Es�G(r����ș���z6tN`ӊ��k��Z��H�vj b���v)�2����9�cOsǱ���O)��["����Obu5��S;QCUØ苇)P/��y4d=����i���->���[1&�4�] �`��'���m�Zj��Q�4E��z��o@2F_#��)�E>���	ޤ�]��v��V2���S��
nk׼ݱI���J���0�0��h��N�����<�4�K����3E�(-v3��d��Q���|�=y��.��m��ȳ���<���wO
�7L?N����n4�pell4���Q���r��e��k�6��ت[�L)��A�*Tgfןi�w�`V��k�&r�$�,}�Y�"wT����mMV�=S�T�|�݁L�=�l�jg�3�A-�~N�K�o~--��da�Z�yM/�w��%�,�=������t��'+F��C��8:S"���>+��bO:fܲ��.�*o�/�B�ǚ�'M��pm�ĺ�V.�u�Ӌ)�����⹐��t�	���{�"��Զ"�(:wn�p4��sG і_wi=��u�SslK�.wM�1w��)����n׻�� �$����HHĒHc|< �u+nMܚ���i�6t�]�EḐp�M_�g3kPM��W�Ѻ�q�q�crƵFZy�!�w��l�f�|"�~���5� G5{�����y�:pš�Y�E4N��!���1�DѤ-G��FQ״�;�(	L#��]6�f��r a����X�Ď5���l�4� ��o��a��=S�|���½���@�/��J��Y������(���tOVK=d6������)�t�a��Ih
q�nL[q�lL��@�K]P�5���G|u5�y���yٳ�{%�e����@�%޶�L6�@�� ǝ(V��n;D�������5��:����M�4�4�gdaW�*�K����\��oCk��Oɪ���AF�	Q�����Ш��-�'e�W�@vlW7Xʁ��W0�{WNE��2|Y�Y�m=��ż�v�Z�v��Ӗ��𛯾(��Ì�����/w �B��+���_�r�-��I����Y�(���Ë���h��b��] ��X�<���Fs�X�|�ث�F`�鼇�`e�ށ�<=���<j��qm�,LHg9����v�]j��eU�5P�،�J�gn�� ��;#�RY�Θu�+�Y��Ss:��#�Raq�� ��N���;��F�r���frf���V��V4� ��E�h�m�*t���>טe�رc3\&��c�յk�̛K��.�g(�[�4�+������}�>W�8����������A�BS��vwyvѫ+z��u:@�{h
u�X���qf5����}ft��w{u
%�r]�^vgZ�z��A��j,�7�����톅v�T���ذ7�����7���ʽ��h�poWK��qb"��GQ�$���CGhL(��������"�W5��hW�uX���B���Y6-=�����rgt��XmpJ���+GVWW ,v�ˣ�p^��V���m����6��z�۸jvU�u6ou���ג�j��yn� ������dAi��YZiXP���6Fh</3�T�u,�v�����0t:��prm8�}n�>�ct��cfݚ����R�x|�w�̾��{�)ev�V��w��Է�s����͇����g5H���[j����l�K�:m��$�]fkzM=�])�.��_����^�˦	�*h��y��JtN���1o��r���2����58E�l���^�Gh��k!�|Px&_ ��0rW��ԊAp�ʽ�)彸�^���Z�:}4�Z��
x���dܧ�<�(Yu��E��u�E��IFG�ͅ�.�2�2�O���WE�&��V
͠+&�o������^�p=t'�GU��x��`m)�@��k�m��S�'iV�;��\��Ngr��ܺ⤌���5���NK$e:�����\��;��腇F��CH���9|q, ����Kr�pIN���|f.`��ff������j�q��EN�b�f-�����pk���X:�ի��).��e��7��ʳ�u7ǤjWi�����m�α��#�7)r�w�6�Ҹa�%	��u Q�VGC�f>��ř��(ù˺��-gf�\O|2G�mbܸ:�V{�b��;3�wW/_U���k�3�	���b >W�`Sp>s$u��nV��pv�ZLE��ﳳ��
ɨ�3aAl՘XYb�FJn��zwS����V���j,5�h�
�O0�<�ҥֶ�Y)�7n!ٌ��}5W`gD�	KZ]w.�_"�g4.ja��Η-��P@W!ujV�t�N��¶ﺹ"�P�} ��
����hŃ(���1_w�vh7���J�]����ҹ�f|�WK�S)��`i�sUE2̳�3�v���0ܲ��F�-a+�Ic=��i�ӥ͜�Ұ���gHܫٲ�L�כ�����(����Se-�+R�QUF�����f�+�ar����JcrմfM�MO���`��;�
sV,Y�a��X��h��1��Q2�����Sb�EQrd��nzrV�0�*�j"X�%�"�mU5C#M8b��`�i�q�2�{3Af�'f�g!Y�A-�#ZO�_�QSI���1Q��(�'�Y�Z�Q�TP�i�m���������GbU9�
+�J� �iim�j�\k]�ڕ��*\B����+m�rTUEDUc�'gf�g'(�2�RȢ!�Q
=j����F�JY]SV��ԫ���J#��m(d������\V'l�q��X�2䍡��V((��TEF=�
m��fb*%[wsZ�'����3�71X�PMZ*1Zڛ�uSiZ�j�h�Gn��Z�b����f��a�s��ss�����ݢ��Uq3�`�Ym���i�˘Zե�,[j X��Wl��T����ro)V8���nDE�r�jnԖ�5�U=(���)ZҖ��X�b��p\���,�����\p]_��m��wv��;�(c�����<
�V���5��%��Yh��>�}���C�!1	 �I �BA�	$��1߸}���6A��I��}�:�l�,+�@��Dk���7L#�;cN�(X����'��a��;���-��3�����H�sZE�&��@ھ��>���U>iw�rϱ݂0��eu���x��,�%����͌ ϝ&�o]���3T��L*6��������|���0��8��	��,0H���h�SO�l����ꌅ���������+��P%���V|��IP�wK�O�83zF�y/�<��l�H��6G|i�g�g�	��֛�f�
Nj�D�0��c͙�P�{5;ѥ����t�c�5�9͎ś;306�=�1���B�G�=�cL1MdG�5��q�I��v�i�qD�)�e���uF��8f��o-��#�Z�S���:�uv9QU��·VN� H��6m~9#x����4j�z�p�nʼ��ަ�of�Jr
J(�4�;c@fp����۹8�����a�U�[q�h��uk$�.��S��p�ã����im��ח`��Ь���ϧ�c?����pn(>��~T���0O�'������ͼ�֪Z��ے���?[��a�[ػ�=Zl��s��84٨��t�8� wZ���E{}식��ۃ���u-�yo�:QQ��n؎����T�W�Li}8�j�4�N����<1�H�@�1 #��||<�gUfst������;zB;AL��vq;��zd3�[K5hѦ�X�1�3��n�c�7QW��fo�6������&s���_(�����V��I+C5Sk�kV��j�=��7V;���f8��NӍR-���'�Ӟ~#����@��.jX�s��Z��<_OQn�`<�D��B5��n��0mS���N�M��KW�t6��Dg)�wo��Ȉpf��;��}�Zk(6�J,�4�aFt���nf��"���-`w�y�����Up,�������=�;TQ�I�6�hNǠv�˖g�32m4#\�E3��Q��8æ68Wq��k��[{�Z'qC�J��m�l�Q��g6�;㌀Yk����ٵ;�Q8�����]u]Z!9��U�ك#�n9��'Ӷ�Ӹ+1�\y�+?R��v,c���K��t�(�Bir��p �W���v���S��5N�i�|fƱ�EZ�צ�c	��[�����p
~��n-���jM�,����l������W?d��.<�~��u�r��~:�G�����eր���.��iҡE5t	uϙM�PT�M ��7�\���wh��(g�z��D�J#E$�̓5�kK����oW�y�Vl>�����S�;�h���+P}���0a�x��89����&����խ���-��r�c�.b�1s.�$?��H1 F0$cF2�H�@�� @��t�W%��h�Y�6;�(�a����3�kf���Hc}�/��4���Fb������7&3�,���ry��	��Ѕ퉚�5ǰX�fc|X�������3~+��19Y�V�
Ӓi�\�X���k
��Bׯ�� ����DQ\�y�t�5��	,V�g3욄a����M>u�aذj�2��.�N4��.U]��5� v:��	S@h�R�X�O�S�ͪ���9w�X��̍���mIy�L�_� NE���X��5:&ۓ=7F&�"���z�����l��&��9��#�Rg]<��)�@��*��MP�B��l[ xǄ��F�ڮd�r��ܮ�O�}{�';��Rwg+���<j59P!�C	�p�oEd����dk�^�Bl�mm[Ϭ���.��s���SF��{�i��e4�ǲ�r<ÚM~P�6��ȴ۬2��ÃG�	 3����N��5����G��m�x#{UGCOc�A�&��s�}�y%\�S��F�FĘ�m�� �6L��U��P�,�k�\��<��o_�8ҫ��#w�!�z�`\H{!���|��v�a�2�I��E�N��ՌXՕ�O=�͉�K憸�D���/�ݧ�>�����wV5��+F3�*yΤ7�R/�F�ky>x����Ԙ߰#ԟ<�,��l-��ul�N]���Nf�xv���qr�6^o�w�6@'�d�1�����$!1�#	'������s�{��^��?s9F���������n�%�Oo�둞�38�E���ut=	���a�hB�x}d�Xcݗ5�0s[[��#n�k�G�7G�+/&�T׬L��)�1>���3*٘�`��ގ!�\����-���	�P��2�ditӢ�����K���Q$�����h�'-��݋{�1�p�D�``�l3�a��x���}�� T���P����8���\F͘�'�m<H8m��p[9���AR/�ʽ��ބ���s*�aP�ѻ�������KTm�m"��'�Hב�7s�m��1w��`%���+3���yV>��ffФ�䣑]f(������$Jc��w��kC6t���B�4�3��|���o���Aףb�����!ش�ia���m����U#���%.�k��<��Z;�1���z�� k�K��1���k�+����B1��=#���h�̓� \��+_%h���̒�f����#Ƭ��0�w�����1�@+T��<��UC)��lj�v�~K�fa������D߳O�w�6ɃE�<=n�N*��m���U.Ţ���׭�l1��gQ�m��g�ʃΉ:Gy�ket����vv9�Z�^uF
f��or.�5m��sO:��N����o(�;���6?��Ha�$�BH� `@c$��$'~������~�u�7�"(�0:��!�X�3b��7�3�	���)��k��ޕI��^�\�2w^�z������	涟��Uߜ]�W.Dz�ح�^����x0��a�wۣ�M���ܜ���[x�>��؄�-(��Y"i�+��>��}Mg�Di�@ǽ����%=.;W����dő!����*t6;jl�y+[ygϾ����qk[��!���ȁ����@H��N�e&�nkM���Ј݇���0�זƝŕ�DT���v�Ws��s��{.cΞq���:����֋!���t�[�Q�p�Y\�Ri��հd�&�v��S���Ɠ���bD��=��P�}a�)��~d.�OU:��D��0&F+�O|#��v#-?�e�4��g ��ai(F�g0�I��q��-�������n�p����_�2�B>��ʆw��S�`�C��;���X��w�ᦃ?@f�z�H1:��r���x\_I8k)O�$�*9�3S	�f��}-m�:`G��C4�j�xy׿E�\�F΁�������h�yMʤS�d��=����#��X�{&i}�v�3�͛�}��m���sƕ�0�tw7������^S����N�A;� �Z�9���D���ް�m'����vuS��a����bHF!$cB���I�HI�����ٞ��������;���d1Ʋ"�Q��]�/�$����u��#��jw��hΦ��wWY�85�"̆�z���rp��| ������*j���l2_��i3fwb�٦~x�\��n�[($BH���"��T��P�P�cI�Y�>������%���nz�ղ�y��L,�i�5[��i�d���o��?��.���+[Hg�hS���@�>��a�s�Y�P�lT��B�E<�QD�E����mX�����.�+%P�!{��X�*4s���ߖ9��{Gb�������QFFgA���?�Fإ}��]
�W+�"؝���3/g���\��%l��q���h��Z�'��do��Zg�#�"���2W5Z�(�U6A��olJy��͖uZ�2�����O������1�ogA�Y'�imx�DW)�wz^X������fgS����y;���Es����Y�N�7�yNz݀ъ�����Z٭۫;f������e�מc��j�};!(V�j�1�a��x4'�>U��Mu���g��;�.�~H�oh=z�5�ݻ�U�]F��NŶ��>��䷜��t���K�Z�&[��@���2p;g�1��Vm��i�.�emq�MqR��a	�Ul���v1\����Yׯ�����<8-u�Dhn��;�a���p׹w���{+�h�f�e	�p��l��!6����I�F$�b@�IĀ�F2c �����}��|o��Ɇ�륧�}��{˔�i� �4ߕ�N�v�&��lfka{Eְ�-�^;W7?l��x6�_\��Pg����++�`�A��'��{�T��Xjϵ�9���'mϮa��o>J����2�jk�Bq�h8`=�I������gS�S�f2�7��Q�cS��n�>č�͋�aŢ�N�K��C0ZCIO��6�旟a�L�s���	W��ߏM���.�T�Q5g�[\��J��i�q���s�����q0�5� �
X��6�qg	g��j�(�/�_D6��/gd���c� �;���rm�p�ê��5K	�؛�ʊp��`\CW	P��y��hÎw,g&lÚ]�Xֆl$���Y�����xђ�����pk)�J���c��oK)b��7���{Rao!����H�'3��d�r�3(Wiy�1���p�f����LK�b^H�����<Ϻ��y<�U,F��w9:�r�h}U�y���������o@�z�&�bh�q4B����2+�
9C�d�\��/�uǖ���-*���쵝��i�Z��Q�+k�}uo��A}\�b] 㱓dV-��F�Sחvu�\�T�wݥ�,���8V,̽w����m�}6����]t�So)qޱ�\�?qg@�4�m�����GN{�t�C�2@c$2@bHHA� cI$??7�/�����~�r�VCA�vC�\�ٻ;P	�a�"��k2����i̾v
Ҧ���W��h��7�I��V�hr�sn��C���M��x
O�nr������[N��?5f�ƫ]�\t�7s#��$Uʹ�0Ϊ������j!��1��)�-N�9�evR���m9�%M��w����y�)�/ܤi�]O�P�^���B�e�u�]C(�� �v^FS���L�L	��c5����Z��T{�=�a��]u#����Y�6Ꚉ�/7%�k�ǚ��nָm;����T(g5��#i��Z�8�a�=�+5�L6`�}�y��i�`٬I��3�z�k"}Q����	�j��s]�8(D]'�ɷE���;��o?7[�2�/fƝ�h-��hr͑�rKpX�M�|!��y����������z���^�QJ��%��E�Z�=8cy�7f&��f0�E�ᔶ�-Rf7��B�ȴ �Ϋ�o��צ��#5��Y�=!��������ti�ՌJ�6D38��Σ|ϖnkZ$�T�3����3cg1\��6�7l��;�f�=ݤ,�M�w�C�i��\��b��ő���V��� [5�=7�����R�I]r���W�+��;�3{�Eّ�G	��]����u��*w�Ō3n��o�$?��adb�#�1�#�1 �|���_�~��������z94rty�6,��|�;�(�1�w��Y��9��V�wR{�Fn�c'u��s�	�燳��a��%�o]>i`���o������35��*��R�i�Ȧ;����I���s��O�/)8{�4j�f��$Ga�s�ǝ�ܟA��(����UQS׻l��[�d��	�D���������J��~t00-'T�^�h���OdzH�'���vYť���gp/�����*�͑&|T3���p �x��o@ւd�~�M�:㭝���j��h�(u�}4f���g��a4�l%yB�6�QX�g10ʂ$^;���X?q�{(�|��ݟ�s>L��ĸ��:g@�u��>IX�MUY'�uT\4�kf�5��c^z^���*��+�2����pK�O�����olQ\ܘ���=T/3n�$㈹�%fl�ݍ�|����bh�29��AZ�-�q]�t"#4�c��Xn�ZʨC�3M��s��nk��fW���]��6<�H�8�vtra�9�"�9�s��_3]LdUϳ�P��Ł^���ʯ �ZoT��=���W\���yȗ�f�l�wW�_+
�]�P�G�`ٔv���eh��ia�i={Nk�l���7�K����D vq{�Q\},����j$��U����A�7HsS9l��v�5;�7��]BE�͖:k��Z68��;����@?�H`@b�2Oх� c ��w�����~���m\Gؔ"����!c��[0�{��މ)���$��y�m;��~�Q����r[5
�B���\�/�h���.�G��'4��>-����9��T�x�b%<���wn�9�ɩ�B5�>4gr������83��<��blq���a�"���Z�������~9� @do��6m��8ڟ�;�����kl2�!���Գ���o/Q}C<���M2lP#��i�C�DPj:ԡۙ��1s)u�;)]�&�{��i���ѵW,���*�� [9kd��b9H�u�Qמ����yM����?{z烺���͡��Z[C�2��1�(H� ���,�Fóa�n>��'獋�v�{?;n�<���e��MXf�Y��M�a�d�XBR./={� �R�gb!�(�1�?��~9��job�\��׵�)�i�sb�Z���z}ʦ�����O��(�d�4�,�_�s���-�o��ˊ78�n���P �,�ouAƚ͉+l(��JzD�1e���4<����0�WY-O!��P�o5���㒧]J����RHs�Yp�"5��3r�Ƙ jv�".j\E^�!=��}�]XOk�R2Jә+�$Fg
Rq@s� �-l�n��nu��[��.�zݞ3��B��9�0f�E�wDb䇓ݧfa����ř�#�*e�(��BSP��B���̚S��һ��C��Y�.JK(WZgF)0Е���J�	�+ս;Nl��P֎�� ���[]���vW�y�N�׎NMm.MGX[1Q3]k9�#��|�����)�� �y��x�+(�G��7N�u*�V��V\ky\�Ɓ����(�z�n��bd��ݩ�+�&?8L��E�	��)�0���y��,{\���;.�V�\��]��1»u]�������[ U��{�������yV��{EV�#�� �X
�����H^`{4حS�q�5/����x�64s:��t��npfΕ/�fV�V3z����h�î��m��Gi'b��D�Uie-xh�����Վ���YBۧ*�<�%w�l|�F� �kr��"���.���4�X����������c%1�N\yu�u;̶��ou�9��H9��JNX+����[������W����@�Rk�WiWc��6����}]�-�`�m�utx�GL$��$y��&�c�xv�"j�f��\֜��]z/.�i��k��[�%��\�����G�~�f�b�JRD
Uv����}%g�
>Y�gw0�"�2v��@���m	�b�T5I�f:��t��7K�,��A�NE̒.�L9��c��mQ��Z���7$ب���j���ܻ�թjŉ5G�4���T/�����:M����8+�86�V�w@r#�{bK���l^���:]�A�۠U�gC�w��[#yvmu�¾�
G��-��&G�K=�m���U�����k�����+��a��gh<mi�+m�.��sT��)(Ք���~����d��y�zg^^0�A��q`���]*�=|
��;.�*)����r-gp���5��V.o�Cw;�J\X����|���(�M�K6oP�x���l�I)6,kl��9ns���̡�\��U��eݪ�$��D��G��1�C�� �A���8�<0�&���G<���SN�y��Y|�L��[�
士�����}�j(��0���SrZ�ݜ7y�6����WzS���2|1iJg��S8+�}}�T�*u���wL޲��r�}Kh%W���~�jA[Ϋz��$=�w�w8������_���˴>S8�G�ֵ�Ԥf:�&.��R�91)��B�8�ᒵ-��ۈwq���,n]Z��\ݱn�6��o�GI-�©f��tՓ����y�ݢ.�����WнY�H�@��&ƥ�V!�ʂ���thd40DU`��
@] !T�X��V����\5z|����a�?=T�[,՚nQW�-�mEjU��T�VZUƢ�ci���5��_���Nϧ#�^^Z����F��hMꙺa���Ģ��k^<��3i[���ඕEQ��(��S��~M�M�m�;h��Q�e�jF=Jj�ˌ�&��j��Tam��Rԭ��ϧgg'w�U�73�Ԙ*+F��[l�Mb�1ٔ��A�bj�®Q-A��R�OM�MZ���.}m�T��Ud�epT�DF�3��Ԡ��	SY�bU�V�'g'gf�#DNRU{�25�j��QR(���*�\k�&1be31j锶���zל����ӓ�yeb�tč��;��;��"cP��luK�k(�ݹբ�k�ZY�.ON�MM�AE�*A��L�N�qqLj��_�Q�l7kr�S�J�㊪�+\ONNM�q�*�������T�ù��q�Uә(���iGj��q��J��9!�Luis�U.�[,��)Y[mEDU2�V��G�-��\j۫\�h��ݷsXt9A�x~t8��zOb��Τ�<_pz:��ư�kO&zC��5�Y��:�uoS�l�;�]�������������:;< ��������X2F�O��HF!#F!2���oߞ�u��'~o��[����~i���B�qM}�:�n#����S%sRǓp"w�q���,Km2����0*��S�$oL
f�6��T��~֐��ȉڞ�ހ����w��v�m� U��4rz�gtQ�f �g��%����C����[���-�<�➦YZ�c� ��Z|��z)6��vWB����'dt;�m��;gsOX���0�k{1�`΃1�����I�:O��;ᾣ�2�@��t�s�g��6�9���M�k�3R�(E]�����A���W� ��W@�Kf�m�:y�'��j��qu#��&�n�j��)�&mc6�
ရ����CG2=4-��tn�����ԊS�f��u��(�dX�Tm��:��/Yw��b�=�%�N�u�M�@������6>���Q�P��T9P\�Eڻ���R6�����wD�Di^$��
�G3�P��)�����j�7���D9{z=n�>3����8�A��w�z��3<�Hnz��f7�)Ȇ7][�r'|�xg+ɻpQݐ��^	������T?�Z�Wq�Ʃ<?mu�5��8���9e�^9}um�՗ʶ���j�whj\ڦ)M�tPg���w�t��s��K���c�ᶡg�4go>��J��A�hW�b,M�-������co�	�A�A� �1��a# �������~�~�a�ב����kdep�o9G�S�t��hf���ǋV��9�,��5J7���ʒ���Ρ�D������ܵ,ms�s����U��dPՔ�'uaX�P�j:��:sb����AN�sH�DK���p&�05��ͨ�s]���H�������u�~������(OmX����C8�h.'T�V�2+�
9����cOJ��SL�F��7�N�`k��9i�S��%0F�d�ʚ����s�uзka�W�Ak�6׻ I�IM�Y��ظN�ha��y4d?(c�	jdE��W
x*��1 �j���c+C���3�!^�t0����y0t{x*�W!\��N�.������F;�[H��׷p�u<��YQ��m%W@%��Q�[j�7<�̱3�����5e�B��cݯ0�I�	E��<Qi�Th�d 2����x�3�bwa�jq����%���o�Z�K����}�Y��iI�f:E��Gt��Y�;�.kE'c+ca�n�ys������K;V�|�f2b�fv�[?��mx�
��=b%`�O1����4���
2�8'ۨ��ڕ%$�r�f����(I�W��vY*K���@��u�s4m��D!�j,H��X3yk�Mk啼�̘Ӗ��X0T���_usz����C�!�#��H1�!$���?��x���o���w���6ē`�l{!�f��Be�BW��^�~R*�oua/6]t���5nU�X����6w?�xoF��v�ލ�cm��d�8�-ɴȆ��޶�ˍ)zX�K�l'j��6�n��P��]"̊[�zO�
�'��& �vbm�[S1���T�k?Fse���ݢ�yjZ�JgP�!��kƇs���>����a#�D>��X��g�"�GS�u����CW�A#r�ٌ�2=ƏHY���z7G��G8�\r�� k�M���lv�ts�o���?N�� �T���S�j�|j�$��: �ECw������n��Jٵo�����dukX�d
�QL�:�9�����Ύ��2�X�l�A�g�����g\t#M��{7������4���_�;'�&(�?J��#�ή%s�Q�?{�暈�3���
��Z��44��Z��Ms��ʧ�k-t�d^T3�ڊ�Ih5-����`�$O7L���-w5{�m6{i�c�F��5̎�H�yM���*�SZ�r31�ǳ�~N/��캔ɽ���쭆1��u�rC-�vu4,n�ϒ��[�,�(%�*�TBgL�% B�_d5�Ϩ]��A��R
)/>���������஧�qw h��r�+��>�}���.3(�*�wXkμ��	�qx�u�K�~��^#�>00�@��HX�1 � ���^Ԥ1T~�(�����Y\<P}>�����r�.���H-��(� ��*�W��,-�eg;n�Cdu�)�ÍJ,�sn[������-��y��l�r�c��f)4v;���T�"m���3������Ìf�;Q&%cG�����@V�����w�����m7�U���Š4��繵P���}.a�򙙆ÐΎd8F���9��A�Yg!Ӷ5A�z�굴eZ�`�)J>�8�mѤ@X�p�67y� l�$ �z�`�d�{U�<\M+T���N:S�ץ
JDȡ��ut0�7��7(�k7�O��e9��#����`r�A%";��ar���x~�d"��CA�q�x�ݎT2���E� �=��`w<�֞bmv�[�ݥV�*�����Jg�����rkd
�)4�ˀ�vzXgs٭�K[GL��������f,����KްLipNcG�ם����C��g�=E�l"��v+��c��rq�ic1�h��w�����sS>��DQA���G����K��p{�<
3�H�-���lm���9�3xk�nd�ܻ�y�n��� H+TL�[�nVõ!���#�p������4�J��Ե��)��@�ٓ�-٦/
���녂%�w�[q��M��m٭kB�=XW��Kؔ��evr����s:��-��JKY}[묰+��k#���1�@�b���#�����������鯳���[�E�O7�i�C��Qb\=��ɧ���NC���[iW'�/Yoy���'Qu�9��<W�o]�Y���7���`Z׈ѿ{�Ā*�
����P�Ql�^�N�2,�3�NfR�W+��0�1/%G���6�"�7�*�A}�t��Z�:����,�k+;�w��z�9��sя>�A.A�R�p)��`'��4k1A�V<��l�'�UХ��V#�e���l־��Y��N�����4j�$Q_y��A�Ϥf;��/� ���ֻ��g2�[�AΚyՆRU6F�KӋ�vR�0ogL
�;�V5��,�X���4��0��&o��r��\�|t�o�l?D������MDy��1���I�����N,��O�C���r���A��X�[�7����O�}�R��Є�k�@�|�_��������=w�G�kC�I��Yb����H�����:�����È��ғ���P��g�5Ʋlc!F��^GB�����
�g����݇s�]e-�27<�:y��s��ë1��+��[�e!U�PM�b�-7gD*��%���n��e�G�u�o���t���]����6�'>
��u�6�5�噅�qӈ����I�Vgt��' B�Ok�ב�Xi�w��Σ@��e��дuf[��V
v�Ŀ���Hd!!���#���Zj/K�T�������~f�dg��t�{f���1��S�fMv��*f�(kkfU-c�lDZ��aب�b�W�n�����L�ό�?o]!�y~V�F� ����ᵳ�>��Ti����r���r�౷>�v��%I��H���x���;k&�(�*
�Ɯ)��4����9�7=�G�ݍ�z^	��1�Ww:�-�=hQ���W��q�u�O(���b�>:��,r����%��j���w�[A��ʟ���ڪAO6oK�y�Z�M?��T�\e�����tOt1cR����d���S�<E	|x���:я�����o����J,�+]���qAZ�O�*�1�R�B'G'�t��,x�纶�k��Ss��wy�LύD��\T
q&��sP�p�(�"��=��e�b���ʭ�Gei�Y�moW��P����;�Q.�n������N��7'jU����Q�]��>�Bf���ۋ�I�[mT�Ysn�l�h��m�Y��]����d���^�4��U�8��Ӏ:�J/h�?ҽ��	�'��&Ã6���*���e��ˈLv�-R��D׼��/E�%m�eE�?6�M��S��׽��-�7��#��8+Bл�۷0�Q���7��j���qI2�s�q��s�\C��z��w�����0Y$�c!�F F2���ݻ�����?v�jAߵ���a~m�+&Gw��j�Hê@w���,�Kl���6�=y=���F����4�{��͵�:%����Cc�\�s�l��#Lj��H��T
1�#A��Myv�n�!6�&��-���:d�F7]�V�����[˵Ҏ�;�K�cAt�s3��1{�A2���B0�q~=@K<{�L2;�.kE'r��j]_�(��}�V���_�!��⨥I�SԸ�&7�����>�1vk�'� ?>kL4s.h:o=��`��gf�eR��6�[�~g�\E�v�.�idz�ڣH��%���l����&A��::\���~Z�^�E��[��##F(�h���]%�(ȥ�1��ӆ=��_��	$Ղ٬��d+�K���k������5k)�]�#��H���m��/�y���"ZF�9�T�;T��C�MsNWS�@�/68�;G�?&}�����*@��ftY����o?�h3�Uz�S�`ndE@g�hSv��o9}e�hf�,0�N ���$�糩�XoL���,7mJ;2tm"O7�Vj�Y�x������:��z�:V�$��7JW��� ����v,��j����V�r|j]�m(;��&�1a��x�c�O[��6	��ݙ]��.�<̢��r��bgt��x��
�Lɚ��1�s��q���&s�}��kGu�q��~�c�1!��BO�u�Ͽ_~���y���?��r�j��W/��"��:kߊ�I�a��K��zi�\���gXu�v>��o@�r1E3 ˞Y�l;[s7�_�m�S��x��OޗN�����sI��A,M�IRB�~����S��tryT���DA�������r -F�ŵ7��4�����έz�n�5�5;���ќ�G���ϥ>�u�.�RQx»׋)Ȁ�a�hƖ�f��M�����ڈ�T|�����y7��x���7bl��</�wX[Lkr���5A�L�O:������ʹf%�C#��
���L_�2#Ta>f⺜!�m���4���ͼ�V�A=W[����9�;c���w��-�����1m��?��.h���	msH�E꒐�:"�CBy�U� ���=̛j���i�J��
��cN43���y��=cJf���z*�O��TUG�-��CS���T�����Dq�+h6t�&���J.�fD;�k��3R�ۗhd����*�R&�:���ƻ�G'�a}�>^N9��a�b[s ��v�o�g�F�f��μ����)��wV*p�(���_�By����,��Y��ma�֪��9��l�f9ڙ���v�O���H��Wp/���$a��tQ8n�ݛp�O�(m��59�@*��5����s�76����v���{eը�����{�]]������ڔ	�E��m���B�r/��_ǘ`1��0�b �}�5�8ʦR��b����j|֘�V�\�y�4�3*~J9�����#Lg<��9l�)&��t���.z@)��l�s� ��ф�DjOfg�4�df_��ݽ�#j�4�9P�;7�	dэ�8s����)����-��,�;�7�;�M�X$]�P��Uy:Ѽ'�!�≌��'��6-���w�9UbD��a>�~M6��J�mw�Y��1�[h}�%d<�W��͏�zˉ�� �Ad�;�N�����Ѩ�0,ӄH<��wh�9�&�藅K��K�O��E̸c�o�+�����/g���@�}��c�Y��+�8S�AR���N�k��-�C3�v�"�E�z9#�H�j��������Y����g*݈V�d�6u��JA�	ƨ
�}�B�(�s�k\�	Y^�6}�ۧb;5�xٿLe�׽�_�,&���.]�)�Z��j��4h;bjL�+#<z�x��v!��K&ٹ�7ח3�q�u�\z�sA���N����p�/�iv�)�LÊӷ��?g�u���P��e�7���ۿ�2�gA��|���k����n17KD^�[f�{>t����?J��{���ο�T�&���M�;X>.S�e���[wui���GN�"w9���ޚ�m]��3zi0����!V����7��>Λ�=�m��ѐb��Hŏ��>>��z��4J�o�[�n"�vԣ݊$�yTQ��F�s
3-D�����P���ϕo��"�Fa�| ���z�K;mQ�����v49>���[i�	�g���m�������=Wr.V���k���IpeL6��6�X�}��C�u*�������@�i��t�6�tE�9�Ǚm�y�7@�B��a�[�fm7�L\�M�0/muA����s�Ӣ�y��̼-o6��٢�4��	�-�`�u��#_5���ddCA���9�������s���8J��=��^ݍ07L�� ��w\6l��=2�o�ozM�0��V���.�;�٢��.�DA!g6��=F{_|^�^=�z��q�q�;�hh}!��k�d�l���fu3�S˲��8ov�1���6�@���0�m{�7�</���s�,D{��Hg&��8bn���}��u���+2�[U��~e,3~y�'2 ��fgd�q�����5�ߩ׭��6)��p�ueD�50^�"�{j9��r�P�`�<5��h�%�����tJ�b(�,�ޡ�=_n{s��vf{�N�d�ća=�G�Q@���wsr����T<V�Ԡ�xV��ع7�}�
�^��i�Ax��HںB[���=�P��Aw�vodѫ�
�^��u��XevM�ά��y���[��G�����Snp��p�e���&�T`GZ����;�
��k��tM�;H
�,��	M��V����DJ[��T�,��!��0�l�O!��Ʃ��=�X�Tن[xQ����ق���Y�7n�4��Yyl�&yr��^k439��N�}q˺���q����{sJ�
��(�T&g�cy�7���^Q߶����^9���9Q'um�ˋ�9�(��q��{,�����Jƫ�<�\���KE��1�j��z5���o�uX��r��+ӏ��GΜJ���\ܜ�X.�����P�f�X�wi�*'u�d�{M!t�
��(�pP�镨u5�ա�<.p{j�tw*osU�7-p�W�|�.�ѻb�*�E�,q��n�1 H�P��ψ��J���0�4&X!b;W���gf�|�n�g�Wfv��=�4'�2��Ԙ6��Okk�����Bmulͧ�:�Ye�Ru58q�3z��wj:���r��Kr0�n��ʛ���ʋ���={���5��B7��]P�������K�MF/��]��/v+Yj�7MIIkpi���su
<�͠�Ԁ����[Q�۫�C\z��w�ٓ��Ytl��
g�D�}��Ƹ�{[��z��TWk'�՛F���M����y�~�Ú^��c�9ӳ6D��,>�kyN܇N	y9pubʋ4���wW|,3�vz��I;�s%1+z��K�� ������f|�^,�I�n��v��I�ľ�F�Ŏ�@ճGq>���d�_=�J�ѕ%&N=o������ܳ�78>i��I�!�.�}�����/��'�v5{�'���쏏)����j�;]|M=�d�j41��dN�E)Azv�C�o���pSS�e��bt{_ ��C��������]�8k&�]Y����[��<�H��;|Ru��ghn�+���zB��&�v'����4f��^�i���^9K9�ڴ�W6��A]N拾���k^�mu3��c��f��EI��R��ٛJZ�[<���i`d������6��wp�+��EdjM�F���fA�svIHno6IC �������s:fnwt�Y��R;QJ�lR/��(]ݔ�\�"����*���@R.0�K��t�o�����*�[�]#g,�2���k'��2	�E>9-s���G7���[�����]z8V�}��=!Κ۠������WJn�T�)t-늶m��+HY���a�Xt����-���֢����4P�@ ڟ��� R�����m2531��Vڵ��2�-e�L�a�0��2֔���s�}��Y\�d�jv}>�NO��*VW}�sF+���n&���M��P�s\��_Ɔ��aU��W榙Vf�Ӭh�2~NO��79
��*�h� �X?'uf�_���0�us+�2�����E8��6�٩����pb�6��kF[����4���]���D���([{j��Qj�.cuj�Qd�Qm��'��g�'"i*��$M�x��&
�aV�Z��f�q���WM�utkzލYUq63�Ws���ٹ�`��_j��QSIY�S��V)>J���e�*��E-�d[e�k+m�0,�����,v���1J�)_w�Q��c���������L�UEuo��l������U%�-�Q��iJ�+�Թ��Yr���ff(���,��{J:�`�WWmT+W�𡩹��ɹȪm���b(�)EVfV�:��zܥ��Q�[i��6ٶ�FR�Z�Sm�J*���
�����M(��S�̣/2�F ���,Qf�auk�A�^[(3TE  b�������l5w.�o
H.�٧9�k �|�ܘ]�փ�Ŗ]3 ጰ�X'�@�w.;_Ͽxxxz��bD��9�n�����z���{�����I���v�	��G�䍇J$zlr��T"SE�.[ҾL�t�>�2��]�R�+I:�0��b6���^ʻ��N�y�@�5�3F�_P�W�P��\.�
�$��Q�9c��h>������a��	�a��Ϻ�F>������Ή��������Mi�6o�@�����?�(DH���ǾPUX}���G�;0ڻS��G+�Θ��n�v/<�`Y=�g�::�,��W!\��^�Yޮ�����6V��.t\8��V.إD+�1�t���T"\����4�5s��zM�C��0�`��d�1Ϯ���Ҫ���7�9C9�l��C�~֟Cp:h�F�v�֩쵻O?�s��C"#)Zq�k\�+2�ܡ>@�c�����b�8���k@�� \��ͧ`N�z6�w6�w;u�#e��1(E+����nF��1vk���t��#�$_���h2g�
Q���*�駸T�
��k^�.��?�S��i-���6� \C����6�������-W�wl�HP��u�H�����! L�ѣX��[��]Θ+��]�]C�u���L���2��Դ�M�<<�r������]k�ئU �±ui�m=s�f�t���o�RH�3z�j]S��OX��5ZM�3o�y�X~^#��b1����߿}����߿O�����Z=ѽ"gv90�J��0ժ�� GN�y/�ă���kn�Oy�يv+i�VT??[,� �'��N�b���jF�����T�>}��8@o�%�:�B��_f��c�����`�j�px�f�Q8b�����Z�|�>ށ`֕U��ÉP�gu����Ikd43b�q��=�DL(� !	�'��Ž2�n����(���L_&,�:'F�5O�Kz�u��� �tS2�k��x�1���@{t��S5W����BkHw�Sև����s�k�����wO���jyfn6&�w������Q�Kc;K�Ȝ��p518�6�Z�e�io0�m���@�i�s��ʤMז͑&Bʆv��Ęs���m���W-6�Pn�޾aCcx�9�o��*(΍�G�����^Yr0�U���b�:#m8���Y�ʺ^-1�^��e��v�, &�e=�5��7]�k��Kx,�V�� �lf�ڷ�4�:r��id9f`��Yc�n�¼�������-���o�|_o���6n� vl�7��m6�t�W|�:�R�mvk��ٻy/����Qq�=�ljz0�����;R|�?�;�`|���LA	O�Jxb�u���m���
�,$��h�|�ؒ�NN��V[�=�}	�r��Z�';k���F�>ܢ�k���f�I�G�ֳZ.���\)W��A����@��~�k����}�{��ĳ��-<�{�H �oL��z�}!�`��ȫ��Ke�5�ᐅ��K����W��eqm�#�ǡ���u'T�B�.e��C;���C�;^��:uga��q��>��##���@R�Y���@�:Exr����a�t����5�@R�.�~�}5�.���~^f%�:a��I����+�Dϫ5W;
���O���q��4�1;�A�**��}����}ȵVW� �u~��{�L���O�)��{i�v	2���,��NsƘ���|���9je�A�,�8e���㎈`l���G.a����H�~5W�̞���"���n�ѭL����d�Ub�\��;�̺Ǿi�(�"����gqh�ؽg��y*���^p��8Ҧ����XI/�3�|�PY��ŭ�÷��t�B�����3W<�>�dX�[�sRߺ������AKY�~���r �08by ��ɧa���}�6}b?/ٞZf��?w'����~�8��
&�I�n=m#S�r}�`\�N���UK�Y���q7u5��/.0۝������[-�:q��m�|3��f.�C��3�E����ʂ9)�����;T����]8+��e��E�����1��	�91�t���N�@2�I�m���K6Fp��EnU�w�m�'�޾����}ﻧ�D��1RF#b��>�^��߼�������|`:Q�a�1^Or�r,=p�b}��(%t+��06n��ގ�]u��g5�;!m,�S�lߛY�a`s�r0G��uʫ47�O3�UoO~~������;��5I���WB��ݏ���;D�382h�v�j��"�
>�^+��.���3�q!�7ݗ��4���S%sW���9ALQ�vX�vT��~��4�h2�5�n�U�7.��6�*m O�?cg�Dr�G1r�9*�l�4�v���@w��H��_���4��OM��sjr8�v�����\�[To57<����h��R��Є��u�Ջ�_9ﮃ��J�_�������A����c�j�Y��Li�+54��7(������e���y��
�w�CR���T��S2�2�<�H!����W���P �������:y�'okm�]#�x��zAuٚ4.�i��b�w�c},�pې�����%�Y�l�{ؓ��TZ����/�rHX�6,^��!�W�x�|س��$9a�Yv̀��]sH:o�0��/l��,k�S�tu���V��������jm9��=�*�R�D�u����kڏ��3jkQ��n��Úkt�
U��c�T�el�cL�\�C�Nr�����n�����6'l|fۜ�j�n����᎝�J/^_��k<���}n�ݔ�?�b1�@|O��> �w��Κ8G���P�+=��}���*8�q�?g[�DiD��H
����8Iڴ5>ti�침���N��47��ǳ�|1@�:��m{M#{`\�r|*��]+I#>�(jA�
~��ݐnW�%�d"�/��,�1���bEϠfuH�:�o,r����+a\�^B��D�u�i��f�����g1���=���e�1��`.tH�")���uqڲ��2�3kZ�a�;�e߮-3�̪zY�P:V��*~U%�\��s��َa)9֝�]@��è����[Ɯ��h���ZK���9H�'�,�EL8�j���Ù�w�%������<�"WK!�������r���T�z0,�fs��l�j�N����ve��P�*6�m	:�T�xGA��̍ch��V>���J/
Z��9V�V��LJZ����Q�ѹb�X�Zt��a�Sp.=)���۝���{aBƮN�r�Y
�Q#꨸gpy���uV�`v�����w��c���&�I�pL�Q�|��W=�)�+��$#�0.��7���sì��x���=e%��3��N��6����������V2j��h얹I����e�u��e���؎J�&��^�Eػ��3��5F�k��}��P�E�]u���vu�����֋;����{%���g2T5�{]�����`10c ||P�w�i>��U!�|�K�!:֟Cp"N�hN�1�Z�@ݘkvݧ�;fe�dp������[��G'�{�������|#Y����L����ȸ�I��{�s����Z&��=�Ze�Z�o!�[	]1�I�0�A.�)[ty՗�z�����`��Ȁ��Za��s���x�]:��
xb��(5���m�}:�idz�UN�v3Qoh'Y������6�#4�q��]7�:Ф�M/Sل������] �ȳ9i��aN���ϟ�_97��#xܲ,���'&j�%F����1�φ�'�%�E8�h��w�N4k�";��r���6F��l�x��d�8�י|5�zm$ݯ3��И9>=�88U�rh�U)�g=����|�r�5a�5:��֦}BC6b���"�kHo,�����"!E���`+�xjn��v2�Vk�7Js���E��,|PZ�N4���09T�K��SC*�8��^�*�X�����Vj��x/I[��U�lT�-f��y(Z���q���:;�q�b���a��gn�o������������ܼ7����*j��En��]!Y:�X���vE=G����Þ�7������m��GGP�f�y��oEu��p�"h7���y0V��}M���jy���x�)���h�Y�Q&-����nR��T;IΦ,a��z�1\ ֟:��T�+��]�����F1�ČH1#b���ߞ����������_��q���h��z��4���y�k� s��񊵳dI��� ;G��^��	�ai�e��1u��Vu�sh�L=�g��5���ǥ�#1��G��6�rځx5E[
8�U=�o��m�79ٮǶNE�H4j�qa4��Ta�`@݈I�ҏ.�Q�Z&t�e=�X+��q��Urs
���m��	�3�,˲+f�p/\�����\S7�ok�v\�������4��{S�Z�c�{t�̎��}"�R��n�]K�Z׀���ȵcN��R�U<p����V��>��;�a�z����㩺X �𹇷�igq����u�s������Vf(ێ���^֟Jy��+z9�H�:E{�t�K<Ϥ+h6x�wwKg=��fD�UQ�"֚vk`�ݍ�K�8»�L��a=y�}��X]zyO -3i�Y+nK[�d���r�t�j)R��~K<6����>1��!�W:}#R-'ח�IķCu�Y�-yl\��ض��繠�1� ޠ�0��1����j$�ɬ���t�Op�W��>�!�f�ab���Re��R2�hSװwޖ`*��ߒ>�b�AWz�a��V�z��70��}V^��EgC��S��e����Hh��۞����.���\A5xIg7�\ɩ>��A���/��Q�>��J��x]$�#�dX��F,C���}�����Ml�;���cf�	�}!��s���2��Ǿi�)����WMs=�b3L�n�m6�Lm��@��-��	��U���b��cl����T��`_�J#+nj��&�~�q��,c�|\
�b���6m~9=���1��ʃ�iQ���JK�ͪ�댗l���v��"^��`�.�x��c"��u������;�0�Eu��S�Y�m�l��� �`�0�&r4�K���Q|g�}^2�P��n�����K#Y����i�j��?W�GC&�&������#LG�oE<{�'QFsf]�q;԰���5�tm-$�X��-�u����H���f\��
b@��j��4�,{Zk��/�Y��6��A��9J�LFq�\FS��؃��cɹ�SdO�=\8�V��0gL
f�fc-q��ga_nTh��u{j�_N�V�&DN��wyD��+�9#�)��%��g1�מ�5x�^�B�/	�iF�!�8������xcoFsSf�&�a6������N�Ұ�#�x�?-n�	{�:c�k"�4�tq��r���hޛÑp�R���)�+WS�!�u����>���ߝ���6I�DxQ�y����L|�4[��o`��y��9bĜԕ�ѣ���q�q�쌩��ʘ��H�g��؆Ї����c*1�������-�M}�?�<���c�h�3�:}>�M�N&�� ���-��}�ձihT����=�@~q0[��H�}!��ͱ1"�HK[sX&O��]��1|������Q�r��u��f Y�[1�}��ç�g/�_�OF��Ή=�O�eV�|��e�8��\m�B.���.}����2C�J��������s\6�W�#����M��2j��!
�%���U��W�����w�������+��>u�pg��yԁ:/�/�uT��^ ���O����g�H4���zŨ�\YÁ��4���.z"y���[.�̘�K��Fߋ{_��Q�{�s��\;�=t#0ù<�؛��s��R2����;�
3��0:nUC?@,�j�nk���X��f;�x�4<h==T.=���c���m\�S�A���+��G5��b �v�@h�/�#X�P�6��L5k����v+�~�S�ǅ�rR0:z�f��#�t����j���N�򴓮0���c��T���i��fKɚ��w�0����pQ�lB�4P��k)捽�>U��[4�t�M�7M��i�[)
��C�-�bq��cS�']N�z��8��	�9�"�}.�=u�9��s1�{�5�73�8�:'m
��������b Ĉ�c}�~~x��?x�C�)>�Mc�(Ȯx(�ܜe1�U�+zfsX�M��ZV:�ҍ%�m^Jv�|e{[� �c��o<,d0�_�F��]�+��c�7 $��]��Qe��3N��f�np�<�@vz=�=�w���,����N�[K�΂T۠_�/d@�}���S�Z��#�&�!�d	�
���U�׀��=�d͢�:�YT2���/8��>��B߀%�t_��F�c�\�9�6NQ|��w����~{�� �\����a��n��dTs�<�p:`S>y��Tl1�N9�a�;\%�+��Z#e�sr:���לl��j��3;�g�Wu�3���g"ĹT@�c=�u�6��k�SbwE�P��=B���!�k������s�{fb��X/�Od@t��5ά:��%I��̼���CCO2Y��(�<FW�#K��R��N����F�U�g�-�H���o�*�/�J�w���Z����jy����H�^�zL2�]"����чy��4>���z�� (�d�S���cF���N9mL��8�8n���]���#b�|'��rӼ�3 ��xx�U
�<n�%�;.�"d�'l׶!�u|[W���X��0�Ň��n���t��1������6�ƞ�\A���R���t� 'PΦ<�*�-�=�9�{W��M�y�M��c���j�����A3��1��H��������b��^��b36I�3�Τ�TW҃{O����	lJ[����1)�hu�uH�]���]�� ��(-���E�_�.\��lӽ��h�y�n�����<z����ξ�q?GS���L�ܥὫ˹�
���]A����}
��ܠ�n����;*=g�Kzv�	uj#�*��]�^��|^t`���YQ�\u��P�4�(��*b�C�*�kik�+2����!R�\k.�U��y��G\�o�}q`h����JV��.�.f+��d���%���Ο�\���W�l޴v���M�f�}30���Vr����r���++�V���+Sd�F��육6�-Ԡ���CҩzR#z��c"��'�k�:�kv#�އ���q��@�5�G��f��1�t�/��wsq��)Q�}f�V���7��*�-z�s�N��N�8UNʕ�pvͼ��MZo,G�=�7�.��9Ren`
�����H���N�r��Eʜ���l�ʻsS����M�\�p��-;���{敞�i��Ĳ}�t�W|��Cr��dρ�|}u��������0mv�e�.��M4���.��ڰ�L���nU�4�>5�J�jղ^�7l�!�eL���@8�<-����V3G#�L&�JI���G�i8�P��bx1��h�V�^!Sus�u��7Jh�ٽ{�me�]�g�p�Z���:.���W0$׽xu����3e��U��QbR��[y���wݘt���Ӗ���n��O�RS�R��g9s3�
�$�v��J��t��	������r�h�Ұ��d�X5��Y}ױ��>PD�@�{l��ͬX�Qk~���RI�W�ސ��5j�4�Ef����SW�]h�y��j,��:����׋�\�.�~^�g�����c�S�j�~.�Y�bh�S�w�Q:�I�dqz�Uq��й���'S6�J�W V��6N������tb�vg*���0��Ҭ�x�n=��j;Y"��\�]���(��	H���N�eJ��VWd�r��̙Noa�Z�t��t�o�5�Mj�:�H�6';�H\�m�/K�ul]��:�ӵh+\	Mm2���oh걓�ߦ��pQ�r
�&�s��vr���������\'^^q�"�Tq���9E�ܣ��-R���Q����Ζ�}CA�����M&�39�)�ݗ+.�MN�118'`����8f�Jsyի�'-��v1�$���ݓ���m[������
���
���a����%⼧���Yf�����L���Xu�+´��:wp:k��9���N��:G�uh��H�v��˧MU�) ] ��Ko��'K����B�!T*1h��"��e1\�j�St�	Z�	��� �	�QT�6A��8�*���$qs��i�]0�����2�t�:�����K�=��ir�$���rrnr#[KV%B�5�t��y�ՠ��+��KZRV�EG�A�U*Q�8�[B�DfOOONNEQ����
�J"���ƨn�{Lʬ�2�N4AQ���"+�YP�Y������Gԣ�]ѽ���*y��Y�X�PF+�Jŝ�(��J�J�������Yg'������;�X-h�&*&+]fLUT��ۙp�[cJ��FV,S�Y�a��JQ�5e�[�������M�uJ���b�Ya��qb1�cZ+l�)��"�6�f"�U�P��m
�����fY�b��_ˤĲ�ϧf��|���)�S5�4(,�T[j�eB��Q�5���.���*X��]2b�]eҶ�Y�������i�~f�ʖ,F�8�)G�L���Z��bL`Q�ִ+sY4 e4aJ�-s+��eL�u�L�����NZ�k[Q�g/�4�X+-�ҡP�%f2�'�v�԰Gv���E(�<�����hڣU�\�uv����Z�5�T��Y��Sӈ��F�)d����
R��L�D�әm-�d�4����\�Q�45�w��qֵ��z0M��Jd��� �V��p��m���vI0��C����Xٙ�M4������*6N����TP7Yr�ַ�f�g1L�]\���"1�X���1`���;�x��7�M��~S��͈~i�'`q���.���>�Ȩ�&�Ǘ��+>�yK�~��{���A�|�N����7f8�i,����:C8��k��Ȁ��u5��B�$0v+�D�t���:Љ^�>y��o�����L{�z�o.�fS��ظ�殁����=��5x{����[����AB���}Lg�;@����nBاf\��)�>�ߜ�K���8��N�����E��B��Û�BS��έ�T���e�#��T����"��hl�w"��7�2z3����z�^mp"Vy�5Ɂ�#&���>j���m��#+�$$3�?E]�+-z�XR�r�E[�[%����{,uY.&T��Qq�']B=�fwBu{�B���K6�[O���KoT��n�Ⱥ�8�O�
a�ڨ�8'0*F�e��v`ɛ*��g[0*-w1f�n��ڇ(�U�C(GE\<�
��j0QX���fEn�x�0�*�nG�3��V����d@�m�acP�};�w�f�>��gdg5�ف�����/S���x�S�*�������b�9�����e��� ���*k.��?<����F�uԤ$|�����U�UV�u��X���P�Xɽ	�C���	}����+n�}���Z�[�Ҟ�F��ػ�� �ޭ�l)�=������21�Q�F1�C�)�T�E��!�ֲ�RP|cս�'�ԧH������t�	����s[���.!zt��/�C�!��㎎;2`��ͺ%��K��đ����^;��ٌ)Q�6�7���Ue�j�|��N�k�<��K{�g4;bg.T���=��Dr������L���!���sm�y��P0�di�גɻ|�� ��8N���>p�kdTd`:{5UBJT�	�C�+��f�9����!�'��s�/`���q�C�@��� �j!��4��4)]E�4�
M+Q�;�7 ������b�Tѐ�PY��kmf�X+�?j�ݹP�8���;���ל�6��;Dx�������9��`�S��nM�>�B;��� Ȇ�,�n���������"�:W^s�cK���<�˜<0��l#b��oǝ�xH�R���k^]�_F6N��&V�2��0}t�v%{
c(|���L����V����No�"�7�#��]��<������=��;���6>M�E��v��xn0�f�51���M��M@��*g���6a��f��*gА-9��r{\��fE�6B��=/^]$��KvWqQ�ؤ�v٥��T��}�����Nu:��p �r�M˶��aD��NǍ�qv��F��*�f���̰�WΔ��]!^�.k��<�0�St͖'�������H��[J;c�5Σ��^f�Q��I^X�ˆ��bV�3U12hמ�|��t�#�6G����lZ5�f��Z��H�~*��I��&����߂{��OX~�O�^���'�����M�j|dͲ��\Wl�u�>��<�|�T�;�˪���Q���<��3�*�'Z+y��Z�kRW������㋏V���c�3��Ӽ��Sa�ϧg�B���6z�ZQ��_4�a�Lr��pY������ƏS9P%F�Vjh��u5'}8�3%��M���sZwC���d����u���@-��p�[M#���3T��LA���#��2/�uA8^�ȅ��N^͵�w�(oC����aC�.޽KVzݖ�6.��'ӷ���4&G7u�+ES�]��g{WzU����0O����m��/��V�F��9��ze}a~S�q��Ư=쥓��U@�ʀ't�l[�6Cl�~c��u�U+�Θm���=fC�}z��xs��}}����{�d\$��P���Z<�s�e��)�N���fl��C`s�][�38��'���Wb�eX�6
U�?DNp���6�F-�C]�ŽAo;4��=O����W��{w*�-�\fZ��wly]Et@e��,�6�ۻx�٫��o+3��^��{���%+���.M�(��|�~�4�L2�z��do{8��i�,�6���F�e��4���6���s7"ѫEGl5/����r�����S�HCsv�|:�T��$i�+��Ur�0:
}�R��uqp".�C��3������vǙ���9�YZ.�7��4թ3���l���CKevj{��c��6��Y�v�ow�9�p��oJ�o[
�ڪ.}ʢ-e�j��՗��9�Fj����|ӡ�ko�,
c��ڍeP7R����9�N�SR�ɨ�����؜3�-SO�٦�D*�]�u�V��߇��k̦g�O	�,���u{�w�@��X�J��k�5���3�8-p/D�J���O�����3 �Ճ[um�ɭ��]9/Ҟ��f�y�cpοS�wMT)k��ZE<����+Zgn_r��.;��.����.<P�����w����yf�/bњҒ����v�_�[�#�dN�'��e���&��`[�;ٽ:�#��/�vOj�t*v^�p��X�÷�@Ia7 [i)�غKީ��wZY�\�zEo0�w�o.�I���_j�A�>�_�N�ge�<ץ?&u٣˭���������٢J ��T�T#����<	�>h9����A:Ma黠9�mv<�Jyn�W��+3z,P4����k��xgʠ�9*_;u�'��2c����evk(�����1q��/;p�,s0fN�U���8��[H�[�n�s+���=ߚ��3<�k�r_���a��iv�-<9��7�8`�g@]��\;�r�X���4����s�g��*�iڤ�Z���v�&�m��Qo]���^�F�}����"�6�sV��oFǎ�e��m|�c���깞�=ͦ+��wK���]��y��'�F/��5��籊�%'c4�3���~�Q�S5]�gl�]d�Ū��⸿��5�H\w(�\�'��,�\^V���xK@�[!���j\��Z`���x��9*�-�'�ή7�6{iNU\3g t�{҆�X��O�-$�(�c��>�eP7o;b����u©g@�Z¢��Q'��ދ��������Զ��YA�O�I9ԍ�NV��zp�>�e�	ũ�*0k�%|���a�:��csM�b���n�c�{�oZ�o�]�L����\��xds��`׽ӯ�=7�- ��1D@ǭ��33#gsL� ��/��h׆z�>�[WC�ym�*�=�VMPm��.
�=X��j���É�hOճ����;���rౄVyD�{T�Ǧ�=05��Wo�ؗ�m�F9�\�:�T��Kl�_V�������*���s�/@�x=%����4þ�����Zѷ�$=�3=��k+������]'����Z�2[j��ұC�|����&9�����d�B��h�V*�rT�X,�Kh�j�3o"\T]�.1"	�ry�1�ܶDjط�Y�}�כ�fV�b�<���I�fY�U}��٬H$����o�3M��N�����}����ѝt�}t�s����:��:|f/%�T�_x�0�o6��UǪ�f���&������M�`�w*�P�M��#�8�G�c W?�WDP�yS��i�u؋�づ!C���ru�>]@93푛@�O@= �1n��+�]KB�U���_�[k��t/ɡ~ܖ�����P����^�^����TG�ŝ,$��|�ȿ�N��S7��8^Tf��93�Mqu�@��x�P�Kg8>fj�O����bP��8e0)v��+�|r>�C�lW/�ESj�܆k��	�> ���j愅f���]�*����f����ҨG<�f�u�f�	k��W�g��<�+�Q5ŭ�7J<����G����;�xAԆG��������;�rT�]+S�s��oK(�ܳd���R+U���j�t�+�6aG��_MNȻ����W�
�[��U�Lf�����?_}y՗�txBLsk�<m��|�l ��p۱���cz�O����L�!`�3i�uOKEf۹켘�[]۷�ӷ[8أv�J�V�L�	�C��EYQ4 ~��l.���3����f�;������,R�=�y=��j���x��ͧ]��<���Ҧ���L\`یUn��J ��aZ�w���'���q��k��3��v��� �F<�BͱY����ТA��9�#ݹ:R�5�Y;�ޱBL���`���5�(	N�Zu07%�=���8�����<pF��a�pj��h�P����
]�C0$���T�y�WK��2kf���U��[�^��(�emv�G���ϟl�]��u�q�Z"�3%u|�e�	�I[��c��?s�m�$�n^�Kᶚ�_rF��<A�rۼO�eE�k�w?wn�_͊�3��;���pݽ��k�&�A@������2$�7�[Vݞ�R��>��d���Hk�9�Af�$��j"{pWN�cᘉ"f���P��;����K}��5=��І��e��x�DU��|�x�(�G�u� *��������tb�:<�5�1������=�����7p�����������H��Tޟe�\���SkFHe��_unV�U�_����<G�i���??QYW��'�Es�`e��oi��vk��M���}�ո:7L�J����h����L�P*C�Z�\��FN��֭K��	�o!{��֤��L�溚X�J��wv��W�����k��ʈ{���b����'� �s��ZU�,��qN��N�k=�={Q�Y�co%�&+qK6 �eM��c]��9!*��uS�!1V��3���,����%�M��+��͉�7��^�_:K|����:pFh#��l��	��}9wR��J�"�
��;Ɏ�^\�{�C7�C�]��/����wK�Yg�OD'4u�\��g_],�Mo쳌?O��w�w��<�>KS�5���>> |@>>#��ֽb�ebk��)׿W��^��nFt,�+p^.x�[r[�8;[�߻d�n��|觝���]#;��{}Gc���{*��szf�yg�U��>½��!��!�:�j�x>J��w'�z�Cl־�{���Ұ ?��:�vd��릾Ř6�[��^|FX �oa����m�IU�|.��lU�;-3����"udeƌg���lQXݯc<��[��V+3u����3A9�a�}�"Y4��ǚ�hxƛ�Z.�W���Ʒ��@�j�Һ�gnyY� ތ���\aV�W#���ߚ�x�c͘�S�}�iRڑ_��o�}rG�����c�������<ϣ�Zo0Sq���-c�o\�S-��aަ6M`��h�M�����������Fs��*�f��p���%8�]O/$��~m�lЖD�a�6;�^�z���3�������;�]��nܪ�J~��g�8Uf�zs��r�.i�nj���!��7KS�"����D.���e�ٔ_^dX3��~�'p�*UN��(�%I��#@P�Y�Mٺp��ۇ����7�j� �8�\/;�C�-{��L:d@���6��E%������~��"����A���������s��4: ��W���q���)r{d�G|n�x9��*j�}�����U��F+��q!�����h.I�`ղ�Cz#�pn��h��ΆM����$R���o�L�Uޟ^pMi7�w�)�cν��373ӽ��i��Qg�)�f\�b`.O/�w�h�2Wl΂�3�{���Z6�*;�]�o���B觚8�5V��u.+�~d�@f��͙U�������w��%c"��g#ڦ�=4zEM��d���ܹ��>Jp'H�f��Բ��Qq}�,�Wx7�G�૫%�}Oo&cŅZ��4���V��vo��O'����\^�(���)����Y�/+i��� �j����0�:�p �!�f�X���U٭��h�~�m�ˌ[�Y]�Cd���E^�ݡT��<.�M@��}.�JZ��K�5s`�]�m����iy�Wޒ�� XF�/�e��t՚ި,�f�b|n�Q
s-�Qe���=q�xt&�ꭠ�ߘ�@�Ä��N.�l�bPP�O��uv��`pVA�X�l�bd��h��}Z���e���<pt��y�o�%e)*�U�l���jHrA�J�x���������V��N�3�tz� �\[��S7e8y�jd��g]�eq\��������CY�<v�G|�Q�R�R�lS*-��$o�4��GLb�\U#�k9�E-r����Z�k&��1Zsu��>/6a�ɬs�C0���j�Y�����.]��!��%U�Z[|4x�fԺa��:6y���*��p"wfZ���:�J\(4��EF���/nm���Ɵ_f[+V4L=�WFqQ��I|�p�O:���՝}�,I*����J���۾�G�a�R�딢���Θh�z���B�,�P��7�]�]W��q�Y� WZ�X�x`�\��DE�^��f�R����c���B�<�\h��z���w-U1��e�%��khY�X���Ӧ�z��\�6�np�A�ЄK���wX���-�}��K*ҥj�5�Atn�l��:��5t޺���-��W9z6�+��*[|���<�&�jOvQ�au�70dƱyk�.��.OE��We^ϰk4����F���g{6W
	ʃ���/q/
�԰{k.,�C0Ec96t�C����K)�l�3�o�(���g:�X#�Y��m�u�[7K�98%:Վ���`���}�WZR,����aD�
8B�wڐ��}��G��l�e�ݼ�i���[Ҟ5T.n	Ԅ�)� R��a9�r�L�l��R�Lqm1�\/$k�kJ�h�8�=*�޳<H��h��:Xp��V3�R�*q�����C�X��S<���iAӨ�<�q�7�����+9�S�v����N<X��X{yb
��n���H�;���˺���w�iod����WeS��@�m`>I����B�!D]>v�4��V�lb̼�ǜ��)�Eɲ\HS�&G%\Y�o�c;������|okc�g>�W��[�6��I���Bl��������0뭈;٢���:�w9t]�R���o��鰒�yQT.���5h��Z*��1_��%u9wcg"�{J���:yɋ�c��n6��74.���e$�mТ���ef��=��%Kv���Lb��������5�EN�`�θ;C��j��t�o���%�T/r­��Y��`�X�9Y��->�sK�4.�VD�V앃r�����6�n���sa|���	�]��Εr����ml|���x��������'/�b���ˏ^�IΚL�z�U���U�[��>�w�l����{�ݝ��wU�M���,��DPϮFa���MkB���V+��jRԬKJ��ٓs��nr$wE,��Vً�qB��)Q�@Qr�J�Cm���b�Mҋ��jDLk8���N�M�F��
Ņb¬UE���B�H�uz�;�`*���Q��IYS��h3�r�OONN(��%TO�b��A@Tb�%�P��R(*��U��+�Y����rp8�2�Y22�:���Ö��)Ɩ�m�Ȣ$�q�����*[QD�[i��&���&�'-Ph���Q�\ʪ �m*DRߘ���-�*-KY��L�-��������q�(��b�Q���-�J��3(��f�pb�KB�A�>�O��&��*��QdD8�3-�m�/3+T�b�Q�G�2�Z�1IR*��*ƥ�N�OM�D�̣��2:j�iQF*[�bs.+-ZbT)�,k,-��y����DbȢ���
��Z1T^s6ɥV(��b��R����\�b���:�V�׻w�7�8�qyJ�^ooLQ�r4Ku�J��O'8��S|�I�!t�{��t􇢶�5��S^���b�1#c O���c���[<�l�������Gyj�/����mޘf�Ǯ��04a��y���:��|� V�m�z7U7H�����xώ*a��\'\ęv�f%,�x�}Aɤ��n�U{����s���98�@a�\Y)t��x��ݷ{�1�qZ�V�_�5��x־m�����c]/�UA�«w��ٞ�� ��,
�b7��ؠ�\yuRHz��_i�T�Пo��z�[���կE�T�y�J��릫Z������!�t,j�ݺg���\�ϥ�nKr�A�ZϤ7A�T<���U����t��h:�
�C�n����kq
�*.F+/v��}},�j�:�TL'�������!�n�vh�1+�;cx{i�W:�bSQJY�b�3�Ƅ�G����a�7���F�g�
�1�y`�K��-��E`�5^��V��L�	��!��s�=�M���/��)P�.�����Ҹnh��7K�ӂ�e�xym^���5�WX��1i��ԪK兓�� �.�B��]����jQj��v�Z��U�L�]�n8d`o�GdB�����=;p/���x�x�EuWc�Q_ODC|�_��vO�3�y*u9��+��ʴ͵L���:{>�����Z��M���hW8��K�ĶA�Ѯ�s[r�ʢv�3M�fڢ�r�FF��^�;O8*�>�q-�v+6<��q��׷1D)���;��w'���U��c����B���wY���=Zr�/�i�gs��拙�]p����V�T\
�o0c���:��=���;Y}&_�4F��؁����e<�^�G���n�dd3
�w4��%c�n�9�5�έe�9�C5_vΉ�7b�`6�Q��o	�\�h��k��_��-�B�*��:��U�J�l��5ٽZ`�jz��uےgl�>���S�aG�[K�Ặ��w�{5���n?��2�AS�9�=�=Vm�4�}]k���s��ݔc�P�o�Z��8g`<3ժ<.c_6��7�2#	�ݩR�՝ob�+�oW�8��Z�CB�tw�Xl$k�{ە�:��֩�Η��g���w
���JJ�5TSSE[z�.�I�Hs��x������	n�8�DS"�v��r{\5�u�����3f���;{]�oZ��a��bяm_m�+����-H�"(#J����������'�#�j&�u�̰>��`�g�����0/wFO��@J��ܥ�E"՞3�թ���nϘ*�ݜ��g��k)	�9�!W��6�K-T��t�>�jdC?KQ�}-/;fߚTԈ�y��Jbi鮅�ʢ�R��pkf�2x�\k�
�k�Y���ox�?�K�p"��`�W#���֢�j#7�v;9��V3�Z�����F׳��7"�x4*ظ�7dt�o�q�ݐ{��Ͱ^�'}[�sꅐ7���&5�x,V����	���{U������ �ۈsB̡��ة�7>}��Ί��d{��;w����T궢��7!�=���mnB|#h�%Ps %�x໋�Si��es������d��0�,��n��z�hc��A��}�r�ަ��+3{d�5���I����L��-�V8�(~J�.����o��Q�GoO�H�ʊ:�Ǝ�*V (���e_Į��Z)f��$R�Tm��)�Po���t�p�Y��(Gx��Xv��;֩t�c^n��S��R��L��=1wY��<�Z�W]��o]��>ɩ\A��6|>�P�������m�V��}hrɊ���w�� ��8ĵj�>�_w����*�h��웄�y�g*�݊���c3L�O�ͽƙ��s�>"@�Zp��̓`Ǎ��
��ڻq6�!&��>�w��\1�4EEV��n�O�{]��z�ր���}a��������(�u���f�v���{�����&����4��
�U2�s�����x�3�7�v�4���ǌ�6.! �y�pm�5dof��{� x��%?��M�R��!�>�gw'5�#rwr�ļy�vlP�q!]����b��Iukn�Ӿ��vE��2�����6X!�	s���� CR��w�JW"�+�<�D���=4e����4�}]��3��ښFV�w��t<�P%�Ű
U�s��*�"�3��Wu%��#�^H��euf��A�ٳ}8��i2xDk��m�%\&oz�_�z�7����%brmTMSO��狶\n�x�0\>%T�&���F���Ǡ^4��qݍa�֩kYT*KJ�ARܨ�;�CK
��ڱo�N|3%���rU;>��V�7�s���7�s�̫���oI��mbm�s��3�@)r쬵�'I8{�[��2�v]r�.|Ս��_|� xR��|h}��=��3���I'�,}��t|ٕ����n�z���x�WG�+������p�[���a��Oq{ԣ۳Ѽ9�c�̅�KgaT,x�Z��,N鸻d� �^PGc��اO+�{�����r��ɥ�S��q��M�C��Ň�2^�xL���;z�	K_oE.�L�����$���ғ�%�fy��ub�4�'^;7�]˷д��}�^;Xc�Q9�y߼�"j�T-f������:�P�i���'����T�υqf�h�"��x2�.Ba5�ژ�
z�N��p�Uy�G���{��s�� ��Go�o�BwA�Ǫ��˦.o�g݋�y�� �z�P�qJ���|9z�پ�ou�P��H4�J���sN�� �eݲ�c��%X�l���{,��ϝ� �_��C�ׅ�e�4D���ע�/-�^
��c�vc�������ϝ5��-��{�9��Ra 3��Y��.a���டwZ��r�:h7�]�</�]�3,Up[}Քs'JԶ+绮S�� ��-.=�%�H-�|۹�&��/�ټE`x��3y�-���46u�p��̍�\�&GS�MZ�]ׇ����ގ��3��=��$��z�$h��j��ƞ�X�l��2�{p�Æ�ͺ�&{���c3�;	���d֊y�,������h������5P�j�j�JYX����~/V�/�l���ZX�����$��8�1�9�OB�ޥ��T]�f/@�2�f�8+d���}}���j���e��h�P+{Y*���B��ґʭ��g��L�N��1�s;�{T����/o��(p-vG�R�3�S�;T���Bs��s�4��x�H����B�q5n�9W�gl\�3�Q�	�.:�ni�ۼ�����%:˛n��:
�ј
 ;�������g45�ˌ�y}�il��|���{i��;�����l������|���WS�Ƌh��y��y��RD03��~Lʋ�j6��|�v����5�-��[���<z/^`�`�{q*�m[ �O#:��������Ɉ_�Y����j�6�E�iv:�n��M�ƃ�o�u���oޥ�o�h7Jt��z�V]'>�b�L�Yy���N�m<�t��MJ4�>��n��ϟ>�&Ǝ�ۀO�ʐ��� );	�Z����Ъ�7����F�Nv�ko���7��'&�( �#1ՇB����^��=�h��=�!;=�,�}�y|�~�SV�z��*N�=�0�[�5�r���q$��#�^��@��B�
����hp���/���wx���z�����*e�wg�j��;Z�}��6E�q^ew�[�z1�{�y��uzc{T���.ƽ�۟P�w3����\n� yvO�����<ÚYt�Cb�|�>.�y�M`�9�w9���f�l���
E��r^9���G��.5G�aWQ)�HUL���-��&+r�br�/L�ͷ|����>�z�RTj�g�5�M��ے]tI�W�:���D��K�( 
"v�IE	�7��_)z���>9O�x&w�gv�M�1n�{ ��IƏ:�~��Vk�)�����������
��\�߸�J�A*���i��v{:j�q:B�����b�g�Ā6�������b��^��q�\��Y�i��͓4�bj�+ա{����~�s�[رD�W���f������𭁊[�U �v�f�qF�&�^�ٛ|j��z����Y�:��o�EA�y�r�m�E۷s��C�z���c��)'��4֮�]��V�v�57-(�����ɼ4��d�8�<�n�`����Au;��!S�?W6�����2�w�'f��m�elt�R��灙s�;�z�$B^���\N�̅�69-��p����'0���)��R���Փ���v�>O'�^�sǺ�d����l�`P��B�k�J��=��:o�x�D�7��#�ۻ���5jg�7U��-���D-��j��ؘ�4VF<�uq��F���.����}p���3�\ns݉z����7�����llp��7���>�e;`���B��:�̭���h2��A��lnl6�X�v7OH�̷\��z�cE����&�D5j���ۑm!W6�d&�bvFk��?���q�����:������t�#ߓ���w���z��{<R�-�����q��� ��ÉR����%M��ˣӳ[�7�R7�3���Ws<��V����bB�n����l-�")DٳO�j���~�l�b���[��o�ؙO�M<Ix�=Hf�<3޾��[�� �n��w�W5^s�A�.��CB�P�}�/�z�Ŝ�����3�w(��a�<�\�n�"�q����˫kcA#��Oγ^��-寵�����p� Q@	�$��W'�V�S��t����^g��pR���"�x��� �w�P*߂|�w}�*kҹ^��
����s�M8�eto�EU el}����#��vڲng�ޟ�Z'_�R[�/�l+�J&7���Y[�ZY
��Y���B�{�1�UƉ}9��g�z��<��ܒU�5�uz���,qĿmol_I0�[�>L>T7u�>�'7�]�H��h܏V���av9����l��a,u=W=V��-bS�2�Wy��apB���;�T�GR��=�Gad�Y�2-�\BLL��h���I���e �;_��^l�z::���kF�
���5�E&캵������^s�8dgׄ0W�턮�����V�)��p�-�l=ַ�<Gp�W��p��G�b=�F��B�!�gT�)�؎���y���9��^w,K�!//{��ݒ�}��:�h�+���9WN ���T��}�nVp:��v#xڝ����/����v-�,�nYЮk�v3�q|0>F�\TN��}��z%�o>��f���)ˮ5#�ݳ[J-��k��ɵ{+4�W���FX�ʵO:���m�p���Q`(��d��>��w��������<~mOQ������,�����\�v�9�:�>9i�n0�UC�n�\7��Ҍ�k�1��ld����3U9e:����J�����3I��,{X�źgC]�_4��I7o⽏�-y�)��	�sE��lwk=�0����f���j��	� L�	y����6ZS.Et�j��1�y����p�k�
���K(�A��{p���M{Q�F�Ms�as�Ⱥ<��Mp�w�Y���>גn�Qy��E�f\�ۣv���L�>K�8��������+>�O$V�S^�C`M�,��VBJ�VO��Ŀ��Ș�6Pf���˙}Ơ�Pnʀ��_a޽�K+9L�:����S�&֎�2.V^ s.o���[��"��|�eϴ,-vA�ԫ�J��t.�_4<����ݖ&2.'.:�x�j�/@�{`�Fp�����Ӊo���\<��W�vN���|)�������Wx��pi�^�;Y��c��d����p׻3�7�yO; J�-e���p�71�2�GfЗ�2��O�<W�B&�"�A��\�_wc���|\Sb���]�X���}xS']�����[|���8�z��ic���M�|��q��޴�}�b;��Yȓ[��x����I'�u��ި7*'��]on����'n����b�_����6�Nk�JL����/Mdف"��Z+c2a�^`溹�b�I
�v7v�ki���+;fWZ
�Q)�j��Ty�\�zc+9�n1�������w��h��� rf�IM�Lv�uef�떩὾���(I#PU��A��r��T�[��&����lVˎ�S�u��wh=�37C=ժ�  �pc]���h(,n�}HqZ�+�{�b�1��<p:�x)D�k�/6J�]�od:[`��:�:W�`�R� �uM�U�)J)��河�s�U"*�7����h��}\�5��K���y9����y8��ڴw%N�vf"��8#h�|�3�ȳXDJ{`d��:ý������x�������#+�������f�#�m�
���ٵ����Q��
.%�R�`�k�+��G��,[k��r�NJ�^��՛ݵi+{)ȴ���^�.��Qkփ�r�އ���t�Gv��\Sq�H:��e2�^�yBsZޔ-h����я���G1])�4�8��n��Ӕ򳒧CK���x��v�x:y�yG+�079t�QwWr��Қ�g��:�D�m�(�M�!X�
�)i!����[��X�1�Ƿ3'93�	v�&
�Ćf�	��Y�rf�`��9ٱ����5ݜ&�����v)�y�wc{x|��+��bK��٫��e�͹h��a�S=��,��J坳i�����)�e$�oM���6�oX�Or�$����ט7�̔V)F�t��df���3vi`)����*���5��a�����9��!�Fpj�y�+6���)���A3V�H��u��	S�e��y{�Z��9��h\�Ŵ��m���Z��<푓w���՗K}���f�0<.�fh+���Y��fj���:-R|r�.9�'C�����f�o4�"��U^ ��{�KX��L�Z�OE6�k���Q�V;hV퍎�U����8��WX�ʈ7(V���\���C57�:�n�=���du�W&qA\(�E�s:�gJ�����K[H��|��m�Gq���:�=�]��H�z���U����9V�w\��V),�]7�Vw���,�	{��V����dEC�<����*���k���!\+m;����Ju���4��ÙW�,�;�{+.�p	n�l�G;P�h:��b]��3��;�ռ�޹ʵgu3x���b���ks���a.>�ݮ.�wY���j�ax�r5@ҦYKȀ�v��Ukh�J���L����*t���ɤi����
]
�)&@T����L�Nk13��DTụ�u��M%��#���ՅƬ<[��1��X�T�*��b&L������a���~������
�4�(�J7�^3L����F$bD��
*j��R&[��������.�9>�W�
�1* �B�Enae�kN6�(��.(�%K��������\ʊ|��2�)F�k,��(��,QW����Sv��k?Sb�3&����s����S���kɁ��n�ff��g�b�Q�Q�*����Ne*��ƍj��#�fX�M�O�'W0�
�lnY��]	���X�"��-J(i���J�Nav�ZU���[�g���g&���^٬�TcZ�UQ+Ƌ�EF5�.R�Mf��[[J�h�h�&���>^��o��Ub�	QB�*Qj�a��m�߉�e���iZ���ӗ3M-�t�(⥊�V*�ы6�囟NN�R�ܔnaADDO���TuB�V�]�~�5&Ϩ
�Q�
�>���WQ�J�WYjek�h�@ˋ�>�U�G�J(��QR��+��M[�S)��!�(�¬T��V���NG�a�������׏sڥ�֞(<��ԆC�� ʚ#�٫��P�!{@-��H�s�]�ೈ�d�5���umhUsv!�S��3�݉�SWj�iӻ�k��# �*���C;��D16�'���on��J�]sv�F���Y!��7�)���<T�c
aP��nlep�Ľ�7�3H	j�׽-��iEnW^� ����x�f\Ĝ�5���U�Aʉ���֑s��RN�n�M�Z�I���� oFV��ô����S������x�ڬDc��ٜJ�j�G������0X4�����WYz"��Y����q�Wt>�S�k�/.��s8;M�m��f�ل55il��cm��
d6��_�n�^�]�ΏUu+�k��q��z%����n{�]V[<#DFg��dlx��s}alQ`�u�W&/==�1Fh���G6����v�b����Gq������ӌ�CZ��.kYåT�6�S���;�ݡ���j���˳W��Cot���1���-;=�ji���m�����1�E�t�w2��+���U���]d��,���Cr�T��'"�k^Kkb�QL�m���ye�{e;<����೽���	��r�<�VO�%�C9`?�wj0�_]@�4y��RIh%�%�Ů�6���v��ooq�H8��4�!v�^�
lj��m�Z�xH�k��ז��>>��ջIDa�7�9�eD�,�'��ԻǛ�x9Tu�?d���Qn]���������yX��O�C��==��/<K�D���2���٦W��W�p\�w�+��\��q[���!��(�����w�f'�$�)�z�)����j.#t���v��_h�=�+$j�~̋�ʠ3{����_l�1��x8[������Iv�;8'ұ�U�
vnn6�Hͦv���g�F�ul)�/�!�0�O;��Z�n�ޠw���O۲S��hk�&��j�9�x�@���%jR�;_�H��S��Q[�R�-�Ӌa�K��Փw]��4�l�$�>`�6�*�L�$��f���k���
b�M�)����q�B��l�Ƿ׆����.m����Ӭ��τxq����D����T��aͬ�^ކ���_ppqp,"�M�+/C$�u�n;�;��>*�V��k^*�I�E+X�v���	���-�(&ɋ�tr��|��{W'��u��o���]܉��
��h�kT��xc�9�е����3�@��&�n�ṽrTVw��61�\�XB�Z�u:��ٮ�nu����煷I@��wamHgM}hõ��q��y���= �/�\�-X���ȰCpH����M�6ktR��R��qZ�'_ө�:�=7�g��g�F��U6Js�^��<'�H���w*D{�����i�ܣW�S��?z���+ߋ��-o�w��f��D�ڱ��>9�i*x��������1!u�{�q �=��º)�N���b�l�� }�ڐ�n)�����"1�J�GJ��km�Ӷe;�^�6��������ҙYE�lq���K����m��wl٩�WZ/D��oN>ޮ��WB�*Yx�LP�M�t�\�4�h�(<%�3r4e�?#���D�f�m2o*���I���k*^�����;u��#��:�L��m���Pݙ��Q{]�>��t,�ޟ,�}z2%�M��N�Y��u�<5�_�a��t�$>���I��]�{�<ze�������t+0c�a����S�d|�]�ϯp�$�����u�'
Q@��4�K�`u	4Eh뭈Z�_pcXˑ�I�����S��Z���R��/&D�ܽ�6�*�	�x&w�=pPw��q��"�Iz;84<���?|��$x�*�v�*�UEF���>�s���-�2�K6EROu˙���iޜ��fn�C�ƂN$��Pe�}js��e�*��;7-���ոI�v�����2�Y�Y��	�3���m����t�a�����u������n��&�u��y�;�����W!-j�M!3������9�f��v��4�l��o0�E��Lsz��*yk�]��Y��7��܇��N�DN����퍟&�A�0�vbmKE��]���U�5��^���W](�v�=�������5�Y{�H'����x5ۃ�!gG��@z��m�я�:_�w4�Q���ݸЄn�^�7v���S�6����utä�])��h�w��[J���Dpp��[wY�����Nc���A�-s�Ρ�*j�vk/2��M��<����d��*/v��ķD���#P�����Bh���f�I�f�qA9ܾ�Ei��/;�q:+epҴ@FǗV�@�ӤZVW;�/��B���(��*�?P���(Ɇ��EٙF�)����vp�u�'N
��峝Z!U۶*;��w%|��%#����MZf�)j�Vfw2M�	��
�D�b3A��$�	#�&����%\�D]��\<|B����p�Le��̫w�b
n R�i�4�	��ڇ��uOew<��M o&��}^l!��],���~z�.v�ϼy'nzuLZ2}����U�3�/�w�X�+_ֻ }I�ի�U6��3Vl�7W�W�\6��n�U���*��"�\��'cNO�C43�)K�m��n�\������v{���J�|���:u& ��ђ��L^Ыg�Mw�-���Egs4w-R�/���*�0�!���q�;c�*����\�V�Į�釧���]���`���}�u]'o*/X����b��Ϩ��m��7,p5Ϯ{��Dc�k�>�J}t�2�O���~aP9ug" m��G�WY�O�}aGD�A ��`�v}z�d�JE�.����F����;���Ϲ̦��BF���4���u�h�_��{�"���:S7�0�url��e�kZWS�ɾ�����Q :�o������o�]�sq�X�r��+��vhƋ��],�޽�l�k,oj�mY\�C��]���s/�'}iv�T�4�;cF�p���'`�{%Hv.��=��b̾cM�
c�ZW���	���ɦ�/9k���7��ߧd�x�ߏ�X��)��}\���ފ���վλ�p2&z��\�\��[5Ƈ(U�,�ڀ�o�Z˴�2��n�庾�m�aE�3�m%�E���W![���:�/�S09�^�P-;-�h����j3�ƴ��1�K <T@�݁����O�h$)����ϛ�F��Z�=�5���*\�7�*jDg8�`�bi��C�m�N8,o��A�|�S�����}9n�Q�����pK���<������M×�YU�z� �nO�͑��%*��r�y�S,�j����+C@�lu��9X�	k\Dc豕�f�v�<��� 7z�@�uJ>Ɍ��O�D���4޾W�8��:��17|Ԑ�}��>p���`mj�г+ܭ���O�o.�6��HB|���)��ɂ87�]�5zj5G�fJ͠o��m̄�٪�Ρ׵4��^l���x�B�H:m�Y� 8e���Oj����V�K�������:�и��۴�\����wP��Wt˹�Cg�����;=1��{'
u�M(��QsW|8���Π��z���l��b˶��Y�5�}�����"�e�T�G[|� ����l[��|y]+/u�(�;��j1}s��]atcu}���VC���)��컵2�]�65����o-�������s�\�Y���`Cdzܱ��.�?b��E���Q�
��~�<���uN�+���y�zc}|�A�9�ͦi���H9���"�4$��)�{����=V�w=Y��0+�r|�= ����z��5ԇ}��u95�A������N��q�}ג5�;�/T>�G�u�0�NV���{Oi5Sw�x����&Ű�-�ې���q�MOY®�q&���;����}�H�{������ӰZ�oH�"�j����&��Ҩx���<��F�c��3"�=!�L\wIk�-H��\��k��ׇȚ����r�� �C��׹�m�w� ޘ����(��>�釖p���C"��[94�������#1W����F���>��ZxZ����ͭ�2�d�]L~�3Z����]�{�:��^2^_V���]/Z��y�C]�S�u��u�r�X�㬣�$Y��pv���Gf>�����z�D�eb�X�o$�����%���Y�e�-�����ǀW�T��U���eB9�4\Rm���Y۶J��wPY7
��T��2jMN��i2��{����Mu��z�Ӽ\Z܃��Ft,����-����i5]�S��w���^�eK�LWd�ж��]$_�ַc�����z�H���c2�'o){;ouo�z3�r0�y����ś�[�+�,pKNu�����-�^f��ٽ�R�䥷tZ����v{ׄ@wK�l�"K�^u�l�+�)M��.��Y����m{�:��뵆9�w6���N�lk�L�z���Y�[����8ͷ�R�����Vg4�<R��}������P]l�%)�׬U���u�v���J���ϻ�ۥ�X��C��l��*�+i] 6U���������J�lam�n�=�Y��ۮߋ��g3��l�'_CQ����[�2#F>��c1��)Y,1�K�M�G�I U8b��4�9e-�������[�QNt!��5dJ$�e��ssw�w)���u���N��j	��Z�Х@�Z�sjoN��n�an���F�A4-�+��=�+/E6�.la��*C;1/�;�h��c]�;���=r�[5M\m)}�T��Z���;�>��{�۠Fi�[��M<��5�9�N�\��qA��DͶ���ד���\j����N<s�ԅ��:P�7��+�-Ւ,;F�Wgz��+����5s�}κ 	��o;�R<�ydyK�}E�t��`)5��3N��K�۪/v��n�Q1�8Q�ʳ�usZ9��Z��<r��u��3�j険�ۙ��SEl����+w�΢�u�y/M~����6i�nt�vZ��eD���ԶE�!T���[��jC*�n�j����U����ݵ�~QN�o�9�S����l
�{Ղ�R:���ڨط�s���[��0N��cv��ȥ;ّ�խ��;g`�{��"��_�k��Q�|1����	{� U�i���,g־SϬ2��J�Fq-��!��N��6=��r%���P�Fj�N�4Rq�.z���o�z�\��z��)Z�ܭp=��#9�����g�e��=¼U'��^�J������ �� �b��G{��퍲:[�FD���s���D9��<�z�*U�,�1>��?W���%�IL$*��j��#2D�=s���~��g�r���;Z���G;DNa^�.��N�7	�7���0$�����{1*�+�r��y�nL�*u��Sٶ�n�ߎ�60i`9s���
��-�x�E��Z�9�<��$������5�����o� �`Uly�t8W�(���}�}�15�t�6ic����7���*�5�wm�?K��̣���/��\)���4�*��r��z�ߴ�{������Urod�x�q�z9��c�61k���m�|"���ɥ�_=�0�����S��Kux��/��=��ar�RR��|���<8-L[NB���Ki�}B���ƱS���L	�_��9�ڐ��Y��,D嬖ح�u�ˀ�*f�5���+� i٩�g<��怜��w�RLK�����Ǆ�n�ݮ/P;��nM8�(T�xS���Ҥ��R�g�_���ݪ��b���H=�_uK�*�����|�VP�X��]���R�4��Wzkt7z*�:��mY�5�r�\�W+K����e�/k��,���ٮ�O�+ j�ԍ�g,��QΦR�<8N��m:��e��7��|�=֫�j��ף.R�^��K�$��4
�P[�e�<�V��W�;�Vl0��^<��ʕ�7B��J�YL<��%.�%[�l�T�泘f���A����'�Zru����*���&�vˈ]b�P˻��VZ�'D&�(v�X��ׯ��A��}]�k�fau4x��IYX�U�z��]����^�{�E�vм�:��������v<��ˎ��cK�/xU�7bu�P�z�vU,��{���hn�5v�9��9���뾮�Q�`n�6����k���#�Nd6����
�r�η֣,r�*h��u�"l�T�@�V*���Q���V嚆�};%��×X�l��]�$�;V��U�d�gw0vF�%�N�\ʕ��Eؗ]�^��3)��:�� /�R&]'trXW���x �z�7[�Xֹ�@M��:jF�=�C�^��%^��K��M����+�D8�K�#Xm�bD3�;Y��Ʀ%F\�eq�A�%����/5 ��.��
�0�o8�`WW��u��p�\�j�I�+�Xu�e�Nɶ��E�ȱJB֮;��y���YJ�
&U�ա[R��
=."�X5���dJ�}�ՍQ���O�a��Q�t��r�P\b��6@��Fu�;�J�orF�0N��b(�OVv�Z)���r�hc<͛ö��6�D�tz�2�_���kR����� .��N��98�-�R([���3X7of-����3Y�*QC�w�����RX��9\m�]�9���f*@e�1�K{��Ub�\锃(,}M��5����0.�x\�u�z��iE2���+y,�����7HL䳰k��r�E�[|@�ę��9�Ӱ���S�leM'{���rEWg�I��4/��x,��v�N
�dK�gY���f��GȾs$��^�N�ʿ�f�3Ktr���|m����Nzl3i}��ǽ|�\�4"|f��N�/^b �Bf��C
#��s@̫5x���e�m���*��:��� �����^�LCc���G�Sv�ZL4muq꼲�h���N
���p[�`bT�]O��3��3+������|k=L�Ռ�K�Q�n�^�.�l�&�*�f�Иql��!s ��X��q���c;�hs6�e�y�k��Wuwn�sV���z+E��r�{CV�Gu�rH��X�G.&������s5��%���bc���$���0ޮ����v6�i��g}�z�	�W%G��T�m��uڱ��E��1>��c�*A��N[Cu�4�C�5���x�H�X�{8�����c�)&�Nrwr�
籹��#����w��7sU�PU��̥Ju���1Q���3��a��r���:�]R�f�Xd����N�/��tst��W�W'����ּ�&����v]\̳0*<lr���E�:�]g3V�ɩ��zrrqR��Ô���D.��1�m�bT�D��p���Mj��s�jV�2n}>��'w��c6���؊�35j���̳v���w������E�����������ҳ�U-3*���U)E�S[V�U-�t�N���y�l�������k���XT*���3)TEQƿZC+�2cZ�ӆ��Ȱ�{�P�����r<,��n�i����-�ֵ��,wM��ұd�Z3�SԖrjrv}9����t�p�4=th�w�QS��GVQ5j�)H(����QE�[2rnvnrN��'�t�V(*��I���4�
:��$+1�!Z��Z�cFT�]�Ć�B�R�)iFӍ�,UJ�Wyۤ�~t0�8��U�-���\;"6uy�T�S�Ϙ癓!U��+�U�w@]�^�NZ�}�c7���F�e>�[�F�k�8_�U��rp����A���>3�x���}�#/g���S�Õ3���~�dO�=��͓�
�g�s󓹗���.��v�W�fo\��Y#U5�fDO�j�I��"s�J����6�jq�BxE ��kqڻ@慻C��ػ}��;�b� f��k)h�6Ͻ�F(�S�hUj^�l�yr��Ǎ(�ՓB��]��tӇ�-M�6x2�vQ�
���<�zDG� :Q��xR�Vf3��s�C��|�p}7tH}C�es����R�[�I,�w�zj�y�,�ur-��-��1��uR��{2s�ok���Ƿ׎��a��O���xF�4���fB9[�c�7sв7z��U>����~�薘��ali~vr�Gu����!�0���K�ף�����7��_���Hm�G2��#5M�c��k�;ftX��=r���(R�ofmd��1���7.���򧜳�w�ծf��|d������6K;����A��=�qݎʞ��c5�`]�Tl��h���D�勛��&ŝN��z	畊`[k�&�7`׫�$u_c�p�<c���|0m3IW]���K?k�>�I$�Nu�.X��;o�s 604�߫���>�wTdU�7$.��5��CT9��W����_N���v�Kg��5��'���*+`(]s�O<����E��f����5=G���g��Cu�Pk�ݽ�hr�.��s��u��E4�.�S��<�V��U=U��d��lz 5T[9�".�^���̵[F��̑y.���{�Z]�]���}x9Ŭ�M��l����5֮�٦K�2��#��.��O�1����Z�E`U5��#V������ӳM/޼3�R���nY\(N�{����j�u��Tr�ZX�j��"�zl�R��V��F�\��Ѽ���[��렽�@8�$�	>�K�+�¦_٘-�8v�ƟwJ�����C>����-i����]�] �i�nkDd����h��S˹u2݁j��ך��B��V����ϗݩ�<�'3��k��a[�X�V�2�i�p����3�u����ur�R>=ں�{�M�"ng2����y�R�;����<�F�s볅���T��r������o;�f$�[]Z�ޚ��:����H�N�}Z�=����s�(��F����c\ �M)i�u����r���
h���=��B����B�^Z��u]���n���1�����e;�U�>��f��i����5�݋���k׬�ɱ.j��{o��s�32�>������-�_��,��UH9y�]�1�XG'�3#�������=����:��qg�`�6WO�~�T��D��N����j���_���k:ԍ��z�9���r����D\�<�d������v��+2��^�Bu�ԇҌoS(�8��3���,&6��n���e�*�L���]s�(e�n�X�����s�3��g�띋d,��| �ŏ��̖5I�ha��kdDG��N�M�MܲG*��b�������{2S�Q����.���޿T��5�k�RtM�� �u�Ү/zC%9Ur��i�h��u3H�2੨�b�(��W�M����e����aI��*�AX%Թ���H�\3U�כoq�d>J�><Fǰ�C����� 御�F��Z���Դ�J�Y��I	�3�t��r�FJ�7�p���`xҥ���;r>�;���#',;�͜ӣ�>�z�T�+1;����nv)roN��to�5�,�%djU�v��$Եd�k�m�mćt��s(�U7� K��L`�pB��#�a(ȝR��}�E��³�w�<ڷ�Ѝ��9n���?sv����P��a�����J;t��s�dR�>ڼ�N�-�ox�N�+�;J��]�Z��;f�:��;�=������ݽO$"I3�m^ɬx���G-�eb�������爮��|��܍�l{�y�m���ּ��J�j�N،�d�R�W�X|�b�3'`x�Տ�_����}��WM����!G6�eBp���O�k$D�"��ݝ��*�{ǵT��N6)���پ�"��k]�8Wɢ�a�mYkӢ�xWO�����Ѯ}���tv�Վn=�2i�x/["��'���:��Ӿ �^)�������o\���<5E?AS��"�Vg3�m3WQ�Qtqȫ"�
�JU������ ��Z�ĩ�y����l��a ;v�;[�4x,|c9bՓ"�RW�r��{���'v��ex*��3�}��	#C�w)D�jN���H��6oc;*>�t��76�#��C�U�:�~N$L7��3������U����d.B�����yٱU��e�r��͑d�����c=D��p���}>�p)!s�	���T���G^����������:w��uK��~�[^��o$��P�Ӊ�0L6��a�}�j���#�G%s���T�q��U�z\xZ�����3�m��/H��Mם�y\}�:�܀�\�'�<	�d��#�Jޣ:A�X�/kvw,�;/_�o]^��t��-�q�t�T���\h�*�횋]l�uv�]p��Pܔ3ӡ�+��]\г9_�<D�O�$��sZյ�s��x�d�:�e���q���Nٌ[��{L��ر%c`l�k���n�5�Uh�l�v$�9��n}���tS��h��F�s��f��yp��:d�_u绛��F6϶�`kʲ|�n] G{���n{Q���9�Z�#�f\s3h�ɏ��K���Y�s�ZGa�k8U;Щ�]p��YO^N��h�R�藣%�I��+�Ԕ<*��(�ƍ 
!NK3���:�P�f�v�� �*�Đ���.����<x_�FoY���t��"ÜP���]S��C/����Um�A}�-��٬�VeH�L'�=���=>��]���{�ŕW�X�/M¶7p�����hds���s9]z������\u�(oClxo�����7D���ıZ���&7�������:�.�/�5ÿCS�ڝ=������\*�5��7��HM��Si��Cz#o�8�"tL�[�dv@;�`������T�5�#;3��2�{�ʦ�c��g��<V����z���m/���Th�)��j0�ƭ:!^�9�(F��j;���F��ZP� tȪZE���Vf�O���ᡳ�򸬷��-��:B�b��s]��D�SA�G�����6�+�����ӥ�}�h&�U~ޘ��a��,����g����]4���Ϻ8X��y�f���>��~<�&�W5iML���Fʂ8ʗ�i*k�j��p�/�/�N6�pa
�6�c�{�n�Y7-]�DE��6��fy����'�z�lVV�AYt�H��y���G��-yYJ���N��n�[ J�YY���l9�PtM]$�f�B��\��X�6�m��5u]��Zj5����c���إҹ�)k��;��W]Kh﨤vg�cs|P�gs�״��L&� �����Ao���}+�K��cgK����M0i�v�dz�N�k�>�k�uP��M�ϱ�co&�٫#��%�i���Ғ��-��үOq�����݇{�w�|�kZ�d��g�e���<��m�g`��\>,�5ILY��c�?g^��=U��v���wR��jk���@^�k�ĵ�F��=F����C�i̘I�Wt���t�,��[˯�}�NX�J���i�s��Ol�`�n|e7c����dgr�KZ�P�Lj����ϲ��c����:��jC�����J�����]5ޮ��|�����jk\f�����M�����V"��1��l���WP��V�kw`���4�D	+�����F���"H8MN��\̯��"��d�Nd��ܴ,���xRT�]�w���䌇d遚�[��l3?��zGr��)�u�K$Ԡhi��coN�X=oE����o>&Ґ�\�-��)(����a���@�f�\���V�h��Ó��tr�pN���o9n�D]�,:|J��n��eI�:��dý.۽��N�P� Z�݌=%�\3�kx;�$��k�}��e�wl*P��ʺ�W4�k���!��e�K��2���&*�1��.Y���>li�98�ߡ(�&z�z������.qV��#�H��Qg�/2
s�t��fW�	zg�^�\n���e^����̫�q��}����n|�#&�.�Y�FUdS3��f\��6uBP������״��;Y��1kc/b�+��i(]*�r�R9U�
���,|�1�d��2K���354L��"b� ��M�SH��~U�Qo�:�:dE ���cDoew�Գ�ޝ��O��9*8j��w�[���ޓ�+6�[��VO����O�{S�z�ҝ�^�v�N���%��Y�2�;o-Z^v�k��9 V;�I�~ʬ�b����ة�'�s����<�_�_�J%d�Vǔ*��D��`{�-y�p݌k���؍��3�V�y��w�k؁���!qUG!���d�YT���B�ajee�{�+�-V�����[F�p��R��R���"D�Υl,�<*T�X�.���q�p�zW@ڊ�a�_]�w\ғ����U�V�na�q;��\�ҭ�ʑ��0��q>3��m�Ckl����K(ָV�@�����1���Q���m��f��7Uˬ���]3]7E�>:��>4�(KRK,-�����o����)�]�(��1�M��(���5�'���4�N+m���־���y��ր��Cc&>����]v-/�6�0w����笷���F����6�O1vF�a�'�b�j\���TE��K�m����ŧ��\��;�
�\ҫ*�jTkڳ�ӿ.f~��ץ�nn9��S走�`Lzg\g\������OK+�����p*/����/%�P7�������<�<�O#9�C2��_TEJ��։����r���Q
��\*�ܿ��j�N����y�m6�m�:�nF�r��:��W���M���2xy��$���y��C8[�z�>Ay��JV�t��-��aQ�K7�[���b�ك������Y]"�x	|�<��ה�TF�õ�WYQw,� ��a����w�U���q�j�����Vp�_mW�VEy�,R�<:ū�ƻ������"�N6�YԶ���N�.��d-���ޗQ+�V>`(1��~���������2�ρ��G�n=7��j�r��WPօ�ʈ�B��f�����׾����U��,��3��o���Ϋ��W�T�d���n�cz�����x[��Voum�9��%�,�v܇[��^���i�l�L�N-綋��6��w{x7s�fn�,�@b
�e|,;��H]DE�{�'��2�tu�늬���ҡfM��p?`x�5g������F��USu|�s�u��+��M�pٯṜ��ݪ�RӐ������쮾���Ńl���;8�,T�9�d�	I,�;ӹQu��#i�16�1<q�������`�q������ָp�ʅm����6�l�7�hM�8�j����ю'^xڦ��9�� a5��u\�Z�U��}�ȩX&*���Oksvi���B2w�� 2��H٭��k�ue�w��U��;@Y���*>��	C� QD��G�BL� ��p���0b�bŐ��! D	'"$�FI!���`�BHA H@(	r B����jkv @�  �&�	%! � " @�� �@�,H  FH n�%  F@ @�@$�@R0�d�@R0�I �@B  f`�@0�I � ��� ��! ��d � 	 0�����@"� E"�a , � � RĀ �X�"B 1d�1 !" ��&#�$F  $`�$�)�$d`$��X�$�� Ā�	H�����I+2a������ �	`'����D7�����	 F B E�B)~!9���E���Q��O���y��g��M����Fm�� y/oS�EE�ŀPV�w�r��z'���C�( ���2�Ѧ	 Np�ޖ/@��ƀO��H��Ȩ�
�"`AH AaH � ��" B
H Dd�����#! P�I!	@��� I P� Y (I �( ID� D # , �@H B �@  �  � #  0I	@@H�#$��@� I@a �$��a�H 2@Y @� 0"��@	 � 2H�$�� 2A �$ �  �A �b@@da��`�) ��n	"Gێ��ATTb �  �P�8�9w�9@_��(���[�rE p����j%�j�R����䦷 PV����mLa U�
 *�Cc��0����!�p���*� �g4����p�!!��T�p�9� P
�
��R��z�@]�B��h��)`����n�#(��m���
 *����`	�v�@���C���9V�gK�1%#UA@Z�`���_R@9 �h�˝Зκ�QT]�FC*�EE����U~\Pޟ��
�2����7@1"� ���9�>�A��y�3FQZ�S�H���N
D��Q*��P
*��n܅6d�lT;gg;\�t�\�H��UQF��G#����s����UT6ñ��Z�_^�zV�e�ٍL뛴t�1��I�0��wm�v��e�ڻw�*2���KY�n��u�f�w5펵UlŽʜ��:6�=��N��	�sT�ۺ�T�V٪���z�-#l���j����;��l�v�[Y�3)v���R	��LY��,���v�֫]�ws'm�fնڵ��\��V�5;rl��w�h�խ�6m�Ejk��[�Ρ;��'Z�x   v�w۵UB��N�M=h:��^�x��u����`��©� ;;wv�F�ɬ�]�JH�Qo{n4+�C�uN��we�׭�5[km������5w����0�]|   p���B�
��=����(P�hP�C}���ĉ;aB�
��}�����kM-^۶�
�cY���X��J4��ٻ�:����6�4�*�ەX5*iln��EV�m���$��WZ�   w.�k!Lk�SB�����6�s�Ud@2��]�m�@��p��M��qs�zj�4��z�l�jڴ�s�ڶ���S��q�SJ�6�Si�����jӻP��|   {>����w`�}qAA���k�UMWlt�ã�����'�uZ)�/Nۂ�^����UR�Fgm�E�R8�At]�o4�����֠���n��� /���
�l�UX�%AT5j��h�i�p���Mrp�5�uJ�u���P*"t��4��G t·�R�`4��nv��^��^��   v��T֊��N:(a��zB��	���P�k�E'R�Q-4�t�)S�ۨJ������wM:���v�v퓙X�B��S�C��   �ƪTT��MU#�վ�x�h�` ��7  uv�P �Ӏ4: ��v� 4��  �� 4 Yy�ûs���ь��m(j�=   t�@�{��� PWg  z�^  e��( r�x  zX  �Vp �wg  ;�p�:v�AXk�n�5���-�|   ��|  ݵ� h� 0�  ۈ�P e�  ;��  �K�  ;m�� Sn�  ���Yf�i�n���n�\��  �� �	�\:  �;�  �\  �{p
<=�  �y�  {�àA��� �F  �O��)P  E=�	))P  5O�̙T���� S�A)J�   �?l�*��2dd �)I4eT� j��_������`���a�H(��T{�yS�w�Gݥ�>���@�__�}�}U�}_}������0co���籃��`��c`0�l`�6��cm�����~��_��������r��ƪT�?Ds�c��sk���Վc���F����<6��{m�$d��z�:�d�u�-��-�Y�36�'tٴۥe`�q�kS57���5�KDf���)�Hlb��e��n�[V�c]^m%nڤ�f��H�4�z\i�3A����J���H���x��a���c-�BTa�N�d�ɕ�wRL4o"����n ��ě�t�F�� ��A���+�!r�4��ّg�d�71۸��Dgj��ӣ�+��%]�X2���f���M�Zr��塷��U*��B�RO^n�a���Ǉb��3#7 �W��!L��Km\�c���%���d2j�Gh]������$��J�ݭ�3tc�:��p��[��a��K7]8@̘%��Ĥ�9w�QJ� �
2j��7��2jy��ߝ�u(5���+4��+�Ә��l�3a7Id��u�(���Ɯ�v��Pț�j�B]hW7Y���l�ێ��k\-뤖5Zq|����y��������������D�Cqc#w��{P=�̫�l^
�ޫd�(�1��93��9'�	�I�vk%x�̍D�3v�5&�*�B���P��ڲ�/����x����	AV^Bͬ�������a51��B��(7�X�8\�7k@6!�Y˭���wJ�= �LM�8�Hc���z��b+x�fn�-`��h����KZ��w���ma�G`��Ո�1 ���!��&��Z�1� "�'Avd�e�Z���YW�&���I4�cr,u���j�66��0;aT���6�V젙ȟ|1��\���-ɯSe&��3-$�Y�u6NL�	�^ޫw@뼡@n=�A%o�d����1=_3z���Ȯ�ƑٶeU���P���-��;Kv�1{q������胻�KT���F)G��[��X�V�	^��7	�%M �1�Ce�w)d%�7�r �]-f���[@�ouk�Wf�Ǡ��J��١�Y��cܩ�^7�
:��Y���	��	KQ���a��e���i�4ǖ�
�4��Xn+�m�ZriǺ��A�p�
��u �\��r�-x�i^�9V�:��*�[u!�"�e?�-�S�f��7�k���ӻC��#�SuM=4ol%pCtU�Pb�mI�1��6-WXȠ��2��v��KlT����Bbx �VҶB��Nc۬c"�u&V؆��,�MǇh�ʶ��zXu_	����hE��{|�U�-:�DM�]��b�*�a�
�P+T���%�q�`1��N<B�d�Gf��< ��l5Dk�[7gSƢ��bm�!>^�my�8$3A���RȆ�O{�Df�[x�f%��*�L�^*˅X5�b�,���>��8N�$��cy��B����Y���փz����2��w#K%�R�L�(d�ɑ�*'��O�����.P���x\��XWJ��B�W���5��j*�:N�
�����ʅ�/M���/11��jĠ�����Q&E�J%������n2ܐ
�l�&�C%�&�mm�̉�2�O
�enLv>	�0�x�lej%^��a4��L=(�l�1;��5�Q����V��)轰���;{D��[PJ�#�M�nɷ+-d
QRWD�l�)a��NDdњ�n�D�]ch����M-�8�C�i��಴K�衳/K.գ`50��/
{�u�`�w�1�]�Z��0_b�i^0"�b7��(��N�w��)���YA@�m�О���mCGXof����j��Sx�!Yj[٩Yy�cm����CtY�y,:Xv�0c�����#���"�[�ǐ��	N2]��ǫ,��wy	f[0*�˧�Ӎ QseeA��6��ws0An'�L	u�B�Lz���A0�ZeJ�/b�T�U�r�ۺ6�v8H!�V�
�5����!����� E�
�<O�c.-�m,�i/�[[I�5-�(V�3��V^w�.�T���JQ/-a���e9�d��8��,Ɂ	++i�k���TB�vdˢtK�P;��ջ���Y�/^�rhj���Uf`�Z�iJ�m�l:0	S�e�go6[?�^:��)�Rwu��u�ǻdߋ�H�G��i}&6M��f"�g��E\:�'�*nJ�T��sV�z��&h�E٦*-4Ԑ�	������J�lX9��s�B$dy����`�/_I�sz��,��.�V��Q�%��YC!R�m[�iF�F��5�H�6^��S�J�";)� 3s�`��+(2�b����{}��� �\������t���kU�H	YB�,Q2�F�u1�$�F�x�(���WD2�з%�i���.��L��)���v/02)'*6�H<�����E��*��fk�a��G�ƉbJ���K��c��9z�GWV�(�.C[yP�x��*�֓�2�i^a-Jx�$�if�Z��tX��SU��!�#/m�w�cZhF`e���T�7l�ND7HL�͕.��r0�Z��6�0B��j�3U�ҕ��a1��r��t<��8�ٷlV�;�f��
��Y`{�i��7vӯ*�
�ղ^��ٔ�UN�(����X�8ïoE�1�bn�&�1D�m��W&�"�Vl�ҷ�cv���qb��ʰ6�lP���7V��m���1�xX�r$ y.�ַS��b��tq�����ݴ���y5��!x�'(˸�\��Ly� &�Ѩ�x�%�[�L�.�g N]���d�_�A�- �������D�a^齷$�z�����)lUև�E�lU�����&�Bd��A�����h���/Jv�0�б%�[�{�a�.��۔��8�ykY	Ǳc�Ľ��.�2v�%zJt��@�c���Cώ[z��L��;�Ә��R�e��Y����hñ&�N�8C��8���j�vD�&�GtXZN�ruʻ��j<�tԘp��Ƌ���c
�����]t-��h�j�H�'ыsG@Ƨ6u�ŋN�z ysT�wl U[��t�f��h,Ӥ�)�X��t9Z��K_1�\#v��v&�ڊ���w,�YW��0��ʔTT4���sBk`Ō����9���^%B|�v�N�y*�^S�����[�����$Z��v�^�OU�2V:��*R�4���,)̈́^�7�rJ�*Ź�H�J����Ba!v��;�x31�a&m�ηa-�iR���шXڿ�yP6��[z��t���ʗI��2��,9m:*6R��j�8�PYK`jl�"�ՠ �k\5��t����eڻ�"֖s%]�L.�.Bš���dIݍ�Z����J�֝@�ӹcK(h-4[�9�^)��`<�a�q�|����4�C�Jc��c2��Qٰn��&�����=�,�#�R]b����,��9Y��z�e�D\�6�ڷ�EA)��yx�T�Ѷ»f^1N\DgȖ�+9�`�t�jA/(cW+C�)�2Pt�n���3Wy	�!^,[�7XWW@�(�!̺NI���-�/.�6��M���/0�MC"��Y1kc[[j���V��^a@#m��r�k *�k[beۤ���m�6��5�V�Ģ�O�a��/�\!E�U�ok	B� b�i(ǰ���ؠ[Z�G^-�tUz+�2�맯MJ�񣊃��N���3L�r�݈ǃ�����b �f ��gٴ�E2T�Q�v6��4D�v�
4�6I�!�⺕�ь=�����̟CG����H�O� ��6�k6�1�0#$�^Dm�	�������N\����( �������l
7y��[�EX!�Ӌċ�Ceś	�m���4j5�]<�̔t�.�ӆN2M>��P��7�zfno�dґy��a��ٍ�4Cܑ�`{<�$��IQ%Q�c�����Jt�"2�e �5n�W�D+�� �M8�aki^։�f�РX��ڸ	؂�b�мwWur�lpx,n��x�u�zi3t�YؚQ�`�6uz�'�n�t��\��	�T$A��v�9���0�ùo.ٳ u�>y�ZMX�[ �+6JP���y3����X�V��b(�E�z�+ͭ��`2�Wd�8�v"�j������&���\cF`{��A-1t�sU&oqGB, �)-�M[���"ɀ�߅�oo0X�SA��Zc (R@n�7�ړk(ɸv��aС��D2��ǿsռ�����cs1��$wl���6<���?`#
|$#�D�4�՘�*ҺY��F���
#/.�P��N�YcF3A]�����B��Q��.+�LMB(�u���E�kp,��P�M�^1z�05nf�JMOQ.^�+�ǫ.�1yJ�7Yb�ט�-i��g(� ����!&~'�7uȠ9Q����m9J��GB6��{�S��-�V6L�L�����d˧H�;;��7������*eZn�11�h��CS[N
���E($wi�#��F*�*�鹠2j8��$�Kxov�A�q%IE�ӀK�1�5�,l%,��k\"�cLѥ*VC*1�]�Y�����R0Q�l �75�ں�3r��b,R�yGU-��4�AɅ��6�iӶ͕J�4�WF�� ����tښP8U�����Gm�*P��q�ri�Z)1`�Y�P�@Ֆ��^��u 1r���ՕO^D�a@en2�&�ȼȁ�	�p �]�Z%�3���ݔ�E���e�� �Sꂤ
�Bδ��YBzj9�3i�kpՏK8�X�p7�dxT7�R�-T�wm$�G����2���LZ�@5�5�XfȬV>ZJB��;�b��6��U���gY��ŻK`;ZJ�LX��'/�c�L���)��%Z����I޵z!��F�XR��!hbYt�ୈ��iL�n��U� �5�9�L��1�F��fVXe���O35jH�$ͧQ?q�׺1��bv�@�ө� N̷�ϲ��͆�b�'V���Lj��ծ̐��:�v�B�|hݧ�*;Z+)�ʽ�+4�M���KQ2x�YP�Li �&�������J�{Y����U�2܄����u�Ķ]б�n<�H�i@on�A1Xyo߅L��{4���X��IV���j�p�9H�gkjkۨo���ӫdh�i���J:u�m^����;�Ap��"X5�kS���e�*5m���Dצ��*�/EmEO/�ǥ	�#Y
�Z�lb2Xo��A*9���G��a�^��&���G%�WO�.m�e!q�� �L�yaLpl����G�MYSF�d.D^�m��ٳl(@��S�f���/��R��ws]������K�v�E�/0�p>��ƞ���q�kvŭ&�#��,�Wv�nZ��J�삨��S����+n�����!똂a���߳1���20Ƥ�Oħۛ[�IzUK�Z�@�b ��+���&��6{J�[j�#�͚�
᱓$�4������p�n�ũ�^:��.�g9�ufc��Aɢ�Y�Ub2��h�����FhA����j�������&��{��d:F��ߘ"a�ޫ[�������1=.�F� ��[��%�̵>ݏ#�0cץ����>1S(����r���z�©k��),eX�����f���!6���<�b+ͩ�=�V �┊Z�Y)��Y����m�ZX�f��� 	�v��hI���f����/wR�3�@
3!��RL��v���
А!�BjVN,���z��i�bW�_]8�}��a�V�@��[/�p�c�Z�&��i�y��k%8)i*�U��A�}1,he@��eI*R6��@V87bɄ�h���Q�&��nd�)�:��9�h������I|�Ԍ�����p�uh]f�-'d�ݗ�-���Up	)����ׅa���N�!*8�VLn��E���݀ʤ� jl���t$ ;�`n��m���%r���Am�c�:A3\��6�n;g�"ˠ�]���kg������\���4ݏNӺ�˄kx�^k�b�he%Fb�_L���|=8�)��!._.D�� �qM�(�:�EE�^����X5��
�m�Du�Z���j�̕�TBi�BK���9�1=e��� �6R�p���-�������u��1��(SVH�z�����փV3m0���p�5�̩S<����n\J\�A�q$.��6����՛�d(��ff*
��r�n�GlY��ı���UZ4��}l<{yB�	Of�CmXd��4Ԋ����+f�����є�1��m���b�
)��Y��f��L ]���2�{�w�xjh�5'��w���*�wD�h�-��B[n<�t��.�=T$�򈽖��kb���Qf*��ۺ���dXm�`OV"#��D~�3���Ņ�z"�P��(�c�Q㠑��$�ITʅ�N�ܳ�j�ɶ����e:G�H�k,,�m�Te�V�v>��"��`£N�;��f���v�Ӏ�F��d`Ez�܂��eDb�8�ܥ�K��y�37s=�һ�v��R��ƃ#�I`��x������m`�
Xd�nVU�RPb�虲Լ�V�D�ⲉq	&�5�:HYp��q'�����m{F�=�͊釰��6seGG�X�G$��2�����f�ɤb�A��8�Nʬ�V��Jh#��+ʱA��n���/J�Hi[�%H5�6I&ۻ��&���Oh�M|S3x���ɵ*�hO(ށ����Q)�P���:v�n=9��Z2"Y��LLLw���Z8�a���3w� ���p�)��Ǹ+��<�ʁ��ѝΧ�-;ݜ�>p�����6�d�Ϛ��{�"�I�r���ɿ"[�ȑr�hN��{M�e�"���n��;Uga�E2y7`���Y[��]�Od$"���m�l��p⽵K���[���מ�o��J5sc��ִ	�Z̠�X��"�Ҍ�\s�n��ֻ˱�B��8m��e��/x�Sk�̩i�.�����{n���hH0����&�+��!�؈=J!|L�m��:5Θ+�CFb���E�(Ѽb�BH��Z�i6O>��q�Ryw�v^!�	�ΤE���:F�r�,��d�t�=�Fl�\T�x�gk�}(� P�:$��v��bФ���(�+�*�.��%L*u���4;a��}���ݶ��;�R�]biՋ���g`� ʝ�:���9����I�6�o��W6�9�����p�.Eje�0�I��Ԃ0]9g2��]R���3M��`���w����Ʋ���o�oF���x`Lq��U@¶�M��,=�*�B��#*�e9��s�9�&��A۞;P)o�J6���n��/�wғ�ܭk��3ܕ����F������T�^��C7͗}_p7n?K>�,�,[�P��嬢^u�'P�;my��@n�29���k��ȑ0�
�`4,9�@h|����I��i�hb���ckl$2�C��=إ%��GM+�`�&�gp�%HZ�&��������H���$�1���^65G�q1��&�r�y��=[�>x�&��V˞�o�0��{ipM����5��o�����^���^��*>��8`������2����|�34I �ҖѼ���8��sO���Uڜ�vx6�q�6�mV2Y۞��=��a�����HvC2�"�mkG&w]��X���T��e��O�lp�������ZW�ֲ7�%���B�u�a.Ʈ�Mk��Ǡ�;�'b��H^�zGl}5o�˨N��]�6!�
�z���oG�M,�a�Yf�^r3i��7��* ����ǂ gk;��߮=����=�~�<Ӳ}�"*��]��2�1Q ���w�gIpK��,n����:�^��/JZ1�͜p�ڽu�A���ĳr��p;��-�U��H�5YǬ����7[ڣDp��+��k��V8��U���� |����+ߒ�9�V�Mm�� ��]����euٱ���&e�`��/(���p|�7v)|�j��}[L%����6e�{;�ah)�]����L��I�Խ����*�βIq���
E=�{87���Ӷ��}�k�IZ\{s�2�$e�plZYR�q����OB�R��tJp�,ݗf�"#�Ӄo[�)�Z�q���,��t�0U���o6��M��[3im��ɦ�˦yη��)q�p�^IU�3MӶ3��������C�AC㩋���,�^�R��[8ξB/x0V1*/�xo��Ѽ1�{����ej�`��8LCr��d���,��(:��x��m���Y8.&2"�d���� |$��uv櫰`�E"F��gU>}+��5�*+�ԉB$
�O��݃G
y�;�)��po������:1��-r�vn��ю��'�@]=���e٬�\-�hK�`1�lpu�:M����*�-#�e�Õ���PV�=�Lǆ��{���RN#�L���kx1�U�-g�Y,N��٠� D�,�0��t��Ō�/q��F�"Kk6��D����yK>�(��3����#ʫkK�a���q�~���$g3)���J!5̖K%v�����'��_�Rw��V2/-�k6�X)���9Wl�*d{�ܦ�t���֝�,]$�ÈLr�Q�7}|�޺Y ��[���B�\&x�w5���~X|��R�4-l�����G[���{��ҵv�u�xvƃz�ipY\��E�fbtC#��{׹�,{����O�%�Oj���խ9y5%�+�T�T�f��mW��ݦ��lK���lΞc&^��T6�V�-�*������Om+��g6�u�&��M�tJS����o�9 �����[�0c�%�7wwRMj}�L�v3\����t����|�� ���CG�C�p�}û�Ga��
�q�w{�S�r=���˰SҲ��"�)��.�qa�tY�^ɚt�>��ۻC��-"C����V���ȻLǸ��[f�Ӿ��	��c��u��D֭����7��I{�PN���x�&I-�<�+��D:č��O���c�:�'��m^��-s���<B.VF�րŢ1E�.��^�
��;2��U�a�+�Ӟ_��������=�9�Gv�.����oe*QY ѡ��3�p�����:5i:�.�l2��VT�� ���Fa�ʌOr�i�>y��f��hA�2;����E��x*`�w�������Ԋ�.s"/D�ӌ>,6(���A�a�{q
�#�z3��Z��#;]�����7�`�P��W���B4�`kr����%�\�Ůd��@,D�Ρ3>���� U���)"�44ʽ����X9�Ŗ�!��mh������t�,5=û}4�5;9܇`�'�]�K;#N���)-dC�{MЩ2L͢8�ۼ�O�s:D0!׹;y��h����0s+���|wH�$	0�H���͈e��x�0��1wc�-�!�g��NP�V�s�����)�ԥ��c��}�aN��w#�����|���8*Z%$���<����	�^*���k~���;��}�ɋƧ;�f�Gfzp{���7Sӗ��wN��s	�ei(]k��}��(Ѩ0��a��PGX~;���~��<�q�*�W5K7���e������+��	�'r�ן1|8�v���@��D�NA�qW;1�T|�*l���[��ʟX����9�>J�m���늭vQ�ܺIl�}x����*/z)x�Z34'��f!Y؃\��/G[�[�z��O)����㱒�����6�+�Si�XeNὍP�7�E3�y	�ʲY�d�^���Rl�Yxn&�$���9u�����G�w�����#xoa�*�C^&gho�F}��xɧh�jPm]n�b�Mԯv�EWR�R���D{k�#8��GJ_r��nRm^�ॴ��V�6o�u��l�z�n��bo��m۳޺��0�YeoP/!�yV5b[»�=Bw��S�w��p
*0>|q�8��u��Anۢ�l�U}��p�<���F�C0(��(W ��y�I�����M��=��;�(��Zx���al���F�����%*b��[ë��L�wc���&��!h�n���uGs.�.����x�����IK��μb̔��݄%f.n-6vOM��d�6��e�^��weݛW�X����YI�-ZxU �i��;lh�v]��6�li�rؘ�u+c����ЕaCF.�y�@�up�����.O{H�*��x�ooI�����&�2��Fe#�do$/tl雜7Ճ7v�"�8j&3��#!�igsׯ,��jA�� ��t���1�iy���r ��h���p�-�ѫ�31�����f��+�s�W [��w+�&��-�³��!꥜�㧔��f��.���ٕ�c��8U��ʆ�:�%y��#��B����C���9�&�=>}�v�@@�`Q�R�z1`��ڒڻDÀ��;�t�f?��K�V��Z��ZFW� �v��DKsr�ϴ���h��U�K�H���cL!��	��tN�U��"�s��x���ǳ��u�E��1��R��t�3
64���vWe?��s�Y��5-�kj�V���z��f�k��o���1��t%*�nv��lJ�l���2E�m=	Z�ԥg��+U��ڵ�+ g��+vȧ7�Ӽ�/,Q�f�mI�L��{��g2���hR]������tg��
��Kܮ����Sx�qhx�P��y��N�i�hd��T�J���yf�s�Y�/�+��	^��n��Lҵ��D�8b�皋�����4����[:˗��^��#���+�[\���5Nq;7|BP���3ٷ1����Xкjj����g���0��6���=�(�����j��
���[�������a�qѸoN��\�f&e5���啹��^8���8�=�8ج]�2c5���	��э��@0�%[�����d�֛.����+��S�E���h��(Ԗ�BǪ���a�R�y�b��g*�N+�E5*�sK�6����u
���|��"��?ug�`���P���L��/ ���]j7�]igۻ�$wviz����x�v�΋��2�윷�v[/,����L�B�,��w�m�(my=�:�����3�e2���%Aa�ch��19*[�s�p�b^���kn���n�S��v�\{���t�D-�U:��ŋ�2�*4�k,oZ<�;������/�YC 穇�!�;�����{��@�(�������I����܂`�7=����d��l�����ڏ�Q���`�}L4������"T�ƶ��p#LQ��3'G�X���Eҍᇹ�<�$��dCv.�w˙ƏQ���n�����{x�@��2�Ńf�g#�/O�Y�p=��>+�>�n��NNˡ��'u�vD����-K��x�[;�%����q_m�-��x)1g����j ��]����zIb�5�!�ZD�y���4�S��ƞ�9�b؆n}���>�v�P���o�ڬ�ٲl��1������N��d�G�s-��Q�.��i�ot֬E
�8e���wßN��w���[��mv0ǚ75��9��_R+�]8�o{d��W��u:��м����:��b,R$ܾD]ݗD� �/�*>ޭ��zk:�<$���.����S��U�$�V	|G�k��-�5k++o�L�g8&ZF�v�1��S�_?�lMՕ�N �u��O\O�����:>m�t��^�ގf����%������i�@9���Ѩ�ݽ���z
��}E�0�=FxǇxP�Ev���h!u1���ᶅ���o>�!E�cz�͓���)�7x��!V�=J(=��E�����U�r���ZYd(���"^kf�����s�\ܜnf�PU�£��HE�K(�r�j�E>o+��� +�Q�O
�D��T+�Q=ym�TT6��bQX-�����h`�6��Ӹ���R��SԽ�FX��E]��2�ˮC�yv�Y�@�#'����!�~>�ms`
��na<��k�:�N�������;h�l�v����I��"�B�ծ�1t�q���9�, �K%�Թ�l��q��uk�[�q��GX�L��vgu�G��)$��Q���|�](��B/��]��^�/V:(v)�2�n-w\�������x{�M�L����ವȂ��a�V<8us�/���^z�O����ڀ8�Kp$�|&
.Am�t�t��@�]�WH�����,�澏��B|1��ɗ�]�iń��v���r����M\�@�5j�i\Q@���scG:��f>H�'��Uu^}t��n�u"p��B����jDO\���R��Ót���ێŢp�R�h(����W�fK|���s2WD��#!$!ǣ6����f�2���nsP���J�x�s�-���G�Dh�Pb���׉Y�	�_Wq2~��<���ԝ�����(��H0	�w�iu�*��V���8V���Uv�*E{EsM��fv0h���,�-s�ݹ�,��!Ir	P�
=�a���t��zEr��P��g	k/���/E�bnMem��������꼩�A����YX���]�;]��8U�҆i�(>�$�fkk�/�z��"Lv ���9nZA��M��rnF^`F���6��O;;s��J2'��9��Y�h��GOK��+��OB����p쥕j/�����?Z��Me(�Q2n��/}�ſ"e-�%[v���P�N{}��K}�1����b�<�e����ټGw���k8j'��c7�7G�]�¸qu5o��o���x<Ov^��T*`V's�E��v���N-��۹"��5�}���:�W�`��2��qN[���Kw��Frp��F���W*���k�B�r!�{�v�����L����=�lٸ�V�̧"��IdV�VJ���.f����d�";��j�9�qB+5vuG��a���b�;��=�s|�@�8���4�q�\�lM�Oi��$�x0ic�1�
��,���zC��V�w	��w���3�2��7[��z!���X]�g-kTS��7������*q���Ir�G�c@�\�,#��(7ט5hͽ����s���h���aB��>Tz�$����	��Ř�����Ѵ�3<�!�n�8er.v�^fP���K'e�`����R9���UǊ�GV@\��<�Mu�����}d���$�#�n�Ρ�PM�{��R�1z�Η��!7������˼��&�,\��|AXa^1�F��~��q�f���J��q�z;�JM�˦G�Ҥ�d�Ӻ���x�ބ>�)Z��c���������6����=�K��-��W�5��YE+�i����gQ���y����N����Ğ�5��[���s������5������E�Ms���ͨ�]v��_"�w�s0�T���A���הމx���f��Ƕ���6�fz��2��5��}|U��/f�n��
�{�U��X,� b�=���5�u�����!Rm�v7�޹���|o{���A��GYm�����J�e3�v�m�����m������|||�����I�2�R_vT�j��q�R�nq�i<�7Ɔ��z���7�p]@��`�/MF��jD,��!�Ϊ���:0�m�$����
�O�B3��k��MY�k΁z�d+M�y�.�h	]\�^��`�����g8�a��^�-&ژ��,��BP�sb5f�`�S�>87~��϶c�tݝҔ�N�3�m	f�r�H]:���糔������ �Q͍/=��a�|�3�WgP`���_?�����S�Z�hSw���-��/U���p����큆9j⺎v�˜� ��3��삘�G5b��i��.U�T��L�hGW#E]|�OU��e�Tٗ7�^8��w��!�����Vr�_h�IG�a픱V<m饧���h�YۯAr��{��EwP�kI5{���{2g-<Tה{q�{ҫS�L�(=~�fmp*4m��f��0M���7�\3M�аv����EN�V�)/�@Q|G�0��Z�6�B�L��y��+���-=7�������9�C���qt��n�}�ޥ�;��7/�g��Pzi����g4�XmTj���ٛ}�'5h�+[3'\��Ke��ԩ��w4���B�_u<��/��c/2���=�^�b�
y���S�xFc�,F&��xb�]n��H}_5������ޥ�v�8���uˊ�}�$�/��"�.�<��`�ެ�l�"}��˷e���JΊ��⦹���7xOFV�u��o1�a�	���nO<�qUH�5�[k&2���!�|t�/y�P�;��.�Y�RU�>ѹ�nbCK�����h@S"\�`�ygmt�Њ��
�ឬ��-�^4̇�ݑTQ�X7wu	Z�+,�i��nr��Jf��)��Ȉ+{�� Vَ�Җ^0�s%��^eA�Gel}�z��2���5{Mŉw3�mn�e7W{9�I��$�s��;�Я����>�T��vđ:/!��kp�p�����4i��[�	�؜/�E�7���G�1tT���f)8��������ͨ1NJ��f3��FC�A\cڮ�6/2�k��hR:��9�=΄dpf#|���d�wW�gf+.X�'O5�8�%��.�p�ӌ!y);�3y�QK2��o�9�v��=C���c��[���zn\|��
����c���B^��ڻ��X�e�H���.�ڍ�͡ܨ�+���.o8�Z�����i� �k.Q7Y���	`ضz���O��ɑ��Q�x�q�T��{e=��T��&_C��)�B;���5�/^����WnN�2j�.=������}4�H@���;2��	�<�AZ�m-��-FV�{����چ`]Æ� N	����4�G&�ҥ-f��#nC�Ρj�|�*C��z���{�"Y�V��{Gw���A�d����xB��㮾���:_C�咞�{�,q��ƴ���k'�ƌ�D������z�pR�e���Ҏ��p;,�
<�Z���ǉR9���.`^�5�k�(;n�::[���7�rUG�	��Ff-Π1��ek]l��^J�,�}���+����d�t���r����N v����fu)���V�7y-L��W�j��@.��u�]���$u����+�� �sK�dH�pG<c�v��)�|z�3�q>��V�8�G���ت��I�0V!Z�S�f`�癕��}܋���C���B���خ��
)hLl��f/M,vd&K�7�O6���V��V@�$�yy�sJ��/f3��i�)be3�3�������P��ʙ�������b�C�u��,��IsTѬf��iM�/z����ڮf���k��3����#WeK����cb�9{Gn��ttV���`�\���t�#��r�i�'�9ɨ��=O�&��a�ԝ�G�(*���\и�ydʡ����	�����R����m�.�6�_�EF	N��ob���n������iÂ�˯ֳu�k;�O.���/���N�V���dYQӖ�t��o�n�٘���v1��J�:��W�����3ͺ�t}b��춖��4�g ����-��vjO0��7��!.䆿t���9��2�a_f�)m�x�e/4�ޛu�
�S�� Fe��̭*S%9�]9�;�Х����X;3�-�t��(���X��]�ZO-�ɷ�������L�a��%��C�{H;�p��8���p��N�)v�c6��HzWh����[�)�Z�zs:�̧[\�c�^��1U6��� ��M���<�c�uY�B��Ew�}���xT[^9N����(Y������E�#Y'\�LK�̮�Ծ�`�J��}�j�A�[S]��g�
�Q6��!lS��z��+��O��ì�8F���C��s�S	���Xs�;j�:Ά��k�ge��T_hf��K�UYӽ�<8{JP�<�{uvJ�~6�*��L�ҕ�4��l��3�)���9�A3ݩ�aYn��sB����4��y�Q�����1jјn��U{E7X�Ů<�̐�urB�'�m����;O#��y���.��%������c͹F��W�v?me�-ǯ�;�"Da�܎M˰�eeL͓�M����D�@��#��:�Z���Z�w ob6�P��~2��f!{�
K&�K�<t"�s�T�]�f����Scq�6$�K��*޽&̀ks�gb��}x�T.PP�*��5t��Lf"U@s%(J���Z���{x�t���Υ�1������S�������[���g��U�s>it�R���k��
Xx+,��g[>
=+=���E�cK�u[җ�:Tf�f�cjy��m8��oMVsuDdo�c�Gk�[��Y���k����gVn��%��ʃ:������}�^�.�i�҄.���i����6��wj0���2�f�2�r�\���o�P���62*v�0𹯃�T���J��6)��b��E�8,z���_[��X�;�:ow8*ի�8Df˸��:��+�Ƙ�-��7(B�S�t�i�Z�T n�j�"���=�J�Y�s������ͫ�xL�A�x��ٱ�>P�Dq������
��[�	W]C��)RS�P:�U�����#U�w:��4oV�K��јs��1�5j���Xv/W-�w�6�h���9�O��t?*��6���N�Y�%�.�ڤٖf��{�V$�l���J|s\���'�Vw\�7R�	�b���J�sQ::��%��1S�i�c�
l
}ԗy�n:��v��ôz�bT�&����:9�f��חc�<��J%:U' �-[ŗ�/Lݞg�^]��X3��~YNK��e�wV����r�N.��gZ
���L\7xE;��X��#$逫�gA+3���|���n�1��oq�v�Dp��k�n�b��)M]���Im[�kW{��}	;��)&�O��N���(�i�(�R�V������5�sw�xT�����(Y�V���ű%|�'�S[S�]�![����;A2<v��K�.����8n�9�`�r������e�z�m gm����]����T�"�F�
;b�K{�E�{�82�m�w����6�W*:�nV�p�&�����^�G%���wd��뫼$��2���[���/z��V�絋�:gP�X^���{n�k'�vh�TTl~�쎸���`HghW�v�"_ZS�ee�LS�*����z!;��dG�~�9���-j�;ϨTr�>�ofpՔOro�Td�R�pS������T˻���j�ޝ�����v�4t�^fG�@ۤe1
���;�2ّ?��N�79�eM]7%,ͻ�ԹK����o�>�l[ef����I�E�߼S�A��Ύ�"z�D`�2�t;h�f�q3�8A�(:�뭝��s���3��1�Iuu�:�X���y>�j>�7oa*Moj���7y�Σ���mI�^o4��&Ӳ�p�!�N�+K-V 3`��g�0d����7�����yw*v�6�3e#;�+E�sJ�O���j�ooG�$=1z��kz]sP�J�ҏ��i��C.�uIs=��^��`�SZ7Y��류�[=t�]dSPX��D�nLH��Y�Xq����q���Q-u�9�y��&֤��7��Z&+��=d/�(k�/(=���Ѓ��+��i]���=���:T��֐Rf��3pQp�E���TqhIu�����9oiy�������1���6#����#�>�iZ����ˁ��v>��d=
s�4����0���h�X�]6F�� ��iR7�m�����PfjD������6��-[��E��.��Ci��1+4n�;+C�!���1o�ߙ�'$�$����	u��:�������t�.��Y�)�ԻD1�cU|uMO�`����%K�̕De�Q�R.��Gἄ��Q�n��97�2����et���P���}5�����_�B��k����^��V�����pд�v���hwFa��ץ��>3��a�R�jl�ޗt���F=��(��u�NP�晠0\�{����Ma$�y�Ż�+UӘ(u�V�i��T�[��(�SJ=�Fq�{�t�E59��L�3U��4��k(a���]��1!��ǳ"ê�C!V��;އ
�k ��pf2z��s��7�b�k��ae@`kX� �O1��8������0��W�z(֛�9�*�BV���]$m}+�G�zy�����#���e��1����S��P�B�P�i3{�,Ϟ���G*I샸��"��7l����l_�5L��2��8�����f���(���S}ċ�d=ޣ�����Ǫ-a�c��/��ٖ;oj�=�קl�c�C�s�3H4�G3�b�����2�*y\lڂ��9<�	��+�1����]��M�)�s��.�wb��Mv�g��fy�xX*B�me�AJZ�|6.�ZD��g�5<�X'�vw�^̡F�e�P��j~T��5ڔ�x�1��V���=�%A�-��W�'��z�W� �UB�_%�:��4D2�z�����{W��:|�4�s���d&��"zh�D* ��+��[�;�im�#F�[�2��H��V����ے�h�I�y�t��897�i!�z�u�8�J�@��C`�c]4�Wsu�=Ȩ��y�$�*̸Mq���Ʌ�����y
*f6���+q8����܀�ɸp�rãM_&�룥�ѩ*��aO1e�UiT�h� �[���c3�;���<�&9�>�0��/h\�8B'��� ]�e�,�I��'i�����e��=%t��p�w��ZK�O�c.j=Wym�lgZ+TC'���ב��9���i���iҢ��T{U�����Zs��㨒ySû�7�.�V�V�B�P���a߻b�ɷݯ���lc,�E
������j�Me�Fĸ�8u��@ˡo_I׻�sD�c��y8��w��j����nW9X�O���;���8oM�WV�7K[�n�/���3Z�`���/e�f�]�oD�M,����'aD9�t������j��-|�Y�u.Ed���2�������sF�X�b��5��Q{q�����T�&��`�}L&��(��i&��I�b�)p2�;U�����U��̙�Dm>o	x$4;�r�N���;Ƚ���J(Yv�<��8c�+2���3lH>,�pp�;����-��{�����f�x��is65JK�ܾ����;�6q�8�wh��K��o��K�G�G�,��[�����j�q
�Xi	ʙ�y>嬮�G��Y7�?Vn��y�`�M?��d�}���T�'|k�^��p�Ԩ� X6A"]��o�9��unֈp�n�ؖ,���%�%���-�� $��b�E]��w]Ê#�:��ƙ��9k�����ݝ���x45/j��y
fӍ�[� W�|�[2�wY��9��Y1Օ0�w1�}����T��ꝟk�[�;��fU���j��j��sH�I�9t<��ϸ&��]1�Tɑ��u7D�Z��W�z��3��Y���ҥ�{��k�݁�^�c(�D	�r(�5��fs���YMMEH���	�Y��7V	�)�m>���m���3�Ԯ�E�i^�_]�fc�d�g_9;X�ef;�D��jfge�#�!�E�/��F���'쬬3]�������c1Z�V!�o���2��
�'i�Q���vMg�	�E���k�嶃.�Ż}ۈr�S%4��Ժ�aq��3'".��Ӷu㗹(�4ڈ�a��9���~ه�_<�,��MǸ��S��<܇r���۩�r�*�����;�6��a�r�gGu�S�:�<g���LY:~Mmd�x3�L��8�Gԭ�Dq��M،�iw��݄�k�������˱rP�um�3{���`�1ŋox�y�v{��)o��b.t&�c�l���WK�`r�|��D�ͱok	x��2�^�5,:Idj��!�D{N�ee��M�֛�}/+�s)��i�7%�gg-�Kp%�b���<���B��3�Ѣ�����N�ghOu�c-+���
�b�y�dk��#�Vة-
�$f*�d�W|�� ���dY��?}����tdt�|��b���49Ӎݹ�J�<�fZ��/6�C&��AYA����9�T��$J��j�[��)�5U����.��;9=�^v�����B�vva�XA
�P����8���ůD8�Gj�R=���rۻ���	��_�ء�޾�i�?���}����麍B��~�{�m���,�{���Pm�{-=4��.�����|1�g������A6�����i���M�c�l�n�:8'R5ґ;g^��Ii+:��]����{u<b�G���}CF�=��^vz]s��XY�#��\
s�US� ͇Hц
�<���2��Ճ��4��P���͖�
��W���W�1�i}l딯NQ�1��z�ްl��շ�kS����Ӆ�4�bZ�{��N�/�R]�W��u�Jڂ�2�u�o�h�s��}xyv_q��6�]-	1�o��9"I�O<�N)sM`C]�{&���m�sN�Y1�O��n(��M��7A�W�Ň���olnF�h�X����+���sKփ�K��B��$^�0&`�%����u8��EwЁ��ց���g�k��f�b���u�%��=wKNZ��c2n
]�f����L*��x��g����6�o;�6�@�S'[��M{�;;��᷽�"T [���b�j��[e�R���.%f���܆M�'{7z���̐P�a+�I�Fa�ֺn>�6i�ʷ`�B�^�H��m6��9W�-�ټu[�S7o�̤��KV��a����$����^���ݹ|���j��}�$y�����]t�JL��V���^�����4��h]ж���vY����1L�D�E�J,�]�2�S�U��
u'wnD�!�G4s�v�Ψ\�T���4"�T%ZtJ�9�r�-BL�
T���J��$����!�9�JEfqI.:�����
�):�n��܂���	��֙,(�H�%"F� �hYd$���W8U.�J��@�q�4�ȹ뇕sS(B�4#���#Z%t"�**���*I�w#��sV�Wt�
��CP�ԎQUq͎�-V����X�
"��H��RӜ�8�0�.]Z�,�%ݮ!��AU�D��4P�YȂ
���du0��X"�f�����U�̽-D��j$r��fTkE£%P�P�d���9�*S2�J�Y&f����s;��-���D4�P+B��eZ� �hs��Z�7���_��ϯ"�͟�D����P=i
����o:��3�%��2��;Q5�%�G�p�v�\#����;�.�<��3(��{ Vں����X*�����C�r ��r�^S�[���v���r)'�P`� c�7@TC�R wo���s�n#���R.��/P��D����'V\6I��~>5���6���qr�E�d	jY+r.i�����lW❮R޵R����W��;=�;�l�qo�s�aF(��;�Y�<�e� ��q��
��n>�^M���4�t*!�l�f��ֲ��[q�r�>�c��{!�S�pp���I?������R�N�k�5(Z:�8j1��6P��H�_N��b�'\:��_h�o�^�03�����v�7�����P������Cb����gÀ��j�*8�3��.2)�Ws16%�Sj�\8z�p?�W���IX��S:<ꯥ�Vc���( �R�oO@wEO�5�� ċ�#t�(h�'N?��PM�R��+%��>sKvg��E���� ��y���ckF2p�6��R.�X�/M\�t8��0KPn��5�F�t �`d�3�7�d�%����u{�KZ��b�!���c��FxI�G�r�[��ܨ�!�.f��.����4�<�ӥ���,���rWg�4�I|g���Η��yŵ"�{حuӘw�]jO�Z�욚������8�5���� �yfK��y| �6:�{M�/��V��麄#T'�H�Ϳ.�c��u�eh���ay*�����B%[�/�W���;�� �l�W�L^�{�Q�$<���V���tɒ4dD�KA1��L.�$V�v�ײ����}<�&0(+�Ҋ܀�@9��{�(xӪY֟�S�?Y�%#��	����+~UP�0;��]�~�s�9B"��Gu�+����RT�\��\G���T��9�t���[�]�1JN��m����m)��]5x;��P�����V��^�@�t@gEv��>��v�/��UwF�\�o]ܵ`���0�*f�?==��;
�
����F��ؚ�Y,��G:����y�Kv���I���[�d�aHsڡ&*��^@��E>{�}�l��a4�e��s�s ^�=�-��
�Y^c~nt��@���L�"��'i��#���'g�'��ӗP��������4䥕�>��X���@�4�Ρ���)��
[��hv�W�)���-ь���j�.�Y��Յ��NMf�V�)N=ӒH��FSp�o��~��������!a����������ٷ'���^� F-�`]T�2�u�S6�	X#�
9}3į��cO�ʋ>�R���6u)�W�Q�^�׺�H�W��~˴���P�,ʥk�ϭ䭕k��5K�i�U�vǌ��F_���W�u �ߡ�l�9�}{qL؍�<�7ND��"�OQsXU�L똛�������U�=���&�~즞0^�g��ct�x��}���|�b�}�n�|�+�(�=snS}�r,Hqs-�ɕ��F����K���ꌴ��?\=��(S݃i�N���$�K�ڸuz��S^�F�c��x(��c�Zb�n^�5<�W�w��\uVl��P,)�{���1��e*��*�.�����>c�|mE1��Y޺����̤��4�e�1���@]5�(`�����G:5Ok�o�fL������5|���T�7ץ�t����Qn��nfV=W �)�a����x���ҷ�����w3�����A������u¾-�²�b��H��-����������m����X�UU�
��a��.{��xꕹ�'s7.b:���/���%-��wk�=O���^�Z�7aT]�� Zf(s�,U�G�����Q��;��&�Absx*�[�2�X�}*ds��84�`Ǖ����(׮ ��\�k;�A��,���Yw�;hb���
\X�|^6������Tzo79|��Y�o��^�����B��bN��]	鸁0����׮�xר���?V,rp&�3�j��}Ǯ�u�k,���ug�y:��a��H\�Sj�}��j����tݼ���j��V@� ?����*��f�ӛ�
�^��4A�Ʉ�BY��5P��"�&6�^��Y�E�����m4��C�8!�ȏM�g'gt��X�!3��͋V�Za^C���6!��Yp���@ƝJ772~��jI1��82�)�ɡ�2�I�d������o"�q�#zn'���b3�]�@�t�?{yr����pQ�v���]Ԏ΄����KTf��*�r�]�2���0�"�ڐ���b��3�s�n�����F;.L`T��'��6�q4�"(G8��ƇQb��w�ɖ!_ѳ"3��L�c��wL2��Prs03^[ˡ\�l�r>ͥ�ev��������θ��̡̞W_v�t�A�l�X��|�T����n��n��S�Dm�DR�V���<|�>�]ti�����"��>�<s�"a��8۫��m�J��8��v��H�2�!W�z��_u=f�3Uܼ��ZƤ޶��pϟ��=�箔4�#�0ɤ�dU�2�LA�.� �N*�4ؤQk'-��֏L�3[�K��#�f�tT�gf��1�Z]O�M������Q����8ܔVpQ�ɒJ� C�x�a��X闎�;�-/���1cG7<4Mrv����*�r4���B�7NJ1)��r�օ��ݫ.���|<�����t�Beu�=rW(~�S����*r4�����R��Q��jݭ�<\}��|�*ȇ�P�d�haa�Wˁ����]r��M��z���Z���V�t����oS�́uEb�V�{U���\�T�k�g�k�6�L!�o1L\7�l���r8��RTTnt>P��,X����u"��1�pg�2�(�nvN��Q�0rn�𵲗fm;eZ����6�@l�*
������=���ǅ�o�u����,����Y]�{X�e/}g�6�3��0���*t�7U��yF��8@f��F.����n��(v.��2�1�더(EDc��S~��ǰĩʈL��zdcOl醀=�{:�:�Ӭ�ܓ��l���K�b���,`�5�@�[(	��7��1������&cg)��Z�:�p-�C�ї��l�A{���o�=i�j��H5u�N��'M���{��T^��{��V��D�a���dmi��.wϫ���̄j�-եQ��������m�m�_pp�G����l�t١�����V�~=Ƥ+ݣ�c�R���q�)�ϥHë>���lWO,g(p��cC�`^�~��׼ t���
:�*�]{�˃7���	C6g�����"�c6Gh�к���A!z�����[V#��B���C�ï�Ms�4\C�ǱuB��hp;U &"��,%�lNY}�]�������ο0kü:����i���-} J5��Q2�-'�W6�����^s���F�臓,;|��q�Z808Gt�^��V���b��̼#e��b
I
���zg��Rq"1��h���%�s�����}��Gi�r0�v���NE��0>�ض*󩿭�����|�]ʾ9�弞�A|K�?*�Բㄅ.{�7ԁUH�I�V�/����nV��H?���W^<iЪ޴��;�߉�9��_x*�ݔ�|,��V{�v�JEYq�hu�|H��K�.:C,EA�£�����9���#[��������M5�e�C�n��t�c���\��VPp�X��@O\n(�S�D{w �,�2�E�=^��0#F�z�K�wg�%� șچ�Z���MO/�I鎚�����U�Ʈg�5�k&wv>0lɓ�i��,�vl�M"��J������W���G7�].�r!+�W(�nж�.=.�n�������������yeS� 8x��yZj�Zƥ��}��޹{�9tδ���?8���: �}"a�J�����I�7�f���T{멍5ڲ��F�G<z5��/T`VX�0ł;
�z��.��*T$�51��tA�p�v�����������b�>,�B���Mk�L uKq%���'�.�FToC�w�"���H��3}\�P� `N��r������_x,S޻��b`ᑊ�'��mO&
@b���4��"��0SYGL\ ^�լ�4��q�Q�;�w�E�y����k}��ʾ�H�ް�	�ϕϽ:��h�K(�ӟD�� �.k
��k�;Z�j:�����8����<`�=���3w����Q�p�`���76����|1Gpf���E+7�=�̐r��$*-��!5M׎��1x�Yg�"�X[o�kŖ��cQ1�c��r��
�� :����n������A��^�ܱ�ʵ�u5$�M��U�(�
�ky�E>&�m����*������n��q��fm71%-z�v���E�M)%��VL�B���ı*�����h��xWʩD�B���R4������Dm���4<�l[nΰ�:0�(m�fa�7_cx9IۦQ�o����,_'�ǥ�7�K'�N��s�f���ʢ&�2t��`fbuRI���*J0G��x����mBE��ٝ��;_t��.����;I ���q8*��ȿ�����@H��#�S$�|a���M��u�'�zsʕ�W�q��:[!��9�U�<�*-U) &  B�"87�`U�г]�%�_L`�eJ���.o���9��\��1?7wї$�C]&��N��x�խ��n||q�[&VZ������h�>A'4�|Z��䘰��H1N�9ܼfI���FU��o�r�G]��a��,E՞����a���>��ׂSٝ�j=U�C�kq�i��&ƈ �$�K��x{7j��O��~Ʉ�K��m�}9\uc����M�+���8ު,�:����
���0�\��XnL1u���+f�zvSn��%�W�˞��ܥp��@��>s<nn���V��G	��p8e}9Ha�0���v�'#�����������뷫�T�˷:��$Z�Q]��'LT5 n�/�ۊ�۾b���f�q'@P �p��k[<-�.���1y�3��w=��Q�$��G7��F^
ᔤ��9�J��aY/ ;�Zu��Z5���s�kE",��{�+�On�2��7o�qUv\�/�3�n��kC�⻣��Vp�aC	���Hx�:mr��$X�k/Baa���ރWΗ�*��L8��i���׼lk<!7�-/
�X��{��8��!�:4M�IK8�����E��ܟX�@�g���Ԍ�'�,򮿉���3��/�F��T�fݕ�ܸ����WQf;!�1�纐��l�Y@���	�o�;p��.TL�2�b����t��T�o,���:�8E�g#O�nW����wZ���
�3���P��Yy���k�z�=y�ʗ((3����C�ǆ����#�N���,F��,�׍�������;\�Tg)�V�t]����f@�q��X�_N��g��{\T�k���M��ٴ�j�3bm-iP=d�<1/�����T���:�	\c,F�i7�SC���)���O��/o3Q���߄��
���h���rR@v<*}��a��Tp���)�"cc�]}ەQ�Zq�{yI�ܲ1H��`����V�D��c�௸[������_�{�|��٦޴�
��
����F���=�Y
כ���}�|�,=�V����'�0�$	ӥ\y�a�Wn!�p)ψ��ʛ�c�Q��jp��qnŤ��M��g+v�լ1�Y�Uk.1.��|gg"����8��v��}m�Y�#��sL�ۄ�[��6W�F�:��|��P3l���IiIQ�2H����p�R�qꘋ����d�ع�#E���U�����׹�wT`����K�x�	��,���Laꉜ;�hxQ� �Y|bn�z/3:��0��nV<�ۥ!<k,㨬1N�W��V��ׅ󭸋}T���	�՝1��7��=�M��g�� ϑ�źV냨w��X�u(	�<)+y��r.y�s��vC�WC|��H��y��g�����]T6+���k���hxS��͔�++�S�;r�����-�n_��碝W�I�}���g�8���t�������ӣSxw�1p��S�B%����a���zy�0k��{Pi,h9�&y�v�vG�)yf	V�8�����c�M�k�
�E�L�{��5�2�Ty�(� E�u"T#!�|Kw����s����P��&Pv�|���v�t�"���_dF��4�2P�/Ot�-Q0���Rl�L0�g�F�0�֊ڿ���9�`?���Km��_�o��Ѵ:���P�,{�A9��'9��nk�&�c0�v�nȴ�0PZ�]r�?���]����i���srҖ����S�����z=[�[�\o_-YkK[�����;c�ʱ��:Y;Z|�7!��<�W��b�nW(��5i�;�;r��^�-
���W��j�:�6�2�r�J���.���y�yW�ػ3A˼_�*{�q�����'k���ѷ�\�՝�� *Pśk�;[�Wh�HurYva�Ѷ�.<�oB{��-�Ȝ���v�F�lĳW,\��`�9ɨL�\���RB5Vt��JD�hk���T�]m\vZx�h��#Z.Ì�ت�BЙչ�-!��>�)�����.b�L�F�+�ƧTΥ8�ñY�������e�S꾛"�������"U�\cc�,�[ʘ�s?J��oT׵gaD>:�X����L�kW $-���ۙ��]��U/�A�[����7]�/=����Ã��ҒR��3ևg.�E�w�Zt!w5{��*�PU�d/8.c6�{0�[ˢ��u������37�k�O:�˹,��-����xtqܜ����嬮)��
Y�CS�H�2�6/s�umn��)�����7p鉰���.�=�
Cu��b��m'p���삂t�L�y1�:ł��V%U��2ܷ+���tv��a]Ry��1��qd���<�+��O��+C�o�1%��r�P�>t�&lu��m.R�{|2�Fw���	�5j 8E���]���ޖ���	Ih���q�W��-^fD��)��%�9�0CfN�4wn�A!`��[�.�;�>�:Z��"�����1���i���Z�T����5�$�K<���eH��sY���<7{��s�e\�';+U�9r���J�r��ZUr�9�!�}��7;���nRuoA�c<��w-���+��k�GӸ�q���`�4L�r�
C|�G����'�,����2F&5��;9=0�>�OC�m�|�=��L���G��\�a轹�0�!.��T���\y.�+�LK:��ީ��u�}&���?`�(��a�8mA�6.k���۝��勲��Ñ��jA�ʏ)�0]�Ӥ˒�"��&�,�!���3.�;
y9�(�u*�]�,���s���S�s̡�_.q��eZ=���\�m��],I�8����,�Ų�}k�x�]�4�{p�֓bV_9sr�[�(C��W"��1]F����UCmM.��i�N3���f�Iդ����p0˾ʻ0�0�+W�٠p��_G�����Ě��d�a�${ê��yў;f�<3pK�H�1���f�^Z�j�ĭE����9pW]�I�덞�o�76��1������[�炚Skf�7׌W��N����u�ސR�7.A�U�E�����Q!*��w+`�3$y�}ꠥ{8z�:wę���W��m��밐Y�d��Ev���.���'�l8��qz��DT<e��WM--�b��U B:�eaR���L��I,D�a��.�je�
&j!p�Ή�f�bWI�z�p���TRt��p�Ds6T*�UU�]f�$�\��L���"9d�IUG.�RI&a�N$��蔑E�0�i�H�r�B�5\��e4脒r���5
���-8�!!��eΔu�Fbe�E�%�*�ڪF��	%�fr�����rN� A*���g*йI�B�"���4�r�R��!hQU�l�#R�*#Gt�T��K�����P�htLXQ�DkH!RS4�PFfgQ(��**�$*ᥳR��kB��2�� �Dt�9U(�fG9\�Tت��8�C�S�F+Bt�R�KY�+�Y�ur��Z;�GÇ����Z�֔rtYʻ�U���ym�FK�6��O�����Ydݸ����찌�f;�G)ݯ�mg<��N�5��g�M��kh��qg��=ü��.X�B>����-#��#�T�{��|~;�z�?�!�=��z�H$��g��;�����$ҡ��O�z����������G�G�DE"-<����1}�qC/��u��y)��T$:�Dh�� ��v�zBw����ϮN��w��}y��?������!�ܨ�B��q�=���P8����?�O}w�roރ����?S����0�o��2Yݧ#,]y�����Ӊ�++=�i��}����?s���{�zM����&���~&�Bt�+������r�A|��s��!;��C����v���˷&���޷G�\�Ǘ�<�?}��>�9�E[the{}��Mz���[ɿS�s�w��㾦�y߿-���®?����&����y��^�>�!���{����=;N�����xoI�'oG���+�4�w��t�_������y~;z@b�>+�'Y^>��=S�.��վ��n�i7��YO�oו���������=�ې��}���󷮎L.�����_cs����vM��w;�ϝ����}O����I�����]��"$G�R/�ߩ�]�[��ܣ}�I�>�#�������oJ�i���~y��4���ܞ��H{Mu!����������C�k���Ӊ��&~}��x���M���� EU�������8�o!�d�s���i������rzq�ߩ�{�7;��~�����©�����C�{C�����.��m�z���x��	9�r���������	7�$������T�Q��|,gV��TJ�^f������b�
CG�]�@|��_1U}����ӽ+�w���e:���8�x�����ӽǉ��~<�{���I�]��i�ohI��9������lDCG������/d�}�������HH}��ߛ�ߊ賓���L,����?�Sr���ߟ}z�g~�N?7��';~��ގ�ǉ�'��q�����F���z��|	����������b���J�ޭ�7�'!{�� � @����D�D DF{]P�@�v��w㾡����{���
���OGߟ��������J��ӷ�ϝ�=!ɧ�?]����!�5Ԝ�&�Bw԰n�{�������}����b�[�p�;���С2)�E8�|��h��͔Ù}3?x�˩�;}�(�o;8�t�Q^��.����XP�N�uČE�L��Sf����t���NyD���:�^$�lS�-�'�;|�c��TV�x�C{��o,d[q���	l��o��Ķ�.v�.������ �C��Ǟ@}~�&�~��oC�]��ۓ�ǿ��}O�\O o����}NO�������9��;���|>���]���r!����Ă��H��G����Q�~�������P��M>'8=8<q��!�=X�ߟ�oG�ɏ�~�����o������m�����]�����l|q��t~�oI��6J�1�ۙ��n��>b"D} n�����	�e�������=z���;N���o��7&����c�C�iǠ��C�������=A�7 x����;}g{v���������������S5q3�����r�!�`��D��{}�q�#�O��6��=&>��
x���ܛ�t�D߯�z�Ja~ ,�y��$��q���������������~��0�V���ߞ�4����G�����h���=�?"i�O��c�i	i��=����1���z�c����w����������$��r��,�_���|Nq��y���?��}w��|��߷����}M܃�zw��B��>�U��*��b&>�߾��]�����;~��?�$?w翾 ����'�����x��?�{�@�|OA����~|�s��Sr�|NS��c�]㴛���J�6�W_��]Sn"p����}� ��_�������x��!���?�!��q��o�`���{�ԓ!'����;{NC������?9'oX������ri���6��N���Jv�>��U�b|�1*[�">�9?S�����M�c��<E��;۴�>!�����J�M�	�q�����~?�	�S{>��O�oϱ�ak��n��7��x���܀����>���~&�<�[��H�6��:}��r�+�"4E�I��}�����'��~!�0�����y�7!ɇ���+�M;��c�x�������+&����=n����|B}|���o_��;�}:q�b�|�����>��0k}�C��O� �㴒��^�x�����ט����?�O;�޽q�!����Ϥ�0�������~�Ʌ?}w!��!�?Ov9��A~��=c�= }I7�/_����+�
�>������K�R�q�f�é� 8��ԃ���BOHJξ	����Z��O��咝�eDs֥������W��ji�����D��*�'us��8��|)#[9�n�Ǔ�q,�vd�V!��1��?�U�I{!KL��z8} �G׎b(}}.�� ﾼ=&������~v�"��C�Ȑ��w+��&���m�'�N	�=���{Oi�aw�����o��D����� ��G�"��Ǚ�>Ն��>R3��c��"=�cF��D1}��~?Sri?���v��]���~�oHzL/��/��bOH&�}E$]��ޜw��4���ߏ?�w`S|B�b<"Ə��b0�����.���=���b���#�>����P��~��C��x�w���M���H~��9K�ߞ`��w���'��������P�����='!�@�>��α�H#D|o�鈀 ��#�4EsW�ޑ(nk�5�ws�u2�w}����"4G��^�����[����׫ۃ���}v��~�!�F�|v�C���x~*aTG��x�q��S��'����>'8�u�H�~�M2"ׇHJ�8V���y��Z��G�|DF�#�c�}��i�߯����o������ۓ}B7�<q�P'z�o�x�q>�X�C�94��=�������"��}o������ܮ���q�M���o��ү� 6o�U��݁{�}@|q�|����nO�Ʌ?{�i��|�8�<�����oםɇ���c��� |I޿#�;��78�ǻ�<v��]����7�I���??�}]������>{=�U��o���2�����ӿ���|BO�o�w�p)��?~�v�x��$?�����;z�;~[���|���9�0����~����C�:d?������<p|g;�"gc|�ɶ�]ϭt׻+ �"}"4A�0�}��?\I�hro�x<�����{>�q��H~������o����|�߁'�p)�7߾�N׫����?�N�?�����I�z���@ G�~����b�X�5~�{��������8�q��zpH|C�ry�o��OI��S�Q��!�>!�����T�]!���w��|1�8�]篿�}m���$�������ۓ}O�}ǎ����?C>�>���H�9� x�M�_��߆�=&��9?����E�o���o�/�r��$������t�qDP��1�>b���������Og�p
�{Iǘ���!�0����AU�1�!U^_�j^�5~�3�}���N�1lJ�w��7�-5@9�0�`a�x�Ġ��ܰ �7�x��p�m<LH��*=�@����Kq���qRm�uۦ�I��0�;]n�䭃�/O���^��%������0�|��1�u���">2@����D}v���3����}�X��I��v�t�������! xts�>�w�s�u���o�������P��ǯ=oj�Sx��眿��S��	?>���?���<q{���ӵ�7���������F:�G�.�i�|D} ��@��q��~&�{�/!������8?Y��?�zO�r�_]���O�{C�����C��+���PrĐ��̈́!	��[�*���Y3ޕ5z9wU�0�vz��tC�W�S�R=�- ��ؘ��մn4��aR��.��U�YYwx��M��x΂��� 5�����U�*����DvO<F��L��\�N����%�q����10�>\�l�j�h�D��p�%�d�ȹ�#DHb���U�:L�N�r���n?�ة	��|4������ϯ�S�{�*����W	���f�B Xoś����B�~j����նhq�~5vy�a�b��e ;��1��n"����{�B�Y�/�k�u����U��R�y�`�Z؉ʆ*�҅���Ѐ�����y�ng!�T]����(MD��kn�bo�&���^B�u��
���U<�̈́ ŲCq.���W��JR�V� 8��nBw���a����ew>��g�ty�_I�j�z�n�a)�E׃����a�ٺ�V2op���T�)�:�u�r�L&d�V6�M*�D��F��G��ќw؏3biJ�c��y�ևU%�fHf��@�iě�W���Z����:���kO���]t�b	�XJ��g(�f��+ﾯ���2�=wYt��)�v��u����;"8s���a�,h9�7��x{�R>�~�>��O,��a[���DT�oT�@"�y����Ɗ�k�eƪ��5�{�+~�4��Z��8�<S��wN ������a(>���we�� k�=�!���'^>ձ�t����mS�|�(�{�J�����"a $k<�m!
�衱�6����u��ԣ2�u�R�ɜ]������Y#l��~H�=e�H�_O:Xr	��aw|��ya���T�^ �4��ݜ-�ǻ��#�0AF�n��Yd3"9d�lͽ��*�;�~ۘ��gC}x�R+���ӟ`n��a3�]����-Ԑ2
�1貄^A���:/e�I�[X��Ū��ٷ�-�ӟ��BLW��S�8���+(����wP@!qΕ*�'���#[�	���!�t���a�qe1� ���D��,�Æ~~-r�=Z��e� �슋���s�u�c-�~���uϭՎu�^�p�E���Y�¸�*��kvӑ4�U�r�k$�՜q�>U%y��2�F�e6���눀�ͣ�N�S�R�1^�Yn���B���e[��p�WJ�á8~��\�	'cn�_4BfM!���9W�|���O��T)��[�9a���8a[˲>G���.\�xT�rn�������E�ߨ�@���D���m����o��uٮ���]g�5�� {��`N%6Asٵk*�"�3d8�O_�bF
�k}Z�N��{p3�c��
�߷�^��x<J���s��1���1��bΰ�h �a[�@wϪ�fّ_7 `���:b���ҳ���Q�������:4�q�[�b�0��O��`\��^G�{]�a��sTt�ϧ'fۮ9&te9+tvM5��)��;y3�b�5�F*4��<`���xtͶ=����Z pu�ڞ��*Ż׽�v�_��S,��қ�!��Gre�Y	TP��l��KG1������_I��y!��|"�����w���tx!W�S���i�*��U�����S3֮)R��z��X�jH�:�������C��d@6Ʒ!��A1�� � m��*�~�k�=`�Oq9���B�Ln��Syp��x�$�PJ������f�3���e��k����[Ec�Q���O�
]w���q���[�r-��!` $DG�9�6��;ݗ�K����N>��h����
v���^٣�7A<k�خH��c�ԕ+�jZ y�0զ3&�ߊ ͥ6���b����:�v�e^i�Z�pݕ<C�	~�����T���xA�<��a�Ӱ���}��D}��rԳHt �������2[5��t�zUՕ����$�B��7+T[��r����u����0Ys�b�u���~U�M��QyUh:�Fjr̚�e�o�9F�Yo	���p����/J�k�/��i��H�'�[9�ѩ]m��T^�Q�����Y.\��W�0���R^ӻ�%���X��<+��Ve����m-�v��X�&84� � ����6 	��'�Qr�h6��څ�/LUe=�&��*B��S�����^L$j��CT�dTG
n�*��81�Q��~C<)Ne*��~t^ʭ~ܷ�mqʫN���q�5��Fq��:�n�O��yGD�7����C�ś�h���/<-1Z�/fU�s|P��3�짎x��|��@���Eλ_S�7�*P<a���ܩ�e*��'g��J��|����e��W|fy�,�����KC�09�_K���u�Z[e���nLXڙ��|:���Z^��HU�ͺ�d&.5b�,����)�Ƶ^��/�z��Q�`�>OAR�!;�W���',r�#�5����Q���cdT1����ߏV	RZ�� �Z$͔-�,.:4���[�\�N�����[��Cs����`�fD\�fѳ{w;� ��I���*�DDDE]�î\9�����tX��-��>S�`�R�?�κ� �v���sE�E&`R������¸�쯴0��9�c�K:_Z����	[tٸ���]��$r�~��$�x���{�8�r��6�zh9l������_5V�vM"�!\{�fkF�K=�/���n��n�ʉ���册`C��8U�)�F1�Kg�2�T<��.�ո���I@P3�M�1)��B2�f@΢�)d��:���Lk<.��Ѕ�'�F�<:�j�/���F@X�j�D�NQ1�Ĵl���GC�d�1��(:�Ҿ��e����|:��-�U���.4�t؇��U�@+wpF}fY��2WN�L������񙆼3��|�	!��W,�.��Wbp6���܁�P�Sy`;Њ׆ˢ��n����ea��b�����`��O	��+ʒ�N�)��H�X�� JrʝϮ���l��9X�J����bߨ���qpͥ�`I�҃�Y����=QS�ậ <�dA�) �����A5ƸD��3lŭ�;ف[ K"�?x/�]�S0�L8+q����@"2��2֔n�6����G-M��S��z��{1[�����ߢ��> C��k��.�S�7�-�:)�V�+�i
��=|<�����B��6��/n�W�_UU{)��
q���ԣ���bǟ�Xb���;��1�)ڈ���9���v����GğC�Θ+,ͷ�[������*r�
���q��@��(�Q@�;#E����V�I%��{n|��e�c�an�^B��	���y囈 ��HA��*u�{)ۮL�B�w��:�ֈ��_϶��<�r�JŜHh�K��ub��+8{�~{j��`�tLd���$l�T.v��ن;3�_n���CC�Ǣ�F*	����,N���������W=�@�_��*g�q����,�7��E���t�TCn�2�:ܚr�w^�V�f�@�.$�ip�Hui�S�J����{�U���y�3�6E��Y�9�|]b�
�[�}�8�܍י� Jg<w�zЊ�:"�����E
��喯���GH��b�F:�������gh���)���iO��=y,�Za9уl�5�BC����'(!q�@�Aҙ׌��(
�5��0�����݃:8G�KB������{0R��>������"�%1
[�m��i:���v�����N12�]�,C[x�CB���n�Mi8�aB�N;L���b<��*]�Уc�5���$�+9�j\��\�T���9Q�O �TOPt\�s�H�W�>���"z��η�^����~Bb5��(�l�Ӏ�n�DT[�"�rF�)��;)IhVHo��oU�󈾝Ù�)ӄ�4����`3h�=/(�o.*-�AX*�]���u�<f�(�[g=J>���B�����9C�ʭ,�U�[����ҥ@b/]!H��˼���_���;�= ��o	�>iV�����n�s�/EШ<Y���<%C��$��ޫ�+�Z��(fOװ�E�pl���;t��|Ԇ�Z�ay������m<Uo��'l&��p�y2Q�Rz��H�k�}Q�$�t8�{\�����w���;��Xc�N�9�K�� ,K1{ʡ��`��m�܁����* ���䡆��-չy<�<�~ov���<6��Iͻv|����hu�9�u�׺�����́P�k��:���W5�a;���f��V����^����Bq��<q�LL��m�P6Oc.776��P�.a�*"�q��|W#al�~�MSGW�Ys8���
;p2ģՂ���X���3"�U9��s��g(�	�si7�bys`��.j�r�d� bor�����W΁��U��u��S.hi�+^1��O���j� w���:'���o�����͋�  ��/��GN	�{ڑ�ɅW�Z��
��sg:nV.���aǁ�]��ɤ٠��Z1�RЫۜVe��>��C)>ɛ	}h�v�_6����l\+�1�d���ܬf���7����w�VuL$:�Z7�bg:��}w�)@��6�l���P�f&3��-�c��'p�A��ӳ�d��݌�ڼܠ�(�(������A���t �f�-}'t���W��e�q%���u�t| ��z�D���*O�����Clf�r��R��Hڬ���+�*Ƹ;9�8��P�m�*�a��Y����m'�F��V4�"��gʋfC��ڜZ��+�����g5�I��v2b�؎�w�;�<І�j�f	��9�6Uf�� �isT�;��_���p��v��R�o>��EY�2�(0#Z�南�W�B�mg�^[}�p�#��ǛYI3��6Ȯ�y}�pb9�U���V%Scq�9���B���e�����qA���]�y6���Nݜ���yI8�cC=��5�����������S9���~(��*}���8���K�������Xٰ/i�`���n���:�O��_�@���H��p�9�p=��&� f�	B�^�zz�5D������ ;X@f��7w�6�	Y]4�v�����H.�(���:&v�n̛��5�$�I���ww�LvwL@`
ѡ�5Y�Eņ�.
�-�j�T#��&��9���4�,0-����!룚hmn�Wc�Vy��bn���[�&�i��+I�@d0�x1�S�%�8���/���"��D��O����|�Z{�Q jr��"r�$*Ü��8�E�ݦ�-��\��ƕ��6dtsgr�*	��$
�����y30u@��O�z���I��,���+�:bű��ī�d����52����<-wP�8�����sJ�מ9	���;�Y�&gB��%d%�&X��Z�u�	�IZݞ7��*�Sk^��<��O�0eN�YiHv;�\�;��ּ պw9��ZR��c���'y֮tV>!x��m�٦ã�����)\�ߚ�%J��T�o4��
Q7O��0tQ8��D}�N�]ȝ.r�L���Ǜ���^��S
�;|6�����c�%XJ��o`�V�Uw����o/S�2_"2�:�G��|.�3b�̧S��+�ֵNc�S�՗N�u�c%YR���.�oE
�VǮG�|���!w��]��#�W^� �L=�S� ��k��L�`����!}�e���];��S<yn/Ius�;3���"�d���yk�4M���ܨitU�ق�Y-��Q͐�ChՏ����>C�A^+G(�r�͖I��w�D*r�*L�&Y�E*AS��L�R�͕�:�H����E�^��������$Eʏ2碝"��We�P���fL��7��<ɑ_-Q�2!VDGV���G*�R�9AY�L�8�U��*��sj�+�y��Nl�'�er�����Tr�vz���kH�P��3g#�E\��XTTI!�Vi��Ң.Ye��5*�TA��(Uȯ9��șqč$���L��je*�V�T�*�E��rx��NsS
�Y��8������	+L�#�PUI�RW����E:�YE㪕^fF,�t�����^dS��s�Qr9"%2��PA���ʈ�VTGu����6��p�K#�aB��X��S{�O<o���f�i�h[:�����Ug�%���xe��DY��E��a�����U��1�]������CQ��}���z�V�)����SY�N��pu3�W2����է��I�GKp�������Xt��B �鍶�Q�_mKu�<wǰ6�:ţ�/Z)��7����R��������g���r�ގ��lq�H��N )����iV�.������V��4b�������ܑ��s+��؄��@�h���X�����X���Nɂ�b�ƳxS=�,J���f0F��®1吤:�b@�]����J�Ì�1WK�����/�'l�����w!۞��V<K�ׯi�Z���a��yބ�º�<1���W�ט^���/�M'��|��.�����}���k*K�N�������!t�1`L7_D�T��9UO�dM�-��S9'"��\��J�S��m4�����k�qp��CRa���v� �rt�%��3a�v�R�?h�78c�R����ݏY�T\ƣ]ٖ�)�ʁF	n�uIe�8Y��Y,DL"���C�\��]���ȅgn��#K���@�rjK�ws�M"���p��5��ţ1޳|p� �~n]�RP����(FU����R!8�=l��ܕK!���x�)R��R;����K����KE��p����� �u����$,�3U��ǯ18�*���^���d�x�)��tl�����m�O�ۤ�d���*r��g�,VDc���b�DoNp��:�uؙ̫�sm�r��b�Y"' f�r^JU�*�٧<���|���G�/g
�_d��璵��-�<�)��=�\:뽓�]o3Ƙ�M1Vҭ�t1�.g�,BͧyEB�Ѯ���V7�8!8��l��P��;������.!�Õt���X�џV/eIb�&�)T��մD�q3�q�<�ժ]��9�c��tƋ�+ő�'��;!���<��K��7�ֆw_��=�~�~�xbGx�˟\<�L\a��m�P東�9EZӑ׬K�d��{f�>��t�ػG�U#j]1�a�����X�5��6aj�|���؂�6ߧNvq'�׽*Һ9�y�.1ܯ�*F�l����#�~9F�yP��mL�xK�"~׭\��d6�۔�DZ§t���	Lv��KF����)��g�����/��tR�J�Q�]\	L�׍Ȇw?0sA���,�Li�"�7\���ǖX�,����B�%3g{޲���Y=����H�c1p��m���C�yqH-]�{(���@�vرh��˼Z A�32b�j�J��w$Lh��+�b���ls���������ꣽs?;��c�l�!5�V:�D[YU���+�Ia�Jً�ι�[u_f^�"�2��0v?���i�b��r�#a� �޸�=��-�_h����^�Y�v}s�8�"���R漬�$h�y���	���0I@u|�ֳ|��e��w�f�gVbb�����.❮R�{�k���i��N�ާ:m�����t��P�M��k�(D1b TJ+�,_|c0�Q��b,،޻�|k�꧷j�;n`��<zOW�b���ζl׾�PT���:Q���'!��%op�0���C�zr�Oq�� gL)��H���X.��M�!g%%�	�+]O<����+Í���u�n�p�i�b���h��G������u��-+qJgG�����Wgos3Z���0���5�C���!���w��(h�{�t�  ÷BEgU�V���/q�j���Ӫ�'�}p���Ez�8��Yxm9L���@�5xf1p���~V�W�F+jwm�X�z�
�rӻ5=m�0s��ݐ�SF|p�No	�1wQ�PV'��;���ؚdR�?cN�8,7cs6��O��WpЂ1��1�.P����ku�&�}Jaھ���p�� 潞���k2.QĪ�\��[��s���>��)W>X�T�������<#+��N�_#���Ϋ�@LЎP�t��N�q3.�_S�9U:}�Q!����d"f�C��@
�Wl�+u�2>�T*��O��װv���c�V|�bV��0Kv�Μ�Y����;&Hc"y����m7��ս۴)$�\#��\h��:H�3���+�z�w�.��+鸣��G��x��Yn��~��I�~�I$ f�b��ww\Uª�͗���Cw"����$W:,��VNqLov&er�̓����=9�2�wNA+BN��m\1�9�f��5 u���Um޶��sx�Mlu<x�VA�����1�#l�?_Kgp2����IS��ϋ4�gb���J��d`:ޏ��iV�����n�s��1*xҳ��5�x�j�tڙ��+�+�h�������j�6ȕ�b$�t��MQ��0��j�_"\5{ԕV)�7�#C�����TQU��y���?�z��"�r,u�e�|fj�ay)d�eҾ�O1h&����{�Vb�y�i��tZ�4=b�d;�滸[�C������(�J�6�s&��2鯸�!
V�,�޺鑽�Ej�"[�S�|6x��3�!�̐�R�t��1Q*���$���zx����A&��iL����6m�/ﾪ������T�}�n��Gf�� T	F'y�0L+M�A7:4\B#LL w\l�lՉ~Ț4�e��=۪�OV?\;��TkE�XT��z��l�:����5��b�wD�	�P��l=�u�]�R0Xt��q;>�ig�L�*����V r�V�3�d�l�[w�Nw�����#8eW�[�(�8�s5���h��|Vtĉ[-��Á&�*�C�l�C';���;xy�S�bk�2��#��e*��<8����\��g��������ll�|uI=���C�k��2xT��B1��k�b6����� g[�&��ۚ��n���7tw�Ϟ�4�
1ı����E7uq�(��@J@�-�j�$c�p�lm3�5��Y\p;�fL.(_�']�"�#���^�Y�OޛB�&h�f��u)^�Z�^�ߥD�_�AZ��0�	t@S9V��f�Q�ۈ:��0G��T�RWw�0k�gP��y����x@��߉��
�
�}�I_>U�b������M�\��Ol��+]��|l*^^�&2b�i���p��6����_Y����o�m\׉9���g)��x��y��4��ߔ�K�>/r`���uڳ�\�Մ�3T�Oe]��T�=��b��\C�i����v51��m�範���+<�x��Nd�Fw����{.5�\�b��d�mG;�6�� lu	�;t�֚�4��:A���̣LA�]�O���.{�l��#+F�&ϫڇ��5 ���+��f�m�i��G]����S�~B%!1;�x{u��X��ٜ#%�!�����7��UP�p��Ԏ0��`ߐۛ���Jò}����3ҋ��cD`��\�f���q�3��FL(ڒ���fē�U�ll�*������."L1w�aY���(2kLA�p�)�d��J1�bɬ��qQ�ʕ��u��1j�CE�V�8�V��/f}|�yh�2�:��^�X
yc����Ǿ���NbKD||)�͒#�3	d�1¨͘�a��)�H{���\�&�}R��Ć���d�1p���������F,f�"2�f9����Qs8�5���ݮ�3c$f��݌�����e�c.�ƷU�Iֶ�,��+6�;�j�}P�S�ka�\��g��p��S���j�xr<��t\'<�v;�4Z��W$Fl7@RNX"j{CvVՄS�����ɰFϨ��{}�WK2ȥQ�Y������/Cp���r��a�زr��-�iev�WP�e�T�#��Ӥg�I����n`Lr�PƇ~S��g�s����
�ׁ���f&#�mړm���Re�a}_}�}T�)	���˴���w��C��E��|����ac�ct�(E9�l^%�yT�5P��7���q���@V�u���� g�0��Y��K&�;H�8S�:��q��g�r�D|���B�t䡂0���K��m���嫘�}7;z��ĵdҭ��sWp��.VmWu��ON����1[�Lv@�٨0t%p�3N���e�j�l��3_{b�O$����wh׻���b,<:_�ހ�����T��#�Y$����^�5cqâ���W���8�����6���[9�1r6 ]3t-u"Veuȶ����<��Ǜ���4Q}[&�J����LX��"$�ٸmP�y@|��y\���V\�UA��^�:�d��D�V	A��[��^Z�f���`ϭ��6����YS6*���v[�u�$�� ��I|iѵ᲍]�u�
y倧V���^2�a����K�̹x�xq�a�z��Ǉ��ޟs!������h,��Dy���e�|�(�����`ة� ]�Z�4/UΣ�.���px�n�u� ����۾WS[G�I����2g�qηrff�ε�l)�LW����d[�ke-Bv��J#�)V�F�O��Q�ZN���3��i�h����9Z�T�f��eW��W�l�p�=� ,B?�_W�Wԋ����+���X@����������_7�����bUg��g�{��3��/�zuo]oS��Q gW�L���ͽn�E5u��_W�`��3����BuE-�g7�%��U-��~"�� s0���o�v�:B;����|�;�Vkv�u:���ؼ���H=�0@}>o S:W�U���+��s�d���r�\]����c�� +�N�(�����f���{@R77< ��(
;�\^�§֖�JY�w��1'�Ⱥ޽*�by&qf����f�O�sV{Լ����o�MW 3�;׏�%��.���o�����c���M�߫$����}`a�j��Ӂ_���4O@H������x�k��)zR��f)^{2(n�ڍT�ㄅ.{�Cq(!x�������eu�XP�N�UoZ{*A{��I�N��~���ҧ�z�r�keg:��>����*~��9D3�`^��њ�F�O>v������'�Q���9�+BM_�������[w/�*Xk�Y��<�Wf�]�iouf��R�u�:V�[W~�9���^���?z�I�_t�N1>��(��Y���n��j�r������̌�
=y�4�fo{�_e��h���g2]����z�nx���/�ﾏ������1��.��� �٩B7�rD�;�����$�ϵ+ysJ@��RIꕵޓ�]�].�|X�LUa�{
����tڭ*�u�>�V:��������מ�m#��\�xd��a���)�A���0;���"��'��^^�/��vk����+��ܝf7=K:��e����a���G9�N�Vy��?��#�E�4䥎���mGK�����H��ҟO�oԇ�<r�f�c��09�A�L�2*�0TC���=�^|��5���ڊݻH{�얊�k��ׇ�*���V�	����>*��וފ*��9�_��g���;^�ᙖ��>�j�<�����*��F���O�*�b��eq�����K��sl2��36���e7�H���r7���1��D�������=����%ا,�q�.��{g竅4u�zT�{���WߠC�J���%�s��5<Q���¥`\�z+YݴΙbĿk�5u�2W94s6q�~��F#��~P.�O+����㰨-��o1�cO��;�#"�&}]������NR�vv=.�g�'�&�h��+��HZΥl��;i�s�w-�L_E��vT�:.Ǻ�o���Q�1Z�r�Zɋe�Y���Z�
�Т�������r��}�r,>��W�U}��b,���������ʺ�]�ꇡ�p�Q/N�`p�yPŝ���$��EL8���XoZ�[�-�e��~�;����l�϶�#_ퟩ'I�Z���R�<��FT�L�yO�Rt
��U��<���1 q|c!���K�QbUv_nc� �	������Mgn����#��9,(0a��q3Ja�T��4��2���j�ƷO��z�a�8��!UOIE�9?"�aw�T��Mx�T�H��K��,�.*����<�2��1wU�ʐ�H�o��@�����Xv�����.`�H;��Շz��<�]��xP���27�S��b�j@zȶ_�؀rQ�5,v�mR!���"W��8k��t�����kƓ�`�)]��L��e��d�����s0���E�]9��f���7]qf���&��G�b��NRND�c*�{�N<fTi�1�N��3���u(��˧s촻z�`P��K�"0��D���P�m[�v|+�+̫�3�G�S��ߨ��V�=�fzK^Bx���M��r�6c�b�P�m�B��EB�g`e��O=�ѷn|v_o����	���F�w�g�oE�4���'k���_G,e����X	n˨��²�|X��[���h!2;n�yK8�� 5�CY8D�>���ї�,�l�O��F���X���)�5X�n�.XIgZ"�n䲕��&V����z�tNߘ3w�y{4]��Fe��3��DŽu']��my���$�L�q���Ɓf���)���]�p�Yt�c���;YP*��y��{��_��"}�"�ݧ��#[FS����ye~{!Û�3�4�!(2f%��q�]�bb7�k��EZH ��e�cZ�Y��k[����M�؛o/�4��\&���>��s'��B4�N1Y�;R�$Y���n^K���M�<����`c��{i䲜1��)K�i��s�s���Q�ˀ��c"��T�W��";&�Q5��ј�9p�+�]�Vʣ�/Up�o@J#�f���x_p��>՚�a�`�mӉ
X��oǰLu�I�
�%���~�it+v l-�r҂�+nLkf���:�f��3P�l�s7t�ʏ{�iM����]X��;+E�����fo��r\
3d�%>%S{�a����3
/q�"4��ft���0;h��+�Ma#Q��	��5+=�o)��
� �*����`>y�d/�K������2`��2��i�qdo=�V���ߘY;1�_�����NY8E���X��u"�Ps;9�$I�70Ū�_���:u���l�{N$�bT{:��>ҋs��6�������Zص( �ZnZ
4.��x��:�o���S��F�� �9��D6��������]K=���=�7cz����QN+�o���j���m�5Â��E�����<0���z��9x��tSV������{C��x�i��[����W���x{\�V���Ҁ
�:cb ��JQu�Md�q���1�V��V˼|�ѵ�uv�f��x��A��&P�-L΃�a�qj��%���%��.˨Nh͜�Oc�a�n��K��:�)ѧ�A��7{��\
��d��X�,h�ul�	[{.���H��������-���J�L{ՠVcq3��F��#K��:�.�%���\X;�흃=;{W�Gh�ѯuṋ���-�uwm
��qݞ*u�_a�2�|�դ�:��q���,���nSvp�Z�T�~4�<ˮ�8b�釪~Bt��9ah&��V��	���YE��;������z�vA�aZ���Y}>�wW��J�:^v+߶�N����q�U�y���(��i�o�>�2�f+��/�7�kh}Ȝ��b�*����'��8k*�P�PGtr��"�9U˗(�=q�l�'qݑU��TQ_��x�J��W9A@�UPA;���\��QU/!�Ԫ:`B.�&DUą���=6���I҈�3�P�K���#X���tK�"�3ID�<ꉩwTD�ux��s�u
��*yB�z�Ag�Ĵ ����.jFi�<�\'5N�2��2��̬��dL�U�e�'@�)K�r�D�LN*��r�D�(���^��w�* �]�<�� E�#C;]�*Q��$��@��

�W(��*=����A��X�t�����G<:��ui|�M�@��)�g:�s���ۇT,��UBHtȥ@�B���!=h�H�Ud�I�ԉ2���Js*9.R<�z�G��R�,�E&bsr�C8��L;�Vz���_)��A`�F�1W)��Zb�7�[��ϔ�R��m����ŶR���qnp4�U�#ﾏ�2��ʦ�)z�P?�������R�f����K�
����Q;(^9��@�֩ʛքu,���W9Χ�r7h@%�	�����(�p��H��*�5�����][�N��	W�zn�.�y�]�>)���Cr֍������`�����o��0���*�r­]�=�Pŕ=PHh�̡��ܪ��ȼ=�S1�R���֧=R��k���Z�V;���	�7fG=1��P�<����E�Ҙ���k��]9���ջز�P�(u�������È�M����-�R�����-���ѧ��Qǚy�R��E!���\Ɗ�X�\n��:a�^�#q�XJ~S�����ڸ�I�M��z��V��������\:�y�:���f����
�KF���eI����uV�nhtݽ����a·x��\X���N��;�Ọ �L���n6o��m>+d9d�߯�X1un���C21�S�U����(Ϗ �^��'?4(����O�������)'SU�<T�f�<��k�bjc7D,�cw�u��ޘ��eG�޾��V�$��SB�1�]���nFI�(��4��J�t9B�ˤ�5P]Yُ�rEt[��ܮ|^�� �ǒv�f�q��Vĳ���B�3L������VQ��-��&�/�U�}U�j ����R�w������1���u��}�
b��Y�#��f�H��/�Wf���J9��s�C]�@u�D��e���l\�3�3;�\�_��0"d��f�F�{����\}����d���@u��r����2�fg��3�HҲ���U�ʷ���0:ޱq	�ry�����1������ʄ,=(p�8p������6g:�Ţ�� BY����j��{��o`�{�=�/!g%,A��Һ����[j�<���#r�� �Q��7�����^7��-<�$^h��Tt�F�+J�l�MU��u��j]Y[TY��XTF��T.vɷ�v��0�Cr��&�L,�[��26_:|�(+��z.Y����]��\�c�����M	���I�eq���w93��WX�|�!�����1��F��L�5���D�O��ώ�X�H��1�eVod��+s!f4���k��n�T:;*T��b��
�k.w*�v�f��W��4|̠U*��Kt�8wJu9�[��;%�V׏Z�*pŗ�> ��X�OF�c�m��x�v�cs�fn����X��y�gr{��UsԳ+(��α�Xwγ�̍��mOPP�Oݞx�{doʹM}K��%/Yﾏ��>��ی�X�y���N㔶�g=0�77�L%Qa*����K#�����|6z}�ؗF=���_�WM���n;U���:F��U�I���tu.p�cm��}7���e_>'��D���d��:�5���*�b����6��������F�Ta�xu�Y1\D�ya�e�W?w>v����g����Ų�D���i`tJ�q�b�F0���ʋ`Įɨ�ݰ�c���r��T�bd��I#=�N c���C�[::e�٥�����.^�_E����1�;���݃X9�j��}pT�
�����}���Z\�Hk�s:M��|}�h�x��E�3��!+�q�8����D7���z����=�O����D@��7ŧ�V-]�>���yT�~�ML�>�x��o�����f����@é<o#���O�u/m>��Օ���Ϳ��;��t� G�O���P;��}�Y�G$*�Y-�C�pr����|�^�sX/�x�
wz����8{�!�tk��ۤ��7X�O<��5m�t'���[Ϫj� �י��s��O�u�W�9��˜ؠ-�S�#�|P,�B�WY�������!Ox��C}3�6��Wy[dz��8���ך�KC��Ԅ���uy�ue���:�T�:S�7���{�%}�lw��ms�=9�]����;f�0�>�OSo��}��v��Mv\7���ġ=�%A�u���-OM��հ�&�Ak>���.��&p�\��hɣ�F"��L��Go��O|�C����O
�\���ťq���[Ni��q�H�2�^�Aꌗ�tvTI�-��^.��iu��3���ϱv=g\�s5��BW��/�)�X*�_�R����*���n��=��$��5b`��*����]n�uE���)G�0�|!\���.�����HZ�����v�W���u�t�_7
E;3B�hW-��泖�]��o8.\:H��˞l�������U�TCw��e�C:�x���y	1�aʽAm����	��PĐ�$='ǎf�m��ߣ�sP���Ά�Y>��x:E㲏����lb-, �kެoeŵ�r4 ۠�A��h�[��ނ�����>�`�AZw����ALŹzE�%r� %��+'p���Y��e-;05�� K�e�T���s�����{Sb1�q�{}>�Y�!b�j�oT4��@m��n�w��*�X:���Z��84���b�ŀ�'1�v�5Hu�=Pv��j�n6�i�=*.na��m:���T�3��`m�A�eE�:��r���f7Tqo7�z���V�D�[cg�^���{��Ο�y6~����B�|�h�[��N�EBs�pg�'F��;)OC�P;��nzZ��I��f��[�V����8�]�|��Z�WRʷh�fʝ4�OA�OcBս˄�SW�o�r�4ݍ���f�4^�A�U-8�SFg;.y����V��i��֝��ֺ��v��`ĩN���@Nl�<k3�'�S�&��b��p�-�,�w��U�<��0���Sݛ�/���	>���rT
��Ky*�E>K�S�ϝ�k/-�P�m	��p:�B��z��q���B��%�AK�^��}}�=�1W��|)����H_��ɷ3�{�Y8����:22 �˸Y�JMz`�w�����,�+����,��ϑ�v��SvjTf��+"���Wˠh�]�����ʸ��^��EJ����fش�UOe��]�R�Y�_PM�Źz�WN��\���}}�L��Z�Ҡ�g�an�C9�u�YW���в����Ws�cv�8����>Ph��	��׺M�y;�d�:Favj��*'��Gv���`;�g�x��CY�w�Uȑ����2�S���:������a�U�+�y���iO&k���Pz��ܡ�w(tUY�ô�M4���������W�'644ѥ���ڱ*�2�D��A�vŏl+��5Q�|��������v��`涧�[���)�nJ��ܻ�=�b�f19���6,BڄٍSq�E;�ɴ�D;�k�S�@_�@W_�l�Eey�;�c�����Y�9�K�}������)�;M�MCX2��ۨ.;(⺷�rEf.<��OE�.)(4�٫C�-�Ԝ����u{�f�Y�t�����[�P���[�ni.�d�__uWأF�ɽQ�.޷�P���=���N��`U�9턽��ں9� J�(�zZY���ܫ��v֨˗�ʐ�;V❊��v�E���d���9��BiW�8}`뼗�ե��bc}[�[Н�-��)�/Mf�%/���
�i#T����;G�П�j}��(��je��|KU�ւ{��U}_WԵ����j��A���8�"�:�Qʻ���6*������+W,S<2rL�s^PތgVs������TmkUg}e��Wio2��=ɮ�[�޵H�5�m�C��n�އ�*�w�'z&)�Xy�u�4� ��L�����_?/H���}��򪽹��:�y�ĥ�����Ho"�.�=W��v���Q���ѓ�|(.��wT�8+���4žW'��tB���^.�}�P��[l$�n��3�fW�w�bd�9���{'��8j/UԈ1]ve�bs��Q���m�)�e!'9Wy`(��Ju�t��E�c�<.LW��yٖ5g>}�"vq�.�v��m:�Ѫ(D]Y.5�Uh3yl47��^tX{�O�������5�g���]ا�<�6�����W��T���do-)q�)�Y1o2�.�Ɲe'�݃���xbB��xz\�ahm�bTY�m>�6l���z@Q�d�o=]?� ��Sei��i~j��,��Z0/1���\��M�>���(��>�rh�w
Ν1���d]���>�":��4��/�sgڲ]�
�a5�S���\�Pi�
Ø�GV�UNr���˖�U8Ķ��8�UMDj�➣��yN
�����r���G+�؟��y�3���1v�X�y���n�yV8�qg�w�zU�R�prᬇ�\Zм��y�}{���T(.:qC�R�N�Te��v�A*�Q��Wb�ڨ/r��z�/7�ս�+l�=EC�g*�q�X��!��m��n��[/eB��ol��{Ǥ����6�+�?m��7����U�-�![���u����^��7�S�N�Қ�㷾[��5�jTI`�W���Ķ���|~����UCz��Ps��ҽ��wd;{P�Z�땶�Ou��U�|�X��:
�W�N��d���R9��p�+�}�i<����!A�{ LnU�M�P,*xa(��Ȓ� ���Wы�_l�M+�\w ���'��N��++�`���nǠ�mz�L��5�����ZcGA�^�T�_�΋���1WRC���a��8 hm	;vh����\��H�����㾺K�g9�|�:��.e�Z%��\���;N�_�]�tr����g��%.��n��U}��_iQ<��ۮ;��We\a��rʉ�Ϯ��x��gL��v h���ve�<��BU+^�a8K�)ؤx��0�G���ek��(Mm��٩ט��ݾyz�sU�}N���o#������*�;nQ��O®9��2.�}�9Cxs%�[��;�uں�z��s��A�T΋2��k�Z�ܭ꽡a�5/�����q�vŎkVO��.f��a�=@%�+Gk:r���i{=�1;�6s4��K�Exb�c>��ڐ�?@]Ds��Vح���eVt��6�2�V�W������^��:�����f1A����j5�nW�l��b:��MCx2�|�qב��v�wד��1��W������MX|�a��ؿ�x�ϻ���i�9���p�P%C�H]����Um�nSY�M8IlNM�^����!K-��'�M_m���,,�v7]<gcmE�O1oiO�R�ε�^���u<��Y�i`W�u���{���t�����e�׍��m��7�e�.�!>�&�2�����suϭ��ޅ�Kad�^w�sh�	��k!f��Sg�K���:�wͧ�I���������}�eeYΫ��Zo�������4�������l.
�_N<Ʀ3��zV�VyW�_;�*�Jyi�ݎރH�=��d���}���.7��=�Uc��A��|�l��S�K�f�t���-�wq/��\D]��V�W֡U|vTD�0R�W�f.2�A�y�S4�N��N�ΗS�.3u-qٝ�8Ɇ黎6��	p�Y_I#^������j��׌V�7Vd��1����Z9㌚t�镐!��*[O6��NH�Y[�1�=��K�v���̸��:�[��G7p�-ؤQ�µ+�s��o]�ϝ�O�+�V�One��/௹����qI���q����L��Y��i݁pE^��4��{�vX�B��;��I��!�O�
��:y��"b�����a&;.��٥���-�X�&�����V���m\#�#
���U�2kN[���(������-;C�b �p�%>91�L��9���^��@��(���1���t��$F$2w=�뒌_H��00�k���f*=�5��eC�����9]LWGy��X4k�f����ǜϦ�n*�U�{��:��?yL������#v��E��]�vۜY�A�+� ��CB�&I������N�?tG\��ΗB:�O!�31N���]s �ED��=���8�9�78d���Q�I!�w#]��F�}١*����\�I�k��>S��J���V��=��Ww���ņ�A������~�@�ŨN�v��!�m�+�UG�[�cX�B�Ǎ��`&9�سH׆�Q����F�L�:<xx�*\�p���yj<��~'Pŷj#���Ӭwm0��8㙚��+:b���\��u����1R�%�1�:�8����#Z#M������E��Du�Fnn�^%)�{��xq���m�c�Í�1�U�7�s��"���wSd��$̺�)u��疘�����Ҝ�#*
Bq����<�m���vu��.B:=��bk��0������H����(��|���ݩ]��T!����I��[4�K-��F���N�<N���y��kH����z����į^��w���>��	��+�6%���/�]�w[=��fD�
��&��[�TȘ�Y��n����u�V�d{Ħ^�&�d� ҷ�P�-u�-�ξS�:�/s+7L�"��Y!N���m9�+v�5��ݥv|��cy:��6O`�;ۙS�x�mr��C�+z1,�%���5k[�&erǯ�G�x�u�W2乣�k����������>Go5��|+K��[6uǑV˔r`œ����������Khw���K�w �/j�R��W|��%��nj�h�
+��U�F5�˷�1(��]\\���C�؁ō���c��e'����
�籱�tB��0i��Z�0�h�7�t�պ#:�4�$cr:'q6i�2뮻`��q�n:N�%�_�fWS6�ۯ{f�#]s�f��.���������j����+��8!�+(ϕ�O��4�h�ra��wŚvc��`˘��t��pj/l�$�5E�F��x-K�s�<�ծ���Dť�,f��ԣu�%Jf���R���s���� �1�[Gk�[j��x���a�;=u$��.d�SM���pzq��G�������jR0h�Q�!:�zn��ڽ���j�! ������>O���U�ŕR��o���u��q7� ��35ꑁow,�ֈo������e��=h���XT��P���b%�nG�2=y��
��
S��
�L���2X�q�ipk"��5���=}]��1�i�ӆCv�N�$���7�mC��vn�-R&�#��E� ���.�jίZ5����X�[�J5Ĥ[�Ği��w7\Ubp��2/�J*�w��P�*V��r�(���r0J��]�(-OA�ݨI�9'˼�xW�q2�֐G�G�B�9��/;�Rj��#�^�UI���:�{μ/Mʴ��dRdt��X�I<��b��!ch�8�������m�/�TQ�.��s�C��r�At��Ե��|y�K��#�*�3E��Y�a��r�S�{��yC���w�D�Ե���(�/˺��<�*�G=wl�K��T���͙�G����vz�(�9ȓ��K�t��u8�ȁ_&��Q#��^��K̓�;��y�^K��Q�Z'"�l���)"(KZ�7\:C�aN���;�EAA�������F�$_/�fr�	��U8B��lH�/�*�xT\*�	0��I;3"�|C���*J�����R����M���CAa�T��c3]�Ngq=��f멂�}in�����<��=�:���.rΉ����c�:�}��^b�y1��2XV����un���kQC�v���{�[�P����پ�� �\�N[�Ho��x�^-�э��6oV���j��o+��^)o�[gʲ�i^�r�����=�ƌ]?�먹Ψ��_c�tu�Vj��|�����':dч��Y��*P���m�n�Է78��:��4���6)�}��J� :ꅒ�!c̾��v���v6�A�j���v�]�5 �T�y٬�7�]0�U��5��3�Յ� O�nuc�wӻ2�f%M���a��&u���zSˌp�o����k���0���uCc���%5<pOT�p��i��؛�׏��vT���p�n1�Ҕ�8�J�r�� ���V��p^�c�Z��rz~;�*�<����鯡K�n;U���S�G	�:K"-��[l�����[�b��A�gD �1q�s*S�B�U�������ݙ1�No��@P�K�8+t@�o+f�x�-����X�m��K}HЬ1[�C���xz[���G*���|O���Vk2l��]����3w�N���9��֋y˱`�/k�UU}�
�_Z�/�AO��VL��Bo�%>�PU��߯����\���-�/�իd,xj��Y��HB��ĭypf_�\����-7sRtV@���֩Eu[�.��1JY�˰J��`��.�Sh��;gI�u�q�ФS.Ca����m��>��Kj�Gh�lS�}S]N���º�����ޠ�T�I�}qN;����Ȃ�nv��#[����-j�Ggc��[Z����J��N�c:�PÁ��c��^.$I��[v����A�ukE��F'��T�n�N8��/��rks�0���Ρ���e��ʆ�ܯ������l[��]KϨ�:��U����bۈӝ�y�RV ���O��0�c��u��!r����y`���V���l�r#��v�O��w�M�m��ԳVn��w��݌�+�B��ե�0�=��Z���t��j���Z��ij���������U��mWA��`�q��7пJ>��*���{1b��旺=������mͬ�8F�ߧң�q�Vx^��P*�.�8�7��T�zB��9N�HE[q�1,B�着��U-���>�����_s��o)�7���SK7�Rȍ���8�*��#�zL�].����=6�}�=Ŏ�4�:E��vl��o6����U�t>,v��v3��-D��#%u.|�)m�ۯu{��2��u,��-�8t�����|��0�|6;+�.J\*-5����}�\�T�+Yt�n(�dK��DRO��ɧM1L��@�Y_OL���as���i��l��	uN�Y�;{����q��&��oD[�1JQ�a��
���ĭx�r��r5��wt�������Ͻ�<hzo��C���[�?R�b��.�����%�@�xpXc�2;k;�g5�K��~9���������Y
�u%c<; �8�G*�<�]�s|�����*Xs�x��ջ�;��N_�M�U�X���^&�ڷ����qz_�ivٷ���񙾰W��Y�t�C�[v��u�/$���v#���(g5<a���w�
f��Rb���K�9��1J�c�)��<�*���:��x^V",�<�Y|�m�J��d�#�)]��w%X�	��̾oX�W΋�+��+����Cv��v��Ř���r�.�R�)���n�){����󌮍N:D�^�2v��T/�,��;��u�����b��\jb��'2gy���4����AU}��8��Ong>oS�7+�㲢+���'���#Pv���.���]�k����z��/K�7>�36��Z��+l�QP�q��m��r�a�7�Ա�/j�|�-�'�f��6�7����Y�o!��-LdɚԪ��W/5mX�V��N�-���71�;��kq��G;[�f��B݁5�3
��t+��-uE�ƺ��=Ρ�p�}3�:^&�OFӝ�{z�M�OX�I!�.�[���*;*TN�]>J�S��Ϟc�Gc�LJ[݉4�P2���ݴ�Қni��_W:��#�G�D�t���=��Cڬ(�b<�1�=TI�u�N6��5T±�l.�#5n7��K���{^ԫ�pWx�U�J/��ox+�4�nY�f�ҾK�[~��9S���֫��%�1�9��Ժ��=.۩�R��S����ku���dJ$�7ՑQ�lU�����J&�.�n��:f�q���4�\?E��9��_Hn��_I�����lߥ؛����=yսC�����ܐ�2�c���:�`���W�٢d���7(7��y�ω��H�{;�ͨ]\�<���t]�0p��L���[ps���6�u��\A���ĭ̸	�XW1��o�þemf�l�Qˉ����VAT������:G��+�U�0��,{w�$���%@E�x#��+��;�2V;>�N��ؿ��e�}�iuE�+zv1`=ZdQJ+�!u��*�K����@��a1o޼�y�ԧ��X&{��'����WD�f�f7\Lt�_j�➳�^Uo����Xۨ���SK=��9{������ �7�m.zuFDWR��珃C9�����˙�\j8����.��=Vl�EZz�.�>��b�z��Ψ�������]c��$
:u�;%�C}3ͫ{�y[w�mUd�Q��c����/*c5=oc�͈���ˣ]jD��緺�,�}��f�ݍ��A�~�!v�������5���`���w'��� �s���@�������nn��4vI:`ԓ�o����Yث �{�q�;1�ٝ�5�1�s�s�އ�������<C]Ĺ��1�_���>�#��l�C�������
�L��0 �:<�s����V��_}U�����rz�_����Oۍ���o뇱*��q�Pgz1<���:v�m�h���z��)��8[���g��ۇT:;6­w9�+���r\���W��}M5��<O�ZW����v��ut%�Or��z��R]NGeIS�k�v��78�B}����q�����6D�bZ.�'ZB�Ez��Wwϊ���ބ�DJ�q�ݏ���/bԚ����s���o�7Jm���)F9��B���זfXW[j�v����w���8o&����k�5�uCv&���`�t�=�vd�2D���j';3���:��Y	:w�}pUÇ0Գ��_m�Yc��큔4wL�.��<\f1c�ד��U��㸄���^uC����*]p^Ng �z�Y����h�L�ƯP<�<�����]섮�Ʃ���yO)u���g&�BM�2*˷x�=;MRl�.`�A;�7fs�c�t!��w̴���o3N��[k��1p�z$ �}e9��'nI+a2�&1rW[I̻�T-�h"�fw���l����}_e0���X�|xtv���hqj�r�}
���yr(�����IY�"����.;(⺷���}��Pk����Z�}5�\)3�718\~��Gɧ�/Uw]�����j�Ψ�9�-���Yf)	�1�Y��7V��"�����zl���[dz����\ⱍ�f����u�t��8ᾼ������Ы��{�]v�s���	TA�U��R�w6��I�o��O����W;�;P��z�bv���e���l�{�]o���L�I~)�Fc����DOo�u��4�{��]�Ss�R�Ց]8�i�y���(XW�����JQ4�+�%uD.|�8��1���mVWKե<�:�26A�sI�q��ᄣ����.�Zk/J��'kV��7���J�����a��r�Asl��0#RkR���(v�i����+�CV��/�>�Q}���͖u�y��8�_[�����}�u�>��i�ߺ�{ggË3�k%���oB%��
<==Wڅ瘣M}�h'o�0b»�D>#�X�����-��=�����Λ��R��/.��={�,+�L�C3|�j��£�'h�dD��g]@�4���y����2�kwax��vh�v�2o�娦E����黬ꖱ>�����{2�����{�lu���;�X�1�t���v�V8�n
��~���g���W����)�Wl����}N�5�
���2�������~ᇫ;F߆6��h��� �{>Y�e\&%����\"r8H9�l<��=n e�=���ѧ���+�mX=��]��c�j
�ň�����O3i[(�;�i9t����_��{�TE�:��r�1xt��sv����*���\�a�V+�Z�P�·���������v�G^�'&�k
1�N��t3�b�����Q[���������5�t�QS��h.I]L�#���K�,#�Ž��^�c�K��|��)�{�. ���>`b^N���6gK8��r�71�ӿ���>w����$NtVm]�[��
��>��Kގꅱ*�֍*.+Z��ʾ��ީU�<�:o*�g4K�++�t˨C�M\�����V<k�j��u{o��V�Ocm#��ȃ���t���~���q��h�e�7�n���Z���� h���hb�U,ũ��f%pO2��V^ev8��e�@�K2���������xI�Ҕ�%\�[�;U�&����h�p�͕H�w����M,޼]p�%���gz'�|��)�G+dh��f˞��k���qVg�h+=�o��t^�'3{�|�t]�`�F{�[�{�#%Йގ1�Z����T�{5�si_��q��t����W�J�B�;��c��<o�ave��Wb酹�k�M+�oB��)r��(�'m����Y�2�r�P�)T�UԊ�f;Udٖ�����p�Gsy]Y�s5��=�y6a�z��B̈́�C���3�U�%����=�:=��b��M[p�M9P�K�t�i��Ý�eR��o������yS��О���T���Uè
�Zc��_h�y��ޑ��q���<K�/���t�޷�B�6�5��t㿃���W_�o���R�NiV�u���Ϊ��ŀ��pb;���RS�v�ʚ��Z�m���8�~ʼ�{7+����")+�z��kK���R���Z�im� ��Tk����^J�2�K�O:�=�\�Y��70@�i���y�Ei��X��G�����l�t��N��Mu�����R��Gq��PuNb�f�f>�p�j:{�~���|�q`~��)�=�c�*r�1=5��u��v�.�?C}�UF�J�b��'�QmÇH!7��k���|q]E�u}o��F:�q��2>많�F�/DL�n<o�3�ޗ��E�ƭ�[w�o'���*����G*��SS;�e�A@ogp���=�6�����lC]��3U�iQV�cMqsx�p1�%�p�ԙ�ĝ�N��u[���t���ˆ��Cؔ'x�J�G��3$i����j�Y���5�U{�����j�)�8y�ۍ�\�hY_7�,����ƫ��Ֆ��;NC�݉�\�L+z�������d�M�xR�8Em-U���S�	GC���
\-s�Z�Ī���Z��&��[kvf(�)�(�O.��ΙX+�
��/�{d�'��麟 ��)��3w�yS�Ԡ�[���\'�-ؚR�W��\!^}\�ya�c�&(�A�iY��]F>��3���j��U��2��J�`�i+I�����o�'�;���2T����u��=.�ݬ�E�/�/�=L+iތ���\/��&�*���/w�9uUHS9�7���d߹��F�i����QZ��
yZ��e�I����J��<(��$��v�+�o��2�W R|dk5N��f�+kgGɋ]��b��v���q;|

'_qϺ�p�^I���dNɺ�Z`sN`<5�헏X̠��ǡe��v�U��B�����c�d��z6.�u�К���tv�7���M�Y($u�c���w]�`���m�=�`WF�u�I���\IÔ�����U�ͼͩR�bk5������-Ї#���ޮ3LȸQ��[M9�*��@����9��.�{��@���PltK����{}��������?J�~��]Z�ǥ�i-'�zoN�*�=����;W�>u�����>���+M�0��2er]N��3�	�+�Wэ���^�q�
}�ח��I֖�'y���!{��5�c��M$��뻸jwSU�.��|��ZٽIrB�*F�v���Д�U7HF�ζd��T��9܈�췁K}[Y �Ǵ�C|����Ê�%����]�n��WJv��	��'&J��tZ6�ή�y5W[�Q��-�V��#pm@����;s���'�ݱ�\����P��ܕɒ�e�ԶO��{c��n��t��k�;]�h����I�+���Z �{K�ݕ&�竚�cu����p�����m :J*�u�9�S�v_8��Q��#o��N�p ��팤.DZ�qջ�i�C*�'��B���Y;�����BʘۙYJ���q%�(!
�R�a���d0N��q%�.>�{>�#�-L]��6Mgy�o�	ܖ�z�=c&��Yf7��͑��4y^H�%���\1�cZ�&����pWimшvGE��뀂J��>���2�7�csUn��;��><m�9�'�^yS޾�U�؅�Zʫ��tM�2
�	A�V��5������Ƃ�פ���:�5�ݗ�Ͱ�-� ����yr���3{�����A�5�u����P=�Dfiβ��$��gL
��#�B^bѕM�tlb9w���j�	Qm'�ak��%�_d��͞�5C8ڍi�w��C�z���?c�E]#m94͒�.j̘*|�*��D���UV`9`p�Y��G�Q�2�m��z��{�u�\��DamdH��m,�}EԂr����W����;�1����v6��9�/bε/2�6��6��8���a=\����#w�wҷ��9�4̴^�G�sڦ+eR��O-� ��(�D����]`�Y��
8Y�e:�U�����������Y�}�a
a�����o�<\�5[� zC��{/{���N�4>�p�]�eg%C앻�d%.�:}�� c���4@3��.��wv�7gO]�~z��L4x�&��I1=�͎��Ov�%��NN+xR����twi	痭WR5rJ�\��q�ݑ�/;�!C��d�R<�zjo���0���G1̊H(�V��R����/!E�WSS'q=\��&��W9i\̴C�v�Pk����NW1;����O8�E��K+��r]��3j%��C�*=�Ū�+���^ty=��[�T��s�I�*�/R�s�%��(�۝�P躲���qۙU����r�2�dd�&ig�*�P���g*���||/��G ��9($"�8W=���z��#S���z�E�=e�e�wy��$�Ԋל�qE*�����^�NI$�����-I:�E�M�����QWr�ZAA�[����[���GD�����j-2.���-�yגX�#�K�����\蕡�)�AR�j&�I"Y
TD����&�C5D�1�&h�~ ���<%��<����+<�9�&��)v�t�h������ݱ���7�*�:�c��j*��S{�j��㹽�	��="�I8c�+x-3_���I���,���=v�z\G��=+܂XdK�p�T�=I:v���W�����2�{dր��P�B�/�7�Z�)���0�/f��rB�CPިh
{hv.w��z�����jwu�-��@��)v��O���N~J��j����'v[�rCL��V����e6�X��n]Aq�G�}o������ΣO_��3�/�Ns���)�#0[�ێ�!�e|���^A�vs���Խ������k~�E�칸O��i�B�mu>������n�qy��J���[3w�qAU4(kZT�V�F���n�yzХ�����v���}��f�m����(/�?D�q��1����+�9�����T�D.��Zk70��[yru�{/ٷai��U�"��׌��}CZX��D��)�w�'�7�����R܊���hbO��ъ;���\���,�&om_6b��y�eޗ^U�ϥ5���{8-<t�ܹ-SN��W7�*~A�8q3��ާ=����Ip��4r[�:uX��;�w����w���z�;%=ص��%O
��uV���F�%�a9;%vO�1������TJ&"�%y+��ϝ����n�b{\v�[3]��)�_tU[�1���	`�Q���\��TZk1p�����Š�{�0���vbY��q�ꏗ�糢��e\a��G,����՘������6ޱO{������qů�7�D'�,���x���j�u��h$�����f��v�F�ކ��w�}N��:Ἆs�>>4�s|'C
��n�32����;4G[��'�&�1��U��̻��MC�n�r����M�-$��7n���/���Ko�g�9�Փ�E.fM�F{rm%�K�7՛��*}�jd�/��X%�o��U�+�mX6�=�.�2o���-���3\�.��A��g2����q����}�}uv����P6��)��6^���ͅҹ�p��SP������B�.T���i��MJ5NLW����7�*;E�G/�3^�!��Jq��Fz����4�A5��:��\@�D9��-�Bt�[�c��1nw�[Z�a�1�!���\�-�(����!iao����i҆wy�WXC��Y�l���v���y�Ў^e(΢,�{���xL�)�7�[\�v�}U�
������kty����~s��j�{�O��0�G��Eֹ�ʄ#u��L�X��缾������\��Q}׼��Uޓ~��1s��;J�����Ĵ��T�!�7p-�v6����Ug����9�>��7�8�fª����ݞl$4��n��楛I�R����=n5J��0^�X��3�8�n\����*��ᐾ7�ʄ��P�r�|���&4E��ya�'�5��ɵ�֮�ٻϑo2�1D6�nw�[��@��/��ם�T���Y�B�c��3�ߊK/L+{5ͥk�ݼq��|)�Xa/Hm���+��X�m�nw��2��`�������W�5��������#�����K���iƘ]Q��YS�]g�ve����N�a�Y��`�5�f�R�©Q�v�Ӗb��k����g4���H�|rO_�m�N�1ם�)�������$l��;�B܍�������m(l5�ݙ��A㼦�7ڵV��H5ZT�N��{\;Wf����_pU����I ��6���K1l�D������ru;�w�S1 �,�G�7Uq�V�'����37�B��D�g����,�a�v�X�7x�^\��N�^����q�C[��i���U���K��ʼ�T�~��b�v�`]o&ˋ�c��
�T�_6��58��&�E�дcڄ���:��: u��S�cP����v_�~Ŋ�ʚk��sڝ���n^f�b����4օ�~<��V%�A�>��z��'�����Nk*����k�)�Ys;����m�����.:qM��j�>t�K
}]�ٽ�����/�����q�Tr�{�R���n��O9��E�u��f��!�2xXw��+��jok��{��v����Y�+�ݍ�Pb��iN�Y|+	:��m(��r\FJ�\��\bi�ا�sߟ��Ȟ��K��ˉ������-�KW��Md8�|�'�Aժ������oQ�[����d�U;��c��~��ҭ�֊�ۘ
�8u��ucAV�^��=�v���Q�V!����\ƪ��zP�NIQ�R�]p�ff�Oc�	�v���D4p���{�y��Ø�����u�_EM��}���C.d�^�Ѣu�,.��]��W�W�e3=������H��C��b+_,]�c�)�ne|�x�r��a�s�{Z�+�̗U	\J6�Zֹ���}�Q
_v��Ȟ����44��Y�n�3M�*��	P�Krf_z��D���9]Zv�z7W��5�.1ֵ��n���T#�%0ҳ&�Z�b�����sue'�wu�8�����z��������n�"�gǗh�=��	��o��J!�����<�j�p�uP��T>Q�	��bvL�z'�*���k���
�gI~��8�����#T�ڇ�y��1����m�� �.�W]+�K���1U��ՠ��F�麉.K}]�y]R�\��ު^l�~)M����h.:|��ROMj�9n�Gr��AW(���������n����P\vU�s�QG؇��r��,A'����J�U@�
�L�B߲��F�ՎX8���<+'j�Y�>���quı�2\a12��{�L[!�)W�ÔH�m�'�I}���w�NK�i3�o�0�֢��{���'�2v_
���?��^0p�=���nq����ILb�{�Ms��J�q�ʞ�oU>��{�[x;x��_Ү�g���ulXt�������o�R����!�,O�>w�M�m��,�����9����T�ݫ����6�K���t��:���^����C\��OvF�[��;7��3G^���u��d�u~�"v��A�j�����uP�r�Ɔmй��q]�s�l-���U���TJQ/�Y+�s�~��"�mW���6�#�+۰�mwS��������$w�Q��#��}���QW��7l�W6�=��^�޿�FS���9FK�Vx��C7�E�q��]�o�=�%_j麟,��{4+��݉�(��0��k[{���b}oak�%j��>̰���g�[Hu7��G��f�񶅐(.^��xl���&�}�ad� bV��؞����̺�����Ώ�N��s�e�r�C-p�N-y�o����X�Yoi�7����b`Jy��$^�p�"�Y ؞�{�/���M���5�'��V<��CF�߳[�����ʴ�%.�&�a��q��#���M�
�����i݊;itSE��uϞ=X*��i�\�K��SF�s�#���B��UH���=�յѾ�S<]���O���F,sO�|�#��0��-���gl{3�nڅ����D2�*�ae���)�]��mX%Q��y{;�3��S���˵mHUT�n\)��K���/-�����9.kuk۷�.�8�٨���N�;�k��]֞ѯ��|eAp���ӨSX'���d�/q4���^Nc�x�vTf�Z�wWϯ����Ё�u�5kL���V�]�ਯ�r�.>x�R�<�}ק}�c�h�Ԣ�U�U���.Yך���7>�wҳ�8���#M�kL=d��|wNdU3��;�ƙ�e��g�\��b�\4��֫�<���V���j�f��܆�8����]74��g��א{J����c��>��pN���_��F��)>|��p�[y�)���T	QFq�b|��4�8֥�P(�ՃDR/?>�5,f_Yu���^��XZ��j�oP�۪�©�`CN�5�gu�v�(�w�,��hND�%��F��f�N���Vq�&����#N3D�e�\8&$qj�7�=S�Ń��g=��ut��'N{��}��[:z������m;�]?+{<�J#[��/sxIr�&�?X���Y���tvA�P�խJ���R���
�1��l3X9wD�klVd
��Xa��F�<l-wave���vW�u��h�虌i�ѽA��9B"�n-�����Q��WMp2�2��M�ld6e��S���]Ux9�fm+7\u7q4��+���ʶv:�	�xѾw-m)y=������q��w	��o����P��K�4�*�y5�v1�]�uU�c�f3ޘ��
�T�Pڃ��|�����0��5�t���1j���W��V��:����g����A��C'��I�K2a#93�:����Qm�|�JŴ��m|��V���q��sI��o���\�-��y5�-{���z�߂�B��n�.���P�A���Vn��Rv���Ҭ�n���٩ �[�N�֤ wT8������R��������W���]γ����<��:�y�tsne���G"����u��(X�>��+��F���X[*oN�w?�U��!�=^��n��8����v��[g�M���8���O��̮��*B2q��H�o��A�g��z�˽�{_7km���`J��ڕ���qxz��	y���˲�E���J��Zi�ȇoi*���_�bS�SoqJ�`�v�Sܽ.v��'�\���Π�.7Sˇ��mmGMs;}Y�
�a���C�ݔ���_��t����-��T�*z�i[��5$Nt�ʨɪ�Ъ��0Byt��a��0���;)p�\�r��9�į*��Tٯ�U޽qx)�X����q.���q�J�G,�韂}ve����';h�	�X�s�Ǚ�5u���G\7�-؉���5�O��I�݇�vO�н	�E��y��[���rF�\�r�'J����n�U���\Kw{���O��K?d�5Q�ot��NR��Ov��{�����5�
�p�+����$��
y�oL�}2:=���v芝=M�!W����SR��u��]�V������Ӳ����M�}�86��*�쨮���(+���hO�F�AY��̌&9��tm@�*L�*;+-o&���@ˠ�d���w��]���3_,J<.0����Zoo$���f��Ʋ�J}Kq+퀅ˢ%����������\٫Q*�D��W�^b�zf/f�~{&�����Y[2!�=��&�m��*��)��E�lyW��/֭�J��:.&����T�e(*^#�ܸT+���u��e�W��#Ҟ�L�鍡���ue�\���Ƿ�!��}���v.a�F�b�Q�b��g}Q�Nj3��s���u)�?R�O[���}}5��5�v�./;�<�	Ց��͝!�,�6��u/;�E�_s�5;�o�趽��D�/��q�=���SǊh^
�����B��Y|�5N�˛ۇ���oh�s�-��S�u��_ѽ�bU�5*N�Qg�nIu�ք��0��N6�\R�AR ���6�m}n�\��F�D�1�M>K
�Y/�`�����ΆL�����i8{��s�n��J��T:;+��\7�FVEw̖aHU�%83 �Ջ��x�h��+�Ε�u[�2�qcCJ;��[�)KH�$J��s��v��H��k�͡KM�h�`Tv�Sr=�aY�bIō�v���u�JL�Y���XZ�q-a�|�P�Ӝ����e\�P���m:�zг��
[e>���b{y��Cm�*��.'Cǋ�V�Ow�Q��7���T�Q�_L+Y��z5�9�5飸{��}x�}�n�*��"=J3�͹��G���{}�,�'��r�ٍ���^r�f�5��*�Z����+����̳ip�z��H����?q���^����lD��������q�����î�賶.bO���7¹8�� �8�����|�f^X=��JW��ɒg]�6r�'��m�&�3�xseoJ[��p�P!Mu�(�4�\��D�Gs�ӱ�L��}ǉvjWI�O
�{o,A���e\�ã7&��X��Y�#�$�
g
��fC�8�C[ۂ�g:�t>U��N�Z��bVC�����S�Dzm��j�2m58����u�Eʔ�'{A�(p���D��r�n�,���m96��Yv�Z��k\�@���k�ī۱p&_FQ����͋/>3�.�`����\tk�����w|�3#�zA�w/�4B�;V�0��e�$�f�:��J��i��&=��BMgyk>��-u$�gX��<�X�}�σsQ]�|��ր��nd�u�Ci�W}t9�x�X�\���y�M�N�XX�^:GJ��p(�������q�Aӏs����
:�f�=ISͬ���̛�&
/41Z���up�
1J�y��F�^����Z����&��1=XT�/Tt��
ү�B�kZN�n9Q���WMJ���7S���V!�+{uj�s��*�G��9,1�wp�A�nu�y��K\u�*"�4�wK/��nݴ4Џ��Ɯ���(�>�6}u)���`��4���|�����u���p��,�X�8{����@�=C���0'���-��>�KIN�tqw�$ Yc{��e垛�O�,�,ݺ��wJ,��v�T���#�P�y� ��7��Aˁu��qw��.=�˕����ȩCu��R�� ��+ws���A���^�`#J9W̘���.�!\���;D^�wdc��",W�f"+n�K@��չ+�|��[���H4��ԃ1�M��d/�R�ճ̪,�yG��Âi�K>��� ���whZ3HT�RT>��s��g3��柢 ��oF-~{�w�D�4�`�&t����}8�&c�/Ꮡ��
� ���UZ����)Nl�LbCX��c��e�z�>�oKA=k,QE^/�
����f,���9K��ea�d �2*��NYsia���LmKNa���(���a�P7N=���I�6l�n5%�v4*jWql�tFL*ut�.='>�	�\�	����܀/�j����.��®e�4.�z�e"���Z���"5�a��밫H���x.�
��g���47���<�wW�1�:y�)ڜ+-�|O��;�\�]� �<��N��(䘐hE(�o:�ĭϏ7����%�r<G$�+�*J�ݻ�g�����*Y;�i��{�9��9䎻�*r�i.�!���(��1��Ǐ�"8��s4"4���գ�.��<<�R$D�9FDKQ:Va�f�gVs"�H�R��.��� ���9s�(Pҡѻ���b�V���3�����
yj�|��W����e�`UIY;����%��z��G<�DC�δ�=O*���EQG���Ww�E�B����^GP���R3�2�<���	$9�&�]#�rH���{�ܷp���M
$�#�������<�O(f*K*��jY�Az��B��Owp�uݕI�t�u,���$dDV%q�P.�h��ؙ!YF��;�'�I�8a�RYx�WrȺ�r+����z�g2�\���*Q%��%n���"˹��(EjJ���U�����&�b�y�e^���� S/��x�{���)�^��zB{�x��E�7�� ��iR����x!<��è��r��6MÕ>�c=���͝k/����̥��^�n��ut&�F8֯d�:J�.m�����:���<^X��=��K�-˱��w����N�o8+q|�ٽ��s����G��=r����ĥQ1}�����,')w;<ո�;�P�ش�EΡ�.��n��]d�舮YT��[�X���W?w2��v�QM�5�w\S��M�����i�F��<k{<%���<��o��\��O���S��Y`���b�v�$q�j�=P�n�׮�sё�ZR�+��>�%�"�������8��.��%-ݫ�!�C�k����˃�=��γޞ�J
p;����ZY��c@��mF����k��i+��ܦkK�:�8���O�q߯����}�1��ԣ�4;�˟WK��kW�������Y]�WמI_��(�s�Q��|�utǑ}�97�'w�K3��]��p��v�6�����U�w ���ໄl8���ܠY�WWJ���Ȉ����~�Z�����e�����9G���-�aP�{�����6X�@(ڗ=�vvZ ���w���y�4_*:'��j��D�<M�@e3�3o97x�>:��_?͘�tW<��m�d�Q������Nw�n�����<�*�y�;OVn�X��:���~�Y�6[�Ρ��v���e:T-:���=��q�.����i�c��
v,/����v�u�Q�>�E�j/BWz��5��;�%���>vzZ��vޭ�;���5����2_�9ıuD}&T~������;��tϸ�������F��br�+fLs���I@P2�?��u@�YRLz��wڕF�O��y�pI��a^�8��u�1����2��5P#���R��v���_wn�<S�*��(̹�Ki�Ԡ���ci�*�v'�R�:�vύz��A��w]�!sJ�&�9z9�ky��ک��Lӗ����l�^sT}~�V�c�o��s�ȡ��6�u���]BLU6���W��i���|�7�iB���R��d�le�Պ�����){� �qW2��Z�뭢���l>Zr���Y�ҹ�-dW//y�YL�_]�(&	�x�?%2���0�֑n���}�k[�E9��g��|���J.�=K�vN���8U,��������x���HY���M�ڄS��������m���7�n��o7n���W�1�6�vZq�C���:���0;��܊�PS/��_Bp6����⺋z��r�=:�+�C�.U�3|�w�HX�����Byơ�m�݆�*(�+��YW�~B����\���%��`�|nO	]��d;��&׸��6�r��c�[���7���o<oz�v�k�Зqy�G6&�{��u�K������?d����}.�KZB��5K3�{#�Pv:}�!�י��W���Q����l�R��o�y��=gmE(��Q�I�;7\D
e2��B��w����?g�ǽ��԰ʌ���1�W�C�ֆ�p�;0�7��C� p6j	���*ԯY��4^{�<ǥ"Mgz.ϣ(Ei��﹄t����oQ=��xr����Cr �]�n�7�����4B�Ϫ+�B��X[u�D�ZZ�Y��*�NmAo���B]^�ܽ��-e`72`�����s��Ij�=�T�>��LǗ�-��0��FE*d/V�:µ��̮���lv�fj�*=	�w0�6�u��*}y��ܕՇ.��"��U��]�*k+�Y9I|��,����W�w"����%�i�6`�vT��.|�{E.�{7��WB����|b�}�8���kؕ�\:���A����F~�!�n���xO�Y10��_��ҋ��6x���>�'�Ө������)/ZϽT���/�*%z��z�2ٟI�a����k(�:���!����i�D�G�򸘘��h�}����VK�^!�G�zT�����m�Tu�Z%��L�n���lM�>���H��#�urw>��t�������+��:�������v\&�����U0�P�����`�*<Ĕr��^�͏i�ݨw��7��3[P�p�g�mUG�r*�sihK
Es�檏���5���=���!%��� ��N�q���v�v�y`vȦ�ܷ�=�}�-W�������N��ݻq^�Q��+��JvX����[N�v���G;���Da^!�̷�5���i��g��?W������v��碻��н�����yGV�|4��*�ed֖/&u�r�����E��^G�s�}��χ{=r����[ �ؠT��wk���!���b�Y��Z��~[�~�%�uv^ p�cj`��k*�d�Y���J][[�Vi{��a�1�r'}#�ycݷwfQ����Y4zT�~��{;��k{%�z��8��-Kq�ܾu���Э@�c��)�E�=�U�WL\dγdςy�S�mz��>�'~�[Y��ez5��E\��46��-�C�Dy	C��H�D�I�`ew��L�d���wׯ��hϝud)���|wJg��{/Å��ld)�,�}�P��l�`e7p*���tZ�ǻ�x*�Gw���>�$�+>��l�x��=�|W�=t*�][/>��[U#�^�fU���7�w��ٔ���J�϶|D<W®��c>�B�g7�4������Ic#f%��+r�z� ͏{2-�����3�}�� �W�dl�*��Ы�v�Xߏ��s�<]]A��{)�F���G���i��7����O��@h�w�X�Ct��ȟ*�>�`���dƹ�h�׃�*�07�wfA~�n��숙��Ӵw�/ǻ��\�+��^x�*�^vʝ�&��y<���W{,� ����ՠq�@W�f��3����c�6�u~��_iz}DEG�I�~�h>�>�>ݳQ��T��y�G%�`�@x(��9�/r����ۄ�߿�9�7P?�m 'A�E<Ya�gq�P� 0��hg�]���ڠ��-�sx֮M֠7+�1i�;]�k�wB҆�܂9+���6_v�Tj:uu��Z��&���L��!�͔��V��$�q�<���om��#zZwWN��A\�����wp��uG���T��zykA}��������)�;��i9�]����}"���N�Ө�g�i�?%~����[쁑�NT��hV��gL:�z��R�7D�?Nu�L�~H~�yp3X��#K}ŋ͚�F�}u0&�^2�ϸ��yW�'Mz� ���nm�^b���V��i��I�:�a�،��w��7�w�#�s�2nz��2W�I���.W R�r��T������Z)�%��zn��Wp���M�}3�����~Vnk8����?%��9�����Gq��y���P��
vf��X޸s&YEz�ޞ������M:���L�S�w����.�����v=��7�\n}�l����x�ت\�ێ�D���D�t�F??�
5�Q^<��ږ?_��d#>gF}��]�=�P�n�Q����w��?w�Z3�r��5Z}T��uR:�g�(�¼^�к�w��A�y���'��F�} ���'�4�B�|f��.���3=g%����!��z۪��D�RÄ�}��S�Hи�^�����ӛ/�x	�=q��v�_�ӷ7��&x=n�xx���ӓP�Op=� 6b�m�M�o�u���������vG��W�׺׺)o6Yuw��b�Z���.�T�7�2�Mq�G�A�>�����,�{'A,��&���"U�f,�;}�I��,�P�/��u����n�\{��p��* �ٸ�S@>�Y�%���&��}����liڋ\=�o�^U��ߜ�*�����e�ne����L�TD�N{N�p�'���^��i�;���c�������ND���tۺ��r*j=�tƻQ��Ln8�o}�V�[^#���dj:��,eBՓ��9זLg�ޡ=6��������F��z;��\w�c26!���c��v����8���������Ud��G�=�"v|��k�U�Ú��y��Z�~ �}��7��=Q���ͯq��O5L0���uG���y��l�o���n�tUwl�	Z`U��l��8�V�����W��,ml��F\t�{&iT��p��\�.��ޭ�G~�<kݝt/��Z<�O�P����c.2��\d�\�痭3n�Ef�U֬3}]^�O�T����[��u�~��%Ҩ΅�GI���=UHz���;T�ǣl����{��G��{�ɟ9��!zo��m���7�{i��;��>������(�=�%��x�Vj掓��_�&|�����i�y��j����g덆��N�������1ܳy����sH�;��b���T�Z��ȺXt�
��.8P��㪗��2Y]����m[Y�8�e��Q�H�nMGWZ'8��6�m�9��б�����ퟬ���Q~��-,�i~��̆�*����x�x��z�dzt|��-o�9�f~T�"���
_������⩁G�>�Je��B���|XϺ_�FDo�_uמ���[��Z3��8�=!\�pc�)��;މ�Jm�5�7@U�^.�6��Q=����Կ:Ħ�,��<�^�G����w�W�[޾=>�UYe����% ��Q��� v#%��T:c7;[���X�]��>�޸��z�9�HE3�o�tT_�܁{��]ƙ�<��Ԫ�~�X��Oz{��\�W\߲��Ai̍�^7�F�����>��Q��>zn�\9�$
��>e��3<��v��(׶�F7Kw���ﲸ��s���.V�ρc)/ZȏU+��A����O� +��˃�Ӿ�HI/���U��0�j�+�ڵ��z'�=�M�-��MVѿ�χvD	c*5+�,d?Mx��ʇ�3#��5��X>��^����#*�G/a6�ɟ#�1׶U��^���/�>������f������J^}=ȕ�7��z��x�����{��fǴ�n�<�����a����VW~�N ]050����Ӎ��j�A�UhC��6��2� 3ul�-ý�M;m.x���a6,��0�%�����#e�nz^'e�&�0�ǪƼ<�v�,���U���Էn�^��T��V����ZS�������Yw�P�d�p<��އ�ћ�leyݖFDzX:k�wq��V��IG.}@-7;,e�z�9���w�o��8l�Α��>�<L�q�j�G�3� (�u(�{�n*���:P�����7z���O�����ث2�{'´�#==��F'�O�Ӡ���ZG#ت'��x���;)$��Ĕ�j�
�>����^U!��Z|0���r���ی�l�p�ב���\;xW���՗�ّ�%+��P�	����F.=�)��'0�����b�b�&u����O#�юk��&�����{.}3U7�i�J ^�vW�_��1�}�H'�%�;�MCk�p��o�ax�Y�Cw|$`��略=��Ou�9)���8Z�W�r�=�H��e �n����^�����9��ʽ7S�dwyy\{�6s}#Ǹ��_Mz��,�d�D��K�xU��'�y��z{	y<��l��5��)?W�c�;���20�W��<��'�3�3 y�([�O����Z}
oꮢ�U���x�l�*x�
�u]�{�H���G�h���~�v�KAӍ|�dZ���V�(�kNo�^\/U������w� U�d��Y�^���]�H5�է��{t7*a`u���u6���`=\�90l��{QN�P��w>��^h�;��7�m��^���ħ�G�挶7��K�N�F�;�;��0=��F'̈lER&&�W��-�,{�n�>�����oFd۷t�o�0�y����X��"~�^7�Ks���𘘧մoK���0��=�|�=���Y�g}����y͚G�΀��.� �#���߮Q9U��csd����<���U�*s5~�6��kOQ�yO��������7�~�)�U���ZM�ωyF|&��:myT7u����kw�_��LMl�i���ǫ�fCϹ�L{�L���p{��l�{�%�������ᚫ�_��W��s��~����?,wZn5ρ��}Ig�<���}+��-�:w�߮T����T�p�%�f=�E{�}'ۉڏe�W���g�7�,�Ul�|���MQӾ��I��騿���������ܾ-v��q碻�D�FYP����߳��u�1�uH�ޤ��ތ�q�ݥt�*�]���վ)s���:CEǚ�hn�t�=7P�}�����k͙ﺺX�O�+wFi\�L��k�l	��2���~�i�t����+��E{�q����flp=qT�_|�>�+�0��Oe�͚���q���}
�I�=�*�]��{WK 2mH�+�2��fW:����*a��E3�s.�Ŗu��r�]���%��\��e�#gm]��:�z����3B��y�ݦM��Uw(;�f�qȳ��,&mE�`����?Q���H���y�0k�Q��"t��-�|D��H�k��<��ey��;�7�|�w&�3���Naj�mWH+Ґ�&h[�7N�A�vh��޾�c{[�;a�/C���-�$���2��Om� �_z?3�da���|������=�>kZ<,b�!ydb���jK5���I��2�Z����.B�����(rt
XU!�#O�w�T�/оuA0��
�V�;L���p�q?К������X�J�e�e	��`��P=B>f���}�2_u�w0)3�ع��Y���L�t_%4l����6m~���s��-���wG�}�	���4P��HT�k���I0$js�,��4i\ -Hm��T�qC����lu�:<q�vVˤ�ӧ�鮗���Ǭ��WΣ+�2�I3$�3N���S��c=�|;R2��i;�����̾�[�	i�PƖ���$㤕���7uk�l��m����-A'+p��>�)vOt�	*��b�,��;7J20�5�r	1���u��%��/6'9� ��j{З�������,^���2��L���32g%�c�x�;��t���R�9�8aT\ҵ���K�"Վ�F<|;�cKiA��A�ӯ�I�{L_Xl˹oے�l��Ĉfe)�ʹ��᝔uC���j�/1�A���[F��U6�5� ��;��d<4&Q�Օ*f )�N`b��U���tǃd�3�B�w�ֶ��ը]%���@��2�s�w��B�%���Y��C1|�̠��F�T�y���Ცkwn���Ã��8��Y�TBap�H��8^衉�V�:FN������v��D<�(n�UAS4K^�{.����s��]mv']��&��<pЙ�Y�MI���d=6i������E�aՆ��ݡ.ĝѮ���=�y��׷�g�=�i���Y�S�7�޴��|.�P��	�y`!U��soaL��5���<t/���p޹�c�)�ܩ�>6�c��nyN �=�L#��35���4_*���o&V��+n�ź�ln&Cy%���w{�-�6�����m�A�z�w��� �3�e�d��b�5�:޴�eo1&sƨ�A�2���qSn7�<�՚gb��lA���J�{h��"څ\��ཧr��A-���I�K��hv_vȞ��E���c�^��T�Jָ&Ի�@9���#�����`�13�Ȇ��^4� Ip���k� W7�������b��	��,L����%����oƎ�ٮ����������P��;65����jɯi]��u���r9����nꇣ����xx��W�8���bt�D�4�'D7\\Oi��t�7e�Jҷ��ʒ�H���J)�m4P$���m5�,(���#��T��嫻��wCq�t�]GGt�:UW�4�Ge�]wELӒ�)��y��rN��n�w-�by�5<<�5̩V�E����ĊSjj(��E��uq��/D�L� ԓwOfĄ�½u4�N��J�/s�LO(���wr�Cq�tP���W�v�O7E�nN�J��B�I&H��TAI�7w#�4P�r��*�.�Jd^螫<��u���J��������rLD�3�L��t�OR��3�.�'��E�J-G=�	KC*����QzZ�ryx�ywny9WrY�G2�B�Q����H�Z���&i��QI%E[���k	w�T���QQ%gY s�\�2Y<�G��x�wL���zr�S��,TTAIĺP�"gh�x�$�i��r;����TtZ-��,K$6�B��9�m�0�Nm9[YQX���hj��!�Ǖy&h�ȫwV,]Y��h@TX����N���I����*��ڜ�YǗ�d�
�ͤ%�U����
@�v�eK=Yz�f]3i[�f�SX��0��Z@S(�'g�9��ϰ���]�m_Tj�(�����.&Gc�|�}~ݻ�Y��|�EW5>DU�G��<��hy�p-�:�9��>�:�\{$}��-e�\4׺u����ߋ0��qJ��R۪�ꈙl�o
�{���x�hXQΘ��O3���(��WO.W����Y��!�-�����ϥz�>��S�H���O$���ѧ}	J#]��wW�y�E��H��ơ8�#�n	=��S@>�Y�Z;���ˤ�*accN^���t�6?Sn��~���t��*�޿ z聱�+��>/�L�TFo��ޜ��8)�O��K��Q�݆�4s�Xjb����GӬ�NK�{�@l[���9UP��۵S�?O��Q1��/P]o9{�3��Qs�25��o@,bTj�^71~�;s�r� >��J#=zT6K�>���p��)������d�t��\�3�Ƿ�Y,\s��yȝ�����4M�{��v����Hy聹dP��7>�#�=Q��L;�6������m0�~�vW������$�Ź��t͙W�]p�N�c�}�9ܼ[w�?
���
��q��/�UtO�'b�K�h�ui.a4�ɬv	�}+;g&� ����wD�ϧd�Ƭb;!�v�'��5�`q*+g�y���a!膾�#̥����mE�u.�NH��[���5d}`G�v���tvuՏƈ��9=o�ق�G�kE�z$�ˉ�v�j�uC͙ñ����/O����g��]�l�K�^��ol��<Y��<j=��B��Eh���<{"'�i:X����Q�y�ſO�o'���������m}��
�X�<z�޸Hߞ+��v���I㣧'�Q�H�ႺhՎ�w��5������ɝs�B��q����s�O���8�G����ym�n`L�t��?e{=�'�Ni�NN늮ny��&u�ɟ"�̆�O�t?9�;뗧n�Ԧ��Q��[t��Һ5��}��oPf9�L��7�M�0&*y/�2�mT/Y�|X��~����kΫǨ�q)s
��a�Gz�:�R_�p;���\��Y�P�SrZ���_=�p�O�-�w�r���j�d��B�F�8�6s��O�w�������1NQe�i���(�Q����qMlϮ�#����ž�m���^7��u�RGޙ<u�x�_�G�r|�� 6D�^�N��k�~Q��#���fv��z��*{Nd�i̍�x�<J�u��>>��Q������*-�9 m�_�ߢo�S�;�*�=S���.5w���
wE'C�;�f���E�4�蟕�k�v.���uҙ�;'f㧽�q�)l=�ȕ&��x<
nT���mH/N�D������u�'%,D��4tD**�w�]��	��3�H-��,�9:&�����+Jz�O>W���++���{'��?JӸ�Q�z��Ǫ���������h*������~��8��~���l�(-���}y^&&)��7�|;�KIU�b��_�8ws��3�c]xv�tjp�O���vp�������蛨{��a�z�MF���q��K�7�RO�x���T���y�E�D?z���u!��{�;��_��a��y�P�g�zFC���h^��i3�	G��lg:��/�u1<o�{n���yGǐ��H�N��Y��ݢ���$����o�Z�p�4�>���)W�<ۚ�3�W��{��ʎ���I=�y���z��&��쓽ض^�.t_�kJ��
�o�o��61<�K+���w�z�7���g��
��fL��Y�jqP��F=ݢ�Ĳ,�����&��q�;�z�vz�{r:�$S�^�ⷽ�~���./F����7�չ�9<�fۢ[7V�Uƣ��:��ςy���<�0�tU�u�x��B��7ק�μ�z��T:�CFG���O�K�&�Sq5
�T=��f*Y糑��E�{�tx]��%Pp�>����x����ܓ ��BXHjk��s������A��ۺ��]��N"�^�f���\�����c��6�+�>�1gL㹘XMq�ħS�y�)�4��9�I�3��a�O�9�E)���';uF+-\�MX�XY/����eǳ������2��^k�
p��=o�E0x��Q`f����ͨ����j�Ie��=����e��"וG�>��}����s}/���^
r�/4�������X���wk�����R6�i�p�y�Q,*x��'�lÈ�x;^;wM��C��鋟15;��@�d��f%#f
n��x�!��o�P�Zp�����s�������������g�����2�O�B��'��(=��LLS������w =M�G�ݖ��őX*����>U�$O��;��R~��n�E[��p��S�2�__�����7���4}ԙ��򾚽��x}���S��k�Ͻ@{�� 
߲�5�eq5^p�6�6�}+;G��s��/ks�߶M��Q��|���[^��q�:���.����5�>.w>��Ɨ�צj".{jr:�����U�ד�Οi2v4���[�S�>��q:Ͻ3���yF�@f��mߞ�s����G��M�p�;����ی����'Ei��?���i�0��#Ü��*R�E����G �dc��+53��f�6{x�Tu^m^\ ��é^&+������>�1E�{2���l�C�x�.��=���<�� I��)Q�vgs
Ze	����f�æo�P����1Un�{�����w6D��g�x����<՜ǐ����s���z�Ѕ{���rӳ�+�X�3�u��Z�d�)��x��ϥs"5{Y>�:a_:C���V���Ew�}#���xk쭨w�z���5����t^��z����w3�>�O���=�ւ�<�8g��B���g�&pa鸊(z��w�����>�Q�iw�ϧӵ>�Ҡ6x��k��9�T�|��q�o��~���^{w�F��\�qeY�!��* �b�́w��g�b�]/���w]{N|�/�#�>ҡի��{e��cvj�}�Y�d{7*�m�^�Q>p� fL���EE�E���,z�������Q�r����SG.�OW���r|RPV����}�w��z%Ѩ= %2G�&[(�¼^��L*y��B�{��W�.u��/޸&�&����$4����}�DmC��#�"���2��T�U!
���Xr ���>��i���R�,�9ܠn���m��__�wӴ�y���#},�z��9�@of�Я����'ϑ٘�t����zw�����ϼ�Ewκ��}����޽ ;�e�ne��GŢ`xf{�C�wb�Ί��&c�a�'��ÿ��q��F������=�slKw��'5D��tF�ܼ���Q�$Y���⦿W��]{�
�.dw�>�;��+��B�}�v��c`�gf�v8���h ���}��'J�b�{�b�}��0e�I��s&#i'F>7�_��u~��=�B^�y]���W3�;��ߕ?W��2x���b�����{1b7�[�Z{�M�y�C���EF�wǲxi+5�񩎈��)ȗ9Ю�Џ�ϓ3����:r��c!H^xﻩ��]O�웨��V�w���j5΃7�ǹM�s�����RwݱO|�>kg�\�>��c�����@�;>�#Ǧ=�[��׸�Gzx��`�����ɜC��Mr����F�Q��rw��<�N��I�>����C�y�w�ZZ؞��)߅���#9�}^�.}
�oV{ �Ns��,׻:�{�'ǽٜ��e����H�ȿc�l���Y�C+���6�f�J}<=/� �c����z�#y⸫�m�7��x�D�g:��qX���ӱ��ϰ�U!�5��L꘿��No�3�ׯ�ߟY�\wǸ���l9qu�2%G�[�I�k(�#�t��NN��Sn{ŋɝf�gȼ�T�:}�>~u�{�x�����WNz�{m%��s[Q��1ޏtU3rm7T���D�M��jaz��>,*w(�S��a��BZ���2vx
�bCq:u����LV�tk���"�y}��{cdt1��br��B�@��e�&Օ�t�g��^���Z7Nv�e�j��U��(�.�Ce�Ҟ^r�F�g��7��T�Go� �3�gWaYc�m�Tfnٍ̲{�eǵ�7F�^�����wH1jx;��z��o�Pn&�����
�+��z�!��TWn�]�]e�1����{�ǲ zR7�|;�5����\��.�4�n@�N��/L�ʙmz���ۙW�ђ�{�E<J�z�9�S;�8:�n�_�U�/A�v�Ϊ�Ph�1>[�X���ǽ]T*�g x,7�l�O[Ȭt��|��zF�q��#r5�nD�^�;\��)�W�H��VLL=�VE3�84�V����Kև���R�Lg�}��2g4����<�f���07�ݙ��4�q�Z=�7P��+���MVѽs�=�����yE�QԦ��EE7����>fx����)�	ٸ�@z�z� ��`�Uyɺ����a秤��^�W�O=�pK>��I#G�lS�TY����ȿ/_G���_ު�]�l{M��C�G{����ED�om���)D�g�y�5�ƛ̿Iݟ�ʘH�{�wp�5�$��>�����J�3��]�����܂֮������;[7�3�n8�-W�=��o��)�7�ۊ�{l�_}k��T�N=5}���[��ˢҗ�/����.�<#Si�n�)�9?����asJp�h�:s=Μ>����PW�2�=}f�u\��e��c�t�Lf�ס�_�>L3T�cw�xyy���;Lc��;��׻�r ���Q��bf��b��:؊:-ut�8��M$wr9b��@k�}��� 	�c�k�Ef�댟
�q�F�n"zX����_�����#rM/EP^��VV׈\B�Gz#��#�=���0��U1��Mib�g|u�1��Q�m�.���f�������S�
@Z+�vW��;<��1otSg"N�0�w�3��dςy�(�9ڛ���������O_������χ�=��C�~�	C�ȕ=&�SqP��������>�>�&�#]�״}T}2�G'��#��i��s�=����Z�2�y�H����gzw�%E�y�X-3���� {�s�s�٠Ѷ��=�����/���O��J�x_ʫ,����}^*�=&zg;�/Ū|�;fH���&�G0��x��Z~��gzs9�~�x?�a��G������B��^�K`��h��޲��[�/W�MZ/��"E���������h����g����@s�7q�ܳP�<b|͘,=��D�>�a�Z;�X�B������Rn�A�+'s5N�{Y���C��V�e0V}�^��3ِE[��*��� <5�c�)�m���
����R�+�r�kx�J�CV�F>��fh=�Yց�5rk{k�L$�b�P�|��vfEZLg(E��:3��g���9E���z���޺5���Y�E�lk�[ᔵ�ij�9ӕ#�T䭛��:s���o������)���@{�]`_��X���nQ9>� ͆;�u��Sv�c�j��eu����U�kJ���G��+5��͛�y�G%�`��I�>%��T��~��ºS��7�^E�mhw�N�5�ƙ���k�e�ϫ����G�I�^�S�/�z}s�u���x��{��?��x���7�������f��	W�<9�z�t%RA��J�N���2��{
�ȏT��dЯDw�Θ���	�7>����Cˌ�qb�f�޹}q����tֱҜ�|�21��yQsr�������Q��Z.<�WqȟHë*�ᬭ�w�z�Ϸ�$����w���bw^���!�������v��h/;�4w�墐{�Y�lY�袇�8�똨���sr{���j�����8⣦X�k��9�~/��q�mW���d�+!�OW���T�z<��+�;}�k:�_{^��o�p�&S������'V&����x���^�Uj�M�b��=\��ձUW�Ӓ�g�9��+��%Hn��1SȊ��-��jX�Ǘ�b3�to����O�w<�� �����n�J ��n���m��x�Q'H�E�5���]�As�E���ɕ�]XB��֍��m�7�EI��	:R�˭�P9�x����'����
Ji�s))��3FcU���.z��eΜQv�te��Sz�w�u����u+tj�#ҏ���y��ok�vn
��UH�D�e�y�-����csې�K8��ijJk�=;O�lz@Ɉ~�dxg�Ӭ�{>�!��%@{qU!
��Xs�Z>�{�=\n�hQ����z�7w8P��:H��(��X+����.=����9 y3�@Ǭ16�@ٌ���5�Z���g��ws�Ŵ�+�N�zϞ��� ?)#~�T��Q��.���t_Ll+����T�z=�}�DS=�7�3�@vu/
�\{��� �u�Iϥ� ���3n�gl��7O��3�]�?�u��ڏ�&:#�r�Ȩ�;��e�]F��m�_����gh�ݨ�Y��]��]aX@�@�q����7S�(��͌���'ä�k�ki�Tr�%�25�^�~����4W��f����?M�;�� %a>>Gzz��q��a�m{��zx��s*CA�Nfr��pپ���=��/e�W���C>x's�T��m��ڇ��3�P�{޸ܿ�T�V�j��A.���Ͼ�� &-[�/��|Qߣ�����B���Z/�=�ǳ���f>��&���|i31���l�n]t�o�L��iY�hd��h��;��ӻ��e򙑜ɍ��.����9�Ǯw7Q>�f<��3�'A��Yu�1���3�����Zf�";z�u#�P��N%�9+��5p��>=�X[��w���=�����Xr����bk��Y��%�)�T�n�L�Z���;G��\�n��vE�\}�{b����I;��Y�f�-�)�x|n<�
ٰ�c�U�1��ow�T��n �����iPg���v�)A tӋ��ޖ8D�	w�f�����h��W���ؤ�[ƴZm;v|,��;�r�4y�98��I�֨+{���Gv���<&i��x�u�@��I�҅^}�H&��W�R��y�A=J��7�8d����,q�hus�ާ�µ��ƕ�A�층TW�&6��n���١����xA����9�r)`��P��3zv�qM�������F�̼LD���:��б����IN{��v�.�t��ɋ��,�x��%��i���vSX4�܂� �e��,Iǝ훮�(
XGR����wR��!�N�t�����5	��������[5��1��e&�A���%�:�m��^��XAo�'Z:�7a��2���R��r�����.�tȭ�u����U�tR�;��TĢ����KU��v�R�KfW8:�Kwۜ���.�&�4����G}Э�Y+��T��8;o�[׬�#@p|��.��J�G��c�w�t�GY���p��{h�V�Cw�鷺�l%�0�(�k>�u�fl�q�w՞j��n��dD�;&�����=A�4���S�,-��>�ڙ׫⟜\JǤqVd_Y�<��lO�T�m&���.��J�F��Mʺ��s^�����G;�#���$M�iMBAf�X��ic.��M��ĭ�5۬�]���V�ⱔRMd��MJ֎"a�Y���5�gC{t+�}��E��0[�2�h�hx���;v�
)�x���CL|6�~����ۡ�\�m[��$,���iZs\ċ�������������������(��Gn�Fa�߼�.�;eૣ���<7.H���Ε+WI�1�^3{v�4�n���.͐�9\�����OeL�y�-a��"�{�X�F*�IK���D�f�.�T�`!���e@���*7Jlt@��eZ�W�nU�ٲ�Q���ET|xL�j�6����%v���v�e�/����t㒤z1-��kC�v�!ʆ�*˩[H&E��R��>�H��ڶ-f���0��F�?��C i2��a�	�
���]�k�I�K�3u͝����s9q�iD��2��,�G��wF�2F��w�lU�5�5�(X�P����Q(̒��DAZa�HQփ�H�f��P�%dkEi!	KV��Ia�2H��ЏC�BE#(�+%KKK/�ܒ"NԕV���rK#���UHY�A�SL�i�zx�C�fJ�aX�*4B$29��ǝ�����&UJ"��BJ�VeH��"�Z��Ydt(��(�$ʣ�E��1ZE�du�E-@԰蒚j��Z�Vꘊ�Ҫ��Я��nd�E�j�\�D'M�(R����!2�\Q(�U���Ұ�u�%>q�ԺJ���E��]hV����BZ*d.N���YJJ�^�3#T��R$�"���.�aal��!jJX�T�:D�.jj�Ⱥ;�Ii�R�O�Z�RR�%,aAM[	^��i�~�坵vB����@ح�'�6򷒦��J����Ga���{5�嶹��uw]�}�>��k�;�#�F��͝�?�^K��R�����|}j3���]g�R��)��aDo
Uz՗��k1dfNN�Aa�>ܙ�L_��'7��k��o�O�q����W>w2Q�{m�a�n������7�%��98]Sn{Ō'Y��/"9�c��:i���4��6�Ϲ4������n��vyQ���R7&�SqT���y+���^F�B��f�yo(z;o�N�㾓�G������D�=��W��ή�c�w��\��Y�P�M7@u�h�5�ʚ�?Zຏ���mG#Q{�Y���A�Z��X=��x)����% ���*}~�<��U�z���=��>�;Հ�2y���x��\C�ZG#ސ�g}z�Hq�UzK��Nw�*�h(r:ט��|`�;E:�hނ�Ӛ_�x��_;Y�'8�o�zG���W�eJ���	�ݕ�@�!>g�&&�E�&i�x��>��rc)/ZȏU+��y�:f�53�}U����E�ɟ};8Z�d�s^�ʉh�}7P��+���5[GY�݂ş�$�2����1�'<�e�� � ���z�[�[wÚKi�ko .�w��{��i�����JNZ�V��*��8j+����`8F�9�Q��D��m�!X���hh�[�cJ��ق�euj�81E �uN=o �z�솓��E�^�;9�"΍����J��s7s#Oyۜ%%��_�M�G���' �@�\�^4�誯#���ךƅzU/�0w�	I�V�ن�6��S�=^��4W���uG���@yg���đ��$�����g�l{L�x��y�4��;��R���>�f�j�Cy��s�>"���������.sǐ��P��QU렷j~[���π�%�/ثC�������Ǻf��b�ǘ9���:_�vⶲ};[<6�Ezs�_�LJ��l�>ݒO����c0Ε�>�Y��,�O ,�_�A�Y7��I~�����zC�oO��:�v��碻�O�aՕLeFMib�g|o\����{}�޳�k.+�+~��|sgЧ��Y#�KGh��G����ym�b�{��9s	�~;����x�y���)ܷY]�?`{���P��/_��{�y�ߣ�^q���>�9D>�Nn$��75y���,WmOf~y:�g��+��n2e�<���OK��v>�I}=�����*�F����}{�Ꜭ�W��������<oT����2/��Џ���#�t���W��G;W�!������ҁ:����J���g�]�>^��^x]h��V�{���WraO��E�{r�Q��k�Pqg#\�'�lb���&iͤ�@�o-;��)�8��A&�4��NN�����jr�Cb�����SǷ�c�wwR�+������^,߾� 6l�m�Hu��h��c���a�up��H�9[�U�_�M�l��ؤd}�n��:}%��������۪Th���Ar�s#g�<T�(�ǉ����x���NR�����^.s} k��=�[�jx����0P{uH����{N���{^���mO)��w�o��؃�5EG��U�=��z��{�\
���L��߁�ɹ��}��so�'����CXs�GGw�&���x\G���G���l�w@z"���f|����"��W�U	�>������ލTG�-Vɯ��>�q�鯒�P�5�d��~�<m̱���ڔt�0,��7��QV��M?E�h�97,m�mhw;�5�ƙ��K�Y����s��8��Mn~(����T9*s�Kl�����\Z>����'���z���wO�'Ei��?���U����bcrb�x�vO��%���T���V&�ʎ���dWq"�͝�yy^����5�Y=�{��3 ɋ(�^���[��y�ݫ�����D� ��-
����Wq��:�*���ڇ���$���Kq��@�wX8b)���`.�EX��7:Pd-F,N�=˻#wihV�bಉ�Kw*76�d�|h90j���}J���-�8v�k��^V.�z�٩��oh�(#;`���nL���CG;��u�z?S�|hM��΀�s~/�����.�������X��g��W�T�˺[�O�<rs9�{Sq�{�+۷q�3�o����cn��N}���c�q�m{��-������qPW�>��ux��F�	@��_��|�=d�s3��ȎsA���|�i~���ˣǸzsΐ��+΄�-�:�V<U��
f��L
<�˟"��ږ=~^�=�ϙ��^����|���!:8��f�Gt�7�\{!��vDk�vB ,ت��l�c�SQ���|s�������U�[��̌�J��EGw;c#���+zwMC�������Cr�P�UHB�z�4�Ч��;�9}	e<U����U�H�s�H�{�������~�x�<�L�9����t��_����md�j��P�AJ����@���Ci\Uî�x����<�� �F�`���9#!��H~'�<�=V�h�Gx�"`���D�)�;��wN��W�ǽ�>>��s��r"VP�{�ї���ΰ5g�r����i"�T4w&鍿��G�.V��wǰ2�J�ö��qf�>�?���~K%fs8ܡW8U�`#�ι�N�h�>�*�>�ŕ�;���F����91�51�b��S�Qy�N(0�ƾyVy]�l���ï����ZL��	�(���\-�k�a:�q�����hP���k���Ǟ�	?=X��{С�]������F�)�Jէ�����U�9��y�/���z�
��%Q�>GML<Y[��O�I��:�m1�گg�s�rcٕ�=�g��'�uq�F9�9�>��"�������{'�=���a�f׸�ɍ��ٗU��6wG�V�A�� 5N��:��/�NO_��݊����}��.'���v����6x��(�g�Dl�)��?T��o�-�� ؼX�������Mgz�\C���~{G�JK������{Wݒw��p������+n�O�����>����
X�<z��z�#�j���OT.�#��ۉ�.Q*�<����|rrp���=Y5��;��!9��#�q{<���~-1F���/z��j�_F\�a��z}��w9QF��K%��98\U0&�X���o&|�ϣ�Pt�+W���|�8�Õ�=�tz;�y�؏e{��U��m�Y�f�M��⩁G�>�JgZ����-�'�|*�����+}��v1#'��ў���o��Q��*��_�}���x�À�k.�]^e����{|�'Yu��F����ϩ���q�􁃾����
r�/#L���u���2.hxj���ۋYZ8�F2U�=�hB�����m&]&��F�c4]f���\��x@���l(��I��p:�~��,g���Kz �z���c����|����v=��kk�nٟ]N9������g��7�f,��&J]W�м��QK]ޠ;�A���d�nmCE�U��i�E3���~���H}�H��.TUJ~�@���7�2F���R�\����4����]~�ȃ��%~sGk�"v����Vt�;w,3ބ�Ȩ�U9 /�Dv�"f)�x�+@b��\=�K�{����ε;˗�dǎ��zggӠ;�+�5�U̐���C댯MV��|7o����q�]�&����<F�v�N��/U����9.p\@��j<�)qU^Grn���n�{�0y�w/��9(W^�6=^�:��p�K�O���w�-]��ߏ�l�w%�ςܫ�^ڝ��á���Q�k�Z{����cڏ_ٵ�7�q3Q�Ż���uG�_��bx�{�Q��=�������xz��}�:,x��DJ�;I���F:����ٸ�Ǻf����������Y9|�W��ݭ�CR��Gv��G��I\r'%���c.2kJ��'´޹�����������O��6�rV��X����=��*H�Z��nQ��Ew�Hë"���:X،��dt�X�Ý�voX�����Z��`9i��j$�pŴ� �-��K��\4�f�j)���zܫi�i�h�g�r0�t�LS�`�{�F���;���[���F�b��(k0y��zt�V7��4�7��P\�r��ް�y�ݵu�zQ|1����|+�������;<��1qtSg$��P�qT�7�zWnʸ�����
>�>����uH��]�~9�u�{�>�uv�����R!�U2E��nv3){]���@��\n�z2g�x�O<�|�
�Je-����õLZ���z�:�ϰ��M̧}�ʭĤ27<g�ݙG��p*�����a����=�ґ�G���s�:������<��gR���,���uP���7��m�H�D�h��c��l����R~��UX���N���bV��DW��Gt�7��C�����3혖͘(=����3���̍���l��Jg/=�k�(�g�W����2=�E�����c��6�L�,��'̈<تD�>�a�נ���N2\���ui�=/�ۇ�����H�gޥW��L�{נ;�fA���\*����~���	��ɓT=���`z/�r���{�ǰ�Gj��^u~9�P��*@�tE���%���?(�s<�s�o�o�f�C�{6�U�d֟i�����%f��^��~�<�}.����i�O�#���ѳF�hM�7\��4�QKa��H�ilI9��p�Xn�윷�V�ȫYT�J}��&[
��辕�b�p����<����w���O�n��v�������7��_"��t�A��]�2��;v�ދ^$����������]E��v���sL.97>y���N��l��f�����fCI�LK��2���:$�Xg�7�:�S>ު�7�F�D?�Yzr'���숞���a�-`xs��
�~mZ�&?.��h���Pz0z7�}�2<�ʛ�mX���Θ� '���B;q;P��ŋ͚�1�
�y�����9��U�x�`W���@N�̕��UHh�����C�=��'�0��UE�{��p�{�V��v�gFO��%��F�}GT���`W�&������<���Z)��E���q�3�N.�N��wۯ}cMO��86�=w�ɝsx}3ı�W��#�/��S�7�yỄft�ȟI�1���y��h��P� ̈́\U0&���&S�������2���i�~�⑓�)½7�~��Z��}"G���ڽ��^�,��uL�J��U0(�#".|�g6��\yz����yё��S+��$�yY��j=i�)��^��tY��8�F��9L�쉖�{�8��Z�r�ΐ�s��{F�7m���lw��;�1�_�=gxT;�L�������!�}N<�ʘb4B�Rj�8�3!�+��H��K��_x��Z�O[;5�A�7dZ�Ԏ�f�)�}c�G�c�v���Ӂ�Wv�][SO�*=)���<܎\⍕bA���'h�߱��۶�m���k���_f�h/�/ۻ3c����7n`�y���U;��V��W���%��uG��H�s�H����/#}�#�z�X;��P��9��Ӧ�Ǻ�;��>Yw��%tΙ/����b���\S��x�>��V}��箈q~��C���:��{��W�H�uR90|6�QN{N���ӐK�Q�x\{#ʫ���Ϥ��Q�&s�}��ׂ�����*�칒���M�y�#�r�ȭs�=����%f�� Tg�qz��+�0mB�;�91��C�r}9��ty�zJ��u>G�麇���]�O�I�t�d��q��y�*:�@t+�fՒ����y� �ל�~���"��	Xo���m�����[�O}����7Œ-��Y�RV=��7e;,�_��#�Q��'��۱B��V����}A��]���b��v���oO�l�;�
�3j�ޗ��q��j݁�Ӟ!G��N��z�T{�V�F�ܢu,3�<OZ����f��^g�����i��<^P���U�����7K��l7ٵ7�ƫ�=�>���^��L��dn��j�Ը~�O��ig�S<�sq�G��k��r&׍����>��z+YUZax0;g�`��L�%9�omd�0V�?/.2�`��R��̛i���3��u�L���2�"���#9���.���������#$x��,P�H&;��Y�{�ݣ���e��1��N��d����9_�OU��\m��v#�e\ͬ�Z�)�l�vOq�^Ǒ���m��-������1s�,^L�8O�u�TtY�y��X��N��:��yϙ܏e>7��ƿe�H�T�U0&��b~�RD�ˌw�=�]��d�>���{Ō����o��:�ޯ�uv���ފ���	@-��O�L��U��s+�(�v�������3�ن�}�Y���W�r6v�;��_��������udݚ�y��8٬Z�|Ϡ�ٸ�#�}�@�h��Pѧ�\U���r#ސ�g#}���yzfi�뱷+�s�3��k���L�ٿ�gn�P�����ә���x�E']~��4Fl럭n(�܇�P�{0�?��救����T�}�>�0a�|�L�����2��z�pq:������V�j��L�)�A����D�r�����3� lJ�h�M�=��MV��^q���go�e�x���hZı��U��p�5�j_�WNG����n��2����uv��L���4��a�7�����k�&��>����G*��Ψ���@�/����8^
#���D{o�xG{cƲ��\�EdxI�K��t1{]Oi�)�L�P}�,OjJ��#f1>y�{Rb����\c@�/��6���Vcօ����.��FOW
�@� �Ar�t[��7�n������(z�������s�GK�qv�#T�~ݔ��c������ߨ6��G��f���������Tg�]�s��T�si�a����y�g��-r�!z�N�o�k	��ͱZ��2�Syfpj����[Yh>t�*�Z&`R�=�YQ9�[�3+5-�Mf%DV#7��(i[���;\�pӘQ��0͉{�vOzN��OrA/&Ō�qg�В���p(�ɧO/V��6ɽ�nd��y
3]D>�z�|;%�k�hjڝ��J����ɛ}X�ڻ04U�w9
7Q��`}��j��_d.�/G"��H�n�A��d�c&��p<OJf��z��(�p�m���M��
��J[3E��"��FNó��Δ�մ���jo\������i�N�t�b͖$M^�{R��:	(]��U�K�Tz-�)o
�,�S��.��(��:��0�ʝ���3x�o�{6��gVnɼ6TzFM]�+��bNIӺ�0�j��0m�ɹ��dXp(x���o(է]%
ڃ��v_Z�x����[���,{M�NޚO�v*a͵���t���{}N�=�kj�X:��ب2�*�F61\(eNװ�t��s!�KT�i�/.�En6]뷸��!]�"�w�����I6�&��Ó_����k6ݝq�C��-�M���γ8�ǝ�Ȝ1�3'2w�q�:k�	W-޽�(,W��-W8m%�(gg��qTWIB��4U��=�ʘ��Cr�C�vSˁc@ȌxL�u��ٻ
b+=��a�y�-(����!WLU�Q�Ath�y��C7�],e�&#_�ȆE�_NÖ��A�/��淌�{X{��B��2�Y��{/�4|�
���jĐ��M�(Z�
N�R's�󅈲���q�͑教F7����n�9GRL�sm��<݋z���<'�̟�+�z������U2��nцF`f*~:ȷ��z�F���<��5��wl��٧�|:�Sz�b̀Ȃ:�>d�ji.CֽP�]��5�ۧ	��plq��O}oV��7sWv!�⹖���6��31�R�8e��o9T��m 30+��b�H�r���v=�'.h%�%Y��٣/9�`��xS����򺮂z�����Gn�h�Ĺ�:�x�#T��ɒ}�su<D��-$qs�u3p�"���F!�2��������C[蓩,��]�Z��dgh���}t~dQ��ơ.��"�:��8�f�I�sNM�ky�z�*a��+�̫�g8/�L�x�����{X�˻�mt�a���{��TFos�鋞e�V�Ɗ���:%�d���k�����H3B�[�+�3x�����ݖ�����D�5r�Tޑ�\U�E�M��Z�߉��5]i���m��a�҆]c�Nswf�\���c����?Q��7*.�+�!Z�QBDD������J� 3N������]�k1Z�d�R(��������CCl�Zr,�X��*	!U��"�ỈJZeUE���DM��BB���e�'�;��%��Jd�v\ԃ�j�C�K8g�G��KU"�=��"��IKeҵ3�"s��x�%򹷝�9"(f|�;ǐ�\�34��C*�"A9�Q&\��]�BIS)��/�u�u�3���tRȨ(����P��w'ZF�:Ph���	��D�-��Y)�A$�Q"�2�%dF����{��¼�먑j��*
�D�Z�a))��!+4����-ݠ隔IVt	8�Q��z�E�J�:�玄s$�R��|�^���x��b� t��!�������vs��3��9����;�E;��s�7�h�XUͫ/2��&sb{��ݯWr��ϩ�e��C��T���O}�= �0�[���i���G����N���;S��p��ʫ����=��j�G�s�M���g���9]7��t��q`O֯����wv��3����9��D���E9���ݸ�죇c�I��}��c.2kJ��8w\����X����zD)��p�iw�y��o���I�j���]�xa��)eS_FMib�g|i�E�x�ꢜ���z�� סT���̐���=�����e���Q���l�D��z���?wr���>WV�=rھљ����8K˪Dm.����:�=�{=`u��lp�!(CU緽�-I�����_���N�����}5yT=�2�p���yp�i��s�_�ujض��}>q��u�jq�6<�{UN̠��E�?Sw�|��2*~y�-������=�>O}��M��G�g�=���-|���W�T�T�h��%�3��¯�x��1���<3�A��}�<����ǣ�s9��F��[�y9^��lĶn��R&	�g����؈�g�2�6edbX�Q�x[Q8W0���K|g�S�k�3u�8�&��n��o���]�-_P���0R=L:�j7n�ǨF>���|ȷ]�voU�l~��,����WTsC�A�,+���L�S<75g!���-����ʟv�.)���Uͳ�C?�}��¯���e�aE��Hy�06�
�b|ȁ���"`>�޷:v��Q�>�U��ʿ]��@�=P�$|3�R��Ϗ��+#޽�{2�>5c�TZ����̖�~�K�o����1�K���Ac�$Ba���>���@y?��W�������͙3H���֌���d���wa�nl���[&��>�|^��+5��͛���M��sfA����#����Jð�O�����,��s^�Mφ��ћ^Q,i���Ǫ#�fC9CeV߲3F���}L��q��Fo�����]�����7��YzO���W���m�N���~�?����{ݝ�.k�V��p���2=:��};>ܚ��pǣ�	�7���;P����'m�~�W����K`�g��W��-M2G/m���H+��-
��Eh���Wq��:�\��(ʹ�G���ןw�(�k�Ξ������#�ps�;Tߏ{cաז_2<�R�=��k�L�N��N�ZǊ&�p�gM�ab��Y9���f�Xֽ^��+�o����*��ވ
��Q/����y07��۝:v����6�]�1��]T%O�m�|kn�ĵ㹆���(]vj��ܬ4�+�Oy������
X�Π�g�����!8�1�yUH�mx[�ϻ��1W�7��΃�F�uה�k�C�������F�n������1��QY���4=�T���\;ɔ�/&|�9�h;�z]���U�W�u�x�y"� ���s�n%*���Yy�)��6*�Sȋ>E��ږ<f��]\U�>�]u�Ϋ�F���8=�u�sޟq�u~��#�Y��qN�D�R=S-�2��7ٱV.��~��]�����{�q��A�y����w��#j/�����z�Ĵn	pߑ�����&­�پ�P��j�ȼن��-#B�ש#��u ^}��4W��w"�ޯ�!��T��3-nN����_�l�vO��hQ]O���0�k�o"�ҿQ��X��@�1-rn/��#�Mg.��^ z/v�H�H�|n&��TDӞӰ�a�%�K�c��Ux��\����`x�fC��H��\.G����P߲���u�"��P��R�o��#�V���;>�V	����<��By���<���2�z�}���.�I��Suo����2|:J�Ψ,��rE��K��-+��>�i�Q�U����yȝ��9��σ� ���V����Y6�5-�F�:h���@_��֍�L�9ݩ��Ӻ&F�[���!��z��s$������]�&6�E�l�ڙ\�x���,Gq����e5�E���,�᝝6�WX�u-��u��2�ɻe��B�L-!؋U/������i�k���֪I�c=�yk��.yW���k�Ǽx� %+��g:��/�r�E?mP��	�_s�T��Xݖ��tʔ�z��0��J�w��}�a�����j�ޗ��}L1j݁|�[�3�*���۞�\A�`�I���J��a��}��=�E�ȕ@f��ux\���U���>?)T�~��|�]<����!�5b�+r���=N�^�_��o�ǒx�<l�C�&��'}1��'7���%qί��]إY:�`��}`�Jg��#�=���w�[e�	l��'늦��x���9�uz����i��bF��Gm{s�ވ]T=U��>gs�^�V�6�=�0��L�I�*n*�Ρ��]�����'oR+����̝f�ɘ�6S,(�~���|{>��Ü� �|���z��\1�
�p-�z���w����?V�QjS.�6��P��q�g���^��K~�ѣޯW��]9�Q�B��ms��_�7��!�읣#�ݠn2Z>�چ�|�+��u�H��#�ɍ�l�\���;Bܷr-z��^F��f
gn)U
.|�d�ә/ƣ�\Ue
�k�������5�:��8~w���o��u2E͊2:W �-��l�-{U���4��o|�u�H�����fy�C}Q�n�r+�n�R��j;���:]<�̩qM�<��v�R��zGF�ie�LnE�ӧ^[���b��z�$��p�	ݨ�etޡ??���~����X*-�9 _��|����r)�x�Ϗ�i�+ӛn׽:�f������s+�ݧ��Rǧ���^��O� W�d�u�@�Q-ɺ����`l�3������넰綏���P��*�>ߪ�r�)ȗ8�z� �@�ϸ댳����1N
�F��]��o{��Zcا���^�U�W��[f��N��ߜ��2/�+B�w�&oH�{�vT�E�3uܖ6����{^)��A�<�~�H�g:��.#�LOlգ�v�ؼ��n-��`�Y@�/�.����$��>����e����Ɩ=�7Xks��n��9Lw�T��ސ=ר�Օ{̆?x "?Vu��=���X�����o�W�)zaʣ\a��#\�y!����B��9�w�z�7��+��v��碻�O�aՑT�Td֖*�����g�|�*��I��mj�5_T�nu6H}���z�!�����IFC�)��'0�\��;�ے���X��F���F��F�֋�&uɔΩ����r=μ�l{+Ü�!��������8�"��cg�oN`��''�w�vJ�W�#1���ٙ�D��7j;6�
V8:����[C�/'��6W�lW�Ի��+̲iy�,��g�ō�9��<E��m�	ƍ�Z�F����.���	g�G��	�/����B�\Y)<zl�s'v�ww1N��ᘿ#�ր��J����	ax��'��O;������}����g��Ne��_H[���V��H�� ��Q`LSw�ԙy4-yT{��#S~��.�Lߜx�_G�e;�*d�9����ߪ�~
r�/4��*@[uR=Q.�&��c��F�������&���gyj�h�{��xƩ�|��#��{#����ɉh��n*�L�<�La$u�mn��g!���_��Pu�V�[��3��E�Do�w��"ܳP�#�'̈<��5>>����U�Lz-un��yl�|���H�dz�_�A�u�^�=X�+�&+޲n�Ӄ#�'9�cUϬl-άP5o���D�M_	���Vѽ>������yU��A�<��� 
��t��W�Ũ��|�����y�Q7T��3a�͒E��MF���o:_ �ֽse^G��?ubʟj�B�>�����(w w���wU��ț���kC��w�j6^�&��Ǎ���:n�`�N;b߫��ry@]��F�Q��ǹ�O����{�6oߤ������<z������ZN$&]1s����)ߐ� xLm��������F5��N�_[ɧ���ʌM�y��+{�<LO�U��t�XOޚ�:��Y���Ǻ�i��DR-�G�qw�݉��Nֆ�Rs��mu#����koy>�K�L��Ƴxu�!l���FI��oid'���O��u '�[�l1�s���N\���~���^&V�'ۉڇ���nn�)A㨚�w
��%v�i��U����Ul���^�|��{��P{�p{�Ew�>��M!pq�8��>r�U�'f=nv�k�5�uH���@w�mg�{��Ty;C����m�l�^�;���T�!�=�E�&Ş��>��w	�O}��72��5�����/��y)�Sf�s��<���z}���5�Q��E�D̈́\U0&/�p�&S����/fC���9
�_��p��7ק��/�#��P��Lf�VYY�)�� -��`MO"+�"��7=M��=}>�U{����������=;���}��_�=Y
h3z❛= -���~���6b���Ӻ�Ww�g�H�β�Fׂ����.���D�=��#i���ᐧ|n��y�8-Ś��y�{N�s��$p��RÐO��f�5M�6l9��|���)WT�!6���wCӱ�=� ��E�L�)�@^ٿ�M
����	h���~5�qV��8}���x*�]@q�I�oN4���۫9��y '��ra��T��G���:�(>��.�л�ڛ,n��o��ԟ�����5�{�����mN����R֦` �94j����W���[�Ӎe��r���,�@����`i��Q�I�Ӆ���Fʩ� o��,��Ϥ�^���Ƀ����=�s�_���%�K��݆/�-�%2�lvQ���w|��;�g�
g<jM�H
��{,u>�6%�4{&鍸�Q�]��yg�*Kι��x�+�\��%~�>��5~U�s�:RY���5�^%a�>Gzn��N�}�������+����(j�c����@�mp|��a'C����%>��ՐD�@J�q>�#ϱ�m���a^��y��>�˝�ћK���x��`	J�~Ψ���S���U
���љqq�9ُ&[�Kn��G�9C���C�x��כU��������Ӟ!yT7��]0��L�8���>�q}�����}��O�Gge����W��f�K}7��6�3������\��ߝ�T� {O������<W~�W����t�X;)��Zx}-,��Vy�&2�Ĩuy�j�{8�Gt��s�?ƅ�н�yՔQ�y,��}98L�2�X�p�Ap�k�ݻޱ���h��L��U}メ�י�e{�ëW�����f��*c�w��5�VFѡҨ�Q˸��~5����V:"�vN��j��ZSI��,=��5�����>P�L{g���v�-�y�����	N�J��r�w�\�v�Cm�t��4�v��/�*�[.�p뛔��;=�^��Yة��Q���_k;�;����kl
��]�,]���,ʞ4���t�^���SEyO���5���4���s"}�n�\�T^�2Ux-�}���"���^.��4j{�=���9�������������,ǜm׸j��B����U\i���<ٺ2=Rݠn2Z>�]p�Ħ5ϫ���Q��*k�w��������
�qoף#�>���Ѹ0[;*d|��XZs#e��}� GL��t]vAsYN+ѵ�����%��iy�7�uNH��3f<����=�n�GvŎ�[^��(���#��te}��c�*�1:~�>6�{2_�W2@���\�C�7�}t`4�IHg��羒c��J��ǲ>��J�Kߪ�G��t��������m}�7�&�����V�Fzpﾛ����V�d�>�����ʄ�����省����ϫ���Qt��W�r|q@��=�`��_ʩ��l{M��C����/����~5�_�G:��*k�U0��͚�Y���t�BY��Ttz���'��H���q���+����q��o�z�r��)�����������V���ҺAZ���f���w>�D-�\FP��UJ瞈+�K49�w钶�G�SOv�����	���QoR���A�3Kʂ�0޼ ��ǰr�ج�$CF$�v^�Z�W����N��t)���l�{ӭ-�ٛq��k�r~��ޚ��V��\�Ｌ鿼��n}���/b2�B��
ҏ��!u�K���3�������?d
�e<��>����ݶx����O�aՑT�X�y�k�'˱���K:=�hz2g��j�7��T�m�[d�z����to}��b��F-�l�U�N�� �'���{/uk�&�Q�j#=u�y3��L�'�]�����>���Sj��ў���N�ن.q.�3j!������JL�+�p�0�nX^9<����]{NF�S)B�"b�\����N�]��r8\�Ss�Y�~�)�@-��,	�n�Uϓ��47�;^Y��F�8�E�T��'=z|Nx��Z}4��~��(�A���m�T�W��o%�3�%�������5�q��>]��vХ�Sfzs9��F���n��G��K��Kd@��j�TB���N>˳[ݾ��ݟAr��,$�Z�R�a��S>��.wpD�^�n;<b|=��4T��c	9�{]����V�Kii�Z;�&��Wqaɖx��cw�[��?}�|���f0co��0co��`�6ь����0co����m���cm�`�6�����m��c1����cm��1���1��c1���0co����m���cm��1���l`�6��c1��31��������(+$�k5S�������
B �������F���TUP�
TRP�J�E*�J���B�@@UT��
	�
(
�E)UT��	RRR
	M�8�eH���k%�(�QR��HUUUI!P�T)@���R�R���R*�R ����H��UEE*T�J"!T��*T�H��R�@"��E*!(�%@�%�
��kU%T��J!�
"lj�ݸ��(�PG  �h�@�6�V�&��h�`� ��`U
l�h)j� (T�ֆԖ -�� LȪ���I��*��p@  �Հ�M�  �4�,k58�Q@���8�ER�(��1�E�F�Eӎ4�(��E9�	(�QE��āER���,P�&�����UA�Ҥ��#p  �U
��`�ecl�6����e5�Z�1� h04��4�f��h�U�Q@�#6��*�Z�  �tR��i` m4�B��+&؀4�3ZP�F��Z�m��YP�bЖY�ִ��Q�Rٚ��V�ڔ[M�*�"V�J���   �֭�hQ�h�Tְ������cU�ZUf�̪�Pڦ�m���X�5Q�	�J�Mf��hҪ���V҅*��Ҫ�%	�$���  G-Z�V�j R��jڪ�Z�MH�e�M�[lP��ҭY�5UQ�F6�V-�m���j�m�����ɘlڵ2��m���$���R�TJN  h�T֪ژ�
��l�Q��ZSQ���[lL[CZTj�[Tҩ�l1Z�ԍ��m �cJ��e4*إl(��)��*��� ��5��m�if����,��V�4�KiB�UM&ҵkU���*�����Zh�ҕ%���-S!%[`5����ئ��T��@�[5
�AM�:  n]
Um��i�Mhօ��Զ�m�[V�mY+��P�l��2�j�a���h�e��R%��4�U �U"��$����@��*� f����!�iK[!��m(�T�[`�T��I��mF�� �fش@M��(b�E]� � ��eIRQ�  # M0� �~CR�����#b4h���AA ���xP���FF�i��"��	QU �� CM  9�L�����a0CLM0i"ʩ(M��#ф0&�1 մ��p�Z��R����|c�0��+�`e�8E/�[�k�N9[�Z�?	I9�
����Aj"
�&�UT��H@Ah���F?C��������BnHBH%C�O�P��@��� �B1 � EP[�uv_t赚�����Ǟ�QP\�mBiig��!��a��'�R�d���#f�{b���5R���lb��}��.�B�ˬ�Ac�(=����S)f;���Q�n�yC)���o-7�ކM2�(;ۤ��F��d�[�Q�Ր�5qF��$��$�e��6����Y�eh-ݷH+ˆӭ�r��zU�(Ҍ=X]�X��	�Tcv㷅٥�`YAІyY�B��-�|�љlr�r�0�Xn�N�
V0wun�+n[�� ���\�1eՕAr��	@�i��%P�.��`���t�iT�
f�]��yQ��aTYR�Nl�� ۚj����-��r�i�Y��8���V����'��`�f��
V�5F�aϷ2��Y�2�̂�F�a-���E��>����R3sԩA�U���*�۔�TU���B�q9��`d?�ͭ�#p+����c�1^E�zC��5AKM�Xv�E���,�$���]�2È��2n,��D��34�j�%Mk�lǚ�)�Ҫ�Z*Ѽ(�ɋl3JKB]�E��	e��*or[z�C���ܲ�c��P������G%��&mַ�����jV#OLJ���Zu42Z̘SR�Q�16e�m�hE�:��X��;���t7�B�c�,Y�a�I�V��۬6ν8+/�MJ��E�Ǉef"��7kMB:,�eÎ�$�EjT�'ţ�Y{)�m�`��w�D�Si�^�U�e�*��z��ခ){��c!�H��>t���8���F\�)�̘j��4��c�P�y�����ek�o^VK_
!Y��kr�N}5���KC�ͫ�{h�Cm�Hj�?]��JS�Q'�A�J�d�Q�;w;���
A��5�um5�8�Γ��w��J�}�.6�հ��ն.dR�d��ǠVf򺷁WE�t�>C,����Ĩ!-L��J��WI揦mG�-�L�v�Z�#Y��+nVZ71K�LYw*b����je��j��MZMl����.֗��Q�bh�&�����*�Y2Mi�R�VDU;���3mN �h�m	����Ca\�+KG�keH�h�Za4��� �I��]ٶ��k&a�]Yj��"X�*%��"�J���f�Mhۖ�غ,��é;t������ o[іmP*�um���eg��k�U��,|���N�P�nn"��܎�]b�`,��UfU�Op�'e����k�-����t�7�4�{���ՔH�J˨6���G�n�d�{a�*�7�_1I
�N��0#r��Z��s+0��ۨt�2<ܽ8�n]n#(6���uS�E���{Z��[@������v��+�v��'j�ջt����U�F�n*l�l��BN��m
���uDA����f��j�om+D�P�E͢w��4�V,��q���\���Q��5�����.�b��fkKA�u�ktm� W��ȉe��o�Ĕ���N�tQ��8JK{yn�y�6��HkԞ,� \��JI �ӷ�ި����WM�[`)w�@(�O7C�=�Wsh@%i��72�*�dbJ�~��X5��⸃v%��H��>Ff��ja�Jޡ��7�6�^Y��4���6��3[	tfT42�R��S6���X�"���.o,n++oV�ٓ5��q�%8��I�I�Wh��]��¦�@���YY�E�Hr�8��-�2b�����4�&2����d�,�"�Ӡ�Pl���T����*�M�m�Φ*�%C�[�Y`�cn�nVӒ�S7-�
�1Mk�5��!�t���69Q�z�V��l�PX7��Σa�$��#�i�0`�@6n:��Y��bL�-��6�Ey-J�f�5jVjB��ָf�1����$&�8ui��{H3�j����e�k*]��n	��`��5�Y���;�
zr�ǻ�٬����M�������Rh��,9�w�U�5h�>��YF�E�v�t�������^۱N�Wv���4ݴ��b�)�Y�sZ���ӢPu�l�J�l��;�1�Y�-��h-�zh�*Bj�N	1Px*���)I�e��A�y�����WU�/1Ĳ,���u�>��J%��3sT�{+9aTǘ��q�t�����{2�Yn+Z2���)���w@LH��sSm^�ym�S.8
�n�L��H�{m|�����.VM���:�����t(�{.��)����՜�Zv�
R��2�����ڲcu��2�d���a�͠5�X�5A�lf|b��r�I���d�s�D��@V�/T�1e�p����B�X8�b����9(�Wk^��a+U"�I��YYMP�:��JV�6��P%1�ӗ�7w��*}fx���B�f-���T��}/C�T��t7pE���[:�&��GdC[2�$r��,�ԎE�Mᣫ�JKJ�3�����&��'���9�&��F��c��5��*��D+Y�^��]�?Y
�X�Y�J���b�0M�h��[���	m1G�z��IK����X�,�ޫ	�8�T�n���Q7[X�R-p���N_Ń�7jc�tI`��l���͉w��g�ed��ʰc.�cb(-&�U����N�V�n]Z�ʻ:�m�%�V�椩D�T-кE� �Z6�h�,�?:��ǔ�7[���MJ�ĵU^����6�Ӥ-�TɄ��n���L?'�J�c�����icy�L�ͣ�����5��)�Wo����;��^ږLM��v��y�#6�,Vs i9���b6�#�#������30��R+��F:H�=�z�$܂�M��z>We��3ZX�B��-��r�˿��	��EʴwaK $Kw��3M�F�`�Z���#V�Ƴ��5�@L(�a�r*0J�ShJ׉J��(��̨P�8T�$8��IkRV����ۻ��33e��=�E��;F!�FW��6�ֲ��T�MV���c��1ff���(�
�V�Qh^��Wp-4�Xe� ʛ�許�NZm���b���V����IekWC �/B��F*��n�.�
	�Q*(�ݱ�2ޚ���G��*պ2�]Ӷ��EVE��cJB�n�`�r�ǁF�I�5��3m���J�v�ܪۆ�i�XV�؝�!�@���z�(�m�s>J�{J,5%�a�ժ�5Y_��]�t��(�4��Ɗ�r������Q]%�g��uf�KjQ��FH��ӡ�I���,HV�i��[�Z32����6&v�h��Vk%�iFn���	�R(���J��6a@dJ�ټw���6J�V-��ڦC!f� �Zm�e2u��4+�SPj�3P`K ����V�M��tQ���(n=��y)�Բ#Θ�.-S��v�1y�*�G�㠒h��mV��3�0h8��Mf(�A�JUdS-+��p�j�Ҕ����y&�D����EXG.�_���+2��&"N����,�EMrm3�V���w���kM0�Vf�2���D���ۑ3l���5K����-M��G�co3$�ۤ�԰���5P�4(="9	�9�"�cq�M�F��ڴ�5N�4u�z�����R���ɓ�L#��,Vں���⣦�j�y�h�Y��"-�2��[++mmQz�ʗnU�'��Q�_Z]h{�545,Tͽ��Jǘ��4A�N�<˙�.�M)(�"�T�ݼ����@�d�J�[:�<q62n�Ya�[.���*�Wm�vѭ��uJC4DiI�
�B�̥�,�m*u6�a�L`0��MC4�oj�5ͻ�wv�]�7*SIj��&�<�
 �jM#/-1i�E�H�e�sk�(蠕������&�
4�Ԭ��*�	d�M�_<���Hs�[��V�����{)�����yQ�n]6���vm۩+H���](I��Yk5To�J�u��t@�1K ��Q��	2�a5 FȈV������Ơ�@坭(���՘?j�edY�*9k2DM���2Ku�2�t�'�"Ue��xXckL��v!صì|1���r'e�Y���rM�B��Y�Yv����r���Z%=�JK�/�5H,:	J
 �y)w �*�ߵ�n��q�&�.]^@�,<�U=
F���k���N�����]JՈK	�%�1�-�2���1ZN�j��0���+sX������2j��Q���B��e%wOM\���d�x�|lTBg�YV��`VM��ZU�(d�w�t요��,ٛ�赺)�j')�[{.�wI��� �@����G5�ir�J�	yu;��{-�"��/Dǚ���i�u1�����0S,^Yڬ_�M�(tsJ��4�M+��&���W4���)Q*k�C�7�ksV�X���FMr�
��I!:�P��)���SX��rh�ԣ6�6H�w�C/�F%n��(��O%
�ܼN]�؞*�,�[����G�vE�
	C{�/i��Ѩ�S!䕄`���̲�Y�^Vlz��+f�C���Ad6j��9�
j8+,Vc�怋�>T�m!�}ib(`Db�`c�t�$��b�d���ÏC��ui�5�D�2h4,�Jí�.�tJsI�fJ8���5�I���.�5YB�*HO"wcpL��U�3r�ռh�8�\U��4U�C@_)@h���n���Y� ��eEw���V�p�Ó�M��M:�X,�P��cJ$������Yj�Hu��j,X�6�T��n�4��Ze�M��F�*�e#�6�B�2@��i��_���7I�l3A�2���(��)Y���Lm,b��[f�R:�_�	�7Hh�ܳW6��'[)�kY�q�1��)� ���ĔiEfcYDⷢ:ǒ^�kt��߅��-]M�Yکj$�݂��� (M�"�\y�lO- �U�2�%�	ح��؉�Ju�魡HPY{����w&і�m5t���ҋ���`��,V��Am-��AM�I�%��̸�X�[l��7J[�5i�	ܨ�݄� k,�fJL��2���4f�z�Q� h�o���x :fG�It�o3>-�
B�{v�Z�$�dXV�Qʑ��U�����L�ob�*�\��L�4�5I㊵d�]9�D�h�f
 H51��a,�؆S�v�����j�D4�ɚ �����;�P�l	�����*Q��� ZzYzЂ�*�`M6=�6��.���1�	z�U�n��Z��
*���"�����J/u���tI��۔���-#cZ�$�B� (d��,( 5Rv;��Z)1	�:��i��-�/t+��ȩ^Ԣ�T�jSr���F#��lx4m3S(��AAu{j��^)[��F��E-o�z1��A�+4}h �AMEИ�^]�vА��6�V)�S*PnR�/P��[H��&:�(^��t���cG�/��uy�s�xdq�7LR�������L
�iq�z���5.�;���MW�a���Q�&�&$��T�y�j�MV�����$s	�����FY{%���k�6�u���/*���V�R�[�e���p�TAi�w�jJ�q�dٙJE��٨2�N�a�d�t^Q�.� ���E�u�
����H�=J�nʺ[��zb�	�Y-��P�;�<��q����M�\Wu��Ĺ9Ygu�M6�ɵ��S5�VIG6�E�x��0�t�LCt����f�,��`�v5'J4�S̋]�u���ܥ�8]h�F�jvЦEbt2ڧ�)0>�n,�W�LX��*�F)b�ك��y�U�l�P�w��*)��"����ͅ�)�$v1Y�K��ͱe��Q��P݈�P��^-��i1)I9��t,HF�Z��K>&��sp��n�f���.%B�;���6�ط�w V[aY���E.�Bʖ�×*2�5����X�5W�a�Hrc�M5�,n���$�Ckf��Ł�Q�J�#���y��6�
mSyjM
qm���si ��f2Ӣ���ڄ����;z�Lٚ^	K)#��3.�PS@@+�s���,-���3�5�ˤ2,�q��,dt��#s@��n���'
$U�se�Y���n��,��*6oC��^���unV�"�úe%�1[�ի`�I�TTG1Y��&���LeZ��V�ј��`lH�6�>���r8(��
�����왵��Ӭp�ٺ�\n0��d�5
#j�&�M��	�7)��ѨV)F���/�ja0 �i��4�Ocr���é��4({�!�t�D��D����
�l�2�[N]c�/jP��(��K�Pf]�u�@��1�I�Q������^��ꪯ�K�za��<�+�:r��H�SdFx�@�fM�l�^
?�?��6�3���I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�v��sF�7��pӶ����ש�1��u�
�6���w-�mv�3� ��AyY ���_qN��[@oP�k���o��u�,�*#���"�r�U�M�X�-D�:�!ף�q��%k:�S�ƅ�{�/f����֋뺷n�#v�c�h�o"�V��*�@��]7���� ���Ow�w��
�F�yg�yt
��o;&�/���D�WӐ�t����4i�9�]�ʹt�.#8�4s�J*XYiv��S;Gv�e����w�w�X7Ш	��Wl\��K�׶=u�

�g�ht�H��xfW��ݛ�5�F��%H�Z���X�T��b%�Vɾo�C1���Zօ��E�坊Iz�e�-��[P>u�ΗW��'V��~�B�s7/� ^'s�pѠu5W�R�G+�!�����N����r�oK3eG�&�xݻ�Hwd���V�ԐNuM�mnN�ܳJ�#�B6��C����k9���]��9�+���b�T�@��y�����EG�<��Ԭ�b���Wjk2_:k��ʛ�R�ƺ0�S[���4�����\kt;ۉ�M{-<Cm�v ��':R��o2]m����6�>K�|���`����]��T�[����Y��WQE��9ܮm�΅w��葫Z�[�$�9�(E�	�Q���zi�ְ�h�[�r��r�l����qq���cf����ً��Ru�r���z���Z��	w���dp3!�Wt!Y�9�ݠ52=Wk,��bҕ���ub��z:�ږ�iՎ�q�7[�ir�&Y��Ϲ��w���v�d$����F�GV%��uu��R��w����RA=��x�x��Z;l�����H���U�چ9
�xG���,X�
N;ͪ��mK|8�����rG�t��o	��tN,�8yHtr���,�s�E,�씔��"�R��s�j:9�X���v{]�48�u%	ͭ"�u�)��n�i]>���_֢I��=����GM]m��k�Ӧ[99M%���Ol�h�9U���Z���_֬���ڲ���4gc���{&D�%�<�n��Wvɏc��1{5݅G�noww�r[x����ѭy:;t�n�6r��[�ֳ�޽0d�`��һk��f;=����kY�E&��,�|�l��D2�]o�L�1\K����e`OoE8�fݻ���wS�.�OK��Aن�#�j�~��>*
Rw�c1p�4)iU���0�o` ��?�����˖�S��@ӽ�tF�Ѓ��u����bn�N�ZΠ3�J��/��+&�h�Sx�Mp]5���vv�7�z���'��3EFj[uvTg/)�j-����� �))|1��뷛��JJ�����m�������Pשͽm�o�Hͷ����
|�zq�٢v��WE�c��sȚNwH�mEAݗwٷ��w��n܆�-Y}o�Uyѐ�e��k�=�����M_�ve�s��QU�䬙�e̓9�ߔ|2��뎋���8�S]t�i���7j^�\h���b�]A�]s��5s�2��A@6{{{A�֌��:�Z��BB�Ow�������g.ܮ�W=��:��CyH����4��ˍ몺w�J^��Z15�n;��C�+f抽f���͔-�[�䂥CY���}{Y�n�t���Ȳrw�1Wfj���wj�l9,)�.�16(����k��ブ#���t�b��)��ꦯfj)_rSoqp����䜥��`}u���s<�<���U򢮞����:����n�(*=�����z�1��6�\Abu��U�gG��j�^���¦�D�K�jv��J�J���n�*z6���"&��-YR��d.<ݵ�Q��3� �Y��49�r.�oŽ8���װ��gL��u�9:i\R��ƒ]9�.�#��W��9weI�3h�)� ��sp�΅c-�k��2�m�#��{�����kj�O,����2"h��j�Y���5����3��o�d��$i�3%��π-��.u.B�C)�K3k0�y�w��Ss\9S�^=P�-T�R���ҭWޙ9f��I�iR*ӫV_ي�;��R�E��j��8���w¬�h,�n�,zZKx������W��^��9�H*WaZ 3y�f�Ij��a���dA������q@���t�7��V�3Y�$K��q����L��G�G��;S�l5ST��mG@匷�j�,�)e\�]��f����RC�+�Q����?�O$�����<���L����x7*	���#���n�|��̏H+���ܷ̔4���Op�F�����np5��XWi7K1[���'%�7?���PgIb�2B�5č������h+�z���mn�]ASO\���d.�7l�sko�C�VK�䡽)w%t��3�L��J�0���Am�1e�ZѠ��w�����u�n��R�|��P]�Mq�p���DͳFpǃN�_�],/kv:��,V6�bܭͺ�e ��],������J����.��6-�\>2>[1vwb�ĥ�.�K���+9]F�D�c���r9��Y�t���z�Y��+�e�3i�4���6ռ��z�TF0�}�����?m]���-t��1�&A��X��eؔx�uҮ���P�շ��(>�C5:��͉���Q��nod��sZ�:�	<�8�u6��Ѯ�����,��F��j�Y���- �i1�Ϥ���4��˃CWU���R�����.S6-�4��Uэ�x��8l�z�ǆn��O�gv:&Wj�]le�Ƥ�*3{����n�K�ˎ���W���9S2V����iuk�Ӝ�C����QÄ��Ӻ�
�`����
p'%H�D�,�$o6�=�-�����(NYYG,m6UwW���� i�<�U�[��Ί�5�TN��ǰ�`=owX�ۙCKYGz˼0�a�9�y�`�D��������K�K��;z��L�[��kݹ�|�s�5|hs�����;�z	-j�gK��_V��G��aݶ�U��ڜ����Ƶ��J��cE�r�_v��fl{M�+V� a�Q�r�n�W��(��>o��0�Q��V(V�k.�'uPo�V.'9*1Y��ְ�O1f��P��%7ո�� �Vu��kUږ���/eJBW>X���LM��5y�qҠ7Kӝ�&��ڻg[���PM���N��T���-�;�U�ϙ�U��[Ȟ쥖D��:�4=r�\�:��v/y+7B>�9�R�i��m�95ٷ0��X��f����d�8�y|�[��n�Ư覷�'!2VG�"�[�+i���,w�b�y��<-�(��Z�9mjF��;$��L��pF���b���juu
�ۙ>��]#��s�B���%�AS�t+�{����ꌅ9����4<'͎� ��/3�������v]!�x/�b�:�����uU��"U���Y0�J����(���\u�֪�m�Y��)���h�(��f��˭/�����X������r�Ҕ9W�}a��f�{�'쨡޻�n�R�������ߥ��b��օ��8�폶ͬĎG2�Xv�c��7�(���ь:�W0hK��9�d��k��[��v�·z��`֏3ݍ�q=�y0��v�`�ioF��N٠��i).�v�Q�Z8`u�ѡ�@��G�8�{v,DK����Wvsj��#S2�R08:��z�W@L��wC�f�FJREw��f��yۚR��Ȫ�h}�l��q����.��w	'��+�uBZ��9����@��w���5�2�ή�����+�iW]b��<�f��
��ܒ��x�"�4����^M��X�~�:�����4S2̾�B���4=7��(c̵�"y����`��	���Od�L"������,u�����݃*0���w���4_sz���H�^��T�x7ir�[/��QuL������{Ko�љ(�V��F�ԣu=�[���q���/6�V���5e������پ��9#�v�/`kP��J�&�f"*F7��ϊOm�nn���
��VFQ �y�;��;@>-Q�j� �}�R��XHU��y{(I�1������L��1�_M֕ݙrU���厠���h����[9UI%d�Gu��5a�Ø��J<H��qgfşj��`^�p_ �o)*�E���Y�J-e뜸�ja�h���.�F 6� ��V�@��=J�üv�7�S�T^�@����ʀ|�p).΢�z�8M��-���!����ǽt�&��@�[Ҽ���5u���;/�B���m���t����;y�2W-M���L��/6�<��VE����֎�k\�E�_�*��ˈ�cP����*�t���9���;�Z�:�kj��9B���#��q�\8�#�U}]��"�ù
c�5M�)�[�Gل��[��ܒo4sݕ�=��(�F.�P�Ù�&c骮��.�0kր���A��]f#��{-��/e���ZW��Z�YЀ`�/0�S� ��(4j�����{и@��R���b�� �ZY�9�\�ui�#��
k�%_}�]�9ǷN�p�Ӓ.Js|��v��Z� v�-�����}:X�K;��n�'J-�iX���K����ْ��.TzLImmv�.��L2�E��ޭ\M_K�`�k�q5�++ {���$�T������#�7Ħ�LK]�Ľuto7� �J�i���y�.��H�9](��e[�7���NU��T;�,��,3��,��q��Jɯ��̺�qS�Hlq��Jyι�����ܛ8��cCnW����n�Ðd�8�K�k��r���7)�;Zܰ_j�=�rf�L�/������jH>�����0k����7f= mt���Kp�W{�|��#w6��͝����D�Z�k(t30�-��v�ҁԠ��1��O�ƌ�!!&=�WmΣb��QopLKT��(YL�h�Z��0��V̽mZ�'�E��7N�U�ʗ١�+4�vuZ|����Ƹn��sZ8�4��'0&���x�����܈��ڰ���ƹ�[������Es��=�-f��-�P�3{�
ʺ�7D���6�.����B�:������#��:g�VT��N�wO�������I����^�+]��]�2hG�z���W��2��� �Kw��'�G3N	�M4�Yw�:��T�3I�8��Õb�X�����pv��(�׷���N���[F��Js��2�2s�܂�e��`5X9�;K/���ޱ�6c�>��twn]��a����v�c��#�:����u/n��B,v!�3+]m�M��l7���烴u�Vt��*^�]�_wdw��eH�f-�}�l��5)g}9dsxc��۳������FeH{��`�##�;Ruf�8p���L=>�2J�Ԯ��[5j:���7Zu���|ݻ��ʽ)ֹ���� �YsA��!'�[��j��H'
�e�]_C��飬�G
[��#G/��mqGV�롔%9�˲��A��8R�����5��-��N b�靾�}7S�����U��r��ZzJ��I�V��+�9�c�@�� �3w^������Y^�*-R�t��L�r�b�B�)EF*�����=�gN	��c�bI݆�7�So���=X잘(�j����w�V�i>w�����ۮ[n8��.��*�r�fI\���C�o\Iv;޳5�3���������;]#-6�9;S\�a�eB��_��>��j���p_�.Z٧����t��*��Υ]\�0�*��7�oTbD�ά�ԏn��a^��n=\���E�.�>郅��n�fs���o����Ͳ*���%C�l±]��X�d�=��o��یw"pw\�O���8k9�϶�s��[�NN��v�����j�:�w)�����֪k��3�=���M������v��:�}��oq���S;��I�1	p'yu���7�m�Z��3{s�EϦ�ݦ}����L�Z�`�!q���Ӭ��ժ�BHP�P5)+1)fZ��"b�xÄ⋲�n½�;���4L�T^����{�*��i��Kmuu�1Dd�/i��j�g�]��;�u��Z4������[t�:�<�3u��K�X�C�T����/+�3�gd��9$��]�!qYy�u�$�*��	�E.\nr�mQ�K�Y�Z�\��6�=������;��y�WT}��N[W;�wr�ۏ�.��r��9Ν;������-^��P7���V�-�.�U�%YW�$�I$�I$�I$�I$���=HT�Nf�Rar�K����B��YA�5�ӹ.��ݍ�F.�--����Oz���fҮy��ڝ{F�bَ=�of�cJ��i���\�������[]9ˊț���(D����I$�I,��,�v��n��A�M�~��*�BA����T]Wʈ��q;Lh����;�q4��V��^��m���6�1��	�mu�r���myUog������i<:�b���1�
�+��V�;Χ+��:eDa�}�x:|u��a�W$�.��M^lO)��i9N����v7�Q�mR��g>vD��ƛ�*r�V���V��։|�v� �T��6O1���U�2�Wǋ�����y9"�;��k�q�*ˏ�F��PӷM�w���9��
	����ō�����QY:�{YN�àZ����M�kZ<�9�+�j,J�m�w`6�<c9�N�mv����{ʓ�Q�u����t��.�
f�Ƚ����9Qe.��J����;�t3��e�i�b�r9o�b��L�ZV�*	�ևi�St�NX�U�pW�;1�x��y[%�Y�iFr����nwd%*�� �:v��NhU���j s�I�OU��"�7:s���H&�ƺQ��.�{�t��5�Q�YF����@�i��h�+�9U�o��AS���F�;���@P�S��9M�I=�2t���T��noE�Fvq�N�Pܥ�I�H��
2���\���W��֝'>3`�X�(x�b��6m;�j*u�Y.ly �ѵS��u@�������qz�����7��-�c$z���M(����p��v�x�Wa�r�S�ɥwe��فj�`i�zK�o(�8���gx��ӊ��ޮ���;+)���/�2e���b�;�V��\r'��w��Jv����n��㳐M:V�j�Х��7^�E���ǐ�ͼY��=ƾ�S#J����K�@�%�y�:�ʔҵa�9."Ӑ�a;�]r���;�Wg�?MnŨ�e�<�/,p�Tf[�,Լ��KML�{I��E������N��$#.^�7����R��
l0�)ʍ!�(.�p�c�jm9��dr�֌Ծ
�+�롔5B
*���|;-�I#�v<K����Zq�8�q��*mt�J��R͝N�ûˣ�z��
ĳE���ŵ����2Ժ7�ۘ(3_^�w�ԯ����k�]כl�b+� @]oEc6��$��&�T��)�]=�b�G�(_Z�:+c�J򆤢�
̈́����/-�&�������
Bf�t��XpA���J�-�n��)�j	��l�զ͉H�q ]�o_;�z�ǚԟn�}�.�
���Y�I�rfN��e���Ȕ(u�]WU %+�wfn��uVM��
��X�\����8V�eZ��S���]r�������=�f�z�� ��F.�]3���S���+{��
��RJe�]:X�`WM؎�1��g�f�(�2Dѷ�u�L;V�C9i�C�5n�ֹY6]07�	-���}�F��sua+�/��meJ���Dp�E3a��Z����x/�w������W���I[R�A윮��#3OeY��pƹ��������Dq�٢X�r@J�w��rq��9'Y��x���J�G;�������r=p����M)|7����uЙ�j �څR|u��Ćo��z;�)�sz��H�Q��7�ruf$���}��+�������� DXɑ�s��12�#��f�Ð31'�hXV�ݖ&�|%�gqk���N�{��Z�ml�q��vipœe7����C���Y�u��Z�<�|	����*招3�۔E��]v��ѕ4�=��]V�y[��J�p��L�}����/jfʾ"l�Eu�2���P�k8��No<I�Ջ�-�C:� �5��2#�w��)'q���Q!�$W.�ŵ�+*#6���&��Vp��j�*f�u�WW�aμ��D̺G��
�m��A��l<�R�i.����u�2��$��<y�U6�À)��p���t�*��?8$��[l��n�I��P�"�]�뗓g����{�l9�XZH��mGhL�LU�Z=���|\��ҩz�?Hjs�f�a	o��K���f� ̿��o(F�D3p��m�*[u�����A�!Kz>�SJ�����[n���X'b��gld��B7��Z�kP#6e���G��s��H���r�a�$�w\q�S�z��O���B��u��&������A樁#u���E}Q��k����c�r��բ]E��ӭR]f]�us��Vz��c�2���,X���r��R;�DV�RUw��fa��$�O5�[��e
�����$��T�*�����j��i�'H��+{c��׺�8 b��Vw�l�*��D�bXp�HJŕh���>f�v.&�
�hZ�1W�ѫt�����J��a}��l,N��2�E�[0ʋ>s &g.��;x��\�Z�ZV+F|e��4�t�U��E�E]�;i5�ܥ���f���n���zX8v���D�=֝.O�r,z�C���t�5�4Ѯ�M\lwt�Qr�9X���j�ɷ��6��,$z�삌��K-�����V�zDO-J!��ZX%��G�j}�Y���	��u���xI�ev�E��K����JY�3\�2̿�3K�1��4��Z����^�w��Y1H��z{�
|MC��mǓ�r�^*O::��[:�2MKw����_�<Xhَ�`tdE`�7��X��Ի/��� ˡ�P��:�̈́�+	M�];�?j���wT_3����*���f�5$��(6덺�n�ڒ�}w�tT���j\ܸ�C�yg���[���'of��ŹC�b�m����1ܱG����Q�S�����[��o���r:��0#�|q�˗���n�8V�����#��q��/%��-5E4��=�B��fM�V�h��*��а��6fG׼����Y\��̥�%���4X�.LY���;l�mv��M���$t}�ڷ��7���JmJG`_#�X��,�li�|X�x��f�w#Yʞ!z_��l�M�4�ʜ7J�f��`]+KS���A�1u�;&,��7��);�t��oN�k������9mu}Eѫ�lEt�Z;V�N��u)
�[kT�s19�u�L��	<4o�z܋��O{4J�-`�\���r͠��Hs�󙧥!PT���%l$�	k����5۷�T�2�{�'�J��'i�"��o����	���$4�#A����t��oGG,c\{��
n]�:��h`��'Z�
�z.D������Y|�>�+������&3v[�	i���l�Җ�V����_J���rn�]�X�o4�!Ҟ*��˫<[{�)�Yk]']s�Z���pp��p�R�j�:�;�7�S@��ފ+���L�%зݖڃ�^�W��$�u��ٶ�[9�=0��4��MڂqRV2��
�g��'(i�{X��ҙϫ�3>|h�S���0J4/N�X9��.���t6��o���e��ޞ�ZZ:4�l��[���vm��͡It-�ܧ)gj6���Ĕ���9�>3��D
��(�'4��rKD��(].�j.xS�h�uR�u����
��5�`�:3K���Otz�&�^Y�K���/N���+fWD��XJ��J/���iz�dmg 7�JBn�����3���b�����\���%�ԟ �f�D��$���V����#z�����jV�����唻��mƯt��V28"�Un�]�V��kr��h�Uu����&�q���n_iɶ�CO`::��э)�j�A�\+w�7���KR�8����Uܐ��$���+��2�S���=�m̧R�^���D]�;���n�gv��꘸Q�����ú_R�)ͮ���Sl�M�4Ί�9�vW�.��nO�b��2��fDf�96YժY��k��zY镪8\��B�q�"ݻ̨�c����:܎���Zu^�p
}�S[��1���խ^G(Vm��O4�a������R�ٔo���S�R]k�k��A�n6��ݣQjf�m*Vw�:��S�8�²�n�:�!�ݴ2��7g��*���W��N��:�>/����9�zϞB8.���]c]e���9&�@%�!�}ub���Vb�{u-�|t��C��1�9���٦����S��m��q�Keś���ӷ9�w��Wm.��X�]Ӫ����Q��ʳ��e�#(��N�v����Ԋ���x����!�џ�l�����u��2���v��������w��M��˔7�5ʙ�V�ګ�O*��V���F���� "�˃�����,��qֻ�l�N�@m��R6X��6C�D���5MF�W/%>s@Z�Nr��ט��{`*kt��ѷY�^����x8*���4�����)�yVݸ
�BA�;�Z]WN�U�q6�Cc�)΁�ٮ.�v��o^)��ش{�:����";&;`�y�^��F�;��u��
,:yδ����먈�9Z��Ð��Z��ƣܢ>����=�WX��D[55Pt��L����<(�4y@s6��������:B�Yk������'"8%ݢ��W��i˨��(��-o$E�н�a�r�nLh�&خ� ٙ,��Y���7��]�&}m�Ʌ�v*㥙�c����7������/�Bʻ�;;��Wd� ����R7)fu��y;2 �E�Q��'�*s�D�yCF&�)s)�gSi�i�p�5н�n!O2�Ә.��u
"�����=�2�r������1QYē�f��uhƵ[\��BªZuȜ;�Lv��5�k�O�̼�]�Z�c�凋⢤��t��*��X_vl2����ٹ� ��I�[��������&���73xձiX5wD򐦻4!*h`����j�r����2��8vb�+��*�}��٢�.� ��x.�� �r�*�.ӼՒN��ۻn��{TF�Շ�]�ї���1��ۂ�G�����F�ɗS3��U�a�Ch�3VT�����3�!�fu�J�G���/�χ�o)VuJ�;��1�g@z����)X���X����5�}m��RṚ��,SC�J��Yt;���Vvd��(Z8OjM
�E2I��i�2���{�7@T̩maM����Iɦ0��.��7/*s���F��-�䰱Q!v�U���>$�]��`�9��R��1e9���Գ���G��i}�R�Tf�4���K�Ww�wѷنMr+��]�&֩TO
�Ee�\{��N�ȴ:�W�����:-Y�ke_t�]{��9��\�-�Gl̻	��{�����vf��pv9��SBU�yAnJ]�#jf�H���f޷��v-�$��ո���k\};nc�A�1��8�^�a��:�[Zl�6��Q�������(L������v�7ˊ�[�w5{rB����m�j�vͫ�j�ܠ@�С�`��Ż���pX�w�);�i�X�kA�����F�h���Y����o�9S.�35��	����z0�_i���6Z�V�ڔ���ٰ�sWM�W�kF�s�D����M�q�4�B����u	wˮ������@
�oq5��?*}��*ړ��!��\˳���P*so�&sFZ*GW[���5�-ybl�gUǙ��o-;[Hب됍�rZQ/������ԯ��G��h�]n�@��X���gpTڼ�Ն��>�7ךw��I���(�Ihu#]�xK�݂��
+s�fT�Ԁ$@�xθ	X�N��S��'>���;R�{{������u��'F�毆g��uҺmZ	:X�x��B�۸�o�|�uڤ��R���2+N��~���3���]�u˷�6�_da��;s�[�g���eJ�-ڮ�ͶJw�FԛQ����n�;��N�]����׽ ���.xh�{M,j��k�Vn���Jiv��,�NTC��R�:�U�ѓ%#���F6�%�".wkÂ��O/�� ��tV�{�^�6�����8v��Zq�v��j;�v:�αt�u�t(�}n�ʕ�JI��'I��z8u��I��)��ʹ3[&^�{1�0*Yl�ޮOZ�R�Ci�7�4��]C(#3��.���U�TJ��� �D�r��ˬ��ĸ��ۃ���D�'6�m:�W��H#}ũ�pj��,�������i�IN*[���b�VJ?jQ�9�JGgou�U�4��f��*I�O9�r��XtN�N��Xz�Q�2oͤ�߇e4
1C�\���f_>=��FC]ݷl*2�9Q���\�N�'%>Ѷ�7��$em$pR�Mf+��]K���*�x�A���^*��:Iٮ�Ӿ3��+VQ��;�j J�/��G����»D"w����-�CR���f8%`��U���|E���ݨkq��P\��^�T�4+J���oL�u�A�/��_>�P�Kz�^�jU�p�|������eբI`�YMჁ�fHS�E�^i���j���.��z"(U�{����+i�ZiY"�}7jV>�ڥ�r$d]�S��e\�.j���YC�yW�������$AE�����χi $x���f��I$�]����فɌ"�B-�;�i���[��}i�E����t|����=V���
풱;��iQV�f�h�"���G�|������TԳ/X�f��x�}8��Li3$u���7O��8aT��Z�]����������޹j=�'c*���rc����&����Q�8M=�/��CrW�Ӯ�t2e��@��/*ʬ�ն�ܾ�unq�|�]����ܳF�gP�f�ԭ�7Pa�)��X��_X�d�Wxpˊ\��k���|�BWN���M�/�xQ��XhiQ���a}H'���"CjV�V�9[�wl]��p�z�I��^�n�l�t��=�d[�Ę.QE˴C͹2�d�oa��̶6�Ĺ5vw,O;Zv�Z&��w\�,��Ώ=:�"a�����n��vY*vt��Dz���|���Q�@W�
�Wb��.3b���X�:�@t)*��%=�pK�]�٫���q�G�rM�����bm�ǝmϞX/��J��4�6�0��G�i��Y!f��U�X�T��|i�=�,�&���4�/�v�������+Q�d��h���F�ޱ`WlZ;��y��j&ѥ���ǚr�y\PQvT���Ő!���I��$���{�⪰�����;�;�v��ʀ�&���	�%�R`*�u��}Fj=Ӓ�o{o�c�qfqaL��$��2q�6�k���t|�S�K�;"s���)��t��G��߾��]Y��m�m�.Z�����������e+K
�*(m$�LVkZ˫��ƌ�1,Rص�U��L��әq�11����31m�fR���Ⱘ��+*�l=3F�X�q1��`*��9����J�H�5�˧=�K���Q�
�X���&%5t����JcP�p���$L����e0T�f�q��UW2�0�����lLkQ\)��TWwZ4�U�2V���N�j�ff0�ck� �U���T��*WN������f2���Q/�\,EQ�,�p�BԡZ�jV�Em����i(�\ʢEP JT|���2@���,�)�����vm�X%J�ku��t�\,)]emTh�\��ɷb��U�ZՊ��0ĩbٗ)���72V��ӑ2�8��-3&��I�c�S�+���Y��6�ފ`m��Z)m��R��b+ҋT-J�UXQ���.QJ-i+�S)�ֈ�\\���X�iKQj����Ҋ+Z���5�~��cd�����uC����*F���'sWm�fPj�e-���O��y>�C�$#��/S��9.�3����wI�TWNQ.�"C������{������3G{�uԨ����/���zc��	��yy��:���_rٺJ�Rn'��-������,x�ox{��=���DX�t�b�+^�M:�o���	�m�:��\�bOE�ު�ަqh�uA�ۿ6)7��@Ȯ��<��^��[�%n��t�:`M�z�b:����竩��q�~޷}��nm��jwAh8��F�P�葓�w�:��w5ۙ~)��`��va��b�ޭ�Ĭ��pd�k��Uz6�_�Ҟ=<�oNR盯�^�\��h$��U��7n)�Q��;�f͞��= �j�퍄&��}ܪ���Knm�r�ub�/�=3�X6e.\cim�K�4�@�Bj�3y�O9��������h{�oK� ��!�g噰/<Ip�%a�b��{o�O�{���=���*m�G�T���X�@���wN)�������r6�lM��(;�e��)O�(�-|������GwC�.���U>�O'T=Ej6�ܨ<���آ��E5���}s�Hn
hM�g��W��3��r�|}���O{����e7B5���=C3�t�I���%�����7.���[��6�󐲼1V[����s��~]�O�VR3[o	���iE�ls��kOyj��o�� �($���ոו��
�YX���=	��[�K:��,۴����גlp�hg���ޛ��ݒcdxw �wWqٵ���R�|�����\tf�g(M̻�AU'.^�O�>������P�t�Ŝ�]�NBT뒭����f���쫧ݩ�;&�9�����N���K����)L+4D�"$���v����غ�r��Q�y���Y{B�fD:�T����V�Œ��]7�Sp�A��sVL���BX�8�F��8ǜfa��]_t�~$Su�M��d��*ؖ�&�ð�����\�Ν���`ު�yaLNʹu.W��n��R>�Z�����#�z*���+�9]ȱ�n��8�>��ăeK9i�ΠzH{_J��u�΅wI}NM���7��]����w��+��VNS��c&=�Բ�7֮��F̘c)ҼfUR�������5e��<���:��7S�\��T^L[���W-߷%
��ZO��� ���D")/��}���EQͪ9r:�P�n�����Y����(Z{��k�q��{}��ñM�'�����$�r���&�ؙ�Jmu�����7����]J���{������Ҍ�����x�DW2cywWk[QШ�۩k����b��_{ԣ�jz|�/��Z�dK�T�;V�a���a��y�O��t��a��N�ށ�L�*q<W""�L��Wg{f%���.!���h��SiS�ӯ9��Χr,v���6����H�뭱!��b��N�Ѕ��4����y�p�����YWh��T���'{p���ˇy��׋�_�{_������Cy17��������]WK{�mա�A�<]jH���1�ەt�Kػ!F�
u�����o^F�{�����K���N�sFdd�]]R!��wK�3gZCmT�0�Tt�g@~T�X+��3�'�y����n��yy(�q�#ڕ��f�����d��Vϭ*ɱJH��-�塦amЅ�E��:�B�y��F;�w͍��}>��ۜ%<�AQ����is<y�!vO��W�o)�:ns2!��i�u`s>ǆzy�t04�&r���	L.9cm=�\�p�PUfͱ<�Eb�-ʫ�&N�'\<Ѹ5V܃qT�D��5M[<;�aĉ�p`�`�]zx˞sR� P�px���1uN�bp�j�S/��}�Ly�.��b*��鷕f[cj���U�;���I&�y�~c*��+��΄���Z�{�6��8/Φ�����Zܷ+������X�/���Ǧ�=���u�d�`랸I<V{^����jX�/7�٭��^k�z��9]��a7�N&��E�;�P���v�7g]qw͌�,ɑw�V�C���h���{�&;S-��p�5��7t�"�-G����Ԧ���;���>Q��"4��l5��Y��[o�8�s�o�_d	ڏ��e�ڹ��ܕ˥!� ���������T��L���5��q5��T[�m�Xz���ށn8<�����V-T�0�Eަ!3�}�E�arQˮ��eZ�ǅ�;�]�ڡ�k�#�����D�4��u7X�'�j��wD�\��1��e��Kf����A��-��W��d���T�+3W�����jL�]sZk�T�U
��k�-��61��O��ۮ�+"�����n��������w�6�C�Î@��/���O�b�cd��e��T1�Ѕ���|���y�#Owa��YC��|���M��1��OeQ]4�,qt��m�.lv��؎RTܱg��tS�9��吋t}~�v#�Aؾ�AOP�
[�wy���ɋ��Պ�!��#Fu�PXI���J�|n[�h*گ?{�W������81z�︚��@*���P�w啱�ǹ��ݚ�Ƴs#�nk�=��q��@���[�38v-������U�+b�ֈ}�nf;]Oz��n���8N��]��;�X�eo ���v�ʴ&,or����[�w��v�%5�PhlcLPN��n�`�7�k���m]J��QصCe7>�tJ3���R���.�3a'����|L%f�6{DJ��S=�::3*?�-G�����#�e�������y]��B����7�һ�
�.nrf��C��o3!s�o(=w�;SŠ{���iogBKn5\r�ܡ�*|wm؜�Cs�ЛL�.:;��t��uU��.�{�Ӫ>ט�Q��ޯ}��.�\��٤�bFr�U�6����eK��wP��s����O����l�rP��!M��_s��b;��n\�4Y�u�'/��O�gn;�4�4���Lư��9}Qi$wj��Q��Nu:��ֻ'j���چ��uI�Z����h&|�֧��R�!��9�[*��SW��N��1I;��>��F�Ǖ��^ޣ��͹�����f�P`4�)�q�
�`Gi��C��CÜ}[E)�Xl��2u�ÝͶ���ף��h˜�;|�u�3z�
Y��μ�����eww/�AR��;S���Yk�^G�,�ԫo��T����t��a�s_<����V��<.�W��t��k5�Q<��
TX{�7�L��^*g�zEN�u�	���o��Jf��Ԓ����9^�<��li�[R�������c�zN[3�;e�y�.���qW�N
I�
��BU45Ў72�$VwO(��/q�#ۼ�.G&)�z`G ���$��B�	徍΍��z��SSN1�k
�c���y��w�L*�N�F��� ��\f6�Wo&au��e�	�#��\�{��p{��'��U8<E�ʈ�O���ʉ�_�E�s��[�d!"�[jGk��RA�W���!�L���[{ |����J۬��\��Ƅ�Zfi���r]��[�yF�ν��򼳶(���ǯv��L���ǜ8_;�e�&�N]��~K���kǗ���[���͉��N63�9�Is|L��\6��]R#��j���Y�[���[Nh���,�3s�t�A]Y���n,\��k7��s��oVU�9��=3WwBk�!��7 ���o��y���[�`��7���a"&�R;�� �t[�;�]��9��V��i��_c���v��q=4\�cZ-*v�t�w��Z8�>K8hw<�l���=}]|�Za��v�=��j;OV;u�_�q��z�]�-U��8[ϻKVuT�k��kÂ�Ɖ)Y�r���z2^���L������&�qݏ�����j��v���8e_��՗C�C|��O������(�����駡)ٕ_��[�T��P��z�*���ӏ����Vsݭײ��mO�Z��h�)�&�ЕMomE���n��3FW���b�|��ͩ�q�21�F��;	��z�t�B�k�ڝ��4�V;�!��+�+=p�&��A:�G*ۥ*��Id-��_��ȍ«Ǆ�ɫ�0%WPw-�C�4l�R{+ڎ�<��zpô0��8jr07��T�E[���_�=e"���?�p	S���uн���q��8����~�����l���r]_Yw��P$vQ�v�E�kI��� ��eR�c:uq��*C��V﫪L��薣\�u7%�jh�S���4{�y�΅��ȩ��\]H�"��`����g�q�f�w~�U<���S�V�\��ܑ�񽻍���v;�S�%½���yڪ��y~Kv��������{QU�ƨk�>�;��xect3�41c��(=w��2+��)=׺^���.5r
z����}bb�����tf�K����m�.z��u���e[�¶�0�t��vP�b�T��g{���'Փ���I��n�+�������H�/lTj�Nz�.6�Ɂ�վ��]�o�IZ�?j*S��ŕYd>��_�����z�{�E����{5|���:����'=��m�5���yP�T���BJ�9�3�j��]��'_3�uZ�<�O^ЅY]�"����U�q8���v �XwLn��]���76�X�B��`�G�x�i�+�i��꧎�nZ��#���P�kXh�����)��w������̼��d��0h���ei<�
ob�ġ����w<����Nۨ�$�/[Y}��l�މ���:»}w<Цc���dʰ70P��z�w�jZ�%YbS�Z��9PVS����殧u+,h�"�a:f��� ��L�����%B���ӭOvub�s��ݑBy�%SB�؎93����S�
l�OE]O9U��r�k" TՈ|�O�7�K`�	�@F^G�yy1z_�L���.�U��!�ߵ1!'e�Ps���氺<5P���w��d�)�o5<�ǥS�[�R���F��oJ���au�w����3���8���.�. �ۡsν�<+-���ݪ��<�kv�5gF��r�B��Cz��J7�����&}I�BVСy�͊|�@�IY�bgZ��:뤷{we��z�{<l�>�O�J�x*��,�v3X�LN�{�˩nR��{A�̛
�i�Xv*ǣ\�I��������U��{ʆ:�V��?�m!ǃ�F�pW����ًaGq=����]Y6	V��N���w_5B���9�SM/�j5��u�����>��ӥ��JO�-�j��-��>���0��N����Ԏ�ݶ�)��`ys+ypV���Z��a0r����gxC2��K�� :�ut���Z):r�e��nԮ��1Wuҕ
6�����l�yÜ��2rκOC�j�s��Q�f&���si����L��-P�$Zw�j�e���� �J�Љ.�i��i̳r�[��0�.4�K�ܡzMf(LR�n��czG�] Q�S1<���0�v�V�Wr+3y��g7����T�)�G�����o�z�3`r�B�Gg�:��q�H�]�{���\�����ԇK�vEr��N�r�D֝��J݈��<ْ����w���J�f]��v�A-a	<��ݻ��l�̕�<���u��E%�ڋ9�P:kmy*g"��"R�o���V��y��=kV��w�n��{Qhٽh�m[��Y�G�8�fP����W,q«7u�a�����z��=��V8�]�+vznM�M�!��mͱ��c'�x��&��j.�{����5yN#�����|��_]Ӳ.>49V��.�N˾U�j�d�$ƶe���j��	O)`�})ee���ܗ�F��:	;t���7�#c�kM��J�5j�Hh
.��뛻�k�4e��l�̋A��:�b��x_���u���$�I$�I.���dΉrsx���JqB���u��'�uY".��u�\�,*�۵�]w�N�8Q��a5L4��r�Q@��ݷ��2Nԛt�nRg�+�u>�(?����Q9��D���������Ρ���eb�Ʃ�����૥M+�6P=�x�Kh�c-H��&�-� +���5j�a3����oR�x��WN����u�:�U�>\H��L�����0��:1ƥo%.��Zd�F.f�{�AWgQ�V �*"F�B�]�̷c
p+ 8u��G�tu���H^�W�RŘ��m;���/;
_k��0+0-\��	�.�A�u��QD4T�z�Z��!�=�x�%�� �j:/e�7���'��-��(K�^h[�c��F��*�Y��^:�(��!��70ҝ��r�ձ����^��=�/ ��(�L���3r���V�Ƃ�s��U�q	e��p���U\�TJ�ب1��00vy8ṝ�+�J'@A�;G�����n$z]՞��Ɓ�6�MJ���M�޼)�o4[�ơ�c���`��;[R�Ͷ&D��BR�Ǎv�:5�qԎ�ۇ9FS���m���ɓ��O:	9�pw���-f&�w>�99�wM�;9I���d��;��Ν:~��G� ���}�W(S��l�MY��UT1�Z�("i+?&����4Z���R�P�]S-)mEEV"�j��t%Ǝk1��L�YQq��T����1W)U3[�Z:j���fTAt���=u�C-���3������[UR����Ɖ�f�V�\\q˖�ΰ��ڕ�T�V�
WmSMb+��s*	���U5EM�) �%��"�j)ir�4�"�LM7Vk*�ֳL2�iuM3�\������V�.V�LKkm�ej�"������+���o�F�UsX\�d�5���$�r2�4��O2���<L\��+nc���0E4�t�!s˽Y�Y����A�i[b:�\���s."e��)Q3y�Y]�]o�e�1�Ze[�*�d��3.a�����2)��̶��Ʃ�0�R����0��net�֋�+�pM&�Qf#o֎�X�l��.Q��fh�����Y�G)�1.``T��JZ�
��[[�FU�\r��\�y�Lˎ-ʸ�	��T<������j���xh�Y3�MZ����M����r���K\��ZQkL�-˅�eʷ)G.�ɬ,VҰ��kF�]e����r��M�(��(�-�ՙ�3-Z�Ub��:Ʌe0ʡZ�.9��|L��/��Ϊj��&wT�ݓ�̵}��O�L�
��3c����٫��r7�u�tr�G9gL�奐�gZU���7)���w��o���IU1�7�#`���vogI�=N�Z�i.q��r?��U��������̋t����Ez5���M�C�6�L>m(]�c�����|~�V���_Xz�'�ۍ������|�p��jM����OFݎB��`���3r��9M}?T>U�����iy�\��<�BӤnl����*��Tr�ow�w����(ρ�O�g��?�����1�I��)��P�;2���-�p���)�ܾ8��CI[F�� �Me5r�hBq�rD���	Wٯ�Z�5I.��H�����sj�*=�?�c�JX&�<���.�L��8�9Yz�e���y��L9n�s��y�=W��~�<� �& ̒3�6U�4HkL�9�^;�e7|� J�ҽd�J���������W���O����ד
AN�y�2��`�Z���+P���V���y���*�\���c�I�:˱j�lԊY���m<������J\��e��0�pG��vܛ�'3��R޺�r۩���Bc�̎��w-gRGVv��6$����m�H��=JE�+�3W�:lڜ���9i���Qܰ�I3�L9X���ˉ��a��k3�J�M�a	��m���ɻ�ִ�~���?'}�{ ��(�m�dO���m/��R�?+[Sʽ:E\ľ˝{ʫ�����j���߳mn�7f��A��Y94��UQ���i*J��L���O>7�lϓ�x�Sw��r���bn�dۑ�A@�.��S�U�VO�__}�3�g7�V�޷��o!�Z�*�>"j�0�W�ت�DP�N}\6�Ƿ>Y�S朹�V�r8TV!��TvUɻkjs�]��Ԡh��T)�4���c��r��v��.ou.Z�����}�!X�Ӝ|�	m����ђ�A��v*#iˮ�j�����}힉��Ϫ5w�/�0�r�*ˮv�E螱�wNk�_ *7���:���u�J�lR�'䌷�6����3ԩn!�x��R��{/y�:��(���B���,`{|���nr���Iv�����{rf9���M�u�t�N���jx}4�o��_p����5E��bkJ�Ҹu���%��XZ��غ�oc�^�Uɧ��*�/Wr��ᕵ�RX� ��ͼs�����.3��fi�%����p:KhOU%��)�w_�r�ΐ~�T��՝4�*���kT
v+�<�'%�˘s+'qZ�.4L�0VuƜ�	�X�®0��9�V�"d�g6�r�7z�ތ����e�:'�MG�]@;��a�r��_�̘��}�]���U=�}�4�|KV^��U�P%�i@�33N;u�˫��B�s�c��M^d�4L��?O^��,+�-�3�x-�@�2{X�W�]6{�H�UK儷nm�9A�E�]&X��5z����c���U��O������Hו��|�9�W�fD�^%v^A���8��6�o��,d�����b��%#��8�UYj��V'�+��9��tG;ꚋ����y�~����S}=�0je߹�>r�Z�W�iV�s�����v��R��V.�|�f螙VUdUS�f�Gr_���rc�h�sVc�3j���t��^�wRf��S����ռ+�ƈ�,`�tb�9ȫiZ��lgJ�ڷs�׬o1���M�t��ճ�u4��9�ޅ��%�6C����4����:x�x���$ߪ7�gm��_y�o�{�'aŕYgχ:r8H+�8�a��L  3�&�k���=K����� ���OɌ��i������|��X�����d�@��2N!�LC���� )8�Y'�<�0Y=E	|���f;�f��og� >�D}� 2 �&�a?$3_d6�a8��|������''��<?RB�~��q��iɾd�,��A>���=����tnSt3����w���QH;�<��S/P=d��7i?0?$ۻ�$�Y=d8�ĝCl��Y��N����$��`i����-�"SlR���}�J���3�xa��LE��	�%a�����'Xxr�'�a3,�T��Z����ݙ��Ŏ���a���I��I�����}f���;��3��!�@}�E��߰�I�La��a�V3�:�N0��dXx��w�2���Z�2�y�?2��2i��g|�<����������˦�� H��G�xD��qY'Q�:��,{�
��&Z�2C�����,'Y4_�OXNxf@��&�a��Vv���^��s��˿t�}�u��~��xHt�0��x�$�����]��N&s!�`s�d�П��2���d���zԓ�޿B�O�������$]�'��=�d�Z�������=a<a�|�m�M���4����x�ԝE��H��g�rݒi��2I�Y��m����>���Ш���8��wX+��MT`�J��L���]�bc�{ `rP���S���s�ΙW37E`��������072��p^:�~��اx�/{��;�)��+W!Ww������޺�m���f��G��5�TyS�F�n�H��;�*�[r����	��)>g�O�� ����I�y����~ߐ��,���ԝI�x��S?{���L�a����|�eh	0�e|ur��υ ��� |��m��%`~�'��&٦|j��2k}�� ky�qY&���'d��{��>�χ���vq](�}5�o������i����C�<OY?}�����a��d�2Ow;�QB�0���u5d=CL��hY'�7�'I2n�g��#�}���B/�����崵_�{��@�&�;�ܐ����垽I=Cg{������C�=f�y���>a?'�,!�B��d�����N������#�>x�:#*�q�_?�̟���z���R}lRO�6�M��0?3_��ǨN$�?fC�~ġ{z�+�u��2OSs�dY>g��I�Oa�Nw>\���ms�������[_>��>����M뺓��?>2q��$5<��m�x�!&�9�~g�dP>f�$�6d{�@��_)�π1kj������߸�����&���6ɴXve�2jo��$��yd��q�!�I�=��������B���g�� n����I�7�˟J�����N�����g��(�N���Y?"�{lY7l���?2jo�j�fs	��'5d���!�Ri���ԅa=�y����by�o�6�o�G�����D6Ɉw�'P��y�Y'ל�d尚�q�5"�u�'����ߴ�z��MY:�����5�s=ׇy�[="������f��g�f�|Ͻ��sP�'���aԚd�Y�k�!�J����d�I�8d�$�>a��<Փ��m�{�C��{��s2���y��)y�r���f�W�F��Mv��wZ�p��\3^��)z������lW{*0����"K��(�W�2�nxb�(N�{Ө��ر��elJ��7_(��.�w_����g��5.���QGr�:I!+qa���w,�k�
쌸��[ǲ��O��C�zɴߛ�2LB��?!ēӽ�i��Hw�I�&"Ϲ�� T5��N0�(�|�u�,>Fﶎ��]K���ݸ�]���e��i�I4Μ�>d3tx�0݀��ɣ����+53�"�8��!�O`n�Hx�m���u���GW��{gO���Y-F�Kͅ�М=�LO���w2���і�������d<M0�M!��H(c'S�"����`uI�Ô��d4w���� t�x��W9��w���A���;a4ɹ��~Bu7��x�Y6jÌ=�u&��I����O��|�L�Gp��E'S��u�b�ο^�s�o۟&1��π��(�x|�������+%d�/�BN�"�Y���XM�04~�''�y�N��'ǶLd�
���s>k�mlW=�/���v�bt��C��&������~d<���0�i��+����BT�w$��0�d=a�MO{����<���}�v����^mny�;o&~1�$������P����;��|�����n�z����I��ßa��LC}�I�!P���P���>a�M!�~���G�U����NT���? �{��p��I<}I�'m���'�8��S|��ݳ��	���Rm�	��߹��~t���=@2w�,�g�C3^_�>w�?w�������4���C�d�h�O�k�''���'9l����=x�c!���Ú��ԁ�iğ��?����� m��Gd�#u���+a�G�~���<d�N�tdP�!��2mXh�Cԟ2o�XO�5���d�~rN�q��Hq������gr�>d|}�;_+�zA�ۊ��3bч�t7Cj�]aW�˲]�&��R|�e~!pî�����o�<������)o���*�2l�<TF�)Y��[n��̓]iT��3�\U�k���,�{Q��N�{1meuݛ�3��h�Ł��0��%4u_cV�wO��T���菽��ry��������	����4,�$��L���"�$���I��]�$��'��~g�i:�Ǭ�a��O�����b�c�����o�O�,�t|}��'-��<I�u���O��5=�
�5��R~E	�g|��nZ�������|(�>G·|��u��������� 	,�|ϼ4��̏���+	��a�و��2c??�f�J�^�I�h��$���2yl�-�Xmg�4��{���^o�Ξ���W��`t�]�+�l�3l����q�m�M��!�8�6~��A�O���,�2Ufw��VN��,<���>�O��.�4�v:٢�i%G3��>d�'r�ԇ�G�����Y��l��x�X�$�S�d8�2M���|�C9aԞ2b)�7�'~��{瑕����8�s�v=�a�~2��sf���F��`|ɭ�����}I8��o܀��M��I�=ϲ@8���I�)���穊n�����z�i[z� �3�L@(��3�XCG?`��~a9�d�W�La��Ԙ�{Bq!��N�i�I���SN=a*J���ǷU����o�{��rE�|��d8��&�~�P<d�a���@�k9��$�&�`���I���l�-��I��&3�	���{���bw�����yU�g>�f��'6�Ny��'���a6��ΰ<�C�y�Y<d��y�*B��Ĭ'Y=��P�8�L�6��5��|�p3���*���o�뙓�����{��d�OP6���G��8���wd�f���u��d7�a�Ԟ�a�d
�Rg>Ȳ����P�:�~���D����X���7T!k���H����/%=��n����6㩧�Ӱ����H��{z�J>���Qo	�:ͻo��/�G��S����3�*���1V���pP�Δ�<�Cd��p�:+&�֑b�J��)qQ!b���\.r�jK#���'� �3vV�N6?{�H���G���$����O�Y?$�,�y@�';i�����~���� ��ì6�29�?0>I��I�!P���ϼ�=|��{w�3�k��*f��i��ެ��4ɣ~��	�M�k$�)&����6{a�9i����K������g�@��a��3��&�>���s[q�>���I��|����{M�)�l�!X|�2m��Pd��1d��Ѿ�E�����O̝��|ï�dS�x"<i*�@}�D��o߇j����	�}���Y���>�d�e�S����׿�Y8�R���'��ٔ��:ɩ�`��2N�$��<�~d�l\��i��~������|#��} �`u4sY̇?Zu'���/��C��
d�&�h��E:��M��̤>I�M�$���k����_��{�~�y��zO�d����O�3�08�Ǭ�倲L��3��<9�!�%gSs�kP�0�o��?0�C]�	���@�>dy��>���e�]og�UlZ_���x�4��3$� j܆��'>I��O��=g����7�Y�O�'9�q�b|��
�2O��@�W��ݐa,?|�֌_.ȩ�V��E�H�:[���ZE�̞��d'���XN'�����|��e�d�g����h��~���Y��" Y���}n�7�M:\��>�Q���E��,�ZIܿ z��l��`u&���蓌�Y=d8�G��C�z���	��r���$��:]����������,�����R�}�#�A>�_�'P���pud�a�,R|��>aSl������&״'�C�}����|/c��z��������f��w�͛���%�:)O�ớU��/3�0��H�G.���4����M�/Y�M�ѹb;�˔z`���r)�dv����n+���o�V`6ƭ����m�x7+�=�S��o�X�ܼVVi�U���u*ũ.�<<>��d/�}�s�ۿ���-2M�����C�q��<���m��XIԛI�>�0�P+g�Y'��L�䓶����2{P }�������X���C�<�=���Q��v���<|>�=��a8�>�O�XqY'����"���`T2��y�d�4g0XN�?�Xbz�s�2�x�Y?w���ks~����J�;IyM0����Ol1��^$�N����uY'r���Z}�u1�L�7��a��z`�{��?�iʊ���f�vkF>����ɶC��,P�oVa<a���m�7�x��:Τ�{�I�&�uI��OO��;�$�7�a��d7�d�>E,bwN��:?Eu����� O��緍Bc��`��>Bu�&��O=�'Y'�6k$�:���&2qO��x��:���'�O�XsVI�s�tw��O�F��Tr��S�WOg���σ<Bw�0���O!�{�@��'�ȡ6��~��|��4�P������:�z��e���7�'Y8�'��~@��}8[�����ή���}�>[ :�a���!��̇�~���|�0�l��O>��E������6Ρ�Ր�
>�����=���̂G��7;�o�˾�����t>`~�䟐>d�iӖC��_��ש'�y;܇Xx�2������ݓ����Ȥ��+��M��zj��ɤ������~����������1'k����8��Ĝ��|���N'���g��O^�:�a�>g��;��I댛��Y�I�~�O��G�������F�z�ͬ���zϽD�!�O�57���2O��?;���<Hl��I���߲C��r�g�d�;��������O��;������a�co�;�P9��]-G;j�mL�p�Vw^��!Ѹ�Z�F, ����V��T4��z-� 0���-<�\�X��
�[#ow/�wܩS��SP�j��Y��ov�t��]6�d}���@N>v��f��ԥ����F_%�ѽD��V�rK��}�>Y"�@R)ȤX�"�((�_|�3����?�Cē����Y�OY6���8ɣ}֤��7��?[	�o�d��x�`x�C�~M��V7���2|�������������>��}đ'�+���Qd�CS��d�,��g|��(�q���kP�`o;���$�xj������i�C�z��u�菔_���﹊ߟ@����>�Y����:��1�����;EI�9�0Y>�FS�$�60�a���������'P�~���~5p���Z���Ͼy�|��8��y��'��<���u�h�Ѵ�����C�6Ɉ�|�u!�J��h��u&o�,��I��@��7�'$��G���y�k��;��|��yk�M�:}̕�BuY��M&<d�!Y����I7��P�'ʐ��C�=d�Y��:�����'��^��'��|f3�l�i�i�s��v�*bN��z���3Y�h'Y��z�uO,�4���$�
�O����,�Ou�h�;���-�9'r�(���M���ҽ�~?XLd�o�'-��
���Vd8�3F���d5�6�`m0��AC:�9z�VJ�r�Qd�Oo0:��G�%Vv\���dv}���Y��@�I�ܧä����F�P�`Oԫ��R�����"s���:����Q�����YtC5�U���\�Yr�Y�W�b����Um�u�o�y�o���߇<�b6�����w��LN6rt�J�/q�7/����l}��j8��uO�P�+m�6�]���BH�4����X���\c�Ve��G��֏A�%��D�qw�*��2�8�B$��Km�,Z�W2���]o3U,�bƾ%�����mu,w�5#}�ݼr4wkS v1:v�P�F+��H^��d���wfs�P�\y���ݚ�A�*��!�R0fq��s�m�������QmR���I����f�����k7�_�HmF�c<�sR�qؚP+(�X�f��Z���]cJS�V���Պ�S�uv�$��o+��N-��K{(�GG^r�.9�Ջҭ��D���m"�7�M-al�ʑ�z{^�ܧ�wӳqe�A������w'3��n�[s���m'��Տ	�-b�2��xw ���V���X/�ӹ_�����|�+�բcԋ�g^�o��j���m�ԦA���%*�4(-^S����C^�x�:X�(�2΍�+Zȼ��Zk���ٵE�Ui���z�L'��]�-I��U�a����{{³07ɮ0��mh�f��K�:��֊��z��r:A/����}��݌��5s�����w1HSAky��s���wl��b���E&V�U&P9��ݎ�H���y�O]�h`���	5<]�бyk��)�Υ��x*^�T����+���Y�T-3S}�3r��I$�I$�����eN=͹���܄@{ƳM�L�NEM4����hZ�pj�f��ۺ��!�	3U;Z͔k`�-�A+�S5R ���;
��Ƿ�!��"_��Rì�.���bce�Y���G��l��j2���+�שq]�MV��6��`�n�T*�-zRN�n�x�lpm�Z,j��a^���):�f��n�>Ub��VU2At�]�ȕ^���ђ\b��֣�
��#5L3t-.��cqh�N՜
�t��(�(̩���"����I�T+�k����R6��������I0������$8�wƛ��/���(��_^NI���"�3�0<a:�]�]\�w��8�#bB�%٩�<}5��kZr�)���}n����z��=�O5�n�8��j'U�T���
\΃09v�:�2|j-�۴���Ӡ��+��P��@�~iV�y�H�@�+l�v,���j%�s�_�qG���-�T�kĨqvb��̡�]��h��䩇0�F���:�uΙ٘�M�k]���^��@eS����ow+H��O�1���e�Y�{P����P�0nvi[�+���r��L�p���wF�՜wv[ĺN�t|���髧Wg%�+��]˒[�˒]�~����8e�L��o�f*kY��KR֥
be5u�J��YW5s+���Q�a��aQQ�Sn`\�wL���h�3��-�\�T-�\1;|�M�r�jŉ�X�5��ˈ���TV�\ֳQ�[s��9j����)��0���L�f��7W#�\�8Q�fI���\J\�p��rֶ��L��WUH�8��6�dG.f.C�b#���[�<��&��7IL����ꨈ��GIQr�r��������[f![���e�.U�֋Zm�\��3-�2��X�h�&5Y5K���(����YE�·)\KR�"��Q]Z��嫖��X�������*��1P�*卙�,̬\�PX2�Yi,[�Tp��f �]9#Qb.҆�V"���
ŋ*\h�ũ>�:���k4Z*����1���J�31B��Z��	�qr̴����YY]e�.�k���֝���e�:Lf��kU���Y�S
ۗӦ�Mr8ϮLj���ոҍ�����]Y��(A7T$���d�Z<< ��f
�v��+������8�Ų�]���y�\�J��-���m�s���$�eu��E�
T��[�g�����bu��w3'���^[g���Uֵ��ʂ[[��A�x������5�Q���lDjI���6k5#J��ׯ�g�vm^dK���jj��o�^���3%�Uߨ��aY�c�"�k�x�T[��tywMa먯v4ֳ�M�4����u�_��uN���3}����UT�cnj�<����UV�C���򠶽�;�h_�TӞ�\Uc��FF0Y33�gsrڧ%jX�������w�0ϳG:r8H+l�<��{�G6���s�-�E����
z�r�NN��KN6����~T�+l�Q�Z.%��x���d���Y&�.�w~n�w�1o�ۘqAX��*�څ}BK�f�UG����Ó��=4�����.EF+��Z��S�r�[���P��*�z4��72����*�21�:�4��K��2�R������+�h����5ܛ
A�YD:S1���ެ�*M�wW����`���l�=�p�W��Ԑe��a�to��������cL
��6��nZ���XJ��F�
����������Ńt>7��;S��ݐjR&P�>h^���at�(��9Ub��טJG���ͩ�ֆ�X��m�����:�F�B6'+�Ƴu�;Q۹o:˫�mBx8��$�j��m�3Uz/:J�f�.�d��̞A�����0^6(pQݮ���һ�|L ������s-�;���}�菆�y=�E�w�������ݪ��<�-ۚ�Uݵ-=����[ob�;8��4��y[s�4�W�P��lXԊ��sUr�yx*�K�K���i?,̚Iey�;��!����&g5���U=�r�^r|�e԰嬱��[בA��B��P��"�٤�@�U���F���&=YRt��sY�z���5��U���Jts��b��6雙rϽ���9�Ce�R�J����H��1��Z	�r80��z��[ہ1�cb�}�s��b�IFU��4m&X�����/�uv�[,��v�ĕ��7�[^J���c�u"�=+%2�>�9��O-ԹVMd�r����D�G�{~��vә�oQ�^K95�]׽)��Ct�R�Ig��������ڻ�{D�_�r�OS�]�aOD�ښ	*���8X����P�S�;�{�Xe����Q���^��oifs]UK�x���ݹ���7��.�����JB�z2���-�֕��zXr��[8�����/WO<J+f�L	���%W��2!t\-��W]�"�p\K����>]9��2��JN�s��y�30���q�&W@ǒ�Qӂ,��M�J6d���U-'�W����d^��~��r�5��Mߝ�%���~��NC�N�������E;4Ѹ<�u�e��'Nٞ��듦�'��A��`�ۍ��.���u�w�,g����=-!^g��6��Ԝ�u4m���s�-^Cr/%����k�֊�����z���;��smr��sbrf��u*�~��c|2)����<S�ۖ;l�ѳzm)�͌siT�jnV��p|�}yF��~�V��0�)��6�ى���t�$0��o����Ŕ�5d�2t��-b��y��������^^��f��q��Ru�7�.���[�w� �Vw)K�Ut*?�ԝf�Yٓ��>+v��94��y_H�B���kkj��]�E��������ym���ջ6�&�6m��K�r��-T��h��k��6݄����$:��U޹y8r��W6�*�	�)�^��e>=��jR�<N��vnG]u��U<�Gq����q�拉2�]J��k(κ�\ϏA�Jo�v�a�m�Z��;�8s�H���T1l�>�u*�J���<�Nֲ��.{��.������������g��f٠y�C*-mFm'\V�yu'7aV�GS���īfS�)r���VF޹<c������]ا3",���y�=��B^-�Ί���*S21*�D��n�T�ij��sf�X�鱝a�vwѬ*;���F�"r��b͐����Vc 'j��Z��S6t(���~ބ����%�B�����3�x\�q򂥭ݼ��9��چ�f���lwN��Gp�:JL�[آtZ۝X�ܣ�3J[Ϯ(��X�J�mu�][0m��$>����S�Zw�#����li��$V)��kÐ�1����V�&&���I��E�[�G!�WJ/r�]*rݍ�Bz���Q���Ƚ��6A~z"Fs�A#w5���jˠP��.-�n/y�l���p���;���9�^�5����i餞n��r��5�=�G�3�׍�V���.@r��ڟR�3�nGj�Z�8-ݹ�Ӕ����r�o'!��ۦ�5��t�9S&�u�b=V���X�=y@=w����<..H^�Q�z���;������VlZ����6:�#��h\��m唪��鞌}ٕ�}������8�˨�R�,��k>/�Ht��3֑�RV���\�����^^zI�ie���9�������U�{A�� +�ڊ�W]��Ѽ����%��	�v��;��9Ý9'�m�<��F�f�����;��>N�5�f>[}�Π�'f��Ӣda绳%%�3"�*קx��i��}J�g"�m�]5�{0�ٔ�o�L�t[�%��@�;WHg�|_}�̰�dɗ)�N�!�zN�gm�A�h �y�������;����=��s�{�{Po~�M]WZ���i��w6�����(�.^>�i�Y���ӷ'�[��>���O^סVwR��%RU�͝�A�_��]��e�nj�/���a�C�4{h5:mv^�Wy�X�;v.�K/�\�/�:C�O��/:)�U�gѦ�r+�;|�f��g��w,�	����B���$J�
�6�-ߦ3y���k�t�Mi1�i������9�oLW�N����D�wΜ�Y�J�W�#�o�Jn�-+�o{�G��Qᩈ���M�!�-ay��5<]��1=W��\?f]l��m��S[��WsA�+ �RX1-�qܘ�U�f�޸ܑ���r�{+i���9��U4<��㞍UT�"�=�޸떻NWp0-f�ߧ&��BE�b�R4;}�����f�D���eZD���۩�š\/%���k��&�˭K��+��h�����ޭ�|�hkr��[�x.j�v�#��c��ޱב�����O#á�F�-�q��(��x+{��gX�oClP�5�wԂ�+7R]���ե��oUZ᲻*��\�l.���ۗ���6�rdR4�����\�O@Ǵ�nLZ��r�s��]a��޼�5��B��6(�4��d���F��Z����_�鴩��>S|����m���\��}+��靥ˣ��k!�q���ⵋ����:|�8̅~��-��욀F�4�+f��Ǩ�T�H~݊�k��B�Q��ؖu�0)f��IT*׉H�t�9&a�n��\�'{p���!p�%m� 򮅞�����U}�r�,��z^(��l�|��+��|�'��"��V�	��k�w��kgU�֑���]�<������S�3O�H�lK�ZfEԭ��9Jp{�Iao[��'��㔰����8f�&P�%PhZw��+:&�Q˰�^t6��LD?jٱ��X����s
�v+��-3>�%ܮ`�9�����M�`�cU�ǰ�f8=j�J�Cb9��B��� .!'|��R�Fv��c�G�i�U}���	r��ܒ7y4�g�՘����˫\LK���S�ؕ_;�C*�*�*Oh�q��+�����B�#���p���r4aѣ�u3�3a�(E|+jn�lC�u:�0N&�Y�,����fw^o3��m_ї�z/9㗃!!ai����1Р��UQ�η14������tN+���J��J��ܖ+���S��h��1��=hcý������o�����fj�Z�tݍ�$^�#-��mD���,��/R�	ls�竻�/p=�Eu㸭*m��7�.ʋW=��V�S�S�;��V盬z�8-�ٿ7�O��ݧbrP��wL�Q����f��Լ$C�ċ��7�h�Oc���v���m6+D���h��V�C���bvf�ٮG�bFo]���ozm��De�Wԛ�}���&l�]��-?9�tبަ;.=C��J�4�9�Uja����m\U�T�s��At�$�`�Xt�\UfۯbY��JӽV5����)ө.c��9�(V64����ym�Et��J1Ze�ڹ�I��w���Gp[�tV�ww	sv�$�ԏT�T6��a���-1�*�XL5b��V;�˛�fdCWdԚ�,�}�)�ʸ��ՙY˪_S�������³m��Ie���JN���F߂�g%�RcзH�+������wp��ꜘ�:_T��C�M[��V͊N�W�#>o�E���7i�9 ��;�+Է��ڪ����嶺���뛊Н��)��Ts!y��V��s8�pe��J�'�̭��냝��CxgѬ ��RtҬY���[����2#D��q7�
�r�g�C��;��2��ɤ74cD����+;�s��g����^�e�s/Q��쩷�m�ˮ��񶫾�qi��ѻ�|Ly�.���"��Xt(̯B �|�y���Hg{"�us�(u��u5�OM�2y�o���k��p�
U�΋�֣b!���ƈ��(e�k�صEbǚ�2�Czr��:��=�L���}�K��n�X�"�u\�"�3C5#A[�z��;�2�e��)��׳f�t�n�+�5��ȴm��� K�Nu�bڨ�A8!Y�Z�/��L"� �s3�4v�6N��P)�e�9�MU�zl��[��ր9����mY��ҳ2]�D%�ZlV�,K�d��`9]�+H�5�*�_
( �#wR]���ܭ}	��՗�~w�C�V�y��HlԶ:�F����C�Y���sؘ�[{w����"���;*6lx)�)3ؑ�Fʧ�Hȷ<�ۑ�\��Ӣ�,I5;��nP��T��$�*5O��q��pi��\�D���
��=Aasϓs��:`_u�!�+l��ݳu��	����6��Uk����GK��P�
X�m�P�t3��6M���*Yǝt�K���9���i��J[1Ѿ�5��R�gL4ފ�F�p��Y��酾���c����N-��س�4�?U���5�.����F��s��b]CK��g�{�:W�杺�V{��z>@��*�6%'�jS3�lSBu��=���M(e1���U��ʲ��)����a`+�Ѹ-3�����:��ׇ¦]���pb��3}/f�o���U{"b�h�V�@��:,ج���|@ǜ���l�}|���N��'19�&�¯V���a$6����˳��#Tm�J�v*s�Z�3�iG���r����GS�̡��T�|�M�R���&��]�ڜ8�.���J��7Q41�6!��"��Z�w�#Ξ�]�.���`����w����S�U�ɿ;�ѓZK%�U��h�Ь�Mf�Ã�o"lѦ�ST�g|�#Cy��+~p��$Y�\��@���b�
��gr����m�\뙲v]��)a�2��Kl���Rfd�h����,IJ��=ڦZϺ��9WE}'#���J�!X8��˨V�/���Ȱd��F�*mt��Z��̺RZ{�م혿9N�z�{f�4a9��<�Gb�}ۀ]s����_il�yt�]H�ts���wB��)nSwx�uF�����{
��>yh-i�c�줦]8Ɖ�w�(��5��j�5==�|�N�>`�א۝f��n\��	z���t�k�3uL8�+6��3�/���S�)l������;��Y���98�Ol>����K�-�C!�y�[}5e���qI5��+"T�it�V��e�)l���p�h���0r�w��]���IcfƉ����.�<�n`�/#�wԒy��L�3��1����Wz{��J� m�!s�*D�
�O;չgWKr��L���D�΋��n{�m$�I$�I$�������wDn��jQ�`�ޥ�<��𽖛	�5���ހٳ*ݖS)��(�S��Z׵.�p�r�6��JL�(A(B#2e ;H��<ݣ�k��s�rܚy�_�#�v�������wJ��y� ���l���Ki`ڛRu޻�8�@u"�N5�E(�A�m��p]5��;[A��L�}��n�v ��"�f���)L�������e

��tM9j�p[�̗-�T�G*T�p�
бnܫ%O,ϋ������,3��V�ɒ�O����]w�y�Ԏh}�ǥ�*�$�oM�Eڭ��R�g\q�L�FV�-�43Hw�*�⮄t�s���f�K�Q���0��)MX�vw1v��z�`�F�z��D��g�vV�CBN�ɽ��}��F�o%Q�d�V�j��ܕ���$���RR��,���U��T�6鮸/�1u�F��	���.@׸G����-�|����HZî�r�v�|�R5܍(�N��3�]�[�F��x����B�˦�sΙ{}��q��Rr�P��H[�T7ܻ�V��qQ(%ҳ�.��ΏzN��z�vE;�wlsd��%�ؗ$��\x��D	"=�L�[j(�(����KmeS�L/�wlb����
UDDD�i�fT��R��QGMPqF�ZQeU
�e�R��TQ���QX��8�P�E�ڕ��*6��s�a��F%�E�Z��PYKTU�(�%6��ҕ�[j��TR�j"�u��J�m�h�jV����YTb[*cf2�Z�i�jȉT�F�7��"hX��KJ����O.8TDm�-+RP��-��+Z�h���ZPkmZ�k��h1EU�cS1RU�r�)�`�S2KiA����-r�Ucڊ"��R��Y�FڮةR�W���µ�)��+�q�U��ˀ�F�E
��Jyj��j:J
*1�9�0W���ƹJ)X[J(��ZĴ<ʨ*.6��j`��Kh��Z�e�`��~��P\i��Ͻ�_v�N�ޘ�_p<�MKw��9Z��(�b�hR:;:
Z0)]���T�\���^Vj텓�2��o%�xxxb�햂ǅS�ʺO���"u'��#���������H�w���U	�3�k��r�Sc}�G�c��9=4եjm�� ��y���t#��`z�ٌӚ�7$m��n��/13t�T���9��Y�u�c��`w.�i��0-b��ɑM�z�	�lVjF	\��&i3՞o�Ƭ�w=�����w�����U6�rgԆ���wkB�"�f>���s/x���}ϣ���^Ew�~B��.�g����_{����5�p��eȶ���ڵ�B��}���A�K��i���7��u
��:��z	��k��=.m>O<v�VF�7J��of��ᨩT_wK�H�aH�>=�(BI��W����}ד���}y7饊@���
�{a�:�z5��dgyKc�����OW3�����'�qݯ(p�w�/#��os�ڋk�0X{����==6����v�7��:}Esm��b����ce�m#8qs�ʲxM�#{X�o��5)�%ʄ��k9Q�7�*��\^�ᑚ3�:�V\�۶�
2j��uʹg0"\�W��m�9�����hVe��i<u:�h'��u�Er���alA�+;R]��< �{z��J�+���]�sb�;�~L��h#>��h�T)��_
j��Ċ�Kv���c�i�.����$s͉uhi+��V�H�;�Ɲ��՗W��ȃQn��T�3��,4��B�нz/K'I��_��U8a�1�4�P����r2y�;7Clő�0.&�TgF���U+���W��ʖg:§N�BPz�X
vmssY�F�n�T�#�OA~�<����r�e\�-ڰ*͆7�3o5���٬�I��7{:�j��F�q���Ć�k���W��n�l�ڕ�K��f�n�]�Um���uT�w����Dֽ�mN	ɚop��u>�Ϯ�^�s2x\j���f��s�-�ᱯ���X1�:�V���S	������;6:�x��ة2X�%p���d��F��X
t�x4��'���8m���d��X�-mlp�ܫ�4����3,�<���"a�u�{/������=��̙�
5���[Y��J�%���+o2_r»��p�\�X'5c'^#o���x{����;�s����c*/�tѭ�po�߇��ne!���{���е��r"�nw/K�,/y��}���k�Z�#(:G<_�Դ9ˉ�>�+��/ac8N&��m,�7VY��y�=zV��u�F�U(1Z9P~.�W-'��W�&Ep{�z�]L^��]NJ�F����$P[ԍ�u�W�#\Y�#��S��UGLlh�`�Bɮ���k&d���R�M��cYH���Nz�{ QL��5�Y�bz"��i7�g�p�)�ou�x��b�z����;6`�N0����bM�u%HQ��Y@��;��B�B�!��aY�?.^	�V:Q�-�O����j�e�`;�RȀn*N�IT\���9���jr�|����[����6W��sda����o��8�C�we�bzC:�F:�a =���u7^�P����k*�T��O늟VB>�!��)ɨ\[����"N�|t*g�{;�/�zYd���g
��لc)ո�K=�5�w�+���/K��k��S�Ek���10�.u�j򋥢�	�Rآ�¢+Gf
2��f	��%��Le��i�'yp���8+�5i��E󁵮l�i���{\.�l�X�}}��2v.7�#.��z�|������X1Y�PRs+9w%�{����sulojs�W�Y�s>:�qCX�!8��h��֐D+�um���ބ��O?m��f�ǫ{�a���_���=GYB�Zi���t���4�:̪��E��Hʻ��)�|n�xL����զ�^����Ώ :=�$�U�ؙ�<埨�.�gpq��HI��δ� ���&��p�8��xqɟ�8%�k�t:-nf�Gz��"�j�˩��nd�f�/��0xީQ�,�7�xpǺ���tV�ۣ-�2��x��2�J;�uQq�:&�d�"��Ɗf]��yX9�6��.؄Gw�H�J�[.#�1t�7�J�x๞.�W.4�i�7:;�D�X�F�X�������C�9�ߜ�"�P؍:Y�BxDc}�s�-կs{����Ä�^!����С�J��`W'yQ�To�\@w����x酜��5�´�D\9f�����q:͍�r�%j���'e����q��Z����%�[�u�;�Y�ΰXI��ђ>;a�0��d�!�N���n³���ю��=�Iu֒z�o�z_*u�P�	�3���twSu���J�Ya��]=���h�.���G#"���W����=�<n��z���yG�G���=��.���
x���xA��Je3��Ǔ\��/�{s��b�v��}�GA��Zd_�R0�A�C�:���l��>�?L񤚛Y�:�"�Eb�ϧ1)���E�J�C��l�f+���#�p,�qLG��'j�;]$zk[��8�hyez��Ɂ-H���$-�Bw����1�=+3b8M�l2�j�=��[Ԣ�^D�S�*�8M8y�L���S&���-�����ј:���n%D���������;%R�?�{i������\��"hr����ۊꩼ����zdJ�y~�,�e�5_���m�`��٢���(��XZ�:*YY7��w��Z��]Ԣ����M�����欘21�^T`Q^2�����0l�,�.�m��\;�O��&�~(g��
�V���d�u^7��o��%٨��>Ua&�:զ�fO&�a�F�8���5ծ��p��=t6]U�N��v��TJ~e������O�ޠ��/e`<6�S����삧kbl���^�_Ct1x�׍�lRR��c�����FN&������_Vh�:��G�Ho)Ήs��j����WuнdWe��O�h�p�t�*�:6M7qp�7��u=��v]�g!B늶�ˣ��8��^��\�uF��;�>���=廙ԥ�ՙ9��]:$u�F$\"�ϑ]�j��C[7��"�Cp�Nw���mOw �R�uP�M�����K���"�5�U������Hw�m��92�1�u?fp�6�t�{+&�Gd.�:c�OJ5j�����G��p�w{G�����r���Y�sstD�^��Ϙ"a�قyF�S�����#���v5�;vs	�)�n�T�T`��̋
C18肍BI�����R�}�f��ֽ�3P���ܜ���)�R �S��UeE'4d"�|�'��R�].TD٩��.�y\O�������1b���[�lM�k���؊�T��U��R�$_�S0hK^C�����ȥ��/8�:�z�*��T�X����I2���1��:�`Ϛ�7&=����q���VkR��8\BVQ�z%��ϩ򢨼<��?WFJ��#�0Vu���������o_Q$1�f������c���.c�f�9B�R�躆�,uR԰�]Ӏ�H�F�t�Z;��4���R���w��hu��6v�b�վ�5x��-n�ؾ�kx:�6౳�%�uvn9�9�]��܇�[s�!�]+�%� �������y]��s ?�o�ct��zaug�}�p�=ՋG�)e���Kn�+smi?cy��t':�j�`(�b����J⍀���_x�ƍ�u�t�yՑs�Dq}��2� ���5�s�观������Vl��p���c��n��u��V��WLV��u�{e����'l���L�5�U#F��<j԰hf�$м�)S�����Xz�wT�q��xL@�J:m�&��J"�~s�ȡ0�/� ��5lOԸ�ce�@gH��O�)�9U��Qk���;�9����B��.U�QH�f|B��hLk��b����q��6ֽ�X���):uD�s���o;zV��PᯛF��R����u��WD#z«s�q�S�RF��eC����"��"��O��Ʃ ��>�:I�"8�i\�^Vg!�]���i�'��[g^���3o�����#<u��/�������ImcR]��Om��`g�-c<=�9�<k��N���̪�>uģZ��4M�U�YԲx&3�Q�wJ��7�{�i[*d�yyPm<g�D��r�����"bݤN�+(�u.���jƼ���V�p��e`�?�o��m�	nW	���n��;��ӭ�x��u*��sW%��1y���V��}�{��^ۭ�gg���D�EK�3�~�<n�f���Pˮ6
�Ӈ�t_r�O�Zۏ��A�P�4=�,�W���Vq>��U��/>ל�*>�������e%W������� ��;,�7Ў �mu'^�Bb����G�y�?
T/dR�#*VF��jp��.��TS�0c��z����ᘥL�"'���w{Y|	�/qT��ٓ'���;*�662��H*;X�!8���Fp۞�A
�`�Tz����h$�0�B7�����Ҏ��֎\K�HczF�ʒ{Uj�~�N���	�n�w�\��5i��i�}]�*KvF��;�p�T�k6Yb�p�MtYuڪƮ��5��w�<�o\IO{�T����v"���%a	+8��_g��m,������:qN�^u����wU������Y_9ݩ����0k F̆rc�(�F�:�5��9��P�����3�!�9u��uXF���|����*�������"|)	P�z,%�$��
}uoed=G��bi������0���´���YS2�ek��բ�>�b�!��J&�WL�	٣:��Г�$������V=��pe\��k�7]��1U��\�{[�s�R�X��6\�m�J6
��=a���w/�������v۾O"d�6�">��u�Y�:޴TGdr��ʒ�*��ߚ<����H�/8�������f�Aa����(���.29���D>�����:�+�̑Q�.���V�T��9�ps��B;>ka��^gykC;<���tu�}2�ש�3������ν6��_Z4�yxIH��X�il6%.Pd�� �p����6���lm�ٮ�wԍȋ
#�<�GLQ�zH�A����e�5���6�7ʗ���s�}9X/38�tg���i�X���*t��.��
�^��ן�a�����"L�c\���2���H�"/d\0#k�3��U�߁N0�J�c%Q�E��ǧ�p��=*b�����g��#|.��ptK�`O��7�����a���K�?qiayON^��횩`�*3=�Z_;���֟���Y4�
"�1Bi'{a�����n�n��#�vOE�ԭFr���F0�F�ͅ�d^E��qN:�J6p�ŀ��>[TDÅ��o�-����9���Zv�6��6��5��K�ph�f�& �Ro�¢ZNX#�DΜ�r�k�vK�����T�T�ʥZ�|�Qʰ�R��E)v�f�ܬ��Q۬��`�H�:�U��v��`��㱵��u>�)�K���;+lcû�с�s�S�m��±���pR9UĽ��Be�.7\g>}	������M�ړLl���G���֜{��ݠk�j«Ð�V��P�X�%G�p�2x��r����zU�ґ�4��XE����W)Ӝ��pE����X���[�7ϗ�\s1u{�Ұ��K��Hǭ�<W+�tV�����+�:o�������b�u1���<�-�y,�-��
��H�]��8�7֎��K��B#Q�ڥ����S��)�0�V�B�62g�6�Q�.TB�;B�(���`��]��SMѲqo=ҕ�r�'���%@�yP�	+b���z�R7.mC�F�ъVj�v�;��j}:��{��G��U�h9�*����C�0��ej\}r���&�{��AGY��;��$�q��nI�IS9Q���Ⱥt��
3��@R�p����Ԗ��M4n�#��ɃB���9P�����ALӁc����Y�t�,��s�Н���$�wF<S}�\�����f1����{E�#���#�ԞŸ)�9[�d��.�ɋEO��.�p������kE�B^���}�3�y��;��e��ސ�t�h3:�pGgk Io9K�6�o�:����б\�}���+P���=yQ�oX��7;��ߚ��ZU���;QT�`��uo�<q�Q��<�:F�n��(�l�w��m6ٗ��W�(�rb�D!LR�U]d��p�e��(j;�h ��
=��r{2fU�Y[["����1uU�m�ם�lb���kǳ�(v�Yu��;-k�ޒ�d�N]A�����&ڄ>��e1P�<���5�_$\15�E��\�J���%��\����|d5��AP[���t*�HѠp���Χ_U�+s:e��.җ���1�TqLy�;Z��q��)i���;P��y$�\�iN�MQ C/��s/rp9���k1�WS�c31a3�fє,P�j�ob��W���]
[�W���7�����D�:Bsx�r�W�!�V� '\�b]ίmj
�Y��;*�싕gϩ]�-w"��{��f_b��,&���V�+�ȝ�<��ZN�6l$�+�D�ۻ�P�-�}���[ɇ�$��|l8�&-���n-)ŝm��S��r'�7+k!E^u��*�6��A�����Y|z��>9�݂jf�N������V>�ھ�.ڸ�\�b1de�$Y��z�&J�ڬMvh1�IP#�|�cer���3$�UkWrI$�I$�I$�]�(v��c��r��R��թa�rwgmc1NStv�Z[)ռ��d�=]g�;���]�w:�*
R�1
an)���s|\�\��G:ݣ����Ma8Ck ޗR����X��os�r����������t��;��-�4g=&��d�*0s���u��8ٴ���yT��#�b�gWzfE\!�[�Y�^͇UΒ+x���S��ލt+�F����C�X\/XA�j[B�&Q���A���!�(�F��SA=��w�#>�R��38�]O�CS�0ѽ\DK7��w7Re�JRڣ�]�=��gIg! �3�pv\o��Sf�-��[�p+��� ��spʏ�Ż�X�	��G&����%Ţuβ�:���d#�<��\�FG��}p�4�_X|�u�fVohr
��^�}��Q.n��ve�������;R��N��K�f���/UZ�b�ᜎ�����b����X��nZ'����E-�3f�&�������L-�R� �6�Xȸd刁��	���v��v-�&酧�ub[WB�\�ڰowdN���hK�$����qe:�}}>[�]ߥa�X٫�N��,�����u_�vI�jK<m�9s;�y�������K�n�˒W�׼��%�ؖ��x�	 �@�U��)m��l��F�R�eV�[R1c|�2�*�*�Z�-l�l��+,T������
%�J�ʨ��7!X��_rc�Z�Z�R�i�-(�jV�R���Uj_0����jVD��TZ�++mkj��R�5Z�ԩTD*YZ��c)Km�Z�+U-jZՌU-�h-Q�
R�S-�W��ڔZ�-,��kZ�PPrʩ���Ѳ���e-mZ��+J�V։AR��Ř�~���k)~�em��Q��TKQ�m�ۓ�m)J�B�E[h��(��ƶ�Tpn5V�#[FQJ7�l(�fLmZ�+���j(�*,Ae�A��r�jPƱQ_�A����F��2T�D�
�R�r�_DšK�b\����L[��ZQ2����Z��eV�5���r�	�j��b[F���[Z�H�[lb���cQD}t�ߞ��MN+����WE@�'��,GW�T�U��T�O��X����ZhWb)q�KJ��eewjK?  ���y��-,��1�K���X=1_��N��W��2"�V^j^ċ�L��w
o�]���rp]��2����{n�"����
2,d���I2���1	�@.F�"8��n3�Wx�c7�Y��u���It�����L>��^ƍ�|L�G�%��2�S��\��j� 圔H���s��î�A��Go�~Un�R�50�U���Gyȷ����Mm�l0��ݕQG�v"�FE��tL%�KC'KBf�(n:�F�F\�O<�����:j��l8�E�m+�7���U�[ ��t�Y��5��\��L.;=���ٺ�c����R3` w#JeH�[����lp]�ǫ#3f�xv�E�l8+׳��*�Ѿ�m��e�h�)��Qq��l2�d-Ud����l.r��m��?9���zHv[��h�Bx��9d��(c�e(���A#��[w�+n&;Ue���N8�n2b��Clu
|�(:�m��jG�������X�M��5#wRvW�	�XQKS�V�*C�r{�<�.�ܦ����)��1M�)|u��#��j@D�Z�=(fʊ�K�:i��ذ>�cfQ���#�Ŕ��Z9]�pn�e�\��
Z��'ga�\��1Wg�"e��[�r��{�з�u��E��������.��g��oLTp(�*���"��8��49mh���R�f�ۨ����E�P�,�`j����p�]�+ڨ��Ti& Y�dm'[���i��Ys0�w�z���ƩV5�D�t.b�s��+A�`���g0c������uu�St��mD18�Y��`i�X�������/���V.�oԥ�H3���-�w4��R�d���������-
̧�@k���V8�91�R�1^Jю�U��?/����Mp�����hJ�"��
�B�!�Q�5�ϱp�Y�(x.�p�:5.����-��ƮC�� b��-u'^�iL5�Ii��|��c���J9�5m���Yuz�Pfs�1"`�^��"'�+����K��bm5���m�
�]R2���<6�1\�6Dw#j�t��}ѬD�Nr"�Fp�>�0t8�^�<V9���l�ף�WzWe*gn%��d1�(��4)�w�
��l���� r���,K�)K�&?i]�Y1;h<B�HI�7n�d�C0�E��O��f�pBM�۪P��b:e��z�%�w�9��e�I�k��q2�v�{p�(t���LR����T�W�Ӻ�vl��i����Ǖ�k��  �=�����JA��`�7���ak��g�5�<=J���yGٴ��ؗn^÷�T��qf�_�����$Oe"6�
|eP�ES���muy|<N�~4�Oz��i�-�;��$S�p/I�F�������J��W���r���kz/�b�+��r%��\�2��!�b�:�J.]U���m_i9�]:^��ǄZ��#E���}����v����vHѥ�[0t�+��<�kι[8��ԩ�t\q��J)9��+��m�ͬ�Vh13����Eq��t��z�qr��2��b��R�݃e�+nG;{,+�b��Tr���F��^s|%"Ǝ�5��W˪��yQ��Ul���5����^�z���4%@���*#;���W ���dϏ/	/Q�"�Q�p?�(-����R<�gv�u�0�e�ЕS����=n���n#!O�����o��S�}(�El����O�Un,����a����"HV���5��g��BLP�^ܥN�>��V�u7\�{���'$�{i���.�Iw��]��������Ծ����b�����Xe��y�޽v��s��yz�u]Q÷�9���-�.��é�K��gD�I�]��v�˔��S��䳰e�r�K>��v��P�`ԑ�����*�R2'Ѵ�3�����3���&ap,��i�����V��8<���	H�����u��lj�ʉ+7�AX)�a�8f(	E�'��U�	�m���z��b�Q���\T�=����{��b)l�	�iS�
�m.��k�:��g0�xa�}�-�|���5�h����q]�E����
	h�ʪ�����f�H��J"_��逕�eN�0a���͖`�JE�-�͚(�s�=C6p��ޙ��_���̑�\!�V��[ȼ"����hj���m�q��͇e��֭�*)�7z�>�S��͖\XU��R5ƛ|�{������&��鬇a�8�ltnE���c�a�Ćh\p#�%3�5<Q�:�ޞp��z�dם�:k �]nJ3B<�S��T0'f��,�<h[�GP�V�,]��G u_b9�-t��KEC��ٶ��ڍ�0��2�_P��&.�Z89��J^\OJ�Ppu|��>�/<��In�4dFI�ױ^�5�c7�B�n��}�ػ�p>A������S&�U�ۉ�6�1Ј��u�6�����'!S�r�w6u�^��id�².=�����t1�pm4�>��Y�ǉ��z����Qҧ}Hr��u%��y^��x��UQF�藰��s|L�\+�ΞPtOq�-|'%�R����dr�ƍ�u|�7�r~�����`�����7g���>�+���(W�0e�f���h\�y�/iՐg�}m!/��i��S%wBN��l��;2,)�K�
8� sb�TWU�Ǖ�r���0&m��7ꇛ6%��A�sƯ��f};�R�>� �������Ovҝ΅�� �B�܈2G:tJx�����>u��?uqt2�WY_3$��r�S���T�*F��Dh5����EFU)J��6^��ZLXoo\�S�LV��K����5 ���ĵ�߄=Ja��Ih�1��p��4����뷷oVr�[[���ɒa�$`9G��BF"�9&$5�ÿ��uH��ʭ�O� ���P�i�V�r�����f��`�b8��m;�63���P�6:pĄ��ɠ\^L�A���U�^*���s8���0ꆑC6�y዁e�ʨ�i�lpq�M������-<��*Wq͠�^zep�e����{t4���W��ޞ|ip�L�u�n��WO�3�ާb�>���"��td0[�kҰn'ݽ1.��7�s��*˭"�k~�C[�[Տ�gf1S#����W[��/J\,���nr�jK?{��3U��0��M��t&9h���J�LU��tw��p��Vz�z0.��Ռ���z�*���ݜ�
��VՂm�����Z��
͖I���#"�ʵ��Yr�g��G]���e��Ԅ���y~����vZ8��ZP�ԴE������+骠��#k�7�ޗ���x�c+L5l�Z/�y�J�N�:�����:2r�xny����d�j^�8�OnWK�E��[��YA�V�,�0P(��U*����u���T��q��d�bU8�oiV8��}PF������;�/A�18����`�5�{s�vN˨�9|�kԏ1(O Wv�^E�_�4��0�	W��WO�CՍdmȩ��=em��@7�����gM�ˇv��_˖�0/
a�upc�����\'��~4�+�%��]3�ZN�t���J����H{}aDZ�3 [��r��_�]q��NAhp�F�δ�����W)�v�U�>V���|x����DR���"B��S�|%S�l�
�c�����f�G���7�У����B���������s-����u�Vb�F��$������f�]:�H�w�%C�ćrj�NX0��DY���;ʺJ��v�T^�֜���L���#��vǝ���Oo��i���%&�oU��Ө̡���r]����7���8�y�N�^�F��8b|���K8 �$c ��r��Bb��i��*�ܽP����z�(�P%�\���A����",4U�Z��G���>;M��Q̊���"};-����׍y�?9ƥzۯ	��ꕪ����4���g�jŹ^�AP�L{*_�������c�ULb+�+���yN��m����Vv��W��&�G^k|�uB����&���`�p�!�|&tᡸ�M�J��,�cg$׺,�i�AvfϤ�N����Ҹ[J���qǏeN �Dc�Ps#H�U����D����\<K�&�]�f<�]Q}6�Cdod��>��� |�)���5�+ӵA���(��H�z��f���y3'8,k����(���@:�#��K�8e�x-��%F���T��<k�Kn1;p�M��1M4dub�@b�q��,�ʙ�9�ر���7s�O�
��0�֠�R�T��^��a�4�{!}8��t�\C"p��������
vi&"	T��+B�� �!�@�e'��.��f��9 �J��n���`�M:g(\�}yy����'��%RMj����H�}��N�*�7z&uj��({���s2�3mD��K�ԉ���������ԗ|��gm�i=��٤Kt���2��>��|<7�� A�z��VF�ꃡv���8�j7������
`#Cf\F?@��1\z�D�������^��f&���'�E{�'f*���/�تR�H�C!��ל�xM:]�ɇ����[�l�{�΄�,���FI�ѥҪ�
裠���"��b\�![���T�d̳����1�n<����.�b���<����E�n�uX��a��V�P�F��v��vM���yV���j�4n&{�V�fV
�y?VB5��H���!QN��1����ϖ�Bf�u-n�v�`�z���4C�q�*Q�YS�M8y�L�ࠑ��/D>X�GA;f����&L���y���Q�{�"�X>�+��IT��p�\��P��,�d�e�$+77��0���dU�+
�J�jZ�1�{I�#6��#w���t����(��r��H�~�[Szx�x��XZ�u�ha�imnE58�����Bѯp>�5ȫa��:@�MmJ��ٹ�&Ӭىě�
�+*d}T˚��Q���r8����so��B���g�l�8�-�}��w7xM����oP��Ď\\����[]O�#Й)��y�1��8�8�)����Fw[X�s����������D���"����ll2�J-@�W4�H��9�\��5F�N:���z-"㫼µ�۸�l穮5lH�\0Gd&c|F�P��=8�
p����٫��!d���5��N��������x�B؞6���2R00���c��b���&F�i�,��	�b�%���!�ޑ;�$��LOl2�8QFȳƆ)W^�\D��UU�O�SQ����6��f��w	���΅p$��:�Z�F��6��n�k]I�������|���y�G޹�%v�Y�`�1�D������q'>TK�ٻ2%!�wë�x���L���3iS9Q��Y�jC1�H(�!$����N��jlV��Da�|�C��'�}z���~5�żgk�4dU:fq�ژrn.L,��r(�쥄�!�5�<�n�~3ŷ�Vb�Բ��{�����f!=���rÙy�Uy��C��߄��&����-Q^8Q�rc��&anxƳ�Bo¸�f�>-����K�ksz��w邝v&��=��x�'&��&��0��ن�����i�=�ąK��
�?fA��Z��_ϣ����o��"m�L&NJ�Z�*��nnl��"��F����0Y�p��mAn������K��W�{^>cs�G��9*���į�S~h�>'��>TW���8F�q.v��3�[|����p0"�N�@�*Y$SFnLP�$Ć��aA��2Zڧ�W>Z�����HVq���8�p�B��J�QG�3�ёfk��0�`�hd�{{���w��u�1�L}Ҿ��2/j��1��ݕQ��'[�͜4u��Q-g!�|:��cj���G���.�������t��WP���3aP�[����l9�L�Mq�yJ҄��j��*���ew
� ^ΛyU��:�����J�����3O_��M1Wϥs�3nE�ud��P��,�[<�v_��3�ަөhu9x��X�E3-e�Mҕ��^�:*FڔUYl�Q-G�Ɋv��C�,:��<\�k/035w]�dL��/��tg�3E�"�*�E�w]{0��w�J0B�`�J[�A�!:I������:��%�D#�-�k�ug��"m�Z.ᗦt��DF��;j.�-���0�\�n��j��/[��_��m�8���YΞWr�l��د2�;x�I ]nڦ�/o����ڸޕn�+}C�nokh-]Զp����w�����MF�wZ��8*��]-�hw{c��4K�!Õ�D(��o)��e	2_vS��7�|�3}��5�f���Q�y�tTUWJV]����Ȭۍ�LB�մ^5ʍgL���k���p����
��B�>-.*Qځ���wMe=�
�)P �|��+y]�.'��Q��1�W�&y��X���>n��`e���о��u�/T+%��4��Lq�og��T�S����;����\2Ά��nY֢SlՂM^�z��d	۹����mlb�9��ܨ�&�jL��Y���WjC��FY#Jˬ=Ձ���os���Kq��K��Z� �O���3�LCV2I�b���aMھ{5�E((���ɦ� �f�n�:)ݪ��z�G����z�V��ٷ&n��<"au�al��5;x�qۡX�,�;�Xi���f�t��N�X+np3Z�Q��qL��<���6���l���i�4.ٵ�)��fLo-N�jX�����Is��[3���1f&,s*$�U��� ��jp��Wmo�K��V{��wY)]L}K[�������:�F��.d�h��W��1�={�֒I$�I$�K������}�K{t�g��)w�ޢ�z��l�f���Kt�%Ճ1Of�$���I�o�,(��b��ѹ]���\I��h�l��X��ec�列�'�%S��MØ����L��U�̈EuLŻ=n������% ��Г�7ԁ��{��\'�`:��ɐN�{G�^��tm���3���#M�s�:�	�..��e��YS�P0r�7���#D3��r���r���ߊ0l��bΚ�M�����ֵ�.V���>��e_q�O0��m�W�&'����,+��co������h��ϻF�R��ϣ?1�H?���n���Z_�I2�"����{e��G�CH">l�.<�Xic]��@����1%e�ҋp�k`�S�UY�Uu��	#�7��av���:~���D���9ێ/�go�
v��ۙXl��ո���((����w�Y���f��� ��a���^_.+Xz�^՚��C��l Z�}�ak���&m`q�yVhWj|%����_L�Fm���w>Ƶ�&�������F��Ȩ �m8�5�ۨ`�gfު3~��Q���WV��ڋ�q�C�of�s:�b��
�n��U����-�P��8)�vF�ol����v�+� mj��s2h��헳/�έ��g+�/zԞSw��x��wH���r��9s;9>�ntno$�+Ė_r\��޽K�r[��jI~��V�[j+jk(�U��մE6ж��[,A��TX*�Kj?��5��02��(�b85�oԱ"�(���T��J�m�����y��3(�c�,���Xڊł�s*,PZ�*�TYjV(��$[J�ڢ��Y�TT��1A�V-A�YՊ*��Tm��k(��SYL-���6�Z���Xa�*n�(�ZZ�B��*�FU�PQGV�V$b��-X#��
�ʭ��
���Tm�E�[R�V���������hZ#iid��,��Z�q�Qӈ�lV�-m���#Z�TD�ݘ�nѭ��f]e�ahq�E��
�� 6��֊��ڞZ"	n�*V[Eb#"�)PʔQZ[R�*��"�TYkJ��D[l������V1J��2֔J�4ŵQ7� ����m>��Ƅm�0�cTmH:8�Lu�a�eF�P����X����X�������F�i�R�{c����Wo�R[����]o5�*A�P��54���:�
zkc���|�Mȩ��n%��g�SGo��MLv%�`��3|#`�<!��0����c>����x?��O*j\�ǂ4���g<��,x��u��/��E�,��'�(K�3�~�0i�)��mа��?P^��:��[��X����PȀaC1	���F�"�JaE
s�h^�62��\i��W�V�*˒z,�6e�8b6x3`�p�R���%	������F���o��[�-�S&_��"������Tu$B,k�;،[8f(K,��`�!�M����j-.vt��Bse�˃��Y˩F&�[�aePgM�!��;X�4S�NW�Z
�����l>�r�$>�2��6r�)�62�3{�LF�a�1�<�;u;.��|�^u_A����|V�ª��WJ�/����ݰ�^�.a�6Yb��I2�Z�U�9��%�5�"�Uϳi���9k�K�,�C��X�\E(�De7\leJsL��V�U�@�ʕ��%�Z--uQCh�( y�t��&���q����^tq�|8��m�і�d��4<T:�����u��V_8|\�57q#�ۜ٬{o�]'\պ�{��X)w���	w��;�X�9Bz���I�?UW�_'r�Q][j�ݚ��>�nQqc��X[�F����������^fdN�0��p�5Q�3�l%)�Q�gK���Y���V�ƶ��>u��3�QQ��}����ǟn5�'3�]�B ��YL��(�P��<Yx�3������Pvi�W��F�כ(;�:rn��%G3�\ApL.0t�rWӀ.2 �2C���5Hһ姝U�Dk蠢3�J=�BP4!�� �,еT���<U����������n���{��[X[��-Hw"m�B��)P��D\)f�f�(��4��m���ttB,8��Qg.��Yj���dh����:`W�udE��A�Y�p�SWu����$=�����{�KS4�.�8Ru�E�v�\!�&,��t��k�
�W�f{�h�K�N�,�G%�6	>�v"+i�f��`6S�3Nٍ;����+8���lڽ�,����3�xj.b�����r""w���s`��[������ \�Q��N�Z��kv����dLrg�l�t���u<��a�H�0��'sڗfuEI�IF���4���d�V-��GU�2$���(=���!FIH&��&��+��b/i��۰c�|��'��0k�{g�� >�fM�Ó%H�C:G5�Q��b�R�t�M��ZfP�f6��� *�鬅�q����D���Wa����p#�#�B�}1}B��$@[Ub9�;\��gPB��xb�F�'�	C�����]%R� ~/�}����<hn��[Ü�S���8 Wl�c���\�T�S$>�rP���K,U��.D�wՁ�͓�����mU��.�o˩�U��x�YkNo�8��t��%���~>�-������c��"�*��q��z{��x����gf�k���:�ׯ^�X����8M�Z>�[|�NP��Gzm�2�=]2���o����s��*��I	��&�Gz؞4-�#�d�b��q�*hwe�M#��S�r�YU�b9l��E:��썟&.���(��x�<�TgKm�����B��p�K����z]�}p�9@�t9j��7Ì�����l�`�UM����&L��1R͑^�/#�u@U;�b�qh�ҴY�:���Ф|�Ŕ�_+l3P*�n���u��s:�s�}(U�����wE�+Sǀ�(<�7�{����$�ePU׏]qٖ�OQ������Sm��RS���Z�-��B�k������s�u&w*jc�g���<|/��uKʥϫ���xFp54dPR��D.)թ����=g:B*4��Hgي�eX������'ƴerOƦ�I��N�V�v���$���fdX��K	-TDf�1�G˄�ps�|_W�a*��
�V]�a�!�k����7J@�ʣbB�`�,���'D�Ir�X��}(�;- ���8��jp�{{'��=�Y*�r" _�x�K���^�Y�|����X��m�jN��z�f����v�b$�C���((d�o�ܘ�N����A�*Ml�^J��Pq����f�ea��X�B(��pmq�d���
�����fYo{o<�TI�����ΑyeDU����!���H6ᎁeϤ���U���wǃ=�ĕ��7H]�Oy�$н�QO��VXϪ;�Z��3*��:g)��6p�zE�E��#;���e���z�ã��)C��ǫ#(>�1`�K:��<�A�x� ���+���-�����`�O�m�9=oYyٷ�<�1^�9�?z����O�H&��Y�gU��z�������2ʫ(��[���U/�)��kE�~��⛴�s��Ų7�D�U���k�]��dY��
鵳a���"؇f���WT�y7ܻ���^��m�s.h��I`�R�Μ�f5+��o��1��0�u-�r�=�*WeֹZ ���$�R�lB}\kgOӔ���q��:#��4
b���q)��w���Z�=�i�"��r���qōr͛��Eۮ�Y�=[0��a9�Q�3��^�E+fa\��{6�������Pq!�Gw�X�tέtH�y���Ze��1�X�S�ϡ�	��a�)D,�8�:t�B!^��Ի�*z�u@x�YH��\ƓW-e��f������_ϯ�P�O}Ap�P:x<k�Қ��)�Q;t)8'�)�m,y�
��]A�u:A��Ъ��֒���x;�-%�-
��=pn�\2�y��fU�=]:zZU�u��+�J�e�`;JY*Y��%�{�i>��l��	h�N�����}��ٓ�Z����4Q�;Lg�3��f�3*\D!2pk$,}����;Q~��&\)(k���l�� '��A<	�D[Fp�T�ȯ֢���P֌�����:nI�>{�U�z�C3���Bj=���wo���CImY���3�بF���͈kW��1=��]xy/wl��0nT�+W!vM�+������;�;"9���%��:������˨Y�褎>����i�?I՞��Q�V3���Jk���<ju�^�d=B������:L9�J1��fM�t�1��+D~׀��
��U��Ju��`�N�ۆ��d1C�Y[b��gwUu䘑�x˗�R���b�*؆
�Õ��+�a<>۶�׵�:��~�Lmʣ��ǹﻭ� ������|�����"�U���{+�E��;B�������+%��C[�ۮ�MT̘�XΖz"����XF��s|��G|�+V��`�@��߀��ܨNuVNd�"eRJ=�ҎX(�Yw�6�VUi����ڦ�<6��V�:�A��T�=���:�E=�Z,w��wωu|����h\��g�2�܌��.U�q/=����,��:]@x�t��?�Dq�\h+$�Se(��Zd9Т&���+|��ެ��0{�裷�U�������.8�`Qf���lLQ��=p�e���ѷ7����9��B���P�S:e�P�!b��<r"�
|$�r�V�ΊNH��1���kݬU�N���Q��wu�6�2!�������c�Vsg��8�E�2�;��^@xǓb�U��W�:R�-��u�1�SF&��K=��U�3�U԰�;2I���R��Vb]�B���TNo:X���]h=n`�-��s��S⯱�wK��3b:��Ki��� �vi���;lQ��A�z�t���}����:-�e��/i<�01�W��N|"��xS�|kʟ1`��v�$���D�d�KX]^ZNG	�����nx�iB����*F)Ȓ�wLO*���3�J�j��ة�ɒ�����l�3c`�21�ȯGu�\Ń�8�13�U������q�M�N��9ǁ��ѧ���uIi:���1�<����F�Ɖ������o����e(��-��������B�����
�X~��b�Q���5��N��=i��H�Ax�����Єv+��eX���Ue^77���D��B`�:;J���R� T����ujW9��7Lo���Z�W�(AՕ�K�ڢ&���W9�:���}��l��A�<硋4�o�B�яI\5���+6h�oےˋU�חS��{C���G'\ezhCM���l[�����NGє5C���o�S�~>�/=T�r�p���"��n�=듸��C�,�8�yQ��)6�
��M��
�5V�5���Lǵ
��]Z�J�����ڿj�7U�7��160������q9���qS�uj[��'�><i���'vZ����Fgw\�a�Ԭ��E��d��_A�N�2�D=�Y��wh!KN�K����2��%��3��ӦS���1���9Ur�Jڻ��o��x�SOp)<���ą��\����s��bZ�7�/�p8d")�t7�OdC�6;�g�5n��*!HCM�Tx�ۑow���DA��oO*�{�HvN�J���pȞB��nzQ�rRgd[О��1=0��#F��]|�U��<�G���=�Cp����*�p#{���Hnu��km�m��Ѹ����S��:_���0�w��/�*g*0[UfE��3rH���#�6�py�`����D�v��� �j���ʹq���LӁ|��5�َKݗ}�����U�\�	�q-r�#5�.A�ۊ�d~u��y2�*�o9]�ֻ��U�-
�.��f#t�p#ԽM�JBa�:�����J+ժ�I��˳��^ ,>���PHPu��X-D�9����,�!7���-�|�Q��G�K}ט/˲��72nK�4����T�
�
�Iћ�9Ɉ��A�Rk���b�v^J�|��(�����GɄM�f���貸�\4%��f�qQ�=]N���o�X�9y�c����m�.��T�aw[nncc�r��')��[s�@w[�í9:�H5K��;��w\��Ζ,���~��m��~�����l��,�j�7�K�T����Y�r"Z2,�9&!�l���$�ں��=>�J���k���]pv��k�O~Y���2�ё��@��eTQ����\ȇ����u}��e�L���&���ʝ5V�62��^���:��*�ݧ���'�G���yI�]Gl<��"2��PocM=��F�hO�,�d����>���t�X�o`��h0A<�^�n/bު�9�C�zn2cj-¬��>ޫ�/;�,̎�{;�/9+�ftsot-'=/��̤8Aӳwà=�g�Z>�\��u���eW8�bv��E2�,�l�g��p'ˉ�3�痄�.�u��9�م��0P(�0ٻQ��Zh�T����X4Ҧ�hu�UtB:��c�s�r�H{ҏ9u��jr�R����~��;�ۏ>�!<2Q�,��(�;(Mp�K��1\��ά\Zy��_=��3m!��ht��q=�)�5�~�q���<r,�!�upt1�O��9���XgZ�]&c�ge��t�g��*��/i�{�<���i�[��G��e�*i�j��%		���a�g5�swy/]�+,���+�-Ʀ�l�;Gư̳v��n�4����_g^	�����S�����$M����]���o6qv:n�,&�T�s�����U.U��{�.�Դ�T��++�C�\8��rG��5�bg��km`^:δ��<<-Q��Dĩf!��4+��Jc"值p�{��;�$z��{ ϑ����`�p�l�V,�6�p��1���r/|݅tOF������â��%��^W6�P%F�1P�9�
8'Y�0"�/g��N߆���w�{�8W�9�Fr����7�Mp*�����x`��:�t<n��e��슰f���J\��%�tnz��Eh�z���rZ|0�O�pA^��/$L���ח>�z��z�������;J�ނ`��0C7��L��[���ʔ��R�[�����֞8x�^��ݪ�j��wޗYhy�+=+H�E��?"Uׯ��M��ū%a+(�WLTEf�.,*�'y����
z뺧<�t�`���h����Bqn.�
v�G1�X#dWR��[��<�[��,絵|q���Ժi���m՜T���m+�Qf�|�Z8vG�9CWf�+)a���ً�5� `rb+Z;��ݷ��޹Lu��Ma�	�hMQʐn8/ ���A��]�ݛ*�b�9�k�Ft �T���2�]1 ,���n�98��\���̮�Q��Эe��y��.���NS�w�[;V�ռ#�5}�pɪ�,r��cf������(2��wԆ��;�2�Z�>W6�&z��	�uو��ax�*n7�����%;g�/%�݌w#F����Y�c&�ӽ+��9H�����)@���0,쩿\	w��vY�Y�mk!xDb��W׫�Z�A̞]I�"���D�%�hɒU�U�\�źs{��{;.՘Ցt�8+F,e�֧\�����FW�7��ۣ�L�޷��yI������TNS8��(h����@�JK����D�ڑ��g ��uFػ�gG�1ݳ3�2����X�D�t(�n��mX�!��C�3�5�ms�N��l��n_^��I.��8�xrɎ':�gZ���|I~V7Q�0VqF�ۗ;�`c��3�U�|���i,w�v���+`�,��r���>roT	6R��7.=Mgk�W�3�]�դ�T�� U����(u�^����c�!P��ͻ�96��nZ�O��|ͭZ�񩑀���fN��}yt�k驈^n�&T��p��ΔK���j�K4��vdo�wwwwrI$�I%W+����UUx�͋���� iYϤ��M#Uf7\G*cw���������{��	9�^�[F��~�<u �_w�o���r�����:��j0M��y�>'cs1j9@s����y�3�m�fĺU�/��x�0���V�Հ�)�}+Eb:�^MWw����J�PT�SmEW[N�Zs%.��)q#]��R 2Ċ˔��C
�W�x+ ǎ1ν˗5�䡜��`����l$�0�m��
ٓBU��#�@�U
��Y֏.p%�vCf
�% �p��Q2��;B�ܔL�T@Āj�x,h�ZX�b��2*p�v��8��\����Jr]7�H*mh�1���t����:XR����8������DD�U�����k0�����h5���.�s:!mf�$��H�Vb��G���d(�ya�T7�#%B}��[	}�7A�d���䉑�ц��nte�ڵ�~6)�}Z�4)�ݚ�PW�D�7+5�qm��7Bn}�&�'��rI9Q�8���fn�vmvԱ�]�j�cFݼ���"��9Zh�{83�7}Lj� |1MI��W/���E���}7�\����{M�o9����uM�9ogl�nr���Ѹ���|��);�w4�>��>Ns���:2����\��D�ڣ���_P��+�(Q�je*�Y�b�%f""�-X�J2�H�TA-���0�Ɋɶ���X�e��m�V�UDDU�*��U�ƈ�.�����c1�U�m�)�&.U�_i,յ��ۦbQ�%T1�Qb*��e��j+IV����+��4���SƬP�B�e`��0�����TK4�& ,]�e���M��ij��jZ�LV+w�Y�\`�E��M&���Zl�ӊ
J�D�.�̨���KhŴ�&;L�j��,Z+-Q���ӂ��4���BiG��ib�"b�-�ISj�E�����(,�Z������)kKjԢi��%Je*��1j�Ud\���,��a�x�VlZX�)�r�7*��ˉ��r��=�t�(���4���3Z�����%�6�)�[r�T�f"H�s�8ۤ��W/�3[������ں��4�gQ�7�uȂ�\)�v��WpjO2iR�2v�;ʷ9!���3���ntw_j�'��D@\:���n�����z��s�����g��<��6W�B��sX"��$q�
fd�Q#näY�r�OR�*��^&��waj����C],�t\i��%�\q����d�4%q��@v��B*�d�M�ȋU�6y̵�h=+ck8�X�]�!鑱�e�"8x�X1(�je���}�v���o���/��>_zI�
X�*08P��a��'A�R�D_�K7,!f^(B�W,.x��=Y�l���(2V�8_rv[�F�B#�<�GL�����^���3��\��v��=W���ᬦaF��E8�8�2*F-piK����nAя\�
�LR�d�f\2���v�l�3����A�n�uXU�Ԉy��`��d�(,�|5����xj;SJ��x�F�Ɖ&�R���)Q����n�H��c��+"�ƉC��K�?�P��5��k�	�z'�?C�ڼ�s��m�MsSYD�����P��dCQ�F`�Xa��sad�j9C���'VX6��Y��w7�Yv�E^�Wյ�:s�֯���U���rz�5����Έ��S���z��Ӥ�;��`3�+���ơK����7�1bO�U�s��(_}=���pz�s����}�[��w��Tw��.?���J��X�\��"kܩ�a���S�6"|�ID�fWy9���1S\`���\I��4P7��EŪ��u;�{"�Kk,���= ���J���k��ݽK��d�wݷ�vcE�#�e��p��3e�X��~(y��Vg��Q<�=E<Ƥ-��Ց\����G��1�;T�6�6
t���P!8P��=}*�s���ً��_��C�^�Y}�,=t6l;�:7��9����:<2��hs�
�k�!���;K%gKޥEf��Y��yڎÕ�nB��oH���sG��(ۙD%J�V��x��˭i�L�%l@��E�W��JB.�N�J��z"�Cr'��"���s��u�[��n�Cu�C5,���k�|z�Dwӱ�*���H���
��_%�9�M'n����=*꣊@a9�j\����9�3Ʀ>�B���ٹ�p*�ݰ<��Y{Թ���!&� �Y�I��ːk�l��M[���~5a�+Q�n�;�C<�Z ��]��nWr�e��A&�|�Ŝ.��Q��e.G.��r�䳏h�7����0����y(o�둷<gX�wE\^�lukYjd;ٌ�١��V2�r	�����rI�s�jv��{��<�ꝃc}˿-�װ����kz��J�ȸ��9�?�R�_˕ 1�ǂ�hX:}��a��o��3���zx��"}g�c�ά�R�$K�`��S6P7��8�%OLP8Q�1�k�El��ۭV\��m�$ʊ�T�,0�P9�Ɋj\EO�R!+��>�h�&�ꕫ��3jjy��U�*Q��i�0D�)I.{�0b��I3rb�9&$5��2҅��׷]�w�횘ȸr��S�EOŎ��n0�K�Wl��8������3 ���B5��f;o���B�a�wMw�/=3y��ClePdVVݠp�+�Pz��ӃG/�L�L�#^����]��>�A��)��v=���]O&t߲��Y�5��3�#�2MŊ,���ֻ�l��ZM�8Ut��Վ���
�{i�V�4�<hr�ym�R��9��m�W�ef0��X�<�]�ߟr��N��N}J+�Qn2�h�Su��׭��m��FI|��;e�Y�,�S�PU����q���T�]2���xC<��EX+qx�'�rp��w�>���$C�ʶ͞^a�C�-�q|q�	q��e=cxs��ܓgN�,lT�J���d������ݘ���*㬊�0�t�ϵ��!�v#����Wh�.�H���w�%r�HkH2t}ܿ|��������2��m�GT(�k��X�(�}ҋ��8{��ً�n�˥ſT-nn�EGXw�*X!��SNhuʮ�FƩ��YՁ��&���u��v�'�q�%�)�梙������gЖ ��5����]tu�Vr�fԓ�m������_1V�`�1tP��.b{��f~�q�荗<r,�"�GJh3 ���)û\��4����Άz܌J�I�J]ĉRC~�X�'�*\��9�b�J1�w�!�v��#ݢ54�V=�_�ݺa��O=�<8Z����"�8�Bd+
Q�����oۭ�V��_da�wG���6
�T���p�jT�ǯs�fS\���{�0s��7�zg�f\9��dW��O��!>^��8򄖨�ђb�ʒ�[���<�0D�r`�B8Uiy�����+�y?u��xL6�V�/��Ql�|���oOSr];�&@tng�\3�C5eix&l�d��FS�o-?Q��V�be{�20�q�ڮ<� �z���տ,�s:Y�ʳ)Zse����k{1� �%�y2Z��w�������SO��X\�۰ďh�ݛܝs�ݦ��I���n������B�K��;���]qa��\����l�ue�ǐ2�V�[�w�3������XE��G~���k���R�9P��К'ٰ�,�Ѹ�O�B��cX�t��fmV��k��0y�}�Mt�9~���u�H�:�4!W�׬�+��p�G-�u�"!�n���<l2�3a��>״��5oa�v*�S;����Yq�׮rh9��f�C���x�*`��J"��ͻ�t�����:ڭ/5�c#����|�,�շ��
�iW�TTi���1�R8�L����]_.�>���^�$��Ǌ�&7UUv�^Ň��3�%�
��%�60	���#�zW�]"6�����>{�	��ƹ�[t���)t� 9s��
e������͇BP5x#��xo]���XR�œ<u��w'�`T��#���]Pfֻʌ�2�/�߾u�ǖ�'���;xz]oqSL�eL�ba�6Q�3�nT��3EJkb��#r!���~��^l���]`��)f��������ݒ<xր�����f��͈Q���p�QGA��aQgZp�������@O7�*�|6baSz�4-c�ރsD�q�Y���3���AZ�L����A��F�mM��������j����M�=�n��㩉s��_
r�l��=����|�ۖ�ul�ۑ����S�ZwS�]��Ȓ^��_�z2hT3�giB���83�t2(F�p˽Z'f��힫����]M(��T�a�p/��3���p���E�L\xߋ�f���j,o6ng��'�夷�����
`���ᘡ(�|���E
�5����*w�x�Aw�9Ҧ�Fs�]ݽ�qj�i�E�LP���U{�k
'�"�`�:;J��4�x��QX�a]t��h�9��X�E�,��Ir�49S���ʗ^� �z!��v�Z�O��Cr�za ����⽛4P;p��U����6���7����Wr�5�@sp�);]������4r��s^��Ũ�*��8=p�꺤��5�(�Seꑮ4���ةǻ}'�=8�#����{�i`�7c&6ؑ�.#�Bf$�p��.�b�Rh^x�sG2�-嵜t��9��K%o�L2�jb�=KC�@V�"�V��u�����Z�'�qa�hTM���2�N�Ey�t7�OdC�6:g�6<1��L9�2�WN�ї�e��\�6N���L5&���v�PMb�kn�r]غ��R��wa��,���=�*�.���-��s���P�)�*��c��w��zN�˦m��k���Wp�0,��r����{��{���?J��Nв��U������SY�=�$8C��S-��e�ԧn(;(ժ�o���<�GEeR��bw���Dp!�r�l7r��*-���,غXy�}cTz�혟Q>����	KT�����Y�W���S9P����Y�����R���ѐ�]U���(pS��`ʢ�x���*�2p��|i��J�>>�%y���uc���0ڻ���Vd_��1B3ա;R���>\M
�]�D��i��ǲ�9F:���"7Ϋ���"�*�!�>�|'Q�|N�*�\�����G7I����b"�� ]�-�b��P2�`ܘ�Ң(	�F���A���X���k��F�ڇ�["&�2$�.3IB�����\T�HW&8rI��u�ee���g[}[؎O��fH��?*�>/MF}�vP�=@v��,*��ɇ=�޹�l�D����	X/�`1#�.�Hm��6܌�A�C6�y዁e͋�b$���G�a�Q�7� �꒡e�;z�*�)�����Տw$zTA֡$���-���W�������ؽ~����q�K9���o��ƫw��_`$�U`�D�P�R9��uʬ�SӨp�t9��(!�Ef�K��^-�oZ;��*(�7��Ox���q�au�F�-��X�l鼦(P�0T�n��ގ�����*�蒬�H��<�Q��ތ]�ǩ��/C�Pf�t�ʭ4kք�����!��-r��3���d���لQjq����ٿ��uN7�a`�M��cj5å(¡z�9��>�j����.9�E��d��+�)l�Qr��cK-�LS��o^le\K����"b��*�	Yb���e�5nTB7�qŁ�Y�oea�Z,��l�7*�'%��n�=����A��2t@p�X>�Ď�U�R�q^�,�`j��ȅ��0���Cmn]�.ᕦt�) ���*4�qU逍K���T���W�34Ȋy�i��LZܱ��<���"�N󨌧尭�/����f��ODT��fQOB3�T���K���s�:=����Ŏ�T���bM�u-HQ��b\EK�3��{KB[�;{�M)�rx�s!I�GL�� ^E�8b�ҴYfpF��� U,�JASH�2���D�jQykb�oT�]������c�����@'<��Cӣz	u�w�q�dB�R�J��%)�H��x*���-u>�����k�4-^�F�	�v�s,�oCM��G��
���{2VwJ��&cn�9���˞\��~3{)a:?V+(�����ax]tg�b��r� �l�g1O}�,��]B#�-�I�8D���od(���P�S!��"�_��N`�B,jq�����殹�O�B���^�=l�v����[x�<"v�し2���AWa��R#,du�+�ӳ �1�z"O8��	Õo������6r�e#��2y)���'2j�����e��p,B�e�?f�.�2e҂��	ά�T<>%�m
��>Ƚ��Fv�F�%���V�,g�$����T��]OzX�ӷSe���\:hDl%<�}D������c*X4l��7��	�#^�W�yz{$99��ى���$��`֔t�b4�'��c�(�F����J��n�3�e�l�clޖ:��V�7���U��L��R�*�=5�,	�"i	k�3�ةDW�J8۩yr��>�;z���N��у�읰.��R�fú.8��.4؈�׮d����0S����y]\�ĖxQį��u�z��2���)�����B��y6���OsS������Vs����;�{�C*�՚��[��^���=]s�Z[��3:v�q��ݓo��ӈ�n��+WR���z�Ϣ-��!j��b���K�.��Y��F����;jqr����ȇ�6"�s
���.8¾�íO�q����3�s�d�D�y���!���]Pmk��d)��{�\F?@V��'�F�fȮX���G��4H������j��|�À�c3T���P�Ȏ@dv	��M��.	Yݭ��^�Oυl@��q!Op΁u�;�7�2��:���N�株":�6�S���<d:�F(t�!ړ�ꞌ�g��1p�<1�L RW�Vo��Y%xA��J�U�c3UWG���
F0�R~.a��j�%�������.���d��W���-9���k�3ZJ�WOJu��b��"��2��h�p6�&��p,M�oI��t�qs'�;&�t�(E���	�%OLXjc"b(�`��/��L���L�$u��^��g��0�dYFz0�E��,��Io�2E����ڜ�S.���3};MTˎK�_�ǩ#0m�*��R{����@߷%
l�]N�=��L����K��}^�0$�^"E��xE�u`0�n*�8�|Vur��.dE�>]ݚ�
�������>�F S�ͮ�[u#+��M��	4��$Ǳ������)�1�~Go=S�̹c�C&Wqy���k��'
J���gA��T�Y��й)2� R�l*��f�Z�vq�S&G�	����ؼ��0�
�����D(�V�4[���v�o*�6�{�MZ|���X�CZ�%��J?[�4q��z��:K�+lw��m�$-�8�}�oc��b�iJ��j�I�R�O)M��Vʹ1魐��aK�l7yݗ���{�S�wj�ѨN����}��i�"nbB���^�l��K����&O�v��ܰҾrE�a��\�O(�!���m�thJ5.�f��4�.�2%���.E���yR�KR�0dCCוh��\�eGjn9u�J�l<js�ri}f�̎ܬ]s)Ӄ��O7C�xt� xSy������k
�R��i�0���2����+r󥮀����i*����ΤK�
�[vs$�Li���dCkV}���{v3��<��i0~��%�l͵��G�X�n�+nC�4NV���tW�е\j˘�.���a:(Џ��
Q��+/vQ �d�o�=Ƭ^,�/@Ա��\m�F�:Pa�B�=�8C�0u]���tE�8��M��3�X��j+�ڋE>{ƒ�zb�א�Рu@[�I�[h/F���ԒI$�I$�I*�گOY]��:A���:n�ڶ{Ժ�:���ǉRӍU�7+uF�y/Y��rzw#b0SU�����2���)x�'�������qQ�en�`� '9˙@��I5T��[i�˨��2�)}��E��
5P�nnw}/)3�f'��X���&�v���*bH:��n+�XR�S+ ��:T��A�B˃(�5�R���ɺ0�ԩ����t�F��η��`��>;`Y�.�T-#���E�3]�1��H��V^�r7)՟��cp�UfP��%��^��%�;o&hSt����L�n�M��+�1�5�k �����
�]���e`ۂP�b�
�}#;���'�K�7t���T����?[P�v��<.�]̛�����ݻV��f�H�@���kj��Sp�:s�7�d�@*x26��z��b�l�dImKp��\��d*�
�b�
�Y�ӝW����5[�@�k�1���U7Y]}P��՛F당�1D�"�lY��W9��/8j9���8�y��n�DWX�eAͽ|ᮻ���[n�������j�)R��A�ӳ��_T��1�"�oR��9���|��9<սq�3�s�l!�3��NN�9s������˓��Ϥ�}ϻ����V#s�������8�u������0�(�7�40���*b�3T�mWv��Z3z֦�Z�*�3tp�Kmb�T�q��S�v�LQ�e��W{��bkVb�Ȼs,�����Qse7�q|��%����ՙ��mT�(�4:�t�f����>�f�!��[�iU���e�ӤK���]f�E%q����V�VQ�A\�ְOub!��UTr�[Cn�m(��d��]&[

,AU�]Q�3c���uj�n65(�3�j6&�}ޕU�i2��-�㬩hXj�-*"e�E�D��6�Ȣ�Z�SC-|sT�eX��A�b��N9l�9pM4A�TQ
�(�&�AEU��\u�̨���(�)���:�#���
:��Z'�Օ���]�K;����%K����D����ܳ���e�X�NS��E /�K��bΊ��U�"-|/�U���.�_V��}1�p�E��i�&Mޫ��Q�Y���@��,͔T)��FM5�k�n�=��mŖ)�)gV�Wr�~��p�}�7=N�:��V���K��Ys}=���� �J<p�a�jb(���]�wxt��&�,OM�3Ś�񍐧�eMꘗ���%��0t��R�U�#�U6�2:
�_������o-\�Pc�^�fo�f��U��.TB��e�\<���n'v%F�=N!�x��ìܬ�˕J�P,D<���S6�Q����dP��9��5����U	Y�w����]�i+�畓�W�o�L>���R���;��5��x�[�zb򩓺c�˵ϞWR����]��wάȰ�3䂍���Gl�(��Duo�i�y�37�ؽ�+fs���f*���ʫP0��2w�
�������N.TF�5�0���w�Rφ5��>nz��+}RӋ�T6"��Ù�q�{,R�`��S6
���斛�3w%�v�QN�4���6���2�ذ)ty2l��{3t�C�����zoX쮊�8c��
8�hs��S�y�������6^T3G�]3�9�C�,���m��ͩ�J��(�\��##�L�U(Z����x_̷ٝpĵ�ԥ�'9ܿ|�����qD�I��e��Á�+EY�\�W�1a߁N�~Qf��5."�
�m֜t��:�U�ެ�o�I`�1�Qy(�4Y��%
RK���d�A�7&#��3�\Ʈ\��ZL03c����v�J~T�:>��8�G~�y/@�)n�6IԹO�8r���h�ZEd�y��*�������2���p�ٞ��6ݨ��Lj� ��i��� �:��H8_:�$s�쌘Ӗ�;�(�_�-_d��N]N���8�p�͞]oF�Z��s)XS	�M�`3י�j�/^ۗ�TQ@�y<I�ds�`(G=x7!�{/T�ڕy!�EF`g��9+�Y�g���Z�e���Þ���^1xx�`��g˵�^>�ƏqV]��>������E�R.BaС��Df3b���B�D#��6�8Բ��Z,ą3U����3�V��Gz��a�b��5�͍�O�ʥ�O����^�g������{^�g�(�B�z�A��\1.{�i�ucEـņ�i&o7j�ф5�w�ux�NG��	�8���gb7'vZT�J�y��k.�s�ޝ��P�ݜ��;K{>��2��Z �Y{];G<�ȝͽ�ҺZ��3e����<ޢ�u%�V7w|�gl�7�OT��+���D�^��*4�qU'�����L�O=�ڧ�GF$�Ӹj�](nc}pF�Ԋ�N:�{��fk���Դ�\)��nX̩�<e�W^�Z"1���4r�%�q�6r�}�R6)M�݇�Y�bv"f�5�v�ɱ�kB�ƴ�c�1h܈��\YflB�,���:�Zۂ#]�h⦩J^�����nu�o���ei�ϕC5B�'i�eK8
+es��X�"�s�9�m z�[>���[�u��Ը�.S'�Jx�d#��d>ue�^�#<������P�
��Ϲׅ#�����Br�h*�9ƽ�r"F�^d�kpl�6;P����l?9�F�*M�"+��4������f��V��f�vH��툞�n��q
{7K|v�kD?�!���h���E�s�*-�d_J�,xj>�m�ʸ���0���&N�/*x��,p���<h��j��^l盞=�!���z��ђ���s�[��c�L��󻥴&)]me��Ⱥ�c��Y�f�l�Ӟ3�<�nz���vz�[r�t�h�֔��%!}v8��UvӆJT�ˆrF�_[�%;79��Zc]��.��JB>ṏ6ȍ�0�q=)U�n�H��;�~�i����/k�D��~Z]
��|�Kk�/�L��6D{�S+�yz'D���Ozz`X���ecy8ߪ��Xe����ę(��t��{��+zYncC �t���5���Q_���/���v$l��(:�x��*�~�Ml�L��Q����/�r�x��R��QY��F:苸o�#/���P��xd�B�H�:�F,.�5��n��2x�
r_�V� \d7����T2(dE �u3n���ܰ@�ߗI/3�͸:�WI�9����W���4�C����u��S7z�\�px���*ϧ[�7ݛV�!<up�|2��+��pb�J�*��0;��EE�=�M�ig��gv��	!���5�zwk",C�n�r����#����I�߂�Omm��>ݵ��n*أ����i���o��!ժ(����4c�.�-p��3�s:�������k��;�j�q��8�3`�8�-��-s��P`�:L��	T�h�q����(�n\q%o�;�i��~�����uڒ}sW]#{wj"��Ct唻ZX���b�-���WX���l4�A��G��il�6�Ȟ�Js��<�1�0�wN��y-���|q<����V޸���I$%b�NqN����i���.GZ��(3wk����X`��s� ����b�}F�a��;3w2�^���)-Ԍ��`�0x�3��җ�����l�a�w��w�q�K;�~�{f�(w��hbS�<em�U��,�jIr�]�W��"59�7����7�=&�]�d?��N��}��]�T7`�;�,�^��qS{u3{mNq�hqep�ⵧ$�� #��%��#��*iu
	��^-<`��ֻ��u5��cVa�1��Ok��YmR;a�7 �u��S��[8и@�E�x����+�|�\�֖�!>���,���zYg��M��:ZY'�ګ�<'����S�@��N{/�
�yA#�JF+!�Q~i�귈�L�Ӄ��
FP��OU�Sڧ��v�y��}f���(�p�ӕ��"�����k�G���\m�~+�w	ےkX=�[s��rڞ
�H���6	;�`��Z��߱p����;ڈ����,�����}c��2l-�o�hV�Kp���'�D�}Ճ�j�j�p��]էf�GJ�PK���<����9i��u=�v��{$��Z��������gE�z�g[���qwR�V6��[N\lښ��I���iE�$6==W�{;�.�
�Oyl7gULt��1������(�]�]��3��>Xg�M,Lj�`�u<���b�ol��(�Es�3�Ř�$s؄��v�\@u@�4/m�;��,p�n,�*��������i���]�E'4dK�a�$�"�XK�r�#��p�N�y--�u���^��x��x�Oά�X�
{�I�/���JY��P�F�K��^��{�t��͖��+�֢�(�.�|_��K���5"��P�^tf^[�"�;7���W4���р�ѕN�
C�q��&����t�
�
�IVi]]M�������������?H��o�5�����)�Rf���ϼlXC�֠=����͓׷C����t*�:�DĆ���gg�S7�Jq�ܙ���͍9�)�ӝ|�V�(���z������S݄u�B�DU�[�t�\-��Ä��վw3'�j��������U8mk��]��y��-��k�7�`�j���J��6��ۦ�3��]&��W��S[l�On�.�G�?{�=���̼�YN�{�Kf�H��3e��G�bZc��
R�d��so�Y� �
mnS����b�{��2����78�wgd���R������JT��q-Io� +]�_*[�S�d��Q�r�Ѱ�2��q�㑌9w��Hݩ�B��"�9~-���1�c*/c=Nh��5�r��e�w��YV����-�p�iª�W5�1<��l�d<��U�ٮ�X�A�7�uF�����lm:f�3F�r��ѣMQg�Ryz��šM�k���&��.�
�@����N�q�s��53K�zwe�%u��z��[ԏ9u�^����`x1�AX d��u�w���s�ی��&d���*]��R$����n6�_Z�f���lN��9G"�2�=��e��+�����Dx�]G��<k_*��������uĿ{��,M��i���N�
�����r��ϫL�DQɉ4V�i�gs�d@$�R��l;UR����%u;�D0�)���ZO��塙������x|7������ݓ&In/SSw����Z��K�����W�־U��O
viquG��;��K�ɓ~��%m��2�U1s��:��:Wo��7���䘅�	�Rv����d��������uc������'2Z+�3�c���i�|ܮ}r�e曙,aD?�]�q�<�{�U+R��E��!��7R�R�3���L=����E�z����s;>�����ǝ�;�Idġ�b�Lfr���dxJ;M��NCr��_'Ʊ�0�!b!�\R��{�Rz�]��I��dE4g��0p8��ᕥg�l��Q��b&&�u�$�Ǥ����ri����1]>S���X��,���ª;"�U����mu�sܝ=<O��n�Dq�����J9�����D��d�ʋ��Wz��/��f�{rh�q&������K�"�$Ru���<f�,߷����{L�Tt�e	OS����ΕGz��#�3"X��N�Y6d3�bI(��t�t���,���}�4s�������f,�6��"�����Zf݊C����$AO:���3��-p��l&���ۘ6n�����S ���P&o�^�:1�D�K��pJt�z݃l�M�姨�Xg9�\wE����x�2�<T�P�����t%M���>�[����c��p��������|��Kʨ���c�XW�5��{ӄ�SE�-b��46���ʔ���b���%�)v�n�[�af��2ҭ�����y�年�k �kumI�N2����K�M\���o��e꣕h�
ë`�D�dR]�/� ��Y��9O�oυh%���rͨgE��
&z#/uAJn>��4X�M��ɔ������}3�N\���ߕ&wA�Kq�2��𒇗���xJ�0�\�y��E^v�E��o��������U>�"Huj��鍋��㳎���,�vB��7���}9���툊IC%��;���恿�x:�0x�&[U��a^˘T���<�{��VW��`05 ��$-)�m��1�%	f��1]ˤY�����5�G��]fu:`ʷ�$��I�"��H�n�,X�A���^�$�OZ����b���I� O�㰡�V<=\@�Rڢ&���=S6Ӎ��kWBzo���e��O��rQ6Y��"��-�e�Y�s!�AJ.���ssz��]Ԣ�Ԭi�'.*ڠr��&���ʌQB�>���p�t��Uӕ�s������n6l�!�4����Eh�U�m�VA�뇵:j��C�
\*b�*�͘�i��pY��7�q��Q�54�7��m޲�Ȟ�t�6E��>��x�k���x ��4���I`��ĝ���gS뺃��|6���>v��:�o��Vv��� v�3:��z��6�p���d�;���b�i<���������/���t��8gM>�cffΖ�WB��8/�y��'ऻ>�~]����}K���k��b�@v�����oΙk��@�!P��`�:O+.{6�s�Q�.�^���Q
��,��Cq�6+�܋�C��׾�u��==s�q�'�Gt�:4r��z�Ћ��/�����.S�=�˦.�+"��9���<lm���������p�}��ez��*蕀��U���yO|�C0�}��-����5HM�ۃ>�QL�CQ&zf'x�H��ي���8̼����ȯ8����˹�;�Yx�����N�j�.w�
���.����6�Q�#���M�3r��s��\1
D�fp팜qwN��W���̓����
���S2�,d�7���:�w�x��P���"�=0�3b2��I-Ňbe1a�R,�2��qObzڛy����NRV=��S��.TU;|<WEqת�C��M��y_)����&m�i�z�-��Ӽ+H�2�Y��P�;�qT��)FZ���C�l=:�U!h�;X'f�*-WK� G���S�4d�>/+�Є:�7OGi��Q�c�ʅWug҆����|�)YH��EjVg=&�wZhx������='Z�����ܡ�{�@�#�L2Tw�P��;sb����4t��%[�@`��n6b�Q���F�]���W=�|��j+�-�K^��I}��к%oF��t�����aܚ݆mv3J��=m��N��y$�"���a�u�k��Z�p�Χ5˸f�	ր��j��#4p!27���o[΄!ڤ�W|{�9�p8hk*�vL��y�ԣ&a�c�m`�\��a�F7,�gju.�9�]a.��k��ghfo7��_W,5�s�B���6��v��2
�,V��� iE%-B�`�d
b��[�D���&�Lk;xS��R���ޏ�v�SnJT�N�5S�H���s���9$��ܺ�1Yz�J�x�UV��rc8�fp���(7�M�id7J�8�M��6�W//ej�jl*�u�a��;A�/ܱ��#��g�]��P���囱(��>ՠW'��-�=fo�л��nZ-��r���#�|eE`�/�t(��nSL��-v�Գ3�����w]�2��e�c
�7�hFE��̶Ub�\�V#�-f��������]}�p^��ڢ'�f��I$�I$�K���6��m9M$y�$�[��K�����o.�\o�̻��kr�-�B�N�8�i-3a܀L9;�f
�`Ge<�~&�U$^
����F��ǉC�t���]sܶ�[x��u�!nwX����L�N��|��ʔ�.ZY.��I�.hb0��r���l$��\���eb��V����Jʈ��**�_,J�R@��4)��( ����bk�����j��r�(vBa��Ŋ��q7�ٍJ*�M!�VwF�<�f&��Z�Z6�H%J,Ҽĸ�Ѥ���"l�k.�I�P���CVtc�L˥��l��Bt'LV��e*M�R,��y�s"�wD�2�+b�E[(�S��5}�'u82���������]�<SC�9)��އXU�T�z�o�z6),�V���;;��(�!Ն��ލp"��-0*�)_���]�X�ki;�&i�m�}��xYP�dTӗB�y��-�L��-[6vkZUa.hP����i��9�v�A�����WV���ۑ�`Y���ރw�������;�a�C'iv�X\�^řǧg(��WN滧E$}�_9�����m$����ݩjK.�b2dH$D2ߵ�E��ƙD��3Z�m��x�t�"J�*GM�řj\̙��E����m���aSX��U5T+)��l�̱q̠�#*73&�����b�����ֲ���V�h#���Z�� �۫����V�e34�t�i�C��*-��2b.�WH\h�	TB|� ����.4��c�J�f;J��e�2�72ڮR�fj�6��7��-���o5����9�i5����0���CZfa��)��mkr�Ir����=ְѬ������iJ��LJ0�e��;��6�Bͮf:j�˘�@�lV�]�ZP�M0�ep�Z�֪bg֦���Ep[EEp�T�r⠠�q=h��t�s,k"�*��5�a�ш�:ʊ[b�Q3WN�!mUnd��Q}�X�`�Ȍ�"�YL�4��h��E�hւZ���--�C�1DCn�,���T����q��X6��T�S"������Lq�U5j#i��Aṃ&��ʁZ����fd����f DT� �&f ��.f����+W��Բ�7 ���ۻV�R�T����*���s|�f���q�g�7hݝVP�F�u%߽�YY�C�3z��+�t(�u�̇�z����)�R�t(
$��n02PiNWӗy�m7��ZL�d�å���$dY��0������7�Ac��2�28LKyJ���MO#yԶ��(�� YS��%��� b���.����uضE�La���n�پ�a�(WZ/��7���n�U�u�lZ�\e��+�P}($���=����=�|�:2r�43e�p�H�(�����^Ň��sH
��'�?a��'w+�q�B��fD�I�-	�Bܲ�m�."�@��q[�ѱmp�m�9���ǎBst�0z�U��W:ɮ�Xb�t�ߋ�K�.!��e�:]8�=�{�ن��[(�sճ��t Q�UG�
�X8���e�`�u��7~�$w�q����*��/�Dy<��Ui���|bԒ̀X:��I<R��uZ_;��-�7*U~���Rάj��p&"�s��S0k_���'���*�7����C���#��Rp��B��9���s��׮�Mû�mx�4�/��6p�Gula�|���_�)�ѱ���*T8�Nk��8�篸Xx�nC|��Om�ϯ/Qg�5�o���q��a�t�'J�xk|��׷KU���;Uݖ���	�S�.��KP3�ѕ��RY��{/w��AC�f�'Q���
a����5��H�6N��>�:�w7H?�&:�:�v��t �ͽ����N�&꯭�6��D�pO�ҍAl�`�X�p��WE�����N������aR#tD����ϑ���hu1pq�g��υ���[a36���|35D�g%q�Oޕ?�"�rod,��ٕ�^�"���F�9��s��OK���>�Qd�6Z1fa�d����p��N�^
�S�Q�+$��|b@���m�o6h�p-D�b����1��o�8`�d3��ZP���*��u�k�]8���czF�ԍ�M1�!�>R;X�^�L�v��Ef�Xw��
x2�T�}]"`��dm��8w�ܩf�l���+ :�V=3��]k׋ic�����Zi�M�F��=�,lw@��6p�J�\E���N	�E�͍Rˋu�>1%D��zy����mw!گU�iS������Nt�`���ڠ͉�2
e9@�Ώ��pO\W���8�p���g,�͌����!ۚ�أ�r�.����b�)n�1z��N�W�x{�L���`�Ϝdsow���L�Qr�ܝ�e�gV��������]�x s��J�N�G#(�N�HӍ��~z�L�7y�GM��sD���H�v֮����3Q�E0�b&ԣ�K,��S6�w"�J���.8ڡ(�������mv0��e첯�X�i��#K�ƅ�����8��Pͻ��VddD�L��wk;B������7G�>un��'�T��DX����}��\vB���a\k��ν{�;�:ō%��K]��
�j��#��}9xM,Wg�l8%.Pd�PS�[������V��U�]�Q�"TC�0kin;&QZ���SV	Xja�Zs��;��>";�)�1�����S�%l�s�G
t�Pr$�hN����͈/���g��
|R����2�ߓ1c@Z�G�b�|q�>n�A�6|��{F�+Ϯ�2-OgCd��LWO{5ф����P��`5��ᘩE�3�BY�Jm��\�V�a���-�ˌ�S�eH��[��$�AA"51A'7�����r��XP"���7v,[빊wGJ��de��	��Se��k��ᾗ�jZ���T;ys��iN��A����X�t/�q�|&'	븵���X�p�^���&.w-M��(c�:��r�p�;��ub)��V&�(��YӴ��sݼ����y�<��c���l~�r�'�̡�����px@����2D�ʨ�-wr�{##q�Ƞ:�.�̻�u�}�]�^4��~6�ԟ=��Be�W�p��dK̋���sc�A�r���(/L ����q�U�2z�>�/����9�.�Jr�v8�J��ɲ�)�O]a	���|pN���4�.��p+4��u��)�m��$p��.;�Q㣧�;ծ��3���W�l+�:m�7�"xH1 ����D�'iOt�Q�&t�6��D��r���@wӄi��ڴo��t`p�"�m�w؞�h�9��%M&x�^�(չQ
�E�qB�|���}����n-��ٓdbv	�z�����
��t;f�E�C�y������
ʩˬ���e�+o��x�ROR\��W#J��#�����y}�)|M�Y9����ߥ͸f�l���oA��f�G36Qmϭ�W}iS9QMM�B,ČtAF�!$R2ɯ2w'��x7�\[�I��vS`�w^>��W��2糞2��ĥۓ�8=�)���c0M	$�x�cp�<�+t�u1��71㳑�>�͙���q�9\�{o�XG!�7gj���)e�	c8���)�pt��,��N��Ƃ��K=�;Ǔ��_�.�۞�L~�n�ʹQ�n=�M8��j8[f�ȿ9f$C$�hB��>YW���O;7��e��˪>T�x��j*T��لBn�jD�R�j��A���G����p]�R�=�A�&*|�b.��
U� w^�2��N�ꇮ��o6ЧeM���휇7+�;%�>�K��z����-�s�:����Ij	k���-����[����p�u�\ ��n�/yQ^��\B�����HTq���͍�U]v^��m�䦲�6�zu��F�7 4dY��0��hl�qўX�n*���J,�kUk����F�C��h�4@���ww���<0h����:y�!T�ȏ'��{z�9k�3����W
3d p��H��S�����F���5�!_w�o�ܸb�P��/��d�{8o�t��}<k֥�Y[L�4�c��U����k�L��Ϸ�F����r�o6�EA��ǉ�6��S�çؼ<Ni�;9h�|����d�<wi�ma5"��wy�l	� ��S�i[�>�*D�E׃:Qͷ�qH�&����=u,��(^�K�j/�F�P��T�K�o��[S�ؾ#�	z��8��O��g�"��J��Pg_Vw�Z�o4m�ܼ��w.\�%Z�ƙVԼ:�Fi��E�V� �n9x��U�g�wJq�ss�:!�(q�21�-ӷ����Y��x�G,��w|�v�Tmm���;\QQ��\�G���AP(|�\��;;��vt���|-���F&LTE�Q{k�U����R<�֙x:+�Tj�Y`�8!N�\H��qe�lq�[Aߪv�ީV+$�DDXnz�w<S0k_��>d�(��ͼ��Ϟ���!���tU���f{�N2��U}���0k��X�W�/:����R�q>��C8ODB�6qyh����lt0[(Aع������RQ���y������-=#%�hDHu�M���S�|'��.�����CB��T|3���(B�6��RB0�ͯ<pY�Nʖb��4)��
#�[��^}�|*���k��=�rWa�Lư�Lq@�P�a�ۊ�1bC" �u�����m�Ou �sr��t�F:���2�� ����dCF,�>�0Y�".Kg�G�ȁR�H9e�[ͧ���/��V��v�Ӌa��9{��^�x��e��*��}�kզ�?=��Ⱥ��n��u�PEޱ�����#��nv�jK?�	-X򩊈����Wޙ��rE�NY͉b0�^ϕ��lrw�U��(��S�()��ɘA��*Y���X{����;��e�8Y&�,���_=�|��[
��M%,r�=�8
؃�
��У�-��\�2�l2����m��}�4o* �׊���wm��7�PP�ī�QA�V��P����&�k��M�t��s/k�Jx�
Qt���6�W��2��\��s�X"�&8����@t�h�ݵ*��f�]+Q:��T����P턡A�zD3��TX��[V��s:z�d�jW�N\q�s�\d7��s>*�(dB��S�����R��R/��F�x��s�<No�h�ka�(VÓ�@{}-�~����[w<�t�a�Y�Bz�uQ5���	�pB�r"�U1+����u��C��c'
:e�����X�1Z�Han�ت�ed2���Z��Mn;&Q��'����X<*����a�����**CS�t�T+����6�K_u���_\p��.uR��.�nN�!L���G5��sYl+�\}������j�ƨ��͓�]�i4�d}}�.��X��=�����_h�Q��6�ؕ܉�Ck-.��˅�6�fh���Q&�|���t�i�*Q�uB���������ёښ^�{&�Xq똺NL]֥>���E�n�uX��/k�g���0{BJ�9�ˏ�ݾ�-K%#XO�/��*�F��r	�bB�Н�8�p�P�Y����sW�#d���\u���&�W�q�K0f��WU�e�0�r�D{S+�K�|+�E��\}~}�эن���"�X<�X=>K� T��[i�a�Ņ��t���
ۛ�֒;�҈������ٜ
0���7&��se��R0����-��5a�8��}�ݙ�b8�Y��U�E�:���V5@���	�^T`�ڊ�S�]/3	��k0$�v�V���C)�^͖\)��Hg=u�-�̊�ݣ��&�Lt�C���A�\I�U���/F���D��{Tl/v_nu֖Yï{%UY�;�m��=Q5��sa�WPUP�;4r��m��إDY��4�x��-t��t���?%8(�뾿�-ff��s=���*%��	c���.��|s���U���"����\��|����Grdc}�m��0��N�E����gG:+-���c�WP���ٴQӸ��V���I_Z�7�WW$x�㝺��!+WA�m��x{�6�T��j� }�.�����M��(ӎ*�҈DIG|-J�x���(?��}Y{�{�>���S��*n����Y8NW�K�,���7B,ZO7�/.��A\�-�Y��;훌��#��l5>� 0���+���VJ�p���&�o�����9�.Ʀ`�f�8p��v��e����������J���vW�ّ�nUf5m��\e�F��Z9P��.})M8%w�-:�"�N���,�Q�g�/��&��v��,c��v�}�DGD�E�O��g���V&"�Јnf����H�e9�vrc:�=�;).e�-R^X��cD���)Cq�!:%[+w���Ә��cw�G�H�1�
#D�T�B+a�`��R��E����|e�C��q�z�r�G���nH�@�� }Yʎ�h����������J����r�_n��/B�u���9u����%�_d�'�3�ёfh>�1>k.���qq"�V'��b�|[��c�Յת�=;ğM��֞���vA�h��V��bB�;O�Xڰ�����+u?��-NN�i���:�y�f�����;��&T��s��2�C�_ucAu�*P�s���<�s�:nf�oZ�����Z�ʾ[\���� �s#�G��σ�EeU lۆ*�>�qF�jv�xѳF�L���`�;�����kR0��o�ቄr��H鼦(f�@�@L���)Tᰵ��g�����Z7*�\x�,�Ӫ5�8ҁ���T���ʭ4hZ�6ჾ͖I��ґ�8�D�l���1�3�$�R��f��ܕ��vb�^?--fx�<LM��>�^1xx��U3�u�V� �j��n]٦��)CQ��d�;
��|L��cZ�F��<=�g-h�����=�q֞�i�֪E秩m���^��(U̞&�BҳӴ�u	��z3x�"#�.!��k�Sك�Y�Ň.��Ί�5Q,�Qx���yM'��v��,��E�x���S���Hz����$Zt."��'��)�/��k����*�=�8��9O�J�X�<r2$磥�,��������'*_t���B��r�#����܀�wP�><7��}�_�yh�+��`�R�������I&���{�ӧ���δ�����X�q����wZ�w�.Ω1u�aI8���w;�f��^m�ҍ��Wq�J�ͷs����� ���fn��'�W�
ܚ!Nr��tF�][�Z+�
y��*�v����6w&]j��d�v�
���&z�b��̅�ߴ;��c����F=k��ɜ�p(�o���x:'�y]�ob�E�����=����˻�B�	�u����Fr"�c�C�V����wU(�l�့<�q��L>l��C��gT�8�`�KYK��o^'؁���[v��Ҧ�{g�ԅ��'�xu��1�C�������[��[k�\͇�nt��f��c�{�
�C�T��ނ��>��ELN�A�J��Ż�'泵�}\s�%�pX0�c���|�Q˭v�� �:�����'}\�[�W>�&�,�S��a��j�G]���Ŵ��xK����2����d7[S:���N�s�v*6JG֗j��h+�8� 
��ا\�
>w�ɮ&>Zԡ�)f���}ϗ,��FI]�dRoX��	+V-҅����@�aW�n�5�C�O��3�7B��I[Y��lb�s�y����A=��5�eL뛕�bM���T�	FvXګ,|]_*V%t)s�|E��J�+\ö6aw/88�>ͽ�z~�2����:M�o����՗*H]u�1�+]�=xl6�D�v�1`T���T�Mv��"��Wx�v��8={ۋ��I$�I$�I$�jwM��0rǴq8C�|�4�0]'M��B#�s�!�V���Cz2M������En����v�+��6�Ǖp�6�]���j��4:bd�<m�2v�hwPi6y�Ρu�;�bRt7�`:�W�M!gV�vp���c�`�ފ�-����3��v���Bҭ��*Gq�dT�N��Mv�*m.�9[{�-td�/i
c�Y��飏6�Q}yHS$�|z<t2ua�N�L0��2���ɽRG��l�3/wu���o6���ɶZ�2��.}
+�T>��[P�8±����V��;�䬭yZzN��D��9���f$�H:��?��:���}�J�Vb�.�b�uLDD�$�4K����xo�[�H�.r��̦����9�u�V˷{�+���l�/c�J�\�2�)��C~�M5�\0�	��\�l�4�I��(��SA
�:tf@qm%��ޫ=�7B�u�z�P�!C�,��� �De�*d������Q��Ф�7N��Kh�ޮm�U��׈�]@:kvE}Ywa�$�z��\�Ãp��d�Ϝ�}o��d��s7�C`�����Q����Y�w<�y������j�'w<7�Θ��*c�$=��U�y��t�Ӣ�>�/�T�y.J�6�$�����%�H�Ȃ3���_l��LQ���1m�J�o�[�\U�uH_�mޫK���UH�Q�1��]e�f��Mj��XYK(,Y���Į�ѫ���ZcK����ke�5�\L��q�2�n�5�ʪ.Zʖ�c�W7f�sm1̸�ۘV�;�F�L����&en�����A�\�\eAW-�[�=�0M2��ޮGEs5��b��ѩ��X)S�ȱj�%T)�4	 ����,[�E��.��Ȧ�10�eݩn�JWc�H�I���˻S\����-�1
3+\)�`��Ŷ*"�+Zm*9k���3*�����CL�E��߯�;1����Rk�&��ͳ��ITvܵЖ���,`�,P�Yq���j���Z�fcm1�(�r�T4�)rəB�-fq6���4����o7��b6���-Z?f.4��ۦ���ZT��LB��FҦ��d�
�3X����q3GQ�V��F����tS�'*9O�ZԸ�p����BB��,�lDQ�q�okm�j�)hޝ��%�ː��N����ɾ��S��GoX�]7��QƴE���"� ǚA]{��>�6[��.��xNͣ�ž����M�����13ԋ�T��ߜ3�����JA����F�R�审�V�ɝ�ۈ�w3\m�B�^4�\!�0c#��'XZ1fcS�Jɂ�G�8
sp����7:�5����j|i���ؒ���b,�q��9����f�q
��yNRb��ő��:��L���0էL�̰p�wO���V*�'}�L[=��5*��l�ێ���n�B��h:K>iX��/�	r?,��:Y'���o#�Me�n��ZG%oR��;ɰܣ�S���|.B�\����91��l���x*�nM��q�]�P��d��V�;�}O#�y����u�n5�#fC8&$�(���2+�vv۽K&d�E���E�E��#�m�:9�t$f{Unzk
NХ��gGvڕ�l�9�����_WDVt���"�J��27"�T��wE�8�.N1F�.�r7���k�E�.~���>���l�.�3R	9 Z}Z�N�r�C�Pհ1�X�c�V�M]ܘwe��a�ci�N��e�j�
�H�%�59T<:��_:�qvs�/wL����f.�6+�ǯj2e�8�-]�-��;6ӇN��w�]P�?B�8,LK.�G|g���Tq�r���GTϋ
�sr�BobZ�yA�>(�hY��xx>K�`�ka�?l8�{	}�딭��I��wVNm�gEj#��mz`hWP��DX�,�Z�o����[�3)m�x}��߽=q	�৺�|�5G¸WZ�ζ��W��xL�͇�����1q����˹),(�Sӥ��q��t�'Zd]*F+ʷ�0k*�;z����~�:�Nf5�<E]8�G<}�#)�g:���0%�����6J���e�|����Nu���Jɴk��;Z.�W��F�7 ��$-:�m�8f1� ��b�u{-rn�rE1�,��4B#*/O3YtCp��z��"͑��H*�fV�ؼ�⺓���;-�'yY9�e,����em�=+�R���H�Фn����_6���0�*��Χ��)̙��Ho�D��g�ǣ�J��=㸈'WVSHW��=�w�VO��wa+N:5ږ�y��ѶwU�}���';_ѽ��+G���8�UǌL���z`��Pʹ��Ky���f�v���%��Tf����s}'Y���;�I\�li���dF[�A$3�����:N���6��z���������c�/�v���6���Vy7`���B{וꍨ)x��*h�ky�!���oc���,�����3��!fNdW5\v�LCS�iK��W�v�ۙ���C���k�W��l�E�z�l.�,׹_<���گd��*эsW����Ħ���Ea���ϒ����-?0+e�UC^�����:��:�mCʨ�)C�ׅ*;՗�<t��e�
݋����Ǧx�Bܢ��A����|P��#�i���s}�:���=�p�xٸ]	��*�����t%,Z�|%/.>s�1�n]TnjM�ԍ��ۅ~[Pf����P��Cp���]���
��XQ.F�Z9Y��=���緤��6�[���`�Y~�>�����J�ʌ�Y��E��9 �6���H���Ԛ�5&����i�{nْ什:��Á����`��̋�'5�u�V�8��Afvd��NAkʈ�֌dx��nUZ�2>u��k�:���P���eh�&8��f`pb��Z*��Be��e�@����+�7�"5Z�D�[�z��Y���].�fonIH>Z�+�|P;��Yy��{�)AŜ�e�dt�t�Gx���5$��p���yK��+�͘yٱ����=G�]����ؽ��{'�m7��>zt��>C��E6�|���V���<3޸����b��[�w�(Vgu��X2t����P��G�L>�KF���1�����H�3����t��d ]x�d�ъ��r"Z�a�zY�͛�"����� ��{�����}Zj3�7e���,���Y؋$Y��05�46x�K��a�ܵ\�����c����ʠȡ�?B��1~,��m;�7��h٣��Ӽ	N��eP1�v<�)ع3n��Nזm�k�[�:ux��9j��R�p���li�V��CW��V��8��F�|��t�_KX'��?���<�A�x�&�F�Q}�!@J�m�e�n%һ�s�<��::b��Y�o^:~?(Z6�񷉇Fm=��<M�g�/D e�޷�w]:=q���Q�Ύr�8�n2b����"E�A�g��hN�0G]K�{o�D�ވ�ƹ�^�,ٰܢ��"�sճ��AU+ФX1o7��Yu����V�V�U�����������6Ռ�2'�cV��l�o�Lנ�[NX3cP�;	���.��Bz��uE��u��ڹr#�siL�@çP�Gt����g�2��˻�#4M�Z��qs��c���ݝݟ��̎ԃݠOÝPؗ[�(�1�=a�A���c:!�w����d�,�y���cmV�T�P2��4F�B:c�*�������`k ��"�)����
f���|�ή�0X]��w��3�E��\)�upc�&���l�O��
�v��ެ�x��W�F�8�o��1"i��\�B3���jg��j,Ύ3jM�]8��xem�`t#Z"�)d@4H��HX��G��^:/鋂��dIU�B���ue��΃f_��A����,�63��?4���{P�����^j��������i�|�~��PQ�y���f8�Q)͜h��t*+t�Q}@��}��{f�˃�M�r��S�8�yT��(WH.'a1i9Ȋ�Fp�d������Že�)�0_�K"h�ҬL��졆�۶s��P����)��mf�_oh�Mզ&/>������4���	�Y<+Q�ݰ�]h5��'~��+ N���f��<�M4XL�[��t9rt��Λ��*�˦�n������y�c\+r֣w�XȤX�>R���9��w�#�g	|�f�ɋ�yw0�d�.K��=���̱t�0< .{Ne���a��ٷ�g#�4/��-PPިYڒ��m�i�7��g媬Z]Ozt8ӷS`�1�82=*+�\��u�򧁌�&��sn7w���R�p��t��{L��wS�݉��N؆dS��ׄ�Pwf���1�7ٗ���{7/n�IGt�Qc\��ޖ[�_*�#���i:ىf�=F�aS�J�d%�j�C��&�H������S:�S��z mƄ�#9���n���U���S��y��8�%��HV�����=Pq�sˌ��3w;��>�[y�Z�ʷ�_EC�
��H��sǢgb�R6h�SP϶�C8�b��ҭ+�y��O/u!��q��kF�@)�*ք�;
x�EhR��,1��"e�c)�{#J�e��+��B�#r"Àȑ��+�၂{k",�f�q�K�\橼�D���2�+be��i��8�:l':dP�HÁ,�GLo�`hA����zv��߰�7hvxVo�llzg��m7�3`��̡J���y(��ʗ[-
;5�V�$�R��	*`�y�(��X���UjٵG����c<�R�J-cr:�������S�9ۻ���N�Lk���Ԕ�eҜ�*�c҇LĔ�ά���L]�w��9�,��Q]܇.�gS��8�N5`~�^���S)XGG��v��%f]2f�x����X{&�2	���9͂C��.,໓����˴�u~��LWO�\6��B�q���{��Z�>��!(f�-l��u�v�v����v�@}܍�K��H�:��gi`��T�c6<w�hMӀ��f9=כ�Q��Q+�{�2���؁9̙��1A�!�,��e*eT�xdf�ܤ�'T1�h�7��e���u;��=��M����Vy�+Ϭ�2޼��j�8�ۍ�v�aL�PϪ#A�@׳g��
���3�u͑@,�݊ƫ��dwX��>
z���9��§MU���g��q�:��C�]��齴�r���7�yw��y�Ƭ����a ��1q-�td������Xz0t�^��
o]<Hv�ʬ/z�5:Yj��]IV���	V��<�:�\OM�e���R8���2�_V7NJ�J3���l�0�L��W�V�a1Cj�����x��s���Vw�iSS$�W ]t�x��v?1�ݷ֒R�Y��2*�Q���$��"���������,)S�h�5dO����M���ɖ4�k��Mm�����bp���	o:���R�Z�C�e����Q�qwm�r�K?x�jٷ��L���,�߬�Ep�P�8�I��3�U���HDu뾶�v���mKi��ʺ���
+���_^�F�u9O�(��~Uz��Ƶ�t�rr��Ib2��=2uVKZ%�ס9��S�T�@�ӂ�G�8sq�X�[S�QQ��4ǣ�6�/j�<��uRsk�,]�o�1)y^ޙz�w�qT��ہ�������72�$Vt�ŧ]�n��&�W�Mn�ǽ	,*{��XTL4���+���X�)9!�5]�ϒ:��ˬ�X�p���L*;47y�k��u���r�4sf�\������	(��}crX��Ĥ���z����� )�řυ֙��˄�!	�]�.�v:����w�2��`�gb�ƒ��(&�����Yr)��r�����x*���w;�#��/U�7�0�!=�s��͢��͠3b� 1��N��<����Hޓ18�q������Z��{'�M�1�sR��u��Z��Z�3ԅ	�Ⱥ�q肫��q��T5� �0*�D	�t�Ɲ�Һ�dl����#7R]�_S\�ã����r݊�9��׻J�&@4��B*�43��iiTP�~=�-p�%�L�����'�W�g"�N̊�M�A�ډ;����/Vۿw9�u����;΂�#��E	�g��ע���E�q�n�F�$Sj ���ݹ�C*���.�#��2ޱ��;]f�����,ܺ�f��|#��n�.��)�&]�Åi��A���t����\!�H��m)Mt�.w��m�]�i��Qur���я/^4��F�7�V- ��9��Em:6���:��{�"�կ��t����I����V��-��M����n�]�U����Ng+b������`�O PN̡
Z]zx���n�I��DS�[Z���L�cQn��N,9�ւt04�R�z��������y�x�^g��%#��������NN�Q/�zºo۽��wj
ܵ�w�u�D��=�)�T���p^=�8y!��-B��OG�-�e�;I��4ԥr�Z쬵L��ym �ܡT !�)b+�)F��PV����Ig�wQ�֥�F߅d���\(C���LF ���-3.��wԎ��*�ݼ2�0NIʺ�z]ur��a	LD��yԫ�;�k5��t�n��m�G�k3W�t۹�C��>�IE���+�V6w{�K���Uw4��AL�=���Yp�����]g8��c�-sU]j�}��۫�%�s~oNS�o!EE�M솫^Jǋ�g*��������^keS�o�-W��݋.[����M2�؜�����Z#�T���u�L�kT�t[�����t1��r�i��6K���r��L�6*5H�S;��g����b�yqwd\��o���{{��Q�G��Ѩ~�g����]�����K�73I1�I�R�'m��33P��.�9u]t��L�pջx{�g���?���?��qS��Z�����4	���9�@QP_rː
*����D]����,�:qd���]O*��\�̃(�I$�"!$$d$$HI	 �I$$�$ .S^����`(�B@�<�e�m���,��rh줪"��F��(�q��}4}k�74�ћ�4�Z��E�+.5\>xᄒ^�ӋR�h��0�X�h̳��k�H(�/���i�G=@ 0����8D?��� U�G��	+C���b�jp���{�޾�$�4����v�x�{"N^ (�.?@<��G�(b tXi�� P�Zz�/��B��K�M� �֡3�K��n; <v�8Ϊ���݂�Nd��@T2�g\�;*yR�eDT��EB��1X��r��Bm�p��S�����j�*��TKq�	;��&�ۍ�t���T��D}�r�~��	mʫ��>���;O�	<�򑗋�&�A�����˜�Qw��j�%��݁�����]���@�}9OgO2�:�$E�j�����<5SJ���xnÚ�*�� !�w�tC��4�1ų���I3��`��@�
*�ي=`(�/������[�����5��'MC��İH��y�5QPU�\�H��"N&�h?�>'�} I$	ɲ�f n7���_<�g�E�10JA�,�B���!�	2�`Z�q�H{ʠ���4��Yݐ�ި���|�B|�5�z��	�{�ߠ�i����?-c�hϖ��Yc�tAB6�W�G'�DBx��'y�)�ݤ�+���TEAx��l6��X��%���v�"���ł�Lb���'�������Mk��A�ߚ�ɁŊ$=�(@Qig��xϻFAk�"��tG���1���a����U�P_���p.�<8$S\�tăo~!B��.�oDtɇ��KE��K u��$"�����S�hmU����Ç`��/�rMip���OL��Y�������u�R��5D�|	 �m(�����w$S�	+ ��