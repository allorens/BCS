BZh91AY&SYxF<�m_�py����߰����ae~>��   /�  ( AD�MD  ��׮sT��F�2�����tuww[kn���;c��5�UfͬL�릀 4 � :��ӟ|s ��(���    @ P      t�  @8)�{��y��o]l�u�������������i:w
+�y/l�z���n�07���a�r��}���'������7�M����eV��vt<�{\�^���]d��^��O{���(>����[�� �,�}��1^��m��wu�Aѽ�:z������s�l���쥽�;A�����3֕W,�� Q9���g���v^�yYc^�V�^Oaӝ(��n���UӪU{�l�T�y�^�֔wgnݠ�n������ tP�9�t��47.��ͽ�q���׶ٯM����܆�d;`vٮG�f��v�^�w6���\�oet
we�3��ma�]sw6��h�q����l!�   w4��s�u�lԸ��v�W-/cv�e�]n(VtL� T������aƞ���!����$�ܷ�v֨���-:ѫkg��4{X1��  4���[F�O@�C��h���f[����om�ы�t�+��xSl��thhBP��]�I��+ZS &�]�I\�զ�x�      �  T�*�* � H �-  �                   	T�&��T�DFjz� �&�i�2	L$$�*��C&bh� &L��	M��%UO�0   ��� $�R�ߪ�i�@�  �  �"T&���bj����12hш ѣ�	�2��6��=M3S�������&����g��F�Yk5����v���x�G�?hy�:g�E 6yhw�߷�� *��(��~���x�	 �?�ZO'���������#�r	�j��?	B�)@��.���k�5�ddYW�����S�?�������UR�(��kQ����3��/��?�8�&���O��xq�\r�����p���x�qa~/��Ň����a�������ɉ���N��A7����Xy�#2O�NԖx��,H�8e�MG������$�$���8��0��}��Ue����>nM1��C�2'�p�&��;m㥑:�^jS&�C��_�}<CȞ5]8?&�U�JؔG�51��DOw�p�:=�VA�H%nJDʝJMl����Ӄȉ�H���?����et��:<䯑ؔq�&�DGޕ�?"sܔ��"k�����R�N7)��D[��\D�MJD�2���͕�å}>���R#�(}��~jR%��R&?D�y+N�=+��%"s9+�[�H����÷r������%"{YXp��G�+��Ӈ�'^JD��i������H�nR'��T숷*�=+��%"s9+�[�H������|ܤN9)��Æ�M;����/8ʲ}vIҙ"7��U�3���Z�]��=�+�fS����U�>����'��W�/̮�%�K9"H5,�;<sbgY\'�$:H ��*�~Z��Kj����G�ķ%"�u���Zwg2{����'����Gb^��rOQ<y���[���U'~����&d�6z��="5<vD݉�d�UF�;"_��URi����2�����+�vAߦ���we]�;ؘ�K��)S"�0�a�a�a�;Q��}��M{���߹zk^]뫽�]b�ō{��f{���ߺ��,�Z�U򯴹�^�}���w�.��V�r\nT͹�����'$�nS��e,��ez竒�Hw��H��M��}�����9�.�MڲD�$�!�OMF�^�|7��R�I��+�|���M�ܕ�<qI�Y�Ipl.�y19F�/�=��'~Ԟ���l��N_�N�'�&6Op���Y-��ĳ(�
�Q"D����7Ri�����'&��F�����A%�m'��o�?9	(߼a1'S)&��ޓ�v�9�W����*�o�IG�v�%���7'��c�q۲M��$�} ��1!���Rz�=�=�Op�=�q�|n��n}�~�F���00�����zze�RB����1�t�p���8�B��DԆ���bJG�#���&�7�a�-"j%�l�?'Q(�H���hh�����?xH�k	�gɌ'0�tG�������8%d�4�I�����a'Nl�&����H��(D�i�['�d���.��DL|J;��|����8>�M&�ӧ[&s	�	Ӥ�H��D��$�X�Ĉ����(�H��H��RaE��:���(��D��ȑ87�N�D����	��'C�K����DI�<h�cD��'��'NĈ�䈔��XYq,Hy:P�ϐDL�D��`p~Oi����C�$L=�>�'N�h�<$��I���:R&q";���	���Z	��$*�'�K/�ɆtG���'>�'a"_R$M}���?p|+	+�a��,r2QдORD���0���a�ؑ<�&��7�l�x�_`�rYۨ���+�LɄ3"�i�ʖ<�x�7척�����:;0L�&���sC	�)��o�,�8�b>�Dj}��aۖ]�>{>OB`�H=!�{��K7e>íT��ʉ΍���zΧ&%��=¯�u+Ȏ%x~�'�%���*DGݨ��Vn�O֔��p�m���,{vd����3!���9���l�n���{Ś=���N��ӝ�=�%�9>G�'F�S��=ji��p�%5;u�I��ݏcꨘd�=�zG�Q:w"t�ϓ�9"Abt�>����;UŲ�p�3��'����R�G�����veO��TN�dI�Q:zD��O����D}�)��*N�D�Ȟ8�$���z�%�JѩdO�w���b7��y��0�N�=$Dp�0RM:W"#�TD\��ikR���� ��	�T�ڈ�6�%�D>��A�"�J�Q�����FUM:7ڈ�91�OH]ϒ�ܨ���/�J�jt�C��Ï*Qᝨ��j"_�A�DG��UR".T��=mN�}>G�d�Y��$G�72�+(gm��k�����眘��#��Q�v�7(���ra�x!W>��O����=��6�ߡ�C�C�H�bts�;�M$�eD�mN�>�D��"hͨ��"lji�D�޵,��}	�p��G���Ld��ټ6C���c\V<��3�Xf5��?�)�v��ԡ�*#����G�iXQ�4�ʈ�R4�%&���*�!Ǽ��ԭ<uڞ;�ig��IϦCT̶���1�y$tk����7n�:L*E`a�Q�ε��cW槭M�2ԍ�V��=��UD[+�J����%�7��YNaU��)R�i:id�ɇݕ�8��7Ҝ�Kҩ���gJ���=��Ք��Tvf%dJ�jz�Ĭؔ�Qf�{�Ux���T�i}J�_�{�Z�MzVo���s��.D��r�jV[μ��\>��\:�q峉�����J���/e��rNp����G'8=�{<eOIr&#�v<�V;R̦�T����,��kqיʒ{���f�c�5<We_
{e>��n��YڎM2ڙSL��ٹ�g'�|���W$��;�V�LʞI=�mg�=Ͳ����6�R>f�������3��s#���!�569eX�+��C�Tv]};8w�Q/��}�.mG��d3���q�H���1�������]8<��d���,����"uex�5�p��GbQ��5G���˔��DGxJڕ��T���M<ܤE�^8U���V'q��~��l��F(��.�W"";4�ϧ��R�8ܤO2��Zxy�_?9)��]�JD����
�W��ܤN9)��Æ�M:<�_'��p��D��H�ܭ8<�}�5)���"&?K�Jӣ�J���H��J��R%���|e}_7)�JD������4��O�����>�ݒt�H��']��&u�C�-U.��M����Õ0��:7r����'��T�3�0�2�vK���Q9R�z#��6&u��}��C��	P~r�����Kj����G�ķ%"�u��>Dweiݜɩ63�2ɒ؃��������۞9�]^�x��U'IGj�4vI���:��������&�4�j���8c �J~�MUW7�����;!�=�; ��vfz;��f2^�2���~/�25����!�P�=Q��n>io�[���غ����y����u���+��=տuy�B�*�Zj���q��'\���{���d��{=��_y}�Z��Z/�k7�	(s�b%rz�h����� ���js��va=�J�;.@��%���������ܓ�fQ}�!u��I�~	߼��2��?�����e���?����~0�Y֏?=)��LY����uc�[7�'�ǜ����!B���ʀ�
#DAg��hD�@Hf��Bs�8CbQ�Dl�
xg�S���9F��г�M�|(82H R4y�4oH4����g1Fl�ä�(�j06B`I��#������8]�08C���&���	Gf����0HA��J�A!X#�|�B�&�:���lN-���:R�H!��Bf� A,h�V�h�HJ�ZД8�V�:Q<pb<!�� ��S���N�	�A4<�a�Ud!�8*/�4&�		U�L�B� bx���馜(�Q��0�`i߲��
4!� gk�=��pD�	�y��h� b��("�:1�A�ADQ�h�G�Ã ��Ȃ�2�!B��X�1(�@oY�i�( :&��,!� �� b4 �!Rw��!di��ܮMDt0�DYѝǒ�F�y93�3�ʄ�#	�{��6Hw�;�b0�0��y"#da����C������h4pa��g�b}{��	:5�R�" ��18�'p�phٮ��C�	�.竻!vF2��v@E����@�y���������1X�04G���0�S�x����Y+S%�n��}�n��<M�Z�oFa&!�<�2�,h����Ì� �+��Y�^����%��Q�@h�6����a���\�Z&ld�o/r�#e�����uʫ�A>���<����b�3�åP�	%8�p���n���L�+�Z.��py.Qr��"�a��� �$�4����U:F0��iu�}~�͟}��?�KW a1$j�:�V#�t΋�xg�8�twè<.����� c�gqO�לYQM�'�u4�k�	��9 �f�����P~GK��A4j���8��]�dY���^��*���g�gS�n䳃5%��/̽�e\te*�óD����rW!�!ά�erU��	�����ŜDA�-y�}�Պ�>�\��&��=X�U\����x���kĚUsc�WS�����aD*a����3}⭋j�K�8��ő��2��/�,�ȱh~��\��3���lΥܪԩ	!8x֪�7pq�&�8���Zy���C�fqf���h��b'$��u����-[T�j�p�~f���� �|����qfMZ�)��GӤ�"��Ʋ�wGQN<��*����Ĳ-�k-VU�G1.�`w+���hs�Ύލ���r��ع��gV8>Q�9E�G���#����^���A�uk���?Jt2Si���\���td�һ+��)���R���^�#ѭ�=`�C[�i��%�7��er��I�M�tsЅ!3�YP��<�מ]��g�zq[0r��J]g
� �уi��.Jy�٭�c�h�<�
���20e��L�׼A��������{kXE�Y ����9�RLG�e�B�kZ!�$�ƥ���C�,~e�qb��1���wG�����:���¶�/ȏ�d�h��2M�=N#X�3"�P�D.0��+C���oG���ѝ޲��,�,�ď,�����I��D���+���E��T��0��9��$[F�kp�4�v��+�ϑ�������Շ�E��K�7ٜH���2s�:�:B�ty-g��q�h8�h��qV�(�,�aV4Z��Ӥ���!���Q�LYQE�<.M:���sɏ_5�=DY�=ɩ;�r�J�WtV�Z��gF�u���N$��=���K��z��8�Y��cę&O����9����x�K�:��<��Z�ϲ����i��:�{�>c�ǞXT~�5aŚ�YL�$�6\I�2Od���ݜ��a��	��Xj8-���X�s���uq�������չ�Π�5eX����ȳ����|:��9�7�;>��ww/���aVgs��>O3���|��G����fw�M4�u�ϒu/s��>����q6��5��"��֔���ɲ:Ӓ%����Q���=Y]Y�:���:�����������P��=l�S��>O}��g]���2�Gs�nx�w8۟#\G��hM���w;�'�͵�]�ǒ�Jew��rV�n���S|x�v�0U��q�j��ֳ�bT�5��r�+R�+6;��ҞI�E�6����ҹ$u�5-97��ra��Վ�d8J�J�\�a�=���N{Ĉ��ǉ�?�?�{�1#5Y�_	,�Ytqd��%X��{��|X�}Cן,�6<�;�-đ���T�^���d��AwJ�L릔��̤�4��%Y�6��|>#*�
,K��%n�#}���>k����%_~�I��嗾'����)h��$:#,���VT�,�MC֌��ԦU��bʴn�c�&�u(�죵��gen��?Jeo��\��V��S��:�L7��C�
�Z�S5�v��_��H�O���egxd�-B���;�S�*\�h��cV�d6\��.�6��j��"��FL��>�p������J=���J�Ͼ��XU,�6ǫ&�X�f��X�a���5��ugx?�:���oH��"�k��H����%�k(��;����E��ű�F�7��]����P�x��u��_�zǒ�6�tq�CdΣ���}Y�I�/�4�ȇ��2�y���.'�D��G��j䉳�\K��y���7G��Tn,�fѓ%j����}Jݎ�����:{+����`�4]5;u�pd����HC	$�t��h�Ň�	%�����e%ő!FC ��@�AB(h��;N9�x�tb��H!���ɟ�����f��8;���?f��~��8�]�DD7�֧����bc���߶tWmbI/{�yu������<�8�N.{��{�z;lF���ۭ�]��~�����ھ~�K�>Ի'9عS��c;7�N�Nl}�J��W��q�[�n���r]�����S��W�#���}��ޮN?=���E���i�_���|�M5|j���^�NOm��r��~cߢ��Խ��ļ��{��9��^�9Gޥ$���)���x'�vT5��b��,�Q�L�+R6����Iom]�(�M:���@�U67#��qoy��S���|#Q-q΢���o,q!B�>���t�ڻ�~��9��ϲ]�歗��n��]���9�X�=&���������$��}/ǻf����s{}�[ʣ|�n�I�V������	�z����꽯���[�Ɵ�[9�'oz^��^+Ӯ�y��=�ýٝ[y��[�{cӯ[��7����H�iW�v^���r^q!��դ�uh��?j�u>��qso�n������q��wܻ�$���v�����:�}o�.󖱶���w��s��˲w�O�y�ںN�7�V��t�S�������������y���kw�;hϻ�u�<N.��V��_|�oS�c"���n������;z�t硽�y7z��Ow��_,�{�.�u�us��[/��.�$��o��'6G'gy�W<�,w�7�[��.>n���z�؟���5<j��|�;�kݜs{�w�Լ�R�$����;�]�ǳړ��q�ӆƫG��N���N���w��ߧ%l�摪u��YH��ɱ"�UM���}�Q��\|��'��z�c����z�s%���'���9�l��	�`�޻Z}�&��h��}y�ts���߼��Ij�'��������Q�bz�/8�=,{�*՞~J����.˨Kb������E���MW˯��9�՚{����Ͻ��y�9���ZD���o}�}�j��z>�{��Mm�/7g9�qƎ�/-���J�~Թ�}���z�[�\H��ﭩo����Y���qc�ީ��9E�ޑ�]�	��ol��+{����䎓]��\����.��iar侌�?���s�	�4�d��xG�M�bBO`����TJiS���#�E�q5�C*V4���£
���v�Y�l�Õ8�I�щڬ�
Ĕ��"��i`[�"F���T)&	f��1���|�d��TGjL�A@ۉ!JCȱ���"�y���\S"�ưB�3�	�\v��$� �"pR$��ƣ�t�Id�:��`6�5&Y���3��*v��F�����cR�)*,����QDd�-���칕(�")�l�	�I�92太�����U��'��klR7��z��Ȱ�,�5a�*j��d@���v&�Ȩ��Q[*"ƴYVX�X)��PD�0iq�Mg��/8�Or�LȪ*ʌKa�<��܁�#��� �F]��DŨd�u+��^{^�Pq%��19n:�=�̨
��g-ܒu:�'�c���I�Ba�d��tFD���2��"*���I`J<>R<.q�t����Ņi����PB��uW\p��Ƴ-�$UV_�7wi�6W��Q�EY�G	��!&����Z�خ/M�'�Oo���.: ޲�*�eXQc�v�x�jBE�+8��j�ۡY�z�cN�9�60��E$	d��Nn@=�E���O�j�3k���n$�������c�J1�H��U�D64���� �hQT���k"),2�`���>@|�����7���<8bF�Aa}!�T3���޴0kyً��9���;��q�,e��$�N/�
���p���i	�-�j�&��5�1F/N1��!�eu�6��q��4B�n$(=0�쀳��(��%{r{ss>ty��+%Q������n�S���{�d�>Iܚ�}�$�ֱ�T�z���ru����q`4�噑<��c��<�Z�c�2#��Լ@��7)���HnJM�Ξ�܇0��]3�V��y�*�7�=�����ܿz���ݠH	_3��ý��@��Xq2�1�����[�����om_ko��ƫۑ������W��_��_���UqiUU�*��*��*��*��x�ګ�U꭪�U|��U�Us�UU�UUu���^*���ZUWUU�*��Ҫ�W��W�努�����U�U�w|u�������UWQUW�UqiR}>>�I �g�|f�Dj3�qq�����Q�KF�E���D &�)U�hX�i �JR&Ph����||���*�j���������*��Ҫ�����U_+�U\ZUW��Uz�j��[U��ZUŬEUWX��U�V�^�J��*��*��ҫj�U�UqW�UUťV���b���J��W�UuUU���'�'��dI�
*� �mck��F��m��"E(Y�h��(u"dB��C��0�H���Z�:Ҫ���U򴪮*�UmU�W�Ҫ�����������UU�*��Ҫ�V�[Uz�*�����|U|�^*���ZUW*��*��x��U�W�Uu[���z�ګ�U꭪�UmZUW�Uqbσ�>������� i��+_h�)�\��������mU��V�W�����J��^*���ZUW�Uqb���UU�UUTUUu���^*���ZUWUU�*��x�/UmW��努�Ҫ�V�W���ګՊ����⪮-*���U\ZU^�ڪ�V�g�}�3� }UR���c#A��
(bA"h�R��u(.J�J�$+�4@d��d�����Яr�@���
L����?���/��@T �Z������E_��?
����3�~�?�8C�`D �B"xDGI�"%��M4L:'K(A�A(��K�'D�&	��D�MD�8`�"'�0� ��"X���&P"C���"h�2tO	bX�p��"A8"'�D�D�� ��"'DD�,R`���8�,���BA(�YAC��� �bA<P���F�i�0DԔt�D�N��"h��a�:YB!�Æ�#R/&W�W��!ᦘ�����)ir2EY�B$�Fx�CJm.,����
���P�- 7e�R����ܖQ)�d�C!JBA�p �B� ��򦐂%"(�QYd�X�p���(+ 1AcU�BX�8BdU��Q�j�2�[*)D"���Bv�D��K�Ĝ(�E�)\����!Q�	�T�
 ��4�2 �I���bD�F�B�,̬���VB���K.B��)14J"� �B�b�bt�(�B�qܣ1		����P�A���&�B9p��yG&�4�:A��*�6EQ�
��!��Q܆"2���
.��QlX�"�� �1�AFA�u"�!-��H1��hq91�:+!H�cPd@�c�(� 87�A���(�� �S��IQ�C�� D)FR��@��֛y	)-$&�%��r���x�h� ��MZ��YaR��@D������)U�VFVЬ�x�2�ʪ%\��B��BcU�Q)V<HAJ9o-��2B�Rc(2� إG4{c�6LDnT�ac%ȁJШ6��Um,e-�XÈԢN��7�kk��ѵ*#B���;v�=d�
c �qABX�(�f]�&��i#*+�K����(W,u�!F�dLRA�Bɗ]�&)!Ȃ�\ȁ�m����ȓplR8D"D1[7F�G1�u��,hPr�9P�![Mʫ�Cd��I��m���x�<�J��CEX�j�a%L��<bT������BH�r��t��PO6���#HO ���R�L�c�[.F\t�Yl����i`"d��R�/��PH܅c�)��d�Dё�`'.%�
���#)B(����ʇ�y�ZV5	h�rR��tHT�5c�bB�h�aqRR7$��Е�Yi1�"]Y�ق���D���	���A2��"��*!d��]��ʺP��VU�����\���H1F�N	��!L���2�JR`�+ ���<����Qd�ʲ*�RH����SA��,�c)D���D&,DɅ��i����%�JT6)V"�*"c<nR\C����Z��b"$!n!�?���jV�)	8\� �.9�F�Pa1���Ar���r1��c!)5q"o`�ˉ�FH�C¹7"�cN!�Ȇ�1!�"�c���#���J��1���Ǖ$b+H��T��2�:R1.L�b*���L)�l�����[RcI,��2�,Q���*$�#�@��H�$F�J�1��P���(�Ʊ�G��+
B",PH���	��F�6	юV�0��Q�\�7�q��㠦5�*��d�`��Y!	V�"\����m**����EQ7�q<�Bx�caJH�$)F����dyf:6�%V)���H��j-&V�X�(K��Q��Ԑ�e�`�p��h�<�e��\�K�l��u�LR�ȡF}]�&h�ǐ���I�H7.9�b���	�v���E�c�`�(�Q�I]�QF"��!H�BcqB���ⴤco%���* �n�p�1A��h�J��Vi���18�0�~��!�=D4�D){������ꊱ%���m�$���B&5,uX�B��keX۬�K�ȇ!R����-�	A�-�����\n�F�S+tRLM�4$�J���*8ҩT4�W���5lQU�5�)eqԤ��v����2��Ļ��L��.d$LU$[B�ĭr�����͘��8�vZ&؝�\��P���UT
�$�buE�%��:+�dՖHQ�FД(��n�b�������Zn��[r�c�����Eq(�%����)]��DB�ݴb��K+U���țMYQ-i̭��ʜqU#jQԛ��5�7c�8��cu�(Ae�؛�H�h�IQ&ĤQ+!]n4$�U�KD[J9#��Ҳ�� ��;^;j[
�ln�1*���r�"�ʣ,,�UU(�"���jE��������X9�:��*�ձE"UD�j�"����
�1�+R&1��'ZN�b"cM�aQ�T!q�X�r�nEa���ڒ)\RD܉JZ����;N�tR�	�,�
860�$<��Xۭ�SdT�iܖĂ;�C��?z�A	������(�*�v�V�q����|�J-�!���֔N����(���d�&L��`+*ECq�]%d�bI(\��#�T,�1U�ʛ���d��$���ʥM<N��c)��X�lQ2FEcQ;H��8�ɏ^T�R�!S�U�����̲�er�$u"��TN�B<J4I"e��#�A��
�[���rl�q��r�	EZ���S����l���H[J%b������������
X*�8H��Ȉ�Z���ʛjei�&LM2�*I�R�!�]QH�#��Z�u
J䚚�ږ2W%�*4�,��TV$ڎ�ڮE%��U�g>�(�}��7��X�����UU�ԁCHB�[���w1�fff{V�����|}���Ub�U]EV����}��}��Ub�U]EV�����3M$�M(�L<"&��D�8i�0���:x��G`�*R�0c$���"mBD5��`�H����UGʊ"ҕ"�B+��&�if!QW��j���&
c��l�D�P� q�Ӗ���	G6�b�.%EP�<w"˔�ERc���!Y0ll���+�2��Sm�Bi��舉T�!��qJш���ˎ�cJ��Q��:��D��&(Q�<)q�n;bb��LQۖ6$V˗# �,��T	�1��㪏 �L**�22*�Gr*�KARڠ�eE�1"�4�V�#I`�"�Q��T�Ȇī�X�X�9�����B�X�I�̢e�d,$E����R=o]�¥d��9��Uj����$��H&�j"U��k���"���R+T�F��ʘ�h�+#�#�UUR�;Sj�E��I8�$aF�)cI9#Ci��G&�)1K,[����7d�"Dmڭ�����%�.Wcp��c�R�Gq9U
"\��vJ�����$ĚؒIn���=1:G�|S�çN����~:^(��k�<�՛�4|fÆ��Uh�8Cx�w��Y�,e�t���:{��ڼv���<��w�������F����[�ǵ{W��Ǻtx��<B[���"��h����p�-V)����(1:T�~ΞZ�����ԦF)KUQ��k0��F�4��ff s1�ή�B�Qh ��\L,8X����T#![��u@IH,U"�l|28H��G�p�"Ra�4}��t0Yˇupb��X��PV" ��xX�A�@t��0�	>(�Ř"h�'��4�8_~�EQu	��6l֣FVVY�U\UT�3g��g>'n�����w�̎!�vbt�˘\�1~����ܔO6I*M�q����(�I`y.�:jM��>��E
D�O1�(�!�p�l��7��Nsiy�C(���-��_\��My6ή�1����cC��ѽ��uI��D�B��:�x��ῤQiAќ:I�M(�D���&���M!���=��I�wn7j�5��$�.�3���A�0�Q��kF�r��lV����jC*x����k��p���rs�Sk�wy|��sL��qb�4��	7ѡ��ss�|����u^���ה�ns�,C��!L���P�ы��E���C�p�д�(.�U��MX�d�� m8s�F�|<�W^��a�(�p+�6�2��@Q:t���Q��<"&��x�(�Haㄮø[E�#�1��g�/9$���I#�Mp�E��ʳ�V���Ute�P�S�Ɓ�O����S��(��[�Ya�6�u��Q�.��E���2��̘\��n��YJ꽪�Ԯ�F�I1�%{�5�I�����]LP�5`@�|W�ԣjZl�aѹ)�IC4����OǄD�4O%i<@������p!���γ�9�td:�Nӂ �mE.�blk�!�C��ż��▼*�5����h\I$��x�x�Ȝ(�	��d,�Dˡ�X��2���������y��}�w:o~;xS�l䇰�Uv��sڏ>y�iV˲���N{e�|�$��T��Ud�\���������d�����a�l�����������u	Q--�7 �kzy{;|�ݓs�Ѹy��j�HL�8p�T�l+#����)��5�����h��:c����N�;��Ă0�A ��t�Q�T�2�H+L��E	���jū�87���,19�l�A��k���N	p���4� ��>n�)�Yj�tE|��gd���Gnﶼ&�+�Md�T*�t��6} �ag�Y���4O��h�0J4�xỦ�p��"s�IS4f6�l�@ƗE"��L�2!b�;��<f��2��UEI5L���]^��A:�Y�
�V���<�]#�e8��(�*5<��d���8RAA�;{�$LV�D(�7�Yw�������=���>�vn�л;0�F,�$2������<Y���~?	�4Mi<p��0J�12(���m��$�HӈT�j�"ѷӪ�g��ϲ�Bmdf��
� � �Aߨ��9d��zq��>�N����t�0�ب2�j���E����<OE�oUxG�M8�r����Q��EgX{��r����9�qqH���U�9a�ޚ����yp������\9�Y��v�~K����V�V��
M@�CC�b<@�4�ĖQ�����h�`��Ha�{�D�շ7�&��'S%�:�ߒI$zba��ȴt�"bL,Qd"E��f��� ����?<H�yc�`�OZD	�Z��J��m��3L�W\t����"���q@\��<�,�/�1������B{�����XaY�Y�C��.��/AC��L�<�L,�7��R�@��WM6YB��"^�Z��C�N�,�D���&��hx���&C�< ���8����1$;���c`�8��BLI!\{�dQ�;U����'9*I$�p�&:s����D"��:'�7E�}EB�N������;Fp����h����Qr���&�����5��v��:��H��3��r�ߡ�q��}�S��ϖ�g���ᴜn�vܺ�s��}~�n��x��a�+��4��
�v\ i�A���m��P����pK5*ج��N�BI$�'��0��c��tvEϼ�ي���z��D��E4��V��
:x^,m��J���f� ���\
��f�����jOsFڮݺ;h���>��\N�n��`�r�,��0l�Aa�a�3=�n�)���	%Y'�4�0�4M��Ha�.r���T��9��q��5�V�9{q��pq���P������F�1��VJ�	]

�%����Y�i� �v�hy����� ������y+��U����D�'CEh�UQ��]]:�Ѓ�WF�<50e	��j�>(�K�Iy%�T���6ҴԯP�R����;��)�Jb���]8�~�iHd���อ��p��z%%�tg��f�Äpf��!���zF�F����N�G��Y�i=$�6�٤h�l7�����=Ꝟ�y�n.�d��/n!�֍�[Lњ5ўA������eA�/[���xz3Ɛ`�k�4���h��4k�h�z<:i:94���ӄ��z=$�4�,���G��z?���$AC$���C����c���0��G��z>��|Y>-�����f�q�����4z>�F�A ��M"M#G����a��^��'�q���ַ
�ÉѨ��ooN�vsrvz�qےv&�C�c5�i-���>FI�M!�i���~*ȖRD��&W�~"i84�i>�Q:l>f��<l7�����=٤X���l4��v'�v��v�n�󗔽��2HG�H���g�R|w�������O�;=�['��۞�චOΏ�=�N_��}w~޸'7p�U��ħ/��?�w}P��}�d�~j���9��{��&��'}��]ryU�޷��6��2�=&`f�raG{����+��>��w��;��No���]��wv�߷����"\�yΣR���u��y��z��l�@�n�x۬����_r<�F�թC>/G��d&
'�+�Ҝ��"j����� �v�>��3���f�����t�̙���BG��{����df����M�ə��4���W��n�fFff���ݙ�����^���y������wvfg}�<xg�x�Ś~?D�0M?	F�0���0��TTV����VY�GbH��Z��1'l�8{-���Z��ᄃA	��K�B��Є^�5���Eu�6+��Uy���5���*����sύ���5�I: ��C�sDgb
 D���i8:b��M7c	r��8R!����QЯÆ0�clr2tA������r�|Tr�d�����#��t|2`r8nhu�����p�9o��pE&�qӇ0���7� ����̅"�4��_3����}������	�j��(�`���'�R@����3��a'�||Y��O<Y�ƞ�� |kR�ƭb�[�TTV���lf���|�����񓡐�\���̓k�<��4��4b?�"�KmN٦i��7D�y��*ft���|�Dnq�����z:	=c�ԁGT>���<LL��A����#�X8����=���F�9$O�^�y�0�'�r� �L7tEUϑ�9@���j\�����k��]!D']�ľ�����;q< .{�����.���	��N �����V������f�<>�r�+�)9RC�v�V`��,�~8i��b��4M�������B3� ���>E��=�,9��S��Y�����3R�b��gPjs��N��]R��WH�*輊���@��4l�Ә$����(��jgC�������A|���=�S�7�ӧ3:Y��d+�sy��i�p⼼��>G>b�/n�e��Ϗ�ׇ=��8{�<}'/�C/\ڗ�b�r�SWS��mM��L���o^볿�ӽ��!a���f�hnp?��*����z8���N��t�ǌ{� ;!"#����pg�Y|El^�9�8P!�e:C�����&q�Jd&x8>hd�!�@z���C��M������L�����ˢ!����3F��[x��2N� .����00+�>w�C�	�`c��'� c&���9���\y[M<1�$���`���qd/1��n<ah���*Ir�6bil� �tGqΌy�4i�r|�41Fni�FE�@���M0L�<��$� ���c&�Ɠl��h="���7B�y�G ��Qјx��N�i���4M��O�a������g��{��&����ޑQQPHQ+*L~$hVd��M01���X�P.&��Ѭ�I��G*�4�� r�MW�|AV��ۉ�@��(|`2<;>33��6!�"D�,�\X�@i��la}c������0�u/A�>a�����o '�G�R��"G~�j;q<	Mt�/�øO�1^�#��}n�'�)���)�+�Pi��jg~�z̓����G͠43���r�h;$`��9g���������(�y��L#L0rA���ǇX#D�w�]-|6��%�&��(d�F+� l��Һ�A%lVJ4L)���� �XIC$�'Ğ���xDM��H~4�x��b̻�6�H���,O����������ʦU8V��}�@�2�1t8���)��)R)X+4�ppA�HD��	q7>2�{	�����]vn޷� R?m�Jw�&h���R4��a��aѥ� tHD�a�v�3�	��k��6A��v`�fN����������@�����G̉�h{Pa�`�2�v�v�+ӆ�Zb$��%8 c�M��R�S]�+�����q�Ja��62��O�,����:��X�ˏC���HN�b��ӏV��ARQѢ�t�zd,h�d��
d
�������8xgǉ?	>?C����xDM��HA�}��v!`��4EAfd@0�S\9h���$(����J+*+�5�ˈc������L:�@h��������C�FÐh����)��~&���Sb�5f�8�<"�:OF$�� 2_�������a���b�0l��f
�[
��[8]P���l�È���M*0$0a�.-�T�J,��Z�)�,�C� ������\5��� �w�$�@�n%���Q:^�eJ��;�[���5� L0Σ!�))4I���E����),jr��V�=�f��d胞(��;c������`@�ũ��be2e�i&�p��DD�44�~0�A�<1���C��4�lE`�J#�4���
q��z#� ��-9�p�7�pcl.��Q��M5+l��u�oF�7Iy����EEEA x��r	�N���h�� WáÒ��5+�3w��Ȟ�|���ܻ��7��v�)L�~��'��bY�wǋ�3N�/C��2N����G�e�r��웞�ɦ��\W�ջIv'�Eٿ?��܃w��(͛�C���]��c�im�
�F9�	�������!g��=�3�# L���z5��F�jNG�4pu	F�0�g%go|��I����L��3�G�i���@��,�ٌ���pJ����?�F��3�iņ$C�0?��Da~d�9L̳���i+:����'���P�J�t�F���%c9ץ��ȠR�@Ã���Y��=::}pLc�� ϰ�NH>�D��v8c�����Yv����m�<!��M�2�e�t8rD/
���i�"Րr��C�<�:`6��d&�O d�B$a'�x�O|'O��<"&���hi�0�a��!���C��3���!��{͵ߑQQPH3�{��|~�+�!�40v�:5	�/aF�x���.�$ta�a)c_NT��ߠ\��p:��r�`x`=P.	�p"�����ŋ��!I���!H�����a�D�B�8�G���C����e

Y�ƚ:$e8%��o��/��9�rp��n��.V�۩.M�j��8�|RC5�HI�K+�VA�������CF.8>�N�1�3�`ry4��쏻b���1�8�S(w*i0��8i'I0����fa�0M4�� x�uϹ�7�Z�z�]J�`l�{�{EEX���S����
�*94���P�4��k��n�}0�4��	w�@T(�x)X�)1)���Б i�g����Ǐ.q�Έ ���:�Î���u�7}�o�:�+�=v�Xu�2 �!��#C_+?T�.⑨l��C�xc���oc�Όv�W��O��	BS�{٫�)�>L/�q�$Q��l0/
JD�0��El�� ��x0.�P�R���Q�OЂ�BI"AAh�aGM����j��*��I�\T�@��ڠ���]��4Æ�?	���<"&���hi�?�rd��A�>������-�3��c�H����`�f��~�Ŋ��@H��tW��P�Q!�
 ��N���fh$�ָ��x�L �|_�
��恢[��s7!�Ŏ���O�	8~*p���)���H���t0�w�w��]/�Ev:.�R�R�XI1� �m�)��Y!0/X��+���>�@ErEj����&jP�|�MP�GF��.�H�����0��A�0x@�b��ME�&x�D�+~@"U����4�F�p���(�(p~CZF�I��i��O���J�h٤h��e���I3L��x=�Af�Y�X�G�c�f�ލ�͋���]�v%�v\���<�҈Ti�B��g ї���:<M?$,�>�C�	�	�	4��f���H��#��|4�=�I4��F�G�4x=:D���҉��=����z;�њa3G�HV=��[zAc��eá�=4�?���O���0�~���ȁ�B4z=�F�K#M#G���zA��GM"�e�Q�*�J!��6^��~>886����*��/���%숗����ٻ<K��vkI��=�	8i�C�0�xG������8#F�#G��/&f���!����t��"�pr3Bv�p��.��OK��b$?,�d��	�O�.�&"�b�D|�qc8}Ӥ��!j8h�i��{��2�H��aD"������t�ל"8|#��<����p�`}	�itb:$}|iFy��Nw�G�����uiǄ���?�.�I&yg�-d��a��e��'_q�xd>�ru�a�؊TqP�:m�՜��#�?%��O85;#ǻ�/��yGU�Tھ�L���w�g~8�~�5#�!�Q;��2 �9��s�p�z������e|q9�f�,���5yk�߿h���U~�!�־�}�;F��w��л�w;w�n�_��utߪ�a<�w��u>s}/�(��|��;G�9z�S�r�����s��T��]�3�1��UQ�lۙ���_r�-o�6�^45�n����΋�w܄���.%��ȖW$�%$j<��D�#i1(D�Q��r�R���e��c��CA�m��dR+�U�Ge�q�;Lm���k���UW-JG"���5ć����������߾��3'332�绻33��������W����߻|��n������U��b��w���������^*��+��w���4��pӆ�t�~<~4DLCM!��ϳ�,�	�_8J�,�2h�D���_��鮃����LP@�:BC�\E�	�,-E�0��pY��V(X"���(,+)��1
�H�&!���"RX;����iڈ�JW2�`�B�B�Nق(�+�D�A��|��[F�ͣ����*KJO��iu������i�dD��2�{M
�Q�ܫ�"b&��Q�Lf�A�d2�+<� �+�\Ed,�+d!U�,��JZ6�X�iv��AIX+
�Z�ERh����"w!	=���DBR�1�*Lc)[G���PHǍ��GrYK����O�V�(�����zR��Ҫ��,�����e5f�u�;�J�[#F7j���%7jmT��W���*M�T���)�-Q��m�d��-��
���UvI\H�l7ZJlqJQH�CDCc�՗uV�X��4�U7i{-ov��֤W�ȬF�6�I[L� �+�y[3�'#�1��!|�\�Y7�C���L4���RYç<���hxk�NC;s�Q�Q�p�U<��'���ۖ�;xS����ӆ���?3y���AǸ#����Nwם���e�f�*���9��f��'^]�{��-6a^�s��cֻO�e��;D!f�s��!=�4�eQ����s�*4I�d��3�0>p�1C�����^B�*Z�1i��")y�t���0i�ǳ�G·�ٷ�ۢr��ߌl8!p6�<��;t8:��T�H����}���e�&L�GqݒGC��Cɏnq���tlp���4��p0p@a<��q�'}�`���}�F6��ӡ�Ȏ�"���y�ӌ>!��oJttW��o��u�1�]H|h8 ���N�U���u'"J��A"�Lz��W	q���b�L�����J�X���@h4|���`������M�����ZtO�H��pHa4�O��8|if�&���hi�0�a՟���I |}�����c�@`l!V~F'l��O�y9�t ��4bp�z<�P,VUФ`BA���jS8,g�.dy͎���Ko�f�ì������K�e��x�U��R��Tp�åp��Dw����K�b!|�KӍ��U��+ʔ�����|��ߤpmO1"^D��&tQA�BtZ6<�ð���&p���Tf�29�I�����t;4������0��]:�	��a�����cL�t �!h�T�����815��F���5i��
����H��A�i�J4��<a�0�x�Κtg��p��MBB�'$�\@Ě�����M1�� m��w��2�q��W-t���&�\�v�F�ǃ`aJT�����s�A�`�	�2�P'o���6����o�BHVX��ʅeYM?�'��afPh��߂����pi�����7A��:���u1�1�49���Ƈ�� �����է��x�֍<;9D��?�cC�zH}=�u���t��
_u=|DU�����?0�z��fx0r����樧Opzö��Ֆ`;|g�9 �[��T��5`ҍ0nE����@�m� �ϙ�'���s333��|�{e�Ǐy63�N��K���NĈ9y0v�l�8�fݛZ2��f��Fh��i0A� �,N�������"`�i<~��,�>��ӱ�c�H�c!�?.�:{C�^�g������]N�n.ߺی���2:�Cpl���Cf�i(�#}��8��Q��&��.��O"cC�<���X8�����7�C��l4��Y;:;���qH��M#�� 9��:�����ހo@ǆ��.�M���
a!Ʉ�����zc�8�*Up�� ~�����9��n��=�c��0�``�ImӾ1b`1�۷c�H�L��.#<2�{'>=�`�ᡍ;��4v8.CA�����Nbǋ��a2< Be8S����?���&���hi�0��8p����d!Y�w��Af�R���i!�sm�(�5B���
��JCW.��*�"����}�j&�i�� �w9��O������:Ә�QO�e<z��Job�GO{�{��}��l�=�Uߎ.ܿVr�8p�闤��K�Ma��hP�zC�7��;��p*|�����o���9ҷy�����9=��_�#\*�"�s�b�ޭ�}�m8��_��^4�;6}󭚫�r����|�1yH̩~-x_,���c��40p:�����d��`������ǁ�{�HL�9H8����xt���;M���h����]9�azD�Ld���щ��O�\�yO9���"�_oRn�O@vA�$���p8σ8y�t�h9%'3y�ptE�1�lyd��{u�a�i#}z��rz��R�C��8x�����D��P�O�s��#Y���۽�q��v�Oi�+�Ƀ��A�����D���q�ͅ)YCw�yp;��Ӑ�H�1Ha�$��G�<i�O�4�a�L<<#��~�g��?D)/j�i��� �S���m����|��9`w��	�h�R<p���E�T����]�T��1\��:�����3���%��L�9���f2�!�,��a��t�臖S]�C.�95ɏ!ӎ�ya=LbY�D'�<�)@C�����2χ��P��'C�=2D��^sO,��`�zw���.Kw�������:;)O���E�|r�d0p�-Б|�� �c���8�����rg�U����N�p4i��> �g��o��������p�?!�lzg�t�X����8�;u����:Q�(�Ni�0��x<t���t�m_�IxMr\c�0 �}� ��m��n��VlW�լm�^@ì:0�@SR^R8.,�n�CۯG3O	��L�h;z�(_(��X|���M (a�}�6�EF��
��-j��\�A`���>?*�-�v�����\�暶K����g������զ2�5���9 �V��pf�ЬE�rM�O�gR�j ���947q�~�A�f3��q0�3�3qfA��LFC�ly|�#�����O�k
X��ұ�����gx~��e)���5Q_N�g8lm�^=3�8�PG2Иd�AH10���^R�0ູ"��u��O��-��������AA��K0�,�����<~?	�"a����?�Q���p�6�j՛nZ��1%�$�M4�M4Fc1a�?����_���%z 9��5�M�7$�P�g�9�5���)ќc-t�g6��̼��M��Us����sB��Р��q@�8�{~�N�1���62=N�ǎ����r���Ǧ����h�|x�Q�p�a{�g��q�\9 �zߌz[Φc��ߪt��S_�҈J��)���r�C0�-�#�>NK���t�����t馆��rD�&CӶ��������><�h!��=�|,A���������!�:�����;`�hw�Ӂ�A,���b���x�~DD�4<xgM?2͒	4���I%TF��@���NBV\G�n&A�?&��Brs�Tl�n��r֥�P��]��~j��i�	����&t�{ك},��o��L���?��[���������6��1�O$*8"���r�����|�xz����՝|z�s��ns�:�l]��w�㖷t��^�s��N[���R�V�6���t9#����О�˫��|$�\�_�j P[|��G.�(\kB�Z5	�-p�E�A.�u�~���P���H|3��0vA��~kn��<0�0�x8`�Cl�6A������ǁ�{އ��� �����Y�p�-x<<�r�C���g z�+��l
{e�#��rB�`~vI�3�����R]XA�� # 샑$�tc�x��0i�N���C�V��4�tK3�@㏣d<1�	�1
_u�s�O���M6�����'�*j��kZ����Û}a�s�8@�X0�.�c�,z��i�:<hyt;�����8Q�r"�N��YG�8||Y��x�:a���4p��iK�Q�K�%f�t��+L��1��0�hnWo.M_t~p-T|)A�'DC!�Π�'Gm�٘�\Mu�Z.)�[P+����KJ�x�DyQS,q5�a��b�k��G_v}�\8��u���3�����A6)��"�WV�7[�8�t�|n&����uK>츙�R�]L#���H0j�t�i̓��8��Nǣ��50�38 ��?�"�E�8�p��2x˦�V<�h�5E�Ʒ��×��{����NН�1��4�a�t��A��В���0Rq>tX���E�	Hй)���ۡ�:��i�@�x�������r���l��㋣��9���`���ᆌ�Tx��8iC�e��h��zl�#G�����8K �4�6�N�Gf���!�6p�4za��,�3�${��iЛ�.���\�؛�4dFX�������h�њ>���z5�H����Za�F�h��0f��Hc�H�����8if�M"M#������z<�1��rI6Q3GF�h�f�#G���[viFt�=!idt}��c�Pځ���EF�G�4�*G�ӄ@�4�4�O��>'�����#�H�[�,tYސP�d�q#҈��D�E�n$����/H�bI�.�Fh�h�=��������ҡ��#��d=8LF3H�aɤ��vi=2��=�B���s�/9�w��iЗbn��NĻ!ۉ��a�濏��Ņt���?��z�������fÞ��Ӟ�I��:�<_k�I`�����'W���}}�w/�;�%���7}^�z�v<�Y��sZ��d�Fn�f��y���_}Y����r�O=��g"a�3��󈨿}�K�ݜ_5ryt�;�����bo�5��M��Hz-���_�g��6��^s�M��o�������|��{�o���sI��_�M'���E��n����'��+��9��~�Z�W��ۻ�߷ww{�������Z[�ۿ�n���w��UmU괷����������j���V�+yU�/��G�<Q��4�M0��ǎ::C���!1����1Z۫6�vKI2��Z+�ӌ?�!�����qތC��fƑ ��EJi_=�p������b�P��>���C���bvz�$R��	ŗ%�j������SE�gE�QR�}J|i�j�Z��9���x�yv��2���!��:}����NS�>68:$�p���6A�@Rđ��VÆ.;����31Ã���2T�\�LS�
0|;���ၤ�%̮�pP�R<��(�fE��Ԃ@��A��"��!#$KN���Ht������ǡ��2|�A?8���[v�c�ݎ�y;=+���wC ����<V�J�P�O�p���~���x�~DD�44�||v�IRLͻ�FfCU&�H���&�~�����ǖ���jP�g�`�H[��+P��b�� �pERb7�%ӳYX�o��t��l7�R��7y��w7J�H�S_.-��՟>�.���,e4`�8m}��n 莅���s��IÉ��4Dx�$`���=�q�;�~��o��m���zd#��gg�!<rB�M)u��<�q���8@��L�SO����d}"��%-vƨ^<�m�C���0)t$R.Yуf
�Z.��S۠�����¸y����C���n#�P2O�x�%Q���><~?���Ha����7<0G�Ca�t�/��Ώ�u�	h�N�9�nU;��: �����|�=	���I
mQ9���QQZ$�
�����|�L�af�-�}FaW����f{�}����҄2.��fy��ŝS��I��Q^-��W�=:BWQ�s�ԏ��;{�1)��>��pӗ�Q������g��mkCkĹ%�&a�5��$X�V��/�[�vF�q���v?c�ӱ�3l#o�tf�a�C��|���[�H���qJ���°��f��z����"�Q2k�٫��d-��l$F��T+텕»���<.�{~�h�㑠�5L;�xs��0���({�>�p?��3y�dRĒka��课x`�>��0���z�;��nݺ�?�Q�! �
�,(�aY���{��G��O�a��xH�C��t��<6�I��
ו��&�xp$�H>,�	>,��4馚a�t����:h�]�%
������QQZ���UO�cL��Qj��b���
��o�U��<��!�qA�!���(�H�~�����F��^��XϹ'��T#�‰��c<���QdظX݊`�;ީ1RA�kxyv���0���3�O���LQYo:�,΄˟C�fS7=�%�  �s!��ng2����d�:l�bƠ[� ��|z{�qؑrrW]�O���`_���]U!��
 �
>$�'�4��N�i�a�L<<3���oXK|_R�,��v(�x��%clm�А��
2�u--�ߡ�)�K��Ѿ�>	�$D���L \�!�:�b��4F���F!Zg\c�̑�OR�]��x,>R��8g�у�}g�v.����`������T�t�9���j��ٷ���C4�h@�y�<{(�����"�b�T��D�T�е�pB�gL��@��j��()V2�+K��R+P
���sҐp���l�
Jn�·�����-h@x]P3�1JR�΅��ɁL��?�2���:p�Ğ,���㦚i��a���ӥIL��H�(ϻ�TTV����RBZx��X�Z�ȗduG���
�����
<�Ph�)L<�Q��|�Z��6�H4G!���uN��,mۥa�Qj�\�l"#tX!���4F�>�ã4$^��"��|�i+EA!�Z|}#U���a����t��"����c��8#���PE�tR��_~�8*Hy=*;`h���C���p;	JT$�Ɣi'M:Y�M4�'��&��C�B����(,.�h�D�4&i#���sHB��]i��ݪ2)*�d��Kr�����**+BC^�rYޏ��t°��&�8f��g���ʽ�r��z�c��I�ۯ���r�={ó>�
-=�U����_+�]k״�&�~�7��7��{��S�����v�1���%J���_%}�ȸox��b�Y���]�h-�*�W�4IMO^Х�3�J,�p3�pD��O����m�A����0��Z��.}��X�D4�P����O_E*�hj����g���XR�H�+�&\^��V������J]�B�w+�ӂI$+�A��F��l�����3�(�=k��~�	CEb�U�Z`�a��4�Y�=�e�2��
;.��D�
SV�T��/-��v�H�P�a�Z�؈A6�@t�H:|Q��	�0�~?	��&	����Gs�	!����h�۔E�I��H$�.#��|����$>�>d���Z��	�
���+T&��A�K�9j��qqqBV/j�Ã9!��*���q?+^3e��f�:��|cҟ<y9+ע��UZƸ.�)5J���R�tg�A��R���ܟ¼(��e�VBj�+�Z���b�,�\���"��	���B��υ��JNs�N̸�D<�e�D�=�ssX0��H8t�I<|t��㦚i��a�N��q�r\�.����**+BA��ۑ�Q�⃊���v�������S8e1rd�,`�?�O��oqpT/�P�]�d0�Dq�n�իL�,�IEASC�����!i6�Ħ��\٤n�/&�#<�g`>
�h~/�IѺ\��po� �\��Z������@1���^MZ��b�i.�ɩ�O�F]������:Gp�O�W_к��K�T�K�Jû����z���E;�܋AJ����	
:3�(ҍ4�g���M4�M4���ќ>��ݩQ�ǟ*p��*ʃUSX��2�ڱ��oq�����	��a��v�=�;��DG81��#��tG��Q�r�_t��hqS2T|1�� y݇\|�b��/�H$�Ѻv{�Ƿ���������~�q@������l=C�k�ัm��b���̕�(�`���x_ ��y`l�h���@��F/uB��C�+E�7i�A��t83�H�5��ޥ��	l@ã(��?�CeG�c�����N�G���a��4�=�I6^������ޏ �a�<B޷vr�'i�K���؛���c��kFkrAM��
���8=���f��ѝ4��H^��i�4�L ���G�h��F�F�G���pz#K#FN�8=,��F�ñ����N�NI�h�f�Fi�0z<���iGm��W ��h�>��f�H:N��#G��H���H�n4z=�pi�I�>7�h�4�0���4v@�	�,�L'ĳ�����<]�'`��.Ľ"]�{���|G��|F�p_�tlψ><3	��&�����'����������A���ӄ=�6[��l7��7��m�p��G��h��L��7bv%�vK�rK�	>1:|5ь$�h��$e�B��iN3�
pgC �A�Hh�A�b8�B�N�y���>?�!h�8Aep����}:2�]��GPzOz�m���e9�!��r�e�{j�)��>�<E5K>��њ��:$���{Ii�
���������>�Δ�o$�:{N_p��xpg
͆�$D4ǧvM/&�J��%<�<A��D� tbqȦ���淶�l����=<��W=�]Q}���*�a~�__%��*�F�\K8�O/�ȋW:����~{�^��}�y,ͮ��[7%T�[W*��_|��^/�2OG�D6�3���U�i=_5�-G*�g������D�L��Yh�]jJ�q)*�x���o��MnUH�S�v4'oҢ��Qmi��Q�#f�s5�G]n�$�+h��G%�H�E������;�(z�L�5u�=��wu�V�^�K�����������V�^�������������U꭪������������U꭮d�V�Q���(�G�<x�M:i��i��::2�G�"`�l�MQN�,)F"�2R	����خHQ�[`���B��p�toť`ĜB���\�t�
:n�1Q��� ��H ��;idd�x���KI$-�J'E�dQ䥃#U�ȃvjV49Ѱ�!ji5�Z��1�n$��ȣ���苐��Q�b�%�D![�
�Bw��xF���VIS�$p��+�^Bb���8�$��F�B�S*���TA�6�R������I���I;���+w �:#�X�r2��B(��0�24��B^\F�%k���-uV[�X;J�I"f�Fi�7��T�!e��u�$�֚�CV\n�I�[6���P�EBm=Yq����8$*�D�D'H�RD����;biar�1��$�M�;K,*�
�N��X�d����!�V���ݲ(%X�H�m&�P�L��M#l���֬d�F"AV8(�jđ&V��̲&��K2�e{j**+BC�����I�;I�f�G��x>S�����^y��I��z��u>��馕�u���K�D���_�]Qܮp��ӝ��K7����������7��>9�Êq�j�V�H�u���_8T�Oq�������Ӹd�7/�{��\z�IcLg��T�	\2��B�jj�����P�!�6��U@��H~�~b�u�O�>��O����m>���o�Bb��:#�&c��s��N�0��s���M�M����Z_G���ױ���`Da���LXŘ	W+�g��g���a�M��޾;��q~�¥��:T���Z�p(g��T��,���C�x��(���4�L4�N�!���!+�n	8�/.��o����	*��M�@eh�r����g��,.�����}.E1�L��V�W`�b�1����	�E�5T*�|	�4
E��p^�����:\V�u3��8}�!���n����0+W����_~p�^H�}4�����q�KV��|@ܜ[*��}B�A�*�dj�@���Q��>:i�M4�M4���і�F�[� ����q� ���"�6����=>=�G��;"��|��:�<�:">N�c����	�U�^=Ҹ�l��J�IR	�2�#���̤U�Ɯ�����?�p�Ꙟ���㻵��·OIy7k�6G�_��B�cD��%B�0c9?G�c�h�����\0S�i�o:<����Bm�W]�Q�����\'s�&O����~���8"q��}�l��x�F�|Q�>:|t�M0�M:t:te��~��U,QDX&�RT��cQZ71`�#eB�_��d$ g�4�o�����tTj����)@pf��/)��DLJ�uV&�c�5>��h·|�
E(�|��u0���#B�.H1�5a����^����"� (dT~6�"�H��jv�&��;���OM�c�蓑��v����;�SOݤq鲾q8Fh��ݸ�い|3��0���}}��Ό��(�F�pӧ�M4�4ӧC�l���C�4:49�q3�����vd<բj	�H��K�x��IV7S��y�|���А�[�g���M�9�����D���������d�=�x���M�gw��(N�g�6�����יZC�$zW������t��es��3z���k^i�rȵg�U9�������z��鼃3��}:�2�#�C8r��I��j�bO=��iRK�g�2L��t��z<pr<��w��썿_=7�AB��R�E3�Vp�t-�����s�	���G�o���KDI��Mm6��^�t��>U�t<�
5PYj��,���TJ����A����=�e%������B�@�L�� ��<$�z���f�>��.��r�"�w5�i����}�`�)8��)����jO��J�.�P�� ���
��"�,&Ԥ��G�Q�>:i��i��::#��
��8����O�TTV��*T�E]j�
�j�D=c�Z���ؖ}Ts���p^�_�?��x:#�?����Z][�rH���3����r��(g�k�
˂���(��Q	<���,ʃ��$R�$f ��f��+��}V2��R#$�hD��"��(��E'x��$�X��"Ι�\A�?,	5�a�MA��v����Z!�V�2r��"pY
�!��2�B�|X:]�XA#<Q�F�a�:|t�M0�M:t:te�巳3�tr�L���*}��$6��,`"=�U_��]��a�H�p��6;u�믃�4;����桽(=�?uq0�����R�"�\E� B>!Ã!�
R�
��gt��6���%����I$���F
�Zo$]��H�R��%`#�������^���X+�c:>�y!�a�GV����2*��#&`��|�+/����<>6pФ㷧��]�@���������x������馟>><p�p���,ah�%�[.1����!�aY_�	ʁ%6&$h�R�b�-z>���!�>9 ��d�9<�"�p����{{x:+o�8��^Go�M�����|0�-XX�]����FR���+���R)xP����>$�DT�S!Mqn-��B�1��/�vK( h�xX����P�TՅ
_�R�ļ,-+�/-
��(:pe�$�ҍ>>:Y��M4�M0���і�{��cΌ�"�g�iq��hStBf�HT�pTќz�jbr�&�źK�)�,�\2��C�b***�&=՝�z�Ȣ�.��)p�;�`����;y�#+5��&+����o��ټ4��gJxwK��$>�z3�4;��>�,G6�[��]�X�{�kIrw�������l��BurryIE�ow�~m{�ֺw�{��M�:�i6�[�n�m�ɛ��AL� �&��`m���Y�4�o��A�9�Mt���ա��ћ��3Y&�x]Yab�uZ�pL�c T�Э�(�)i"t7��:3��t��๢�A��ߞ�X��X��T��8���V۠ް�%#9�q��AC�;Za��s�܀0�n��T.(G�^^B5%M�p��B�!0ļ@� ��8x����M:t�M0�L:t�ΐX�6�4�l m�%U��U��%� d5�b**+F��1���>�����UX8�Z�����^!]��8�8�uDz~�T/k��,�08Ż�tVVn���B��H9GO�+��p  g��$]\�yx6ê����~� �&I����Fݬ�r�Z��4�KL�?a��F���dΊ�
J��CGFP4�:�}��+h�WV����kᒏ�`3�Ⱦ�,]X�.���Id�(ҏ�$�����0DÂ�DK<"&&���'����AA��rD�8%��<'��0M �&��`�&��h��i��"	�YB'�"a�H'��DO&��DN�����x��"C�%���"a��(DK�x�!�h�d�!g�J�Q�8%A0CAD��K<pDӂt��Ěa�<i��44�H4�J4��������:XP� �h�A��3��s`����֭��NOyX��s��I��X5󍕽�KT룏�8}~=sY�;����۬K;�+�;Ggoy���;|$���ٳ�S�ﾱ$��u������6z/ܬں�9P3�+�%�.�s�۬�OP�7�j*�摮�u%��|v���y�9��u��l�ɭ�ڦ=�q4���^�S'g����*fG����:ʒI{��}������(�W�}�F���k�U꭪�����������U꭪����wwws��U^�گ���wwww?~�U꭪�w�����Q��8x�Ǎ:iӦ�i��aӧFt�g��kH���	�}ߋ���2UIZ��!�('����yrl#��FX������L���cX�RԩJL$g�+���ڲ!µ�� �O:F�!�� �1�H
W�����Y�9,��#粥�%�t��I&{$���1@j���ׅ+�pe�QW��������a�0q;"������rQR�ZV3�Y��p���u8��x����R�VC��I"`��=��R��,���4ӧ�N�i�i�N��8[k
��B!G�V\�c�ʢ=�1�7�f&�t��xsAF��rĐ���+�Ԯt�Uz�z�lt�83¢��4G���⵩�F]�`�4��������3H5H�D��д>Z�L��CZ�p<3���H�8�.+V5MXP�Rq�)�p.�{��t��pF����0,,8�b��ac-+��GB���><�dc�Y����|����59>]
���E/�h҆�b�	UԬgT5����M������t�ㄜ>(���O��4�L4��:3�8t8SX�b:�ZB��њ2hR�9N�
����nH��;
#��T�((�u�kclm���e��(�YF��#���?�a;�f?j`wOaw}�2ef�w�^j��r�z��?��5C�gOn��N|=�o	��;�p����>D�]���]������(�M�'5�k�\��FQ9�p�xɶ����+��׬���Y�Y'�9ωw����9���ϡ�:1	>���y��Dv����eO�D|dn��:���G�`Ih�xZ�t$f�W�X���bl���&�D�{b<�Y���$�8J�_d�T//�^^�Pφ�T��@If�`�Q2�"��I����m�IƄ$�A�a�0�ಾA7U*��4WNR�eH�]��	$ei�NQ�L:|t馚a��t�ѝ ��QRI,�t�R��\Y��=TTTV��l���?c8[b6+`��qzt�'\�_>�'Gc��::��̉���;�J����H|�^�#�jk�ϑ��}	�.�ſ.�M�.���B���C����$����hu����ϾDU@g��_W 윢���%Z��O�F��)4t�b\0]<��ZA	����>1Dn&�O��C��à�p|Vbq�84��X��7���Ձ$�>$��4��N�i�i�N���r$�f$bB����Z�׈���	�ʕ�wwWv�߫��¯.��
-u|@ފ��v�:��:�1�b���
R�T�a�� ��"6�l,���W�A���+�>&t)�1�L��M]�6|7�q�Lب����g�V�\��|o�V���
 `Y��.-_BʂOJ�" q�����|Y�J����Q�����-a��+�E���3�$�ei�O�:i��i�:tgH,;�B��,�1e0�h����'J.�P%h���UfJY�23W�n"N�ĪH=}tz3ҿU����p �RE�괇��t���U�(�{���/��|�ܡM���Zt X-Mx,��)(^Zp(���ǎ�p1@�����a��WHx?Kad��n�]&t?ip$���j�h�RB�����04$��:
;�
��Y=V��CBE�-@Ŋ���,�K(���Ni�0�N�:3�YG
d�@�|!ADC��쀑Je���Q���r�v�X������F緤TTV���@�=�bh��p�{��Å�dA��Y�:���7滛��:o��+:5�gN��!Dq$xߎ���V�p����a-��W����X���z/�������R�a�N��+9��w���7�=���9�Ϲ����fO���2�[�҉h�_������A�jCEjR��"�`�HupѸcL�����81=Z-2�!x&���lmr��Ǒ	I��@0�Z���$$P��Fb�|.������Q*T�2��f��A��~2y曎�5nۊ��!~�[�ЈH�k�l�8��ˈ�{�)�1@uL�"�N������~}������,�'�(��M:t�M0�L<t�Ή�7�S��4:�K�Iq]�# �kO"���&WŐ��\5[�C���0�Z�ӾO
j���PLWI~�t?��p��k�BjKi]�X{ƞ0ngEպ(0褠��-eP2dF"~$n-�v*)4p^���ߔEU�O,��x����kd��=I,�w��\9\"*Ë��/�ZPP�����cz1�w���KB �߾��y@Q&��֛���y!uu|RxHΐ|x�K(����N�x�L4�:3�4Kl�6Ū���F�j�Ow�m��Л5��צb���s��:/�[n�Z��"����Z�h3�jC���|Px����^\u}+�h���ЂQ��jA�� ,ՋD��@DD�!�ؒ��L��Y��,(P 7�J�7��[X��Nx,�0�B�A:1��7ab�H nƝ�0V���A3^F�$�L��x/�>:��E��4`Y��=߸���<I��|i��㦝4�4�ǎ���o �dq~S%���H �Q��∁+�bw�!_و���	�]r��kE}�����tl8��I��s�Ӣ�&"JRJ��:|��~0��h�feQ5��d�db�T�I#��q&!$.g�m,�(Xdr�E��<�8+���թ��GW���:���
:`I���96W)�R_/o���⒉o)��-j�ÉE�N�"#��/��8Pa��p���~3����4L(A�b"xD���x�G�
AA0�8p��'��'��&	�	�M�`�&���`�t��KDO�pA���xM���X�8N���:"X���&D�&	�8'�M�O	�:%�K4��8%	E� �!�A"pD��O4�et��Ǐi�� ��Fa�a�i��i��x�8HA����������4el38IӇ�QG�FoQ���iь�B���i�ш�B$��� �(���	d�	��KNf��d6>�ey���]���)�ݺn'���g��'���e��$�,:�nAG�|O�E����QB�~�h�O:C���4��h�i��zq����̸}�Yy�ץC�u����O�黦�|oW�D{>5����F�����(o��CG'H�1ȏ�R�d#6">����h�#���S��L����W��Z|ϗ+^|����;ν���W�u���w!�����z1���O����ϧ�B���s�����}3������/!���n����c�Ƿ�Þ�ׯ��|����N��+�\M�	�R��MI�K�ܮ��K%�WF�ܱ����bq�ěcݹ��lcc�)E+N�)�J��%0x����wJ�h╗��+�ufe;7���洪���ww��������ߩU_+�V���~�������*��x������wwww�����^*�ww��>�HiF�pӇ�4�a��N�i��a��Ft��o������!�������!�I&�<CY)(I ��c"����H�B� ���()!�"Z�2�!���
@L�,��h�[�
��"����ڙUq
<u���2�N��"I\u(�ZYj���;V\RB����oF�q8��R'Q��V�C��Bn�L�$ �(��d��;#ʱ����#p)Ip�R�X2��L��(2�2�$�����
��+�d�y�A9&G���@���!2��"�JWq��H82
�72���%����,DE�I���JME!M�T\q܄ɒT�I:5�2�,�ءH��"BF7nL��A1$7J���7��b A7���N��U[����j��r4�"uK]#�F�r\��e���\lc)d��n�0lL�":���JيY�E�,m:QF����J�;8ƪ�Dʖ4�V�#Q��X�"�$u�epiU%TBph��'$JHBHԍ��DIA����(�#H�xՎ
�]RѲ�9m�����k�iT��#%�-M�|����Й�gs�8C�������ؔ'g�ae�0y�;�c���f\i���9ߛ��'+4K!4�I�!��x�>�^��x������r;#<�y'���ٞ�%�=��<99���sC#mQ�r7S���go�9��<��l1�sw.���z�Tꈧ�[�	Z�՘�j7sNV����B-��uK�N�?H<,R�А��xl��!gY�B����s* �洁�V�X�,;|�������r����#��p<�Ưh@����|)�iHE 8BBǴtf�ioV��q.p�x�P��n|&���@�
��IdD|��i���� �ğY���M7���L4�8C�l�BS�dV�6�Z&)�SugٴTTV��!�`L�٣B	2��<b1*P��ܠ���X��R��L�(:P�t=��EE�OQ�Ӹяε��೽R�X�R=>�Wgg�����yaN�qIL�V�BN��!�G����Z]��+Ȃ��Ȑ�pv���iֹ'�P�+�q���єJ��Rq���j���VXYBŇC��J>��������p&����2I�$���O�:|i��4�M<p��g>62R�BE�%I.+��QQQZ+��T��	���
��ǰ���L�\��!q|���E�WW)�O��B��ˉ|��!q_;�KxAc<sĘB��kZ�HJ����'
>�V�?x<�������>{My@�Y�R��5����zJvtmݯ(��	)�m6�h����R�R��$�"���Vv+��W �)gB�I��t�N�x�M<||x�ӄ8&�U�l�$�v9x����[��4���К+�4pi�ȗ�h�X�)$ ���
�A�9����g	"�S�]V�C�F����ͳ�Η�k��!s3�Gpʊ�	`5�ƪ�ٷg��-M�@ԇI!�)K�z�������e�!��?�&XfF�����ݜ�l��61����0�����5@x�4�L���Dm��!f.����)��,>Sg��3�a&x��M4�f�a��t�ѝ ��,��IC )�� ��
�(2~D(<�T���#sJ��t��5�5^ruA��N����%��+��'޴TTV��a�ܹ�ٕ	�x����O!�u��=ތ�Ga���K��9O�O�Q!�Ü9`�nx��G��������]����ga����=�D�,���9\�����S��+<����*�9�༌�։(_g}좫�����TL˖L�,Z�/�*Xt�h�Ѧ�B���3�4 -�џ���v�t,���G��^�ꐑ�i�->�ґ˟� (]P�X)z�]^���Q�[��>��bD�\-J],���p��!t�%u�6�}�d`|qW�΁��t���|$�g��	t(�tg�<C�O���i�N�a��t�� ���X2>.�K1�R@��	J�WP�Ԛ}��6WJ�k�ĕ���8T���G�j�D��,\�uHA���/Ǌ��9�m��3�{���n�]����5"�j�֫V�,%+L�
È%��c��g_��g�3��Q))bY�Ij,y�������쩣;�v����7\�>�pcn�:t���oWE�
�ѫ�}����}#f� �Kdt��0�4�Ɲ4�M>:x����ӫ�"~U�Yl�R��cQQZ���	�Ҍ�����9WG�DA��x<,��taA&����M�f�3��ezw(C�)�������Κ '���J-I����p���c�qWwA�X��i�0��(oO��J��q0��cv��>f�uf8�V�\�<:�G�H�+�f J��S���y���X��p�tો�$�<I�L><i��Oi�4�çHtM���9ua��C=�����'B�?n��F	�J9>��|):6���*�$�h���jHq����-���8ʯ�����ΊT ��%�����K1T��Ⱦ�p�y�,P..CB���,����LL�EJ�W���D4$أ,��pѺ�I""BE/U�H�&IV�!|δ?@ttvV�G��ՕW�ُ�=9;��A�2H:p���><i��Oi�><p��g� CGDHBB�P��h(�3F*~�A�@La��B�'ަ�$�Ns��'G$UU*D��$N����X��6a�>��oAv	>0�;OH!e4�y������6z|p�O����M���������w>��1��Ӟ��q����Ow»{H|�ϻsJs�:��>j�s�Ϲ�YO����þf�^_�����bJ�̗��<�}�8�v�p�c-�ɵl4�|�d�ŀ�5�@�\V��d�,޾�6��.��ϕ��t4�b�㲺G!ÏS��ԝ?6YjB#������Xaի����p^%|����Z���&*��L��&��C��
�8m)������\E����b��5ū��p�t� ��9���|'�4R���i(��i'�Ǐ��i�M:a��t��a�7��A]ʶ]Z�N󈨨����Ғ�T,�+��:x�o�+U�{?G��|� ǎ�!�o��0��a&����`<�%X��ՙ�Ǡ���r��p���ƮJby���p`\�g)oM�i��,8[<.�-
	]Na��t�����vp�S���9x]4��w��-/,ۧu�Yý�2�@��A�*@`ub�p���|�Х, ]\���,$_�t5sˋ�I�"��d���φa�:|YbYe�� ��""&��"A,DO�""a�:'D��!b �tJ(C���8"tD�d�0MDӢh�D�4DD�å�DK:P��&�D���%	�DD�ı,K8&P"B�K�0�H"%���&�xN�a�:B�+��8%K"H �xD�8�tD�L0�Ex�GN�x�L4���C��b"xD�?�<~<~:p(���������A�5:sN͎�������<9g0���9��+���vE�w�7�ե5^�]��7�y��ä\̫���G'>��i�j/F�<�a:��i����v]�G�o��w�=Q�~��1�·�tNr�w���/Wz�F?Z����󦬦���.�0�x�O���g���9�GT�����&v�����w�a���{������9;�ﯦ�z�~����s0�o�Ӳ��'=�;�=�_h���b�w�UUťV���~�������UUťV����������UqiU���񻻻���*��ҫwwo��4���i�Ğ<xӦ�x�N�i�<xg����b**+G�R@���*�]�9���&�a���y>�O��0�)t<��:]��_�������.v����A`�F��П�^X�-�3;��j1P��?-V�F�O�0��c.)��� 7���N�b�>���Ůa�����P)�x�cT�����>���>o��$���>4�0�L:x��m�Ʋn�5.�(��oq�NN�R��纊��є�!�J�%!��b�T�F3�1�kG�v�0�d��t�|�%�]��ev�˾��۟�Ai�/�����KF�q���%��z>����̤2<���>p6=�~�:W��~�`z�������qo.�F�����W��΅��Ե~��ꘐ�p\�|i�>)ԟ0����c��Moɘ��83�cvI��i��ƞ4Ӧi�O�8�}��(�M�bc!�H2A�Q�e�L)N��X���4��cn*ԪZDR�H�!%[�wh����9�e�DC���C�G��~lWZ3�;���z&C��҈�4����<o����+�
�Q����o�w���ßr�|۝���q�;����|�L��6��g3��a(HTU]��G^��W(�s�!4!%�;��T&��8Pj�g�""C�(X+��EЮ��x2O��{�^g<�ǓPd�6�σ�4`S8_	����LZ/���K@���$Ꮻ�.F&���>�,d �"Q����
i�۶�z0Ղ�b�"�Z�X�8!�`ǁop:X�"��&�i��t��ƚY�����!�ܘh�vz�L�F�(�������s＊��єg٬�W�]sʏ'�h�^��͟���Ť���B�b�U�p�"W����(�J�0����Д	�����h�Pt���<PETi͋Ԩ�j�^������9{xtx��zuz�E%%�+�'h{���ӱ������|�yk�b��3��������d�o�N�|x��i�M,�M0���<>%�e���H�1�:A}�����p���el�����؊��5���)���ރ��Ŷ����E)T��4�Q�����]׻S�r�!7�x����v.�:��k�B���\�@�A�F����Za)��fxJJ��x�����!�3�ŉI<W��*��,�49�'�UК!,.����)X}x+�2H��$�&|a��Oi�M4ç��ߋ�v߫*}Z�p�]�5>�QQQZ2�_�qP����)^yxV�U��t!����KK��C�!�	��Mf��Pˋ�8���w;������x{���?=)�p+��G�F���LI��t<=��>���isJ�^�P����e�d��X�?NRʗc|�W��J5��U�WU�ǎ�,�t��q�6�V�1��ĺ�j���>�@�#�&x�0��ƚaf�a�ǆx�k�C��A!��ѐ��*�G!��4��c�y�Q����p�kY�NoW`T��7���Z�Y*���Ee\�v}�1QQZ7�}�ovo�3�ag���������L0�*�L�=k�wy�F<����E~{��K��e��e���ӂ�7;DY�>>��F{�����}Y���p��7�G7~�^�$藯<���5p�w��SϏoT����{�:>}�N���%��g���ɑȞL�Q.��YŢ�V��łk��T�""H��Z�q���4�m'qh�1X�ZuuQ!�����S��Qþ���J�\$nI0>%"���ش8��h�?��kP�30��ӡ;���U����ci�tG��I�b��d�;��\2�uŊd+�Rp!4g�=d��R���|�z8י�l�J�Z��2����N�Y��x�L,�L:x��m棕-�3v]ʶ˻��Z**+G�~�����c��Ӱ��2J��޶��{��H�R`s|\�.�/�DGW�U���5��g�^On��q�,THPy�5�܊:�0���_H�|7�rv���#JFV
$f~L!�0��{��MhME]H�y1wEO^����|���A�C��U������\(_t#�upT,VH�#���	:a�ft�������!�ܛқ�,���ޝ[��RMJ�{�"���f����T�&�f���J굂���Z�h���Ν�!�DU{t0����Aж�(��rz�t_/����%��u���Լh6���j���Qƛ�s�7P�s�"HX#o���w E��m���j����Ep�J�����=2�Qf.�ǡ.b숇�@�:/)������>L���wN�#�����(xI�G�Y��x�L,�L:x��c��r���a"�Bq+�X�co�?C8n���������<�Ͼ��"��K���FH����0�b3�1�N��ϙ���9e��8Cd������56�|
��Ac�{	���S 6��i;��`׺z�7Q�hNk��%���3��yj�)��ձ�g�O�,Y���4 P��a��W+a?��vxL:i�t���4O �D���D�8P� �tAġ8pD�8P���i�h�`��h&��h���	�J�K6ȐL(A<A�%���4�"�X�%�g
$��dDD�<P�$�D�D�0N�X�C�!��FK"H �xD�8$<%���(�:a����O�~����X���h���tN��$��Fhhhhhht�f��~���t�DR�D1��L��t��!�;�!9�!D2�`���/N�c/g
CMd"���H��4y��4�¼g�i¡��xw.�Js8s�4���w�g5�����ny��)�O��tB�������S�}��Q=������"�B�1aHʊ�S�}��{��wHw����>wxt��E�^<�Fm\�i������a��f铆��nT,�Ǽ7���a��HC�} ">eA
 �����}��|�M�ݾq���������9�����so���|W�r:�moy�59����ۙ�뙮��Tw�K����+����\���{%W6y�rےI�����^���4{�9=9�O&���Io��Z�'`����KvثM�ے�KI�㩫D�2J�v�#�Z��I*�U��	���բ[��X�m�u�F�ą�RrG[v�,�Q8�D���*�	���%qG�¿���_���?����J��ݿ�������U]b�wwo�www~EUWX����������ߑUU�*�wu�����Ox�Ǎ,�M<i�i��N����(�k��F�m�1e!F���1�aQ:�H�"���$�cŔBL��	cCK!
ȱ�yK
B�����p�TbJD�Rʲ�TDCbl��2�HT&�LyP�H)��X!�����!�U��M�Wp�x���ŷ�DU!c���iV��ݸDY�#�V:Lc�p(�FPU���ʣ�\���F��(q�Hhز�C�$+��5�K	�\eC,��!bl��"���`�."���*�)ih�1JZ�,)�B��B�Q\������e���e��r�11�X��&�i�X�- �11�$�DD��K �H�i(G*#e�����,mF;)*$qEP��b�����$�6�H$TA	Ñ���T% ��<�&�K���Q6�e���B9F�3��Sb֪�-i&�je�ܢ������"-���$7SJ�����e�ӐR$�e��\�ˎ7#�:�,c�Wv[en[��������?���5��{�}ț��^�ӧ7J�t��Q�V�=0��#�1���'l����=���}��N��~�(�}�6�gL��}g��wt���˨ʜ7c6���&m�����a'�������{�s���8/�>O�s�}��M}�")U�8�X`���b�����఑��k��<���x[��y|*b���|�(]!o�x����>*J*�Ì4��u�-�L�O������M�>;��n��d�a���ի�>���Шi�Zp��DA䘄p��/��~�Ҷp�z�w��'�t������
�	�VxZ������ q
�a+�`Q:t�	<Q�O�0��ƚa�M0���<t�ӐGq�۰�y9�r�Dr&��w��O��Ȣ�����~���gEtf������H�X*���M�ֵ���|sNVa���9튍7CK�x�N�trT�c��À�.	�R�����N��+g9w������V��Us��˃!���)�q��Qp���5b�Q��G�Ч�a*�xTU���p��i�2��>$�4�M4�if�t��:I�0lk���c��3Y�qE��U��0�N"r�p0j�#�V��`s�jE�M��Ȕ�h`X�Z�R�g
C�]~�M��9 �H��D�|MUAT�°_/�O'�k��C��GEk��wN�x&�/,��h�؝.��x77Aa"���{kE×%*A�ଋ8&,Pd��l���PpP-~�,0��,�I:Q��4�Oi��i�O㤏�au�Ǯ#5fu���.{�(�����{_xT�.�q�1�x�F��a#4�P��wuk�1�#$"$6+)�2=0�E�}"�%B���8e(�Oإ`AŊ慢��a���+V�*PXp����qq�`�&$�1I�xT- ��R��ܺѰ�l�S���Ib"��"V���*įL�L�\�P���"$�'J:i��i��4�K4ç�����`�'��D�����0e?X"�q���:t�6غ�Ţ�M�ڢ�ql�$Aȣ�t�����OCą�DC�}��z!�i3��8�#�3�9�L��t�i���;�� ����_q�����g�7��#�w�z�'tZ�t݇�.φ|Q���	}/�7�/q��ݥ���Bޔ�����x����Mz���������n�-L*��qu?���Xt,V)�=�P�)/0�t]�����+������)ҁ���S^#M��D:�*M+��Ö_�y}G���y^M�X!�:�s>	I�rt�y����(G�ȑZ�I"-B�A��T���BJ��K$��<igƚx�L4�L:x��$�p��d͔��T��kFy�!!,7�/���`�qG����_V�8�}aai����w�QUV�^G�t?u��0z�����:�x^z�EQh�c4bl9�΂��p\�� R�$��i��֜����s�4Z��K��:�����}>���J�ok"((<�p�x/
�BDa!�ʽ��U�6a<�ֈɲτ�Z�N���(#y<����!�id�$��M>,��Oi��i�O㤘��6	$TC%S��ܩl=�����S�!2"
���͒I}PR*��`�4]Z��FWA��tQ2ô�g�ZZ�´~!^�U�ؽ�Q�q&�<��0����2��Ç8������ڮSHF2n�-7d����$p�_��8m�h�B!����r|Vp��17�H�R, �Kఱ@��4%h����+E�R��*�i[�u��0�z�<u��L�z4�ñ�v�$��t�	>(��i��4�K4L4�aý$���PT�ɻ		
I����F��1��X��br�!�/���ix,��c �XH��#<�����(�BgNswk�����}"ғ���y`R��`g����w�մ�)���o�XH$�m�Y����ދV�v;|�{�t܇F��1�2�ԑO�.��/����Ux\Z�r(	R
�R�,��MXp��a'ĝ(��Śi��4�K4ç���	�R���c?3�N�pYI�4����6\�	��<"�Є/<�&X�ڊ�ED��Y�ġ�4c\�G.��llm��Y�<t��|S�
k�/���f�9�,�&��=���ܣ|	�
޿WV�y�J���3���y���ɇ�%������ʙ�η+���&�;{��3}��T��$�ێ,�s٫�^{�g>�Y���.�j���&� ^E	���k��A�'�x.��\������Ux��efp>��<}?�:OW*������&�\^O�CRv��C}~
0~�����I�X�`yyo�C��:�sU.��Hs�I|��3w4��w��A��p!h��pi���d����$�F�ag�x�L4�<xg��U�8zH��5E$q��$�K�!!!,:>&ߤ$)Zq��5�uq5��L~���2���P4l�WLѳ(�Ml>�)@��U.������lgl��ފ�g�K��ij�dM��Bp��P����G��=�ɤ�хr*���9ƃ��Z��pY�^P�>�a��h�F�o�P��r�m�Ȉ�!�)[��:.&L
��R�|�T./��dY�
0�Æ�tӂQ�(���4O ��"'DL4D�0��
�A�'��D�8"Y��M4�4MD�4Hh�&����&(DJ,DDK4C � ��:"a����:%�g2NA� ���B�H�b";"Y�h����	ϒB��(�YAC��%ܟ$H�a&A��N�:t�M0Ӥi���tD�DM��:p�ƅX�3GZ����+_�)�sq-�'}��բ���UL��uG����gɶk\�����l�G����-��ɰ~R���.�}������"���7w4_s��o\x�.v�(1��|���N{�N9y^��;g�;�rM\Kv�|׻��g=�a��q�y�:�T>�Mn�ܫ~s�<�ʊ���w6��'3�;WY�u���+Z�;����ɧ=s�˙�a��zyٶE�܋�1��6ט�^|D5��9���}�����&��R�s���xN����h���Ϸ�����}�������U���񻻻���*���V����7www��ª���wwo훻�����*��*�ww���Ğ$�G�Y�4�L4����!Ӆ��`�#��BBJl��Ȗ��Y�W�}P9Ml7]�ީ�6�a��	�]kG��X�\<��H+�4+���,>:1	"����&��.ݺќ^�;�$�hW%6�ƐDG*+h6?�2��*���^������C~<�-�\%�N�E��WTH!��{��GE
��&��4��4��0馚a�a�ǆx�'
�%Ǡ�f �&&�m��`�b�Do��跡�S���Wmvs���O$d�ˉ��HR��E���_g�&37.,��)J��g��(_-&�8����O��|Ӵp9��ϗ�۫}���Z�����E�&���ǃ�"�}Vd�s^�"!/`C
]�XqM�
(fId�(��4æi��i�O㤐x� �a��JE���� �+rช.�M$I10OF䞨��,�F�+Z�9+�Q�1+aUt���m���dlfԗ'����pS�\��=�z���3��U�
����_�<��xJ�ܓ�syOxt�9�nļ�$�[��W���Ԯ.��_=�ߗ���:3�x�&���%��eD�iH5��s�0����R��T)XZoE����|�ڤY폦e�G�s.,�������M-�M�ʎ[��Sw"�]�P@�
4����v׾�����X/����Xh1qR�wF�AA��(��Q����9�%���g�!2H$j�Io8\�kbW�sY��ŏ'\r��Qz�����@�b��4�(0�%�aFif�t�M0�L8t��:C�3���X�fژR�}�$�	�;�:d����S/��fa�9�o�c�����������rB
�WE�C�eh��p�W��M=�<�-��ހ���#���*�6��x(GB�+!s����|#�!��"��xGHj�o/9Ҝ뻻�%�����$T,��D>�\]�!�t:,M(T�Hb�_0cRǙ����l���>7JR,w��>m��&`�(��<Q��|a�4�M0��ǆx�#T����L��몪���u�j-Fh�,�Z�������e5z�p��x}^�����J�̦C�脘��yBfPXH��H|1`�ۘ���jdɖ(��[T�*Y�'$��x|��A�ñ�p��<x߈�]��#Š�D���P�:�c��v����l'�����qѪ��'è�qA���p�'I:Q��K>0醚a��p���<t�Dj�S7���:�UG�c����<;��h�kEb�����A���y�<ѥ�kst��z#$l�i�2�C��,Tix).(�7��l0�p�ptE�Q�ǈ^T�C���!akU_N�L�=)\"�\H��j�S�:2���G#܉�ڗ L��� 1���Р����A�3N�a&�i�t�0���:3��x�'��A�!��N}:Q4�/Q���)R�;č��8"���tĸ82$=�f��ɝ��AK
H(��׺��$�Go�v�Ɵx�i�l��.>�G��؋�>z�T?{|(���Y�g�O;����l4�3Y6|tgt[���f�>w���H�K�{'�h�l�i
3�1qҥuj����f#�;��K�gl�*��?�D����k�<��}��$���!�l4�vM��|bş·��`Ϟ�O�d�	z`�i��P{��bBI4�> ����C
����<p]\�m.���p0�Ҹp��|���Ū��M���Ӱ���qСp)tX�R^K��T���A�KDQ�x���cٻ���m�����j�W�������0?����0��|a�4�O�x莜&O��w���+&��x���m���/
���h�V�u����˔X�H�;�N�~��A�H�ڷt:*8�XԪQd|zaH�X��a+��h�9:�gٴ�t����fe>ɟ4GO�:Q0h�J�{;>����N�'%�7N~���<%�B��M�^PÄ+�p5���-���=���b���.�L��"b�=xv�qa�#�%���ǅ�ŊV�3�<I⏌>,4æi��4��Dt���|�Ɵ��,�"�fTDU�A��$�:iރ-y��~
�b��M�(D(��:��6�����(�M(�5�(c>�uȹuB��.��h��T��j�E���@t:���ñR��k¢�+i[+�~u��k�M�MA$N�T!:B�_4���o�J�E�,��$�&�j-3�̏�T"X�	�RB���ʓ��d:l��g�<x٦���4�ǆt�FC-˒eđ��!vkRI$?t����5/Ȓ$qq?��$i�`h|ag�	x�Ft��%	&p���1���kU�9��x*�!�q��IKBNزK8Yͳ���\\\E��T��C�H��;\1���=�y���9��|6��h|Q8MpW�k�B
;�L��D��h,1Z���E�tK�k�O�Ț=�0�ն�����?���O����\?��֮��	DD �N��x���zLc}u�P�R%F!bD :�Z�VX�-L�)��I&Z��)JI�JQ%)$�R��*Y��,S)��S$�L�)L�)�L�)�YT�YL�)d���*ܒ�Ie,�5&��)��d�$���I�)I��[2��iK(��d�I��Re*[4�YJIK&J[5&J^J�%&J[2Y4�&K&JMI�R�,�L�JT�^<r��JY2d��Y2l�i2Y,��5&M�-��&�Y4�K%%Ie�&M�&��d�Y2ْ��d�Y,�K%-�&MI�Rd�Y),�Y2l�2Y2d���dɲd�Y2d�Yl��7&��Y2d�6�-��&�ɒ�dԛ&��
�2Y,��K%��d�lɓRdԚ�&MI��%�Rd��5&K%��I�Rdԙ5&MI��I��d�dԙ5&[2jL�dɩ5&L��̚�%�ɩ2jL�[,��&��d�I���4�&Sd�d�e��Id�Y2Rd��%��)K)$�ɖ�I2iK&�&Ilɴ�M%�%)%��SI�%$�2�I%�)I���[4�L�M%�R�&[,�)4�L��K&[)4�L���*�d��eR�%&R�S*䶹Jl��)2Rd��&�ɤ�i*M)e�Id�RI�)��)e)I2�l�$ɤ���iT��&��e,�i)%2d���fJRL�R�L�d��,Z��e��))Qe-K$��YK-K)d�YK-K)dɓ)e�e,�K)ijYK,�,�,��YK*�,����R�,���YjYe��U�k�efԬ�S @�0�
@0�&0�"@2$	�C� dXRZ�M*@ʐ2�#
@°2� @�02,rlӆ�bH����)�02�(�°2$�"@��@ab��@���
@ɲ�dRQ��`aX 倆 02 �0�*�2# 00¬�ʌ@�@�$
@�@�"�� @�$�0�"2�
�ʰ0� 0�0��Ȅ)�2$ @�@ʰ0 0�,�@�����$���(00� 00ʤ���@���@, �� @@��R�ڕ5YSj�*�"��@@��q$Ie�*j�5eM��V�6�T�J�R�P��HR!�a�!�� ��Q����!X``aHdaHaHdHadRP�FBBBFBRR�!�a�!�a�a�!�!�aeHRE�T�Q�P�P����T�G�e�a��f1���B��,�2�,��Y�jY�I�B�B�Xfa�Ra�a�e�a��a�!Ba�a��R�a���VYe�Ye�j[L�e42�2�2�3
H,�,��,��5,��&aI�F�B�B�{�Rfd!�fa�a��a�Ha�a�a��Rk,��,�ʖYe�Yf�$!�ffffRd!�a�d�e�Ye�j�ie�Yha�d!�d!�d!IY�fYifYK2�Y���YY�R�KL��)M+K)�,�R��YR�eiJ�RT�eK+L�RR�e)%2�R��Jm)e2�))e)JV��L�)*e2��%,�R�ҥ�,�����YM)eM)�Ă7�j� �H!����,�V�SJYL�*���eKJ�2��2�)�)QL�)L�)��2�)�K+M)e4��ҥ�ҖRV�K)��%K*T��2�R��2�R�����K+,��e))�Ғ�)�,����ܥIL�R�%2�VR���*RT��*YR���J��JUE2���ʖVYR��ee�,�i[,�e2��,��T��R`!�a��	��Zѻe`&0�� �T�����V�)JYSJYYel���,��Yee���)[)R���J�J�T�l�e+)R�T�fVR�ʒ���VR�W���VR�)JjRV�R��2�*̬�EIK*�Tʔ�)�)je)fZ��)I�L�RŔ�-JS)JI�JY���Z���� B�v�'�3�e���qN\�������EA`�E����?A�~������z����g��@t����s�W�?���W�?����$!�^�}����?�]�����B�_���(�����G�g�#�}+�r7��I�p�������WE��W�?�������'�	 �@~�ѱ�?���� ����O򂀣��I��a  ����*����ʵ��꼾�߲���W��z���$��W���G_�@p������G��X����@T �������E���t&��q�?��	t߽�~T��a���`���bb�;�N�\q���ߏ/Q�jz��d\��נ8M��"_������{�����$P@s�ѡD"�P��Da�TVXEQ�Q2A�D�F�������"(��y��_������$Q=N?����<��� ��PJ!Q� "EU	�� hD(�U������:�I�(���eτ��u��P�'���D�ں�����O�|�*�?Q����'���R(�������ۻy��* b~� �#@~o������v��o����?��q���������G���?c�� �	�;O�)��bC���#����?�����G���ߡ��V���
�濲F���V���3��a��������	�)T �[��@�?G��	_���?�d�8���A����?�\F���'��/�H�%��_��(���TG߀co��'�SO�((���&���?AЧ�D����a����1�?o��S] ���Z�A���jZ(���B\G�rk�!?��E@G�������������yP ?_����2t��� �y�(������������?�ph�Ѥ���#��_���q��/�;�������$���6���?���	���P ?#�ڟ�p������}�X�TX��Qb6-�TlE64Q�F�-c�Q�EE�h�bѣE�Q�Q��b��Q�Eh�Q�Q��Dh���#�"1��b��Q�"1�1Db��F(�Q�"��Q�1DF#Db1DF#Db,Q�1Db���F(�Q�1DcF(��b������#F(�Q�1��1Db���#F(�Q�1Db���#b�Q�1Db���#F(�Q�1Db+F1F(�h��#�F,h�F(�F,b�EDmQ(�h�cb�4Q��4b�ъ#F(�lE��Q�b1�F���(�DTh����QE��Q�1b*"�6���Q�(�cF�*4h�DXѢ�hƍQ�F�64h�F�4h�hأŌc�1�1EX��1�����EF**(�Q�b��hآ��QDQF1�lQEQE�b�QEQ�QE�lcQ�QDQQF,QEQEb�(��(��(�QEE�*,Q�X���6*,QQQ�llb,Tb�4Q�b�����X�b�11Elcc�cc���Th���(ŋ�Q�j(�F�1��h���b�E��b(�Qb(�Q����F"�EQb(�b#b(�b#b(ƌDb#��1b(�Q��F#1E�1b(�1b(�Q��F1���Db�"(�QE�DF"1��1b1Eb(�h�1F1Q�1�Q��c��1������4b(�"ŋ،F�"�b,X�F1��E�4lF#cDQ#b1����Dh�F6#�1Q��b1#EDcDcDb#�4F�F��TTTFŊ64h��4b-�Ɗ-(�#F"��F��h�(��F�4F��lFţ���"4Dh��F���F�(�Dh��(��4Dh�����F��Dh���#"1b"1b#�#DF��"(��"4Dh�4Dh����"4DlDh���#DE�"4Dh���#DF��F"4b#DF�Ѣ#DF�(�F��"4E��DF��"4F"-#�,Dh����ѣ6"�#h�b4EQ�Db�4Q�4Q��h�Q#Dh�Q����Q#QDh�F(؍�؍���Ѣ4h�4F��4F��#cb4F(�4b4h�661QDTF�4hѣF�cF��F�ѣE�ѣcF�ѣF�ѣE�4cF���F1�F��DEF4TcF�c#ƌc1��ƈƌh�h���c��1�Dh�h�hƌcF(ьF4hѣ111�э��Q��#1���,Q�F1#cEc��F,Q�1�"1�1Db��F(�Q�#�"��"1�#Dh��F�"1�Db���#Dh�Q�1Db���4h��F(�Q�4Db���#F(�Q���#F(�Q�4Q�1Db���#�#F(�Q�1Db���#F(�b��mF1F(��E�h��DTh�-���*1Q(��cb�,QcF�Q1Dlb�����b�#��Tb�,b�,b�(���DTEc(��E�X������F(��6(ѣF�(�F�1�F�1�F��4hѣF��(�F4hѢ�4h��1�c�1�X�TTk�����b��E��Qb�ޕ�_�����;|[^�D�D?����<��?4��1�@z��C���@~|�R�6a�>?h�`I��{މ]p~#������I�������+���6&?τ��]�������
�)�c�/俁�c�/��������.���G����<�_�����?��RC �?��G���G�;���zT�����G���
��̏�5�D��������w#�~O�v
�柚L�a�?�//�盧�?cב������M�a�38S�����rE8P�xF<�