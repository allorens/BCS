BZh91AY&SY P��;�_�py����������  `��>L �=P
2+@ ���ӡ�����  �   �   W|hp�I�Q�ښ��
  /���UT>��{�^�t�t}�{7]�5��-N�X��P���E�|�pb H�gW��t�6�:��� S�4�
�d[�zz����iv4塻���m�����Ho>{½i��v�p�Z��v;0a�	ࠕ^����'M�t
�8z�:n�ooGq�yU���>��8�5f6�����37y=��e5�� � '�e�b>O������k�z4�&��=����p���|^�Zi�Ǽ������,M� l�q�'b���7:\WMe��T�;��A���n�ٍ�g��1�&��9;2��]    (
    (�J  �?I�Ԫ�M�0� FS�BR��� 4� d  ��IRTz�       4�(T�4bi�10F� F��"DU	��h�MS̩�='��4y���<P@�U(�S�`5z��� �!�M7�?	����?o�?i��F?@H�5��?�(�)� ��D?5��*��~��_���c�?̟�Cq`���I",��o�k��e�p��|� H�H�Y�ɨ�I$�I '�@*"���c����I�k�/���~�mV���<v���ݞ���f��x��k�C�U���"7^���l�9�CL��r��|�\���LO��4��;���?g����b�W���b4݈��kE���o���J���o,��}�`ۑny5�Y~���S��`�s�Z�jz�=�#s�_��QM�yWШW"x-���M������j���&�!4�֢�<�m:P(�=�������ꗭb1o��,��
uQM�4�Q�siȽJ���mN��F�Q�l.��o`W�5�a�Mm��?ח'C��mh��u�:V۷v�n�&�8)�w�j�ƶ���M���k^��X:@���ױq�1ab��]S)�q ����C|K#|[Y䲤�IR`�
���q�"2�p�lxcr4��y�5�[�v�x�g���Z<�����q�ʇ�Y#�;�5cYn*�y�6S��s����Ǌ-�b�n߭��	�x�x�c�&����?pm{��)�CtDb�\Ax�q�!W�[�mz#��M>7���Q�9�=����tt��8M�B�����V�`╷v��i�tc������t�F�(�-E2Yo�6zݶ���؛F4k�~�Ŏձ�	�y�3ݸ1َ�o͏uz����K~�8�Q�� �����ĵ��({��o[�����mS�� �X�z�wn.ޫ�hǈ׆��%���~�D|H9�vX{8{8{<{<{�6@��k�GzLDb�b	�:�q��<D�D�%��a�D8�a��8%�1Kl��<��-�T�K��&v��*{��o���N���4��S�'<�B�#�~���	
�t�@��%f'(XԈi�l�ι�T��TD��[%��4ύm�3"#��x=q�X:�E��Ǳ�ML��-�9�S2�b�t�y/�D[L�x�\:����M��1ۈ�0�+G =�x:hѾ*z/�?l��3���s��b�b�xخk_3�5c��^uM�8)�-�v�F��q�od���yt^��tqz��ȻF��C��k)�2t7dDMDn&��p��g�!�Y,���,m,g���`��[���lM����!�c�]��v���F:�cc����c��[)����ö⛟8M��cF8�X���ݸ��-���p�~lo[��L�t4�����=x����#X�z;��,�z���7M�i�i�M�m��k�u�`�e���;����1�5�5���q��<�n߭��!��bm	���m�7p�Ʊ�����1DF���D8�uN�,�h�-�y��D|c���aDE�����(�q��m��R\��pُ�^�1�����je(�	]T�D3�Y�8<?/'�r�������=�g��Ƒ�DU�/ZT�* �q���>G�O[mʄ7l^���#�>b�"
���8����N������ϭ�zxyW�s�I�Lq
o��_��֏V^�e�)d��m�F�6��ƙ-�E\AX�Q@��k~Ɉ����q��y�+m�1�Dy�8W�d8�1si�%i4��'Tm�zҠ�x�y�ө���$�+���'K;ْ�!��J�|,""�q�K���R&�S�E&�p�^�o��˚.x�?x��-� ��:�q��0q+e��lZ4�ޡcL��"� �q(Q�^!k|bB®��'�+�%}�x`�T����[�p-F9�0!6�
[�m�[/Rkb���x�KU.)Aq)������x�Z�{��U�h�+F�F�Q���S�Tߔ��E��b�/g�gC�Gt�R�Q{�O����op-.#Kq_
m�)�*��"�}=<<��爓�)�B����Q��V+T���}h�#^�Fד��r���'�E�@�U��M�$ZW)y[BV%�X%�Zߢ���yR����_
��3�V&,^}"�*����ϲ�D��/yx����5-46���i��L^X-�2�(�h�k�#b�"���%�Wt5U�9C܃�����y��{<u.KU.)Aq)����E�b<��E�T���T�v�b����qh��*�J"���y�^�{�y 3�P�h<����ڡ7G�V�xC�i��ț�=N!�'��F�8�Pԡ�}B��(."�Q�R�֎5e�,z�{[Y��k�a�B�V��׆ث�,%�<ܣȩO�>��%R��4%bX-Mh���UJ���J��	��*LG�6�LQcz*<���h��m�����X�V�m�Lw�xSsv��m:�����崮��M�%4ko�;����R����M�,P$!�yȆ���:��
��W�g�'�%{�ZB�&+𘲄�"�
�E+ԁj�R��W�1h��!�G�G±P��h����X-Q���_]��6�U(�(��]�^k8��~��ܨ���2��o�K���y�M����տ�����4F@���#0����ؿ-��%'G�7�V:ჂD�Y_e��Tm���g��P8��������v���ӄ���C���Nn"L]�؁�p�"B`N4�0m��JmX(zx��˽�r�Y�@���'�<9�oL��w�}�F{^�An���l��}���hD�_�ߋ}�ys%}	�n`<�z�k��s��{x�<�Xڰ~�U�>��R����rvZ�`��gP��"|���lT�x)��������uV��wPo>ӳQ���J�'�[�k�-�gg�~���m�{S�n3F���Y�g��S������ݽ���G>��J�׽�xNJxe�7&砵[���/7kx��ooe�{J9�exxo�ާV[ dDE妟c]�<t�r����q�H���n���i�h��}�7�lӓ4ڢ**�sT���f��6x�81wz6ꖸ�V����z�nq����ިN��o�H����&^�[5��%>���F"/�W�E��j9�?�1�Ĉ������C��O�۩�tZ�9U:Nv�]���$'�nj�i�V�t��z܇�/��S3�0���D|G�ox�ϝ����}��9�/�x���ov���a�F&��u���L�i�W���5���s��&��X,'�u$2���ڲVBb0M)b
'7�ǹxr:�+Q66Y����/i>��N�/ⶢ�ꉑbW5	�ő4^C9�����>�=_�±�f>��������Rc���n�A�o���;�޻��o���������&����'�5G7��5p��Wp�/%��5�S�6��뻼{����6ZUq�<^w���ۯ�y�y�\㈎k뭎���N7�� �?*��X��O��o��<11��y��ߚʯvx��N��s
ە�/�W� A��1f<�h{�Y��x6o��
i��<d�;\�O�6���r�.�2׉5X�분�E臒:i��{��k��~őq]��ꮿJ�M#*��)`;�;1�j���yv��@�����پ9=�f��g�\��R�8t,�.�w{mews1�Fa%�u��Q[���0�uq(Ж�Ҝ�e�;U�
�ըOoI� ǐw�Oѿ�]<��}*�"u������ʯ�����;�܊�
!��_����	�o�G��K�6ܹ<gs��K��|.~��g����u�%~�I����&��#=s"�$�"� ��< �����M�S�#�����:h0@����¡o ��	@BĊFt�V��Wo+jmT\8�Q�^Vd����Deٴ�q��Ŋ<�*��#�u6|J
�s�+8{��^%�'�Ǧ�K;5��"����\��p���d�߻J�baSǲ�(�3H@�_n�豬�`�t���t�f�]��i���s��/p�Jݸ1���5�E༲�1<&�ٗ�fO9�-��J��RL�Ǯqt�G-��F�w!�k���}z�@I}��{>w��腹B�u�~N�o]_y��o�|�#{5���I\��W��z��n��ʤ��Xt<��h8MÔKW��fjr���>+����8��-�O�n���C��$���!>˜Y�em���T�7]���K�������d}�R{���4(�גro�+�ﴪ���s!&5l<n�ǽ��H��q�_�<��_��.�o�YW��ٙOղ�L�x�mm���y��U���d��\��9f�L�}+Y��CHT=���_�̢m̚vm�f����Lb9:�l-�!�>�|�Z��de�!��{������/8��3K1�s�#�kv"~}k��)+�%�Gn�����5�R�p��1�tɆ�L�˙�wvֻ�M��OO[sG�n��}�o����ѳXrp��+6��ak^͗��{�u��XW��[�:�y�7lX�om�0�٘puV��Dh��q3nӵ��*<�[�Lc�M�����o礭�H���>��{�; <M*o������R���F����$l�ˎf�=�eZa������0OY���;��þt�{U)��Eu�v��lH�F�T@�$E�U؞��G ,COD3�ǞwH[���E .Z��ٌ���lF:ߣN����o=�,��%o��ZeQ.�7��$��F�O�B����ݻ��ǌ��eO\c	O3pd_;ٙ�Ӭ@���8o��3�܋u�����������d�
��9����ү�ֵO�6�י��h'�0�����e%�K*|��(m���۾o���΂sp�v�C�\���)��{h*�\j�\7�k�鹄�0AU���.1�쥢O�=�i����9��l�g��<і���h��koy��C}!��N׵r������m[C�`��
����`�v(I���$�.`�#�p�vc�}.���V�w�����b[]����φ��M�H�MH�a��$��O8�͍�Q���{�NV3�_�������EH�������tؐ����e�����$��?��>��&��_���mT_޽��2wv�+Iq.f��ܲ�e�1��}�3�x�::\R*XLq(kb��6���6�����Z���}S(�KR�-���K��gV�C2�lQ��JtK�˵�$c�� ��j�f=�y,�J�v�wz��{�n��,���YDj�E%Z>�S�fN���!p�Q���!����Q��m&���	$K�ێG?:e4D�Q���n3�� ���qB⎒b;�M�H ���銺�8�puڅ�y78Ŵ��c�;]�[�D���dj��x�D�x�F X,�䎖��;��{��7436uL�H[�V��~)�];��D�P28��J�A}�D��{lG ^�Ok�L]+b����[X{:|ߝ:>�O��鷵"�)��QT���B�)F�-�����_7G�-����eM���p�x7����EI�p�5G��J�Y����H�vvUԠ�O�IE�i�"[�R��}G�c���B���Y�>�SnД^P�f��VP��~w�hĲ�O��K27k\Ԉ�V��O�
�M�u��w�8�ʅTR&/Z�"�h�7�n난"�d�PAI[�����v>x�����&�Hk�I!��E��ThQ����	(��~$��|�A�\[yH;"&;!Z���ea4��)m�h��ػ�a5Y�A��[��\\������Y�V��]���7N��}o�a�->���/��͈T����o��a��
�k�H�s$>�3�m�/�/tY�:,�c/«VcrFjɒ�j�@A���������í��˳p�����\5~mQ��k���#4&I%����M�����?k_�t��zEk���I�Q��~��G@�?����?����9���I6�?������+�~S�_���� @� �   � ��6H@@  A�    R   P0��ݍ� �V����EBAP��J�s���;����`�� P�x , �  уa@ H@@  �  4�@��  
 � ݽ��h`� ӹ�
���5A$Q��s�f��  р�Ł  x ,@   l�@ H@   � `yh�  ������ @ դ���JI���K�K��̼��� �`    
 � H@@ !  �  X 
 � � �� l n�wt � YN���m}��}�z�� ��� 0@     
 �����  F �  X 
 �`  �    Y���wtF H?%��d��  H   `�  ��$� 0 �@
  � ��  `x  ��ww@ ]�I$���/�$�?��U$�����������'���qO�?���Ȫ�C�l�$!4+HR�*B�,B�b�/$�6lٶ��xa����m�m�m�o^����6��m+fͦͪ!�B�*B�b!j+V��B�����P�U�T�K�i�4�͛6m]�i�o=v۶�i�+f͛6��cli��m�Ok�U���IF�{h�Q���U&-Y�&6�maψ��ZB���I�7Z�5E�5���j'Cp�7q�L�כ5m*4�v�fx׏hY�{��5�b.�B�D���G�b ]5�����	�Z�+U32kR�;7��g�l�at���	��`��Ra��s.�~��|qn�^�Dhi8�2D���e֗y.Z9V���	�5���.��MM2�j77s�l����2k���b���c΄в�ABٝc_X3mj[u�Wq�{���V��A�䊉Y$f��M[�6�c6YD4Օ͹�,�t��"�{����|R[HDXF[t/�JY��g_�ɭ�*U�v�y,�2��آ���O�P��1Q`)�%��3�= G���%ݥ�D�f&�i��Y�R�h�|]`�ٲ�ji����p߷�[o��%�}��}��33�;��I|�I'����fg����^r��}u�\{�[�@/9y�{z�s��������^����9��zJڬd�a�8��3��2����~ލ���fm�j�)�a6�5������f�F���6�˭ZFӧ���#�5q��7��m}�V���촅��:O��k8<Zۃ#���Nf��跓��ceJ�%16��֜4b@���ӗi��Ǎ�Ɠi�&�p��tɣ�&@�Z]�6��6�@d�5r�{Ǌ�ROq�2NgrC�J

8B+�q��-�m\�t���o�t�$4z����G��T$��]H�Ç� ��=8q4��,u:��f��\�MU��Y�曭�uY��"�~��f��wp���H�<��Ix��4��7����S��ŗTK��GI�eN�a��UǍ1�w'w~d�e�K�]����p�0��Vh���'e��l�UIU�d�i30��ݔ��UR��7���駔���NSt��b�nI;��H��Ek��j����tS9n�=M���z�	�������6l��(��w`姍�J4C8����&n�w�Q@�L�Zm6�;i����Ѥ�qDp��(�oL;NS�9Yv��"v;q��Io��xjQzN��S�&�J
�����B�݁�r��qA�?���:�B��l��L�<�q�^7�j|8UO�[}�Vsgr�]'Ǯ�|Kf����d,�d��8�n������3(�J�oy�O3�ez�3�FE1$���8ۤ˄��A��T����UU*��&i��6�7
L�9Ī%4���b3���ǈW��t���;K,�0m$�ئ
q���-�UJ��jǦ�a�U���M��fJ�2��D����m86J�Q0�g=t�6P�Qd���[�3`{s9�7�Ț�Z𶨚8��t�t��=(�%ԥ���L���N���i%��-���ڧ�y�ZAÖ��OX��s90��U]>,��,D�;t�m�a���@�#�KK�m�kz.]ܲ�R��)x��܊
[ƅs�Hh��M$�J�
��s���p��UTL'�['��av��h�Sq���S�L0�Ex�M4�M�j�d� ͦ��/�����*�Ɲ��5m�B2�$��߳~Ǉ�$�*�..&R�������=8c!��b�$��7�\�;�}5��������8�:j��k�il(i<aąV�QEΝ1l��KT�������-RQ*�A)�KVX�J �� �ttӈ��:v��P<!�ș�"=����v���k���u&�?ODd5���݁*M�2c%��Xӵ�A������Z�~�Χ��Y�I'h��#,�bH��uf�/L�[��f!� �ו2ʕ�K�}�F&}�:*UIK2���=8p��\FGQ
���Yn>N�g}��dש�=��k-���L��:Ye�Y�*.�[y�0̽�'���pǝ��׷#<[U�뫺�3*��b�q\�+�i��&�Έ][<CZ�s@wf��%�'�9���V�w��8&��m3����i+�[ ���k?�]`B�B�^-]��V-^+�J��g��v�qeq��^+8�=^/k���q\|ǫ�⸽���\tʸ�Z�+�Uū�qq^�忙��Ҫ�����������|W�q�=W��x���^/J���p�-^1��W�\^/|���J95|�r�b����˗�lDF�Q�����y��П&.QhQ�Q�˙��x�;gNe�4�^;VqU~H�#�>�*�q�����>�:��c�3�O�U��_�����������ɯ��?"<XM��q����]Ǥ:�-B����8G<>���]�R��
��h�}G&�.�w�����.�V�Q�b�8�P���I��g�}˛�<�/t���f!M�K�
y��[��.�4l�H�#�������}\��Y��u]#�|�?n`�p��ks�wjpj���3�=���o5��߂)|��;��fs��7����꩙�{��JO�����g�i�~�}��U3<�{���9��;﮺�s/5R�8�Ejj��i��|�׵jիV��\�F�;�OUUQxJ
�*'� j�)�.Hr�$�*�VS!rm!����RD�
��j:���9����HB��b�XUIKl��X���B�1�1���}@RE4b��@͕����7�B`t��"]"p��Si���2����q�#QF,U'R��x��$�KC�>/q�f� ˦H�cȣS�4�Z4쭾i��i��m�ǵjիV�ԣ/�28�s3�L�����<��y ��R	��19T��-p���M,����s9px�a����4��b�:E8����s}��af�9>kqS1���%�a���&'��I
.(x_���4D|��C$l"T�RC+�=b��5IvU%R8c�45柈��-�.?4��v5��=��ZY4h�M��~+�ZQEQ�l���z+��[n���~�|8u^�s�r�Yfݴ��2��_r����1��|���YD�i�vʭ�͙��C��zU�95����|�B>sf� @�I���2HPq8Ƶt�r��.:���1S�eTK�D��& %g�+�R�r�U�6$b��/R8�k }��0�R��� Ƙ���/�Ř�+�r������m���u�~�2%q(^���$���5�����4G��LM�#ؗD��D���Bө�pD�7@t.���Rq��h٢�y�x$�?!|��G� ��<���hӲ8b|x�k	"� �,��e��0y�#�ˑ�G��J��;�\iU�K�q��i�m������j�^/o^U�V�Zw���#���DӾQ+� l��;eėM�J��	Q2�J��kG�jJ/ Ĩ:M�)�8h8`�Ds�
z��M�C"}rHI4��"e�O����Q�o�Cq�ݶ�u7�%�C�F_�>�Uj'�SJ����H'H�.��+�&X봙cga{3	��$��%�� ��Ŧ�▒>�>� e��&�L�C�l.�D[&X���+1Zc񏞴�M4�n��e���ڷ�7�V�$$)�4����b}�M$rޤ�˂9#DC14��R[H�@6����He#۬���I��7�QJF+O�O��&&�#�jW۹1e�ww'j�~zG�$Kbȥ�RT�J��Ӷ�L�)خ��%`���b@�@pMw7R��QzwΝ��<���+i�L?}��Ԣ�/���g��[��g��w�!@0�!�!Ã0�,%�G!�P���޴��b����֮)��_��Ex\�D�GNIeJ�H���l��nIj�J����x�b�Ii
�X>>d-�sZ�<I�1�\��i�]��P�+�4i*��T5�� ��c��n��zɦn�mYYv��_86~892�:K�u4t�4�i��ƚi����uw��N�4%���c3�%[p6�yo���i��P��蓕��%���J�������X�k�LV�JD�-e 7Y�OA}�� 1�3E��_bX�%�lU�V^i<M6�>��Ύ�3TUS)�������I�)��C�]VC�Ҍ����w��v��h�N�|J"tMFk:p����[��q�~w�ŗ����Q�����m�������c+�-�N��Q�o-�/6��.�*�E9N%����+L~1�i��g5rj�ed����	"'��y�Ii��Rq�̧�=!2&��Ww,����8K���l�p���{��������P	x�e�6���m��7�n��9��;�R&��v0V�������GTż[��SK׵{��x�.6��v�)��;�*&pZS��/i��d(4�i�Lq�1�;��m��de����\�mդ�x��7��A��)<O�4�(p��zqU%Q)��i�i.0]��Ѯ���K�Ss����,Z��ZU��2��,-v�6!s��yr$�Ng��>�<Z���mŵ�>q�a2��I� q0S��&bq�7юX&����߱�S敆��1��1EJ T7�%ѩX,Sk񷛁��ԛl���q�ǫ�:C���-����	�[YD�������c����pV�`p�a}	Xf�4�K��?3i�:d�e�&X��M�#���P��x�5���se��o�RBLd��1`E��=<���||���5$%��*U_ʫ���X�~U^.��U_��W�Y1�������Θ�_����/�������q\]/��x��Zg
����qg��yo̫����OW�q�_\g����l�_���~^�k�~Y����Z�,�j�j㌜^��WN3����rv�B��F�qɉ����-{_�k���>��j���mx�������x펜��i��*�j�^��OY�����.g�����Ne�i��/�
�x�c�qx�|���*>_��p��mOs��u8ܲИ��O�o���Y�n��p&���-�旒`vTaH�=gm)3P�R��:O����&\��8�F��3�%vŜ���`M����2GN�D��E�J##�Mĉ��Ƃ��S��$Ff҃�6B�KhF��k�ϩ�����8�͗#�zd<���!�R��2��b�/��a����J��mD!�Em��8��c����ܩkq!�_o���S��t^tb����y�������r��c$��o��Q���T�!0�P��q��3��JO%�xc�;7ۗ>Iid=��ě#���/�o�[�GW��B>�E��<7%���=~�f��w�i��y 6���ݱ3>j
E�h�_c�NH��L!P�� SH-k�������ԃ��7��5�v�Fۡf����E�}s������ŭB����17�hV��AR1��B4����̒�%�1�P�t�LJ���}�Y�:���M���Ki�T��m�U؝
"�#��e�5�	�����=|M���im���nSK�oԟӒ�{os߁US<�qɾ��wUT�.:wϻ���uS<��q��wT�]��.:r}���뻩��C��w{�.wDA�ir�&�MD&�J/�ɦ����[:�n���mQ�Xư����t���,:�`ᖔ0!�M���f�T���E�%�j>���u�Avn--]4K%h5""�X��a���,� A�w�W_���G<w�e3�l0���fS�3U@e+ˤ�e�/A���� U=M����2��
;wR���D8�0�yӹןGg']․��(�@=�M��:��\�8���9�%�Os��3*�׍�*e.�K
6B�4�����4�?~�i�G.L�d�u%z���,�[����.'q��'�`Y����>a�����!F(m���D� �Lg�u���%��2�%W"#"I�|��6��NU�P��sXwRF�\Rg���@�ĝ=¥Ė���9�A��]:�1V��
"S��'����,_Gf:V���f�x �p�Te�}.za$`��$��el�'m�&��)(��0d%䑖Νt ���iv�*�$٬L�N�L91䶏J����Y�'�,1`���u�L��k�2p8��踄�OYfB�@a�&&�9�/ t�m&)�/5�%:�!!4���m:!�8T��Z'�y�rh���G�ÝM�����aZi�ti��Ɯ����k��Z$鋼��i����0����R��y���i(����Ж!��w�ap��wM�m���5�^ft�i٦�M��җ��	F\�HH8	���I�;a�7M6�Ft��$у ep4PX��%���J�ÏX���)�&!@(�i������MLo�9z*��R�$M�c�������`�6������(�c^���Z�Ui8�]С�2��Dm�|�Ft�sl͚���*1'���P�>L -sT�����t�.��孶�ϗ���߱\��d,mLp�U$�0a�ړ��/!���SD�HUg&í�Ghd���V���i�������P=��I"��@�X���H�`#p	���Iyy�(�0٨�]���Կ�ak	\n֫�/�nBi�ܽ��z�D��N�X.0k�N'ݺ�����}ta�Ⱝ4�>4ګk3��,����&��4ᮝy�0dĐ�Y12�r�Q�*�a<�,��:�9tbHV0t�4ℏ��Sf�& ��qճ(妊��$�{������H�&��ن��)�	��/0|頴�jI&��
n�2��5ޝ!�di6C��;�u�	�1^��nH��ZBi�C b���l{P��5�a@��	�e񖴛2��k;�́����m�W��� i֛u�!$&�8��}4_\%�K2e��`h¥jT��-u�	"nmvH�L�E�IuD��ɒ̿�Г�#�:s�!˺.��|�xx����ړ so@�맚#��mEdLb���'�;�;z�+M1�mU�MM��+-\��N�;ܹ�I&L��2S�l����<y<vdF\���e�̱I��N���x�9�<��M��.�4�Q�C6�>�ܻh*l>s��f�У�G� Qp[���	��oq
&�JO��8!����d�ou�:��c��Ϧ0���´����Q��i�N��4g&[d�7q�c8���r�i�����FJ��[�	�u�Ju�C�4�e�"������x���;�:t�/΁JmB��3*�I�LO�;B����ԑBgߦ>�O�c[υf_�	�L�I~�	��8��/9��ߢ��s3����֣��w����n�Ή$5�2��JM�I��fM�cFS@d�V@�N&�g6�/O_��|S)IV�>H8x�����-
}5PZ��C`ù~i.Mu5~��V����cLWƝ��O��U�P9�M$M�i��ϓ.@������j��i����M��B9rn����x�T��	������i2Q�����u,��
�q))>}�<m<��^B����#�냑� 㮃��N����ٓ\r�4�Ljd��L������Z�U]�W3~Z�U^/��q�ⶽ/���\W�k��+��~Y����Wk��*�-_�t�*�j�N+��VߙV���Y=c����x��k��i\Wg�l�������V�����Z���������\y��}Q�����(���
��p�E���q�^�����[q�^>g�e�/��㦪��^j���xW
�x�4�goY������:WK�[��/
�x�x�1�qx�]8����?̯׺uBTק腢�,�qީv�;����I���,Ҙ��z� ���%{{;C>��hr�T��=�4��x���rw�Q���_��}L�Kĳw~?)���1�s�݌P�w���Dv�ǂ`��}��k��ߚ��E��yȦ�cn�j�d��ǳ���w��>��we��r��wwOe��r��wwOe��r��wwOe��r��/9�s�w�y���_�q�aX�8�Y��e�[�U]�vdf��-?5Ո�5�t���\�����2�8y�@6a��#�}2C�i7��@#kO��gwY�s����۠>��$��*ڔD��9M�L����I�fhQ[�梎u��M]�7����6�i�|N�|B�B͐���Bډ�S7|H�c �F(��-��������x*]�v�%�u�����x��"K�Ұ:ն6�n'$��D��3Y��b�x���@S��zbOW*U^�u�`g/��9u�р4zs�%�xe&�,h��e���
X���i�Od�p��ꊪ�:e�y!���)�R���aX�<Ui��N�un�5����{0U��f��5�≛F9���`xMn�#ic,��cj��T�r٬x�zq�ZY��S���c���6\6,�q&��}�l���Qگ�9K5h@�c��庺���r�0��=�I�i���H���1ڐ��V��.��Jt�o2UW,�Y����18�)��N2� }ìBC�HF^:`x�LO(�B��֤�dp��N��K���	��~L���&Su<&��V�ӵV�*�Ҥe$R�E�%h9!4�w�|D�`������T���o8��jq��h���`p�RyΠ�.@�Z`#��G�g J=�rMԪ��chjG�_>�l�m<]ͭbx6�7�BL�=Z��������>�׷��"jg7�k����)M�+
�,�!g�!�۝���͂u�97)���!����	�/Y��ƀ�r�e���+�����w..���_�>ЂO@��|�w��^������Q.X�-�!F� ��䓽;�{��NS�I{��#�N���'��};R���j��в˲�	��ܤq7�I�)Zpkin^=O����Z~+O�\m�-�M.����c�>�Mw�.[�w2=3�_@�s8�3�!%(�7��(�t/�L]T�����zq���U�ӗ� �ZS�UM���V�4V�O����ލ�Ƴ��'F�.T��+I1
i��UTl�d�lx�):���Lv�+�V�Uq��γ:�;S�%�?�w��չ��K�iz�r���өl�Cz�U�Ҟ��|��F�60�n�m�'���w*F3�,��6�j�G�P�B���@E�o�ŵ��P����&��Ck���jc>�iˑ�j�Y��KL�Bb8L?'�����[��i���x������W
*��4������5;?�S;'}���f\�q�� �eʳ�yڳ�Ŭ�y�_�Z�毩���b�t���W��:QQ/�D,�*�|ݵ��{�V%�6�|��'�U*K�J<� ˁ��qk�6!6�Ɓ��S��'˛ҩ1���&@�ix�eſ,�y|\X���}Z#oqSQG$�P����7��ϲbƷ�>�l�iH6:֭2"W�TT�Fb�1�k�GQ���aX��UY��֤1R�i���<�e7�k܏���&���Nd�(HoV��y�zٽ	������f�j�[[�����]��EZ�����<��dI}ͧ������WWtU�������1K��bI<D��� vx���k4�8�rh���-->#�����+
�l���6���g�(�r~(�Ws�bfs=�s�ZǂJe"��y�4��A�Ft���%��v�~�*�'��xm�8�� "e)�6e
&�[���U��R�B�Y�Kv�l|P��8py�TL�&@���-;!+���m1��VO� Q���ύ�&[m�,�	d�t���*�Z���Uڪ�Z�-Y��*��W��\ճ�g�����x�ǹx�W�8�^2m^��^�b��1���W���~S��j���#�hk�O��Ȩ�����z�*��8�^1�z��[�̶��%�Ū����+��ƻ_��q����?#��/3���#��:�f��<^=c������gn1���=q�[�x�8Η����V�/¸^�X��=^޳o�k�zg�ӌ�x�W5nb�+��x�\q�^/��T��˚o�[�S�i��ڹ�A5P�i�k��˴�@��U��eb�ԐA�-'�C��1N���"[�("_�����)(Tq'�uW�',cH�h`�n��G�:`�dpzk��\���N0��Al�4�f�Z����gК����������E3Q�����꾅���2n"�h:$uH�k�[�r�B4w!��q�uߢ/ݢo<c�ߏ�Ə�*Y��YA~[�Y��1r��Ȑ�;���P�X�M4�"�m'�9����W�R�\������w��Wb<)S�=[s�.n�Q��+�88BV��h��t{�ͼ�ݨɶwT�^-P���8�Sd�p��8��"�i�n�˹�sUqUO��j�UEJu���l����y�
�"aKkJ�-����0��AQ�Q�����t��I�I��:)�Y�\V���~�z�cy�5�f�@�aKb�2V>KW���\�ұ����0{{6l�Zv�,�h
��ܯ�ӻ7�;5"��N�N�$KB찚�Kn}�����g𬻺��������������������ꬻ�������ꬻ�������ꬻ��ܼ��N8�+æ�c��ˉ>�tV.�|(T/�Ivm�5��m�s|��I���i����h4�Ɗ�&�
%%�u�nw�_
KZ�0�]�V� }I�u ��]�ۏqت���#@��&���eIJg��oS��W���ʫ�� a�:��yɓt�>w H{�����hU$KsR� �|lj�k��6MJ��%Za2RP�x&\�L�`w��>�{'�u��^�cbWA�I�|3�S�sx��O�2�X���:�ic����F:V���lc~��Z��2���o�|Gi�d�Ki��[t��nc��j��]���ٲӯ^6��	�COqk[X�M	*����9ⅸ�ٙ��]��T��� �@lom���$���i=$%4ᔅ�KK'e��:��;�ޢ���<>:x�� �� ��E�p��h�j��Z>�}NS��6��ɃM��Wɾ�f>t��s���UJ��8�6S�zM�}��3'lJe����"8�V6�?>/��Dv�C��z�ޕTQ*�lt���1ɑ��IjYN4�6�jB�m2�@̕ӵ�#BV803zۖ���dÐ�F

(��F�QF�&�9���ç^׸qK-#m�O�x�y.��*���(����g�s>�d����!��;UJ�UZK`e�Ĥ:��׹�$�Q4l׋L|I!���i���H��)Ӧ�q��i8�Aa�I&�:L�t�_�>2�����Xcю;1����gS:�k5u��Y�+d�,�"��\�VN�=���Ѐ-��)��6R<��.�Lj�W�
Hd�`�RHN�� 8u�cU�+*b7ig�$,2t���]����YC�I�"e0��&8�M&M/)��u]�Ɨ�z4�|Uc!�oV�+$#�)�s)�UIzN%{��<�ڣ��$%��TV��6���h���4�BLƤ>̪R̹5r����߭ϙ?z����b�Uc�lcvGV=���S��n_	��d���ī��Ws:�^��!�Y���U�j��cA2��/M�˒�q��Ps[i<����tm�t�Ƀ������n�������'r}�����X�5����m�L��`<�2��0�!��c�U�ݱ�q��~y�5�}�� ��
6��I�/���]8��g�����W�ө��	�QDL1i&����]E�v��8<�����P�&�o�()���{p=�j�i8[���ߌ�<�$����uy�2�8�9����u,�X��G�<T��\�za��1���a<�����+�/%3*�c�f7>��bB[i���iFH�֊=jG�,>�i�#	T��,�VDq$������l7�R��?'O6��üϤ�7mé҃����o�rR|<M�9�2'�t�2�Rz<����؝w|v�b�Uc�0!�R	���I,~�b�\��b��Wq��/�n�
�<����;���*�F��fee:Y6J�FQnD��fS��;I���bc�/��g�І��uF��I8�'��#i�f?!i�0��]�S�8}�QU�.H@�<KN�����-�ې�e)2��$6��U��c��ĿwY�kź�F��$d���0"a�y�N�<O�Ҩ�\r(�8&p��/X�絜Ŭ���~cwB���5_l2<Q�W��~WlW��c���f���j�UN�ٖkXcOb4�卛(��ť<ҫ~�1�q��?HK_��qnR[׉�Ǔ��Ī�:q�\K��1�ȭdj
KY���[_�y����^ݙ�d���Xӆh���s��Z���*�auW�ۮ��3J����ͭWkWkV�2U��~Z�ʪ��b�Ux�/c��z^׊��8�\c��l�1����ÌU��⪸�x�x�U�~Z��ߕW�U��|�~W�t���q�/��Ŝ]�q����|_�q�W�WkW��Ū��+�ۧq�8�����q��gc�7+W�T;Q�!�X����G!G�(�ی��~_�g���[��:_˥~չ�O�U�^-^���/�����[ӌ�x�i���c����j�O�4y#�|��Q�4����}?;�����J=��Y.�E��H�σ�>����n�u����qC�*aWj�����VΙ��ſ.���uo���
v2����x�b|;xPj��Ǐ�y��a�c�?���ez��'��>���Nڪ˻���,}���U�w˹�X�����.�s|�>���˻���,}���U�w˹�����UYw|���ԧa�WX⫳��u������d��I����%���4�����H]`�I�3����"�6�6(�Qu~�b�'�h�hp���d�'��QU�[�ȝs��Èy�ްHI��$���#Mj0�&=Y�>x��UXګ����3*/b�b%D�5�$�JY���x���w�ڛ���>mŽ��$0w�U��]Z�N9%jT��S�[iJ�iجz��?ت���.���\&���z}#	h�<�t�q3��}׾�vu�����;iï��WR�]�'-Ŷ&\4�h�ֲI��ܜjG�n�c�������}T�vn��jahܮj"�i����T!g���7�t\K(s{U`-a,8`dcf��\Q�!���^e��0�O���I;�zp�B����MKbKZ-�(��HH�O//�
��UC���@���	Ep�2o��낂���%��C���]m)�i�)+��n	�lJL5��$�������^*J%ʸTeV�6u�1�m>rt���Z�Ͳ�fh�x�1\Uc�W��.}�}v� �䐄���jH;;B���:�we�_���Hso_�cR�>=,��A䲒��Ҫ�OSW-Ɋbd7����-��=��+nC/3(��c%Qp�oX�G^%�a��d������-+灇{�[�L�M���((�!
4B4{�݆�X�����l�>�I+�r�t�8�i=zy�B����s����D������ʘ婵.*�d#w�<~<�f�Rq4s��Ҥ�0�3A�B�6S��`s�B���]���:��:\�^|q��p�ltiJڻUc�Ǎ9�T�����cT�K����3=̲�
�	 � �Jg���P$m�[��Ejn'Q�[��s;�_#����3�$p��{&�����J�i~'p�Fu�Z%��p���^M:R�W��v�����<�	i17bަ���Ӣ�l���-v�AE~��HDq��v*c�!���62C:��c%��p��suְ/��4	��&Yt�"a�,�ko�&���F
_D�J,��KM�Ȇ��(�3�r;�lp�RC�Δ��ц��$$���ϟ����׼Gؓ��W��Vm���n��.Ϥ!a蔙t�_�i/�h����6A��)$�ˌ�M�R��я�d>�cO�N���|mJڿ*��U�w�o�O c�m0�F�+�j5
�HY����ҥ]�"a�%��1���%�O�[O$i/�I�G���ϫ����4�|ֹ�����T�V�*^oi��%'pbC'�a�A��x�U8�_rc�N�븺���-�	���L���Ԣ+�	Æ��ݼ�t�jߛN�P|jh�Q�%�.=���e�Np��y��т�,QK��������ٳ-&��^I�HH�ީ8�7���U��{��cGp7#'�0h�+�z��ʭ�q��P��#����h�:NJz����� 3���F����mw�ƅMbh�
r��m%F��8�!i��H[��NUUR�j���y� z�N��2����F%�QCi�3�KgJ�G�Ŗ��m���ަ���܄ۓ)��HO����$'J��U]-_UW��cl�8W��*�^3����^�K�v�_\d⸻8��긽�8�\q�x�\Z�[o<S��_��~Z�,���~i���z_�?+��8����m�6�W���m]��U�j�j�m�a�qt�<q�\W�e�|ϟe�+���nޟ5뼾3�r�=ge�m�^�gn3k�����/e�8Η���Lc�����*𾯭3���=q�.�e�8Η���L�U�_��W����6��_��~B�N	�~"��̶����i�s��KS���d��+jP>m	�-���st�]���~��s��Y�R�ЊBo)oNl����7��4F����Z\B�x��D���*N�j
�~Kj˗�V����&�j:�ۅF*S
8	R��YD����x��Q֞^94Ր��}j�g��T)#�z��~�հ����h�<�RЅ�7k$>c��q\;�+���I�	A�ʯ�dMQ�~6!�����ܞN�lp=l��p�l���_THzwbi��\Qv���M�J��F���ɏ�N��u;HK�3(M�a���`5�Zt&���ӭ܃�*r.H��(]�S�I�\��7{mqwls�,���`X:R���ڻ]�>rz�g<�R� Ҁ�-B�dyH*��E��	?�ZX*�OH1�e�먚��ƍ�s $�>CB�=n�[��C}�x��R��!�;,��}�� mtH�jXH���u��CH�c��vh���ꝭʪ�������ꪬ����[��˾]������]���}��33u����}��33uܻ���%ɤ�&�M|�/��2m���n���p�[ݕ95c[�)�D��1$vO����*F36d�ŗ\^޺�vX�1�8���u�a�蹭QE��ʨ᡺T��a'�KWMY��V����S�f*���{O;v˶�����/m��B��m�T�n��]`:�JI�̾��c:9l�\��=�%�p�=���Z>�o� �<i�O�B�:�l��m�!��B�1w�W��n�������G��U�U{9�5X�4�v%�\��GO$�巘��>�'L��A���i0=D�MY�ǱYG!��1uuA�ۦ�Қ=��>p�ߍb��q.�q5��^�>��5K�:ԭE\�x5�W�O?%���yk�m�Τk���a��9$��hc�5
��<�ˎ������U�V=U4{��j�� q�F�X�IokG}ڦ�Lrt�v,��M:k��֯kΗ3C�u�q�d�͒�'��i�}��$*�����^�:�F��R�=r4�d�j,W��N��ó�+�mU��_;A*�L]=����Q�ǚ��6�v�\�[�?,ˠ"���/��g}�B�W�}ͰfM�F��ڙ�	�	�g&�ӣ"$	��&�&�*���V������3��&Snh�B���>=��y,��QU1���%����B���^�"������i����M�h�t���\p�P��%"
��d��J��ܟ�L�ճ+��IH"Q�m6�M�?3k:��Y�w��!�<�T�F���B�Q+JD�,��zw��wv�5��''��e���[�pΪ���M%�.�$�U]&Mt���UR�&X����~���Q�qHm���u��IY�.�1��阮�^\Q>#��z��h�+��RI�$�ey���:�f�}�\>���+���1��˙��fX�D�,�4��UTT�n��6�T}�(��$t3��sw�;0��J��&�'j��'���O�0�M8��J_.�	���n��,���j2���}�Yַ�躬o:�s)8�N�_�4���K5r,O�x�p��t0�J�M��ǌ��Y�G/vwk8�J�xѰ"n�$��M�$7�Ht��h�z�J�X�OZH�E�zCPQ�F�4"c���A\�U��ԁWI$x�bv����:��w��6�h���R]\8Dن&_���:JO&��Dէ�<ΰ�Y��R�S�?1�m��Tr��T���&���Q���w]��Sx�]��Y�`��hZ� Ӏ8���W)��a���P÷xH�1*U2�.||��=��=����,n+��{;;dd���3�v�L|�|��|�1����\�Йk%�%��������H���d��b���"ǘz��������N�R��n�ͮԷ��t��!CdZ���Q2J|�	4ڋD���,����N;�\8(�6�#��0��I�O&�$,�(�M���:`d�S�*6U4��O]�̜N; ��~{�Ŭ� `�T���l:��Q���Ӿ�ާ����Y<��	�h<@�(�Ep��-��I.�����G�JN����6t�_.BB�!䎗������F�e��3����xQ��Zr�˕$���Tj$"C^�t����5Wwd�Vi=���C!'n�&�>$�2�|��Hd;i[0�����f�6��mҶ��mv����m+fʹ��6���ǧ��U�N:q�n8���o��;m��lٷE6m���n��hB�K��^^V�J�!
бo�|��޾m��N�v�m6�lٳf����Oz��o���M�[)�!!	�Z��*��~5W(��=Ɇ)��bY+١�
�z�Ҝ`rQ����߹���Ѹ�k@�fC�;������o=k�a��8����;�K;��� �m�ۤog'��=��ׂe��h�q\
�{��u�(ۚ`��Ȍ1�o��w'��I����������33}˹�����33}˹�����33}˹�����33}˹�����33}˜��⫊W�c�I>u���I�����0W��Y�IOZ�}�I��-�U����m��,���w�>Jp�H��w�F.�����F̹i������'S&�N�*�9���vw/gE��p�+��M}�x��X�wLw:���*�R�����5�s��L�#��g��t-"u����A��-$I8m�����ճ�1��2�	�*�X���0_((��(*���HM��Ǉ��`�/]�M�}5&%��l�<�Ns��S8��*��㮘m��a"u��ӏt�!!�
���i��tyB"n==$Q�<��qx��>�i���ۓ1QX�k�}�k���m�E�>M�\�mem�kp�n_bXU,�LMbؓZ��Og��;�gSd��Ś�z�(�:a�f�cϙ��wB�g:!��S\�UZh��-2�́������^Ou9x�9<��HHy�p��6�����7F/QJL�q�(W����@}�gi��T�*�lm�c�7��uֹ���͙��Xǅ�sRp�O'^j���ĉ�ԗ׎i0�"x�i��{��:�"\"}�e�X/��e�t��s����'S;JH�oi�uۣ�4�~����w�՚0��4��JҪ�1���ޘ�3G��ĒI$tg��I����}��$4���E�Ѥ�,�i>KO��qR���Η9��o5�ߨD�n��|���͚pY��N���Æ�UUUEy2�a�ʔѓ�����J���Wj����6��ϗ���w��+λ׊�Nqc�j����ӝK��ϗ�@�r(�1��&X�
?u��)j�|y�*w�O7�ˋuG�쫯����q>��>��1�Ff��j�$�#�|dɳ����p֓I��~J-�d��ͦ�&:Ro4B A�
A�z#�~��޲�W6���~]:��{ ��6�k��&>3� 甔��KF��6��2�J�k.c�Ȯcm5��Z)gC�Ī$e�e��R}�N��N�
a�t���(X� [�-���k�f�E�<�U۾i,�S�I�񉪅T�ݶB�}�������Ԅ�E��F�&��g��3�Ecʪ�=p�9�=�/����ʐcB������k�ڨ����2���c0�:+�
�U[c�
(������똾)�&�'�FGI��W9$�M'�c�3��q�e.���Qm*��ۓQ �K�����1��Ư/Y�'��>k�-2��-��y�y�[z�����kQ`�pn���d閒�s&t���'�eHC'��7�~���/��Q���T�UX¼T!⌔QF��eE՚�L�0386�����s�c�p�gqw<��x��2糋��Q�����s8���ڛc��;z�$�d��Hg)����0Ém�4�n�4���|U�/22N&r���4�N@�z�1U�Hm6��Ce2UW�m�1�\��c�3_$����q{�����=qq}EԶ�1��i���6`�I��tV� ��ve�$4�FI&�{T�MF����Z`�o�-Ҷ�>+�ip�x5��0��W���?F箺)��f<)���|i��q�c[�m�m����m�m�ٳfͻm�xxxq���qƹo�;q�O[m��;m�zٳU6ڶ�M��m�m���P�Z��J��,BՈZ��Z��X��]���m�ٳfͫ�m;m�筼i�M���gM�76�v������ͥ�e�%&�����Wz��ۦ
0�z渴�����ω�;�I}#���h�fDK��9j-��dh��܁�����S�8�&��	�M�;��8��gX�]�˵��JTQ�5lK�r�_1X[�3�d�o��ϴ�&��/h�5�XP�C���&�}n�3�%��L�!��~�n��7�h+�q!Q,9���}��s[Gp!䗶�w�r1I���N������5|ĒX7��74�X�S!��
��A��-����Ɉ��Z\�kv�f�	��(�@��F�˒˵,x#D�qH�e%�u�xN��׈/�߉$;�'��$��M���s���iec%��`o�1=�bXl�2*m	��N�g%=��ݪ{2?���i劔�,Ui�	��ث�p߮CmŅ�T�o]�_l!.��C)+��4��XL�$4���k�΋�q�-l�z���H��u�憷���x���kp�P�v��fM�Fظ�a4ŉ꫱&$K�xåL��ic����uO��m�����~_}��337ܻ��]��337ܻ��]��33=����.���]���wwL��g.���UWWU�8�1���}©�2],�i��(��ꗹ>m4�^��c�	e@3�N:<�f����'&���6�� K)/�=�!W�+��bB�~��g���3y�xg'�y����c��^����xK/&��tnZQ�;!��pq=�:��O�}��H��f{���Q�-NQ�r� �q�B311<S9�����z�)�Wla�*��c��v�3t�*�nRR^�N_O�0������ʯ�'��6jI&S�&�'8CuUƠԫ����.�>����q���-H��y���9�z�~�!1AU4h"Y^lö� H���c~UW�6�1���X�5D������	i�˒���.�fIR؜:��ێ��||�\�&�:X�pA\��Edpބ�����)��g=�cg^}� F�o��#���)�s�%Q%[��#���e�y<���G����*��1⪻c�0����TV+���`�8M�l|�Z�'���L��FE����1�!��"���-,��U�m�9��4���&�e�x�=�L&�x��.��	i��"��vj��Q�]%�d��RS;iu##�zv����Xc�Uv�lcw��\�ff�YF��|Ǳ���_Kuַfa�:�/���'��㊗��v�b)dg�Q��MU�c����.���:�qb����C��_����O^�	�A�ԁ�yHJ�7$`��[W6��e2�;��ɔô�wI��^�sp1����^/���&O`�d9i��� L�BUQ&v��4�+�<��VJ;%�ې!-M5M�^�V�ɧ�����%��4���0��Ut��c�fu��w��5f5т���e)�'1��4MHO>�������W����{�Q*����6q5� ��⫝̸�._�~�8��1��	2�%q1�ӗ�6�fM6���~�:>�l�w'#�g�L0ƕU�6�1��[l�-��o��)�s,��"S���p�~�C�uWsF�Ӄ�Ϩ�� �_�2#�ƿ�a�b�1��$��x�{�SIM&�<5|O:h�%���s!	$:��t��8a�<UW�c�{�|�Wz�k3�����ouJ����zl�C�܌�=������Y�����°�(�h�~�����|[G�$�`J�=0�O%���4)�S��<��y�<%8p���"��T`�l��C;U$�VH�OZQF�$t���Ae1Ҫ�c�1�\�;�53�ӫk]��L�J��;���\�S��5N�Moia����_]s�%u�|F��i7�>���w��UG$���-��~1���RHS��x~(���3Mn�UJ���|�o|�u]9��(�)��=t�|a<sx���7�S�#6��{M���:*BUUL�4e�h��Lw��i�Ca�U�c���^��������l�q0��7���S9Le-���,ƭ-�D�O!	*��)4��ۇ�י�:�L+��ꋬIX����p���mɾnT*����vr��I#r��H�CULd#��r��z�����w5��?+��I���8lٶշ��m]mv���q��+��8p�j�������q�\^>w��O\m�o]�Ҷ|�M��V�i��6�ͽc��|��^R�!Z!!j�j�b�*m�M���V͛6m���m�x��nզ���f��6ڶ�Ǉ����]o�F�����(������ۏ�bk�\Av}H]ٗoXQP� �+c����$F^m\,p�~�r��*��6�aYΝ������O��G�$y�]e;�`GU�~*OL�7I
x�I��=��$�۰��˻��fg��������33���t���陙��|�{�wuL��t>]=ϻ�������:8q�⪸��8���IEpÔ��J�TO4Ľ�{�����;դ,^}�=\u�Eop��m�-��)�M�%Td���Rx��:���쐴�x�!m�������<a�4�����־����F�`��Y�3{]6���_f�U�BϘ�7�.W+��ƈ�����BF���'SN��I�O:;y}oIN&�j��э&L�>4\t�L����I�����yz�)�]�G��)�a�*�� ��}'��6/�uu�F���׈��[�kV����	�r��0�� ������i-�'eO
�U �לl��gK��X$b雛nϮ���n��'�G3���Y���F�R��^2�7�ZL�?d�?��18h����#�a�Ii����K:�MF��4����=c�i�+Z̬Y1�"Q F8UP�/����ۣ��0�j��1�|�*nf�[G�oA�t�L�Zo	8Xb�����ok�����LO'k7�:����$��!�J'-��������7����u..-uw>��F\=��
b�K��]b���_��ȍb�>��ơ��_si;�zs�J��_:�0����z�1�ۖ���v$�����^�	�`�;4�8����F������Y����-��Z�k(�[E#c�C�C�������U�[�+7%Y0h��,ۄ��N5!8n�U&�	���2n�����O#!��1ڪ�c�c�}�WX�1�\������~>4y4�޺S�%�J$��,�J�[8�ۄ�~bd���a>O��l�߱�ۧ�4Y��	T�`j�ET���g#Y	-�>L��|&H�(G(�ơ��/�0����;c�{{�i��ܫI�
��fܠou��(�8�ݡm/_f3��mu��qjsz�h�6�2`8�˽1h��;���U�.K�J�'�8�����E9�}牄�If��$��K���a�䳧d�t�y)9��%9ϰ��6�$rH=+sJ�m{..>�;�%c��	�q��w8�����3�#x���cJ�퍱�u��z˚�+�d[m�[�'2fHG&����w/OoS���S��@T$�vƌb�E��q644��lO�}@]e}�q}�k����m���-a!����=q�l>�og0P|((c�Ut��>���B�~����Tn$�u_x�G.�鰣A��x�M:m:� �/\�s.�uwe_�5�)�����)C�#A J�4�:����IE��7U��Bn�'��=���L�T(���n�`�IĘ2;a�<UW�z�1��Z�uoZy$ц�r�s'I���@�w�+SQ��E�+���lb��#���0�r�Op1Uḛ���Pܓ��/�r������7ޛ�Ze��ު�*���p��ot�Ou[�WR��NuJi?W�����A��I?I$�I$��UTJ(������?�p��X����$!�  ��ҢQR	�g���5+��]�*�ʕG���d��#�
E��"�PR,�R,�H��%�A(�X�Ab��(RRY�QbRz�dB������,H�Ȋ*H��(�"��kԈ��"����(�,�QIX�E�Qd%�T��RXEBQRJ)%bʩpdQf`ȣ����E�-(�UQe����X��TT��,QlR1Z,��,��,�h���j��YE�YE�,��Qb�*FQQG��օ�,��,��Qc��|�Vy�UU�N�E�*�Z,QeQe,2�d��E�QE����E�,Q�FEQb��X��,Qh�E���YE�YEYE�,��)%�,Qd�eJ��,��Qb�YEEQb�(��(�E�X��QEQb�(�E�YE�,RJ�,��(��,Qe(��)%J,Qe(�E�,��Qb�QE�YE�,���YE�,����J,��,��Qb�(��)%EQb�(��(�E�X��IeYB�(��YE�Ie(�E�,��Qb�(��X�E(�E�X��,��IeQR�(��R�KI�1 ăH1�K*Y*%J(��,��J,��QE$���,��,Qb�X��IR�X��(��(�E�(�FE(�E�X��,Qe)(��(�E�,Qe*T�b� ă1�1`� ȩeD��b��,R�,��,R�Z%��E���R�*R�Z%�ZZYK�QKKD�YK��J�����X����K���$�J��))b�)d��U�,��R�(��R�)b�(�L�z�2)d��RR�,�Y)b�(����R�(���K�K%�*)d��Y(�R�,R�D�J)b�K�R�,��KK%*)T�K%,R�b�)%�R�*�)b�K����,��E�U,R�KK��)d��U:�0�R�,Q,��K%(���)d��U,Q,R�E�K%,R�)K�d��QK�R�,R�K�Q*�JT���)d��X���(���TR�,U��UU��H�j�UX�J���D�V*�,U*ʲUJ�b��b�TUU��UEX�J�VJ�T�b�U��T���*�Y*�Y*��TT�%X�d�d���U��b��%T�R%"�R*"�H����X%B�J�����)H�ED��)"R*D�X�H��� �Y	H�*H�*H�(��I�$)IH�)!H�
E�H�R,�y�������>�~\�hJE!�����i@X�Y	ERI$0>���'��}�5�'7�{�_��'��A���1����Ͽ�������~}��8g�Hb���'�?_��_������H�?���!�}���:�����)��R~���<~ ������>}��?����ڃ���$$����$�H�����,h�C�b~#����������?�!��1(R����������?�����B�h�Oȇ� ?���@�������Q�?儐2����|҇�0������V����w�"RRzo��i�k�k[�p?A?j~g�5���k��3# ���������@@?+)#�H�$�h`��A!�b(6AQD/f��!kL��]�U�x?��ӓ��<������x(�F �Z*�����T��EQ$�h�"DK����!��F�м������+�6~�?b;���ο�4,���_�j�?���
EUD����%���Zӯ������?��?����	���\A���_����~��D��&G�	�������U~O�?���?�������UD�C��$u������W�?i��zl��0��J�#��" �	�O�UD���'�����E]��l2�I����i %C��
U.V�T��W��Ԭ���g��	�,?�G�6	�rt���J!�����4	�89w�?����-�k�����#�	� ���ƪ���]�������
�����2��I�	���S��a�S��������'�6	��?;����'�
O�O��o��rDO�
?��������	�ª�'�R�G�)�c�_�C���l�d?y�v��������~��O��PC��'�<t?���H0�!�s�G �2C
,Z������KH���|/�� <�!��"Y��M~�����2
����Q?1���ф��O�?Q���(l�X�c�����'�s�����P9�!��s����������~�*
LS����; '���C��O� �A��	P}����G�ަ�O��������_�C����=�&�����H�

؀