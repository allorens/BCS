BZh91AY&SY����%_�@q���#� ?���bK>}@    �_@E+cB�[h�J��(�Jm�����6�J�R��%�h�f��[V��4l�kJ�Z5B*�6XҋX��[fƶ2�����scI[j���6�[3`Ҍ�Mj��mi�Ej����S����l�Y6ի[j��f��IbZL�Ԫ�,��i3l �)|�z�L�4�Q.sh��m�(�mu���Ѳֶ�pU��-imC�9��ѫJ�m��ZSkkX+[+e-��j1�j[+kLj�ef�R$�Y��kM���i��>�   �k�p u�9�;�4��9���ڂR�cM]��Kg@tֻZ+2�  uT��v��)nn�uF�ZKZ�r�ml֭m��m�ʥiV�   ^i�@n)�`@fr� � �X� ��˲� sr����8� �N�t �w
ݍu;� ��b�m�,�ƳQ�k`�o   ���  ]�  �c�� `������R��  j��: ڎ���,�� ^��^y��Co-ހ�ХA*���6�Y�23`��  ;��>  >�ds����� � �������j�3ǀ  ���z: �\p� ��w�� ��<p��'z�{@:k����U�P���6ef[(�SE�  cx  w����@S�C�\s� ��;�}� zù���z��{��� ��� 1��� {�� @Wz��5���K6���!P��   �  ��� ��
 ���  �4  �0 iws��  n����}�`�v�p (7F�dUm���Ѷ�3M<  � h �Ӏ �v�   �M�  Ew@ 'F����4�(X�`6�n( ګ  3U�Z��URl
D1cc�   ��h��6�� �Uf�7p ۳ $ws\U ��u��1`C�j0 s�b��[j�(R�6�ie���  ��� ���� `Ά��a@PN���w [� 4t����� ����F����2�mljK2�A��)�  �x@�V  �vn  n\p �h n\ �� �( m�� ��g(   ��$!CT��fU%TF�4 � �#COi��%Ph�d� ф	�&��S�!)TP �    E?	�)TP 4   h ) P I�4��L��LbI*z�����'�� 54р a���6n��:�S�x�-[�3\�5��;�4�[3+�g4�����Ab�2fT�u*���QYAO�*
����QEx�V�q������]�	B�檢���]U�r��+�?������ ����������C����d�"<J O�Cį�C�!��+�Wį�_��� >!��!�� x�<Jx�%��ġ��x�<J� ĩ�D�"x�<I'�Cĉ��"x�<J O��H��*x�|B%�Cā� � x�1� x�8�<H!|B ��S�	��D!��+�� x�<@�!��C�!�N%|H8�<J>!�ġ�ĩ��D�x�<H�$	�T�"x�<H� '�Sċ�b���|@� C�	�D�Ğ$LB$��C��P�x�<J&$O'�Sĉ�D�(x�<H�x��<@> O��� x���S�)�x�%<B�x��*��T1)�SĠ� >$@|H
x�� ��EC� ���x�Q�_� D|@��Q� ��AĢ���AĠ�AO�>!<H�x�A� ��S�CĊ& |J����")�ESĊ��T
�!<@B�x�A� ��T�"��O�> E<J"x�� &%� !��DO> <H!|J���+� �$Jx�<J�%|H!|H O��!�Wǌ!�%�_��� � x�<@!�Gġ�Cĩ���x�<B O'�S�D!�P�x�<B$d��~���������/A�R�Z��?�C�y�L����P�M5YCj�6Z�4Z���EYr����D�:  ����i��8pV�V7Lo�n�4��Oa�	@��;`�����B34��{h��˘�Y�t�-��Ć� �c.Rږ0ؖ�*���j�\W�(�+&RR��0u4�wEKU�o
�V��E���$䰥"超l%Q�l�U��|��s*��C ���J%`C���t�a;F�1�=���+mJ�	�:��� %T���zvCz�KI�N�e��r�h��R�įM���
@��(�{��q����eաB-OR��,��ڐZO^�{Sr�F6c�̓qx��iab���-��-�4#�.Y�X�/E����OV)�/� H!JĶ��[m����{V��o�Ϊ�`u+E��Z��Mʓn��6֨r�Բ�l
I8X�Y@�A_��w.�v�S�m�sڱ��� 	{"#*<�/4dPř�f#v݄v���%<���`�)��$cg�U���%B�Њ�qʆ�e���^�G�x@9��b��Ĭ�47*�1P��.��Q�4:�jJ���9��*�v���iY,X�V.	N����HF*�ڵ���/�4$�n��9qR{A
9���`���(�U "�EyX�U�D��k�p�+��/U�X11�v�2�`��ج�t����
�ٙ>o\��<�a=�#��E��`*00������48��!�4yC��ѱt�����pU��n��$T+r�MI6#M M,������r��� �Y��I��;��e��m.�0�vB~ה�:k1�W���7v*2� Cb�����K��m�-}�F/f� ��������.�ř��x
7��V1R��MuYXN�l4�֬es���*�OcW�� �3&;�tP�O6�jI��V�n�� "Ohm[&��9�a�)�Ք�Սݳ���{�-��ŋ^� ��NL�?��F2�w�[����s(əYWM�����Y���,�9���]Kx(i��V����5�'�\�u�J��6]+̛��#��Ivּu&u�m�4M�(��͹{m`բg�"/���.	JP�\ǰ���洴�vT5��̽j�����X�R�`T �4#�������U�Bh#Xܺ�B:�XmՠBu2�R�5�Z���A��\�كC�Y�nW3�U��*J�3��!�rc��Z���4%^em�ٓ[�l�� (��%��`���	���sw���t��a��dQ+�]%A��4��4t���ˡ"/C/v�bZ�!�����Ŷ*<��ݼy��n��f�"�/j;��W��n�1���֓��2�X�#��wE!�cN^�I/I�V�ߒF�R!Y3u�^�u��t��i�u����r^ye�De,��qJ��nh�v�Y���t��>-P�bR*��ٗx�*�o��P6PM�Ĩ���z��nbo	y ����ha�$�shn�Z�� ɲ��
T�'H���Z�L�(:�4���M�{wr �j�3��5�N�0O�eǭ<#]n�@7�*5�פ�Y��Szq*)��]���T�"���I�����!��D^)DML[�V"wktC��n+���i�vX�ܼ��� ��]�݄�+R�j����)�䲤�]ǭIg]Lxى��Ǧ��r�E+�c-�e,��"%O1�ק�iGB}a u��q�N�ǈ���L;Դ���F�m5�6�dLSv7j�[���  �8�p7�۔��j�H;��^� à����f�s)T&�Ÿ3a���ܡ������&ޫ�rh�egӭ��,(�Ŵ7ٮ�IY[��!O@6�cSQ#L+���X
O���V�����b�Oс�SN�ň���b˩X�mY�>SrP��ʱyZ�"�m(ލ��]^�̛/N�������Ѯ�Ҳ�'�l�c];�z��d<��Fm���5���f��Ȳ�$�6(۲��6�l1T`���cV�$�Z9��t7�0�ŐmHi��M	I�����0Sd����&��6�0Q��-R�+o1��D�T��ܰ�ɷq����9J��$���!{l�13��PZ���^ą����33kAB၊�rGHPw��h*�:��#5�O����e]M��w(Z�`U���+I%�����]MVa9��:�k�#J�v8��q��Blm�A@U0�[x�NI�-�䌇X� j�-�F�a[s4)t�f���q�x��-g��Ӎ��Xj3���t�*]�к2�r����<Տz�iޥ��ȓJ�8�)M�c�kiZ��FM��-D2�sH��e=`��U��
�oJ�`�7@q��P`%Y��:@�e1 �[H�-�%�\m��׬,ԯk*�����n�;3I)^bt�{$t���^�8-���Z��5��ZӐ�WS͕�i�CX�Ev��*�� �V�ܫK��(ĝ��P�tunj�v��핛*[�ęXV�C#պdaϴG�!4��XD���!^Q�X�97f�`�ݻ�B���n�躱l�q�md�G^H�m�a�GҷC)3��[E���"���
k�O�F�^��R̆�3+VݶkelZq,qTgvi4(w5����DT	-��[F�Kw���(�]�oq(���ˍߡù��e�ѹBl[[���-��a���Q@&^�7���#��+CR�Q�U[B<��XۙLn%�Β��3b���,)���a�Xn�)�if��De�/�w7,yb�k[��
�<(jν ����ӽʛڈ_G�CV<eh
�(	����C�NJk&j��b�ʬU0�"�"�EXN����S��5���.!Xq��N�oq��ґI²e���m��`�I`e���ī^ҿ��+u4c?5���le����lfF�Z!L# pf-B��o\�1H+!TOd�Y��ՇL�O�"��-�wE◗�楁)V�Vv��ƒ��(b�C]�Y۵��Y����.T���ȭ��
�3�S	� �X�2+(2s�G%;��K�m-8,fl��qk�{��{{XԓDC\��2�]9��d���@�mVi����]�d"�5����K��1˅V�ͫ�*�^�ǥP����H�Z�2f-��=�VLו��Z��f��)k���؅%�x�[��O	�NCr��6�Y�/BلE�CV��l��W�:KX���VvRE!�B%]��
y�-Sz�V�f,�����`�ٯ��M՚�*�O.���>쉶۬D䴯U^�0��s_����+Z=�IڲH�m�[wB��ÛtXʃ@���+��D�d�seꕏ��h�V���|0�M�kt�Y��N�[1F����l�5�G�v2�iL�oNn�b�5揮��6|6��q�u��"��%�̔�e,̷`٭o��@j����̱�n@�Q��R���v|�U4�k@�.-�Yl�,@Ҥ�![��b���Ǩ*��22yYn�4���m�.K@4���/6��`��ܚ�X6%/p�`�y��σ���ƒ̧��I���f�8�2�����:A	2�]�j�]��ƅ"�j��|8��	�U�-��DިpX��jhW�X.��Ljۂ��mV�	�M��6p�s1a��h�2<s0�Ze<T}F� �u���c��^���m�v�hd�;WE�R3�]��c@��M�)7��6�,smUՁ���9L�n�oKyj�@G���0^AM�4ҥ�i����ȩ��7k"n�i[�\ywg&��L*hgfY��f��,���mp.���u�P)�.���8�k�*�4�t�ͤ���a�����Yn�2o/p%�t)�����I�{/"m!t���^V<�6*�2�^[�G�u�
��X�9��Inc߉�d�:?:t�L�Gk3$��+��b��%Vݜ8e��:]	�r���swrf�	VP�b.��lR䚆�6��njg@EC���&m��9v�k�RT�� ޼ �j
J����/h���E�Wt,<jnc@�Z�cF�J	S~8�f�k��q������Qte��Id
�X��pԙ6��:"4�l�i��UnҒ�b'pn��b��a8�~�ÎU�߅����!��l���x���eˋ��=��c/z����&v�֋��w6n��j4%�O~B�[2��YT�l�ȷs]�u�iӵ��=U�b��I�v:Q����
MZ�}��V�2�K�<-`vl�ӭ8��h�!���#�Dm�*�fe;��eJ �B�f�tMz��uh�k)(����*�%�"�Q�s6f6������R6
��=ZX�D�X۠.��,�&���y[M��M�[`6�v?�ZS)є ܢI5�P�/�V�Gm�X����ֻM��Z�r2<w�)Рr�J3@\wXD�ַn���r��o��I����6&�j̩��kgZ˃4iǚ�f)z݊��A�@�h�Y�G�,�؞����rV[��X�4���{����c��t�Y��3��ٽ�Ȇ;ff�k�%amgآ�-�("D׍T(4B*Ӯ���.���s-ek̨��7
i�gK�� �o!;p��(���V�wE�wD[f$�Ֆ�����q��$���f�yKj�T�)�N�m*ʲ���/A1��%{���x�44�B *�ʴ7ms��$�ﰚE>{�;JV��0e��-�j�ݕr��S�J'&��r���1���	����ur,�ֈ�͕���Ֆ�a�b�8�O#JV%
Z��S��y�3D��t�Sb��z�5��A,�(��+ɳ��`l�a�Kn�6v�^��o�l��>��`_6 ��1���u2(
�
�`�"�`˂��Zf�9��.�3,2�]Ͱ�=N�%�����swjY����2^���PI}Ăxm+v�c����[�	Un7Cr
+owV��:tS�l7�)�Xh�ۻ�x��&�r��R��V+�n1���T�y�(vPJj�'R�N���pTcEҶiۇQ���O*��VfJ���I�k	YXES!n�I8�������z*�h���D^m9���j�쌎�]F.�Py���f��X�O+uk�qګ4M�z�hj5��y��fʈ�A�gi
�6�%��ad"��p��.2�6�d�F	��.@���t>�{I.��.�8N�b�ݼb<�w���E�Yb��r[�chꡈ8NhD\�&mѬ{M����&�-iQ�X{����y,�J�IsS�Q�n�����K7���0̔���)�dE<��<T�u{R̽�� Đ;:�t[�Zor��J��
zY7M�,�l�ݠ��y�T 0�(��۬:�e#R)Y�����܆X��EfO���5�ocgI2��S�-����`ei�oN�Z�x��۔�6���^8�4:����z����G������hJ_�b�e^�2Q�Ț-���(V���\��b�Tpf�{gc��<&*z�����<�+ ����(Y�N�2��/^���c�����eVC72D"���.��$�!�F�un�d��l�y���h�ӻ|E�̀l�y�r\�`���P�S�sZ,m�@#Yl��%�PCQݽ�9�ݰ� ��=XѾKr����j�[�j���%D���g7&<�F���ҘkN��FP"��U��jS�7h"�D�5m�ҦK�Z��l�	[b.ﶍ]j�u�.�gÐF��4���Z�E��V�A�:1
E��2&�ܷ��P�3�ڴ�&���1�+t`Zdu)m̢�6 	Ʉ�6����	���y��*�Δ#�A 4a������v� n����$g3t���z�4\Y�8j���<I}�P�^6Bz��g'p��;��*��]��YT��� ���0���TcC�h���A�U�ncQ�[+[v�l����L`ӇQLܨ�)4���/Z�d]<H�l�
b�n�o)��i͢�p�ķ�#fLʵ�5�()��l���5��Z�Mޭ� h*�rb�[�˭g,VeO�ڴ�Y�&�8jM���m��,�ܲ��o[�#!�$�r�Yz2m'Y�����n5y[nݢE*w����eZ�B`�zK�_by���;�(�j5+JW>Pһ��Z�A�r[��b��懌
��i��L�MC����`A�1����)k@<f�� �V��?��`�����@,�(��Yél�FF�Vj�鿯O�2��� �[�/k%fR�TOba��	f�aG�fL�^��/�K�uw��v�T�w�oi�� ]�����ٰ��.Q"8�'p�d�&����]����� ����U3.�,B� �����Qs �b�0ɢ��	T�z�¯�BȪ	���8�����h�y�L�twr+�@=+E��xY��i�`�m��Y�}Wti6��yGS�Fk�I�v
5jIz�`P�r,���ot�{*n-�(�("f�@$׹%B�*�e�0�h-�Z�R�v��n�!|d�M���kv�kb�Xӳc�0\���ǣAј]<�u�<��l����U�D��37m�M��+\���4��eL	awN�ۊBBB��w�Vj�d��F��c���AL��Nh�Ӕ���̴0Z��Å(5�&S߷w�ʩŭ��J�{���1V̎�a�ea�D�'l3��`���ܽ�$Z}wZ.4w`�U�n6Vn��m�,̫����!�4�*Ԟ֑bD�G���2��Zڳ�&�� &�3�N����]Ҳ�7�V����[���}�h� �؄=Zq՛���^5r!��6B��&S��4n]hh��$qn꼟52�܁�ZY"B�;�U�V��׀9����2 ��(�

[.�Ɲ��H#4�b������ɭ�|b
�n�J��@<���7����[���j)��e�1�Cc�U�u�j9�Il=2vV:�{pXJ�<��n��n�9ݓl'�>P���gsj�!
�59�@���l0f˟;Ğ��K�}�"�eJ �7���׽�Z>�7���A{8�0�A�]��e��9�u�|
@KʗՃ��n]��9�H���V��+������M�$���TRx������M֌��y��\�ʛN��]��4���s�ͻ�Q��I휵z�s���\��6�et[؞ݮ�v
�My���S�m��[��R�}Oy�7.�SCt��A�(u�M�'�d.n��r~���[��s]���ԝ�.��P�l�r��bvV��4{��瓁���Ə����t=�,�` ��G����R��|��3X�ۇ\�ɉq�V�Zo��a��ٍ�U#D=� ���*�N��7O�2��;�wGX,��3�|�>μ� Ր��N^˔��g<���GL䜳�Uc��|�PK0/��O_.Ty7_U]A��Rt[;��b9Sa�㧹:�W16-#eܽ�F�P&f��x5hh��W��S�K	�O3R*g]f�jX+����u1����B�b(e�@�)N� +��Q�+�m�(uh�; ]��5=�N$N���}��1\��fq�X]>�9�r�ql,�g�.�q�Nr!\���c����6v�{�9����TFQ&nnZ<�$��ڴD�L���u��s"@췑 �9~�:u���C�-�~��4]'	�|�NZ�,��!s{�7�4��RZw�H:N	%u�u�=Q�KX�{8P2�,Dbf
�z7]�l��X��[s�h��2p�+1�CH���g�o�S��+ұk��� r��*s�h⋯��x�l���][mykt�P7W��跌j�z�	o��C����RK���5���[C��j��ނ�\�+땖��;Nf�߰S=Vsx��.,#�&6�*V�]��a�uxWT�N�8vN��c��ʒ�{	�0e�6똆�f��j�w�J�[ܷ"+Yw]j���(�H'�jp�'�`����\���Y\�؅�-���͚�d�Ⱥ��e�ܼ�|#�"xn�͖�/�yˬf
<\��ek��d:�>�X��\������Sa��ݳY:*��V��j�Ԉ�;��b��Y��HN�|��փ���\��w�M��Tj�Ƈ �so9؇o�zi^��8�ݓk0��1��=��o��$,؎���s�Ԡц�ot)�z�Z�Fv��j�+���dSXS���Dh��qq�sp���%<�b��K	T�����h�g݊��A�(/U��_ޮ��ZzB����]0b���8���^�#���ԙg�Gj����j8GȊ&�^��y��VGk�p���ڵ&kn��t��{��ݵ"��e>��Y�/���`Y\��bf&3L�]�֍��IF����gP�T�}��CO\FK<��QI��YNJc6N��S�Lǝ�L���o��j��fgs��&<�1�n��ݷ��*Tє8<5��	u|��Ԭ��kS˓�F1A5|:��s�{4�3ke�e.�j��y*92īT���Y�V�:5��ù)�n�����{o����\Y�[��MF���^nË��� �Z�9cN`���_#\L�7/K37�YNB�B�V+Rk�3e9��o{�Nu��p0�[Ш�9E��̕a.k�)ؤH�J���m�(Vյ�_W�!f���!3��E�ks�\=�e��%��S]�΀�/�2��M�7J�Zè�ؑk�x���ŵ�o���7��w#K�b��N5���)�:�4f&87f���3k8Ekb�z�r��`�8���qޠ�� ��+GC�[;�!��.{��6hI��о8���rZΊg�|�_-=�=/���ͺ&�ܱ�]�{����2�s ��>�q�P�����ױc�4���[���_CR�۸��R�h|�'��R`V����:+o�	���Qeu(\;-�5���6nV�p��̣�m���nV��=�o���ݫf�m���l<�͕�Q����M����::��\�im䠱M�g6�=ɒ��+q9q���,B5��ք�Bv�A���]̦r���%�l��uG3�n���<2ż���p�9ZW8��&r��O�ٟǕ�//��o���E��y	�IH+�)�H躳�-tQRu�05��ԫ�L��ʹ��拨�� `����y����
�Y�-]K��N��t7��������X ���[�'Q�l��WM����&v|'�q�
��*�@q�Nn�c�v�p����L��m�HôX���J�����9ѽ�`po
�.����_]uҮD$ܫk�k�m��೤�v���@`���V8T�|�J�ڄS�"c�]*����1m��y�G�Vh����F�	��]��8�oR�^��&<���xLμ�9b��I8�Y��r���}W�2��*U�d�oD�8΅J��r�Z��&�QN������a+��`;��L�3AU2�-��d��4��A�w�R[jc�s)u�PA-�{��YvD�KQ�;VT� ��X���fu��kRe�&�gX��S�J$Q��.� ��k�Ͱ��Tb%��~0��J�J���Q؟)���rR��|��Щ�Ib	vj@��ڡ��R��S��g��we;R{�%�A������4=tv巹��F�돣��]�g`��K��Y|c�kΐ_S��ǔ�Tlo'P��.�1���:�;�/L]�,R!�v���r���b�p�*��U�U���Zm�Bξ�Gt�������Z"��*���jQ��n���ݮ�;5�zf��x�D%���f-��l⬘��9�4�뇕��"y��e� &�t�
�����F�}z���85�h�����\��/�{n�r��8����mUʻ���ڂwP��h���Cܚe.�25ài�*�ـ�ov��L���7��"q�:�}��"[�v��X���('s��n��h����N�
��� t��#ǳ��y�����Aov���]�Mq*�c�I����n��-l�X�0V�a�:9���"�'�������D}���3z�S�J]Ch-�z!��NԹe����^�F�ș-'����x�����!�Ws�}\���
ЕE�9KN��2\z݉���^��e֑ړ�J�&KΙ�0k.�+�Qę� 7���#_Re�m޹��3�����Z|طo,1�:te��AB(f�@^ \�3�S���*v7Ǒ�mي�|�;Қ�K��{n�qQS�[3TkBLx`ՙ���;y���N*v�a�C�u^�+��x��Ut@�H��:�}&ٛ�.�I�T| ���M��s:]G�����`�vr2��O��tg|p�.\۶,�\C7��]Z9��K��X��V6�X�"5��+J�>B;A������l����`|9��x���#�(�M�f�eY15��]/&����z�=ł�QT��:歐=
i��i�x��$��@�� �_T=���i¸�"��:��<�U��;���9;pD��ڔ�t(Z��%+�.�5��	2Oq�8���M١3�-L�����b2n@"߱饉��ʯ�v;��9B�R��Ut���ՀC�s=~�U�&������)S�u�n�']x�$�:>�����M#[�5����/����l��p��r�U.�ʉ�{8�p#V� c� 2�Mc�(A��wm��!�%�ڕq��k�ʵ_RV�q�-a���V�${�2����f�[�'�Pk��@P���ۮǷ�d�H�����@sn���x�4F���|3ԏA��1�o1$���ٕ����k�m���k�v�	9�U���
��󫫎;�4���X��z׮��y�o&�ľb�.t4_N��N�ޭw@M�n��Y�č$��.�Z�YW�gs����c%�9��l]�K���11���(����kU&����V�W�$�m�k'#}q
��u�6�z�'8����j}E^�3x�u���1�9�����p�����sp��ei��ɔ)_�!�Q`�]���_��F�"�['m�r��ukB	�U0�ɔk�M9f�̾bR�p�Kq�^���6�$A�M����΄',aݮ�p��e8�� l����G�k��2g.�v�C�ު���).x�G���qE�i�/�u�d��fS�!���L�*��M�]*�����َ�
�6��fK8����B���	��&X�f�⯶�\�RҌ��V<f蛍��Kx�f^	�J0�wf��]ؕ,u��`B�ԛ�;p#˘@�3\���s''v����T\by0���8�E���2�G;m�����S�ή;��e�)'��E��bdp���u�Vc짹4�����Տ�j�������U�O��Y�#{��0�
;U�s`:;+fe��T�O@�d�"���z�����A�F�.8W�y�3��J����3{d}M�2kCk yN�9�-��\�-���6�ͥ�/{������-/�զ��:��M�+P��VvX�+cu�R�H�c���������s�2
�zT�We��]@rS�m�!8Z������^�u�w_)�*����bS�K���8�P�q<l�M�Z� K15r���[���ݺ��HMr�U�]:{��"���wȧ�C��o�X�et`���I���5T[z+E�0�WN�}�D\2�i��C��$������o���}xYd�,��hV4�/jҷ5V�9m���N�љF;Q����-��������x��M��:�ټ�[�gf�2������fw-�Vڠ��aQ���7ک��=*�J��{/w5:f��Yqr+thߛuɉ.泗N+<8���j.2�X��=@V����;�*J�/F�wc]Q	�%��V^�$����:����)��"6���X^�\K�[uݕcFC���t#{�=Tx!),�Ջ;�s�ʋ1t��1�BSW��-��٦�vVSA�J���W��e����B���ZEE-=���䰘�Y�����w�4����=V��p�:�n�V,Ԧ�9ys���;�oJ�1̲�r�m�2��#V�Y�e��$&^m���fpո�ES7D�$��\�Z���+�І�C����i���G��!��Wv*����K'S4FT����Y�c:E�H/�~s7����gOU�[v�^�cC��n��g^2h�#!D�=�d�r��Ⱥ��a�:��#�@�Q��.��^�,4e<aUsT���"��Z�ٴwL[��Qə��b�9Vm�u����D��m�0է7PmV�u{��X�+V~m�d��z��Fn^\`�4)u��)*�����b���vv����.��'C��m�X5de��S�K�D �N�W9��&�s�A��35SsU������.B�J>��3�N#vFc{�Ioօ��{B����칵43��1Uӏ��)7o-@B\��/�켚x��<䒞��)!,��ԑ��<,��`�疝2�^F���kjY뙜���{MpyBN�V�ު�\�sz�5lumK���X��WH���-I]&k�ۀ1�`�y��<��tKS��!\o�gtTkL4@kE`��+4�r��
^Z&�T�wuB��+5���%'C4x�h:y�r�A*t[�۰~�e��=5S���ol�|sV�N��f�S�&��)��`�)QJGuqnR�0\�0�2X�Eå�D:o�����l!��70�[ջ��E��hd+�S@=�k���
���(WG[��K�3"�]��W�E)��X��E'.)�T}��F=�6u�bc�fk2�ʎ���x�;Yn���0A!��
�ص`R�vp!��[ܜ\Y.��8mGP0U�RX0M�a��w'�5�M��k�Yn���n*:ˤ�7 i���8�S*��.�C��IL���Q��K����A��ef5��������r�#�eu8m�݅�o@v�|�G��+L(�5�g��ɹ��	�\��f�^wd8_ˤ�}��	��rڲk�]�{��e�)
�Xd�O�h��ڍ]f��fmPj����v_rр�j�'֒�~������u\��f��7w��w����i����l#�]��0͞4�q@6�αЅ��7�m�w�dV�3���bX�k@�����=Rin�c-	D0��p�b���M�D�[����X 3���l�5��̱�h�<�����)[��u:��'�;/r��j�ʻg�- ��OW.�^��ZYX�.M���c�AlR��Y���(����VZ�zLT�
[`wܥ����(`���vM�܉㲥���+-VI�fb��cR�h+!]�ñ[�����U�ģ�z`���� \�h�oD�#&r����è0\�ͣG.��kkeGaV�;ֶv�>����s�>�L���:�����x��.WW:�Qrd)Aq�`	rN��<�-�M����r��x�\�����nQ�.�7Xr�ɤ�P��ڒ�9�X��ݜ�J̔\�g�F'�VC�L�҅��7�U��s�<�N.Dxv=q1��A���!צR��j�=2�(i�oa�V#�X��U0�%B+J/�T�|���;_GR_oTĉ�
<V�\�m�}�'�YAR��WC��ۏ���:���r��p�VIS`s'� >�`�˯_�EQxsC���~��z5��3�F�c�8��UDk�8�"�W�X_<!��xh�dz+�(¢>�I��t�Y?A��m��8���0Wf��(JN,ܪ��[�}B�r;d�|�U*���bڣ��~d������ӛ_��{t~�>��HV����W>��PP� }��b��+�3��j��h�+DMWդ�����:_�:=w���x?�?/��Q��4A ��םո�4��������|9�ݼ�*vWklfu���)+�t��RrYצ�Ө���e���L�73��wV.�R��А��u9��J�л�n�x� Ƃ�NSN�׻-�\��w>�E12ҩr����%��5�]&�R�|�g4'6�1��Z��(��������΃��7������m��ʀ��˺�h��� 5�Ҏ��kj�4��ǽRս�g0R��%k%��]=����'W`�j���n��P�{��Q�Up`��f5�S�	K�%��󰚅��r�;%���|����.�#�)�.ӎk��5h@q�j�]Bը,�jp*��٬�9'������T�ԥ�����ܮ�h��%`��v]���U�6�`��.��£���+�//x��BB{m�w���8e���O93O�"��w�88ؼn�FZ����t��{{�,NcM��������/vAC:�Z��X�|���Ӫ���U�:Ќ�3uK�n��`���LF���|q�F�aC�aX�>뽄q�X �L�|c�w#�*�j��Ɩ<��ߠ�&���غ�sm����>ڇ^N���7��vآ� ��*T�tWq�����[4��Eu��O�`�P�}΍�{]�����k-���״�NB�������ZY���9�L�S���`0ǶӦNm=(���\��S�\�u$��63�p�$�c��|s�KyQP#��^+�2��+z��tjR�J�:���p�Ç<8p�Ç8p�Ä8A8p�Ç8pᣇ%J�*T���VU���f���Jn�
)6��c�-s%�ff�{/�Jݖ�;{S�R�Z*��r��ǐV�9Ʒu���'b�cNT�a��d���l�U�h*��Wc? �c|����1�����锺���8���A*Kqީ}+�Y�V�\凕�R���[��D��uۮ����y�s��O�Ӎb�9��k3bl��������x��C��}7���#��������͍6L��ܥ�즂ۺ7�;:9�~O{�B	u��V����Wtu���SZE����C4�j������sO\k��^%�<2���2K��R�V�w-Q��=�~\�J,�a2��[:gH���R�Ċ�#+7�2�f��cl˔u���zh�ቾX��RQC�ݔ��}H�f��}j�Z���6�,�/d�쉈�k��Y�3��c��{VC�*�n�(M���O�S��+�5g4�@�2��1�Z��9�ʻZ��M�СϦ�S�m,��sJD`/]X����d�Ĉ	{�W�b`h�5��p#P����K��l9C.VrÑ�0gi�6�f��H��qt�Gmv�A쬨6��Ԗ��Ң\�P?h�%�6�!/:r�(�:.���Qd�as��y;�u.�u�u}ɧ7�w2�1f�$����-�Z��V�(EZ�Z��ՙ��Yڸ��W��*��y��)�8p��8p�8p�Ç8H�Ç �8p�#�8p�Ç8p�Ç����8EO��Z$e��5}.IS�+`T*�`������{R�*<�-�E]���+���<�����p�	�_#4�m>����D����� ���QWbkG��i��H-U���,2�V�8E3ˎ�%l���sBs6h2����Mi�z�����j;۳m[�y��゜�[���k����QU�k��<��:c����l���ئ���J���mh�}�����d��*��R�	�6���T��{��n��:y�M�8`/r��u}As��ě�k���k=�';Uk�6�����8ڙ���Z��-"��cd�܉2�,��uenȓ;�����!�]�����:�N��D�'n���G�����e]���b �"T����V���̈�b���ph|��^ ���ba ��]G��Ӂ<�Vߡ���)>6*��s��,tz�%u֐��{Z�\�8Y����c1f�z7�qA��ֱl^RS5#��R�kX��ֱ�\���>鼮%oj��'x�j�^$j�B��K�,��p��pa��($k�:YOkM��>�E4��e_}:$^ϰ9� ��ފ�w����O�G22�:�k��|��j� ,�ZW\�a�MR��%�.ħ�<J�\\O��yVQ�N	���-]�ʁ�(�(B��B�X+�Ѩ��F���˄�C�t�Q�N�J���#�8pჇ8p�Ç8p�C�p��8p�Ç8p�#��R�J�*VWc��}��v
,ޙ|���	,�#�v��C��&r)��f�%�0W׎`C�I��k��]{�3��>b:Y�l�q�P���UN�{8�K���ur��+!(�Wuw�T��f��2���c$8�⥄�-;hإHb;��n�����iW#+� ��9ط�:ݘ��4s�-���KX�Żc�]�fﻗ�v" :��^�LrYv&�"��j��7��5wq[Mgj�ލ������n�6c�~��bwf����gU��v
��:A�Q[��� ڷ�b��.������Z�i<������BfHm+���X�4���Z����j__�$���3y)ARp��&�*�L!�r���)�ӳ�'Ϭ,�b�7}�����ωG]m�&�1ɥ�����˺��ءxƚh�t��3Av���ҳ�p�`��4��`N�Uՙ���ĀW:��쫩.�UL��h�fs?��( �@@(7�u�h�}�:�L�5�0r�@�n_n��55⥬�4)�
����I�`�O���%]>L�l23{iv�r�l�vZ��~d��P�o#�Q-P]�,:���"�����T�n-q�C~+�����߹�cN��.L";��}�	D����(I��B�:3C)�gwr�r�_Ws�3%Eq����=ޔ�l�S�JWJ���o���hew�h�ԊE����oX��L��BD�0p�À�Ç8p�À�Ç8`�Ä�8p�"D��%J�*S�WR�J�*T�R�J�ܩI9�	{�9]h���"�@��:�����Lr�K���L��f��疲���f^ʀ�������EZ���o]�.��ʺ0�xF�u�(D��12˧���	�X�w�!M��8��Y{O����gtN���`;%`д؉aF���R�A�����)n^7Ӷ����+�1w2oI�"�B�O��jح���I����v&P'Y�� �-�Z-�����&nNn�X�a��9��5��+e�L#a�]���oE)�Cp�٭��tn�f��v��v��μ�*��V�.MV�C����Y	�P�M5 ���M�W�.Un ��řf�H�*A��f6�P�P��=������:Bq�Q�;;�3}r�x��īŇ��ݢ5�|�4-ɦ��y]ؐ����]0����d�9�B�hFnk�	��ʝ�x-ۉ_H�ֶ�1�# �Φ���u�Ⱥ�֓��4�>�:�d��xV,�Ή(h��wǴ)B�U���`�����E��O �����3e<:Eo�����ⲮJ�p���*R��h���ժ���ʠ��ۂ�0�1��/����� (�,$9��yL\��mp��I:����}�����"��֖}�!��Jm��N\�t�^�w����:��b�������	�i��)^2Ő襘Ht�6�v��5�r���]��ɗ�I��K)�O`=m���_)��MMVF�6l.,���z��7R���V��s��rLOe��J1c8����:��fDV�Ӻ��AɕۙS*,�4O��d�m����05+�V�j�P�C�6��9m�y��Iݱ�k�.�٫��4���B����yqH<�I�H�� �fc���ʓ�D�
�`����l;��O!Ck��ڭɵ�����@�KV�fY�ϭ7Z9ʎ��6S�+19��#��2����86�[�]%�keѡ�t'�8˫C(^���K_^�8��6�s!�k<�W�(�v�t+�9!Տ�Z�|�M��S�ċ��ʾ�ʺ�[��<�<�
���	yis��qfR�՟�*�QJ�t�����"��(r��Qf��`�S��`��q�F�	�԰䲺-�p�}����U���L��+�%ӏg����������g�e��*b}����7�0�)*�;x��7G�44Z�G���+�7a]�|9P�7hk��'���vSt�[�)�Sj�s�zZ��Ru�aX�D꼄d�VxMZc73l����fO�t<wn�?�̊c��]�V��-��}Z]����U];;e�[v�m�(5Ope�)NV�ޥM�p0D<�u�.�S�غwm�^޷�q���fZ�n;�)�q�E����Fv
��x�G3�W�����\���j�*��ݨ����U����q����[�̭�\,'�����RP�DYL���m��9���'DdE1p^`i����c
��L��4��+�hZ>��DjX0�v�0�r����l�Xm/�2�	��9��t`J$<�u����*M6J�_+G�k\�,
 (�O�B��J��6y��I*HҠvP7X4Z��4�x����feԣoj��:�F,��'c� 6��-���΍t�e��1�
��3NH뎺���y!�
H\Ƶ+�|��{._'Z����R�٪���5����Z���SFTx��y�&��P1��j}8m�%�|)l�Ν8������eCq�X�69�b�&M�X{����
��1�-��,ׅ���or;{ϘήVNm�L��j��bu�0�d+3~y�PM�8%���e-9d wWC�'�@��ET5�.�6b�X�w��W%S�}R���y�mٺ.'�ٽ|y���)��I-�C�Db%m÷�V�W�otİ��ce�m<"��}0$�gf��&���+捴޺{�F`���:�ʰ/cH�i#8|��������GAe�@�|�(�e�uk�a�
�̶�1݃e��\�*m�HT��P�}Z�ZM���΀�X֘1��Re��2�k�mC��)�@�o�W�b.m�����$�x�VBZU(ݑ@�Ok;r���A��v(�ʰwz������#O�䛙���X���Lg/c��ۮ3�Z�D)�j�պ��4V�u(C��ϧouT�B�>�|��F��0{��G8���� ���hj���cqg@O{�I��&��z�
Ô�nS�+gF��"@Mm�O#��d�!�4�}a��ms���
M��VeѶ`�'��O� A�Ʈ�NE���c��f�Ҕg�oK�6��Sn�9�T@���� i�B��0�9e�dt���F�M5LsQ���' �R�O8ʑ�Ox��	�_nN��ل=*t��Floh�j,�i�r��/�L@\��bmsn�X�(�A �G�ʛ.h�ɗPW)O����u���rnV̺��ɚs�b.���7���+�n��1b�� �o��a��6�%B��#��<d�/�EǱ+vqM�_f�c��*4���E}�qX� �2��v(!Y-S�fuGY ���uiT��t�׏{L�n��:�%�Q�S����_P��� r7��)یV��I�*_=P)�����
�<����T�P��̀q�ۢ&+:�Ӿ}��{�T���@�'�!�h��&g&�c~�uښ�v��l>��k�8�MZ6�h��Ư쿆�LJjj�wa�u:���� 9���Ώۖ�Z��PB��*v�sf�ѽ�s�6��!I��'`S����m-;ӂ���bG2������V��&�R��+��Ț[�`/20�7�覘*|I&�U�`� p�����Q���1�R���>�D�)��C��V�h��r'@�7J�tcx;,٫륐*ɯ�RQ�G�8AY�/L�f�s��	����W/����䇻�^Yy�VĀ������\���Lz&�2���%�C�f���m�(�� m��Q�촩-}�xN2s53�(��x��*���Ɩ���u��ʸ�a�5b�f,4r�YqiZ��S�����-9���S<���*�׵eb SzCo	f�mk�O�`�ՊTJ�ffZ
�K�N붃�EA�."��GQ*^�%o��w��j�W^���X��v�B�������u��1��*����<��K.�{�b�bVә2��wO���|&����2�nw�u)�z��WB�����h����P^���`����A��+A��ЌUč�1��F�Ss;/�B�捄�Vw2�k��޾�v��,��tg�8��]8b�`��)��n�U8��m1EJ��fB��fF*���k��6�v��HLZs*\�k��uӎɝJk�a�ZJ�(�Z`v��\m�3H�E��U�b��\�X��/�B�Ύc�>�l:�!9ven���=�LWZv��F(��D`��� N��b7���--=(cǟr�B�g޸���sz�S��|N�й�6��tr��Tvrܲ�%%7v��%�=Q�]�<�ʝr����4�50�>'����ʫ<қ��>˱�E���hQ}��=Ƃ� }{(-&j���K~}��*�	�m�VnZ�Vο�Z%-�U �PX)v*\�7>���D��,r���w�4-u��1Y���w/�7،<En���-�v�X|T����A����6`��ZM�����p����)���0(���l=���J�u�R�t�;��A�v��7sjrް+C��=���i]]�<]�M�3R�a3.��.�����Td�R���y�7��U��j��b�u��S��`�k��9�c����~�bg+�3�ɲ8�M�˽���x��Fp���l໏gd�%�.e^ΙR��;���ݶ�p�l��ͽ�Hr�Q�
�J٫�aG`T�%�<bgr���hO�**Bb�z�l��a�m���v�dG�t{ɼ�����Zk�z:��:6�8@���/6�����MZ�"�ݗPV|�Ɲ��kӉ�*�7����ɟ�V���$'���ZK\�L��OpL���)�j���Zi�jMq%]N���eʶ�7X�����<�$:r��J|��6��b��,7b<5�y�]1�r�c5Rt5�-�+j�h��ڮVB�(^aK�D��Sg�Y|e��lU��P��B�R�@t~���,=����%*ۭ�}d(���c�L��Pm�����܄�u���)��X�q+N%J��Y5��T��V�gJ��z��(� �������]��`	>PF�2��������m7��?�}7��L��v�̔�GNMr�z���g+���j-�A#���Ed;6����nn�|��tN�5��qS�Ŋk�om�	xC�V^��U�7��������֋��䕊�[w\m����~\U��Gŉ���l�fP�ń4����'
eְ9�����jش@^�N�P��7yJ��Ǉ��k:��n�Q���^=j=�햘ٲ͞�0�|:v*�ʉ�TX��f�SG+�����R�@ ��wQۨY|k�x����"���']˞B��U�n����3���upN7v7��v�f͢��S�Z^_;��g'�Y˂��u��X�r�n+���ׅ����7�zJ�o_T+�Ot�xpP7��Y�R��Z�����SW��^ˡƃ�0b��˝�z�@l�Xf�]f�A��3vj�ztK7�ʫ�O*JnP��0�4�LQt į@ʽd^d��-�ۈMc�De�r�M1>���z���C�$�ݘ)Z�"�`k�;�x9�N\��7��h5�#��.t��P̸�����NF^�oV�K*�H�!e'[4�i��S֞>����� TNK{|N]K����a��L��w'\��z@d����it��#*� �ȷ5T���Wv�>x�*w9m�n��su֚�عW)��aι�q���j�"׼kv���hݞ;�޽y�I"��j��$E*A�CTV��X��h7F�j���j��N�D7I�HR�[ l���v�"���6v0���X��$Һ��-�eP��oE�n}�����x�ظ�GGr{��Ƿy�����8��h���
&��Nؚ��؍>�v4E�[jj����
��[kA���|||hڨ#X���AQD[t��k귱F�k�Sm��L��������&tEA��PU�G�MGF"1�kL[h������4�q�����[+��'N��tDݍ4�t�CM1Q�P�*b��i��|||||�ET���U_^�����f�0AAEE[
�ţ�(�k�=4��1؊��]�^ڢ��&wn�;b�5QQk�{��V")�n�Wn�k�h��*"(��:=۶�TA&رb1���c5�h���q�у׻f�+mQQ{��h��mP���k`�V���f�(�������%�0QD��z7cG��$�1U$E�F�?!L����~�u*�#����z^t�J�	���
���ե���n�
{YK���oT}��#'B��!�C�07�`�[�굹��q�n�jZ:��ئ��5N��y�}U��\��M]*ʴ�`���O�CU���"��en
6&��U��{��"t����Y�]=��3o��9���>��}�.����wV.�
9��_�M��v��'ǽ[8e�H(�g���.US�k�'N�e.י�������b�����*��f�
��p�{ۥ$8��{���d�:���P������?[�ZD�eJ���3*���g��ifΛ�φ I�)���п{�0�@�Fa�_�W����3TϧQ��� }��Ց\ܕ$ ry6�Rxi�&67<jO8$�eו���.��{r[�}P��l�{������~�;�J��@w�����{����
j�A���}��)�a��伽F�{�*�4~�J��L�}~�N?.��ӿ<��iŜ��(�^A�^.����u;��R�vR������3�$���|}�޺[{�ј�.���Z�F�re��:��}}�{/k|7�V�F>����w�:��nSZ�ӕ��h�����|���k���9xnwMOr�l׉�,,�P5cr�(�I��G[���O]���Iov�,�Ҁ�:ʇ$����y�΃Ǝ�W,�
Nvy����?=���:�ze]7�F��T�_��j���Xh����F��p=�^}s��f}lf�1j��eN ����L��O�\g��lo�8���<�X~�ޯz���ي�)���^���y(u`�f�!���V���wL�EV����e{�Y������6��'X�-͐B�Of%�1�=��̥bjU���}ڗ��|���gr��=����Ξ�=�X��U��^��;�3c�[�7��s��bW�u@V�^�HB�R��>����y.���W��П<�SLrr�0J�����҂���'�u���ף!=v��J����̡�J?U�T��"?�K�>��:�� ��À�^�'/پX'T���������{k��^�y���W��C����h{k#D�o���<��gS����y�F}�t�����&��[|�����ю���yW�om6Z&��(��s6�,�7��n�J��
*_j��������}W�V�E��/ ��B���ٻ�8��C�i�~��[�5�{��:��q��6���&�vUF�IK�L#p�������x�,=�b*O��{@޽BH�F�9]������ڝ7)����U����5�T��_jR�6���Oo���	<�n���Ѷ��:��'l3ޯTᾡYhVb�,�=�|^���v�z�w���}iZ�&n��5��6�Z܅\k9
�F��d�	�	7v��� ͫ��k��QM��)?v�WK�z�DWo�n���鏫��|)z���57˟��zF:[��-����|�u�o�enL����5o�_�N�ҽ2����u�R���NW��^�
���%��.���ԧ�*1w��46rLJJ�b&=��q-��$U��֣[���n����1̔���1�R��O8D�.�[�%n�n�������(K�T2{�L����l�����>�[�{z�{�J�+�����y�gk�`R�\]�0��;��W�w�ϗB=�C�c}��o���V��U1ꪎ�~�U���{�H��)�:�����y��}oK];�о�fQU��?<z��V��s�lU[6޼3nn�V�]/o���>w��~= DN�	e���� p�6/���ix�M���ҷ��A�8j�%Iv,J7H	���v��,ۅJ�oo��z��h�gc��P�9_��;8�=�g[�.�b��6ۏ�JNTQ�����y���� �h��j�^n�ID��T�M��~ӽ=;3��􆠕��{ӽ���M�jc�Ճ>U�:(@4���B�=���]����ЯV�Ғ���\��V� �>}��˹{�Q{��ž��G�YF���U��?^�N�$�$4Ҥ��g��U���u�-�eS���`�Ľ�����]�W�fT1g�x*�}��7��]���Hõۜ�o��[Y����^�o*��W��	M����T<f�^5�{�w)���oL{���z�j�l��^x]�_H���l���Wd+�̍6iz����T��9|/]��ukw��/+��wK�I��n7����+t�Y�Z�*[=�ʇ{�X){n�XK��J��X���j͜5`����+��*Av������w�r�o�+sf�ˬY�w�GI����o��Wq �5Ue��P�\؞Ot�r�Q+�A�Z=����[t4R�9��@��d��(v~˦�H@��L;������o�f�F���AF��u|�Y-#��m9Y;�$��R�M[���%�QA�܌t%.�}�Ow:�zU����iW^��
�����t�N��2�͕�IO��]xu.���/I�X
��K��e��q9S�>��nm���5S�)��[Ћ���C}���u�1:���iU�q>��{�'w�=]}Ջ;i�/{W��u/wh��APK��&�KM�mAʂ��������r��~Ul����gk��[]	ɺu/_yV����z(nOׄCH߶]��޿m�A1�Rr�hPΠn4 3�+��;B7���@J��ԮWe�ݾ�Y�
}1䡔5��ޢ�>���U����78^���X�+�$�vڋ]��׫5{�ɖ�2E�9pס�*[VD��dv�sy�{X�3�<-t��0��gv�=q�~@GX�c�T#���<�}�+�{̳*����������K~���=����0ה�f�*��:�Rb����*}�Č�|u�Ր�K������"�M�"��~�w��fQT�����7�S�z������&��)TGK��:�%n�3Om�KQ��j���6'd�y-�v/Y9� �2]a*ޗL�v���*޾@�IԭԻ2v�ZƏ9XC�.3i�	��V��ڞ�ל�/�mӴ�|W���6�
��k��3��N�=�O=G����뽫�����9g�7)u�zW�.���Ƒ�*�{������Ӟs4gM���:٤jU�^�@z�{���#M����m(��9:yN��+�����S�F>ۻ~�4���j亵�:��W���r���J��V$��n�B�����I�kW�|6>�\T+c�V"��W]2�{f�)zo/:=���?M��׋3�<�9�HjU�~w�V�R3�c�0��:���=%�{�i�9=�����3'QU�����j���j�ٳU٫��Q<�9=�I��Xh�F����C"�Fʧ�.�z�^�M�C=:�_�'��ŀ`�vv��z�1ʳ���TJ�C;K�{��D��W��^�F,
:>8��U9��6�s4%B�2��v��D�MC��B���[΅�qԦK�z�N�r�-[cF�`=@_���P;ڥ��W�d�y�GQ��QG�R�
.':�[ع��+��ww:����b�C7�@��oBxђ��>�S�vԧ��dM1�NX���eE����Υ�:-^m��t&nU��މ��9R1;�U]�{��G���"�|S�k��Ǫ))V���F�����_!�]g���{{hq�K>�+�-��.U��BϠdUi�[�D�j���*���z�ә��t�j�T����Ͻ��{�`���٨��p�6�'g�#/p��X�H���!���m|֟E��y�������y��t��&����V@/�t��U�>��5P��}[�3���_s�ޞ����Wz����!zU���)~Ϟ]�>�'�M�
�� ���'k��}x����/�]��Nl珇�W��,�})�s�/G������sڮnݦϧS�$5�9\^��o�1�k��o��n�yT}{}�k���n����t����M�C�z������V>bй�
�J�
�W�x��+1����|����5k���W��^�+�g��d��NH���1s���f�V�s}l����B�$����������}jkn�:ޜ�t^�\ᴺ�f�L�S3�����l0v�5��ջ���t7Un9.�NN�е�]�����+�[��N��2�l��2������]��[����H��]���Vϰg��g�����+���T��0�f�璦@;�O;&����;4!%b�+��Jo�
k_�*�{�z �A�������;G�:�u��?Tw�6�t��[gĿ�����Nj�s�V�)%yZ3��9ME�����Y�>�\truu��t;�K���}L���M�ǵ�t5��������R��=1W�qgG�������]��=�������JӎT�!	�[��߸��	+EH�zw���;D����U��{��_�(�ӥ�𞬯JC���oz'v�]��R���̄3�}�ݒ畾��SL���f*��ʞ�T���S2�C�w����zޙ�Z�=~�ۦwb��Y��|ǲ����n�U��xV:=[��/k�Qq�D�&{e�~W}�����T)*�[8ձrЦ���5NR�g
݆Kff�R��kޣ�3�W�}YV�Y�C�o��#�!��Z�RꬺW�O�K����`3Ӡ@��2��MO�kg��2���GGu�w[-��ӖV6��;;_���܎�s��d��^]�z
rAm���9���Ն���7�wP�蟂0ۑ�=?	���n�W}�?�/%�?N����͠��s��������;)��r�'�N��Ts�p�E}�W���ϨQ���S}e/m���^y�U����#��NFޣ��V�%No��������I5�����M�{~�J�\�Y�rZ�� ٕ��/p��o`A����=0B
�DXǯ���ݭ5:t�[˪�M���*t�_TSi��d��z� }\��}
���j�F�(�%N{9zM�7:� ��9 �Ǉ`�_l��|����b����-!�{�33��F�OVN�{�� ���V�*���﮶=���[骧��?(3���8�D���f��s��^�nyW�����"��3�w���`/7�_V7��B�����b�J�J�Y����+�M^�\b�zc�����1�X������]� N��/'�|�)a{�4a�����nf�ؼ�)�}���5M�A���3d����r#:���|�<n�����;f�Ƒ3���W�)s
�uU�N �`�����Ý�mt�$U��i� U$��s�*���h��!�np�ջ.߸������{��%���Rߦ��ܖ���kЏz��J�}F���8�[��Koѿ'Ѡ�}"�\��u[>>��j޺hzf]R�{ۧ��Z1ɌΕ�6���V��9X����6����y�G���HP<~�G��GFni�:�(n��ʆveZ�}�qk���l����y���ˡ�V��B����6�b���*ܜ7o���U/]�o.4-n���[�^��$}�Q��1*`�j)U��O]*sn��OQ+��9�߇�Ɯ~[��&�6�ᆕ5�9�zY�=9W�;��o�[N�Nh�����ujO�}�G,�sW�[^�N]Q��鍾�C��m�X���K
�,.�T�y�Gh,�9���>�/�?o5p��}��nP�����1b�<3��(}���^�@c��"�q^u��^ g16�8�s3(ǡ�Ǥ#��Ѷ%�2qx�j.+f�¥����eFWk�θ&1��j#Y3V75=srA֟S�V�S���^ҡ�!|;h;�ï�À��e���Swn�^�7����`L�&�cr���㫂sޣr�%�J}j�K���͜hN;e���CCwun�I���kF�����yE�m����"��z)��[��� �x�؛5����)˧=e��G��Iw���݉v��ݫcn��E�Qs��S��>;�(՝�,�[ܘ�m]8
"��	��V�&����[9�1��`������)M�vn�Օv�H�m
]q����m`h�x�sם�=�BTE�r��ՙ�m�ׇ;/��H5��MAY}0�B\�$��$�5ZB�-��G]�X�T7]���w�C�b���:,a�Snk\�j��Wyo�ȯv��N-�Uɋ��]%��2�^�:�k=0��wS�)��cx�q�K�k��u�����[}E9*�Ԛ�B���Y��T���S��{����w/nL�`�2Ӯ\�^�i�ʱ>�T2��^g$�vvԥ��3X4]Yg+�d�e.]�Fy��Ͳ:2s�.K9> %����7�����K�<��+^ Nr�Z��^��v��%Z䬔ä��0lF
�kN���D�Qn�F�J08s�H�K�o��]�o*8�%O�p�^9r�5�J�׏'�ٴ�Wˎ^]:hڙ��j;�ܯ�QW�Ξ�h4/F�ě�A�r�[�
�;�ʝ�3�U
�����Zzm��-�$�Ov,��������Z�]ս3C��rRӂ�;7h��-�ǧv>֫b.�Z�:*��z�:�[#���4u��@��M�R�����j�Y=h�34� ���#�%
u��^�K,+f�]���,Ii���
�zNeC�q�5{��@hMY�%!��xV.M�Λ(���kK�"�e+�m��{���`�� ve��k;�r��)���3aqގ]��� Vl��\0�nо�c{��+3�ī�0�r�˛�{��+b��EAu�P��0Aw9
��i�f�u��u|v�|��|:��W�.�eu��d��Mp�5���t��9���Pbb�	�!����"r�y�X���ܬ|���,�\}X�P7â!�5�a�t��T6�W �fI�`���Ʒd͗�Q٨ ���E�V�k��謳b��J�y��[p�K:����f�д���jA��E���/U�$f���lL�Z�M��w@�N'�~�ي��\�̖��$3Ls���≼8�S3s�ʽ���z�]�1ɲʬt%8�/�0Yi�nY�q>�E�]���cv��ibnQ����݅�,�u&јw-�3."
qJ�2 _�kk�rO�:X:���[�Ci^�Yu��u���Yw�$��V�n�(�/1l��k��*�^����s�7����(����URTA~�i�΢h��b�*��o�`�(튊���1��?���o�

_�cc�)"�����f>������Gs��b��8���>>�����*��1�"����$���TU����^��=qƢ��&؃���������4~Z
�ֽ����mb ��"���ո�v(��F�q������b�>>>8���ON"=m�MX�݇��� ���^-�����֯mv5V��O��Z���I����b�mh�˩�u�u3�:�k[��Wm�lZ�m���{��ň�ܚ��w��m�׮�[U��j��X�b4o�=��/�*�S�͎�˩�E[a�s��>���g����1�w��6ϱ��;�4i����5cE�lj���t�kwnkE�D�v���j1�G�Ʈ��m�N��hgb��ZߛQ��;ݽ�����#�m�E�1��h�����7��^�-Q�Z$���5�m����������QE�U�4ii4��[.lM��<q�5LA��Q^�}u�b��]�kn;�&4!�۸tG`����7M�8��\a�	r�@�:���5+����
�.�֩���~�=wA 0}ݗ䫄���x��)�+{o�����ؐ�s�1@!�ʴ�G:¬])Jj��#��<�?J�#m�u� ����zTW�r=F�m�u���+�_z��R�r� ��՚}C�o�b���J?���s��Ʌ�Y`�*&-.*}>��U�¸���>n�5���;��{:#�$�^�P�F�-�!|=�L�����@�px�8
F�����g��`7�k��K�L>�E�:���3utp���q��/�]^���a�2���,2=�xM@~���l��A�� �c���s����jٖ4��5m��ϩ�q�d�x�,q�,՜&h)���1�p����vԿjW���^��9�(�Δ����[$x*�e1��	����|/���\����x�H߹����c�g��<�2ڨ�NФ!oԪ :��(.�n�|�m�������t���|�v>����x����@���A�_�	q�[\#�v�E����1'~�8�7�x��s��F��/ۼԖ�p'zA�}}|�F	(q����οU�`�}�FW�tv����L��%)�.�D���K*��4a�k�Tէ��8(1aϟj#�<*�]^�3��t�����&��8����]R���mf��)���ȫQ�mͳ����Y�.q�3i����z��7^��"��5%b�ڢ��fw1%fK�UWK��'����k�\�>$u|�����0�/�k�1�+�|\��:�Ӟ���ɉ�w��������;��7���i7kF�R��*f��:)WQ�?:Di���5x�k�{��}W�8�|���R�wB���u|/s�S}�����F0#=�v?p��^=��+��$�s7�v��+��m�������sj,xx���G��$txЭ���r����@�����ء5+������G����X�V�XJ�>QA)�"4r�W(dl{0�<�g�Y�M��6�? D��OA��8~���xl��9�W[Ҹ�p-�^��Q�Ӵ��ùؗ�D�E�}��>�0�b7�5�U�&~�R*��@������?VΤ��U߫��z_�V�ˎ�z(�oq���������A�=���zFGŚ�d���{��}��x��¬Ƿ��2���zf}C�-b�ߢǔ�����a�8�L;o��Q�9��9%X��$0�z�񛃦B���eR3ϣ�A�rf�0��_�_ ��=9�m'�b��(�r+�rK�)�F�՞Ð����״s�����=^��t�����Q5�Y�3}���>�������>��ik�xo>���gn�3J�c���)+�	�9N��r�Ǳ��gP��3�Ht�W��,3:�M�\Ӆ�|��v���\��+�u��<�9)��Iu���j�g�:o#�w�ɠs��)x|������#�9�tX��S4�ϛv1�;L��5�j7β_�"t{��/�=��|CO��8O����6�w�QE}����n�=�>�4=������ ����W:�v0��O�,��#`�3���b�OA�W��8���P�y��l�i�LJc/�+9���nZ�Oʲ9��dt=FF��m_'������Ԃ���s�m���b���x�����]Q9���/����>$I�R�8�N�+�`S2LGx�8PV���:��㪴���כ~�9+���61�H�W�KH���1�t*�[C9`��c�8A�"xn`�Q�A훦36���y�c�����Tw�����;]�xt�ϡ�=8��FS��j��&��;�T)�6!�;+�ܪ�y�	� ��exm�C�u(�݄㦰�b'�=�^0�ｓ�1ul�n��<=��a�r1�G@*��
A��A;���]D6^wTh=z��~>e�K(��U:��w����a⨅���U1_-��t���i�XDM�#S�6��ˬ�CDZ�`'�k�k����g�=�����(��sf^��ٷ"�+]e�&�@U�Ǉ+���[_����Ƕ�<���gt�u�fs�����m����e��jW^�v�Vs����D5Ћ�SV�ot��e��Q3���n��Vw_��۳:���5C�$[y�^Fx�[�;��܆"���P��:���G�"`1����W�9����b_�ږQ^���5F��?�ei����5�,3m���J�_d��T�c��N��¤ќ��G����`-���d�>��E�W���E�T�[,C���-�n� ��d�y=���y�ő�v����>V
�)p�������g���lp������T*��&����3�Y�v��d����lx�����9����������9�Dz��Ǔ�k�w��\��f	�{��c��99����g�萆�����1v����<=�@c�t�B����t�p�t�q��"�eK7�bE1����3}�����������cP�Ԥ�e��UK�`q��oz�:����F���^j�^��m��q�v�.!C��׷C����m�䋿�;�8����'*��'�dQ���w�y�t��Q��3X=�����P����[V���W�
0j�X���&�9�*��n�q=/S��MC����S�d��ƚ�'%2kT�y/#�^��6�K�w;.�^�:�*Q�Up(���}E3��ڊ�o��5���%����<�\�����.����p �P��D�D�صgoCNU��w���Lo:T���:������^/.\�:&d�=�c;����t�$����^�Z����� �]OJ��욄ͬ�&zW~�`����~������Wt!���T�U����p[���m��r�59Tb�b׷5ܿg���G���>��}^?r����Q
���
����H3�Z{O0|>�����v%������[�^s�͸���j��${!Oԁ��E��Jo���l}�	���k�
���O��ː�����=�.?irm�>��*!�@to���Ć+�}f+�ta��f��Ԗ�uE��z��8ck����0�t��9�z+�|�gXدo��U���Z~���H3�ѱ��
��$����gJ���Xf(x����p���'�s����U��w�e�o��>�;Ux�{5U�y�`
��^�l{k8ߍ�c�Y3�FD�-��<V@o����ec�tu�<�w��҇�ȎF����ul�>�@O�xg�8l�9�'��
G��jz�����D\/(��jv�wWo�d��5J�XS(29��jj���d�x���,�8L�R=��U��?ts�Ѱ�J��"�����A�Q�o�ۀI���WN;��6s�;�&�W�L��75��ݼ{ �ǭr��n���[�w��e���Ԕ����n}��ĺ�&��ޗ� {ݗ }ڻP�*g*w܁K���O����t�v ɧ�#�Mp��T͞}�lg�=�]��@����3��Qc�i�πS4���.���F}=��}9%��W~�#ò����.�b1b�"�uDu�[HC�*��S%��M�M@q��n��@���ysu/�;0[/�7����x�}?P�9F��A
q�+k�z����f-'x�:���wy�%��z���1�,o#AZ�K���Oހ�g�_�
l��w�]=�o��MX;�m�կ�Z�[^2��=
M���ĎЦ��>�~l���tP���\_�8晎x:�`�W	���O��y��3у�R�Yn�]�m��&#k�P=B��ޙ��b���0aJ������
����j��t�pGa�о\������������]9�3���/ofasL����jxPu�	�q_I��p$���B`����B��>�m���ױ��B�ǬBC��=X���A����Q�S�+6�l7��#�yyX��V�ZU�]�����W>���������w�(�`��z0N�˺����pg�\E-\Di*���̔iǵ�s,V�AJ"b�G6�e�%��q~�5x�����Q5 ���ۢ%H��uY{\�߸�e�=��;U��_�[�y�7Н�Q���Qw��T�RX�"������phs-o�jӛ�*{�;���7�Rݴ���x�N`�$h�`告V�B��EO����^�|�M��f��W��L�)A��	���4p��/��B�ݭu���>�3���p"ק�!E��R����md?pY��d���W���~����b��9����4�Ï@���	gճyņ}�Xf�Ȩv}~�j{����뜒���xF�au
w9���
�~�OMe���^��q�Z<T�O#L��X�>�J�ܙ^}��n��l��]�̼�Lt���]WK��Il�������%�g��2��cR{#Ǐ����Dq��q�[ê�a�uհ;Mį*�}4�E%�F�B�B+9Q���ݸu{N����ֳ��O��E��l�.VOW��O��0(�!�'�@IA���#kdT?h����D�cw����0��O�bU��~����z�����<`Eǃ=4�#���Ś��.��ϗ���Q���;�@g�񘱋)�Y�t�X�`8$�q�������9�љU>��C���u�E��a�	�^|�,b�+�^�v�c��Ю�lE�?e���窇F!A�Pj�� �?*��L:�k���zϮ�p�ޕ3'��X�U� *�)�H$�3��h8அY�l�:�����z\U�v^6���˝w/�82�q(��l����	��K��F�i��j(z���=ۤ��N���n�9(��ec�^������rBp��dd1#eC��v������ŷ)��"6�������������K��@��	� �Ң���U����ﻅ�
�v.z���[*C�ڋs�F��w}�_�ސ�g?��GE�
����x* �@64K����4����Mp���s����=���(�Ʈ#��jfc�-���dk�4L�U�|�	4Ϡ�
^�t�8��r�s���������X�Y��8����_7!����9�٘^� �!H�.O�lb�.���Q!��e.9���F�zl{e�j�X��X~W�a�.:O�%��I�L{g�/\�i+C�0_�'�H�w����*��}�W���cS����b���xݭ �C[��7�G��*eXiW��ϐ:dީ�.ǧ�(K�ExT�0�~�Cx6��)����gF��m�1�ם��=�HzC�^����7�b� ��S"�>�R޿���uѹ��QGW1n��鶽���O��P�fkK��8N��W�oN��9'�ƀ��>�"� �5D�U̪��	ګ�$�`�ؚ�&^s�ʮ���΍$�zV�J�9�GsR�Oۂ��׬��j�MY��Y%���-v�Wn�l0
�73�T� ���ق
�*�P����ˮ��lTeVj)]��ZI:���(2o���Ԭ�R��gfi{�c�������7PMV� ����j���
j/�:nn��z@���W�iؑALG�EO`ی~� Em޸�N�-�tX�BA�[)X[nMN*�\�"��\�:������=o�*�0f�.��Q�d�^��{�,5x\�z(K��WPp�nX�-�$]�N�M��q����t�5>�j�����eGDE(��IU[A|��~�Fŉbv:�k�e�*�G����Ic�Y��������;'{���#|Ǭ�)���2;d!��+:~!��=SQυu��e���v�5�gyi�ؿsU(!��Qc�Z9g���[n�AG�s�@��ʨ��R��c��r�C�ޘsk��_��b	^W?V+�9�>ī��UtZ쨄��1�DDpD�Z5/,f�9^l�u����t��0����-�<
�;�=�?������R#�Q=�fc\���E'UϹ��!�h7�W�]Y�h斗�ZO����R�7�bC��y~����B��M���.Y��O��|_���r=F�mv��g�TE!��jϓ�@�V�>�o<pi�p=��1S6)�$^1�z����r���C������^�(�E,A�%na2g����ٷ��>˘F
�%��l𧗾��hױlװ@�u�J��sۛA�VX��r�ˏn@�wfɁ�1�.�NC#���:��#C���;��ö��H�����U�� �����tH7�z5�cb`���]��'g�\��(�fȨ�X\��u.�9��5�^�8����x"�U�^�o�61��2�&~�#"Fѩ���:�@m��k�B�*���o�Z�,�������T�8������O��,.�x��xe���x��ş%<\MG�Uo��J����`����X�+�:e�E��j-��j��Oa�#ÎAf��'�g+\z=q��_j�� C��b=0z��h1�{�x�c�i�ϔ�2�>�p��n23��WC�.h1Qk'��Nk��j~	19��|+dWx���Y!�*h��m����c(3�ҷ���1;��7v�.ąU���Cz}�ϧ� N@�b~��󍝞���G [��.:Ovd����w����~>�8Ƞ����hz܎��5�]@�@�@��pt���=i��g^;���Yj[6�ϡ��}�\��n�������gĎ�4LH>�C#����b�UF;��&c���RW�Ƙ��H������l�`�T��u��#����+�"P*}� }�7�#��|=�Âvv�2C�p�����<z�ًD��;�/"f���E!ֵ`l����3zW�A�]bhQ
��v��+�<�*"��g��t
y���
�7q�X"��b>ÅC��(V����.!��[��Y}$�Q-��o�֊|Gd{�eX���of���%�1�[�1����Q�n�mss&�`U�ă�4,��;#O&���� �}���w��W*�ySB�-�mʃ��aޙ��%%b1}��� �̺��t�8���SC��g�@R�A�d��Y����_����U0��X�VT�[�`��;��dQ��u���� ��H;���ŭ�f]Nbk��m=Bu�s3i�6�.�n��]P�F��m����,�M��[�4=�	�5��U*�$��].f+3�;��M�W�|��9( ��Ȇ7��n]Y�s���9�Ã+:���k�;vF��U��Kʋb�-����c��*�/�Kr.�W*
�ywlrpG���v`��-5�m�Ŏ��`4s���`xe�ܽ�f�!X�4���l���ݤR#��"/)�*{+	����a�h(x����,N��)��AͮY���`����,����pM�L>k4�3Z����6c�| g!��Kk��� �.iW꓌}�F�b���=/u
)�Ί���N㚊�YG5�8�����H�vP��v��(u�hG��7�(}`�D�^9sA_|�Ğ�8in]�巌�ʧ �!:�"���I����b�z39�,�w��M��ʓ�I�aY��U�LN�4*~�]3��K��3�Սl�D6d��z��8M��M-�� �Q�5}]:��^jx���s3�)���Uq �����(k��>؜5/Uk�[�����o]7r2E����-W��w�)R{u�Aa+\zDl��n<�k��Jq��}%SV������]>�>��$8���`Vu=u�"��w� ;�6XGgr�at�eC�[xy����
�&�dpwVn�ԨL�H�i魀+EVK7��Шћ:J�+{���s��2�hv�r����5`�X�Y���K��s9�]:�_=���� ���x@U��VWl��,ؕ*�I����s!�n�8�Ǚ�7xM$��$N���qKO9}ڨ���ƱRH
ܽL/�u�*Q�t��t�r��>�1�仯M���k=� �fs����������j�@�y��Kk �g[< ��.M\����w�lӂ��Lj�<)�v�Q�,�3e�ɺ�m&�ޮpQVx��n�����<Gۊ1V��0�I�#u�t%�E���e7�,�Z/y��LO%]��'T�Qц���˽x��c�Z1`XǠ��Z
 !��W����ft�E��Y��l�)�$͆��5	y���.��.y�K5��ԟR��$�d3����.]ήֺ�=�*̭	�� ��ړR��x|�Tj��J�`�vE/�J�@���P�1����K1��sk[&�rh6WV�C�l�m�s�������u�j�lb
)4wb��:][}=$�j���I���������M�?ZJ+�ű������
cI�"��������SE[��k�F�Q�h��h�&�A�J��j)��ю>>>>>v�5�mv�F�]ڎ�����ثF��:>��)꭫5-SE1h.޽�!T�om+��뢚
t�*i�LIZ(66�h�$���=�%Bo`�l��UACTU�F�Ѫ`�F�̔�\IZq!QO�P�G0j%�:4�m�J��Jm�ӣPhŠ46�zwd�UMS�]t4��@zzQ�4�F�4�"H�&�����qw`�B�J(> 
�Ҙ���}z=f݋��Yu�-f����
��ߺ�1�&jsM�Dd�xh��{O+Z�ܖ&Z����#7ڙ����9u7)���2�
��]�H�]��#!i��5��
B�>��B��ZǯL����1g8�ۘGlv��p:��;�����R�谏`?P�c�n��F�ٯ�(fy��@�؟G��Ǹ���6ǹX��+l������ؠ�ۛP��ډ���<<��p��6�i�cND�����bG���Կ���P�<<��U�F��D+����ɷ�y�'5�\>�������.�Тe�&'FOA��}S��+v~m3B���t���3UF�Т)�o��(� �z,h8ҩ�ǣ��M��Ρd�Ф
��[<}{R�ېf]Q�w���3�/4���SZ��
�%���a�J���E�gØ�Q�F��ڿ�ώ[��U=��!�$�����ׂ>�Tj�úXgc>e�o��m��
=�#޹�+��Ƙȭ�By��-n!��0)
�&��_�4�V��q�/���!��Sl�U�x��q�%��ks$��,=�hg�]C��9'o'�h���.�2�[1��=�u8���p��3L�g���9r��l,�b��2��YԮt�	��
��9��G�(!>���"�����Q�"�r��z��웩��xl�ҷ�07E���������S�OqJ;�u��۾YKEk�P�z����)��Л�����!1�w�⌻��E@�&��͚`S��ng9f:����<������\;v�D�ħN�����c2��o�ʏ�Y��)Tw���mH����򮮮�������N�i����>������e�T��(�a���H�O����=`u�A�jg}�O�������Ts�L&;��V+��%7�2:(=F��ھ6OA�@��,�l����1�s�?;>u�Z"��\�;�u�ť��W}�����?V�B�`hfI��{�|c�kZ�NК���8`[���9S!Fq��7Ū��J���?��t(��`W�僱�¦��qu�u�k��V���lG��c��D)p��
;�`gg����C�z[)�ǖ˴���*�׆sμC��8���
D�4�`�|ʿ��!���@��݅bN]w$��Q�����#���;s[m�e�B�-GAP�dpR��Y��=�z�!�ƻ�}��R�ul����JW��8�{�����b�U�69ULR�9��(�4L��Uh�#���*ޡ+�n��ש^�v�>9���P�w\@��ӈ��	a�C]3^��u��56DFty�>���^g�xH�9��qf�=�L���w�F�zl{e�j,/K�~�a��:W�VN�q�|SX�u<�ᱛ=�Ӛ��Y��C*&k.�>��yQ5�p��+v��u78��Xէl�8��M1ʶ��Z�NQ�0U�:/~��Q����]�{��५�Qܫ)^�I/�MKfe���	�{#U��0C�i ��[ɸ������]}u]]}P �� ��b�K�i���&zN�?�K� `-s&��\�>����z/[���[,C�~�n�G����&<����[���͚?��h�}��U�_��|"4��:�7��.��9	q���I���$�����������=@�Y��?z�u�
2��^�|~�jB��*z����1Yϡ�'Ьq���ϹS���^��{����d@xw�-���k�j��[�ϰS^��Y�#�DN����N���T�~Fj/��p�6����Nqc2��v�S#��f\\y���5q�n�(B��(S��qɿ���\x.�-�f��XWP�r��"����#��򸊿#�|1`FE1xK����8V�,Z[NH�����8�F'*�A��s�<d�b����a��P�� ��;��d�b����f��ʜ��y/X���9n�냦��+9��g�!�����#�E{��'`u��L@ �={uq�*�\<�����Y�����;����sP�*��nR9f��ߞ]DoH��=�h*���v��9߽�wO�OO9�M�S����I�iؑ,��ںxQ��WL��o%�
�b�+F�|s
�QΩ�L��.��0�v̽���u���؃������j���b�t;r��(Ғ=y��@:���p�ltˁ�0��qr��m|f"�ű9�ԃP:HR@� @ }��D}����i��ۈ�}��]S��9�>ī��ʫ��eD+�N0��" �
A�wB�i̢�;��Rޝ�!ݗ�Vy����v�F���-�ޅ?R�ؑް��ԴNB��L*�ut�����P���[�æZ�H�y�_M:�pmϴ��K�~�1[Ҕ��HHB�-�7�uj!t����C:�i��Lܞ��3�\T1��NCf��<qx�=�WV;Ԡ-��1+�Sd�{�[�����:����U5�?_�\(=,)pc�eǾ����u�q�گC���^B���珻w�1��Q�j�C�9F����c�X́�xe��Y>2,`-`�'��-�n<����VY�gQ��=��و�w.o&���Ѽ�qo��S��]>�ȫ2����a��[#re�.;�̈����ey`}���m/�a������6���ո�{G��pHk��hR(�=�ߺug�?�W�c�O�L����6�=Լx�e��)�egϨ\+�q��#^���T)���l��?��$���D������#l
��l�qS$W˭�g�f�NE�{�2��x�G^����p3��-
�@:������u]������2�hc�c�Ű�$s��V�Ư�oPai��m�+g��qh�y'V�:���'$�92v�A��%�^���`�SD[0��QHj0�c9/oq�A�.��O��KL��5���<��yR2�4@����_}��J�
D Ңҟ�W��~��lG���߹�@�O������l1?H>S��]X#�/�~���k��{�%D�d�V�c�g�m(�-zs�~�H��hu���)t��r��8����q���l��:�%�7�D��'�N�3<�61��rm9�6�#��5�1?t�	���� �z+��+���/f�vGc�8�Wb�Y�/
2���c0ySG�������wU���b6�`F��-w(����}���H����u�x����ˁ�h/�����)M�_���f����<	 zVϻ��3�����24J�*�c��g�{������!d5W�;��!s�y�0Zx��5���wez28aA��"~F`�	PbG�ʊ���m��ou��_yyX�b{�W0���W��<����x�!E���Z'���W�Тe�&'FOEMKe��F�[�e��O��s*L��˳O���x��+�R1�ס��U1Xv1���+�hY3�U1>�sP�z�3�}���V^>�=����������k#V�`�^�!E�����l��C����d��'����M�`�6i����zi��$��K���J�k7|����H��^Y+P���{-Np4�=u�:��s�(�����Ǉw��)\9NN�-��9�c�uyZ�
gsi��P���1�хQ�E��g>(�9��C>�\=L��(>����H1*D)�R�Å��W?3�W�	�4$���]VP}�鼋�v0!����"��}~�j{��ԟ]bs�� ��� n_I���z�EXL���F+z�zK㧥�zpr�e�����=;QU�W���hY�n�ˀ�C�W������bT}!ʨ����+���C:�tX2��77{p�y]��/��r2U���!�3[��]�Fd�zw�"]����E'�a�F�B�B!�:�h�m��_Dg��~�wД�68ж[��vs�FY�o�KO��������|��糟�M�1c��T+�+����`	VCE�##��27��=�'��BկM�%���`��J&,B�}sh�W��Ӂ\1S�1x��5�'J=�Y�b3/7�]�*lEz���8f�Ő\ecjP����s|^~���|�t�}}
�w�0H�Ł���|js�����0�|B#�����Hr�X��ѷ�V1�.����_�\�{\hK��7VY�{��g�P��}��*��	� ���E	̭��{��P:	)=������0g�ʕê>�\[�7Ut>����t��8f�{�8��C�t�r�E�~��ê�\�!����ͱ6�B��-��3*�w:��A0A������Sn���&tOsl#s����J���'s�e�;���������ߣ���F%H�b��)@�D��	k�\߳������L��"��+�谺F"���I;�H3��p$������RG��C���㈔o݂�s�v��Q�*���U1KD�+��dklMɠC��^�V�``��縄�C���Ð��5n�@ខ8���	�7!����)xNC�6fEt����f+����<D����JGn�<r3���g�@�h�J����ҿ�ލ���~03���+w^�>���(tDb=���	p0Cdd�U���}�^��H7��xs��6�nׁ����Qf%�ڪ�^ic��m� �z�eM�w�pe�r}���
�,���s�7,w��vOBm&����U�w�Q���̾��.��~7�b����8���������*'��ܭK �d?��7�(���N�,�N����f	�{��ӳ�k��!gm���b�^;���hq��*Bo��HB�s���[/�3P�~���ڧ�Nq�2�ev*U�s�r�������#*e�H��r�+[)���5�6ˁΥ��G0��c��l�.�6r겅F8�� ��k�i+�8����x͋�Ƈ~�4H�J�,�ފ3
��s=����Q>Qz�k�.��ݧr90��Y�O2�Q���H��%<X�%	�<[�u,U|{x�t�)�d�]�rMǮ^��\��lG2�(�Oca�Ƴc��������/�H$J�B$H�P5�� �l�>��q6-׍D@�?�7��#�R��뮠�Zܱk�rE����)�zO���)S����ꅼ#|�힓��A��A��@��@�\lW��v:���x)W�(�YB�0�m�'s��]�Qu|�j�4#r�<����.�[��:��QD�H"~N��O�!��۫�ofg�FL{)���<��{�����Bs���K��ܤo2d[����F�N@=C�@�8t��(O"���b�!)��݉��rT�$o�Ր�S�!�Y����ʫ�u�BЧT�����O_�b����H��i&���v�#��"7:R=��H�;�SR�9
/v�$1�����hf<�ɢgp'A�SN��n}��%b�� �>��H��	BG}��]��f�)&�7�jo%��g���nM?MA�%EC+�$�6o��]ΰwٹ���H�w�	��V��������c�R���6���Xf+�5pOZ���֎c���ˁ�c���8;~;��:g���Z��m1����c�X͏�/�Q9�FD�����l*Ϧe!2~ɹ���cÿG��̔�f���b��o�T�^���+����&*V�n�25�r��33�c;.�\K���te3���m����]�����yVf�<%���[�C
�h�m��۹�ewn�Pȕ�=�~}���ߟ���[�����H���B��JV�H����u,�LLLA>��q�;�����'��q��QcUl��������p7��h0&�<�}8�X>���]5G��]_���	�@L��hj�X�;辙a�c��4q�W>���`��E��a�+�=O�< ��P�yK��"�O�Et�1����BΥ���e��3L�}B�g^~O$��N�c�=�X�~��-Ǣ�)%�?HhM	>��Kʈ��\!��0Tɑc��_��o��M-y���S��h[[]��]>Fϧ� N@a�� \n����GpTj��^�;�g��7��=�F��6������>�����Y.�EL9$��<Zc������s����������yW �Wљ�M���Óa9�6�:&8�����wZr�ndM!�[���H�1e���Ų�R�p�Uq~ަ�Fy�X\����}��_�a n���G� ����&<�C��H�}�RcO3
�*Q�\�f�t�pFF��~K���
S}����t\�)"�����W��ǬI�^��:|�
(I��7�0���+�T�	CGn�'��ߑ���X#㯽K��{����}p��c��;�q�o0=5?u�bX��	R����9^�J-�9�5�`�I�wd�r�2;n���Mp���E���w;�K�霧�3-&�6��v.2���Ad�n�����&A�{��j���#/�TL�O� � �B"�hF� ��
@|" ��nsu"���1��kc�q�����H�0t�<���~+6�l7���q��9;r\N~U~���K�}V�X�����)h�F��["Ib�h��5��_nF���ʲ3���.ə�#��:�sٷV7�#�Cm*���c�2�E�
E[�$H�wq�NEwF����q˼������-�-zX��~�"�MV�����=# �i��N�S�q��@h�kٻhy�,!P�CE�Ln��3#(/m\�E��ϖ��"a�}z���u�����q	����o$D�H��4�����;7�/��zX��9M��!�ׇ��^d�ɞ��>�ߪ�﮶����ٹ�=�f�Q�>���ُ}��(gS��;�Uf}[X��zt�R��s5��n�<���Fd�zo`�1/����	�0�#>ڔ!�$�vLOy�?�K�M-DG�G���J�~��ϸжm�V��t�a�"+}2"ND�ɑ����I{��Ա�O�A6ȨKΦ7���bU��~�Q�����GA�F�����7]�1n��k/2�4�7��Q�=q� �r���aιK�Y�aՎ�=�@�ČI�O��z���H|;&�W����V�Q�+b��^u��S%�.F\��Κog;s.��Hc7U6�'+zƸ�_X����V3
�A�� l�C�8�k(:E-�-��t�Z�1桝�[�4�q�v�Gs�[Z3;���U�-)�*�z4���ԫqj��}y7&ʹv�9^�m�4�nɵ6�V*X�͇/-�	$�����z�Gj�;��m�ǚp�|��R��"S(�ϒ��#�f�������p���w}�:�w� u�Nj���bdi��Ɍ�S�J� Mfk6j�S�I�]��.�ѭ�Һ�\{R�32�];������@��6���֪M��3�Z�`�[���hHR�{�s�EdW��;]�L'[M �yV<��\ۮ42���P4 fi��K�n��,�Ep���ji<�>�C�ƹ7r����8r�X��9rftC\����22��޳��{t��t��%3��e�'�s=Z��2�,e�Bud��X.`�ohl�>\��)�O����۹r�ɸ ���c٬3�cw[��)^#�;:�7YQ�E���δ]q;�qk��Ԫ�p�"������t�B�}�f-δV���6�^d��oC�M*��2��0fqY볒��|���zi;ԇ,�ѣ�v�ɹx�hx"�h��y�1�u<5��Z�srk��A�h�^˧W����̉��39��m|/���z� �#F`'眐�{sS����[g���|�^Hvv�X{��k4��7�k������K�#�p�l֙A8�pŹ�NqR�T�f���x�=��� �v���!��o#�ijBF�o(����D�,T�v���s�&��!�Fd	W5��̎�,���`pq9�S.�T���]��x�>�qQR�r̫:��J"��/<*I\���U}�"��*[`P%�Ѯ���4���vlƳ:��s��Zj��8������"�&�nfq�ɼ�=9"Wt����"=P^�v����FK�Ӎ�.R����W\�Uz��:��A�vAa��Zܫ�dV��r�7��/K��������aN�C�+�7�`J���)�L���BOu�Ep�	-�k=[�������4bne�f���n�3Wx⻗4�T5&/:b�ͪ9�U�w��a�8k��w��R�^7�a#��u&�`�0��k5�s�f�٬�}[���m=iꥲ��u�o�4�T��ιV>��p�*���b����/��7#::����ef�jԚc�s���''���CCB]�����!r��x�~�[O6�(���Ψ����s�7�� �d2�N�(%Ip��(T._=J�v�ǝ�	]ό�{c�;0�_1f�;��vanTE���mn�� �2V��7:hֳ��[�%)vJ��L-m�Ñ�!{[��������S����
5���"��@h�D�3D��S�A�ӧK�����������}v�a�4t��Z5���q4��C+������������4�I�h5�Q�ִi�cm��DZ�q#֊�'x����>��(1������Z(�&���U�[o�/V�.��Q8���~AOZ��5c)��ΫT�q4U:4�;h�i�ɭ&�m�F��(-b�lP�32D[;Z�mj��F�m��z�DLX�[m�@[	kSTQ�DD�DZѱ�4PbfJ���t�Iӈ;F�˪1�5u���`�'�X���3�TPV؝���c�T��DT�ѐ��+cZtk�uTU�Q��F �F�b��Ui��5�[4��4bqb&�����J�TQ@D"c��%�o�����[���J\�)>�gR��s���s���]����CD�à{�Yp�#rv)����e{���<چ�CQ
@�*�"�
�*����@��?_����?����]��������BK��sl�YB����]�T��b�l�'J�{fnQT�T���^D{˻��i1��4A��G`���s�o�ς�X�©i��O'�y�P�|�\O*�C[�W5p}���������@��`�wѱџHr�_��:6���<��>s ��껉�?Thcs����7�s�(>�[�=ň#��**A�*�ۨ��G�f���_��u��;��~��C�^p��{��"�Ӻ���Z:�&�Ȓp
A�\Y�du��ߥ�p��1�Q	�1��֠_(Hń�#���_T�|�NB���Q���>q���+�"#D�Q�=�� ���p��	4��l��ﻮ H��^����1]S��5x��1��$13��Zȼu�c�'DЈ�B}�*l{�٪9��{g�@g� j,w�l�A�ʛ�'|'�Ao���/�q�v��_+VT��YC��X�;�L�~Q�F��+ݾwusq�l1WO^vP�%kH67� V}SrU���?1.=�R���<b�����s���L�W��9��u?� PM���sI�Z��6��B���`˞oo1r���t�1���p69ma�9�����gC�o����(�KYHxz Z�N������p�	u.���է��0V㛫�c����,�ή;u��	��w��d��ޑ�����B ZQ"U�$
H��V��i�B����#��� ������5
?�����T;Ջg)��f.��`x���A�aNC�(%�o�c�L��vg���^dFpc��P�*辖)���ebt�8�i�̟X�x��o�Y�����ԯ������Ʉ��v�
d0(��"�pF�z$1C9_�7��/�#5��M�p9J�"4f;���nbӸ��z}�bsq��D�1����(B[%���43��p9Դ[f�Ti��z��
����	�"]G1��}4���q��s��.:�u	mХ�m�x�����U�{��[y��oR������>�p�>���i�){]�����`k�h�i��S�jbf�=��n�c�ړ��H[��l?H蠍�g� �bv}��������:�E,���n|m�+�������zp7)��碀yu�n�}� G �a��b�Uh��'�ځ�0�1�E|�b��򬇂S���C��q�_W��Uк�!hS�%W���ꉡ��8Vwp�"8a��kO��ۘg�v�F�u4{!Oԁ�Q5���/�����7ם'�#!緯�L^e�(%�.2���dP�W�Lv�:<��P��X�)��l�=�3�����o��;�غ��\�K�hDA{����;:fXl=�.��u;&�T/Hõ��:ߞ��م�3y�z�!��S��e'B����� ����hJ#��
�￀�@�(�� ��%	� �T��B$)T�Z�$�JTJ>��D|> �[��nY��13����v	1��%p,��Xn�#�sKi+���Ґ7���DA5#��X�g�}��"s��f�1���� �I[�3�BTTS�2>��s���������o;�{;�Q��q������1�RA��X��ư�Pj�*"��\W�����r$���L]z���S�x��W��$�#���;��X	�X7������:�T�9B���':��.��Z�'����x��OՃ�^�φ�����E��'^��g�����}�c�Q�ѳ׮�^!]c����p=s"�:�B.�A�Xd1�j8۫��ո����X��H��~Ls�P�r������sL�z�Uۀ�(!�{�,�Z��V�_w������g�aE�n�23��WE�}9%q�$)�rs�����`:�L�w��P�H�N���7��Z��|fm}ϰ��o�~�B݇��:/���l�~;_@��,1?Bơ�}hB��]�v�R�n�r�BG/K>����]�?\��N3���"��>������z�+��>���� {��昨�z��cs*�oC�a�>���ty����0nj�7��������E��A��EFn�d����O!5ύ����������6��F� WAϖ�g�x9Ago/���U48����{�C2PC�{�IܛkM(�j�퇿�}�U.����&h��"A(B%BeV�b) �J�
h�
�R�H�QG���@���Gw��K�碈��5Nu��v�����:M�)�q�t�!3D�;����˸y{��1�������B�_ҕ�?oSg������u���#�Y��ь��n��N�u��]&#��8�����cKFx�;���<�@��B�v������#w��c�|_�7l������ն$�ZE�eu/T�+�9�t��֑
�l9؈��fC+5OTm���B�:΋E�G"@�0t�f��K�^ۡ��u��n"=i{ϲc{7��_���"��N�Xգ�����_-��M�^�L�D���'��Q�{ye����"-�˃�4����ط����7^�"�U1X}́ưʽ�d�D*p2/�R!g��F�τ�Ñ���w��f�-�[X~�!ŧ�BS�:=���T��tr�����|l�G��	L��}�p.�(%>5q���b�a��T9_��_o]^�鈟fg�����0UE�pc6��* ��*�R~5��q�5�Ë��Ɩ!�֪S|l@&��w�,�t��ٛ
��X(U�1�[���K�������:���#�bO�[��if�BTY��.�K�0������;9���scJ�%,��M��RX�4�t[ͫ=8,�
חϮ+j2�g�
�R���3l��4�.��������������B$hDbi(X�JAb@h@h�)T)��V��(D�}��G��������O�{�ŧT�T?\�p뜒�zv��]De�
�cjLp��>���ßxv��5?�eƣ�f�X۱�;L����
�ND���}4�A�[FI������縦O��s����ǀ�n��A�~�Bٶ�XY=^F����6#{�Y8"��3����7�����G׷AV�0�:�C:����PGG��׳\sf)C��N�bVIƠ�d����|:��X�X��m���O�ŌYM���(C}��i-�~/�2����n�2LD��� �:���d8�o/��cKH�	;P�Q��r.O��1�^�����b��
��X;8��`@�@�wѱђ�V+�tm�+5O���&�4:��w�/����cH�qʖ����ϩ�@��+c�6$�xO����A�),�s�1�uǫ۱���ۈ���pX�n��z��S[ʦ:5t�F��)M�
A�+n�`Y�����33\]����A*�T<�j�F��àr����rpQF}�'~������6���F���ܙ�y�xf��eh��(���>I-X�HP�o�[�Y�j^S��� A]j�X��7Em���2Q�ֶ��_]롚���h	�*h��d�;N�����h�V����8�s�33�μF4��g��������}� �@"�ҡ
P	@�$B%"#M(�� �����X�>'�"�̘�}�W�����4��$�!����Y��N/�u�+������w_�v�U<<2�Ԇ��hr*�O�2�kY˹������GzĠ�xy�/&..�Yl^x�A��W�P��=�9%�9ᢔl�>��	I��豫�?�G���i��4�5?j���7��-��P��'kH67� Pʛ��f��b\z+¥E	"xǇ���J���o"����Ű����BB\{��	�jų�S�X���7C&�����vj�N��U��o��9�F1�I�r����]�K�e
j�Y�t�8�i���}^���2�6s#�g�.Cr��Z�BG�%�#"p��*B��萆r���T�~�CE���V1��;��z�y�" �`{��h�x�9�>/�;����>=EH-��b�Mw��p9Դ[�ĉ�2Θ��u�GcQoS��jzʋ$F�qL9��<����+[�-b�rE�h��;��ʣ�R;|�K^����
�R��a�D[ ��}6.xN�^�Z/j�+�=���	t
\�^%�Z�$��ܧ&TNp��#��gUX���!�9>5/+&��UoB�A<�x^��q�:��q2��ak�5 y4����ېpuH��F���O�N��&U�4��x)oSkt�"<�_<4zK�bՋ��S5���?��[�¡�b�F�Z"�F�$Z@)F���B�@����R��@} ���h<|�������}G�{��sw�c���~�v��:+�l�=�K+��Oʡ��B���)R�h�c�{⺦�'�+Q��u�9l���?x���w�-���
<��B�;��fGW�8`�k�����6�	0�E꘍�u��Jv�z�hJ����WE��Q
���v�:<tO��V�A�" �A�ÃBMi�9�0�Xݡ��u4x#��yA����8��wd��^�q���t:h����O��)&�y��}���BC�~�1�Gi{����d@�]�{�tQ���s�7��0��?V�ܞ��,���'!�uӞ8�d��T��}~W7)wz7����ۈ���J��a�j��k���o�5�cb`�	�c�ˍuy]0k�u����6�s�8�߼u��b��ʫc�Ի��[LC�u�
-5�Ƕ���2�u'�T�\����׫sʼb�D^�''�B�ۿ@o>ۛ��r�s�1>��U��|)�z�� ��܍nG��	(���0g�&F�����j_�!ާ}�L�ȿ�MCGuqlZ�Qw�J��5b��xghDȕ���T�������	�D��%�ܣ����k}��T���ɳ�v�q�&@1��<툝�۽{yg�����Zb���Du��N	���s��Ѯ�v����̓Ձ��_�����߇�����ο7��r�HJУ@�J!@,K@B4)�J- �H#B4"��HH������p�1Ւ�3��E��<hY�h"=�i�X�p�PC:W�e�Y1��w��}������x��[�8��B��j��ޮ�>�����dX��#lV�v��~�9�Ab[x�ӯѽ�M��C�۾G�L�)�H��=���.�#g��ځ9 ���e	q�W��5&c�1T
ڷ���r����Y�v���\t��%8�?|�L$e�4:�}W"����
~��{8�2�+�#/x{��%�`I����5	����q��g�Vћ�|�X��6��gĎ��1�ҳ�]��8��������o��k�0�>���Ԩ\+�R����M��j��?b�b�^���s�^�����U�7�8X���p=C��&4�n�O�;U�G��t�+��~=���H�R2 d�5���e��?��ƶ66����&:��A����E'c����;~�bz��d:�2�{�=�ފ�vH�#��@�člth�Б�H�(�������������,y�
�`��38�B�u㝝B�����*�P��#�D�7��KdI,@1޳_^N��w���2{2�;	{yK�>�-�Xζv�B�9���C�Y��L7o���l6�oec	�m�t�&V�3�e��X9�[���鹐.D��X��M��چY�M��2�uӀ�M�d*�ø���Ҕ��%r�4&(�㟿������~�����@**D
$B@� %��P
(R�R�]�?�������>�Gb�Y��8�u��+������qcz�����_�*���ь�k����tC6�Y�0��V�1$�8l���v����r�+��ݛ�_�e�E�K��~�"�j�Z�n�1:-�t�xo��:6_�_�ddl��`��I����U��^�ȱ�Pgc��ݴ�vQ���5>�{k��^�8�\�`U�Z��������<H�x���;7�/�l���P��~���=�]o����Zho��[sh�
�4���{��:�$�>�4%G������:��xԥ�:ᕞfcz�tXS*8��V݌yN�#2z�)�(����νK u7�"��{������x��؍��B+9ъ�����!�o�4-��VOW�тg|fU26qA�wސ�ߵ�Z�����RX⯮���ם�Pκl��!��,V�p��f��ʌ��8K{ �G�"�.�6^��|l} ,>��v�L��_�Zϖہv1S�1cSf�Kݽ˹�'����}ʏ��?E��X`_&#�����ߡ�`!�#}s|^ ��1B��.� ���Ҧ}��vh�9boe
��C��pVP<�XxJ�w[�t��e-�.V�+��ԥ�2�tar���>������v�&�.[ı��qyVʰ�ȥ�t�ɕ�)LY}��,����-�կ�������s��J��߭��;���D�J"I 
bH��hE(�
B/�菇�����'{�`~�{���[���+M
���8b�/����F��H�{�9�wT_�p���10z��Y�.��r���Nz�+b��t���Al�.'���N5D��`[']D%��@�M�Y��q���_ܮ�������
R$��S�;�NGy8���{�ըH,�?������G2�����yz��M#ʌv��U0����Ѫ} �!w��7�t,Y�p1Y��@p�]m3�_�)6w�p�@�nCJ_�q����qA�=�wl��.&3A��6k��"0x"�9�YK1��e]��	[��bU�R��Ʊ��g�4r��3²�/�z��}2v˾!��8���W��dO�|��B�R���t���T��(��j.�Ҵ�~�o���ʛ���b\z(xT��&<r�i8øv$���]y��z�	`wQ�b�nr���X�s��Z�ci�kGX�D�
V+M�W���w�y���E }$r�����Ȯ��b�,�^7N�ӡ{>�x������c�ܨ�mL�I������9�9Z�!B�߁��B`Ens16�fqM�>��*U�锟Y����Y{tB��^(��w�l��|(�ЊI:�o�4qP�nރ�ř�t�1O"���n�D�S��Ƿ�s@�˅��Eh%�B���6v�� 1t���h�f]����|i؛�t�%Zz���׀�t�1^�-�W[.-ۇX�o�
���h0Wb<����m[Jj�G�q���<�Y�aB(p7m��pr%�#8����˹r����5]mrʵH��骛��cn���]$���}z�O�#� �R`w�o�ލ�f�%�`pw8��7��rj{S{�,QU����{��mܠ�Lkhی5.��oT� P\3�j�
�c6��f.N�ڈ��6��
��x+��6�B����kXE�f����T�%�yG��y5�z"��ͽԑN�N��i�b^ù���f��Z���
T����za"`cG/- ��pA��S�3wmUۧ/�f����[��v�1B�����O��R�Co.��n��5�B�(7pu����I;��Wp�Δ�:��|\�2phlp�y{L�Ę�Ϯ�z�z�q(J�����[��*�+���Sz`�(�<d��7�٘j�7��5Nde^��id;}t���2]�-�����U7�!lZ�-ڋ��]*�p��(efV���S�60N���*�|�,ȶ�x'�<��T΄�I���iXP@r	j$S}��ݬ�F�4P��� ���8ᕳ0ɭ-ۧ�C^=���9Q��\,V��U���l��v�f�MY���eۦL(�ي5��e>�����p+4Sv���*�F�=)���9U�,ҋ��V_fQ9;`��Ɗ���N�O�d�P�/NKH���0��W�}h��4�Gm��$��yY�[�6�wZ%� Ѧ�<�I1�z�,:��^��B�wvCV�Vi�����wԇu����K<45�n7"�6����H�`��i�K9�2�5&r#���W�:+��hR���Je�U+C�ae�ܴ�ШO͘�_,1�4��ۣ�Y7�b&Vm+�{�)_qt���(`1p�+�B��,T������Y�nLFְ,j���6/#���[7>��fM����v�*�r��C0'g���"�u�+E���N̷�R�h���첯����|o��͠�}����$qi��5��4⢲��e��x�ʙxr]�JuM�	�G����N�E�\+���:/�C��ű6s��9�AZ�\�*��s;`BA�L�{f�PV��
.=-k註��#ys��Z͹����R�MT1����X���.�8ܘ�`2ݧ��B���e! ��:��}�)g3Q�Ӿca����9��oN�H�4�6�L�5b8	�Ƕ{M��E�Ǽ�d鐘鼇x�n�Wp��^�%�wkP�k4��3� ^g�_pwfdQ7C��]҆��v��䦥�FD��ә��Z���((��ˣ��~~?������k4RQ[Y̵kTQ�G�hJ��j 5�l&�)�A�*�g>?����ɨڰAIl���$(5ӊآ��Ղ���[kI���4h���||||}�D��U~l�QF��6��k�Tm�LI���A��Qbu�+�i>1������h4�gM&�o�4���OF��qBj�TS8��TQ�Z*��<|||{�b�
-��:i1[h�T��rSZ��]��iѶ-�F��M�Zu�8�i(���DF$#m:ݓ���f��cJ
l�h�l�gC�f��GAӢcw����]�N#v�UDu���b�6�QILZ{e��;;b�ڢ
.-�F�F�j�+Tu�SA�5�Wc@h풒��vƊ���b���5�Pm����U�b;�J�cZJD�md�l��3=�;V
�;!Tbmm&�h�6ڣwu�4������Y8%����c�`����-��>F`ͨ�<]�ގ�Q���"ff���s#�� k{h��M����VO�F>I�Kͤ��죦�݉�1�q�9o7E��E��A?ꪾ�uU����UԢĥ @	BD ���G��#|��lO����k�Ѹ�?h\T��;�!�_oL�WA�\S����Î�r=�)ݝ�\=W/ ?��x�9�,�ӱ"���!b���7�(B���
v4yc&�[6�����֘���ߚ�v�to�u�7�z�c�=eE�	ِA��Ø�E	�.:zC��-��d{̍�s��DG��c>�s7�I���I�m��NT+�I这A���	�����	�;���f��e�������Q����=��39;Rq��v;���#��6A�="E��������P.�u�x/�<}�5ӵ�p�����WSӁ�H�g�@yu�n��=�!vXY��"A�8x��c�Ez�I����Y)ۅ���`J����WE;��MT�����|��(�cgu�Ȉ  �%�BMi�9�0�nȈ�Φ�gЧ�@��f�޻���LͿyG{�������a
�L_`�
�h�ĨDj ˛ӵ��-�B�3ѭ*���_bS�L7�����+�]fh��l�����J����J�r8U���C+[�J����fjJ�}��W3����U��:�'Ζ�
STیt۔�.�ՙ�_7:ཡ��\�٨���~��vTǭP~ai�W-K�P�'
Hm,`.��eO��1R�-�ٓV��;�O�v]؝��O�T�/w�9������ځ��- �$B�A��|>��>�F_��O�:����;�߷U�U���_�?Xb�j��k�����L�2�@lb�Vm�]�ҡ�(�P׏8Kxȷ������S��{3��w7q�m1�נ(��^�o�mc6<o�
�9�܌������`b��H�)����
����7��B\{m��!�}�l���Vo��F�ʒ|�4%��yE��xe���x"=�P2�B@ֽ���S��2�"�MCE��%/,�������s՗�����'a���`>.�%}N��)�#�p�W�!c�I��\�?=�io�Ui��E"��qxPC	�ո�)v>���|�*������o_P��^0�ƽ���_vf�uU@�XS:�D�	Z�ϔͲ���Ź{}��]>F���v�	�����{�y����QO�HF�[^�G>]LP�S���)�u��h$l{S�����z�j����l^F��`j?�\�(Ic��3���W��_Fey[Fs·C�'=��>$t�X���܁"�ETFg����_�&4�0?{Du�&!��]��R�p�})^F`ަ�Fy�Xk�"QV�������dO���;ܝ�*��q�r�Ӕ��f��KolXRsW͊5М��gr٭ZXV4+��e��#s�3��c��7�W]nԳ\�%�6![�i�2�s��%��K�βk����0�� 3��~�^�{ߏ��������%%�(B%
V$"@"��_��Sn�`x@�?�b��v6p����)����r7& t>3�����XǅӁ�<7��]t�옏m�s��#q��X�u��}No����a
�H�����
+�'c��ۘgM-\r�c�F�Vg��ߊ���Bl��BGm���/�FƟ_�h
����%�U�x�;������2��%m���{t'��#�/+c�Z1a*�QIOI�N#�6e{hQ9����TU�m��������7jR/]z7
�������q{Ըņ���XiT�>�f�@|��v��~]��������'+ƕ�Px)�X?x�k绅��e�B�br~�#��ܺ�WR�c}��b����YzFP2���g�H��-���VPK>�M�^�A��<�o� z�5�t!WO�<�Tu�Af���n��ap���_�ER��u�+����r�����1���,V$��#ǩ��8��-�L�ʁqa�W��Ľ{%�g���%��Ҫ#;�/>Yx<"sw6���<��c�ͥ�.9��M�Чi���2#~V6����}E��~�u��4�����g��̷x���G�6�:G^e��Xb5�j�ux�^�7�Rrf�"{5��k�۾�f�s�0�DC�׻�׮(���z����l�\Pu7h=׵����f�(]�05�7����C%m�z7���W�*��� ģ�4
�����>���z�10#q�M�E�B��b+9Q��n�2'�"���XY=^�R^e�Wtz
!a{�����^���f]"G�	�P��=}tF�ȨkΦ/�[5�7�h���y|=���e�m��p^R�>ʽ6=�ȿ�!�(Gq�����W����p.�S�1��\�:4�Ū�����>�^��N��~��fI��h���;�8�9s|^+��A�^#�ݪ��'^y��n�E���@����~�~��(�� �� A��c��\)������S��ugN\�1Ϲ��
^�!�=9�r��#�
��迸�'�r�G��L��i��g��E;�"��S��֠tX�n�τ>��Ϛ������:h���A���p�R,s������XC��;	�(���C���ö�:�z��9M#9q��r�^���w~Hڔ��'/7�w��2
;M��Uh�#Ri�@���C^�$g�5cz�=��	BG��P3W�׉~�W����j��S�o�DA
E0qs%���s�#=�>�d����'|,�6=諠��ʃ���N�����#Jz��Va�y�2S��ki:��Ho�E�D+��7XO��=`ԃb��M��q��!�dx.QG�J7��b��b�a�N��qMK'�5�*����WwgM���֊Z�4N3��~�����߾����?�"D� �H Qb�:h�4OM��M"��Ȕ勆�7�%SC��)+�(d�&伮V
�^�ߍ5#�Y�y1�eg<���R�l-t���i*N|�X�c��x�� ��GV@���W�Pe�q��a���=UJd�勞p��a�"l�-�x��e�dG1.=�r���T)���3��6<o�_De����UM�a�����E }u &(w��"��t_K�`�Xr��ÝN�1�[*9J�I�1�7B^Y_Y���8L��?#��#�7��oz��̤PFcc��YJ�x@���z&�V�|�^��NqeJ;�z��pr�+b�;�_$te
���ْ������h���l@3	g�a��*/��dXhC����'�o��~|\T�u���{�%n9?�S	[�.����)�z19P��Ԥ�8AŲ�	��@.6"���!�_QYi�k��C�L+��ҧ 8��c3�Nԛ���qU�ވH�!G3d�0��ƫ�L�����[�,=���;O��\k�+��C��z˩��Ԥr�s�A�-]��us�j���ҁ)s�r����~1��P�m�j�.����)�&���P	󗋬���$��SY�e�x���fzb�kI&�x����hw�^y9�D�/�*�qOXՋ������r���)�cm�9�f��^+p�ĺv.R�����X�A��ƽ&I�~��߿/�������!J%� �Ec��Zuo��@����ycK�����ud<����9�2}�/�~"��o&�S?~[��D���1�N0��" �R薍I�>G>ۘg�v�F�Φ�e�J�Y�ys<���ې�����M�KD�(��&w�D�@�Ȋ�u�ୟin������Y�62swK������@�H��$!_r�0�E��l������QQ_1�Q�������K�v"����E�ߣ4�Ū�>����C��q}�P��a�j��hf�3�YCBe��=츗W�س?nl�+��='��.j~�}�U�����i�w�:����~��}�Ŵ�d�Rw�	k;W�ZgϨY3��=����HmW�7�m��_w!N7>�LC�ƪ�;6J�*^*Xn����T���K{��n�W<�K'�(g�����e#��5(L����h!c���e�DW�MCRX[�1�sr<�����_��WZ�_}3�>�㐄�����#hl�1�*\]蠆���7��
Y�'pop�ĸ��4����V�.j�\w�ޮ�Ӓ_�B����p�#\��һ�e��ؘ�ξ���>�w��Q�9��6�>}A�f�J�<�ҕ�V��5Qc=^�zW>�P���6 �ي�YM�8�u'����]���;gUA$�QW���-6g;�]��9�k�'�����|�,�~�������}�����#��,J� Q�|G����{��kΦ7DOD_�*0�D���g�f�OÍv��E��9��tt�їOT�������+Ew�ơB����=S����[9��S�\t�	h�3/�3A#z���U�>��=�n#��>��9�c���RP�+jj������3�*h�9O|��9t������<�<����̚����
O���,��4$�<��3��]�R���ަ�GN,�NȮᑿb"]����ոku�)�s�� 7k�����(!�<�	1�Z��X�G�;�v�b�7>rgN����}�5G���a.��e��{���c�w��z
�NǑf#�[Q��1j����ۉ+�P�ǝ�@Xʫ�`$$v�S}�<<T(�H�3tOA����r�.j�	�C����;���u��yyX��V�_�TB��IZ'�5�SX�׋1�ys��J�ygc�� �O"�]z7
������qcz����Ca�S�w��6s�>N�]��z8��q�4<jL��hY3��U}LW�D�����W�ٻ7跲�"���2�CyNx�n�`ٿ�=������=R�HOz���+��H��ԾN�y�֗5խ����;��2�x�cXL��+��ul#yT=(5�8᛼�Ѭ�K��įM�GK�t[�݅���Ҋ+�pt(������\C��~��|~~�^�������*@�F$}���@�����v��yV�y�_<5,~� ԯ�K)~��uU����F��j���*�yߵj��C5����DL&�_�ڞ��_޹�*�DC��0M"=?�K�Y�-z}����{5�ڮf|C�P©H�S��F�i�oځqa�W��뜒�d����v��8U/�{�]�ߦ��'�k�C�d!Y�㣉p�D�<�m�ǔ�20��ޜ�x7Լiz�wn�Z���q����� EmJ��a��ELw[��2'�h[6�a��6��\�z"
�t/�:	���ݑ�A�d��렂6�"�^u1�g]6kTF���F�L��W��w�B�7��c����zF
�1���P��c�m���Dn^����赏ޅ��;|�Zf٢��5�҅�h�É&"{�|k��h} ���d8�z�qc�a�θ�n��z��ݮ��<��S�3v�^>��X-����9`�Xp�?i �v:�����A��2����w���OHP����R��C�z[)�)�@����|p��H���+J&�^��d�e1'�`w�v����xD�y:���I���b�iU�ƺ}R4�G@��G֯,��ه�JD�֩�*R�JZG[��Q��т�I��[xMΕ�w;�nJ�)̳�,�T�:�srWU�z�u��H+w��x�c��O� �b"D@�}z"��R��ɩ�j�p?�?}C�⾐}�on�������݄Ma��w�7ܪx��-�]ݡ�z�<�g����t�%�r蟔bg�V��?�uDu/Z���1���x������Ӫ�ozg�.c�'!i��'~aH�'�Ԛg�,mez�u�	��\{�����E���
�-��X[#�P�¹�����Cת����R�4�c��)d�,�C2��J$Aʼ�w�Sت��z7i�?t��Qw�m?Pb�i_�Y;e��NI|j����l�LVh��]S�k�ۻ�q�����\�_`�P��Fjt�v���[��� ��Vx^��*�n���@��7�}�ݞ��LxI�1$J1Cʼ�g>۠�d(�X��v}z�8~~�L�ޱ���75�c�^;��9�ځ�^30i�q��Ԇ�}޿���u�`t�Nf�X��^�s��yHg�p깤1������n0�Ȑ�`�� ͎�HB���+z���s{���P۟{����.��>�ìB�����Nq�2πӱ"���P�p��B*��
���Ht�����oATZ2��̓/a��9	�5xo�#AW�]Cڒ�6
�S���<{�Yn)�(T�k)x-�����>��~�[ݲ�y��#��U�v�9n�	[5�;��m3RIc�$��m��B�f8��՗V\���JX�V���V�[8�-�g=H�F `@���s��c�c1�fͳ�3�����n��c��=eE�Di��7�x���a{�]��6��k_�����=�b��2$���;�7��8�F'*�Rz	 ��A����V7��w� PT�{w�`�^���*��c3��&�9�*�[��l?H�l�T#pb>�܌���{���#�P-� z~�K��W���d<�[�@���{��#�i�����U�B��,���Pf5��@.��!AxO#�bˊ����}Ր�	N�,����C&�c����ލ쮝_{�zgcv�!q�9�" ��H3�~�h�9�6��z�]���Ay/�/ҕ�w�y�̀՞b:~�8!bF�Ah�0���ĘU�D�@����A�8�}��;m�O�NǽX����}N����:�ߠLP�)$$!\��P����R{ ���F�U�)|D���w�����NB�V�x����^�+���P��5*H;�����Xf!i���&6���?Vy����������,�k��>���a�w���b���E�׬�;�g����w�k�Ŵ:��mq���P�
��m�Ü��Îl�gm�jyV�wigm��V���iJv�q����Zu�.!)VRZ�lM^B\��xC�������ّ�#'l]�u�W:����ڠ #=��6
��"���x{�����bS�f�Z���;�Y[���LvVBvTY�KX����\�#B���n�e�RnP�p"��X�{��sfp�%�b�tL�5�/����p�q��Y\{R�Zx��w�-�ؾ�F<9P���or4z�ci4��a�X� ȳs闒�3lM��᱙ne0]Ö4_x���.t�Y�m�*1*>���c����1��:f��h��sSQ1��U���` ZY��fL�`Űgeb8�0e�p�)�2�P���-н6&�I�!a5B�m��rY��� t'@"��:P�a��\iZ��<vR�F�5*���Fw�X���&L�{;;���J��MνR�Fѩ��a��ko�q�2���B����l�΅�[{1c��P��9���uy�E�㉙c6�]h��/w�E7t�Ծ�U��ڶ^[j8�_K��t_m�O�u�]���:N��$�l�����4D6��WV�ڎ�K�{{5�B��އ������Ú����)Új�a2�2y�ؗ$g,�&��P�����LvR!�T][be�y��������% �]S6�T��7l-�Y�q���ɵM^�'^��[xmu�//];P7J�n��e}���z��N� �-�Ɯ�y�;���u�h��?aL`Y��Am�[��4�Wn<r����ό���Bpt�2D�H��&̍�ǳUX�nNU��F��#����mk[���!�����g�M����@,)Xt��!���#��Kً��h�v�kbu7Æ	{I!L9f�x�ؠX�ͫk�X�/�@��m�S[:͜*\o_"h�i�z��^A,��P�	]&m��uxl^`���ŵ�}�8��9;W�r���Rǥ$E��;��!}�3`�ǐD� rŸ�Rj�����qQ�i�m���8%�7z�V�@wStK���p�\��]��O7�\''U��t�p�槅�=�hi�l74�Q%2�\r�]�z�{Y@��i⬁��JݵfV��F��d��43C���$;N�l�{�c��~����b��ku8���e�w׶t!�� 5 ��IW�bW���T�js��Y{�
P��1����Cn�ߋ�{�&F�p�ޣz��
�)d�4�P}2�.���I���v�s�:kf����h8�n�5
��;��P ΢��v�n�ѓ_ה��͍HA��l�;��uo-��"�dlM�[a��݌�qV1��
n�쎶!����뾰Z����$I=y���I�"�p��嘺��>�w:_v��B,&:27��\�J4�&��I:˽�4�e�ʱ;Yލ��k�S].ݾNJQՌ*G7,��r�M�����Xﾻ���Y�ӫg��`���N�I��AZ�h*�:6����JجǏ��ﶪZ�[��V�Q��o��C�ڍ	�Ӥ(h�	�C�������KF4le�(��['��A�k�T%kc!F������E#D|x�����&$8�ӈi14�v��tn��mT&�ح�EӋZ�N6������|��`زQI�;gZi��wV�(�E�i(Ť��%Dh4�(LZ5@TN�5E�tht)(5���1Vκ7[IGOA�Mڒ6GX��A��PسZm�u4X��^��i�ӡ-����M��w]�JC�ESĵK��q���Q�Jt�w��Z�K��:]j�LlDz�lh��(�Q;cN���4���*��Qu��HF3�ѥ�[clb+A�-�K�5�эm톒�D�?\n���~�?�)�������}�RT���v���V,i[����x���&�]6�7g�Ah���X��^��c�%U�W꿪�����  Z���#��O���u&G���59?W��y�B���B�vk�!�Jˀ�׵c;���n�!����w� n����,���d0�P��	�HH^�Bǩ�D?\���V3"�U�]��Ӛ�nAMF��7W)�q�3�>����E�c�¡T摈��R�?u�}UI�_S�V�B�C= ���(�x)�ed5B�T��}=�������dl����7����B��tY�Dfۈ���`-�P�L�K��g�L�)��w����|��}?���{����g�����b~����n����r)�Z�b�����<�������V��7��&*".b5��З�5"v`N0F��G���+jj����:ش<��7��Ó5��]������F���Q!��®LW�>�"��B�&!��v/��"�l�y�p~�N���Tb[�\�7ҡ{��ӷ_K���X��b6�فG@B9Se�x�]ކ�&E,�v]�~�h���3��P��v�W׸)M�XG���1�`G��(K�T��e��?E_���8�=9[ۮ��S��c]��
�ѨϮ���榚��h�=�G]o'��nL�̊A�}��7L]�H�Gx�����y���K_����u�S�5;��$:Z���y%� Uգ���u��|j���yfv�oiS5��K��� H F��>p|��^�u�"�|�	��m�!�IUp,$$v�S}
8aQ��f�����\�G�n��@S��A��=�gu��C���X�V�ZU�#��A�R軥�o\E��їv�w�n0D*�;�$��Dč='����]z7
��}#=��*��q���13J��g������!��u��(�Z��|��'�1 ��4p]�}}�Mdk�l�#Z��U�rX��G�]<pǗ��XIW���Y=# �_6L�
G�xKf����_«($��J^'��L�ѕ;�Az=\��;��a��"�����A�=�追��+�Dy�#(`��=l{r��VĪ��0�W�E��q�,C���m��U�n�@���+�}s�_�}��`�h��X+r���	��t�������c��������kJσn�<�23>��
}�T�p�*#_\�w	�~���G���)�+�B�ޣFr����h�p�}ƅ���)��#�_V��3E�c�W��>�0(o�Hc�
ع(2�+�4"������κl׷�עH�(�g,�~=����;^r�V`!K�[��h{}�����<$����@�����3Y�P���c̗*�^}�q�wɄt���={r7�׵����:�8I1m�/,�l���|�R�R���V�%*�p�oN�۩��r��F�&WtT�D��@� G��l$��o|	�1�s�B��Q����E(�`Fǃ{�	(Gq��6����Ū��"ߧ���E����<�*��i񘿆,��bt�X�`S2LD���� �6�Bd8�{�+_���ɝ�ǑM���F~����+�^��@��Щ}n�H #�Ł�3�@���甽g�Y�Q�'�����C��r.|6)PQ��B�|]?�����r���s�P��q�OO��H]��~�xw�����g�1!�C�Ϣ���U��B��Z��~M�Y��p51����pCW�C؎4(����`]��_ۂ`Au�P�g��:%��3�{=u�y�QC�֠X�4�X(�F<�Z��Ó��_�tNC���Y���	�&EP�>Dĳ����k��*a>���Kל�ޮ�]Q�k��5'!��Ϩ�/	�v:k��"3�H�bqB}�l슶�v��[��7�_w�g��c��(g��5ޔ���1`4�诲vˋ꜒��U��� Oh���h���߈�xe~P��U�Ϫ�W�������A�ZX����-��������Tܔ|�J����3x�񕛆[����g {����d��/rDl�t��c��*m�-�[�Y;f�o�Z��J�rj�k�Yf.�k��
����3�OB��OV��i�$�O���M��d̆u��(p��W�np ��W�>v'&�[]a�oz���0�D~�@���o˯��G�A��	�Q�OF	"Y�ν���t^LGO�[��<�8w�X�e�P���i�@�O;<7�8^Q~7�b���9�}�R���s���b�%Y]��A1;׏��c���3��㱸g��>&����!o��HB�r��o�|��eL�y��u�ݤ���cQN:nn��zGʖoNĊ
b=S.�}r�+�I��̷]�/3���s�Đ���J�H������v��c�O@�V`�dİ�#ї9�^��6Vp�I�*��u��T��,Zϖے/��h�;'*��'���-�w�B���\��N3�J�B��}J�׷V��J�E�/X���I�{��t7K�:#P�t�"�`���UkH,s�D��@���^�ښ�{�u��x%������R7f1��>���G����s������WQ�
�	�BäbyxI��d�w�OyVCϥ;p�6�����"/�(o�S��mx���}^-��h]��)� �D�H3�Z4���}���>�.W��{؏@�ۻ�����`�'�|]�^5<���s�)��a{�fx�[��w8kvn8#�	�#���ES^Z��s���천��f����e�}�C'K����%�^�����G6 ˗9l<71Ȯ�<�
$�1\CF�E�����F&r����������>��j��?�B������?J~�;���h��`�\d��ЉP(h>D%=��eu>I�۶�\%m�y%���)��B�m��R�6���r�/״��Ids�*��(N��~�����8�y,�99	�������B�E�u\EX��@V��0����Iͬe���������@�9�0�d���TTW���'��+*���y�^�|��v��;�^��W�
���n�~B�De��`��Y�Ǎ��(��Z4''��;�@oh���S���.a���$�c���5wl!WO\1�|et��t����F�,9��5 ��	�d!�q�J�"�a��z�	��1�,i��g�n�M[�'��{�9��'#��I�L�ȱu+5��=��z��^y�آ��ͥ��f�l�e�JMP��m[�r0W]tX>��������Y�����ygp�0y�d?��DzvP��m�*d�]n�>S6�S�4-���д�A�������_�����4O�
�v� �{Gmz-�f;�fҜg��	��m���=
�\t�8��{peB��\&fK�b��Ē1����0ђkE�}��rq�,�k#���}~��	$�b��x-�QI�
{���ǳ0ۘ�G�<�\A-�_�7������g*��]�s. ��1��u�2��JN����Y���@��@��;��M�f�߆�\�A�| N@U�;�~��|z�j;Gk���*h�c�*"��W���=�޳�c��,�l��#�)�bGO������q1��\Z�B�f��onAz�����ѷ���u$z<ԫ4����b=�g	��ف z�#BLih�򍂹W	ю�������+ڨZ��X�;�]_^�7�h���&:�X�"t�ž	^�4r'j�=�o��������Ĝ��a��;�yX�~�l����"-!#�#[<<TyB$W����]�s*����O}��8N��=��U�"�w�iߥHj�?r��8r��;�#�8��v�;Y���	�j�x�5�U�"t� �=_�yv��\��N��}�:���KԦ!�	#�z~��g�۞h8~�8��\+ҵS>U�I}��]�����ҷK�y��J6��،�'��f��n5�C�D(��!�j�����z@�,��nfr���*�߁��ۮ�I���+�ɏ��3�0�x���)A��l�-Hp������g�-�0�9��Y�_�c�ۍc}%�2�~��0P�{�b+U��Ol�	���A>�g��;���i�>J�Y�`��b`Ωo<�t�2�m�6-�=���۳�d�k�T����`�tܓ��y�e#�k[1ĺ�����{Z*�����&j9��|��ˮ���e�� � @����q��<���!�"�}S^1A�l8��R���b����/�dE�yj6�z/��/�߭��T�]v���/���*�2���b���pΕ�b�6|�i�gͻ��d\�+����z-M��}��v���K�S���^�� }�"�ԡ��Q�"����n�?d8N�D�]Yj�w��C����}ag���l�3��%�'�_IA���#al��/;��p|̥yg�W>�N�
jM1�Y��FGE=F���j��'��9�M	�B���W��b<�3yB�Za�T��H��R�]��b�Ŕ٬N�+��فA�&"{�|h�k��	�}-]s�~�d�SKs�4�ȍ�E�Ͳ�~��>.���v�_���g��`(�c�8A�4��7}���e����{�P{pÂQޮ�<vG��ǅ���C�zq�H�`�=�	�S9��^ы`�O�}�����)<�4��$2�n��m�M�HC�	LEzwc֎s�%l��Qt�w���=�G���@*L��H:�`���]D6_L��������FY�Ra�㉎�]~�G�6=(xܺ�-��j���ִ��90Pt�$
�&�v�K�l��Ki�IW��.��5bv���D��9B��}�5��;�������[/<�_�6�}�%ô�k�t�,�/^�.�0��s�/���2�Nb�	��4g��� G� }���Ɩ����C�1��F��
j�-�{�dkM,)Z'�Ԛg�/k+�WC�c�K�8),<�<}n ?l����	��E%�Vb��82���C���+Ɠ�J򠄛��=����~�؇F�M�2g���r�L?�E������A��}2vˋS�]����}�gq��d����'���� ���"�ޫÕs辟T�F�!���X�c�[��iznu�ݾy������b�K�>}7tOG��J��'�P�Cx69	v�P��1�V-�>��ʍ�s�y]�9ۧgV8~?�~�պ��A���"�������޿���u�},S����Q�x'.6�?F��k�ut�B�O��;�Y�>&h� 2�>B�w�B=F8W
��Y�<;�E���{���
j/�:n�۷�Nq�0%ϾӱA�`D��4�6"#y��>R$�h��t�������gZ&��l���t�~���;�=��S�TX$F�tz�/���=���(�͎�%�(4
��H�L-��m�"���c�=	�	�R��a�D>��ś=7������Z- s�V]m��p+����K1f�b��u|k�PN��vIL��^-�r��󃬴bޜ��-�R�������Oz�[)��j��d3u��9�v8�Et
1�f�����L�@	ٮ�-�� 	���CE������H� "A;�^�?��~���}�������L��BP��cn�����_�����ړc
�*�n�i:�\��f�������{��X�4l�9�H�;T��^�����\�(�|�~�|���1D-��Y-5�ԓ�b�A���%��o�pm���WF�����g����x����������7�r�����W%=�)GI�fʫ��eD+S�*
A�G ��-�����5dMg`z��ۉ)��JG��S� o�H�$k�/�Q��L*�d
�����S�Q��X_g���p��> �N��ϴ��J���~�1������.�GF�l���ȉIۍ�^wg]�=0t�1�������򸊱��j�~�ŵJH7*g���)j��B9o7���٣���aԩqP�.<'��+>������z���#�m1�4F+Y�Q�s���s������T����uʩ�k(T�W��|a�u7w��vV}�5�^2�y���ynl���J5��p��U��S���0�U�G~��e�#�<&�e}2k�N<1Lz����(yL�V]J�۔1��yIkނ�eq�;^0M���.d�����_GZ�wX2V�o����ߢLD+�ہh�����N��y����Ð��b_�+sz+�0�Π�t���{$��Ds7B���V�ͮW��+q�y���>#� ��mG:�i����!�R��PdX�5��yM[��=�迸�hYC�4,\�o3ҭ�i_m��v.���@�蠅�O���2���f�X����7��#>�_V�Dq�.�zg̪�������a�zʾ���_�FLG���Q
��LC��`>�Hj��/�3l��"��l����+<��#�x{(4_�Y��}@@��E'� �.;�P����Z8���aq��m�j�g��b�jsF�����c�4���P} �� /���(q�5�VMGw�l]M������p�Қ��֙az�Ói�q�ωJh���A�,l�����I�y_�n���Y�m����͢K�P�����;�qlT���R�M������{>��b6��!1�S3�zf�&P.s�ތ��q�QL-V1×��S��s亾��k�~��}�$�WL�d���C���¨C�,h��:=��s�О��m���U\HH��p �z�G�;+�/ûOub�Hc�`�._�=�Կ{t6@%b��[ʭ��!G  N���:`���U�����Vl��8CK6ro��h0�9�gQ�Sv!�_;V2E�͢�1��Խ�
���T��;4��.oV<=I���Rq�V�"Ղ-}K/�ܦV�)�<.�%�v:��2k��[�A}�@8oP-:!�q���5��cAt[�v�E�.�`Z�w�ɡO�=�wl�7hc�R��{ײ\�� �jQ�Î���[�齶_#f�r�)�+#T��l+*���N�r��1��Dw�c+�����A��,2�=���씅����ΐf�
nKk���k���K++\v5⥸�V�}%�!�����l�:�����BQ9LՃ5��5�;3�T��	ז:�fr�Ǘ S��q.�3�9B��n�7�����Y�_h,���3d�N��T�AV�Bͫl\,�����嵐���}KV��xR�F3�h��l�GxK'��
����u�ս�Q\��RJ�&���}�\�
{�m�����jQ���f�8�ax�a#ZD�D����+dlڬ��`P@y��>�=�N9���a�	���]�<e��hX�u���C��f��5����7��Q{��5���t�����Uu7�Jt���<���+�^9�̜��U�y`��{E"7n�m�˙�� f�D!Ϗm+cn���&���o����ra�N]���;�J�����9]9G�:��=]-n*0q��b´�t��}fkk:r�nn����r:���R$��� �M�˸ U;#F�e����Q'�[62IˢsgJT�8��r��W��5�V$��Wb�ɍ�,(�|��EdY�6.�[��Ζk��.����[}e�7ETRܳ��u��K'.�t5�t|� :&n���ԍ�Ɍw�����݌��Z�X�P݅f�.�%uk�ԛ<2胓ZU��<.k���͜��{�J�/�QyO�Zl�+S;S�#%�J�fU�Z�%e�ϰ�z<��m�� �N����P��PQ�h-��f˚���t�ӹ¶i���]��.����1��1�G�]����Vfs�+����.��(�$���0>x(��v-���((�AXjV5��fV��m��v�󫁪<����ZN�J�@H&���Y�Q��S7��ծy��e(��4޵�Y��(J��ퟁ-�uJO`���mX�y�U&���D<���8>���ș�:��1L�)]�����	�Dx��P2h4Z:�iVˇ���3��c�*̬��Aa3�tN�z��H��e������& �Sf=�5�}P_+t���G�ɝ�.u�Ӥ�7��w-�ڿpS+��¼�/�DK���f����Z�X�
v�k�sz�wЫז��˷KVf�lus"��d(��ՒG�\����6-�v+����u��2�}]ӵ*���"6�j.rS�OZ��(�fs�;Û����$�t�Ƙ�z�P]+N�����Z,���7�=���g�t[F���^��6��n·��.��:���(���?��||�4Q}�kE��V��M:��M1�J�Z1_F���j*+���d�?��WUI�Ռ��Tu�ŜCF���ich�ɵ�CZS@�?�A�N��ք���]���������LElV����C���������E:� ����}�u�EP֍��&�C�
և魵Gd��B��ٗI���Z4�ѥ]����
�&��F�4t��tZN��j;c��Gm�]t�ݍ4�h���h��M&�����j� tm��'I��v�:�F���Z���b�f�l�lU���=h)(�4����ƫlѷ뱢�ѫVM5M6�v�b�DZZ��]�4tT���k�Sr��p�P���]�(�Z�]���<bou���{q`0832��Բ�)��n��z�Ƣ��$t��\�x/��YD�	!g����J62CC�?�1 @� �������I�8N#zk�hQ2"bF���R�x:�[������۲���7Z_�%X�~�ԖB+��+-�`-�GIL���c63��e\�'�B�l@�7���d�禜r��Ǫ���bK4�@�p��+����bXoԄZj��g'k!ߤdk�	�����u�u��Z{����<����^�ݕ鼋�T��� ��0�\��m�����}�rW�H����TZ�u�{w=��4Mi�<c��qc�/����=89M���o wjŀ�+�2�\�_�Z�ۂ���v逸�����z>���#�_�x��_�q�}2᳊f�X۱����t���1[��.W���y���;ӑ2�����bv(	-�+jxC���a�3���v��Ϸ��O՘���S��xжo�+��:	���#>a��X���렆�dT:���M�b݌��5{����������6��4Z�68y�46����<hr$0C�@IB;����o��� {�k�{��K(��o�-gm�.��o�N*�Ƹ'J��l��d���I��
k����|9��e`�@�J|��#]D������k���.<L�+�� i���c���
d���*�x�.>�X򼫊Z�;�[̆��^E������1��bR�}�	���d����eMMʎ�RK.�9;o�G_��O���� � ����翁�*�Ѯ+�+��XU-#1'j���U��`PG,���G��dSP�1@�c,���HR��+����jv3�]?���l�n��S�V�U9�������Ģ��i�M>�eA�� ���#Y�~��jE�&� �k	�r��?f&/5M^�����ީ���#���P�B��
A�\gp�]D6^}�ROd��
�XkƪH^̽�_c�du��L����J��-��t���ē0�Uh�#BM3�������nbW����39J�c�qFzq�V7�$�!��}F)xNC��Xf��"��S��y�h}��q?ED��������p	�ޠ��W���Tņ����\_T�3�_j��J�"�����j~�~��l~�Qۣ(o
��$�F��ۘ�o'AiZX��?X��;ZA}ho�㉹q#��K�ur�'�@�=S�]�6n
ǣ�J��H�1^�^��n�:,���x���^��q��N#-{V��~�̱�,W/X���`x��r �}r)�!��w��"��u��6��g�7הlM���.���ʿ��5�zL��N��[��Nh�p�`����VG:�����CK��a�yǖm��s7{)�y.j5����(m!lH.8��)�7\�Gu�zon�;Xq��8�3¦p�~Y���E
����:r$���&�'宴�ӂfN�
�3\^7N��Zv3&=^�;�,�x�.6(�33N:��9NWwEݑ#��!�.�����%2�}�)�h����cn�N",ʔliؠ�G�<f6n�����[�JX��c�(F���b�M}ޛe��R�o�3p�=럣��*4#O����� ̘���8��cP�\�z+�bz�V�X�ܑw�'}&�����B}*OF��>�ck6�gɄb=���FD�4��� �@��`,N�X۫e�z�K�3��%s�UEs���1N5Er�c�_ڤ8���{��'`u@��A��uq� ��%����	�tq�����B�k5��z�r��9nz)��F�N@=� E� �^\�Ɏ.+jb;Ž��N'��Y_0v��<�����sy[���Wa����M��]s�N6
�����H3�^�����f�F\y[��9�xv�q���!:Ǖ6Vs�0o�L��H	M�KD�(��$®�&�ny���1��}:�@sV�gf�]l�K^J�*�ߠLj)�	�]f+�ta���1&�+5��؝����Ⱥ>��^Є��Gu{x,���mwz�7�����<_��y��[�+\7FM�z��g�/;�~->e�:��R��65#ʕ@m��˰��WQE�Y���~py���beZ7��"�9���:���r;d�� ��J"ߛO"�^���0VR�a�z�x:�`���ϔ�=��u��o��WzT�PC�W���=�P���پ���ѣ���s����
��+)pqH9ء>�YYw^/�z�/���Gn�g�ɯp���ע1Tq���*C���йe��g����(�� �'�nr~�ߣ�7�|�1��~�r�>���'���!�8Ul���O�r*̣���a��|<&�a�z;fy�{P���{$p���`t����4y�W5n3>��E�� �Vp�Q�~��7uq7v��hH�-��1������Pb��q��4�g�L�+P�M�qpw'c}U�*!.��Us�_.�������F�FE})�F��z��X��S��d3l��ƅ�}���y탗Q���V���#z}��>���	�bf���?p����Z+\�v)q�_�EtŻ�2,W-�{a��~9�Ƃf��hu��W�����;$��V��>8:�W�ɒc�d8%��t3�yϢ�㑰��N{��|H�
�C0��������H��<h�y]H���:��k�/]�o$����҆�&p2Oo���[���2��{.��Ҥ�[�m�Z�[N#X��:�L�>u���zkF�tG5o��ʳ�'y��EVʼ2�6J�EB��
Q����5���<�|ӥn)�7��	�LjV�NN�n�Y��W2H'�Um#��~������B�^����*��#3z�=����u�����p���b��`�s%���F�8�`�vLE�'��j���NX�;�>JW׹��:u����&;�!�~����r��chk����'��z5�u�i��+b)g��Up,$bGj�.��k��'��T�,n�Po��w�����?p��O��K�^ۡ��u��yyX��яE�4�s���3}��c'5�\?�Ҥ��C=f^Ȓt0Dƌ=5-��9ew������j��֧�Tn���`>�F�^�#������1�k�Bɑ�U1>�''!�}�4���I�һԽ��3�/?�M�,-���,C��������C�H�,��d���=+���+�v��O?#!�f�L܍O�^�ȱ�,3��-���Ȩx1�̓+���7'o���{�4TgM������"�h�A�G�D�1�u����|l�!���m��U�n�@�9��+CՋ���L��uz�$�@>��'��\�fT�b���p����G��L�(����83Պo̬3Nn�$�]�7���=FK��`�@�Ė�5��m���UolI�6���b	E<�x����BV+�aW�׽'��x�j�cٶd|�
�::=�o����]���F�]M���FQgNö�A\�,V��������
�vI�����q,�=}�X�;|jE�S�P/_��|�z��_�Q��iv�F4Fr"f=��E�������y�����}ƅ�m����6O���1�*t�%U�t8"O���ӗ7�.ߣz�琘O�\���3Y�J�/�##��z�[5�I�<k�D��O�UÎ���LMe�Y��b��f@{�L���X����_��Sf�'J�{f3$�w��>���sc������0=�pǪd(\z�qz�G�b���\F`\�@�}]
���Qt��z5oz��2H���8A�gs��h�4(:O�(���T�±]C�}ʅ����C�zp�#��uѪ�xpO�u�dL�����
q#��_)8�'�6z(H>e^�D=�������Z}K,�L^'��~�w)ꍶy�1&�?7u��t#�
�
&x)~�.�3�{>��Ce�l���k|�����#��V�[sH�)1�u*��NB���Q���2T4O��^��f��O�eׇ���Sۃɸk)B}�Č��`ޠ�6��W>���?t�����}T���`�ו~(X�ȾwՂS`~�$X�������0h�-�/����g�#�\㽠�f����� �(�c۳*��Z�(_v�3�f��z�ƃ�YU(���.l*kw5������%EA�W_V����Oa%�������
w�t%_kO��uhs���8"}2��7��wg�C=)Q}�AO���W�VN�q��(�I��
���~'d����xJ�#L��4��Ȯ���z,kt���v�)ջ;��އ��K8nc�Χ�?T�.�E�u�6�����¥E	"xǜ��T��B\nVw�ۣ��1'�v�t�E�v�E�UOݗR{����,�B�^P?Ɵ�"���� {L,��w��uF��y�F�'a?��ebt�8�-@v3'��7�|e�|L�#"C?6�3��}��W�(�nm�+��4q��81����z�
l���4X�P�6����Nq�2φ��Z�9��~��&d�Y��O�BX���m��މ
��ZiUJ�Ì�+���;	�����LB�Ewp8�i`}c��<���_�rŬ�m�"��N�M��q��	ʄEB�tY��TB�s�H��`qL�H=P'��8ؿ���u���
])�=��3 ��I�-����(LƧ����\�v��ͅ���;�O�Azz���\�(�r�̮.~�b�ÕՃH����ī��ͧj�(5�Cf�ȎԠ@ܭ�΃fW^e���[[sت�d0y�@�6���V�Z]�4+}Ǧ�b�������>N櫯]ֶGsk��/�-�l�sxU�x�[�s2�k�s�)�9�zoTĜ}#w����T<D�<���#Q(��T����G,�觗Qc� ���P(G�cK�f���vr����{��vm�J,o:�y*����,�9W���o���߫�P#��*�ƋL5��T�	�lv�C�.MY�q������:�\J�q��h�C�B�0|<�_^����s��\�x���y󤂿�|���N�����`�\E������bߺ8:�0x9��� ���R�z�Д79,�8��������ϒ�����R�/5k5O�{?mCb�{m~��2?[|��j��k��S
~��7w#�^��7,w� �U�j�k�_m�V]mF�05?���A��OO,����3��y}�.�I�=͇c3�_ҷ���9VU�,<���'#.֎�so}.��`�+��(d��,'�|�n^K�q�x4<-z�0o�^YW݌y�,`^�J_J�_w���L����Z�7ʔ!׉�*��dҲ��ˬ��Xg��MS�ö�<�&�m���Rt>�M9or���u͏e[�k�����5r����1����Y�\��Wn۶��Ė��-�����̣X�sQ���k�О}��dc]�L�y�w��&*>�"$����-h]�Ћ�2؏a�>@�������g�bq!u6�>F⾊�t��ӊ|�&�QK���־�M�^~O���0��fxl��l_��O}{;i՝��fs�,z��b�o g���uo�����_��(oV�>������z��[������۽�}�P���6}������G�0�]Hw��q��U���ܼ�w�p�Kg�>�Ξ��^�~�}�7I�?;��ہ��8u�..���{���86��!C[�h�$5�'��C|��I��Z��u{�)��7�_���Q�~t2x��Z��F���
<9`2�`A�}��Mu�z����@�/���S�{�$��!�3��z`��#��^(����:���4�q��&9I�ힾ�7�A��d�_b	�|g�Z��f��T0��-��Vz����Wth�MU�����<k��{�hw.�x�.�ӎ��j0#Lbcb!�{�jǪ%VA��&�/��<�>y��J�����JZݞ��+f��{�c��i�I}���"���U�� �ut�8�[�{M`�K�sq�#ZՐ��寎�"/t��-`V�f�L#��A���mMV��(�b��ȕ�+W��������+��3�4���c	��}_'�����v�<��~ɡ��zV����_h�O�2���||k5���Ap�������f9Y�^��u�D��f��+g����d�1����e���S��<�*i{�w,�yr��^] ��Ez#��m��x���ڳב�K�2��?nG	�{��|�˹�ʄL�zl���d���W��Wgq��7����c�1�����!�6"�r�S�!%��@{Է��-��q�M�����*��0Ǭ��u`�#'�3}�*l�ōY��K�w��no��.���}ޝB66D���P�؏^�5�	�6�j��ʲ���v'ƅ���~O��z1b�a\X����65
���5��uW:
�/|Wz������)��׻��/&�nzĸ���A��\�81Πr�m���r�d7�p��@�B��6���P��+:+uvRw%_����3�M(�����xN�cF�7n�y6:�.Q�׎"^nA��.�_:�0�M<ީ]����`}#�h/�'�5DDG&��u7.�M�L��}�"�]Mޙ�x�@N=�h9�d} �V�ַ� ��A�j`�@�;FQõzEEml�t�N�JN�b��G�$��Pĭ��q�Tu�ڸާx~���'�i�n�k����
:�\�3�f�⭷������w�vh�4ʻ��c�� x�ٶ,mnl{V��\9�[Mը������t�v@u����SV�k�Nҥ�D�ɛ�6.,���r��Wbg[FD.�'�pͣ�ˇv���:����:�|�lQ,���\[����g6�
(���a��b�畃��2��K5��5��"8�-���ػqu,AڨCFe���[���F���s%m��0���vlu�HU�^�'�/$*/��ܬ��u���K���	:�J���n��e(1܋�+8V��Px�r�ns�ʐ��N��G:�n�%��(�&��Gt�KC��}Q��3*r/:��ZW.�WKa��r7)���/̖��u;�'�n���� �jS�]^��/�"@���ֈ���XyG����Mlx��ۅ���dx���|�m�=�	��лW���48`�o������h���Sѡ\�Z�����X%��b���*�q-�rgs��^�w.WZ&��T�t���ܱR�]Y�x�O�k�ǫչlק�*��aFeCp��Po��Ӭ{��X@�ʺV!)d7C>���EMC���=�j�m.S�L��W����ܢ3v���!��՟ekri��K4�5G�P�q]RP��ݽ�+7��D�eN�WS;�5�D���� E�܎f�I6w#F�ݸ4i�#hΦ�.�O�+��`D1�8z�S�ox�Ә�׷���DPe^�`�AXҘtx,�7��-5J�7F�׽|��R�t�ԡ��c�G �U��n} Æ�nwc��k-a���-"�H�A���gu:��IZ�k˱��`̕ڊ;����=g���Ep�)����� ��j�n���~�܏M�o^N�o_ϟu�4�B�Ѻ|�D:k#��J%ݼ�O�Qa��t��I�UCRS��P�ΩiS�0���iV�7�#{N�n�U`T��X�[���h@cT0d�ݮ�Ac�w����d�]M��[�d�J,�:]	�Ҁ��^���;sH&�W\hRX�C��K�*�-)S�K��'ul���N�]J1� .B!��L��86<�D��v�e�8���6i��}�>#*���jK�Nb�X!�2gF'8Z&þ�f����ٖ6��
����`��C�r���eXE=�݆�=j���;�Ã��囨��@�}n�ťɼ��ܝ4��\�t����`V�j�tm��[G[���f��]�ҝ��WC�4���Z-�g�G����QSW�tm�&���F�#m�$�k7��t�qO]j
J48�5�1��������|Z�t�4�V�2Dm�[l֋X(��j�N��Tv�ZM[v5�Lq��������b*��DlkFm��%m�CZ�+Uݒ��1iѧF0e��{�tc�������kA@SL��}��I�j��Z5E�mQ���i����SM	�z�t:4DL��Mcj�k�Z]Q��wS���ֻ`"��6�m�jŤ��5Z��z�v����t�ѪMa��UQ��Pͭ0mTb��ӳ��1<l4v�SA�������*6��t[QZ�Uj��kg8ƚ"ڌƴ4L�j�f)��:)�3��U���v�E=�ݱv6�U���A�kF��=�ڈ��Tlqv�Q�q4V ���.��qm���ۢ�*��h��wn�
ر�P���t��M^�0����.]��޵�k5:H�;�!MU1{Ф���;l(�:�H�W[��'	�}z{��D������LDN�����wP�b:F�:�oH#�W�?V�.�{��'�:��?C�L�������u���k�k)���H3��}|��t��..�:�p�,38�J�p��T�}�;1�w�����t���4GW�Z����٫�&��6g����{���9�H^��O&�-{uG
�r�,c�æps��f����w4g�؅����gs��-F���~����'M��@�������R�5��''+�6���8�{@���gzֹ!�ռ�|�ʤm�ʲ�mAa���'��=�w��q��u�����{}��;;^��5N��]�������ae��HzĶ+d�Ή�/2;���3懻��
Pzi��w-;�w2��at/ ����S��Vl]�^�>K�b�шnG	�N���������$�m�FYy���u���+����o��ە�F;9�ϒ�a��	�����-�ӝe��)�X�Ԥ�f��	��$�����ק�.�?�nV%�B�R{���OVD�S�,8)�\Ë9��:�u�]���T���1��q4Hn�`�zf��wӃJK�"��J������=����Wփ���Zq;��q�s��D�~Ӿ"���3��woD��P�&�=%���5-�V�����ֵ���Ϊ��To1o�e���z��[b�Α܀xoV�'ObW�k��{�0�{j��r�)�C����Rݠ��|��@!؍ﷰ�Pڭw����J9{��m�`������c����WW�=�t=��{���xM|�.'�k;ͭ��U���Y����U��P������,��k�/����ޱ糋�dv�]�==�F���xc�b��)~�~���6�ԅ�Qޠ���C�g�O��� O�}�u��#����{�x�k<�w��)���A�5�X����Pۊ4���M�½��fC��0PS?1�7�������=�N���c7���B�{1�pm�/�[��*��2n3%w��)^�������\2t�������I�o��ɬTޒ�[�� �R�	Q��0��f��x��ڗ�9˻h=y���PfLt��{�˛sR�Q?���yF���\-�t�2V�EJ�;��!+�����&t�3��Q/�Jfv�ۉaq��ISvC�sfM�:Dn�F���V�� �zB�����:��4��}����uA�aD�j�Sv}=�sG�.�����O-�:�+�N�so���+���迂�{&����u�l��T��z��c��B^T�ZǆK��ia@|��Ԣ�m?�{��>��툎Z���	��X�D��b�Z{�������Վ2��v�gL�u�c�v棛p����_X���yekϤ>�-�@;!X����Sn)��OA��(�F�}����Ŧ�}����U� h�t�z�3�2�C�R_u��p�ܗ�z=���J�<��>�ާC�:Da�z�9V����(�ܵn ��>�����T/���m���u>�`��cձ�kMDc��ƾ���<�-�����j��m���NC���
F�KǺ���������ǽ$ju=��*z
O�C���.�+����1�s2|d�\+��w{N#�J,}��¸���x��7J^g?g���7�A�(����]֣�(�1�<�|�Y��x+an�;w/R�&��h�W��7����^��V^r�g�;*��1l�n
{�zx�;Ҧ�FF@�7]9�xU���ҩ˺)�ou�Vǁ��Oxw��Ձ��b_�<<!��v6���9mMX��őp�K��8�clE�]k��]?W�j�d��XU�Yw�2���:�zX��}�bs���.��t��uˌ���x���q���T��уW�VL�Uu���g�����P�+��ß�񲽿@�׿hb�f����Ѽ��*�]U�����������
��Y���'���C�����nny�0���cvM�;�;n}7C[~�;�*�ӧm��������/�<iRَ\���ML�1����xd�	���o�S�A��[�����ٳ=�+�/y3ޤ���3?n���:2�����ؤ	l`��"��X6O��ٻ�{ݙ�t�ZI�:�&��]��מּ�b�b
\������{���q�߽��
��l ��=�R+>����/~�#״"�{�����v�p�l ?Vq[�)V�qf0K̲o��wO��	u`3�gq M���*����nJR�C@B=Ĩ{�g����6���hs�K�u�J�+/T�u���	(�5@.ݡ{�)��K�Bk�b�#�u:��F�;�e,���wj��3��EIZ���O�1m!��t�/37����L>=GV�z���>~�]3w"9yb9�_9P�j����y��O�V���O@��f���GZ���[�U~���6��&z���7j�b�����)��_E��3�ī������������~o��_�n�o�S�Kq���F^�F�7;ܱ.�/���u�H�|4w��'�#ξ^��2�*����.�R�	�+͎S���o&�C�#�ޝ�V����
�i�fW�na1[7�[����(m�xz�k\�
������
����1g���
�¶A��c՞kp��9�\m��/
5܎���[��"�z���y�(b�o�����7}@�/z������K����ZڼTZ���̗͋b���fv`�n3%g�S�~�Y��~������Mn��o|����K4ʹ&L5��k�43��R�EX	f"�j��.���'T�O�xC��'Y�k^Z�z5��O���d�Swñ˻�&H� �ͮ*�;��&�0�.�Y��Ŧe�wn���'Ke��lT�`mC2��˔x���VNf��|���G�����[@5@���[����#��絛(p�rZ��cy�x�;�(��ueP��X�/�_}Ӹ9A�쿶��z��ׯEk��殱e�CT���n������p�U�^Ӽ���^�E�^���b���bQ:����[���!KOg��o�{8�귙�My�OvNn��2��1���� Zq?v�O>�m<i�ò ����]�}�5	��!#۞�q��!���[�����[�w�OK��D�����������\�7ܝ>_�����H�3�{�)��wOϛ�뉍�g��w�)F=�P�ϻ�>ۡ��6�̡_�Z�}�B�+���M{���#�z�����i]_U#+��gk~����h>�w��{���EsS���u��=���q򞯖؞�N�[�Fs5v�;���`<v�� ���D�Q�w���#�FM"<A�7��V���Ұ���1Kwk���v�ϝ���z�&��m�e�ڟG{Ia�ΎC.Ն�z1���Q�.��X��R��F{���'� �(�#��S�ʷ׆���<|77x�!�#zA��C�o�m��X�ԯ�w�)�j���6��W��f%��T�ǵe�>0tk� ���O���n�}ӽ��{����0r�0��#i���G�-颳� X��6�ur�G��r?���0�{�tP�S�=����`n�Z<����4^z��
g���s1����=�B�}��w�}_5��S�䘮�9+kBk�^�u�~ڃaf�۵�� q��T��2=���c��~���?09��[�In5ٗ4Q�Swں��yHqյ��4P�V%�O1:��Y/vOySVt�_T����g�ؿa6��[��X��}yH��RCN���?~��{[/z;\ש��Zp���:]~�c;�w'�ˡ��!�݈��B�s���N�������{�����o��{|�JƚT����T>�xΌ!�2Jhm`�� �r��d㾪��<N�|����8*�%3GK�Ӿ��v��J��1��ܣk�:���Y]�=K��5�m�f	n��)����˩d�3b�����̩Pd���T;)eæ�d�s2��=V�P*Ph�]����\��V ] �3����{�U��V�#����3퟽�6�?o���b~�|�N�tw��ߎd�����+�~���w�%��[c�)X�HqW�O�snW���>}�&��;��*,��.8�����o��_�h�m��s�����{�������6���}nȝ�L�؇�o#˪��@��G�����b���O���.�������"=�}�s7��������o����W��r����*�.�+���7���+{��	�R�U�X�zb�����o�m���^�(�{B'c2�S�~�`���Ot��BiGZ-P��U	�,3��w��fb%�͊���U���Ֆ���I���>�]+8��?v��VZ��=Z#�	��w�u!p����F��pʓ���.��筅�/0�7�P	��9HH7�U�ھ�#1靘c��a<9u�8�D�n��߬p�
�:q�F#k!zX��G�=���x�]�f�
�2���)7y��t��2.��Z������L하#3>E��DT��۽W���p���N����9�;=
�����6j�s���doMmi���Թvb�:�u��ʱb1|;E�,�;����U�Wг�?\���̄��TB����}B9�T�w��[��H�W�{�\�/{շղ��W�Vg�W��>r��.���6r�����s�r1Yڇ�z�j�m�r���o���z~�� �3�}٫;Y��]��y�>���8H��ݔ�qm<i�o�G�hE�U�}�T��**c�47�5k�6�U�t�y��o�.�������x�3�q^��Eu�^V���<�1�'ޣ��}��b���7V����~�ܸI�O^�]F̪[e�ר#wP�`<�zD�z5�ze>��1w��s�:�W,^�_���>�{ҫ����c} ����P|D���ݪ�9W�L(}�;Q}�߳���X	w[�����ۘ�u/=O�t� _l��㘯0Zƺ�E3`��ܛ��ڿ�>������ڲ���t�|���z�v�C\2�&s�w�d��[�!J���F��u�ל�|2���wU��Ӻ���;�q�4��b�P���m�gd�(gm݁��rYٵ!ˏ&M�LØ��;�Z�����ۜ��]B_i�;���,�{Ҥ�(���P<BC%��d�T���N�)�5�� �7_o����)��#_𾯵aU�-�3N�T���^s���P���.FFz��`���>�H&��>��B�&��Y��/w����a��1���C��϶�/�n�<��v.�L�D���nZ�22�����fF��w0�]�#���_�"���s�5��W�T�o��=��n�{q�g��ʲ�j~�Ԟ���&�VAk;Ϯg+�풻�/^�݌j��}��\�Y��l/r�������n�?U�Kf1)���W��qv!��//�v����V�6�w�`�9
��ʵ���!a��C��Ju�M�*ަ���-=��I�"#0��6����5�b�|��.~/Z��^z"-8픛�m>�����t��F�:�w��Cܺ�s�}7�`��	���ܤ�Ͼ���f��e`9[���@����31��qli˨�U��rV1�9s`��:�V)p�ctJ�<��u���v�L�-�o���[ӆ��ebJ���L2�;Oۗ������y[Ͷ��Cs��YW�8�	���B�=���[��Jɔ�.�R�멂�Q�ɧQ�H.����ܱQ&���Z��bl�H�{�V^ǘ��Tr���p�3but��_�%
P�ٻӻz��f�L@�ѡ:-�M@�#9�����]A����4���*�Y"��Uc��B��nK1����m���Z�<:R���ȥ�6.,b��k�6�G�jn�Θ�2sLh3���u��Q�L�-�{����>޶�#fn���
���-�.Ӓ��I]�kb�sH��Jѹ�h�y�riǔ6(���`����5\k��]�S딃X�)���Mo\�����w������y�T�x�(����ko8�X�@��#1�Cʕ�+d��Z�z���Z��qs4s�;%q9v�.R܅�}����iT����\�#�и2�N�PZfF!܉po���3�V�m��\ِ����:&��f��F=5έp{�V��q�A����9����y����J�W�닧�Ox�)f��6ĵ�nj�A�:�sVa�t����I���:q���י{"9Ӷ���E�zofg.���՛�N�h��A�̪�U����r�|j�<mt��n���s��FWn���ͬ��0N�<	����Lf
̚9�oI�`%��FH'��}�g�7���<Ku�yL�t��ЮTn�i�cp�$u�E�ݘ�#дձ��{}%>��vc��E��Φ�q��W/�Ēy[%!�\P;�  �4Ja�Yv�f@�M��`�^�v��v7d��KM7�z��E���V@�p����n�q\3;�s���yn����!���jul!3IӀ��7jPi��jd�3q��5s��:OqmJB�_�I�Ŵ�"��Pd�N�>{Ql.s��p��8VJT�q�@���Z^]i�w>��]v>sNک�bÑ�sWY�@\��\�sқ�&T�V�L���H�W^^�r�#�mYs2�j�^�cCy�6�f���,�����h��g^;h���Ρ*�c�	)0�hΫ<]=���.JPk�뾤-��ٌ�6�6z��J�	�!���hq���	�"6/����AH�^�gi��@f��7�x����V�1��d��2��v��VL-�}�`�ʭ'�]M�u�e�x�F����r�����fql�ǝ��Z��W��ý�n�Q:!9w�It���v�uS5X.�#�1���<��E�p�Le��G��3&9m��l�N,'-_VJaX����|�PpR�.��(�΁��Yuw\{S�S�d�t�)�N�wM�Y���&+9W�|��s���My����\{Νn�l�}�N��$ՅJհ�	q��]��=������?��}�l`6�#i��j
�h�E�OZ)h�UZ{��k��DSZwc�����+�裂4Q��PTT�Z��wQ�K���Z����{jv�l{����,cM8�������A_����룢��.ڠ�����S���m6Ɋ�k�k�㏏���}�Wc���[QUl�c�M����QQ�����30�bݷm����.�i7f�8������5_N61%�AE�#Z5fْ�c����
�&";kV���Q�z���hѦ�llgj���A�ƶ�ڌ[i����WY;[���K�"(�DGZ��n��SFb�ڍF���s'A���SAu��T]�ው�3;w���Z�k�6�b5��펌Z�Q�=�ݺ�� ("+F�4�z
�m�Tn�:Ll�m�Fƶ1��Ŏ����U8���4길�.�.��hv�h�v��vh��n��&�hڱ�������	4���
 ��So�͏[�n��L�d�k ��M��{�m��]t����jUέ���>raj����*���;b%#ȳ8��N�XYgl��a���4/%hx^��0]X ��t������m����7����a�@>G������@�0��P�w��|3�I5«���u�kO�?_6�<ӽ�%��\;��cz`ov�YU9)��c7���,^�ٞ�=J�u��ol��˦�W7��??�g�>���稺�d��4����Ϥv��j�Oj;�,o:���z���Qk5#���)@�x�㮯�/����W���W;�����k�B�I�c�nO��:�{��-�o��N췜1P�F�'�;��/��7{�g;���jy��������t�i�𷦏`��`�b��6�οnf\�#��#=��.�R���R��Cw�O��2/��fʯE0t��9��VN
>��1;WC{���(���hӺ�i���݆5r�o��=O�˯��	�iK����t����������~9��_���S��?h���ʠ��S�[��{?~�㍄��|tU�t!���yA�����Iٻ�����ƙ����G��N�ʱj��e�B�Υ:|��v�Kț�:v�/UN;�`Z��'�4 \O;�����,I�pT�����b�s�z��w5]���,ܾ��U����d��.�ڟG�kE*$�p82���ܼ�3^��{@ia;���w�������+����̏+�Փk=�_{燫�Ȑ�!X��o����8�mB����>�ж���T�!���s�b�N�����՟HC$�<tp~�3*�U>Z��*��|;��t/�Է�/��T��]�c�:2�a�����C�f��d�;��b깟h�:{s���nl���vC�}��%
~��NT{-{s�Y��-�O#A��_�����:�������}���D1Ǝ��oTk("	���E	�m��.y�Z�*ZR��o��ޜ���إ\ˊ�����������͌{p��h��@oI���o��)>�z��cz*�x��������fv���ݶ+�b:G}�H=�������=�t�;���jW����Z�Ӵ�!ڑ����B��`���u��q7~�\p��N�6�2�L��p#���V�h+�ˍ�?cbn��Υp)f�W��CY�R'!7Q�q��e��љ�K��Ǘ�ӾWQKܧó���4km�}.���݆:�&k0n��i�'v.�'�`Ǡ��]qkp^��q��n�v�L�t��
F,T5O�S�.:+�b�q��^��R�n0Ƅ��u��{_Q���+W3�f��=G7�B~]�y���PN�M�>�zbw-����L�C�3;��V��n��wϛ��m�>�;4�V���d%��y�~X𭘼�w��r<�'g(}ͿmE���ҷҞ�-�[m��vV���7����d��wJ$��q�V��Cq��&ͱ[�y���Zw�:����W�v��ê��������:l��(w�Ge�;ݑ?g�!��-5�#-Xm�+�����}��{�A�ty�q���sn�����z��w������z��;���m7Ɲ7ʣ״"�U�o,F:>���^ל=V#�X��^�Huw�5�w��n��|�iA���U�ڜ����qG;�D��/�Y�z��A��j�����Zz_?{��n#LsD��`r�P��S#z)d�c*�0Gu��h޼����ԓ7:�3�+K���m��,Z6_2�0J��c)�ⴿzt��C�o�Uo1��4>��/c�;��WN�[:�:+/p2⭻�<��H椷	�bc9�B�+9Tx�rU����}�p�z=b��K���k�X�vT��0cf��dz��kz"���^�sb����P,o�!�p4����k�K�ޅ1w�Y��-��΋�]ڼ�u4�K��79�:�=N2%_�XT�]�B��+-V����=kdwP�֬y6�C��]9Czv�V%b�e��U-�^���"���DS�����������ܩ
�����}���d�,��\��vx��7���ē��F��2�X�g���Ӟ8�F�B�m��*����X�q6���Sy0���%XࠦC�nŇ����lL��}����s��`�~T߃R�on����w8ͧ��fvb�u�ܜ�W5=/S�5]#8Ϲdz{���>�C˟r�;���[ɢ�mE	p�s2J�͸ߺj���^w����'kש�x�;�as(]YTz �����̄&�L�Vp_.wR�8#\�J���l��<*�P���)�}-�J8n�^��o��أ��ħXf��d��D�73�����6+���z�C+�wy�k�5-�o)��V�wg��ה�2`��@qZ4B�p��}pS��H�4GGlI��m\;Ҭ:��9LU�`Y��U:T: ��|����qa֩}a$݉i��w0B˟-�^��y���_mć�7��-��'��U�M��-X{�|=���h�2�5+���=W6���z�e�Cc������@��{i'��=>���Գݽ��'��0|j&�G�ۍ���}���ܪZ\A̝y��Q���]37�>�ҹ_k��ThRZ��=�3�@{6״�bg��+9w���u	�5�YZ94j߸�庱���F��������%O�_(ܯ-@ȈlKT�^OS�{�����)�utʩ^�wY�ǲ�T�s�؟|�����u���P�u�)��+��u��<�c���T��a����>�<2�rpPPXj@;��CC��؛���-�RG1�U�w������7����7F:��F�Hu��7F���7n��#:�A�V�|�䳑�}���SU�;����h:����޹��cI9%N�Q�_{����{���/W޾�Z��*6E�cOb1n��L˲�����Ln])2���v�<8Z��M�r��g�o���gMi�;�?A)�����g6�NnD�mnm_gt���������i��xZ��=C��	b�~<�v���@9S��b]Y���ʮ�7�����ӆ����~�����A��LLeM_��)ƭ�8#<����t�gO�rb�c��Кد���eÍ�����ܮ9{���=�P���2��~nǪv�ro��^	n5���ՏՓ��(�����c����*�G�:�ļ��pׯ�/vO@�Myz3�k��s9�./���Y��Ֆ�z����ׅP�~��e�i��G	�}�����Ȫ�{\��ޭ>��a�5���V��:�vYt7B����=<�hWdLִ�UW�,h��7��Ɵ�%���/��3�ф0�eW�^e:����~���ы�=]�޶�R��>gg���5%�39���,e{�E_~�x`傲~(kٗ����������ܧ���`��nǡ�lO��;���:q�X5[����[��_�Lcd;Am6#F���k\9N�q�Y:�c���ǣ�	��%�EڛaV C�D��+���N�F>���0�c��:ו&�>�XC{��q�}�'P��[9^�va�ՙ�F��0m�/�w�s�'�;��G�F��.X6�]�+VR��o����XLRV���N�*�������Y{���l�7�6�Ow�|���'޻�]^�L��=�8nw��I݉}�X���GH�o������S�sr���{��~:����v������]쮱
z`��#���d��=��7���s��D�����z_�dwӋSp�\����o�6��<2}�4����:�_t@�W0e-7x�}�S��'z��7bB�3�?c���4���Db�id^O�!b7ê�[����Uyv=��z�K�`|��+إ��,:cE̟�=J=�^��1��ĤE����]�}7����sٵ����D{�!WV)g:���z(�74W�`a��?5��t��8��q~���8W����=�ޠ���Jy��͚=W0�~r�D�T�DncNv���{���)]`���|�L�(�Xm�8wqz�y���A��sw���RzwF�j��(�/*�<H(�ԥN��μƩ&09g2Y�u�Ghh0]۔�;�
�'&g�;�9j����|���b�	9T���d��Jp������Z��[Re��	mSn�\�=o�}��{�q���]�tg�3�o�Z5��� �w���S�-,��}�7�z����Nx�������������(J}C�_/u;��@���u>Y��^����U�mK;�	����^��87� �}C���]c���'�<��;�#�����Ϯ��U��فc��H����6�2�\����V��]�-������6}�����ޘ`'Ӿ�|�����ot�N\����Oկ_�%�n_k�C�;dER�"�Z��~'�~���K��
'�@�C���[���V!�e��:�S�{��<�72�-ݰf3ӹ���A<��f��H��{�$���*B�GE^�߁��_9K��iGx�~��:��g�+LXA��eڱ�C�߾H)�c�O�>�{o��3 �!�6r�h����G�Y���� ̸h�ېVE3�Qa�/����Lm��T���:����"�)wk���1)��6�N��FJ}.1�k�gI�fgu�A�q���5��S����y�}�4�%�aMQ�����Z��̗��V�m�:�]_�_��~�n�F�*�t�c[y����n�Z1}p7���c�U}=����[X��q�6�7�Q��)��99��ǖ���.+|pw]���ϫ�������o�"��[��*���c9��N]}~��ڹ<���=����b�w����؛��u+We��.��3P&kUA�����q��"���]?\�;8j�$t:�T���&��v��7/||L�/�u��%чm�P������%��/y{z�x���'����؝�ǹ�]�R�-vgP���l�e|4���t1�"ӌ�SF�	��&wk�j�L��@���7��:~ݡ۝P�d@���}����ӻ	��~�+�	�I��0~��_�{�K������3��q�ߵ��(�{!�r�ī=K2 ��xR�Ĺ��_������p��_��*"���"��|/ �No�W�o;���AAJ�-ei��k�jh�HvR�,�,b���CH�컹+.2�+JT��d@�Ҙ�h���Ս�o{��˕"}��i.@Ҡ�;������%�q��M�,[�� �a��[j���;�3j�楄�Iuy;���������W�� ڭv'�P=ַ�_�HN{�x�s-m>�#���tF	��7�y��������7�n>Ot�,�7�{.s�11��Q~��Y3�8��H����O ݞ���o�ѵ��t���m]��E����xҘ�ww��x�F*b`��t���/�y�|��u]��k(\^经,��0Gzu�I�A ���dw��6g��0K¢lh��y�z�z߳_V+}���>�K�~a�}~�����,�\`�Q��x'�
�Z�H"��hEߑ�=����خ�:��_ɭ�����"�x�Xh�I��6:�v}��s)Xw���º��y���r��k�UN���TFV��Cד-��yU��b�X�ʕ�~ׯ�|4��mS�*�"�/�t��}�-t�����7������$"�B~i�����^��DA��7i�W�Q�V��%or��m>�Ʋ��B�]S��OZ��-ʽ��Vk ���)U���dh>���͵+��āF��N��L�����h��"+ظ�	�b�9VGWA�[x�����&�>sB�/Ms¸B���E"��kWؤZzv[g��E�)#|���Ӄv
hsF�����BE��.	�W]w;�����Z��:���2ʹ���1Yֶs޺�a�}>*G�Ŋ��^�M���8�O1�I��G��n��\5T����O 4C�ɉR�lx�
�N������t]w|��V���ͻJ��*S�c보�g9��U;���r�<��C��l�ez�0�� ~3oyi(v�[�P��,b(nܫ"�»{�t��b����Y+9�z0��g��3�	d�����bh�A�F�q�i�v��0VAadcE�t�W���7�jޜ�v�[�E�**c��/L�vdGpEXqXV�Nw���ۚ��\�\7���'R�L��V�����&U��ta�,F����jV�w�lT%;�M�����u�:�;ӻf������n�b��aӤ_E\�MU����st��%��y%�oz��f��Fc�B^(Y�<�,ȚMZ�v�7�n�ڨ��룤9�W����w��)�o����e�Y	����F�S4�qa��/j����VaWt����[E�ɾ�BXF�=͌�[^�ZJ�5+\0m�l�sk���lL�@��\�Mn�bv;Vd���X��WR������8�_	0�u��,ф���+��V���s/���wWYHP����>�[BJu����/Tֹ�V���U�GFN�"'�-6��Jth�s�p<9��N�����F;���k�e�훮�*�18s�"V�KCU��S<c��D� #I��yt�6.�DE���WI��knr,S��D���sS�K ��x�#�7jܛ}��zud�����hN���x�@�� YJv�"�)�U}9�5�'K�<y�䇴��+qZ��r�(
Pk7h���Yӭ;����`�P�M(T7PT�"Ȫ
��n ��=Q-�O	-����mo&��,��s�[�V�b$���D�@����+��!�olʈ�ne��;f:#�C���g0;�]u���f�y�P�� ���Es�o13��k�F�R��w��&�4.o[D��p.�6X�uy6��P���San���1��ra���i�(���uNa�<$.��-u�v�b�t�rU��gAS�� ȳ��wf#ǭ�s+%���pޅ	ut�͠�^��1\���m���#�T���p��R��#���W^�G�*S�a�,m��y:e�À�Ĉ*��k�<��ո����Wl'ݏu�+I[Yp_��X˽��j��_o0� R���a��;�B��s�u�Cn`ށ���-�����+�����h��*��c:5�6�q�\���j�m]&9�vu�~�������$֊&")�-��:��b�=!�:�*64�;f��rc��������_F���Qۮ���h�5�E���
Ӥ���b����F>>>>~�$���q3ET�E����*����@ELM]d�m�1Ӡ�(�||||���;��0Lm��7cwq�It�)�t�Q4j--SӪX�Qn��t�t��WFw\�F�UT��tu�{5�w��4�Ez��k�{�GZi�����몪;j����x��Ʀ^�bj6�G�P۱�lEZ׻t�4MTQS�L�aւ�Fwq���
l��5�D�8툮�TQ]�ZLִ�C�**��Xb(
i���Ѭ�i1�1��h�5����L�Ub(�3SFՌlzL[h���E5Wb���(}U���G�pŏuSpA���眫��|eԴ3�;)�u�["tMv���q/���(ݽ�t�E�7�v1�7��y>Zk�Jr]��?�!�4q���j�m;���]D	d��!.�yu���s'�5v�ᜢGu6�,>K�4�k��w������'��d�܉켰f�mo�=��	�/գ��.��f��:��y�;/�}ޗ~�¤�!>��J�qѨ@��=�<5�ڧ��VW_y�x��ܧ���c')H�������i��cL��=�t�_*U��	]{Z�~'�7ٱ����>�{ҫ�v�`��� ��@�,p�PD�`Ow�|��ɮ��Z���}��)��o�W�&�һ�P�u�便���������Y|�<��̓�v�C\�e�7�%<��P��t���M)b�Y1�$U�}��H�F�M'�ç|�T𯻆���W�呗w��D�F�v�i��yݜ3avu�\�l�rϽ���Bho.B~]�]3��<|c���{l�œ�:b�_�#Ψ7w�x@��᳨�}�R�t�u->Hym�ۂ��]�oЂIɻ`r��,��$�t�ɫ�/tL�=X�N�U�hc�ҷwF��p��I���z�-�szI�(ё��\���<��1��](�.�Z����N���ũ9�]U���4=l+^aԓ�
�Z�==8������B�'��n�/�7������V.>5�|qׅw=�I*�\��gu��n��
ӗ�7ޅׂ抯(,<��T�O!��5�n��=ן��fs���IP�~�MZ�J}����7W0��i��~M�����g7�lY�s��ջ���a��r��{���}Q�30)��}��W��7��JC6P�עEj��a#���4�^��ę�r'TFPC���4se��h�S��k�
�[t�8߯��]L�Y��,W1�+��W�t���}�]����@�}_u5A{+����k}����`�Q{c����c�o�P�V9wyt=�@��� q�@��g^�	�L&ϳ3*�F�h��1�P�{{弲�r�cr���K/h�o�7�@���^���A������^�T�;�um�]�̧�׭�<k�ѫkqW/N{;6�=}�b����mȱ�;E{���,��j�9��`i�7�o �a�ո����'K7�"`�7Z혅ٮ�z@�����p�[z]�6��9��4%\f�_�g�*.�u5e�QQ�]�M��V���~������m}� o��eًW�|E�u��xPp�S�;�$,�c�~M�C���(����]q�Ȥ���V�`�س�JoDj�XQ����;��xzE��r�(Q؟��f)�Ύ7� ��WU��L�lJ��_W�x|L`b�ъ~2�_�<�}�:F{�3>N"��aR�+�٨uF]�Yυ}ˢ����O^���>6�m^_o�Պ��{����>���QC7|&�������m��;0lw0�s9t�~W�C��fwfYy�2|�g+�7�Xk�x�'�3��*ʡ��+��*8A�x��*�P� �(-�y'õ��۱�S�}�����̯l`�Y� dUx��Ggzt=�lO�5�ĺ�R��I�ۿ��9��cW5k���TnU�Khz�[�={ʷ���7BI�2n[��7s���ϕ�I�s���7
�8�@舸b�ۥ>l�zhR˲RJ�vw��jd�_`�մ�Ьzf:�c��1��.��1��B��5���'�]��waܦ�F�o^:- ��s�2M�n�����N�t�����+��w�ux46��Wt^c����NMt�kZ��P�~��gWі��l���[���۩2j(����(��F�_�k�9[O�[�{��Ρ
7��'��3�x�6��צ�2�/gw�7V�j�+^�i�ޥ��M|����5FB��3���Z�A�D]������"y|ht�L�;o��R�5o�yn�X������1C���o�ǽ�w��z4u(���U����@�Z����i]]8�}�'�!z�Ԇe�͵��������;��R�[#}��[��Dw�FT{$G��#j��}�Yd�������#toA�GA���'|�m������茉t)U�n_
���#];hw�䧪V�!_H��!��H2�_cs�n+�6aZ�Gog�Z�����Y�ky!C䂕�g�-V͞������~7�����$\���U�����М��V��i~�_l�?wř��Ey���=ᵛ��n�������v]-R$��g
��PR��VҾ�s�o4X��d��sNm"��]�����M�Sd�fs{E��0�#t�I�I�Wm���d����6��G�_U�&�uz���\��Ş�m>��}�%���fn��V,�`��O1Q��&�~����>lW݌urƓ^�bf%ڟOb����w����Q�a���2��$^k������A�&��9w=#�s}ݵ�^h"2��l�7��ʲ��;��OeJ�#ZN=5��O����[��ӛ��7�u޴�;��ne���2��.��$D�*<1�6/�����2�~���x.W�)+�+�'j�m;����Q���o�A#�f����ϵ�l!�����j��H��}��Ҥ����U�{�Yg+s�
����C+�9��@w��݌�׭�J�4�zO��ϣ9,���j#un�>o�q遜�,oV�>��~������͹V�^���GGp͜��o���3��e�=���ʶ�_J�����S�w~t��+�8�Q��;>�Sb��m�?{�{e�&�{�>��ԫ�oc�FH���b]��3���6��i�����L��ӷh��=�&�+;�߽=�pJ'���[բ�[d�j)�f<�V������'KGkT��vvc�n#m��b3�̨��@i�g$(���8o�W8���x�k//ݻ���C=9C����-y�.�+��=�b;���D@C��.v�@�^C}�}��{����-��(����[#��
zb�´�Hɦz"Ǽ��p ����n���CT�᪹qZ R̚��<�`ɻq���M�ʦ,3��)�kG��9�Bk��hL�ӱb{B��n׷�Ռ�(c^VNс-I�j�U�����筅�7��z<���G�eث��]�/ҳ�x]uFa�w]3��ww�LsP��h�WR{X�Z÷�z�z^}sEW�`*r_L�>���}�YW�Coy^��#�x�&���^�?��r?C��ܣ�@����'�|����lt�������z��қJ�\�8\��c�,9��[l����Ѕk%%�op��r�����c�{�H�T+�M!��`GS������f{މ1YT�p)�����m�x#L����b9R��%����֎w��jwԘ��vG�U�L:Ѯ����Ȣ���A�;����fH��-��HV�td�T��[����\�ƍ7��J���S��Y����dQ�j�U�Gh�H�ܽ�֫�0E�WJt�-^�����~�����O�k}���؟����R�ӗ��%���֯k����W+����g�j�?Q���MP^��ܗb��;�P�������ƾ�m��>�]���G��`?F��WG{P׎�V�>���>�����%|���������u�τ�Cz�Q��V��+�b�oa�����j41-���u��կ֗u������뎡I�۸b��({7xo�1C2A�D��=���m�mt��;^��7ދ���eOn�0n������9�Y�g_�7^���z�r�4z�]
�����-��y;�z��}�j��.�`�1H2�_�=M�Ϧ(��$!��A�����6<;)�5�jlP�蕢��4z����C�o<�j����vb��^��Us�Ǟ�&��]C�hB�I�{�htٝ�?X���<����qvj��{�VIj2v�g6GF�I�XN� N����!��1Y��`�!�x���jP�o��Z�v`�4P���\���nۇ����+��[ƣۭ%��
p����WF��}�af�5��֒t���ys�{�dP�`�U�Ԫ����Zç|����z�	l%�/�b���v^��������{���=�<�ڛxԲ��O�ޯ{�lj�R�����r��׆�����/�[��+9�,=E��zҼ�æ���&�3ޥ���ߪ�[v�V�u\X;%�<y�O׼����J�#�����>�{ݽzwk��q�V�%��ǳ��e퐅�i�������ZHWW�9UM�xr��\�s��q�A�v�s�l��c��������.�c��u��%�t^'���ּ	�O��Q����Qo.�2��u轟,���l����S�;����z�4z߸�-Ռ���D�ג�`��S�~�ƨ63f9!�V�k��q�K����˒P�7뉤&(xvo�%��B�B�2��ߐ�9e�#�\���h���)��-�~f�w�ޘ0%����D.��������7�qEW�Pݓ���9բf�՛�n������9q�Eӭu�)��v("�A���·'FiR�צw3||/����`t3��%�v'I=��e��6���.����ng:T�w��wy���{��������ލ�S��W��o	�+�]��O����=���~χ�D�+	�|��1WX�4�;�5�.t��DP;/���q�k=}�;�N,|*�JB�AJ�2xZ�𬞽�"�}s9�3���R��f�4WH-'}Y�Y�o-	�o%a?0�5���3��b�
DW{˸M��w0Ǉ�PG�j����Ӟ�١��� 5�[��Iv9�mL��,dߞ=_G}��S���J���R~n����A�+����Fߖ�u���ƻ3�*ʫ;��_J�\HR�y{��B��J�!9܇�w�*j�t�Kꥹ����"A	�nrG��3l/=�U�ƽo���]����t�:��i�c��m����m��=S�j���to�����/Ct3�Ou6��?>V4ү��ֻɁ���2϶uǴ��4�-Wo�툥��@��j̣=3�8h���)p�`Ӭ��]+��݀)}�Y@�m��M��ug��-�hʆ���"��vpR�z�Ym<'�]Ŵb�9�&ܧ�]�`��1�gE�&J�-vu���)�I�ケ�u���P��JZ�|=_��fT=�U�c2/[sa+|�n��{�j鉼{"��P5ru{i�ގ��aA�AC{f_xC�l_�������fXv�7�W����},��j�O��?���l��>�_*ڭ}*��GE<�����'��}[�sۿwR��p�3��N]��}��HC�(o@M:57��H��+&�۵�n����Q�'����m+/�B�]b:{��~+���ɫ��_8�@��]��=�˫ɴ�e��G�ڮ�`�'���9��=���.���/І�E�ks)&��pŉF��U��p�FL�Q���~�	��(�j��?zc�5��t�e�f���=�N���XJ�fΩ��2����'���g^��c�:ӕ��s:-O�1������^@}g��� GN�~ڍ�-�䯂��XQ�c�����
��G������������UUE��Q������*-�����6'�>��"%T` 	 B@��P $	E@��P"��@������$��`%D	PN%�G��E��U��  ! 	  ��@!�� 6�G�1�QD�E"@D�D��DQ
�D�DĢ�DDAQEA
 {�QD��E�1 �4H �( E��D2��aU{ eU`%U`!U`$U`%U`! UXUX W�����
�  @B��H ��@@�.�$^$Ap�������z?�D@G��PR%2�����Ǽ��_��=V��#��$utH�}�>2�y�?e���hl�k��UV�3��?_��UE�x�Q_xtt��$6#sXu���6���*����SH;��M-�'�0�&� ��>�7lI�@�
�"�(  R��@@ "��@ @��*������*�*�(ʪ���	
�H��0 �*�+"�
� $*�����H?�\@   L
�� �
��������O����P��"��ؘ��1:�h�������Ez=dЗ��RD�}�����O�TQ_������Q����������ت�+����A���~��c�TQY�hC� ���a�������<������{�<���O���|?������Dn>��z�w�UQEnU��d����c;ͻ�A<�x>���v>V�%UV�8#j��+�3�E�Ƿ�$n�`���>��:q�`1�ʪ(�B�A�#�w��������?���#�aUW���I3u6���+(��];*��2!�����)��F: ��8(���1$-�}JTJJ@A � PT���HD��*B��T IJE*�HR!H��"���t4�*�B��!(�>ت��B�H��MTTT%BPu��.�"��QDk@"$�QUI��J)P�@��%J��� @,�Q%T�Ѥ�TI"������B!"EQJQ)J�"T���ET�UD)P*��*E@��J���EIJ���١��R��  a�k�u��1�].�kv�j[�����p\����t�v��5��]+mN-m���I��7Mh5��[��֡��59�um��lq�*�J
�l$(@��   ��
P��B[��y�AZf�)T	���4��RU
Q��H�����V��:[�R��2��[PݩM�-×wi��p���:�V۴��کҔ�ݻi��i[k��HU(�PAN�R�x   �ך�[�waڌ�ݴq�eɷv�T��2�֚�w��ɦ��pg��m��nۨ�ή�]�J,ni!V�W9;��]4�kû�����u�4(HR"�@DDJ�  ew��R���:�75m�u��w@��۵7www8S�[��U�����f�4�h��� *���5�-����$*�.�:�%J��*�(�x   wo���p5ERuM��)m�v˧C���QU�tp����� �;��TV
�UP�����$%*�$���E��   ר2+E�� {�V�V*��s��HrVU0��N�T��Z�("��Uk���vU@��T�Ek(Ai�  �������4Z�A��j��!B�b��� �4n�+`5EUխʦ����(��r��P �GD��AD(�H�   {�� +�i��U �&  р�P]4  f��@�F M	ҰB��LE Z�����II((��U"�Q)U[�  ;΀ � �Pp;:P ��@�7A��:X�
1�  V-�
;�S� Vd� 
�bZ�R�)QR�UJ��  ˁ� 3F  X�� :�:�(�[� 4)�0��$��JÌ A�� ���r����"��JU	� ��E=�	))H  ��4�z��@ �JJ�1 ���%J�� %<�A1U  �J��3D8�I'�gy����Ƥ�A��
���(�^!�yet @�������������8㻸�?�����w�������N�;����������;ϟ�_����V�(��8{h�ȇq��y#{V��m���u�(k�n@�c���Sh��mAW�ݻӪ���23����bYB62;�.X 3�-��w�C��A�vɓhe@�"�����%
�/�*�V��i���z���vj?�Ь�ZeL�pA@:zf��j�ME����L�>��n%x%*����6�a6r,�����2�\�����4��
I.�Vᤄ[.��OW�*H�jR����;J�R�fIA2�kJ�EG�%N�6�YX^�)��)iK�7.�cJ���[.}dK�h`�!n�Q����3.J-�F.P�%�L�Z��N��DF��*Mմ(
�ī2�GmZ�Ѭ�VF+��\��yb	��0=�۩4��S��϶�i�uyb�,�۱)�"#hҬ�N��X^]��[J�<�s3w�z���ab�����M�T,gƃ�J�-;���{�6d/D(D��cU�����l*��\�el����Mi�� \���M�!P�/1Y������(�V�T6���sn-�K?4^RT��+&l�OC�(��k7��]�����Zp9�\̇i�J����!��ǋ��r����*���Uq���T^���W1�U���R��{�%�E*AL"t��$�6N��z"��&��l�*�봢�W��\�
u6�R���4����n����ؑ8����#��sE�Cff�e��ɴ&�[��v�#[���i�
�cC���]�W�`ٚd�ő$�f��Z�u�Vi����pJ[�q�ŋ��M�5�i��
��oI.�t����� �`)ѱ�Tt���7(
-J"bx~Ɲ�s�̋Z�e����O	��m���b��ܼee�1��4Kr��Y�^�)i*1kY����2���O(�}	*e�_Yw�^l�
�Jkj���L,���pd�^ڲ��lc1ٷ��t�); �m��v�ĊJ�,8�X?E�6���n��0k�vat/.�F:�l��X�Ƌ�7Y��Qytj��^껑���&t�d�ɣ&bD�!ȶ�Z����mfh�r�[�Jkq6>��
Kj<[�(�wE��<�ٶF�nܽ��B�B7P�Ŗ7r�5B�gj�n"pe��$V
&���X3f[��p�$֛إ�)������Q
X���0B�ac?3Zr�Eb�J�ACI��X���8ʤ,UJx�I,�C\	���Y����ҕ�j�B�۸tԧ��	�S0�Ez4�oof�G,��/A�U'�kQ�����Q2�n�="��-�JIAEv,�\�CrP���]XQ&`�^�4�J���t�J�V|�<��E��6��:s&�������4;*T�`H�ZP*�$����Y�]lոn��ܔ5(���P�M�٘E�I�U.�իV0�cP̛�������MZ�l�/2��+i5��.o�n��O#
�b� ��!�2��
����@�i��v�ϝl��Rz�Am���l]֘pZ�See�B��0�ܒ�>��,�f6ͫg3#�,�8�����7����&�۵��QCr�� 
���5�j�4(�V�ej�ֽ�׉����Z�YQB�n
{��&f1R�ܿ������f�C+.�;u��.�j��/5���L >�ؕD=��K�tV�9��m�{c%]�r��b)�C�Tr��W!,���E=�F�m���j���Zӥ�*�2�t¨�i�sB׎�R���DZ�SC��Z��xu\�V^E.Q��,bKU8��]4��^���n3%1�b־�
���ڙ��Zt�t��̅��S�Uq�n-W��h+̷���d`�p�2�I�K������b��M��z6����˦*F��T�V�h��dQY�]��� �[!x�㫺�T���ݹXf�]�.8 D;5�j��?�lV�K
����f�������Xi�іE��X[�̅ᬌ3��cl,Z�ةPtr�@ڬN�N�5�iM�1�W����*��,�Z<̈���E�2�KSjM�CcR ̳h�$ސ��C{ 6Qܛp*�0*�"��=�{(�6]´�(m�.��d�8J�c+abe���[��-��׷wf�0m��cu���R2sqD6��)#�B9[��U�"��ޤ&kFڎ���*"X4u#4�203`�(hݺ��-ݰ^1��H�HܩD
��TUʑf!�q���5�֡�t��4+� ���a��@դJ������NH��zU(f�[Goq�k������v�A�ksE�V�lV��[YѸ] ���x~ٯut�HU۸��	Whd;>��5i��Ѳ̽���k�	GKDZ�n��ۈV'���Cp*i\��Xʚ7vYX"rхj�tf�M��i��3iZ�:�"�U�\Bdd^�o6�b��]�ͺ62�"M�$Z/]$���/k�`��F,�Bĺb ���.ݽ�Ϟh��Y�;pQBm�z�nY���@0#Ѝ�&�ܭ'��ϥ$��e傌�Ӄ�,�陆��w,�F��!
S�H�h��yuV#���E�N�ʛz�teKx&M�H|X���a��K*�2�w"T[���wK�X�
[vE��5���CE�٭��l+Z37��&fة��i��6[lӇ-�vh���m��Jʗ���k��Ĕ��ǩ����,��;�eeF�/��M��f�N7��w]��@c���˙Lr�&l̓�����^��fU�4.�)�٠9���kVe��31���]�X�Ӹ�?0f҆�f��ͩxi�.ؚ�%�c��e?����.��W��ۂʺY�Z�f��r'չ�S��ʬѯ�oF �#��*�EP(�$��Y /���cx���K7�E*
�L��m�Q�sX���;M�m�a�Wu.�S�.(�'I�9���
i�Vu#qKu�Pߐ��/rک��;�غ���7a����4�ӂ�00�խ��ه@�ē%�F��B�.X2��[x*7�m�u�0��k�T��YLm	����6�Li��lj��&�`��F����2�OB/Zu;7sG%�^�=-�A$vb1@l[�N�=���uf�(������Mc�[���r��j	
�����u��������$U����a����ܣ�*4�i1�Z#2��̵�_٩���)�L��ߓHY�1�m�V��Oe])l�lMl,�R�`�)7B-�T�)�Fe���ʹ�7A�'�c`��dP,��F���M4�
�H�Z8�M��YWAV���t�.B�W!1�4PYoF���wn0�R�F���4)%z�%!��5��+u�k/Uµ:�X��OV��ˠ����_כ+X-�S�gE�4$���"����ƊѥǸ�^����>��m�!�T��)|(�c�sK�s�j˥�P���#gpؔX*P-mD��J�t��j��`��+Dtf��Ku��ū[R���ɔФ�Gh8x�唎�	�\J��^���ͫ����Q̧pk���&��n��/9e�����66Z�7�?l�t���e���aE���ӣR�Oh�d�ս�A�64��DU�n0f¡ˣ�h0���%�ź�k�A	7N����6�3x~[djX�V 1䑑2��U��U��/q�,�-� �m^��5��wx3@��Jܔe@%��-&�nڠ��[a��kPx�=d݄�q�����*Ǆ2�nf�qc��{�M�"�c]��2�q�FN��5�P�(a�}���3n���+�9w+��0<��(��{Za�Fͨ�v��]�lm`�׺�rNZB�&�M%5]��!�S6ZJ�n��+���@m������E���vt*zCǦ� �̶�YXbaAX㵡0ڧy�C� �I��b�m�)]�Ú�ҫ+E�zكk�lYB��l%n��)�)kw��)�24�JR��/4:��a5���Q��f��R�I1Bؙ���\��b'5c�%޳b9{Ec��`V^]�	��B$TҀ���I)n����M9hh�-����52�ۏU+ bܷ��@�b\��(J�If ��[�Z�%,�,cӮ%�u���y����ű;���@����*��[����-&��E�V��t#�O,�Hc�f
0�#��%rS�1�)a���X�X�X�U��i��"�O��R4�vY�%Y���%�B魸/X�D5�Y:	Vn�Z��u�̤B�s)&�P:�'4d�����}u��D):?�qiu����ʈIl��s�U�X^�%�{�Xg5�R�o*�G�%i���
����6���P����5�c�-�1����֧h��{.�҉�e�b�[W���H4=�]5YCc
�˵1DF�ƅ�͘��0�)n��l�`��.̘��ѧ���.��6��2��� ��of��ɱnf,�s0�:�x�K@��6a,��NJ�&�{����^d�1ǣ/uV)[t��y��p%1)�0�2�Ŭ��aT��z4V�EGдJ� �zw<H86�0�4[��.�ƫs��ˁ^�9��Z�f�H���m�Œ���㨔OI��y��Պc��Ў-�6�d7DQT�J�K>-EV��B;�d(�����L�Z��Gy��4.�9�р��q݀�eR�[J��l�����,�'i\��C�����2r�d;���=�mCaԧ�Edw�h�T�ڰi=�wzF*YV,��ߟ��][���+2`�v��F#f�jIS�\�6M�ͺ��\ń4����-R����jb��l�؁�u.�\�h�rG�HlP3:�0�Z/*1i,!�B��E�� �������Hɭ8��{mK��Ѥ�D�DR*Q��2�|NM���^PR�LhӸ�c��&Y��	G(j(��鴾7�i��۬���3FZ�Z[��P�֔�
��Q�qVQ*m	K[H�Kj5��t]��K%E�Kst�S�H*N�xXel���،��AdU�z1���K���T�ٖ ܔ�PcrY�t��	�%��ƶ�5��L^�!�רV�z��e k&��xXk�x�>�m�!���to��.���Fҭ��p�j�"�)M�a(����BѬ"ܹ���i��x��Ke����>YX����-���Κx�ӵ���D�%������H|W�c�vsr�9d����:��]�A٭׺���-�Vd
�9�+F��YXd���k���IC%��<u�*����i��mV��� ��R���ѽ9Z�]0�;/h���x�d�������wWVɸT�y����UZ���w\饐n�F���9W�w��#��P@ۤ��X�[&�y��,ہ���b�>�;������\��K�5+ͺ;�$p��u"�9�Ȱ�1yL&R&IV�Ɓ�E�>��C/b�S���Ȟ�$jKŸw4���It�5o歺�C)��H�O��.�mlIS�>o곊���$b`-Z�!I37/q�o�hb�//1˓%�l��
���Y�@h���2HX��W��:el�8��B�b���Ɛ�^���:6������k5����It�:�ۥ�Q��o&"3W�J�fԫ�/Ż�BkP�v&#�6�����F%��.:��e�jwp"�q�Y�zoEֈH�.)N�u���E^U�f�H
	D�j�I3._��GV�Q<`��e���$6&^��rk�,46|i�)��� �����KrF��]���&	������ ���1[h0n��ܣ�(+YYN妵2�fbU/C�N���J"Y��eӅ;�V�$n�x�7l��>{L�n���Q1��D���N�Y�XPd�߮�7���0�jkVM��v
��e�VNM V��p,�k�r���.�1�=B�> ;D�#~�	y�����A�q'�6�vXM}�6��nJ�EҴq]��pP�MA��Il�P�-ԍ9����J̫��З�%�i.'x�������BH��r��J��5V-�p����*a͖��ۙL��Rq�Ӭ�V����L�7-"���6��i�&��a�)0����	ʗ�SK5�P�ln��=vh�5�ۥ�p��z�DeǮ��P�����;��re���W��͔�SAlX�ݢ#kh���.��i��w.03[u���b[oW���D�Z�٩���b��*%�I�G�@�)�'d=Ioז^L���
�4��X���+�0e���bjn�p��S۩nPQhGqX���7�ssM71J�����˺�k]��
�����&6�|�TL��৖�b��%c�t�>*��m�n�+p8ͩ�t��K��V+�-Ѷ�a+ius1um��@f#W�F���{rPZ[&ėŠA3⒁�)3B�l4tp�X��>SdO#�b�m�I��Y��ٛ׽�8�<z*��LԄ�)�P�"ͬ�Y�1Q
�d���b���(�n+D��aة�3��&��r�e�E<Ɏ�F]��ff�D+��V�GZ�*vd2� w窋�[�囲v��ne��5	�S��O-�Z�j�x,��c�jS��;��h[
kt��{
{	����P�m���R��q�W����mJ�S��5l-�4ԫN��2LBU�nAk	�W�C-�;������$D����w����>P	lVVց�w�04鄓�l�φ\�k(mcՈn�GXN�̕��K0�`��\�������R�ێ� I03s.{�f�3P�n����\<�J��̈́�V�5Hvol��y+̢�mcE:+o&�R6�GH�g2�qR�*вU�˲X$=(ǛA�(��_�Z;wD�Y.�;�Fh��r�J���ʳp-�hhf	E*fk�nnŭ�GՑ�'U�:�s�Ṋ�9��ٱq*ܥd�w�q��m�Ny��A���5n��V��m�����*p;۾"��V��+��AG�4쾓�Q�۹�E�	����ݸ/�q�������0Ϋ��k���Fn���J��7���3;�*<WL疤��C�V�Β瓠��@wh�喴�v鬮���n�j���s�r�rK�ڶ������ᜊ�Z$���E:�wT�ҒØ��{>�ji����U��u�\�On����N��� #_v�W��m������_!/�;��>�+&P��r]�A2��1�9�o:nhd����
�,���XF&�|՗��xz�'B��5xk�
�;.S��V� �
Կ�.��X��y^�A��t�
��ja��u�ֺ���:�I(:����Ӎ��Y�ZՇF�=+g�W	7eg+\�KO��mE>8����n�}ݝzZ9��9��"�-Գ\=8�67���kF�&b|wk^i;3ot}Ɔ5�Lz���wn�a��\�Vu�������oU�[f�n�y�,�QL�fo4������u2���L	j�C�p��3�q��NV�{R(�ZGl�T�5�/�/��'Px���#̃8(��l����GMA
�Y�t�$�5{��l<㲏A��K+�H�r��n�_^��<�i`��e�fd��S�㫱r����ocjC7kkD,���W�WA�qh���e��i=�Cb�^rt��4���oP.�-wRW�c	�g.4-6�ӇE�l|���\kr�	e�D�3�'�]�+&)�D�w�4������ጭ�D]�l�݃�!�ӆ��q9Jg%x(��̳%g#��w)�2�j��lH�S���aT���&-�RVt����޲4�����Ί��wbO�w!ނ���?5}e���I����RB�����2B^b�ԖNι"%�,�q�qu�<��m��Oe��w*�s.r�d��w���ݬp����]ҭR��rT���]��6����2ŷQ����ٯ�o�q �R1Jq�����{��q��������2{�j f�c�S:��|���X6x��䫛�rB���/�V��;w6���{��w�!���\܋�(�u�@Ru����eb,�fc0�t�7jvum�{G�(��»�Wf�8�v��e�O-���_ė(�Nm^�u�x�����6���<�R�f;m15�f��#��^$�,ܫ�%�w����&IݺMK��齣�F��+�R�Y�JSJ0P�3v:�J�뙛o<L�Ё���'p��و�]�ȋyWF<�'>��-��X�p�v��H���a���3�ֵ�vw;���7�sf�&iauj�r3;x�.�2���u�V�	�:A�����ђCҒuyF�S���J�e����u*�
�[�#�E��n�*"�;�
��7�su����K��شE���cC� `��������G����IT���K�T�Cx�^����0]ӳ��w���.
C��~�0�QK8~�ۍ�p�P�s�Ju���8�cj��Ob�����v5b�Q�F��TMW3�j�`�u.Ŏ�n��LQvA�)�{��$,X�&e�%����9n������ӛ��{go�XvYQC3��U^@"}[.-�V�[�EE[���+��6i>��x٣Ag*�J�c��-11Q<4��=��� �'t
�O��kK+�E�*Q��Q����Wd�q�x+/�m�m ��&�w+E��A����b3{;#:�N��:�J�ڨ�F���TZ�9ZzT�Y,��J
��4*jn���n1h<�7g��H���܍_�B�͚6���sa�k;Nm�e�J=���*�	�.��m��&�����G�Bl�ɝH{��M������'K�$��i�m���	�I��Y&�8��Y�¢�����&Yd�ޥ{��[ǲesC��dέ�UF��B����73����7Ԟ:�B��{�i�{,r�0�|���.5_<��zC���������b=��5d�N��Z��.FVG��m%;���Q�xc*⿉ε�Idl����嵰VӼ��׹z\�FöM�sԭ�xK�H!��`�S�Jf����ͽ3��YY�w�ݍ��3f�u6�p@��7�7���b����`��ͼ�^P(Q�r�f�<���<�:t��]�D[�Ҡ�ֱ�g��4�D�7kF�#�f�:�f��t�O.��ޠdV��8�����~K�+� ]a�Z�NQ���Z�7���=n���t� ��7,�r�c��A�̵�́��.��Az޽W]W�oS�!��Sm�W��g-���rx�k�Km����-WJ�����f���Y���׋y������3O5�v�D��{ҍ��a��D3�5�q��դj�GN;���b�� {']Cj�wB�$&���D�W�dX2�ف����+�G����%��v��9�ζ�v)���L�ݖ�V�ˡڴ+����FN�[p��]��@U����r��0nb!t��4�vZS�m�K)`RD�5P؈'/{VfpfU+\��us]��k���j�%2����RԤ�������+|�eԻ�Ɵ"+����]E�fB$t��es��x��@�vzi�c�W��hخ��t��ulΨ.YZ�+�ץ��h�ư4��x�wK]�|��Ֆ��Y����C�iu�M���Z����S��T,i����ټ<nhT*R����v���xN'Ӯ�j�sOQ%^���8�tiIإ�
����+n��\X\�RXf;�P:��֝k�Nv[NX\ml{��1s��j�t˅(o��s���k1&:���bܴ+ˡ�r�����=�{�h�i�2�׹�^��i�Jb\~��7��őÀ��%:�㣔@�����u��!ɚ��O:�.{�J��^�iYt�FT�v��#y�]����8�n<uf]<�K�L��o"�؍r��ޭ����=2�#��u�h :�]wֲvv^'�h�_���'+䟼��r�%��2�;�ks�:K#�	�4�����꼇/�I��.�v�b�K!Íc�������Վ*���!�M��+U��u�w,�{��'���p��ܸ)ۤ�d;V6�ɽ����w���}v��K�/Z�/�#[p��۳dvw!�w˵�ѷ}�:m�S���3(�d�QJ�m�ʾ�-9w	�6��3-��ga�O�J�$+6���F��<A��U:�d�,4�u$�Lob;n+��l�h� ~+���Y����jj�tJ������uuF�N��9�D��N�U�M�H�e��h*�Yk�WٛNj\�1��[,�Q]{GZf�o(���i΀>��j�#}�_:�7b��T����0�U+4��V�Z�c��5cF��G�L��Yu�&���0e.�֣�-ή����X���s#����[�Ա��!�4__�vs�X&F��'Jˡ���75+��|��e^j��Y��'ZO�MB�bE�ފ{l���<E�Uiosr�j���˧õ)E���d���6��ث}�w78f��)S�3J�3&\�7'WnA���/�(�g0�Y{�� q1�u+k��V19b��[K2b�Ϋ�`�L�M�-�T4��̩v��WY{����ec�G 晡i����}ڥ
܆m�b�wu0���J��շRy�:e��1���Q�7�{��f���qU�G�i��̾��\��>��� ȓr��S�WC�%jV����
�lX�6H�H:�L��ܻ��3�x&��a��g[�1�r�Vl�)^�����q�6���ᙬ����VzN��L��Y4.<ށ�}�fĵSp�:)�F����.��Zj�����5���G�R�5	n�3�i󻧜��V騬D�P+i�)�QV����*u�̆f������w�F�4H!kv���CR�]M:#r2G��̫��7G�����*W�7k��'}CS��ƮVd�3�Qƙ˩e�dC�oUw��Q�w���*��@����V���-��~I�N�� e��=�j.�wȮ4��5��W�غ"�*R�m�}��L���M�UcY��:8陽\���p|&ʼ7QQ�o�ݮ���K����sc�^��\J��\_G�����=t��sc7ԫJ������S��԰�H�\}��M���ue*PF����`�J���zX�pAS5����k����#�2�A6�Vcx�W9�e�Y]�W&tj*�ႵR�aNs�Φ����]����)�*��ל��R���5�M]�2�[�xY�O!��� ڎ��I[�-v�1�(�a��uת�"��n�̡p�t�B��泈%v��3{\�zWp�Ě��}s�Y��Zv��F�	�OM���}�|�a��3+��<u�Tф��;��[Ԛ���.
R�����xtL�"��9��v�k��ض�[��3
oz�⴬�n�wU0{g�+@}�I��J�y�Ǝ��ɤs��бi]q��e>���g	����1Ҭ��o*���(��:���ሶ�������u�t���k�kʕän��n�2��2d��J��a@�בT�i��b)@�f��[��uҮ��Nm>�js�-�<�;jN%gIa���&ݣo�E�P��rU�xQ���7B�SZ&��̢6vm@Rl!e���g���r&���[4��5|��'�p� +N�d �Q{o�+۽.�Y�K�0>@�*���s�����Z|��B%��}��l�K���_ks0�ss��L�	�*u*��r��ei�RC�Bŷ��m��j��.����{�i�क��ʝ��[Y�����]r���+fL6Cҭ+[����h0��3:�S��EE(+S��Nwn�Z��j+԰>����+��M̥K��^�`����ǅ*}�B���Zɓiv^�/k1��Ot�c���یu�Y�����gmB���]-��'�AS�/�=�2]p� \���y���]1���ghΥ]��@��1�1 �A���wf�:e��0�z��x�A���tssvֻ��@v��)�p�l$�
�L���R=J��|�GF�S�D�D�$�-�W�eS���j � 3��]=�[�ܔ�0Zܳ�7�\�cw��N�űV�Z�Y��];�t�TĤ��_wט�6��,���UÜ��r��YF�hE�E.,@r�G���竸��i_gT��.�n-�E�˾w�$ �1��AU��\z��B�ʰ���(ó�]<!���zK���8��Z���ƛ�9�����̩�3YڲB,����ّY�G��5��ۛyS���2!A�"�c]���%C�ӧ��K�Ŵ��Au&�ٙxH�F���:+Cë��@��v�+�镲���҅
ˑwU�x�&�bi�� -�7�n�^�m�8.28��Z� �kw�D!뷗`��#V�Q^�y-@6n>�{K!카:�l�@��N�87>І��:&���}q�d��(ћƯ��Zn�든��.��{;�z^���&(#뽙��G/�.M�.qbu��Y��F�fc7�s�Z�n����8�>]�����51�k�r�L��vqwWmW	�l^GgI��V����K�Jc�t�[R㭌Xy��{�G%��]nU�h�x6�H0�Q���0<��wZ'n����h1���JA���:��n�	�ށ|
������ַh��u�M/�pX:s{�G!�"AyJ�,�R���y��i]$�oszZ\{������q���:w��3c7���s��C-v�
c}+�}K諉�r�e�H�}��I:$z�;�ϳ��zu�spH�ga����3h�V6k��mhCt>ȘČ��B�� �������	^�qe.��I���T��VVB1GJ�o2���2�P���}c�yQع'Ln�+s+h��VDţ��2-ϗ՛P\��1���>#0�X�`�*^n8�vjC5��� �K{q�+FhD�j�����V|�'o�p*f��i�}��Wsm't:}옧^�ւ[a|f�:��:�9y�jj�o6k���9���/��-�JO(���Ր2���VAܩ92J�<��Ov�}��EF7y���W{Ղ��%SPBL{�pE�4JOT������(�ُ^)���wMb��U����t�J�]Ҵ�e����Jm��|0wf���wI�25u�2s�+&ۤ�\�1�u:m�
�
�ú��k$�V)��ٟh/�#XTց�n���4�}��wi�2�������j�EKbꔧn�"i
4m}�+<��/0 zܜ���T��s�>�;+g����S�W)7�-�V��
��ܡ]�t#x�`���V��D
��ʁg�����׭����m��`���PU」ʡdy�ڕ�:��o�p�:������׏�_D��/X��6]�Z8Y��D��TJ�/y������E{l@30:K"��v&l��dk�[�����u,6ֲ����]�)�\��w"kv�^����-���q���f���6����Zr�#��&s%��*8��Z36k�����1�����m�w���J�<���ec0�:���^�9�g�m�3�?�N�W\��T��1R�#gh^��%�Z��};�^T3W;tn�"�bٵs�\'�aos� ���w�kx�]`W����k(+1bI���8��A�ҀH4������n;�Er+�1��z���ܱ�z�_$�>�v |y�o.��cF]��t�����̛;o6uΣ�Eϐˢ�*��oBsu��縱:�q��E�Z��:���!7bQ�6�nl�%v�g�p��`����6C�*v�ܶ X��|:�Ǽ�����/^�KU�.ΜK��
�͎����_c������i�Or� �p��oxٜ���Wr��{wwsv�׵����  D��"  @���" �����]}	c޲ϬNd�~JD�P��On�Ε��	�(�_s��t���tۍ�^`b'��/����B[&!��n�\H�n�e�M=z%Y��`���!{��6Y�oz�ܸ����v��{5���p;����z�j]�K]o'j�������K�<3�+���r��"_Z�e^�339�6�Q�'^�o2��'`H@�pv�X���:4ko���|�bם����h7�2�u7�z�[��l�BݮO��8ݮAaZ~{@�����׆��N�ĨA�֍f�J���yM͔SX�Ãg;9SP!!�R��nt�)y���eF"L�.Е�JT6���#h�i��!�g 
��z��Sλh�%i\����I��IKj�e����M�ؖ�J�0o�ח���u��gʁ���"�NKs+S�m@�	[ղ���
�Y���B�3C2��ہ�Є�p��XA�����W�l̴���Q�M�:�Sd̄v���ٛ���O~�ř]�{ܨ�Z������I��{�p[�Y�8��8/�U��j{D�Y��иow0�B.�͡�5GRǃ�]��~`����6��U�����f)�ܻ��T����C�6j�|��v�;�$WI	��}���;�gM�r�Ҏ:�͵X�{�1]��+Ew��Α^�ӠD��^�O<�E�k!8:'kCD�fQӕw3�#�ː�ڴ�ˑu��-u DS��ϥ�k���իN�6pQ�%af�;�C�L�/8�܃+�`"]N+q.,�|��e	C�l��\7fd�����q�P���1�u�"����WΉ�s4VtǮNO�3���5qh�9x��{���Z��+�4��t	��:���83&�������#5g.�L�F�lս鍽�6���I�!F>��03mfp�b���#�)W$ܭ���4�	9�t��Œ��u��s�8�f�FCdVX�cD��כ�X�>t�1����y�b��v�ҽ���hcvJYpR��s��#E���ʔm>�lS!�t�7����Vn�n ��A�l��� u��e�Ջ����m���]�����B��o;U����j�S�Ը�u�V�X��!n�Bx�����kM0$�^ -��e��GԷ�
�
#j+k�kyC�!�(��e>=ETܼ}׏+���Ż�h�Kȝ��1�n��N�ab^M$��o$	R��=\�G1oN����͆,��d������F����]'e�hr-A��{J�:�yX�wBy@�Fu�t�=f}�F	|�2n�f��pљ%�i6FX����i��:+7���XW�vH5�� �}�.\�:�4X﯉�G!�gF�R��Al�ۭ�RwR]��݉�Zv�FZ�F��:ujّ�j�
�8)c��c�x+����e+=�n������Yu3e�h���ES���6���:����l�9bǤ ;��[A,�6]�e0ĥ�
�Ź�;T���ܷ��f�q�	�z�q��-�\kK�<]�nr&>/8j�P������(������E5;��F:t�����G-ó;��R� �9��sp+T��z�oN��G�*��sq!h��#����/7+�AM�=���B��L��e4.�ݨ�����ݬ�����-�$���q+��n�Y
+�u���F��\>]q1���]��f;����������)b���k�²��쎶�ulD�uu��R�[�9ؗt��H@x��.�3�%�4�bÍ@��QCwiR�SZ�A��:|�(拣V��;�U�zv��}:�ݍ�Ӂ\Q�� �WgP��Q� �v�S�t�++�e�@ #:Ν�D�A��h>����f��o�[���K��v�8�+s70"���l���&�=�F�Gڎ٭<�ђ����)�x�V5�$�����# ��X���|y�0t����ã�/�w�NE���v�gl�sD�*����sk(�Ϸrn+Ϣ����E'Z��;"��Y�'�v⾉mc�\_MM#s�܋����]gsڧڪ4�nD�i*͜*^�M�Yѣݎ�6I6j�IM���09V�����Rgi5�r�]���*�<��õ:&�LT�����Vk�]a��^g%c��VNJvG���LF/�r��8ЗZ�	���6�s��+,�@7Ջt��V��Ab�+d=T[ʔ��!R���$j?�̜��Gh�w#4}+��S3:�C]��֓�K<�ً�O!������XoML�nl�H��.�mږ�����z�*�)�
�-��
�r��lQN����R��$}�+���U��6:?���ҎfУl�+�K��K�uʛ��N�Ύd��'�NF�B���|6���j��~a\+%_VN�b[���-b���
��]�n�N���)��c#l0�ч�G:���)g��Y��!K�8�g-�e2ܘ�4��5u+�U�#2��D]S:ϫ��¶Ct�B���P
��������;z��5�˖�e�����t�8����;Muv$z�K~���L��9'}X������p8�w]Ü���[�VT�T��.�͗|d�P�3�'���wS��恮����� ������Y�,�ʽ�=��R����k��	\>���}��%[�=�(M�fk�j&�w5Et%֫��"Hr��Y�)��*Y��|0�uj�v�s�����)��]�Pݬ+mp�=��mV�"�����I�fc�o23:����^ZO �k3Eb��J�Ş��b���9�J���:�`�"oC|U��q1,�YX�c[�e�,��4�\�gt��&�T�����
�9���"�;���
��@�dB��U�E�ħou�<�%��	�O���n���m���� ]� �}���U�߲�����[|o���h�9	`�/��٨�u9r������WS��h�Ƀ���/	�}	|3��I��y+"����U�W;�yRʃ1)�#�D,*���1������"�X/m�Bq�!�e��I�b�����/z�]�EGw5��-�{�)�����2��N���A��e5�7@r�R�������lP���R��ؒ�����Ձuz�U�-9�M��ϲ-x�%E�G�C�1�3��y���7]��:�!��Z�h���q�*������;�M�u�l 9V��t[���ĵ�`�}�q�����v��]����)o	o�xP-���Jܜ�ճ���u�n�E!�16Yі!Y�����M}����[O'���F�huX4��v�BT�¨j��n�W'�Э�V����c��wi�55<:�TM�jY�^AR�f���A5u�L'e-�a�ϝg"a����=<(澚�qk)r�8\:�G��:�;����\wV��^R 8'J幝����Ya@�ޭ���ec�3qW�������v����,��{����}ݶ:�Kv!b�|ԩ�-�̺����K�C��kv8��ˑ�/R�꒝�xe�ѓ��Bx����S#5K�wә�i)�S� ڕ��|��\�qɽW''RjgGQn�]ţpR��]FwVr�p�+� �jYf��듻�T�%M��oS;�D�Pfw`f������aC+��n; Ⱞ����hds4�m6	{�
�X/�uY��r���{�*s�۾�r7�uW�W�BotV*(�ܣ`K���BOw�gr�ۊk[3]_qȳ�_>��l �V����-Q;°��cQ|`�Nc.핆ڬ��e�0�X�K���TTf�������[�ެ�42c(ќ_w.ç]��3�r�����'��[km�W:H���_-��?�oK�����}J����쮏��}uKM\޳�f0��B�Hww JQu��R�aδ����"�V��^���n�x�e���ۢD��D�X${��������mU�w�0��E�r�b��:�|���j��-���������qj͹�j񱸺��Yn�;M�U���5�:����|l�t,�yk�����Tsu�dݱ�]���
�gs�������]�b�e��Sl��Q�����eD��MoD�y{���0b�&��e����m�=�H�>�EĪ]20ur	�f�X�苉�k�'g���<s��.�Mw�o9��y��|�*�Oe��5��gG����Jκ�j�1�������R�½�FpV��h���k�NoW.�L(�}��E�F��S6�+�H�nh�\�⎛r�H(P*w�5��z��1��šdX^U���A��{u.�0������pu��(r'�+V�Ý,�k��-ذ�+D�`b�k3�)�O�84���wt�&��N+;�EУ�+����X|�쌪Fj�l�,	-� �����AXcs����ԩm۱���'�^�����m����i-�k�9�,lQY���N���ˡ����mSb� ��l��ˎ�V�:�3�n��  ї��uj���W�����Qj똇����Ɨ_'�j�r��ڷ�;���gC�����eb�ޫ���o�l�3�s�u�ӗJ@��ѱ|Q�z���Td�x��r�6�J�1��*Ԯ�7���W]��KXp����(�!j|ސ����Lx�]�Q�w�/_g�&C���j�Dȩ���y��NhKXK&�F��)i*su�"��/jK���仗p�����ۼ�f���v<}�ؘ��[v���^a�L���m��EGnWuR:�� A�M�V���]d��2���ז╻ۦV%�n"|�D�^R5� �z�ɦ����3Q��^p�Wvwc:�ꫛ��|t�[9��[}b����`�9�V���k�.��
،��{�w��NM�ѝ+� 臷��4h��.�msW(;!�0���D���̭u�w�s���5��%�%��ܵ�(s�}�Ȫ{�E�Yw:������ok��f�cuX�QU�(�MȺ�he�������\OZ�fY�ۜ���˩�d-u�m�I�.c=�bc`0o���eՊ�G;�j:t� ��ƥ*9ۂ��k8n�i�V��v+��;�O��x�w� *�Bҁ����\�F��7����ڀ��t�ZLdfVC�&��v���$^�ˬ��ö�z,���[�2E��]�2��铡���R�e�\�n ���a�S1��TU60��2:���������	�|��FSŽ}���귱�@S�n���{-�U�Uƹ�D�����1H���	s������O�V,���:�3�	7�4�sr�N�sW_o^ҕ}��QI�f�4���ogp�[�2�"�gCؘmi�ulY:��V�k��u��\��ξ��M�롈��p���汜�j�E���jt"�Y��a�Մ��P��\�C\闹nQ��K�k��v����K���9�Sz�s��/j�_W�jӹ�(���ʙX�:����y
��e�V,����#涮!m�K*�j����0K��.A�o�WN���G}�ʱנN�z�� �h���Ү�6eff63�yhP�x�vu������Z���Z��%��ܢ	�z�_5�M�����w������6��.���UË׃��]i�԰CSMn;Fӯ5�����6�*a��&���:S,J�v Z��X�����h�t��9��p�`������j]��=H[��J'�<�i�^�bQ�K�j6�k�M%7RXּ�o�v��X'R�oj�|m<f�q�'�qqdf�Y͢��X�豤f��k�׬`�� ��Vi�C/�j����6!��E���b��(�k�u��r��&�-FӰ��6�s�i���G�W󧧢1��^d���4e�Z�3�M��(@��y\+�3����BN�j9[�����r���H�.�}*�f[��4A%IU�E�Y]w��@�
�0�ɘ�8-ٜ(�Qv�Mv�u"o�A�6�sv�.|���N�u�����J�y��KiQ�*�͋uK��E�Yykuz��V񃸦񻺁J-�DU�c�֗����]h[��,�4�r��k5�udM%���w'tB��đ�7�J�) �"�������Y[�UB�Z�d����Z��*Lv�ڲ�9�U>Lٶ�5r�d�j�;;�q�F��.L�>/.�n�ޤ���3B�]��Wp����ɓ*D:��7�o/� 5�;�-�;�s%�fQr�ʹ��w{u��(�z�Z�osf�
�ҡur�P`Y(�82��n�;ZXW2|�&Eo�Ѕ�9����-�^��w�:N7u#���4"��dR��p�&s�Ƨt!�[b#���B_}���$m��]Ȝ5�Ϻ�rC��.��`s�jQ���f�C�W5PW-5lw
�j��u����#h0���2��|�`�;Y8�����A���k��@Xf뛬7�q<��y��ٽ�qT���3���w�`���C0���V�ê�z(��r�(��{���\3.�e6��C[�+�����:�|�V+	 � 'u� ���wt�?�IK���Ǆ��{Q�͞N
������iС�o��A ���R��4���t]y�z9�L�3��wfTQҤ���u�*9`C�ԛ[W���VqϺ.q�hB���+jఅ���%�iy�n��W+�w�x99tD�o����7i�Z6��7ln����ejZ��)�o%ʑ�Nm�V�s�J6���F�8Z�Lս�����ȶ>��Y�N��bPKY�nނr�)ݡ^;M��o2�X��-��ݼ�A�<*}�A��Y��/�x:C ����-���WA�8�;�V�Z�	�_8���X&�Ҝ�ϸ#�������+�s�X�/V��Fcj�>2��]�]�T���0��]�ПM�q�5�J���N.��@�|�N��m�vMr�H��غխ
�s#�V騥v�
:$�������d��:�+:"V{,0�^����,dbk:Y՘���^A?gީh�f�g��PD"/����R��������O��l�H�w+
M�bkÚ���Ò��*���]���Q��G}:Ѿ��n��y��8b7������#O3��U��\s�j�݃�av�ٰ|��o�����qIkӬS
0*�hJ�]n�a&l�a,7��@b�ڽ�{��c���rXN<��i�w��o,���e58��D��5�o/�ڶ��ZG9�h�\���'/�������J�v�M�u�c8ۈ>P$���<�2p�D�[�3�S��#��/�g;�^�9_eZ}�8�W��)/����2�����=HQ�s�Wnc[��;p7P]c���G@u&Ђ�u&a���;Cŭ�y�![H�z�­ܳ���5�%q\����R����ܑ�p��&��n��1*�d�z���Y���z�;�E�����+��ӷ�ީ7��RY��HK/��ʦ	�и�ۣ�c��\�4���B�K^mX��t��-�z�l�Az�n7���{5����[� �4`�IQT�Q�(A��48�+
��s5 ;�q��/J��'")�����Sk��"�c�c�GT��7w�z�q�.�kŭ{t��\���Է����P���$��\�̧ۍ�Kŵ�`�5������lh��`:�֧J}h���J�ag�����'��pcJu.���r�qu��Y�\����Vz��
��Z�cz 9TJ��W�>�T�y���1t:L���ReȪ/#��۬�%yyX��.�C�"���2�;	QQ��睰��C��J�BI�[�
.T]15�)=Bm�Y�F3�J���1d�rg+��g���aqr'ZwcBSt
�M7T2¥%r��T�ʈ���4(���"�ͷah�L]9%zT��e�"dRF�J3��Z�bJ��V)��.+4ª��v��u�Ϊ�=,��3]J!05J�Q.p#��%$P�M�&��M3&HT�8Qɒ�OdFXV��i�r�7,%20�&!�i��Rh"H'�#��ɢ�*�T,��V�����U��ey�Z�X7TLR+,����#M�λn�A�i*l�6��f�y(��5�0�[s򢂂IN�*T�0�t�Ԙ�4(�
[u�"�<ȯP�G����wܲ���o/U5;��:TG�JQK^�F�%{׵�[���.��ߏrX��U��X�k�+S�V���kj���ԓC�=*:_�Wm�yYB=He�YƑ�u�s4{����b�k9��7z���68��X��yAx�,�Tm��'=�v���.�cP�DmԴ����RŚs_q�&��s�w���7J.w�Tp�7Dqp*zr��ƪl\��'L��:�Qo��^��ϵ�Z*Qq�j�D���������M#�҉�����6\˸��tN��X�a:~q'C'1O���2���Q���MȦ�)x�0�U�^�͕��}����h�
�p:��)�`xK5�M��(*�_�K���+��M����z4�y��1U��'�h��(���?XD=,L�� .\]���H��)����1� �{īF�V����	�9_n��̹D�4�Ek�v�$,�G�Y�C}���+���Rተ�[�>��:㙋t��ϮtkɥZxq�\�]67Ƽ.�*,�aMԬ�<��e�k�tK�;��C/�i���u� R+A�x�� 8T5o�[���0Λ����XfϜT��PW�xpѻ��Yv�kW�-��ֵ�����}kk���z]�2#xQ��л��-�݊�
�N��{���o�t�6&k�n^���2֥F��N��x;z�
X��ޛ�mh\�+�n������+cС�ެ�ڄ0�8��G��U�r)����ֻH�s��\g쯜��IF����JVg_b�3b�2�(�T�q&9�:��#�'8l����oM�zs�:���P_(�v���u7��ڣ9|�5�,� ,�ɋ�j���u�p{��j�Wh�MZ[�O�PD���g�	M�@n��4��\�s(9.C$��T�h�{s��Oud��pQ�����rk�����{�2��/����y�P��8@7ȧ���|�h���
�C��;�i��BB��V���ev}ٳ,�d�M��yv.8�$�:�<+(xA�ퟒ
���p�x�Ӑ@�{�yQ��v��w��J�29��=.�oUҡ�����	�Hng*Jzgb�1ԥ�[���P�1��t�؍�a��_:}�����5��k*�\�� r�:�+�E���Q~�p@�l�qS��g��@�u_��W��#zs���&�gX���n܋���L����{U�'0�7G���E*fS'��_$�B��-��F��wov#����ZN�̥m�7�sk���ݩrz����ī�h�����r�;� ��Z�Wng%X��������vd;.�H�z|]�����e�&�ט+v��ڙ3dA�4�8P;B��$%J9��w;�H���a�ݒ���I�.�	,�G>����U)�F�X&�]S>'���u�Ec��l�5M�fXJzބӛ�4�9��<K���e��G����0ϔ�F�ZH��%����v���Ex6|�̝�͙��}�_+�*�7���m�ed;w� �xb�)�h��OI��-�g,�摕�48ڧu�"-�n)LP5��l}q�!��`#����fو�:�F�ɮ��9�s\�m�S2��Z�t�4n1]Aw�p�J�05rф�N�s
*��C��<�f�+Ϗ�o���_s	N���Vd_p���KuAg}㻯O�bn��ƽ1��=I�S��mk��I��	n͕B��]v\^�gޭ4T���Z���1�	�ݦ#ǧD6q�Vq�n�lA�2J�pjR0� ���ֻN`^z���b������	���TZs!�.m��M����H:�C
��o��]�=�^�q̹R�^��S�1�DV����i��C��Zv�)U����;"��RiN-GG��h��
d�0�e�7F����r�z�h:�5@C)���{y$�t�jJ#-�I5�����=��˱���E�)�2WU��a�y�g��#�=�.�2)VW "#��u˨��k*�W y��M��վ�L�F�R��!E^��Ư���{û��Ќת��Q��)R�CBڮ�A'UAL��&�����D)=�.�Mo�����>���-V�0��+�)��^ۭ��Uv�%o���g��{z��NT9��������핀��׊�{#B�Y�6�7<ok�g�J����;é����GP�<�"3��md��זg�e�W���ҹ����TDz��cУ�X�N��$��F�LwU<u��A��5+�R��DV^�k�U&Y8(b:گ���4�vc�|���%��K퉽��wo�NE���ޔh:�C\�l�\i�b+��X8�<'�f)�1�l4!|2��y�}�El/�ʼP�n�p�B�T�w�2�K�#K���p������4q����Z�a<�S���|��ܝ."�8�r��x���>~��v���.걟k��2��n;�`��x����ۋ{��k��7@kIm�N�{ڍ�H��w�����|R���+خŉ����p�f9��M�ީj��EJY#'��i,�D��h{f��Ӟ���o�nf��:j�e�!�T��~ ��Ƚ����ݎ��Sk���4�^�wn��}��Ub�V�"d�L��#��[6���w���u+�"I�1Јӕ�B�u��W
1���Z{�r;�������ִq���m�\�]���@Q�f�n�`_V�	�����ߎb��q�^̑}�j�Χ#[(�[Di�K̄����iL��L�l�I~�T2o��c��]\;%;l��"��a;�C���<��mn��k��,��~���'�Ω��/�;un#,;]�.c7+��ݲ�'�=0{!Ԡ�+d ��)�g��g|�������S4������x�咢Fv����fڲ6M��	@[�2��r�p6�����C�p^TTJ��;F��ۄ"�S�c!�WF�P�;zf-��Ju�i`��,+ʱp�����妎M��;�~ەŢ��|��bT�ɶ�tV�^�UKDc[�|qs�%X�ןw�A4�Ҹk´#�?qk�^�L�<w�h��ǭ^RZJ/�Rپ����ٕ�(�{g�9�hB�1�\(�#XD�Q�R݊�;kp��3�@���n���qS�~��É��:���Ce�1	��=�Վ���J��h��⽁������QU�V��n'f9t�@_*L��i����gr!]}�}�w��op��V��V3�Q�n�]�ju����<G�ޮ�����oA5�(^L��e_N�F�N��V=�ݬlR=��R��陸�P�򤩇�Y�O}�"�eڽ�Y�\U�
�6�U�X%sW�β�(�����yu=�h����x���6�m��kG�[\X�R�N�ZX�9��K"8������E}nSsۛ�3[�Ch���˩5T���1!]��Fڷ��йp���es�����j��ڡ�D�7
�SG�� �^o=�����?pyx�0�K�<>KON4�
��뭍�^�
2��r"�
;�M'��K���T����2�某ڇ�p������ a|]�L���A�mV����vn&1X�~x굜����E��X�q_s��j*��6A��5>s�D�=���
��jH�IL-$V̶�t)��'\4g�ڿ���7��o��t���2�y�[�Y}\��(Ly�%�A���U�1���T�y�pe�D�=� �5�I�P�s�5���ր�s]٨�k7�!� ��S
�+m�����|mGѨ�3nF�xؖg��VѾ��³�J��ě4t�,lδ�cԡ�A3Pz~���U��������j�u` ��jM5�U#��_r�d�&������5	+�U�S�k�:t�9���ᑬ�T��1Fc����ۓ��:��2��`����5%od�&r����v�9�.jf�e^�0Fu�����I[2u��N����O��]f��V�=әʔAݬ��h��J�Rٲ�����˨�ioi �h�+�ݸ��iٙF�(N}5�;�[��8���N��N6a��WP�wh�>�����׌�x�%��!�Wq�u���-0����s��9�;���U���a��<&/vPw�C���.t���ᵕb�aDv� F><=��y��@#>p3)0��(�9gZ V�a�#=�s1���y]�r(�Z��<-����В�q9����ꏹ��U`��'r�H@	��H�*��b�Y.�
�Ip��&�Z�����pd�h�g��Iu�qGg[��u�Ѹ7�[7�&̖�i$
�%jҘ�{˲��s��\t�.��^4+ZH0��vtu�%u^��P��(��ku�g�a�Y�	����ƗL�eY�n[+>v��:s��<j��u�_Sd�u3�:�fV���Ò����;(�q�(�폵Ô-;P��}�m��N��;W��0��,��H+�Y�M�+�/���ԫ�ʾ���?z�!)r�=��Ưڍ�M<�]	䖔n��vtx�\.zEѦ�I���cK��6����
��X�\In��͌��0bK��VW�䤌�����c�N밸Q��4A�+3H�SPΰ���6�إ�y��>7�dn�a����Q�%��uc�R�ǯr۝g-,��Z�n5�0r]�a�Ϧ����ψXj3���p锆�nK�']�݇e<t�u-�=aR�ĸ.�)�\8���2���[Z�'P`�n͕B��]v��]O9�m�Y7���W��i#�\��9��o����Q$�8jR7�v/�%�ʆ����7�c�Σ��-����Tr�tn��Ysl��V05ζ́�E!���5ۥ��Z�)��s��na�-�7��ѩԇnxT��<��k����.��ܴ:�\��b����$�@��T��. l��
����e*zk �CkU��ZN�2�@Ij�m�dNQˢ�ڮ<멱��6�WCx��x"��]z/�>�u�r��r�b���6�����Чh-�h2�����ܩ��4)��m��3vӷ�2��V*ī��7Pch�n,f�y]��]V�Xp&N���捵u�����V�f�B�?�����7  aB�31o�;a���eV|{��S)�K�C�m_�}9��F0g98p��
-����^���w{ɽ���t8���6e��L1�2��t��5=�
��/w��X�V�t�Z�����㈫���Y|��r9D�U�r�1延3�wRlK��
P�']mv��*����D�r���n�j������Rw�(�.(S�%�We�����@��������9�4�W�2��z���`�ټ��t�'�zZy�H3(���� �D]��2΋�T�"�]Viuaf�_V���l�u�������F�)���q�L���h
��q�=HN����6>E*�c�w�5���Y'w]刭<ջ����с��vd�(���|�¸ۤ��WpY���?r5�<&�l�fd�ߣ.l	����t���u�u3K(c$�4t��q��w|f��,zN"��{��"j��F�%���˘c��rm<w#-�#5�u*�=��z�m���U2JS�����<����Q���� V≋���S(��Ot�6���Of�b��J_��t�2ytп��C�#,0����.��ڲ�H��_A��R�u�[�wN굔�QY8�%[�٧H�rk�\b�z�w�\�/�z���2\�ʄ`.�B���6�_5G �qDE�?n�"��'(v����lׅ���\+_y�_��K�q�GN98��tz�Ag��>&�i�$u(9%�
��!y�þ���s����ώ����;� ܩ��6��}�̩�V�xw�^^�u�s�B5�m� ���0�8�˥�L��_'�z��9Bx�n�Z06-S+�o*x����^R�:q��he�n�F���o�����Po&��b�I�Y�2*t� �:�����Г�[�+�yӂn�J� l��7J.F���]��Hq\*zpyF��ҲP�I�]z��7�Z7����{�ٿ�m�Șxc��G�;�=qY��� ����驇�}����4^F�{�R�0��S�~���'/��`WѸ�C�w^������܋�
�"Ɔ�R�}�wK�L���l�Ѕn��N̦�����ʓ2:��M�*̢�����ҠFK����_�������ɭ��Q)����6X�5Z���.�}��Fg9�f����g>Z��wԄuϞ�1}{��r��N���+�Ζ*�5B枩�l[-q��������Oaz~ae�;��\:Tƚ���11�N�L�!��}�c���������J����v*F8:�ƃf��ڕ�9�C/����r;�CI3�lEb�����"Z��TP��-Ԩ���̰<1g8����UZ�E7_��ca�v��r4�8��NaKLLĩ=�:���*]������� o$\I������a؝p�[UU�Y-{��u�|�Y����G�0oHZtm$�,rX��ŋ:nld�2VI�j����:�ݕ��_G�%���e��o��+{2�v-Jkb�P9���'�q�z,L�j�b_���1 �!��#6be}����)K�v��ƺu���Cw�J@�{��dl�j[R�j!v�%�۩�a���Ф̔��>���Zj=����)<�p.5и;�.�gd�h������ł�g.Ӿ�5S���0��B��՜Q6���6�K$��T�����z���^�����*ή�'(:�I��j-����G
�Rq��HA�d�תl����H-\!Px;r�6���h���hR�8��z���U�+��4��q&(J��Yn�̔����v�2/�a_R���$��[�ŻDa�.e�os4&���t�]�nѨ��R��Lw�,Q��c�W�y�Ǔ5L�g
uɁ��T���T�ˎ2��ӧ��q{]�`]��,�(o����'g�����=�Zк��Շw��sSQ�1�t�X�~Ү����С�K��V�;5W9��^×���mh�|��$ʏ��n��d��Z-ݾ�>ֶd]/�%5N5|v�c[�(�/	������_K[YCrgi  *\�Q����']˫����09ݱ&N�k;t�S����-ZFv[�Ms �]�%m�/l�vA�:�&�B�ٖ�=��tiV�b��Z��f`�k���>�Ѣ't�vն���"�� e.�1���W��5ev^��kG6�h�ǹ��e��TXÆ�Z��]$�W���v�U.���\���l��P�:�`L�n:�ڎZڷ�WWl%\KG�;�c������7���s� �.�bh�s��M�[�Tc�/tM�]�>3��z����>���B�Ab� q^N����6��e c2nO���f��
�T�+*]2���|Н;)���Wx^�6�[Z'�yڃ7Kй�H�y]wpXu���I� �g";O��^���|5��Y���]oݾ��B�"�@1ܷ��T=]��]�ǯz�ﱆZ�m��`:��(z6�:f�����V$�v��n�79��ڹm$h�H�x/.��u�Nt�'��m�q�b��y�v�U��D]�8]��:�ΙM��Z��@\b�^����S�L�3��U�W�+�*��u��st��qk�T�v��m��"���������ڴ��+����sj�p4�S����6T=��:K-�S3�}�\ L��n�*��U�f8��o
X�;;�[{[]�jS\U0�"�����m�t<z���\nt��4�t}��5\'���JU��U��_k���x�]1wGX�#ô\6���Yt���`D1��9�=�^���n�2�yu�2f�k���0�D�.�k����j�k�3��ob�$�L떔��F6��͝;�on��ܺ���z�אE�������sۚPj���qfl� v��B�ӣ��G���)���Hi'9���GS�fFeU��dH�TI�$��Q-�4
#4M+3\�W0�'II�%Ғ#�\�5�@����\�H�4�L�K,�S.�S32�s+�$�B%+sS#-�m<�����DBM3Q�2��,���5Ԕ�Ha�	�zfj��F(�	�[�j�&*Q������&"I�yy�UV�^G��E�^��(����Q�Z(^zd�irnȝ"2$R)]ITдʰ�2S4����T�#�)=%�U%$�P�E���4M$�JU,(�]<�$*����"�\�U\�].�%R�r�R+ЊA,-��2�3s\��=TSJ=2�����$�D�2�T�At�H�Q��@2��P��UT*�ED���+\<��CQJ$M#)43��mb)�ZUn�D���y�Z��Bf$��S���(JY�\k�AD�����/c�J\�"��m	w[Q9�[y�8W����p�h}p@&���ki����Yq+A�b�k37�j�5z}��k�"1&���!��S���2(I�����'���p�2	�C~Q�E��"I#LB��(	"�8�nw��f!����b8���@�ϼ���[��W��tnϱ���? Y�d2H���$G��b��� Q�1	(��?� �'�p���y{�ǒ�����Da�mǄ�`QC"=�`I�#�F�(����	&>"BN�f��ט*Rb��޼��{�@� @}�Rr�Ov{��o���u�����'~Bz{�t���$�HI=��_?c�!�����x@��</��I�S�g�vCL	$�����"�D*@,Mm�Ư�q?_��k��߷��a�,� a�f�@�0�1���Ɛ<DI�����"H�nu���f�C>���0'�>?�e�q����	���쾮�9��RDɘ�"H���I q<|���逬��f����F0�""��R���I�EԈ�|DiR�j �����ޘ�<Dc���G� 2 /�w(��<!�����#����}���#�3 xjf>��� �;� d�9��>���B1
P��$���W�����1�n{��'��$�d2H3	"8���#�5!Z��B��U��,�Ŏߦ"�Ř&8Ł�0(� !b�s��Y�"��Ӻu�s�q�1P����<`IDx�������=���xN{�ǊϷ�hd���Ǆ����vCͰ}L����Y�E@F�Z2��0"> "=�f#���1$z�)��`೷��US�����8�<|Y�L}�I�1��0�c0$� �G����G����{!���8^��������yN{��=!�;�v�o�ߐ��D�#���|�'gog������#�ȉ "��"I���g�K�Dk�F>��8�Q i�P,Ǉ��������wx{+���;���߈
ץ@c��,����(�Ƙ�C�(��D`��ݽ%��!�/����7���b	��x��Ѳ�	� #|���!��Eo�$�|��F�ϭ���~{��������?���*�Ǻ{�z���z{�9�ou�c����vL�=Ȉ�?�M��}X����w=u+ע���-`����U2�w��[B��1�η���[�z��v�;7m_(��ڢ�=~.�@VY��u��J��%9�����`�-�����{�[��mr)�nN"�^��w\��f.Y��W#�Q�K�@Ke+잕�$e�ؖ���=H@F0��<�R��DI	�c�E$!�`��}��Q	ށ���|b-pzߴ���2}N���߿n~O�>��ޱ�Iǧ��������K#LC �{x�zR��>l}r������0�F$�j �H�	F �ܱ&#�b')�B:Dd� I���1@��H�#H��� ��"F�b#�G*��Ǩr�n��VUo�x��#c������ H���#�3�=����'���[�"$���� I��3���
"_��]�����=����w~z{��=�s� W�#�2!�}��gW�iW�����v{ӓ�����{'zs��A����8^��(='���C'y�PP��10ԑ ��"(�d2�� �ߔC�"���DcLB��Di��e�$��Ŀ��ޯk�ח�m�}$������F��1��b�� #�!��d�D26E�
"�Ę��`���������g������S�Ј�H�
1�!4#��c�������B�<��0�*q{�v�D} |�3���H�D@$
}�����q8�DA?�wL�,�1f!4<>��{�'|BzO��q'd��<'��;�w�3�4y{� }~��Z3���IʄfY���� }1�3�T\��zUE�����$F����BŁ|�	1��2�=��Ő+{f<c�@f����;�w�$�o���!�?���
 !�0ȓ�D�"$�����1C1����=�%I�7[��ߣ>'���+���������{��1&!�������Ȏ1e��0&P��q�Ӳ�
1$2 Q�1����(d=~�������~}u�w���3^9�%lץ��S��O__h�Lq�v|=�2~��������{C�p���A(z�x�ȀhOH�D���x���>1Y�"�〈� #�"��#�@$G�w}1#Ԅc�9�1	(�2D�Gsk�k>{�ȟ���r�1f!$"K#��&,�" Q��F$�&��!���`24�Ĭ�"1�i��,a�C�~N��x��x������$���=���H�{��~7z{�'~Bxz�~�$&����8��vL̀��oOVy�_WkKglf=����"o�����qE��pv����-�A�����)}�q��ҽhv���Âs��r(Y�۳X�!�'e��b]3�ǫd�O��x�ɝ�̂h��s���Ʈv�gVb
�V�=};gv���}���P>���F#���>�	�1���G��<</y{�<��I�<�xx������S&C��ޣ��~{'���?��p������=��g����Г��1��<>o�C$f6խ��h��@d}{��� ��aL�G��2DI;�(���G�t����eY0<�^��I���0�g���z��	�P��f4� Ȏ1�����6�c�}3�L�~ʦL�[�����Q�R���x�ȼ� �LA �'�� x��}N(���~1�f���_(��{�@�	$i�m� 
H��d���5�>"Hf"�1~��W��F�q}�}�^)�^��#�`�}		"I0",�	Rx�QЀ��0�JQ"H��I�1	!|1��1���������u���~O�c��C"1dabH�H��N���G��F��^ޕ�k-�=C��sǄ3����N_��?k�{������P��g�~��{����B1_!�`I�1�8�?��`��|��ۅ?'������vN����0����U��x�M)o/-��?Er�C�NC�S'
?�z{����x��+Ą��S��w�7�ǻ� ���$��4��|߈��Q'�G��+���|G�a�F=HM]�M{܏�{�垀H�b,�1�>�
"|�0�}��& $G�0��P(���q=��\z|<g�&{�==��&x�ק'
��)�G���N�{�ցF8�����H�	��t)fk��?a�g+�{krw�x�ȀI!W�D�����G׻+��?{��(I���q���DD���
"�0":�|��7˃��/Ou]ߟ��<���q�I $8ɂc��"2���sH���)]enn��A"7�Ƙ��mz�c��u��#��	�#�?LF�4����Ēc�!00�ﾑR����w�	=��]�n��d�	�3��F '�T@d#���}�s���k�'�]ö~@��"#�C�ƌ`w��xN���<~x��_pw�|L�W�"+P��i��(����8�3c���XI0,��
|� Q�G��(�?�@B�9���xH.W�@�A?�P�)rզ��C�^0�WP�j��kzP�
�<�j�o��PN�6�ݱ3*@�W�o]���i5��+/@�WW.Zk7@Aa��u�
��=�q����`ݔi�	�W)�sx<��c&Q��L�����|����Wo�`i�fL~���DM���;! z<F�}{�'�����z��S��~z{��Gd��_�ｿ|��^Da��tD|@\�GC��Dq��|C0,6�08�`3�{��k��\�%u)ϻg�� LA �l	#HD7y�wx{����L�/|�p����/��c��GxC=��ݾ�ǻ+�c3X@B#��s�b�=��!�`@Y=�����ng��3���l�,����v�>X�L|bQx�6��������ϗ���*�;�=�����8�����l~N��S���i�Da���p$��${1� ����O�ZŚco��g�o~b0�0�c��鈯(�ȏB��a���9"> "���W� Sޞ�]A����zC�˼'~L���J��)�S�2y4{N��8��G�!� af#��ݽ�|����,�w�����Y� Y�cLq���$��Z�$�����
"��@�Ę�Dq�#L��c��"'Tw�#�w�$�G�7����<=�;�i@��b4�"Z�#�PxM_3�Ҥyeu=�S�����F$� "K#�H� /!�]SDif1�2/u�$���3ѹ���� LG6� |E���c����"0�G�V�a�G �#�!4#�goM��}��v�g�gC���� �b&0�H�"0�LYf,�"#Ig�"HpΞK������P���:�G����c��n&��U��\�����Mzm��i�.�c� �Ŧbiϕ/d�5�4�Y�����o֍�S�:�3-q��H�s�ҙ�^8�+������U�.ڄ≴6�����s�G���x�S����Q˗��5��<�y`WO�N9��2�Y�Qq'�w��\��k��_P9&��R�����G��jl&��s�v����<s��h�n���H��!��ST��h��5�x� 	�r��ll��HA�nvq1�vQɨp�V�^ 9����	|�`HL�JWsܜ��� ����*]c���W���۾۵Ӫ��Ͼ���0����a��2k�A���}�Y���zP�7Z:�N����Gz����q�ֵ3|���tƇN`3P4&�R�Ǚ�/�?!��θ@
ElEb�-כ�i$ǰ�v�MK����2���V��Su�-�.�i�#J�8��:6o$�TYx<z�k<C�Z�6;�e���o;[_d�]얮}���kδH��ki�3����ֺɗ������C�� w0��:rU�0��j�{B��6x�Z%}���9��9�{&ia�iU����]<���(�R;�l��u(.C&
��0vH��m:7�\�z�{/j�Nm��3����-*�&�u���D!@b�֜�ԡ�Q�R��q;��N;;�SX5:�<(H�r��\�7���m����&�&�p�o�OG�\P�dkL��5+:2�oplW��-�5�~v�'��م�U]BI�q��~rjJ�	�م��^�f��Zcq�S�1��=�w�w0���F�t���A�a��O��WOm��}���ِ�\��@m^.��/iRz6*̱�QyJ�W9̾�5��F)!nn�U��1.c�Y������{ըt7��M�7Ǜ��b�귊�y�\s&�v���w��T�zq�V�P���H����O�p�9KwO�K���K9�"�������DDo�{$���鼃��wM���%wI�0W���:�:����V�o��Sr'u�3�PF��'Cc=&�
?{�m��~~i�����>��Ť���X��m@�ޙ�=���@p��vH�W0�L����s�R��S�M�'��%�7�j{��:�z�R^q)���v�kʦ��̠��Y5�9L�ߞ_�uÞ�p꥖7�{ t����~�6���z�oh�&l;�uJ�.+�b�:�\it���eal�y|���"t�Ɖάjm��{���� �hA��H,��1Q�]t�_en��_jv���������zy�*
�j�w���L�<~a���BzK ��l�ccu{e�Ϻ���T�����@�(v����1trY�=iR��0�)��@�Z�Ƙ����7�2�>
�����;�uu�+&�X��K�ێ]>;��p�^�"��/u��F"N����Cz��������rT2�N�?o�\k�I�D3�)�Vۭ��(�W5)�K�Ӻ������L�t辷�V�΄� �!�ǒ�kPӶ�ow���v��Q��҇%�t��̲���:1��gNw���r�hMN�Z��pt�'F�|ڱcw���5(��י�Bu,ߵ<�!�_`ל����${���8�����lߒ�{���꯫�>ʎ��q�spN#Υ��vJf��<Lg.�+#y�<O)� ����[f����4��%R�f�����ʠO���adV���mP��g�s�-	���R�w0/�G
�8����ݹ�ݛ��)4�-q:�Z�>���ub�/Yzpp�Y�}�wzF7p��������`��~�m�K�ωj`n������K$1�P]ډ��$&���H}n��́��V��P�f�^�UK&�dΈk]k��X:S4��
vx�`��0�:�k�k[�lu��������S�i��l��V��rW�{���S#��ʈ��p6hg@d���	a�
1����iD����1�T>�T�dࡈ�j�ގ��B��w�SN�%l��&u�$#g����m@o%xԾ���-�'jԎ"Fs�\W�z{�x)�=l��HKZ`��o|q'�[���C��V��tW�XP�RX��TY�Յ����T[�HD�o{;Q+xūU&�oc.h��L%eM5���c����<oW��0}�U���vA�{��y-X��!1�r��`���Ќ��橯4$���[[wWi]:��n��h��45
	�Լ��k��Y��ha#��)�h�^��O�H%���>��0�Mpd�ǃGQ�Lc�J�i�I�� η.U��b���9Z.՛�Ϟ4��ʴ�E� ��z�.�{Y���wD��@X�|��86(�.8�J�3>0�n�+A��Ffӵu�,�C�'8��ǾР�Gv�=��Y~@u��kC%ss��� =���g�.YK:y���M;�tx?R��p*���&X�!�c��@�V�E�4�ҙ}��e��.��EEk�J%�t���P��!�kWȔ�ޔ�&,oͺ���Ơ�ҁ��joa�WK�ѻeI�^���D*G{S���/������r�a-�,�	ڞ޵2Y˵�i���q���ce�MDt�v	�x�!!�<��=�&����L�	>��w�������'��<Jq�^Qd���1jW �v�ޑ!�M��]1��f��f�Z�����结��ɶ|2Utn2��4�.ho���O�,��X���6��󶌺~Q��-,�5��oqe�e���Ɗ�̨W���\�X�ҋ���Cy�PqK��wT��U��;z��s�-z��|��Y3�%wJg��}�)�zb���W:�:���4�n[K}�"#S^Zpʃ�s�@�j�O v��cE���m�5b{���Wv���g���G&��`�\;D�����Q0��.�dYz ���E���}�.b�_�t)���-�Jva�E��_�瀛HWQGP9[�f�:�c�珮����R$Ng� ���u�;Z���a�c* �d�rrO������@Wۍd1�����;.u7=N�����/�'k�&(Ø��U�Z2��W��P�7T�0<%Y�M��(9���"�L〺�K�v�NV���:�4�,��,9�}8��/������v.1�t�<f���&���h����
�E_.���O?
���5[�nF�ȸ����ѕ_r�Jն�ޕ��mV��Ip0p:q*�]��ӣ���H�t��ț�9@�H8ť%m����۽�h\�`Ω�څj���)��6dNjV��9�9��6�u� R(�]��f+��� �ˤ|�o3�?��x"p�K�gju�R?b��{�n�5�l��mk���s��q��g�Gss:��2^a\�Y�\l�&Z�89��(����y��μ"c���FD��楍�"n�o��ʨ6���x�S�>��&�Z�'M�g�`#���0y��]s�5���zfA�]h,��uj�GT���uZ�n�134ۭۨ�0Y��~H��"bVӣ�i�yx->��:*2>���6lW�:�z�x(��S��\S�[�̼�K�-19
��7��˚ܾ��c��I�HvrIWWU��b,���ݚ:�J�vv�􂛶E4���Q��V��{c�h6q��w�e�m�}���k�~�"��n�fo=����W�ј��*�%7<A� h������S����w�,�S�>�Zx�WtedJ+�i�z����}��4�t�އ�mT��d�&����9ú��b�$GWS3��o�;(^���R�V)��6��Km�͘ZuU�-�'v�c��ɨy(N��H}<���Bq麔�-��/�=��P�	�Hnx���/��!qv��y���g��Q�x矶�n�z1��:1lC]x���=�j����B����\~ܯ1�c���(z����-���P{ֳs�VLXhΝfq��bᩡ�o-|���BJ�\Nd������5��m�ܴ��ngfjY�9��41i'�2�6K?Z�֕p���t^��Q>*��-՚ޢ���wu�����-����7�)�H�l�
�%�MG9L��h�놽��U�yE����S	Ծy#V]FL�{�4I�Q85��2do����@�����z]0C�g�n[+�����(J%���5��G�f� ����l�&�ZF�o&yX���OPez���T����}T�_����%��ng[���W�
޺%���%��<�P��ܝ'P,x[�/�g�Zue���̗�Bٕ�3n�c�	íФ+4k�/���X{��_XB���]sj�	:s_p`���YWl�#��8QK���՗��nE��7Ae�k2��\���Ƅ(A̘�n����l�v���F��Cr����z%����D5�����޾��)G����+q�Ե�[�BC\87&��#��qr���K�r�Z�oe�����U���zN�E��!�{���`WC�۹��d)r���QT�|����n%y��ڳ�a�g�j�0�=[�uJ��{X�m��Z�)$5����J��lֵi1��:X�d�B��vZj�EЃ�R�����\lWq���52����XA��6�\IVm�&WM-p�zX�āY�Z�dCY+y�D@T�,xE5:�5fgt��=���XCKZsD4�
�3�u�;Ք�=k�yKb�]nEb:��i�'%뿁M=�G-`��c��%t]-��d��k��fN���d���K�W�ǎ��[��t��KQZ]���yN%��kj�X����*�w�BG��b�,����v�fVs�w4EY�8���C4�|yk�]�,�|���Z���h�>�W�!�|�v����W�֎�c,�9.YSp�Ɲ����W����ݻ���Utu�WG��
JD�/�{J�����]��Z�r嵶�k��,��GF��+AŅ���3��a��,�u���_4�L�*��G_>��kW[�٢����ZZqX���iK]Q�e��˰�&�K�t���2�[��p��9��I�Tg3�5�������r�a���˻H\�]�_Ho�]\]LkT�Z)sDx���W6
���/H�����4;xT�B�WPҺ����i�Ps��q�3�N�N�ܭ,�U�(�r�ERTd�����k�u5����uBd1�@(�)Q�J��~+��t��Ku�B}{�� �Y5��G��g�0����yx%��X�/�m�X��1��c���̲[ݮ�=WBĠs�Ǐ��Z�8[��Gz�nղP�7�5Q#����w4�Ģ1]
&�����&��4�}�ۦ��t�T.ԫ��Yef�F=��V�J��ѷ�����y7� �`�-Z���1�`e�܋V^�K����  ��9].÷]q����;��g}���%�L��]��C�����y�A
	i��j���#"�B��IT;aw"{�a�GPB7j�`�+b���
��E��0V	e����r[)��8E�<���e��<=G���gR�ę�%���Z�����G�\i�\���փ/0o"�2�I��s^uY�Sf,��2��LӃ�^��2�d!sf��*�5�R5�rڦ+���CzN�҆c�2��B>[��,v��a�ʵ2�,r�Ú$�Ww�'��ח��TV�aXy�$�B���������W���TW�[�j��aEh��yUV�-��2�۫��ʽ0�X�f�	�nFf	Q��en[�EbeEXJb�b���IE.K�Ba$��-��0��"MJ�BW2Ԉ�CO��R�r��WvPH�F��yI�)�g�Hd��F(fUI	V����ey"f��*"!ZAT��*H^.�Z*jD�Z��I�=��2��=7P�*-�Rr�B"���+Ƚ�Y��jf��dYj�!(Tnia(F�+��&�&T&�Z��UU�����xF��$���X�cD*0�3r��=5O0�Ip���C-52C�J��2���"S�P�=S*Dʕ
��"ȫ,�75,�]$�S7L���F�YF�b(�(�b.R'���Z�f�����Rafe�Q%Q��P�:"�Z&n�"EՐ��)�q-%Mك9�СV�O���j�dG{��:�vP���'
�������[5붼/E[��D �����~ #�k��_���G�;ep
���Bl�$qT�}�p���v�su��D�X�]}#����cI���85
�B�mj�`v4Ɩ��T��[�d�<�bw��꭭Iv��ݪ�o�n�u/�t&�i3ب�~o�|��Ʈ���ʋZ�2�Õќ��w�L�^��~�5��}I:H�:!���+�����2J�t�+��2w�9
B���ݬ @6xGI\pf��3zx�ʎ]n�f8C
�d�S`GEtʱy�+n}S����cI(C�w�v��q�B���T�K=\��B@�ޥ+sp]�[]�a��,�AK�y���UTTr��	��煯��>��.�V'���8]��n���=�b�i�v�꜡c@M��|KS��bo�YV�,�|��Wj,?b@Ýu�bW�pԹb��dmz7�1�HA���ʩ�����d:�MBs+��DTaD�@69��0�s�Ɵ'�8�b)TS�8�yخ�$�b�H�V�Tͧ_4n��ˏ�z+�0E�GKd��-!�F��̬x(;�^��!��!Y�"���\�HoD��8�y(?y�㾮�͒Td��t�0M[���:��m�|� �݁�r��9@����|2^��be�\[�)�����.fٗƕ�o�wƳY��պ�9���.������>�"""���*�7Y�}�qYU��[%�����j��L�^��Ͻ��f&+qX��������ק�*��I�{�[	}��6-�a���2�Z&�g�@�t���ܓ��v�T�jp�b1I�c1_a�p�@�!�B�҅�*KS��+4���9��n��R4m�|�KV�����g��p�YSMvĸ�4b��x���xޯ+�l|�n��jvfا��J�oJW�#x1���'n��:�j�Y��N-Il�c�A\�;�^��㔺n���J]ݩ~��U���?����!��� ��ީ7�Ƃ���I�u��>�f�e�#]v���!�1���V7�}I����;��\��"�#^:�{iQ�|'�Lꩣ/q �� �:\�q)W¾�)�# !�kWϥ;l�|M�H�9���k.����6zzp�ܫ��{U�GRe�� �E�r}[#��j|z�v(��]l!s <p���X6G��Tp���m�ƽ���s��E琐՟"�]���5���U�;�v�b={�8$��ĳ7 �����>��x9�Ѽ�P���>�^w�V˧
~6�圿zTdL�O���`����it��f^�;��`�=ہd-'`vq�˩VsEv��&Y�2��%+��q��=/�x�PT@R��K�֮�k@��#}z���  
�U�w_�V�����D�ݞK�y�7̑$�oHD8ũ\��a�Q��k����0�cOj29�o�����6����Utc�����X���'��� ������V�:X��w�:<��WY�f��tÆ
כ�	U��z��^�Ba蔍Σ�!nI��U�t���Q�u8}=/���ҙ�_"a�Juq��D��-.�Q�D�t?wa�{�(�#P`U��^��t�������7*��/�p�:�p�^J��� ��뻝|�GHz�1���ת��	ƀ��U�P�i�Vo�k�����{$#<��r����mV
����]6w>�_f�Y:*3r�T�K��.�6m񖫬T��>|e���Cv��,�����c�"�ܮ�ψ��Λ��1�-�z���Hk9	6�E�O�MT���ћ]��ja��`6m*��]=9��=�lJ�쉺���Z2��ܾ�c7��Fv���@I�2���κ�a��S�lȜ�R����x��g���V�"���A1^8��GQ�z�N��*����4m��f'Yԧ.����n�'�<|��pzd��sqP���G�I�`iY���-��D�u��2{��Ӊ9Z��6�6�-�ʺ�5mu<S�\�X���Z���a�Y���j�D�im����U��Toh=x�۴��
O��(	����锏ئq�n~/���㞻H�V)�<˷a�`��혓��dw��zq�#dkT�D�h��������-���F
�	��S��Ϸ3ݷ8�8�[�~Ә�����<�u8�A�
�:rUe1���W�3�&}��.UJ\�p�	>�4RmZ�n�0�Pd�� V�%�,�T�F���xkGC��_o��>���{��Z5�Ò��?�� �a~UJS��R�<=Z�^�=�f��Ֆ3v�����npP���=�+��}6�$r��M��͋��#"�<!e:��F��Q���5Zu3kE1�mm����'���KMDj��I:�0�����X�S��MЙ��ǧl1U�y2ȗ�a�*�e���*���^�a��xMJ���ұ1c�_��������OM�Ss.
����ޭ�&c;���ZԮ�'�^�BX�RH�9:�6��ʌ��-7�֌����p����'\�4df���m�H��D���aa�-TC�C�cUi���14/w�7΀�-|���_���*X�p6�>L�ø8T|n���,mq\�63m_@�]�v9�hY�����J� R9�^�*�s�2�g��&d�kv�><v��֣])[�k1�G
��׳[�/���[�y��+I��"�M�r�iV��v���=����""���֜��lH��3���I ���y#�6M�}}�W����peLV�6x�Y�r��eS�y�/ ͗�����GW6t�Ϟ����̸
�%�MG9L�ח�nxF�è�J0vmf��hs�F��0�WI�\�C�+= �gh���*sd�&=�1�\�z��ۖʉ۲�]�Y���Fu=���>�b��: �H;�P �<oc�l�0^w����޴k�;xC�K{Dt�����m\>�6��(G������G	�WP]d�b�j�:bԍǸ��*�!�9:0ZYMȎƼ��1�yk�6�5�`��b[��ܕ|E�� x�
O���
�"�������T�+��8q*��/�pW�O� 4`ǌ^�-CH���nh|�
�`�3-��~�=�.5�$�#�Έl��r��hpAS�VY�<��Kfv%���'0�5/M� 	Q�+���ҙ����r�tS1�EͲ^�cC۽{ ��ʚM�H��)���	��@����8�&�e�P/ڡ{��r��	t��<�g��{Y��l{��%���P_�$�w�X�}��[��6���h�:�kp�/:��6J镜�|�բߌ��<�*V5�����Gt[�ܲ�E�-%qF;�wW.�{�]�ЪS�W���خt0��vt�W����S��6=�F��"" 	��-�qv��h�;f#U�U]'8�:�Z�>��R�ubU[��.�j���w �_v�v9��`kz��,3I���s��K*E�K$��ʂ��L>y�Lc�6*I�mjY9r#��Z.VK���*Wg��{u�P.�ʘu�4)��m�0o�^��}8��]���7"]=��)c�xױ�*u������.+�bm���]�/��3�bfC��K�zX0׾&B�:�l�v�_4���x�"b������,�5��W���yY7
2�NO�b��gD�0�F�8r�eH-�%�^>��{���R8������5�bʌ�la�t^���4S4�fMw��Y��b�+���+>s��t��i��@�x}���As�>�F�Br����pk��]�(�E H�o&�N�s8���7�뗢���a�@�G��0����p�k���C/ ��N�zn&�GE�8�J����`��<|�Z������鬶T���d=?iJ����co ��ީ9�����m�ef<~a����[�Θ��]�{Z�R����
dZ�V�eY���Woc}Y �w��>(�;�5�|hs�O���|��K(s�u��X-�j���y�͓WEћ���@��6u�͚��)ʦK�X��E�>Y~���!�Z=fs�xo�5�渖q�"m��'ذ	���|{�&�)�#\<w#*�U�rsC	�YS޻�꼴�Se����Zѧ�0f̦P�������z%;l�A7�"�R�{lnn)ys�oU���5�ɭ���[��)q�m����&��G�����P�.�<�����;�öo�{��TKh��c^�s��W@�3��C�Y�i΂�W��8��V_ҷ2��wDá�{�C�=G�j�/ 9`k�"��^tE-<N0P�0��[ќ�V��6.K�Ts��C%�n�!��6����@B����eX���'��ŖGuLS���jPj_���h��a�k{[�r@�ߒ��Q�8!_'w�s�t��~��'5ֱtۣ*쪭F��kRw�P���9딇����o@ _I��j3���zb��⹔N�`�pQ�Ⱦ�'+9�]�>��Q�,5��Fq�ʜ��D���Τ}��Cz�,��tEF!�]�'0pҺ����E��n*��
��k
K����<8���\��_��yvL`y3��71�p̳L��G��g:x�Τ�c��._Ay�(�Iv��|���vKl��jʜ��'��*v���x��]����Lbk-�"ذq��mef��.�Y�#�{L�➤����
F3��4=�Y��"zf�u��{t�'ﵳ�e��=���g��{~L��9�o�Q-Y��I:!e8���S��c%_gs��%�gP�*����-�n{~�\FT>�<s�?Le�gާ�+Y�8�Cc�ɓУ��G*����}P�aI��@,�%w����u�����*c���GR�r�-A���u�:��;^��G��L7İw$u��C���`�=�K����^�!��>�?!�Zܩ�qowUː�,¹�͌	�v�:I(	<��i��׊�Y�������V�q�����W�pU����i�8��P��B��00"s$ҋ���Hȶ�ݝxAR�*�k��+'79Řq;����eNn��}Aڠ_(cP:�"�� �v��[�W,GE
���q	�T�Τi��ƣz�\��&���"a���m��� �7V�w{;�CǾ�4*Ά��rU�Z=\���Ѩ˄��M����4BB�Rd͔WNɷ��K.J���Ԓ��!s���_Ƈ#�ozWOk��D��d�&�����Z�3Ə�Ӳ&�[cu���;�.:6���r��m]�ߎ2C�,����	��3;k� ��I���t �v�|,��ש=Hq����N��F�"�%�t�ώށ�ʠ���]�{��=h��E�P�x���}Jn��ˡ��33.�zqe�|�7�v`�c	3��,F,*��?Te-�5<�c_k�w��Rֵ�oC����K�+gtV~����x��hpy@�Ws*�*�U��0]=��a��FLђ�NFpkU�s(X��;�:�ϵ����ʳg��@�� ����B�y���*�	�k�+����z�Q���e����9�P�M��8q]R�Pǩ]�SX����*�$�M:����L��x���<���&��ضnU�F��e�������&t��1>�u�`X�2���u��7�t�4of\d�ɮr�|�cS��b�@3!&2���G��<Q�ȓH��X:VF��J|�����K��+
�.5�@�ۃ+�s���K��-����4+X�Ѕ�>DtW ��������<W���{g��� dI�Mn_�n��Ң�Gi5p��?T@�82Oa��s��L�Ds�,]�\����HqJ�[�u]n�	*X�me4c>}'_�c��˕v���]@v�\��������Y2X�]gT`zH-�mnshni�����֘�� �ѓ~�x��L6�W'�,e�Q����؀�[�x��;��C4�w6i�1}��ͮ��h�պͨ1=ٸ�XE�T���>u(����Z}׵��ʱ���ǣ��K��'q�m^\�� ���z�k��K�H�{2��b}Q=-�p��؄�=���U��'\�峦�uw4��O�w�5�i6ay6UZy���qx�n*����.pCg!�Vp۾����.U�3�O�s��I-��K�U	P����+���ҙ����W.�E3!��z�h�^�	�G����ޫ��9����&�u�X�ȭY�,^=�z�Hs�)<9�o+�X�ʽ�ծ8��&�%J�����ď}�Ҙũd�8�@�=���|���F���B::U�bk4�9�]���n�2�@IG9��_�卧�R҂C�Aȸ���b������%��\��;��2�X�2�,r�n���_'1C��D\aD�3;z��h���H�h����QӒ��S#qL�V��L�u�F������^�'��?q����ɾ����!Y@ُ|OR��ǟ��r�rZ��+;hw�\�&LH�t��;qQ�&�]�Q��O�����U�t+a����q.D����6'�uӑ�(�a�1E�
���-0yS��\�|�wu�;�ݽ�SrK5�,�;t7��)�'j�"��:E�49�ec�-倎]�<GU�4�ehF�v͠@.J��cfí|�zC�jĔ�C�Ez�$V��-Xﱍ��{׀�ԛ�,����=hi�.�E���=0��\pL^����q�Q�J�zT�&�q@{+�pewdצQmp�
8e)c�j�/�Q���j�z�W;؆ɮe�6����>D[�<<�	��mi�EY�Ppso9�]J��7+�v��C%6+'ǭtY���`�.���#f�G}R��d��	u��Ѯ������Ǖ��qtQ��̋qu��*]U���`��lݼ|�
�5�Aj�лv�,Ȝ��y�n��g���4i^�3))\"���=F6��6�Ӱb3�S�5l8�1�0
���ǚ�k�2��2{n�ڜ�l#ݭh��k�U֭e�|�%��wQCh=U�@<W'׻��Wʻp�e�>��{�l�#�7'��$����t=�`7������+n��}l�����L|)^���h�uGЮ���hvf?�k���Uk���X�+&ΡY���{)�{��qJ�GwJ��:%*	�$
G��Qd�m""��:XQ��U��pcs��.�A�ۑ�i�� o2� ���o9u6��ed����4��4Ȟ. Њ#b�}�傯l�vּc-�ד,c��[���3��WK*�T��u婃X�,������QC��4��i�쫠NQ䙡Œ�":9 U��j���4���*������hw�[ڱP�}i1�h^�uչE�`b��Z���׈:z��(jMf�\��o^�gpG��Z��4dV6�Nu۩u*�#Ѫ�r���#��{ ��j��j�,1]j�M����_�s-El�����ֳuw0��h��+a��W����d������2��g*"�N*��2>��>jf���9}nWM5{�kl�2���¹ r����!zP姹'�^�7l9��7���\�j�k�v�����h[�Z�Ʀ����E
WkY���TB���ޅ����Se(6d'��L;�&���w�x�iNy���ɒ:�X�\�4m�m���U�
y*^,#xӲ�*�.�J1��C�Nn�.-]����hwV+8��kF�˹��Ds�sY�9R�;q�;�8�qc��CխEI ^�i��oq�����ppӔBΌ�E�Ff�6�0�;oXvK�gT�sv��}�S�,���+F�/V|0�;ow��Dqye�o^�f�q���2�O���������f�b#y�k��![����{x��F5�����ݽ�5.�~�{I���lzc��Vb�-�y�*1��y��+i9�V���N�|�bg^Z�Y�A��3��Z�LA����Z�#��^�y�o>�>�w��,��$����4�C�P��"<�7t��yv�TDda����Z�j�DXi�UE�^�aX�HE�%�yY$�EV���F���H�nJaW���!I�W��R��F%K���慢�%�&�E��F�6(bA(�$�W��z�g���C\��St4#D����t��LQu7U�=<�$�OSp�\���		̵��T�ńQ*�������"ZzQ�YbY�b�T��eV�����9��
�a66Q×]#t�0��"����)��m��!F���|[��Ǎ��M�	UFq�hD���h�Q�p��g�OMSM0�P�J;b�����\ŶMK���e���y覉���y���ec�	�<]:�:��������[����Y'��O(�N�+;D$�A� �s3ki���K,矲wwu5{��Fwgo\�e����#N`ۣzcZw����ء*obk!�-�Z��^�}:/�@�3n���ޖ�����U���0S��6뮽����>o��,K��vWR��䊼���P���Χ��kL(]�(�Y�#d���3Ԇ�VB�̤�n�UZ�j�f�v]�iJ�B߸�z5��-F:ju���S�����Q��|��u&F«]U}n�U
�J�+���PR����/��M�ꑷw�r.�C�/%�����V��v��q,�q�����F�zw�����7�a�Ӑ���G>8Ւ:F���{X�p�<��e�#�4V�b��P��ы��d�m�軉)Ȼ���n㓹U�x�Gp��f0Esu�e�
Z�e��h��v942�G�j|{tM	3ҡ�[ڴ�?'����ڲ��m�V��֬$3��Ba�<ש�Zl��\yU�jU��1Oz�W��b��?W5L���5��PDON��2��F=d��IƤ��u�LU�=ONF���ݸB+S�cUtn2�^��[�C��i�:S}رkF\�q���:�5���vk)ɵk8�J0����^�SU��B��Cځ��8��r�Obܴ�ᕫb�gX�c�o �[�+��OQ%{x|(�ۙA�Ubͥ�ҭ��3��S��.;�H�+F�-�:IZ�S�5ok���7I?z��o� D 2U`7}�7�J~*.ƅ���[5�i��=��ݔ�n�����|���uC!��Ŗ�E�T[�Ǫ��Wh��ᲨZ��^�z�@�}&w�����W����Ӌ�U��vr{z�c���M!�n�~z��l�������[?4tx����0x����������n'P{��^/,��4o=7�H�z]����JcK�;�fp㮙�ļ�W�/;1'�{@hq�~��3!Ru�R鳹J��*΍�ʝ7g��O��
����Ȝ��{��V�ֆ�R�,����$t[���źb8���j���H\�^�`q�゙�x������Gڹ;���5�gAZ�n��������k�{pً�Ҧ95Sќ,Fi�ہ+��{�������C��M�H�J`3��jV��s���P��N�>�zY0L��?1�k�����Eb��$�#rv-=����'�`f�����b�e�:�8�;��._�Q��W�ͬ��Q���6A��L`D�H](I�<��,�����m��fk���ϡ%�B��n�3��%#�{��a����Odƹ���o���/n��b-�#4+�q>>��;�!���;$����؂&�fL������"J��c���-7H�{uhw]�}/�eks'u�.ʥF�9ņo����h�J��E��� T.�^mwv]f�w���[W��w���']Ľu�?/���@��PXMn�a,%��8�����Uu�E��0��f�V��0$��8��"bᘰ�m����H��v�iɋ��)��#�v��[��pzH����\�z�#��ƴf/a*�&�7\��E�B��o ��n��`��.��Q�Re����#Y~���U��ѽ�\o�����H>��%�{y��ڷm �V/�[3������7 �Zj�+Uq�ͮ�xA��kl���Ox����r�zv���qr[�3'��+��}�^Y�N��tzV�P��`Uc�z�Q\�I��\�W�l�BNCy��h�	��C��O�1s��,�u�ڇ��Ŭʜ7Q;������9��P����b6K�,��Z n9�9gQ��Y��SCt�nO�n�E�D�:�!G���%��i�U1�Yܯ���I|N���|���ɷ?b�iN����,+�F�֣-�'r� �OI��Jq3�j���2�N0;U[|�\�)�yv\z��uU����a?$��y���dr�3��r*uvi�VwE���Լ�ޢ��d"���[� :x���9gH�lj�V�8���<�z�yVe�*7ΈՍP.z[����]�T�zX�@���G3�׬qO.��t�z��_PM�9n���-d�_}�����pT�5��!��M�ܜ�& ��Ν�S=,P��)o8�|Q/�R5�]��v��q���G�×�>?K�aT(�o��P���^�x�"5*�^�gL�_J�Ԩ�\Fg_�\:Gǉ�������H2F��Y0��ŉ=�wUM�z�Z��#�->���Z��>�Є�i�v��R�Q�`0�׮�P��>��>���L�p��QM��[�Z�(�y�_p�O�&�[��e�>;��&���ꐝ��K�Yٝ�驝�H.r\a #�T�A�2������_rr�P\���76-��M��V����g�����j�EV$Oi|��0ǄTuJ�c�eƞ&2�u�?dd�Y�i5C��|�ƸdP��rZ5�:���|�&�u��!�$T@�{L^��8L�T�BCp���iL�ÂdÎI٢وƄ�B�x@�(���u!0�$x�/�xȾ�ʶ���sKF�4�������I�P�E��j7���?�����-�X<����s�yZW`��U�y��@�O�[�n�=�w�8�h\����'gu3�k�v���:���u���Ԭ��Ρ-ZƓ�Τ]C���n��Y�^u";�vؖ�;%���úe��8R��g7\uqMp�;l�$��V�B��>�3v[��:n�7ӕ���lϫ�Q��N��+�!vGu���VK�r��(���säQV�o1&r�Yυ>q��MYQc�XfTK[�u"i�(f���:{�bP�2��+���[]z߆���p��NT�ى�7�wb���gMb�l�'�,�X��2�[��8MV�|���SI�J�C���d��̍j_)�{l�L��a�~�jV�7�n�_i>F��\ǵ]b\gSTю�5�#s�6�ך��*����*&~�X��*+�4��	�)��@k�v��\M�5ƥ�������z�=~�ä"ۖ�d;�a����F�>L�hR��w�Vk�+n$����*v_�l|�R��8�z3\L!���[i��A��w+@��t�<�bW�9 +�z��KJ���!r.��-��Ar�+�D��/Ds��m���Zn>{�#o�p�g+�><��H6;�����,�u��N���8��CumG�h�'��\n�lq�0&b�l5Z�a���n�q�!?���OS��D8��,��Qa��������p.�-��ܖ�N�)��;z��u�5l�{���%�ݾgX�)>�ƹ�-�ȃ����=�|� a�"�F�U����FmFt)7��\��ٷԋ��
��X4�;:�L��P�VQw��r[�A7g
��w'�6����V:�8��=n�^�� ���2���n�����*�ܼ1�;��W�<��mj���f�Q��C>��Pƻ�}س�;f���F��6�p�?cK��0�����W��?)N�ҹ��}(-�O�&pǂ�<vkuBGIus��\k��W!��z��ԲZX��3�����n�R�$E�Y`d]=	+�xY쨩n�Nm�1�{�Ej{lgͪ�7��@A2���ಬs����T��7���u(�?	4N�6-����~g:pwe;h�u;�i���0<�~�k[ ��BYN�f�l��K��i�J�Ƽ+B1p���5�ǻ��gx����ۑYb��S"���+�M����x�������W�s'����7*dK�w�ȝOy���3�d!���1.u����uo�yS��CD>(WR;1Fv�5���:��T���1|�3#��t�ܥ_f�����r�MKT��mY�-��Oj�� ��(T�ސ�5Cꈲ�"��T[�#�%�8���/[�)�r�AϞAJ�u�Ry���ul!ߟ0�T==%���uz������ӕ#Y�n�R»$��$��vh{�3|ln�&��n��54�|5���%]'&1w.^f��_h�\���W
�&���CEm7���sgY�9*�[X.�ۥ�~.����DDDen�-���ֲ �TXI�h����&4(J�;C��Ɵ�Yp���aw%�UI}�-�e`�7Hu�����oIg�F䷨q��)=�K�}��3��t�ڵ����]%��A�>ck�p��h��l= 2>%y�ȍ2���V����%	�[�n�ڿ���/�Z�#��i��z�*�PS�t���С���ݼ��wO�T3�c������ҶoV�������9fQ
{��v�c��S:�R6�����r����Q���M+�7��6�Cob��\p�t/g^�� ��5+���+(0��]����h�\�|���Fͱ��W:3���ʚ��t<�&b1���[�snM]sٽ庞>��R�s��݃�1|����e	n8�#3������u���D�s�F�ܡ�<�5�/��m��R�-�녮�Pq;��~�G��K���$��r�B���P�b���.�9�WiӃ��d�����ڶ���7��6~w8��R�|��ҋ-�r{ ���	v��;�v�U�$�}�,at��;��K�����S�D��V��{0�WqK���Q,T8��m.�9n��u�$��r�`�|���}U��W�|�ϼ��s�9ݿ5�Ƨ�ӟ��u?m��5�\H;K�-ޛ(�hދyP�Qⱶ�e�8���]>mL�G!>i��ݽ�vn5�J�ޝ"_>P�
�.`sUs��ILu��D��B�N��1:��9{x[���3r��VYU\Tr�}��juCW��
��-�i���pP-J��M�(i��i?���͚���/�@�<k��Ρ��ϋ�d�J��ѩ�����ھ#25���p���K���v�}�=Org�Q��lT��km^�޻�r�G$�\5k�p��M=�H�`j*�n��읪���EMhxm�AԷ��O9�Z�^7�r��B���Q׆t�����+�Z�� ��բ�4��wF'Ơ��o�<��<g�����Lb��2��Y��~�R�Q�s�z��M(u��ɬ`���Ee�g]�sʎ��7:��\V
4���]�ӱ�ӷ��Hc�[܍y�
Kv�;�sSv��X=�F2��8f�b��^��JT��v�Ⱥ�{[��<�H�.r�M���<�Afw��L�@�\�¬�]��nwH�{޶d{I���" +gϦ�=\�,���ٔB�)F��Ou.�Ϡrx��h�]O�H�jD��Ԓ���`�q�;CV���l���o�í˜������tSܽ���1�ɱ���؎i����k����D_!�kp;�Yra鱨K@�,sۢ/R���.�:������n���5��u^`:�(�]&�
�����^o�G�g%�y�)<��zp����~�2���qCO�z�t���b�gjS|S�0-:���m�D�Q���sD��WQ�� ����Z�r�p\`��p;S֖�<r���BU�~������*7B3�嫏!H���w�����5��O>>!mOZ[C�[���-�^��'}LFk�R�B�{��(���~���]�p��h�����uMYf�]���̭�v��=�S��oE�Vᬶ��uϬ����@kT�\�={�v�wg�>�zi]l��ֱy\ $�αm+�y����m;a�/&M�9��S�^ߒ�d�b��M�K�ܷ��`9U�|7�B]nl̰�󸵤�j�ԥ������ga�d)�b�D��g)kr���ZU�wuśݫ��  �K6.k�wO��U��שl��=���yxᬸ�i4�N����%X�q;��f�[
�m����l����Rޚ�)<�b�e��홞�����&�h�k�K���(t�wˤ�!&+�),S�ҟ-�S���T�-�"��m.�j9V'����(�ȅ�wgŃ-���d��c�U�:aWE��v�8�3���w�d�*g+�,�!O�)Tz`��o{����p V��gQ-�U@�}�������;A\q*Q����9�[k1�B1�&�3�wkr����}6���x��	��i���7	�c1�>��W�AY��R �n�;�/s.2�l������z!c�5��qY5��.�1�О��w�3�6R�^S�(�x���~�r�q�틀��d��Zⵝ[=���kB��> �>��zo֗⪲s��y�W�ݺ��b�j{2�f�ٕ |G�s7�I�-��~OA�耨�>��/UnV��v�=+[p����:U�Gy��d�{�Pv�s���KGf��о�]z�
Ew�*��I�/XF�ָp�����;�Գ޶���1ٹ"�ms}M�X�6��*�#��a��N�+X��ov��BM�S���a��؝������ Y8�5T���d�q
���A����ģnR�,��FS�Y�'Cܗ��Q �_i�m�����!}G����im�M֡O�z�f�	h�x��bo�˜x�����Z�]Ȳ�г���ӂ]lT�m�R��j�gƆ��㮮�.;w]̽�mW��.���Jq���ę�i�|��:�ۑ`#�Ph:�Xu�����d�����Wg�X�\�����,:5f��,s��#n���]��纭smTgb�4�!鷸]���ȵT6�,�x���9,�
ce:�y��J4I�r��Q9���C/lb+�Sz�t#J��9�ˬۜ�G
8Q�u�������\+U�s6V�w�VR�|U�ՠ��t���﷮I[Kw:�hse=�q��Y�{��\7�ܖE��ܳ�v����ǵ�1vS6y:U�l8ҩ�5JFf2��=�iI�R$uݙ�b'�;J��IB�r+�TM�W̌��$��ʛ�.�9P�so'V�w&�㗎G�2�7'F������:6�	y�\j�� ,uY�0�;�:vy��z�SW'n3Ǆp�<��(��;
S��1lhU����,�]ʴh��{�Ҥ��c���u.6ٝذ�cVo9]��5ip*���i���Jd5�v�}GJ#���ڴ����ʥe��k�����
����L[�����>��GEt�-k�y�F;9�e	X��[��C%%1�p�t����:T��f�u��eĭ��l��?n�Z�u'����h��0KnY�^Tm�cb�vͬQ��$R�]L���	�tt��.3C��n��������
�/&�2���NH��lQ��H���Yx[{��K���tm>{�&�Qyb�q[P�m�;q�d�爭il̷�X�u�e���+{�hÝ�`S�M�ũ�RTY.�5���д��(ޱ��k��;�I$�ҏ�޽@V�۝j�T�e�owIm>z๩�q��/i�gf�̵��������:A;�D�����ƓnVr$���Ele�-+ۓP����ۜ��h�|&�J��T¬����ٙ�{�����Ѩ�x�/dK��+n���[u��,�O*�Ҙ�j�N��9��5$N�*ѽ�����.�)��օ�{���l�����J�]�z+.V`���`�����Z�b��f���WqZ���˛V{T^�Jyf�sxNȕ���s;��F�sC/El��WW�����K���i�ّ�u�r��9�K���.�i�M��֔ޫ5���yD�N]&��0��>��z}+��j�8,�K@o*�N0��/�! ��N�P������"|��d������ʋ�1�"J�"[[�NT�J����XEJ�R$�byZ�����&NFW�鞢�a�E�E�a�V'��P�>w�����=>�zXXd��Qm��n�a����n�|3�zTa�(��IHZ�����!i��bdW�RPe(�^&yX���(!Qf�S9�\�<����R3Fл�n���[��Q
^�R+��Y�D���$a�E�Bfz�9J�E�i����i��z�#�*�JIW��bx�
�Xe�a���F�$a^���34#D�=��T���C�bYe�Vu/9
Vj:F�*ATyW�yMHf�D��ؒ"IdyyDx�j�jD�"�4��V�Jz����.W�¢��\I*r��$Q�I(�=��y�O3Ҩ��U,�#�5rHL�U��%w\%t��4�"�����/I/h%���h�$z������:����H�$��H�(#�]L_��S��uy,���J,�ܬWe��]ϯfk���Ci��.�:���4�^�8l�/�L��įE�������5���)�'3�N9��Cr�9ٺ�3*
s1T��'�0��-9���Z���v�{����2�/W77�����9Q�fToD
�K5o=��)�HuG�YI9�U'au�q?_$�¤�-��D�'�Y�}ݓ׸7a��'��2s�A`�g�Aj����\%q�z������nSo�%���n�2a�2��3}Ⱥ��ʨ�@l��r�ڗ5�ꀫ�F���5�b��$S�5ʪfnn�M�a��w_�މq�
(>[%'Ԩ:��K�W6�=z|�o����tا�����-y�8�Q#�;��E�j4��n�2L��a�BFܻ����\���e���q�Oʇ)T
���0f�;`hP����gN�F�oJSw���ف�V'�p[J�ո�hx�lC�e�8����(�(��MB�����sΈGU}����_�;�f�m� 3������ɩ� ���gW�8T��:m1#�]n��uwd�
@���}�gj��R^�j��ժ�9�\a�$���7-nt=iܘ�M����1I/�<v�rd#�������oS����oc��}K{��m��O��Ȝ5D@��7Cp�*{�8�_J����ek���;��F��.|�w��P��Zj�;"��,��6~:rV����؍��jzݩ'��*�+j�.V��w�	��k@�F�"c�ف}���{2�������%��Q}���O?������Z��C�jʭvn�X��%�R"u��okf��ؔ�������u�ܬw�_\B��k��nrٺ�C�l��{�З�8\�E�;�>��ku^�q�m;�L�G暜̬;�&�
�;S]ǯ���)����Φ�*$�:𨟯�y!Ы;j����G�KZ����w_��މ�d,��q��iԝP��c6{�Zu�D�L���{���7�fz���x��%�v�9V�ru@N�85=��ˌ�K�+)�a|-�W��}n�����v����'���WYc��MǂRT�����s����
8y%.*�����{�[����f�~�7u��a�NؠBͼ�.��S�5���tʃD�*S5'���-:����Ԓ�B�*�Rͩ���r��{]]��S<���Yd����h�:2r��r���������������;���lmD�F�S{����ɧ���j��߯N	�*�(���=��7^��8gv�A�Kzh���5��m<��.�LřmZywԚ�����S��{�^�k3෫�_���۟'�%�VϷ�l=�(�g��!��@���>J`0b
Z*4�y�oTb��C���a��8��6[��pU���9����*�(��%*}7Իw r{!��eU샰&�g��zu�w��|�vð�C���t6� �raJ]�$Lfn�*{q�J�ͫŎ5�龩��昚��o�O�,�:�Y��Y��]�n��E�u|��<���;�:5V+IԬp��M�ڈ�Q���M�H9�J���ۻ��ۑ-�o?EU'�X|�vz���C^�p n_g��SW<S]=.X�ڨ���+_����s�2�6�ͽa����WcQ�6�l")]{��i�de���pm�耞�d�x�����E���a����{�:�'�;d�;E�*z�b��tƽ2|]�v���u�@I���ݖ$)�[|/l�Zr�^��v�8{�U���U4Nr��fv}~5b���} @���ޚ�ݽ�fW�h�~��H�}�����*������B�>3�r��t�ֱ�:���5�t�7������{���=ih�V��b��-��LԮ�O:�6��vaLT4���^��s��{�L��S��g����(��Eý��&�.OK�Е�t�b��X�z�s�5��x��2v1���'9�o7���/��7t��@w'&d�]����vr�O/��4UI���X
��E_t������R]�2ސ���8kI�og*�M���^�i
���zbӼG*:Z�:~�I_$��I\.�w�[�,#{�b�[#��7�曌ꇌ�9Fb����KE�M`2g���O��6**���g.�I�jۂ�Wޥ��
m��r̢�F��EP�:�rUu�s����}��������i� ��8Ū� ����U��ͧ�R�߄{k��~���0U�I\��U�d����+6ƕpc������rŚ��p�W�j���q�]�����g��B]��e� sd�35Ô���z�u ���tVu���=�K],��ݎ}@���������U_KѤm�p֛�@럋}5����N��龩�i�p�v���/��Č����=|����6�V#ڸo�+��7ε=vک���i��?b�s7o������u��r�:[g�Y�;\֮�һ�F��Sn����#�:��އ5(�}<�i�i�̫=6��>Bs��T��[�==��B_��bw�oN ��O�����VN �>��p���k<�ݧ������b�]�z��'X�ģ-�ЦSc�����O�[:���y�����m��5]lu�}79Rv^|�7��9�y�Ή��5�<^#Ed�F/ޞ�񴡫<e�	��^˙:�r�3�Rk�ܦ�-V9������z�X��=�r���� �ڗ5���V��`l8s��2k o{7nb����'���C��T��R}�;ü�b`���JN����i��d��#[�	W�C`��m�,&�`�W+�h9E, �0��%N,ı�-�c�gw��TwW]<A����С�L�Ƀ^3���XM�3��\�XCt;A�EN��m�W��՝(�uw�Q9)���L�!���.^�)н�8D}��]NOq��o1���}^�W��ה�~�{�.O�'èU�ᣱ����^�n�m�x�>}�t�S������F�����\f��r�r�@��;��U<�@ᢦ2.m�s���?�ԳެO��i1Z����,�Fȍ�w���9z�.�w�[��-l�m.{��\v�i_���cBgTj�r�ڥ��6t�~����F���T�P4��һ'97��K�ٺÇeh1�����C"�_?��E�f�
q����\�n7��s�{��R�Z���ev>ީY�Jj18����E��6��\��Y�w�k��}��o6��W�sÆ�\f�֪�p�����]A�w������O'�Qe8)=�8�&�,\�j��<�]�o���7+2�����t6��U}
��U�LC��3.�w%����Jma�_��T�VR>���➾MV�N���d�:�31��Ɏފȱo�_,��V��镍�{�1m
ZU�|w�{��l>O<�̤�����۵��jwW7��]����TL��ͼD�e��O���e<�n���i<�	ڠ;�0��;���W�R�f�L���޾�J-��,ɥ���T�4z���]���	�U>��J�`�l���}%1�TM�B���c����nWW���gw��}3�2[�g������s�i��N�j�4�V�y��T7���"��[�s���:��]��r���w ꭩrbj�B��m�\�ڽoz����Ҙ���Ym����[1�g�"�N���Xv�R�ŉ#6�$���:���joo\5��c����_/�6�4I�Lq�;����P	�pB�?ao���zw���v>�8���b�B,^^����}��:~��9����h毂ެO�|[�O��<;k(ˮ��W�������g�B��)�_�W<���q�4�/@&�f_����:���s6�3���R��>���۹{�Z�1�*.���n���r��)�@vð�&�<��Ά�3q�Q��*�xNq�����ɒ�9{"jF�q�*.��o*qW�܊�c�)�Nٴ½���A+�-,F��F�5{]�;�C�Y�ȴ9����7
}��l�I�S��jV_Gc���`�ë��a�97'Y8�j��@'N���}Q�é`��O���{W��e�}O;x��/�5Pb��c4߭��!�}��؛|9�4�\�o0�Y]����X�'SP���yFjb�9E<��f�jܓ�S��Z���Ƕ�߳�ټ��u��㔾���]�)�{'2/dù�ū�z8���H;����=�iv��ڡ+g&�r��"쨣z�-�N���입���m�M��ᪧ�-�x����Ëk�rh�])�s5��'�=�+���S)���ͮ����ݜ�c2���`p��N��{���y��V���%M�&��[}j�6���휪A�m�*n�<lٕ�҆�.�U=5�\F�J�b��e�6�[�}pkt����£%�vn�h,�:�+�c�{;<k��Q=��7}ᬼp��Ib��PҜ�[�������]��t�U��=��RK�ToN�Rx;E�&'9�~&���f��R�v�j���DXhG�-�®5ަ�yg�{B~�my�)�7��5�ޗ�{�O6��)-�tt@]8z���ں��
"
Ya��8����vI����ߟ��t�?]��f%��q�χ �����Ý�x���o�����t�/r��P�d,��~�)T
?wϤ�!&4$��U�{�j�T^c��}�x�|���S��We�od��zy�q����p��v˗�g�+v{ӼzA	=;ݶ�k�\sit�&��,06��g�B��R�Ƈg)ŷ���D��p��g5�C�ޠڌ|v�sV�� ;A\q0���*3���^rr����
��ꚛ]�{����u�MsL;��cyƅ�[����o9]6Ȝcd��w%ne�W=���[Q�븆�N��ܪ��諜A[X&2r�)Ss��^}=s*�=��f�ռ�IΧ����xD���[}{��ㅽ]k]{<���ݧ�}r�E���U��������W��9���nRv�^�7ܟ���+'�:���޶�>,[�Gn��U�)�;*���Qt��2��W?bN�x|BB�|�4�퓢�-e�������.Y��ɴ���}���)�)�t;�.�z��h�����{�}}6��f�e*{�{�4���/�ULV)+$|m�맭�2vN�ԦmM��aY\����@�g��9���&zL��~���>�6��͡�*��G5Ss�8}��D��Lڤظ���J��4qf�j&�2�C0�S-aJs�(���.��`UN��gWt�+`�S��9O*�6?d،o�vu�'�ve@Ule��Γg8ۋ�����}�.��=۳E8/�[��QRs�'���|��}��hk�W�2u۵��R����S�Y��BOm����ƹܣQ�=�b�j!�-�6�H���}%F�n�Сb�'#b���T�izq��:�K|k�-�_�������)P��-5�{�#1�ku(_Rpaj�imd,���o��V��܈o�W�ݜ�6n,���i���U��s�\E�>�#A��ges�3�.;Q	4�7��,�sh�c�anx�[;;��j��p�n�'o�FN庼ސ/�zj�[���;��P�z�k�M�ˋ惸�;��%O��*���{-8�ؽT��v�30��'����,��,#�1�T!4w�7�+�X�J�\�G��w��1F�yub�ɿ����WQK��[rG�m��؟<'^��yx;���id":V��GO.�[�\Ť��E5F6q��Z/�Cb���Y0A��SY�ã�'Ӭd�nu���z9�L+eb�;]LG�+5��hݚ�L��.�ǩ�݂����&Q]ES�]����`-\ Ȇc�{
�1>ݝi���s�m_iL<�j��������Q�^c��E
ۉ�/A�2�/gh9����+�0��.��T9�O^I��d&�,$�0[�\U+�wm���M�N�Z��]l2��#'X��u�V�C^�=˅O�^Tm�����SÀL]ijp��k�	������+�Nt{YФ���J��&�|����:0L�3U�A��a6�R47����<�-�vR�$��|4"�F�՞�F��.k �;[`�s�0uV<�H}r��9��yc{���22r�@c�G�������m���'�����:�&�CA}�71�yȬ��ڛ�k�̆}�������<��P�Vk�
#W���ʷ��G���|�1&��m��
RKJA!����y�����]���"��>����O)P�QYP-��t�p̰���Tz�}�m%$F�
��
?<X����J���*x�8v�I���F�:)�Y����ZN6��GyK��{�k5e�����A2�Z��L
tV���f;����U��VD����u%��O��၇��Ư�)k��ȹ��G��'\ y��D{��uL9�V�L��ٳS6C�����7R��	oP��K�����ڱP؈�g%���r�J��3O8N|�9�<f�F�m^վ-�Z�r]� �N��D$ ՅM,��,�}��&�T�����k��͒!Y��"���!d�k��7�����[xl,Y����s���k�C{,�����h
�e:�X�<�.T��M��חh^?���$�J��$��ŗ:�opq��������*&Ό���'iY�e���T���hv����;x��1�<���[�_m>\2�|�� ֈ,u�(�8�R�@H)��ܘv^FBFM�|�6���R�l�+�����P��3ݬ���5u���z��#�b�s�T���$wK�rU�R�@�,���e�tY%!�ͽn]�E�Y��F�Ub���-T�LP֬7�k���D�ޘ~\��0{�]cN�\�����:J��]��l ��Hf4����*tj+z�=��ѵےS����/�sҩ�Y�*�ΰX]����豔ۼ��]�ԓ��T���T4�WL��.K�wS�OM3�5w��]�$e�mѹ�=Ɲ5�,>4Lc���F���މ��S���y�\Y}8���Z�o���];6Dռ�R��v3͕t��@�������e�o�l慝�؞���(�[��a�;�}x��.r����`� Y�E=;Y%I����srQ2�q*�qCB�(*�&�ڎ��y=�j�؄UV�$�(�\���7$�Kt��(�U5vLjv�sQ�T�i]�REE�k+�YΙ��[�cm�*�J��x�O(���xT�(�%U�Y���ѳk&�Ԧ�ѕ�Q5d��J�UFTJy��^z�S<H/#ȯ*9�-�X�g��J�F�g�m�ծ���t�
#����IUAr��)�d���ՠ�Q�<�"�+3�Y��<"Q<�"ˈWE�بznJ�*hvɒU�I�����nVb��H*����ԫ0�j�)%<Gd��D�aY�Qx��n����̔��빉Rr]H#2 ��
��6��Efzg�z�&c�M�I�R���v�EL��*m����R���\Bgli)6ݕ���U�)�hژk`q�0�QtQ���D�EY5������x����өn����[��u��kΟ���n��٨!�a���Ɔ�>��as�
����oQ�{��ﾌ���|�}�g�f�M,�&�7�7��-�M����,j@N���췭��qu�N�΍U��'\�Ô�A��uѮ�c���c*�H���-�c;J�<�gn��6�9�녮9��Ck�Q���a��Ѿy�����љPS��f*�{RV��m;�L�G��[]K�Pێ�o/z��{м0�:�_9W�ۇ��\(ua��$�G��q�?�B*�K��n9��͘������wD���E�؜ĸ�c;�ZRi�q���Q	&�!�}p�m�O׶r��v�x�|�ۍ�
�t�kTƮ^����k����nˆ��t�\��:�G�u���;�5G��=��n�7U*�*�+�:�R�Z���\5���i薰��"��tO%o�L�䂽z����{�)��5Rysƻ�H=��P�v�n�e�N�G��](K�e�O�7Q�y]k�<��U����%'WIɰ���$<��o�iu��!��A�ǝ*gT��{�E;��l�{-g�V�[�4�GkS��:�"a2��/�+>Hr'�rY�s��6�ǺIiQ��nY���Ԗ�$�R�5���y��N�):Xw
�G�����Z/�<�d�X���wF������J��,*h:}x�X��ۢ�3���]�%QKF���f�Y)��W6%0��ۍ�I�3�����w��9����æq�
Y��`���V�-ۻ��+*�'*.�q���\�|�l;��&�1�����O��9%j�Sq/�:��k��K+cyn�_}�MsLMCn5�7��#ew|�kQ�m,��e��� X��
���2���Y�o��:���7�+�r�a��{��%f�K��}��	d_�˙g��ZS~�%3���<�r��ܥ�+[��TNB��Lt�O�dR�nC��^�c��k�7΅�5=���3��
�;[�==p���5�馦wD��;eWk6�����|.�E��|�V���p����o�ǯ���[��a��w�)���Z���}�n�g1�PU���J�!�ה�����%s&����_����1*m[Z^�ژs�/���Ӊ����/G���\��o�K�WǏ�y�Eع�yWv�{�d�R��x�ɢ<8�����yy�#���X������ը��P+�t�Ej�+g:YZ�e�|��L�R��]r�OJ�;���i6���Uٷ򾟯l�LbU��S8��}���?Q�C�+��z����^�[������>����/B������Nw��Q��>�T�Y<jv�T�W\2�^8k)m*�2�ۦn]���=�ۏ�[�(t����+�6�%��:��](��՚��]����������/H׺ʌ���w�ŭJ�ૢ�9u�ϻ-s��F�}�;����3�Q��
~ﻤ������[�Qr�����5��V.�iC�J�p�8�9�[�m�ݥa�
�4jV,iB���O.���:n��\Ն�;��W�wX7mm�]�E�5t��%�9^��ɥ�]��kE���MDsL5���ӽ�;ҽì��wj��H�p��mU�u�#�El���=}���'gbo1���v�U�D{�~�*�jk���l��v��A��@�g.�hp$�ku��գ	�& d@�V�u/񭽭8;�Ƨ"��Q����Ypu>�9n��<%���'Qw�0�dauL:�_P�e���7m�����S��z��V`�!��+��dO��L[_�������\]v���Y��_o'kAW�i�&�k�4�s��Vn�P��3o�왅؊a^�;֬w�1��u���
e��u=ʟ�ޢ���;O�!���kݪ��Vu"yb���3��M�TIhe�s��i�����U{_N�$�e�����h�lqA86y�oqPg�=ih�.N�8��z��䙵I�q-��U
رJl]
������0�^�ͽ��H.��`UN��T%i��)0OD��we��>Z+�^�>���EnGm���@l�r-��'T��'iMŻR6�Y�[ϒ+)���^8k-�|�=�[�#��T��l��m�n�_cn�'�?���T�GRyѮ�p���/��_
=��i�V��v�cL��UK����;�ث]�K|k��e�<k�5�mC�r��{3WR�v|�Zհ1A�+�1Ԯ�&X��T7��t�;$��^Cj���kzӦ�✬��`�4�TI�v�H�va�5u	�����%�@իk�H��ag>̭���)�q�fլ���勀(N8�b/��j<�j���+�\��z�WE��!yd�M��}X�{��{��?���]4�V�k2ޯ�>ۏ�i_�ޭ��G�fo���|wD��&�Y׳�@w�S@糲��GUb㴓K���e+;|��)�K�P�����*��=.�YB�<{�v�����E���Y�71S���:�{�қ�ᨴ�
�~R���l� �ߟ�|*�_���=iM�&�9�����SK9���q��56/�3M�5�3e9��x;����;���y�e-��yګ��k�4�A�O*�ٶ1FDڃ��gӐ[IV�#{iv�Kk'���y�>s��j����?m��
����6a�����$Nҿr�K���VU)Ք�������P:8���u���پ$�}��w��i�f�<�ep�7�%1�TY�Yi^��g�w-o��5<t���?Y�j��wH~��U����0�^H� ��=�RO��I��[�����SVC��K�`�t�[��*΁�|�u�5,��7W�VNh���ؼ���4�Fm���X�2��c�.�/:��䷫)u㠨�y`��G`8�9���jr��^�=H���8�k���۔[lPʗn�t�J%vjv�-rν���a`Lo4���]�QӗuՌU���m���COf��:3�5�7X�2�MDJ�
�:W[nˈm��t�Y����wg**S�`Ȭ&D�˵^��$�\�����;��Z�ۍp�c���i�v9����h9�wϫ-�n�p� ab<�3�����	;؎x���0�Zs��m��8Zw��GKQ!\wϤ�!-9�෪zU��;�6�{�dcq�~�^oU������<
�*���״$w�I����`ØÉȻ��k�JN;��m%޷��
m�S�e�
X40�D���E�n2�Ml���a����G.sP���;a¨�R���k�)�]W���<�b��΄���ӂښ�}�q���S-���昚��k��o�y�x��C	WV��]�hs��Z�eY�~�s��#X��K|��ڸ�{s~����>�}&Ȝ骱�p����+����J������)� �2|nh\i9,�|8CٮP��漦��8`��t�U�h�����5���e�����U�ujH2�ة������c�8�әCF��f�Z�;�eo�X��9�$�1S��$+)�Ǔ����[�N!o�U�{��7��S;^�sڍ�Ǭ�t�q/6�r[6�Zv�dx�I��O=�s��H:��Y�ګK�m�	X3���ݗ[�:�9�jւ��.D��|��Tz�5��`uqؽ&u��6r����x6\�a\a�i�y��֮���u�ٳn�Ts��%q����9`.��j����TJ��;�
���k�%����U۰�v���dd��j�V[l,�2��A:=r�ڗ5��.��E�k-����2X9�}z����Y�<��&i�n����0S�yTK�ˊ�M���R�5�m!���v��sDvk͇��{f���C��A�mJK>�A�բ�uǝ��Ypo7/�5���<㔥*;�}��Lts��t-����=n�5c9s�7�z�4[�f�nBq���(�"�}�K�fa��𢛗^6�^O9߈I�#ҽ{Xӛ�{
�Ne@C_L#�f�m�Y(����W5��56��%�~�j��^uZr�T��JEJەU�頥lt�M���L/����k��Z����nx�ݮ�\����5/�'��u��22m(J�2�����`[Ջ�n
iXw�C��l�C�aP���A���Fv޲������`��k��ro寜�;���6�z�*z�p���\����W�d��u=t9��ӝ���]C}SQ;z+��v�-GN�kFPȵ��
�a:#��man^FW=�՚�y!�֮��˻q�]��M,p��q��
꾍vD�"��WdK̝޲�k�Ѐ�{t�K�^=~s��{yn���^�����<���*�U��C��k�ڥ%f�����{�Vtv�~���������k5�ڌ��vm� �6����i~���I�8���S�w��2��W'9���!LQϥb�r�����{8Ig�P��Q[�G��,�/��ͪM�������C |#0I��:�:C;�<���z�}~�8��a���nn>��b�<6���krm��5Υw�k��s.��k�esεެ̲�+:Ђ]b�/�U�t����nK5v�K
f�+�S2��>�)8�>��^�,��#Ư��WBh��5�r٩��|/�6͕�t��u��_v,�|�k�Ѥ3��DK���e������q^��Ww=2�Ԟj�}�~�O3@����U 6O8��r�w]�:l����{א7w'�����X��s�Y��:y�C����M�A��csV�3}�#ju�}N�-��Ԟ޸ko��j-�ۃIT
aؐF]��V�p3�r\�}I�pB�5��q�������g;kTF�ͧ��үu{&3���v��\@�����0>Ih�<�g�oTb}�����/|֬3:c���ݫ�����&5q�����u�{��>���_u3:tE������i�9���m����;e{ ���zWd�:������SEjK�L��Ӊs�ք�q�¸�(��Cd㪹�����M�ᕸ5������Y��pکY�OBl_P�M���X���<h�6j���7�Bi��²�{�Ѻ��Ub���u��Ú���'�o�w�P9cËghLw	�a�Gpk�V�������*13��4������M�+A=³5�]��h�j� 郧,�z:>׏oC�x'�p�}W��^�R�oB(s�5��#6��˝6*V,����q��%��u��� �ֺ�ܷ�.K��OeZ��g%;������J'�y-�����zE�}�3�e����D��|5܃��*�Bq���F��c2�9�f*��zo��:����J�1�O-Z�r�E�G��6�tļ�ʣ�δ�q���Ëp�;]>�hv-[/;���C��
y�k�F{�Cϋ!g_��q�Q�ײA#h̚Z��[|�ea���T*�خi������$�fB����K���ҭ�Y�4�΄�-�II�ȝ��ѥ�Vᬸm��t�	�sC�6��n�H,�:�s�����������J�joo\5��ж�q҇���+NdeI�íu��4���@t�W�£w\5A�D���)<zm�ܾ�&�C�y��+��7�m<㔥*�|�J�-��k0-�p�����@�7t�b�V_���
�n|�诞3��e��0`���$��s{M�N��k�u<��Z
Q ('e�Ӿr��e>���v�T91ÜRa�
�/'G2W_m�j�E�-o"������!�X2��yv���v_^�W�ʘeG��V^]7}���Ӳsq�[i�B�-�4m
tj�3k!�A����a��� �Kh�Җ�&��Xgk��W��u�`-\�9�TCF���y��������B��v�c�HQG��Ӛ�΢���e���M��Z����wON�noT�(�e]�`�ԇk�V�����((!�;젷�|�MXV.��X��ɬjtk �����z��U�U��x�LX��֜� �+,#:N�2ȴ��+�M�7k�T�-�`rY�S����#�p���`\y]I>���3"ɋ;�F���v�u��#���+�jXr��徇�j���(��
����ڸ��}��u(��-���E�zW]^�{ʤ��]+r`N���6��Dw ��3	p9���Υ� �y��[���Mv*�CZ
m00.��}3��#�ӣ6�bH3�v�u��4��N�A�C+x�VEfkBb���f��F�F�δ���� �P��=Ѣ���mھ�YY$vPL��p�E��ar{�do�<���ώ�w-�֞�\R�[�B�l��vK웰�1»��[���C2�����9�%���Ba�K��M���u����W
�v�a=3w�"&���IV�j8���V��C/K`����WO���H�ɓMN"3�t�w�i�]��r��E��0Ҿ�?2l_+�ݴ���u�֖d��&9��D*�q�����i7�G6���Y޵zA��m;�W�k��n.�bf�������\8j�sF<z9�����Ս�r˧@�Q�"��']m�^LP�؍b#�ʚ���k��\����^t�t|�o'z�[29Wu�ƭ�JYŀ�&-�ՠ*ۡhĵs\�h�(�3�	�Tf��N��R;����C�^S��4�˥��-�O���)>��%r�]<��-NY��4�}ۛt�b��e1�1�Zܱr` �bFYP�Gi��U���9�uֈ�쥅I��a�8��Ƕ�q�����<��%�.�y+�4-��u��Yd�K[�,�˦NC��r]A��}Ⱥ�9�:0(�*i)��wKLt�nӺ2�D)Ѯ�t�`����Sreܝfẕ�.wy��kZ���<��u���Oz�#�g:y�j�Y��V:�C�M�mq.����E�֝J����ޡ��B��
I�e�62`���]]F���6�'Mn�9<nW,� .�v�hG5����.r靖����w�VPђ�EX��s�a�4��˺o^�Rۣ��ǈ��R�8⤬�X;�-d.���O��0#R6��ݎ�GcKh�+pKxmS/)R�\䬑j��x	Ì/��2�=�Q�Vڜ����ܣb6�e��slf������D��B=%�.!3��%y�"��� ���'bؑm��P��(��؍��-3�vS@ŝ����$��e�'�Uu�䫪v\��5����md�g3\�-�7,�fI��A2��hn�8I5��BBI�䭮s��h0��yG2mI�5 ���4��X�^2t�Қl4��x��q&X�lȊ9�WC#$���`ٳ�d`�֐�U	�^QJ�f�&f��<:���"ӝ���g\�L��wZ�뜷\B�l�<9�E���.�Ml�WW"�����ɗ���(��3�m5���dR�D���4�s�[g�S1B�A���.� �3�Y3����ً�vգ$PBghº؉R��l(aQM�]��H:�Uk�Y�KjrI��d"��B0�o�޳�WZ�YҎ��qDO����6��	
��i�T��uΦ�Ԧ�z|V����[ɡ�u1k$�塛;%v>���W���v�b�ɥl޶�X�m�S�f����=�[�[�Q�r��sA��sN�ݎMDc㜹�Bo���a\LB� 짻�1<e��
�Ҥ�]|��96�j�7�֦]7�5�14ۍfH��)ݵB/b^Ow�mz����{K���z[�O�q���������o�1Y7�2S��^Q�5�jrݧ�/)��j�)��s�T�q�Ǖ-�{P�<�z��-����Z�μ�����7Q�d�/��Q6���R�á}�����8�(�z��k'�fyٞ}M
����4n������o"n�u@���櫪S�����:�¢b/�w
e62j����'��-|nk��k"��3ϧu��G���
��)���b�%�֫�e;��g=��N��ajq8��*x.
��uTmK��uBZ��-��^��
 `J��1]G}id1����/�zc�Ԇi������=�c�tݩ�U��PEYR�UÈ��݇�3eX���ށj�c�|��>CۦW���+iAz��M��Jެ�O#İ6/�DX�t#��:|��f��i����-V�������r���)�>6&�k�s�3���HF�����n��s�<�k�ܓg軙&�^��s�L����F{����)��dずN5�ٶ�H�r`uE��Ohg�Ioe�s��$�>��m<㈥��O|�`����X����r�k�7zi���z�>4[�m��q��ߜ�1��-��1Qb��{��Ԝ�9+AoV.�i_�ޥ��
��ˢ�݄�y�P�w]�jnK�y@��qԹ�B-�����=Ưޗ�w�OMI+f�F��[;��cq1��v>sk��]�{��kE������dV�{U����mL����q��+����6ۀ�J���糮*>!��ٽs,��rc'�o��̟r�s��������E�q�m���V(��|������n?��'�8gN�µ×�o>�_j�z�E�9��:r���5Q���GS
a\)ܮ����&�\�tn%�EOf����[��6��J{&ž�f���C�j�V�~wa�]��x�J����3���OE*η0n��/)>�w���xf�
�%���vD��ޓ�,��r���3.�+l|;���|�[���o��5I�^o7�F�Yyj��M؞�t�a~Q�b���v���Z^�8��OZ*ug�m;�2��WE��s�QQ�P�,�I[�����/*�!N�WÎU�v�ŵ����Q1|�26�e�f�8��\+�8��zs�3��Ő�����O�k�n��I���8�I��)2�V{}��k��sgs^>��S�^Td,�s�������]��:��u�=.':�%J����k�ކ���F��{s>��n*<�Ie��:T��V�%Un�U:����:�Έ�m��վ[f�Z����h��B�����3�ق���kJJ�V��-�s��k��i��]��U��M�J��q�������-���z���C�׊8ޚ�^F��T��Qʱf���u�s�By��m.{���l�yN"V�����X��yPƤϜ�������ցc�O۫����Q��w�<1�/&�%	�t���+#���o-����S{%n�6�w'm�rX��0>��)����`���\oy��Z�ۦ�;���*�;�@o����+��æs�Y���h?�i���7Q��g6���Qw�.7�����	s��7����q0�1�l�����ԥ��@�ۻ@dn����ʯ��im^�����ͪ�����n5�#3십�r�e��q�$�@��� _�s!RȞ̬��oumj�V�����s_<P]
�'�c}}�C�E�y�� �q՞��:�%�����{Z����z>��J5[TѸK4)�.��I�P�K*�Wf���K"m���9�,iy/��W\�q*��)��q�j�̜ϵٺ��3(���MÔ����[�=X�l-�V��{�j	�g�G��ș�&��yE[k:v��v�7��E�g"��S����_�\uaLW4ۖ�n�¾��l�lR�Ъ���*�4���zA{Q�*j"u¨��^�D[����:{ԣ[p<���!^���;�!��s=u1+�ˌK�k��ȧ�s�9�q��Ǿړ���c.λ��a�^�gP�W���F]gI�)=��;o�*��[D�ط�����%�๗�SY�쫬�Z"�]�}K��*�8��`��3���;���M���X&�f��|�}N��O��v�z}�j�{?�sy����ᬆr�ً��+E5��y�.ۃ8��������ʎ�=!�Z{�W�x��E��){��̞�Ry��/mD)J�Pߞ�A�#���]�QJq���4�>�I�v�E��t��p�r��!O}�1��a�t�l�-F4��C��d<�[k�J��oRc,kok�l�!sS�]�v@T�C�Wڜ.�q����ל9<|ob9s�M�p��&��ē7!4�Wu����^��h�q�57�5��2�ٗ�l��e�+:�x�[=ڪ/R��/>�o*��_����[<���씲��P�z��I;\uL����n6��ֻ##����t�w[K_Ni#��(�kZ����ueG$�����������B���3P�l��r{Z�l.������ \������=����v��*��/�isPR[��Z�Y����y>*o�_}�P%Թ�9cx�� B��.Y�F�׽�z��:�{îT�25l��ry�	ϋޮ6O+���w���Y�yغ'��j��(N|���t�.q����/{����3��>���k~�VOp;R���ז"�0k��n���1�*�qWT��DIhU��B�M�8�������}<2\�9Aڒ�/����/Jz$�hfs��*J�����b�i6/�m�/=:nc(<�8*f��k�Rq�b���t����KsS���v�F^k.@to�ba�q��Μ�6���l�?yQ���v�p7���c<ɢ�m,@���\�_v=�?��ˌp�^5��z'{E������f���oy��#{�.��d��ٷ6��N����[�s��Ih���>�sջJ��;6�%U�pq�vt��O�Ao��ۉ�s�m���h�M���]�:1'�v|�O�U�zǡ5q=S��i/�;�i�	���ri��R�����~V�Z:�u�l�Y��.w:�5k��I�{���#�P��輝2:��9z-_!��KD&��׃|�-�Wtfz���-�Aݶ��J��cuw2
/+~C#m:�r�d⅔�Ŏ���lsy�$�UxnF{���`Z��v�j�t�נ��I^�fG��ܡ��)��s:�ۥK�=˙l�<��P�2ب��F�;@󯆟��5=��s�n�[�J�d�%{!Z�Ϙ\=��l�rL;�;
�~R��:�ܭ�n���*�T[�d�[��h'�r����1�]�������~"�S���o�x�*���x�|��������-]��9:��k�/�s���f�]���r�FQؽvq�����yL��	�VO;e����:�r����n{���}��9ۓ'd�կF�imL�J��\���X�N��C���s��9��s�.�ͻ�]ہ-�Wo뷈��#;��J+h�?�ڿX�;)ꗛ��l�U��j��Ϳ�j���Y�7�ߚ�����T�Mc1�ONP�g�Pv޽};��z�[^����|*���&��"H�#,^_��^�ɕ5����9ҽ-ۆ��o��}p^*�cMrU�r(�k���*��k�o"��<��"��ӝj�S���F4�Z�.r��I�f��e�c�*�w�ܫ.�;'���]")>���� ��s���*j��՜�"�>�;	N#3�N�],�W�*T�q�d�v�,�8��񤳦���ud�v���K�B�%�p`v�mO;���Rw��᪋p���4{L����=����z��:������}�%x����I嵍v���RF��ԅ�
=�*��9՜6��o�~1�뉿�ex���9��q��\�7f�)��|�sݩ-��X�Y]���\4��?47�Tn�#�� w&"��D�-n���X<�Մ�MB��u;�˸o���K�G\?z�#Ǉ�_�+��{޾�9�5�'�����.<�v�,�ټ26}��U
|+�m���ޗ�{�j6�W�7��������
sNfE"�Ndij�A���%�3�6������q�R����_���ů/Y��}|���Q��7��y���۩Ch�>�(�Q&AVc'��\FZ��Y�Lu�;�d7븷���x�kV<��D�uߌ�W,�U��	G��h�f�Y���Z)�.�����P������Y�����5��ǌ������_{�����ʇ��M��~ڰ��E�l�v�^4s*�W�٩ZN�ag�b�Q�G�6�F�m{����BR�n�}�2ݭ��@3�vwqT�ա��t��F������V:��P|��ŀ�o��{����� ͜�\�ecm�p�B՛ȕ#�DMv��lQuevV�xN�E�n��=�!����Z�^"�N�h��&����Iw+Z<ǳ�Z���w���>u1��Z;���,9�/A��II�vʋ�~9욠1^d��{���wĳ��*Db�2�d��{"w	b��Q���̟�������u@<�r�{Fz͍��F�)�`+�����?�\�Ǳ�\w9�cf����N,�Y{�N�h�����g��U�3�C=��a���~�J�z��;��ٷ��FY[{�k�W��~4�-�,q'p��>T���T�ӑk*����s��F:S�ѷ�g�푸�ڴG�����G���c�MQ$��,��p|�+�H��;4?�� �l���rʟ��x����bw�s����F��|n#ڪF�:��6L�q {��JBU�P���U���9�Aү'�3��oLoF���n'޴�|}9����ʁ��L�G�y9�+��u)�n��a*b�`tm^z�d{�j��ϼ|6�TkU'�l�G�:�;��o�{�zs�FP�{�=��]]f�Q���)w�d�L=�I%q�Q֫�퀥�_��r6�5~o�V|r �q�ǯ�&��So�Ӷ��ل�,��V[=�|;�̙,�Ov�`oZ�,k�����A5���,��4�x$M�a*�Yս�Kv��KwrU�-�U�y�E��U��%��� �\!�;������n��i�E�;�)�+��� �G ����޹�ݟ���x�W�loP.����?I����5q�H;����*�X��h�!��=#�)�x��=d�;g�kb����T����(v)���M��{���θГ�1������V�yئW{G�*�7}@:~���{*�����O�T��;0�'՘E[J�h�~�S��ֲsӇ��+N�eG�9z��D>��S��ʉ���Q5�,4rP���w֣9��vԺ�W��[^�^���)ԭ'Nj�x�vڸ�:�����VF��;�&���fϕV���d\J׽�����3c�)Ф�*�7�X��#�̿_�~��V{��zB��pY�O���;�j1�"�T�qœ�fb�>(e~��%�]���'~Z��������|;Fۣ�属�/�+��֩}��ՙ�l*��+]:���f=�������o�߆���Im_x�n�x�?W��G���Y7\\�Ȣ�:k�+ƌ�B�3�>�5��w��z�r�g�ƍe��[��}ݷp��]{N}����>�}p��9��7\�6J�R�&`�G�f�����fj�[7s��(��a޳3����Xr�[I�8�+��m�ɡ׻@X{F���hʷ�h��AJ��bn��$�[�P�D�s���Xo�I��^n;�t�gwMq�����O�����B�\CrG������Hj�;/�
{Bi���s���J �%X�;1�[�^B�YPP�7�xY��^�a]�Υ�E��}{s7�.�7�|UC6[	�*gK�]���5�5�j��E|�ձ&���`�c�	d)�L@�OYy��3�@��u���nlv
�ۢ�J����/�%_ezP~��5�t���t�>䅛�yw%3x�ӖD8�)�,}}}R�u�f���ddԞ�R��]��I���mXf1n,�w�b�>˵�6o�r��z�n�k��@�]'O%��L��H�1�72`B�;*fJTv\��X���_N@�Xuy�n�Hq����Z�3�7R\����b���Pu���9�-����E-N{�kq���t��4�	9|G��Jդ�7��Zko���Aa٭>�vOv�4�A�մ��z0��@;f�`�v���Z��a�'fX�b�j��Ab�ѭ��G�S�(C�Gs��Yo7T-�yw�Lu8 宮ɭ����k�Tآ,_ ,����a�=Yk(�0�( ��JD�
O*����C2wR�r*8k�ӡ��iW�/3�=P>�)F;�L���`���]�[*e����!-Y��Y�x��=��j_	�YF�%�� w���8!����;N�Y6}���*�od.�mH�`�}��K��)p}�h�v��&8E�ݪ�d�E\y�r1g�H�qmi#	��Ju�m\U��3�;W����Ӆ1�j�o�g
͜ȍ��;�L9���3}�e3z2����Cgk���W�9�2�9��g���&�d<]�]�{�Co�LyS.Ր�fǫNI�2�<H��{m��[���*ӛ�n�Uq5n�S,��̭���oR7�3Gs����/,^�J�gcr� �lw�ݝ��{nYX�Zg��ُ���]�S�γj�$޻�Y��$M��A���d�t��q;��gT_�����0V��-͢*��K81t%�Ԫ�O��&ٮ�.���ԍ!^]�>�U���}��6`�t��z�k
�3��k�E6�GV��]�K�R�vVDփ.5�Rf�1t�c+f�3y�0ֻ��m�)��q ��c�ۨ�^�S:�h�{�X�	՚��]�]F��\}}eu]%F���(�}r�mb��U��b	�-6�Z����?�۴z��ںr�Nj8	=;K��"6�9)ӣ�ٚ�#;/R�F�ƀ����7��(\�坃��zP�����M�s]�1�����X��.��T��!��:�uwtV�Yɫ�Dd�
�:Y�՗������|�T45���Ԩ�k�1���P=P�у�r�>��q��RB���Rq����Ţ�اW�D�e�J�XyQ�S�6nvKB�d'�H���V�R�;�z�dk�vs��pۗL�-�2k*"�Gb�6���ɚa��yY�Slg;�cl����F܆[ik�Q2���l:�j���k����Q�I�E;a$TQUUh�WL͙CP#JH�9�J,�Su���J�rˑ���S[j0��3�ҳT�b:L��	�ʃtv�m��%�L��ʄ�b�V6ɬ�T-�ʫ�!"�2���n�1�"�1 �=%4��n�U�;��clS91:ÙI0�i�R��Y�E�X�I�ZT� ��Q]	2�Q$�2m�MC2$���ʫ��Td&��g�����]�S �j6�t�%�4]�	����6���UEs�Ð�UUzz=r�Ԅ�b�Z�	ΙR�Wklؠ����0�D��%F'���/�[
_8y�n�9D�S1<܃�"�[��s�����un6�Vԉgi��,UҠ��Д���W��+�����3]�;�]WzP����ި5�ߴ���<_�Hg�ڮ6��.��F�?8B�\��;�^��x~�π�t�3�3U�3�S�!7>��瞵�c��U�}q:��N���&.�p�3~l�z�ߖ��ܖz �]C}$gL���G\j���%��}�lf�L)�ޭ������=�Aڡ��#�\�P�^$=�rUu�Gݬ�<}R0Vw�T��������}c��d�<l2{�~��Ӹ�O7�S;�8]����}�*�����ǲl��]�\R>���Q_7��7μ����}�@u�9���tW�ex�����G5���/ʦ�7�Qhz#*_���r��?uǲ=�wE��tW�ޠ;�]����dҘN?=d�q�5G�d�9 �_�l��/N�������k��y��чމ���`�/^Y��O��ixC�b����ެ��r2ϴ�.�Lu|2p+��������c��w�^����ktX�]���ی��]s�����脮��E������%ݡ0��j�K�����q&�s��Pk|;W������u^Q'T�è��vwf�e�b���D��P�E{U�4��ࡘ\Mi��5�R�up�����\������\���	Bj�����2�a6�{F�.�'N
��Z��ߍ�)Ī�z�4	���.��4#ݺy�{kw����w^rʻ�����^���=�<+=�!M�A�xj��NL�|=��Й�+_��i=k���@D_sY#����z�鿼�h쇵³�$�ܲ|*	vh��/naCrm궷���؛����e@�r:fFS&㜦_l{.=��+���ep�ӍY�\�Y"��~�z�X��g���}��fULN�ңW�������#ޟx����<��7�׎�W[~��zL޴��p<}�H>�>`����J�2)]e��<�^=ޏS��w�g���[>CL�R��+�Fw�ߌu���B 5P�����Q��s��#��4���+c;�>�s2|u���j9z��%CJ���^R:vF�4֩�A�J���q*������G"{G���?T;Qw5��׊�9�����o�\8��o�G_���)������A^��tL��U珍��WzTg��o���u�1���>������{޾��猲I�fR#yO�B����Ȟu�M��D�W�_����/��|�F�j�F��|��>�s`?�ә�V�g�w�>ΏǸ��f\�z�g&�\�>���b3�
wV�Lœx���s�7h�P� g+4z@�ɺ+�����Vm�w_��K�Զ�7@Aa���(���d�M`��gU�r��'L�����,s�.�QR@�qNF�w>�J_�)Tt?(/�4�)�?i����~�����Z���7����h����_2�S^�٭�=衔d�a�;C&\	xb���\e�~5���\s���C~���+;���Q�8\�SK�[S�X�o4X��T�%l@���wL.��[�┾>IW��y��FH|��QT+��}��g�z!�RGz��,�7׀��
�d^}������++���Tr�	�LdT+�f�;|�wˉG��[7���U{����yK�ۍ��]��9},:K�]��_����D�P^�U����H�)�}�.}���įJw>g��y�%���a�L�Y�;���X�Q3���x��L��&|�'F�����l�\iw�n����׼{>v�;�Y{�^&&h�zzf�G*z�z�*Y��(��b��g�u^�u΃/"8��=�g����o���Z��t���W�lc�/Ю�ό�]s(�I�a�����U�ϭeAw�X�bT��6}�6k|I��}��!��ǲB�|�l{�}7<��(�,���8�a�Keⱹ�͑�_H�s�u��G����Z=�6Z+����v1��/�Z�����ٚ+� K%+�
�O]�H��Q��ԥ�]�٫��8cN��˴��]\;UvWUe��)�T��$�좴vnu0��ܤՔ��c�e�w�o7�;j���d`���}��e��$������\M�w�8�#�{"7��~�R6�S� yJ���Ҍ=Qѳ���M��}�������E?+�>�$G�����þ���m�i����,��3�c�Z����#�Q[��p���"~�u��L���<���R�/�ُ�l��3�Mǽ���]yl�m���f0���ޔ��M�����`��k{\��k�Ps���|�F����}�gƢ|[�ɛ}�B��˿v[J��w�j2uz�j�����/A�1�/��n�Z���1��;��Ӥ�'�y����v��B��%�,~�f� �~ːj�z����eA};�~ە�ԙ�>��b�.K4��swi�|�����}@:���}�3�b��mH/��y�c�g��Al�
g����!�6�zǗe��h�S�7�{p���v�>���u_��-�����ҹZ���u��M�;>\�Q5����!����\VR+�q<s�_��m��dC��q��{Լ^��������]��F ��f�����O�g�x��,z0��T�R���j�ny�xgΩ�<�u��a�gU�V^��=�
8��Y]o�R�ɱc"��1�����bQ��S�.�!�v�<9[;��W<9	�ԯ��3.J��,�ԠC6�[G�	� �U�V�P�u�v�s{ ;�zZ�[����38�R�fK:`��{l���,���_lV�T�l]X�M�-��npV���o�ŕ:nd���a�|'ȱqY5��]呦��������;�R�����|��]��[]�ީV���E���<�#+�X�^UP�'Fs���_J�N�j���������}��#~�눿W��G���F����qr�<jJ�2�{.f�����^�ڧ�۬�����P<n5��y}^ӑ����7��[�ɺ��l�JX$�����N�����U��;�ú�r�Ż��q^�X��n��#�#���ίj�}�q��מ�t�D�nM�a8����L_�}�@\��
S3q�[,dk���z�����{�h���=]�}�!H凒�n'��^1��>5
	TQ[�#�^s��炸��C�D����=LJ�a����J�˂�p~����{������2Y�@n��11+��o�Z>�j9���ۏ��������:�!�Gw+c �ԉ�|=8/ޜ��ng�*��=$��&k\���͔��Z�c�ǯ�r��7�j6�~�oޤ����}�`eɜ�,�e������T��{Xo����~�N�b.͏]�V��C�v�_�N^Δ���=_�Q���/]���az>|ṽ2v�#���W���i�#{+q]78e�˛30��.��Dq��D4��ľ��޾k��ӲBW\�V_I8������g��1�kqU~C�j�*���r9K�|��Ͻ�wF��F߽@w�<�}�&j�|��c7�4>ix�����>	7�X�m�s��Zpn������u��o�h��D���l�<㷛;7���!�#u<�-�->Ұ��(�P2a����"��tJs��Gu1���ᐽ^Y���Q��w0#|���->���~�V
���P���d��A�^��a�e{�Ժ�w5[ >��Ǣ�sNdK&En�����u]}�;�/�uc��d��T���,���U�.��u�ia]e�VM~p$�x�o�9��{��� *#~��_�'+��s���k�gNIۋ�O���/	�.;�k��id�*���B�}Ѷ���9P9�>�O���/K��z�=������m�QӒt<�8��׳�Uʋ�K�N��)�7���9C*g����J�P/��8���x�9���dz�Ǖ���=�ٯ.L�f���#��f��$��(	�h�}t��r>��Y�n�M�?_��G���g�^3}%�=����/w�n,��Q��7���F��%���K�"�[s�����{8H��!z+ٻ5cӰ�3�,Ėl���>�W�r�죙�Q�&��F�Y�s:K��k��u<��J)�т}+�֟��f3Y�xY�s=C�9k}�Q�{��ZU���r�Z��u�We�]3+���[�S��V���w��cΨ�c�rh�9�����m/ޑ����Bt�ΝC�%��ʠ�10[�&����bI�L�_�{�.�wm��n>K�ğyZ
���o��p�}���z����2\� �x���o�l��Mqʪ�=�=�W^�}�W�ݏ�F��Q�߭��Ӽ}㾝����|�zs�Y$�p����!_�([��8����
�WM�/���#Q���Q�~�"|r�<O�:�)�C �E�	�T�og�{�fG���L?`U���Oxк�K��*|n9��z��wF.���&_gT�Y�,�Af�+-nRj���MFWJ�$����L>��1Q-m��s�4����wzu��h�qdzv�Ws��w��=ʇ�n=���>�Y�@gޖT�?�� ���.�;�^�w�<��)s$Y�f��}�����ᐝW�ȇޡ�K}V�~ڱk2�f�BuV��m�{�(�}���W��_��Ǻ����ӑ�}�}���!�W�����P��#��'v�F��$��KN�����s�l�ͦ�݇ǥ�u�Zn�|�G#f}�y�x���P�|�{Σ�|�x����?o���b2;�YCK۰qQ{���+O
h%���G�u����7|F�7#���V���VѮѕ�u��*k9ʎ���#:�����dď
�S_p��t��Z��S3y�)�M|*VVX�b�}Yo�N���p\�\��b/Fμ6�Va��\�7���?�fm�N'E�L�wR�迪])͙`-�B�?����h��Y3=j�M
���G.��ߕg�TgeN��>'�/ ��TϨ�Es�����i�x���8 0H��n�oh�|;к���J�f��B�F����0�AR�Du�*�ҹ��Pu�^o�EuwL��]��+�"����FF�'��}�_��l{���E�E�UD�O�CޮgΎg���r,��m��+�r����^�\Mķ~Ӌ�<�}@>7�hd�7��@�y� �W��+��\����B�ݏ:���U�n<g�y��r3����#�Ӟ+��H���\���4��P�tԟ
�ML�gx.h>�#I��t�8yjP��I��:�;K@Ϩ\_��?ߩ(���.�������2gS8���M����E��|��2vs�5��F�ܕ��ˎ���^����H��X��>���y�u�:�E��&az���}^�VK]7�X��`Z�<5F^f�s�פ`�Fw]ȸM׉�|=>}��`�� ҖOP2>ʊ�պ}C����n�L�;o�]E���$�q#�xj]�������є������WbG���p4��p^��@+kys;n�:j��%z���P�Ֆ#�6�[����{��P�ML(��6�>��Jt�m�C��ڭ��I��Y���N�N&��·:�j�8Ҥ�v��M��@g����������C��>�g*���ڐj���ɱ�>ʊR�܊���,�p�R�i��|R;	O���T>���/� z�}�1;����&rbCN]ݐk�L�<�η�>�����)U>�t�Gt���W�S^����x������a8H���RVX����3�0�g�Ggng��@���(踩U����L�;�2�~?!��˨�'jE��������ۮ���gJ��aہ>E��ɭ7�K�<�4���>Z�7>���;�z�������ҿ>�x�wHog������?��YU{_���w/p�]��SE�z�Zkz��v��z�C�/�E����~�,��&�}��m��$񯤯���B�DW���#6��]5�7�zP>7���ϸ���#}#��Do�=�9��ׇ���U�螛�C�g���iw(^�I�X�.���n|7�wG��ޫq�߸�GzG����ǵ\>v3��[��eO�0�k�~Zk�`��e�0���-�3]�x���Rs�Z2<��ѕ$����+�u~�m��1J��x��skE̫���/���j�.T�xك2�S�$E��ZLNj�̛\��ܲ���3�У�Ewr��cLʹ�r�U�jn�ЕR��\:�aݹi�좄g��m\���E>�tF���u����	���{����ZS`}Eṁ�9٪�g�f���ULÊ%�������I�+�w~x-~�4"&te_�z�jf�-��X�Y����Wq7���ꯧ�G&�H�Ot�/�9+%v����R:/0(Κ7����%�#�ǽ�la�������V�z�q4�}2��ٸ=$"���ϑţ<'}��P�*>��^=y�z���y���m_������ 7��N�ɚR��}�����^��q��lz��5��#��O�Z+*}�{��7��q�y�QOex�/ސ7� <�֗�~d������n�C�2}��"�����wR�迶�_�wKң����o�h�|��^���Ν>Td���b��䫯�%�6����p�q�*�L5ckC��i�t�q=�wS���I��՞�G��c	�T��s���{yP^�ޚ��
����-rWu	��Awhs��K鲮���$x�w�"v�j� �up�:�_3;Լ^}�V;�}�<+=�#d�l����Cׇ
kp�r�`m=���$�%{M /?\�Ey����}9��͹�>�殢�%� `}>S�����(�Xe0NtZ�9��-_E�%ӹun��iaa^W��ӊ�Pk���č	mn�\k�;D*B��[�����(����$]��W�#nQ�:b�<ɼ</u��[�h^�qg�@��n�M�ƩyK<�-��m�A��T}n�Y$r��fZ�J�%�S�Rk89P<��[��OoCʬT�.��_d*�1܄�v�&����[+��5��hapt{)�E��}.R�˕{�q�(C�}w�u��Z�m]F���ΉV�\����f��+��� _*Y�n��m�n��BǍ��ަ�.��f��{F�f��E�����=f�OFX��G�)DNӌ3]n�%4��y@-��ˑŽ7ee��]�%\�;�X�WI���bZ�n3$nU��,���
��'ac���=���������iJ����S�|.�=qfQ])RM�)�����sD��Z�D/��ҭN�s��r�nr�z���U=[.#b������"8B;m��b�@�뮼��r�VDz"�@��U,�y������c����#EMc�2�6;q��n��{U��#��������_ ��p�.�M<�QY�%�鄽��dgjN�2&���D�f���n�AH���C�Y��f�i�[�~�ۋQ^EB�p�b�d<�}�5{x��p���0��ΎVpܭ6���-�)�)ލGLu�ʮ���@�9V�XKBsB]oAu����Ӥ�7�>�f�6��9��U�W��&�]�Q� z�qݸ�p\�T^E7/�W�f8�U��l�����<��0����F�\�b.�AeCq�S8]�Ϻ�����J�YmnJ�)���W++m�;p��ͣd�50@�)���p�v�9��n�=�����y��3:�8��wq��Q�M��re0R �Rw�]�<��� B���&vT.ʝ�v���P�]-^�jB%�t�i7v`���b��u��N�;J�V�ە�����qf���%b��w���_q�s���rZ�/+������.����v�v.�(�xJG2���:���F@/�f�.Iq��Ft�J�Jܙ+Vs�q��cA��%_[q�V�Iaq�/9�l�;H��r�qM��k^�)Ӂv
�P��A���Q�>������8 UR3%k_e�\�/�֝}������s7]`� �5�{�<�_S���n�%uA�6K6��9Wq�5���Բ�.���X�t���W�;�L:��[ը�3]gj9��r�f�4������W\OX�;��>���_i�$mj�{i�5�y}�"A��� b�'���Ʈ0ji��c'$Ĳ«�+���Jw*�d
}��F�޳{��P�ɽq���{.d⵽���������%���{*Q����h�cӜS=e��{0�Ǌ\�Ƿ��,�RҺPݷ]:n��N���Wz:�i՛e`���B�}o�~:��=�fc�V�:u�0����V)��s�71��.�o}�~H!I%�TB�Լ�ɞm�;��(�L�$L��	�;��iu��H���B��ڍ�i�(��iI�Iͤ���g���W�a��53::�!�]4%4Y�Vmh]���#n�DA�]9\ٗ�������he����cl���ʩ[D��r*:�u<j�F�=�B��65�m��ժ	)�����%yyI�S�3�"`�m��ʈ�����Hu�2J��Z!�$J)YbM�ۑ�����k��{Y'���d\���Ps�6,�v4�=�t�I/I)rd�f��T!Dfqv�b��U(���uҠ�g.Bs�!2i�]g+B����"+Q<S�k��i�m��(��CtD�9����kN�5���v�&�^�^��CB���UqOEvLg��!cP�b�n��%q*�b((�P( ��W5�6R������B�,��V���G8>�x�T��!:u>�\�ِg]%���㝖1�{�������<�R�}���V�]��,�|f�6�[��uҠy��q���W�����=/�7^WH��]I�3q��z�S\����I�+K���%�=�����t�����<�����g�x�9��>�\�G�ŏxe&jg��R��F��ͳQǰ�7�����b��]x�Z�,�7V&������A�]�Y�*M͌[�{=���w�v�w��;�v|f�a��䢇�+L�$�2.:e�9���>ԧ|*f<���{�]i�����ѐ�י[�z��~�BtۧP�\�j>D@�3In��^�OL��]�Nt��w��>L���Tj;�*�Q>��2���k�p�o�ꑷ�bk�2\�" nNb���L�D�gG)�G����|�}���GZ3���#�8���v���|�s�_%�}w�q�3*'o<�^D�D����H-��B�h��
_�ۄ����?O�>9Ӟ'�Df��`�(�7ޙٯ6��lҙ��ǧ~30��X*\����K��ܩ���������qÜ�ў�<1G^W���e3G�vϠs�f�8�̓��'�L>�>��ތ�u�5�wS�R8S�j�	��m���QC&Kı��qݱ�/q:�'��`��4�:��N�
r��Z�3�w�"�r�����*��<,��.�^�j	Eau�x�&Eȭ.oGv�e���]���l,(�k�$ށ��P�zCB��5F�QY�gb�^CG��p��M��>z��4X��T�]>%F}0��V靯A]�;y�}���y�������oo�!z�Ⱦ����x�?mX�Y�#/e���8���5M�e���E_�u�>��my��ԭ'N}��7���!�W����B���ܽ��9��uXdOTV̋��^A'���rϊ�
rgN��(�L�����꟏��gz=�p��u��q�TT�E����貲e��Û,d�g�>���])͙`+�.���O���.Q�^����BMרor��/�+��v��C�MڱK�ڄ��Jx������/8��:�`����}s>�
��y�_�#۱����q�<� ��]�(ݖI�0�AR�Du�*��a���{�>;���o]�=����~�
7�>gr=�C��x�k]<;@�Z�5rKd&8lkh����⼅��v�������Y����u�u�ܷ~Ӑ�#�{>�� �ߵT���S��S�a�_�X�Vϣ�Z���������>�y��#�O��n}�H����?H���\��/eGAUWa����Ȳ��s}��=��ODV�b�wMMl!I�ʴad����LI���$�h�"�<��>(N�cMd��ԱK�oW:B�$���[B�u]ͨr
;�OM��n��A �m���Atՙ8�t�K�; ����]�$K��2���S����}?�
���㠆}R���9e����s�޵Hv}/�ٌ�Nu�u+)��]Y�ǐ�Ṱ�ͪ�y�Z_f�yCf~L���t����A�hd+t�{`9�����Wbw����1B��Zͯ57ޡc�y���>�d���x=!ξKC~����H}������o|F���u��H���٧�nԆ=��E������f� �����K'�����B�3;�fH�=�íU->ە�՝����_�G����=� ����d3�b��R)�*��S�Z���v��)pmx��0��S��m���v����������ޠ=Js��eD�����{��9��dm��7�;|�ܦ_�xh��+�l�wY^j��<s�_��ڸ�C��q��Ox��R�y��a�̠]o ��_��f����G��ۙ��CgC��tlT��N�`Tny�x\{����"a�3]y�W�h��p>����C�X���1~��)N�0�"�'�ڗ@y6��K豽�pf��{� =�i�����{ǝJ��y<*3��MO����qn����s4��b����X����xg=�������4z*�-v.�ʶ�i õ�#���\�Km����R�`�'���Ӹ:�4D����s����ƶ��p�%�3��������v� �/�;*�*�U�+��+P��!�c��f';K��ъe�����<��Y���Om��<��]��&���s�g�����^%��J�}+ݿ�;0�Niɸ����wp��s}#��F���S�z�xvD�pQtA~�񾸏��L�jA_����(}Q>`5Q뎺���b���ޫ�״���|C:��Ҭ{^s#$wa��,�gz�\`�� �,��x��l����r��Bn'޴4[�o�Up�h>�ڮ2��J9W��G):U������a���B�T}D�I2��v�ݖ��X��&�<�5��/`c�;�����c�������Aڨ�~��\�Q=�^${��C;�B����w��ǜ{xLo{Z�-?;c �ԉ�|=87ޭ����Y>�[�2=����8ɬ��]���8^���o��n+��z�T?�f�[U�/�x��XC�re�+���*�dL�Z�Kę����`��]Jgh��/����q�������M��P�B������a)����W{�Ҳd�tǊ����tx�{R�轷��Y�O���n7�aI�^�z�6���$�_�~�I8�u�W^ս��Nb�bP������P�u�ZG�G&R�y��/�Z������}׶�\�
˴z��T�)�nb�+Y]�/t��RI}�:�$]�%�xl��`���j�6oJ�8s�R��ft�3x�,k���=��[Ӣ�_����랶�l�a�7�q�*0�Z6�9>Ӄi:�{#����ʏ��ם{�UK�0y�%������z����B����N`0��N�9>�R�۪��ԔL�w�����
�ܭ +q��ȇU��g~~���<��q�<:3�R1Nf�����������^�9CyV�p�J����h��k�M��(�r��9�W�5����ݓ�gNI��s����@Ͻ͠����}2���C�UTv�}��tσ�>��_���.=�+���F�������f�x��1��|$�$�K�����J���S�0|�{�a�W��������]{険�M����~�[�K ��{�v��X<��J��-ee��;f���ӄ��r΢'i�O�����c=���\?;�v�qD������bK�"�[s��~;S�0@[~on�{��~�ފ��$\��џy�y��'{'��n�C�+���A�e1Ǆ�=_[�����&�X��>Sw�'�g|VǦ1��+���yb�^G��F�����m�ުbj�r�n9�ߧ�1<��瘶$�d�ahK�h��;ى�����tyg
�tF� �o4/�_q� V�PL��w-f�*�w�K{o�
�XfW�fS墈3���s3\���\4���H�+�s�Z�>����혧�ow{��q��nn.P� ˑ��O*�x��|G#F�j6�o�����>�߽;Zǽ��=<x��1�;=�7h��u���g�\�/M���g���}�B��G�l@R�n7��m���_��>,���}�B�W}�kʼ������L�CǧL�/XU���xп�.7������nS���zs�����/;4}����3Q�}fIϑd�a��'�b�Z�ћn�Ɨ��뚟}�0}��,��:���]п���K��ļ���M��zYS�Kd1�EޘO���?Q�Α���s��yq�=��W�ö��:���>�Y��x��ՋY�#/e�����eP��Yd�������,>������7����5K��~�s����9�u����@�g^���v5��m��js�K�l�;s>�EΏ\VUi�%x�n2e���Q������=s��(�4�O������z1��}�d΋��Z������_5f�����[|N�Z��*G�� ��ˁ��ipv���{=j�b1Y�S��|��,e|�b㮫�g��\h�epة��nP��9X;/$k����g����B�a�ܬ7����)��ܻ#�!��@K؝���}�1�
eb�2Vqy����j�k�m
��8��wVu����V�Ь�D��5�:�R��4�Hs\��h�Fj�
@�`M��T(=	��P�V�L�K;{�+�/�{z�܏z���]!�o�R�F�$���~5�LO�`����\ �5���ԩd�]>�ʃ��Ї�#�^��3���P���qϦ炸%E�Pw�"ܟ���a*qp=�����y������u��Kw�+�yν� ��{UH���0���xzh{r���Dԫz��q/�d�9MD�#μ���uc���Q+�z�#��V��#Os��M��>���u콐rmJ�H�t׌��2��[�"b[��~,b�瑿��C�_��N[�@N�����O��5����3�M���Uxȧ2Z�50��� ��43�n��hs���5�0c)�l]8S���N�H~��ȃ�+>9ӌ��Td
�N�j�z�L�������E�x�t��xg�s��^kr�{7������ʪGB�����*,��.A�,��C��sۛ�>��lz�}�o���G��{NFܴz�����~󚢾{�տ_���g*���ڐN�D��Q2�lY٭V�M@�|vp;�[��ۗ���%/����<�O�h��P�9쨞�bO�/v�� yP��0�Yȅ�s��̮C�Z1EE�g�s�5�B�.#u5*l���;n����-�����ʵ�B~j$��>ޗ�8dd��ϖ^�l���7H�&��'7���E^�s�z��ONH�� ��J���K_I�6��������Q4�n>S�O��r�G�
#�߆·u��J��#�_���=+����Md�\��P��!?�z���n�a~�w�?Vic�͝G�go��6t99'F�J���j�OȎ�K�N��G��k7���`�Ω,�;�eg�V;����ӿ"���	�,_ՓZg���'������|g	�=���;~��W��<�P�<�xg\Κ�r3�{ӨG��WfnRH�����W�^��wF����i����K���/����|?�Q�u�m+���ߩI�-b��>P�d�$k>�3�u�JM�],o[������9����7�����þ޼8Hgʣٙք�f$sB� �*�P$�L�!����T��l[�>7^�X��n��;�<_��j;�B�$j�=���|,�Fk�]�s��6
5
Ue����-�3��{��ߗ?L(rs��?+1�ݛ�s	o�������W�|������L�(�W�	I[�"�ey��Q�G�"�@��T��y��a�m!��� �i�?WbU_����;��)�Ot�^$< v�����]��l>�LDd��p��'�Z��N9y�Sz���-
�s�{s�7W�g=X����cF�az��v�2�ՑӨZ�|.�Ӿ&W
��6�*����Qt�������I�2��/�N�8,���:�Y�ӆV>�֧٨C:��y���ܙӦE���i���]{����^/�&5�k$pOΘgޤO�zp2_�8z�q5���t�/pI����#-yC^�8G=>�*2�[����f�nW�/ޔ��x��� �����+�EW�FϦ2��x�o�L�.p�g�l��Q/�E^]/�������|�W����hڷ�i5��;C/�k�k�,��]�����5
a�4rX���V�O�u>7�;ۇ����\��eO*�yz��s�\c7�]{e������Y�;|J�0������t\Ru���h�b8�/Xӱ��z�G�?}��p�N��zGzS��X=q���|��8o�,n��sL8p�ѵ�$efW���2rP9�V��׃��j3�~���������Y;�Z�cت.A�#f�Poyסa��93�b*gȕ�i�*17쑎���g��z<�pX��8����{��8~T�������@p��X�\�u���P�,*���|�3��=�G��^lP��G�������^�~Y?W���>�D�ip�D�����5S羠\޿U��}^�Q�+�M]��1�V{��p����+&�Cv�[q�9��ʓ:`oO��:��z8����-��u5�(f�8�n��>w!6�z	`��ن�)`��U������9�,�b�[��MƝ��vS����>�6�A�j7���L��C��.�<X��2�mFMW �9oha��ҼV}�wXf��#�e�rA�2��ȱ}t��i\�m?r�^��8�f]={i*^�>��C�G8�1������3~0��rQ�GĕPe�/L���i��ӗG/ou��i�ީ����勵^��=�2�<��W����7�C�%�(���Th��
o��ŏA�<y���3��~W}�h#�#�ӣIQ��HۏU17�������'zhʼH{��O�4���"�θ�2�����r7��o��p};��>98]敘����ೆ�������t�3]2KDI�Ξ��(R�h�����5p��QI��L�z=+\�s �ix���N�|vsĸs`l9�3"�g��`��=�B���yʟ���ĭ�%E�{�qNF{�޻����>���f�8�̓��'�d��>���e�l��fnx���+C�9�p�=w��o�t-�:������,_{*A�_��B�{]{vo|�{j*�sߵ�^A�i3��1^��i�_�+��q�{~��W��}�4��`��~ڱk2�f��Q���-�0�������9�ŪvZ�+�[��1��}�f�b�N-�Y�iG�L�����P�"��vz�krg
ԝ�
�J��'�x.ؤ���^I+rT�iS�qm�!d��O�N[ٜ{������Ψ�˥�&*�M��-5�o8;�Uգ-�{�iR����j�<��z~�+U!�/�A;�Jl�mM���k{�vL�b�ł�lts��͊ؽJu�fuu'+i�M�!��f���g��wS�lz�*Y�\Y��P|`��&٭�a)��+2� Zx���`�s �*r£�z�ա���ho�\U��b�]t;�`��t*r�խ���z.:7���7[V8�W��;�Ջ�a��z�i)���'�E�V*��A@i�][0�u�V��^ �t�G����\���mfv�F���&Cm
�+�$���%�!U�A��ӝ��ᔸ�rp�)U�f�����Q������ :���]T���7%��m���v��mK�nN]q��V9aU����*�Z8�v�֔�&S�؀ޏO
K�`������N���Qm�/��n�K-=���>��׀��s���"̸�@��7Z2��.#��+�D�fi���i�Q��ș���nTu0�v��c㪬C-�ٝ`����]���!�Za��9J̔�J��ӏ:Ҹ�T�)^S͔�+��?����o@��$"PjF���3��Ц3[�X9wj��w��z��fث���uv�sSZi�pPY��Z��!1�.�2�:4��.��̨�f���G�ö�\���$���G�ӥ;/�<�^�\.���򿆡�۲֛���n�Ԉ��5�.���mmWل�@7AN,�<�ۻg�ZV����s���&sb�c�e���t�p��iW �1�ʅ���A�v�k�����ctz�F���X�5��������%���n*����)Z7Q����Zi�Sr�/�t�C]X��n�zΦE����bM��Y����U�H2L�i��Щ�TS�G+��n�"Ѿ���[g��J��A����I�Wt�\Ӈ��֢���3�좳F�'KqV�ؖ��.�!]u��m=|��W�������ywܶJ��d �,E�W9��K��M��wA��an㵴�.O(i��e���]���$�d������Χs1cQ�[]��hn����{S6e��8K<ˏ�I}8	�+m��A�6f1)���ܸ�k|'^�z��Lڮ�m����Qu�����wgB�U��5[��{'�M���gv�n��q%��f^�V�y�䵾�9�[+1e���t�u�'5x>v�q]W�d����Y���v�Z�:�S��>mf�ތ�����,��k7:�SxgDm�iR3�Yʹx�R43�O��WpC2�O�c��dL[�}Ʈ��O���G ˤ����Ke��	Oi=.ҵ"��Ȃd�\���NfT`po7;���G�\�T����P�
d��s;�jbрe�G7r��WA�h�H�Q4*�B�^���nWc%h��I�E9�W�\��E���ذ4��,�D@��1QL��͙��B�4���4�ʥ#Et!ڃY!궖��(�v����a��X�2q,UWd�̋U�h��+`����笙&T{Tɐ�L(�3Č52E3֦KF��ɷjW:��0�&��I�%��6©��c��.�唙l��!Uh#)�j��v�b$cc5h��l10�̂C��9��Vm=/T�R¹���,B¼�4����^Z���͙rR�&4�fa��.U5�sd٨��V��l���56���=$-�����"�t�U�\�ۘ�'��a"�lJ���jv�;ebF���K=�mNmP��J�9�w�n��j��5�%�dRդR��^F�Ξ�c0���LG3I5��h��T���#��l���U�w}�b�%��D����)X���X�v����آ��ú<��mM�� i.ގ�ġ���fkxɌ��i!2����/��q.��d]�����3�S�'N��w+��Ϊ��g_����wQ:��:�s�~�M�ػ�|�i�7������s���YU�I^%ٗ�y�{"S��&� �'Ү��������p�*�5��΋^��ne��x,���t_�.���,��L�u#��������~���w��x�W�p��Qn0Id�Y�2��,\u�z���&�(�W<�Ϻ��[מw��Xz�~�Jܶ{��C�>3|aụ�Y'���^�O'���y[�x.��fא�]W��>�eA��7�!�>����O������z}7<�����s��iaW(�6��\�z�/�f=KU}u��������Ku�+�yN��� �ߵT����K~5;/��-��Ū���T
'}� ~����ׁ��-��k��G���&�޴�Nx�2��Ξ���X��u)Y�z����5܍�4̲Ag!A��"��o��6�V�Hteo��WtM_�����K/�Vc�g_�w�;�߽����^2%��50��� ��42�^=�XҌ��xIZwp������ǀ�j.h��|��˔]vu�����F.����iW�]
iЛt宱*��f(����K4��ݤ떚���GV����(̧�EE��^܃��y�e9�|qů��a�*a���^���:�"$w�7�[J�'&��h�Az#��G[j��>��<m����uP���L/`��B��]�i��^�R�>T}���y�z������~Wr.�x�g�=>}�3q�TC�\�JY=�*V�r;DÏV!�{����eA��p��s��ꇥG?u�{�j��H
��~����=��z1�eoga�Y��ސh�=��4�[�:�;E��	K�v��<��v�>��R�}ԧ6`y��q9^�W^�%����f�>��¿�:�W��*|O��~7��<�ٔTׯ���I/c�����Hǣ�R�}�;�og�3�����������:."�W�wׯi��xKfGeEz&_>j�@{;VBe���]s+=�ݟuo��T�Y;�fP�"�ݞ;G��&�.A����_�%�ʌ� b��iX�o�FC���9�z�����'�FvT�,�-e�:Ͻ��u��>3u��Q߫��}v!�zȸ�K����^Y�C�d�pDeoј+�[5�j�_���32�%��k>S	쎩�?4�q\�ۻ��}^ӟo�x���Ǽ���^����V�Ǖ�=ŉ�L��s^��k���KRk�e)��ֽ�֫�X�#�xwt��\����U��3�"�(�r�8�&������Yh�6��%��0����g�E�7VQ�yb�\��,I8��ȋ���e�7R�����ƌ�Ž��`�ԣ��'�/N�K�O�ʡ��uMφŻ��q^�X����v�����^]��{�x#�����}�gp(s�*2��
W��l�����*ZK)��
���{��'�9��Cy�|_zF�q�������w�P���Q���H����^g�`{�ly��]����MN��}�CB�y���ƨ���&����~�TMC2Y�D��\���s�ɹ�)����}dǧz�F��>��l3Q�Z��sĿNM�{ޭ���q�^N�6=s=�f�׷���37�d=7�DϺ��R���P�_��j6�m_�����@����W��ڻ��\��lʚ�j���mR�5>'�'�!���F]/�������}󻣛}6�!X*<�P�K�&��}@s�s&��mLk��^|p|��[��u�_
ϻ��ŝ��>v�t΋���}تW8�>Wh�C�Ez��e��~��|}�p��+�0Ս��}�E`^���VH�>�v�۩^W=%z9S�n�xd/W�F>��{�z����f�F�N홅�,�F��}��߮��8�N꫙���'��Cet����+��6��+�g/=����w�"$�Qd��h֖źO2Nc�,�3�Lq��-�,�V��I�^�"ͥ�b��<�f���έmχeN)���.V�E�P�g-,��7���IWz��z+k��J�s�V���~�|̿Ox�)��vΏ}�ʑ���9��4�e�7��	{I�2Ϣ
�C�ʭ72�J�,��&��2������}>ntw���jML:zzg�1x������OR�iu/By#j2����p?rэ�=��W�ջ��`Ё}$�S��{���ﶾ��ᾭ>�MY�\�Y0ޟ�o����T��\�k�Xojqێ��܉GA��[W��ݡ��r��+"=n���ٔT[�Q���X��u㋣2{k
zR���޻���ڱ6��ޏS����_���ݐf�a��B>$�2���t��/�hG���o��>�鑤���S�w�AI�G�י^Rp�t�\���i�^��ͭ:����~�0Ğu�������Q�~W}�h(>��=�?W&����o��`=�\�k�s8�z�9��>� �K�&%��o��}�G#q������G�q��+�	�y��;|r��Zr��ޭ�
s�i̒ѳRٳ�D�/ԅZ�h��
_�����;:�;�.�4�����b�R�'�����r�̥]M�6�s��sI���ouD��me�o��I��$4�n��z��t�SD\����Ka���:HھX!W��>�Y'�Fuv�1����>�ַ5۰�(+�ݤEd�o���k��k��)%kރ2�9�6���-ͤ�o�T}�̟�~'�����|�>���lo�g�a�ϔ��t�rh@��U0�Et�%��4���ouH�����ů?Y�q�O�w��ʎ�Y�i�L1�ԅ9��~����Ą��gvV����}���k;�î#�ކ2!�]и{��ߧ�Oy�
�O��Ў�g�i#�U��z*�u�[�Q|}����v�߆D/Uy}�4�7׀�~ɠ���Σ��ef���ڔ�zC����pwj���Խ'N��_��j�2U{�οT/9���4��u��Q��Gkw���D�,��S�r�X:v�/���wYU��W�G#f\^u���4'�αM{C��KG�O��|{>^w	d*�6?D�w�l�%�l%��_��>k�~�ӼԌ�)z�i�<��a��m�~>>�׼{!ڸ��X�g\Κ�r2�W������$H�Q��gs��j���P��8���z|�G�n[=�t���4���!�'V��F��y��u�?eo?F���a�˧=k*�)��z�(��O���P���c�rnx.�R�=g�]ur�_;���c�p��h�ӫ���V�Sr�w]vt�]4Z��c�bO�)�Л�[��,�z����:��$՚IB�����=��>��j�q9B�I��^^ϭv��,v;Xw#�S@���'��+۾0���cZ�bĥ��8���v�����<}�tp,�P���������{�q7��NB�9���1���lMM��-g�'�L��/�,��Uxu�d�� ���$7^��-��hj*)�\M��֑+�G,1@u�ck��.��}�R4��T��4̲Ae@�>�&%��x�� 瑶<|vEz'��n3���w������L�q��<��g�̎mv��,wQ�E���rj}���B���U�*.��w�σ�*���x!�>��<m���F@�N�j�z�0�E�����c�꽘��؜�gG)x��tf�[7�TǮ#��G���μO���g���`�rt�w=���y�%I�g���7�yP}ӸwnS=Y�p�����~�:�7}@:~��������J����T�S���2������6׫t���W�K��YP�"��#�rW�2;
�%5+�݊�>�~��m�N���z�oc���PrXWgC�����oo�H=�?�O�dӶQ>^ݙ�C����{�o����f�?36P�����F���?ײ;'�����������\�`�e�w���E����1��q.!���9Ϯ��7��:=Z��������sPx_r�I��`�/:�L���s]F��g�Gy@�܍AJ�S�)t��$M��k��=�r��׺��ܻ�|2eNus�p]����}įr��w
S�x���2�须�ռb��S��N홇��������<���^�*�Z,z��7=@5���F'o�FC���9���:�3O<��S�������&k5:�<��N_���_�C�UTv��y��b�z�Q�~��߫��+և�u~���z_�<j��U��^�Hwr�<k�-�T�Ȯ�����7��������������Č�U��ۃ�4���!���pW �*��I��%�?l��ʙ��+�S��E���_��B�S��}}�G����Hg����8˰liAʠ�`)^3q�[,m��H��vi��\���F{e	-�c���ޑ�\{}q;q�a��D( $=$i�ύuvV�ب��p֋��#�3�S��(��C�O��>ζ;a��������PO��k��eg�5X;�x��L�3��n���&&yWQ�)j���z����'�la�����{Ӏs �Xr�ϒ�쩾����9K���ύ��&_W��-�U���f�[U�)���?TL�Z�*[�~FEu��$�7y}٘��v�@]6�.�����묑	+�V��bc{+Vv�®Y����po[���NX'8Y�q
j�Kw,��1)�u	�q]ɫ@CA=�l5�B��*�<KFݞ왺�.�������5�:j��p�q����e���ld���I�S�x_�|Tਗբ�2�x��/��?uǏ�6��99�Gӝ�g��\uz���S�M��@w�<��dɥ0ʚ���G��%a�Ѷ��*�����/�I>���;Z=(�5^�{>��]���^�~�by���Y�*#��T2a����&�*�Y ��m���Y׭_�(M�w����۽����;ҟz����B�{*p�d�%=ή�,υ6ED��Kw�Y��1Ӓ��T����~ V��9�V�)����:��r;'�ԅ�55|zw�j���H~���pf=��U����qS/Ĭ�LQ��d�w/ޓ>�ǳ\=�������|?UW6���`��
�:rN��%������B��]ѿ����93��z|O�<
&���߀�}�Z=h�z;.������d���V��I�K��A-���J{���+����{�Eu��n�d�E��sE{E�s�ې���l��n��>3|P�2�Ź �`H>E�n��N�+$_x`�v�$�d�\}}�x�Subo��Æ}ޏS����\?;�v�w�(�����#߼o���%���en���V��p�yq%�U�'hp�iFgL.��n92�� y�|Gf��%7��*� n��|6�-���ܻ�9�xg�*c��@�W7|�V�f�kw�h��\{8������`�5�#�e�ތ������M�s���s������)�nTk�������"�^��=�2��*:U��Bt�:u�ş&���^:������8}D�3L뉳Ҽ^�u��򸛉�� =s�u�ti*g��T���N=�rv���R��;�T���2}4����"b[�㌴}��r:ј�o����M�2fS90��KƸy��>���?V��~2�s$�nKdq#"_�
���G�o�K�{��tN��Lȹ�׾Ө���Q����Nx�dX|朤L�]�v/-�X�G?e~a�M���o�����{�{�#��UQ�B���7��>�އ1{��2MD"�����r��X��������c�kף6�.5��^q��C��So��'�<�E���+�,^ͦf���Ӱ��f���#���wL9S�v)K��_��^��9�CƖ}��Z�;j�{k��W�f�����h��T���x�����P��j^��#T�����g�:��9�8$��e���I�����}�����Z.����j�R�_;<��&���-��xey��v5��t��"^,�ծ
'�m����m�~���{ݹ5�δ�^��i1y�Vd�綘͜��Z�7\����KHe�ᱚe\�zz�P쥝a�X�N'�Qj�o^ygr[��a��5�ӣ�'O�A��N�2I�S����n�+�Z�r��w�KgMM%us��C�C��u�����X�x�����^��Ib��EO��Gv��h�*B����o�m�����)�ޗ~ש��T��]uF�u��u���,�+�,e�"*��������#cs3��}�teL�>��2�#���ȍ>�/=�7ޟx��x>�0�[�E��ϧ���~S2;§�Խd�5�vtN����Zʂ�)��z�/��>gw���l{�^%[�i�٩��������]���@�(�qD�W�a���P�:�x���{�'�����zG����uAtn�٬�S�V����}��F�*��Y
@SQ%�0�q�[/>�V9~U�cO9��z�<ۤ&�7y)�4F����Fx�Fz=4̲Ag!A��"�[�㌿4��)��kʞƷݳ�ϡ.�8��ن}�m���;�����'�#�^2*�jo�S�è���z�ƍ���Cc�{J���CѶ���ǌ�z�7��u���2����N2^|=Q�*:�E���^3���Ǘ��Z�.��ӥ�=fS�ݪ]o:����������v�|M�O�" �� �� DG���;����wu����w���;��x;�8����wpq���㻃����w����;����ww��wpq��x;�8�냻������ww�pwpq��・����N�;��x;�8�������w�㻃���q���w��d�Md�H�	k	f�A@��̟\��y@��T����T�UJ�%(���@IB
%EUA$%�R)TJ(�)AJUP"�U* U"J�R����j��EET����"��(�EHR��S�T	#�UP��
��UP��Dlʔ��D�Q��*QE$�7�"��UQ@ J����
��.��UD%BW�%�*���(U$�����"vd���*D���I%5��%UJ�=� rz�ZS�v��Suպu"��V���)-�5�۶۷kmrn�e��[tt(r��l�7D�@�Q9���N֔������T�!42UB��P�  ��Z�\魷\�igC��q#:���k� �Ǝ�Ѡ( Φ�(
(���e� h
4Q�n��:(��E�g�
 s����@h裁�TR�W�J�OMR�O  � �=�"�ִ\�Nµl����Pf����.�4��]V�ۚ�lQ��)����m��N;cT5W$U")Q�C��R��  � z���c��Ss�����q�@��֨tq��ꎄ�K:tջr��Eݳ��K[knPùmn�n�8���V�mK��$JU$R UR�Y�  <�n�9��';A�ݻ�u��w:R�RUp7K�pwgܥ.�[wn��wl��[Wm���eΔ뵛��r��j�V�s�wV�9�źtv�6�����aVh)(T�x  ��]��n�ٛ�nѫn�
ڹM�ݪ�v�l�ڮ���,w��)+�g;�����gT�vڷt[��&�ݦ�kwV�fI7T��ۻw[m·;e��������x  w/�V��7]c�u��jH�ݎ�Gkl�7J�s���.u��F�밭ͺ��JQ�;���滮��AFڻS��g*Vݶ��N�v�+n��:ȥA$	QE�R��O   ��Z<Wl���C79�n�ج�ζ
ݻ�]0��Y�h�p�Mld��Vt�;[:��Kn�H��wn�J�GN�u��klʋ'nj�n�:�v��
!H�x   X�Đ5n�eW]���u�����njֶ�gJ��ƵMe��R��m�ո]:ʻ6�7�˶�wUR]�;���v㫻��XwM5IΚ���T��'($�"�$�U$x   �t��:�Y�;�م��wjXӅJ��]���A�8M���[���k�M�[i���Ә��u�k��Y��Wnjum�[�.��v�� 5O���R�  S�0��T �a�OS�5=  E?�P� �?!3*���   $�T�1U5(b�b5s�L�M!���5!JP���rA�/SO�~�Z�߽�y�߼�_�B���bB�	! ����$�	'�IO�BH@�$��HHs����f=���<����S���B�L.��B�)�]�jo������@��դC[s%Y�\�wkhd7#ʶXK^j��V�!����f�u�j̔h�����/��H�ѵ����>,�k"�H]،̖�*LX��V�i�W�Lܥ�F���gd��$�n� ��E3 ���죄�ц�w,����(r���(*kU
��0�m���K+Ƣ߳j�AR�C��)�Cr^2�Ef�U�d;%!{j�g"���	�661$��t,C�swp$2�?��d��a������(�,cCm�Tֱ{���I�좱kZ�8ۊ�ϯ.R�F�䅗��-�%m��Zl0&�y�p4s`X�K)���n�ڼ@����R�˚^@�X��J�{��B"�j�Sm�s�)a�[#T�pÖ�LӀ�j�!s.�FV ���Z�Y4c����KD� ��V�R�.l��[qz��7�V�
_�4��F��; ^�knV$��hhrc2,�t��ƴ�ӊ��6�^���VQ�2���[h�8Ƴ
���ɭJ�lHt�V�v�'T3fQ�nEf����U��T�t�R���rL6�m��:2� y%���6p�]E�T�!A���˦���fHab�m\w$�
��+լ9�X�7G(S�bz��y�1�]<ĵ��Zr�!�^c�3@�R�d�%��;��1"<�[h�0b K=F��Z.�l�3�������]��ص3e�v�M�3-V*�VF�E�͕-��7k@n۱���,dI�:�OH;O���Z ̇j@%��
��f0�%X���a]�檺V��E5��p�r �GtwN��P��N�1n\͡��а���^�4�ر���m7Xb��X
�n���!�ׂ؅�L�D;�)`�otٰ��QۚX�c�NA��n�-�ԷNd`Z���~������qHt!�H�Ч��TnlL�{��n���e1�cCH]���Ep��^ն�?�i�k�w*�9�Z�S��9�F�
�-R�I^�ة��$�#�l��j:i�1ۼ�[;��XT�e��!��f�-î��6`���ē�'Qh����x�')L��ݹ������h7���$FX6�2 jd��P�Se1�uBc&�l�S]��Wb�\X�PCԔy�V��E�� �ӂԂQ��nc��ZNŢ�֦���ab�ɚ>PJ���n�VKhդe�{w���� +�k�z�Z�+�F����
Yʷ�����6fd���&�`�h�+ᩒ�#Q��E��X���^�Je] �m����ĩ�U��f�
�Kwú��KZ��B�G�M�j�d���h���i��o���m���n�����l���=�Zލ݈D�N�!GM�bQosR�z��@v�ǀ�[��/ �dH^ާ�yN��oF���7�I���x�IުEFe� ��m�!*�^������u�m�%γ�)�B�oR�m
�.�R'NK��T>W&˘�MT֢�����pa�2�t���F�7��h3f�J�J4��I:܌Լ�m�l��$Ռ�J��MVLȆ��E�{A?�������]�$�z��{C%d�iܽ�2R��	��ʊJ9jV�^*ݙ���R�݁�N]/��F�Z-*����-�[����k6�˛�I��$J�����-�ܕ��;`xS�t�U��(�`1s0��o���e�X�\���=�4�'w�� :͎D���VY��Z���n�`{[Q�� n�7v�dҶ����I[��ج
Z�Z�`x��z��(�;&��;�ZU� v��LZ�lf����B�m�8`f�ͨtS-`&膋��:IkKQ
�*\�v�4��'�e�ڍ���S��T�ˉ�Ӷ)T7XӸ�(�`�ek�@����ְ�I7K	�%��%�`ޥqi�VP����G2�����wq��� �h4J�bojl���w~{�Lf�ݡ�T�F�u�64q8�pj)�������Թ�{�"�4�t1+B��@i������7����5-�M�;	f�e��&f��{��sIJ-��MV�"!��k\���� m0��lB�9>O+&\��d�1|�aڄ��T8�w�ې	��iI7X�ܶ�wx���˦1��m|�V�6�B��)e��!��B�¶���	�`����e�m&�b�m^z�h����Ihr�Ӕ"5w٤����ѕ��D]knU���t��w{eF�dᦜ�h�y[f�djhc^�-��Zi��Zsq\6B�|v�S�[Y�.����&,Ł�� �3/-oh볘��j�&LE�/T��<��6еfst2�5J�m �ڔ9G��'��*+`��Ց�n@h����k�Ѯ�C��ӳt��+�O����[�JK] �ku	@IY�Rl�P��`Z�(��P�,��<�Z˄Z�e�H�3Sk���FU7jVj�(�@]�8b�F���P�q�7k^m-PE�ha��,�R���^,bi Ө�Ӽw�Up���Q�
���!�H9NdÂ��V7c���;P�R��,�"U�ikQ�9/��	���6��_�[X�f�Ƙ"�J,Y��l�&�⹚��,�a�5o�u{V�k̥t �[�+Q�6B��+-�(�`�A���jLu@l����eѱZ�������H�ᶶ*[�,d����z��ef8��������H��y[�a��A�(.nP�NnRrf�C65��J�0;���o&<.f�1�̀[�B�����4c�L�=�E�����(DY��8f	Pk5ch�%n�7��Y3S���K0�7�������z��Ռ(�)��jU��Ww��hd�l��4��xN���6�=1f�h;D5����<���1+�Z�l�ÉX�Z��t�,=O ���#H̰��Y�U,߆\�Mi5��@-aݲ������m����9�J��FHMu�P���nd�Bd܁;Z�XB�֢��Cuj�cn��mʓN)ԫׅ-�4/NҚ����M\˹��1n���-�ۡ
T��qhS,m�ģX�������R�2P���U-�*ͺ	[�Ɗr�T�6N�u^���ܒ�� �oC�j ����g �+Y�]&���5�5E^
u"���æ(��ژ���X����e�W��K����b�'�e0�W�Z�H��H滙ݢ��V����x�2��Q�ٲ1�B�2�⊥��P9��3t
:�;�Z���&�=H�ReZ��1ƞ%o`��B�0�ևR�,)���Ӭ��t��5�(��5��M5qY��qb[���˹v�^�ւV�DV���
�YMn@�Y ��gʶ��ˊ�Okba�x�2�ZB��]��2Ë�E��m�B�*kJ���<z��fM��F�Lp���e��P�AmQς�:���iH�Cz&�6H�����[[�(ԫ3U�,�����,jh�	��w�bU��M[�b�u���F}x�b4��a���
a�Q㫔��Ɔ��F�n���J��o0��e���h
�i�5KL���:ɨ"j����e�艻���4G�V��5�CJ:�(a��jZoAw���/(]n��Y�h	���U�Y��h,J2d�1��N�ux��G����V3�-��h���e.�ۢ�U��&�n���&����߉�`�*L
�Im*r�kBջw�t�wl�����M�,eKN�7��e�{D7J�䔄�)��� Y�4mm �FZVmފL���Ե�5Su�4ޤj{j�t�&�Zs5�C���9P��`���4�)^�����9M�k���4�TpUӱz&iH���Q��G�C61���$�5Ԁ�%�M�#�.�H�۵R�^��1�҆�	�4U��j?���7i��=496�0RY��;~B�A,�m�œ&�h˲��E����0��|�Ҩ!�Z��1@H
��-�u��`�����r�e�p�E��M�-���Œ��r��k8E�qd��#�����.���NV�RA-*�4VS�UwgE0+^
��W���],PRz�[��(=Gn-;���H+d�]�b=�um����Z+m�;�)�je$1��k	�)b� �4�m�v��Y�j��3w�mX�Q˥ y4����&P&�Y7�bI����Ū��K��:��[��P�������A4�`��0�/.��,�y2�V�[��4�����#�̭E��
u���������ͭI��7yP�/ʺt^�,AsB�9�1�d�ǲ�$f'�2V���؍]<���MP
��Y���x���8C�>{f�,Vh6����gU5yDf�v�n�;kn�N��we�b̌�.���3죥mK[�5Oz�a���okfk`&�ƕf�]D޹Gd�'	�2�f�h|�"/E��wS�]#2�Q�q��^f�$5m���qn�A��e���CI�S�)Dn��tV��SEA��3&=���-T*�6����х��rf�f"åKr�5WF��˶u֫j)���E���7�z��R^b�*��inN|�Ix���\{�w�C{��8N7K y��)
�X2�@^G>[��f�c��@�l�R�)�6��C(������Rm� �����Ռ�r�
���o.��AI0�6��̇A�ܡz��j��n-��*����f��u�=�t�;x�J*,�t�Ս�:�D�Äz�w��l���f��䧵���*T.�6�;rh�t����N;J;��=+�iO��2ȼ��c&սQ�dúl�ܸ��s/��\ʄ�V�fh{NhĶ
��ݗK��1���{�!���ʴ��f����h�wW=��0T�S��L�+�W�8�T[�%�X^l�1�v�T�.�H�B˴��O&��y.�թ��`3`�b4��6֡�kV�*�wN�Z^�Z**7F��Ɏ3*P�v`��ULPV*����IIYX)���"cƆQ7�+:�+�ڌ5��ճa�t�TV��N)��e�*(-7j�k�g�x�q`�q������dgWC&�jՠS��]�"踒�5W�[j���%��,i�V)Νn]��� -|䊹4�5<'eh.�L��IJ��ѳoV�AY�3q*�J��21����x��ۚu���"�F���
	�b�	�-9Nd���6�Zg:�]-�>(���6e��f�֜L�fjiP��C+nlV���]��Vt�4��r�Ш���v(���!�P!Y����q"5G�\��N�ݧm�ܺ�$_kM��k�iȆ�#�!�F�/H��U��f9�Wb���aU�4L݉��e[�P�P�!쵪V��ʧ�ʫv���%YA��@m�Enb� U
������˹�i݇ZCf���])YF,�t�Ѩ���4e�v�ͩe��6�&u3%�
!�8�����Y��djC#4sۻ�9���z�f�R�t-�rP���l���T6��^�zMT���+i=�ki�n\V�#t3��޹r�K�Q��AǊ�T�
i*�Z�(�kD�;�5��e�G/t��e��X#�ɹGƅ����t��i�4uL�9&'�1��h5aLg4��d�K�E��n���D<��G2L,�F;�0Y�m����ϳCr#A�,�t�,8���݅��1�ƫUj�$��]��WD0��r�̗.�1�h-Y��E��mB%If��-�ɐ�0&cu���ցJ���0⼭7p^f�63��4Y�ۻ($#���Ēh;lVPV,7e}r����ҴJVha�M�PV���ę�d��;�B��*|�*`��Y�������������T$�{J|�ŗ'��	m��\*�Əd��p�,��V`t�;i�yMڕv���'v^�[�����uu�(oAT��	o\�$Į�2�5�&�J���t⭩W�] K������q��A�����:̡Ff�bX� ˎ^��E o��[w�Km�k�̩B�nk�����CB�)�nͭ
�n��^k����n3F���u4��c�36��lMe�C�4��Q8n4֥�쬽jb۬�d�[Y4\�ۑ,{-dkڗ�h�Z�X�� �kkI�3t35��.ܧ����ן�v�i}�O-+F�7J�r�J��SȜ�k&��)���|���5`��IZ�I���+2�	W[��K0��F:���Qm̬�a�m�j�oM,��,�F=4�]k�I˵K
�so`�p�Cup�w��c5{��O��)sa�'c��Tb�G�I�Vn�{a����'jX��$Ƴ
���:x)6���k�kŌ��7@	Z]��4`��0��BY����W��v��Ukz�cU��/u 2K�PXۦ��	[�+4t�p�q*N�{�+
�pe� 曶)������2TKIb�Q��}u�t��ؕ3��/e�nG��S�d[�γ/5�l�?e'pT�ֱ��9�[a��V����	��mK�l�=q:�j�1�m� ���B�	؂�sMB�|b�����Dk6T&�+h<M�l�!�J2���ۡ$��3���é���i�v���-X-:x^n1Fehv��1M+��N�Ѻ��#R��Uj[+Q^�r�n��Z�LyJSB��_G&�(�m"N��CX�f^Yt�9q*���t��C�KJ��x���M���t�6q��$�*���M�l逇29y���!pVXxi��d��e��u����[����r/�K��k~�Yyjn�����ή�X��aO�SS��eCɼ\>Kk0+X��R�d�b�<�H�u���WYJ�8Vq��멥�4�WLδ�3�����@q��(�\u��������+���і`��H6&'_����g:�_`{B����<wl��2�J��Sa����'}�wTv�>R����̮��*PV�h�Jb�w�9J�N���M�G��f��έ��u�,ggX�N��frST&�C;{�'����N���D��s�=D�\���U�#%�s*�U�9�pk���f�w`��B+.b�PA48mE@�lX�����oS�eN���Z�ȯj�9ŕ6������@P(k
���]#��O����ƨ�]u�ӬhvY�Y-�9�{�poQ�h�� �u�i����H�<�����4f�]��-�,_`�ꗢ�(7��\\�sNh���4%�y��&ww�!]c��R�X	��$�Q%��2r�4QO�n���="糞��k���U���y�,w9��H�s!c5Z��S���.���M�w�n�7��D�3fJL�(-8���vR�M���V"�z您f�d˾�걼�Z��"�/�@�Ҹ��y%ְ ��-��b���j�w_v�`���J�btZ��г[S*����X���̷�.��t�v+M�Jպ��ͺ��˝��{�i�DH��Q'��z�u-�`��V9�Og}ԛ������6�E�2�n)ۼ
U�]��]�]j���.WQd>��R����2��R�+ �:n��Ŵj�qhދUv�X"���:&E��=׈oJs�IK�����[u˻6�S��jY-��j'Z�qpe�t.Ŝ��ŷ�m�d�����۽i��a��^j����r�ɩ��_n.��ͤ��8�ݎ����S��9�ŉ)���sZ��#�1�8w%�7:�X�M�𽤷��{��o�q@jj�G(ܭ`sZhew;�'\~�������2��W�9_fPH���Mū�F���J�M���yeoPK��-�1�خ�8��]�8sqN{�S9�
�e<j�03�wv�яS��^M]J�ڃ@0�̭d�Lb���]��y�CZh*<�г�S���n�aɮr�zv��7,>��h��coH59�	�^�o�d�ޠ��8�g1�	�\�d��#��J͑�^v;kd��W��i�x嘰l\2����qmf�b���n�����jn���픸�ڎ�:@�c�1�;J�]�zk���>6��"#���6eut��5ы�i����՛*|Q5��D'IZ�/���o\۩t{Z7��I����(HUW�aAc�6%n�,�.�ގ�|��/)� ,)˩�K��h�b�{{���<���������������\�i��-
4�ڷ9p�oǗ't�LK{�ם�:�T�q>	�j	���wu*�p��mmC���Q������&Wv�V����o�{<!�I՞:� @�{w��ڂ�[Ѭ�/\��^�b��]�-��fq�����)�5*�Pj�Q�^�׭�3����.L�k��3NJ�����!W(��ˡ�F+�;0���LG,���0$�K�J�u%��/��93(�mQ�t��H2�����=>����yLA�n�(Ksȭ���ֽ�P�7U�/:X���r���� u[9oVӮ%&�|U�04Zɸ_���|������<k.�*P��d�q'��GB\���[��ZV��`B�r�q#:u�lN�"�ǜ[.ha|�W#�l�L�V�Fp�,�fܥ����sհ��|��xj�Wcj�����1��
�d�F�BQRt����I;L��ڻ�..�;3��i��q�YB��Sx�z�b�� 6 �u71k	���Z՗�Ky��������>��*���ڸ� �an�,C��VvJ�dAԤDS7���ܕ�fL�إ>"I��u�0&�C�P5��<�����h���oc)�+v���G�����-;��G�d�Vघ�r�i������D�v�p���^+���qS�#=ТE���j-�3u1!�W-J�y���.�%�w�&��mл|7�wi��cc#u�`��΁Y��,��K�S�b�e�ەn\}�В�R�[[ϔ}۝����$,Ӷ ij�߳Վ�c�z]1��Ϛ�G����y�Km��V�+��M_�;��δ�9<8&k8�8u޹l柯l����X�Q2Rѩ ��V���`]���-^WwR�ԗS��r�z8L6&L"�H ���v��4��YVRo[r� ;�+!��d*��u|Chd4B�lo𘃩%>�sP3{���mokX�(��8\�V�ooQV�s����=����4e!+7{y'}�gō�IrzB5� o.�*���X&�jr��V+��q��ܾ�r��<��S����E��A�Gr�ɱ��S&2%���wj�9]΋�-g1hVtU��`�!�]N�F&���o�N]�#����ީ�r���ʓs��Wg���9p��bR*;�޵u��.S�[���$�j��J��ڈ�C\6��k:����ч�A�yuvY��s��j�c�����]pp������P�w��}��]��O2��0�:�K�G�s5+A��.�}dIL;�u���%�F��yEq��f*��Z6�����+���i��uu^.4����29�6������P��|���xa!�X�*�U.�/Vs�]��6(pͰ���;�W���oz�]	]�D��}����4B���d�HU�j�W&v��Jt��;�;{5��a��*(����W3����a(�\N��t�XI��gP���˓5%k"B��ŗ|�<i�)}r�ot��0u�#Y��h��t5�A�o1�i#���]y��>���ih!��bn�V��^w_da��u��)A�v�=��#1��P���C�}ۡf^}�h�]��J�%�sHǇ�8�۸�ݲa;2l�����g-���R^.xLմj��c�㫾�N`]XM��f}�X�˶�I������<�;tj�Ҝ������I���а4$�7`�����&���.�q�g�ґv�Y�\=�2	Ncכݫ2��A:������u6:��Fg<5��J��KgL��>�]QXQ_�W�@��a\�A^d��XW4�ܭ�E�M�V.7�!�y�O�X7�M#�p�s3����wʶ�dI�z�8�n��(!��5v��C<&H��`ul̾]�v�C���ff+�~U�^���<yK�\��m-�:��:���]̀x��yk�����iݨ��+���f�$R��X�37�o��Z��V>�����bP��Z(V������;}K��c�Օ��d��*}�P,^����œ�˩7�P��i����Z^p�x8����s{��:(���s���Sqnō��1U�#��l�
*�TWx3~a�B�{u��eX}��0�`Dr�Sܩ����:��Ιۻ)]s�-+�A�A�9�S�cN\�lW��,����ۥ��ۊl�\��_bR��I�oJ��b���t����n�ә\��
1��b�S���;��۠i���2�*̎�vk)J�]�<�%RO7��̱��{N󉋲�]�WMK.;����6�N�C拓)g2i���][@��m��L_&uB/�hSʵ�Ω�m��M�̹��⹄�x4���������Gy�:v\�[֟��}x��C�v8��=����.���C�A�zڣ$��^EƁ�:k�L�A��P;8����/���2��"J���u��#kjN ���]��������
V�_ev4������W9^�z+��J�� �5K��}lu�r��l8�Hf�b��q�]B胘�^���;\j7�j>����-U��	\% 96��s�<�N��@��UՍm�����������ⷷ��D6���@>Iغ<@�sl3�x����T�+t��F��s��\+z	��h�]�v�������ӽ�A�ha�*�X�]�铞�哵,}�y��:֒+h^�uf>˕�0������K�nt߭�-�w6� ����Jq�j�{�������c�:���5{P�r�ǺBËV:�n�7yQQ����si�0� ��yY���TP	�uK�����s�����Wh��+s�����Zf*���M2���V�U��V���6v�%�Ls��a/83@q�y�1nMҊUeᬙK�n�Tu��J��ܵRP�Ꝡ	{1����x[v�t42����cWI�C�d��6ޓ�]��$.�bE�֜O�d�3s���RL�d��Ea�{��Թ���!�%��Z��븙���m�5�w�����Ǚݥ�� u(^�K�Y��rQ��K=�]l>*��᭿����@׻ݚ��*�α����ً�w��i߆|N�"�ݐ�r������ך.g	7E�K��|�����l�]k<0ɵ�ofk ����Ѭ_1�Ə,�|o�N��O.���+���.�L�9����rd_Z��2��P����5��Y��_V+Ov�Dv���W�;r�����#Vm*V� mj
���7DVGB/6�X&�\쪹a���p��ض�LB�XW^N�ɬ�Nuu�#����&3�3w�1
�ɚ`=��cu6�2j���G)�"=t���y���������k���^%��Dqh�c���ڊ����vnRȲ�FO��
�G���bn����G;%S嚖徬ٯL"��V�?:`��Z[q�8����_;ko ��9Is��]m�u9��+w&,�H9�%�NӼ��0�����Lb��U�".V�"�[ؓ=�� םu��<2��(8�ԣ��G���j��
F�+�vo~b��9�F��[�v1�-Zu�ߎ���O������ͳ�;%�uwf��K=��[���G:Y�3�C�YK���孲��1ɽ\�]t,���D���7�㥲��=�tۣB�Ao�A�tu���E�jJ�(�<��Q��{+2\��ڬL���bZ\��	�+:��%]s���B�zT���yJ���fwF��=�d�L�Gp]�dx[�e�GHĪ޹�U�ǳ�CRmbPc�n۾�����ޅo;�4&_i�/"�\�qRŶ���=���M�]�[\d<�[B�G��C����fڹb�-Q�Fl@	Zr����}dQ�����o5��*�{���̴vZcɎw��gC������'�8yփH���^R�k�I*� ���wϲ��Q�D+/��:6%���'!�Ds�ze�\W���"��L_��}A�9�k�WmoDRj�:��|��v��y6�DҔ�lT7�I��r*�����q(����^�r�S�ٗ�$��e>���-����Y��٥|Y.H���D@���Ð���4���6���5�g_������^�	�$�,F��ӧ_�cqIc�qc3(���5��å}CYY\���9�zG�X�n�P���u7ۑghX� ����J��K�c��P�Y#����lm�ꆝ��3Q�û�����\D�5ؾ)�����%
@����.��7}3�fŝ��ܒ-��궞�ӑ]��q���ç�Ƀ3���!�F����j�1f������v��cD����ۡ�y+� <�>k�\��]ԫ-t�g;(5+
4b �:��ML�A^v��O�b�j'���Y�D8���ƻ�|�R�kD���C��:�1��ﱑ[>=#�Ms�!c�n���W"�����k�5�kުi��)��:�o#�c\�� �q�͘Ȩ�:>�*��P�s�f�#�t$�otV�I�J�k[�y��v@}��!�q��,��g�h�&SiFO��`[����{�ʜ�ں�ரeL
[u��P����N�A�>1Jj�� ���%4#����V����+�]���/�l��y�.�����1v�7V曅���[ ���|����h>�Uz��q�U�tK9x���	�|��X5�[k��k ��q�,⢟Vr�NJ���w¥���t�[������Ģ�T�6+B�}�J�������F��ʴy#^�GxX�U����)p<�lGV�i����^?��;$q���ڕ�:���};F�;[��a:"�Kw�Z�ʩ`��3����t
nU�o�R��3��օ�K��F��N*�e�·(�ʔ�Ţ�6���E���i��]�e�K���R
� Gn�v��*�]Zǵ)p)�L�vjM}�U� �YVG�0���]]ZQ�"�����ͨ��f:�����x�ت�e�ϭqp.*�Td<���^\�o17�����fva�Q��V�F�vF�h͚R<+�z�]]���~�|�e-��MŲ�G���YJY�lQ���S��ty����}��Kɏ}p�Azhbu}����LCM��SV`[ܺ0����w�g������+W�Lp隻�]j�ðN)Q-�2���+ˋ�N�B�0�v���$<�G��C�ЅW�u.a��v���ۧ%P	jgu����ܰE��W멊���gPM�����֞U(���F��wyG�&��4��Z���Vv�����m@o�Ol�ڡ+*���۳5����lҫburӼ-�V����sG]٤�-���Y�8f��� a��v�2Z��t �����ǵ��gTܾ�#FE7z
��>p�W},m.���Zt��dݩ;9��>�զl}�ӮS̊�Kp3y����=]Q��$�;c�fF�\!N wʠ�ٻ�����6���؏5;mh
��h⦧[��u���+s�ؿ5��^Ļb��{��~|> }�!��$ I=���w���~�S��������Ý2������� �o>a��[���ws��fS�����,�r3�[&�˫�[SO0��[�1n��'j����Y�Ł��T5Π��v��Yڧ.�A���d�^��E�Wz��#iV6�C��`��s_e��A�N�t�Av�;]��nn*'o2֪s�r#���-��aٮ�h�}�2�����&��l��}��)R���r=o�i��{\s�ބ����έ4T��sHx*���H��N0=��1�RAd-u�A�B�/bSX��՜Ң���VsR�q2x+w�u*N�}4'cB1����FD�<p�7)�v��[�Vv�J�l.��V�q�]�9|�9 ���Z�e�������-k�M��,�5�vs�trP�$FcrCJ�W�y��`5���;�&.�#N(����Q&]�W`�I����V_=� ,����P��q�p�C��3����s���L�������M��G@=)٣(*�3�j�)J�1��"�ǉZ�f��~C35�x/���oEirb�}�(�h�<�SE��[��Ti{f���2*q�Q�W�miw 	�X���w�a":�n�v���_Ė>B���ϻA��2�Z�^+��õu��n�k���WY��]�������q	NZ8.w۴���Tw��襋�+��SHGv͖��<A��A6��Oa���� (PG���╬�R�QQp:u�8e���dÖSs:Q����s�ޙ�/�V"�� na��L�Y��ci��ͤR_JX��P��'xb:�{5<ݴο���g.�:�]�;k̠�b�j�����pA�.Y��A�Y��M蚃oq`c���gAp��O���|�[�tN3�[63�@}{Ln��6�d�:����LJ�B�n��A[05��')w [�_�ә>��A�q��;*�kv�$`WoC4�Й9oW%�t&��v{(23F*��3�	 `��0��ut͛!G�<���$�B�N-����1�W;;�.
H���Ŏ+�f�q�>����b�՝�uJL�!^ΨC;;�*��0+�`�/(����m^���l#���]I4l�B�����(��䬸�t|�:pr�|>�N�p�鴯�-gT�	.��e�t�.��,������#Xr�v���i@�܍M�v���(b��t�-�љ�QFR��2����a-���B�<'�Z=���
�aL�	���-vXϩ��eϷ�өܬ�&E;;Ǭf!��P�!tT\�oLꆕ��&��a4����P���ԡ�=����b�l�1ua磴7��g4*��_���9�X�s���ƹ3b��H=�tDl��p�����*�s�e��\|�����Վy���c��O{u5������ e����[ZHPx�P�(�	]�ԯ'>�x4�t��ѩk3$b�\�ݸo;*� ��?n�$�@P�}��1�h��\p�n�<�+K^\�
���it��=�Ƃݣ0�f�ox�:����к�2�`��r\̧������5�yC���C�[�vt�r@J��#���D�EZF�+�b��wDP��(�n<�",�Г)�}��(z���*����r4�dxkM4�BC��X�fԗ:���vd��\n){���	979�F���޼�kf��_%mi�6=�oG�w5��*�;#��f앩Vq=em�f�Х�u�|&�@xj���^���Z����l�I�gM#>��ٯ�1�M��W3yӏa������`v�Ж�,mh*�<���:
Q�s8�-V����w���\]vv��U�CY��Bw:���0��os8�yB!���t��|�q���Nou�W���V��;��O6�*���Ʒfa�k-P�W).���J�*����*w.ݬ�xe�n�
F��(�J���QOfv�.t ���8�v鱎��;�y6-��b�W�u�1I*Ż.Нr�:ôN��;zR�lu
4��+0��
ĻQ��, ��c���n�;�wyL��������@qS�{�u�d���;���P��iB^r�D�k72�eZC)?��태]c1�P�`𻲪;�,�$��6��6�:����o9�'ǺZswn��w��˴It��;�Q���iU/��C���-XZ��h���e�G��J3I��c9�X����ur7{���-k��@���.zѬ��T��m�ܱ���n��P܏L�w1I����-�뷆�e �6ga�˗�ʼS���VSks*eL�7�N%�XY��{�yQ�G�2�%�P�*��78�M)�#O<��p�D�VZ��re�J��n�>"���Gq��C�vi��G�w]#O��Y0����D���%"sἮ���r�7�.�(j�;� ���%[�A^X�R���'>���.�EXKW2WP��`���+����je��g��Q���f�R��W�n+3zT�	Ҩ�VhS���0l6��۹�����dX)��L�	|���ȑ�-e��vz��s=O[ĳ	���Z�;�4T$��A%�n�%C��ѡݲ��=��^�7�֮2ضڠ,hI�W����+/o�+V&rS�ٖ�Q����`���s����8j�h�9�s+��@���"���%7�7��FQ�)Z�lN��E�W)uВTaG�c7���g�|2�O�:�ֳ�ڭ�0U��[��H�884'��	݃��E��_Gp�R���S��:����j�ꚩ���`�L��JbR�y�w	�d���sms9uj���=�m�<�̙��<�G��*o	mj�w+Z�=��ޖ��;Nv{���fY�O8��wIz��D8�NK���7�ؓ�����3:Ӽ�;�_C6�h5-��ݏt�����l�c�%�#M-�>���]�\w��ub�)�ė�g�Zn��c3�=�	����y[JNp�U�r�{[�ѥ�o��ѡJ��#=v��v�t;
���@��AJSG
�Ύr����gk�A�e���[L����T�j,
�*�_[��w�w,n�
�ˠ�
P;��Z	y���[�lJ�9�N��@	���@��Բ�T�xr��$�[s��tu�.��A�Z˅�OVc^�[��^�`8x�e`�m]&��٪7��a�ofִ��E�C��]�h���f�f�q���,T�KR����͂����V�t���Q��%���Y]��Wp ��v.c�1)c�v��wad*)N
/rv�`ȝ
�0���%�	�Vu�HJ��w��2�r��RXJ��Ҡ�r�N$�Zo4k��1u�F�w]�R����I���_f���)t���}�>�Kz�&�7H��,<�2�\|n&���jb,�b"m�Ƹo
�s/��Cţ�,���� �
�dQY"��]Σ��Z(1x�����N�����gu��W`M�i\��r�*�,-Ucs���-��c1ewM�W.�yYz
a�w��e�ś3c-<ܶ���3�F���P��0ЬaI(���蘳דX��Ij������9�Xw��Mhn���T�xɓ:��."���+�k8p�]��o��-��`хev��%d�q0�����*J��|���V48aFt�Gv�<`S��B�ݭ��l�G�}J�c�\v�}U���	��&m��ޝS�_�;1��0ɰ3ښ��m1���ǰI\�̭���-v�5��%�"뷗k\��L��2&&*�	�	��p����+V�+x�o����X{���z���ɰ��u����<wXC�уR��|�247�$��amt�;�W"ޮ��f�e�y���K�P��0��9�ys�ġD������%�������7��;�]1�8�Ƙ.}j��`ܾ�L�"W��X�� ]��=��*.�d������y�UӸ�r�J�s��C��U��jd��/#�6U�twCB�u��R��=����nP,KW�>볺س�+wZU®�'E��,#n3[r��:D��98ݛB��n�^u�Cr�u[���M[�T�vwC�o(j��c%+�Rm��<�N���K�I]z�{�����W�!���>�L@ {x���4#dѽ���k\@X�]ɭhr�3լ�ݴEw'`Zhi"rŋ�ـ�n��*�]e`K���[�K��X��k������ڻ3(���R�Q��G.���%v��YP���r�8���4F][�����T�KT��� B�Gyw��m������u�sw�I�i�=29�W.P[}Q�(N��A�'u�u{Y�p)EU�xq�e�B�X��ّ
�3�Vu &�*��ZSm9�|�@ �0�s&�e����K�<���Śn9#���+��[���75�>�+yH�٘��)��أ��+��Wn����1�[bs�N�R���٦�ӛJJ�/Y��rjm��U�J��ֱ�E�n�k�A�
!�+e�ܧU���'f��&O�wk��ݣÑ����5��+��s��:ne�G���1����q7�ys`������E�����Tˠ/�*��SE`�p�j��Z3����5���5s��u�Z�t7%gnU��v���7����e��#A����"��y,:XU�n�Sn��GXSuM��JEJ�x�%q-wvm��N�������SL�1�GH�ݔqf�"�hGw�����H�NwCϑb�o�6��]��=Z�O.��C�oTA�ye��&�՜��U%r�����b��5ګ"G��Յ,��+;�&��>���v(�;>�����^e�����𝢵�џbHoY���v�op9"9[�Of��]� }Zb��/[���$Bo�Xln�뢣�m힥
�L�G{n&K��d���,��B:���y��qWf�`�
��S�]8{�����Lf�3�Ԉ])�T"�����cp���Wv�-�V,Ksy�89��$ݬK-`�c
HZ����z�i�	��g����S�� ����fV5M��Wqg;w�n�	�lr$p��3]-�' ��[Q�*v�vj�N��]W�w4"״���Ƒ��yhbGK�-Vk��Bյ�N�t6�5Ϝ��}eV���z%y�둽봍��]M��z�y �d-��pp�9ӞY���oF��G�l0\�Pt��YV��\��"������[���g]]7�S5ѱ�%�\l�B \�̣CX�����GQ/9Z=���K�Ȟ�U���yHr�|�����@p���nVAS9�5W\n��"'�A8����h�t���+�h��tf3�]�U�3��rբkC�wl�}�6�l�:��̗ЊH^���Wq��I���q�ǣ��-���ՔՂ�t�ĐT�m�SOj���E�j�'|�
!�����}���ճ�Y}�N�w\���g!Yô���$�eK(F5�u���U]8������<�Ů��'�V`�V���.����Y�x���_��v���c5k@�\G�J����*)ѷe����v�Ie�9Q��a{�NuM�¹!�}ʃ�o�wCF�O����:�ԟ�W^{z��Lz�#������[���<�m�r�$}k������|���=K|ᬪbUݣ@ �S6�Eڜ�)t=L��"����]�P�h�J�R;��7��Η�#I
=�:�Ι�Zh�4�$��|���7�*G�{9M�SVz�q�2�:�U;3�o*Y\-.�G5�9�I�*�)������Ճ���H�y�(�n����7�.�U�����7��DL�+��M!�ݨ:+lj�^�ή�#Sdy���3K������N5�ݦ7���k1UGK��wT�[�:�s7�ܥ�=V�e��ux���#zVKWf�id
Q�(��D�GN�ۥ%2�ϒІ�c��w�8��:��i�J����CպJZC�zv$9mq}VY���^nPU�������H�c�tvM@�fI���Q����%ݏ��a�am-9ur��Rt�lV�w����`�Jr�����$PF��ݥ��f�ɛsj`ޝ.�vw?�Ts���P�-��`S��:�g&T�O"T̮2P�Ͱ�u� �֤�LMP���\r4����E֤t���q���C��̙��8M/���b!b�.��KZ�.��]�j��nY)�:�ʇK�u��x��ԗtf�ϖn�<�.�1KS�u)���ɥ�	�Sa��x�N��2�ģȧ�^�sm�]�yn�7��=�у��OEF�(��oM�(+��)�U��܅��as4R^!.%)f�Ʈ��״ 5�[�h1׶vш]����V1�eR�Tn��}�gG��ͭ��&RG��Ֆ�U͵�9����W�v+γN����K��趺���UC�3+�z����N�8���B�)��/sb7�V���7��L\�
K�w+�W�D�9A��y]1�Nі�KY��N�1�A}�'d�y0��Z���N�2�}��3���8�
��Ȯ؎A�(·WP���ј�Z�t�
�-�+s����n��d�LZY|�,� 0�㗹��\�nl�����v�z$U�ӚGU�2�wf�$����*q���Z;L�;6�H�Z��Cn�)G��4&+us�f�O�.Ψ6�e��Xo+;z����E���# �e='x�Jт�%I��Tz��4�x��e��n�1Ks��T���:ۼy��IB��r�������^���w��]{���ù�/X;L:�gip:ws��k�3[OxΆ����F�Og5'\:6N�G��v�L��UpZz�Y�B�p��yNLekA��uޜק��ϵ�RB�rf��/��<ֹ��x���ӳ��yL��=n��WX��Ś�\K����qu�2����˽]��)������׼�� !�Ǟ�օ�֓]v�yg�̠�VF�f�-��z���#�S�5ΝZ��=�����꥜V��
�QT�Ew[��Đ�5�:��w�έ͠o9�Y[Ժ����*Œ7��o��|�Im[�]	��V	��y�]ŃWWfD��+�il�K���S�dWs�i��&q�։k�� ,��m���-�nM���I�3;�܏;۽����A�~�2�<���X���{1[�Y|z��vf��p1�a���������7�Ѣ���]��u]F/#;0�7%���;]gs�:�f�W�Hfu2y�4��"���j�Y{��j��7ՠU��eM��K{s1�yH��y[ڪ ����NS��u*	<�N���7�����N�|�t�U܋����J�0|�Z�Y#������Pv��rv8b�;=�e�wpΘ:ԩ0wNJ���5q8(�"�u��0���35�;�l���^�)��3x�ϱQ�!۳�rl�I_t����QӢ����-�M�3#T�JY�Rv2O�N��oz��mc�X'kj�4�৷��EҠ�N����7h���Aʛ]H�e<#��In��7�;�3�*�c�8ggܚ-�(Ԇ���Am+�؆eԮJ�{I:�:�'�޾�ŵ��W��I���'�A ��TPDP-�h�dU�6�UDX�#Z�ʊUKi2�r�\@�E"��,PR�QP��B�%b�XV�**,QHcF)+DR�,Qd �*2��XV��*� TY�PU�
�Z¢���J��%H�Dd�YYq�T(����l�mn2����"B(E�`ցm��1�I��� �J�2��VV,+��*#
��2W1�$*E�X9aP��W.d%J��& *����j ��ZY��$�Y*AL@��d�B�
TU+����)���R�s)��ST��2
�b8���_��I.�0jz�+y˄<r���-����wn�8���Y[N���R�m"6�bC\5M����=�k�yTu�^_}��{�zE�;�p��]0��|�V�F��D ����T�ݧQgI�m�-�o;���DOT@^�{��_�Z���$�g���OB7���$��IV%�H��w�7͢�owBKg�K�|U�~-S�k�\�0�4K�w��3�*��v�עy������m��7�N�����w�jNx!�ݞ���[�+��H��I��8)�J�^S�*����3�XCE��n#�^�tϵg�7�/"������>��}���vg��v�Rv<�r��z����>�A��P_�Q^���{�ѝ{��^J��fb���mW��|�O��iz/5�t�i����H3��d��W�H�^T��[�-M�t;�_u�]3��u�2É����K�����j�ѫR���lR3ŝ�-���Gvo�,lV�7v_�i1�%��2>ڗgs�|/�N�W�s�Ѕ;�n���zw����-j��g+T�-�:����V�pҙi֖e��� םX��v0��(8{��=��@ۘ�7������g\���|ʚ�I�5���*Y5̧h�X�E:Hݏ��i�u`ӴVr�{Y������kK��r���D=�&�gd�<3v��?�y� ��c��c�zH����:T�8�������g�yӰ1J���x��ĥ/;����(Ȱ�<�JK��Uh��.�Z�5���QE��L7�S�6w*�,�˥16������s���ۗl�\W��MxȴUW��dU��l�FE<�;�k/C������7ܟZ��x�������%�n�j���b����	߶��o7$�c�#ii.�wY�j/%b׵�OB��j��qs�/B{���/6h`�}B����FH�[VT��������ޗ���J�gr���Vt��w���߅@�.�n��am>�V�)w.��_z�P����Bs�Xtw���=
�
(u.�}b����52�'�$�=���[]uA�����^������Y~$�Ϡ�g����D%����$m�ЇW��,�>������;Vy�k)�r3�czX�{��_'�=Q�ag>�dT}��ȋ^�N�.�x�)�u0�rɞ�^�I�|�o��`����J��=8K�=��U$��·�g/%>��L���r����LV�;(�Xpc@�HiY}���gwE�-��2vN҆<d��g:�k}ыj̼�A��6Jr����ޔ&�&����yA.YZ���^��=����(�x���c��q<�\(L�5}ob4ݬ��Ҭ�r�.��<C�8̈G��l�ܶ�9��kv�9jY<�bkrp��x`w�g�]����1�Dև�B��\�(^W6�!�V����ɯF_��C
4�><uy�g׼���r�vz�՞~�,�=����[�tN�? ����Ǣ�б��Li7���/�뀠�$��6z
��%5/�s��^����Y�Ah�/��7��W
�SV ;4��4����z]T;�!pP��ME�
d8���ǂ��-Vm�w���[0uD����6�DB�P���碖�$�z?0�^ L\八ҡU��I�^G�T�E�2u	�-���,kX����K�H�WU���qhp��id\�oە���)��|%��Q1c��o�J��v�a���>K�`�������1e絲[��3�n�*6�S}�V�F`��i<Z��q��лV�Gk���r�y�+�k�c�}���%9vP����=i�۹��V���Hiq�#�"�䎡�\rbR�XV�.��ʱ��Dწ�5�J�&�#���
+�7���y��<%����]�:���I/�U�������ڧ��xt ��dӪ��������z���8k��:M
�6���#]A$��(��̣�d��]_R�ͼ{����)`j[v�k�N�0s�|�l�!^�^�̹;Of�۝R��]�v��t�1�58��[D���P����sT��u1n{&C�XP�)�I�uL��d3�_��ʺm�1}�g���1?@�,�F�lv��bJ��q	ޱ0T*]{�Uo�f/-�%�I�kW�N����6�{7�Y1�5�u���JIp.(^�ܢF���j�<�^��C��z	/���!�����{���������N����Kŝ��O��M	Ȗ��&�u�;�%]�eΙޮ�ʭ��EB���1�1Gʲ!om&j��
)�o	�k��<C�_ϮF�{"&'��M�@L���y���Y���	U�-��I0@��5�µ&Mu���#�}�ix�W���8����o�Uoi��o�jg�)U�,p��|}�2R\0�����-mqKμӃ������+�z/j�[��C�8��������6낇K]��e.X�s�����{�)�agx�5C	7����V?D������ẗβ|�>?h�Ĉ��Y�0f#�R�{zmu���+A���$p��K=.a���5Q�qߣ5��L�{c:hDl�;�U;��Vz���ma��!X.n�Н�s�j=�6�����U�ǈ9����F7�3����3���!aR��X/�9���/�v��(V�fb���Ou��K��/�͖b簣���N��<9:f�*�8�� �m��7"���˩ցw}"b�0�Kn���������5�}�ɋ�q0�����>5�,NWs�̀�
��Z5H�ݣ�YPx��"9��nL�x:�4��L��0�_[ޔ�y�G�����}j��=�h��t��,�5ΔF�\a��]��փ����J��{�rr��k��qoM�T.���@&T"������٦W�W��u��3@�={���@�f�1�������|3�[�ӝ�*Z�˞Y�*_�6�/�,Pk�k�������B�m_6mRΔW>�<qg��8���_zڵ�g�z���R���{�]\�t��D{�ů/�D��-������A�s����h�V^V�9ެ�/½h	մ�8�La��N'�0�hu�����U"���E��#,oK�O#���
���	v6��Y��­4]p�&k��<K��񢎙��j�_�<e�H�^��W���8�4続S�y2��y�mC�q67:w�2��&�ñ���"����}/���t8��jS�X~>�Л��;^O��Λp�Ե�J���wb]u�wim5%���%�㎭�ڐ���fe�"�E��y��k5�\`��2ThI-��.�>�*�Tڎ��e��
/9^RO���ٹHAW�\�
���5J�l��g�E��;�E^~]�����p�Gg�ϖ�J��E����	��b�>�V��ӷ�H��S����;�Ls��d[a�e�n⼡�<�ن��&7l;��Jm�"��fq�/e}|)���]k��Wc\{`M����p��Ӯ¶k�u��p���Ƙ����0=q:�/��3˖�V����Ffz��j��AW�����L���1˜:��P�'.'_����kG.Z�=�}~� �wm���Q>4v�(�k�ֆ��u6|��߹N�J��QVI�I����l����I��N/���|�����`����P�R�VH�b�^�<�6�϶F�s������҈���0�Pc��b�pb��<^t�:����6[���}�;�\Z�NI��gb��*�;G&���$zD�Y��ܼ&��n����;������Z3�S��]�g���������3�Y<�}���@�=P�1�6f`wX�(�Խ{�bZwR-F^�i����,�o�=��C��#|�.^��Q\���Z�hNgf�)�T�p�u��ͷ��yO]�טj`����}� )��k��d���������� ��=�9r�{�79��>��3���u����I\۫��^�yۗ �5�95	u����־���:��I^�^���9{��%r��}IxϺ��sL/�Ay�j�f��.�����v�ـЩ$�n�n���y���{�c\Ǧ�ghb�ȧ�o#�]&��>�9�K����׎�Q)�_k[�k��OP|���<��
�Z�[A��5��ܫ�
��������;5�˵I�o(=�t�s籛��.�z{b=������9U��z,�Mz�^xiGW����\���wg{��Ж-Ni��n���Ytѕ|i�����1Z#�\=6W�F�*m7�m�u�}��{���e�3n���,v�h{)��>�"�*�$H��κ�{�1��0�P�:pǛ�ri��v��"�u����%3n�1^���Sz�VB�ma�����'�{&���V������Q��չ\i����9���+����e���r��W�o*G�7̮��-���5�����k�to7�2" ��İ��w�^����]�bRZ����㜨��I�!���>uЯ��3 ��u7�����[_��㹋}�g��{�ٞ�u̓�9�lU�����/�S�t��F����_Sדk�S��<��D!�`�c�s;N�9��������wJ�U��+�2��Ὠ��3��j��I��=�a<�<����_<}�%Ly���Be��{�1ֻ\�\8�\�j�+b�D�k<h{�R�����Rn���lw"�e=�i�� ���T}��Ć� ��,J]���s�q�s���}ޫ%t��3��Hn�k��w��p<Hr�T���>�e;&���������jk�X��헽<y��q���Q��^�;��7W���s���=Է�gi⼖�r�>�S�=@<��
lt���v*�-h��َ��s;X�/����ļ�/�5yQ��LX��4]N�fYӵ�z]������w)䏖�iz��K�j9s�I��A����uF�b��)���[B�<Lj�0��������(��E�0��!ݫ��;e� $�Q;E;��(��[�pc�"B��4�k�Šk{���1	5�=��ji������銗������o�n�k�dC݉�G��?�{{!
��y��u�]�����4%Ev8���ٗT�-c���o���%��D����m�nƳ+�
b`_<������O�����2�q�V�|�]�n�R�W���H��A솂��E��[<��NG��ӏ���g>�x>�1��~Y�����\���z�͔�2��%&�/{P9�w��z�F��(-��v�u��sZ����Oq�́<��ėf�+��/�z��y��ْ���tG��k�s��mԙ�f+��튞��W�Nm}s��R%�NI��"��'�y���<uZ�=�R�G�S�^��p	S�E�sr� ��
D���g�z�
k�UG�����kd�ꂹ��D.p���(��z�� �A�:KE��������iY�f��M����sa�Ѫ�O��+��U8��)͹�(:��ko���^x�G/m=����'�'2�3�î�R��ͱ�]�qF����$�x���𛷑�.��ۘe�S�ȷ}���MB��ޗ�.]�6���һl����?���0��3�����ʶ���;]f�ԏK�@�|w&�7s%C�5�ܫ�<�~&��~��<2�sh{��w ���NǺ �p�Pj�"����;�iһ��G1�p%Y�[��K7���])�ys�%��mu�_z^]0����ֺZ�W�Uk����ln&6\��A�eqGg��Z�i+�m���W��Q�DH�wOuS�����Ab�\Jh���c7'����Z��G9��*�#��̳���|��K݆����ϻ5�V�����Ǹ&�ۧ=y�7�*�k���+���[���}�Ɠ�@�al����Ӿ�A�A��(3+�8��ϓ8gm;_1���=튘��s��C}�#k{眧�c��h��r緶ޙ�'���,W�c@{���A�h�Uf�9]q!��4q�%�	�8���2�u�l��^H�*o%^�K�Xk���Tx�Ա�:/��������.@&,�MT�c)b������z41Ԕ��2T_cˡ¶���Y�8%'{��U��9�H�
j�n浽qn���o�['���9Pt; z�����*Tr�]e�Ի�"�q�,�s��
.WVcq�y|H/v�t�;+��8m�7]I�Ȟ;K^��|�%͐��f�)����x*��K�\3�J�GG�U�<+��&F�.���/�b�v�$��΋��J�cJܴ).��3x,�<��{9���Xe�螱92$�Σghh�5'e;�8nQ9�-��qXy��.r���Xp��6�r*��"U�W[�p��s�[x!��^�S��wCOx\U�O���Hf���SjSS4��<����8�*8Q<WZ߄֋�IK���5�k%��`]�t5n9���ÇdC��$���s�U���aA�3�+qY��n��8�N�tM-*L��=z�2�,� �ʙf����}x���r^�0�à6��J�-s�o���[��-֕�����C+-�Q�]�C�±���5;Mwje_ g^��˞�(����ٖ�V1b�XE񤓽�ۄ��6p�2�
��7]4�(*�I<�o�4��ⷪjU�8�S$���9��oV�w<�=c�:�k*�=��0iF7t_�k[��Zh�v��#����!����-KW��;8�~�`v�{fvp�ξd;�Ҵ�l���@:��:��.���0��Zu��㙯(�1}K�4���-%�̷�گZ��ү��¢ Uܳ�G]2��] �R��(4��V���[n�'���>�X2�u�	�6�����yݚ�́�j&#�G]�B�r�rٯ�v����A>Ynۭ\�P�O������s5�]u���[f�X3-P�/p�������[��:����I�{��Zd���)=��"�t��^^��/I���K�K��x9�c;:J������A	Y�h�n�ҕ|ܨ��E��i�w@w3�n�<���W5*���Φ �T�A�%dѢ�<�Y���S)$�I�s�5���\�s���j��Sj�$g��'��+�3r2�NR�4^���
WB��-��2�[&쵅R�8̓2ۅHu����ٮκ�+��3���Nt����RQ :��ri�w�����V�)�tm��2G�-z�.���dc#�Y4vAݎ�u��Us�|#�4��p�w�������f��C-Wt|�ƅG�ǔг[xz��w�����Gud%
F�-.���)��Êk�/VWq��-쥓55���-3$ 5��]c-�f�RS�'x�G^�*][���iPo��c�R�s��}����Hn�7�\yɕ�cڷ����Z�zL%���?�<[8=�ݓ~_߷��{��}����Q!X�Y%a`�q3,�mH)*��Q`,*��LKi*Lb[Y�
ʁl�[AIQdXUH�J���[`��J�j
T���m�Z�i1�*V�Abʋ%b�mB��"�e`�Xe��V)+[`���e�b�&aJ��YQTP��*�� X�m%�R� bLd1�!��TFW9�B��Z�Y*�Xc�Z�
�ĐƠ��"�-�Z�R*e�PĊ �e@U"�"0U
�(VR"�d+R
EiU��E��$�Z �KH,�TJ0���
c�HցAB�_==7�Õز�aP���띔�7����]�P]�3�������N�#j�wU�Hj��9k��
3���Ki��׮��0�������+�;eI�9���#��� x�@�p۱Y�e'��o;��j|��/���c��r�ʧ�o]H륙�k��M]��[zn�����<5��|Zx��kw��s����T�a��UK����!�vB��k�X=��Zx6 ��r�u��&n?mSnʤ�/c�ǂ
粄tN����Ow�c��u�|��C�����:���f��=w����n���W�]D��g�y����Q{��Bq�#�~	���W��3��$�q0�p<�)�k�mh�9D�5��{A
F@oۙ�"��z{���ވ��q�1��g}JgaǷ]�� �P��_�_��z�K��:�����g/u��+p� '��6"���c��2�_1��2V菎r��I[��:J���e���:D0����mG"ջL�gF�ܝ�{�[�QU�Nue,�l]wrwr����\�h�kz�[�5�\l�$�i��@u�OK�5򕎱����ߓ̡���2�����ߠ�uycĦ,v��L��-ݭ�{�����.�Z�\Ohڗۋ�Wxw���./�XD���m����|�c��ek�=�zE�d�Sm/>/t�F{yN�j9Y��q����(c�����ޜ��yWH'�ΧQ�`���ޝ��ͺ�������C�M{�/����Y����<��)���y�ġ�t���̓94�GF=�}��iu�x}س62�6 �ۮ�V����aչ��Nwbq�Q�o�Uz�X1�=�p��o!�sU��������q��]Xw:��b.�Ì�1}Up���]pZ=_:#����|��Ne�f�s��Ҿ��4����o�~�������#��ϰx8�����W�eKj�nl�*�M=5vdR���x�U%H�tN��}ө
zV����o����,\�w�hjs�=O�2�܆�,&��;��؞�Yk}�A�Y}�p�V>(�0�~S��F�nznlGݔ�l�/�J�k48�Pu���b���D�� �z��[t�q97t�i>�g;e���Cgve�/�^s��6m����,�H|����W�v��$��^�ʢ�����l�E"~�[��ֹq¸�j �$뻋=X�C��T��a4r;S	�� �)�k��ȋ��NF�w3��1�y�p=:��IG��Ĺ�|�AN�V�ޮVxK�a���#����uwB-#=pLyW5��������[��w��;&�5Ht���=�繞.��Ͻo>Z�����V�>�;�ZV���
Z+q��3�'T�Aoo�z�>��6�<���J��Õ����Wjى�ɜzg6K�o�J���΢���&eZ�Eо4ײ-L�p�o_l�ˑ�\��>X+�����N D�ηܫ�4Z�u�uhf�y�	�Rr�������ham�x�{�n[��>j?o�o���u<����Ī�l��^�*g��{b����(�L��J�I�v���{]l���q��/�g5�>=�Dv�tv�+㱓� �w���w��Λ��`uxT�*9t��9adT�Xr	O&b7�ri۬.��X]J����
02�u��8w��+!�i.G ɏE�iakz򵢸��z��`V`I��nՎ�wЗh���av�H_R�Ҷ�u��W��ڷ�q8���/�t�.]ɾ�+�u��
>��Dv�tG��,P\^�k��^_��9L��ׁ�޷�k���3^N��s��.KV�$�u�7�'�m�۞U]�Pq
Y��"�`ʗ5K���x%Lw�sr���T�� ����^��W�t���cQ�wuy����|�)G`�{9��5����MUMtVop�򐪢`�4��O=����4�Y�Iqٔź�4!~�yU�b[��4&��EM;&p�^�o�}ȳ�G�\�M�U�{�N��zd�gv��Ѐ�<(���~�/
?}�?yRW�I�}�,���k�2OSS�2q���ǩ<IĜֿUw�k�3N�����t��v�l���.�OXT:wxu�b~�u�h,NwԜI�*��>d�{�I:ɩ�2J��9��������,:�x��Z��k?S���y�;Ϲ��gCq��|�l�'�:�������.���OP���Aa>C\��q*^w'�6��T<9`x��'��g�'4{a�Y:��߹�^�~ߞ�\ۆ~������a=tɴ��XOS�jyCI:��kx|�2q����'�u��/�k	<C�jo�:�d�3�}�Y8�	�;�@�'�Rzj���F��Ͼ7�����U�W���w��O'�+��ͭ��a�.�t+�ly�{���,��YЌ�|e�9:��o��<mѝr*R��������|�Q����-I�l�srsb݀��3g�n��Z˃y��çCun����܍us)�S�ut���䃷O��/��F�q�1���C�q�I�,�$�+?j�Ru	��d�'���>C��J����:��?d�i�xϹN�q�}_8��~����#Yls���͏��{�l�d�ԝ��$�$�њ�+'��zԟ�u�	�c'Sܳ�&�T��Ad�����Adѿp�'q�5Π>�}�� �������v/�6��}'wy�Y6��xw�8�z����̓i'������hz���CYd=O̜MLd�!���C�,&�����N�`]jy�~�>�m���%I�M2�O{�'X~��v�u��3 ��'̜��N��nwY'M���IR|��-YY8�"���q=�Ld�!Ɔ�����+ț_��o�޿}LS}���u�����w��ܐY:�]�ߒu��N����M2t�܄�6ɩ�d+$�?��T�$?�hVN O�jʵR����?�f8���@��̎�$�'����M2Lu��d��!��`z��N�C��p�'Mw6��O̞k���x�����'L��aXN�|޵�߻�=��g��}��:J�����!Y6����q&�m�I6����7l��ߔ6���C���&�P�f�q��S|μd��{���'�4�������{�ᦆ?�i�Z.'Ӯ���a�����z�﵄�(L��%d�VO�P6��6�aa8��}�Z�q��_Y:Ç7�'^!�w�M2z�o����o���}�����߷�>d�'��I�~d��;?wu�5�`,��~�J���8²m+%I��o�7��q���>�!�Ru��xs�]��vk��٫w�{�3�����s�gM����vs�<a�$߃�?2q'��C<Ag���P����2N���d�*I�^0��|@�Y8��'SS��8�y�޹g�J�)�E��c֎�w��������WV�i�����a��(-���iګ�T��O5R�PCj^%y3b�����o3�sF��V^�]Kd2�<����R!�Ζ,uq�:�t��|��ư9�u8�|�Y�O-��}U?���o5�o��z�ɶM����Az�L4{�u�bV�9�Xu���;�I8���l8��>�p��ԟ�k'䓉7�%Ւq��E��������3�]}þ����+	��i���d;�<}d�zoy�i��y����ϰ�$��d�N �5���'>J���T������ߏ�h�\�9��g�4s���\��$��(O�|�2Ì����写:�~<�S��$�M}�=f�8��sxI�a�Ө,��S��J�rs���'�X?��?s.?�w�0��罻7��b����?I=d׾d��&�8�a<}I�je��3��,4Ì&�O��'Ru&��I�4��?}���:����B?}�6f~?���n�����yc���'�Y��Xm���`x��'�k���N�5�'�d��Ĭ'�R~g�g'�S��:Ì&�XbN �o�'�u��=߳�����{���^��׽��M!uM��I�>�6ɿl'N��:ɷ��������d������Y?0��!�?2u5�q�z�?jÈ)'u��_��K�?q�Ž߼SX��� ��!Rq��Y���N$�~ì�	���&�M��u������d�d�t���u��7C䬟�q����ϡ����b���~��4?:y��k������1RL��zɴ���	Xq��Y�9������'Xl/0�'R|���2I봚��I���f�J�����w�A����{���? �����T��OS�LI>Cl���SL�o�C��J��ԕ�Y:���{�'P�k�;�'?2w��d�'���̲>K%`Ѵ�u��G�Vf��M~x���vs�IXx�~���I��!�d�h2��m'_���4�c��d�C�s0=d�'_P�wy!P�~�z����b��{���=�[H:5ƁG3,ʈ�¼A���#�ug��5z�O[��(�z�#+n��j�ʿ>����j�V�=r�ǻ����T3iҲ���a�y|(�-�C���dj/	eQ�b��Q@�7�	�C��F��}�'��S��(]����]g*��5��������������s���o4�I��2l�&���d�'㟲J����͡Rq'�d�N2u50�M��~�y��i��<��2u�!�s������{s9��������?y�}���?$�=�6��O�<�rN�Y<I��k�	�i�S�ȲN!���*
>�hVN�d����&�F�M}a��N3G{���o?xk�y�~ӭ}��~ۭ����n�x�N�ɶI��<��4��	��:�����I��'�4�5�	�4�����{�d�*I�^$��J�P6ì�=���ϳ���>���k�I�'��R|ɶ�.�4����d�z�r��u�p�1�l=`w�+I�;��N��&�|�XN���*�����̬����ds߹~y}_�%d�X2���2q���a:����Y:��>7� �d���I+*s�:ì��=��'R9܂�z��{�*OY9����ϱμ�~������Z���I�N�����ݑd�2��&����Y8�~��Y<d��� |�d�o:�c*�αd���u��
�+���]����r_��u ����� d�T;����N~�0�@ެ�VIߧ�"���N��Xq�x��<��N2�����0�OM}�>M2u���u��@��XA�ϑG��֍���>�$����Y>J��l�'=J���V2~�Y�$�&���_)>d�<2����I�,8�<z��P�N0���������}�v?[�ѬCs?3S�ﾇ��=As�I�>a�S�,'�߶q&�Y�w'�6���ONP=d������I�M{I�Y:��є&�Y4�2�2OXEb�s�\%���f����ԇ���}�~�i�O�Y<?{�|�q�~�q'Xk���i�x�	�d�N2��u���?$�TXO���VN0?Rm����!:?�l��s�o�����l{8����x��Y�噆��۪�����@��M����g�k6�g���ߧ��v79ӝ��C%����t��{�L��s�����Iz�)_/+�6b@M��6�Q�A��%�y��F�E���YS�ڜ�}�k��^�XL�}ޯ��W��&���=I=eOƬ>b�3��Y8�ɭ��|�:�<�Y	�a����i��7�:ɿl'��p�'Y6�����}�r�	��:�M�����V������ed��hk,�����k,�	�*~ՇRO���'R�7�I�N%Nȳ���?a�l��<9�u��W���Eq2����5��?wճ��w��O��O��I�I�Fk	R|��l=J����l?$�4e�I�La�o�[�q'X�¤�'|���r|	����l�~U���{��ſ��n��&�v{�ݲ|��}�$��'XVI�9�J�ԇ��Ԭ�Aa�-!�I�k.0�I����u4�?:��8����7�X]�)O���%_�{�w�FO4���ܐP�����'?2y5���<I�Մ�z��ԕ$�����V,&}M�Y8��H|�:�d�a��'b���Ef�s��Q��F�o��_߫�>��o�!�������}C���q�ם�ox������:ɦM�	��&�k	XN!��쒠�2}M�Y:��fs��~�r�w���y^�Ğ�m;��z�l��m�I��dﴛa��ì�׌<��OXMo�q�O|��|�:�d����w$:�I;���8��k��Oy����ۭ|y��]w�{�y�*
��T�eI��Rm�����u��~<��2N&��H/̝C\�N$�x����L:�9�{��'|��;�u4��6 w%'s�O�Xz����@>������O��d�*I��ĕ&�Y?e'Y>d����a8��|ɧ�N�q���^2iO����Xh�p�'RN/;�K�&�_��z$q��9ܻ�/��w_W��r
2z��w��|ɮ�̓�5�2J����vE�~X���'̞��a�N2����2q��@��d��{��ʷ̌;{�09�e?��3R�7l�.�y8�m.�*�5���ē��[�y��Gƻaz:펢���0����-їk9�=��գ��O�)oݕ9GAȕ�������E�P#��2u�A�b�Ďt��KU�1�@$�}�_�s�{���2LJ��5�I�	�5�a�N �4�AC���a��)=d�sX~d�a��2J��9��E��R|�~��I��k�2q���}������G�-���v�k�#�G̏�{�8�̜C��ΰ�0�st�$��9�d�\��8��T;�B�����d������+�$��&�Y:����/=u[������?$�>3��0����z�̜ağ��<O̜Ay>�z�P�����5ϰ�'�4yܞ��O�P����~�Y�I�M���sZ�3�ͻ﻽���Y1���XO�i52Ì'��jyCI8��kx|�2q���rO��'P_>�x�P��ru4�>g�>ì�J��y��Y>����7���뽼٤������#��~�/qQ��~�I�R~d�VC�q��{�q�z��C�:����C�'Y4�$�2u+<?}�8��js�N��'�u��[���xw_W�������]<d���Ì�d�Ԟ�̓���Y���u��t��'�eBz��Ԭ�	�?!�I��d�&����8���ß�3_�\w}k���k�y�����a���s�I���'_M��8�z����̓i'f�J��AC�VN���d=O̜Me1�|�SG�Aa6���6��~y�������{���=d�V<��6�l���������]��a�@��'����I:�ɩ�d�a6�3Y%I�C�hz����#�=����Ѝ�̝D�X~��ϺϵҲO��t�&�'�S��6�Ԭs�P:�ߨ}� �u����Ԝd����>v�L��܄�6ɠ���!}}�����I���x����������B�i�m��:ɴ���>I�����I��P�'�Y8��h}�u�i'���2x���ɮ�;O�W�_�ʾ� ��~V��W��޳�:��zZX����\(�PmtO�s�a����u�S��Z˾���<�>�*�<c�F���\ʓ����a���i�+0���<�qooE]��=B*#��d�ATmD.�u7*��i�]ps��Z��X��v��ztI˱|���ź�����x�5������eT�8�W�+	����%AB`yfЬ�Aa��:��6�RM��~>�!�d�g=��N��;���?!�o'>a5�gL?}����)"c>�s��bF���c8ɦ}I=Ơ�Ad�C����2}x��u+'�m'm���q������$�4s� �2u��o2N�C��������[~����5�&�?0��>��M$�ý�u�d��<?wu�;���8���d�+	���
ɴ�����d��j~��d�?{���:��=�~y�;�Z��xw7�d�0�w�>a+6�S���d��{��N$����c'�,�����&�|��$�M�$�RL�^0��|@�Y8��'S4~����\*l���OՇ?Ue���W�G��&�=C���Ěa�~βLJ��9�Xu������N �59܂�=Af��)=I��~I8�z�]Y'��x�aFK��@{�۵�g��]��_��>� t�'M;M�������2x������Y���p�y�I�X~��u�c�7̝I���ܞ��'�Xw��I�Mw��:z������y���Y���Mj�]$�zr��������$��5写8�y�=N�i'nk��4��/�7����o��LN{N�q+��~��O�)������S������0���Y?���N�k�2J����J�i�'�{�8�|Χ�?0�	�kx|�d�N����h~d��~$���~?�v��g��|����H���i�ɴ��<���z����̟2}��&2q��OɌ�O��x�&�Y�I�T�ՇXq���I��_���p��4��u��m��2w�}� i�� ��N$����i$�7�:�Ϭ'�~Ì�d��OMX��?����u���k'�CS,�������8�=J��o~~-P��c�� �k��3k�6%s�4� V�L̥����(���-h.����A�x���B�O*>E�K��MJe󝝣s%+���8fW`��o��	��
}�/4�)���p�W6��U�q�&*-s5�L�w�	���6��.�71r޿����7Ee�NB���`wcpS\RG84cဳKtѰ����Z�m�rW��+�3�8��Ԛ��� ��ה��SV3���h���W3�L�X�Zҽ�f��v6�J�|S�����W�������yX-3���U�_gu�;� �9���*N�N�4mds��=m�_��i�EZD���To�ASuxr�k���Y�(��V�+}��pC{���/�:���+�:�|7TJ�`��}�R��^7\(�5��O�XV���lv��0��r�\5mG�k�ɥ���'k���1���Ζ��r�1��*���b����ut�	�]g2L�?"��+�}��m��:�\�y����S�=�	�iDl�Wܩ5��s��"�+eJ�Ҳ��w
Q�'��=yWq�V�9��iX��Y,�P���3LiFo
y�[�0󝵑ڰ��ňk�DM�MN�W+�
���"�fn���[��Z�*��0��:�`�v�ٜ{��&PV�t�h,���F��Es2�5ج�ܮ�l�R�J�ϫ�n�il˥{XV%�"�8@	&����86�X;�n�w����Vb��1⸵���l.��V���X���#2Y��z��������J:aU�岦M��-Ul\���w}��/���>M��r9���gD0���	0}M�y�w��gB�1���Zy�C�:g��y:���)3�WN`�ѱ]��|mb�)�hQ}�C�y�)k�0R����nR�g�}��g-kS���c�6I=o�ԙ���q��G�wa�4�5>\e؁�7���p�LQ*a"�ݜ�sD�l�-��sݒ�����1R�t7D�v	�=�B�r���^v��A�c���w;�wۄ��!<���ըi�	���m��#��'T=x�Y��G�GU�Տ��`j�LyC���;���J'#��|5�X�%��=ѓ4-xU^��Tɨ|�X|�H�
���+ ֻ�ww�����ǭ٤ƊR�u��ʙ�E��A��������<��֧�f��Au\�x�vA`���u(U�}[;�5��+�����UvDP7n�*��ъT�\&�콱��Ǔ�u�"R��߲w<�}3����4w]����1AZ�cɦkȓ�}�>���3&|E�4����4�t�n�,��]�f�2�f��/�i_5����#��|��,l��}�"�(��芩�W�j��nl��X/x_1��Z�S�@��8;�x���1@��X[��
[W����;�	�|�%�C�YF1;^uգX�n�LWl����/�s��7f�OF�T�4��l�QW߿o��~���شek�j)X6��2	��Lq��)�b���X�����IZ�E+�U��«�T�J��¢��h� T��"��6�XE��UT�ʒ�T+	�*��2�*B�Ym�$&$&"ʐX
-dQAB��P(��Q@R(��+Y
����-H,�YX�
2[B�YPR�!X)V�[ej�b�(�ъ���V,RAIP�ˌF)���*�T%���P��*V�D�L�
�V�UH*�	�9l�bQ��QT�,2Ь�VAE��F�kAE��Z��P��"�(��X�FeAJ�-�Ib�"ʁX�*��P�"����s6��j��q�gW ,sT5^v5	Kh��Ϡ2�u5/zPj����F,RdΎ�ͫJ�:6�v���Z���p���}_U����ږ~�������P�OP?�=�T�d�Vh���:����L'XnӬ�|a79��	��&jɶI���VN�77C䬟�q������ۮ��Mw�ٯ�����2z��q�u�S��RO�U2u+�߸JÌ�J�s(C}���N��y�Y8���O�Y'��79���'�u��Ǿ�\�s����/�vJ�L�m�d�O���8��M����|�Y���M2Lto�C��J��ԕ�Y:���{�'P�,�Ԝd�ɾ� ��O?k?so�֜����gw�y�>|{$��'|��O���%a� �XT�Aa�i��'SYLa6����`m�I1ѿ��s�!�3�N2u�{���O�ם?z�d+�;<~���GO�C�ȏ�� ��M0�w��N3L���B�O��d�(M}fЩ8����m':��Y&�B�����~Ȫ~��f+?�nCy�9W~t�y\���
IuaNK惦��0��������������<�ś�N�s�v��m�E�`��Ñj�"���W��;܎'bD��J�c�d���t�����>�%(��{r�����3sMNz�������M���;vL�r�wV�~�m��:�݄�#�e0�p<+^��J������9U��v�u�W���7ݲ�zx�{��:�̿{��z��c�f��H8K�E��ދ��J��I)�|IX��0����-�,f�;� N,i�;Ӥ1��x�R	�o�Tn?��oM����Ք��V��uo<�n���]����C*3z�q���Z�{ê�ܒ橃g�I�b$z��}_}��t}�/ދ����S� �^�:͵�.!N�}i�W��|�Tι�Լ.$J�9iܗ�=C�u���g�mb��/�+o�ʎ󷀱��t]�U��eפ�o�bؠ�+n.�b�e\����hjƾ�2/v!���.'"�o�!�}m����3e|��.�\+\~����~^�XvT��0��S(�Z^���ϔ�i{��

������w�w��$퉪������%M��5y��Yq�L�i1�
��P�.t����zo����lu(g:��;�E�M������{���l_
��se=2x��(Z���s��zc����̋{^���tv���|v4=�hj����.���/���+��:��������� z�~#x��\�\�<ؾX�g�����ST�Nd7:��ѯ�s��rZ�9/�.����U��4d}��C/�F_TZ�۶n�S%j}�[X�o����8�����e�0�`s��Z^�n������nue�	L�g���+;�G��{V_E��<1��"�.u��+ȨocU���l��6����
&�f�b�v핂G��快ﾡ�Bf��ty?���xk�����nT�~�7/s�qj��\�}��A�+|��������=�{<��boӆt�{�O��^�I%P�,�nͮ�}��&]�n�.����\����o/��]Y��hYsTP=����$�ēW�T_;&p�~{��G]��å��~7ެ�3Xi��#�R&���c�>E=%�yOH�{8�pU����D�\�ܝ�M)���pNc�b3��O}�qϲ�"_H�����u�1lY�`Z�.�9�n&/�y�ױ�3���7�ү��w 2r�W1�\����y�ӥ��y�O���c4[̻��
twث��D���I��JϻP����]��h\��1��
�D�89拞���~��2C�^��Ms�>V�yC��C�Q>4���,�%�^��xNq�<�B�x5�Q�N�0���]����fj�����YW��v��>�P߂�ɫ	Ť�ϰ4�s�}ƀ�f�����\IbU����Ӽ���Et;�A�;��MhT锒�s�Ŗ����${�ArR�����I�����H���r�}�����\߽'x�?��r�LjOd���Y���>1�^�a-��ӯ��s���MmfW�ϓ�PL� ��I���L�O�Y�>,zG��iu�$=/���vO����˕w�:䛟l�S�U���q}(�lڅX�(7�9feN[�7�{yu��*_uG�k�{�dy9�u��kE��b�"��լ�z�N��Z9N��y�1�}�˼ς,М���ܷ�L,���z� ���q����y>ۋU�9/��#�k0�}�{�x=7��k̘UN��<��v�W��ۑh��e��}��.u'��˿G;T�֣�8zy��MNfw�\v���93e�@;'Y������v2"��`��	;�d����;�K6x�'����tMS򞦢�+��B{��� �Q����ܭs�.�-�eG�	��z����s�P�t�g�z#���V�ot�����*r;w.����W+���^V�u�M�V�էo-§y���׹ە:X���C�O>�F+��gY�m�昖Zv�^n��������9��U�#�n��ZV�w�p��'CK�X;�w\����> >��y�q�пͫwǒ��G��|��NYV�ߝwA�ǃv9�+i-Jf�dN��^��+�n;�E��MvԜ��_z�K��Co����Ϻ��s~Ia��>�C�ﻎZ�+�?&��������C��O�\^q]��=���ہe�h�ƚ�T;��g(�����9W*f,�`C��q�΢�;ӲÓ7ˡ�4�8Ky�2���H�Qw��~����9�
cա»e[�����v�}�v����J�늕�'��P,ΰ����l�y�ޙ=��J&�����׼�[��r�g5;�r�#��G4��{����{����<({��+�W��*����w3c�7[�R[�V$iDu���_����O���,;�ex^{V�;���	�J���uaI.�)����#�����J�'h-�N�g��j�.�]��s[�m�G!sS��_:t
�J[(�w�L�=���h������ׁw0Y��v2yb�����rA](�һ�[�U�p����y���v.����>���0�Ѻ��8��I�V��)�r�\s��U��W�pg��U,ut�O�����}*c�E���%b�HD�R�7��ݎ@�u����4р.ޫ���͋�|�u�}"��OpHkrn����@gh*��z�ׅ@�7���M����Y'A��a4܎�2�ݪ�3J5F�RPe��s�4 �SY7�n�x��;OݟQ�#�?9�{Z�o�tU���Z6�v����$
�V����':ʹ���n>T��s7�.�ϯ2�_w��wd����z���s��p�W��&pv��O.Im{5>�yEns���9lż�������ʸ�j��ʧ��+��)�g't&k�Xu�/F1t��[1v�.�d�8:��s���nզ�D}�=�v�z���y�f�P֯�����A1�Da�p����v;Ӳ���[���v���5��c��Q{*�cQp���۞?M��c��Y��\��a_*�H�J�u��^�0�,���S�˨S�w,F����z
ͥ.����������m6�W=zx^�:#R��\�}Ք�h+��=�y$�I���1���4��\�ɇKQC�{F�8�M+��6���՘��U����}����;��5���;;㚚z����s������k�����HvȺT�\JLG/�l�ɳ[۟=3nY֎�4��\���0��Gw�[/{��9UQׇ�7�l���ˤ��#��7���ԧ�iKsz�l�m_ro�\76�ӣ_\�u�T��<�W�p���Y+e�t�g��>�:{o�Oג�3*��n^���^#�Ἴ�W|�8��*c���s�կ��?f���O|lO�6s�	Wn.���I]���#5��n�����5���:�{+��Z���a��Y��o��;�n��śt�p<�&��h�ÇY{��먳!h߽(z��X���홛�ƃ�)	��)�|�y��zy��*�x�A�̿Vd�ԥw����ޚS�=O'Ǧ�gk�Y6D��yL9Qxx�^�1<��{��ڍ*?��m�h�,I��r��4v�k�˂�3�X�4����6�!a0��h���vȭgk���ʖ-Qx���t�aC�ͨc�'���m<��bkW]���i��W�Q5غ�	&%og�����ﾠ b�k���_���-b��x�Ÿ���"}��W�3��7Lz�z�o[�p(nޘ�^ȗj���Y�Ztjb�f�,j��H�1T��;�w��W8<vJ�s�miYSP��y����+���P�*�t4(�v/[�5�G�k{F�^��=m[��\��ќ;4��|i0����V*Vqm.�ͺMo��#���1&�\A��̗3�<���;_�3�|�B��B*��wOu�X%���!W���;��L�"|���U{\��ٗ�4U�K���4 1���[�͝rM͂PS�U�';���u7�Y̹�ɪ��4Ttli���_xs��ʐ�,�s6Nw9�;��=�4�,Eh�����5S�$"2��G��y���@m�i�`Oe�����׋���W,�E�7UL�w����Z��M�fψ~��]`�&����S�����}�Iҭ��R9P��s�97>vOvS#syU�ա�*n/u	�1fs����L����eG·�N@���l�c��0+������u�~��aw��%�M��z�/�1���H��ۺ�Z���Y6����It8V����c��O,�������fw3��j�3[���.-rV�5D|�>�xל�J�{]������n���K���b{��krj�Q;'�����M6}]����)箕k��/m��/�g�������8�eq3��맾��5X�4\����پ\�W}%��y�v�}К`�s�r�͌�s��Uu�Ub�m��ür��u����y�!i�y-��1ϲ�\���{X|Ӻ�39��tҤǦ�^Wر��q߯{֝ڤɦKǞ������o/>OlMW�I�{:����R���I^v�����oV,�i���S^q�9�z��x_{[\��8����mZƌ�|i��:��{
2׽���:ػ���Ah���\+��QK��;,93lU�%]X��)D/r�(��ٞ���>ZN�����[6�ޓ�q�1��Y�[��j���U�:l����ߣ�[�|IdK����r�k����ohm:�kr�]HP5��>����fѸ���AU�
���O'��{�T黗�	�&LK�aG�5c��9so��W`�]ƏWT�yu��z�e+kƽL=ǯR̷��g�������]@��MWV��#�p�^�k�֫b���zd̂aM�aY��g<�}�}ל�5��Ǻ坧Gh�l�K�9�T�r��Wבdlw��[����A8�ꙮ�;�j���Gs�D{x�@�Þd�.�W����T�~e~����݌���z��u)%�N�_4G��&{;�=BZ0]��~�uo���l�[~�89V�S�"Qʿ���i7�g�z���)�0)�Jo�l\�磭|>�%(��)��^>�,�2������Q��3>�O��zצ�B��d�S݄������'3U�ۙg����pn!��hu����y�_?vQ����Fv�?c�f_N�7�\�9��Ao�r)�8
w���d�yom�}�<�{ĞO�ɉd����wA�#)�zn3�Y0u��~�P}{u��H�øugV��F��u�\�m8f�\5/c�O	�"��W:"�;�C�0H�e�B��K�'Q�=[�ʓNo(x�_�[WNlGu���H�tH^�ݶ!�8�}�U�]Q���7M�7����:�yYv7Tf�ד����G�^�L�=Jt�e��C,�U�
���@�����_>�,z��PPFY�	�#�����mzO�0j�_�l��Z���r�$բ�r$�G�I�ё�Z9��E��ʦ�]*a׌��s�۴[�y� ����SBH�Z9j��
����9:o*]�S�/��zr���H�Vܫtn�����uc�yz�u��Ǵ/	�`�I�-�Ӱ�h5�Z;��V�s�U܊$�(c���
�rXJ����QgT�E��l�8DN\;�pJs4	1�ݭ"�{�e����<)2S���'mG����At]!�ɱ�����\�Sv��w�x�N�@+��M�� ���.k�!ŕ{ћ��)ؼ���M6{����I�r5���k,���mM��4�w=�ռ���"��� �u�!�v�N2���ih;vrq���@�ʳh� �Q�Kl�����uq�����~�iw�X�
(TNf�I�̥��٪j��;�ʔ��J��O2v�����gY�R��&������6Eb��5�b���w���6�dim'��٨�K{fKX�uq��M�g��R1�k�՚�#��ݻ׎TFB��ո�{�«��9u�zy�};F�,<w�R���Y}�ayfps��$�u����!M]�A�3�a�������dU��:B�`۹a��t��C��<D�U�K�޴����������n��|�P��y3�u|��T��k-ݬ{�����y��)C&ܽ54���;j����g�� �����;�f�G+�,7Ǔ/�
�.%Y�(F3xg�B��;��5k��^T���u�[v1���`�>��G�Jh��Zݔ^Kgp�75�O8q���99���	��/Gu�VfN�k�D%֌���h����QL�v^oWM�	Φ��V*��0�(8��nl�������X(������I�`��sg���m����;[�ܩ[-U���4�в��M�C�і�w�{�u��)q�7k�&���(l�hwc`j���"��	ڻ����]E�nl��T���μs2��#���]k}R�m���Ƽ��^w����� �r=�{B:gG�n"3��ط�xE��9Z�Wv��K{���pM�����K8>pQ��-e�{�����IK�um?�m=W��^��c���* �X��1޶F�{+"�m�;�n�t�Ո*��wP�ݴ:����7+���r��컾3/��a$B�2ks�S2�����Z����g~�(C��}�5��6�A�8���y�C��u�[Ú��N�L����t)җOv�[z��O��Y�(���� ~$EDX�)UE+���QQE�Z%E��0r�"���J"�e-b��ʱ�Y.[@�D����*¡*�[�F�*�Q(�E�XҕR()�ʑb�`�E�Kl�����V��[D�[j�ʩ*,P���(��V��
J֪9K��R�J�X5��R(,��VTXT*B�IZ���V��؉�*��`�AU*T�ԬQ�%TQH
EmRQ��� (�D-B�6�Yd��YX,�-̕��q��X-@Z���)mQ���U�b�*�#-XQ
��r�,�V��PPTV�kQT*,-�R�+��lD����*���mZ4R�T�*�TTZ�B�EQ�
� EEkV�&e*��3(��㇛��[noz3y���������������1Zx�tˡ�Z��9k����=Ք�����J�+���v��|>���GI�U�����o�b����ױ��ٚm��݈��l�{ϰ�י�Kۆ�M��cגgH�+�q�&I�y�"R_s�ש{u��L�Or�����񦽍�b�F:��Ƨ��S٨;�<Ƕy�u�+nMo�ǆ���i��3� ���\+���jb��m>��~w��|��A�nX��;'��OP�:0Ǟ�h{�A�.���Ȍ�@�}�����y�	��d���ǆd�ӣ���c�n�#K�ɜ<����WY� �U!��S�spl�]hw:�zY��:#r"<����8����xl��w�2�v`�9�\�#�?k���}����]���SB�񆇣�:f��x��m�,����[�LRhTu^�+�;	��{�^�۠��t�B����]�b�gg�����ϳZ9~�����3�q�:�VP#���;����l�t���������nZxՑ36�q��y�����4�v��a�7[)nk��6z�	^���_V����vĽjc�j�*�0�͢�'N�y�k3
��hͬ�2+��c� ��H�Ӽ��z���bH�zL؄����ƀ��HS��Y���]�Y�ys�5�Oۼ;>���8:Òm�.������I� �$jz�$v��nu�;�{�������+~q0�
���S]f��H��-ՈM�y��7���]���S@��,oM(>���pr����6k�m�{ﲖx���#���.Ͷ�����w����yA�����?iY�U=�-U��%�擇�/���E��N��LX��깽��=F1\�s�0��}�Y>n2��&�+�Y�3��yᯔ����R�Uϳ��fv�{(��<��}="����;q[�<��"���,�����Ke�&|��K{:��^�z�u:X~�&�Ϋ�h�����:у�u�\Ujttn�V������	]'Lon=3n[�c�)z�z.�Vr�rQ���jTwuo]&P���a�jaV��"7^b4oiV�f�:V�� �[�r����m�ˤ�pv� �]˰HQf8x�6jWn���6���}�ٻ|�޾��^�mr���AZ9�N��7�`�6�V�L��p�y*oR����꯾��MX�S��V�|a�@���lU�yu6W��I�6	_)�*NkV��x���n��G8����tv�3�p�|�]r��2l��~;�^�3��w�Ybs���:��U$jQ�(���|��J�m�o�~���P���KJ�����V_dr;�R-�
r_4=�>�^|'K�|M�J�ծQ@u��-�7`����,�Ŷ�E�Rj� �;%}��~z�ExG��I�]�;4����1	.;2��}cC�W��T����G��3���A���S�wu-���~��lE��-�p?-$x;5�V�+��/}��i/i�9�n_IY��}ީ�	��b�V�E=+5�;�uSE�{Nv;ѷ{�8v�T�S���Gs�į�s���X��=����v�MK�=_<l�1龼�1c_e������t�}�t�u���v���Y�;/Ќ��vއ|��5E.=�u��tr:XVc�TyY�%�r���7��t�.���$�m�N�����Z�������q�c�]���̧���N��p)�&�w�|�]�+�67V~��ˠ��.�����}��E��S�z�^V:c���8���P2n���Y�0�^����Uϡ'p/[��N�&b̡�b�]�������&�ۋ.�vc�Tk��#�Y��5f��ZG���=+W�xh(5���X�~�7�;-ɛ��y�9_��}=�^�o[`�Xh��r�k�����{���=d{E)��6�o����9;��˂q�M6���2`�S^��[����_1%�J�UZ�u�<�o4]������ӏr�Gh,Q�	��[֯J�U�5	Kn{s����Og<�8�S�ua��W#R��7�y͠Wa�:�p�k����*���R�9�=����s�ꤊ�NI����K����B͜�t�~�y<`�w/�$���>�ĩ���Y�\Y9�H��]=gd��>*��;��\�%i�J>���l\ގ�|�`�q����5�0^4���R�æ�}T�6��G{WH��nGF������=OO]
�Ǌ��vΡ:�gv�f�h�V�]y��̯w3��Ag*;����\:��C��+�j��R�ȷ��UgB�g
g��XƳ��۫i;rv�_v�`d1{�g���\1��/�Z�MR�tJ�z�{+���I�[��[�c���3�%v��w��g�6:�u�u��D��Z���S�Ql���=s���5˻-��`�s� �xWA������ʹ�_�"������_^��'��-���ҟA�y_9�M���%�l�g��fj�6�����@��J
�9�o&=�t��.gn��7���6�i��^}\t����C�k�|�SY��qQ]��3zl�A�����k��}\�ը�u�4ײ"��c´Ff�oS��5�Os�=�3�E>��O�ہ�;qc��e}�i�eE�ƅ��˄�S�K	R��Dz/=�I��0d�I�ߣ�ϧ��i飷���2vis���gx��c���ع�zd��"�g|�����#���,yP�곶�w��)^����)Ť겎���B�kNU�!�fƊ�ҵ1X_N��nt�C$#7IWQ=[�������-�%\Z�A+�9y�{�J��K��)o;��fG�Jhi���:����"	��&��}gc�f��q��XįMك�k��<��������"a�%�z�����͡;�~�{�?	_)�*���r���,;�Bh��;�6w�����9�m6�L���vgӣs��J~��~����׊|ib9vANw�6�ܴr�tG���s��J����5�J�fVOA=g�4Rk��L;���{@6��aH��Mƾ�N�)�؝���29H]�+��n���d����{9�����'Y�c�e!Oj��ھ~u�k[���{��N/�Y�K���Áؒd�*��2���x/{עё�&���]�Y�{>�Y�GĹ�d��aº����t���҆a3�{&�w�qAc�W����V�z;�K�ziO��|�pNc�x�u�X�գ�9��v�@�նo�^4����V�������=H糔�a�-f닶~�Gg�ʥ��=Ɓ[|���ly�@��G�km*���Q��?�~�D��,�*��=�+�ݬ7�L�_�Y(�<�	ۙ��y�N�~zѠ��F�֫������r��۬�����A���{�E&�o�*x�=u�ϐ;]{���/7&�Ɇ��C9������}��N�l��^�"f���諭���zMl�~X�n����$���+�y��M{b_y�#M��y(ɗ��浌�&G
�8'/5��5�ڷ����g�f���ꌯ�ѻ��_�_s�\�L�p�;g��u:X~�&��|��;r�(+�ynY��W�\����,/Ǡ8��9s�C��!���g�2u	a�.~{�e�*b
�]��SV�\@ڠ�Jkk��U��K�Z��H��5f�&!s�!]����$c8�M���ՙ�i��0��
��_�&���2�K�3�e�{<���=���u7� %yt�׮�Ű����a���_�#�H�x�|�5�(P�b��L���Y~R���쾿IZ�<�JCH\��⤥�JW%�aR�]+Ěq}�^g�J���B��z9K�<6Ԟf�>ir���y)^�1<+=�T�hϔP�%��|&Dz�%q���'.���A��(S!ҿ��k�����>��gˋ*+�%��Ć�W��[�N��A�=�
E�=4)��(�o���͉�yO�:�y!v�sYQ��t6�bwBJL�׊�%�V�u8�٧���B���\��Y��%X3{h�/J^�|\�]o�t�M�ݤᵽ*e���㼊�����{��}hs�K��4�j��;���c쭋x+e,+���˩�]}��}U�}_o�x�������D��GCk�E'K-��q>�1Y�ʤ�.(i˶nY�yz������r����H@���/��;b0�g�G��Kʥʮu�R�p�8�wKE+�RiX}�Y��)�r>��MN�5&S$Ƒ�Z�'zאx8W�L,{J��[I=���"�^���#�g�zA�)����%:�4_�Z"b�%W��j�_�b߇ZW�JK�����Zןz���*�~}s��9����6�Ȱ��9��m,��v�CN��䙱�"�8��~��{<�f	Eof��W��8<��1U׵�A�V�qe9�=�����~C����n�Iϻ%߈����R倹�[���Dx�c�e����=�^�+�"o�f��=ެ��!��u�Ft�����l��VGL��H��MH�K$qQCS)���M�ś��v���3Z�K�eկi�p*�t+Q抬��z"<8�z�L��(�-Z���x����%��!�Q�'[��f�X&R=b]�Ĳ�>K��$V�įŔ+�.�����~~��v.J�nW]/Z��U�#��Z����i�t����DXV/g%zR^k{".Iխ�G)�s+ܱCO�e3ֹ��ڱ@��qWP3PX+�u����5f�v�I���ˈ�7�;��C�I���.ܺ-��N�[ﾯ�諸>�5�x�ɸ�?T�¯�!��^�]eo8k,�\s�VxIl�G��4Mt�;���'{�����z��̝gL!��:�И����^i��B�瞵�ʩc�;	�g˲�ԑ��^/u��� gٴ�WU~��R����SJ~υKZ^�fw���2�=���2hE2��w=�s��f�I����Z���S~�X�y��O_�?3�ҕB��S�ԑ��ޏ۹��6���l9P��(Gt��-�x���o�}�����#֥,��޾ѽӮբ��O��\���&�!��M�T�*��f�Rx'ϔ��r�D�E��2��^/m)�ݜFf��J�܀ѿ���n
z�J'��0��7���9�<�d�Mw8%rcd��ݶ��ν��
�=:{i�zz���ّ,�ŝY#�oj
���Uxg#�|���G@�b3Ԕ�4����nd3s���_W��ߞ�iz/5���ǧ���E�!Lm�#U�e�\lo���G�.V�| ���v�{�[����6�F<��G�#Toz����K�P�%�Y���ƀ�z;kk�e��G�7�s	�nV�#�]uـ�Z3�	���Y�C|�A�%��;z�We�$�E��d�n@�m�c"E�.j���:1�m��<���ݑfI�{��'��c�e�άA�o{Y��}_UW��p�uq��]�2Ml~!��-T֥q`��]�G�]�j�T,�N%LVJT�i�:\�Һql��M�xeD����<�gr�ц�5q#��������Bf5W]�ҧ��ƪ{�G�>֔�j�,�Jw���!��q�;;L�կ+�juMzz����o������z�����48�^%��$�(��l�a��MP��C�Bn	���Eq�k����	5�O�{��X�*�I��TEp��X�Ʀ��b���K^���23�
^�.%���Y�M6�_{�,�.,���3�a��LB}�[��ׇ��O�{��.)ԁ��,s�3{=�^f?Z�#+�I>ix=�D��u2�L��iI�ۄk^�����5)+���g�������6�}^^&]�Q{�:�� �f��U��$�,딡�V������}�ۓ��m�BOj�Ү�y񔧸��Э�;��F�����K�8��tI1[�����t3F�y���#�g��7%dA����paƪ�1���)�u��;{��:{2�Hue��Wu����L�|����}�N�G3��dno\�n�����̧�1�����	έ�v��K�.q���/����a��V��N\
���۫�jmʱCM��kwyQ�p�)P�X��{u�� YJ�M�{f@���f�W ���
S\� ��F����<	v���q`�FT�m7A����p"�E]Ȏ<`]u7��<��"�7>�8���۝�}צ��kYB�l�g"3��P�����KpP�U��(OP��m�J��Hp�����ѽ����G$��싛�)=�&�5�2%!���(ν�X����'4�ٷ�)i�����։N�"�GV�R<ðM�ygxC͂�q����s��*ͤ���V��k��u��݌�h����=L;��������Lx���)���[�:6��i���\ʅh��&^�LE1ݕ�\�<��$�W����i+j=��*m^��GP��[Pe�Ė���r��b�cS�Ѕ���HWg�c�ui��"zڔ7�p/�&��� ��]��h�����3R��dVkW7��d��1���, ��9��`:<�X�|�{b��ʷr�v1���'�v<�9���ܠ��˛�8�F�Ewv)}]t����g]k	��[wnb���2Nt�{P��A�&օ�l����u۶&�t��)�Vg<0ܰ�V�VyLn���������2��C4Χ{��_CwS~��t�Ԡo��s�^���	7�zaY���a�[Zq"f��������l:�o�� of�@�}�ʛE���`v��P�"��)<�Źz�wY��v��V{�����c��i���ѣ�j·		c�ɏ�5^u*�� �@�W��"l�ہ���M�i���$9[�;���O��{�7�2�(���BQ~0���o�y�F�Z����;��E;�3���yfH;n�K»�-�E�d�E�g��9�N��]��.
m`y-Ip*ζ�v����˩5�\�ض�e6��
���O������>��/o��v��!�+�N�{�����8 ޵�Z��KR�u:�{�oS����Y5[vM-Q�T[��(���f�N:��ڋ����`q�&e�Gd�,��l��0dTe���h��/�,P֊�I�l����&#�#�~"^�T8��_>�}������������"[�������p�ű��c����2Α	��[8��ՍRzɾ��x7�i�����;׶�=է७�c�ktK�H`:J�,��u�P�K=	�s��(wz�}>|��\It�Z�������1�v;^��h�tz�%sӑ��MDo҈�T��lwpp�mv�-��5λ*���~>��r��M��a��V">m%3�6�=�cϕoXל���Y�Om%I_+�����Y�ǀ��I�p��6S�j۠zu��#�c3I�Ssw|��}�y���b�`���YPl�XVVfa�V��V�D�2����Y*���Q�b5������!D��j(�2 ����+e�(���-��m+RF�U�[h�"��Ńmk[[
�1b�q11X(�H�iUE��уl��+d�dQ-!�`�q
�bմ-�-eDVC��"�YX����Y""�fZE���$TF*bm�q�2�+	Z�,2�(V�++-H�hQQm(���D��Cd�E�)����*���VLJ��
P��b

�c%�(�%���H��̸�X�²�
5�B�1RVQ*"֭j*���TX�Pl�+A�"5��"�*[V��X���*�$U��*����E�0FVU��JZ���ZՊ�X��т���++YeT�E%DF"�T���˽�o>��Bq��2q�Z�ˇ*���A������;��#�aK_ts�]��D�#.��L�{�q��ﾪ�����tK�CG�u���u�E�_I}�9��ΨE[���-jϜ�t�^�>��'ry�����{Լ�:"������u.�,vUτ���y�B�MC���ɮ�r+�mb<�_F���%9�巵ıFj!~Tz�Q+O�^ś���e+��3*Ia���r��|����d�>�����o��z��Yo���xd^u�ƴZ=B��w�Y"(��my�o�	ְ�T(�{�y"���g�ۢ��E��]=��K���.$�Q�odޙ����8�Y{���b���Փ]�55�P/�P�0�k���f[�id�#c}岫LKB�!�ޤ�X�⶧\8�)��u�f�!�$h�Q
0n��y���=+��uZWz꫌��]�I����gޔb�'P���4��7@�8�K��C�ՂRg����C%�[L�����i�H��'m����L��	R�U�:̜��x�8���l��kN4�K(v�Di'�`�	kS
��ڣ�ܹ���;<�Z�i-\�{S��GN��ըK�h[�rm�E�҆_G!�8wS|���dh�S����ftP�wy�MR�m��"�t�ĝO>��6�Z��L"o_p�=L��u_S<|(���Sx�"�\­�V�>�b�`^mn�1u���@ӕ�V�g�W-�����	�-���}�Df>\}���#��;³е��3藁�� $��`(t�cp,���}��cp-xW�f}�w�֡���B�g"��R�\%�aBY�k�x����[��mSM����(sW������zG�ĥ{��Ao��^��E�X�n�Pћ��f)�na^0)^�yUqJ�gho��/�>��`���	=0u�7X'��7V=��D�G�˨����=-m$=�%�,� '|B�d�ͪ�l񳶞�Y��t��Ↄ�9`U�_Y�/9M�v�x�`0n�#BJ8_F�V�6xO������K�s�"�k�����g��LWA$�y�bǨ�Y4��K�L��:��>ˤ%�ؽ��
���,{sב	�&&��SDy\�x����[Y~c>�0��|�4^ƼD�u��
�v���[���+�>��bN�`��wA:{��y+������_���c�dR֜{-��v��߅:kW�f�NRΊ�kU���v���1p KԷ��b��=�"�\)�����>�\7p�qC��G�.�48��s��tn���_���dV�8����UY��39<�VѾQ����I@i��D�HH��b���\�X�#a��o�j״�+��n'$
�����Gw�,n:���U��]���픇<}�| ��ٌ��;ԍ�<�����[����MiV��5"8�ф�4���^�;���x4_�H�]�V���|�%(ϋ�X)q#l��E`�=Am',=5"W�O)�Z��^�d��홽d���Q�q��rs*����.�j<�EVt���(=}���M�7��c�K������&d��Q�'[���m`�H�˴x�L��"vЃe編&���s�z-�Tg���Rկ��+ə�};���q�N�d�Ϳ�Z<TF��d�ǣ<��ƊKA�ݐr��ZY���u �|����U�kZjus�Z�J�eT�ֳ��@�QmrW�ϒ�v�3�J$�1���{��~���g;�ꖴ�>�g��y,����mz�u��0vS�0!5夨s�ZI�]��=>��ر�z,A&���z�������?Fyޮg�<��(���B���{µ����N��U��Vj�D�J����b�{�S�ʂk^>R��ܤ�JpS��	����A�S���{vx���x*�i��=4h%.�n�O������c��H���8�u9�7Treʎ�_$Qn��Z{����F�/W���Nu�ۋ:^5��`� ?��(֞��ô\�Iw<�c�*��凝s
�C;����b� J�};(�ua�Q���?�UUU�,s�w��y����x�vK�綰O�����`ۂ��҉��4a���׶;J�י~�{~S��L�����Ѡg��ѝ]�c�cR}
~��g)#��BVaX�3�����\�Z�z�4��(.J+E�qpr�O=����_t���߽F����M��<���[�x2�&"�U�[�zP�-��:��q3gM?X���u�cιtк�҉��\�􏼑Q�	�-�#�/vR�jԮ,��,�*��z*
�\5]����7Rm���A�p�\�1�;;�si�WH��U����U��%ff�>BF3=�3�=�=��]bP=4�Y^,����P���ί��
�N��ϔdh��{��f���s�I4Rv^B�ez�keC�4��(��f�ST9��C�s阎��m�*Y��\~�!��>R�"��-��U3,u�E*���!?L�l�<�s�����k���g��ܣ�WI�A"F� ��5����.{��7��vf<.V)�Z�,��,�V|��\ �a�#�kVY��k,Zq�||m{A�_�d/�Z(b�	%D�΢F,e��x���|����Mv�>�/���ڽS^���{CbV#P��k��\]�O��o k��&��2�ͨfoZO��/�Ƕ�:*nN2��ܧ���}�i�:�L޿f�����|1�a�C������D���h&f����ڄy��^R��`�=��ݸnM�m��KIVt��w�Ԩ�(߃!��$�E׿�yI^�8U�+%�63���P��� |�G�+2�*��Э���-
F�u{E�P~�á}EDU�͓��\����8�Ř;�l	+"�v���PêZF|���j��1bC���y���b�t�pt$��/szR'�|T�s��Ck2�V�H��yJ����#z2�j�C����<�����wz�&@[qN�MU����سއ�:�Aa��`�Y{�5�>����>U.|��Ksǃ�O��}��e��>�^���ڭ�/������"�p����z��Z�{�`L��w������1e�/��J�y��^����n>������B/�Uvu�-�ȇ	�k2x�od.����<��0۞�vM��ZE|�J�k��m��QzΎ�/T�P�1yl��Ն��
���ރ����ב�t;�)=���ڼ�fFMv�}y��k��o�G5څ�����)*�0�6���皹�9ڴ��� ����:1[�b��de�o��4�;�u麴AL�Xv�)��9�nl;����UU|x�_��#s*�����uL�ypP��
�M5���+w;!�sPֆy�^��l[�8��d�w��T�+=�a��.�=�U�O]Uq�򈖭�IOk�C�(�/��Bm����l7�+{�Z^���]G�7����f��IP¨�'�?�/�"�t��
s~�"{qװ�m���8�X�����M]�d2��ʜ���|��;U��\��KZ��
��ڣ彷NtiZv_�+ވwY�T#��{.�6Kf����˜�
�Bה��%�FU˯U��2o����s �&�;ۋ�+��/P�n�i�?{����.&n*&�N�#�:S�slh����I�q�(=W���>ir�G,s�J���2��[�/�0<r��n�U�^����V= D/��Z\R���i�_�Yk3�ʊ�����(�yuhm�b{����$Iy��|��ez��I[�GY��E&��z`�9T�~��`Yk3/hS�2o�T�f�}��ȉDq?�˰�kɜ����J�л�̦y$"�ڂ-�{�5��EsX������_���9����R�޳}�B�7�&6��-����x%q������>V�!�2��u8�@B�J�5:�P�|]t0��՝�e�Lܜy^V��7k��OhA���Q���c���}Y��Y�� |2���Eˏg�ux���d��Џį�������mx�Z�2�1�Y��͟b��j>w}9��:^�3���k/�`t0��@h��;����ߺ���o0����Ӯ�fw#(�_>���^�R�
��[G�5�U�!����5����~�̦we:fͮ8��5�m���oMi�g%�2R��U�(u+��]�s��@�����3��q=N����4��O5q��j��4�5��P�k��8�ZV�k�Ԉ��Fo�:f.l[�g���2����9�RޯD$[���F|]
�K��g�"�z5���}y�1�\�=9.z���e��bw��{\v3ZԵWKP妄6I�V��v�~<�#彋9\��d���My(��3}�	��ƵG�o��Fi�\������@E�N_3��7�P:{��̺��1��Y3���XC��r�ޱFú��y"f�5�o���.�6O>�mv8w�7ir6
��q���l;y5D��`����s�Z�L����9�w��X�=�*6O8�9;�`�n�to��.�z�ڽA,Vُ�JP���#t7����m���o!n*�n^�'خ�A�����U����Қ-M��h��º���bRJ�g1��ֱK5s��u�-`Z]�>�{	0�u�>���/���N����>�
�<���I3�
Aoy`:��}�_���,��n^�Ѝ[���f_�86��;��nԿl	u-d��夫�t�I5�����ary��������X��Z�N{o��5kOai3�%^�\�#~�(D�{�>�k���:����}.��:�n޾�8�E�O�e��:�4K�w��p|�eu�A���xs�ro6٫^/t/{�����$��껲]�`�܀�&�=K���Y�ο_����Po����+}G.,x:���O�E��؆|�XԱ�*�{2%|���g�t���gWF��ޫT�ık>�C�חL�ͻ�.����] C=���gQ�©�/b�{�@�����6���c�	�3��O���sσ��#��O�}��+��|���7���"=���Pɲgrыun�QiԪ$|EhL�+���z��������7�~a�`��K>ܶc�vg|����uhͦw+-m�WR�B �j���Wo�oaYL�:�=��m�H�}�#p�P�b�z��!v9é�9"��&LN��ݖ�2�x�.L�z��-��Y�ӖQ(�"�m���e���֮k��7�Bs�HN������v�N��d�[b���c�Ѱ����h�Y݊ ?��P�ĩ{}���UU}�IdN{�9W���C���_i�_����M)އD3}��a֩��Z��i�ւ6g'dr���R�`�C�L!ǚi0��S}��&3T=��C zhMƕ�}oз�*����;"@��#���r���;.ȫ��X�Ʀ����s�j�ȅ�cyY<�����d~��������4�oW�����f!|�̕U�*U{�<<l�/wX~Ϻ/�u`��xV\R{�^d��������������3;�Ҝ�"$AWI����q�i
�"��w�7)=2]�.b~�� �erY�.���n,�sU���ĸ����lM��	�B9�b*kK,ב�.�D�(�'V����j��'��U7�]�*Rz��	�Go�$Q���t���%dA�v�p(|0�phL!u�8�YN����b]�F��B���ix��s{�|n�{ґ/ڼ �`����Yj�6�m���0���Ѿ�>�������U.�,vτ��=% �ս�3޼`H�h�+;mb� b�B�^�&�����;x��M���
ө~qsN��b��e{rL��<�#�裗q޼3�N�<��\��.�ݗ��V���4��jU��/_bI�4!��Qq�䢫��Jfm��\.݆l�^E��,�6��>��V?���}�m���b�>nƃ"Ƽ�ijnmß?R��<�G���U�vk�#���L~��)�����ahN�J{P������z򹵢��~�P&�=��$���-:��w���G�����l,��ዖ�B�����g�	�8�^�o�i�������|��8=G�b�-E-	0x�~�-L�:��t?B���֡J�#�W�u<��������{�d5e���(I낅^��\���������:�y�[,���y龔�����C���Cs�~�*���U������ �#�|����><z���1Z��u���h<.����j�v����P�j�R�//�a�U"Gx��=:�`�ǅw��Ժr�~S�K��w��	C�ßN5�QC|�N����l_R~ms���8��{�V�te��]��Z��%���]<�}s��Y�Z��DB��
Cujǘ�����r-M�ɧ��(P�Ug�+�M�J�3��B���S���f�KD��+p_4�WM[n,6wۘ8�Kh(L��YS���']g����s�q��U���8~��p�˕��tKoH@�{-���,l�/�TeJ��V�h%�P���;�c�'¢���Y�y��4i1-.طO�\���d�a�rhX+8�*:�w���pm v-�c�+d�롼���N�]�B#��)�%���l�)lF0 �z��C�����k*K+��Sa�q_t�m�V~mLB�#)�t�^�!9j]G��+��S��q:��X�;��&�ń�*n[��d���VSu)��b�e��4�bI.�yM ��*�uu�E�C�o)�m�6��$�!;4�c�R¤iB��*-��=щ3Ac:�)Y�xs��R�S��2�_b�w;�j�^��/_��{�W��}2F���fI��
��G%�+��Z�r��Uu��[G.뵒�1`en�R4�1��е	@�Sy�ts4&��2�cl��;ƮWu�eNu�/�����X��u�Q�ұ���;�3\�V��eIJƷ�� RL��1��طx����	j;r��F�A�
��Y�7r��-�^;J����;���z�����h�eۗ�����ܧU"����O�U��#�Ծ��ɷA�r80Q�ĕf�K�ۈ�R4,e^�hަ�lֲ��d��#���]�߆sc7�I�������\}�:�ur�KH��p�_jUz��r�+��$��𮜟��bT��YՂ�oÌ�Q�Q��xP��`:��KO�������N��n��7zto�{i��K��Ʊ4k�ߖgcb*��s6�ѷ���ϰmc#<��Ŵs��v�T��W$�#�x�����!���C��n�@FE�3;��;W�{j��^0�:��¹�Y��<�o1�Y�z���H���ɦ��m.�ԗE׽v�ň�He]Ǭm�d����/8V�zP����U�f��F=�!W���e��x�=s+(�҈:�o����r�>Ө4�>���e^�,�*���P&����U��A�\N��9�T���;L�
E=y̧ٻ�>�H�����G��cv*ŏ7�(P[�Ē����HعR�Y"��2EDVu:ysX<7SM��Je6�����Z����D7�gt�o�RT�p^E/7���&�:�470,s��$��V�W1@z��e�
$�*�A^�j���(�2+�{��溉�N��u)Q:W��I2���u�;�u�K W�*۷\�eB�cn���!K�X�VE�m�gV�%��*�J�0�ޮjʾo��]J��;��;�����:�u�=-e���Nu-Y,e�������������GF����s/f��Vs�Nyʵ�,,��*R[J`������5��F��Viz9��t��L�����@r+;���};c<�&��^-M,`�d���:��7w���v�v�O�gw�Ă!$���
AaRKhUE*��E���E�QUT*����`��UFZP����cX��(��b�J** ��UF"1H�\e��ƕ*Ƶ�e�(��EH(�X"EQ�#+QEX����m��؋��fE���J�db��,UQF�J�(�,�ʬ5�`*�TX�Ѭ�*U�b���h�TDUґdX"(��(
Fҭ�Q��UQb���j�T���`"���DA`*0F.Z�++"Ȣ1b��Er�jPq�(�"�Tb�TFDB(�
�VW,��Z"�Ʋ�i)UFڲ���?P(�}�Ǻ�Z�v{��`����m�[o�Kz�^���o��3Sg�aO3:�4[+i�-��쫻G���������J{����&�$�|D;� �܆�k�q����{��Ao��^˔���N������?{��=r��"�<I?a0V�Uy���ȿ]���	.Xz꧘�~�S���N��r�Q�U'�B��W����W��GY�/-��K�,_�]n��bɹӸդih���Üޫ�����(i0o�(������N���<^ʔ/,A���0Z���26^�5�x�n�"�qwJEp}0�hF�qq%��Z�^_E�
�+�m]l8��+�l��U�1[���	��ּۡ�/��P!�{���=����j�x+хe�uOum�"��ވ��{��S�ZJ!gn`g����LxnX�P��추�S;�]�x��/�7	[�8NB��;�	">=>J�ȗ%�/9�P�v-�,8�S���_{/l�F�.Ж�^��K�Z`�v�jћC��!���ե�E�S�>V�5�Y�<m����~�g?���n_�V$2�y��'����*�g�Ь��m�D�z�9�<��{&z���b�~�/����+�:�.9���p����g)S<�.y��t���Ak�yk
듳i��I����D2]m>����>�A�'0��t�J�S����O:Gf:�X`|���G���A���^\�|q����/����s\X�c���4�~�z_��v�ե��jZ�B�Z��C�U��%y�B�mT4��?O��3��р�����n�&<�5��N��њm`�H��v���s�s��|;16OL�m��q$y�٘+:�3�|��؉ޱFú���S,��O�0�syaU�$��y�Y�h{�Dl�� ���2�xu��\�`�[<�Ө �;���p�b�,�ۇ�Oj�u��d9��yH�s�I���_/�{U�Ρ�j]y��V�?.�O֍��Γ}��i�PIS��	�1d���89�-+��%/���{<��d{(��ky�����8{�V�xI��6��B.`�/疒��N���x�+���"g��}�U鱰s+ǭ[C�i���L��^*�%����}���&��Y�vZ��*�+rk����PR��
�� �6�{Cu�]�K��{p�_<�_8)�](�qA8����K�Ժ�=�9�^���k��:�#�aˋ��_���������Re����p6��<O��{ ה���Qn�`�r���V����G,�E���_%^��h����yG�.��)�ɻ����WUɃzB�|rj,�-�m������b���	��c*�Y���O���tBvl���GT�Y�vj賯��R��m������4Z�̽��7E�D�:��e\\T����S[��0c����q➼���u`C n[�����߽k���%a�k��m��O>��������]���z�Y�g�B=��/�H����υ͒�������<��J��)i.#�fmw5�.�X�o�F.}�+^Jj���w����o�;<-ȧuh��v�׌(1�]}��Q�s�9�Gǯ�i�z�B���+AG���i�_���Jw���!�읊ٮ[�&�v�,�[����K�$]�R�l��3�UG�R��_����_��(�zY0��MP����ʝ��y�,�Q�`�F<X��{0qvW�4x�Ȳ��?�b�źV��>�y�<q�}6�m��j��l�ט������p��_���ѭ�E�+��̱��T!�v����z��T���^S<x�.s��-���!֙$?;��J.�]�B��,4��%bۺ���^���\��B6{Ug���6r���2]�*�@���!}�5h{4�?c=���0
�A��
0����7Uo;Y��t��s�����@{�*�LN�M]�C�$5y3X�����^����4E`k��'��)�f�WVE�ߒ��m�	��f�gMmZ���]i9�Ƙ����H!v���w��ta'�M�iY�`�/��{k� k|r��[�����Ušm:�3Q��	�J��R.0�^G��p��D�y�KױUqo/�w�1��BiaH�ڧo\�r-[�0#bJ���ę�C��}j���HKAk]m��FƉ�
���G�����1sj��ܡ��zX�y*O�P��#��z3\�{z�{�bDN�-(]���@T��|��:�w�c���g�����,VU��2M�T��^��!�9^kR���-��R�9�B�ȶHG<'�9�)���.0gm�G�C�'��A�BHNb�>σ�o����x�Hp���[~���P�ά�:��(}TY��mf�`���P����~62P�����f�g�)��
��E*Gމ�i��p
�R�C<���Z*�������e�{<��s��*�攩o�Dӛ�*���:�B��4�XZ�.�k�
h��[�������ke�a5B.���2�����=�v8�b��e����K�Z=)���� �#�3��my�0��ҷ$�]�9Y�s���L㣱n�S�jV*�-T��'S{�EK��?V4GH��x	�UN��(�k���@�h&��&��-+Z��TG���Õ�Jm��+�-q��Ǩ�j@�:�]E��w�.����M�x로f0�p��_T����yΣ~����L��B��]��*��O��ꅢ��/�a�^��{<�~�=�[��$d���/�s���C�Âq�2�Q|ԸKb��M�ݽ.���qu�����g�V�Fg�%�.j��T欧�Z�^4�oR~�v�oО��k��G��k]�(k��,�x��d�C;�4�9ǘ0)�,�����j�W˪eb��z}�2t�.���PCڼ(s���;������%^j������y��v꺵�{d�X�A}l�ɂ�����:Ri4��W´Z��}�q��Wz�~���M۱ޜv^��C�6�y{���1C�L��t�_�T�"���j�蝂ǷrX�t3�o8����IO��$����F���N���Y�8z_�J��#
��0�ݔT�q
1�d�8cLwKE>�M4'"z.$�H�)	}����!�+���넭�u�?��`�B�)?���`[Y~��a��j���3��Xw������w����dl_��V�>�YW�:�ƾk�<�[���Njh�}���^W����9�9�2���\j�r.}1 N�d.�YD:�ǪA;s6�S�5�8[��<;�j����g@ܷ+HK6a�6�����S�\�X�	)'u�R�������蜗�L��J����L:��o�o�2k�V��u&v����w�s�������k�h�,�}ޘ�Z������Oj�$Υ�*�@m�q`�aūݦ�R�iK������۾�������91U��p_T:Zx�倹����;)<��o�����W�*�	��r� ��'���'����b�zy��G�w�ï_������t�K6���MH�)ğ��_t��x��k��Vq�>L�4��U�W�å�x�&�2߯�
�s�Ug/�8�.���� _c��X���|��V��]�k�F�l�ېM�F�	p4�����k��~� �<=w��R}�)	�{m*h�3��.���Mc�ު�t���D��)Dl� ���V��.yp�[#�ЯW�Ot��j^��{������G3�SCyL��@�J%�T�k(/�ڨw��M��CXsb}Y��� ����r��<uߋ5�C�19�ʘ���A���_s�Z-r��*���k�aV�}��#B����禖.	w}ȡX)��2d�/#�x;�.��^����Cg�9�n���k5���Gr��r�aBV:��ћ8��=iJ�yv�_�(t��$yPf��;l�p��]���
����v����e�PNN�!t�k�N�Z�Ro=a�|�&���B�E*鞟v�zP��\P��(Kyi!CY�1U����oT�~>h͍�[:�\h�{��;��^�,:��V�.��_c��iY���ި(��௏4��'B�+s�W���S�X~������b�=�h���p'�K������{��7�q�XB�ІkZkg�p�2���_���8���@�)�Iʕ�[��ջ\��֙�ǎ�-sn����J�L
���^e^%_$`' �ۺ��ʲ�����,ŝu��){� �c�/�+t��lo��}ة}^���FwC�5�{��l��Ŋ�<�G*���F}W�y�%������d�0R0{nݶD�dp<�~���N�"�K&+L����f`w3D;q�ݨ3i�-�w��S�!ñ�N��$mxAT#Qu�L�]if S�>u,{W�W��-��:�?T�Y�u�U^�ԕ��k�	gн��z����w�K^Ҋ`��a�������s��Q�S�a�Z��y��Pu�_����
�7P[$8�˛|)
�e�X�'v��]�ǛM��&{�7̫�:g��ElH$,^[�z��h�wx�HŔ��F͔�V��u{����6��!#�o�W:�z����v�S0�Y��=�-I���Qw��~���`K��;5ŜG�P:=�>��y���I�,{���E5e{�E7�����n��g�}��԰w�c��"QC|�ѭ�E�qqe�u7��2U��!^�{�w�핬�Y�POBʹ��7^�uy�Ca��kW%��˳�j��{��݂,����`�yZ��n�xK�=��i�r��ϦK�7�\H�h�P �i����*�TߠҼ���r�g��R���<��v#�ҳ�Zz(oQ�P�7$&H7�����S�H�B�R�R����}���OgӨ�]��ǌ�S��3[��mܜO�5�;E`�Δ��b��'XD/���GE����:3�}d��XӒ�2��S�泩��Ȩy�	(��Q>;2�Լ�@T��SS���ߥ��a.�q�������G��fF�S�B��!��+Լt�Xܨl<��gP��i��J�o�=���fk~J�D�5�o���V�pu1>�JjBb�>���-�C�[#�$w�y���խ =YVUiu-�j�H+��7�-g���.Z����N�7�晇�{�����n�KA?a��G�#6�z$v�y;=��W_`n��K^���%K�ײ�Y�1ڜ���k��36W3:Wu���u������.E���ũ��Q�c�v��y|x��6�T0`\���:�6�E�^�H��z�����=��(E�55�bp(g���/:���S{C@أ��fS����5�*o�O/��Z�-ή�F�hYN�2�M#/�^�T$�`�7���,w�/dΗ����=弸R��f3:��� c�M֊�I�K�|zRX�����T$�K�������;ʹ�Ũ�
�l�<�2u	o�3�8�������|�&��^Z9z�Zq+��y�؟_k�ޮ��]T�"��J&X�;�߀�9�3���f��ʈ�'R�`����n�2B��6�z���K{�W_[N�F�j)��ʄ_���殞G.s�+=J��F�[*tMO^�s+չ�y :GA'˲���a�Ϳ;�����C�`�"���t�3�-��ӝ9V3�-�}�h�$��#Oi��f�a��\f��5�U���I�pu즣��i����A�S����&
����_o��_�}��Z-}w�<:�X����+؅��|�:W&C}W�k/��Hb���ש��m��,���3D>W�����D�5_��zh��r���v#t0�2Z�W@�ܳzur��7���{�6�l�<��O@՟:One_2ɷ�7��2�M{�3(r�l+/�95���R��̳Q}}�NϽ�B��9d�Cs)%C�ʕ�R���+�m/)j��Ҡ<y�POW�߁�N{k�@��S�0m�$`)�9�󴃾����S����X�9�7�i���B�R�U��f��� �*�w� Tu��t������N-���aQ4�2���J��=U�U�<e�wF�ǈ�OR�]�^t���݊Q���7g�wy�
�lnZx����xz�[-��<[U�du~0w���-qG��V+�tos�?[�v�Ị�`Xl�U"><M��K�痂Ҁ��/r�e���4�}[��{AF��\M%�������yKhm�4�>&x�\�S�
�a�XeFq��#~4�0��^P�L)�a��<j[���q��c�Yj+#H�WK֧.���C�w����|rׁ�[�#�MH�K��������f��*�]-C�.]ȵb6���-�w�X���"W�W�oZ�g�~~�MC7>�d�.!��N��њmP�W�都��<-���6�z���1}����<q��6$j��Ao0��{l�E:��2��(�L�d�v˩��ui�;-,��0���<��c��CJ�u�P�e���&�79h'I����m�:��>o���7�S���7��M�)Y�͡Y��GP��\2����pدC��F�C��ft!���e��e��B�v���v#Cu�����4�0���:�,��15��6�Z��r:�6؁ay(U�Pj���P�	t��!gf�)"���>�2E@8Oa��03okel�z"*�7���F�s��<#
���_'��l��@�	�+N3c�b�V�Qk3E� a�³\������7j���2�׊mn��%9g������*W�j�6�HX.���3��ǔ���f������V+v�jTf�� ��I,�V�~�����p��Dn��B#�v#F��}�,�.�7�(��'3�.�ӝ}�eH��M�n[�H��b�����A�'6��T��<�7u��V��i�*�%i��O��ԯgt���=��&��{ǣ�5%��ը������Gә��M(�V2m�Ŷ����K�&m�x55\7s��f���P@4KL����[�;W
���OaΥ��Ġc�@��,�ݮ�+F-6,m��V�"��|�gVn�*1�j@��ZJ�0��B���|A�������!]m�ۦ�rL�X����v3mu ��;�_M�����3`W,���W-��J��������:1�q7�*��c;�a�`�}����-2�A���֨�\��o)5�nˬ��Pynsk���h��YҵJE�/S�7��3VS.�>��s�
Ǯ��P�E����R����2!�Wx_	O���K���tf�w�"쨶�#wl��f�"sd͐n_)%ۘɾ2�Tۭˈ%���5�̻�hu�Q�p��)�A����3(�H\�L��Ý2gs�N��*�NT4�.��F��P����,�5�,�yi�;�Ȋ��.s���I��f��:�U.�p��F�IbBWgfE5�w�-%�ƺYw���|�e������ ^��������e{���n�:�p36��k�AeN0��9̽�̩�� �(���
 ��z��d2Zά�$`V5E�m� ���Ǽ;�7{mT%c|��+u��:<��VK����n�7�u�6�.#j,1��������a�؟��b�rQ22��������A�P7�Fj�g'R�WR/E����f�Ś�RG�f ���a �쏻��b��Nr����x��Cow]5�\���ưnX�XI5x6C�x���F̬�pd����TuL�75fh5+���nB6�M���۴���GOqϯ9v�b��ꔟ�/���л��/������{-�\7o�5>c��{8���$H��m��ł�1��[h*��b�,D�
6���(#"Ȩ�`�[iY+���Dk
�kU�l����Z
�kEV1Uڊ"����(1K���*����*ņ6*�QUFڂ�b�V(��`,b�-TDUb��U%j1�D�V*Wت ��""���Db+V�E��cUb��Qam��Q�X�EĈ �b�b"ֱ++0QcE����@b�EA2�#DTAEk.Z
� �*,�TUU`� ��X*5
��Z�
��*�)h��Z"+)je�[Q���Rڨ�̥�1���Z؈ �	� @|>m�n�8�"���Gf�v�Y�z�M]�]f��'5r��d{��ͥ�+�M�(�ݐ�W���F�}�fZ�|7����_p�%~ix�_xzC�{H�����v+�&x�y��#�Oz���c��e�SS���;�9�.���x��\�����i�-�;�\�bd���Ş�A"�����UP��V���
�R�Zǔͼ�s�I�ցA|�ڬt�
�l҈�y�Zރz|3�\�%�_�ꖴ�j���LB�2�,�����iz�B�{��3������՗=���4�.!����̳��+P�1&{�G�ە�&
�yi �5y9�N�{������4`���Z�k��!�M�&[�ay�m��OQ�+��}&VMcUH�<�+H�>�&�X�O���9jR!�?{s�6��`oL���4o��`Ҩ�6�U-��y�u�Y����;��m����f���^�k��qpu/�E���σ�cR�Mg=�۱�d�^��{�A�3�|"�gTv����#5!�#rǩ����L�ͻ�'��.d����Fj5xp~� @��{-�ϯ�8��6-�ᵇ	�g�0z��WxJxE�a��#�jr`�W��t�N��v��]:n�F>��3��½Ǭ���|��N�ٸ�y_YM�D0=�Nv� Iar73�G�>&�q,�������,�h�xB��r�.�U�}�(�Vk����������ǝ���"�8�8yl.�G�N	��%�k��pu�q"2��>6K����cx��ڤ�w��^��ey�M8/贏*��M�P�p�S�f�1��=�A�Ov�ٴ���v��S��"JS���V����6�3���C�
�;�;M2�}ZY��r���cڽQ���Z�'4���~\��jEu֗��xhtp.�$��5��˩V:9�ľ�|e�D�sƍ�hd��_��,`�{�7��=U܃҄��=eiam&�<dZ)*��ؤqn��,��=׮�u��'�q��g��(�+�J����ÅB;�kz�b���Ϩ&`ҮV �yJʹK/�F �߅��&��B�9�ܦn��Z������JǴ��v�4��lm�EP�.߭�3���>���ӗ��nU�9��w���;}���\�d�־cV���I˒�{:�(pM��[�b8���ZdPޢ�}�Dͻ��=���uG�W��'�I�x�)H���|�v�ȧ"��s�=�)�]I���ٔ�u����b��-X�ދf��!��X�/��2���G�l�P��m�(����p�yG[�{��Tz��>����7V�j���Nè�X3:;��Z�c �K-RN�Įb�7K�l՝b�8��z�����q�Lr����r �B��T�W)_�.��n�e�7��L��E��a�#c�WXD!�2��~j?.��Pu�E�f3J^�Ek��I���Jc�"����6���D銪��{=/��H����n�Q3/��7|�z{|1>���y�u���yzވ�@� �
�?b��U^�k9��8�X���γ�WrOgټ3xqF�y1G��<2��Ǽ,����ڄ����O�?f�m���_f_ri_��Y�����L��J�CJ�.�<uzY�1r�/�P���{��J�P`��O/�k	]�@�r8�*,��iuP�J�A��B\��ئ^�3)�������u��yF�?9C;V��U8�`�^�LtK�K���(^�>�R�t@�o����;����/KMC:i��3o��"�}���JK�)%������r�6�]��� �~oI3��E��ҌVd�R��	�ǵ
�;EP:�伔6��o�=�k�Od�]f��=H�i9��DL��z���a�8֙E�<q58�����=<��?-G䎣�R50�J���땖�陣����KvȪnb�P�Y^�2�m��;j[!*>����Y}':�y����N��K�&�{*���^��#.���t{{��1�����<�*��r��G��β���;X\��KkR��u�Tp;�o�V�Ff�a��y����е�s}[�:�OT*�ù�UH�H� 4��2��+m����g5C�>q��d�y�8��jF�8gEw������aن���O�{q
����y�2?m.�<R*�f��ٓ��E?[��zTž����&
�YH�JM+���J�}^�9w�1k�63OY�z��7��0?v4��R��9br�'�i%�)��)j~�����;R{\-/������T�,J�����y.�7]�xB�{�g��k֮�˙��o��.U6}��*��\3NC7b��},�~��pS$�x�"Z�i�+��@�e6��! [�p�c۟y\�Y���V�קP��֠>/c^8��� ��׬��L�7g�>�y�Jݺ��"���,�ޫsƝ�I\.�-����l�^���>M�z��o��~��l ��޹�Jݻ@u�K��ٍ�'*�����z��J�>t$Zl�Re3^��7:�qW�ge�oˢ���u���E�k�vzQ�Q��
���$n,�=�:V���45v�PݛjD'��a�y��.�Z������.��V���3"d���1��ض�`ҝt���bp�u�5q�S��m��T�����s���[�C����r�ix�[�:ҟ��x/4�3�>�k2���y��,���g5���'��	j�t=�VZ��E4n{�f+�����w�=FC~�c�.-���� zjD�z\"é�'�����W�9�z��Xݶ\�)�~�we�X��J]t�l��
:q���5�l�e�|=j����������.��T��ݰx���H���x�Zi�a.!�H�j�������Hn&g�l�E{K��`�f��������/ի$X�ެ���xؖh�iD|Wm8�]h<��ɪ�mk�m�9u�c��׵C�б��z����`�X��7�@��J$���3�G�"6Q�h���kϳރ"�j}NK�u�T�Ӎ8�T�-=2�)���k�t�Hs���m�;������k�\�e��\�|����md�P�*�ޔ"��b]B"_�ݷV�xm#��>{v�[�.�� +�o�����5�W���軫�u�bU�]����.�5�~�t0�/Z�q�����\7�8�P��p��Y�gm)�ǩVV\�Q��m7H%Pc��Fv�=�{�lX��X�폺i�D�{����-5%h����er�����d�v@��ͷ�)H�m����b�X�5uJi��A֥8�b=��
' ��8��MC�vyW�{U�'���u�-����I�Ȭ�[Ql�s�pg�͏��h;�{�I,����g���3��L-n�^+��ݜE]:���~*Z��ͮy��G{�Re�o�=����t#�&? ���b���xe\\&�]	�"����;����˯�+H���O�~<�\��޲��X`Wh�-ΗB�<��U i�X7���ɘ�שZү�T�.x���Xq"6�z�>�di�q{�~���V�����ޘ�ҬR�"�.#ʾ��X�e���S�`ܶf;��|:Xz�Is���qg���Z��c�!m���9v3ԣ#���5|��[hZt9 �Z%�s��i��V�e�w9B�����n����ݝ���o<�ả#@�|=��3�H��]1C�5���QR;�U�OjJ�鞘���3j�yM	�3�(�G���$�͍�Ku2V�{NZ�F��Ǡy��@a�OW��1X��%�|a�'��hk�Z���b�+�����ڛk0>
����WU�df(�_W5@����a��a�|Ơ�f��&��{��c��u}n�C�3�����yң���]5�s_c]4��v��L[4n���I�7;�-Cy7��е]���P$zN8�{��Mᛵ�Q�Ž玼!e\�f�(�����"�ĉB%�n���ǯN4x��^��KA����+�]������������p�2:��ə�=��+؆o����=H�t!i���Q��B��ꔡ�y|�G�fi� ]L\S�㞙�5G4ʵ���Weߌ�;bZ&Q$k�����{�P|���7"�Ө���s0�{wo�fy�~�^�~><�w��#��oލ�	�p���敞�X�j*o�ǎ4��̝b��=��[�_�Xq�-(l�����E��8���ahʕ�ȩ��iPw��3�Ը��p�)T�W��@�_p�2�g\�/������K2�<h=���R�^���#Ʈ�<�;}�ߏxY�b&��	!9�����[n��/_�t"q��d���l���'˝hp�,h�}�s5�ua�CG�x�߇Q�Ա����=�;}S/Փ"&bc�%~0���A�K�L�������z\�#ZJ�k]6��֌B�����Ve����4cϹV�Na�X���N�|e�s:n􇰼�������n���p�/@�H���a҆ӒY�4�M������1�{���j����dc(D��9���k6i�]���[T��N:ۢ�}ׁ��\��&���^05Ղo?
��]u����&:|�3藆=DW*�����z��t�k)P���R����'�m�8��"�]��<Zm���3x�7��㬘�9�[�z�-�����l����B`j[��#67�mu@ꠗ��g��������aɋ2G�x�)���a��D�8ОX�/�3~�5� �k��,�����'K<T,���n3�B0%�p6�]����}ow.j����1ɷ�Y�F���K����o���Mc��G�L�G�;�����OP��A��Ϲ����W��'X)KW�隈��K9ǧog��3�؞y`7r�0����Α'�/�������T��]L��H�ޚyߺ�ܔ�|&Aj��L[��&C�>Cba�k�&���u0}��3����0�ƥz��3o�{�����准$4ܕ����.����>��|���gfx�I�$��zE@+�;�vy�m�7��U�"�vbLQ#A�9�� ��lݾ���m��γwK�N5�&M�j��@��{SdO^�5X3"�+�XJ�P�{(2R���b�ч�3��ft����gGcve�|�}���{�omj!�U㡽�@�wj�ow��V���*��a3�ɛ+!y�r�	0�%���iu.� �ڴ@h^N���z��Zf,��V��B4N�)�|��Kܕ�)r��t)�~�si��ЅCR�����->���ƫVZ��*������^���(׻N�瓙�غ$4��{E�-[^��V��,��9�kƖ�
ߒd�Zא���*�ث�׼���H���;C�^1붖R�޹e+w�0���K��f6	��c�\�r�~�zTch�;�{UK��8�B �[aşS���	�ҹ�p�-���+�R�`�5�^��V�r�}��}/Q)�t���q���39��<~����H�W���ଵ1]v�GRh�4�C��g�#��Z�Qu��x�;MH�}�p�u;�.��㱚ֶ9iFLZ��m�Ī��EUoǠ���-CC�ܔE�{�p��ߞ��o�ل�.�YGq�t��JŢǣG�G�{��e#�.��t��K�v#��/f�7� m���noE�)VoXg��Oٯ3[΢D��b��)�V	3�����Dh��zx��0����������U��{4�h������)��ԅ�b���m���#��־��!�	�,�Ύ�*x6f�[�}��j�l�a弓�p����(�D�B�aV�t�h�Y�C�gs��-����M��-1�NM���
���p�Q��j�r�[�KSTOA�Go��D�o�z|z:9�^�.T"�Ա���٦PwHiD�T�j�#��x���1��s��c�G���C�🲛�C���KZo��j���192�)��<�C���e.�>�����)Lc_��ҝqj�P��9w��D��0��J��bL�J{A�2��C*�gd@�N�S)���=��+.3���47՚�>輭�^1�*�.�����+ַ��k���ˑ���!ؑ�%	�+���O��]�·��x:��tO�x�R����x�j��]��-����ak�
�S�z�DN��p���Cֱ}qpu.�/ǎ��׆���S����\����=�:�G�鱹��f��X}0*�ڒ9�<~�Ҋ����^f�3����P}Ҵ�����cK=+Z�&V����}��n�Q�z��j]h�Q�k=�V�{�j�J��C�����P��۷L�s�u�>~�?�lSL��{ll��i�NAۦ<c�!�7��\EڄyU܋8*,�N$��1��.{+�������R��fM����WP�J�.��(hmX
��Yӎ,�2s��GV���f�*7� �̱��Pe�����v;.T�hf�G:�1{dL�v�V��)t�n�=�븱v�cb�)z���ʌ����mmu�]ڽ��S*N΍��\��컦�$�(WDfCV9�����6�屔��K����U�
���ɲ���s:P��}D��;�ʔs�[Q��X]u�-Ի-������W���#sUw;��^/� y�Wt�t�ȍLL"]O4ei�V�~{���[��U��׾dms��_� ���Џ�3]�(N�c(of��-1w&ҽ��qUQU�7�Rn%k���egl�:z}����
�i+9ޤ��»�I �C���d���-FMk��b+��dLpyJ�t�'xV�<�t>�b��q�'��qF�,Y�v̲�4B�7�=z�v��ݜ���rp�RJ�I=����+p򵹇���k.�U�X,��7��N�l�r�f�\3>̛���C$��>�r�ˬ�f�N]�īc�[ܩ�P���ɺ�Z���tV��A�`�2� !)JJ��yl�Qb{��)�=B*�+)�P�\���Ѽ�TL̈́QB���lTcC��x����S�o3�-���h`Vɝu��ʜ%c��^�q��\�� '��gD����3/qu�h���].�[O�1���]��p9m�A��@�*�I*��o*
��w��d�sڝ׹�x��D��ó�չ��ZÜ��2.��s���kU}B,�3:��ro+ޙJd]Xj�0I쫘�vm������o�y+W�hw\�����l���r�2z.sX�6���W����Cͧ-��la��k[ֳv�>�t�t؛N(g>�+�9�wm/֏XU�=U�����+��sA�����`��7Eu4�f�`���N[��2PQ<"���R�����+�.�mj�F5Kz3&WI��[�mX����)���� g�η��T��j�}Z��Wn��I����Έ*�T���"[:��|[��r�W�������r���ق�G�Z�bo+Jq�O^A}�4ݺ�-R�*�ˀ�ED샵�L=�ԧ��u��%u��уWn���������ڋ���yD1��t@W�N�������]�(jUͫ���1O��Ԝ�K;����+����y���h�H�Н��S�p�i�*�X
�!�Wp!4-wW	�f����k[���e=�Uvk�N��ܭ�=v�Guy�`j���;,�`�J�����V�����X�n��;Œ��b�V���շۛK��r�su�*lV��ѫOS�7�&h�Eb0#�� ���غ��u�f�����雙 �Z�x1*>��ƍK!�!S����.A4ܥK,9��"k+���ة�����!�{]�����u��Gf[Ak]!Q��o�C�ϵ����o�o�5�ϔt2�*#�����HV�j*���DQ�1QPDUUb*����D�UQ"6�T��F
ZbAq��̪�EQ�1
��#b�DKeUb1T�
"�EQ����b,*����UD�*T���eEEQTV"ĭTX������QDQq���J�E1��&P��B�-��JV*+XV�(�VQ�TAE�J��icAUE[e)kX��QUT��Z-��*,�T�F,�E�TJ�Q��R�lU�F*��YL�-s*�G�pJ�ETr�E����U��k�(���b��Ŋ�8��KZ��#QDQ�ch�-�Vڠ�ڕm��`����QU*�*�cU��!���h��"�ciq�&%1��-�Tb�bĈ��b[bʶ�f"��X���X�����naG-H�K�Q2��)���5��>��u������y�a9SV���]��s)nm*/�!YXU��a�XOݣ��]�&�x�n���2�G�c��6w���޾��}1pȣ#���	��G�ƴڮ*�.���kif!�W\��ke%��e�}5�k�<	��L��a}���*լ�G����%��ҡ�&�|���!��u�X�����'z6a�z���(pU��҄�����ki4A�"�U\a��z�OrG%<����TEJ�V�E5{�b���<�`��B�#CSK����`�´��i��z�=�{҇����[H<�bskD�,��s�+>����x5�'�ն3�k�%�{fӮ���0Z�i�-��؟�.j�k�E�e9|l��Μ%�z<�5���0�zߴњ�C�����#�� �e4�
\�e
g�w�%�6�x'��J����֍�o|���G5����=g5�0(���,��$�iqYI�ׂ�>W�o�zu��{��G����^���y��~煊����{>��:,zu	i]�x�,����<�x�o~���I����zv]�'Y�3z`��P���c�֌�%߷3־�X�wE�.D;�B��o���������*Ƿ����):W�W	�>\�U%���ɦ�dL�KʱX�X��|���\��Y�:hKz	������coP���2��u�(:������/ޥX��D�q�ǔ��ݽ��6�K]L�&>��_G��nVn�⏏�)��{۞/W����I�*9a��Ƽ���r�˸`�ܔ�=E}{�U,�m�(e��+|�[��o�:����H�Bs����2�[��u��a'�\U_��m��͞�t�ᒗ�h�q�1�x��pz�������oyv�����/ݣ��K�`����^����7(úU�Uz,�Rƫa�|*�<G��.ޜB�n�1
�
�ur�kg%z�/�z���y��ŉ]ax;���Ic>'�	ʞ�AFKt�/nÿyTq�7/�x0d�&��P�<�R���'�m�8��o���c���q��xv�wW,��x��|n��LW{=���c�<�2u	a�'���7�e?���^]�Y�����4�����2^|���H��@���ȑ�Ƅ��J&c����P���k�A�k~oy�6�Y�6M��$�'{υz���rw�6QM�	Z��%����yźC�*�t�M]���ٞ�y�{��ɞ�L�v��P<C�j �>g����S}�J�3�� lJz�%ȿ]�o�7.E��CT���0�o��a�V$v��5}�5��uy]�9#�>ѕr�2�p�+UuLp:ʘ�`pCKL�3i�Q�OI3;s��Hӯ�ս�5T��Rl�u��*��9Vm	Ţ'W(�y��MB<�z�����=M��s�B��޻F�L�Ϯ&n�aBY�k�x�@�����+�#�T��/g�oCo���:��%+���}9R���.6 �* D/���$�E��b�w��e��p9�MA1�������>\Y�^LJ��R��X��O
��RK˗_�M�S]yΧg�Z�b��u�U�[p�Ö�x7e�=ҒA��U���<�G�u'�f����hə[c ����.��R�k�qp�8=�� ��@��F�х�6�T����_�wE��&k�_;�%�ؽ��V祅Ϳ�+�I�^"<�=n���j��zvƶ�l�s�񞎻�
=�mg�Գ��Un�xJ��o0�K��[�5w��1r��ߕi�L�l\��S����ֆ?a�-7�{-��M�{�P��@j�L߽��Ƴ�����.�s����Ǥ�/32<�׵�1��Ë>�3���z��n����b�A�.���er�Yq�bK}��;�ܠ��Xβo����	>��O������{脋�^:�s7W�n�WF�4�z���Q��T��{�+7[-]uy\��N��FvH�S2/:���~�o}<.�l*���1�X��qJ Z�{�w\2��6�֑���9��M퓳��1d�M�lڼ�s��p<�wIYw4<�]������Po;y���[6����X��\)iuH�9)s�_�u��x�+�/x��z뇞�T;�/*�eZv��Z�V��P<�1].C���7��u'b����@Q�L��=5�}�	�uY7�DJ][d�׃�f|���O��e#���G��5'�~H�j�������J^ldT	��b����&�%�� ل�7�Q�u;�� �z]#�D�D�:Qx��C��mЇK��T���b�������؞�Ө1��z׀�P���:և��t�89҉{}B�K
��*�0�4%���m��x"�w�����Ȕ:��-ie�,�L�~ڕ/�,P~��(��L�S$޳qt�o/���x���S-XJC9ɽ�z'-����l���%���|�ډ��s������}��T+�ݴ����%u+��p��Vj��u{�x��ak�*t��ة37�Y�{z<}��gh���!�%Q��p�CptN�+j��W���tx�]4�h�g�3�{IX�,O|��0PpS�w��,!�֑s�Cֲ5���<5S���%�N֮�B冺2�vLͻq�n�����K��6߲{RWMC}�gHiԯ[&�g�˂�p�a梍�AT"��&V�%xV?KC�Ս�����v1�ݮ�Yj��TS�BR���r�R�N#q��:���;n]���c��T�۾���t�Y�[��^�wzGN�,oD7޷�!I��E�ά�ӷ��/ɥg'�T\Z(�6��ʬ�q4�����c=�����PJ�/��X���ƖJֹ)����o�\�w��B�vR׭Gh�j{��֝R�cg��O���[k��H���υ�&�}��Z�ד=�Ĺ�/w�^:ڇ�s^2��/�GE6Y�R{ ��f��y�c�����N� FxܿwOLX�߄Z}Գ��
�F髉�C�P`��*��i��G)�~�'6nn�N��KI�C�J��~�x5E�uFF�G��K�EV��C��qOX7���E�ӄ�/�˒�OR��L&jr���C�e�<x
�\mm&��W���2����t��+Mϥ�E!Mt>���M�l�=q��y��qA��45����	[�X������>���AAq���c��5�竢����<n�sYi���0�Z�ҲX|�����$dIx�����R�x
fw��'��R^ߏxS��^�fڼ�H�y��@9��,��|=j���Ĳ(m�X4��8{��ʊ�T�Ė�5�n��}d�ٖw�g��a�����1nk��^m��BK�}��6G8�,�oCnu&�%��9������z�J�e�e�m5]|�c[�)�y�xgT�`�F��s���Q�b�l�� ���Q+��vB���\J�G�|�G��`5o�'�Yk_��?t�Z�ô��rz�6��lKD��6I�t���Rqu��|���ȼE��>�s�vn�������o`FEq��}��CH�0Ú%�a���h�:���3��Fc�K}�N��u^�T܎
�]f|n�Y�ȿ]�K�'*N$��(�hr���2�~��^���^���u7���"�B�ͦtg����ޗI>��9C�9^kR�t�x��nK���r�{��~K~��_
�2���S<΋�V�s�a���i=P�=2��ٔ���x��V��#�Ǹ&��#��9�lT��5�x��������fU{D"�2м�;K����;�Q���x�2j���b�E���wU��b��.����}C�n7dL�wC��{ȷ�=b-P�J��w��^���
��/W�1�,gҒ��j��b��E$����ԃ�~��YL������oW��mP�"�P�m+N�V�A�.�s��ȳLz-���<ג.�e!{�mo��j�H2�^%���z�\���l�A}�g[�[�Rcu�F�6;����}}F�����E�X�Ѭ������׀��nA4v�c�Eڷ$n,b�uZ���f��\������j�I-Q������$�:|��������W���B3+��}����mW�*���v�r��<�C��^�P0~�H�����٫��'�lN4&z�J&,s���J��jܫµe�S��g
�8����C��Di���0l%�L�\^_[�Eԩ���n���7!�/������k�0^�xVz��׎����0k乨�՞���۹���]ʹ^"j�A����y%!�/��1%K�b�f�KD�D�:�&���xPqyC�T܏Q�{�KnL;n��k|��0k�y�?|eՁʘ�=�!ÓCba�kUy[[���%�;_Bu���C=_<�|^ȿY��O8�Xxb����x`r��0(U���/��_�^w`�'ϑf-Z)\/L���a������sл$���0[�����Dc�}٬>9�T̻��\V��-yT����E.�Ӄ���2����K�cG�?w���J��9�u'�g݂������!/�{<m�r�fKsƝ]���+�����ś)��f�#�rוW�9\{�&��U�fv�5�qΜWl���~�'v:��z��uBc��L�/���j��\����)����95і�r9xѾ��r�.F��ЏlK��f5�R��[`�S��M�Ѿ�{����5m����{YtYPo�����8�z�Ghҷn�&ط��+�"\/�������/)ބ�{j�x��2��(<7,z,��oe��M�{�
:hj�L߽JJK0��}��\�̝ܼ��8�k�}���q-���s0{�8�W<�� t^R���4kY%�Q�.�N���ʨ^%�JܖM_
���Xۦf;������!"�HU緆]hْV���T��pNEXZ<|+�--���H�H�K�_Χ`��o��tW�W�6G���{ZgњֲeC�+-r��#�;�l��
:12ҿ���nج�7��WJ{ݛq��9���>S�����k>�H�˴x�Zjiq�DsV/f`��ջ���A�y���2[�[\���V��md�`�Rѓ�#�
��"����ɪ�Ex��;���E�%Q5�'�Ul��i��!s���}2��,u�ݚe5H�5�y�n�%9����KOr@�oy:m<(u�*Z��={옽1>~^��
z)˚���O�k��!<�4����:�`�/~Tf���=�y�����qw <rn[����2k���ߜ-���v��vX��w��*����Y��A��V�(尹�W�W�>�Ѧc��=�d�`c����s�G2�T��u�+zWu�ovA˯�s��ɶy�.ׁ������Bե,�=�oh��OB߮+P�*���9)���k�����h[��>�Bxut^��g���r��>o�e���_��tY������ɵ����^�բl���*�&H)���6U
ɡ�+��W�{U��D-�=W�O6s���at~Q���n����)�"�%.�]��>�+pzD5�����J�|���v��)]��w�w.� ޖ5'�P�f0lOag}qߎ��ިB!o������[F?��z�گ�@��b�ʸ�KɌ��ؠ>�ZC�({^�iz/5�t�i�Zv�����N��&�/;�`Q ����W���i�:i���<uU������D�̋�	WzW{�z�j1��߹L^�Lۨ��UK��L�%Ryp���=��m3:j�Ys� ]%=�+�Տ�����\��g�Yh���,�д�rA�2�K����l�TgFXyHzp�n��"�qJ��S�:�f�'5��������i�e��})Z*�':�V	~���SipP>�`/�3�������,�ǭ��:�NR�KzI+�={��/�<����-��[��o4.Ѱ�WL�����a��.�E�秗�bC�At����/u�6�z[4vB�!K���.0�����ܛ���ܺ\�<'-�TN7;R�B����<x���59C��yM	�&c<r���4T(�*ۃ���?�����I�� �0��T;c�")W(σ*zg�l�=q�����bqA�(�og��
���v�����(�E�)��PL��9�uA�bsk~�����w�)\�k��.�cۢ�㒷	�I;(v)���T���$���˱B������T#_�E�g����>| ��f6w��0�.v�����38߆Kx��!�t!k5�\� ��|��\��wYM�u�x�q���w�*�Kό�~�OB���-à�s��]#�:�u�N�k����j�~{����Ru�>�`F䬈<$����c�ë�im����9D;I�*A~����0�Ƽ�x:2��u��L���B*��`�Zс�N�%���ו:u��{68wվ�\�(�{��g��B�6���yzފ���) ����lɃ{���*��Wa�Q;���`BAE�eb�f��)�gE��~8�Ꮲ&����S�~�p��{)����d����ƚJ�5�)�ƧF�rR�<�gK�ꎍ�e��j��3V�Ԙ(.�����<����sZ�Ɉ�]�Hr��R�k�R����s�Ĩ�o ���}�I��J�� w�ՌJW�7��9�1%��p�Sb�h�m�8�D����%v�;Y�76�XwA��ų��������F�U�w��S�Ruw�a��e�:;�X���43[��u��Hz�5��U̗�]��KE�̺�,	�%����m��<u���ǵ��g����K�FJ�H�wo�[��_e\\K�γ�6�P�ĩ�ݨ����)�g`˭E&"<��5��9X39]�@�sln'.�Ν�4(�����4 ��s��d�a��%��]n��Ň��}O 8(u��4O!�).ճ�^����5um���;w*M�Ly2>�,R|�Q�]3ul�8,�c{��xҢ���:=&L�v���Q��P���aǜd|�9g��P��Q�s0�h���S��n,'�u��̹��<ݕ�3&8r�ױ@��_� �n�_W]���r�9V�*"�U�r�*�c�׆t�-��"�/�}
�6����������TH,BIʙH�JTT��rh"��r���ǿi�v^n2�ǁ�F��ǣJ�k)�b�}e+s.C��hW��_>��L��e������.=�����o|��4E"��`Wh���5k^-V��p۵Vo)�f����5z�t�Ճ�ECvu�Nd���oi�e�8�V�r�[W!��F�]�o+�t��݃��;�uY��G�P�5��IGjug:��B�:[����h�dAr��*7K�1�rf�ػ{z���)bI-��	�e�;�ś����ӧH�jy���nܬ�!����V������fr�	��ѓ��⡥0]��	�f,`�K qh[�T�YЁ��铦��cК��/q�����K�k��2��`/M��B��������CTd�t�}�;8��='v�V�ie:�{���l��tP��q�D�%k���6���k��7��;�v��6�q�m�-'�U�䯍�ǱVA�&�:�V�c�Q3��9�G�������ngS�6�Π�m�V�0�Z�`�w����I�c�h���ѻ���|���sr��0<�#���v�t5Q�9�����#��y��D�Cr��13ǐ�����͗ك3���I#�[Gb6/O
OT��ZԷfL�T%cj.��xwr��y�#��ȇ�R~�j�ZŻ��#����;�l	8\H�T���CD�ͨ8�y��9��;���3h�n��T��6�B�r�߰�S)��kl!���o���e�CQ�۸�uϫk�9gC�u�JC6��W���A��X�]�4�{�l���U�����e�j2���i�o��r��N�	F�y����]�h��"i\�ޏ��v�=�{�߾y�,V"�9J��*�A��$Ɗ�QUQ���",V(��*"��mPA��PUQ�Z�S�[E��ePYm#V�ŗ��D�ƪ�ĤjUTX�DBխ[�q�U�����Kb#�Q"
���U32d�+Tq,�(�[m-V�((,�bc�����"�Db$�*��PiciQF�b��X�L�����1*"�8�a�E-0� �"�E+*�(�1(�*QPKaUDQm��R�����-J�F+2�ƱQej
2�c0U\�V(��Q@m�֢*Q%�șB�aUb�R��+"��h�T���"(.R�eDP�4��0��d�)h�d-)ccm*��eQPbȱVe��p��b*#��ڠ��PTY��
�pr9eA�E��*��fe��G-U��\���AdUQk��"�\�1Jĭ�1[d�������*s1�j�J�q�jT���<�k_��ѹ�
]$՜-��t%�d^�Dd��=<�fo������I�I�JW�n{�R�Md̞�v�G�=��\"�]�~��lvpL=y\�R'KڱJtb����mH�z���u�˹���x���s���L�����ɨn� �ú�QgF�]�������A�����ç<��f��/X��Y���jf_�Կaσ�/}sZ�nk�C��j�ʭ�	�1p�/9����oo?WZ�Ҽ@/�y&�祖�r����`��T8���P�w�u}�m��v��ٌS�{eT+�b���Q�(I�H�S��:�fS����b�]�ǋ�Ş1hO�^�ҩ^���U�M)�uYh�.�]�n�D��ő'��y�d��zu{��R7���.J����՘;�w,�Di��6��0
U����Tqܹ�/T#=]�%�`�D�Y��ɘ�r������m7�7�v�L�vû@��0q.jg�(N�74u�l�*þ
7��Z�#�ǣ	Hi�y���,����Z&$��P��噍.�R��3*Ͻ-�U�j�*���S�K�5��W���2����L[�ɐ�ɂ���DߨT\&��-�w�����i���n��J�r��o1�t���{�E��}���:�k����6��Z�)Pj]���s����*u��3(�O�<��~W¬ټ���]�`^��хo�tОܙϸ%\���E�3� v���o�m��󆭗�p�RX+Qb�3/��oh���zz�W,<1!��/`��x�>8� ����o�J��k�L�Ob��qV�69aأtZ����vI�ӽ���wU�e�����!��甴�X�^��_p���B��6���p��n�w�T��b;��c�*��A��o�MN�5 L�G���8�r����Qmi�I��.�^=��׾]�b�]w/5��M�E�vF����}Ȋ�v��m�x:Ҽ2|���X���xήt}[�7IUS�w�`���Ƿ,z �^/ҹ,��;����(��'E���O{ok3���l���%>Ψl}���q-������矽/���@/hgw5��שMo���A�gŬ����R倹����D�ǢlT̶�����Qޕ���m�����[����u��g��V�^/�^��+r�4;8���ԉ`�]��ų��*�a�R傤ǫ7��G��c5�dʇ�VZ����}J�̽�P!�%y{3���L���P�khd�}�G�=��7��Ƚ<m�x,]uu����92�vp3r�`1�+)�.jt���&Z9ʵriy\�� ՚8�/G7�aݽgZ%� ���eQ7|^w,S��\�-+��.��r��CKӵ�sFT��=L���C���)�k�:�+����+���pd��BgS��f�X&R=b]����P	q�DsCKU���X�����x�1Vzo� �C�����ޱFө�X$�E^<v#D��^�9�5�uI��hVuO\��wN�ó����ɫҫbz��t2s���eB-_�X���f�����f���\�kq��4��iX����dz����:m?K�u�
�zYq_�OT�,�k���D�Į/[�9�]�S�(m�Z��H��P��w{�.O�{d�Y�P��	y~����^�HV�>ݶ�t��i�꥕�L�P��(K-$5��z�q�U���|���֩[y���o�)�N�������.��q�OQ�C���edCk@�3�;N�.���ߐ�<���<{�{�O��#3z`�a�H��I���O}�:������kh̭���'n�o����.�����:%������7��KAb���8Y�ߣ�(m�uҹ����_f���V{o��o�y�x�1�.�@s�i����igޕ�rS�UoC��h�^u㽇�)���@k���3#� De���^��s	�a���^�6k�m��,������y����}喝N��P*yT�ˇܚF+x��Ƿ�6�;{/� /:��+�\��!͒n�8�>f�]�.\t.�"<yTb� zN����tk���c���#�َ�L0+����ӥ�c�������T������Ǡr���:�A[r������f,҄{�7NT7��Ƽg�p���M��VS~�W`������ۈ�2���׷�������^H�u,�9�^0��?�3N�*��u
��b�����^3�zߍŌf�d�P�_ե��iN�8K�����e3�+-6>Zj�҃+[���Ξ
�ۻ.�C���BX	�[�QE��L6��:��3禄�v�Ѭ�7c-^{^�}S��zﺞ�H,�I-/n�����+9�᲌W����0����"�^��c��I8MV=ɣ�:�b:�b|
��@�/�٦�<-�'6�OB�9��*�C#��n�'EU���^��5��C�BH��]�k�\���e����ҏ���(%㱱{���4�s����c���.�L�7��!@��_}��J�s]���!ا�	UVUk�c���fI�\)��w�;��ð���8'�[�(�ب�EG�ZWRqu��*���o+L�峱�U�@,�l��$�/-�n��RCu+ ��z"e��둣�(2��yƯ8㧁j��|�j�X�ʏ:�� ����A�r�-F*=�p.�����fXJ�2���v'�-e�:��}h��DGQ���9S��9�s4m���7�{��Z��9�VD�O}�GA��%�a���觏���<A]�ջ/��,��G�kQ����V^|;�����{�ʄS�0\��`n 0f
J�Xx� Ky�ޑv���6{�!o�(����m�g�ס{�W��@� A�vm���9!Ґ��o����'�o#��do�WZ6}5U�yT�I�h]��We'�tق�TJz�����}fc����(I
LOO�w�|����fϼo�o���C��uCF3�6��S���v���7��r��J�&����4����[�Y��5M�m���N{i�9��C����'&�Ȭ� P%�����/婙tԿa��^�k�*��b�@|%����o}0O���ح���4��f;`B�P���2��=t�s΢P����'�m�8�J�'���%�u;���,u�ģ��k}*����D��p�IC��[>��:1X2u	�-��'yC��_�ޞ#�3�Ma40ʢl���8�����@�wr$g&.��e{��t��'�Y�_\��7pp�z=8G	��~[	O�%�b:��7K���%��{��6�i��cRWM ���_�0����c�fDeB��(L�J�ͣ/1�gu7֫Bw����^s��܀�v��e��juњfl=AM��z�6��<�>Z�{��Wɕ�f��]޹f�F�y&��)��qx/�⣁ܹ�e�UYs��Dx��>o��dd��B殞G.7xV}�Z���SK�� �7��R��w�-�[�fg�O:�F\��j�!� 9ǘ�}r)�X.&n*&e�"I�7ӑtx�Gw9!����X�����T���Y�~A�zܩ~��r�r�CR��;;�kf�R�z�A��h�KR�P���ٱg��~���O_�\��nJ����>�;k��������:� P�H�%Z+m��b��j���W�qB��B�˱<��8�t~{~�$`)�9檃�ؽ�2�L�����'
Y��w�ܪz��
��ʱ�7�[��{,�N�~%8)�P��q;�%�١
�+?o��+O��3_Y�k
�o+�����O�J�J�Pt=�?_���h��Z��f����Vb`�~���)�:�p�\����qyib��5��������p{
b~�����ګ'��{���b�
eb���;�V\�A�ڎW:�����]	�g"��$Uj[&h��F�ߨV���V�[Q�{}��r��&ԓB5�~�����n�\��q��ͮ,�]_lx�xv�87su����V�)���sj�,��J58jR9�n���q��30ws=�2%�	s���;d������qpw3�����ܨ��������r��ૺFWZCb�!��.��l1r�\�����'ݏG�����<ݾ���]<��5p�7ig�m@"����+-Edq�������..��`]�D����j�T�j;�f�ޙ��N[�d/w ��ϳ�ĺ���gM:8p�I�EVz<��@%�b��჉R���r���?�i�����o����jZG��.��-5���b�3qu";�c����O ���wə��f([��F����
g�b��4L��+��*�S��^��>�A2���A���MQ/D��ΡNw��2��K~��k�7�.��Y�Z�H�.�>�ICt"����si�J~�R֛���^����i�^�V����][�F �����(F������Ө]��={�.O�'�ȡmx��)�{�����Ny���V��%��u�xL׽�Z�w��:����0�Z����5��q��)��d��7�ɇa�3ȿW�\�{ک�km�i�Sc�<X4�=&��}ŵr�-<wQU��"%л�*�
�:[��J7�*ԭy�_�Aݩ���]ۄ�R�3xKR�v�S{Fe�ڃ
kbNn�#�d���Ԫ��U��;�y�V6������Xt��}S�h����U�N8)B@J�!NɡÅvyW�{\�r�>��9��,L���a�r�WczX�/�ۓ��1y��pS�z����a�"��l>I�E�`�/=���V�nn+L-���ݜE�=�� >��=���YՂ<GMZ�/�y���w�Z�{�T��(/���ˋ��n�/�_�==�=��v5��
�s�(�Yֽ+N��_�"� =�,v��+\>�J�+��Go�E�����ވ_��B8���ܥ��##wC�K�O�ڭ��E�jԮ$x��L�*r+�e��	T)���������@6�.�gptA��wR�3�T�=�)𥶅��r�V�U���[��@)���_���Jw��Si0�ӵ�UZ��:.^�y��������hͳW�f?n�!�U"�,�Z�sQ'�Eza0�jr�>�yM	�&c<x����Ms5_�'�y���1J\�,��\c��슿������E5x?e�i�C�
��8�	�sv�?O#5�f仢�|c����3�S�z�2��CY��Y�MdɱJwӞL]�B]�����w!V��v;桒���j :L}�hvu�sG1'��I��[ m�bV8|8���2�9軥M�F����5��20v�Ƞ��m�ѱc��u�S��/\��K�Q�ʛۡ��JF+��>����s�5��?!�:����(YO�4'k�^�$�0F�������m�Z�Aڸ���h�(����̱޶��&�#Z���Mܝ���b��Nw���qFGVt�����	����r�B��K��R��s��J.�t��f����Ǵ{����Wz{u/�pOB�����K(�HZ�q^����+E�q���\��>I�'�u�#�<P��x<1'��#�xC�U}59%��Tz����=���#Å\$h�k/T.b���X����{�zN%��(�h╯���ҫ�������c�7�VZ6vV�*o���g����V_}�<��E^�}���[�eK`�Fŗ����}�ƃ���d������	]h���W��vP�%�Yᛉ�_�}��	%_rmg�9r���7y��V}8�V	��e�Bք:� P��U��xa!��)Ov2�L��O6^+��Cg�ǈ�/=����[ڦY��n�_J�^\���p�q��okeb9+�8��x��"�_X�������`�ҩ��k8ؑ��i����o��&��X��Q�b�s��M<�SaOQ�m�U��V`9ðu'��^�\]Z:q�n����gw�ϋB�`�vz�x���qq�d�	�3@-+��㼨�i>�ɩ�>�0��T>�~��Z��u���/}bkP����5��z8:���/�<Y�;>R�`�gR���_
�I���+w3!�T�������R7sīɻ�\�+=I���ȳ�-7}U\f\�h�P��H�WyшI�#�|�Y�،�LswSn���0��X6�v*��O��.T_R�//�a��E�N4&x���ߵd[:(�n7����|ߙ�J��q��L48�4�K�`��DW���Tk�]��y���'���s�ͽ���������@\��Ȩڲ��k�K�u^�!�O?L�ƥ����p�_6�U���9^f��앨g`���b*J���������},�/:����CW�+�j_�+�0�ğ����	��1y��<%��򗚃�y�E쾹p١֩��j���i�zѥc�H
�%��Z��L��-[�=KɁ�˱�\ĳ�Ӽ��m$6����wi���<*�I.���+�����ñO ݖ��t����W~��z8��QM:�F�&?��e�CxeKC�B��ؖ�U�kHs$`��Qh��T�5�XK�c�io��:k\0���(U��#s�����)bx��w�q��M����a��x���S�ocĦ��t�f���/�E-������N@���u���R��( ݶ��S��»���mʼ�b��N:l�渐Q���Lg]�	�N��'v�r}F���zm�g�6�����/f�Vn�R���m�Mv`����8�鵃�b�Wc�pM�ߘ�u��N�{�U��E\e�DVSV���N�����v᠛ά�3UN���rrh��P>��q�x2������Vɲ$$�)�ަ�µ��� �tG9�D��]b}|���2�IM��R�]��U]�U��;Ge�u7�n�䲊�����+��5���V�%��TRq��&qXD�+�J����*�w�Z6J4Juk��Dͺ���̅�ƣ5�@�t�;u|�8hL���ȭ__et��ҟ*�7,�@�h�Q���,�Y�%u5��|��ŝ3�v��6>��Gu�ǯ���]h͍@8!d�b�d�(�Ql�����V���8�Z�J�%��:�=�im�u�N�-��L� t�¹����4�,L���YDL���B�ڒ\)��!Ѻ�'���5�m����3]����,$�S3�#s36J��V�뵑��4��O]k{ڊ��{���l����e[��V���]eJӺ��(I�'+���y:��ok/_H�t�1�4�9g^9J<kD���3gÈ{�RE�v�۠4*��{�򺖲�6��K����M�e�ԧw\2�{��w
Z�,J;sH$l��x��xQ�2�A�]jT�9F��c�u
��r�}X�P�w�uZb�ǕՅV���e��on9����뽾C���I2Ǚ�g�� �T8��JE�jSch������<VCل��9<�k_�:���t����]2�u��}������!�Ҳ�1�c�`e��r���k��k�L���3TO�ji��W*U֚��ީG�Lp��_8JzޤG@�^��y�">�y63;�,:M�tN.1\�׈oV�؛��5��o�jy۶�},�
݃��*T�7*_]���Y��:c��+�qA��:�n��↺�V�-%B-�2��p�d���Q׺Nd8ȥS�L��b��*�@d�|��]�^�����Z8-�8��KnbScT������
hM'�������j-�{pdp�i�A:���=Zz����3"�F����$�e���*�sYsT7@��a{�q�sU`9M�Nq�һ �P�3�l��vW��^���,L��^ݴ�}(ڻ��wj��s��m��xo��)䬬�����',b`�ܭh���R�fK�y���]]HK��ٛ����]H��cEs��b�%���z�̭	�H�+�Ƨ-`��V-cQ�I4�{՚rմŌԻz��w��]��YiZ**��Ƶ�a�5�
Q�b�1�XF�,�c�cXVж��2�ƣl��YP��e1��b�����Q�cYmƸ(Ԣ�
���qS1�LFق���jШ�ʘ�kP�,��
�U".V��K�)3,�\E#Z�!�53
��. [JŊ"��*q3Y\k
�D�V�T*6�ZT(ֱLn5fZ��e��e�jVTĔA��D��Z\HTY��Ш+l*6��V��0�R�ʃhRՒ���Aq+%�Q˙J*#s0�ar��TE�Q��P���(�L̘��9sT\h�Vb���\d+F"����(��L�EV2"����Z*5�mEAaR�DL�a�UH(��).2�KJ�!S-�\EPQU#2�L@�
�+J
����m �"���!T`�(��DA�B���)�?�燌C��n�KiK�4�+��N�i�M�{mV)7f:��&�Q%Y���ϵ�:�I���^=��T�����k�{�Ʌ��g��X�%0�s�R���I�=	�3]pR)v�+��26�{���x��:�q���׏��d��ЏĠ�IB:��;���
�;���S��p[[�2����xeӥ�.r=�ko�>u�!�@|P{��~y�lk�WرlËK\&�v�e��+��,ي�+O�$�k�+^B��D���^��wP�㹻3�v�7�:㱢�cJ����eg%�d��Ϫ�}wU��\�P��p�mq_ը9��v3������B���VVڔy�V�	��[��\:Z蕏C*�,�mK�I�oWI�5S31=���D�W¤���Kz�".��v5](�GM#�S�T�+�vq"�N�@����Ew�r\�{�l�E�S�O5Q�q��jL�{e�B��A��&�=����ӕJ�o&�^�wX(�1C�_�MC7e�.P�d��|��F��zU#�����3�췧�f8�7�tH��%�v*�����癛�l�E ���%>^�^�ތ�O���2\�HJB�Y|�z*޳�yǇ]猁H�����jj5���u~Z���@)����]�G:X�����8��gM)l������K<�><^e��-�v��9'-���=ros�̪�=�M靶�� a�emA�i:��na ]�w4�O')�;.�@���u�b��'����]K�:�l;�5zUlOV������zק��������I$��U���>}u���5�ú@�JQ+�f4�d{��V:m9U?0*Z�ꣷ�ȧ�o���d26����؝�f�v��(;<�s�ZK������B��˵ᭋ)/ty`��6<�q���=��<a��/B'����{¾�w��:��������g���/^�'&=}�q�N�2�]#"��@e[Dゞ���%Q��hN�r���wˣH���菕/]V4'��<�k���0R{r+<�����.�O�Y���Sك��6����x%�Y���G=zR�^�8�s�H	�յ��?6Y�pS�t���{V���^8R��LS�A}
�2����Og�^C�������,]b�z��{�P�t�� ������Ya�]������������k�x\��t�_����[�,�ndH�{M����O�پ_�׌Ä���n�
��o�>��K̢�� wQ=Aqqdw-��@��q�RY=������ѕ�Ì0K �����9�V(��\��NH+s+q;��;�ֺ�td�
X��4��;xe[&S�ީO,oR=YPm�i�;^�����j��UX5��j���e�`���}�ך��9<罪���R���=��*nӽ�v�׌(=4����+ش�a�wyO|R����n
`QO�p����L�X�,�U;������qv*׏�5��,8%w����(�O����J�b��ֹ����X=0�l59B��C��[pv�U���t�����}��o�|`�5�a:Q+��%�oݗdU��l���j��1!q��㴟�(#�_��=�cS)��<��C���wkU��X�W
	�|�5��x[�Nmo:��_�y�}3n^�ڊ33��Yqs�/g���BH���j�6��h&f���/�ۏ<���t6mz�n�l����V+/*K�t��	��<2[�(��B�D��5��3���{�X�ϧ8��^��z�(pM��>t#`J��������E�9r�ܙd�(�4�u���J�sU��2�)=N��v��Qk0G0#rVD��o������%tAMfwxCx�T�"u3x�{ƑC���;.������Yx;�����{�9P�NY갫n�٨a����R���6�t�Tk�+9���"C\��{�Sa`N�P���OZY*�R��1-��w Q�V�mvW9���1����@V��|��tt�n��)7d�⮾�w]5��\|*�ܙ\`�:;	ĝ���,�����^�2��``z7�Uu�gҵP/�#���]�K�e��� m��@W��]�[:gމ*�h2,k�o���U��/)�uU�G�K��
K~��r�lx��s'
t���:p���K�Bbz}�ci����#��`��mK�Om��K�z0g�o�6�<g<oꙮ�ar���u
8^Ƽ_�5�`�ú�QgF�-Vwq�k�[~r�am���5eF�&����-jf]5/�q���^}��kqY�MM��(/�`/67:bX{�_���ߪ��y\)p���$�]L��s2�oV�ܥ^��OzVKR��7��$8���������I.1��M�P�w��ϼ���g|f��^��O�.M��h9�����AcZ��@�ļ��r��R�.�]����H��Q��=�/�M����o��~Se�$�3~�5�q]���(VN��9���+G(~t�ˬ�s�Y]v�FQv��P���Ɠů���
�=^��;�4��x��Ed^Mb^,�hV]cB��w��'����-�X [uz�0P�n�:�������oC/]:5Е�����{6�f�gP���4���(�X[�5W�����u%u�-�I�l���Y����P�D�j�]۲,�����8��U2������Y�3x�wԩVkPk>�z�ז1���B�y���\�g�}q3w-
:����^N�g���������"M!�(8�7��|�yF%����\�����g�e"�
��cTT��C�0GF�0H����/�V���&x�/��-fŞ�%���q!8��𪺊Ӹ�r�Q�}I�Ш����[����":�^Z):K�������1��o5�^�V��ve����jHc^;>.탎Q#���/<�>�ZI��R�{XgW<C^�����מ=[�0E�bϻ���K&��,8)�n:G��L�Z�>�[�'��{(O;]TY[��/�Crb��y��-��<��:|����;G��ORϣ�E}���wq>d�s|�X�����/ԕ���;�Mu�GWk�^����p�%�t���.��q��]^�HX�:0;�|�|*�V`�gRȡ�}��\D�:(�c/�7��7��O�/tc�+�o�N|7K�S���JJǡ<p�s�R#��񄝳�[�-���)l�]WE*�iT/��	>������Amv4х.��A�5��e+����S�a�
�:)S��mxr�=��:#y��H�VS%ω��V�!o�I�;}\-3�����	�2LڎG`uY��9=��ͬ��tM�)�`.n�f��܃FY���^U���<".���Yj/��שz�Ϫ_c3�ӛ�[��rO�{y�.�X�����u;�U��3[�&T<��!妃6�M߽a�χ?NdWU���������'����e����K���>5�K�@D�x�%�y	���j�i3�����H��ؐ�����o���HOy
:�N��3���~��J�?<*�a��^G�m�'ܔG��,�qv�Z̚�%V��;��>�V�'WR�I=���������_`�Y��Lۺ@�J$�1�����6��:�U�zvӗ�^��}%��W�q$`�s���/�R��ıA��x�^/�T��(y���:9/����-���pv �}��s�î��g�2���2�&
�$�}��%b�q��u<�Kr�>�}����3�.�x3�輬�ј�0�2��s�=G��TD)�4%�������M�ُ�X�)��]�C�:�.�#3z`�a�H�ᖘ6৩t�|�Ьu�gՇ�m:�gf:�Ĉ� ��Ϲv^��wa^}c��.�糱8H��MA@H˾�|�s��B��6��u�WK���Դ{}�rWT�A;N�x��:L����������!��,l�zS�]��؏veB����:���J��z뻗j��ܽ�����CZ��C�e&sVZg�ޙ�]h{e%�,U���Iڗ�I��ޣ�x%}d9����o�P����T�Ex^qp]�ɯ�\�W\���կN�n���b��ޚ�i{��x.	��;�^�ݰ+��T��yi�/�S��i�SI���|�9y�������oTg��I}��~�7���4�|ˬC���C2�0/8Z��ڼ�����H�#7����̶����|,	�N�W�s�׌+禔��-Í(�5�5Hr���$��=�'�z�5��L�]if/�S�Q3]A{󷣐*�֓�}���z�^Ǐe�V��P�<1C�5ߞҊ,�L(?N�7�����*69Ji'vt�2q�4�W=��8+q���7�\dS䖏kHR����}gk<���)�%m��ז�	��r�ֽ�߮��!},���ݭG�,x�.$3@�y��P�j�7^��u��m���ܵ�F�T����2_5�P�K�D�R�Z�(��������'y[^ü�ϫC��mt�ʧH)��[�hN�Ȭnq��Ghp��mo*��W2���Z�!7;�1T��j�64��_��y���L�.oqu��)]H�����R�guŔ3B]�°P溸W39Y��)�-�7ir�Μ�.�iv���\M�Ns�[�^����:�gpW;�`��Ιq-9�%�X�:��������R��V)�̔�l�\[�4��y��J���]K���o���ۖ�g2���J'm��s���D)x���]P|��7"�Ө��>�`F��� Īz�*��\��p@s�,^1o^J�| ��=�
�p����YT�pt.b��;�Ř7�
J�r�&=�6��ܭ�b�����>���H�ҥ��h���@��|�.�88`�|)Rx̓c�3�6Ƿ�i���T�S���a�a��Z��t�Xܻ�>~��3�{P_:�H��T��35Y�����Ͷ�����.>2�}0���	!̧⷗��^�kB�U�0x��yVk�j{/0oOuR��� Y��<��˖n�G���o&����{������ԨF�#q=��y���%|dZ��2+��&��=���`SR���^y�5�F����Y�;���S��U.���Pߙ�=�[j%�� �|`������!�&��:o���k���_��m\�n�*|��t��"4F��9� �Y�d���:Ki�M��P-�>����Pxb��������� X��q��ڥ&�]J�JP�����C��:��3���h���}�a�,-�vn+����m�o{Y�N��x7���Ϸ�~�����P���󺤰>3䖏J~`/����;��������/�����e�[&Wz���bo�U���sJ�M���1����|M稙��x=~{��WN�Wo=P�P�S�J&c��۔9�98�rɆ�F	TN��9��[lo=��l����z.��n(��Eө��Z��r�-~G ��Y��k�{�q��D�
Զ��3��{ۀ���#'ܵ=Ұ��q�S}���t����b8Ȧye�ͨ�i��H��}��O>I��f'�"N�Pqf����T�0k�R�Er��V���|��̚�=~s�A�L�;ÓCL4�D�^L��d3�1�|���hK���*y����5j���uަ��u!��z�c\Bw�邡����x�\EpL�ڬ�)�����;fXH5^�Wop+��}�����bL<H�t(瓴���b����3���7��%��8���g2��VOW>2�},�ߝ�6�(G^8��B_݋���|��Vv��u�PY��Zݲ�n������`�}�t��pU�Ե$�뭼�X�kEbf�Jl��>v�qmب�*��J�d�byopͳ*9�%c����o�Yιm�`���AM��1�����:��;����S=χ����=3��j�$Xz�C5w�h~�۫���Ɯ�u<o�!��z����"b~Kc�Dm�[�u]S�F���w|�3&^Uf��T���f��[i���s{-��bp>ڈ�U�o\�}jz���ʦ������Y��~�g}�r�B�]�p-�"�9��7�s*�yt}a�yJt�w��'J��~�>���+��K]��e.X�̛�Gq*ӯG}O�b��\ڦ|I�U������'����C4
��6���p�yg�X�|b߈�!t}�)3ޭ�XMH��R%�T"�u7�ܩ��;��Cʩr���+׺��pg!�-eΒ��[*s���Q�KC�P��d˔<Y�'�ڟ9KH�K;�U������.�����3��K#�{�t���X9;~���3;�HOy
:��z�|E�U�C[`R����j�NA�x۳D�J#����]��� �d��*�'�OGC��֋�����WtI�����}��O��{SpU��_��~����i���}�s$��!$ I?� IO���$��IF��$�$�	'��$����$��B���$�	'��IO�BH@�p���$�$�	'���$��$�	'�!$ I?�	!I�IO�BH@�hB��B��LPVI��h��a�kw��A���y�d/���,/�x��t( �
(�R� ��YT)*���
Q@)@P�0j*��(�P *�����F��wa��*m����4�wuUY2�qKZ�M����ӭ�݂�����K�n����p��K��\�U\�  r    ��˲��c
T�5�B\�"�"�ws����nwwiۻ]��gI�U@�.I۬�wgm�U۹�w�r����u��$P\�4��ۮT�2Iv�7G:�;��;]w&T�"��jٶ����U��i�
մ��J$N �٥�m�Yk+e������&�%H����kel��k#A�Ɍ�ԉ�*�nK�cj�Vص[Y��֖ƱYn         �x�e)RP&F  � 120 S��IJ�OS	�&�`  LCL`LM&L�LM2100O��IḤѐd ��4����a2dɑ��4�# C �J&���	�A1je3MMM)����ߨ�f>�3�k>��E�&{C�I	����������K$�@��B}d�	 Đ��'��m>2@$ $�/�v��a?_�G�~����?�1�B~�,���(���b�O;�@����=����! ��>�vA��� h@! �Q��Y��4~���P��W����������+��I$�I$�$�I$�$�I$���I%I$�I�I$���I$�A$�	I%I$�J�I$PI$���1�c��!RHC,��	$2�$&Y &XH@�X@2��2�0�`I$���M�)$�J�I$PI$�A$�IRI$�A"�I$�$�I$�$�I$�	RI$�$������|��uF�O��O�_�_�%�G��I��o������������1F����=B���������g1'�`�
ɘso4\�OZKLB^�%�V-��HN�6�Vն���U�W�>�W��B��T0��{��xƚ�(�`�lZ���f�E+x��U^j!���Ħ��gu�3w���C"tlՔ,\*�,�'�����Z���a��}���<��i�ȯ21�[3 42���5��YX*�B: 9V8��ߕ�5;P�u/K�&�i*5��e[RV�"1���D���S���n�n��:�VeM~vڧ���
|r��,,|VU̊%�B3�n����!G�k+s30��N��Xo�1^��*��AWY�1�cn��&˘�Z%��=t�J�D��5����<l��I!��S��KeF��I �:Y���.�KH���C��XFZȘb�V��vv]�t¤�W�h%��
�;�,�U�7a7u��v�\b6���f�;{%�M�N�!mwe�`�kBV;ru�v��tnŠ�V��R�X�y���wQ9*,%��H�t>�
i�3-��.9��5��l�ہ�j���Q�+rJն%[�.͕ �{vIHP�vK�m��&az,�
�b[B��+NdJ������+iP��1 �X0��(�YYx�Y�,��]�wDc�����:�]b���u(�K`:Cx��ѧN�[E��]��F��;Nd���Vd�U��M�b���ON��Ff���G��w�5��Ͳ��Eh�k�9��t�*�6��"�c�BC�z�iٺk�^��F*��-L�"�Vo���ThS�����v��u���ܥ�=�ᬟuu�D3yy,,V�9X4'%m����e9��7�ʙY��#��ˋt���cY���2��.�������FC��ub�<ם��R�T�ҴA&�n��:�d8�CS9�n�,L2�7`���T�G����$�zae��o^��F����)5��A�]�G.d�] ���)�4�cD*5ذ��(7��h ϝd����e�L���7�Ә�_XN�:�i
��3� [�����M�h��������U�}lg*b��0�e�¹�E�{A�K� i�/�ʑ�-'�[�3s,U��ϭ�7�&�֔.��XfQ�.Q�����VR
�n%׿^�Z�D	�r��Ѝ�0̈h!qY�y���ȟ�yd�k�'E��w,�.]��X��T�Ւ�wI축��,E��f�Ww��&�[�Օ��ذ�֊�9u`�Yz���bh���j�hU-L4�Q�b�A-��)�CAŘ�ԁ�vw�)�Ō;�M6)׽�ee��o#V�Fk�m��!"ѣX���n��Tכtnɳf��kLe)��Q�mP�C۬j����������p|l��6�ׇo`�����VaeXZ���n�~9�h�1W+��Lv��e�l�B�!�Gzn�*�i�rG�&X)bf: fY�W�<�厵����/(X9%i��ҥ� ��tM�vq�kP¤�/k"źZZ�&�nS�ī�f�!ʚȽ�bց�f�k�e�-�$��w`�ܺ(ҡBk�*��Ыh꿱X����V�5a���÷E��R��x���V�4�`K��f��N��B(U��N+X�Gm���h5����nܫE��Hh�Z�%��^
��M*�J$)�r�K.�ŀ���P����-|�Q�j�t]ꂳ	46k��i�5����b%�aJ��e�U�Ǌ���t�����ոD���^�qX��Zce�n�\��.�:�5y6�Eu�1U������h�Ƿ0Q0�G5�Y��ww3,����@�����/K�V5�зm�=F�5���]�+0Kf�m�BȲ3S&^���t` K����j�L�+�B�
5]�<f�^;�0����0÷��iV�4H	�	�	A?����ռw�N�v�gm�����Mc�8�3�E�ֱ�}��?����5�s���������=�S�!`��ԇ�����1��K�<L@���J�
�����Ѥ����{3����0�jb�?b�q*���7��WY%��7fjk��|�a��%�[NY�'m]�}V����S|ʦb�3x��^�y�l5#.%)����{x�9�WX*����ԝ:�fe��}-i��q<e��́gG}�QxnX]�������Z������x��T��,680��,GW|�v�ʛ7S��mqZ��M���wi_h1�%�Ү��Ɣw�0>��<��j�C�R�2�r4V�h칶1qU�ئ��S"���,�}]7���:8�E��`�E���� ٠�G����j�3k�S�0E%�^�su�Gr��i�P}�7/�T?�������\� ���<��\��j\φ�3��ޫx8ݓ��9�G:k������(2�VR�$�|�_t���7gw2���� �W�j�~/B'5(f�n��{�"\Âm�)�b��z�%|2�����m
r�dc)��S���`
r�f�mD���sS�Rm�s��Px�v��e�2q&^��13z����1. �Z�S�6����-�:��\/2���J�8����nāa<���rK�Ř�4s�6Օ���������p8I�p�r��D�o���h�poT��K�J����Y�'w��۸~�r0��lٻ���&g�ng�76�7���{��r���)Z��{\q�>�(�|����Jr�J���S{����E��ֺ��q�˄��}N�B{��<"��T˲p�k:۵���1JmT�Y���5<1�u�vH�0"+x�f�/ڱ��E�j�2�s�sV�h!{�i��DT�l%�Kn7\oO��]�� ��u8�:��%�/6��+���u��q^t��騝��p� �����
��+e��x��u߭�2c���4�t�����JFv�z�`Թt�A�ᶹ,����<�p��;Ø_�9٪�3t���'m��{E�ՍoP��ӥo�w�}�O�%=�a�pj�@wY��G�nɽ�s�wQڌv�1����g:�`��k�Y+��5�R�^���ty�?�>adz�"Rr!�R^��y���	��/��a�@����)����j��:Y<E����^Al�|~YJ�מ2�'ή^`(��y�uTғ����dKyc�4�PR���{te;�[�xp�rv���m�2{����W�R��9�s�f�U1�t�,�qí>�.�h��=��J�d�v�FiĨ'#�T���*�탵�¹��`8\�x^�2#Z�N��0�v�.��VvT�yH���y�s%6�\�u{%b��K5���7@�X|�U7���g,m��Ysa5�3Db^�D;��Guض�����fg��`�1
��NƟ��;�Ƭ�W��جjE��f�7}X�ה�̼3e.��ut�;(�!#�O��)Hr�o.�p�هou�j��i+R���2ns$ܒ��CT�Ɣ]��F�Ԛ�D�ܝ�i���r���&����1m����Z/��^�SR��z�E�������5��H��Rrni�st(z0���l޺�7`Kf�pT�^)�,
%�S5e��ײ��V��e\i�3��2��Ӯ�BVh�Q��qi�u}�<�{A�u�+,�ۤ�dΚEYQ� �])du�wij���raݤ�ܠĝS,d���3�P�t�te#Ƚ��\��o8�uN�(�[�3��i������#�`���FSR��wVgn<���4�TP1���=};"̎�d�����|��<�*I�����C��Qk�0���!:]Ax�i���<�Go6� ����\�-��A���2v���݅���Ϋ��5rE���:�	?��'���W��}g�3=|�W�>����~�}1��  �>P�;G���͒��_O�����{�+Z����$� ? ��'��������V}�9�}d��gV6r�m�r��1DL�,'z�}Բ�oF$��(;"�v<H�ԛ�.p�uw$w�,��1kC�u>sI�ne�%�7B�^�]�P6�2��mc�)A9�c2�˺��yf�bYQtc����ԙZ��Xk*�wv�վ��cz�AiZ�o��ǳ(�r�nK���*����1�<p���#V̑����be�D#rL�I"��I$�&fI.I$��rI$����K��<�r�BU��"XY孈�����J\x�WtZ��T�ۼ�ib��]L��x���Gb�{�O,���o%����n��k]#����6��9�ZPѹZ�g'��;fv����^>f�ھ�4�cMSU.���(S��|.�'_ݻۗ\>
�W\*�v/5rރ0y�Ӂd�^�uo;Se$�I$RZ����	*��I�I!�M�I�q�P ���f%ø5���鑰w+�X�$ٵ��frS9se,d����e�
kgi�<%��,6�X��[��GB��et�tk���M��]k�D��v��n�آ�
��[�U��m����Q�f����Z/;��.�,e`q� *�glf[9����$�&�$�I:I�gnI$��6I$�I����{]֎�/'7Xr���y	��m�T�)�W%�ʻ�mSt�C5wG��/(����J�[��
@fv�[�V���eZҰQ���[�qM�S�X��,�u��s;��[�S�9�c��L���wU��!��P5�:�ƣ��F&�Q��j!KEX�)��X*]ۼʙPk�ݗ.�ڻn���[rT�I$���Hd�$�����I#�$�I�dk=X�$\2Ÿs�׻pfl�߮���7n�U�+B4���J�㣰���[����Iup8���R-��JWM�e��L���fD��;S�CJtL�N�'+�]�uzs30��C�qۗBܪ/^!���ֲ_�43P2@���CjN���8EǜS2�\Q_Sל�
�Ԗ��`(v��Ԯ�Fև��E<䜇�st���tf�n�U}!�4Q�46��}�)�t�T��ϴ`˲:W"p>U
��гhY�u7f��]��@�z�~7`
�"�=r�̩��	�]l��-gZ�Ѐ��ct��y5<�*c\�ry��Kᷤ:8��هR.Xn:��AH)��ucL��S�I-ʗ�p�[�I"+�c6�ls�$�u	V�˜�Q"�Zu�L��QA�_Wo^��M�*+�;[멯]��VU:�V�WtL�L�&�AGP�wYW<=g@�#���P��O$F����f�D]Y�E��n��
ڔ��b�C�#p6V�}4�j!xcy%�ݾm٥ѵ}���+)����|-2��{�	%q�<Ɯ�25���!�w�w˯;h�	�N�Xʻhlj���mJ6ʁ�����.i=!�f���[a24�Z���A�A�X�br��L<�0�MC&b��>YȌ�[Nƍ��-�Z�I]�g(=9�n9�ʋ:��G��^1)krP�c��[����ꔞe[��QT7��;���N�f\���|
 �w�b��k���s�/*k��ȓ¹ r6�Avn�I�����Mf�&��6�s����Z鬸QrV��ůr�*ЩB��}���;�C�����N)0;['�m��z��`Y�J���������Ye[�7:j:��!LԬ�G`״a��Jw�6��]�UG��hEX*�u�4�Zܣyxͭ˚�Z+Q���J�'�3�ʽ��;�y�] j��MO�ZtC���"�a;_WX�V� �n�͚��R�Z�Z�l�ڦ{2��ԅL������H���gNd�[Zֵ5+��h�J�2�J(e�).��6ͼV0eβaX�[������w	[E�t;Qwon)��d}��3Y5�eA��W$��΁��K�s3�J�&���}K��Â�i\b�y�{�o�{�ᇬ�����'В #$_���̀���|f����|���e�W����Q1����hЦ&
c��,�)I@��6iS ��I�	�!Si餙_�;�D5@���%׾�4>����*�j��E�ڽ[]��Y�W�v����(�K�W$nƑ�a;����P5k$<�]"NJ�iR ,Txk梣�K.i"�B��ݝS��D�U�,N����)=� ��Gt��R����:*8�;���Y��v����ǲ��/�T.J����pR��ұ��tG����U�(�>X�0�wٍ�ڽ�S�VL��VAUTբ���5���j�1Jj�[�k]�zDQ�*(���}��EkD�Tkb��n��gB�QUL����8�-���0Z�ʒ�E��[F�,�,P\0��aW"c��b�x�����͝�ww�c�X������%��YP�2P���aI�_����K��z�����/j��s.�[��D)���s�1���s{�VN��6�/!zR�so/t�J>���ع�i�̈rv�ŝ�"X՜.���a�B����ݾ�:^O7q��!���WY�&zE�k��_f�A�/{Y�C��u�]Z�54�[���V%2e�a�*B�)_ԇY�a�I�]4�轨�ZG�G)��xwk��e��*v߹CLD�8����䘺Vv�kqwC�S�]װr{u��.c.��nu�+�95%.i;oM�G���Gڡ�Z�T��xS�Vߜ�x���wyݛ�-f�F�����������>�9ˆ�Hcqr���ݺ-�����9�������_L�Y���s:.�s��t#nd��Ղ,X��6Δ辌��ɬ֟_T�\�L��KY�'5��I�\{�=Hn��l�uuoT2���Y]�̌(�-�ce���ˁR��̹1�3j�)�tœ�u�R���
�Yr�6��Ȋ�U���o^�)��5�fЍ~p�k-]�j�#8�Kq��Jx�*x�J5e�<�n��u�![w�f����T���c��:��j������Y�*}�rz�����Y3',����3f���T���>���x>!��kKAK����D�O�Kr<qI{y���J�k8b�z�����x��D�5)f�㵣/���}MdO;h�t+$}g[�uN^�v%R����U����X�R�3q�ZK����ͺ��o�x�l;r�{L�̰�`�{pXE��ʺٷV�3�7`��L;{�:C��ϗV�����K����2�����Y�'�v�y�Rw�ූ`����6�]z�]];�n���+���j��݊]X�G�h�A
�Kƛ5A�#��3Ɛ����}Q��Dbw�y�sz��0v��˻���2��w��>���~�G
�f�T
�"`��xUX�B���*��rb�A�Y3����2�e87N�C=y�=���x˺v��	Sl��A�s�����8�ݧOb��"����?�`�Ӣ�V�+�"��51��a�r~���X*c{B��&v6�Ж�ܬ,4�I# ��ݝ:x���3���"���;�=�'oŘ)3�񮖪�,1���g�*�F�x�>;u�2�.���Z'��1�<L���A,fa�J�����H�f��"�v��N����9ݗ�2���2˱w�hX�������
��F��3�y��sF�����|I���g��B���Z*�w:t˲�٭x*wC�x����(x��:�X�|��0�u��q�*�}/����&�9y��8�V23��h��un�W�S���a�6ΰ��w���|�q坪e闻�00�u��0���yC�s��S��۶i��U0���}�SW3�o*��}�����̯�V���h���b�MA����Γ�V(�����8�=&n��μָ��
�;M�|r����Z�/[ٽ��q:j(x�8�1����7���t�ƯJ� Vm�<uΑ�`�r�A9L!���15_lÕP��Q�7j�%leS^��uym�?_MU�Bɥ>�����wvK�{?����q��z�SxT+8����V
�,}���VφY�
����3��+��P�!��h��>�����ɾs�:zE2��J�ǜ��]y��:Mr�7Vt�Yǚ�	k����Ѫi�ř�8�'j���8��yל�oT�||N���R2�}��}��}Bҥ�:�|����|y���FkĊn��(��.7{N��k��u�Ǯ���R�)��5���kM�W�(}�3r�m�Iݕ��4��aU�t.y?b-��7 ����]�C���HQ�W(�L(9v��8g�S<��(��ݸ�w(AW��8�EV��k�C[�����(k�c���y��G���˙�퇌�eϖ�p�+G�����^@M? �*�B�K�`�����4'i�l�a��k��o9��զ3K�zc��l���ь��1�h׊*�U�b�kw:��Ң��`��<ɬO9p�{1:�;��`I���;�=�]o�c�Ok�6�џ˳ku2�� �̇�3;d��).�����-��5;����Wd1�gßYy�M��b��9�ذk��i�T��%�K`�*eVusM_\�����'�!�7���Ը�\��h�fa�7x�0�q�a�������կq�I��=]�!N@�6����M��S�+e�Ǩs3q,�k�N�+8*Sz�Y�[�乙�˯��~��T��#�%�GV�g���R�B�
PWʱ�:�Û�<�T ���u��Y�'��@�VrVۺ(�r$Ƙ�;��Y��uu��'\O鋥����n���NDG�1�ޅ�}��fWu�9Va��׆麆�db�c�$�]��� �-�o��s6���0up�@�bD�Ǻ�Ν��[�]o���z|O
o�z�+R[�L8`���k�r��Uh�YqK�{�]gP��(���Q�[�kZ:�hb�@�H[�kZ4���RM2�C�J V���D��0ʷ��T�����"֌0�ᡌX7D�)qEU������Zm_|gf���0d�26�����4�{�xΞ� e
��)��w��{��5
�x2b�R��:L97t�|c�=�9^wN�C�ȝ;p�lFaח��<���ͳ�^S�M�xͦ�t�����y���bÇG���±��K�T�6�=f�����,���z��u�1�q�C�ٞ�÷~]��z7����Y��^�m��L��"cg�q��wت6{���|䊇18�����c>y�y_U6j�g��4f�S���x\��Ze�����h�d��ݤ��̯�7_� �^zӽ��8�����F���Et�f>Z���ۗԹ���v�y����Ha�=|aY{�!�2̾�Ƕ���L>�?l���b���u�~�@��5B��$V��x��P;}���ί��&����3�k��f�N�2�N�!�\��bfw�m��L�x8���k6r�l���a���ߝ㏻��v�;j����{��6��N�c|�����:t&|�8�y�$흺J���sΊ�V��.�шˡ�Q�G���W�Q��ȞZ��2�ɵa��،��A�6g��k�(>R��K�:x�����}��g�}���*��ip�j(�o�>��A��<d�z�v������ޓx��4!��o���[�>sen���g��o�$�:<�����~�Ru�8<kӦz��Mf�N_{k�j�"ʯߏ��ժ(U��>�>zj�doG�f�ڤ*�B�}P!��ߟ���F���ةx�?`��*���pl?W�i��|��
���r�=���.]�ϕg��	�i �z�>HvJ~�RF]�|�&�q��}/�}WG?ez`e6�3��y����2��1uM���gn�9g���ל�~l۷mb��q@�ͪ�p�?R��U�h����4x|��PT2��<��]3�o�SY�d��k���~�С��P�Y��_���{��z��p�G����8_��V+�#G���xW
@��EU�</��\*L�;�DXv�3����|�:N�;Ͼ\k�r5�?T�`����+�EKߪ�h?����O�\��N=�$s�W�E�fc4uz���k��}U��{�>�uF�]<w�]R\���u�}�A��4�ѳLs��՘͞yq�q�W[�1c�4��8���p&���5�{�Ol�q��4���Mj�{p���h��Z�^��P�;}pÌ�(��������_Z��4Ə�C��*�ی�~�B�����i��tWղɼ���,�6�~_Y��6�����8c���"uQ�*���~�*`5�r=?EO�?SVL`W
����M�������:�uU���?6�K������<�灾oy�T*�K���;v���]�r�5b�����?ƌ���F��~M׆��5c�����~C��&����d
����W�Ua|+�5^/��Ǟ�w�<�ΙS*�=Nӱ鏼6��=�'2�f�>Zf��2��,�1�x�۶i6���x�;M��9���]�|ji�0�i��x��n��<�G~����]����(�p��u�s����8��n�3�N��]"~7�5����GxQ��0 È<��WWd v�xٝ��`|��\y/D!yi.?G�G
�s��R�ʕ71�}��{�/�<}N����5g�Y��=�}�|�b�v b�sfn�|gF�i��^��C�Sh���ߝl��_���V0W��ٔq�E�/��Zμ�]:{j{�<�N�=g�[Ǚ��������o����&	�7�<Ϭ�pʝ�Ǹ�&ѣWB��?;�?9�V�X�����ӡ�Y�R��w���;�v�Ker͸r��1/�߇+?R�P����*�1~K1I�����b�w����G[r<qI^�}����\�r�<j"������W�g�ه���f*W�U��
��+��s�)�ʭ�_A�;
��x}3��<�܍/��g�<k���������P�W�UX��C�[��������{�:��6�'x�����4����u�^�i2�'�J��c�c���|M;O��<Ոȵ(��[���C�OuL?	�)��3��鏼011LU~����>�f������_�e�_��<��8o8(O�w��JnC���*U(+�v�ڵ8��m��OO�b�O�nT�W�9�Շ���щ�0�7>S�=��f���/��>��㮃�Y���t�'O�Ǚ���Xכ����:N�?�1�
�>��y����f�
_���3��+5��k2���1��Ω��:�N��w��3�z��L�)�.��S���ϻh�}�U1�k*_�޳��YNY~,h�H��D�T�!�w����S��׿l/��
0�Γz�)�T�.����g�}�Ȏ#ڑ��s��r�K����-Gr=T�g�+�Us��f]'�Rv�{�~d��<����{�=p�J�^��u�w�ěr������ꇉ�����y��C�<g���a�u�`���7|�x�f�v�<ko�l�������dd���D	�������T����ez�T)��eG��=?A�P'�S��}o����=���e���V{�<z֍3��i�z��W�Ϸ��9vok��OP��m�`f��:E!5R}	l+�Iw1nx�&�`�U��c^�YPd�8|�e��7&
1jЕ��n����v��G��7�D.V�D��F:y�Y{���e.n�\����n�d�.�l]N܌�W�5ɓ:�}��qv)�h�܊��m����b�s��.�͕R�/:�T�*)�?)��x/��d���oF�cY,�Jg:q��k[��u����ن�j�@���C��{�S�ݫ��\0��i����]���� ��Q���t3�0~�i,�nd7�-csL�ٽe*l^���X�BWM2�-�}a��K��� 6��|���
8��&�����ͫҢ���'�.��1�u	�=�˝p������iwӃ�X�l�H"�.�rL��-�.𳜱��X�Au�&�����߃�ߪ�o�.�aǛ�k�SI�,��q�kGN�
�Ja�q�k]m�Db�au�kZT
�"�K)Z��b�QEQQU��(�,W1L4��0U�E�kDiI�b�,��DIi ��"��I�9y(��0w�s��չμ���Whr��%,]�F��@�|�:��8�&��	����D�-�W�s��:{jt�L3Ԩq�����������'�6γ���t����i��:C.���u�~��SSlG�)}�9������2J�^�}Ɗw�|�qE ���R�Vm���!Xq���ԕ�^���*�v�)Y�)�H(�P�J�Sf}��z�a���a� �m8�(���R
Aa�a0�R�O
,钲m�'hT�Ȧ:�^�gκλaĕ ���$��R
AH,2¤���E ��- �e0�y�
Lc���:�/{06�������\�`a ��=L0�
�R
A@QH)��*J�Xa�f
AH(
)�ݛ�n�� ��,0� T���
����0�^'l0�AI� �i*Aa� �
A@QH)���d���Z����g(k�S��;y��8w�:��2��'��K&h�ڔ9�=T��u���W_��2�	$��6����!�H,���^�0�L+
²
�PRE!R+%H,2���:׽�H(J��T
ɶT0��E�0�ړ�T��E��� �h͘H,4�����Y�o<�J���R
��R
AaX{�AH,���*)!Ƥ���'��aP�J�P5lPXa��������@��H,4¤��PS ��H,2¾�*Ad�J�Agl� ��sz�ä�Èz� �`(
(t��N�f�VaR
IY�QC)*AH,�%H,0³���� ��
����� �`T���a �PP4�E �tʐR"ņXT���*C7�:��`(�"�XV ��=�2�R)
����d�AI��P:=�e��H/L
��a
�AI�=繻Χ��m@�V0� �JʐR���Sl�$=��A@Ǹ��� ��g�v�q�wԚa�
��ha �Q+�J�AH) �0�����H,9�$��aR]w��\�ĕ �c
�IX{݆6�R�T��Y���(���\0*A{C0�P�)0�Ĭ�����^[�[���pu�V�,Y�����,+��:��x��!��u7#����sg{�z�$O�	 ��V,:aR
NЩ �=jAd��Xe�H) ���Y����wy���yH)6�a�Ł�Rֽ0*AC�p�R
Ұ�$��R
AH,�� ��z�gPP!�@08�t�L�T��X�H.Cޓ��槩 ���Ji���e��1�[����ԇ�X��P}f������k]R�+*�f����w���k̜gq�(h�8T�����B�~�ʼ*��\8z|f޷}�~��o�a���M��/I�G��|�m+�ge�I��9������M@�%��>+n��#Y������_W�g}��P�����.I�*��a�x���a=k�k>x��<ه��x�+Ç�1HV
��Yr�.شD1���3Bnvuk���݊O�vp�{��$�2-�G��9b�NG|����9�3�)�z����{u�4�\-]����:��W ��c�faf��w,~����^�A��Le�:�VXiJ�)��X�6��K4|Gʐ�u�?����֨�=JF{F���ܲx֨��Yb_<�W8���ט�Gv�u=\Rqn��7��7�c��Qx*����˹7�`�4z.����\�S-�n��ɩ�6����Yb�����>�EE��݁����7�W%���xZ������`�Xl���$�T1�O�cڝ��WïՌ����=\
/oTp��Mՙo�A}�]�uKf�z/A��@0뷸�B���a�����W�۷�v�OTb���˱�Q|u���C��u���ĬJRk�b�4;�y��0�o��^��ČƩs@��WWj�T���eI!vD�e�NFNO��`o�w�ο�$�C�ףٌ�4��sy�{D�!��$9�*Ĩ��X}�q���k�������Dk	{�3�M��^�X��
RP̺:�3���M�pں��w$:�!�ه.�N�K�B	�gֈJ�j4�<��}��g١U��O �߱�v�s�i�\ȭ�=�A^�S~=����l�Z{�+5ϴw���3WyP��O��^Jfԉ���'^`
�[���Z�'�$}�V5[�𧣇F�dqx��ms�x��-x,�����s�7Y��{^�]*���N��mDM��v�F;��a�6��������f�������C7�]Sû%���^V!P��X���g\�v��I@�-�(f���Ox?��1�[KGK.}G�ja5�H�b]�K��;�7�ľ߾��\�՚��L�'�5c��b8��w.'�T�X�Q�@�fê�s�5E��i��W����U���r>��w�a81����n��@w��cN��3�'%nQ#�	�]��t)����=����� ]eRݭf������%�����҉�f�5�Y�h�����{)-�3B��CY4�%�#�"{����O��;��u}C��eY�Hr�ܷVri��(��G>Y.���>�9t�f늋вuihï
�G���ԯ�p�D�9�#"kAnՏ�f�_ep̝�֪,�Z��C,�f��[U�n1=o9��tu�x2�)�^�1�#�����̱(]�"�J���=���0�V�S�q��Y��k�]݃	�v�Oz�acf� ��B���ژ�����ű���m�w�7w.�R� �I�->����9�δ������/� .����N�f�����[S���M&����͔�Ѯm�*�E5J�=�҉C�q�e�oi�͓��N���⋒��Z�-�Q䮟�վ
�.X�!���'
�i���f�"-q��@nt�
0��{�I���޻|�5��LZ�wv��������}Z+�"�)qE���c���ZUQb�5�����Zֵ��k�-���kZ4X�iH�Zֵ����Ub�Qբ��-�q��*��j(���L5"���Q`�	��"�B�X۽ya��_e�F�AV�=0�?���]�Uv8N�l'P?X�Ov�雐���[�Q�y����d#r.��r�b�)Y[���%'k�,V-8(�qh���}��=L��k�N�4�D��2�-dZ���b;z�v�ܕ��/xo��cj�|N����bR�mq&H���}4/&.ڋ�U��4�po�{�_c��K�����uu��~�����c�����g-�zb���w;�������ӥsW�its�2<�sS����BɬKG�0��xw�h�c��x�����s�w�������/^MT�Y4�l�3��Yt��R{��\��?>��t<X}��z�KdC�n��s:�,Z�J�E�����_���>��f>������)��3a��Q���xe��=�b��z$�]�+����Fh��w�2]P����ޞs�t��m�8:t^$��s�ə[|�<��[m���;�;P�M�Z7�y%���~g-���v5Nk���������0��k=��N���ܕ��V"��pI۵$nu�E���]s�s��	I����g�9��u䝡�������zj��mA<*��4�& W�@^윝{� 9E��)h������ʽ׎:{k�w��:��N��{���ysFG���׮Cc��}�����灴w2��6�6����!m�s ��ct#��ɭ����?C� �)!!߾y���Rߌ���z�ֲ�?���s9��| �/�u���V�A#��qC���ԕ�z��#�A�yJ̽[���a�#��W�I˂{
�����<�s"y��:�^�y�V���-ͨ.�Nue7m�=z3M4!��̱���F���h^��i�7�|B|2E���9�o�����Wx�nb�����`U	�;`��T�7��<��V���ש�~{��Lc.nGU�NvW�25��s����9F����|���:��xVY߽� ��j���=ơ��������02:ֶיu��KO�ˑGFO���ia�rPs�Q����_�~�	 ,�R L�y�<��:{���2������*�in�{����5h�J�%�''����>��]d�soo�+��{H�yV����k�.*��C�k�;�r�8�c�|Wﬀ�[垸�FX�Y��m�2�a'��lm�ޝ��,�|�R��خ�粲�-Gr>O� �� ���;~9���:|u�yN�Ài}Y��7��>�΅Z4,����.uZ�l��z�u�� �����~3�����xo�@yp��w���Ŝ��5x��"f���aۅ��c U^R�Ǭ�_x�j��-��9ݕ�k���=s�����9��`
 ��G�	���ח��տ��dܭ��1q���QG�o��e�\�����@�g��&��qOp�]��w뮴�K�N��\w��`hWT4�g-�;ү�$���ќ�NY}\ѿh�5��3�E�u�W����H��S���ֆ�W-�筻��:�w��g���|>�H���}.[W��*����}1���98Rz�� �q?��<k�w/8V�_`S�h�j%�y~��w��.RjYt*�>�����ي�K�M#�ę/�ѧ���H��yK�
��U| ����=!����^�]b�٢���{͔�*R��f�b��Fb�۔"���Pv�A�R�J�H�5&�dG�
�3�*�-�[(�w��mY�h�A�\̧�P��i+�';F���(ް/{tF%P�sr�E��Yn<*h�� ��C��ô��Z�Ҿ�]�xS�艩�N�_��Ov�gEދ�s!s���H��Ʉ�¤��o����-����&fM���V9Xҷ#�7kz�S(v!�m��)�Z�_ ��T��!6���)=��%6,���uȌ�Y�I���N�]�[�6���e����8�b��rۨ7:6��V$�2F��I��U�I4z��B-��a���A��8[��F��f������S�a��5t��٥|;Q����{�������>e��DP\�'��z:X� �V��5�k�0V.���gB"�V�ZPWWֵ�D�0T�b �Uij�5(�T��YZ5(�Qhأib�
�����T��(��+[hVȰ[Z	h(�b�V��*+A�5~�Y�;��|#2�N��W�ǟ����N���e�r]\�/�������f>�f>�韢""�3ȧ�G�l����Z��GCʣ[u�2cG4�ҹnyΛiZ��s�	�������g~�0f�i�r'������ĕ�#آ�@�}����i��IC�\f�ݢ�W/��9��N]w����}W���~�*.�^
X�{ͫe�Մ�j��dt�y/��$�t m��ԝ�)����y��߀�N��g��]��}h�m%��bë����1���Z�:�U�@Y����2Ou^������7�U�S{�yೱ�v��~�p����Ԅ<�-��Y��5ڦ�!P�-��o�(D�Nh�q���zV!�q��'�q�����씆ZS&]�7�|9�wψ�H� R <�y�����G<??^ڊ�y�$\K�Z7^�ȡ����Ǝe����ы�;��:�%ٳ#�0%k٭���6���>�贞dҬ���y�g��Ǭ�z���,V�j6��4��<�e櫸Ӎ�{aE�G��"�]ª1̾�$�L�7�_1�o�4=s�������	�`G�[}߮�?]ف��o�A����87�w�h�]WKִc��5ԏ?qdg�&]D72�s�����vR�?�ʨS�\�O�����e�0��~��m>5��u	Nhy�F�� �����`%`WN"fҷ�=��1Eh��I*�Z�.��:��Ùc���"5cK.P��v�rW��(
B)�Ϟy�Ϗ����k��߳���A>���ʪ������_�%�'{��`��鹉�Y���F��6)�"�s�� 7WC-�.E�Ni�=+^�����N�#���v:�wbۧE�]��l��5��7ી,A�ȸ��>���!7�S����~Z[���;�>D'�$P������_�u�"��O&n���T�4�(~G�s�yt#&�ՆƆ�LB����eP��<�EMʾ��ĴseŇ]���a9��"~��K6�X�u�It����:2�m?te���^���P^O�6���{ebጔ�ah��*�ȼ�n�FS��]s���X�;�>@|�
)"����~x+�!ȃ~WGF��^�T���@ʊ��P��.�+j��v��{��>�r�7�P���Xؽ��_�P5᫼}y��J��g��!��G���;�[F��&o�g]ж0g�@�����^��ή+[*q�	~��6����H}�����c9eLl�6�aa��I�~������H�
@���5��g���'nq{�:���������Y�I�]��R�|��T�]��w��O	��?�߮�����=팕	ϫ�Hb�ַ}@ܑ)�����_oj�ߗ5����L�����Gg��-	m)w�#���o	�}�{W���<�6w7y�LP=��6dgcRmQ�$P$Y �Ǿ���מuq�.��4;��]���|_B��S��1���o�K�鱤�M�uۊzn��U4�wo�u7vrc���W)\J��)�hv�^�fښ�O����н�X%ߚ�G���R��Z��ʄ�pb��j�̼f��K�I���h���r�F�n B��>��o��|޻�7��"Ȱ�$�9����O��Wn�����q��O+k�/���`xx��|�Zz��G|�	���\�W�X�̩ܫu�ˈ4�e��ΞC�����Q��k�l��3s�0���)�U�C~�7� �W;��K&j'�����u>�wY=5;�XʹG!�����V��z.���^7']�
�$���68f��a����f�(gV�зP�N �^�2�:Ê�e�M52�u��Y���@M�\rҬoT��u�y�R)�?j�����H��0^n�H��c���@�]eDGVfŭv�'h��y��j�;ٳ����x��s釣5�Y:ja�a����5�_b!�������As6�Lu����N�[�g�{o����%��#DY�r�u.uٹ{�Qt�̚P�J)	�%nR�˵T��Z\E��a+��x����ܱ��5r]M�6ٌ\�1��kr��"�%w���rj�b�����F/1?�9��wZ��ƭ8;�`��|e���L@{�ш�Q6[��Y�,�@ >
"��#"8Ƽ�Z�ե�F�Z��[�kZƵ--�Qe�����k�kj,cF���kF��T�R��U)R��m)D*T���Tm�T)l�ƥKkj��kie��V%�
�EE��j�m*���Q�[mJZ�Z��m-����[jJ��M�4>���~_�=6���2-^�2�w�R�^�"ff&~��x�e�g�Σ�\V����;|����W<<�#�{�����@�}����SD��K��!���`�ԵB�x�������7]�\<�%��-�ט��Zk1�YMF@_�I���`�)���֏U�JB(�6�V�2��M�P�(h$���;yP���������}�<�|���@X)$9���̀���Og�G���%��Og�Qo��[_}�|��ֱ�ጀ<��xJo��-��H��'����c��g6@���{�0>�-�.ъ�f	�Ǘ�n��Ն�dgv����71>�]N��5�~�0t����i���p�wwH����� ���v#��i�+����]~�"���y�Xu����]�<����.s��V�P���x:c�;طy;w]�y�{L���/�g�T71\`�F��t��T9�fa���/����E��Gӯ.���S��˺f.��R/��g@����W�u�26�(�n��^W>���h?V7Ve���܆�(�^=%J���HL�VR<��?���wW��{��5�����d߰�"fM�y����'�K�λ%��3$+Lj��6�3T�TQ��@����n{O�������@��W�+�t�3AU�Sj�K{�8��E���T����dB� 8U�{�{jq�|/y�\z��dK��6(����
ZP�HGb� ��.��6�q���wWS1��d=t�?����6����ޜ����q�VTv9֌���P��\��������ܚ�������$D�h�po7���w�G��Z���a�.��H3_�I"��ژBKo�nv��yBKtl�0$V��iݹ���K;��?f�5�zWb�.{2��w"��>,���9�ݝ�k<��)��?��tST!`���1e~&��Vt|a�ݼ��e7Nr��Ր#�o7,e�{ֺ�n5Y��扽q*�7�9X�L��v��=G���c-���?7�:�&r��Č��X����[���Mm�"��8�sܸ���g�(�	-�:���}���>$�� (�)'�yǗ��P��V��\��*�(�S`���q��n���]]��K��;F`���5=
fw
���j1��)���f�tl����~W�M��x�/���$��g��}�zH��.{��3;�t>�D)�;�h���:��æ��iOwa��p��+'<܍��c8��m����ӱ�:�{�|˾��|��,�Y!9�hA��:�M~4����3KUx�5��-fWU4�k��x\�{N�N�S�O�Nx(��܂��É��ʃ-�Oj�j�1sCS�S�Z)�`�۰��*ϼ;���X��u�Ӂ�vvN}�4K^f���=Օ��J���ó��]�]�3%3����}n�k�����s��dP���J��gPj����򍛁�:)s��V��uT�1f�K��x�Y����[�Ӥ':5�!�Q��4^7�X�1�\��PUs5V�����y�5��$}���q4S�q~?O��]K�{>��s"0K�fl��F#7�O�J��>�6�$��I�$̔#-���\��E$X9�<��-���g��y����ή�2�حݔ(g{�{eh������V[����K|_��'g75��fþz��_U���@��-���F9�/2"�3��*x>���\��-�G�+��%�mcp��!BE��]�*%<��;��S|ldܦh`=��W�����tH���`{,����u���ƒw�q��ȤY:�[��#��K�N���ZbSg3eq���T�"6~\�e� Ȼ)�Ua/��.�u��f���Ѣ�ط��W8j���e�E4�q�����9ԮP�n��Y�7%)�+[|"�E�='nruGz�;o9�Q�EL��T��{�v��ӥ̎�U���U=7�]��$���N�'�v�5l��L�^Z�t��Lw��If�4��GfA�8y��� �k�u-&��������p�P�6�Ʊ̝ݶ�c'd��|�d�3T�B*
���a�cZ�B�_Iׯ���l�ԋ�<�}Sat���+�W]�*ֺW/�گ�#�R��w^%�gջb�Z]�TEZ��B�b(���mV�o��t��"�T���QeJŕ*�U��Z֤�X������j
#n��u�heF���֖���X�kZΦ�ԥkX���B�����A��ib��6�m,mV�-m�E��A���FЪ�
�X5J�j����j��-�����ֶ҅��aD*���F؊2�hQe���clO�PI"�Q�X=�_��di���dr����e-SfY�R�.��_]U]�껪�wUU�9:a����`֌lν����T ʘ�׻C��`>g#�+ٿK����f�����֎W˻�0��dԞ�޹�c�Z��gXʗW�F�#7�]�D�g7y�rK����IU�^yj�}�Os�z�W�3X+�J/j0b[D��7����\7bC;��I~��3�L�����]��ƄGW�)M�����団�z���]{&�OT?�S�v���w�a���~�b�	���^�8��O��solk/2���gN��O�y���Fbs᝞�C��c~��>���2̂������C�y�{��Oaz���hmΝ��ff'﹤�w�U����Xk�暠ᖹ(��T��;V�ڋ`Ac�(Q��ٝO4vxkc�i�Qc�^]9�jw�Y����]xw�:}�U���ƨ1F�[�c��T��:�5�7�NJ��n3W�/>]�<�����['<�P����mV��M�?'�]��&�o:�s�<����x����]��G��C��B�J6���������K�����8�;�e��j��v�v����*XyyUɬ�f�ىť�a���5U8�����˙���wBxz'`�y�[��ᮂ�ڥ4_���U��)�[�_��ʱ~��VHl�3�9�!
�<���<ـ��-�o9E'�N�����E�%L�|�U#�>o�����b[�&���C���Em�L���`7���� �����<��O����|BgC�fN�^j[�tn�����LB���T�γco���KxΖ�.��K�x`[B'����\9�y-���,�����eYa�*I�3{�/٠���|�G?�t}F��
��ϓ���u<�^�x���/4��"Eݭ���}�z��h����oS�`�3���d�	�uC5&��Nލt���.-N�3=-��ǔ�t����nʩ�ݴf�i��:ҥ������X�ˁ�6�ۗz�j�&.�/1���j�fFv8��QF�/;spm�X���)��^�!�>����A�FdEǸ�}26@}ۛe{a�s��p&;ο�<oػ+=|E��Z��.�+I�BM�⌛[:�^�y��Y��;�S4ݼ�o��*�Š)�4N�V���upu����]�K������%�^�r6�r}T�,�6���N�����y�)N�5
���U�u��%���0�FPė�2[>�n(�헸[ᘜ����c4wo/{��1��`��uoBz�b��o0��Ay�t{��νyyW�����^fb����2)0�Y�K6�[�<��:��I���a�� �~�[qܑϪ�RlV����O���γ��W+�����^��M}�����|�/���wk�eCl��/_������H�[:����u�>$���%�B�� �)�}�PwA�T}�r�{۽bWn�UA�-��S����p+��4/χ��1��_����T�eL����v�F;��a��������˫=ߌ޹����I�1�������`��� �vY��7�w�E����7�v�1�36�4r]QԷ�*,�G�T�>#J�b�u��>�<�k��� Mu�D8˲�K �����=
)n�o�^)wx�Շxt��[��i0�\�@�r*�cwr�
����ɱ#՘��6���u�\
�/�i��~�,,QmMh�I�K��rrЎ�ڝ��o#ڵj죄�^@�&�0Q�����I���]��  �/;�Ԙ2��!}N�&U���DŴ��xAIⰺX'��@������4�}mV.���J02��v5��+���W4f_s\�54y�4���U+3C�s�B3��������eH����%�ߍ���$�NS�%�'�6J����k͡��Cʷ2������.5��w_
�3I'F���$Bg�l��E����y���"�G.I���f���\�6&���/t�\�ۚ��Rv2���Uy�V���+_VH]72��3�+�ܪa�1���V�8�Q%c7���	��D��GĒE
��T��㮻օD5j��Z��R�im�Z։֊T������V�n��kK�iJڊ��KV���ҕ��Z�t��+kkJ)YQ���*���EQZ���F�PB�ZZ��(��TlkPm��R�UB�[QD�6���Im�*Z[h�Q-Z�[*�q�s�3�[גӽ��mEfI=U���P� `�V�4�TL�VJ	�c�g˘ڑ�c��ڪ,�����T5��t%�W�P]$:5a�����ֻ��#�3�0�{Y�`wҎͮB�=��7@�
�{�Q��&a6r�����Ӛk�H���gTޭ��F���v)3L�m��N���d�GR����N�Y�f�T��Ê���	���p"����ގ�a@N��A3��{�~��U���<�1�;���OyK2��fۦ� :}�aӻ]ao���i�]�����"�;�������咼)޽����wW8�61܀/���6��n_c��Z���i���ޜӛ{�^�Q�Nje�v�����Z�`��H}.�
��/�{,���5Z�շ�ɞ/�=�sդ��Э��
9�{mоs�-�2�����.xI~�tF����V[Q�N�r�I�X� kM���E�z�x��o�8j$d��'2���� ��t�j;�ȊZ�npr7�B7,Lz���ˉ�pz�Ԝ���r�7!��;��Z{zw�FU�]f{c9�̋�n��~yy�/kmSh��;%�&���E�VU����e�璚_8l��!���	��w���Q�7���h��Ζ��$��B�Mq�Nэ��[��~ҌȴEluT�� V��^,�h<=����lz�����2�^�ũ�0Q��離~x�p�+��[s*)��<5�USH�,��n��A*Ԯw��t.=�,H�xp�m�?2�+�F�W���zW�В�9g5�]Eh
���o��ctE�jr[�!���כΫ��d��q�\���y�Z�nW����3�k��{�z�i�H���V�����W_�y�dB�mx�^��t',N[�b)�3�2q� ��m!ϛ�ͬ�ì�[t}�ͣ��F%;#u�Ö�OΑG
9���(�R�U�܏qb(�����f��_��ƷǷK�ݼ�1w�����+���Jit:UmR�n��s`ynxs�վ{ǘ-=��1{-b��I�~���ǤS��q&�\�k���u�뜭�~>yb�5��\Uk�EG��f�]G����^�{|)�eL�!�h�*N<K�.�5"��i�v�}�OGY��)j���0�4�R7����:������?�%*�{Ge�s�K\�S`��V�C~ ���C���ډ���n��˭���2��¼��mp�ٛ�wi��yfh�hvEW�f�֋�n�u���,(G���]���g^�z���-Gr%�X8��%vמoTͻ��)Q�.�\t���c/��8��a��X�Vøb�v+��<f�U�j�됞�#�B�)�7��w-qi��A�fF�X��ź�C�s{��қ׀Xu�#���ڶ��8�AH�ȩ���c�'IBU�n$d���A����w|�t/T�j�.c8�{Xt�>E1Ie�
��{��&"k��L��5��{�?z��W��77 �̸�nK?�"��L���{�|��uա��î!�[z�n� �\z���o!lYX{F��LB�w��=�Я�d�����p�N��؈'{��j(�2�u���E�t=�:պxiQ�������������e�_�8�-i�����R*���V��r��dT��tN��?]*
�cN '!gt眙���E���R�Wå'��=���M.���{MlxQR�i�����j�oJ�4]�j>36���kq��Gu۶I��v�\�`_\�����IPm1a���{k�m��]d=��C�n9���u�={��e;� ژ�HUu;\�#�vr���/�ᱤ�
��h\ؕ�-[j]�9�vP8ZzS�pnXB�BbQ'I��%���L}Rr�,�ܾى�����p�+�Æv���ZYGht�E��s�s��� j7՜��_�jѣs.��U���d�+���Ӎ��j�ƋB��6�Z�����<�SQ�["�A�*�in��hЦ��Jڥj5m�ֵ�j�VKjTe)F�kZ�ѡFԭm���[[F�[DV(��X�ڈQB����[j%��e��V�J�T[Z��cY[H��+A���ux�j������cwP��r��sF��
o6�w'!��o/������6����q���p� ��X��7֔X��W����^��\N��Ӓ?�|\�_�I.�ݑ?rU���)�5�u�6N��{�k匧m����$3���f��j��x�F�ʻGf���+-ړ��vO���c7��̘��u�2�^���7#�������z�۹ō�K%�%9��������0��RU݋��#0�H���u���77�u����w�uv���5�NnMRs�sTapUΌdu�|LT�4��3�|^���`)#>�w^�<B�h�Ys�K��`^�z?]i��yv�J��M�cx;w�V�Ι/��$�t m����#�np[��eh���_�.ڛ�E�Me^�M�Վ��O���׷�����ӟ��=��՜=C>���K��Ԋ�η��<�����Z�B՝�����;#Li]�<�
5��}�ܗź.QV�+�,O�;Ǳ`�w���
���t�\N�U�R��$�"�����S> I⧉a?+�9w ͙��?b]r%xg=K1Y���4gSKrv�j���{���j%�՘�/u�I�#��ϯ���n���tݛ�j����Ј��6O������h]�r;ݭ�����vL�W���̮5���J��m�9�����!���\܆�y�V&��v��]�����7+*y4���E�h^շ^�)\Hz�Q�E�ߋƏ�`���{]WJ�{���^�Wi�^VSc]�{Soiiev	�0�P���ȻyW��i�>�o'%L�T05�@�����mE�%�����jli�?����ڄ���{`u��G	]�,�g���Ȋ��:��k:D�ȷ�92�í�]�?^�j��9��JӦ=����η���܊@M��*�vuX��f��{yd���U w]�Ƽ���<��?[�B�vd�^;��>��:���E��j�_y���CDѾ�ۯ?Q��qaf�]��!��"܏N;i��o�u���܃����t�������8���aV��q�v�Xyv� ��V9��ч���,�kEC~(��/5����-�2axm�'d�KoU_R;��=�'����;.wq�y����
�\��:��$|�"���{�N�m���1��̉��E"l��>t
�#r`�^e�$��}�dTT�Xy�3���Ҟ�����z���5�q �v��x�v��]��񊵴�z�`=�{Y>wϨ9�Fkf���9�P��Գ�Ê��/�Oz�O?o9n�c�@�Sꃝ{`꒯@(���cD<���WU�ցC����e�*Iv�;�	�k��y}��
+.g^5��4�Zi���̳�s���|ݯ��v��)��[7U3����S���˪��u���}g����T�>�h/
9������O=1L������v9�O\���
����}���ˋ,f��?R齕��c#�t�ٸ�{Xn(�C$e�;�;g{y��(�$������A�\pRÒs/ޯs���=FFP��Q���������N�(��1S�Q����Z�P�^����F�Ǧߦ+�����E���8�e�����o�Mcb�8��G*�\�ř��v��S�����$&��r�y����jİ3��� �fՓ���կ �����.���P�^Gf��Ӝ�����g�0:[���:�Z�k�v���*�ЛOX�)��:�6mjż~���=e]��Q8$�ۓ�EjD3�Q:껷���EЈ�l[L�7��\�ޛ�)4y��u-�H-�n�f}�ȣ��o��PO��R��]u�uIu�ke�4˝kMow:
�����#1�h�'Kz��]�.'�d��.Y��\Y�fK�+v#��=����U��ssY!��`�A��Csm^"b�JG�����a@.fa�sf���PG$첳6d�
[��ֱ�+;%�����h�Ю�4_
��]���>�6b�� �P PEk+V�}�{�ZT�h��R���kZ�kTF�����kZִ-��kh�kKh�kZ��t�iKj[K*V[h�Q1i�V��ث�L[-��JZ�U��0�)Q��n-�V+Z֥�A�6�V�h�[p�p���e���TUE��百��No�u��(��׮H�*F�fg߶��s��q�h3Moҏ��	�yt<���.״���{B��D[��&�.o��J�:���
,�lC6lYgUK�p�`�]�8'����=���8�&�;�F�s�Ȗ��w��n�m������˚Ҟ��ǖ�>d�w&��
=��{@�KV��Yh�����ă�z��۪}�z���`�
�^�$E�k���u�q�|����X㷸�g<���wyb7FMH��f���w����
��͙�^q���"3
t��y��{0v(MC$��;]: �<�����;��I��ڀ�`�n/��X�/9 �"��F���y(�X�e��DE&U�7DkG}�6�^]���mM��֥o���ok?�e,�<x���+�k��Ge�(�W��s=Wb�Y�}�:(���>��R-�b��Z���i�{Zx^��A����*a+B{w��a�9s%�=Y�~e��b���o{?y��+��=8��vKn�u��5ҹ�]��k��*X��o}%��SQ]�/���~��t�9�w��ϧ;�j��V����M|���?�T�Ѽ����y|V��ڛOnj9�V�<�i�r-�,�e�Z-�uMq��	�uo�������I*�M���'RY(:u�\�K�V[R<q�ݞ����_�-�ˌD�j'1�3����Ԕr$v��'g�I��H����k!͢뒨�Z�xs�ʭ����f�h���H�([]��ۑ�6�1�p@�+5�r�x���{w�z��)���޾���$7�T��/+y�2��_a�$nmw%9��=L�w��7!�ǅ׭_fԆ�\�=Z�'ݵ�a�=��w�{pn���k��}���8;Qz!���mC�y{��eD�����1{:7�������&j:��g�v<�y��'��<���.\�o,4p��z)�W�[Jy��-�N����_KX�=�n�U�`�H=���j;��?\�پS�Tڰ������������w�9�0���a�~�����T��C6w��1�c�7��QYP[z�����<Ng)d�`0���~�r7nU�Ic�����y�L�ԓ��. n9��$�CǪ�Vޛ��(���(�T��3��Ҷ�u�N�"�(J�#i�u%��������;��0`,4h�x�����)�cܘonK���ћ����/��1O��;�'sI�{�ݴq;(�;j���#'&,�����j�*���V�-���]<tyz��_�}�2�"{�*uv���tߺ���u���4:����寂'm�Xٜö����5+�r~��3��٪�?���{�*q�t������
�°vS���-�]�'��h�����:l.径_�;�.?b/j��M��7b�n�7v�|�� �4d�e���<ѮC��l��?'|:��;��hу�z�%}P�d�w��n�S%�OwU�
G<��Cd"y?M������̯_��F�U�4-�t��d���L"��OAJ����.B�i����^p0��n4J��@ڶ�[	�z�w�gU!K�~7C�_��s?D3�OZ��qY�r�'!θm�E�����y���s��owMϚ�3���0�����'�~��}�
�EQb���J@� J~��$��������!  |C6�,�?�L`�b�S�L�x>G�M@a��������\��f���0	㤓9
@`��
IJIhu�%�I��$�,��g�Йp0C"ѳ�I�$��!$#B�$�$`-�KB�(("
�PD�,AAPa�("
�YAAAA�(("
� ��AA���G�	0��J���l��,�S���a�R��P:��JM�p���O���� � Y1P�|���7龾]~���|��>�`:�A�/ぉf���?�~�f}��0tXp̆v��y36ц�ae:0l)k�Q���'�JY�a������؇�\�B������?��������@
I������  ��s$�� PYHRL�	���^���������	��?�u'�0�)��I�?O��u�>p� ���B��d?����p~BDbC���L�����N�4�s(��O�@:H�,?�{!����c'�'�������1�<�k�?i����+'w��?�	�4DԳ��i��E� p��,�'hh��c�I_�g�3(��d�)� c��L��=�k$&Y$��ob�E�^�f%��l%�\_������?�D>t��'��G��� �!B(�hBB�HT$-h0�!��>����!��|:�>�����HC$.����圁�}a��I�>b2���>�?Ϡ
]���4d?C��?��O�q{��5��1>E"K B��%�0C��'���H�&���������fB��O�5���!�ؐ�7$?��E����}���G�>�:?A� �|=�O�����gg����3�!����I�~�����g�"?�z|uf��6?�%�����B�JP���$��X~ ��!���Ѓ���O�(-!��!����@�2I��S���� �4B8M�,���&@�n�	>�(����C2�)��H�����&�!$��I:(�>�}���h�O��S�= �C���?ҁ�@� >;	�d:�1�g� Ɇ,'��t)��x�@�! aO����΃����l'�$�d��� ��$Cߤ��RC��}& 3�O����>g������y> ��d� �	��C �?X}�|���?$C ���>ट���O�!�� ��$��b}BO���'��	�3?��,� y���tk�}g�% Y +������C��d�! ���@���78d��?W���?T?��}��}�����}d��LY�?yߒ����r1��3�� Q���ϟ��/��2}BCf��0?O��|�$;����%��>_%�����{�����_`'\�����,ܒ 	���'�	�k��Q0}��|��}V~&�"C���Q>��>s�|�=O�I��
m��4`��́��'�I���0|��I @�!C��O�C ~��C��	�	�����O?���� ��?T��&C����i5���@?˒����0C�1��?\7���������3�$�/�����w$S�	O=�