BZh91AY&SY��`�W_�`q���#� ����bE/�                  �������H�2eS���+jڒZ��k2kT�SMX��,�f�j�*�����)��U��Rhj�*P�D��v��5fj�h�ؚ��H҃*�m�͚T&�ښԐ�V�m��SL�KKL�lR�lƄlh
w��/�R���k+U� 8�.�Dn ����Tի� ��Z�)R� ,�cMfKQ��V��f��mf��F�j�٣B�h�(T�[g{�� ^�ԥ��
P@ '�R�  +��"����m*;*�+�h���mz���kZ,�����#omqFm�c�t�jޘ�-hw_o}c�R%����t�Z_s	km��Z��e��_>�I  {���+��+����=Q"]Uonݓ�z:=��t����� ^u�z�z�WkvB�[����m@�ݫ�z���]��{mhi��载uJ{�sjʙB�UX�dA��I( <;۠]O�����{�@�խ}���}�髰7�3{y��R���<{��[��Z=�=�޾�U ��=y�E=n�t�<��^�CE�}��|�>��w� {�^�Q��ma�-T��T2�>RH� ���޴����[W5�t� (x�{x����7��v���[]��
v�S;���4P�]��ݽ�
����3�q�En�f��U���T����w��Sw�[6����a���e�>I$� q] ;��@}��ꪊ
=OyΔ�
�ǯx�C�����w�[lon�G|���K��/��:��'�נҩE�����Uր�{o
UR�[��0��M66�mbf���%$ ;��� ���΀=ׯ �ڽ������zs���$7c��5n��e�Z�g�(�Op �z�Y�6�iFU�m3��IH ���> 3N� ��x��^Ǹ���W(C9��ѯawBj�v� =�^^ �Z��� �yU�I�d%kS6ƶ���JH�>  λ��;u��:�� h��� ^��� �����
��Ǡzz6��� ����;�L��V�2�ͬ�V S_|�R x9����5)�� ti�w� �����-���6�ݠ 5�{����q��7z����t=<w[YD��h�ͶU���I 7> ���@ϻﷻ� �k[��� C�� �]�w�vi` =��o��(m}�h}%@  �  Ah    �JR�i�@0CC@2�S����CCFF�14�i��4�� ����h��   ���ST�`4� i��JBeU&�h� h  �j��RJ@M�zh������ڙD����o�?o��?o��/�e�~���1O��Ȧ�׭X�|�u��9ן� �����U^ 
���_�� _�4��3���?����O�W�0��T����U U���I$��T_���`~JAD肨�/������`ɋ�/� �`� ��b� ��#X��5��]`�X:��u�5��]b� ��u��q���x���5��]`�X:�F	�]`�X����u��#X����u��]`�X:�kX�bkX�5��]f0u��^0u��bkX:��.�u��g�1��M`�X����u��X����u��X:��.�1�Xc0bb�X:��.�u�k�X���&�`�X�5��c�:��.�5��]bkX��5��]b��k0u��]bkX����5��Lf�5��&�u��bkX���`�X����u��`�X���q��bkX:��&�u���&�x���u��bkX���1��u��]`kX:��.�u���.�x��.�5��]bk��.�X���]b�X���.�x�bcX:���u��]b�`F�]`� ��b�X:����u��`�X��5��f�u�q��X:�5��]f0u��^1u��X���.�u��Mc:�5�kX��5�k�5�c ��b� ��]`�X��:���u��]b� �.�M`�1�.�u��]b� �.�u�bkX�u�`� �.�u��#X��5��]b�X<f�b� �	�X��5��x���`�5��]bF��.�bk ��u��]f0u��^0u��]`�X��u��]b�X��5��]a�M`��X��5��]`�X���.�u��`�X:��`�X:��.�`���X1��]`���]`��u��b�X���&�u��k���.�u��M`��&�0u��]`�X:��&�u��]bkXF�u��`�X:�5���X����u��]bkX����\bkX:���u��]b����b�X���.�5��g:��.�u��]`�X:����b�X���&�`�рk�.�u��Mb�Xk1u��]`�X����b�\b�X���&�u��b��u��]b�X��`�X�����.�u��X:�5��X���.�u��]`�X:��:����u��]b�X����#`�X���.�5���bk ��u��]`�X:�1�.�u��X���&�`F�u��X��5�kX:�5�X�0`��u�q��q�k �.�u��5�k�]b� ��u�kX1��u��X:��.�u���b��.�u�k�.�5�b�X���.�u��5�k�b� ��`k ���b�X:���u��X���u�k ��]`� ��5���M`�X����u��# �&�bk �.�u��X1����u��M`�X���cX:��X:���u��]`�`F&�u��`�`kX�b����u��X:���u��Lc�CX'��u��b����u��]`�X���F�X:���u��]b��X:���u��]`��$a�`�X����u��M`��5��M`�X:��.�u���$`kX:��&�u��Mc�cX����5��`�X:�׎�1��M`�X��X:��X���&�u��`�X:��F&�u��]`�X:���5��8��.0u��M`�5��]bkX�b�X<`�X:��.�u��5��0`�X�u��CY�&�q�kX���.�u��1�.1u�kX�bFk �.�u�k �.�b�#X��b� �!�CY�	��`��5�k ����0b�X���!�]`q��q�`�X����]b� ��b�.�1u��X�u��8���/:���b� �.�qu�cX�u��]b�bkX��5�k�.�u��5�k � ��u��X���`� �.�u��b� ���X8���]`�5��\f�u���]b���M`�k�XcX��8��.�1��u���]`��!�c`���u�k ��a:��.�u��`�5���]b� �.�u��X�����]b�X����`�5�15�k�X��5�k`�.�b�5�k �15�k���P�\Ax��`���E�"��#M`��b kX��@�X�X��]`�� b#�Tu�.�E�":�WX+�u�.�E�
:�X��]b��Uu��5�&�B1A�
:�WX��]b#�Tb k��5レL`�X:���5��c�#X����5��`�X:���5��a�]b�]`�X�1�.�u��`�X����c�:���u��Mb�X�u���`�X��u�k�!�5���5��]b�X:��.�5�1��x��.�`�X��5����:���u��]b�X�u��]`� �!�]b��!�]b��1��X����]`����]b� ��u��X��X��X:�5��X���5��X���.�u��]`�X:��kX���.�u��]`����]b� ��b� ��d`� �.�u��X��5�k#X��u��cX��?Ә��#������_�����0�b��������_K�WI;۬�N9�-�M+2[Sm�˶�۞�nʧf�@�A�1mh���.�+A�X�ܻ� WG��(<1�(pc0֩mJ�擑mZ�0뢣ɇ"zbec�{H݌�4���p��VFl�kn��d�	;���)�fU�u�:t�hͼ7M�ԣ�1�ᒪc�W��d��-P,0���Rl	p\n��(AՑ)uk,?�H],�������Q���������U�q�,�n��3IثF�0�x�N�Y�J,H�Y�5�ÎJ����V���i9�$��s��&�&�����Kw&PgL�v�El��抎f�2�`�N���1r��Nm�������a2����'HB�Yf�W�Z��,�����bjj��_�'u3n���*��Z/i�f�; �z�n����.dnR�"��,��{Z�e���H��ʗ�%���˒��&�M��a�*���җ�n�ypB��9��`71a4Xۊ���x���#U��ѳ{+2�Q�b��AߍҳOe�ă\�[1&ȵ�c�ռsl�f�xT�U���U5��ڭW����*�׍���D^a4Dۇ\*�2���}��ɘv;+3�A��^B�Oa�R3[a�]�ݚ1D���\c.����+]���sSy�U̡Sm��,��m:t�(#��r�R7q�U�8��yo���G8���xkG�����II�c���FZ��Ke��/tFѲ��e�ě�j����14(��w�x�n%7Q����,R�r�
���i:&��w�p'��	��v潸/(��7*����D��f<5X�уCxr+��1q�m�1���f�]�;��q6.����Sײ�Bo2�R�v���YH�����&�/v`D^�wsp�ڹvt-��F%J�Y4<���.U��ι��kI��7�7BSr��2Ru�[ia��I��N��zR���R��~��.�R��r,��<î0m:�.f����`l�j@�0S���mZXx��]eZ��k�j5r�㪵m����sR�z�/]3H�­3N	Q+�t�Xy�V�T��%�וU,�z]6��n�w�D����#�V�.�)m�ܧ-�T�wpI@�ۦ��,��Q��Z7�o#��L��S\��1Ul�On����t���){�J���K��-NëPߡ��C-��cR�z6�d+q�nF�7O
���IW����w1��I6nM�مǶ�!��읨&��)62U7/3PX�̍�a)cF��Zؤ�út��,�z�KJ�wYN��i�Ǻ4�2�"B��
v�"8դ�x(SF�T���om�eb�w��c�͸ql~.F-T�I `'�e�L1f�����V�)�֊uZ\��%�6�4w-���mҨB��F�N:U5�j�4^U�{� �X�L���x�,���"5F�Ǒi��[3^�z�<X��um��l����͍h���޺�R�)��6�L��h];�y7f[,�K
U�%G�'��̔�'���u���U���TFPK��+E��Yf�nB�k��~�Iʭ��sM�1-�i���$�J�LИ��%u��ra+wcN����0=��h��$��ڂЍ����۫�;��i\B
��$�ѡ�kj�ּ{b�9.
l���.��ܗ4Pw��2��Ex�f(���pGk_�8ibn4T7I�{q$,�y��4�i)v��U��%1�ԅLg}E��e���M�j�
��1�LG\ڂ�g(��ì&HJZwP���<��u5��m���K���[HY)��j�B��L�rj�� r�r�%y��ʐ�[2���;wMhr�I=WnPå��`�d��ӫ�b�7���$��QG��j��[IS�aj�U�� ��}��t$:�4�Uf�&��Y``��]���n����nV�����c.��KE�&��/d�{X�G�m�ʱf����\�b�
���
]i諬Fd�r�B�^H`�
�vm
#��6`��Pnջ�֬e�qٌ�r�ȓ����)�\(���J�i�\n�aʘ��N���6=tt:�.�bi�N��q�+ǐɗt���j�:ɭ��,-�T�݉��U&ɬ�.2�n�8�+�RY�)	��M���pG��X����unF�����M�72�N����1��c{3�V�f�-7�3e��J��V�q�Aˑl�jf�-�&�]�C�dۍ��D�k��[�a���31Z�Ԛ���B��Z1�ȋnmQjVi�e��N���z.{))�,�K]�=��ˊ��uZ[�E���SN�m��9��Kj�zQ6ubI�m1��ʽ�x��:��J�U]ܤ��ɬ\%�l��T�f)r޴#aP:ow��u�B-'���E;׋��!<��~;!�q��H�wGD̤��t���Z
���K�W�J��w��{rB�[G]�Kc���N��i6�4DW5OJ)�si�y�ם�y�;T��OeRYd�4�8�&�ܥ��U�L�O0(FP�%�m�1yc,�ͻ�T��a��O3f������BIy��⼸��yXl�͙̉j��im�T���ab�]�����]Ƿ�oS��� ����uM�J��oB۠"u��5_m��r;ZiGlI�1Z̻4��t�0��S`��u=nU��b��]^k72�����?V+��u/�-^�"��m��ˑ'�f��^Ki\��&:;��6�_Ki�yRrwGbgde/"�SS���l�nٕb�h����t�i�)��^��e٪���aI�IVD�B�
����tF����U����5�ԞӘ���� d����^'��̢����u�6mC*�Q��V��z$�z"�S���A��IgS˥�49Y�mU+O癸J�Wa�q��'�l���"� �Eq��{x	���[�c/Dx,�*�f�aݼ�kT�r� .$*n�4��Zp���hZú�z&�{e�W�q����	J��E��!b�6���k9FZ�0���a&���YZ7��˼���]�&�$�iѵF�BbO������z��Į�d�
#!bĊ����f��Si7J�Kw�6�k�;{Q�ܫ�P�T*�YNmMId��ei^yY^�Z�r�:X�����ǐ��_3���H�M=uXmG�!ī�VaU�('�1W{L���R�8h��z�Wߴ9I�8��<XrM�n�(n门KP5��K̵ujKŬ�;uw(�����u�n���k@:q�����l����35����[�y��ccPL��(�oM�,!&�IH���U�����;��qf��N�ȭT��A��N��"ukx������{n��q�e۷an�jd�b
4�ˎ͇���e�R�uD[�ԭ��X�(�pb��K[�5��pn4Q�j5r���fQ9����1eL-�A��ճ*�ɘ�bf��,yr�J�)��9����u.z���2�ci�tRuM�Vv�[ˀ�n��4�`����Q�*�ּwzZ3~M��e���܄1�1�Sȫ]�h6��k�+۶���w��U�+^�����n�Z������œI�Tg$�.R�V�X��KJ;ʊZ�~��GE�ř	Nc/-Ջ�2��V������7۽���ƶC�nY���l;�/*��6�Y(����A*�^x�ˆ0�,�k1��"�C#�v�a;���F���^��h�%ř�yPdK
YwN�k�`�#ɗR�f�δ�Rc/]�"ّe'Ĉ0ˢܻהD����&o6��a���=GP���&7�4.���4�Y3j�[̩��I������o-�3*�d�2�5r�7+kX�Pp��cQ:w��jЇ.�B�WZ��E�i����$�I��^��'Ƥ�!93N���&�o���^n�h�0���[��=b=:���i�lk�&��]�͔��*�k��T��D�ۘek��,R�V!��Gx@t�gu�U(�-i�#fVB���\{(��b�5y��ܑau���<����b����Q�&ǖ�3$kV^���p&	XZywT"XÁd��yj�a�!�j�w�����q���2޺�,-%jPՇY6���a1ݽa'� e��ĺ��(���k7#��C�J0�[��J�8eSA�n;�-��Y�Y}��3.��pETh_]�&��y2�+�S�Smm�Q�;�AlF�݃�T����1�E��2�&%�+q)mF����ON�q؁�|i^Q�6IY�u�q�_M�� ��mÐ��a7��y�h5gS��,j�ݦ2��&�(mO*a��5�Ki�Mf%.ZZ*�Ԡ�"&�f66^1b��F5��.'F����MAn�̓=�iN:���q�I=�V�56T�T��\���b¢�h���Z��[dɂ8�f&��T3Z��;*�!�i$q�O�92
ʚ���B�K�!��U�*oi�Y��j���vF�V��\l�A�';[9٤�]j(rв�H2���d���0fR�����\kc[� ؊�?<ɗV��ܫw�NW.!Vl�QGXD��D���5[,m�j���̵Yk!oV�^�n��SU��*���g5����kSiVnI�Sd橅`')
Y��M�j^���l{�:��g�_QbR!^���,-��"�[mlYJ�06�YT�p�;x�n��CL+�1���#��N��n˧�ͬ��&5��ux�U 0-��q���㰍�ʰ�jX����Qd�Fd�囐�*��n��R�&K���b2�����wT7�p�A�&��MhMZU�fy�63V�h��R��j�4!Q9wL�Ĳ��6�ݑ
�"r1�:�`mͧ�����g%캺Y��2Kt�,�1��Ԙ\����Z������6�؀���^ˆf�4ti���z�R��ݫ�ۆ���ҦmnS�5�$���v�8� ���lU���S�3h'�����7��ed��يV�5(�R�fZ���i9d�y(-F�˰���y+iV��-tޜڍ��m�Ii)�Mq��Ă�"�Ñ���;O�iJ�յ�X1��s�aiDgj�E����1PJ�f,���KWbX�+�螿��j���DR|��ح%IVL�h��MO�֗-��X7��dE�h�MsT�-6��"-h��2ͅr�^uelNѴ�]���V�)�$�OI���Z�I��h4�j=��[�ƛ�Ŝ�%K�mO��ؾ�x�˹\V��ؔ�Z\��α6�J,H�Ҁ֤�D⚲�=\�U��+Y�9�'�"<]���K��]学�]$��a!u��b`����ί��Q(�-u�31�q<Yj'�+���tW��MTF#�4��p�otŘ�T�S�Wk�&����UZ��Twt��V�I�)f�堜]��T�0iZ�I$�Ҝ�'j-^-o����䜕���6�"̥֭�hN�[r�R�ijU���KZ��i��R�F���B�V�<�R�\؍�
JS:��u+\���-��$����sN
1���b�m�n���c��"մZ ���mRX䢻]ȃ��U�M,\����Z�J��P��V��1fL�Ÿ��H��=��w'�Lx����e$ִb�sM�	�RGVg_V`��U��\�fs��[Ir詧��f��) O%�m���]�D����j�L�őe���:��{S���L˒x�H�A�[��g&,���ՑE.��؎'���;�y+G�I%iX0�۽s)MY���R��<�,�Y궂�:@�S�kT�����S:,���Qԁ��X�%��NE�;��ݝK��[�mU��1X;I/��~U�b��.�*�Z����Q,�DAƟ'��^%I�ZqKN$�jԻkKV�"�.��su��VE|���m=]�jV���\�s�QKQDkZ�J�J��@p}Be�s�5"ط��nP�,�rV����l���R�X��G库Q+�ؓQ�Ě������\��i�*j��Uʹ,[����JM+J�k[�'#u�Z�O�I^�j��}ĭ,Y=���h��Z)5h4Ҥ�w/ܓG��ܱ�i��R�㥺�+ib�I%kb��1�����1$�q(�UJ���+x�M���TRo.�x������j�Ujb�OT��MD:U5(��jmZM��j�X���8�drZ�#J�$��Ž}��nB��`���iZMug왨����9e���5'I$�=���Z�jT�-�z��ڔ�\�Z_j�}j�JK5X�/�f���NԵ|�)H�ƚR��vb�b6�����T��o:EIb�R���)6�%�;���R���-<�Uj�Rե-+V��x���=Vmj1�(EV�OS�)V&3�n��`�*�q+Ob�L\Ҵ��n�j�In閳Q�ԫbƻ��+Yi��Z��E�K-D�)KZiRT�Ez�PI�x��嶳��I�՜��Ě�X�J�jY�-LS��Xk�-;O�ıp;���8�i^��uU�ĢX�֢\��IZ4�.ɦ��5.X�5o��j�]I4�8�iZ�]K2����U��k��Z�b\�[�ye	�iO�ڨ���śj�ȹu#j� ƚX�Ŷ�������V��W5q(�Gr�J%k)tY��IN#%QkJ�i�1J[ĹZP�ZȳR��U+��&�.�5o�:�'�iNW�M(�&��Q<T��z�*�A8�9Z��sX ��(�Z�R�]+O�7��t�{z:�&�s!�-�4��iZؓK�����[�-&�)-i$mJ�j�@��w����-T�$yF��{�T�����Z�+J�P&'j4�@�\�b���Q]'5I0z�j@ƚ��!�w���O喚U�4�lD���E*�Q$�Q#�Ҕ�Lɇ�G�`��V҉�v���V�Ị�iR1F����W�i4�*V
H��&�1���_oujKR�8��������t[��@����8�)j�<OwK@�Ě�SZ�k34�I�&�(�5ܯU%�+D�ґe�t�KV��Y��&qZ��-4��2���o��#���aϾo}� �7z~����0`���V����'�@�l��v�n�K5�������ub�w�ӡ� *��6g.�d��G��w��Ӧ�̚wBV�r.�����3����)���Ij��u�M�����tƝ�Ia��6pUO+�u�)Vn�4��(ov���0s�;[�^�Ww.�R�Gm.�5���Y��[72�.jor�1��&��o�tz�W32�d�\ڪnp��'�9R�Z����Ar-����Ն���WY]a��B���s2��o���y�+�]/�;#�[��Ms�U����]u��9U6���-3�׼s9C���uYؤ�:�snf��VR��H �W*d�ZٛI��1w��❉_�5���1[�R�{S��"�Q�_c�rv�ԣ��������j����o�eYN��/��CUh��W����;kUU�k�Rt�KPQ�Q*��ǪUC�׳�����|(N}g�v�z;�bar��۬c;"Ne�L>�ܜӹ��\�5��	��D��g;�=�K��ĥ�ұQ�q�x�r2�=�v��xSZ^J�.ݜ줝if�(��W
�D2R:�.�:��BGem�dl�6�Ȏن�]��4SB]U��6#�:�6�'J��5ڣ��ǟeL�d��!Qv�Q]!��F7%E���L�h������
m���85���}�V����j��S\/�8To4�r�d��u5�����y
���wM%��U�<�W,�j����lb�y��M���j[!���� 7���:��2��x�Q�:5c �F�.�a�(G]�����A��BP�[�Ӑ�p��#2�|�Y�����^��A:��7맋��z���]��o/�}׋���~w��^p�W>�)P��v@vpc�b���Yh�96��g��m�i����t-�=�ٝف;�F���!պ�r��[X��wW.RB�����|4V��8KR�͟l���KU�S�q�<{$��q1Ļ���Su�u����R-F;*�>��Ϲ�pY؅�b��Mŕ!R��3H�[d��f8$s^�i�s&͸�V)V�2�ͷ��n2�ۻ�O`$�v_���%�#�u����8��m��)�P��,X��Cz�n���Ҽ+D-i�6�>XK�74T������b쳯O��U}����֪G���s��N���a)�ݨ�g7v���/�nQ;���Cט�f�����6V
���F7��-J��V����ҾLnB�׶�����ݷ�r=�@�����{��xl3���]�i�ob�:��h��d1�7�)1IehiP˚X��ҵ�T��wYs��[�"����%Ԫ�!±��u��QC����r�w2K�;��6Ug9k���|�u�Hc����xAH��ٸ���%-U�}�ո��u,�WpT�M4i�m\���#w�^��S���^�p������I&�l�7���ڢ���i}��(�Mܘl�-��(���2uo30����%��LN�5S
��숡q^qL���tc���B��Z��ξ�n^��l6��z�nb��&�gL����>�5�pZ�7>���U��
t����f�����bb�)s�2u;=;�w�)E�[�l*�Ϊ���C��Q��-N�y���z�#(����C��z��0�Y�J.�m��TP��ю��gD�ޓ}rbc$]��+&�o:��ž{E�<�_*��mrL�G�:z��jEQLN�YI�>$��ۍ���`����EX0KK�n\ۘo,�����i ��ײ(;��xnm^Ѹ%��@<�f^��4h2�����G{Y�Ϛ9�H��YP�I�9���k��y�]~���h���k)����X�u$��l�U�}[���v�-��k	\���z��<&)��6.��/dB�v8�(�N@�T����o^m���W��ĥ�y�љ9!�s����!�[n�VN�v���	M�����{�Cjq^dP�U�[b���go�S�5�a�Js2�oL��F��`�9aM#V��{/&:�w;p���3�8�a��eb�X1��ܸ���Xt<I�eV�r�X��7p�/(*g��s6Μ������L�"��~ޅ�÷l�5{ބ�w>=��Խ{;']��*q�d:�XDY�e,)�a����2�ʡ�-�}���.W�x[��8�8��#b���O&ڰ�g\v��p��c��U�X��;z�g\�z�epkkf�v������o��E ��[j��l}J�\(�9aꔝS����T���Ce^�c�ӣd��.+�;)�b-���6�������`�MHj���V���`��u`�ve�Fs7k�E�/��+�������M�礐�8�D��zH7��8y�~XJ�]�aZ�5Y�����a3/�S��kwd���*>)*�m���2j��}iu9�s����B1b��f�|%Zpwu�[A�Ž���f�[�eCpW8����R�P�C�O`��l�vK����l��X���)̩�X�R+n���ǲ��uť۳;�#b�h[��3�8����:2�ܾ#6��=Q�-5|72���pJ����4��*�fgy�D;�\�4(BW��1�թM��U�enTGo2U����˗��Y�*�yw)�<iƩv��q�<71v�U�l�u�]Ś4��t%��-@�w#(�Ux&<�J���#o��ב���BL��ji{�e2؋��mY��"��p�2��[�´p�ͮ2gR�Z��X�*�TZS���αZ����^ꖆĂ���I��tl(v��ff��:�ʫ�Q�Z��M	��}��'vv�m:�{ޝ]QސohF�[ag%�j��*Y�t��晙�HVzk�L��q�����8R�vip��C�9m�ta�Rx��9�5fsà�|�3�;t-E����7�86�Ҿ�TyFѺ�
R��{�DbZI82��[b���8�|��s�9�s��MQZ�z�E
�׷��1��=8m+���*���z)��-����1�z��X�gG2s���a�n���c��3���E�T�Mh�t\�/-aP���{�n���r곴���F�����>����n���^:�u����fI�{�H�Y������B�4-�P�R5�V͸�& EeQ��=���7�i�%����Wi��9��-M-lα��%M%%]��!q��\�[l&��;�!���Q�<roL�]�3�j9�SQ�bA�L9D��e��dm�f���Ի!�w��,k���D�Tİ�g�d�VFP����7�,홫�WFV]zn<��ȸ&�s7���5�r�ʕP�e>�o�-�oj��S]�E�d���N,��էqJ����3/�s&ґ�����k�`S���ճFty7���B]-ƆK+7d��U�]J*N�kI�v^���t3�T���TmG�<i�k-�Q��Y��L���~�*�9����x*�-4��6�5]5d��]�+W�[�3���Iٙ���ojz�oo�:mhʽ�2�]�S*�n�O*r"�Њ����r1���\�&�c�
SU*��vL�������t-$K���8�Tծ�[�*��uI+���b��X�o[C��׹����H;";�Vd���b�wn�w����{E��ٱ5�Vj��sU��B^��.���c%}Y��s�������z�w�f��a��9g���φ�����+"�6�<��=:��Է���d�g�m�pmh�lUw�;_[��ё�=�2k{�)�.��������;��-<]p��g/�Dܪ�F��Ϊ�;�tF��g\)^m>:�L�\��Ϲ��s�'j��YؒνUnue��m]+�t��5������#����d��Kn:V������T�]UM��t�]`J�����
�+@���[S��1�o���M�����Ŏ�׫��wޫ�h�*�u�5*t���4Ej���{-��=j_=��ۻKj,���^m�b��l�]pk|�Zd�9�s���)�Tl�E�LΠXu�F�6�՝��K���Y�	oZ��VVm��qLkq��.�.1i��/*�4wb]���7���S�UN\��th�[B�v�u2��nv�a��ّfN[�l�VAȄ����n=�-��إB3����zT�/���Uoo-oKM��V?�<���קhc���t��������kh�X��ޅ��˫{�i�D��R�|7��9ɺw�;(���8W��ljI�^v�ϝM���qgQ���JB�k�c����KT�j��#��J���3�t�k������A���Ԝ��iG�%9O\-ݸ�3�mZ{w~(�n�bD�n�E�{pZ���Y��mѸ$b��w2�r���yop�;7bnw�Q�=qn�w�jg0�9��}�n��B�}j�.���"�l)a���0�/t�v��iv���nX���f]�kZ��a<�N�[}���_-|­j�9�]uԪ��u�{���.پV,�<�Z�^Q��ӳ�u&�j�~�� .�k���H:�]qS�n#ݓ��y�}8Н�<��yu֧�DSr��ä�����t�_v��nwwRB�/l�9��#V�G�ҪC��lp.
��;�ҫ3�R�p�j�$�[���73���z��KMT��P�R���ІAp,�WAm�(J�l�*ި�[J�ܵ����*tl��k�4e��ۊA�d��+x*���7��ST$�4�n�8[��
�kjosJ�Nu�_ua����R�r]>ZD׼侕]V���3igUpo$r�����Q�|mK���;�E`��ggӝ`�.ۥ�l����3���О��j�]�y�T�#��ˤ��,���ߕ�,4pm�ZU�����U�����7}�,��Z�}\ʼ�G����'^qo6ՙ�h��R��wWO��~ꚅ�&t��{���e�3FN���C[�t{ju�䭪�!u�2��T�m�|�]ޓ{JKN��W����p���ɽ�N���_N���5�G7u#��ot��V[�lN}�qSc�ޢ�4�ep%��n��ͯ�_pT�9-��:U6�"2֎�>E
�Ӆ;z��{�f��˘���lp#��,N��6
������)�ʵ�ƹjsz�U_n	��'L�'3}����]�p��j��:oD�0��YK�̘Ӈ"ss4�I&� /� ����G�b&�N�>C�b�0�@,z�����5/�b ",�
��xiDE����+�g"�@�\����πϘ7s瘠X���ߘ�۟:���}���4�z| ���u(i��Ej�\�s���1�F˓��#�My/xx�'���P,vO���+���zo��u���?/�y�n���M�{���D@O���^�u���|�Xyp: �<�{�=�_�:��!� w|���0P�Yɼ�9{Ë*/Y�� xr�Y�;X
s���:&E`����7Bs>Gw 	�F��������G�0=�4}� ���| �1� ���(4��ۢ��@���O"�=��@`��X�o0S�E.���"|�fO� �X�� 	w��τ����������@�=刮@<�sLw޸��( �������QO���B}����?��G� ()������a���~������|ʯ�F�c����3q��Q��f���dZ�7��f�PѴ+�sa�w6e[��Dz>�:e���}��*�����J�n���L�vX�r�K�#q�2;����雜_q�$D���̕���N��y��ӧ�l;=Z��K"�Bl���WQ��M�>�ܻ����p`X�s���Ƴ6��\�5�D��9[�����w�	S�6'V$��"�	�GC����2�vZB�`����"��]ҟ3��ާ�l���C�h���ƧF�\�9Զ�+�=�T�6B�9l_t`�el<;9췤!t�LG
ɒ�D���_"��k0v�W����j�:��0��_X�Y���Q\Ie�YW1LnݎwX�r�Zf\���16i���mg��%�C9��5�g�p����*�mw7��M5V�-���`�p����/4M�~���`��oǖ�4�ܧ�6,�.E/mŧ(1!j]e�����.�	J�t�S����i5���.6��Ñ��B}� ;oU�O1[�ʬ�=.W+��U;}�f�s9h��6�Ʌ�<v�y�þS�-[k�b�eǛ�����m��
�޿O_����{�w�ݵ�5�kZֽ��5�kZֵ�kZֵ�k�Xֵ�k�X�ֵָ�k^�ּkZֵ�Mk^5�kƵ�k^��5�kZ־4kZֵ�kZ5�kZֵ�kZֵ�{k\kZֵ�{k\kZֵ�ִk�k\kZֵ�mֵ�kZ��5�kZֽ��5�kZ�kZ�Zֵ���k_�kZ�Zֵ�Ƶ�5�kZ׶�kZֵ�|kֵ�k�Z5�Zֵֵ�k�c\cF��k\kZֵ�mkZ�kZצ��5�kZ׶��kZֵ��k���w����q�Ml��N9����]�5�[�͆�Z)��Ϋ�N/���X﵋���1x;&�Z�Ǒ�^��ˇGwk9�aʳ�;�LO1��	=�ܜj�ə�D�YՇfT��M�i\�d�/OfQ�e"*��q<����_-�ņ�SW����.g��rH��e�r��k��oj\�h�5�b��h�(0bw&�	5��/룸6�Ьn>&��p7����x6%�E;��	��֊���R�:�����;�\�h�Gv�b�qf6�eM���K�~��26/�N�xGo��'�)N�rd:5R(�]�T�%`��s�-�i>0�¦�3�ɝ�ۻ/�QH����r���q�(��]4�%X7w)�ҳJ�:C�"Jŝ�y��,٣M9]�'}M�w�g����V�9\��ynuys8:\���n]�nvl2�.�v�s�TS����d�����|�+�59�*��w����M�>}�%���G�,Q���ۥ{Ԧ�g_��-�S����p���Ww0n>�k`�u(���[�TsQ(��7��z�=�|{|kZ־4kZֵ�kZ5�kZֵ�kֵ�k_�5�kZ־4kZֵ�k�Xֵ�kZ�ƿkZ��_�kZ�ZּkZֵ�cZֵ�k�ZƵ�kZ�ƍkZֵ�kF��kZ־5�kZֵ�kƵ�xֵ�k�ZƵ�kZ�ƍk�Z�Z־5�kZֵ�mk�kZֵ�mk�kZֵ�kƵ�xֵ�k�Z�ֵ�k�F��kZ־5�kZֿֵֵ�=<xֵ�ֵ�k�k]kZֵ�ֵ���kGZֵ�Ƶ�xֵ�k�ZּkZ��s��s���0��9����kZ�&�W�7�öi'��er��[�Q8x�ۛ#��t�����>�朦v�o6J�s.:[Sxp�.uɷ��+٤�٩d|Np�b;<��Y㈤�ؗC��ޡ��b�d�� �B/%�V�
���gAҧR���HG����f��
��8艅ofR��M��ws�:��>�4sƅvV�*����Z�ԥYsD��턫�{I�YO���K��y*���)ڼ<�=G��yb�G]��k"���+,��S2er�Wx��ޞ���Vs�i��\ڋ����[Ͷk@���k��dЂ��R���M�0��*�u�'*��+�f,�-iI��qv�LH��}���=Y����	�`;�7ci�h�i{!��ফwq�l�JX}֧e�y:IAt�6oZ+���2��/g>�c[��̻:�}��/2�r+���Τ��H(�q��u�i��S�{[��-m��4֥����I�m��V�:�J����T�u�K��˘´:<'01:,�j=�]b�E��GhEhp5P�S�����Yݺ�w��z+�gK�]�)�۝�g_c�^����kZצ��5�kZ׶��xֵ�k�ZּkZֵ�k^5�kZ�ֵƵ�kZ�ѭkZֵ�hֵ�kZ�ֵָ�k�k]kZ5�Zֵ�MkZ�Zֵ�Ƶ�5�kZ׶��kZֵ��kֵ�kZ�5�kZ�kZ�Zֵ�Zֵ�MkZ�kZצ��kZֵ��ֵ�kZִk�Zֵ�|kֵ�~5�k�kZ�Zֵ�Ƶ�5�kZ׶�kZֵ�|kָ�{k\kZֵ�{k\kZֵ�{k\kZֵ�{k\kZֵ�ֵ���kZ�{��ջl'��&��R���.s��w$|R�;c첦�Ib	:�|��*���gS�ISm͗�^���q��'��v�]'���R�-�l�W[QS�2�E�)F�bk���V,K%T��il�V�:ѹjkk'j]9������}ˍ�}���9@r�/�ۜr��\��'�с>�tnB��]s���|�!�叢v8��G5M�T��YĜ��$]Gu&���Y�T��ySA(���찜�"ң���U����ĵ��ɦ�.�\������͒�G[Wx��R;,*͸;o-��r&���2���U��ާ�����T��>�f�+w�0gD�(�=���WS%»����=-^�7i!�xa���O���,�r�]�2�~����{+���"C�X������X7�&�m�9�ʂ�װ����d��{�h=���)�YlO%l����s\j�ݛk����_�ۻP+P�7t0]t�ө������MK��MȰ�n��(xg�9�9N�*u2v�>vK�`dbn�U�n`Uj�Gƥ��]w��g���]�R�&��Ǎq�oo�~5�k�kZֿֱֵ�kZ�ֵ���kZצ��ֵ�~5�k�kZ�Zֵ�Ƶ�xֵ�k�ZƵ�kZ�ƍkZֵ�mk�kZֵ�kƵ�kZ�ֵ�Zֵ�Ƶ�tkZֵֺ�~5�kƵ�k^�5�kZֽ��5�kZצ��ֵ�~5�k�kZ�kZצ��5�kZ׶��5�kZ׶�kZֵ�cZ�Zֵ�zkZ�kZ�Zֵ�ֱ�kZֵ�Z�q�kF��kZֵ�cZֵ�k�F��kZֵ�Zֵ�k_Ƶ�kZ��37ɽ|ݸroZ2��*6ɪ�;�2��x�7-��I��'L��r�D�plX�Y�ͪ\�7��4�3��;��{3��I&�?���Ic�aaۘ.�s��a�cb�J
ҳAb�w52Gb���湫ݻ��J���]��O:�Ȝ�I�i��?i�i���Y��K�ȫ0�G!0��A(��*݄_e5ÞJ"�3;���'����Z�j�4�m��=�& �t�S��՝1q�vWF4���j2RsL�b�U�BV���)ᖐN�,��s;��gVr�<ӽ��s;"p��n6�r6�uP[7)(w��yhྮ�M6��̻{��,m���B4)˙�Z�H��1�5ˤᛛ}tј �<�b���]�6�Xy��̧ӃJ�P���r.7�:ۆ�U,UZ�5=�@9��\�mMS����SO8���k�ݍ����n�(�G�!���6�MQ/ ��٠�F�7"f亙K�p�Uw���kh��M��|)X�Q���Kor� ��lW����&�C�|��}��m��hW�m�V������!�y��f��}g��{��Y=,-���Řy��{�w!�^�	ư�0�Bٸ�C��I5}�9u�n��ن�AQRѺ�4:����wi��m���>b�fh���E��	��ч���{U �-�ѼgT����	��yl*�4{�pܘv�)c��'��=�w�P�z��t��If8��]��$��Ij�7+U���x�<�q{���=�G[�m]Y�VOC|�=�˪Zl�S�04ON�w	9';
��L���]�D�a�
,�S��^R\��M<���6ՂA���pf^,,�l��՗�b���3u�!�{��g/]܇&��MdY΂��e��7��K�a�z� �&TK���V���b'�@��|t9��P��H+�Yw���5��eY�D�2�uSG�y]c%��Ƽ���S̮����{�qhaq��J${R*�`���-W�2����&l�{�+7���b絻7X����2MU=ӓ�Z�x�:�`�B�a����N5�)��g��-���o��u�z*��w�N
t�2�qa�"��2�����U� ud���ؽ��q��e��7^�ػz>yםX�T���7�jƓB�mA��C[�����Ҭ6�s6Z\-�9��Ǟ��4|=�l[�R�LqQe��İ��8^�t}wx%�K�4�����u<^A|��mV/xV,)�����z��à�u��*B#Y�|r�!���Qi���쾮ͮkw�lo���K��Hr��v:�ן\����ڼg05qVܓ��r}���%R��$�.Ӛ���!q�6�̨7x�fW�i2�)�r�Q:�M�^:X{x%���@{��}�NU�c�+��=�
��k��oa���8q�9�rɮ��4��N,�ƫ�(�X0c.��1�#ڝ����t�ż^]��cVYz�:�fN} ���%�B�Tn�E� ��2֣Rn���d�k�3m�*��u��X�B���޻�9��1�Yn�hS���54kz:�v+�ګx�#�G/6�b-�Fl-=׺'K����I�'���B�+.�PxĻ5��k!�x�ނ��7�)Zww6��&��cʻ�W%�lJ�����6�U"ӎ�y4'-{�����| ���Z��2ּ;]ĺJiԲ�Cηh0��b"#���8o��)������P".�A�3i�YY�W��p�[���j�7;{���$j���Z����5w��N�����3:��7�$��D�^f	s�*޺�j�D�2��C���#�EQ��TVz��� ��sQ5>����W�%��][������\ɗ��)V:�ǀ���Q1z��I6�e75`�r�cw-��Ĥu�e�k
�:���]{mѸ���%����\˵�*�{��[���ҋ8��h�bB�H�QQ���W�\���jmRU�vi��l��{�$vP��]���܄�񵺙���e{�~W���n���Fu�7��{:�bL�>��J�rpYt�G�i���f���E��*r�ی.$P��ۡCo+/�h�R`�\-��Տ��H�R�T�h��_I�\�Ҁ��x(�3��PCV��m�N�������n��-�w�q�'h�U�p���3mVlv+lnd*�gS�[�bt���1�j�������[�d�Ͷ�{��_}�:���Kj��"�0�R:o[��}D�V3!� �]�i�E�\�<���5ùvpqwX�y�е��5�DV��w(bY}���U�d1&{�q���$d\HƠlC�`B�:��&�&,��m��Le�7w�%���.����O�	Q�j�8�g)m;cX';���:��Li���t�Y�n�4;^\	S�d��wLk�������T�7���~[��=v��̮�T���1��ӵ�`��]R�fP�.X�P���I�[�.ͪ�ׇ�t�B�����.t���n�>l8ҩթ��#��"TQ�i���`�h �������Kt�aU���g7Yܴn9�vL��(�K�o��f��].ec�ӝ7���Ÿ�k�뎷�V�f�%��GK���-p���W9��Kg��Sj�����+h�y(��sl����q&�1�q�2���G�Wp�#��Eɭp��T�^�s����C��!Uv� ͽ>7��1��y"4�n3B�"�8��J�qɧ��d)�(���1B5�C��P�}�6����I��J��y��ڙϣ^�����	I"�Պ��J�Rs�OV�p�j����:���Ae�m�u^s�CڒJ&����]s�	%p�R[�wP�����9�\\�-��R����i9KE`۬�Z-�f"Tގ����{ruK[;��׈�zU}��{-pK��>����qv�^���g��Gc����J���������3�B3y�Y���t#zF�-��{�m;͐tGh����hw\�����w�}Óki��uyyn+��V�M�*'iM���Ҹ�l�m@��-�2i��Q!&�s�
{�a�zl����J���]��v\��U��X���F�K�U��K���Z�ڻ}��wG���y����}ohސ�+�&8�{�-��6�
@�V\D!���[�����X���4�OnU�[V����צ�i�2lo{ǥ���[��n-�ӱ�Ҿ}Y�Ui�D��l��cF
ե��Ք�W������&l{۔{p��E�=n�Ή.:5Z�,'&�P21Aai�w�:�qUd��k
�����5��`�=7��z�1�/쑴6�um�X�#�WAM�N��]fu��C�����W�;�}�l��×]�9Ǡ����cuRN��ގ���Yr��I��mu��O��"va�IS�`6�j8e�ܨ��{��sc^Fs"�S���f,�y6�Uʅ.u�2y�g3���?p� ��Y	���~��~�������W�O�o����<C���'�y�����w����D�.F�d��[$��!��%�)��@�I��i$��_�m�Y'B�q6�0��#b�E�qB�r0�r� Z@�Ar�_֦e%F�B4����9e�& ;���y����ם�R�Cp��$�($����)�0�$ A^����MH	lA$�Q�H����1\��FR(D�����h�l�K�6ȑ�!a��wM�4�P[M�hO@�&��AA�/D�F6c
�q�b����d�T,�
Q��,&�Q��>�E$QȐqƄh��$�AZ����E�^PqQ��JD�RA)���m��4Y@Oߤ��
&OH@n$�
��T2�d�AFF���)�xE��e�H
F�&?Fd3Nc.]3TJd���*�)"PXA�!(�B0"�a6�-GQ�b>-"	�(�d�	�І)"�FBH3(��P�H��-B��ry��\���d�h���e!�2٠�I�������J��#3�	�CV�V���q҂��	��/j�o��8z)�z-��ή�fe�:�wS��]A6&��Ѻ�i���ԝV���jH!�����`5Ъ\0�#���ɉ
�sN+�
�i�fn�ݔ��hU;�q�Q`��w�d�8U>�]3�M���\�Ns�Ώ�Tλ��b�_&�Y��Õ�A� �S2��U����n��t��ï�9I9qf�}h�\�7��٨8�[9�$]Q������*��K��'1�+,��uu4�	��ʭ��T�JdK�
�#U{ٛ��3c.fՓ���nfn�|+i���f�اW3Rü¥��̣6��8IxD���P�}	��mŃq�ԣwCH~0;{��2���i�/�a�o�@�d��]��aZ[0lt��=UyR�[���8z�Wc�b��k��q�+��-h�{�n�Y���r�O���n!L��`��V�IIk�y]:�� �c�#�,��r�>��6�!���Ow1j�Ǵ�B��0��.v��_U�x�˺��7.�%djlc�Db��$�l�ZN!d8�&@��ƌ��@q��f!RP
�E�J" �B'#"�HRx7=�3w]������p>0��!R�$�	0��`�Zk�4ȶ�T�e�?@ʑ"����j0��#�)b3��,&ہ��%3���qB*8c&$�a8�m�a�B�dPN�iE*I�-�'���B�2(S �B$Z��d(�!�e8�e8$����#BH�IH�$�(��p�b�t�J�^>pĳ�s�+x��y
�
#߮�+CNxT��
��^.4d�H#/�H�b I�G"H�\�(;���.�WΉ�/WzV&/Z��s�b��CWQ�}*$T0T���%�R8LQ�q9!A"�&2J~)��2&��%01�=��Q�(�}!1"DK���1��2�0K@�I���0�JI��Ԡ£PB��e���B8DaH��C=	M.E$^%��A�$n$�~^!�Z,�M2���(�XJ�f6�����#&�Q@�-��f0PA�fHIP�S��0�3�&$���IP��~Q��=��^"��	yω=u���2��b�[D�zHZ�E
d�hE��@��'p���
$��0���sD2�ь��m��&B��F#1�b@��m�BY���E�`i�d��B�22�(b\�:iF	0��`�Zk��1t�l�H-B|[��)�ۄ�A������PD@�$�mcqB��4ɢ@���s�B#F��8���ңW��7><�^wq�'�wEe�T��)���2�	2"L(�p"de"ϔi���QP(�)���Ĵ�̔�)BYHG�)�ٌ�.?F\A�DF� �O�`��@�I����.	J"b)1e#10�L�>����"%�-���5$�Fق�	�B�R%&�r2�ELd��"#	$9**H�p��b) !�D�yRi�H�FHqYsĂҎD���2�4�n�(��$
�>H�
��@�2G$���w��TE����l��T�!�,D���R��a���$��>=���|kֵ�k^��ֵ��뮵�Ԅv}��_�*+�[�(����AA(��-��`GϦv<{k�ZִkZֵ�{k\kZֺ뮺נ:�3 ����d1ҥ2�*6�W!:O�"|��:ֵ�kF��kZ׶�Ƶ�k���z�pd2w2��/>sb�Uh�a	$\$�1r�<q㯏���kF��kZ־5�kZ�]u�Z��/��**�N��
g�c���f8�s�Xwt��D�v���!F�Rwy��a)\�򍎣��E��bnE� '�.TM��'�(� ^��j�m������,��N~?4��z�12
/�'�Y˰
#���3��zw���Qr��y��i�z_�����l�^��H��T��g�=�u�ח�Fw<�Q9��r��G�ylba���ls��W��l`�כ��<^�#`�åE\�)�u^q٘N�0wwc�A�ؿ\��޲��d����v3�㻥�6.*y���y��R�!#�t�]ۮ�c����6���n�|���<����;^�����o�w!��_Ͼ�ŢD��˭�8 ��u<�G\Ȣ���8!%|u]�ψ$��[�������B�
>G'�^z��I�鋣��q�G*0���!͊�I/�(��� \����{�߹%O��e��$�I�% HL��L�~d�� �&Cp[P�
�L$$"Da��dPH}a�s]�LUx�3�L��<s���ȁ���TI��1��&7��sS��s�u��ca�z�s��rY}�důM�7$�7��r�\��p�襉٧0p��"m����M��(6
�HJ�l2���l��D�Q� �,@䀣 r&�O�)�p��s'OW���>x�t����Qry>tGWu��<���/M�L�$i�y�%F"��`��H�"���Kt�p��$��	D-9(G$�0P$�B~jJ����<��G-��G�/��.D��L$��!��QDy=^]眝�wx|7�3�s���Ͼ��EuC9�Q����Is7r)OF�/����*�ћ�H.�S��0�X�o"]�d
��n=�B��Ǖ�պ����������L�
��ܦ/��y�~��le�T�{/�g�s╾�D��{���H�.��k3-�
���E��+�Aʉ}�|5�Q[F��yը�'|�׃/ï]�P�xjC7��v	�,R�c�jT�ب6��79�Lc�L�9Ӟ�S�؉dT�Y�;
�T�zS��]�sN]�[R]�-�moپX�o�E���z* ��1���˫��P�G�)#6�ud=%�X,��h�v�'�X����w���z�{�y�r�ί}���}۠�H�vz� wQ�fQw��vix�.��X�>��#Uو�d���{�yN��GF��w^�6�I����Z�NcL�H�y���'�q�X�z�K����s�f�8��7s��ut�e���}�@#XeP����hG'�x��t�>���>j~�*�^8���ٽ����:�M�#*��[϶	��5c}�UK�#��}ώ�;� N�! Q�hm�����ڬԺ�,F���o�nT-u�uʃ������B�f�O�iڬGp�˻�x�|||@>#�_UVN�IYu$(��!oen�y�Ϭ*毑�	{a$o<��{s܎�|:PP�#���w���}iy�mx�߶I:����pG�A ?���jf8&���ia�x�w�sټHn�{�{ܮ���bHe�E��Q�_Z��(��?\̖���tZ���g��ߤ�:C�2fL�g܆G����WYI�~����G�𣈠n�+5���g� �_�5���׼cn�^�/�y�o;3v�j��'-{w�S��:>�)��������N�K�n���P���0\�3�v�߱���ӷ�G����{F6�|-EE���K/}^���$��VT��;��T皔���-v�Еm�E� .����:�:gͲ�%�k�b��}����|S^�*P/*R��S��op��X�Y����(�>Hh�ud����6tl�mq��(�fN����q��ZG� "�N�[Ӷ�ޜ��=���;}O��[:onwwXȭ6�m\J��ђ��S�޷<痻�l����Tu���Mۻ���ȑI"�D^{�@At����$x ٭Fs=KM��o�ldTA�|9g�}��/�>kY#�z�']H���*�E$����*q!whk<U�Բ���ʓ:�������(��d�����e�=�C��
kh��B��[M�ޖ��j�9�+ē�p�z���/\����%�)��N�!������k��@���S�g�D��#E�v�t��\��{���^���*��9�I>��B�Ü|�:O�w>��D�7~[q�|@[~��\����'�69���u�k�1i޶�3}4޶����MB�vp��H��f�����Z�˵��N����5S���3��;�6>�C�ך�:P
���|H��skij�*x�7e-,��BՕ.f������@�fv���߶�y�H��)�~l��6�^���1a��W����a8&��˻;�o!W*��)��H�r-�V��>ղ�B��9��쭜� k���	������y�i�S��b�pc�jq$�'��5i�@^o�����bYkm9�a��?���MR�qQ.g� �(Afݺ�2�S:f��N4N�xB��߮tԓw!j�o){U���[)}� 6�}&��6i�PLJ�~��?��b� �s瑓�AEK���.=�N��k[�ܴxԉ;(h:�>��/�[����󪼤gͲ�&5�-T�MW�����ʞ.�M��\�6Ϩ#�Qq��N���mر>5:L��u圦���܋��L~.��G����-��Q7p���n/m�Uhԁ#<ב������������Q�0�-�JJ�Kڍ,^��[xo��wv>��<1|y�!y�
~Y��{�4�D_�L�9U�;�<����nm�齬������7��NRmq�/���FX�n ���9!��s�ID4��,����,�ɕ�}#.G�ڵ�V��I�"��,rA�c��ι͎��Y������3��W�瓼�����+��^xd2������W-���������W���bKP���a�Y�2`F$`FO>O']�ߝv���qʶd��NY�ױos};����ts�p�f6���c��+�YW;%-��-Ű�Ӫ�[ⶻrs3iL[gk�mtH��^�C&J}@A����}�ff��` #����IC(TX�.Y��q��?�)�a�#m���Y����(a�C��ח��h`@�!Y�"�;�?��g(��i-�#+�@fJaz�&�{k�ǡ�����7�%5�<3�/�S��䔠{2�}�n���j�'��j��ug+�U�J�L=�ZԴb��֯=ҳ��ѯ�����>]Q.�qr��/U��������	oR����Q�o]@oN�:��fӒ�aR�pك�Q���T��L����]��$��8^�������F<����1Uf��09��>���l.�|����� ^Ǒ��Ö]ޖ5��l��*vh� 笭�M�y�Mz�E��y�rA�ȍ�ao
���a�ٯ�gu�A�R�U+p<�����j���L����[w���Z��z	B�A=��E�u�������6'sg��^'I����>���*�H�:�n��*)G��6MP2{�k�K�ޤ�:T�s!=�����>>O*�L*ħզ�oԞI��m����������Qxח�����P�Xez��d�ذդ�a�@���J�U��w��ɜ���M��v�A�p��o��}u�X�N�I�zTd�v�8
F���ӗ�(H�A���}�`d�4���CDޥ�n=���䫍�����k\*����e�\];pn.�ڻx��_g�h�g�>����^��Z��{����͚�8�����^�tm�aW\2�J�סL�a�6�2�ʇ�M:�r���/@�{ݿ3�faEߡ�Eur�O��~fX&(Uy^�o��Vߖ^"#�%I�5�wr��Zpҷ���YK'J�`u{+P���`���>����y��v��Ӌ�d��%qG;���V7jgj�����QJ������8�T�Y��]�p���|@>�>@�<֫)�+Y8\69e��YCu���8beɢ�I\�n&�)Ff��N��링��1�����9�_<���s�dv>��fNm����4y
y�P���N���mӒ �u�'	��qH kx{����z �W��F���Y!j���Q�\�L��n�ӚQ�
�mޣ��wg��kk��I�n����C���Okμ�zcT��������RL�����M�SmRZM斍�1n*��l�uMJ���:���/|����b��z�x��WD;C���Ɵ*�<~'^��d�h�:q�N�_�`�Y�վX#r�*d�+2��b.4� q�4����e�����7���<��T���h��$j)k6�^�Q����0F[�)]��VJP�kp���֨�����i���֩�ͧٮ}�'�Wƴ_ޗ]��q)�����6򃍹j�rZ��H�S��f^�s��W��,g���x�,qq5L'�z�=w�y|;�[��仼KK����iQ�mt�5۰k�Ə�3~��0�B�@���_J�]��s���#1�EV��=f����/nYV��{1��d��4�dx_3ɞ��8}���~ ��jt}ݗ^:�ה�߆�{��Klu���J֖��Y6�5���@`o!k=0��<�˱0�L5���R2hmŔ���K�S<D���up��!w� ]� 2j&-my[�kIQwAA��I]#s�ᚓ�L}��@׽�g�͍͹���Ѣiz�o�����&��+��^�~�7G��oɹ��ژQ�N$X�Y�+��VLi��늃�h��z�噿o�:�UE*�5�����z�Ⱉ�Ϝ�M�}�m%���}IT��ܡ��=��D��(ʪӰvU˚�ɡ�.�Vf�j��Z���}����3���>[8��d��e��j���uz��;[,1�S[�wfuј�u������@�P��N�d�����g�[U]5(+wA��FX�[�h�X�D�U�~�?E}���6��W� �E|	i"��U�K���:g���k��gr��u."ssˌ\�]�'�@��.*��oou�k`�)N���}�_�3���$`F$`�3{���2���Q��Φ튎���g{{*~�њ����"����aeot ��ob9������}g�����;�����~�}Ks<���P6Җ�zq2rQ�;��ξ�h
p�	�O7�>������z���<��?}�ox
����P��Ѡd���}�4Y^��f\�?v 45�s
\�b�~��ۖ�և�R��j=:cԮ<Ԍ�s�� f���ZPq��Cp�5	�����������_LCk/��T�����7������	1�f�����O�ҿ��`oמ�k��|���j��WO�t�{qf�lf\�ϰ0��Q����BQʗn�
X�����o����R}_^��q�ׁ᠄�>1D��� ����;�s�B^�K[H����.���y}ʠ�����Z���`�1k+�9�LiҎc`�jp���T�D
1xo۽`w|P�e�(���dp��h��AC˳�V�xY�ڼ���*Mou�"�z,9�W	�k�<R[��^^��ny�Ք�/�=t������-z��7�;#��i�9YN��z�w�����A���g{~|��;޹��3������Q��d��k�E�u	�Y$��n��M�Zl��csG��lf��o��䯳�Ч�nL��)7qv�}ΆF���DC��KN酞d�$�o�;1t�����"~�о�jǎ�o(R4��;��|I���ٴ��3X6���#Ӓ���Ǎ��J:�0�_1D��i3���6�Ϲ� �۶��Of�m���Z����� ��Ѻ�K=3�*}I$�U:���_1�V�lTxZ!��d?���	d>ژ�׵`$�;̢�ڂ�a����1i"[��Ｍ���4n������r���o*O�I���2UMB�w�f���01�x� ��q4ػ�^t�N��d�����^�x�F��Ƕ="K8#_�;�O�=���"�����9g2v�<&&���{$?_���T�X���cS\�ϵ8���9���h]u3;*:H)|�R)m�I�AqE�H�3k��n���R�Nt0��K̽�pMԯ�
!�S�V�w7�,[�t��\,e��7Ҵ����;������ȫ/NWd�$H�Vͥ�̚�9�w���(�r��r	��gwZwƣX6q�;��X�Pe�Y}.�Յri�Eza�/��V�ޏd�s�n'dm�_XU��X&��:��Z���n�HH��.��f��|P�CG6�]L��6�I�9���X��nɼz��uە.���Bd`͠����\uud�Mܢ78E�6�T���&�=ǵ�в]����q5kr�;:�__[�Ws̒��e��}��tw��m�3������:���,n�	��Y\��9v��d|U��xvh�ئ�",�]d�]�_��dtǛ��F�r��{�e��7�7�-$���4�"��u�;G�K
�y.�gp��I��Puܛ�qެ�#��NGN�j�1u��(ߩWU1;%�����@��D�������Q�C%
ڧI���_4�ؚ��G��tI�W���ҵR��ŀ[����X)��u~0�a��rş9(��A�+N���2�qA���3�K���0���M�N�j
��K�3]A�O�q1Će
��yJ���bP���~�?�k�<���kR��]��T��x�(d[&��۬�FԺ�w=ܪ���xխi���\�jӒ���3gM�J�Y]�Zj>صu�g}��J�M\�9r�,g";�n�0ַw��˶6g�W���ή�z�q�չ2���c��73�֥�s�r3�7������_�z�j��w�B����a7��d�Z޼}������!f�8�z;Յ�&���J�x1_vJi�D�.�U�u���k�司;�L�&�t_=�Wz��9����ђ��L�CΑ�������SVZ[���<��kv����S���!�iҝ� �/zd��[�tŬQ��X=�Ut��TW�-N7�;*D�=����D��;ۧT9w��]'F�ޮCg'x����R�3[�cᎴ�y���I��-���u|r�5�Bt��UL�U&=K�����G`ڻ	;�՘:��=�K�U�+=��/I~�y��na޼�_Gd�]���V���'Ů�9=.�G����:�J��K�S̱,Ҕ�� �>��:
K�A�0��H�9ˁr�i�>px�L�OIs��&��oL>^��ݽo����oZѭkZֵ��cZ־�뮾�Y��dE�h~��?���$���wr��ʪ�_̫�HN���D$s��<u������Zֵ�k_Ƶ�x�����=�;���#��x��^����u�ʪ8��S"�0�r���.O��p�$g�1ǏƵ����ֵ�kZ��5�kǏ5�z�=��5G;�wLK��(���y�)���p�=yݗ�X�W���>1�>:�}|}}}k��ֵ�kZ֍kZ��Ǎ}z{d��J��r�G�9�'�z���EQ#�yЉ�K"�֗�^D�S���$͑*BeHNw*�Т�M���VQ��^��2���*�**9]2�Y�YE�ڔ�[34H�G�;�RAtE(�"���U���g9$�v�w���H��}ޯ}[��bE�TC���PDuY22TĔF��(�6
���֐�1�;'�!W"� �Ȋ��#�EA�z����Z-�'ZQ����M)����;�u�oH�Nƣ��+cM.�+WtN�����۵�n���/�N��}��Hz1�8��8���c��[���x ��z��w�V.�r�hd�6E�7����p4��Д�&�G�S|��T�ab��_���<885Y�������%x��;�?��}�1B�I�cm��y��幁�xx#�=�����G���zn.���L�5='P������H���^�S��l�ĭȾx�����x s�܊N�$kՆ�s��,�J/<��&�W>~��4�;L"_̤E+���!�w9�ە*��8�S����/��E)?ʵ A_�x�#<}<��~�@}���~�|��G
9Q�"�o0f���-��{�� �z\�rSՋ$crz�R����Ɔ��{�6O���q{��$�7�P�0�S�>��3	{o�a��0����?�O�E�rψt>� ��̋���~0w���k�:	҇����41�0�|���Z�XAnW�R+�gRa�F,�+ӔOB}����R������;����<�i?W���X���4��<~ _lUzc �� �-���c���WjR8*��7���$�͇���r�8o5��/��}"d?7���O6(�y�izۑ~?A�]��p�[��R�<Vb/W�mk�Gd���XȤ]k5�|y(�XT��͞&��3B�{�c�~޻�ܚ���hא��8���묮�T�r�f�Ȇ
�3O��pv�
?�{��`��b�`����έ�߇�3
d�}�
�.g�}1�0�9ϙ���?�����뎗#�[�������g�� �ybۮz�N��A� d��z���,!�Aj8�g��;���1��<<=V�����ޖg�'�֊g��Y���y��0���{O�����ϝ�����K��V�u�����᝝��y���� Mw�� u�%�}4¡��M�%�(�ϓ��ak��4���{�{{�/��h|��4�|�x~?�2�t��؀z��Y<`�cǾ��:U�0�{�m��'�{`2��&�z������=��:=���\yx�!�[���󽼉i��z�l�����NQUL� V�ƛe��L��z�����{�ė�1 �Ңڜ^uN������o2��cb=]�4��L j��W���M�C�/Q�M*ux|���:�V|,�|�3_v� ia��ǆʹ�!~��_��C��&�z��.�>��6<�e法c{�e��'y%���O��O��M�U�� ��/�������A��&�x?���#ܛ!�a�5��������ư���m�ݧf�V֭� �N9%K���-���T*���3:bb�=%l�$�� �J�=:��+%q��i�H�3lۮ�s��ͳ�e\9{ݑ�/#����J�;�{��Vz4�����!��⇏��>^ 
3��'�G�����w��%Y���6zZf��L�z�5
�mUld�F�
a�N{8�;AO�����ڕ2_�����>b���E����o��矨��`�y�oS
�F	a(c�R��y� �� 2���Ͽ�,����D�a���3�+��`��A�  �4��f�x��-���W�{�6��|�v��>��b���>�2w/|��i��?����4�O��F��lE{��x���X˞m��.@�Fp�y�68���ӌ�������ɮԘ
u�b�x���L$Py��쏩f- W��s�7t��\�=2ޟ0��,6�����0g�=+E χ2sQ��;���~����A�G�[��Q
�f�#}Z@��U3�z��5.�MծY��-��Ǵs�;��&1��-�1\Ntw=���5<T� cp6�����o���,��O\��f�������@t��lM����	��0W���Oj��ۭ&!T�\�r��T��e�"�n��;�:>'��0N��a�"�@e��?�V��~��2������e[������~�D�)�P�q����io�W�`_�:O�z�� a���w#�閭�����JO�����cj�V�h뾙�]Y=jE&f�5WF:����&��������,�JM^R�Žj5�r!;:%����n��<$���|��)�u$���kz{��r��#���q�1�`�~M�����}���y �����<�����ɰ0�
���	c��<!_�Fϛ�b��]y�����~�jr�^�*3������b�s��K� p��1B�g�w��������H�_��JG��k�o�y��8�1~#M�T	�P�\����J�M�v�-$� -0vwv�3�x=����k��4����	x��	Y	�\jr��X�g3f�?f��[V}^�1_�U���%~:3������=���C�[�Ws#�T# Ojݝ\�����)�j�������
h��V��?|~�����Z�����鳱u�ip e�w��eT�m�soO��= [wwIn�/B�o	Ys���s0�Q� ��Iv��2{d��V8&������������(�|aƼ�`+���P��S�f��VZ������� �c��#��g�wϜ�r�'-G?� ��ϫ�n��~}��z���IĴ�7st���;4�����������|��8�}�  .��֑}##ݞvOV��~���%������5(+���0�3n_~YYһy�@[��C�φV[>6
�ܨ7��,�{�/z*��oW(���B>d}�",��}��`R��**R�n��%�)��X�W��V�&,���qT����7�xoD�1ノ0��88�
K瞍ĐS�z+����4o�����6H~i|z6����>>���O�w�JEp��Y�{�=��kp~�4���Q��!�@�K����"E_ަ=E�����7��]���kz30�]�:��]8\Γ���h݌i�>�m�^x�Ѿ�x�р{��������J��"^������&k|���)��@��C�=����!H��Y�;E
	wA�
4�=';8���KY�D�K�H,��|�U�ޭ?�{�����E��֎n����o6)��m��cm�e�([�B%���t���%뽑݀τ�W@��0�pE�2��β�9��7}o�p3넼��o���3ǬF���Ʉ��us��$<�p	Hq�6�ǁo�O�ed��\�9j�~Cg;� ,���:�E<yX_�(�M�j`�l	�KJU�<��H��u�-U�{͍)
rW���p/�����ƀ��L �>~�	iگ��J�?W��ȯ%��'���L���ۛ�ݣ�<R�0�#���󁽽4�T{���=Щ���v�p)�P&��cZ���`M�o>کx�f7!�MA�8O�ܢ�НY���w(/�7I���3��&n\�����?Zw��l4�w�z�͗�-͂��xƦv���X[���B�K��;�f����V�r������/����<�7�%b�� =lk��M^n>����[�`Иmcχ�x������`��$����Ke�����JŽ�?�h<dH���%��<�W�W-�[rLg<����o^���Fmy��:j��/�~�j��q2�i�_,~O���|>~~�����6x���WˈkN{��<��ס�t�%!��b�h��?�n��>��:�jϟ��4����<8!y���CGW�����2�}�1ݎ��=:ow8M�ޭ�@$���g��@Ƕ�`���d����ߏҗ�m�ɵ�JŽy��l���VF'W�r=
�d�O� M�t�[A��*��T�;�Y���U=���˕#����ɑVr���S>a���C�������C׫�F�R}���"a�p���x2��/�Bw���^��.[��2ߓ�h����h���(��ѹD5-���&��-����g�߈a7ֶ��Û�=��yO�<'%ٓn���Wa��W]����{��m���S,��j��Zh8�>��j���^/?Q�!?ۃ�����_����Y�j�(K˛�r�w�������j�&
b�o�f��D'��2����вz&YQx��AŎ��=�w4�;����!d��۩�kee���&ql���N�̢�K�t�7�2����0c�8���3����71�f=O�'�g-љ�9R��u�c)<��KH���1�����{ԭr��l���?v^]�nM�a���z�>��$
Կy�x`=�'�#1]&}����|~!�����_�3�Q7	)򳷌����cbqm�9�7�=���דl��\[;ly��h @A�}�jk�ch�`�̼��@{Zi�:���?2`)�k�hv<�ۯ,K����z����@��n� �vP
��i��x�����P`�Q�����ɦ�8�!����Bg��exo_�)7���s=�~�����͛�m��}\�E5C�y�y<��F.yק��8X�6
��2��D>=��=����ם^`�-��}�Y_O��x��w�>0;��>���q��wȨ<�7qr���+N��{[P$�<����|��İ��G�pKӭB_��?���j������Oub����g���`7�b�C}������-����n��� w��Bd:�٧�p����v%���H�!$�zS^IXG���H���\�9bB=P��xa����fc#((JT�]9����;`[ۋ���g���=!��Iz7�H�Ç�/_�����|���t���5��G�KA��z�l}�K�a�׿��)��{/�����8+��ĊA�t�y�h�T�+�z��X}�P���AF\�t�ShP��c��p�=/��̡2$�Ӆ��=��ݾ88�0c�8��I�-�������?����g����8dU04ɻ�ouDI�@���z/���\y-"t��۬ypÑ-�L�	����>�3M`%�`/��ۭ�)ڵv��.��̺����{a���o[0i`����y�y�zy2������~Kme"@��n�b��Kԭ5k_�w5J�=r�Ç�{?r�w0��~$tC�"�ެ���a�y�^���8�f[�ej��v~$����А�
>t��>c���$k������*�|	���x����E����C�[���Z���ߢ�b���T|s��6x��v�V,�NAn�w4w��<n�f0&e�dZl�����[�jW=�\A�G��l���1��Sࡺ����S����M��{SWU����>�}���-������|#��=`��0����,>��&�<ǥ�έ��J�<S�/�V�.��Z�&��/�۪s��ǿ1Sp+�d�r�4L_bS�x�q���Li),9�txN{�@�z׶~y��x����~Q�\��|���\7��6����n��h����W2�f��ߝ0��e���|�b�cwYW��cl����B&->������C��B�q4;��I�e=aF1.�wUg�L0o
�BV0�����s%e�����Dڰ�<i'���zy�<���'q�۰q�v�� ����o�\�a�z�K�2 D6㳆|�1kdy��&�ۦ)�
p}G����X�Ű�w1�^� (U�MR]��.���f��dr�o������(k�s^m^�n�Z�T�Joc&�;�`
ЈS���mn��Cp ����>���y����=9vnxp��#���}mJ<5�+c����7�E[���Y���p�݋�B�_��/W��ߗ�.�&�� ��zzEW���z��.�w*%��7�Y�߿�\>J�LO�E��$�@lA|����=��|��Rϛ�g�{8�����һ����&��k��u��z#}�W��(����~9ȁ��~���.�e4���݈�3�l�A������~"�ޞ�@�L^�l��J��C�xV��[f٨L]ͩ����Мf/���rS�z��y��њ�A+K=>�W���!�c˹��C[1��܊\�Y'xp��oA����{���`�p��}�3_�wh�G��=˯�n۰s.��\�m�QL�<!�[�X�,�ڼޓ莋�eI�������n?����[��a��_X���|��6֯���9|�R��>���F�<�8�;'u�*}rb؃[�2�:ma�N��Z�f,�<�G���V��ڧ��!}�ݻ�k]�"�S����T��}�#��ǀ�x��z= xoxtB:X�w��P�-�->�s�M�AHa� C��&*�n�<� �OG��"*!�wkݪ��f_V��������֯#��Y3i�S:�xυ;Ň��~N���C��#VA�n9�sn��zW�{|���C�
��j�E���@3�����#�VY���S��~�|�D��ϯC�*GjS*��VҀ�8���<;>)����t?<��gw�@���5 ^����Y��hޫ�/��.�-������|E��!�_��������>�v�|�|��)g5w<a<W�kѯ����&�>~���6�"C3G��Oc�z��	��[�EFd���.׶�j�K�ߡަk}�����ܩ[
�%@2+߼??5��d�/�<ڞ���-�sh��Uz�㈭<���Q�[���F�3M��.@-��#=�9��q�i���8�r�in�Ѐ�O�pr�Mr*nb_u����?&��+ "���w��
�t��(�[�Wk����oJ�=�"�a��{�;��'��z��Ld����xiּ�s��	�D@��:��������*��d��]Ůi�ɯ"���?hk�}��P�����o����Aq���pRƌ�r�hQ���QJ�X�P]�F��o���pXK��!�Lu���7HڶGw^�f�M��\��-7�+��ܒ��gc��1�V�˅(9�\ζ�:)�@k/�LT�jp�f�$�w��b唻�^L��W��9y7����v��+*��D�=}|%��6��}*���
^Ɯ㼔33*���w��'�.c7ף�l[�:%�uu�,dZ�Ԓ�r��+�V�#��|ɻʺ�����A�<@��e��7�s�ە�Xݪ�9M}����l��y}8�!���±��)r]0�Фz�9�ҺJ�C`���7��:'NI4C��(�Є	-���,��T�'N�߯u���D'IUWӝ;����K���j��^_�8y8W}������cB4j�^l��9��r���*:����a�˅�	�����VT��<ވ@�7%P��u�ҏH�fH�k��J���e�J��fӡӻN����m��w����ԕ�":q��>hԪ��q.�K�J�7���9^uWb��҂��wmB�h��6�a����B�o�k����AGU�]���$Yƛ�%a!)U���k�i���E?�&�i��j�P�j!�P�J�M:�͙���a��)[���->�FI$�R(P�QhO��ssJJO(��P�;�	�e2f�h@�N���xF͸ޙ-�w��������7M��/�Qڿ)�vtc�aOl>ő䳃a�0΢i�[Ȳ�P�ͩ��#�R,��ωK���p���P�QF|�hW�����ݺ+ ��p����5���u�Den��Y�'|h�wn\N�:���0�W,QjnN��V�̯M��!4��{�E���H��gdf�hRӡ9V���J+"�ڍu��N|��r�\��v7J�ǝ0���t������OZ��U�Ԏ�M��7���N��Č��"���"n����)�`�wn��Wy�s��m�J=w�\�뮪a%Q�p����i�u8�/:J��]��ī���Mǽ�ؿ�q����t}�\ҫw/)����# 0�wb����d�R�N��=O�e%�tܾK�)���s8ں��Z�&vlO�P�i*�*�2=�'̤��R�w�XIK��ɻU1&�9�1���˹����� ]���vnS6�������IP�egG'K;]	7,N��W1Xv[�(U;C��5����&���Xc�U�^�3�V�)Wt��6�hպe��?�Ki"",��r!0�~$9Ȃzo(WȅE�?;����P��D��3�y�;wg:ݼ|}|}}}k����ֵ�kZ5�k�۷o������J����L���(����ȓT�E�B����c�x����������>������|hֵ�<x�׮�	3�V�����ң�u*8O�"e�gC*Qa�2.DH�3$1�ֵ������}}}}}}}k�F��x��ƾ�l����\�4N��k�E��;�s�����QVD|ε�z�7��ֽ��}}}}}}}}}k�ֵ�=�}߷�}�,��9G����*�@��ABIEʔ�����H�mPN��G�@��Ƞ�m�(/�
DQU��x�!���.qG��uCf"�r;<���eDp�VSđ:����$ADP�N�*sT�)ƎܪT/ȦUʊ�=��EOM����GI>t2*yG|c�)�y.I_T�-iE����DUr�<��s1(�{�������wx�>�p�/�:�a�A�DĀ���6?Ta�)Q(���$��ㄖ�	�i��P�m�QL�$I0�r4�d@�~D#M���b�����RM�;rK�S[�wgKOv���:_s��Ocw{MGz�Wp�}2^�y۪����?(Am7CE�|�83�Ǔx�t�+!I������F���I7m���h��gБ�"�-G-���CHb!�`D�$-�E��lHL�#x�
�h0�� &A$��~,��18�tL�7Ey(�DEQ8�H��,&(ĐPD�~�&l��m�⍘cM��,�%�NE�Bm$�!'�!R8���'8~����N<2'3��x�\ �� ��"=������A�RF��s�Di��Oi�_oG�g><�2���b]]nLS18���0>��e�'t=m�k�˯��~���T�m��^� �)~\�g�]3��./����j���vS�AAA��b���/[p-��bأ�+��(k0lo��vp��ֿC�,�'o]�T/ݐN	�,1�/�Ʒ%����ќۼx��g��:�@�|�(ƅ��4�ֶ�1�̧���,S���"M�w@�;�����fM���.���)چ�ן�lx[� ��>��`&&={���������kzRȼ]z� È� < xI��4��K���G�[���`,!k0�a.��rt𩣠�V6u�V��A���pȦ=�E�3^�G�����x���B���PuSoku�@���8O���ѐ��C���}23�t���3SH���޶�Y�)旟|��������|z���|����w�up,�7��un����� �m��z4/=��z<d%���_�nGEo�v���oJ�u�O}uj�K�.3vFz�ޒ�Y§��?h�I���|�~@h�Bƈ#]���ޑ�S��ۋ��Sڕ���^eҤ�|���}(��͔}ܬ�������?������f�q*1:������w�����ɧe+wo���u�[���Q�*JiGk$��]|3b̗'Ppi��B<�j�@G�=7751pgs��6��Q��q�*V�;�7��2p�}�]��/9�)��o]�m�>R���D��q�c�gv����۰�v��G���	��gwOpڨƴ���2+��rU�C�b��{=����c�?�(�v�[�M0����f�h-N8	��ݧ{J'���b��nL�_r��z/؀���@��7���mx�������Fc����J�W�7ThS������in�Z
��ෆ@9�-[Q�����.�`E<7��;I6��ږ�T�Ec�r:�p,7���2��!��L�I��q�=�z@,&�����?�'�o���c��Yc�d��n�b���<=��5�k���;���Q-701���:�����k� }��s�L�kW�3_�~�Ft��{��t^�g�����u���"Oؽ���`�o�W����}w08bէd�����t���!w�'��'}^���!�Kٛ ݠ��������'�ʖ��9�s��e�ZPL5�a���@̆l�����w1D1V���sh_j�����L�]���͞sN0v,w�	 ��*!����?���Dz��e�;{�&5��*�j4i�{3{���o�;���n��;�gȀ�7<���(n׫���!R��DSۘ��R�ou���=��:��ڥ����W���+�u�M��}.HWr��"/�>�O#ݤD�e�>�I�$��AE}�U�ݒ�;���T�Mf��zy�i�R�ȹG�_V�,���m���XP��í% K�� ~5��@y�1��W1���^8Ǐ
E $�Q8g����r��.�35��z�Y��о ��|}��b��M3�������x�V���a�k�x$�����cz �>�y��k����+�%�c�����B!^��s�Z�����#ËM����8�K�c���Ð���� �����(�/�́zjN%���@K=L �0���d���]�{Z}��[�p:��,:���f*��+�(gȸ��_~W��=�=�0�{�&�s�R�<�<�;Ĵ�<r��s�|�����'�ώ��q �Jyv*{�|�}�����$�>C�ޝZ�S�~�u'c���;�]�pю7�5��|���7j5�����r[b���09�-�؟i��{���f��4X���0�psυ�#��=~00�')���6�����4�6���hov7�.�\�����v�� �@�5�C�X����4࿘����`K��O���q���y�A�>���Wشf���6�������}���|�7�RA%��������i�Alot<y��p8Qm��b�\�}P�8s�2ml��r�< *��6k�m��8Fb̛��7����Ս�<Ջ�����O��]�]ǒe���_�7�,�-!����cՕy�� �4ҕ q	^A��\���7�R����4��W��q�n*��4����=LI�}2632��Rvޱ�Ѳ*���2~8���ǌx�P1�<Eq�<@D����]r��ߠ�\k�����>�!W���g�~�vf����#_��6�� V��ώ��CKsٵh�<Cl�{�07�R��[z)��(3��333ςIL���	�� O��Wm$+��}�ǀ�a���!�lT���>�J�\_����=K��.�4$�5{8眎�� ���>��Td��%?|�,p���Q3���V�����^�����G����_?���Nj�5p���ސ�q�:�o�
����x�����}�=����1���F�6�1r��;΃G��a�@	��NZ��Ȁ�]����N�����2��P��K������5*]������fo�����C�b@-������ΕE���c�%�=�O���.������.�:W��f�c��{$�����g���W�u���Y[�*�_�;y�=�ݻ;x��Ү��H���i/�|ψ��9u����K��*1��#�Z�XB�eb�}~���kk��Qȃ�l{�m�g���p�[@
n�.���!�oѭ����=���\�%ݐ��	�Ǯ�ׇ�u��*�lM-��ܽ�A������;M���S���sn����@ֱ�3����D�Q��x�����[tzáׁ�>���q�,쵾�yv��k�ny:U��|���s<���{�΍�⯑ �q�o\xǏ\xǏ C1����B"EUz˙�d��9��]g�}ܼ�$�d��/;u�F�Ik�N�)d�k$�o��+qҌ0�g,놺�����K�����{��)��7��0^���<�B9-�oV���X�b�
Ul/�@a`g�~�F��ȿw���N~>ŀ�i����O5�Y.~K7*�� �m%�<0ɠ����L��3��a%�`4S���9�!�	��z��$ZV��;s�:�p.�����;�_����}[�{��!_ /Ω��=H~:@�K������@�Û��_L�"�pƚ��LxN>Dz=�#'��� w8���u`+�1��i}�J�Vi��z�>��/�V���y���<[[6d q}����W����Y�;�c�:`�i����!! 2��q������&��i���& <�z�E ����׋��|�:g�;���=w!H���Ȗ�)7�TTw�'2.3v���Nlkkn^��~�
�>������bo�Y~�|@�-�[�(��V!&�s����J~����kq�s�~�k���G�|.��"&=M|�so1�sg�ګ"i���	�ߔ�_��f�'��|+��x�n�a���H�`��ߣ��+�U]�r�pf��p:j=2)zm����L9Lpk&<:�)��;F��DF� �~�ql~��ڠuaXPq��\[���.Z��#ڽ܅�|��ǗO<�k�nf�/��>���_;��חБ����J�k�l�|k\�NF��3q�p�ˊ	���'��.�ꨁ�(����^@N8ǏC1�� �gv�91�q�Cl(��7fi��<]�(����8ҽ0t�~6g���^��`C��@n a��a����9����u�<�0���F�<gG_���
�e..}����XS>v���(]U-��r�ꜜl>����Zx?G���c���������2��n���_,5�"b����b���=m罉PM����ߣgHצv�H1dOĎ�ӟ >�#V\X@�jo��T�fY����=�8�e{	��ܺ�{���dL^��4����V�Ur%��SxÁ��`�����\N�~�P�O{����c�@�iY�}���7�;������9�Ti�ە�m-�����$�E��O0�k��>�~z�PXA�a<��V���m�*�*��������@�L��_�[w��0��4Gs��,6��o�*�Xu�Ζ�������Cc.�-�3�s�p/�ާr{�|rs�{��7�X���lv� �Fz�w�=�z����t�/�_����Hv{X#y���>Q�~�@N>��GݡH޾�W���g
suA���y�=}&ei4O�Zy�O�.�����o8
ǃZ���r�=�eA��A]�cr�n�t�c���z3��:�#���\��n�^D?c�\xǏ1��D�1��@�D@HS�|��Etp��www�D���s�X:�hi�w��(A�O%�����H׍C�ݍ�����Ց��g��f`/}���f��<�}�fC2�L&��A�O�,2�]�p @��u,N����xfmч���9��E�~p�)��3��>�a�ǨG�c���	m�Nی{����%&��`������W'����R�6|(�ʌ=<�g�c���N|�õ��n���@y����L%�$\57����x����C��|US���>^2�8���߸��y�����皪u�ٛ���x��M��^��2�` �N�*�C�������~V@��\��f�+G9�W�{Mp�-8��j'��d~�W�� 0�L��1�P���My�Lv����z��I(��n�爐�� ���X&u��=�m�j�=���y����GtqU��[=������I�4�SM4Ua����2`&�	���M���|�㢛����¼����8v�dp���8�(3} �~�l�xP��ЪSǵ��u��n��Ks{O@�q�]=�n[�>U=��)G��Gj
	��K�'�J10K�p)��.cw�o�`���k�h�%�E}&M��Z��*����$v�\�C�v�N�ٷ)���L��}��7�[;�|�\?�X�x"��<x��<x��#Ȋ2
-gr{�˸kfע�����>w�zhB���f1��!�j��/�"�r�E�ϭ�
�ږ�)l|�{��O�.��-C�KF�ia~_�~yd�T�1*�����*ϟ��(�w�����X��|�:q���]'���f]@@��C�<��0�VTx<tc_�q�3��O�k��l䡙f��S]��W����]�p�	�_1�p-\UR2�-� c�i���	n�j�{d�9���>��=��D�#m}\�����?U�|~�<��^���z���cw����75��L8J`��������9cD��;�\_�]��}�ύ�wA��g��M9P�w[y]Ԁ��R��It韼�� bP���i�@?���r|.)�B��3G,���y�6n뼗��U�Rm�8�Iٱ�0��z)�X�����K�1����T=[�^O�TxB/����
h�.<��4[��r΃m�ڲח�8A�<��C��c=���3��:;;����:Uj�'��k��n��H�4{TU��k&<�|�{gO�.|�>���a���*�%e}^�v��Ex����x
��������hƂ�;nZY�}]��:��L��v}d^����°�30|'U8��5�-Kf��N�S��*fm���W$�-��9E���L��q��� �>_�q�[��vې�k;�Ż;�`T�dA �C�}:�׿>{םu����C/��0�rO�[�u�1,�|�g^�b%�7nv5��.Jn�ێ-L����� �E�0��l<Y��b��#����,ޔ�%�����ʟ�Y��2.ar7��R0�c+���Ƹ��F��hP�u��q�#ox���x�^�u�1r�-;C��� ��$���@A��.�Sh)+:�f���o��ǌ?~T����>|�%�t�| ��^)��M�x��R����sҺ�q9��i��%k&�d(�@/�c��t$;>��������/�zz|�-;w�;�u����ݐnu8�H�JE4�Q�.��r���c�sl���i�x5��G��<1�ѡ��u�{1�Rݳr�,���)���1sH�rza�8c:��;�pဖ�ρ��6�]*��{��u٤��I�׫�Mכ"dT��м�nj�u�����nhw+Ϭ0�c�:sO2�;٪+L�՞���_��^�(35N�`x�l���&���������:�ip%�-|�W�fN�l�{h�D;�y������C��ls�	|n�`��g�������sg~[^~�<�d���K�]Uv6��rM���{�c��ׯ=.9���=�kN#G�p
�?Z�}�����W����{Q������g:����������ɶ�;ra�׺�OE�mMz���݋�m!gޢ0�D����N'^ce�֕L�C{������u�Nd�.��ow�	�RGB��;z��t��/���2ٳ&~���>� xǏ1��W1��D�y���߿:�ovy�����1���'�^����v��)�:�a�u8j}y�׵J��gT�/�;�5�;0ĸv �>�`'���}�����F������ۊ�����>3�@;n���/�����}���,�y�k��m�I6�����5`�5�}n���G��Uqm �'�p9��Q�A���W�Lp��cC��l3�(��G�a�q��y��z`�����@c7�G54�C]lyel� y5�]�l����s��ϟ��rg�O��?B�@#�	>G�~��
2ׂֆ���y��ܱFe,&�Kĳ� ��M�oO+�`)T\<zEk3�h�釯�Lw33P���-ư�7�.���݌Xzs�����ɍ$�sz��.�8�ZY����H{h��;se_ǖ~uu������7���R������m��|���=�
k�T��dO`����,k�o^�����S�;Wz#����{�\�HJ X��������	�.����z���	���-/��k�U���jcy'wH���`ӄp�ڈ��bn`�Y&�QJ�j��l�	]3Q��4�)/l͒��T0�Bkȡ��?_�]�̙͹*Ȉ�έ�z:���ݡ�/E��!�ݧ�96�!G������-�s�L�:�`�9Ǫ�US2l	�zV�\ã�u�LUgy\��W�*׬��:��*�ʗA9)6���cw�,��J^n�$>'�Y;˻JL}z���,�oe_�M,s67̢�[\nA%���L��0[+h���}$����j)ɮŕ��[g�`��ejf�N���.=lG��(�iF�gw�[�"�Q��R��$���u4�K�87@��Nl��bn��V^����ˁL	�MV����G��,�3{�����VvӢ\["q�xh��em��y�ٰ�ܼ���h^Ъ�԰��o'H��ygMZ8Ky}�
��Y8>l'��f�;��Krm��e��}��ȭ	EgG6�7��+�\�������K�J1�Vp@�q*+��p�j�ȝ�zQ,��V�L/�%s�eb���N�,��WݯeGe�Xni+����Ķ�#(n`3_K+�[�VU�<`�6��y�=<��c���G3�҂�iJ�Az�������y'L�/,#	$�!XETd|Ā<�K6��k�Eg&�n,�Q9Ǜ�5��&���T-��c���l ���l�.�"ɱUu߬�(��d��"0�r���l��l��ې�Tc^�
���e�@)�(�5C��=��#�8��^~�}��I�V�q�1�ڮ��\���X۵b��J!���/���mP:�>�y��-y��[�ƚ�r�+e]u�c�(2xw'N՟�r�0�+����8=�X!�݃R¥�U�LXN=�0�M���N�i����ʆ�QԨ���R+��a�nq�"kJ,F���\W�+/����t{��ӗv�ܹa����@��n`k�J5Rv�o����^���܇Ϸ���<NL�f9�s�yHLu��U�k5�ȧv�V��p'�t��:9&����Z�*
b��u�X�����N���G�D�X��]����s�nwtn�r�;� ��ZA���&�,T�V�]6�9��9��uhq��gv�A��]�v�n�k˲���f��WS*2on�U(B��9Tם}�3���R������d�A�Pٹx;ئ�|5���.�c�j0.���܇�kf!R��[<�]wJ#�Ӝ�V-�M�q�w�lULo�9c�f8z�����
�)�pR����C����d�ES��k݌O�>>$I �������G�`;���*"���)7�mJ*�t=�>kN:�ƾ��mk־�������}}}kǏ5�������̒�PQAȮJ�r�d}�\�HA�d��<xֵ���Mkֵ�����}___^<x���o����dT��G�s�9AG"�đ_ԙD�s�w�HF$���I$�0���Ǐ���|k�Z�ֵ�k���������Ǐ�{��E?����UDW:��UUE?uʵ"�E�REo;�2��y����۷����o�ֵƵ�kZ���>����x���{޾c�XE�꒷�s�=A"�I�*U˄r��q ���Az�m�> �'����Et���".�,�(���h��B����gS&UUEAD�%Qr"9�PD�ԧ8����ys�EȎW#ZEUʬ���(��G"5�,�r�*ΆK:�q')օ�)��T9AG*9�9U\T�����փ��9Zm.E�"H�h*^)� ��#�Q�n)�[P;��0i�e3jɩζq���b��P�ʄ�s�>��v�~yC-�5�C�wy�]�'9�
O�׊	���c�<x�
(�����/�}�0��N�[r���?������t��/��0�8嵽-���w�2�]F��1]\�����Y��'Ʊ+_%��!o�CO���į+�q���ֶ��+�վ��+q�[�ݼ��#� 0��(�����7�'��7H����}N,ڳ�w0�B���Β�z�����榯*�f&���}�C���R��d;yN����LCc{�����n�z5"�\N��enf�g�h�,t�xh� ���s�#S�Cq>w��^����N{�v�⃭�6N^�^?~�'Ґ��g�V[�{��,v�:sC�I�����{`K�#�O C{C{����,R�)Y�l�e E� ����rO>�Ӧ} ;O���]�V�6�R�OV���g~�	�G�5�B:������SP��\kdٝRo+���M���	��>�̳�ݕv�w6jݴ�������/I��V��~�,
��|�����i����:�����\n��7b�������o= �%��_�������1�-���û�-��EkQ�KߴB1`��]�ɛ�	�l��̷Y��g�UI:
��īs��f/i�4|7J����Ӹ�%,�>�9c�+]H�,�<&>�E�mKo_�Yw��"N5��գ�� �_�����xǏ,U�x�1�<���#�����CϚ"�	1�`9=�>��?|��Z��4	��)��i��Kk������3O�r�x��./5;����Gύxc������Il� ���5�h}��Ɗ唭 1�esǇn|�}ܯ0f�;Z�B��֩�Ey�v4�&�+)�8	<�h]~�������+�_V�F���㱝���[�a�mg#äTcsp9�k�u�ئ���t������8s�r��>�F	p��O�a���]�9�'L���@)q6�c����cJ�HK�6�U�����h��5�}�SI���w�-���0f��~�-��9墚��lj��hhh���Y���u�nY��,<[��M/~�4=�x��-����)�p�k�v����D�LO��xP���_%��}�A�����[�Al@_G�o�Czt�i�:����kt��OS*��a���/�$��Tx^�YQ�ռgv�x3�ងv<�y�x���vM���w���q�m�F0�lx��Yۡ�/O,驏�Z�N{�*�[�5cG��B����{b�����]����+d��Ӊ�vҰP��#N�AM=\Йb�\�{�:]U�U�drD��{��iޕ�P�b�T�uSfUFU�����FΜa;����ޯG���
<cǂ�<x��DL��o�����-V
�KU*���\����参��`��M�a�#�Ց;o�\(gT���=4��u�rݢo����gÀ^[�xQi4/����+�D?�b��ߧ���-�=^�/
o�"�Q��PsI�6[������>�@��-Q\F}�zq��ўo4��d�0>[J7e�>6dʃ���ќ'�Bo���a��d���-�_��X�ӞzC����>[��j�鈊���|͌4�{2�p��F�Sjǂ���'�^���L
w���d��U��v[wCj4Ѕ��k��~?��EQ�߯��>q����]ΰ�,0����$�'�[Ó�`�O<6�2Oǒ+xm	�}�8A>��[��9�薂,�43�/���b��s_A�mdf��gz�����;,ȩ |A� �yϗ�X�<,��.�~�g����GG���:�E.w;h_�1�Oi:xyqY\�ϷoP�����2{�Y�ݗ݅VF�]�gtY�b3����VS�-���� _�u��,)W��y3k��\[��= .i^z�7��|���&�{����1�ܰ�^y����]>vK����-8c�F�6�}p����5����k�͓i��`�S�c$���\���T�/m�/���]���
�?��ľE��3n��(� Q�͌������l��Y��2�,w<P둜�����[r�f�\���bN^�=������*1�� x�ǂ!<q�H�q (3��۷�~�ߏ�"HY�������s��&�V�Y�����͉�����v�4�X�A.��N����y퀏k�q�
dǵ��j��q����d�=��g6�CCI�.UI�;M�7t\�D�P5>�D��G=���z\n�jEs>���F0��ǧ�_qgw}m������@���A����(:�_�g(C�x�/���z�BP�5���$�/S[�N�7x�d���`�� ���:��}j4> ~�C_:.霼�[f��o�����x�������T�ހa��b����?4-���ǽ[��}3k?}}�G6�/�0��@�~�"�k��;�]Q��|���=�o ��ZF����0Nk��x�E�pj�CC��=	��O- ��t�8��P&�l��2o4Y6V<N�Fu�G��Ǟ�]��G����z��5�>��z��?���@X3W�$Zv�}���������M�WVS�P�C�U�����=��-���ic�c����ac���O~֎�o��8���OϺ,I��ן?��R��,p�����=O�몃I�ytВ�,���xU�����l4�ح���ΐ��-]��$=�r�����}Z���i�}�J��:
�����ǂ�x�ǂ$x�ǂ�x�Ǌ	Ƞ����o�����!�N1�����;QM�z �y���������@�{�?y�X�|@s{���3��p���>qެ�#_�)��������H�@�ܜU�7ױŻM�J��|d	����66� �^U"��* ���|��ye�D>үB�~��-�|�_kt>���HA���Lc"��i��˫c�Ny�DSx��{�3<�Mz�Q���+��|�4/���	0=(��Ņ�<�.�Ö�Sw:NX��I�3������'5��������c��0������T�7���[��y��3�%ݺs����3����[kH/N���姼s�¸|�|��Ɵ���J����-d%x�GU[H�Rƛ�eWU?�P�=_u��@=S��L�珫|�7/��
`b��is��9��*I����Ɓ[G�8�R6")&�|�^<>	�_5�硯���yO�!��g`>����7VWXЀ,9�9��}� 	8EL��x���߽H�x��G�P�,��|��L��m��w���ɲC1�ln�jV��v�:���wId��]��/�]/����J�WZ�W~J��j����<|5�?��� �����9�E�>Q3�Z��S���뻭�t ���5���/��*�'P��:xs3�K���?G�\x�G�xǏx(G�x���9�~������>�p`_�N��d/��¾�d�"eE� rV3�&���ra���W�Us�[c����W{+���!T>9|c���R�0Z���U���Z
�����Ԥ��҆s���#���Ŏ=w�  ��&�h�	{�ܸ�"���m�:#غ���껨H���n�0�]����-�0[Ӻ��L��G����@4Èd�t��u�욯z�1j�������4�����M+ ��Ͼ��>��RԵE���りm�z+vh�U��iW��D ;g�|Z=�_��[�:=H0jL���5W��c�/l�����as�/��8�
����6��������� .:hL�㢜y2k�\���!�H�~>���8Vk0܎�S�W`�÷����^����� L �����19���!ι�~�9���N?Ta���-�WC}����Vh%�J�E��>~a/p# p@�6� u����W,���[��e�J|n�.���5 >�y8��7`>��H���8 C���u�i^T��-e����n�ޣ�ʅ맼��6�
v�Urp_j��n�����[��2��裉���AH鍗:�>=�wy]�C'pk7eL��2�WE����7���{5(��ѩ,l�y����+7_]
'�>��Z���ACx��B<x��B<_�����������uw��Nm���Z����������*��=����)�3�F�	;B����F�:h0�п�u�{�]�5FG#��F������Ί��2��x;�������G�zG�ҡ.��I%a���d/~��5������f�l�Ŀ�`Q̡/�(�A��g�i��~O~W�M��L30`L���7(������_�x����`,C���cC3L�+��K��󟋏;�F0��A�jOE��Kd��/��	���" P�;��h����y�9~N���4z���Z���y�;I�߿L2wIT�A�|=����̊}�
J�.#�p_��_T�k_����ߙ>�NY�eS�M�)gFi�������(f�o���q�-dU����*��� �����-�e�'�����r�N��/w��ψ��@B0�1�gB|��9I�t	�a"���������Il���߿_���H�����f����<yz��2,���`_�VW�A�M����ҕ�����JR4Ì�%>��4_�%?C���ޯ�^�����=��^T �эf��[�Z��üK�V<����3�`������T㷛�� YW�ش�V�1����y7�!��n���r��؅2�/���u�um����w��L��V��ycC���`�]j���{����M`��eǅK�{�6����ݷgm�c&k���՝��^o:�)����I��~8���R<x��<x��<x��@~���}��8���F��Q{gh��vC�s:
��*=D��K7���������L.�q���NlǷ��ss[X��7"����<���ߕz}��~������c��h��[��=��3?�4�O��s�G���4ޡ�1=�x�=���_��+O6��E�;�kt��H~���%��1�sIp'�1��k���8@��DE0n��"f���s���0��jn�S�{�M?k��ng����\�,r��gw�ƼU��WjJ��a�'�M�n�GX��{)��_�7�HW#��j6�N5�nՀ�T�r C�}�p�Q��<��昤���;��Ɔ����>�'�w��?R-ҷ���M4�]�F���5Lk3B�����k�n�� �������=���.\rn�r�e#�iV/@ne�5����F�3?��QQ�!�c�������o�W鉧��rr����l[�כ��5���[�����{8i�|��71힑��Q.T��m�h9��1�ͧ��|n���_;6ozsX�]�^�V%u�"���j�ӡ�۝�����n���Q��(
#�͐>޲�R],����1�Hu�PNT��3x������ߕh-0�1���{N�J��o8�����{��w���ݻ[�gv�n;�kpl��9{VwUΗwp�1-3.������)C|�_����	7�@}���~��~��Ap1��#)�Q��"��;�V3�N�"�\A���@G����+8;���C]0�U7�a��mJ-˗�yp�?9��}G߇XF� ]Vh��H�~�'�f(D���J^�J������T�4����.:P����e.����u��G�S$?� ���~, |fcȲ��;y
���m�:�fU�j�ߠb�OL�}!��yR`r�ƳQ��=��t��: S�'^_/�R���GN��3�;d&5��^�0����AW������"I�����
���A�@�Yem���l��k+�t��`t�0iÒ��;��-Ҍ���w%#<B��5=��m��ء̶̴�1��G�È��'�/��}������>�ig����{������s�W���U7k��y�o��?�K(�c �R�o����!^0���vv�����S��8�������s��h�T��p���M��a��ɑ��+	xk!1�%������N+�AYb��L��w�m�v�Ƒ�7<��BU��Gc�fڒ%�૫ɒ�_�b�u��2��8}�2�D}	 y|�/8�����Fu����!q�Ύ������\.�5 ��<�^�S���R^���|3?AC�����B<x��<x��X�� T�N���w\u����h�a!=ϟZ�/n�	_ 4�
����k��,k�K_u��K�5��Y[��W�g������[޾���l�H�2[�пXO���M�3����m�A��z����.����qs3gx�{k跐�#�l{���� �n��nM�#��sW6)#<�F�����ܲ�7_~�$a{ �d�*��e(�
�4ʖv�k���D��0�R��j�z��hj�}V#󸦈��G�-s.M���l6��Z�Q)�y}�ӑ3���>
����̧�Z�^���2�}���%�����{B�-$C���b}��/~��^u��
�f����_��3��5����ɵ�Y�o݊{��M����6z|Ƥ�q��f�	��;���ŵ�s���j���[>]��H;u�������\Ƶ��BW�)�zދǖ�[�c��C+�v�����maxFzA5��c�~�i(E���u@��	�H����<Ǽ<< ?��d�|�p(���Y����c]�0�)���=�mJ�}9Y�Z�TVmN"�޽��(�="�i�w`���.�]��x��P���aFLU��])�^p�KcMl��ѝ�i�o�g+��B���.�΢{$�^�˰C��`:�(pZ�����E>�§��:]a�X�zD�n�\��Ua!�/���ʂlX�+3��]��C��)Q��ێF��.V�x)>���paG��YM�����w^,f�w���L����i�:�28+j'L2�-�m'������Sgrњ�Ѓ/U�>�����L]�cVM,�wI����]m�d���Y�}R��]����\q�Ϯ��t4̪v��;҅�t	�z��\T�3��Х#�x�ru�m:-���aH-�wx�����'���0���A��]�(��QȒl�gi�]�r��w�#E*��Ƕ�±���n_s��,����#������{�֪]�m���h�έ:����v]6��p�S�ʧ:�I�n��mY�8�Į�-,tj��UL����/�P�ŝ:�F�}�HaZ�Ũ榻V;�P���NY Ү�J�a�n뛔�˩�F���u� �Xo��9W��:�"�@�v�L��W�#v�0��gK��1�[,v�1�HX4����-�
A�ַb�m�/W5������K���e����c���)��$A-dʁe��*�Uű�k�K��sV���l��C1nX�5�,=���m����3pf�\�nLpկ����G��e��a���wX�חh'�;Nk�!q�s�EP��e��Nu���;��o�x����s]u��xҎa����w�mL��/�P��_I��J�q\~.���<߷���׻iT&�7ՃU����R��7��t��CD賱��Rݳ��j���3Rcjd�]�Z��XGjo��_Q�\�ts��\]���j��<��U�U�'�$WR,ڰo�S�_���Q��dM��n��襑P��,V�{1�1&V[�'W���*4�[�s:��ٛ�0^�JNw��Z2�-����T����8ּ��.�cþW�F¨��ꏫQ�2R�7:p<�.�6Ɨ�^	�ȵR�`̦��bM�w{^�
�$G���)�� A�����u����+;S��'�9:}�D��l�Q]�UeoQWF��L,�V*�{X�q��)�E�=PJ��z�G���翟��w�WH�H���$ȫ
��Vd�FI��Ʉ	�q�ǧ��5�Mk\kZֵ�mk�}}~:����{� \��r*"��:�S_zGG�\�@E'��=~����_^�_�kZ�Zֵ�{kXֵ��뮾��'s$2a�d�a$?�y������.U��r=BM���E���*<�g[��_^�Z��ZּkZֵ�cZ��㮺��z;!$�I�23�,9�(�Qr#�
����U��E�E���ַo��Z�ֿֵ�Zֵ�Mkֺ�뮾���Bp���a	a�Vm6j	9���"+�Dr��\��۔@T�_]'���֐U^g��wNU� ��.a@ʪ��t��reE̖G*����"**�3�!�!r�U΋J��W�(�(�TD�����r8UQ�����AUUXK�h����UTW �Qv�@�bUS�(�*���r�
>�9G(�(�T�\�yNDQ�D.��^Y�������c�z� XJ8�nI! �A�<C�i�-��*@�Q��`��	��D%!Q��q@�NL�rBJ�i��9�<�:�IGtx���H��[��]~�����Sa0JLǼy)͸�<�}�W]��f[��L�iw��{�(24�B-��L���%����%AB�(2�m�![�-7�M�\�-�
��Ď�HP$a�ٞ^Lƽ�2�F��-H�%�K��$����bJ�8�i�i�&���R&&�F��@�(Fh0Hm��`D�#&"|�R beEmai��"$,�ў��I��@�AA�i�L?�x�׷�� Ǐx�<q��|9�f(�.u{o3KD�.'=�<W{�����3���`��`.V렫�2�:W6m�}�]�s�PF�1���傢5$��b���E�X�*ay'\�S����^��O��M��o�-��<�g���B@��1͖���Ňy�-����z������a�4��W��|��(�J�r��c���{N�뇮n��:�x
찥k�S�H��ۅ?�ȁ��y|W8�ʛv�Yۋ,�B����Z��_�P6B��}j	Ĵ�/�g�3��4��)�R�S�h˲}�V}�c��8��&���0���T�����~n��	z�@O.�n�7���kq�˰���<z��k�^�9����-�����4�UR2�Űs��P�h�&�y�7l������\8�yb�P�2C=���1/�3]�{��?A��X 7��E,����f�.���ݸ���t�����A���B��>7e����ȭ��T\�wvw�B�G��7*_��hw�`r���A������M�rCb��*�\ޞ�l�)Ut������ve��oFX�m��g���c��t�sT�>)�~F��DrI
#��-��ˋo�t�JG{�1�X�v�����]�x��l��]�=�\I��q�a�@d"i I�~ik�a���fP[����k�:�6�>S9���,�j(܎��j�A�q�];s��������!<q���'�����=�ԏi�����{�g�>zv-�C�~&t$m��*�s�L�RÖ���]�v�]���C6p�0y��<�~D�����@���I�Gǻ�����$�~xIA�/�=���f���ᩃ3pR��}�~����&Ց�O߾A��aճ�<��{��-a�����j�7aWN���Pb�&E�ܧݐ}X���C`�tk��%p1}��i�_c;"xt,|j	흥��z�G<'�.�h��l=B�9F���Śf���9�a
���+��>����[lf㶾���!W�,wt��!�q_+k{�S3�e-�\8p��8�^qz��g���[�~�-�Z��"����y���Q��~ �BMeU�d)�Cw���0Zذ	�w�\�7�284���6��0���/;�Ȗ]e�L��cD$�{���}�CHq|�ӎ�@��9�\l�=�1��^t�B�!d����o���M��>����ցNX�ǘ�>��Uzw�cd�c�q����G|�芺�m5ݙY��ˢ�$_C��o
��4��1h�<`�>��I��Yf���k��[��8�Fϙ�#x��yY�Vm؝h�v���P�ا7�T�N��7�:�7�^s��rd/�s뮺>d�9��Oƽ8��1ǎ<<x��#ǎ<T~w���_}����I3��}��(�q�f��ff�aa��K�d�0���>k�x�󂥬�0�,�}����߲����j�^{(n��⬈�<�š����J�i�0F5	��;קi�����4<K�I5�Y2lOA�bL#���������-��l��ٽz�t��R.[�P�ٯ)�fƟ�>���)�K��ǟ`C���h��K����7��)��{�Z����_�5�z�	��b��p;���UaX���ќ��:�@f�dp�a lE�Obj�j�,�9�8���6W<�pYj:otno�
����b��o<z,�;ą<��>��3�T8Y"�����-$���~�T���a���6���6�1���O���a�'�,Py�W'C�g�}�C6�NX�d�JNW�Z��*�)�)w��E�ك�&d|�����=�B��yq��~x\�:#���z�~~��/����J�`�UzF3���^z~��P�tp��3�$�3�3m�j�y��-n���{筕J��Z�p~8��6�]���ooU�-)A�e..��[��x�6�t��a��mF�"�D�^�$���(B	�'ҷ�l�}�6�fN��B�Pj�;�u�v7��'�"���+^yբ��_H�ݾ|<����������ď8�#ǎ<Y��y� �%c������O�}��ݼ\w�B\�V�{2�#"�ﻜ0n���ċ-�����n��׹q����|;}	�~;�������O��v�~�#\pf=8��?S��������1�h��P��_���~T@�L%E�	��p�w�
�s�)�9g����W۫M���?gAl��P�G<0�wǰ��m�.:0�p5?T��^�Z4�xg���k�^|̌)ϱ�����>5�������-?3�K���_�/��g즚5.��o4���B�-�Wy�S���^�'�˨�K�s@1kbL`�Ն_�W�>��5	���M҄~'��]��<�pUi��}���3��S���z��u0��|��y�z��Z����ݳ�s�X�Ba�'�f��O֢)B�c'�W���g�̫����]�d��'o�W��8@/.�� @���5��������-�@2��?vj֞�Uv<!�����!H�	-@���e{Y�'૕������A����C:Q�3E��w���l�-�ME}#;$ᆻ�뗃"���;D�՛p�gO<�y�Z(��!  Jhs{���,Z|������DPbt���]��k�L�6����otu�:$2ogq��<�,$�C��� �8�����?�x ��59�"c\f�[7X���j\}��u��OF���ȃ�+%�\�e���qc�.c��ܶ�6�'����*�l�F��x+��~@�EQ�SVYYa�����	T���=���wZ{t���{6c�k�ā�~jGP�r�*��;��y�a��n�/v�=����������e��~^ŗ@��{�	����[S�+(P]�;��6��-f�s�Cl��'��͡9�`��]03Ly5�{h|��c��=ޤÚ�R7���ݟ����&7�ꉟ/֡$���?�U~^B���,�>,���{��X�Ag�}Jk0�C7_n{8�����U�0��dN����-��Z_R�04�c��<<�섣��ƫh�۷�r|�^��s�R��H�HX��/��_:�<���@�p�d$�Z���X{Q;�/#m�Y����>�N5��mt>�yw�Vy�L��G�7���0{�{�'���%�%�\�3Lô>�Ý�أ*cXcM�#'ư��s��\�|y*�~c��:jn0�� @> {g㲢�{����Ŵ�=gM�a���[����Dn d3���1�ܣ�S17]����F���Mc���6''r�=w��BkǁNc��yԟG{��O'������}�;�~=�D�(�"�?�\�Qr"���(*{���I�$	 �WB?�n-�[jj�}��f�I�;|#ǝ�a��Wl�w�2#�w*��GUv�{��"��{�����#ǎ<X��<x���}���ߑv���ޟϾp��+�l�k~i�`<��P��f{�Z�|��"S�:,��Tk�w�ɲ�L��	�(Ο|�Dry��=	v����I�F�� �&� �S33y��������^�T�{� ����`O� z}+�>��>�7һ/��<�5�M^�����fI�7��K#m�G�n巍��ǵ�*Q��~f^�����N�˯N"x{��c��"�V��Y�@�׿
�@I�֍��{BM�7�6�;ӧ��b&=�j��Xo���~�LN�v���F����X,cB�"��C�k��.=)���#�O�vCy�na��y��^>��_N�n#��v0�p/��`+}}�����[~�C�H���C��ڦ���Wp�+9l�\)��L�+�.:�-<��aVQaBo��~C=�!t&�iZ7����g;
��)QΆ�_[ZF?��g��}����Z���b�\�!��BK^��_�Z[�ֻM�����*�J�i9&��Y�ϴ�HZc�Wc8(��\`�AE,͜7q��5�oa��37A��J{R��%�S����Z��so��*���S�ޖ+#�WS�^�/O��N<X���8��� ��;l�5���w���X)���D�_[�1�j�Ԙ7�Vŗ������L%�<��Q܏�^{�Ѱ���R�.Z�n[�X<��
7f�F%�i���j��|�&���:|Ϡph�6��72fhڔSmΡUq��
�Ɋ�*�<��頴�����t�UYf���	��`�������06�m ��as�L�0��0������ͦ��&.��i�<TO�[�{���=!d����!�vO��I�kvLo��m��l5Cn-�5~������񿕍��2!�Oֽ[M���`��3�ɝ���V�L���Y}I�?5�2|d.o84���|�	�b]2iOA�a�׆v�l�.ƨ��<Y��m{����0��ӆ��1�e�%�o;��Λ�Z��5׉��]7h���s�����/���h��L~H�_/����b�r��?pY��U��x'�鮷�u[�4�t2�A�8 	x">'������~���>G����^#i{�mi���Τ��^�v������r��uu��"�|�^�yKʳ�Fu����0)
6�˞���P���-���`�<�t �Y���=�x�����!�l�D㇓�l��n޹������$x�ǈG�xOG��� ��R�w��!�= �l��x�b�9�$�c��{��͜�DcI�UzY��a�\����1�?s��'=>���]:��v�R顂K��p/� �����;ъm�ݚ�$FCy��;s�7]�����li��͞��*�����'�j,�b�o���މ4�a�3��V����3tG�q"@��)�������P*��+cgMl[?[DF�-�5n]���ߨ��8/������E�A��#��pl�^�"835�l����gg5����L0����5`���8|��Xo��_/�A��V��z��U���t�^�.bg����%cDH�1v��p����������}�����э����mm�rپ0X���c��,
Lmۓ�3���[�?��^�D1�z�B�,�%��$6�`��Y��)�v���ӛ�v8^>�ڧXH��J�U���a�QL"��j��^o=���օ�sQ�Ԭ?H1>��}��+���a����W-�D���;;���`���Ã�㙙���'�6~����H�`����Q�X�	y�2Ҙ�D����;:�E��l�]���_+�cҐ��Y�#�0���闩���N�]��[ǳM��wL��&H��{%H�Z1����<����m��	������88マ^^c�]�u��s��1�P/�y���������Ѷ����#�l^:h���B��VB:���罎:�Ň2N��5�W������yg+���K��e���X:$�֒��Pc���EWT��ނ�4�@fq{�&�_�}b�ڪ���ϫ����q�>�ae�4wŞ�ܙ��#-lO$O�v��\��,#�I��	��(��Y�����BY�M���[ݯ �ݹī���0!��o���ʳv	�x��� 4_���c�y�4��,�WO�nْ���FLȤ�� �}~Oج�ڞ����5���Iظ}hg�c�0�ps�p��AѪNN��[3Տ 0u�"�xǱ�6\�����	QaGb�e�;�v����1�+�.�h@g��;nib�׾�'"}u!4�G���;�������ey�m,��\���>���Y�E Ʉ5�@�=!س�{h�"��VI`�	{1+*���:�6;ĻDo����%=��B���;ͳ�����S��ǆ��G�����n[&L��X�-2Ut5�QW�6�{��Xuƞ����ˆsd=Ӭϰ�Rq6"���P�Ƿ<���izp4Ͱ|j�pw�l�Y�&��e�5r�:֒>��K��&�[���,��C����_��zXB�K�����'w�d��C��Q�dͤ˵]}��%�.l����޼j+����3��K��{����y�??!��������yR:�W�žO��µ���X�S(��N��k�f֦�Ɲݛ���@�m���a���(���-�u7�K�����Y'�6����'ѻ����X��� k��}�켶Kd��$O�	�|���ư֛>R*��Sվ�uwP%�436ϴ'�~��r�Q�R)��я�3��ͮ>��y�w��bA�y^G�>\���_��&�g��u���z�4����,��s~LP�.Hr?��42Ԯw��B�l��t��矮���l��A]�&���#���ߋ`#>�����A~	�G��~�����g���s%�u�K�D��M>yph��07kk��	?Pf��7�$��W�}�̋��ev4���9�gz�u������/O�nJ��X��N��A��a��[T�� ������h���]��1Y��k&v�{��aR��>v��a����3����9�ڡŰ�wߧԒ��>����ɭe����������z
Ԋm{�M���_7�{����{�̪�/+h�	���绎\`�&�d�:��p'�/����`+"�G�Z�i)�-��oWW�e�H�#1ѝ�KXy��/e7m����ɖyv���-4Ou:J�v5v��»�83.`|,�qf�AT�]�NBQn�+V�N�@�]��a���WzDR�Z�;�ќ�Th8�8���ƺJ�fM#eq�����<�L�7���:��X�� ��H�/xn��ʂ����p�;nM�i<Ggf.p��ݾq��b���t�q+���Ag�W�$o�ќ�:xB��&�+��WJĆwL�--�L��]^��?R�o�ٜ���r���GJ�c]��bք���B�_]����E�����6h�w-͉ԧ5�v��8�M�1U�����W!7�r�N<b�p��+����j^9k�r���}�=9�@wZW ��GL��Izk�U�P�Z��}-����U�e�<�<��tgx�cܮ��Wewrj��]��C��^�Y�A޻ ν�O04�g��6f�|�eڢ�1��n�O-vj���ٸ�2���*󹘪jhL�Ĳ�>��ό�gbP�[%�6�>w,��*���1�ُ����!��m#M�LϝC/M/��&wkD�Z�`TUعMT�B�b���(e����jS3�t�6�b6�Ԥ/��G��=���\�^�9�[Q���h\B��O/���K��>���w@7�;'���ΪҎ#J�C
U�ƙ5�,u�?�\xqͺ�I쉵����j,��C7*f�p6���� ��wcX�);�+�oZ��bÓ՝����B�����J��a#��X+���K�QIx��rK���j\��F�;���9 qU�=���=�PX�m���x��+&3�46�yU�%�W���-_ojy��ީp�d����&�fќ'�)�B�.,���O3d�{�\�G���R
lY8���)ͨ�����8Ӄ"�2�����&�v�o�!9ac��֩�^�C7��2�L���p�lVsܕ1`���}p�IL���b���I�wv!p�.�p˪Ni���$y2:�:��:��S8�֩@�[n�5ق��&�'p�x�U0������\������/�p���n�Z��=����8Z|t��P�/{��Y�q�%����^@���c�j`}M�����{aA��㱋ʖAe5�����)1��qY��L�X�V���у��7Y�*�cEjW/�Ͷ���x�����&�2[����f5��Ƃ9^��\���j;0\����|%�M��G����j,��Z�iǙc�HZ���\���ӫ�W���X�d�lU���b�)�|O�'ĔTUW
������⼮Gia)�+����y�o��z��kZ׍kZֽ5�kZ�뮾o����젨�Bs�p���[�?��p�-dE�,�r�c�]}}}k_�kZ�kZצ��5���u�׷��I$�"��h�wph�2�\�9fJ�.D��U:�Zݿ��������ZּkZֵ�k�k���y�߷���]����8y�r�'ZY��(���s���Uɐ�<u�������Zֵ���k_�k\k]u��_^>w߃����_���nlaS�� .<�Q\��U}ZsЫe�	s�QAE�r�3TH�RԄ�B숮r�Uʌ�+YE����=$)ΔUZ�T�T�ȂQ:q"�(��M
���iA~V��b���\���J���B*�(�;4J�S��ʫ�y	TZ��UETEQʝhQDA����Þ���̗MG4C}�%�R�$�i��yW�_��3�vM�R��.�T�Ng��p��vfz���<x��<#ǎ<��[ɯ��M�S�Dș��(���~�"��7����O��l�[O�w@��!��
=M��L_RKL{��F��a}S�QJO�\��rW	��d=?��!��fM�m���Y�RI5�,����BFK�O^�Pm򃯬[}o 6
p-��iw���Ls��wN&�_i��#�k�X�<룃ϻ@��涸ܑ;�p�F<�����k
z�j��x��&�!�g=��C����c�R��6�}bܓ�;�7��yN'l>X����];����������DC��6��`j��z�Zc�Z�	�]\�iU�f���ξ���N8Z �m�u�x��=�^��by����[�x�-��x��ܟDg7�C
����,�Q��mc`��Y����gp�֎�Q�
�VG�Y������q|�q��,,c�]�g����P�/��V�O��sk�>??��8����&��������N��U�$gS9T����&#rr�nʏ6�/vs1�5�'ywA�f6(����@D��ezA�S�0��+��M�P�r���C]���ҩ��2�*^7�;Rfg#y)өYx�5;��Y���}�	<q���)<q����=�~�����W�$I!$$Y�=������{��I)�HS������f��Y�m�+/��Z��\ۘc�����)5X����;�����d�B0*wg�y����q�3��sM�}*�CJ7�7Mt�O�p|rL^cYH���2���(z�>����G�.�]-�"Q�8Mנy��{c���ז���װc�(q�=\����E�E�v7k{s�ʁ��&){D�D�Kn?�`���!/�������3N=M�刌���V*�5�.�S�J��G2@'��h�k{���o+�8�X/�b��b���U>�^�Ǌc�Z�f�v��׏���^vOW�P��$B�N @Ƭ\kؒF:]����L�^�+A4Pm��Խq���;��A���J��`bc�U�S� ��910�h��Y�YrT�~[S��!\���p8��B���3z��ـl�gR�󷵉�U�����X���p��|��M���\�������y&f�^v|�Ω��}pq�q��9�韾�k(���dM�5����f����rI���ӎU�Z�B�`̘'N�ck�n<Ѫ�]���66�i�7gmݚ���ߚ;'�d�w���g�( :���rS(K]n�����jkT��I`{hL��PKjN��7C�^��c,��x���-ū�G��*��t�ǔXA@`T��B�����U*���|�vY�l�t�4���]�z�z�<a�35v6�E���316�U?�L7����u4�n4mkN;e�b�;/2�s�]b���[����U�cM�P��-٬��]R��sN�6b07{ v�������8T�m�`�hS� /ƃ��S��.���+Vѿ6�W��.��@�LOb�#;f�͑�Ki�����|�M�1˟^G�ܞ������׷���� �*��v�~�O7��A!�>��z�����q�+nmXvO�$��������N���sD���z/~߱�]���,��S�b��(�����'3$ۀ��������E0a.�1U��g�YWC�oS!��oi�M�����s��}ֲ���L��gד���cUĎgr�J�}��[��q&�^�q�#33��w]Ӥ�[(�2�:�}zu��q��<x��y�Ͽ~��7��B���o��]֏sx����.�GK36�*�$:O���z9h���6s�i�:��}C��&1��'�����jW�ޗs�/�OT�yZz�f����?�� ѷsh�^��@ey�>��]Bq��+Y�`���Y�3���NA3����*?�����T?&�+�)�%Uot��CI<�%�zR���k4�y����$��d,�ZK��V�M��6��-���$����<����]H�lT��3�~f��}z�8Mq�f^fz=���������l7��f��Rݕ|AD��r���6؝��Z=�&�Lr K���M����l��1fLe����I3,���숌j��H�A	@B8�1���Z�{�0<����}T��J���w/MF���k��Vé`�����)�o����s�K�>�h'6kQ�U�����V���C�ד�=�V��`w���=Uw8�f<Q&�i���R�pېU�߫%��{M4$)^وt��GxN�k
�<����s��lSE�mJ7}��f����u�fg־�8ノ88�����Uߍ1{3��B��p���'`P�?��|wX�-M�nJ�-J��޽�=�M�=�沿����v���j��+�K{������$����|��B-��l=N�`�HE�\���^3&�ޙ��W���YY��0dGv�I���%z{���0Ѭ$�n7��器��O�w�&�ɰ�^�`��̐}u�W��S�DMo`����J�����-;]��
�s��	ϯ}*���}mM(�5��&�9J��ׯ��*f��P�oi�.e`	���Io�z�2�D����skfR�=����O�����n��MZ�C��y�#q����7r�}�X`���Ü]�==A#��Ky�k�v�-Idsϻq�Y���h�}�;і'u��}3ߏp?|�J����
���|f�n��Xb��+N����d�(न����K�q\H��d3�ďa�}�gǅU>�y��`2�3�!�#bg[I�̂Yv��Kwt��_kW����sp�{sX�>����������������,���K����3�'�X!%���"�"z��5�X��p0����i��� u�v��v����}����/B��[�5M�]S�\e[�N�*���7y���d�g�_O�>�^���M�W���qE��yӇ�����oT�����l�v�>�ӑ�U����`ڼ���P�藺5[��t3���<x�R�)�1��8����<O�(�ݴ1���戫�z��e�k{�w��=�_�P��4�W@��t�n"��v��u2��(ԋ�~���V�~C��O�0����z3;�f$:�B�{5�/,����Bt{��]��
�9م#�鐢j��ԥ��)��w.�7z��0i9��#����筼�5���p*�Kj��������g�)U��#o);JCQ~�7�1�(	�O�UE?�;�1���{%��Z�ͳΝ4⋳^=x�V�Y���͇�oK�t����'�B�I�֒�	Z���qZ���^��}�3&��3�pV�-��9k:��~�!���<�������u��e~���U&dt+^�$���x�OLt��e����޷�M�e����c����t:�er��ݔ�fnLwٙ-T��r�5�y��k���{`�p�k���6 �޲��g_R�+�z.�3��''�SK_���a���G�Ty�`��i�Y�XU��ǯ�iƈ8�c5�h��y�n>�m�.�^2�Ott�<٢x�zױJ��w҃�yf�贖�iƭR��Z��S?O�r���K�%�x��Z�۷Uk��Z�^Iz� �ϳ�x1�ڛ�h�"ޠpN����]����!7��<��"�Ym�{�"eoO�S{��m|��^��Pj'�*����v�F�+��9ث�|�-�W��_�u��^��������l��|�1��H~�T&�V}����f�����-�r��='#N���Aw�6{)g�o>���ؘt��?K�_����W�I�d�"D�S���{s��w�E��üY�A�U�VO~�R��w+)w���Zٸ�ͯ���ipgb�Z����j6��F��p�M��߆�{�B�K�Q=�_u{��ָ�;X�qw2���g�+��FN�n�^�u�y���%��9��Y�Ϭ~88ノ88㏧z�wa*$0e���ΞY�Z#L�z�xS�E���R��_&��ՃV��}ç+�7n7�O���t�xz�{����ކfk�?���c>�J�+ܢ���ة���n�K3ub�Zy�V}FJD�Oj���S�C/��V��6疲՛���?�h(�󦹉�f����k�����h*�Wqk#l���{!n���)����s=��<4X����&�u�X�[����I���9��$17��R�}�|�ϺE��vZ/�"�&�����X��!�S���o�A���w6yS���`��o�����0����F��IR�.ooh-{�Ϗ_���}Nn�]GW���T�*�99-F�:��@D�%u�/!�|�n�%��$%j[Y�Ҝw�Oٙ���-5�h�~b\J0(� ��ff�޺Z��@Fv!��e5i��k���7;����N;���T^���W�n�=�{n�`١v�m�㎜;M��jͣ16{L!��A.�Q�D,=�t����l1�杖x(bǮ�L}q���:�uG)�ޮ�x�#��?����yyy//!���������|Y�62Ԧ�Q��������ڃ_��ؼ����ݐխ���T\�h��t�=�-`C }���e�`@t�}�����sP	f��?;l�Q���q4�,��Yt��0�"BtS�ֵ�a��fP�֍i���P���ߞ/}^S61�S�0�{@L$���ϻt�6�U�U�����AH�<��q�ك�5�X�`dlf�`S�#���*�p�מ��o~�yQ3�}���|Mh��v��<M�A@ܢ%��]6T%�ƶ���k�a�z���֪��w�Li�;�/����|K�[T�>���%�>�k���3U��jIzr<D����ͱ�M/,JwIkVB��|�v�-��ɻ�f_�FE�[��(#�:!�}�hǪ�W���6a����&�(�Z# �V~ίC���R��
@�X��ド��D"
̹��(�٨��y�TǶ5�V����0<������+'��ve���T��o�VXF��4G��3�w{���y��d����k��a�ɵ��b���91��/&ǽy�Y��/���/�|q��88ノ/�&�.8��%�採|��@��zN�]��5l�pO��Lp�ÕZJ��B;˞}dMς�'<��Wwt������nS򜸋��szY���[�U���r7L����x���{��_��L����Ng^q�<F�XH��n\��~���8���5�3&�����cz�������b�e抑���w���L�9�O�t�a��v����0am��=�!??�ʞx��P���*����.�[��Ǔ�������W�x����
�BZ8vS=����@�x��=���`s�M�w}7~�n�ꗖ{�^p���G�:����h<B����ʯ>t��20l�enf�����*��8�,��"���� TWvK\�8JL\�u&�yujъ�tߙ����4]�k������%U���H*xW�٧��E/Q;�b�o1r��vڙ�ic3T�:N��A^�؝hwҳI�V�xs[ܛ��ɻ,�ݝNW5/O�Nf�k9�k��.����*n�pE�i@��#���S2�nADs����%�lF^�]]h�f��N��X�L+�5��}V{`kT���Y<����f�幽���ޭ���)M���M;�nr}Uٍ<`����97E1�1�:�@Ү۵��6
��uV�3�\b[���.�Ǹ���s��^�c�I��V��٫�9��UZxY^�'E�KR�$��*�H��_M9�-U�^U	(��G�L�Q���T�y.⎉���en��p9��.}�{���!�bǴS�eVn��\@�{0���sån��5���%+<�&:���-I�yQc:�e�ׇ�SqW^V����˹�Rv1P�C+9���ꔱ�^�s���r���M�OU�F��NO{�MW�𗷚\G9�z�7��96����զ�9�Â�Ԫz�S�P�J�*��Di�.ۮM��GV[���co5�L���̆r�yX���vwd����ʢv<��'|I�m(�,�s�ҝ{��>�?��FIUjqF�8ݫ�B���\I2J��8|�P�ĺ&�'��vCm�y��N(�����&? |.#�	�/\>qp(򐖪���4��r�K�.��q6	�아��e���qc6����[5`s��.�n��d�u]\�$�b�� u�rhAo!�Y7�����U��a�m�即l6�=������+�ie"��S�۶/w ��sFEf�Vt�#���/mI��u�8����c{��K�ӯ�=�2Ω�t5�"\}Z�=o*���,�.�2RyLv�ո�uk�eU	�WB�=��P��v���@�@vd�Ǥ�[v�A��q�r��ݬ�*+G�2��/0�W5+�'�/b�g!�<��اgv_��n6M8uJ̪Ow��r��i�f�6���f��7;�X�����:S��	�d޾)#W���c�|�36t
����"���u�:�	��`��+lX��j�b\��̰S�0�I��f��|��P�*��(������c�a�[�VJ!����h训�fl;V_Qt,_e����|�z��u�++�{Zv��Hd޸��ڪ�[��6Eњ��R����ս{�e=���Q�9�x�C!�^b�l�Rكb;���3��[<���AED�A\(-f,��_�w��$���t��K���|k�k]kZֵֺ�~5�q�u�뮾�{�HBIHȟ)Q��(��<��QaA��$�"�V<I��nݼ߷��v����Zֵֵ�k�k�k������{�|�r�(9��A+��<�.�r9(����𜋄X{2<��	�^�<u���O�}xֵ�u�kZ�kZ׍u��㯯ά?��֨G2L��tӦba	�I����Zֽ>>��kZֵֺ�~5�kƺ���y�o�?X�U_�˄W�Ъ9�C�TP#��1�ߜz|W��#�O�y�������w' �4ZG�����o��=q"�AU7:EDj_l�)M�i��iVM󣐒���l�Q�G:AȮ$]dQ�S�L��G�iQ�R�U�Ъ��!9��P��L��y�P�N��AU�J�$�r$�Z�Df~;�Ȋ���������ʧ�Ȉ.��yAh%<�y^v��T\,�������@�^B�W��L- �2�x<G�'�w��x�Z���%	�D��$Fp �q�>�	��1!�� "!$ (�Q�K�E"��!��)���EȈ�8ח��a��{�woj��ۏn�;P���ӵ�!��3��m��k�Wú��
>M���&6�'�(�%0�R�0�~P�H."�`�!q�#�1�9aF�`ĔQ��q��%��,"I����n@\i�?"Q.	�jB�E���x�%�% AA�QP�l��H�q�"4��@�A�[#!03P��Q(���b4ёD�h
��S��iP�@Ca�#HH��6�E���AC"d��1�9���pq�q�7�����ϖL��ߢ�q0�Bs��]{��xT��=�c�E����A���*��s�F�S�D�u����j����}�Z����n�P6Y�S��}>�&����e����}��m��9�h�cR�(8 ��̩}�1P
�,�U]�!s�UԎ��ɻ*���L�K��/Y�hL��&���3��WY�[=�	�z���8{��'��M)�O�WBƯ��~���_f��'6L��?{�x�Y������8���V�P���֟0�`ܙ�^�U;4�=�Z��Q���tT]��{��`��-W��Q�p���Gg`�����7Q���A�t�MК�gݛ/ùk��}b
G��K�ج^R�N�T��xgI�x,��?��VpW�����/X�ˤv�x�r�g:��p������+����8�@FNf��H��\F]h�%�3}�LubR+=�>ܨ�g���dO�Ѹ�A�Y�d3ʮ�r�p��_K^駹.�n��{�����ZR��,���w��X�_i59��~�qYMl�K����Y�Ȇ|���in9ݦ���e���<͂s�N�y�:w\1����ͭ�
{�_=Y.d�+jq�FL���pq�q<.����F���׺��G�Ӎ����Nk�k�&��eT�șq5*�����/���}{I�0�՝|����ƓlHX�7� f�mǴkn;� D@������3�{������o������zl��D<���-9��Ҵr��]�>��!��ϳ�Äj�θ\hT�if��i�N������[��I�A�fye�3�|93��;{ЧSk4dӵ��8��Wh`��x�W�٤9��NȽ�?�f�M�9r�9���X��<f'��b��G��#w�z�ø(���r�ж檞��.����Ë���>��%�ؙX���"�x��dJ*R��؝��\�z��u��L��k緭L��q��m�̌�J���Q�F�ew�Z�� �)�qlgf��?(��qWPϡ���[�ԎV�,N�.�ŷ�:�\�x��J�V��gr�<Xk��#HU���x����F����
������:�_/Ċ�:�8�\f�s29�&S�r_�⮨����g�y������8��G�w�w���}�X4�35Ȓw;��>�PL�9�ҭ�*=q�g��z�-��۫��e�ss�&E��6�m%G$�pspn�;{�^ɷ��a1Q���#Lo���8<��N9�9]��!.���n�lvg�M9���h�� a�ݲuD�Q�=�A-��}�Ђ�'�_}�Ϸ���.�q2�M ���jf�__����v���,5��Z�=��r�>Oi��Iir�����e��}�����|�{���n�a���t�z���2�������Q���Y���|xB��3-���vn���ӛ��SZ�����fb@��?��x�L�<���Q�1(�N�k;�L�}�]D_�����3�00��N���>�P�jq��AC4���$�����h�3�z1hJ��>���S��;�'#��{�38��Vm�>�u�1�Fi��YN^(�E���]UFr�{��uD�D���nr�s���_#��H�X�g:��:��v�5x	�&��s�.�"�_3���SFss�^A�G�*t�V�/�};;���ノ88ノ8�wz���ګg��Ϫ��C�BԿr^ج�Ol&5�R=�te�&�DM7O_f��I�6�nR�u0Cv�]�\�D�wG�7O�9��I�Z�1�C������q�ͥY@2��z
ǽ��wPz�0�S+u�WN6nxZNa����b`V� �{�NԼ9�gP(A��)��0�r�7������}n
��~}�}���#�O*h�WP�v�bl��ټ'/c�"�����\�Ł�H�����h�4E*�O�4����ϐ�q"�r�rE�U{�@�7�ǖ1���x��-s5�W�X;��od�׌���3�@�7j��;�c�"w��0��N��M?<@y�?`�D�]����2
�trE�1�k$0Q;�p��*4z36P��O>KvV�Ī��-=�����﹕�ꤒ�o쨕����3m-�1i�RB|�x2��c�k��U���k$�(C}g�� @�.�QUt���\9�]�aUP�ä;JYp�G�V].�M֭M�5�A�R��M��V�S�,}���^^C���yyz����o�~�j^��S16��q�"�Y�y��u�t�}RM��V^��N���L���g�(#��JMǘd��1}G���v����N�[�nmh��CTUT[0m����Z�o1v*"�%Y{,�#��sS����+x�
�-�F����F�xC�Ku_O����E�ϥi��4��{�s]ڤdy��h�[u�3�ۧM\�ܟ5���tvn���k�8ݚ�no�FОc����=���,'�7�2��vط�r���05�p�(7iQyñ��a�Q�Eơv�����%�0^מ[���_� �`c.��)���wtn%p.Xϲ��f�{cn���0p.�&����r-�5��Ia�{�ym�H�?G��`��."� �5ƻW�(:ru��������t�y(�|3�����|Ws��k�*�����9G�������T�����n�\�s>q`,��ؕ�n�Yz�Իuh�F:�u���>�ȿ+��z���6�tS-��+WzF��q6����5����6�
�����.א��e[L�E��h����2�&
���7<8�4|<8�44j}�%uԦ:ñהg,�i��1_f��������)����ܝ\+:^����+냎88ノ8�g:�;�<��.����}#rܜ2E���F=Fk8~����f����G�^u#s��ڷٞAv�7A�Cm$�Ceh�u�?>0}��n)���F�s�{�r��DHx��k���s���Y0��!3�6@���1�ay�[�޾��+5cC�{0 )�N7��QӀl��!*�n�3��:p�-I��z��Wȓ�}KXs\��$�_)�7�MZ�uw#���a;����^�m[l���3�ˌ��ZC����F�{G˧n�жh�f���;����������g[�t�c|G��ot��7��
�����_g��d���#6p-��N���w�_rƞ� ��ahC��cr\'�[�Jx�g�F�Ѣh[����2�p��_F%��g=�C��(~�l�y�����;�/|�d]3��#�I�}a�=�z~H����>���俒��Us�k��'����F���KF�X�̧��6Zm]�x���9�;O��}v<b�ˠ�辖�n��F��T�-J�l���Σq�q;�c͑�lW�sC��^I�6��^J�?���C����^^C��������}1z��SjOސv<����a<n%��I�o���ff��Q��	];,�r:6�ffn�{�r8UZ�r���0i��,�v7��Q硛���s�����,��	���V�Z���s��5�`v$��W�Ei�\��jiԁC��]fr�(���"�AK3�z�;��f""=lB�P�q2���W���c�7����)�kf�s��թk!�}��}�27��O$�s��I�\u���������"_>�
��af���m�c�ܞgʍ�}�!�{�I$	 ���Oޠ��:c�� ^�;�<`Q����H�p�n�ޖ�"�[$k��\TEPf8�r�P��C0Ţ���$V�f����(f�c50�;�I�kR��,�V?f�dw9����{D*�j-��1�b�өG.�$�+�ؗWd�?-s۶��|��e�wռ�5$����]���I���@&{I��D �l/�NY,s�+�oQ�������Up�nA��z�M�����u[�I�f��~� k�F�����}>��������?�����KQ����~	Ks;�϶=-)Fy�[w��`ˋ�7
�aa���>�f\���HH�fÁӆ>�;���?ߢ��}���W���F�o�ft]�_[�~���7_�I07���{�jaQ��4�m�2E�p�~G��>����lD�|��$��m{�l�<M�����O��HI���j�_��0�i<�<h�����L,�Җ?�&΅����5��O�(X؎᪹=l<�MP��]7�UD5�C�l*�t[35����Z�S�v��z	�O�g�3(�Юv#��N��b�} L���7�&���n�ױ���8+��}�k�a��e�a=��Pu���ۥʃ�Gm`��S���{;ړ�>���>�y��lE\�YD����a0jQ��j--nY�FȚ�9$ְY��,*#]��sk]��&%��F�7q˖�)��k��*��#-��]�T������l�{�\L���릶�����1�%^���s����;�d+���pq�py��<�7���9�Wѕ�kt�鎓��7*�A�.FN��&�p��v�����G;G%39���u-��n��6+scr��� �[�rl79M��ݛz3q
�W��꓾��u��>7�q�x�U]��3ǟ:\aj�� 4ۣ�E��ow���f��ɷ@�c��1a��@����4z�j
��s=^��^��/��H<���j�}^#q��<�YVcw5rG`�?�����~�KwA�v�C��k��k�Ǝ�YaV���x{�-�ݙ�Z�ߗVt�?�H��FV*��i��{��ǲ��; �=��*~9�{_��#�y���WS������e�k�GZ�<�ئ�/�t}z`�f��~l�q���ó�2wd�ܚkV�}7���]�H���0��NǙ�6�Ӿ�u�X����n����~�%^�Rښ,maݫ9{c_4'��/�����5�u1$�u�wߕ&�}�gc75��v)'{���zԿOJAX��r��@p���W��w�7��-l�x�^���L���1�Q��- �k7v��.rC�e���5Re�^�u�)��@��Ly
����U��X�뻸�����m����6�pjKOQɓ��˛���8��4?zz��������^^E���Բ�U�."�	�:o}�8�(H%@�Z��!�=sY�Smi'�4n�E�$�����*~��K��k�{��m�G����N�F�����N�DS��.\�EO����=�q�s�=��?>�j:�[�v��$�����x�L�|��>q�}��o�D��E6u}�4f��`��� �s��$�r�P|����l�P������Q�١<��>\�,�f>+�qT�I �6߯hk�[>� ?l��{.�N���hc^�CD��}�<��bFJͦ�Ӈ�|��f�4ߣm����pq����㺼��|���l�%�t��z�u��r��r�������z�=�����dWa�W�*��oN������vj���_�W��g�4#ͩ
_wp�:29���PG�ѝ�맊��ۼ�V�$/!l�,�X��,�q뵦8rg�xMo;Ȯ���j���qՀ��ys%����n�G���r»��k���S[�-#%���n��$�no�誅���)��}V��ˌ��2��j��!|�5+��/��6k��U�v`.�ZЭ���Q
�F=�T���v��z�PQy�p/@�o�_�Y�*�������P�ِK���b�Wj��]WV��k�(�V3f���z��r�h�^bĢ�WyQ��]��,ꭤk�Cr`"��ĵ��R�,sd�Ǐ%j��8\B���N[���n-K��ell��Բ�X�t�Z�򇷶Q���S{\�ܬ��Ek�Wݩu�չ+����l۹���}c���qɦ3�=W/	�.��Y��껵_D;ғ�g{4K�<#rc��le�|�'l-AH㊭�H�
�PQ:o<t��䎊K�<�[6�c7r��k	�x�U���ˉ��B�S�͉ѹ��k��ǳMc9=�z�Bb\g4���K�X5�\o��Wg�^ؤ��u �H�f�}6.���t�&w�e��Q�16��]A;y�qL<-�0ݼN�!#����oje!*:#�v���B���	x��ᦜ�|�'Km�4��a��P]���i�߷���9�ϝ��'dJd=����aߡ�]l�J�vG�R�B!r��P�\�[��j�͜o��C��Y"!���\C�p���܋:b����
��T`��P)��W\��Cyٝ	˪�m}��j�9MQ���a]��wX����2>�펫͉����/�l[��3BJ
����ë�����b���lDvA�[�6.^[�ii���;�}-Z[SKǭv���	�܏�k�Ք�X�J��]��UXh�z3,��X;O�s�Ǒ꒱�A o�mi�r[��[�WqD�wh|���ΐ�%W�d�;sZ�3�Ib$�4��K]�.��+�%��C�����{v��Q&⠳�TuْK#1#��$�r3����L��Q2����X����E�Ȧ���ېխs:�+��į�f��ݒsL��R�hjۓ���f)�����s�s��n�G�u���a�)>��j%-��`����Qֵ�i�ø䩐��eأ���6EǝL[/��龘�u����?��ړ�u�ȧ��E9�~8l�� � �@�IH���E*�W�*����}����ƽ5���Zֵ�Ƶ�u�k^5�]}u��;d�y�3�$�ޒDϪ�r-Xr��H+$���!�^<u�|z|}}xֵ�k�k]kZ׍u�_]}{�ߓ��UW�(��
;���W.��KR(�?�޷o7��~��澼kZֵ�ֵ���kƺ믻��|�0��R#�\�W.U�>�
dr��	ݡ�;'�׏}}{|{k�kZֿֵֵ�x�]u��ף���I$!	GeQ?P�aEE���z��=".U^<z��*��TDA����QGĔQ��.�D��wR��Q�*���C���E�N��PQ�m���y�&ϸ���������K�T|��∃����"��+(��֙�C$�|mO�~��54vd���_Z������B%��2�$s��غ7)�5D!�d{���w�R��/�|������<��������?<߶}�*N[�-�vٙ���U�Xu�7��fh���>+�aDާ������	����g8��)�S����@������4� ;�/e���9�]�� =��K݀l��k2Ox�%N����q2��4vL�k�3Wu{�F��F{;���Rh�=��A6*u�K;�[�E�I!y13�!�G&�2(���
���z4YЅE�ς�(��|��I�6@������8k����1��U��x��f���q�� Oq2���uU�y}~��vefb��;����:���/\fe�j~�9�j�R\bt��	V��w�n������C������r/�;t�9:�̮#���y��jN�Un�������.�a2b�Vg#�;�>e8����5˷��c�8��r]��prNS�_]�kT	��}��#�f�g�zQw�N�H��vz�ӹ�I,*x��9 5� ���,��5���3�q�R��ƹ�O��nv�������B�*�ɁIA����^7u.�Y��m~���!���<����󁎚R�K@�z���t�Ɇ���(���4�[{�җim�}�8af1YyI���NN�G�c:?�O���,}}�z�#�31}�Z������;e�X�+���2��D���C���M�3���u���7'���8�A,2�{v��P�[8�o���[�`��m�T�e�i��퇯I��0f��2�'��Ʃ��V���:�f30�N��$�5����Ot���u9iH͍��;�ٚ�(�b����Ԡcy��C*6�t}����[>��؆�C��A|�\
���t��6��I��{�����v�y� ����@F����{�66����zD���'�ы��� ;�aP^0{��r�z晃	NZez����Y	*��w�4j7)��y����	ګ��c�ܼ2*�����~��>W�U;צ�+���f�ٹ#z&u�I�S���Zv�=N�)a'�,$�Z;[���<�UīT+�-��P=� 4����I���qʕ.^i��_VJ��>��w����^^C���������.��.e\b�y�����ET�Xqd]3�7q����T�;��\�u�zC���Ua8Q�����\j	�ʅ��p]Q��n%�3�=������x�54�T�xR�q(��Ri��V�{,t00Jf�񙋱,��Ԝ�xz����FꑻFN�eļ�w��.����V�[��5#��L�n/FڏVv�>O�ù\^�5�0B=��/�=��Sf3C�*@]O�DKf�Z���G���d�� /5��y���*
-���q?˹��[=� ��E��f��#�C�b��?�k�n1��ny��^e%���6E��`\8�H��}����6�=׸os���W^��ڔS�|��� 	�4o�]�6H��*cSPw��Mu��w���t՞���k�<�i)n��>A����bh�)�L��W�s�,�I	�~V���@8cqtM���V��R��j}�����MPVo��PCp��B��y�/ntv�J��r��:�`tzK���S���V�h���*v�u[eN�刳Օ�����3g7�W���Ulw�%ǜ�;��y�^FA�u�n�y5'lS�Ҫ�F��N��G^b\��ѭ�if�;"�7�-�|���m��I��8��8�l�X�mv�x�8p�Y�ǖOK��d�QO��n�d-ޞ�M�k5�,�F��u�b�k?�١מj�>a�������������n�:hճ�P��+B��9�`l���TH�@�]����E�uN���iT!8m��楻w���R�+�q�k�̹}^�	�H��gY�LG^�K4��oso\�&�
�<�FwAp`��������3��^�����x	ln�奆W�֊�v��y����Cz����d��^JW����//��S��P.�f�n=>�g3�A&c~�������A�e�4�c�k8骏j����w�M�H�����
5���i�6��6�39)��|;�H� �<������[�+�[��:�	m�{`���8I�O?�e��_�׎�WX���z.�fϟ��]�X��&���V��QQ�X�xdA�����\�*�)���i��ZMu��*�ԝ�?`I�6<�c�|�	ǻDC��U����'bު����_`��/9T����z�ߞ\΍�������<qq������﫾����0�#����*t	ۀ��~�-$ l�@�a���e�=�7��kw���@��Le%�+�Q�;=��d玬�Z`�=�j�K��d[BP<E�l�Q`gd{ʣ�ɢ]��w	�끻�H4�7րc�4W�n��17G6)h��w֞�j�f�t�6����^��G֫�@��$��x#:ut_�C���קk��W�6�e��R0c��������\�l���+z�J�C9"�<�Ӏ?�/7�^Is�c�����g�eK��GJZ&��>�Y����7�g���q�x7�`����8��x�u�D�T	ݝ�j��!���>�W-�V�8�W�E3�ĺ���fOv�7���>��#�2��ّ��ue��u�F^�o�g���Y}�Ww.Q��C�V����HY͹��.�ד���w;߉7k��2 '�� ,���a���c�U��y�Yb��H�m*���U�����b������Zu{�y�=zq��q����d�{BG�d�����1�� �$��OC�7���~��%���Uoef)T5��w�D������/M������xp��+�.��m;ҽ���-��D;0v����������	r�eV��&���-�qȓ���邢����.����*zBI_���z�Rc��]=�:{cW���T�=�<s����CO������
�={�{��r�'p
@/p�ng4�9�f�uҤW(��P9Z���7��i�������MϹ�@�7}��ȸ�᭫|���~~j�e��,2j_�ӓZ�[�I�pfk��i�����0z�[u7�*&k7���8�S��������6MVNҟf��"�#�C�V̬Z�3yX�� ��h	R�b�/N����k��fƗ4�ߗ�*�;2���y���ެ�֯fdL��*e�%��B)��s�j����Ԋ88D�J��לoM�L���[҇�Q_V�weG�q���G�3���h�}�i�j��[��m�S���Ι|Iզ������u��]u��q��_��su�����k�"�������M�W)}�џU�\�=y�q���o�Oo�z�4��M����C�**'Mv�˩�nK�elS[]];����;��>u�Dw���0V,�5�&N�f����:56n�ʸ��%v�>����f�wP��Kn�@rY'
�	5�yw���-f��,�!�U{lF�oz+�=oTr���h��7��K��G����mG����`,l@A7��\O0��Ӽz�duJøkd��K�@�`�<y�E��g�_)H��H/�{|�+w���U����Q�������~�}�-N� {|��qR�(Qf�P[/���Zq�3�`��ͣj*��Ӱe8��\��'tT�|�����V�u�zw��"}�1����4���N�^�A�nD
x���{�9���LĆf�*C3%�WU����mǮ:�<c�)wP��!5Y�]�rR~�)i��0NL]�^�m��U䫑���w}�7-�X�<d�}�����#�hOGܡEG(���ص��#���wm��O�Y���gɂ��#��z{�z���'�){�rO��Y��o_'�F�&��;9Ҫ9¦9\H�:cI\��C�\�O&��r��ϝ��L��ۋ�88�c�>g<�Ė���������p�1���8��֡���!5�fEζ����;��
���^�˼Mq�oB��@�ku
l}cF?��ٻ��L�F�A�~_1?ߘ�6���銳23��ftW�*��+���Z�qCZ.�svۖ�_��0��}�8w��W�P`{P2�ܨʜ9z͂$�S�:I'��U�ny�wG;�Ȓ�W,�m�Qf,��J����F}�
Pd-��0f��|M���Q���]nd����������]�$�i�[E����z�N�� ʳ�z�Ϸӣ#��h��LmWnmd�ܹ��i�n�~�n
������	��~�^�f��p�3ߴO1�׉��\�s���TV'�P	%��D���|va�ã�>��5��H�~�N`y�;(.��;�yl�"U�+˘�+�wV��')ЗՌj[کnN�����4ʑr�"���gK��ixa���t�_��>]ݶ���S#���kb�[�9�U[֢8�>�0��|�oZ�R'z�
���v�����8ノ88��/��,���|����	�[Mz���
q\��u�C��%�W&��9��U<
�픮UF�#WH[��3Oi�pU�^�Ռ��Z���TE�К8x⥎���_��rdϜ򭦿d���%yă�߿7D��%�<�s���aH���'abIH����o23��RX'�������6�VyTj�cPr��'^�s�(1~m]9��h���nx��fh����VE�cz�P��ff ���p�z{�U�vg/"��+yCs588���P�͐\0��zj�:�c ����SYA��b�
k�{qT�w+�	g�gY��������➌�ͫ�̞u�/vSܼ[<��@��_�*����=Cj=��P6/�z�8�Ƴ��t�.x��4�r<�ݍ����0e�V�_Ɵ���SŇ�X���p��l�+����G&�G����169~/SBT�5�QJ��������3��cD�s�+��5��IM[�7�p�N���}bWj_+F[F԰�*�O#ٷ�Ϝ�?D��.8��.8�����˩P#w˄o	O���3���� ��jz��c����;l�ⵘ&g5֧+Ъ3͑t�s�wɴ���Q�*�;vwY#o�wf|��Y9�ކ뙅�t+5&��<^���똳��Ŭ���J;z�Qm9�}� W�g�fv��P�&[!E���q�2��tӋ��O �� ��*�����l�����^r�r�;:��Z��*�<����Ub�j�e�c����#��G��8�^*��!���}��(�B%"B%�͏��⯅�n�%B
�m܍�S��wY8K�9[���`�^�6��	���:�dY� �zz�K�Ƕ5�lZ����X�P�*��ff=޸"}���-��^K��{��w��.�\nq�@5iY�g|�Ƹ`"�k[ڢx��YK������������S5����\��.�ec˧�9��gI�L;<��1�Od�`յwG8���u�e`.t�gM��6�ۓx\��^�]�L�c�*�B����4�5� 9k�c��r��Wz�n��2&`v��)r�pt3D�2T�U�w�s쳸��ӛZ�H�t�<�6:g��\���nf�Tu�x��Ǻ���£����o�;*�N\VN���*s����qWU�;m['3>[��l$3�9%�71,�Ya���|v�킗6�wt�:�`6�b��x��i!^:[�0M�t��^�nQ��Y�k�'h�uLj����ñΦ�ඝ��U��F�;V��ɇs:�|��{	x�L:/������Wdʥ�`J
C�5s76��96L��,���0!��1�F����:�<��3�!�SF#�b8�'v�Cp�sF-�kgi�|��%S��!�U]�γ�������-��}�[+�;핬[}�.�YQ��j�G�:���宨��	��'Wj�M�p�r�pEEPA��������nL�Nu�R{NK�<�V�9���U� A�h��G*�n���o4���m�WB"'�BWWB�O��#Cl�-�2��S8wՌ�0ޫg◳�?U#kp[!7�h$�^9HSҴL����i:�q�X�8CH(8K.k�K4���eQ����|pU��d:��y�1ӗ6�6�!(�M��Ǎ\��m�v��3����+f����g��a^������CD���� PK���b�4Iɲ�m�.ity8��o;A�ƛ�뺧6��.;�ba�:�r>�.�'��[�x*!erᤌnk�ͧ5;�v��;��U�o�hu5�V�Z�>��ؔ���Fy�Z�8�
+ȰY�ơ75�wv�`@����7g#��Vdz1fWCyc2��`�m����a�{P�LhOߖ�dГ����ը�k��,�����M	�+kwf%V��m}G�+�,��xi���e�T�vf���n�^�I�}z�4����1e����.�]��n��!���ސؔSR��s���x��I]�B�ס�m�47%�u{��]]�\$�(��9�kq]o6�mI�L�Z�r���-4��k^)���I�IS,z��\z��8b�x�Х�q�»���o<Z���˱:rtV銯;���:�Bm�0����!t�9����°�}�j�1vGB�Ϋ	��3�=�Ue��+&f�]Fi����=5
�V��rH«k\�Tn��sxռ��H��.��٨���m]�S)�OAH�������G�rhO	 �I� �H'�P��D��B=��_��Zݿ���_�o��ֵ�~5�k�kZ�]u�__[�䄱��c��3d�f95Si��(���ON�ַo��������ֵ�k�Z׍kZ�]�o7����o��C$}�r���
����s�;�'zݭ���������Ƶ�kZ�ֵ�Zֵ�]wy�o��|����;���)�t$�r�B�8�kZ����Zֵ�zkZ�kZ뮺�����#�AU�w��!��x�_�(s{ITEAy��I9ҹA�exr�z�'��:NC��q2(��8QI=�սD�Q�t�D��G��2.U.r��oi�"#�x�w�%ޙ㋬��*�L���ȎW�+�}2"/E��*��>�*#��r��UuJ�3��
:4�1�11�$I!r"*)H�F$�&�r�P�Az(�#�`�2ϙ�m��*̀����|�rY�-�	�B2(�&L��E�Ya �d6��\���T	~��$Щ��K:ڲ;���
������I6���Ө��4�ȼ���������6
<܁�hڞB#⮡��K�2����$@JbHd��.(�aB$(Al��lu�=���D�y�;�<(���$"p%�!A!	�#QBP$�R~1���!H��#U�F
��}�@Y���*�l�}"��ry8����ŕ	�&p6����眅�d
Rp�&"R34P.J�#l2�d��D�����<�4���߷��5�mkC����>�d�7�e���䒨�
	��aI��)�5�jɷ�; <`��O��[d�6��xq��[�qU]�\��:b��e`�8l��r3s2F���DW��.�&URwb�R�J�S�������}/�C?����	$��k~�ѽ�E\��[|4ϦFS�����W��=��<uzv|�xbU�Ң��/g�tۻEWD({[��L��T��+�o�n6���0��nΝu�\`[�}�j�_�W+�(��ޭ�=0K?����ߛ�M��N�����Q�r�{�qq�R���O�]Q�/Rn�:���O]Wdǚ.Y��`	���J�:}��Mu�;F��4m͍�PU�>\�C�l���������/5�vT��!5�Vl�˲ꏳ��Da���쿴�L!*����Q���dnL���{�������i�T]{Dv�T^󛋴�����l����'=��������~���B~��m�`�{:_ɺrg�v�ռ���ԩ��Q�����\�p�6�op�(N����+�Ȉ��N����+�y���,r���%=O1i���K�X!���r_k�1�Qӎc���o�v�<��l��8�xf��ִ~����0c����{��q޹~�t{�_�9��}��Fŀs��6�5�j&j�$r_ڎM�S��8C��7����Z6�ף}]�eTS��}f��kQ����[W�򑫹z�A�������<��y�x����[R���6�^0A�L%f<��K�q�ٙ��c{8:`�=`W<=�@M=7O�x�wY�K�褦��q�{g��ofZ��$��f����1�0�w����6��~���x�����>��	8�з�������oʖ�ӳ7�z��"ER�pZ�a��<[�s1���-��V��H�j�h�w�����O�s�5�4-z�d���y�,��q2"=�1�����|�Oy1�xg�Y���7��Ƕ��#z�\����Ϙ>��5��F:\u�MR��kX�,�bos��u���H���BEU�a�����dv~��V'x�u}��m����}��[XO{�Y�����P�o����x?h����m][/Q�0ڭ0��/xC�!G���@1Tu%��%Ê���Df����9��oS���Uw%Z�����	̩;�ӝ��o}p�\`�b�g\��;��׼7z�&��$�}�o�^&g�]��wlol�-�dp9���u=Tks9h�d�.��[���oയ�=�1';mI�a�q�Ym��O�o�߯�=��л�I�H��=�;�Q���>p�2xȷܽǧ��ʲׇ�m�c�Af���E����/rں���p+���E(EM�#�X�xfw�yͬ�V�j:�3�p��Mz�ܳ�^>�
\����Γ�U�fW�cz�Ti��۹3M�j����Uӂ�'�j���H�����:=8��Qx�To��+�r�l�cnWI�F�B�9
���8�����̒W���k�U�y�Tw�ż��-�yڸ����f^�
!��@%���d�vh�#Ƿ֗b���/{�V^W�4�A>��@UٔpΉ�5�5t�7s7Hl�~�ǝ�J��۸�t;7��G�89���T��Ӷ��RI�2J_JV���ι�����{�$�c�~A�=�[��uɡ+9�f�D쾬�(���������������W}�Խo]0�X��X��V��y>g�y��2m�˺[ϸd6�a}�>��� ��ـ:6c8��3�|��$����]������i�^r��=6�����w��f���B�Y����oTz��ج����� �o����9�k;M��]���7�ґ��۹�Ʈw"��c���'ν�y�͈ЪUܵ����H%�񩨤&"z��m��l��Z�g�p�Q玥Q|��f|�lI0���Hk���\a^�㳽t��ڳT�bT�,OA% ��@Q:�|��FHb�����@^���-��q\�ίʯ�"vk#��^�8'r}��� j7a�Ɣ9�OT��:fj.'�m�^CV�(���fs��w�J��7�p]1���b�^��͹���̖��V�/J�`8��V��� ��`�#���)�M����k�[�:<Uۚ��}����k�a��oURK�r�����`��PɑX�x�wY^�QE��~�gf�޺y���^ɬbMLZ��������RA��pM��Uf��d��Q����?{|G����o0��Njd7U�T��
���y2���qvR�N��Ž�R_.u�r��}/&��PG���Aj.��ٷy�:ی�	#�[p����s��|�]�վ��PT	[w�30��~y��Iƅ��5w�(�@��O(��>�ޣ���5�B��kIj;�7�F�9���J�1��ңӾ����̛���l0 u��yi��%S���l�nj���������7M��w�y�0 2�:y/0�4(�h?j!}=�^�`7�{����6�F`n5?��߈�����{�ådJ7��zގ�3���g��+���F�v�m�4��̘[�p�J$�v�xϣ=��DL=�H�ۇ�Ϫ�荒i5ˮ�P쯭~��p����!��q[��@?d5�H�7r1�n�g�,�;1�����.XU�Wg�މ����\V{��dFk��\p|B�s�ѱ���~�>�a"�K8H���;�.�v��.��E�7���i1�Ŧ�3k�΃�Qszr����3�^�ݓ�#e��n�u����/�"�|Ǚ��6âS���O��t����^q��Zl�5��R(ļW7�rf��|���w���E���'�6��Z{�G����> x7��+�J���]���E� Hs`�N��8��u=�OQ�q���O~�C����*��o@�"�hǲ��p�I
;W�wmel<K����:���>y������~�*�6��F�d��n"ĵ�D�a9�=����0,����������Z��&����n{�����l��F��[�kl�G�חV��u𿛒����UN���F�g-5Z�o�A:ff5����M\9�W��}���� Uz�^�wjƺ])��FX�����w����Z��)��O���[?g��~�ψ�5� �}����z�<�� �xzA�)F�Dlu�z|Py�7�\��ׄ��W�nK34G��?��_ۓ�M{�V�i���Nw6�����q�;��m�\޸�ç��CE8��!Ր�����B�Ev\�%����,ωD<*��,���[j���<�_iN�^�ir7#���uok`K�'4Cj���+�ϾՓ�@�Q�����ɪU��B��eLH����7�
.��O¦��c�e�Y����٤�<�[�:������߾���Χ�^���YQ�3�LUxZ�������>M���Л�Xgӝ�w�&1���&��D��lܗ��4��{�jz|��{��Z[q�*��|�~�3��͝}��#�}d��㵅�4�=yR5�|��a̐�t{
'N% �Q����h�yjQ�Q���5�&��[$���w�{�=�@���ZzE���B�'�� %�%����d���V������oU�Գ�&1��`'�V�쇤�ۦ,S(���5�o�8^�B��Ԗ�����;�G)_]��r�.\�-��2�Y��������m�Xs35�'NT�uz���E���-���7�����$���}�_��p��D���->����^w+��e9�=Yun�-��';tD��:Oo���4�4��o=7.#��c!�nNP��1$nCU��]+�e���W��jmy���_�H�ꤺ�=Q�v%�e��{[�;ݔ�Sd���q꫔k��\<r�v:�6��5+�:Pʹz�T�х/w�{�L�4��������\b̽H���W���K��@��\y[ J�C_7�[����RMc��p_�:`��L�����-;*|������8�^�ٛ���j�M�.6��Z�7L����u�pd>�UNg��_�Gf�a�L�L֋~y�=���J����Cۡ/��6|�� 6k�Q|[t3���ft�궓&�i.t=�c��)�oo��T4���?G��!�H�U1��G�;���V�R�q��x���1*t�'+:u$��r"$C�z�ϳ~���v�J�Nsʣ�/��`��G�DH�;U��C�8��Ek33�U��_ ��
دp3��/����x\�{�w�u�SW��z�oOh�h�h���P�\z�T���^t�$_Eom�=E����@,��S��Ϣ��J�o��l�tz��kFE?�iRY�e���[+h���]5_U���%�����K��r�`0fUN���:<�ݿ;׳��l��`d�$��$
>e�o#��K"�o�/�ҋ���d����oNL��rC 1�j���ކ�ޞ#���>>����&}�S����+>��t;��Νڵ���.��ӷ�Sw����㢲��NNr���Z���!i��}��/b�s������t�N$&��^'�7�&\��U�^``���85;"��q�߅��󨙃w��������4ݿ�!"r;�,V \���^y��L!��Tj{���}�Nڣ�^��P�=�ས{vU?���ee��&*�1�3"���,P~�Y���oo�#��[��B ]�\�Ç�_D����K�&ٝ�� D�M�d��Q�3Y>C���ĴAS҂��e2k��*3pZKS��S(��T�n���'��N�XkL\WgF�\����X�QZh����1��ucw���w�#}�զ�Wǽڥ��_R�|�Wp�6O������Q�6e�8�qÏ��\>+����_~�/�����4Yl�I`Dez��X�_`�O��f�#u���3 �7���kw���y��k�V�X@���J��Ag@
[m��_�i�V�n�^V�Z�2��u!��h�.�{��7�eҸ˸�V��v_Eq�l̾ʨ���Z��+p����f�����vr��y����D5�ԛ�)Y�㾙Y��7ü�K�~gЌ0c0���j�+_9�ou:��d��]Nfk�~�v�R��U�Kw�1;]��ۉ� {��D��DnW{��u� ���@̀�/8M���k�����V��;+3)˽M��\�\��æ�:�ǫ�9eJf2��ޞ�k���[�6�2c�z��P`^g�5����T϶z�6�>�o@�������|�tLl�\����B�=nn��wr���O<��a�r�T#�������}َ/��D�뱚{|�'��3vU.��tD˄���W$��9���z&�WB;��:�����~��qg9U� ������ÿ]<Ș�|o���i;���p甚h���$|k�5�?}Uz��F�'x׏�B��X~���J�s��ު�O�[����*���K� ;���M�]a�i�Lm=�λp�w�n�6�2�ph=g��!f�M���#"-\7u	����v�o��k���+����[\���!c4�9qgJ���}���	*�NV�uh�X���:旆��wb<(��k*GN��`�E�0�Y�B(]��]����˲kW:�
=��`�Cq��s.��>;7''f�a�|ϝ?Q�λyn��}�4vrس2���vG{��j[R��h`��G�u��XU��˳�{O]�m�Wb�p*�p�1�x��"q�vS���w�u%���:�|h�_�'��%��&+ Hܫ�aȕ�N�dՉ�\�v>���v�`��g��Y�U�Ȇ�qŘrm��%��\<��κ8�Z2�d.�ujY3�iWS�ޱ��iq�i���z���1m��0j�TYy���5u�S�6.��c�ɋ��Zs���0��1O������|�߸״X<�
�w��R��"Ť="�r���;�q�������v��-T�Om%�s.��KU.<�:y�5�o��^5wl�����Α�4/�M�ag��p~̻G��p[�bG���tF��Z�wFn��5D����F�FR7<�R�lS�l�@OmHOm�~�N"
�y`�)
]�[=nWo�;Y�7�/ˎ�7sU��K��;�@�������l����\��r��t�sǝJ*��c�BNw�9��-Α�fZ�L�*��G^t�����t�iWr��9�<u�bpqi�����!��R"��p��d�p�j(n��]�k�or�2�Q�d�z6�\���R�;����Y��՜�E	$���I���]�m�M֓��-�䲑��sR����0Ў�|mt$89�K�`�ݣ�j�,R�ݛr���ǅ�"������a��FN��V
�S3w�M����{q�U;3��c�e�qá<��R��fQ�)�ZUvNj�K�w%pnPP�
�ރ�WizћT���&c#�̧צ3�ei���'պֵS�J�t�����R�գj,M����R�u��7Q���$����<q9H��p�o�ΓgLػwSp�|�����W�����Up躖8X�=x��E�R�:��ل�&I�N��^]g-���;�]{�gvB�L��ȫ`���S�R�{��M�P\�:*�pB2���)¥Y�<|����9G|c�G
�s�r#���OM��!��Ǐ}}|k_Xֵ�k^�ּkZֺ뮺�נ���9��ӷ��rNo:��?�GՐ�!��'�ǒ�I8x�:�kZ���5�kZצ��ֵ��뮿w�����~�rs�'gs�U�+���"�Q��fǎ<}}}}}}|}cZֵ�k�Z�Zֵ�]u־��$�L$�L�K���^^e���#�VE��u3�e�_�N=��X��g[���������ֵ�k^��ֵ��뮵�B��<��I$���y��j�h]����§؜�H�᭢�'�{������+�8�&�Ao&\��a$�.Eq��E�^nIS�A�T\*�j�U�(�]P3P)L��Xym9h��Ȉ��$*rJ ��r���ME�= r�^�w�AW�~0 �����$>���V歽���Gn)Y�33�W%�yn�02�W뻞�Wc�=���ӯ������n������������x3y��>��ؚ�fx�����Ȭ���v����q4��§�;��ۺ�DnGQW�K����8����Clﺂ����5��Ϡ�!���M��L;��̀�0�Z|}O}�ٺ��-sd���q'�Cnn*ZM���y�>�^�C�bô<unݰ=ԫu����Mu�0��[Jƞ�̧�������0<a��B��ٴ���.��%5��3�G���͖�_�ڶa�)���v7��Z�r��]V���y�v9ݓg}״l�L:/�3����mZ�f�gp�XY���W�Ւ�g(���P1��Y|^1�ު����9fxqo��2���b畱���6s���Yه�٬�e^��tG=\��nM-���o~����|�|�ϸW�h�xv|�	j�JK����J�x��w�lޅN3:*�+����gau���w��Ʊ�-X5Î��{f�Om�p��m��vk{�r��Qe"X!�������Gi�So�L�_'|����`G���$`��j�Qu�_�״��������WR�?��Ş�OhÎYx�N�j't-[�0����"��w����/s&��
��h�nY/J��VB�5f����!�L�7���3�������`����,�O������z��d5�}���Տ���2+�B��ԵG��6�n٣��T�Mq)鮤�]w#oKγc�*��/yH<S��*��햿s�6� �A�ڭ��Ҷ{�	��s�������V^w��1�ws5�I7���c:t����4���h�e���c�j��Gf�Qw��#a5���O.���O�W�xfk��yUժ�-�0{�� l�����j� A��]pN��ao���WiJ�z�e�	ⰭZ�)�8s��)KvU�v��<��Wpp&ݶ�s�K�A�z�z鱄,R��zZ���e;Ѷл�*���d�:�w@����b�!"���!�RdP��HUd��zX�X�<��GtacU=�]^���Kr@�F�G�1[t��$����۝d��]�I�}`F1�`�O��W�]ddۯ�5��IY�$��K�{}ܰݼ:c"�����f��;7̄������ڿ�;��oM�z�N��9/8m����ae�Vף9�wf�J�O'��t	��Z������t6ɍt��z{{����q�8ځ(S}����c�w5#ź�9�u��k�Ј
���������.��NQf~��H\�;]O�ڶ$�D晐Ľ
�!�q�p���z9Ո��t������ݰ�<xtu�<gctK�UET�X�Bz���+2�f��! C��rؚ��7��C<�]KbxW�1Izmc\��3��M���eFNw_��i��bV��́U���ܩ��l����7��i'���u��(u��W �V�f�%\��y5m�}�nɸ�{���,$
!�"�g׋�S��W�`P�3��ս�,`ՠ��Dd��a,)���n������>\�`��'��%G����U�xŔ�"�6���"�8kn9u�`T��{�*�|{� �����c>�s�b���WG�F�x��0���=9��Pi��J0��&��q�ft妆����B=<y1���W]��p7s+&'�Ը��ѻ| ��x��o7�y��(R$�*��
����V�7�.:�\]K��h�ڢz=u���Kv�j
���4�l�	s{d�2����-îm��n4Z�a��3���h��1*�̻��/�p��}ٳ�Ԗ�[Ϩ��	��
��iZ�0=�P��]�*��!v�������!�	[u�g#�}�ϊn��rn(�n���>wۤ�7��)�"e�ݼ�f�n�RDL���^!��hn#{Qs�0
�����]�3~U�� ]A��h薫v����e흛��{�v�UO�����o{���b���)_����լ*��v�56G=��l�ᨘއ�;9����xd�����*k5YڻX5�z�n���đ�d燁�?���, �j����y�J�հ����9]�E����f�z��g-��z�څ�od���K�<��"g$vraך��Y�-�MZ���<��d�Ds�q�,k��깡�Y��"���V���W\w�&w]�#���+�WQC��6��r��J}�S�Vn�/��i�� �3��޺�gE�f|���<�γ���B1�|�"J��g���4�4\F�᪉u�O��;d��)q���廰Mhל���t��[Lco����DEUP���y�wM��=os�n��ƈ&�Ӧw���eKî��PsO�9{:�+��h8Ȧ��znq#[��;�\:	��*��s�L%���ZS����������
�8e{w5Q]>����9��z|�ע���Wv�X[`u�f�FmWbT����W*��4�Ӭ������>����oQꎶ���w<�-2�q��譅#!f�wy��-s`5p\ c3%kF����`�V3�1�;=���j𾈺�6�-��g?E�77�j�Z]t��8�H��޾׿H�ne��܏f�+�����d��GF�][v���7�tyV@ܧ��/�z5%�4�m�ҍ��>��n3pd��p�`����f�gl�7r�
."ݮ�2��^��:�٢��2m������6�lv��H�:�$��,e�}is���d�����f���u�����g��y������M��ӫb���qO�ȇ0� ���M�L��WP P��h?WC'���}�nY���(���3��ěJ�d(�a>x�MHz��U�gi�x���R�\3��q$67�'���`�&$��t�M4��b�Vv��&Y�c����
m���*�IFq�L��ie�V��o̟�0�.:�p�
Y1C��ɩ��n�s{��_dJ��(���8ffj����2�k0(wXu캊�O�����8�Y�k`��|יv��v�tG{'t_�Z����G"�]O�3𧠕o�fYuGNb�Fs a������Wh���u{�x�xL�Y�].�׻���Җ�	�ۼ d�oU�G�\׹]��w��0�����oSxw��On4^�x{��Eݝ��3�gH�I�x�:�B��q���Z�/&L3���'�b+��I�l�Q7�OZ��i��[��Κ�#�or[c<H�<! �[�@�mU��ͨ\R�D*�Mn�ީ�p���Q�g�B-��5��oI��f�z�v�cO9�s����c �׹מ��m��ϸ�]�y���g�h�j#Ϝ�\��wIU��S `�;*J�Lk�}sGV�[�QL�G7��I�>�<�KU?G��^r2�w��8�3���i�\5Mg-6Ӳ�˖.>%+A�m��/�>��@�����ۭ�S�	��=�n��{�}��u��n�yKx�a���l�D��Mb+7��x3���H��ꬻͶ3���)zv?d<�-���j��l&Zy��c]���p}?0��ﾑ�������	���\��Ǉ�}ߗ����p;~pn��U��ص�����We�vFk��<޶�����'��F�/f�S��E��n�>�W�Y��V�¢d��3hkޏ[�FS?|a�Ћ�6.|e�K�Z�l�uSdż�üP�;g��A��ڙ�^���f������MYs*�X�����^z@'�gfA��0��<a��D����-n����Yt6(�Z�k��x����E�B}�iaV5�2�������{���r���6&%ќ�ȳ�N#Q}�2u����S���!=a��b"_=[�Y���G�����Z��W�l����|||��޺��G
��0�C�m0�\�>]"�	�R�̧k���{ �Y�-�)TK��tNYӘ�Aq�fzDt��>X��F�l��JBJƳ�ɋl0���ٚ�\���x��ˢ��(g����ˣ������/U��L�D���Jz�{��'Mr�3��軿e[�h� wtȅ9��s�ڋ�ӝ�[O�f�9����\]K32�So���|�W�!���h�w�{ڴ����&;N�m���dd%�o�8PT�ê�=)���'����3
O��$�zR�V%#g��%���1��1�Ȍ��/o��R��p#���T`T��lG�a�K�B[������۷�'�^m��B���W�x�37e����Dd�^��w>c{��8O�ı{Ӥ߾|�����=���)~��$�)�}I%~�B��*��Ѥ������������{��r�4�K��zƛ�5���X���<���4�I�d�o�K��S�HB��U}�����r��"(.A"�*�A��}��}�~�g��.�K7P��} ��֞�n^6��W@�r�1�w�e�;����x���s���%�g5Rԗs76��E?.��];�35�k��q��Ƕ�M�kLN��&��n՟���+>���=��,� ȿC_�}�P0}=j��cٛj���={{Ў�z���L��p�s���_kz]�������s� ^cr�O�iu��0�]�O�a��*7::^C�>���ϻ[�iB�T閼�����G_��,����o���	��h�����v��xun^�eё�۰�:�r�^���DU�A�������,�"����ㆊ�A��V�ܞ����3��W�A�aǯ��a	G�Ͷ�,�͓���:�33յ&
��U�Ս状~	����>;��N�߯�gU�
't�����dNȳq��9I�������~�("��~�����LH`ޠ'9M2[��a�!����k{����yT�����0<M��I�c1��\�>�7�}�W�}�׮S7V-�� �g��[��WY*�M��f�cz����k]��ʬ�\�©\Z*���&\S�(:v��I�s���㷹O,���5���o7�Z���Ԉ'Ԣ}����B�}~N�����lFh�-+]����H���L��1�h|�`矟ȝ����m3�6�-�;�q�kZ����s��ye��N�������>�<������b�X (�6�y�a����5�f>U��&���و��&Y�̯!�\{y�D�6f3t�??��[�vT�~��Y�����w �y7<�"<�G	��,�y]�Hu�}^v�`F��NV�Q����h5�V�9�
�ݶ�$o_c�n%:����=��n�e��,�`ǮQ�Ow�uR\�{��z��Us6-������x�^�q{^����,�K=�L2z/�y�N��i#��s�t������R9<TL�z:I<�hS�э͚�"v�3g�{���p4��ϟ7�������ۘ�� s�`����?����� ����'��a�l؃ӽ��`}@k9 ���#R221�E �����##B!�1����a2���#�#�L��@Ȇp���9E#����##H0���ș\�v�&S&0��+�1�##�20@ 1P�� ��@R!#H �1D��B �A Ń 1����D 1D��D"1D��C 0��T 0��B��B 0��HD 1��@��BD 1P��BD 0��BP�� 0@��D 1@��B��D 0P��BP 0P��B��B 1��BD 0����u��BA 1�� HP 1P��B��A 1��B H 0D�����`C a���d��B H 1����`0P��D 1��BEH 1��BD 0��B@A 0P��B HP 0��B@B 0@�� 1��BE 1��B 0��BE1 �UM�U  A�1UR �HE  T�0TR �EHE E\b��*�� < �0 �P   �0T �@ Q �1D� 0��@�@��"@(@�@�@@(s� x@�@�@�@�@�@d**
(��*Bb! b b�� ��d���(b�*A�"��@b� `)$�q�`2H X� �V��00e2�1�dC)� t�)��d\��9p&9�G; ��`L���r×�a29r3���g.\�3����������?��PT	PH� 1?��g��?wN�������a���q�0����0@�����������������J�������� _�x�P@U�/�����;?�?�_�O��jܪ�*����	��?���Aϡ��'a�/��D�@���!���$��a �@ ��Db! ��Q"!XE �H
A�A"X�E �P��XD � �H�D@���$b! `�*�B� �b�D�$ �@��
,�$���2*����EG"�H�*����`�D���FH�B"��X�D�H�E���
b! 	�@��@��Q��"!"!`	H A
HE�b	�A""U�&��	�������?��TI 	 	DI����s�_��������CA�9���p?����y��a���ω������S����U U�3�����?by_�TW���������?Q�(�/X�yB
�'�����-_���o����C�'Ñ������*�
�����?��g�C��w�U@i�������/���'����~���o����@�'���?�;��U@i�?��?����
���w����$L]���`v�ہ����������U U��IǷ���  �?_p8��x�\K�����/�``~?4Q����o����1ޟ�����)���\?���8(���1"__/�_T�Z�AM4�C*�54͙ATEmmU%��,�سI�R�T�QZ����IQ�2b���k6�¤��ڱUIl�V�)�����kU�ٴ�ٙmjٛJ�i�m�ma��-dKZJZ��H�kcfmh�6h�M�L�Hm�ZKV�jͫ6���v�e!m���)6�f�!�����Vٙ-b�L�m3Z�-Rԫ4֭)E��j��Q��ƦcX����U�l���Vٖڪ�����ͪ2�j�U���ꎳ@Z��<   n�z�[jRڒ�-JR흫kmKZn���J��]�4�5��X��m��ku��ƪ�Y��)J6ڎ�[JqM56[�5u����0wRѭ�VС��k-km�-�   ׸P�СH����J$P��С��OjV,�����j�,�����R�Vjb�ݪ�i[Y�-���[m9�\і��۰ݭl���ڵ�vM05�j�Rm-T��Cf�D��U����   ׀P^֭J:�ևY�کUQ�QE
�r�QE*���N��V�Œ�B���*����e"���nu�TJ�ٲ�l��[l�(*�T�0�   7���hҌJ��]�ݶ�TԲ�hU6v������ְ٦����\nJ�k;�⊒R��fb�'5m�f�4��H�kf3T��   ��%WZ�wuUU)��[�@���+�T2ݲ�І�eV��J껰����ڶi�۔WXn7"umATN��L�a��-�f�4f��  <�XoV�t��� Q�Y���9ҀR�9�� 	���`�CF�Nh(P΋�� 	��f�[,��J��J�5���  &�)TP�m�J
�۪� ����P ,���A�vr� 
,� *V�` jAn��
 wm�
 �3�(�mlm��V0C�  �xe@L� �6^nR��4ڮ�B��+1� �&�s�Ѡ��
��u�PU��t�P:s\� &Q\�0�Z�*��e��C�  W��P[�n���]nR���`$J�L�I�pt 3S4 �1�����ä�	vۀ:(
�8�`�m�iPhj�-���  ��@ ,���q�  t�r� E��P*�J�� :*��ʹ�
 �uL��(G9à��U�� 
�6��JR   �{FRT�� ѐE?Sd�U0 �b*�	*�#@Si�@i�  �J����CA���m ���a`��"B �5q���G��y||}vͨ�g � \،#��{���Ͷ��ޟ?���6�ݶ�1�lm�6��1�����!�����1����{�ff���1_��������{����85�7F�l��6�۶�����T�kXSV�ӎ��r����4���K�( ���܌"1Qte5m���01�p�kcM��K5bk�L�M�J�)҄��`ť(�����#-Rz�����nA!�����i��	��N��^�$��q~�s�6�ǻ&lg�P\��7�D�����F��hShf��c��-uvݼ,�tjd��I9��`������"A葫�7t޶M<U��X۱!�Ӵ��V�g]
[����[ͨ�D�&~��f%zL64�!S[�vf<��*�q"��s����2�zں����X����aה���;4�Ҷ��(�tk+1�X�O��ý�v� ��=��0�{�����u/�;p "��Uw0ct��6ԍ��OUe����EV�7n�ɭlj�`��8d]Ĳ)OqSƈ�=D��I�V�{�0��$#IZꕢ�oe�Z�k@RJ��4ĭ�$<����nEoiSݣ �����%��nSQHE�8lҌɉl�n���^�/r	&]�
8%, ^(��B����N�\hm��P�̩5Lf��48UcRlj�sd��W��٢Y��m�P�x��%�]4����rR;�h�e���x�@�f��w1jkFYR,-�n��#�4��VEګr�����Qk�xi�Ze��n[0�7tV�^�̚����ǙI����]80�[�s]���2�{T5�4�v�#OhjJe2�ZV���R�0$zh%Z�;4��[�e݉X(��K3�XB�m�v�ƞ��7Jb��i�ʻkQV����������u|�'5�\.Jh�Ev2�wF����ts �����.�8������A�Wu�QVFK�V��x�����"_2�M;HF�nR��&A�����Aw*j
�FC��J�ԨəYA�Le��y�dK+*U�sZR=ߥ��I�	hۉZ3&��c60��ݦ��pHM�"Tb��eX�X��h����l�����M��b��3�48�e�)ZG+6G�J9qZR�Cv
n�gQ��0k<<������q\x蕳5�Z��\%j��7�d[��
����HS;m
��r�ݱ����P8��n�S��&�4�r��!Q�	���6t�����
b8���3oK����1�S'�۳nڡ]��-i)@���Ve|Ekņ�2��.��,:�4ٺ�5M�׉�ÿk�zV�;@YGm�@�YѠ�w#�ի4�dw�m��-8s5��"�S��Rl��5�j$�w�ީ�dz,EA��O�Mc�)�{x�4�m:}dB@z�w[L�d��̷�-�d���@�:V�,f���GQ��-T�u@�U{�m�ss1��ݖH"0#��C ��Z{�Mˉ�^�B�k5g�i[�<�%i+�����%��[�"�֕U�Yo4řYc*�ڴcɬӵ	6��1c;��3
��b���1Rf��fc7�R��(�YI}��������Ɩ0YzKJ�G��w�I���͂�Y����֨����0b�骍���wK�XT���C#jA0Suqj�j�Ԣ�陴�0 ���o)=�`Bڦ�[W��n�s�Ġ`��i��3fU֧���oj )��7��г݇�6G��4, �]9\�I�F�1u�;%��I&4kJ��#U�Je�aG��Yv�B��I��m��ۈh�YW/�8�Ⳙ�SY6m��A}�G��G��D�C`.Ym�!o��EUp�
�2��L��EJ�Lm2��b�wYb�P%��L5r��-f�b&]��L��@���6��j�.�}oNV�G5%m	2Z�z)�۰�d�\f9�)�y��@�v��n��l �r�٦��/j(�e�J�U`#���ZJ�j.�pj�����vZ
h����x)Zh�(1��vP���.�N}� ��>9U�Y�d�RG6�Y������f�d��7�&����2m̺�0���ڴKYV)�m7�E3ׄ�1���ӕ4�a���Ty��гn�n1v� �Ǫ�� %�u�	4�ۀayo!��lqT��id�@��^��Һ�G1M�_0s\������E�;�ٻ�� l�b�xˉ�
�t�5�F��:��c��S�dQ��[�:͹��v��Ie�S+n���$]fU�8�$Z��d���?'WQB�Ƭ�smm��i���Y&����l�J<S�8 �ݍ���а�K�(�kQ�M���n�m*������3� ǃR�� ��p�A��-�sV��7V�+h����lQ�ܛbʂ
��ҷ��GT�a�E�������2�Z�(n,H3���NyB�Z�7Q���:��ݖ�L�ouPS��Wn�xq��P����ZP�`�!x�R�,�.h�Ub�3�Y�m��uoUGk��E�����%�v��y��d[x�k�;.�/4I����)F�v-eM�ԍԓL��q�8�p�Ű�0�Oqᛴm#�ю,�!�t�b�᫺O�Cwa���K�5+j��N�\7s~ЊiՄ�;�t
u�h��F\�w����CA��}�9���4��o��j�����gj]�� [�Zk�֕%�i,�V�u6���Y��te[h �Mݼn,�vͶ��!��Qi�m�&��GV��p�L`n)۠�z^�L�#0|���4r�����m���;��nc�V.�Rh���aGMVn=��M�Ĩ�Y���°W���F�t^ �Z�Kt�.��j��wQK�1e��R��7�"e!X5^bl�֋в (G�+�Ș0Lf� &��a�&�+��A<�Y�`4�,J`Y�l[@���Vdͱtv�j�!е2��Y�i�<$Z��E�v̧"�B9,�֕k3	�Ea��m�aa�cA��JؙF�ˌlȘvFNT�0<^nB�v�����Dď|���"��9x)|�o�O��<7�>�'�d��kmЂ���B��Jh��,:"5�-4R��]�P{�$K�ws-Zw{SX�ˬ��1�,��`yJ,��U��=8�R�ُ1��@���*F
N���ܨ���ȴ&E�e��7T[���DkDZwG9���N=6iͳ�(�Aʂ�T���7����q�yZ��T��Rt��%��&���4ÐѢ髇e^А6��op��=��~>�}�4�>��n��>������fr�������(��YF�����E���J�m�N��F^�.kn3`'F�kP���ڸf`�cs��$t.u�ƹ�е��[�T�g3q���]ȋ�׆Z�d��]Xz4$d���j�11�)�O4���V+%X�7Qw���DD�h{���
�+oР��2��l��4����OR[о�f��� �)n-���O>��7R�Z�N�j�%��SD��h�sn�۔���Ʋ~ې�� ��a,d�h��N#%XT#6�M]=Cr�k��.2�3*i�X�I��Y�wI"��bK��[X��qkt�p2��S8��q�6��V�ܢ"��Ļ��Q�U�oV
:�n�le�OZ���ۦ���Iu(���-��e�����Y��آڴ�@-e	�C�!/�vt���ByOmR7^�.�z���AF�d�Vɇs.�/�Jw[�l�H5d�M_%m=\(VT�YN��rӵ]6�C\8���@P�w�n*?�b(�i�����U�H��ɷ��n�p��t��j��.��1R�7XU���X�8R��Aj{��l~v3m#oF
̢q@��I�]K[V��̢���ö��@�X+e"�lV�wY�QN��~�g�Ҽ Q�ǩ���iХ«p���<�$ƣX�"ݨ,ѪZ�vn T/�lҎܑ�c0�0U�ۥ�K�k��"�ݕu�"Ӆf�N֣A�V�E{��d8��A�����Ű��.MP�;pL�H��
�@bL��8�A���4�b%��ͩ�Y��
^�lŎ��pS~:$��a�:�w�����媔 X1ŷ����U�1\��a�e��ҝ�)6��=��ie@����`�H�.�U�SYbV7�Ei�?e�zAa��ktP
�e�ن��y74%���Y�eˆ��{N�T;E��%F�5L�w	�3�X�zN���t���cN8��ٔ�6�,�l�T:��{W��$	ZÄ�zҶ,�,��E+����]�"�g�aշP��D��H�m��e��n �<U��Qf�����X�n� f㼡����!j��,QY*ȡMz��1S	��<��Y���@��;�K5��Ur�aۗ� ��z[D�.nAz�N���ؖ���ZԯK��u2Hգ�B&f�@�_]��Cll	L?qs��t1����wۯ٧xÖSlkP����#�]]�V2M��qLA�jV��7���Qs�/�u02虊<���Y�#�k$���wV
sS��V�a�\�S#hc(�`:a+�͢�.���'�+v�J�r�O2ƫ�i���A-���d�D�J�ݡ�����VÑfWyv�S6���#���r0��4�=�Q"�\�,UB���@l��c���,�����:����V�[�JV��ފj��[m�/V��e��4ޛ�0�>�eaِ!2����s~:f�P�2��ٗ{��z��E��.�8ŦMD�H�@�dڕ� �x��:UhThh['�ƍ2�^�����w�B�H��>�P$i�oa�d��Wr���9�ww%�S���uv������ǳ
�g�I]m��ݺ�â/��yV�X��,�9[������l"D4�-[sr�ڱY�n�B��7��p�����Z���F �Hd'�G��=�Β�g�.��S� �)�d�Nޜ�{r�efD��$�ݺyq�F��xeh&�ΩSU��z���#3%���aZ45!��:g1[��?(`��&��*k�?�y0`�/?%�M�䚲�3r:�s��(�\�C�=��:r�y����B�c�3F�Ɠؼ���=��c� ᧯bz�_���Ӕ^b���1�t�����b�dZ��mĚ:k6�pi1�T��u��������.L�5��q��^4�b��Wi;S&����-��/rI�ۙ�`0i(��M9����Ɇ�qI?7�谰��;��1#͸F�R���c��V�"w
I_K�Q�x�T��Ҋ?�l�)R��҅#�+R�k�ê+4f�JL�-�y��^�̋ �V�ɡlJ�T`	#x�V��a�F��V���;ViJ��i���J�/m���M�w5V���N�Q,�;tw3Fi�2�;���{���R���ĵE�'�&��	N�U*��a����ķ�}�-�<x��ޫB� bR�``K6�ok@ז�Ӳm��<�0-�2b��ɴp�OaU��� �vȭy5��If��J$nY�w ̗��cX��W���eZ��MY�r�ز�5�l�h�^GV�F$/5���PT�.Z�IܭϡV�I�Q
�eݩ�i�*2�Z̦�Z��.�L
jͤ�7�� Q��d�e+
f�hv3q�5��F�i�z��37Qu���E��mEX�!�R�r&ᡧ&��~!����)K���ұ��1���M-��kY�?�ŐTt`���֬3��Ld��Sz�:0wn�h���H:���5h���藃pا+,]����D0!�4v�}��!���ۄh�&ɹH��JF�v ��m��!�î{kMыW啩��%��(�=@vwg����!�}��Ix"9�K!�in�r���M��hب��շ�X	�Li�'�- c-��M���%���{�h[M�m�e��V*�m�cZu����]�Pm�E�����q�`詴�I��ѻVki�4Xw1n< �6�-KHt�$�J�[�kt�nl�m�ӗG�ٴN)7L���!�&E�rJ�T�*T��h�T%`A�nѽ&�7��K�b�+jpU�v��EV b�*�����a�P�[7f�f�8��Y�!�>���3DO�"�Xى؀����b��V�L��o2��M�ME��2S���pH&���Z%^ld��V���� QB�Y�k&�F�%^@+q���4�*��e��z�����5@t?G*�u�Pۨ���5�p�����=��`���kE^̩��,�V۫ۦ)��weɹ�orY�i�55<��*�6�6�p��x�r�n��lMB�4wu�r��<u��I�$�gl:
�s�/n�6|�W������y����1�8�6k�����|�����k1�)����b-132�-0�r��*�$@G4�A��kPDA�x%R�H�[� p�J�kU	�h���9�[d��:���@�.0�.V,t�Z����E�7JFv\LI��r��X.��
,�Vf��q��V�X� �Y0����1Mf��� ucr�c�©L~'M�AU��Se\m�����"�Rl45]���H���bh��^��Ɂ����[����鉶��FɉR��z�S�J���W�8� �::��sVV<W��'�%6<�TRefՍ�eL@�n�"��X�0�&�V&�YP���N����@tȔ����a�LrHS:6ܽ5�u�*���2☣EZTw���y���&7�7��yZݹdNɴy�4�f��57����{���j�w�Eh���) �XE�*_Jg��θj�u�U��w����ۂ�3��BD+�;���a���.�AY��w�N��ە&�Ӡu&��3�?]��M��y� /K��n�d)�a��Ϛ��/-\Gc�㍄�\�%�*��ҍd6�H	yt�E�6,�1g�x��5��ZN� v�B�\�c��/����h
�[�c�O��3}<.(5˛#m��]���jSv��O��D_m�@.q��_
��V{q�2g��ڬ�t�N�]�\�ͅu���ܴ)]�|�����+-�%,�]��m\-wB^�<.�x���&#��r}�]�_68P�qSY;�e-��DU��B��?1��`�;�g�>�F��y�ͿX;��q�x`/q,ޏ�����n'ڲ��1O��Oi:�-�eP�}�;�h�fpN�x�o���s��a���v��
�s�+g����tE�Lμd�"!0ç��le��5I��|N�b�U�v�ګ�r	�<�ՎV�_g}Ѯ�4aC�C���Y珃NUW#{}��oC���KY��N��螜k�I�N�����̬f�VjYЎ�ڝ�#I,�R��)��F�rrn�T 6փ��tq��	�f��M�ނ�[��Z��⡝J�EN>~�q�{F�>y�������.���R�?��wgK�z�9���NN{r�8���.����"&����z)�Ej�|sF��%1}|s�|����Ø��Q��<�a\&h�3���=>�Ң`�Y�NAX�4�8����]�*x'�fw�Pנ7���}�5�:;m�u���WX��N�+z�9�6�,[��<=0�a.��b�q��&h<J�7�ݧ��0e�n��-��{h+��|oa��|3��o�^>{I�]M�%V��'�{]��y�RS&���W����I�,�h�cؽ�iW\�t�\yu���u�Ta�};�>�6�����|�����ډ7���2k�#����j�n�W~�v$y�^yd/�j�S*�;��@Wê�q�@Ax*^̶���Z�#(�=`*G�	,j�*��&
�]Yߺ�py/�F�(t�QMŒ1"wuٗJ�M�#�u8��P_'	���A\�r�6�=������B:Q+��� a�ȷ�@�>u]��T>�=������É���sc�Y����ɾ�8�X�2Ԏ��Mٮ�B��F�Vmk�+�[�{[�i	�V8�bp^��@�Y��F����v4&b�fe��%���.��qU���ĕ>9a���(-�Y��$�1"�]q
�,�ܻ��[��~ކX�R������̒��46.�W/Jw+M�.�Y}F9�)�P��t$R�g���%!��;�WZ���ɝn���d�ۭm�
�!.-6w�G�귞ooR�;3�����af���ѧ�hȖt5�@�!��
ܸ�A�R���ą�CjR��-fZ��]l�1�[>�����Ob/�)�v�@{�4���3m;#P��-8�����R�`k��W3�gk<�!u��93U*w�cVs��`Ze�=4�^]�����	��#��,ew#�"ۊ����#Պ�o��=R�*��,tJ;]�~ ֠R�o�a:��2������X�橹�)foV�1`��Q�,đ���-L�}W�B�����']Qw���u%i�n�'��;87]�s�q�:,���*��پ�� 0��mí�т�(��=sJ�ܻ��0��Z�8ɼJ�W����j[[Z��٦�N=�h���v�F�o+*P��cr�o�L ��`�o `TU2��,:_<����;�����xFnԹ�w�0�f�[�Nk|#��}��v37	�/nh�\m9sZ��(����p��8�����>�<�k��M@�6���b[y8�`j5 U���[��=bR�ـ��{Q�q������Z����h�+���q��՞ w1��#�׻�����&c���)�Mѓ;87[�`%s_˓򉒾�C>�D7���p��o��zI�L'ؘ��gS6v	�Ly��6��Y��y��&���{��Y�+��U7��/�:V�wa�'�5?5ag;Z�hM��rTÛ5!)���Q�ܮ?1�^���6o"'��,:7j�N�.y*�%e�no�ڻ�^Z�S"�ʫ0[5��d�8_u�2y
��ʿ�G���f�jc�]�gJ9@Hs�ZS����l��En��� �A֬η�C��֛d>B���;=G�e���{=�ݷ�a;H���op�Ņ:��ru<�z͢覶�I��~�zeˬ
����7�gZT̀����q����Ү�e7�@��{6���;��|����a�j\�(���V��W��A��1����pa�]:�7 b,�EL��	���2}�!|��9i��Y�D�r�Y���E3+��|$>jq�`T%�'�g]������b=M;F<pT#���p�`ʘ���~|�tkB�_f\Wг�Q,㮵��Jy�c�A,����d�*�&�͟_����X���:�Ӽ;�k��Hy�g���=��ڛ�>���4��ZSN��[�W��M�3�[c�x́۔7*W�ݕ���Q�s��ڡT(bK�ŉ�����Û�/w"k��x}2���)H�����UQ>�r�^�RY�\�@c���.��2�bz�$���*D�,���}V�M׼��Vޯ��*D��LE��Vyo�J3t]�˝� ��ɥ{.5��Llr�_���:oj5�R7�v�f@��e,�g�w���3�"7���q��)Mt8��gO. � �'�G��I��D�3Un��'Xe7i�2�����љ}ðoK�_,]���wG8SˣB�OP��\L�W׃b�1o��)v绝����9n�V��5��SÅ���v�=u����^@-?q�rQ���=�jڌ\p�_
q-��ՌIJ���w����+{{�N���J�8mb���2Z�����b�#7�S����=���N�|"�DMS�s��xN2�l?����8��R/M:��;l�X��D�ZkB�v�gKfNI�5��"�"��u��}�5ok�������D�mD"��v ���z:'���s�d0��6�;J`8{y�gq*9dK��a������ck����G.���&g%kzg����Z��w�u�wI��$X�9��f���y}����pe Z&s3�u��nn���ٵn�RmTY��ڐ`N�}��r����J7�Ï���	t=�r��˭Zu���Q���qa� XΣ���Z��C�k���v-�ud��h\�
�r�A���{|V+ݬ�%�W����eV��iz�z\������}�� [��t��=�[�1Ӟȯ3g��T6.A����7K3�{��0/���%�]�N諘n�Җ- F�J��[���w|)�ɳ�w����T`˃,F��9����' ;řa�zE�Nw�"�Ҳ��X�-��+;]Z�b��ۇVU�;�tW�',A��s�};=I�qS;���ܮu�2ڳG�o�;�������t;��C��w��җ�R�S9���8��J� ڧ�5=gm����6PGdTS=j��sY����Z7��;%ȩ+f�6���^�)D����c�Bj]s�x�-���z�18
�K�X'=�Т \Wk.[7�w}��6'�����Y; W0�v��Պ�.�H��v�9S|�^[, �z��}�A��Q��2՘w\�����͹u�%Ew��#@��%gq�$jS��J��5h�y�'�,��ss�J��h3��j��N��hWn�/��3�QQZ��+�鬙�����,(�����
�3��aՕ��~|�/7Aw3�J��~�����6�'[k��ީPfq��"m�`�k(k�Kp�.����޲W��]��3�|/!��C�z��;�w�w6����Y#+�����t��*�m�P�V�v��k���]0R�h5aS��p��l�7pGG �Mܮ��y�7,l��d�۾��FD�^�\�ޓpd��8H����q�
������E��.;|�`���9SfƧ�d7'�owz��	��[+��5!.��J��`�1
��q츾O�ڒ��=�4�p��q��"�Sz�J���|ѭ�Ul79�&E`#:!�e������V�IΉ�h+�1]m�߬�h���=	�^F��}���ihV�oo�W�c��
W@*X4��;D�t�|9X-:���g:�νr�ʝkZ��<8P���BZ�57Ѽ�T��~;�x֝� ��b�"��6�T]�	W�dx������嘟dm�㵄N����B�4��N�^�Wo�p����plx ���Kf�wK<����wr��]��nX�[�Uzs�r�l������ίV����>�Å�}�
7�/����P7�@Q��Z;�ou�홛���oB]u.@`v>������70g����b�l\�Ǻ\�6PV@�8��W���r"�pz�qL��r��r��|E%6�8�;�u^K
�z��)wZ[�_�:w���H��a h����8��G���{�G�cwHRs7�jpz�>������3�-���uƨ���v��!����έu��T{�ȼ��d�dp�]��&#�M��Gu�ݣC�-!R���udxp������p��1�R��~NͽS�m���_�z m=�Yc��f���JF���j��ve�I�h�f<��O�-��i�ں=����� S���n�т�ѳ-��m�
1mu�F�B&��h�YD􉫇��D��)�ދRZ���X�@x2�Ҽp��W�k���>W(�[][��"��]����,�x�=8c&�|��N,~y�t�`��:�R�r� �k������bw���6ܝl��=���C�h�?x��փ_���ji��w׵*��\6 �Zµ�K�|nn��!V5�x�C�tR9\�>�֝��v�CiJ���j��z��f'�)��'G�p�YɃum^���[�׬��h�7� Yd̹��r���e_h�:��%�p������:�����qӕlvE-z�S�,�F*��z4o��J[�x�)��f���� �sb�c�������qy��@�/{^��bv-͗�n�ո�sЬ�=dɮ�+��N�\:�v�N_�m-u{ӎ�����<FS+G%�&^��L����wNU�~9ۋ���K��W+Y]���Mqя1`��*���� �x����,ځ�������h@��v��;
j[�4?SX{�h�o�pɷ��4��ø���/GVWm�[Ԟ_+3��=�;v�e�<�������#M�=�G�#��y��i��׼h�����vMX���%���D��<�8���YS��+���:���2���ܤ�'wx�C�ˡQ"�]z��w9�����o%K��Fvc148-0̼���d����Os#N�7�]I���H9�R7�;���ǦLN�(w.�]vk�m����R �y<���V��d�y��\N�AP����$w�w�i��@[N]���c�)P{�Ȧ������W�µ���	n�hF@��{���+v�v��a�b�e�Χ<� )�W/o�\9�s�jK��v[MYvk��>Ӟ�1w���k��)�%n��8� �!^�ӻU�^���U�=���1�k6�;;�K��6�b��Z���A�4y����<�K��4%�]JDEI���8�x�\�.ag/�d���/���h���C��]��,R���P�V`y]���Rb�wx�a��8P��oa���{fk}S��)��q1.�2M��P�$����npN���Z�ۧ�Җ��/IʁM����N�C����ƥ�:�5E|BC9n���>{xܲ>�9��n��AK jM��/f�+�惒pW�R���w��$эd�vC�? �s�i�{4,ޙ�Q�s�l���_v���.غ��&_Ib��ۈ�^��,dL\��o�q��{;}����}'Z�'����}�kZP=������R���ȱ��	�����T�¹ֽ�8�o]6�����#6�;����٠�b�&H�A)��mv��@h�d�)v������c�8�T���ubs�݈
����Z��MD�wta�!B�Y���Y�"/
㋏v�z!�ő9�d�LwN=���m��a��5R�u��I\�ƶm]��	GmS5�ķE�2�uY�g��� T��,�d�,�tL&�;�-�}(��d���	0�@�mO���:.X�2-���� �Oc��́R0����w��"|��X�O.�-u )*}�7����~����,�'h�Y2���-k4mۮ&(sjGq/q�˗�@4u���`�#x�Qt�%m����� ����X��؋�e�����s�7�� *��z���F"�r�Q�4�,�^���i=3l�t�މ>��1�|ť2=�Ż;<��������zn�{�8ۑ�T���r�`G�W=�X�� �q��ݩ�P���P]�;'l��͠��<�����R���Dخ�a���(v��2�U�Y�Ko<��ڰ���$�e_�`�-߫�n�H||Һݢpjt������!�,Z*��$�]��]ZW��5�/�2���;�|`�3t.��WW����s�6�����^����>iCb��O-*��\��8���s�}p�P�}��S� w�9f�(M�l����z���٘�M��D\V�j�X.:��O�]%��p]�!lo������Rh"�����%:"��a�3;{�Z��E�c� �±��wd�����VR��`��	����K�[�ݓ�m�M������Cn�a��F�~+���Y���S���5�J�ٽш߶���W"YIQ��ݔ��ڪ�e�z�xk9���.��Tzo	w�%�<6�c� ,R�jY�e�sNz���r�Վ��#Q��K=U����/�=�e������[e�'@{���ϟ�m�6���m����^�|8����3�������3d'��3�:���Fv�Pc�mK:�r@3sy	�rg��>2�����:uܡl]ۣ�����2+N ۖ���W�����Bē����7z�ё�$�"�K����?n��NAT��5��z��	@�):0�
8�>�P_�0hذ��Uw;D36�����N�oq��&a0�,� |�#�2շZƦ��D2aJ�yc6&��y�}�e�ڠ�MS���
��������d�9�z�=��Y<�z0ocQ�|h�Ky�v�f���+=����Z�Cp�&���m�^��X����=��q+�fq@��W�`�*r9�t���qҧi.��r%Ō!?���4�x��U�W\R7�%1�v��sdD%���+�b���;����6 �*;,h�V԰�,��L���9���%u�X�Z���jȆN�I^�pT=�:�J��/�́ko@AB�,�Z��*[�1��b}x��+W
7ՏiTs'bmo�,3ž�i=�㺉�n@���a��l����ïuYT��v�������=o{�����A���}�i�Y�ϐ(k�]���fwi�(֍�-f��x�F k��p+Qm�L�L݇kg*J,��H2sE�s�xҰ8u::�:ߜ�7��Rj^�g0��΃&����HW�D��1L�L�ܭΩA�n��iB��<g�υ�[�����q��:a���(�K4i�*|�#E���Ȳ9�Њ��U�����c����CZ�M�/�j�3&�S7eY�)����ZA^���!r�s����S���no)a���hL�1���<M��(���+]�B�70��t�;-p}���P� %4-���h��
%��ҟ�]ټ2惶���e�EZ��\�	�xw}A�������Oݶ�=.�t��E+N����QD�N��f]ó�kkz-� 7ҷQVK����d&���5��Y���~��nׯ2x�v-�_�-���kޖ��EAL���t�H��m��.X�I,=���S�{ZA�؆�G5�#��0B s�}HpH�2���g]'�۵(�k2��	׋���N:�u�[s�s�A��$���Y��xڸ�x�e��;�b�[��GTd���]��]�����n5��5��?�%��qM=ih��ўQ����+�7�
,��E��xcz�#<�W W�f�g���n�N9y�#�A�(�-'C>#1��p%�����	�ஞ�k��AB��G�i�k �EӂS�1�Q|EoV�4(��ґM�.+�ĥ.1�"ek����0pWx�@�W'V���<�pg`���4ƕy�X��)J��7��k�E����N���Ѻs���=� ��E���_��c�"1�f�\�>T''�@U}��Y�6�����yn{��G���{�R��o(fФ�kng�p��ݥ�e:)�X��93��-&���7:^�+�������<��ס�f�)�&ɾ�L�a�F���K�Zy���!��L�Q�\oB�Vww�^+������5Iy�ST��[8z��U���Ɯ�Y�n��4�9`p�V���^5`D�H)9�`֜�KO㆚$�4�	6�V���8f	��:"IZ�T�����$ ��3:�&��W�\(�|��+:q=vY��<�{�[L���eI|��;;GWA%�sԳ�3ޣ��V�,+��,1zkQA�l�E�՗\[�Âi�Ů��Ph&�C��u�1���ީ�-��׸�mPm#Ws�Ȧ��b��9rii��Wj���W`-���tx8��OU�0ч�G]CO�1i���:�g��k[���A��E�e��u\����t�z����]�J�d���N��ۭT�9Q��u=X�qA�yԱ���/a�m,Wk@FVm���>��"���U�#��F��ٸ��:�O�*S[S.Y����V�SV�m�X4|����B������k� oocb�^v��40(�n>��R��"�&��(�LV���7��ǯ.��jq��u�$X��`�]v����ׯ5aN���gXæ��j�h��2��c�:((�{u�.�nK�W��O{����fE�s��Pd7�c���;��{	�z,Y��ٰ���l�����d�}�IS�ݻ�85b�X6��:�qZA!\���;��X�5a�ή��{�0�t\�sB����Dk��(�r�^���U�R;���A0�����!��M�G�oM��v�n��v���GF��9Gw���b����f�c�xZy�]Z�����N Μ�v;*�+$]��,c/P;�ԣ���k��%E�NoC�%h���C@������u�ռ���8qWEl	B�%��q�w\��(���h�w\)9��ni�	��uW�d�hWT���0��Wk�l��Q�yTʙ9��Eڭ�`ĉXN�k�*�Q����WV�
]|ȻH�����#%�.+s����}�[�������^�8'Q�aMƏM	�gH��T.�����.�͙�FI4+�1�8˰���"��3�tg�4��5������h##��\;C�m�+n�����N���Z$�N�؀yä��~|�*8h�����
��:�R��]�%,t��LF�����U�5u��f�9��!����#-�^��F[���D�,&-�X��k�5n�\x��4E�� ��/ۑ��%lu�'aE��tN���ڒ̡%�Cd3����92r����-���.<ʰy����̤�:���ɿB���w	����g��-�t)�N�-�Z�^��4$�.��w-w
\�T�����n��i}s�3�GXB��_yQK����Id~&��M�aov�<���}�=x(ri�>�,a�������2�"�\<���[a��V�$���z7i� �Pc�F�#dT�j3���D�wa��H�`"W�j33SIMy���y2ĻGk�v���Eږn�r{�ۧ�7�{�U�c6A[�tg4l�;�IH����`u�wp3��g)U����KY2�����j��g�s�v:���;J�-i����[8D�7�W�����ck�c桸�P:�/�rv��M��%��� ��A�e��(�r��ô���M"����^�ΘM�O#�ؓ9�R}0��������"m���ٳ��:2ѹ(�I�3WIR-�˼�n�.� IW3kMr�;
Nڴ�FE�y�`���wI�W�����C�7n���
��A�n�(LͲ��
�0����H� ћ���9҅�/��	R��e���I��}|z��Z��b"���毓�Je���������F��p�\�ҺO�T�ǙV�x]������M��޿t*�K�3�4��Ϭ�h����d�*p�va>��m��¼�� y똬/�T���u,�}g��2bb��e³�mR��Oa��
~�jܶ��3�Ԟz)7�U�z�y����y�#�>�`5q������3��4I�\���ޘ��5>��/�_��v1�z��7��,�[!+�'���x�clhnm#��^𰂢՞���򾬋	X% �u�{os�8�.����z��_�ߊ�Zyu��
wq���[�Ẃ�Po��8�����W"l���3N���
h�(j�oy�]*k)��R�:N��+��ظg5�DQ[7]Le��
R婊1�X�Fվ���=O�rWe�jy�ժ�s�]7S���3��(IF����J�D� �KN�t;��xi��#9��+�����c<�W`Ű������Fq%����� ���@^��E����#;c��B�ڶl!N&�=���OE*l�ѵ�[����-㞬�C�cW�Z��U*�a��;�:aR�}0{��硜�Yq9�Ș�]P/A��-��0�}�ǵ��ed]C@�b�������|�=����>�g�ȬA	�@�ʬ��q5huX�"w9!�GD�U#r�*�r��]t�����|�Z�zZۈ�	���̊�74�̬�si��ɇb�#�X�E�GN�k-h����y�e���Pe�ϼw�ݾS`��{��KU�0l1#�f�z'�6=C�,X��A��_@�+Y���6�Z��S�y��F�ۅ�k��X�f�m�}�x�96J���0��ם�2��g�]w�
�6D��f�vB���K���S@]��":�r��\�;�Wv��*Ǖ]��5R�i�=^3���+���6�pi9-��5w�Ґ#�f~�i��m��,�E����ޘm�'��1����C/��qp��]�/^�z�;Q�Q����eb�\[��gg<��`�]�.�=ԥe��T��;J������Ph����so��>x��9�+�`�ƃ�(�V.��g_h�E`����q��;�뮮�m�U_[��(6����%+X	�<�k�@��bE��Vq2h#��ӈ�(����Zy`�;a��Ĵ��(u¦#-��^'u��ϵ6�Y;<<'p)O2�^�${�]��ij�Y���M*�#���T�!:�����Jj�gK�S}|���Jo9��#���%e�n�srI�ol�=�=�o�G���RqḞ�s�$җG�a�4�D��c�Ie�<�c������i�Gΐh�������U��ҶQPq,����:0�z��k���;M�Z�N���ܸ�gy���*��u�w��{ �%�7d��dC�Q�9#kQՓ�|:�Y�c��{���ŤVȔ�.R��P�
���팫��-���p�n0�g9Rw6��Vb�%W��d�uoU���]�����{�����@�ży��"�+�I�NB��U`\VykŐ��Y���ڀrA�cV�f��(
Mސĵڮ���W^B�k���5~�N&:���i��:IV�u�Vq壻�=t[�Sp˱�%�I~��6LT�Q)��z�ǬW?��
F��y��}�{b�L�����s�V�%z�.�+����=�3),�c��͑S2ԡez�7�'�9���#�..LR��3�sY/��T�ۤd�f)}'�RL��o\`��zK����]�8R��C�x�<��a^�:T�+�)@s:���������OZ�p�?!N�H�f��N2xzf��+z־y2^��Υ�Qm�J3S'���pV�fj�]��m�?O9�b�+[!ܽz䊷�ܜ��(�ܥ͠f��xS��F��u���-�@��H�{rs�޴����p	Hw-��a*=���a㪱A2���;S4�^�5�0�^��Æ�j�Nd��6zP�8,v5�AyC5j*V�w�e��.wZ5:U�'���	���n�(���y�W7�u�S6V�Բ��z�(=}�����g=pռ��pCra�˞�y�͏dÓ%��_ċB��1��/_u5�;@G�!Y|�~��|����1�Zha*��#WUA1�,��n��+3;j�iJ���Ζ21t,'x�o |d�Է�.TNv�=��ǆ��)��OH��ݢ&<8��O��r���hzn ,3k����EG��v�?u;�z��O{�~ȅ4�U�8�gE��"�Lu
!����:s��r������c�}ä� �dy���Bb�n7s��y]�ѫ�͹6;�*�(�Բ��@��n���{�	�j��1D1җUU��(ne��W�cC!QM-KZ�T��e��?#�b�:B.���gj;�)uf�k��W���ti�՞��;`��.�a��ט��"q�c���\�t����6{p+�
�*Y{J����#f��&�uEʅ�Ѵ�Zj�z%]!���P�0��]ckr5�Ұ'L�d��]�0v�W1�b�%����-qX��e]aA��zn��1&Ʋ��tl��|�vm�ۖ�����se�v,�s�P��1-��E�Z\p�;�]C(����'G��m�v*��ʾ�&�3
�u�c�U���=6q�w< �nݹ� Ҟ�$�eoz3E�ClΜ�'M�D�&xJt�n'-�i�����"��E�8���[�)��+e�_����H��-Y��	��������:7M�o�/�������o��K�Z�]�|5ܫ��O�\��ù	eO�J�X�ܲ���ub�Gc�¸"7��t����o�Gn쫕�}u�9��\6�݇�Ĭ����w��orå����go�a�;W�{�W�֬���R��C���G�Ӣ���[��o��ܬn��`�z�C|~����{/+h����U��MHN�m����q�H|K& ��9.w�������sod{�����C��ȎR��f�%f���F־SmS皗^���Ka��b����;#>f��z���z^��D�<E�2��0��Hb���u����\:��8�v�������u}9�ʱ��5	�;�ɳ��W.��2M�����og��Y�I�9<G�֦QЎ.��w��U���.y)�O|L�K;nv�47�'o-^��; \�չo+�]�"M4�"k�7���ړ�Y�cw[�$t߷�8]I,>I.���n��˙RZ-Z@"���#�W���!� ms����M0�}o���O��6��;�P8�of
�[�9��;�3�x��1���N�'�����\9�K�:�U׹�$!CԒ/G��P]1�e��K%c�v��.I��2��j�P�	�����/�ܢ�\�/#BЮ����|�sӾ8��,Y�t��S[V��r�q�d�#&�2��Ǿ��ۑ��8�W\[�:�a��A���N����h!�ˇ&��[5C��J0�gc'�W��es�7h�Y0���]{B�����h2
?n�/�s�����|�����z�>w�K�"�Vp�Q;4��A�.�����5��l�\� 5¯�j��߲��aѬ�*J6O�j��V��@��������o{��Y��l�u9��M�{x��P��T�8C�91�\l����y����6�? >��a1qE^��^�*��,6C6��m_w�q/� ,��]b7=݃u���r�:Ĭ
�oZ뷘�B���>���Hrn_�k\�?=�<i�օ�=Ko��f���΢I4*�by�wp�r:UE���d5��+��,6Zt���h�t�4��Ye���x�oTr��eLl�F����#�������=���A����	�:FOX�=��.�F�YHr�p���qm�\B?!��z�e�>\��"*�y^�O�U�|se`՘��s�>a{�Q۞�b�V�`��U���5b3���J78�����í����qB�O�%��ݸ���:���So1I��sG��H�2��w��w.8�g7�^�"�C�7:�8�a�f�re�©��[��A��(X�� T��*Y/v���OeҏM<3���rZ9al���cZ��t8O�F���,q�!�p�y��Ȓ�+�ju���ۃY�:V��)�n�'��']+J�>��p{ӗh�5&�6�P���q�H�ܛ-b=v?^V��2�T\g�S�,�Sw��s}e���}˶ٚ����^��.�����F���{�m��Z7z���TrS��!0<�\D=׈+�y�ޣ%�����P?�P$Q �PH�q8��+�
V3JN'QL�D4��� �\�(�J˕Fr%:�QaA��59h�2�l�$���.]"�
��l��2R�t�e+�H����ȓ�HZj���XDDU�ISR�.��E�*%��*�V�C��H��"�(("�R�HF��JЌ�HD�
.U&I9WHBJ�!�c�CYZʭ%KZ\��qJ��1IKR(!:�#kY5
��J̵��I(��2U�{�q�+t=�QLH�䜱2�������SKd�U��+2�4�"M5�$eaZ�uJ(�K�R\��snW$� N�d��l��Y�J)Y�*l��wk3
�a�l���Q�B�%E
3Ԝʊ��D-�F���VAT��Ԣ�U%"�����'�;��Q����B�'�\�ݼh���S�M��YV:(zMH�B%z�ݼ.�h*�cv��y��i����|`7'���n���y�����`���Z��u������������&�"�m%��܋HCY!�����z���R�LeY���w���.��ҧ�y���J͞���b}O6�J{n�
t��d�)��[#�J�U0��@�)�v.SV=�{=E�w�՘W5�:q�����Y]L�:u[~~oΐ��:��m����v=��G	3O[��iY�<�B�G�v���K6�F�{S���b��KPO{�)%�B̚nX��}�s�ۛw��Ơ!&�3�1�ܻ�R�v�Zi���Z�Tyn��o:��䵏vrsu�!\�33~��.�Q��\��Z�e^�yg��H���$d
���8KX�4�&<�_�!�����!8����54�]B��^˼:��4'�gN\�	��b��N/c��L2|3����T 3,e��Ur��4Qƛ3�Q�@��ovay`��'Z�Mt�J7D;Z���L���un)ƌ�&C�@{��^�Pj�����M�) �g���:�����CYt��a�p��7Kb�ߝ^��B*�~�5�������hL����"pG�������F�[�
��v��U��J+�Ca�π'rY�uw�q��AD�uܦglx���Q�cV�}���1+/��d��N��}��RB�y)f�v��Z��� ���*Y;)�2T�@f��Ӥ��}m�rǵf�{.�5��0�HSH�Z��"4z��n����(�L�?�y��Z wc�W��g�1P��<�������Iĳ��.<^�ž�$�8����{���T�|8�����.n� `����8�d�È���*��xeK
�گ	���V�L^�5�#kQpf��6��Ц׽'�<����+��%�]k��%xm�7��3����������Dz�Wq"wy����v��Prc��-Cƙ4�?Õ��c�_�����5�o�R�TD���HL��!����`�ͪ�l�����S¸ZȜӎ~��`t�^�t[��~�J��`+�Y^�~�� ��M�k=!|���g.~~�*�5̑]�+0���j�W���ߞ�K��mW�g��}�u�mK9o5��8ܭ|d�����)RT�X��|]P;�������,� �p�J�������J>@�����wjmF9��,�6����v�+��n��ՕZf�C]�����x��4a,�q�¥��4�r�up21��8Mvy��S�ʄ����΃�뷴C{��륗w���f���ϡ0ASh�*>���E����^��la��t+�ee���z�a�|�wG݌.ם��)�m៙���A�-[��#�)b.��Cӻ}V �H����W	U�]>e�^�fn9�����E���/���2���ɪ�(dG7����˾���~Si�'N4Ƒ�f�;e���Y(N����L�r�b�?P����No�G<~Rs؅A�J?	L��L(V��U;�R���e1F�
l�W�[�yy�k��Ȼ[9�ٹ��}\V �����-%�|�o�+o>^����n՗(s��3R��jKH�mD\��mR�%�<�d��[f~ih����O],<=����|�j�"_7]]h1V��M{傐]��ϔ�|���]�AЋ��pnqxVU��0?��lv����2��±��)���U4�\ ^�tb���*����<�VY�����i�3�8y��2�kR�P0��]Ȕ%6�,��򗛢D��[���(e��Z��#-a�<y�Av��j�<{n�Ҩ!~
�S-M,�ۻ�5*�q���^�2������
�u:�^�Y��Y�ܼ{
]#����.?S��~^˺�6�g��x1p1޾{����0��=+��3�����D�k�r�	S�`\�tz(:g;��*��TT�ڲ�>���ꐎǤ�j�C�-K�co2�f��Ӈ.�5�������O�<:+�������h<5�$����W����v�T��@�}�}H+��ٗ}���d�4T�q]��
��]PL�*�s*hX�C"+ֶ��zdUxu[�B9�>)�}>;�b�h�yn���>y�
�P]Y�Ump��2͚|�T���[�L��v.r!<��So|��u�;E
u�W�݉�Z�(w���Rq�����Z/%���I��3Eܲ������b�S��{�(j�Ҕ[�k�u\u�U���ٮ�@B��zm�#�>����z���Q�3�2�YԄ��{�\�^��A�F�R���3��T�ft�D�n{�7���^m�����W��:P
����j��|����^CcEJ�vߜ^��N���Y�h
�W/Ӌ�&����c�k�Hxl�~t���;��}�׷��z,��	t��N��gԲ<u����\I����Ƣ����i��h�~�sej�ȅ�*�N��Y�[r�/�w6(���l�n���"�.]�Lk)��-��|��Ĵ�М�4�.T[����6%���T^�"�u��c��u�k��H6C�ڗ�C�'�Y�;<�� �a�.����z���"bsط�iŏʇS�����5*v)�;z��W0�$�	d˝[���֦���lIU��x��� :*���<=Gr�s�!ϑt��tq}�)s&m�����
�`��ז�/�������Rz+U�@���s���!��ڔ�ӣ���S˛�����T�䡱�Z��J��Y�BL���d}L��0��ܸLs�����b��x_�i^�R�{za�(�f� ��6x*TжdKǇY�T��u��bM��FG��#����t�(��k���^Y�f����X�V5�۱r�b��zz�W{q
`z��Ώ7���S'�ɽ�kA�X��ܨ�*�����E]3��{��T�p���oq<`#�k@÷��yh/��^%�_��D�?V��D���LR����o�=�V���*�U-��k��C�@����{X�,�P�U0���ݛ{��]%x��^���y�^���q�/ս|�x<�/��V �^�i�xP�ry�%�-J���"__{r1��L@#T��-m1zco���Ah�4�)�ǧUqO�G�#0Қ�m�j�8Dk%30R��V�"i����΀�y��=�(O��-hW��-�7"�*o5#�ך�rY�79�:Ȗ���L����[���$��rC��#�hnj����`��w����}Z�ɂ�X��Ze�5��^ι�m�t#줝bN�m�v��x�XQU��J��{���>ORi	l�6l8�oK{b���j�f�:�+���y9��|�e��G��Z��o���%6<@�]� R���,��ܼw���KL�⻙�"��L͸�~��+��e��7�'^O��)��+�pQg����3�/�_(�*�;���n��Sq(�r���d�^3U�����ʠ� ���/�MiN������p���K��<�P�8��*�ja�[�	B�k�'{�xC���`��d�x�>X����I�v����̮�~����u����d��Ch^�YP��k`�A��υ�ط7�s�k@��'�?�� =��S�~�vg�}ଙ41���&�㊷�{�Ƶ:i=�݆}�F�Uzၠv�5�r���*��\/c�+W=A�m��ּy%P��0�ҎͶ�fd������J���ʀ�Tm,����T´K��,fS�������z�z������;xS��<\ߒj�v:�Yވ���.�"�u5��i�ǃ��|К������^A@���x��
�/s��ŭ�����>]H��.��Doh&�:Ŝw^Q���,-,���$3h�P�Z�{w7J��9���N���5+
�f��=��\���
�)+��>�f��ۥu].?��%^�nR�x�˧���jeno�1��%y�\����"�����\WYz��7��9���,��f`4��<���	��2����G�i8����=�L�'��e���u��Y�����e[pp��y*V�
��Y^�~�� v�Ʈ	�z�[��'���z�1�k̑[u�y���`ݮ�p���c7�g������)�}���њ��;D��c�,�U�]�3���q���/ΩEV=�nR� �|7u�^�t}�C�Wi|���ru9J�ݔ�@i�L�x��+̲��=cB��*4�MM���EU<��?���Ga�e�%V�}gj�{f���N��t��M;k,/�}x��J���<�=�.]�`��d�Y&6��I�}y��/��e�<�(k�v���Yg��u�/
:g�2B�n �Dk����̣I9&�˹}^B%�Ĥ����S
�����JW*�ym��r���e�L�wu�Y�E�g�S.�f�$��� �J�8-�VK�z�Cx��L*��¥�7�P� wR��2ɲ)�Ԅ�7���E�B�cͦTKyl��@��s�4�W��֎�\�z5�Ջ��~R��j0��ި�9c�M�e8V]Q	�p��Nnܭ�h�p��:S\Y�
z)"-���� �#5���ԉ�������b��c*���7^7�<	�����A[���q���%/7��>>�e���0}xg^��'��ڀ���-�5�-mh��^*ϔ�@��,�:��Gi��c�&�A�mV��5�FB��]�������=���#ܶ�����뼛�"a�Vn�z����x΋���N�00��]Ȕy%X�P��B/7D1����+�1!�������H����xS�}�ԴG>��i�{a�
�S-M)M�-��N�Y��SPu7=�o}�.#��͑^��`gq�G��wF�Z��?��h:�<<R{���觖J_vՅrO��/r�-��@�q�� ����3�<+�վ��LQ�ߍ���x{ 7���U���{���-�~�i/q���9���]�tn�����n��pZ�nd2ORzn��j[.�^���y�n����q������+��ݏ,W�i`�lVȫ�T�|��|� �V��=s���j�7}u3ɋ��f	^��p��b������{�����Sܖ/���!�|�]��g���U�ڼ%_����x��~��b}-��ؔ�Pd��n�]��;OP��������qaO7����3=ok^�{��y���Ph�Ş:��F���ܽб�������=�i��ͥ+���AX�gf0rW�����}Ϯ��������6��ɆP���-�+���������[�f�b�!G�b���u���^N���#��?ː��V�.m>5w���rgN��n�1]��y��b׾��%8k՝��׭Pϗ���>�3N>@W?֐��U|�����{��[6�#0{��OʹG{����<v�^3ָ�ҹ?Ճ8ԺeM)�Q.֑��*����,��o�ƺ����R��1FS��*l@��1*`�����60r�dܢ�"��]�L�25�lK�b�/�-��vOױ�]�<}cU�)��COJ(h����U=<Y@�n�Yל5`��ج��NLl���pZP��4���UTD�Q�W��m��X_K7ގO|��N���88�Z�	�F;1��6����C k�%%M�׷�/9��ږ�xT��H�н��+�������'�aP��.C���=�p�_a�Xf�ɔ�7��]��	���"�y�~ty�#?-L��u��Hg労[���~�)زJ��N��۝\�
D;����\1]�(z��e��`��99���
!�#I�wcn�jǵ�LdB�MaS8)͝>f{�VI�XQ:y�/l`����^��h~�o�)���q?i��8��a睋��<���v��G��z���:�q`F#r�ޡi���'l'w8F+�oD⬬��NJ�'��P��_Z�y��v�Z=��b���h��`yC�@��$%�Y�yT'��F�t�����V�v�m������n8=���zw�����E������=�:C�Ո=�$|�ۆK5��z��{�J
=���q}���kX`�ܝ�/Lb-�;�q���4��μ�m-	�~ݞ�7:�9�m	�aq��Y\|ڳ�)��V��C�jB��ad@M��r�ǩ�5�{L��֛0����Xu�R���l��wK��|����Si=�_7�������"]X�J}V����npB���Ĥ�~�����v���,�y�-�G�HWT��V>&��{A��f�)��jY>_��sD�����zsv:�U�zyw���E���ǈ1^G�`������!��h2|�i��QZ��pE2KE��1}�����s]���v��*�*�T���S���n���|v����,���a�T��b�6+1alhV��B�8lwxaPH���!��%����9Bޫ۲0'f��b���-�r`9{�HU�R���{Lک�m�`ty)���n�u���n$s�k���us�ih�4��O`d{�BG��%�G%�ܜ�Zy ���X�ݷ\��t�#Z��u�ԵޛF�;+� �0�3oBf��!ڱ��p����l�?Z�����o�Xԇ8�jd�ږ���X�{=M�1�����XW�I�Az%��<|��;0]:��i�:�ky�.>�Ҋ�'Q��~+�{��W~;�K���>-A���:�qU�󫷝��a|(tВ�x�h�����Ǜ�-���ݞ��s�l:aP�YO=\�+V_#�N���0j�WW��`�'pu���E{۾{+oc�!�<g�^d���j�<�\\���K���j7u�:���Lz���8l���r�\�h5�K�r]���1$�^�v'l��2��ﻁU��^&E��ǱWv�*uI�sp��2�:=�&�J<љ���W�L�Z�;����Q�m2T��[L�|�J˂I6=��7|�[�/��%Ί�p�kx�w+v�Z��	����niفC��-�Ǣ��	��I�㚹�9\�k���t�u&��r��r׌�r��
u��5,�yT�lA�b�,��m�~�㽁S�j�����z���&��'�\��{��NR|i��:�x{���e8@��3}&���z�y���A�x�a���=� �Wj	kq���!Wt��,C�U|Z�7.6v=]9'�h�x�/�¶>RA�w?��m'l{�9o�N��/{���E����Շ7���6v*���!��O>�$���z���	N�ä5���s]xk���#�3�U�@��Ҋ�!e.�nv�����Sfޖ�����];.�a�}:��(��M1H㗭�y�k-ǯ�gwQ�Co��,G��Z�v�(%F��Aj����Y �����͋�7�zv�=��UL�/ ��w��-�1Xn�{.%K�o$y��|��6>��)h�7��"n��W�m66�wsr�r��Y���ׇ�۹<֭�5�K��?0p��lȚ��;C��i�'q�=ǂur��'~XwW]Ʒ]a� �}E_K����1�q�.[eˬ.��<��Wpq���c���2�G��(�n��I�g��y �.^°}٭+��8�P%[�u�?EE��ζ=ƙ�����]�\P&'+��{Zz�
�E׹�u�k����:�`r[�i�Z �Y� ���� �ё�m��8�<ͪ��}�}��Cqx㭱�h
��.c^5rΫ�3�kpA���|+�;��v��{���Z8�N<�u����=�;h�_q{�N����ڻ;��R�}\�W.jVQ�]a`6QZ3{NR*�Ô�U��u����˽	t�ۼCk�/��Ő���%���Ĵ��ɥ�mЀ ��>�a����b���X4X{�w�ƮԽ��e�^�G���o���!�MT�(\�h�@� �h� ���12���!�gY,��BL��T.����wR���e�%6S��WZr̪���뜼)D��T)dE����������"I(攫H"�4��YF"Hғ���էJ�!5H�NTʣ �Q-,�ًC�trNUEȹÔ&&vF$�kYtjY�2�^���*��DJ0����)IYk*2�UR"�$�&U"���rZID���r�SD�0��bs5!V%ȒU$��g**I�fu�Z�&�+B�hV����D�B�F�b�di!���,�Ĉ����,А�U�hQU(�ӻ��%AKE�ZRI"��ˤR�uι�pԈ��U���Z�a�f�VgÝ�:a��"����ԃ����	Ee`�Y�DL��9��,�)de)�hXd�dT��p���P������f$���D���2���������N��&a�{�,�E;����smb�F6���g@��s_���Q�����b3���n�,f�G&*=�ptsF�6D��[�����kv���y��]����O{BO�ro?�x<Vˤ>?]���P$��:|�~[y@�C�G�<*~v�w��ɾ!}�n��������'�x��{|�۴�zG�����qp�z�&{p��5;����;�{��yݷ�'ӷ'y>~��Ǘ��o�����zL.�Ǐ�Ŵ�I���d߾�����`���}�c���y��þ�����
��+�&��������?���������"��~��W�ї��s���w���n�[�oW���'~v�����)���w��y|��N<'���o)�7���0�c��ô��~G;�[r���~O��0�����}��ﾁ���c�S�M��mv���1vkv��������s���ؓ�aW�	�	��׾��7�99�\s�w���yq8�������P=$��=����	4����?�_�O����\yw8��8v:���K�}�e��rW�����k�p���bW������Ϳ��o?!���[�<&~q�}�Ǘ]�90��;�QC�r�>��?[.���}}�(Rv����ޭ�I={�����o���*2�g���١����ݰ�����_#�[���\N|O��{v��;I�7��ӷ��C��c�}B};VT5Xo020������ݼ����>���`��Y������:�����eS��ە�n�gC�����C0��fkI���i��ÎM������+�8�\�q�L?���}!��!����;]oHy7�y@���;^}��������:����18��|�x���׎R^�6�.{�n����˳72P�����v��;��1��_I�~���='���7����v<'�xC��o�<S���λ�n=��®�x��<&�������HcĠ}I��O�=���˰���S<��߷�p���UX�*��~8��M?��S_��{>��.<���z��v��?���zO�q�]��~��on�zB�z<~�\Hzy�O�8����]���xq��Ӝ<[>�O��t����M����;�'d���=X;������ rN�ǿݼ;��n@�������i>�xBM��zw�����N'
~�}O	������|�������S�?u�&�B����� ��t�����fQ�-fN�}��c����h�&� �׬/�F�c=��v���nDw�f�6
c�2�K��hen���~a�
����
<��NA��A��c�vGS�Ӯ�,ʃ,K�$���L�X��V4�Ç	�q�9�}�Y�#s�sTw�9������N��S��A��O����w��~v�[Oĝ��m�������k��������'�o����C��<���H{w��{O���߻�`��xvb�hvvoz��d�;�4�oa�ܽ���0x?��2����̝��z��(����y�#벛��7�P��}��~v>'�7;��m������>�_��vmv�@<ݖ/-,�pk�|�V���/����raO�;��ohHy>}�x����}O�}���ԜN<������v�i'�1�7�ӂq�!�~M|��{?�ˏ'|q�;�]��w��<�ڐo0v�U`p��2jBuT�����w/�����������̝���<��?��>����<��}NM��>'�y�㼦�ˤ���߮?�9$?���xw�v������P�s��}Pާf�of4��b�X����@����35��_��`x�b���?���~�ǔI���;���<&�'�y�~�yN��}�w�V��O���<:v�i��������x���)������Ǉ����uٟk�莩�9Vx���N��\r~=F�ORC���ۏhs���e����~��yw�k�����; rN��߿��o	��÷=�1>C��Ǆ�~~������w4�LDI��k�8#;;��90�?s���|O	���V�c�|w�?��|xL.�������|q�9���{�ohI��'�w���o�rs��~����q'��ݼ��� xK�ULW��TG��M�j��ۿr�׾��r��|C��\N'{q���<	���>(�q�;�bw�6ܛ�<�����}C�>��.?;�ra~}��>'����_�r����}��Sc�wmݡ����g�b��w���8[y��_n9�N�c˼;׋nq�����򛐝�㻴��oh^w~�{@��É�O���~v����
ԟN�=~��aM�	���m�<��N�����z]���P�����{���Uwg��O����m?������������)�����c���������< xIߓ돛wx���>$�ۣ�o����lw�$���z�(Rw�k����?~B�r�=��"
MW��%}�>Y`x1	��C�k>ٯ����ݥVzm��^ d` �ڝ�i�j�R�{3�ވ~�gK�W^ݙ+i��x��v,����)t�vh�'Gk1�Q�̕g`D�#�1wA�a�#�`��j�Z7l.�dx���NYl�q�N��n��}La��ȟ%S�h���bJ����"w]{�<�)��n��ZчǤ��jS&���3��ք�5>�e��`W���o���G����(U��9^X�z���_��[-�_13Bi	���rXֈ8ք��2ٔ�Y�O*�`��,6�hc�D�k���$I�ε�g��y��Lz�;���5Y8����[���\]Ƞ6���S��w������m�=�������W��?<LS��x��k�k��@*Ӟ����4��:��b��Q�
�U�E,cG^�ܜ2�C/,YQ��\3���,�L�tҽ3��u�<7/�:�m׆1�5�'�꘾��xy{w�0k8���p@�����0�����f�qJ=��H��>���\��Ry����2�̳��LQ��jn��P��cT�p갮���e!Kߊ��g��I�d�a�R#B�U	�3I�ylP����e,�j銚A6�xv��������#H�ȱe&;����>ܳ��C���r'�)ѯN��g*6ƥ�-IK�*�"^�!��Ɛ W���v��RyH>�z��]�����]�>�)�p����WwlxG(�*�j�qaVa�Q���0�u��پsR�M�L���ά#��J��D���6**�b仯j,#4y\�&+-q�k#0i��6oY=Xce-K�&�Z9�+���>��R�Ї}gX����O�"2�3Jm��a���
H
-E�z}���Z��I�������)Eɝ=��vN����p�l������vؿ.�Wv �E�� �>E��;S�y)O�1D�D�򏄣�h5�;��R֌.h�jTl�ƙ��H��y���$x>�*�u��CA{�x�G����I1����|�3m1˶���O&�]|԰��+j���6���0<��� V=�b�C���<w<#���W��
S��3>�UG�ѯ�#	|��zw�b��mQ~���5��ʈ��s�L~(�nߢ��^�tA��9Dd������,�]nN� S��T��(N�#P��������K=�hX��j	���̳΀\kp��������Vx<�xJս(S����?$�»�eN�t��b�+�ykM�Nd�'����Γ�aYo�����ׇ��I�����Q�N����P����"]X�J}V����np	�����?��^��O������~��j�z^��f*�Գ��yj�0'X�d��4����w`�]���4U-��5?xͻ�������w P���ƴ�����.�˻�O��Uŧ���Rh�o-��3 �D	����7Ou͇,h�C;O�*���{ܺx��)ȭ�XW��H��e��2q-�S�-�Բ|�7Z�(���:�{u_%��[Xs;�0.�E'�*"G
�<=�
:uߜ�w'�~5ᓽҼ!�}u�`<[���M�nYy�s��f�t� �' �k���]��J��3���u����d��xCAA��*�-���s'���{�o?R0U�h����@o��'�(V '�q���5)�=�i�c�U�Fz��/pO�C'�;\;�v죆~e����T<_꜅���C=��ЯXV%�+M�Y�� bŵ�]2������Z��&H+���=]�h�j��ʔJ���{��0�:Y�h=�P��.�K1��M{��Σ�]~2�ieF.{=\��#��P�I����DP��<��:֌��ޱ��p�L5���d�c�NH�f�z6�=�(5�R�Лw�`����u.�i/N��t���b���zt׉�1�Ճ��L;�]��z�{�$Zty }�>+b&^�Nz0�Ŝ֝w;y�}J@����4;@(Wa��a�W�Sv�&y䩹�����ˬu����p�%���y4ٶ���j�M*�/�em��˪����C[�OpcP���K^����u���ƀ���Xi~�z#�Vj�P笾͸�:E�﷌����"��ǋX��ss6cl���i�&���@�Ͽv�xew�8=֒9T:+_��5�j���8X6�[������$�f��8q�$�4������/L۬`ڏd�Wmv��DFe��`C>dxH��}�OJ~�ȹK��gxV�=T�߆�Z6��LT��׊)�e�;RQ�[��|w�>}l>D�c;����g_����tS�t�p�Q�>�d�D�|�d��u^�x����x�:�g��qrz��\��������c��o�Ʊ�����^�_:
���l�y5�V8L%�m����Y�ozuM�@�����x�*�J=���aB�������Jx�"�`<�5�w^�}b�Q�Th��ֺG���0����{k���+x�iU���޸��31~o��x�)�����E��ݑ�}L�f�2רo�~����:ŝ�a�M.�_9߉W;6�]z�j�u��{M���
t������)�y���û�y��x`^��+c'��gW���5���<3�=s��^֬�
�9�������F��pR	</�H{�j������[G�Y��0w�s$��W��,�N�'^c*�R
K�/������F��/�V�6/��n�>�ۑc�VV�>�7�4kѴ���(�D춣�5n4\�L<����[�v���(Y�H��q����m��")�������^�y\�C��f�C{V�\�<�H�X8mT�IM��)�!Ɗ�Q�yDd�kF�L��W��H�Ł��/�!8��x�p��Pt����P�iL���T���r����ݸ�:��$E��1sdVʢBbB���Q�~_�]n6����7�`>�am�w���p�/~�Z ���~�״[���s��q��S*Q�vc<+��՜Wu��]�^a����a�A��"d�.1(�iZ�>�[�p�J̐׳� Ĳk�x"�oe#��>��ǡ�6��@t9U3�
�ؗ��"/��G��]:^˃�Z��=��Ys��˻�����p�h���|������Py�
e�)�m���4%�cLFc�t�bRlRN/kN���*�ܑ���[�?/S ���<��	Kzg�y�� �ɴڌ�(�"1]�=:��
b�vx�%��Ņ�
�ː��>w�t�����90h�[�
Ӯ[�̌��M�s5KYV,��j�̘�,�M[�LE蟟 +��Hxm��^�jz��`�kn��.�ם�p
"�{���N��S6�m3�]�e#�{�W�P)S�9�c�=kڶ.��l�E
�(���:�tn-ƈ�����<}���d��1��{�ҽRO+�^�g�fX����V���}x���=Wy���RY,oV��w���22HV�g�zN=9܈B�� #�x0��q:��Z
T�皹�3ޝBK\<s=t�e�>���e��
b����*l@��1,�p�&n��k�~�9�۽4�����Yl�=ų���8g�p�7ڈ�?޽�h�����Pb�ty�Nd��'�;Ӝ}�X0�v*+���[؜0{���Z{�p�{ʰ9�:9Ky �]J�N��Ε��c'p�4�Cպ��*���6���XY�	�FScJ-��JC I��q�>��$N�6�^ey�J�����+���`puD�!(�
������A��mu��5}�}]��P����17�E�
�;S�2R���fT
�� �(�rC)b���}�j��.j����^��Xu�MT3��������^B
���ĺֿj$����W��Fv>H�%�ፌ���b��-���kFg <�w�~�6.W��!�T'�J�}c����Y*	�7F���G�[vnѪ��=�<��ύ1^B���o`5�����He�t4��^vf>�P�Vw�Ba9(�^{u$�W��<i��Dܖ ����4-�b���Y�ʲ��$ݼ2[�u��$�2Vhπ�!���q��O0(��OuΆ����ou�N8:d۶�(p-��u5P�1�Nf�x@�EP/v˘��aC<���_��~H���SV��|ʈ���A��8�C��v �Y��{u���9�^�W0 �Z�8���.��Dվ�:��zG&�̿�΀�[�q;1��!��O<r]�⒁�M��mn�ͪg^3-z+}�zL_Ob�}Y��`7��쬔V]>@{]�RMRm�9C�X�p���yހ+�� ��4����NI�Y̯y�_�~G-��Z��
�-!�����'d)M�[{����������tM���.�f8�2��~SR����ֽ$� 52�. 2\��^,�v�}Fa��)�M��e�%j���)��|e
:uߜ��qB�OzQ�OAEhB�>��hMx�RLJƶ�oV�V�2u�p>t�솦i�mB��{L�5�^�5�1����D����V���]�� �=ˮ,u 7��'�X ��ioAqʧ3�H��&�n�'��k���"^���0m5�L0C��%�Mv}6!�_<�Q�^�Gf]w����P�.nm��e��9��,źm�:�Z�`�=��Ҕ�!��hq�Hi���.����2��yݬ|�-3C�M�d���C�]�+�����̚�_�d��FG�֦V}��oSN��rؾ���wvIc'�X��[�Q�ޅ/���G�趰���&*"�x��8��i]��\,��}���-��Ć*�͡zFC���oy���2���D��xWR¯;U�/��<��;xS�{�x)K��U?"�v��$�3W���0�ȿjz�h��ЧH^8�m�x
 �`T��!6�-���ޖ����o�:�|�O<�5=vpz�=�8U�u��(���pK6+�TvfKVǐBg���\��ʇl��"$�l��#��4D�[������CYfç��j~���[pp��y*�ܥ�����g$} ;��ɾ~��ZOt��{�8'�E��H�u�z�5We��`۫|<8~��a..G���ښ[=��^��������jb�~_��rT��<If]W����8��B����p��֜��%$������ ��MJ�5�<{�{{<��^ˬvHX��Х�@Y8ֹr�h0�^�]��~x�*�N~�=A�B�,�%k�있�O�l�[��a����Ji75Z����=<�v�8W��������ٕ 4X���@p�/��{��~�5�	�{hQ�~.K��oH����kǙ��N�O�X%������ڪun�J~V˕ݩ���Viѷ�U��`
�D�����X����2��j���^�<��|pL��o�V� eS�=�b��ң�`}����1w`&��Um�`�wz��n�Ğ�cf3��9a&�.�����8�R��bIx�w���+�.���^�'gZ���1�<2we�+��y���;��>��ķ��ق����1��̓(�Z�ǉ՞�en���܃\�xƱ��s4՚�/F	ic]���wu�`,�s�TE�FQ%9����F�͏ѯI������	���W���ۤ�,jI\�^�T�ɨʢ���MOr��6�ƍ�x�Xn��t�;�u{�J��9Vӡe��V�1�;i/�r����q���,���ٚ[��Oz���"�����Ja��U���5��@��ޛ�p�u;�V1��f1xC�1�tN���¶����[�ʳX�ز]uL����AE�e����^���1�̮E�R��q�ͬ�54Ȧi�44f�NK�ύCWxC��� |r"��з�8[Y�m�wb���z=���᷃���,C��d�a�r��Ґ���4%R��}��F�}�5D+�_c1�m����G����M����Ɇ\��\�>^����c3�ݞ����*3|�GѓP�z��a8��' 2,aν��G���)�KKW��/�,��ŀ�7�*��m�+\�W�"B�_
�c�O1<�X�\u�������f�8P���y �o����|`Yծ�^]��r�����<@����.�/�0���q@7!^���FM����T���e��I+xl�R�W3v�$9��Ä>�RK�-�L���v���<�*�w�Gj�O����[��q������zoev,�	(��U^����>�.;��ݾb�.z"����]��h��"v��oxI��<�}�d$w����;�lP�����;O���오3��Ѽ/d�8�V$y)�`�7q.����1n��:�4� ��9�>
�Ş@�P/<�籟���i)�}Ҋ@̠���5p�����r�En�;��b�2�Nch*ýT�%=�"7�#Ñ���ޑAb\��c!���k���,C/�Hy�[Ĉ~�*��Y���\��b�R���9����{K��&5��/-ޯе�W��f|mk%J�� ƶ�(HeI�TƸ���Zn��\w�����W�b�ۺp�kY�}؜~����\,q�W�%��jo-$o�X��h��&K��C�s��	Wf�9*�}2��<�:�*�6��<C���)zWk��o�PzOS���N��
�W��g�2v�H#�k#G��
����c(%zgzʿY��R��
�u����ɲ���ah�X���I�{���{�L��)�=�j���6�5���3AIsR>�ڒ����9�>X�>��zh��\�5�8��Ž$��۝��$�}�{���TF�I�Nd��qũ�V�J)H"���DI%���AU\��Qil#	
�g(��̐ڵ"0�ӡQ���%JP���VXQt�Rp�Xg*UUK�Z�*��( ̵*�ȳ;��I�,�+�R��L�%e4�*͔GC3�Be'B�.EWD���DI"�D�u���Pr��۬�m��M��,�SKha�WV�\��rH�;��Va&TNt=UC:JU��A��� �$��B5�%R��*��"�*NU˚)X���B �H���+D��$����Q,*K�aX����ʨ"8���T�K��YI�b+R�iXYr4��Dp�i)e
�R�(�J��EA
Р�E�$e�J����P��2�VQ��U��顈z8�.qE6r�̊$��	k@�R
�T���8U�),$(��(��p��"&��CEM	:L��G6V�\J���
������B�$E����0�H�$��U 	�h	@J3Ĳij�%j�� �v�e� �]�m��W˩w""."%X�E�R0/+0�ㄜs�5������;l��G~�7��ԨS�B�7�&�c%S�p[�d�� ���a�[@Za�r����WnU���^R����c�`�2�}�T������+�j�$��5+rVEL�A��^�g^ԫ"�I)��Q���m�|�oW�ՆB�Ucc��6���%�cJ��X��I�YL����82��1�$�����V��s�<	gGe���Z̖}X��'ISTUce>F'cE��Z�ɤXA�;.C\*W� ����QW��/�<������[��qG��+\����4�y`e	��u�d��ae\�Q�f�D'��6}s6=ɹ����ڞ�?w�m��$-�1P˹�j'r�t��g��	z�)�����KL2Y(�Z�2���iѠ3�9*�J�͠���ٛ[d=҄^���ę���5������U^�`Shၦ7�lМ�|�7h˹B���
���Kt�Om���	x<������"�G�P�O��v�ٗ/���[m1*�br�J)����Ѣ, ��k��_���u�z��`�I��,�N%���/��H/�7W�4ؙƜ�������F�L�*��K��'o��S���8���kiu�3��5Z�-��m���a�O�uJ~*߯�8�w����ӓ��(�ɋ\�O�Z����Ϧ�^,Z��C%���f���ԓI������7�.��A��Y6���iz�U.�� Ά�Byw+]���d&h%*1*��2�`�%��QN[@��Am/SQ'ԓ�6��ꎝ��Ռ�"[J*��VSYgl-eEܺ�Ճ:��*��ο{��}���%����֦(�&�u���eU6
s4u�%7g��>^�k�C��x){V����gL�l�GoX�ڕz,�JMF��*�\���@�^g�O/}G��h䬿:ʫ3�j�=;��W�h�y�/�<�����03Vr�~�:��P�BvC���\|�����ҥ)�}Ŭ��=Y��חo(�i
�����m�Z!�e*�����"�;�O�k�Q�0���7It��<9X�3�S&�{?{%�����)*frS�q�׸�²螔�.��H p�6*.�4O^�-���U�Q�9���9z*���;��{�G�[#��N�z�ؑ����WX�d��E_�����2�I4�X��hCf�sL擪b)�*O>P��;HN�3�=���"����do=��'z��m����^�JlE孖�4#Hh��34x\��	3�|�M���w��T��5*+U�*���[�-Vr���1y�j�ۢy�'��A�r���)!*��̿,�Q&[���k��q$jwa���+Cy����(�~@b�o�~5�=�V�r���>�m��ҩ8�2��oYIZc&w��v2����(�ra�C�r�G�Xq�s�})a��e/�
�42�f��j٧�e��R�7Ud�ʱ��2�]�
5J 8��v3<a�e�}F��˪g�P��HӦ�ī�Hµc)�[�"�s�R6��ې���<�r���mg�MY�~]A��'ͥL�J�+u����l�L��گ����]�]�6y��8ӟգvmL3Q$A^�Ec�!��.&�K[ds=!��^��!^�w]9�S6��ץ�x����}}��ڭ.Q���P��	���\3bYDV�����=�A6��oӔ�;wv�L/#��#����{g��I��>����US5�\	�+Ɠ��t(^Ɛ.J޻�&������o3y�X�>���N#~m�:K����/��x��;~ɹK���:�Y�����뢂��qͫ$\�T�X)�i����z����)�e�Xb�C�R��jDTZ�!397T�=�)��I�E��ӥQʙW�����ߕW��;��D�QMS�`�k�D�!��'��(Kg�ˣn�S$�M��n�"���� �f�u�V�.�K��4據d)��R!���~
�Rw���s&^Gx�W ��S~������NX���SuAE��7��N���ɲ�ăv��e�l
��i�kT�r3NAC(Q2�bM"��������ӎX��RS�B4j����O�Ug/3O�,޶�s�m?4��'��.^H�ě�L�b/P���i��!���.�sȚ>����HQ���Q��ۜ�ةd(����J����.��`�Ľ��؏��Ul׼��uh���4����{���3QrDܩ�F�69}/et"9���I�{����D
�V�h�l>z��#��q`1�@KL��u�$���a�=/�A��q�&�x�	l��$;J�D��aZ��Vs#NcHf�3�2L�_W�}U��1�=��j_7�	=�Z`ոgF��V���[�����S?{���3�/Ef�|�kk����6�-D�E�e��M��,-;�c�-��w����$�*�Jr�[v�s�){*ܪ1w,����h,v}p�}e���'N��Z� �v�ĺ��Z=�=]�1�[�f1E8U~�Zi�XݛSL�m��X��A{�̻[��p/YԴ"��W���H��0Z0a�歠-1�"�Zp�����<����������<����c˙>�|��{�T]'�%�������^��jd����+p��*ȹ�)&���h�Ӭ�3�ռg �GS��7R��=$NL$cs%ͫ�V<�O��eF���G}�a��iZ~�͝��2��g��Ύ�U����/�ӚOl	v@bX6���gҶ���K&V�C��B�z�<�k{�U�/�sיHq\T��H`��8�m�z��׆=�����:�?n6����(6zxf����(.N�8�N�U���W%�̵�O�S�ø����G�KMA���ο:j�FW{��[�-Br e���[9�ڽ۞����CsO8..m@}~�9���f�0�r���I���e�i
hozx:<�_�{e�������,E�Y�H�	�2�i��� A�^4����EO���2�����b|�&T�2J�w�7f��R]����xmr��%+^�m ���t�4dak��ãκs�ɝ�Ɩ�V�weR��~(�S���5����WM�i�Nk�1���8#/�e ^E�|Ñw�
���
Xu�=�T�an��lTѐ�D�Ѯ�m8�RWtF~~M;����G�LU��w�K�����ؙp+L�(e;��j�ڍ1�OӋ�>b⯟�+��ڬY7���ͦ�b�+e'ʆ��D�ۧ
��kd�[�an�f1*�ّ�+R]���X�/g.gIQlBƓ��s���UrZ����"t���5e05�gp*eEܺ��}� /����M���׽7}�d!�4ꑦmLQ$K5�
*ϔQU����O�0�s')R���;���Y�Z�`JN�?���w=�T��{vy�,���%���mi����=7P5Ƴ�g�n�՜����q�#|�LT󇺢�������'�w5fs���r�n:n+o>��Ý�N�u�3�ʞ��o:ά��)����33*�$Vnv�}��1<�����T�:f6a�#�lu�K+�wOh�c�Dt�PU7��7գW�76�}=���β����~;�ڬ�����ϯ��ăE��F�Lޗ˷�Ф���>ZZ�l5�BvCݎ�w��*�!�]W��3%�ii�Od�uv򒶐�!ͣ.��cP��;	�9��=��n��ޮ�X�5ތՎu��t^Z��'s>�8���V�R^I��Pql5���--Yp�e�6���OJlT�SC2צ�i ȼU�	6��R}7�h�)��e�V��KY�k�3��d4��R1t�#b�6oQ�,�pOV^Q:����s����ϖo;����`�Y��T�S�{��׺L^��x�z�c��D� ���I���֮�,|��Gj�e�9�I<�e�p��Q�֫%����7�2�j/��A�wc�t�	E�7�竏V�Y2���5��3�8���G��c��Nr-I�cRa�I� sox��R�<�� j����x��^���/w�nSőͳ�=@Ѕɴ�۴x3|��8��܇;f5s&��Y��ˡ¯�[�/�1���C�*=S11�K~�7���tYNɕ�kt]���֝�j���O��Ps��~'�&:��%~u�m�V4���2����3i��b�ϧ�Ui#
Ռ3O��j\DU��5x1I��diq��h�[�e�����QeVY��!Lf\��S7$���ܝ�۴51���(�7^�[,�MHݟZ��H6��i6�Kn��hM����/B�0��X-��"��l|5p��QO�6r��˫Sx#�7�B�G�g�����P)f*R��Y��L�>Y�'�ү��&���CK���bOdyW�,��޵�
H�JK5i�j��8ϳ�j ���l���i4��p�M���>�qd2�JO�B�a̲2賌E��g%�j1�	�ڙ��xV�,ϫf�������4�i9�e{����Y��C���{��#g��N�������T{؝�E��_��R��.,}{����ffYǝЦ�������^7�C�F���/}�onW�`�xB��Kr���8�>Sb�	љ�3���˨���������t�)	���L{�`����� 2N�&Ȼ������Hln]�3�i�����Y����C9��7��y�Zg���\��2�n�45�"|6�x�s��L[i��J[r�{�����r�8)"%�MJp�a���Y����O�h~!������D��Z n�÷�������k�1&�FS%��-�5q��C1W��R�/"����)�o��W���R��Pr�s��|����{�MW� ���xf�)�U�I���&�L&��,щ�l���[F�m�h��5�d�ʼ`�hRل�Y�����:䠚��1>�����y���u3�ƻ7͇K-�M� ,H�b����Tj��(�� �����=6�P���>Ƕ7ڵ�#�},�o�ɬ�+bue��fI`�%��2�B�{��;P���e�r�|�FNOR�%�$�+B+HW�������0Z=��@6P���yjN�E4����3R&鬲�8l�E`�2�}�YAe�N�K6ǅ3�޲��U�Ō�F�Z��u��gr�!`����rf��d�m"R��A[�]Q,k7F̭�e��RzhҪ�ci����`�s��� �^��[����+	�̸r�U~��û[^��;������)��Sr)�{Ú>f�{��^�{
qj��w_4�3L閍��+r��ڕdXPJy/	m�z����f{�ϗI�^��+��H�}9-R����WD�yjI��>���s�ֵ^�y3k�8��������T;
𣁑��[���ڱ�Pr_\�t��e2�a���2�A�$BFÝN۞u�y���*�� �T��wY��/��sͶm޾�:Mj���J��2���[@c��3��T�i`�n�s�OǼ�8�Z1&Қr�V@��)�JkZDRצ�#HK���b|�Ǵ�3���%v���^��۱
�E�CX�a��E�-{��xxaQOW;h�ܓ����W_w�!��nyZ��C8�[E��s�+��d�?�P*���:m9�55��U�lW�~8��򴺑��9^�矯z�v�[R-����%&G@�i25����+����&/��뎗P<調�r�5so��/�ab�Mz.o���x^�_��cȳ�m�Ц����Ժ���.Z�6e�]�!�2�މS�T`�92�r�е|�Y��b�ua5��@�n��b�+Z �.�B�+�L���R��^�4����+�Q^9����>�q7���:0�G	�� �|�wV�XzB�<�L����U��T�H���u>ZRq{��Ls��j��U�ח�k%�z�tdO���k�@���Q�<lfeޫړ�%[�:�o�JҎ�T�������fAb�XD������dL6�;w<
��
���U�{&��q�ܐ������N�|�p�1�0\q�[��i��6��oq�[�K����ŢB�����8w]��z���tѨ���s����Ğ�7[��
k�ۍCF�GD��3+g;���<��o���[`Ԟ۹�3�#쨭��n�>ˁ(�xc�5�{j1��e
��S�w2j.�e�%����Fr�wT��y1��T�hh�X��;�.�Sp�Ī�==J򑧉�p��u��gnl��)adIE�c����dYwPE����N�gi�%��AZ��>�]�DP�Һ�ͭ�GM�p�x��bl3���Or�j�賄+2��={{T[m]P���=A�����t�*�8���p����wBS����L���d9��M���9[r���ۋ��cS��24�`�,MPu�X�i�n��:dU�7���">\5�;ޥgVaҟex�*���W���m�t����泄,|�m�Ғ��7�V��u[�ڨ;u=�i��>�lj;��SF3�~��[���7�i�7��;U7�o���)���[8�'4�&g*�^��{c��y}�Kc%�^P���vPm׷��PK��D[�7M�Ԇ��Z'��� ! s��E�=V�n�IK�w� �A�\~y���VRO���L���Y\f���b��A���@6�/����^{u�S����m��ி�b��ܳ�WY�M���b�Nw]��(��0���Q�=A��`�`8��w�t���,�.V>V]u���-�f���@`����,��e��d�U������Z�!�j�!wC7�1�x;�t��3Ĭ<�r��52VR��6Xv�$;�h�F�썜~�{*���0K��qn�(��\��6�@V�]����x�r�g��"�
1nT/���,.fJ]ME�[w�~��^���0	<}5K9L��?�:
���s��6�i���c,�jV���{��ޥ��7��b�|D�7vhׇJ����x9u�k,qE���ۚ��Gݢ�ו�K8�>�˅�E��&9��a]���V��p;��ǈ��n�ྉ��Yq}`�ɬ>6U�D�Κ�&֩�9�˥d�T�jL(�o��i^���VJ��Ʈ{|��v�=m+,f�3[t&��y�^^^��m���۾|x���J�EJYXU�2櫣�Nb�*�+�A�����&�ZX��a)JQ!��\ۻ���Q�l�$
L4E�9,�!O7*�2��B".Q�SYI`��*QW%hE�(�պ����%r8�Dh�
��aQ�*�-LN��(�Zi*Z9�s�t(N��".p�+6��2��D�6���W*0�p��K��B��B��EjT��$nt��V貜������Vh�
#�Y��Ys�G#�Q�92(*er�D��G�W�Z*̒�ay%4M
�0��
�֎�iЂ
��+�֐N�VJKQI3)�r<�Ôx���nW��6P\#��TV������e�u
�.t1��TT����9VK#P���L���w3����"��P���J�,;BNs�"E)wnE:�.r
L�ȅhrO]�$�.d2���dTEK���r����Y`@�)ͱH2*e+Fޜ��S���b�rƃ�����4.g��V%�&��$*�����p����L�	�Ke`wj>�7��{�g�E@��n�ݦ��Z�����~|��qW�����YW�\���:�o
��s��鵊V��V�c�/��X�j�w��(�!�PiB�F0}ە:������[��Yj$���U(Վg(�Y�rj-���S5#�?[�粽^
#��̓���9(�$�%��EbU�i�ך7��1Q������~��Ϙ}{V�o�$�d�2$��{Qe��;��ۛ���@�Vj �����0s��yŴ�e!7ō��v�so�-��c&1̕v�0�*���$�l�C�j>F������G4Yi��;��F���-��p�gM�Y�p�uv�u(X0�Q�E��h6D�db07-�u�NV+-�3�3�Wh^j�4擢�֕'�(H�s�n��N�we�9��m�N��g�xjeVzӝ�)�
x�%6*bz^��� %�ae�5��5#�\�WܻOB�ِ���&p�V��{���Ϩ�ٶ�8�=y+ǪCSA\H��J�&���6�M?���ue�T�_�m��m�Mfε</8sN�$HN�k�F�'ӮN�dn�ݥ�pu�(պ�k/����x����ͩ�ﾪ�����ȭN~�����=v��9�,\U(��i��KiL3gS�2�t���gl�[�i���T6�hS�v���qq&p+��鍺��2SIi��#���gݏ}���)x�=m�bO~�V��w��y�\��V?)�d3өC��H⥰�*�bSR�X��`���܉h���F���Ƈx:�Wk�\�}@���fr��􊧋�2�3��~'�ud՝<x�N��g�d��j�T��>����:q��&���/ �:l���d:��2L�F.�m�
ق�f�l�aD�>Ҋ�eV1��m�-�aѴ�b��^�lo>��Nu�u���i{zS;��s��ذ�Cn>`���­5���c�խ���E�Z���nZꦙ��u�1md
�cgj���IԻJm{����(��,ys'�O��u��eJ����O�(���un6�"z����҄Qb���%
�7���DM�D��PE�g=��W�ڕ˱���ڽ�R�ֱ;dѼ*�A�:�wc&�A��eu����\Zj��i����B]�`J�tW;i+��S��=�4m]�_)�
(��{��3x�P�%���Q�R�nʺ�zZm
�JMi���}�Vrn��̈�Հ2���:Y-Sjafk�D����'���c�I�۱���oN�9������)`�Ke�����Վv�O��)�
���(7&UڧV���աPx��ː���]�y�'}�f�)��L)�h�j�KU�]�8�`u�v�>��{eQ++���Y�y��~E�Q��vy �(�T�������׶�#@Cj���b�w>h6�Z�DE�3.O��&z���E�W�&�yi���J2Q{�[`G��,�f,���\*�S�bX}�{۩��h�=ֵ>�X��B�l�ةd(�kU�MM�`]�צ��J��/��{���*�^��a�:YK�R�:0��aZ(,�Su0Z��y�}145���{�M��s��V��k-���]H����h��uZw���~�?��(�cA\� �Ls�d��%?W��w�C�G�d6��V����s��8������u�GZR�=�������� ��7�7��֪�PޖDj��ȹ3�N|�:���H�����'V�j)5Ӡ2Y�i�+\�lN{����މeM�U96�;��z�Ya��j��W� ����[����g��|���t�%�z���S����IX���H�hB��ZiPv��|+A��Gkq5��$g����F�+�^�ne��w2�C`�a��^�O�/Pq�]Xq�ڦ��K�]lQA�����{��{w��ʞۅs�]oш�,�ן=��UL�ټ+oN��o_kϺ�|�n%�g��2wA�n�Cl:Ɔz�%�NL$6��ͫ�EcŵA�0>Ͷ�v	��x���3q ��>F]�Y��z8-��j�0ֳ	9��j���͸ɣ���)��TΥ!,u��Z���ؗ{�RtH@�b�U㹱i�J�(�p����8�jZE4%I�����WY�Í�*5�MI�sD2Vm�����7�F|ې!��x�)�l������̼�{w�<�S0��m͚�l
� �q`v*n���k�*��
L��u�l�4�#t	������m9��<2�SL���w<|�r{ɡ3nhe�mX.��]���o����wd}Sz(�Un���d:�Zn���%��5�.�>W+zw��9��������'Tf�)f����s{f�A�Qu���L2R��Z�7��&����wt�x���j�%����.�R��~(�S�U�=����O}�إ�)7l�j��Ҫ=`T�6��Qw�Э�l�,�|o��4��yZN�x��>ٳ��:D���(�����=rb�-��\�՗wZ+V�4���ot�kN��uvu��6�J��6VLj��(�N\\m+1!dT�z|�13��jlbSZm��`ر	f�:H�W�����*.�LQv�� Nn�9.���G6.�
RЙkg�X5D��w����k��]����"��Nk[�w	�w��`�6WM�[�M3H�j-����|QY1&�TU�f�[F�Hl��X�E>O��@��//f�ꪭ��a��to)\�����D�qY��mz�:�,yu�G�e�5��sը4���(g!]�~�k%�C�y�Kl�:�z�*R��-鋅�KZ�j	\�h;D�G�N�Q�xh�`�3%��+ď��MP�aӔ�b��3��,=V���1ڕ� =��SG����N�o��Ԗ�C�5�i�V�/�\5=�r�7������1	���jk�mۢM�RO�Ф�����i�X�c=%�+V��/Q�1:�,��*�����l�[:�yd���A�s���4����+��#cZ"�s���ZpQo�U�^�<�����M	Ry`e��.����6�S�S����ix��To���w��m��;�:��6"��u�cJ���S�N�e���ɮ���h�v�4�gyf�YT�y������_
�\�֔���	��{֫:2x�K��R$9y/�{s׏�_���^�ӽ+�>�d���[�g�ǵ�(��@e/Bu��z+�k�X��o���X�Q�,��bԑ��qS-�V�%*�F�]��nFRI��Ƹ1��Z�/��'3i���o��S9x���_O�e9ZKhz���0F��7�f��F�BK4T\�F2����f���bi�Ӧ�bU�i�dlA�W�8d~I����5�`/����YF:	[L.�J�k]��&>F�>�U�����ԝu�̩G]�)��d���Z��:���.WO�����ŝ��Q���we���
<��F�Y�
��='\��7z�D�H�K�o37��3T��ʤ�R.vEvU�DU[!�l�����XQ(KiER�*	��˧v��l
��-{���b̔�eE�όQ���l�D-5��jmi��xz�U.�#�M`�"�w�̏�T�s)u>0Z0a��a�VS *���T�=l B�2�Y:7E���w-���W�ʄ�9���2��:�Ҟ��VT��tJ���L�1��]n�-f6��)"|�:�cn�oZU����G7 �	���3U;j��y�Hm91D+�}���3��{|-��N9Sn��>>��WSև���ͫsv�Y�c�2�ԩ�x#�quᗥѝ^�ez�(h��p_����]�y�w�Q`������0J�.=��k����=4#HK�[MD�t;#=������Hi��;T���i}�U�$��қy���2׶�hU����a˽���#C�<u�\�޾{\�U�������sr��J�zOR��
��k+��F�.Y¶r��au�l'�{F_���1�H�M ��ܾ�����Y7�i���+~�b}��̨9�>�����k�cc6*m9�:�����gY׼zQ�bx諭���J��n�Zk�<ٷb6��.[-1�cr�)���E�em����J�����I&
�9�d��}�Zߗr�Z�����W��x��0��*{6�\.1���$� �c�ȟEE�BOse��a�ц�g��w��Vo]�-������|�^�X�tTy1>�����l���<3b��uuZ�'�A�ʌتx�s9��U�.Ya��j��(��BL\l�c���ƣ`�e�OqKu52f���wUxĥ��$�j��t�d!]@��IcDB�pj�l�&�m��������5���H�|V�B(ׂ�T�-��"�e�-�,f-���؈Kg$��t�X}&Ikن�w\��\����=�sJ�v�܄��l�Q��s�i�5��1<���@ҩ�t�z5�׼��r���-iC/�R����H�Ǘ��>�,����P�ӓ���1��XDy��#Q���d��/����}�Q��F"�mB��P��y���/��Nج�Drܫw��j�u�`f�#3pRuEOs4lW�����R�b\P�|�b�8+��Fq�����8�ut�Z�L틽6��S�V3�GL��)�&�E�>��/~g��U}_}U��"�!$voK��>O�ʇ!ͣ�g�a��0��Y��j�:�v[F�if���o55]�V>&uI�%m!R��6�!S/�`<��R;�k������z������X朦�^Y)N|�,6m*�hKȔ�E�8@L6���Q����:Sb�"�k�G��(ij2q2��J�y��'���!���ٴ�!��+���i�JQw
�S��U����=[yަ��o�h�r%��֮�,�w⨿S�X.7<ָ2,�7�^���b_la���@Msbᘪ.�+z�,)as*Z��V�V�lb��Q���E�G3t�H��}^e^�a�=G�LU��\3���+ �\4��l�%mrun�T�oUd��f��2��d ��h34���3^����VJ�ߗT�]O������7ɪ�>���.�)oΏh�:�׋%�lg�5B�Bq/;,Z��T�Z��ೢ��؁L�f8����� �#���X�򥯳)}c[v6
&8ņ�"��5y�_\�{̜�x���إ�m�=e>�r��z�)��j��v]uD �{�^������2��enO�f�y����"�;��F�@�ڱ�-�,�#J(��YLb��l���h ��w{8�n��Ƌ��(-��4
��B�R4ͩ��H�d,U��0���ɷ�m"�*W�+M`�R�uߟ�RÜ�h��~oy�-y��ق��^g��6i��T%�S�]��g��L���i�YWβ����:zk��^�Ӭ��b�V#�uF��gG.�X���PB!����g!�P�b��o�J���-Ri�	��S!�w-��Vβ�Y%m!R�Ôaї����D���е���*Ȗ{Fj������N������`euʵ�$`����l��}T�N��b��ɪNu�n5�O�����f�����"���}�7{^�ǆ�	�������k�|�{~~��L$�:�y/�ߌ�ӆmp�SR��#+^�l�M���`-K6�ܴY^lW���c�X���9 �uŻ:�FU؅�c���dI��t��S�#;��Y�hڱq���5�u��Ӻ�՗۴��;���yg��v�5��g϶�H/t���goC9���c<��m��G*���]��Jv�4�w���ttD�N�u��k�cS,uK|�%�R7����5�R-W�4Tڼ�f���0����5YOBL��{7���K�P�Ĩ�#������-Z=-�Y@����j�����˽ý����rzͽ-1U�+7�M���ҝ��Ò��%eXe
É�������ig�jŷ�tsA�8|
y��]�Dw�F�Z�s�m�]3�;�5+�Z�[W@��G��i�����a��3״�7��=0�W���#���
 ΄�Jg<�$�"w��`�]&���Md]v�Jȩe������]��W�x�W��[u�$&�3��.�{)=��3Y��r`#j�sZE5��������~� iwi9�+�F<���s��5��L�v,��q�4�����K@g��!G��wͶ��&*�~�{�5}��qC��gQ r�f\��	k��z.N���
����Ȱi����/�L�;;5��A��Z|��h��@>w��q�>|ؚV������s��n�h���3.����e�4����YL�ԷE)��h{]���2�ƫ�4}&ݘX��&�Ŝ̝3bG%b��r��çd�Tv��0wU�L|�����\�o#W#�5ݰ������s�I3��y�F����\�T�!F�L�l�T�.�5�f��S���̵x�c@�tQN�yu�G�a��R�g��y���{Q]�x��Fx^}��FJy8Ӏ��p�`���uvS�F��&Sd	p��tcZsF�鈤�>��=:J��c;�:�,���2�wݷvp�U�t���0XM�9,�%�K��質���ڢ0
��4�"�+� 'ؒ33(��hX$�H��8��Λ7����U'8� �H�ʎP����v�ى�W�J:4U\�Z0$A�7��D�.��d�ܮ��)�:v�<�+��X��4!n�������	�T=WO�fm{Y�,��].�/S�N&���(=��J��lΜ�}MM���~x��쮴Fn �up�F�f�cV76��pl)��7b�j�Ul�9؀�o/	ͩ�)J�GLc..Y��!7 ��Tuj���h!�]�=0�%m�]Fb��4�Ou�Qs�	5�T��+�vx}8�}a%{��6�:���q��A��+wO@ش�1�UbQ��N�gyÞOr�`�����MA`]ݚ�m�9%���i:�ub�0��2��xu3 Iv`쉝�B{�aNp�&75�2��&�^�g~���Yѝ�a����B�(X��6|�!JU�im��8��˼E��E"������t�'��6��񞷇l�T���&�b��q��V�n�K�R]]P%�~�K��fZ�E�}=���`N���p�+�j�EY��U�wu:&Uӡ'iE�BFdA��UL���"$�J�4B0�N�E˓��'P�0�hX�z�t5%(2���U�P�s�UST��j�듔T�EY�(����V�QU�:U9.t�妲���3:jS8\�Es��H�Т�DÑrΑ��I*I֑'B,�(9յ24YEB�PFiT��FaTQ\�.�"�Y���#�U��E2	X�M2���N�Zs�Tit��Qd!TE�6sZZ�
�BUʹ�HDDgK!I��p�PG(�Dt��3;PC�3�D�IQUr��s$���U����,B�*�41
&E�r��
�G+�&e�
%E��9U�\"(�hT\�Ѥ��U�D'BT9�VaDi�BJ�.�Y��,�� �9r�%EQ�U�\�.DQ�r��TAQ"QI�"ۢ�K��@~�h�?v�#Y���#yV�<J����<U�]��h�������]vaܝF���(f9䩇�s������5����{��7�K!K�R:�2��\�� �(���dj�m�j���oƱ'��zz��3h��ήW���q�tyf�X����'�U�5b��N�8 /4$}��SB���s�Ջ8?\t�����>���r��􊧋߼��(��\MY��5`�U3�J`��A�BU�^��꘺���բt�]����Y{)��,�wV>D��!��sӱ/X�/c��f�m���P�d��`�B�u[[�)Zk&J����+R452��d�pj��zs�&�w.TH��9��W�Nik)��D��U�Z���y�.�ɇ����;�h�\���.�OPg�'	wr�u��V1R�`�2�G�eAl�v��@�p�V6�W�{zbU����#��i�f6�ʺ�zZ�й�)"R�Q,kd�+v�f�+��Ϝ�I�~���U�p�ӓSfZf��S�:)>S�-sO".m����ٳՙQv��M����ʤ2|�)��3���v�[���N�����=W�/#w�g�]�t�ս�����_iܔBސ~��E�Sη�إ�oR�F��8v;aܜtb�e�٫�n�S����ⷎPΤ�4�l^m�:����ѧ��ff����2/
�d�0=���}ް�t@<�{��U�^u<�Q��J�����l��9��>��yk�!O�ÝO��ü{�I������ӄK$b��M�6�M�z�L�5�b)�'��i	��{|���
��$�3_]������W��L�}�6*b"�k�B4j����S�Ltӯ�~S�od>Qx[@�^�ōq*[\�e�1,nTe2Q�Ƚ̭�&j��U���wý˻��bz��<l�EX�~Ю[56%�E�VP��\m�K�P������'���H�H�˙��nC�eR�|�j����*/H2�#R\��k-y�i#Y>YW�[�c0MP�a��Ź�髨Q�xA�R�G��0ע��5�z�5���vo�U��y��qW�<��x�MZ��uv��T{H�#���{u[��qV0�,�-���	[���,����9��Z[���@yBz���0��W��EC�o$�������-M�b���7�'���yʮ��l���w��(��a�wzT|E�s�y/��z��N�ͼ�	��؃�4�eʜ4��{�oTu������:��V�`D�MNё�3�U}�U<{�*QR�FWF2Sal٘j$�ch��B(�z��[�d����OqF��<�ح�O�Q9ɐ��h��ie��iX�Y]6D��ڞ��Ta^�R���a��f0Z0ay�ٹ��SL�ُ^�WK^�ֽ�f��ܝ�p��r�a�={|�}8����s��y�lF{B�`X����Xi)U��,ʳ��I>K)�9�|�;m��	��n�50��K麲�눓i��c�sI��+i`�!a��i�m�Z/"uM�3e���VӒƥV+M��9��n����������DSC%I偔%�í���}�J�\����w��wLO�VP����~��_�w�{ެ�����x22L�Q�a%�@�P�C.���7bbť�xmr���3X;�,����Ą�4�{��+<�:4�f*oF��A����q&p+l2aM�V9x�m!��$k�^65䈋��V%��v�:�$�L��^vs������ �o za��d�X5��ٲ�)z3����t����?{G��M�8���P�X��MsF+��W0cֹ�T�^"�ͺ�b}�n*rp,@��]��o?�}�SxR��0H�52�{vm~(��T�l
�_�e~��$������ܴ�u׉[F(A�ZZ�W�e�Fֳ-��x�MJT�Pz�p�6���ܵ� �VŜ�ߊ�'������e������<|�/kϘ���?b^�U7��/t�b����T\)hM�6[b�8��4�c�/��y��A�I�2Mn�ѹ��3�g�z�1:�F�4
ق�m��D��TjɈ��7��U����ea64�w:c�|�73ӎ��ؾ=�#��6��[��p��Y@�c�c�+p[�j:�eA���A�u��?	�PM�M7}|�E+�-x����Z��^���*�N��}�h䬫�Yfx/_/n�^�b�QɏTz���)�uL�r��X���z�,�C�j=���O:2֧�/$<��ry�^�*	�L�]߰I���$���*BXs_},ȼZ6�J7s2�Q���;4Z}����[�R�V�I^!�p���[)��1�+�&O%�^Xiٹ�����`���
�[�>�|�u'iIm���K�1��{���b��ǻ馎��l�A:lsܼs�}ՙ�z���|gt�Lz�U}_Q�пrPsga�y��n���ʖ�shn�s������W�{4�û�`yf��lz��6�e�~�j��C��,��쨰e�ON�H��͇��M�erƓh��OM�)��u�d��]�qf��$��g��k�c����u��Q�TAGHz�L2[T\�k�B�5P[@Zݪ��k����bQ������<w�:�V���3]�����@T����s�w!��]��b�6��|�	=ϯ�6��Ӟ~��)x����'ܘm������R�ڄ��U=��y���K���?l�>}��O�{�Rdi�A:j�i�\��������8��:�5uL�sX�Xi�  �^�x�-4�4�8�D�IB�c(վ�cr��@��,vB�j-�o2�R�V(y9{��(,Z�U���J��T]̱�2� �@���Zg}�R���vr��wJ���֫��`�5y�sUր)�R;���J-1 �Yj��_�Qw3X��ށ��\�r�1���}�t�����ک���P��XH6�Uec�&L�a%D[܀�Ciu��-ھ����⠬�|��v�*-�2_7�9��y��C��7T����Ɇ�H�h,���`�U`�)u+����s���6뫼'B�{#��1h�锆�z�;�]Y�,�JU�����ͅth���ݎx�W��?����!i��fr���^���,Ф�[vEj�|�o� �
�f����w����Yƅ��q�2��܋w�-V�e�W�Ns֥ak�<�E͇!��u��l9�+�ڿzm}�%�v)�u�-��,�GKNS=־��J��6�2����_�re�ue9������5i�&꫁���r��L��S#HH�u�o��Q��r���4�V��Rk4g͹2�(Қ�����Z����,�P��R.$���b�i����.�Ѫ2�e,���Mz�'-�?x'^�[����5Ѽ2��w�k�=���~6=�pn���6�6Tz���r٩�R�Q��M'�	��]z�#�.�]��I%֭t&�{���n�����C���t\'�M��F�[:�3�V�uz�,���Y�]��Cy�>���r�A��q)�J�%v�[�,s+m��De��$v�k���v� G��Fr�L]Vh>a�X�����2���-S����D�@$k��po6����Z�]@������p[�IG�u��x��|�f��L����̦}�i�e�[�U��gW��R�&�vz��x:ޣ�/�Qvkq�D�1*���%�f��d �Bt�ܮ�B���i9�^nu:��8�oX5,C`���X7�̒�����1]����%������O8	�`>^�cvmL5D��V�"�z����U�=��w[�Z��q�v�]����prր��H�7�H��,����	N�<ˌ��h+i��+�|���R�F/,�n`iU�30ׅnk�W�X-��s<C���k�^Q������o���Q9Ə=j�r�%P�a�,VF>�Z��M�m�ݺL�ǟRO�!E�0�Y.ڢ*e�@�T��������d��0�s%�V9�sI�%l�P����i��������S�̕3A5�4Y3%�Bܡ�"�T($d���"/�C�%��̊��)Y��q
�/��i���4�M@��(�]U˄�k���Ű��]/���[W[��B�F�k�Nd�i�@��UǪ�_�܊H�ͮ����8!��a�i�ݚs�m�f�sNSZ�)��RyfP��g�q��l\�2�@���{�d��M̚�Z�>܁�S��M��DR��W��Ӈ�V��� ��w,�L��s���/b�Fs��[�}^Z�^�`󷃙��+[���bc�e=E����F��H�e���T�{վ��U�ZN
�ջ���d�a8g�-7u*��`����U����J�/X��/AԫZ)mv�=Yȼ}�+ؗ��d��^��S�{^e���mQ��&u�����x�R�f_5BNg֘5xlXZXi�M��j�/kϘ���[�z]z��ӥ�ǧ�"y:��bɵ���?�P|�7'N=���ñQ�"���-�0^t��k*�s�)ek���(A�h��-�}am��Q$O�J*gQ�m���^�mC1�W��Jl��k;aW�s,`�`�u�}��H�>�m{��:�N��ް�ަ}s�y%��G�>���>f����He��	�x�.�57 	*c�Az4�n��I]��JXa��B���r?�����}|{�W��t��y�y ��b�VǕk'k7D�����mQV�K����Z+�m����oy�zI�����u�W����M����s�C`��V���7SLY͞�x5�A'�l{;�u�J�T%�l�Z���TkC�dQ'$���Z�sv��O3���T�-�.VY*�i'���d�Ե#��S�z�t(��c����⬫3��禸||��8�+�ĕ��H'�zܚ��}5W�ĭ��t؏<3��	�c��mv��M󏩚��X晜�tF�>��u5�kZ��tci�7���D��>+� ��<����g���67[պ�6���I��{��{��	��v����ͪ\��,�w��ɏ:�!]޸ת���oJ�;��ŵ�j�4<G����D���{6;��-�e�IC�&o|��Y�X�ߋLA�Qx�FJ5uKl�@l��i:'Tčǒ�I�n��jZ6��,��>�U��y�צ{^/}�o�Y7�~2�LD�H�פ"�*��l��j���W�uT����;\����VEC7�h�ǹ@v�R���5����L����m�7�A$9�����{�fX&qhp����{Xzj�.�Z,��旐;��R��3.�qb*��A�U5��R��[;Pg.���;uHA��V�	�	��܁B�Г���R�z0��T�R݋M��0s6v�d����\��\��� |�C�y�f�����Xqo���.�����iu��m?iWЯsY��U^�����W��b�P�a�o�X��تwj,X�-Z^�u52j��(���IYf/e�V
���\�<+�#7�-,�<<�Y�G�'_�53��/b�%��������T�,w��{yueN��1�y+T�}b��k���}���;�'	�{�>�������X)�����J�<>lꃈ��9�S%c+~��~�9�{�dY���2Z��𽆽��{��oە-�͔���#�ve���O�a�z�ϧ'�6ff��RTa�0{���e0�%���1�YL��ạ.�z�l9��	gKf�˴�uQM�v������V��z�^uI�yd�C��D��|6m_������5b#�~����e!�,'�X�����t��8���L;l��ݑ���i�o�z��|�>$���wq�����~[���$�o�v̾�'+��)đ��{�{fx�Լ_"��~�В�p\f�Y�x�1 �K]�Y�����_J4(�t�Q5��J��j������\���7�JTi���6	n��oq�����0�"(k��G�:�Ȧo(��I�]���s�5��
z�T�bb�w�}�U�oe֙�����1?�Sn����3�!&��D���q�{��%	�+���$�����k$�;U��؋����{��67��p��R�󰂻��=`B��h,���*�Y�
%�&� z�ػ�xfh�i�*�aH@���)Xw�3��ϯ\�w�����m�^�s¥HOL�5�&ݬ�}�`Z���(�W���n@t¹^c���#V�2�[�2��Rf�=�T�>���V�2�}�������[���>K��	����q�_2�;7�w��W3�Bar3��iT���Qk����₼�WM�XV��pG��U ��[ԷMh�������!��?[[;�q��1+��O�d���@^�����2��b�E.����U��%��ا��ŽG�4��Y�]��,���-8���&�p���Wwy#��t�Ow��6�G���|h}�@H�l��lX]��sˌ����/�n3��r�WF'�/;�8pg�[�{�-	}hG��ܘ���-P�u������m�fRLm�5��-Ӏ�oK�Vt��'8��*��z��J�4dh�ˮ�J��e��ĵ��Fʀ6����- ��
�FX����v_<��o=<������!��Bk;�'�$v,���īaݙ��նB�@�fV'�S&UoWP�e��6�m�5��豃$*�g����	����F����:z�/u�^?&�]eY�_��S/�����(٭k%f��*Fipyp&K�d<k#�w�Q��5�U�D�M��%������WOM��[4�V������2���ю�2F˒���j�c��ͱ̰�15�X��٨��2����)��Q�h�H�T�%D;��4�һw��F�w�\%do}�
����]����Q��f��YL�9f*Z�m�v%&�C��[��\��dZ���%{�wO���=�9�hc^/H��n� ���]�:�=��xa��8��8Z���@��2�>L܋�=�j�W���q��Y��I�u�L�#ܽО�9	��<���G��Ҏ��{�2��f�Ҳc����"�<n����чl6�ǰ��kOHW�g\3�5Wvw���-���=�����=|��!��{_��ԩ:s����k��J2��m���R����`PY�H�y-�k0�Mʑ�p�Q>Ʀ[����SӅ��H��W�o8G`�K���qG���K��������3�X8z�d�@o�ѻ(RX�]�󊼶ED=�*<���(r���2�B��	8YI�YQp����B�N�,���gT ��
"�E]G<��QA�S.VYq-&UW8�Q���$3V�W<�UbGL#��4P����9����XKT#"0����TbXr�㧷��eIʊ5�&����'J(J"-B����q��%.DD]:\�ʔNDJ%eh'.Rʊ�)�Uh�I�W�*��U^F� ���EDEÐ���ETBs�W��(�5J#���ʉS�]��"�����EQ��%�*����f$jUr!:I�"��*�̹UG�UQ�R+�G2J �R¹Q��TA�N��L��]�'t-D(��; ��]���2(�TkYTAV)hh~@4e+�w�{)�K�.a��T<�\B�t�Z��ٌ;�*��+d�\6�1�7[8�h���z8�53��Pحz���4��(�'S^�V=�2���MH��d��B�í�#6�ܫ����Q;���/��ͮ�>\};�#(��)�o���Z�����⧌��}�9>���P��W�����q��[Mz�7�����y�,�~�|^52��z��$@]���Ė���j� �}���~�Pt����o�b`y%��%3�lL^���w�'܀H�^˙\ͥ���������*��j�.�E��'S���cP��zD�^���b_��
f|-�u�9���pJ~C�^��g�@��$�0��Ne0����R�~SSϛ��o�]�j�q�#m�8�M�%	zL��u�8�\��;hsI��pC�����oSE1�EB�/݅��!���j��@�+f�ݭ��Q�:F���9�%V=�b,���w=M�\�D�zҔ�^Y<�i�O�[Gd��}�wyN�C�#v�"�8��9�� �f�L����+明r��AuXf�Z�x�߰[m����`����ut
���	B�=�;,�w6Q������<���5eS"+�q!�g�+ugW�9�e�#�����s��an�=A�-����}l��<����K���@3���y-�P_hA�&�V�&uR��.q������4*jlE�%dP�޾3t][h��Ի�Q��6�T��+�B�l�P]T���ՠ� �BL�7ոZ���]���=4����Zhrz�]�-�{qg���ୄ���*��xS�^�q·3ޝ����d�J;@��^��/K͟���� ;(iC��,s4�+�\�x�6�6�E-x�p�*���9ӯ�^���p�-l�}M
'�T���c��M!��[6ܶ�i89ܿ3
�����&���K^Ht�OF����|�d)��}�}l'�}�(�6�%�ͬ�r�����o@�He,_|rE^���[�ښ.�o��_y���J�gD�\����j\�%aAܞO|��3���DS)�u�+����טc>��3�au�:����Y�!�p���N;5i<�v�x�Sy�F
��9�@ൠl��ɜ|�L,`\8s���D���܉��y�9��F�k�ш-��~�������o����& ]g��e�:�,k���-�ŵ)��6Z���qc�u�w���d�ae0�x���m�'��m���|�������u�s����l��x��g��c$k�`�v�YN�(+�M �^�c��R������|7�"W˻HG�5z���M�����7�"�W�� �Yy�T.4p.I���R�:��/�!��ti���mK�[�wqC��/M���Hk�כ���^����7_N	�"H��Nd�{Q���S=1�Y�xS���o�ݫn���G�*�l]H���n��@K�%�3lI��iɒ*T;�d��)w���*L��L��j��i���x�Ϊ���j[P�}r�S)�B��*�!��!3�)�#��|�	���$
����V��oHsSϷ�7Z��Fr_\� *hR���KV4�Y��������6r��Yo�y��i?5�i��c���M�l:m���F�z%;�h�N)�,�}��twU�������Q�)�SJ����'F��ML���u����4;�W]�TGcMۮ�ٱ��������Έ����E3��i�)��vu���ģ�
�;�=J�+�$ptB�(�u_k�#�QÛ���0}G��f��T����UW�<W��y�c��ӎ��W�3Z����x��ni�#�[œ�~���t~�V��J�W��#�g���
\��.��UL�Z�X�]8�x�~mW\��D54��_�"���h��B�,��xd���߇��ˀZ�[�&�RW���S�67*}���A����3�G�(jq�s����Nq��嫸��s'P����5��p�R�3��h����p,�S�s���3D��޵ش�p{�*s�uܮ�@t5���	|L\e��<���{�S�Vfjc�@��c)�t��'�w�2,<�)��3��E1�������xƲ���q{�1�#�����L�i�极EG3���|��#����@�=s�ـ�~Ǒ�[YD:�]&2����`��m�����c���z]DW�Ep����������x{�-�:���q�Gv�z
x��99��z1�d'����NB�q�g��یK��_�:-�^�����7n�}�v4�l�.&sb7s��=��NM��H\��N�}�φ#Pz�O�*"�m�i��y�ů�����t��7m�@�b�@��_<��^t��xc>����;<��*mgq{��/�y�X�A�����jy�s��I糧 kڼ�G(�{�Opl4 �c��Ixqܴ%Ng\��6����g��HC�]+��MJ~�Q8E3wG`�:����Jҟ�	�v�O˕�(�_�.���#�L��E��?R���ISE3,����ʛ��t�ף$!]Ѐ�73�Ǔt�̛�Μ'.���昅�� ��r��LS�g)Dny���i��K�
�.���Z_����+�q(��s-
�ͳ�����z)ܚ���.Ɵ�{Z߮��@��_3������ө[B�1L�߭�-���&�{J'���SM���x�Su���`�qZ�K��QWx���=W�]Y���_��i*�]G� <������L>~~�>(�g'�Q,��q�w��kLAu�٪��SI�y��f%!�׸*I���:��wz�����$�V���~ ��rl3��7���Q���Ӻ'$��z�����MՁ!��3�)�u�ots���d�O�������t��j���;�y�:6[^�7q��5��Mk�Gz�{E01�_ ��ۼ�t�p�: 1֟p�sL��Ⳃ�Nt7d�T�F�Fv�]pP�̀�|rfK6j�XQ��ք���H��>�s��ǥ���Έg���T�#d��>�3ɷ�Fl�mqϓ�6���0��j_�)��w޴)��7�g�Q,��}�]7v1#�� wm�9�S:�-y�3����`���7���۝.��ɧ��o�.0�Ï��M���\���>SV�\Dg�E��ѻM�������V|_�z�'%��W=��Ev���r��Ay�3O���{�S�#_L�%�l��\Ff���3�������x�Ίh�M[�\�!�Mҧ8[.��'7��i�f�k�wf�h��G=�%晫g�U����L{(W������xq���o�����	���]-�H�L�t ��+T/{Y�V�l$O���J=�#϶�M�����4b���V�t�Q���`��ӳ�ul<��pk���4ji
֮Z�=� >�Bp�b��Ͱ�-o����Mf�ԾX�/y�F�Fժ:��t���{��w�x3��p,�jZ�)���91�3+��tN>4Sui�iDŝ��&��ND��r{"]f�L�����Ԣ��LS�nXCWwmA�\�L��pƝer��qQ�� g���񚟦L��@w�cC�JϜҔ�L�y8�ԟ���s�6��C��u�,Ěq���
 �(�L󱪛.D,��P���꽆i��А���I1�R�WQ����Q�Gr��X;�T����'�m`+P��G@.�j��X�.
�/3`��e�Uk���ۯ;Y���VA#pc ��0��*h��쨴>�Q��!���f$��_1m7+roKvڊy}=*�CPY=�Ҏ�/�Xf�Up�
 !���U�w2ڃ�D�!�t�ĄaÝ!���K�3��kג���_^����Swu63�����tRժ�B�o�0sgc���.��LC�E�h��F!ٰ=�D9�Ӡ+��|����S/K ��~�~�p��"�mM|�d���Q " �k�ه�FB�P��g\���06�s�������\��'.�գ��}X����HZ�S�����v���3�)��*r���0M��:WN���� �������g�x���w��bȋzF�=�u��	]d�w҇JC&]O��av���Yuʝ������M�>K�u��z4O�N�7��T"�W6J��N�_�/u�ϔ�>�7��)�[Df���Mle���#c^��r�$����X�幩���;��Ηx��|��#W�����pA�5�ɜ|��X��6z-�{{e;�N��O�D��.���SFpY�;���}��{��& ]g� ?>ƿ	B67)��]2B�����_�����l�w������Szs���N6�[��2�W��f	?Z>����ؚ�|ޒ+L盄�	z���������ju����g1
�4�[�1���q���r���䪜nT�����q�-����U4�D�*��O;���ڣxEzL��C���[;Ͷʽm�Ǿ�H_wms�omC�n�@)�LZ�*�-�DY霡��潊]ƥ���h}8'֝����M��%����\E�rͼ� +�\� *f�)�}�U5��Y�����5M�JE�+�n�VF]�Gz�=�٧�	}fX�8m��M�c����h�p���,��彣e8�b�;�&s�?E*ʢ���V�sLF�E�
~�2����Ttc#Svh���������r���S{��cۡz�����k�w�=А���*�R�Zr��n�1LB�"Oa�(���^ n�]G��<Gx�����;%)պ�Ը"�δ���v�
��.�r��R���=ݾ/���y��ێ��ji��jJ�+4��f�p��S�����8��\�Mim1�i�.�388�\wg(n�S��vu����d��
k�#�KFmlf)�;=��є�p��QO���z��+xw/���,��h�g�i�]�	l�ro�1����)k��s�^��`Χ~���JR�g���'����rB�Z��N1�
kǆS�= �M���]�!�x�)X�ZH��k�}q��m�[��SB�膦�2��sO�Z'��2���,��Ʋzg"�BiSKt�~cՓ0'�a $S%��l�ۼ�[���
���ߠD��bަgV����������7_����MKm�[�G@ң��h�K�{���j"��~0�`�G:�0�?s���[�����@��K3o��L즽�uYdW	��W�oX�=�d��Ù�f;%:�k6Q�;��<rx�O�'4T�����rvSх8�L��[q�~��0՝��On(�Y}|�o-�T^%��|�Y��e9N��)�|OL~ _���#PtpF��ry����Փ;��dnQ����u�6�T��~���L�����pT���V�[�-9���d�<��m��9wK�1�AeNb�v�m�m�D���1�܅�#�+�̼������k��v���l���&{<�1:�P��o�Y�Ǵ� ��/�?wJ`�)��i���@h�}���t8��Q��݅����.��k�~��-M�%��jy�q��9����u��L��7�2�|�g��St����ᢺ�����^؜���3���_J�Et��5)�qD�����R*en����3��8�"�7ouf��o��<��\��C��-/I)hK'��m�r��6Cu��nr�Nе��x�3Ҵ��&� �y>Aߍ�i{ip��pw�|�u�)Dj08b�d��s��
�ۍ���\��\��P�竢Y3��w�a��@֍��u^�8����f�vTF�cr�7cDq8gtG{�>T�Rx�wL�R���R�]k��^��i��,u�s��^���J����=��Gtt�f]�zbxN4)����dC��FZ&"��Fȱsu�Wc������nX��e��I��v���\�n���7��L� b����eH�4�,�2�v���lWy�	͛�NL�i�]A
9�:�	ki�t���:6\���L��x�C���>=}�_�o|JcD=�ĥ�����>Nt���1٘ym�/�w�O-�/�	���lY���(���)m���I��cU�l�3V&�/UJwP	��!�tK_��7˨�+����Vl���	YNqy��9��z�쓆f7GF��C�]%�]���!�s]��ۣX�`t������0������:n8�fY�n{�����>4	�u �C�ٗ/����S=�k�2�X;v��L'-����Ў����&���y�}}�k���1��[��sē���A��ݦ뜜���l�����+��񙑐iENr���؇2�.����睿gU��u�=�)��/�A�:�M73�p7������M�ε����?Nd�SC�S�-t�9;�O��f�k�wf�h�9�x/'7!��,����m�ᠿJ���9���m��頪\-�����u[��v��!P��Y4�Ҳy�M��+/�{��.{�J�ӑ$A��dK��L�kzZ0Ԣ��LS�n3XCb�#v�vLJՑ�ۓڛv�,q� �Q-hS7D�c�4�Y��Z�0��tK�)♖O!�Yv����Z�;>�u�Y�[#��4nN��#�7t �Q,��cU6_�B�S�P�����>�Qt�]M���[����r�@-��y�ۦ�?[h�SZ�w*+�0��F�aO��SH��~�	Ux����a:8��I�}��@��݊��zi��~;~�8�[`s�C?~���Q;�3��_�?���/dç����ӈů6�ӎw�Λ�m=Stdy�e7 S#�`�Xn�]�_op��Y�XRz�ʼKw�eU�ݳ���O	m{HE�f�޿��,b_$���qJgZ:a:<X���l+˶�D[�24xbUӯ��a��rq�(ؐTVh����lv����y�D�V7zk9��� -�=���~^֮�mе�ȯ�{�,�Q�"�dCw=X�o�</+&lhKCy'�i�xL��`�� \\�� ���3��w�w/���X�dR�sk41���Q��B�x�.�ni�d�I�x�2���r�E2��W� ����W��6�'cNm����J�ـ�p���z�#oչ���7����̡(CԷJ	BR�;D�r�GZ��o�-��\v+)c�2Iq�s�e�5a��F��d{�`���+#��^� �Wo_trv��������n�w4�������n�}�X�+{�=|��)D��5���]'�i,��&GЀΜ�w�.�5�n��K���i�,D��g�W��f�x� FvD�����zd�]e����y���j�yl�؍/E7��I]�wq�鎥�0k�[A%�œ��s.Y�|7��Ӛ��Ұ�,#�=<Ⱦ&̋��Ïܯ��_M���LB�l��Ȧ�|91�3�d��H�8:����o\�eK��C-�{[1���;=�/�X��+^Cv1$&
��y8�c%J�l����7��s4�*�UY��K<^#丼�U��w��umh%GN���"$���6��7V�m��y��N7��b�#��H�{��Hs��h,2�|kj|>7|ؽ�wm�4�ea�Пy�q���kB���{�^I�����i��;(���S�125�of4�<����Nt]G�Գ@���/��EE=����wC�3*���k�H�R}�ǖ����\��s2�q�ȷ��tq���Ɍz	�s�����⍰�d�Ւ�.im&В܉o�Ꟶ� ���^]|{\L}7��瓪�"ݚX��K�)��gz9&����s/4�W�4�,�{��3���C�!�>���~��:�y�ejsEQ#N�3̢���s�̶��徻��vͫG�R�:��pN�s��4k�-<\�x�,��y`�����m�k�����T�~�>3 �Y2ھ���D�˓H٠t�W)p��{N�8�m�8���;�I����u���z�x�dU=^�H��2nhsr�5�|�t���˒��!�J�#,S�oM��z�&��4;ŒwA�]����wh���ٺx�j�UD�G�+~z��~�&�{�6��',խ������Or5�u�xP%oϛٽ�<w���w���b�i�;�7M��ܧ&	���`X�4Y庽�a�cY��ѝ��'��_f 5�������I"�Ć˔\�:w,H"*����L4���s�"4���L�L/D�"�U����$�"egwXU:%��������><:�(�Np�r%4��%���k#�HW4�XG8W�r3�r�8A&Ȣ�H�BCe<D��YG��E�y��]ݕY T�W��*"5
��B���G(��G��q(�8�Uw'v-�dil����D�r���
��Ku�����k�¾&���i����ԗ\���������(͉Ȉ�CD�Ax�!DW���𒊧�.���E�����k��G���9�sg:��S��V��8�wG(�h'hEۋ�Dz�u�՜��RIh�u0��*)<���HNZ���%zY� B�(�N1x�Q�]�����Ԥ �r�k�U�eCi:v��cشx9�d&2N�u.�\�9���طk����+��;ח���NT�1��S��;�����䣴��U\%g�4;��r埮^��r�v]�1�mӹ�8�	��@�^Hu-�:���{h �W��M��}MJ����J[J����O4~�_6G�u���Ϲ��.��Tb^͐��:!��`��{L�����u�6O{�]�sj܎jw������1rd��)h��h5���W��}r�����F�
�v26���f� �����a߫☹���w�^E��-������M!`���e� �:�	���Y���bO�͕�9�їu�t���L=���U�r<�����i3��l$ݑ�U�_4z��;6�_{	g곜^8�k�a���u[3�'�7�}7���Y1�� ��u�����b��6������1�9����5��'!\��'�x_�s��o�^�wAn��-�a�Xb��0�g��H�ɸ����d�x���;ک���΋c�o��V�Y�3{�㵱<+�Db��z�Ҷ��\`xC]������.9T����� 9�
��~(�]]��0�ږ����[�=9��1mI�P[K�A�}�\�&�[mO^�ð ��w���#M���ݸ!�������1��{PZ�\Ouduݛo :a�Q.U���^��=Q�"��>`��{��T�y�Q����\�i�k�Q�4ӲK��'+頶"_lgܶ��v��9� @��B��U6\��!�9B���"�5�L3�E���.&�t��~�����S��+�Μ����S���S�4)N��Ѫ��b,�U�M{��Wͦ_'72��p�|�C�B��4���HCיb��˕7m��:��1�h�p��S��<��l5����α�'tޅ�9�nC@(��)4�jy��GB X�݆�2����u�����ew1~�{)�lE��f�:���bK�:��~	�pP�k�~B�'g^�.�|���
k��:��(���/q�u��H�h���νa�(�X��iS�?l�x������Z�@�����H��@^d[�4u��T)���E�[�D�3-��@p{�xx�Z���_GݰK�v�Kb�׹%�����hM�ϻ���B�膨3!��r�a�=�c(GA��nmŦ�6w����[��xl�vL�����t��_��w�2,?(���jGm%�#�4�[[u�vd�ѯ�:��X�&��ߛF�M�?�������e7���
ݵ����E1���|*JV�6]���=Ք��`<dT�Ӫ�}m+qޒ��|��F�S*��6v�ΐ�&������<����s��³�H;6���[�~���%��'I�}���*��TSB ���H�w{�wBޕG��e�X�D���F����ƛÔz��pcԨ�{�8�~�YW�1�{�����OL��M�Xka+F�V�'��'�<�;���<�������z�'�^x�o�e��̞x�7��2N&��SQ�ž����y^%��~t,��]���m�Ͼ'�cN�}��1�����EEGn��l��F=����1����~*t}�����)�KS>��f	�|��\E����S�{�şg!ߏF���fy��5<���I�v�l�ג7�S8�M�e>,j�k�g��n�n{dƬ���n��V	@�)g�Z���WJ�m�R��NM����R#�����:�3x�9j\��D��m1r^�f	�P�&��MO6���Y=~\��_��n9-a>�����SQ�j�o6�T �(��,�#PǶi�X*b���r�/��hČ�0��e�%]Y�ֆ���F�GCĎ��4�^�p��R�D�g��4���i�.�]Ts�1�bn^��T���S\�}�C���0�^��O��Y�C��sD����g.�V&ú�n�W�2�t�1ujPܣ����a���V�/��9���:uf��P����}��ɥ�6�5Ҿ�m�6$U���{7.��"-��x]h�c����,K��M�`nf��!j�����d�}��`�����ԺWN��B *:Z6�V�9���;��E��1�����`�-GN8��A���5�i�L����H���:K�\q���_}WlL��.n�7Nl43�1׏�ٓ�)��B�xM��Ep�ƅ3����l3��O��n�OwKX�'#��P����+_��NlG" 5�j�XQ����%����,;�}]�MUs_" �FZ;w������Y)����|��.׆:ϝ��jI��?L"������sx�}�V��V9'�g�먁,z�����6.�4������[&�={z'Ck#rFp���3΄v�ә��!�[��5WȈ�r�q8n�t\]�� �M�p�G[�t���S������zߛ"77r�}�}�<�V�^�ǻ�90e��"Tl��4��Y���\�Kձ˝��ܰ
�	��vY������9�K6�>K2�����ڍ���n�N:��D�7���Ǟ���T91X�z��	ޝA�+�e5<����o�Mڶ����2hdC�Uq��r��@[̢q�\A�ӑ$SJ�@�6D��L�kzZ1�J*/�b������p*�V��S^g�:Vq��6�uF��-�!
�/��V6�7�au�[{��gb�M�b�q��vq��]<s(#�ϟ2ʮ�Y[����%j[�L_=8�]e`{,��.q�.b%��IЮ�wCQv�hˊ��҅J�2��V>'�B�OzTp�u� *eև�Ɉ�)�C�U�\׳��}iJx�2�ʪ�{����+���DtvI~�!
f� U�ɞ[cU6_�B�L��P��.�kƾ$gY����ʮ:[y=X�jg��n���O��|��^��J2�b�UӗP�b��$�e-�T'�iSO9���]���:%�"�p����+�w*{����L[.�df�`��U��ΖGX�]^�[��,��l�Gh�,3z��K�)���� �l)���a���np��,��(Z���(�zU�#Ϋ>z5���\�wu63�N����b �@Pt������z���}�jx������@p��4R��.UE�?O٬���C{�)��Mp��V��Z���k�S�}lO���K�'�7I7�Q��,^��t�Kg\�Tnܝ�W�Dۋ&�7��@��\M1��}�C�{��3ϹM�E2���1m���g0W�,"m�o8�ٿW]�8����dw����tE�kޗ~����3{�_)���U�3�!�����k�Է���\&TI`�W|9$��=���L�(С�׽�o{bk�𖧭Ir�o�� Q3\�k���H�gXh�d�M	��$G������p�����M<�)�0�w�$7]Ǝ�ù�9v)�y�$�����AD�K��h�`�����"$b���j=˅�v�Un~���&��3h���׼Ө[-�����}��ɈL�P���5�;�O����~ O߃�sB\�c����_��Y�0��Q=[����ӌ��o����-�1���3sjI}�I�������ܡ'��xe?/����W砍�|�ms~ϣ��c�nÞlj���]�]N��wE����!P�&���T�S�$SJ�~5���gإ�nM�"*vu�+��,Q�ҥpV�i��7-����O\�
!��Ê�d&r�5�t>C�3��:�zꖫ�/�{.�}	���p�0�j�NQzm�9[7\� *�)�tj���B�K^�emG�k�[?A�h����P��SgM<��HC�2�1�m�*n�a�hu���Z0#�����v^F�#c��{�IqL�;!�b	��T�jy��GF3#vh��<a5�Z�`\����5�i6G~�� ;��O�t�@tmw�@{�l��kI�נ�u�(��OA�U�n�=������aC�r�4j�Z�g�V%ܼ���,.��qζ�]�	l�q�2��ܚ ��.�1t��+�_qӉ���\������b��������G�A�vf�~��P�̇T���ʉմ��$����SƃpWp���'7��xg�5���͡M]����c"�l�:�ulUȫ�h���&�Ym�S�K�u�n�>��i�v�dޘy�Aw�c_ �r��z�u��g�E�> F��0��Z"��:��\�N��mD�M���t˫'�O���	�[�>Bmߺ��d)��j�2��DS����W���d�]L�m�SY�>��bxe'&`O�ap)��w޴&���dXy�6����t#����b�`�],''����0cƨ��l��[&��oL�i�M=��x��y�20;�s���E
��}�v;Q�];�����lA��3�o�9�}�4��;)����E2Ȯ��r~�ƈ����'�+�X�J��{& gTC��p���m99��F8�l���읔�aN8�v��-�{数�O��7��^�(r�*�X�ޗ*{��Y�ʄ;U˶S�N����k��b��5�1����}���Ad���|�|�~e�<A��o�ݷYl��5��:s�?Js��\������c�y7z���t���.����r�������Ni��/}y!l�q�m��*U�:����_`���*��C�J��zVy�UjWzb�W�Oۊ'���h��'���U����5.͒�����u+�p{h"�'\�s�#Ӥc�;���y���xjW��T��e�w�Y���K!�);ǻYٻҟ`s;���7����^!G��1��U�}��$�TzβKe����+��wR�G���_w-�ʊ|\����a�J�.ܙ��3�o(�uM�'�=�\�����C�Y���i*h���ѫ��bȬmT����Pj-���ͳ����4QP�L�S��h�C�!`��֩�(A���(���k�a�sȹ-�eD����kR�0����!V��ʮ�d�-�Ɲ�d,u�ds��B������M7b�o��:]���}���+�L>T�Rx����sD���/p�A�*mkcQf��d�U�e�hw����J��@,E�����>�T�	�S '�U#�_�!ܖkV����=������:"��Ey�׏��2{E� �W �p�w���G@�[]ǩ��t��ڦ��6v8��W�˂�,��v���${�$k[5ug�OM���ST>�v���ڐ7�[Ծ,��n[�g����]��(��ĪY��v�1�|�|%Wkh:��1�]�[�0��r�Ww���wV^Z(s.|�ynWQO\����q��)�,��)��jS����r�O+/{ۚ[V Q���Oӱm��^nO���."1�E�����m99��,��΁+dU�c5M4��VQ�3.=F��y���m�z���M����F�zt�J<E)���2������-(��&��qi��BՑO�j�Q�^=������Wlp����xr��Rಭm����T�f9uάMl�8G������ױv4�/@NF��Ip�G�_�O�epW��w���:�������Xr�|���Co��YX���{W�s�K���;��M�����*b#Pw�=9���g���{Փ�5�j4hنt��5-ݱ9��tݬ��d�����;�1��-m0�m��頪\Ls�wM>:�.�;M��/��*q��.vz,e �"��ŏ�'�S�=11�J�J_��J�Ԣ�V�/��DO5g6�asK^���j]�PGP@TKZ�ՏsdW�T;�����ޒ7uծ��{��W�lv<sb�ÎuR~B�:�k�7�Ѐ
�D�g���M���T�s�-E=�oZΨj���+Wu��qsٳO-}	�R����<�m�t���"�V��ʃ�N��5S~�b�l�6�(̽��ޱDt�#P�5T'U&i�B�p``��0����A_�E��Mi��W��}=q���@��b�4���9,��������[�b���в{��U�S����9��;�y��=�w:���޾hwJ��%�ˎ�>�S��9y��N���A`���bfz�7cЕ��R��lAn6ؼ�>ƽ�,����z�1�l��y3�0�_T�+mR����j�>�iA��L�U]�?%)땶k#1��_f��<�͸q��D���ҽlXy<W4.�1��� ^�0L��(���n�1����U���듪.��?�j�}�3X��~7�]���0��Z&���l�G��Ϛ	�y������M�/��ɼ\�3�'|7���-�}l)�Ut
h1 q Dk�[0��u�,�8Zg+T��8G4D������ؘ̭Jq5⫝�rqY���ܦ�"�LS��4DK�X���5�vw��`�M�Vf�7V#�Gax㮛���׿0>FU{>`-�}��1����y�+��*���^O�O���n���r���i���i��0W�$%�jYV��M{�:�؎y��Ϫ_~�+�;�.M�j>�O�.K͸��y�(莈��@<6uմ�`׎�6Bw��d�+���on1<4��;z,S��\����Y�C����yV��읁���<n�s7��G�{%;ǭN�y�oj�qB��3�<��S9m�Km�Փ;�Tw��tLaQo�ڶ��W���!KNNL�M*��d�B��0Z��]-�k�~k�:"�zI
�L���崟��a�n�@
C:�e�*�����WO;���s�ǝ��Y� �sa�{A!T��ep9Ӕ^���}r� ���w���H1N� �b�m䯰��o���ݠ�{ՑÎ��ӝ�O�b���Z�h3���W)�E��s�}ݳȅ��i�qZc�*ւ�O�u�ޘ7w�_.���U��쫉Y_z�`^F�?
������d��M���M�+<�T�)d�k�t����>�H(4��5/����]M3gYᢳ �O�L�������L��c��x:ʊ�h�����͉���jnfq�%a�j�u��!��ip{��6��AWX(�ᡢiE�M�Z&,�W�0�qa����*>����K����\gc�:�պ���f�W\�81����,��@O�W{�; ���k�ii�h�\����:y�vv��o�;E3F<��A@6U�Ֆ�>Ǘ�����&һ�X�[ڠ�'bǣ}'��k)ZP���WhMaE�($sgf��h�$�|���:M��p[qs�B��d�C��,�*�>Ì��V+NVCx���#:�=J����i����!�Q'%hbQ��z �����_Ow�cxz��wl��>7*Vީ��({��"R��y2:X�n�l��]V����0f!������U�s����di�\sٽ�c�"q[�U\��p�h�,��b�.E�mH�U�$�<�M:cs�|_��������fg�RKYW-�t6��4z��Z]��N�T]��畺|or�뗈���yJvS%L#�'$-��vs5�-F�0�*D�}�JҠ�:fn�ڜ]m��k}qs���`k�C�IG,���\n�u�7e#o)^nv�a.��(`�r=e<4(=7u)�K�e�k��[�{���f�A�J ��wUfu<�WU�����/�ޏ�}(d���M"p=���;���1 ܨ1Ҷ�۵.����f0K㏆�d���4+�J��6����C��\r��x�c\����f��J�D�Єy��'7����,����e�ֽ��ܷ��$=�w݄��7q��+rƪ:ىY�1*=X��uΖ�?�ic��w�8�7װ>�-��uv���V�A)�;L�Z�{�צ�Q���:����{g1�Q�Ge%j�{��:�2�*s]�)�c�*�s}z�:���a�f��8��9Y��YY`�u�������^y�d�������$!(�i��bxw�UW��	<��Y3�L�]+��^��z<Ǒ���廊֕{�8|�����,@�c�2�u����a�5}�6��W=�(��7&��|�jr\����b�z^����0�4s��G��J���������Y���XW�!�{�=g_ ���:����Wh�݋7��+���ԑ�ֻ�����{�{�Bs���jf:����9�q��I^�m��t.����z�L*��x�ג]"�Ǵ���E�kDLN\�t����7�z���Ŏ��z������X�\�ܝ��;�|��g��Wώ��3:�B5�I�ȎY�B��*� ��ȝ�U2�$�G&�˕E�wN��xy^�tr�	�fwVf��u
���i�EAˑ�*�=XQq�*�D�]VRa�N��z9T�rD�����\�/K3n�*p�Ե'tp���NN^V�-̫w/i�hU#�拒����z�	ʰ��$�s����Y��#�.Ufr�UܲR��
��DVy����R,���)6QE�GChs̝�㇎t<�	0�κ$Q�˔AC��.nu!��E���u2�%,��Ь����/GvI��
j�NM
���8N������*�%0�����/M�Rp��4"	�B�ob ���۲��`�k��7%\��^wonZ}`�����4)�;�s3�ơ��Ad�:6�ty�qh���s��8����?԰
P�4ʞBڄ��^�HC��c�ߗ*n�6�^��d^h����г���T�K7	���9�Iw�h����& ��yr�M5>w)8
00u{��F>(|�Jv`���Uon��>��DGO�~�}ep=�6��=㲭A�����C��5�3���Ck�q�f�Pwi��fOJS�?W�(}�VXkѵ�0�ηn]��$ҭs�n.���Zm[���y�5�
�.��z�����)���E�> F��0��Dds?r5ȴS�V�2A���>!Z�fI�-��\+u6�㭙	�y��
k��d#�Ngyn�D%�Et�We��e�,#�:#mFP��[�t�ɘ͛��It��Zn��E���6���Cj�������}7�4�B���6ž4�y�d,�R�V��4�����������o$�]k<�����F�/� }U�m"��mu��j�pcԨ�l���������{��"m�P\
y����V�:'yi�K�%���E���]?|^鯯�ǚc��s��k�^��������4�(g�[\�I�!ד�VdYM@�*����\Cs��W���r~Lf(�P��z�L��N_Uӫ!�P�}�F� ���Q�&�Q��j�8-c�Oz&@�h��ප�k+���|;=(-�Bhp���N/*�/�[l7�9mt�Fi���|�s.��-��~��l���Qy���ܖ�73��. �9ٞ�J�[(C�4Y��<�]߽9��Lb4���O�-u�OE>��eN����Ә8B��ɋ<�;�+nzz��~�9�&~C�ͨw;Ѽ���r���������հ�^H@�����{η���'P�gs:\�p�O�昋0��a��<p:إ�=jWzb�W����D��z���%�!e��J�mF��ԇL�&�k�B�&.Kצc��p�ﳩ���T�^Y=��r0�����kh���}��Ǵd��ЀJ%;�h�C�b ��j���c��'��v����=�N�7m�h��!��/)�WSv�@CZ�;9T�ɞ[c�;��� .�E.��wܥv7Մ���L��1����L>GL��n��V��ʊk�r'�l���=��6�3�ٳI��Ds8O�U�c�4��`"�t����M�5�B�?)��(]�t5���|�܍��w=�9-�*)���׏��'�W���������|!�n�>�t�,Dv<�v���P��:�-���N~Ү��kP��ſK�:ļ��%p���zA��U�=ѽ�
J�Z%!'�� 7�K-�A��Q�4��r=:�ޗO�����|��{�h��������N�<@Q��A�m���'�j]y6��\��`�q�>H��\)����RpU�.�:�93�5u/�G3�c]v�l7�ʩ�.�����%� :�[�'�#ݤ�4C�v"�?��|�}�����4V�\�)׻�q�{D���}7��b��K<�+��>=s����+���������?[~��-cWf��X�潉�V���%�r5��%��>SW���r�q+�v��rs�����QN�Aumus�Z��C��9;)�
�{�z]�������u[�uM�g�N@�~n�J�e�a	�^�o���O=�ɔ*F�+g���eN1y��Op�.��%��\5_��%��S���~!qXl7[�n�F� �@z�@�y�����P�b�w�[L7�Pg�AT�Z��|�Ǔ��q��\[L���/����Rڎ�0o����"P��iȒ!@�%��b�w�k[��Tq���̇���q�75ɛ�Y�J6��s7���������D���:le4���~@w�þSU}�/�ѹ+w��=����6f�x�Y)=2��^��/��2B� Q,��j���<�7:c?Jͯ(w�q��L�7��3#ec�q�����HohGԙ�y��vq��sԪ-�D+�`K�L=4(W��ݿ=�W�R��Tg,������3�f�u�魴��iAcE����tΤ;�J��>8iM�(��|͹y�:Z.����hw�!?W�M<�BC-�J�g���7I��DX
�i�;��|�w�j��ͱ>�_<����>��H�9���L����(��݊a�Zzil��ÕVoTq��D��[�l�n|��ζY�ZP�N
ث��&�C:���Gh}��s�3c$��{(-]<���|��q#�z�� 7���y�Z�x������__X�K��ߪ9�M��=�,b4�9H�+2Z��}JR���K�#�u�`pt~���{D�TbY�>�}г���bj ��V�jm���$�9������]L2W@��'�6�z!����J��r�8�����db��(NT[�lL��u��w���D��{�|�7��1O`���;ں'�z#+.��̿f��t�lD�v�E��R��t;�kwT�q�bq���|��{As?ݵ��KI�= ���g*c��p���U����y�P[�:~����9�o��N��0�7����էz���v�F^�N�b���:%?���z�i���Xg�����y0��oxQ���܂�F����Q�h|�-7��0����.zLHJo�h�i0�Y��A]֋70�<SkP�5�����B9�⠵8������S�� �[oW6�i��S�!��Vl�x���:���uJ*����;@���J\t���1o�P����t��n���`�����V����ʷ�wd��a��s�$�/^���s��)�=juÅ����-�;�ܸ}gt��&}�����o��1��ov��"�� ��5��n�T�M�ɒ*T;�۳�HF�6ם��u��.ﳐ�ǣH�1�"�i��-�����s� ��D/tJ�ƫ��P���fVR�Y#��>��;��k�ŨHE<���\7NQzm�9[u�p�³9v��sү5Q9<]��a�˘�0�2d�+�6�!L�Lp�eʛ��)�7������(w�Y���m�q��R��הJw�Ѳ�W�b�j���~j�SI����Ttc#oH�M���7q��%��!YVj4N�Ά<�.Bi�ܪ���δ;ظ<!��%,7��:d��[�y���������d�Eqz�Rt
��S=J�+�$p�P���Y`puG����iT>ո	�u�Gj��1l���9���~c
w�����)�wN;�������(A�4q�p����0a���Ƨ)u������*��2:{ON�V��m��'�w��q)yϒ��r�U�(�-�p�{6.=AL1�&���W��x,���F���H,�1�Ij	��7Z��n�k�YT�W�E�ks=7�o'��5g`��,�xqq�wgN��Sq��gt�J�C�������\�v�wx��홨7���\��~;`�:jp],`����=�LFj��mc�K6s�)�ɘ����C�qBm�xȰ�s���w����õ�/�>��G�_Fx�h�6[�������/�8�����4�o��
f*9�6R{Ǟ!UsAkR��Pw'��2R0;�TDc�0�m��޶pc��7c�%�f�=lvS,8��aD�$�ۧw���:���s��4��yV��& Om�x5����'4B����4!���)?a�訃Kt��[�F�8��%�v3�>wU�RnS���,�%A�NS���8�t{Uz*ϻq�R�����*���{��^1���e>p�e�<A��ڮ��/�� �~��m�c�+��W��W����ONL�L�9"��&s8��z7�љNP�5<����Nkݽ[ �S���x�pۜyUn��g8!��3���xҾU)�r����O��AU���+�p�������XcW�����00�u��{T,E��!�B)�h�C�.K�L����6u5<����;���tK�\�ڳL�x�g"��m�M��~ђ�ŔJw��cߚb
f��筪`�q�&��7�<wa14���e��hpV�_�}rS�̟,�5�I����nt��gx+�9M��sK1Rv,�B�VPX�Ou�3��u+"Vqή5��v1���v���ue���.��^,�2٢}}�o���.ct5�О�:��4�ޣjN�꿼%�n���~�����e��r�P��StK&y��N�ᐰD�=`gx��dG]�ba���UA~��8��T���%!�b�{���L��#��wr���9��ܯc���|�6�Df��9��^��q��+�Q��=;����[(��˺��7T�	�S 'A�߸�L6�eq�d���	1� t=Γ���T�?}�^^uY��3�������+nn�.5�,`V5e���e��!��fr4)��ߐ�r����w���tr"_�WPB��q����mWiv?&uz����Xw�Q�2�u�%1�Q��g��d>���c�úO>�y�[f�շ���}̉�ي=�~2���t޸���h}�JcGֵ���v�nΥV��bm�_Q�<�N_�v'�O�{�=�����Ll��2T������V
�>[���p���;���c뙳���,t�@`�`�26�����xv�s�Ϋ}��{�S�#a��ca] �V�����:��$"
l	�/�YS8��z{��}ӽV�-�����W��k�^݁G2�fI�/2��շY�-".������߇��.V��T!d�{�h�ƥ�]�6�J�h��Ή�t�߁�~�d��Q���GF����S�i���F�JТQ��a�n�����7ֵ�VL2��J��\b�+��v��|a��R�O�G���ش�sd[�|j���������ֶ�N����U.99|UB�t�5����S���7u[��jڂ-�� ��N>s�B^,A���"_�b�wQ������K���ʤ�E�����
����ڂ/���Q-hW�'��1D �Tm�鶛�Q�A���s7���i޷/�{4�|�<S,�C�7U'�T�{�����u��j�J�g�n:���ǖ�+��c�GLF�p����1/�}	��(�y�y���t���E��֥�ʋ�3��I&F��3�v:1����aL���kUAuRf�4.F�v*���-�٣ԿNȫ�ܭ8�^(s&Aq�5���:��J�{T}��M�R���d�����ߑ�vJ�i����Z*��2�vX:�Wu =��@j���,�>���qN����Oc���u�9�u+�;z��C�2,�˥��ut�(Q=��̇Fۄ����a�.���q�¡���C�SD�[�h�x~�S:T�
�G;�'��|f
��T�8���נ���>>U�M�_׸�u���+߷�a*����2�`����O}�;+u�@}�����R�8s��e%�@~\�8�����z;0c{[��s4����l�1����'&/�f��v/b縖���9L�������#o�u��u�,S͍��0����Հ�\����>��,�jy��\(L��d��󿒟���G���cަ.��c��9=����`��X	�MK*ޙ�z�ߠ�.��R�^�#xZ����)O�b׮�wݧ�}���z:�L���X�\MK*���׼ӨZٞy4��t)�E�K<Ö̫�fN}]ϟ1S|-��1�� �l���fzi��2��5��'�)���a�4��7s��d�l�Xr���JsU[��m�[�\d���g��H�����87	߲��(�vn��D߅�nf��>�Gٞ�B|߳�g�߉�=�]�n�+�ok����2 ��YY���+s�f�l�6s�W	����z7�T�D+S4��q���zf��s� ��3l#�k;:	�<Lm�9�|��"/�4�g�+��qC�Z��W��u�ۤ��q�r��(�	Oյ6)E��G'�]��`	�۾�ڂ~4��.�?L��-������}j�G,�Sv�k)��T=�bh�M��O�cuŸ�G`8HAw�Ѳ�S�Y Ѿ�NTi{�w*:/�ᛏO5<�D������"~�4�1˙�7��'��8잀�r�9�f�T���S+ϸ��V���V�y/C���-D����{^��U���p�D�H���=�	D6����=k��S
T�%�����@n��
�4��`����ݮ��}��9I���UÜ�&Z/��Upn�h�*�C�T�]�և{�W��Cj⟐Ί��{�m]B6�S]u?x%:�}��_u0�M=J�+�$p���ʚĻ����,��h��1ѽ4j�D*�-����.�	�-�ro���ywN;�uu�T)����P���@=�(��(�fa��N��P������)̞�-��\+gSo�9<S�w]s��)��k�L��ޚ"�y*����û5j�|���C��t�{�P�V39ᔳ��>ͅ�H�K��zЛ�r����W��X���2�ޭ�/�#��v1���E1���pວ�)���W��5���;i<���W5"����XV?x\�Ծ.�a�8����t�޶pcԨ�~m�|ȉt�0:�:�5��\�VwsSm�nn�.b)dW	�n�i�ʮi�L@�ې�k�'t7\��C]�Sv�u� rvx�sc~�/ީ��eq�{L��1/ӱm���WMY�S�����Ĩ;M7�_*
�eױŌP�Q��~�9�w ��<��ֶy��jb�]s��O��� iQ�`���a�%����S�h�z$U�M�������{����A��r{�a0�kQ�K�,~�렊�G���h�-�#���q� �+��a����'S�m�ٝbJb�^�,� �?m�Mi�9�g�?)T�1}�c�p�iE(q�8=�^QyM;�ޖr5���G��eA��-z�/+қ.�-2Y&�Ʈ�����fV�5ws�R[��5��.$\.�Ug�_yx ^7xU�.��G�:��Cr�w�9�w�^��W-=�Ӄ���)Q��[�Z�Ax��9���{b�!�q�� ̛���v�%��_Y$0F֚��N�Cݩ�,���8)���$��u��R��u8aVA�i��oS�ho��ή�nG��1����]bcY/)�_9�^�멋�@c�a4z�7z�p�y�dG��_|xV��	Wg{z���ˇ����H�N��p�����@��ü2���ޖS�3���9���L��yJ��;�����DU�-'��Ρ{��=و�I�@U�oI���t�ۑ��o;;cz��"�	�'u�i�X���l�6;��'�i0�>� |���h��l�XO`������M����&�ǭW35���ڞ��5t���\�N�D���.j��V|íڻ:��U�Jn�b�.��/1�[�����OG;np�
�թR5;W!;S0Βԛ�+�ƅY��3!Y\���z,7wu:UmD�iy+g+��Mv�tr�� R�B�ؗ��-\jK�Dh�y�G�	���\k�u����Z5#�7��bL�'1�q���38��L�f�}��{r�s��|�
ZDǄ����˸R�㵢��=�%G����WLu1^��x��_";/�;:v��jpD����k���k-�*�I�cr�: ��V�� z����k�eb�4�3��k��UF���QA
�Hbc�l{�F����샔�`ơ� l��}v���P��q ���:��Q+���lvq�W����"�*�o�~^WVx� !��{��>���PiF*�����繫�Q����gX,N�mF�C�Ұ�9���wX��1�_�$��"�����c��,�Y뇟L��H�K:����a|$�Z������E��d�!އ�U���;��vM�7�;v��H�\s=[��h�%�W%�+G�bw�M�s�qA����Z��˝���Y���!�/�
o��g� �!�}�Oi�r����.i�����O��[|�����e]�h��5�;x�c���u�)���-��̉Y]����S���]HQ��ۅ��y����e��aP�ݚ^�3;]�rvs�\1�E#�O]�<xsA��c�;��i���oaC)ΰT�A{�0>�xo0��^X
Wu�|��E����YV���X2*�؇o�nNK����Ρ})m�S�6Wf`�YqP{��9��1e���]ŨED}��`�S;���� a�]��f�]W���ɖ@���""P��'t��T��l�'2E9��%�Z��E&b$�]�a�V�Eʠ�	�0�\Pįu��E1�J��ԔZ�(�[���$Ȋ��҈Ԩ�(�*��(�-Yr9%�	��z�$����EEE7V��r��h��U�R*(��W2����b�r#L"PYV���(�4YEE7P9��*��XE껻#��]B'PԨ5u"s*9Q�)�� ��Q�˹4*���'�;�����RwH��t�̮�U!UA.�	�E���RLŧ)�*�&E9��@���H�Us�=w.uEJ�*�+ç97CI��G�d�fAvy���DRK5�fDW*���������U���QfDE�G+2�a� 3w������Dv̙56�GwgӶo[��3��ԙ{�,ݠ=A��k�ڶ�/9��E��g4�r{�4¹��lQsɜ�k�xW��ƴ��b�F���������o1	��MO>�{�����y��k�=*�6*%��@����r���n)��b,�SJ�F1���,�jWz�]+���1�o+�~�1l.Zc��׺���#�tvB�ԇ
�M�M)�ත�H��[
��ז���9�H��^�&��h�R�Fߗ*n���6���p@,�%;Έ�1�!`�����4h!��v���Y�.�x�C�:r)��F�j����/)�WSu�h�Z�Q�L��i��@�6�P�����C��v�����K���H�=)��5Gh��=���S�=T�+�dtU�wr�U6�f[U��z��ܛ63U?9�䳵��g�Z.F:�����!�n5�u���0���j��ٺUi�e���gX��1�ȇr�a��-l4S��x��2;F��!aE�	cxTݩ���ax��Q,�K�1ټ��2���\˂g�a��㵚���m~^�O4�!ӭU�E��=�p����a������#�%1�{TT���l�	�]t�uѺ`�5�׼q��Lw�u"R��[���a�X��7f���W��5��g$3��j�X���:�7[� ���ҹ�N��-�>5�p��ۃl�Fy��z��t#k@,�Ӡk���@k%y5 V�˫��U�Otϱ.��:���s����fU�u1^*9�z�
i�\_%�y]$]W}m��Ə������n� |eØ۳�[����|yl����Q8*��ЊY4�;�9=�J�q���nQn ���푵ݮ���If���eӳ�*F�1��;)��#�Si�w�ݳ<�͝V�M�u�g�����\��� ��H��)~���ך���
���l&xk�,�����Np�2�r|eL�2j��7��o{5,�_�^j�|>�bӹ_6E�p2^jb�c�J����z�����NuL�\j[�ַmZ;Qԇx�I|�SO�}ڶ��W6������4�I*Y�H<E	���-�N2�w��;���h�TS���l�=ݵ_\ �(��+�z��"��6��p��v���|�󽯚�?آ_/���Y?!����r_�FHB��W�K&zj8w���k��їren��|��#pSLAt�����4��А��(�y�y���?c�"�%`�O��V�b9�M��G1�.�N�(���e2���u"�����W�=�<�^�U��K��+�/g6.�ؾ]���"�[�+H��Iy���k���l�t6\�W��;`��ե�E�wPtٰo�j%�����s8�bm��`�B�����ޭ�a�Q��W̍�<��|����h�"k�o �u<�!G&�e;v.�������cF��]c�ξ]O�}C���_�:�s.��;=��pVż�vɭ���d��;^^�闥��㷎��@w��0��I�b/6|gޤް���P7�`? o :��.h.�6͙���~������3,t_^��lg]-
'�T���WŁ������/��Ob�>wPkt�X6�,نa�ON���s�ryjw���aP��A��#^;j�h���4���8GC�lZWrۂ[�=��;jy��U��:Љ{��,�ܦ�";SlC��{U���'���"%�_b�d���W�,�5,�zg5�~�K:]�{��q����;.��9)k�i�!sn�@���k��u���<��a���8���#�5�4bH�UU3�D)x���U����>هϼ���[��"n} -�����:#�a9+�Ul� �\��k�3�"��n�ea�ʵ�1<4�oU��{���v�xt�ܳ!$�z�M��Q�:Ǯ�j0X��ۧd��8��Ÿ~��L�!_F���cE��jۂ-�\`o�[0W�%SL��b걪���]��0��c�e~�L��{�~��on���rV,X�4���rS�O�ϱ��	�/[^
�&!�G)�"!�I`��{��mY���i����}�|S����x�}�V��M��&�I+���geͽ7L�j6��N�_R�z�"�b<�o^6�Ei�;F̿�C�I�~5����b�x��*L���~���i=v��9��@+ŷ e��환�؉};gr�H�n�4�r"ȯH,�dG9��֡!G:�L���6{�m�oJ�������MAp���,�5Se��Y��4�IB�A
�:i��$!�)�s�FNT�B6m�gN��pj�{�|gj ��'�4j�8{O�.��zS�P_K��T���\�m{��5�cvh�]U�����p�Zhw*�vu��|.g(oZ��z��ʟ�F�Myf��rGI�/L9N�_���/�X`֞�M��8U�v~Ub]��0[.�g5�q�ṣ�Z�I��Dw�'�Mr�%��u�)��_ ]�n�����^�2W�E��~2��R��5r*�/|�0��yf��B)�?p��xe9��%���l�m��_�	�y�w]s�6�Y��0kC�>j.��="T|��_W��4Ό�KDg�a`��R�&`O�ap)��w��՚�S[��-�e9N�'����!��;F.����)��<�k�k!`Șe~ޙ��_��0LLj0-~��Nb�'O/���\�Z^vfT���O�s�@���k����z[�=����[C�k0�Ƒ���j���!�Y����͆��.����IB�P^�.��֘+�����T��{�k}Y�n�f~2�j��cI��L��і�.0�!�;�=rq��N7t�-�nAg��U/��d`w��s'Ǯa��0���ط�Q�7G=�N�!��&b����׷�l��j��.�	�9�-8��:ۈ�ݷ!��	�ёz4��nGMo�g�1�M���}o�_��^x�=��b_�bٳ��i��-���sb7_����Zkڍ���ǻ|&���<�ޜ�Bx�)�᯶y�F���e>p��<A��o�ݷYk+�b�Ԏd���Dݙ�u�Ә)�J���M���L�F��g�Ƿ�x9�NP,�jy�K�:xFHi�v"�sZ1]+{�g 'Up�S8�M�e�i_*��{���=+<�_��(fvpR[�)�9�g<OMh�}^O8׻��B�!¯(�uZ"PǶ��/L�1�E�r{F(��6���Y�o�Y�-|��3M4W�J���ʛ��t���!
� �!;��1�b�3���4�n1���I��k��TӮ*)�"0�T���/+˫��^�!���ʦ�L��}���}tڸ2f�y��ľ�0�	�D�N���<�S�3<����ئ*z�<Wt���T4�=�1u@�kC�
�+�����"?Y�����T�!��4��b�z<RT�Zp�C.��7{�9����z*Ϋgv�c��#ϯ�d�o�=�����m�sDA�0�_#��MX�0]�,�t|�q�)��䴄�
phg�x���=
3wK�Y'�w|��0�:�g�=�!�֊�n���f`�-�t�e�A�Umú��M��I��n�X˨�#" ��*�%�ȇr��E�Z�h�g�*��dv��1�l�R��;m�bm�z���+����;��|������|_u,�8*��p����0��R���'i[�y���s�@�a�����BZ�{�Xw�W=��~6�D��0[6���U��)��E����g��f��fa��_�(��}�d)���g�WQ �D?q�������n%�"|b�6?h|?EU7�ܷ�jy鷢pW�z]�Y4�;�5�>SUq����\�MsqSb��$բ�wF�cs��*G`+�>��N@��OK��ٞy6��o�QH+iUw#Y��Ѽ׽N����-�ˑ>��ךi����6<5�TDj�g�8V��ݐZ�6���qn׉�����[�7l�{�vmF�Ιs��y�p1�C�t�Y�n��V�T�7�+��m�a���!l���7;��^��mA�� G�[�{�J��P�ʄ�F5;ů�i4M����@򽧆x,���-���o�ҲA�>攀�FU��7�c��}Z'U��%X���1eJEVG�,��}��/D}Z��EQ9�n�ծN�e�C��j�<�V��jt2�&�R	U��@,�c*�A�cʹj��ʠ�7��og@s��Q�]nw�����L�c�*/�b��p*���ݵ_�� yD���:m�s5xYߞO�����g�z����J�4�iJx�Y<�n�O�_��K���w Y��M�7V���_6Q9ş�0�eȅ��b��.��ϯ�!��P����EJ~�7Vy)�0mLVb�����T��0�'|Ѫ�S�,���j���3O>ͅ���#U�78�����kZ6�Y�·����ż!^���*k�w,����4k��)�S�A���26�6M�ɽRm���7��0�T;ؠ���L6���K���ߊ�.�h���:�L�-��W��F��]���̹{�{����D`{h!aE���M������M
'�SA�G����~�7b鬊>۝<)^�Gջe��D�T"f�~|Έ|f�Ӡ+o:�wδ)��}�}l+Ъ�3A�����FX�y��RIؾ��y0�ё�e]�v	�u�z;v��\�z�/������i�Oï�VC����Kv{.�5��I�룯0�~��3�a��z�~o���g�g���=ۡ�d�ů��	��i���)u���pV������C�8;��^'Am�ގ"�s�e�
Q*�ROk�����8%lp�� 6�,]�7�3���b:7��}�Z�z���3��=�û���*[���&�<p�gQ&[
����+i���}BA�CD��z �W���%#SoN@���1�\�~�4������0S`\'�5,��G`k��$��=�WT�:�wQ32�P�)���R���\)�W�� o7�g_��3�4�`Y	�L�z
/��s<f%�	e��;��y��e�\�x_�q����/��;�~t-����v����eI�F����ǵ��\�z�u�Ϸ����+���~&3Ǣ�i�V�j� [~��8L<3�;8T���oQ��M1qt�;�����)w���)��!(�~���K�7omC���vO5��En�Fv���g�x�Z�&�-�DY!3�+"9�b�{A!⧝p�t�\ИAp�6�a�;�0f���R��m��p�2��j���64�IB\�����HC�����uuſS^�0ket!�Ȫn�6�[h�p�5�!¦��,�6S�|W�.��xS��3f�)G�Au�{�V��^�GF{�^n�MK��7k�W�@w�Z|�}����b�q�d�'�N�K��[:��t��Q�k�)��SGp��}j��5�w/f�����# �f�q�Ċ%���0���#�[�f��ʰ�V�\5a��!/Qm�'�����U�)c�c'Ǯ�?:48O��&e��%�ک��NsN>�;#�Nk�Gz�@������ם� �\}���ЛN�X�8\:���V�f�w�OzG5��ٝӘ;����q��W.��;c_|aN�X��3.��z��������Zr��i���i��;���	�y�\s�qn�RǆY��1���n�ߜu�!6����W�F�a�{�b��R?`?-s��zd�)�?h�Dg�a`�pʀ#}���s�U2��&����6�����;��"�}�c�e.��z�Ll[�������q5^����e�>��0��ܲ�y�[V@n��Ӱ(�s<m1��n2p��u�[C� �ߺ��ÂS�ώ�z��+����6�s��s�3O�MѹMW�/��"�N�u4��W4��ra�jC��n��M���*��쉙���o��'���眝���
q�6�����;��M�ymw�sb7y�m��k�>m���a[�w��w�/i��ngHDY)�᯶y�������\����y��H����[��k��73����2U-vr�I�8ݙL�Vz�� .��|�f[H���<C���y򱥸���V=�'V���nޭ�^h4�s�n)��"�5zT:1X'���N�x�}����<��D�	���t�u+hIw/k~��cV.+�9Orڌ�� )�w��< �;�O�����&��r���G��\a;i�+���O����Ƽ�.Xta��&K���V/gp'��K�:�w"� ��{O>�f��Չ����c0K
۽:X�4!�b���MJ~�`���-֤8T�m�6��1�.K�L���i��]����.�I޷;͛MO>�J�GGFʛ��t�ף$!���Jw���>u�#�,����# q5s{��F���~�~ᾓ���Q���m7d��˫���\�-g+f����_./�f�	�?{�m;�� XTs��8�5Oh�JC������Od�(�&:�q����y���� ;��hq��,���S8.�S]F:�ON�`�-GN8�{/*�Z:����}T��=|�SX$(��%R9F �wΌ�ka���WU^^y��0���:��s�3-/O���`!�@7�m�[�o�=z�@��2�4����b����;�r�TLU7q�h��zL����fiJB��gδ%����Xw�Q�1��~.�_-�rۉ��ۜ�n�"*��4Oa�	�S��;3;}/�w�,�4دq|�~U1���?n�*Y����1I��i����טc=���_��?	�'�^���,�~��n���r|��������U��Y_�,�����-��QW;*fZ&wK�H
 ����c�dݼ/w5[Wڙ��J��:�+��G�l��ދ}�V4Nӛ�N�e�L�t<4j�{�v�u�`I.h^e��믧���v��b��.�Z�s�Z�V�9��fT
:�����C{1�����u��f�U�V�r�s��2�(�j�u��w�V��,��fgsշ�h ۠볞�*�Y��;�ts]�9 ��z�ͮ+�:���V�T\�*��o8�c4k�G�z�6K��W<N��<p\r��^��;�Ն@��]U��TK�(�p��+k�2u�-3������9'a��ի6��[����y��z�.Yk�ǆiNBf�+���Ù}l��3֕����;�X�;�xh��{�V��j���M�#;(;����~��7��L�n��3�rm���gO����́K��ԝB�n��3��7u9n�A�̶�W!M�}�}q��\�x<s�=�	%�U��c�����]xvq�D����;s��'Q�U��ˣ��=}6�z�|}|;��+<_V�V{�:�w�[�@:m�Z}�0L��U�������,��"�N�]��H:}�e�g�m��w8e0s}�-nh6f͌�A6�s�}�rG3�)�M���կE%��;؛�o�G�ک^I���^��|yRޘ�/`,���l�/`k�����Z��6λ����[3�0��Tn��LH]p}�v��Ֆ:����lR[�D\�G 6��SFGv��U���=u|��h*�ҹQ�1WM�$�^ǤM�jZީ�^��hQ�y�I�\V�\^ f+�;()������k���X���X�┅z�mn�N�X�9ٝx��EM;��D٦bW��D �Ht1E0��δ�����jN^u�p<�9�����\ҋ�W}G7)}��B�r$�dݜ�\5�,<��|�cM  �&�U���]�m�	�(�A�b�V� �X[�1r��<����-j�����QtJ��%�v��%�4b��)� ���5p����w(��L�#=9C�X�����j�iPa:��3Ǌ>]�8x��Zr󮔼�DU��N;�u���,�1ҋ34��ن�[�2�T�wg'
UÔW��v�:=�[�lRyt���
���;3Q�V멳�]ncɈ8;O7��,�����T��.��-�[�,ee���gZ妖�ćBk��;����c�����#����!d��e��#ɬ�4q
����Y.�.��U6���dW����v9��`�_oggk:ztr쩯�.��M����K��GK�Z��U��i�e�,�hF�)�]��^��/��l��b�<�vp�%z��qp~�<�w��Z�:��'u�c�@245�σ2���-�˵��3���Ѯ+yN���ҿF����=���7u����x�J�&�iK�w>��Ga��t@�u`c��r
���eED&�ﻹ8DQ�;)�!QE\9tB�q�**���DAG	�9r*�:�y�QHD��.^tM�QȢ�p����Dtª��8$�����"�ES*�: ��&��"241 �����QT��G`VE��Ut:	b�EȚ���:T"iGT(��hf�"!� ���8U)�*�TdP�K�t�$�r����\�w�B�ͮ%$u��()��R�B"
̓d�g*T�%"U`E�2���IQC�iD�u��lȢҴ#5�se�"�UI�RVEqE�Y%�t��(��I�L9�Q����[���D�fZ�p*Sݹ�je
%BZ"P��g�*ͅ��b��3C�UI0��ϓ���ǿ>zL4y���Zۇe���M�~I��I��|ePue g�ɢ�[��B��Y�3�m�}��3�\Eq&-����Q���Q��[��(ݦ1�v3ސ���F�rX$���؎y�6��`L>� �}/����o\�w�x����D2��y����g��TDj�������}wwd��kD�&[K��C��O�T������y1�7�C�9��[8#�r��.��G�>�Y�1�5�}��9����ʗ����o�^�[PE�+��|�(K�#�;C'���ѦloNة6s	lN�����;���4Q�EE�����`�j�wmA� �D��wy�v���Dپ�[;{�4W[��_
��~T�0��tK�P�,�C�y��?!q�%��d�/�>e5UMD�]��� "Y��7����!`���r��DT�f�o�!���q�}�����7]*.�q�o����:�y��i�K���n�N�U0��X!���Au^�4�ٰ�^�v��������Dh;G6s�͇j+��H+~�x�i���̻�g[,���CE8+b�_�{teN�{��R�:��-}t�S�/�;@��a�3<%סL�)�4;�s��h���:���]�y���R�c�����Y�vŌ֍̩o�>r<M{�T�D�apݩ�礆��9!�k����L�����'�#5�&K��Ž��8����)r�� �J�.[�,aX�R��Z�Z4��f�U|6!�h���ч�M�����
��:d�'c/Kq��`9��:��{d B��+�����}M� �[���\-D���X/,fh�8p�ѰP��Fk6C�����Ѡ#�uZ����E�>E!,ų��d�TS��vjߙ9��I�����9"�Y��߇iH�m��1U��98���y
�T5��w7;��H/P�R�����{��I���y�3�?3��\L2��z�ߠh���-����M�Wy������j_+ˤ`�dg C���>F?�8�M0��p�ɩe}or�wg*ǻ�uXS�,[��{n�ri�-l�<���T�׾�o����b�� ;�ο[Y�D,'/�c�����+������M�A�a�%V�1<4�oU��v�U��d��,�,�I"_��qn��79{f]i=�Sd�z�뇖��L�!_F���c�[�v��!P�O'��B����u��+ݼ��-1q:L;���w2إ�To���%��w�m'J�J�Uo�c!�,��>�����[oğ��8B���EHL���6)w��	���p2m��3�Yq�0.v%��j�ȉV���u��uȆ{��ᶞ��C���5��f�{����owV�W���ޕ�u}�G�^��]�E����V�5Vg�{�W�ׁ�$���kG�_\�3��r�7ޔ
up"��*]�VM���T&���+�i,I�9}�9E���r����m���"�5L��%�s��aF��](���c����aZ�M�X!��Cm�*n�6�[h�p�5�!¦��>Ѳ�S�YM1�G5�Ѵ��7vfrJ�g]퓽ON�S��GF#Wa���]U���E��Mi�ܪk�.��hw�\�uk\��{�.뉧�DG38:\S�*Nν0]:��v }}��EOR��n���v~F��nx��I�
�X:3M�;��`r]�\!��ڇ{@�gl�׌)�=�5�
]Ӯ����hl�|lc���,�)��β¢���5�P	a���8��F8�\*���2z���
����M��9�{ӭmuOy�[�wK�x��8��4��̎1}N[�4cDg��a`��xdr"�M�S�u�o��㶵�	ۆ]��p�w���r�~�L�jGm%����+�k!`K�HFX�F�kp��ƈʼE�9��y3������x�=R�_s8@u��}v�+�ev�����]�ֱ
��|�3N�B�l��uK"�N�KFf�yV��& O�nC��R�����1&�_�Vb��hw��d��M�>ޫ��5tXօ<*�L^i���n��gpT��M`�2&����N���jEN�?�9��k5=���}Y,ѓػ�&獽oR�Sg4���<��'xx7�����3��<�K��q��.��\�:_N}��.��ٯ�;َ2�'��rvS���f���n1/ӱ�)�[����O=����[����p�$t���C=�;M1q1�w i�S����=�A�B{᫮x�9�aF���x�{�n�=�����zt}c�)i>���R?^����xލ��28C�nN�n��R�1����ʓ�ޜ�\�^H@��{��2�.b,�W�C��'����>�i뻋i�{�]����0C�%+��MJ~�`����[u�(�u^��=���~
z����ד���ڎj�p�K天�dttb�,��M��m�$!^� �Q)�Q�����B�s�ٍ��sz0[��#pSLAt��4�
����Q���mvIx�K����\�2��Nu���E��p��g��1,Y��za��SLAu�꣝W��<�S�3<����ئ*Ƚ�]P>GZ��W���>�����b� w�"4����Z��@x{L��z?��`�,���'f��a���``�voy8�;�i���M4)��*��-�!�ˣ- Z�h�q�b��ᑞ�I���lg�6�=m>����x��]�0@���c�H��`��Y��Q����;�盚�5�7�с�rR��ާ=�����)��EO�K1��Vѭ��5f1���l��==l~E���½�
�ho
��"+���D����@f��:\=ּi|���ik����#[���@2����	K�����o���|� qA�U�z;b�.1�����Ί5�������=�05t�Ϝ��;�Xw�W=�̇�`D����~����ř�۾ȳj��~h9+]�|�b�~zc�0��/��G;�[!M6)��K<���� ���r��	�;EC��K���6sg�~�������ߓ�/~c�J�8�;��l�̧��g5�^v����e��%�o��\��vW���g�NX}�y;)�G`�z]������d�l,q3F�Ny�dj�iu�=�)��/�ȅ:��2������W������|3�������l�ߡl��9�KoU����xt]}�lZw+�ȷ_|�ճ��*�FUCŦ:���lz�Mi�.��̦�:C=zR�c��}�V���&T,��W����OŇ�����r�kCOϦ��j_��zL?Y��*gxk[��L�e�b���XCSwv�m� ���4�Ş���$�9i�� ͿLE�M&�d.u���ZҔ�9ޙ.��G\���vy���6+,x� �W��������ˀ{4�����a�:Q.��u�Sso�j�!�-бYl�+�`wR`*�xx�XI�t���� j��Տ:��0����^�h��jrr�ng�׫�e���j�����*e}�J�4�fu#բe^��������A%N=��i�`�3��ɸ���_uM�0qP��3�lj���H�� �(mDXb_�~lR��QV��yhiE�6�z
޹��Z��P���{���F�aL�H�j�.���;��H(��V����[UX��]��򧦐V��­49
�s.�Y��;=���pV��X=�vncZ����s=;]���,��~J;@��a��U�\(��&�U�w3�D>6w&���M�mA]f�h����W�}8���{h!l�E����BR�����#)sd{��y�Q����6���t��_�U�<�E�!5Q�{6C���針=:�u�hS[��_[z�����Z�[X9e�T��x�kA����%ۯaϢ���M���.3\Ȉ=Ee�h�~��v��{���J~w�S�@��i&7�:�g�~f��,���8_��[+������9P2���"'���2��a��d`���}m|}h�N�#^�p���d��><��L��女_6�h�b"9�y�������|-�W��� �l���a�/%c*w����|�s}�4�b��{��m�;ת��.)Q���β��W;�7f�S;]�G�+�e�%��<7�i��Jb�6J��j>�\��y��P{�m��Q�p1�1،Y:�u��p��#2��9�4)���Ľ�{/�n��2�ʙ�ZO`�p]��{����S
'�x_���ӽ4����'`n��g��e��s��
��Y��׽�<��<O��z�L���:�巵S9�Wѧ�߉�c�o��*���HѮ�d.�SD����2�?Jk㟟�t���y��;�Y�L�����^Ή�z���܇�����ߛRʇ�W$LZ���Q�9B�#�ױK����=���C���X�Mi�V�R����yN@V��)�>�o�?�wҲ�Wʣ>�W:R�U���|�5�~f��"�b�ᶹSv�E!ŴF8B�h�p��%;ϴl��1d6��]3k�3�S	4�2�0�B�t)i{l�Ttb00wa����\�E��Mi�ܪk�.��`q��2�������n�Q߼./DS8\6�qN��1�>����u0�Sԩ��@�V��{"L��j.�֕�����g��b%�]�û����m\�����LaN�Y�5���0QD�V����^�s�_~Z�1LTP	a���a��h��8�\*��dtm=:�G���g��Yuw�.���7KM��GZ;�mf#�L:6�Wu�����?����=�>^D>�2��޵&z� ���:�F+�浽�D�pW�V�w4*!N8.��݇�Dg�l�Qc��D ��k���
�v����Vѫ��= ��b=�J��E�}�@-/��ւ�ڲ�/{�<��������^s�R�Ϲ_�A҇��:���Y���9��i7l���s�a7���d;@�^=�＞)ߌ
[���	K�?�S���(}��`��
ī���c	~�&&�t���i�Ts<m�|�n20;�7��'�a����n���e�Z�TnrLeV��F?4����d�:z��e5�C���"�N�7u4��W4�n"se��*�쫶X��{�������u�y�S�`91�|=~��+z{z/�K��g
|��M� �w�J;cKf�2݋Ȍ��g���M4��
���Jwx���=�A�B{���k�M��-v�7۬��9!}��6�M�u��T��qӘ8B��i��!3��3�P�ڟ��9�V�e�
�{�[x�~3:����|�f��z�{n����3����e>[J�T~C܅�)-��?����듷��F��e�/�!^+�p�7MJ~��S�SwGh�/�Hp��&�V��1ޢ�m�|�xዪ6������1��.��*jy�ZJ�+�'��m�*n�a�d7^���7t"OϏ�X��fa���Q/ao�֓t��3��!v>ȟf4���[������w�˫DmpY�j�%<H�㋻pyf�g#����b�d�#�>����vȭ��O����!�Ǫ[�C��}�s�LJ���/�Q�7r�3�5�/��������c���!`���j�r�zLS�g)O�إ�e,�x�L�WSsCfގ̈́����Vf�m4w�C��L�Y3�lq�z��X*b�U�c�S�3)�6r�>(�9&xt��U�Ϻ�,�����g��C�PZ���[,��\!���R-ў�Ѽ�c3y��H��
Y[���[�#��=�zbxN4)��*��0s���D�"��E3��d��+����r;F���n#Z��Փ�(�`��|&����y�����=�_J.�[kk��H׾���o��Y���E�]^"9�,��Ӛ��s>rxjln���@��2��u_�Fu�+''���^;5z��_��c�;[A�ߘ���_�l�SM�n/�ϸ�Tװ��8n��݃��WD�����}r6.�y�v���|���+~O����=�����t�|h�|×��$�̓�5V��Dr�g�7i��rsHX
l�F�|��N�����*/�l3	�S)ܡ��fS���K+�`���B�|�^X�9Nܡ^���}�V1��]7D�E�y�/���D3h֙.��k^ 5o��Xf�Jَ�g

�_t���Id�V��d�`��s�G�[-�
�;ys�yo|�j�zer�q���qX�ĵ{���u��K�����d��e|$��ie��p��ƺ��]�yCngoTߪX<4|����9�KoU��v��׶�ͨѹ.��`��L\�s���&�iT�!D�t95};���(����׻L7�x3�AT�Z��|�n���Y0A�����ʗX�y��cqfd�7��t��有�M=A��tk3�5��h��P%�k�����PDU����N��zv�� �(��+�Տm1Dpw+[&��Κ{J�ڞC��d�h�����Ս����O=Ny������ T�%�<�ƪl��	�29�u�f�o�!��N��l�~��(£�}`,�O>�M�~�`*kR�Tt�5S
|���"穘�%��~*���f��J�Vv�^�@��00wd��(��o%_�>����=���",�S��v�2Wdޖ[j9�S���@���v�}��7�����B�ܚ�W�K���PL��qȌ8qD��/��i��=}8���ry`��
n��z�����0��;���΀�z�^|�x�>;�J״�py�dpw�Fo��ƽ~�^W���lcm���lcm��6���m�1��m������6�덶�6��m�m��m�1��0�lcm���lcm�X�lcm���lcm�6��A������co���co��6�鍶�6�덶�6��m�m��m�m��co�����)��<���,l�0(���1#�� �U	 �*� J� �P (�� H$<�E  Q( QJ�!@������Y��ͶT��ִb�VJ�4�}�(�[Ma�m-k-����f���*ֲ0��:��.����kJ[��kR�kX�*l��6�MV�S�ݭfV�l�*Zʤ֬��ʬ�ִ���i�#Y��i�Dɥ�՚�f�1�5*�mB�kSm*���`m��Q��bѶ�1Um��-[[J���nU]h�Ɩ�� w[�(�_X���]{��h*�m)�K�6�j��!�طdp ts��w���4;�e 5v���\Ψ�i��Z+ևb^��Z�[l��M��m��  wW�馺5�O�=�GQ�gǠQEQF�1�@QEQF�LtQEQ@P���QEPox}�袊(������Q"�nF��(��^��Ҕh���V�Z�@���d[bD|  ��Љ�m�>޹�wi�nt�{�]�^֝κݕ�/m5���*��u����zw��ٷr�/^kԶ���iz�ޮ��m�v���[Zv�5u+�f�]jڽ6T!�֩R"il��|   kҺ����]�K�� GJ���Ϟ���m���ڻm���V��T�۲M=�K��:hu����ŷ-lr�,����/n^��"�Z!���ʚكmQf�n�R�K|   ��w��V�4��ؗ[�껳��W1k�t[v�"Ϋrcw���Ev���hZ��ۓۼ�f�rی���[�۹����j�t]�8n�[uһ{Tي��#(�"ژ�I>   ��u�Z��wW3�]�Wgv㻻���ou5����Z]�N�wSNi�p��ٶ��ȷ6�m7r�Ӊ�5f�uз7��O]�Umgl�sR��mkQ�z�u�R�K����f�BٶK6�M�mTf���  �/|�j�n�glw4���m���n�W���{��ݥ��v�RU։۵z8^�OMt{�m�����ݻ��:L;��tr��:����݇jG��W����O=\+55d�e��Y-��[MZ��  ���6�8��ݕ�v6��z�]����]��9[l+c6�]�b�:��{m��ֻSv��w^�{ղ���m�s�W���7u�Zvw]�-�Ӭ�6��.�Y�n��Kձf�[���jJ�-���  g��Һ�]:������I�f�u\wr�iwi�W���[oM;
�]��m���u�XZ�[��5��s[)V��T�u��w^�e�MG���
=�xVFm�c�Y-�)�+h�  }���ӭ��mT�飣�N����4ݽ��WT�Svr�����])�t�ꄍ'E`��9,뮆�;���RT�� 4 �~�R��  ��Ԫ(   �~jR�i�42j����UI � i$�l��� �~��������[�Rڸ8W*Y��u������g���g�H@�s�?���$Ԅ ���$��B��@�$�$ ����>c��ٽ�z����o��&�	���gc�8���s5�+�c�)b��"�f�؝͚.�߸f��eC���Y��I�<�B7�{Z<p����.�PD���su�\k˫�������i�M��=���,c��lL������CM�M3��s!������[����|#��62.���<1��2[��>�䴦8gP���>d}���N��켕�h��z�[�_ ��${���e+8��Pb��Ӌ�`��k�׸���b,+؞x�OvO���u�#����f��ӳvS�ǒ/G�av�c�>�斞�k�MG3�Ǽ�W��/I鸦N3���B��qf1�@�Kp躚N��t���xط۷���p��~�(V���'5g�ZT��9r^�;Pj�v4m"���k��,�y�PI/].�PT��ulY��0���\�5�:���(\�K��-�	�;2\�n&��},��^�(A����`�y��ѭ��Q#]�SЌdr�����U���=��*v��y���B&�Z4��E�^kٶ<
P90�y���>����#���bH��݃���j.�k�m��� I�k�֢̨rY!8\E��g ��3p�K%�xv�)�o���#ufCw5:�B�8NR�"�).xٕ��Kw�cM�w��=9�5a�zssWd�4�r}�%�*���cj�̰��V�s)�B}��l��bdۏg*+���W� f����m�Q��b$��X\���4�C3	�;C�Z�ֺh^w3���p�5x�'grFn,�ܙG-,�{�q���l�遪E۵	b&_T�u��q��twt:�s2-]�:g�a��R˘JU�|3WD��	o�FB�ICD��������q�cQ�!^x�5�ԇ���n�i��0��ӵb�Pٍy�Rp�ݷm3Z�Z.���
V#�fe��������^+LZ;�zy�Y��>�+��r��%��jM���N��f	���8��v��N�nʹ�e�4�)�[�xi�*�ܓe��1rno�J}pj���9$�'��[8���Ǚ�����*0̲�D��e�oQ�e�+kg���c��q� �̨�C�VEa+Z˲լ�����1���-ڼ�fra�Ԇ�B�r��,��J�y-��䩆dR�P�6�^�}���uP��g�x�q91É({�]q�YH{�rЩ�{�ɽ���=@f>s{;S��C���B(�]Egnfj��b���;����s*���y��;�MXr���ie��3�g�:�ٛ��kN�g0�μ?c�!��ڃ�L4��R��*��ǏN���qj���H�&85��E�ނnn-�u��	��}�JQ�>�"���b��j��ө��vS���'>A
v��1ooN�Bô����N@�1�0�i�wu�|���i�ӓb>�5�2�ͥ��7Jw[�c��<C�g��"Cvݤ2�
�g�0��e���wd�H#����~ݹ�'��
f;2a�7"���vl	9�w"�����gV�ܴ�/MR��a�w.�L�G2aU�;eM���k�Bf$�tU�+9L�k"kc#^��L6"�ɻpci!I���]E�6��^N�ǆ�粨�v��b\l�d�Z��rVdN�ZCcsU6�BE-9�pl�(�g�(�b�	ݷ��.x-m����rvŸ�;��$�L�r�
�k�Zޖn�v��<y�k�p�CA��5R�tN�c�5z�����v�N�j�E+m;ɀ�XZ���Zm��n��'	��zK.�N���y�\.현���K�^�$F>��zCM�֑p)��1��ST �wmh�c�c'3uǹ�W�0`C3P���$����h�w���=���:�'h�,�u�����h�:,s'L��#r��a�����+ў�wvgY˛j�Vґ�������H�K>�$]���.@�3��V�7K��Q�G	�742�^�
��ya:r��?�Z��[#�.�Rg�w�v��U�]ݰ:Gm()�	35���J.�H�M벖Ğ�Xl��[͉�[J���X[i�Cw�8cO��o�:��y����;Ea��F�wol�ŧ�G�s����[h��4t���j"�q�������������0q��-CX��:��J����
�nu�.,)ɝ�P��]��S�ǽ�k�1�WQ�ә��M^�X�^Q�q[��ZFE��b���Bn�q������R[�X�4�`㽏������
^�5�U��b�$ntM�����s��F����M��%�93��/<�]8�m�|]�����2�}S���X�yӪ�^e��:���#T�%����V��J�r�*��,͇q�y�ma!V ��$6S�%;8����B �wI����-ct�"�Mq`o���H3���7�Z��ߝ��V�'E�Jw�C�_��Sծ�w5SxV|'omҹ���0DRЫ)T�%	y��i]�L��{�c��%'8'}q��������v��C��Ʒ�,���N܁��)d{"��[���s��*§�+"d���L�����j{�^@f��Kn�B�B�.��f+��m}� JV懌�����5�N�ovnb[�Z�3����98�s�7�؏2b�F)�Av�/PMW�4��B#����척��[����O����z�Ś]B����onm��8�+
��n�؊�'�+��ǥ�����齲�P�U�.9ջ�����w^E��U5q�^�(���������E�������<� �U�s�y۹θ^�앹��Qʎw7��8�>[��K��Ԓڝ����V,S�p`6:�Pk���o�i.L����lѻ�5��f�c��rKY_^�`�l�Fk㕊=���7[לp��Q��*[o&fȈ��I� 1�d�O0�^��L����=��R����Ζ�=�Ԑ��0pg��;��S�hvA�m��핔��&H�&�L�kB��Ʒ0�2)�Rp��Z�Af����SE�d���ss`�Xv�)�,ͺ�'I;�(l8L��{M��o�	����0�L��e4`{ġ�v��5��Gw���{F��s�j��*��0�޷NZN�"��v=/`z�k�"kcX�tc�Qɷ2�Q�.�rr!c���P_aY�oq�/ͥX���*�L��a0▀Z�v�,Y��yۢʒ`�����'��0���6v��ZN�(Ƕ�ѝ��s�4��7�r�g�g�<ٷ���SV��Z�B��7wq�g8z�*�t *\^$��A�:%�-�vb-�[j�����ձj�-b&�A��POdW ��f�Y�Z�,u�{#q1����S�2�m�ϩ�]������+p��7s����_Ǆ�F|6vꗶ�}�^����4E�!֚��g9ɫzmp�=x�b�~���w��vƒ�1t3j�\8ܖ$���Q��s��Ա�!뻆�*� ٷh����fn�OPGgc7�iz~�ee*%��`���rL��8�ɨ�&�6o=�ɕA�3�}�;2nSS̝t�KYz�q�.cgB�u,��U�۽��[�)�b%"(�#&��3�n���θ��ɽ����w�����I�[xѨmX1]���$D�U�&[�J���3$�y30�tW�܉�p���/�yy߲�$��,U��4�Ȣ�E=LfiCKHMV�:B�N�I�ŬUެ�a���q��M�`�f���DD���NlO��O����;];s��@�<8�7���P��0L��yeu���DWE�v�1t��'rɋ�SLt���yp��28.��UAh�ݒ�-z��ݿ7�#�X�ΏH�'RZ�
[Iw����	%��Ci���k�o�7��8���Ȍ#\�=g�R]71ɼ1M|��_��J���]��r�u��,A���D�F޿C�nŤT�L���Ӊ�˹�
V�B,2�V-��:��`E��=�4�ܩ������3�͒�2���c��`��E��sb���b��83�:��9$y�o�s�^��C�4�C�l�Ay��`�iǖGN�X�V�̗%+�E3���K)P���ٹ��d��N�jZ�B��u��M\6
��̡+Un�-�]�m2˦(/�k�
Q7�����h�ӈ�/+��Ʃ��%�z��U�����롈�7�{�n����8�`�=�oXa�6����FK���T�a(�Or��[7�Ҁ�on4��CQ�A�K��3�<��.D$op[(�dy�Ǳ���/-�-�Ω����pɃe�aO2�6v֚�6�{e�d������f.<�ù�B��za���'Nd�Rt�.SP�Y�DvfJ��wSܡ�:W��%�D���;{f�=IƢ|9n[���f��d��^lfu=�8%qv.�ڞs���EDI��k�ݜ{�9��B��1
���'l�8�cʬav�ɟd������� g�������t��ԺrM��[� �9l��8�Y����"���y�j3��`̹�Χdp�e�tZ��QR��Ñ���_^!W2w]H�o{{�&q)룁;�.ő`����l�*���rB[���qe�Г������4��9���ojw;��E�y
��p�ES��nnk��}t��P1C��I�vh�Iw�,Z�&��b�!�Ϩ0Q�u��u� ϯ��Z�a+�ofV:6���C��F�D
��4jz[��v��.�ĤI�E�ݡ�(�qf@i��m�h*Lf3f����ja�f�F�Lz:���k�d8v`��6SI��FɈ�wb���ݑ��a�Ҏ����P��E�W�d*�sڑ�7[WJI%k�lV�Zmݭ�������n�7Lw����K�C{ӈG�zre�ѱ��ѻ��5l��d�o]2��1Nu����e}{�{�'�V��x�u� ������N�z{��"I��FP���^�ZF���K.�+)#aӣ$L�@=!�M�{��ϪS4b��]M�Nr�7��f��e=/y�S*��g�^C�[?3b���f�osݶQ݉+B2�9r��@��!V�,1�؞ߪA�״)�;Wi�Fns����6�W�H�q�Y7�i�rܚyˈ#{��/jjq�>d�V./J�c=�3������Ȉ�ߎ`^8���B�΃�%2�1ҹ���8L��㛡e\9�ӓU��"v���kQ��O���e탉�����q����c'z�����r���e!sn�=�lGyE�^������4v�в��?�טj�D���2Cp��Yf��0���ڳm��5ҵ�v9[j��N[�����΋]���gnL���芪wwNv�������b=���W�Q���z��[{����P�pKt�,�H�6�-%�V�Qh2ɬ�0�	г���6&�󪁬]�W�h�[����s]�jغ�[��]�@�*b�N4�@��/F:3�����`�����M�H;w�L�z�,�;���ܪ�1�ˡ���Y˟mssn�C#N]�m��5��v���4�*�Z/��=���Z&�֣�f<]�3�b�B��S�[aKt���F�k-�gt�V{GD<���+�y	�5bޥ-��i�u2��q��7�|y�i�B��"��I���q�g,�˚��pfC4�4��U40�j�b��f�����s��K�s��r��x��wq�Zx�s3�=���_r��1H��Ƀ޾�A�[���1e�K$-M,G�x���6�r�r��N̪.oK)84�VE�K�ك����Ǵ�9�N
ff��Ww6v����Y�L��=�W�U���7�;x�N�֎�=cZg��L��+m�d��#}�x��%�ő9�u(�s'floVmᮙ�� ��(\���Ҥ���&�iu%������zT��%��^��w�?��6ǆ��q��ږ�'���1&1B�M�ݡ����b��ϱ�y���[���g�/`H�ːv���|P[��1ʑ3z�9��C�Sb5;w�ŗ�M�r�%8��{�{:�TA�`�Ѯ��V�zGN��z�i�v&��VXm��^��	��v<�8<��u�8���6�j`�Ba��Љ�f.�,'m\�4����ja9�}�E���9KM1�ǯp8�;�-8�acDEÜwI[3۷fZ�B[�D��P�{�)	U{�VzZ�;����̘.��߬�Z<��s���`��u��R\8[ז�f42\*��VN�CD�q���m�Z��B�k����x��]֚���SP��$t>��	��z"L�f-Gt��r�)����%���L��Ƥp�w��p������)Ȗ����b��.���.f�&V"!�U���i�[��;�N��:��`Y3�&�Ĭ�fф�IOffQ3���P�=凲q������S�ʡ��)�3�#��p�`�U���c�"V*d�O&�]3Q���EAFGGH��s�G�q��S3ݺ�k%��3�~Wn-	]�.��Ijke�a�L��\�	ۮ�?Bؑ�fT^�k�w���0�BÅ*���t�[Y���0Hh�:^�3����h��ϛ�w�Z�G�V]�-jJ��.9��'�1X�)˨�}�N-�"e�7�Έ�:$[%����cF�A��K�z��f9��#�e#C��Cv)h�Rj�τ�@�r�x�8kYO_����/	�Ne�a�p��foX���B�%�2���;�!,���Y7����m�nwM㜳TČ]@L��|wJhAi�4���0C�����m��W�{��y+��Βu��#�{#�O0ޥXmٮ�gm���'�;�뵞��ŅkN��
u�{ث*���$�;2Q�[zr�4��ڵgPm"�wӾ��pN�`�ϭ*U	�z�syp�ͨYs5k{�zv�	�+���U uXV��=�j����5�Y�x��8^���Kߧ1le����`�Zt�;���զS��:U�y���x�%�Br�s���P�R�$�Hs.�L�#"��5(�Qm��AQ�z__MȾ>��gh�b<��a��ݷ�%�-�pRx�
��k�mX�z7+�2�eFy�8�0}�
���K�l��+͏�'\m���	X�0O=�����+(�$��=.!���#Mr��n[�:�0��lY�J�����t����������,W���+�m�e/Ey3�^����fקh����/-�1s��;JX�|(0�� y�ڼ[1��<U՝��L�.sz�|8��z�&heE��н�
���d�|4M
���`����&�J�DWD��$��=��S�~�b��{ �Dj���X�F�`������[�N�M�&�D�zF_m5�{Mr��,a�����&P����Ѻ�Z{`.�n�W�t����D��_J�`[�Dܵ��_*��dG�+������If�P�k �j�9���&]�}��a	o�f��wCQ��}��i�d�+{:R�*-T{;Qΰ��A+����+��h���OL_���x������gv���%�k:M��oN�Fl��{�*�a��'�"��i�vM�첝-�|ޕ��:yo>
s����i�(#�Ž��#�v¶_0�J̬�@��}+�'{t�Ņt�U���9KN���Ӷp�\���B��(5@���1��c���d�����I`C��*<�V��Q
H��-��"��/ٹ��eld��������Yݝn�����������Kk�ېL�jtA�o��W�r�JK�#���iPo��^S��D�Jډ�WJ��&�c���L.lB�F.v��CK�Iݺ%�����%�~��=L��df���7�޼dMV9F�*E�ʴԼ���\��t��S�,r:�q�/HaqM �����_vvX�g�'i��6����'p�u4hxh���Y6���[���Z�&��]�2�����m -�8�%�V`�U�=tč۽u�*��ܽ\c^-n<���������Ubj�;<���u�u0^Ė�۾��t����W[}��$ȱgH%�폒��R�j�K�Ŕ���Wh�Va@��Ut�,�������n�t�ʎ(�F֍���bO,>�zQ�{-����"���RaY}m��K�]ƊW�uP�;�-��01ՙs�Vc�u��%��Y�j�(v�((�n��Q�G��Ƴ+��)cҵg*V�V�AKU�[�$�i)̺#r�>K�+Hlǈ�ι Uz�n��'b���A�x��̓	���Z��wu
5�*��F,��;i��fM�e�t�e.}} ܺ,XJ!9bh���䩜bX�'��Zo����i}
�7<�żz��*M��lI�e�q���c�[}�>R=
���nX]��)OqF���<�M�D������OG�|�x������^�
��7%���=�����W���\l�w:]�2�2���HJf�kog����ϖ[/FrG��Z��yZ��َy��Vv�%�3���:���� U$AU��Â��k[�Y��sN�o;��u�����RoܵE
������Qg�z��e�U��Q�9n��QeF5��\���^T�����X�\��h>~�^�R�^x5]cWK�k&��&�{f�@�u컬���`��8]�C��g��Y���Czv tuʼH枕�]��=8Q�Dnç>�eD#�qt�e�F��C�Do�j!A�[�dŷ(\��u���
T��`Ⲙ.�Qj�+�Ѧ��7��p.c����53y��5�g�2��/�M�J�� � ˨ %��_��-�)���W��@�X��n�Z���-�)U�w���o�wUtaM�4XŴ���6�5{���Z�l��7|�!Q��bQF[�sRg��z�w���6N^�L��2�Μ��!}�5�;rq�,$�v]�	:����@�)��-Úy�Ǳ����%�|y{Fx��J{�����Q7��Ը��U��bϢ��#0SKVM�iu	8݂4�qr}\���V�e�+�[�t9��V�}I�q�h�)���ic)��dս���}�NA���/�����l��Nͫ�i�A������I�� AR��ĕ�fe6f�Q�.&t�Y,�GoV}N�����ݛsL��ǲ��}r�Q�Ҭ��x)˳n�7�媙��=׽$r*�:�W׬"�=8�Pk�4Dc�Y:=�}f�ピ�R5��	�{��Pk��R�ɟE��}7�F��௸�\3)�l���Bس�Ĉ'�Ѕ�]���	�ה�Zt�*��}�
LJy��w(�JG4�M�᫆��]�����fo3nFCg`.�x��]˩�Iۋ����Y��ClH����7n��]���p��/#�M3v�h��b��9C�$�����oq6��)�;�L9{��'��ކ��=|���ƪ�<.x�Q�����@ܥϵ�B<��Z�MnУ2nl��V�~ʬ���yh�����8�3�RU�Ǹ�<�zT7�Psi[��i�����:�_Bt'2�z�
M=�qC(�ǲ�)uCJ��d.����$��mWe�YLGG%�H��֬Dw�z��px&������T�i/���q	�r������r�-��)03X�_s���8)]�b
�}R��;/�2��v
֦�ɜ����EIJ�$�T6��G��Zd�-[�5Q�����|��[_�f��E�:\z�Н���w]+��n����E�RN�%,*V��0��k�[��9��!�,�7�w�_�S�|����DU!�"�fHգ�L�x�έ'�(��g�qP�)vF�c{����c�/.��q��\7���Zʔ	������H�.R�e�Y����+�f�:l��<P�ۢ�[�{������参���}�`r>2����|�|��V[�}n��HG��/ܻ(G�2|�9��[S)_��RU�Ɔ�ۜ��n�<�bų-㧂Mf��c���6w!��]y�^�f*M�����w��f��J�m,
L�a��@���wv�pd17J���8��@ާ�j��\�ԧc�̆to;d�}��8��w�"Y;�fG�1��#�wvזl�4�\�-�;�Tw��);n�X(��s��]�X�)���5��UK2�S����P=�w�ӕ��\��;�a��Թr����9���C[@�b��oqSu�<u����=�0e͌8�Ө�=��|����3+3�37�*U�N��v��V�����w�[P���j '&���AX�G�ĺWT��j�!\�p/��ѓr�d!�zZ�5���S9ǎ��*ji�����]��m�[��JR�P�F������TKw���G���"�������$��]�}�
7�oD�(-􋷛R�gu�SQ��<VVTt��Gu�u��b�!s>� H��:�v�m��ux4��v��&��Ys��+>��E�Ⱥ�+�Ӎ2�#��*O8m�˚�N;�`�Z�c����C%;�}�!��ۆ���Hº���k ����]+r�^{0�~3±�K�e�tK(�䬥��:�T�d&_�}ޭ��1Y'65�M��M���fn�a��n웰�U�QQˠf�³����&�ƪ,{ĝ��z�Q�Ә¢��1H&wu��K����|�=�~�k��,�f&g���1��k��.�E�LG�����O�����Gm��Y�i�*>EAv�.��ɇqaChV��e�86��]iTu-�uR"�l�;��&ĳ'M�X7�G����x8�u�p7+� ��<r�=M�Y%�^`�Y�1\��]���F;�CPه\dmGք<ɭ֞�9�4�z�|H�j�����v��v�l�CA�U6���s�Z/��x�A�����;�Hth̜�	��E�ߗ�|3s��YaNZ�I9�G���{��C�ә����iV<�Z�Ж�qu������!��љ��(�H�A��f�ݙ��Z��)[}���Wʂ�"8{vlr��,�U��q�B�xZo6�������'��]�r)����<�a�¬X�clbDF�Y16]�@\՘��>ɤ�&���䫺�a�O)�6&V�q���C��c�f7A�e�ȷ+xV,���m����Ʋ*���5�*�rB�k!}]v�%鷚k!�n�ޡd�%(��UsU���-T�Z8�]Z�z^�l���L��j�$¡L��-���q3.��N4��&Q�Z���˽��I���M�����G�H칬�Vo"�����"��;/Q�+�xO"b�D�o�a�P���>ϴ9(��xl��c�������%����_���heu�q �����.�MG咴�F���#��]�·�vj�m㴫[����2t˵+��b��K����oU�yԴq�$�;�&�f���9:f�K%�zTZ�ՌF+zRC�˪�%� Ҹ^ٽC���Ikŷs�絨�ۖ�k��*)	�ʉ�l|��Kθȳ�n��Q���C�<߷q�����^ܽ3�������]U�7�ee2ɬ+�}88R�.S�EӢ����bl�[�CM5����N��t�W��Sp�?F���v�͸����=8a�19����D#.���ki�ŭPn�')�:X��|��>b���Xr�j��ڕk6s9�V�Vu�l,ʹQ���R��le��*�.޽s!*�۰.Q��<�kJ���{R/�)H����VM��gI/�i��5�Æ�qo;L��-Ǉ�W#�zoan���]�&��BV�R��ٛe�;-Lz�yW�uB�	�n�����b<�Lz�w;v�Ҵ�h�q�kd��ǿaŔ��k��?3!V����ޢg���UX�U!�۳��{�&���dY�mǺ�w �:;�ڰ�Z�T`�'m��V��������tk�W<F.�%ua��*�Fh�c;wE�}������+=L��%ܖ�m?�X'L�����{{*�I�"�{��gl�:$�<�����<�YYp�='[+��ֹ���Eփ5/r�����j�b�E���)�Bl^��'A�]��T���I�,��� ��π@�/qe�q<#҃]���]�u�V�ύ͂���r���/��E���+;��.���㚥�o(�����r�+����W���GsJ�e��4��CB�zQ��Z[�_(yra�v��O>��x5c^�g�dդW*�뷓W	�w�������ίi��A����W�/7��Ƴ]z�����u!]��4�[([�,hɹ�xk��]\�s�(��B ,�u�)U��9!�y�Y|��Js�n}��-�J�97���⮲e�:k�/oV8��77�=~Ni�=��¬�k=ɝ� ��Z���o77�'mE�B#[G�v�A���`��g5�T��G���}��7�J�*�T[�/�/E��r�{���4{�m�s����=�7.0i2b��u_[M���U�}��T��ȷ�J���vLO9�;8�3�u�T�*�4b��j�J��K,�4ꏧ A
Ov6&�"t�nu�i������L!U�e�Ҥ=�g��ݖ�]�S��M��Gd�4��n ʜ�+0�Xe�X�[mt��
�U�w�G*��J����D�Jn�<#�Z���v�m�9���Zs��W�v΢�ܹ�����(ͤO\�n�2n�;�I)�Qԉ˭�@����9����^*l�Os �Y��d]�[f����ggu��W`G-�t���z��H\�J1m[�����]�u�y��<7)u�u�Q����Q�
����Yegb��to�f�� tO&!{҂G	�=31.ӮT��l@���@������\����>Q�=ڧ����׶���v���o9T%��/�9SZ���U�U�٬l�a�.`sq��5�Ft�u˻�yV�0�/�Ae�/V8÷��Uo nr�Ҡ�m��έ�j*��,��K���z����˂�C[���l1'r���e��rx��tb����]L�p��F�Y����Y=�޹"�+�Szmm��X��+�~�I���؛�4�s8j/
�n�\�����k��y�j�e�S�C�u�I�����o̵;��/OR���WЉ
��Fuj���}Zu�ڊ�:sfk�$�hs��C���>�D*�1���Iw4��V����"v��ٴ��0Y�I�->9�)�9P�60q[����5z�F���^��,=jq�rj��|4�������A��H2��h��]K���f<�vI{#�Xt��mj��vJ��Jʊ:���Qg3��q��=��-w ��yY�Y2��*����˕�^�NPC����f�֫��'X+p���v;�}��-�MJ pj��I2Y���A,��G��4�/$��7W���:�a-_`g%�zoJ��yq��.��,ޕ8'�!��P�t4���� t��m�ɸeGX����D7�H&d7�ku�J;}6uv�tQ��G}�.GGgbU�c9|f��Jޜ�l�#�|������ � ����g#w;������z��ue�iΡ������B!!��$�o߹���9�s��|��W*��������C���Yő�ۯ2���b��M��]���=�_�\�����t�;��e��حͥ`U�HsJ5�7C���Ϻ��r%����#4��}*f<�u$�]��"���fb�Y�@]��7H�J��l�t@e���v�����6���(�OHg���q�0*��|�rZn�kj����I��tb���y�ysy�zG���J}�j22m<�&��Z��ם{nJB{)_��9B��	_-�ҭ�9�by�V�p��'X���G%���$�p5�����ǈ;�l��� �6S����d([����s�SX`�_�x�);�]���#/�W�e_5m���N�����Tra�����s�AL�خh�.&,�rn3Y;�ӧ��ڃ4"Fk�~*��]���.��Ulr�Ҡ1G�˳�Ԝ��,��ʲ��kf�\�8"����C;&L��VU�8�{��{��K�2-5�LK���i�GV9�����K�{tf[��WH|�6�_'j��ً�GQpu9fI`Ӓ�d9$��Ѡ����=�3���	�"gJ�3#:�8)9�5%�]�u,�	���o�s���2S����ٖ[��	�=��r/zgp���yDLю.��^(�|�3Y �x+K��ov	Ɵ6v>�P;�@�*�}4���&p�1���C�CN�j�O��>�)�Ž�v9�&3|��x�;���p�̇V���ɇ�N�tۯ���x"	��Zl	u�,E�h�wQ{��0؁޾;}��� -�`IYAu%��WU{9�^;9��т���k>�����algu���M��u]��ws��챃�d�b���q̜G)̍�͗�:��+dGI`��5�S�l��BOq.����'IƆ�VZ�1 oAr��#�K`����ޛ)�"���a{z��p1��7رf���б��x%Y}�w{�ժ/{�^0c�:I��\�����	rzuoi:��x˭ [��*̝7 �GT�|Ae.�߲�cs>�k�D+=�avӼ�h�]�R]6aS
�y:�׹��o�d�u��<h!X�nܛZt:,/��
O[� ����BZ�U׀,�NAq�Gne��"܆��i��a.�u˰/���A��H��.:6xZ�}b֡0f���id���LR\3��H�l�̝G:+0�}D��Q��I�C��Ͷ �j���:֖)�>�9���q]�Y=<Q�X�z�ԣȍ^��*nu���x��+�R"�Yp� l57�*�|���&�B�9
|���;�� 'ëZ�3�4躹��:���C��N�o`�wz4����ړ�H/�K��}�e"�B��mr���1}�uXՌm�H�l���"[Ij�ԙ�ͮ8��<�J�)����B4({��f�w���wF�,����%xW���[,��5�ے�k�S��v$��Gh�;x�e�)�3��%�'#.��N	ne��Y��ԑ�(a��B/��u�oG���Mn�K��r�Q�1<��>U"�"��խ+g3�ΛV>���7x{M���pѡv���F�H<�F�Q5{L���M�W��_<j���V��	Q^Ț6�3��ghV:E�Z��ǖ!5o��o�3H^�LQ{&��l{�E12�����+k�jz���1
���� �S_f�4���u���b �ޑ���8s)#�i��r�-�+Є����9u�Y�܃ߓ;Z�,�Ҙ���Z]�4��r�5_Y��t�$@�gU��qHS�
���o�a^�l6_X��>�pV�e]�U�q����v�ќ�C�=�4,�{�F�-,�y�t�w7�GZe>�� �\P꽠�Y�J�ڜ��A�\5/��`>+�A�Uas0�V�}�:n���?	J���	��,ޱL�1Y�pL�n�<��4��iG�����P��v��3�?(��#gTY=��~Cp0vܗ'���;���Á\T&��5��^����\F�k4
�"Fś(�U���H��=)�t�L��*헂��׳.��f���=��E�n�u�TOo��͏}n����O+���j�,D+�6�T��b�G\r��0�L�{�6>0�H|�p�^��Ө]+FL�t�JY8m�>�6��׃T\�|]>o��)>�9�E��DAܙ9v��JN�R1���q�L�<y}�0z͞<�wD�һ6R���ҍ�e���:��W ɽx�8h�
	����}�N�"$�;���a��Ȑ������6�SsMa4�v܃�}xKX�����6�'u�Ћ=�qݘ�	.�oT��pv���������c�l՗YR�R�g7L�N����G*��]b���3�
45��O��Ǚ#{�R\�
d1:^^�)���ɞ��'�Yӆ�K��)��r
�G8�� p��cI]ؚ���'x^.{ُq8���1��<@\H�{�F��=�zKq!�9lQ��v�ϵZ���yyh��ȷ\���*��h����#�t�9�!J`��$��:��j�U�z�%��ҙ����+�N%Y�u���_*,�#z�Lk�O.��Ϙw8 w\��M8.c� \8ٓ37�\7��|&ֶ�x՜Ef�z�je�.�HW7��<L{�*�J�����cne�&���{�H��1�d�/8*��oh�����!��}��m����1\z���;N����2�r}#���������T��k���e*l��ŵ���P:4�������2)���⽁�O�jDB���<V����E�9W�$w�Y�|Q�{p���H��4���`���o�ݤ�Q���Rda<��y�-Y�I�)3��pq�
�����z���'�2�^r����1��� ��uwg����䖌r;����Η"'���F�~�Hn�Ƭ�=�+�#o�`V(��Qٹ1H���:ڭ�]�]qv����i�ѪM��ǫk��>�掫40���X^w�ER;�hת
����-{�z�9��uy��b�;NS��� �S�p����̾x��kuQ�L�_ZR�"p��+��,[5D��w��3a�kR��'�ν��4n@f&{2E{�ߡ�+֨��ɇ�2���X��v��s�\���ߌ����UU\��j�fB�]Nm���^���ā
���/����vA���ѷ�C�q\�^�I��eg`+��s��shN�u�d_=mnc2h���y�T��]x�`4�v�WZ.��5"-�G���;3;1�*���fa���čù'��>�U 匑-e�2��@��a��G�ӣe�X�R8�}F��R�|��$�6B�ʋ͖��p.���{3�Sx� �pǋ���o2��"D��R+�P^����%	�`���z� �P���G���sl�&���A7�f��.
�<�K�Af��k��^]��j���Fc�°�vIEIh,�#���x�ՇN���|t.FKU�~�ܶ�#���G,<���Mޝ72�(H�r��YLٔ�C�]��V�db�G������T��+g��j����
���0�qp��R���	��	J��3��ԝ;��2>��,N�6�SƧ��%�X�.��x9�`�w[I^C���G��%ɳ��U�X���qϦ˘��7݌��1G����;YY���|�^���OVB��@�Y�y��:0f\��u*q{�p�GI������Rp��D�3��.�VdzQ�����GhI��!ݯ�zc��dw͹.�n��j�є���� ���	uSZ�פ�%ӳ`�fh<}��g�y���у�sÔ$9�jNV�-p�}���:	��:�bR9[��Ϧ0
��j�p�FT%����G�\�Y�u���|r�Z�"�Z��|/2̾Y��q$�!٥2QA�1>1,�`���Yc�ƭ�K���w_e�W�.�R>�BAN���X�@�Y7�ӗܥfj� ƢGvF�1b��;��N�(^��L�	��6�N|.�����wmusPp�ַx��k�)HtQ v���y�گ�'�,3�����=�X�T��%��^�E�ш_U��7����s^��7�/K��㋺__`j�d�՛��t� �δL��P�sO?����Qf���y[J�6�q/�����̣ݴ봺۔&�N�^p/O���l�:��FKn�Ǭ�ߡ�Z\(���:��V$/ºԺ{F�u��e�W/��O\��������N��,�J�\�^��*�.�!�ko�����us:1|}ݏxH��d��jJ$�$՘�P�w<�Y��˫��.)���a2��넊j�b*<捃c�C9�L�<Q�s��A<�-�0���mfw{ϳ�36a�6�ע�v�7{g)PS+�Υ��/m���!��yQM"H�����B��	^+�Q�s"fI�Q��2m��F!��]슛]MV�r�7ޙ[z���/)��nZ��{}�N?i(��a�9��:���7
���i�u�/��k
���z|��3�`'%X���m}\��<���ŗr̒��o��uvk$J���U�έٍ��f�nb�F���W��2U��oni��Y8M�-�X9DzN9Z���֫�W�)V ���C��o�0ǃ~zu4Ɯ��x+�a�2A[��DR�dךs��F�N�s.�,�����;]����YY`@�<���Fr6�J��qwosV�S��@n-�"�Tו�g�)ݦ�ǲf2���ʹ�n;>o�n��`L�Z-=�J�Pڝ
�j[{���=�OP�~�9�B;#Y�Ĳ����m�7�r�����㚄�E����/\c	��)��]G(Qþ��3�Tmr�]�d��R���"�q���MD���ەڴ�$����`���9b�MV&-v��q� �1l��3�Fk� i6��#�@����*=�� �3�]�M]����@	v�EQ	�J$�ʫ��	�;jH�=��+��Wh��av��/�����E�aNP�F�prƾѹ�v򐂖�th���Sv�m���B@ݨa�j��pt��.�ַ�����Yea @DH�R:2n����O�E�L��x�Yp��Nuu��5D���_mL46c�^ҭ�{���:���'���X�#98��!�9��7(�ul�<j���k�j��q�V��U�1��3��]q�kc��EW*�q]�L]�k	�Xk5���+�׽��x�Vj��×@
a��@��\�[1�ۨ-�v��d�.eAC�բ�mpc"h�6�A^a#s��rEۗ(XŽ�NÞU��݋T�����`ޏ��Z�=L��b�w���A�ғcCܽvǋ\}�t�5�*'�ޯt��ᣨrM�=�yX�x���_^��ul��G	C���-*��qV���8m<Tҍ�Ϸ��2����y��+��4�b��U�)ܧYu�}r;r����'p�ѣ�������	�ǩ90���8�]���b�=J�r�v:�7B�؎d8]�jY��-k�55���Q��]���FRJ���~�Y�(*o:��=�e#e^��w=D�E뻡w̛4�m��]{��ȱ�aZ[��Ys��F{y(f[�h2"�q���ɬ]���}�H���os���cWtm�R��rJ ���ݛ��`��68�zvGk�@�9�,��x��nI������8�H�Cg	�Pn�#fѥ�#z�v�C�ǩ̅��!�(u��"n�w�X���̃o)g=�u�ӗ�4�u�Nj������F�Y>
o'V��ԋȬ�V���D,���Ō���R7���5�Os^��oR�����F�r�lev�u0`���X�}a鉆2{e�-��3��9��z$F+��{0�F��iN/�����.\��������9�k1A��n����t�2�Y�Y�]B��j���/P�,����L9�;"����
j9�6� �����l77aj��z����,̝_��"X��{�}ǂ�/�v[Qc������p�R�'�Ή�Z t4�!d��w��n}�g�H����Ž1����q�7�����0�����I;��u��Z�!Sky.�Kud�i�yCnR/�Q�0#Ώ`|VQ��=i�^ˌ����9����{	��R5��;I'��,�0�n��dE��kr� �	Ջ�� eb�6Q�Q��N�u=��]EK5�g���3ݫ/��;��Kv�t�vmr���i	�5��Ӏ�pN�5�ѹG��kqx����u8���Nv4�� >��2� �2�Y����t.e�^-Y�5��.3f��ͱ��T���@Z��2��LX��;������)��v��.!���6tg#�Yj��>n�4�8V�Ëޕ�:8�5��@�#�9z��
�*Vvi=�+��Jf�%�2������J�,<.*e�=�Z�8��l�������hnu��eLp�okN�}&ԂH5zD7��{`1'O���@A�EMf�4V}}h�|��iU�uͶ	u��4%��a��eC��zqCy��ܯ56�Z1��D�@�ٓ.|���u��n����	�On�t�Ĵv6�+�3��0l��눎��v,��&T��=�s��os	���F�޸��S��mI�p+r��ؖ���wM�mR�p�W��S�Ш������yK#�m@��Wp��8���9f���u7��*㉩��s�*��E���Lʅf[��fni,R�Ѕj̂��+�$>�����`��Ð�/s^�Ǣ�Qeq�.�`�:��r��7T�����6�L=6�9Ӗ<�٘���r����\ћ�v,�N�}fqi�Uf�&��xx{�ᓋ:�	B�S�TXw����f�Y��as|��k+{�Pto��Yw9����N�ڳn�������E�<;�j��<3��i�L��z�uh�-Kh-���㻧����X,;�2��Y���#Q���9_r�-�|U�{M.��7+�K����ؓ���O)j=[i�%�F�n
�1�b�-K1h�rє�<B��-�p�=>�Y���m��7v�gf�G�Rsa���hޭw#\U�ˬ�m�1ptU�r�B�v.�_v<�#3wQ��ۯX�(=w����������8���.Sr�@N��	��\�Rpef���I�����V���gS{�2�K�S���W5�K@Rd���m�Zۮ
�wE�fr���85�W��u9�/�O�Z�������Nt��� ,5x�[����1s���,mt�]����v�2�uo#ƽ��[˗�ma�'p���l�':5{���rī��.Rm&��/y���\=�2��#!�u5l���s\�8�{Le�&l���|m��]:�D���+��Y[i�{Nb/7Rܯ\�Pe�j���d&���\�%ϻe���"�.�����n�*���s;����Y�y��6����<M48\�)	�M�N�Is��x����se�6�$����EۭM�v�M�Q6�ox�����x�v��}��m�!�J��峵"rF��AB��_�v("��VҲ�E��_�\hZCr�XVQX�(����m��j�ԣ
�DU[j9��DX�ll)lm�2V#(T��d��E��Tm���h�UF��[`��6�-���-�ej�������*.-A-KeYbQ%ETFڥ((X�ZR4��eʍ�*#VV�J؉�P�aF�֪���10q,�B�V���lU�E���\Q��*D*6�jYQ�h�Qk(�-���Zմ-,�*�n&#h�R
(֣Uj	Kb�J(5*�#mTQj4U�PU�R�e�����6��db�����5(�ũli�y���y�y�{��,8��	X����z���ՎoS��#�9��s�%�dR�3Q�%��nݲwCww�(��/+z���L%*z���~�������*فi趮���� �n.��jx��u���ߏ;��h��UN�UP�mu;�M>;��	�_H��m���1U�����L�b腼�XA���l��/s��i�p�5�:K���a�]b�[; Z�*�{X�)�=��ӓ&���&$�u��t��u����a=^<:�)}���EV+�{�b'؁2�f�*Y���q��[T"�;g��H�Xq�Z���S~�y����$G{╓{��Q�z}ƒǦ���{{4Xrhs9���*�8�7��L7�f����In�J1O���č,ǻ�vB����'R�1M���,>g*��9|k#��ȵg�|Sc9s�Z�/�U�����D��Rc4�3���^`T]*�D�o<�L*���ᜤr�Ca���}�f�t�o���So�k�*�
����#�83F�:�~�fX�(b�VrZ��)Q��T��Ǔ�v�gcΫ��Ma,u�#��>�"u�w�R-�'p�r��]vH�bJ�H��kz����k^��Lݾ�ڙ�s7Y2�%���=�bq�!�'/}�yM[����*㊄N�j�#|����F�nҚ|Ɉ滑+,Uw<��oͽ�4�(��s�Vؚ4���YO+՚��b;xOn���i�޼A���u7n��P���q*�\���fm�ɗ�۔�>���3ȩ����Y�sީ�z��FEI=ّDK�ܚ5wk�k���.��Nk5P���=�ls���T���%�ҭi�3��E���WZ�B��ƽ��ۏ;�3_�ߣ1��M_*O��a���-Y��e�M�+'�ʑ\rF'�b�xʬVp"�^r-�-q���#�54x�%�<ve�M�Y7Y�������q��Jv��cA���v�֊�M��5N�V���r�fĬ�]b[.�8^�;}��<\����r�/9�wgR8�K
�>�Z��{w��uG�{��k;�I��=7Vg�pB���u3\s�Ւ�B��k�PZ,Ij+:oY:�|��|��Q��N�fF]]7�ڶ�s
N�D��ц�.Jtz�o���+r�)lH���=`r���!�+��t�mM�Zz�M�Ւ���\��2���QKv������z�[¸ݪ�a�8��Ϫu뜗&�}����	ń�[�}Y]j��F�s�����ovfJ���f4�J��w��)�����1��)�zV9�/�$F�W$9$�S��5�,3"9+{{���}��r�8�ر. ��+�3���+�jވ{i�m�α�G)�J��Km�}����UyM�F�<�҈�s���gI���:UWʫ{z�\���6�qN���nfr}�q�W�\��SG�+Q1�lG��\�u�!��h�)�WB޼A�������\2����g#/���8%��]n���&�T>2-5�1*�Z9>O���ԡ��5�
ӹOx�{Vg�6ĭC[p;&�z���+��\+5T�� ��\�+�f�v�yTs�V��,tFRG�8ko�MqU��׷	����mM�9t5{���X총������tR�Y��cv��|RX��D�mխxq�N��I6&ŏ���+n�ɾ�҇Y�7�e��&Z�/��3a�5C���)-�����j�L�w�m4���	U�kXd$i�͗�wS�������cUs�m�Ѣ��'E��N����s�S��)3�!u�,�eH�9��������&�e=��7�;�Oі�s�Z������SvL�3Ʀ_d߄�w�+g��F���o:�T"�3��Y
�כ@�$�P�$��ST��a/�Vk/kFs�f_tp���{9eS~(v||��w�)�H����]L�����ӭ�3�[�t���K٪�^�ʴ�71�ت�^cgR�^v���7�P�Gm����Q~��x�s�y9����)�D� �'WB�l�*�a�v�K5�t��o��=���:��QY+�����_�+\cx�{�1z�õ� �Kͪ��k�g��U��gX�瓮��j_f�����n+����!Y�yM����z�n;����C-����,^�K�s���u}%�Ns|��{�U���i�`��j�"3z�V��]�̓|*���Zn���h��u��!%������۫q.U.����l;�y�O�ڜ*L��:4���R���+Ɯ��B3[]S[�s$�s�s67@�\�,�<�g��愴�f�U����&�9�� �JJ�:mg.��w.&��u�r��4#ө��Hд�r��u��lK��҄WL׳M㕢|wne�c�Ŗ5*�em��W�q�/��J]��!��5tI����*�?g�cPί7n�����]�O<�������\3��~�W�6&��F��>��{�NM���6���(WCZB������=ŋl��Nf>��`�v7#�UJ��Ľ����n�G�-na��/ewS\��u�57g�V�Qn��+�-�-W7�J�B��d�@�e�c6����	%a���ܛE��Y��;��;�)�M�*�t�g��y6�`%��̞�zћ��L_[���U�%}���9Q�}����Q̨HԝA�g'��
�zxu�r�7��Ub�y���F�Ń ��
�����O*�@�_>�Xk�����X3�C�m�C�-KUO=��09m�sw�F��oخT�D�$%ҥ�]/7��پM^b���V�S�I<z�2x�ȡWBļL��A�nl^a����'�7G̒�շ�g���*&mv��' �j������]6�)�>{Cv*m,M�=��An��о|�3&d���^lK�Y�����g���^`��K�ٯ%�&���pr�����j�Dڒ����_��~;���{��uy��{{hI���#��h�|�˪9a��~��YLP�hP�S�st56i�{��w{o]M���q�3<���[���oS�͋�؁:Я^&k��yJ���o7���I+7�r35+����򼝹�GU|iP�'S4/�5|�U�T����u�=�����Yx�Ͱ{���(�m�\\,١��\j�J���g%�t�e�܊X��oX�m���������}X9յ
��I�V��/��Y~Ħ�UzS�lr�a�ddP�og��_zcTY��͉ֈ��5�̮�_W�n�9��S������t��'*��ִ\�!�Zx�KW��H�(���
�ۍԭW9vc�iz��L6��-�q�B���f�'���gO�H����3��)���H�qTO�囡�sh˴�5�{;Q����{"�rKO�:�b�b)�fK�.w|�����s$9��b�3h׮�O����gQ�1��8���!�/t_T���r��9O}n�W��$Rg�L�ɿJ�ʚ�1<ۣ��Oy+�<��/�'�x�9��=+���0�M}67U7)�e;ͷ��Y�|�MڇLS;�%����=S%H:�KL��J~�=t�ٱ+"i�d�!�4/w���f.�#���Gw���M��w�#x�ӰU�c�S��S�Iya�M�1�J������^eU�����c��:���;��-�M=Ĺ�����5���":��w��p߳%z_{:������3M���M���7�{���{�I�psv�\����ƅ���d���y3w�oR�
�]������#�9������y:�V��j�/��H�S}x�1ڇ:��1��|����s��ꚼ�wѶ�uW�ZQsc0MTHʥ��on������ԙ��#���By~��y��S\�R���W)�qC�;�_��ʝΊ�]��uP!�-�8yt;D��v� a�b�����	HT�{��gP�;�dE;}�>ו�/����飵�N`ؓ=%�w��c�f���r�lF��$��"��R��*(����Fn�}��j�2b��Gn��\�;�N�D�c���4tZR=TB޼A��X�ul���܅���-wU��U��W�ӳ����5��3��K܊@��\�+�.��Dwb!څN�b�i�s?t�҄P�t%��k�����wxԊ�X�%&a,}|r��ô�r��<�g�T�M�T��b��Ȥ�p����N�k:-�.�M켰j�u
K���1=��S�S�'�W����+��d�egc5�":�'71����V�w�����N}�U���ЇC��p
�x��쓧 �8�4���IU�ɇg�V��y]�z�F($��g�XM�w��?`m78m����,�g#�Ȣ�ֲ"q8��B�/y��0&�:2�XD���x����C�׳ܚ�<�]a�]��*�f�6z�n+&������35Ƚg'خ��Ï����,O:��<���dHjڡ����)u#�zD���Wȍ��(-�(gf���+���p,�n�/]0ŋ�ۄ����>Uw���xA߃�TV*B�[����܂�;o'&=���ߞ�u+͡x��[$�u_0���g����N��SW��O)�@��/�b�a�{���̃���{�
3�sV��sٚ���e��oǤ���>�^�����y�uy��}}�*�͈�5���d'=��q�fB���ʴ^6;��yM����z�~ԓ�O~�2��έ�����Ď�d�D��,-�~�S
�p��l�[�]1�ӧ�\�"�����fO{U����{�m�]b��4'S9�䍧�媺a�2��	�n���D�Ե9���sd[�y)��s3�����78�$q�[K"E�|�r���\ݍc�oXΦ������&�3���.�l����Dթ��~��՚�=���+��gV;"[e-a
Ӑ��t���{��T��{b�٪��No����������O���h��Z-9��<p��\�[�^-�ߡ^׋r9j��	J�Ъ�^s~-�f-%�#f� 3sx�����X�̓${���8��R��η�2�)�+]�Èf�I��+*�.��ʇY�5w]�&���Iqa C��w���{wU�V����`�����������.$��y;�u8���*�����rZ�7{T��������vM�/-���$b�e��2�o8�,�s�]���އn5��hux�&W#�t׻UҘ��u~���{k)�/yTc�ڇ
�R[/4rBwN�XK��߽����y��J^X�M����N+SdʛȆ)����Mn�m�8��ۯ'�!Uվ������W�7�rʯ�3�|���h䇷�Iaɮ�M��&�m�9.�O'�o<kB���f����3��\�$V[���j�aҭ�^�t�v�;b4�*��m�Z��!xнK�ަ�<Ov_I���~����.�Ar\W�y�ʜڮ���5x�¯43�����n�a�g-@��5��s����ګ�	۝z:x|iP�L�$n��p;��[��os���[���m�)�AE(�l:��m��ԕ�����}������s X*n0#�l���]��8V�k�o7��9O������.���뻀[a�P�}ؓ�u��J�x_P�ni�2Y�V[*��O������+E�4i%x�jڛ-�F����i��r�<��$EX��t�{��+�+h5�ꌻ���h�\U\����qp��;�i*����$]1X(.�#Xw.dj�Ŵi�;�=ً�E�Y0c��\�w2ÄR7�F�`Ҕ3ۗ9`�}�h���,��F�;���7hMėT�cfɉFg�[�fg6��_v|�zqz��{�p��|`;(˴�a���J�Nk"i���b���P-a����6�o�"�����W,����l�I:�O]OEq�cx�%�ݤ]vr�㙫�I5Fu�vʼJ�_j7�]!�%��<��H��}�����3�
�M躌�wTy�k�c=�,+E��\O;�@^C���^oݞ�^�g����lp*rXʴ�^e
BX��&w<ͫp%j�r��!A�w���}�䠻0#�\��+;�X+��V̙[�T�Мr���2��!L3	P�\߹�J��*3��a{�TH���e3��l�K@Շ��V�<�C5᷺��oCe�t��wgV�Ƨl�6I�#��7*>CXC��0�N��䳪���c����HdUӋo]�-�f9w�.;s"Ru.��{؆��q(D�=L���!�껱z��P1cꎡm����[j�4��M<v��6��2�>�BϏZj��n�d�>�%b��N+nݷ�D�����S�כ�T��Z������GJ�Z���goJ+]�왜���L�r�+��6�!���BX"�!��'�@&�*��:�ţ��S�w,�F�I�JK�ޫ�����e���9k\�� ;��52v�8'�ͺ!�9`��w&0���l)��,��[��/��lw��{,��שӺ�KP�F����v^�ĹdR+&�Z/�W��Gh<�n)4��êӗ���Hx�љϞ�fN�O`׶��N)�/�;B��
1�Dq%�>t�͠Χ#�0��vjZ�8znd���u�JⰐ���,(6��ot���vF�s����P�_%��-��3�0v�Q֒ve����E,�WZ�}vQ���G��)W��6�s�gY�!WM�!\�f�.Y���Y�Onə�G�k�����.��=��j�ڸ����7kio��qѝ
�ӄ�І��jɃc>:7���璍�}���S2ۥ�/z�C4`�J�Ԣ��bAV>������`�x{��D��U�r�W���uԶ�q$�}�cص����S�S��WU�:2�
�m���E��jY�Ě�j�l��P����B(J��fN��6�fK�ě��M���&jh�Q^ܬ=v����tZ� ��Q�zw��dN���rAOT}]Q<gA�:.�Y�{wZ�xMkCiER�l�0r%�JZ�4j**T-���E�V�bR­�ʅKkeImEe��f.f(��iech-m�X�X����m��Qb��eJ�D�q���ȣ[Tm�@���b�%JZ��Q�`�2)R�h ��\�ŕk*Z[j�*ZX*�J�J�*�Q@Kj
�Ҩ��1�F+���ږ�V5�����[hR�+[h�(*��e��c.QB�+j�kAh��l�F�Ũ�(�4��������j ԰���kcR��`���cTC���T��J���+F���Uh�jմJ�YRƖ�kk[Z[B��Z"�eJ�ֶ�UA���meB�mQ����\�SG�*�"��j<����5�pٖ�6�L�F2̝�����[�d6�J\SP�Gpu��"�6�� �q4q��emk�Grl�xR}N�t؇��s��<ZB޼A�ޱ��4eG�+-^�o��WzP�!f{�9��#��r�Y����.��gV; �K��[x��m�ڹҥ�D՝��B����������Y��=/zꪥ�f�V<�*q���T��5��"��=f�Y5�V��_[7ůzܝ�ܴ�r�R食�{e�������c��2�<b\䬟[*��by���Ϩc�N�G�]������������bY����𪛔�����?D�}��%e�ӬV�:��mx�1A"�6�(L�<��j�+g�W��[�aU��u�툑��u!]�a�$q����6ު,���=ɤ�.��0��U�뚦�^eW�=����خX��G�e홣�}[7��s(�Q�s��^B����o)�r5�����	"e��#3�,��e�z�-V�V�bf�j�"tޱ�g,�EҥMP+3��r� z���/��h�ƌ�	��4��ȫ0:��6\\����G�1��r1���XE՚��bN����*F���]���a#�ʷ��[����3�I	e\}�Fܮ�%E^�ɘ��駹�4����*�VR/���
�v_�|��m׻%�d�o�8�m}P�����b�8jv�g}Ӱ�Urcɬ��H��M���&����p;{��W���m�h�(��'���ȍ�����c�h�|١��j❱���ov«TR�n�k�K�e�Mc�]E\X��/lM�l�$vҞz��oX�m�kP��W�k����OAO����hc��)]�W[k���c���G�OtI^XM�v���/Ӊ M��Vv:[��C�-��]=@C뢹�4mc�:#;w�дYU����NL+�+}�6�+�k�����A�ZB��qU��i����-�u�.@�)��q�!f�����>�O�xD�g�	��pA�p՗�Z�����wq;"��pLSɛ���r9j�2[ڇC��&���" ��w��T�p�+�1묉��jz�����Cjn�/M��5�	�����V�u���\$��C=w[�)c���:�o�g��C�x9ߛ�P�Z�lz�qa�>3����EN�8]5 ���qU��H��A�[r;��D��V��L{�)К-s�3{fF�ț�����Z�<d����'̞��a�!�I_P��N0=C�<�@�C��i	����T4��,���C��Xut,��d{�E���20wϯsc��������<�8��q�g��q䟝&�d8��57C�ԓ�y�z½Bh��C�1���d:�����l�AHxs�
�Y=b̾yn�{�u��5������똏d+̝9��x�>H�y%��>��E��hsXN�q'���VC�ɯ(x���O7a���M�Huf!�{gRJ���~�+�;��U\i����PR�,Y�� ���ϧ�G���V�!Xm�}�$���w��K�u��a*M�����O����f�)�u	ĞM�z���'_��q|���Gx}��~����*~�8�|.��RJ�ݟ$����9̞��'�6w��O̞C�o_2M2s��K�I����J���ù��P���z�8���X�N������\//mW���D{�6�$��t�h|�Gi��$�<��N$�+!�l�N�z����? ~Iü޾a?07;��'�$�O!�rE��`v��Πv���\jed���	���!�!�ן�<d�'��z�Y:��=��0�}N&�&����:���p��8��O��=����~w�}�'6�t���1���/���_Q�����M$9l�!�����
I��:��wa�N2u*z�|ì>N&$�0���N��}�|�Ğ��4nr����֗T������>�;W>l��!��'�v��(|�|͙��$��i$޿d8���7a�N2q*y�!�N���8�d�a�w|�	!�,}�Q����^௅�y����T�Ԟ��7�$��f��������'�n��8��>gr�$���Xm4�>|2É>e`h݇�:�������ۋ�~Dr��w�M�@,ت�*n��u�/�kf�Ἇ������c���%��B�=�=��jQs���k�ۺ՝�xv��Bv�ifu.B�uo'9��k��g|d�M�u#�U�3�5�諶:��`�4�NW�V�c��g,�t�۝�_�����ӯ�'Y<�0�O�0��V�6�������|���	�C�9�h����f�d�72�I��}�#�~�?K����-Cs1u}���݉���O�:��i�8��������I��	��l��x���p�C�>g��z���;�u
���� |G�����W�4��Y]�n���e���a�t���I'��X~d�삇>I����8���S��	�O5�?0�u	�޻�?!�6�}��q'oRb
��?j�W[׏|��s��*O�Rt��Ԝd����|��5���8����=��yl�Rm��s,06��:������&КL�����ȉrr�:�ޓ?�o�	���;7��J�$��s�*O�Y<ֲN����N�XN z�����P�%}d5�`z�׬6e������i��5���8���}�"H}� �P�C�'y�5��<��J�$�߳�+'���N�|����'=M�x��q���J�d?�d=C�������
ĜU�J�����? !�6��>A`y�d*d��w�B���G;�2N��纒�I:}dY>���wXN�|���{��ɣ�t�y��Lg��.FJ���GE����s�!��2C�k�q�T��q��,r°�M����T��k�ޏM2y�{�+�$�߲E���k � D{�G�	|9�׫�Ǐ�ٮ���,���͡8��6�i�'M����P���Ad�3���'�;�6��=eC��*M�s����&�<�=�+�	DW�(���7ھ�G������ig�}Ӑ�0��7�C���)�<B|���q?!�']��OP�?Y�)&٣��q��P��'�:���'{`~d����S���V����hEIc�C�\��ݙ�2�^������2+�֔��:�c͇.�n`x/^�#��L!f�&��JJE��v��w&X�y�ft8N�.+��V�/�*��u��m0_[4	���r�}Č���m��>��l�.�x�ɽb�����H��tO�a4��H�����w2m��ɌćOC�z�8���잡�N �{B|��|Φ2O��0��|D=.��_L�$gwF��ܰ̈a{���'g��̟�~w�{�O����M'��$X~O�̛d=C�11Y&~��N �}7d��u�=A�G�����sv1�y���_�(t�8�|��O�>v�s�������t��N�~I���7�OXNwz�HO�w�"����̛I>B����$�~���"�LY��8�}�R]��#����Rzʝ7B~I����'y�d�N�����@�O_̛��I����y�Bq!�s<�q�����H�P����"���@�&2��Q/o]<��'9-X�8�$ǧ�>d�����O�:��hn{d8��'_RN0�}�8���	���@�O_̟�`�C���ޡ:��� Ϥ�̀O���}�wo���">y������y����?'fSORm<ՇɦI�P�'�R���O�;���2q��/�䓌���R~~a7ޙ�B>��|	����}�j�k	����O?}�s<���t�	���
���C��:É?3f��=Mya�i��<2�Y>v�yhq��Oۡ��!��Ը��{���NG��Q����:~SK������yQ�0��2w����h�|�*
A�2|�d����� �N$�͘RN$�5<���'�,?$��!�X$���!�������ϛ�����߿u�٣���q>��>g�M=5�!��d��d�!�w�ԕ�G�ì+'�Y<ְ$���SsV�������3��Dz�x4~nvw,,�-���Ο��i�fY?2C�4�	��S�q�2u�Mw$:��N����T�'�w��
��VO5����2{�c	�M�;��_���?+�yr��
�u)E��e��Ռk�j�>�\p�w|B�l1����z����eu�*nZ�׹`sul�Z��毶:6�5-��1�gXu����"�Yn�.�X�q���𣫫�^��m0P�b��]�Y�n"��=�bn���E���Z��#�d����̆�N0=a���:�mߟ�x��)��T:��<;ܐ��<;�5<I:�p��RT�'_�d�� ���6L�?�7Z9=N��zϽ��ꃳT'=f٧ԓ�<a�6�2�oR�bcOl�I+��i'R>�!P�'�Xxs�B��&��z�$�IɎ|`���O��a��~�G����}�v��u���m�6j��i��<z�q��v��<d6��z�0���Ad�3���'X�<>��:�� �\�`����ڣ�i�t���N�?$�����I1��7�Wi'�NfIRm���X$��bC�����<a>I�:�٦N �m���N���A�ݞ�����Э�����_>�"�>�!��?%a�X�z��w���L���'�M'ydRm����`z��~M�Rd6��ĜA@�ݓ�:���r���*����T�=�>@��RI�<�|��VC�{�:����ӛ��?2xs���O��ߴO�I4��ȡ�8����iX~LM�Ra/��zf��R30��L]�⿨��{H�>�G��2u+<���'���4�m=�d����g:���ON�$��O�5�m���w�|�	����C�x���y��~������D��y�xq@�� Y ��5}C�'X�x���8��П$�>�����<�0�'_XM����??$���:����s��'��׿������{��.t6��|���H��x��ngp�I�?3�	���:����O�q��Y�!�N!��;��8���É??$�=�:���K�������l�/��2P~?{��>G�o(���3�Y�8��gل8�>M��4�q���4�I>}�2|�����'Y8����8���~��q'��ٺ?{xk�j�f�:����|F�ͫ>�W]R��	r�U�G�<�d#=i��V��#�U9a=��	c=�Z\�gge�ds�f���8aݬ��a6�%Y�oq���.9�d��\��a�/u-�_Èmz�����"�������R��V�/�  �C7���#�?$��l!�~d�?w �=a�x�z	�Cù��T�AI��d!�Oɼ,�䞧�|�I>J�Y>|H}hq D{�|~Ϣf>����E�¸��[l:{z�$�O5̟�~x�i��r�q�d����q�{�IPP��8�d��N�Xq�����q'��,G��}	9�/����Zs1�|{���C��<x�r���>}!:���2~C��N�s u��MÝ�@��C�{(M�Τ��%d�Z��G��3��-�g��nm|��U�>�8�a�O��?$����������̰8���:��G���f�u��wu̞�4
I��z$A����.t�c�yz��W������d�VN�k	�'=t�5a?2z�a�CHq%v��=����~�u!��4��S�$�<�<�}��	�J�~����ߞ�9SP���I���{�VVG;�IY8���5���?:M��q��h7C�ԓ�y�XW�Mn�!��C^�8�uEr���dG��t;�j������wE��3��|��,��
��O��d�H�y%��;�?d�'��<@�O_�X�^P��	Ğn��=O��2<> I��1H=��|]�����v:{����
IS�a�O�R�ORq��V;�!Xz��|�I&2l�=ԗ�$뿳	Rm��尬�x�=Y>��H���G��)Nˊ?dEc՝����~C�~I�ﴓ�:�G�q$�����N���ORu��V�0̟�<���̓L�s����I4�v������w2��3�w�y���n���*�����U���G�d|G�d�I���M��9N��&���rq'Y'=��N�~$����'�甏���-��d�z��j'��5O+�Չ���zo��,�4�4Md��j�����L|d�Z�ݸ�O[
��H�#�K�\ހ���8�D�L#�T��j����3�6FEj��Y8�Ay��-}PC^�cu�ޖ����&Wgd#�I��_f������ZIrg.�W�x�Y��t��x23d<M}CL�Ad���:��/�'�8���8�d�g���:������Hg�����߲@@G������^�3�󰞰7��'Bz�=�(~M$9l�!��x��t���q��|���J���0���${��>���lxx��1_Zӻ�|�������8�׌�>�I��??�^d&����LB~C}��(|�|͙��$��z��$��$�+�݇�8}�D~���>��ä��D�uԜ�m��O߹tt���|ÿ�2s�	�*�ě}d��rN�?!�l��N�<�y�q1	���!�<I�7�f�'��Նҏ��`�2<���	�2�Gi��L[Ҿ=�}��u�?xI��YG�}���>��o�'Y<�w���	��Ł�_̛?w�=C�y;��'Y]a�1��,?_���'�Z�q���{ӷ}���:%l����<�G�28����ǂ>�������N�q���@�<�����Ms�����o��!��&���)P��{��J���{�P��Aa�5���Ͼ�����q ��" {�|0���1$�ve��N��y-2|�o����������'���q:��nk��3i6w��I�:w�3���ϻ�����9%ABt�p�¤��'��Ĝd���XN�z�P�����,?2{��q�6�a��8���u� �i�dY�E���U$X�ݜ��מ�t�Tzh~Iٜ�@�O�y9��J�$�y�q%I�+&e��>dۧ�XN z�����O(|�������=z u!���Z���ޞy�{��}���O�:}���x���;�	�>d��QI:����J�$�~Τ��{`o�a:��'�N0�@�zn��O���>#�x��z�5���d��[�]��/;��È���1lT�$��g�=>m5Җ�qklm�n��׵>�y\���l:sU#�n��o�?n{5R��x��d�2��k���,�T���3�׫Ay��վ��i���GW�����wަӥ��^�oA�xB�yҖ�:���� I|(�0�C��^a�'Xs�
�Y=Ag���=d�;�2N��纒�I:}dYǀ��H���D{O����#}Ѫ��<Q���Wӎ�
>G��|4��'��C��C^ӈ,��{�d����:�l�w��I�N��x�i���I]�N���H�~݁ﹼ�אX���սQ�Ԧ߄��<}���>��)�>Bq'��z���	��p��*�Y%O|�̜J���2z��?2����'��=���$��^�yݚ>�o~��t��f�J��t�쒤��ù��Xm����C���z��$�݇S�2qߴ��:��u�OY���̈ z�{>�=����z�i?���3�~�������#�|7쯈���<��tO�0�Os$Rz�`y�ɶC�?&3f�$=O�i��,����d��'�8�����I�w^���|�;:5����u�]y��+�g�dA��i����I�� ~d����}�'��~މ�&������̛d=C�16j��Y&k�Y8�ɶOXq'YS�xU���N��_�[þ��q����u4�~a�s2q���{�:���'|�uԞ�Ny�z��|��4���H���`<�ē�8r��,�\޾�o�3U����6�]�{H��>̏q'YS�П$�O���I�ٓ�:��n{� u'��M��'X�~vs���]`q�����H�P��u�cRt�$����角~}�i'RO�!���X�'�:��ho�!��g���_�1��|/W�������;�z��JC���{���wR���5�/�+5P����ˤ�szl��7�~��Ca��n���.�1z'4���gn�qx��]~�I�qr~��yĐ�Vk����6��{�5xsy^(өF���G��Y�z��Z���V��l���+%Aq�/z����M �KrH��K�bv�F��������}�TR��E���4P�Ж��/k�������,��T��O�������`���'��l)艥�Mx9KHW��H�xV�2T���w\���r]�pgO]o���6�r2*�72�&�d�et�]��k���<M�}��]oc=[�T�y�b��:&�3ƾ��������a��7���Io�����6��B�E�6����+	w�h�6���֓�h�Q����ٿJ˜x/1�-���ǳ�
�+$r�AV��X#Od{�EYf����w�`��k=y�B�ح@��o�\�õ��|�fk�cY��{�v���pz��]d�yHe��2���Q[Uy�����mmf�c��w%�C3�w��ԟ�M:�:��@8Oi�]?I�u���a�x��,Ow<�W.�t��5�z�+\��}Kfuכӻq�|��h�qP-�53������'l����sY��)�4v�j''F�d�s�[���pmPRƋ����{U\� ���`�5}3G*��9�L���pRV��ؖ��N�����q5z�&�h�Vӹզ�T�^:�or�1�s�|�-�R�WL������Tƽj�Up����f���3z��l�57Z�yU��.�;.�6�u����:�k�:�8�QG��p��K@z��
�Z3��̜���L�;��J�Ű��kz����\6Q�,�#sMeVV.���C\\�dR��xL���;��i`�j���q�K����}����y��A�|�����W��W)���*לhlV���P��(�6!'���*�R-T!e��d K:f��b�kov^��P7C����TA�E�/%7��o�(l���;��a,�0;.��G@=}�����v)�B��E,���)���oy�/��ʕe�s��Z�
�F�U���RJve;ȏ�U�-�A��CO�`�Z��gq^Z��	���ۗ�z�0�s�tJwuu��'��Mw[���xL�3%�J,�l��{a`j'Hح����]i�8��|��𐑢��X��&�5yyٗ��x[�=|���kB���B�K��}\��f���Uih^�v��Q��oD�ʝ�ڃ't�s6tҦ�훅�c�����]K/�ԫ�]�W�${Jvebۻ���U��/27õ�UL����u&�oP}�J�u��N�M��)J̺���^\5�T��w9�6t�ݳ���>��"�dq賜JK�Ǯ�����2L��e)�m���akC��兑���u�i�p�l}F���b#_rc���Z�sH�Y�w�0̳5T�r�j��X<]{to���>�d�A<���Z��)���RisV��/�+l,3hUo*&�\�ŁxB����,��iX�h�����7q�wK6
G�|bA�M�L��&=_^�I�0����"��n�QK4t�J⹮��Z2)�I��.Gҝ��Ut��n7�����f^�2r�Y�)=�r��5)���^��h*�w=�8JS�/8.�+;.�DP��2C��S�+)0�Jc6|ںѶN+|��qm�����mp��Xҹo���Hh�F-m�m�ovp#|Q���D9R��u�Xk���4��x�i�J�j ��X$/��z����y9Im���v�{o���pл����Cj9������cg`w��%�̾����P��>�E�k��	���#�Ie��/7��qV�P����ʹ�>\\�\�H�Y\Y��y����QgUً6֭�,5��ZV�l�<�H�G����VW:K/�q�k�F��k��WE��u>�]R�/��ü{�iu�9N�u��q
�Sݦ=�/.L��o3S����m��N-�����Ǟk{EQ��ŕ��֠�kY[JR�[Rҋj�֕
�DPb	ceF�F�X�Q�Vڍk
��mQ��E��k-b�e�+D���0C30Q�֫iF����ce�jB�k)b�
�E�̶���mj�b�ҍ���@j)-�T-)ijYQ�!YVڪ������4iq����XZ4F#J��R*�fQJ!KR�Um��*�
�Z	Jֱ҂�Um������A�P�+J����)J�h�
�R�իKZT*�U��b�K�Z1+kQjiIe-�iZ12�-A�
���cZ��[b�h�Z��h[E��B���ҎSU�U���+k
5�JѫJ�-X��`�KF�4khZV�m��-�-A��J��j+lEE[J��kX-�m)h�AU���1E*6���[jƴEF4H Q$� �D�Ǆ,x�ڕ�N���˩d7:�� X/�(��6�[0��.Es�'�J[�p���5ۡt�!�Y��w0	�S�U}U����ߵ�'������K$��⫔������Ҝv÷:w��/M�����"�s�-�1ܦX����ܪ����9�D��W<����Od`֩�6Yݚ:�b�����o6��0A����^�}�Ҧ���U�ƽj\ERˋ�S.��(��[|X�<4��t�;�̄֌�� �X��y�mo���9�\F��!�O�wcX��K9C3}p®ʍ��t�d9�M���Y��&&��[�,�rc�.TK���E��P��K��`��Wڶ��k�ص����S6)�qm�����o}�пyGQ#�i��*��θ�1��l��p�)��v&L�Y�0zn�:.V̫9r���`���O4����_6�y[4;�g�F�/GyR�]Z�;��e���#�~.��#U�=R���.a�O�wݱp^uYI!�M��ä��haUY#��׆hTx��M_#����Z�p��>Dcy$+G��9�9��<���r��]{6`��8fk�H��FF&�f���R�j���"$oh(\e��{�#�e蕓7�\E�8!v��s�D��/�v�( *F�VV�͹��a��&����<��2���(�ԥ���_����7"6Ff\jnv* *#��N�y�QJV��uں�:Q��ɞ�=���xU���B*?��{�j��C���u�������׭C�ߜ,b��,��n���J�ݚWuOR���O�ʠ�u�>=�'9��~���05U�f���O�|�-@��K�Vn��"c{R�Wn����(64�b^ڸ��E�`=��ss]�ܥ��?g�����ղ���o>f6]�1�9����edi��p�EXܤ�u�tjy�g�f1���z�KLW�$�T���r�Yz 1�>��.���/�������w�{M{b��h2RҮ.� �.}&�^�@���<�ASe��p�-��
\�t"�'��S���Ki�h��i�^P����oS��)���6�D��^'n��]V8�A�D���A��v�_�w�F����a˥����6۶uë�yͻ����@�GQ"���@�M�$rk��W�����W!8������<t���8z��[*)Ԗ8�e��R���<���<lk�f�1YTT@u)��Wz�l+�O����r��k���	̵��c{tܫP����i�E���c�FACkk	tc"w[��1n��5�3u"�Vոhڻ����%Gb��u	�W#h��\b;ǽ{m�]��[��נcbѸ�VB�ّo<3�Q�ي�nmG�Is�wk��{��:S8�	.Y6�;?{�{�^%�1�\7�/v�>�K�X�;�A�sM@��짏�YK����۽�3�<�!�k�
|k�,R�v	��ʈf�7#C�^�J7�eKQ���(/h�w-$�âQ�����+�<��b�n���#
ȰR/-�o�[v�=���:q�S��(�,Y��&��8"�n'��C���k���~bc�]�?R���_��=:���TI=�������J/����	�I)�H�A�=��-NF��u�,kJ��<��1�e{҃�RJ�
6�>�J,I�Լ�Ln��,Q�U�*���j>+}�����[��hϊ��V���i7���A؀9U����?h9莓o��x�Ⱦs�H�����������8l����m��C�ΗC���kvG���{D����9<zU�� �W+��JӬk�8���Ź,�i���S���^7(}�2�	{\��bg���.y��tT2�Y{��27�ӻ����j*�y蝇وK�QVVl��m�M���Vn?"���6����k y�(֢qW}Ҍ�H�ݩ��Y\�8��L��`S�K�+���C!�՘́u$��8�t�w�yh%we���fhP"�滯������%��l��u��n�ٜ��7�o��I�@렵�\\5[��� ������v�;������[�F�6]=�Qgq ���ګ�6�;�Ϥ�����p޻���Z�9=���z"%�$��ً:� V�\T��X�w�W����TQ7���T!HE�={�K�z��X7˓����#��Hu�T�y����� ���Kޞb)<a������sd��uΘ�%��S��\nS^f^P�Y�e�?���K��"TX�:t��|� V��sX�"�?
�%!�T�k��3�)���A٫��~�~��K�/��ڛ+�7E�2�c��\����4�6M��mlx�lҩ��Q�?i/G�5���߶y�o:v�ձ���+idVz�6��LŘ�&����&.��_q{j6��������_�V��w�����n��C�A�,O%,T>Q�J���ģ^Q�^��o�\�o4R��p�l�ֹz��+��}���>R#�L����^g�_n��'/��`��&f'd���R�l(xkJ
aY�Fa�y��ڠ*�S��  짺��a�a��l9���V���]�r��7�>;,�{lj��Uxv��%*�9�����b<�YXՠ�x���x�vmj�r�5j����#�]��]ׂe�j�p�~��>��A�[�NQ���о���=v{2�8��,��iVvF�elv,���V������qڔ.�$�\��yQ�B�:2�n
�pл����W��B�]Bh$����T�o�J�֢X���a*�$c��&�֝���s��"&n|��c����c2��A4�g(Fc�R��;��utE��L��Ry�'��84׻C�}�aɋo��hlYۦ�������Y��%WF��@��E�b��K;��gJ.�t�5Į��/�S�¶xr��ӮL�RS)s�R:=O��������u����9CD��>�-�8��k���n����ҋ!X/��}^X�+)���KpM��69mc�S��O����n����0��D�����~9�kW*�V���D��1hˆX�Qt �cY�Ң��h�&�Q��f��ق���>O���\F�)�v�B��ъYzlfZ�G�x�vcn�h�/S6܎Q~|g�w9'/k�fʉr7���h!�-m!�39D�fVnvM5f2���]5�Wꫵ/���x3�Uͽ"����`��^��>rZ�X	f�]�M�Ǖ��]A�0ol�q]�B�g����7k�k��?�{}�AZ"qN��N�G�W^��:�e�@n�r�I��܎'Ǆ��$����W)1`xH��0���Y&]qJ��(�W�r�%��s��͝��<*WM�n������<���}��`oށ�&�B=�0Q|���r�eYϮP֟L;�-����o��@�ˋ���U�JV�g�R�h	�lF�0Q��]�j�`�9dV�,(Ή֜睉Ǘ���U;wu&��^7���r�"�}tk�5���e�R�Ԡo8o����#ղ�UTC7	�A�4�0	����T�+^x?�<�YG�����t�Yř���[͚����{J�F|'Z>��j�,.�Ќ��K�{�^��~p�����^�f�zM�,�/���|��8PU��9�qxNh��;�9�iJ׼9R;��_/n:�ú=mks�l��=]�+j���H��ڷ�c�������P��ΖZD�
��@�T`���xsm��C���Q��baС�~HU��)#n:ݎ�r�l\cY�"Ax�/F\4�2���t�gm)�6�N�@��;6*�ʾ�(���E��uG,s���F[Z�[Ѷ�5hL��K%���"�y���e���p�-���(Ы�r�3k�O��qI�9�I���!�K�S�6eF�Jy�̇
(D2����s��"��z��E�aa\��ʯyE��M�fg�����o"1�}l4kl`6�C�wGs�"�'nd%��9���
ʝv�oPgn���m�mIQ��W5$��Ŕ,�w���d���� K������~�T0ߓT�;^S+��`ҝ���OT��I�'J��|MRb�s}Ͻ�V�kC�S(כ�fԺ[�z�u�y�S/�)�Gٲ�|��.>z�Wp�C���<�\�ai�{LP��d^BQoe�P�rc�V��a�&8_S��wOlfm^c����s;�}U^8���<��C �<�p�T�m�b�>SE�ʧ�i{���ѽK�Ψm?v���Ю�.&ĩp�}B����D��'��ĸ���5�=tߵe�۾g�QU.r����( ��<l��I��j;���rP��������W�w�5Kr��9:D�v�a��~c`p�lI�g����)��]Vx/��\F�l��^�G%��S�B�Z�0;��o��ـ���m�]�Ѹ����"�u[|�Ǳ^��<7�[L�x���z��1<��$���c��.D|v�K'��N�'�$���!��\�E��G���'���y7�t=��8=%���X�P�[UY����(�^�K������%@�v�f�6��xze/[ۯk�� �nyT��o�Ʒ:;�	�,���5o����̙�!=Z]�ko���VS�cC2�'�Q���N�+����5�ǝÙ��	܌t��[+:�z9f7�Y���M�:ba�׀5C�Ef�˹�şx{�����-�c�g!r�e���k率B����{��Ӧ5I1�r�$5r���\d��J)���R�̌S�l�^V_Ñ9�`J+�-Ѭg��S��Z<��M�h�P��O�YB�d�hn�%<y�V,��jb䣛Z
hg�W���`�����rgz[�{8w]V�5���q�g[#p+�;���q�5�,S�<�z�ޙʱ!I��v���ݶ��y{��F��9�(�r�F�˧��g�[>�
����z��r�k ���2�\̐��Q��@y�������,M5��+}U�`�>v8��Nu��f�����`�\��U/'���;`G��BFCR͔R�±V�Bl�|nN)�z�r�º��bTJ�L�g����Tuu-qQrN.!����_���l�2�{%2Wh�ް�@��c\����<|*P|��M��#^S�(;.M��͊�}{�	�Դ��d���p�}r��b��.Y�_϶�&�{�(v+��z��.|��^u�F�ƔXEnآ����d=�rVNQ�f��+�E
��x�(}�S�l]{�9���A�*2�IvkY[�Y94!-r^�X�4�TGx��u�2�uu���qzΧp�c=X9��{4NQ�>�F�Z�[�xJ�!̛?}���}�gdQ�0��k�����x_�<��{�^S��81{)�c�y'~m�X��v3MM��5F�/��5Mm�)�46���٭�^����T�r���)�{�\,(�$��/�N��m�K}�ƩSHB}�|�)��έC��E������7bJD`7%O+����՜�z������%Ņv&j->���A���f�E����S���=��C��t�tCFd�I~�Pk*��VZ� ๭�k�{>����/���Uo�܎�I�~��aݭ�aX(ǳY0�ؗ�Z"�G�(��>b`�K6�H�͚dez��R
}OgVڥ�=΍YH譍$c�fw8��,�9p���	�������Dor�\R�[�������ʢ�}w��BH��/�%��p�ͽ/�׌�5*�72ꩼWϚz�e݊�0�9ID�Y���,�YUr�cS�чJq��0�W�D�mԫ�l��{�P-�S�!.xV���[��z�D�R%=\EWMu8�TYG����0���j�u�Ɩ�{`�ͱC�Kلj7Ý+��7�1�Y�����5�in�SG\
�S��>7K�g*��Z��e>騱��J�s�j-;�L2��u�7[\�ށ�㔯7ch.� �L���ka\O2���cN�G��ӣH�B�Rπ���/{���@���~�;��̂�p���3����������;X����=\k�U�[�"a"�&�r�㑪�zĽ���Y�W�Sj-���|�M7Nۮ�Q�:,U������u�9۔jp�1��5}�ͧ#�X|g�n�O�?L�A�r>��CNd��OK��"UT'���]e8;q�B�F}�P���p�soH�+O5�,�>��@����^�����<����'�z͈7�#�\d:5䒏^�Z�޶o��M�9qa<I�>���ڽ�KQac�Ɓ�%��?���� �P��΁=kb0�E���#�`���W,˳�U���S�3��Ps�A�"�,y�cI��%/(1��_b�`vhaU�b>�B�[�!!^�UV�K��.�VtǦ�H��ub��0^�0�#�y���p�^�O,Q>�Q��%缞5� ���/U[��]	fPr�"�Ϭ���]E�;Gr������j5�m	���s�~�����u�W��9|IY)Q@f��8��揍��х����H�߾������%vַn���T�\�b�l̬K�FG3I�m�r����p��fmF(�j���ܡ��_U.X ��SF�5�[x���'+6)��fL�鳱��|�5+'���'�W����p����ߛ0��c��"�!ǅqc�k2.�n�v��`Ŕ�sŮ����]"���|#2���]�3����2w2Mڋ�ll��W��[�Y�����=j�
$LT�v��`ȭG+Df�5�r;�m)NY�֙j�=�8yϩ��o�LI��ir>w�{�h��f��b�&�c�e*
��O���wx��,V�s�a䌃)܁^�&]\^j�y�ir�: �yz+	C�VR�0��Ɔ��ux:�̺Es�U���ud�ɉ$p�V�y��SQO���Of^u�p�nó� ���	��sVK�UL�� EG�e6��_�K8\��]<��x�;�����a���7Bc�2�t�ǃ�����B���|8�*x�����>�%n�A<��8dUr+X燻�g:H�^V���%"�
����	��ž�V�f_Z�]X��ܽ�ӧWc�+���/*3.�s��a�ϻ5���������R9,�!���6eA�9h3�,�4�stm���0N��#͓�C����m#{.�M;���/����
�X� r# �ڎm;����-��)(
���*�b&�f9J]Ŵ���Q��zf�r���������{30�c�r�YFo�>�){��=`̙�GE�q�$#�_K������ONSs�7��(Һ3d�a��ܓ�P�nV�|��Yd�y�3��7J���B��1��W��֑���8Ө6N����$䧺yF/$��XQ���o�)����\�9��Z3�ȽX��(��e>Y�)Gr�eY*���ժ�7�Ά�R�֎��[7��J'&J���_,I�Νa��XA&p���𭃪�H��]q}aR�(:}�V���, �w�`�+~�>�-���F��í���{��L�d�n�@V������*�=�6:��yǣO�ws�I�<8�{����Hvj[�O����I��Z����\/����6C���;��7�� ��ٗ�(�'W �u��Q�ž�u�ݜh<,�\��ٲ��6Jޮ��P�˪�(�1K\�R��9(��輰���-�ľ�7��`z�6*�"[}�C���]�K�֪�����
�o'+�Z�˝��D����������`�%M��h�ɩ�0>�:�Ϣ���#�Y;Q�[�;�u"��K[]Wɭ&asu�;���Vka����N&��]w�o>�6�A�-i�fo�c_��t"i�wa��%<�қ�`��\a�n�/U���8�IΧ8�%�/k{mu�r0$������݋�U�\��wސ/WWCN^I�T�t�ee��c�̆�%P�6���u�����?O��--E���Q+Kh%�R��[LLDq)R���Kh֤iT)j��.ث+Z��b�[l�1���QE�Т�ڌUF��+l*"�j�����Ҵhʬm*��TP+J�*��cZ4�#F��m*X��VQV[YiUeJ���E��V9��J6��m
��Kj����h�*�c�b��V�,m�҃+Y*���e+IY�J-�ҵ��FUP��Ԭ����-E��(�������U�\�TjTDm�EKK�Kk+YH�ZDUAk(�ZX���J,*4R��*F��"�����PQ�-��Tm[IY[h��mUjJ�b""�b�l�
�Ь*�ڵ��ƍ�dE���XRʊ�����A-�(�ƪ*���X�JU��ȱb(*�[iim.!�b�)l-��V�UH6ʖ�-���֠��
���[m�D` ְZ���F�+�Z�+TQ,�V�3*���U�VҦ2\�b�%���l̸�e�5W4�r��F'���кѷQn�V���F��/K�N��re�YF3(丨��r���6�h�H�u�Ι���� �W4���6��t�*�~�&/e�|�Ez

��ğuz-K =��5�٧�;��9�QY���|`����|t}�����:���LN�Z"�	�Zi��G���o8�Q���;}��C�.���]1F��:E�0�تG/��@͖�߶Qt�Q�:l�x�+���`��T�x��t���݁=��s�l�:�ŏ�&�
�������x�ݮJ��>����y.�M�T0���j)���0in����i=S�*h",MR�oc���0�I�)����y���	��
�E�O��VGb}�m�:��������x�AY����񞒳1s'�ୌ<���L�1^#�,�	'=P�(w����1�+�1��/l3���I��3	{����<�"����\$9�K�/�q�.���O�{P�"y�9�\ޫ8Cy�~�3ZA:�z�:lU�g�?���oer\�\;�*Xu֣�Ui�]Zג�5g��e��ڛB��fW�6�uM����e`�x�E$g�5Ե�D��
!�ӻǵ��U���q���-Î��Z�G�D9�y��Z%��eleomd=Wv�c37��Y�2}2�P��oA�*��^�*�
�Li��#{�����Ӣ��r6Y��\]ʢ�{ѻ2H{{�a�Ǐ:��Ea2h.ƍOE�s�]/1 ��l�Í�,t�<g磌ﾪ�2���G��X��Axht;b���ڗ`p��)tGA���)��^x/X��~�n�a�,�1�����s��w��Ob�`�0쫲a�a�o�����S^��>'ϙo�q�W��(Ӽ�5�R6fhs�2�Ħh��7�N�-vZJi�+��	#���{�Owr��\HÇǚ�Zr ߘ������[UN�Ԩ��:����7^��A���TO$S��7M��\#!?;3㸖.`�'د�/�/�PZx� ����Z��;� *d�7jչ�pI������u�:�X��yY|��+�a���ő���s��S�=0}�������%9�ٵ�
[�������ł����b�7E�4,�'�7����ޡͰ�rKN'���y��Wm"7cEF����a�t2�+�27=�u�v1��6�(�Od�p�L�e��Cf����u����h4.1È�(�ʩ.�� �{q��Wxl'��W����畽��A�{:2�Vqk(��I��)��;�����y�K;юӽ&�:
�A�R"�%�[��rw5h�t��b8�ٍ0憺�R�7M곬�y��.\�g���6n4u߱�n�����w��j3ђ�X�/��o;������B6�$��9������,�$��i��q��E��Ȼ"�\]��������D�`�c��5Y1� �)sL�
�%\5tb��0���QoHUZu5���s٢��@"�)|��W�VY��2B�)`�k��/(K�<����ڌZ�<�������%Y��������Ӯ	��y���D%�D�����k�a��Qd7��jy�s��kt�1��՛(�-V�e:��C$�~aw9��&٥S��2�� �7��Fw�.��̊�U}�
*��Cf�f�+idV
T�a�x).�>��:;Q��}%��l�����*#�Pb�Ѡ�\�l��e�Nz\�� �3\�+�0S��,V)��i;t��n��P�3�U�j$�t$B_���ᎋ9կ/P���Jj���7IH�m��C��3ݏv�Q��u�Ǝ�Iq<٣���)U���f�j)��؞��E�өx��T R�X̢M��Չ�e�B`<+�1,��T,ݡ}x�ʷ}�`gF��⽰���W�p0^%D�/b,5PD㽱&�֝���&3��AW�&���#!�bNT�'`l�4g�=��a�Av�5���_���^��x���[�?zR�Y�E�غ������,aҰ��v.�z�]Ƭ�/	\�,ǹ�8��uӄє���w���uwTr��Ɔɘ՝�vtй�bk �&[�|��}�W��8X�z�\m�K���b�F(�X6gqS�[��� �i�O�����ۓV��6t;g�jm����b�9�S�\rߛ�߲4�+�"�V����DPX���г��Z/6�!d .���:QB��W�C����\W��Z< xxG]�/�}.��[V>��l⻜��B(��X�D�V��fIo�C>W�`m��e��N-��^�]X�����R�X�%�
���ԫz�m��E�M����3�J'SRt8m��\>:g��̍mƨ7�ە��YP1��G�/zy�:ߦ�4ڋ@�2���9�������{3FRV�,��E�Vw�z;���E�m"��S���<����/�.Q.GJ����m��:�?+��m͓F��ǆ��W�b%ڦ,ҡ��X���T����j��h�+�0��/Rާ��J���Q�$p����zhKC�*�K���q��\5�Vw�NG\=C)I�6'n�)2�ء�١~��O7��>��Γ�(A��s�ߋ��ӑ��v\�˜�H�[3���Yy��Fj^�`������iW���z��޽�aMhw�Dl�������o�3�ּTp4�W�z���4���b�pnk8��_*�uo��o2�
\��`ƙ�{P��B�gN��HX���'��v/'������|�1B&��)dW�P���kj���m�85�~���C
ȳ/�l�b�^aL��$�EpG�4���܄v��Ѕd�|̬������>7����(F�O=�ɯ%r~ǣt��?(x�Dk��	�=j5fQhFv��1.��mI~wVjx�q3���׻0�⏁�[g��׾�(*�68�C��揍���b,#��	γ؟75���UT���&
͜�B9W�ü�ۖli�H�m_���[���	�@�;/�2���E-�D��P����Ζ<>�;Q�w*���.�hp�����u���J��������z�'��s;��k���k�Y}�^"��a�Uqx���_�����ǹ�᷺Ʃ�4+���T���S�a��j����\�C�g>v�
���@�ژ#n�&��ک�ct�1�.���lt�SR�5y�2��6�<5�&�5��\*��kͤ�.a���j���CtlE�p㲑f��S6<�����+���襺�e8���w�a2���*1o�ԙ�i>��T�=b�t��Qʹ���*��s�ﬅ�Mڙ+^��o,��.�5OԻb�:�anb�$o]gS�����'�k����fR�.=��O1y�
ȁ���n�(��ɮs5e�e꨻��m�So����W��{��k���ݜ���iq�9)�`l]���Nz���g�OAXv��=䃜��W�{:�V�N�̧�GF�傪��/��:��Qw�}W��q��`�V�^�է���)�@!oN��UPn\BL�H�u�V�>'�1�.���O7���6�2��7��Sb*�KR�X)W,���yP�Y�>'���K�]�O��[�w��⣡*��yyӻ��6��&�a�8໪R�0e>��)�U0�߀�!���+s���vC���W�N�6"��jQ�o8�,g��z�]����N�z��T�ת�����-�;Z�3�]e��^(y:�*ԓ�>��(JaƋ:'M8��u���Jx�Ə��w�L�J�ϨvDp��`��Ԙ�|���.I:�R��:��ŉG��U����N�*�Ǧܢ�PdD�7f��L�?v������ڷÁ�ސ~]�^��@�)�?�s|fj� �Z�"2��w%�G�kĞk���_�E2����!���z��8�hCu��!�HnV�|1�=�r�uGT�.��W�o����8�_��-�4hu��3-�P��@�a<��>��>u��KyO�s����*����Q�Ӭ���V��wt�P2��H�B����Z���ta�rk�ܓ��������m��Y��P�b������� �x��r��OQ��&��R�6ݡ��=|�`Cݜ]>��cyPf�V�p}��i�݆s�Ěu��vh/�b�+�<U�Q��q*dj�Ù����j(W=��u�
>�J�w��Ja	�z�ҥOUz�dQ0+��Cz��D\a�d��q��\[}��͛�o���z�������)̲k�{P�Ξ��`�����j��<�nxz�Fe��י����㧎=��ST�0�aՕ����]���(
�FB*�턎j�29���gg)䝱Y͒���!��/zpr6]y��u�L�8�w�Pe��`�����r���~P�7���W�iuu2�����M��I޿k̀E8d e�u��VW3�/�
�͋����g�4�U��2x��g�Y����l�z�r��d�mђoֺ��A�Eor,!��;iROu�]bE�o�������,��ԭ��X)Sq����f	�����j�}w{:@U*~Z���#)2<r��aP��٠6{Ӓ�gY�f�HWK����CRĵ(�NAo��	�b���=y=.�	�M��������!���S~L�;�@��~w0V/�<��1����wLB��q]K�	Oax�EV:R��m�U�!V���i3�7�7R���*�ov���1a��X)㘶����}	��/W�_}��r���z����$��F�����"`�,`��ˍ�^�;.x�����
��λ��7gY�5{0~�}?l[��`+j"(B�мxk������
�>Y��Vo�T���-KR1��ć���;ރ �v^I���4&�»Y�9�p��B=+N���w;��S�\b�Gb��5������0���5PD�w�$��(4b/ey��Y�o�,��k��k�>���;[���e�(g!������w�H!���[�yw�,�{��C��TR�٘)t�g/j�:24�*�U���7Yg!�̋�t�L��f�#&�*���ۙyS�ih�g*�+؇;��Xׂq?u� �N��;}y%��2���LL:�\?n*��������<_xV�����U�Xڑ�uH�z�������߰lb�{�1�-�֩��6Y�Uv��6����Gz�N��������lߦ/J]�yur�7H���yL�r4�C�m��5	{��eC�[BW��}�\F�)����O�f�����j��孺�W�ۋnm���9����ru�Ҳ5�x��`o���79k�/����ޕ۹]��t����F���>FjI�w-��oB_f��;�V']�����r#N��PF�4+-�·/�hHvbʃT�sV�=��n�3xx &�Rq0Յ�+��؊嗹��5}�̈́�r���͖O�?L�X*%�פ�R�5�y�/��N�sO���Ö�b��&]�b�k�ozY�}\D�n���X�Q�GPy�;n�NޑZ����.���t��I�U�bd�٫���~O˞M�c�c{;#S�O6��
���u7����dBm�87)R��V�Γ�>{5_���o%s�����Ѻ~P�u��(F�,X�&4����$�~pk�o�^-&f��U���r�vi[nc��L�N�~�֌�	��pO�]EPk���`:u��sKG����49��N�*��{�:���)�'�ӆg*K�k���S�Τs�5f��m�s���5��t�����N��o��^Q���~|^/y�E�I�Anlp�C���a���N�{{k@���"ĩ�^f��&��H�z�Z���ѕ�:��i�J�Ԩ�ۗ�n�[����RY����%Su���'8�<=�{=lN�p�0}�]y�w�/S~�Z"�`���B�	W+�>w�1�G�'b��߾�W�\�A�aM�����,�#�'�p�f�Q0�0>�7[G����rkY�wC�6b%u��Ɠɚ��^�\T�WWt� ��I������%�hQ�]��NrZ9s��}���)K&h5!뾉��� t��T��
�F���2��K��ݯ�b�������i�2����e�5�p̹|�f;{�X�U5�_�U��-�`=T���i�O,i`��N��z��S���mʸ�6J�֘���uӀ��Qq���)u�K���T�9ܳڝ�6x��'�wb3�q3���[���^�6V
*�xf�c�����'���K�����6۶u�y�S%tt�H�շ<�A{S�;>޾/�Iq�]Qb���#b�Or�=p�P�&=i����wS�٪�UQ����y�H�9�r_�2���r�J��du��
y���͠�4e�"������.;EeoM<����tdmbJ�p/�\;�*Z���.`C��_z�z�A<�P�O#�]jh�)@E���T��r�q��C%���7�9u9n
��%aE�$�g'�ZKM]����;���f��Px16+��ڗ`p���>��*aleb΅��7.����j��Q�/�6+\��K4wMJ4��e��:�%��,5=�-v��8�n��R���Q̂���e���ݓ��z��5��lthΘ�b>����ZW�x��g��Ήc����t۹ׇ���	���Ն0a�Qc뷢��K��ڕ�2!�;
�a���4�9N��`�0RY �m;��c�j�m9�颮�Q��w��|(��#��L6��a��䲲���b�b��2O:��7�qU��D	+7Ԫs"�ʍ�z�s�Էx�����t�w�O�fn��mހmj�����d��ّ��F��(%Xi�y	�Q�LVR�<���̀��ΐ%�������}�o�|#�~�Lv����0��	�fadJ�1�t��i�����wvh�`귗��1���uҲq���맵ppd�����a���l��z-�����=9�.(�a�݁�N�6_S�����8t�/T/p��V^�Wg�)ਞ�1��wHD<p��u��!]�$�2�oϏ�ȅ�����I���`��8R֩����%��v̤A�Y[�Bf�]�rh,@/�u��b�iwF Y���vk�Y�v��=6-F���WB��=����N�n[&D5�(h��i�pM��Nb�8|��(o�]3��$��zf<�ݡ������oT'���=�&7V�U�M�R��5Q���Zc{Q��lFgm��*�j�X�@bI���0v����Wzvi���4�@�Qit��o�#��x�>����m��t,{L*s7x+=a�>�T�Q�����ҳ!�Z.��	ד��{dgdKg-j�V_
G�3Ds�����uo�0�s�$�]�*=�;!젴�)Z\p���N�@�
9�n�B^^95�p��bԫ^k9�r�C9��ڲ�N��B�V3�7r����� �^�K0�:��\�m���u��5r曵1<uvS�g���T����1*a���Vj6�b�\o�}�/�b\m5�_l���f0Ɋ��9.�zܦ�m�8V*�*����v���|ل:/�}�'�����ܥ1ðU�y*��j7���nf�i� 偾�l��tR��L[��؝�� HVc��%�]O�h�VRpU�I���	G��]��,B�u�)R�R�[zE$U�p�F���A�-� 8�������&�X���R#{'r���O|緟�xJ1W�@��~��m����v�C�U^�űѥ4T/��ڷ�Q��\�
�W�D�➸�4- 
�܇.��̄��]]��G;�#PX��;^Z�P�f��R�Slk.�T�B�����]2�i�!^Q癠�H�T�NE���
�G
�묕:s��w��gAR�axF{��j�N'$��gǸ�°��30�w/�)Ɇ�M	oG\(�{y}wK��ڏ$�W-���ג�(d�x��:uCL������l8v��19�27�yfwN���R�������h��n�Ѿ��jة��z����x�3���>��E����[m��,mTU��-�cl�(*�"�R�-m�VեYm��TX��(����T�f�Q�m�Jڕ�ʊE*���QPF01FTTH[V�؃+eJ���EL��Qb�ĢAAE�&[2��EQ`��ڋ
6�JU�j�Z%��U!m���Z�5h�T`�0U��DE�Tq�1j���m�mh[eY�*�A@S)TR
�����"�P���b�E��D��b��TEUKj!R�(�*VXed�-�+DU�P���\�*��`�#mUDX���PưQ�֊�Qm�DR��"e�LJ���-�X�4dY�*ʋQZ�$R�U��!m-rZE+U0`���b�4�AEU�c���m�
�UE!Y-�E�DeJȵ*��Lj�����1�E��kJ�J�mQIV��\�TR�����V-ˈ�4`��\�LAdKJ�)m*Ub�����V*�b�CT��YZ�k3.%`�EE�+�(V�UF#��U��I*QE ��++��TY��@�_ ʹ��R3��X�ٓ5I�5j��R�Qӏ�VSA'ώf�����6��q�Ƚ�y����u��^U|����%�jqg�=�����M��3d,��S��NTq����2\t�935�k�c��/��ڞ@`/;/7�}�nM^�E�3ܴ�3(�����.9�����r1���1��X�Nۍ�f�M���j�j����rcvX=�b��0���3�VW�j�7���������Y�aj����r�d��H�)���051�����{q�D oc\�Æ
:���*?&W�˳�yƦ?M���F��8hv�pm��݆�N뾱%��ű%�m2���=c��-��KX�(˹�>kj�#!��oK��`t2�)�F�֝������X��VO�>�Tܸ�}���n��Qx��"Iѥ�<�(q`O�D�F����c�Y�ǖϷj�up���k��[�*SZ[��gpM�ɗ���)̲oT$�kOqO#�P+`*
������7{�ں\�&nG:4�Ï��#AMR�Þl:��O���v���^���dU0�'w_g�cy\��	 �ŊV9�nF16{�č�^v<!5	��H<.S^f�yB|8{�-�ߋ���7��������9һn��C2=��Ju��q^�|�n�Q��{ ��v�O�0�ȷs�Գo8�L��ew[�|�(���,Ń����x��C�9M���#�Ե{�"�5+���6��AtLYi^���ƾ���aoW�UUQ^�w�9˔j���%�W����,X<�o\��z� A�!]2�nH��**�,��=M�l�i;��q)E������L�Ef�6)j�k)�(��2J3n�a��$�%�/IUoږ��Lq�ϐ���禄��<�R���U}B���+��aQ��H���f��{wۓ�����'���X�����U2�OL�GƯ�7��*�}P�f��.�^�g])�9��EXz�ظXS-%�E����Pc�����꫇�������՗ҝ��Xf�Cu��¡��`�r��-�&���k�v&E�����j�q`��V!���6�����Φ�G^*��N�\I�H�L�&�k <�BVE�2�n
�p䗹��e��̇k���f�^��ŝ+bk�eG�FK��$�Z"����;��L�)��6���hC"Y�(�3�a��^�����!��b/ `,��uğ{i��t4�}dڬ[��s<�&-D��lW^H��Xφ^���EJx��u�n��C	s#��'�?��s�כ��E	�qw�+2�4��X�P���)P�;n[�����Vwr�oV�z+���W{3�$�av\iL~ˮwvD��Xk%M��T}uy�&�:�bК�A����4��r|������vfu�����:<��i2�IlUԫU� �v��%K��?x��u�UħS���x�k�8����x �:�^S�yXt�x➡絻�]@�ڿ}��.(�}dALu���[�y����jDKΩ
[�os�&ox��Q�!����odkR��QG1�̂�p�U��3֢u7)����n�q[N��L������"�(��e"�)Q�[\{P��<�lM\h)���38T��&ٵ�A�����::,R�ꫪ
6\F�^��,ׯ�����Qo��\_Oh��-�1f:��,�ه�&u�Z�� �Xx��兴��u�&�SzT6��w6􊒴�X=����ґ3ܞ����*�3n`mT($�VFȄEq���5䒏^Ή�]�l�D�t��b8c�=�r��J�&��!\XOc��>��$�����(T>hԼ�p�y[�^R�^P��[�~:/A0c�({�@p\�E�,X�&4�����7�7����5�b�`Azn�S]|�?t��8�>�������.��%@G4UD"U�#�il`R�u*��h�_��M_y]�.�{�y2����X��b�(�XP�e�V!�{��Ha���3���+3Gl�]������gm�}��Qջf�/Dh��0pG��ޗ�]x���"��ΙFL���RRw4���S���_e*imd(�Fmm�R����Y[�{�{'6��on1�x��$S�a.��t:̠��E�:����]E��M��g�t��U�o�f�a[,uK/ztT3���,b��1��IP�l����sG�؁��Ϻ��ܨ�[����/ޣ<��<�T���*GsՀZ���b?���P# Ao�8�TWԕ��ǶHVҪza>��:��b��Ζ<>�;U�q�x^��c���DG�]���o��úy�
DS�Iq��w����WӠ���e��V���!d���4��vҸ����>��d�����c�^��F��=�a��;��x�`	�#��p���=?��0�EP,��5���Ϟ*�+�:��ˋ�Eה��lt�l&��v��{r<��#�c�΁7U�mp�w�����cL���[V!�Wފ%gyrsŞ[(�)�B=x�vθ����U��r��0��ۓ��mF3��#s�Ҭ�v&1w+�9��yP���]��w��rj@��OAXvGp��qу�rʪ���g�Pօ��y8B*�c�Ɠ�]��0gq�b��n�J��=Ŷ��cAP��q
S�x6�y�P�:	���Vq��l��[��+X}�R�`��Y���H�Y���d4v2�q�>R���(�pE ������1��f)�9��y�E`�����߾�ꯩ>7��Qb*�N�wM�������P�F�7%D�R����:�Q��!���T<#��[��g�l�U�8*�UFlkԵ<.y\��
�CH��tE�ԵǮ�hcdb�}��M<��}�t&��G�x�/o�<��n8.Ի���)�\�h�>ts����W-��c�u�.�<	ӻ�C	BϘ덏lV���e]�}���w���s���V8�F��Օ�:��,�W���C�\~���V{7�Il߱�8��=�`�}�v�7�n� �7��+ks��%�ⱿenzfkX��Y�4�-�gF�j��}:±��)jĻ��#��Ǳ,Q��O����@�����7]�j�D�'�"�J��0���+�,�q�jc��3X�2�+>��+Q�8]./M������MY��r�/�&���4;[�6�hn�y���9��&�oE����:٘�����#�*��R���.�/�2(/�=�Rg5C��p�g]i݌�q��^EnD�
Gpɐ��R�����e�ޖ�^��t {R��U��'.���̏2�Q-�J�V�6���Q�K�E˱Hks���7��\��6]Nݒ��`C]!��5r�q�(\΍�v�!�����Ù�^vLus�E�Ԛɞ��A%+j�}� 
�%���QBѺ�9������|�*|�Puq�G�F�F�˧��p�=���x�Y7z%�}кԐR>�6��n��y�L��e�LL�h^�$����űY�!أH7W{A �8�x�/(UWt1�%�����
�#AMR�À6YY.i�ʺ%P�j ��,��l�S�j䱒�Z�5c�+zGb��9��:���Be�C��*G����7�~���r��Co-uj؇�(����t�,�M�w���#@p�@�2�oER���U^$:�3���F�'��X�(�g���ͤlR�l�S�Q��d�U���DRz[=/n�ΐ��� i�=�	��Bx�<��J㛊��{��S\�����㹰u�{�I]�G�:�p�+�|y�M�kR]�#)?��/�T�\u=0{yb��߄�$�rF��9Hs�.�5hS\+hv-��)��c�H�[~|)]%2��㪶�"���͂�Zj�vd>|$� pGÉ��D`7%O&%���{֒��\�Qx�uR"��#�\35��g��n�����C%��֒��������o�������|�
s�P�G�<$E���H�G�7�	
p���9��E	Wxv���}Z:�-�ƩS����A�]u��4�I��;�t/wdq�C�����y��MSǝ�b��� *�n���������_�E=\
�O�]�Q&��8���eF@aWG6�P+�Z���N����:v��V4<w{�F��2_,3�?�Z"�G�(�;Ś�q5☴�K+��wv�Z���2��ɦFW�nѱ�2���X6gۊ�E��g�<:Aȧ{�v�;�x�]8 �4c�k�o��m?�R>ݪ0�˸�^#���+����\�Nt����$�y��3*����QM��35�.�k��0_�=������G�	/`�^M�����uO9�I~���)��;KF��68V��K���c��n���S�^�kqəͽW���0�bO-m}���j�)Y��+�DZ�Qzp8�3�J'S|��[[Ĕ�oLk�u��-t�EgK./)�^R4�ж���e�u�mo��|��=՞�R3�"M���U�4����j��'n�s���Y����5}�ͧ#�X|g�w9'_��V�Ffn�ܞ��:6�x'�B� +KŴ�ة{��ڦ,�ҡ~ڇ~���Plz�՛W�lI�o�����Jɗ���2͊7���Kl4�I��v͞���98j�y�Ft��7���F9}�$icެ�;'U�:K����̄M�x8���U<��*�sٔ�x��n��a��'FAt6��Y�|��\,�*Y���\�F�p�D�G��+ܟ�Zܖ�����<F^�aLL�;5e#�̸�l���Ffo�z&֚��uf_P֘��?O4����R�6�/v��kI�inN^ҽ���3$��0�sՖ��&׶�)��PB�B�Cs�1�����&.���໇���a��4��F?x��[������k�5� U��_�A��lT	�^|�-�3�	7���m>f��]]��C��i"���N���]���$e��o��Qfg�	Ր���Zw�w�=38T`�+&�K+zv����p��{ΞJ�%_g

�lpb��hn�u� %�}w?!CH�2�C�pR���,D�}[|��^V��O��5�4�Yٸ��r���z�x�*�D01Ψ��[kϳ����j6*�!�f�s�kPc��ؘt(C��ES�k��|_>��6��^��M�=���Ce_N��=1G�Z'H�q�f�*�͔����y�n�5�]��\t�)��6Qu��s�� �S�y<{�'�8�E�c�r�!ެ�۳�������y�����hm�"oPD��t�[ܫ��'���&�[��.��+�y����:�Ʀ�f(7Vr��_z�$jx��T�	������h��;>���N�_7)��\��nI�/7�������]�D_y,f4�R
]s'�?��i��f^]�ޑ`��LΖ\^�.�R����aMK��r�k���j���Pal�;�1�}�h.�1�ZO]k*�� ���_�zo{����4��xX�I診����k�\1��ͩ�rw������o搮&p9�»�a��!w�~�F��*�"�|�`��TqC�Y��VbLp��3��䒅�_]�Ms5�.�*Y�yخ�����۩^�p�7Z�']K��dr�@k��U �#�^R����*���ř����-�<��Zs1*�#�\�Èe��62�;��NU��M$k�/Υ��vkt���+��:u�Ҙs��F�h�׶"Q��,�^j�5b�#v%]�� �j׮�>�rڻ�f�P(������C���� ^�:w�F�|,2789���~�[w��pno(/�z��=���u����c0k�۩�Ǘ}�U�'�_mrR��y�q��F��4q�a�+�{�Cl�Y��>���(���EmnpzK5Ɩ7��?d���oVz�\j��g�Ū�+=�ڡ�b|ƿ,W��|�2�T�j.�=��X���Y�7t�:�����E;B��%�)#�H� d	�L�R�J�n����B�Wl���|t�������ν*q�R[l'�h�������&����.�����
� �7����}����3ݹ#f���Υ�s�yX����G�rp�a}yj����J����J֗����5��� S��)�jcc]�	���lQ�lPrgv������.�_�mN�_zT|ovh�8l�U�Q8k���ov��7w�<X$���R��B$�i���Y�͎��TyK���u1W�����2.2���KX\�]�yv�S\u���n}����Eg��P����t�!��|�o$��ʐ4.1C��r�������>��g���w��b`F�U��h�\�Y��ܞ��Cb����O���<$x��w��zu�lHyԝ{[.�"�*�Nۆt���SZ
h�4�e]�H���e�G�Ǚ���t�N��T��¸���^!/zs����Yf�Ȅ���z�<ǱE���=�^���e�ODP呖2QU��ҍ�|�`,]65�;��y���ѵm�]#9D��n�]^�i��|�V���|e�Ô{0m3�͔tR�l�z�r��d�_Ԫ�����/���\@�[q�{�Ѽ�@��Y�Yx��'�67�7�f;��g�=���bf���n�D�q���ᜊ�Ks.<��j�f��j=Jd�,��h;BA�üV����ꝔK{��ٟfbF�ǘ.C��.�wf3ݽ�Q�f�!�)�'�&0h޲��/��H�g�ޤyظ,�ƚU�έ��.h�A�ia|M��m�i*���;�[�]G)�%:`7|x�Y|2���(jo+-m1�'�j'f�DLa�z�L�jW�39F��P�u���g��8��ӕI~�pm�J&�����
��ǻr��TT�6m�|���#>�S��i@F
�]x�% ����ٲ���ĸ8t�(j�1]�7���9��u�:�@ˋ���v��۴�'TL7F�n�Oo��S�ݾZ�����C��^;up��6�e:P߀Ĵ��p�Fc3�G��$�x"��;D>ӊ���;�n�W¯;2cF����6
�0��}h�v���F��7&���L���
����w�ˋm�T��d�9l�)>��ͳ
n���rU�o�g�6�OqWL������2���)*k%���ɂ:���b�DDE��M��;Z$�VZ�����5�	2� r��m�<�v���4�w���x�g�Ɠ,A�-[c��e��FNG
_;Ťv0��(n܍�d}�u��G-ی873r^Z����%`t�R��]ZY ��4�먃��:|d�¦��QI]bN������|�G�#yopIP��q�e���yY[�9ڋ2�߃<ąmpbbb��L�@�0V����MJ(��[��4^��v�9��M�5ڳ&;�z�G�k���@�m�o�9��J`�_B�����QQV�MY�a��l�t�s�Il�F���p��j+��;o��Y�"�g�܍��qG�̒�K�p��t6��;K��O��J���7�m�	{��Y&̥+6"����+x�B�`��� ^�C]�*������H�|������H=���sM�Ź��y�3&'�O"��&�&�ob�-�y�������R��Ǯ��B�:�=� +K��FMLn󘭦�cG\íQ`�{ϻ�;v/J�L=I\����ai�/���sj7����uT�+�c���w8���FJ�.RyV��X�a��Ш�/�bW��Q���!L�+���dY��e�5wI�"v:����d���3s'���^�<��G]�i��]�s��콻Ǌs���1��9���5N���W�c�&f�v���R�J��p\E��p���Lu�B�%�[���G�*�aHw(5����<��r��۬��m���u�X<�t�Gf=��S�n����6��+!{��S��|���l���7Yb=΋��Rt�r���,.��W������:�z_Vę�;Tkev[�Y���ϣ\�����]m�׉}����m��OkcQ�| ��UAEPQ�a�0W-)@r�f\pE�AI���,QE#iU��"�U��R1�"�PPq�*�VEX�+
�"**bB���2�
���\%IF�(,D���X��rٖ��X),X
�k
�nXQ%J��VE�PFE�m�m�A��DQ�R��X,Y"��,Ƣ"�j��b�E�����`(73U,E`�����PX�KlLKQk(��k���,X",��,`�@��E�
��,q�(��T�cQ��U���",X�*�(����*��CUT\��b��ň��V�UY�,E�S-1UX��U�mE+U��U��V�3%Y"(1IQULB�����Qb+�QU�Ⲉ�V�0Tb�
T�[Q�EE��(��aZUAV*���2���*b�R",� �	1ap���G��uo y����vES\C���M-��q�iv77���x��NJ'O$��r�p{�H!-�Uw=���n�r��&��ֺ��A@Ei�z��U��{!�9��]�����F�}z�^'38���s��Ϫ`�,�Q5}-jN���������r[�8yL���R��.�G��w܂��j��fukEu	�e�p�1�]P�8�ߟ
D�yE���㪟+��򊢲��L��w�rX���wp%"0J�R��O޴�-p���2���"����+�åة�t睞<<&����ڼ
�N��@y)���U����� (J�1�0a�
0E��7���:5y��u��i�g�X�p(��H�|��%:��I
^�8�]��e��*��8��6�`��L���GF@ʄ/$c���{��O;�����כ��۞r�#��<0o�g���9��fXrf�'�#��:�W����x�4�<��٦�Y�ρ]B�E,�;���������`>��S��q����]Mx'�� ��cY�&�phZ�U7�^9��:{E�Rd�;�s���gH�}�Z�Y}ʲ�X2�r|{DZ�e�z�4�k�D��N��Z��k����4�#�V��nj�;R�`�r{�=k6��A�{ƍܲ���Z�\����;��=�vm�,��Å�*,|k9]˨*�&���K�ά�F�KΠ�	o�0��h�X�I�$�:(�͟�����'��M�Od��N"�Q�B��)��>S���I�O���z��rc��q���MޚҮ�>��}v��a�D�:�����Hҍ{�m��B^���<�M\b����8_f�����U��j��c�H[WT:�*�"��Y{��5�,��r�4���zN�}�#��Z'�	Ƴθ��j0j�<XA9ki�R��.�1`�,��S5ШD:QxE�f�ph�
��*�bϽ{���@ے�"�H��O�F
O���o�?��;5yZZ{��k�탛mkϱ���jw�Ts����u�v$.}� �sDuS�w�gj���iӼ�iY����>SmݱH3�c�U2�}�=ΡϮT"ԱcX�H_�a�I��H�gJ�����Hk��)�9�xs����A1���"�6�6�Af`���n�I&�gw�(&�궻ǞSphyz�3I�q`KGGY�w�g�C�==���4x��#�r�C�Qܧ.��mz�;a�8X��:������g;`�{�v�Y[}�i�!YV��{`~�<3�J9�h]�r�0�;B����IIp�cǻI/dJa)����+i@�{��W�8�����U��-��˖�_mm2-8��өLh��²f�A�=�*_���F�+3-ɹsfh��T�q>�UQe����4fj8��]��^՗ro���=T�����|-q�щ��u�x��f1��g��^�X��@2s�Y��	�C�ݝlN�p�>f�s�m5��_���ӂ	6���o��/'�2E�JF-�}МwB_N�|�e�<���x�[h��Yfz!�n��0�<��po�(�N��t���}��44��}3�p��9,F㚤ٰܷb�.^�X��iЫ[�uYҋ��Eה��o������)���f���隕���Gi����P.��tQ]v}G@晑�uI��a�,t0ʬp��K<��ثƜx�7F�Tf�u,щ�����|}�[�b�tr���.�ؔ�]
����F����,���6���X��X[�b8�5����8_S��T3�UT8����*����AI֬��bv�\��)����)�Ͱ�>SE�ʥk�nB��^}��_����}����}x�Q����o�p���;��g4�͞�yO��'�!V:"�5��Mܱ9k���7���k]u��j�t�ʼ�ݽ#�q��m�)�l�iFC1�a2�k%F�;�9Mܖ�d���̡8�#�gkOČ���p��ryHp�ꆺ��BX=�<�+avPNБ���5�[�`��\�S[�2s�5b��wWM)�=[����o(�1��-��s�u�B�{�����/��P�`�S6����gӏ�us�[l�����7�^���n�]�^Su�9�|6�:]o����3u��Y�\����"��ڗ�(7��,���n�^�c0k�۩x�y<�I?����Pt�,�Yd�鵈�o8p�EZ�B���:j'j�-%�h�����u���c��wʜ��:���|Ҿ�}��o^��:�wR�`N��I��ıA��5�_<b���sUQ�W�r���F��{K�������1�}�[9đ����51�Z�M��l�sc���~�ע���/Ӆ��D64{-�P2����(w�t��:'ku�ݡ��=~��Y��Q��0�=��Aq�I��o���43��_�^]�,�!^<Ut��6:q�S#Wl���F��\��{]�䃺V����kX���:+��y,�j��R����>6��W����U�Y���c��������1���[x\��6�&XV_�Y
�/ �xH@f�c�=Z8�W`,}I����1؏Uo!���7U�h��E��ީ�^�&.쬽ʻ�v�dT��}N�q:w�^ݓ�Ӆ�0�$0�R��.������Oh圥#ٲ"�ē�o��1;D3�Z�`�L'_��SU�f�7�N�I��ӝ����W�^�ڹԉ܏Ũ˗��X�w�3�l+�� ��La��ue`�4�e]���L�17SX�n�o�;b�!�aE�� ��1	{Ӟ�$j�VY�)�������-G7�����'�z��i	�S_���W��#/�(���iF�>X0�ע'7G�b#��8�4X���y��G�urY�ʕ{mr>��>H�`�g�f�7KU�Y�u�2���T�ӫLbͽٞ��I8]�4M��$����
��C���1q{�P��!
��k�O��.A=��|K8�Cc�/e8,z��#��6�F�A���uZ�١��ޝr���=megu�/�]c2w�����r��Kb�aL���v"8��~|)ZPc���������j�*Q�˸��Lzk��'�յ)���g��D�`�朗����z�P��
/���y������;׶F���\}U���@V�p����"#=�N��{-b`�]D��ӛY��zlٷUeWM:������ݪ��,�t ���J�$�}��O�ֈ���{|�V��u�v1%w;ф�z�!�q��ù����1���ݖ��5����:s�W\�
g3����;���^lT�7Ku�v^$�2-�p�w��|�x��}6i:%��<�WG�u���'r��}Lw1��:���r�����1�"6o�oꪪK�d�z������n�x����$D���`?7�t�{(dW�^θ�]�����t��{�ٙ��CC�]<d�{�ri�9��������K<.4�r���悏W���]4���.�t���+g\;����A�kŁ6��N�1����YMx'�C�2dh��{��+�m#zt����H����`c�qߏ��>��dAL�Y���*����m�o���c�%}�v�.�������h+���j�)Y�W\B	t7��O�7K����C�ӺvS�%����K���I�����0I�/�i�:�|���u���疓XW�t=5 Z`t���ê�Ī#|����1*�"��,�ͦY�_m3a9��\��ʂ�c�F��A&���$�Cה�-.Gګ��r��Cn��&�j��ҡ��N��<�2�j��VQ���%���ؽ�\=2�6�ȴ�=��."�J��o�	��,��ο��y��k���L���<�2�uG7���>ːk֛"uM����xn���*
 �H��s�to���J-���˛�WQ���J�9�u6�t���Ֆi�Vxj� *��{W����"�@�Z��V�|/e���-�*�6����v�1��F)�fA�Q,��lEX������˓,�nh�
wk{�Ǯf6�� L�lF����f�0�m�A�T=Ρ˕�,X����5��t�sع{0���V8ۚ9���_ش��«"�}f�3h����_�A�����Q���s%����Β���=9Vס��he���E+�X��5�����j�f���=]ef��N	<N���:Z�-`��u�=�j������?�W�*8PB�|_[��u��n�Љ&������##z�B}�B���^Y���B����o��׊�̲�3}�l�:Q��r�(�Z$G��v����u��~��mޛ��;~AgϚ�]��mr�Ql�����8���4���¨9�.��)#���М�WN}��mh�#���<�^`݄�t�:>Zv�zr���y�.3�uG/��=�`=T��@y<{�=��Ԟ��k|��76A ����yL3~s��,u�:p��E�s�])�yg�7b��^0q��Ӫ�cJ�6���X��g�I꒔�F��"|�qq�d��y>�f��pM��R;V�f�N���nNWqq��^^��M���W��PT*'���e"�0�4����mG&)Y�p)��������Y�'>�&d���u�1[J�jZ��`��(�auՁ��\=5W4.q�1�����g���-�蟶sU�Q�w�;��F�}ȗ�*�(�څ}�bG����bS���e��a�\|�B��%8��p�[v������h%�6�b(w��Zp��3���χS��z���ꪇ���.��ӓ&��XA3��e/Mt���|s��;569�\ޫ8"ν�tdmbJ�p/��<F�4�Dp�Ƚ���á,����(��.aы��0{�i�9��O�L�,#�%�����u5�I��U�!>�ǱR�]U�O��[�ϗ׶T���M���8��-�|�ov���	�~'L�$Uε�?��j����+�k��q.��F�'���0��s+_:���'f����q�lu�L-vF���m�ֱ�5��Լ^<�g�jK�	���CL-�]����vU��U\Q
0oK'���ڄ���h���;��u�n��7VƔ*�u�+5ËyH���yIl4v*�	���7��:]{�vŉ���ql�х��K�OG�n��W%���y�lʱ#�8{�ސT�/i�@���E���j##��X�������G��vgt���#�Gul���Db�:a��|��������)4����g)�J�<h����^<�ل1Զ�	�xax�����TVG<Gރ܍n�^a=�C�X7O{Ws�������z�r8nM��3��#"��rՌ��ˌ'�y���a��w�kt�d?��AA��G���x;��JӃ�{@Cj?x��YI[�{ �O����-�~�x�p�-]!y�]?O1��3Y�S��JB��Vyy���6����YU���fU���a�]�`5�]l[�z��5+����8s�Z+�����9�u�,>������T�FgLp�����>ٶy2����9�C��"�ͽ�Y�z6�ӽ}�ۂ!����M58E�9(��`�z[�M��8���4�L%P����MRԜ��c�����#y�;�ǭ�1�${�A���1#U�VYQD j��8��x�V�t-z�v����O��5l�t��Er���J*�+J7�O��˦ƹ'�)d���y3v[��OQ�F�}T�nzD���T#ƈr�f�>�Y������cV�7xsg=���ڙ-I�}�(I��%��D��q�?��ج=4:�{sɏ��9�C�*<˗4�����#���	��R���9�>�����eB�Zԝ��I�G��c��r�F^4g~K�f3�%3(���2{.�G����p�xI~��2مg��5)�"b��'�f���r�ԇ���c��|q�K����T����p�Y�cA���B��^F�:�
���{tG8�'�O��]:������]��C�w��I/(��7%��(^rZ}n��P��oz�5\�<��ظX^�Ic�H�]7����䣭��e��2�η�}�	E0:\t�Q���C;��p�$�FrT�wbx���apS
��_�6�{ӧ��~�΍~n
Ue��c0��<��@Uj����S)��l2w���Ҏ��M��3��Cv)Eqy���a�^'k�[8�vM��؇���5����<�9��o����1�^�1�*Y�G�xU�2ߛ���2�A��`,���"Qgsk/5�U(�̝;*��L�2��v�0���L[~K6��i_IÙ�:��i�q��%R�l5۴��r�~�]�[�6<f1�u.�ye�m�V�N
�D�&]C�1ƕ>�.�1\��/�J$���r�z���:S��W����,xh��|�!��v��~³�w�>�x��ѝ�W�k('��@����(����tJ{#Z��,�gv��"��x��'���yw��E����,t}-j��g��:_(��uCT3�ç�����9���y{k.VC�]v����wC%d�j�x�[�sq���o*܊���pW��L�|�$�ZAݖt�gn��;��lq�M�k)E}1�2��2+t!�u�pg��W]n�nwv<��2��K3����� f�vY����v���C�u�,�~���p�UV�-$K�V�W��-�tG	����&�vXi7��]*�nե�G�3�Z.��[�f����rӰ�/�jmK����pl�,#Ы\�3��gl��h��q����L�DF�ę~�����q3�XFؠ����ۮ]�6<VʮI	��c-hU���5�D5.;�-�Y��l!1�)�	v�YR�F,u;5�u=�EI0R�1��RdS�v�i�X�چnSï�,ޭǜZ��mpf��12�[��K��mދ�x� �$W���;u+k�	fC-٭�]�)wC�u�k��ܓ��Cwku�]�rRF���@+����`g������2�to�MV��c���ŵ�BM��L���j�܋�:� �)R:�U�y9��sl�Dm�h��Cj$f�5][��)�Sx&�~������{}�J_3s~!�O�T:�=�@㷝��K�R����R����5���M�,7w�q;��VocO|W{�9��alAB�`�8�O}�>�K�<�`�/��o���k���S���L�F)d:�t:ɱ���G�s�K��t_A�P����ƠZ�w,QN��[��s6���J�����]�nb��um"ٞ�w�X�K8E�W#d#���R��e���5�T���`�5Ks#�
���v8���_\j���r�7���D���;�����;g*�7��*ɰ�,XԌ��/!����DãHðf�r�:B�ѱ[If w���v��z9>������]En�:��SG�W�`NԮ�+�wwkc�Gމ�MO��M�Z�O��ٖ/n�u���Z��7�C���0�}'hEB���$Thu�K��^	����o7���S�^3sC,�Һ�Y,V�{Wm�T���L�R�X.�����a�a��QkTMx�Y������W����K��%��]
�1-kr�3D��\
�w(�{��2�����:�|������N���^�u�n_n����#&�k�.�G+1���x�;�0�5e��GA�v.B�����d�2b�,��f�yv�|�Ʌɚ�;v�w��[��5<ŔKŮ>�)Z��%̼�ng��d��SM��ޗ���ja�˸˭t�U�s�|�!�@��O��_=��K��t@��f�v�vY�n�H3���Ys����3t����{g�J@�
�XG�k�k;�X9�(�%B��m���:z
<��T�o2'��a�w�z+���*�񊦫�+�K�kY7\q%�r�ᘕ�7N�qCv���)|�gy�f�Q��w��2����S.�sͻ��0X�tёAA`�e�k)R�1IZ4Q�,-��,��+Z���0Q`������"�(�0U%[
��6��*��T�*�5bbҊȈ�)��+Uc1E�X�pVcS��1QQV���!X�+F
����chV,��jA�"�j[Jad�*�� ,�EPD1+
ʢ����*���j�b�,cTV�EA�����R
��#-����E�Q\(QU�UTc�*"�QX�J+(�b�A*��F�E(�@Dcm�Tf�R,b�Pb���U5�2AQ�L�Y�1����U�,D�TQ�8["�QTU�V"RV((���i��5D�*���+1b�E�Uee�,m��*R�IQ��-TP˙1�"�.f(
�F*D�9J�(�D�Q�E1�#����%DVDb*�58H �@%E��*���ɦ��z��ܽ��-j��e]��6�ӳR���r�����N6l<��[�d��"�1���q�+f��]���f��_��y(+�����ݷ]uJ>%��x����5��v�،�q&���EX�S|jE�6Y>���*%�ު�ŀ�r��b��'�]�b�Veq�c'�z1�{Z�Zf�p�mi�K�س�A^��2�.J\���=��."�����9��v)	�>�{�㙓l{�P�ܕ������[2���ӓ�bn:�"!)yp�+�kTk�糺V���h�r	�،4/6`�z��R5\�.P����B��z/6ẻ�v�%RV%i���kŤ�X��+"�|+��Bb]�8E�U�<Ȧ�φ�n�x9�`��(�Ga4)6ilT�Q�©�42��_՚��q`I�8<��u�Ac�؟3�{�	�\������(�b�gh�T�g�E�v�����<��c)�i;9��8s�lP�ʸ
�GS�sG��1�0���I�>T��-qʽv����}7���J�WH���/cE*�J��n_��玓�	�C�g[;Yw�����)m�+�evo�b�U�H��v<�E�b�O�SB��N[08��� P�[R�l{��j��K1�jsf�=��GV�ӆ���x�Q���2T����rc�nQ5�9!h��L�2X\f��p8��!�y���]�Ĭ�&���va]�+J%�۲t�7���=ݤxҝ4������d��nRF�n��NR��WӦ�mt����T*X3z���]P���EL�7��e�c6[�ce��x��1=�7j5��S����y��*�������a�\U���������W��/6���|e��jԱ�U�x^;�C��L��˫y����o	�4�nho�z��*�hO�C�ˎP��dĎ��	�"7���P��/�*�ơ��7l��o�mܝ�,�B��FD��Jp5�ySI���x���ݛN����g�O�z�|��Lz
��=gtI�:�t`���UU7FAƯ�s��Q�Vi�2:�\��������VpD7�?A_m���lIQ.��d�TX�ٳ�֎i������tS�Y��(<�i��림��Y�;n��+aW^�F��$\ț�sC�n5!��R��j���[���}{eA{axx16+0�p�	�$7�w�܌�B�o�R��)>��7M��^7SK���#�|t`�'�ƨ�Fژ��e���B��_c:2�wX�`ѝHT��7��ڻ�ɫcѩ�!b?sY���4�Q�����qِhs�ɛa�=Z� ��ԥ%�wB�.#�:��A��Z/6.���� c���Lᐵy3����.��o�{���ܶɅ��h���T��S�T#�2�°2\t��co�Gl����z5D�ٙb�|��U l.��J'��څ��IFv�؊�k��w�d�ٵ�ٺ����p���"�gHz��f��DN�	L8ȋ�^V$�쿏bX����W����͸�����H_c�ep9������zA��b�ڨ�ܔI�S�DdpםblЮ�aK_f��MVZ�f��Q���7BTq��E�Η\�4;[�/rFd];�]��UDF����a�V�Qa��X�n��ً��7�}>��@߈�P��:��p|=�s���_��9�bDR�DcwZwc��~kX��Sp��YN�/�*�U���8}�/�i�@�����u>݋S8Tt�Cp�=������g$���M�ɗ+/�be��C�V���Q'*�o� ��hO]r��R�=���,�Fy�:v��F��)�8�ug�:ekڴ �+ŀ�m�O	y�(OW��ڞ$d5,�#���K�D�Uu���d�].�h���6������,�4[�%dk���w8ʚ�x��z�pM�趯1z7G�F�[�Dk�.zXHk-��8WcdU�51Ը�`��*U^��/���gD�]���.t�U���|��Kn6`]>���8�õ/���'I��ɓ�2K'�JeS'(9�}J'ᨴ`��	VyAYu����Ot��C{Qv�)C��d�̩�D�?ĵD z!tbD��.����YQ���Ϧ�iZ�6QD<��eH;i���!�U  U~���Ȓw�+H��2��W��6��N�%�g(�}9��'g����yv����<*`�"YDྖ�'w|FRdq�p�p�����5
��]˼��1��6K�1i�J�����{�9�*P��Kb�k��,w�K���R�� 9`@���������b(�W#}�vTߺ�
��n`��ܽ�5T���!���|yVޫc�no�x2§0����()�g�hfY��j��T�� DF �i��Vd�e%6h�e����!v)Eqy�p�C���3�yU�WB�sް<�Z��� �C�6�v���K:�9��.w���9Rͨ�<��p�����C-pc(dK{*ߩ	����T��'N�r�nb��u�C�ܸ!{�}�ίfXrb��ZY>�b���ב��Eޥ��,�zQf�F�g;������PH�2��Gݼ��,��X�c��O8s� ��o���Cy޽ri����Vs�o��g�u��=/1ӷ��:�罪�mq�պ�8��ۆV-�"������e���Y���ۋ��	�u�4S��Ŝ�+�p�|;6��{^/ܫ�N�1��ǼR�N#�y_��f'��n�ޚ�*4�O�*�)���Nެ>=�`%������gH�I�I�(o�e_n�O���ה�e�U���Q�;�R�E�'ܶ���Od`�>S���/y��/{sS]���?�r�mj�C���ӿ>����&\2��(��[|J�2��݋������D9b�=�Y瞚�қQh�L�:Ī#�����W^������a�*�[���Gc�X��X�!����(��D�'�*%�ު�ńӖ��۩{�P���r��5vqvz���G�p���+D���z���-���H��.D"7�r3Lu��\���Z�P��7r����e.3��ܭ�Vp\��1&��l>��%��fN�Օ��R������I�W��e
����&Z�Xs�͛�!��Y��!С��V�S��]�y�ڄ#ng&"�҈�R�wr���ZL�*�,G�F�3]��'ȃaZ�8X�PS�k-��^�4ypڭ�Ae���*w�ׅ=���^B��-��m�y.
Ys��U���(��XY�o��VZ���Sq���e�ْ)ԅr�3��2nG }�)��l�%Q�&�p��jtt�˘���=0�a��Z��X���z�4�R�n�/v���)��m��tf �΁�9���y�7���5J�,	:��#�[�'k[ͥ��6�µ��O"��d��j�'�� �|�R�s�G������t6���W�l� ���$��N���j^���Ln�,�g��I�_Т;5e3=��	�7öf̒㳶�*�Ҷ���$k#mS���qа�^6&�,v�ו��匈�)fq���YY�ix�����+��L�s$]�H������@����-;`�㓰��P�h��R�N�z���R9^��(6[�ceI��!��/ve�fT��ݍWv) ��sj����\�C��ſ;?ex��@�(��m"�K�e�<����Pȸ���%e
�^.���S=��-ۚp�K�����:T�l>%��a�ߛ=���_k����wW:��p�j�ۗKc�?g��E���ˣ�*��\|���9������ܦ�X�}S�a���~�N*��7���'��z�����6�K
�Z�����;$�qĤ9�;>	�32q��e/~�t���[�/N���0�����d�Ҫ/q��L��Ȁ�yB�s�\�H���s�s���JO�፞��PgE�R�J;4�҅;��_N�K�6tG-!whJz���Yf醌�Evc�w�;���������ת�y�b]%^�L�����:����4q@�sz����^�;O+zu,�<�Ce#��8�o�/uj3뤸U��uk^K�/�[��.^�Q�j;��N���*J�5���z"��}
�<rP�^��|�®/��C	�;x^��3���Z�f���n��t��0*}�n�S����iy��t���0�r}ʚZ6�v^��ll7	
����ك0�m��vF�vmxv�����zfm=�\�z:�',�y|kce�܅347��G��6�q���|n'j�-%�h��0�Y�|5d~;x�[��Bç�I�~X��Tƒp��U(:�F&�dI�d�h���3�.����TO��Pz�|�C��K(�v���LW�Q1#r�$Pk)�^�zJ�Sv�8���nyL�p7D�/gm�,xzw�,.���Ʊ�������X�d��.*>��SʘM4#&&�u�����ł�����9���g+N�<nP��g��X�H;ͩ=wH�K�J��;���S�)\�v˧Q=�օ���q4��-�+����.3��h�0M�6Y����s)֬7#;u(Ƨ�n5���닢��:ʀ��=Y���kg�w�*���F�Q����uc��=))ғ4�uw�mu`��'37B��42�Yca�O27֝�o'O�E���yM��p�L����"-�f_S&kw&�sܷi�O�ķT��{�����g�`*��ݺ��l�f'\Q��Yy�Zٷ�ܙ7��� �������/�MG�?i�!��e9�#�
j��V�e��Y��wb請8u�OM3��%P-D�!d^B*�ol"Jޑ��%�Ns5vdR2&���̀�uΘP�Z	�!�^O�Qh�|a3<���v�A)�r�F�n�.(�Z\qՁ&��� ��N('7��p�@׺e(�m�T#b}����8D��|c��j��6��FL�Ԛ�J���5��r�����2M.�$�V؁!dP�2����y��ޙu=[�̓x�oM[:p�d3BV��x/�E�L��c(����&.��L�*�/2�kp{+֫.d���rℿl�t���8��e���p�S�<��ظZ�i+;:���z
��;��]��"����)z�����N�W�V�stn%"0�J�N[lED�������~k�{-Yݭ��A ��d�[�u�4�����}���8(��V��dE��iŎ�ؠ����*��B�&7���n5w������1Cq<����1N8y38�]Φ&�C���Rt5�vBG]���f0*Hؼr�I��h�]����Zr_Go����,�M�|e)��(xkJ
aY�~���E����S�]�@z�W��G[t���ݎ�RAPz��
�.0
��W�Pf�~]���,�P{
ߵJ����no���RX��͜���O��DW�#�\�13�,�J�{<�����!��Uxl����4R.�w�2R��;�A�/:�"�-�z0C��\ssm�r����>g�0�~�r���^�(���A�n�Z��qg.K��yh�����kŁ6��W�c�3�?M�]�{�4�R�8�5�>T���<G�$^�Oa�)�lg�:�;N�xG�c���d�H��u^�)�u�+/�V]`5{R"X�"O��Pմ��Od`֩�jmu����s����{y��Sn/K>��%M�4�."�)e��2�HҊ�kfW}���t��%�
��s�,�c���&�4��3�����B��v�u����E���n=ox�Hl�8`ɷP�LM+������wּ8u�A �\/$4�-�^-�[���������Ոk��M#	���x��珉��#�wg@�Օo�^�쮏��N�m=-�����Z��m��9�1������`��;�w-��T�:��7���a������,�Ђ��Ɏ�Q;�Ү�L�q�?*2ݗ�1��,;k2l�oZ}M%�^%`|o���\���l����/@��L��-r-#yX/p�h˖�;.�3e��>�#����GsՂ�c��r�eY�r��#;f��=�e_=�WZE�s�䁉����7�ϕ.f��֓��=���`ͺa�R5\���,��z�,�Y�l���0k�i!��$��\}�s�ey.7�@���Q�z��<ssf��E�-#TwT6C:�d�pB�h>fV+�5z��1��y�D>Xj�N�(L����me�w�5�Ҁ�Z�8�y�����]E��;���=�Z�i,�xJ�����N��I�k��-����Pg
7��b���9��~��"�0�v�^c�#��Bʔ��ŗ�ɝ��=۔�ݹGN�Ĉ�6ո7"�'(M:{�����Η���7�N#��z���b��)F�g*���š�/	�E=� 5�w��vyHn��쥽�*X���"������,_��H��0��R9^��(�l��Qu��_:`!��&7Q�c��	���MM^�c]&���E�!U�?{��[�ۼhs�Hwז��xdS�o�29�AtǴ��]dpZV��b�a�����??A�R�r5'j�\��.�*����fWv"�p|��2�<=�(rq�PL��� {)�o���}[�&����^X��ՠ,7��U���N)V;r���KK�=��vDS�!9>�ak��V���	 �{1l=�t޴�gN��r�Y1��"���6���:�7��nnJ2C�{_`����7�zd:�{;����,t�C����i5t�ν2�kVf�n�&��(��P�{��oq�٪r�l��s}.���i���u�cp�V�w;���(��Z�ٻ���'t���b�:���/�F���Rn+��w)��oS�gQ�[ٵ)�L뢬F�sf�v��:q���Zl_.�P�I�}�AL��9�\
F2}�i�p�i΃q��E�o{�qLK҆�0<-���X~��W�}�g�#A�yƞ��*"/Z�'�{Y�����q�GSV�|�����x;^i�&7\rQK6�����jzÈ�)ĥu�,=����(�.�i��fN���v�&�# �P�l�=�z�]i�2Pe'����otY&�QDU�����̲�q)i�fZ�Cx4�סh�O��p��bWe���ڰ�Q���j�P�&�̩�{�A'Qd����=�D��4�5���
[�[��:���Va��N��4�H^�+ѯ'���{�H]��Q�l�i������]"1i	XcLNi{ɬo7�b5}�C�F1���g^�>��g�\�7i�:,4:w*�um�ԁ{���,�|�|�b*d���g�&��R�����Mܒ�lr�*̥.�=�A��U��iv�+�|o�R��	��r�,��`�NJu܍�`�j�lic]���z�����m�K��@[�7�E�?*�~�n;N�}A�9)ZZ�qR��9�t�����[�G��e�f�l���e��E���aֳj-k��y��s�7��.U�no^�{.��xPR�l�-�-ˆ��U��N��������W7PY���ƭƭA���P6k�ˣ#{�9^f�8�`Y޺��'):�\��J���w��c)w9Q`F���N�� �֮	YŢ��j[�x�v|r���sQ�5x=����Ӽփz8:�n �R�]��n旳�D1:�q�;Z���i廂��֩d�JJ.ՓH<.TАj�N����������jO�jM������pClW��('�fEF������ʚ^�3/xO-։�&6��5�_�-2�����蕃�Bf9l��J�OvM�!\��M�฻;׷�g*E�2�<�m��,]��7�m�@˺;�?��1�}c ��F+��%C��_gfl��8ȉ��2�̘��޷�[��<�ni,U�_l][1�AA�T��5mQT̕�Xe�-�U��h+l
�*
�k�EF��ѭF��m(((cr֥A*1���"V�n5cl+r�+11U̦!�UFe�ª.6!m2��R*-j+YU	�Q�آ�K*��+X����UTU�+**�DQV`�)X"��VZPKe"�PUY5�[H�Tpj"��EQE
�f-��,��m�QQ�Y�PX��1Q"9j�.!�`��Y"�(1QF�V��)V�*�R"�*�&Z
L�c�X#b
�m�h�*,E�T�B�2����"�F(��YYb� �E2ئ4j�1�Z�c,dQM&���1�f�b������\D@\j�i��(�5r�Q,�(��FA`�2�E�c���8��dR2""��DUD`�+�V�F2c5�L�������/߷W7�d�o��dW��+֦]&m�I��&��Q��Յ���$d=X�SY�m�]���T�9����=.RTa�Y�,�Oyb|!��x!�ط�g*�'] o:Qqci�Kol!V`�7b��-3k�abN���>���=�W]�G@�AV�*Ca�)V�`\��n���St�NFC�eo��
]-��'ٶݳ�\��sn��s�mFx�Gnan��R;�U:��2Z���bg���E�%oi�Y��i�1��I���N[��)m�:��W\#u,w|�ъ$&�U�i��ز�Aͺ�N?tLex�KW���>Ԗ�U��/u��L\�P�=��9t�g�K;@\�}ip���t�=�4�������P�ܫ�s3ͥQؠ�˔�B� �2���LK��r�C��(^�b�R�{QP^�QB�}�����G��w	���ɇ�~uJ]��� R�ў�mN:�]g��uq*���;�_�V[�i|�gM"4�VjY�7�U�3�;*�qvF�n&.���}k����'Oʦf�/���k�3�٫��L�h�
�S4ZtN��f�eDC?	�Q
�ݚȅyu�:_�Unu�6k��=%���,G^��m����<��9�yv���M�T���S]����_�GSG���άF�#�!#�d�'V�S���aB:�+�����y�V�Lǝ۫/8B���\�Pv��o��"]�ݏ;zV.r����6޺�e{�A�V�W��B��M('R�"'C#z;$���|���Wz��+���rJȿ:3���VS(��ڳc��D��HƲ��o.D'SQ���=�T�� �����5�e�'<�J5��o�X���%a���``=�J��XeЉ�]w���R�,b���%<z�X�Q}�+�tw��b�f�J>�ʤ��2�փ�J$r*o��J�ip�b��TC�,��u�v07����(�V��)qd9�5g�_`���dy������q�X���'ܢG*�o�.��(����'[xdr��D�<������<-c�s�O:o��2`>��OW ���q[qR�7X�w��p�+��>��yv�b�j(\JɄ_0�ʇ��]�\�k���O(r�A[�,b����tͬ
���4z�[0�����~�5l�k��<���PGyZQ�Cdj��L��1�ָ�*��1����c\��c^d@8d k�R��M*���0]/)�ϔ�v&�r���]�/Sfi�U�����ҷ���2��3Ū��b��W�n��Z&2V,�"\�X7�|	���� �{>��p;�f�Km�J��3rޕ�+t���p��׷���qN����Nˮ-�Ztu!}j������t���U����8�i:���i<�c��6H����[��Ϯ^��P���4M��$�8����]EeY��Κ����Zzk���o ^B%�5�!����+*n0ñ(���'<�m�+�r4=��RWw�զ=��*25��cgK/:{��gX5L׹HV��r��b[S-$=	���[�^gOPH�$B|�?
D�,`��d[R����y�_�R#�%O/v���9�?d��7/�2����v'���pR����3�C���_j��F1�7v{e�љ)X�0q��A쵈L<+�1,��T,���q���3�����V�=�o��˼���C��'�;�O�Z"�����18���y"&n|��c�۸;|jn�8������H�F�8�Ŵ�C�g������ݡ��݇@�����������m\�)��ӇHC�E��uC/��]L�ø��|,z�h��V'�mb�FW�K'��9wt�#�c����$
SN���5��W�M�5;}Jq��d�;���`�`�������^Y3)G�'Q��ANy@ƣ�ֺ��HY{���QV4H�9�b��g�*5@��E�;7�-¸j�q��e�W�|V���p�*h#A�g�ݥ�aM�&�"�'L[��^���+6�[o��yJ;�ܛ�o5f�v�y��R����b
�����9
�k�{R"s��b�;{�9ꮞ���Pq��=�X>��2@�s"�n���[�W�ϼ~�xªbN���ļ��������Jf[x�v���c�E
�`l�sX��9�Y�W�
mE���+��$*i�m�Z��W��etݟ{v�V�5�۔jp�=�Y��g���,>3ܷ�'ܟ��.�Q.F��\x�Ӟ�"��bV�����{�X��_�ϰ�?� �,��S7O���n����'TX�K\��ھɻ�%9ݩ>�x�T��*�Єz:ĸ�z��7����ٕg��`��SD�}׳oFi̖��7���V:d��%U��<
�����;��(�ق��rR5\�!��S�=���̈�P�w�HX{������ן7��ZL(a̋�����0'0*�ґ+�5X�(T&�/����)�UD"U�#3Kc.���g���lf���.H����O�s�:������R�y�����l�}j5f�����LK�{�Ta�)��Z�U5�����rjژ�r�w�r�h����B��)��JX�XUT��C�ĩ�9~h�&�3K�� �c�L.�+;5�r]����f&����F��y���j���q�.����K����`+t��h�Nj�9r�ˑ��2`�{�^.�!���3���(*͎�b���9��5�م���9:�����;|�WE��9���#_&C9W�ü�ۖpli�H��V�/�W�԰�񹹮Σ�uH�F+y���q�����^Ag�k��0�P��X#�$*�ێ@j�ﯸ�	K�-�&���+�<�dB��5X=^�|���ZE���w|r��<=R"�\e��9��WLZ��T���*���+v_�Lw��%e����݋~v~�4*�@�B.!j�sA�+4`��.��ۅ1��ʡ��/#PyL�c�����6;h�2:���P�y������Q������~�J^R,ד�fԺ[�O�m���Ku�)�G�6\/��h�X��sq'��N��+��Dl[
�b��W2Qj��bx�5����3 Щ�,�R����[hmz�r�!ė�_�6%���^�<�|��Vm�t��,�U4$7P!?O>�W�g�?�����p/��.AC�u֣������`\a�!��x�������UJ������	�43=^Ž=�s��0|L������29<�*ܪ��j!��Por�<~8��3ۗ�w~�.]d\�oc/���7�1���Yo���^�ӎ\��A�'$�aX�_S \h+����v�8�yN%��2�
�G��wTU���1]Md�!c�A$k��Q���䡽Y�B���}�z��mŉ뼧���!	U�C�>�4���&��\lI�g������<�«�2���oӽ#�޾�~380j��,{b�`�0��%�L'��pE�N�<#��W��+qke�<M���YPsw���b��3C\�kǪ�6�q���O����O:II�fT�^�坨J�(���c��ܩGj�l;��r5����}���QbS��_�1��/7u���������w���'إ����o�I� ��b���mg (��[K����v��k`>�#���:�9<ו�9�W(�.�!��۞�:�S�=wz��1o�p�$�ݓٵ�M�h��X��	+N�;;�7ژ�^����f�N�<nP��m{��!� �z�-}Ԉݍ\�t��a��\E���WZwc{\Z�+��<�����v�����OI�������#ܣ}ʩ�t�1�,��[?3�i(���J����śXq��}�p�b��~�*�j�{�g��n��s5����Z��^)9n�d��.چUs����[���K���z�à�l��Kox_m�ۦ��%k{��e�G�6Cg���7��a�*}0�e����F���?g?7�[�{�ۼ=n+�:?Uj��nc>^ ;<"1��w��
�=��%����:�[)v۔U>�%�4���)a��-�ϩ�3�]�娃X�,��EW��I[��Y�W���O:�R>Ω�({����U	�.�)b�~�5l�|a;�Q�����CvDN(*�&(�*��\�pO.��$�XיPp�@?�)�S]�f�,��Q�U�޷rV��"k��~����Hإ�٬��s�+�������PM�4�a[1Ę"W�힒F�w9q�sz��������[K"�R��	x).��#Ě�\�b��c��g$nZy)��ɴh:�����Ξ�gY�g�P�z��n�S5��eNh�qڛp�m����	�M��^豃�U�P����)��k���H�4f�V��9S��o����/]���Q|9� �e�ǆ���eႲυÈ���ʭ+8T�K��*�s�1u�/�1�,�A)����0�b�>�BVE�єs�P���7��ƈ��JpmTt���f��
Ǌq�2���+/I�CD��xy�1�&�촨��B�U��N)��^L�B~�����W*��*�	j�ݪ�a-�"3�`�G��`��O��;�G�m�kg��_>KyQܶ����S��^�o	�^��&���Z
4>���c���DVG�(���3^�vfOfX��o�.8�*�aқ^�����ݾ0C-@�������R�4b�g�<:i�������;ȼ���ݘ�s�ݼ�5)t����LÖ��/���^�A��\�gT>���|,z�hὝOϓ�|����ޢ��%z��~X���k�S����- ?�i�([͏����o�^U��R�
�����ۮ�rAZ��:���G�ëD�ũ�J&b��]-�7�R�E��G-��N��NN�W��dTU��K�w�!�J�%LxfGw¥����Q�(�MI����b�\n��ꉚ+�'���:����t�[\qy���Y�P�ڋG�q�TGy?����}A1��m!�5�S�>r��m����\�<��I�W0�m��q�j���ZW{��a�����(N�i��]��{�f良���f��S7O������X�Q���<N�ڰ�W�s��䓪�-F$p�����C��k��l��E�[���lʳ��j�w�+��|;~T��*��{=.��F�R�Ln.��..w�����/*�*'�'t,�mi�G��m�B*\5	���ֽ|Z�q�ز��n��Sa���l��L�Y�,Z��u�L�خ�sC�wƦR�[�"�N7�t7��O�7��i�$S2�/7��Av�AQ�H�H�v�A*ג�8Ǖ���2�����[���{�e=
W�r��,�"F�;��B���n��^U7��Ť���+"�~��≻eڝ&������H��f�k�Lӂ�#�U��B��il`�^��^6���N�v�X�ScO:z��_�+���c�c������s�t��,��&�;��M�R�ޖ�U��Ga<�y�n�:'��(���p�Jg�*� ��f�g�C��揍��ݖ<pVX�I������{��6�V��ג�����7*Y�li5����ڑo��&����Q�d�{�w�����t�>f�Y�r��2�171���!޻���K.o��.S��/�׷��J�v����K����-h�"�wvn��겁��n���d�bs�؝[������Al{}&x�ʮ�U�C/5�8{���]
[�(9}�4ѷ�	z�_�?t�pӰ��Ṕ��a�ڧ�����0in��ލ'�hBT:�<Aw�L������l�l�bT�1(0;�mP�����'%wo���P�����sm��л�L�γf�=��>�:��n����n��wc,��/5���Q��0�W 컻X�Q����F.w0�=}:�l��V"`趟h}��b�K*3zg9�'QOY�Ϲ�l5��å��'����E�>�o�]-���5�g'yL�)�G�^֐�i/����q�f4�9����v�L��L�1^#�,�!(��{L��(CX�:E�bp��\7�i�[qNƬ�7�uj	ޘ2���rė�(���3]񋽋(TSͺ���I���j������"�K�z^�>�wh��\����]Jp��<����-�̜T�u��ܾ�Z�P$�]�`��*哞0�X�D�H�D[�j7>�P��rP�k�WF*�@{��ޘ���[�'�+����M�÷j]��� R}�o���*�����̷����3�ʕ�v8FQ����t���,��u���[0`
v�L'�Dg��v�t�<Qi^gy�6X�k�3�]V^�u�(y<�I?���nP��h������N�i����`ۧe�=�3����QU��+ks��[��C�mUdAfЀ��QbM�Qx�������ݾ�\�Ln� �%�X3 j�hϊ9\j��M��c���g�}Z��y�o���c^#�OoS�������&'��Į���s���77i޹�ea1PE���\{tw E��"�N�iss3�����	���vxRy1�0�l��fQܴ2����):���Q��O(���)c�r����N_C���@�z�AkOl�x7�'K[����hJ�j�z�I�i���t��,7��&IZX։&T�/�]0y}u+ /E�͚X��㦩5�e/����UJC����3*�"�{ȹ�s04Z�#���R��m���&��0��}�	k�������F���S�<~s�,�!ݺ�Na��(p�
�f3�XݷKz�3'�}�9��w'd���JH��vm�_y^�7q�<�F�Q�P��.���K�g%��龡�z�L����Q":�4�:�F3���P�
6��6����,�m`u�u�ԃ�	�B�a�fp]s5Gj��&�s�@Ҿ��Զi���Q�s`�~�܊}���o'bk�h��+��8��9$�*�ԓ��!�{}�o	g�e����ϟb.a��Pp��k��u�p9F�WN��܎��z���%P�-k���a�h��}��לxԛ��c(�vzvWP�t�:P��f����[4N�ʩC)80 �eWSH��԰��t"�{�8��خs��zNm�cF�N��̩�e'��촌�ΰ�̯��G���~�,�f�8�W���r��Z����gي#��6n$�T}3����̗�܇�T��a���鏪P��E3�\Z���Ԥ�v��̛�;dΙ�q��۬'rJ�J��mÍ��C.�6d��w&v^$�t�+��ӂ�	-
}Z���B�}*>�a�,~�2O0Q�}pM��Y�S�6->$g>�\�q�u�n����ij�J﹝���E;���R�qRX�N%�F��ִl<
��&�tmH��ռ��Y�}d�r�gu˽�@*�x���0e,`���U�Mxk�<A�zz*ZWuq���F�K�/R�1nw
��sg+�����978n�vwK��	�(����É��Q��pd����#�Va�D->�r�^�����ۈ��Uʅ��7��Y6�(B��'l��:k�7��э٬ޒ^�L��Vr�:X���A}��T�{�۶J4��Jڵ:m��3#[���u,�6ܚ����X�[Y*>hm�v�)}�+�ާɃ�.�צz���� [�y�]I{wA�X��a��ޗ�Ԃ8{<�8��P��f�����e�W�	�5.M�Ʃc{u����~�>~��.�^W;�ՖQ�}������>��3N%#=��wjgV�>Wn�z�����m�v츽�4�3�F{(���@P�߱�'-�@�x\��<�󫬁�>���a��ܶ��_,��3-�*Z���W_y�ʵ4��֌ܮ� �jZk�LA��.c[wێ�ʀ����DQE��\ �����l�����!hX�*���QAQb�Ղ��V
��*���ˌč�J�TT��ʈ��j�[D"* �D
&Z3��X��E\��e�*2��UQ]Z�*��Jj�H��e*5�"�R�1(���b�L�KJԭeQr�(,�Qm�bcUJ�Ub*��Q�""(�e�U�����Q�Z�E��YZ�K�ZF�e�"�,b��Qq��h�6"��b��TPE\����uj����j�Xµ��B5��8�Ҫ.��3IE
,tؙJ�+[K-+M4QEf0�%"*+Z
"(i�(����m�.���Q����2��Rґ�1UA2�R��DW�U.f
�>�x��E�k��݃/�n��a�E_Ws謎��E��Pq�����\U�R�T��3�Z���b���Վ��Ƶ�U�s�C�ݵ��+���Ū��w���$�^V_܉�+�a��qv�Zl9�#�SC�g;
>�{j�~�ݹ4O)�az�A��hn�q�x5����M��\��WI��	�}�tY�$ꬽ�K�Adb�28�.���\E���]i݆�t�X��=��vz��f���r���������<T���g<|m{�O*�v��p�=�����Uw�n���c�6��a3vf����V`���12��],�g�F;���
�=�İ徣���ۯ7����=�b�v�7�ST�0�aՕ%��WD�����B���Ǭ9�8'1ʾG��-�8�k��6X�$j�:��)��7��!쯗���Z0m/(K�(+7"��Wnsn�h�c:�f���`�8'�M�w�y�E8d z!(͑!m�L"]�X�Q������5�W�dI�ڞq�KU�YN�Fd2J3n�k�	;��!�/<'�\}ٲWj��\����YG������ňr�vD���l�jV�Ȭ�M������ew՜V3Ή���]
�C�GG}H�4����y�}.� 9r��2tk;*nc�}Zg���jx�(w�a��.[(����L�S{/	:��Jܾ��mt�{^-����;_����,��鐗����y�Blyw{z��]d��s��#;M�RN��,���I@��O��V������z6ka�9.Fu�T�r���N�������']��U��N�I@g$u*��"�Uq�Vp�Qz��ίT��k �p�7yK E��Wf���j�`�3��M�wu�*�Md�(�:�v�aa�b��uz�2�"(���]�5���)�^Dɦ��9"�ubp=��	��v��(3q��@����~zh��7yݣ�{^�&��J-����O�ֈ����.w���9Rͨ�<���R���{3$�>��H�����!���d�P4ln*q�i��t0���M��&�Bm���U���UB�������ϭC�����1垗cY%̏ø�բ�u�t�3cz��d��x --����c`��ǼV}Mx'pTid���Ô��N��+܈9-�j�Y�hL:�\=�\y���<F�Z+Z}Y}ʩ0r��D��R$�\~>�gOUGF�Z������s��-0�HcZ��Es8y��
mE����Q�*h-Ϯ�:m�D�6ފk[�^�u8�#��z����1Y�ζ����%�n#�В�Gv.�q��O6�G5	�+ޙ�@#��a�C4���p���w6δ�T�zs�x���;(�J,��%.�y�R�a�K�iҨ�|����+^�̧^�I�H�G[���R�{��{��18r>�eS���[|uy���<�]������`��HTӈq>���=�/V%�+�vХ=[�y��5�(��o&&��[���Yq��E�f�V��I�fSy���Di�>3�Ö�b��&�j��zT/�P�ͽ"�^���V�ǲ���B�R�����,�]�������uJ��Qѭ�&L���"��3ާ<�h�ܦ�$ܾ�1����;Pއ�x(+}� �sDw��#��*^�P5��t �j�F׽��ϟtB˛�����JhV��G+�9JYP��$ƒ��o�wr���]���ey(,Põb��99��}6/w���E�����k��87�!�U��XM��sN}mzx߆�낊I���{��m�G7�o����")_,	b��5̠W�2�9'6�J�P�����%����Q�m�y7��^{������{ΞJ�%Y͗��C��揍��wG�XK%�p�r*��c�gE�(���u�{�\r��b<�y�8<�G�A?>q'�^�Rqt��:�w�w�����&<��R�[t7LL�#ffS��ի�����#~��.�7�k/���
���&i�e��Z乔xf��- ��z�#�(Aw�N��n��aq��f�M��RC�S��F�%o�9�-��{�J̊t�˾؛KӍ,��M������G��M_�/�,���]�V-u�~HU�w#���N���Y��{X���kpǛ��ʾ�/�zb��B�wvo�H�v%��D:(��f�q�@7=^�V�x��[T���}ӡ�������t��=sjr��bE�팆�]���|'75�t�,j�\X�EҗP͎�C���s�guy�`�ݹ����z��da�mg�%��;�Ji+F�C4��W�E�"����.��b}�m�:�+|8�����k��8u°OT��a�	6�B�����2��!u~��uP��/X�:Fl��1��q*�a���loc��N:0`=P�YUP��g��CZ!O<�"��8��gF)��"Wh����w7�O�����7.!a/?�T�5ڌ��.a��θ�T�/$F9T�Q��\*��lCp�K[�YN�d�!W�� �����R�vH�v�:�x��1f��}��7OMi��\__��{���6+��ڗ`p�lI�g����,����6K�]��y`=�lI���:�#�h�v�rPnb�U#\�=݂+��tuJ[�0:�m��A�Z:���9.�f���K�/�Xx	�Y�bK;78@-�&�E��w>���#Aԓ2��R��h�����x�ek��^L]�$�Z�;�t��=�[��A|N��|�h������ ��o�-�ak��3D�r���gf?-�IA"�T���kX�Ǭ=�q�C���������)�,7P|v{WS�Od��y�_�0-�Is�$�4��ܩGh]�y;�E��zfk��D�T=f���
��̸����V-\�rX���9���Ʒ�������n&6�"�}���.�9�;f?p}<�Y0�:D�A���1����+�{l�b��������Q�g��ڑ��j�s����|x=�.�:'ku��hn�7<z�X�Q���b���<\��-lҙ���5�w=G�mV�`�p��*�K��ŗ�27<����7���X��9�c&㓮��,[�2���Q{R�"Y��K�ʥg!�_t(r�F��t�E��t��(>�o�m"{٪�p ����Gf��f'ZW:'��x ��	�����4�q��b�i�qR�����y�7��4�Ì;��*���} ��(�h�d���rG9k�b��bJe����x�%b�[i<4�֐w��-gzB��uߥ���庼���w"X̧�t�i�|,��5����ʰ�k��p㰺��#|:�Q���r��v�}U�@� �R��9��#��E^�
��0d���/f^���6�x�eAk0��GG8�nV2��I�w��lH��Om`�({���7�J�2��R>+�:��`�^P��ۼ"�h�U��)۔j��c%�^���'��$�l��Iޱ�3̲;�)F���ar̹�\۸�W���B�Vg���ͤo�2��P�(ȷf��Z�<[��th�]�׳��[�4�lP̊������/�oo�%h������X)S6o���=�(��m�R�h�X갢`rZ��w�a����^^���/zs���.��r���8����FZ��\�V���ŋ;IYؑ�[�
WIA��vS^8��Z��xgp��2�tNx���t_W��t�4�۩S&��z̠�xk�n
Ue��`�4��Y��&μ]��l.��Z
�P�D��w$_&[쵈L<+�_�J9�TΜ�r)���+����ڣ���Ƙ><Uep(�͑��a�I�ֈ���7;13᪖m/A���4q��v�ھ/Q����W���C-pe�@C��=�\:�p�mi�2�ޓe'�Anש��w��[���]�s��*y�U�/�&�Q��	�2�z�|t}��N�sfZ,��a��<w���4��È2R�w������-��pA���1=�=ҶK@����ůcm`Q��sw�Ky%�(+8��us��NC�:;���%#p���1�_�#{�3���XF���r]�k9rW�P���1]<�3�+�9��wb�$X;nt���WL`@��敔����.-���W�M�a�s���Iܧ��[B�S�P�=q����E��"
c�\��9���_=^��S��c���K^�Ak�oHx�k0���T�H��b��.V���q����M�U`�-�Ɍ:ۙ��O��v������]1�_cw�ۖy禮5�6���G-�{�6�������޷�Aپ�f�-ݎu��+����Q�[�e8��x��sS�.�ng��|	����uAkR�>*� *Mi�l����sL
����Y�c��wc�F�7y0w´�|�٠�јE�H�mQ��>UƷ֝G�f
/�[�=RclWZ<�lWUY4g�uC�o��A�RODS�H�zD�3t-��׉��'*	�s�z��UF(ݲ�m �j�*Q
�J�	���	��WT����)^ɶju�JE��0�8��fm�7}kZ�с*ŋ�����Uznl��Q�3v=L�|�ڙ�#�{Cdٷ`V-`JS fU�:�w�q�N�饓y��v�bS�j��j��}�щp�P���۝F��K���*k4�I�;Yȗ��5R�-�3u'�gj��;�������h���NqT�@��ӯw��-�j�܇�F�&n���p�u��-�����W�O�px:̠�@��\�hC��͈RHj������x�݉j|Za`��5!�����՞_WՐPU�q��Nh���V���u���K
ȋݢ�60�*�rN�q0z�d�{E��X��*Ь�Օx�=w��\Šsq"�M[�GDL�`��mmQ�>{n�x|]�`���t�"�l���P
�vt��<��zX�]�����r�_���Or�b��'H�8��f��GZbP�}����t��6�N���OM��s��x��O,�=���=}+�,��7�9^�.���khK[���U�8�����ˊ�W^�Uߺ]-�gS�gw�����9��{{b̎�]�|9ڍ2VQ�8��X�@�(����d�tr�G�K��b}��3�����y�-��W$���([��W���}#�h�m5�/���3�ߵW3O��EJm8�.��ؽm" ��iE�.��9�n���\6�y\�T��}���Ƙ�QF�[��"�$�Eofq��]M����a���%�7�^�=#�D�4E�fh���hT��q�gdI��|�U
�6x+k�_ۡT�f�a�\o�D9!�Bp���_��Vȟq�i$�s��ĺJ�R��س�"���5��1Zg69��B�g;�8��נ_n�mrTK�}U��
�م�e�g������R�Mv�8y�/ #B�y��:哞q�6�D�K��'���[�(b����hG�{�Nn�r.���)��_^�����Sba��r�K�8\6>O�<	��5�׽��ӑV��WB�*�دc2&�c"�9gM�!�;`ԣ[ά��g\��ZPr�{%���oC�P|��#�fѝ����u�n�#���=�M�߻���؞�볢�J<�%���]`�'���P�4Y>��W��N�evy�M����bP��cY=�P���l�48�M���:���W4ԁWu�ҳ��ؙ�w���+ՠ��^Hy]]��t��`�����2eRw����m]Fm�u��B�w�1��xmr^g�y��B�w��I�o2���X�Ŋ�kՙ��-��^k�u^�4޺V+���h����*\�f;'r�a�mo�������.8 �K+���>h���	�0�I/�gm-	���W7�1dc�R����-jl�c.���:�3����1wNl��p�嗇z����Y;˱<~�W���-q43�4'��^� ��y�d�W��6�eN�P�W����u�y����C�3�˔X��6��(��մ�h3�(����P�^zV�<BڮT�aT5N�|��g9�^�WFn�jm��u��Ws��[y�k��R��6'J��Cf������ˉ�[���ֺ���R�o�����;�����v�(�X<�Y�R�s|5}̑d܎{ҵ��=����3�֩���3˯��u{��P�73�>�y�t%�/��8�j���UJ�޻������R�57��Œ����O�DLΞ~�Ť;�/�k�T5��U����<�=��yP��ɔ&ƻXD�G�	��~���eH�9�����jH�E��KS<#|��!��D�J{P�KtL�g�	��7+(<ڸr��S�X�k*Q�y3[	U��7�*tl����ۑ	���9z�oW-����βs���:K�7��H)7���Z;67Z��(�`�iT�:v`]58l��V�j;�\�vz�ᓻ\ޮ�h;��Wl�ɑ8m�XX�C�uwrp�Z�{�Nϝ򃬼�V���;k��*��0=�����Y���:�QNG7R��N�x��.�Ff�(���K'­cShz���{�_��>�#<(қ�j[���Tdiy�$��tV�[3+�9:�i�	��Q�P�ag"�]�U*$0��!+�����C+�̨n�|눟F�^����˾)
���g2%��1��'2wL������p[���8�w��h��O�LU�`�0���|�g:9M܏��
.�	[ۢ�^��p+moq޺wt�ot��|6p�S:�e���I��l+�I=b�����
�9k�V�n���yҴ��'{O���f9��*�)�ci����ڙwW,S+=:F����r^�ObN�͊�I����|��Ӝ
u'�)����3�"K�_x9�Arm�3l�a9wK>�c��3z��ݭ��{{��^��K��Ytn4�ӨX2��O:"���e��f˩����^[)z��%����#]q3l��>�7׹f±�:3�5h�{8m��#jq*��`*W=Vx�N�C+7�]t�񢲵M�Z�����h����k4l��aə�Y0�4�'��;�r�|�K��Yk�c���J�e��&�#)N�Gs��V.��M�Z�ũ:�r����|/o�1g���܅N���P�2iJ�Vy�ۤ����򜅝��o?���0�r�wf
Y��]����*`K�W�Ck ��l�L�MX�Rb"�Xe�u,I�����:�%ӹ/���Nk�q�@WֱT�7B�6B}�M��\�3d݆�9v�[����5���}�=���#����Gq�rhEB��}X��6�Ü2fZU�̾�ޔ��(�
��+i}G���N#�f��ڱ<���R�8#��&M<R]Y\;�/{�+�+�mdF�wmƕ.[��L"T�ɎA�FN�f�︧�u�ޛ�M�\՞�Q�8�D�Y:���쳡��JS�`Hm!2KUeeKS��7Zz��a��|��l:GT=��θ�(�B>�����*>����6����;C�"�vI�|��T����}8�#��J�0�`�>�(,I��IT�ŇX5��z���d';픣5y�<�������og��lVC�kFոB�������m�B9��Ȕfb\�)t�6;p�e;����u䠱6:.�����`{zS�2d���B�`��GE��8ŽS!�Φ�&�]b��$%�'q��Uϻ��wŅ���Ӡ��ŏD1^D�<E�K�j������pz�}{V,�Ȧ��.�H� �ܽ��4��]�u(��j%~��o�/��yosX�Ffc:�o�eJ�UDEH�1V�+F3�Z
��DīTD��P�b
�*�-.P���FE�1DL�EjUAq��&R�R+�.ZT��V
�TX�X*���Y��Qb���jDC0�&[FFV��b�UR"AkH��"��UB�TT������*�5���`�1c1��Ub,Kj(娢*9B���DEX�2Щ�\j26�b�\�G2�E�"�V,Q��U���0[kB�dEƊ�2�Y���&R����+V�,b��j*��DPX6�TB�j[q��dQDEFah5*���)��#+c��5�T��<�[�\Rʎ㾏:��vi98�"�����wL_u��X�n���/0�vqμ/y����Gg^$�H{��Yx�����ij���a2�u�r�U���o��yb߻�Ncѻ��M�f�;�č盺aQ���]=yu��㩮֕Vso���{����U��g6+ܱ鶎c��q�M��Ć1��{9=���q?lysQ6���3����X��y�BD5�Yz(bn�>ٗJ.��*��9���w����/����u�����ۜ�KA�q83SD�̮�1��+��z&������Q;<+ݍ��]�Xz��t����ХO9-��>��9��n�6֎�iBq�(ݬ�&�Nk]{ʲQ����rR�wm���ov�\�T�,6:��Y�bY.X˜�O)�XA���֍�睧��:���aۜk���WIu�Y�/���~��ܕ�;o�M_3|�jw�A�Qn�(��Yc��oJ���V�M8tv�z�C�vu�ӄ�6���n�l�t;��R�޴H�#/BN�����.�So%������$�F�+��MƖ�sc7�祈m=�/m��M�}��#�r�wa{Rґ:E@���:v�����9���ɇ�v��s&ՙ�^���������Ζt�ts�3N���U��Đ�V�b��� ��9��[�%�xS���,�YZ������F8�5W�^O$�:�Vw=��}rLs������2��2�0R/��n�;���`�t��8�T>Z�}	eT6�V��p'Y<���Ux�c�ś�6��T"��T�-u����+�-�����MM�q�F��h���9S3f��9m�+4���6��J���:�{)�2BwO$�2]Ƌ�;rU�M�3���T���+g�Y"��N#63����a��T���R�	N���|8d��4��є�h��]@�w�/��{F�ƫ퍴�-P��ż�6ǳ��`Y�O��a!�t�ڢ�ӽ5��bf׌�E����gki^�k1��}���y��'RVG^7�L����i�G2��Wf"=k�o�o��}Cʽ `��Y+["����uB�6HY��{S��L��B��Hێ("�]�p˶���{���m�1:3�E�y��R�$ʓ�jac/jR<1v�3�ۛ�����3���l_v��F��3&��ԍn+�o���QY�0�=�
�v���kϯ��[�=�{��}<��4\��)/e:؀'9�ٛ�>ޞ����:y���_�3*��X�swA��������^T N�o�<���c�X�h��jξ�W:��棝Ex�1�Mqi%��M���8_z]�)���_ti�H���^����Ͱ5�۠��{{�b:�	s��}>�����y����auؾn�����u�c:�;"|�(W��ګ�r��V���X��B����y��n`�O���j���K޻mH�DM.:k�R܉��X.&���C�WXJN1X�w�!^���������+$��A��ly�ɽT��0U>�
�S�M���]n�*F�,6�"��io�}����d�����#�#��]�>���z�e�C'�N�q8r9+/�w�;�b��^�Z�"U���/��c�����.��F��t�u��/Gd��IW$^u�f���N�mJ���1faȡ�9��������΢X��n�:�j���$6�+�#�k������,'tq�˓r^M�B]¸0��ZT$jN �<�2�%���^r�nHo�9��Ԯ&G��f?Mu��'�υy��5�7R�cF�'�.UȦ�C��Y�8��t�ֻXg8�_:���,���}�)�׬B��+=���Ż���H�6���u}^���z�O��s��ee���h׳AnlN1�f2{��_.$�>C��P���[b^Me1W�
�-q43�4�=�Y�D��Q&�Nb�f[$םn&���A��ŉ1�
�L�r�r�Γ:-j���CȻɂ\��^�y{��^Svr��mW�/OP�o��F�s�yG]�`�Z_�(Ws�K/Ϳ6�T��(�~lN�y46�����K�t�;ػ7���c.�6�P�[؃��z��^
)B�y.�sd��/v. ��x�t�j��b;���y~Ħ�H���&yu�Ց�k��~��t��WwU
�צ�����f�y�T��poj�]�R��@�����:����(B�SlmA{.���:��~f�"$����_^t/���641m��i��%��#WG^7:`#�^9�2is�E�&5T���e�Rq���vv��9g:���� fH���Q�wx���UzV��������1z4:y��������-=ABZB��Mk�;Xy��n����a������Y;�:8 �]CR�&xЙ]���V�v��.�c��:[R�b����BUB����d��ȿ7D��x���V�+�T�1m3��eY��w�= ��[��:T�b�KTL����i�ܗ��+��6nn·��^���S����ø�Б�N�ߊ�n���܃�5^a*8M���ݜQ�}የZ��P�M�����k���|�c�I�a��U��Н��h
s\u��2z��3C�=7v�n̸��"�R��I9���ewz>���]˫}��{RS�QT'L��A�n2�P+�U"��e��k��k��X�y�S���ck*�r72�yn����[B��}ˏNʘ�˜�y���� �V�PO>V��o{+p���m�\=$�o�n�d>E��轩���J�R�uv��gtv�EJG.�]�&�f�����Nc���H:��k�8N�{���¹e�W�2��ɡ�f�2t��p���T�n�긯�&w�>�Wz;��F�<Z4"�yJt����serLFnj��Rf���,	݄��`v�mU���ب�D>(P=���k�؉S��|�-�[8=��lq�o�x��s�[�L�m7��w$�^遬6Z�]��Ó~��*���2g��ӽ9z�5�h�Y���Uf�64e{�V�Y���U�:��������޻��_+��6����_t�"���..;�N�����/E�!�xhp���+�ֻ�Gj����t���6�ۨt��a����"�Q��o��i2�v_�,�eL���	���1H�Ɠ�[)�z��^��eN|D�"��,�>�����q�l��M���g1�k�Sʭ9�Ǌ���2�y�1m��4�d���P{/W*��h�I�+O=���
�t-�6�"@��z����Kԇ��k�k1)��ۥk`�p�Z����5�+J����9M����9}6��G�}kNʌ�8�O�G;Td�k����Ӄ+FM���h�Y�}ܮwtx�/]�����b��� :�q�\�X�C��S�I�Rl�4'�]0�w�{|{I�H�hV`���<�U�/�rVϪ�E]���1�d�2�fi���ڔ�U�fB��� �Д�M&��j�Җ���{a]�58�u�hP.��^k�c���%�*�Þ��=N��S���\�y��Z�����r5��q#^Y�w}��/��J�+#�Ң���c��<�ِ���tXum��sz���b�ݿ7�A���f3�⟬���!���{ui������o,6�Xt�,].􎛞�6H[wk6*[��έ<WeyP�'S;Fw>�qM�s˶s]^��#��a֘č���qv74��E�
���خ�\o��K�ӷ�*H@˜��;�X��.���g��6�r�Y�g۾ik���޸׷Ֆ˷Ы�&ʵ���ϲK�D�jo�_����;"[e
��e��wW,��Tb���+]D*��u}G�e �pڵ����+��a�/x�ʡ��$��=�G���mV�f�w���Q���m�ڛnl}����;6.�Qyp���;�y�*c���+�f��	�Ύ7]�A0μ��e���B>7�N(���q���N^�����S�y��mH�DM.:Y)T����LԠ�t�������%��\�nyj��M݁�M�	g19��ĻupX����*�r�Lp�^-�p���;Θ޾�(}�Л�� ְ��P*ɟ.G����+$]gU��v\�OX��}�!'9+�w��*H;e�j�:�`�%��=nf�B��U���=����~F����r��K�x�����,n��}�$�bs.0tk��u���L��\it��S��N�}��ב��{o�\�鶎O�����s7�0JM^�.��=fzU�9:��Ȭ��R���b�s�����>�{��y5��N�^�\�� �˹�b�ί(�ە�YHP�hP��泒*��=��D� �|�Wn) �~�yA2�"�%u�����~�ߢ�S���+׊/W!�A5���@4����3%ؼ�;�-<�_O�KZ�莍]tVY�ے���f@�)]<9��7E���zh�п{
�˭=%S��
E�ϱN�����}�J��땮HHO��;Ls��1�Y�����u2i���l��2���+/����!2���XgIC���]n;{�^W����mW�/�"����_$z�N\�\
�>�d�\���ƹ��ۼ^m��Uj�R�lFo�OdH�{n����� �F%��;�����_9�P�[��A�߆��۠��!}	t<�u�31-�]Y̓˶���L��c3|�b]Z��޴�.�c:���`�s��问b���5��q��V�t�+j��wc'�<��M�{��jb����{7���x�+"��m�Y5�Mk�k<�Cu�m2�
��7ú�+T�V˱��7de&xׄ��Y S*��by��D��\��G��Ѻe��T�7�C�!�&C�x�>��{�Ω��%o�[��a�wɕ�6A�K��}y��rҦ�/�H��ji�[�1��y���x�_dD�N7����'R�6�
�t��[���v� 1�a������n������S[N782�Y�6olx�^.�K����vHJu�J!*�>b���;u��)�
L�F��<t��5r�NbrcǪ�{VD��vjq��q'�.��<�S8�4f�3d鸪DMS;b��*�$��q��^��t��a�o��"���ʫL� `��rǦ�9���؂�Zڔ�6k(�0�Pu�U�}���xz>����Ť��PO�X�8�oQc^m.��{�'���z�l�C��4���e��v��<�{6u9<�*`g$i�̾{����gD���w��LO_Q���*�u租�v�7v�0��M���]�m�F�<�ѽG�l�\w�Lg^7��JR�B��\�ڧ����i�`v�T��+Q�̎ꢷ�S�z��)�w#4�,~�:١|�=����R�"��������n�%���o�k�f��W叺^�U�V��|����x��U�jr�cv�ګƟ��}5 G>��6Ď_ܮ.j�֗bո��=��u��onQ\d;G	�n�QvȮ��y+5�J��Zge���5�~}�]�$ I?���$�����$�XB���$�؄��$��$�	'���$�؄��$��@�$��H@��	!I�`IN@�$����$�@�$����$��$�	'�$ I?�	!I��IN��$���$��b��L���H�)� � ���fO� ė}L�E��@H$�$�Qm��Tklh����l
$����!Z4l�m6�)F٠�
�*�-��"U��	J�%YKEcljT�����+*��*�k&ن��lh���&�֥[Z�1U��L�1�U�����Zm��o����Ɩfi�Z���k b�7n��ˣm�&��m�d��+m�Rh��Y��ј��6��V�a�j��4���f�����5m�f����ff[-�(Ҷ��5���mPֆ��;���[iC[�   �p�.�RD��\m����\��)t�;b�KmU���a�vҦ��)]��u�r�j���6�5T�m�Eu�
��t�la���Siq6l5�лFY���ͫl�x   7�"^��)�vei�+]�q����͎�Ӷۮ���wm����m���l���qm�
ڶ�s���:���\�J�hm�t9�7
(r4�q =�6�6�
Y�Q�  ׸t�B�
(^�gxz44CCC����
(z(PС�80hC@ h����(P�4(P��Н�� P =
$���[2�ƶNM�i�٨��jUZ���k�����,ⓋJ�H��6��lx   3�V�oe��n��m+�sSnn�vvƭh��ʫ�]m5.��Zj�*���PV��ˎ��*���uJR�n4��T֥*����V���t�Ҳ�h$�����ֳM   =�lkU*�Nٷ.ڤ�U�8�m5�K�.�ճU���R+��һ,wL�[�l�9aҩ*t�ZCVڪ[6����Jl*�J�%]�:"[5-�E�0E34��<   �ORR��=N:�v[T��κնk�*��p��XʖQ���fe;3���T��v���ԥ6�m�I�]��QV����wsm�2�]h֑U(�a*��  ����P�wC�Q3�  nٕC��V��U���hH��F� 몡!j�nU�t�	��lјj	P��  G�i@�Wtj�I:X+CZn��T ��p4 �M�GUn��P(�t�Ъ�CU�ڰ� ���Qf��m������m�fF�  ��(#S �wK� ]p(Lk )�`��F����.��P�ӆ��ڎ�����I��ZԪ��Vٞ   ��Q[�b�bUՈ5ۧX	�ctΨTж�\��wj�UӲ.u@*R�뺊�V�ڵ��v�@4��'m��*�*�U��b���4RU#@24Ѧ�S����i� #L"��)�R�#@T� JRH� �x�4�d  	4�eR�i��C�+��B"�2|�BG��j�U"(Ͷ���q�s�Ԏo0����Uh��	!I�! ����B��`IO���$`B!!����g�kD��F��?������v��,N��aF�1�q/�/9wD>�{

K+,�*��/n<��R��2�޽kv��Qx=�L8��^m�n�4�ݍ:�Um�Ecf;��(��á*X����-2C6F��m��b`%7����D����`�ݫ��\�Wu�Խ��bT��հ��G�P�ٰL6@�LlJ�L���ާO�܉u$���F}��� x�t�9J�]ij�3+^)��Pp*���35��! )4"׈���)� �oi�(e�_�Lr�[��SmP{0G@�ȹV8͢C��3oB��3������*��7#zQs2dbͽQ�UL�]ɓ��5-
f�{O^�n�k6��ަԧ��`Ğ�afrM/7���z�ܚFܖ��sT�Z+3P�N�5vѓN������2�JS�u3`���#&|}��v��W.���I�p��I���31�,�6�ʒ݃�n���AdTJ��óI�z�<;[4eI�nY0m�i��0-9�0���vbl���py��K_��1��8�Յ*Y��B�ًM팀ڣY�3$&�Vӫ��� i�%(Jsm�e
פ��e�R�a*�Z���������Q�oe<�L���;�4Rܸp`A�!Ȓ9�Y���zJ:wV�T0j&bf�N����hX�IܺυMu22��֩�R��-�v�s�z�Ā��k�����GU;ͽ|5C`ȯZ�@�n��P��E֩xNYC
��e-�R(ʒ�ķF��f�R��b�LzSR���V�]GM��u�̫���N�#t5�IEF�+~9�XeR�𧦵��O �a黻�4Q�ռ�Rk(,���<9O[vZ��
`1'v6k�q,���xt�i��-��t��w�Fݐ�pjP.��S�6b92-���H��4eʨ�e�u.3tJIC���]j�{�O>.X4ʤ�����V۬4��:��RǶ�˙�ȅe�e�ȇ�[���E�R�tn�U���<w{��F�3,�Bݕ��G>{dݦ�T�Z�2��f�E��j�U�R�.��i�l��V
�p����I̴�V��e�	n�&i׻���j31�F��`J�
Sae���z-!�ˢ��}�n�L�\�L
Yb�դ�OVFcv�F�lLA��[�AJ�,���ˤu:C.8e�ǺƝ̖��)���dUT���U1b���h[5�a2:s�2�)M��:q}���a�.9�h��Iak�R`��3��e�@�qD�i�Uio��wR�H�kLo\ض�\1�-R��s �ѡ"�J�m�#V�r9%�ԅ$�ݬ�Q�-�Yӗb�p�3J8��:0]�w	�ݒ��x�p��e$�,L¢�z	q��R�ɗf|�Ab��ױ��Qy�JX���$Z�b���蔶0�g�*��W#F��K��*y���U6��XІ�I���^�sJD��j�s]U�q�yDd-���4���1�k1S^�<O�w�� doT�>���l--��%ش�U��ZZ��ӐMT6M,�Kne��_Ү�K�DL	K�;���P��$x�CS����s+)�rl���e�I�di7��HZ�Pդ�������b�-Z8�87��$Ҁ]��������?	FL���U)���]�p\�wwZ��Y�i|��y
3N���dيjo&dutk�$�M��V �Y�����s`�R���-�m�L��~Ն��:qf䳯�ܷ�0ݍh�	�r�xr�ޞ'�I�&t�����]�Bm̺�욼$,Oc+
id���6)н!��Z�1WH3wtV鴞"k&��50�oH���; �!8�Κ�K�4���Ҥi��5�Ê���K/ej�o%&T
^$Q�-�Щ�q��;QK�b|#&ud�c�y�A��L=x#[X+v�W��ӥ�[lj[�Onƫ��J�v�L�:V��v*I��0����m+�����b"�Q��5(����X1�2�{!|<47��x��x|��&��2�K��J�*����J#�7�Y�%��Z�JhT�ih�&-��Ŕ@Y5�{�mL�oEو�W�쭟�9R#�F(A�6�Z,�w�]IM�ugr�iV�x~��^+�r�"�h))�:u�Z��� �{���)�֢�{BCr��em������G.�Ji#�K���"�uh�	]ܘi�2� A1Xmnf�F=r����m�,��t�,Z@��rn`���S,�$�uϭia*���"a���氙��tD�&%��%�ΕL�e��C�c�[�t�wh�:��� �����c����x�&1�Dg�a���SSQݘrn�G�(Z�g,#=8��)���w�܇�#� $����h�Rȯ"��u�S!oIѷA��;:бp��oX٘���ID%F�4���>V z�8_�e�F���uq�(	r���ò�Y�2GnP��c2�)��CZ�SVh؛����F�R ���SS$�U�&[-�(��(��Ǩ㙴B���ДFͥOA�0;��j���j��r��q��)� ��yY�)'��xY�a�R#{�*�m��n��"l/�G5��Hj�3m�V��`</0\�!Y�,�HZN6��Akj�v��J�T7�ix0��`I��&/dm>�٠�4�ln�m��SD���L�ub���(�Mڨ�Jӫ6���Tx�v\$kU��yu�����U��[Z�Z&��6H���̻��(U��l�c&]����˩��5�e���-̓uL��?\�k���s$����VùN�����hhG�0 ���0C�1
�����?�5h1l`�@)�LFN���JA���f��ec��*Y�4���mXM�;GM R�R�X݈_۰�~ŕ*=���v`ۡ�`a+�M�ؙW/^!sMm-#���5�5�L������&���1!X�\�/Brk�GS3!��5��\�k�l��{��������#a��'��mPh�$�27�N�i7l�ne�I�*cn��5T� �/�\�U��F؛b?�o^R*�2V��p�����l�%U���DAZIz�<�����
���)�x�X�U]8��f�2�-��Z�����J�ı�Ѫ��.Y{���j��o�����6ڡ ����u
݉V���/�,L�X�գ5��m�.��t����YkmA�Vu��r2��:Vڼ�[e�*#�
de*ip�1�*c��֝2��E}���j�U'0,1�y���졐����6����a#��(k��1	���ؖ�l����˒*��'�	j�vjk���=�87�sR�9��XB�&�&�薺��5I�����	3E��)M�i�	_n�2������n�úɁ�&� Q%��o�JОs��Gq䦉	:�Z`P!�b�
0'v��V�l���c`{\ ,��&��;��q�j�	�k}���I��ω\q��ln�ٚ��D�jƁP�����W��i�Yb¬e�k5*s^���{c��������%��I�SE�F�]�J�b�mc�e�N]bO;#�{���L��h���Y�H9��^�M�O\w<m8�dVJH����&��R٤</s#wk*��&�ݧF���;�[8�v�e5�h�2�A)��W�t���y�*V�xV`�ԓ/n��� s�o���	ݓp�q ���{��͗�bƪ��J��l�{+G��8��#�L����]�c�y���Mj�h�1���v���+b'.R�)#�7"�\�
���me
,id�IN��v����>Ŭq�QD���?U8=}�v!��� ���Q���X�R�m'�u6H�����g7��f��"]1xx��7$Y4� �"���z�AWRf�.����i$��2mhđ̔��pˋB�/Dj��0kÂ�;����P�̽T�P�Fx����W�i�E� ��>F���u#k\úJ�B	/.V�ֵN����Z� Z��;��[�j�k�!�4��̨/s&��ISb%%���H���z4��d����q�v�90�%��b)Z`+%I�8��3te��X���,��m���`��v�k�V�&��I�QJ�������<�S��,Å�$2�H�dK�wg���˵�Y��:�E���`�t��g>����Ge����c�w��p��Cw-�wi�.]�q;�L�BRK���	/�2�o�(�!�Z�J�e��^�z/(V��fB��OZݨiњ�8cݡ�Q9Z/��5S1�M�{��C~9��륂�������*�z�L�勶&�5ZPQ��]��P��j��u�9�:hn�@g���8�[���bU��$-;{���ʼiY2�nm*���/%��k2��40���w�>6h=Ô� F�X@�[S]�D�eI��ge�n��I�HcR��9�'J�{i�t�R��&M��0�����s�L�ˏ{���#�2�t�Ӷ[�m�!�,\����t�ܴ�jF[��sD̔���K ��� �Vƕt>*���(�6A�=�u@��pE�8|�rfa�V�Ү-Kf��Z�7b�R����V��7+[-|Bg]��/S�C��	�3ZʺR�;��se��s�Z�6,�F�j�<7��<:")Ђ�ı�/S��@;6\�G����4��t�������p�F�Yl*7u�������V�����Y��f���!�;��;�T&�2-�'؃W"��*9J0i�ہf��(�uV�4�\��<� ȵ�h/�[a��:��rV��J�Õje��6yn��\X������m�T3,K����i�7̼�.U�[-�hn�7���4Щk�]�p�wA�Қ�ÐH�f6M���[{xV�Y���Z���ѣCV��K�`ג�A�`�Bڛڻ�3e�()��Ih��$Ä���]����f��5��z§�+8XB��x�+dɚNj*t�p�uq!�ݚm'����Ҽ�����s3R̘�ݫۀ�c�n�jY��S��l-[���ûB#b�K�3kBx�+U��p�AU�k(��Qch+����1��8j�b'�-�+��%&D�x�ٓh�qɵV��V��V�²��n�����tV��8-�&�Y<�\��sq+8���򜷣������ͣ�ʠ���[kDu��n�U�'�4�M�&�-�F�3�ۚ��C�Id�tLm iBm����ie���@�-O�|����;�:8���]�y2�OB5V���v6=IIpi�.a����d��v�4�������%z��k2<#$�%[[$���;��oN�ɧ(Ҍ�4�O"�P��Z��B\qd.�[P�vr�ձZ��.���6��$Q�pa��ś[��YTh(D_Y�%�n�wQёA�&Pd��V��HJ�5*�J���JSڗyx��6��G��A�ڇ&$`���l�Ɇ�J��:����V5��q<��L�#ܲ*ŹÀ�-���b�b��ѻ�Y��=:	�q8�$YB����J�5�4I�t������L��U����sk)2t�L������5H�ƙE�
X>_+�9nm�f�!�~'%��[�ћ�q�:��m�����ĩ�(�s\7W6H[�4��t�ئ��.5�e���!�gD�$�G&<�����ɹ+nJ�W��*��yo,�T�lb�%;��T9n�\��4T��#��U��(��olk@ݓ��3.�����AȰ��"JL��U�=>x��A�t}�=���QP7Om��.���nS+^=z��	N�V]:PTR^�4e�wM���g�P������;H[0��t�V�����jL#�A�,lk����c���2�4ܤ��3t�	����#	��3Р��rH!��}�ws��L��am��k.'�e%�uUiG��T�{f�H.��	nL4�.[�eM��+6S�i���BIu�)�
U���c�F�*�h�6E@�*`�w�A��Z�R�M�1aq�_Mt1�Ōۭ��KNbt[T4���i��t&�&�86�����ڶ�1����{Uz�*U���)�Bl�p,��&��I��cr⚴��;�j��*.�����bYy��d�e'ld��.Ff+��Pn�����̖�X�a�'E�Mb���e�M^Ih!i\����0kQC�u5�,�٭�.��F�ܷ�8�	SmB�i1̂��Y�;*2@кw�[.B�6k�5�)Ve�I�SYT6Ȱ
B��8�۷��%�T�F½��DʐT���h��mK�l����'ȭ��dK��̭���ԡ����Ŗ7E=)� ��V�>�f��դ,��6[9c��m�ʺj1�F�Ɍ�/p�"�e������IGV�����0(��W�4a��eش݋��ۉ�`-�;�v��
����������.�<{���U�Ë�-EuUPe�ݲ�b�r�p`wF�����3�:��G�0"qg��#��9g��=�F��+��O?c,�9���ܣB{N[Ү���G>�B�)��y�dk�. f�H���cd��� �������7� 7ڽO-%�Jl������gV���&�W��*�v�2�6�Hܠ���$
�
��M�ia��FV�V+8.�Mb"��۷�Q�7vT��aѱ�L��Ua-����z5FmU�3p,�Ȓ�b];T�U2�Z��t�Hd/X��X�B�&˹zkM<QѬP+��N���pj��@����m��.Y��H��||�aqd�9�Bo��xx����9n,���3}�j�eT�+%w�D���PeK\)�b䫀����{���]}o��Rx�1z/�1�Iy��D��e+|�k~y\nQ�ٹ��=�.�}sǆ[�~�m��詢W�1j�W^�2��qv��F�{�����0��vơ�J��\�&G"v�o���6�O.���0�\���ArĘ���;q��F�#ܥ��/:�xӝ��W�_M�]����Iq!�X���r{�\�8]��_�hi�J�\�S�j��]w�ߐ�,� h���^���Y�e}{-W�//V�;'��U��H籣�^����}{yY�۰����D傀��k�4��f�scΚ4������77_Y"�����j7u�3�er��>Q
���+��]�aZW��(�<���m�G����m�p�����@ut9sfԾ��k�q�8�WX^���Y���/g7��J���;ݮ	p�l�k�'�uۧ���+��y{��5�c��{7U
�y������3�W��UD!#�*醍;��)��8��%m<�ٲ�8��!�e���R�w/H
E>�ay\(�n���P&�Tѱ��==���FŢj� ���:���o��&�a*�{��Ͻ�칼e�x�v����Q�}4�����嫍��Fo�^��qZ��w}.A�}ώ��'���Y��5L�dv|��}���6]?dX��6��h����T2�$��z|p(4b܉l�]��y�SbX��kbEu�W���LwXb�D��~S�Ų�'�lC��d�o�f�.kh4��0�����ի��N�NM9�Q�9W
�v��ti[�q�8Ї�o���9�o�����b�sz��y�#��a��:~VLM��g���>{����[�2ȼ���LG��g�a�OouXǬ-*�k���}w}{�zbB<�{�9^v���j�r4���
��D�6oL���2�Ӧޑ� ^�@�3ts��(WVD����Φ�yi����A�G�8|!�����0r�u��^� ����34�S��.�{�;|M�څ�Z�\�Wd�\R�Ǝ�w-�Z�q��#��v�&?q��&��^��W��YҴB�i�ݻ�/z�q;�b�:���h�ȵ�*�X$�,��v�ã2��4�'���k.�l5��8��S����*%LGP�����j�a�;Y`h���U{�c)��NԻFw�]~���+k�n6}lk�^t�� ��v(m��:՝$����V��qu��>�	�ϸ@i@��g����qn��{%��Λ��
�#�)T�[kv�h�pHnmkoe:\�$�^[���������gn� X�w0�dp��x���ғ"�M��O{<�$,�ϊ�v͖�}���ϵ��t�N�s��]g0����W���Y|�Tt=�7^鯍"��N�j�m�Ie�ź&+y����ʉ�R0(%v�U�Նr�d�G6�;S�^Jw��ƨ���:�j�,U�K�/J����\��sχ��E��p��\�0U��_8��蛧+�Y�Xw���u��/+�9�U�Jڀ��<D�.��8�rR[��A�mRs,��9kU�FI�K�}�Js�f7X�:�p������hL6.�b�	`+�[�ug�|��з'<�C5��&E���Hҹ���#� w$�E����O���%�`��ž�5�#�	�y��,\<3��*��5"�����wp�=�9��8NX�J�2�����;��T�~K���G�wuR�s�����3�_b��M�d}^t�$�|��s���m��wt�,<�G3���ɣ��ܡ�Ҷn�n(q��"0��������p|'_t䳔 �m�p��2{�}��r]B��G���z�ǜl>��g+Jv_%�H�WU39�E�7c�\���%�K��F]:��w]��ã�R�C�J�x!jHY���?�Ӕ�Lմx��:������>�0�/3���mu�]M��Go���-��6�f�v�ꕏ��%`T���Yz��NhC�*f�$�df��.���;�u�&�;���m�ޏ��+��I�y��g���\��ye���>��M��5�[m�������T�ǆ�vk��/J}C�v_^۶�/�M�z����=������yz&�M�,�Vj�����K򢃴�a\I>J����e������֌�	��{����y�P�B�fo[̌{0kwC�F#�-#y�I�T�%.���.�K�#�h��i�2Us����_�
���T��xV�#�y�U��̎D�
��,�min�%3���z��x�Y[����;z�6�^�3J��|oG��0�p��(����K�O�Ep���yB��S{$��s^�L��rU���S���l�櫏n�p��/�i���K� �f�9m.���-�NVnM��}�˴�_��f>�I���
e}얮zM:���#{t;��ram`i7"R�D�w*�k�s�5�����Gm�t�I��TUsIS��Gݞ����E�g�!�߀H�GvG��{���A�j�}��L.h�f��ޥ<Q�,a-**���i5�����W��3���g�̥����L��v��+*PH?���V��:c`��|���v��m��B�*;����t�u�1\�Po]͖͠�t0��BW��QK:���HX;p�j�sg;8N��*���ȿb�jZ�K�$ɇ�|����c[���נ��U�K\,%�Ҩ��z���AX�����4;E���]��nY����Cݷw�<���H)g�Y0)4*oLT��5wں��k�kTW��������=e{̡�d��M!yk��N�+��XZB��XI�c����O#�]�*Ю�o�3j#�.�3/gV��﷋��Ni�:U��l���C��mx��8��N�F���Q�|�
em�ړ�F���8�6|�d��K�Cs}ٳ%��&
���Fٽj�2#W`��-ᐹ�%*�qH݂氶���FT������:54�^���$���j[�D^�W��˯<��<��M]����*�	;5�z�:
giVy��N�f�OJ{��F�\Pd��F�Ⱥ�i���}{����r�k]jT%/xM�p'�,��wP�q��y��*�.}n�׳�q�R�䳪l<zgBP�@nm�ϻ�Z_2�̛�b����\�W�ZV^KӗC繍��4vS��6'�+�V_�WҮ[[{]bAQ5�:���U�Z��p?����r�r��ǹ��8�5�,wkՔ��U��u<�'"���{<oW�����뭧�c��P�!�ݭ+�[�ʤ~�os\��<��@t���yob��w�,n��7�n-�&����nS�#�L3�yƈr���ĳ��w�&��,��B�ۍr�|W69rl���M��G���ԸFK�6�;���eX�]����og�v�}m�N圲��ya��!��eyrW�ա7E�L�T���D䭠į,�"gpҪѠ�d�7����7��/T��/w���A���!��i��ڄK!�ؠ�ޑ��a�غ/bS.Z�n��y[o�^����.���m�댼~ig �3�w�V��ޙ���Hƒ�D$�1DR9�Pl��Y�O�4w�\97�oh]W�Ys�Pp.ZPW[��Fi�U�9i.t{��CE;�m�pSg8��]��-G	e��wѣ'���@���n22x�r�;�J�t�W����u͹������Z�(泂�gQ-	j�MH���:��Ӏ�9���:A�"��ѵaJ��N\j��sR�e���V�Y�0x��B�T�/�,n�A�um���x$ven���y#��O/W�B�d�4��i޾�ͷ�y8�Yx1pd�lkvuv�y�m�T�X�W�����q�KV���U�	|���x7u柷��&=�j�B��{s݂�盬1���3�)���o;�E�
��0��K���6�o�Ù�P"�]���aQ�r�������Fɗ\&{��o�o�>���"6�g�9�"գ�-�h��,%lYv��ζ�ӛYG���Ÿ'eH��DG��Γ��{hEu��	�M0���dX�Ɖ8�Zѩ�ũ������]+���3�F9�wxg�yRݬw��ؼ��)U��vZ��W&s�����=��D�n��ݼ��A,v�C{c�Ͷ]=ɈIDo%�q�5]��Zޢ�����u����k�E$p@�b�Y���0�b�ʕ=�{���W�hc�ݓ�Y���ddu��z�V��:�<,���6뀋=z_[�Ѻ�υ�Я ���Ao�p��{p����R&ژ���|n���4y�����b�$瞠=�uLQ2q�\L�����<z̊m�ٖ�ջb�(ڃ)�G�AY=P�s�|�gRU��s{,�xy�<��{i�
M����IL��+v��Y#8��ېH|�[4��l�[�6�n�d�*G9l�'���fy�컲�a��@찻{��ʼ(�8<y�r���c[�L��L��u{�1vؚ�}vn�ے΅{B�w��B��j���̓��`�m�+��Cfk`��+wR*�i��ؔ�$38��V�QM������F��[��˃���.�7}�8�^ln�׬W��K.;�b�B�*��ZN��ev˫�	�����>��%����J�\�Gf�w��ـ�;P�z_N4&b}�*N�Y�nGAڕ��m�i��P1��5a��n7�utZ��;L�뷎�0rܺW׊Vl,P��]ܖ+ڇC�m\<=l��}s�2[�<��&��9���A=�X��$,�5��Od��ɋg,�2ʱ�)�i��C��)uIZV�ygz� Z�՘���yb��L�C#5��fsj�՗��$;��V�������r�Ce8#kc���$�T�M
��=�K���:��*^��ha��ג���S�1z0{��B�)#��y�Z枝uz�눜�_b�
���w�M�l��笄��.i9&��%��M���߳��R��c��O-�O��B���Xn��W!��\Rdx�<�y��	T�_P�w6��p%¤��ZD���]�r��
.z��n���pj��uH�B�ئ?
7nrL|�G`I�ŭ�Wcq.�:��7�>�5s����bt��5����v�hb��N���[(��3E�&��3E�wĚ�U�$f�ve�:.����w��oz�۹y����@������E�C�LuÛ��*��ӗM+o�E�۔�=��[�F�������-������k��8�S�f���'{�.۶��#��a��axӈ�P���qq�,dY�r��P�zUs�~@+�J�o�;�4my,+rR�t�-\�Ի�-���!v�S1��MK7k��w79[s�ɍW�x��
�)$ǧ��d�'6w�g����q��Y&ZI�����R��I�`�y����j���걡,�ty�RP�m��R߬Q�%�Ƅ�o,�N$AY��lY����C���0�㊓Ȃ��̃9�;m6Ǒp����Bd����w�@죖����6�[J�aب��0K�"�h��§ۅ:ȃ�b�qc˰��A� �z���(��/_�jL�9���0�8�y�g|�'��:�I�2��(����<4�/��k3CI,~)��^���l�Ɠ����x�J*k��u�V��^�Gr��^v*bH3m�,"�B����|���(��p��1��3%y��i떯r�����@(eA�|�n�A��2��n1�zT+��*�j�o�N��:�b����HLy�ŉ,j�>���"f��6�1�/��\�_��~�8=�w�Ѭ<����n\���N��å�[�G�P^�]c;+�Jy���c8�ktv��,��;�I���_v+�㳸��qǪ�n��)�:3���pr�K٥-סCeO���2��ݘC�C�Qh\�=��11v��ڥ�y�r��'B�w��ߕ-ɱ���d�B�>=ػ��#lQ�5v����(+6�yJ���J��l�ξv�u�hҵ2��먏.}��۴�]���U5�=֕R�|M���+�+��M)���eK{Qi}R�n$�o�(@ת��.l�P�%��zA��w�ַ�3\�b75�o,�O�U�(�/1=ˇ�e����b��7�d�#��d׆@��{<�Qm��[���]H���r.����l�ϙ�ݘ��@�0g&��,Ow�����o�0�8ӌ�f�P9�WTպ�f�2-X�[Z��l:
t�+�GUZ��׀"F�ܬouև�rU]wJ�p�iv�+�Z�Iϖ��M� ݼ�u�|B)ڀlVC=���}a��f
��y=0�ݪj�Y��fW�jB_�h�=���5��H 7݅o��(�$=�/#C��2���{�e5Ё�n��vZCY�푆��c��FU6/��я;��*��Y��R��IVyZ�bc
æz�m~%�\�i����;@&�;_##�3����rf��;���0�#����V�h>q/U��8�f�M�y�eEH�9Iġ<�f7�fI�|�M v5����Q*�U�V��v���z�����ƕzaw����n5�o�Z]WeU�Z(���:l	-�Cr�1�������3��\�5�r���s+h���Ok���-c)WV����	�Զ��3��9�;E�wV�Bt�8�*1[��K�#(���;�Z�E!�l8��Ԯ6���{�k%��^������Nj��zWs��z�&������A�9�o��I�lf+�G�k�3���+���#�>�M]����X&{"nU��[2��]}k�������� ��<����
�r�����U���l�Rʂ�NR�*ۭ�)k������f\T�D6ԇ���x�� }��'|:/�h��{Q�՘*��O���c��AN/1mag�����1�5t��y�2;sT��07��;�*��Mo;e$i��v&t[�vm�pP�<��M����IW�=�=�Sژ%�)+�Q����%����T�v"�[-u"�Ⱥ�|���^ʽ�ak�Wt�5�/��l�0h3mk��~�3�" T�ya�r̽���K��S�QC��j�S/\+�S��yo ��g5��X�ݸ�ᎍ�箑ʰ�Spպd��gz�8 ����I��z`S�*���/ X��!1�TD]��r������´ke��b�k���K�6Jf�\\5r`��!طN�#2b��͊����WmK
�eZ;VgoKZ(��c������z��9�ƙ�]��{_�K��A+=��TG��l{�X��b��{ɠ&u�i�ty/p�^vD�K�I���I���vJ|bR�bM�hv^>]\���Y״��K��mޙm�d7�����Ç��xea:V�T�����N�zEB���I�X��|-:训D��u��7@�mhn�h��<:��f��F^�d�>bΥg�9�YU=�X�3��EG#���.�=�^Ǚ]�];��hP"�#pa�j�*��tv}yvnȳ�3�bj#�L��ݓ|����Qp��0nQ�{����6��_89<d�B��穒���Sv*g����L�K�����0r
מC��V������Qb��,;��xc�In�i/1d���:Qk���p]NZ�U����U�ZsP���NWl����Y��81��j�f�����j���D�_�����X�F��e��&��w�c�l���e��*q2dQ��UĶ�HT�eIP�U�{�b��u�u�`���J(SƇgq�A��Fܣ���;�M�
��:^\.�[���Y�:��D~�y���q�>��@�^�Gi����|5��չX��b��&�+�k&<���1��9F��v�v�A���~gi��r��z�4]K�5vhێ�^���v/]�S#9B��iai�u]s�/rsH�WK�*����^�`�H,�W��C�S�����w)t输�Wbn�y�a�Ƨ@#<������a�m*;K��T�=��eݲwY���gtc�(�04S�`�884ڮ7Őf5�����_n���A�����K݇
�
�6{u���Z+�^�������B΋�9Y����o���A�r�L��'a��/��+{b�:�,�]�z֫�.a�`NA���9}�Md��Թ�F���h9x["'���vu/<��7LΑ�[\6ݴ_ԑi0][�HYΫ%�z��Ѱ�@�{Z��!�_n�`#�mpi2���w-5m^��+F+R��@��/�zГ<���1λ'D���7�aj�`���ל
,G�i�����*�i�ZVdeж�F5x�-�ż�sťRM�nƊk^ɠ	#���ûG�Ry�o*P#�|�ˮD(B�R���+�i�z��u���]j�0��67{�z0��{�X#���]Br΋$]����b����%	}�%uu�g��F���`����vH�-z��V�E����?l���i�-2�;��%Z]	����U��V̭�w�;8Ƹqe��A�vr�OY&ef��p���{�ѧ=�x��p��Y�Id�9=Ё[���A����CZ����s.��C}q��ܭ�87�z�dԎNm���(�$����e�{K56Ӫ�����η]���������Ϊ�MAW�'��u�f�AI��?U�l��y!��w�aH���z�n[�Y�vB{�j��k1�l��Ţ5�	 ���GL��7�2�UX�M��t�,��l�T�H�Ҩ�<ymZ��U�A�����R�4%6�7���1<zX*��,6Q��GĿ��ٰ��'v�7�k�"��{�7ӖW��}u���h�'>��^��p�B�ް����-�<��A�w��j��N����6�wr�o��G2[H�X��3b��:V(Q�iM��R�.&��S��父Y�Jk�po�s��I�[ׄ��1��co-���6�kD�����i��
US��{��@EVc�p<��etZv�7;�I�afoiB�����HPS,@��v�K]b��P��<�P+m��S*-�.�����]N��寰�,4��/��t0�#�1 ���ek��uP��vB��wmbj1��B.������|99�<��w��|�w�8,>xE»0a�pB=Z��͵�Y��_ͤk`�]c��G@��u�f��a,O��r��C�{tU�"s	]W1i�2*(b����CW6qr���X�I��iB�7k7�=�I��;;wS6� �o��<���1Y$��J`�gq2�p�o7�H�XTR�6�׽�tz�ɛ�į��G�w��oZyju��
���.MFk��K���B'�K�~b�36��-p�8g:�79C#滹���wT��-i�Ь#1���u�e26ېX7F�ˤ{[��͔�`�C��1
Xaޏ��Yh�����Ç�� WS3�� d��:s �)vF��on4���aG���C�E9w��>݋4�-��3o������*;��u�ٜ4R����2�i�%滜��C���t�
>}u�n��i�=�S�OQ�Sn��Ɏ�)�ە���L�w��C9M�R�1B��Θ�$^-HmPX�_h�,��S�*�ˀV���jl�Ƴ��6�0i��	+~{��g4Q^B{�:L��n��=�����+h"U��I��%�Nh���yb�}�/�9��В�ι]iΫ¨'H�办O�4�˽����h�B;��8�,�2d�i�э$�b3qعt�t�Ѩ��!����K����n�Ŷz�dc��u��b�h��q��;�陗��֝Fj��[q�[��t�C�(�%-}�1�ͬ�
��{�&%������X�άfAֳ�0!�;&&`�=�0�P���|}��~E�nk�9��v�"��AYLu{F�U��E��N��n�V�ؼP2 q8Ujל�mp���^�/���D�R��M#[�Y�T?TN�.��ƂǭPj��uCm�=�\��Y�Sw3�}�`ڈ��m���NR��s����xh��Z��E=����.)o�9A���ޔ�ߎ� {��oQ�!-�5�b�jf�{r���W���'rj��}�7�������< �OW��x�=K��l9�7���h���]�%�7i3Z���9L8��:�]�	������X
N;X�J|�5V�:��ۓ;-��Rg���;��8��>�������v'��se��b���׺��ĕ���h�[W,�(�"�}!�֟��?-e���J���%=��T�ܾZ	[ux��B�3�k5�����vm9���Y{o�٥�H��0	�H��n>���3N�=�w�C��u&Mn��[��x��UOR"@���8�D���6�6��`�9����Pygr���g������D3w�0ֆ�b�m��O:����5b����H��c"�d\�/�u��6z��;~�q-�����2��S�t�O�bl�C�g�ɻ�� ���E�(|�umFnV�:��n�ݱ��3Yv�U�}�s��or)�ޘ�R��2r�N.(�Jj��'�	�˧i��ys��{��#��H��3>=�vpZ	�eje�U�X�"Ɍ�~�!�Br�3^���b�Κ��c��y�ɴ'�a0�7�u��z�R�[�4��ck'�[���x(��f��S���/�gi��Ѕy,Ֆl��K^
ۨ*�*Lt��e`����xP݈�ekID��,
�5��q��X&�v,��TU�ԗ���Ң��n%�!�g�>�<lØ�J�`�b���N��U�0]#�r� Ր>=��R�=�a�zk�`N.nS��8�:y}ׯ$d]5�Թ�r�@[�u���u�Gt��iO�{�#��tЅBw�oi�r�V���˖9v���-2�����(����.+	�1�-��iv��]20LL��������H� ��='pk�} ]�>F��犊w���j���wi��
��n�����0�H�ڑ���W���r}��,�,ܫ���boNKP�:;Y�tEģY| �E���`����u�]L�M�fM��2����[�j��`�n�r����Qh'�-)�����&�n���(D\�xr����!Hd{�G��MY������]�C�zC\W|{k#��6���(Z��m��7�v�\�rYi_d귈�PsL �ⷆP�5�8z�
+L�2b�yz�vqrS�O.Y���,�Ln�=� 1�N
���Du >u�f�ɹ�ε���Qb\֗�VYHӓ��hb����(�a���O���.�v �r�8̰�`.�t.� �F��?%�x 	P����Hv_�6Xde�P��W���]&�CP�]��J28�}�,��uu�y��YEr��U�,�֢�Qy���^�/q0�=T(��;=(�A�TC��;z�v��޵z0�處n�Uq�� Q�XU��Hv��.�_Z�dGݰP�Z}Қ�z�
�h����C���A���n��l�J�<�Z�$���3c�!�&`�����ǐ�s����l�Z�v��2�o�Aj��=��푢��ܡ/;]vv��J>���U S+Wr*fx���2���\'��X1�wm�2*�'�z]�H�Z�vu�#�!�cd<�R�4������,��fПtrR\���I���G����x����ɢtC'Z�����wۆ�б�T��VX%�B�;KQ�_v�v��l��.��.��#�o�:��M��2���;U�ˌ0�voX����u'uJTL	˦#g5��^�ۼMw����<�ʋ�{׫�ny*�0CO����P�z�8�t��A߽��0�D�P4�4F�ʓ\�h�Y�ֹ9�m�2�5��F���v&��RU�/+�a��_X�jM�*��%˹z��=B�w�&�z����t������`J3l����80��jγC��%+��c��#��S7C^QEԥ�I�J���q0��-�Ѽ�D71_��B����R��B��{24��1��ð�id˦�9�ry0�I�N�q�%>�'�Wt��(w�Z����7��l7��m��{�M�^%�t,c(geb6��9�Ciŋ�yc�i:���u��F_p0�$�7sb����%�zq�b���p	+uV�c�[�T8���O�fE������ �DU��e��>᳜;Ԩ�V
�sn���������ܫ�:�J4�r�����ŝkg.�V��^��Z%)s����w|\Z����qY�a�Ь�8���Y�ΜF^Ž�E���Ѹ[9D(CvX�9��q��&�!�E�zk ��ay��H.Y�D�隱fC"��[-��s`�X*�$H�kV����B1�0���CF�V�tq��}mGo��	�� ��R���q���,��w2K=�j����2�hǏ���a�'m�d&���s�`.�������3�K��ul�ڵJ,#b�^�R20�V�]�؛���w?@��n��0�Tf��Y6�8�B����G=�$<��>|� Gf���ة;NI=H<L�ѹ(�[�yb-`11��y6UȪE�gM���[�]�y_G~Y3�>��(,,w� <d�;��X���g"2�]9n�4]�	�e>����;�b�mn���'��t�vV���t�s�YO-r�I*���r켧7ֶ�j�@O�1f��/>@]Vf��Q۪��<��*���Sz�7��KS�#u��h�ך� m����k؞�ӫ��n�c j�Ω�u���	Lzlcs6\�s7��W_8���ڴ��y�qw��Ͳ,�Z�a٩�(0^���~��ZVy�U8|�6*ѱ�qTN��M��y˨�yc����ء���z�,	��C�)����H$�!�ǖi��y�h=\�[m+c����D!�3q�*{���\���mue����R�s�!`�%]���(,���<樆��+v��X�n�h�1��ԩ5R��3F�v��];���X()�:��/��'�36����{נ�Ax��];X�٨Hu�'�=V����Y�E;^��BC��[�08��zH�`�N����i ɻ֮to;wBũ�4���^������n��v����x���H|�K�L�ݚ�Q�}����0����yi[O��5���}�`h5pt}TU�4��f���O�Q�1v�zY��0姕��YE�
�� %yח�lѻT\A)f��U���5�g瘤sh@tf<o��^�2��o	vm�N����#ܒ'���P�~�sK�O>��)/zF�h��q�����݄e�B����d����f�����?_Kk2� O%��[���r����
m�g`c��
�&�ʶ�4_4�>��5��L��_�rx�{*�ј�\��s� ;n�Yn���l��\3f=��*�Rpn�Mr�H�t����j��� 
��27�"��)�j�x����X�4�W;:�{{7__�dq��.I�f��"ާ*��	H�Y�rsN�ƚ0/���y��F�gm.U'��:��l��c�(g:���~��z�����i��9�J���|)�0��(���p�j�\��7����к�6��e�׻ݟ��=��z��v9�Z��,0v7i���4��9���&ً�K�L�d��L㴷�k�Թ�NHZ�\�`�����̥�fi�앛q��Io�u�+4���&k+:�%�7g�;��~3G-D��ރ�	nR�u�@F�M1�Y���z��L3h�WO{�ȈL�����;"XQ���;��t"[ �wl̴��=�އ`$u
M��&��^Zi�{S=���YS��R�}֞+U�'������J����1p�\p�h�.�u������f�(y!��8B�j ��&��a,���J��Փ�wº�Ӭ�b�۩eh�XGC����
����^�:n(}�̷��׻��P�
I�C�J�l]�E��y ɜ2��g��^��|,n�f㭉dmo�(]Gh�ʠjG������n%]�m�ã��v�G������m�g����wp��^)ޅ>f�>|���r�6tT�N+��^/xOu^����Ko����cդI�~:}�	؆5���u,Ҋ�nrN�=U)�o�.7��0sQ��s�gaj��]؟�m�F{�}���s���D��#h(s��"@��&�u�!�:э��{1��ϙX*�N=��|.��u엀WQ΂\ ҳ8E�7��t���̵�q6�nN�m���F����y�稌�Յ��nWhm�-����Z�X.;'�}����=���X����*VZ�$U-m���X�����Z#V����1�QTDD+E��-�-�FU�X��UKe�*T�����j�XUm*Բڂ[E+V[kD-����j��Ԣ���UEV ��[T��,+,��D���(��Qj��
*�֣X�(�l��l�V�im�U[mJ������1kTEDQ��֭�J��Q�l�� �B�F�QU��j�Pm%V%lR�TRҪ0�lDP��� Ա���Ҫ��UF6��)R�T�P�UA�Eڂ �V�K-���-��kJ��Z6�X���U���m
�TQ��R��ڊ,TZ�m��Z[cJ��YY-��)hU�kliam��!mXT�Q���BѢ��R�QR�@��*�4���aiZ�D�(��[E�ZУ-�X��E�Q��clR�[��%�(�mRZX �mA��Ԫ,X�IF"��A�1X���R��J�Z�ґ��(����ﾽ�o*-��z���9��Xu��g4���t�q�8��}rd:�{M>w�~jŝ�ݒ�wx"S�6��G�y�s2��?������oH��쳷�:��Cun/���s.d�[�~~r��=�������E��~�����r��`�Xx�H{PC9fv7h���7C�U|�b���ѬM��+W����S�C�;:��I�^�Ȼ���ᬆ�6j�G^�T����a��*
b�B�J�G`Lޚ��Ǌ���ǳ�Ȇ��qN��.�Լ)U�۲Ýϼ�heL��A�>��?S�ܸ�.�Ai��������PZ�������eF��u=4�2�K��TmD��E�Q�4m��n��}ı>��b�"�;qB6�gp�w��e��Y*����1O�>m������������ӹ�P�4�E�u$�{(�l�j�vn��n���	t�f�8�SVk�$�˪�f��8�����1���+ir�����4�&�A�F�3K&�`��#�#�Э��u�W��6]WO�߼��h����v�]nh�����^V#�ɄA��zU�e�X��Z�������$nr�u)k�Ɍ�Ԋ�́���ԫB��[0ÅJ��k��y������B6�׷�8�|.s�a�݌��n��]}����F3ӻ��1�K������x�Qg��nk����X2x�:�����Ö���ĭ�&��Q����tNi^��a�޼:�c���4�\tx��WUY�y1F�g�Ɵ�v�X�o�/I��%�%��X������G9���P�g��~g��q=@ԃ+���lV��_����؞�+40��Yk�ssF�*�:�7��˃�>دrRϷ��j�G�,u�pJ��\L#�Ç���a�5�o�1ٿRW3����G��ו%�����Ք��Ӊ"��(�g**�1-͆��Zk�?9�mLjS�xt�O��A妁��:0m��-

�ןLaٷ��k���}EJ�tk�_$z}}6���~8��4�l
���
��Q7R."���={�{I7ت���S{!C�5���j���T�A��Ҭ��qFv U�F�WL�{��rV��y`J'g������dR�S��``��|9s��Vga91@�*)8���>uJ��3�pouJJ����f*��,��!X1��9�y�mh�n�1;:"��ؑr��gS�Imv���E�i��1g�-��/��t-���1����!iv�S���1��,ފ���K�xbK��{��<�H�����+���ܪq��Pޕ�>����3��o�\=�/!����Bm�!�&���W�[��o�)Aͧ��ԧB2���R�սփ�ʙjXۢ�=<��;�܆��s/.=�ܷ{7u(&�g[�r������}�}y鄵_O0Iap9� m�C��h���`Ks��oԺ��_�ό֯N�Z��wU��tAgH�,jf0T�8dU?	�@�x����]��r�+GO^#|�Q
��c��1aTC���C�0(߸��x�]���A���������;0qȨ]���n�*��Z��'uCE��C��n�=C�~Lװ0���>�¦7�mHiM��/d���UfɻʨQ�fa��b��(�y_���͝��E[�VVͣ�[�ƥSW����&׃͛jX��Wz�������2vSb�%���cg�T5�0v��]9�XǴ��R�g"�{6���zY����=�c��3Rq�U�p�^��]�h�l���0���&E_����6|�͵@?l���B�QZg#���&�x�y:���|�C���<��X)���$tmm_*Q6�ګ� %\lD��E���|͹*�3istz��j���6���m�.d��<3�/&c�k�c�+�& ��fa��pV���T3\�M�c�p��+yW��`8*����5�m�ۭ^�q��t��'q~�r�V���������Y�8a癯��i�e�W�Li}�D�yP��|��#��W�R��%�wm��ok��%��w�n�j�raz�`�9����y��;�����H:��{X<G�k>�\��[=����GF�ɝ��&r���i���6�*,c�Υn���>�	����:��鼯�]�����$r�>&̨��f���Z���`;�e�<;'���o�'F�Br�x�eA'�]j�硑����{��)�H���1���m��W�0_sD�xϘe�W���b�`V��T�pk��D�,)xrl���fm�\���9��;�:0i�6U8�i�W��XE�m?��@���Ws���G�5ƚ�K���*lG�>�U�X�_=H��,��x�2����̫帰h��q���2h�ʗ�^��
���7�3����6xgw��@�1�-zp�����V�HQF9L䘙�ܝf�4���lX�gՒ�%�;�����FI6��5	D�kM�5'2ESp"ͧA���;�,�i#֭��{j(r�?VI��{ں�.��g��BU^,��VD��j�}�P��$�\�r��������1�ȝB�4�c�!L��{2x�
��_K��o,R�L�us<Y����� TO�Y9�@�Տ�cv�:�l6�p"j3�7�T�XmD�Ꜯ�Y���quՄ�juwj�9gV�;+zr2ƚ���& Vl]�w�d{�D��8Զ��0t����]88�%�xi�f/؉@���b?�����x�Ox?�|=�0��W��Q_b����|��m�8m�tGIަ *T�W1�X}�z�ߞ��f���/�^�,����z����	���p�,���P��c�R��ȶ�8	xz1N���=~n�IP��!�"��]٪i
7�j�=�q�2���������jU�����jdu�E����%���;v�njн�s=����Z�k�z�66с� M]�Ga`V��BS}?G�{;�v����D����{<	{Z�oԟX/
/��ϸ?����r��`�Xx�Cغ�s��>�$2��y����]�ʭTj��ԅr�9�~j{|`�,�y���q�q!;(mI�)�4��vBVx���w#��(��f�м�<T|X�=���|�#i���qg�vYr��l�}nk�1�Ne8��Ϫ��7.,K'4�*c�h8�U0����1�{�s�h��u�h��ս����h�
2"e��O�� ��g1YMV�,c.}O�ͭD�z:�Yv,T����R�e��.��Ś!��]��U��M���sI~���_<�W����W�M��Q�C��]�'�]t���oީ����B��$8i|�N͞�fi��e2l�`j�ٜ��ot&�ȋ{r�{���i�����sfu&s���wY`����t�b;7~|Y�:	k�}����`�1��8�$}۬9y;��i��
����(�%{��I	7�SVm�>ȡv�E��ʃ{E����3�7��{�{1bJ�Q����<Aݤ6O��
j����	�O��^��e��>"ꛝ��m�l�ߠ�bg.�(ފ�ֹ�� h�8�l�I�a��$4!��-H���WdyM}�2�j��U��ڛ.68Cͧ�7|������ �a�Պ�����k�Z9�w]�Q֘�nf���\�R�"��E�xb�s�B�H2����ݞ���ѩ�7�%)�sWsfە)ENr���YغLޚ�*\�b�
�����x�V�� �թ�N�Q؀�����SU�����P}n�=r�;7,Utc՞��}�kY������*�zø���	ֻ�!�l�jht��t�� \��4��3���+�{k�8*@�������2���\�������8ڐ�t[�!�xB��Q3 �	�d#�[�8�f������^Vn��K[���)��Gry�2��"MT�^��=R��Tttm<W5�#��7_�:�d�h�g��1��LrM֡-�U�b�vU��7#�.��}�m�zRSŽ%b�k��>]TC���Б�䇵%�.)���ɧ+��]�6��G�7u�<����5�گwG&z��;���i�X%ӊ3���F�Zqo#�<��.�0�;��̩�] �:����Up����'؄�'T��t���7��^-mx^L>6~��6b�Ze�=�+�����F2I�n�1;: <��X�d�ט�U0wdqC�i҉{�������,�W��Z�u��E5!-9Z!����s��x;�[b�~�gD$�"*xB"*P�jܴ:�l�,y|��Z�\�E������V���x�Z���[ހzO{�8�y���i�jyX��cꮌ�-w���k{:z�t�`�|�zk�����_k'�g��;�0{��g�E�x��߉2u��˗`�>�/1�G�E�{��š����9��̯ee9=�Oׂ��K8�*ހ�����Q�P�Z��3ѤfaA�q� �0��+�y��C��gu�it_I9y������z��8FL�K��W�C������<9Q��գ�-2�������=�ե�#5-E������%8S7�K1�>��W�nA|;lB,���Lu�V�K`X��ͻ�^�9��{�׉`����VT�NJ	R��ܘ�����G���'m+��ϟ�s�h�.�tF�z�/�D+�E��V����͈]M�#�ڬ�ё�z��O�������K�3M�,��xe{�w��W}�OT�=��Kd��l���M$ߕZ����"��=j��l|r =Z�[}�h2��s,+�{B�ιB�����C�^d&���L�� teeo�*Q$[��S��ׂ���La�����a:�]�qY��-�{fԈ3�9|�����˗;k��Ҙ�;C�l\�\s���TV�s�LԛɈF���XhV�#M�E��u�,g;K�����{�������9��;��_U�`����	���q,j��=��)�s�.,�ݓ�T�#8l��GB����1G���*1A�}0���)�qt�5o��b�`ߗ�^��o�w�s-�}���o�ź�~v� ���L��;�|��8��$���>���.n�Z�̜wז����5u{�La��.®�f���C� 4��N�����=~���"Гփ��w�'��wy����lO+K� ��l%��<��j(	�̸�Q[ޣ�8�TrĆ���so�ژtΝ7(slZ^C^�@��������*�b~谏R���Km7Էǘ�wm3^��ǽ�pP�w]���AWYE]t!����1+�S.�$�ջݔ6�bTK܊MY!�M��#��c��8²[��jLz�63���q�z�}��t�g�,��Y��6�I����*�wR�z�\��_��I]l]y� ���lq
Ӥ�FŌv}Y!̒��q�Pci״��9�����<ká��uIw5��qVכ��o	�ØTl^�v{�ǲ*r;��1�g[̌wx�9�V��6�Q1p*桎t.����U�3^��cW�3ųѕ(F7<ٜ��ǰn���R�e*���@3�M�������I226gG!^�� ��W}-��{�3[�T��n��Y:��c��2�!I��ED)�#|�Ӛ��N.
f��;���͞"�R��V���S�	/��W륢f��6���j_k"��;����:��v�bbb	ɬ����R�W�ۭۗ��Di��|�Cr��6,}��]܊�-ɵ#��+6j:��θ�Q|�(;�|^�.^>ah=���c|@`Mz`�Q�FK��|�Jbl��dnb���Ʈ�2�|����"�&+�y�,CЉ�9I�h�㔇�qKK�.��j�db��}ȇ�+ob4RB�]w�7�.	wyϤuZ��U�n�E����F����UW�����A��?U�e����7��ԻJ�x���h�������a����e#+���[�1k��g_b�պL}H+�d/n��ޓ�������e}t��7�a_�a܋R�H��t�O���-���D�茛�ȸMkıj�U�3�����tk����r�q�&oM%��#J(��V�5qi9��kw�6ϟn����eYKثĈ��7�)�d�/�g�S�ܸ�K'[L�LX4{/.Y��0�a����p}S���G�]��6q����u�2b���O�x�	���d�1$�!���T��8_DVaءEF�l].j�]�x�mu	���H���s��uW�pm\M;��9��r��i�ɯ�d�����o�0��׮O��U����Pvi��E�;���E�}ђ��)��?Y'2�A3�^�b5���{Dƣ��+�,�Ut��q�a5ȫt+|Rɓ�]ӏ�F8F�Nc|; �umʵ�t���6-H��Z����8�j�Aۣ.;' �5��p��J!�Wy9�q���mM�b[qם�8���o�	�9}̓�6���
֊ߊ�2
La��ѱ|ϔ�Ӡ� z�)[��%���g��iEO�]��T��s!�{����[�L*��iĻ9�Ӛ�]��t���n�����@���R�z�|�*Q����:��5��}R�S��<7�4�������!��"�1�+�������۞\��y"X�Wz2�;�(�����z�lfr/����pm����0m���T�xP[�i�.�Ԁ�b�'v���qg� ���6{}�t�6rH�#NE�!@��H+G�9� ��*]|�%�}%�SԱѾ�]a���#�em�ҵ�M�^��S��WH��
�S��M�cCz:U�:���v�B��Dj�q��a ��Xi!���JAn�g2�g+5db����	��=3�-�a|���^�H�iQw����C7a{nU�!��� ��d�ew3F�s4S��n�-�깤n��b���r8`���V^�F�؆�j�	��[2V��k{f�M�AgZ|���8aH�fQŚ'<���B+��������e��%�@���5�d�"�4X���L�� g�Ry}"��o|�s�� �D�tO0vE�-Eϲ��k�!��豹�70\3>@�|ӹ�R�+�E�0�q
��2;k��r�v>��P��,=K���$݊:�����抉+�({�}�v@�/*6��S�hH�E�R`�Ӊһ�KY{�$����V�W�:
VN�'}3�o:��}L�j�"x��.+䑳�V�į����t�h�X�T8��An �(&�lm�}֕L.��q5���9�Ds��Z��kr�䭮��pq���;�R�U����C(�P�,���a�u;�9+Zt]=����l�ِ:
I�R'kjo\�)���;=u��.�g�	g�tf��=�ǧ7�s%��>�K����r����5gy������QW'%<bɒn���xï�0�{������Qޕ11#��Ke`u҇YCh]Çaf��0#V�	Y�hҮ��Y�d��Z4�P�]R��8���|ɽ�A��Ց�k���#9m�V��;Z�%U�qj�u���Ѱ&t�э��zk�<��H2"�����9HC|�l����߳��3V>�G�N��G�������*�_\>�M`yO�����;iP�f{ۋd���ہ2�}�tr{�W�k��*�^����6����s�'=��0�Z ��8]�B�5ZSxj��W�oT��*c]I�����NG�8��.�K���9g)\<���]�&N�jk�F��R���ˢPɚ�f���x�鲿Aʑj}�rݐӳ/�u��n���hΪp�ʠ� ˻[�V�oZj�ec�����z�jp��\�{���^��f����̨p�PH[�ӊ�V:ZG3�Q��u�
G#�(j�z�sA�8nn�]
=k�;���7�F�;���a���i�y����s�������(*ZXV�TШ�����%B��[h��"���mj�����U�b��jZ��ъ�U*���H�m�Tj��RŃl(
*(6�*��j�UQDm�kDX2[TE��X*���"E�ZX(
*EAEX�*
�#R����l�V"���AAR�V(���#R�b+%aQb ���[T*ڬ�iFҊ,V"5��UdUPX%���**EA(���""[,c-*�QV* �1B�ŭUKeDAV)b�#�(�%�QU���A��
(�*�QE���mAETE�������*�X�mUVҬe�E*[j��De����ŊҖ���X��bԨT�X(�UQ���Z�Ab[A�آ��UQ��
"��$TV*1EUb���AF,ETF(��)T`�b�`�Ԫ�*���2��TU*Q��EA�QU`��EX�Ub"*�(��"�(��
 �UDDV"
EDE������o�_�o]5	��:����~9�W�V�N�a�tn(Ki�~#,��N�ͬ�^�A�6���ugC�v�uln�:��ߏ��U+5�驆��J����R�"�Pdu�AMf�=��{j�kN�1[���^�k��r章WZw�P}n�=K��T��-5���/��5g4���7i�r���ѽ%�Ƭ<��`\x�!�ɍJ{æ��D�s�`�ϝ+�H��p��9U.�5�x�>c=�׹��]bS��#�U��8ڑjG@��("`��h���N��P,lNu��ζ�J1]�"��o�6�8����{P����=I�+�S�|�Y���}�/��/2�����ъ��-"�G:�.vUYys���p����.��U#�GE��_!߼�<>b�k۔�ÞR8h�p67d>�O���&��5�X�v���;�m�J>(�e�!�>�!.qf����Ͼ�O�Q==�Z���{㫑����2��L���	j����畆ܴ9w�^���xeז���7}#|M���ft"]E䪒��)��)����@EM1J�������R�zF��^W�VG|:;�ۅ?e<��WP���.җ���8��{���O�|�S��u+yV%�(��Y�(�o�qP΅yl��ZC���+���\xH�n�4�F��Um��6-������Xwwv+��6l}���:��l�<R���u���������^u(���b�;�)3�6��b+ d��N����py�x^�v}Aw����O2���D#T��pT�Y�A�qᙒΐy�b\�gO�Ĩ��ؚ�N�9���\��j_>����Wq�u��F���7Aq� ���+󂸻͚��ܻ�Ʊ�v�s�0&þ7�?
�E�;a����>ٶ�ǆJ��q����)k]Oi�/'.b)��ې����[>�A���X��f��4��V�z޲-�{�w�w�N��*��8��P�bp�	~z�ǈ��͵A�e�z��]�b�c��R��f�*�Wi�y�^�1��T��Mۅ��[/"GF���}n��^�D��,q��̫�=CB���|;&
��Y��+r9Õ}<�-�.mR9R�!�ƛ��u�
�j���p�=a�;�l���i�j|�B}[4�Sf@E9gy�:3��������o1��:�m[q�Q��(�b0��� B�ጞ�� ���ׇ�ezo+���k�)�`�{�aZ��e��
B"H�S�G�6�+n����)V��T����<�~�����M�����_6��*)�Π��)����љX���<��l�_�ӕ����1����Zi�[;���7E�{)q�u�j�Y��j����͹ܳ��:�#�,X6e�\Hgg@����F⅄Ϧ���F�>gD&�G�=�#����8m/��zv����N�a�K/����z���3��Y�~� 6����S���·�v`�=��:ؼ~���>r���ķA�:0i�6U8�(R��n�a.��tٴ��u��ʅ)���'�ʏ���a-���P�(��hs..%�=�Oo>���ڠʣ�v� �ʿ,,�/��cC���W�j"@s�X���1�H���{:�j�\�q��r��׾�d]H`"��
�f+;>�PB+$�b��f#*�s�Z�F��m$�X�|����FI/����	F���iy3���n��Oރ;�f<iN�ˈN))�J7���<�0l�v��W���BZf�״S���0��Z�~�=��{@P%/S�jߜ�'2*ߡ�n
�q9r�}�㝊���fhr�|(\Sfk�9��a��sU}m�
��G��Mz�R�?D}=�L@T�s�����g��^f��,�du�#T�;��P:��^m�x�ɩf�DX�yKL�UZ�E%p�ؔ��ԍt��W!��]�f�q&����=�+������ݟ[����KGjUd�2���V[yӭ�|�'k:�!z�˜��V3�g���[y�����0+$���:NU��߂˂�X��x����P��B�cY�'a��sM��9��n����(�3������qR�Ä!��{�Q�%��^#K�M�c ���ػx
��!��xe����uwF����!b{N��
O��Lʗ��z�h����0'L=b�yoL��7�_�v���'�Fk������o=�d5J�B=�O�6+�;D�F�Ҍqk{���g���^G��RwZ걝�	�]�Ɵrذ�Nù�(!9t��C�;:�y�6��c�#��y�k�"ߡ�Pp�CS��l~���ێ���y.x�J('���*(R�/�S�����V��L^�?�<�D�S�.�,��z�,�Ӭ���y7I'��e_m�M-b�:7���lg�V�+'���h��V�3[�_�fb=tKXo^���`�4J�|�vKޞ,ha�.�\vn��fV���}�nǠe�j�ښ�[2I��-u�^��a�~��"�Lo�$$�|`�՚��'�]WK7���8�3ɢ��8�ﰹ�(c�^���-o�+��2w�-��3�,Q�{w�9s^p�X��DoR;"������_n�.�[g���5u�ҝ�K1[fA�)�)�����+M�E��bm�OM�ka��[ޞ�E�^AVyu�Ň��ޛ�ģ��{��M_6:i8�����>H�1�����᪽��kI?*���O��Wq;K���x:��"���zRJ�����F�2�Ƅ��!uE�y0��i@=���-HH�_]iVW��y�[�!�^����*? ����ʈ}�w��茍��Cjh�;�@��m����8m�$�x�6 kN�Ց�Rc ^<�/���t�
�FA�ʩ��ػJ����@�����$_�*!k
����R�����߶+�G@AM��y�<̨���a�WV��<���t��֝�Tn�
�v.�T���zoʅ��
_q�ʿ
�����˧�-�"��"��Y���V_C��
2Ca��B�����N����%��eK�~�Rk�|3�u����\��7��=����+k�K�v$,l�v�@����ܧ)�K".|ТX�3UU�q��{�ۿgKKk�w5�7J����d _OR��:�-Q,R�~�2:C�G�͊tS�3d��9s�
�r������j2�]��ўحJE^��7��X�zMׅ�'1m�N���[1b*�gE��tt�5����Y���}��y��Zsۼ+EJ[�qq������}h�])��W}0������+Hx�d+���� ��}/=���*��9ϸ:���	�ԇV�������6bwfTP�]��?�l���f&[�U�>{�P���@�b��i��a�n�(/��<���v���~c
��&�C8��!�>�$9J*.���T3�ǍZŽ:�_:ɮ芹}#`W��!�&tE��؊T���P6���4G���͌���Gf���δK���f�چ��չ���@D)�.m���RG6E�0zH;U���h�����1�6E�6|AR2&���B��-wD&@�!��Ru�L�8v�]家��f9E���Մ[WjR�*OyC@���C��}�,�a�3^��-�ݡ9�R睟=��}�f���m๔�\ǡ��0Ki�.�0�e"(�G+󄣰b�zpTG>ַ4kBU^,��.:/dU�1X1k�hM��m���W�C�q�v�y:��0��NU�}\�3i�zf,\���]��z�����=���kޣ�
7���L=_ZxwS���1��n�.�S�ۼb�yy�fK߀\�@n���j����m�~�G}��!��0�\��'��Ҥ�3Gj�����S��#)[��E_-}L+V��r'#��\�J06��w�0��B��Fq�
:�Уuڹ;�^���}ץ���<�YBJ��4մz)ub������d�7���bT�gTX�M끣0�4t)�]c6&�v%U�����Sw}��4���Y׵=`m1��Uy�˅.�%1:6��r�}n�b�ұl�e�k;����H��N^�7�����-�lڐ|5Q�����ܨ.xL�Kۧr�P)��iֺ����>g��^�,�P�	���E��\hA[4�z��NY��e�@;/��n�y��<�t�K��Rҩcv��Aӊ�B(�hi�V2��Ƭ<ry�(s��Ѽ��fc�HA��N�����w�3%�S���xf�#p�w���^7�"N.�:���?@}��_]@*'e���Q�.���3��]
��}O/�a�0A��y4"�FbN�D�ͽ���63[���;�7<V��ޞ�+1p�.���=�\F�e���1-�a�@gM�N$H�h����d.��mlTB&���>�'(,/ʾ?L7�7�X�q!��������G~�,�3��x_f[�eۿQ8�x�Y~&&A�;o�X0&xO�C6xu��B�zܕ�t��n�.R{W[�"7�Z���L��Aw�0пT����%��5m����vjyU��|J���	�պ�Jd˼��n�jt3Nr�Ǯ����?�׏�8$���A��,��L;,`ZoS$�L=7��P�_^f��n�wU�Q[ )�{Nd ���j}����uَ=X��8^oW�����[��o�E>�ԍ?�wl8���s��	f�V4������S�f�����{��բ�:d�U�LVGG��L`s�ry*w|-	i��b���.��J��n\��6>|l�o�G8�y��/��lK�O��̦��q��y)��u�����ޕ��ݶ�n���"}Ԝ�ζ���p�O�9��|O����|���N��U+ �TT��a���!�a���z�OY�<�`�����h��v�T9�B�zȷi�pD�=�Ft\+�܊�����/��I^����=�VTP������q�Lt�׊�d���[W�����/;�d&�
�A{f�_Ǽ֯@����06�
���*�G�E�j'�Y&�����m�t�Sp��V���J��<�z*
��lWj��3@�Q�6/�b�役��L�R�Q�nG�f���X��~���_,>�+����~j}�!񝅝A)<O�����Vj�b�s��:ƙ��g�WHa�@1���W���J�ş~�:>/佞3�Y~{d63��S�q���3]I�)�K%�����o�w�t��{�/&z�jF��u���`��zat]9�P_uN�v���}>g"h���Pɛ�l�����{����(�B��mո�QJ�9�_`�#9\�.ɽQ���u0/�����Z�UO��BKhZ���Kq|���}h��K��^�S�֟yx�7@��:r�����۾���|��э?jH����>��'�r"��.<@ѴdD�z�*��5N�գyE�-����8 �B�"��n(A>3�غ]b;7/�Řmu	��}��tc]P�l[���L@!��#����<hs�6�"�L�$��<pҽ�?m���x߇��az�'��+�idMl��X
�����=1
��`߹OU�#S�D�����/,"r���N�}�>s�"a�{��r�ͣAۦ�,&v]A�f�L�hD�����;����Q8ަ5T�2ʥ�LeNz9�A�L@9.��Q��C�茇i�� ܩt
�@�>�ҏ��]�<�e�P�i�Ӵ�����X^<��\��
!CR5�z6�h�u\���Lkk�Ca���Ev��f.v-8��`�}�!�x��z�{��2T�J�f)? T�������*E�8����K�J��A+�1=��g�W�w����:~����ܿ{�u�C����3�}d�Y���s�x���i
��^Y4�����'��1'=����E�a�
��;�����J@Ŋ���2~�R˛lI^�c0�d�>௨գ{�K�SH����]�:�ᒮ
���g�892��b���ni�JKI�G=�;�h�Z�K&pN�Z9*7�`T1�1�9�뗷�..$a5����e���1�����'{clL\���V�j�<��f� �>�(��M0�~�I6��q<2��+��Sa�08�<�q=5��$��O%�J�2~q��f�A���������i����E4�*J��A�yG����Ԇ|V���~ܼp��Y����x�l���&�~aRoϰX�~�u'���S��8�~�@�O���y��ṳ+�g�ɷ�OS��=�L�%2k(���O�(�G?d�G�s�|>���2��7��)s������VT*C��{��eg�1���X5+5��N!�1����b,�
��z��J�;�̓h
(|�������>g�5�:��kV�:ǅǲ=�� �~w�A����φ�w�.��4ͲT���UT��@���F ���y5�o�,����XsT�Ͱ��C�*)���l:�C�ug�Y3���fӏ��m!���b���}� A)�X��!s{��>����ss�~�� d�c 3�TP��a�0�s�wk���iPQ0*q?��J��ɯ���)
����>C�H)���?:IԨ���O̟�`�L������Q��}����P��������@�5�a��-�r�i�~T�'O{��d�ʘ��aRu
Ɍ����a�ϻ�AՋ'�γ�((
)�&o��q��7=�:ﴅC����Ȭ����^8�
=����s�L{���yM�� ��
&����f�,</2݇�B�xw�wv河Hg���"��J�9�§�:�$٭`kv��Y�=5t����+��_��=ҍ����;�G���2 $��4��$��1�2o;�>��aY�NwXu��T�{>�M����d�u�8����
���&3s��� ���]Ȧ��
�����w�ϵ������z�2��E>a�b'�1��d�Y�<ì6�դ�y�Y��1}kaS��c��a�a��S�°�u��~��-`Vi&�w6�������X�#_	��i��gK}�������e!X|��YuI�e!��?$��OR���ɉ�'�0�ޡR�O7��w��ݾ[&�����^�b,�eN���}����Y8��:����L*�Nj��s��7���~���z5�;ld�X�j.��e �u���=.V;�#��qI����6�m\Z���2�`�	�ݩ{7�"���i'45�T�U�ڙCL�ú��`��6�A�+b��+�j�	�F�u�cr�f��gt\��H���m�W�\0�*��ZΡ��r9pE���麒�a˒u_D)E�R7j�H�g1Ϸl�0[N,�)q��6������)Y3Gm��K&�(�a t��r��������ӛT�ge�-�y5N)�-Y��]��o@��5n����v�7� :y:��ԡZ:����arӵ�@�.��r:���������|��)�Bk��K��ʱn��A��},l؊b'Fغ��0"���L�q�un��l���:�����h�v��4NԷǮp����.N�r��oͰ*�(/H��N���Z�ue�K�T��V�V�<IΏr��Y��QJ�yJ���e,���\�u@�z��tmO�D��>S�p�h৸z{
^����c��lL������1mx,�7-�6XVu��fw5�ڎ(���x��(nwEr��n�>Ě��*��3}�C#h�L�7��<�4���°7���v�,��}��(�O&o�b:��|�1�D/�K�9�a%u�#�8Ȩ�!�N��:Bc��#��N�$�f=s���N8�����L�=�rҥʜ�v-��y��HKn�%��՞(b4*^�Md0b��'�./IS�1q���W���B`��R���e�.q�(���1pK=�.�(���*xs����7'	���Ǣ.�����d��S�8ʴ/�.�c݃�\<O/x��5�q�g���*�*�V�m�z�-��m
��n�/�xҋ^������X�qK���/z�;����+{v�ɸ��*I�N�T��1I��v��"!57y7b�j������e�q�,H�ƍ �+��Q��D+�ᝥX��o���9se�<��\ĩ����R���gHU�.�uҼz�pb���	�[Գ�CQ�u����i�(�ئ'���[JŢʦ�jP��Xo^PNP� ���p��ϾQsk3U�Jf1su���_o4���V�_6�y�l}��6�c�h}AvШ�jgt��D��uB�*�m�LD1{q���ٱz�I��A��}�q�Btv��+��aׁ�q��Ljmn"��r^v} Mpuv屝����kp�<R�?S�z�|M]��CiMY{na�2n�mNap�ǫ0��{��>"^�D*u p*ʝ��k�}W9����f�w>�Ț�/RUEV+Zhm`��_7j�n�G�9f+�vb�\ȗ-��8�NǞ~�A��7	�ylÔ�B��W$Qcz��Ho�]d{C6�ok���tz�A��gkJ\�,�Lz�ޙ]��~��/Kok�Sǘ+ΘO4�z��,�����=("�X��V*2(�d�������Ԕ`�
�j
�
��"DF,QAE�0E�QU�����+U���TUU����`��d���E`��QQb�(���Ab �U��������X�A������V"���DEU%���"��
��*���ATX��"�+QF*��ł�"(+�UUTU`�����[b�Z���QET1PUQPUc"�(�"�*+R�Kh�DDAb���
��*"�cF�QDZ�*�ԕ� �E�"E�%�PE�$TAUE,U`"(�Q��� �QUQA�Ŋ�Q��A������U1EPTUTQb�Ub1�(*���T�2+��*����APb�H�1�:�4�\	�3x�>�d�<�3��.���5�ľ-	)-��8%\%kx+:�kyZ�˛ݚ+� ��N]��8�^�5_��1vl>s�g~���3��&�SC�0��*O�o�oEd��R75ܟ0��'��X~݆3�J�d�{��)=@�<фⲤl߶N�Ê�I��7l5��G_���eQ;\�{?~��+�ks�� $�Q�P�0�x��bԗv��Y�����C�CL6w����������Lt��\��6ϙ=����0�³l�<�|��d���iU �������<�痞sg/����;�Y�?%�HW�>L��y���}����TRs��a�����}������y��0�C�C��ࡦy�ɉ<�p�,6§��xn�'�VayOu�9�у�K�oV�����r�4��q�c�P��~ݬ
ϐ��f�PQz�����Rm���d>f��+3=�9����(��4�$�4�'��'̚q�/p���M�T������Xj������d��MV��������Qd�*~N�3	��B�l�5l�&0�?]$��>���S��s�|N�T�}�rm8����,>a_Y4�����d�g+�{������_f���1��7" xD��X"O�� ���y�,=T+<Y>Ձ�YY�;����4��a��:�>��3�0�S���ա��r�=Ld�����J����_w���ӿ!�����Q�k=�w3!X|³����0��2y��EIUR
q��T��8�^R�7�4��i�i����Qf�*i��z�rwi�%Ns�Ù�n`]G���#g3�����!�6�ud�<;�"�l*gl</2m'P�4��u���Xq�MO9����`Vq<�rAAE��s(�*M!�~֤���B����wI��=F+��~���
;�<�q�늁�?oH)�N���1� ����񇻰ĞOy���<J�+9���&2��8)4��T6s2V[g�La�޼ɴ��m!s2q��(�=޸A�J�9ym}sH��}�(� 1��'�;@���a�
���w^�h�3�J�6k�|��S�<;��=VT�9��H{�T+���9����p�mE&�{��J��1=C��ٛ�hZg~��a�k(]�po�����V=ٝ�l�}B
r:�bd�w3���}rm�<e�)ClT�Hx���˦\۶\���w��"�E�<�Ic������/�O�Y��wVf�?�\������kaF�ں�:g���]��iq�����b�NjM�� �a���2|¤7ho>�i�:Ɍ�B�=I]=@�=��Y�M�p����0��o5��u�u��bi%UH>��GP6���N3ɾd��Y ��k����^����|;�G��e�{�1�a�1P����J��b���P�AՓ̱f��1���r��Vo�LO!iXc
��>��J�a�����
ÌP�M��&=F2��߫�b���u�{� ���7�Ci�I�y��~e�!_5����'�s,��c?$��O{LE �2{�ٶ�*A���I��!�~�r����yb����(�v7.M�ןK����@���S���Y�g�La��T�A�OO��uf2T4}�h�O�'P+3,����'�v���i���ɿ}ÞR?2W���n�AM;��4$ⲤϹ��髋�g��s6~E���>���?~�u�C-��W�1�CH
({��>v���bm�O��ă톐ٮ�E��Hj�A�p�4�M2c�4��WǬ=��i?!Y�'��!Xz³��j������|xf!�ɓ��������ǾHi6���k�bm�Y�!�2�R�<�3L�x�ݤ���Y��!�+���H)�3}�=Ci�k"śLa����OwI�
�wd��o�{����_�����f��@Qa�<������;w���P+���4�Rw-`]��O�4�����sy&��
�g�h9��/��s����I�7���@���CG��M"�S�Xo��'�y����ꨭ~����0ǀ�/�}�m1�����tu@�V~|�0�@Qd��ɤ�)*O���d�e�u�����u�o��svq��xg5�N�z�~@���i>dӟY�כdԔ��U��{�nV���i�#	7���~�M8ɼ��^���bOU�%�~�<�;�04��l9q��CS�퓎���1:�רm �a����,�
�֟y�gu�}]�'3���Z�l��cި�ާ^��+��xw�q
�a����B��
�u�����9�<ԛOUT��� T����H?RѾ`,�m!���%f�|��̰�g7{�ߑ�S<f'�y�,'SGv�#E����+..�8݉�BKvAǲ<�W5j�kqg��S9=�s|�A��9Q�t4OEpiW�!4��xd�TŨ�����:ѫ�<,�y��d5#�<�r���F�(mX}4�ë$;�{����l�bGF����� z*�G'�5{��
q���hq1H<�9a�,�q�0�w!��?!Y�P���i�a�wz3�I�+<;���a�5�AC�嬛5M3��"�o쁤P ���z���Fcc��*�b�?8ۯ��=�l���4��e'YǺ�q'y�d:�H)�{���\B�~��Mv��cv���m!��i*l��U&�N��O�IRu��'Ϧg���,���7�!w���?=���PY�~�~g�̞݇���=d���t�Ԟ�G�=J�|͞�q�l���䒫O��q!�s�U$��=�»�^)��bc��ǌP<>��@�Ԭ��'��P�A���̆�gXT��z��J�:ɞ��1�+�����O�Vu��0<�B���Ý�l�����s�T�%T0�{ǿn]��}�?�w߇�E�"��G�����ٷY�bC�������>�I�4���&���COq�+i8�g�uI�+<�=��i�C�|�#�� d}���h����w�a�������a��E����8�h~I�����βT=9�4��+���x��,��{C�M0�?e'�P��I���m'P�7��~t�x� V!�Hg���,x_�
�r<e�����~�7�ݚHe�m;����IR7`u��������2z�l���<a�&�m٬���d�޵�i=d��������S�O{u�B��
�*�������ci
nz���k���ߝ&�2i1��*T
$�O���;����T4���P�Vx�2p����Y�>���1H:�����gXV.d5�=I_�=܋���������U]�~ᷫ_O]���wHI���ɽ~������m���@�>��Y*m����@����c:� ����2m�>L`w�� �L4����
���5߰Y�?��g#L��z�7߯���7����X�i��=���Y���ړi��a��P1'���M0��(��0�Iܵ9�&��%AO�>���M2o���x��d�.��y�m��3s����F:����rm���x��+N1����!�5���U�t>�y��𡯞�;l{Gk���p��� 	�V���3�ז�`�~��rל�G&c���H��.E�*�Րaü��?��}S�֨[�V�C�_�Y�,s�wOiv�W�-+������&.�?_UW��5s_�{���?��
�Af��L��?%E!��֏̟�`�B��T�����m~o3���)��2N��IY�l���8�l�<9��=aRu<wn��������_�S�S{~y���;K����A#��BȄ]��$��LC��Eߴ�a��m��&�H)���_�7�P�T���Q'��4�R3�C��H{i��'2��c��`q�Y�s�|�߿{�.���tk����=Cs�w��~aY�9�y�$���{߰<@QB��y�����?!^v��z�T?k��g����'����%M���3���&��}�����]��Q����?�H� �:Y���a���h:�E ����f��8�0�9���JŚO�����C�I�+���yd��6sX,4�{@Ĝ�w��Y�-@��e��� Y~kc���Y�++�n���o_g`|ϙ*���Q0*q��ĚC�d����ԅa��l��C�R8��w��?%E���%O�?8�x����~�bc7��H}l<��E4�*J���w/�s��>{ߵ�p��Ͼ�����?2zʞ���5a�4��-�s�d�a�&�9���l�O?] (�Y>q���$�
�'���ṳ+��٧�O��>;��:�_̚�)��`
|�F�7�"ӷ]�s[����N��V~H<�t���8�T�����eg�1�¢��R�ɿ�N��1��3�0�Y��v�Cԕ�w�d�@QC����}q|�eY�M氅{��|��}��|:�T�c
a]�q�4º���2T��쪩8��{����$S�w ��?&0�V� �l6^a�>B���i�f!�:�3l��%b�'��������}�wt�w���O=p���3߬��������{�!��Cm��6s���
��ns�wk���6_p�(��8�5I���G�rk��a�!{��9���O�I��N�E���a����wL���]n��x��G��������7����ć��y܇��|�*O{��d�ʘ���:�d�[}9�+&�q�Cs��PuH{l�*
�m����N T�B�8��3�U�ߦqv��`kJ���{1��^�o���H$e�e֧n��z��_l�'^&޽:o�Z e�v��/KG/�z�6���=�e��`�#h#GU�t��dJ-֫�.�_h�C5̙����qܗV�),%�gL�ř9k��� <W[Q�U����!P����6�Փ���ed�Y7��>� ��
&��U�H<�ya�Xz�T�Ձ�YY�3���,
Ԯ�s�O�uI�k[���@��>���i��W��rj��`xL�ĕ�a��Pѿ�M;z��6�l�:��s x}t°��'{�<��c+%M3_s&�R
q��2i:��Hw�p�|Af��l�� �idh���^��Ef��m������@0�Q@��c�m=C0/�Jś�>a���#���Ɉ�n0�
���<Ci����&�V�\���Z���M��m� �9��'�C���[6�~�����M�����Y��+�Ͼ�wI��C�kZ�$�ğ���f����z��38�H>�7<�a��bCv�d�VqRVj{a��u�:�o�6��&=�74(���g�j�8���l�#ި��W�{���[4��a6�����i]& T������Y>�d�M�>a��OS����g̕�ɿ}ޅ ��<фⲤl�����qP�=���Oˣ�c�(�qɹ����>"c��S���x�����Ͼͳ�<OP��!��	|���f�;CI�a���ڞ�b�l��)4��!��a�g̞��OM٦�Vm�s��͐_8���7��k�V��OV�Xh��<�!H)�;��I�>q~�?R�:���y���O��P�x��*)=}�����4�'�7��~�V.�<�Om!��{�����&$�k�i�(��~�}՛f�+7yY���ã���q'�+^S��L:¡�9���`Vq��^0?���I�>�}����
��3�C�I������L�N8�IQ�{��|ɧ��&0<!H�\����'��X2%�Z<��5u��ҧkv���۠x���%}Փd�>O-&$�
ɾY�βc�}��'m!��猘���g;C�ӈ'�uܛN2~s��K���Ќ����!��/�wr;�E��ﱜd�!��r]�H)�&����eH=�9������MY>Ձ�YY���mE��\J�0��C��ya��n~�a������d���� �DW�����N٫6Yw��瞵YM��xT�A��Sxӡ7�Zy�85�s�P�@�m����G�X�I�yٯ}���ŔEK;���P��e]o��������Z3���;mZ�u�9g�I2��O�%�r�b�+���5�������{�{�:���P�^���z��|@���u��Cl�ɬ�d=��
�����~�~�,�'u�*J��S���*|��\a�Xg)
��͞}��ZAvSl>M��
�<ݓl8�C�s����9r����������Ci�%N�y�gɌ1!��O~�q��Y1;�"�l*gl</2m'P�4��u���Xq�Ms'�����gl4����'�(�*C J'�����N��\M����b��}��Ǿ�����I�9���3�O�IԺ�H)���ܡ�P����'�=݆$�{�n��ViXy9���&2����I��B������?2c&yf�~A���ݼ�sG�־=�ߵ�������*�v�$��q���P����r�����W�O����|�^��]�{���!�{��'�ʁ��0�ir�J�|�27`cY]�w
��R\�n���G���=��3��+�Vi�&���7v�m��14y�8¤7hl3�&��1��TP�%t�~�	P��&�y>�i��+6��d;�a�a��M����ރ� Q@'�Y�W������y!w.sﾮg߹'=�+�/u�
m!�@�}�4�|���*/��1+Y�h7�!���'�b�'c�{\�����H��T�l���T+E�?����x�ex�1��^�ؼ�5u���O��gg��&�PQq�a��I��ud����~5����'�s,�7d�~I�ě=�E �2o��� ���i��!���@B?x���;�z�0%��v��Ҕ��Ā	��<0f��~D�/?�c�NˋZwe��f���lX�g��z۾̓���M ��$C�9,XH�8>_{a�%o�[���Y��X~cy�4K?Bc�Տ��ﻙoz���w�g���2L0��>*vb��MA�:R@|0����fJ"�)��:c�¤.��V�&1�nk���صa��mAo�N�.o�R�ݓ\��1�6���LC<B����g�/j�pb�GV�����D�3i'�WWʵ+\�$����+��-=��r��Xv�Κ�;��,l'hj�On�Ѿ����2��e}�{�d����r��g�}Q@�ѕ,���D��N���Շp�z�B�̾��f�����p�N]T��03g��qP���O�<����ni�_=lq� ��M�%�=����L\�T��*(���|���C�#�ep���j�ώ*�.��oa��p��a�T�s�W8ެ���������ǎ�6���%���is�M<ݔ�5}.L�*{����'��K��Dg[�a2-��vgh�>,{���@�Hm#m�UP�6��tK{K��'��'&��8�D%7���q����;�aWEG.�^�6�����8s1,��2(\��+��~6�ze!�]Ha�/P��7������B
�� `�?4&��)�[����_�7��ig�䴚Js�8�V}�RX���ێ�&oM�M�*"&8�W^�|�,�x���b����b�>5�6��A�H��ʷ>4��w�z�Z����ɱ+!�f��}D��	3�1~4z�US
j���j6o�
�z\{i��v��=�SJ��hJV�~ش����b��_��6��ڻ�r��h��-�L�t)v�q���g�-ᆟ�w#�hd\��^���<#��y���]��k�iK�w�K�y�8s:F9L�/y��;XB:m�$5ӻ��	3���k*�n,�C gu�G��=�K3v�nq=��n�/�I�~���7��.o�ł��t��r�<Y��SH��ٙ�8v�����<5�!���Z3|'��mP<E���RHOpc�
j�z�<$��QiL��������釽�"��eA�6�uc�9<zbvS�lE���ET�.�-��׹0�OS�`�D{⌱}�22*�]Ss�6�!m�s���8��ܘ=������v���*��q*�P�|�!�7��5�W>�*>�p��J!�Wy�l�\�s���1�9�Uz�:6ޡ�4Bñ$6GXjl#�b���ȼx0_3��^EZ��[0��{�z�4����7�9�l��k��j�\�XN,�X����϶Yqu'>v�r7��'y4���!��OPڭ m�[�7�-�M,���B�%S��8�3��N��}Бq�5{[�)}�e����g���9{��ߏ��\�ԧ��4��uR�)��}�j���X��5��D�٦W�����>��./�g���*g=7CI��(aN��X�����֟zzɳ���uxmƟ%GK�+4��1I���}r��O�&:5�=�F���U*|{�����Υe�� �БvW
�;�Vydw�ӲE�j�(�Nܙ�&B���=�8^+�!3%�N�pϝ�ݎ�ǺIJ;>�����$��J&X�G����z���qSB�sg���AGx��mW����wzp�Z�$�'�_MC�c7J����F��#d+�ъ��$<�)�W�,"r�*��Yv�[n��1��ָ�3~����\�a>3�g�=1<�Ƈ����ꊥ�eU�n����x�y;��fy9�{�0�1���̾:7�;>��)����L�[�Or�Vնms=~�Kg:�O��P��:�=���za-W���k�]�6N.8�P���͓e���Z|��~�ډ^��%w���B�.Z��1�ǐin�ĜL֩#]`�DH;U��VC���>3�����e�xP�����Kl���5E�7}��K�1^�4�)��Z2}�3|�[��Ϛ�U
�ܘ��B+�!�=�)�u|�/�J�N7H/&
����'�1�{a�����=�NO���)�X7@���i�ʝS�� T\Bc������6tC���J.}�Ck�=�Ơ}�mK�/޻�9�R�udמ���;��b�N�>��I��D5�_�ѧM>ś5v���O qj��κ��p9�w\$X���w�W5�KuP͇kv�{�J�ԔY;d��0�K����-�S�#�/Q�^�%7o�/$��X�5��|���W۝�s��F)��W�{��v[�-7Q9:����Vp�r!�n�V`.������k#<ث�xf�*�ٽ�7}���f���է�V�'�k�M�/~pL*�{�����7�VXo{ʍ�+��+�Řa��ʹ��6
�a������=ci�>�^e7n�Y.���3i��UY�*�~��m�{�*��z�E���"�{
�R��#��崭 �S��*��})�o��N�W��~5����|�ҟa������E��E�|zx�{9��Z.�X�K0l�Fg�L��
�ɝ��ʛ�1.��\8<���!=_?@.!Ŋ{��M:���w�<i����+��΅+G����ݓ�T�+}w�lbF��3�`S��1��x�K��y�I���j�x�힃�q˿utu�1��S��_�#Z�sB7�#1z��n���r�U,oD��Vq_�@mQ��o�U����.�_k�'�?y�P�+V��9���_^y5�o�ӥ��x�y֬"�6�:Ȣ.�RpK���za��"��l�c�~�W"�a�cl�bFn* U���V�i����E�[�#wfĦp[��7|�f���yE��� ��/"����B�2{_��c�nR�1���c۹p�m1�����ʝr�WV��/U��������Н��\ �p^��)`��Z�-���<J���;��y�_^&�J��PwJ{˫��2�r1:o�M�y�n^b�s���aAu�ij��?�@���Re�_A�\Z�6��r��f7*�N%�v��i�1�֢�@�.���I�ta�XJPZ��M����I�+T�x��ۄt'�@���쁇R�Gd<�������2�ѩ� �^���F�/(�vP�H���/�����3����wd�W8����[�Rk����V�M�X=�
�o!퓠�cm7��+r޹�Z�WDh�E�S��z T&ҏ ���E-���9�dܷ�[�;�2�\ϑ��Ll�f�E�1K��o�XmtD	&���VA�Y�w��8}X�;qјE���%rat��e�֨4MǄ.�� rqVmܚ5�nQ����1eɡR�6Qگ�\FC:�n����h^3��o-�:���ŹާWbE��2�ي��Q4}R�3���/M>�X�U�S�i����,����ӕ?/y����Y�ʌ���7
}��܇FӶ���EN}�1��@fڽ��G�
Pn��l4��N���e<ԇOBo/y�j>����b�_��R�5���rX$["�������;�R�3wqwW*x��=GEJ�w��tc�f��lo`;;L �X.���ӭ%�z�:T|��r%N�j5vҶP��R�d�]��x�o�\q��d@6���x��im�b91�L0�K9���F�K>�z�t�pTB���%��c� �c<Q��3|{U�@�r���L�ۖd��_0��{�\�j���{m�Wui��q��k;t��ʇ2�Ԑ�w
�%(�������u���u���j_���Z2���d�r��C��>������4/R����ȇ���k.���8���#���v�9���o��\I5y��ӎ�b�����LDl��{���1AXP�U]&9�!U�B8gPjT�-����R{rS�s��t�n��q�X�s�]�8�8��voqGnĳ�vd�a<����j�����{�>�N[/{Є�B�ws�	������5ȷ�xvlWY�Iޚ�]�s<��WX5+Δ��h�a%���N�3���5����PϹ�ObAyQ�8�&Ujm��F�Yr��չ�Ѱ�ﮅ�-�8Z���k����oy�O+f�V|߸y,X�Okf��E�:f��"|�����=^=�J\���(ؐ�&y���(3�px\Ȫa�r4�B��^�p��,�ۏL)+Dݍ�^J�p\���/�m��^l|��җ��Oc�[�m��<[��g�J��}&��u�`ODGl^k�ׁ,���*׿{�����QFF5����1V�* ԩl�UDDE-�ʱE)l��
Db���H�m)�H�DF�V�
**���1+%��m*UV`��*"""���b�1aYPF*5+#li`�"(�Q��,UX�AX"��b����V�cDb��mEX�"�*E���#PX�0UX��رUb�E`�TA��� �"
�TeUTH�ETdQ�b�l�k%��EV �1UX��1X1dE"1F$� ��bȨ��!mb�b�(**�EDPX("
��"�,DDkV,QV��Db��J�`�U�TF*(�*���h�����b"���+E��U��*�"��
�PF$TX��((��TU�UKJ�ұ� ���LJ�+"(�9C�
�"1E�m����b��������/����J�9Ï"ց��;܇�ޒ���7N�������D/��_i�t
ڣ[88%&o�7WFev~����<���������� ��2��#O� �ʾYb�_��cC���L����5�.��a�m��p��@�ň�>�zU�Mx�C�5�ƃy3�F��%�N�t}{��|V�X[���ԁr����"�J�/��8.��>1�M�n �A,����Q��5��]ד��vݽ�(�/Q����F���z�L ��ʶ�*vc U�Fs�u%��7����.�O��?�+�Z�~g�����|��� ��fSIA�O���M'p.ܸܞbn�V>�HQ܎�`]��>��0����0�d׫��ה��K7��Gn�r�	�~3��.���9Ypէ÷�5�3Ӌ���3�������F��+��|��_3��=i��2�)�[�f���pX�l(2��b�R6+x7j$���QqC�����x��X"\��Ջ�4�::_E�F鍊����+S#�2-�>���W��)ql��
Ďɋ�ӳ8�K�MC�q�묂?v>˫�z�d%7�q���噧ЏEB��k�G�;���;ւ��:Gg]�jZ7Ɨ|������jn�_����2Γ�ǿk͐��T��rm��ɲ8����j���?/\o�wQ �S�,@��S6�i����ҝb�F�֕i���+�O��g -��#c���Qu;�n:�\!����{�NfF�u3W��;�l�N���K�!�\F��Vm{�Ņs��A��P$A�;;����|W(ת�~3��Ρ>�zM��Q�:��_�h�y����ƶ�����[���Wƃ*x�J(��B؆�44��H��*��!�^3��f���C�.֝�J�"]c�N'�,4�T���q�US
:rQ�B�F�x�C���{�Mz˪��l����/f*[��vU!�	��&�+9ۊ06`���+dbrd�f�N�\�M)�l���z���$����z|6c&�@ȉ�s���qo�2����Y��ҧ�Kp�O�y�v����^0�纬��Q<�ߨJ�zxj���-�xU.�,���F�z���v��0�����nwf��-�4��!uq��\n��U�u�4�1��I���rd��cg�A�9,�!��)����k�kЄf҈p��Mf�+�N�f7Q-E��;X��g��cO��x:9��6 kN�VGJLa��h�wND݊�^߯��
#�tS����9K��{�!�īXA�f�����B��1��A�s=j�a��r5]`h;�_�b������.മ���;*���*���1��j=� ����x�SH�ڳ�7b�Z��$3k��5UR��N��1:W�w� ���ui<��슟��6!*H�+�����_���;�Yؖ��2����ѺxuǙ�P�*�0P��ps^}�(��ו�{�͊�Pp9���шw�{���{b�%�����J�ٱ�N��#(���GARF$�,��`_��l��GL�L�����
%�|������@�5�6
�D�zi�W0�/�|eͪ�.e/d\of��D�g�qp}
L�rHy!@�!6+D$*#f�R. �77HP�����u�2���4p�3�fq���j���U���Y�_\C�?M��r�/��L�^FB;~tiR���'��)����/��%�;ɖ3�qs����l���,cG�kPGd��Oi>��@��bQ����i��L��1����_�0T����
�+A{91��ڥ4� ^<,�V��-�t"}�����`��	j��`��M��;r<�g�o�p."��;�6M��_W���,�n��EW""1r��qϤ`��C+�F�zލ^��ĳ��ki��v$՝�q�pW9�gn�4$i�����e�ZN�.����J:A���/���e�K���;��&��R���9�R�Q��;t��ᖰgRv]��GB�C"�'x�Czz�7�.���w�d�w)�߇��{�ح�s�en�:��gAT�M"|�v���*���9	i�yP�p�d��!�Xo���������;Q�� �5$k��:��-m�"�j�AK��o�P�Ş�{V:�6������M�bý9c�RL�^�/|�W�1�{a�����=li�a�W��^�E>3��N��gV�8�W�?�%{|(���Jm#����Kğ$U��G����ÜY��F���tÓ�Ђ��r;���]W�]�#�^BC�5�ZԮ��h����<a���+�	�Xż3T�e�{��R��y��/n�{�7+V5�h��6��p��G��tZ�s�(@�Ο6��8Y�!��-��\���k`ۻV�2	cվ��eq���=7��ϨP��͛R4r�"o�^sބ�D��j�̥2���~�׉:Vv��l�;��[6�7�M��7�Us��ut���^s������@{�B�G����-��� ��B)�����֌�z���#E�F��U�p
;`����]���<N��	��1F�����۳����֮V�ɐ�Y|�pĸZIAl�/o��	�s��6�B>�hU""����DV&FW&�N�.�5�&vTf��Ӂ]�~�   �F�Ne�<:/�u�����r�\T��.0]�U}ҋ;��_��㻻2��������6Ϸ{�̾�JZ��#ɿ��x�7�}�Ys�ȧ��� ڧ�B'3����s^�ܣ�X��w���l/,ʴ.T\�77ȤF�e�WA"i��ɻ��ry����q*�<R�w\ ���N~(@�N3�u��Ѵ��@��bR��L6伋��4r�����Vڇ<�V�c��ߊ�L��Lo��W�����W��/�Ǖ�DJe��j��Һ�Ž�5}N��&| @y������^D�!��h��X�p7�1{xsVu�5���%�cz�/�]��ש���P�.X��f�u�����7��Q�Ae���2>��M>O�=�ķ��2�	q�0�lX�ݎ��c�2L ��ʶK��Ж��|�5W��A޿��-;��#���|@����~{��YHF߶����hD�oj9T�*��S�U�ɣ<|;L�w�E�l�Lw�@=�3��\U��P��O>j��k� m�<��o�0�{T-Yk��O6^	�t2��慳M�+��Du��{�|��W��������d�@|3{�[��^Q�֫.R�(�]Yǲ�ŕ1|�ׁ�u���$�V�m���`���]%'^]d,W3P�#+9!�r.�R�{�����ַ��2Y���X{��[�=8�
C �཰X4�])<3��|������Jͼ��t����߂�-�vC�贵s^�����z��ƾ,m���(��a`�wu8����k��EYꁰ�*,l�=~��D{���d[���`�R}��)q`2+�*�oEn����ڻ�|�LR�1T���?v>˫�z�̄��O��#X�nY�}�TV�9�tf���<���}a��`z��I¼h��A!�65˱u���Ņ`Nù|Pki~�.ng.�0s�t*ވCD->�,���6�נ�:�q����C`�����㋫��"���u�9�}��ޚ2\�F�P!8!��GJ�1s]��aֹ��)M�i���N�<}Ի%��b��Ϫ���qa�8!�[S�U0��{{|j6j�V��}}��2j�s���`h��b������x;ʁ�D��}^,Fm�����2��G�������7)Y~�K0�v��r6"P�5��QaS1�8�%^��Bp��mp������Dy+��	u����B�O�F�)�a��ȼ���8��^@�Q��i�k�ضri�>Y�A!h<y{m�ι[ST3;f�Z��=����qj��mo��[��j�3O�R��;]`L��aq�+�ޝ�V���;���+JK���$,�D��^�z�.���iA���_NA�t�*���"���I�����e{?#+�R'��ƧϞo=C#"��G�2�捣F�ncBg`F�1�Г:-vv+y�j�`��tmC=�-)��t��7��5�W����gǁ�үw�iW{h�t�.i�1��w��ܨ����Cjh�;[#�4M6ӱ��#�����Pi�OCA�̼��ʓY�l�f��C����ca�[�����ؿ6,�Xѽ-��yOB9����t��wj��B#�HaM{6��'����N*��=a;訷
�p�a%��*�.��sd�7�[��8(�kʭ�4~�-�YHi�N$�)l��BŴ�+^F�J�ͫ��zۣ��Ճ���'Û�`����[���Ӿc�Ar��\�l{�Î��sguF�x�cP`���q��|<���aw���N'�%����dڐ�ɬ��d8�p�T�Nm��B.�o����~�栋H�*�.�Q���F�V)�7�T	�*��+�ma�}��+UX�ތ<!��b����)B��+w9=��>�r��c�Ј��.1��s3�7���gARA��O$x���ǵ��k�������Us��Ln�wa.�&\��'f�6���g�|���c������6����ݽ�,Ñ��Y}�;����7�����.Q�����= ��r*�>��BsP�}�8��d��?Y���vc�47����`�1o��T�FӀvwd;�K�z��z�__�\|Q/��u���YAsb������A���
@L�Y�l���x����g�lL�Й�s	k|�r����d�/w����'���M�C�&��_W���+�oԺ��[unb+� �C��7�ɞۻc�Nq���^4l5����i �W����Uљ�񜄴ϼ��+ʽ���&�ֵ(g$�(�g�Q���b�L���g��*�����j�O�."�I�(JQ:���}Y�q?��p�<=�,��^L�{D���'�1�l:��7Ǳ�GF%с���/��rU\�y>��gR�8�@�~pWy��^ȣl�Ql�O��F��^0�ds՚�3U�V���!G{��H99;-X
���1���ޗ���7�C�Լ�N���Ą鼿IGXQ�+2^_��o}��f��v`SfK�\5N�O����f/o�,�W�/,��oFN��mP�d�m[�5ۨ���WF����Vs�j���\�bw�d;x��4�mh_e��!��J�.��p��sH �裚qa�>�b���҇3U"�y��\&����8]��̽�H{���N;���t�C�a�)RSP>ͮ�>�F�/i[��8�(��r>Y�4������r��7�t;����S��S��tmm_*Q'�����p�����]XL�O��y{ʍ�J~�l��N�y���r�+�̄�AsΙꗓ1�+c�Z�$���Q�4�W~D9�{���j��V�zt�2\��GEU�;������p��>t B��4�)Ok5Ea�������mVxW���ܽ����V�����$r�_�]�č�	�Lj��j�o������*���N.�:�)tz��8'�]j�\�3O/�a20���^�alE}����y��0|'z"gxϘ�,�_�i��	��,?Y}l�R���ϱmN�q�b�6���*��u�ޖ���	�{εaF�g�pS���g.W�����J�Y�V�.Ss]��i��ňvHw1�X	���5]���\�E������oAo�ٌ��5����61��Й���~�އ"l�Ţ��ˋ�N�<�ފ�0r��7�o�����VµJ����Ǌ��w����@E�jؠ��O.��ܡ��K�y���5t�2��IE6�N-[�&Tq���yv��έ����.�Ҭo�V	�A�_���]9��A�T:�:�7��`F�% ��7���Rf�y��׵>p[����h��q��{a�%o�[�?K>�I#��(6���Δ��>��V�?}��e%��ᅻ�F=Y&s|�a�J����rj�1�%�O{6y�>���i�J�T��'=O��Lal�^B6�����o�;q�o�\�|��ބ}�u���b�"�g��h�����W	n����pE����z��jf� iw��7��5@l<>X�Xo���u�
C;�����_���÷c���@�/_p��FR3>cr�eX�E��q�^�S�s^������8�X�c�8~���=6t�����=��!����͋k�V�G_�"�ܾ;(�F�aK�3�8����F���F�]NFd�
��(�t���Y��{�A)��=�������ӹ5��ɧ2�mc�T�J*t
�����i9I�h��R��a�/`V�W�%�Ѿ�*�1��;�fG{U.!�������!�7�ڡ�ACP��yB0� ����))2������*��r�C� z��9�J���K�g�U���}�3���,�Z ZǛ�0����z�y:�_��&/-J��y���t�a=�-��ь�}������IҚ�(ȝ�	r�����U��KX[�[��b*�f�Y�_�[U)0m��H�$AڹA^Za�:E��p�K�(�[���7s4
惥�%�~0P�cc�6�����S��y j������K�����$��P��8����4r\F��V,��mǛ��|�h���/����FiW����,�����u�V�#fI�B�7�m*����j�*��罆nSw��уxnǽEU�(�I	�Ș��;.d�%�Jyv4�9���K�-���h=R�RF��rI�:�s �S�5}}�HKq5����6U]�\�Q�<M��՛b�;{+iUt� s��M�	K�\�.�<��3w+�7�8�
a�j���*��'T\���9v�t���§C�I!p��d�q�'�׮(8��q�ԍY�=D{bc:�w(�Jo��ٌ���̷L�zb������^�.U�V.���vS<��œ[�m;�M���@����kG�}&�͌^�h�@��.�ORY�!ݖ]Y��a�x�kw��6مM��Y7���x��>#Z�<jm雾崆��춀��ʝA�/��:'��,��A�s��*�
�|�e=��x�c(i�	�<;u�;r����=n�&�e��Y0�.��!d��E��ddoYWf�M�t�5JM�흭�x��ʝwe8*�w�u�� �į�@�/Rϩ�t\FyT�x�9|����wv�OK��;�.͝�����հ黣OC�Ut��Y��{$Z��K��_�<s�(�8V���w)9ma�����ǛZ�D�76V���AG*	$�Պ(S��;��źv�������&��7FC�h������Y��gR�[;�s��w��	p^1G�Q�Ꞙl��┞'�����7�ܤ�?d�5�]�ި��"t�����YJ��+��^Q�p�N}�惆�H���Z" h$�����&�w�H
:��Q/+��=Vk[W�Q��ZOt.z�	/%�p�d��0�+ؼo�\��c�=��$0l��Vԫ]�|ҾM�R���wkJ$]��6{ ���9����1�n�a^M��ֹ�#��J]+�m*�_���%
����Z�L�}'��is�6�K������9),ee��Cb#��pvi����;�����XR�E��61[��+��,�3J�+�	�įj��;�_KJ��ШZޤz�26N���Q���7B���L1�8LІ AS���MvQt�^���� ��S�<�&5�T����=)f-���o;�� �uǨ�$�K]9->na����[�������߽��EE��QF"�>ҋ=�Ԋ
���T�@V�1�TQTX�+b0��QV�KJ��$TQAEUҪ����TArʶآ""��j��DV*�X6�`��eAT��DQ��b����b�h�ĬU�Q\�*"�TE�����r�S��QDDDPX"�fb�b(���Tb*��DD��bF����Fe,KJ�U����Y��%h#UB��1+Aq
�Ң
�E�*�J1��e�TTQb��+
�\��Kl�����&$*
�""��QTF"�DE�QH(�Dn\eB�bJ��i���X�YZ�b"9h���Q��1+kS-\�VV���r�b1QI��Jت����AIQ�UEXֱ`��TF��-��ڵZ( ��D\�81-(���AF��"�-U��#Z�R���*��-eTAE�T�b�Pm��(��-��*�ږ!�`��b����%ه�׫��1�z�ƙ푔�r����WsE^��0��=���e���8ymĆ;}������^-�lA��Pf��_��B�x�� ��`��j≊���O��~~d{}�\�j,�!��:����E���=	ˋ�pE��꘰h8�ySG������C�dt2v�����ۗ�����h~����Z-w��z߁���+|��Ń�>%b}�E��ދu�E5i��������3�̭��(~�&"G5���o��\�M�]��2��[��m��Փ25�4ϊj�u���U��_�q��9�:�fG��T;)�9y�dV�\r�����/�5�~�1�����(Ѱ*���Ss�6�!n���M(�R_V��5�}�������h8��F�L��Z#�w7��4W�VeG��N�i�b���X�T�d����!ߕ�C��Agyi���*{�Y�s1��5�i
��-�qp�3�J�Z{���*�S���6�I!�#�CR!c##[��]���}��;U�V�#=�qs��>�	�Q�E�)}����p�x��ڭ m�����l�b���GԞuڡi=�VVii��LC�J�̃�?����7�hb�=�	�����qF��)��0��t51��h�v�©��t{�7t�FhѽeF�μ�Oj�-�6��O�<���R����K��e�玼o)���T,�b�\�;�˓������&��.�0���YJ��l���zkʅ�P}s�FQ���q%ag����Z�Y�n7�j��uJyBR٠�O��P�'7����ɂ�4ϫ�z�?��s<���X�o\T=��eF�C���S����K`PD6WH���K�l��|-W!Ǐ�Kש*W�38�%�3٦-4|�k93С���i�ϗ�Մc�!�u|�4b��Ig���+`���x�2�;��J�l��'!�9s��Vd'58�E/'!���ݳ��Rx{�i���<�'VR�|j�缅�D���D�ޚt���:!C����~C2���8{�rm�f������
_	sK3�W��@p�*���g�l�`���p���;���~>g��;�Z��$�9��nZa�l��/��9J��]CY/�u�M^)�S���=��n.땀\e1s|�b�S}�)x=#Aگ+�Ȫ�͟�L���Θ������&Od�X{Q^�tK�w�`��S��h��{��VF�v���]�/ʇr/u`��k��S��}�Q&����MWkb|��O�1���*���_Q��\����bpr��^7}r�	u�K:�xO���h(D�@|��WǛ��[�Cfb�P��≚vĞ[�������P^RN$�G��FN��J���yZ��W�^g�>��1Wj��6���5���~L�^�.��1�1��u2��k�f�͠y�\�eT��y��E��1���
!�r�8]L�HprEF)���`4�72�n�en4�k}5Epܩb�N�ᒷ�q�q�p[��gZ�k�U]�c��K�`�{����}�xU
�kx:ļ�4���m����Om3U�y�M�,����DN����~�k��������~�]R@�
P{&��l���hQ�)=2��-���x`���K�m-hܓ{�ז�B�]��1ѵ��TO[��!W�@D#ׂ,WVD[�:�}�m4�U����[�/޹���7��o�j6�9���(�83�/ ���[B�HH�֓��K>D�����C�с�g`e�~2\��GF�ɝ���T�tK���"(����^޻�i��y��B�����Xx�W��u8FF�ʜa��Ĩ���m��ϲw�7�pj�|���zg�Q'�L@|@�.4y{�����>��k�Wt.�(�ȅ�7,l5���LMS
.��T�b��2�����~��5k�'�����o����.&��ι��vSd�Y<�iǸ��oa�˪S�b9z��3P�����nq9Ȯ��us]��v�Af+H2�R���2�;���)R����oh�m���#��}V��6Ox������ri�\a�xU+���z��j̯Z�	�T�@m�LT����0i�6
��
����vz�2k�YE�*jQ�h-�t��.k,�ྊ�!&���(B�B�L��X	留WC0���W,�1nF�fvj��V��Q6�}%P��Sz<�~��3k�ț1�-��b������ѓ'�a�ﰻx��lX�g�FPB2)��f�^����7��S�uk�sڕKR��΁��K֖��v	0ܻ�8h\��m����
o�l;J����X�^!v�N����_�υ[������$�������[=B6��s}�@-���Qq��'�Gޫ=ױ�x�b���3�Kx/����,�|v+���P��`O>w1Yt�t��k�σ��Z�X��ʈR�F��U+=���&��ґ��%�#�e^r\j��=a'(NyPǱ�l���.��n����-OJ��]a�Q$<B�C��{�c"��
�y 	Q�jn��:�+gP���pN�Db��o�#���+�����Y���	Q߳{���ݶ��)�ꙸ���e�uݾ;���oMT��N)�Z��gn�X���;8�I~I����j1|�8�`�f��u�  �mޭ��_d���П,#��4tӅ�����}Jdrt���`�Gԯ���W�.n�P�:�b��=h66р7�צ}�����V��BSc���c�&���1�<�jxD3	^)�`F�.�^��p>��I�>6�4G�qo�ާ�*�jiOuu�ᢼ/l��Gb����y��a�vu%�Ұ��U u�a��� ru1<K��8��`'�F���C���7���Zd�J��O�<r�����,��챻��/e��2�b)9���zϪ���qa�8!�X�����h�����~]��&���\���j&]�EZ*<tm&*[�خ�b<�'8 ��G;qB$v��=�<�!n+r��j�4�@��UC.^x�F����#oi܂6b:�9�o0TXT�d�mgk�֧����+�Ot���HH7DaMY�X��,W:2�S�����l�Ҡ�����:��j9k��gf��xj�x��j'�������(Ѻ��Jo�Yc<��\��w~�۬�(n��5����=�K��ݯ���=�T�q�v9T�T3�Y��l>ZQz<)TD�rj�n�~e�{�ެ��D�K1u�I��9�ƽի�zs"����BL� �Ѣ�px�ʊ#���-�ۤ�gm���gt� s�{�G2��df!��r�3��_��6-Hc��Bm�>�-&�˟Q����&���:p{J!�Wy9�q���Cjh��ؒ�9~�&��sE[ع��F��2lw��?\L�ME����;!D"H"V;ݞ���}~�uv �P8ޞnp��){�syZs,:���J��E������4��^16��H|�%�,�5K@�t]���;7꤮g��4b�=�pPoMyP������z�P�9K���~K�ވ��W��]+�g����"�LjS�xt��.`���4��0
��+z�;���6��g���bZտ{@:��[�f�#ثS���t�$,lM�>&�4!.l���/�o���ncL�J��ۥ7�0Mt>���Ud�l�w,������qa��b��Z[W����'�y�#�y$�\Գ���u�r�uϯω�7	ɊYQD'!�U��)��B���'p��˨�q��f+��-�0c�b�C�c"��Zl{�0�P؎F��Ӷ4��%�A7m���R�+Hb�s��AuAn�[ݛ*���vֱ�ĝYs��;Ԍ���x�5;�j@	�C�K���ad�S���z�o���t^�Dy�z�{KgH�`)�%a�d<����kU��{w 9��~J�]�˴4}�ޏ�N�L}�O�p��M2���1gԀ�%�g�~�5�l焟5�P���k�r����н�y�/gp>��KU�����hu�M�}��[��[�.���ۨ�Zs��'J��R����-���X�4l5���D	j��謇�WFa�f�Zs�n��O�&\QW/��1j�yk�� &@�<���e� ��T��XE������!�(���A����Q}j�|N���EBY!�6Y��~L״0�Ϸ���x�r{a���D5�7�7{�n�J�l��D�oB�gܯ�\]�Έq{"���n��=�$�j�9J��ٌ�?n��<ٶ�ǆJ�P�Wk��}k���^��{w:;\or�Fv�;a��v����d�Hc�T��-`~bu&�z�����On09�xf���]�g���$<�{�}�66U���c�t�xƇ����|���a�G�'�W3�mz���c�M�ڝv�<�C����{}|�������=c}g����e�Q"�ة����:�-�2�芝YF({(��l�,��.��-(t���Cfp�Y���d=\��w�Z}��[�LoC^�t�������<����V6a削�����\	]�L�m���[��'�LVU�D���/�A��ˎ	ۈ�W6��vf=5ֱn��w;��Ӑ��*��@��
��/os ��E��L�K���ж:¶L@>o�rk��9K��Qb�aA��z�;̗:���Z�&v,bg*o��1,*q[1��������)�=��!خ�\x�u���yC��}�Sy���>��31f�w�)8:q<B3+sTP�#�B��D�]L@���>��|,��e���/�+�q{�l-.|�x�ϦKm���#j���+F��3*�`�υ.0�o�U������?dk��E�WZ��]qsϫ��U5!؇D� �zXj�?#�8�y֬"�h�`MdQ��ŗ��Cj�P�q�!T�L�>�a-���
�L��Lk..у����)�F��E�v�Q&�^T�7��z��Y��64MB	��,f���^D�!��-�SU�eZS�J{ՙ��!��&db?��x����v}G�A�2K�/��(1����FI;�����V�Vf&���"���EE{v+�?1���˹�\��m�p��C��pW�k
��9�`�of�쐺9�����˧�_&}B�Bє�6dĖ]�~֥�,�&ֹyx�}I关F�J�!��W�p敬�Kq��%��rX��v�=�=���;���z�f�T⎠�r�$�o���3\�C��pҸ��EP�B2�ڧ����F�u�����_]�>�Ж���SS��pg/�Vñ�	�E��4�m���#�����w����)���}RQ�Ζsw��H��Ę����(��b��Kp���.����Ʊ�<簭݇��=��)��(���Py;��Zʊ�F�	���{`�`�]E+�U]���\|.-�ڟ/���B���|��WE��*�Eu�ݨ��
2�US%m��n5H��4��*Q� �����hb���?�V�GZd[���`�����*�S��Z9�%/&p�K����P�5J �z��������΂R�~�q7�q�/����`�r�� 뢣�@�Sa�>�:M'('����0R���sɺ�R��|��lA�ٸ���a\�;�m>!>�?5=�>3���O7��S�K��]l�h�Q��y��]�{7L�w�z�GA�6�.;|��4/%��iE�L��S5J-�\$�Yg3�By�<O��u�ld�
�>̧�Ϫ��7.,:'_�g�b�����v,{�'�=i�r>K�r
]^�ՌŹ,j���>\���!s"��l�k0P��~�[�t���t$,E�d�Y|�}`��y��kN�b�o���Z�t�����(g�v�ǿt��o��˂t�ͽ�Q��U�\�WxT�7VC���D�'�N�qL)�\���ǒ�j������r�X/K�4m2����<K�!9�s���8��=Z�erq5Z��
"͟ �K�#�w�ř����Ȉ���Cn!����ڔ��7���u{�dY)��I!'�� �+3��F�Y��N2��=�Z���#�-{���-n�x�\E3t��cg�qB5���{Dƣ��+�1f˪��߼���!�wsi�q��X;�!�+�s�� �c����P��KJp,lA�7� ���i�֣M �6�`���juZ��C�X dt!3i�;]�;N����!m=��O��,�{����ݶ�����{�n���q&2.>̾g�{d(�@D5 �+�����>�G_o.Ķ��:u���n���*;����ޕ��Ŝ��8z�8r�A��V���U�x��bv��H����r�%�V�`��Na�~p��ޚ�o���\@�ةy�6�K������Q�m�{���Î�
2[�_��	��W*&y����C�=���Al%�E��AM]p�ï3lnpI�QZ��N��������'.�dq�9��o.�w4f��8h���X{Ts&����[q�t\u#̀��]�����	��)f2ُ
��0�U��ҫ�|a��2�O
8޻Ica�OZ��7��e�Le�j��A�/S�z��x<M�]�uӬr#��/a�9-z�Q�jo�W�9�.@fc���'>	A��`8�W�]��8��L'"�BL�'�V� �<�_j�Bk~"���%�+�1/���m6�3=H]�-�˹z�4��;m�3f��,����r������{�����ES'qjQ����I�ct��g%��;n��+��Pn@�V�\�JB��d��<�v�z!�N���y�(��책���l�wJm���Յ�xz����oE�VY��ߗU�J�y��}nOíV�;���:`tn�`>�j�;	�������e�
���:�3�܊R`X�$�qa,?�վbw6���SB�NM��*ܤ��-ͮo��.��H	����N��hឣ��U�;ׄ�j�.��V�d�%����y$@�nx��������)���0�����C�i�l[���T���UU�Z��,��H}o��`|~�7Ҩ���B��	�N ��q�����Z��A�-Kö�R�
6�6��`�.��wx�Ŋ�3R�c�Ou�B�M�{@��U�Q�{�K/��DUX�G�b�~�Fx:����	�g�/|�07�wE�+Nh�ܮP��6�k�Q=�l���Cϭ��z�<o_U͉��G�1���`���P���<Wd�݆��޽�rJ��3:�b�*I�$�6ޝc��Ljɗ��
$�]Lb��ל�2S˦�X�K,P��{{$����� �x�9Cۓ,�ݠ*�[��]ԲԮY��p*��b�w��.������z>���^�A����Z�N_��Gx�w9G'�{ӹۮ�O.]�x����o'pV�[	�8��\t���gL�a;��۶�:��{��4�:���T�7p{k˱��bĊ������jd2�n��P�ʕ�9�y��sZ��b�&9}���f���i����]����ݏ�$:5.&�U�*���"���=�����i4��W]�;�f��
�D�% ��*
�3��{j�rb��D�5��o5�%��2�j6�b�di[.*�����"e�w��yT# ���Dޙ��>�Rt�GQ������=�
�½�n��D;,I��j��	�ݯ����eΣXs���?5��[Z�u�\{|7�.M�\Z�����c�=1�Su�[��?���%�zA)�*�=Z�AY�z�ٌ��:#��ۑ@����lc��\�Jsx,��^�9��6�l��XP��L�s�z�m=�~��5�����hUV�b��U�Z�*�J�*X��E�Ʋ�F(���U���B��-k��� ���V1Q�%�s2,&\�b(�*˘�j�մ�+[[`���(�8���h����EUm�k�EQU��cZ���!ZKJ��e�(�`�QR�Yڋ�1����
�DD`��eZ�,P�UU-Z�֊V�EV*��X�աQ*���lQ���b��U�mF��EF�J�kR"�h*(���-�J֊�,�Z�����F�A�Z �mUEA+-�--�
Ԫ֍��EKEV
�յ�DQ�UXT���*�-l+%�T���֢��B���Tb(�J�+-J*�V�AB��QIiA�U��)KD�Zѕ�keX�(�$h�V�EE*TekDmZ�mX*��F������'�%�� �R]jx�ªyͪ�m[�:�:��c��h2��P�l��m��Is�Kp�;=�*t�..�s�d۽��.�H��_�[��y#�_��;�~8Я�!��C>�P}8�T�j��O�0u�҂7u�<���H�Md7�u�im�ԙ�Wt��ן������+oMC>,Ufk�M���b�ӠGO@���\���*�9�:���lBrKuN,Zg&v���^w��ͮ���6~����Le�4<��у�����fy�����}܌�ȧ��ESvG<��D����!�>�K|Y��Oжs�D�(��n�^ǀ{2�z����=�w�(j�C�L�EM��DC��"��:�&�����-�R��R��,3]¢����+��<���Q�1��0=`��^捆��bg��i �S�3�.�TO*��R-�^X��Țم�xjf�e&|0k'������ ��8����g��*�Մv�����=y��9�wv�����R`L1�ቛ,��?&`�h�� �O�x�s��f���Ϛ�
�5���U�0���0�e
!�_�.�o'}��)����l�um�sK���^hT��v�*�w�z�0�q��vh9Wi�IW3�������q9
�hU�8��׻\�}�o�s�܍`/���xq�}.�5�$=�ؑc��==��������������6bq�ýB\R�Œ��o
�z\�Shr\���^״�}+ޡ���[���=�P+q��G���~R?M�VT�ƺ����@�b�CbNNӠc*��0�&���B��鍅�k�ɶ�*Y��\���ν��aT���ix�P��>|fڠ���m
='��#�~�smhNFLt�����U�Sv�e2�^zf:6���(�n��^��^��`E����ܓƳ�;Q���ٵ ���m�Ê�(�83�/��9����kG,����,�m��FjD��NQ�4+^��#b�Y�cN�� �~]�Do���]�AEP�w=�u�h�8��DP��b:�$!5!ه��M����b�y���]�j�m�e����۾2�Y��az|���`�I��:��7���q�����Q��˓R�T�՝]��E��1lz�_��#T�hE�F���,�8��$�����.7縲�ᠮ�qq|����ȣWW�ؕu�)�]e9|!рLੲ�Ă T��v-lC���!��r���5�/�!������FU����K��,����������V��'ܡm�Gz��P�ڰ�s�h��5G���O�\D�ΊB�[����T>�k|F7�������>u�����3�Z%X��uW.�\'vvڮ2�DF���G��ӻ�G��:A����yW��{�a-��<P(z�0o�=��u]F����9w�V�0����Υ�,ݓ��4t�������C6xg�އ"lUS'mnh�C��J�b����^68�7��a��O����X�<�(n�xώ7^�zX��R�[��(��1�n:I�"��K,_�Ơ�a�_�a��p�l�٨��Be� �U�DE�X��鸜��{7�v�Jn^����zV����I��0�o�lOzi����I�j�Sq�k��-ԡYJ�!�P�Mþ\�jg:I���<���FA�g��7�O;z�Oğ'�e�������x��`etB��L@(��Ī'a�]S�YQ�5b�fӫ~�K�T��Y-�}��𷼛y�b��]-��Z�/��g����NÂ%���;*�Eu��D�ތ]uG�)���-��\%(3�.�Hۡ��f��%���is�M5�)�hN�7��L�rY͚>�D�WgT�B�%����>�C�ƃ�zScm�|@Mz~���к��_2���f�E]�F�U���(�sq֞{�5t��3mwdl���f��y��3%�
��<P#��(y߹����'�y�f�A�Jy������
�P��Sok��`�l�1N�|跃#��܉�W�ɜPw
�@~[�"�,�X3�u���5Gm�:��Mv!>V�WG�޷���Ν�<�z*�@�Sb�C��荱4�\l(�rʳ�+�Cջ���t��E.S3�⌦.�2ذ�a��T�H�;��O��>=�C<ޓj��AU�.�$,��������)c���cӞWHa�Ca�+����B�\�F�PN(5�#g��+'.��{�'��U����ˆxdD	s�̧�Ϫ:�j�Gy�z�*G��ݺ�G7ρ'�����f���l/�E�q�h(#&*[�q�=T�{!x*�����dyڧ��ǁ	�˳��[�3�غ]qٸ�x�[:	��HLD��`�-fٷݞRbn�ۇx�=�G�����J{�I	>�<aMY���"��9�vT�n����\J�:�v��Q���� ǘو��e;�1���b5>�O��4�����f����%Ͱ��Y2v��q��n�����#��+�/��,lZ��7��&�#�/�_��/3��3)���Vj�D�p��Q��C�茍��Cjh��ǽGn,�מjg,��G�h�[�22�ҭڱ�쨯3J�c�]R�v+<f�]��n�f&���s������B�
������Wp��EC���|ݾ�fͭ&9;O ��(���aT��0X9�O�i���fi��V��\��I�&Z�W���p��Y�B�j��&2-<��>S�zt�'˯�0���iz4q:�9m5�!*�gzً����ĵGT(��_a`N�h8rw�M�4�U3��u���s+)��*�#J�fv��w�Pm�g�\h�8��d��^_�n#�� U7�q��e��Y�#uF�t+���'Mޑ_�;��{æ��Dޛ�w�2��ʑ�^��3�����<i�_z��|�e��rU/d\|�S�K��C`��*�FM�Y������㎖b��D=g��ɵ!����mW����=K��3]�>z��\X@�����uR/v��.v��|�h�OX��� ��\�����#�}o��7	ɊV+��1����{�W�E�^N�g�;�7����|����c�bhcK}鄯d��={|�Eh���ۈn(�F
���~�¢���\X�<U_�b�t"sT���ǵsr���&�"=o�_��}�vK[<�%����&��&�>���nr��}ͬ��P��D�qj M-y�<l���j/�>��؇�V����x;��|*��G`+��)�Utj��ϮsJ.���}�$��5���٪f��p��i����ܫ�`�3q.lZ�ٜ�#NoEY9�R�2ؗϠFkʹ�@j�_q�	N��Rt5kZ��~�Ȗ��?
U���a����U?	�@�v�ɚ"�w['�ץ�o����
���.��"��t��E���e��5�L=�x"3�y�[DC�|�M�%��mu�.�"��ܡ�Y�X�<| ͖z�0��[�}$g�]��lB�]Pڷ�^f��/�^C���ݛ~l齻�\�8�B�
!�����qw�#��TY�G�=Y�x���Z��ϻa����P>ٶ����+ޡƾ���-��Z���D.�P8T�q�"{�p�Wh�
�u��?��j�����Cm���ԝ��d��T�{�*��8b�g��=�2��U��נ/=��/D��|F��m��(�6z��Y�k�J6ˎi�N}���t��#֧��Z���V��3[W�T�M�>��^�r;��j�mQW	0�)m�97��>�z�Ks�6�j�~�\�)ҋs��ꗓ1�7Ì��n�/N$'�1{c�1�&-�AǊ0�0����������@_z[Y����UyF���9y(%���.��-�Cx�S����{F�~��^ۍ�	���W_�S,��9�,���Y�nyk�F�K��z���F�f��Y�m4�a<�W�W�@�F����2ЩIgJ�w�t-#](��o�:YEgc�㓞^o0����V\ǽ�x.���~7<\��-1
�d���Y"8�(��yNX�z��65�)�|9�;);�V�gg@��xf�r7,Ϧ���F��:��7����.6�xT��R[<����₯��b��.z���б/Z`�WFL���,�\��b�k����M��:�<u��o�躾��T܇b ��
�*�H>�
��_N��A7�^#�rIwۼ�r�K�V��~Waq��'�̈́�3g��(z�0o�k�ˊ��b��]7�{��9G\\?S�W�f+��q\��3�|�������myN��L�Oz�qk<&i.���Ⱥ2�^�����]��W�>�2�^�.X2֚j�UӅ��<�����)(oP��%�/��Q�ӽ�.��Y��{)ʇ/�Ц9}�p�ך��(���c��a*vb��MD�1MA�P��I��������M:�[��G����Nd*U�C�.�4�0�<�Z9�L�dl�r�/�W� Ⱦ�j�GVv`�U��[P��L6h�F��vr�(� �{E�,w��+�����}��[�b��,ȅf���9{l����2eCs��H�gV���]t��}2����竆{��p�n�f�K���B�}�
{P�j��y��KKAY�!'5GG�z�tO������#�;���*!K��ҕx�h;�=횕΅N��ʮh��S�Â��\���'����"v,�����fH��r��U
����7P�v��g�P/��+��s�u8D����0��Z�ň���
z(6"\pDJ�J"����������у��5KB���[�P�.�!�e�Ӡ-������p��ڕE�[(��h�M>�U�6�^�Y��ݮYB�tE�d����WO�m_?Su��T-�S�1\j�=G5gt�]	V��g(�fAEH�'��Ђf�iGs}(U+�*T�j>�����;U<�q$cOdgR��ȧ5��/�H����P��ۀ��u{x�"��\�oF��pKgݵ@u0�p�v`D`G:��1bb��_�,O'#%ff��Ve�8�Gdh�:2��t��V��O��b�!��R�#X/����@G_k+4�f��9����9��Иo��v���z3z�1+uYՐw��V�]A���E�:q�
�W[.��/0{�x�nK����fnS�v�H��L�D��&�)k���Áoy��J��m��<WR���-��89�SC^��[�̫���TF�J�Q�<����Rt����91����q^|6h	{���	��A�Y���^���k�95�־��6��lg�c!u:"�ޓ�΀Ѝ�ç�%���2�>S[�d�N�u��F4+5������{T�aTI�V^jx�q}�uS�2��A�w��rQ���A��A"����-�MvV�ƭ,j�5��:q��+p6K�~��|.v�P|}�#�f����C�<���q�K��w�LE��Q�;�>���v+�p	���ή����)�/�SW�xXSN�<X�P�Ӈ�J�l.!P����|%X�x�9Y���{[�]��רwu�/�ww�8�|W9y.�����
��7r5�H���u;k=C�F�9����muƱ�ܑiA��(;X��.g6m^3]�چ4�p�5��YY�3�.�-��[i���޾=��]�C�*<�	���B({��> L>A�ΔĻl,G�j��HJw��ݮ�Ⱥ�7z-���X�&�z��:��c
��˓L�Ռ-'{�,T�9�Zk�G�I�X�(`PgM���H^�O۾�|%p�%��[O_�Uc�Xվ9LOB�u��T�{�1=��=*y@x���]
�H�����v�x�\ບ¥�5��S����k�pO$NP���t.N)8���=Y�v�7r%�Wvbh���P��젘���	>��P���g�anI�1)�}7s2{�Q�ZUS��Bgy�D&,����6L����[1v�n�њ����8��9�&q�G��n�>�籉�Lg1uX5�RTb�T�ܤ��.u��(�G��Y��9J��-��Z��o��^i��e�tF5��Y��#Ro*X7�7�M	{��չ^�yr��4(aA�ʫ�,�z��9�n �	Ux�;^��Q�k͋�§%w]]eQo����7�j�3��G:J�OE�vow澾���+}/��_AK=�c����Ut黴�� o����вu�$�����L��?[��$�N��J��κ5�d�$m@�����+1�Z�1��Q�A����(��F�K�r�N���T�����f�ݴ��)�_ �6��pY}���\�ތ�4,V���sh�tMU�Yų{4���2g+�f�9	\Bmػ&<|hd�T�O��"�)Ӵ�a���2}�E�i��4�ڗ���+�6G ��
"�)�Ef��N��;-��[�V!�[�93V�Y{�5{�5z
u{S2��S^13�`�{&�����w|���,�1�����g���x���������.�{��t���, �4�o�U_@��c�u�m_��m�B=g�a�ǌ���Z���wQ�S�����}h��� ��c'r��>,҆���b�}u���I�Kp��]���u��S�Z�;���vy��}|��i�+�]#H��S���ޭc
5RK+Fp������tqa�S��.�P|�ɏ�fwq��'Z�4����~��T�Z�:�1.�,����줹��X�"�qv�gb	�gh[��'3��
77nE��[�rN���7���l��60���Զ΍ѷP��c�9p胧�D�	��ֻ�-cQ��N1|8��N,M'U� *K�#re�9��{��7���m��Fᣒ��.G��(��o��YEi�aW��_��n�q2�~��2;Ѣ!�k]Oz�ǯ��B��^ēS�2}���B��k�f�4n��V��v]�N��z�CO��k�9�",��y�'.%1�Y�����o6DOgP���GAa�څv�N��_]p�,�j�L<���,��ٮW#�]�y�WB�sOitҡ��*�mk��lޛ�UD�)L&m������c�Ǿ���6�ط,�9~tC�bnuUn��ΐ�⭮n-hkKv�<�ɂ������6��ij���J���j+���=�[��P��iW��V��p�j�=�Wu
Q�^���c�o�t&$��w�*�M���Q@��W�6�z�k<�����;�B�����edG`��9��0N�2E�F����O(Qw�9'��YkC;|����|A)g+����r��W��ȬSk/c���9N�[R�ݖ�Vx{P(�h.e�������l��Qە؄�	b_���<�P)g�I�����j0��֎J���F��C��'P��5k7V-�HLK�|��la����8C�o'`
�񥻷����_\��X9�4����JG�_E�N�Ds�b��Y�w�O�5�@c��+��޲L���F��r�A�}�'���{x�Wo�AV�eԫ���}	�[�*��OX�6���C7�8?ԿX�}:���ǋss�	�k;���4�G����s*���a\f��=�n-�b��Pk������뾢^��fy�Þ�z#��7f5}��BU��������C*/k�޹{՝w�Z����k�D�s�'����Y�V�ڈ��hQ��KZ�"�Z؃AFE�-l�U�mDA��*Ek-�cch%Q����-���+�b�����l)jZ�-B��������P�Fڣ1h�F*��Kh�Klm��KZ��TQ(�mU�V�V�����ڭE��Jִ����b�b�Ѷ��Q-Z4�Ҷ�mi[k�m*�iJ���QU��X�Z
 ��Z*�լ�-)idJ2�[mm�QV����,E��Kj�����")[J%�������mXض�ZZ�5*�X����"��-kl-T[F�m���Ej+m-F ��R�Z֍�E��(�k�em�Ԡ��m�-mE`ֈ���c������z���N����oyVQ�WL��]�@AY'���=��MzcR�@��>��A#fq]W��2��q�ޅw(�rm�h���V�X�7�ҕx�K��%Ga��8g&24˅/v�5EXy���twav�zmCV��{go��.c`�XXA蹌�f�R�(�	�v�⺼	���58�rh���n��n�v\R��/_�K�IC܎eP�ȕ��+����%j}ݫ#t�2��3!TR�c;�?K>�S`�5�
�74��CB :�U���Yz�u��k��C�"l�{�<���n��Τ���-# �����5�f�P�p%��s�y��qwg��=�=Z�	V��8��EHN,����T�K1�2�T+u��a�eY�Y�������n�Ն���N ��X8Vơ�v���S}�rE��k�
>���[�����s$8��&�M�n�Q5Z�u�1�fkm�fP��t�#)�4J=C7�z߱���8���7���/?%��|�����{'�,T�l�1A���I�J�7���	��K��kw?;p��{�c��ф��A��_��fO�y�\�]�Z�R���}r�3�`��5�������5����J�_o.h�'
/\bwd'i��V�)�=Z�	�r��q�D��9�˵��ˣ��al7�z���;[���Ҿ�F��6����*�8٠%���ܫ��]7�o����9*�s���zCp3���P���9U=�ץk�D*����Z�������̛��TOj��#7�f����}�^�s��>y������V#X: Z���v�|�j�n]:T����Lq� �5�QH�X�[]<������EW�V����zÔ�s�vlU��p\���(>�b	�e��:а���f!D��y�r�b��TX�P�.�*����E��P\FWi�N8�9�K����>��/wa?,v�C��@l&e�}+�DQ����f'+�"7�J:O#3�G/{��c�:f]�=�lpzp�%^l[J��� ,�{���3)K����/[�����-wV�HЛ���5(��h��+��&��<��y�z���������no.Se��),�7��8ք �-��\s��K$=���y�i�f��Q�^����o�u�����$����Xz45)�Մw����ۗ��
Z������i��͕��54�Kx�:ݵNuX�k,���a���`�o�3�m3 ��2:�q��r�|�#ug��UK�]�G�A���=v.W�]���އ5bH_1uY���Rk��@�ʐ��m
�{C$���φ��pKg���T��v������]���F<����BP�D�e��Bۚ�Ҩ�e��x�9u��^Bj �
!�;�2��-F	�qMg�5��
̻V�9ͱ55���LęruƆ�D���پ~ۦ�vS�91�D�qU�L_��x��Q�K)l�����\���b���>包����ޓ~�;��w9�a>���ךƺ��d�e,�b��Ǟt�hW�Pdm�ʞn��SO�ח:�k�O���5/۵�:��Fk�)\m4/��<��Ү�62�J6R���aTZ�k�Nη�
��l"_�Ԉ����]#:��}B�.0E���j��'�ۆ�'�%��t��-���J���+ӻ�2�n�����[�r/��6#T-/� [g�N�!ݧ�AM^�.<��1o������)�t�f�w�,�m�xp��������-�n.PS��q;�S�=i���ʇb�)�x����
��Q�vp�,�:���z�8�W�k�}��=�\|�pEW`ٻHa��醖,]T�Ƽ����:��8��>��ܾSжɡn��zgz^ƀ����l̛�!1=����YZ����VGZfU�e8�S1*�Ҳ�A!S�˼�ｽ��aUP�մ��e*��cG�r:j�L'z1�(�=����2�R��YQ���V"a�81�ݦ�ur�U��yn�!o��IM�	Zy"S��U
��qءr�4����	�4�@�e&�6j�l�)���R'cx$�p(J�Me���8A$�ö��'���I�u.�tFqdh�Ћ�a	�-E��͒%fp;ev�Q�U�u-�AUN�U�ݿ]�*�`�l��@�s���&3���*6��>��#�ri2�;7���m��Įw:�r�P�(]"އx���a�A�J��E��wd�vp���IW+�Zw��40�M�x�cY��lfH�ê���X9��H�a=.d�4.;�co��Rw��±�%Y��vpi��<8b���>����7c��gwY�v��7G�HW��7�gk�k#�l'��_>��t_C{C[�	h/����7�TZ5�啧�/u:Y��%��m�9���~�|���j�������f�������]!���ofwEݗ+��
uԡX����n���]6	���՞�b�C�y�M[�}9�.cJ�x�q�pY���H,w�9���������z��0x�w�c�Srj�v``N_�^(>�p�Y	��KX��l��rQC{���*��'[WoD��n��m}����/����]��q8�V�Ј����A������^���?F%?�&S�g�m8d�Bk�����ow����F�a��iܟ6̻��������&;Q^��1L�n"2�rbN�=tUr~o���H�>M��\\&�dJ���(p/rN(�B�3S�R#{��/�s!�"#�Vc��o�]�5�с�*]�/�K��O*7y��Y6�'�7��{�HZf���>R��o�x���s}C\P�n�ܬ�|�l*'!�S.�����鑗���%O���4]�⑹���v���ߎ�V�S8��*rw��Y~�G��l�/��\��ϣR�1����w|pe<^�ک�݈u`���&�������{����H��O�2|u� p�V����3����\���lk�Û��8�R�}�ʙo����̫nh*��oD!������(Ͳ�r9E��6P��/��*��5���x+2��[.�R��@̲�\=�Qw*�}��lmQ�k�\EV8ه�^�ܫ��=�[��ՖA��;]��V�<���[�g*�;���yp3BVm��`<5TL]��K�����E4J�lvj	Qy�Z�����lP���]�������i���{I9ΰ����/4:<�b�k�"���5����Ȝ��^-]M-�Ө���n֩,���'�\m ���:�!6ׄDj��e�#�]�Oh:=u�meו=��ǣa����/r{4W0Y�X'ؚz�G�*l�\4`��Ȕ�y$L��"�$c�K&<����V/FEKGt�%ńY���UuN��,�J�1Wob� 8zތ�E���uWŧYԖM9Z�$C${����9�u�9�ʺj�$�ɩ��qP�W�N�)��d��\ėK����K;U+�oyfZ��V���l�%��;?{�Nv(�2x���yf�ҩJ6��^����z���X��$ٖ��d�lpd*�n���owT��2*\�\R��cfr����+R2	���@���ӧ��\�TR��ʴdS���[l�`�o�3�E�d,�v��i'"l�k�
�FC���x�A���z�R>�eߎ�<�~�g�EI�Բ;�E�fˣ�u��X�/�!���\U#3hwu�kV��%���Qk�*b�4�5�,���8���fP��ҫ�f�CH�w��W1x����w�EKZ�C�EPhk35���.��u�vr<߻ϯ�FNAotD��1�ge:#�Z���O��h̺�!xCW�X�N�������l1V ��)�C�R̨��piS���y: ^�q�2���Ҝ�(��57C��+kwy��xz���˺*���V�CEt
kӏ���ݫ[������kI��U�=na�]mlb�lD�-�+��������b��#[�g�}�ci
��<��.�F�ޓc��Ojl�w���'ʓ�7X�%Le����s�]!��Ь�F�)w�8�p1�f������rb�gU1��A!z�T��5Ք�:Z�u��Q�
{�*��)>Qŋ����	_OX{�J���`��*zV��J�P4L����)M.؝���/����Z�v��}4p����	���m��E���T�*l���F"��F6Չk�C�aOE'�T8,2V��E�c���E-�J�G��걥����58㏭[���=jX��[�=8ힵ��3�`ю{�(���Ϭ�VN7awV�� bw-�V���ؒJ:a]�u�1M{���Z%��%P�[O;�Y�y;<Q�5/t��[�D1lggk�Ӕo��B*S���dQ�n�Vm�V:�]�IW�ǴŔX��_P�QY盁��Q{���q?_�=�[a��<X��ع�oqd� �}GG/�8u�Rk�5>8���s�k7{=j"�4f�s���({��>
�7��C׵Ft٧��鄳=`a���>e�����bց����.�{�wo��c���^�J�qEǙک湺���H"��J�W8���/��K�T�tȊ�f�q�t����FH�����@���	"��@J���[��k;~�$-L���'6��wf��聈����(LYj,Ml�;��-�w��u������ V��f]��J�[�<>�bhrcS�N�c��x�^GO�Uْ�?�myQKw�U�t}��Sc ��/b��d(��y�}:�7���TG+��6���B^�����t��.�,��b
����nƤ��e�{���Գs]�Q������J�ht�v�'���v�齱��)�IȜ�e/9P�}^ϻ4�R.O�0�s�^V/p���e��k��
��n8:3�y��@�F0�5�j�0���]<������δ�;�T���J�I���;��.�����\F��M����0�Gg��sί�T;�r����.�q�!��Jе�{�A��;`���[[�OP�{r�0t�q�]-���z_�u��=�.��о)+���v��M��f����O`ҝ���֭N��P7unK����ѧ9��!�����k'S#B��KyN:��@A֖BnV�Bkz%c������ɟ����(�
	��ث�ue��5ٚ34�Gt}���~O�.������Юm���a���d�Boe�7�/->��Y��w}s��m�v!9��WW��xS�G[dT�����V��5����w����,j��J�o�sO`:YQ�ї.kvs�{2UV��u0k��Vk�t���BU����E��EHN��푌;h%�N/��*��M[��D�4}�)��>�m�:�@i���y7�ѽ�µd~�`�۫�~syC$��°9[���ϻ�QT2f+���}l%��':�]�%�rJ1����Sw����*�o��A�Q�4��$X��KXN�j�K�BwX���5�"�ƽ��ǂ�*�a˩q:9��f���6k��=�>A�e*<�ڮfpk���_��2�Uz�EJ E�B��9j{������BU�Vm��`	P�6�hB�q��7�;��Nᤉ�Pv�Y��w:!�"�)S�%��vE\@�g�G]l�]Z��rE2��J�w,��;:n���w�w�к߷�Dw�{L�菴�Xq���Gb�e���1G;&��d������f:����F*��!��D����\�f;���ǐ�ꙌЎ�%ܪH)�[�L��11ޖ>�W-}�7�i굘� }� n}�o��w_$��<���ě��WՈ�6���� t�Ot̬Ղ^�b��V��7�}�ҙx�
<�c���������7hR�+�m"���l[���۷;,@���4wR��5!ұ�s۲� �<�\��6��9F��)"�����'�KB��i�K/G��lB��'��f�ry���	�B�\D�,������T1>��I�@��q�S����hZ.m�m;��@�4R��4@�
Ȟ;`�jZ'}xhқ���(N<�Sa�x/k���w�Ʌ?��Ծ�ʂ�{�+�<�#��d"q�yO������D�pw��r�77Cv�s�!���*���4�R��+�\�\�����K��9A�y���-���-ѥ��t'��nM�W)���u>�ږ���1�D�;D�Kz�3��w}k/�.�F,�����Qi���	����Y<�c;�݇2��5��i3w�����wJ�����y�hƝ�"Y�z�/��E��'�*ǌ��@���`KA�n�����a֯z�����Q�[����9ZC���z*�T:�G��5�V��ᇎ�����u�d:L����?Z�ǜ���sk��n�5���#R#�1�u�2w'We�vR���j���F�ᙊ�X�-R�\5s�r-և������|1]��}�Է���� Z��#�u?	�����eڳE����3��^��+��2T���^�z>�1�����~=� 77���5��l��u7yr]
��9���a"{_��V�k4�ɗ�ëu�9".���ݧ�7>�\��Jf�a�R7 �
S��q��T=z���M���������"S���	ek�H}�И5�п�3[�r�&��)%F�̵��+�������M���=���Q�ȃ���cBr��ކE�h˕x���Y�$�H/��Q�d�n�(�OM#����_wd��7`ҭپ���Fc�����|uՍI+�]��멊s�xI���m-}Ox�f���M�,.B��)���	5�D�#p���B� ������֖X��{Δ��J=�۽��rj���#�-!�4�����=�eb�൒T��5�p)����+\Glb��͈ab�Ys����� �Y]����% u�{�7�(��`vZ�X�Fv�P8����S�Cp���k��������jکF�m�m�ke��DBڠ�D[lKPU��m-�%"���j�Z"��iiiK+)E
*YR�j�Km���-����j�(�F�[e4�Q���Ы�Z!ED��A*�mkm�Q��ҍ�m��6�F6����"���mkm�Ŷ
�A�ֵ�*Q�ԭ[b�+hڡhږҕ�)bQ*"Z�b�,��dUJ�b�-JVV�-����R�Q���-iB�UTZQkm�Z��F�F�ee�X�ƭ�eT���VĪ(Z�[U*Q��%�X���+ij6�b�(�Z�KKV��*6YkJ�[m�+X�EQ-
[Z�JZ��Ym(�mikj[F
�m�Q���QDK+Z�����[�=;IF�!�N��C���#f��a2�]�]+����;M-|*��.c�-os�Z<�`�^lR�-5Mq��b֔nդ�Ur��7�����包��|+�ۀo�0=����h(cj$ss�Nb��٧N��qLf67٨"�G-{��w�E��E�:0�F���V7�HN��7X����C������^�s��7�{����u\�p��+��cw��;�A�/�������&u�HθF����x��{���6�6k�Z�MIp�B�ج"pOX�_QAuJ������������3�qM[��=a3.8#+�DU�w�ت��j`�=[��߆����#_��c�!���)襰c��
��^:y{��y��V��o,�V6Bݡ�#�Z#%7:+le�S����)�	���U����첛�wJ�Ƚ�WS	vʆ��j!��*FWK��YQ�"D=�b�>�e�;O]�Pj�ei�q�����{ރ�OՔf�(,%�����Ѹ�E��\���a>}ė�H\9�����2�"����!Cdf�<�v�r�τ�Լ������<���4m'�Z������T���:��F��[�������p���Ts6T�y��YV�{"S��q��1J_'/ހ`�Hi����X=s�nv3��Mp�϶�u0Ȅ�4Dsr�����Y�-��LR�vz�������T��D�+�"��j,NqTCY ���R����X��]����8���z�t�t��v9�LcQ3��):cF
�������N�ك�����L�ʻyrތ�(-���K�֋{�[���=ȷ�:_a��V�\4�A~o[E�7Hf44b�u3y0�r�dr5n��bU^��׽{TV	�p��3BWu��U�C�"z �����i��=-���n7}=oz)X��Ve��������d ��D�OW�3�GL�}���峤~���=}8T���LT��Y���:9EXy��+���>�E�&چ��>��ѩ���Kͧ����ܣǭ�9RG6�­���� ����t�۳J���}e���Z��S�|r{�^�%�C�q���ǽ5Za����k����έ�Wx����e,x<U�s�j�ee�)�Іu*A�^X��_��:����V�-���^}%
7�G?mf�"|+���v��j���K}j�r�[ݝ8)��㔏}(%ї	����y�vu�[vu{VE���R�v]�P0�s����s���T��75�Z��U՞���gꦛ��N�����>�v\(�.�����@���dFv�q!�}��V�!\;����������x�ޞ�Zy �����W���wB�d�`�˭R7�T�iYc��+�9{�گu4D'��btRp(zP�2M�R�
wq�h�7�G�y�+��'y�=�f�����e����:����svR��G)���ps����Fޚ���GU���*eM����d�=o�@6��+*���d�t�m�eZ�����澉f��\��|�mQ�k��'�F�z^e���į��I�o4gob�Qg�[!|̃N�j!���=����#Q�V�Ĝ��U��B������R_�彃Ř�h�&֢�Zљ��pv��u���;I��û�����YY���ij�=�g����&;[�0E*K��_,��wU����j�s�r�OQPS��XϗS��r�����S��ɫ��2�v�z0l������(mo�8i>�|�׷�f�9<�b��3��3�q�}Խ8g5��DL�gRt�r~�+�[�m�*���������՛����;�ב���8,O[73H=7Ù�Zm��֕�O�ln�B+��%*�,�����av�C�U��(�PL�v���\R�:�F��+Xy
���l�Շ|w��h�n|���`G��v��@���Ry��,o*�8��m�aF,��憄@u��Y���@�z`��������ް�vwk�qZ�*�������m�<u�(��kbg:�9�Goo�;�Uk�*�_�8E��
*B�4$ɬ<�r��X΂���E^��0e#�t�mT�n��W��WF""��5�J���NL�yd�W���X@@��ʓ�ER!Ր˗˝���Ɓv7q*=�f�x�v���FZ9��gUvo@ׯ�s��z��a��V�^_�n�.�gTJG
��Ӿ�� �b���xZ<���l-����f�$�iaۍ5+WLR1�]3���飸�^��h�t��-�:�n�ᬝ��N.�m��c�G!bk���Uș����Vܝ��m�ju$gR��h}�*k����o1C�CQ�hs���\F�wB�a�	u�ۡ��sθa�5����VP��vW����7�03ķ�8��ex2��s�R���s���ws�4m1^�����9T|���v��ҵUs�yg>�
��i�U΀2őm
���F�'y�]�T�df+�T�C���)�;��ϐ!�]ee+���A��x�{�6�.d�yd1Mr+��/6(+�����#�1�
� �P���gm�N���/-p�v�ݭ^N$S�ޑ��8�׋ᚶMbq
��tguWo��YDu?mj�N��}i�}��to��}n�P�W���Ϸ^!�(Zs�x.R!t�N��f�+�{Γ��,���#s��8/��tmŨ5�O��)]��Q)���
_]��iT�%֭b��>ޣ����լ欋��	n���P��\�u�*VT���q��r�;G~k�~�S�c�"+�=�p+5�>ɲI�P�]�>�ו�.�Ɵ��� k�8��-��aOE-��&2M�����4��_	���^�8�v��#��Z�fb�A�쎨Z,7o0>��F_� >��p�$����n��*˟r���%D�sa����7m1{o���4����n"a�j���7��Es0��j9�����{�Fy��%8
aw8�r�SG�pj.a��b���%�/F6V�{�D'������.蓺��-�AR�;Y){��/s�7S%\˶]gSѢUpr7�EKZ�\��ܮ�ӱ�W��)��ޫ�Y�o
�F��@��͎LcQ3z�d�`\$�ٚ1��+��	R�o�}��+2�v��6@�B�����WS��N�-�U�د�]X��}Z��U����R�n0�w�]!���b㡸K�����P��8��]&�1�dtZ6l��{J��攬VZ��5�W��l�������e*���&C�F��O��a8\���&]ۂ^%�s.�}�Һs#7h:֋���N��\[�}�1����YO���	2wU­j��s1���u�m���&�n��O��f����@����PKq��m���(V!/��E���Cw��ފV.�f^������|���v�[R��W/��ћ\}Ǹ��Y˶w���q�����/�Lz�1�t�rj�]�&Λ�^<k�SЛj�-c�C��R���zۖ�7%W�Ӽ�f�<�b��4��ki��hbq��Quq����hs�Sf�P��Yӏ�*({�c����P@u�]�d��.�n1o�IO[Vm��Z��2|�A�װZ��D���Diz.]�[ޖ��=]��DO*�a�j���U��Jp����л=��o��鳓�'�C3��v�7t��S���pi�K�9®p7�,�;&={�ӥ5&�0{�s�L��l��h'c<��&��}�kn�Z��r�:c�*� �ڛ���y},N���xoY���.٤��몡�{���b��'8�<��j�����Ŷ�09�ɓf.�[�ܭ0t�p�F9��������(��� ���mu)��A�ڗM�7P�w�\�vN8%[��c|;��T�-	�LK/��-�;� �{u�]c���7�*�lIr��}�6�> �ѻ��=�NS{g�9�s;t�k����O��؟�6��ɡ�"�s�fgwVe]�m��!Vq��V��v��7��N�Xb��vҢ��#��k�z6n^e��^�YA�)���:x���6��� 2��Ε �r�WS��3�G��i���O3;�o���=����WϔSD�T������Y��Oyf�{����8x������$�:��	b;�-nN���:�R"<��+�蒱��O<�I>�	͌uf�5R\Y�gk*����,�tj;�$�ث��Í�wF�V������IE;��Zv�)�������9�l���7w)���;��P�j���B����9C�2��(��z�[�+�r��AxIY��i�Qr�>�gpŌ��c͍�m��@Xp��/M�K��	��K>	/�g��������-��E'�����sW��=�e�K���!|l�����Gf���U��LoXX�x�}�ɽ�*ҍU*�s��F�+Ҙ'�v��i��n��(��44-u�;m�ٛ�u<���n�Je�=���Z������е�H�Mν��r��	��r/^���Wy�V�"i��ݷ����*�XL���,��q�ǲ�M����ev��D�m�H�}�U<�zb
'D�Q�����s8�~�Y$Rp+҂���xv$U�}��8%�W��.x��z�o-P��]�xP��׃�"s��U��e�E#���B�~,"�5-�\ݓ�]��X�,W�9��91d5&��T8�v��1�k]h�>s���6o"�O�
0��)����GÙ�q�2K�5kSP�\o�{��w7���r%���kp�al��WS�-��!��]!k;R&{��>�u�n�Le�YTS0��hP���O6������3���Ԝ&�,a6���t�ǖ]�k�(��7�U�������fm?y[��ε��c9Z�T�~�ֻ���ŲY8��[P:U�x]�o�$5�[�y�g��.����㽷
����'P�i.2k�WV�ɡeD�7�"��ݩ���]uWٝB���>쫬�nv�hP��:��*�ؐ�#�,��ڵ�q}��ڼa.�>y�C�����=uamt���hq�z�mi^z<���{�F<Y�]�����ΰ��f�e�ܹ��.ud��VUk����)��(�\SX�C�aOE6Q����n�^�C�.b�]�,�<�_s��P��F������6�Z��[h�'���JկB�f/`'��ºtY�b��E���6Bݯr����ǝV�sR���R�b�����d���M��U�R��\�	�O������~NU�R7�5���YQ�;��{V-��+����}��N0{*�����G�Ղ��R�s<����	R���zүm:�i��5����,6��j��F�Z��w�k�z��/��aR�ﲎ׷0����ˢ�C��˼%JRoh0�g+`9hu�u�h[j�>hc�D���4u�&E��|�˃�XǏ�ݓj�P����a;ތ��2a���}]�S}��ι�w��[<.N�0�Q��d�hhn$x�2��`�m�9,3y�
�	�A���V�Y�B�ēCKs�n�kU4�ՠ�֦m����ώqR���M�̲��Uo����;�kx�Ց���������3 X�U:+�^me�2HԄ����s��ac�l����\PIEӽeJ�|�/�^�y�sW�]}�|�h�����1`�y���Gl"��nŤw׶⣉�X�n�V�eÂ���Cb-�=y��T9�ݭ�� l��/�����	 z��f��Oh���<��L����,m�1n�k0��f���zӘ�N���;
��j��M������<�!�Ѷ�����A�S*�p�|���A'��f��CV��]hN�b�u��a8���㒯����z���rb��\�A�Rd!_ƞY�¹�(�Z�)�x�0WsE�N�@̻�Zy�>&�]5���e�qڗ�8Ìc0�^�Eo׳�ɽ��۬V�����.r9k:��sxx�o��s��4F�k�c�օ�Pod�,�a%Ö�\�>��}�:�Ƽ�d��}[��>pk���u~���_jheծ�wu�k�l�'5�]�=r������ ���<��V�}޸�l��PF�3ه�<O^9��|�6Ѷb��;c��Rեc��;�{Mo-�9o�:l�����q��ף4��`:�Ŋy�\X�����d����mۚbv�	wB�P�88މ/�
S-�Uv���L�˽Ê�oj,6��l��VG-\ܿ�!�Bu%�.3^�@iVϻ8��b���c�yܹ�{j�A.ں"��U������(��IY8��u��S�:j9�T�K�^�Ȣ����zTc,)�x���[\NЦoJ�l=t�iuJ�����O����֜&�x[�x��NT�����,	�v�:\��G�@�e�۝-얨���ha���	5�ze�!��t��c�,!���`��ݡ��](5&C��j֎�u��%���g�;�5l�Pb��Ӟ���b�F�v�k�^L+Iʅ)AЪ�
�4H���'�9����mA�Q�P�*�e�G��Ɔ'��B��A��D�T�3oU.��Z%ʭé"������C�]Y�L�Տ�#�ٮ�Uȃ|���R�v����APh��|�+!� O?)g��[���rX�"��﷡QӉ�QV'���wckd�FVV;��A�4iȞD�o"ۓ�m��r�C�YҢcVp�Mb�	��R뺴����Г���6�n�4�{)R0�Ǥ\+	��bӫǫf&�,���{/iI/��	����N�(:�}M�������''��9)�����OB����^o-y���%�"�% ���P�V���R�m���V�*�[�j"�D���-����-��
��,��ذ�F�P��h5(��eQmKX�le)h��X�,hҍ����#J�*��ZRն��[U�-�DDiZ��B�*�+iU����hڬ����U���ڬE`T�T(�X�iJ[F��mb�B�V�J�eE�l��֍������4�Ա�-��U)b�6Z��m��,b�T��E*Z��V �T�YV���iF��m�F*��,������VТT�-�Z�[Q�؊4�("Ե����[
��(��֨%����F��і�QUjXQm,Kk)h�Bŵ���F��-�aU*F�U[mTm+UD�e(���PR�D��B�+T`�F�!�`�2n�UK�v��\m>]$u����NQ6:߽��U�Y��c_z���K8�u�;�����`�dޛh�c9���`��p�so�1�����b]{����*X��󉱯��xvf���̣	\�m�Ve�@�Tn��(p}������EZ��쒷v]9�{4b%��ׄ-�y�̫��鳒�Ylm���
���Tï��j�'>����#i�釺rr����hsv�Έ�Nlos��=b�]�Գpw�G��y�
�I�J9�Y��;:�$ð��#D�p�ѯ٨5M+w���OX{�C�Ŷ$�ں�����s�0��a�ҏ.�Rfd�2�.S�w�9��ɦ��}�:*�ir&I���'*��z�p���k��YM�r�;��IU�
L(����V�~����82��"}OkǇ5z_j�N4��×��hoa��c����[
����Ef{;|Knz���S�V^��[ń؅fz�XY�����k�Ņ'6դo�Ӯ��4�������\p�w&/�V�)Ӳ�*0��x{���"�^!�O3޸�2�p��ju�Oo".�m�k&⅜)��E�3��X��;�܊C�}6���>�r{�vx9|���O=�I��(;�ZU+�������D�D���dD3�s�F����ʽ3y��q��X|r��T
�ד��dQ�zĭͻ�xY�Zb[x�:Ů{�Mc����8��D�s�Ԉ�6M�m�N��5r:��82����������4�M'�"XJ{�+۬K��v��F�N��Ijh(�t��-��gy�����q���KF�rNu��bk�%Tk35�bn�5�YU�ށ�����7/K�׽��/�hMn���ɡ�"�ƽ;��Ve]��R�k�Db��<k�t)�R`�N�[N�O��9�ָ�Cy-�zpd���h����6G�l�֖���W�������X�Us3�l^�3�l΋x��U�;Z���fX�Tv��0�u��F��^h]{%fƊº�P��XF��_�]2�Nд�F������C�v0H�J&�����e��i�j���3�A[�|�R��#�s�۝(�tI��ȡ�|4l��-�vL��Mەn6�{_�uGG1{Z|Ǻ��p�wP�[�r�m���ݽ�r�=Q88��3���t�����y9�洩p�w�����{Vh͆�So7��q�䣰�����s"�{|9�����Έ�^�=0�bY�t+���b-_(ܜ֔;�*�U�����A1E��Si�7ԕD��{���-��.�������B��(���P4g$�\�]�կksl����s�#�>m�v!D�d����sk�pM�e���WP�������n�wk�qZ�# ���EK�eLlɳٲ�)����'�a����cgۺUk�V��9n��=�s����'vT�8�9C��7 Q|L6���^�ں87�[�bUtFۧ�.bVC��*�uXI��'�����"�#E[X���Z�T�L�r���'�ٞ�N�b��74F� ���H�8wu�X�O�g�#+Wr���G��#w�dU�hۮɯ�Wu��殺�����\�� e\�x�>���}]��w�^�Zz��YN�ÝyxA}�+ =���u�lE�>..wtB�o7�A ��l�c�WO9Z\BY)WNDx'�΃�91g�F	�s��q�fr��]���9}��I;����J�2�al�H�Drch����*'�ʑ��ccU�,Nv�I�K���F�
���t��-��/Ns/m@�縘�(�wc�o���u99��(Y��o�b�[�s�f���8@u���'*�;5�~����YH��x�Z�a�t8��޸)�&�,[{�v,��s͍V/O���/�_��\����sWL�o2i��F����0���]����}N;O�P���h�Y��|��5�s���ev�g}�qMc�}��)���]�����^=}����8���*��v|�=�������;m�1�tÙ�=�)�8��_����*[��6�>�>k�6BݮY��ԫ]�X�VY]9Vtēt&��Y���(��j����Vw(�k���L�,"_��^��	�<��.���� Zw&�Gyu݆��g���T�]�G�`I�˹�,6�Q�twy��ϥ�fR;e֧�cȑf��	�u�
���N�d��7�L��~�fJni�K j���MUz78�-�t��� BW¶�\�3e!����d*S�'dP+F�!���ݵ�to�ׯpI�:�]1ڙ⇄�bu`���"��^U
���BإC"�&mZ���+2�=dhگXi��U��0�Ոi��1���yJ�f:�df�5U��x��9�p��KF�u����b�Q�_��q�;n=z��֦�f�F�c����YY�k�F�� }��c�<��Y\Z�4�Q�-c8�7/TEW����)�%^�鳒�e�*����m;�{e�4�ģk�J�kv��s����6���n�.�o���ʫ�y�B2H5t�/G*UHV)vȾR��ڧ��;<�&���Fi���%,�>��u�\������Kkgg{�z(+A�V�D�)"E6�e�QcW�`~c��A���C^��&�hO''��#�'����b$����4�����6c�N��a+�\vd�����A�]ݾH��p���	tV9�����F�����Kt�����n[�
i����Ks6+�R�f�s�?�贆'�V����W�ɒe��gH&��yl����l-��;�w���X'b���f��؂�T�&ڱ-c�9�
����V�:�,�J��r��o�v�)��w�q��w�p�'1b�����l&-;N�Q���:���E�ej�Z��j)�"Vu�`ry���)���yq;��2�BsO`+CB��o��̪4���/d����Z~���u���7�(�FBn^@idW<�M���+|��5�K���v������Y�^�o����y �J-i�hR����(�;��Xނ���t.Nq���D`t�g���3r4�n�.�x�T3��]g@�ᬺ;�(d�u��`t�C{�U]�D�ȥ��F�u��b1�)E��l�Q�"p��ʶ�ҫ%���Ix :~�o���&@�V�ETY,_غ|Ύ�lu��U(��ټS���x���0�5�]C�&���pIWqh5w�{bgD��x��. ��rs�-f���t�ٰ�(&�Jf�iyK]%��c����8)ӏ#��"����#�7zf����o149��ŉ�qC�k"gwVe�n8��T���3l��V1���
�K9��U���mQ�sZ�*�ѳR�m��̺�vm�k�Q�O�K+K�ߙ�G,d.���;ڮfsυ�!=q���f�y�k���.qeՊʠy��#3PG��ob��׳Y�:o���%����HQ��b�Z#�8D�9S���;@�;{��T���N�ۆ����I�1V�ݽ��M��>��qF2�z���7���d�w���o�[�Yؔv���P�.�C�XD�;Ol�~�݅�$��N����}B��Q��q���ջ{e_��PN>��lȝ����<vm_4�K�X�l�V	z�wN8���[u/������Jv��fͣ��)����eH�_�8W�j6^�;�ߎ��#�Z���\L�`��(�Ѩ@թ!���1G�����"�G�˩�{�OD"���Ά��w��wD�_"k&4	�;���2��M
�n�@�u9�j�ѝ�}��`��u��v蜱��xm��N��7Vն8|pY�3
c��V��;��
�D:q��[������?t��J�M2c���wJ����}|[�X�tm_f���'��;�dT��p�� n)�"a�82�c����W8O �&���U�Asi��:��H>��P����C'�T�nu�t�N��q��^��KkgR���9�Ƞ��`o�𙘐�׺tL{�w3�d��y��cy�B�-��9�"������Mc����OKp���#��V����t���.�ܘ�#�3jݿR��sʾ�C=:�*]�Sw�Ặ������-���u�C#n'���n}�� s���̸��6���BV�Պʢ�t�hf����FX��D��Q�����ϓ}����ެkҰ�Mo�,b{����M#z�4�^�|whJ��X�p7}=oz)X�)��/���=}%q;th�+�=M�c��f9��9�J��鮸%��_����urO�V��yR�+�����#�-9C�cI��i����qv漀�z`T�3�RޭP��op�����"���cQ>f͸����P$w�<�]'f�o'a|���	)l��f-����P�*������7�!��c�mo�h�q
�b�֊�g!���ݩθf�m�sw��.��{/�`��Z�bm+
z+3�V�"WE弽��9���݀�D�7��O�F��7ߗ�p�\���N�OT���ܸ-��9��Up��V(�wKWx�n�]Ԍ^��OZ�Ee�8[��ѾFPnu�K j2�dJ�ڏ��o�dQ�XG���@�J"x�L��uϭ�7�:�;�� 6~�ѳ�}9�{^jy��[Nr����R�:��Y�u�E�z��z�W�0�b�����P�q{�DnZ�Vt��)'NiJ ��K2�g����q贌"��@�Й�L�EK���cD�w��o՜JѺ��p�������)k��]���Mؕ��[c�Ɉzz��en�:�a�*��4�B�<�Ed:���|g!�}�C-�µ��ٞ�S�^�ns��<�ت%XÙ�c�d:Wys��5�'�=�{8˃�4���J�ݷ��x����<-	������r��D��k�w{��s���=ʼ���ƒ�S�a�ǭ�	m'W�ˈ�W�Q�{^�Wi+d˗��ڪ�����q�fV�q/�p=�6��"�<f�Pm�!�t������4Y�}�y������29�!��\���>L��{�������u3�Ϳ<�NK��)����n�!��L�0��<�]C�~�>�
!�r�8]L�N�^ȣ��O������>ٶ��cK��p[�ZmGG�w��t}���쯇ӑ���N� ��������>��9�(vE=՛���s�Gte��1�`�:��w�o{.�Y�⋼�f̗�.	�à7]����{��px;#׷.�y���Q�l4(���ϫ������39��l�T�b���s����oC�b���0��ܸ���Ϲ�����ՃA븃l���R�� ����|q������p�����Q���C	ҋs��ڗ�f:%lqY1 "%G��X��jDh�)��^�ֺ�P����NA��{u���T�"�XT⟝��hi�R���6r9kͅ�:u-�s(���aNB���LwK���;��s��͌H�P�&}1C�C�_}��Э��y㌘��ڒ����{ ���Q˒чq��a&�'��4-�9�G%.�h�ce�)��(�/�;qPŗ���=B��d��v���`�p*j�Epp!�ڸ�=<r�Q���{"�Н�׵ʵ�L�x�ʗx�j=;2�]�8��Q���9���U<t{o/A�7�G][n�p����ƀ����O		��|V<����D뭑ovfTo��j��4PV:?O�Q�I힔�Q�Pԩ�#:d�^����M�=S�&]��rZ[��o3R��y(�ӳҺ���=@
�|����P<_�_/�z;�}ÉrhGQ��H���o�&w�Kw1��i�L�*���^�<l�Q���sM�/nr�e����&�}tN|Mc)L%��=gz��.������ �زEޑo�&��)~@���Q�w_�y¹�l
���g;ݷ����x�#ou�{6�1�ac��5'#I����=�iפ�;�r�$�����i3Y�pK9���ُ {�u�f�AL������a=�򘆒4�����KV�5�)p�\��eE�`�y��԰{gМF3�-��95&�8(B$ܟF��]�$�D�� hY�y	�mZ]7%x9�d^�����z������Vz�B#g�z��wˡ$��YA����j�~�x��QѦ���^t��w�h�q
UsNa�4[�yh\v����R�Ԍ�[�#����69�+��;��7VXv�k\�HnQ3䕗��äTX��Ze]$��oM8㝸�:��\��.�E	x����WF��.��g\4��H��׭�c'gm#��^��X�נŠ�_^�q�$�i��z� $�;��iNTw�-���^(�떈њ��$/J�[%8�u�	N���-�^��lA�oY����1��N��ȜHȪ�e� f�D��R�T�{�r{ �$��H�=:�MH`i�����zOo)j���l]�j4������A��FWaމ�N�/.9Vm�僩H'�����|�h���خ�2&8��nG�� ��縺)�2��m��\y�,@c�#���@^k��fu���I��S-�sǻ���'����_&1��o�!�Dq�6�+[�(a��[(��N���V"����+�̧qj�Uh��t�q��rw��[�04�Cݢ�G��$K�m����~�����	�F7sUJ��WL����n��T��2�k/�u�m"�f�/T9{ǺU�!�|�^>Æ��`�[+P�=D�w5�Y��k��o�ˊ��K0�)(G�����f{�Ͼ�����o��4�i�J�ݤtYh7l=��Nw�Q�f���ٔ"�M��ܢis�͇s0��$ő���������E9������5QG�Ң�|f<��*��tx�J�3)��yvB��0��w�e��*�r��U�!�T5wZ�rN#lB�Y2������2��_�$"AD�PI%����m�����"�������[#DT��R�
ĵe-E�V�*J�V�V�-���m�ڨ��[Z���UeeD-iJҪX��J��JZ��R�RTZ��Q�U�k[l��UV��V��ZQZ1�V[k�J����-�J�Kih��F�kl-��"(�j��х-D��Q����$PD��ح��Kihڶ��0U���QH��h�����T�R���m`��QF���,J�[aR��ʵV��VZ�l��mh�V��F�(���"�lPQ��m�����TmZ�Z1b"�h�-���Q��6��jYJ�X�lZ�U���ږ���P����������+h�+U*UD[D�U+)PD�Q��TJV�6�"6�QAkkJʕ���TUV��mhQ���|�'�D�wn�t��f�J����Q9Î�]@���M�i�om�:Jj�M5�JQ���֞d���G�}RvMM��T5���W����IKR�Gҩǌ-���c���V��i����0A�O&�aݙ�#�{z7R)>��#��x��3�6�8�� 6��a6������>�կL+�cڳ��]��閎�n�Nw\ ��8*lN$@�T=j�4�L�
br���G�}�\/$�,9=s;�W#U���s��(z�3�X	留s/�N�rf�p�?�i
c9��k"T�
����������Y��f�C��>��h��!�^�/uX]����3�`�OE�����k��9A�d�,^�P}N�S�$�"�E8�V��q�y4��HJ�_w&ƶ�*�d\d�Øz62�#{�F=^�0��S���S����/f��u$]̭�8�V�m��]T���|1�o.a�bO�N��_\|V?y7�|��#{U�q�pδn��	�L�w�E�l�]�}���Af�\U-�������w ���L��A�z�m��fc1D��WD%s}�r����$��Y����3HgsQ|}�P:F��I�G���WJSޭ>9�����I�=i��+h��}��d����O%en��}���L�^1*����:׵{U��K�1U-f蕋�h���z�y�]4�f�>V0{������}�y\�٦u�Ų�J�K%�1��_{�<�r�@��zB��S2R����6���v���/F)Ъ�D���D��
.(vPV��Dt�X�]dG���N�Pn�ڇS�\�W��T���,:�K��N�K��"�B(]��S몑����9S�]�:� �\�w][��4BS}.=�X�nY�|"�&8ɜ�A�)^t:�B��tWw�ODm�i�,<h�b�a�/P�� ��C��ԅa�H�ڎ�������!��5�Bヰ��@���T砪X�ǐܘ��ø���xS�&�9�}��B�K�!QA8��i�Ӫs�#i�?�>y�V��.ު��q����Uݒ�a1|�����j\\�pE��4j1���s'��VVdg��K8�0�\3�RT��3_���5ן!d{�f��;ʁ߷��.}�� ��� ���t��+y9�z�AY�(z*/� �ӹ{f !�!͍�
�T�dߡ@ȉ���d����ik�ݤ�(�(�a�&�b�	�E�r,c��߶�g`W����Qmd��c��]H`滇��{*�}����ʡ��u��\@�.�>�}�܃w���vȳ��^F�0�Тum��et:���W��.������e���h,�K>���q�w&.5��11*/�
Շr	aN�4 9P���!B��_T�[=�)>Ma���"&��Oi�������>l^	�G��[l���Jo�Yc��;t��u��ݦ_	�q�E�X��_X��9J�e��
�A�7��4��=�F5�������6Z�F������{�����u_l㔭��A��c��%��t4؁�;HSVGQCw�^�P0ݍY+�{�����d1�QӰC�"�ec������|}�;	���ѽ4�gP��87���tev����<`HaK oj»Q�b�Ut
�N�*�Gӫa�͵�#���'��x6���1����9��Qq��(����*q$B��G�nH�u���t����vty�]�9/
��J��.zl�ezi���}X����k��#����^qw�s�s�+Պn�>��dS��@����+D����@�nl�RX&��1x3`���9� ���߲�L������R��F��#d+�xlآ����"��N���M��B�\����1�+X'!�G\��U��	�X�uN/�Y>8l���f,,n�.o��%~:�Q(V�۫%\%ż6�ˬ���v��b��i��J[�K�+rɥٝ8� ��1�*}������gmu	�x�2���W�W�Ր51L�g�|����·�m���wW"�+��3��!�3�y[2\�z����v��"ء�<�+?1f!�����զ��0�P���̵h:��a���p��O\	�
Bd��_��u��E�a��)�m3�;���D�u���j�P�%�v�r���ɢ��/���)V�K�Y/�t<�o��S˛e�3��Q��a�g
srP��Ǝ���O�i��y3D_�]��rZg�T2�<,�W�U3i�Is�8o�E?wG���G����ѓ<f�Pm�!�t����nLej�
�D��ұdl���H��2)��K������>�}/�Lny�x}2/�[����Rk%f�>>���U\���P�qBC�x+����l��(�7Cf2|C�F�l�.Qy2 ,J��|�j�jܒ�8'�݅��̔�N�
o�^P!-w�3Ϫ�k����rfX�Ǘ�}�J�<8�7��(�KPf�zY��iႽ�Ob�Yz�kf��g���=F4I����턜��J����և���ʹ��zRzes>[_c�F�3���8U1J��ѥ�AeןP�����ݽ��&���4��|w����c�F��%�+V��y�V���f�Д�lJ�ײp�ק�`����2P��=��1����ߜ�J;���6/�P^�S�D���3�0�eo��6{6���q�3FfE�%���Ӿ�y�<��R�fp��������������6Ϩ��-�)�G��G����rw�Z��P��H{ˌ�߼�1�XH�O���d�ǎ
J��3��O-g�Ny+ٚa2
x˰���Z�ъng"��ԥ"�S�"⏝`�G+��_c��|�����9pl�x!��:���缺���b���+����F⅄Ϧ0HۤwRǖ�]R�xEQ��N.K� {���ڶ8�W=���[d`��˾Ko�+s�4:|f�L��>�>c�����4�R�`�r���dRʈu/}��F��ѡl.���]pW��[�m ��
�R�F���ʽj�/捧3�8)���r�T�N����;n��jb�P{*"si^���D��^�x�2���̫�,�F:��ӽ׉�5Y��	����61�_*���� 9��Y�އ�l��E��x�=zK�ǽh�b��ى�� $���v5���֧��؏??��l8����n?K%^EޯpwT�1߱��8:�����r���0�x�8��iB�Y�7[r�4��9Q��nLl�cz*���m	�a]�aG�;��<��������=�	ޜJ�ny,�a�P5��n��OtZ���O���隞s��R�?K�p��J� u�)��Q���+س��,�lX�ݎ��cՒa<�!�T�nsd^�Fu�Ƽ�]iս��!F��݋����%�xj\�2�4и��~�&f�9U}���[��M�zƧ�5z�r��U�E��I���=�0��W��g�5���2�C�0af�&�^�d�+��٦�f���������V�QJ�.F�Rg��|F�r�'b����W�u���B��O��2y�D[��82��b�
�tO6TO<B����Y��]sF�� �暛׏��F��,G@�gG���Hux�eL�����qإ�O����./76&��B�-ә�:�FU�`�B� �&�6^�;���@��K�q��&��sN�K�ٜ�uQ�N��-^�GՄ?�١���i8W������.��Þ^�xr���3Vd[����}��7��	��2�	|�:^���B�ڧ=Q�8�q����C�V����;���UhF'�Bc��4,d�1�4���pC>Zdr�V"6��A�SpK|~g*��� G��=�ww	ަ�Q�j��3�X�f/r�y��&���.����Լۚq��nm�9T�j+�����;�kA�9l��ӛuiև��g�'lt�ܾ&7�q����1�4j����_.�f:�VfE�n�"�O��o�(����	R�ٯNzz�,�m3���˙<g����捦i����{�ә4��U��4m�1R��;����yX0o��\��`ϋ8|p��y�t3������_��p��̭��+�~�&"G�'��8�?ChqJ>7i���)%خ�hT֬�����>��f����],пT�+����?i'����6q�v��Z×�������^`�����������Y��}�7;�P�a��6��r�ʋ��3(���^�qFѼ��92Љ#`w7��4W�yY�':��;�.25�m��U(VJ��9���v�����cN\½���t4�GN��:�(eIw�;Ѭo�l<��>�V�0��d8�|�jA������]�}~��ܽ����;�k|��l�.�@uԓ�����6Y�����:�8r��6
�Wj<D,u�sҫ�WXN�*`i�@��F�'�·��'y>��ш576�	�;�P}s�}�zv�#��#V }�wF�\���YZ<ʩ*��K6��dK�5N������b�\�F9|C���Gpcx�n�\�-2�.��9No���u��D���t�jy���!ԋ|����xb�K8���e�{Hl��gj��X�<��<."�fN5����<u�rkGZ�lqM�܄��%�5����>\��4��0W���4�ߵnsӺf�:�t�$�7�	о�Z�f޶~�Y�S���t
`PD6V*#f`�����!E���r�E5՟w "y{������@M�cԙ��)��Y�_\C�~�1W�Q���;r��(���ŊWs���zu���]VC���[�p��rb�VTRqQ4FG�PeYx�VDc��-�VR���Ty�!X1��1f!�5o���NΈ�t6$P�b5C>xlnE�s|�~����������,����8��؉�PjC� �=��M2l�o��e��|��w���O����͹hu�ɢ����[��~��5���^D����f������5Oz����*�h�k||���&�yX��u]/���3�!�,\ӽ�4U���Zf��2u��Q.�����ѓ���M���	��H5���<�W���M;��n�}�f�Z| ݖz����{���p���O���f?l��u�Ɵ�v�xދ���}����[����#�����g�"�Ux�z� 4nrg�Vb�l*.��Jv��ɜBH���Πv��:���r��:�߽L��⪄�˳q�碰[�Ԃݛ�F"��4m�謺樳���bb�k�q� �(�y_�.�o'a��!Ḓٌ�G'�u���u�~�$�Jz@H�B��eK�*�ԏW��}\%瑬�~�u�1��q}Q4�/}�2��=T*q�7��T��6�M2�&�����@*+`��|z:,�,p��oy����:Ā�oW����j���8
"�)=5��m�6��t�0��ٺ�{���� �V�:2��OD�n��W�@G������d���4��O�s�35�q�|��L)�#\�m�s! �(�.]eKS1�+c�N� ��ᓽ[�o7{\��thc��~�G�TS�|�&v-:�^�]�O>`��{��e��ׯ��s{ͧ\'|�.!��u��C-�Rc�\/�yS�����H�P���Q9{E�#!,z7�B�����
�>�Ių��
���.3�a_���zv��}O/�����K0��I���#A�}i�_N艝�>c����ri�P`��nn=�H�f\�ۼ�݌���S�����,�ڴ6��(��kr�z�o��a�m�U�W��"���X�Y�Mu3㤏!����y��Ї���qFK��n�SJ����ؽ�f�N��bn����T7Ax�T���1h�՜ˑ>��G�<�0#¤�}�	��;���h�'�chp�=ޖ���	��GZ��h�s=�%��M��gs�Y���rBL##z��b$;D�i`'��x��a񯛙W�Y���B+���P{3�j�q\�]�6'�V��~�އ`��H��x�=g��د�ȓ���l�h~��Nc��cج��PB(d�,_q�P@��^!>1�O2.�s�H���m*m����n�Pdx�N��c����k=���h���S���*w�4�*e�\Dm�p��7��3�*ئ�h�2���$���$��'�4е����L����G{���TS_�U�u�q_��k�8���ձ5�W��q�q�3`�Y��t�sJ�%��-�!Y�R��p�QeEʠ�vU�=��)���BFn|D�#�]M�aS����7~|<v�~��{>Θr��/�
������:�����ګ5�|��^����g}�DF�w�Y\���_ڨ���1]5!�?}�]�s�?o��z��$��B�� $�	'���$��IO���$��IO��$ I?�B���IO�@�$����$��IN��$�	!I���$��IO���$��IO���$��IO�H@�z��$���
�2�˚M��������9�>�;��T�P�WFA�����-��EQ	J�D�����lŲ�[�**�l5�)R6�aKV�R����%T�,��H��4ԛef�e���Zԍ�K56��듭��j�M-����5[k2X�ĴcX���e�k)-,�4dm���i���kY�*�2F����mwn�6�1Oq�3fX�j�m�-l2��`��J���!������a�[,�m[&�մ1�X���Ֆi��m��ƥ�jj��a%fͳkjee�5�6��F���CCfٓx  9��|@�h�>������=۽^źsWu�ac��H����{y���w�����M=���'���s%�\�������i��흍�ӽޭ�ҡ컶E^�Jj%�2�hb���G�  v�;��gGk����y�v�m)�]�a������ҧEVT��[�+�N�v<;�z{y��P�{vx�v�=t�yu��Mz�	�����kwk���)�����J��J�5�k0�,&؛|  ���X�Z{���m��۰���ly����m�Z�����Wm�V��f�6�w��OKڃ��}^�QEy�a�@wO7E(
(�]�P 
( ��Ս�5TŠ�j;[%mY�G�  ϸ�    ��z(���8q���ޗ����wi	�wx��`�N���=ꨡ[Nx�^Δ���ګ-������x�r:��ݦ�mmV��i��k-��6-�  w<|@�N�cEt��=�zuT���:��E�u6�lޯU�P]�]{����n�{��=���]�L���Cޱ�����շvu����m1��[�   �����Zm�z��͘�{ױ�]����
���{��� �{׆��û3j�qX�{���[m��յ�][�������wkn���M��Zֶ�6�[fֆM>   <�m����w������C���{��;]]Ý��릮Ʃ�;]ݻ���ҩ;��yuզ���^��Z�w-�v7^�-�on�����ܭn�W����zVZY�=�孥J-j�dP6�  o>�kEm�V�g/Uz���gU�sx)�h�v7w��wl:�w��w�kn�w,ѽF��T��7s��ݺ�׭r��MZ]�3���^����g��c6kC�wzV���ًհY�[[l���  ��}zmuGz�]�޸k[�x�oS�K�{E�O7����ۮ����@��^��z=���zײQ�e����W��ۛ޳�z�^�u������̎�rӬu�[cZ�+[`�,X���  3;�F�С{�9�ow@�T��s{I歭s���wV����=����i��=WZm����˝[���k��*���g�p��4y���=e:��O 2�����~CR�� �� �6d�R��j���"��	J��#@T���j��@ I��*STi�4x���?�������t������?��MY;��sj}����g���|��$��/���$�B!!��$ I?���$��ID$ ���y�x�ϧ<�����4R��V��t��wq@KN-���#�i\�(Al�Uk��J��B�s%1����a��Ð�ܩ��-�[�ن�7}yD�9Q�a�@]Ez�"�F�lԊ6få��I��B�˓P@!��e�,2�ѫ����QT�+	ɴ�2G���-�*@3M;0LiebP�tVȠ���B�^��[v�P� ����5Y�圏lY�D���י �� I8E�j2�Xr�ۀ�@�����5S��]�"C�Z>B�7ta֩+iE�e��Y��V��h�oZ�I�pQ�c���*6ֲn���u�r��`-�e$�wF;��Xm����.��C;B�B��3[#Y���8��&���t��p9�+I�j�ۨ�U�%�u�&P%P��nö�r=��&���=u��f��A����,��r$�A�n6�	��;W�`z�W �������QҠ��ԍ�T؝�:�u�VR�{cU
�0Ec�u2�['!�tQq(�eicr�z5ϐ�hU<��0j�*�$2����_l�KS�oj��9�!E	B�\���LJH�Ce#YLV
)��tƳ3۸vw.}��sD�1�2�P��c%]���i92�W��&�-iɤ,�+RY��CB�^�7��ɸ)kx,M0,Kj2�jOu�Ǫ��;$e����W�lxug��gX"#6*��	!�i�y4�A�q�e6�h���'GJ;WIh1�kI"�"i�z
�/c5��^���SP�u����2	����f+�7�ճ�z�D%&��W@�Z�˽nm�3NK��أ@���S#B��q���O�����2R<�����9|�WQ�)�cUh�.�sn�ݝϮV1���qZv�f�ƳRf3�'n��A�f�F�l����&�7eZ.��M�����6Eŷ�LR�4	��TF�,+����ni�6���f�djV9{%�,Y���]�3q�X�
��rX*����R��=�%^(�8FQJy m�p���VQ85�Q"�)�m-�5P�3v)Y(��K٤!JćUf��� h��$Y�t�h+��3�Ė��j��յ���hyE[�
�Ij9��VL4P��2�&��ܛ�,f0q���k��wWi�<�,
D�k4M�xl��r�B��L�E�r�")���Y,��3rTX(]��Qw��^V;�E�-ݡ.]1���C��|2��R�0�_m�c��
aU�:e� ���`f���ی�3x0ϟ�O��̘������B�{�E��d�l�[t�Z�(�b��PSj�JH�^��Q�7��'�5�z��}���p�^DFW���K�Ʋ�n��tqJ�Sq����P��JT���F�ŗhP�fY�2���'��B��ʸp�����=�6��a9@M�7Y��"���*?Hs������=���O�x�E�Պ���Z�a��]ܧ�j�m���SkB��z�!��1c�L��#lsV���"��e,�AC.�eATV�ȫҫt�3!������(��[o!1���е[�Q�C�{��g6��)m�8L��6�Ƙ�r�/U&�Ш�	���lh�֥�hzqք�Ѻ�f�8>nn�*�W���a����/rݕ!
`!���՗f޷�di5HM��M�tbl�BfY92^-���&@Cv�ѷ��<$����x�+b��a1;"�TS+6��S���FJ
�7[�L�f�t)���@3V^Q'��S)�R�c�$���`�
�XTւ�#2Q�j�)�J�6D�W��A�5o�L��\�&�0P�w2H�0V0��OW7iR�D[0R�� �,E>�6��A�b��^V�ŁPO!���詨Ru"��(u���wP���mŢ�nm��S�[v]�ۦnYi�q��V*m;�d7��;�ltP��0V�1�jM��zhF�"���77@Ռ������$�@����P��������h慃@��-0 6鶉o*]
9IJjݤ�2�kR;�Ap4݋c*�������hAɭ�9��o�Qe^���&Tӑ'@�)fJ-bL�xn�Kq��-��\92��wr8��pjR��Yvr�L�pm=e��O]:s&5|0�ɋQ��8fJ�b�aʂ��k�T����Ǹ sWro�q���c�·�kx�9��ۥ$0�@E�Xѡ�G6�����=F�r�n�Յ�C�Z�@��! J��r�ӳ��M��`�\(�)���
���ڹ*�;U���O	T�˂���Q�`a�����ޥWs7��,�F�-zb���n0�eh	�iJ�-n�˖��@�?ko���'Wf�d�d*akL��+n�Nt 9����0�:
�{[N�.ӪZܽԝ���ʨn\`G���:l�E��	W{�[N�
���O�����͡x���9��b���/wH;e�D���+%q;��r׹p4n�x-b��g���B
�*-�1GKf�5e�w&��4�N�V�[OlmhK��{����gy�Eq����!ǈ��.����(a��Pj�m��0�K���ƣ;7t�hC�ƻ?���+��k^T��qы+d��.Ȉ�u�SÂ�#뺳M�����hf頍�ա��JZ�p��ukV0sv����X�cر-{��M-ɒ�a�Ҍ"[CkpAuq�h�[#�#Z�Fng�Y6�Z�1f�6nڸfk���ɶ��D���fܺI l������bc��0�ち����98˺}�[b��5˟((&�`�%HoГ��z���}�yr]�p�kHz5�
��x���6��gZ����|����Z&͉-�U[bl:�h��Y*bQ�ʗ� �l���c0J�Z�i�%�Y�6+%����:ͪ�� �2�����׸������9�wE[sq'r�� �,�2*�3*񸮳\����oHi�X"�
��A�;!��{B�n�mϦ6�l߼���a��xS*p>K���qav��kF�bޙu&]�Ժ61�Q]0���lP���cE�]��$̗p���K���s>X�=R���	�f�٧�i
���aŝ��]�1�$��j?<Ƃ������x��]6��x����zE���L�b��$�,�W	!��.3��!�'[t���Y��	n��rf� ���t�Fi%f���1Xd��t�4x��%y���uϓ�kz�֎�n��oޗ�k�T���T�1�z�ɫ74�.=AJ<�pR���ޔͪ�YLތ��ƔWs�i�X�V�B��ռ7*ڡ�w��{.�Y`e���%����ҽ��b��o��B�������{�B���*�XoL�|X�Z<y�ʌ�s	�qȾ-]�RT�f��㥹��]!D�0���#a�5I�+m�P��U��ͣ�mZGޅo�*TH(���0-0iK7Z�SJZ��������)-���@4D�Ңqj1�3/)mI���ƈz�1��fКV��ʆ��ɪ��	�ӳ6x�B3$Mc�#6E;��uMT%��r�ٷE�.�u3CDݚ�Gz�i�h�ЬA[������ÈJ�bv�#8jÆ��n�d
���t��BP6tmM4 ���໸mel�YA��������"���9zl��)eh�P��>��?���a�,���̠1-���J��7�R���d��VP%���BMP�5�@�y��j%�IC��n� ��w��R�mCyY4=:`Vd�̚�H��
.�ZNJ
�����M86�A��E�\��K�*���]�s���]�n�F'�Z�g)�5��q�����KS[�XN���y*�[���׫r��� 	0�S6Ք�z�j�X��5��#"�=�&���>%���Q�ke����	L^��#����dvrm��,sMK��14LۻhD����g�(Mh��yiB�&�Ѡ8�X	���/E.С�lj}���˺Z�H�ka�2����\"��U�b�e���Ȅ/BuÓc�j���&�e�U<ײ���Ǆ��������Ze��17*�͵���EC2� 9iVֆc��n�
Cx핔��{fQ�I�����7�)��+.��eb��q�z����*���P����yP�ּ4��Lk��Q�t�Z�E[2<�lV�)2�cfқv��if	�-ä�5�ޥ�K���L3�X����*ҜAr�أl�(��Xp���XI�+�*2�9HD���.�7uBD�
�0�lQX���"�
��U����*7�X����5Zm�E�T�ъ�d��g�`�rTx��%3(Kڻ�YqT�v��n&s��i�d����Զ�
{��;t�fe9w�6�͌�5d6MFjh��C�_���aL&N����N���S
?�b�i %�4t����LM��-T��~r�T��+;-2l�
۫���U���q��4k�ĸΌ
V�IM9N�PJ�l�ć�o{Ќ�&���]S�hYy{AP����U��n��yB�L�1���U�F�5�2�BֲZؖ^�"�mY��[ŵHcVs
�1e��Ѕ֡%���&Q[�v��vCEn�̃p���%�����u=�F�%�&�?4f"�ű��g,E��:��_E)�b�K�� ��S{1�
��1�L���b�[yQv���w��J0L�'gZܻl�A�6��%��N,���9'�0�%�V��d��H�+.�:^�N5X���4�B����Y[W6j�*a?�6F�e�*����R"�͛Q��D�i�О]��1�:YQmC"-*�Zm^:���wZBD�߃���
���VV6nc$J��׎+��0��؉ikx�!�
�^�<x(�;����6�w�" 	oSJ�;"!�%��X�����;�f��2d��^�@���)&�Ɏ]%MEt�T�㿎�ͱ��C� =	�QĬ�1�(@�3"@��P��[n���Zء+r����Y��ޛ���n��� ��W�.�/`t�Z���u=�C�Sm�TŰ3X׌RG*L���@���nfb��	E�v���Eݘ��Ei�n�Eiu���f�۹i�������S��^D��qNM9�E�H��O��e�Q֫{�N[5%��.����.[��0�lX�����m�Ƀ�z���l��)�T�/6�1֊�P�A
�ذ��ӊ��b0�;��lgM즅�/dٱ+�F���eX,����RE?���y�W���ͰK��F�óUl)��Hթ/R'EXݫ�G1k��-�G)6
���eXj=��г3+V���ˬvoT�Ԭ;�e+��)�[�w!�ܲsV�[��`����t���e^T����6���R�ޔq�i;�i#OopdHze��)
��Xnnш�k)ۈ��"�aTK&����
���X��Nm����0�lt����uu���F�Nm�
V��d:�Y�i7Q[S��g}Wb�Yp8n,�S&1��p�"��l���!��S�q���f�A�[�j�l����fͬ��P
WbX��ʆ�M���T�ޫ�"��,:�ʩ�-��cw0�qm\���H�{{�p����RI`Q�ĕ�0i;��s������i�r��My3q���ʎ#F=�YX0�R��d��x��ā*�Y�Z��h���nh51	�u���%O)�o~�-C��6��I:Ia�p����e�
ɻR��,xi�R�	l;Z@փtգ��]�.�tf��kUM��7Al4��18���LU��Pٙ&m� wB��[��nмQ�Z.ί���z2�E��M�*Pbe	nj����hCI�B͉�۽�pcф���1'7M�%!.�V՜��HO��܉Գ���fG4�ދ�&��$�=w�0�A�g�E��\�	x�c�9�`��&fOA��y�ѐ�<G����7�D�QZ�4bRS��:j={��HիL��SU�0�[a+Oi��¸����*{�5{t��{4��MnH*avag����iٺ*H.�Ǭ`uc5��SZr��N�w[L*�@�/K� 9.���wD��;H/���)M��;%���`�Gl���6h�r�^�V@��j�]Ō�P�m���Y�)d^��v�?�V�81ݩE9m��轁dF�۠$���l��9P����"���V&2��ŹM����n*��:9d�km*|�(P��R1��&ᕏr�D�l&��J��V���w�ܹz�F�e<�M(��30Iٞ��J5�I�2V��V��GT��6��0@(jztY�L�E��Qt��۔R�̷�RzZu�b�Hd<��u[�ٰ�[c�7n��Le�+*���{�	;A�Vm3��RiKі�z,=�Iw�nd��F'x14(\�e�W��刋Y�J*�r�t>5xؤ�Q�M
���݃��s�H!;���X��j�%k�0xK��_RS:m[Y���)ʲ�q/�U�c.���q��A��ݧ= +��(dTr$ʳ�4UCd�<˫��V�q9��X�UڠЫ����.�ڒ�.�K�JZB�e3S6]��i�6C48�� ����6:�D��&A�w+�ma�nI!����XǮM�Ȥ3ba��E���W�v���g#��4"�@s�ljh�ݪ9*8�b�l'+J�,��W���I�c��kN5AS�)شZwB�h�H&7w�0@5;�#�[ׂ��ё|d��mb����T27��0���uR���ґ�E�%*ƒ�/�*�F���a=�]Q��6����5s�+:ͻ}B!�vy�r~�D,1bn1��<�|�JÂbA�M\\��Q9V��ǚ��) �%�����]��-j�Z�o�^�Fwq��Y�n��VH�89�e8s4�<;�Z����yӼ/ST,�u��;}�.��=}��-G�c��C��#�����Wi3[r�ܵR�V��s��`��0�XB]��j�;}^��E����k�4e�#�I�g-�2ՖC�]e��Q����*1��*(�V_׭d�M�UF#o��}�q��o��{���	��!�謰�jR��a>W��{�rMi��� �����8.
P���E�.��1�.��y�V�Ss r/�x4��V�uu�Y��Wol��mL��ڹC�a6��k���k�t��G�^��)��Aa<�a��LRЬ#Ua;��Ǔ:�]� X�ۿ ����p��<}�2�l�x�ϰϑ�!B5ه�_&W:Ø��V.,��+^�f���Jbn��9bj�ڏ/�Wy;#�/iL�GL6-�E�,^��cܚʣɝ����z����s�8�LмL^s�a�U���ws���!L2��t������y&�z�GžWl	R#��┶<ث-�]�-���F-���%lKh���
9�����f,V�:�\�p�-�����ip���R�)n&ѓ
��ޢ��ow���\�F����!�/O
���Cn�ѽ&�w�/k��yߢ�~�E�{�)���wi3��ekD��	\��jx5m��6�R��Lq��%L;P��R]�æ���ѧФ�6��xxe(11M;�
o�x�������x�8�Yk�D��*�LM��*fwS+�2��q�]5�|z��G�B��R"X�k�S��X���U���	�CRl�{��ϵ�=�3-�!޸ꕁA�{�3q�)Z�"���X=O!�{u�j;ǹq£��R���%�g��1�ެ��]��d�� u���'��N��0�s���15S���{�Tcq��\�j������]��	�Yʴ��� f�e2�U|t�i�J��c9�ͺ�Q@���5*�.��̎)&��
��o_l�H�`�.ƞд��|��q�����6SV:}B�!�V���-�P�ѥu�ب�y+*��.�k�G6���t:B�k��qY��=���G����\-a�P��R����,쾜0�1K�26��t:E�j�H\$���1�VΠ;���ΥҐ�Ucp�YVÛ�z(�]���B&��oh�����,������ZÙПh�N5-͵��gQ�4qwnַ*�t�k�����v��O�u�q[i�ܡ���N��k���4Au7x�^\��
ҵ;Ih�zȁ��4+����Yf��*VfA����hה��ٝ�l0W]v�v����/d[7���Ff�,V�Y�*5��b�1��6�n�e#m�=�}�����z�cgp�(V��*�+�Q��X�m9�sCP��>������[�	�So�(l����"u��7Ϩ�\��L��`���,�}>4��Ʃ�L��N( ���{̳8�HK�O5P�H!�/2�q�vxI�8/���;���ڟr��22��k�'	�v��>�|��ȭo� +Jw�3yz�,�O#`�x�7��\��B#��{z�Wk]�v����vr�;(��\�JJ���5�5��؃|zZ�ѳ�@�&#��ro�Pd�{�A�;��Y�*��ܡ���F}��٩a�s����wF�֤W�:G��>.���G5MW!��ͭ��-�\͔�2�R;;�y��x����X1�O�Ju9�:�����]w�I�xv�����O#�hi�AĜ݉sO�yU(�`�o/E��O���9F�cög���:��}��Hr`N�3�دB��6%۫3������HyO\�ᦔ���htƮ�C��x�:uuw�p�v)%FY�蕓!⦑QTP�Jǈ����t�Ƕ5.P���gF7�W�(�˚�g���z�,=]f:��Ί�8%IX��-�Z�)��KǴݥ�vLq��v��s���|޾V
=k�kC�zۘ��kE�Z �6�	n�L_Sx�q(�Ѯ_4T�-�#͉�	:���.n^�'8��4�P�m	��
C�H[W؁J��]��{��|�n0�Z���
���i�^�	˫�N֏ �XY/M�R�&�x�$R��*%*�P��1�qo\�8�)�A���;î�c�����w����qg�c��R�ȐwSG��f�ٍ�K!��+�V����.�2W����o�%6�/��i��ʻ]�,���<=��%I�mq��<��7���`%sZ���u	o���{�
j��#�x�S�(: 6w��[�{�.Z�R��Hr��{t���}�5���ٞϝ����s��}H�3Ɯ)����*���w�g.G��8P�/��y�K\�U���qz��g�5�5���d�<6N�P6���s���;��ԓ�MކS�l���T��hku;��xI�{�ֳ/��^ٶD��uЁ�j&���cm���R�
W�;��x�T݋J����u=�KB�t�E36\�E�i���V��6r���<&��}y�q:��Ҡ���i`���k`�$�E�BF2�/�i���e���g*����[��gר�c��!Fb��1���oq�N�EN��8v��}wى���Y��e�.�6��VU�Fgi,�a�S����GcGK7�0�G;�Ceb�h%��s�C��+j�$[J�Kr�x�/x���l�
�%��jGl�t��{�iU;���!���gp81:R��h�ʵP@b��Ha-�i�>����Ё9}�Fܹ|_w�U�9*Ro��|����[_��;�d<��j�&�&��;�t��d>�2J�he��S!��k�o�H�v������:��I�[d��ܘ�q�}7V����8�E0��Ƈ$c3�PQDx�����oq�t]aCl�:��6�qCk�9l�%�}�<�X8S�ͅ�zŔ���d��NY3V��c8с��7a��B�.=�]�Uw��^���5�Oo1��Y��
f�K�'����t�9�ur�M�J�|C�q�X�ښ̊�曽��`=_)�'r�`m"�Wh�Wja�Q��=�Gv��� 珟mε���P����7���{���ك��'��a~�Dl7��-;�f�}\�8;���¹�f��)�}�|x>����8�qb~�ɘ�nf��o\Y5�Ӡ�u&�른3x6����l�u�t��G���H��m�YEm�&ʜc_a+k���B�k!��D�eYZj/,�#��X6�T!2=6��VsM%�_+��j�dA��� y��A�����OZB���3Y��M*�����V ���=ʃ.� ��z�1+�"��;���R12�Ʒ�kݐ��9��+tf#C��ཫR��Wھz�.RW۽RU�����!Y�w`�Q��<�jRz��_��I��n�5�����Ӝ����*6��auL4i�'�;K��f�j\����U��c�y��5.��ে�<voS�l��.[É5��j�W��*<Go+��Fi�k�R�Uc-�V2k�y�%m!�T�'���IL��;�/!D��܉����
��݄A�@�{NԺ�ln�E��CR��}���n���r��ќ�A�<;l*&]�w\ۮ|B��2��-,, �$3 =����G;�m��0G��UE-},�:��/���ؤ��%f�+�A�[��u�vcA�NMp�m��
ˠ��bal�굯s��
�e��63��:t�W.S6�0;-$���W����X��ޠ�Q2v��.�`K����13J��ڐI�u�)���ţ�݃50���G9F���q��
k��]odG�^���-�5�jp��b�T���mLJ��ZX�Ө'�Flү���t�'����}�3�o>>J\�&n����xp����d�Ж��;0KI'��h7j\�np�$�1��%���#�������l�$/Y�T:�s7D��)�ݔR�w,	;�r�m �ݵN܅�wP��TO&�,{���6�I�C��)@G)���Wmp�H&��T�K��0e)=p�-�5tU�-��c�%R�Oa+��ܕ�1V3R���L?;�J����j��)��q�M,�wsp�d�C������==të].�Bk���Stq�X��-)]q�m�?f�9�V��4VS�{Qo��q#��]Ak�� EdxM큽Jՙo�AF����h�+vZ*Ta��g{oy��6Xv��}|�����=��</�F�$�wztxN�|P�'[;�h�J��z�s(��,�������P��D�x~�աm��y��S������%�������~�&>Jg��駭'��;�>C}���G�_B��կ*�/�a>�f�B�=��-eu��o;+�/9��ι}�{���8\v/L�cg���t����7S��	C����\�3�����	h�Bs�����n��r8�+�Ώk���R���%���k&����s8���݊_Eo�w�@��Y����i�6F�J����x	W/T�h�`��rq{�B+o�At���ݺz���0i�&�ma��);uLe�7+Y�@J��q
^�~+�����OqZ��eR`�9�E��6dѹc�71D�	�,�,\2�ڈܘ\Jau-��ݛCKC���
"6DWx�+��k���Hf����s�V��uis��-��v�:�H�����M��퓥�@)*��&c��R�pVm5��'���	'e�m�>Ӎ��l1�-Yܶ�e����s+�n�P�@�`��^�W�LG�O݃��ی1����{4��}��
bc�����u\�n$�&���V�W�ϔA��E��q-��ח��v��U�|�Dy�⚭����7ގ�*K�g�xD�݃�����*,����alU�N]3нS���g��yc�㶾�a��T1%�X��.D�W�]lu� A;��6�����h���|��%_<ӤLlW��:}���Մ�Z���S��%�PP2����ϫy^{6�t��P����fw-�;��IL�Cǭ^��h��}'r`�L��[����N�;2S���[��۵xg��n�6u}/�:� �[�����t=
����Ǽ2�n�U��_,L��Z6�:�YE��[�b�"��
�>�E��_]Y�iܩ�L딥��WM+��&T�Ħ��B&�-�\,��qK����i��r5��K�}ٓkw��.]͉�s\�CM�WM�6w;|�鷬[e(6=έ�)�,\۸ KNQ�I�K����kt�b>��c�wb}���=�@��(�g:,⸷�t��m  *8�a*�8��\w+3�+c����2*��dR�g5�����q�ЧR�����gJ��d��۵�_o@l���9�{ه�M�S:_#6�r#��*t��� ��	?��k�w�n��^[B6y�i�����6��͒ �u.M�X��ViLr�n��Y�_JsF��7F��g��Žv�u눆kiL;���#jQ:9mڕN��Y��C��ηV/e��]&�c��&-v��Ō�0>J�(}�}���X{O��ޏ|o�41_H-�.F{zQ�r�������}N�C�Ldfd}���i�C�]��U��Q��Bs����eg+��}�#�ِDu���3&颫0g����ї6�3�b����t?p�wM��;of��e����g�� �c�]0]��I�&��Y5>��O-Vl�r��a����dB��Gq��ŋ��%�KQز�w1`t�VNY����j���)Z.3s�/�6�\�՘��y��dD�и��b�{��ZA���:U��Pݒ�`�ؔ����������V�֦�=�:vCu��4o�7�L�z�jü�&����Z����O��-��Ns-kB��*;k�^L���z�=��vxWQfܔ:������2,�Fgd��XY�iI6�ɕ=���eA'0%]�i�ݠL�TmS᧪�.�����vTzyA�r��g��.v��J�{���hJ�&�g�3ۖNę��J�K�v�,a���5=tv��WKl��4*��w�o6�A�qr] wNC�r��ɶsZQ���oZQ��7	*�l��hc���;�j\펺T�׺	�g���:Ӹ�$���H����<pj=�@�Э�Д�W}Koן�H��.1�2��݀=���;hW^.K�R�Ga�9t�p˩��A&�ы��R������)4��Yf^0xX$�b�.����Y����	qr�*!%4�x^'��(���7��7���u�N�+w�ZNT�F��[rYkw˹"2s�^���6���p�*\���m�� xw=ue�I0$zz�m�����'`Al����;
z�i�GL�F��*p ��=7V��:7j�pfR�Y���rP���V��g��#��Ύ{� j��,��6�P�Gu�A�.1Ճ�����$�:3w
�ײ[B��L�W��s��θ� [�m��̻ƶ��\҂C�,^w(��hs�a�y�e�dԠ9R� ��#s@;�k�����h4-�vڨ쓑x:����uk�XxVe	�ʨN�xhƠ��_1$@�:��w��f�t7B�������)���ɗ����X�_g�6��v���wskH/Y�e�p��ҽ���CL��}�35ו9�:��X^	ˇu�zz�馩-�6�;nJG�F�:]�Ƽ���<޾��BB!!�!$ I;�w�s�1��~��mr�[a]8&�WbaYJ�\�tl�*��Bc�f��ȹv��3���kið��*����-���:V�dC�\+�i��L2�SP���(;�D��'��h��B�BJMM���|)�r0�v����e�g,�(8g�{ڴ���X�y���{�Ҁ7��ԗ]���.���7��M��FuKù��QԺbv���g�Flsޭ�����*��b� ���5t34���W����,���>���-�^.��6Q%��S����WZᲃ�����+�K�zi�#+jR=��Lfh<:��M��)�iT��}JS[���T{]�S(`S-�gLH�����H����Xuޅ-+Yy�-ڔ(��ϳ�A�R�՜���a;$30j��0h\ҝ����=\�C��B��{_G��b��������DU��=`�}����d���2q��av�K�7d�[�t�,�6��s�۷��*�
6�[sr��2���z�;�A������S���e�ʌ�Cv�g=����]GV�7��w� (m˳,E���Қ:Z�볨���d�n��9�wċN�:
]
�9J���Պ���]����md3����'K�I{�]Ӄ��I�Z�ճ�a���I$��n��U!˿j[�E�}��</o�-�#m�0R�B��l�f姥���)K��WPű2����v)!�Y�Ѿ�(���u�ԱǶ��F)oqQ�(�h.��r�����B[zܾ���I[�hw�z�3�.�1��/��tz�Xq�2r`CYZ$�)u�l���Kgr�nwu-�=]G��h0�x�m��m�e��� S�@�n0#�;��YjV�؁d��U�J�Ѿ�@�&޽����œ�oM�;x�Z4oXsud}k���+���aGx:r���v�Z�uݻ@�6��<9s5L��բ�2\sN�۽�3�!V��rQ-w�:!Ӷ[��v��rM�W|�i�oV��wo{F�S\7y,�wE��c��L�S|/e�8+R�����l�2Q��ܦ0k�u',r���&�7Q�0�J/uUX�@�u]����4̯�g��\2�jw���K�ZF���	��u��v�Iɫp���㵣F�K��1j�M�l�����ѝc�;�w���ٲ;i\w+p���B���-@)�7��L�����ٚ����9�w����6b}w�Z�A�<�E�����s�vݭ��9��v��w%��6X3PSz>�\����gZ���E-NY�̧�]�{s�
�0�k�9�J���#�)�E�N�Oh�r;W�]ty�[��2� :�~I��k��Č|rDy/��e���,W�(;�0����.4��:�i��V�I!�F�s7��'N��Y(����{����Vc��2,Yr�3I�7�`Ծ��r�x�rX�t�Iw���Ot���D�'$�W�[��.�s�~ԫ��=���7��/_vLj�控1kc��_@p#��U�S����y@�^͸�	Pf�"��]u�y����xqE��\D�n�6�ΤR�w�d@�b�仚u�A5҇f�i&q���x�� i��g[/47C5I�������GF��fŬ�$��s�"6���I��s�W����V�!���kK����ħ-j�=�ܠ��w��a8����j/�<�a}T~��s�����J���gCzvNs-���K�k~���5a���yV6R
	#���E�J��k�
7A{w0�i$��Q���Y��fb��k ��Sh'��aX4�j����L�4�0�����1X���D���F�g{]s�򭷸�u�i+ȂSiX���Ϧ�D�C��D�}�yL5�cG�ʚa���C�&�#�|n1=|��j��i��j���S�)�`��Og]��F�+��i�۴n�umųhn�p4x�M�Gg~�DY�����)I�t1	��S���8[����If���	�%Cws3��qK%�oJt�3�%����q�� t���BrܗO �8Yd��@��m�Z�b%S8�n̇t�����=a:�šN���V�����u�)��G�#��4;���Z��!�?\��'
DO�7r}��g� v'������u�o�9�4=<�c�0���G3\9����ش3�!���[ܼm�Y��9���r�؋Ч��};��/c^,��k�S5U�� �ï6�.���&TݩҌYc4�t��l#�L��
��Ԭ�Y�_+�E���*�hw*k������16a:�a~��\��e�ٲ������U;�Hl�����������o�rᛲ���<��y���P���x��]�=�n����8��,�"�y|2�I����Oj�n�纴�х�6���2�Ik���t�DFfa��e6�����b��+�o��ܚ��R��&sy�rm(H���yC^i\��wB>��P��#�ܹ��k��w~۹��>z�����e0��}��r���8�hH�&'�ASo�,M�u��,&��]�\���(�i���� ���y��r��s +�I�u|�1��ìv.��kW�����N]���Q��Tz�SjRWn�Ds#��Ĭ`�*<���蘵Q޼�y�I����Ht��Ʊ�΁Y�����%�1�\Gd��[�&-M���d'�	ۜ0�C ��܈��LT�;4k�oB��/��U�5R������J]�֑�6�c1C+��w���2�hX��8ݸ�pD��ݵvF��Zۢ�9��]��&e+��˘�0RY0_����FC�]#�^泂%}(��D�2��) �5zj�v^\�&�d�� ����F�ۍ����A��v��U��L7|�jq��G��Q���xX8ɾO��w�V7�Fv�N����M^��MX`��n���T���ջp{x��Pf���O���NnRS%ļ4�|*��F<���W������|9뷑8�}o�6��iQ��w]d�,�Swr]��H\r�07V�ۊ.�Q=����[^zuR�c��#�7�e��s��^>�Sm��v��9h�΅l����|�^�>0Nw���{&o>K�yڧ��{��vC:���曥W��&��ij��:��V�q�yt0�/���Y�8�w���(#7�JqKL�_�nn��JW�c6K���e����JZ�|Ŝ�uձ�Y�͕�	q,��}�ނ�I�;�=���{�O;��b4X�Z���3"�ߜu�
�v�q�i<�7@z�M�s�����l�F�ELgj���P�i�2��}�4/��j�7�=�f�WQ�.W��s^��pWڹ��8��4J�5�LQZ����:N�xY���FSޯ�ò�n��ڧP;�c8��bȍ��]\
-�ȎM��[�gI69�WnvfpTW�V#���iI�(J�A8�[h��Y܁D���7ނ����6�
�$,��X�N�nA�/3��6Z��1��#){�]��a��^�{�v.��`[�ز�F4R�9�F���Z�}0peT�����܆���IËa���hj+8\�
W.����[�p����������-;�_@�5��tEi�#N�4�	A��t��:�K)M���V� �̶����	�R��G��ӥ��g�폫���R���>�tkח�4[ɻ	.�5��)���yd������g&��rZ�٢��&P�pVL���r��H�k�� �7X�wl/�nAx�^��R7����9�b���"��o!�xN6(����G,�W��;W6$��U�����ה~6ɣ+۶������$.I�k|��4>m�뻲2���I�e�n���ǡoM]'eh`��az�m���Qѩ���ij5I$��.+������ew5V_��;��ol��{K��x�j��]���E��oQ%�y4l�Hǩ	2�m�zJ֒�!�S�{+�vQc�CM���Q®^�0M]_�W��Od�L"LpbA�������Qv�7Q]Ֆ��ԋ���T�]�\�_yg��;�L{o��S3T9[�5�#W-��EbͲ��/�3_�ۦS��!���gy�Pn�[t�">��v��;:��WyN�d:�G[�:u	j��T����\�^�ub��Z}�f�Y\3@�e	���ކ[˳+.���Ҥ1֪�X�ő�!���>Y���R����ӳ�%r v;�F��8]���.9���w[�b$N�7$ݭ$!:��D=�N�0�4~��%�h�n�.p�n�o�m@�R��R���9G�t�q�w�}L�ݗJcȩ.��e��J�+P�kvCs��˻��|qV�]��ĺե��~$y�uay�Z1�!�]ޛ�zYn���9��"x&�K7�*Ր�f��m[˱��H��}����Yd,�}��[�f����]��|d�0����'�h�N�����6��&�i�}t�v*�,�k�����{�g}�m����,���67�,�*�/��2[}�#�v�^R,��Bk���E���}m��-d���z�\�pj��3�$��[�sc�OHߤu�4^�	 :n��.�&�u���.<ڗـR�U�2����a��K.˞K�v}��w̛���zu��`v��Wl�r�\d%R�>>��1�`��(��rq�Ư���9��2bC��[ҭ��V=A�#����Xo,CA%����'��
x�����\�0Y�\֠1SSzӝ
|�N+:�C�zA;)��9�����������E��_7&$�ae�a(�� �� +
��[��vc�FQ�h�6����}�e>[4c���=t�Xv���eS�3��ͷZ��+]vbu��.&Ό'�Rr�<B��ܸ�����p޺�C-�5 <
>�XF,�g���yI��^$�jn���B�1��^�f.{�(��S]ȦH��Ff�i��߄��8�r��Y�@�^8��Ĵͬp�O���D�����e��A�f�o6upS�tn_z*9�3xD��zѷ��19RoE���q��'6;��fT. �-]�Ge�u�^��+��z�mD�,���f���w˷��p��r�f�"U�(�(�9�I�cq��&���P�o*{Wv	�l����o�r���.R�^��=��B>�6��v�v2T�����9�y�0���~�̡�Td(�p��j}�;�#}�wU*J� Di������أo�N�)�6*����w��1m�=��-�B5��w�8�(��"V;�$z�H^�+Ł�]ZF�B%�4|W��Mȳ&"=���$�pd��K�I�]�8[�'����ʉ5n��G����}� 0��W����u2��f�W�k�+5v�-7�=븠w���*���������~u�؇ի9�ٜ���1�"��@ٮ�[��Yp��}�.uL��l��FTY���%�(ڻ��n+w
�w2���6�'J�L���=֨��j�qb�<PkC���]�˟��d��Ym�\=���u�e"爧VS7��>J	t��#9V�Yy2�ڻT>��-���rh!o;�����1u�����B�Nf�v���EY."H�^�3[5�g<�\�׉�n1Up�ʢ�K:����,�͒������ݍ�m��d�W]J{SKww!I�(e��1�n'�����dY	�
{&T&V�ƛ���Ҳ#k.�� �w:yʦ�*�s���n��n��W|y�� �����{�8'�iV�4�53yL=�Ǹ�v�V5i]����ͷ����hv;�/�m	\�^ՈRUc��u=8�K���m|�LT��R)y!�Xe�y̐����5w��"֟�똳h�G`[�+���R���J��H���CpN��j����va԰�&�xy;٢��O{�]�Q��vSm���N2�q�ܚy��D��SJU����+�;��۾(o�Y��%�0������`I��'�
q�A�x�N�^�3�m���S؋�އ��:��ՋHȫO`��Ĳ�2�]H-B��z�$���$��^�q���9�u3f�Y'y4���Ӓ���Z��Y��"�P�-�5��k�0���8�
@��w�����'��95�M��c���ـ��s勏^�/�]4��NA�6^7���;��JcÕt���N4o1���juĩP�9����+�3+U]� �i�P�A�t@.����ǉ-��}�a��v
���+^Y4��2l�������o%]"�^��E����;bޚnJ�� �O��f�ֻø��HF��;}�k/ A���@M�h���7CEFOgl̘��)��a��]:��ZPB��+:���<�a鵉���M6+���[B�u	6ݼ
�p%�	bG�҇W>�k^�[�����Y�anit�fS�	TU'X�j����,�vJ��Z��씊Z╴e����'�n�<,�~��Q�9W�.�(����ׂ4X�_��}s{��*ۻ�����ϻDvnH5�0��ނ�;)�G�ϝ8�����+o)=�}��QW�v���H��=z�zU3V{w4ˣ���Q��+�����"��hcV�	���GZ{��A4tS�]��Y��]C"s�F�Z�����q���<k	���FJ�
Z�!����9�0Z�f�7�hN�l�ǓFt]'ٵt�W�/��"��V����P�W�/�X�-���8!��1���&J@I�W79&>P�r��Iˎ%���N�'u�����=���nv9�����p�q�����g�D�n��yu�fo>�Y�7�|͡���wse���X'���׸��h,��
���SMެ7�]@D���oWu�{]�Ēh��ob�s��C\��c��e����wVnp�:�C���5i���6��֚BZ�H�0^�I���SC�5�)T��2�=/vQ�˂7������t{9L3f���4E��k�y<�|���ϑ�z� �$�[C9�(��n��m��vs�V1�֩sd���3h$`��ǰ�汱+�ܹQ�0;�*q�WTm ���I�ܫQ�5һ��u��j6�k۵.ֽR6��a4=��v�E��št�mՙ}�ew-Zx��5N��x�V�ef�:�SKp��\�G,'%�k��Sq��N�n`3�ά�v�4q�?���)�y]�qS�c����ä���V�����ð���ƚI�OBc:r��+��۸M�!�33�rѝg��LS[K��PX�&��9V;�;�ŢU�1c8�bT�=���qt�Qo��/@����F�n�-�=�ص��>�%�ы�!TF�ɡ�v_	��P����V�SXij�B(1�!�o�M��;�o�wW0h�J]�3<Ի�+��[�i��mh��y�){|S�}�(�8h�|�@ޯ� ���bN��vn����8o��/OK�v����Ǵ���{�~Sl��ڱb�Ub�*���ѭ`���EQ`(�>!Tp��֬Z�QE�-��+0TR5�QAiJV��(��"��kEAA��*X�PF$X�hV-B�mV.X���U\2�A�mB��ii������Xa(�kA`�T�YZ��T����lmU�TV,��*%F��1V((�AŅciQ��VAbR�2��Ū([��**(ŐX��aF���`+JYX�m�EL&(�Z�
Db�%f�V)�J*b�)Qe�FE��`��j�b���H,qQ�H�(
%�[h�+(,�,\2\Zņ-�(�����5�UV�@
 �(WҾ�K��ތ���P�r�+��A{�`F���%�]`�|�\5��eh����g-�SJ�&�����m2N��/��2�-�N�5t�:�l� �T:�9.���e#�_��g���	��S�ش��R�7�,1EUyF�c�tѾطlH5��`y �c/��!1հ-^��}o[��;�>�8,�}B��&V/��S~�m˞���8=&�ӾnQ&�t��r����a���:�I�8.�������9;�{C��Cř�;Fs.�[DUj2����]j��z�����X=[9��5�u^0�gJ]40j,e�N��]�B]�rvj7 ��{Vu�*��А0~�"Wr��ڸ�=ONz��usC΢v�V��\�����R���x��4`�>���.g��@�I���9$u@��r�NQڛ��������ż��O9Vu�g6 �֓�BEgnT2��&:��-a�_w	H�9/M໷΅`8����8:A�t߽PD��A�J,K���%Q�J������a$j�[]7��Y ��t�'}딵Cc�U��^
o�C,�`l�R��|�+}14,2��/_�<�X!tϬ�;�9�hq}���3�Z�����SQ�5��[�~Lo!Y��Y�e4V/P��ĤԱض��z�7W�]�j�S�K=(���d�w��P7�ю,:�-S�YB:O{������ᖍbZ��1��i~co]"�	Vn�R1@2"a��%aUr�lF�aB�V��9
,i<��t�Q�2�ɰ���[>b��ڪ�YS��/��L`�j��3[WHq/�5�[`�ULz�]��ж�z5N��v������ғ�-	r���X0zn|�[ꅸvS���9\�n��]-pV��]qz�UC�&��c'[j�%�;9$f��σ�MU����y�l<��Z�v���-�`��T�՚�����:���~�0���[[Ed���3Hԫ`Nf�#��ǐqM(��<&��#'���W B�1;Ғ���̡V�1X.��"{����J��K�;��3 X3`��g�\�qU�d��ü��wRfS^�:9g�wL^����1O/W[����ӷA�&V���8�{��w�m���hpu~TÜ������+��������4{��^���D'�W�@A�(wU��;KNE˹B�Z�	��鎍�&o#��|Dl��V��s��}�呚iL�I#�<�q�ul稁���x�W���m�����6+ּ;veȁ���KB�;�1�v�N�B�;U�]Mco4��K3�X��$�};�NjŰ��cBMu�Hq0»�'3]ҷ�շ���Īg�wa���r5�e���:�8ρ�V������������R��;2�%�+s��Z��-���/�u���X���׭^�M��ݳ�� �Y&�DQ��q3�z��	5y���1IF�Ѱ�Ps�o�@�Z�6��,�+w&	�ո���.�τVQ���:�wםH�摑G���c�pv�6����fF����,Dƪ���`���vs!�՚X�[�s�&�h�:�����|mu�"��a^ǲ�(Sw�r�_����
�)��e>Z�������S�K>�pN�.�WV8�7>�pE�j�5ηͣ����y��l���i9R_UoL%�#���*�6_�N�*�w"=aઘ��}�a����Î۽�Y=�[�{i5c:(v\q�
J��砦@�ku�ƺ�Qw�i�^+���&3r�Oz�H��H�i�N���څ��1�%�f}�qN��,O�x�%o�b.���Vk39�a�sA�R��9�ª�����^�̿���U�W�C�EHo��₻(�X��;�����Ey�M�m����5\b�<���Ȭ��`o�S W�k�R)L�z�A��������g_X�񈦒������T�r#��{[n�=:�&zE��H;��������%�*m��.�(���gR��`w�M�AwY]�,s�������p�-�x2ڴ;9L�T ��ڝ�����o��&����=�3=y�鎮/��%�q�E:�1Aq��~sN�e�dT�6�1X�X�)�i�ы�]f��BX^�![����:B�l���t�,s�b�53�;�t˳�n�\D*����e��#�\�Ɲ�ږ��d���J�QƄ�*�	.�R�6a���j���R����Gpi�i���2/T0m�S�f:�S>{P��B��<�^��(�(�9P�n�':o�Q��]����NG�/��}�X"���͇Q+�4\N�x�d�!u;����.�l���<��y�Sd�Z.�����0PXy����uV��1|��;wy;+V��r�ۇ����8Ç9(�sd��PQ��m]4<3�z�`zC6N��#ض�ƥF}+��%YF.�89[j}�0���(:P�t�),�(���Z��^[�<Ӥ�j�/OPn�+>�]	���K�8Es�9�2%��3Cv�}�QU]�K���(i�`��b��m&=7�򫵧����VDo"������;�� ����%���!�}˸X͵��W��/�N&t��3c�
V'�p$�Λ8u:�L�^�W��Ý�SJm�Yw�op_)�ۥ��w[�uk�2��@H1�	��d:3�NO-��=9�y"/6����uS���BM�Cw��1m�}�H�t>J��|��y���qv��hW��஥|�*��T �g��&{F�2�x�.C@��{�J�hG�!<9�2t8�m ��U��LX�E�H�SV�FW;o�h��7��[�Ν�
�Kj��ۣF�C�*���Ӕ^�(�K���o�g��R�&�VU�Y�{}���ٕGؤ��pzG��P��8��LJ�"�uxު6�WP�]0�=�R�~W&·��s"�T9�8Z��Ʀ�i�ا]ƙ	��3ڪ ���I�2��H�>^�����y��ܗ	��Q���R�f�%�y��\r�ި�lH5������m��u���������A|�+"2RSq-�s҃A�p��p�-�I���ށ;�ms����V7����OW���G�cK���hk<40�{�V]b��Ř#��k�����1-��Y<ɼMr&s��W�O2G���g$p+�C8�\�Y�$<�����o�8�ky
K�B�	��[�!�������Sӕ�{����z-������Ӧ#���Z��X��O#�s�!�"6�ȶ�U�ׯ�e�/�S���ڟҸ�Eˊ_��v�y�k0���sT�_��_Z^�t+��}kUODV�-|�ï<��(=�w�˻���X�T�T��+{i�fq��&#jB!�`=Q�ZJ�S��gB:ao�0�u�AK�a�U�����:�v༩{6�-��"�Jk6GY�.�r�lY�LpY9�a3^NX��UX�B��'�\@tGW���T�v���v�M-Wny83�Q<WW�d�S z�YPD�xK (��C�9���UX���nݵȻ�2��Wcqv�D��V�B,�|����=�j�P��V�|�+}14�IU򪽍���z��P��;�U�����1F3�������q�@�� �yj݃��1ݲ;��^Z��Q/�֙�F,���}�Xt+�1�:��>�K�k���.�^�=
.' �n�x�*"9<�Қ���i��ϊ>.Pe��y}��[p�D3jL���3���u�
G�v_�]STX�j�L�7]�E�U2r�ʤ.��&$w?S�2.��9�onZ �j��mA�qf����=����^��X_g<xz���So��)�AS�I�fu�~ˮ��z�@���ȾW B�1;Ғ��Sa�O2��,F
�'�#pv��ΛX��h�O�j�cbOV�]�Em=�
�q�K���n�^s����4U��A���f��ػnowɥ���xp(`�=�b���;��e�)W�6vp���k-,��T�AD��Ù�p-kaS�)�d�9��Pj�uZ_{��3��j\f�ZRK��C5L�3�h�L��"�-�M���ư'u]u�9l������y�-�c�)P�ݱ��*$����qn�-VET��Z�Sr�)�	�(�m�U�YY퇓��44l��C!�<J��B�.�@�����=g
g.�
y�a�n1�㶫|�P6�<F��=L�Y�vY�Mrߣ4Ҙ��H��a�D�`��V��Gl)�M����R[;@^ܿ3c�%��g���~��ڭ���S�g�J��
&L>�E���=V��:=Ft��{�F�Q^��|��O�N���L��ٸ$�^�h���O`xw,�!ގ���s0Fo�21��R��y�~v�{)��
�S�6!��w;�r��5	�j���u5%�1#����q&��^{)���9��K�o��h�"�V���q�+|L��Rt2�s�u%��5:�|t\�M5]k��k���į*�wS�](&�=W�ĕO�a��ۗ����-H'Gt2F�L�ɍ3��N:	yXQ����_��j@��J�vZ����㏯�8V��Պ�m�~i(�����}�x�k7}P��� ��}H�:���=C�*�4;��̰mA�k6]���㒱�}����W�C�f�mx��{�sX�Բ�OL��Q�h]�iM�����Ǝ���U:���*K�d	���u�ɬyS'����</r�U�W���ظmYj4���P�v�6X��N�>a��,�6��4���L��6NI�'�S�2��}���="S�i#W�E��S�%\l�'&4:�L꘿t��,E��o#����}Si�]ֶn�`~������W�W�h͐�m0'%2{�k52�Q3u�@>$Lr��cs�f����b������t!�p>���1�7�C�z���7�K	K��nמ�6���V�2�顼G)��l��n��P!�/�g�-�m�⪰�=�/����%3њ�2K����)L����I� ����q�<
��a�K��T���]�K�fM,}*
ǰ9(��هS6�r͎�JW�Ԓ��ڄX�v*ď3W�ijQ`��ƊuuG�����N%ܥU�؄
sH�g��-�\�u+�4Y��3!O=���p���$�H��{��~�n��w���	(��}H�	���B6{�1W�T�
:�Y[ ��Q����V=��pEz���_�$ߺ�Fߛ}��*`x�n����EJ�������t���
)���d���!����vlvdf�������];\����K�+Ƿ�u�Tw����j�6�~�F����a5�+���ܾh�
�ms�DEҏ�J��g�7��e�5��.�H�)8�����p
LưX_M��0*8��M�ۋ�q�c��ݕ������po��x:�7^bk+Zaw+�J���`�N:�L�1������>��V���*�5���,�ı���W�ל�MP�z	���q�{�k��C�w����t����د�2�swvS0J�=�m�i��E|6eњ.�iݵ�GǞ�u�S>0S������϶�ypWR�QW�T �kvp�t/�R�1Q���,5K.댖;O�gA�q��egZ�<��w���Vy�qC���B���1���j�ҋ̼ى��Zfkѯ�D�F0A�yw�(�'oi9/��S<�W:e�&^Z@�m�W��T����`�o{#��ẓ�<�%jW��I�+�fP�϶�@}}2��ǐ��ub��JF�̰ŕ4܄��m��S��L�A��fAw�W�FJI_���_��\T���u@��\�ߔ�ٸ�u�c�p���4o��
��`e��ڷLB�s��J;��Ɓ����Փ��I�����՘�$'��h۞���du<�uu��7'���S����mX8�@p@���6;jqs�_J�, ��G1����ڷ2�j݀Gf���ɼn�p�V2�++8G���<LU4�=�
e}����r'���nBsb��qw�����Kn\������N���aV�9˼Ʊ�V={9.������,)�tg�Ixn"�|��`�we)N�z��Oi\��bq_����m�ȝ��9���'ڶ$X�w�����gM��!�`׺b�i�b�GəӍ�lP��<.!3@�`d�v|�aj2u�ƭ�ׅ��7�ӫ�v�Y���u�Z`N�J���&!]�п*wl`8@�I����H�����{6�uL闖�ӝ<6�@���1�IvN\	��G�S�/Ϊ����2|���8��Ø�qv�*���U\�c"�q)�i�F����:n �y����J�����躣�A�󹹘����-��n�%S�g/)�~r����Tv R�����V�:���b��Tz�u�M�"��C�t
c���a��Z�>���1b<6�{1����|�2�+B�۷6��z5Ȱi�\�ۉ�{�i��b�}(c�
�:̙���+|�V�{](�tʭ������Dd�5�U��#��̫g�>WE�ν�+e)V�	u�NV�Qg����:�9��V��gR��2
"����K��kR����%���qc@l���|�j��W@ +���D�P�ol�ҷ(n�vi�2@��oY���@��u)�
$U�ľ)=<���zl}r�y�W��O�iC.����Z��u�iǁw�c��7l�f����+GpX�;�e�o!�we�,Z�8N�._\�:$*^tFq�P�W]/ZV��6��{p�����"��[�;sgpu��*�
)B�X0��Vt+ �.�������V;�C&Nv7tiʎD����"�*�>մݞ�� t]_wT��V/R��2.&m΋s^��nV�`�J��}x�]E1�B���[��voJ�T��՗1$���\�|M�7c��h�õ�RoT�R}���>��I���$I͝�.����rs���	C�l-{�	��±u.�x��'$�M�V�G�����/VW2�4Ӕ����Y`���{�:��®T��"ͧ|Ú`VpL%�:��5����5���3F��e�C�����e������uD���G]<� ����9r[ ����.�ĵ}�}F�`'�Dn12�L<C뾆��Mɿr'G����9�E��ξ�ҙܫ�)�5��Vx�A�-d��'*����Z+t�$��;��&9���2�^X�B��tU�Z�\:��wL�ڸ�e5!�����=R]i6z����u 9�]q��i����U3��
����v�HfGժwu��ČV�����֮У���>��GDii�rgj�Ecf�W�v5|{ ~�q���t��txV���Y�i�Y!�vaB�s�Nh4�b�k�&byX�]Z8;��I�4�����y"ޱ�@��z�sV��I1���6PhY���ɼ%t5�)թ¹�F�ɷ�#v��𻼼v�;4�ki��$��vizy]Jgn��>�,�\�{��.`���z,�Ji�ƛj�{��W��۷k"��r��R�Y��0�]�l����܋�%A��m����W� ���3NBS�euE�Nj0{|��8�7C��o|��Ų����k���8���v�|��~/b�c��$9+�O{Q	���YІ��D*N�)�"X��-"z��O��0�p�N���������u.Ý�#֩Z�|P�����YO�]��	L���圵[U�V�B쵠��E�4�9,�1S6o5iG%�9oX�k&��p�;]c5����N	�q��!xF}'�UA4>�wF�OP>$��6eu�_=\�})K��6�L�;ٝU�b	�=�)���v��&F��^�xz�{ʥ���y�e���5�՜�HR9��d�M�S�,Qe�_l>�V��f4�]�$-��z����eof���R�$�>�'�Z6֤�,R��X�PU�+qG�jA�i)h�`����TH�FŨ��b֢ʀ�j)iJ�iV��mIX���m��E�%-��am�j�h�E,bZŴ�Э[K*V)D�Z5*��b�X)�bU���,�ch%*��6�PR�dJ[E`�j#*D�UkUkZXTU������Z�l���0FJ��hV�Rض�iD�PX��,-�*Xʣm�)XT����������()X"�Z*��ma���*[b���+cJ���Kc�dX[E+D��D`�kj�mlQE�eJ��[%TVҵZ�*�X+lF�T�[-QEڊT-��Z2����J#ZƥF"����%+Z����T���X��h4eU��IJ(���&�Z�˦�oǰgT���|A7t������o��\V�s�~6͍�z��K�[xngS�˒��4X�
3M���o*)v��G�5 j�U#Ɠ�3���<�L�3��M��h8ʍg�J�4a�����Q���Tܞc>4&eMU�f�qq9U�c��mW���"���9l�B��螴\���s�ƴGYN*X�ƽ��O��c]j<
8�De��kw����=Kkh��#��
.�n�+y��sap2�7u�X��;
"�\
�\��IIF��<��� ��{�yl�1�=���K����3TΌ�U�碮@n��D��@�J�����q�N��Ua���:�]�{�!�_v���&TIX=�8w�;�D���mX��48_�!P�[�-�;�)�hp��F\9�]�8&o���	�VBc�#���8�-9�3�3.V%|��bg�>~W��-�c��4mS4�ˌ�M�֮�%��-� �^68	��ڷ6�vTB��R���e�1���aTzZ��C}�ٯZ���s2/�%E`dL�@�f_�N��ve�M���B8�YEt�D������өL]׶&˫q	���ϴ�Y�����
�;�mu�\B����C������t(�d��K��s<��.�).����b7����p�1��j��P�LC��fy�J�
�����wY�)�8N�9�C%#�<�zNÈ�L�7�Z6�zbn*"{�"G��{�3���wm�F"�Hc�Tm�3����[��
ﾢt�l�8�NR���iuNN�Ѿy9�����
��O�����igWT���b���;{~�x�R��=iW-&oX&(��6[�X+�
��
�gp53�S�E����d�,��]�4�&��3�>��%����@S��%S�۔��Yl�5:�U3�G�6�\p�++N.�Z�:�2��ۘ�����Y�$,5\9' �@�ku���<�]_��v��v�hr;�c6u=>|{�O�˨|��P��;���%�fєf�c�;�E!�MRPz���en��R�w%D{� ����+��5T^K�P��e�S�6���D0͒'Y.qN�<�`��u��o{8h|tS�k����ӕ�d�t��*����5����OT`�A=�;ҝ"�S4;Z�!i���:�	�7�5���'�o�eZ���M垔U�)�����^�Ӏ?<� Ӗ�V9NP�[=Ed[�$�@T���(�\;��T$:K�W�,h�7�	X�>�[��Ýpl 0�n-O�n�aL�xɼ.�����.����w�b��j�fd�A����s��_|��ۤ�=�=�|k�9@6���6���ʹ����Ց���,���'`�Y�6̢���;�ٛ��\�Zp��J��㋷���̣�M�rٛ�O�5� �U��Bxr��R�1x6����G{�o���[Z2���M)��cX���Ԓ��ڄX�v*Gw�~�2�d�o�4�O�:��[3���D¾�08��(<�]���:�U�y���|*���T	��f��rE�ݦa-��m'�B��;LA�Ai���L`����ʑ��T�g9�\
��l�~n��i�S�R�f�mxmAF�m��~��麃��@`N��*av��ٻ�,�H`���ҷ�e�X!��uP���o�hJS�ͅp1���L�ٜ�]B8_wl�-�8,C�
n���^�@	�s��rNQ��j:j���&hm���	�m*م����F)*z���ux_+l�_���,�3�=g>�NF.�F�|"�T/�*Hd(��i�=S͞t_��֖pS����w��5�x8+�_+��uB��h��:�G<I�Lwu�[G��ѓ��g��l�Ӻe7i[U����F9��ut*y��}�A[c;O}���VǊ�֮� �}$��1Q����8��C<6��q��ɜ(Y:��"2�;|�6b��U׌�oC���=c��x����j��7p%���[3�w
bV�K�>Ku�/�nⰝ�� `���'�ҍ>L�۹�7��c���T�xx��<�Vl���9�F��C�'=vӵ<��|Mz��O	��UN]�Q��J\uO�\G+���F�~9��i���V��TKH�:�m��6=��_�b����].�o�G��)��*h1���m*ᮝwg
�ϰ˽5��ٱ�.Tg���t{SP7�{q��P*1W36���u>{�pM��z��=�w&i>�yg�3w7�L�A�:6+�dw,�F���.�2RSq�ۛ�]H<c��)V�@�0���8��2N�nx�A�`X��td
���>K}U#��D[J�t�k:�&���Ĥ�յ:�^���W�H|6��"V]C�<�v^�L�a4Z�p[R]$��YK����C}�aB��q��lP�;S����r %pr��d��[q�|,/�GE��{%}ݎ�׵����V�6��n�>4;3r��T� B^N�͜�:�������lw<y�*���szns;��Z';��h}1�IvN_��f�S���;�;@:7d�.�\�����mE�'�K�Q�T���'q�0X�^�k��>��8�E:���+R�C�ǽ�*��?E��f��߬�����/'v��sV:�9ј���ņ8��z=@�r�͵ �G�h�lSw4�ք��}���y�h�����" �Kw#��$O2�����z��'��'���'���lL�G�/Y������S�{go������hh������g>������5m*/e�P�����˪�`�iݩ^j���9+�R|�C�`�>cՆ�V�Ϯ[���V˶Y䪍T��>,�U��f�d�<�3���2�w�i��#P'��u���D+݀��sw==[U�X�AÙ�)1�4���^��w��v��|]��3���7Aʩө�k0�6�� ���+�2���1�s,s��*ڭ�9	�q��Lɸ�f�wp�@�B�1<�)�3�Yt��.
�aP'�i�>�Z��u�
�q���ai��+-��d��oZ٥�wWE0�p�fiu=E��d�^�@_*���Ѧm�P۫ߛ�q������l��S����^�υJ�Hs��⻉��n,����#=g���!%51�6Ӆ�n�����f
�r���N��Ժ��d�]0�o�r��Fm�����hpׄw�����M¥�kll�q��x�3�Pc>qN!vS��8�黫9��\Q�J��w�h�ϲtr�|}A�x��(�R�^��,]aR�+��k<:��Ќ�c�Q���K:'/�W � ���x�>�o+/F�$�t;��Mh����M�yɗc��q��E�c�f��CĬ0�ߔ�����z��Tv/]�⫳�Ȼ7ua�/�w(W�[�!�}:��U�
Fމ�]�: U�c����ыtt��J�[��n��
�Āڶ�t�c'T"��+��V��>$��z�`����>T��y�V��vWC22~,,��^����i�<�TO��Q����7C��6~�qV�s�)���Ee0���9P�6)x��|��X��?=l����^X�4G^��>��DY�3�n ���Zκ�R]Lhf{c���A�s�~'�y5�Պ:m�I�݁�%#���ƪ�y�.P�o�y��@}�@�c`>ӂ,^��Ct:bm�������.ل��mY�'���;�Y�B�y�d�s�����]=s�n0M잎aoS��8��ɍ���\Hxk�\&�T�5�}��7��4��:�G2�)g9�y�T�M�A\C"wOeKNߵxR�X�i]���~2��)�;��w��[�1-^�	�LꞨ����'V8Lu7h8�D�(��U�ĕ#R�[w��{5�=�U؅�Js������
t�۝P��9G���)���=�{�ry܅칅U�|qH�O������;5�$׊\�K&�i�V��#��Y}�+u�Y��/���6�ס��r�������&�A�cj�P��\��������x��(�$���=9ﴎi��m�����ٻ�b�=��W� Vr��k�����.���f���!
���#��t:޷�_�����!�r�~����(�t�K�C�,{��)u�	qUc�!~e��Vz�1&�*CcU�{o,�ћYa{}�����PU���e�N�^9l��O�-�����	�U�Y�ݑ:�*H*׮y��a���?Ur��U>���+�`��-���X��j%���/��<}#)E.<���\�GIfp I�7\�~�k3����͇R��E��w�S�d�1��o%���|�v~��"~���F2�g=(�&|�h��&�mӸF
<,����8��^u�"���/`����B7�Jp�R5��1p�"�nl���j
5ںhxv*�����Tk��Ψ����c�~*p�	A�)�C�T1jr������6cU�藼;k.:��g9^�3m5]:Yd�n;&n��}�@�����&\�r,��A{:���1!����3Kvq��}�z�Cg��]1+������+Yt����O v�,��8�M�JPPr��6:�{*�;��}v��SQ�z;����������bg�NX�;뺩4!2]	@	�b��$���k��K=3�K��CU1zն^u��4݇�dڊ�t�߳m��e��wvS*�P!��BH�N��[�ȥ[��v����wF�킘�\Bт,���d��bp�G�ĩ4�3)�������SM�ݲ�-7g�մd�v|{��~���ցz���(4�r\Q��rv6>$��l��呃)�B�e�T��<F�9�Ƽ-O%�(�m�S2V�lv�4�eh72�`U��I�f� ��|5��U�Z�+�h��Xx^�+��A~����o���5V�t�DW9�mL��FC���x۴;b�wd0Y���o�Y�a1M���+*)�P�Dg*�X����7��:�p����;�;z�1���^�j3�^�lPe8OWF�p����6��T�k��)Ukޕ����U��ջXW�Kt��S�!98O�R�5��0,t�:2IxcK����9��Y�=\�f�.~�4�z��[^�!�dOfzݯz�#c;��i�u��Yb;�G���e7��3�z����d�{[����*[;���V���j[�o5�j��n&��y��o��G���E�zŰ+ZǱ�͈ބ�1b��Z�C-`���'�z=v7:9�p�T������3pq&�kV{��ݟ)bkbG�?a���	L������U�)��������k��jӐz�'��Cg;�8:�d@K�r��-��|z���Q7�3�̃�ū�:b���^����N���L1�b�]T���p�
��sg$����NG�f	\�{���O��v��@����[1�d�	��Ge��UX�^�e���ʨdٲ�)|�֋��m�v��/+�)�vsx���M`K����bQ�Xwx�n;�Uv*Y<=[�~>Ԡ�~2�	wta�
4]�eMVr��s�yO��`��Tl�
D_��Ѽ�n��y���r�Ȭ+�zC����cȺ�q��L|ǫ��u�*՜��xn���{0�;S��ձ����R�J �O 
���M�:�3Q��v0J�
�:̙/�i�}�k���%«��Zn9Hܑ�I�;&_�1��UX����O���e�;��Σ�����:��*�˟l�{P7�,k8�X뇵-9�3��q��&�	�S�ĳ�����b�Y
�5�A��!$Ћ���9)vU�lUl
bl�Ok��w�.[�f#6��]��'�Y��-A����n������ڴ֓4�E	��>;�O,�I9�}��M$r��m�u����6������*�{i �'F���%��y�^m�iѫ���[9�CK�=A�Eg��Urqxء�L�z��x���������X;��[�:����^	��;@V��� ���+�ʖ}��� ǋ�x\�W{=~�>y�G}H������u%g��o�Wq3�]��2hu"'�y#�0����oTt]�A��ψ�BDnl�S��D���T!�w,�AuB�g�\nC��g*�lV��]��V�ī��Hq�b�_O#7:����� S^q��Z�g�q�K��`Mc��e�]t�z�i��uF�>�6����B�Z��0���д�֮����ZS=,�G@Vq�trawM���=��� ��y=D]8(=�j�,E��_ӦJR��O�΄����k��f�sKwFz�VIX��
&v�DQ�6"�4v֏"_9a��:|S�u��S���u�T�l��ʧY�{ױR���7~DtYb$g��Xf"�2@�Q��ȩw-`No9��̸J�WV;K�� ޳b`�V�í䵃���x&(p�6���@��g�4>�{+.�?�-�����KC͋HSP�W��<s���݀�x5�cl݆C"��g��押�On>��{E.��E4�i�P]v�j�3L(Vm��+v������dTFd��_6_DUM�0��[է@PC��ki���C$�O�h#;�w�n��Y������~pc����֝;|@�l��J���ʽw#>{�'�i�z�[HܥϺ�>z��z��X�h���<��m���Է��H��̨{����Wq�L�^(��p��|��}b�[�j��D&NV��M��N����t����i�V���&����H��E��7ؼ����/�������F��;�Dr�̍|��P�;%%S�J��w��P��F^�m�F�����(SYW��Jo�c���k]�'f�t�U�r�LP4K*��o�>��u.�;�aF�<B�r���)����f�wi�Y��Cǧ,#��� ��걦�<��!��Qz���"�>:��+���������6�]�F�rp�{H1Y����}��/,��
 ��+� �k��L,.��y�D(�K�vi;�B䆡���B~>3�!���\��W��\}�t���ۓ��j��G5��ǹ���x���;�2�I9ʳ�Ԁ}kp���)P��;oO����˒�}�_���w�U�B�q`��ѹ�If��`�2)�-Zڰ�2���?'J]6gL4{5��]�r�ܚ�~��̋���$Agt�^gr8f�����V�.��"aS{;���������@�!�0�,��/�r�M\j���#��qU��޷!�rA���y��kz�=/b�����	�X�yf�i�J�a�V�O�GK���Ǭze�S����+�6�]��y	#)�T�݋z��v�Y|+�s��N�,��?��h�8k��DB�\	�U�h�#�ќ�ײ��\�r�ϹU�̱9,8���v�K$(_�՛���u�K{����T;E�G����e�l�Y������˗��ݶ%B��άz���5q��A��u{�=xuc�bb�m�u���2�ɽls�+�*�k�{�Hkjj�t��.�Ǣ�em텫��pc�%M��j�/33P�g�z��WTTҤ��d�>��ΆȌ�ՆW`ܽ(W7:��T�G?�6!{�}���bE9���wɽ�ĚN^�dە�܋{<v��,�nj�oI�k��D�g�oOdw�����+�:COnR�y��^���������c!dǭ�o���6p�K�w������*�f֒����e=S´���>�k����]�U��e�uڶ�$P�Eb�t�{8��N⻱�rh2�b�%����+����ByB"�z�r�>��	4�hΑN���Z��yg���F��d�cͩ�������$<����n�n�
n��=���;q\ u>EoD&�;���X�ZjN�v��H���ـj[t�M �V���ԔB�m��KAQ�)FE��bV�P�#iV�0AeD��0K[b�[F"�V�+Qj
-TTQE��Ym�KDek%J�Р��c[m�E��,-���h",KQ���jJ"2�m
�ZVh�E���m�T�U�UEb�k*�Ԫ�����m"V������QQ-�եe+b�mUU�Ńl�2�����j�V�Զ�YF-)b�(��-)X�*�*������[DFЕkR�ʵmaUPXƴQAm���YU��b�Z�Qb��F�XT)eh��**��kiR�TQ��Ai*Ҋ��*����Dkb��ЭQJV�A����V��
 ���DD[j(�mV[���V�mU�T+YmUAUA���j��lm��"��V?n7څ�7Ҍ���׭Vr�g]��Vp�2�o���(�Q�1�
�@�bo|��]AѠ�´�vg3J���J8ޏG�6�֥C.�U�d~���׵J&iKuT �F�p9�:��6Y �P�T�a�5��Ez�/ˡ���꼠�ho��V�e_\$�}0�r�������B��[}	�����:�Ü�h&�Uq3�&4dYxj2��Y!�ip��bj
d	��X �4v���\�op�,��J��N�3��p�DT��P�^����Qz,��U��v�ɬ�[A�6�-u���d\s��^{Z
�-�����W���X��U����:�;6���ʑ����+@뫗=��97��#���q�h\���z�@j�6�	G������rVb#d���4�R+U��X�[O�#��2��}�����n�s_�M�ߕ̥�L��]��������`:�/
/�����AN�a��R�LI�
��	f���r��iv	N�O:R�����V�2�'4-�̿FO�-������4'�R&�u+H_ObiWV�휗Z8g�<�U�%b��T�{����Ӽ����ޖ"��j%S�(�AN�����uŕ�����?pb�٘1�ye��2fk��x�iR���##��[' �m����W��b�G_)"�;�Д�f;�}��$���r3�37U~�Ն.��&S�ؤ����}��;x]�Uv����0w�p�;�d��^������
���c��#o_���.Y�d���C���}�`"q�t�e`�{�3��w3��1�Д6����-�b&���j��,����h��P��i�!�����)*
�hj=�K�z�q$p~:��[�X�n�
L��"�nl���k�ں�:�w�u-��S��%��~�n���p-5\�;p%^*�RuP�7!��TД�3A*����\/�T�z �V��}�lA[J���T��)`�}��"$�e�*;�ަ���بY��MU����"t�5V\3�=�ٴ0^S���L�m�Ұ�)X"��m�p�SL���&w7v���[��<p� �Fo��/F����U���3&h5��*5ĩ8�oBmN\��+W��NE#���E��2j����k�2t�F����fx0��8mE�3��_H���~��^V���y1;��Zfk���H�c�yw�a�%�4=@���:��ԟ�[�[�=ӸP�)�F�L��wA�����7���aݪqi��r�H�+��|:�b����l���2<�z���R��W���+.n쮬����%Ǎ�)^�\g���=���3����}��>�ٸ�M���x�2���w������4���F>G�
��������o��YրD��jt�f�"�r��q�}����I��:�����a�kʔ/�ȷ�~7�(1~*h1�����ݡ���8t\��cA�c��UB�W���(&S.bQ�P;�a�s���U��,6T��8�<*=��˃�pu8�
_as�O���v�d�SRB�](����{��I�V[vx�7߶~i�k�9���:93�/&pI\�����x�O�Ɨ�Ѵ5��%�Қ��'i>����v	�8�i�<oؤ@J˨~�̑�%�^��c��Fux�0�N�u�š.���>.uZ��v���b`3^�"Vr��2u�+����+f���E��|��6;�����k��.���U�at�����S	�����]p\���S�[��gXD&Wr�NQڛ�A��6c����0��Ge��:��d:]E�E�oifj��쥆�
��'�k��	�C���Ut�����%��t��op	��N����t���ήH^9���[hxO�ex�K�r���|���3�ڢ� R�ȼ�W`D4��Ħ u�^����۠dʜ��I�	�j��q�Yq�|��e�U�j=�v�n���u�=�y<�[^��'��7��mh4�ۘyv�n%{y���������1mf֤w�ڤ_Eu��\���˥��[�չ�_����&�W)���~�T	�F�֧gLS��SS!��4"i�������!���������4�}zt�kj�\% AE�ny kc*'c�i��#W�.�	��Uc��N�N�y�9��=�I���f�%a�s�5۩3	��Z��\f_T���]toY[]�o�kEo'࣪4\IVN\����#��7�cY�9�9�����t��e��w'��w���I����ƪ��Mx��Ǘ@h')�z����ء��,�GW49�x�.�U��a�9��"��g�{��������|/�h
�k�S{�9���!�RTvo����W\�sanD�P�����I5mFvy��td;��r�@od��H%��3#���tf���HM�iMD���wXԺ�w,�^��=��q��2�D\��}Q?z؁�Y5�ay]6=(Y���Fo�:��,pL�}��4'�W�B]uw7_t��c��Q�6y\�G���TV.�Feq��xp4'/`�3�`�жxR7�t�u'��W�t�.b�M�q� *�%��|y'e�J�Θ�# ��v��L�T������Qt�Vs�,�c7m�q�'��+�O�0���侾^8o���vUv�[���k(B�Mݓ{����7�G�-���!'�M|k�[�{�o�����}�㼺� �����\i�[7� _j�Y��{���>��钖iv�16�U̾[�ǻ��oo΀5�b���F�4lEN&|,/v�y�Ø�V�CO�4e������N�1�~RL�R�D4Jb�,�+(ɀ���9PĊ�8�H��H��c@n0��;#ZpwcN�J%\�N�Ӛ�`�y<��>��LhuF{c��X�� i+�]�^�B�~����&��/�uBi��a�,���ܺ��§B���~�PW@ʌP��t�b6>���!�I��0(k��h���/ �Yހd@�>_��^��>Y��,�eO6W�T
��dG�4��,b�V�,v$f�.�^U,M��8��6�>C�����G�X(��[H��X6x��vڇ�<��v;J� �E��T`�L]'�,�Q�d�ۼ9�G3'u�A\���K��Ҽl�߱x5�Г��vv�q��цW�!��~ݮo\�����!��⁎�
����̆��n�m���(�4]����k���a���د�ʝ��,�x1%e?z()��M����jC'oR�f ���I����Ʈ�z�x1^�G}q�.����G��ٗ��y�DM����u0�^J7�X�w��#K�(�z������a��cڢw�Ob�+�DG���Ő�s}Zl��q�cQ��h�UVg�1T[O�:\��A�E[c�{�ս[�&c�)��r�\Q��6�!^��
�,A��\UX�p�H\2��*��'�RW��#8��Ӕ̃X��\V��]�6˳�X(�:�q�[3���x&�GH�n���ҍ��[�*������<6a�b�֪SJo��0k]Ҥ�^�����FKt��QX��;���J����\�Ͼ]'�f��H����|E�,6�^=2��=h��:�mʑ���OX��l�b<�[�B&��n��B},�"k�(�^+�;LE�f��ll47Sɼ��������\Up��׭C��u�J];�r
�n�v0t�R鍌�CL�5�pSfy��Ihٿ�菨���Ͱ��d4�_S�N�����%g�yl�u�'9�k$�O';�ɤ�I��k2):���e��:oގ���V|��������H�B��������4�i�C����gP��Y�����e�Hg�0�JΡ�L�sY'Ry��2]Y"��[���_;�s���ߞ��vOY5����2��M���&�c��C�J��u�B}�1!�q!��|�:���&Y�C'��"���7Hu"��z��w������#|��V~�,z��v���9ńۡEw�8X"=�w
�z�u��);m��%���Q}�����p����[�\E��~�S������\��x��L�.d���{%�2�WuͲ��Gp\	�/LŎˏ8Ljݓ*���DG�ޕ<�8�9��x���s��"�N�i�L02o�Ra�l��2��<��*2d�g�'Y�k�	�C&��<I8ϓ��}a5��i1Û�Oo�~�צO0�h@�&3>�|�(>�rJ�	�x}�I�0��hx��0ͳ�����}�f�4��0��<d��5�	���DZ���@s���jm�F覕���e��4�Bx���z������;�'������	��O�T�]��L3m9lXL;>�O�c�"#s	�1:O}R�u�}���G��x��v}d6Ȱ�>~d�CF�O�I6��{�'�{�2��Ou��ԇ������C�;�hm�`y>�&�3F���F{誘��m���9gF8�=bI����|��>@��M��T',=N?0�'��u'ܤ�jq:�yI��Xi�9�Osx�C�CL}�V��,���v.�}ֺ��_���`�2q_�&�z��0ϒL8�2e�C���d۶xj��Xf{M��=��>z����0�q���<Hu��ۮ��W�+���R�>��]����`�;9��6Ͳx��5<� �2T��6�=a����2��i=��i8��4=dRq�HT�״�l'�ӌ8�a1{��z���<�pc:>5��s�Xq=d�s������̆�;�
�L��$�l0�+��dS����$�{�0d�Oa�0��'9C)
�B�m�Rc�.4Cω��9����<@�|É�C����6�2vwX�̆����8�o��X|�Y���,�N'1�q"�/؇�J����xb<�q��	գOt�ջ������w�ć�g�O<5O��:�i=�!�8�2xs]��$�;��'��ӝ�X|�^�x{�H�,�x�5_U\+��"���1{%F'�*��(k�J���;�r������b!�l�&ĮߓW����*�p��;V�.?l7�nO/*WY7q��{-�c�7M���4ҳ�'�h�q��o�7�9eqV7����)I���v9ĤA^o^�t���?fqUx%(˱m#̏���{��6c|�޽�wd�?	�bI�C��!���=@�C����6��%��q�d�f�Hu��39d�a��{�<z�=�ƲE�	�O��������ۍ�������t}����|\�x�6̗�>��a��1�u>d0�,8�a���Bi�s�:�i��C�=d���q�Roy��	�O>~�qoT����Uo���]{���{��ǀ��A����@�'9OK��c�:�a2�Y�!�M2���P�:�L�!�8�Vi'Y�C'�:�L��!q���Ʒ�΋����ޚ�;�E'N��+$�O';�ɧ�%Oy�I��́�Ra:�O��H|�l�,>Xi�CL���4�3L4�f�'�_�kOs�ߓ�xo��}�֎���a!Ӵ8�l��L��dY0o��%@�;�/�H��q&�u��gĆu6��H|�j�!=d�b���=d�=��VZ�~�n�T�8{�n�������=d�g���2�	��q"�����:Ȥ���I����ua0�>�$�
�`o�<`a�S��q�B|�6㳪S�]�۸���ҍ���=���}��+=|5I8�hd�2�N0�+'_P��ΤY5�'*Y1�w$���C��	�k��O�T����?g�{�o{�{�o~zk�Y
����0Cl����(i&��ٚN0���N��dP״�|�8���N:a<�8�Ԛ�Ӕ q���w�$>����Z�5�`�gn�+�GOu�9���G�{�����g�e�����&�z�;�ٶI��0�'����u����d8ȡ�l��	Rg�u��RO7p�Ěz�o��`�/����}�9�7s����P�F��{��ԇ��'�Hc�M!�e�i�{�l'�4�N��m�g��3�<x��f�ԋ'Sl�!�E{M�I_	�T����Dti�����gq2 �_���/8fF�I���t2c��k&u^�b�]�S��B�VU�ix�wash ���yv.�4��.�˲Y���5l�ל���\y���m���P�Y����T/W2I��]�t�j2�gyX!�w��D�#r�|g��{�� c��9�9��_²o6�l0�m'�s�<`u��ӻ�d8������d>C�8��]2O|��0gXM'��1�i�C��z�d�,>�IW��<�s�ϝ(�y��z0DD�����E&g���L;`u����4�|�����&�'~�g�O�My��d����"�����I����x}�x�J�k���	(�����=z����N���) m�Oy��'����8�ó��q�xs��8α��'��	��a�%f�x{����wy�'�yW�#ȟ���M���|~����	P塦N�d>3C���=��Cl31�a<d�՝gY�&�L��=d��w!�,<;��O��Y���`χrh��X���D}�ȤY6��cܒm�L���I<�2sVC��HzÉ�{`x�����`yl��C����n�u���\�@��<����w	�S�����#�����q���~̋&�{�"�d�l�/�	P6����(k��|é�&!�'�}l�!�8�:���`y��>����o��xV|�Ri�C��a�&��M��d��s�i:�r�R,�x���qI��ꄨO��'Sl&Xy��a�HOC5Hz�!�/�/�]��F��O{]�V_ݿ{�Dx�X���&��C&�q��+>g��q�Y2}�3Y'Y<��s&����9�I�N����pL�a''��x��>���	�Ы8����S���5�W˾�p��h���|ć�q�C�V|�a8��d�0�gT8ì��M�8�d�[�J�u�����"�7�L�́wC)
é�.c�����?�\�໬��D�Dp��V���=1a�8��f�q��=��g������L��~�N�I�vR,���$�C\�d���{�o�p=����k)*y�h˳C�Nm��.*�F�>:��Tʛ2���W�;9�C{TDթ�X��y����}�ͪ`���`+XF��[��c����
��v����N.��l-��n�0��Z,��QGCE��_k��P��d��VWR��G�z=�{�\�z�<ϼ���L0?s�C6�On1L��嵛Bz�X��:��:ϓG��4�&��x�q�Ru=B|ΤY8�&�0��L}���G�����|�^�������$P7�b'�&߹�>a\05�$0�!���b��'��b�L�g���q����t�q�Xz�t��b!B>��1�#�f+Pʑ6ܞ������2y哈�zy�d'�9��O�L3پ�O��2��w�!�z��!�>a2�;�L�3�u����>�	ċ�`����}��^��c�s��Ǻ}٫��^p�ē,:v�I���@�'��w��$:���9�O=�3'̇�5�bM�he������ON��6�3��3�xͰ3���0o?s���]��oy��y��d��wt',1i��"�'��'ݰ��8É�ONg�!�'{�Hq���y��6��g���|�Rq���̓�KἺ�3�r��/�N��h���<a>N�X�Ri:��6$Y8�MR`u�i�Y"���'XL|����Os�!�qn���<�{��m��q'{��>�~�.��)�t�K�N}����H�����'�>g���e�$�{�1�i�Cٛ2��'9a6�a�6�	����'L>�gY�O;�Cl����&o�1[���k0���[Y���#DG�-a�Jͤ��q�+%z�RN$X�CIē��l0����P<d����Chg���M'Xq8�z��z_�u���3�7|=�]���|��vw���&d�>̞3l'��`�>IYԞsX��,�x�1�q"��ݒ,���4��Y2�xÉ��($:�}�Ϻ���v����[�h����C����݁�8��y�w3��,<;��'��	�;�dRa:��l�E������K�wd�O����SL�)Ϗ�2W��~�WeI]X�QAB�S0�D����9dRWv�w|;�s雰Ϗl|��
���؂�������*��:4�|@OHz��Q���<�����z��	�Qr��.:���<��Z/��9�1�8��#WL�j-vS�.k���0EF�5�e��Gl�oO���G��)Q�q�L�,i�]p?-�%�P�z�'�e�*��W�%e{A˛�t+�ɔ�Q��ޡ��ǔdNV\H�t�㙓y��)_;J�Dt��:��oH]f}zX�+7���S�.��`t�L����]ۢ|���\x{�/��y��ͧ^Z3�9k۩�\��(v�G`�v^�N�É�nN����8�lA��ڥrC9�����@靅��r띔��k�&+@�u�\V�V5���;K:f�c���Y���e�1�4��Ԭ�0G򫡐�@���C������]�o2N��Qޯ����ӡ)Tn���y��2����X�g�nÚ����r��%<��9B���f R��΃���RQ��w:��[�c�&e����j�J9K��|��ע�]w�ٌ_r�l3�7W�|߹�K�˅��ѷ2>���]+nv^�Ћ�Qm��KU8�����'���hc[��A�$��T�-�0�Վ>�a9x/v��d��gLu	�x8�l�T���ʹ��Z������X��{y �r�:.75�]�
��q_r��w��h�0*삜�2����V:זE
�śI.;�ZVdP]y<)F/)����@n__i�/��#nu��[�s�z�"w���IH���>+��O�9�̟3�Gg_m+}"�I�r�4�Z@���O{�B͊�a_K����u-���/mk��XIpM,t~V�2s1��yʣLֽ����r]�t/[�;���@��Xt�$�����m�����eFc�o��y��8~}���C�m�73b
���ۮ��Am"�;6GU�ю��謅]��(�%�]�^S}UB_a��'��پ�8x�c��O\>��-@�X�6-U1�a��
�YË[R+np��
1.;�J�L8{����]�n���l>�1���3�u�9t�S,hI�;�8؇��4�@ɼ�1k�i>�y��+&+�iL��d*����x9���؆���E:�Խ����;�Ĳ�͘�Z����N�UňtvwR�w�L�S���^�4x��d�fu���p�\�*�l��< Yݹr[�h.C5��w��Am�pu�A(���;!gJ����/m����ۄ*�7�S]c�
t_*�m��lV5oq˳�.G�&��o��&���ҽ4^��i��ĝu+mG�[�C�zb�YU7Wp�4���HuK��@�uVhY˱�+���Eڢ*��L�D8���N���w�h윶����m@Ӯ������N�TI"��,���PTF"�������
�j+�A��5�1X���V��cim�UB�bTV����iDJ�R���Q�QE*�Ŵ[UQ��F�[J�AX��bȰX�l+V���b*(�T��F�+j�h����F�ш�QP��D�#j5V��%��*�TF�ZŨ�j����PD��DRѥjU�(�U�m�Kj�AF�E��DKmZ�T*Q�KcZV�KV�kQE"ŕ�eb�-X-VѶ��QE��QZª��%J1F��JX)F6ʨ���Em*(��V����`�����(�m���R�`��AE#hX�#��
F�,ej�D-��J�(�����"�bTQh�b��"*��"Kh,������(QZ%�Q��*
,Q��F-h�j�(�� 1X�����RTm��iQQ�)UQ��Z~��(��3.zgI����)��[��nn��PU��nT��iGM��rEՆu냚�R���EX;�3�7�ԇUfX���� }��QwGO����ό?c�3i�q��!l��f�:͡�����3��3i&Xy��2x��zƳ"ɇ�w�����ó���Ts���?T�ڿ��d}<R�^�]�2��>�|É�!�����6��l�!�8�5M2u��Xi���<��a�L�f�N��9��M'RN_q"��Xy�y��~�O�;�]|�u�~��5���>�;y�'�����	�b��u4�xg��8�P�VE��=OY0�$<=�������"Ƀ[�k$�Os��_t���Zu���oy��]Y"��Ěd�l��u6��H|��1:�d>d�>C��	�1!�q!��4�:��O�2�2��q�I���~�8za��5�W�|oϷ��"���{�0���|�Iud���M0��w��0�z\`�R'��*2d�b�L�=d�>M{a8�Hdՙg�'�}���wq����=����|�OJ�����"��37@�1�s�I�������M0��M��C�6�;�@�!�y;��d�d�4�a�%f���b��w����\��Ӟ�e�P�,��$�S�M!<��dRi�OP0��Lg�w�OR�qSL&�}ğ0��~��J�!���1L&{�k~w|+��^�Wf��7���O���q��+4�j�|Ȱ�:��:��t�'ܤ�M� u�]�{;�I���k��'��{��I�!��	�6�05�{���d��}�>��s��{�^OY3q:s���/���O�xȤ�m��8�a�q�	Rp�Τ����� q�����Hu�������!�:�3��{��y�w߇�g�����4�zù�$��3,�G���L=O�q�i&��'����E�n���u�}��d��g|�	�ɻ�8�d�w���W��-7�sGC�鏕��NjZ>��t���"�A[&*�)'S��b�Q��٢�՝�aT�ghv�[��,�Ug#bɊ۫.��~������������36Ko�ܩ	�>����5��ľ\����ɷD֒պ��
{7�����k�z����k�?	����?/{��d<��rf�<C�<� �2T�y��OXq=��!���I�s�Y4�H{��)8�$*�h����W�j�V��kz��1���zV&XLvN��|�d��|��8���Cl�uJ��J�$�w���%fn��N2(�a��I�|w�Y;��2s�<��}�c����ݖ��Mvz�l����b"$z>Na�D���|�i�CI��8βy�b2gP�/w�|�0��+2Vm&�y�E'���	8�L��!���0<��S? ��@K�.����<��zG��6�!��Ć�ɋ�l'�j�3�u��zj���f�<滙�I�w?fO�'��
��J����E�d�ß�>�?�q���.���Z���c��}��,��b$�Cٚ�=a�����g\&К`j��8�2u3St�Xi���l�,5��2x��eQ����.~Ò�^J�N<�"0{�y�>�dRq�y/�	P6����XL���>a����3E��&�z�Bi�}gYX-����H,�u'�}}2e�騯�;R�>�:VV��=C�s3�z��9}�Nf���pL�a����{��l|�Sl&Xh�q0�i��Ϙ��3�=5dY��&��N��3����>�ۏ]p�q�5�t=a�J�!�`q�I����N��;�ɧ�%ONgi's`y���@���q��>G�u�	���:��!�0L�4�i����oyvn�G.�W�G�{ޡc�,�C?P�2W	2�:Ȳcs8a*��I}�E���4��Xs8�$0é���H|��Y�L���.5�s�$�����v�U/S������=�C>XM0��MS,��m�S��t���H�u0�����J��;�E3]�d���g�wi�L02o�Xa�^w[ˉ�!c���jc5�K���W1��w�_P�Y,6�6,��Wms��SAsW|rs�l\���꘾W�Q��w�n���!w �8�
Y'��n�۠�w�&����M-sG����^՛��e�2�<�t0��7h���N������*`���k�o`q	���1P���'�)8��J�_�'u�g�'|����MYԋ&�d�@�&4s��H�d�{^����۳�h�Uq��و�����,�;'�*a���Y
��v�d>N�P�'��	:��J�^j��"�=�S�I�6����'ذ:���9�""�p�ߣtA�4_��c�����ćy��?0�g��$��!������=g��l�$�;�i�,���u����j�q�C�q���>N�}�I��y�a�'q������Oj�2����	�C�6�Ϲ��z����3���1�&��2������0�;ha�d��癇̞<Ha��N���!�E*�r���"
izT�_���0W�_p�>Մ����8�I�Y2��S��$6���y��6�|�;`q�*<�d�0�9;�Y�I�瘆Y4�!ﹽz��}��=]�޻��R,��É
��=�{��OS�8�a0�7`u��z�\�p���=�_���mS���!r���+F�/H������{�c�[S��(���N�֒5�����>��`��xF�H�m�f����7���x~+|����~���J������y����V8d�c����mǛ��m�!f^O���$7�Zqe�Z�����ck�������p^��l�r�.�w�O`������O�-�g^����q���_SZ�aF��c��w��|��L½��j�
���u�Nn}k.���.����H8o0��Tی��an���Y�}V��oK쉹b�I7;C9��U��Vsso��@��F�1����=�^�M���Z*���}��k��x�`���#�~>�{��v��P���;��vx;����9�w�I�n�`�ӓ8���|� ^>���݋�n3�3�׃k�9�T��	����{�='a��c�ݺ�Zį{'D��}Ux��\=iY���Q�9�^�#"���Bw��=��n���S<�@��sYEK�s3�9.�YR���@��W�MD*�x7o\�\<��\�݌d?7��v_@�؆G`�O)�{&�iy����3o;i�}��\�-����z����sj!���P����:�pr�xf[8��X�+5�n*Wp[��^w�;���Jי98�y��c��2.,�y����k����jn?B�C����7�/'y�wnչ��m^���TR��J7�8���΃|�^���������}�/vRW���ك�U}Κ���4������Gv��-&v9���*�HX
�0�̓c]3�n���cҽ��+H��tK�0b�W��)C�J���S�������<��UW������-����-��}G7B�ƕ�[��Ci�w����/�#�h��Ğ^If.��{�vKͭ�$�����έ�Qj����{�����o�Þ����SDO��W�V96�&m+���U�Imt�<ٗ�~���p�����M,����WC3�ƺ�3}�G���N+~!Ew"��k�ɶ���v��V#�x�_E{N,��kg65�K�CC3In����q���j��Ʀ���Z{׭�*���FN¶�$=�f����)tv͹�e�j���J�j�h\ݏt md�̫���GӖ�G�OU	$�Z��1O�1lf=��viHy	�9
��=J�~%�ori���ej�y#�>��j,3��B�&�i�
0LLTᖷO���gsc#xWK�Ѽ��]j\t�}N�S^�W��}���e]x�:�r�_=y�Fh��\5ȋ��Es�V�l�Vx�s��N�E'5�ͧu�p���W��O�*�
C�nx��&g�y�M��¸ :���b�U8�t��B��e���OD��U�G��� ����[<,RQ5��9��U�c�D}�zB��k�P�6])�*%jQ�9�+y��bӦ�-o5���B�a�f(�Yzd�"v��\�I��{�w�ԧr!���諭OmI�I��H��:}����eF�Ƃ9�S/d�X�Tl�.w�����������t5�{�~{շ�e{z���$�8����m��O����u9�ɓK+.�m�lwN¬�5�Z5��+��ͼu����}�Fm�~͸}ے�eCY{����f;�%�_(���a�ɫ�Ά�d�����)�a>�M���SDB�LjM�J�p�C۵���Ml��N6r����F�#86��9�n+�u/*�5�H�f�Ҫ1.�F$Vv��~�=mNE���S������O���Quxognrё�����a[�&ۙ�+��5<�W���΅�MyT�#����a�ݏ=��u8(d%њue�ŭ�E�u��X�y⮏T6/"~\��<�n������.��x.�:%��h�W�4+���P����[r��}��J��z����v�D��=p9B��y��c9�n(.
2ut���,���7��P��\lX��e���˺3���LsD/�(��)O:�'
=W��p��$�7�&�D�FpŌ�ß[Ϸ��m]>� ��~��ǿ��|�|׽�~����~�t�Ù�h�9�2R�t�}58��'��Ms���*���ڃ��}ê��f�^S�k�2Z�v�}4q�)��]�3P.([��O�uW�dζ���D�ؘȯs�4���u��˂�?o���oxS�b�4��v��z�|"�������Q�:�UCذ5k��r/7B8�w6Gex�Z�Z�k�T�3�n$+P6r��s�	&���{�>�6���$���.�����++�/3:b�Y���Z�~����ݧ�vݝ|Ml#�%��Ļ^�/�:���~>̒׫�Q�̉~�Nv=��Ŵ�sҷeX}�l�J���p�"�dM���.�}zD?&�a-F�����|մ����̼'�ج�q��Oj�ҍ��p��_8�I�A[��}P�.�-����)ӥ.p���Ų,炑F�[35�>��wjJ�bj'a�Xk�t<�6�)�[��c�F)��$e�3=з]N��ٻs�����U�U`�kx���4��aX�d���i��j�%:���E����������xi���{��X��v��lOG��b�kbfҺ=1�ZH��m�k����ʊt�,�J6S�F�7�u�`n���\�WO��ck3U��f22���%�p�q^���S��ߒ�7�"M���C9��r�o��=� �W=�OV�ݥ�Qu�Nʽ��mK�:0���L%��Y^/�n��o�<����j"�u�쁝��^>��|�s�9�v�AU	����zX�;L��ڦ"%���]�nb�T\c���u��	���b�㼩v{��UyC��zD==�r^QŕX�]�'#��a�k��5v��
�f\�w�������_�,�v�	�*�����'�'}���
�
�"�Yx���2���c"��g��M�S�|Wo���y�L�orUڡ��U{�rc��ԅ�M@�
�y9�w���mC#3n%X���7*˦��u9���~đ���sv��} �Y[ʳvg�HoqN�5�"�[t����s�z���
��xN���}�m,�j��=SN���SoZY:��0g{%5G���<=���U˒@�.�|�[���:�<�ZAa(��QU��{ޏG�kv�Q�E�aO��eF�cA�N��<�q�vj5�7H��:�ԣn�&r��/�7]<���^�q��[����w^��w���k���	������u��C���֡!�1J5���U{m�V��j˷�Sɜ�j���t�̺�L.ܴg�I��7�^E򉴙�v�2�}�@R_��|_�f��Lt���}Բ)�&�Wec�kfm+���U�/��gm��7�Z���.a���ᣛ`0�ٝY'�D��qU�,�s���p3R��2�u���晆���,���jp�\�ϻ9�Ա~��c�Mx�[z��gVƧwڲ�55�;\���[ﻆ�s��e��Q`��?z!r�Ys���Լ�X��ܥ]5
];G ��w����{�qUC}�U^Ƒ��>�K��׷1O�.1Lf=�@x6Ĩ>��:<ϫ��*�E�]������!��=��K=��!�����{���%P�Rtuj}!�t�k'<� f%2�kE��jZ���]]h�8X��˺�������qv>��G�,�cyf��=[,JL��*�-	��j�R=WYf������V5Y͞��׹߼�C�s%+������*k��vMZa��-��,\�y���S̾��!�:Q�ү�Sp�v"��8������n���ͽ��"s�lM�#<���q����<y�}`��C#r�ⷽ�R�ifhq�GS��.Ҩ�ʖfq>��׀�s�y���_:?LL�m���3��Ľ/�zT�>���ȣ4��sy���A��v��u�[��ک�=>������Q���lqx�}��K��_M�
�x�q*��>�Z���{��em�nW�A��u�)=cbU�Ԏ��[��3Z본�?��cᵽ�{�|��lõ���$#��[:�� I���3UǛå���K=ۮ��s��m�nDSDL֘.�T�3	wJS3������f�������F�m*S�� '�E��m#���Ն<IVe�Ql�0��J�ʈ�ʵ`Ӷ��&�,QpB'˥,���su+��Y��K�h>9�v���0v�r��Z:v\��sт���V$��ӨS�6��\�C�q��ʑen�x�I��ͷGN#l��gOUn\��ןJ�(Q�xZ�K_ڷ̫TU�[���Cq#h�uԗ<ua�{��h��Ma���n�X�9^���O�� -]&�"챼�\g�;�e���*�+��QJ�TM�}�v����m@(�zn�Xr]��|��%uJ��d���K�@��j!q�K�ci鸻pԮ�G�wZ�ݪ�-�Qң}�-����2�k�3��I^�P��,E�q��_[Ca��x��q�{M�6K�Iz:׽LR����,�ܻ�=`5�}���)�3�.�/2���=���M��g)���*Q�|�޴�}ynS��`u�,t�g7-:����̡S���M��<)�����.gO�⚎ⳢW#�p��খ�j�����SRf.M�0r��o%�zd��㼻���Ц�X��q�T�Gsф.=|�]��n�֗2\g�S��պ;�kޤU#z�|^.7�qQ��:����������4_P�Ss\��*�=W��l�}9_�x7P��N�sH�ǐ��y��ƽ��f���[�x����G�]��\��g�O�v$��bL*ÝP�m���6*0wG,w��vT�a�9�kfO�u}k�۝�Pݼ!�諭;�]0{���z��E0K3�8����Y��7,��\�W�O���f/n)��k���)���V�# �$�.Ө��r�*�w+Ev�"hw[w%�|$KVg'M�7�8���h�����	�1V�0�띸Z�S����I�ywg��&�K�?7���{�������=S
Lz��}&����2�⿻J��,��C��P�4�]m�Txiv �-w�����nTÍdhPU�f{��6���Ov%d]N�r���Pυ���כ�o�fE~K�2n5�&������kLrt�Ʀ9�O5����(�Q�kcʻK��������6nI��e��t�j��]���׺1"KNx�.�4L������e�Ob*��ܳQ4a�r��w�����ţ��� I��7�o�m3d:A}\v�������e�$��Rh��������a\��\�v��ã]J��w�p?`��2T�%�q��"U����X��8�lG/q��M���
�IB�^�w�0+<����=�����24�v`!�B��CY-^���3r��ɾL�!��[A%He�	�շ��#r�i��
���LO1�}¤/��\����R�k=E�h��m�	o1��e.kw"���t�#�]{5Q����y�6���Zڛ��3�+������K�nO��{��
�UTV�E+m�mEE�Ս�Q+(ȌAJ�KEA�iX��iD12ڨ��V�Z�ckH��2�J5�҈��--B��VQDc"(2�UZ��ʣ����K�-��QJ�X��#+T�
����[+F�[FT�"��҈�����Ԣ[X�U�`��Z,[J0QA-�����c�T`�Q��F�X�ZU����
ьF"KlX�"��E�+�F",X�ŊQ
"����A��*Z"���V*�D�U����DVڑ�l���QEQT�JƵ��j �DA��b�e)R����Ѷֵ
�2��F�,`��5*��V�֥c��"��m�ԱAEDU���b�cV6Ѩ���[�Z1Ub�KE��EDc
4AX�*��l�  ��aS�o*_^.Cb�P�^=���Q����'�%������@h��^�hi)q�����ι���<}\!�;���}�v��Ώ_�G���$u.�����5:y���V�h��0��Z�۽�><��p/vh�jܛN⫂��O/٫)cR��e\؝�Tn>�W�ζ����g$�n�XtI��4��C9�˒�|zc��*��٫��R�m5޷�>�/a���"K8v��uaF�Įظŏ7��M5r.Q�eGut�7!8��}ʓ�s8��4�JV�O��3��iu2)�D����J̻]p-��>�h8�a�s�#nx��;P�|�#4Zlts�2�Z�nc�����vLƦ8�v�11q���yMѦg���#�N픫�8�~�)���{sy#��o�C3���O�����|��h�ƽ]��M����m";(�Q��d���T�K�x�q�U=��j��OH�ً�����e���k/v]��Pm���`z2��fIEg\�P�l�/A��gJ��_�x�����H��@�P��v&��5������n�<��k���;e�z��-��*j�ͮz1���7{l�Z�}�(Cy�K�>~�J��U\I%`nڱ,�����;ZчN��������UUWit�+���	�����b��Ot�{�^���ӱ/+n"]��Eu�]T�^�P3���Ԋ�pվ�n��]��eX}�l�MyV�#�����!Г��잖"2��сN��z�{�T��[��}�-0��)���<3Caä�3�nM����_(���܊�W>z����6��Nf��s97:��	��z��j"���U#z�C|��n&��-�!�.֥n��T�ۃ�g�;��S�����)fʭ�]�X�͎�����,�J��I+d�8m��Һ!���ߒс����,�v��]�揧J-�-��v`ٔ��Q�駐_[�u�H��Q���ۋT�J4���|��Fm(�x�|5c���W;�3��������Ha�z67�s��Nu���ꋌS�μ	�TDw��O�_��a*J�wn=	�j�F�c߄l�
b�s,%�H�7����_pW}�4��>�9��I���5�#��i�8�I�V��8ֳ5�I����(�WX�S�
X����agB`�	�-��{�ĝ�F9C+JGi�:�)�/�U�i989m�W�}�{ވ�9��U�w���h_t�ŕ5�/S�&cyFs'���C7튾<��%X2�.�����l���Һ���\���"�SB�=�������+z
��}���6���^8��D[Ɍ�Tm�#y�J�e�;*��2��q⍤����j:��^�g��^!&{�lݱS6q%��hmh����el�h#)��_%~��N��c�K7�"�g�$A(ޤ�����z�8����ݾ��ܛ�٦�Z9���<q47{�oה�k�B�P}|�c^�ⒿB�{p�Rg�����zi�d�tՏM�[��=~���3װ�m_�㺲]�I��X^5��.;(�zs���������R�Z�2���qIm��ZԨ4絩���Z�p%���>N����6�L�R���}�u�Fo��7��Z�V��pSJ����g�Y�i�rf��!7�nrlݤ9ݬ�u�)�W�Wͮ��){\0�\��-��dA���n:C}�]#���p��w��8F{���\��_i͒�-*dm����	�����;VW!�×
��mN�����G��Դ�>�?x�U��/5:y�|��Zѡ��	Qk��;��)����m�C�K���#$�d��`}���r�_�N���~KT��kLj
'��A�K���m��ue�ŭ��U/$j����)��R��`S�K�eggIN/%a�6����h�ڰq��x=�=�����5 )���1a�:VV�i�u���R=�y�ڙ�����]t��vS��
������Z�TC�C�����!t�׎j:d��@3���{^�ő����P���ޔ�ծ�r�I��Fy���F&.���P/�-sG�؉�����Λ�V�/rrk�T�k�f!K2���la�y�=��̹G�P���lMߪN��..�J�����qyZ�B(�u���,�ۤ�t���ɕ�w`�M���Օ�м���W�����r�c��l�5�-ލ��D-��W�yw���7�ԝ4yP�`s���𾽜�����$�:
�N�M�2R��W4�&a�=u�z(�=��fr��9;����[G�w��3p��eg
sy�h����,��V\k�t�S���=�\����R��"~�����ZR㎫}#oѾ��Բ�[���lV	��9�sV�q�b��B�ķ�n��H�o��ێN�-�ۑ+vU��,9�Q+i���nl���s�����gf��^I ���ϩ6��)�'�u��e�ʜT0�«�i�ޮy�����򐟕�
�i��y>���h	�dz�6�r6�@9VV�q��y�r n8�)
��9ݫ�Cո���fȬlq���eh�_Ӡ\��}1�Y�.������Ͻ}�L�݆����'�v���W�����{��c����!|�IB���.���V���C/��?h}=�G�R��I��1���C���T�]J��9�Q�;�5���=���[�&	U霼%X�ݐ�ӓ8�p������k�{7��oNb3��Ps�i�ar��KP�r%n���CI������W\�L^���f���E�D��l�A���Ov,<h�jk��W��@���֫��5Y]��kǀ̋H�����:�.
����|�,�zn��+y&gj����H�K%G��H�z�(��7���_�Lfx���6��x�Ǥ  =���s޸����YW��\��7f�}�g�c�.11�Q���$� �aV����B:�9A��x�4��-�s����(I��r*�(?u�a� �'v0���:-@��2;(�^��&�F���1=�_+�K���Ʃ_7���zǞ�<�k�:%�����5;R�NTa�w�/�(��Ʊ�z��6���k�n���t�K� �˳�y��-*[
�h&�X�ooW��վ����[�b��F����7q��Q+�zw�����g?M��gA�_(�լ�$�!M<��[M�~�$1yu���+��yo{����^N[�S��7	V>�Q6�5�*����O�]��(t�_T����=�������+N��u8�fҿQ��i#^�N
X�nNn+�׎;B��;�����ᣪ- x�7P�8��M��+��=�k� [�W���P��g���ɚ/e.e�����?�v
�yT���Yͬ��|��tT�(A[�5��G������ǔk`�A�q�xԵ��]�Wx�*�Z��z�"��-�wlb������O'D�a6�D	��z�2�諭��y�z�ψٵ��������oF�o�t�{ғ+��u��}4-�FMlt�_5kf<�>\�`&l�}m^Թ�R�O��>�]�5�nrg���n͸��s�y>��:ԫ����r
NKyW(����e���d��#�]5�^�`.L�=��l���̰:W��v�WZ,���r�&o,��{O�2T��+zX�l��r��֕��N�`�F�F�z⦝�BC�VN�p����X�P}p��l�ʉ�u�\�=-qR���o�rB�AOx{����1M�sk���V�-����u�X��q�:��J�s*7��f!'����c����s=���NKf��K#���n�ݢ��nt��+4�{�I�N�{�Q���e-ˤ�]�IJu��v=��"�d[�Q�UG�۷��w��ݾ	��0�>�z���o�]��$��W��s���Z��C�}��.���d��zv�f��d�n��OY�S+\8A~�]�h�t�-���se�n�����_k	��л��W�0����) ���8q�9U%�јL}�8�n�V]��_���)f 5���g�P�?�e�}t�a��Eښ�t��U��M�nD��W-�g�I��n;�2\��E��3KmѼ�ӂ��� ���n��>�M�����T�o~�U���@�|}�1�Z����o[a�@&�V2N�zp3^�>;�@���#jVF�f�s1=��F���$���{N���U�,��N��ok��F�P�BA�ݞ���:�PK�мhddK�xk��a����{uNJ졩�j�X�ӝ���P7.&��'���̝�P�n]u�[���Q�F�}��S�8��!Il|�s�W����8m�c��?�
8��7��z;x�rv�6�_�-OD���S���9�h�9��)Xu2��X]��w�v�k{^�v^(�~�PlRv�0{a�:Q�ҵ%5�N^[�yeR6��K�}��u�XT+�Y��=!T�n��S(t۫��� 0���e�S����u>�4���pj�i��K4��K��0sA�9 Y1����O����)c.���J�����g_�vm�xڽ����X��֡�N]}un����8=���&2+��t_o��}N��3��I](�����܋Y94�\�F�FaK)1���Nމ�ؚ���U\�����q.�Tbs:���qm�vL{�5J[ymל9����)#*�����y[~�c+ؠ��QuW�-�Y�;�U��y���t�y9��&��f#�$���?G�`
�h�o*_�3A�`n&�i-���mӋiv�Jݕq��x�J�W���*�i����q��5kQ�iW���s�M���h��֘.����UO��
����x77蚇�:��ZH׭�^S��'�F���s������fG�%cxkD���K˓iH��V���jo7��}��u1A�Y��SC���h5/n��L�+O^Cq_��L߲���Ps��DI�9#wG�z��e.�Ia��>�)����¤��I�%�\`�x�����MV����t�]B6p��Z7,@]�hȻ�;"9��.\B���"����l�H�G��#�9��O�M\x����媪�2�<3/0=r���&4-1�uFn�Ga�&�h�d��G��-hN'mj���V���ߒ;}ue�b�ܷ�=�vv��;��;��5'����W=9
];G ��7��O�-��s�o���'WCa�;/M�m�o�z*
7���;���3���sJd�~t�}"Ѧٺ��{E�L���ٷV����x6���èNq��sQ�%�{���Ee�:���Ձ�Q<�;�j �ʉ�yx�[t�B����Ͻ��zm��:�@tix���sc�D�{�;��X�V[7���xz��9^��*M��Q�]�}�q�闖�����s���9���*�֧94�K͋��$'RU�s�%�����R_Z�����q�<����w���1rSȌ�V�+Zg�9=4u��,�}����ݧ�S̜zM8G�K�ٞ��a��[�W=֧�X��s�{�u���V����iv��+��ʈsъ]��+��Y/rb癠��n�]��c��[�F�����\y:���]٢���Av��ӧ��/S�ֲ�i�4���{�����Ջ�G>"�;����.x-0�Z�!(㄂�{�����Cr��ϼ��컿K�U����*o����q��N-s$�3c�jٷ*�� P���B��H��l8
K�L_ϞN��X���<�H�*�Tf��Usi-�ePKhm�y�	+��pA^��ƏKL�Oys���S�F�^V�b�DE�3,����U����:��D��O~2��uAVcx�n��5]s5��`)�y�{0���힐��Nd��1���Vh�#�,�Oz=b�C)�Փ2�6�aے�0�W�C�2�M�r����ս��H�N�~]%Q�~'2h�{��2E�ݿ��v�؞�\��(���o�|�;���Y;��e�8��j-�� '
�޾x8x\���c���v���E���G�y� =�}3@���1L͉�:	v'�i�3p@�+귡��-Ξ? go�gs4b��D��$���m� ����@d[�`ok�|����X��v,�es��V"��Gp�ɫ��<�l6�X��U�U5�[r�~yn�7b�V���2[p6�_*�]�8[���ὀ=7��.��3U�����yF�V7���4r}��{���՞��bYj��AH�E�hØ����v��o ;"�k�4RǮ!������k��7
o���b�[��/��5,(����Q��<M��o���|VZ^��캺�������D�W�g�ݳ:�g.V�\NKh�}ׄ�]����Cl�����SP�kWL� Z�b[���&<"����8 �:BP�OEx�k/w_j�8K��V>���	Ym����ձ��p>%�\]r�U ڜ�9�O	 6%�Q7c���.�4��A�n�ua���A����%�Fn���#�U���u��b�»�U����;h�T+l5d�8����aV�j�L��-9�ґN��&����.��
�$�n��;�ڼ�}&hC�&.��#ap�d���'�LGI{�a��\�(��v�7�QT.���WD�/���E��H�}��o�$�">�|)����Y���<.{Q��N�l0��|xc:T�pj�{��6`K��#p�J�c�@�R���Y1�P/��5v\�"Kl��%�x_��r�h�&Qb��j�i��C#u��o�'��"k��}�wzv=�侌�8�o}���i^��-8�NpƁ-Y@�����f��0vQ9�#�/M۞���SN��H�3'o.�	hlM$��9�|��u��s��iOW���1�_�t��{;�-��2�X;z_cJ�h��~�����|��^Q(p�C0^!B`�=3;�,́�l<��$�]t�mm�ckR��0�i�q�SGeaXF���D,����j�-e�J#-UE-��k+�UF5P[eTm�ª�Z��Qc#��F[EYZ��Ab�*(�*�cb��E���2�ȋ�խ���U��Q�*�"�֫[
��`�X�cX���l� �dE���մTQH����b��[KH�A`�Z6�H��Q`�Fұ�ʕ"��#"�1�l�U��E�E���Ċ�A-,UTU�"�Qb��A"��*���6���mUDH��)�EX�lAVE�6�1�E"�TQU�,X���,U��BڬUQX�1+Z�1TQTUUD+PFҪ�"�Q����TQ*-iF0��*
�TE"
��*�V �YmDQ��EUb�QTDUQE[J"�TEX�*�Qm*�b�X�"*�"�,A�"���QUKJ*���X��MY�D��!����F�����)C͔�Jb�ޑ	6�qU�۲�[:��x�V�]1�NY]���*� }6~�b��_���E��jTc����Y�IR�yp���i��˝`�so_��3�\�G�I���sW�J��_(�I�A[�^ �oM��������YYn!7�K)�!r���Yn��&m)I�.��9�f�}���'��C�;n!�j��W��GTZ@*-D�kጮDd�ܗ�,o�<fi"M�C����\>K/5e,}5�'��~J��E43�ʩ�Գ���ݟ#�9�wӁ+p5;�[�U��];�O`�����X��z����*�
��ވ\�R/��[ڋ�s�y��:IW;s8����:��O��}��t�x�I� �t��^���޸�1��ƼA9�TO!�NزLO8sss7;����׹�ÜsNd�~��o��^F�j^iY��$=I������_V	$3�8<6zU��4����z��>�r��b��ێ�����$N��X=XS/HX#&Tly��ۯ zn6�/<v��(SbRen)wZL�A;�Z�qM�|���eut�{(˞�f����x�W��^�g���U�l0�W�k	��͙K�[��\eљ]�P��}P�n��^�7)���G�}�r�s�Lbc"��3��������0bv�0�3Hͩ\c��jKSY^Ҳ���R��N5����D��9���,��N{^���{���f�~�[�W�헍v������6�E]9��g:5�D��J~GzjemĬ^�޺�:�+zݾ�kvW�5�}�:y��xɼ�f﫽!~�|��o�k�)u��o��P�wV�j�`]�N�jW��/�I%��£u�{��[�J��`ݰ=.o��J���Ybw/��ψ�.w<�s�M��-��u��2���⸙��q�B�!(�w�Τ�e����̭��VI�oN3^���ܐ�{��}���V�(����-����^�)dܻ�]�q�,�f��N���F�%>��u"�������p(plT#�.M���0Wexjwگ�cSNv�5+W��3뼸��� �N�f1���CBh���e�RQcy��_M��;�W:���|<��p�M�W��g�bf1��Ǒw��~�ܡW�y����V��G[zuY��`�B�g�X����0���&e��������q��ܬAoN��/��XY��qa�&�q�zb����y��@w�w6�t��GF�S����/a��J3��� �mZ�<�~�*�}w�sb�X��gk��w(�c��9Pi�h\9Q2R������*k��^77�7��m5Y7o�JL�.A�s�����L���y�۽G#1����0˼���z4�W��Eҩ�/��{�v�.11����E�_�,��|��8����lZɌ�U�r���)fRq1��Iu��P�17X����˪���m"2��*�V'9:�;�q��di1V���\˼T7���N{����fqF�~X����U[��U��^�}~�b����9�W{�\�2�so�:���3�5�U�����t�^K�up���B���I�OnwV���Jݕ~����sƢV�wXͧZ1NSWtM]����(v%mn��@\�����]_/��]�y�.�@���!��fܮ��k�����]��j=u�=�P&�R��SI*a��� ˶�[��D�Z�C�8�H^�c��w=z���n�8;N`;�7{��nDG:�n�펏{�.U7iT�x��$�
��rm�nE4D�]jGEH�'��m핃��gs�$��^ڼ��l�jH����\��у{y.�X��o�����[�0�"���R��JGw��Uz�Yq��C��&:��Y����USR񬮧���1��-y �g�n�^Ӌ.$�wR�LO��_��]2_�*�Ҍ��Yi��ӝ��ƇQo�T>�Ti՗��yrE�$Ӻ�
��F=�-���ur��
�-��b�c��9�8��A-�ޞv�<�z���Ǵ*O#���9�w�9�S%+��cۜ�
�����}S�/�o���ҧ�Ix�`�Q��aס9�.�t�o�Z��S�/K�ٚ�%J}��/(�YW�����vn����������(�Rq�/uǫ{��$���MeS�`~>�^w�M��s���`OYwZ�t���v*�-5)�K��Q�ٱ��WF4ǽ��O`ǽڱ0FZ��{�c$�1�.�c9A��0�|`h�m^`�D�]��VJ]��n��!��4H��Gl=�7#R�v�ڋiF��r��w`z�_��#>3�*�rH���ĝ1iI6:�-��8i��&0ּy�j�ͨdw��;���z�
�|�T˰���+b���2��7vs^�8���si����'��o	ܜ�]hh���p~&D���+�+ic�O0�{�Q����=ӱ�*����#Y�����֜�Y�m�ש��L��qɖ2wk�su����u٤]������O�˗;,�=�b����Y��2�5RSMf m:A��9�zo�����̼Rmo��*�.}|�m$j9��.ba�uU��zq���;�j��Բ)�&��V[��q3i\Q�N�v�HR��k
��x�k��+~O��گ��h�HŨ��*4��+�޼�]�Ϊ��ŕ�]��j���M�M���2��ֳE&�YWu��8�0	����6�J�s�Gm�Ι����cj\�х/'�@-ع\�����p�ъk�pxXzv3����Y
�|f��U�R��,&�)���κ��0Iṋ��9�mAv�oNou��k�pcvș=�����7ښ���H}/al�	��{ZS\\�Gȩ�6�^�k '�.2�
\�gr���d�@����&7���o5�Oޒ.;��	mz�<���s�s�3��B\⪩�7I�V2��n���`�K�������)��g^���W{q|*���OK�Ѯ��nq�GL����};⼲�r^����O���W���9f4nA~j���ȧm׏P} �@o�μ�M+��ue���f���	!�k�\�����z'�0����^w�0��U�z���(���%��֑��O�&\���gU���f<<�0�X�s�;�p��ۉV2�9�N��ⲽ���(�Rw^I�9u�H؛�p��ׯ���/.�$M6{f�VV�K�Պ�|5pVߛ��X��\ᵧ���Jm�_�nt�oӷS��b*ڱ��U��ul����R�J�yF���>�["�Q���ɪ��iy�� %�~���T�5��U�"�Y41+Y�E#n�r�������h���f���Ə��� ���<G����
�w\���َ��i�{z�8�'�Y����Y�AI��n!ͻ]|���	�����P�+��CZ�����hi�NK2f��w]m�5Y���!aiIw��n:p�l3�ޚi ���}P�}K)�$.�zee��V6۷`�[�f�p,�������.�yN"�L_uZH�����'po_�;rBh�)��P�[(��{�	��OWv��ܹ7�덮��ifjjl�{�~ZY�y���"���8g�<׾�����2�Մ;K��* �ۖo;�(�߮М�κ�v�:f�5�ӽاw5�z]�.а�42�ܺ��nv�C�{wHÈ���{��mҚ�.��9T7б�Kd<xbrb�׈���8�E@���^�����;`�Cz厕�/	T�JW��S�Y��M$"S���j�Y9w�ꑛl:���9�^Nr+���t�j�����%\(�B�[?����D��^=��vL����9��j"}����<$C,d�R�.���ʳt#����z+W�̫�9ʍP̦
Nz��!)R>?��a�t�֦\U�n��9����pȮ�d�9�2�"C��ɨtLP�;si������W
������!�tJ�Z4�rN�E�\B_|��%m>q�<���yf����F�f����q}S��J�kN%wW�5��u�C��*х�x:=�5��y�ee�gd���/�\��&3jcr�1@����Ʃ�<_������NGy�I��Z�(aVz�`��r�}���Y��05.;xv3�r��S�������=ʩ�����[U�q��2.5�L��2�
�����S��e��5N�Gll�t����Oi�ҹC�P��g���e	��������z��t�WP<��������Ͱ*#QV��F����:RSq*l1����1�)ʒU��8'�+}����Ӕ́J��!�\��$��R"b�3�J��)�U:9d�kXB��y�y�b}C�y�f������{κ���Ҳ��;%uƆ�}1B��G�ٚ9�]QނX�V���r���෶�@�)FLBU������^s+��Y��x&��� j���yF�|Dl�GB�ֺ�Ɖ�L,'�����+W���BaYؐv�̜�}C3ǘ�<_n�~��=P_��1�e�xs��P��┺��� 
)�qh�ڠ�a��Vi���
�9��1�h����)ւ��x�R�<�C�X��CDm����5z�ޢ �M"�;��f�έ��ŲZ+�I]=�^���e���^3]�e�Hk]6��0u�2���I�T�����"�X1:�{s�^X�Y��$���IH3���:=YEIz��O�O�H�K��ܘ'��V���69QG�S��J�H%�a>G���'���
��e	�⍲�$U����t����*�9��=�+]��޷g�����"��H`g�cW��Ŏ�V�8<��y�%Z�:��e�*��㮹y�D����s�59����C�p�Gu���r춲X�^��ze��mf��W�\���T�sk�&k�`��
X7�r�Ę��{�8B��y�$����u���i�Ռ�H�5z
e��P��V�岩_ޔ��W�Di����ƶ{�����E�p�C����s�K�^�,�+L\	g�eX���L��杜~�b������s&ǹJW��;>�z����j�,>�U5.�+����T��<C/�|�� �㸒����`���W=�ޚ|��Yٿ[�U�D
��qH��Ua�ً�!5�y]�V��ڽs=l�3����r�y���J����kQ�Q�
�d1Wʀ�P��Ӛ�X��0tB�kQ�M^��ޛ)N-�V��.���z�E�<�q�qJnT�iv����K�������}���\-��`%6��O;���t�Ѣ���m�=�GncTν��~�3J�`�3�2/DF�n�-�V$��+��leX��Kz
�/U:u܇;v�����ǫ�#�U9bOx*C�5��G=F��sM�Ȫd�S$u�Xz�z��~��-}-��&i��zU���N����/>���W֨I�N7D��ǒN8�Wڦ��śQ-\]�pf�#�>��o��|N�;�����p	�Y���(�Kpe�4Ϸ��v�l:���ޘ=�Ն�2Ի�p��/]�W*F�2I��f�]��C|9l� W�v���6�O�NS(�el�T?n�f:�n`d-�����H��P�s�R��6Kx6��Po�EI���A�n��:6<VyX9��EN�f�6���Z1���Nf�3���hJS���P�t�>K,�lp��]dtT{��˃iRy(��b� /9�dD�#�6_Ҭ-�b�5V^���u���iFq�Gc��h݈0T���j4�MxC�}��
�����"}��Ǣ�n�&��z
�t����rR���i�����ᶄ�஥c��VT0'[�\k�2g�[5k�]K��"�"�s��U��5jݙ�I���������`�}�UtN��`���T����hֺChy3V�\����ԥ+� ��ul��z��܃7��h��RHQ|!H����a��ׁ�Q�3<���d;��Wv͹Z��^?Y^nڣ��!v�uiC 3O�Ϙ;b�u�l��gk	W�������1��z��l��J��i�^��{��*�/l.np'�0m�\���3Bz�����V��3�`fd�ou�od�طy��,e�CN�����>DvW!fV�L�m'>���F�N/kx�:9���1M�׾���f�M����>�wV��F��U��H�E7������z��ö宰�O�+��\���d�����c���y��/F��ٹ�#$�hK4�����wy'to 0 ˹q�1Z6��q�9��o���<缼�I�2U�(�X6������mo�ΦQ�Y
n��ym#��?&���T"v�'íZ�h#��5��=��M�G,�w0Ãh=�5y0�	}�/m�yit��*�}4�J�q���)`�gaC.��[���b�V1��f��{v���L��*�pTN͘�11���-|'x�<<R�ഺ�G(�t���vʾ'L�aU�Ht42S��%��F%��4`�9M|4�
�}��ۇ�Q{��=C�3�MǾ�K�[�O4m�pU,�9��8f�{��`ulA�+�{��k�x�H��,'�e�_k��y��aV����f+c#���WRJ:�OT�{8��`��aP��=5�0��fQ��8*�቞ɨ�b��#�X�.|%����;@�:<QY�K�ξ/y�$�+��*�b�Y����pS��N�*�S�t<�ɔ}�D�#����~�/���.�
s:��\��2��bu.ꗚ
�6d�Z�E3�� �m�%�1�h*�{�/1�լ��b]JYB��(�>�b"������05;�H�V�1����*ת�4G	Ut}	'2m�$�场1�:w���{�2�flL�u�g����s����t�Q-#���',!U�7��hM��[�׮:�y����s���n�$���G/-E�%�ܙ��K~���Ŝ�C��z��et�p�F�p��bΉcB8�#};��,��P�9,��jm��5o��?)�Hp���o�w5�����y�_H2����A��R��]�V{ͩ�!	����||�>�=3}�ݣw&�~�jG��fЯ��5�80����i))Σ{urUo���nrȢ�/D�w]p��ɶ�Z ����a���!)��d�����[e���;˞ء�BQ�d��\�H}w�2�cB��%��S:���f���\��t,O���Ѝ9I�%j��RF۷ARێ1�}QV����2�]Nn�:p�Ҙ��V�h�6��r�����-r=O��-^k�4��o�{�<���}϶�Yb1V(�h"+m��cb�1����b��Q���("�UEPU
�T��X*(�DAZ�++b�Z0DU��QTEX�֩m�B�e)`���EQQF
*��űb��X�1H��X�F�EPTATQ���AQ��"����EYl��EEb+UTDb,UAee`+Jب#( хm�E
�mmETTX�b1R*"���kh1�"V���B�aDU���DQZ��(�����Tm��+X�X�E+E�TE-�YX���TQB�����,�,�H�e@�* �6�A�bEV"EcEb2�*��H�m(�XũUb��j�V ��V�R"�1dX�6�%���X�*"�D�F(*�"(�"2��"� V�(��b��YE�1�Q�����#@X,YZ���b�������g���=��ee{��=-	�=��s�|���%F�;����*;[Pp9�H9:�W-�@e�����ӛ�r����HO@�8��r�u�\�)��^���)ش�0on�ӊ -�{a�ܝN�A%�V>sn�F�+|�.����Jn^�/�3�ڙ�;�-mj�=����u��Xm�k���.u�i{�U�������
��c!�;C����Q.��ŉ[us�W�ѭ��!���kn��*ю�wG �4d9�
LR>��=њDK����:��K�}�M����:P�.%]y_�:�����:bA��alx�(eS�~����=���L����e,�XGhf����+���OC�A6�KV	*$��{�Tl��]��nowp )�pd@�/ʒ�c�x飞���oJ,��!\N�i;��vH�f���y�U�/�Ɂ��z�Z �k�D��Yc��.�O�|$՜s����;b�r���������%ԡm�m�.�����چbUttsߖh����]y��r=}�VCry���0��U�C!S�b�G9,+�#�v�+c�$�V������M��V.JM�#����:�K5�V���Q=�d�w��=�w˳��;��;��Y��k�hW���/�$���w�*�|)���Lj'{ΦW-�o/x��h�|�/����x��N@�~�X�f߶:_���R�O��2���q�hk�1��v�B/ܫ8����	��TX�N�G$G�L�%a�uu³oLL�8�[��)s�MV�;U�q_r� �Q
�>3�z���^�HX��Ǚ��C�X�T�m��W,�-?#�0���֗���^)��C5m*/P�V�|�+�&� �у����[��n��e���0�j׬��.��N��x'��\�Ɯ�ɛ��ۛ�vk��gxH^
͖�'����c�
��+�6��x�ƸW�e��rz@n&kx���]�G��:S��L|����.Pag����7�B.�L�[[�a}탲���ЉB��7T��}Qb�mV��n{����r��B��IЌ>��B=�Y��wz���^(���`�E�X�%�mՇ�aqє�����Fzm���#�����b��oa�@Vٯ\ޔ �(V�ݮ��0�Zw��C3-E'hjjLs�j�t)�Ț�o�űb.n�ۈ�XХP�9��)�w&�`�Wy"��'�!坎�L�&�fJ��Q������V��u��jȻ IaJ�h���ޯw��ܞ�oEK2�Է�$3h�nIי�x��J���|i^���/'Y�j����Qr��=n�U�{-X����������=raU���J�2Vs�#����>ǊR���2���5�U�0����*�%u��*-�E�Z���mf�ֹ��=��s��zuz(Y��)�8�N5�vP��8-���^s*��>f���}H�}p�h>�\e�C�{>�y��.�,֦:iL�I#�|���d����l����Ηڨ�mfMM杓�*E�n��g
�3�m̔�}���� ��}(��:�����K��r7�`��ɟX^�X<�rØ���	t[�,M�V���7��^����s^���9��C�0U���<����@}#kY�^�:OX>�ba�aڙY4əʎf-3]>��v�P��Y�}켳�TXa�{c��A�r߇��9�Ĩ�P?D�.�^ʛ�}q��eS�#�o�y��@���6��V�S�:��C|�j%ֻ͎����fM��GR �N��`Y�s��9�-H'��
�n&hE��l�,�̓�\k�F�ԗ�WQ��B�^Ҡ0�bsХ�&9���փ&��I=L�d�!��¬�ӑP|�f�Ob��T��5K�3������;g��1��#�u0�p���	u.��8y�zXe�'P�8����2c���iR��R{�*������+Cբ�+eۧӘ�:,X͂�o/���]�9+�IZm�ã�Y9A���ݍ�݇��g��'o�>��8��%�e��4@L�	�l��.t��K�.��L��zEt��ՁR�q�_W�����Y��=�Z���[��T����}R�`>�[7j��ztEs��f��U�_]�DΩgt�q
~.��<ۿ4aG/�.�ź7�}#��b�i�Gm:"&�a��y?J���'�m����y ��"��m��G�lAnxo\Q�ߊu����J-�aJȍ:�eù�G0�=��f��gz�W��1HӿJO�-)/�Я_O#7�&k�� �U��8g_���k�luk��+̓���4=t ���Vl������u�,ى�%�|qt�$T,D��"�Rm�0�mM;ͱOi;;-����Ѱy;��6'ԧD�S�f3�X�є�ra��X���v�q'���z@�9�b.`�[s�Y,`ê����o8<vj�^�uKg�79���"�nl��f
<o�A��>N�.����~�1u�Gv٩�Yak����ً<�l1��
��vxv],�K������zOM�]w����d�Ei��f���e	}J����K�F�7����d�s��;��bD��Ԭ���<�j~9}Ġw��"�*�*��7��m�- �V�e�̭59�v9WJSu@�'��4b���-%~jV���CŎ��t�,��V8U�^]����o�H�ĬCF����</1���K��Ts�9�=P����=2�F�Lך*>˖���Ki]z�P:�
ל�/�y�P����3�,��C��V$g5��W\�&�=��ӑ�>8+���ꅺ�8By
���,�)b�[��6�vV���S�iF����c%qG	���o��cz8O�*������P�ܼ�E^nh&`�4�>�n�ҋ̼ى�s��^sn��<B�;ٍQ�I�WC*5��څʥ}`�$��+�ITv�������Q�xIw��&
�([3��\mB�͹}��C�أY�����p�PB�L�crw�i��u�i�<[Cِu��:��2(�zA9�����wT
�L�a#r�����MJ�w�����D:��h9|R��S��u2!m9��u��ILM�[�A�1¡�'N�I��h���1j��Sz��Z�a�z�OUj@��R���e6���7����rj4va�]���)�r�Ȭނ!��{��;�X8����4D�	ǶC��颾�W�m�7��yH�Ǟ�t�W�aL�*~Ryp&gY'Ͻ�뷵��؂ջ���;W��}C�������Yxd�s���(p�XҸ���'60hգ����M����{q��"H]�Yΐ=ؼ��ꆭ a����+C��k�3��s<��?;�z���>�������֜�AE`d�v�U�'`9��,��O��~E
�q��ҋ`�0']���8hwf�s2l�[�͜�:�-u�<�T1��Wo��^̽�����glz���%��@�('3l�)�тO��Q��v�s�#6��\��Aw�fO;��l�S�@1w0D��d�d���C�s# �u�� �4l̋��N�t���G�ʻP��[8/+ܛ���6���&}���F`��dދ�-s�uoO5[�L�	�H} ��24��X^E��8xg���[�����r�z{��#��7��/`�mUX�0����*��W2c�u�.�������e�T�R�f��j@Ԥ���+�籚��z��Zj��|h9��-, $:V����n�9�����2� C��Ҥ�ʾ�X۰�B5[����3%zw)g���N��(�*]�"T�%�ީQ����nI���z{�6,
u#;nͪ=��iLL9�J<5p��ȇf����=�sf��9�IuZ�8TN%�|�ٵӧ`����
�1��uL,�����n{���n�g/̪B������Ga��WF5�:�u>�8:���w���)1x���뮅��sǇ��ʟc��龒g�7���O�M37�l��rudÛ�pƻ<�:�Ww(�A�:1ݛ�K����j%�@9��S�r礚�{Q���b�\����ƅ*�|jw.~5�굠rk;��U�#^���2���!�,�^�ėC|�O��J���;�ʷ,A���J�}���g���@wB\e5�9�/��h%(ɈJ�����<6V���{���q_���3D��/;�1eeR5�w~(Db�WL�69�`Z���v�t�Wg���[ZM-�]�l� csxlsZ�<)��п��Js_H' =�@ot:���օ�W}�U/:���J���ߑ��S`� �����K�q�E����F�����Μ��xn:CfA�I�.P�`Vs�m�Y8̅�t���R�t���O�<:b��GaR�ܞU䡋�JMK����.�t,��ȩe���ۇ����Ȩ��k��N�p��8�;�F�w)˝��dg]m�����]�g�M�/�2��<��h��-R[����lC�5���XD\���>
WpZ��Y���y�������=�0:��]�0�С�e�)�+۳Rw8>�s3ӹ������H�Q2��)�"�1�BV�皜��`�ce��V�S��n������1�L��hF�+��,�T�Rv�γd�G:�-Nx����!Tnu�j�=�'r[�E-"CӜk�WP� ��֗K�X��s]h6r�z�1Y:w�����s�0?N�j	��=��"��'t�-�B�2���lic����26����SWw����*#�{�~B����o���<]h5P��\�{��n�j/z��{��]bnub�������с�����W��5��n��F���s�S�z:��c��х��ޮ��K�M�8�U��Yno<��hf�U��_U�^���=Tai�ۮS�c�ߴt5��-`
QC��Q��녲��+"�1%����Xs�\��N��z�i��{���]���fQ��l�g�'ɚ���x���=~�$���@C�	�=����{s��^����trN�fE�H�h$�w9�����͛�G�Q�p؂к��uu5tfm��<{vx�X9��6��Ĭ�>�.��;͎����� ��nnUghL�0�3Et��"�R�Ƕq�{l��P6�/z�J����9٥;��{Ά�ؽ�F�9�kkD�~iM�p��wJ����L��'�}�2�K0�h�A"�:t���V^��:���R���>Xn E��A�e`��J�������i��W��$]��f��]������D���l	N�(,<�W����� �[��2���{&�`�+B���R���1jr*Q�nl���j
"�daY؊����D���-�O���	�N�Ҵ(f1^N��3���:���8\�V1��m�G�ڝtw�{Fwd��RW5e����5&a� Ns���p��J��[��Yv�z�Y������U��_��ڪ8�u�|�7Xz������oY6=��G��^��gSK2E��jy�΋�P�%3�^����v���hO �]K�EZ���/I8��г[�iV��2\gǪ�p̝:
4�R�j�!jf0Tix璣�xe�W�,�Q�h�����~E�ȭ��L9�F���x�Bw���Kˉ�E��ǯ89|��ۻ	�����͛it�\�Ē2��ڏ'�I⤾�P��`�o�������8v�S��2�M���\��v���ه�!NW�E������5�mrrÇ�֕w� ���$�ƨ�'^�a���#s��/8٬S�3!�u;��sL>���o���q���5���Ps����}Lެ��͸)����/`�˳]%i�)�n:e�/�f�ۨ�ʴc�:�4�x�4e�u\6q��ɺA�o:�q\�oFq�@�.0��07ة�],$J���θ\&�yN��c4oco*D������S1��o�4\�خ�gr�t���ILM�i��1Â{��`�܋�x�鷼	�t�7<I�� �b�6,4z�i}��֣�C��W�����#8z��}w]�����!�5Q�,s.�X9���3����]��W��»h+�]wݑ�;�v�9G{Qj��<�ߖ�b���O��5nD�㣥�}�%i�`�c�e���أer�E�t��=�'�E���,JW�B�S�c  B�n�76rH�� 3�8���)�!Ih@�5pp:�L`�%Y99E
N�G$G���K��֎_�R#�𚔝����Q�,�^��Q�6�d�d���*�̌ �G'N����|^*4�S駷���,P��J�x�-�(���\�P���]ϥ�:�9r_|�h�@�)R]�����	K����F*DK$��y��[�%j�v��̣w�8��.D�������|���S�!�{ir�l]��u3�KC�.�������KƩ�LN�˺0j�h�'�5hJ�c�ת��H�B����cb���g���-�i'�N<�e,Z�#s+� }C�n�ʌ���G���vL�.�EiC�)ɯ>��3�����$�!@�{Mƃ��$��/Rl�l[F���6�w�c@����=ʋ�+5�&�kA��@�f+��1w�6W���޲�<�OL�R¼U���I�Q!���M,�h�6s�a�$��4�_������%l���/o�]w����F�($؈\-$��Ս�^AK��a��K����B���>y�����=S�MO�s�^Mm�V��&�F�o .�����3w��|X�V�OQ��ݳ6�4��J�e��f�c���k_f�H���
��ccA�j$��u 4ac�F�
٭%X����+r���u۸����mƳВ��efLu7�����p=�ξ��u���A��F����Np۽Txc�TX�,�lr�r��-Ü��0��:���hʔ��[�,�A�j�v�����XRC��`к9A�un �흖�*7>[�^����%�jY̧��TUƨ{{jx�[�}��)n�t�os1{v7���
]\3�9G����ftՎ^[c`�}ו�^>v��j����������z�[�9� ���])0ms�M���u>��F�[pU�͍���N-��2���R����R�nĨV��_( M,��n���R͔�S�������M	N׽%$�Vu�(@�-d�۷*rj��%���+`�����<�*<(��F;���ȴ��_U�h<'+�-;��S�V�B���h�o~�p�֨����P�Tޱ5��]+*�l�0u��՗ml�Lgew'�mK��<����}�GX�Dث�Ww����������u�x�^�
��Ba�<��\N�{�z�%�>��x�}knn@K�����,v���A�p
궹�� ��	��:uk�+.t;h�֦p��S������|=A�_K�v�w�8X�.�;l];�N���"v��Y�"S	i-/�wj�"}�G�v�h�u��چ��.�.�YV�F}�� EIC"I��ʻsi$��T8\V�*���x8ުH��u�����	u��(�ߕ�3s	5�:qv�6V���P �[VMzUǙ
@L=�)�A9��np5��;#u�G���h��_���!���vժ�{D��:Eњ&�ũ�݌uF��[_�}ô�F���o��v�~j��o��W��o=n�']�gɾ:�N��r��w��-$�a@P�> � ���A���U"��Qb��V(��ŃR�"���
�TERVV"���X�)"(��(V�YUb*�"1X�FF�Vj�X(��X��q
"��2��E����IU�"*1J�X�*�*(��`����E��*���RVb�Db2#�m�RlR6�YmPGR���(**�qj�F
"*,T�"�1���TEqJ��QEF1TD����U�-i`���)F�8lb����E��EE��0b[F"��Tb����1X�Eb�c�QX�DY�VL4QF"�-F*"#QLXTE`��V1�U"�B��E�2V�DE`�����������b�c�F1�)T���YŪ�VZ���*�m�Z�b*���b��UE�lF�J��d��*ȱ-����0���)D��i�0Vs1lv\��]$�Ύ]��7�)!b��?Y�/9{��`|�LaӲDϧ��ۖa���bn*/5E�"w^����������'��1��v��9l��{��r����ToP�i���K�7��������V�14XH�s�����ʲ�\��욲�×l�s���($;ڕ��5P{<	�м�-���0��e�����dǎ��l~d���ut�Ŝ0��@�8s9����I+ԝ�syz'=θ̸��uh(��z�<=�3��Ǎ�9I�.�6M�l�P�8��,c9�1�X��O����t��ԑ��6f���D+���8�9gFuا1�v�}�k
�>Ls��E�����ۼ�-8; GEJ�۸qݵk��e�]�u�r��ֳ���� ����vyRu��Mʛvx�!m��it�uگkM�����T���:���g�.�^�򉞘ХP��|��w=�Գ�A~�������W/����N��Ɏ�r�5�Ρ@ʣ9��3�S�����У�7X�.VƨG=w#X=U�~�z��vX���/��Ƅ�*�a
������;P��N�n�]�|�ɣԭ!�a��ì��D2�j����Wjtj"�����1�3�9�̛���ጽ-���Ĳ20Y�M�\/�*(����wq}���������Pb���㵵o�}r.���]wE!F���}b^���g�����=��zˋ��R�X����M�֮��������: U���T�t�#Uۮ-p�uoވdT=�7#����Ԏ�u;ŵßj��gc�[R�-��TT:_*�ľ|u�R]��[����EX6y�z��Ϭ/v�"_9a���g���}��6�-o��oT�1Ogt���ޡҘ��+(�=H�*E��tgK@g<y⃪�,'}�c�%�jf	|�>���%�J�^��䵃�h��AS�Dk�Xb�\���x*s���k2\�n�뒑�g���!���p9�:��S`��E���Z�O2�xk���%yN���]�k�ڙ9�R�T�cS�*5�#\�3��u�Z��3����ͅ�"^%v�]J�hܫ��d5cC�㮔H����9U�CV:�%�XB�r�T��·����g���]n�4*�)�(+�Dœ�X��N�+�2����q�FQ�X� �YSN^1<�4��N��J���F��x�����4��{��U��R�U5.�+��e����RO�LJ�Fѧ��p���(]�=�o����z	\�:��/��SӺ��j�Q��%�V!�5r�ƴ�;��9	��˩��~�0���7=,O�so���^�u�v�&߷3b�J�}h]�|��u���΄���F:�դ��.ev_XΒ�����Ս��qA\�)�e4�s!��ٻ�b�=��C��w1��;5�8��cDm)*���Vc�p�9:<~�n���j��<��e����qgDfd�},���ױ���X��t"��a ��"�$v�8�tĚ
���Q��{q���K�i�8ɵ�J;/4�5���fQ�N�c-�Y>h�҃Q��q�<
��$���Szm�p_r�e����aLp��*^�Q�7��5��RV/{�i�KQ-���
"�fQǧ�N<ц���1 %fa_��Y�Z;w6]Q�oKT�b�iN�3��^����%��c�f��D�I
= a�bL,<�u�w�q�Å�!�Y��ͅ�y�ե@Bߓ�B���f��E�D���k�ںhxv*�el�R#D���Ϙ띹�<p^�yX9�ѐC�T1jr���2%)��¿j⸮ܠ�6�<��/_1Mu�d�"�G;��4!2]	@	�b��$���]��g�nݸ��G����Z���v�2l���{�������hF�6~G*䳝��Y���B_]��k��xWb^�8��;�Z�� �#��sj+k��Ϋ�V��dthpR�hK�Tq�!�*�*ӛ�Y�Y�P�=��o0��x��C�6��h�;��8nYn��6C�6yt����xpC�-��Q�@rhC�}��!�y�#m�k�v�Y��qlwփ�۪-ϊ�/9��
r����wx��'k���B4̅t;���y*����O�]e��7g��[FL:>=�f�<Ri����O w�[��uP��!Yƚ�c��WOBH̿xؗ�9R\|�R�o��g����5b��mɆ���6�]��1�}Yh'i��(�p�{W%�I.�j9/��{�(wj�9ZM�U�Ru���S�X����/����J}P�Lgu\癸S,0���kn�cN�j�S��L�CFj�`b�=
5�;lK�]E3p"�.5i��U�3�Xl۫�;��j�7�5�jsjh��L����W��,P�D��ۘ!D%: ���wq��������K�CʤYy�<y�T�����Y�)D���0,t�:"Ivv�|��UH��	Ҹؘ�MЯp�Bb\<�=�,��Ƒ�˵}ΐ=�����$J�X���V<#,h\o��H�Gqy<٩�����}V���'� n���D���)Y-���Zp�Z�>G�Lμ;˸�[�JQ3�^�j�}�Z���׶��d����Kty����6f�RBz�FM�o1P9s_��`�h�^�kA�����O��>=M�=��qඕ�/y�|,�u�:+(�݀/XZ�I�j�zr�z8܁8�̵ܘҎ���66ۨ>�K�����}�����61+���l�:�Z&J>H�f�eW����t֠S�.�=QOӵ��(�mM��f0 �/xڕ�����-h��JG�j��s���	�7�C��ס��֫*����̨"c�Y�T	��*+���m雞�!O�#�wb
�z;]�s�ESU�-���7)�uT����M˼�\V-o�IԷ�3�M�Ԍ�|��0-N&�Uԇ� �?�FZ�>�o�J�����m��)�'��k&ݘ'Q!j�V��M��/`-���8�e�F���I^(;Զ����W���c4��s�ĬK�ϵH�ԏ���n��s�3:�	�<���MuU��u��}e��9*�ˁ_0P��M+��ۨ\NUC��f���ze��2#��˭�.��9�+&Jh�b��2��T��F|�3���2���
�q�����NM�9�}���j�S��zwSz�j&��ԁ���|Ҡ�ݓC5����1�י�e��˜=���yAY=׎!z�(|v�fS���`�/X�a�R�R���]�ֽ���!��Xw�i��sq�4ag�{�X�T�h{-�ώji�s�ij�ܥ�e����È���{"U�r��ޏa�P�[�V�SzP���_wZ{��n�/I���{�b#�xbR�`q.T�P�gg��gFS��r*��H��$e5�X��Q�+����0l�s��Υu3�:X���t4�\��Ρ@��q�汜���Θģv����顺�[�F�B͌u����������+!qu
�pz,���:�oj��05j�Ҏ��.��h�6Z��0���N���kWB��
E�8K�c� ��d�;r����%5K6�@8��Z3�g"��o�^��E��"į���N�)M~��e>׺ ��	݃=Q�$�P	;�F�h�T�g��k<�}n`vS�3�)�oH�3�ۜ���s�ej���kQ�󝊖X�C}�GE�"FI���TE�H�#kY�s���8wWz��^�'�ANX�N��`⭷F��jKyb�
�o����
t�򕸖ZP�WVr�9v��%FwU�|�*}P��	���>�p���
�§B����or�]�lO�6�i��U�J�ʖJMf�^�r�j�Y.֎�HT�:�@q4%3��j���`j`��V۷ֱŹ�û�j��r���b���b�;���x��q-��vOMZ�A8�f���=�581t6�@�ý n�ܒqK��Բ��7.9;G�Q�K�^��S2s\�漩��5;�\��+]a3\��'��`�c���R�h��6��v���C�<�z��`H�&`=I��bkХ�'��`�5u���J���f%�i���d�7�2vٝl��=�,a;��ܝ�Wei�f�@�.��U7�t�^�ד]5d��ndM�9�����E\���.S��4�Ooؼ���K9P��vV��;	2���p�X]z�F��(�`���e5�wd��n�X�v����E����J�	���H�9k�H��Ua�:b�i�Gm:�>\b�>u{T�<�j���L�]��r���!�H�5��W�*�r8S�.l���5!��[jO7+�x/�}}ѩ�6̉���fQ�������O�)����Q�CBx�C��#Rv����g)V��r�@�
a���=C.�6W�ŇWu��u$�|��<�Z�[[^�ܹ8�/6������xd�C�MG������rx2���a�;�[�V�n��'[f�h��N"�����C�a�u��C���8��[Dr���0={R���e�
֞*,��=�Z,���F�����9���'��DnŸZ]�J��YT��mm:�Wܩ�����Y��%y:w	n+�`}	��(
��-M}W�-&C��<�ͨ:T!X��"���(�0�G�Q>��0PXy�,��+����h:���u��Ȁ)n��eW��.M3�"����o�j�xcȈ�s2zPj�qn��~� ��(sV��\e��(�c�؇�Q�Lm�	JC4M{�x�k/�Ll)m���)�+�QŃEJ�5�R6��'�x*3��!�l��^r13C��n����o;�U�J~4:�j��<�b�r��^"s����)X"=�m�f��.3�C{;��V��8,`"'Нԇ�Yy�,���>����B���+�K[���T#̣�ޫ�/�9a����oL^Ts��HK_-�����4ڮXW�w�:�0�U|.�}Lkd���v�XP����V%q�i�r���Ƃ!G��e�AA1;s4�@$sd~�֭d�p�p�yS>�m��[��=�֡ݪqiX�L�\��K׉�$��cQ�-F�w\mG]$g9�mL�ũ�nCn�4�Fu:|i����ۼhe�=j�9u�e���r��=���pc���E��e\��B�rcn\:�%���9�z��B�}���0.�̥�]���V���U.���3���M�r���)��ŋ��t�1�hR-�3xI%��.{�R�{�y�K��t�\hr�=�$���n�}��ULK��GD\�Xi��U�W36��ͺ��θK�Z�۫�GbZ�����?[�$�V�Cj�!sr��|�/
JbT{%�1orO>goM����֔Į5"t�}�$�PN���т��7S>J��R:�P�C7357a�-U�����O��r}� >,�{1�����0�.���2G��CJǂ}�o��*�7�n�Z;�p�@�U��\rz�'���l�괱��1X�"Vr�������}ܩI����Gl�Pp%q�c�������,t+��
��!Rt@nuO'���IJ�]u+��!GwTS�uϦ@��d�:4�ļ�;r��.��U���g=��ws�>�8g�#�l�s#_�s�S3�&6*�����fT��,�P%�5xT�`�#��O�����P��v<̭m��@�⽥���q˧��.a����\!�
������T	�F�׵;:`#a��WRd4=L�8*rV�yHnW���|����Z�z�\�y�gw,��Z�v���Ϲ�|l�	7Eg��&TLQx��� {%-y8ƾ�3��9{Ԙ(Cc��,l�9N�s�'��즬�y������.{�4��Q�xq��Gd�`�]Ú��p@K�H�{I�A�D���bx�{�d�(� A�)`I�Z�ۉ�u�e�Z�60k�1��G)��S�se-�$�ǵ[��9�\��K�%��_K'd˰��
^��З+�pt~ru��f��h��j:�E�J�r�|�[م��V��5��T����P�]OL�� J�Fs�����<�7fC�n�N0�
詌��R�V�@h*[�Urqx�(tJ[te�q;�{'vܿf�;�6�`����,^+J�G��[�k��)�(:�\��ʼB���ӻG=/fe\�K�Je
jP��c�b����te:�Z&M腌7�����驪l��l�C�HH���J���;�.��p���5�U�0����D��m˝���<kv�+;UX�qu#�c��^�)�d�.��2e!�hO�2a
���d�U���Z�
M��P^�]�"(��]�-U���h��N����t�(�1l�,[Nj���ӎ�ӻ�ڷ �|�~�:�r��o�Q-^��e꘬�x+�
�W3�hR7+[�
���/6��T`専��r}��l��Y|d�>Ļts!,و��pffI0�<~�ONg���ʉ�L�h�뽫j�E��
1*��v�W+��ESJ�l�Y0𱇅�逽ʅ�Z$t�J�d��s7��<D��%e.�	|��i�)��3p�D���u�l�`��.�n�>i��I ��b5��ȝ-�V����/�m{�{�K�Em����I�>���Y���F�>��֤/wM\���g!��=��Z&oO/>�t��38���o�|�((;��w]0�ɜ��n���\x��i�_v�!��۱QL�HJ���d���uޣL:J^ְ��5�Ѥx�z�c���S��@���Glc�4:�%GEc�(ձ����ѥY�;cQ������oNƲ��VU�y�,���j��u�1�6��Zl�==:w\���D����,A�r�8;�\�n�����Z����gj���wh��ai��m�Nr��ul���ф�U�^ &@r�r}9.� m:��3u*ܥz�V�hM�O�s�8F��I�`�V;=뺚���˺϶�Sj�',<l5��p�����~�K���5�PўC%�w�*�B�y���ݢbEk��� EC34B����3�`n��B�z�yQOVE�t}>铯��q�b���FG[f�f\=s�|�yP�����Vg#�E�p �$9nFf������kv����{�(.7	�(�k*j��.��uj1���ݺ@�ӐCM�#�'+%���#̡N8p	��oT4�}|��<��Db��sa��k �d��wf��y��5 �����}�YhT��,R_+J��M��!��%�g�.�Y�e��F�F�6��A��O�B��k5��1z0̽�>҇'�7��{NK��L�Yד�f�'��-L�Np�ZB���o��@��3�^�g,�-�;y�2�|/�+3�	��M1t��C^���� qjK�xa��X}ۼ)��y�K~���봢j���a�#�ץZU��;z�bS���w4�sc�a�e"�PO^ᙈ�4�}�͹($d�oL��of��r�;
���7H��WfΝ���D�ED�K��;r�! P��jE�'K�-a2�PJXl�-,���`)
87/��)۵A�(���u�s2�&����
8�Wq��m�T��$N%�t"H��DzؑI�9��Q�to�yS��-@;d�co;���ʬ�еL��s�|ZA�m	��9��M�:R�ˊ�ʶsu��²Ѭ�T��c��uq�}���6�4�N
fi���._��\w����`�}vۡ�L��D���:�N=�COs��(�BŎA�O:�I��S���bmD�g���p)����/���S�}��)�KfL�F���v2;�-ɷ�j�M��o��2��Ap��Mm�a-ޫgw[l���k�";J$QAW�K�`�E���F��ETŢ"����*,Z�h�".����ԣQ��\`�+�J���)�q(�b�T�Ya�Q0�
�6�c\5P`�m�T���űTTX���Ve�+�UF$m
�4TEU[Kl���X,UTH�+J��\Z����)�f ����ʈ�T-�¥W�1G�T(�e�.-�"Ŷ�R���DdQ*V��#Q���"��b��L5�V"EDQ�"��YR"��ᡆV�
�(ZUDT`� �j,V �EE��EEFj(ZX��F
��6�U�ȂEQ	LZ���%l�1�����Z����D�VDAH�*TS$�Z��"-�R

�kF)�DdkAdW�E���ԢMQ}��n�]�qt49\Y��� #�Էa�wq�'��uDNs�ѹ��2�
���jjB�5��Un���2��ڋw�KƱĬV_I'R�s?$�� �d�~��E���π���z�������4�b7�~���q�t��u펒��C�SQdVQ����e��E�f`R.��5L�j��}s���@�yQ�Z��T"�Y�3�[�+��O3>�i��]Lhtg�1�Y[w����Cw���?Q�˃����n������_T&�X&rϰ-ˬ����5:5��Z�uW��9�t�b66+ɪ�ePPמ��^r��? 
�N��`Y�ɔSC���f�)pR�t'�xs�2Fߦ]��|^ʺ�d���K���*�&�K 8��gT�Z�V{��չbn�8�fOo��~mo���O�Ez�������Y�:����Q�������'�6���ٱ<iYS����Hr�ld2�։덖�Ɔ=Y�u'g��a7���u���
��wmh��8��e�^wK|.t�5}v�VH%U�1.BR�y��;��D
Z !��L�V*���+i�GK��q��ni�h٫��
��o��6���� �Ŭ�ڝin+}����f���.&i�"nx6f�l�+�jS|��X��33(���h^�C��3 �CT�ѫեST�i�b���C��3�y�_V�iG_bYS���v�Vv�Yr!lV�jy-���7��mPB����5��WU�G
t����*��&��$��To^��S2b
��V���;�l��E�F���rٛ��4i>�5k�9+ΰH*.�<��;�뫯<���/�>\�U�J�K�TiM򿡱�)\]��ntdF��ef(�b��zT�ٝm�i��+��Yx	8���_^�&�Y��rTPy��Xe�EM&����Їn�����낏S��1�E�Y��d��G�&�l:y�[���͹���)|b��]{�Tft`g]k+Ac)��(_�M3�"��sd�0Q�6��<o �9�k�3Y��K�����\�����p�(:�4b���-NPu7�4%)n�Z��{��6wi׾3]�Gg��vʧβ�_�)���5%Д ��b��I��^�4Ů.����������`0�B���F��>��U��q�5�2r4�Mi&]��:�uw���w&���i�܍�4@E{}۠S<BтR�w���S���V��L-��J�/�(���MR<��1W�<d/�%�����M����cG�,�[^n�Q}Nw$6;=���ѫ�ល�	�1ݓ�Bh�����y_E{3�n��=���! �[�VuY	m�wB�&�Q]S��i �l���=&b�=�c�X�̥"�Ucji���Gv�Y��[p�>�Ga��+%c��1����)�Z+��(PDŇ�#�2է���^*S|����A�W���(f�ң9]��r�Ӟ}h�6�H	��,Z��Q>����5�����o;�j5���fAӶ�hr�_�A9JS_�������P1t���<��)��3A����Ɲ���4L��\+Z�c꥙}xk���.�-��ǨT��]Y~.�yЬU��6����������y*��euv��ʰ�7I�văA���C��tlW	T��U
#T�J��wr����Y�޻HN�`W^^ܽ���s�d�h�%x'L�����R^i}�)�6�u����d=�o�-��CM���:ޕ���,�#2�E�s�+.��xt�$_�v���h�[��k�N��x�Ֆl
�xp�g��x9̆�wZs���1^J �b���T�*k��5�xX�Of���>;[�`XZ��cν=X*����:�]	\�'�@��7�e����S/:C�&�>��`o+���[���! �7�o���zv0J���M��[��ܙ���=h�`�pB�5�
�:�c5j>G��{]7��c�t�
w��YA�`�+��0�{ȗ�r��"���<mz�\���~~��[j)�f{�W�"1Н��\�ڭ�'�J�8<�U������P�yi��a�v�����2^�6��}�H��(y��O=6�U�8���Wn�_Y����j�qܽ��mcӝ���lT6H�J��-:��%H�j���V�/0�阩��۳�r<�Q�@�����A��ၰ��^Uu!�@3C�6�e�#J��	t[��F�T)��,\%U���Q`I�Q�����:�3Hł�	��UK]��jk�
j�(�ц6��P�L;��O&6Q.d�?*�����Zů���	�Z�R�z��ԟ�K��%ʀ���X'��&�����p������Dk�ac�-;��ȭZ�u�95fZu�d_5S'.T�e�����u_�_h')�ҹz&�s����[��k�zn���{��5z��+'(��j�n@sH�ú�,ed�^��)�(%b���Õo��_Vj{M��nWtߥ͇���P�E�LF���RU�v=���&|.]��/(�&��]P�wg<w}m�a��**��[0#��a�J�t[�FB�՝���Yh�b�]%O'z�b�8�N�(�(晷u���\8�o�`�=�c�+C���m��/];Pj��өmut]�qt��6VH`C��G[GM�;Cw3��_H��}Ԅن��J��w`/]8&W$��8�-���cػ�Y��_c��GgoS����s+֥#7���,pL�}��4'�W�@N�/���]���3ש�k��Q�_aqFp�r.�
��ƈh�d�ZmkWB��H�ǁ9z:�Zz��⹊�z�Y�I#l,:H�l��$�mo�XKW��Kb��:� �q��,c���6�%8lN˜�q-ӻE� z"�H��"|(-"��gFz������q�q/h'!WU�g��\oh� u����SZ�d9ةf��h��e�e���p,3�j�e��D̗��-wN��j ��_5F�SKp���6&t�q����R>�C��{z������s��5��$P��x=٩:�&w�X� c"5�ˁ�q����Z��X�A0��N�{�r$k��N�d£~f9�:�R� 3���`a��Ş�=��r�}u׉��WX�M/�V	]7�K���/CV&�Y[��U=e��G��[NT��&)���,��vu�'P���|�4�J�K�*��z��S�u��Ldm���� Z7n�U�,����A�@3�ו��pG��&߸����g������s^Y�:k8Jދ�pU��_C�r[�X�άwq�B��t�/2�9��2g��Ρ˶UV M�:����*d��3�o���Y~���*ռ��o���+&�Eh�x�J�.MQl���x,&wJ|��jAL��K�O��o����E�{��N��(�mB[�]1~S\�xD0�r`ãӞ�H���~��Uq��W�h��m���3��F>�y��)�`Ld�@�q�g�H��Ua�:b���dv��l�.1vhNN�#�l�*�~_��Sk
�����8��L�1X���}��WU�D'(/2��*aE�:�K���\�N<��&:lX���j���XR9�2�bub��fp�����qiKi9�yX&,��~�=�Rm@:ҦT0���]|M��q�t+�C ���Vl���Ԓ��|V�T��6���t����_��3W�m-J(�&NP�h�j8���G9<�ea��n̉�㒅>�J=�-�-N�X�T�l����[v�'�2��9��B�&�l:w5�ۈ����=CT�'��y�����1Cz���^:�YP��Pn���򜊔o�͒��(�K�UA@s'���R�Q^X���c�w�F\���l����nւ���%�c S���k�u7õ>5^?Z�}M����{N=ϯ8���^��jGxo��O{2^�`��ll/w�9�-��v�r�$d�t��s�|R�,�nN�7����S��*�tB���,s;�Q�m��|z��XR�S�k���(�c��𜭏5��wQ.�4�wo���"5,g�_t�>��أ��]
쑴X��K5Ě�n�b3�m����z������K�U�.ʋ| 5V^E;�Ul�Q��3�6+ϱ�]a�E��*5�+���y��6�P�`���)y�����UYy�,��赁���{a#��[s�}�N�vk$U! �+h�{�#4���225�5���'�,�Vu�]�5�|���_��t&�����VLX�E�^�d)���0N>�T�o��{Zp�M���xyy��v�z�����&2_-L�7�}�Ỡ��X1�ۍ�,wL��K*�Ŷ�g{w3Y�*�Eb%��h���
.�3��7�S,1p�h0�{ڄO��j0mOJ��q�������0�>'����R�:|e
�7K�L�r�����R�e:8f�]C���{�q��Y;�a�a�/�ꈷlH5�ӱ�xNi
��(�r���S}*{���G�f��;<ài֠�A�7z6v�"'�}��=⨸7�~�ɉ:�t��d�+�J6'ѝ�{1MԜ�A�}m\:�_G��[=&�/���J�*�܂��:6]�(J�&�ng�.ްq���ۨn��G�����2�8�`��wA���nY�pw���ǲp�6ԢMx'L����R^'�[���m�E�F]M���\xٿ��`moJ�Ř#��w��EÝ {�)bkbD�"������S�2c�k�k�j���ѡ¢WU�����uX�
 N��LLj-Ȁ�ٜjd�w��˪�c�Ar:݃9mƨ3wׇ�u��i�4��:�]�N�)��;R�ꖽ��*o"��Dk�=��^{�HMO{ �zc윱0�6T�f���o��l9ҧ5O�UY�� ��'�o��:���S3�&6�q9��ʂ-�"�sD���i�$޴��(�=:�ܒ��*��-��VG�fC���Y�S�8�E�������u���=���[j��/P��·�@����<�C۔
c�^#�8t�@���ZlK��{޷��Ӿ�X��w���N�bx�(J��<	�!x+eyU1�aS�>����(�R��S��PC�1a��D�F�&k�WH_L�7�r�$x碓�+��-b��|�'����ze���o��q��+fq�Ӑo�{1_;%g���E[�"=�s�����l�o�o�*���w�ܹ�$�DҊA�z�$(�5K3$���K �]{C6�z�Sn��+]2����GB��I�����.
��VR���&��ܬ�,��3-�a-Pag��`�#�M��P3�����R�g=���.6�<���R5q�U�(8M��j����sU2q�(Wz�2��� ����悯�������ȓus|B��Z�VXvX�N�[1�p/R׌���=x���G��(@�ʫ\�g1��/���FMw��փ��XR���6�em��"\�(-���j�g�.�B�����w�}r]�d���7ڀ���#n�J/�/�>��w(�C�B�;��R�`��I��Yl��#w��C�����9w*�qa�	�_m��:J����A.2��5Kz]t�層;C���`Y��k�g
g.����0��:Z�Гvl���GL�����^��g�O{� ���&n�h:�z(�����éj�\�"���rB�ء�Y<��G`{#G���R��N7\p B�� ;�P@Q���/�7����+�W$ϭ�r��lZ0%1X�ɂ{�un!�9ةe�7�(��r�H�8#tVvq	é
b�(��v=�N��gs������D�!T;N圮"?�w��ɓ���ʩ�}�n�C�(I[=�纍�X��z��@-��;�T����T��Cfht�۱���{聾ș�EB���m��8[ohC��r���8H:�Gx���>6'�Kt��͉�W�G[�k>뫥'������bd��uy�u��R�R,e��(?n�I�j�L�)`j����p/�k�OY�B�Z��Rsg��m��|V�*Ŗj�S�"��v ���wI�&S�U>�OkW�Y�������G��*�Cn���N�KS�gG0�lL�1���YWP�	ip���d�MbQ��j��O ~���Z
.�m#��`���Y�n��'%}�z���y^��CnG�y09��I� 5��`�\��zg��6���(:V�h+�^�s��i�~VOw� Ǧ(�z'�ɹil:ՠԀ�LX��L�Lq+�����Hj�8�t:+�SK�2Χ���7�+����2�>���Y %q����L��5�锊�Ua�7�\'��+5��4�Q�\�����S2�1H�Q��֣�F�%{T�bt{�����
��AN��5�F���7�#����՚�Ӏd�4�/��eq��;��r(��E�F���7?{���ãT��<,;h��>kks6�;�^���E��)�>���nP�`2�%1�DT���tb��� k��FV�pc�A�$��pL������ұ�Ͷ<��(��3@�&]C�ʖ�T�tŜt� ސ�����g-ִ>�"|�H�j�k{k�����+p�NV��i�K]���[p��S$id�l>Y�>�7ɬ�A��Ŵ�����^�淲$�[xT�ӡt��X��u·Pt�
�T�Z��<��K{]�`7X\�KGV�,	���C�cRy"����f���I��+����<��.{����|����D�;��=��d�6g�j㳙����)v��av�xW�Ή3yky7�ݓ���ץ�c�|Eok�Y:��c밲�6��p��"z�����چ� ���Ύ��>�b0���xFac;MaT͎���h���S@�,�9�b`9���Cl��FS��0�'����p��ۗι��ZJ�q_Ra�|�'R��M_^uBL��\��,.s!ٹ΂.7��*����#ٝ����n4�����4Ui�Y�S�1�*;ur��H3_W��j��>ʌ���Wڔ���PB_a�&�f� e;��=�c����W��n	Rw��txam/%+{��]�{p� �S���{��5Ԣ{>���r ɬ�W�9t��7y� �`��^1�fl��ZO^a��l�{���Q��b7ȸ'���_y
�g�΢�,uN�[v�kj>�]E|s=�f|��rc��U����Ns�iqׂj{ܟ3�m�%�p�������.u��g&�4F�Kr.s�Kە�k(r���k$�ۥIae)�w��,��`6^ú�sˏ�_	�{2���B�a�=sW\D�/gP6�с�'�b2�y��5.���5y���r��F)���pC�8�\X��[�FC|�1<���o�r��g��M�zM9�W�gv�ep�w���:�g���7�gb�q`v��^r�}��'�= ս�R����}:s6�Y����c6�ӆ*��k͜6ƃ;��&���u�ᝦ�oJ����Yr]����+E&�w��Y�V��	�Z���ue��Kz}{�f2Jk�=���|Nb�D�KV�J�
��ڻH�i�ɼ���7�
�����+C*�R^��U�d���w��|�R���;/�.�w_�,�<8�jv����^�`<ʓ�B� �\�,ˤ�	&�f"9�Q���A
���଄�p9�WT���y\b�O����6Vf]����i.V��]{^*��oO	 WQ��)�[��.���:6�'<u$+�Ѕ��M��`�0���0�d��k�M���O@v��,�.�HYG�u�b�^T�xK�c�ʹ��k��ݤ�GSʼK,�8ޞ�u7���E�� lj%��IY(
b*��;#�S�����(�澗�&��k������+p��s*%�b�X3h)�H)0�X
���� ��ATUQT�����m�E"�1i(��&DQATP�n,��(�ҳ��ب(���	TPQbA�ũdU�
3	*",��*�Q��*�QA�QQVa
(����)l*����\%*�����*�db(6�H����QPQ�mf0UX��*���
)V!U��.�c����H�����V1"�X-jR�8�0�QCb[**[X����e`�Ab�����b�bň�������,X,X(((�������U��*1��l}��W��:e�\�7�jz��٘;o¦��69U�.�5�ѯ��w�Ծ��n��ma��A��L3F��ul�*.�.�o�%wZ��{��z/O�.|���L4z*�iM򿡃�ҕō�V��v�q��.:v���`O;r<�^�E��&L�P�h|6_q�|��"�ܧ{\ݬ+3oQ�yw�OeF��̅/[�iVݳ	�T�~�"w(�@��t����wv�NﺟmnF+ʌ�S�M�Xg9��sD��l�Uc���%bRY�*�i(m���d��;�<�й:��A������;�%��Nf}��w��2���8����-��^�t|��/�)�������WB�$m!2\ �Qi��h����y:;�I�)���@��&hm�-\vL���\�7�8!������ Ur�Μ�<�S� �!Dbrp�,`"'��۠S+�-'�9ߎ���b����N^q�)�518cz
���*�b5�8d_��5����3X6�:wL��\��ީ���+��KE�4����6��
f0W���(�b���~E��)���I�g���n����H�|s��;�t$�gpV�+vw2kt�W8OV���ބ�#&��*b.Z��z��Ρ4xŚ��;���<r�1_4;�� �:���.�g��K�&�8�9��܉;3�a��J�,eG����|�X5��w�.�hbU�C�%�A~z������r_-L�6�}�����sa�{��j�;e���잉��%�xx�����(�׵
��"��y��S,1jf��]Z���O���������`���!~6O�ЧGO�(n�e�����6=ױP��;Ǫ�u4�G��j}�u��TѾ�văM���2�ۘ+��;��"(�w�cw�7|�6:m(�'�n�3��S��*_R��^{'	�pԢM�p:y�*K����`켲�0"��_��UH��m*������`����G�-E�[&A�8��y~!���=ࣣk�a��C�U�s�3��8d��ᨱ��Gml�l�4��(��j�O�`����:�n�:kŵp/�Sӕ�ʱ�T��ga�gʼ,.�cn�DJ��Px�m�wwc��H8�: 76rH��S���گ�@��.�a�O�7Y<�����5r�e𞕣�v�S҃uU�����.Q�^�_���l�ѝ嵄xs�E�I��4��ae{xm���K��`�u���W���x!l��&[8[C�Ϳ�J��;���联���W�w����n����A&\Χ܌'k���X^�"ߎ�7'��Bq��ؙ�юC��sɥ2���U�&��SY�yB+yޟ2������!��O�*�y��p�F2nVF㪪C�D��3/�����
�D��]�\��G}�t�;j�\�c'��7CT���°�bh��u�ћ�UX�W�]�y=�a�WJ0#A�M�a���/��˶pl�B�:�+�`'�B�V��t����i�H^yʫ�� u8�B܉�����L�ԡ��:����G��'`Fð݇3-ٵ�6�v�r��XR�8�@A��U��(zm}�'�W^��g�׆x��;b�+�-L�e��3g��0���گ	/t��䑞�>�j���5�CK��PT;Y�~����Ġ�y�f�{7��U��Ȁ��׭��0��ȥ��V@j�kq{�����^ �>2���^�0��M\
�T��KJn%M��<�m�!�T���v=��E❋�h���}�?,c�t��Ӛ~����H���dJP�0Қ�S��@N���َ�$ܫ���%��SX�Z�ݱ*��w5��ET�o=u!
�s*Ԥf�upX�����ob�����V�Dp��/tM=�gPwv��K�&�
Er��b�v�� ��I휝�.�'WN]��t�ɼԞ\�*:0��q�������aP��#%\��S�o�e�lc'>Dm���$�r��c��{�;�kNǑ�Z�6�kwQ�R��{�t��%vg8�g��PP�E�(wU�Ჰ�6S..�
��V/L4r���i��/v�t�qIhQ8�kePl�Hߞ��]�: B�����ҳ� �[V`��/˺��۽1�X�m-�E20Ȼ���[R�-��TW�Q2`>�E<Ѱ"�>���E�1�e\�ܷiLڻ]�֕�Ɩ��n��%*�C~���P�FM>�v��!�u���fs1!IGh�3��1d�29�z�>�T*�'5���[n��2[�[�b����t��Ý�zL4D��7�f���-Y�x6m�9x��xU���g��A<�k9�^�r���\���0�2P���FP�,^�5]�
�m���|� ={Kl��	wL���'00���XJo���WE,+�s�'����]��Y!�&��J�|�m��;����\j`](��Gy�K� r�T�2����l��=%�'7e�Ǌ������K�u�?C3�b�Of�Fic�;ųbxҲߦX��\rC���6qL>�Lʛ4vf���q8l�:���+�aNA�3ukD�v� �Q"gGy�e_\*�/H���\�EY�q���{R/��Fv�E�4=+L�ӔnÊ���"�z������<�u�G�4U�%	��㹗����*ĝ�����G�VZݰ_-.L�:h8O~�_+�=	~������f�0a���}��դXsl>�=��&�����:Հ�d��Y %��،��cY�{�R+!UX}��B���&���[�w- 2�ݵ�i�Z�0���U�������Pc�7��XJ઱Ȗj�͜y�j���Ot���Ł�/�QY�4!�.4�1��kȣXR4
;�X�r�(���{�V:������~x�Gp(jq��<P@��O �l�~ىY5S|�cY��L˕��y�r�v�[�������"睊�#����KR�f@n�� &��/L�aYל�¤�����=�Cxۋ�^��4\N�1K�Qr��}o2!�:h��=(�&/Z=r�$"���w���2C��"x��v����-�U1��uV��c�B����#W��*�_�;.�3�t�xúI��	�we��1��,�������p���-��}B�ߴMK�w�oR=�˯r879A�۩�)N6��Ҝ���b����S�\�F�
��#���Q����Z�z�}�}����So�z�a��.�|�-��S-҅�:��SS�ܹ�;N+d{V���g�������Y�^���8obd$淞/���y�ڃ�g�ͱ����P�9,dOi�{�9u�i?kuM�ս�Nz��Z0��ǫWr`�_��^����$���h�P,�	�l�q�3Ϧ&���Â�S'4�Wts��w@��>h=J�
�m�KM
D��<���"xh�N��y���=����mm�f������Y��Я!o�JHK3�X��ѳ##^ѓ^ϏT3X7�Ǖ���=&Až�_S���gZ�m0�j�1p�cF�����6�ō�FyЭ��T�_���k���n�sbS2�Hh�<��N���v��/��g�ϱ�R����A�.ZS��n��u�&���)ݮ,>��pU�u��赀��c����m+b䡇1�X��s��wϐ�P�j�F�i��qӾ���W�K�>�eޚ�\���uxK9���ܞ�I�M�h5"���eÔ7���s���4o�ݱ ׃U��!��WT!����r+�h�O+��ޏ9�C
�l�3=[�B�z������e6#�����!ҡ,�����U�]��&;p)&�����Au_M˺;aq�f��݁���zVe��#0���;4;��%H'$��۵��]��֦�*��γwp��Y��%ڝ{/�W}w��!(�s��mCz�U����S�1��"���hf
(c~'�pz���~�nEN��M�u坾W�|�B�MT�q=xeI�^�*	9��j�7��.Z�����L@^��/��5%����к���p������:<�X�{S3���Y�'ݞ�@���Y;���s�o������ɰqw"g(-!.�#�SӞ�����*ǝOV�ixa��{YSS&��J��s��j�ӻC�*��܌$v���q.���&�V�8C�n��|\Q���V֍��jj���#
T�����r@tz��P��n�U�Ujٌ��Npp��Z�Ƭ��r�y^e[� [J���+	�d���C�9���UX���@nC2���DZ�9{���=B��š��3����0mm�;)xj�־V���>�������/�Rs#-��p��H9�]��e�W��Y�����Of3�l�B�:�*���6>r���(U^x��[}������\j�v0O�V�dǎ����>�/a�o������]��蒝���%VZ�o/D�'�'�Z�3�j�g�Лt��{]+�+N�4�-�V��H��MhB��Gd�ld�mW���Gκ��u�AYo/(u��z��}-Ćs�s��3��d��6�Jn]cOH�����,o��.�n�A��c��A��V�һ�)�vs]����������Ĉ��y�yv�I}�:�:΢�*�{ʞ�8`g�A�>��J���YɎ��^���Ct���qNޜMYf).�XY���h動������Ug�~���(�9଱��X�c��QKkh�W`�/}��+]5�V��7�[ά�)7(	��!똝�IMʛry�*ۦ)�������)M7��+����sS
�7�ʼ�t+J��@��4)UC�@u;�
"wV��gxt�ǁz�i���6T˜�����ʎ�:��sX�ET�o.�!^�1B�JFo'Qa�	���Hb�L[Jw9�t�����Ĭ0��@^;����X{�g
g.�
����L4se$U A���e�|p����R]T�:���Jg��H�I�pS�Us��6��� әۥ�=nF�a���t�O��x+6�d^2J��
&L>�bE�W��gF��ɘ�f�^��q�7^�*;��`�����{�0H�����k�x�G�V���������*W*z!���#�Ga�J�}���ٽ���B)��J�^o%��}D���2-�+���M�v\�V��p
�xP���2�(n����e)`N��<U��k:.���+�����U��(-�J�h��T��9Pkf%�OFr՜�Lr�62�C���������P3@�Wz���5:��,�%���=�N�&��F>��g�~}���6��6/��-���17�]F�S�|�a;��R+���U�N�\�i~�=n�;����鍀�N�xSMWCE���U&��@sR[�yB�{q���k��q杁Q	�"��5ΰKS�gG[!Tm�eٌ���S����by�s{YR�h �C`l��Bk�2�u�Ʒ����m#��V�!f�k����x���^�%����ś��{�7��2�FU���gtȸ�9��Q��D��5�k���Fr:f����a,	F�FQ�y�6P1��tΩ��L�s�ŏM~�7�^��Cp��R#5 �������w�#���O��q�ht�i�1)�+�k5�)����,B�R${�r�c��΄���ĩ_Z�^��c0�.�%�W���J�j����r�,$:�f*k��Vk5�8�n�Ŗ��[=Ee�bMH`��2�e���]��p�/��83r��)���\�Q�(k���/�|٦��y�E�t��	.��^0��F�Jɉ&���1"����Y�mM=��\�qw
��3���'���f��KR� ��2`T8���@-Z:�H��J˱�������A���(0�Z`�w��2cYº�*����
��|�<ZР{��k2p�T�g4�5�Ϻ�.��W�������*�	u��.���5���*6���ͺT2�a2���8���i[���h�-�Gl����p�ۖ�A%*gJ����F����2���y;��)xj-�4�nٌ�},�c���`[��&J���7������B��:��Aa炅�u���i������B���f�x's��5	2t��'%�����f��sd��6��Qںt1S�j#�`zv�n�����1��´�
x��hi�G�9AҟkL.�t|���t�),�$�
Ϯ�)����˸tS[�ok�9�T��	@	��)��rN^�^sG��g�L��e��ș���x`n��<�3�k+F����G�i���W���W�e���*�,z o�p1�g,�H7�Z�9�۽�rΌq�V������4̢����~״E@t|z�̲�s��]����O[��6Yl���@������cDk��o��SV�F�E��M����uM�}��Vf\ٙpۺ4a!x��k֧�x�4=ST8:���S>�m�ǽ���U{9v��ɪYobشw���4`d�.��り���9ڭ��n2r�?��������$���$��H@�XB��!$ I?�B���IO䄐�$��B��@�$��BH@�$�	' IKH@�z�$��	!I���$��	!I��$��	!I�!$ I4BH@���
�2�� ?8'N� ���9�>�]��<IE*�T�R���$JI*)J�))(Q)J�!ID*�@QHTJR��(T*IQ�BA"
�)�"��T���* ��B)U"HR���T����T���R"�HR�T��D�T��IH�QQ**P�6��åPUU ���*��T�RJ�JHE ��AT�IB�!�)%B�IRE�	QUIIUE*%
��R�$�
�  �`PK۩�իV�b�@�[`*�&U �V A�  f%�����@ �
-�j�D���%IE$�  7`$�D��*��F5�R���U�0�)�0Z5j� T� ����D�$$�I%TD�  �j��2��1H��Ұ�5Yj���z��V���̙���5�۬.�'Q����(Z�eJ�6*�l �(�TJ�PH%�  {�zlt�X��N�SV��%�
(;�0�P��
 �C9t �B�(P7kp�B�: �n��: P�B�
ꛅ
 �B���.�n(PP�B�
v��
+�p���$��UTQ*��Px  s��PQ���r��l�,�i�5��� �v6��S���Ҕf[c@����jt��*�gXR0ΎU!M��*�PD*�%Um��  dꚶi�cL����Iv�έ�:t8��+-��dc]5BT]�g]	]�N��a]*�uFi���nF��m�5�[J��j֚�R��(�P65!$�   ΁Ka��¸�&�ڦ��bYT�P�U�(����wwZ	��BSX[YeA�5��[V��j�����UJ�IA���(��  i��-`
��A�]�Ra��v;����PL���mqLt.R����2��k)5��1���t�3�Ӭ:n�Fҕ$�)*)��!Q�  ��E�%d�hlA��u�n�Kl�vҵ2�i�AѬ���@,qqV�V�L�UJ-�ƭ���2�[��	]�H(	J�T�"�   �(ӧKm�uݴ�����۶�jE.4�֨�*��3+��V�a�@������+h ��O 2��A�� Oh�J�SF@#O� 4�  E?�)� � 7��*��� $�DM�J���6j��UE(��9b�O)B�nT7��2�#�����CX�UV\`�#��z=�K����	!I�$ �BH@��	!I��IFI���=��������ssM�XM޻��S��j��KR�pZ��	M�i�)\��zU2��J4��b�fi�M<�t����x�CTNͨZ!�WL&��1�t�y�֥��0��`̏kb܎* ښ�5���R�`�f$6C�@Ԏ�V��KKpUn�i,��<"c`ޚz� ��,X�C!�iЙ*K��;[��*S;{x%d/Ztiҽ4�hZi�v1�9�ʚ�::LV��e�ό6��H ^�&7E�V V!6iNb���9T���5T�tR��f^�*Sn�T�)]�z�J{���VN�k0�,�W���QL�$fЏ�M�9�-1V����)�j�u����f)���
���Lւ�U�d�K�n�K���6�=Hbm"+���M����h�
i�V�ͥ[
��\�-��ۺ����r+Lݍ+e�\D.�u�N��,f֧%��e�"�$LMʰ��d{�Z���va�0���V`lR��9>crln�a,�(I6�{5InVEYřV��=�7�%Ϳ��P�N�����i������@�N���;G!v��.���Pm�I��j�,��5e"�b��x~���nl���EX)����%=�ƫ�m�3NEz�в	ȘE�d�)���(����uxƀ3F�Ykdլ���-�3�3v�w#L1z�ׇ*Iؠ�K��!eY�+b�Mވ��v�v�C5��!e]c����f������v�l�j֬�E��ACu�h��'��u�-$4�1�@���K�QQ��Q��%��^<U�Y��`�����B�eI��+ܫ�f�j���]޹�J�))[�1�m�{j�q��Ț �r�[cVm<�Jsn��ȱ����b�{�S�����Ö�D"��V�P�%�(�0�f*z�I��VF����B��7�7�	ا��dT�md�7)[\ �^X�H�E�_\9�������G��G�\�jj3G�SB@C%���lйsH)d�zq���Z6��X�ym��{��a������,vޝ�4lL�-n�`�[�!NV��l��Z���^��xZ�1$6���n��TZ�[[�H�q`�VA(U�a-�zl5�v^�e=�+6:&&�ګ�sB��Oc��w�o.�n^���>�p��yc�o,]H~�	z��Zq-9��V%v HJ��ݕdQ������N4�����e�-\B�ܛ��ՅYCNZ��ٰi�DR*mZ	Q��W"�c4���p2`n��S2\��eH�n������ͷt�n��^ˬ�]�m�PyX�v�;�^�l*�m:SV[���M�h��ا���Ȯ
�\�:��xn;'UC1�v$Ĩ*1�w����heB�kj���(�ZdsZtܥ`��b���x7w��˳��i�iE�).���D�<1�Uy�K��+�9k@�c�2:KE)_i�fnf^��ml�ֿ�nӏi[4��2'*�9�^]:Z�=?lf�w^ف6���Oq�1�70�	�d��ٽV���K��ʱ62A�`&;LV��*EeZ�4Z�{v 0�њ��\��+,�y&P3�W��f�Ѷ���X1�¡�Vf��.���)֪��i�JA���
 sp��v�u$��U���V�GVNնV��a+0<�wzO��N��حtjd�jݺB_L�J]c[X�jˍd���NnMR�X֨�*T��Ƴ7kC!((���-�=giG��T�G�mGDư<E����аխ�QQ�-̈́�5kN��6e�j�Vt=����j���K�r�]ᠷ�ʌYzY�ZH'��ـ�`̡�����@1�&����iJ�I��Y,��ɉ��Z�� T�LM��Y+�ystS�.EZ�Eb�.,:�#]��k�" Jq��ߞ���X ��Um���C�EMU��tw0�N7���V�n]�h��*�m*�ѓCn�gہ�A��Vh��� �؃���ũ{����M��:(L���u1��B-�/��p��n�Q�6�l���Zn�k$����ʺ�;D�2,�J����w���c)��G3nn�.��ͬM�9H�������v��f�Yl�P�ȃ����m��[�4�z�2oT�n�6��������eh�^���ٻi���sp!�Jæ^b˩��v=���R+;�U;U���2����t���Y�#Y�\�l9J%jX�4����L�*^]�j�"��@y��kߊ�F��S��u���v�5b[[kj�Md��-���Z9*��n,leU�̔6�b�Mq�K��w�F\@���$�i�V9�nx�aI�w���Zm�)g�G�V�+���t�(�%�n���8�j�ۣ�Ph�δ��d�c�1+���ZA�G\ujm�N' /.�ۺ�?�n<��% �.�+q쵙0%(��j�A�ֽ�C�7wd�P�k���=��B��@K�a�|�bZ�I�̫qPG2�{�جT6�n�`! Y{>������jf��HX��U�+��@6��cڗ��DDݾ���Nw)-�X��m,7��O�=�mf�CI��Y΢�j`r��+e�e݊����μ��l��-���nѭ3`�ɠRD��h���=7�Æ�M�wN�[WO+07z���� ۽II�we\��F��ڛ��e5��Z��M����z&� �*Tl��m�C�!lA�@% (FfAgm��؏6���yCe5q�lc�J���ׂ�#sYb�;-�c
4,�(�1���$V���n�{,��`�R1�B0R��L�K�I�1�M\$��T��AQ���&.�#������{�/O�V��rȹjA����f�yj<O6��ڔ)�x��I�B�͕��8f�9�Ț�I��F���N��c�tU�B/iI������7Y�K�(��yY@�@\�"��t5��躢ie*��JZ8���\�6e`�ri�6�xU�M�%�<9���`cp'�1�=���GS��[3FE��DK������-[���q�ZtM�Mm&�:5`��,�����p�XZ���0j�j���&^�]ZT���x��*�!]4�Pe�^A2(DsL�mJ��w�������!Sѵo@�tа#��O�*��I��L�,
80�km6�t� M�0����E�V�sob�Oc��m ��]!��z6U��a9y��*�ս�P��&h��j����N1���g�&�Q�/��16�WG@�l������Rbm�VY��;e��Xra�K۰]�aM����Z�I��-\A���f�v�#�]���ko^�:^:+3*�F�5`y&։Vs���݀���\&	z�&te4��sf6��]�pV^�V��dha����f��j�p]��K6�
���F.k��;�3oMmܙ�*C�l��yK)Q�љYu�|��Z*�.�B&ٷ�Ԅ��v�*�����A��mcû���)[Z�9A�2Vm����3kA��(�w�7%���9E0�I�� ���ucj`/�u��G��љ�t��u�B�[����RĬ��UJA�2�7-ho-�E�+pp�܈S�)2
ɢ���C���s�N��8pģ��$0���f� �e�n��[6ĺ`V:��7�a݊V-5�)�K`[�kN�᷹�ͺR1i� ���s)����oh�ٰ3s@�"튛/�<�����[L�h�Qѭ�*���ՕC_�*�W+St�
V�u�d��Gx���]��!Z�f1�`@'�0����7lE��h�����rە�֭՘������7���(%�J74*X���:��a�"!�f�XdLϷXU3#iF�d��N&���a�3ib�f�$̷Kwm����L���V	�I9z�8(n+� ̤���Rnl�4U�Cv`�n�x�4a����5w�d�����ؔN���z����y��eI"4� P0�������H-�mPW�e�p��2�:���@}�.��[M��
��l�D�DXH������D����WL[����`N�c�t���NJ0N�yX�Gj��V�u�[wy� �h�lPV�!�F�tkK9��4�d���k�]/.�o)P��f'EQ�ʚ��n���.��ŀ��2�@�w�ں7���mf
ժ�mi/q%��[�q��5�DaK�˼�j��I�%m�'2�QLf�tbۊ��1S�r��V��1��d���Zh�`���C0�n��������V77�i�3el1��L��lܧl��Y��b����{��úa�Ӹ�b@!��c7s2I�����H�b���n�w�����y��Z	�y��"��u���|b���l�ʼJ��0Z�@��З�s!�(e �隱���i�V܂K�o+wBN�z�����Rx�nb��c�W//nӔ�O��`�.j ��#��FR{wOH5u�⳶LY��zt �6��L����`A�E���Ĳ��-��ɂ�{Ʋ���^�9V�FC����Cg�t�ޚ�d 键���WC �5�i�����#c��YI0{Za�ͻ�%4��L���u�+����n�4�5Kb]��a,�(�Ɲ����%e���	d��42��a���\��Y]]Q�"����]��ֺ��c�m�u����By(�	�MV�ѹ.` ��n�6ېR@]㤴t���H��uY���ܬ�8Z*e,����x�
��6�ء�^�%.��h��ٙX��!R�)E��3��ݬL��7Yl����Qeh�x��4�(��0!h����1p��M��Ȇ;���
l��Yl� �`����b�hƃ5��N&5���ɩ��i��ޗ@ZZE��Nd [*F���8���'��&FY���l�t�5.V��5�����'��Z�(���Tv�B�c��G�VS�BB�r�[��P�-���+M#vn���*V�o���㯓�y�1��Um�P)qe��7t(ػ/���DCv�R�X�w!��;VŠ�Z���qI���j�T�^Ag��P��1�����:�{&.C(��l�ۧZ�1<&�\��ߝ֌c]1&H
���w�Fw^�	�,�b��z�[�\�i����I�Ҋһ���iDf��؁�5�#�6\���Z�T@�yte�2��ɕ�ի�&�IK�����Sx�4���v�	P��)�c��V�6���D������B�G �𵵒�;ʕ��I�N��R݁S�q�f��72XѴ�p�
כ� ��I�J�[b���i���S�3,��B��V��;i]��5p@.��wW�v�X[Ú�YZ�I&(�7�ƙm0�E����bڕ
5�t戦��sj9o�����X�~pLӗ��
dT"�VH��2m���f��*fDBwSF^0�,�8��z��	���Ŋ��I�&bծ�c�R��Hl�����ۏ6�p�um���! ��ߦ��-X�hTy��m�cT�F	��W�#;	u5 ա��c�2� b@�ݠmS���ySuޗ�m�f�/T�A��f&u�0f�%a.��%���i×w�+jP(Dr����G)+�1�ɶ,�hᔤ�4�*�����`Zn��Ui9h�1�E�,�ܮ+�>�V�3�eͪ�A��6+R�����x�E$U��0�i��JE��r��FԊ��q6����X���"�T�ת�$�H��7X�T��oj`͚"���d�T,�[�¼�&�6�m��a�&!a݋,�Dbz�@�.X�ѭ�r[n�۟$u;�i���B��F�e`�F *I�Y��� 6�82����vӋoQ�5U�`f��e]��[X��l�҂���Ȇ��(Jڂ'f��/A�� ��wz��X�vc�i�����%ެ��QPw�e56cM��5H[��г+@1�Lͺ������ccM�N�R�6��QV����]�4��U-7/U�wz�]I�^j{t�����	j��CM�V�oI��Ŝ=��B;�2�)��N��M���.��K��V�=J���l�r�Hf���5��f[��T�A-dۋ@Q\t+I�qyy�d��Z!OH�@ɏJ[h���*Cn���-S��PPn�Ҳ�(A���=�����b�>�r���e��M�Z][#��H��DB�`YX ��ko>l���#ud��Ҕ#���w��M����d�8բ�W�8�`�*�`1�Znh)ژ�	Ln��cن����CN�OB��e��M�kX�%�e�Cv��έq��H��Pl��lF��m�/oCX6HŌ��L�Ln?��BTN�hV��Cr�6��Ӗ����@醢�xj�c6�=��kj'�ġ(�Oc׎�Ec2�*7��\��CX
X�f;�I����b�Yf!��*$V������nݪ$%tJ��ڕn�jrB��Z�4��uzܫ�؍|H�2�	sD�Hk>Z��&���՚�W"���ʼ1�׺��:	�A�t�����uN��f�R��.L��!L;��ɪ
Y�IB�%��ӽ��X���J�C�(�#V�����6�̧dj���e��iO`���@<!U�Z0�Q0 (]
���TB��x�Չ	wV0?��u`!��%�����9%��r+�[��WX��G
���?,��a�N�H�Q+��*�cx���Ƕ�ډ,�X����F�&�����{�:YH*�FM;�3h[�J�&�%Vl`��]@m�eތ�օ�yhր:i�n�*�ͫȺ��/[A^e�7�U֗L$í8T��B�V؅9�0�������:��%�����[��0acL򫴉S�j�rH$w�q7yI����E��nC� �Am��Wt�ӕ;�GC�Ӯ]�`ff���Z)z�۱�'F��P^U��F��#����v��ڳ��VL�zڇ���i�C���aN��,��l�[�;��.��K�%͛3�A�ǬuλU�Z�9�St t�}�s�+�K�2����|{Z��ԇ9�a�W�q�WJum�Nn�a��ѦU]���ԃaT'eN�g��E�.�s�j����\��k����g��ڏ��"�f�h[hͨFWiSV�eYW��rpgQ�`W=��B�p�i^)�K�ԭ&���a�D;y݃L�� ����=�n���!�i��\a3�r��2��D�`�����ucP ��a�Ȟ����:�`�V��%���������m<{ǁ�/�����{RU�;P	��VK�s��g�3v���\��Tao{{N�a;�2�WmXN��f�X��>�D^Ev��6����mo�o����C��[��r�)�D���'�c��vm�ϐ"'��i�ڸ�r��B��J��zk�nw�}xUl�+xj끉��'q1��u􎶣�J;Zy�R�1mv!9��Q��
�Wي�R�ࠑwv�4n�k5sH:dv��+���i��9�8ć^�8���;v ��)V�R�|D�8��b�;�v�b�V �m���8��w��Uo+��֖ f��Ŭ#���2�ꕽw���ٓ �,%G��$Y���0G3�h�B�����K1 �*uio��evJ�2���gr8�؛����,[��	X����u�{���#iU[j�X�c�2���J,e�B[+r��NhsNeEX:�h����:iՈ�H�)w�n�8���x��
�^YW"|Z��S�f���rQ��s�<TH=�K3�8��he��v3tn��V7�T��AL:f�Y�����p��8��Fq9o�a�Z̮[�vdݩm���E+N(TƯ����	vx�nƱ*�-�]Iޕ�Z9ԳU`��Iu8$�K3�P�yN����#�FEg[B������
�4F
���.��'���A�{>�`͇����%d�4`grCP碅d�@2S��\���չ }du�@���%��.��q��vN.S'7vp�KV2���\ 
��o�5�2�]���?��3����mmM|O����6���yz�	wHpu���U���辝]ǯme��bq����J��:���9��oAD�e�a���l{g��h\T���&�W�u7B�[ܢ�6��+��)��I����� )J'�-�7F�8��6I�nY��4��j���t�� 趮��WO,�rX���1��b�]���<<.��-��{��Fޞzv00&.�M�=}�2T7n��Շen�sn5ϫ_p&��,��Z&���ܮ���\�{B�2�ZOBf���%��ī)��d�Z�{ׂ뮢��w.�v�@)���*AW�X;�]����vef�iU��Y��sZT+ph�Y���M%x��b+�C�͊hʕ�;OY���R�4ީa%8���Hp��Vk{��,n@f�
���gw�oSTM�SN�fm�&�]��Cm�s�Wj������[�H�Y*�#�{x��
�+P.Ds09�*ʼP�l�w��m�Xp�B�����ͫ���ޞ�W����N�y�<6���N�.�����`+l���N�LR-�oI;��p>Ι����*q�����N-�ˌS�^C��⠤�)��{i���f_�����(���ZI��ïEn5Y�A�h�]Ռ�TWϕ1��on*�ޠ�X1S5mq�9��E���|��Sy]�)n�M�d]1�W[ճ�&�LQ���8�V�K���7[m�R��] Mޅ!5�R�@X,l[��JO����g���toQ�z�Z�ޤ�Rh��W6���a�ȴ3���Z
f���燂�'�*%]�3�vWPB���Sä6*L�idg��(E��v�0-�G����\��쎰'.;{�/78!vա;/s�-��`uw��L�M7�l�L�|����Mi��.��,S�GZn�>��tkh0�>��l�`k__;s��٪PNrM���{�o�����R��U�	A�0�bY��t�s��@�E��,cwu��qz�<=e��'u���4,��9J�fv9��y�@�8���K&q�.-�EI���� ��m����I����R���uAp)����E�h�[.#&U���.�7��\��da��:3�J�v��I����l�]u��I3���l�n����.�T�f�N��y�x�T7��F�w>�DI�E�,��+!��r��#1�,*���vc���8ܮiJz��l'��S��'$+Ga�T�����<T@Yb�n�����̳�C�����u�<��P�7>~����Y0�7ʀ�ɞ{��p�����Yez������T�n^�+'�ʰI���"���,WYQtIŚ̷��NPu��
\׬&�RW�P��<��9�4���2�e�S��w97:-�w^�ز��s��cV�I#OH4�U��)|t�nkQ[��>�;Ere���j2¢�'Z9��X��Z��nwWV����E����]�sK�����]CW�-ٮ�JWL���zP�� �v�3����%aue�VBLwdS�����Vv���m'f\�[\yd2FJ\��vV�4��7��jޥ�r�g�Qp��fA(��
٩e�(7��82l���wE�W����Sp������"�xg]r
ZB�;��Q�6���Q{S�>��.�H����y#lj[�+����;W�+�*�B�\'��Q#��X� �Q��)�v��h��]մ�x_ڒ���@�
�>�]���j���WJ[�s��"��pR�؂
;��n��:,���w%N�PRw0���iB�ZƨR�ъ(����Q��St�~��wB���Ǯ2hu��a�I�\�Z㮮�k]4f5�,[ұ���z_QYǨ��k����JNeD���pG�m��i�Cs�ys|�Z��Y�ý8=��}�D������n����0���>�k#�z�={p\���vU���t;��֘�ve�/���f�D�k���nq���k.��}�a�g�л����3�8���z'P�h�v��b�yg�ȸ�WA=zqX�A��T"�-So\V�ٴ���/�o:Xɖ��EG�����0d��m&��8�=_^��6 ��j�F�e�
�O`$>�]�:���z^T�1Z�-,�ԇR"% @���V Z嵺�sw*i��j}a�x3^��'IQ{.c���vAm�or�E]���(��e�6�hNz�����\�_���:�T�n�c���
�Mm��_r�Й���d�=�*Or�aL�%�^n���؄��Z� ��&��z�l�`g,�����7ژ�כ&���8%�:ˉ��B\��0�'�͔t�aR�O,f�����Գmm,�i��Y防,��Qm f��M�����\(�]j��	t����䅦C'1Ŷ�	�n8+��[�:�v�G���XƶE �t�s�B½���Wd\2�T���s��M�!�L�6�f�V�0��:���*<�3:��j�[���=�/�Y�bݲ�=W�
3&�ή�_E�M'��Zݲ�;�xbWC"��o\̴�����J�5���QK��ݾ!e�E�m���'�c�Ac��8Xc��[n�IZ̋�WBe�Mi��!K���.���$���c@zU�t�RV��а�mm܆Kj�vZ�i�W/��>�y���N��֎@v�¨�)|]�[s��~P�e�3���	#6�ژ�9�'q�'�rE�]�[�j�=%a"v�E^�r*]�$�K$�Y���]�Դ�ya|��Ҡ�%b��ط�(6�!�����8)��4�_C�!k�dfw0��)�����l���'F�.n��rt�%8(����*\{��P�y��d{ϫ��D��ەs�j]-�҈�}k,���z&:�LJh����}�u�;7��`�U+��op�L�}ΙdT�muݴ�XB��	YޜKy����]p\69lfe�,��h�:N�ִgV������M����	8�>����������u �m��v/li�����t�n'i���C�~!�N�M�-�' V�����m�s�u��6
�'�9���QI�ק��#8�Y�`��KQ7��j�;	$+R���r7�=]B���;����2��7�G
��]��pt�}Z�%�f�1�^Vk2z�[���e��r�a��=\����&��Y�	wɥ]�)���d�qֱQ�Vd�fb�6#��\ˢ�5
��"�ɷ�:�:ڙ�<���ǭ���%�{��I�K�n�.�鐮tT靲޹��͡���=R#�ٜ�N��U�0;9l�V�}�u��KZ���ۤ2�N���y�j�!�B�![��/h����L�[��F���T��,=��72�7�NK}8n;�z�͹�61�'c�t����'}J�f7C�m�y7!�s��.wrR�D��#�K%`�+t��\Ω(�;��uLm�i�	S�V���R��f�}(^�=iܫ�}ܬ��TШ�oR`�"B���o��V�wX�V�ܣ��� T���ȷ�v"��)��)�l;�S19}���ґ߉w]������ҙ��+KOD��X���lV'��`�1�E�tOs9��=90kao�<l�Y%�CV�@�Q�fc�6>�˩X�[ �Qc��7�CK��.�1Z&S�Xm�)O�.��a��X��|uH$ͽ��C���rC��:}L_	�?-w�V�eGybpV�R�,K�;J��5�^����[�].�����}5u�YI<w�Ae��*�T8���hY9բw�nJyd�]���[����&p�Ć��Y�xaeWJv�U˞W@ �L<U�×��Y2�����ƕ��g�p�JMX�\q����������v^�� �yVv,�9�Q���*У9v5��of���)Q̚ŵ{Eu뱃���׽{�YY��/gw�vmh��'X���>ht4puKaܭ&Euݡ^йx;Bv�\X����2��gan�Ä�����@J�I]S��O;�H��a�,���G��*�Y���LɊ��B�QZ��� â�u)VZmT�L����:j�7/R�e�o��s��[7�(�JJ=� �K%��+�b���;�����fo�A}3�ע���ض�ރb<(���L�;����Q|NH�wq
�s,����{�V�X׆O�̾��5���]���ҳ����-�`�N����R�+u�]�'c���u������h4·�k'(\D�Q���$����]yjS3�f�EYz�e%v�m�����*��묀4�Mo��oo�[)
��K�C.bx����\��2���Fu%�k���Y��!mK�CNA��k�3^��7Q9�K���1%m��n�4Z;tW!���/W����'�(�^���WV��s<9��H��y��	.���k^�֍�Q���I]Ղ��]�[%v�����ճ�R����%���(�4�p�-����N�ov�`#K��&�Vl�'M]�J0��uc��j޶{U򅡨`�s�T�o]��cij0����]4�KX$�.�{������u!w���jm�2g}L����ɝW�Z�kNoZ��2�a4�NC���Æ����ϩ�#�/�g;s~�7n�Y��E���/X
�����k���ܒ��d�t�ş��+�u�I���
��HMfVM�t
o
�8�]kg۳m-��ҷ0Z����Gh�X�i��]k-U�{tz���k��4�|��v.v�E�Z��^�]����p�V���s�X§V��w;"�t{��hW"V��H.t��MY��Xy~�ڻ�b����'d��z7�aD�Jh�X���sݢA�a\�B��kg5��^��Sʻu�5�K5�� ��Z�V%��]*�*6e��:�������ۺJ>�(U���p+����Cz���P�F�X"be�s�U�]u�m�� �|tu�=�g�J��&��y�)�kʇ2�A�V"�����m��[?Ej����ﷺ����oi�s2��ۭ�?$������}��X���\7:�Z�|jn>����3������'���sE�JM��2;`Z�a�S��n�bdɘ�[7^���`��X�l��D
�8W���-0��M��dovm����:�Đ�<���qC�<˥:�nK�ϖ�\�K2��칸8�Ú���7���%=�b^o��ס�v6���t�X9����,:]I�ʍa{���b�����(Pq�kv<s(sa�'6��a��A�-����O��" Џf	.���B&��Oii�J%>�xk�D�Y�ɩ��)���uݖr�;:+o76�7I�E.�*X�����`�q"���S@ KZ�7|%��x��J�9���f�e��uC٫�l�b�
E� !V`
��Ղ���RT������L�Tt�����uْ�Y����\��X/TdS��<Y"��:�^�ε��h:s��Ύ�������y3e��o."���k:]پ�W3���ɀM�'�k�ut��gm�T �Mf�$�/���k6}G�N�}���9��J+�jJ�@V���d��T݃g�?S�t�CFAs{x�� �����bM)]]ݽ�y]|
Q������P\��9�tJ�n���mE�E9u���.5��u�&�^�C��咗Fz`%1����V�.��$b����]ݕ�t嶪�mꤋ�����\��Ş��=jf��S��p�fe�9�So����%[[������foy������z=�{�����|*��ٕbj��}�n��)��=�b�#0�Vb������.Υpd�;Ϸ�%s�`�+숣`��ѡQ_f5�o0��]Qi�v�u���ҫ��]�.��`R���PO���ػ7I�� ��ǎn`�6���w�]��h��x���6�"���U�
'�#�=�ȡr4t�[0���yJ�BGZ��ոF���e:�H+�۸yЋ�P�2ɚml�Pօ�m6�d���*!��]�q��]�D����82�����q�f�V�m��S(*�J^A(L����)n�r�����Q�"t�H���u%G��Δ�8�-�ΆoN�x�;rpǨ�+o4WM�8:X4���͙���l`���ƨ�J9F��]�L����q��N�MV���ԥq�WY#�]�<f�o+evL�;������7�*���<���˛���_[���>��9Z5zp�_K�J��g]�}�ѥ�Z:�#a��\tN�[�wʕ2�
�y@�
�:�6�쾫�gmuv�I���_V��� �/��7@�`�[S:�u������Ql��D��ܟ���I
8+C���F���v��#Sv��h݁�]�����f�Sx(i<��K@���Qԭ-	إ�����CX��8l���`m���OSfệK\Ge-�Pbv��Υ����
�	*XVv옰����2�t���6� YQ2VYh[d�5\QT�+t�b�iJ�5���x��A�a��ZQ�5���W�#�.v����k)pu��p<�Z�-Q�'Z*�ʓMZ��+^U��4�	�,�ΐ9o{�۹5oӴ^��Oy��]'��q�dX��M��q�xBu��q��y�I�2�su'V\����<�����k�oL2�3^�h<�Y�������}Ǖ3��da����]�w\a��U7]oZ�P��=���9^%1���5���]���YH�55�F�+��a*T�;����V���c�y�����,��tFU��x�e�y;2���*►B�HAO(�8f.T�9ES׋K1�B�N;;V�U��=�Q鐞�}��jhǨ�*+#�O]u�t�Z��m%�`��w��'�wT�7H�C�d��p��qVa=x�n�I3o#����l#Զp�2GR$�|�V�FWT�ܽOi֩����(d��	T3۪췼�:�a���e�1�ܵ]�*�ˋ�N9ـ6�fV�5��Z��YG] ,��܅l��ac�Eхhf.X6(s+x\4�o���3��n�BU�Eu��=�K7Sz�jJ��W�/�\���綱*k��$�ӚbЋu��w���Ӻz� ���Q�.��"�w��y��[��(~�Q��ℷK����ŗ��[�LF�O�����̣��t���jy�p!��r�ζa��w��<���6�U�U�[:WX��9[���rюh�3}ϫ7��eVV�5n������r=�o�L��{|�j������!ެ@������(�A�e�ɜ۠��4�<-��^�8 �Cv�M��P��mYƜ��ܳ�f&�F�j�zGfTl�Lrm�Տ����Z�M���:����/�����l��v�{���2��ߜ�%#�\�j5Cxj4�>J���d�7�Kr�����N�q�R��/[�I���̶hj���CRG�=�bV��Z�
L:�T��0�!�����SS�3G*Iw���ǌR�']pV��ݺW}�<YZ�*;ڨ\�U���1�2-�9T;�+�әY��g�)#o��j-��܂јjQ�V\z�ėi�I�aj]:=%���ޡ [˔8�ޥ}����� D���6��x4n-H
�OR�r<�r���)���hN;�V���"��<���R�4�T0�qu�C�Y�V��d��R��@���S���t��e�����6�]/q�Q7���*e\�6����Q[�sv:g�:��A�&�u{O[u;���$6���*�9JX8�^�}�	��rw�SC%St�:�`���������`ƻU��ں���WGi�\�$���P���JԵ���xP�ނ���H�D���_uE����.mf�7u��@˦�\.)sg	*��C��Qd��K ��s4�t�u^S�#T���Nq�9�W:��^j�\Zs&lu�
������q����ﮌXfl��'�p�N4�p�܊���{�/&��%Nk�w�a�!(PN��6�mN��8g.v��^{p�B�.�̏7�=zȺ��s�u%�]���|�4T�j��2���r��u(��|I�i�*�T�C����Vʏ`��hm��sm��)��N�)�^H����_̭��+"�T�2+i_3ׄu�圉�ŕ�Q��}[N��+�qr���m<�..Ρ�÷)�a���{i:�Yس-*��#w�y�?*M���5����
#zmk)��o�X���0���ĸ7����<)pw ��:\�tv��:;���E�D�C��g6�`�vC�$��y��FglQcEJ�رWcݓ:z4�q���(4.А����0�2�;1�@�_X'J\�����"a�G0% !�BՑ k�9:Dn�Ngn�ѾH�H�Gh�8����Ƅ��TUgX�-<�i}�0���t[y�Q��!�i�$w�������݁��jۂM������t$�뢫�G���J�0��;�mSµ��J*�/T���<���cUeu���֥��Hz��e�wY�(�fV�M�:=�w�@K{�V��,`�����+�ުZA�E��g���ve���Z�3^W$ͽ��ؾ뮧JRS"Z�KNU��q^��7
������U��t�T��N��n�d�Gh��M_�0D
�no�{����	�<-r�h�]j.*z�R�fά����xn���'�i�}6.s6cW�|�������;�4m>��Bɗ�I#��#��.P9t�sR�m�~h.���F�#R�Һ�w�@�y�����Q�w\�����,��$�`M������H�ֹ
���;e�smOG
}׶�PB�cz�+����nF��=�.	�d���,e[%ꤦ��v��Cw�v���ɪ=����cJm���c��(������*�(A�b���nP��uYSmB��uL�ƶ����T�{η��,gb�r��k�T�,��LO�sw�n3����5�Z:�J\�`�!�}2H5�����q<SC���3������;�-	��iD��XXx EWR�6�䮏���ó.)n�7A������U��e*Hw|`�}�K�v�3�����f�,���m����bgby�F��ѳY``�z(*�Dю��X�w��5���F�Hv]��; ����m�֒�v���\��u��ڝ����.���n>�G�j1_e�`o(D���:m��w�71��}���4�4�4�$��	��S8��k��`U�L� ��@����G3/w�L�.,:N�l���Q(�+qt���9n���\z����p���:���v������>b1t*�)�yE�+�'E���j��k���e)=Z9�5%y��d8��|��#a��]α��1�-ٍ�mp����P7�K̤��A!���B
F����nv��vN�q�{op#��c���5���։-��;%Kc]�oVn�f�Iκ	�M0IЩށ�Gvn�
�H�;y�E%�6�\ڛ�	���S�Y�eh��L�Q(�!�ټ S���!�7S5�t�Uf��`"Z�Fi�о�y+�!�ߖ�zXfT�[ݸґ���cS�1l�;C�j�t,]�z���Q=]Hs��<�'�e
�q��X0.��l�s� \-�9,�K$޹��aU/;�v3F�s��bKT[˓ &�}���z(��W����f1�#�^�z��}���;�;��L!����r��Fe_-I�����-� �V6��[�X��A���iCome�;՟K���F��g>C�]�$j+��;��^�[��˻fc�{8��M�T%��L1Tau8:����o(q��[���ggC�R�Y�_ۗ��͸U8,ZH_q�é���oFϦ1�{Y��ީY�\S�0"�b���q6%��������$�s�X���K{RӾ��O��2�mJ!ξ��E�v�Y���V��-�@A<�*�W^��֚n���y+\�E�t�1{\�p��"����أw�C*,�O~��iV��r')�d+�	n�@��pZ�NU�Y��Dm��a&��s�aN�A��2�T��4�T�,ry����Ķ�p�t`i��rlu�q�Y�J����QL�2U���)%M�!v�ݳt�^owbf�Mn���[任D)�!�&wU�a.Q��L��rXw����35�;{Kk�b\#F���}��Y�*��Ц�5(ؾCf�e�F�t�c�5�S�G]l H��DjF�Bۭיqvut�5]��s�֩�Ȭ��e'���g_bWj���m�o�Lf��r���Z۔��6tѮ�L����.���ʹ�ڸVR��j�(�:7n��t�̕��U�ᣑdM�j`�Su'�h���]��tr#\�"�y�O��k���YVGب�����,]���]�ܱ��.�EZ��).���IYs���"gc�"���	�ls�^��6�G���Ov�����S�����r�z'|��ʹ;�c�+NY��0a�J>}S�V4Χv=-��b��Ч�ø�Z��<((	��@�ވ�C�4���ՃTB'u�kMʽ�7\���JK���F���Ψ�}8�1s���_.�u3'[�}�Ì�z6��2,�T�n����FgL�W�'�p��2���i�9*��
�{��d��L/�>��kQRd�$�Okm9y��z���gq��ku�3v���r�J��_ZlfȧX)�c&b΀�ee
�热����X�9�^sN��ά�G[7C���durv[̂Z� ��-��6�VCz�G�m��]8f��R3N8k����[�G��[��n9�R�ؾ��l�$ۀ�5O�S��7l�v�e��hE�]��Xy Xۺ����-i�:���x����K�E��+(+ ܗ�KN���7,G�w8���<J�e��s��J+�㔀כ��¦t�o�ѵ�h�WsJU�{�ևs�+���F��Sc�t�S�R렵�+q\o��(�-�,Z�t5;r�!�YV�+*:0s� �n��)q?�G������n��J!�v�:/�pe�)�Z���O/3%KU{���0���,�����{�d�����}cX�}�+<;o�Ր�/�̀l�Ѣ�׌�w�)()�C@-�G��L��H���)[sAEm#y9��]���Z���H��w�ֻߒͰ�/u��D�loSh�rfkf��P�F�����y\T��D'[����*�*3��%��o`��ݱ��l��b\7uΊ��9�A$];�3�+b��v����W��4��	�vf�A�c�(��sw. �-��������<��r��wm� �&^ޞ�*�����"�A\�.h�.޽r�:�H��w�Y��������B�d$Զ��/�t��|OX�n`� �R1Yb����[J��r��o- ����CA2�\�ӳ�	>a�Z��
����c�l}���'2�v��l��*�@t�Nb��i:۬T>}qj�M6�2re�z���n�C��OE��C�F��!z>�yE}��4z9wn�G+�M�XL���Z��(��2�&:d�t�k�-J��K�#���u`��=jT�;&��j)g����]1ݫ��zR�젦��6<z-�����s r<��B:d�]���FV����2Z��c4pkDӼ�F��:p&k����vS��M.��&<=�Z���Z��]cQ��V�2��M�Wg',�)gs(,r�Z��=�df�:eR�7,�7[�Z��q�7G�0�-�(�M�K_�9��w�f�{m���y�H�wܶ ��)3���0���57�y�#Ƹ ��ˮ@��WI"�tt��p��:�}� V��}JWJ7����E�)��+��U��Q[�|�&�V)vĹ�+t.T{ "�����J;xv���[Ԡk��E�u�X����H�[�rv�gD՝\��U���h8���f�����VP��]�4��6�*`�gU��Z��0L�VӐ=�pa�'P���[05o�&=���b�pB��]��櫛�y�N��}�V+:�H����`=�(T�:*����Y��uZu/��\�w���}�t�aY$D�)]אLљV��{�Ӡw�ޝ��9�"�K�>@�u�s[��$����6]���	��wd�[̕(���MP�m�Ax뮮sW6�uh坸07� ZU����6����Y�[�v�c�J%k>�t��I�:Ѻ�i�.�@�V�-pq�S��j�#��[�6�ݴ��!G{���6X�2�4z���Z��Fm�aYf�i�O@Վ�:U�-�\0u#���HI8W]Z	q�ol���A�36���ȋ��ي�U�i��ˇ,l���b�GRvgn]�BBC�L=G2ث�����g��cUoN.����bg1O�K��l����.��#7@PV��1�v�I�mr30N�Ѵ���ի���Dl�+ŉi��rW:b��L�!���n�<��Z10+Hȍ�֑�+,�Q����B�}����P�l����Gj�)����%,�F�%�U��B���������Z�<�����4ƀ���
�Z2YL�R�l����	�I��
�n�7��� �,��.����ז��n��$�x�ڏ�LX��*�u�u�o�o7���7����5�r���a{�0;��k�t�7��)�B������c�.���
9�LF����"�L��]�q��1% ��0C�Z�ܻ���*.�@��&L�8'\�@L��@b�\�<��{]��Rz%5w=�V�o(S꿌�۠/e9H�zY��sRĳ�Y9����d{����ߑC\�rU��^���5S�N��T�
�Xt������G��{h�����)jĬn(5���N��J�ù/���ٙ��R鰒���4Α����R�8Y��*�+z��	��H��u} �{�vܜ쮭��[]-����8nW�V�j/5w)�f��A7*B��xH�&䶊�֬sV���.��vF�\;Iїa���F^�b��
�(���GF��V���_d�Ԧ�ۢ��W%c�#�uc(m 'V�iV��Nqܺo� Ek�t����*3DTn�L3�Gin\Rn ār��q]FE��������wd�B�Q�ʓd/�.�Lͩ��mN�5�37��`f�G0��Y28�_M;[��Ù�k�u���G�1>�2s����?Y�ޥ6���#�t��\+r��Jz,��/�3���Z��)�;�V��X�u�/MyչmZ%��Yu�w�6D�`�1��T�w��kr�nu�(㻲B����Պ�b�U<En$��,W��t�Z�A�� G� G�Ll�UF�H��X���-J�Dj�DU�bɖPQAQrʊ,Q�������"�cZ,`�**�f%��1e�r�0QEAV�Z�jUDDH�Q`Ŋ�J�
9m�UĢbUA�TQaV�ժ��bU�Eb�PTU���3jF"
�j�PaZ(��(��bEXj�Q*�����
(�j֡Qբ�Kh�Q.f+IAU��5QD�E��"Ƞ���J�b"S�"�i,Q�����QEb
"�U+R��UUB0Qb�`�,bkT�V�1b�%"�"�4�լDƠ�"�b(���(��q,`��խڨ� �e�Q��0�"1F**VQU��e�����(�e��i�UDU5J��fauk����(�2"i�"�DF.�T�����K�(�S5CH�q�D�U�V��+1�,RVQD�Ӆ�3V�b�*+$4$ g��h�[��نq۽˽�JË3�$k��HG�Ѯ����oV���v&�3w.!:�1wu*Y�����v�[)t|�8m�]/��֬�����t�_R��&w^�r��K���\q�H��w���E{��{� �V�-{U��+R���W�V�b7*Pd���O5�j�%Erq�zj�P���=���N�yV���5�p�B�u2�rd�u=�込�B{���T*Kb�����*��n����:����|�Y��Tb�"�ڂ��X�[��	B�S�o�mOm�u���)ӄ�&���s�|��wٷ�&� ,R�L%^#5;����p���_5Xx?lTZk1t��z�o;|2^+V9W�l���oR;����XU���]�.w~�}1Y��1���bFm��z��]ںj�'	���lɝF��JgRt�m_B��dO�X��h7�+�{|�7��G�(�o��l�ٕ��W[�_��bw�[�[�O���U��-]y�ׁJ�P�/�:4� �2��T�6܆�1���w�;�^D�P9K��si�HFNZ����$��W9R���e)���0m:����[= w`�*p��֭Q;մr~��3�^�jFW�n����>�\H��H�ٵ��7�ӽܣj�2��e��.k��!|��C�����Ҽ��G�Y�t�H;7�:�u&�f��@��hԦ��
�>��x�__�^]L���MZ3��9���bs�K�n7�C�'t�7�TL�gH�KW!J�m��U*��eW�2g�⣭1^\������r�%%�;�琓Ɯvnub�usq\VeU��Q�Jc����7*��}���s�iw�2��q��_�k�o��>��Y�z���k�X�v�����Fz_T��O|���l����Y��]��Ț�����m�Au[ýyy��-�m��\�:��^(�{Ӳ�ku�vJ�v�r�>VR�g�ۃ3�ZO'�"�;P�z�<�+��;�c�l�n^
��ְ�3���4VT���Cױ|�z.S�ڌP󭷵;u�clv�C���Z�{��,q�H]����*-Yy��n��m��{��3��Ͷ�U�x��+�f����Z΁X�	fE�A�o ��)3po;��\���.�k\|�Rsլc����9�)
̓h;c����|�J}{���䱨�|���r=;�+:*��_��{!���,�q��o��s�K��"w��9cNmp�mUR窆Bw�n��*�hJ�t*�=b���\�Mf��s�5y�V��㯥��oφK�sP��Qq_m�;~:��ﶺj���I��)��|Sלs�����y
����
�9j���Y2����߂�ȍ��]��1nݞ��l'1�C�g�����Lpߊ�z�!���8���S]5t;��Ř�
��lJ��%ג���èF��=��3�t�F���|�vQ�u;��s��lgE�&q9�ĩ�!�H9�r�C3Eͣ�����VUk�"b��J_e��Tݬ�ǏI�Q���S��0q"�����l����X��WF�a�p6�
���c��y�[��í���N2�I&���,��o�>c��)��]�c@�����rb�^3����7$���X�L!�Y�W,4�V�n�u]8��W�����E�?P��[��zŨ�EPڰ�L6$�t��ؖ�a���1QZ�7]��{�H�.��\��sXh1F�).[�L�����z��jum%���(��X��c��[�uU'�:��'ڐ�M�x�9��<��f�|f�i�Zt䚕`����pqҺ8��:�9�\�Z�I��׽6�.�>�V�*BXNw9�=zv��f;�5`u<�N�'�G)U�S��j�@ZRH���WMRVi'�Ů{�]�Ц��OY�ݧ'��>}�}VtזH��������
�5�Ѻ��WZ��N�p�5
�CZ8��=���6Yww���%��ZΧ٪�<����ݸV�w��U��=��^�*7^�N�#6���%?ot�f��w�F��%⹤�ʸ��P�*�p� ,����%i�Y�Lں��>��Q9Π��n��l�B�S�H\V���S�e�LU,6]E����Zʀ����l�OA�ٲ�;����(�)���B6Q���
�/�=�y[�f�UK����)�v?M���\�7�/�i-JKV��tޗ;�"���U���l�[����Y.ȅf5�ND���F��D�U� �V+�!̢��Z�wf�\]��
�F��gR��Fkܒ����ͨ �9Y��Qk�Ġ��	o�R�;k.V褒�j;uXK�9��.:��>I���oko��g����I{Xlz��84_>ﾧl���Μ�;�8D������Wa>��L�֦;��7��}�'h��p��{�LR���v���J��s���ܛ���O�剗���i:YU�KMDk�-�SCaps���sÕ怽��U,��^s�b�̛�륕Qn1׵�N��1�U�����q�0���Ӗ��k0c����猛�Wq�ZŬ�jB|��P�h�N���:}υ���B��������_�g٣��k�)d�����U���/g;�H
}-ô� ������1���+sVS��K�d�lV=�Sf^�����X�����=YޅԴ,S��O�W���.��U}����*��=�h;��.WW=Z��<��k[P[�
Ԭ�/:���Yn����-��\���=��w@U�J��Y��Pbe��,���R��N��6��?@X������I+x_��(t(��ʻ�k\e�[}[��ݔ���Y�t�k|M��M�ZU�@<�P	�R7�>Ϋ[��]�]��:s�A��g��,���]3�x�9�b�����q"k�x\͵�d���?�<:�_]�����b�Uzs$����r��I�{���%�r?F+3
��E�mW�qUu�U�[��l�=��\qY�4�ӛA*��*;.\����Up��[<	]��u[�M�]��9w|v�fK����z���o\�N˾�'dLRc�}@嫇[�F;��� c'p_!Y��]2�ej�����P��~st��&#�+/��;M:ُ�g��|�W2���^gg����';T��n*!hiԼG�i�9�"E�.N����a:��[�̪�ɘ�P}��u&5pw��8���f'm.��]o9QTkl���@Q�αyjn�F=y���:NM��n�V��Ȏ���gT>0. ��+N�[vA���o���ջλ`����26=W���K-�rb���f;�- V*��&.����d^WL�6`�M�s������%��;g���yw.GE�1�Z��l=H��rut���z�T�#�AϷl麃��-��g%݇�ݞ���8!kz� 43����Աto�7���rw_��	�M�<]�^tҳ|�<͵4E��;�Jn�n�ԩ�.	�`rg���8�9Z�TB��ս�K6��zz��F���w�V뀓k���� ��I*�O:�*�1<��Վ�׊�ıN��}3bQٮ�:��S�.(���օz�*��u�UG�vW�Cζޣz]�����7iͮ&�1��uB��P�k.1t�<u�z$m�a�3ӮDLɍ[bW[H�kf�����X�_����:9�_]���=#V����'6�y@Ui��m�6�d��sI˕5��+n��(Q\-U�u��5��}�r��5��:���'����Hpe���/j���\L��U�:������{�vuQ�ٸ.�;"}I�7l�����,��{�%UK�o:���]��d�c��cbT��)�9�q��vj���ӷ�BF���쭇��Uf�6��Ֆ߳՛�1lWy���i�����U�*�}���uu+�+�TRI�0�z^�`�'=�fdrK� L`:z�mw3��h�+{��AR��p��.4�ǒ}L0x�>�[b�n��Q�}϶����Ǌ<G�����kJ����U�<�]��;*��ƚ���e��ƫZ,s���,���u_e��Pݬ�Vc�Ǥ�(z�n��K��[��[��C�/B�N��y�m�w��?o�5؎k�(eP��s�S�]��m��!�b㭡^\�;�\��V-���N�v0��^��T��P��!��SX&Ԭ�ؾ~�1�H)n�U��㽗9��sZ֬3s/n�b���֢��d�����*�s�И\�Z�T��$�$۸Fna;�;�B���?䟆j�_��:��U�Tcx�u���>��ݽT2S:��;ьuPV���!����G'�s�d#S�����	��<�m�]K`,S�Þ��*S�_
��Xr��Ե\�v�6�w��o5���:����n��,R��a*��:S�9:=��m1uz1xgk��S��\��֢�����0���E�[G�c¬�]S56�ݺ��ܦ7w	����఑P!(#ܣ�]���j�;��i��+��(�v�ÝϝL�)��{2����N��"Xk�����C���9�hә:�&���0��t�M�����I�_7��}5����J7���ɇ��2�[��AR�RY����yո�7/z�}�q��Vj���E=�p��P��3վ��(l�i�B��S�����߾��u(V���Wo+���U��ק:�Ǔfsj�6��N�+�j-�՘�Hp�+�=�y[�\U��by�\�bWh�km�gy�4�T+E>��z_ҥ��G��11¢e����1��熆mB��-ݧ̡�:&��Вu��8DƸa��vՉ�Ű�e)qs3y;��'|ɘƧj�q	���wN�7Z�u׊��3�O4t*����^��k�UGYڵu�Uk�׵A�������9���yd]�ڊĘ��@e8��/'�)�Z�{�q��LJ��v�O��d�*���l���U+�m�Om��
x��WGDZ�Z�+ڐ�Te��:M)���_T�Þ
mr��*w��ي�&[G��%'��U+���z���r�Sg#b��J�}�����+�Cq#�����\[�����@�_<��o����z�t����4um�I��Ւ1�����8*è_nd(��`�>�d,��.;�ʛ��c4��mBq��������ƫB���yST7*uh0�ӛ��>32��R��:����=���:�+J��׉�q��w���[8���$7���TޭN����t�-�Qb��㪢P��S\4D�8u��%Vv��;���z�ov(y��kjv�,R�cYv_���#.$d��(�=^��U[�ڙ׶Z���it�En*�{أy��������O��I���4��Ε�<D:�௮�.w~����s$y��H]ʑn�!��c�Z��FW�~�{��Pv�Hq�=o��2��g������z��}�u8�X�M��+����1�V�
�]A�u�¦�I�:E�T�،��]7��EM�r�)��e����Lp�/�e"��ޫ��L��3��RX����u�&6%LG1.�)M����<�Xb*a���C2:/qؕWL�O&��Τ�k^>,�J1�%m�iX�IΨT�L�iĪ�9��/v-�f�or�U:��n���u��fu5۝���EoR���C/Z��}��`S����qN4A���T�պp�P̚�*Ŋ���Þ�^��(��T���uf��l�H	+e�0�+o+���+M"a��6����!��#���n�e*n�9�>�y߂�-������T1�Nl��x:�N���b �=�ut�T�f��c���eB�[Hm��>F>}�>�l���y�r�#]',�h�����9���A�X��=�.M��8U��Dr-��S�&����I�W�y��&ܡ��Ɯ�[[��	��y�G��]y#b%�Ik݉F|3��Y�{Tk���ɖ�<ُo\5 ��W�]�ȱ����x���]�[�p%'ڣg�����n,��%�k-������X�ha�ƙ����&�v����E�:YX�Y��Ư��a>ES6i��݂�Mi.���HΑM��\���j
��Ԏ�Ν�W+o+AY��n�G_N��������ǋ�nnZ��T(�6qE,������+/�E��q��
6�r*���"�4����+�`���db�eF���|�;��;���!b�d=��#(��I�h=U��]ڎF������:�9����̦���wS�_�Q�:�b��g�w.0���Ӫf=��M�U#���;	�IW�z���l��7Ѵ�aq��90o7m뢱uЛ:S�!�!}S�K&�?F���w�.y���OPL�sD���f��q�*�9n�QȮn��̫t���dI�f��@c1��}��;Z�'kuN�Ft&ĺ�zi��Ս��� �я����.{q�}9�J�Jx��8fi�¥�e��}�rdk8�8��mk��6
�y7r��������]7-*��$�m���B�I�>`r�X�1y��Zς]n�q��C1ԗX�C����*�^>6�h�-P�lX��̣WVT�xtv�����]��u�����}8�Y*Î���p0q��tT��Z5^]i�֞�һ�󹧶$�e��>�˚B^KP���2��U-��U���S�Y����v���5>=A�QJ�m��7��ɉ��Y܀l��9mobB�c*uԻ�0p��x�'Z�PJh�˥!��絸Yg3�a
�Ϸ�ŦH��L36��gD:��Ah:n�o)t?_q[B�gEl���xBj
�h��H3Su��@"jĬ	;W�  ��Wq.��F�u����g2�v��z�o��K���4�"�;�mS��Y]��[9&�Gf�/.ov3Zs�;���尕
�uE�����Q�E���@�=,jb�"DV��_�"���W��J��a���c]�.��7��u�3 }����U>޵�\c��:nw�k]ä�\��cN�/�}����+O��t��FFe*2*"�
AB�řj*�X�QQ��������l�eJ�+2�)r�\eTc��ȶ��F(",*�:�����1ա�U�\�Tk*,Eb��U�R�j���`ڕVJ���IE�f	��V�mGT����1��Z�A�-B���*�4E���TF"���
����]:��ª�*��Ն4aV��4ؠ�T�MZ��F9B�2ڂ���H֣*TTU����X�QTAb�ZʢcTƢ�fUEJ�rرq�i��n�b�a]]�UX��b�D�.�G-UAF(��EUt5`���h�""���u��J*�V1�*kY�h�ZWIT\�����Llˤ�b:j:JVUȫE��1���\J)�6JKJ�j"�T��SM,)Xұk*� ��U��[�Z:E�EP 
"�P�S����^��
R����a+��4��,v���k^��f)3��L�]��iv6уK7�u��Y�L�c�;��:iȺ��m�վ��ʱ��4'�>�o��3��ڥ\CqKC�N��9�x��ޥj�quQ'�8����XN��9V�"�*�&�td�I��2x�1�A����0M�� �mWu�u��=Zv���\~Է~=K������k1�Z��U�its�͑��?>�Q���,8Ջ݀���
x��Y��M�7}��O��gs0�ǻ')��M��=U���M�6���2HW��-ۨDk�����/u��7T�I���{Z������CK6�^����ԃRaf�����O.��oT�鬢v�/�\�{�R��m=X�����J�Ν�[>��7Zs��<�*z�!ڡ�L��9ޜ�s&W��E�,�w��ʋ��NX�E=V6S��n�)�P����H�
�T_5��]����{b{����}���z�T3=�u�W�����U�Е�U�PW�as�K4����5,���;��3J�p{] v�C�g	V汝ry̋B�6/�=�	涘�#`Bp���F̩�R&��nvJ�:�#��t_t�_��*㬀�wmiZ�7.�sb�A�v����h>�㚉��,�Q>�1,�K)����[����'�R|�|2a⹯'.T\j�gs�����<��&	��cy3��ǈ��Sk���NZ2K�]�Ns1����id��4�)a�̨�B���gUA�هҵ�s ���	��@m��М��2�@[�'l��X�YoJ�ؕ:ĺ���Ԓ����w=58��l��S�E��{.*_P;J��1��O6%;�k�ˉ�o��
�X:|�ӸG��!��V�;v���='�6��e輴�vCɫ�P����wF����n��T;^����I�y�uBz��J~]3����ތ�lTu�*1���,8Ѳ����:�I,�O;�=q�<j�����u�q��Rݻ�OM��{�J��/H�:�{ޡ�^��^53FP+x�Ư�yTk��hO�'�
�3�Mf[���oJ�����\b��<��{�%B�gb��4��:�:�m(6�r�ʖZ�	bږ���B�����d�wJṪ�Z畦�qo�u�;*�!o��*]v���:XLU�q�w�,�T�r	J�1��yr��:�*J�%}�.�Vf�4R�N���+���]����e]v4�D�~�n��˄��_�����+�'����aC9�o�] �f��Ԡ,�y�*=�u���u-��p���S�⯅酙}�3���w�s�T��*{yv�ި�P��M۸��	T��j]�N��6��U��*AŦ���b�Uz^mBQ��x�r�*D��AX���&�9$۹p*��p+7�Av��bs��Q9Π��S���)y6��L�I�UM�[e�҂-E�K�[�][ʀ��Q����+���7-?Ryc�ڧz����.�CVb�4��{oc+p������U�u�]x���U��z�Z�Y[)Ĺn໇L�1¦_T���b�j��T�QUz�ͪ����x6e�(��'�&���p�����d����̹3eXwX��]5���=���.��١=:��Ȅ�Y��7��M���Bx>�U�u�d������d��#oi����3�15��;���V��[n<���K�Pϕ���]�aFjWkV�rJ��j�5�0�#W��/����	��9��3�s{�Kթys ���S�!1QC�BwN��u�p:��[�KOu`�G���LZ�5�s9V��*�þ�[��hR���Ưv�
�S���͋�#�����iܰ�kn���ю�\d�bb61��Pdo���k�h�Z��d�������e��ןǗk�/Y�U$�a�9���~���D|Wmw�f��ͪ<��~I�f��f�л��NM��G�����ſ'�irx�>���<�ވ�:�����s�7j�Rz���p�F��n�'�z9j���=N����;m�WgvE6��ld��tsnt����5oz�{��I��f�P�Z�-�w.����u�ٝ��K&��kDr���OX�|*�Y��-.nj�sέwH0�%�!�s&���E���m�@X�F��hI�`�}w���>��C�cb�\u�(U�a���Ӝj�����i3�|����z�m]8��3�9x.�ކ^t���
{l��u)����sɕ�tY��b�Aj�f>Y�Ǧ��Τ5s\J\w+��3d�D��| t���ڔ��uֺ1O���Y�-��Nvc��V�l���5�3�H��[v��u��b��Oh�+�=�P3�ө5��~�������O<^��:�wvou)⳯�NuTA��ߓ�U�ba[:�v�����yg������ΝW��N�/��qV������Y�����NȟE&8T}�u��tI�jkiEʷ��W걓�X]j͂���K�%)ߜ�;G���3.�T�[U;(��w���Wob�}o	���̫�!�����d���KqlfS\��+�eV�a�u�u���Ԗyѷ:|���w�W�gި�-�j�j��^H�����p�3pzri�����w��?hMq�KOQ�g�V���m�:f�48�����k�u�+7�ki����`+x�|z��Ŧrum��N-FuF���z��V�,�v��KYsR�u'Dy�;8��:����S��e.O/���CK7^t��CcoIV8���y����t#��/Y1�ըJRC
V�f��ܠ���v�7�����h���HM��v�)�3hF�;.J�ݣ]�_k+k�sR�2�,L�lmm��藃���+;UӚ 2�H�O�{�
.�'���\�+KS�!��`��[@C�;;�K'��J����:xNA�2�����r�h���I�-s�c�����u1��U�u�W�v�rd��z{���i��k���)ۿ�v�B�B�=b��{F{���L���գ�v<��n(55������%7n�]4%P3�:��+�����\i�T��Î���[����O�5���I�7��*�˞��FqW��ZN$�J�6�ҫ:(WS���'׉D�:�Ox�p�ᘊHp:�\�P�)�$����[���2�'{e�^�S��<jt�0^CaVM�0�Iͭ-��C�_(��qߣ+p�����1�s�Z�j�Vj���oet7��	z���~��J��+���n��f18�������Q��y@Qƀ]0�;�����uӗ�fuP;v��Y�g��kK�f��Й�@�����d��u8-{�N?w{M�~�	.��)*���䙶��)򷞲���ꍓ���ߩ�n����r=��Qs&t�t�@���΁bR ��8-rV�W�i������3@��se)�.nF��3���:R���ǊW���ۏyv^�/����ʺ��'tj9���n���9�.�vU�qlL�|�.i�ʯz��^�6S.c��*�����@�_T���Ϙ��5e���u�-���\d�BU7���wǦ�T�F���5�[<��p�8Wz̑W)Ej�0�k��hJ��U��δV�O&��oQ��r�i��ߨ�Ư�g�f�:��K'o�J=|L�1-�����3WZ�C��˱���6O}]�t}ggvh�d��U�Ui��{�����*����u����΃��J��͏us岵{#rjzy2�J�R.�y�t�i[�.�S�\��<��ᒛ�
Ԭ�٪�o��u��bf5�6�Z�v�o9D��J7���qω��C���2�(��8q�U�ν���u��먀�n�9��S���=༧����<�d}�sw�}���[�؉�B��>��[:�_k5�IW�F���W;$�M���9L�&�:�
U����p�ɋ*���J�P�_t��;G����@g�o��L��7���b�բw��Ӽ�}3�b[�@wb�Ej\�\��s�y�]�����b�0�\�-P�*��p����^�[m�i��AU&l.�O��̖o7�u'f&�*����2�
���lwN;3P�]7���?lOJޥr�0��4CLp%����b�7� �l��ݡ��
iz�cbT��BI�9�w��u�9}��&*Lr���U���TR~�.��n=&c�ڧ\Bb��0��B�pF�e��m���QW�)���q�]:�U�˜�ZzkTin:����1�����d�V�'Ω[�TV��Xr�0/i�֎�񼮺yUj1���}�-T[K��ݦ�§x\�Z%��{�����V���Azs�h^ڣˑ[X1u��S욄��4�?F����x��c??9�y	���5^��3{G�qPsI��]��k�R�+�F���5��G�����
뛵Wǹ���w9�G��p��
�f;�d�ۛ���]�`�Q�+�%�p�YSȉ'&��9޽"YVrJ��݄��U��E������w0B�V#�K��0�)�U���mp���*�h��J�t�Y�/1�E��8�A�j��w���-���t��~|2�����ϣ�-���c��u-�X�u�5`U
�&&�7b��e�Q���^.د_%W+�9�jެP�5�
��y8<7*��ԭ���iS��r�=�����_
�Me�.���\���������[�
�;�3�K�j�]��l:����w��0��&����̻94�cn�F�6�#p�b��U�=���\啵o#z�M3���U�������4#�ÞW'��)���i�*{�U�¦WT��7�7�ɉ���j�ᩡ�Ͳ�a����T�~.���&"���3�"7�W�9U�������"�d���VO�%Ls��JlԽ7#��3bw_N:���2Q�J��-P=_\	Y�=X>����/�j�G�^�8��t�{�4��C]����.�Ρ��{�RY���N�x�Q�vdŴ�[��D��M��/�l�foۛY,�KW��y3FH�I��Y��Ȯ�q�yi���z[��٫�&�ՙ��0�c��`+/ yQ��=Y���L�Us�z�V=
WP�Pՙ1�s.t��>��[��b7jToʌ�g(�J���Z�{�jT�g_>dv���|��{��p/j���9�G7�fT^��7��v�M��b�m��8�hW�c�\w��f߃������]�fz���Xҧ��^)���ъ��V�%Syq�W:�Ǜ=赇�OU�gsFٙ�����4�6hύ�u���-F��P�<�x�!���-��1�ݐ֩�gU>����N1���mk3xOZ�O�2y�r�X�T6������5V�:ȕ�ު)�w���{U��*򞺃��D_%e=����n�9K��q�:�8݇�p��)ۿ�wT)��w	�����=���OB�$�������w��oT5�X�q���ݻ�X�\	Ft-s�!�(7h��q�M��T����}Y�e��O��|2a⹤�ʿj�=��'Փ׽��k�ʉ��i�Vm]@}z��U9Ί{�;��p��`K�Ӹ|�+MT��R�a0��x;8f�&K���||:��`�����|N
�e�[h��K$�HpI9��\�O[Rc�`*e㚧E
���dCx�:<����?n7Z[�Y��Wv
��s���ܽ�OT�2�V�|�R�Z�j]7��+�\�9�l8�o����?8���X��yK�WV�9�\���dPT�p�+��`���6r�h*�gGL�Z�.�#��V���(ԓ�����5��&���]y��6�4,�}�V�)�V֮��ڹ(&Z�Ȏ&����Yq�h)�Ņk)�']u:rp���-����Wz���/ܤ�Z��;}iB�i۫j.`tx^�92/f��ó(
P����6��_mt}�:��[�*�ŏ�Iڻb�1�J�9�F���U�%LWWu��:K�]��t�P�g}p۱՜���{����'&�Ԭ��ɣJ�����Gv_n8�np�4t������uvo��K�l�|���6�A���1t3�l#�6�s���u�9KcJ�&�����
쁔ռ� �WLpWŚϱnޱ�;��Z*�t�7�Y��{�%G�h�dݳԎ�ppYRv�κ˫�nEʫ�u;L��{�@�o�[t�*E�̃��I���) �JW�N��C�֔�(�c��W �lR�������u���d:���Y��MM����.���oa���M'����툊u�]t<�yJ�p��5�,��o� X;���Ӧ��P摶m���f.׀n�j�����w9�am��s�� H ˝$x�QK2�>=�,*�kF��'.������Lu)}�W^�����u�b��u�����[����މvȨk�ۏ2�"��r�C�4���L���X��;���ei�Q���N���^�����Gw��3s\�^e
�v�G��88M�2m��<�j��y�k��P��ٹv���Va����
��x:�K��3��!�4(��� ��J[?2���5�O�]��]��JB���'*(霭��!�*��CuԎ�����2��w�rm��a[��Dv7G_}�+�[��t#t�2�������o-mv��ZUsJ����y���`<$���`���t�;��p�V/�銲�%�]��/��u��S��O;�B� R�=��D����V�������ⱥ��b���u��Őb�Ji�~�5N��8������\I��sN�$]J�����V������]@`�w���d�ݛ�N�o*��\\�"�5�C����L�
V��Zݦ9W|kS�	����[�JޗvXڷ�޺h-jH 'miƸ/@l�n���1�m*�oPޚ�
��� F�`��"Gwd��{���s [�c�%�����L4�P]�4�G����Y7��Ⱥh'*�"�.�W�B뚮\�<��
 P> �ϩH�X��☕�1�-r�&��mE�X9����Ap�J�[5k�f����	l++KMe�B�V)R�eb�]WT�`���W8�
�:��PEE�QV"��ь��&ae[E%��cidEQ
��U-��"����-Km1��MTY��R�֤s.��H�DX�UKF�Ȋ
��KDm�B���TE
[)E+*c�%�C

��Y���k-,-�%�X\B���e��n&i�(��H�KM#�XҶ��Q�Q� ���U*Q�Pĳ)�H�*3V�Em�@DF�+Qb���R�k�8%eTiB�X���i�A��YZ��Dժ�(��dm(�)1��*+��QC)DC-�KN<�[����n�Vk-ܭ|.��2TΞ��f!�J�G����:�9a�K�2�D
}���챎�����o3�~��<� ^�m�;BG�)T����-��hqu�/��s����o5�3)W.�6��QԐ�FWW��y;eti��K��q�p���׳��f�=칀�%&j�6D��=�R�� �+�:������ �n��p���P�ugzp��na���S�v�1�]y��3��=Q	�"��5�=�s���3�e)B#%������;�����ۢ���ɭ&`_岷�Ψ��:��̪������LTu�*8�O+7��-vx����]Al�uH���|���~y��
[��ݎr.��ո��;wʊ��f�D'�6�<͵4E��jZ�+Z{{LQ#�]�=�t�p����^�&_�ͣ�>�%�f��x��j����ee��V�ԛo�fS�b�\�'ނ��]���뛵|{�f��!��zpl��G�p�D!�;L�7�Ⱥ�b�|7��� �/�(#5��4(��^�c���	[�>�]
X�q�j�d[�z���|��tM�Uv�L;��][�����Ke�ֵ��j6[U>�g;��)i�����xe��E�q��W��}�:��:6>�ߵ���P�rzC{��m�]�V8y���֯�b�n��P�$;�}�.�Ʀ�C�튋me��x�ov(y��bn�+S����9������k���z�d7^�h��+��Qw��o;��j�g� �{uι+=�iK����cR���W���b����'���O��SȜn�Y��aU˛a�cV2��c�)jo�dq��{=�jڣ���W�Y�ǈ5�d���	�����Z�N&�͞��9:1�I� ���5��և�k[$Xoإ���짴�wQ6���D�Ʈ�q*S���4Dǻ�/s=6�ޒ�f��
�qB�0�L�،�M���Z�`��!����5N��'\�e�M�CJ�O^Gp��i�R�pK�~�9x�{�1��mS�!1P�9���m.�#Vt�'r���xӾ���:�<r�N\�Zzj5F��㭠��X��VGu��σh�^�E�����(�HԎo�BX�5��{��)�OQ�ˏsЎ_v<�tb�ΦG1ص�d���Is���nu�匮<~�,����-Һ���9h�r�����W��Q�*o�Ob�'\E���C�<��:W)��6�_z#��YAg8��a}���Ia��$�C#��N�7��O*�F:אI��X^�� �R*��Q�FJ����k�5�6Z�{�d^�)�0n�Jf��{F3�⊻}؃S١-ޭ�[%���T��kW1�p�_$�f�ɯ%�c+g�+�amg\	�=�u?QM�O=F�1����N�
��Ozz���9�س_Dw��m�;�}�������y��ڞc�C��u��}����יޝjZ�}�Z��u�c���q|�z�us�Q�z�<����a3]N ^�>6��j�:���!���/O{��>ֹ�����.��O�>��K�݆��0�Z��U�	V
�vC�����b��ex�J��T�5��V��<��'Ⱦ��W*z/��^��wg���NK�Y�h�>�=�ʱRq�f����O!=����2��6g��Z��Xl��t�ıv�oE�9�-�=Ku��*]�_]L��� x�B���9�-qid{�;g!ѿ.�>�\���Pw�+r>ڐ����w�I����@e�v��Z����bvms��;n�>�ȕ��ݫ���ZY�V��mR��S�6��j�=�W�G�J��_FR¦�frͿAW>�n{:�E>.��	���sg�n`��5d�ޠrݺ�*�f,/cڲ}�*c��IJ{W����h�wҪ���Z��悽��~P:^@���}6���̥�:�w�q:���t�4Oh*,>n��8n��\�ݴ�"���v��e���%"�6�h�K(�OSAl8鬧o���ѯs�o=Bc[�y�o/�Y)z[~�����T�v�F��SAm�u��,9Q`͸/���r��-P�����)]�qW\Sګ��Q�+R
��窣���S�c�[�Fy��u���S�Bj�����hɾ�tq��U�r�Zʅ���������	�!���#{�K��iuʯ#ko�k(��u��FO>Eo�<��3R}���{ޱ�3_��:ܻ���P�^S�Pzب�J�S�Uљq��D�R�zb����{>k8G�	~��x\���ݴ�(�IE�=x��>�Yn_�+w�y����NQ�~V��0*]��.h���� ���(�80�FV�D��-�&	�xr�=p����77�����,�b�&H�W[�w	]�:ݣ��%_NK(��ꯪ��%���jpu]���P�{PS�p)ۍP���u\�
�%N[���ת`�{�z�;����=�X�q�>0��ac�cBU���bE�+��W�RU�C���j�O�5���-�ɇ�漜�U"d&y5�rm��L�ʪ��\5@���Y�?�Om���U�D�V���'X˧����$�q#��85-W�iu[�Me�N�ʹ��糨@�`��,n�MT��h˝,���VD��(���ǲ�
�z�d�1f;�����5j�k��7R{��S��9n��èFȞl�]K�v�����`��J]�扜�v������&���:]��0��B�����}���Qs�U�Ԙ�r�f��MZ3��b�q��KuИ���wF����nM��L�y�9�0=������|�ݡ5��Kt�����e1^������/2G�/�'#~��r&;'�쳃�#*_�.e��5y�2(���j�n����w���AE�R�MZ��'8����C��F�����w]���kr��U[����\��0>��aC��J�Pֵ[o��X�'(𷹵s�s�gN��}�}�U��k������n��Pڑ�¾2��{Uj1�k��HO�7�-�+.稃���ʄ�j#-^V�6i,���6�џ����ӧ�����֌�d=��[�/��~�=���)��y����m�=j�1�·r�Vr�t�zu%��sʇ˲զU�'�z�
ҸSWm�jr�M�`M�w3�p{�u��\�r�Z�c�}ͽ�+�XX�[�$rc�r'P��d��v^�]�WaɎ~�w�½|�_�t�S�Q�z��u댘MۭtX���IT��Z�M��ӎ0�Yj���ɯ>�jx<ȘC�++B�T���>�r�^Z:���X��o�n."�[l{�?5�Ϊ�gB��d�3�,W��.0���iB�f;�}-k�^�o8�뽠�6�3��b�{~"UΩ�+�1�&/I��M�@�^����jU�xs�Ks��X�[7����O�0!P0u��M�ȗX6��NO���C�>ۆ3o�߭���z+�(�o6����c���xqpK��H)Q-qʔax�#N���սX��Wc+���q�V���sl����Y|���&�����YK�&�'V���4B--�uǵ���V:n�Ðp�We0a�D�o	4���\jwu&�9��=jq�{�������{��*�V�_n�S��HP͊�*5�Pw℄���b��ԓ^e�p�RK�B�@�=���byt���S�v���lEΞ���.kK1�2�q�����<����6�0��6�sV�)���Q"�����U�g�,��+:2��tz�}���m�����,����M+wʊ��8�jA=��D����V������
���j^[�`�0� g{Y�Rp	��=U���)]�J(LN����Q �tJ���^� c;���+y��پ���]�����4�|�78��#VuP�oh�N={Jz�EI�(Ѐ���Š��e�ER����i�1y�P�����Wz�`��z�����<�f�!N�7am\;�vfjڐ�x�>�
32!���U�r��<�Ӑ�ת �����D��c"U��7�
�y�n'��,�R�ɨ1.v>���2����{s�]�S=>z��7��a�A��*��JM����R�����)P
�u�(�d�>J"�p���a�k�袷�P�<[(!����Q7u��������p����4x�{R,����l��ڒ�Z�v��td��wε[yj=�9�w�OipM���*X�u�^X�����9�;)t�J]�U��<]�++�c��Ջk�\Ve�ϻ��R	�%��y��K����"����؛l)�����)�ø
aIB��!)���z���ɀ�x�E���;<�%Ҏ�gws;��!����op���z��<s�c��4*����&�����s��V�uگ��Y�~�C�Y���L1P��	]y���-���F>�<<9�և���q;;�7��P��{��,��j��B�������7<��!;�9�B�28��k�n���*�t���C�6kC�<v��VN:��٨���yןګY�e9藕�}Q;��m��f�8�)h"�b'�'�'�D��'���6]U��}5p�[I�U����C2��{Ue%RB����]8u��U�c&I��~�
�<5!��b�S��N���\��]���]FW-n��A,z��
�<������8��o���/�:k��rW�v�w��

��g6Z���P��l*����A����c�EG<��z�N����#;���q�����7���e����7�:Pd�e�Q�����F+�����`T���.�1r��{�����mи��WÛ7�vuJ��ڒ��ۏ]z��ol�}�Wd�(��L.�n�vM8�i#�s1ut��EvNi�.Z�U�үB�YM�wK��ʉ��U�pS{rb4Ɗ</u>�#���|:���Ll�nb�_G�ވ�*˓������&��R*'6�E�Zb��
�f3b
�!�g��T}:"����3�p�U�n{�;Z��[B�%�c/�D�c��X|*Y���l\�^�U(h�Z/x3��Me�1{\�H��~�Y����;ьOY��V�T�&�JIm������o�:��U/�ain�T����7���?��ξ���6��2"��7�s�PR�
�OK>�`�0o}Y��;;��Rvq��71�
�S�*1D���ݱ�,Xb��t"�T�b�jv����s,#6�nE�I�t�"^a�L.=���cxױD�p�����c��fB��QTg�����-�{�%�kU���پ���<��ۅ%鍄�pRr	����صֆL�GY�|�O�A��A��z=kC�*�Ҩ��.g/�y�vC�=�;�L�
}DL���7$;6{�\�qe�v� �iԴl�%�����������y�,>��j�Nͻ�v��S�.:s��.l�'y ӝ������{�h�7��x��k�kkV�7TgH/�T�xxfɐ�L���ZԻ�{�οM�,�`��+c�̓c|{{�$�T�G珏y��6�K�m��Y�]��{Bv��z�]����I)�O\�<�p%w�:u�N���o7_W=���-�·I/�Ề{q���u~����D��u�7���~�ȣ¡�jbQ��u^YDJ�y��q��Al�R��7!Ğ
3�@ӷ'#��Ԭ�q[,L�e1 D�&:d��*!�b�~S0Dk�GVDLv����u�ʔ�"q�����Q����Q����wئ�;bǐfV�i<��a�� Wm��(�I���"@D����ޭ.wM��LW��'j���(�!�����vq��]��V���&�*p�3�٦ϩAO�X�j+�o车	W�a���Uk��\�f�ݧ�cp�������3�F��q�mL\%�t�ٱ�
��1!���f��S�p�Q�b�weCx�4�9��#�����	7X4w阴`ꐍ��dP�3�hdlt�����7�\&�uP��*(_�\�
��C��\��Į�щ�#f�|����r�:(Q�\Y��ݫ� Q���E^Uy��[P�KÎ�TCvƋ�6����ۢ#�����Ŭ��^��A���]]Q��6c�Y8�y^\V�� <1����.V0-��Q���I��%�`dJ��Ԁ�|c�)�W���� *���n݇�̆�F�D{��EEJ��">A��[��K5l7�l��
�n�x�V�l8��k�S�9�!}bG�
�Z�u6X%����si�����4%f<�[N��'	���$�r3�V��ڼ��do&jfV�̻���˪�]l3�ÛY�t���;3{�=��펑�r����Ӿk;�gZ�N�kyrU��*��v�)�X�W���"����:���7����rdY�[K����o�6��WB��sE�o�}R�XQ�FU�:��2:��nh�� �M���k|�WQ�����ں7:G�*<$vG��E��&E]y�P�&�Z��Q:��v��9]ø+[�*=Y��䒯�0�|m�v9�Q���{-Vȥ�.�Æ�H���m�M�j�{�y�\��B�T�aҹҴR���O:��6R��V�go!J�\�:B�w6��9����+6��FaEd�t�����p�~��{�+�]�8&�M=1G3/01��$y��s��qk;/���=��x,ޑ+r��y�j��E�T�R�U�Fz�h���cޒq�=V-�e�ye�]��WY���.e����+��:��d3,v�Gn�p��e����Iӓ�IZ��Fs�A�C��(Vs]�3�Y�M��T@\</Ng��P޴/y��"�a��q��֍�#6��	�x�y�\/o�6���D�])�I܇S��,�m�+K�t���ha26�\󳺬���3��A�dٹF�t�#���.�I�gvK�3e�Y��7�f�>���\�g2��Y��kecי�:Df����T3��A�db�m����it�Ov�z0�cz]�V��&,{�4p�L2��;]��TՅy���[{Y�o�!z����K�}��>s[`G�n�8������7�!�H�{��1os���2 .����6��oEV�6-0�ӈ���7�=�z,��q���홖����Ĭ�Â�[t)֚�I��-�ǵ*1�-�,d.>Q����=;9������4�dw�׹���j�U��p����^��Q��Y4�N5��M�i�y]8`?�"�sQ��i͗�|%sU%�ѪN��}t�GwM`�p��\x�=Y���y�n�����Z5���9�j��I˘��e��F�^�l.��tN�uJ�a�cI�X��,B1��t7~����3x)L�m	�൙A�8_W�:���f�Tǈ�O/u�����XYw�78ɽ�� '�-�];TϷ�rT7n�fC��	��n�������Ck���Fij�N�)���탍h(�u�v,v��ء�Ehb�m��V�9&���8'��Vfep�j�Z/-͒�9��'�7u�Lom�Y,E��ˡ���k(p�3��h9w7�&F�n�������P���o/�~������Eb��m�TJ�[j�J
6э��ըe�`ѭ��&*`�k-K6�.kut��\�GYLf��e���i���4��#��1�LF&5km�m+PX(嫕E�J�V��R�+U-��Z�
�ұ���ab�R�kml̡m0��U+�cPQ(�*-A���FL�U+�3��2�R�E�+m[E�nfP���TLJ$1�*�r�Y,YX�-.2\��ƱV��+
32ॲ���XV)�Lq,q�5�X ŭE��R��B��-UmG3ĬEU��-��6��Z�h�1*�ebܦL`Z�ʡJ%��X����Z��m
��J�����11��G��4�dTf#lƸ5+R
#D��;�;0��S;��k}1�%����u��v��Nf��q�h.�rL���<Z˦�o�P94M����-�u�B�k]�ĿG��{ގڭ��ӛ�&����mD�~� $nTŉ�d�}��~K쮹����9�<��nr�nmc�I	]�/:Hx�bsN���a�0��ޒ��8"�G���aA�]wHoT�t�1�Ea��S-W#8X�*���&Һ�qԴF�>�]md�YyOI�S\�%n*�{�Ezm��.��F��<��%̀�Df"i:<M�R~����ݽuui���s��N��*p0��ō�(g��Pw		��X�9��v�=Kf�Zfs$�Mα\o
}=X9;c�W��}7f�eE�S���'U��e%¢8�r�*��Q�.�*�����7��2WI/֢H��v��3��V��t�~�=&k�>sU�Q�$����i*2u�R��m:�Nj�KˊqjA=��.'�Ά���VNY��/��@.�z�E�ˇ����F�ZK�}Dvzl���x�T����Dm�TE�-���0���G;u�(��î�ю��
hϫF�jY4�|�f��u�d^��=�g5_���:岐�%p0L�zPv��U�¶�cNVې�>,����[B�_3Ȃ�X����Ŝ΋�n���bt0T�[�;��� �i�՘���v/�*�}��z�� ���Ì{��HPy��u�VTb�u�%w5��{�m'J�.�-�Zz��-�ge��(�}�{��z;:���d����k���[.�e�M%,F\+�\'�.#^�Q�bڞ(��cEfZJ��x���B��G�ok�$�O�dG#Q��X�aC�xT<uສ�˼�'<nfr�:g�HN1�f�e$r!����X=tx$oѕ<��0�6S��|�HG_B���h��tݽT:$'��p�w*�n&(W�TN{,J\�x���mTU�]j��;��D;n�v�\t_ѻ��=�����J����JnU�S�d��Y\N#�Er��ٷv�A��ۃ��}�5;��(���#i���ϕ��(�B^�,
3��T����=Rl��t�TY<�̍�=Y���L1I:�@�Cܩ%UlS�p����;����5�2�X���W\&b����;j�D����X�:�[�>����޼�@�\���(���=^�<"��0��\=����,�:�Zτ����t�mof���]<m_���&�!��.���	c���+����w�����f�;n�{q�Ro��:�l�c�CJ�{u����ͤ�21�u>����A۪]+Y�.�yH�y���lg ���p�Z�.ʙ���We=Y��C�����g9qQR��œ�x��;���=(��]��ny������ƥ2F� g>��ꯪ���u����˖�������*��ڒb��a!��;w��Uvx]ྜ�%�X��B?|�NL�M���T��]X��({V���]���V�}[�G�J���\��׃��J�Jљs���!���:��`\)�]�2�1q�(2��lA�*p�k�CU}�|�[��(˰h���9�9U�pue�˜�Q����M{���9Տ��F}}m
�v��ևW|��z��dI��s恼LU�>�PU�\�m�A(��9�r���-�z��ᶭW*+��s&�̈C��ˮr ��z���~c�}�}�W�ċ'̩�o�;M�T����u�|hG�\o}��|
��nEOt�?�=�D�W?<t���$�
E�;�8������;��I�X5�{́uC��g�5����AN�4��+�k4�3���W�(:a�:�~�c���ϑ�[j���&v�e/�{���;��Y6�=�Cԕ��'�9��6Τ���]�T:���>�0���AAH�9��q4��S���E'�ی7��㴂�q9��x���H� ����zG���F���=�����d�~a�1������Y8�N]1$�5��Èi�5"���f0�
�}a�{�ĝB��&��T��ԕ/)�;v��/���+8�V<��>"��<G����u�U�7}�E�~~��<��䯩�2�'���1Ğ{CXu�8���6�S��8��!�Z���1??0ě��"��T�xw��&2�zʛ9���'�:�Cٙ����%C��I�[�����a��e*�=�/
����y��,v�0�IU�8'�oHЗr�'0�Z6�]���-\Ԫ_"��-�B������L�q��5w��r��q�U���TQ��|�xL�k��6���yQ-�EL�I�+�I�v� u+*�t�7j�y��.+.��)���꯾������O�<���8���'�_�h���T���m��
�ܽCI�'�� T�q%~d����$�Ѻ��Ă�Cɺ�'��o�λH}hq4�>����D; dU�fB�9��;�Z����j��2i�'|�&ݧ��I�z\Łְ�
����&�j�kD_X��Lȡ�J���N!Y�O�O����JΦ�C������S��B>#�7Ct���5��ӕ�G�I���;=�	봂�|�����5|� T�~f3�� i:Ì�<����Zɹ矵6�ĕ��y��!Y�%M�8�a�<�g�XhG��#Ѣ��O<w���������=�'�8yC�&ЛϲC����I���ns1*[�'T�2��� ~d���q�=�ی'��݄_Ddo�~��dw�>�`����n��"�ҡ�:b������>�J�I�>B���%tͲT:��d�ggP�ɱ �u�g5��Lv��Y����m4����o!�:��d���x���#�D�M�<_y\���ZJ�X���$���&�Rc�Rx�8����i�:`q����B�q��c���Iל�Lk���T�6�jy9�4�q�Xh��iI_�w{�����]�4'{�!J���"����k�!�8������x�� ��t1=a�u���bu��c��q ������I�%C������ALa�bl�p�<C����3t�|\�o\�6��/g��.�VN�����gY6^kRVV0�����N�Xxk����C�{�4���|`_i
�Y�1S��ɉ�
����o�N�qϩ�z��I�c�w~"���k�9{�~"��A�`���1�H)�:}̟�i��0<�{��������E��C�k���M2�g�bz�I�>C���:�8�*y�8�I+?8Χ�0H,�=Ͻxi�xq?m}�W�)���X��	""���I�O߮��{�i�W�<�<~|H(=�}I��i �s��yI��(=��ć�������񁦰3ۉ4�d�*znɧI�:�o�>�珏�>;���R�em�-�v��2�<�[�,�צb��C�bNI)X�9��+-�_�7�g���ηI��uٓn�3�Xc��X�9�A�y�5�*��q�֮��h�kHI�hKz�:���S������緌�X���׼���̛r�l;|�s�%鉞J���;��߾��������BJ�����a���~M�����`)��q��q%z��Ӟ�<I�
�0�ξ~�*$�֞��֩�y��E1��㤞g04��T���j�D`"= �q��DX��:�\	�����������ơ��LAC�P�=՚H)��ΐ�i`|����L_RV���B���y�L�ea��\���~B����:�6�P��,+�:d�}�w�w�s�=�]�����=מt�
E��ǳ��P���|�n�Į$����;��g��ͤk��?����O'�;a������.�P��;��֠~J�MsyIY8����~��{��ܻ��fg�y��n~��"�zDy���X�����/�p8�������ԛR,6e8�'��8��ɔR|�N�sۧ�큈q%~f�(u���PSg�1�O�ɦ��4����R�T�|Ǖ���f�%���x	�d�}��4D`�k%�=t��B�q��Z�Z�gb^��`u�>��P��1& o/ �_�R;<�8�!�J���VE'���&����B��9��~�=��n��ח��9�`�!tc��3�#�G�8�t��~�i1��ɷl����tΡ���&}�i%Cg��R�i8���?jx���1��٭d���|ISyd㤟!Y��=�������:�l��ך���罇�Lea�w(�}�bO���C�>v�@���3�6��8���AH��8￰�X
bts�6�!��%qgw��I̤�g�jc����~o����LĂ�����ŵ_=�����n����!�b�D��=��x�2�0>j����yIY:�����ɴ��>�CL�N��0�]�hz���㏒�0AH�|��i1���P�N!S�'���z~�sdf$F.Y**SB= Dh��<����>$7��Ę��d�혜@����y2��Hyi��Shi�ư���] �Ь��3�������螡�Z����M&$�������yup����<�>�_zj
E�*��OYP����{�<I�+=����ϩ
���4��1�V�n �S��t�����
���,Ӧ��+��:�`w�9��:�-���R��ާ��ܜe���ȅ�S<JX8��+���DzZDGn�e�`���ّ_��֬ͫ�b����Y��m��7���ܗ����(6z��]��u�֝v劒7�G�i�ܢ�x9�P
�>������9��%��Dz""]k����?C���9���a�6���MÜ�tɌ�_]���I��3_���'Xy��P�{�q6���=q:�_��q&����t��d�
E���lڰ>��B_O-��8��.�r'�p�Փ�\N���iI̡����x��PY�3Z����VLq�Ϩbg,��
(m��j�֠l׸i�J��]Y=f'����}��i��!#�=Q����������;�ݯ���%IS��۶x�D���O��'�&'~��LB�P��r{�� ���Ϳ�4�t�S��
�jOɤ6�&��_�=|淨�1�Kぢ,DH�BEo}�}`G�0�������7w���vM� ��:yN�L
���g��O��[��!�N�$�o��:AH�eM���=eC�~�4����4�~��?$��t�C�����bO�ڤm
��M������ɯ���f�~�����>ޯ|H)�
����m��C��.3�8�d��>t�PP�~�f��<��C��LCo�8铬�_P���=jN!_';���,��G�[�V��
�j�
�:M�;�I�d���k·�4���N߳H~IP�î>˭� �Pўd��V�a���4�P�Y:���T���9���fݤg�:�'Y����N8���"v>��G��D {p`����u���n�ox��Xt�̟&�uIY>|���c*|�$��9���q8�=��I�=IRy�d�z�Dn�'̩�N8��|�N��a��
}~��{�=O�� �+�F������~�~�AH�I��i;�0:�Xl5����d�9����m`~o��.�ShV^P�4��N3����O�M^:a�
�LI���8�"�<q"��T>L���ι���xs:k�s7���|?t6����<gL�=I��R��2)4Τ���ϻ��
E?0ٝ�$���N3N08����i��M0�3�v�PP��Ѵ<f3��z͡�b����s �'!)�2���_��=�#�p��Hi��R|�<����N���P�'����
��8�C����1%C���m�PR)�^��:�+N#�����'�ߴc���}k�?���Qu�9�j2o�h��װMU��OƄ��/<�Ε1��Y�v��<�|}s5!�޳h0뽈����@��E��t�j����ېr�W/{Q	彜�s�;�U	Í+T���5؍D�I۷̼�p��7�-��s���'>��]ӿj�����)F����v�~��c�?�La�Ru��̰��'\a����6��Pu�_�6��Y��=M ����9�f�>eN&��VO�?w��m$�l�m�|f�(��o���z��y�������?_��VM2��;{�m4�Rq
���I�]�>�&>2q��%eAH��m�8f���@������Z�z��T>O�}�v��PS�?����� �c.���O��'(����~������&!Rt��>v�L*q1����`u�)w��1"��T6y��&�] bN>�f��Ls�����$��O�ڧ�TAH����)�i:�d��$��q���ÿc����?�{<��|}����7���Cn��SL��O]�}�Ohi��@�y�N��b&!��o �O�Ys3i+�I��g�H�q>��T�h��!��Ӊ����Hq%C�3^������{�w��[E�ݩį��A z:~����b�����m�C;a�;�=M�$:�C����4�q ��i�jN>���:��?���j�7�
����['�P{O�7����d+������{�<DP4�?P�O����g|ͳ�J�RW�Xi��:�D���i�S�79�=|O*N��fi?2kۤ��}��q����x�CH)�=s?a�:�
+	��W?Wq�3�$��h����z#�f�<�&�ĝ-�k�ALOS:���|=�gXm'P�xXz�T�by�`x�Ơ������T�&2�ݧ�4����pP�1'�Q��~���#+�&�j{��hZϽ� ���O�k�l���M��!�=|H)�{冒z͸����I������֤a��J�Y�ě>�����by��=k'Y]�������D@z+��\�M��܍���V�b�O��4ԊN�{��l1�O{d��f�T+P���9�h����{����PY���:���`o�È�������:�v�P�����f8�LĈ�=#��R��K'��w.��7���_:CI�N8������`~jO?w"�Θb��]�i*)+��zͲzʟ���i4�d�)�m�����&���u���T�'�"���,E��"=��?}:-%�v	�a�.�t;�o�J8�^=޾!��*�J2���	)XS��Uem�y[�����m[u=v�v@*�Z{�ۜ$
���%�S���s\��]��a���q�-rk{),���ֳ�M�������V�����[Uص~����{֕lWms��~�Cޭ4"�4>I^�q��<�&�R/P��a��� �䞆w����>k��T>O�y9�'��j
xw[�m��Ve���0ĜB�@��aX�G/�zw���'�6��S;����D;�1�ʑd�7��$�_P1<���:��;awaP�J�P�\���i#�9��&�
|��d�O��o9��i��s_h��R�S�3�U�AQO�:eo0�~��DCf3��&'�f!���x`u��O9t����8�a�Èi�5"���E�a�=��ӽ��N�X|���wU<@�u%O3�zÏ���?s!�+8�T��~�}�g{�����]�T�eg�g}�w'�_<��'�����OP�,:Ԝ|~��H)�O�w<���`u�y����bM��"��T�y߳l����*o��Rx��A[��q�|nԄ뷭d����G�IP�:^d�LggY<����d�*o������
¼Cl�yt��S�J����^��CR/ɠ�_��AN!��'��l�3��ZCB"G�EM�s?/2�~�Mv��m�ơ�ߵ��+&�Ro�ɷi�m�$�=���a�=ϰ�4��P�y�_R,��2(x��|@���V|��?S�P4�Vu6����Ab ���L���LIsO*��o������Sn�f���i>f8��	봂�q;�=Oj�9��P�P���vwyI�f!�g��0:�M�<���.$�y��O����l8�W��B�A�mnR�3�3�Os�?r$���.'��w���Î>0+<5��E���C��CI�eg��;���4�Ă�y̝IwI�c��[�4���ٝ��Y�AN�]~��"$z!�7s��=�c��
�mt���&�B�a�t݇��:��y�,�ed�5��*m&$�7�é]3l���AI�q�u�&��'YvsZ<d�i��vΡ��'��0�y����J��s����O�f����翾��]�8��PR/y�蟟��AN;d�i1�)?yg]$=�4�g��k�V)�VN2���8�ΰĝz�M�1�:��S��L`u��5�B<��~IV�w�V��<��Ohե�vZ����=�9oඟR�v�K��ͯU�y����.��Q�S{	�]���Y<�]��K����{��]���ѽj��͙� S�\J��X�=9������$���FM�ѵyV9��������P�#g/;V�����G�����7U��CWN�&w&�~B�䟜�ol���J�&k���ﴂ���������H���I��{@㤂�h=�S�Z�AAC�P�$GD>��$z>��Ў�D��W��ξ�7��^�M����o�=f1}IY6w�.�b����2J���7�{�6��Vk����C�{�4���|`_p1"�Y������P+�=�똋g��A""�ƥ&�&����+�^~��|�?$�R|�q|�*�C��a���$��d���O�1��s�T=0��;�.�<J���~�6ɦVL��OSi1'�~�k$�|����a����#�����z�~=��{��o���~����AH�m��4�2~q1��	�N2s��=�$�$�XxsXx��AACa�p��O��I����O�1C�܇�$=�?'�ߚkf�� �Ь�eO����O�﫶$]��[��}�X�<ǢG��ihi�ְ�x}f����������T�?NP��C�+��z�!�O�Vq���u��!P�%}�0���Z�l󙤊c��I<3�OP*O�����k���lQ���Z�,�Dh"= }��<Oj�Rb
%C�o���AO�q<���m`q��~��4��%a����N!Y�Y��4��Va|�揽�x�����!���A�_��Nn�+�� �#��Exi�AH��=f=�oZ����.d���Į$��!�Ne'��y���íw>����H)���a�l:�C<���@QC��<�{�0:��D;���
��<���q"~�f<G�c�x�}���u6�~}9ܛd���%�.T��q�9��&���8�'��8��̢��*u���>OlC�+�7���

|�x���i���sX��gN���y��DA��#��d\Hyht�;��<`u�����
i
��|~�jjq�a��w�m�ְ���C�Ę�^8��~eH�y�q�C��댊N!Y�5�}����9f���?N��|���n����4�R|�T���ȤS�������M& T�����>06��;�vΡ���K�P�T<��+4�S�8w�ڞ!�1`u�kY'��\� �F~n>}X�Q��ɘS�{c�:�4X.��QZ��uc�&��QdIWx:��W7K������鹣]�f�㶗Ϡeư1^�T�J[a����)�,Θ���-g#���yy҆.�RW��٩<ӷ���R�b����S���@,D�|���;��t�ߣ��G�V�C�M�uO�{G���=�����2q���ٔS��I�.�����P+<��u&���t���AH��8�;��� W\���y�'�\C���C�9��L��Lv�PXy�t�"*3���?p�p���<�'��q��!�t������2�08�g�`=���ef�YS��La�_g�'S�3L3��$�+8�����LR,Ѿ`u�Ld�H��~#$}�:x������Sl�����
$����R~q� ��o	��1�4ɰ��N ^�~q<ˌ5!��SHc�a����B�v���1��:�;�螡�Z��]"�'����\��R>�="�H�H�O�栤^2���a�N2��J���^ x��VzwϴO�>�*O�P�?$��X=���OXbuӿ�'P*�E�t��Y>eq��SL�te���+Z;�F�\/�� �A�s�l�����e��2�޽>��ׄ*��쪋0�������	�i��o/��o=��m���oR^ZS������_G^X<+U�\)�c{��ʨ˫�ՉI�������]S�h���C�y�i���_�/f��;-MAn�.2A���H�3IoBZ�Aũ��[�Ɗ��,�w>b��_�A�~������9�_��w7U�a��|<e�K��S�H_�SQ�ʣ���ωuܼ*�Gc�����y�~[�����3t��Sw:��ŵ<^:7�xMO��y\T��dG#Q����r��ȼ""L���-�']�'3��WF�Wh{�d��d�R4)<�|����h��-`[6D��<�x�M�`��>��C[Q�U�е��(^+wq��95�vY���z�M�a�lp�09׏7v����tlL��1]I�l�WC�XBZ�t;+�n��efb��!pf���M�G��1�.�t�c>�}}����]Z��{.r����6jU������F�Lr��i:��+{�|����nn���bJ\�x������V���2p��%3��Q����c�gvq}'�����]�R�I�XWN�a<8�H�e�2<�t:�eb3I��3G��%|�TT����(��4x��F��gsN�0���Mrd�58�;R�]n��|ޒ�����we	 ܇���.DN[�I;%;��,τxLVO�#p�zu�N��CS3)>�5wv�|�Xz���
���j@�*���=�J���ά��V�nvw*��%���A�
���Y虡S��m*�;�hS�w�ۋ]j�Z���e�õ ���L�0vP|�얝��gLww�&������;j_ "8��Uk9�L�v�ӱ]	���/�U0R�-Ws��LM��7.,%gJj�#���[��]V\ۭ�ј��7�٧�=�������pyj�CA��aɝzH�X�JZ4�o8��U�7gi̬smS����w���j�E,����|�t�=Ʌ�M.u���޻k��2i=V��ŽD�z�t�N�<��wȌ��,�/ts���ܜ�ԆY��
!]��]F�8Ȝ�G��ұ���=	�n�mí�U�i�[���J-}xO5�e$�FZH��Aof��,�o�����������J����RP���i���X�ָ�Whp=�{-򷔻2��\ᡝ��W1�L�r�`�lv����_��K �!��;V,r��ԏC4X��EF�Q���׷�zӴes������'[ڲ��&d&�:Kr���.tA�+�٢����-��L4�۽Z�j�)e#B�bZ�d�L�b�7�e*&�lD�i���sv�л9���G�M���d��]_;a��.q"�aǷZcu�ubŠ4{&7Q�<q��*�j�l;�0��֐��澎�)��W�q՜�NR� �[�TAU-�L.�r�.һ��"�j��1$�{W�7��^[��szN�·e�Y�5���J�r8�'�G�h�l��4mi��bn.���&�e�}q4i���&[��N�t(��|��r��A}n�e����E��Ôv�n��☠�HvS�wY��u��Y2�p�R��C^��ݺJ@T�N����ժ-����c�x����d��}bC-m	*eX�\u\�2-B�#RSvh"ev��\6mZ���� ��.u�5I;<���n�;���{k5e��1�_r�Ss�2sK5\�j]Ճr��@�!W:u�����+}�E	��,�D�g#�o-÷(�c+�MNv+L�,��g#e���p��?}[d���J��AR�eO�X֌�Z�TU
�Ԩ[Q�˂�2��ֶ��DJ[Z�YAb2��Q���&1���jʆ!L���Z�eb(���*KhUJɍ�Y�L��l�
Q�ZʭImc�(ⱶ,(����ҋ+mXU�����&$���i�+ �Z��*"��Ts0s1���Q�XT����*���dRV�h�AD�
��E"�q�)�Ajl
���r�Q�JR��*��H��m�m�+GZe�DV��X�¤*�Qeb�H�P�YQ�+RT�
�e̘e�R�P�-�Jʍ�-�,VՕ(�T�kmX�V���V��U�9�eq���VVZ�mZ�DV�UP�PX��R����E�h"
1�(�m�*V*-��e�5@|E@Q�D:�sɹ�+��󛉡�آ��A�*b]uܭ����o���;B�s2n����ރ��^!+�E+�i%�=�����h_Sz�l�|u]��y>���䎢�qsSa̪W����nK��s�Bl��I��"��;vv_���T�a[Q�AYJ���q1B��@%=V6T�dߣ�aA�t�=K�ޖ����"�F���QB��^��9���a�S
J2���z��Y43!Թ���Cn��}�{�g�^��:ΈCc���P7��>�6����ϗ��M��]��_*����>y��o�}M[��~�MO��a��}x�>R�y0�Nx)Q�F��*FkR����� >����6*�`ژ��꫙�W]Iǳd��D��a����7<�� �E;ON����}=N�Y�+��8V�G2����+�u��VE��(=�#Ց��n�[ٷ�v9iq�%Y4�K���wRM@A��צ�p�3a4X�%����}X���	i�>}��s����`Ȅ0�ot���j2L6@VW���3�l	1vX�us0;0g�n3嬾����&k)����� �텲C�����<YFz�rÞϹ��w�#F\�ɱ{O�ͽ)�Ћ+­�[�]�*8�tx�k���̈Yn���f�@|�{�٬;�x����#���i��Ba��Y�
�W�Y:�[��Ζ%�X��3 E3g:��n�}��}�ٜ�m�b���	-4�m��x��Ν��s;���,N��w���}U��UG9T�2����Bl���� /)�mp��E*�((��������[��B�E]ݡ��I<��ﴛ#4�t���eF���(2j8�(�*�W}�xJ/c��O�9X�g2�q�e8��6�T��ڱ�ز�µ���8�̊T�ٝJ�#��_l�7�V	Y�Z��m
�=ɴ7�z��a�VkGR�Z5w˓������_�R7F���[1p87�o'ͥw�,o�/��x�³ɻ%�x1M�]�ޭZ�[�;x��myT�0�-�A�6��zl1�+�".�7���4R�	V�8=�-�l��m]��P�\YH���AߡLhCQ���z��c�e�\AX����iU�t^jr.;�ZzE�p4;�&C{Hyl ���imt|���)1}�}���.�t���Oh.�ew3y�;i��N>�l���� yca`��x�1��L����;u�Fws.#���=�#��BtSٱ"��S��p�\��X��1a�	C��l���s��Ҷ��`;s��t8u��� ��RZ^\�;4g�WZ�Y,6o뫂a�Xg�A��oX���[��!�_��ިe�Y�]�T���.Q���Ȕ�ّ�C���Vr�MX���m7P��;����[h�D�bH�ɵ���{��Z���R��g{�6��jc��Nc����Ĺ/��8M5j��j
�>�J�%FM�<�h�|�z�&��n���6."T�f/��{�#Y;��15Z�:�����XK���Y��qF3[0��;"�̇��%n�!��sf��n���tiF��N^C=:��w���5F���y��g��*�)*HBc�K.��a���^�ӹ���;ݔ��В��q]C�񓯎��μE*�T�]
�v(n���b�ysi8�Yu1W����Q����ì�:� 4IU��ბ���k�i���f;��%��?t�����͕y'{J�A>;k�r�г�E��ee�R�N��46γ�����a��y��&� d�y�LFL9�H�rٿ7:�Sί��U=���< �Z�򺜮ƥ����	l
�i�`1�S8��:aW�]�����g�^�i��6f+��zP���9�f�T��j��(E?V&>TfI����y�u�+_3N��]�G��������;{���e�>�0�=�#nQ��l���4TL��yzR^vy�����;D�;�ͣ%��&c9�Hօv�iQ�M�i�A��W���[u��p6�C}����4�V����X#Ur�ḗS�8��m��)b]IX�M��=f�r���>�����舏G���Zӷ8od+00�i���1C���qg�WU�+��-R����p{��d��z��s\���J�|v�'�^R���(��{�j"�M�l��YC�9���e�w��Y Gc�|��q�8�T�n�L_�\�&���+j$-�D�+��Gh��� ��b��^�ۢUԞ�6s��������ޘ�G��m���]ŧ:�P�=0�d�W���*o:U�Q�)���i�r��a��<A�҅DVK��Fp��Ok�b�W\Y-'�c��)RB�<�'|��d�Ur���eA�
�fb0t���L�n�aш�P�{l�ٍ�+ܼ��HsDξ�}�nu橺�Ig&���.2�Z�(;�BBenwe��=���9�)S�%����*�%�8��C����m�^��u�5g���ea�@Q�z�^�}�.2��"��3;�vא�3Taߑʒk\�)�8Q��B��Va[:�b��2��xK����m��ޙ��2J�kd���y�ƹ혼����V�UG�*�Y�1�S���%x�<��C��[ru2r
ú;��R	I�EJ�P�E��ʽX`������6�7K50�����0Wf��2ӛ��D�+��n�]cn�,n�[�:W*���˅u�Ib��A���7�"&��j�IΔ�u���R��P��5�._{����Fts���֣�t�ke�,Dm��.�{^\�_h�g 6�Vu�ԥ�{Fz�;����წ�v�(U��6���Rɥs�))��5�q�z��U�_7��#n���Q[0Ȩ�{V�A�l��W�����?Fˣ�Q(1�`@m�(��5x�v��[�IQ]?F=��q�jB�83N@�=��&��;�����#��6�����s��y^<1c.pf}�3�g�̛[����O�C�I�F�!c8�\�{ihYZ7��M�����)z)�7�����!����ʣ�a���PR���&�&�퐯�W3�ꬔ����s��
�����p���gؼ[��p�BSpZ�T.J�f�|9U�}��0��d�"��݋�!
�s�a@�������ϺWU�mڙ˲6Tkl#��0�C�J��Q�%qy��f�\S�b�u�NC�v0C0�֌��S��u�Z�t"apΩ[R�M���	��RCk��O������w{C���{Y�U�'>�ϣ�.w4���;8sE�����hK]So/�&¶�E�{w� �]���@x>�:hm.ʉ29f����������T�Ի%��'��ȫ�>�W������Ӯ�+���U�����STJ���I/�#ޏT��R�9ɻ�G�ζ��B���/�������=Ect�梨O�$��sA�^��)�N>��L'1�b�Knr%�y:�'  ��]&�:>Pp���tjg�^���۝ڟfoF���D�te(��琕R/=*B7RLT7 ,7��?"UF��J����_�%3{_�q�f�A\��R�h!Q
D��|�]��FvLTs�*�)�y+!>�B7V���y�Q��]�Ѥs� �J NS�.8��C�"4 �8gM�Uk�i��Z�LI�/آHp�
���@ͺ�ع��Qf9L��Y��>�q�^���S����
�&b�/�U�>YR"��#6�caOT�y4#(�1Qg���5�h0=\ ���e�������Iza��mΣa�LU_�b/��hW	T}n�]s�J�)����]�w�X�+��Ъb�q�T2��1^��,�*MfF�cx��	�B�B6�X�K�ݸ�;�ef�]��YaW���W�Oꌔ��0��c+��Ҫ?O>�QP���fi��o<�}�{�fϦ(ƚm�kGR�1�t/����|�:�>�/)Wa�z�#�J��HM�R�g�Xte�m����������Et�@�e�Mp�������Szs�T�ى��Jnob�������NM�YWa;�9����M.��k���m�_/$�ִ&����"~?-�|c�Ζ#/���s1A�`��������}�&��P�d3�+!�U�� i
��?-����?��ƙY�������+�i�Uw-U��B�n�pM�5Ք4��U���$3�i��}��jf��7�_5�{�'�r2�T�f;�|'Ey�ؑ^N��X�Y�<�EK�P�9���x{Q%�l*��z�uHN9���Nr��N��LŮ}�!�T��׸�p�UMۢ6xv`�X�^ԛnܾ�APB��<3JF��S����䘫LR$Ɏ��nh���_��(�\�TT���ɇF��1V%�h;�]���+�l���{/��Α�]��e)�$����q�[����1�f�u��"B�%��W��X�ȐS{��ݚ;ޛЎg��*"�wR#d���A:�g�\��雿%F�7Tt���UT򥐦w;B���<k�e�\�,Tk�#�x��ۦ}a�|���W���v�缮/^&��4!s�����׆��mn�m�O2<�9��Z��r���,��r*�{�zX��D�T��Z����u*�Yܮ�����ys�,�[[���ʦ�;�L){)	��ظ^��'��9w������ٕ���l4�����z"&���4�F�_�GD��
�2R���ƪaQ�-�4(��0�29z��]��}�_Q���#i������[7·ƴ�c��ŵ�t��b���%3{)	����qj�vb�3��}�G/g�"{����w��6��	�SV�}���ˏ"��eha���rc��'���m�����c����c��Pa\,ؾu}ƪ�;uλ�}|/q!���-�_n�U���C�]�^b�mB�j��Ω�=g}.��6�X}Z�m�*p!ee*:܁#�N;�-�r�&B�^��#_'��� "��W}��Y��sT߱HL\k���c
ډ
��@H�j���&���DQ8��+,�+��HuU͌�5��|^���r��⻄�:���gD�T��	BdRŰ�71��Y�%�b((p���
��+�:�d1�\��D��u���r�@]��#+j��ٯ�x�۩o�����x������Ln�i�U)�`��Ӣ�9/&��:�i^-�A�HTs7ӭ�\b(���6��(c�^��K�V�K�Ҳ4���]��?ZU8V����.���v�}М��I�`	����z|U��r�8c�������'��3w��o�Hb�'NL��_U��ӻ�W��֖��9'
l���x��j��}0�en�99�(= D��P�k���U'�g�w��pr�^*ҕ��/әQM]I5���K�D*��~��r0�ʳ��'��o;z����"���}�ӎ��4��~��y��i���m�Ȋ���hp��ݞȰ1	c��wf�׭�˓/g�*�ʽ��&m�8�m�K���/�F4tyK��yQӷ��	�O��b��r��F�cj����L�]D:�ypj�V�|4P����]]�J��~�6�=X�ʄ�S�0�y~��)V��/���p7�Oڠ�8��ް�"K6My޽���o�����e �f�½~Nr���1z��"��mD�V9�]�Nä��#;*4_��uŵ!C6/N��>��{^�'gڊ���HB��o졽Z�(��+N<�L5�xىؙ���ɸ"Z�}��:�κ�2���'�u7|�wݡ3�:}��&۟=S��R��P�R��<�LP�� �u�J�qT<H������c"�0ڹ%�M���Az�SJ��7�l]�K�w��47��_*QAj��gU����F�G��+�U�k�����x&IE׻n*0����l;K�W��q��U���W22,.�3o5Jꏓԫ�e�㷳�:���A��}�+gN�����J�3��}݁X}�\�
���W�p�Q/6q����a�0��b����[\�'�M��:�v��<����p��e*8m�!�9�0�h}h��M^mÜ]�J�[ɹ˟SK.�uB�J�&�Y�%qy�Q&�_��0��
zf<(9Y�z�\��ȨCusb��������貉�fB뇞��bX�N�WUu��<��2��ͦ �������/������q�y�7}��Θ�-��ǐ��꾛�Lq�qQ־U��Z�������Ѣ_Ç��Zk �c���+�m4��Ӗ�s4���Qqy,;�K]B'K'Β�E�ʇH�I1M��~���̐��U;w�y5�Vj)B�gC!	�8&rP|d ��cԔ��<���Ï	aT"=��7��Q?d�h�r}*�S��AN��qA���"O4���W[�Te!�eNj$�� +�6���]&�eRO��]	���Y����G�r�{xX}�YǕ�nД�r���75nn�/��)1�Wتg(���C�ƫ����n�̹K���t!��$��`n�l,�ۓ;(MX�ٷ�6`	xzS9�&3����O;��-S=hL���*����dv����q�{	4�����ٰ0���CL�D:F1�Xoq
Ζz�BZ����!`r�aݷ}�xegd�uPX�����]l3[����.�����T\��P��ᙝlGS�O��C�%�x��q>��	Z�{��&'m5�B6��"Õi-R�b�cB] 1���h��0Wm&�׷I����� 4�u�u `�1���j�����d����4m-F�ӫ�묜��'t
�O��t�B��co�=���v�+d���L�Ț�Z�Oj���5+][p�]G9)Z��0 N�3�Q8����w��*I2q�]2Zt�ӼUr[���dZ�H��4��9�'sE���ۜO��n�˻I]f3ع����t-[���'L���US�e��RJ*!]�8�v�,�.����-��ƻ��ʞ�C�:9��wk�}�2�L�<�ɬ:�*l�m�N^�	δT��5403i��MU�T�v,�*;�����Z3��7��:s{\�ă�J��u�7�0+$8�#��<E�Sg&�'p��0�A��6�h�谁<�wH���6F�6�ʒ�Θ[�Y�tD��HT�����i��%I�3��>j�>@wt�֬�{P�G)巍G}c�hL�b�N�k�J^�}��%/=,4z�E�m>�4�7�>����9W(��n��wO��jl	µO���ԥ�v��uۚ��|f-�V��u��l&��8ŵF�9s�P*���]ޙ2JiV��"6�r4�I�X6J�;��}���p���Y:.�<�V�:�u��6)-kwN��,K�nЁ�㶁�5����m7���X*����ܠU�hkmҽcU����w�b�Z�3 2�t*&�*��Ze��XT��YÛ��8�μBm���zQ����:eӑ��@���V��V-�@�D�	����3:���[e$���G�Q���`�	1\��ⲯ�]@\�A��̡]��(��WP���}N^��!��[�1�媃��<�\�A���z�G��^�}���f�a�Z��f�nwZ���y� ��{�z��[��`ZHR�-����n������I��{q����6�g_j�k���81u�b§WW!�N�>��Vg>���+�V�
f�2᝷� �p�p���[��rv�a̼=�<�i�j�r�6�J��n��P>Ū1��nr�֕�	֮��;��_|���[��D��\6����j�b���$�ܣ�`⮝��������̃K/�@v�Erv�P�t����^�X�Zr+�*�/��s�8���v��p�M� Z\p�=˶��b֌K��/LX1I�"��X�Kl�b"[E%J*V%�F��j�j�%A�Z9�
cUm
ZE���U+ �!UR�Q��EE����P��bZ�E�h�e@m ҂ZF*ַ(T"�2�h�����5�`ִ�1b
�#�R�e�ĨT���*��	n5*��#�E��U�*�����m�Bڊ�)hQ-DkjE�B�j��,j%IKJ�`)P�jԨ

�iV���F�#&5b��e̕�U�m��ԥQ���b%*ZRU�Dj)UU
"��
��U[ih,
�AFF�-��m%[*�j��db�G-��iR�j��),1.Qj\�!F̵���V�J��V�Uq�Tf0�1EQQ��
�Ҷ�6�#�T��EƲ-H,m�1�8�m�kmx��`��  	0J'�v`��Hun�oe�21��oL�h��f���л�c���5< �7��ts�Y�f ����,7�m-_��軕3k�dq�<{k�'�#�̈�5�Fn@t
�-hi��}��:�-�Ozo`�.I�����H+��lq3�Xo�Σp=5S��E���+���݌�r զ:ϵ6F�d��Y`v��ӗeqa�Z��^�F+Âw6�|�Wq�����z-	�o�uӭ�9�]J7�*�]'�-߳30��PY3�24����a��0��c*�4����5*[����R�O1˧^������Ӯ
!�%��*��UX��:X�PX��7lw���X�\=T���a	����B1P@"���=<� P�_#���7�>{[PRc�+f��sjL����@����h�;�8�v8��s�D�����C����C7�T�n�f)����9ͮ�5zi����>��#!:�E`>�7:+��!i��)�ܯyaV�;�5��+Fq��S޿T��1q�Gi�b�>ܑ^�0�t�'�z9��U�b��j���V�)���A�/l�^�a�B�F�F1�\�p�䘫LR&u,��sy����
oH
�
��:�y���H�¸�53�V��P��z�yu�ɒ�� {�v�X�޶����� ��7tX�T��Y�{;!.��-��;�l�|򃮹N F�<m�Pn!k�V�ulB�+��}������r����c]5�ؾ�z!��eorq*�$}���5�$�Q�fbԱ�a��EfC�S��u�^���ۄ�LT��e>�8h���*�\:PY%T��3.�"�i}ή�c�!~��.�:U�8�Y{:ƫZ.k|p6tJ�TE*ΤF�|�4D��j���Ut*5�
v��-�Zҽ���;y@[�A�1�am�E;��7��Dhg�$�<�b���,_�F�?sљ�Z�]�7���lZ0�0깛�h&|v熮V�u��p̬�c�1�vv�Ļ��[�W=��-J���8��(TZ��߶b2vy�η:�����NmL[[GL��86 ��j�q��`�4<�S#J���x���_h�]���u�ru�E��]��5�T����B�t�;S\�8#Y��}v�A�[u�5�4�ʠuشxK὇:�#yy��Dݞ�c�v=]�hl�T0�:}�m�Ŋ�x�7�<��گ1\��ci��:�s��$��Qv!�3�w���X�[�r��`0��4�x��8��EΓ���"��~��k�
�S�1���cd@u7�_!3b��rA�p����Pϭ�I�\�d�=�ExX�¬���p�kW_}՗�fZ�K\8���ӷ��M�)�9Y֧f�huq��oMӔ݇�ڐGzpZ��;�֤�}l.��򪪏���bR�w�z�L���@xc����c �:C��P�s�aD�Q#�٣�7[x)�{d��]k|Eu�n;�s(�>�sp�H����/�κ�@Lɬ�Jln$j�*�{*����U��B$2�C�^1�P�VK�r3��b���7�l��;����B�JQͱ�/I����0�/)�Ӏ�xa���O)`�a��F�r����d��毮J��Xb&洒���u�>��gјm;<=�
B�������`��N�݊C���ೢC�
7�TT/���e�p��c��˴2�hYS�f�����g3�A�8	Ǘ�yw��w�f%�*z��y�f�ôr����",S,p�;P�97ezU���!Q5qP�p���A���3�ݞگ*��6Ìm�K�Jq}B��'[��e�+�����f,!8n�b������b"��2o˨�^ח������QZ�h�`)��x@��\��~ٯL@��P�[��^� c�m1�Y4�|�@߾�5����[��z�e����1w$�XT�:��֤�\3B�*�(�:�!]9_!(��4�@��y�{�K\VE�Ǖ� ���L��D���"��s�[����M�ӝ��>����=ڡ�j.�\���*4���-��p8$t��i��$4����^��'���7o�T��"�&G�O(������'(�<sH�(�tc/ک���m�&q��l��!=�������׵�s�!�<�^���Q���M+>��x���yW���'��K�SY��O0��>�k��'�7�Qf��A���؈	n�nv���]�$/B��*Xw�(B��O&۟=S�f����RYJ����b���X���=ez�2�]�Aw��n���Qs�q�8O�D���n}�[��p9W#\#�A�\�.���W�F�����ڵ�hz-',�Tqh��^���f�
��H��b45�Vmw;��5(y��}ƭ��ԦWOo]��
���SuG�-����>޼U�l���y�/r[�����q���F>��Ýև	q�\�qye��]�u�z��;������R�U�pjy���� ���V�J@������a��D{*����vwF��7�Ry�G���#��*�]1�`�i�w>^�A��獵Ex���{��YSɼ�S&��oeAG:��ݹL=܊ҋ\gx��Օ�����WY(���O+�t6���J��<K�+����l6��,nڣ�x���v��� ���L�ōݱN����7"�nR6�n�J\�A�,�.��R9�'�����u�뱉r�==��䩬�,Fɠx��C���2���Lid�ג�E�:ˇp�T�܁�w׊�b�n�Mġ/Z���g�_�����B�xO	E���c��"X�BRC�'�a����U����v�2_5�YM�l���9N��E%�I�A�� ��t��A�ޅ{o��U|��j��!�͈"�ʜ:����I�ʡynUEVˆ�~U�^ޮQ�t�˽)՗\�vh�_gK�!��A�*D?u�/,y�a�փR�������ղ�xչ7U��=@"���m��a����l;銌s&�eH�.���
��SbS�}4�`U�J;�N*gK�4.�uC/Ѳъ����I����cx���iٔM��j�r~�e��e�b�Z��$�Ά8{j��X4V���Sj�xh1���"쎔)p���r�gzթi�z�
�]U�9l�Q<K��W�P���,EF(�3����a=)�V�z�nPDĄ}t"�)�@a �*�*牱+��ҭ�Fǣ*������K�gGó6)bU�d�6�&��&�.�7��"ʆ�ܧ���e�[��K��Us�;8r����l[�Ƀ	v���}�ׯx����u:Ky�*9qp�S�
�D������:�+k����k���%����Q�Xj1}PD�t"ۭ=Sص~�z/��v���q�{v%��}D`M�1��#�0��?C6����,l,Q��Q����v.�땹��*:N�Jts7��,��y�3�@��E����$f�r�31�s�$wSJ����:O�<-��D��0S��y9�W�lU��8�%�я�U��[ޢ�f��TT�)������ۃ(el���hl���](��KF������
@f�{М�h�5\�^���4�f�3O
�Ȓ��40Qg��S�}���Nq��c�ڱ�V�i�C��h:�xk�+uO���h@S �����^_����g9�&���ؕY�Ώw)��UX�,\)�""��|H����{b)Uz�J��F� �P�Uq��Xxr��H%	���DCv!m�f�˸��ōpH�T�����������_ME8�K��J=1Q���mSg��f4C
1��M�۝6�T�=GE,j����C�#Ni�����A�rz���iw1;<��[-�������!�(W^z����6+�C�	��nL���H��T-f;ɽ�X�ZIV`���ʁ�1:d���8/+R�[�O�.p�,]����7��&g*�w�D��lBkJ���L*<��A3F齮�nQi�w"wN�.�%��  8�K:��Ħ[��42�����Up�3{�V�,��<�^���0��L�7�aVˣ���=���u�f��ݻ�^�g��g��}��KJ��7��yX��L|��8\5�֕of�f�g������Y��L�{���lRp;._��_��^��U[08�@S䍺��^��(�+���wH��U��ͻKSg(���zn5��"����*p!ee*;�� ���F�uDT6�+6�����Y����~s�eK�z��k�����b����+M�yld��/��	U�w8-B�Wk7f����w��dL!�;�q|�0{5��D8x��d:�PY{,�W)*�븐Ա-�74C'F�?:j9�F�5�j+�	:L��r�E<n+q�mW5l�ӓ�tz���&/I����iT����L�p��U`�t,k2�a��o��8�IN��C���1�+u<M��!���a��R�����5����sDt�lvE5������q�7�1!?$6n%�G\'�$Ֆ=½3,p*��;�x9A�K}�-{M�D�����>L��G)��Ga����n�@���A7|����\6JWyEՎ�O�hiA���#[�Gp��^Z�}�ji�P;�ۮ%�ޘ��[��X8ё0���/�0Eo:,F�Qqd�%���ծ�f�D/��������ң��Ε�Zj�._z=�V�ç������#��߽ҍK���W��0й�u�&,*,pf�c�g4|���z_�N�<���ߢ�Y�S�gO���i$�C��Y�'�~�#�ٯk�Oa�2�x5�-[��R��,�4{�j��>v����I�c�7�T�.�2�Yu���㠨X۾�V���[��xX�<�6]ry�g�������1ԩ�p�|��>��|�g1��qy��xX�\����9���eB���Rr�!fw֧�K���rz������_S��y��H�{���-�o�5�֐��y��6?/��tiY������U\��w�V��w)ɟ?>����^�y:"�Yz25�D��TGY�+)�uw���-�۔D�B3�Fgy8}�W::9'�℅Q�������8�1����3�%�J��;�X���t�.
F�v^N��6��!Yd�b�*��GJү��5�^��s��9\�iV��K/��Bj��*f;�vϴȐj6�3�(uE��r��p�T#��}Ƕ�*�$:Q-:��J�9��ՠ��B�=�[6)��+c�2�>��=��<'o`N��>�J�c8�yZ�]GD��;w8�ݩY�V�m&p�O�jwk
�X4r�59n��U¸S����e��V�wQ�|᮫I/�މX�mS��^!_mX��gG�=�����}MӪ��|B�nU�u;�Õn������gI��[6���v�S�����!��P3�B�d_ |r��\$	��'m-�9�'��^��D�< �O(np1JQ<m�1���ٹ*�9���0�hs�N^	y��v�LN�rO�vC���1Sʛ�ȗ���d�2x���\dc�,�zyu���cꋄ8A[�w��2�WM���󤪑x�,�̓r`{��t�l��ہ�������ݯ��:�?���O+	;|?:�����BRC3P�=�3�U�0�V�I�+)X���;$��n$���>�D!��9w啕��4A��@	�S�&ң=1LmF��v��n�M�O������zڳ3Ԉۇ�s�eS��\���*�`��R!@��v��Vv��X��xhi5�6�u���W�eH��H�� ]��^�'��TD��:M�]���ĘvPz�7�"qa�nuu���X���hV�Ʈ�װ��R�w.=�N[c=2[~�c��@ޕ)�ۿC'v��>�=�uyw�6X�vT��<��!s�&vNe	G�b@����v�m���
���/���$��*P̬�*+k>��%@��u���*P@�����Z������I߿}�[:�k\Z�3#��+.gJ�8>�T2�e�Ez�md�T&�#sō����Q՜bF��/�uX�G�s�t{7M�!gQwT�W!TFKjXzh!���`��^��0�;��Թ�E�#��6�)��Pd�Y�U�*����Tj�"��c�x�u5N�7�+#$^��c�f:�b���x0�F�b7f���
�䲺 3�
�\p�^*g��w(6b�tƣ����F
M屄�RU鐊�@s�D���������D�+^�)-S�Sb�e���}Y�K�	H����:+�fĊ����#�����a��B��s��Uf4E3ОndF��z�Rs��Nc��'$b}w#mLĺ���2�>�tU��t@Dªʂ5�M�"�/AB^,������ʽ�R��Eޅ��ps��T�W���H��M�Lpc�axm�hY��^��p�B<&yl>�L�4��Y�\���.vh0��-کo�C��5���;>$��y�u��5�YXe��7��,��B0N�ώ`��5�i)���<�}XF�״�������郛`9��;�uegn�H�eK*:�A�L���ly��ڗ`�c�]}��F���2|�:S���]���4S7�� M��Ɔ�1I���Y`�ї�u27&=�#.U��1v����8����4a�g�[�a�ɚ�_%���"Y9Q�n7�u[��ÌC�����:]G��6�s�{��^�Pӹ�������S�=�n�#�?�P�� �R�g���ԭ�E��E��l+�n�<0Aζ<�{��.;���m�i`b��K�;r
�(0�����JqfSK5H��*���u�������4wS�7��qо�G������Q��/h������P�Õ`��I�`m�j�����闶9 ��H�t*�^�����o����Bv��/���~,�
������nv���P�`ޢr��޼6��aa��i,i!��,R�Ȁ���1#�oλ8v��]�t��5-,�ι��n��[���`��#j��ÄR��cL�u-	ť܇if���N��3:>�Ὓ�n&gK�M[�*�Z��=]�RﭫB��[�V��I�d�����%��D��]��WYQ�#|>�)�O����0S�s	�u�m^��}��j.��g)���RӐa:��9���֨A0Jv�ٙ��Nfp�y�1ZfͲ��	��lĺ���*S�/ᓝm�7��Fp�4�Z�77'*[,�n�8���v��\��gr��U�vp˒^�(�8�Ns�K��^*3[S�����sF�m�{�f*�-Do�%sCm�+4n'�9s�C*c�[kϜ!��7�K�S�È\�s��Y��6C�}H���n��4���I@so�� �}±�Q��^&�r�����V��H&v�V�~�������!,�O*����n�Q]���k��	C6��C!�K�?J�⣂K[�t�s�4p6��[��F��-T���0,�JU�>*�Z�C�Kv�>]0MG �� ۨ�ٛ7^od�O�n������%Giz�<�	Z�7cQ��"�WG)B�h���\cGC;��nM��)kegƯF�-c�ƞ"�!S�=b��fͺ\�31�����	#�9"�K/2](�Aw�ݰ����m f]{8ժOE�SB�z7[�@;Y���J�:��F��o%�I.��3ֶ.Wx6�=�]%�Xh̬�b� IȰJ�67�N�b�XWvu^�qL���#]�iL=f�ih�s0�2Ξ�7qm��F��Z�b<!����|��;��'0s�|��Ux�:c���g������Z��n�_G0���;6N�8�%wS����.�>�D����3���j�̠���2�|%�^�*r��I6p��n�`buҮ2�m-�k��6�V�2.Ul��&raW�jv�l-�Wv�{S���~������ײڤR�EE��eF��°��7Lf2�e����*"(Q
��6�s��؉mG3�EPEJ�,��b�,��kUl�*,cY
�\rT3�X��&0QjUʶ�([UTX(�T�B�"#PKh��"�����ZQb�akm�[2�,R��2����X"(��� ���J*
���P+UU�-���kE���XdPc���`�T*F��$�R�Q�Y���l�(�*#eV
��E�Z�L��5�(bQ.c���mQq*8���V(Z؈,"&R��-Y�A���R(`�"ۙ,�+l,��`ŌT�jʅQX��e`�F#""(�
��Jň�Q�0eATA�[iV��mL��b
�+1�1ĬX(�q�H��*�\Q"((��k-mdQb�11��[U��*)QVAd�V*"�,�X�R�REQR,1�rʊcZ��r��}���{�߿ot��-n]9i1�qj��I�=�R��M�=Bc�K+��5F�]�NA��lQh�
X�P�)Q�k�ވ�RV�gr�G?\�e�u�Ȫ,"`���n�z��ȏZ�_e��L�Z8i��<�܊zމ�Iq�FW�ݡc�3+n4�]��pŊ���8T p�u��<x���C�;z��e?E��c,1�X�M���D��:ډ�8y�/H�hH��`���RϘ�ȩ��~�s�{"��q�F�q1;)�)\�M�����a��$��i��No������wM�Y�p��@Y����q��1������+���LOQ���f_e�IoQ�y��%�̭��Bv�t�{6�Jl�.��J��_3Y,H�h�o���\vZ�
;�X{���/һ/F'Ԩ���5�#��,@�L���UD�;\]�嚛��U���T-R��k�#T�cD������Gq�Y�% �Dvͪ͞��<]{��{6c{�;c�d��`l�]JϫݥoM���V��\�=����8_n
�W]� ׷9�]z�"Z��O��c�ӟP��"uL��L|���^\Mt��7��@����Ja[Uy]p"��uDm%�s�\bz!^��χoh��i��N�X��Q���<9`���+hJ=WB��6��B�2:WϮ�X���p��̭W��4[�f�O"�V]�} �{�O���J���Q�"M:�I��z�Np7��V~�z"����y7=�Sc�sVO
�p�oI��ŋ�S��w�(W�'�$�3*���c�KoiZK����k��t~�H��W��9����h�8��(E���tƆuG'=��&��4C2������M\������b�-'*�|6P��<%\�3��0�vx{b'V�˃Ҙ꾛��tĢ�c'�yl�e		��c����6���8_�����J�V�Ob/�E^)�}FJ�g���ib6	�q��K�J��y����&��Y1�C 	�r�G<�Ub���*h���ˬ��:
5�dΟ<����[!l�y<���8�}�٤1�L�޼�oU�U�R��VNc�C�����|��*�l]�gk#�O����Ux��sJ�r��ļ����+g`�������Ɋj@�q��t���Й��s��ah��.A��A��P�v5�{��j�}5��Hh�]�9�`e��;�7�^�|�F��?n�%
f/9ք/��Eƽ��~ŵ#V@u�x��>�7��p@'"��n�ҥ�jB�Z�h�C� �T�X�8ͭ]A��� gjg�Q<TI:\��ٱ���uM���A�M#��)�=�f�i�-�"D�s9�M�]��ܬ�U76�G��3O0���2C��1RBEֆq�s#3�i}�7F��;����v �-pEo�4kUW���aC�xS��,���G\b�:����9�D�Y��N�
����������7����	
�S�l���1��]~�Kmh���V�Z8:���}��)�_�N`dײĤv�*����*��Z�C\;Db�{Ӑ��Ct�Wm�/0�iC[m��Jb��&6�]se���aP���ig\#�^��N�a��p#nlKW��] ���#*����_��EFt��!Ҽ&.	��@\]��!�],�ğY�g��s9�
��qY0�6난��uA9uB#�uHB��l�M��G��O��5����箱��!���Q9\��%:�\'�f�JP�پ���1^�V����Є��#���5�m���Xw�ޓ��u��F+�ʛ��Kʀ+��I0�'��{"b�X�GkQ*���,C�6/3�C*:&�N�O�%T�stt���� og���2��rL>�a��-y��~���b�`�6�������� 4��5�=y�9�F^N81���uzg�K�����gdn�+�N�5?�I�ӫ�;�WUԥ���AW�tA4�3Cu����1ݩ���[Y|�	l;��qZ%r�Ŷ����@"���!�Kp-�<��[�B�I�B�q�����6�_��Ud$��k��{�c����"�D��Y�^�ΈB��ߖVV0j�n�bλ�S3ݱu�S�J-Q���C�GK��DL'6 �w3g\6�m�#^�j�&�r9KE����W�ӎvɼy�U��3 8s��G|���gA��ECYDf�@`ˈU�!l7ݱ6��G^ކk��K���8+u�EL�<7��Q�]16�2Orʑ7m�YG&L��wIַ9��J��k��d=q,>b�v�g���H�ɵ��I��������¦i�l��z�ܶ��)���d�)��k�/N[T�W!VK��L>�:)N�3��Zv�P�!9י�)�ނ�u����RX�I(<L�w�ZU��u��Rxz���)�����V��:�TG.�M�z�^v�E+ЋnC1A�4����O-���_#<���}���e����q��.mG[��5�%���F
M屄�RU�L�U�1T#�H%.�sTţ�'�m6��j�6t%����Y�}R��Di�T>��͉	̺+��3&�z���xY��z N��	����c�7� �e�	t��ڽ弚3t�@5��H�C��q"s�Ӣ鞾�2����̭���$��󩠖n����VS:y��3M8Q{}�~ެ�Jܬ���LC�,�)N�z���\\+$Ɗ��V�ǜ�#8	/b��j<=9�0�h��V+��:Q�ѓ+9�>t��)�q<����fHT8ڥ��3�g_�@���N;2}\��I�n���E@c���C4�/�u*a��j}S���u�uh�m6���ߣ�*w���h���^F�}+���Y(��xR�{+��
	��2f��ĤvN�N�%p���6h���x�m�t$��y�e�dXM*���I�m��;��q��Y=T)�<vWs���H6|'ܕK��"6J>~%%�U�֚�3��_$r���ER����=z��B	8[ULp�f�m�f�˸`Y��$�T����}@7�g�d��A���>����E�鱂;li@LmSdq�Q<8C���o���3e��cYY %�[j�&HPpC�ڑ^����P�;�iw����
�[���+�IȹǬ�ھTW?_NmLZ{GO���{6iM+�|�:V�3�~멝�oΑ��W٧�9�pf[�SE���;���N�*;�+�Ɋ!)�p�P��J��e���p&I�P�;!�͡�8[�����W��:(J>�];�"�32�m_�8O
at�W˵+��m�ͫA��O�͏��l^wR��Ͱ�*��>�H
)��ћ��+�{��r�w�Jޔr@���EDa�����1�ԥ�Υ��}��*Wf�.�Loݵ*K\;��]��!>�Edl��P��.LP���aMNl����,�t4��S���mB�j���\��)�.%N,��Gq�Y ��uP�ol݄���%6z!�6��4j�P�}~�ҷ��HL^�Zn[�c<V�HY�m��u����+桛�g�<�e���}�����*ᩬ¸�S=�徒!�
�N��S꾥��_J�����#����J�ل�%a�O.0��c4�U���ah+��]�N��d.xlGu��	)�\w����v��'��75m2��k��F�.��'�wM��5�o�s�=���k����N�o��"a[��n���}2�c�ZY�u?#�׍����3ʹ�r�d]²�7�b��.�5'���4���m�Nq|u���\3:�g��z��.t{���N��*�K5.�	TPbᛣ��T�MK&0Jʌj!C�6�(R�Hq]B�9Y��΂�F)�3^���%�/�h���y� �������ޅm�B�fE�:�b�H�}"|�x��k�����-��l��Q�xU�b�� �>ᑉ��;�����׫.Ws�u��k�d��k�N�ޓ��7ڸd]կ0k��c��`x�9m� oC�d&.f�>�����}�%���1�H�,���}d��S),Z�8Jv����I�>Uc~N�b���W׽*OZb��F�tBq��bm*��������ٱ�xO��a�@_�?
��.�N�qu�9�f�%�d�E>�
�]g�jp�{�W@���岐#b���5��xf�Uݚt�f�* O�9F2���5�1���Z�yQ���u�-����<&��t,�ݚh�bnj��g�n�8��[Ș#���U^�U�5���Mu���Hm�#YH�b�y���-o���y}�OV�,JK]��:;�[Z=9�%=��s�r�6�����N�0iZ�jK\��Q(���r�07P��pDr�/W��kG:�Z5ѭ�=x�?q�(b�az ^�|m�����p��K�sCبj�	�G��3�;�W*�u�0��Ar�&��f�V5��\u�Qp6���&�� ,s�p6J*�gP
�Ҽ& ��p������|�3N`˪�\�F�p���s�K�Ç�.�k͏�`��T/Z%U��Gy��fR(��wxjKq�t�E����r�q:�o@]
A�;��`ƌ>��X�&2����hw!¤���Z�eiKuZC�f 7��Gz��U�M�S���9��d�]��
o�&��G�>ۨ{,E��]�Jq�;^-�r.V�Nv�����+�d�ʻ��K�|퉎{kʽ9\��u���L�#=JQ<m�1��~���2�_���un
�90�����lO�9�>��0��1�b�'�73��� RwRL �,\�� Ws���$��,����!
�#�מ2�W�&�N�O�%T����B����)U7��*��r���@�;�~D���]F��`�'���e!�t�( ������躭�N�hR<�IM��h�F�9ĎXs��F�;�����j��j�n�D�Y���l�ȳx/m&�� 8��l�Q��DL'6 �w3g#\I�H
���ۨ]v��b���k��%�1��вe�l���L����s���"*�#7�0a��SS�|�䅞�\{�6��s��>�N��,�g����U#<7��0�'}��d�H!3Y��Ec�U�Y.w�M[�[~j�*�NXA�tN#��^�T2�e�DpN�ad�V�1.�≾���z]�:J�*�ࡼ~u:��6{
�I��%�x]C�}+��U���B���c7�;��+`e�~�@$EjᲜܬ�+ӠD�����b328�Ɋ笓t�ؚ�O%�]��3Z����+"��ϝ!r�`(mu�3�e�t=��2�u�N�3����r:i16t�ݭ	�Z�ٷ��ur�b��p/Fn<آ�/��L�O^^�֥N&�Q/�"-=sq���!�j�B����<��ʨ�I��Pa>͹���j��A�d��%��n�뙎�����E�!���U�`\zVW��Cu6f�j��];�Tj6�ar��5���u��#y7��x�
J��!a�W����FT�K���"�ӵ����C.m���TF�t��n�K��i�_���ؑQ	�:+�Y������jh3��ܱH\u�`�~1c��%��������cbS��o������/���	UO��(Yed�� �%©h���5�L�GO����2��珵�F7��4$���t�V�e��rl��h�;�q;T���{>/�]>������k)�}��`�=:����ܕe�TĲ�!�D1P�����=U^�7����{[j�����^�\}�Ui:ő�|���8��h��J/"�NU$>�*"��H�?�-��[���3�˩+Fs<��9�(A&c
��v���f�m�f�˸`Y��$`Py�ׁY�6=��\z����V���&g��w��,���B�[��i�3���WTבټ���Y�����2�v�	�zf��N��''�;Rg-v���u<�ǴYj��T�]�%���7�զ�a�k��iK�P}�6�.������˼Տӄ�X�����{:��,o�"�D߇bc�Ĉ-L(��`m]�[���ϴ�<F��W�,h:Q\=�,m�Da}1;)�+��WvePI��R�I}]˟Zo������*}݌����-h_��1�SJ�o�_o�7����NC��MȹxkL.K�9�!�K�/B�N��zf*-LS~��b�W�BSd�B�_���5�ME���z��dZS�c3f,?.��r�+��'�����5QO�7�S/%B��b�mN���p�F�D?\�.�j��G-�W����r�j�L`�S� �U�n�Vo���zie��x�]�9 qyN���p��Eԡ��}~�ҷ�����yY��ю�����s�Yz��	����<l��S�QjXY��C���/�Əo9p��t��3�.�:��e�D;���C ���d�N����V�pT�b�����(mO�%�%`!f�x.V�����;�)px{GZ��ڧT���i��>Qp�m�U=b�k��fj&�W�9獨UY��ATͼ�ը%�t�m��x��e��%,S���R��i�n�B��S�*\75+�f��nr���L���u��lE�@�ӱ[�n�b�&�����vDOO�����s��
��@c�(��wX�'�:�����z��cmZ=M�{{�V�,��o��f��Y͎��q����(J-pP�s�u)K/6�N�&�{ӭ�\f�����{j���O�]�K�%�V�O���̗(]�Vz��˗�hs�y/*}1Q��E9[��ۉb��}Q^�ؽgu�փu�^m�8���6�	¦\�*Wp"�ܾ�-!/3e�hZ�S)��M��Hٗ|��^m,vi3�B|[�NUd�g-傆�@
��qw鹌��%e��D�`������ ����V�� ��<욲�i���m��](mvվ����cX7s�c�T�"{4����§v!h,OF�7f��g�)e�h1��d�ӻX	����DЌ��H�R;����Z7�k�9�Դő�8��ԟe��;b���ĈxZ�;�t�n�5�;f��FL+m�M��[�u��OHڗ˨����Q��A�qZ	`
����%�5�)uՃ}�]��T�#\0#�܀�Mkg]������;���ub��sշRf�zƹW�^���U�]�����!{V`�ݐ{�!X�p�.�H�|y�ڙt��?a��P���HR�WR�{���W\�.؎f�][��N���sCR4Ƃ�Nu3oz�ܻ�k��<.�V�F�����tԺF�k2nس쉌yZ��v�IR�G��FO{{�5�Rͧ�]�E�1�I4�l�Pn��qo[��S3��y��,L�Ol�=���;%Q��S�U�!��N¤݅yÛ��z�l���gNeJ���2�tʓ���n��Xd�u#zS��ݜKG#ڷd7�@����Ky9Ӷ���.�no[�o���������g&���K�o�r&1-��:�ͽ��R�բ[\��kr��V*���u����y��8V����ܾ��_ �l����̬��E�7*u��&��ҕ�b	�W�X��� ˼�P�i�b_ml�׶��	h��v=�S5i2YP*V�N���u��y"s�ؤ���kՙr��7b4������f��;|��ءR�5�x^�֏Q�c&5/o����5��������m�y���� �h��bq�߈�o�T8�I���Vu����S�ӆ��n�;�m#2s��em�S�5��Ɲf1���Q����%�����7_X��oq�gL�	��1��5�L-T!@��=v��.i�{�Pz���w1K���eȸ
�I�"���f����_Z���md�1��-})�S{A�v��Xd����z���9Z4���O�q'a�K���[���=�>=�安�\R�җ��74��ų�i���'��A���7�N�e3��鷵y�r��C(b�]R�P�)�p�݅�����E�s���ه�XK��(3�7uwNĺƈ��eEX
#�fQ&4\j�
�-`QX�Ub��CTX�����EKaUDPR%h��b��ш1V"��(��R���b�B�1�����9j�2���mER�D2��Z$�F,Z0�j�W̲��",ĩ����X�Ҭ
��-*�Vc0�¬EVQUVe��m���
����ʋP�
#r��	m��H�m�W1ɕ������C,b(�Vնۖ��e�T�T���n6�&"���*�1����L-E��XV9���ҭl�U�J,�p���D�m�Em�1ʣj�[e����Ĩ�2�"1�i(���"�"+kk���cAUd���j�21X($\bV-K�#m\��TjQdLV�����Uq(���Q�b�5q��B�QX�V""�-�\B�kX���1X �.f
�2��8��D�PAT�EF
�#R�b���X���-������m1��V�J�[�es�5dW��aə�OB ��S�n��]�e����Ϲ�������j�o��e�Gwk�^B�7���ob�������L�}{V�h��t�Ju�2�n�V�x��U!����0�!��8r���ai��;ftl��Q8�&:�l)b�f(;����ļ���yrM�=�}3,pZ6�Ng�+{�SQ]��uE�ƾV���C�Շ�,�����p�E-���'ueE�sL5Tb�����&�B�QX���wg���Y�S�gO���wL���YH�d�>�{�V��i�u��EV�ŃE���\�*�X<��A�;W��Kq��x��:�ALsro��ў�	��=͑�=r>�<X��A��<�۞O�
f$lZ�1���t�*��ԯ���� �D=��&��}½��7�F,���I͖��)�r� ���U�����/�*��\l�ˍT��#l�_:Ї;�������ڑ� :ѼB��4�����U�>S�~��=��9��U^�r�ߑ�^����WX7���G���}2�7<�(��#h�=���Wx/�2��(�L��FJ{6��꜆a��]=^F{L�o9�z�ޔ���LU��.�ǐ�d�.L�Ú:5г����K�u�[�(��pt�#�z���SW�.��u{�,ۣ�ܘ�T�_A��~%<������C.v5�D	45�٨�t��٨Xf�^��a�Yؐ����K))4��b�txg�R��J�Ĥvω���E\<�v�~0�a���;��92�r@��7��~�{�W��\�d��:(}΀|��jQ�&����yH�����[Ɣ�!��߃��ƻi7x=ac�+%��t�	��lu���*��M�X��k��g5�G�ͦ/��4$炔� �/]����.�!�T��1�Kk��vQt:�8=��-��q峕̔�ОP	�e)D�f�j�F߷|
����<v��V3 H<��>��èu�F)ng��T ��;��
���s�y=|0s�+m� ��B���!_�l5�tkȃ(etM���[����8.�Q]����X�_N�ɺ���a���߽�O�ٞ���]F��E�Ѷ��{)�p��L��G&M�rǭ�V8Ȳ
i�
�<�!�$:�R=jU//����2�O��ۿ�k�Qn������ڵD��̀&u!|B,��"4 ��<�î	|U]�>�j����J��y%iSF��S��1z���L���.;�tv�餚YCw1f��nIC�Y]� bƮQ��mv֫�n��M���w|h�N��*P3,���ӫ��͐Ì�l��qm(���MUʷ��\�L�s��x���'u�d�����>��x]w�c(�AdΆ �5��F�x38�A�*DW��#4�Aܒ���brv�cC;0	�i܃�4#"��^ƺj
��0����x;�ؗwu����1�7�?-��֣�m
��^r �d핗3���9�x_��UC��GB�����{\���{�q����xkQ�+kD33C=3=�
�[T�W��
Q�y�k���o}�F���?��|a[w��7���5M��M���&U3�z�Vgg<�S��F�9��kYV�18u�X��8�3��:�c�����f(0�F�vX��o��+��ۑ��9K�a�^T.5��#ǱD�~��F
��[�RU�C�1�y5�Waܔ=sU��΁*���K����5�*�d4զ�1�6��s/A��͉������3���n��,�l6k'�!n�0CC���seY��'9�\JuO^,�[C���8������e��m��n{�\��Dt���<4L�Wu�<|�<@X�M��[#<����[���U�԰k-b1�o����Ƹ[ ���jze����� *+��ˡ,Q՗x7&e�pj��1��6�n2�I0_q�9�p��+��
��wP٨�uSP���Ѕ[!���m��̱W��W6r�\A�����:��TĆ߱e{�� �󈁓�U��e����Ѯf���®I�2�{�^���d#��Ű��K��y��^P�7�KI�m�t�����m�����V0@o��#wޛ�H�g^�*HB}�%�p�Bd���BJ���z�!���9�����N0����pJ��A�����v��I��mݱp �[PY�O.��8b�ؼ[9S���CK9�=1dHe�.��йټ/.wM����Jv��/�8�&�p�#F�[���b�����t��r��D�Ƿ:n�h
�]R�O�4��ۋ�!�"Ϸ�Kw��|�3��9Ԍb\WN#��=w�l5؞���Cj�vC��t�S#J�o�_X��++q��^~N�g>h!�q���],<WXy:�xdq�J�NTw���X��LQk|!�H�z֨���3Yk��C^UCW���޺��Pa�A���z�Tyl��U
|�������suj�j�����r�W�گ1�f)xq�❱��*p!pVR��<T6zܵ�BӘ�9����.T��qh�CEc��ͭ	:�F�J�]�*�U�S�P�ڀ�v������)�SCF�v��e�H�\�`���p�3Z����T��)w:�G"��3��R��j�>{��%�2��I���9%H%��_F�=��k��ڢ��e�����z�Q�&}F�w��k�Jޛ�b���V\U]F1�r�*/c	+no��JÂ��C��2F�P��&��p�E�}�:b�p��}�Lͧ�M�cy*T"W�g�ם>g�I"%㻅�uԡ�zHB�xT+�}zM��ŋ�������v&YS�op^��Y��&g ��'��1]+�#!�h�F}�[Y&E�="��SSlr��Ea{Yz��u�b���ưp�:OD�:s�ހ�m��NgI��5�#ׂ�p�|���v�a��ٿR��tsa��1A�BBf�^TrwRNŖ=� �5I�;D�{�$��A�˻C�l���óZ}�΄#6&aWK5-)�s7FT�L�S�Mu4�d��\+ZMXC����u�
�v{"�|o�"���j��:d��Nuһ��u���:�Nf���Μ��{A�; ��Lp�j���'���*B�����v�w��C��|K�!v��p�b�Ph�13������p�:1���Z���o�e��;緦�S�z1Tॷz���W6+g����-�7Mb�7I�<�)����{޲�]v3k�G���]ܚ���R��l&�v)Ͱ�ov��L;�9|��tٸ���
����,����a��bt���|���a���*ڤ�M�o!3@.}Z!ʖNB���Ӂ��#L�M���G��O\H��.nwj��t.�	`�1� �ښ��l�1����1���E�^�Qœ#�B�&x%q�J���K^Q�y�ǲ���旱�_FБ�^�g5�X/(���ٜ{�s=O[�lͤ;��F�:.�rX�s��;�#����Y)��7>z�[ۚ9Ճ��U�ު��W����&(����\��ɸ�S�^��GJҡ��ӓ�)�������q�:(9�Vl�n}�8�҇*�k%g1�C�t�Z�5[�M!<)n�'t>c\$�k��g�+��tG
��x��F�Suc�9�%p3�n��1uDN8Z�p�W�6�/3j��ͤ.�ƊI�9��eп'N�zƆT^���-z��3��2e�{�E��1ya�>�����kʽ9\�ħ\ ��@\�j��4 f��v��I�;�M���:����+�.�WH�eyןժ��ܝ��a���ˑ�<M���)^��c��wau%�l��3}��A��߼�ŕ�{���$����Y�FbW@��*<��`��N��\:ج����E-��:��\�E�<Hvۥ�u��oq`�2a+ZW��`��璟�Y};Ss9M���'+(�����j�0��9+�O\����I5O!q�.t1~ã+��p�:1������{�����b��Z�����p�|�ʤVC��"k� d;���g�l���f ��s�d��N��ڴ��ok{�RF�"�AC�䤇I��x��9�*�eϻ�i���5�(�P�qp��ˍE�A���S�/�B,��#�E{�T�q$v_�U ���<w�8Jܓ�pj��C:����e����b�A�^�l�p���gA�*Di�s�}Q9�&t�K���D���r��A��!�k*˸�@mAA0�0��7:�J޹W5�r֍+wʊ�q�6Kw2#F���s�g쨖
�kGg��{��|�B5Ӹ�#�:��O�j�0z�J<��
�s�t~�n�9��_�;��!y�g1k|\ʇ}3mb|�+��p,7�XZh �%vdBx�x�D#A-�I�ɥW#{8-��u�=H.�y�T7n�B�R�V8�3��c�&c����܆b�0�G�!9��gY�+������b��~��[{���`�ļ��9^�q�r�.�����!Ѯ�����DYkf�����9�{܇M����f�GuC/�.\��s��;h����������쾕��u��A��{WD!{O�E�N��j��9��-=#��#���� �,��\j��+��5�X���F
M屄�RTn^�T�ȥ�kP�Q�*_�@���0��y�c�+�g���F��C�:.�ٝ7�d{��맺Q�x�3�>�>�Z3PW�1��;��~��9�bﺅ̇o��}V�R��V��ݕP�㏁�u����2Q)�<>���(���i.u;sr�wr�Fp�S�ظ�0ً�s`u�yT���@���]&��6T��D5�b�K'(�쾌�՛���ƈ�tgg�MR��^n��ה,���ZL�߇J$�[`�o���j�Ėg���Q��	���cE����e�w:�>�Q�ԈٕT���q�:�}}��f:��˟ ����;����C�pG#�<�aS�Ɠ����w<��x��$1EH.�m�q
��bt�7X��5��;��q��\	�q��^���\v<DX�U�J]S�x�0��Z)�ƃ�Q\:υ��|�i��Ԫ�ǘ�L)���
�9�(���Zqub�`���vW�F����R�suP%��sn�Ř*%#�j*��B@���9��1�'\���U��1G������9�9��wmXs��-����j���L
櫘�. ��c�#&��Gm�wL�{�s����N��	Ea.!����7�Պsjb������U� �g��q�����5��Z��gr3�V�ۇ>B%t��]`\��:4^�O�����d�b�����g@��l��A�̆�*���ң~�Q��J:(1ޕ�z3��*+#f�}�E3I�O���y�]���M�7� <,�W<ʿmW���T�=�P�R�*U��>�"o�<Y���9a�V��t۾ *vb:<T�$G�ICW>�V��7�@z`r�nI�Տ0��Z�i�\������Vq���Za.�/�S�XY�0�Q�+2�$'ݝ��j��v������0ywK��"&+�X�C"8YЫ��f	�5��G��i�^o���z���ik��B��6���&f�c��zׇ��:��#�L^��SsP2�ͪ|�7A��R�n�����wx*�Lhb�`�5ʘ���@f�n�V��R\7K��]u��Uûr=޵�1p���ؼ�ED��b�M�G>X��
7�yQ��I7�4�*�"J�@d��J��-���2��㐪���xWr41���>����jgo�C��*n_J�(f7�N��������L��͐A��g%MR�V�;��;���V������uֈ�.t���� RQ��F��'q���@�c������^#��O�|�a�S퉘\Y�z�E�/R��UMָy��}f�%�����������	E[�<̓��O�X��^N�%0B�Y(���Ȱ����[���m)�M�9;f//
�pxi�N��*�x%���3��ic�j���H)����E;���>�{^]��'[;1~ ^�D�s^u�p�n�r�:V4wj/��q�W��'��&�O��Ӂ޺�25d���C��_�.���Q�]e��m�=�A��jLh��.�`�ɋ�(���|�B�F���Ͷ#y'������E^s�:�!'�<�uA3�5���JϽt��i>����׽:�E;p)%7u�C��ܗ�#�>�_N��Hl�dl2�[C�]�%M�dQ���<z
Dd��͋�r8�vMZקX�f�W]k՝�q	m�<3Ϣb�J@Z��Ğ�ɿb�+0���Ʒ\E�39v��8��b�{Ӎϴ'SB�Rcn5PW7�@>Z�4:-%�WQ�>��Vm��eF[_Q+$���,'/Er����ۤ��rnnw�aU݃���+G���h��]
�0c�����]���eΊ�2��x!�eB:�*�K�[-#�p[��8�5ϻ(^���?D7Gv��r�.��X�ؼ@h�{Cq,޵�h�ZF�&��G��E��ʛ�~�f��.��T�n�	K;U���eɯ��x;S��v����<��Īf��3���/im] �����ᓴv��V� �og8��0��m` ܢ��X�|�9��
�s�ۘ�k�O�����N���R��uru�M*k�P[��Em	��S��')坛��7U'>�++gPS%D�wk ׭#O��������|�Ă���;r��nۺq��C,T� �+k����y�^��)�`��V�[�]�Fg8��`&^��7zn(��m�A1ֽ��p���D�g<.f�K��8�<nE��Y����p������b��r�����[� �8w�٬�k(%9�b�Ǫj�gY�q�zMJ
C9ė`�	"��1�Z�|�����c���B�
�_��G��]0�8��Q��4�P����T�����b��:�wH[h,�B��A��F��zˮ�t�_q�+vˬ�>&�]#��q1�gX�,�:���a�R�<�(f
�<��ԣ�lu�{S��W�a:�T�X�Z���\�{�Ȫ��1�ݳ��T��k�)j�p�VL��Ώ#=y�_��T��v�m�Χ�^b��af��=~y���k3�N� ���rr�V	I�Yݯ����Ku,�v��Y
���� ��t��S&��6U^����n��[4��/�Cp��s���0c��p��5s��A�#}ۈ7+MX��ڶ��s!<xl�A"�hjZ�ӏ�s�c�>�O���|
E�ò��"�ފ�Kl4�ޡLj�b̐Ӯ��.�Wy����]��:��<���lG�*9WJ�؄�{n�t���l\�Š��e��z����*����V��Aou����kA(�P���ۡu"㗊�����k�v�+˜�r[�EgfZj�3�]9��n	�Z�a���Ձ,K)r�j��gr��x�Vktá����ϣ���gY8�5�5�޽t�g���Ktou�Wcd�k�+A������+�V�S$u�lo]��yS�<P����4�-�~ޘoN#޲M��`����������y�*�!��Mhi��p����x����;-u;���얓����es���iU���)[v�����J뗧� �Sfѫ��+��)iv�,S5]���.�)7��|�d�lK&�N/��lH,�mj�۷c��=Z�nn�Ά��n]I��<Օ�|��U�PdW�.�v��>s�ARu��t��W9�Bs���9���h�os��Qۍ��Dk*
�QĢ���1�F#e��TV#(��*�1Qb��1TYmU�`��F
��mƃl�`�Ŋ�l+QG-b*ETR+�E��.aTD��YU`�!mU�J"PQ��Q�QA�TX��XYib�(�GY�-Fuj�b��EETb��)�,AUGX\j�������F ��f�T�Q���B�k��QQv�Y����FE7B��Q5h�"�(�`�t[*A��-b
�Z�XZձ�KEZ�Ҷ��b˪`cF�[cmeb�amXۘUĪ�YED�V*"�c*��Dq
�,�pj�Z�5b3ZV�m��V"Qbj��+Z�浚�9Lp���Q"Ԣ6���T���**Җљ��-**(�ʈ��%�h��UP�U��UBձ��*[kQZ2�Y�F� �DQ����EG��z/�일^b��h�w���v����|��/�M���4mf�K&r��!"��4�8R}���`;��t�nθ������sNu׮�N�hǮ�̈́���V�ˆ�EFt���r�xD�w7m줫
�`

�%2�6���Ci�h���pR� ��]P�*�z�����QQu`�>��w$4z�d#m+�S�~ِ���[��s�̔��� �:�9	d*Y�/gg�B�(�:�Ec�4�뭬���܂���}s��t�Q������:���N�$x�f��{��X��t�I�����!]M���N�xe���46���+wS�P�F
'˔�)�e���&)�����=�=w#��?#F���z�O[�?�_������z���$��R%�RRC�'�a�#;$�pJ����n|V
�e[�jF�����EI���h�{VV3h�e�:#)�,��"���PQ��ՙ��F�X�$�:u[MW�M��q7.z�2�YA��1J��6�7�^�c�5STls[:������Q���w�:Ь�;�5�b�=�?�W�
C�k*Ϧy���&Q�N{.X��]W�y�����u��+*kJ����Q��\XP��������lN����ܕ��]³�� ��<hm�#Y�Y�NG���r3�Dt�wh���	���L��P�,�\�v�ϩ�%����u�F�sy&.NZ@�wr<�s�kPɊ���:�]o[B�C�v2뜈:W��_�=tj��}���hxu�`��It2uEj�\m���m��&��7Ō��e�֬VW�M�[g��9��R��E<S��]][nr��Փ�ḇ҂ܛ:�]��9���b:�F�[�7x"�x('uW::g_0�F�D�Q�]�*��¨Ѕj�"�ı��ݱ�虎���X��\7!��(�Yœ������8�e<�/ӹ\M�d���oj1�mAb5��#&��R�R�})���	k�rɩ��i�!�1���*
��n2P糞��͸W/LRR4�0�a)J�����j�5�r)�BC�UN��|�Z��J�Ub�(�(�ѓ+:���h����Eu��=i��T�+؞�Ӓ1[���hH�nKD&���
��P�{Q]JS�WH�jmks�!?t�.�S��(�f:��Н�*-1H������=�9&�v�����\�ƋQ��������!�A�/H���\��&
/��D1^sf���x���9��w���[���tkr��d~�d�X�d�ډ��{S�_��\�����w�\WWpL��T`��O3�v̘�%�Wv��S�L��#Ő��aN����@����*l����+2n�q��Y�U;j��Ν[K`��v�:T����]�3��*�v��\�0+Xe챃|"BIe�U	�Ȫ,_���27��z*����9�r�ى"hr���m�d��ymY�D�g��I<����v�T��Y	���.�{�%Z�TUThb���H�PT���ζ�:\<��c>�^�O ��x�c�m�n���d%��-x �WR��Ś�9ņx�0���h���ì�[3���L��iv���\��`Ks�
�)�+�lQ��m�d,=Z+�knے�UC�C����Lp���ЮB�<sx�EuV�.1Lj��Tv�:|�O�K܋�5���Z�3+Oe	�h{�Ų����h.,�t"��v���UR,���쪎W�F6��0T.�tPc�v^��U�V�;��P�������@�,l�i���8�#=sȭ���[P�5SӬ��;cD��Bf������u����B���GS�J=1I�T��Gs��~ڦ9�MM��<+�Y̜3�5�Whf�7�[V�HW�@H���d�>��R�̘Bi�n��k���A�L����e�S�π�˶�,˳�/����ӭDաTaK.�]&Vƚڽw�]�+�V:�P69v���RլGW�u��|���<�'^�ޝ�ۄ�|x]w�κ�c2r������އE��VM.�:�\�a9����I��N�z}���I�UB�uԡ�zHB�'�B�}zH
�P��C�y�:�*Y�[Ju˯�sph~҇TA�����u'I���Oo�J�W\C���^��Eu��1i]�v�*�eʧl^vV�����Q<���� E��1���1�n�e)�9=��(T��a�+���L7R8ev�7;Pz@�G6��bC҂����`�%J�nd%P�r)o<�d��\q��	(p�3�h:��*�����\֔"v&aTt�R�n�1�*�ee#��-\*�F����\3�$ג�MX�3��V:��dX��X�u���M� +��1�k��oz\B�%�����'Ӎ�� Nً�®RX={�,�}gV"{p�;��S��kf�_V>UHDu��.�k˱7��gf/ᢄ�� 6��O�:>~ͬ����.�y��Z�Aژ�W�-�#c�S&��|��a�k��"��jt�7�w�D�^7�U�l�&���z����:@��g�v4�� �6]��H��Fٌ�u��yQ���u�*�B��Я(e��`u!y����x���]��ö�:]^k�%���㫡�oR�au�K��A�B���q
÷5�
>���l�C��_2p�k��+�J�)�A�7�Ff�k��#ۭ`��1�ܹB�u!W)w]��O;��=�M�g���E4ɑ��Z7�xMI��+���ـ9S>^�+
��U<�v}�ɔ�-�Z�jw^�9i�me½����z�����b����3q�<��!�hS⣄➱ێ5Gf���t��!�+k֒�Txd{iS�s�=�%#�|M���l���͕e�57y��Q�7:��C�ױD���n}�;�wL)1��*�-TP�����ܟӖ��(��;R�U;�9��AF-��r�1\�x�P4c��`m&�҇_��#ǡ��A{S?�򼟻SH���K&�0l2��>�U¶���)�F�I�9��eз����*�tYo��s�T<�@Ω_��l��8�o���nB�kʧ+�)�"ܜ�Cz��Ù�����r��`�JY<n���ɹ+�pn�	A�NI��9�;�޺��9�c�X+Յo�1V���0�'I�\l���������Q�tk��=��j|Ү��IM���-�"�}��E���s$��ra�|��2��������!���G}7&��,��;|����yh- ��$�&�$I3I4�2 �nVX��%[�;7���́ˬ䒲���vޖH1L�Į�8����Y[%Z��Ֆ�L�����sR�c��s���A�3�o�k���t���M�:�bg%���P�R%�T%$:O.��gd�^�VMĹ�fT�������,�|��"83*��76��!���e:b�E���DLBsb��8D�'u�+b��M�OLq��Z���9�p�.c(Ք�߃l���L������1TU��h��Uլ�E`!�e!O�l��`X��b�1WL�A�B���tXљ��[�R3��Ds�s����ߌ��^�x'˧n���j�ȃV����
�Y��W(�9���3��s��Ѯ:u+Ãy7'�5i�َ{�Ҷ��(ۛv�"\F�gaX_so3]�}`v��
�u�U1��%���Jr&��WfD_��7���!	�q���r�'����3�L͎&�U�eTs�Q�
�,F8,_7Hi1�x?��C�K*�R����zE�~zz����&��/*��
���F(�#����g!�`���κ�F���� ���q��1^G����F�u�Y솚�ڽ1�0�[k�Q%I��b�bdQ���᷵b���a6�Qo�mfB'hF�=+]%�m:e��c%b��q��r�a�"�gu�����m�E���+x�/.��Z���Q�h74H��׵v��_,��+#�i�������wӾ
8���esXWwr���k7�.��VpX�@��T��>H�O
Aы�X�����ըNLB�oi�=n%Vw�I��.Z��n�1_�fH�Y4$q6�Z q0�L�GJj��ڄ>Ώۆ㴝�y��� P�pe�S���N�b�L6bเl���@u;��2�U��e���W4u2o0�ɽŀ�R�ʾK��hS;"��s�^TĢ��D1Nl��O��s/}�}��I(%^�~�.�"�ջ���k�Lh�!$���T'q2*�þ;.L@��&�7!�'��qN$�vz��q3�la���g��9�F �1�[wl\!ipw��n�/u��kl^v]���,V��8Qr.Y5�g��9�l4�y��:�>�:�S��<����opqٽD58�&�B��ҽ�E�x�0��Z)�,h?�W�9�dnC���'	b5`:�z���DZ:��d�u��t�V)ͩ�kh�C�C���B����[V�5��g��
��A`1�3��tƫ�tv��D��a�,�
�:�xpΙ�����\I�в��M���v����ּY:�/D���ކ�R�[�]װ�Vo�xV�M����C��t���h�V�)����<�G����n������a<ܦw]�רF���b@	�U��wa�;s{��E�U�b΂�'��ZKoe|rv7X�]����(E}�B�2MP��ҭ�ޕ�����Vj��=r�u�!�0+XSJeVb�G�QO-�_w���$[Ǧ7����
�U=7�r�j�=���Mq��ԽU�h ����n�Vl�5�O]S��&Q��#�r��>8�P�6�y�fҧ��ƨ�}S�@Xa�\�7-居mD�zd��j�_��j
�p�E�gtV�+n��;�͝{��`��9����1z}���I/�,uԠ8��Y/k�}�{9����~ޞ2v��a�T�(Ud�7	:L��P��D��u�d3-��̊s�����o�ʉ��~�u�ae�-6K{pe�41�0u��:q;����+2ʕ}J)] m�o<;+&�~����!�{e��L�i���2����W����Lxp#�ED<)��X;���զvU΍�x}���4J*��u�먬�u��>N�𥔕u�k{+��
ߺ��٥Jkj(!p�ц�̒�dŉhfv�	�;�uU���R�v�@6��/���v.�o¶����{s��w��5R��*MA,a��-eM�ɱ>� }����]�9�o&3��b����U)Zmu����˦��p�
T��vŵ�`m�I�g4��"��u_+̭�duiA܇</_w�|��P�I\E���'U�(:�'l�K�#.gC91a	z^�P-tc�p���k.3����@l��L�]D:חaN�Ŋ�&'���5u�G^{x!t5F����8:./&(T_H��LV�^&�}�����w�	�gcXev��YQeǡy��d,���fCY{�F��;j`^�tc/U"P�b�h@ǲ��t������{gh�]g�=^u#VZ7�>��$�m���lϦ1��u������[��]8����ͬ���G^*#��r�s���U��G�g$�e�(���E��;���X�7�.!)��9�a��]~˅��t=�9���u�M��U:]��l�����qs)ZP�:ͨ/6Ss���;�����A\�j����YM�VZщ��5C����\;ƮU����Μ�p:Z�VrUc�a�PHt��t ֕B�0��4�t�J��&�i���ل"o%	f04�pS��vl�eZN�y#����$
/(�ٕo�So�b�3̩�v�}��»���n]�tS�˂Xܸ�����X��О�n\�׶�iy`T�Fg7�r�G$s#�u�&�F:s��][�����|2�V�r}��s��YD9¶�3�{n3�Աmȶ����5L�ۡ�'U�;�tĭ��[պ��c�WϣA�Ø�hp�s2�I_�B}׶ju��S���F�KB���R|�&�hA��@u�9�D���xߜ�t/x8��=Ec2�M[H�=1�Z�\'����s���(�	�L*1Q���ɹ�99�r�$�\p����!\EM����������5M�� hU��ߺ&�N�O�%T��Y`;G*I����+�_�¶J��Z����Q��Il��k�����Z8&s�H>"J
D�ꄤ������#��Lu�=��:7�v��}6̱T˿<���o��g% ')�,�>�!3BQ�м��u��qĞ��I,�c=Q�I��5I(��O��f�l42ެq#C�۫����Ũ��E���"��m
w["��y�b�kC)^8)a��:�~۶ >�k�������&�/�h$��2ˆ�Q�}15�6MDrʑ��2���5k!�N
��Nvs.�5�	���e��H�ɸY>T�J���p}����z�W�t�����-�ׁ=z�S\��yn��7��$ʝW�[�I-�C����(R`s���KQ�@OE�6�8)��ں�n
T�#�K�wR]�sT2t���͗ʶp@�3��ն륅�E����3��
y�$ct���Z��r�G�Z�mN��,'���!SGq2u2���1��EX�e�M�D�[[Sj�wj.�P6�1%`냃��U��(����,��6�qAn��d���:Bb��p�ھ�ް�S�x�Ƭ��EZ��cz���صmvΖ�өYK6���/Y�{6�˛�������X&�d��Z��GD46�a���h�GU��ݡ�:����dglb��Ɉ���ٱB����<5�Z��z��j��-CZ�*!yo�XQM8lV��S���]q�$�*RN���٧^��� l���[�ǐ�|�sޥ�:�;u�Ǚ΄�>�}���[hkI����3Z)��WW2`Nk��{�%�����{]c��;�غ���ٍ�nV�YY���k-��a\��"[eY�U���]�lƯ���y�P�� �TFPx�dn���
ƕE�͚���9y͕�۩��Mj�^��15^@e�GNTã��g'��YSL���hXiY2M+ii�P�}�q0FMN�e�2#ku��yt]Z76�F&W��7��Qz{�����,.�hk�.�il3yG�e��骋��'H#w���C�_k�2.���NN�b� <�L[�q��5ۺP��8�≷]�p�(4�C��� �w&N�R:a�*��8V�������铥�B-�'_S�F4>�U�ݹ��	�:�+UЭk-6�*'����W(Z�̾}�� �h]����J]ΰ�:n���<'����T$(D3�vt�ꮑR�dЄ<ZNRk���3~�c�]/I���:WJ�rߕ�N�|�2%������v�mD.�.�u����l9n���CUL�w[��]Gg[���ˡ��
Yz��[bv�K��S<�+Fvj��ά�7ݳjGI�͔.�
���א���Si`S�-�(s[@Kz͊}E�g-�+.\U��X7hs۠weh ;+�M�(��Z�A|ױ�����Z��W���A�w��XE�F͊wH"r��9GP�x+�X���2���Ν3��o7V���ӐYY�n�os�ϕ0���G]:�LWK�Ʈ֌k4�xr�	��W!�r�mtɑ���͍\\ޭ�b��@�(�nj��=�awK5��kGt��ۿ�a�t�W�Ρ�\�V�sFe ��6xi�R��o��.��N��7F��I��c�t��aZ��B���F=�QCGc�{�fd��Wb�پ� ���IYpR��4�<G]8��1�};B�\/'Q P��,��3��YH�ۺ���"���%�U����X��#��u̺�o��]�7�s��7z-�m��H�Z�u�W���a-gz8 �-��Q��lQ�QUQX�i�+VZ��JتT���հEL��Il*3�U��9J5�,b�Q�QAQ��[b�"Ee�t�-]U
+�� �Z�U��4�Uj
������&�V,Db+�UELh�QM5E"��PD�Z)TUX��V�TU��"�X����QH�%q�U(���U�"�)n�F*	QQT����QAMZ(²�"����(�C�����(��:eU��B�Ub��b�P��*+*,Y�c����cUQdTPQ�-JU"��",\���EjUqV%��DPQ"�R,���X�ESZ̑B�j���TX,Fj�V[3,T���D`�EUX�(�,X�YJԭ�B��DTb��h�EQ`"V��1���b�UQ��`���TAT�,0e�(��{�=����'k�'�2K�2��{0+�b�n�]V��7n��ųoh�@��«t����M�k�Ja��xY[:u4��ԇ`�҇�S/fP�G,�����WfD'�j7��]����n�/z8�ޯ>���������J�?fa�.x.ʨ�j�B�j�#/��5��YB՜�ьw9���fe�K&��P��C1P@#J�,�����ae�T.5�{P������jqE�Y\���RkUi�yݖ��IW�B*�9�b��$QS|N9�>�ۅ��-_5��W�-�8�|c0�{�|'C�BF'T謀|���P�s!ًuP��8�=z^n��v^�n�ͩ	�=�TI�s)�`/o@���C��K��&��j��!t�pרA)������PB@�Űx^l�.�Q�Q��w����D;��2�U�6���΅�W�l���璢�lc4�I�qs�b�#l�>��E
�=eɂ�s176h�7�;!7�QVqR�J���<��3�}xɪ.�w!l\�1>����c��O�d���T'%�TüH���f�%|��GCY�.������f�"=hkM|�B^�VxQ%U�u�O�U�831��3hVM��e��y�qR�*ĉ���t�I�%�ws�Nh���A)��:`��KOo�~����<�T9^mұ0���ߗ�yh����M�Z�q>���.�s�c��]�;!�SY�19\o��+�r9�0c��{���}��8f�$NƂ�e�F�˸`Y�����l;��\咍�Qv'^���X�;^ڜ+$����Y�8��/�q�Lp�2�2R���OR�N�cA���C��[��	K����F����&#'e�B��;��C�����9�1~kh�T<9�&�^o�=v�X9��=ѕ!��PB�q�������>],<�,�
��b<8gL�`�
]�.1^�U��� �K�ӂD���A�UG+��Tcn5�`�B�A��A���d���+ۮt��X��Ԩ���5Q���dQ�WmW��[P�U=,�]4��Μ��u�ɂ�Ȋ�[lh(�C}e*:܀��PҮ�����L5�������W�S��.$�nspuy��S����F�Zn%��3�k�;�������/�U���;o-�=ޱ4�i�����hx���L{y�����]qԠ�ITd�Q1'�7pޙz+*?(;�H��(��R����1�P���f�'I���ت߈�t����$E+9�,��|d׺'��(���*i'���ܨ7=z�W��t�6�}�*�OE�3��oSN�a]X�gn�дks�&o��>6����1j��P��}� �w��Y7��Ō��i���μ'Kl����b��n�.{��w|�A��2�y�m�"��+n��l��j�F�ŶQ<*d)^�F���T�Ju�3�j�����Ƥgsޮp���k��6�6kC�y�e��DTKQ��/j%��9�.C��Ɉ]I��SYI��H����J��Ou�K��4���E\�/�^#��7�>C�ﮌ���hr�}�?=N;!�8j~LHc��чh�I-LXʦ|4:+p�U���㢖*���^�X�k��nC�k��\�q��U�^��3m�Ķ�%�8���8e�F\DΆ+�5�ㅧd�&�Iq]9f��P��`dmSr�7��C�yp)�y��R�h�19�Hv�)f���gf�}�	����
�)�-�������gZ���V=3���
�}�`�IVԷ��ء��3�WD�Mr�Hh�]{Sh�}���\F�D�B6�ed^T���e^�������ٹQ���uŵ#Vx:Ѽ`��x�W��L�o"`�F�UW��z_I����}֖��}�=Y�C��̭9'DT4��dk�x�����uw��U`����`��Ҙ�+���&W�D^�X&콞��0�^��-�k�^�'}UÂ9��R��k�/�����VAai�	w��0ޕ�	��"���є�̒վ,��X4�|��;��:U���9W�y�\���%f$��Μ1M�鵈����g���cjn�x��о:$vy:���f����bYJ��}(�@+Uׂ*B0Fu�HL�k��J%�t�ن��C��b�{Ӑ��Bu0��Rcn5PV����Z`����g^�1e�Mz��q7�<�e�2P�b�S�o�@ю��I���cbjR�s�3Wo[ɹ����y�%�St�d	�7��n���)�VU�磗GȞۘ��}-nդ�n`E���J]P�@�¨�#�kZ/�f/,4в6�����Wr[���j�qqיE�m1'rf�
)J'�Úb#4�[Y%Q���Py�K,>��9
�k�Z��6x�=���1�b��73�u� 's$��&�jW>�~�T��u�E@�ޤ8̓��<��e����5�c:��,�:J���,q�I0���}S�1i�5/�fcȭI����ULfb08�8&j2�u�(�JD��S˰�9$�E�#\�B{�$f���b�ܿK�v�꼺++�4Aܔ �e:c�E�}dE�˫`[�Ջ�ˉ�KH8�+��ܬ�Q��\��Dn�{�F��tm��l����$#��j� �8z��\4&zgL
���-u��Ӭ��QT��VnS���|H��4�]˱�LV@�&���#*Wu]Ԝh8�V��_7�\b���,ٻcZ]/y#�Ws�o.���v�Bq}�8Z�G_AT�s�Psr�d\�Q�(=���(2TۺQs���N�S4��4G���xq�S��W2#�#6ǘ/��2��|��uO0��Q�(l�`�Z
��^�����U�c͚��f��5]�2�[������;���v�}UKl.z�+Z�˅x�ɬ�����<��|��>�n��Ƣ�t�{(��7n�;�'�z9J�o*.�V�x��O�L�kSڒ��r��1]�e��[�k	�B�+<�g-O+<�m�O�ɉ2�-;+cqRsk��Nc�N�j=Q�*�W��ˌ]1�r�S�z@�{��L���ԁ]��f��4�µ+��U�u�=b�+�^��/"&8����ӻ�i�
�8���o4�d�W5	˕p5*��S������^���p�}|_�&���E?U>���)���8��J��eOr�@�+���J���1[B�ڤ�5�P&�
>��.�]D+6�6����Yu��n���;���黢���K��n���l��yt��R��zX��9	�p�AU��,�IԤ��[���]�.��G+�vٮUS���X`�u�BmwN�]bG��v���U����{���UM��;a;1>���V6�幅�����UR�yו�z�*�N'�dlJ����ҥ;�7u6&�iu9��S(�D?u�B�2���Nw1tV�X^��+������Nl�d��b�ƽ\.���u��#T�۟ �PZy�^ߩsw�Ng����=��x�C���ޖ�|*�>N�f�����ױ��o-KH�ZW�^�(�Ro9��E�A�)�G[B�px�NsÞ�W��,2oWXSصپ�-9k(cK\%�m8��^��Z��51*��*�pj��~�r�󺈽c3�r����Z�6Qf�[oF��Ԅ�����Bw�x��f�\�c�2�-O!G:]�:�$��h�o�.�Y9�'�et�+Db��]�o���F�gU��=���:� +I���'���%���Ն��s]ѪܽRɴfk�E|��>���>[�+���F��\Ȱu�#�����F1��C�[J��}.Ny;�Z �@�/���v��U�4���y�`�ˉhdL�J�[�,WV��~������rX��`��Vz��;��wd�{�s�bb�7�5Ga���z���+�B�8�l��*S�U�Q|�w5���N����U�N�jި�:�Zڂݻ��J��	CKT���ӓ�6�#�\=�ʻ��w������{�F�|/^+V9Q�!J���l&��]T��T$s��x#k� >w��+5ǾI�7��=�I*��l�ꍗ ��{�+�׫����yg������1ٮ�s�r|k-U>���1�7�L����ʋqkL+G�D������¯�c'؞m�s�ܾ(FywQr��$7o�BΗ��j��}K�"b)1��_kC��mgː�a���aM�zݧ�A�JS�7M#ae�*_W��Ws1-�+��T[O�頝k'l�������wM5��p:�k0�X��o�gJ��{x�gE���ݷS��W�c%���LR��1��2��5h
�!�<]rEq+:d����@�7K��N��Uy������Ng*쭿J�F¯J������v,�=�����y.�ْ�%�me��檈��ǘN�vLV!�Җrw�"��ʹ#w�xS��Ѻ�į;�l�ќUc�5�G���J�\JC���2���D����a��l�9��+2�E��ge1Q�Х���vh���j��|��./��v/w���<E\��{U�Q���jC���NJ2�/dv�O�U{��޽�ZÊ�uU�ؒ���Wr�4�Mqٽ%�MQk��̾���w�����:sj�k|gd�v蝝K�9ͳԼ��i;�qk��w-W��X�Si��oB괱N���	B����WEd+V��Wg\A��Qi*��N�j��ي�k*Q�Ӛ7�:�@�M�k���$���ˈ�k��C��Z����-�����%��F��+�&�{�Ҩ������
��@�M���ک�s^��X��o�} �r2y&g��K��/�'.T\j/O5 ����l�{�Xļ �������g�f�	�*{�i!¼媈��<����ĻV�R���>��e��.P�:��(�z�@�I
���6@G�'em�s�= ph�6��뼡r���o�2<�����,�}1�vDI�5�P�7#�k��Zu鍌��V��AK�F6�wG��yQ.n�޲Z1t��fη�ܤ�{���(Jb;:�&�u���1��Peux=�5o ӑb��V-y6��g\U�8�u�WDk�)�9�t��1͞�n'���Y��J{����� �]p�n���f-�3�鍉S�7�r��%�W��D�t�7A!'�~��v_��@;v��=&�vKu	����b-���9|��پ�QgF� �U�~.:�׾9��+2�<;�E����w7SQ�;:C�z)�X�NrÔ��.q�oe?cu��'՗�}�'��asY��-چ�W��Ǜ5���w��L��]����z����{�lN�>�<�5�kAjw�|�Y���K*��6C�}�O>Ƨwӎ��'o��:��\���>]��0��Ld�*�QȽiG�v�Ve�����N����;<%rVy�r�^��;��,��;;ܱ��x�V�^ޏ	�Ӛ�j/C�|M�{�d6����z໼��'�!$&fT7���T%d���t��-���]����θ�b����ލ�|a4m�J�r�0�I�}ۢ�D�\�m�����.�g.����=3���)��n�<S�����W���x�/L�%�o�=V9���Ecc_�-3���:�s!^��&v��*���C�S�!W�\�1ZC7�Z��tWj���'��{5(�k��d�W)�*1r��U:��'�i�Mhn�.n�,����K��r>��Q9��{�1i��T�-rl�ѝ�v��B�Y**N�<�e@]{q\��g:p�lߋ��N�SP�8���G0
ŭ�'P�̥P�enuc1;��W>ؕ:���J��Y��ut׼%Υ��*
#;��2��R�[��+���^LFĤ��ܩ1i؛}i��8x�z&yiCǯ��K�!kS�*�K��F�3���q��H��mw4�
�)��T-:���������:��Z�A��O�'�"f��G��)�!�P��Y�ޗ��~��{i׿~]���]!$ I?�$�	'�$�	'���$����$��IO�BH@�����$��IO�!$ I?脐�$�rB����$�ID���$�!$ I?�	!I��$�؄��$��$�	'�BH@��	!I�	!I��
�2���dS����������>�����>��]��f��l�`	245��-����&��B���VmL �I@� (昙2h�`��` ���S�JT�       9�&L�0�&&��!�0#� %R��i�&	���i��Lj@��#��0�bh�2h�%A2ħ��`S�6�dڞ�iN;�਀��A��* �?h4�Q�D��� �YO����OԔ�8Ad�n aH!b
����b�||/�O��n	�����@�ؔ���ᰣ�|��u%��PQB/��SA����le�q+��a��!]��O� ��p���̸5p�,L�S�*i�s�VD�",���A&�M���[2sᒡŅ�]�)���
���q�o+�b�5J�Ɇ&@q��H�*ڌ�k�3B��2n��(U^
�9�1r��%�7qNc.qK5r�*��5s19p<�!��e@2"e\#v�5��@�s)�*]	��F��/p�E��r���P�2*�j�2��V�H����
��0!�(ڢ<(-�Ĭ�bfr���(�TUR�m�(w�9�xU�:��7WN��K��LU]�Na5���`J&M�fT��S79'r/	
Th�V��P�V�&��ۛ�xi╆��E|�;��������~�t8V����r���R���m6/+K�n���~<�v����B����89WY�����wy�`p5���$�i���֛m���m��4��{ul��L��wv�i�;צ2�-���(�4*���oC���t�{j�nΩf��ʭY2��zn�oQZ/~�ȫ��=��;����(k$D̢^��2kgn�mf3vo�8�ꡝ#jDY�s�OwsuI���F(M\=�w^ڄ��u����YbVa�D�fu;	ƤYy�f^�*�≓ZNꣳ���m�#w	Pޚ ��NM��j�ġ뇅���
�+4��nq�Ķ�F ��˵W�J �qgf$5ε�F�W4��QKv�Ė��;a�X���[�0�l���e�e(�Ɠ����
��s�մ��#Lk��ւ�:d�����"�w�PP�\Na�T�0+&�}cZ�����W1�Y?��X�u��5*4i���"�V��I�ܪjv�q��(N���hex�����b���k%Ѩ�.��i���#%�ȷ��W;���:�LZ�56�bP+����� ��l'S���F�T T�b]�St	J*���!�b)��͗W�5C���b��Q�\0�ffI$mL�S!�R�����B��^`�$��]dT�3z"�D�!��M���ʚ@��-e�a�s�T'S�Su�M� R����G �1N�s	͵�yb�0�;%�L>:MP>��*�jl�B��P�*�\]���S2�B&�X�I�N94l�e�@S�I�.hd����7e*
'���َ��	"��C����GM(�;�_����M��Ùi2�����hb[td���8��xG@��ª�(�"(�UTU"�1`,:��Z����ͽ��E&o���:)�����c����n���F��O8UB��5���(�t���F��F>q-a�	�c�9%җ��Z�OH�#�G;+��sm�y�ž4*6��@�i/���`�h�9��;�i�C�p�q:V�GKe��[#Y6�^�5}xYDEVWGdOob:��K̮��IJ�-�U��u&
��@�������Mv���z&71۞��t�P�T�A-d�c�=\GZ�6��3Y���ٱ���Q?~��=�����*Q~�+�-�e���F�^�Kl]6�s.Nc=��a���`�ӝ����Yg3&�,k����!S�t�P�N�8��>
}��,F)"�(���U`�*��s~�6^�y_z�~L9�Y��{:q�.�.����k��z���>�j��t�lT7P�����fw3�~�:���1�X�[y�G�o8ѽ�%�5�mz��=����f ��G����O5�ŧ��w���Fo�^��E�Nb5�h=����e�½�����>�Ff�aN��׹�t�K��g����n���Oi���kj'����Vc^�=����Q�G���1yS���8���v�C�9&�^���+��>s||���h�����7��8eU��U�:}58�k�}Y�ae�fJ%'E��aN�U&��;�T�IQ>��]��,��z�z���L��Y�+lʩ7���Z]����(�`�Y ��{~���uo.�2c��}���(��w`3ôFur=�4:�������c-҃��йҎz�r�6-E�蝌����T�_{�[{��t��lv��v��l<y$�Z��M��vu�6����64��nM���d�f�K��5[\kл_Q�t�!�[�%`�<�p�rB�;����g� �e�XI�.�Ep�  m�b�+I8fٜ��N��㓱c�ҹ�1&s%g)!N$u�u:�)�c:�b�˭��X��/����y���%zX�"��b�+oLc�sC)�ek���;����{}��.�OZX�d*c,:��^Ҷܻ�X�_[�+�9�WJ�)���@��Y9[��SS�as4��3:J���;�2/\[�]���1�-j�ǳ�ox����=�o��}�F'������OQ�̗\E����W��e*�{��ۣ�WW.��Y	\uFhOus3Ѡ�s������6����li��u���I��88��1�d���b�[y W���p�;z�b�Tn�0��C�m�v�t���J�Lgi�\���}{k0)�J�Ԋ1ÝOf��ƛ���ww���������X�="�\����!����� k�mMQR���>�C���$�|J���.�*��ݺ���J4DH���7n��:K���8��B*��M��[OZX�Z�ce��f��4�<��[34�r��#���b���t�Gr�3x��A���ĕ� �Бw���v8ˌ�f� �b���ʭ8�#d��qr������0lF.P��$��G�9�]���]�`��������	�p�u�r9��/z���g�[��g�	$�B}�%vjJ��cA�Q���@�7�0���pC�:��*^��Pl@�DY0����WGoV�N��g���U����h�D�,�2��.�q���iv�O&�?/�x14at��E����z��1�[ư�P`�1��K˿DD@����y*/���Y��#4�!3#,��#�ꭚ�}��rDl��`��P1����KtF�&1�X�����բ���S�=�=
���*mD��ڊ��/--�xqL��T��)3�[oZ6��'q�d���sUթR\��ܼ�M���?ώ��w�@���4j�r�{رⴢ��X�'��	r�4kk׹��1G<`����� �P��4��K���#EC��M	����DF�$������ O��ya����bт��+ɍ�:̬ۮ��D@1[��3Ҁ����P��(�6"l�g)��P�Ow����|~��f��8��� �@Gkތ:�4��<�"� �վ�s�g&��/�b�qbu�#L�Dɷ�Úk �{����G�|/�+�/jB$?����Q�./�T"��z;�2L�ʯ}�DC�#O��#���4#h����a�� <!c+���go��}���[0xI�Ɠx���y���0h"���݊��=�~������!b"h�&J�J(ǔhU�I��k�qS#��f��/�5���UWC2�/*�Ҩ��y���y�m�M�:�e�l���t��@q�f�#gh�暼�/��L����m|g�$$�m3Tw����ү�>P�M`��Y��/X���k��]��"
�#��4G8J��h��Ì�<���T�)��l��Wy^��ߤ��(�=g�bD^��XO���i=�����w�y舁\5Ja����$��^i�TbDǱ��`B�u�߃��>zfG����dM�Ѫ<G���N�s���/�����>4$R��O(�C���c�/��"�¹̺Vn��<w�;��=��}��c��M� �Z@6H��gZϨ��x�� �b3���Q�1�p����z�E��2vW�]�o�BJ�`{�����i�e�g��Q�^�n�[P2���Dt�:�1���`�X���<����p+�/��}�׶�.�t���9����X��"&����iaw�h��A�8��3m�6�h�hm�k"��i��ȫ��Th�r��p�p>G���瑠D�Z�-������I�`a��E���_)�Ʒ�u9��$�����0����j����\⫹^ɛ/g,h�(�4F���N,0�&d#듍������A��R����c�IP/��>�{z�/`P�,k傦���I"A�39F#�bDv��}3Z* ��(��:�`���C(�%���	���ŝ�4��[/�:��|Ֆo_hLf�0� ��f�P��:.�r��a�U�nr(q��w
VV�0�=,�+�:��!]Tt�-�}�-ŇV���[�9`���䉷@�d˅h�Zo\aQ��a����wcg!��
nmvU3gi'�Km������I f$�X.�$N�n�=z�I����   DUDXީPP
 � ����Ӄ��s��G��38w��ˍ��N��{�8�L^nc�J�� �a�ΥUe�6;;u8ԇp���}1���Y�ڃ7�T�Ԯ,�)*��ŉ1�N@��&��K�[���'�D��Y��z������S"Vn'
yv���)C��J.f�F&X�%��d;�y���k�1�Wϗ:�R=ۍ�G-�|�;�,x�����.����L6�͇懮pa�#�Xcu��]	�<���<ӄF�Fa��{��=[�-�+tC��J���lT��CK@n�Å�ܝ�[Om�-v]jvW�35$�hywgV�Vu�r���ێ�8EEUUTE��DU��PX+� ��n��t_�8��d}3x�lZ逳A�]��gqf��2��k� �S�!
��V�wj��;huk�mڲi�ƞ�
ٺ-_W#�y�[���k�7"�j����P�(�嗚c�+�x�y��^S&�L���,��8ɖN��RI2�����(@֒�n�\�:��Mv�d�Y(�u!M�C���q��
ά���,ɆMcv!vaԳ�&�
�����p:�PRC�u��C�Y&��:�Nr�
a4��"��fPS(l��St��'i��|�o��3���&P�6�e������� i��087��j���������{)vt��W�s��4B�
u�v����f�]юtu����$�}���@zW�T��Ҫ*��TH K4|�@ýh�( �󄗇�S
��*S�E���M��m�mt�Z��H� M&P�;I�CA�o�I/�F�P=�Ȃ ��(�i0���=��K}s�1��=A�J�����T���cU��8G��ac<�������Ƌ��� �L��=ڵ���`%�8��?�����dJ-N�?�]؜(��e��H|5V��S���X8fJ8�* 8�@�֡��$;p� ��
���B���B�f+�)}`���JuV��~��ݹ�&K��Ju��2����K��5�xU����L �p��s��cʴ��[���at�+��B��x�������6���T��	Ʈ�P6�F��r�>�����C������hi�#E@��4&k��M/�/���5бZz�J8� �^/�.}GHpy'�r�Ht�~{t^e��=�A��� v'(���q��Ϥq�,Ԟԇe�@4Q@j�s ?S��Py�}@�#Ħ��dbY(#��E��(���m��ǠZXP���d�t @�d�I�B��Zd0�p䉌SIQ=�23��}��bR��qk��}j�� �����ۨ�8
 7}�R�0�ͯ=�p��~Z'�� ����֛֢>���wQ�=�k��C�s�9� ��ԯ�~�)��� 2�d���'�P�7�B`T�y�����`b:.�X5�=-��XT�s�B�0�Q��N\��t����G黷�aB��im.� x��qM��$���}��Þ!� �'�T��n6��ł�
zX$�� ق�W�
�����yl0��D��C��x]��Ǎ�!RlI�Z��W�<�ROz	�� �d9�����H�
J�	�