BZh91AY&SY1���f_�py����߰����  a~�               �� � �
  �h  �(  ��I) *
*�� 	 }>�� 
��\���^�w��z�x����!����o=�����g��p��7H�b��Ѫ9ǃ�����f�j���1�zR缪��On��s:j�Fڮ�Po ��� g=&�{Ɨ���WoNm���W��<]��%z���Y���N�����uS���ӣ���������v�ѽ:g�G����=vw5]�q�v;������f�o<DQK�{��c�����ݝ��uܵ�����=��׸�x���v9 ��k�ѥ�j�z��;�˶��m�]Nv;��Uy���g�u=�]zn�T*��E	UDs��]��lٳ�����州�[2�w��p�+��W��KM��VmV�v뷼�6�4;���q�[�C��۫{��������J��@�/ei���vu]��ox�ʑ5����5�rvkٸP9��u���=�۽ݶz���;���y��ͻ�zφ�   4              � 4  ��1�)R�e0� ��a2�� 4��$�Q� ��  �i�M0y��4h i�� i�400I���*U# #10 M4�`@
�� L��4��h�z��6��L�
zj�@5*�#M0	��i�� ` �<�NǚcT��Vs{3s�9;�\���6i����NO�36�ٍ��y6��f���?�qÇ����lm�7���g.|�;;�?�����&�]�Wc����u<�H����֒�w��6l�9!��P��Up���6ͳf�[7�C:�9eUUU^<�����v���};|�����_?���v��}.���;\quq��u}ˏ�c4�Ց,��j���2�$��Ζv\+$P�]P0x����0��J%&I��.�C�ZiC5&h͗H��b2ҫd���:�C,�(��,�2e>�d����5�f���&=�>[QE�#�+�-���{�g�ݷ��_m�a�s=m0����ޣ�)�C(��2Dh���	�C��,��P�{��
4!+(�҇Q3��U�u�QҘ�	�1}\�U�1ꡛ���B2��
�X�Tq�J��d-Q���i�MTD*��$}L��D1��L�vb��z�RH�ȓi3Gn"=�1賫�;I�t}؆H�%�Ό�] u��;Le6���1ܨ����8Lcv�����̅я���ڎO2P�)��Qm$�u�#��`Ǌ35��M|Ti-cjN�C�c1ʆtr�r	�P�&�r����1�Ap��}P����2p�`�TX�5aCQ��R&u�dF5QE>(ђ���3[QF��|VX�Ҏ��u"F@��4!0e��>�Ԑ>`�ĝ)$c��;�h�1���|o��	�}V0x�̅CT�c��]�QP��H|'�T$'؎��1!���B�8`W(d"(gFS���
/z��X�X��1�����,��c+��c�e3F"��5�h�臁�T�h�e�_Z]��d�&B��I$\c:�It1�ǣ,�4���2��x�RD-�L�ص�]l*-3�dQ�!�iP�P�i�`�!8,�p�GZ�lgJb:.��:ʺ��c�`�;H�2a�P�Ш\|�	��J�+'�P�KD=L�ؓi)�H�0�L'k�z�fmB��.���1�cK��"�"�)���N�t�t�Όw�і7��c0r�f�2q��$���@���n�2Dd�qDP���nax���3ǏV2<t�FQ�<"�� Fmi%i�dt������d&2�Ů њU8T2�3HdЩ\��:�L��I�P���1�aq�Bc݄��F����[��q�і�4��©I�N�"�2�5�naID��U
�:>�&u�l&1�#�çz�e�l��Ι.Ѝޑћ��3N���T2��)�넇�Ζ�C�K��u,�d)�0����Pk:Y":�(D�)�βA=�p�兓*``��@�n!A��j�a'G�&tc����'� i�њ_\+d�D0�]�'ڄ����=�L���4{�L҇m$\�#�%�w�(o���I�\&t����i�Ib".0f�&�{�(e- �o�������3Y��|�	�3L�
�(�����aH�1�a3Fw�	��p��YO��������!3�,$f'	�#	"��1���.��C����Y	����p����4��cv�z��;zD�d3��fkFP�yd@�ŃZE�������Z2#����gG�GG�Bͅd��\L谲�!�c4c�"GA�q���2�|O���c&3�٧I�EU���#8�(�ţ䌁��
��\JO{	�aYP�c]���BeW��d2K:2�Ώ�amoi,:3N�¡�2�z�a�1Y2�I,�d2F]�T3L�F��p���Z��ȋ).�&�.�����Tl($��\�0`�q���0�F���p��mL)`�	�Z1ӄ�"��ӣ��BI�t��n,�Lc����X�OD����=�L�B�1�BcHcYA��L��z�c(»��dW�����9�I.1�W��1�.N��1�0C)� cD&1��F1³��G�y
�Ӆ���dH���!���ǴD��F2&EdE�C��f!�U*�Z�L�YV� c�Q\+:0e��cjΕPD�J#0}IP�H`�'J��3M5�Cc+U��Y��c-�h��C,��Tq�q�#���H�i&tg\�c4f�Q��p�
 |mGH$d�P�te��є3��R1���ڊ(�ӭ$�`�KC�.2�>:P����](b�1�w�Dc�ьT�@�N&3Mx��@�b,�*�:T3Fk�I�bx���`�Gg�F2G:��'������Le��n�tc,cި�$s�8�yMD��t��1�ڈ4dh��E��G8��Qd�2_T2�35����i��:"M��3���f���ǵh���Y2�#\C6�.,LgJ{�C d6��(��΃:�C0g^�c(o�F`�te��!�P�&"��"I:�q�S%wp�̱�DҴ���c����7�$2a1�DH�n#�����v�>�GS�h�ih���㸂�����®b&R��}��V2Fcj,Ҍ|LэҌ4���v�R!�\A|q4���#�m@�hIq�����G֨�与@�K�ƅ�5j)�a�Er2 %H��#(e<���Xλ��Dl(��)�*Ռ�،b�Ln#-��ы:S�d����7*,�j8��A��U5H���mCc] ���9Lю]��C�fJi2|]�2�K�c�{*0C:4��6����G��6�	w
�oWF4.>&ZR2Ii&P�t��@�c�ަhǛ�:i�4�R�
��j�=X2Fh�"ѝ�Q���Q�>2E<���%�v��.S�H�6���2Mx��Ԩ�1Rd����P�Ճ�����=�:�C0x�c�(�a#x2���BgF;qa�GOE�4{؆!�3�؆2��'�&Q#$q�H`���I�2�I�fL���e�CF>,4f��GF@����+�g�&�4�`_��h&�>Rd�}��_�v�g���_�������E�n��@�Q:Gd�m����[��/��:�))9���I�K~�ț�>�����ܭ5���s�)=d��_-�90{{���1��������2����Ν��3(흹��D}RN���K�h���U�_�ӿ�:/z^��oG�'3d�ڞ,$�G-�e��{�����P���^����-^E�K������yv�J}�Y����:��]�rv�2�b/srSm��\v�Vf�D��m̏�q��3�ȷ�ɛc�Yl����dc��U*���s���L��.�$����yl��G���󸲟��=���r���?�4oc�t?~ٳ��~�<]�[�{�Q�O\�y_E�GL�麱��fd�m���~��5�� ���g�����`�o�7�-�a�Ƿoi7��	�͛�^�&��������˙�s-8�;���u��&�njk����c-垜
b�l��o�_x(��1H��ˆS�m՗;�_���{�S2ಮ�����:�2=^���&'>Y~Y'�5\����w~c$o=�X�P�*�+�z���� �S���U�m�OG�B�gJۢ6Zc��e�b�dr�*����=��n��=���i�kg�o��^��B����{�Ε�G��,X�ոgq܃�\-��E�_wy��,��.�7\��[��v�m�Ց�Z������C}k����|>�<�����Wp~=����&{k��p[;s,��}�d����s?6u9��V1w�C͝j�[��3\j\�����4#Y�	��������ŭ�spǏM˛s:m�����ݹos�M��p:8�R��e�"k깘��߱�:e�y]����Uv����#�/��>�龥��؜�&�]Y{&)��}���ߙ�@ƙ���8Ι�����������v9y�l+����	�͛���3��|��i��]z�\�}s	:�wn'1�_�y���ױëM�O�����w�4��H��_�����E��J�6MY���LW����uv�v7�[���WE��-���Kgl���:/�����Y-^<�Ƒ��]�s��ޞYq~��}�I"	�1O���C����s�3�5�{Z̾ج�ӱa�M;Y��2�����Z���KT��L�)�bn��S	��V?��1nz��B�<�?[׹������ޕ*ڐ���W�ل�^��A��Ya��������Wje�����O�E{\�h|��.�*�ڏY��&�A��I{�2F�oj�5�S1�ΫjnXN;(5o���{�������>2XɆ��a�n+$�MO�����q����Zh���U����w�LPLX\~-7���;5e�w7��׹6�gs1�jǳ2V3Nmˎ��pݥ�js2��՛�d�w�aI����ϳ��,z���������M��i�s���UίY��䊛4���fw[_}÷�'�P$���M}��́�<;����N�a�W��T�ܗ���&�v���Pr!�j����쌛�N�&a6��3r��==.Gڽ���@���㿗���'���\��
�fw���ks
�v~��l��VO�����R�`Q�~k���fP[Q��i���ن̿1t���T5�ً�h��|����v�?vb}�m�|ÔC���qC._d��l��_��S6w���}<�}�{����%�N��L#�?��=�=�̦��M���پ찝�����'33�o�,�Z�=�=��\a���Eq�����{e�xg�ٜ�d-�M�ƾ~7鞟Ͽ���P�$�צ6���rm��8����:�)oZ��ɓ3'n����6=��3��f��hg_kR-�*��e�1]��zn*&��IY:�p�K��ɚ�f�02�&����to�y��ޘo���w;N����[1D����V��C����P�ٖ>�5�D�E��)%��e��;�[��Q�7��\&�z���fCI�������{�U�{$3ӽ]Y��t�2l���wƍAu乊cV�E�)S�ڞ,t}��%�l���~�ʧ�_�h=�7���f�3�vI����%��u�[�z/{p�^�n�q��LQ�z�x-jF��w2Y�϶ż|{}���[6��`7�o���Z�u?�yO�{_�ߵ��Q�ކ��5���{����z�r�^Ǚ�s(�{nco�Yuݙ��v;�]�f�&N�٭�h?����kY�sz���d�r��\�by����Yۆ�2�{�gz����Z��i��<���oX�e�[׺�����{��)��4�����ŗ�=��s+rf�fn�ϰ�����Z��窶+��]�2�˯&�����]�U��s0�2�����[wqٜt�e���9;�;s�o�a���:����$FY�,3f����J}oۗ&d�t�W�fN�i���墹�����O�L�N�Oik)7��z�й����Fw�3.��m]���(�=��N�@r"R.��y>;ߟ��~��ǰ�[���7Ϳᝃ߾�}�RtO�I#��mݿ�\���9{�UF�UE��)�S������e�����Z�&z�f��.����!�c��[���u���-��u��m��W�����E�WO�ɞ�x�7�ϛzӹJ���5��g��uoA��{;�c|;\���j6�����d<��e��>M���;�
6(�	�$��P�]�N^����{G�K�
f7.l�6�w�w-J�,U_zU;�����̓0G��w?{���w&f7�o����K�Fǫ6�W�{�$�<Ηw#�ܲ��V����u�6�ѭ6L�J�Y��،�?�{����l���/�M'?T��u��-��i�'
~���7˾���=�S��N�]�Ƴܯ����6Z3�.�=�k���z*�?o�����qϴ1'��ݝ�:z��'��;���w7�����8O����lEP�2�L�i��!�f��{�)���v����}'g^@��׸��e����S�f幐��(�<nw}��{���+��;5ڳ	��e}�{��g��=;����lG�����,{�oI�t�ʣ���x��G�k� ƿ<=�h{���/w�/ؾ�] ������S�;���@�
�˻���o��������)�ҧ/�?�~���[۾8鞗_W<ݻ�v?���W7��L��{�����۱bz��7�֜���,jXq�fd�eoVܰH٬
��l.���-�p&q�� �1��f7�ғ)lM��׫78���]-���X
<h9�A,ծ%�n�]r�2�-��W�/�Ե�d�s7S���}�U�����e��^&������ٺn�%���_����;�Q�I\��A7d�R���ܒ766�̒.�������X�X�.�=��Nw�{$�G�A�T�i�o��׽� �V�E���C�p�s��Y�g���gq�꓃���j�tn�]l�;*�*m���s���`������RϏ�D>'y{ ݣM�F�����wB���Z�<>7~ͩ��o{B)).�Џ<M���ˢׅ��5������{�V�ݭ��Ѽ�P�?8Y�9^�-@۲���@�>|���~Z�Q�]7\[\5�a�5b�^��=�.�"E�M��s1��Q0�R�Q�e�Z�m�(/bay�cu���.��]����m�sv�mҒ�gs�f�Yn���C�6�n�7-�1�<_b�Z[�BK]�s34�f��f��-ΖRf��-6��B~�m�ٵ���0��PjZ�u�M���ͮ¼!�MGV@�QSJGc�6���QH�R�
�g鹇ŵ*nu#3Yf�Ղk"��t>d2kH�9X�6�U�([�y��m�	!$Q9.嫹i��hrWcQCG���k���J����I⮷ �m�՚�5��"�޿;޾�:�D��R3+╳:a��h�K(Jv�a?G�]��?5�S5��8�Zs�TŇ���pȡڳֲ�'�ZƁ����/ۼ�N��{'/^�4��`FkK�^B�jM5��Y��3���]�[�cE�[L��:l�==}ޭ�/��qF{�=#7�ˉ�v��:�ɐ��u��{X�xXV`�枽�3,��,��Zx�H�Z�����4����	�����!�,V�0r�u��-,Q���s.���D���l3�{��ʱ�[j��",�;�V�Y�T�h�J�w�܌$D��EcM��c�v���*�G~�k�1�u���+{��삶��B�k��,"�QqWP�g0����Y�0��"��T��Uj���K�J�Ek����A�-y��0�R)�"2,�"{�,~3��������,�譪�SX���.��TY�D��8��_��g�)ʯg���G�q��0�g�ݽ{S�p�Kott���w������g�Y-�pH�9�%Ç?w����c��^���c�Snm��m��m���oZm�ݶ��۶�m��i��o��7m�m�m���m��m��m���{��z�n�p�m�cm��ַ9�\9ÜK�8s�@p�8��\�8 K�]m�p�n�m��9m�����6�m�p�m����۶6�m���m�nm���6ۧ-�m��n�n[ww������6��m�m�n��G9Ü��[o�m�m�m��ۦ�t�o��nm����x�6�}m�m�m���m��m������m�m��ۦ�o�˻���m�ݶ���mӳ�-���Ĺ�!	\>�8������m���m��֛m�m�m�M���m���7M��ۖ�o��M�-�ݶ�m�����oZm�����wv���oX�m����m�n��k��8�s��M�V9,�YY�)�����o^3f��Z�o��^Ͽ��~p�cO�~����t�'럤�G��:3N�3h�0f��2�,�Έc�tgF��`�igJ0`�"��H�0c�(gJѝ�4��4f�њ3,c,E���iђP�:@�P�b,��gF3�&�2�ь馃4f�X�,��t��h��tc�b ��!�1�1�3F3F�<x��yO(��y�,�$�1�C:!�1�1c�b��!�1�X�єtClO��}�5������{h熛��W_��&�+���<�(F�Ыl �D�xH�
e�1�oqۉ֪"��3j���)),і�v�ԛS.��P���1t���m��6݋u�ғX��84L��&��^�LQD	�����fX&A��3;e������69��3�(��v��}_W[N�VWՅ�^;*I�$��e��-ڪk6>_V>���/��i�.U.6.kT�ᣭ��Y��Se&�g�u���]]fw���Ŷ�<7��A�^����L��p��I��6�Ku-�J�M�^L�b0F]��$��l���0�If�����[3��Z�5p_�.���A��E�DV�Yr���"���8.��>̢��1��7�	��p���6���|��0̤���L{j��e9�8<���I+u��|�&�l��H��g�eFh�Gk,�[�n 갵���,ά��u�1�R	@�<��/�l|ehD<6b���ٶB�����Ma-�sBݱn�n��i��m┄&��D�UtzXM6`4Ji�:�3�R�iu/��z̭�9u�S̷�u9
4ؚ�y�I.qg����6��g��s��8n�?/{�m���ppỸ���y�o3<s�9�����y�o3=�r"!hy��m���[Z�yלuǆi�����o���tBPMJ��L̕�DD1K�Ÿݨ@��f{B�v�Z;=Jm�c#�j���M����14v���b�k0]��CY�ʶSj�Z��B֔mÁ�C�Bt$�ϢP��XV6X�sh��-�e�WD?�������Hz>>�ơ2�4z���b<�Q�Ñ�6Z�M����iá�rd؃��i�n1�P��oԢ�uz>14�=���8�8"QX��5l���4�䪦��g��4xSӆjt�É�q/8�.6��[n�Z��0�3L,e�d�Q�b.1JI!�y1_<&��O`���8F:6Q٨N�M�Ce����Xh���X�B�T�s�$͌�A҃#��_$����������5m���jT�-ǧOyL	�^Cf�}��Y7�ͫ&qtm�l��6%=<==c4f�јi��2�2BŃ`0�Âh�JnִM�w��֜J��Ճ��!�a�QC���?��Ac��pR��S�ч݉_��m\M����6�%�0���L�0��a�Qn-���4�+m6>-:M��:9;ղÒ�xF/�D��,4�C��7�f>͔��Ӓ�QCM<�N8ۆ�y׍��1�ac,c$�t�b:��*8����W�<�u�!��io�,�uN�����1��Θc���"�S��g2���)�ӑl��=橾�p=�NOMȟr�4c8L�8XvgG�D��G�K���NP��=�>�͡a�\�4�TK�6ga�X�_4�jG ��:t�����3Fh�4���c%S���e3Z�֩�(���Hu�D���j��9��j�\
mx�#bS^� r����o� %9�k�^����ܞ/���!��m΋Efk�r\�K�lY�>�Y�S�JI
OD��&phIm&�f���14��.�ΏH����y��Y�(��a ����;;���*V��p�C�)���j�o}��aΆ���,/{	8y�a�o�bi�	�D�J����_���LI�L`��7�s��.�̥�Y�v�2���LŢ�e�N�&�2'�SfΚ4�Ɩ`X�h���1�ac,c$u�F��ʡH���	�yI.ân��8��a�s����6&Lނ�m�UG~v��gM�O!K���z6)���a��t�`}"�vԩV�l��($��3����o����9��5���(hC�FC��m��8^9�D����(ZI�4�~�$����3ƌјi��2�2N�W@�*6�\'Jh�_Kx�6hNh�j���N%����ꡖ#8>����s��+Ӿ�I�z�O6�[��@uн�cCCjqufA��i4�o���>�t
a��R|}�1��,�S�ɭ� '$!ŊhJPB�Te%@�$T���D.�o"�a���T���͚4����G
Io !9���4�Kf�f�њh��ь���H"���,��T�R�:Iժa�b�f$���1:%��w�Or�Zz�<\�J����������I�����[��4V��E=�	�8��J�eA���U�l�>,�'{Ɏd��a ��1��Q�dae���3Fh�4f�����I:��|/��Y��T�D[�a3ek&�&��o�f��д�ڛ7>��[`�cA調6Ym&L�&f'fW �z��(�rF�#��["���׹��>��A�SRe]��_�q�����UQr�]�%�Ľ���etD�+��h=$��v��i�����C���j��Vi�i?%�'��ɡ7���Ra⤰�N�!��p�J�H)���N棱U�����B���0DC���t��%�tz3A}�>��M��>�����p����&K=[�4�b9|;���Hj�'x_:1�1�,af�њ3M�4ã:1�G!P^��m�]���G���P�/Bb<�|!�̒�7)y�qi��|��,d?n��Z��j����,���N���cei$�|�7TT�D$��`7��}v�ml�7��=%D����[�`YC�=g����<N]�G�g��3��`�|a�%�L��giڌ;2�f�ߠ�WYVSn����*�o��~y]NԶ:�O�iy�Zz�u�<��+��WR�u6��M��^&�ckU��e]qKM�S�m:Z�g�SqS+M�V�4�eJZ�I��m6�Z�����<Y,�>0�<C4�Q�+FC�A�Q�������^$�#'�Iј��)6N�^&�Ka�mL�V�mj�UŪ�i�x�-XNSi�V�y6���Uiqj�Kc��j��c	���[*��U�\Z�ձ��p�Z�SeZr�al[*����cj��ŧ��ʲm6�ZmJ��	U�L.���G�G�_��K酶��
[6�M��R�u6�M�\Y'Ԕ��_�_�H�dt��>#���<(^��q�A$Lg��OfE]���	.�շ�W@<��X�cv�_�s���to��S��,̧�����+��0��[O�w�]Tn���=ȃ�g٫�6�fg�n��{���癙���z׽�{��fc8n��ǳ����nfi�I4�N���Z�yo-疵��Keo7���WFY��UQ7F��L��UU-����R�*�	[QIIK��i#���`�&f���~�A=���מ.h�"�erD'd��LM�(�#�J�&��9�w�=�8*݁�p}��gkT@�Ӄ���A3�0ŕ4X���Q�t`�����D���c0�D�+R�fbh�I��ba0L�Vb��C<�S�P�'z~0�d��q����B��
$M��ͭ�$l�:07"�qIJRt�Ĩ�`�������RhCx(�ޚ��DBe�'$�b!���&���*�u0�I0���ŚY��Fh��3�4񕭄�&٦���̥)\(i#p�҇����f��JJ<�0$�$a$�I�Q�ӈ2�)�1'DO>�{Ȣ��}��wN(��p8�pc�cN� ��I\�q+��*&�#	��~�I����6|Rc	�~Nas.4�3D8!���	��e����URɻN�#bK	K����2��������-5����7�JQiy'���JXj�Ku�-�i���O��5�H�peO�j lA6m�J�;<a8j����H�:05؛����L�$�L<3O��>�4f��Fi��<t��M�Q3b'�]�u<J�p�"�ƴi�ʪ�A��YV���3K*R��+�e��L���	l�9ޔr=nAcMr�<w�� zے[U�R��`ز�C��O���ao�I}*,�̉�_[���~�� ��XBS�,��[���V\���;;2����ovm��M,,��y��M)�i�ق lM��Q4�0��<wi�Djah�%,��\��0�\K����10�=�z0Г��B���0`�D�3ds�����/�B.9���5�a҅&XDNg&!����ޔ�sF����;��2&�"bO��LL����!F���<~C�3�*@��R�t�k*�rJ�ؤ�\���R��.a�-�'c�с���i�
�mK�JT�l�,�0T+~O!���0�'P��b�[�>[k6�μ�μ�ޙ�-m-lF�Lʨ��n	�s�9(Ȱ�&LR&ZK�JX�L�M�-�P�I�2|'<(�~���)��D��B[��!�)XRRܑ�k0����\��U0l�X�.Ó
݆�F�3 ��,��1�1�xBrO=\�0�`�Mh�$>k�4Y>�Z
q<L�d�B���zϹ���	���#T�QDDNl��S-�3�RcPD���I1�a��jkL���������{
@b�$�0ܼ�9�iMZ����h���'�N��tdЁ��֭�񽆘�JY�y�Q�r�º�LD���AOf�!I�Μ0D�ɇ��k�+j%U	�[��k6��њ3Fh���<Q�ĕԒI"R��mO>S	*E&#�D�JH��7��n�l)�>���hs>=Ԃ"&$�%a��0If��M���'���Da5ҝ�~E)4%�~�V����,�I�
"s��a�bJ��TUab�b��?	\2�,=\ĥ��@�sDXQJfBp�Bga`{E(��8!�i�8��NQ:ũ�@�{ᲈ��Rha�(T���ہ��l6$�@�*Gm�A�E8��D`ꎯ�㙃���7!�'�J*M%��)RQ*Q�jF�Ko9D4I�0��I�y(TҜ���K2�m-����?JV�����Y�Y��њ3Fic�<Q�Ğ)��tk��`�K�w�\��HB9ߒ�h42����g���diDJ$�4+��o� ��H��/��J"x"ş���Ǔ��1'wXbR�!��H�l���fɠO�,<T<��,ٺ(0��Rh�O`������8S��I`�;
i�7
��pI��Y"���YP̟q:b!�I���0̰��|k�ܜ'��Xj'P�Ad~)R)���ϕS,A���გ4���aa�!�A��6!�ᢆ�&�$`�����l��)\�6����6LDRM�T�0�5�%�X�>0e�x,��4f���3<x�ǉ>����E�;��HQ"�q�ȭ�z�t��M���(����N2���m����Ќ Y�lg�n���ȵ�Uպ��7/Emy��vi!7+�p�g��y��M�
J�yj�VH�J�VB�"�ɖc�� $}��[O�zb�9�3c��n��]��s&��W��KyLa���>���ec%%ĸ�R�q�T���jXIp�l��}1$�>���=9$d=�Ї�b�?��A�a��Hv3!B�0DѭC�Na��H���)d�f�Lo��Uo0jfj]K�1(j�!䣹L��L�M�Qĩ%��M��\�;�*��'�D�Q?;|�>9��60�=��`�H�O��lA���0�b��k�E0M�)�&5.�r���\&�g>��PS���<5ND�'��H ��B�c>���z��:�;.���[��6||h��4���(��K���#�=�*�2�-�#�d")��a��4���K�4ɸ����
�d�
�&A?	���>������M���'���T��7P�Gba؜�����}
O����jE<�4&��=��JdIza�0p��LCPMa���x�{Z~�GW������Ob�5�y�+���ql�Q����h��2m(Jb-�_-�!��J�LS��.Q�E�3l��d)B#!Ć�����<)6!�O�LEVp�Me�F	��g�x,gƌњ3Kc ��Ol>�h�UQ$���0�'�pe��P�W���N(��!L0�SQ	�d�ɧ��C�~��a�v7f��0,SG�C�B�%�L7*�X7�*a�&a�!/v?O�H,O,����Sh�z�54�%�LzS�&�(���D�����T�����n���A:SI�{��s9�D尲JM�2��ğ=�\L&��N�ݲ�qi�M�	���ɱ��<ɫ�Ї`�p��C�/ڥ�S����;"O�7��S)fJo�?C0�$�]m�>q�םyםm��-jZ�+����n���������h4P=��G��"�D�0���JL����̺O��Mn�����ZKn�c�Q��x�[�&�s�(��KQ[�$��0��di��Nd
&ć��
].�J%.F����Ӊ&QI5.������)�K�aOXhPfLR_q2�f%��$L��;dW_��p�$�!>���p�=�⊉j3I�<�n��ӏF]�*�����!���J�j���j�>Z���i���c���j���i���l�i�����j�;SKRSi���lZt�I�xӲ��>>��&/�f��
9q/���mj�i��ajJejJ�f���e�����1i�<3Қ�g�W�o+��J�VOi�m�d�e=M��aT�&�Jص*�[M��Z��M���T��+���I���ż��^M����[�[���m�[
���ե�֥��겛eX]NR�&�SKm�[Kem��U�ֶ-=b�ʲ�jU-*���}]���UtT~>���-�R�jV�U�R�mT��8[�]M�Ű�M�i������r���ǋ��%�������9QQ5�T�D�[Fa���5�2M�c]S��y��BW0X�c\�,��]�'�>=<��g0F_a����c1�C�fgv��3�ϻ�0�x'�;M���U���$BWF,x��Q�-�ɫȽ��K�~;��̴���@�ۻZM�h�c�������DL�1ߍ�+�r�'$v+VFڷ��ݺ�kj���o��9���g�����a�AQA��]���ܹm��k�.䕏$�����|ަ�x�*�Q�X�5��v�ߌ��!xm�eK��d�ɐc�6� QcJ����ܬ�������|�d<C�������P0��}R��Ďm�*l��%oM���f�EՏ�1�>Z�'G~�u=xN��b�ZחY��÷�S0]0�bXLt'���T����K���ә"�F�#�� ke-d����n��%��P��sX͛�e+cF�Z�kF�S�����7��z��+Pү�72+��E𻘂G�|�O���L����r��MPۯ{�m1S����z8!0м��*,��YAUY�������.M������ă���,��Ԕu�L}�=H�Kip�����m�c��Kri��\�����Tʬ@��J=����B.��;A3����Vw�y���{ws33�m�{ۻ�����m������xm���n�I��4��4f�њYу<x�ǉ(�a]�q
&i&mՆ��.���BU��M��yOys�P��Kv8YMk��=�RROY�Im��0�س1�,CZc5���,�� �{d�K��;k1عa,!��2��e��[V^��Uf'� �x3�앙��Y�L��$�%Ȫ�ɽ��m��js�#���a����%��1E��y2�_���5*L�:���QIJ�b4��,�6Rl��t�V�jFsc�Oɦ�=�">|�1q�?Nꢥ_a4��7U��i��=�UVb4��x!ËC�l��%����h��Lfx^.�hl�
>��·yU�d)�ی�������t2���6,�Wo�͕�?$���4y��E�3*I�r2�[k����[���L�Kqo����ַ^u�FigF��!����|+$���e:ê����B�y>2v}0�n@�Lף�l؆�{Ms�5m���K4Q=�)�0A)�7��(�6�u�>�'jNCpK!�g�'�M@���<7�4$��,?{<���8��%5�a}(i&�}
��K{�bap��r!/�E���7ǅ�6�#eV�ERx�v��\�I�g8M4�C(�0��3�N��3���)���������&��C �"J���B��eL䊄�R�QI9����ɦ�G�i�{�O��,0�d����-�ˮ<�󏍭n��μ�m<ykR��;\c�L���K��q?!ч�"�ᠩ�^�mu�:%%���0�R�W	DF�0����I�0����Z��al�ɔ��G �2�f��\iEo9q����O�d|gĘ��Z�1ҩ�X.�Cf�L5;�؟����lL�P���(�/7xtF��a��NB|y�B�kI���ؑ/�C��
9�C�Ec�����9o���JeSgۆ1�4�e�����T��"a�AF`Ϗ|a�Ǎ�4f�ta���O����xį?f��������ɩ��Ba�I��z�c#���8�im?����Q\)$u0���1�;i�$�7d&�fIiL	���w��9DUt�!��;8�A���ÓKn&kXr)�!R[+`ۑP�؄T{3:a���<��ۙr�����&d|�C�h�Cț`w�9�����!��hѣ������5mn���L�����C
}��m_�7�:a={��`ę�*�q�>|ӏ�qf�-ם3FigF��rH�TMD*��i7��ZXb���l[J�р���=_�]Z��5ь�+tڧ�嬹�F<�p�ET�L��b�n�2�s�,���E�S�dU��m�ܤ�JrF=����e&��ij��ʺ��hk�!�� I�{�O9�tI�����M#v�UP��p�����V+σ�Ĥ�u�T�T�I<�33�iN4-\`�a�fR��QT�5�OM.�ԛO��Ha�FC��k�����ԔA���r��I�o�,7J|!��ؖ��CBr>�9�A0���nc�ڍ�3X��z�> �2�<{4a[4�tZ)��F�QN��n�����j6j�~4P��<�T�Z��h�-�%�4�-���-םyםYу�'��ٛz���LZ�oj�8pF��V�|8s�UF�����Td�y�!mu�	%韦�3U��KęZj#P��=	>�TfCP�CP�p�C)Q�_Ə���A�zz`�]�������npڣI-i��T+Q԰�4�H�Hk$�;!���.�8��߶G� ���iѺ��mO�ma�*L����� �z!�ҙb���	eK�)#������6I�a`x!ӟ^ۗ0.�&!�i���|ڝ|��q��t��4��3�<t��~%-�O3EUUR��i�0�;�?$�a�~u+\�D�� C��2�P��Aa�B�Cه��m)�a�N¡Dq%��a/Ba)Fx�w��%��s��*����D��x�{̷�ƃ6l�I�&�j�:�� �fѪa�C��,�C�ɉ<ᨙ|=���Ae�����P���_(��@�dK-r�kj�_�]�B�[Ԅ��� TxCFߒY����=�����Y�؂�C�,O��2�uM�KS`�[��i0�0����L-��E���pu<�
O�P�;����m�8۫|����4f�њYу�&�q\̓�UF��jxh��XpO�(����{#5�V��p�\0��e���OA/��/s��<��3#I�w��;K�[��Jb�-��z=���Sή��e�����j,��th�I�q���F��0��+��o�4�ئf`��Z��&w�NOtS
z%nXr	��u&��o}�I�&>�f&>"N/�b#�F[��jp��d��ҡ�g�����9q,�O4��>[�6���^u�[h��G��N-Ȕ��O�L�WT�BBZ��H�A�S����$���Ĺ���i��8��dm0Ah�TD��؎�)H�*R�%"�*�I�>��ge�-نV�2�HKJ8�T%I{Ό y!�Fe� �0 $�4}a,<XB\Sgi�-a�,�m;@K5����~8 i�+P��
�ϡP�>��2�5���;�[��v۠��(���VNGT�L1������:��R3���O�����������C!K[�I��y�zfK�k��Ô��3B�u�O���O��[L���:ɳ�[&N#D������_�0��&'��0UC9i�5я�/�i,:}�P�|s�^����cԘƪqL�,����2���<mkun��ζ�ǞJ���k����f���2K"{&�L(�҇�Kӆ���2O�A����y���v	��l񍓟�����3&E6Q��
	�����'���Iu�����}�n��?�8�\�"%x�"/��x|x�RF�I�*�}>�f�ð��Q%�=���&7r�7Y��,���EY3|�2�T$�jra�m���*R>&�.=��j!�%3Q��hC�Pa��������â��B'l9���13o����O�i�z�:�)�Z|����Uo)��r�uj��ܩⴝ.�&�S6�-V�-Vf����F���LG��/��J��e,0��O����S�Gɥ��+K-��\Z�����o*�kW��M��'I�j��2��f�VV�e<eT��+-R�ص*י�i6�طi�Ui�eu>W�i�ej�j�ک���W����qV긵m:r�r�J׉�iu6��ͱi�V��VSl�e�M�kMM��[-��r�Z��Zz��16Z�Kc	��WS��U4�&ZRS�V�Z��[5Sj���0�aV�M��j��
���m*�U&ɲ���>NS�5?4���+���<��M�Ͽhӌ�!��h�Ƣ��v�Өs(g�8��x�L_,:��;���+���M"�d4�P�a�I�3,*HT+��J��I�E�$9�Bo��q�8����c�v�mp	˞B%.{�+�z�>�������x��v���ߟ~6�~n���y��y������6�o=�������m�{v$҉4��[�6���^u�[i��%kYM���2,�n(|m��Y'���%������:���	vN���'D)��~��Du�J|Z�43���2��{�31�K�u(fR�g��N2��W�fS-�.J쩊D+$J�>fq��%�e����Q�'a�fO'��é�����
2OO!���<����eG��'��U]RR�UJg�C�
�T����1)L"YɆ�0�T�J1	��)�*��$��a��8���ַO3LgFb<x�5%�J��:I�
o�UD�CӦA���ʚΎ��*䣰g�N	`���aȘ��;2OM�-p�MA���C�{/�����tI��c+�>)8�j"/���%����v{&��4~,М���
�7�0Li�����,��	m1q�D�ĜeJ���fRURq�feL��}
iD��y�\��+gFҏ�)��,ɇ2,�I�$�a��n������z_ng'��a0��Ϝu�<x�ƌ�Yу�<lW�	S,i��}ٳh;���{��®���]��W�/�l�B[kպ�ؓqK���4V�]�z=�ad9��r`��wr5�V�U��Om�+�:�il����8�	��G_y��(�*�����%�?  ��M����"e��d�\,���JS��l��}>rE�O=3-1��aԹ����LL40<�_&M*[mn%CF�r	�@�d����lf��!�,����?mЕ�lCJ��rZ�38��RҌ%�����q0�N��S���b�,����J*$�`��`Q9�ߍD���j�>�60D�'D�A���<���=��hN�y��j�6�0pd�#dB��U�E�6�^����:�pޕ�{l��!D�������?kc�F�$��+�"ǚe��-ǛJ���y�^m��<��l�1ȈT��L�nÕ���R�D�d���"@X2
���E7�*���CY�Na��&0��I���7�`�9�	��~=��)�aa��JP��{�܄"tN��k��\\�,ĩ��+��z��"0�[mhIT�WlB(F��IX�Ym�e�`�Tcж�،JZ�Z�Z�m������%�/LJB����ꑣ�Y�&�.�����D�YkIDb W���)=��/*̜��AR/��̯��z7!��N\��A������-�A�Y��F���1'RB���w�#2*b'�kO�d�&$��2O���m�Vh��d�Ah��Q����j.����ꛦ˙mf���4ִ}<��22r	O
n��%�KE��Y��Dꥇ�0�!��74r��~�-#)qp�C��4�8�o�G!�T�!gĒxg�>0��<i�Fi�,�ǞJַb�)U*������Ii}ǙE�9]�͚z|Sv'�$�7�EaOڅ��'X�=�w
����5L���%��м�[�ȉ+�����Sn�bk4�S-�U�y'���D0d���=\��8&��`�g=�[3�8p����2T��!`�?OHK�M	�K��s!��|�i�?	񐳂G���
����"�D���<(ta�4���{*8�L��θ�ĭn�םu�Ό�3Ǉk6��O<�"h�Iw"W\0�y�UV#!��aN�L4xP�pOD�����C�d0��4$����~A�,:�8�2�Sa�'�C��f�D�밨�KВ��b*%Ĺ�ϡ�cCIs[�C'��}�wI;��	�p����ӳLV%�L�%q���6�"x{�����<��sTSf#х�[��i�V��J���y�FYу�x�M+���V�ҕD�!�	4$��������He'�JINŭ�æ����9����:%.��"b�rJ,��7[m��ƪL��[LFufW\]
�e��� 8����TW��=�C4V�ƴ�Ub*��6Ogpή�e<6&����Z�tl������Çe�l�y�D������؞)D}�t����b ��'=t:����sx��a,2�R֑�K	Xp�~lD��~�5��D��)mJ�m
�paT����-�T<돜�4��S���[O�}��U'H�V�ַyǜK康^uכi��%�Q�l���ĥ���a⏺c�p�
���"
|�\�M$Ft��N��ګiLr�a�_>������jd��ਚ��� �{�>D4.aB<"Γ�Zt�;�b��cGnJ���Y�U�i,8�T�%-�fڞ���F">q�)X1�9����<��{ʥ9;��Ja]i��[�Ϝ|�_-պ�Yу�x�pd�'�$��0�R|k�)Z�G��<�r_!�p�&�Xu�R�n~rjjqƜI}u-CF��i,������K��k��o)�P�2���=���"p�~޶t9��_���-��Ӧ��}�x͆I�?$�X)=�%���5=�v*��4���ɔ��2�354�����%����>w�4��N6�����%�-պ��Oy/-mT���JXV��m:�*�y�D�Iu����a�!�}<�e5͟�e_+��Q�."�ץ-��wb$G�sG��|#�/f"z`���c$��4�"����0����yL�xN$��Q"3��}�R�k�1l6�Q�Ӎ0�1Й���~��X�34x�&���$����>��,e���(��/	i�5/��P��u*#�#R��-��q6�'.1��:M�Sj��*��j��<�|­6�'�+����X�����>.�����ZZ~/�(> �Y�6|F<iH�4��Y���-ڙ�m�u-'m��)i�VҲ�S.1���$�j���6�ٶU���l[������+��J����Է�b�Rީ�e�[���n�i�r⬟&���i��ŭV�a6ʘ^S�M��R�j��m-�&Զ-j��gbV�Z������+T�L���5S4�蕦V�R��[2�bXU��M��յ��mW��}]�>����~������~:|O��*>'8Gq�MG"Z��{u���~�˯[in����@����}(\ƾ��[1 ��a+ڧC�L�QN��$6��f�H��L�-YG�8:�m��UL"����7+MUJQ�L����45l,YV!fE6n+��i�B<Q��Z*��`,�+6����@�����N�x��&��l�R�exD�R���<m�>j��L;M�nn��K{���e��=�֗�5͉LK34ȳ=v�Y�<�'���b�z�Ai�k��푻Hª7H�����P�M��Zc����Cl���6޻Xݷ[�T��\�*l���|K!s����6�o/um��/��7%�S����O�\-��&�2�ɕ4�4��O��r5�u�1�f�.��v�T��������y�|���7;��CW&����u�o���aތX6�2�Mvu�-����R94���;�S��[}�i����,H8�,��n��k�k�D���8պ�56�t��m����a�eQɮXֶ׋gm�nv���TN`G�#x�.g3E�i��qan�q5��5�F���譻L\\�m��vf�v5��\�/�x�2��Ezdʚ9^1�"_�)��~���ͷ��������osۻ�����m��n����^m��=�&�i��i�#ǆxњh�:0c�"MG��|��Vx�����뭕����F̬u�o�.ۉ��5���M�WR�X��b,Ĳ݊E�G�URc��1�ƤR���mM��[���9%JV�T���JF���Bn��� pB�PO@_���Q�äs-�"���,���啩���a-e����e"4�������
�!��$�3|�Xպ'd�7�xy6�ӯ�m��k-}	�FҮC4qu*'���gDOL<��6%����Zi���B�r5cg B����Z Uo=����U�Z���Tҷ�u�neŸ��yŸ�����Oy/-l\gЧ7333��S��I�L�߽���`�)�m�D���9�O�-����@❲~�f�d��}�����؞Mß+94y)D��e��M�X�uWWl��o�\ˌШ�5ӝ�p��tFzQ5�����>�t�%:p��OX���د8�")�q�]y���Ϝ|�V��4f�2Ό�3ǈ6�x��1���p�� ��xЯZ��ڪ�>�Y�Bd9��t�lû'����)G�z�^I;rbk|a)���i�a��O�f~.y���N�dX�6��j>����O�fN�)�щ��}�TMuII�'�c8�)����!��DO�N��^l���ʟ������SI[-�._�R�GJ�iu�vhyd�|3�>>0����Fi�,����OOO�xb�[K�*�Da�E�{�ff� ü"���9m�5RZ�d�3aIk�Jby�ĥXٷY�Ya��[t.���ڨj��D�-�CRa��|�pD�y>W��~Jm�T��L�艨krt��n8���H��Gy�=�F���,��Yz0͓9}pp�Z槫B|�*1�=!҉���M��W�J	��i/F�����ì)�>i�Ϝy���Fi�,��!��F�D�5�a������a&$��U�y!/�,��C0�$ݗ�8������>�̾c���{�&)��=1=H�;�a����L����m�Yg����O>�Tm�JM���b�]�ls�k`� ���5<J�"�uAu�.-ԣX���IL����52���r�6�N�f�Y��f��Z1{�l�x`�Cp�m]O}�]	�gL%p�m��UL9,�9�k�<��w��<>0�W�e����.��Jn��y6�Lee����N�bXa���M|�~S�3��o
�5p- 0���6���f%���=�&�a��6'�X}ӏ��±�1��\G�e�m4�帶 ��3MgM1b���������Iq��,�p��
E��K4Ӎf;3�����Ĵ�XZ�C��k�nrpe��aa��%�'	La,6l�[���j�QD(�DQ?j��f��[�,-��� Q[l���\ă٣�_N�l>�l��-�Zz:"׻�N��L�*��0�0ӉO�N$(�K���E�>:||3�> ��3MgM1c�v�D�uJ���V"~���6��m��b�fΈ�22�8a�xs�}��34kG��8�!��J��v�q��JcPê!~_��� ^ �6)J7*$v�
f�s"5O'D���MA;�s�1:l�G�}60�#��Ͱ���|�W]�E�X�b"H�NH�)��Fe�K:�<�\�3=T��6�9m,B�/D��N-N%�1,�a�ᴸ�Ft���a��xњh�:h1�g�Xk�U����"'�E����5:lM�0�9{��r�)��b�K�@�u�)I�>�<ɺq���k��a۹��yԵ
���C�F�崷�u����;�R��i�q-����|�;�����Fj����U��H���Z�(���p��[Ū�m	����O-ǜZ���[�gM1f:�DȡNt�I�ZO.[mگ�=�<3�V�Dc	�C��;���Ӫ�`�ɶ�>�%<�0�T�8��:�3^dRnb�i̒H�͗�G��E1Q����D�V0�&��M+�;:b:����'hX˸���� �x��:5�Z�V*���h����\=�_�����Y|!���?)���<U:&C��᩼�4+�l�������<7���B~g��C�d��=+5�sYkF���%ؔ��S�/����4�`9�jdf0؉�~[|��֥�p��ߗ�z_����0���iU�Mo�'jh�)�i��u���� ��񦌳���2s��׹��y���MC��х&ᇞF֜i,0��6�t��uԾm2��<Ӷ��g��%+��O�� ��Tώ�l)؞�����Çv�a�p�=K'#�aD���npµ��{ie��9ֻ*w�}�m�S��Λ����:L����[�CP�~[��K�VsZ�D�a��n%1�1���-˩�|�ކa�\/�u�Ωź�4f3`�0c��h�,���2L)��h� c0�[x����yL��$�Iy)y�Զ�Z�qm�n4�yםy��4f�IӣєH�Id�`��$d1�H���f�f�1�4�� f���P�,c0�$�4фcc��I1�c$cьC�Qd�3�����e�%�ǞK�yN��@�1���c�C�$�G�<x�g���CWx���]�'�4�����2��6����۝�-�dܛ=Q;\�۱�EW�|��w{���������9o����X�`ѽ���oqm�W@�N<�y��f���6�=Lϧ��̛h�I������_ɳ��w}��ckU�O�g���y0�����os=�����m������{ޏ6���n���G�m��H:ˮ��kqn-Kyo-�^m�OC���$�\Bq��L>i�D�U�0ƧDM������4l���ɪ��Cie�rr�1eӍ%������&���v�z����I��v�uJ�x���ЖR¸L%�����4�0����Ɇy	S�ʛe+w�T���'P��\m���4��3|8~���z�����(���9�R;����Ĵ��_:��yũo-��ʹ����b]K9�6������JaY��S�w5im3FϧN�'����A`�"=Ӥ�ѽS�4�Oj�0���k�h�t<:u=P�����tu	\��F\d�9e!�hy`��r=6<6pK��,3�iJ�^��/��Ul$�Xꡖ1"m6��6|�g��ᣆĥ1���ϛy��������,��!��ޓ��V�"#�J �T�Q���d�A�h���d�{��s��9���ڜ��<%�T֠�z��O�2��'����K��aU`�r�rQ�p�nI�V		�m,�k��m+� !=�\1)0t䉑�����lV���I������%�0E�E%���4&O��c[�ْ��d�qItj"�Me��N�LN]m��q��S�/��u��1Yb�)m�.��&�(�X��O�U�K��eO��2�iu�WV͵�ҏYLe�<�'I�t63���)��Ӈ���US��KkbfXy�iך[�qj[�yn��m:��y�T��Oʫ�D�Ó���`��o��L�*e�х]����:����qK��p���oDq��-ˌL����I���M���pʙ9L��fR���`��ֱh��n�m�5v:��>uؙk	KK}�D���q�	�8V������ C!�R��Oj�E]�LMT"\� C�����0�$D;&�v���]�)�h�>{��TL�:��q��E��.����yǈ<3�<i�,�&!�����I%?'��WӒlD���97�.8"j��:3�E79<�~�&f`�O�=5�Q\�,>2���z! ��h^_���d�XHH)���K��:е�?�͞���l>6Ju��(�_L��+I�0��T��X����g���fQ�>��'7S�Z�F�:�)��,>Q�a�E�&iX]��u��|�Kq󏔷��ƚ2Κ1�c"{uf8�4L��I.!�g�0�7��M���#����C:���2r�%s�1�\��
�&6�jq�CJR��R�ii��"���q�L�
R]�bf<O���K���bϛ���e���*9n;�(����"R/�ʄ���p��h!���i��V��:�ZyŸ�-�n��gF1�1����,�);]��{:q1ci�Wrv��rj��4gq�=pIn6 N��̨$�9�i��h����%�����uϬ��ҫⷓ�1u��|Na�X5;��ҦSiO��k�kao^�v��5�N�WN�� 8!I�~hډjpP}L�����J�Y����3ofknm�j�4���G��V��/'�?�pD�>և����y����n�.�t��0��s�R^��p�K�p���i4tD�S<)�~�>N�8l�l=�������C��F	���-N�!{�&����`�XUk`��a��0f����d<�v~�	m*�*
9M铱�u.���ç����Ǎ4e��@�W�UDDѩ�&�Cʔ��M��rt���,8m&ϼ�zffT���s|E2��J'6�BRd�V�L�f>�BQ�5��az���=�b�-Yn3��b��t#}.�~3�,����崧��a�4z,��J�;����3�s�&Av���5�`�l��Z�[�qka�n�2Όѐ1�K�� P)�����S3$�s<a,�h���M��ˎ�ӛ��z��J��E��Wܻ���Ԗ����3'���V:�#��4�W�ɓ��<�=?t���3|�>3��V#m?~E��������8�ff6zI،�K0�t�����E�0O��?�٣a����^}�y��m��i�Z�yo4іtf����=i$�iUĆ�5	K���0S~�jf��X`����Lƅok�	�&�X��q�4���"��}��ҟ�3<4�V��O�P��b��5���jy���rx���0]����UIU%rp�8S��WPö�ѓ���j�����م>Q̷"9ϒ��<"�h�0f��3��4�i�0���`�1�tgFY�:��q��x����yL�/#�$�8I�R�#юţ0�ƞ<te�l��V�l4�m��a��Si��1�:!�e�f�f�1�Ӧ4���2�X�,�+e2�1�C�3F1�0d�@���2F1��2Mb$g�0����`�,�,�<�L���C�2�1�gD1O<��al��V���s��V&[Xq��N���[��`HȢD�����j���|�Mm��o�
[%$D���G�^�g���O,�e������'��h�&��o�o�3�7��z�w���B���F�}�F�f1i�㓻Y�TM;f4��Z��]�Acp�\m(��ږ(�.�������v���!��.ooF�f���+�/�T�	O���16���>]��z�����K}��F[��eQ��#��U���z0ɬ,���F��ZV�� ch�$̩,���m���ix��O�����T{Sb�%������2������V��h>l�ɲ�ߜ���h޺X�-����.sƻLd�k��q}Y��� ܏h� ٿ61>���ġ��1��J�HWZ�
��I��'#�����o�m���"�����o�?_X�}�B����\%�,�9+��U��r�Vc�Qdt5�7�'���ݱ��)#5/fo�m���X���pܵ�+��_���#��e3��Ѕ���.���,[W<�����Ϛۙ�^�ѷcrMĿp���᧮��1���H���-Cr�Iʢ$+e.�A�R`U�b:��!7��3�2�]AnG�֣����ĐB�Wܯe�6�{��[�����m��{ww���>m���n�����ͷ���MS.��-Ÿ���ַ]y��u|��|����j��!v�V8@�1�d.mz���,-���4�bRn��f�[m��m66��p�2ʗZ�4S1�)��˰R�/׵%]`�4r����;� !=`���Jk�[{u�͵�J�`H��*T��%A�ب'�u,�TL>���P�8ˇJ*&0����B�R��Ҿ�1���3�O�zg79�%s�����$�<$���Q�e�O37���	v�\�,�<~�e|'y��7 �O ^P���W�%]%��OCF͞
&�]�Y|��U3S5��:󮴷a�Č��ƚ2�h��&Є#ت�&�z�?&�/2NCFCF�a��!�0��rc�F�R�#��*	�¡;"������F�4ns�n�qa����s3�~vb�s(�n�1�bL����z|!�gb�����gD��Ӯì���2�C�����K��g>4��ώ�a�$g�4і3F@�)%e.\Z?*��C�pٳFh���o��l�M$�rfqf4��%�i�L�&}�iSJ�u�*UJc��fgl�� o��^�?��'Z� C�}���\2H�U@(����"'�O�I�N�~=��������鸢�C�4	�O?�+�S'��,�3N�����V�C�іa�y�u��J73ƌF"g/0��7%�]mז��[�[-kuն�<ç�0�c��U�ºH���p���h�/솏����{�o�N?�����[�s������w�xn�"��T%|�p�%N�Ia����7�h�ZN��4a��,�����g�'qp�b��^T+T-Q1�	Q�L<�:�m0��-�\mn-o2���V�μ����q�T�z� 8Oy69  JK)�ڶ�D�ٙy$I���$=Λ���KS�BOb��u#5ɴ����je!�ƅ���3��b@!
]sf�֐�Z�'$n�^E�� 	
ڴځB[&�K/Q�X˕t.�>���ذ�S����	�0�*0�<�;���\�}Á�G�R�c��P�9(֚;hrU��K�{��+)����b*%�^�x��o�&p��޴�P��c��uQuv+�Ԡ80�t-�S4�V�۫oa~
M�a�sw�3�G��Yc4�ǌ,��Ǐ��ь�yu�P��F*"f�x(C� B�q<Z�6£�e��Xa�wfZ�{�&��_y??(�?d��e�)�c�jU3S_b&_-�t�b|�d�3
*�-]m�X��{4o�S���r,zr��\���06q���Q5�a�o�4K���OB�g~��&4KzLN�1���i����[�4���Z��q�^y�Y���ت�':4��n�R}��~�y�LQD�)�>[�/��I�m��KV|�ߋl�q�V�j�O(�$)$�y��Q
%�̾�LQ$��'�8C��=�ٙTʖ"�6^��@��RJ8�Ƴ0�I��K4k��p��cPŬõ4i�R�v찉o&���L�FqF�˚R��&�9i3nYu�#��΀�q�3V�1��KYe�����lB̳X ����Wkn�?�j�Z�)�~i�.]x�s5�e�v�W�w���?6��4�7��4�kcF[w��B>�j�vԺޱ���~�(A1<Aֶ��K"�S6q������gx��!�yf!��LӼ'��i�>����u��0�-8��q��Z�ik[έǝy�v!�A)%$G$���VE�����LT��c$���a�
�P�fd"�N2��td����	��&U�!L4	���t�,�|�z�KN/ꁅ�jHؔfSFY��j���d=�,���A,b{M��-{4Zr{/�ђ�a�yP�*�GTF_DI�e�8N\8��w�q8�!QI�"e�F��yKZ*�lٸ{���ha�8SL�|�n���qm����ַ�[�4c$�J���.�*u'�wS�����(�u�c�~v���P�J&���'��<�I��M�K@�jF+��z5V_b�F��g��#�EJ��I�k��ڴ��K�pRE}.t�]kM5�\rD'�<U���@ H[�	� x(U#r5S:��"9^mdԛAz}����Xt���Z��ᇇ��*��-�釣�����r	4�c�eUL{�a�W%���%��I�SFԔ������pf��l{���rϥ߸hQ}�
�'��2�XO'�~�o���˘e����>��`�t����cE)�SX��,gŝ>�`�0��<x��<`��4sQ���S �J��rB�ON��Y��a�p�e�j��i�]�c1Pө0˞��T���Y�N�:	�^�Ξ~�������g����nM�ǜ���pJJ�)*E	_4g0�EѴW�r�1����u���e�ZrS1\�C0�r�Zq��x�^qǜ3`Ό0f�����Β2���2����4f�c0��2X�1���0��IGIΌ��33Fh�3A�i�/Qe����al4��ǞK�yď�te1�3Fi�c4��ic�c,��Y�tC�c��6�C$��1���tc�(e�`�����0a�T�Oy/)/:���c��2�0a#�3�)m8������S��50Ģ�3)
�V���y�Vj�2oVg��4�X��c*ORz�m�&�G����dMj�VH�`m$�d8�J�)&!�%I1I���B��i1��mb�~Gz;�N�"=��_�?z|�{�������O�owsۻ�����m��g�w�����owQdx�x�Řx�Ξ<xn�ǝy�^�ffd�q�j"�Is��C<��C)�>�����m(�c��%o6e��*]�?iȲ��jV���O���a��\.;	G�/�����2i��ì��!"B�E�#�P�jd���̷�SU,�Ѷmǟ-m-��2�<xgO<3O3F2M�������XS~,���kYQ�aHؒ(�F�c�3��"�A5�Ү3b.���$`�O��fá��Λ=�t*Ƨш�G��e�j���LL�l�4���	Za�5�Ca�Q,>�bj�C������3���Y}���)��1�i���k[�qm����ַ�[�:�_(���M��2�V�nÐD��h?,l֒ÂO)0Ǆ�;K��m�lY��	�3y7h?3SOE[����6R�6�$�ː�-f[��4��t2C�"0YDk5��T�0i��⪠�����42�GLº��M�YfH�F�����j>������mS�ڇ$��8S��l-N\)�LL�!v��Q���Xc��tѥ71}L�=|q���PTf}��i1u/��$i�3�{�_�%�d]��n�~��m��1>)����:Mj����� ���,��O�<a�,���:x��x��1�wt���T�U�'!�,�~��h���>;CSR!O��Knюe��l8'NC!����71�KE�T�*��Ѥtl�m.
�M w:��GZ5[$D�<
Xv��9Q2��l�91258�9�S����r�J�IR�jx\(R�M_~?L1�)�6l�C
h����Tl�L���j��n0�n���<ه���ǆi�h�I50����w�S>UUO�`�X�鰦��ҧQ+���\��3�E8���1�ɖ��0��ZG�sWT��M:[-iM1OI��|d:<<�}�rj��iI�#�K�5���I���>�/f����_
;��K�n�V1�\8u쭎CLF�Қmn-�2�<xgO��<`��!M�Ptc�fQt�M�"�� ���&�iM��?~0�h󏊕h�.U
9���-n��{6Cή�>�h�֫R����{Ko'C��DBV��,��TD(�3�&)(�8�*�w�4m���*t�O���ӹ�q����L:��������yn<��8����[μ`��.v;Ɉ�&GI"&#"��J�%&������uId,)�cl[ñ- Y��4I��w�ySQK[]2<NH?�وZ����~GD�K���f�(34�13�MuXd�754ݽ=�U�=a[L�ز�� �ǳ��.�p�"*��[Uu 8�U�Y��F!�`��fWɟC��g���?E��4�>��Ҫ�cT��ᅵ��1|�F�"D���ȟ��y��=�Ӯ�:�����M)�U�E����U�4�H�1[Shm4�Eո�/�{������"#:I$�e�[�4���Kyo:�u�s)L1g�UPF|�l���jy�S�}��ٚ�.Sl�p�q���q.�W��y���{7���s���4*҉Ѓ�N��|������3.��20�,��M���Der�ʕ�ơ�ك�F!ž�f�}s�U$�e���y�ύ4��t�ǆt����ь�߶��"3c�;�J���Nxt�yQM�p�}'CF�]�����5̇���	�`Ss��E;̓����ݯ�|]�Ԕ^$@�emMM*��u��mV���<.�0G����F�D��^D˓�p�÷���8�18��Q��I�6��,����xf�0fd�U���MS)��Ua��P�͇g��t�CG��m~4�7�w��~R��u�V9����E����S.;B[���e)_2�q8���$۷3���m2�j*,q�a�56	��5�U;V�Ӂ�DU���e�!�Q��yٙy��-}�Zw��C�?%��0��4��3`�`�&h�(��ac,�$���Fte�1�AgF4.3�1��	 C8��2	�:H�tc,��њ3Fh� �FY����e��ژR�-iyO8��:����1�3F2�iјј��u�����ѐ1�����1�t�E0c�2�1�1�q��Ǐ0K�KǏ0a�T����0f�dd��1�3FH�C c$��ļx���W?d"�B��
�-,�4�x{"z�de�U���JT�k�g�>�P`h"�-+B����`i�x��sl
j���,�"����n53�p�D��"�-e��I-r��(����Z��!�yr�|�5�-�,V�euZ:�|��V�Dc�����R�i��3�e�Oaڭ�V�;�לyu#�ǯ��e�vfB�D@E���M�[/�q	�Y�U�~}��Ůl�S*�oMϷ�4���Y��I���{�n�,#�[~� Ϟ��g���m�;-�،���M5�XC]�}Y�f-�eH��e�	K,�7U��Y�g(Ѣ�j���"@��&?�}�f*v����H���X�,G���4�6ݮ]|�!�y.�),D�����=m].	��G������rl��)�ƿ���}(��"سB��%3R�%���fq[�Ζ1��'�)��B���o�̴�e��R�p��}�Ǜ��ۥ��E���͛�k[5�Ƙ�X͍*��0c �i�ЙH�c*fx�]W	���2�9�������F�6���*�%�͡A����P�3�Rl�_WD5z�f1.��Y�R_-{͙-�3[6����O
c��6E*o�7G�EY�,�]55�V������^o3�{�{��y����g��{ޯ7��~����{���3,��<x��:a��<X�������lR�"�����=H�#GYl��駯�K�ƍMt���*�ZEQ��Yl4���m���,�	����bRm�q���4����n�6��m�q=���ko�`�)��;jD�:ZB�[t5��mm.���9S���  ����(�k�����*�l�M �߳wY�'/������)���z�
��0t������7'��~0��S�)��#'~�E5�F�+i����a�r��jkq��̶���b��$|��t����Ӯ��_��b#�*�9���wh��i�d?mw�?����&�
O!����FT��=8p���8x��x量�c<3O32JV��˅��8}⪠�|<;��>e_��Ҝ��Je;JTɇ�\���|�[|�.�mJ�<8	���V�Ԇ�838�خ̇�D�k����ΘwޱF�PT}����EH&�"��WZtm��ߖt"W�Z�s��l094��mnd�V[K���bx	O�^�'���0��~��&y��L�<Ҙ[M�ǜ[N-o<X�������BB=i$�T�,�NMO��e�bt)�Y��9��p�:��Q��j��Zm�#��������Ղy�(4r�4��5*���[K��o��~�aã��?~�Kh���NCJm��~㚕15$�K���Ҏa&��ý�g�fe�Y�:>���؂a�'�a��3�L0���Y��<X�g�=<==0���i����j�S%�X��s<m&����t߬m�<���cx� �7@k4YW��+ܞPY?���,������ӓLV���Ç'��9*��'��u�[4��G999
L63xi���E7r���/�uFN>`Y��0��>0f�0��3������E���B��L�r�him�@@�-v�m�ܶ�N.�Xm*�3@�ڮy2��R�i��a��Vi��d+y��:�e���.t ��:`g~� $#��-�������j�ľ�_Bx��>���8�3�/ܵQx`I��x~�I/Cn_e53*��{Q2ۋi��г�O�Q��.�W1*���sN�d��=+���5��=3.46�{����QF�P[�fTEE!���PM��؋�xxt�Ų���\yո����y帷��sy�!��>Ҫ��M���+���S�RtS-m֟n>�4��i0�4ŮfZ����\iy�~����_aa�t)pٟ	�LA'�a��v��Cl۲�4�\����ƶ��y�h�2l�<_�~��p�_<��Fh�]��8�MaUyUn/��;
ql-������g����1�B���HMGw=a��/C�a�}�X�3��Y'��h;�be�Ję��p�^Ց>!T����
~�Ɋ�q̈�M(D*B����P.|��O��y�m������S�����zd�1�8Y�z���u��D��#R�c)KG29V~�qn����䯈Q|��������=	|�.5��6��غ��P�[ϟ-�qn�ż��[�-Ÿ��0�b�fffI\2�)"�Ӫ	�7k���jO�5�~Ģ�݊�쌴q����Mz%+��JfU�S5f<�K�%�Z�+��8ͷG}�댦���-5^0�IT�-�513�Q��a��C�:#=���MI�<!ED��:�:��q��<��[�3��1�RQܨ8�q3ؙ�E����|�tIu K���d(�J�%x����h�M}I��4�0�tD-�bX]��M��v�[ikoS�~ !4��U��v�E�F�ͺU+5״���0�����r���㇦��
�7�"-�Cd��&j���p�o&���T�.��j4R���ja���>��l����KX��������)����:n{��SE�
}�
����<I��><`���ym���[�qo0��fffIK^L6��m(î�\�q�5�a�.��]�<�D�O)M�p�p��vbf��V�p�a{��*�52��N��_����R&.�&���)%�Gx�(��6kG���4��i[j��V��<=����Q8%�	�'���T�D�N6u��y���S�:tfј1�#h�(��ac,��P�d��`�id�0`�h���C8��2P�:3�:1�i�h��4fX�X�y��O0��4����Z��ƒx�㧊IY�3F2�iјј2�gX���t��h�&2�1��Fa$2A���33P���C��DQX!�1�c�h�"0c�C<t��j��.��/ePc�e+��NCZ�0�r��M�����	��s#!Fg;(S��t̘��*��������{������{����w�33/��{����<�̿g��{��|�30��<x��4��F��[�6����O%)�����̒��O_����Mb��9�#4�ɻ2�jp���lv�,=<t���MO����;l(�]E���S3U�����Ӽ1г�#�G�%LD("fS:Ws(��H�W��|�-��h�6(����P�����w��賕���(�����3O4e���y��żýTMR�{����I�Gש{�[�����28I�D�EW
���n-��i����艬���4�QK�њ�����{�̸�:pNC�ӐgS���ߛw<�Cǝf��V�v��f:3ʩVa�X ����Q�0g�3�3O4g�ጳǌ<2I�uݛ�r�E�Q��hZs-�9���ml��KP�^�Z0���é�=�YvRc�� .M�&�X�8��&ga�L��VS��f��ؖ�nlNo{�Dd��bʇ&f=��-�)Zڳ� #��[��Q�q	�T��aH��cYs�i�F���ð�zd?��C�hJ_���{:�eZ�d����6K1NBٖ����a���8��������_J��w�����J���uE~�_ќ�u�T'��MrdS3T_��J)�	=�tiP���몆�z�b����i�L�3O4g�ጳǌ<2I��t�mu���UA'?5ѳε718�����p�Ӭ�~iIdʜ}�q7X����uS�Na�KQ)E+}EY�]�3���*fJY�I�O��S!I�7疮%]�k8��z[��y\��xq�ac���g����ԴY��hFf��sp�4xQ>6;�a��QJX�QL�Yr�Q�v"W
����iv�\|�m�|��[�:��g�a��ǋ<2Jh@��/ZI%$��̦u�O5���Tb��Ou3M��p�L05yom��j1"l��B�/�wn&8��iX�35L����ih���jS��с�Zn	��-_!��9��ǇC��a��2k���QÁ�a����R�vbM�{y��Q6�8|#-\4�����2���-�Ϟ[�<3�,��'2{�G�$�@͏���j��4zp)���j��}
��x���B_�3Z�	�֊�Qq���y<9)�9L���{ga�hbL;�|e�!釁�F����|cŷ42y}Z��n��<5�ܞ͇;��-y78y(&�!�F�
kS:r6al���q�[�3O��4�ǋ<2y�Q�ډ\K�R��20뷏v#�d��H���k����ǀ���,
6V�L�N���^+s7�۵�7��9z�6Ҁ���UsMItՆ%\���0���+��WG� ��t�A{cK�Z�k�X�������ci?V�{	E��:Q\0�o5%A���o�L��ó�3�Ԝ)�;ߙr�EH|0;��^�lJI�{�|A0g�������ޠS~���4��ce��J�u2h+w*~���{��\̼b��k�)'SZLޡ����Z�yǖ��uo8��qkp��Æ�J2�_���kŧ`�EyrL��Ƕn��u���-{��)w[]C|]	�8�Pz��d��v_���Q
%G���$s���`�'n��F�>c2�N�7���ʆ�k9�4ȥ[��2xzf͙=խ��C�a�;��x5���eg<A��1�3���-�\Z�Z�{3�%UN13y�:��C����_fz�b����e�9�U��h:N
}��/����o�͞ü<I �i������(iME0
*aEsnPp�u�^�x&��=��z5ë��c��z�I�Y9�S*��a�be�E-�!��%�I���e����qkyo-�[θ�����je��,i&�uU-æ�B��;0�g��ym����n����#Ph�L���9"��U/�-27�7�׫}�72��kB�O��Wϑ�e�q�GsC-�i�R6�W��.2�C�;�6��Ħ1�.\B��gS�ݝ�Nן�m�����iK+���(ѳf�Ç����S?Vv������s��g'$�8p�׃l6v,f�f����?���מr�o�G6H�A@�C�H��-�D���%'d��	I$���B�I"B�"D�!!!dZ$H�BD�Б�HY"$Y�"Bȑ"Bȑ�H�-�F�2D�#H�mD,��#H���"B#Z,��d,��d,����5���D��-)��k""�i6�Q4�dI"ȒM���Sh�ɢ,�D�D�SD,��I5��
�$B��D�D�i-DM�DE��k&�Id�Md�Mdh�ȓZ4�,��E��ֈ�,�dD�dD�ɢkF�MidH-2Mh�1�I�4�!d�E�L�d�$��H�H�,�$�"dKIY"IɒH�D��$�$�-$�d�$���K$�,�$�IZI&Y���"1
�o
DDSIY2I�[K$�5��YIiL�$��$�Y$�I$�H�ɒH�I$"I2�$�$�,�2KIY$��d�$�D��$F�Id�$�$G(8�$E�$�H�d�"�D���h�Id�#Y$�%��Yɖ��I"�I$�%�I-$Ii�H��%����$�i$�F�KI$ZD�p�q�&�bL��$��MdH�-,�$��ID��i5��&�DII&�&I$�I�I,�I�,�I%�����ZH��D��$�I$YIdšh�$Y$�i"L�$�i"K#I�$�D�L�Ii"KL�%�I�L��D,��H���i�YMi��#nKD���kDB�dMh�[F��H���D�0�D�D��5�XJ��C]�n"b �2,Ȃ&�lDe��p�D�E�-�&�L"a�M����8m�ab&ȍdLD4M�̎|��-��E�DȌ��1h�Y��Dȱ��D�[4[3D�˃�9�F�l�f�3E�#h�E��&p�#h��X�&ȘDm�9C��[dLD�E�dA��L�"�E�XD� �m��#�8٢�4L�6E�M�m�Ƌ6���8C��h�"6�"2,ȱ�b!�L�l�cDm�d[4FD4F�l�f�f�b,E�,4�6�6"Y�CDm4[4i��"XȰE��lE�"�"ͣ[4[��!�h���ȴh����H,���"5�H��АZBB�qhr�!dQ#Z(�D��dbА��!h�!h�H�Yh$HZ$HZ$H,��H�Y�"B���"F�А�e�P�h�!dH�,�$Y$H�#,�	�dH�Y#HH�$H�"4B�z�"D��H��$HYD��"BȢ#HY�d$5� �H�u��!h�""ȑY$,���",�DBȑ�,���A"�H�[D�!d$H�$�D���"B�$$Z	,��D��Ȑ�h��drFp�!h�!d$-"D��"BȑY$HZ$D,�"G7�DHY4BА�!#Z"h��"A!hDHYF�-"BB�iDDв$h���Y	Ah��D���HYh��Di�dH�Y	�""���DD,���$k!"�Z8pk!#YD����hi	BF�d�dkhH-	BD�Y��"""#H�"$D,�����B�"4"�H�!d$h����4D�!!d$i�d$DH��3�����ݬ���rgM߸��:nt~�+=��m�l�ٍJ31*m�g�ǣ//���v���޾}����y��?k:g(����;��:w����wbOӾ���<]������Ni�����6��~/g��:�x�����̞-��罽�OC��v�����˖���8o/_w=��88zf͛����^>�}��q�Ǔo߱��0o�Gn��X͛7��p�K5�7��ћ�ߚ����3��c���߭�p���o�3�73�o��{��֝���O�3���1�6h����__���$tg�����3==[�ݙ���vnMe���v�����8�ѝ_��a���{�t���GX����<vq��^�[vg9٧)-�ۮ���tpF���qra�f�3nZ36.1���pfr��n,�c���vur8�DR�D�>S��`����~s��d�#�s�ϭ�n��k�f���
$m�H�(��Q!�n!�j0lq��}���[��4���۷}ΞF�~�ȷ�u��ӷ~��އ\9�8p��v>��l[��_���^��N�6lܳ�n;\�����C���gn�M�{�S��~�G��#���f��q��o���#���������΍�e��yӽF��IǞ>}��%��_�z���lټ����v߷ߴO��q�����w�ݮ��}��8��ޮ�6�m�N�όٳ|߉�oיm����}�g��r���vc������ݛn�����Nܺ�3�M����l�vf�֊ȫ��*�z������~�lm�����}}��l݁�����v�yѹ5�p�~��6���73z��gLv�n7�M�1	�����4$=��C�?�6lٸ��o?g��_��}o��ۯ��f��gfo֛h�sս&�G��ɏi����O����{[��g�zNY3����[��o�=���oi�w7����ۏ~r��8o��S�z��w�3f͛��-���7��D�}_o����6n�{�{���������<���<�7�<[9����>���Ohv�4��i'����n�`�Υ\�1ͯC|����G/��g��w����l�Gs������tΞ�ܝ���r����1�6i�:���m��s�3�3ݞ{��M��7 �x6�.M�n�|=G��v�nӷ&=�ONޮ�tl���o����6��㞛	���[>��|��������Q��GV�{������&����N6���t��7��u�`�?ߕ�՜�#F��:�����w$S�	ja�