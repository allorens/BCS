BZh91AY&SY�J���߀`q���"� ����b?[�    {��*B�H*� DB�QQA
�T�JH)��)%U
IUQDD�BJ�Q!UE(�R��U
R(�
��/m"�mU@UB�"��H�X�DQ �ԂT��� ���J�I
*UI��*�*J��*�Q	S`85H��DJAU$�
QT���A*UJ*�
P�	PL*��M$B$�	(D*T�*����E!m�
��H���C� ;��Tm�FT�����d��ꩧ�wL�����eշw]�M(]wv��v���W;U�R�+��u��m���u�B�u����C��T)P���%)	_   �w��X�7DèA��S:��R�vϯr�B�*�v�Vka�K��ԒT�Kq8�lE9+����n�:e6�WP�)�U}礪�R�D��P�H�� ��J�*��cN�Jj���x���֔��7Gm���\v��k)C�UU'l�۴��Z֭��n�vQ"BCn����Mɫ��[iO�yPPU@�J%>ڸ  gw�*R���8M�%R���Y*�%.�*�V�v�t_w��W�U��gS���C���T�T��=�QT��5����|����U6�S��Oq��Ԏ�BQR�PR��($��  <��T�;q��iN�s!J���<o�@�4��t��J=y��RUv��+{�(�N�=�EA�Q�Ow{W�u�ev�u8�tԕE��uRJu����E"*B��>��RQ�  �� ԭ�p:jv��c�*R	�+�m�QP���J��n�u��n����wJ��ݳ[p�)�Wu*�,�s�R����uUU(��"D%%*<  8=�uݻk��p�t��Pq(Eíʔ��[�]v $WI��u*յ��n�f�7IwN�v��}�x
=;����EU[���(A)*D�*
T|   ���t2u��0�S��_OJ���r���+r�
tV�"���T���U�K�����C@}ޕ �AJJ%UT	I0  s�ą�8kt
�[��Ԗ�+]Ƶ�����TN�ܪW@@@n��.�]�J)Vr;] 6���TB��xIE��PT�TTX  ;��d=-���U7!��UW]��PK��n�UW5�Uv0��U�c@(��8zRAw%܀o�     ��R�A  &� E=�	)IPM4`F �i�� EO�C�US#P�  `S�A)JP�2`b4�h56�JU0�  C` ���ڑ&��6�z����&������=󼼽�����.�oz�/{�m��v�<�ǯU�Ͼ�{���
��]~j��A>�W�  �'����~~U?�D U���U��PW��J���"�?����x���W�C�?���fW�e&W�2��_������;e{a{e{a{`�G�@����L�����X^�^�^�^�^�^��^ؘ�^��^��^�^�^�^���2������=�������l/o� v��W�@�;`�P����P�P�G���������(��Q�D�� !��� !� !�*�� !�@�@�@�@�G��@�@� �@� � ���v��v�v�(v��L
=���"������(���E�P�"�l
�l��l�l�'l��l�l�� ��  �	�(�� ��
��"!� 	� 	� '�
�l��l �N�U	�P�P�P���|� ��� ����
� N��E��Ez`^�U��E� N��� v��m�W�W� �;eN��+����u�_l������P��=��l3	�+� v���l!�(v��l��!�0'l��W�+���^���W��l�+� v�����ǐ��i�N����~C�b����Op��+iF���B�Y�KQ1k&���Հ1R,���C��<z��j�J��w�ø#٠c�X�h �V@M˫�v�@��qjlFV�ڙ
�nʕu{�V���t6��Xn�#��㱦�k�@U�mJ�'A�3q*U����^���5���j�
����le��E�b״��!��jz�6�ZK�۵wB��&�����6e��$ IV�Z�,���šއ��n��K�JۓF�R��*o+��� ������\%C#9["�R���/7v��R�v��xt�3�Z�Rʷ���i�F�d���JUpE1ko�W0�z�Ф)^�1�]DA���M��(ܔ�104��<@�NP;��qܺ@2)M��Qx ��@~o(éZ�X�V]M�]�C2�Y�f�e�r�ʶ)�E�%H"[���l��S{J�7q��أ�v��2�`�m��jM
��/1D[�A�/t6@-c�p��Ε�Y7m��G���6^�	��ư*�j�J��A(�vf�*I��H�"�2DD���Xu!;)k�5��e��lj�������>�H��l=`�Nk�K4n���	tl6Hnk�զ�QK c�7rZf�j�?l �Š�=��jP� k�%�h�5Jn][���ViaM��
b�R0�r̬�ǆ�D�#L8��7��b��H����,�c�H��N�G���'���1YYa-�x���6V=�n�݌|Ӥ6;�4f�Qz/7�o *�q����Sm=�!��&���z[��� �U�a:q�v
u��hEmaYt�i* "��9{K������� �v��<�z�!��Z��2�b�h��pK� �{ji�P����{{�-��qU�"�y�V��Q�%:T� �Hu��&��ra����P��(�&��V�EfY�2��H**ka�b5	�e�#뢮!S1�[��ښ�묘Pt�"�Me@��m�����l=x�`�zA��׭���Mv�L�.�¬���@-��� 5�b5�|��j��<�Y��Hז�ۓm蘒�X� d���)�L#�
6��2�lRRd�nP�^�ׅ$��{D�%��X�.�!Y���a\W2e^A+X���Xݦ���EQ\��%a�,�V7�&�"�`彺*΃WVՓ�Q(�m�wo4ֺ*�Zɑ��j'���idA���B��B��̱(nb�4�*�(��5���6%m*;1=�Ŷ)��3�I���Lgo�;����Q��H�Z�Fܫ�y `{[#щ��&5�n�#�
�����%)*�.��-�Ҋ��vdy��������J�JV�x*�.��Ţ���J�8>�¬�.�7���SU{�]�+5V���7�TH�n�$�4f���ͣ�9�ED8-���a�`B	��IBTR�D�n��-�H}j�fh�����i�Z$Gv�,�0V5Z֖.�Z�ݪ�[-Yi"�U��e	�m�����O+@�r��I�.·z�����;�ƳZ����{EMaք�HѺÔ��NU�"�/3;�Y,L��cUl�OU	�T�#��yy�X ̛Gm�:�cR�ZpPM]eS.T'4��Y�W�n,���la3s��Y��7*lRmc��oE}�%�O,jV6,2�ͻ9�b�F�^鎦�%C !��F�|6��"��iZwjL�sP�b�"��ׁ��fӈ$U-Z������]�&]�,�N��'m�skvT�\����4F�z:;�b�Թ�M���Q�5��SQ����S/y3��k$���1��-�c5jj�۫�g��Em�`ۻ�h�"*��:oNJ�N;Je���9n^0m�T��nE0Qv [V�G��ĳbz��d��R���L�X�FXK6f�'ܖ��lH,;iL�+����[��Ƶ�&3��bG܆�/N��i�R�|�/v`_M��;N���,]"��T
*�j���f<��U��ڐ
b��r�U�6�!���╶�Ze<Ѵ��m;�o7�1����T���ǅvՁ4�)�*�u]Z�����6�qֶÄ�NJ2T�/4�ݡKE
���5��=Y�b�� Bj�'���=,b)�ufW��j{u� �u��Y�iR�m'��4��2,�(�o]�v�VXՙn�Z�I��뽚�	�b�t����J����չR��Jka����5d�����ˢ�*�>�Zi���K�1�6�q�ՠ1�@��#Uh�AD�m�۷F�Ů�f�ˀ�^;�n��g��	5h	���fF 4�&�Lc0�D�kHY�@]\��#�>N�vܽ9�i�m�N�ܤ����6���=�ۅ�T�Yn»M�y��$��#j]�Fl����kj�9ٷ�3���ږ�@P����\�ҵ�����Ӷ0*���f��j����p8 �-Xv�7V#�IsS&��찲CYO.�b��ӭ���6�h��Z��CL�͙�s�^2�G,:8�-'φ�lf�!�Yeg^a� wS��UbU$M����u�^X��:���x�QSU�7�(�KV�-��L��Zp̭@@awE��W1֥�����tM�hp�[�����aL.Xj-��ͳd�L�4��ۻ��ʅ���m�%	d����AV:Ӵ嵋d�n��{��
�'�a����ܲ�L��0�Wx�Y���Yt���p1IY��Q��ҍ��ҍ c�%� �s1*So�iEdk�N�ayL5`áf����MLӻ�7[�nU�����5��[�4�Z�ֈ�:T1\Pe��l\̥�&�{F�����&�iзW�*ӧ/)V�B4 e��Kb`�Ƭ��ѠsAS-�@���x�8��.fK�^ǈ�m�A���K�y�ہ�V~�L�~Y�hn�/鹲��P���q;:wc7���]6e<�pT���ݻ��MP��`�ܰ����w�clG��b�m-�/A��F��&�Th;`��ov�mݧ�U����E]��ɹ�L(Ѻ�N:F�1��k2�N��Xe��z��3���0N�f̭AT�S�L�i�r�yw�3^����&em�fݵ��Z6F��	1���T�Hpd���;�@��%4\7V�t&��EX�NEyM۬�*<�2�[�ڳ(���Q���*M@:��W���7W#�`e;I&n�v����ywB���L�zK%�FnZ��Ju�밆��x��d*I�����V�c��F��P���$�VIPR���"�3�ݵ���5�r�S&ʔ�DJ�R�ɸ�̺�^��^�&N����<܂�IZ�2bè�,U��6Y۳�X��A���It�nd���FK�ӷ�:a4�]
LLD���Z�e��L��X'��^ȩ�viIH�zQ-��� �T��h�2� �@f$Ψ����� r�h݌	�oU��	0�aa�4��d�q;7��N�ĵ'�wP���sVn����.��Ŗ��c]Ԍ�Y�ȁ�\lƮ���L�f��ܹ49R�w�1x�]�c��)n�43rD�n*4>�[X�Z�ۘ ɵ�l@���ҷ&��d�$�!�U�2�){���0Tfb��-1'�\$3Xw����8	�p�m8����0�V�ݦ�Qw��5�L)U����/�w���85Q���U����.6#��`�5�����l�B8������Mʺɉ%[��q+�P���J�JɛSn�ZlV7x�$�+"hK9���*���Ƚq��X�fd
�]G��{����`�m6�x��� 7jĖ���@)͑�Zr�^Ka!z)�Jw]���ճ�]��\�Ӏ�z�Vs$b���F���E������Uq�T�ùOh�Zi�Bn����1�j�Ic�V-k��'j�-c1���1�h0݉Oh�jF���U��L��Y6�;i�iц�e�:�C��j��H�1Ն�,;w�#W#+l7y�Křc�F�&]c3� Q��ww5�L��c���fe<sށ/�.�m��d�����*f���[����7D�'�]YCl��+ym���he1���L
�)�6f��A���7yn<�7K��]KS*[��Kx%a�Za:Sm�j!��܂ޡ��C�bo(�+�=�X�=VK�Z�J"��-�x�9MGn��[��u�mi[R5�D�&ږ��Y�l͓
]k�-��2�!n���ݷ�5YSH*U�v�Y����X�J���uoR�mZ��I�Z�R�y��)�a�泖le@�lYRޏ�������o�D�%%J�6�'��d����2ۂ���Ć
;�F�s\���hd-��l��eՉ70���,�lʰ3Z�[.T�2��B�8�Z��K6$��,��j慅: c�x�eF)\���+��M�'��r����a/3M͛w���!E���1�h�)C�ԃ̶-�"�!S��+�R�Wr4����vZx��vvd۲�e�(6����b.
_ r&t[{zf��V�2�m�+@V3iMwJĆ$���=��y`˵e�!�����r��T1ш��4���i�;h�7�f^���Gr�cYJ��/Q�A̭�����uE,Ǒjfѕ�e���T\�� L�VE&�c xe���Q�hT��ѕh�$v�e������2�{�1��K��
��������B��E�k �W��ⷛp\�4�M��*��ʈ�m���ߘ�.`��Cn 4d��	_R6��5�r��[20 $n�u�N}�j7jB��Эɨ����f�,���/r�a�,GR=�Յۘ$��1�p�Y5(JŅ�n,R<�,5P�MU�5:Q��b�G>B*�{#Xmc�ZBfe�����@1��SX�m0�\�/qj?'.XK^A�e���MR�����&U��Ū��B6L�B�n����u�UХe��J$�𼷡��f������0��P�c7�EӔt1�V�5�C��Co,Թ�ۊX�f�g�c+l�m�����ʀ���j1ؤ_��Ӓ8䁆VA{��7m6
��:`6P���vͽ�V��ܵ)m�ӥX�\W����A��m
�l�hX6��d=��T�l�<T�z�V��/2�/!�w
����š�cjD�l�Z��Ή�/p�cqc�vY�B�E�N�zd&�\`c��T�z4K݈��W��h��]��(�!�rjx�n�.ݛY�Ñ␍�ǳYt��"��ܫt��A[�pĮY	�,ȫl4JՄb{�T��Ɗ�i�H5�@�.@Y��RC�b�b՚�
�� R"�/Ej�Jֈ�;T�l�;u��/2�,f���-'kR8�ՙv�yx�*T���f��lr�5�r	��
�x6��A�k�ue�`�$��0�駑jF� �ebU�V��YZؒ����hXס��N���b�թf�D�Î��)VM�%���ʆ��Y2�K���0ˢ�H�	n�F
[D@ѕK$j�K�N	l��w�`�4cԭJ�tL�n´e����Y$��H�F[�14�F�CLZ�;�� �ֳt�;���)5��;�Ca��A��ӷ��U�a+"���y�V����I�d���p�Ȍ�����KPܻ6É�U6��  TPr3Q���E�+o+ƥܐ[a���t.�ё�ypn����Z��2Kj�
�mS��e�F1Mx�L Q�VsoV��R���T��tw�U�6Rɭ��e��(seL�+NH�)U�dR-���q�b�*^��	�svi��u��n^RF��$��+v�����������kXB�w���T�����"�ƥ�o# �xjS�4ҧZ���81@��o4Ll�DQ���1�۳m�W���J8�8�t�c<w��q�f�٬�z,n�yJ��e:e��)*�)Ce��];٘�7^�^�feiv��ˈ"QA���{�W�+,�C%�H�b�n$D�Ҩ���`�(�%w��(���,*��	Su�UZ��hI��kMAgujԵWz���U���fb���F'�ɳ�P�b7P���(E�
y�0����^���I`�mk"T-�@��A��B�D����TЦڢJS���Gw+K�1���2!O4ķ�Q(�����Y�]y(u-ߥ�k^�h���hc;3(�$EX6m�*W�nZ�R���-ڼ�I��PUnD�B�Bq;sn�- �N��x�����Q�Yٱf<X�$Kչh��c �)eG��5�)���L�[��Ӭ����n�M	�B,KŃ�4�H�sZ[wkS6D��8����2l���U�ѥ	(���{�[;"K)�E}���������wkE��Ar5��0��*��h� ��l�9`ѳg��J(弻�^��ԝR0fQYb��R�2�́Ȫ�)`JIj�l6����x�镑h���r�W��Ա�Q%Ab5��y��;�\r���Jەr����↱�GeD�E���c�ChR�Т�.��KNY�h�x���"� �/�&}�%����㴾����,j,�e(5+/�i�M�3K[ 3pFԬ���ʕ�\�E�ot��vT���ҕ]$ub"GJ���b�=��|�q��C3 ����)�Ɂ�K*#Gq�����ˬ�B�e�ַ�u��Z��<]�Vԕ�*���FAzq�oa���;�Ϋ|�Z�����@�Ƹzf9�me�ӕt	�?.*���$Vr����Nbf����,�ܣᆸ��E|���B�� al`߬P�UK.�� �˗�c��J�;ő�k�Eɽ/hڧP�~0�7m�S��4�=��W�H�1R�V�݊v���RξDVܲ�KJ1h�V�k����A��`WB��J��D]]M�4��k+Gs$zm�U��c����ٴ�5���{  }*��E�]Ыh�w%�e�u�Ѓ�X�=���?�<?=��f}��?��~K�^����s&OI�.��7����[бo��&�PU6p=Y]:1�j�qf�+i�2��a�*� J���}t�	��Uu�,�����6 #pW<l�=��j�.�{���|qfL5��c&1iV��0r�]������U���	xu
�*d��������߸d�c<f*m�n�̼�s�A#>��G�n8��4�Ҵf'����sm͸�%v�_۽3�L���s�	wn7���4U�`�,p���#~�f*��xZ���J;�s.ԥa7��Ԝ��mr3k����`����s��Б���Jmбl����Yo��`��t;���5��V9i����p��)�)v��8XgjG(Q�����KɈ��X�%Np�o��+8�Qחܖ�jX�2��d�Wk��'n2)�,;�Ր�\�cY�����|,[��ԸJ��}�۠���IGWq��[�}�r��`�P5�B�%WcG K�PZ��� w�5�v��j��lȻ�X)� �V�4�С�Of��R���e����e�Wu�|�&�ܚ�2�nn�bY�U��3��\4֮4v΁N��ϱG[}�jr,��H^�#m�H���>��B|�uZե�ޓgq�bBG�W$u�^̓OS/N�{9�^8,�5�����6w`�mh�Il1ǎ����:�5�Wu��$W}M- %lb6#/�u��S$�X��:� �u�e����ص]C5їh��W�e�K\$��YBKY��8�2�%V��wM�؆�=<+��WRW�G_"��itě���6T=@Ԡ�_m8�D;XN�Z}�c� ���N��WH\��w-Me���:i��:�����9��h0�����lG�a<��<�3:V�įq���0�g)*����8����=��U3ݧ��W-GFu�qJ�o5
ʹ�K��6�32�V�%�!���r���N06Ò�-  g^+��{2uFk{ھ*�J��4c;\�ə���Ⱥ�u��{]&���6N+��Kyayn,zݶ.��j�]�v�H�̕����_UiP0��ԬnT��#�6���})bY,����8w��2��\�%VP��A���f�o1 �\��'�t�{LsU����b��,�qx.�Q�D�ooWhu�XR�X�[v�Íi��N�h1�QO�=��!5�G 
�*�v�J5��ݫKh��x�H�n��x�]�����"-��Yo���S��½wpԡ[�q��������Ec�*���"�R�9���>�ł�^�]�)S�Z5��9�#�h����K}pq�k2��E�kj���Z
�N��R���2�6�Q��>(M��Ix7�CN�ݸw���^��7�؍w���CW����ꬋ'�R�Ono^!>��`h�)vY��;�Zr�\�oR}�D4�'9�1O;��M���Vf�٬���3��2��r�$���Y�57�k�ɣ4��m�۩�N�]�JaP8�dލ�v��"�]�CI��z���iN4�M��l��q�qǧ�r��a�Yjr0r�7R�,�s(n��T�Z�\a�V��	ڀ�1n撮`+����v�ns����lҔ
}�Ck��4��dS27��obۇ6]���Eb*�d�JO�^��7�cN'OL�Ѭ��4��'���F9w���[��g��Ө�W��&t�A�����1�� �V�_NV�)�(WE(csE�<VspX���VY���mLc6�#ջ�!`3�>Z[K��۝�@���nX�p_I��t�{pB�q�V�u�8��f���l@�7������t�"�}n�1�s��<�n�Ŧ����!&��]����cO�JC��I���b�z�vJ�j+��%�d����هgR�lW-D�d��*����:}���@����bs3�
�Q�o�����8:ʤ�$���֫�;ǧ��^�BPa�y��-��vT|��#�^�;�emL�w��yT,�;c��%�n��َ_@�Se����Ą��=�
���to�c�PA�
��v4��+���6m��IQ9P9�v���ixT�ͫc���;9����a1;�2�u��*ֺ<779,w˒�N�-I{�Vs�6\;�&2���@�[��O�U��X�ۣ����[��'»)λ��=N�ӥwrN��4��̝�'\mcYV5dC��é�0s����s;����TI�J��IY�J�ۚ�����4�����<��k��o�,�3�*Kˮ �6��Y�(��_;{[-e�,˜�4Ԛ���a�n�J�$��ۼ�b�Q�=���C��tA��or�v��Z�}�bQ�ة�#U�|;�n���9��B�X{t�t�$����MJ0��R�..�osX��c�UGˀ�]�3 ��BS:��K��;m����qB�p�p�>��J�ûտ�e�eH���چ��z�z$s7��Lp��$�LVf�9�rYy%���|hgN\_Qdp��#��6MՐj>��N]�S�]juwʖ�^VN�Sy��(*u�M>P��zz�c��?�pm�<�{F��Xqڤ����9�.���h=UsYe�Ygi]���k�ݙE��ep��dyK;��-�-yPX+T��S
�wmgL�X�Gq����v��h����y���M񺮎k���jct�n�B�0�\��T�T{L��wtu�q��Щ=���(Y�j�\9�nsQ��&�u��O\�V�:�N��
9i�W�WgZ�&��F�'	t�S��҄vF�`�T�v\�*��I��H�o)��x���TS���zMl���:���'`ޗSX��R9;v�N֎D�Ce�vhJ�Uƴ�E�r
.":��V��;D�*u�j�Ry�����.��)�EȤu�XT�m�s�3��R��'Esb�����M���zL`����*��_q�Y��%K��1���,A9S�{G\�J�i��kM��;��ƌ�A]'\�Ͼ��+�[���w]�)FA�*�F��\���!�9�V$�tA�[����iŐuXhډD���,׳���m�b���κ h�k����@��8����X��Xx�u�F;��#[�Q�X]no���=�0g�+�V�o"*�Kae=~�#���C���RQ۫�b�q�
�Xc���;!ߓ��ʓ�����(���-c3x�*��w!w�^b=7�ڼip���
B� �ˆ�U��E�u�RYX�L�K����4�)�aԠ9+_7�,EA�4J�TP�;�.��5evݱ�P��N3 �Y�M����,��k2	Y(p���gK]	e�˶3  \i�� ���-���U������얮���ܨ��B��;�����ǺE�ݤ��ڪX�v&�������� �����؏�R:�c�����;�A��<"�<|MeG�6��^s�D(ӡ��}g��[�t�<y��j�����Q���u��A��MG��Nn8%��5��V󓱎�[�v[to,�(boiꋂ����4�Q��ͱ�����7����12���v�� 36<P��\�!�$���O��X�R�R7k��W�z6��,9��\f�f����>;�f>l<��!�Y���Q���N��|�qhR\��F]Ʋi�����|J�F̓0��Op��N���������Eaq���M�v������'��ݽ���o/�Ҿ5�~Tݨr]˱�0�>Â-��ɱU�-�w�v;�z��5a�*�Ro[���p�My�&�w��P��_�/x'yRZo~���lݷ���*��f�����M�y�8��U�`T_rնAO����+m[�{WlĂӈ��A�w�����d�Vy[ƛ���mubZ�����+h�Ү\��7�l�rc�x۰�]CÆ�����N����}6�!.���X����̺�bu�.A�T�4qX����U����Ct�K�7]��́�2��ڮ�u�rs3�ƬjI�Ъ�����Rq��9)ud쾴�*
de�I5����`�uǷ�p,���)�;�d���O�`}��4Db����oy�(�gYO8ᦪ�*ț��GZ>��Z�͛�h����Kp�@�R|~V��rfV��_�WZ�L5���(տ��VZ �ε�
�a��,b��M����O����3*�U`v�*f���q�wt�K�+�A�! �g,�P�J��ק�XFo��h��G
ǽ�8 ߰�"�D��`��6r�b
��qǁm�j�J ��33�Zq,�RW�#vk���ꛝܹw'F��6J;s�H;��#Q��wP*�M�ѥ'�����F�K��\�X�Ɛ��͇�BW*�\��=,�y�\�Gk�=�Θ��
�����KD�OX����OKVv��ٲ�ڦ?۪0�w����9׃c��pk�$��Di]�A˚�2�J�+b��_%�g:��\��hg��u��I�ۨ���@�w,R����Z/�ѡ�^��e���;of��VVj�r�'�\�?*ҌE>�Q���*�;�偨�`����iм7�q�OhG+>x6^j�gl�euD�ul�*��94�51bJ��%�B�ц";�}�=tU�����M�N�κadgW"�]04�7]Ӄw���4J�֩wܱ����52�v�;� �Ħ���L�}�J2.�̼Gr� ��Q���n.�2U=��s6ɡˈ�V���.+�ujJՕ�*�lݼ��O��{�&Q�}����wi��D��9�����I�; �u�!]JJ�Q��/�I�z{-��b�:i���H/r�z�NݸbU ��;yɋ*�D��F���t��p*fa�k����[�j�슳�� p4�H�y]nֹ���ʵ��ݭ�y�Eem<i���Ǫ��t���9sa��;����C��,;R��<��yݭX�۶ՠt�*t�����^���S;@U����dm�Ԩ������s�[β�w����b���[Ŕ�&ͧ�-gG����ہU��\�\�Љ���π�A.��a��[�|q��m؟�P�G����\p�.��2�W����Q�w�6m�İ�'��d���9Q���Z5�~�3zT��n��
�\����\�-7z�"�
o��j.��f��7Ep�E\:bǝȤ�*p������n�gq��<'N��`��l��.�����`�$�ؓ���qe����v��6�r��X4��Xz��`=1�U�&r�v�<8��rM��W�T�r�*qO*Wq��-�ۺ�)+|T�8e��5�8.��Z:�.#n�Y���i���*�A�7���wn�����B�&z�"���2��j�Y7�>��`����O-�>Q�p����E��S�uB.�|ؕ0w\BN9/��r��4#ˬ�}���\�4�ɽX��MC�Ӻ�i��Rf��x��s�7���i�yY�1�ڛ�+:��ڵ37&�ۉ1�7�y�md�"[�{�W�1f�k��Y��2^ig����e����.���i"u��kh����&:��&5����5�����C(u��^�� ��R�������o���t��������|��Y���t��ȫWv˸�����.-�6�gb%�K�����-�����gH�C�N>%��KP��~ XV� u8��)��]�l��N ���OU�h޸I��N��7t�p�����`����ŧ�ޗ�.�6�vg3Mv�����8g7E��.���n>�T� �i�X����m�[������`cߠ�3�(�_zɻN�.�Y�p����RH8��2hy9}���P�s�N���B�{G�<�Z쩣��U>��_v���b�f�G�Z;�;�wc�[T�s�|���a嫷Î��yQGN��TRι�U�p#�^�]��Ќ�ȹ�F��
7n��N��;���O9��G�� ��v�vWV˛5PW��R^��B�j�\2=�M:Z�fnvP��M��n�i�V��䳺�M��m�qv�sT���>6۔�5}Aoiy�띙�Ґ}#��jU�w9���%X�=���F\� �#�T\hҡ �x01c��(����zy�J�6_=�h�J_[̥뭪R[LF�AP����銹,�.Y�BL�՝Cs���El��t�Kf�w�vvK��K����i��f����R�9�b����u	������,����s2�׃�\���V�0�����ʸ1q�JX�: YW�:�/bp(��'�߀v��m�&��[�Xг�v1�Pڋ,e�U�H\rqH�2ͫZe\�����q�8�[n��a�;�Ee��3���v�I��D�D��T�z�u�#9B�X0���宖���U*uev��7g+I#��RR�M{�KX�	+�ɇQ9���Xh�'O�:��Ժ�����Kʕ�k�%)	y�A�8p�'y�������o�Ww��z7�wP��r�:�+��Ɛ��٦ԉ��Z쇻i9�����B[�\�R��OH��]���p�ۦh)ڑ\ȓz���E���{"���\��`�3�����$�M�������ͼ�l�,��0ni�}��O'Wm����v�r-��)me:.�-�]v�a!wZ������"8䉞q�:�n�WW#51P^�������X�9[���M܂n��n���B�W@{�h�r��)��-��{�8di�8���.���]w��U���՝��`�e�N��JX� �8���f�V6n^�Y��u���ni���@���QR �.�
��� �i�tC���a��d&(Q�S�Y�C�h����e%D��D��@$]rI&}|�aEYt3�QF�0�D�`R��P��')��-�,��@��L��A�KL�舍9���5+F|��G�+[�#F�1|��4:���B�:)P�E�SYmQg]sk�E������PA�}#���"���(�����/�z��_���}<r>��]�q�0^W�e���+_c=�Gt�d<���l��X�.�%ʄ[��7Ff�Wh9���Z���=f���]Z���/Y�U�ibBr�:�v�˱�Ix�u�Ąb�5o+s&U�M�[8��M��=;�H���%�U��凲�Cs��5bwK]\�p�/��I��n���ʼ����3��ɍe
)�V�q�J��*T�Ӗ��z	@���u�r`���:_ ����Õ�X �጗N&�o�a.�4t���fʩ�K�&$(�0U�BpT��m6�][���.Ӻ�<r�۽ sA�֝�*q��ib��u�ը':Y���W�|����v��oF�Su-�.j7�{�5q����R���s��6%������=����Hz����b�ĠU�^��|F�^h���Q���c��pw͜�Ћ�i|�BF����Mgk=�1>޲�v��[Y�������gq�8�g����Szsg�RJ[w�]w�KR��6PF#w�CK�HunĖD�+-b�d%Kkt��q�d-��E��q�VL ?�[7����hgmT��;h{+�Qy��ݥNVb�5��L',x��m�ъ��
a�2����D���|�;5-yTӏ��{��m�SI���:@��f]�e�[�gS�ۡ8,�j�E�)�'�@T�o�7��]�}��b��5���.ue7Ɏ�-=�̓Ad����ok�PV�G뼟If�2i�4j��ɫ���tJzM��*5�O�u��X��g�f�����}-���K�K�ޛ�Θ�W�����3o~<�u�5��Xթ<�`�5��hp_v�U���ʵHqŕ|�v^�|�ɗ�v�jٕ�#�h�޵B�e>:Q��rU�R�q$�Yb��4���ǈݭQ[v��� mJ���N������+(R�O7�������q��q|l��)P.����#���R;���%�Kꛌ��@CS���`X#Nӌ˘��=]g2�-����|���]ij�*�$�Q�]��4�
4	W���(�s�\��]t���ug�M��Y�l�N�
%�9 ����*��s���Eq�)�-;�L�q3b�;�����m���]�:����crȬ ��̓��].�#�s�^�alt�&�mX�49���
����Syu����/+�9��n�r�ˣ�m�|�0r�U��]��h�*�VX��0�g�wS	�RXJ�RE�,�w�6���k5%����d����M�71�4��k��3�:YAa�&N��4Qa�5wA���(EJ+4Nܖ�����TN��w�s�+�5WО�fȣ��;*9r7����k�X�C��
�a��2��V즷��O�}�+�|9uM��o"и��U�����R@޽ig:��mtk�=&e���yv9�)W;�R����#�	Sq��P�^�[�K�g;X�v.�s^�!� Mwimv�8�qT�V"�n|Z}��bg��cu�D	\]gT	��xƶ��|^�p�C1�'��9ZV��kvb�6G3k,���=QZs�7v� �g3��]����]RqG-v���v�Q7�q����{[��SGkCqJ	���޺wG�3dO�4CZQc���;��ʮ��iŮ��"��@3j���׹�2��7�u��k�N�A�1u� �+m����Y@��b������sTfT�֓U�J����0%�J���#u�rn<}F�M���ֵ���Zs{YY]��խz�\ǀ+�|��Y�\_ә�:!ßTٶn��*�L�wx2�&�D�h�@͌���tY�,�H:3��d,�Wl���]��z魷��$4��^��p�+(�����x����8KWOE'Y�Gt=Ӵ� �J�[�Y�ƶ5��qe�"��&S��8(��(ѥM�ߦ����N�]�X�ȟm��"\x�"�6�ϫ�&rVn��n�v����e���'6�㠲��.�����(>�e��V�̫��r׃N��]n���A�3z�^��t�oP����޵�l���L4��l(d"��p���pr�(���ͳ~[y�]�0 ���.O�e�{1��JVh�{>l��,��֨����m^��z�;&9��m@�gJ���KwV�h�]��ޤ:�^$�ݥƪT۽�R*�06x��ú�}��L#,ds��/!��Ѻ���mh����@�����ͣ��*�n��K�:�T�޴�,�qT��dL�0�ɿu�M&�V����P` 8Ѹ_7�����̢*ޘ��6�J��J��S+u�z��bu�A�����ɗ����1A @���z���y��Ӭo�eU���G��^`"��{t��}�a�q.f����T�NJ�ͭc ��GfiB����鑝nr�JP��9uh��!������r�.���=U��n�_ F�YDB4Ê�F-��^X�y\�M���6���]�}1�p��i�ڕ���y�B��
T8�x3n���o��9ic��r����9�'^�����_}�Ma<��)cG)��S��P��G�w��r��z�������Gˌnl��3��)]w*��t"?D���eu\��N<�sI�
���=�f��K�Y"�ܜ��R稜:�,�xv5��r���\pj��R=}>.�j�5�|�]uhV��>;q֪��++u�2�{�C�%�J�o���s&jG�����r�7tZ�L�4P��
�'3IX=lS��=�%4E���kC���^�ŏ������;������k�f�`�ok{^�X������Z6e�V���V�#M�d�92Xφ]izR��<W�1]nK�_<ܪ����ǲ�H����%Q�`V
���v®<6
X^k����n�,m B��kCT�6}6`Tu�{��c��,%Ճ��C4�v���r��/�u.7�AN(ۻ��]�{����Zs#%;l�ϭ�B��J-V����:�9J�F��=j��	:�Mkz��ٵ�}uu��#nW(moV�Ϫ�.Ծ!�o��G1�Q�Xu�ST��%�zjek�u�w�Ś�^��z��
X�/��Emg[�S4t��F�&�yXЊ��Pj��N� � ��L��r������e��+�p��u��I��j�W#wg�y(�X�v�d�/P�}��9EI�W�㹍#��G}��27��VX�,�꒴,E���5yi�
����\������72�`Se(�3Ù�'�f[�+��%zU�s(X�������μ��:��fM��CGN:	#p��j�0sKΕ���\FZ�T�Mf��:��b�����B> T�$%pC^e���Q���00*��
dYg�a�\ķ�om\�n��yS��tE�]��b�k�[V��R���'t����t������m�r�
OT���5W[|0q1�VVV:�.�rN�Q�
[�!��8 �Ժ�d�غ�v�/����F+V�#Z��c�NY�k�,�)����+n�m��y\ӭ{w�(܎Gݐ��ˆ���v���C�ѫԲV���4���$
��%9u8�|(P:�e⤹�y����@�whwR+������b�b^y5V�ޱy���X�hH4�4���V�'Ԧm���W��5`�������M�W�8IR��IK��܋i��1+�-�w�88�:�2��oQXz˳( ��K���k�Y�{�3E4C<쳌�(>qa�[]Բ��m�EZ�NcD`a[��ƚ�*
��3fBr�Ӌ[[Z4v���KP7@ǵ����u��3h�ؘP�]�A���Qt�7+�m�:�ޔi�����y�wAf��9t
�?��0�1������f�tvMe7O� �O35dȭ1��h�ʞq�����k��d��U6n.�ճE?��F���G��k-0�i��*	:($��g[��<�tVv,��{;/�����RU����u�(��8<?s���2�"v�4I�X덅{X���e�g�*�t�mbu�.$7K��1�%Z�bD���ɑ�,���8��*�܌�}��	yǕ���lv�W��D�wo9)���h_;��ͥ�]�2R����Cm���kF[�)n�VWnv�)����u�F��
PN(�y��F��ګ%�-�=��P'��3��9gw��͑�ń�'�u]q�1Э�n5ƦNE�MQn�	���;��D�mc�L�u�y�X1987zVZ쨬Tn�ʴ���[�U�yXܥ�r���'rA4op�Ʋ���.Jt��2V �!`Tȫ�y@���Υ5��`u>�g�j����Q�lJ�ac��XY��J,�CLW�h�N��񙜾�r�"�8�dFY��t`��7�f�^J�o��
(���Z������srwgSwu^�͠�k{��RӍ KX��L�֓#4���V��lb��V���Ή���4w��]��\��W���5��I�Pޛq�j,3v�<h��!j��c{`�_#�sVxa�}+P'�wE{zٷ��Dg����mu���K��?rW�#|�To[�S)vִ�4��<���z�@��l�����\�K�]�I�N��,`q�+�냢��sTy�1o0��� �<ô�b\)Qcx�[\�9��k 4��Ep�����qz�՛�]�N�}��qcѕo�Ǡ�f�4_!Q��aawe�ҟ^M�u��|2�_J��Xx�1n#m�󭩍��o�-p�!�]�'������Y�G(�+j�POkNg|TJ��+k��R���f����)���*ޗ�g��Lb����Xy�֍Q��܅���r\�Ga-^n�k25��ią���y;�9f��`��s{�	�X��>���Ą+ ۴Ͱ3X��;���yu�wD
���Gi�p9+/q�X�Pe��R�諚h�Dv�y�/�v�&c8��n���.�x.�$Z��Z��
oh={������R��Amյ5��}g5��xԪ;Iȷ69�}�vs����
nu�.�Ȃ��R���{�<�^�ڍ�t���uc%I�k�z:�.�k�
c�:)g�I��ڝӢw�*݇n�Qav��A���E{���9uۖ4�]�u�Ek���+Sr���/g�����d�6��Zƹ(;`W���N��m�8ʺ��]+v�]��TOA��PE��j�Ϥ����n-N�voe;�Ck���i��T]�mM⺬ip��h�R\Uj'[�jipt�:+�f GD�@�>۰�L<6�]��QTGU�M��������L�X�F�QgR}{��̊r���[�n>nҐC���6ᔐ�	[��֙ne٬�z��s�_n���n�a�܂�ݙK��e����Zb�	z�/Z�Ԋ�� ��T��1D�P��=�,�H�K��_:�����O^�jWc� �a瑭=Gt'L�䆎���Vv>�4Te��aq����gU\���F�^Zõ��uI��gG:�%C.e�yV=�E�;��Xz>*���T����{eٶ�9�P��� &� N���.U�D�h��pR�ڮ��4�3u�-�\'O�Ȳ�G|�:��}��<�1�Y�0]��BgR)��4��{��;(��;����yĪc��U��*�t��lu�,���b�rh��d�\\���Q��K`�ާʂӭ\�������[g;(���R3	�[����vMXc��f���}N:6�J�^�)i��Zی�����B볃��hrgc�5qd=���T����ݿx�B*Ą�hk�ИU���t�@��wui]7��f��H\�y'�8���g�^���m]c�l�F���wn�+\S}���ḪV�VP��hgCk�l�.�8�,gIzC:�\���?D���S�M�T�����H��*վ�U�d6jse�̛�U�'U;�� ��e뫎I����}��6٭<%���4�g�*���wQì��� t��.�J�X+������q�:�m�ݻ�U�7��u>��7"��oh]ٮ�}��S+f�eAN�����20�{u��e����C��Q˵xV�+��Z�L}�Á@��9�Es�YW_cxŧ6ط:ld�ݟ_,�i����w�p�i��^��A����xK�ώ�狸�0�TjJ2�G(]�u%��p�D�!'�Se,����fY�w��FZ���}X�����L�B�w���1�~Fmu;��{PNs;�HFk��t:-�z������Ė>�Q�H�
W3SnP"c��jE�.R��1����<iTU�&_:5SN뜛Q5��汣cn�r���EszC՜�v��9���Jed��|�	WL�l�^���bB�Uz cz��T[
��s�}��,��o'+���C%���w7�0�7���.�K��b1:dJ��N
z�Δ2���r���y�<��C2�ġ[��t^�gD�Ŗ&`hݔ�řq^�o���Q����f�E�(R<�Nn>�㶒U�[,�H;6��ӧkS�=j�zrh_�S,��)�u�Ŏ^^���d��Kڝi;Zr;�@������usfN���9Jł��E��`YA�hgx�m�xP*��Rz�g+!�y���F�"�u��<�� �8ۢ{�*��f�s6=/��)��WWv�|�ͺ=��]0��T9�L[W�:VҵD��'��p��ו̝��wX/����9]A�vs�K����B��;YYEP�L�話����<�:U�*p|y�&��Gm�6mr�/)���Z:U�l��p�F����e� 	L��Մ�nK�ʦ�mJX5���f�ݹ�Y����諥��X{euKWͥ�d躣i֊���Ji࿐�Y��y�h8��!E�Jl��
ݹ��Jj��q	UX��ѝ�ȉ�3�VU,���~������� ����������������_������?g�������������=�����ׯ9v�\�!P��G�t�N���R�'k���bɪ)��+��w�)�*�i�]}����Ȭ|�ueb�v�X9tHYZk�iQ�P����Y���Ԕe�_*G�p��9��Y)ڜb������KL T���ҥ{���JS�t��E���@����r���ϭ������y�Vc�vͥ��V#�t�%m�F�w���u�x.%`͂F��ZwP�E�.������P:c��۠�|�!�
�h�)�9�vE[��w�i ����tɥX�U����׺�5��&�ʑ���V)-��bΐ��.p؇ 欳]{�.�V��Į��:h̗V�\�@�w��sCv�IRJ�\C��X��Zs��L�yWjn��Ԉ�j#[+PSZ�X�oC��:��ͼ1�|#](��lo:e��r�m؝���Nn��Hv�do@ b�2����N1����++r��ιy�u���8�,X{/Mur7r�qc�T����M5x��eL�Ca�׵��:�z�$�f�3��ۡtx����T�*䔀[Z�[`�T1ev���|ۭ��âu5V���r)5W$�u��;YF�p��@�K7m�G.�7K�L��;�+.��A�Ĥ�z�a�h*Pͨ��T]b����r��r��&��*rK�w�2��o9Z�ʿ��ؾ���:-�R�h&�e d3I� ��E˨���Q��U�"���<E�Z4D��ąkE!M�vƨ6��C�ml��i&!�t�����l�B���j �h
i�))�))h�4� (���ZkJ�B���h.g��E"QA�5@�@i�JRI�*�%�"����Ji(H�A��(tWJ�h���F�h�)�T���"(
�
����)�����9�iR"�&�����j�Ӧ�i����%�"cD�-QE(SlQ�h��h(\���y���	��<���q�6fq�ܙ��H�X�W�\�,\���0o]����^s�s��zw��s�4Azs_Bu|���}M�)���2����yԭ�X
��U�_?��C��p<}f�����{���=U��>���{6������v���m�7O�ﵨ���J���=_�j^6|�CFGv�� �z�k���w��>L߇ˎ�]�'v�c׷D{h5�4�Ϡ����0�7ku����������Cq+E����O��[TU�w�O���3��gK��먮��A����bg{�V����zE^�{��vi
�5@�T{�׷>��w��]�G������o��i��&k��1�����6�q���\׶;(9]F����-(��3-�C�,��	������9ŏq�L��e���ص+�����/��`W��m�>���L���S��r~���~'t�9�"[�{E���L�F�z-�a�uV�׻�f? �<p����'}�����J�����8�nO�љ��Rzz�7x�E�aN�K��~����Z��ǰ��ta�<*Z��A�ͽ[�y��n�&�2�OR�����gW@x���B�N]޷בm����J�g����u%]&��^���!n���t���n��g��[ڟN��\�ʷ���*.��W��}Jd�yRc5�swF�� Џ��.���o�뭦)�s����9�=�/�W��]_���)���_W����-�{l�s��!�c��5g��)z���kr��Z���@��3=	��ןi����@�kM��,v�[ʰ��χ���i��t���֏Dټ����ș�n�D�<F�M��L�z�����u,\DZ��G�g�:{��G�6j�o�a����{�\x����E���׷q��jw�ZC��!6�]�ِ���6%�H�}��F�Ƅ#AˑM�~�����]�y+�2OkA�R���=��g�m� ��*_�Y�b�=v�{�2kk�&�v�3�$w[�W��l���o����l�^��yz_�hq�ہ�zz�9��'{���g.w{VB)�����k��Aw�R�oSO���}k+ױr!my���ǭ�/t$h� ����B� �������[ڛ@��)�1�7�J'j|@i,����1�侥�:�F5�|�)i9��/�!�}V����F>�x�K닶��W^J�R�\��hԡ������[Չ�m�"P��x83e��{���V����^S~���ng��ĽX���t7���h�_˫W��}�H_e�}��xO9]�fO?,��}8��\p��� �ҫ՝ �����nߛ���9��ޛ�\w�>�c8��vx�픴����b�X��ݣ�ؖ��7�V�����3im�fd��F�[�����ft���{�o��\���T)����_EҞ
�V |m��@�'��c�daݺ��q�'F��;�N��讐�r��f���.N��9���3Օމy��}�θ�Ώ+�{j��6�W���ZN��ao�TOm���"��Z���R%e��Mx�8׊C�vz�* <�-�Nc���^߼��P��z��g�j���Nu���)��(T�3M�nv����k2�`h�ϒ��b�Zh�v�~�UY@J��7)y!������ykQ��Oָ@S���Bi����#��PW;���'����o��|����TX�1�|�=��e݅�2��$��ǎ�ޙ�h��������=Ɯ]��伸|��&����إ��Ջ�nq �T�i@���g���f��j��`��[��pR��ʭ�{�*�X��ft�����������~��;�V���{3����O��;�Y��[�j���_ZY��x> Uwm��3ŵ�����U�y�/eoԵ�&r=��+��Wy��q���*�+�4�z{ʒ2p'�F���+>=E�g:��~�߷�n�����[��NC|}b��SVU�w�\�Pc�^�oևW����)?t�:w]�nV�Y�xP�p�=깞��ܸ�6���1�kς�xM-�M>������al��5��PZ�,���PǛ��k7e�B�c�������ַ�3��s�my��g�x#I�t�3Gh�M��c��g�Q݋t>�E��k�y~^ɻ��%��Gxd��(�W{�r��yHg�����X�]���� k�Oq�j��1= ��bĝ-�l�"#0�&���v���^����ս�_#�굹
�z�Br��5�-���}'Ly+J;׶h��E�ٕ�bu����ڎ�88�b�q��$.ni�hҔ�(@��d\�ͮ�@Em�(P6�7z������X�e�	�H���6΁�UZ`5�t��Յ o�t�b��9�1��]��B��|Q��|�CN������qZ���]��F��{�z��^U�@�{՛��)��Wp�k�+�Y�׮r�$9n�:y�Qj�{M��;N�k�C6��Vd2�kͦ8�	�v0�fߨR�]ї�7�.�s�C��}]�7ê_�Hn�q{R����V��9FsH�tR�Q龍؞���ɶ��]�{ާ�SՖ���@���zЉEɌ߻ޏ�׳������x��V�W���c��\˨^�/ 3ǘ��ƅ��}3��-Q�[6r�a��6��v����Y��� �}�o�����y�r�;�U���޴�=W�����;�{������-�jX�;�|��}����}J��u�����J���A񵵞�ߗP�:[�-�HP�@�/��ǘ�p����{��z�7�߭g[_Q"װU���������ka-.\����p�E���bJy�r▋��<j��|)_jT����n��	My��M��"��:Ƞ�꠬���~�|�;b��+�1�8�ٔ+x���%�y�o^��܂�ܜ%Cp����d�q̦���1M�O�кtB]l	�7)�ً2�$`��f�.��C0�St� ��wg�M�An����?s=��_�Sjh�>6yv���T�Y2�/����:h1�<�p�>p�f��p[;�c��	��uWw����%#]��1�2�Uv�8�A;�,9�-.皟�wj�tť���Oeo�C���K|�״ݓ��?u��7�����eG��1���ʱ�����5n'8�+\[�-}��%��b�R}��{۶W(f?��^I_>�L_�>v�ys��n�V�z���m�l͞�7a��[x�	�u�͐��DI�v��N� �ʪ���m�#���$O=�3�]�5�Ô������<Ǟ���0�]��hn�g�9oS��{�;��udw��Oz�o����{{%�f��8ř���y|�ⰽk\�N��N�B����M�UT�ܣ����מ��}���9՚����8��ұ��gr�B6o9�8�"I+>rk�#/����ެᄍLT�T�'�V���e�7[Q�Ǽ�NKu�ج�U��M���5���g�� 7�����
����Ձ�,���^�~�`_n@V�9���1k�>|k­>���*7�W��`�~T ���^Y��T��O����&��vz*�{� ��6ϼ��"N��W�L�s��8g����$�����_�>&���<��5,�:Z��-}D7=n�=j{}P�g��
����n��d���9��y�T��7A����}|���z�7��uB���0V���m�|Xq��/'2�Ƕ}D�ֳ����K�8��{fDs�:s��Gڟ��늋,�j�\����[�LF"*ZƵ��D
To6�Z'rvX>j���+�&�zv	{eN�4��Ϳs�߾.�`���[��{FUz#� b�ھ>�i?uQ�پ�h1v�9^\�i��x�Oru=��^����`����_������$�� �H\�N����짊p�f�q���͆#la��y�[��~tu�A�S�"�8�ǙȮ�D-XŽA��fNU�����+PՕ����3��.�����R^�3¶�6]>�Y�NJ�R�0�u���k�w5�m�����n�u-�����2��V��,��rK��a��l�j)�$�9l�
{K�%�d�TrZ�T��;�L�:�_��{r�{IL��6�2j�a�d/.�@c�A�d������t{΀�u��^�Sj�����e.q�T�p]{:���sϲ�#���9�͛���N�M�6��F��{�e%�9�� ]&T�7r,|�M�EvP���:���c>0��CWR"ɘ��l��06N�Lc��U��E1�:5?��X���g�sP��W���K����o�3/5�����i	�\Ҭ�Ɵk=��-�5be�*��_�>K��{��ή�;I��ɋ�L�5��4��f�ygxT�lw��8�߳&���{Ւ�5�՚Ѡ���؎��Nh�{��[��~��su�n߳�=����r�K�W��q8,NW���waK@��m��J�<!v{���A��L�:a�,�{�k:����<-Wʒ��9Y��%i�;�QӧX�x�uo����<��t�&z���]_�'���b#�L�
�n��p%yڜ�7GנVөG�cŦE]����7d�0��7��ܦ�uovG�f�0v��c�b�*��9��@�-9��+��J�x��#���I� ��.�UgE��Q�h�Y�V��|ܔsK
y�3h9�O��Iy�����;��Z�%�§9ȝ����ݰq��}���sf�Ø�ڇ���ʕ��o{0��`�)��{��/K�}ۢs��[o{x��T�μ�lg�Lp-��o��MNֶ��wq�=�"�����Aw��W
�z��Lv���S���^0�۬���8��%m/Z�X�59^U�g�ɋ:zz3=VW^��{CҗA>��_�f5���Ϩэ?J����>�������Z�kv�������>t<�P�>����޸6���(�C�N�劮�s��GP.E�<�#��#�[���9[(�nJ3�˧����sO���r���"s!�Ɋ$\i�j�{��k��+[�*���N�}Duwo���2�_y������z;�@��X��g�>���l<��醲��g>�k;�ނ���I��h�b�gN�yNZ��m�X^�ƾq3\:��%�2���96�bC-o��_�/b�6�zگR����g5v X{����\zk�-��R:0���Ld��,���R�;��_\�!2芈Z{]/��c�FRҕz�g7�{v�/�[W�2�Wql�}ܓzA�d�7��3��̢w_�J��	�U��}(������ҽ8�F�3d{aHX���e^ݙ"d�f���#�Q�:jv�n5qB�Ե�C��<���9�>�/�~�%��_��� �{z{v�5��7���y�g���9����|"	���Mk�T�ڋ�ƀ��NU}�?I���?M�U���}�e��=�i�o@�.��9T^����=^��&�!obJת~f��N��� V+��J�Y�s�sڈ��=C���I��+�����"��yx�I|��j��n��|�_��Jv=;>�~��Û'��k:����#j!d��-�lEZ�
%���}���7���O�S���Ws�M�7W>������^�ػ��#)��2�'�d�/ՏN��Br�y{�����=��G�����w�����������6��5��l���V;�ےe?�U��0u_�vX]&�<:���Zg�lufx��u&���p���ʱ��(�ͭc[��wT��+U���R��˱;,4%���]���g��
�W���GT�P��]�TY�Wn���S�g:wt�ά���6'�|*ܭ��X;Nbג	6�,��A� ���Z����<7(Cp�g�iwQ}��ջ{B����m����!Sc��M���a��)���ܖ�_(��X�.�M� �+3�s���MҘU�t�淦-va=��uݕ�/k��!��9�'��W*�H�Y�^���2�w��ʦ#�����.�]M�m�D����>�č�M�\�+j�����o8�v^.k#9�v}�:�e&ZThP*E�h���s�w��R���A-�.��ʴ�v�c5˪W_8b")�\%�ښ�%$K맹ے��Fu�����e=�V��n.1<ή��h]�ޙ�p������^���Y�DAt醯fj�y���q}��7
r7���Nȭ˘Ld��܄��V(�j�#��Ȣ��2E)��+[|�#o�}�l����MV>�߃IZ�[�� �Y������U�e��n��E�N�U�IJV�ggp�9kMaռs#/�%)hX�'��MX���0�^�Lt: 6<��+��E
��V�p�$�T��}��>�e��၆^a���������ˮ�1 ,5���KF�#[����9|ה��Ǚ�/ޫ��%[��>�H�Q唠�W�PN}]$Z�J��*���Ϫ�cܰ�����(�n�Ħ�܅e0���%��pY׉��N��_.Ke�X3"eW51�wu��e����M�)�wq�ԍ�E��ԹwP[�:�4�}y�il�p���Ǵ��
ފmK7\��C�w{v=
�^����l��cC�cC����:v�;ht���*{u�j�IA��+8�M6q%��1�v���W���2� ulsnU�}uЙ²�ή�wmk��xo7{�i�\�SK��ˍp����F��ɜ�O��r�+��;�E�7�+6\�ղB���2�nm��iwq�;f��!c ��绛bP��quZ���e��`<>-����c�u��� q�*���cR�U��tో6�����9�Gcٖ�Ǖ����}2rK�����%��@+)Վc~|T\4�[�i�ۂqK�]��ov^�p�O%7�W=ͤ�����V1���d5�z�º�#�����:�<�O�dW��nQ��'���="�<����,�p-����������_6�l��.m�J��j�Y�;ձ���go\&�wb�u�]E�Yp蒱>B�^�QCJ�v��"�oc�٤S*jc�����'S��Ip��zwy�/K�0����&����ۚv]��`2�l��&/�e�7w���
#XJ��J�^<|c�]z�����r�� "J��4R*� ��IT5J�QK	M[j��%�O*���4�1:^I�ш.g��9!���˄��i1�#X$'llbf"&�4�%��i�bu��m�KHs��c�L\�8�#r9��5N��A6�[#�r�F�f�љӋ������2LA>����i�,O$�p�2f���`�ETm��F���=u�n�p�9Ñ���(���6��U)ʃT�ֹ;�c�4'$:��Ƒ�(w76hxFۨ��\�ͣ���4'%�Q���-�ThMr5O\�Fu�r���A�4�&�A˜�6^�$둗4u�+��AW�4�*)t���y�4�-	HruEUHm�'\��#l<�)Ek\�!����T:"Z&71ʢ����h)a������_���9����Q�e�JӜX��Z�E"���f��Kv����$,��G�����ۄ�+ bxy�����~�fl����s'Mxu3�ne�(�N�Q�����59��$��:����S�0w�)���5)��Z���w%��#��xv��;w�n��[hZF���=5N��nayدm@|��Bn�+4Pe�˓x�n%��4]���PY�,{'��G�2��xӴ�6r�am�l)�PP7)��棶&6{��@�{-#U����U<�T��x��\��|bS^��e��Ty�k���)�^ھ������L�rK��^R,��>v^�Θj�;�L=(a�0��^��Xy�g;��D:��#$d�1�ǧ�h�H��r_�V�i�nyd�m�Z�.�wj�ܝb�֫	�H����$B�ݹE2��׈[�j������E'��)�A)�{J1�͇eT��)�^ܑEA�:�i��4=��ߙI�v��a<FI�o
�R��1%�2��mE�K4�g^*����=�0�������0ܳ������^<���D"��a��{2y�s���5}�]6�EA�i>�@�hm��K4U���ف��e�G��D`&H�c�s��le%ۙ\�@B�:<��{��y�ݴ2Rf��(n�Q��r�9��B�ؘ��5#H\o���;�e�l�똑S�������u
���s��#t�t)P栻y]�!z_j0e�%�2ܵ�Tt#:�U��>U}؉����G^�[��M^\��8ؠ���Z���RVgft�f\��Y���^�OI*Ox=���w*\׻(n�I1��ֆ��^Eq͟B	���/�Ko�o����mP�M�ZniF���l����迎�:&Xz��SHf�L/ϯxagX
~�
�n�������� m�J��e0�1,c�:�zTn�cm�,G�`-g��,�;z.��u�f���k�����»b���u�u�E8��2-�6�C�3:�%�M@`��9�Va.փ-3�ٔ�{xZf*+ڞԦ�!��b\��٩CKԓ�Y>-��>+.�Y�5K%E���	w���N\eǏ8,��a�����E��P˸��o�o:�$��zZ)i�z�2�Y���T�Aǆ8c
&�<�ex֠���'O-Uߍ������rL.�~�;�GXA�)��7�c5�FY��zYءڤ�����Qz_������ƪ30Ձ$�7��%�sv,_)���w�R���6�#����l_*$�v�%�d9����v�B֯rV��gT0ř��}���8Cܔ7*m�;U.|���:ׯY�o�exVϳ��CEv'sVa�7���aP���H!r%,u�}�7-��r�6�=�-088�{'�E�.�]�j~��ދ;=��=ȶ���{��F���"mէ�����u 0uwÓ地�����8eE�W=�Rܾ]�'���V���Km��}P^p�"��|0���^�.��Z�f$�:���Ʀ�����0�3y�b��l�Q�m@i��Ũ��~��{`%[�/9!�	η�mnz�i�����-��g��#��M�f]��[zv�ŋg�!��T���wH������A�:��
�CVe�YN��f�q�2�2�2� ��c����.�K1�q�2����]�n8'u�g�ݯ�"�Ƭ�xm����oO�"2��b��;�f�tR��k��g�r�&�Jb�T�GD�u+��9*^ԣ.��6X`y�e�����Tp����p+���Ք"VƢ#jz1�v��o�.�2|Z�0�b�f~��m���4���g�m\�hI�sb�{�8Ь�%R�c{�ߖ�k��w-o�ҍ��1�,��3
���nE��Z�
�;�$�`���	k�����Ӵ[ĕ�3��j9�-�tI�!�Q�	����R�W1��y��6c�X6j.�f�"�7�86Ӑ%Csl��h����6v��M8�l-��RN`����xjY��ȅ�^Bv��ץx9k.{Pt�Zcȷ`��e�O���׮�I��
);\x��:��3d%�A�ۧ�a��z��S��������Eu쐴:�<�y�M�L�I�ڦ
�3vS��f�(�]�j��ÖȂ�>#[�y��������n��t���&����	<���s��`8��x��
��o{����*���1#9ofJe1��K;�
%�\�G��Ar��HS�:���2_f�p5�<��s��S��;�ٱ���n������B~�}u��Y".�As_:n�9o��s��i���m��F��n�L�WO�����k��M��D����0�"��P#�u��/�4�'j(<K)c�e���Ly�(J)���4g�B��QWB�綬*
����5���;Sݖh�ќ7�β$
i&ZY
v�M!Ȉc09�����f.�k�v�p� �*&{5�0(܃�³���f� �OT;�$�7��	��,��-09�Uq��!��,��Jt�2�ʼ����H�2�|��zT����N#�Nx�Y��oe��	�>���=>w{��k��+�A�:���OR/nbS�
�-ܔ�b��} �۽4{H�Hw�8ݧ/���$϶q�Cݵ�F�b�N���9�T�}��?��`Ғ��E'�Q���c��pa�`��Np��Z�����O�_�I�!c��PȖSت�;	�D����	ts���y��6�"�
v�˰�/4���a�˭c|�|\��+����=Z�cbS'$�qX�a3�����4ɻ����.w��x�Wō{v�ɞ�7�͞9��5��uR"��z��2v)��f|�2mt����=�q��ںv�`{�utP�,}�1�mqG��m�s�np����=dl"����x���1Qkb5)�P5�jm�\kl���Z�S;.��n_��Ym����׋�ņ�E�˼c/��cF����z8
d-im�y]�a+�Yr�\c�g��/0j��0G����,y�%Z�x}� k���s�xŷ�)ՊƩ���dwp�u� ��4y���Y���3F�� ��'[5����c��[�U
�̡�3�R�W���lF��A.��6���]�f�h�rW����Ҷ�������E^�B��-W���Mt��u��ɷ���6��"+��5F�܂כH�G���cV�8�]�x�V>�ꗾ\E��+/�Lةiӌ��p%ړ��?q��鶧Խ��2��[xöp*Pmr����0P��5�э�9�&�},�C��Ma�_�ք/�"Y���G�^]
�Q�i���Fv���绹��f�M�$�6����k�K�{�N�� ��sTQ�Bb��"��L/^���"��*���^ú%u�d�j%�bW2�VN5M��xd.�7;�X�k!O�<�e�WT�s�fy�ɗ*��f�@�6�+�7��8G���Hf�jKTsre7|B���_)�m�I��^�{��,�q��4$B�I��ﶣī�ɎSp�{X(��iV9��k�gan���y��g��=����ԉ�{ƺpʒ��ILY�:�X�CZQ#nt<Bz8�� ��5���8_d�����W��!�S��~Jq���N���Fх7��m�u`�(]2xJ�w'�i�V��GCT�,aC�J.-̪<��Zrpj�}^�X�Z����BլG'F���:��zWS�L{��,��{5���[���h�E�X��i\v��+�V"%0�0%�񺩞j�Q�6�ڎP6$�C�`Y��C>k����d��^]�vR�Z4<����dmU�'ܣ��ז�'��f�H�#	4�
e�ֆ�!�y��lAaI�6qp��̊�������z�SBt�X�:�㩞	���Zӽ�|`��4ߪ��B��A�]=y��Ӥ�κ�lZz�R*�%Ra���ӫ��R�sP;������3=a�Ѽz;��ve%6.�I�TΙ��40�1m)�t��5��u8Ҍ�m؁�؈�u�1Ә&�Wc'�i��G(L ��a���])�[S��hd{��X	|��@�u;��%�̬�[�A�s�Y\�
:4� ܄O���7�\5�\w��.�z�I��W�v��c]�����u�{1�їp*g|̕�D[u��7+���k���Q�~�VԦ�x{&V�8���$L��Ch�a��/:�e������%J���T�΋��e�wHw��K��<]�;rLF���-���L\�cZ���o�w�][;,O�.M����%ʥV�x�`�7Oumw�O���=ڋPk�}j^�0�o`�VQ�Aח+`\�g(<y�fT
aB�,�~��g�r��u�vE):�9�5>��.�\�>3nz1��Μ�(Φ�LyR�7/q)����j��̦c ���ڨz܂�����9ôоTI]�IvC!��;�nkx��O���g=���BTE���}��s�}�U-|�A�<ҊN���9V0��֒3�u�/������?,��WS�-�Md1�>�tLG>�6�p�4�^?7a��)>�,�{9W
7%EB��l�ݙ}�Wm�㗑�v/!��y������S{^��g���/q\�k�2Y�)M�w��N91F�A�\��`��M��ӕP/v�9�6L0@�o#F�ݐ)�sPfc"�q]j��:76�9v�����v9��)�?bR�a��P�5��x���o@�� 盰��l��`ד�l@��x�1J�5�����D��B��y����;�з�W��6F�� �8Y�x�ޛ7&��1"Pjۘ��(����l��Sn�4s���D��q�ҝa��,��
<�l�� ��G�տ[��2��O�w�����٣������D���J��m\�o_�c�D����U�ڹEIb*2���+�r?6��*�=Ζ֚��iK3.�j8�w���q����L��9#N�	L�.�_�K  vr�WVb�R���G�%v�ܱ���y~�^:'|)x6w�k���bʅ�k޵���?s�䤰km�`���[�UGH�M)���6���� 3���Q�����S)쮲޲uP�Jz2�^��"o'(��|ͻM����Rkn�zc���c�-g�r��=�0q���\�&4:�s%�6�u��|:�"އ�W�8�=�5\ϏF�KP1ba�8f�6嬿�j���E����3����e��9�MS�L�:���8����c >iS4wLsA�LO@�]�.��1��(�k��ț���lޤF�R���-d8��Y
��'�����d(-�,g)g����L:�U���vV�����kyã;B�4d]�b�G[Q����C��9Z�î@���Ss�ISۛ�s1�"�V4Gd�N�~|N	��k�,S	��Je��v�)��w�&�o����B�.иx�w��҆[���*���G<L�ZY��,11����o�G���WF3hL��^-�޷����r�c�0�7��T���p\�4Oa�MQB�K/7�Tު�0<e4��l�i��Y���1欳���zđm��]�Gҹ'���ܤ$��Q�b���Q��us� n�<���g!�q`��V*2k
��qQ�,�R��H�ڃ;(`������kFyZu�VaL�U�ŧ��i�iH���IJx2Wc�f�O/)r����e��S.s�ҫ�~�R�o<�qNz^y���u��w�do>f�f��9pc�_ ��-�FwH~�(�s��;S�ܼ��U����m�^�>޲'w���i������z�d"�]�B��2h~�XM���H���J�|�B�Ơ�;�I��se�E���{0�aΩC �txȵa�=N�_Z�Ck�{"Xϳ�\0�5�=B(YU��PK���OQ`�.�����3�lxp���|����6���m��'�rbwqQkk�Ԫ[:�)�Ⱥĭ[D�ϰ��	���PZBֹv��y�hj�tX���2��2M���򠸊���}��6��K!ڕ�}�X�,�;T�U�D��c^0����h~2[aUV׵���*�{�>Cq�c(��W�b�>ī�Nj��kPz�����LN�`-dϢ��t����+���g��5�
�����a�-GW��l�����oI�܁b5(� ��b��d���{c�^8)�����!�Bؼ1��~S�۶��3u��[Ih�6�X�L{	�����S%
k���mvpG�w�Fj���g�lmw'��-�{ kxx�ݷ�:�|���#�P�4�/yL���UѮQ��l�Y����/k���%l��O�p����P�/�2���N�M���1ŉ��v������>D c96�	v��dF��*Fe���Y���oz�un֜Ȥ��!�[5(�񌞀��ɘS,�d
ݘ<c|�=�4� ����숗R�u��2�E)i�=b�k7'i�we&£ݫY��ޕWԋ��0�3�����i�j�ض�h�x��/�l��X؁�u�P6F�M~d1�ɍ������ֵю��$��tL�w�g�nɭySWtyT^���iݮ�+��>�;AX���^ފN��1I�l	l�T�;z�B�m��[i(��Pgw�i<��_C=����RM4�v�� S�y�bʮan�aO'��NNj�|r����1��ٍʧ�����nNC�;j�;�Y���e���uJ>Yb��N�*,�(�[���LC�up��i��#��z�e�bF��ie�:�؆�{�E�#]�a�t6���̽s���sR��&�����tm��j�2�L�ñ^1�[�07�$����B/�]���l)������y��˒T�jcl�~g�ݏ�w[_��x&�mKZ�[������}>_�����|�Ƿ埗#��|+z�ڟ<���/d.�Uv��8��Ωs�<�0SA�P���.UǶ;�>u{f���V�q�%X���#��d��k�F¥vr�ͻ��H{2��P�P!"u��.����G p�siw&k;�X���VC��J��Z9�'gsGg�-2��:]��Ov"�\��N'm��lu҅����p��mW0�M�f%�� ���б�B�h�~ӕ��޺��oץ�]�S��d�qt�`#����EZ;�k�ND�s��W/w�ZYϖZ�]\D5�t��C��h1G+���,{l嫵�̺�4t�end��M�Tk�e�(nW��\�ՠ����kU�z���7O6�w�D�ỻ�#h��,ILs��U�!#��S�HY珩�C@
�]�J�=��;�x�C�K�AU�wh"Ђ3���P�:�-�O0<��y�˸,#a��$��_-Y��B�� ����8.������e���Zǻ�1���[D���6U4��ZJX"[����FK��j��؛���
z�@��쾫�)��@�uϭ���Q����9^�����v˺:6�w"&@�s5rl]�l�Wd�sl�V��9�f�{�,����i�Ǘ�'rW0]):2&����W+?f�!or��]*s�_IN���vH!(�e�=��t|��X����J,�Pڮ@�4�鱫�T�;z��u!L�}2��jp���en ���P�Zю����{����+Vwd���R;]W�Ҿ�=����F$�g��G 窲d@���;�V���{��I�w*������?|B�*!D�3R&����"Wq�V_c/�����݉ ��Gyb�jڵ��a�{��]L�y�cy�WG:�ǻ]��ܹf �8�$-���w��m(��8AI�;�.��Q:�դjBr��a���5��	g���e�|��.,\}�5F��%���D���Ѥ���t9��α��M�v5��*x���WFK��u���;wt�h>Y�g���+�z�#l��Qf}��.�M��g��3�"�|iu�q�0�u��s-n�G^�]�KQ��b���T*��ְ��9�s�N�ز�/�;9�0��`����ݺ�E���,�r01�<�v�M%�B'�N��Z���bһ�����e�Ւ����� i�iwC�����qJ�8i:�'�"�b��d�V9Ox��/����r��+��i�M�7f\��[�1��D|v�C}Z��6��{)�.TƗ}�(���V��fwM�1�w��/�4ΎX����Y��K7U'�kxl��MT1�۝�.�A����ޤ#�6_}�]ўj�����j�n�kN�:�I�m>1��ƹ��=[�X�*�.�Ǻ��_r��3�����^�t��a�&]����,
�]��3���V]䮗��1��s�G"J�V1X{.v�p�h܃�L�����SX/�6O^���I��{����1\�[��7޶�z
xq�s�%�6��&]��o�C]k�w�y��V���Op�����Ţ���e��^��cn��mPuM?��(�H$�D*��s�p�Z��|wQݨ��`���OW'��G5��M-%OV�$�3Ɉ�h#���rq%h~ 9�h
�h�kKHi�" �(��X4<�4��1� ��ܸn/$�DRP%PV��ʒ���[SUF�Fm�5;!(��Zns���r��Ӡ����,d��$\���h�b�+K���� (�$H�b#��h�7.P�9i���9��TBkE[b�'	9cb������C����%m��
4%i�5�nc��J(
H�4�M)��l��9�Ql�5¹��$��cF#D�I�j$6ՠ(��l�:9r���6�-�������s�����>i.��悖Z��X�j(t(�|+��Ъ�y��\Yk:ho��:�3v�r���j�:�4���t�\�!�'L�y"���Y����*O|fkʞ4,�)�1O3��,��]f���>3��6�%�3R�ֈ*�F^�Y�A�9�5�M�\v�zO��Go���P4�# ���j�_�'I�bv�ܼ�Cb��`�������Ŀ�ZE�~hn�d�#5Xs�6���x�wۮ�x�J����n��	N��b�XE;�#�>B�(��!��<౳8g�m��K61�v�z�cL=����	e:�1��	���&=��Pn�~fҘ��(��.�;j}�l$<�6qZ2�(�P��u��������Jjs�
r�n��i�v(v�'����Õe�\E����N��P��G��͏ՠ�J��ߴ嚏?Q������Ai�x$�<�a�04�s�f���#���׊������a�*=��*?{�e/k�����c
n�ܻ�0F�*�:9��n�Gۤ�z��V���d�|:&#��ġv�t��[Pބ˞�ؤ�C;�1�CB̍�P{x7��e��TFl=�pX!4�W�-�M��C�0r�mV�n�����g�;�B>������0Wg:�[��Y�:��Z���\'�^�"�\:�t�O�iz7?iW�J�z;�DQA^���W���~��k���$���8�ɭ�R�.ʧ9fd���|�K�orc���Os9 ���ׇ�LZ����u���U�Ϫ��1ǝ��������ț�b���eG'!����)�=��*_��O�3dէD(���6����̶���r�/��:L�ݯ�%>�W���w�J��,ʯɽ�����r����Q-s����l���	�N9h.�g<��2�i5)�^���L�oJ�l�:��O��Okv�Qg�w�v����}-=�^�jcÛ�ױ�{uE�\�:�xd�Lc�����>��7��4�f\-�֚��tz�$c3����N�q��j�ه�GgJ�/�jߍ?��9/mG��ɬ�vMD�D��}3��v/�Q���^.7���>���jsb�m�GIoI�J��T]yV�t^|]��m
��7�Z=бG3�$�ڀ�zc� ���Qp�\�E�a @}k��'W[��K`h��7m&f��,�D����|{5\Ϗ^5R@j.��@o���t���5�����u�dUj��� ��2;7��������;ʰ����>_@	�90t�R_m�;����(�;ǧ+����"TR�/e���yeV���ӏ�� �B������� ���t�`N���S���ؠ���V�-�ʯ��)ƽ�]�� �^�=���-g�ʲy���:���z&´��Cc*d����\+�.@�]Y������������>���v��4�t=%J�ݸz�55G��n"�����+��t�����ɻ]{G6%"������U���qŞ>yr�6F��C�.�z�zl���Z]�mG��M����z���裌�f�&i˲OL$s��'�9�b�t�cG��#Z#R�ڽUM̈́:lk<L�%%!���҄�:v}�ԩ�ܴK�tP�X!���Hr:F��3�������+��2	C'�xn�����	fX�v�՜'�D�L�����t��\�TKY�&��Fm�]��x����<g�4���,�ʪc�sT�u��`�B������5PKO�>�����ְ�������Z�1�4Y=A��*�v/	�B�̬�l�S���-�l�a���"̻u5]v�<�m��9.��'���	�v���Qq�iQO����j~m�&{Z&K@�*�u��'�n\�]�5�K����W�;k��K�b�i`��1B+��\������?=(�yo��c 㣏M�N\5��7Y@'��5��M�7���W��s5�+��L�@O�Cy�����[J-xC5��;bp|ok χ�ޚ�Vt%a�7
��V�^�a]J��
���lQcq�	o1 oC;P�W�!�Q��� ��h�V��/��=�o��5���K.�*��z���1[e�J��׈8�]��t�%�M�{�sA��m�JS��U��$W�=��%��(��x�n�i�sr~-��m%X�yO6��K=���9[�[��t�lm��-��5R��Yr��r4]Q��ȴ���q�ŵ|Uƨf��Sq��6y{vS�z����� �r��%/_nޢ �`]�y�	��JOF����W�P���ӯ����XCR�:�OM1���S5#ٜ;eHg`�!۵��t��'$�	q�Q�H�n�����;m�s�-�ML'�h�^���R�Ű���o=��8�t:%`�����pz���eTC�d'~}g���R�����˽��5���XS_C8#��|�=�����yC�'�c2�RFuLGXx܌���!��_�#�$%)��%sM��]����u�0�-:KU;�Lݑc8KgR�5��ff�j�]sR���;aM^�ɲ�-]�b�ƪ���xi���A=9쮸��\ǘ�*cm�T:��8F�
�(l{��c��C��ϱH�Ģ��%���"��t�����띭�z��t�����Oz�;z.k�����Х�Uw>�� C�X�NgS�`��8��Ǜ"�q�Z���^�����[G1���ù�u:��UҰk��eS�p�9-�C�b��7�Q�w\��
�A��޽}ʄ�Sd<t�6�����sq6��9�8�<�sɦǮ�ϴ,�Eް�m���WI��0Q��dy:Cc��r�%��� ��lV^�N��C��?����F����b��>�/'�n7T��b�K^��醾l`�/!L�w�]�V�BY(���� ׶%�2Ĭ���ܪ�}"&�T�k��y�P���	�l��pc_�ݻAf<S'e�IT��]Q�F,tƶ���P709�����S7[��_0�t\��ٺ�OF���L�=b��w�="�p��P����q9/�`P���	#Z[B���������s����+6�s��Ea�2 ��6�%Ra���Ӑ�g�tL�5����{����3���_�9���I�k��2�Ū\v��zO��Gh=�q�2!����mx��<�f]O*\����.H�S�cg�cW�f���,�r֏S��G���Ղ�͡��nzb��Yti�aSL��u���r���9��B�ϡ��<��<ೇ��1�6�z�5A�F���lF��a¢�x��.�^O N v��wJ�u�g&�˅e�\<�V��n:�ۇ"{a:u
2�·�f<�w��ꦢSHwX����F �L���;ڤ����<�Y�}橶�{�~���Zj�wA�7���]i_v�Jpk�����f�v�y�V�<p��q-����OJĩ� ��j�\�o۟�o^�O�=.���� �R(��U>�v>U5���o"�|����؁]YWs����;r���������I~���*�F(�h.>B�����mF���ל�ڬW*$�ڤ�m�f�	��2`��Zҭ˚�1��'�(Dx؇a��޺\T�ܕ�O���r��vyyS�F�[B�w�F���*�L��zs9����U��b��4!��?��as��O�����&\�ڮ=%Q���Q}=VAܓ3�����=���-}e��M��P�H8�nY��mPŗ�.��I�T�>圉�5�|N����_љޮ�4`O7��_l�s`Q�D2�= ��h|yC-���r�������d!A�:�3OoJ/~s2��	���%>�Y˭�Gg��!�G4)�!�B���b�N��q�K��2χ���VV�0�MJb��ϥ2���
��*sC�n!�k�^�X�ͽmk�-.� �T�~l���f�VU������Sь$d�X�0/ҊM��U��M�Su�,\E3;s�k�g�O�vnW�s�
�U)q��=N���n�R9O7��3g<�B��~Xjg�
�?��̪�A�0���6ld�8���b�5���*���~O��c)1&^p��~�~�f�U�[З/U�Z缷�㋯�������;48[���Q����5���E_�9[�����;72.�����K��u�5�f<�Smgu[���gTCK�K��}u�ڮ�f�9k����.��c�l��dB#���{�5sm����?a�_Y���SkP&1��������E�a 86ӍB�;	yx�%���02��!�����@9���S��N��^�t���T���Q��K}�s�sy�*�,���%Ի'L&��-�:��wlr}��lx��)��h��LJ��g�#9��ƾPLZ�Y�&wu‘�+[��v�����,ؕ��}�x�w!���AQL	lAΉ%�u:�ږ®�%��g��S�8K�Ϛ��/85��<&��E��t�ݪhj��2�
�J�p]OCII4!��⯆���|}0�u���C/�}�ؔP�~��py�����ZS4�fb��7�+}Z�+e���v2�q�����[,�N�w<0�4�����)�C��{� ���ff�J&��~��i̠���T�Ǝ�
Y>�SL���Cz�D�]�r��=�<MQf����{��]���#��n�)��+\hn�U�20�0�7�S-��S.s��ֲ۫��z�q;��@�n�m�����-�m����:%�N9�Q��'7 �;L�u�XOt-l��l���q��]����֑�$xaȅ��|k٤iY�O��`T��Բ�`�����ǳ��>^�H'ͤ	͔�����kr�<ڮ̘��3���[M"�E�lH�p �qb�,�J[]Kl���lq����;Ra @��Ս;!��s4.�L�Ww����
��q�@f�[�� ���OnJ��n~D�&w�@=r-l�6X��V�
�͐:��[�A�8ͪ��a0ؙ-{,�uMKT�r�&��<�������m��c���@:mCt���(<�Rn�MIC��{����"���=���1g[�[Fk�KۊǬ��_/DBm�m���CL�gGW>�3�J���:uEܶ3���r���qa��1�n|�ن�k'��k^ɸi[.Sh���Jo���j�7���-vD[@�</S-�[�lEv�e�
��A,]��ߟ�Itd�֮��O�c�l�t��1>�e1:�/~��������ȫ.���s$�0�=\������}#N�a�:�ZLN�H�F۠��hPڳi;S��c���4�vN$Y�=I1|̛����ʋ��wl;w�>s	�{ݓ�r��Z��SRE�h�3eù�tk
&٘�@g�w.h
�fE'��k��V�//�k���tb��V�0����,�Wg&aM����X`�����!�Nq���+���)�@W��s�Ѫ���
igfP��.�����0K�ԙ�f=�ː�և)��VP�%J���<����6�t��ޯ+a���ve��k���E�@�o��8.t�����X��h{�.����7w�r�͢ir���=���`���� �ؐgC�h�g���Ͱ�͉��X�R���lt�%�}}pX/u��|dL�����`���ji�6�y�c8#C�TxJ�:/�u���5z��i�n����嵭v�u˶�l����,�-U%|3+�h�81�f���(TpKO�"{�|u�d��<�)9�ڨ[m�vl�M�烒�n��Gn^��r�0����H[ȵ�Z�ӊ9���(���*�;�;���:�΄['���B1ؖ�yJ����)���
i�d���{����B�Y�V��}�\���DR}�R��r7d�d;Nh����{`�ln����ŵ"�
���:Z[���e��56d>��������f=��dᰳ���S7[��6���sSEv�E�YʏVlT��ا��z���О�2Ynx��SMY�KX�6	�v��^�Ӻ��ț����|`d��+i�\���B���͇��Vl�.�3\�c�aJ&թ�S��..��4ë������g)�T��1X��GO`��N741���x���T��΍h֑Y�����fh�Q�c&���f[�S�+�e��_�* Z~�	n��]���v�2��m���L/z�v_�i�:��%�+�뭊�q�_kA�z�.qs�[\�75VҁvXXf��;�r�wim����4�3�E�_���7���<Ge�b�$+U���p�o,��(pTH��$:9�KP���G���倶�6���i#99x��
7�ys�����¯R�"�GKz1�7���'���d6�\�d�IR�.8�@��wq3[B�%^ՊY���;�j-A�ҹ��x�M��Z��!7�г����U��ŉ�9���M�xV�Și�
͢��'L��,ؕ�3�Fm�s��C�]�Z�xl�7Nv :{�&��]��Dˍ�f��|��V3�MQ��D�sMR��F���ÙWL�'�y��p�>�|�G��e�#�^�XfBT���eE(��;�1��㹺\Τ��Zdٮ�Sj�ws�����:�~L�?/~/���u��.�b�pkW��f_f�����W>�7dE�)�^i�.��v(�vC<��ײʚ%3�b�fI�q��U��Od�fV^W�2g~�o�̢���#��kǫW�6�;V��	��ˊ�sF�%�(0Cw��=h�N9t�=׏���a!�9�^)��ħ�*�X��u�p��o��x�|�/�����|�_c����?�x��˾~��\��#��pA_6У5K�$U�Z��Uc �X�Řu)����c�V� ���|ld����[e]��KNS����E.���e�e�%�M�R�qYUв�eY��Lp�|y+�M�:��b�0���Y����[v��G7n��_ʎ�Zv�b�6�UY�]��O\mR�#�u7�.����Ss�v��Hv����[��WR��i�������9���wp�w��{C];�\��X��f` s��۝����u����k�(&1��F�Dǽ�8+�i��4�{kiL����Q	ٹ���[�����lU���%�:��ۥwW��QS����-�q�]���z-�����].m�V�o7U��е��N�3�,T�93�٦��tV�0���j�!jw]e��XɽU���g$�+��;�B����W&�p����k(Z���p.��5�ת���n����<��C�eXظ�[9�7;�U�fѠ6MyL*p3YZ��G��Iݤ�6u��7�-�[cfn�˦��SG�CԦ�`�ogp͕�;ls�}�}����m�\�X��mf�t	��A��*n�(�޹'�G[e��s@��e�편vVV�}B�`c��ycn2�����aM��v�Zh=��K�bv��#[Qlz���̡��,�-aGs-mh+J��m�F�`�dXz@H�z�>�YX�0��(>��r9@c�������2�5Ԟ�-k���;7�#�d��:	�޺�^(z��=S��H�圡jV�Zi>��N
ظ�SS�.����ϔF�w}Xf�7/�,��]\:�KR�^�j�qGJu>�v�Vo\��Ѻ�Xu8��&��r������f�='{o�נM��73�֝��(�:�gܱe.�]��+�yHN��YS��5eY}{[K�]nt8�p����r-΋�I�X��u�WS;y��{��B�@Mܭ�՜U@���9�v��{�6��z��&���B��MK�sn8\7J�U�S���`z%Ez�ثS�S᝵÷.*|�f�Y���3[:��=�!�=��ψ�Ƹ�))b��Os��S.�Rs㧜��v��ʹa$�i� Q�8)�-��c��r++:c�;I!�S7E��-�
m+t�F�}�V�tn�����mY|u��FU��u6��~u�jf?.�NLc�1q�iޣ�{Q�u�Ň8���]��	�l���.�[��)M�.��6]<���o>�f�ڬ�����
�0�ڙ�M�v����&1u5=Ws���\@��lܶЩ�(�}Z9[���ɗD!�-ի
Gd*��oT�ޱ\�`S���p�Al����・���y2n������@��l-���m�ͥ�����'9��<׈�ӭ��jM�V؈�60�UZ�m�d����t�g͡��9Lr5AE��h��]�A�H�naҗ6�d��"t;j,cEZ�-rNZ��mM�**�Y�J����4�v� ��-��6�M\�I̓E1.v��66-�<�l�k1�(�W[�SCȦuj(1QZ44m`��<�#���i���%����(���Hڍ�Ί4������V�Sr����a�c�V��kf&)�N�m�g��s�h�h1k-ͨ�ŝ�l�iqD1i�<�UkT���'lcf��h�i3Z�#cF��6-nN(����4� ��'�	"�	_[����w<M�Q���g_�]��qW��N�cB��T��C��9���EprQ֤it����6���y޼FQ���}��}�� <=б���ݖߎe��~xb��=��?^L8x�&)��Jc�}.+������[�זE4^�-�5�S4FəZ�Ox�.�� "��	�6i�EaY\P��d4�ʎa���n\�o�^Us�M�5��,v�us�c��؂�fb��k8���>��Vl����E!"2�k]L���W5�&�����q��ǁpG[K+h�1�b,O��g���I��;>���'�r�|sk�X�����7[�[���H�cе�tj���cɁ��f�mK�ะ������P��N�=�[=��k��dƍ�s\_ַ�	��<��X��5�&��f����V�A���S��*W��"RB�/�[M�BA��.�-����2CkȒ�C�f��L�a�ҁ^�m|b�)�vI��&�eɊ7���Z�}5�R�E>�k��fK��6	v�bl�ZFy�Ww�o�|�[��]Ey��g��:z$ƶ�L$C�P+�Qg#۴�v����^<s��Qy0�U�.}����k�偮HT���4O�>ݯL�
I�N�t�x�W�ZЈ�J��#ڶem���uUBe)��$U�|�;/��z��W|,\͵:��IN^��dwCk1���᫖��.��n�*/+VG�Qʔ�f��V��@��S!W�� �ф���yF�n�c ����k�A�g��?@�R��oc窃���r�,^:���xx�4w`�ϵ��`�i���&�W"p�_f��ùV`�d	��X�-r:��l��za>�s�\a�*����k�Y?X�4�lb�omx�������;�~���[�����^h��"#y�7��.Ʀ��1�C8��8�}ax�̱��s�T�u��a��̘�-�0-8q�gs�����/o��>���	Ʒc�͂@~�T��<�L)*����n�|��fTdBv�m�!�L��k���s�7y`~`2)�3�i@�̈́;\6�#�9�=�����M���p�dft='�V��zSP���T���ٟ�û񶅎�r=O��Ue������-�e7��m���v�e�!�Z/a�貁�pv=66�-dH�Ǭ��_ �=��t�)h[�����Hňd�&��`\�����J�cj��	G7b�u�k\�\{�k���1W��,!��:�=-yN�5���㦩Ȧ�}���4S��,qd��s��kP$d�71Y�4�i8��H]6i�=�k�^�۟�='>��sI�6�p>�g��>�b|�O�ܮ���{��a�웵{�'*V�NU�t}�d><��SvZ�口]���X7�ɵ�ڂ�]��}42P���������|.������p����f���n���}|(�׍k�Z�pg�[ܕ�+�:m��[�O5�~:��ͽ���J�`�WVY)�AФ���}UU��"���s(	c��2ߘY���ns��k�C�����v�l1���]���X�Y]&]he�$��ut��R�Gc�W@�z��TPE�CP�-S���E��vܮ����ъY��^<z�d�&�Ǵ�������#ag��w*� -�<daD� K��xhNSĽ���4�P��'���,�Yx��jckV� ���lU�=SK��Ph�&��exӈer��WU�i�"�N%��5ۼ����k��P���g�I�_Z,���[��b��{Y�v�Ŷ�0���|�[^�ёL/�I��1�a�7���t4҉d�M̶h�ց^��b�ɖє��Uȗd�����!���!ED5�P)���Q�ha\{��q�k�g��;�9KFEf�T5p�W�2a�Z�h�k0ڬZ���&Zd�v��7ʹ��(��{v����D�z����d�>z�U뢢ӓ�U�62i��l>��>�ex�[̼t��/l���yǹ\Fm�܌�N��jJ�[���S�vJ�y��(u�UІ�w�dTE��σwz�oPI]T&eђ%]F���R��Q���zpn��98c�V�[�-�	���M��L��������
m��ԘsR��oe��J����p�k�ٛ�u=�ǭ�]\v���*PXl�7�L]6QU�����Pڰ�U��6> �>o`< ���{)�����u�ö{s�KP&�Y�Q�F,tƶ׊9`���w�ϭ�k`�NwJ�]V�T�{W'��͘�9�!�+�&�y{	����dwj���3�)�+�Q<����q��#�Z�;�g��pmҙ�����=�ĪL6�)�t�6=�ڙ<gF��5C?m�1��8Ϩ� Xb�X=��S"p�Iֻ�C*�/����-a����C�6�Z��(���5���fq�t`w�,���ĳS��of�ϭA��)�]�Z�rt��S\�T�`�qf� ��n�k�a�u�µ���S��L��	^��Ҽ��z6/��^D8��ui��x&�3F�3`�`�z�MAnn����z&�����Hn�~j �x����Y��im����i%��M������S�[�����tYzm�X�Ϭ�s��n�N�;T��;���)���OD���r^r�����Q�<}��J��ev�g���p�k��T ʹH�˻��	�T��օ��:�i~rO�$�/\9���e�P�w���A�O���de��}�!@��?)H���OX��ޫ��췸u҆�rj�n��	��;��1v=sMgu)��}�7A]L���R�>;�½=R��@t��Y�[Xjrq��Fͥr���^�|�V�N�<w�xn�lΠg6*�;Z%9����c��k
}�/�O�����ot�כ%X
��kP���P��P�w��=�����_?=W��~4N�@��T�L����UÜ=�Ԙ� :Y����P�����e�x�U.�7�펷2�P�.���R~�[B�ʨ݁r�䰈�-�g����YSG��b=̞�Z�ߤ=���m�+�L�{UcktB��̢��LɄ�c�lU���H�Z���e�����ռ��oK�<�=Y�84�m�R���t��>�S�+9t\�Ȏ�E�����V.�f`���X�b��g��ن�ei@�jL4���>:�29����[�a�cpuX�c[���Dw�_�@��[.m��&b�q��>�QB����N��f�"w� :L^�k��ϰm�?��O��`螟-@�������[^����ó���+6v��3 �,ט�מ��a�/vl1���T��[J6c8�Ň�`����Ik�X2��پ͈�+�	�E�C4�pv�A7-G5�U-�t�:�������@��t������m�ժo�U�6���W@��q]�����~x�ޑ�J�hzv� ����P���s�iܢzq̻�Q1��n�:�#D͹N�o����9B�)�F��������	�)C"�]}@�P����;x�:��yA���X;Dd�\TTo`3B�9��ItB�{����r�B&BB�:�o��-�����{��� ��0  jvR��~%AJ�0l6�	[�˖e�m1�b"ؒ�ٸ��d7W[�wΜM�<�We�D�Hه�'xk�:r�n��:Ui$E�����8��yPկ�ߞ�16X���$�O�蝡���:��[��k:2���x*_�*�+�+Ã���46���4������o_p���]���4 �=}H(ق�{��b�R<�x�@z}��h����~�Of.v��ݍjP�Sk-"I�!6�*�V>���|'kȑw��A�`���UX���ҧ'�88��k�}~�A���jFD��@�X�7�����4�o�{h�b��v�
��&�����waa	L���x�4�4��R;��1�z�����^%��]�L���ⱺ�-�ab��h�5����L����b��ِ���kH���4�uϸ�<,�A�R/a�Jr��U%�����{]��;���1WŭG����4ѤzJ�'�E����d
q��ei@�͎�����1�z��4���W�i9��<<aƛ�����8عƻq�\1ib�m�Y�.�Xz�[�\ɝ�[�o�2���(vPjM7�lv�l�G$���{C��v��\��^�R6��C�Sm�G�#��Z39���XT�EE�=���:��>�[L9]�W��\9۟%u�b�)��:���<���c 7��%k������zW��/~�7���~+u���B�*P-#���� 9i]��d��$��+�{�zTP�\�è%���C��>74��wv�c�|6|a���M�t�h��/m����U�)�
s�L�ف���Q��o@?>�m(��ז��)�rl��mv:�y9Z5=q�"��;;[H�y�ܧ���-@Y^v�&�Z�H�v9�np)g���߱��gj$Cq�@���0-����Pˌ�� ������;YhUNS�7/L�^�@�/�&��\����Z�/;�[���	�ָ�9�LQj:�<�:�s#[��V��<?ikeuΩ�`�<�O{z�X�x�G^C
��V1f�e��J�-B\aQ[�Ͷo��F�:�
�\6:�n8[;�f^<�۶�ר��{�����}�<`iD�"]��3��L�W�qCf�*xN��B��1���!�"�6Nx�{y`l�m�aL�����X`��!���fS�����ez�����C/EFc��{��&�u4��|a���)o'b�W4�z�����ou��ܱ6(S��u��k�B��t
�"������H��V�����D�l�����G�X`R(�B3*�6�G�s��6�����гu�+�QZ�E�z�*J�mwf�%*g��W[%+�8cj�%�G��b56�\EP�ǽ!Ǜ�B�_w!����#��S���6���XW�]9��6GI��ڲ�L�WW^<���D_�
� ���S��>�'a��v+%�	!�'`��; VDu;�Ҁ�=��A�x8�;���{1�I�n�A��Zaꍎ��]o\`K_fi,.�5�V�=V�@w����gJ1�`dph�S�!�7o�[�R��	�mɕ��:�������-V0֯q��s���$AM>�0��d�T�������XS��vu3p��,Yzj�t�TR������@,[C�J��@�h�Y�B��}��=�*���~NgVFC&�xln�1.ټ�A7+���.�!��A]�:�����NAV�-��.�q�M�wړɆ�����ـ�Û0�²qP���<ѹM
�13�E��ϒ���m�۸��.��D�:INPߡ�!
8�4s���������.�0�Q���{�ն�8�ok�w���z'�j��ZM��gR�� ��U��	�5���41fǆuFu
9:ҷ�q�ƄyY޾��'�z��Cu�1�K�rY��cxK k��Q�Q�� �ʞ�f���a3���pwhu��];���.4���x%��93��o{�3H���[\�c�6N1_	rmQ5g��������EwCds��ݝ7�����wf�V���$޹E��O@N;v�#����u���l$�!Yh�9����X��dv+:J�x��`i�!��k��4 8a����ύn�����߿�����i��Vo{��^湬)�yM<�޸f�;�>��U���3�߳Qj���S80�ov!l'��283�bj��â��K��K �-���Of<�f�pJ�͏^�#�$��2��{��_�.sk�M�����i�zכi���*�8�����;��a�2�j�'4.��r07��Z�"���s���qj��٪�*o��v��6v<��o?��^��p2�G[�<���J�a��t��a�R���ڸ6m���u�(���&�W~�*	U���u�4G�`�B/���Ù�y�U��vyѼp�Uf�C�nBIlk�˞��'�+h^��q'�zȩv=P�`yo^�=2�����ӗ���Qa7�
�3H��b��*�X~�I�
5�m
ǐ)^��Gka�c�0��}Tǅ�	o&w�xq�A4��G�f@�48-9�3!y˴�:�iAtS~*=��݌GFM�C�c�{�`'*h��O\���u�KL[�0�G�w=yO=�b���QL�c�)�LV�e�%�h�$e!9�5�ƣ��R�x���g�,��9�;��ڣ����թ�G���t�N3=�9%��b�׫�sY���-2�ٖ��J�T�b�Lu�p*��Ǆp�y&;}v��u@���D.����b�3��{���)j���:�ۼ��2R�UrU��݁!18����h�h�i�Clѽr�;Ӛ��x$�YE�t�����SC\���3����?����o_�S�EJP�J�7�0�����'��������խ�o�䵻��|$7Y2���,Y�3&��"�[�����gݛ���Ii ��|��Ȉ�o61}��|z�a��Z���lǰ�k�"ñoa��9�O�l��u�m��BwTWn��Hw�P~|�?�����Rc"�G3�x�Sk��_AvŜ6�L;��P�'z��~�k�pp�B���}��}W4ŏu*-��f��\IbXn�g��>��k�N�x����Y&B2���-�O9i.�Aח*��`�lS}�H�0iqX�k�f{��͘��B��e&�Z0~��nSQ��C>�;��,U�:��7�k!
�-��ߟM�w&K�g�Mqj�B��n)��5S?��8z�X��%�w8�+��Âu�~����.��0����IY�v^J1��`���!"r���p��,��`�y���d�2�2�9^z�!4�i�cz���q�$+���҂�},�`��a�i�2��`�1�W<�G��u3��jmGC�3��kɫ�M�o)d���]�8�� �6.��ۉu� ����^�W������G������7���l��9,v+��F���Qky��N�w�P�K�X,��A���a��P����6�ޞ� Fy���yVR�\�/tӜr�̙�2\@*�����{�ҵ�T�e,�s�J����J�:W�n�X�9�[zL)�d,�w�u.U���徫�4`G_F
�]�:dn5�����OO<�E�&��v�B�lsm	��{EkS�[׃�i��LJ�'gwf!�Y1WdRJ;P��p�C��Ѧ�qd�_}uĹ�mj�Y�,�mv��1ҝ��ugZ��a�Ũ�W�ӟF���X��7�X��k*��]O�,�5qeꫝ����!�خ���]]K���j|�C��^Jv܇o�{�K�4uwPV�Ι�P��]��JY*ƭ��w�xm�v�s����8�46�A��lٚ����n[� 5!��=�hD�Mv�{���^�����py$�86	���z�`�M�̻	���:�/R%�	F�	��v	}&q��f�LM�ذB��C�d�/A�p�=�'�;��l�P�Ҕ��xA�R��ƕ.�8��Y���v�m[z��B�^������GX�ܬ�Kq 4KY	Pg�8���n��-�lZ�����"��|�d`�u	!�!�#���d�;�P�!���8�ڽ��1h���F��U�����(�lva��Gk%��Xq��_5Jl9.sR��T�v>O�J�oIvbY��|$+x8;�Y��jJVWn�}س��ir��ٳh�����������N4ޤȦ�s�n��pT�5�,�A���:�����PoB�/�.���Wb;Lpͧ�ӗL�A>v�����X�ֺ�b����֮#��W停xb�}:�Lٮ��]Q��]]r��vC �b�%Ck�/���!��[���wvlY�@e���5<ȟ��ݻ�Q�Q��̉eÎ��:�iA��-���,䨬�����P�	c�s]�`��z�7�UZ�V�ڨ��%����@�5��n%����6�gWc�kZi�
�=V�i�z;����M[��>�a�W�L��|�Z�l�r��;�8�B�η;0�ojek��M7p��F�K4ܦ�P�)�C�,>��x�aMy!��d���Ұk�;�̻;�Hf�K�=Z�̙�emZu�OyM�6c��O��M��-�g�W$�S�e��V� U����|8�Vm�o&�7�s5s�Ժ�dsr���t4�9��עZ]�i5��:p	
&Y��ȕ�y��u�}Z^^�m��ܶ��0wr�s\�'���"�N�B�aܣ�A�Jq��/�Ζ-�T�ʳ�q�.����+V�`?0��sVzq�sz�U˓��ц 懝5;
��l@s���{�ԥo[�C���vm��Q�5�{����3�A#\v�ƒկFYk8J�uR�]G�9���W+ޤ��ϡ\.g`9�8*�
I��e��Zq�X�T� ���^��ܝ�ҷJr���g38�j�w^Q�n�
	/��S_ś*�BiF�d6Q�&��H��Q �>N�MF��DkEV��Sa��A%k	�m����`�i��
,y����E���Qe�-�����K�J����g4U����m�-f*b-���kcZ1U���bq�6��&-�m����v�E�j�Ţ�cE�4�U�E��1T�sl[U�����Q�툈�mDD�h�k�ci��ED��1kE0m���V4kUE5EQD�m*�f4���5�TD���m�[�j��cA�*����F����I9�ʶ�V����6�b(�Q1b5Mhՠ�U$S[�`�Lh�lmgm[Z �t�b"��b�s��N��N��5�QL��U3U5�U�ѣm��c0i�A˜�3D-U5Q�l󚚤���f֢��9�0@Q5_��]���u���}�5{�%.�<K�
���q0N�s�ëPa���#�-ST�V��nV��V-}��Ŏon�����Q|Wu�F��V���W�\�{�� 3xJh��9N�� �8P�K'9�f>q��~�4��x�7G��Wl��j�n�)�K;���31{u=59�a�O=Rq}Ln^<M5�j��svmQ9� �]�|K���8��93v�5i��k�mX�U�Q�:�~�u������＋S>͗�O���ZP26Y�9!�V�m�Yo�ً����t�<���o_#�ui�k�GE���w�mz_��C���L�������k
�oH��3b
��(.���c�K����bY�Sp  Bv�4��n����OUnV���L��blz�[$n*-lu)��E~�|l�s�[[J-xC5�4<f4aF5S^����C6[��/�`"��@)����ޚm�S���-�|�8MV��B�z\D)�5���v�� �e�]���ڞ�fཇ�+̰֘c�><��#q�5{)�Mfi�	`�$u������b�:�L(���F�u;�[����F�g|s#�P��t�0�1�*'������(sC�"�މ�(�ߌ>W@�z�Қ���������{�!���#��I��
¤���Oe��0�un����f��b�-/?j�na�Jv{��,|5��sf#�����}t#��SQ����jyy[�#��8A�������>���]�4:�!j�W]wS��Bq%g#��*�n�D j��K�̉r԰������3 (BaJ�(JF�$��o ��S"V�xbf��h;|,4�ץƵ;���~+
&�x�j|��L�Z1kX�y��V�c9e���[��W�NNUCP�*���F�n�b�S/_K P�<c�`��ǑP:w!���m.��SL\$�/��m�7�+�a�O4����nS8l�m�u�;�׃�����?M%}C�=��#3�@�`l ���is���U(dq~�O�����4�p+y�)�\�u%7�$��KG/~�љU���,P��)!J����%%Ж�PZ����˃�&�� ҈�ڦ��]O*��]y(����E6$�1�lk�Ӗ�f�-y��`i�=�f��+t�ɨ�*zFe��LR%��Rv`ɧ�L�{�Qi����5�j���{�NC�;˦x�4��^]���m�F
���ɡ�(L�}���=�Qf.PTE'�IP\�b�A\�i���[e-�D��\/_�H��/<a�"�����l��M�.�r�=1��
9`�;M�����9Sά��1܆����:/�`"��ϡ�er���&^�f�4'�����yUU(�]A�Rʾ��.>x�E��u��ڥ�}��JWV+�:�����=ķ6.���]J�eB+�a���N�q�.��y�ۘR���w3jY�yt�#�&�Z��"��C�� b湳v/���hMGun�v�IO3iÌ��գ}�z��|��x�z��?BhX�"E"@�
ZX��ef�ǎ�y��%��>���Ϛ)��0���@������4;�|���}��}�EQ:�0�k���j����骑v�*�^WcB��u�R�Eח����p����I`᫁t�	L��xc�\-V��dv۞[��ަ�6F V��.5.�4z�H}�UZ�	�tǴ�lg�vjLo	f�}d��0_���������cȞ�`�y�m�/�Ln�ap�:D����d���Nx�78QO�WZ�6�`���[���f<���Su����f�&�e��&}�-A�t�h^�����蠱�4��ý�$� ���[����'K�[4�C?�
�R�0&�n�'�3IY���
ض�^�TI�Y�}�Um0"�3��&�[��9VPy	��o� �(��v�<�C�C�`��Y��
�~Yzz��h����&���bMn�����(���@m�& w��0�y�O��cZջu�d���* �s׭E#s��9�L!�����KvS=5/1�>@�`gc����1��q�ʗj'��b�h�6t�^��|�9B�)�q[���-�Ūo]�-6X���\��c��/��z����&�7Ǒ&�%{ܻ�Y��_k��R���S[�L��R����	����@�n�l={,�2V����r
N�x*�����wP5�Sν;A�ٌd�m��/f[tw\����Cv�(~{�@0������- L�@��R�_~IrIƸY:�[�s��m��lβm�L�-`9�I�S�M�+s�̹A��k�4��C;$���ꭝѾ���2� �F�#��E8��9�3!y˴� K��O,u���t�.�YQv���B�.�]!�	�،�M��س2���7qRW6��V��0��\���0��sGTJ{YD�c���AD�~*8�Q���orc��M��-��sf��a���(�ΰᛨ��zru�WK�5Z�."���_ui�i��]E3?{l�-��"&.l-3L�J��ss�yV^�$Ф8��������#��kd�,�9�C�@���0f�X������V�~�k]Lŧ2����[�N���ק��Ƥ��Ǧ8`i`٫9�7Y^xT�n\pm<
�
���m� J�I՛�b�+`�g���><��,Зn�a�M*��,���;.�,�嬸=�:V�M�[�0�v��W+d;��78\V��e%X�;f�Kv���j\���<�ONL>�}�g�%�g�g�R�6�d_��>���4�]��^5��]��z�%��W�ܳqq�Xu1N�%|n�^��Z�B���N�薑Ǵ�p���Q�{:1e.�,�
���>�x�F%�Ք���}Ӊ�N�)֜t���f��%Ѱ��S�Z���3��yv9�����o7z�ʆ�s������u�� I`i* ��"�b$�����}|�4�\a0�]��A��H�TS���'6z�Zj}`���qP��퐦���1e��C�ұR�ik	��g��*dp@��U����a=0�u��9OmzL#��F��N4��t�֩�L�u�T��;P�Ҳl�	[b��$M7�eD?4��V�����	L9�4ۘ�Zŗ[� �+`[��.�{=�O<���n9[�-M����,Y�X�|Eԯ6`��ݮ�~.v�l�2dD3���j����0�����3�w8�6�F�$�W��v��Ɇ���Z���YX]����I6���	�7a�:v�ˎ�EK{��V�9�uk_dFS8e���΄[R�l�r{]X56�@����-�)��}�����Ŵ&Y^S=	��]�&�gǌ�A�%�sJ�vO)��j�n�˨�H\�]�E�����m����9�~Ab�d�j��σ=�����Y ��	pJ�Oa���u#��tcs�M5���r2�&�օ�㥣�H�	��H��ܦ!�{6�[Je�&6RQ��c-+Z��Xze>e�b�&i��9H?"W=��J���j�1�}�@����i{�m>|И6�c)�[�Ja�g����G��p}׻�wv�oZ���Xr������s.Y]�iv�ke=D<��+�}��E�\�ow��:�u!�d��9������u�k��v;����Q� ����3 ���ČT3D�ϋ�w>.��_>���Xf�p`7Ϻa��)���Ȗ���c��זW�U�
����Qe�y9�k%�C����H��`L���E�x�S[�����O� �f=q�<������]�Œ�7�X�u��!G�l�'Z+'̙�ϲ
le��!�qxK־3c�k"��H]c����B����5�jn�y�c7 X�5)�k�b�w-Y �6C(- J�-d���B���g'Y�x�'gt��75{�˷T�[/����r� �}�<k
%ڨ�1���j�0�tS���=Ʀ)xd&�q��Q���|ZfUCP��N�C�J���[a�A��O	Y�gL�7S�rB�y)�Iy{q���
�2^eV�FV��w.f�ҡ��+,���^��UB��F���7k�wB1�M�M��⨄�!8�(J�38򦱖���dBǆ�e`�Qh�B%sSR�YT�d�k]��w��nTL=��p3D�] �&�[ ���3������n�ٷ�[Ί�.��˗���k����UFg�˱��%�/�W��\�,��wsL==w�1��4�D���W�����������ת1�ד,��v�Xۭt��kR㖛�R��m�+XQ86���V;��Zt�m*\�8�:�ƆW&KnFp�좋���s�X�L6y���;r�}���X#\\�T�jRe�K��\��ز����+����" *�Ŝ{�¹4��a��y��9�]�S�|��"�OE0���Hх�-T��A���ن�[F\����5��\6��Ƴ^��;_rTZǜ�EC'����K�X��Z��g`�E)R�V�f�ٲ0�����hlg��̅�YegBh��]`�܌_J�n�u��ʷu��ES��GC�$�����"� Eq�V��b��e��Q��\���{M���VΕΣ*��h�F8������gD�z��-i��8<����0���faCl	YP'%��ۼ)S]	oB+��wb�:c�ٯ�r�y�ڎ2�?WQy�X�]1l��57;�7A[�*.�JݹF�J�����K�[PzF�U:��Y@���8*$@�'~
�~rZr��.�F"ϧ[��ʦBC�~���]��6�9�;<^2��I�î�l�cAΚ�M�(khcهdN�u����~~ypXɎ3�7l
� ��ٷ�͊')���`(�CPK%1ԡ6��5�4�E-�kf�)��OiD�1fA�A�Z��t���heU:v�V��Do?3Q����e=�.���M[M�O�?�$j�nU]����*�Թy��\��	�m�9w�bV���>t�Q�4W1����ݥ�n���S�2�o���';��Xm�������:�й�-˰����k�,��Ώ���%�u�|x�2�-�����}]��b�w<��YW����¾�T!���"!���y�������.vo�t�b�Թ�>k�*�N���]��6������~�������y�ʛ���Q��x��Z���xi�C�:O�@m�"<�;.*a�KC\�Dw(Wl^��M�gFM���jX!�'u�� ܌	�7#z�E�)`��ug�#
�d��eY��H~��◽Э�y��U�\P��G$a}kj���r���J[Ә���yڋf�*���&��*����j�]��m�4��X��I��̤���O�61[5�B�e�vi�8G-�*�QG��>��(��YYN~����� �/��i���J^��.��S9��ӻ�nΚ�o(i��|{˻+�+��8��xt3����1�P�2��ǣ(�����m��C����Fy�K�T�>NԪ�{�����8�5�ܶ��\���,Ŗ&�%������,�74a��\s�(0�ɝ���COT!K�OC�7=�{ukwP:���s,m��.H�gn�|ks ���]�~䗤�Qũ��w�_�G�z�9`�b�C������n���Fu��iF�z��1�h0a�ș�Y����ύ�txh-�#�f�VɊ��*g}��m�M�/o�g7��m��j'l<F�J�9��n�v7@aͺK�}K&^n�d�C�PN�$*�X��Mg$s���o��bY{X
�
�(��׃i#t1q��fǜ�G�Ot��E30��:�,f3�@��W���꿯�`�y�y�x3I�:Zy+v�E�7��)<C�ڊe��[�I�cR�֣��U6�cˡ.�L%�u�oUv�l��������
Ϭ�iȕͯ��X��}����݌jDҢ�P�:���=�a�=���n��|6�,t�(�6��G��iA�L�-�ӝю�u���Q���������udE3�� 縪xmQv�?���O�_j灵\D��͏,� �c��5�C=Xŏω�j����{��ڋ@��)V0j�%�'6z%�
�5o8;��گ�b�}=��b;y�H	>6��ڦ����ڎ��՜<��Q �ق����]5g'��Y
��L��u=�)���M � �LD�^%T��i�V@M�VP�{��U{TC⤯L�a���t��
I��M�0��T�0�c<F�z�{Yn.�m��H�4�lb�om�z3p5�W���t���ȅ<�Yp\�$�9� &������ܝ�@!�Z���K��;Llؓ�E�j��s�z�ڹ�}@�7Q��
�>ڑc5��Ї��p�&e�t3�n@,<�s�>fw]B�fH��q��f5�\�#B%a+��g���{�P�2��2������)�.�.���%vc��ߠr���Z�(�I��L$��t�}[�c�*�d�:���X��˷3�&^���Z�a}b�LqXx�&���e*����R\���>0�0�L�#[���D�,-.�,J�mUo��m����h�i���khX���1[Rxr̢�%�3]͎�	�*���'汪9�����r�q_��_^k �q�{a\^l\��!9�9��n�v*���b��qn9�s�y� v=648I�Z�4�w:�Ne�z�-�K����E��'Z�T�mb���5*�#n(�%ܶ0PZ������0�6&�lt�j�����٨�{#�iv|<�Ml�^D��3�q��Z�C�j����r\��/g�Ұ����޿s��@��`���0-����r�!�^�y.n}�V�9�=X�t԰~�5�W��Lr�½�s��[�N�4�|��g��H�yTs�V�f\�V��H�x̛�ƌʬ�����hy��a�f"˽ OP�@��0�])�DgB��?/�_?��n_�|��٨���./��͇m�vC�}�r[i�7Yw)�	ԏQ6�e�C��mM2����ȕ����8��yC�l�!�U$YU��e�����Kh���tl��?����|>_/��{{f~U��ؗ�ӗ½Fa6�j��[�`�}w��\�]��r�H�fsW%u'�{(D��,.tfv��֩q�[�e��C���3�7W���m^*s �r�V$��1KUԹ%��[DwB+����De����|"`�=7{ %q
��D܎���ww�3�s��h���7C������� *�(C�w9)����;��F�]Y�F<,o�ǴD.� �t����)՞רn�[���}I�N�ٸ�U��!�Ti%���6�F�C��%��6�n��f��Mt�'��v�ا@��kQ+�.$s�)��xJ[�`��Sz}F�>�N��q]�u�u�W�W2��\,{�g�߷D��k��c0�m�-T�=k�w[�.ܸ�5����;t�3|�ӏ� ���@vؼ�6A�;��\����:\]�#l틮��S��FK���aC*k��Ab�y�J�ǸD��[�EKr�3���g^#��r��]"	���+2���Ұ\��+q�G�J#�`��W�X,�o�&��:s���0k�kiuKQ&������}�,�Q���z�]eXJVp�&*�����(�X��%n��Q����=��]��6�m� <����Z�8�ep��{Wxi��!8�5*���mĆ���Nn�qK��X�pm���ve-W�.Z��=˳�qg=�Iƶ��WG������m�Ti,�ŋ�Q�t����Z��������fGV1f����Z"���}�.����O�7�k{1��9a�ʉ�����un:��**���w��`	,]��re��1������g@��Y�E������oj7X�Uӻ|S��Edm����;FgqI��b<�c|FZ �����!�%GA�^���5�pZ��V������J�h��@�|���6
�̚B�[�/�Na��p�&D5_.-��	����an�v�҅�@.�!�fU���ZcNp���ܙbە��.�� �2��}.k�7iθK9�/����F���A
1F���ޒ�m�Sv$��}�εՅIf��%*w>2o�6����m_��3�Y�"��`%����������f��\Ϸ��X�K�}]dji8��άSm��jG�bp`b-�n���CR��V҇�{R�(m՞��v���Y5�6v�?�Q��ʅ1h�]��{u�1���ï$�R={w6�NصkaΫ��n�������I3`�<��ޜ	�|�t����n���9��u��T��OJu�����\���jH�T'o4싗��%;��h�ʅ�c+�-'�k@����5�O��췫L�N�s�5���cj�ћY��7;�a���Z-l8��2��*^p��)�l\�h+o�,EM�w���)A{P��B�������F^�t�4����2	J6Yn*����P >#�� ��j��-m�Z4h�����
u��%METTQ6��PAtkDd���`ѣTM1QV�E�PEU�j��KmP�έ����"��614�I�����1DTI[h������j
i�ccD��DEPSDQEm��PT�LE4�U5�UUU[j`�"� ��k����@j�B��֢�+lP�V�Ѣ#A����(��b� ��UQUEDQUEU�Tk	F٢�
((*���f�"��b��QTET@D��-��v�1AkV�EE�[����&��F3���������-8��ED�ţIM5MZ�TQ�U6�kS�4փDDEUDQIQRձ�!��4�Mi�%T�LEPm`�TS��Rf�*��$�h�m-��+�r���8�xTSM�j�B_B��Nm)�R����1o`�7�x��Xв$���J&��R�h~{� <����.x{:y�7_�²��8�^y��>Ȓ�f�t�W���$�L���+"��C'�4E��m[R*�������zw�����i�h��f�:�`l�~��ĝ�e;�k:�'��k+��ٶ{\�ND�6 re���-vUl<�0��!�����#�ݮ���3�h"�e�%�Sf��]t�x8����'��)9�n;����@�oO�G�χ{
�\W���S�
���pئ	�ׂ�*�k�6E�
y=�(���ڨ���a��ⶶ�{�㡷ܵ��`Ȝ��ڋm>�B��ڸ,�{���݉Qcp�*/������^��m��Q���IuGV=i�۔�C/i�}@4F@V)������ɴ�yv��UM�5�	���sE�$k%��pil��:ƥ�e����=ql>�q��s
Eq͑+++����Z�x�k��|2�m��F�6r&sN>��\u{��&�[�8�@O��}`��x�>�pc,�i)t��J��y��x����ܡH.TXn(�t�,��]Tc@�sL|���|�Ig���ƻq����������
�l���k{㿄��p|�Y
���-m��*�]^+c���\S��5�P��e��ƆWm��Ug���GU�W.�j�n?rv:��>m�j�6F<w|�^gfL�[6t�}5�1�8�T^�d�\*�1WJ�%���N�a����[y�\���efu���| ���%�R3�G��<�l��s:�n$hcP��hSZ�L`g/@��ffͱ�&�咨��飢"�c�[�2�2���v?�P��M�N�\��3���R�"���q�p�v�;aĻ�1YZM���I)1'�;8,��:P@�oE�M�v�^̭�l���I��o��'h�=IWkgLM�K����e1���&�<\+(�.V�{�Tڌ���g��Ӗ~s;�)fwz�]��3�����2Zs��l=3-ɂ�f�sя�t�(Ρ1�K�Ǒ�" �q�u��P�x`gR�u\G<�wAt`n�E@6���|�I�;T��Ú;��᷐�"��ʣs��>�@U�v�켘].�֦�Nlz�Kը��ee�«Z��n�H�$~젰f~���~�����8}�]�|'��|u�Mxy����f�P�R���� Qk��8�K����Ϝ�<|��2����D���5(�-ѝF�'�J|��V/^dQ�k�#1�K��FMv��3�븷4�HM^2��u0�ݑHhg��̽y˴�ԻO0�e������.Ů"�!D`q��Y�[�3�����Y��p*,�/�me�'zؾ��!�zo������2�ń6��%a� �T{d������_3:un0�[N����Һ���������ڻ�;��_:Y2dDs��5(֕ڮ�XgS�CyV;b������\-�c�7b��:ڨ�ίgޜۑ��;�0�F�L��v�:0��	�:��k|��+��_��X�ܭ`�5T��|QR�x��	OQ��^�,�w��c͔�lӐ���0Dj��w�o[NU�~2xVqB edqG-W0�2X�c<�@[l��͡م���0�[{��+)k��k若���Lŧ[Q�ќhU{��R�oN�X��-(�	k���s0m�|[Ƌ�z�a-V��T�s�<��<KA�<yӲ!���'^H�c�����mj~gm�ָ�;�����������k~�mYaJ��dgN���Ց��$*���y���*�V�E:��ֵ��v��0�`M��p��V�E����C�d�m5���2Z�m2챵�$�7��=7��'�U&��wT�Y�˿��a�����)�nn.�V�JĬ�[b2���f�O�ȶ�/�y;.��h9E0m1@4]0���m���Skk1�Tˬ�w4��ME��ʌc[���G�����k������$�E�brϤz��[']#��!�/
��qwKGnH�Ɓ���7K�G�l��W׹�B�`C5L�wK�a�8Q���V4�{{n��^sG<Rzút�
;L�Kr���롽0�6]���rJR������+�L,��/��s�F"w���\�N��z��~�3���#*KC�1��*���i�V@-��P�}V�$�vN�2񗵒-2��\�z��2���)hr:�k��^�<Z ��W���>R�c����g�N�q��{z��R������F�z�hv���h�,�sI���p�H끧���{�mjq(�f��ͺ��e�sJ�cy�l��'4��i�^�-P�n�t6B��� ���]�3UL�t}[���~`��-݁*��]�y�	�l����� E�$��K�t��'�7��w_��� ���;�"ጩ)�u�����y�N6�5أ�.[ɛ��\�(K2�iZS3��Z!����QO�BL6��dK�b�oO�	�^%W'�PK���w=.�nn͑�J�Ɩ�|k��+���;:�8GG�`��^D$ԅ�F����Bi��8%݊!�0�^�2�;�齲mﱉ�iև-����.Z�s#�n���cO4y����٦�׾6�jYB�Ag�:��EU�!a���5y�>�E4�H�F����-��U�~�i�F8诗�+|2��ƤN_�V�5��<yo3�U�-�B���^ͫ�{���z]�l{��Y4ڙj��m�,��Eu\��B���i\
�1kh���uk�_����Ү�b���)��7�<�(2�f��\8\�;m ξ\��˺����m�}�v�{�78��l���-��8s8��X��H�[���hY����EDvyo�ew�f��s�i�6���Z���X�}�GHbdckX���7Y�z���;G��O�H��E��"]��cDA9�Šg[;w��ր��Ǌ,��e܂�fm�l�.#�n@�d,.�8A:���&�nEA�+�"�y=��K�1h��h�>����l���Uw���h��U�Y�4:�f�B���s�Z�=��g
/�V[8i��B��i���o��0%԰�ܣѕ���[&�9��k�O(�5lѶjV�.�+����v𽷒�&tǜ�,7��{P '��BUjG��ts%
(�����qە��(S��X/��,�n�VֵߗN�v����e��B���Ij�yn{����Xf��)����Ll�,W\��Fī{�c��|W�p���ʨ���Y6�*ܷDK���i�=%�=��/+��n��k!Z��V.��$b��g����q�XShͥNdKf�����p���zro+/�Ӫĺw�~�e��t�/���^�
D���_vҠK��a꥘�6cr|�E�E�w��7L��f>�>�t^h��v:p�Be�CJk�R�K?me0���VVy*a��r����^-�}5�Ǝ����f��3J��a9����q�p�f	S�.���=#m�g���]B����2v����{��rށa��7R��:���V�GH|7��;��a����M�-�S�C�ܢ�cĻD�}ΫiS̓��+�/ܟ��ݩސ��K������ew��j���Π�����0���Y��ӯtz]j�M%��,�Ϡ�x&�[�%�?yW��O��H�(���5����{'��J�F���]��i�f�6'��g�4�W5y.q1���#��Z�r�/3�o�3Y1�Q�e����>���cO>vW`���o�Ա�C�yUV��W��`��:��<ѪS���3�c�o��%�5��l@/G�<��k�T/k�mC\1N�u;0�8\�e��=����v¹ъ\s��Q9lCY�!����ͽt���N]��4�9�^t��ɢ�RD�q�&�E�5>�p��*����8�W�]BW�����x)��w�����1<����#cE�G%n3��Q���	h�i�WN��*gG��ӕe�&<�o�-������]+3�`2��UC�YK�P�r#Zj�Q%ڤ���r�o��n�q,<��)��j9�wt�j�&�����dܮf�t�
����-����2Y�����SU{H`���Ë㶟7�wV�j���aK�,K^�]v�[2��v�'N�\��b�o;�͖����]��9W@B���u��F"sC��� ����͇��0)�?�*��4mo�r��F[ȹ�a=�N�����֢�핔+oÕc
j�b}���Y�{��E��H�LCg3�b��y�e��a'���@GD�|g<\Jg�QI��e�*�\]��0�]n+�՝y	�/Uò����zk��$�,
r̤,�b�#��f1�p*|�IK��۬��i����{"��K2�Xθ6`Q�Bf� V�4c��nodS���C4�yJ/��ք��^�U�e�4y��c�	���Q���3q?6[�w�<Y��مI\xu��d(Takm��h�rI��#R�����2<�Kj}�;�ό�x�ޛ "��"w;��5R'e��:��/����V���G��5h��Ot�kwY|`��1���$S5�QY<�M���{��p_5�t�����Ί�����6.��P�oS��,��r���}w��g�\U*�i�s�X70F��Xv4���>a����TS)�ްJ�iOE�Y�k�{� \#�n���6,�jZY,�g��`�l�k/㚁^k~`���m9�ͱ�ь~�{��p����������"�)�9dZ�K!wt���{ Q�9��X�bÊ<��U���7ub���0c���
R�~�W�-�0ZG�ʝKQ3iT\�gL����d��F�d�5,�iN�87���6s�:����^�����]a�vI�>5)�@]ǩ�C��������j���s��~;A�T�&�}�~;{U��Z�7��CH��J�=���u�K���8�h�8���"�l�:ϡ�s>�`i*�57,Y��D{a�ȉ�8\OaE�(��*"�֘/y�M�3fd�O�`�~{ ��Z�*m�H�6П��}u�� &�^6Ft�b�h��ة�I����騵��ls'*�[@�,a�A�BD�U��ѩv�M�,E��o�m��G~��Ly��lJ����L��4ĥ-1�ވki�й��:��ߙ��|'���uǨ�V@��Wz���`�fiii=�Z r2�s��^-��Sm�����7%<�9MƵr��ɚ; �����T�����I�o� 樠L4���i����״y7)�i�ܕ=�onu��3<�s�U2os�ۨZ���fD
��W��r�0.w��덖d�t��d�ޜ�7*��(U��R�^S�	L���n�,���iI4ѤK��.\h�:�1��_TA־���Z,>6���xb�׸�.ʞ/�l�6'��I�ְ�H�g��4,�˿	u�Y���Cj�_	�\���b�b$vwZő�YI��ŝ���Ƀ�m��y{t�6v)-*�@�gׇ�gٷ��H�-qs,̗�k�-���˒Z����'�R�7��U�
�,�|���:JY7����Ͼ��*�~���Z�|��i�+v��N���7�7J>%V��. �\C���Hm|�94n�U�-�<욚�<��c�F�a <Bm�mصE��љA���:�m�'��\�e����'�D�kۅ
H:�.�Y�3B׃>�p_�Ϛag�Ml�_U��8�a�bʅD��b�}C�3܅u�ЇdE�{8R-��v��;�g�y�P)��L"�kMz��
$l��Q�9��ɦ�7j=�R��}�7�����!J6<��'Z[;;���c��x�"�E�!|�k�@���� �ס������&F�5��Yw'�`��.��3���v�MI4sE��V�;3���,�y�1���d��c�$���w�n,�4���RUD�5��܏p�ʕzwll�:m��n<錖����x�=6�?��e'k�͂�EJ������缉iREE���nL�ۯ��+���	��
���=�'�5�t.&�uJk՛0W3.�[;0ͱ���O[5�nyC��mz&�5d��[�w�DΚsTW?&8������ק����J������pue(q,���Ѽ��y�sޝN�=�J����U��QK�`�޽c���`����i�Xg#�<#�w�^�;�%=]�K�0�u�YO�����������z�Է/��>��j﫻YN��0:�͚�s�L��yh3ʉ�}+��x^<�� 4����[����D�{;2j���M��U6��ƚ[8�l�{k�e��kr��L����~���(�]�9�n��|�X��)ֹ�fӬ������4J<���\�T�ȍhl�&�C���}e�ޖn��pk��]B��g�����+�Ԫ�c?#��޵OuV��k��I�sR}1�^� �̼t����5�X�rRZ��\���}ސ�����S#g��[�hU:\���7P�O@�����/�����^]���!u�	�[���9ݜY;���r!�7����B%�#[hnF�q��cl)��ƻÈ��ڭ��]ʊ�z�Fz��̦Q��}xul�|dwj��mG��2Ij&�e��t&�Pm��q{�ᒸ�܉QYQ׌�f���a�8�Y�&sz9�ȮXǌ�^W?y��j8�@i��, ��c�{������L���VE���X�z����0Sϳ����c����5=!��Uk�1���w���,�O]x�롗0kffe�cId{V4Q�O���#tσ���iy�c۫X]�Ǜ����<�����^�p�{|�o//fx�fڙ���
	�R���bx����)��+e��[s�^nS�=z�*�J#��D��8�OhQ�̾�a��ޡ�Xz�p{e���b�KU��È񝥚ظMwB�9���$Z�k�$��=g���#�YFb^�{r@ �p�������ad�v,_qq��n���(��6�f�e�F�|�:�-p��;j�b��h*��9MoiN)3��(�㮯]��{��3�1���7`f��m��X�Vє�9�с���Ƴ+t70����1��^UŶ�/yeܮ�����]?6���z��_eԘj�Բ��!�/E��O���͜oU>e�R���:�7f��*�iͺ�N��w^�9����W�ք�ԛKKSв��9���Ǝ
��e>u�4��!2��X�Le�:�R�eQ�{"&�qw
�Z�N�we;J6)��ams��	W��P���t#�b'Ϻ'����E�ϐݞƎz�Z�1ޕ�������^�x��
����ͯMӽ]*�:�����Xl-��G֒u����:�d�)�:΄:�8$�m�wv�R��Fn�B�4�&t��ѭf��i�C�kl�]���"���G䈮���_w(����C��7g|���,E��xjs������vV�Rt�����]d}(=���$�ޟ>��� o3&����/ ��0�k���Q�F�۵�M�R5א�3�*�K����C-dǝg�t������HB��tبjt�$�rj�L�o2'�4A4�TG� GD�M����Eݱ�b��7��8:iO^)��t<e=��pXt��&�%�XB�
���ˤ${RLr4����w/�{��/>����-;�FʾA�ش7��J���O�gq�Y�����q���d�k�ds]Y՗Z+4s�+wB��g�%�m���9;Ϲ��J�*�"R�rǶ���%�u-2X�����/MG�V�Cisg�n���K�[����t�t���)f� ���]�}���B����{Eh:�ouAe1�m�%�����"}��4N�VE=5���V�>S�{Q���]uh�4���1b��ݽF��]a �Aл4���f�D�gQb��ӑ�.�.ۭ��
Q�)�.l.$Ï+�`��S�ihf"��Y6����]vZÔ�����)�/%�[�`� �<U��b6z�>��:r���8j'w� ��tA� _c�\V�Xydf1ܟv٩����
���A}���΢��O_q�8�I���j	�W���*Q_n=�s���gS,�E�0��f���A�^DV���'� �{�r�����i;<n�e����x�e���M�O)]�G-;�SZ��k���q������l�ur�t�&$yAe�+-�����*�4ˑ_^S�R@d�q�Zu&��[����b65�h�,]��t�Z�u��:���N���n��F��X�4�QN	*|eB������TZ���Ԅ�(
 |(R'�֐��
*�lU$UNت�
"�*""��lo��Zi�+Z!�j�fI������h��)`��E�b
)h�
i��"v(�Ѕ�P�Qm�Ѧ���`�5�4S��"��(�`��(������@F�I�Q�PDSCN6��j��1E��QME�UUZ�T�TDScX֒"&����	+k)� ��
+A�lX� +F&�	�.�sgX$��IQƢ���������)f�Jtf���-.�������MV�=l�6c`�؊KY�)����"֊J
*-�KA����"lQƊJtb�Em��$m��"$���6���N��5�j������E�����*�>��$�Yro)~�]o�A]Z���Ug
�@���uc���k�d�h娧ZO3�
��V�N��b��5K�h (�D�;��)چ��~|���rol�k/�8{y�����[l]�M�'3��+&�I��8�0O�Z� /ekA׆<`aD�ǋ�e�.V�z�T���y�4�3��l�t�V8���{�γ�F6=�u����g��nWG�TO��(�%�����-���d6�_2��D[w�\Z���FE��V��n��T_*$�ڗ��6"h�>���av;��ڿEE�1vj=���bk)����t���vB���zl�+��m���%�2꣌q|v�f{�Vh�Y�k�ܟ#�.�AAO"�[��56�E�(��x���6�����5�=Z�E8�m;	��#�PV>[���~����M��-a�Jd��L��kb�0UFdgUA���E�����p��i����#F���Hhi�p͔�8�����g�]No=��K��Γ<�x�J}���7�7�Gx���,�?��(z�q��6�2�
!U���Nx��V�A�m�Yafa0=��Z�<sm�Æ:ȜR��d*�\��y�=a���tqu![���Sp��ͼ���C{v�{s�lU��Ւ������+<C̉GNz ,�}\�£���\C�@U�|U��Q�<���v�J��_t�e�S-m<��r�p\2+�7o�_*��zJxo�~�ֱ�bR#�ɓyo+�r�����.���N���W�����[0����������� ��2Y,�ѮaI���]�=����UjM�Ls��D�Y�e��1	�T���G�g|U(q�����Y�2�RXe���۷u"��,�¥�=���kp�<9ك1�o	k�!�POE��p��bQ�q��mY+Z���\�sq����w�"��1�,5��-���<��m9���,k�ʝ7q��g�L���8L)�cZމ�hǠd~���4��"4��!�I�����i��ǐ��h��ڜ[��-m-	j�����8�g�0!��T����wU�,������k���@��p�����G��k"���ݾq8g_���ԌT��Sm	��z���Wg�[��S��lF���������9����<��˻�Ő�}mF7�pl�l ��I �1��Yؠ��֋&�*z)���I�eG���|o�4���L"/�d�QM���[�M*�&��t�g6��u5�=�#�ψT�;�d"�S���	�@�ids�,Xbc�����1tS{���鬳s�H�6'�)>���۬�o���2�}���h'2�S��q�w9�qS��y���K犮��P������Hl��%v���ﯥa6��G]!�R�%y[զ�>s���.�b�8�e
׶{���V)��
{6���?��GN<D�]� m^������@!�SZ:��Z�ܕ9�2�)s�<��	�ߊ�d�橶ڵ��)(̈y :Xhs��g��Hk�Y�y�)������n�t�u��H��LI��U%��U��:��Sy.'^6��3=�FwŬ]�3�ö4 �چ@M�b���(���q|��ת9������:��9Y��r&3��=rGC9�s�����;�h\�g"�7!�����׀�7z3��Ϻs����\^p�S��gB��f~x�cp��Y��PA����6�e�6ױIjj�5+�j�cJʉRF���g#�!P���NYcT;a�׈�s#�i�Vh�)��;j�=镍=�hoF⪹�Lp���]%�(,�;R3:�H�v40nc Df�����/T"����4���@�e2g{�A='��]C��#�q�g��DeS^��)�֏��,׭[�h�68�؊Ue���b3�9�N��5�L
�4v3��ۨS[H��	��,-J4�:��19B��cz��c��q�ن�\��`�z��_]n�I�p�4����wn�m��
�{(Rx�m4���G��N[9�
��5cHx�Ʒ�}/M��޼]�*k�c��6�mR��׮=cB��+it���<�����v^���	B�B��1hA��?b�g�.��h�l=���g�A- ��:�GbR�vgjr4h��=�ȃF,�m���5�c\]��#Vqtm�hTG��MDKM�'m�CP�`�Q�٧�����j�JɘS/f�4v�C�2K�y��P6�c#К�u[�0'���E�����k���=�_{�d7=�FK6� ��6_��PX/u��u��/�<樣���zBh����!K(��/(6�3�����Ӎ����Uw6$���E(�M�	ʦ��[4]��5&���A`���cAwv��n����o�����"ۄ��m̊N��TRs��SooU���N�CF���=њK�j�G��mR��n?��<º���ʣπ%����x�n�;T�TQ{����cw+�l���-4�R� �U�?uQp
�_7���\.1��p�¶�Y�σQ|�����ܨ"��ht*���vW�#��.z�ld$�s!s� [spo;_!����׹�,���\��:�r1�tƶ׊9`߂q���9���`s<sH�+��;g1^B1��؍����u]]�������K�9<u��3����U��� ׹�������W�XsW�w�x;";۫P�x��w�TFf��1� ^ L�S���ݴ6��=�����>��*���W{������C��K5��Z��9�c Ơ5+f��r�xYf��">N��"���eמ����~*E1�_�\���6�1�G��(Ni@ݤ����p����-ǁ�^­���gF�;�Dŝo���qG3�#�k��N[z��1�{g�����d10*܎i��:���J,�6G3�vN��-�<�����u8�d�i�c�Z���Й,`-\���c��9�P����X6335/1�%��jքQ�kװ/�c#��#+Kԓl��A=z���K�v��a�Jh�0��M�e�8,�����޺L�ۗkʪ���n�q�����j��i�	�����3��Z�.�\��1�Q7�\++ƵAr�蘶��&`���\��F�v��fjYx'��&d�^y�j�g�Sp��5�*��BF��v�u�"'e[���k��=�bH�����C�]?�`o?��&��TI]�Iv@d9���T��Vʯ:Z��־�^�L	w�.'�?A�O$��1㔺�4�53Gʻ�wF�Ms�d�֊�����#�]�l9n��=5/1�>@�b=��J�����Z��u��m��*Z[]�Lْ=��򎰪��l�]��uS���f5�AkRD�>��.K���S��=�~]!in�������D�u;���VY�G�Sw;i��A��ޡxxł ��pgi�β��O{dy�2�U�G�:����ַvᬒ�[���v���T~�}6͕O8�|EE��]}��^݁�]��W��zc�[��}��^/ ����t���<�+܇�LI�p-���9O�61X�z���a���c븦F\8��hߑ��r�Pf�;M���]Y�+�m�^VM�̀\�'�3(���)��ܽ};1�z�%���`�r���y�s&�ݦ5�7`�cK��u��ǀh�`L�m�F*S#�tO6�
�h��ѷ�6����|�����{�f��EK]Ln/X�����4���6eŝ�\��2Y&1�;���>���:��yW5h�b�뀱�ن� �ʄ�s�DLe��zh��Ը�����u�q��Ai7t��.s!�z�u�J<`a`��1�����	=��Sub��oO�o�P���?]��fU]���B�ld/#�u�U�����@�U-#��φ�ʎ����2N��`ڔ����i�|�̵E���y�Vz�#���W*|_��k.{Pu�j��a�B�m�wY82��9�Y3�0H:e"�:ݫ�-g�/����f��h;)���b�.v ��P �/c�Md���s�j�{ {�m��)�iZi����4��u.��n����9��ƆnR���0e�J���*I��n`d��x�2�w:�F��]���#T�vU�-?�R:�*���ڔ�j��"]׆M��]�|�;������+�N��ӕ��P�I�B�K��E����Y]�q8t�W��P@o)`�g)g���wC�h�	��v�`h��b�}�&2��G;ʣ���������,e�A���P���Es�B�\�YD�댊�W���V8
��p<>��sMT�7W��T�ݤBi~��;�;`�s�����\ba����g�$]}���-,�r��!a�#z�N��k��/j)�6���>5+��\nl���2���M2���EfX�v�E�g�=�ĵP�a|3�۳�^�%�A㕿���ۣU��$A\�؞a��bS 1��1M��V0I��z�TPw�`��L5�.�і'%�^�׆9n$l<��������� ��ӑm��kh�I������Uxj�{^��#Zb�K��[���&���OEŇ4����*<��S�o0��x�d����;oGo�(�r��?8��/�w�-��V��Sm��a1B(���8�ܔ��h��{����9LF��0��4�%��P@�������x���]tkK{�n��>?v��{t��s�}KZ��T�yf�6OƳ���C�Ӓ�p���;Lj�>�1b��vV%���3m�P��J�7���jtDnr={|�s�b����rQW.�85�4WTC��h	�)@){�^�s.���O8�Y@��:p�.^�>�a������vz����t�),WC�n���;e�n�qa��
��L"��G+���1�ss4�Z�t�nJ-�i+����Y�Rl�H&6A"�ר�z v<�5���\�JG~�����>ӯ�G�����s�U��w^9�|fvA6��i�1���K�Y=|OVT^�ZmH�F}����F���{sh?�o��>���o<����4�u�z�O���`I��se��S����ûwN���Q�9�7qC�!5���:ƽC?���T���;��^�nC�F^p�~������8�������;�d�hF�H�lR�CY��Y}q���B}�,�7�Wuv5��&Uya
'�!�
���l�m�����w��jdװ����w�i��8�W+�'��C����
�%m�W�̥��1��;�!��I �b�c:��Lh.���^�8�1��Kla��,��	fV6u�#���%����1=���ЛmK��"{c.nx���,��I^�h.�������kUo<�𻮯aT�0��=��(%�O���u�-����Ֆ�U&Չ�6���;�>;?ہ���[p�c3��K�*H6�ڽ]/y����j1�W��!~ �F�d6Fm����5-����&���W�pv�P]vh*�����[Q{m���r�>T���P卒�Pl��5��o�Ws^������j�Ø��own�F������k��wG��y@ɵ:�=�d��p��C(�{�g�*�_u���1�^Q޶����ݐQ��<�62�i�,Lwtc������{5ժ�ՔL��M�^�mʾ�ø�W�wV_��Z�"���0z��#�<��w�gʳd���EDn���U��f�qIn̣ʳ"�Go����V�����1d����5���n�	�w:�+��L�ܸ�x�-�yU-ǆ|�,f����NT6�����>��(��F"�Y�8fw~����Z�������-l=C�K5�J�����W��:��լ*���o�@EO�\��Sד�X1����E��;�K��z�Z�Hܥ�{����g���[�S���v2&x*@�q�"b�ږ�z��'#�b|�aĝ����a�Tp��N��p�#v\���[d�@����j i]u�jp�i�wV!�f��c������=C6\%✅����$t�1��ݙ�2�KIڝ�{,D�N��,�z��4>���iUQ�t�"��}pfKϳx�QHd�Z���Ϫ�g&�!�Q��~��?M@�����Ǭ�j��}�_/���G"��)����g��I%M�(���aM�ǵ������֔��j
'�IĜ���[�.�����_1��:�I�k�-ш�hC���I��ү˟_���hɇ��R)qvޖl�ڋ=���(�mR�8�d�Hd�!��^�X����Y��1yk�(0gF�ѻ�%�gbUn#v�xƤ5�$An�cݱ&N�ϯZ;Pab���S\x�\ls�ݿ�U��3Ms�s>g�����"^�I��R��2Wdo=��|q֝�o��M"���ױ�#��B������4���%E^1�-�/��ͭ��b��ه��V�	wW�c�OryUK��	�����htşr��O���^����=�j��R|�ZĀ3�����~�W��������w������W�
Q/S�f��^�r����3)ԝ#�5�ݷ��ɱ�|��G�_%���έm1{�n�BY8����!v]3HM�8��u$�{]�s-���R��#��uyO��kޝى��{�B�ϫg"ڬ�Ⱦ�v�z5fX�ϙ�|�{�J���k�.��V|�)�Wq����2gG7"P��v�l²��q��ed+R�H�Z{»����j�ne[�����%wT�)|�\a����g+��K4;X�,8��:R������[ݫ8�瘂�e (ZN����Dg^�[�%|����jCO�xK5�n>����S��E�g3X*�XnM����f����Ps��������\����]t���vr���=���uf�\�[�+��}ZI�r��<D���3jf`7����LoK�G8�@rY��?��X��unin����&_[{P=�����<��wQAӴi#�I�9P	��U��`ԥ3U�򙖦ֻ�����l�J�ҸK�ƇZT��;��ÏO*�+���[�R;!x&_&�7-L�P�[�����8>���.�9�)�j�9αbx\*��.u 򚺱B��:X��nP-bͳNe7��en��;>ʹ�p���779������,얫l��rIث]��r#Ւq;C��:Uw٪A��%�	��^V�}Yo�Iuy�h�uƫ3��-hOj[��5���C�h����;��/=�jX!io"�@�^qY�p����/xY�#n��k�uHi���ee���b�#2�����ܗkVP�WZ�$��L34+z����G)Y��k��]|K��\�/l]�r%�{�����b�A���-uk�Z@�[O*�dS�4�XcMj�`�gz�5����a�R�z��a��PV����ݻ3��a��./����u�+fF�G�|u֭�ܝ/yn����໻��Dlb�9�cE1���
)�#B�c�_���F���vgr.��;��z\��K�@������`�6�.以h\�ӡ�e6]u�%1kƯUu̾�6a��ė3LF�ή����h����y���)2e��{o���t�U�69�d�V�oD6�:�*�۵q���w�n֤�q\�.=��4�p4,�&�@�Q�%bB��<5ud���4�v��4~޻T�I��7�a.w�"q��-��BG/=��3§"H���e�"�s�p���� �Xb�zk�[��^\U/�Hr�E��6k�����]�eg�'\��ˢ9eb|%��{M�v[�֙��%��Ώ�&k/y`3��u�11)�wX;��m��kR�k�3t�S:���nk�܋j-{׺��E93-��X�gO��L,u��WF�˛������-����}�O�0D
6��v��|�/_Y1�Jo�;�b��`�����Ԙ�L{v�p�E��.wr��_^�IA��&f�u�J]�]�n�\ �F�珀���q�� �i�R�|%j��wì��E�f�sp���iN���a����q���5-��σ����UPTF�$[mi�b
�h:�SED��ئ���FmD�L5�U	�6�%��TP�ت�J�Y�ii�a��Zu���+c6�Bb�:*�h)&4�m�!N�Ӣ(����
&H�j��J�c%$K��4�D:�h�PSĶá�
�����")��ILMS@QZ�DR�j!)���"h������TUQERRALQ�-��SSIEh1)AUM)6���Q1IAEUP�4MPPECM�h
�ZZ(��*��R�ꪐ��#���4(�*)��llF��f��H���gPsj���b��f�(j��h�Zi
(#lWYuT�T�%/*�C�AQ5M#B�ؙhh�@�PRU��|U ��?������<]xb[��Yta�K�n��-�L�s�2�)���]�gR�3mN�i�Y�Ӕ;4S�^���gc��.���F�g�=3���l��`��Dj4*�R���q�5TuCT��\�K���׎��:ӝ3�ܱ�qa��I��f���r&��=��S��荥�����m� 4���al-�e�׈���P%�x�L:��{�j��\O)��0�~��Kq��HcA���߮��&�I��a��j�WY�߯X�S�"l�v7ۼ[�h�f�� X�q����Q۔+r-B�~ʇ�ݒ�ʘĞ,�Wg�'*(f�H.�;&c��SZ��1�[��L6��L�y�#���3�s�)�/��A��+v����C�f�N%��6-�����:@��Heu��2�pܪ^���U�!FgDR���T!4s��\"��� �Z��f��+2��q�*�k�v�K������\By,^/��AIY��pU{�%EJ�x�(�,��v�=c��m�X��OW,�(,�Wn�e�p�+T
x$Gm�q��rh�-'��4cFY�%ݳ���[gt��n1�l�??�7D�Q/����T��bĸ"Wb޹X��ݥv&�ku'S{8�����2�uk�u%����X�luʵ�8T=�k����)6���o�N����k��j�:��[�ť��sʒ�^ӞJ�|��'�uV_:��X4��9X���Pg���pBپPav��(�ǁy6�?���J��E����ަ�5�ͭ��9��]
�.D��8.���� EG߰	��'����?x�grQ�ȧ�'B	ܠVt�fv���Hz�Ƶ�TtM��
d3d�f��u��E�lO#~��%d��K;Lz���7������"������� �\b��*q�s\�O8��E��ly�t08(�19L֭�q���5=�)[f��a�a}z�/�Pi�i6ϴ����F��u�>}f&��Hr�Vn�v-��݇��ZG��m&�?)��}5�Y��V����
j��9fVlA«���r�g��3��z��h�*��]#X#Ma��O1�p?wy:���XG�6��3�Aa�2J�H�I?x���n�RГ����Jm��*��-�Xє�+�(�\��.�c��V�-��X�4v�a�\��Nu�4�u?�B�f�Ѳ�󜠰�ͩQ�P�Ge��5����u
�E��h�ܫ�ncg�P��1�,���\z�y�U�=2`]r����h��b.��ݬI"��aT�h�)቟$5��\	�i:�9ݢ6:з���7����Q�@���L��{�KYjS�f5�*�M�m���5�Z.wҫ�ݧ�n Q�e%s�8��Mm-Q7�oX}/�3KLQ�b��8N��mϛ��B*={�ݰ�=�/uZ��Z��z�U)�"���k���H���5w+����\�������8�Y�64��lن6�CmSOE��y~��f�l�|�ݩl���>���N�=����o ��'�5OW�%��)[�[U��:%>�}>g����T��_f���yZ#���vN��.��+7v;xq:W>삍�m�E`e�Yrt��5�lۜ;|D���ui3��:����f�R�%��ߔzЦ��f�v���m��3�8�R"Ҙ�F��m��V\�|�vѫa�=�V)�ȡWS���Z�d�/"И�Z��*�;rj������xU9���*Y\_l��W�(� i�*�����C6E;�fL)P�.��d���v��"��VI�n��F�"�^���>���w�0����ݘ��79	�V]�z���Հ��ѭ�QD*�"�L[��k�׻��>|�93��wZ�uf�Q���)��1����+Zn#Ͷ2;ڣ�1�y�1X�Ќ�Y}�1�]/خ�4U�?1��-�]�I�^����F��v�/��;�K�%5i~�O���w8��TY�C����ɖ�N�����k.-�M�Q�s"�tM��1w:����5MY�St��I�	+:�G�S:����P�0�X����������:"g2��ѹ��4����n=��ї~�i}���%���r��p�Ќ�v��ت��槫�����.��x��2ܿ�Uw�DVe��j���v?�&�;y����&Uٸ-3�=�d���Db��N�X�����9l��w��`��$YX�n(P�є�M(W���UOJ-���3[�@�D��J�Q�yz�1�al��!fm%�_Q�k"J� ӉO�^^e��Sĥ���-V�j�r�dk"���7�����mƹ̣.;Ƶqw�З`PL�J�(YW;�g3X�3G˦]�uz���|���F��R���|�@���L�v#H���V��owj�˗p��]�W�p/ ���xM����DGG)��%l�g6������i�=ϰ-���65�o34�o:�5wH�㬻F�%@�E_�J�[���ڇ�䍃vm����J	�a��݌y�dG�ެ��?Y���Z�'�?�j��'2�ͻXr��l��[�4[fxCv��a�.��n#U�����Z�P�R^j�=�S��h�~t�X��Sl�̀���o`}O��y���Ga�١������%�Jr��q��fu��kZ�Yڻ��-1�/e���l�SL�x��3_
�9m$��CǨ7im,0쭆�g1���{��[;KtEt�=�MK��,���Nf�E��7(-����c��	����`�sL!هβg<B�c`�}�v'�Ms�ǹ�
��C
៳��99�N�$�f0�o�����5�A*bl�_8�����+�[S��a��@Ds?Ty|�f��������,�y���L�a���v�mz�ҩ������iu	#WGZ�O���݊�����MS" ά%�=�X�+��6Tk^�볐�#�Z"�u�:A�L�2��S�:�f���qF��{�V��`��?:�T3��ɣ�_1 &T��E������96�u�W�p�Ӓ
��j��֩�=i�Q�p:�������Ud�oEos�ӍY\��3�+��:�yI�K�����5�eY!��ͣw��O�~,q�ڃ�k��]���{�-*�jnI��$�o���˻6��;��*$�MB�����Z��W.���W�����U��"���Lc��<�S��U>#�ּ�49�Z�w��.!�ou�d�ю�<�-WU��X���R�+RU��E��7m�3��Z|���*8��s��#g�6Qry�5�v��I}:�b䕙��g�:�D����*�B��A1�qc2��'�8Ԏ��J�����Z�bl��۳qLl���ȴR�[4g`b�c;����[;�|Uɼ~��� #;<Z�/����v����>��xq���f���Uh�h�<c�����N��ۡ�yh_e��4�ʠf�kY����_�Itt5ȳ��V���]VE���96Bqc����+_]������}�[�=�b�U�n�;���j�����lV��K�ǫ��mС@�vo�;��^�Ax ֔��O�Vlal����gY��#&w�S���[�l5�w��n�pϠ_����S��\,9�x�{�׺�_L�ﲸ�4�N^ō�Ŵ�E �"m1�N�K�����cݘ���f0�C-�8�Ki��K����ߜH�*�d]��x�}:�y��q��j/30YNf6��ٽ�+֔��-�$�.t��
�h�)��� ��ٹ�C9Y�-t�Ѳ�62�uьU>�g4�Wb
$$�IQr1S$;e��M:W,5h���L<��1U�hre�Uפ���m��+)+�*����];!�v��U�&�uS�й�D�Id�3��H���SC�-�fN���PZo�2kwk��,�U�P��V�d14�0SEpq8����];�q�g���	�+k$�P�W"��oR9�w%3�t�\Bخ��j��ə����g\K���M)f������pX��3O�öj9��7J�s��*�:����ּ�:V��{f;�����w�$@�5WȻ�Q�,<���*�<�ҳn�2�{����R����C�T��Xz�!��F"pJ�a���ܽ��ɡ���Q�va�S�s�E�-�@1���.-��.��3��d�f�Ƙ`��0�n·�MP�%�� �/�Yڔ��DI��fo[��Ckaj��sY1��덁��a1&�*�J��c�N2�n��T��;U|�ZR�%߭�_�л��9<����Y@Z�3�ov�o�D/��34~ؽ6��3;�j�l�{*��⺣��J���Ov,��7U�筣�E>�\BZ� tΣM�;�`;��<��1S�]"�C;�yD�8�f�a�*=����s[CnZ;ri�5�zxa�E�/��9�Է�X��s<���ϸ3Us��5�c{ ۄb{bݯ�<\ANd�
�5���e�u�9:���]�tPźJAHE�G�������u�^5\i�=�v�d�OEzf�
�E��N�gP�{ʏ��͘�?g����񙚑�����n�1k�N�҅p�.t���B��M$m�������X��z�t#H{}�& �;�7&菺��Ǒ�ܝ�狳[��t4��uj��г)|�Gy7����IM����I�����!�}m�/x$@��~�1_�b��If����kk�,��!C4Ԭu��x�&'^ݶ�{�u�~&���s*ɮ]o*|��c�on3�]֤`��-�9�qo�ܸ��mW�UM��R/p��V�5�fͅ$+�eey�728ὗݓ�z��yU�J�|��ȫc"�o"�k�ђ�3=6�;D5�3^���6Qy��%I�f���Ķ�&��[�Цާ�{ɭ[\Ouig�u�;�<	�Nj�4�%+�1��1n��<5�ڎK�dC��o���"��*�'ѫ{�E��g��J�ܯ���W+f�8�E�=]<�����X��C�z���l�iK�5
�Zk�^�̈�޾Ƚr0��㘲�1�So���y���w��!�l���s���Kryϲ	�ffo+ev�(�R��{ѝ�^hi��̎$#�R��=�=�����Y�k�E����p���7��.��-E�&��n@�x��x\�s��)h��m�;��p�Clxw�j�b�@�]��֊��9�5eeI��T�۶�e*�%�*�q���g 5�X� }����
x1��woR@a&�Ε�x�x$�s<+<�U��9���� �{����:[J�T��5�ʸ!zC�����/H����t��bz���E9�$5���+�D�=m��`����.|����DX��aT������'�.��d��V	��٤����6�g�j�tVDٺ�=wr�*Fh�ti��9+zP+��q�T� �2���!�!;NzE򈞡Ly'1m
"�g>��c[�L��cx���KkltӉ�&ݣ[�3M�Ww	ê+:��)��"��5��ě*���+yK`ޛ[$�W{���mI�Y�ɭ�r5�l��Z8D�2͗</��:�h�KW�9�בp	�]݆.��ȧ��]�1}����n��a�-S� "��pQ���t��:�K�9��;�;��1�v����m�y\�����H�Q��v�ܑ����s���|>������o�3��ǿ<�I��= ���9�!3Ekv�'l���PzAZV���kQ���ݡָkJ����5�<*���m��)�=�B��<W_K�AV61n����e�����GeNB.貒���(e<*��i�;��T"�8�J����$�"y��t���O{��A�K�G*e鳢�m�Ny��㑼YSЈ(�d���)UнW��M�L�Ow���:眫Qr]�<α��3�*��0��`��%M�7��9�`h���XQS����x�N���JV�\S8L��#�M#��m�%*|!�n�X��%YJ�岏LQ����s9ap�T.���c�m]��qd�k��mo�LN�GuȂj/�|{/4b�c���J����;Q	Թ�z������&�-�|�=y��l��w�X�Tܰ7]����'�p��g]dKf^ۃF.,��Pܔ;r�x:���X[�kθ���a!yS�Fvoan�[Sp��Ӆ����׊��hKI��Y��XǳAyS]���zǏ[|��tݔ�>�k��n��#���W����ƚÔ���po2��NF�J�c6zi�;�2��.�\ZC�Ƣ�zr�����b��hͅ�w��8�,p�	n�w#co:��/�7Ҥ��Eu�>7It��Z7'�(.��L��g���P�]rG�ݯ���{��;ܶV�ܤ��Si���=Ld{����p9W
#'Voe��Kl>�����"N����ejj�ݗ��o5]�lӐ�ۭ��1\�.�c���>>�G��w�ܾ�4+�R|a�t����sa�i]-�V\�l!T V|x�#`�t^d�y�e�<)��Vۭǋ���=�>�}�_ݯ���M�aos�p�U�������]�/Mﬀ�kcv]]bX;�(3��G>�N��[�'d����3g8�7J�z�b���[�K{�uE�%����V���dr4�G�M��y	�.٣;sm����b"��}�ż��Ņ� @�������ݰ�{Sw#��X�ߎJwQ	��U���0<=������B��:c��xx$:b�x�`�U�H4o`��n��TܵY��i��X $9�tf�Kƣ�һ{-hѥ��WY��Md�m�u�w��*[Ww�.���2��7^_ufpg����t�Q��~;�#
�oohb�1�"J�8I�ԛ��-T9_sך��z����|��?�C��uXξĊ���K7���v�cv��&r�qa���:_NӲІo�� ��=�y� �wÚ�7|ĭ�h��.��i�+z��,�X�Î(��͢�e�+&�C0V��팉�`�l�y�	�������L�V�ܲ�p�������^���k���.
��K'e��^k��rG�����Cw���ҭ@31l縖�4�@)�~=�Ӭ��Ǧe�jB/��lM��=�8Muw�{i��CZ��X��no�,V:�A��<0�`�n,��a
)&
�$:$��4B4�P�x<p��.s�r蓮�������P�U��&ڒ�l'�ryRDER�QR�m��%��-a���cLMTU�QU5��!PcmTTh�6��4�DR���&
b�*)����tRSI�U�LEP�u��mF�4TAED�4�P���QM�14�F3Z����.����
��Z��T�SD�;����KF9�
J���""��
�i�((9rNu�IG-����h�:�0�T�sh���
�nd��$��͐���IC��I��MMQE%&����JT��-)[���`��CMuj��A��ԚB�S���u�����一������*�����"
*�F��KUO$u��ff�� [�y�����;�yQ	*2��;nof]�{����N ��AV��͒�^�������ūUh�^����o6��ju;)��-ܗv,�Q ��CPd���J���hot��;m�k�e��z�|vz3��/vx���6�R��IK�+���Ɵ��ΡE�;@m���?[������z�|�<��P;:du�+�uA.�O��-�sU��We���t:����NW1���؛W�>��^٣��<a{uZ�k[(ǀ��ys���=�W 5��2%��B�li���-����=p�!9f���Z��_�LXm����ws�.��6�[��ufSE��DM�[(�V�ț�-�&��ݫ"�nbz1y󷢅-��{bD=ur��sT,c�����vχ�"� %JX�)�lR0_=z�n����b��4TՐWfn�`�-/ ���*��#L�Æ(j_p��|�:��^�h�,^�����
+2DM����Z��u���s15p�����#�e�������^I���`'䚸�i\��'c��s�&�5/�P;�u&aH�G48^���P1�����n�cwVl1u;Q�2����`��C6ή�I8N�1�p���K�s9V�E�]�uR����o^y�%Ȼw{S��5��<֓�U��j���&Cҫ�N�q:�h״�N��t=��Y]mT�.�^Խ{�,�ɏHk�cC��B��[��g$z�e�'�u���k�5�9�ms*����N�ŀ�-n��+��ŝV�{���m͢6�*��y���t���hq:j�\ѵ�ݾږ̇)�`���:Ҷ/o$bMD�D��D{2����*��q~���K�Q���47$���:�cP.�>�{Sr�)�Y��b��7��\��W�����A�:�)���ym�S-�)�37o ٔ��<f�cm*�v�U仉�����پ/'{���9¨;A�f�`F+ ��Hߧz��7�[��kf���D�^�׮G�Ќ��~Պ{Z�m����/��p���X���nZc+�lS5+�E��F��6��M�O{L���8����K��M���Q8��P�X�1�5Yr<ޢ{Fk�a*$�E��~���ޖ��|n+VR�p˭�1�R`�3��)����4ɍ�.Vr!�,�OO4q �Ѽ�9�q5��p�����uE>蘮��Ɵc�dd��l�\��Z}h�N-!��|��>������F]���V҈^��\�PӒ�7���ZC�0�#��}�z�kn�Wkh���[g�L
0(Q�(�:�^b�Q�����vÛ*���ꭚ���8D���W)�i��l����AT)�F���d9���%lQP��s]w�{�g��dJ���f�u��{��٬�QB�:�Bm��Ƣ��f¼���f�-C��.r<�T��~����-%�w3���h}~�۷Q=L�`�q�W��+g�u�_�Dy�� q4.��w��t�����Jg&#S���������R�Z��U�P9���Hk��Y��bM�j���$�J�cE�-ۢ���� �S��G,�60�면O���n�E^�)UV��F�O6�"�w{ɫ�2�i��������;�T��/��@�j2j��;P�1���Gb�#'K8�䨚E[)[��]fD����L��ě��G&�R����;L^Q�)��U:d�g�sPG��h��%���}&u�>'+�F۹o��ėY[�8�#T����
�:�gS��\w�t�{��o�� �aV�k*��u�W�j��)����m��e�՞����u*� K{���� U�Sѕ[��+ƛ����Y=}�j�v�ZN�A�t���=��0K-��w+�{i�{WC��Ίm콌��*{X]��^�1�wV${���G(��
���-��͊~ݝ�70w~qs��A��+�+Es\��r}�q� }��6�
O9*��9���Un�����5�[O�_0ά��Y#�m.=��5��o��q��~.rg*,�rFW�Oo����V�jZ�
�ŋ��������h�k1�9#��6�M2{���s&�E���]�Ye��lBӂ3�_`}���Z�=�[P�����swqg�� �X�޴��Άzb3wXu;/��;d;Xf��vy)�2\H/]Nygb$f��������k:0(j屐��$eӰ�c�I�e��Q���Uh,�	Kh%����f+w��7V�=��W�I�������5̵Y{��wVsz��Lx"��4c���˸Ѭ�Ƿ(�<\րL�LgP�{��mwQ��^4�"�G[�ϔK/*�7AW��W2�M]��� i��a���>�Yo6�������m�]\8ZÑ�5Ō�\�0Җ�J�(��]-N�]�����}�O��wB�e��'�+�rZ�UB�g�F��z���9�ث烼/�g��]��Z��'��|�X\��~����T��/�Yن���ƚ��/,���x>kTN4s5@�o�r65���yLj�z�"*�v�%�MôL)�^š���/*��R��y���[|�͌���炢0���v������qX+�AJ۫΋�-����@.��Sz�1kl[��S$�u5t�:+^��S��I\���7e�W�G{rC*�gj+c
��&��v0VUdq+s���F��)�;�ؚhj^�٬������4�ZG-���5Ә���4���d@��ߎ�A�
i����������ѷ'&�o��K3�xw��Y�-�2#���)�����YǫQ�w|2����׻���k,w�r�zϘIm�X�_�fv�uףΞO1�����[��B(��[��V�	�[�0VR�[��X�z��샻�#Ѵ��ήχ3���y�v�}|ו�Z�J�O�%p;���7����F�z���V�W]͊�\gE8jb�.r�8[��A۴���@Q�u��rWV�E7{7){��d�,�YD;��2�~E$,Ё�8������͙��#gÝ��1*Re�ر��`���ړ{軎�ıh.��Ok�Ry�)�"�HY>JݠEźP#T�UÛ�&�h�2ok^o�:��ru)x<&��ga
(�p�t�T�"]��ߟnY�ԡ�.���r*[m�a�޵ys���P+��2�v��]W���W!~�����YݳjO��φ��e��p��h��e/ӯ�~A]�Q`������x�V�lܳ�3��NiY���V�A�;�|r�=D5�I~p�w�u�Usw��ƪ��$h1�v�Q�f�h��G1�ڐِ�5޳]8���Z�BÃ�e0z ��{�x��אsJ�,�*����;� W���XS�x�HѼ��C��B`���m�Y�+��1I�vJ6G��݊F<<�9�fP���Ъ�1<���.���5d��t�� ��b���|{=����d]O"7\�9�	�Z;um��>"�#&'S%�}t����(w%k/�Wr��I3mi������-��� F^��:�$6�m5��-�N�����Q8 �]B�0��p�][Ԏt�е�3ñg�Ǧ����U]�L׮R��I��Lkj7w�׎Oc��5��>~��h��H��kۛ1���}��_�������p֔ �'heˉ�u9gh�D�\{;��p��6���t���؍d�&!c�9�k0��ݓ�9�@�(Y��S:M7`�i��ͼ��d�)�a�������*�C<�t��҆�ҿ\���~���� ��8��s��E��`��t��-Qun�
1���n��il@D�H�N�l�V��H~�T��G�h��׏6���ywe�٤��R(������Δ��ܽۃ
ٴ�Ed����,ү���a<���hk�ʲ� �Q�Z#س����L��̦g����e�@b���D	�ڿ&V��lVY��n{ͳ���1V�M�wC��<��lq��d�`k�Kb;��k��0���.�K(���1v�Ȫ�1A�S�J���h"+ؚ�AWV�v�v]�a�8e��0���M�=�W���ٖ;����|z^�r-OD�b-:]�X��ȹ�E�Y�(�y��.Ǧ��NkU���=�J�O�������q�����Iu�R��^x�����E�.��Z��Bd������4�)�,+�cup��\���r�JD�*����U��X��6�	����%�g�8�c��3d��c�C��iR4��S۷��w��D�'Q�N'^���l*6����P�N�~kt1��@%EdFCY�2�Bk[��� ��֨AN�r����K�}yGk'�^�.^#2Y,T,7q��nr�Ei)`�e>Os3��o;mr�c,5Mx��N�c5}
׳
Wd��K�%��5
n�0��v�k����ğS��9t��qF�y��NFj��l��4��Fw+rO���q���e1ZFV�Ɲ-:���}m^J[�d^��m]C>m�Z�D_�謬{���d�x��qyƸd`>٘
�ؾ�z���s=����Ǒm�/��`��©��cB���̦����+�Q�R��f��s9�ҺLD�iW�����s}X���	�`��J6�^ۂ�>:;���z]�=����>bf.�;Ov�P�Y��:2%��33��C)��4%:�jo�>�{ЗU�6t�X�TY+� 4H@����n������B�e��F�_7e�/����R��X��g��K��}_����	�5�Mʝs�hg�j�B)����_���)�0�p�����n����Hl����L����u�/���@�gfLЋ�W�"F�.,����u�������^�
(rY!Tvk�N���=oS�˚�ls&��p����Ɏ�(ڽJ.0�t,�Au(7@�[@��fU�'��mc����s�a����\�:Mi,��ܞ6:�	J[>��lE���t���h�:n�j�ɼe2�?%�3��.��t�6 MT5��lOu=���s�IzG.�	:�	�޻sPt)�?�Z��{���+߾`�T̍d5V�̭�ۙ;�ύT*z3n�v0��ȴ�t���d%]:��Y���`乏lVB��Q^�Y��|)�+K:�K3^�;���[r����2p�`����}+\�wAP�|:��}ږ�Ȭ_�{�37�}��r:��2Ф�~��V+h��~��Ƿc�SYE���mC��F�Z���CX��m��B&du6�in.h���qR��#���nSӢ:7��锊�w}�7}*@��4&6ڙ^�O�,δ�[CL�ɚ4���Xd���>�w�����rT��ƚ�oAYgX�S�u^n{�+&���V8	w�hh�5�c���1��3r�cNׇ?b�]�zƴm�(��&�`Q�LnSO{���c��!�����Pq�����T�HE�2B�U�LZ��YٓFq���^�PV@m�ՓP��Wc�&��r�;'�A��#õcmrw�XJQe��6)�d)X�e���˩��"*�<Q��̗��Ŋ"�i$%nЍ2Q"�s1�L�s���� �����^��3F�*�/���
�2J�]b�N6��`�_MlA��hrݣ�X���@-ښ1D�z�cؒ��@��}����S�L��{����I'*��מ�����(7�.Qk{�c��������|>��o�?.}�o�~��5t���܍g�u`����u\�.��Rj�?@�p�������s�hd�!ȲB�j�5�x3/�@�bO�3;i$�uL��Y��N;�*���98�+�TX@S6��ƭ=3 ���,m���|��v�9�k�CZ2X�y4�Z��kP��f��$�T{T�{J���%<���뛄d��S����x
���8�.����̇~k^ѽ�1�X��f, �VM]`�Cb���ޕm�����8
ӎӍ����˙��Ɋ�*���:>q��0m`����e�Yݪ[�ɓ�ųc��ckqI����}3�p�&4�y��Hn�זyA�����LN�����N��v޲�Z�	M���A�!	�e��q�J��}�Z��TcZat��#�tr�+.�;�
ɷ�u٥%6���3�S�ŏ��i�wNs�!#0^N����^<�r��)���T�)�hp���M�i�D�.����.ح�li�A��Li������
P�t�B]&;�s�JJ���T���d��ρu:���:\9�#zw,�[CZ�(�*ɬ}�:U���W��v�����j�8y��o�N��YB����K��}$�TҩK��a)/���� �f�W(@��QE��͂�i�#V�nU�i>X@*ﲻf6�2ٺl�2�^Ω]a��n���5�����<��%X����%_�
(�{��wWn���ٱGz2m^mZ��-�͑9�;Χ��z����C��W��I��M|� i�F���u�b�9���[�y#ef���a�Vy��m��ą$d�Ъ=\ty��>�d']/f���ا�;����w){G�G���7��}�yN��1���x�Twzvh��r-�:V�ʺ���t�ݕ6��R�7nő�$���19¦�1�}=3�x�-�j��u����◴��x���Y2G@Q��1��UtIЈu�S[�{8�ѵ��S3���%m�Ӳ�^m�[�T.��eK��<�y�����>��rGK���"wK����"�E��f.s�2�FU+�'z�ZW�z2�M&x���J����Tx+�;�������y�1S�'6�J�`�&��$-ԓm9ԓn����Q:2GST�"
>R�tI��5��`�,��ptc��buͧD#jYE�*͔d4uZ�lK/�q��X`���+�t��i��ҊOo=}bp�h�R�7�<9ɧ{XҘ�ͩ��W�f�֦!�@�@�4U�$q��d���ES����`݁CM'��]�+��6���%R�%�u�Aӈ+��z~{���j�:LŐ;�^I'ڨ)jТ���E�����\�똮�)�q�YhZ��b'�k��Gzwf�"�Z㡲��3��K�b}6�KEL��A:��(G�f�eNr�X�ΚpNle_C���k���s+ѽ<��60;f���$:f�)�7 >畼(֧l;�涛��*qZ��@�}UH}L��b)th9AȤ�JPP�b�[���9.��(("JA��T�r4�U7V��UDT%��� (q������:����������B��AH�G'AAH6J��
J.�bP��
bJ��F���4[bҘ�Ѧ�Ͱh�:v�
��:��4RU5u�� ��SGP:�jd9it��4�t���ZH���F���(b��������(ZH�hJ9�h���)(�(iZ�*#�ht�JJ
�����j*h(�����*(�i])X$���5����(�B*J(hJB����)ih4)�(�֓E&�:�8�I�&|�O5�Z����2�(���&q��%��w��w��0e,��w�a��z�MZ3�w���SPꜞ[��Gef�Ⱥ�]le�l ��Qb��2���{e_�{���J��K*�l�3��؂�^c��m�`g��	9ݑs#����D]i-�,�ȣkQ���dkfk�]�U�Ĵu_o�N�Ef�C\,�d�tއ[�}����"�2��il*���M'����AƊN�NX��抭�3��_����}-`^�.uǘ�U���w�$�U�u��1�**u��=�s�Xf��}����	��#�Հ�g�L�bh���0k>����f��صB���:���{x(�qk/x����G�g%ɹ^�h':|u��{�����r��I�5H�~&گ���i'6-���&p��~'�е����6��ӎ1�m��N!��nYȵ6�ۯӰC�;7kU]�wn�^V큪5i�u���)2�E����;�F��&�ȁ��)�����}�lG����BTY�:��;i�S�j��e�c�]���fᒦ����ݡL%�{�xz!^�׮�Wk�&6M�����v01��
T��c��ɬ���޹�,CI �mb��t�4w9��k{�$��W&
��P���a����<�!�%LD\�9�]��g�Go�\5��L���M���w��1[źJ@��ŉ���+"�m˄��bH֋�cf�{(/~x��(�
����7.�SG8h�By���9�hr��L���a�Q�vބ�~.�")����5}��p�Ż,�\ʧ�a�U��e	��h���Ɋ�wϏ� �q���[t5$�ԝ�7�UM���:��t�m�v�B��A׎�t�'m����!�in�:9��%.X�5]���rojz��v��u�L��)��Sd�+fȭ��7�.��a	����۝�mŇ�����%NН9nd�^D�G�1'�ޤ�H���v�7y(2��#6SV��<\lx7y�]�f�n�[�v��A|@��#V��D?t�n���A�,��t����Uy"Q��B�}����@������Q�/�k��a�7�Z���ͬ\7B�j�mk����tq�I!Of��Y����J��k���Q����U���.�	b�c5�ˮ�X�,>ҹ�'S7��;����n�].��,��ۑk4��f�G���M��-�6�`n���iۏ�ۨu�Xw�ơ	�;4CoOUc�h��Z})B�j�$�}K���%����R&D�j�k7s��"����/��6~t�kK�b��ܵo�=��1�9=���M�j����:i�R�TW�i�K�Kk8��s�ҵ���mVx�'�;:���<.��9�<G#A�O0O�!Ƃd>٘
����z�l�~�����4g���7S{Q�J��&��h�v���Ȼ�7T���F�9�3/~���
�j�Ke綽�b8�i�'�����Fb���-�ɜV�S�1�>��C�G]S��D�rCdr b�c���i�X�V�Ʉ���_��X�NL���"��
��!G�R�����1[��3Wbm�����Uo��K�M<�|2��^E@��=�)����%A�ib����g!ho�!�w�o�@l���a�2�����U��l��gX}�5�)nm5�4�n2J���A����9�i��+H9JnOm؝������RW �m�<�	j�7a�y��;�~���M�W�,hUxes������f,���k��}��i�D�jp��R�������N�p���+�P>��P�-Э�Z�/v�UdCc�dn������t�^�e�׈mM���
�b��G81%��+<H�����IŢsԫf���z��6a1�;��T��U�>Bo��F�'�uhaN���&�r�@��V]�
W����[,�c&����g���uJ�µ��4e[�ѥ#7yC�˓�~˞+�G�������ɿ��{:'�o��xvч)��`�ݵ _��D��%ܭ�'�Υ�F7�^��L�'qm.�\]�,�����zWY�~���"y��z�)�bȌi�i��jn��dy���#1�g�*Ɲ9Z�K`p��ӯ�:���v��l�3�M�� �\0���p��^Z����r9���D^��w>�{k��=�kZ��5֦��ݫLe�P�+�{UB�.�5�ǻo{��1/�o|%�⮬�m���'lu5{��Ɛe��3���ZژZ��p�Į�r&��b���}��fju`��2������U<���Q�X���j�svj��K1����������K��/׊>�5*�f��0fG�7+���Κg
[حG;�m^n�(��K\2L�5���G87�m�6�+��h_��kwe�����s\;3-*ݭq�}w�J��b;s��h�g�J���蛣u֭N��O�C���Y��ۑV��sz����A��X*tPh`��1�1�`��wu��v�v���ç��t^�j^��$���W
垆&D]�cP��B�p�*�R�K73����65�[�h擵fNв�h�T�3�Q�B���ӧ�d��ܘ�	��A���Y��$E^Z��Q�0��G���Q��;j�۸B;�8L��n!� [�-|�x|�l�B���xFj]^nH���o�Z�"��"�*��"��i�V�	����q��CLT.�v���	�WR��3�eXv�Lajq�{�iy�=E�h�ɹ��ˮ����+��J��<������{��G&�ow�=�}���1�H>n�@?���`���ƴP��_�����aߝ�)�6����y��2zI�/[T=fV@�p�9cEŅ��S=rqr=�/ڛ�j�{Q��e`P1�2ݺyZ�� +M.J��0���� Lb-X�닍Y�}��G��k�(�^�Gl�p�k�N�˪�[W��ih�jٗ�����>����Ўv�����s@�ּ��ٞ��nR�����L^i,�!�@=ڲ�<��6h3; �l^�^��������B]����5[/�G-������`h�%�;WIsyZr�F����5i�t�~8j\��ۈ�z��x�x�XIjOl���s�<�yL��f��:���Ip5ֆA�,���?1��+��|��j�^ٲx�~�@:���D��Uy��jp��S�J���cK� ���.��:���x�; �A�d@S;��Q��5�u�������A�X�hf\�*���{�;/��nD��deFf��ڂ�F�M�UC;�Kk���Z�W�]��Q��/z�s-S��ϰᩲ��-�R�z��US`�2�R�����yd��dD�t�mg���,�(�Ȳmi��{��JD�*�4Y��HB+��K�R��n�7��e�;�I�yest�R��Z�n�YU���L���nVΦ�Wb6���)�	�F�Z�p_<���X2��齏����?���-�����F�wX޵�ǲ����UӅPл���eAx�^̕j��P5� h��������g7}5M����Kd�+f�]���]g0�f�x�i��� ]�OwD���SgJ� ���٫ǟtS5H~Kj8�c��_j��dFhھ��}�KU!C�f�[|�-��gu	�YQ�:qb{Ţ3շV0*�p�}|]zGn��)w%~eܶ�pr�p��ս�]U܄VPeyv[n�l���.���Kk[X#Z
O���۫-#�6�ܼ�M5��7�w:'�nL)'}݈P2+;�rՅsV����O���kʜĦ+5�\�5�ЋHlJD��r�b�N�\rؽ>l#bV�u����C=aZ)'��ڽ7�y�pp�fDfl_F���Z���5�V�mE�9�\;��e�N��%x1�ѥ��S��.�Z�w��\Z���`�WU���5,J|��[���b<�&��Y�K�\�2Y��d�q���>1�tu� ʴ�Wƻ9:wz�S���9�[�(�Eе�p@_Uq���<Eɽx�����#�R�趆^�H� i��@�/<���͝AV��R5�o�ՌL�Ӽ��V+uV4��[g�r�������d�l�yե���K@��H�W���C�iP�ӳ��n5��B��|���{Ĕ��Cy
�����2�l-񭟰��F+��Mn��Wـ�ra��F�D�/�x�®,�V2�v���٢�j孙ћ��W1D�I��<�\��W$��x`Ю��SJ�}�KOu9��5-��anيP+2�۸���j��m���T��o��aN�w^�TN{��;��v���3&N�8�r	�U�8݊�k��dj�Kg��a���!D��I�ѳSSG��4���F�݁���@�\���Y��TS�ٱ��09������F�23��wk�ˍ�GVyv�N��s�YMY*�ħhWY�Yn�W����M���#s�<��W�F��ʎ*��l7NO#��4N�^Y�n��e�mN�{�1�{���l��PK��n�L����H�/�Q�j�;��M�zm��9���\f#R����꡼�!�%@���e�Ǐ�A�^��{�2O۫���s�k�,�bԾxhe�u�6��K�%���p\=�/��R�d�K!���1�*Ūm�V7�[lԧC�eV�邔�v�j��5	�|��v���[KV,Uw�j�5�fvL�s�jS�o'}�*-T%����X.ק�
�������kvPm��1�g��SK��P�y�m�m೸V�|�{��u����l1�m�����F#ٶݰ�TOqѹŻ�Z%�U��xvv�n﷬��8�!�� ��[�bTaK����%O����/xy똼OL"��P;;_ӧg��D�*R�Y��cz��?K���&o.�ڬ���`�v};�UH��D����9��Y8T�.!�nZ���ϒ�H�_����}IGH��|�Qe��G�h�hy�v[��-B�>�l<ݦ�vX�&�h��H�ɏ+�]8c�s�WcZ��ok���$�*�J�
��\��{��]!����t4�y�B�@Qe�:�c%IA^��ɻԶE&���+2��cG�=��C+4a���VC�����cX"s� ��ar���`d�I���۳��<������i��U]=�����n��u��d<������:�΋4ҋU27���������B�UҞ��djrn��+�^�I)�.k}��)=��"�y�}۴�* ��Ӈh�;2�A�+�����ۏ9vZ8�snp�ީ'�L�g;����{���Vz�k�;k�Mo	����ld��Zىښ�z�cBoN4��Q�gN&4�zןE잛y�d.s����4��5�ԥ�2�n =o>C�ijp�mR5� ��
�x9�u\d��m�O̒��w�p�֫��"�㯤작�t��(�'q��ò͟Bސ";�%;u�[��������]v̐Ǹ��̡Veׁ���Z��9�n�g�o��T2,6������a�uyk
��"ol�'��"�*gd#m�{M�i�y=wF�?gv����d֠8���jH�isWZr�w��s�-�����4���ᜂ2���Q�耕
�?�ӽ/������������5�\u\�P��f�6*~���[E��V^/��˻.G� ����rn+u�X���P�i�@����Z��@���w������������v�}��@]�(*(��}?��L��l ��������<ϓ�8VV �U�U��U�!�f��	�fU�@�e!�!�P� �  �*�2�>y�z��p�0�0�D\2 �　u� 9��EW��0�v å� � ª�" C �C  C* C �C
 C* @� Ȉ�(����(�(�����q�W Cu a�U�@ �  � � � � �UV@ �  � �@ � �P �UV�E� `XeXdXeX`XaXedY�a�``@��U�� !�a�a�``X`VV@�U�Q�U� ?���l���7���PiFdI������o�_�������������������o��D7�6���'��rWN���  ����/���A��" *���� � dܟ�/�O������W���}߁�^������z��!��|t��0���X����D�) � � &D �UY! e 	$ 	UY� %@A� % ��ʐ�) B�*���H�  R� &9�,?������H*�- )@Ѕ�Q��������A�����`~G��}@^���y�_!�"~��?`?������?AW�}�:~=��'�T U��@_�C�a�0��("�����J��� 3�����C��/\?�7��O���=� ��@[�������
�xzJ�����?��>������?x@��|��(�
�~���D U����o(t�e��&>�X='���O��=������I���" *�O53>��d�:�z���ޗ��=��QQW�=0`�>:EEu�/�>�����!�'��PVI��e'8fA���` �������g�>��J�T�))QT�A"�_Z��R�
�"D)��"�! )	!B�A@�IJ��*�DB�J�R�c,ڴ��͖R����j�Vm�A�:�T+�����(
�wsZ�%fՍ�TR� *��m��$(�J+c����Z
��J�%%*�mRSYDQ��U)kJ��J��VU
J���M�I%i�h��D�%�Si� Rh҃f��if!$�B�DHB��  .��v+UJ�vWhiJ�S![M5������e��H&i�4,��r�Km��&�u(Cm&��jR�RͶƔ�h�QJ�5�J�J�͚o� w@  :�� �(P = 7�=xt(P�B� Pީ� �B�
ڻhci��m����*���R���h�ն�ۜ�sZR�ж�����Q�D��L�J��+T3x  :򂕱Voq��P�*�G[���T�����*٪��f����V�i���LLP���U3[i[MVJ�2�ڙjUR�Lvb�M�F�UDMjP�^   '��iScT�/N�mZZ��LP6�f���5�m�4�Pmd��iMFV��Kb��R�I���j�5�3.�@ F�ڵR(�YH�L�EZ�*�  <�P���*	�LP �Lj�@ڰVRk�� �l� ܸU%!s��t4��]ܢZ�V�fJ�E-�44��  {��*�� 
.�� �V����UUrh4��E���&]� Jukm A�TL��\�T֙)UHV�  ��{t�cT
 ���+j0���B 
nX�@Tb*a� h� 5@f��h ��) i�T)�U+�  -y@R�2��  0�  ��  ���  6�n�:04 ϳ8 ��ۺl 0�� mJ�R�A&�B��b�    �=p���h���� jaC@�V  YX ��X�@{�  f�  e����I%4fժ�i � � ʬ�@�4  �{�@ ]�w��(�L A�L  ��
R��` �h@ �{@�)J@ �)�IIJ� *~�*��� 0�~%)P  "���F���zjd2I���*��� M}#؍�j���mVw��t�%�r�rM�+(�>��~g��.�s<Ͼ�'��	 BI�g/?̄�!$��BC��IO�BH�B@��$�$���;��������_�qk��93�QS#X��#�˫6)�Е�@��Vsv&�5�h�V�hl2X�Źdw4m�a��Pe��S���I:Y˺�z���m*T ���u�1�Q;4c�V��J��eh�>�!Ki���Q�5]�@��φ0�P�ۇ#�Z\���;7�:�������`qEL�S[T�,MU�yI�S��
�����'q1paB�4�쵿3�hh����AE��CX�`6�r�4�m�$�Ѷti��!�m�a�0�훺�%�����tHRQ�τ�Cok(fU�kV�1 �52L+�s?�pl2Ys*
qQ7�Z��q!R¢5�P�[�[|���4�`t/#�HwI�C͔��Hc�X�4l�"��T��J�W�U6�`ڰ��m�VlFl0���XQ����ư"�F2%���v�J{���ڲ�$+�Lef�G\�XJg/
vr[��*u	@bV���T����`�t��N�weCpeC.䠎,f��� "��ԏ-���*ܣ��q�/4�g4�s1�nV�K5l ��۲��h���v�)�C5f�Ĵ<�GA2��
eoʰ7���ݕ�(1*-�z�,*Gy�^��Dh��`�L�L��N[*4���Hvf��RZ�-�~�Oj���-ט�k���Y/"����S�fh�qS���L�n����c2�[�ج�-�,ϴX�%,
����UaZ�a.ރx�\���^�4.�5@�5s2���XU�$M,�u<���'�C�xf�j\"E��]fTz��T���26��FQ#�2*`�֌�˭x�f��r�4��n��bw�6���,�5��mn�%$!�5�%�1��ͧ6K2��O-����ٷ��=��w>4���^�6�#骟O�e��ЛCfl͵�[ZN��6
7�<�M�h�������T-Ԛ�V����9����I�X��B�j��nd$'�^��)Ի7��Z0�ڹ-
�$����w�ެ� �P0@0M!g.��Œ����x���r�ܵy�LەSE�T���AVE�kwo��7gPO$���ȱղ,GJ���C�������3\V�Xكn��qH�����%�����u%�j�a�R��6H޸n�EDtb&+��,11m�At�=��2�L�L�Xa��k��3d[e���	���ĢR��̧�)=@�um�:ʰ�Xt�	M��x��C	�ɥg�%#�n�%a@��(j�(,Ƭ&�	X��,�d�vl�f���㺙b�,�j�WN[�mAXH����n�!u��˘��їr+��&�m}������
L�*�;(RGk6�En�$� �j
�O�RNYGD�n�B�*8�i��O��Aȩk�Z��sN�h���f�ڢ�H#L;ո��8�`���ݠ7��ˊ�*5�ʍ���w`g���D'N�*۔�cm pmÊ��@�h��dN[-�����K���S̨��li�]��7�6@�mj�4^ǟ�B�D����%�{2��n�zK��(�jR;KL05j��A�^k(]$PF�׷4�%<M��@ͻ&l��U
WY��w���
���]����c_)�K!-{�97��h0�9���R`A�!6��x[��A�j0k)\�H�pm�T��+�f�#v��	�W�U�M�@f���� x���F�U�-�`�[C�mm%{)|yY��ǓSz�Cr
r�X�fܰ��or�������t�4Gu��Ӱ+4��\Wuop���T�I]*{tv����� K�3ϳ$M����8 �a��MB2�9Yh+�+�@.�al���ŰL��"��x���"e!h< ��-/���AK2n,��-�[�o��Ǯ���[I���s)��v㱩\�`�|qC�b1�r	�p���,B��Xu�F����c�3�rٳ��ܥv��B�[�����b�\K浊+u���J1-ԀY��R�t֨c�Aa/2ڬ��Y�L�� `{�7]"à��Xr/��Cd4-�r��\1��by��ƦU&��3*Tj=�3�T����n�A�E�D��%��"��;M�2kT9E[�gt��͈PV0Z�V��2���iyb�vVEOZnÛ�hh��2@���!����m�:d�bt�����*��%e�so�����j����hQ�LӃ>ͬ�Ä�/3)��"����\.̔)��=�oN�:y�mnK)��������X��ԃ-��Mةw�j[�Nf��`�ub��6����Y��6$3V���&����ᦖ���1�w������en��K��@�-bt�.(.mK�oIۭ"
oUk�$���Cj+�����%=
��Xr�t������1[KM�-�W��KT��I�f����d9{�CT$�!�V��2�Q�o�"52����P��	ŉ�Ԓ�������B�i#D�v�m=wqm��Ӕ� M��.�QxڭĘ�(,M����q�uVE���jX�'-jB��T�7R4� /V�T�^
s)e[R����)(td�ۦl��eJ{�*��(&��ѹi<��E ��fn��ѠV���;7W�����7�{�af#WK��f�")k�BF�R�]c)#39mD�BӖ�v��aR.*'l^ih:GT�oC�V��56��@
�$�5R5v ���d�pn�F��j�0Gz%��=�l�+([��1��m�8�ӊ3iA���ZNؒ(^��wL�-6U�-�;�xN�Kg�t���qcrK�FŊn�v��M ��&�;����>���6{��w��G��*�4#�d�d��)l����ҠI8"����ͧH2��O0��wj�%mH�Yȷ@���GA�^+�X��
�2�m��e����)�$�ty[r���ҭU��:5^�Bf:5��nG�Xf�[[ui�D���2��y��u�+Wo"��M�������w���T�[ M��D���3,�7b*��ff�S���k6)�$BJ��D����#g@Z��4(۳{cknf�;�V(�Ю@WHa�S��l���B�<�,��j�U��0�(��jL�2���W3�V�^-q��U���Bаq!t)�%Xژ�˫l]U�Dw��(\�.kF�4m-0f5(<k&�n�:�X��u��[��up��ug.�l�_n($w���ƫ:�&�z�3a%�-қٷ��Z�ٕ�0�6��[*�6�/��4���8�j��\8r����/ar#A-Mf;��r�ީ.�Gub�m������&��9,��d�4һ�
�Ez���k.���dCqK�p�X�cSf&�T�9��f���aw"�t,�V��K��"��4r�R���fm5�MH+JN�^���o�T©��,�;z���<x���;"�0��Qlr��Ƌ+n�ubPV�S��Sy�� �h����:�E�,-�̘�\�b�L�Bڀ�X�ݗQ����eJd�����0�f�)��x�u�ہ����� Uմi8B�U�ؿ�<�[�J��e�lD�6���[�]iˑ�`�h�W`�����ܥ�L\�ਬk�8Rumn�{*���̎��0�$��0�4䄛"��A��6�nb(P����e�E"�����җx��n�5`,Y9x��鳙�iM��h+q[��vD�h"N��b��++�
�2�
�[��n�R�;�B��էc������u��w�#��J�B��D���h�戵��wf�Vl�
]cp�)L�1e�6K���yd��)�����F��F$�Y�z������*�X?bMhF+B��-ٔ�*F��{eXmh��v�!K3J�YG6�����9}m��訫�،�j�|�Ie�2�l�J�[��Vk�d�:�Z�L7b�w�`4U
U���[D^53!ʄ���m���$�̊�5HV=�� {n삍�թ�H��*����-bc�Кzp\��F��*�J]i�z.Q�Qؽ�TgtP�l�u�3M�YnƽE��O)�t�ت3�j�鉺��c��W���&��V l����n�>$ șXFQ&�T�>�����l�ƶ~�@��j8m�*F��E�����!��Zۨ��Z����S2�9DB�4L(U�N�J���ä�VGA5Q-:�!����:����2��S2�T�$h���"�9�&CA\Eٶ� l��LɊ�`�M�a�9��"�ie�v�Tx��)=ceemGSon:9%�(�tI�-Z� {$*��ݡ�ZYX�c�*	��@U�ޑ(�T$!#�2�[Y2���[�;�b�
u�e�ZZ�Q��@1r:�ĤY4\�u�0��Gomb{w6�H
t1,[%7be��	�ş"��ݳXV� K�x@��R�V�,���B�t%M������	����jz��/\�.U�M�U�@��2�H�f"��*�Ã)V��#5�n1z)�;��h���B �w�{[�,�/r�b\{���"6`���x�7�d�YJ�j���UEtj��&�m@�h�h
��W����/�vB�X�8�K/�J쁢���IXd���ZvC���ڬ��f���4��N�S�C,��v�{���6I�(�	Ѭ�ji�����є
��)L-�X]�4 sqj\��i�zݬ�Wi���vUp��Vf����B+�^�4�;3Vl؆��8����fʺ;@Z��u�Հ�1��.�������O`�޶���'e(^QU ���	={q\_Y"�3vm������v�N�X���]Գ��0N�kRȅ��5�d�r�=u�Ѭ�0�e���Zub�-}�i�kEf'(�9�2�4m+̸����P��̢vGV쏮����(R�B��3�u1'�JoL���{f:t*�1�ʚ���U�m)�1+�j�!fh��i; ���������{zU!���q�VZ:���۷vn�;Bh�PB4SJ���W�wE��a�W5��сfbwN'qWX*ã�;`�bX��զ�J����2���k.m6f����cF�kd$�հ�Q��cp���Z��̊d�Rۡ�/��3"��� ��Ó(���pbJ��Q�%"p
���j�ܸ�&U!�^�i�be��m����ڲ��R�Ǔ��0'.Sg ��X� u���£��F^��oE
.�X�`�J�J�l�=�,��z�N��tcv�]⩋�n���a?��15��C@8&���kv�t�!e����~��C42���H奉<L*�bѩZ��&
�Zk+U�Xɧ�d�oX��r]ڛ�V�n��	�N����U�"�rO����IG�E7v¶ ;�"U���nGN��Ah��p�v����V�
��,���zT2(�~+Q��	��	��5M���0�Bs\H��JEbϲec�Dl6��&�w���8�E�h�Wz��5��Չ&5tM���ܭu5aG�P�@��2^�J;+.�Ձi�t�# �2ޚ�h�
�t�K��yN^�㒰'!�wF�Z4�7��+����ĕ_őH�v�� ��N�j�m'O�)D�͠S�6q5�IWr����E*r̘��u�ԇ۔輻I��e��`��ne5z�ܤ�Y��n�;kS۬�B�����N�T�yC��n�F����E1�X[�DѼ-`@-��4�k�J�n⭆š>ȃ�3v�WY�-��J�**��7n�S4^LnFN,���Ui�E�a��`.@��qX̷��6���"�V��K��8,�YP�A�w�U3�'����m��A�5�8�S�N�y����D�J��]�%��`�Cw�Wa�{yl�av�G����3Jb���ʑe��M8n��&n�;56^Cn�3V�-,�h�YSIKi��t) ����(����M���F��ʵE����l}D0�w,j�R��6�#s���*ֶ*�#��
���4�	��
TE�W�n"l[B���t�a�ƤY����YE���sT�a	�A���O+w�X�pMV��zԂ��2Ģ
����WLS���X���\H��\�w u�'���&�@�<���D�N%%m$oHqګ$�\f��_-6��*�Ś�hѱ���Wc�� VU�4�Z\�R0=̩�
v��t͸>n,�x���oT�݂�Ҷ�E��V��gsU�zX���yF��Y%��heY��j�b���j6U��в��ݫ��׌+�i�A!֎�N� �x,h(;XFӏ p�f!����ЩԺڅhk����yYA�b|،#)Rs*��i�X�b��������x�{�aS
F��n:نk���M�d��]�pS"TOۅ�F^��8Pu5@���9bV94E��it!��J��0�Ԯ���sZ�\tr5ȓ��踃���{A:r�ʴ^0`�9��oh�Щ,U�H���V���-v�˃(*7�����e�-Ct�۬�N���z�i����uN�O��-*��୛V�����@E�!z�5wOfغ�{�YZ]��⭤L�&�"��750P���w6�e�z�hd�5�蚇L��Z(-1^�C
!�:"����KX��:q1���X	�+l=9v�Tbz�#Bf�Ǳl�;e2	�0�1�V���Mf������	�%n�8��65�ϓ�a7X�[�J����6,ǫ5-؞���(J�
X^�¡��I�=�9d�fM� �.^S8fɣ.�]7YQwNSbJ�7)nnݟ�h��R��ꨳV�a���ԨQ���ܴĳ�fȱ�4���\ET{t�-�͘�8��0蓚ݽj��}����j(-.l�cR7o<}�mn�v&�3�Ţ�1��铖詐uD�̹����ꂹ��T����3d]M$��9�O��K{�W�Z�V���բ��U�X��_	݁�Z��l�%��u)f�:��teȽ��^��M`�ϧ�g\W�%ps{�J�u�g�q��^:�	J��v��G�\B�4��o~�@�<��5�؅M�3��9��B��릪�X���ӳ�@5R��Ң����ݴ��}ي��Ѷ�K��38b$�[ۣoUn���,��$$��|�J(X����GN;�S"� xE�>���s�:�*Գ/U
n�J�&��7"����;V���{w�xp�>tu��t+'W�v�a��؝3c���F�k��f]�X;p�D����fs�c�.K�c{^��"Be�i�)�DТ���z�u[��{��d �mJ������v/4vjM�f�M��Ԟ�c˼o/��OQ́�{�z���������Fb��s��J�r�jn��>� ��+�3jP��bQ[ ��T���]o7$�\w�S�A�ZgV/^�!g�מU��R�M���e��l��`Cs`n2 4912��֭�������L� w�7
����M?1|������PЯ��6�>O.]�n�]<�)ٕl��n��wh�Ŧ1��
�u��}EeDʎ�쮔�)í*�>ͼE@ f�;C�^��Y� �a۴���{�.�%o 3b�$�ݺxq
�w�:�k�,;C:��ʹ��\v��Ue�X~8Ы�h�GV�O0ҭE����f�Z�V�v�0���Z�X4�\�F��aʕx�p����r�^�@4d9��ve�5gmZ���j�W[�����Y��Bƻqc-�W�.�u�]����]��`A�&�S�v��cJYo�̩IWJBpPã���3�ĻU����01���m'wW[�ޖ���m�w]W
�fv����:ʀir�ǋ� d!�����3)��sXkl㦞��� T:`�K�w���9i�F�Q��d�n$K{����;�4������\p�t喡��Fӳ�J�s�GT%*;���Ԗ�γ��.��.�_X�Y6��o宷cy�nq\�����E&��T�I����D���oYޠ;0�H�-s���J��܈���xn��Q�
��:^�\=H�@���z���ީ�D �x�yݨٺ{�\�V_ù;��6�<+\�xDTw��]�	�-{�8_��l��1:��>`���#*�ߖ��R�yR蜡M�2�__	y �;Up�GV�� ��dǨ�ybn��m_]`'���=}2��Y�{dvyy������Y��d[�2��.��J�6*AS���uxy;�_-��ܒ��Yʖa<bj
\�Hw`�v�|�Ї�z{��3njjJ�2
^8���.(Ӿ��ؙ�|��y�E�l]fu�S/M3hݧ�m��/�Jf;1�Ha�g��βu��.LQ���a�a�����哃U��]�g���Ńc8p�2r�vu@�WV�{�\�l\r��"�a���uk4k{;s�Gn#I����x%r�6�>K��+�r�,���8m 黈W`�M*�L���I������Q��Z%vL��{s�S)ZI�N�t�19P��=�m!s
��Ӫ�޶�k��h�h�C�?�'#&�d��R�=��g�/���٪1}<�=*T�9S���19D�7W��P3����ǈ}\QA���d��u���ؖW-���f���օ3����O+,�b��Aݹ��Ա-��¥��2�i�匆�]�}�6F=�Ð���0�K4��I.�QHh0�B:շ�WI�Gn��N��� 8P��T�k��V�m뜾�'c��Fb�y�IJјW*\�GW�^v�EjJ�4��+�Dus�X5�T�Wh=�Cs��[j�p�t1��[�+;�����$���S�"�u��e�?a�sX�1��Ze�]�wW�{StL��X�z��c��ŀ㇫�C�Ե�H�o��r<�תQ�|(5�����m^;�V�B-���$Ш�郤s7�jS�C�ͲEhT�A�:��Kw9��`���s䮧%�����A\����[��ղ�H��'´c���
7wL���Z%�l�}�Yu�=��ގ-A��7�Ժ��EEy������2r�t�������k6[���C*]
�p8�ᕧE�b���c�x�x#����$%��[��)k����#S�[&"ym�!W&��Iz�)9���}��^U�4������g}AȮO!����w%q\��$����v�f�P� ��7�Oy���,� ���G�F�ɛ�q��N$䬰*�H���Qi��fAghus��.�e�ճ���mL3lb?޶�
�޲f�G��'��HÙ�D(]M���!7X�R��wu՚u���-4*���o�����W%H
��n̮�8H�K�B�Io u�1M�|7��|�"e�'w���r�$Al�%m�k��.�7��j�|��̱�LB@ʼ��b� 	�[���0˙\�"6"x��N�;�[b�ή��M��I�u���튽���׽Ԋ�]���U%��2���
NݩP泴��s�V(J��V�-�Ӕ6ݨ����4���s*�=��s5�2�bY�w��-J�P�T�ޚ�̮����u��[g��o*�ÂP%�΢rI.����}WM=Z��Q���i��́�w��}�&��T�_tҲh�X�Y�5�A��qN�fk��F���+Q�v]_Pj�X�[���>,��X���V��[�m�
C�$;��
i��9�a�V����uΕ`!ֳ*�܉�˶�F���*��My\��Lt��BPZ��(�O�9�Z�kH�
��Քn����A2�U�%�Z����V�W��1Gr�d��9O�1V>��$�J^ڬe9�g����e��J�|�{��/j ���e���8k�ʛ�W��_-�ƪ�6w�яB��]@[�^󫦂��6z@j͗}-2�W-[u%�	O7�>޷�h�.u�� N�0ؑ=xWL���X�$��ŵ�f>X�/�0W:=��޳�L5|��h��O�A�����q�R=R����Hr�mT�wc-��ݚ���K;�T�P���?E�6�"���������ĝ��H�`&�$ۺl�ܠa0������;�f��˰I��c9̅�3yk{��厅v'&�t��k+��v+�E�M�0ʵ�Bp�
�nHQ0���f���5���"��Ո
t�8��T�qU�o��T^��ʕ�ܔ�����;�S�����|a:yGB�ŷ�¹hÕ�nT�T��=�m�*�P��}$N��g�M�Cf���c�[��v%�A�
�2��������c~�-�f�C�o�j40ͽ�����6�g6z�5�F�U��q�[�(-U!r�UmKY0b�C�":�l��^��s;���>ؚ�k�{QV�e�y��.��%⦉���z�=r��D��ۥ.�N�&�C�E���t��8K�Y����̷g-
S+��Lսi�w1εΦ1%]v`�^����~�v[�W��*!��n�I��7NC-�(�O'3A�x�'m��R���۾X����n3��hK�PU0<8c8��Ђa��:�]K:��{�]?k2�.���P?�ufVp8j��y��B����{��T�l��mW�kK�V��p�W�Ц��BF�Q����'n���L`�l�9_;�4Y٘���)C(�Lv���wj d�[K�+F]�Bˢd�nV}��ڋ��x�9$�z�UeY;�f�r��Է��=�zt�ǫ���'v�{9F��Rt��*�*|Ԩ�fZX;�V���� qw6����U�%�Vd�4+�P ��J�&m����v\^�15VB�
�o��GS�20��4�Q�j;o��xs�9l�/p���|􀯅��S�y��d�g����Ӹ�S�,��;��m�3>E�LiI�4V�%R�WB0u�ݼ�d]l؀V�3fC�*�Y���!���<����5��dҵ��R�����)#3p
q�"���ES����4>�)��VXϦ��l-G�`�T+x&S�{m�ʵ�����bR�.�X�S<�GN��f�M:v\�Rp��#�����h�(K�!��j���	�)KZ�H�ilb:mq����Kq�s)l���t:�&$�������5�Hq&XD���⮧h������;���Z��I�u���ӓ���,P�X�n���{d�_�1.��eGY� �oj�_:4��74P2���nm*VQ[VV]:�����b������ى�HM��m��R���ʘ���9M�a��*ϼ������O/�G�m�V@�[�B*�[�Ar+b.����N�����VF��A'S{���ƶ�9���O2}�e�[k�Յ��:�z�0.sW��~k�Ǹ�E�#����ԋ��V�{���畿��������1�8圕kO=oFQyUb0��dySA&eI.���	��}W��6�/8����}�:����[H���Q[o��ux���j�2K#W�ݹn=s7B��A��v+Q��4�����Ӹk:�%�ѕ�>�ٗǄ�� �U{��=5��𜵎	X����v^�nx	^=uy7j�����4a8���y��F��%Ad�{@O�D'��'u���֐(bs��g4GLéjX`Y�=���R䌮�`�aN���wN��f��� ]��9Wa�ϔ�>2�4�[��oPƶRc����B�d��+-��-����\6�. á��h���c�J��ζı��T>��W�iy,-v��٦r��p���N�aChЊ�)6j�q�v�\�>�{�q�Y�_J�3e�p>���(a`��o���bJ�pt�Wj��HP���	��n9�%.M���`6-���#���^����z�
�hw�
���0:���589�$��+'�;6C��y���x��Ö;�q���.7u�>ζ�H/!�p@�ܲ�@w,�U�֕ɴ�s:�)(\���-q�c�+���_V�)��T��b�� �N�97;Ki���(�%�|.f���s*��+6�o�]���-:���]�b�7Ք��g�GC��#e��"�n+��1��P�+�fc�7;8m^+\��C��(�j�m�k��n���ZZ�wv�ak.��S��������
�y�ai�s��s��8��ژc���K�P���Ӻ&V���iq�<��C�v4�t��23�����}��PuhZ��_˭��V$g� �傐�S�v`���k�j
FgD�����L5 F�
=�\��9#
6�3�*fAL�L�غ^�Wى,G�$��z�s��%m��Jͻ��X��|��x���)�JnQ��!��s���yF�A�˹�����uJ�"��5u�خR�\z�Z�}x�;8ք	�H���n,�h����}6:��_I��,0�>c5������I�/8����՞o��u�U���^pNK�y��+C�:"z�n�K��㜫z#ZY�\�Cŗ:��S��j'�)�7��Wu�@�P;u��ݫŹ¦a�i�<�J�l�;	-�s)F�9W�^R�3�).��S�КQK���ьr/��� �ݙ]��!	����)��ө��2[�����;�ݽ��u��d!L$j*�.�S��Tn�q��ĩ'����ZcĄ��eHH��EݻV��ۋ�WM���m�6���w��{����(^�J�6�:�������3i�(e�Z �����H�4i���r�;��+�ڝa��O��ѯj�q�zާM���(�ι��k��lNtk��v;5*�T���#q>���<���=��T�@B33k��Vv����vӺg�g�X6d���:�MWwc���N].}b��ֹm^qF�)X�$���P���9�]d�1�V�*Y���e=
���G=k�vR�n�]�[-��j��H��42���E����t�.*���Ay�⁓�sn}�p������\�u�5�:V�8xd�u��$l����#�V3�_�2��]J��u�J�.|�6�B��ɶ�YԂ����K��!����[i�}oD���.6����M�z:izl�FT�pH
 `�*���9{�M#Xv*a�9]p�	�H��!9�e�i�����ݤ
�\�F�'wV�ҡ�:x�eq(Bz�=`�z�KЎ�MR�l�C3��&7�c���bM���6�R���<�Ԗ����`Z/�r�$��@����5��7u�I��d�b`�r��h] ��;:���lo6�whޛ��p���u�Poz��,Ć�^�{�l�/�5�/V� �53��5/:�n�b��tn4�𝹚Ы5�t�sa�8���b)���{~F{�(�c�2�IN@��D0����^G�
C���>��1|��,K@&���j*�\�o��e��UĦsFա�q�&���@M>\�9��������8L5�w��SW��/��A��`v�7��t��<f� 8�c�r��R���V�!_ �&h�.��WA)�=Ѵ���r��n+��nJ�yw���;��ñ?(�oڌf�z�oG�&vc!t#�R�/`��'ݗ�<���6�i�eL�D�K5�<�{�;Y���F�݈��!q��ck�w�`��+KY�kJ�*-�͏H3n���/O7,42�&6~/v]�V�MF����*��u��eЙ�����C}<k�Wpn��
��}��M�ӥ�{�a��2������V���A�Hk����c��1����	��ƔH�m��R�h=������w=}�6�z�>g��T˭�Nݬ/��rSo��wuH������s�X.ڮ,A���]>�
�o�}��Ͻ����$!$���BH�w�O�8K7D���\��9�z�WW#ټU��իk��q3�[�M=[��e�1�:��66Ӹڑ���5�-��|:��,��ⲇp�
�+c��t2�o�3vh�j;��6>52�C\lku���G��j��םy�4��-�Ʈ�G�<�Բ��������>��w���I
�ֵ+Yq�t��̀R�T9S	� {�6�����J�ݩX�"&��}�ԟ
��"er���x�r͛����� �l�B�����f��Np�1<Wr���8\5�s���ayxc�M,���'#A�b��7�����oqz]:����k��.���:�e �(��s���"����E���*�)	���n��v�	�����q�k'e��n�.�v��GPG#1we�@���3Ȼ5f���(��[���R:�H��`��r0��{GGD�Z$9�L��v�V9V���z͚�w��혪���ZœZq�<�Y�޼+�6�.K��oB-��{kJ��n[u�)jS;'gvȳ]�e�t��Ƭ�� wa�uM�sCh>�����!LN7I�ӌ̑�2�-{t�ر$��*F�q,�
n�|�c���Tb͎Z|����CA���a�F+H�n�.�'T�+��d�'N[�=nRy{)��i��m�#��x�z7u�[���;6�<~��,�/u>sk6T֘3&&�ʻ��f���һd�iVG�0�C�,.k�n��x�EF�Tubm��P���;x��v���
�ʖ�0s��ر���ͫ�V��+;[�&�B��WR�P��c�.�J���#��ڣ��j�wʓ+5�)��h��C�5��e�D�:.�,�ܜ��**vr��J�a2��i�J�ۑ� T����+���� ���kr�V�V+.�ω�qɕ.11`����ۜ���)�����v�Щ0b�d����.��,���hͬ����G���@�k�U��j_+��ڨ�e�{���_I���c�ol+��Eed��TP=|�b|��EÊ���t`�. �Jۆ#}�s7�Pl��¹m��-�.�:/���dn�jb�-�p�uD��>����i�����l#�pE�^�4/v⺶%�۠.�ao�n�I��#���L`O�7yئ�׫3�m��N
�̛q�w$~���(��n�mP:ٖ8�p�8�]����	��h���|��K6���R��{yh��۹gSAҶ����ĺ�v�iʒ�u��4{,�x�p:�:3&�]�ކ������7��-p�	�F7�O���EE�'�&���Pӭ�V�B�vl�kh�_bm��1u��_n�׷�86�+����'W��m�Q�!�|TU�!����&)Z6���z�=O.鬴�S����m����qR�5q3�S/3G2��)��r��/5kM�s�`����%�qSH���������-
<�$�;C%�
�Qu|���j[���Q�|�\
y�R�t�胚V�s�C���I͸�+���+&U�m������� ���L3.�^��H���^�P���J�P��2��.MmG��7�tf%	��0u���K��\��k���	�Or�X��[#�t��g��Cy��Z9��u���o��묭T���m=��T�kH���V�K�)�r��E�ހ%@%��O�sVv>(�F%`J��'!�b�Ի㑤�8���:��ѓ�ށd��f��I#�����~u��uթJe�ϛf��R뻊�9��tz�d�}s����F��v����S%8��j���Z�n�ۭ5���4�Z;{��P���+nH�:3�0a������8��*cl%�f֙A��wص��Ղ��w�F�엚�1�cC+X������Dj`�z�wϷ�M��*sS��쮏�u,i���]bn�u���|�KkqM��+9O�wWm�B:���fjS���:���ݼ�Hy��@���s��ӱ�}���s�1҃v�Y��i�CH<�:����!lg�j\�����g-�7fGԫ�8���ȗ�r���ph���]�v�S��/���6���+�}o2�ﲮ��%piB�k3 :z����L�Yb�w����*%�:iW}��t�|ͮ�g��N���zEJ-��hm������w;F:����g/qu3j���Aor�L߄D�C�暺�̳�A�h!�f�{}z���1-�̴i�ė|�2�b�uM����{��DJ�R<�Z�L�0����;+�r����lp���>W /eE�2�Q�c2/S�4��\��`��\�ʄ���,��Z9�⊘|��	&>��ؾ��k�q�V'��*���bBH�@^��PSvȦ�;�`)�ڛ]K�lR��=T�k 2D��o����['t�Au�����9�%����#@��D��H�\n��&ɜ�r�FÐue
��@\˽�9������9������_e�ojte�}z4����t����i
��
tՆ�|��rWxu`[)p�6��p^�����Z w�&� b`,�2�JH��Ǻ��.�x���k8�º�2�=��_s��;7S�Vޗ�����ȯZ�tn\�tZ�V��GN�
���`<j'�\�1j�O��'����xu��^��xP�-�WD޶mս�39R���cM�.�� ��C��@7����e��0�B�A�k�;F�� �_cN�e��X��*&�t�d�T��Y�����������r�j'y��q��`��]��d�g@튉�]������K�w$mp�ɂ��=��z�Qk�,��T�.u��wJdyF�S���X;K��Zz�[�0��U��z��*۩��5��(I)�fβ���n*.��;2�k=G%�Ӳ��)9�F�̂��WS���oX̴ܬck2��+(��<�6���;�U��^��(�2�['�k��B[v_<)#-p�NcU��NY+6�5b�)�6`|/����΋V�5.��6���E��I�U��U��U(�u�:�Bǹ��mۦ��n��v��:��B�j�'8U�nB� a}C���]�d�)˩5ɖ.���ҥ���wÈ:��;�0Q���]��nwثЈ�=�!�u��).z4PzGw'�ӛܲ5X}݇;��ض��ú�mt����[�Q41�-�`��� $LTn�zԾt�e
]��ڹ��Ӡ��Ufk�)�>f�-�;I�ͮ���ϓ�U�6\3�:���E��ݙ5��S��[�a�F:�@f�e�[Ӟ���h��ݧ��@J����s���սd}��!�f�5��V�e]q]8RC�k+8��rv���Ut�0#oB@^�ޫ�;�Mu��)���i���݃��@�;���݁"VjU�qv�N��'.MP�ni�l�dZfnŏ� �n��4eX��t������$�w��ݎ%�j��{*/�� �xpWEƄ��)�LGkN��E,&�{p��t��99\F-���
XÊd[۽;V疆7�L-���{���ɴ��oso{q5����XY�Gճ_[zR�vJfYh:Po`�oq��J΃:��6��K`�wZw���((+z�r����oX=�PP{Ѽv^�(L� ]-ξ�ǖ֨|3��ڏ�D饑�e�F��[��Agmp�t�5�[��ŀ�Wdዷ4�Eԭ�8���	s(w,�jR��A=��<<����[DK�hRk��Pvjw[�8[��ۙ���"��arl:��ܺO7�)��<���% \__=���"��ʉ�R]�xz�F�;P�;;Û��;�=���r���[��Π�>TU�(���W��Go"{�5��+3��Bl[Yt0U2�o���#�*7 �t�9XJT���2��wsI�Z���Mj��'.��3���cun"Ɏ�m�\�����=��j�uγ+���gBׅ0slN��޺q�dZ�ij4�]��TE�;h�O8��NQ�9FF�ȭz���.gI�AO���)X�a�F�5�`��Kylw��e�u�-�q��B������5|2���6���RS�/�� ����TL�̨G`��p��8��*ns�u"�@g*}ɂ��u��v��<�ZV8P�':.�1� #���h���PE�J�mvHsM��Nֿ��[OY/��������vK��]��d�����CJ��ӟ8�?vf�EW�
{$���j���f�xM"I�9���nC��p�۫����7)�7����`Tr�:U*��N���[%�z4��m�uZ<%���2��jڲ�°�J<6�"�4�t�{�gr�e_vW�:t�m\��Rf��K%Gо����c�����V�v5�:[�������pCu��6�s*�d�]B�+|c�o�(^�=��ۂ�M�ض��\��ov�V����N�'y�/�?��r�R-�}b���pŜ(��n%��q�N뒡���|����!؝հ$��6�9��hjS�vVP�`��jS;�r��
�	�"�}�ќj���4*
�}��$�7F�3.�h�:��z!�[Td�Ӧ�W�R�}�.a���C�����]�uf���d�}���"n��7�Dk�swi��ltp"76�SOS��[��wNP[�it�r��`����k��Y0h
\��l�2@b���X%$Ci-���{�E�fS��YxtR�G!js��=��N��ۗ�Ƌ�f��9�O�E� �	���ۭ�l��8`����b�Dm��T���)[.�ơnT����&��@)[�*M�1�Xt/S݀�G�т��Xlv\��x����W;1hee�����WĜR�*�_9d�+��n�4���:H�7�	�u����P�5���vԩZ�Z��V�[�y�E�ʬ�q�\.�S����l��P��TYb'����w�x�(�ӷN��
�:���N�8sW�r��xvvHљ
�mk����r恈��F,�����#�4F��Fy�<������N+�&����o,s�'�O{�^r*���`����$�{�N�Wp��W������}Ymxp�j�Nx�ֈ�mNۆ�{n�g���z���뱪��N��b���ĺ���Rb�tx���wOS���Mc��!^��Jb�{�����g���2#�+&�g|f�FQV�|�wS�Vp�sw��Y�9Z��tB����k���Q#��n�ٻ�N�R=�1���
�� �/�r��ck`ъ�U�t��伦prr�QAT��}w{�52��]t�@��yz(���N^�����8�T�#��沩�W0z��ǳV��w/���duc�(��F�6z�41˫��CK�äȱVTdJx{1RXs�I��s
��x���\{iɷ�\�Q1���캎�[��K7նq`�"�=��'�ܺ9ݼ�(���	�f�:�&l�A�ިgb�^  �^��)��m���>���ɫL���4
������أ�;���^��k��w�85�r��h�I7ה񗺭<���yF� ]`�v���]�4�����[��މY|�94��*:�#�i:���z�ZNZ��.-|��L�E�P>����·r�]��C@hw;F�ud��tY��������0X�`i�Ї(Ȯ�=���q@6�\��O�Z�]x2m;!K����}�9�	V]ѭ.�8%�b۰�e��Z|j�P����LY���ZL>�99Z��� +���/���o&��'i,ƧT!��9�WdN�u-�����9��g�&k���b��5;��c�٠��Eݐ���#I��r�7hr�WY�����aǘ�|-���6��º�2��$Y����J�yi����9�����짂�;KVwn{��9I�q�f`yKU��mw:�ݻ��h׉{T'.k�w�K��o+y�(kb�Bt#��k����O�s��<�=}֗m�W��S5�w����4���X�XC,J��R
�cp:���i�y-�t��vfh��vʸ��n��rd�.�\롻��,K��>qJt�\� �:;�'�:��{��U���!�D���<S ^ۗ���lm��Z13y�l� S�1�JW1���=��nvui\�-�����m�����:����+�������c��Nq9N�]��Mp� v�S�c����kK���١����u-^�@�ѻ�S��gr�o�ل�.�R��õ����G��u8v��Mp��j{}\_k�.���yn1�J�?bPM!�|�/ <�����ˍd	u[%]c1iUx4��9�)SL*[{��U��̥��d�)9�P�����7D��Z)�� fA�å{���t����u:��l��&]�sN���k��ʹE7���ĺ���ץV�V9LN����W''h�m^p�^���&��٨�)L�Bls3��ֱ�l��Yug�S7�!4��2+9��+\�;�%�%���C�,�ګ��N��v_��2�m�8Z�q��/+��_K��R���#�9[�Ai�ӄ�}�s*�ѩ�i��wB��c��a����"�')�INt�n_c�@����gjd+�fn��,�ڕ��q�g�mD�y*س�F�-�^C�ի����l#uc(Wa��א�K���+��CI���eDڳ�X�}�z�+g��*�
�k��ԁ)�v���^�tl`�l�Y�e���>�җf�/ �!��$u���ؐ��M�ȫ�w�:v2�1k �h� I��k���*dc �-RsK��{t�jf�)T�&�wW]c�s�\������f�k�+7�e>۳J�C�u�Y�D3�aTU׻��f��t��m�0;v���Y�z���um�k.�R��K����}��_W�}*��>��z[��NDj=h��([���XnW)]�H���1aJ���Em���=z�GG�eM��%iW^]��j�[Dq�������q�s���w�gi"_٠^p�|)�ǎc�m$�9 1m�j�l;�c����l�˚�^wv��W)�v-K���,�Z���9�����-��X���x���ܥ�Tu�j�4+7�+s+�r\��.����@�T�bٝ,�����A���	�9"8B8�t�|U�ߞ�$�d�S--�D7����W���(au�{��v�.rѽ�t��ëzo�o,B�g3|c;�Gq����S6E3/jݐ/l�*���p���ëh�]�[�;/�v5�M{����G6��r�5ݳ���ЪȴlWo�Ө���HЖژ��%�����ڮ2��ˏV,����wʬ�ѓ��@+z�-*̮�o�4b_�����6�պ�l�}��%�i5˄��/xr�������[�~��U�Ho j⻳}5��+�8��������/��"�anKJ��2��'�k*ږ��C�^i ���Fr�����ⱳ�;��7�q�e���,\x����v2�P�n���j����b˝�x��{������W
]�}�n�g�geҭ	�X��u<|_]��q�>�Dq�9j�y��Բ4���iK͛�+.�v񸢘��!���+�.#����}U�UUv�(
�Q�`�1*EX��`)PPD���
����[@�YPX�QV"E��"����b�)�U� �,+Q`TPU�(�q�H"
�PQE ��X(T���a�%dEE�k"�J��mE �XE�
2B�%af*�R,ģaR*�`�bJ�2R�Jʑf�
ł�֩����1TF�C�)��d,�J�b��R�2��H�B��"�,R,MY*L�1����`��BX�c*V�`,��U�,h�(�2�Db�"���_+�.��|}���N�Ơ���^&�T8��<��c�ٶ���X���@,�Oq
Y|���;ޅ�ո�N�uW��-UQ�\{����LT����d��_4��,��
�V}��Ӯ��I�B知��<^Ke��|�ՙ�,���P���C�n|�T�F�爿��3;�`q���w�7E�P&�6k�[.v�s-Z����'�|OX>cC5�s���:��c3yci1��_/9�n:���[��"��f��b�!���2p]DX�R�n�O;�v���dᢻp�c�fT�U�Ù����s�Y�3]O�y�[�T�����R���j�[��܋�Z�\�2_a�l��f�k�j��DJ��(_��ђ�5�a�Yw)�����'{%���J��ã�{���PدO,g(. _O��p};<�1�sW��2�E��z����'�{�����q.q!��}'Ρ�b�;-�NIB:�x�ך�c82�j<3Sq]�S��!����NDq�GNș�(�o�S=+�Z\k�W�ʻƬ���5�NFɍyF���J���щ�a!��:X骮Vs��e���
���*k7ȿ�xVZ�_z?f\�fP�`���a�8]�+N�T�2��G�%Ɂ����ث���&A,M�S%�)������&WX�y��#��z�ŶEo�)G�n�T���W;>ʝ��و@�.����3mt�[�Z@9�{�����\�9�L,\�p�4��{�)�����Vhl�1$�2�u�}W]3՝�h<�q�`�6��:�����C� ΁`)Woܮf*Ӿ���-���F�8�ǰ�Ms��r�X0:�h�g�jg�� �K.Ո��v�L��g�YoA�7֞$;紤M㩗;���;�<�~y8����	[5n�RB��\�]oF���ؕ9��K"�)���J3���'z�=]��Ź#�	a����"�r<�xh�C��:>4�e��{øh�5�r��u[Rcp��%	����j:Z��A���-� t=�E��Fʥ
�$v�?��=\f �����E�W��gP� �V�Tbu�#"�˃��_�x��t�h��n�_zT]�*�n�Or�_��ZP��)4I�4�,����(����e�Ϟ��d������i�p)�aZJ2�"�+�^VٯKU�/���SYg�����9)����{ΘB���_q�Q�i�kԐ����s�0F��x1�|�ͨٽ	�S���B�/;ʸiI�l?^dアx�`S�ä�a6'L�:8�86f����Gml���-P5�4��D�x6YX���ux#��V����?T<+zbVE�c)����ԏ`���&�z�q6��bV+圪+��L�kXcD]�-�R�j��8��ѣY.��z�ZC���N��3�v=u�Ė��o�]���poy$�>�YW�(`u����؍����+\.U����^�b1��N{�Om�x�v(��5����)�m}��^?k����gb�{��*�,���PK�J6q�)�Ϛ\��8�J��ݹ	��	#�Zz��n3�P�+t�,������^r^���)�e]�k�j ���ϴl}��25�|Q7��>́j�Vk3��'*#qV˞�Q�����L�H0:4B�b̄��Um$9&M�7O��;/��	j�/�C^�=ٺ�e/L�u��r>����XZ�G"�Fs9~�Pf�h�=�Y�5�"j��}�%&�y������8���;P>?e������/#齮�.6�l8��Gw^��P\��S�.��X�O��y*#����Txs��_Q��5(Wцg�	g=S#�f��"�r�6U�r3ưV�>J��d��:LF�]�EAw�@�z|�z';ޢ�+�Re�)S��O��kFČ�c��6���V� 	Hm��{�0]t57��׳X���Y��X�1V�Z��D֜T�|eM�d;�{��˽I]�&�d
`5B�[���7:��x��r^9�����R�Fm9F9x/�� ��M�9�⛥�P�W�=��h�t����i��TN��x����N�K�R�N{�M��SS8��a�n��L��a�C컼��x�ep��k��^���Y�e(��>�y��9b.��,��c*���8�L���̳Ks�_l���4[�Ʀn_��w�`AJ���F�7��=�fS�ͥ��U9#��)��<ZM?cޏ6:u��4��U/k���5�B_�*�r���1����+x�V�->7���Qz�K2Tǫ�wau^�p��.�N���gW��[cF|C6]ꕾe
ދ�i_$;P.r�*���k͑8����S�x��:���:���Z2w���AL3�V�OD&��z����TD�؞�*�c@��ܓ�ۘ����|"�����y|���.Ϫ�ꪭ.��j����P��WP��A��Uj~���pSS�;<7Pgs�v���;��R��6ݵ@�K찺Oh��ₒ�>�����-PW�!1��ϳ����V�	��M���V.A<܆��=%.��/�2+%rk+ �)L�	�
�x��=�d��ՊS���N�߯��@em�:�56���O���O�����Ey��ie�c��U�1o��x�g�`�E�f�L�Vzzl{#���H�'��ԋѝO�c�_գE�Iüp+g^Xs(Dɘ��8���z�v(1�ү;(�Q�Y�r�|rtU���TZ:SIfF��6%�IĴ���-�3
g����6)�!�>��&�2����eN�9<�髂�$!�U�l���ҘYe�
w� r��U<[�n%ٻ�/��g�R]� �Z4�9�������x�9	���y�̈���  �/^(��$��-kp�QP��[*,t�"4�J[�bL�j�-� �{2��dZ��L�X�����R�::cf ��H��x*T�^3>�^�p���x'�4�7�������kӊ�
7v�`d{�4(3^l��c�[#\��pv`�Q�"f�읜��Y,�|M������!*�lc���� Rt�]�
s7A�忹�~({���v��l��w���g�S�k��7ۿdCU��lp�O�W�{����s�{M<<�)���H�O8��ÍBC�m9���z����s5�q���u�����zj�[ۭ���΁X��+����{:V厸8s
�a�� +�-�UN�"W{
|�d�=��sޓ�<�6��m:!:�^"�7{�WZE��	�>\���bO�+< ����ٷ�C�Xt��'�-�/��h'<�� !���}��CV���{VȬ�g��lIկ��H�C�t�Y�@t�Gцmp#�z���GPYm�5u:���,��&P)�v�Օ�afH��u���/��\�C>��uZ������yO�M�v�8*��o�D��q���-w-�J�w����A��/׫3����]9(lM+��/�c1�&��7g���Yh8j����7G5JxOn3�o/���o�U3ҺZ\k�`^����<�����܅a�5�6o~��\2l"61��9�Tt��,ڙ�6���{k3��Ť�h:t�U���u�h?�t���v%���d42KGp�N�c���6aLr��!h���Q�-Emsy*���[A�@_�
��L�E�}5$���t��tZx���W϶���0t8�4��+Db�~Oυ|���؋�ѠA���"N+�"z>�쑿'֤M���%`�����K.�Y3(+V�=]��WX#ƱѪ�)�a����!ܦ�sP�9�N�S����c��TV��2K�31p�	����JT���`���]�vBc�&q����M+���C��`q���m�8귏��]���X�:��#H5�eҏ�9�ԕN)����y>:��o����f����uѮB���3:�4�"�h��V�ѸC�횑SⷛskrWB"�+������y��5%�fٯ�r%��:k����F=މ^ʸ���B���땆��4Z�wVk�]J�Uf����=\�m5��3Lt�JG�x��������kS;��<>��)s�
��.�2�>N�degG��C����b5�\\d��a§�ڞ�ޒ�窹Ռu�E�8X!Y�/ ���E�j������J�,���xѵ�蹾����c�`�3�~�Uٮ���^y`)҃�
�k��$zѕG����c<߂~�}��������}��j�:Wꗦ�P�k�;�c�й�ć�v=O= �g�W�j{�ڤ��َ����q��٦GY�5�:ѪZ�CT��p��R�R�K��85�Q�jSH�>�:yz#��=�)C�5���ve.V#G��huH��K~8��z!�����Vӧn}�㑐�������OV}�C=b�Ѻ�a�}�oU�|�9�����UX��Wگ����t�J������dwC}���#o��"7j����;�ch�,�v��Ӯ�]��x�����b���v-�j\��R��}4�F|�9縇
�#�'gF�nHU[�NDk�R��b9�|�RV@ϣAav���O��P��F6��ET1٪��R��X�e!���;�����ʌ�r��*��I��Ѻ�9\#j�^�/)t[�y��'����ʱO�nŋ}��=K�����d�����ͅH�H�As��!�vSaa{�S6�����;c�ծ9a%�ڻ��	k6>����}=�������6Ǵܙ:t��_㠸�O����I�cص+"r�r.,�U���u�w��+���%w��:v(��WQS_L��6�է�yC�/"gôHko"��,U0g!:F��NK��uю�*�3�ĩDz���۬!ݜ�K�pz���@t�FI�;g�ړ�ʷQ�:�WU��A��� \F+` .�z�ݨ�ξܻ �V6��/�q�@��F�Ps��mOdc씝[�j�B��r�����bg�lk���}��$��-WdWg�刺�\+�}��î�_�qB�֗�(r�h%�A���6�Фg��\��C kx#��<2�P�s�5��=���t1��?1I�[�v�d�Cu�҈��r\wLj#e6�{�C��?��5/�>F�#����a	i�Z`��q'���gv��
��Z�Ybq��'�8o�y[� �l���E�o��x�q{�!��N�c׾���fU��n.ev����.®��O>5�S�� �S���y�r�q�4��{X���]�Uڋ�C�oZ�=d�3�{��6�'Ұ*����R��`��/��:��}�����^@�Ա�hc�2�lqk[H�Х��0���3p"�=}��k��ɏy�pv}�*�^�K�����^��g>��,��Pf�9�Ց��E9����#~��R{�X��gP�����E�ݫ�Cni!�B2c���ɰ��P{��.�F�F����]�����d�Ҟ=���-RN�qGs����2w�J���u`l�UBaS���u�
;�YPF:��%��SH8\����͹S�Dڜ�Vȭ����<���
��
C�z�����l�{����V0r]�OPv���=�#])��;x�6ܠ�fk��n��s�>�u!�cIu���U���2Ќ��bT���)�B5�VX�s&Әq��RDBȝ�s}yqڻmv�7�?�ŀHz6�s��ܬ�k>�s����U��@��������C8KS��1;�\EEAWh����g�"#p�R�v�R��W1l2&]��y��-9&�pG�!I`��!�B�֊�Oi�@�9S�R�F��Gs�f�Lt��mfҸ҆��D5���o�|�v}\��[9U�5׽b��5����9l�s�u���;]�y�K��7s�_:0Q��큥���Ҩ�uhݩ���/+R��)��t)�� �<g�v��w
5;0���uɤ�qm����Gf�̮�;��z@T��8�� sn��;�l���]�E|�)�BK��w���ΣV��t�R��tr�� q�θ$��')��Ι���f� Ҕ�NNIҿ)�t�zr{��a����N6I
����Y^��8k��R!�V�Ęբ�ޢh��̕�o�?�)B��)y����@B.5�2��{~z0U� _A\3	�ϼ�G^[�s�n�չ�\*��TV�WˁN�� ����s�Y�3�N���j�9\"�58+Ɏʒ�R�ū�G�S��bڗ���AaYuk��X�4�ȍ��
U�x1��V���	Ξ�w��w�{��.��0��}�|�Ww��!���=���l���be�o:�\|��g�k<�$���z)���2�����2�.qJgG�����u��2
,m���M���ӌ��,�p�\R�9����8'����m���A�� ���]����y�9��n��w��_��ѐ�6����J�Q���P9�3D0�t�WYQ�D�n��ImT���wP��2�.1]�ye�����s�w=g�.��J�b�V*u[�.��!z���T��x�S2`@W\ ������獵 ���fh��"g'菲�guY��,*����<"��K�G�I�=��[D��a���a�qТ�rO�j[���� J\�֗$���Pt]>��=��0஦�[��A�0tpSҺ��Il�ܗ�b�}��=��ƕ��������W �O�W��׽���ͩwS�{�����*�e�u\i����miYcvZ!���֛tq<�@qZڴ�黑˜�+a��SN}˞Q�������dk��PS[&�k8�^ё�
�G�6N�z�a�dP櫤_8�wz��W`B���Mk���5�г��P�;��]v�<
l��%2���R�=eT����o2� ���#57mK�f`�,N-��ZK%�#xTBMЊ��Y��秶�i��Ckr!�E�W�D;�S=k&ƧF�� ��6�b�d�G�JٟG�3��X�3���.[YA��z��$7���$��|'����Ǧ���"ӣ �'y;�q�ͺ���Qq���7v�ֹ��)Jgk(b��S��ZP:4E�duu1m��)!]d���R�^]�x��1jZ�"�Huk'c���B�`q	cqv�3]��p��cOD�p�*���	��_T��;�U�d���TGhU�]���I�¬�;,�-N��L`_P}�p�JLO�3�� ��oH�N�0�G�]x]^�MG"��.s8�꼃��i������6�j����7��:���x'�����0z������* j�b+����kN};x�Y4�:t�ѝ���h� ڶbܿe�k#�����y�:���I�Ш���=Yt�&�KIۃ1��ӮusC�V�<h�!�6�D�N�K����"�4�ܙ��,��Kk6�.+x�D��-n^�&n*��]��Y�wm\�)�x�/��˷ �Y��]�.��#R�c3���W �Rq�75A�si�d��,�R,W6;�]+��^�L:��N�n.B�ޚ�4�����r�e]���Cr�6S�nv��������1��W=�BS�C�jΧ���!���Į1i�
�vK�@�7�V���lT�Q��U�
֪yg���̮B�:�c�ݸ���9d��B�$jà��:��(��ÚW1�_(-�o]K[[��}��8%J�:�� ܞtU���p5ϕ@�U��}�Iܱ�ՙJ��0�[N=F���w� �Jw֩�3��KIN���_+�uҠZ:$�2��ۂ��G���.�ڎ	<N��#o>�H���	!�� �@s-�C �#Sl�Kp�m���5c/�v�/�.���Zeӧt�҇{B4�E�N����@�*�}��nD]�4dz��E��W��["'vm�԰���U�X���:�;���;�Ӭcj:k��^�`h������E�
ٱE����@<�M
e	��Y�<�+�rB�6.{)O���ڃ��2
�-v�Ƈ�V��o).ub�o�O�yj
/�Z�	�W�׊�����wP��s�vN�g@�\�u�i�౦�y�o^���_X(����X


O̬����++FT�#@UZ�UAT"2"�Z�V,,X*-aFT@U�E �Z�I� T�&%B�*AH��@DY�0S2�r��+TƋ"0@�CR�(,�J@r�P�&$�`bESZ�`�k5�bTY0�	�2,��$1�2)\JȥJĴ*���R����*�X,�11�E�dW,m�aQea&$��q�ꄨUd+X,�Ԇ�VC-��e"�)Qq�U����
��QV[T�V�(�PX��bCZRj��Uw�e��9ɑ��)>ީ��<5
V��T�0e.��݂�g{��5�ۛ���ZW�Wn�c:�d��(��w��N�����k z9I�w<��x�Y�?���N��H*��DIǌĚ2�>�*N'��|�i���:���x�!���M*0��=����!�.՟$���q鏶\ß������!m�Ϝtv_�o{��{�8��mLT���M�Y�%���L�%g��C�;H,�;l1*f*Oɼ��'���C�v���e��l:�ST+8��z���^f�
��+��燜�����{m����{��u7����6�uC?SH,��I�����O�T����O����]��t�b���y�'ɤ1��HJ��Q�fE�q�72�0��Xf���'���K��~�\�����������8��<q'��c��Z���?8����CiXnv��I:�`l9��~�:���0��w�'ɶJ��>�4M���1�öb�����je�Ax�2g��W�M�q*,���������|�����=�>�|��d�6���'�+���c����~�bI_P��o)��0�9��I���A|�u�����xsy&�X����bcgy�gY�bq�bg�㳽�_mѼ��s�~��
�z¦��T�H/�~O=�j�RT���RW�i�C�T=Ir�=~�i'�Y<>��>\`bI|9�M��<�2M%C�1Rns����X
M�������6`^z=7I>2K��s�O�	�� OO���SL=g��y�LgP�1��`m �N&�.��=C��hi��d�7��SI?!S!�YRq
°���kOP*N�S��&�m�,��1T���w��C�`ġ�络;�QEJ����7�f�*M!w�����j�Y���!���&>0��!�8��xk�H,�O\|=���6�U�<��i'�T�=��uC�<��g�`O�	�Le�v߽�c�%���˘�v��;����g_�1����Ajzɛ�?$�R�Ü֤�g������4����R���'SM{�4�W��{a��� ��y�v�9���茊�hV�wz�ztLm���왟�~t�{9� i���ßh�3�11���J�Y�����C��
��
����>CĂ�ﺆ+?$���_HbJ���g��q!�K��2T�!Y԰&��7�s�]����]��H�#�+XV�l�k$�P_u��l6v��9Ztʕ�eB��Wy����"^��݆��t���԰�T�K9B�:����*l׃� ��,��=x��止ܖ3��۶��L���y������x��6��3n_�����~C�̠~x� �?}�2x�3���H)?}�:�a���f��LO�|��3��Y�3����x�Y?}f!�������Ag��1�ןq�ݜ���~�{o�}�����i��1��C�vI8��a�<����6�~g�y�X�O�~fd��l��!�O�����$9?B�� ��}�m9Y�X����>�Ӓ���k���1������LI�
��H�2|�ϓI�ٴ%d��oY??$Ǭ1Oh�^Xny����sXo�:�6���1��g����|&"����j�z��81��-���=����6�~d鯹��{HT6����I�SI��9AM$�bJ�H"O�S�U �`T�S��6Ϙbb{I���C9I����)��.����f#f>��K�Ӿ!u���Ⱥ�\�x~���0ҳԕ�Od��>I_�����a�LB��%����I�+<>׺�y�!�q=��2���H�S�%J���VCIKN'|¸�s�g|�ì����������s�o~�������{���CL���p>Ci����g�q8�2~��aPY��L���M$�
�wy�M���;�%@�>E+
¿}d�4�ՊL@�W��,4�4�Ra��<�������~���{����O��R~B��x�w�2���C���SĂ�!浇���1���f�?%I�<9�N2~LC����C�Jɹ�7��q�:k�*�SU�!U¾:~�,�}K��a*����߻=H.&���o�1& k}�H�u����L��O�=q�_�J��W�>�O0+>I�k����v�H/��Z=d�):�C�Rb�O�D{��ُ�f�"+��򝞸�C�^�WŻ���>M!�����ϙ�1>g���m ����Y��b�u7�C�Vi%f��!��I_���l4��T=Cfs�B��
��0�&��`c;��4�ïΒy���y����s�=���?k��߳�Y�%J���}�ғ��?d8�6���y�M!�>La�<_i�C�y=����$��Y�?&����T����a�R�����4x�&�u
���yvz(*_��x��Y�/zǴnN
��6	d5�kklħ3���[��-C��w���]j�ON%<���p�Č.�����#ɍAT�Ѷ��ԇ5p;ګ��P�Z��H����\���k��:����7O�F(�ݽ5� ��l�,�s�5��>� b����}������~�zk��f��%@�W�=�4�+%C��C2��1XzeI�/�'�\v��|î'����m ��������1�Ϭ�d��&!��}�n�'Է��r���^���&T�
b*c�%P�� q+{M3L��Lz�߷��U��]s�l�!�Az����B���%I��LE������q
�2z���d'�����'���E_�۾���{#[�z!�O�4"��G�3����:f���V!����m �Iӝ�N��8�3�13��膙Y��/�4��AT79�u���@�}L�!���.�R��J�0�6�G���W��4Ƙ%]?�3d�	�)��n���ߗL�%�����ӌ���]!�}�	�q��C��g�<T�B���i'��c�+�P1�c���S�� �Hy?k�J�'�1��K�#���~����۾\}S	�LF���wVL�����5`�q*O^SI��LI�+�4�J��g���V�}��w�6��~~�ٷ��VJ��:��d��V{7�&�~@��z�8�mo�\��j�ԨRt��
��;>���&'
y=����s�1��V��%I�٫4�y@�fƇ��b�s�p��$Ǩ{���g��X<���_|��6u�����O��O������-G_��1H���ϙ�(i'�*~d�ͫI��|�*i���}��	��k�i�z��K�N:O]�`"`j���Ax�B���c8��y�9?zb)R�j ��3�w^fǖ9��)���
�֞���ĝ~���8��!���C��y�̛I�*s_�6�'�9��VK��̺C�J����I�3��*jn�f�'P����_��6u���{���$�<La��L�n�`T4���:ϓĂΧ��f��q@��1Ru������8 �[�ܞ q*K��&?2bN�-1����k�9����Jd	����c#�k|��F&��%IS��̕T�q'�^X|��{�I*��>e0*g﹇_q8��};�J���}����VOR����Ci�'��4m�>�*��@jb����F1��gZϘ.X�K��ݘ�݌r���нy͗������ե����b[w�(]�*
�3���E�Z�R���_oqYƭa�A˺�U�U��V��Ɖ�V~�����д[�x�:1N�pZ5t$����؄Of)eb2j��3~��_?}��,��>$�i٫4�U�M��Rm@�e1�:ɟP�&>哉�Y:�x�{�&�u
�a�{��s�`)1�gr�2q1��S�1��9M0�oP�4�Rq��۞��oُ�>޳c���w�����*AVE߰�k4�_��q�P�~O&�SI�3���6�CĂ�y���N���2ɏ��+=O>� q*a�;�x�dĜB��y8�~Z�Pپzs���=�fUE�KF\�C��?)��C�N����?$��8��=ש��S~f�f+>d���a�8�&0��j�5�P��7<�u�4�Y���mɴ1���1Ru���<�0�Ax�3yq���=�E����|nϡ�L|��Y��d���1'fgt�aU�ɳ�I8�J�_�;��rbx�$�y�M8�QeB�I�/�O��.�����7�=I��*>!�I?1s?}i��k9�TJ���K����L}�I>���+'���2(i ����a��0�w�6�YY׉1�w�� �<�{�\��1&��=Ld�P���.�:�O�M۶J��@�S;~�U+��~����u�[��33I��~t��]R�{�z�W�L�4�}@�q���g{���Ԃ��s�4$Ǭă���� /�m>C�;���x�Y�xw�LC�1g��B��
b6b*DVZw���.o=���;��}%!�Vvg0�@�T:�e�=L���)��S�^5���g�粴U���^�MBj�T�vx�Ej�0�n��SK��o�n�����³|@�Y���X�	ϓ�S�%���͖���s��A��-}�j�Z��W��X<��V��/�������Ξ��Xo�J\<6{+"�����j�V������s"��N�ip��3���O�����An{��}z.@�ϊӶ+н���V���Էt���4�@
��u.3�[��o���n9K�t��؉�F���/s���[K!]6c߬u\R��Fp��5�_\7�t��NgR*W"�e'���|o[���*oc�h�}wVF�E�Un�gJ�h�6�%ˮ'p9�u���G1N�S��/ܸ`��:sk"xh9>���	�.7����Z�.��Qg"5�&:�s,v�t�Hv:�7+F�r��	�e�A/��k��r�R�ҝ,��z����I��eL�]�x[ϞA��,J�|��t�ϩJ6�u�W*c{�=�[�b�Q�|q�����;�A���릤�o��;F��:�:6�o.�����<�vU�g�����蔭�f��t V�>��C_ӥh"�f�TˇM��t�jNMX�l�ǭH�N�zL�7�v�B��u����S�u� $;��fx��NR�F1�Iq�K��n5,Y{ �'�fb�ؙ�( )�
]�?a=ݭ��k�nwv�Lڻ��CC�o�B�e1[f�����2MW��~���2���.�.G�J�ۣ0H� B��j�s�&��BW�����O����C�"Dӿ=�Z��=n�vڦ����
u-z�v��iZ��)�P�;"w�4��x� ��H)Y�fZ����+K]��x���Wt��5b�<&�U��e[�\���ԙ��ǲ��.�&:7F�q��2����W�U�+�	��ؓ�(�uw�I��)�|t��A�S�sI\�S��w[�WI�@��o�s�Ʒ%�
�6�Y4�� �>^���`>�و�NJX����J�U�9〬Y*fk��n\�טhG@�3�̰��㰘�>���!���y0��y��\���iX�j�������u����w�t_2�Nvt̸�͢|]B����܀���5�x�<$V�W����S�!��qO(+��G�8�<�bTs���Sθ��:k�hh�ȊU�&p0ky�"��/U�8Uh,ڮuj�Χv|S�!�6;���-=Y�;@�V�h-U\i���O�r��U.P�7�(��������Gl�5���d7MyP�W[ΐ�j\ V%����1�ęم���ڙ����h�+�&aU���;.�+�Ⱥ�6�Bn���
�<ٞ�69VJ�9�D�g����s�e�����2�h�oW�,��iXc�t�k�ߐut���tm>����'��N��� d-R.�꼖��B4�/���������5:�F���w����:v)�ÆXc�w��ܗ��{owp���1E�5d�+����gf�OV�>��]��_1M�x�e�wiM���4fP�V�}�VӾ�un:	y_��7ϗu<����H`�k���/��V6�n��͑�i�7u����k�}�����0���vq�H&�]j;��
�%���d����M��idVUt�1��2�C��X��Wj��[@ܜ�퇗;��
h@�疀���)�Ȁ�茓+E�S�'i��Q�H�]S�]���X]/��7]�ׯI�H��Q���/J���A�=��⓰"�.i'x��c9��3E������X�:uc��x-�����G]�������]���:x`�h�3ٍ�ȹ¹P|���/�0f�W2�«�xX6h��D�˟�ϯ1�^S�5�;����h�9{6�P� Zk���48\�k���8du���2-����9qT����3k[/�uT���-�Ǎ.Sڪ�l���g�"��<���ue'RE�OgW֞�h���g8$`�ζ���{�����
�t(}~��Xz���rŗ��n�d�R�HrXa�cظ7Zxte5U�8C����t�"��U�S�h��:��.�OrN�6�&n�|#��˪nq;Q][<�0�Gy�Y^����ظԻ�ϑ�1�]��k<J�����+s5�9�t�kO���ePVSz���� l����\�GF��.�sn�/�v�l�mk�9�	5����a�'u��ޭi#�N S�x=��YukO�)��[#��8d�1\R��V�c�4��IR��M���˳5݋�o��S�Z�&�¹I����eq��z+aG�u��pg�"�ɞϡm��6f̝���BT�]�U���,�$���a�1�xz��	�I����xj����h|�ݹ3�Kvp�\���YVyJg��.����Q�\ϟ+��F�r��E��CR����Jb�x����3
mʦ�[�v-W#�h�ޙ]]u3��K�rЌ�U2o�I6��B�M��ٍ�f��;pv\^>n7Mm.AȨ��Y�� �to�T9��nV}�|.� �B}d*���Ty%�Q��GUv�"E��q�DY=0�TTFZ��������3�ƹ���3���$��"�>�Ү�e�8c'�7Je{�C�W�xT�{NJH�炧ڱ��x65
�k�z��<��ʝs�5$��+��+e�oߝ;���*���p��	���j��^��g�oh�׶��h�~H��
&����L�ca٨���Y)�ѿ2��t���D�]���	�՗o�\�mhtu�-�ݲ���;~d.�y����J[{��5P��*�'�p�D����^�}����6͝,;Լ�^�] M����S�Ľ}�ï`�
�5���*�lT��|����W����Ѧ{U��b; �����ZF�/|�yk�8Ud��6U�+X6&wSt"ܢ3/k�	���'tr��8Y��t��i�{���<6��ݛ�Vt��%�R;����ŏ8�1N�x��W �Ϳ]x_ܭ�
��`���}��cU-�b�X���W=lQ�ebu���< ����y�֪��F���r���Î��nn�_��]�O����.��0ʤzϺ�o��\�y�4���Lv�H�Б����IH|ۣ(����5���=�>q}@�ʮ�e�����u�8�V�4⃡&ߞ��.�%�N�;
x�dC��Nc��r��h�� ��xh9��zp�c����Y2�s�F����
:���>)�0��j�M�"6�\J��V��1��/j۾�3�QZ��5��ͣ*b�1]�x[ϙ���1I�!:dn�F�s�/U��U��o�P�:��\�6�͍��Mp�\;��{�`S�Y=9���*ީ��.��X��i}�=Hc�ґ=x��9�X���@
%*�B4kF�y��$�h_=��2�Nī�L���H���	�)���M��M�{��WP5xj����a���/LAs*:<����}:c��_*��;��� ���یq�
l0_��M[���WbB�T�u�c$;$�;�$IЏq�/+[�a�o� ��[�u�3U<��܃ڶW�k׀cV��n�t�i�3�	vSN��7[�tCn=���U��
j���m[�ޗoHg�8������6�ob��,\:7���fcP�@��IႸ���jO�5/��-�q�W��F~}����BC�L���1[fܰ1@�.���X��	#&���.:��z}=ו�_�v)��tkl�����ߤ�ᐅ�jX��o�|�\+���p�0]ͺ��W[�WKhʐ���y�n�e����1��`�z�zV��OuR(Vӧ@�uO[v}3o<�M{��tl�v�����c��+�]*�{�,5 	��^^@$��N8�Ҋ��n{j�m�H	7��K�y��l�΁���:^���X���X�k÷H�k�{éQ��9j�*��7҅��0���@Xu�4��xOX��r�0O4�yQ���]ܕ/?k���#P�T�{	x�ٌ#w�<���;�J}�u�Y"����4x�&P��}gg��b��[#�2�{.
����nC�h>�OV}1��)\�Y����_!��7�O�AW����߀_ET��̳+`���ϴS#�M�#��^�ͭ���1͗V��9!����w�]�6R���>ٵ�ύG��@�τ�������fy�~� ��e��y�up˽�|J�G �ڤy��ۨc�ew�VG`on�����J����*���#����t;^)Ӄ�	�ժ�
�|�M��W��]v��X<j�|���ah�C�Z/�U��ܺ�Tk�
u^� �v���sє�+�3.h���Y�ebN.u���w}
#[7xP�Ϸ�B�J���ټmw&{���:A�7�f�u.��8�Uz������v����ʐ�샲��o6nA�1b':�u�M��!*J��u=��3����Ϯ���j��pq�����5�84�9{ݏ�qq�iٯu�3/tX�}�&dQr��J��h�f�T�9-�� kMZ0�ݹM�4�Wg++����V�x~����Z�HkS�mث�K)�Vl��,��x
�:��&�tu(E��m`zu�r�%`E���V}s�N� �* *�	+��yF�.5����ɦ���Xee#�WMn�m������ҙ��ɬ���6��u�˷1gR۾ɜ��X�,e���$�+����zV1�PJ+�ek��^m�Yb���1ڬ=�>���6دV�,en�Ox�x�=T!f�Z���+����ZN_֨k���8�d�+~�J���+�)���U���$wLr���[t��ShMY}"�[0��ҫ�h���+�XwFK�v3�$sh��!���
Peg@�Rlޢ�e�6A.+xA(����#�{j�#@QMp��}a>�L�4��&���{����s]�����H�5��K�gT�]�]ٹlX�Y�"�o>�Ib�s�8�Wb��� �ڹ®��O��f����i����p�e4n\8���T���Wb���0`d�&]+��Jl��X��.��(N�PYF�Σ.����$�B��\��pѧ��ensu��nDw�bB�cB����]7���.OJ�Y� �ӌK�.��{Kt��X`p��94 �Z�,h�9��`oy��w�.Q�9W�Pck �v����ԢjU�+�!�p
�չ��VX�&����TJ�P���jh�]a�F݉,me�@vl*�1(ǻF����jW] ���rd݇��+�a>��C��k ��V��i�{JO�����CP��8Hk����}�RňزB�V�d"	��4kP�B�­P��%:�Y4s���Q�)�Yn�(�5ހ�1�^�l��ɯ�d���03�uݖ�B�S���T,X��w��2��F���ݚ���Q=W�c�\G��]j��Y}���+���*�l�C6��!b�L��ïx1[|s����x�Z���ݟ��%bߦ�v���@z�*.O,
�$#�N�;6��}W�n�a��ε�BP[
�����Z�+��G��T��c�iY�r�Qh������p�Ӻb���[F�~�ߘ�V�*J�*ԭj73Q� ����X[aX�Ld�6����!�TҖ���A� ��T�Q��m�m�Qa*��ejH�U�V�V���P�I.P��YX�Z�+�S��QA��VT�����IYSI�bKKl�+h��4ʬ�b`�Y-j�)JB�A��*��mecj2)TATm+�1�T��B�-�ƴ`�R�Z�VЫmJգE**]\�aUAPY���Uc[lD1V[e��Ub�`�,VDXւV%IX�R���D*�f��G2�b�J%E���W��3֌Ue����TbEc
�X̷-dPV-�Kj",P̸j�奕�V((��j���\�D�Uuj�V:��,.�Q���5�1.��)�[m�B�ň��@Au�����u��[«fm5�ˍu�X�ؗ�^v�U8t�L�:'���cs;����z�(R<�s�u�?�̋?�}��6K��=��j>?�_�\��lL�d���L�]q�	�Yp��s�+j���B�;^���j9�p���k�^>�t�4P�U^}�s�#��_(�J����>�S�q���J�;�[���� K{��Ժ�/d�p�	����ỔD�J��Bl���7��jj�ҟU��۶�&�PQ�����$1�Ned�������IϤH��j�R�N`��4�jǳ�L��T���N��6��m�V}]%�uQ�q:k���܁Ò"f�E�l\�h�>�эR��Sa�xAg�lԎ5
{x'�u�N�:�)+��8Y���Ohhz=�X�Vz��i�� ǵG�8�M*}��w��rƮ><�4n���A����wnY�ڵ�r� �D|���A����Q�l��a�x��C������1��t�a__������
���{��@�x����nx��z�rk]���̇�q�Y�t?�B��	��-�n�#j#dD&�!�J�3�ިS�NV��b�@�͡����|QnK��2�N�Y�:jtA�#�W�����%�о�
M�is΀�Wo;c�v���찡�Ȯ�W�%iKj�s�*�*�_l�x�#pҸ�WD�[/p9RO���n&OVowt�n�[ީ�w�$1���U_W�X��rj~�[k�z�����	C>=QwC�N�0�KK���9�Mݬv���6Wr�}��M���K�����3�[nw6���`�Hg��qp��·�Z�8yf�^��T�!��ݥ�Dd��3�Ps��"���d׆U��v���]��W�Zs�J;��E����iSƣk��ޮ�&qI�*�x���Ɏl)���]��e�"��N�iK�Q�Va��$��˸3���s��>�of������ܥ'��y�@a9b�����c$W�E�����d46����KF>]Ʒ�x`ս}l]v&+' ���3ˇv){
Y����/��|�:��/\����7 ���r�����L)�����v����)�k!;��/0\c�FK�����c��
�����т�	O[˕�6zcd*'A�r�qB6���]idkթ�����T��WF��`��!ͭV�dF��x�=S�<��,�V�.s/�A� �=���������@�VVT����~B����V�QV?w����oiE
����3l�����:��9uu�F*;�oy-���b�i]��u��Gr&��1s�-ޤ`��ݨ�ݒ����15r���4�#<�� Yf>�oB�A�Cz<��g,�#����; /s���K ��a>=]#��l�J^��;?�_}��W�'��4���s��eHZ�U�cWD?��Z(�d��v���ڐ���9�tj�Y��7}̲d����1I�js�������Q�2[ɱ6�	�?s��>�s��&�[�݋̤�LǱ�uf��n�a�*�g6��;M�s�>�ə� 
�J�4Yv;9M�8k�mfHx1�\���W�Y�,���>�G���E�qu�=��ju��IYtl\�G�޾N���(��;���Ϩ����)���)պ�f�]x_����e Nu��<���&���5+|���[�n�8}���aY_ +�k����mq]0F
K`�:��ͬ�-jbp֎u~���˱:��1��o�6+�;� FMaJ�8X<[���ã\���2�r˟��l��C�a�3����i?�Dtܤ�Y����{W^�䔾Ž�ҵ�8��B��$��*�m��z��3{q�C#>aOK�������5���Fw��ɒZ���yj���|\5Ʃe!sUBc ۼ��0tdBt�3��:n�yHf�w���dw{^[e4�<[x�Sf/j�|u��[��{'����˷,V�m���4ȨJxC��7���E��G8ͧn�txM3^�vM��1�wG'��W���j��h~*����oFC!uG����ͻ���*=N�������w��Q�UW�}T2۱�����3����@V����f��mSUؖm<��FNCT$Lᛮ�7:�wsC��!#[�����VDt�2��2�<��K����%�;�Yy���獵U����f�v�Jng������gi<{t�1�dO�
�RȻ6"�v�l^ ȉg헝m"�#��^��� �R%}��gfݛ��M̮��]�ަ*3ګC���;'i���: H�ߥ��o��Ƞ�5`�����O[!�G��ᢕ_��ؙ���,<����"τ�����	}�@���/���C�1t�Tɶ�r��NLfn�{V��U(�A�
�ӳ��u<��[g�W�CW��5%leBc��F��":��]iD�6�.����F�aJ�n�X��"�!�GJ��^ ��T�)��}�e�7&qJ�y�5;��N�Y{@;��i�];���6��u�*��/,�B�J�󭴊�����d�DwK�K��mRw����Y�p�{M��]fU�_�]E]����޳��oTf��k��)`���O��]C�Oht�J�`��R�R�u���}�y�C�ɖ-op�$t��;�����-��䜭}���f/���b-l9ٳ���9&�M��\\q�f	Ł�b�{״�3[c���ꪯ��#���T�R��N8�f9��<@U��F��(Yq����^�C�
�:χ��ƚ�~��%m
�pl�,�����F�|����i
P7�ߝ���<�;V��\*��f9���iϗ+4xk�'g�ZY�S�\�����*�96;B��&�=�w��b�.wSH�� ��FLd�"�%7�*��Ä&��rG���[�:V�d| �E X�����e�d���d'��hdP�#s�o�1�l3� ��ڙ��]�*\�	��}�-���ޱ�_���b
�I �KH�DC���VeN�#e*�\�4Vz��@�K��9tϬV��G\�\U������j�쇱;�9�~�F�Uᕪ���T�N���wT]�(0�j��B��)*ߜK@ȼ�av��@C$��|�F��	�C#[����W��T	B�Q�(�.(B�{�a쭫��Ƽ����T��<���
�d�3q1���,%��U0g!:��B��n���s���Wi�q `�ʕo�e�*-T9����0�
vg���c����t+sWBiǣ�m��L��{Q낯v��;���?#9���0p�B�O�pn��7iV��?z*\����0y:`����M÷�x5^6��s��s�f�3�v[���^Tn
��{���[�j���ݺzu��d.�M8�V#Q�>�>���"�Y=�)dR�]B#?w\��r~GI���;>Q��/I��B�S��4�tpj�/!^�t�&v�
ce�7�3�j[����w�~��ِ#_�v�Z��h�
�Zz���>��_
��)���:�>Ξ�+&���T���Ձ�W �u^���d�˅A�=x�u���W@����$z��Е�2 ��Q�p��%�,bW���5]�Ϥ���P�|hǢ��k�6^GTm�ao;���v:ZǊVԧۊ�m�J��y=�����4�1|V�N<����h�<��v�>�Պ��/�o��B�*/f}k��+�O���+;�玂�̉��u�<�=Yͳ�T-�D�"�����t��{MpwQ;<%�^� /�>�7����\�򋓻�'�.wWvv��v���>�$��B۳I1s�U	��aM��Z��/F�R�[�)1=+M�o7���ҷ90w��G1r�ڞE<�c3ְl��8o,���%^����s+�. �@�k̄ƫk>���Y��]ƶ���K���,dVJ�ݫ+M�~��i8��ARA���Nm[�[[�9�0n`TNu�WXP�z�ӣܵgln�ѩ��1m�Z�zA=�Nx����i_e�f/�];zY�%�E�����Q7 �-������d8)r� nk9nM�$�U�`������Y�I�DDV8���,�L��}aL�Y�S`()SR�)���:lh�=�XSO��çWZ�g��cY��l�
���=��˅q��S&�Q��)�BR��o��{��k���S<�'L�[��b�������`r�s���\c9𪀌rO+�>�oy��d�.5��:�U�|P��\���B�q�T�V��K�r�����KGYn��;��ϺHͯL���׹�S��A��L�_����1`"7*�W�s_�v�Ucx�V��|U����5VB�NFOC}x�§s0J�ٙNo,J��LM@�$᪨�ݛ%��\���]iy�tۄ�O^+����\j�V���zew���7��ό�)�Ե^�
u�]��<�
0=�κwYjM�|�2����<*�#�)y���X�B*�]�l@@M�;T�ǥ�Vc�D�3fP�@l.���f�CWg���_����V��~�ᛲ\���=���~ޤ�:�������
{���pϑ��n�
OӳZ5	�f/��*��o;4| �_�T����Uw����O��˓	�P7ݱ���6,��KNҸ�9Wu4	���~�������tg v�笨��j,��,,��y�4,:�7��b���B_ȸy�zJuݽr�����-�;��2ͼ��Fh �����ɘV�_3
�l:���_U}�W��w�K���|s��'
�m/C��r��Ex�89r������8��Wlˏ=�=�N> �u��|�g�E���t�qڿ|��vĲY���������Iț>�����\/�1%���u�<d2!�j��1�AN���`�V�l��*�]M:�_8�T�Q< ;)�}3�z}iq�	U{Ώ��U����!:L$;A�ʎpD�Y� "|�:C�������.E�cՏ.��Ip
���2֎��͑��������Q�J�-].�[��ΐ�U"��[j�VO��2� 3R"|Mh�]x�e�@(��C^�W��&-�R�فU;/>�p9b'�x��c>ȟ�D�ThF�.օf/����j��ftu_V��d����I�pdOE'd����Q�g�ش*n!�c!D��"�f���5es�i�s�/�kAP�ډW��sC"����/�-�ڙ��yb���	���L�<�y���e������xу��,�vx��k�����m��9�C~��2lk����A,Z�G�T�/� �L3�g7Ry<��¤�����֔l����=�C�=�W��V:^�*v�j�U�x��ͮ��S�۬N�7uL�<�$��b��=nY�Jse�uv�9*?������cט;3�x��?n�#�����-L^:�Tn��HS�Pw��6�Ԧ]=������݄,��ʝXPا�����4�ں	���+�x��Eh��vEPwT^�,��p���'F
���������E��@�/o�J�A��ٟR=�"����]��V��WN����c3���wH�E�3(�.w�Jo#�_��%z�����.Ӈ�{\�Ws�U�?%J��ި�Gݼ�ެ�VY�8�fN ?��@:��[���B��0���@X�M��c���'-xX}�����I8E:�܍��Y��Vp��9��b9�w���ӱY;�^��[=�7<�R�De�K���w�zF�s�εr�pu��AO�}m�Ed"	"��Q��n:��jןb�gLn������U��ZG���/�ee��fsc'�fP>�1��q9�>�"�n��	��o�1������d�o�Mf�5�k+wם�V�,�&fw.���j�)s�j���>�<#�=���6q�u�sL����}�2��K(F�S�:-�

43��|F�񭣘-j񆅿R���O�t���<"͓�}��Yv��&!�t�f��=[zox 5�wn9�r�$�#AҖ��+��s��ژ���P��w�؁w�C{�7��i�{+:�kA@�����>���q�:CD�Y��Av�9����Ȅ����O��g�F��s�DH�hY�)�L����;�]��4!�m}S���D>F� �#�	�"�Ȋ�2�J��愝2�/@m�`���t�	.D�]Y ˿����*dD)8/&��E���U0f/;d�2:p��k�v�� 9�[�oۡ3�\kF:T�|�=%S�^!��5+Mp���w9���-��e⽨r4g���Uk�z�S��:M��qأ�^*-��A����ǈr���];˜����?@��oK�Ϗ!�P!�y׋�>��ّ�L�ϫ.;��Z7mֺM-X9Yh�/k��8A�:��zr ��r��ѕ�s�|�A�P6h^���d���(s��&��(-���*Ҝ��냑�l��������`��r�U!.Dl�5w$��*(-�I�:5oo��6�g�K�l�F�G���ZǊV%���"�y~.���LO�Y*�ƺ)�z�RU�'n�@FOK�;q[jw"51[��q廋���^����c��K�zU�����8�@�V�3^��x�ͰδxAҳP�,���
ԭ궜�u�[��o��`f�Dz����L�;0#��_v�M��%��w``v��0�!�!J	ݜ�`��w�:^v�72�x�Wu��:kw��l�Pk9�b��sd�WS������0��9��d��c�xq)P�F���r���(�b;�uѥ�άY]u�]1��VF�P�VR�9!p��X���D���Z��2��ǝˎG�\��]p=�a�\['�tU����_Z͗]W�mȎ���������<v�a�s=�)��Cu5G�|�nA��R3��'�ER�޳�z�/:˸̾��ю��|Pw��)rã��☎�%�FA��<fK�qv+Vᬍ�[�����v�#�2g��c�A0�ҩ3����;�ktaN���iza/%-���^�T#���uH4N=}�\x�di�	3gj�� 2�V<�&k�Nb��ڲJ[��f�ү�%̰'n֥�hj��k+��3�:cG�X��V�鼖4��d���������S!��ٻ*v1WөN�`�')r2�v�K�4�j�]g9�T�v�H���%4멪��y�Fm̈��H�¹�le��K�#��3J�����{o��թ����"�iޭ�],�e�A�ո}�h�鷌3�D����m��(,��Yg2]��3�;�<�m..\�2��H$�=�T�m�۾�!ۙe�<���tu��Q&�]����l�Pc�`��ͧ��Y(AW�t°i(�-q/}[��ܽ���(�1�_n�M��MSy��@E���kZ�Q.Ӎ�àh�u�ط��Ŧ�D�V����Ի��@�w���rd��>"�ſ�ڞ����F7K����I	���4�z��^A�Yo�`��j�<1k�\q�y��`��ۺ;��Iw[O���#]n`�$� R�v.���P�uċ�h2�\(݇Z�EA��l�'d����Z�cPY���6z8 =W+��!43L9k%�i�)-��;qePz����xg�ʖ0�v*75��g
/��H��ĝn���K[�!ё�Gn�p��s{+���2�K�A\xKYT'�U�UN�e��n»��bk�U�00˄ hخӬ�4����%*50�!��u��
����|"�;�t��N�]�`��C%������^���Fo*�3����9�[����[Z�cKne�/pۇd��AuH���4�ޅ-���L
�1]9gI+�{�A�+Ws�}��⠋���|+r�(`���vq���k�N����V��(���8�yCAz
�@����aӻ���1��8ie�[���v����]�w�M��H
�ա���|�mW�I��_]#���'�A7Z�������i�k���>�o���i9:͡[����?{�}�1�%D��-j�kQE��R�ʭ��iX �DD�0QV#kJ�֌�E[[B���F�(�*�����(����k1�mEJ�ZԪ"�ҵ��Q���b1jTD��,[J*1B�b���E1�S-AF�Pc+[mJ�)JT�B�*eh��%l���"U�UT���Ĩ��UAdKjY�Zc-�U���%mUEQcV�[-�X�P[lPm�[-��"����*cX���PL��c,�X��B�EX#[mDU��+E�B���.J�l�H�����P]5����X(2���QZ�EBڨ�eh��(5�m[j��ժ��+l�j�"�DR�E�TDZ�cQ������*�*(�(�6�Z�L�P��)\��f�uef�mb�̢�E&%�YB��p���`�T��mD��Ѻ��Y\�������s�W�q���U�{�wl�k���o�+�'i<�%�Zz�p^��B5ǃD;�F<UwA7��h� r�n8Ε��G�G��Av���s��[�����d�|�V��Z@�.��^ث��Y�v�x:���q��)���8���m�Ze4��L���1j��{fx�g)ܐ�1B2c��;¦��S���Y�=w���ֽ�M`�W��j���K�F�.��o���gԷ>�+���m�RZZ<;��u�¬�
y#���d�>��\t̔ՙ	�V�}����6 �r��,�3����N���}��������z��_(΀��
x
 )�YL�=A�b:aN�:�O�V���m���$�X����p�h��g�
���W�ƺ�{���($���e:M{N�Yʴ}�=�
���F͐���AO��J���F�C��NUâx]/�.dr�*���T�
Z}d*d�V�"`"2*U�G��g����ag]�����9λr٤J�����K��xf^��ACƼ+~�{N�H�'��o����f���#5$L�3�Ռ��)��.��L_ND6oa��qU3%��iИ���+������E��X��B�N㓝�֓�d��X�e�\���WWZ�
�<خ��o�gvc��K�Ә�X���Y���U^ɔeiN<���n�d��H��5(�jyv8�-nR��3�,�
m6���E���GPb��I��h��;�UrF0�꫼=dN���Y������_W�_UR��;���o��k��}c��G�Mx���|̮�X��Ȭ��`ƪe���<Fu�yN����ς#��^'2�
��p�R���+�N�)<����˿��Q�@' ���l��cә5���@�˫�@����=]�qXb���Yn� AOh�^��4񊣺:����(�7��0ẞ�����T����R�Y]h�1�j��]48hƣTm@p���f9��3p��{��u���v����/ir��W��H��u��C��ds�οZ�u��//om�e���C� 5.x����U�=�v���5��Q�k��>�S[u������b�86�����*5���������D9�QNc�4��T�v8]F-M`y������ TO��Q�HC��UBc>+lއ'E�t�H\՛͐�3}��d]B�:u�s�fՠ��
�<7�G�h�N�6G���3�KR��5F�J��]��-V�<�7�/��p�n�K^|g&���)X���M���K��|{1��]���"�"�������v��Q�R�o��؇^8�bE����W9�_Ƀ�Bu-�ˤ�������v�t�U����"�݃z�K!`�tU�S[��{:���}(p<���ۗ��G�{P��P�L�se]����b���ÿ́;O;���JHy[�&��V{��#�Չ#�if���U�S�[{���õ�L�'�a��6������ĥ�f�5�vT��,E��:�m�ysFA�����W6��/s���>�f��鿘�*n�2Ȗ#�t=ػ�鹜��|�(���Ϋ��5oF�C�b%_�nK"���c��!tC������M`\��S��i\�I�����Ut���3�R�ѻ"�@Z,�/�l�9�U�:�g���y޹�w9%����u�#H5�e�(�S��o�TC�ؼ��u�m�g\�����9t��5��#>��/~���.�|��a�kF4�vڨ;>��c��̌�ʣ�%����[O4	~��Zn��/o�J�&���ё:�v3!�n^;f֫��HU۸�`��
�� 3O��}�mv#g�^�u�s���i&F�ZyEr&��I%E}Rv�P�j�������}j.۳ݕ�L�u4�3
�����w{'4IB�/r��:�X���׍,����r'z ���Grw�M����r����c�����q��ef�������Ր�&M�Z�E@�Pp�m��a?	܌M;�q&�\;��pn{Y/��.�������[�&?Y��|W�+�����T���f�䩩3���Yj�9;n��p�?EU}UU�Ͳ�N�ǈ��Y��B����\����Q;=x���4�b���fs�"L(�{]��+��]�PF�X�#Ga���\F��Va�.P��
*����{2v_ Q~��i�g���H�/�M�)�I�v��{m4Df���>���i�t� ���H�?b/բٷ�vC�K�]{%-̊�h�$9=�p��v�hV�oi���xR춋3�R�IY�U���.K~. �s7�0��u����!�u
WϦ��o<��N��j�x��mߑ�m,��&|{��u� @C������C������%_&
����q{5��m�L��oOuҁ�@{��@tW�ÝEH>�V+�ٓ��i���EdUt�.�)�zM����2\��ɓ�
������9�D	\kF}�d
�Uvr������ֹ�1'�ʬ�Rd��5u���b �2B�L�	.���F��8bM�]��:/y� V�e��N>�f{��ɿ�w�k�r�o�S�.�b�O�ӛ ϒ�������|q_c�<�.T��V�ɷտ/�	 �5K�
�Z3tU�a�������XTL{ܷՑd4t��������'� +��f^���>��w�XNe���Z�ݛ���u��NT��ςW��V*jNޙ>E�(^�bƸh���]���a�4>��:����V��$��:Ҋ#(�W菾�"!��Ǝnsh">�s�B�ާ0�k����(W���tݞW bP�@��s�lv��cdTnH˕�IX��7�M�x����
wC>Y]�S�>�]۹�g�J�I�:�U���:�LR�k,'W�v\~UtJ��#ӗ������Ց�O�VA������+H@V`/_�Nf<�������R<��$g�x��ǆ�+|.Zb��^̪�Ca�S'��w����l����-�0�鋃�;����Xb���������蝞ү1e���#կ�W��$���V�{�u��12�z �Z����f\US��
)^wX(�=�2��DS��5�U�C���{�X���I�����F��]�	�pg��v粖��9�n�\O/&1��ïC�.TYꑏ?=�*�U���x�j̄�¶����hȂ��v93R'�Y�\�H�]�a�����_�����Xj�� ������Ah�� �n��6"zaOp���|r�~M:��ݼ��+�G�Mm=�pTq����A�\=ƥ_ 4v�	�#���+3��V+��s*{�\��g{E����_��_�ME
��DE��د�C
�KS�^k��,U����DVX���Y��i4ߵ�-�	P�U� �x{���D#Yj�jh��U+�{ZC]QTz���c�&�� ��&�z��b�|��}/s���f�)aeZW菾�>�Eu�2[nq+��*���Ӓ���@����7�'�AU����&��k{N��kg��L}�qS��i�BKͼ��ҕ[�P��r|�V��|O�1U��*�ԙ&gTJ̄2W	��EQ#��5y1�d�ΙY�v� �p��ʨQ��(ێ-��=a�SQQm�X��2V�\)�w��u]�q��@W�W*�q����[m�:+p���Â`z�p�tW��5�x���|̮�XAU3|��&�e�d�_Gv�c���{�ŧ���I[�Iܲ�V�[��K~
�)ef��{.�4���w�o)��$�YЪ�����ᐕ�9_[6eP�@t-�N����<���^J@z�k��/��]@3�J�p]��1���וsM�~.h�sk�^�c�J����8��~r{.����]1xZ��ȉ[���C��3ݓ�^��,�GC�5�7�f���1��w��V��s�ePZ@�L��ζ��2�R��]�]O���A��6���-Cv�� ����)G8<B�g��s]X��޿W^`滖�S[�Qt�.��)�]� C:��(坳���5�����X�v��c��hH�(���ά�b�>�R��۸�2�uekrW�����Gp"a/DG�D}��WY7h�38l�ԗ��R����O�5~.5���k�;�'�����S��*c� r��(R���k�Wħ%����T�L˓#��3��F�!sUB`ӫ�@`�쫢��1�w��+����9gӕh�z�_+�@�I�ю������+���R��L���d�����*+��ܾoi�����r_P��h��.u�}�)d���r.	�V�-����ϡ��|��g_#��4�wh��3%�>I^���dN�[�O։2r>I�7� �ae����,aM���@�H��T�ݱ���#��SM b���9�}��7Wp�ygsY;؅)�T��glBvd.��=���]�'9M����N:��Dv�O6ȥZ';c�	ɚ�����+��Z�$�=-�aT�^n�P���\�������w	(gl;C�l���F�u\c�KQX�iD����_V.�d}a�[�5:��	���w���A^ž�r�D��w*��u���ءv9N���3U:�������
���G�M�.��f��m*��E�e�"l�,*0v[�|�9Y�a�0K�@����4v��UU_W�2�:�8��ԏ>޲��$�j%��V��7�m�-���>�騺I�{�RK��zEF㊎8�@-��!����v��`�U'��6��]��p�ι�n3�f��O��]YQ��9Gj����G���l�����0+0�#�'b{�-�}9Ѿ���q�ި��rq����z{��e�P;{�ޖ�O�����L(CuP�Z8�ڬ�U���ս+�g�,{w��MU��ܪOi�v�/�>2n3$���x(�j�l���SEtUn��â�'Oe�L��k��e�����> (��4C�齐���3�.�{���闟pkrI�m�b����*ܤ���nck���z�L��)nj�_YL�*ic�v�jt���ՄT�/h��qQXg{��z
���JFn1���E�E�'>NO#r�� y�\T�qU�iI��}��y�8�u<���cX�e£�y����]8d,�S/a��f���k��� I�nGgy�ʓJ�`{F7_u�de����ﴊy�a-N
�)��F���Q��wi��B0(2�m��V�-�A�ԯ�s�3-��u����}���}��Jo��#|�д���0�\J��D�s"Q��ҝ����Ⱥ�%p���s�:S�%��1V�0��	T[ɨ�DE�G�Au��R���̮��s�y���v�}��m[���F�1���u�nي�NL�vŮ�s%w*U�/�Q��n&�4r�rd켤��^|�CLd��!�&n:w�]+��g5�#x=�U5���ܞ�ar�?�>*��u&�5⭷�h�=v�6�7j���3��f�9�7��]��׏��^w�ݷ=�����1i
0,������] �V��O[������Ϸ[��/m�W~ci���ކ�5ײ"�i(�Wy/�uD>ΫOF�=����.2����[��M������,�(FZ����f��){��m����8���|sPm�ЦTM$5�gl�u��f�4�'esr��ݱk��==�A1�$�@Y=�@�B��5�z�J�����ؑv�G�h�t�c��fWl�ܨ5Ճ�R[i錪X�e^���K��L�ˣ��mvq[^�R�BNn�ɠx��65 �yx0m�ь:���|1Ƴ`�Ô�v/P�Ll���8��6�z��w�:��̊�*����}UU���5�M��~���h��Fw�ѽ�֯�!��=.B����Y��� ��z�w�j����Q�ŧ�Y��ry%#���4��n>H�o�Lt��zs1�	����� ��@3��i@���aJ�,>L���%c�r�� W5�6�5'����Q��,o'�+�F�TqBFL}���!�u�tv���^��+���d�O�j-�Nm�ba*�a*����k��h����:,��8�%q��2i�)��?cɨ�H�ވY��G��Q���b�hޣ����}��O܉)����n�'�W�&��L�U�o`��>ّ]�i�p#}�R������1�ٶ�T>AA��0o�޹3 ΂�ٖ,̽Fzl#�-vl�x1c���\��su�x���q̋�1ڊ�#���W�^}����R�+�+���E�o�;[ɒ�5����e�T��1;�ϟgE��:�{'R���ͺyLi%f$�<�˵�[*5��^gtq�}6�J�
�U�vͷR0^�z���w�8/�'Q�9�[Yy\��3\��H:`�jqZ�<��P5���G*fvtj��R�9���-1�o�'ׯ	��/C6�"���$�4�T0�)5'2�Eݒ;@6�f8څ�n�嚌�2���YX3��1Q'C��t����9da�Vb%��/��{9��=� �vZ�Y*�-w �-��5��<b��kY�)���=��,��螡�^}bL'i��+v3GpU�IM�BW�ME����m"�x�1��r�{�on�n��N���=�.5����7P���[ƀ��g(�ZC��Y{nv�Y��R1��*e��8��I���r�X�\��۵z��	}v�"q��_ ,U��I��'U�"<�G7Mm�A�^���h�qٔ����cX'�n0.�
��׸��ooW5����W;y�2D]A���u�1y"������N����r=lg>�%˛�p�>LLV��7���u`��b������Ơ��V�v�!�r�Bos�.��풂�.ݮV�i�i�ٻ-#K�v0��r�`i�z���@(��Q{(��w-�Y�ppL�j� ��«;v�޵��S���5�����;���)A�Lo>*ٕ���Uk�hGZ�J�[����e���	�V�AH�Cvn��Gn�sP]��m�N�6kdpCM�5[Xi+��wpn\�A�W;��[���dk�H6��V{�^1��*��Ad@��6��)'_t���k{�_�g�Sl�;���bK�lt�N���$,Y����w|�w+�b���O��6�����]�u�������am�^�KA�ҶX��𔉡��QsN��v��ѽJ� �?L�s��[p�h����=�1u�]N=�����Y�Be���H<xK�(��֛���wnݞB�s��Gs����u�G��|��V�2���p�M2��;�R+7��7j�ݝW׎qmV�ш��fWĶ#�#qvb�Q�	w�n=����
6���R�L�wE���
��&I� k�A0�I@3�(Efh|5j��z&�=u�{��m]�,ZC�#7�hJ�=e��b!FMz����ɛ��W��b��ѷL��i�N������x7c�{�Z\�bJ�Z�ʹرIt�D�,����c��Z�=��O���4���NbƹY�Ec�0N;F��z+���5V*u�{��9�p)���-Z�1g�H(�w����t�3y�5l,\����;�����"��&���/0�b���6�t6ҏ���ed +8b�3e_l�""�N�z��V&�IF�Ǎ��c���#9gZ�T�H�}{E����\�㸻Y��V���q�	Jsi`�*t{]SZ��c�<��t��vH����ﭟ����[V�U-
֤�9J�F(�J)mU��V�Ķ�
�ը���,G)TZ�U������j��V�(�-j�"�J�b��*$*m�iH�墱F(�S���U�TDEF���̴X���H��0f��11+k�`Ŵ��ň�Z�6�-����Q
����:h#����c�j6�PQV��QY���%a�,b��(��*1QEelDH��V�E�ER��R���R�*���1�VV�q�����
�QD�EmQ���EDT�1��K+)Z�h��KaQF*��PEFУ[j
�jb��m��fQ�ffU�,���M4�Q���h�*����f2�-iD��`��
�A��PF�X�+cAdU�E��1U�ȫ��EVD�"ţ���U
 *���Y�;	��Z�T�(P�/���tp[:�HR�F��+#,6�����)�v�)]�&gV�ýL��+�G�G�|���*:����%^Ҍ��3'. #�S�<��zQ��g�sؗU������y���O�fK�1�,[{;s���Y,Ȟ*�nVms�q�]2�"�ʤ�^*ۍ1��A�N\'��A}��鵙�rwXz�%s�h���&mVo+z���F��o;Q���h��tڞQ�a����{�Ӯ���h�����x�a���ÎK�_aM�>l�Vlk��ǜ���Y����I9��=��_5x
z�5��75�o��f��G�z���4i�U�|��B�Kt�����;�=����ޘS���5�r�G�=��o�[w��r�
�9��M�=�S����z>��;qq���->�K[�{^�:N�#Y��WY!��mԃ.u��vy���j�y�DK/5A1h�a2s������d��He�ga�H���ea�p��4wV�>��Z�Z���ޥ��{��І��V��BK��ܮ�W�Y�l���Ig�L�_ o����y\����~�Y0���Yk��|;s\=!��\6��*��+�zk]:�w-@��P�Sz̚2m_S���}UU�=�����7Q��>��� ��P���;��5�{^s��bw�n�
��K�-�7Zq�̸���E��ۛ)��D��S#mUE̡\��O��9��N�C�V?���2�7�R��v���81c��X�5�ñ�t,v�v7�Y�\4pn4���a�n�*��Ȇ�;�zi�Z�=���D��&C�ҙU/���5��{o"V��7+s����CmR+:��ޏ��>;��O~+���;�6#�y�5at�q��e�[;������KǷz�#iOv�k}C�߂�h��@���cZ�z����R���/Q֭�{��~v�k�v<��8�l6��h\v�)��v��~5=O"��<]��D���A��^����Ù���8j�φ�v�T��E�V����iA[k���'6�=��y���6\�=o�mw\'����H7_Ǡ��)��<�a�0̞�k���t�$�ͮ9m�c'l���;���3��Wmh�j=����y���{��jճW�C�/�f���P FU�:.�]���ZZE+�f�w<��3���J	Û}�;ꍝ̂m4vN���BQ�S�B��tֱ��gO��ﾈ�I�SZg�7h�q����M���V.�}���2�
��mbڃ�+m�ׇ�%��YG�0�x闟pkO���{�z;gK7�kv��^oY�G�WA�7o��Q����~���n;�vF��yy0�j�tBl���6�ʡ+���'a+�uQ)��^�.�V�'bZ�90yL�P-�����=�!���j�l0��	u�J��L�#�ѥ=�}
��vA�Y�Q� �QHa��{����A]�Auf�<�5S2mI̟���>��$�	Jʄ�Y�o>cK�`�{6�z=p-t��d���iA�i�"�2�٭Gw���������(g ��y��MCNL�2r�l�ǝ��^�1yٸ��1�]g'����-�8�o���BwH�0�D�1��Ž3;�m���3uf��t��7��D�,�=L�K�ޝ#F���yٵ�g7n`�=�T�(N%i]q�E�8����U�&*,���u��{yr��{%�3��[�ہm��!^�Gy`Ө>�//�hfBS	o�s�������Fu*}d0��1��.�U͝ef�[?>h�b�%nN�Wt�f~������	e��}e��;9~il�d��{Eb]�z�]�8n�����X1�����X��Jv �gU��K��}�jͣ�o�ض[�(��2�ҽ7������\���=8�w<#�h냓���t郜����XN4G}���5.�5F���8��K�ϓf�=z�u�fI<q��צS��M��dwek�d��6�b�\��8VMf�N���5վ��rF�U,�Ϊ���%���J��d�����K#J��-pkr)�';6���hֽHd�9������=��
I����W$�Z����Q�榖��V=�'�R��#e,���'��c>���&���I4,°Nc�޹e���kC!�I�4�{Cm�uq���*�����0#jމ�U�SO����Lm�k@��9�zeg�>�W�j"� ~Gn>�:�(lwz]D���W��h"�z1i��m|7!9z�J��of�'�u��CƄ�>��e�ź[��o1{׹8��k�m#ucb����A���(�Ķ�{J����ٗ�u�u+{9�f������s��(+g��O~�菾�����&bEt�"�{�(���KLk�R��«u��.���X+�WSUn)�ns�cx��U���[��ݑ-�I���ͼaC-���<��JH����
0\�6T���ݮ���_}~���yJ޵������Y@��ZΌJr����Eê�G̹;��Gc��b}\�M���u�؎x�Թ"Y}�>��)�:���.����v`�Āw!Ow7���$�IH��qA��b�k��x���-~���E)^9�r��YV^�7��G��^o�ұo˩{Z��;��'��A}�Κ��;x#���ŰE<E���ȥ���V(ĹV�m%8�������o�^�L�S�Ic�x�̓�O]Xm\`ׁ�ZjMl%i���j[.�g3�QǊ{�������I�@Fz�_5����j��%��T��a !���gl��&q�p���A�iయ6���ع��y,j����w<1�tv��Հ�m��B?t��hȘɈ��٣�����xTF1��8���Iv�"Gb[��������E�� �+4Ώ�ږ��7}�K�ӻeC���b���;����Wu�r����]�C���'a�A�˥��G;�+����Ά�;,ݬ���Bv�U�i������қ��6Wg�T�qS��@A�E?�m��ΏB[:��1�V�H�̞�|�\C���9�zn�9��77�Ot$�3\M�!��gҋ̃�i�	��t��;!�';���`��u*8��T8%ɸ�klBUj���!Ή)�i	|_�L^�^H��b=߳U�z�W�ٴ3���f�nl���V��:���׳Q �=�J	V��M�I1�nȨ������r��_
b����poRdos��iXĜ�Bjϕl;C��܀�M#�Ӏ�a�PK�u��mƔ*4�)�Ĭ���U�p:��ܬ�����n�Xi�����+,���J�p죲i�M��zy��Q\q�j���q��yu%)��:|������{+/��A��-�OIgϩ�y9����]u@1{G�P��O&eMI##�y��[�VđX�ؤ~�+7xSpj*K/n�Y<;S��}{"�y�!�l��n��ø�׌�[�u
�u�Z���c�qv�0bo�G�}�Q{!�0����D%'$�ѯ.1�������q�fe�w�D-���������<;y{�t��Ԗc��v���Q��ƨ�|�p��N��=����m��R��Z��
�e��G��'����Y:�5�*X���E�� %�.Um;xw�[�i���Gj��rx�Y=q���	��'3Wc�qBg6���Z�g
m�׌�@Vu���`0�q�P�j)�3ԋ5�:褣>�']2��|�"w�oj.�q��|���P-]l�3�G-�p>���k1G(���i(}+�5��.$F�6np��Vs�|q��鄪'�+�U���E��i��H���MLt�3QY;�Tc:�y8;CUn.��{��!_7L�+��	Y)��Gr�=�=�X�ݪ��޵�����./Γ��+ǓiLTv�o��E�Í�'ۆ��I!��)���q5j�r�x5_bb��%����;�7�(ތz%�c:��{�FǬ�sO�`�u�h�Gé�L����������5��v��O@�]���$�]Or~L��Xx.ǂ�yV�H���x)󦔖�w���ij�a�?}U�8��o�L�G�K;��v&����kc".��1�p�o��5]8�7�sw�Z�G��ٴ�ʹdE7������	X�I��aC8�a�&{�Bb�8'�D�^�f�$[��=���<�|�{5����|Ě��7L��Q�Ӈ��5�M^�S#���/>�w�<֍�җm�ˤn'���9N7�a���ygP�C�P^[ȓ����������c�ͭ���:�
5�kw��?v'^�L�'���^�+˞oy�O[W�l���E_ ���bYhq�.��J5v����sqt�?w�ߟ�K�{P�Z8�3bW��=`�����ߜ3չݴB�J>>������(�zv��b���������r�3%8%��6�utg]��k�J]��3����;J�
���	e����:g��^�j��2�����[��$��fS;��f�C��������Noh(]��6ݛ�w�닶�d<��<w���a�B����f���I�:oEE���`'z]��eq�z�l����DUf�xm��qjgQ�KE&�طf�1s��))���9Oꪪe�<s<���L7��b����!@5:9�'&#
W���GJ�v.�\
�=gb��7z��:���;c]i���L%Q=n)�JFf��{�7v��JȾ�2�+g;\s�Ql�)��3'�C���ݤ��Fa*���+M����;'��I#X���fF��������Y�s�f�K���;5�ghlJ�t�ܿ{+��v�"�-ϥ�)�M.��sfIo�-��I���<{7���v���g��#�U��j��L���	0�k-�Uu��}N/_O^$�_F�L������Z7��s>�!�.^���t�W;�M>�ju�鴔>0���&��'e�]y�f�j�*]�b�
)�wl�]��-Ʀ�4�s�����w>앖��jn�58�M����U&��Is�[�dwێ+�6���`��wC��s�`�Qeåq��9�t/er�����Oz�����Z,^U�8r���·{<�k͸�g`��}���!�|�&�4�R:�v��w�Ŷ�/��c8��̠r(�=XV�"� ��J����F�ͪ�,���fW^��nwk��zq�[���V+)R�W���>;E��+��K�MuDq9-����:obo�:�`(��t�/;ڬ��ڿoGYąʏ���Οb�k����K���f����U���M���!ۆ�m<��3{J���T�;Z�\�X�2��V�r�����4��l�̀h#=t�_5q�����s�����H�u��;y��w"l�x̪9{����ls�P+���H�ht���kI<�����/%�e�pgs����7q�[ϧ�mX����&Q�L�{M�Ev���P�*QKj�_Z|. ��3'�>�I�rc)��;���&I��n/�����,�}(�ϵA����d�єE�=�:'I���1�b�W	S>�k�سU��y�(��M2G���ѧ5jަ�,o�o���.�=�c͠���#��3K�6S�qR�H#0���Ÿ���J�:�p�N�Y�S��z���-����ɏ�t�ܡx�m{W��t5+s&_;�F��e��v�sK먻P�@su����,i�<#��ֻ�6<��c���}}�˝\������#�N�z��˭���+��`��`v�vq�w�}5���c�2���:#;�iy��TzhC0eC�/�U3y?��Ļ��V����]G{�/���.�Z�܂�E"��{���;�k����E�
�
}lQ�s�}����xf���VXK��;�L�?T¢콞�
��v�w�u	�+�P��A�i"��f�����E˨����.�P�j��ϟ�@��� 9[�ޚ�lbt�lC��8�Е9�.�P�4�7V��Ѳ��Q�D�v�fm�t3�f�v����2�s��Ov;V����=7����v��s<`��TGfّ���N��\���Wi6��@�k\%`�!5/�5efu�̡J��0��j8/�S9��zF.�H٨zͭ��S��S%_��c�{`��C�������xw݂Z&�N��m�J�n�r8�fG,U��Ӫ+JVx'�ӫz�j��n��e,Ñ���Z���Mn����Y��dl1gk�C�W����\�y�7��.��b:Q�L��K����&��|���y"մL��1��y�cݴ9����������,;�GS}emn�4,u
�u�#bam�v�S�F���3y��4,��%i�p=�Qu;m!{.Y��z��a=��+a�P�
�o4�uis��;E�W1b�8�|�*ޡǺ��x<p9wc&D4ISv�!s�!�GDӆ�5X.�ȅt���{n��kS�iw�ea�Q2�qI��0�T9�ʾ�nL(�}��XN
��oV�+���J��@��tt1Py�伢L����ʲ�jf�u/�>�,v�shNŐE�z.�>�ygE[x�Q1�9e�5o�a=W�-�#��4�Ȼp��q���={h�k���wM�<gV8̫%����n�0A����I-��7�]ϙ�H��㗳r��q�|�:]Ů�������{���mR6VXC����\��(Tz��ý|�թ_m�F�;U��%�>$���X�>�3�V�ΔN�]�;z�n"Q����ghX�i�9�W#A%h��tXwvU�@_9ien����qn��n�/���w���J�s�X��mos܀��5RٍpJ��m���1�̨�̧Y*ʝ�iǻ�8s��o�e�&����2���u�������,��6���U���2�X��;��/�ξ�2�=�TR�@�q�Z�j)WK*��X�+m���"�Gψ�)au1����WuC[�ۭ�O�g��С����]�E-�>�`�F2��|�ۗ�v��V��Zu(qt�ۃLR��f6�]��O�u�6��ڴ�'ئ���j��=#ms�����ujEkn�`��q�H�JĶ�lq,R#Y1@\IP���UH�� ��*T�EEb����"�X�������L��()
+b"�U`��D@F
ը��X�,t�բ��\q+�*��LLq���ʢ"0PE`�"�b��T�j�b�Ř֥eIX*�UUH���DdA�+j(�����Z*��5J���DH��0ETQb*�PPKJ�Ab�GT,TR ��-UD�"��VT�"�B ��F$��
�Y�`�1� *1V*�Z�V ʒ���,DU�iAV�*,�1U5j�TPģX"
�EaPPX����"#*" �YP�QTQb�eT���Y���)\j
��JV����tCw��cz�J�T����L 6�MZZ��r����irf�7*gs��^���y�6����?���%f8��L�����JڜLXJ5�{җ�<t?�m�/��l19I�o��_/1p+�����+$��5���P[r=��:�NMu� ܧ���ͼ'5��Z�EiL���5@�֢NC�w(̡����;�|^�I�5js���W���x�����<���f�P����`'��V7�q���T*��ϊR�1�ug����AISΛ{�c���n�m�G�zE4�����,w�՗�ei�f�5F�S��vj����K@�fV����N*r��Bh��^!�m-�q�'���=V
9�}8�oyYc ����dAMͽo�b�rx��	�6�lh���VN�Mq�w��۔�4�Gj�1ԭf��lsmvŷ_|���Y���szlȊ4(���j�t%��]"�E�=�+2�Z�bS��Y�G"�ױ6���"��[��#ܺ�f㮹�����r�����'K	�H_bm^H�=�s�ީ��1Nm1]���u�ixfv�rWh���5��쑷x�Q�d*����T�:.5����e����Uf���+��W^{�p�y�5�@��}��Q�nLP�]��!o��������-wa��4)�Kt����ѩ�S��A��4����}0UDOBW�3h�_.����kv^N�Gy�Ґ��4����nиn�Y	u����T�rx�V�����s���;�Y8q��o><�>-�͒��q/.")"n�6��M��Ke�k;�K[�^w�4qѶ����of�Sp^-{�~Zw�EQ���?�⸌2>�v�5>�+m��;���n�N�y��#D*;#�B}�eٙq�����Z��=�V�uq�����eԙ��.��$p�4dbNNq�b�;���g�Wp�涆�m�J����#޵�����+����cn�)8�Q�c����4�$���el���ח�y�e���^Tlj�D�Er]���b��y	�#:\s���^AmO[Z=��zr[j�+v��\E:=�f��k�Vk��ә?F�7S�="-L��R���'�u��kϥ��oTp�S�� u��<�+%I�7�_K�i�we�S�d&��%E�e��s��[z�>��.|�c�&/]L@	�����"㵸��[g��}����N�ħ���Z �ݫ��}��C���촶���ۍ4�(���w�r^vk�[>�ٴ���-+A�wR;VEY<`u��Y^�g)����.?S�iϗ77[��]֞���z+��P�c��Fo��=���g��K��k�/��\sz�K=i�P�tҍ\�V��k{���My���ʄ�HVuc�/��ƒ���,us��1>��.;ʓԙ;��l++�]���)@�I��J*y:B�nT�$�ݳN2�%&�b�?>].۾5	\�U���Z`F�t�@���p�;�ZInF�5�������.N���'6�3	���I���5���EE@��U<Nd��"55cHX|N$�K���q�&R���в��2^f�ﷵ�.��2)s܉�{�2�+>�sfIˇv��?`l ��b��I�qf�3(�@���E.ڽO� ����w��龔�rq]wCl���vυ8D�%���&��b�8z��;�.l:F��y⽶%�ܼ����y�:�7�JHP��U���cĵv8q����)w�\�˴���s��d�:A
��<gq���y웷	�ڬ��ʗBǹ5iɛ�3��\fɨ���k�|�/���T�����#g}��fz��:����V�ᜅT�L�;(���E.��҆�{U���l�Ԅ�Os0z����[�!�
����Om�J��fM�����X�Y�#�x�)�+���e,QQ�u��>��U�,[{:D����\��^f
�+Gޜc����.'�ЬW�]��;i�zzW���qכ?���|/|��R����s`<g>��Z��v�]��o��}���E'����y����~��I�5��qh�o~��3��U��u�|�˨�&%�Ť�Y��/��g����-}�ݑ=+�TR�|�Q����W(����v�����沎�];��}�����k9#+n'L@1�WQ����N`}Hr�KZ!�o�p�~�r�e���!���ސ��9+i>��3��;���R��.uٯ
�3��*�J��Q�s��T>��	.5�>5T���3M��mNγLr�C�4Y�]ː6ή��1��zc]o˔1�^�� #d�2��A�-jUr�V��j��dYfk�aJ��F)s
cc�Ƚ8޾�F#'��F�U���9�uz&����Qk1G+)��*ic�[x���ݓ}
RX6A6�nm5NM�L_D�$�͟���}h�a2iA{4iHkk��o��Nq�p��_��"a��J��s̔w`�&Ɲ{�8�ul]d���i�q�%�a���*�u����&a5��K�h�YPq	Er7����	q<��cn6��51�l��)ce�[��� 50���� *��K�|�R\�iP�\�Za�T.��w�W�;��]�o�����r�W���>c+
w�W.��Q<^S;��j�ޙ��a���%��Uߪ:�n2��y����g�9E�h�ͬ�kt���V��GϘu<������ߙ��|�JŴ���
.��̆%��p�_%yJ��wR�2��U��8�h.;G�>�>�V�@7%�O��S dLv}�]C�
�_{wҢ�GV7���++U�k0����JZ��݁���z��v�/u�_A�^�p�)۱�yR�4�u)���vk�9�Lj�\id��M�)�\|��7��lۥ8o'M�Z�N[k�G��u��eZ�<��?��� ���<�R����k�$~�>�0:^A�CiZ�������7t�ZoxF���IrZny=�dGS��z�u-ބ�vC=&�$�ɜ�ߥ�J{F��3����ѫ����c�Z�g90�\6e���Z���
���ƗK'1�`uH�P+�^q890�8����=���t)��#�՘�L�#(����6Wd(UQ=�"�����Z�Pi=B !e��7{�eTmY�y;��ԥ���w!���H8l�ӄ��}��W+p����\]7:Λ�Xtk��N{Q�n���mʸ�Knwf��H�6r�:�og�����G|��o���gINuǓh!Q� �B8�
;�
1!����Q���)���p�b�d���;�|�D�;jYo޴T�E��ߏ�VtY�.�r���V6�v��2��9�|��J{/{l��~p�EJ�7m��=��������>N>=d�f�g�Z��ݩc��b��ۭ,���Ck�;6+�80�(3n���&�K�u�ea���(vΪ�R�֖o���"��C���b�X����U���]�A�l�{ް�q�%Uh��+ưg�sn*r�~��fʕ���e��6'�T���ص��n��¢5k����YOo���3J��������bz�*w�&��9+�~]���}qˤ��c�W4+r��-�O�p�t^���<��'g?4����k��=�"�:�R��(�.��؋5�ĝp�\29����Ge��g��5p��UOZZ=� ��ض@sa=���I��^�n��[q�5�j������ON}	�\s�5`�RZP%m��}�ӵ�qu;d�o+U��{J5du'�y78��Mq��#������Tݩf�S��c;�q�$�Pc]�S_8o�D�e�y{�l[��	���e��]�qv�\�[�<v��FEsW
Y��OS;��b�i<*�c����nz�Ev��;��Qt���9'n��)@�Iʭ�Y�&`Q��x��]��nM��/$������u�xܭ6;���2�h-^(@�?���6�Feg�%X)��ṝ�e��d�Yr��ex�5��o_={QXǦb��bNzA������n^S�nK�R|����<�7=�\�Og���u=[�9��<��9v�k7�c�2�!4�) �ih3NeB����ܧ7���*��o5݄���I5(���m�J��1��F�0�5�'g[1��.5UIg3�E榖4����zec��ѻWҖ����z��!Ja��g4AufDR����it��R��.J���V�k�ws�W<��������M�]V�E.ڽO�[6Md�+&x���C^���(fVA��f�ce��k�3d�[�ԡtL��&M.@�S����kz���+�n|��Bj�UN�C�.N�;�F�L�:�����;�W�W�hi��;��CT�1=i���̜���I��8�N���9�����[�]�.(���Nx���}-������q�{{���]�N���������4f��_oS��z�˝و���'�����&��b��<�խ�m-���s�|qv�=�������w���'i��]�XP;I�y�4�ݕlV���Fe&A�.��!�'�lU���;7z�ͤ�cu HlN���"��C�P�yP�z�n
�#!ѽk;G@�KJ��^��1ڳ�3b�έ"ٸ�;��N�&��Sޝ�с�kuT��uwlD�=;z�7�&�Q�1��M]pߖ����fx_n���޺��p-�]&�>O�[���I9�l_g���P�n襓v�U��������i�o>���ɶK��������i[ڛ��姈�r�I9�)\F+�pKj�5��v��������y�7}So�I�5U��Mē��Y�9}i��Y�2{����̭��Me*�L�����U��k�z��U�Ig!gT�q�u�[M�7��^1�F_f��Γ���ګj�y0�L%�j;�Gt��}8�]��u�*���*-k"����3��'Ю1��ZRf��N��3f��r��)��IWȹ-wlJʂ�V�Xba���f�ӱ-�]�w��eV]�2�V�Z/�=�n�����V��+m+p����5���؛�;#lw\"A��D����o�S�)�;扫��r�̝�n���kY�b�R��B&�!S)]�V�ӧ(6����V��A��\�t�:N�ȼZ�^��7H�h6��9Ӛ���t�7��n)�dU�Q��R����s�r��.}��)ZF&;�iQ�ݹ�ٕ2��7�����?ks�F��[7�f��£VȨ�)��Xw��ZpY
�l�1�n���� s�z��׷�hy�S�OO��~v#՟8}�3������v���m����<tm{���z�E��h����w����&~l< �E��'�Z�z��'F��K5�3;��k���;KGmč<z�[yY�5iS�.�_lgjQ�?^�(�����<�ߩy��W�o�B���rƊ�n-u����u����w��r976�ܟs'W��g�7����^N�Q���pI���|�N�v���ZϣC;��{^>�Yp�Gn��9֕%,��#{ �|E�(�*/��Ӕ�.�>[���{��M}8{]��/S�OJ�P��%G;�"�3��:���t��)195
�	8��[�C�]ٮ6����~�J�zgґ��^\v���e�il��W�i`uZʋ,Б",��3��eok�,[�H�T\���p	�����炨����HX���l��3��I��׺�k/�Ր(6���p��֭���a�y��=N�P1'R�`,"��K��7t]�5)�o:�u�n˂3��;��j5��0���)at��M�y�R3Dt�euM}��09�j��c�W|�Y��(1�YO4�M������U#ٻu&c��9�;��!^���@_��k2]�K��q�B��o��rwk�ҡ�P�Ż�nP�
� q* V��)���җ}�Qf37���͙f)	�͡��\��n�ϾQbʥ-,���E7�!�1ft؎���vV�z3{$�pi�&QG�����{K�lX2\6&�ЄT�%�ꆠ�3ב�
�j���\�v�n�͡m�(ن5����),ѷ/l(pW֝fwGnQ"ҩHb���$�e ������.>[ێof1�$)5|�v�B��4�X��`-v�>���ri�L�l�B�򒻢��X��y�����vD���{0��nE����	�#�f�2�!�	�B�̥���Y�09N:���f�Mԣy�J�6��K��QO���ʕ���ѣ �����5�|�\���4���a���s�N]����q�,SE<�@����4�m33�}��+H��뗹�����r��,�Q!uӋ����S���h'{vN�/Z-����ֆ�� ��s=؍��gy����n�bP�km
F^�`Q�����U.��W�᧖Ø%�Ė��%�]�b�?)1:�܍�Z
S%)h}���5�m�Tz�˫"�2l���ߜ���]��;����\S�e�m>\�Z�8�[дU��e��L�!{y8�b�X;[�Lp%w��v�]
��,�w/mo5J�_f@A|�&���3R���u��{j<�J#r�E)���:� �c�u*��[W��!\��x���=��݂��nY���M킈pHW�#����ے��6����X5;yn����,�B�����Ck��d6�ݙ�`I\t(G,m��y��/�F����0U�����xev+���vBZ�`hl�T[�r��ouq�ո��E�R�����R�Q�3���0e-�a:��S3����\�j���2ص9�uewR�\y1{[\�Y@CS�1�����
j�lP��n��%bq��o���t�����m<��h��zv�m��JU��N��hj=9�pW^Ry��N��4�<����Xw$f�MTF�8Nj�w�Hӭ�@�*�nee4�0H;��K��ܩ�wd}(����e�;�>V�?����hz4�g��3��h��qumY�a�j��hk�R�ݷV)�V�Z��*�#�&3 �ݻ��(}�G�կ+ke�v|�Wt��V��Ոp��Y�q�1t�Wf����z�}�=T��DX�b�J�b�`��UQH� �� ���#l�-((�Pm/�""�dQb��* ��U&�ZJ�
��*QQX�ZŬ��� �����[`��"��Ab�KF ���QAh�Ř�Q�P*PT`��9ab"��1H��\�X*1E�EU������X)UH�*��3CU�J(�����EZ�H�c�(�QDLjAd-X��X���EX�#"���X� �DQQ��
0QT%J0��"���Q`�DX,(((�T�E��(�
��`����,PQD@PR�EDQ
E�Z� �QD\���EE���X��d�QD�,PF1�
��EEm�A@Tb�g�>�rc9�[�����h�|K���K
�}P��Z";��cf�����d3h�R����� ��;�N�+�t5|�Ο�«z�p|�����2j-��>�����Qnи�酓	u�!(�{��a֗���wk��wv�}g�6��w��gINuǓ_Z�#�o�0�V�2��~�w��^���g�#Q,��Jk�Ѷ��,0�͈�����iS�=|��<��=;2���^9��Ƨݟ�ұ���*�N�7ґ���e���f��&�`��gn Z��7M�>��'����A4�yGA+�*�*�O8Ĕ5��h-L�лn���|�_����G��%@B<�=�$��if4@pu��yk$���5��x��V���ø�����ńp��x��Q�w�N�ߋ�<�����=��;Wc��k�mg\�[��x�o�q���GdqNo�3i���p�gAf0Q�sYL���N;�q������9Giڳ�Vrvqsr��������U�N�{5��.����&��Z�����z�Nξ
�SA�YU�냹��?y��zŀ[�wb���;u+{��4��ז�%a��t�wH���Yz+�2�w��V�79�v��kC�b7ѹ�P4npvG�ڇ4��'{��zI9�+cu7_�z���=���q�v�c������C|�%�gU��lM��yV��TOrO�S=Mʭ*�'6��t�EsW
B��J���sF�l��f���������<f²� �.�P@��o��&*l*E�ʈ��~|�S��B7��ȓM-�����)�)|Q�̐},!bQU���O5\�X���{��Pj-SK!�<�Nt[��5�Y�wg��[Q�x0���#U%�ϥ��n ���*^t���`�G�m��ܳ;Y^֒ޓSS��%^_�0�\zQfE.{�(���K�VGCi�\_Ev �B�V5V?�gJoa[���a����>�k5w��h�4��ΚvߟM�|���ں�f�t�;�������.،�2�lg\�<`a{��<�	�W�'�\���ͦ��T��0M2�����<���i:���d㹔��q�JՅB�w5\9;����,[�5��\z�PEQ�)�[ýXQ1Fw)��
��հ��������Ww���zW:Yu�̓�{}@c����V[�.�\*���v������{���T6�a����� ���+^Ȩ�)��n<��,m@�j�7��[�0r.��wLT8��\{��B5�ANڢ���Ļ���c��ƫ��.9:�s�\4蜪E��h�8�>�X�.:|�JŶ���>�rӛ�<#+a�WN���X��xq{��֥��>��Tv��>���\|��zи5߭L_����=U"wi:�$�y�P�Z8�߫'��uq�v5eeiܼ��=+d_�_xu7P����o��'�暒�[$>ug�&2F�m�r��6��6_HƆwl�{��k[+���d[Z�K��:���9��dW7����k�T�v�	��qΌ\��
�o�Χ��t���.=6�[�	���-�0m;뽪�V�\R�o�۱��R���x���WRTN�7�K7���PH��`Q=}L�j�.y�x�fH�����|G��i]ʾV;�������-��U���u#I��*����
��b��Ȩ�72I�vع΀�B!�X�S�.-^�l�MN, ���w&k�S��\�e7&v�=����WX)�$����	��mŔ����h��疪�ad��ME�T��p��WQi��u̡��B�ZE2G���gIOQ��Z��;�rd%Y��������1�nK�8�s�'v
Έ)��fۛ,0v
��V���XW�vp⎾�\(���1x���W`����
�F�&4���j�*����W��.�Cv��cc�����,�����o
��b��pU˸j����l��a樒E࣫cyj�NSp��@�Ϋ���О��{~+��H��{M��cll������)�ʥ����F��bg��=���GSܩ�Ո�����8%�ɮ�͏}�Vr=�9Go��ɉ�X�[W��7҃�u�������e���UW�c�Q���r��{�z�[K�{P�B�!9�Y)WJ���@=g�o`ӱ�M�8W��aM��ҕ����K��\�!O��vPܳg��}��ӫ�/���ϺL�%Z	\�@�:�n��V�f�9�A��ק���b�+|��u��oP��Y2��a�YJδ&���f%�4Ż9�ر\��=��]N�%�tN�\�hnָ��#���wR��_U�f��V"�d��N�'�ϯ���Μ���L�ki�,�
�9�#
]��r�!�\#;Wk�� `s�&��L2�j@1,�9q�J�\��\�8�/�fU��F������1��J1<�>]X7v���E����n�Y�v�o�4���U�k��,�)����g]�/x�ei�2�I-}&�J��9�ryg��jݫoY0�<���2<�t�Dշì�14�v�y]�癥<ii�ݙJ5V��դO1���&��no08���VdR�=�q��)�����4ʫ��BnX��۝��s���[5i	g���{��:K�"�xB�/�`��˕v���U�&ߝtT>�[7����4�ѿb�_b��5��z���^wk���T���3���B&��9avز�#7T� f#{*�1rf�KnNG�c�7;��̘�p0�͘Ŕ���T����o'9�+i=N&����z�M8�߁����u�<���d�Eӕ��a���]�oMq�]�M(�m��{O ��kƾͳF)\�W��H-��\��=��"}�� �<��=�IH�ɟ�m�j���_ۊ2�c�Kp��������ĺ�V�A�]^n�8ͭ��)�Q��i��j���m��S;�I*�U�����OO\���۫�w���F���A<���f���0��/kbE�jl�r`q�9��w}G*2������Q�9;9���S��+%k$��Wk��e����S�����'���m������J	�'e=1��aI8l���g�硢w!��s�e��V�c��b��:����[8+3\j���О&�rxͅf�9l��P@��;7�̪�nV]�Y�sy1�횲��ex�Z���{s�MG[�쎕1�c%�QۑY׺Z��:�D�a��ꨉ(�3}�`�k'J�Ou�+&�٧Y+�P��x�k��BL��z�S�q0�DJD���d��Q6�&b��UJ�w��M���"˰��2Uމ�aK���u�wE���=t�Z�c�����P&����EXܰx&����l!>�e�kTǹ�C�h�&��4��ǜ����b��t����M�ѺdKZc��ΐ��JX��[��9�Q�-��=�>��zaی�Oz�j��As�ni*@���� �9K�gҎ�ILB�N���s#�%�%Fw�6�¸ǳV�zo�{nQnE.�yÌD�kW5�����.�h�-�~��>�3��q]�p�C��Z3N5�Q�M��m�G�'ٍ����A&�Rv�p��wL�(s�l��?���d["�JiS膨L��yN�݇Pr�ޒ����Yhfˎ3;wm�N�v�ބ�5@�6�B*ٓT�G���-~Sy�a2�Z��W��	�!X��$ek���yWJP�l�<�ʞ.~�9�~�o���<���V���V�WWXo\�;
�����H����v4���:�?N����ĭ����lG�k];`���Ʊm��"�s���8�S��)�z�nŮ�OWc=' ���"V]���ye�,8�����&�z��ڼ�V�<n`��}�+��#�Y���.v.G\��9t�ִ6�XŹB��@�A����^iVv	��Wvj�k'ۇ���2�U�8z���o@�3�� '/tT4yC;�W\s+��=�7)Z q}�*�v��L��+�}���ہ<4Q�V�K[�"⛯�,���x��v��#�C|d��������%I]�ۙ�P�)���=�zvy�Nǌ� Ԟ:߀�Wup����W�O��B�u��;aE+&d���RV@�u/MF����0&8Y9��2Q��'����M�K��ӆ����6�[#������;����e��~K��{!�M��a�Io8�{�Y�����7�f����}��H�Z.*�q��x�-%ML泫��^��B��	���7p�����z�Ho����c�_N|�*�}��B���`��#��������?�����N{!?ds�+�B�m�Uz�į{n ��j~���D�9���ι��z�1��<{m�F�����s�[͡ӿ?U������LY�w��x�-)
je˩�lZ��<��g+tB1�4/�>�V��a<��ϏU$vǞ�Gx��e�#�Ǿ�&�N/vd�w�\,M�E7*���P�/�ݸy���8�,�����vR~U�Wcϳ{�_4&aaK��-opH0mt4(Q�6�6�N}@f$�uE[�8NL��=zT��i��xs�%J���y�Y �q�戳�U��q]�CI�p*�}�E��ͨs�v�q0p��V=���!qB��J��wY���sH8�}g1��A�'�c���w��اm{2�#�����#"<�og�!�T�p�z���+���"���{�j�{=���*� e����zf�]��Ȅ� 'C��_7�8d!<6n)џV�Э�����F�d�r���Z#i�����}Yʜ��E�o�P�/�|F���^��D�^�Ho����%�%��^��P�o>��*�����j��8�ɗ�}w%:�S�~ �;2L�j�_G�=�_�ؽ������k�Kўk��4HȠ�U����mW1���2"����:/��7ڷ�T�}r�eI�ׄ?{o�By�zLx���A��|7T�N���ҝC�zU���! M:��X���^-z���_����XR���<5u��.�c>;u^@$����SW�Q��Y74^���l�g�$�?x�{X��7�6;��o����*�=�D�bH�]UR�>���W�޳���|"m~�͉W�lV�lD�M�	��Q~Ǒ��zs*E��~멭�\�#k|�<p_���o)��='@T|7y[�dF�����e�~�!V�P��ׯ}�fw��/1T���R�K�(��i�L=�Q���S5��5˂�J��_�'�t�8꒍�!5Dx��1�d{oz�6d�^�5L|6��a�m�]�\��{,�9IgW8.�q�vi����;�a_dU�^�L�Qn��o �]�
3��ׯ'%ߩP���:pG���2�V�����=��ҟ'^Aϫ��+�򊝉���4�����r<���Ĳ�[�26*�*��y騯��^�L{�p�W(��f�ҭ��	j����0�n���Gx�!���ϖ���fo��&׽t�ҷ�d�9����WP�i�_/\�t(������lx�ZCa�դd/?d�Cb9���_ �e_@�$���S��{+
̯yy�31��Z�����spSª�U9�{�1�wN�>�T�~��p������>������?��h�(Ex����y�x=5��פ_m��)w�==�Z��������X�r����O|#�q!7�.��##�z(y�Ȯ���|�h��S=���9�]o�N|�ֈ౺�=����q��=��r�3S�˅Ŭ��?h񪅃��닌�X��&u�X��z��C��V�E�j����ܓ�ؤ��v��G{����\ �VE�>�w����U��,G��N�!��'˗��{�~̎��c#|k��g�:o�Vt���(,���W�&E�S�1�"c�͏��Ҏ��;���Kg���	��W.=�|�r���(�;�(ml���9��f|��\)�;W��8�J�g^�K��q�ɂ������:���tc���F�G�0r��hq����E.�wT$���;ݙK�ޱ����@���+�L�zVX��V�7�r|�9| ܙ��1�=�r�XC��:[��� ��X���+�)p���#��07��b����{H.�N3�>E�b�P���݅�]���)q�xY����~GR��1)j�T��}[�K=���Aw}�q��\�G%�Ttb7�v�c/��:�]�k)l����J����kfԮȩ���v��{_(Q���Z���h1�m�n�N��
+��Du��ܑ�����j1���d][���+h������S��Kvb���Sᆬ]r�Y�psYDf��njxE�u���Hk�Щtϣ+3�h��^mpW�V��iu9p��Xl����R8T�\�H��Β.�X(Exc����� �
X�C���.x�_7j��Y�kj�6��WB�m!|���v�~P�|���G�H|���I]-�P4�ǵ:<j�c����"J��7��{�;�(
4p�����Z]����(,���J�hn�Jƥ��/�s�ֽ{٣��[��+��[����e���)�9]/���KJV��b��t����c��]�Zs���&: G7$��+�,W,����� �J����1�����mS�ɥ1��!ʰwV��恕}W�$ɓ)��	�Ǯ�h��C��凒N�O;���+li�( uXR�F.�AK��%�-��:�)�ˬ��t��Ű���=��KMn�[�����>K���U����i���])Rr����j��8e �}Z�Q���V�n�Vf`�K�O�we*E���S���Y���_C4�ko�r�}V1�0t�}7iV��S�`�sjeM�x�k7�;k��`5�����wU��%j�P�����j�>W�1��qG�L ͊���U����r�\s9r}�[`��dj[I���ݜh-�;��tW"�x�gb�.
�^�Zw�ſ����],��<s0�b���������|�n�`ed%�G?ؗ���xς�x>��:ҳk:��PES9�v���l�s�Ƈa�q%o�]'G�Vx���MD�� #��{�(NW�����r�t�����A��4���Y��Q��s]w;]�t��{rݽ���V��N�M��݁����HZ:���M�Swn�f�`|�C.`�ѫu{�,�A�hv펱]���r-�+&Fi��!��5�Fڄ���(<�t��V=׎*�Z��;����8:�JC���wEL�>�U���ٗ�r�-�ޢ-����e�J�����v�]��Q�3�'�*�a���\�*?G�,��[6P@�zi��8�*d�	��r���k���̗�o-U@P�#�J -J*

)Z�*�"�Ub"���YV"  �D
�$V�0X
5�A�`,Y+)��R�ŀ�+QAAUV(�-kl�%AU)*�"$EEQ�QH("�#iUAAb�+R�H*(��Q�Q����U��H�e��b�V
E@W)U�H��"����( Ƞ�b��� ��@TE��TX��$QV
������b��[bŭX�b�)�+Q-�,EYP� �X�Z����5����E�!U�(�E"�X*��(�m � (���D��,YAAE���IPPP�YYF"���T�H�X(�m�P1+U�,�"H,T*T��U��P��"�("�$���+Z�>���6�[�쵔Wr8̈́��Bl��u�n��_=�<,v[P���dYs�<��5���8��3tA��it.*֮Z;af��:�/�/�.��/nW��������/C���x���c����e��1���N^U���g�=�oD�]&)�ļOا�*��d{�Y���Ȋ��#�܈�;��{�zzQ���|���52}�����4zV깒`����ߟ��������T���z^���	�B��:�2�Ł�T#B��C۱�!\c��O��yt�Y�Wy��OY�~(���G���c�����y���ܳR�S�'��h����yL1�#4�g��4z>}呐��~2�����y�o���;�%��l�G��S�#l �cL�d��_�\{��c�ǘ��|1?������|B��2��|��J�g	��1�b�dGF,g&�z7Jw^S��&�
���_�
�=��NF�7~P���ʝ�T ̂���y���V���������oeg�N}B�8�2/ ۟_��O�!����r]���n=��瞽��v��X���sމ}bb��f�>#z��{6��\f׸s�F;q���V�=!�f������U~^�urN�*re�Ý�V
�:^Wq�{I&�j֓��8�t��M-u~gN��:�u�D�  �c��#�x�8�u����z2M=5��m�u��٨�ts�l>*�}�Ya�c,^��!�@�#���|�Ӡ����/���h���x���s�޾���_�47+n����o]�����A���|笚�'3��/9���� 6<9�3��X�N����h��Ix_�/�[�
�-�k�S�+}��^5���²�B��G����x�W K�� �M�o�뇡m!��c�Fx��s��c6���d�Z6��F}֮W�ת��׳�7�������j�~]a� h�Q�͇t�w�X�S������єX���J;2ԳN�^��-���D{o�4�xt��3�ޯ:J^��5��,�B�x�Ynf��7�0�������v��4}rLL�unX�o��������z)Z�8�e�-�R����}Wj۴h^�9�JG���/B��2�rf�v��QX����xlx�9'{�3��~�IU�{%�� ̷Y~��ڑ���{��ᓢ���7ļ���kbX��\��H`~�Ac�鮛�糧a�:ϤL��*�W�U��thb�2��O���@������߆���Q��}U����F�pM����8�U~��K	�-6����e�>;?-��z:p�S>�2�sb�v�j�o��{z��n����u7��fYݙ�R'�̩L5{�Iٕ��w}�^�d�i.�}mM�0��]BΉ� OHi��7�Tcn_�N�v�5�F���b�����5�I5�6&�����~����2�}~��N��.=~�J�������~�閮F�o�5����2�8����4]B�}��"����ds�I0�Θn��~���8��#z]��<F�����F�̯!�R&��#*��ee�9}�Do�о���I����@����>3~�mO�}�c_�s �u>�=�b_�(!�NO`����p�#z�D��9"�lH��������G���O�wt����nd{e��}AȪr�g���S
4��G��^��)/9�uZ<:��U��[��������#��yX�hx�#~q �?�:�G%��9�};�W�fӛ���a�s'{���:C�oܲ(o���u��u�]��ِY��y ����n���� ��S:��i�vW|��n=���o�Ƽ.�ܽ'�/�z�i���[�I�(= �C��Ֆ�6���~�˄��V�A�����]��̪���'l{�ߐ=��������4d��UqA�T*�\<�|${�72���y�0��(�M��P����뎦,�({"�:M�Xw&gp�� �d�缗��Q�1ΚD�p�3舚������/Tj��6�V�%�n�5�7%�Q�Z�[}/�`,�m���M����QM��%uA�e��[1[}����P-V�7:�xNb).���ߖG��g��߯��T�c��Wr�bd.�'Ցa̷j��U�n�D�3��`>�Y�R<���7ג�O�#ڇ���4$lw���^�g���R&[�6���n�-��۾���;��˛��ͯO��lJ���B~��o�����Gp��<�⛗4��U6�^w5����| y������lv�;�5�w�yb�Ϣ�g�N��փ�WW��շ/�Ub��Q��.�jdxI>>݊��WᐶC@��ז���f��@k���>ϡ��
g۬�L��^�D��ͼ�|�qz�{�]fC؏{ڦ}��7��1Hڦ�Ȫ�d^zj-����M��v[�8z=�3G�'���_�C�\ϊ�2���p��H��J�Y.NF��^��aG:B1za�=�݌�����Ǹo��~������}��c����]�UzQ뇁�F�+=4�zN��ݍY�N{���F�1W�W�
�ϲ!�=�����z�8�!�ݙؗ�4z�Ԑ�7+�c��pc��w��P�?E#�9?ү�XU�_�S�������B�O����wWp������:��ş�:js��ʵٻ����*WC�$�-1h*x"NX��3O(�����i��Rc�8��ٌ>�F̮�����w��V'c�j�����E%)������rB9�B��o�o������
��e^��`�G|~7���g����������4��9�������3�޿P����ױY������^��Z��U��Ϲ����3�}g�[u�.��:����X���x��gLf]��磓�>hC�{�<G���|��>�3��>"��F�88w���ՙ=�5ց���#�7�ߣ��o�m{����}w!?g�߾>V�1��$d{��ӰUmLѸ��4���c�{={��w3� �mRt���5�{.���`�ｵ��q��-��q���^�/���^��3�c�YS:����/�;iKc5��B^���W~c�ЂТ��67�+�<-��ܠҬ�qW�wlC��\@�*��7�мo<�W��jW�����L�WySn�ۈ��[Ի�]1�.�������*���"[� �uJ�h^��e��_sȕ~��Rsc<��O,�ş6*}�[8�8{mH~��Iy����:b��"|��2ش*Lo�5���.��Y봊�0%����w��^��2���y�o�����*T��ϵ�����ج�\�q���k�U�|T�j
��SA	�!�;)BZG�<\�(Z��Lq���e˽�����Q��*كhE���ۼ�{��!!�w;Z��ƅ��	>dUY�o7ؖ�\���">�r�<��n����wj�-U�7�!9�s���mFƄ�p�x<����yfxlz��=C��2ו�*W�3@�X�[��́��Q7eo�и_���^���R�Sqλ��|1��7~Q���|�~w]>:���b�Tޛ��Ѻ=��@r��4V\5������s��Y��:�=7vEi15Y�Vo�{�oyJ�H5��͗���5\o9~�<{]����x�{�S�K�nf|��>~���Uh�Y$�*�/d����9T�{��ɹ�٭�>�F��ޮ�z2#|n�V��x�A�2�rR3���W= ׼qL����|x�>Ȗ.#�N\�}7Ӌhp�s���6_�*��U�^���d-�4��;�޿`�
g�au�9�>��{��'����"��tA��'�c�-�R�����lƟ`󐪜�Dm_�Uʣ:��u��y'a?g�g����H�	��A3c�v�뜰�{��;�ǘ�8��[ �ߦj2���޻տuҗ��d��^���������G8̘���VQ���آ��Ǩ�;Ϭ1`P�
�.��]<�n��B��_���=;��6�%~�NP��ؔ 0�<OT�����X���P�.�*���t&��
����K ��ࠖ��m�C$�>Q�Ԫ�L�u`�&#u������e�w]ϔd�K�?�yr�Mm=�gG���Ñc���Ͱ�o�n�r�.i#�"`]\�iҴ��^s��4�;��d��R�y]K����s�m�ex=�ߩe��dȜ~7�+��D��/,�lO� �G���ɞ�����͏�ܰ�D�S=2�w�깡�/��\�<;�~Ź�#Щ0�|r�Ȭ���!��A���`s��B~���}@{WՇ�ki/���qġ��F����?ؑ�\7y[�ϵ��ح�,t3�~C�e�^�~�����;��k�b���w}���QP��,Qn��N�R�Ѓ�)���Z�Txe/Uo'�gV[�n���y���
��B}�Ӡ���Yp�׀��j��}μAؕN{!��c��G]hˍ�q����=�ף���udC
gޛ��+��(�����v�F7�h\p|=y�(\^,=��<������G�S��wH{Φ|S�̟N��bmz(!�T��|+%xomC����ͮ��a=o��y`�l��~Ow=;	���C��HdG�ّX͍}AȪr�f��{9�f�<�v��q����;�[+�׸6���Wg�<~~��ap�9�y�
>�V+���Co�=N�D3B���X����'\�I�\־�s_b��p�bo@�E�+�;�{Dsu���:1u#j���cC�fR!��$fQK.LK ��;��N�ր�Vr�ɝH�{���cP(v�9��Ѽ6��i�,mf.�%��_� K��̔���:��[�c���:����u����9k}�y��
ע���m_g�^���{�k����F�!H??{<������;�-�5���h{����!m���k�eh�߮����|�mWxg�n�y�A~ܔ�{�L�{�*���N������^���fJ�ڞ��Fd�B�d�\?Ֆ�@�<��̄�w�kr(Lel���tg/f6!�=�Y�8���ez}E{۪}=3JNmM���ȫ�3Qg�z���9���,{/����-_�yvdy�ߖG��=o�Ǎ6�_�ʧ�ꮰ��u3J��Fd��}>��,V��.u2Z�#ѽo��*q	�d{az���d8����?_�m��'�~�P0�i�Ͻ2lM��>��\�@U�m9��ؔ�Y�0���R��w�g��>r�j_�S�
�Bчl���åc�[������*�u���Q�3�*ܽT����P2\yߣ����w�����ޱ+��2:Xb��QP�\e�"�ٿp؀�iϓ��϶�~��NM�O%)V|�3�VociHJ=�3/}� d��gt���His�T�~׌����:�����ߢH�Ep�޽Bܷ��O�����3�z�9���b�&/T�����̟u7딄כ�!�����b���*�9��[�6��X�_\r���:�gV����F�6�F�8��[=w���n�*�b\H�?6'�A�����1O���w3�oί�eg��0M���)/ò��N��Y
�R�>9CO�Ǐe����֨\p|���݊�p_�`�~w3�m�x�t��^�0U��xH,:PQXԫ��K���9��!W��W �}��;�uʇ~y��yӢ|�w*u�^��v�)Wk=�&��^��k�{6�o�1�En[�PV�cӾv^�� 9�����huK���av�����x~��1Fz�0p~��=�#Ki���~���ow��$�\�ػ_�eovy�k��'�h��x��MMƲ/�!l�pȠ�yl]��{}p��l�M�NA��g���(�w�_�V��˘Y�{���|;���k݊L�jw Cz�΃U*|����o���VV���J��^�O�#n��6��;	�<F�׼��A#=o���(-ꙥ4M�캋�n ��=�����޹�U�>�
�zu�Q�-�l'�͛�~�F�{������,Yu���39>������{�ý
�h�D�]v�l��������{֧��1Ӿ2��㛤Q����yt*kf�	�h�>� 2�*g-�[���%��R
���C-N���!� ���m�c[{T1 -�/W-��d����Y|�Yĝe$�� �^��C;�0��c�P|�hs%�*�+p�|�sm�����8�x���������WU�#�ONBߘ�A؇�X52V]�ŀ�@dh^u��e_k�����{��go&B��9M61W�}�=h�ީ����Ý��1��-��[�T#`/ZѠ4=��֜��7�t`�$��^���59^v�ߡ��H{8$��{T�}�zr���������s��>�Ac�c��	Um,$;���?�(y��y��~�_L���5n�Ѡ��Q>�W�j��j����yM� �W�����*��"�9���߽U�z��O�ed{ۀ��w��{=�mq�\\�yP��Q�vEe�N���EJ�]�vy[�Ջ�.��Q�??d�G'����ݾY���T���}/+�v����z3�Aee�Y}��פ��:Ew,s�n�˹�E�o;����kK�/��W�{�GW�^�����&��ihȠ�쮸^�����޿|��d��eT�ژ���ol��_LϷ��\���u�C~�]){ۙ7/$d��7"����u�ё�7ڍV�]�iiZ�ۅ���RP����̮�_�??Qa^Ȟ�.[٭��h�T�|+�ރ*.*r�~�e][J�θ0��U{o�)m҅�aqv�}U���t檖�1|y����78/�ht�3��������@�\s:v:�Xnh�tVt8M�̃��+!ޱX�}t���++].퀻dMd���.˺Z.��h�Q	�,��w���.���k���c��+6��մ�w.]�T������t۾Ă�����=�����[bظXV���C���S>�\�R�aC�&�7�TOPɺ(b(9�ڴ�d�gG���k%6T���9ACI��JS�w8=�l9�uŪ��c'�^�y���lr��|�w�B�omՐ���b;������ |%j壮�J�x��E}�EM!]\!u��ns`v=��OWm��T)���]��"���>ᵷj�m�F'��k k��;�v��`adbT�0֪ɂ�,�i7�$�9���Kȳ��5u�yb�c2�mHr�y�qa����V0nke�����8nc9��|�b��wt&ε�}�pR�R�HޱCI(��b�sgӆ5��D��� ]g�CA�P��{s쫼���U�����R��w,
�Ҽ=%����	e��7k2�8�����:Z��`=�GNwk��ʊ.U�D󾮵P�r-Y{2���-q����_ %�f����Z�U��'Oxmގ=��R�7���q]8�wZ�P��� �=��a��~9ܳ�:�ꘝz����@N[�@���Ҍ��\y�X�(+�fdok9�.��I����J��NK*��}�������2�^���Θ��U����eu�r���k�(��G�U�� �W{+:�j�4T+���Q僇�'�����\�.@��󶅲�:�6P�v뫜cEo,�c��{���Χ&A��	�ǔ�WE���a�S
�� �k t��L�c��=]�@m���++�V�B�M&��kUݻ��DAC%�e96��
e��u����k	�S�g.so���r=G|��w-q��q�U(�r�K]n�jJ���z�ޞ�=�9�Ⴂ�V@��*ȕ+�ǝw���]9�xꍊlw:��Sr�|�Ô�{y�'��pkC���u�-��pL��*w[��e��+-l6�9͠���k0�Xm�t��ݶ,41� :�gi��B���;�Q9���Ω����M�-EWK+6�hA��Z<��;cYj�Μ�t1ǹ���jP���d8�'ۙ��k�1���tT�D;��~��_��*���.j�uj�諪q4雡S#*tN�%6�Mb1X�����fLг
���Z��tײ��F�uF�w�O�4��Y��8�iՕE��}ה��-��Z�֮�;�&�{WX�(k+q6`�	���3z�x�-YWE�X��O���ZO��z�~��ƙ�(��#(��H,��aV"�U�`����UQAB(,��PQ ,(
�ň�b�Ƞ�dX��(��iFAH�V* ����F����"1H,��H����AH��$STQaj��dEDa()VB�B,FF0�TX,`�
�EPX�b�0X*�V,EVT*�U�",X
-j,

KR�
�(���KB�PRʐ��"ȱA�,`�`���Qr�+�b�`���RJ��,���Rڢ-@�ER1X(��PQb��H��#dZ�QH+A�T��
k$�m���kJ�w��|>����x�m �;ۘ������v�OOob�Na		_�� ���T��< �f��,H��ʙp>��r�[_�O�k!�Ѵ�VG��u�9�<B��^��!��;��D/�+�bjo��oi�FX���U�Eە{W���w�:�Jt�߯$�'��u{ø(�D��<z��#�=���3Z2*yxJ5V)/Gz8�C)��9v�p8�R廕/K���¼�L���>�ر_v1w�������1�^A�+s�*����eۙ�P�)���C��9����ӹ:���g���fB����@yJ\���9	UN 3'�Wj-�@&�W�� ^�1UC7'�.*��גȖ.1{�b���lg�Ӕ|lN���=��6�H���2�UN�����`G"'�P�M�j{���Hȍ���g !cK"�)��,w�l���<��z�����.��Y����'��w^��l��w7א݉W�V�7��RW�þdC��C&��fNw�v��libgܭ�@�7���z��@W���t�R��*��B~�'kֳ�R�uq%��˞�Y˴G����B�镐�l���-�����o�E�]c�פ��U��c�uf� �}=[��	���\
/\�"�}2�ojб�2.��:�o' �J�I�FN�=�X�P�h
Z��ڶi���WT��t�pb�|k #�gc���$�B﫨��%�﬊�$��A����yZ��� O�9�"ؾ���j�[(�6WN" ��*+��d="�qq�T��ϯD�D��=��W#x��/'κ(tϮ<T���Ґb��vV\3��!�Y��w7�/�ߜ��U/�\�z*�����ߧ>j�2=�s>Le��X�BT/E7*�����'clw���-�����]ލ�G+da�Wې�2��N��wL���"��v�z4f>���q��w�9������^�8=F��}��^����|j���M���o��`g��<<p�\/gP�S�
��OM��Ʌ����ǉ�1~\2R��r�<=-~�!��=Nd����� ڃ���X�@z���N��cN��z#�e�k�dP��*�9�W�΁����2��'��n4����Iywo�>i[@�WJ���/|�#7f��������}�\ǼDt�"<.z�������-q�Gg�׳&��������{o�r�b����R��B�.yR��2��5���W�n�.����{�sX�:,/|n��c��i���f�Ǎ�T���Um�����
�{�ܣ����fk�ݲ��}^�f���#6�>�y!���<���q�A�F����^�g������#�}�p�x���r�)����1�h��eo��*QӔ̽ģ��Tl;���t ��zV��
̂�2I���B�:�wvQӢ
Nw�Y5u$X�o+)��]�����~���vI���y0�B[D��sI]Ґ�	!��M�T�tp*�GP���s����}"g�_���u���C�1�X%�X�k��#=D(q����C=����]�Mr55�G��x�Ě�N@��yQP����_�/�`:^���/7�����'�˿s�
b`��79�`ϣ�Z�@�j=۱S���Q,�U�h�k�: �q��7�vS��em$�)]�d��w�<R��^w�2<�HY>�0]W�(���=��J����?IƧ�-�����C=�I��X��)hwy����ٟyU�/S��&+fe�&����^��엑�߇���'ócUjX�L�T'�������2�F|������F��z�A�7w�=�`y +әb��d���8� -xR��DVS�����6�¯��
���N}���{Ϊ�B�+qx;�1�����+��p}���h�)��P��f����+��z�������n��=7[�<��^��}�n��<�d���u����Ѕo���`������+A�)汜�g��B�{�F�q��Q�ng���;���^�'���s�}8�k�dPz<�"���o�{#�P.�G?w5jsW&3R���a@C���I!�/-���6�on+yõ_�Sz����R��j�"��o6��.G�b<����ǀL[v�tW�%� 5,p�3Z�K뤶�Z8��iswZ��t�X+�*!u�\Z�QW��m,tt�8����O���_\�-4��!s���֠ϝ�'֌������g3ք���.��B-��ޒ���o�(MqY���ξ��|MEP���o�5�o������}�l ��0�^~�L� �u[�����}��T�v0��f�'^����5_�'�+��?x"7�^����w��yJ�%����������߀T���eZ��W���!{ا�G�٠�(&�VF]G��"���4����@y�:�u�;�52VE߬L�����~�+�y���z��6�x�m}���R�;r��D����N����"[� �yv�D�R�^]d	���	~��w���p[�q��ؐ�ȧ�Ho��֤?�s��#޿��"|���S-��{���O���+�߶|9_�L�7aT?Ҹ�}^8�6#նd-oڦgݵ�ю�ҡ���#ӑ�ș��O��)��.��bj��7A���F��pr<n�1�o��m.��W��_rx�^�vWj2���#J�*<�ee�9��ļ�Os��;��d7�#q��ʆ�/a�W�*�\�l/�����P�d�9�uF)WW��]�J�I{�E
����d�m�
o2)��͔�3���� ��M��Pӡ�F�a�;s��
O���y:ݷ�42	��GC��^��!�͙f<T�d�.�jc��#\Q�ظ�bī'�򢜱?�t��й�ئ�{�I[�C�M~�]t���ۯ �m r�ᬍ���k�h\s��Wr�>6=D�Ǘ��u`Ђ/�Z�n��d��7/##��y�D/u��Б=�3KFEC5�k�����=����~���܉��⻙�^�33p������wL��>��~��M�G�M��P#@hoEu��|�&�6�)��端o�-�w*�<GWm���"y��Qf��\O&�z�o�`5ƯʜJ��̕+�������;�Z�1��=�ϋ�IG��=�H�^�$y{�E�.��!ǎ^�#UZ��Oh���d�S��j�=�Q�n�3�)��!}'�A�4�����۬�t�oz${�A]�U`@$�H=v�p=�\�[�jY�w/����`��Y^�T�|��y�sﹻ��=��2)�����]  hyYv�j.�4&�s�'-ﻪsY)wk��D:~�5;��}!��IU��5c>V�:�u3�'�Wo�=>~��5��6O�o4� ����?�l1�lo�3L��BvK�{=:��0�D�R���{�'NS�;�
�t�Esku
u�9]��I;��PyǨ�X冇�ޜ��=�����`mҮ�S��<`�-H����ژ�Y�v��^U�A"� L�x��=�G]5Q6�=�#`emZV�̻��{�r��E��D��]�em�{�9L�؅����^λkWy���~wx���_7����@B�1��@�cb|4�C���Q=�ڝ�Sj;�4+�j���΋�)Fw���H���e@S��w2ǐΐ�pݎV�3|�Eg���c�Z@Bx�{¶�yGW��vA(��/�����w���"/te�-���;ֈ=�~�,<����]m��{�J����Fe��u���쬸g>��m_X�==�y�X٨�M3@o��7�y�sǪ�d����z�ϕk��dG��H��?M� y�ˆs��	��I��U��8z��<J��h{�1����ҧa�צ��������l}�>��rPCs�'�'�ϵ������oA�	z)�W�߫��������Do[#>�?+���'�~�}wt�}�$\?nd{e��]��{�1[��+c�D��;�U�\9����������ƫ49�:W�=ޢ�"�X���	BR�	�-�;�z/�����Ez��DW[��ھ6�7�>�Sެ=Nd�Ƚ�עaaƧ ��ul��9u	������x{��Y�Ϣ�]�9H����-�x|%�����8�xw��p�3+RS�5�[�\,\+f��&��B,��#�4��2�U4���c�[�In�"���fil�}�z���~l�w�Җk��1�qw���]�[�S���.�;ʶ��O:�����A��qݮ��C�P��	��M��&�ڽ��e'�_�޵�'=�7�C�&ߞ);G�! h= �C��Ֆ���r}L��ӻ���y����k ��v�?g��_�=��Iȧ���c�3jV��T��A�T�y�f��0���x�f�3㝐�6�#�d?^W��-�l%��lʜ��ܠh1э������gؤ��l�ޙ��dΪϬ����26�#[͚c~y���H/uF���Qc{fg�&$嶧�Ή�����8��2���+>�e͇M�Fӟ1�Д���7�	�ׂ���^9�X��v������5S��Ǟ�{��w��r����C`�o�����~�� �4�� n�N��E�M�z��=>aN#�C�ϽۑSq��2�h����o����z^p�\I{z��_�X�}�Լ��l)ߣ֯<6=]jB�{���}�n1��p6���HiJ�{$u�2����m!�9�ZF}���X��u�p�׆)�^w��T��FfJ�=�&�{� �C�Ӧ�|�UB��ީ��²vN}�b}y�����2�FCx.;���g�k�̏\Ϸ��}���9�b�Ƕ��*nq�֠h⍫)��>L�J�SM�]��a�i��n�c�3��7r�R�����a���F��Ia<o���纕�����i�]L��$]��w1q}e���������s��
 ���9a]���0l
r�Ϣ��+#z�^F�xWrE�!ϯ��v=����D��w+n|vj���>�c+܇�3������=|ƺ�����=�f��u�E\v㙍Y���^��4��]_iǒ�����6}�G|��쫚�~�} �1��so�9�ޫ�~������{���e��d�z�9��|�Bv=���?��k=nכ�g�W��U��~���y���uGb։�ֽ���K�]+����=/=�����f�}�jR�ڞ�|E���v�F�d����IQaYjt�>�C+�X�:����Uβ6�Ҙ�o2�^��}^�f�1�����w.�6���⡱����W���/�o�^�iw����5~��o�=k��W��WX�,z�v���3�2��g��S�dv�p0�B�L�U9����C7�Kcz�g���>�|�8 ���������
|��ؐ��ʼ@~��Cl1~qN��52VE߬_�6����ڢ�����<{l/4�}3^���58��w�iv<lO[�{c�5k��lk�f��^sz�ڧ�^l�e�p欷VmgR��+lv�0=j��6�0aQ�YMo�k�T�x���.�6���1��4û�t����+vC���y�R�1�z�W1��=s��i��;\��bV!H�)�Y�_Wfy�)Wh�.�ln�C�֣�S�}n�#�����T�Ɋ�:0���X�M��\��p��x=G��F�@�E?ZCa��H~>ʓ>����B��iǫ;��"�����^���W6=�Z&}9�&��d&��Y��cնd-�~�3/7݂I�����Lǝ.<z�Szx���C�Ut�2*�_جM[�öC��>S��;W~��c�+�_OFMv[�s䏀'�+�� -m:`�hvEe�9����\*y���Aο�����)�3Lz*�T�΍��H�!ud��Vú��Ctǝx�b��9�mv����5��D�L󳏅]�^ӄw>�l�}��8W�=�1#iyUϽ���"n<�ih�7��ٷ�!�{ϢL����<{]-`��2+��3<V����S�������s�[=��7"��?%�o���3#s+���z3G��ǲ7��g�=�h���+��~�	{v�������K��$蠩���O�Y�<4[��B���86��f���L��C���퀴cН� �&���T:ۻ��v�5��pV)/E{�(�[B{�}N�AȻS����Uި�u)�7��;	�=#���5\k�^���ۃ���Vأܭ�q�5�:�_.�q��E��|/?tܞ]Z$���%}ɼ��w��"����M���Y��--ܛ}d�2ܝ�Kg��QWhL��㿚z�d�b�#�uf�v�vK}Q�q�1�7�\��ɵ�ٸ�\�<�¾s��㳗��R���!�1�#>W�{����@HdS��r���FQ�s�s�(��R�3:������ί�z3
�Or���V�3��W���߈ϩb��~8<!ltU '�*���]< N̬b�ub���OpC���b�����Ν�<f�}�������®��vS�p�>Y�LU?f!1C4���3�EO�y�e�{u�I��!����Gu�'�=s;5�g�Κ�y�'�>�F�`g�z4��NW�&[���\��)��@B�Y�S�$6� X��WN}��W.����=J�xQ�Tϡ+�>�-��/���|y؞�(��4�.3�dR�,�D�O0g{���n#H��k��ߞ�xf��?��v�Б-�1QP�\e�*-���߇�p�A���ځ�X�����vW��Q���a���V��V{ݐ.ߨ 2�C��3�� �W�'����>P�fB��bL���-I�=�j��?U�c��k|���=w�'_����� �+.��2��b5Cw�79%�g�>�C���OKO&�8�v�y�ϖí̟K(O/E/>�o�՟R`S��ݠ2�Ζ9l];(t&�`�+���Wg��×1�4t���Hp�0ZY��V@����]ű�MR�`��n�D��k�	yչ�
�z���3W|�i�K�Hޮu�)}��'5��͐Vջ��+��5/uq����	vZF��frZ�Dlِ��M;�'y�0�t��q�����[��q��9ԕae����Q���հ�����M*ʝ��Xޥf1J�lY4�?;u;��h'ؘ��������Q�ӯ	-��#�����<�=@o$�s{�M�&ل��	NH5�I-�Mn�˔1�}�4�n���e�N�]EZiX	��㗫�|7�;{���ۆe�uubU��J�B)��:�뭾,@�yn�K�2x4q�kR�K 'nr�ɝ}۵�[��T)[�e��5&rIr�	�+�6]e��d^��މvI��Z�$��{Xל�.H+�1�Dt\7Z�w�V�B���v�<���V��pեf:��jtt�����1�j}2��Ƃ��+y�v`��a�WT������@>�u�%���Fui|yr�St�ÖfŃ>��l���,c��I �e�'�&�;vr��fu'K�P��X+3�/�v;�[I�ʹ��H�J,X� 2	������i�_	O�[D<�2p��e-�k8���ղ!�`���ˀ�1�]�N�����6��b�n���X�\wn�S�S#�b��nJ�X��T5[�C��}/���8��2����qGl���m��\q �����[Uh.�0 MۖOV�a�c�Nk�,�
�¶���:�����7�v5��؃����j����'��.�E(I��%Yو>w�	돤�ma�5%��Yd�c΋�+T�5������E�r�hs��3�7/%�D��{�,�"���-�l޳#�{m:�Go�*\	t|��R�	c(�Y�i�wH�օDF٠/5�jZ��FֆzF~ۦ��۠
41�]��\F����s^�o9��^� �Ȩ�R��OH��OP��r]�|-K�5�f6�yz�r�L<�=�;s����yel��k\k-eꧏ�}��H���O^n�������$�Z�2���qNI}�6^��>ˏM��e�t�\��ge����V����R����s�e;2��W������^ev�iW#Bf�+PwJ�Txt��$��]u��L��S���c�5��a�\HA�;Mk��$�_z�.���&��;Dxuq�2`̓;���|b��%}p�����ẋI	S�L�>]��w�JP��M�����sNŐͣ�G�!u���$��^`N[���*��E1,���"��hK�X��	%ZY�P�V�K��ڛ%��;J51#��9q=F�.:&5b��t�nF�^��-1��c�~/�6�_ʳ���قwoiN�	v�J���9���O�D���K'QEs����Y�|�t%��=o����5�n�����r����v19U�nG���k��@}@EbDU`�`�,P�~h(�*(�� P���`*bJ�"$U����
E�@���%V
�U$U��Q
�Db�++AJʑA�VE������,TE���V
�
,b
X��(*��Ec2E RDeHT2�X(,,�c�FVH�`,�+l+ (� ��UAAU`��"��`��a+"
�XT*(
E����Ȣ���"�E�����,X�!YE )F(E ��T��dr�VD@U�VH��1E"�l�Z�*(v�']̥�[�`tze5r�%�������_K�!�V��#���Xv�wrc.�olk���Gu�(e]�4��$��Y-���dd�}��s��K�Pc�Ti��ݻ���]ߡ{��(��Ya;��J h�Uz_�ӝ��q��k#����=Nf�o�=��e����q��ZWv��h[���h��z|?}�CZg2<?	����:٬{�F�k=g�Vr��g�>�^nX|��p������g��j�#��|F}+�Ϲ�ZjWXY�|������ui��ZY��Ao�*ܫ�(�V�,�JG>mr�L�e���G���N}����ю̜~�R|���f�^ z����M����ܜxWY�q5>�U?��v+�݈9����u�:��g������ǔғ�SF�|J���~��OVl��c��N:3I�?m&G<�~��#�G���l%���������5�����9�U�Ϻy	��fK��隋o=#Ba���HC!'�z�m��"3{��Ud�z�'ϨY��mξ�a��&[D�]�_��Xh�s�;Y�*ެ3pSL���^DWU_B��(��>��&U�7�S�������f%��ꊆ���o���ܢ\0}��d���-~��@5^���cI���سv ��d�eO)�3�)��:J���p��}G�^S�,[�,�2����3�-;�-!0M=x�P٧q�E��}݂^l��oa�E��F�s�6��Q�'v�v�}w8K���,NG�l}���Aa[v��t657�˖�������V�0��t��B|�ݻq���Ȑ�슊���-l�c�'|���Z$�B����[�g���S�z����ԅ����o�`N:� �S@ޗ�36��
IZ����ʱ⦢��z��Kc�MC��?M��y^xlz�ɟ>�2��S�q�F��hg��ͩ]�9����T��d���6U^29�<E�/i�����x.�2����=P�U׷���K�����j�� W�,9]���������9�Uqʜ������c ��\O%��Ú�_�]G���F#��z�F~�|7�c�������<ck��s�d���+��
,�绎����k��ICF}�X�l\�}�Ͻ����G�}A��]p�6�C����lV��ϻB��U>�<�L�Ϡ�zf�^��'_���Y��݊js�|/�>��]�(=XM���|}��������\=
���vpg�j�{��B�f��~��>�������-OZ�8�6׺���>,8z,9W�2�ެ��,86� �~���^�G�����_�NH�ͽݚ��yi���vfb��L� �M��o�[����^���9�Z��3��G�ېYԻ_�c>��P���$>0e9]����*��[��VqU��㼬=J)OKl��m��ݽ��xi�:�\;|~��.P/�fT�i(�HK�>�̈́�T�+�NT�T�w�F��u�4�W����y��Y�ו+!h���w�lPX=�T�Ȥ�;"�>!F�O����+�;ixʿFG�����Ӱ�l88����T�SI=��X�fUw��2)�=��Xb���Jȿè�@ԉ��:��#�u͟<}~$5�7�>�=�R�}�ns��6H/�'V{=��Ab��KC�r��VA��żMhڹ����K��<��@>v#�D�ǉ
��~����֤=�f���=���{����0.p���"v�/�*���l[2��@��U��o��E:��C<��Y��3-�N8���k����h�Z��ϣ��� ��P��X�`�ސ�;��O�~���z���v�i�wC�[�'�P1���*��\��� G�P1U��rr>�X��p�_��J�=U.�r�dّ�m
�Ԑ�g�;�<6�a�� �0����@c����.��Η�mzM3%�00"�"�.>��H�xᒝX��add?;�i{j��_X�7S4�eGeu��'�CG邕:�n��О����-\.��ܙ7�j����=�q8�7��\�B��4�����ř�^ϬE�/�E����f���Xss�J�\V����
����/z�$�]p��4�l��ƞn�@:\�����|q^�oe�����O�8j�;��/6#}�d�ȳ~��+=�����Ɔ�|�J�~�ɩ?z^+�������ix�(.��y�E2FPpguB�������s2Wk���XCW�'�ǎ����w4z*�D���o}F39p�꾟t��#�*�;�]Nw6�!h��s;�w�;��/�ZB0��{=������Xg	8���!���/ݏ4ʮ�p����������ig�Y��S��߯$ޟIg׌��X�vh�����,;2��.���C)��9v�k(�9�ڮ~�Y潙V�*��紞Ck���=����fO��
������vǶ��Sőٱ�d�BϺ*����U9�[?2�ex�T�>5�Y[�#�2�>�}����zw�^yӱ�4�;��NS�R�Ut�����tE���@�D���>�ފ�3Qe[#Ba��<�B��G����M�R�6g�߳���O6y׏�·���/�\T^�'ʬ2�d_���v�g�����7��K"���C���9D�;1ս^��q4{�ϱ�N7w�bD�f�K�ъ�n :���ʟ���y�d�����=����s�1��~������F�	T�1��N=�xo����e鯭sc/0܊�Fa��6ܴ�!K۝�B��}ȏL
�`ȹV�#�҅L�yD�:�X���^U͋�AC*L.#�c{<�� ���eS���s��	3<�b�������>���v� �8@�疀�t|:g�h���n�ݽ��r���\c��э>���X����C^�Q��L����oo�A�����;�s�u;>�W��
���c��NI�w��n��C~���S��Cf|~����ϒ��+��o�)��W��5���s������и��z������zw���y�ϼ�]ϧ�p�7�����K�t{ı�>��R{ VJc#{�o_���#�!�b}���8(��#J�*	١�/P�V� ����މ]cL��<nR^�R���ʖޙ����>=Nf�q�t{i���{���u�M��ry�����=��M�g����<2"�J{+�������:��_A�������Tf�;h�g�e���Fk�@����2�dV}ϲ��[5��UNqF��r*}���1�kg����x^O��Ó%���r_W��d���;Rr�����N��g����6.���iv,��>��л,�}�\�oݙp�E;�#���������_����g��3jW��jc2���!�C�*�J�#)�Gv/���&�^)�&��{�[8��vgǹ�G��\+鼻z���Në��+Fm�[hX�e��ެ�z=j�媓e)Ů�����`_a���)�ME�5+Vf��]��tCo��{pu1[/E����;cQ��ѧ�r>�u�tШ3;e�{Ba뻅����b����l3�㾕;��'���wמ���+�7�ul<�S4�t��g��[y�F��d'��>������F&�]=ٙ7he�-��D7L��y���*�=��2ؿ������7�t�N|�k6%zt�ʼ7kggif��p�f�ϖ��;�ac�8<��a�NS���"����\̯��"xk�찲Ǘ�����fܽ�4��PS��h:�^{�b���bC@����ߥ�(@́s9���ݜ�^�#�{ָl���>~�B�G�^xly��!ǫ�Z�� M�� W���N�#�K�U���`�UL��9���o�t��5CO�fs�W��s>[��e&�{bCU���yͩb|�T���*���o�?<E���3*�[C~w5��t�~���N�5�ÙDzû�� c�"�Ґ�޾��]�W��
ʜ�*��w"�9�r�\*.�w�\�*��F��Q�FD?vdz��߇���8uz���ٵӬ7�]sG�#��M*n[�C�݋��5�.��#�.�.�]�·�_Pg4
���a�N�[tZ��|��ԝh��3]�)�k6t�Qa���b�V���e]V�go��\D;��ގ�N��7���r�k8hҘ{׀'{�L�ݧ\/5���F��Ҕm�L�V�w�M���^��37_>�O}�/���������G�PhvW\=Y;������T>懛}�u|3�L�Ϗc���ׯ�%�����d��b���|/�d��A�bh��q��nty��C{�pt\F�\�5Y����K�`���<C����fM�<Rd��4m۬z�C��ຆ+3ｴ���΃Y��fC������Ldy���~���^�Gs=�=4.�����(�q�{�{�4l �H�W�H9v�k���zW<�ᰯד���6�z����_��C4�����\v�0�:�i�S'�v�k뢽C#iKc{��^�}*���S��R����[�)�O��>���5z�FE=�G�~Ur���T�Y~�QQ���Nv��>�ؙ���ڽ� =����dʼ~�59/y��D�����]��$Ku���ܫ�'Ы�
[Ȱ��r�]�ڭ��q��`��~�*�=lT���m��:R}��=7�{T�q.ϩ�����r�n��B��$� L�;\�������t*�����6��ރГ�ig�G�u��aߚeP:�S�m��.�"�_G��;�Ƃ\���5Y�~��ӿ^�d�{1�����4+��74h�Ń���v]��B]�g`yH�ʋE.o�-�,oi���m-b��
�����,=F�wwB\�~�v`
�b��jt��ݿ�{̉��]�� �����M�xoH~�B��^������5�B�^�WД�/^�G�����Tʿ{pok��P���rs}b^§��w��^�o0��7-�]�7�Y�\=�8.7<����~w>U��}���c�-(y.�����Ϳ;�~�E���K�$�m{��z�H�A�>�� ��&�{cc�ܥO�W6Z�"k�)�Z3����A(�[��yL��������g���D"�-�ʂ�����ho�}s&���ɹ�٭�q��cޛ�ړ�׃�fzWצ��I�~a�=V�d��<�sg��bH5�/������R�X͝�B��[>�m�U����s�]p����3���u�8���IĶ�D{�E˟ߴ��:��g�0��f����B|�+";ݔFB�� �[���i�����ʦ?1�GS?���*~�|���t�}����x":0r	�^G�Wc<\<Oq�/+e7�[��Ic��#4廟o���ݯ,�r��2_H�)���{o�g��dv��� @��
��f��Ք��G,[3T��K�Do7R�Ty���e-.?�L��@�x�9�OH�:��cp
��z.��;��j9���L�0�s@�z9�j��p��e`!��]��w�����El�Çn����N5�PEwQ�v�4[fOi�Յ-�L�V@�ޤ�o�u�W���4��;慴y_��;R�"l��	������_�P�C��0g�K���<���ݠ6W���"P�~9s�l8��$��8'��q��3O� n�v�=�f��l�Wr�ϤKu3�-�xT�ݩ��@A�W)����97�޳t{�������ٜמΝ�W�<�2۬�^*����n�r�n���4���~�3#��
^����관��P!�F�pM�;�A %��**��X&�����h�3= ;6G[]�Ń�A��i�5�g���~���ԭz�~��L����`[��E�g՗����wC��s�V�V��z#�"!����d��=�s�[�}�˩�~�R"�gq�W#��5�+�X/՗r6��{7�h_�ׅ��7��9{01�u3���O���& �N����Ƕ=u��|��0�fu�~o߁��׍'��0z�ې�1>����wt�x6''�*�no�N��ˇ8�=����WX�Xa��J���sղ�m���<����tǭL�<��R�R6�]��z��a�l����2+�5���qE��p��%-��UV��̎k�4r��Xy-���v��)[���v��D��9�<�M{��ˢ e��0�"v��"���;	�`�հǒh��g#�**P��+*��:M�Fz�'�S�2=�⮿{��8�'pϩ~\2,~*�����𫵝Q���v�BFo�/�}'iJ��C羑��ä?V�gܲ+��l�pȠ�ym۝͎�EXu���^ԛ����K�>�w3�`�nJ�f��'#����t�~�Rz<l��4��t�z��l`��ӧQ��2�7��Ֆ�6����vfB{^=������Oö3��9KqON_{9h{}7]]
�z�[,��=SF�()J�G�vϲDm)W��?^WpG���l%[M���{��=�-N_�\����z��k�����3�?z~Z�K���Ǽ�GaA���|{��#��C�l0�\W��~5��șlI%w�~˛��49�h\���O�pb�̢��bkяئ߽m�~R���ީិp�¼���!���V-޷R���=޽z�x$==���w�k��<�M�^_��ǫ`ul���d	����vC�|��MD���KѻjЗ�C�-�= 4;��v���;�c!�ِv�3��W�@�$��BH��BH��	 BIHIO�BH�R@���HIO�BH��	 BI��$�	'���$�Ԅ�!$�	 BIHIO@����$��� � @����!$��$�	'�!$I?�	 BI���!$���e5�6�o�#U�!�?���}����k�x⍵Ag��$�f�3\�R E@(���    U?�J�  ��  �"�( @    �`&F F&&	�bi��� �T� L��ɦ 0��QU�      � �F�M'�d��CM�F��[� >Q(sEU�~ph#dڂ�UO؀��S��?ş��(~V������*3����#T�Y"2	h( b�����,�߳�˷�h���s�JV�i�1���y����eV�A	�����I
a�T����+�U*�l��8!&�0`
�rEY��F9E���C�%�+s�w"0]	�U��f�D�n*��\�T9xr�gcB(JF%X��Q0�Sx���ɲRx�u5U��%��E���1w&jT
��1V��LD�JUB���%�n3��#�+j�)X�sV4�Y	lJ�ʄ.g�`�S����,��R��7wy�.�\N8�
�j�Me�5��18��_f�_Py��f��S8`�
I�RA��  ������W��.?-��CʙF��ո�Wgś�����ה��ڻ���[��b�`8�$��Jв�\
�5V-nd���̓,=�9VN��6�l��4/?2j����%�5��E�0������9�,d�B���Z��g`ΌbEX����ܓB$�r�h)�OgE��Q~���t<[�n��9E7m���F�HT�+ pA�t�dd`6S��j[y�gwĦ��N*�w"��7{�ZJ��S?=�{��&�7l�����RZ�]ی�)��gP^��G3>��RW�(�[e�)ŚDW4�4�Z���� �c���LSls��(,�4���,&1"��Pe޵c�l�.,r�jDua�#�B]K�.�M��]�63w.ر"��D� �f�i:�p�5�݋t�[��:U���*q�X��I�WA�5�&��PR�	e�f2D���"�H�{ШUI�Ω�ZB,!�/�
ϱ�.��e�7V��s�tܵ�;S��֔��9�#"٩�]4ٮO����M���P�:dT��nu��s�؇�S��o֞��������{T�ѳ��%}�9��0�r#��Z,�1v.r%3N�75�r�g#�Z#r���ՌǑ!�F�h뀣lL;Ij�םXl�E[�ӽg�P���)����f�+�����-���n���k����"bJ,���D%��|9��}���D�g�u+.��<��Ul�0f4q�
��}�'8�\��|�lA���"��V�j|<|;��8K�~�vg�|:�Y+�a��[t+��o����>�-��%�&��B�n���[f'��~��q�7���M�u]xx#�$x  8�xa��?t������f�UI��=U�l�7���=���i+
�`�CcAL�Ƶ�Dr��[��sk���M�pn��E�i1ac�qD�٘Ҫ(@��Ò�'z��MEnv�c}{�tu��=��l�q]�քΫ�!�g*aʱ>�c��}P�+��H?Kuuv�Ÿ�lp�����1[�(�U��]�\薨���0k��ʉ��6�9o�f[�98a��vX��n�잼S՗�3v�v�ݛ�1F����jz_���B��&�}#~�?FR��+'T&� �c�1��ܺ)_g�F+��m{�Uw�Z�Ь�P�u>����,�D����m�}a둑���%}�l]]��=4A�~4��Ģ��L3q7�r�@4����s�v2Q�1�:�*2��^"�N�̊��E�W�G�0Ww��2Ľ�6���в���$MV}^�p��AZ�j͖�/��5��/��;�ylZ�f���b�:�hs]��yE ��<�f��p�.����Ф�/K��ʙ��CX:GMaHb��R�o|��u�V� /�LA
�/G8���L@��m�@o�F�LEmy���s��1���CJV�RA3��)!���qu�WH5a��9q*`%6͐���G;�*P�X2% s��e]�I�x�H�v�F��UU��Ħ ��j�$V�6.	1E6��]��y�Z4rlk1Y/y4=���}��"��Ye������и�%�0��毜����b]\X��j��[T�ts\��R��<�<�`�ɇJw���Hb��e�.R��g�Δ�s�y�v�X�k�$]:{�b�C*ݳU�/����m���Yi=&��dё�N�#&�mm���]��v�j��+U�61S��dU�
�Kl��Д$��j��u����ʑ�QQ>��7�2��u��̘�Ѭt�ъ�)�oI1lݴ�v*jx��wģ�Y.�Qͦ����k,�z�4+T�r�/���NEY�3un�۵�D�%�ˁm"̅Cp�a������f��Mb��b8i쩟������<�X��X�7Zrht�dS�P��3k�0�=�$f�ַ�f�'$51�5*`HWQM#ti1E�=�v��Q˜y�
�:��:���+ur�D��Ox�t��>�++=�a��g�"���K&����Q�ɢA>�g�a�Y6��۴�ߠ��5L����Q(
 ���s���PW[��i�>"HF�m�	�c\��m��{��{y3�HG)#�,�G��KI^
���  �(�Am�s� Ӥa�G�ӱ�n��{��ߤC���AG�(>s��>�R.�������YX�9�(Y�&�ǷO�d��x�ӥ֜�V]�sH]�Yi^��ǔdS��sWPSvX�wNLDÆً  ����?"jP��@��T~�0�i��Xb���xz�( t�!��@#'H��O��p��2*��iӇ��:EJ�Fr�a�I!�C9�TX���Q�R}E�^�櫺j��d�.��H�D���q��ϙr�L��d�;
�"��C���[��ae�)�>b"֫���nL�p��B�Ѱ!��Mՠ���iE�8�)&%��!	���jIj���^Y8���0k~�7`�Y�LMd�t�+���8�Ve))Fƙ�0���5�A�s:v]�eਭ���Ӵ����u-��a�6/-�u1��VT{����W�:/�&O�)>~,���>�DV�3Dj�m]�)�9qhV$|4��� S�*Ԝ(��ޚ>
�G=���T#���a�j�)Q8���0�W��7q������X}E�0�,:�5<��2�F�c1l�@�I�xL�mu�tH�G3L�U�SҐ[�Rr��싾�X�4�V�����K�?@��}�n��u�̧�!23g�#���Pqf6��"���S�2�����J�ĝ���h�9�����f=R��}�����b6/�݊d�WSS��6�&
ntֹ�6�U�ވ�d�y��c�����2͝(�W\f2��d������#.�ִ좪�0:�!ь<���Mw>�=�����f.Jj���N����͵�WZ Nu�92��o7_^�Zk�בK��� INm�~�����8T�B1UUz�IP�31a��Ⴏ��(舫��HI��R�ib�2������c���[XjCIB
*���Kded,ˍ�6������_uQ�]��Z���E_YM�(N�w���ϚlMsvj�R�ߢĩб���d���3(b�3jcM�fq
,�P٩w+��-~)����m����@�zDUP��U_�:�(�;M��[�:(����>)�r�붹��_��.��y�J�H��� �үOld���_q����H{�����h������up�oÑ�ˉ����W�1J� �DU�^k�V�,{��芽�}��ai$SK�
���e�����AȺn�;E]�Jt�N-��m}�����X7}p6	m�U����|�hy�5�y8��m��QV��hʯ��v;����S�}�ߎ4���
9��_3=�a%ӊ�����=�����#�r8�w�d��<��G��6�3ͻ�I�5�x���T .ʽ芾���{�wФ���2kP�s2.�\}��P@�}d���jԜ(�3� PnPndAy����Ю���i)
$=�!��P�(x�k�M2/r��(yeE]�wA�x�/$�DU��;@��I���DOC��?v�^&�>F� ��ǊT�o �j3�uBI��^���~�ڞ�Y�+���-�}�zO��g<��(�?_�3I�DU��\1��ڟǢzq�'��Tޛ^ ��>�SL��Z�o��
�ge9�!��@�9��_ǔ��g�ΦN������DU��:����GBJ�e�&d<r
ߣ���0�Gm��NY�@�%��� �EW�0_1�S��y�ܺ:����#�8$��:��8ova��D/�|*�na7���Ƞ��6������ܑN$�_�@