BZh91AY&SY̔�Q;�_�py����������  `�~��  ��*�*���3�             ��J��(����@ �i�|T��#o�}ﾚ���s��+ny��R=�{��JPy�>;�Cl4[Ϙ�[b�w1Cf��\=�p�қh��� ���q_��:�:�;�nt����݊���hm��Ġ�|;�U^�|�:5�hWCaj�e(�ݎ�� �|v���]���ho�;ѭ:zn�P�uRS� ^ ���k륩jv�kJ֢��{�G��M����N� */���i_m�kGw'MJ��{���^�Ǽ��˝�q���Z����ઞ�5���8 �}�=���ǽ⽴�d�y�ȭo ����kFy�r�N��-4���;��n쭘       	
�@( I��=&����Bd��Q�F	��� 	�d��~��)P0 44 ���JR!I�  &�   ���P0��2	��L@�� �$4djd24i3TzOS �Ldjz ��R�Cԏ�0	�4� �h��M���'��	��R��6R~������1�Q F����`$: @�z@@S� �b��'�
w�_�������������C����H~Q �@t(���d���*����?�Ȋ�'�p��	������I$�51 �"�bG��������������ɒUC?ɇ~�0���h��!:3��9�xb+ǻ������=��I�*�l5�ȗ��<g�q��g�g�g��$�#�%�{<����/%��=�5��N�<5q>��w;�ſow����������&��U�;v��Mp�:�f�U3r�n#��Ώ�9��nç�'k�ߔ��l��Γ���:3�a9_ViN�N��y��s�^�\^�S�ո�븻����y��q�D�NJN=^Y���vכԟZ7�,�$�%���6�c�MYĝq��wpW�v��fdF	�Ҕ<�}�A߳�$��%ޜ�u�Y���7q,Ý
�r;ږ{�G�I�p�'�	����)q>Ĺ����H�{���o]K��i[����9�p��ot�Ǝ"�-*��B��Ğ�x���K�.+����{�#7��<��O��N"�/�]����w�*��fF#۩w����8�x��֔��=N�'���0��.�UG���}���{��R<N/$��*�8�Ԟ�W��s��{-�l�ߓ�gz���N�>'�梱�W�w��Qи��3��0�Ԟ�w�����3O,)iǥ<<Gq�r'ȣ�Q���g"���z���m6�0p�"�Ǹ�r^�K�仸��3����i]�ݥv�܈{�*ёSOM�~N��}�;,��%5%u%���=�݉v��Z]���a�xn���4�Ի\�H�D���C_S�z�6i�R��.=�',)3W��!Ήj8M䓿w%���W�W�(oD��[̮'�I�̏q�K��8z�Zt������|��ԉ�J���"<�����x^�>��I�4��r�V�'�{���O���=n`�]�D�8cD�.'H�{��ό�|o�a��jR�+i�|���A�ĜG�$8{���/�᷹,�{���,Jk$��L�S�{q.��
�M�j=���q,ĕ�*OPOSʕ�=��_q]�}	�|~��▖�J��Waޅq>�O#�{�%�ej=���ϊh�/x�Mf>G)���»�.)x�<�K
�8i<GR;��O�Z��V##�v${Ǽn�o|��.�T��
�<0���<Z▚�,��}�u~��ޯm�.�Z�����{�F^+8��Na�>�+������d�<A�.-x�N��w�=Ǒ'��|Nj(���Gx������+�'0��;
���+��N�	�|N�Oa���iW���Y���s�\�����s���5�|ΰ[S�M�i����⻍�)"���Y�0�u,�K{�{�Wx�<�^���͔��<4�#�é�N
|��2�n/c;�ߞ��^��D��.g�+����9Ȯ�z%�ir<OrK�%��2�=�-��+��D��]���YL�i����Biv��+��x�������[�?�"�q�|X|g��#�f�w���\3�+��[��ܙ�3�I٦Wh���q_��8��q���C0��ἒ�Ep�b\;�.xUؒ����\���� ��<R�'�R���G����Z3��;Ğ�����A�$б�٩vx�9j^\W�8�G�ؐ��T�R�{�ږ	���I���G��R�q&���L$�EQ�$����m�za�;GC�q_�ua��gzs�Ko��'w�y%����Ļ��8fޓJt�b����I��VL:�S�� �c�����qZ2y/{��0йNq^��<:�>^�.Κ����'��qB#���$,*�:�:��)�Vg$��;��r+���wh�A�$���A��u�e}È�x��v;;L���gS��W���K;�p�$�����J�����*wbWh�u��M��/��C�E����G��$��*���:T;�{����;:�é�R�vBu���YW	ܕ���n�Tzw;O������hX�C����`�{	�Ƀ����@b��#�'O��X��DŇe�\:�tzj����T�G����Ҽ���}:o�Nu^q��)�'mo�5΂u��uW�7S�N��O�������Їi'>�I���'=���d(�1.�T�%�qC�È��B��W;���g�����Ԯ�\3����IA���Y���SΕ�|/|;� �IЇ����%C�E����+�(v%�¨�yҐ�	��c����}�\�/�AtI���w%}�xn�[�U�������>�}���hX�A�%���N��4F:�~�P�X<O�V�閬>��:���Y����U�U�Q�S	D����!7��D��d
����ҝ��v��c\�vuWw��_��K��'��h���P��h��|�Κ�G`��zJN���ǣ�=��qvt�O���G�v�c�4\��&�L��NY(�'e�����	a5���&zJ'I�2nʇ��;rC���3D:�ٮ���t�gx��Y��Xk5S�:�v��!i�Q?��e.'{�1�B����6}_����������ӿ���1Ij� ���b���0m���ф��������]�ˆ�?��_f(�?�B���z�Jh������n�=����:E��iַ^V�y�Lj�3����s��Q��Zޠ]��Г�7g�i�Tb�2��ԜŜ��^{��~�ŖVmך�#t���nd}���;Ķ��@��͹��*d[��~+�ĝ���XF�0����-7:�Q�2��ot4��q�������OM�<��?I���՞5��`Y����B���Ix�r��f�����l�0�ڃ\�m>�ˎ�����>�p�+�5�j{��][�{6��^|Jx:��:Nw.��a.��CZ��*cV�s��,o��t[1�[v�x�k7�q�����4�df�,��=��G4�z�R{۟f�Nksۧ7��s_���exuW4B.��ũ�(R*m�����x~���Sz�m���8�,[ڳ='���?���g�<������TKj��13r���r�N�Y>�0\fF]cO9G��2����3�cH�4�~�4]H�����}����+:$�_���L��w�l?�^��!�y�w����{�y�Q�#�}��䌙��\�6唦����<�G�C�|�0�Ą*<���.��2���G�nq�s�^����K�!���b֦�#3d��7���Ǜ��qǀ�T"#�%~y5�O�Z~+�B���/ĢO��/e+k�*�XW=�Ų�D��|m�É�~>�wu�P/f��zN�1�ٷ�:jF�^��z=���p�u���p��f�}Y��̋����'~ɘaV�N׾=7r���}>6ux���[sƗJ6B����.�M,΍����|�tKd�=��3�IzӒU�Rz�~�����\Qm&����=�����W�;���g����=�FY����O
��k�(7�s݅����L�ٞ�a-�W���p�����e&x-��Y��H6l r���5��������/�-J��ѧ^>ѯ�2[�i�J�Ί±?����Cs�y���,fl�2��n<��׼��K�3_{%�0Y�l�'��|0�;=Tfm�0��ю��M��$�~sf�'��h���p����?�Ŝ�����"p�;�H��=�������2�VG��O5���$��肑ㆱY�=��g��V �����ּ�g��=v���_w{}�ˈ�\Ӿ���YH╭���}sÙ�{�cX�x�X��Mm���}����������No���x{���,^F����'廄���P�Ibq��0�V�ұ5���{=���5ع����~��6ba���b;�$l���y�sI�����~���j8�d�I1g`N���	�������n��y���'�{ep�+y���{�������_��k��.3ʼc%	�]u��X9�埄�S���r�G
���>�)س��~b���ɿ��kw��APR��\�ϳ	���wͣf�6��fqz�H���o�{��0�^���l/g���=����ӻǎ��λsI�,��K.s~�a�fC��/l>�`�����8�~���XeB,&����x�q-�X�X�9���l����9�+Z_U������EO�Jd|�Vg&w{��0��k�c,��GL4�,C̼{�˦��+�k��#���ι)�1ˁ�V��{{NXa�=�Γ�&(c$�r�ۧrv�~�r�t���p������1���3D,�v���從�Lҡ�WUnO\A��g3j~�do��{�ݯuYR �4{���}������<A̾�Vs�3_+���<:�#�/	4n�r��v�}���Vw��{ѓ�u,r^�"{}���f�m*#Yܞn�j���I���U���s=�.{��� �iu���vZ"��V>�=�ҙӸ݄����x����Cͪ�@�L���6L�uB���=���ڇ������K|�Bl+�w��vi{r��S��l��l/ޚJƐ/���oG��33}�F!G.8{�D�����_=����&����a!(M>��l�c�g�e7N��p�֒�sJ�:L����i�W<�.4uO�3ߑ�����w_1���_6aˢG)BJ0��X�`�l��� �XGa_v��#˲��L�
�N�~�G2���CF϶��][�	�;F��1���,h������	���P����/����@��y�ҝ�f�4ަs�ꁶ	\�����{�2Ƃ�*z;��]�չ�*�ܾpbP�k&�}ݐ�n�{�Vݞ*	���L;��Baף n�10�'[k�}���➪��Τ��+�כ�o���x���n�P������g�Q���n(WIl��J��Q�2A� �wp2��sQ�*&��1�=��R�͊�����u>6����Y^���BegT�M�c�e,�Ӛ�o\�Y��E݂mA+0�~�"��I��9�0Ԯ|��z���?H"��<��[d�c*��*�쾿(��*닽=z��K�Y?o����6,�_���U��GM��e?M)�M�'��/�C�$?l���P�~�e���_�V_ڞ�q������N*�,5��4��z����q|H���K��/��J�%�p󀋽�5�7��*�K�fXGjˏ�C�+[�� ���Y,8�9W�B`�!h7$I�	���*�K���i�'��S)�bF��!�Q6�!A�0�k	T)�'��#+j
|n��9�v�zkʟ#_n�Q�\B��Z,Și���\ǻ��=�C�͖��ZjZ��������e~� ����&�l[H��^҆��>�z�H ����a5�R9[���H��ffw(D���r!��}��N�"2��\Jt.ź�V����>���g��� Xh�0��R��G�A
d6����2H�a���m���x7��<�	���2��SPlၺ�C:�H��f����J��EԈ�N���>�_.Fp��@{�xvϮ�@=�1CaD��l��I8ӑ4ҍ����U�Q���sD�~#W僚>0%�����$�i��QHd�H��L�a,t�ځ�ZşT+@�@�4$�$�n�U��bM���|Gٗ�<Q�O8%��� ���}{|a��г	�Um�B�6Zм��A���|���T�
��h���D�a���"s���O7�{]M������>��MR�����x-����oog�D(��`@
�2�6� D��t�� �,\���.���|�M�DW��sp@0��JR|�H�H����e����-����z]�k[�C/��o�Q�K
��@Y���0�J
Ǝ"���f�f�oǢ�����N�5{���*�oi�n��B�E(~�}/�v���f=v�b^䵅���\-b�!d n��\Ѧ�s��
��X��~ֿQ�YEk��Г��� �����w����'���������ϛ_Ny�ԩ5^O<������|�����h �e�l ,`� 6 X�w{�` � 0� �@ =    � p4 � ���{��@� X�w<�y*(��2�<"�*��  @ �  p4 0C��` 6]��0@�6 �`� , ��  �@  �u����N����{������sF�++9�  �   � J  :P A �� ����� � 8  � �@P H    �k��{އJ  :P\�˩�Uy>&�3�@�4 � :@       �@����  �  t� �  p4 ��� �   � ��{���  y�W�y$����� ` �@ 
  �P H ou�� �   �  @    Ҁ �=�@ p w��{��8�Э�<��ԒO*��n��J�<�׻ �X�` 6 X���� 8������h � 8 Р �  �A ,`� � �����ޅ�z �7R��Q���c��Q BI$�����o��������?�S��?��T����6l��m�i��vm����o]�i[6lٶ�������=|��ۦ�v���m�ͽz��Jٳ�f�V�i���m�n�6z�o�c�m7Bd'!	�K���!.rd%�\�m�ح�6l��<x��޼z�m6�lVͻV͛m]��m�ېM���������a�hqVY��6��V����b�
5ȇ�&9�S�ao�L�B����'��fK�2D�J���2~h7���h��p�*lB�(���E&QC>�%���6qu�_K�|�x�c�B$�b�%���n����c�ۦ�m��Cl�8�ZE2JMk�me�c6k�~͊x�DGk��G!e��A�zrҡ-��R���Qfk7hf�If��(�[f��F!��]��}+�RQ����n�`���@��3%�o0�26d��j�I��@���8Z��M�n��Ŏ���ef�A�:�6���&\�!4_��H�X"aC01��Eտ&
e����>����
TP$�V_;R��Ջ���#gྔ�ٚh �y���5�m�] ,6�b<�e�:��[�e�K5���K�%�{���g��$q/ ? b)�6Zr:)-�����~���:{��^ A����{9�q���J�
�EWm�����i��$�Wm��ئ��I<��V���kO�'���*�����7���#8�qU\g-ċ���*>~�7�Ncx��.�/1�m�.m���(�;Zղ�7ơF����D)'�b"�!��L"j�'ji����Ѥ}�m�30�G�=��+@�ɗ���Qh�|�5f�H�l�[�UU	RU�~��~�������O�:3D�ݗ���i#ǉ��s��l  ]ʪ��gY$�M1���Q7Sy�>�n���.fBRX<�ժ��q��ѩ7w��Gl0�Ex �(~[:g@�=��2\�0�x�`�	�����<�N��䢪QEz�-)6i�R�m���r�ѥS����v�.LꜮ���FUѮj����Xn�j���q�X]�SX�My=N�;<a�<UW�bۧo�s2M�Hd�L����ui7�|# �;�ѝ��eH��6oJ�x�t��SڒS��u&0J�vJ%��IGh�`�_5QQ�:k��v�ˬ��n	�&\ntwc�--�e6tNDI\u'1Q$���AA���!h�<��f�,�WR��cV��ܽW���/������1U,�bT�R'm4���'i�i�@�r�����V��J�;�Hp
��jF��5Ԏ^Q!"�̊�ߞO�j-�U�P��1ڈ�6YCG?�}>��W��f�kM}gЅ2 ����~Q�#;](#u������M�������L���w�[纜i�����{Gq+f�Z�;�R���%��=>���+M��h�C���wGƪcY�Q`~�/d�=G ����[��A�UT���ώ��ar��A��^Wi���vK�Ȭ��2�v������S�J�V�!�4x���|��m�U���V6��q$����x�LL�葘�T�%&ܡ���p;qKv�S�%�J�MѢ�Zd�R������`�C՛�i9�rBC.�YL�LG��B��E���-&��z�(00��B����Qg�I!�1l������`bB��5��f���USUAzx�m0�;L�,�Pq	���*:M�6QM�;�����cev�M4�M�Ϻֶ�7���"t+���� �M��G�F��y>M2J���U��n����2
�Yiy��i�QIޘvl�dӓI3	^�L��|m8��a4e6m)=��kY���T_|x��,�;鑉��ETb�M��>U|�-���Z����).�m�0��l����L�)'���σv�VUD��td�ae��P�:,�[�o7�M&h��+U�����O�x��f��H�xM=��y+@e{��HL��J8��4�-������C��9Vx}���$F�]��앟&S�)pl���IǢm<�i��n�	aa�	Q|	Å�Ye�f�V�.�K���%�Ӝ�㦾!��A�N���cA��ZO%c\ۃt�@wI���@L�}\�����������gI��g��R��D�=݋N�ѕizvɗ\�$%x��<���~���A�qQ?�D?�O����D�D����:x�BW���6D|>��=��p�X�|(��>�	��t�$
>�%�������^׋8��W����^+�z�t�6�-]��U���`�Þ�O'���,������_����I'c�,��t�<������:>:OW$���6>��=!����Q�'��ͬ����~�p�6>��Gx�A�>|��	������O��|7(�e�=�٢�~��"���OFr���Ӟ��g.b���;><q���0�\{P�xLJw�O����^
�,�؇D!?j��0��>S�ɘr�-�8>�x�2�;Gt�D������U�]\����y��{/s�]����55��'ǳG�>�����~�캙��D��>׿~޵�k��ޒx��ڹ�wlWZ��*��f]�]kO������bӪ%*��33��)Uo���ŧTO*FFjOg��{T�Qq��i��-{V�Z�h�T��I�ú0a���Bi,12��� ���dx�zq�o�܀_O'���8b�dj��$t�ѐ��o�̳�,K4�/�HX�����QJq��1= �fI2����ı�Z�(���K0L``L�Pj&�H�I��A���}ϼ@�)>hR��HN䔧g�iWV�Wi��i�_=��n���a8DQER�T4J#�9j�Ѷ'X�+@m"��S���-�P�9��K���r�Q�#di줠�S���M$S�!]!	%��)�D���yI��L���,�t�e$���܍��n���;b9�ʩ-�@N}	$��%��i�v�I93М`Ri#�iBo�	
�@L,ENi�Yc"�GƘi�][�_�,��?uu�Y*~�Ѩ���]�$VH�?,��h��!�AE���%�K��3�75�JA��6&�=���z饬m
�$�a~�����K}҆J�T}����(���#�r+�Iw"F&T����.���5R����VQ�(���a"�VF����^��e�f+'Cʛ��ZV���"؍��B�����e�z�TRO��a#����j�q�D� ������Le�e�X�TKC��.�@8�+�� ��M��5���X��h�-�>�X0NE0�i� 2k5[���X�8ے�DET�R��Q(��Th�����Dn!���ѹ���w�<<a��t�����M4ѣ�;�wY:7��EE��%'�Ȗ�\n�Rܱ+>b�M�3Q�X�0?%+L̻���I�E6GQ)�Y�`.-	Fkh2���u�AD�Ӫ�$P�u(n'4�$R���1U`�,�j�9�������oOL�yJ$v�-"e�5c�%%d��JOP��M�����Dr��G^�#"�M���JY8~,��,����k�A��n�mQE�T*��t�(h�U:��2)ai4���5)���S��N6���014�� pA0�	�]ܪ���n"��V��.ah�G(��M���2�Ym���FS|2�> 77$x�LGN
 ��%��B�R�$8Yi�T�w��@6�=h��IM:L��U�S,<�;����x;��NΧ����0�C����,��1��C�t�I ,@���t&6�v��0�(���x2��/�u��UU��u8l
�g�ݬ,��~!ߘ/�]�i�a��˷,�2ڎ	,�Hk�J!���N|HIKk�F��Ω����J������xf�$+�sgѨ^So���e��H�h���.�'S�O:�)�����n+1�c�F�Ye�a�~>�����e�n#�r��h���vL�.���uJ%E!���$"�ϓhn�,h��-d\l�72�|�8|��Yx�U%1����yO<v����}[>M'R��f��.@���UUJ��M��XN�e1��Ł�tg	�L�d�&T��\ ��\��6k�Z��u�d�I�����JM�{GF$Y#Q�x�)ƃ�,����^�wt�XV�c�m�M4�O-��7p�Y4�"-�>���GkF��2I���)�@Z|rHz��(8��S���{Ǔ	���I��9�	%�e@���M&SF�yE�,���7`Y�I
+�Xd���0���^&WNY���h�t;�|��������FG�!I���[ǌ��!��(!e�Q����B������]���sP�"D�1$���4�m:��G5�)����֕�u>vk	�u(
>9(�|0�#�cm��S��F����L��:�L�����0�˜��N0���|���Zd�4c�´�᧏�c�Ŕ�S�UƊZ�'Z�vKaQ7*
qr�i��$�I OG�I	4���Q�p��f�]�\-�V��ط �$j˫�)��E?EQ�Oђ$�W(�e@>#_��I9�X%����I��ƒ���4d8�q��k0�	� �m��/[\����lͲ6t�8���n��F�ME����ׅ�� �,�O�Q�4�\c���0�q\x�c��xN���6>6x��O
�x���v�[Z�kW�U⫌�u�L�;c��^��=cj�<t�GI�������G�|(���ׄ������d���<�����t�:^�E��>�g���p�G�����=�ɳ���CLH>��'�lf���FM�	���`�,��$�W��x�c8�^/3���u�����oUk��"�-�����(�M���V�.:�CՑA��m���̫6�ǉ�����"��r&��CM����~�^����-�	������C�]hE~�"�J�
�%^G!��ۀ���l��O6�y?P��w�l�MYO3c��A �Θ�y�c�"7�]���D��2,�1C��[ʧ��V�s֖���G�by����������Y��kb'���Qe�MW�sXt�����#͡"V��w��hT`�78`�r~�њ�ˣ���#o��]mꖬ�?GgY�]��y�+����b����#ut��B�O!�3N�$ǆE���sY-��3�0�U1<���j�Tf��>J�A��C#��.�RE,������Pl�9
G �+��N��ߟ�n��$XQ����ن0�q�ПR�D�ADU�����/0���K�,##�K>�a������P�T2���	@�A�a��PU{vk����VO̴�0��H$�c*.\1g��@��s�o�����uD�U�ffc�Q)Uo���ŧTR��331�TV�Z�w�U[�ff1j��%H�Tԕ,��Y��!/8k�.U��@�K��{�km���m\�*��Q�H�1��Y��u�q4	ff,�w�=ɻ��j:&�x�1�"/�FsR6�2����ZvV_yO;2���>aT�����p�֟�p��΀����m&�c!�#A�]� e\�ÔƉ�e(¶i5�~�^��n�%��r��||?F�QEUB��>�Qr����&�Q�{_�'30�vҝ��攎4����$/�:�뭾�ԉ�M��F���,ztڰ�4�8i��Ɵ��|��3e�.K��_8�8;@x�|��Z��^N}>��v��sͽN�KP��o@m0{�ٷ��Qۜ�gKEʗ�!z>- ⎹ift0��Uj�[wm�"�i�������x�ɶ���m$	ߪ^�� s�UCN{�O1��Km-Ko�Y\�;��sȱ��+
�Lc��q�cMK(�%�-�tj�g�ig��
7Z����Ukی�d��.BKe�� 6?&Ϯ���=��s�Wr2
��E�yEF���j�|��y�g�ğGcѽ<H����j��#F�L�CE�]��#�]��t���I�/�a�q)zN��W����d	IGmQ�8px� Za8�<�e8p�a���p�òD�㌁`�'�:��a$�N�2X!�Ā�Y%�<B������^_�c��s��Q���J�~�ʜ��!�5�9�r7����_���b�0��*vn�K&��'N䓎�X��_��r�8�:����̰'�y%t��t(��G�0�v� J��E����L�[�F`U�4�̑*$m)�a��}�Y�B覝+
�i�O\c�D�L�҂�U}r�\w��������&o5��b�]�R!�Kn%Y��MVQj:�b��n�[.oqMh$\��w7��Є�lMF$��2�ݘdʧ��/��L�`�Ap��n�U�.a�P��$���Qu���,X̊��dȿ������F���e}a��H�HI�?������u��z�Wq��2�1+9�3��Q5�)��-!ꀋ��t���ܯ)GX��c/����k���~�+i��Q�͆W?��Ǖ��WV �����?\C�����ut:M��+�;�ǧM�
�i�N*��yɟI��0�e��F�:oG(+�kmjh	F��*L&|�|$*i�����2RXq�m-���<�9
`T��q�9K�i�q�����a�m��>�ZC�]��h%���X����Lx&& �$�!�q<��Z���j��j�wJ�����D��u<�V�}|���Յb��D��������Q�(��5D�wx�6%�M���-	@y�_���ۂ��$�DkD�3���Q�;L��TV���	�i�/,�220I*IU!��(v��IB�2r�Nf�[m�5����+&�J������!ħje�F��Q�j�����զ��8��Τ�7�-���NՅb��U������/���/6g��m�� �-2qƓڽՈ��pKe��.F��ߟ��N^% 怣l�M'M�M���&��t�[z�' �$�@�at��>��$2a�t��an�a>/	4���d��<|x�����t�g��&�#�÷�±Z~+N*�a���i�,ݑ?^&�Z��	���:x�4i�A�6!&l*A\i����A�B����?5":]�$�����10���U����j���ψN^n�^
&�ń&�l�,eB���I���M��6�Xf2�̴�2��-�k�zy#�:#�I�%�e)Zf� �m>H���ۧh�+ڒ3 v����i5��`l+)ԏ�X�+��
���ɔ��?nW7��eY"�?�lG�D7E�Z�	u|�oՌ{;t�+�
ӊ��j�JEi��aU*$�n�ꦁ/4� �'���:�MI%T�N:������6�ϱ�p2��Q2ZU���a1��h�2����wG^~��L�̦�p��)��d�W�n�e��J��{L���^9Vc3 �T��I��$N�șo<-��y�]+_j�G�����GGB#^x(�D|&�?G����G��c�p��D<'���Nxa�d�Byp�|)��^�'�4<N
'W��0z"t�����d��ñ�'��ׄ��xN����ؘz*>t	�Q�xk�xl�<j/�d����9_������4N�Gd�|p�;�I���'G�	���>&�����h�xx�6Y68l�>���lp�0SĲ��s��\/��3���x���4~G�������;?�u�e���s����b᫗;_���w{wq.W'���&��?<Óȸ���R纬v\/���8^� �N7��]�ŗo,G��~��7.sn�|�rOMgf�����-�33>'��S;J�w���-S;J�w���-S;J�w���-S;J�w|��-S9J�w|��-S9%H�Tԕ5*&�xD���$d��㕇���{㩀8���V����_�ӷlL9N:{�ӏ���W�l�B�5x(�%�oR�'���%�xt|S�� ��~N��M)�-�f4�~w�� �9��0�N,:B�O"Y���f�t=�]9���G�|���d&��δ���UOs7�&��5��cqQ}Z�Q����C�ZN�%���i�5���]���Q%k(��(����I�-t�m\ٹ$�S-܄���.'��^wN�Y�ZS�j±[t�<Y~0��2�ic_s��zϰV�sZ�77Bh�X��C���Ex�fRإD�q�m�`c&2b��kg��aK/�GѼK�h�O�N�$%�,���9v��q���}��A�8�|��~]��ʫ��������P�k	?��D��&�N��m�S#�$�&]�6��˖��KrrN�>>O��'���8Fk��YϪ�*�wXī���b�.&S��7����e�Rl!aa�� $ϋ!��o��&6�G&����6_�&e��O>L'��BB���a-�@<�2�������D�N�4�}��oS\i�DA�&4�!��'�zp���z�&����h��W���Xh���2.Q���耆	 �0K8Yt��������P�����$Iy�rt{�����U]˻%O y-2g	�8F�h�樫H��KlDbP��`y:�O��vL2��]Q+�*I?2��_O�n��F����/�.M�vF���L�'j�J��U�ͣi��e*���P�}�f*�h�H	�ag�B>�͑�2�V,�'�xz�Mm�)�Fw����~�.R��A���!y����,F��F����>M��9Oo��UL�J3$#���h���w�ٷɗltm28x�C���By׭�|�
-!o�!YL\%9��l Y�	�agB�Զ>}e�z^�{ַ�yZ�P�ĥ�LQ��i|�t4v�P��c2 ��#������V�f�H��K�����pb(*�h��6
������<�2Б>(G�٩Q�/�Q}�(��i>*�bo��-�IC�:��2:�G�z�#'�[��ꔔ��گ+TJ�!Y��ߝ6�cC�у�I�i�2�r����ި����E�BDHq\�V�F�����tt�XV+㦟��8pԀ���L���B�QFާ��tF@���]�M�SF^�L82fI!`m�i�ԎޖB*�V��lk�>h�Ѡ8�]����]��^�t�p�������%�'1M��� �-�SNZNV��F���O0�Cb^��0��*K�W��UJ�@�rZm�:t�p@$dM��I	��=r&�on8&�;��jKpR;ϋ?2�\&�+��[X{����O�:MQ�k��t'"��� ��:�n��-+Olv��Q����G��Z:;~V��!�D!��3RU�~cLn�s!k�d[jY"�6]�{	D��@.���p��.����s.؎2���-5�2EL`$�����'���at��Y��I!��	 Hۍ� mQ�N�$�2w Ri�[I���&�@`�S�I�29
p5ͧ�.Tn��	D��O�4(�N� �����~���*���B��?��������~=��O�=C�A���	�O`�Q8(�yO��اHO�~������GD<5�����z/VҾS�G��g��Q�vC���x�|O'�����j.���|p�:t�'����'G�	��m|M�&�������<	�|���������lp�0|6>��M8�^��q���^/��CD�U��\~Ð�P~1�^(۬Lp2U�m/-���]FFcr��%'��vc;Pw�WWj���w�/3�u�b{���H(���Ƃ��d�3Pyd%��v�ّj�6z�J�05n�D��c�Pf=�(~�4�g�͵�I�\iD�aJ&K����@�2%>���C�{H���|�8C#V�AF4fP������f
�\<�XN�q������ �	۬;,*��)����VtRV#"��ͮ�����^YU���Q�����de��8D���9�7#±�ް���o���dZ�1�Zŏe��S�=��oqr쥒iZBd�Ѧ���^S+ �;(O2�$���Wza�o�E�[�����iL�/�a,�T�!�nP0Q�	�*�h�9�B3�������b<�iP�����6���H��~������Z�͋�pKa,,��)��!=v��h�3k�>O�|��`O��b�wF������s{nh�lթ7Y��5��~-���$V�iA.��Y�Xgj��|���߳�k�P�;0��fgb�3���w��b�<���w��b�<���w��b�<���w|�b�9QUn�����y�N8�+�v�1�ro�a��\1��]������(3���m��vD�:��{,���<{�c,��Z�G��c�^�1�К�,�Xi��N�FCXJ1n�rb72�X�<y��~i0O�=N+�c��d�m�~z�m��u��~���z,}�:�@�ٟ;7 C�&�ӫ�RzӠn%��v����4��x�����賒z$��yQfH%��j�=�x��Y�v�S��Ǫ±\0����9���Yo�[d�(�ɛLi锃� SIi��Rn����i�v�-`�%��h�~.��K��х o����Q��}ձ�V��l��bR����RMd�i9�a���ܕwp���'��O�'`���d���9��X`!�A6К!���ͱq�y=�k;Ӆ�nBt��|x��u�U�T�THn�EhC�G�j�P����(�%p�Eu1���]$tջ[oc�J�:���ݺ|��aDmE|}C�����,�>ʴ�m2�nIn̎�����c�n�6�{�m�4x|�1]�⫶�}�d�l��'����),x�f�(>�:�����^\F�l�.�fL&дӴ�A�g:l)�{�&.�T���1ӫĿ��o�h(c7%�UQ4�'N8N!G#��<}$2H�2�ݘ4��'�L��E����'gG�cяU]�P��:� q~�/�UV�(2��B��Dح~2�"1�0�"�k�#���ԐX��k1neR=�bD��o�s�nhB.،���Kc�m͟rH��:ǲ�n�u��4a��b�W$�0�ii�)���O�Ͼ��Ѱ�@o�]�0��8�����FÎԾ�G	i�@�@ۀ��}�	R�ϠH�}4������˦����>��.�(ɜY�ڝ�֓�!Y����T��T�&��hP'L<|�K�PB	�$>4t�r��K �.��äç(WqI���y<����VY�>����`7IOL��'�'K�	w��~�?����O�fӊ8�d�a�`����)������!�>�e0��N|H���
��zG�C=x����Y�����b�Uc�VO�C���T& =�G����� drn���!��5nq�$!>+��;a������� �ե�V����QjL�[�&�W�_�Ro�s���;%_��$!
��$N����i�;z�0�x�S����˹R�t��B��O6�ω$#������3���l�M�Љ�c���v˻�}��Z*��ꡰ���]u8�6u7�Va�tU>$oRd�v7�K O�B8�Y�l�m�����~L���*�����N�'��-2��t�l�v�v�>���Jm0��d���QRRi0�T�SI�f��]�)��1��U�ʯ�;����DİM�)���	[zh�ç�Kk��Q-�Ǘ`ꦰ�CKZ��<�s����3Eu΀�[�BcM�J2��]n��}I%��fK��9��e�3G��F���~��!����v�%��F|�L5Au�o�ϡ's|.�yGh!�Dt��ђQ���s�Ơ�tv���Ci�2Ӆz��t��Qt|��`�y&ILK��&��'^>/�
�����3���42@��$6"|>p3'�մ�5x�i���Z⃩e�xZf�� �J�����q�D�j;M$
�6����i4��,�M
`쒲��m������֟����~E�������˖���O�x׮c&j�J�q4��a�{X�d�&0mw��牗WH|�%��z~�m�v��WLm��eV�����|">t5���G�x`�����6>'��xz>���M�����,�\Y��6���V֫j���qv�����z_���ߙ���4���<C�|>=�G��xO'�G���>!ӑ�<t��/�D��<r)���x|t�x�_��t|t�&�����`�l|Yx�����Y>!��l|n.&��Œ%W�U��qq�8�^/�w�~_{?�/���a4��~}�H��y�xQ^u��r�\Q͖y}����~�_�$h�5z��Y�~P�REU�?�E�_�,��z�P ����Ԇ���诊$��N
aV��>B�ѵ��4g�n���Zr!s�4�g^��⯙$��uҜ�hw�"T_|�z�C�<h[��5S��B {1\p�.�B愈Mjp~��G��y����Mg�w|�"�9QUn���Ūr�����1�T�EU���c�ʊ�ww��-U�Un��Ū߇8��*��W���uȲ�}�
*�i���aK�����&;��ˣ>�	+�J�~H%��-ȘK��Ē�E��맨�h�C�.
F�ja1�|��W��a������a<kޠ�[��1��[�@�>������6�b�Uc�W
_��z� s}��)i�d����r}O�=>�M5խ��yu�5����|w�F}�$��M�x�1���oI��!��у���Q�n�g褐"H��l+�)|]&,8���y:l/'��UT�y��	��Oe��~l�'H|"p���2vϳ�Ր<[��(X�C������r]�S/��{ܘ��B؈e��H���ޥ&��a���`GE��0�Xl����%�.�H��$Z$-�b\V�O�~�Q�����0�����lp���L0�9P>�G�~�E^{���Q��@��t��7�Hc���/���Ycx���Jeܺ#UA#:�͆�>N�G#�Ԋ|�i\Uc�W��n7'8(M��D�g������i2�L?l ��Xp�,8��l�h?�r������A���	�UUEUT,-�����Rd����7�[_Q��j���.����_FWG��JV��V=U|��l6����_�MCy���q�= ����$/Hl'���ԢbI�N:t}F<����-E	��Ի��vL,�d̙��$Hݝ�5�u�F���[~��I�M7������G�$d�tn����©�5�������SGjW��U��\}�{#.*�@7F�����E�E�,�!��u	Ju�9��˗(�((���`�Î9n!ΟQ���,�_Qa���ѳI���/�f�l�Ʉ������٪:��Xn'�'�,v��yo2�M�%�!Ĵ��-��� ~N	��/	˝��o��%?���/fU-R$���ڦ��i�Aԭ�$�h�0���Yr�hu�@��_�kOu���X? �I
�qF�f�N!$��<�U���jH��FX񷱓����GM��##�����g�P�O��4a~O&-9�H�O&���$�m4���|L�7v��o�I*L;%��!�e�(�Ƿ�f`�^[tt���N	�8}�6�&a����OoKz$<�q뎙N���I$�4a;�o*HIF#�����i8�r��&ZO�Gņ)��ZP_��Ϥ�}-�t�m�z�M�7��॥�i�Q�n��O4snB|u�!�t�Ԗr0�G��X�z��HpD�k�f�u3� JjQ���{MzB"wI�'��I�5Fz�_CT3~�#\��w+�� Th��'�':���l��%a:��q�-:p�!kG*{ͦ���G�����Uҕ�*�Љ���o���ҭ���}t�0U�~ ��r:�I!���@�`B���o�(��|���u��j��1�]K������i�?	��%g��O�Hy0=�y W��D�4�h>�$�-8�d�/E���a�?@�D���G��I!$��	ͦ�`��QQ><JD��x�G�#�DO���c�d��<H�'��xtx����xOG��6>	�A�h�C���x>��D�'�<*�zJG���Y1�z_��go�~~g�c�q+�|>=
'�
>$|J񨧇�����>'NE���<=\8_Ɖ��Ӗ�8C����|l��'G�Hp�;'��������c�U�x��8_W֙���>r;!�qp�0|6>���#�O
>��ў��\5�j�\�3T�[�g�p��L�?6�p�,�T"z�aT���v<�}7iAO3�E온B���.:_�z@�.M�s)�aa��M��O-i��!:mZ�az���n`Srs3�
���G�D~�
H���)#��uB���8�ǁ�6~�n�vDb ��A��c*��0�/Dȧn�b{^n>YVH�'�!)�/�0��H�1<��fU6ߛf#��Z�Q�D���O��Th����"*�̫D��� �'慫�k�A�m�se4���т�r�B�?H�Ϣ�	�$���T,�F�jT�c��e&�I�:l�){F�}x�P�"?;���$�#V�D�_nЗ������=�.Z�E�!p�J�ˠ�e-��e���[(�����_M�S��F�&B�I������C��z�o���5[b����1�U�*�����[ZU��{ŋU�֕o{��Z��>�����x��
�'�	�<"C�'��ռW֡��Un�RX�f�E5���1c����c������i!
�Q3�֥t6:�;s�и�5%40�o�$�R7X�⦏Z��a��x��,�T���FL��I��d��?�&SG�����@�C�����:�t��I�z`7�Y���{��$�`v&ҞO��!�o��uX��\,����ۄ,*:,x�A؉��/X��Q_�6�]W��H�y,��I&N�ل���1I���ϙX!Uڲ�&X����j�CF�9���Ji	��#�I����\&�:�Dӂ�{IăI����u{��U�+�v�C�'KG��]]�� �L;Gh���!z���^@����Ň�O�|@����Ϳ��.��E��L�V1.ىx��AUZ3l)��z�yÌ:�WE�h��,�Kk�!�dp�M����zY�Z�����b"BtM���Y�^ޯ>LL��˓2�,c�9��KAL\�;Д1����AIA5!B��ݤ�.���ۉi�p�蒡��MRZo^�i"YrC�f��_c$���׭v�I<m�m�w�GL�%}�r�U�c�=a���B�d,[m���9I���b�EH��0�%��F�JS_�$�i��M�J�4�!c3,Z�������*�5"���h�F$��V�,��ƽI+�O�˩	�g5&����$�}T�q6�`THRu�v��EJ���\՜Hd��Oxƀ�����[K+4oP�=wE�ɫ��������:h�)2n5���:N*��қc�0��'���i�#n�NWM�>�7kƷ$b]U�Gu�1��&��׌&o4��n]'�N���(o��m�1��e���dQW�ˢ'R�00Ӭs]�b�b�zN&��u,͝ZO;r�;��l:�
|!���6>���fv>A�x͵�j>:Q���>-�����c�UI<Ji8�����ڟ�"�˸��h��(�I��U����󧻋"y3�BL����Zm)���HC���Ur�J���g#�O�$;�4��3%�W��Y��'H�C"@��h��!�.~�{{޲�f�+L/:赶I��rI!���c������#�xH!K��i�����X�`�4:r"*0��ꮕһ����)���C�Y�0���_lֶ�I���]sl�Igh�i��z��f��Ǔ'���'K��B�@���>!x�r��q_�.�\�M� &�Dak-<O�1�L��g=�ﴐ��2?%L&ߘ��R�hXQ��1E���#�"|���$Qy9�Xh��U�BI���!.2呖 �"b�i]n�|~����AfïC��nI�z�#E�	��eu�'�&�<2��i�����~)��Mg�O��=����Mm�@�=�ބ��z���!'�=8uD�~�@��0�B�?z�fH�I,a"J�qV��U����ʯw�N�I.W�;��u�`�Rc骪�0y�e!��~0D�>�*�$�L�&�L��۸q���u��1�p���(�	���~�n5��[V�bdd{4��N�{I���F��'��@�t�zzz|l᷊ٶ�ci��6���co�|�M�͛;lٷ��6l�����N8��qx�m~x�Jٳ�fʹۦ�6۶ݶ��筶��<vӦ�m�g����;m�o[z��v�m6�lٳf���O�6��m�i��b�l��p8pC�p��ɶmPӷZ�n��Y7|G�_6!嚇%����w����^��)�l%7=R'�o�h����Ov�e�ä^�I�ێ`�w�l^�B��6�|�]{JCr	����u�G�����{�5%w7���rw~�^��kuy�������U�J���o�^�*����b�z������U�V�{��-W��[��o�^ȂxH���x�!�Du��h��[)�ˤ��誔h܄���Zm}0q���S���{)����ԍ�u��Y%�X���p�˫��Hy4Yi��W.��7d$-ц�a�I)�Z���}��Z"i>N&y_�����cJ�鍱�x�75 ��̓�V����h�4J5E��=�M�*ƾ��]6�/▚�Φ4�G�@b%ć�G���=E��"���2*����u�9D���U�&/J�HI��N'��O���B`���D�x�Zx��ke:}<�����g�q��UN���!��+�'�{�t�,���ql>|��I��<�a0��ml��6�4%����YkdDa��:f�P��4�n�i�'l>}��[�J�o]w8��G�=��%����)�FR�[�IG���o�䤴�G��H@���⌐��r���ii�}<�,�T���!L�"��]�P�`��6?6��F����6x�mU]��Cg�nFi��4x+�"�M�u����Q�̣&�Է�G-�̥u���'�ݦ_�)�{����݅Y$d�BE�n������z��[�}�X�팕e�ߧӳ�0�D�CD!�y�w�ӌ��d�7�s��,6ՒHZe6e2����^]�x���v��[�'�2�Y��Q��2�cl)!N��G��M��$�6�N&�g@����q�R`���Դ�₃ec���Ǭc�>��j������,�-x�(yEְ�M�l�g�Mˌ�@�p�Wh��ߑL9F7��l��	���ٲa�'������V�M�۾�<t�tS����Иc��6i9�$��1����

0DM��Cg�dk�լ���$
C�"����8��c��B�g�n���BR��6�j����$5LDϱ�Vy���a��Z��6�jfJI���'
32�YrĹR#P�ʔ��U�)+tJф�m�є��!���TQ�bH�G�!��ӧd���)i۳&��U�J��0S�0����N��z��^s����$8�K�N���'�����wE�#��y�ԁ�>��q)�|@��8B�yy5~�����8�y����c���IY�w����̘ČG(ѲQ�>�|����J��\+��J���uU�	��M6�}�G0�y����$Z��=D�WT~�5��~�|�E%�>�ݿJB�����5,z��׉f�La�>U&�x�!��]��E�0��&~ṙ'�HM&�I����p��xs�ܢ{���~���3���cV[��M�\�t��!aG���E����G�IM�N&�$�M��!��E���<���N���0�U�1EK����0�Lg��~���v���"d2ۅ��$�&������JL��Hʣ�u�m.N%nI�y=���:80��<z@�غ��ؒFrD�ӯ������]ѣ����᳆�6ڴm��t�m�m�>m�M�V͛6�[6����fϏ�+�5�XK�c;�2�fFnT$$�	J�m�v�n�x�珞������N�!2����'a;N�L��K��4��f͛Wn�v�Ǎ�Vݱ��b�lٳsk��m��v�����C��O��6M�$n�!�t��p�$����4u���Z��;i�KY�N̗�a!x+�����@�!D�bt%O�'��qҐ�81��kq0\u��NȳT�����b8;㛶�$y&<5���<͚3 p�H$��M���`<A� 8�[���׃9�>8F�5Ϯ'L��K��Z�b�-�ɤ>Z)�^��{NE-��6����f�Q�c���(���3.��?��F�G$zq2&�g�x9\6�U	���*�d�>Q].{1��Sׅ��X�*�4���%�PC.��L(�oV$���*	�Z~�q��ٕ�"F{�<���V�;h3|��g��U5,��.�%��1�.*	�O�phHℂm~���l27(���dHF{��1cE�� {Q0J����mBL��Ȉ1$�;1�0X����U$� ��I�G��-����&���(�L�#�~%�0,�e�v#��?r�7���f{-�ފ��{^��z���������Wջ��{KU꯫w{�����_V����-V�a�8��1�1�?�ۗ^]�5ĩq��v��
����`�v�]�z�����mY�k�
��]}lw���]4#-�ec�%5Y�R�/7�'�yL`)�2��4�i�� 0y�?A��	NK7M$Op�q�w��[�{��0���L�5<J%UQ*��M��kI~u�4�;�N9�`�
2����?���YgΗ��0cЙ�w�;o#���a��U�aE7�z:�fkt�����kT��17�/.í�R���+�;L��&��Ē������R6Gu��=�n�:v�՛�$%vZsi��I!f�S㤐�L7쩞�o�3'Q�v�ѕ=8�|������C�����^\�+W%���'��CG��A������]��޶$�)%:
��S��k9���˗�E�Đ��h������U��̒�ӏ�P����i8��>N8�*BMQ�7G�݈��Q�s�V� C�"h�HB�Đ��2�+�	7���}�5��hʲ��Y*��Yud���v���M�6�O$2��Kn�P���m�	��>��?9=!�~�tĐ὎Ӊ�����;�^�VF���c1ꪻclaៗ�F�ڣIG�in�k�r��gmy�`�H��&6�h�0C��[	�@EϓM�,��L-�lƒ��;�_�����3D]���ԅ߂�}H�H�.X�chh��$��&ZN����G<�0{[$�ޜ8�L�<��VD�	'�!P�5(,�u�]�0W'�y)5�=D��It���FA�n�ӎI(��72p��4��^9�L�(2a�>UWL|�1��MUSZ�V
kr�ܡ�c(���Uۣ���,��'�H�o��Pq�S���$�M+�]Y(�Uч(h�v̑#�H[���/++�!\{cY��M�u$�Ԗђ�ө�y��d����D��:M_w~ԗ��&6c|����w���h���V������@Y���Y��0��1}�7���]��	F�9���J��:�ӔI!Sn�ܿ/�M%�y۔�`���!��0DM��C�9;�n���Ӧ��z�9Ь���*F#Li��N�v�6�̄�����'.���/cc���l�D�W�F��ȣ	Q<��$)��q2!��S&�ߋ���2�=����>�M� @����!|{L�r.Ú�E�F�	Z�A)P!|��Ö"�Ō@]$��P��������rv�o��=.t1rU�x�!�AZL�a���U���z���
MvH�%��rm0�Lv&���'��UR��:�Ϟ|�/�L�޽�}Gi/g�f��#G�te^d�|ҹth����2���,DL!���x�7c��:U}r��p��I��i���HK#N�2�%D5��pn�]ߝu�h�&f��������Z�R���6�|�T	����I)�'~��M'���WTK�%�^x�O;:�5�J�ӣ���Ç6�[mZm��tm�޶��O����f͛z�_����V͞�Wk��\]���m��^8�\8vl�j�m�m�M�x�箞������N�m���m��6��Ͷ���ݶ��m�ٷjٳj��N�x��ݴ�M�[t��6m�x�M��k�������H�Ŧ�����c�"Ԃ�o��͢
���LO��X��u�5Xe��B[��-��_+F0V��8<p�3��Xi���ٜO��q��]�)uX[Ѕ����g����575��7貿����6�E���-%�����Ut�Q)/��q������r��۾�]��	���p���PϏ�S��~[v�5�����>ɦv�S[�e,ʽ�v�;s_׹���w;sⱿ{˻�»�>���w��wL}U�n�{Z��������]c�Wm��֫�t����u��df�Ԛ�DO�CǣFGଣU]���QDl����*�̔�n�} �Z_�*��Ų�_t8�sǼI!ÒC�I����6r<�т�G@ZQg	&���I����lDO�4B�����-��d�'��J8V�M���S7;����f��wK�F��Va�%Ub#���ͥ�)��d2�)6�z�I��G��$���T���7�	��UT�&N�D�W�O=�Iħ	��ϯ��]	Z%�4 @��D��<~٘I:C��[�m����%��mn���cL?7�!Mh� �K��ne_�$4<�k`��Sc���ԉ�c�پ�:��vS���>����"�����N"�=�;SA*��a3:Q�i1(��"D����0i-�O=L�(�V��n�����	$j�GM�+t}���=��Z��tl�y�;M<�6�bR\��R����c�φ������$�Q;
H�J0G �����g�#�����d��:B����5n�:͙{��,��zλz�6�!<��O%'�����o@l�K:�ٺlR�!�.!�t���k���f���9��#3�Y��׃��ۃ�t���g���Oc�ure�w��F�a�*��!q~�O�z�s��r��FQ�w�$~�[�IAf��@�㔴�`�a�.���g��[��7X�wu��5�jP�Gy�O*j�Q��`=0)0��L&�;�x��-2�:��'F�mU^��1������*)ݔ�*3(+��~��31�$$�6�ve��az���^��ļ��)����wm���;ܯw&O�#D>bG��ڤ��'�&�� H��CIF�);���Q_�Z�<�M'�l0��Uq���5��?*~�K��ޏ�}���A��r�]Ț`=�f���s�=І�_h4�?8g�qP&�`O�ub���'���S�qRB��
�MFoV�-�\�ҍ&xڡ)N%��������0�JKL��MRy,�d�ɭ�S-x`�0R�9�)��!l��*UT0��-2��>6��7�Y�
?�Fz�(H�A�Q�����g�O��GQ���0��cJ�퍔QE�9 BCJ�Zc���-0%�R߰{�N�W.���G�Zv��(�~L9^����a~K�A���fi�[t�YR��,�^�M
�B@�4�־c��i����ɇ~J��Z�N>s����c�Ut�B�>�C�r����j^*�<����OeײRq�q2�����q<������o��Y0`�2d���:������S��r�F�5�7�O��;�ǥ'�7���i|]dɑ���a�0Ǫ�鍱�k-�.fVbl+�l�*b��x<��TH$ij�*�Amy$��n��d�5#Ľ��Q*2��~M&�I���LfJ*K����%�x���i�a0�s-KO>�	� ��Kxk�~������	�~rI$�I�*��Q�������p��Xy����$!�( .��4A�C#��?cxKa��w*���UQ�BR*G�Fd���PR,��Y�a)�����T�EIPT�EIHRPQAE�J,�QRJ=R2AEAE�E�Y!EE�QdE��E�QIY!EHQd�E!EAE�a�#"REE	EEDQDQ`�T�)&*��0d�20Y��(��,Qe�#R�YE�-(�,P�R2(�X��,Qe(�X�ưj��,Qh�E��P�E,2�dQh�vF(X��b�F��3�J��ʵ*���F��(��(�����R0��*Qb�(X��,Qh�#"�E�,QeQe(��b����)E�-(��)(�E�,T���-(���,Qb�(�E�QE�,RKE�-(��(��YI,Qe(��YE�Qe$�E�,��Qb�(�E���,��,��(��YasYE�,��*Qb�(�E���,��Qb�(��(�I:ɂ�X��,QR�YI,��,Qe(�B�QE$��,��(��,QeRK(��YR�`�`ă#`�R�K*X�����,��,QeQe(����,QeYE�,��Qb�YB�(��(��(��(҄�E���X��,��$�E�,Qe(�����b����$��c$�J��T�R�,��X��X�YK
T��X��YK)b�(�(�K�J)b�R�,�YE���R�(��YKK)b�Qb�)e,��QD�K)b�)b�)b�)E�X���ZX����Q�L��)ie-,R���*RKK�ZZ,R�%�X��ZZ,R�YD�K(�Z,R�b�X���)QK�Qd��%��)d��Y)E,��K�Q,R�K�R�)(�R�,�K�R�,R�K���Y)TK�K%,R�,��JJX���b�K�R�,��J�X��H�Qiib�JU,�R���ZX�R�JX��%��R�K�UU���U��b�U%X�%X�d�d�*�TUU��U��U��T�d�d���V*�UVJ�d�*�V*�V*��U��T�d�Ub�*�-Z%��U���J�D�UV*� ��V�	X	X		X	 H!,Q`��R,�(�I)	H��T&I%"Ē�I%"Ȓ�bE"��"�(��)R)"�JEH)��H�@H�@H���`'�k�(��_�.�4%	���ޟ�~�( ,����F
 ����RW����_���������w�N�����1?3��_��2��������?��O���3�Hf�ߧ)BM��o��zgg�(����H~�����9�ҟ������~
G����T~Q?���9���������������✓��I$G�Q���Y@���x����`�����߸C�I���B����4�Q��O�~g��O�~G�~�� 9�������!S�s�(���BHJ����҇�[��h!@j؟�4?�������M��"�4~�k|tn�����3W�0E�S�,����x��LoE0U@ʊ�@�P[,hW�E@K�?%Iu`D��D&�t*kL�������?��C������~C��Qe	��Z*�-HOhI�UH���
#/�?֛�!��[�hN?�/_���@�w�?�N�)�{a�S5����jj�����sO����aAQ-?s@r�k�?ؿ����<�:���?��?����k��!�����������C�D�� ���~������_�����D�1��I���
*�~���:���e��������;�gO�!��K�肠�'�?�QU�~����������E]���2����&��i<m&�Q�?�?�@��e���$!�q�Io瀏�[訂F��d7�覈�'c����J!�������	�˼Q�l���k����b	ȼ�àUTJW ���I	������Z��
*�/�e�"������C�~�X������n��~��ҟ����=�g�u?��~���������$D���G�w��q��O&UQ?AB��~B���Ƃ�O�_�(���i���6o���Gh������p~����q���+��a�C�s�G �1�0Yb���n���-"������ �_/~]Ж�������UD�q?P���h�#T��?K���
 ��~��<�??�����,�楯��޻<H�y��c�o叢?�?���+�G�RJ?����"m?`���:O��pP��a*���K�������:�0���������R�#�'?w����H�
��
 